MPQ    �=4    h�  h                                                                                 �W=T�(���C����K�rŽF��4;&�b+��"�eڂ�L<���g]�{�v�f�0!{��Xy�ELce �*^��"�-*�j!�ȴ���0�z���לt�}�n�lL0��S\��Q���玀cQu��Yʚo���K������7��.�����L�q߾$���}�P6p� u�¯U��Hړ��,g�O��فβD�X�TF[��S���J��9��ɞ	D�E����uF!%��LQ�,b�m��J�0`�m�Xe�(O�+��m�ߨA�Zw���F�T�;�dt���L��fE� ��v�Ep,a����͝6H��<MZH'p�(j�
E��
*J*�����iV-��F�
�'�ț�ˍ�� �q�9����Hf��P\]��|4�s�`��b�Ov(�7h1�n�@�0S�C=�}>� ��w�%Bp[�.�Sh�f
jǠP���9��Wi04y>Aũ�����d/��.�Žٍ�F<.��.{���z�L*�	�}9��N7O�eq����D	�A���IB�mTfA�Z��U��Co�O���C�U5�vߗ�`/Ζ��A&�Qm�]�t����T�'G���#�ZrqA�09	�f
?��Y]L�� �
1����v	������wT�VR��j$]s�k�X��cC{�����l���v`x;�b>V��&ȱQ(��N;.>�P�l£�����<"gz�`6�set�a�NU�D��ӱ��s�,�6*m��B�kʄY��wqb�S�ӛ�.T�`���8͒:.���ܦ����Z�Oa��6��l+p3�㈧:?»��<CL��4��-�&ɐ^Yղu�0�M��QRV�\O�#O"_r+�f�zu@G8���*�&���ϊ�a�;pX���c,��=�H��Ի=\=����$2�|a�D0
1�A%Mo���u=ڴ�u���h4M��'���]P�R�d�����%����j"9;�fHi�(�+p�^Iϵ /d�����iu@�n+4��DCT�:���6'	��%IU=�4Ͳd��ʟ%S�B���o�8)]*Y��(\����-�u�ޔ��' �W�_�6��u����k�L�ɞÖɀԕE6,�Q9�T<����Y�*튌Q�͊�
�R.��`�z�d9���"z�X�S��ptU�=�}M�~��|��%�v�����}�J��C�&��1�n,�U�S{�n?چ�؛������bdvɧbܣ*zy��vFb�5��{������lp�FrU�%���lc�����N߾m�m�_��-�a�w��F����~C���^����=D� �<�):�	RЗ���=��?c�=6�O�p�{�HrQ�Ju+��U��&��&+7��4v����_�=2Omi
|\�刴w��6(7Yi%U� ���S�tz�*�"l�!�_�ah;��k��*�H1/x �n�"��?�(Wq`_��5TG�~����fX0\��"�V'�r+���~4�J��e�(�A=LY]�y����K��n��D��7����.{bE� ����v����j�S��I�hXvJb��D5n�90� ��F�� +�����Dd�1|�|lK�5�3�Yf��+ݪ�H�@��=m�:�ct�숊�0 ��O���!t�q0����>
#F�����{��װ.)��4�k?<B5g�C��񢺍2<��~��� �+;{�[L\����[���V_�գ��D��]���	���.��n���T�]�aS�v�HD~%ǫ�nW�랳�(���1��7��t���r�q�f�̡���qS�7͸��|����0�������|5��ѧ�u�h1^
�����'E++�h��v~V�\2�d��6nӅp�(IV�Y�LX��J�b	�M��A��ˈ#s[ŋy�BW�X7�'Z�k�O���M̸��46�tX΅a���=G_��{.cf�lb�4�TF�:�yw�a��ʋ$�#�"�F�:��|E,�oܽ_K��N�76XĨw0��24%��]����2�F2��c�h���'� 7@(|Dh�g�0����Qη�m�ԕ�)t5��m�\T�+jG���#��r�J0NS�
����ԯY���h����v~�Es@��U�D��m���5iv�t�!��f	�)-?[E�G�ԞN���{��/,	ئ�V��G*J�OX�����$���`��_��1o�+@=~�V��=�>k�i�緫��{+��FL�q��RS7���1�ƬK��*Zv�$�{w�t�>��:L:"\�h�y�Z�
�k�mʉ�	5������B.�	���c�f,�\��>��̩HI$����FT���<�z�Є�ςJ�8�?d�����o�}���(�"��Y��7���H�E=n��Y7�%�n}r���ȊA�;�{d�O�f	+3��7"�h��~B���y58��6\-
�Zr��rb� �jے��QÃک$��힐�Wh�jc����"���sȶ��F)/���m���ؠ�o'w�>�dZ|��0�Q��VF�
��L;�&�4��2�@�J�����+�鲘[63��ȢQhw�@	�>B뜖�:C?����O�����%�ox�H��Ld:G~�:%T3=V�B=X.R��a��}�w�_q�
�H�"���d~!1W2Z*3��l��?�@1��?r{�3��c�i��Ix��n��%؎\2P�)wÙg1�}U�D�,q���;K�f^�94U��h� i������<Tm/����Z�\c�X��1���X�~A��NP���\��f��(�כ��UXƄH��\<G�ށ�t�3�-d˂��@��as�=��[<�ڜ�yY/2}���l{��]#ʲ�}���J�(J���(��>�� 䞩sK����0��wT%��Y4E�Ŷ����C[����e�e��㨪����W�o�<�>���
tvIȎ��\z�Z�?U���}�� ,~�771�X�c�K��E�֦�vr���Z�KVi���?=��B��_��l"8j	臂�B��J!����y+	�r��h�x!ăz
�u-A~	Ƀi0�â"Vئ ��O�?��#	9�OQNuT`�����n��fYR���r����D��Bi�+Z6�ڜ�`����k�:�y�xxJkP>.`R¡��⨡�d����-.��w�捥�y������W��U&�J�dF漏c�>A��qP�T�{��ѹ�2�M)ty��g�D7C����5�P4��(c2x*�*�ݮ��y��]�B��#�M@�`�����i/����p<�B����|�P�Ij�e�W�6�@��
��L?�a?vo5[Uj���(&�( �h|J&��q��Q�)S`6k�ޛ}�v���8�髓W�&m�֭%Rl�����^H!�A)=��H�e�Aʸ7��v� $C�����؃�B��  �u��he�-��<��)�#�8�¶���N3WWi� Ki�M҉��$��jWD"�$D����a)*�J^T�8�i�����*�)�W˄?��!�?��s���fe��� ����&�Gx���[�(-�}bɆ����ƻc�n�����{�,��|7��z�![�t����ͩ���8����װ+�\�F'0�ѻ�=�>[�N?���1�f�W�8�t�݋3R�܏��d^.u����x����v��éZy����T,ʛRP��j�~���
:�chP{��T�J�̈=4�`�kb�sG��
���`��W>����Ǆ�|�Q�`g�cW6i�(t)����
NP���A�ӝ�C,)��*�7HB�����5w��S����l�`W�M8�-=:��\�tĉ�.J��u����^��p�F��-�?=���jL�K�UI�&�kY0!�uXj.���/�-zS\�k<O��+��rz�ٯ8y�4E��aŪYna �0p��+���5��!Hh�X���1���k�$m��|��h�? �1'1M*yp�:�d�/:����$4��9'v�FXR����<q�}��:79v�H
��&�[^� �T1��0��G�I��;T���Çm	&��%�[�O������zE\��^�6��3E�*v����.��cl¨qru�����B ˀ�Z�#6S��s�k�̺�D����a��<+,�0ͮO���,�_��	O�lO���H�-U�䛦$�����V��������1��0�M�PH�9�I�=�_v���
ڸ��MC��۟��HnK���5	_"����;q��ϻ�d�>�bW��z�߼�iM�Шϋ��;��PB]p�?r�R�%ƵU����f�ZN�g>�ȼE��w|>,w1�Fr]��T�K܉��^�R1���~k<�_�:VR��P�ρ⇩�c�|���$�p�e�H�raJ�o	��v�v���B�&&A���Z�A],�X�O��%��\"@����6#wiq�-�����J��T�*vLrl��5_�n�;�b �!�H�� Q�" ��,q��_���>�y�^zX�q��=�&'���_Nv4��Ɍ��<�^RA�As]����/�
��I�I�
D#�7s>��/�b�7A F����g�G�í.mI!6X���Sn5��0��Y�*�i��|������|d<US您7��5�1�t�9¦y��#)Y��d��| :'���U�KdD��J�a�r!�A�0Z�1�97�Fx�W&�{��+a�m�v�(�<ݙQ�>������������|��h#��
�\�!��N���͒���&���y]���D����L���q������S���(�~ J���5#�DĖ���<�k���t��r~�@���ܽ$�]���2��L ����ɀ��>��5�h������^�6��uP����+!�ɇck�V������6�n�?���B���3Ls��Jv[	b�#o�*L͗f�KsVJ���l���XR@ZW�&*�ک�2+�d�v6�����D��xT.��_��.>��l�����+�F�U@y� �>�$ؠ0"vg�:߯�|�WowP�K��&����X��0�:2���|�k�6�ؐ���!��3�h�[{�Bֻ7��-��D�괜���~Z�Q)��mp;��D���}����BT�wG�|�#�1rAq0	E$�?�
�H�װ:Y��h>�j�(O~�n@p��_�snޛ���ty���a�A)��SE�O�ԹM�ҍ����u,DE�������J��H����\�v�W�:f1�P�@�n�8��V�q!Z\ɋ����2$��V�����hLJ\��M������dج6ʪ����+s�WR��Vr�5U�"�$�4G.�u�1��!�m�g5	p�8v���F.]^�K��c�������~ ���$#�1�A���]d��5����Ņ@����'Gx�
5V����}2x��-�RBH�^8�EM��=����nnx��+��E��;��X��Rjf䴙�
�Y���~=�̱�46͇��\HLWZ��r=�T���m�C)���t��Lh����h7��j�i]��߹���Q/FF$ŕ�QÈ�G�#Ko���>���|8����2oVA<ωS͋���4��t2��Jh䭌+���<[1_ͪ#N^h2��@$�#BfN�$�����r��=��n3xQ��g=MG����RTnD5��+.MS�a��V}C�&z5�
U�p"���d�3�WͳP3�P^�l@�D��}�͠E�i��x��6��}�����Pcl�ô0j['�t��,��{��z+a�9i�yU��������;����<O��/z��Z�	p������򍐁�3��A�4�P4� �WH�f���(}�7�	��Y��_���_'\׷M�|^~ 7-:��ˆ���D����uw� �t�2ؿ��wfj����-�}�����(���#�+>=p� �#hsf�A�Q�l�R���?��4�zk���T�߹��씀�p�,��c���E��� ^��>
�%��I�p�'N��վ�Uq��� ���~��{�k,�Ȉ3K˪y�Q'�vMP����[��̅^�EH�t�l= �j�����}��@໷@��t<����Π#�2x<w�z�
�-dKɾ
��^kuVӂ���6w����#8��Y�0NP�+��:2�	�f  �����JD�'B�S�Z*�������k 9ݺ�aixHPY�BR=������&	�'	.����Aj�4^���-�WiX&[�=dY��*�><��q����6I�aPLG�2t��t���g*$�C��5��g�P��(~g�*��݉k�y������O����`v��)��/����m��<�0��S�	���Ij�e�b����
�%�
�6�Lz��?��90�cj�}�(�� �^K��0�L�!Q .U`���ޖ|hvi�8�7y��8u�qֈ�f=+�l�����(�!1Kw=r�Ẁk7�3���Qǹ$H]l4���fB< �j_���ڔ���R)&I�8�vж��hN�d����;�q�ȷ����b캚CD�K��o���[��٤e����f���`�����%i��@:
��-۰C{�lR]e��T�h�k��[X&(��k��[ЋL��(Ն�P_�@��Xp�{$��ּn��z=|R��z;3��O����)0�]r
�3�O�n1���܈a`��L6=�*�ى��苀�f�=���K���ic3m���0]R^	���8n�F�ov��ީ��Ň߇TG�hR˭j�����/����{�O�ʥVM��ց`��b4�R��}��1��:9>�6��"gk�7�Q�egp�6D�<td�V̗�cNK<Y���U�I�,Dw�*c�BmѸ�ϪLw��S�叢�q`�/8�g:$���b���͘��m�޳��jp�&�ӽ?�no�NBL����	&�γY��u�OIO-�`��\�*)OX�#+:�z+��84��`�c�MŅH�a[|p�O��ͺ�X�NH#]��s
&|����$�k}|Q:e�:0�1�@!M�s@�U�3ڪ�<�4ß�'�WS�BRz��^����y��^[��*�9��H�\�!��^�y� �eݓ0#_�_�:�$Au�U�T���־��	��%�l��j��Zf\�U�#ɡ����.��*ѯ �U��1a��#3u��F� �^1�U��6�e��.�#k��qǿ����w�T�,+/��J�X��E��F���#Ŋ@�������ך���0���
��Ҕ�3ӨM�B��t���خsv�5seA��C�Z��'�pn�p�����"����Պ��d���b��|z��U�쬌�kS�����ږlژ��p#f!rK��%�����߃���N�0�#���Z�����w��YFM�~����$|$^z�-��D��|��<ٵ�:��R�	��
�u�D�c����cupUo�H��SJk�C��j��X���2��&!k���(������s:PO�N�6	\]����_+6i�-�v
�b	jO�*Q��l0�_%��;�"q�|�zH�dU 5S<"�e@�� "q�_]�kc��t|D��dX��T�X��'�s��:�43a�>��ʴ�A�V�]xX��Jp_�A%�$'�D^�47���P�b�w< #U���3��!)�	c"I\�eX������n��f0X���E�i��ν����dטb�}_/"X�5��ďx'�!6���S����z
���P:��U�bB��f�������<ɺ!�0��R�4�/FodZ� {:i	צ�-�H1���y<xԾ9���X���
��2�	�����������@��K���ZT��:{�]w�Y�}�F6C���3VX����S7�>\t~����3!
͖���ɗB�學;t1חr�h������ٿ���-5���`�>���!��H�5�a���y��H�^��DdD���J+<�r���Vv���ھ����!n�ڡ�[���4L�]�J�nb�r��ev�L�sQ�l�F��uXmkZҠE�Ω�g���hP6�4��; �oӅIJ_���.�Ql�>Ċs�F��Wy-���u�$�=?"�:���|��yo�K}�ښ�X:j�0*�2*��W��q�h/���:$hIW��]I_76�?ħD�K��K!�y�WQ��+m+�_����� �T�vG+p(#��-r���0�V�
�R�����Y'fBh�3t�Z�~AJ@+��zJq�vc��}t���\�)�WLEew���l���Y��m�,ґL+��췽JS�YV4����۸�c�1���@RO�3��VPdE�k���筼'�1[�mL�f��H�'J���-N�Q��� ���~����t���0~*"M_��Ҹ�R`�aP�m�eC	�8��Vs���g.gН���c̲׿u/Ŏ�&P���$�.�<�Nٸ���|1��#F�@J����W�b�ϥ놫|�[������"Z�m�ؒ�GlE�K��x�
�[�Mns����E� !|;J՗E�uf�^�E�����~8Ħ�/TT�B��\c�zZh&ZrMٴ��|�� ��_�ҧbq�;c'hR$NjYZ�n��N�y�쑒F{nެ8x���>C�oΌ>��|s�ԇ VV<����m\��F�4�"�2�-]JC:=�f.^�[,��~h���@?�0B����$��,漠��>���d�x��6�G�)�mrPT�k�x:0.H5�a5�}��@�D
��P"vK�d�emWh-�3��˂]�0@�o�4�9q0��{G&iZ�x&�������P��ϻ��X��O~5,��n�qʇ\��9�X(Uh�*�9*b�1���<���/�4<��ZD��ik�02i�$	��A �OP��&�R!�fQ��(8��$k�����:VY-�\rH�w�[Z�-�����y�W5A��9�($c���o*23R�2��5�ʨ�}}���(�(�PĦ�>�� Z�
s��8�̏K�-���z�~4{L����,����T&ڔ������>G���ڤ�r=���
*��F�B`��P�UL�C�� 9;�~�M|�e@؃��K�u���!v(�?�к��nT���[��m���DslX��j��g��ؕ�{�ʷ�n�om7�($
��T�xWJz A@-�i������S�V�~t�=�>����#Se8�2<N+���.$�F�f��A�O�O�_�<DQ�B_ mZ�K�1�5�L��k��ۺ/3:x�D
Pt6�R�����8�	J��2p.�6 ƜfA�����Ǭ�W�h�&6��d� 4��l�>7�5q����$���=��2O��t�|�g�#uC���>�P��N(��^*x���ds�y
��o/����`1'��Dz/���HJ<?̔�x�{B�IŚ�e������6�N
��_L���?F�+�jUQ/(�'� �tB@�
�'�6Q;R`l�Zޑ�8vrg�8{ͫ�9B���cbxxZl��!�t�=-)K̛W�ʮ���,&C$��!ϐ)���RBt�� �JM���0��ɍ���)a��8Mcv��x�N���̃V�"�C�o��nL���cDX���	�Z��ͤ��q�.T.��33�XT�_�R�z��oؗ�ڰ7�j���?eų�O`6JO��<�&h(D�&�B[�t�s톱t�{�~��v�A�1�P�e|mK�z�d��*U&�6�j��u��.X��fJ��� �|�x�ǔ	=�6��-/�&��f�����+��3��֏�$�^���	�W�ᅋv��u���BTb�RF�j�"[�%9���2{�'�� .�=`�)+b�
�� ��5���>�ٹ�}i/��D�-�3g딨6;�t�J1�2��NF�����7��.,_g�*��]BH4X�
i�wB��S��?�l`�P�8Ě:��l�mp��H�� �~����ypd&�ٙ�?3�%b�L=�����b&��8Y�]!u�=Dd �~�Z�!�\ 
�O�R +z�z�l!8��{ (�ۥ�`W6a�f�p)B���2����|H�쓻�����欿�$�`S|����5`�1�oOM��4�pk��%���-4��W'�� N�,R��:����{�^p�[:Q9�oH:�I�b^Z�� `��Kku������=��'�TUs�ֹ��	�ɔ%z(%��@���� �0�z�R�l,��)�|*,���J�8�L��u^��J � S�P�6	l��阈k�p�:��ZT]�F��,�M��E� ���[����݊��	��{�U�5v˳`1�jB��g�������MiT����s�v����ȏ�{�C�$)���Dn�`Ƭ$?�چ�q����E�dǈ�bMM�z�P�' �������I���3jp>�r�y�%|�I�NxМgN���~���	A�47w�F(���ʉܿd^u`a�xb�7��<�+�:VPRar��Ej��߻?c�Z.�`��p�@H��J�X���~ꙓt1��E&�p�E�����q�{O�{���7\�T��HA6'i'�ޅ1J�)���i}*, elk�~_��);�^��hHb/� Puz"�Bչ5qq��V�o'��oBXa�	�s�'
$���U4n���s�*MAN��]39��eh�� ���QD�}�7�9���bVط ��<���=h���x�I��BXG�~���n�{~0�ǣ`P����Θz�Ly`dr���x6c}�5=xĪ1]��ٿi�f�I]����:ݧ��O�Ё���uȄ���!%F0���/��F�p(�5�{U���!&�#�+�14<��4�@� 0O:'�����!�璯��lo�ЇZ�&sժ���]R��������x���:��GSRB����~����Ri��͖�������h|#tLxrt��O��R�"��V�(��ǥ��R��-��1H5�z#�X���9�^7���r��Xr�+W�c�Y��VQH/����ln��9���_L�YKJl:@b�ၤ��7���sL��¡Fs�s�eX��XZMk���ҩ��%��e�6�ĘΖ��*N�d_�T.�T�l���%��F��*y�g]��{$�"l_:�oz|�Bo��XKx�j�H��X���0E�2����2�ׁ��ǐm�����4�hsG�x�
7��]�m�D���ɿt�2Q�	^m�h�z���s	d��TTp�Gƃ�#��r�?0��
�w
�ｍ��Yb��ht��暬~��@�x2���Vi�!�Q*9' �t�~&�W p)>EE ���﫛҃՚��/,���*��qJ���i��B��lIƕ�d1 ��@��D�.7hV�v���Q���e�(u�#��<0L���Cmj��b(�l����µ�(�i�by�+ǜ"m�����=��ܞ�m[��	�	nW���.�c}����c�������/�Z��$Y��7����������킻.4��_�ܝ��@��w-��3�ɸL7���zђTwzE�j���b���nnq���sȻ�l;�ٗ�'f�(�����91�~3������'�\~0FZ��r�������y8���j��ͺ���hm��j�j�I�I���zȇ�FQ#��Ǡ�:;Y�wo�)b>me�|����"�4V7^L�	.��WJ4fq2�'J�\��_l�\�['p��Xh�K�@ZfB\���Eڑg"� xC�'<�6{�xǍ��OKGxf�H>T�o�i�.C7'a�(�}�]?�
K�"Qd/��W�3�ʵ��$T@bgbO�����Vi�iM�Rx�������m��P�Q���%`v��*K�,"\��:�W'�9U#���T�
⊅����}<�M�/T���Z�ĩ$l�K�&��|����A;~PjA%�MWf��t(���?�O���$�hR�\���r����s-�w޼s���~j�β�c���p�j��2�|����PQf�#'�}��1�=(�ۦf�>�' ��s�8��Go��aIܵ-�4>�����THkv˔�@�"���������d����
��ȿ ��]�8�ˉ�U'�*�.t{ ��~�9B���>4�K�9�G�iv����'�ǎ�q5����ݐ5�ls�qjz�9�lS�ĶlM�vГj��⃔Š��xr=vz{��-ҏ�4�hؔ\cVɚX�M��p��#nC�O�sNgӌi���?�Bf����u^�N$D8�B��Z���l浏�Gk�|6��$�x{a�P��?R3���h�B�]|E.��~����������K W_� &`d���`!U>2�rqa(���W�V�B��2*d�t*��g`C�C�ҧ��,�Pek�(�1�*�>�?��yX&��.�i��2�^��`�o��_v�/we��#<=mc��nv��I c%eF����;��b�
��L�_?�7&W�j�DD(W�V �a����Qv�u`nތ�Dvͅ86���ZW��9�>6Z��*l�9���{!罳=�"̶c[�)�Q���$���j2��ɢ�B� QJ?��bڊ\:���Z)��8�o����ND����3�q�{߾��aCf�0[�D���%;���t�
��e����º��U��υ����uM��4�RO>�R�B�b�e�޸���ї+��=(&�Hj��-[�������Ķ�4���q��ь3��C�0|��.z1����D�qBYǓ�V�)� �$�#�\-)��2��B1)={b$��ԧ��}�f�� �InW�C�3�Tp�&r^����D}5�|v���k~���n�T}W�R��j��ȬW�V�46{��[%��n|`�cb*�m^��=�n���$>��E�؋3���H�gf]6�Tt�`��2�NA8ށRIz����,zw�*Y�B#�g�EG�w�8�S�wt��u�`�Ԁ89��:R�H�Ɖ�������.�o9)p����?��=�Lx�Ǥ&\�&���YA, u����|������\;	O�95+u��z�e*8�� ��Tj�;��a�p�pē���9��H�����8/�p懙�$v=|��&�0�r18��M[�L܋��ڠZ��`z49�4'GСI��R0������S-�Q�6jV9'�H�aZ�H0^��s �a�f�s�Uc���v��]�T�p�ִ:)	7�%%5д����P���wb?+��`�$Yj*����u�g�O��u9��L� ��:�KO!6d������k+�ǵ��50ԁ�,a���@�D�=U�� �+]�O����P�Lm����=�����?o,�ܰ��)xMD�h��qp��cv�edp+�6C�L��n�=L�?�]�}K���4�L��� �nd�]*b���zy�2�b���ϋ�?��LGt��܆pYƜrA=�%W�k�X���7p�N�"�������<l���w���F�@�#��Zݻ^p4��cˬ��Z=<��:��R<�?����z�c�����?p��HޕJa���q���#?�h�&���[ŀr{���Ok�v�V\����BW6K�i����쩥D�?`��*��l�vA_[TE;��2h�H� k�`"�P�Քj�qL���u�j�o��Xsˎ�F'�����=4��x�tF����A��]�95쀀��7<{�D�c:7D�[���b�X� w������������Iҩ�X����4UnF'60λt�{>��1 �s[��u�d�)�s-���5�����
���ڴK�
n�58��a:8����{6МP@��ą�!`u0+-��*~,F%����C{p��ל�b��Ԟ�l <����/)L�X�
}h�']�������<�G-L�-ߦ��y���B֣�A�X�0��]-;����z|K���fK���I��Sm�g�4#U~��޼Z�:W�Ɩ�K�M���#`�tgm`r������*̍9 �.tܛ#b�]ʊ���m��Q`�x;�5p�@ѓDN����^
����l�lz+r����3V,,y�P](�ann�-�����E��L�uEJ��}bups��*[�7��sG�>�����.�YX���Z�U'��92��5��6�t���^���T�_|�.�9�lN���b�F�f�y�Aܕo�[$)ش"��:p�D|1�^oH�Ks�֚���X��u0`{e2 ��� 6��$퐞�v
�٦�dMh��sۓ��7,��zSaDTn����o�)Q:e0m�/4��,���js"T�TGa��#��:rR�x0:�%{,
��5�h�Y��3hQ��~�J�@�UD�����,�b�tJ���R=A)��=E�&��
=��h�}q�,�L���K���J	�������t����˼O1[y>@���)
�V�M�u|��/��Mݶ�
l�wwLܓ�>� |f���(z��c£����&0"�=V�e����HֺWm6�	!�	xŖ�$�.��|�c#�k����ؿ̕�D$�%�2���n���f����݂63 ���`����۸�r�����¸l���F2����E��b����Htni�<-��v�a;7�f�;�0fu.��z����~.d/����͸r\�ҹZ^�}r�Vr�V�6�p�ƕ��]WD���Xh��jO�N$������"��FG��b�w�x��t�o�#>HP}|��Խ�V2�d~��64.��2���J�E�ܰUչ["��4Ehc�p@uh�B�"����Ñ�~+��[��~����x��o븈6G���#*�Tˬ��h.>Y�a��}t�!�AD
�&V",YUdj*zW���3����w@�j�!g���1�i�4�x\���E���OP��(��۳��8A,]���hR��9z�EU����o�{���f(�< �/�	��jdZ���߼:�f�����ܥ�GAv� P��H3f��(�bs�Z����D������\�ɰ�m�C�-PFE�ӺM�ҩK��lZH	}�eU2�
����k�ʞ�"}_XSl��(�}K��D>N< �q�s��_��nM��O����s4�O-���P�,D����ѧ�M���Z�Ce*ߨL���
��l�z��x�r�FIUB�iT{ o��~����(����KƧ�h}vމ�Fq�������V#�KF}l�j����G�,��bD�ʥ�e/V��$�Tl�x�P�z�;-��q�o���/��V��X����+��#�A�ʕ�N�W����#��M�f�!�\-����DS�BU�Z������	���k�N��5|x6��P��ZR�?,`>��}-����.�Py�R�݈eU��
�Wڍ�&�Q~d
;Ҽ��S>-aLq����g�V  ���2Kte�$g���C�����@P I�(��e*nL���vy�iJ�ɤ|�隞�u2`����z�*/�����<x�n�$��q�
I{K6e�������,16
p�6L+j�?|�(!�6jX�(� � �6�B��[qQ���`�Y�އ9�v(�n8�������??�*�lU���FD!B'�=�2��я�ʤ5E��C&$�kh�J�ė�B*�� j5�0�W7��@�)�x�8������gN�B�CB����|�9(�<8��k�@D�����(��M@���R��$U#�]S���jL�ͮ�p�QY��mk�݄�e{)�|�l ��^�&��X�[!u۷i<A�g�M��ʑς�l�/�������|���z�'T��vԬ���.�P�$�c�s�������ኽ�=V��:���\,mf�c���/c���B3��q���^���O��+v�g��j�Ÿ�>T�� R<E�jkFF�����Ϻu{�7$ʶ<��)!`���b�)}9g��xq��U�.>���3�w�h@�cV(g�E*6�
Xt��h�N<�ꁭ��z��,���*�E$B�Y焀ELwx��S�����`Cx�8T�:�Э�#�<���јV��J����xp�A��/?)k��L�������&���Y��uD�y�t�2�I�\v(�O)@�+phz<8e����z��վa��p_���\3�iS�HTl}����y��b��$Y�;|"p��+ �1�.M$�ܦ���Pr�;��4t F'��D75R�(���o��ꌿ����9bHpC�N/^jS �W:��[Z�������T��T֯`	��6%�����Ĳˉ����ze���Y��s*�����U��A7�u3z��� �ٓ�F��6����_��kF1G�0}$�,�ԼYH,�ꍮ;����8�ѼH��_E��{��0��U�k��:�A�����C����z�M���%�����?v�-�v7����GC��^�ns:�z4�ut��wq��zuջ�d�RbC^�zT����6C�<��XڧdQ�<�pt�6r� �%2A��������SN�KZ�4ި���bw+�Fޔy�@�5���+^k(��>���9v<*x":)�R�����h�3Xc�U���p�L�H�6�J����L	�	� �]$&�9��$��-pG��~
O�zQQ�e\驴~d!6��iݪ���)�_g'���*�3�l�[_���;�"���uH�$� ��"�K�o��q�Ў�<�M�eݔ���jX�A˩,7' ��ˍu4���	�v�AW�]�Z웸��w/��XDj�7ߴ-�s�b�. 2Ɨ����3U����I��X}%�����n��0��ţ�LY��z�N\�d�#��nD3�<5�d����+Kڏ��E���F��Ck:�ʸ���[з4�kwo��m3!�J�0Ʀ��%+�F���C��{�v)�kO���!�]�<Il�*���i�<��͜-�n�z�Բr[��u���.��+�"�����1�\������]���0o7��t�g`
��S�B�����~l���������$5ɨˮ��ct��Prj���]�&�Ȣq��{������oP��	����d�5K�θ��oۂ^�g�U΅8+�H�O}�V0���܂��n�g���g� ��L߱�Jb�'bPU��r��`�sB�a�Woz��RX��ZC`��q�t�p�оn6�D��L.����� _�V�.�>gl����[
+F�y><��*��$D�"b) :K�_|lD�o�ڌKnZ����Xk|o0{c�2�~?��Z�"ۆ�9HG���K�3hz
$ۮbz7�۽UY^D�/��{Sj�<Q��m\�����i��NӼT���G�
�#��r�Jr0�KE@$)
�WǽC`�Y؋jh��搰L~R@\R:�˦Y_����ċt�>�M��)��6E���%�f�yz��X#+,0:	���ϭJd�L�q����b�啦k1�q�@#�X�$��Va�1F���"�Fj�����$L�F��9Ƀ[���G��K���kI�k7���Q�E�`�!�u"#�� Vظ�s�қEm�	\$������xs.x��7�3c����[/�����н�$��w�-���ɝ6�!z�'���WX�����D��v�)�m�Z���������2��J6�E��)<��,ʻnd������1`Z;Ro{��|�fPդ�Q�o�~)�ݱ@ro�s�T\���Z��r����,⧯������Ҹ�l�Wh�ˎj����m���PyȽy�F]!޽X��3���Do�@�>#[�|$k3�X)�V- ���ϥ�	�4IL�2	��J��K�"E�m�[O���;�hY�@��HBRT����\����V_���*���x=�����iGn?��5*TZ���I&�.9�'aF�}/����
A�z"d���W9Z�3����n]�@ض��������i��gx�G���#'QPO��� ��V(��D,����By�MM9���U�L�ٴ‶��A�J<;� /�$��ZU�c��m���Z�y�(��vA�m7P�,
�Cl�fbNA(i��u�R�EN���,��9\C���h��l�H-5P�7�;��qA҄��@d�d��`$�2D�n�c��Ȇ�����}:���f(QD�z>�� �vKs�P��=�p��^g�+��4L����V��
1�u���.��=��/�~Z��C�˻�>9
;#F�56���VU���yU�u��T� 
�~~�����ش_K7_�=i]v��ﴁ|l]f6���|�����w�l�`�jp!��"� �,y����s�`���9ռ�(�x��@zq��-�;�ɪ�r��ͱV�2u�N�U���#�_�EwgN�h;��+2�u�f��k�`b����?DnB�E�Z}Y��42��Mk�@ �@g�x��#PŲ�R)�;����oŰ�oX.��ƭ,� =)��%WUP�&�c	dE������>(��qԍ"N;��8�Y2��t�%�g��6C�X
�Oq:P�F(�{�*餾��Jhy��h�dog�ߞS�`ba�ӕ�_/m�I��"`<�)��l�I�S�e���2���
KnzLf�A?YS��jf�N(ͣ� w����ĖQ�~f`=eނ�v�"�8�a��Y�Ð��=�)��l�i!��p=^�}�������$4����B�M ǩ/�K<_ڀq�����)8���~��N�!��o���%ߴ�ӮM*즛�D)j��[��k���B��_z��P�8��	&g�0� �k6�O����1��c��X�peV�U@B��̎���&y�6�Wč[<X��}�B��,��j{g�g���B*���|�U,z'�@��7����R��@��}���)����̈́��8�L=1��u�����f����O��ܪ3�|ۏ;B^u�n��A���үv��#�!ws�s~�T�U�R��BjFԬͼΟj_{{�o��t���I`8�b �8�*��y|���>���֎0��#��~�Ng\N6�"�tP$��9N7�ӁD�5��,���*O�iB�ׄ�c4w�S��I�P�_`�;�8od:o`��YC������dB���%�hp����*��?�TR��L��I�\��&��/Y�(�u�j������tj\�g%O�f�+kb�z���8 w�̴��6��C�aG�Jp�����!��ķH\x���X��l�=��$� N|�lH�&��1Mў����ږe��r�4�`�'}�?�SR��J��0��� x��)Q9��mH��t
^kO� ��v��)�K�@���8�A*�T&�֪��	��%���֙ڲF���������=�i���*=ݴ�{0����Z�y'u���DW $�$�A=L6?��Oka�ǫ	��G����a,�iڮ6H���W���y��󳕊��բt������+��V��?-���^�u���M�Iy�`���DA�v}���Ь��C.C����nNW謵�|�T��*j����vPdh�b��z/HP���ү�=����������p���r7$G%� ��X�m{�N��揆D�FO�w�y�F��B�{�"ܐ��^f<���!�h8S<EN�:��R�l����̇��8cޗC�q��pA֘H��JW�&�'zЙD�֨�3�&S(�Vm�脈��*nO��*,�d\I㌴�c6
Ri8�i�bɘz��Vy *��Ila_��D;�b͊��^H�O� ��%"�R�J4q��\����`�'�%N_X����ę�'{������4=��+�L�A_�]d�k���-����DJ�7z����bg�* ��5)����6�uz�IH�QX~tּ�n�݅0DI���z����)}���dC���i{g��+5nF�����h�j�����kuf��E,:���N5e��8F�������;!֜�0a@�� �F�U���w{�eDג=Ȧ������<�pϾ%97��f��bW�H�(���ɲM(>���|�c������}V�и��wb��&]>]�
��k����������M�࿱ES��Я*j�~G����l9�`���G���噇�t��Ir��8Y��,w�d�1��_�15�*�d�$>?�n��5&���	M��
�A^ �
��]�����+�����V�S}��{��=Nn����J���M#L�rJ�x=b+�&�Q_~�mRs=� ²3���UNX�cSZ��9q�?��|4�k�6|4VΧW�[~��R_r�:.�cyl�/���YF��y�V���L�$_�J"��2:&�|��o~�Ki�C�Y��X&m�0�k�2�����B�]����� L���%�h5�X��U>7"2 0�D�圷��e�kQ�{�m\�������)�T�G�~#�t8r,0��7[�m
vD���"Y�uhE�
�b�~�y@o��Zw��Y��>z��Kt����HX)O	0EQV(�@)�����3��,kGY�=W��6J��B?+�'����Q�����1щ�@��v��V�mVѝ��,�^ö�:��9%LQ��4�Z��������Ū��F
���s�����b�"~�M��)����l�MJ~m�	�]�?x���.�����C�c8��aU �`
��{$*��(�B�$�u��c$�B蕂,�ܚa{��N�s���h��DaU�}5���>,���-E_���d�#��k{n_�r�����_W;mf�1Wf+F��1���
��~$�(���.h�\�v�ZT�Qr��˴̜��J?ʃ�K	���'��h��4jE\A��A�:�v�X\5F�j�N���Z�c�o	�j>���|_�)��v�V(k�/���5�4d�(2���J���R��&�[7���h�z@�d�Bͥ<�\h���j����|�G~Hx�����Z�G�ۇ�ahT�H���.4��a���}�c���
��"���d�nWW�S3|�[��)�@�.�:*]:���'i��x�w�z��~�P
���;�юV�q,�TE��H*H�90"dUT�������~���)<vg�/%_��fZ�LQU������`�z�KA�K�P;���>Ŕf��g($Jڛ������ƦM=�p\����c�S�'�-�C��R�̺C��_�5"~�=�[�2����'�ȡd2ʔ��}@��e!(�*3�
4">� F�~s�'ϸ�������f�94�ұ���e�eU�@%��֡��Bf���h�o ��o�׎H
�r?��p����ߢ<�VU�� ��t ��~���S��o%�KR�6���	v��������1�����C���l���j�8�����g���G�9�[qe┥����x�ֱz�Zf-c�����e6}V����ߝ����#���x#N��w�x��սf�"򙻈�K�sD�5�BK��ZX5��.���k�Ro���>x�w�P���R�N[,����ְ.�.�����z��DG�3�W�2�&���d����1�>#��qr��ݯiV����2��|t۝�g1b�C{�Ւ�CtP�d�(Q�*d���ҩy	Pۈ�Y*�E��oP"`
�ӰV|/�O���U�<��ZSg�.I1|�ew%��*ݨ�".N
&LNL�|�?��sPj��C(�bI 2�,_+��MlQ'#�`ؐv�}W�vޠW8ghū5~Gh.��q�dWxl������!�Y=��Hʚ�p���$o�;�L���B�!� �	.�f�)���Ս^4`)M�]8�U��y�sNU!%��B���v�/M�����k�D�A��&8����G����H���D���2k�f����؃����{:�ӛe1L{(��@��} C&�i��P[W[c�_�ņh�g����b��ѝ��t�l|�C�z�jY����"�]�d��t��5 1���ڈ�]k���P=�>ٰ�
��@f����Z�t	�3�@����L^P����S��M,�v�a��|���.6xT�dR2Jnj!�q��(�${��4�l˲���`5Ҍb�Ġ�`���Q���j>��Q����޻P�@=g�v�6�ZPt�W�̞��N2���c��@�,�g�*��B��6����w��yS�B����[`�Y8�p�:�-���ى4��ճ�2�����pP���E�C?^��*�L)0�����&��YRWu�d���jJ;O��\��6O_��+f|qz��8�����K��?���a�O�p�H����<6H�kw���9o�n��-$�ut|X�=�!`h1ImIM�9n��s�����V�4��'v:.RA����K��ꂠ��ǹF9�H�ٜ���^�T3 L�������eоk'��|��T�)�֥�	H��%fW��L�����ʜ�y��,�؎����*�82�6���7�ڜu�46� � �<�;6u�����k|#>�&���ƃ�2�O,2�1���N	��GV��(N�y՜�O�q��S'ס��������pF~�-n����(M���yL�ߵ�vxa,&��g�CI����YNn)�����Z������]���1�Bd3��b9�>z
0W�ݶ�r�g��O�]�+���5p��"r�G�%�Fs�	G��1!N�����+����w��yF�𛄶���+�S^apI�t�L�#W�<`DD:|VR�U`�1��K*Qcٖm��zp�>H/�HJҪ��h��`�9*d&s���������9Ov�o1T\��c��6�Xi��B��������*��lW�_,Z(;��*�C&hHN�� �="���%Ɏq�_�r9&�[w��ؓXM����&p'�%l����4ZI�E� �B�A���]��ш��N\k} D�֩7�����b� �}�P���)�حP�I�=X��KַxTnW�0��T�����}���8*�d����dҋ�'�5)H7�V�9�E���C����gI:Im[�	�R��\��a�
��{4!�0�����F6�a��{�t��0ͦ�:X�8�<�J� ���;�c���pk�(��ec��-���B�8i�s���G����]��H��TMۼ����[Z�zjS��ᯥ=~"��g(Ƃ��6U�^��T��t�>Jr`��G��>���� �i�n�����ր?����5��D��29^�2���I�D+�J��E�V��7�;����un�;����J�v2�L��JXx�b�褌)~�ds8���_�NX��aZ9�L����Q��{6wDx�-��y�Ф�_�a�.`��l�_�đ�@F���y��ٕ��$z/B"X�:o�|���o`!Kd�D��[�X�}�0���2��e�p񁘧�o����n���h�!��h
7��N�D��R�G`�QK7hm�Cf����_O�T@��G2�#�{�rc��0k��v��
�PϽ�w�YN�Th����4�~�@ҫҳ/�U2�޽����te7�C��)�E)EI�[�Q�o���f,�t�SA��ZJ����	�B+v�X?��\321�o@YM�CxV �����&�����x���(}zL�{�/�T�N�x��+}��R��!�pM
�{�(�+?"ٖ	��Ƹ*ĺ��m�:�	ҶYڙu����..�<��TcS!¿�n��;S��Ff$$ň�#M���t��m�])^�� ��<o�܉�Ϭ\��c'����8�Q��jŒ@u�E:&P�L�b-�nZ��M�-ȧX;�}=��Q�f�S�l<O��#q~D������^\�xZ�A>r_�@�-է��O���A�n�a��/"hم�j��l��߹ug���^�F��scǠ�}-�;�o���>���|���Ԏ�aV#"�uo�C�4��2���J��{��dn&�[�E��h���@��BH��7	��SS���Ƈ�C
���x�T��	��Gd����vT�֬c�./�a�m}}�P"nQ
7�"��^dA�Wom3w>6�$�@N�����،���0�i9l�x-�_�u-��5IPŜ��V>�L,1;,==�x8C�9�dSU���C�vg����X<�Z�/�����Z������.�o儥U��A'J�P֗��9>Lf_(��S�����;+tƁ��T�;\y���^"�-�rR�m˅�����:�OI�|��V"92�uB���ȼU���U}����(�1���>_(7 ��s�&�3-��t�Eܡ�4�D(������������"�ݒ���������yL�����
��Xȫ���ɚ����U������ @a~�4��)f�*�Kmy�3ʁvo����,�����4�g��|8�l�PGjf���~XĢ�����VB������x�I+zg1->g�� r�� �`V�J����\�#��t;�Nr�c�U�j��f≴����kD�~�B���Z31��X��Sw�k�:��)pxg�P��R�Ҋ�.Tܰ��K.��Q�c4Ɉ�li�NlWK5�&}�Od��ּ�3�>Y�qͅ���b�q��.8�2��]t6�g��Cv^]�6�PQ�>( FM*ߵoݫz;yD󡈚d������m�`��q��6�/c3����j<)fI����b�:I��ie2y��E���\�
J�L�5u?M��gjR�(CA� M�o���n��Qb�'`s�	�x�v9?�8"��P}�,֪��&�l&T��!S#�=԰i�"Ԅ���s�$������68B;$ =�0؁
|�vw�9�,)�ȿ8T❶t��N�@�t;��Ypߪ�r��֮�\D_9��Z�!:q~����h������ ����f���ae7b	�>������Nׂeʲ�.=N�x��&/
����[r~���o��sMĢ����s�]g����/��|�Q�z<��q��]���g������
�Ht�W��.�=�Q�����-�.f�����3��/V'3%���^+5�0�5�� v�����e��T��aR��%j���C���O{�?'��B�ZG`P�	b´�"�)�Z�&8�>����DUŘ������gR�g6f�Dtƪd�9]4N-�9���D����,��/*E��B��1 awIVS����`t#T8��:�� �oo
�'f=��s��)p���`X
?��L���Ld�����k&��VY���uu~��U}徱*�#\'FO�z+a��zM�8����X�ŧ�a�ٛp0���	�z�dH��z�������@}$
�|����0�1�<MG�����ڌ���[�4%��'���5��R��>�V��f����@ϝ�i�9�HA�� U^!z3 j�ҳ~�AQL�F����v�T\��֠>�	�j%!���  �<ͭ�wΡ+IU�sw���9*�O��������\>u���q�� Zt�7�g6�k�����k�̥ǡ�V����m,��{�,Ln���S��)�n���Ϣ*��86~�<���QRu�+Ρ�H��BMM�����f�zJevsE��M��"��Cd�h�	n�D�+�lF�>������c��k�dN�.b��z�7��N����w�ڸ|)�m��p�ur-��%��U�DUУ|N����E����KB9�`wyvqFoN���Ǹ��^\�	��X�ޕ�<{Z:|U�R�^˔l߰��աcԵӲ'y/p�I�HJ��JM�����ϙ� ���@�&�A��^���mO�h!�3\�7/�O�P6 _�i�G��h���L�i*s��l��_�F�;�B$����H	P ���"u�d� ~�q8a���&�V^��ۂX����Ӹ'qv��\M�4��Q�����XLAw�]�|2�� g�#��F��D�<�7��sԶ�b�� c��k������+�0I��@XN�;ֲ$7n�V0�V���6���6����s��dy�X�_I�D~J5�i��1���A�� �E��v�2%�ߩ�:�����n$�����m��^2!L��0�����F��0t�{ܣ׈B^�j��X�<�]�ɒ�z����֜~ϔ��j��" �3~����3;��.Mt��L8���]�Z���D��Æ�^�x���5C]Sٲگ 1(~�]�F��K\��o_ɹt"�/ht�Sr��?��Tz�y�>��v�m���`����Z���d�5�֖��h�@�h^��f�����+��R����V����<��s�(n�չ� �ɽ17�L0&?Jӗ�b�뚤�r����s3m��h�USXR�Z�?|'?٩%G���4�6rt6�]\?�ѓ��_h�.;.l:`y�,��F�QyO�X�[xm$��"�ʼ:�~�|o��/K_L!��/X���0�ۥ2��y+�ӽ�
���MC�\f�h��M����7?��*�D@3����[>Q��m������0qߥ�T{�G��V#��&r���0&ai���
l}E��3�Y��h{��&R~cP�@�u�#�ЩFޘ� N+�t����>q_)�"E�n�v���a���,��5����Ju
a��]����L�7��1G�@�k۾��Vr�_w�ϋAD���ٶS���c�#L�F��*Ül1
	�G�����?��yO��.���"4�E�Q1��2�#�Cm��i	0�u:���4|.�$=�ha[cn���W�&���́�$`���̥��X4�R���x�n�"�ɚ�4�đ>�G��^_���Sh��~���ƒ�DE���ڪh��cnU�N�>\�b�];���'l8f��*����@p�~$��Q��ͤ�\�ZJ��r:��B��������6���됝��h���j;�d�M͹�"nȎ�F_��Θ��d^d�3�o��b>�;�|�]s�)rVc����¥��4��v2z��Je�k��5a��\[�}:hO�@���Bè��I��/z�'*��Զ�ʑxn�D�$��G�tA�UT���2�.*!�aWO}`]�7&
�r"���dV3W
��3r���"@	u�8SS�3͝�iti�xȠP�pe�4m�P���q�����q+�,IEi�H�>��9�ƂU����ۨ��o�����<�mJ/[4m��
ZfGL��^��2u��8��0_Abh4Pq}��4��fs5(��Q���\�����\	���\L1�Yz�}�8-<�I���f�9������}��7��QQ�2U�L�f��fxʊ��}˧�X��("X{� p>�a� �D�s#�Ϯ�b�OK���`�4��}Ek����俔=�����[�`�/�&�Iۻ͎;
Lq��fFj��l�2�Und��U� ���~ԏ�	�����K�6ȧ�*�vJ�p�2^.~����Z����7�Bl���j��)������{��} ��Q3e�J��@�x�ܬz�'�--��[�X؛g\V�s�_6��N#�y���NM[ ��p��F�}f���q5��(D��BA�TZM ��������k��a�Q��x"�BPO�R��:̙k�i�հd�y.�=ƾ��Q���iG[W�W�&XYd�/ �g�@>A�q(m�S5����?2q�ntQ�gg�qCq��`H�P ;(;[�*Zn�݆By���5�8�!Ԟ%��`��a��6n/�6,�j�<d4%��]CI�,{e����`�����
�g�L�?��c{�jw�(�?u h�W"rĵI�'Q��`H��s�v��@8�[ګk���Nօ9��&l�*#�.!�=�ŵ�=�Sʐ3M�N�-$�gq:/�B�*� �(7؜�V�񀤍�	)��58�Զo�N�-/-W����%~D��K��WllD�P4��8�|�9W�"G��מ���������\;������R����2�e甉�T����s"�&�ʪ��}[���U{������ϩ;%�Xx\�S����9�|��z�-�L:/Ԙ/�ǚ+k�������VЈp��==���&�p��&uf���uS���;3*)���q�^�8�k���?v��.�2\�Ť�T��R(�ij�ެ~t�;{�׵�"�U�ʚ`kf.b��t���dR�����>�K֟
�T��Ϫrg�'�6A*�t8��7vN(޶��g�fRT,��*�S�Bj%G�l~�w�T*S�l�a��`/G�8��v:�
��c����������K�6J�p�<��{��?���jL�8T�-�&�DY�u0�Ǳ`St9\b��O��g+\Rz�$y8Qe'iNy8�łPa��2p�h��0�դ�H@끻0\�e�κ�$E��|�"�� n1�+M����B�f#��4`A�'Nv�0cR���{��聥^�x��}9"9N�`H�W����^|�� �Z����\��!�$��LNT�DR֛�	��{%�.�'O��#��R�Yf*��,���*NO��@��ӗ�u��`��n ��(�2��6+2��K#�k��U�o��|[�Ԩv�,h�Ю'�^����o��Dp��o$o���s8���Oų�mf�4��uɘc�2����M�_��t����vn�k���܃C�ԟ��[n�m��fղ��G�����2է)zdig�b/ �z�_U��{��}���U����(�p�f�r��%�̨����>��N�/8�x�wTw�$uFJ���,b�a��^W8�*L�����<��:�NbR��攧#1���*c��u���pr3�He��J�0�����o�ow&��g������0�	Ol�>�\����*�6�3�iI����h�˃Ǩp*N�l�0=_bS�;�⹊�D�Hď� ��"��o��R>qs������Q�I�6M�Xß����'����7�v4�ڌ{sX���Apl�]����ꞥ9!��D��87K+&Ϸ�bx� �������@��+I�?�X�GC֭�5n`.0ut����s�κ�P�B�d���Z����y5����L(��~�X���1r<�����:��~�;��#\�WUV�9	�!�S�02�]��F�Z�/dd{����u{�E�䓒<<�>	���������̜�	G�f豲�N)�n���4�<��v��]�����q���V�]t2����0��}���*��;�S�»��D+~��x���^�-���e����ʲht�drV^p�ɂ�̴� �5��
���$�e�[˦�u����J�5��$Ѻɱ��	�^��Z��h�,�+���;��Vs�w6��3n��!�[�(��[1LK�AJN�b�=�Z�>�rs.����@���\X*�Z/�o>�`\��<��6mĐθ�㐌���_��-.��lu�l���6Fz��y�e�>$�	�"N�3:���|X1�oOeKZ2ښj�XW�?0�Cz2�l<�T���v��~:����6�hf���7�����D{t�]�V��Q�mH�f�#*�U2���8T�Y�Gh�M#���r$�0�R���
�����Y�(�hJY�|8~���@H���77AKA_�ss,��DtQ��9N�)`E��ԑ�]�eD���*�,/����ɯwJбRs�2�x߿�Nz5�͹1���@��!�	�V̈́D2�N�\��
h��.ri��c!L"1��%�.��*z����}����B��I�������"���eĸM`���qm}�h	H�z����b.�w��# c�-���|��D�̼��$��?�k��5׳��%��ǂ�)2����@b��i�Y�c�U����S��*#0�64�E��I�ey��nP�v��g;� ���f�������ܻ~$������_��\ ��Z�,r��}���f���L��$뵐X��h��j�m(k-���g�)�LF��n�)_��K�oz��>���|D����V�f�+P��x�4��)2�Z�J@�'�\�[	?���(Hh
��@���B>Zc����+�­��ڶX�Vx)x��?�GZqj�TF��� |.%�ya�P�}��R�b
-LG"s+kd�EJW� h3m8_��N+@����3Α*�x�Qi���xce��k������P;tÌR�B���L�(,�mɄ�w19�9AI�U��2��-j�l�9����<'� /�����Z��Y�8"���e���B�A��P�u�/��f���(U�ӛ�H�1�{�7���)�\����T����s-�/弣7p��� ��'V�єO�L�}2���O�v���B�}��Q�#z(�����!�>�� w�ps>_�)L6�*����	4��}�x*��v��q�ɔX���(�;<w�jo�߯e���>
� ��!����^p����UII�񐕈 vP�~�
d��ؠ6AK�=�)��v%��m�=�p5��5]�����y�l��j\�����P��^\�LD��֬��V�x�6z]>�-��ɖ�x�60pV���6��t�#�1=`N(�L��t��2fط�̻y�|X�D�p�B�70Z�q��Q���{k�H庬lsxݭjP1��R����<���ð��.�A���f������WA�&3��d1�=��7>I�q�t��(��2$3�2L�t��'g��Cl䠒�z�P�}{(V�%*�FQ�a*Oy��+��ك{�����`Nĵ�WC/YZ��E�5<�"u�+�SX�GIB�e����{���M
��*LR�?����jҘ�(�^ ��g�+ӵ$�Q�Ϲ`����n�|v��U8������y��`ͷ%;l\!����!	l=J���XL���]�)>H$ �����@_B�^, ��AطX��l^���)��8�[��jx�Nf���w��~[ߠc®���쒜�D��g��F���.��,�=�w�����R���RZ�W1�e�ش�ʰ�[�D�Ee��,��s	��n�:&���C��[�$l���熮��!b֝��SnѮ��m|*�z?��'{n�Ӌ��5~�7�FC���Wq�9�֊$|%=�	��a`��cufz��kֿ��O43EM���^�B\��Jn��qv��*���X�_mT��R��9j�O�����1�{Ǐ��}�׈�lS`�`�b���ٱ��	�\7*>����������ꏹgH��6�t<�_�o2�N#,�t��!9,x?*;'�BEh���^w��S�-Ţ��O`��8�A�:�(��jQ��塿�]��~?���ip�㖄?�:�_��L�쿤���&��mYc��u�g!X.���\\��cO0A�+W�Lz��8J�8���7��]?�a3N�pfL��uY�0��H�Z��K��O��TL$��`|)���0�1Z;M����-
Sڂ�=��74�!�'�]�+>&RR�6B�������V�X)9�wHwqx��K^�$T }kR��t�7������-C[T��֖ 8	Y%�ʧ�B&��2���-:��+c������I*�
k�gV�	�Q���u[���� �{��-�s6�!�սk�~MǗ{��W�h��,�}�"Ы�_���x�M�_D��{z��R�Z�r���
�q���=��~Kךg:MfQ\�L�����vvi��=�sИ/mC�+����n�
b��-|	��6��nB�b|d���b�8�z��L��F[�C(���S��n�D��pip���r#r�%y�k������N�����gߨ2Fo��wo�F%j�gZ��� �^R�ޑ�_��Ts0<��#:rh*R^б��e���c�ST����p-=�H�<
JCx�����0���
��&�:|���=��v�KO�����\5����6�(Ui�PυN��暦B�*)e�l�x_�d;Ƣ�TEH:o �"k'նG�q�a��C�O�LT͖�7�X~�r�0��'gw��m?4���v���PAˁB]Pމ�"�������D6i.7�����b�� � ��u�����ᑶI4�X� c֨�Pnh˦00���s���pΕ@u���d�5��U�a��i5Z��g�����Z��2�l9h�oD�Ս�:ZQ��:(t�>�3��\� �!�%�0��?�l�FGG���{b�~�$� ����o�<P�L��^�0l�朴c���W�������O�Ϝ��Y��wФH���ت?i]O*f�W�"�Z�x�5.C#�TS�x~��N���������Ah�o�E�V�t	0}r�ܬ��Ђ��V�з��ի�~�����ނZ+5��b��ݮ�v�o^����W�u�l+�އ���VN#G��8�쩨�n�i塶�g���SLf��J�6�b�iϤ=H6��X�s)�V�����hXE��Z�t��������̓6h4����G)%![�_^�.�6�l����b0FFu�y ��#$˦�"�+w:���|�|�o��KU8o��K;Xp.0�62���/��IJU�@�����30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���șs	R�KF�Ǌ�pxC?�ކ�m�$�������D�29쩑�G]��f����qm�O�2ڡ�?|�>jGG�ZB�x���;�_�K��@T�V(uz�;G�7�L.���S���,\b!��IeT�������懎'��3��~�K7$�!2"�fyŻ���r���������������C
�P߯&��"k��������;i�M�'Wl��s��(��-�XD�2�����b�3VCU%�'��f��k����D��z�0�1
b��{�Ug�tjx�Zg�<�(ݶ�I��6��$i���-z�w��'�?!~�0�"�+�/Q�Y.�*	7���g���wE"OxQc�ݦ��W~D�]e�p7��<�E���ȇ���� _DT����a��8�����+=(��?8ۦkV@����b�v��Pz3�P!����:�~p������fP*�{�J��O���8p�tI=�8>��{��5�xRd��ԇU����銓�R#+�3p�ŏ񖊋�m�X��їП?�� �R�6H�`rGd���wV]8=����]�����*����
�#;o8��,٩��+������A}��D<n�Jq�wFtUu8{K]�:��G��)�:n�ǵs�ˊD������{���%�=�`r<��Au�����9�C"G��QSF��� í�?�^1�2�pZ���zg7s�o��pf�~�Z�]��F�-�&�׹� ��G��c�
��Ǔ�����.F_�8+K+AX�,w��9��6N?^�XHTb`*1�0�����}����x�������s�B���'��
W�|�1}�ˋBĚ�O�wN#�W]����
_�FoC2�`���d)��8�Wb��\�),��w�r�1�w�S�~d�|	[���^��|�S�R˨���1J[Hv�!L^z�����P%4�Ͼ�,��9���çSev��lK�v��k]�p��d�$N&�o�=��Ϫ�	���r�hbS�ڷ�^�ު>���o�	�����@Y7tr��&��)��#y%�؏����x��Y����;HP˿��Q�Z��̂��q��^)�a=�7&^UH�^[�ϕ��Ŭ=k�k���\sI`�tZ�&�#
~|8�e�W���!��/s�<T��.���4 ���MM�J���N���>�q���me��pjM���)YY��J�'P�7�3�E7�?}��C�K�e4�d�U�`�'%�Z,�ձyε��D��=�X�4����N�ƪO��i��l���d��y�Fh���"����D.�I�#R�Ո���U&�W���td��Op�5u�|�w�ie�П����=0�UMw�q�$
��ô��l��?�x08_��id蘱�|�v�s9����y@l��;#������f���},w'e9W�3~A{��	���/�8����ƁU��b���M�� J�O�pS�B���"e6�G$iR���Ő.�۱ �E�*�SF01~zm}[��r��<ǿv�t��6�Ǉ3�HcUz� ߗ�-�+Gj�g���Dcw��B�̘�o6X7o�]'b�ԙ�y��zf"L�EդY.�ed��y��)T棧�s|���p��{��|���.�'/Ny@l�a_Z���\ )�U{��� &_�Ajf�ᆩUN����ʈ��7�{� Mj�yV� �`��_BUq�t'�J�&	{�/i�q�)����G�F��DIȓIFG<�5]�I�/��4�f���^��g�	����P�<��������@��/��dLs��5�	2h�Nv˜ۛ`�Z}H��c~��§U�86{N[�y���/���7R�鑡�4F�h�i�5�ʳ�����C������v�X2����S���=J���+0��N%Y�),v����͢���"��։J,�
�\
�u��ٛ�v7��-����_X���\���(��qH�i29ĥ�xI�n�6�f���
_b�bq�춸�fC+�����#Km�uL��6�;�3㾨����/?�rX`��Mq%K&���ٝ�X�\"B%���f���X��2}�È�^gI�ɲ�ɿ�pY�%���#/��9��N��{4ـ� �ǳ7��&�?�c����~�-J����0�̢Q�"ҐL��e���r�V�������^�}�:f�P�Z@m���@kyQ�*�F*�F���I5����f���K��x�[��٬�Gn�a"�����8���4��A�~L8�29J��ּ�`PR�:�ijt���� �ۍY1�R��D_��^�Zg��s�<*���Yd�,�p���tE�ӕ�pQg��l����@����A�>�[t@�	�[�Ǖ����Q,/�ξABĆ�C@���B#`б:�H�Β�����A����(�	2�f�{Y^��^m�|�,#���uN6%�%(�fM��G���P������cA��]��hk����iƺ��N��P�i��k��a:����3� ��T]���d��KvL�Ȝ�!?\`��.����j�Jb�ׁ�]�n�A�M�U6r-D��8ҩ'�D���{yOL�L�)���<]@6�{w�U_H2g^H��fz�@�����psfk��e||�$ZȂ����.��� YHWE��8����'z>��[�^��G���6��0Ͼ%+�	eH�z�"߈�g� �(+xb�Ըך��+�Ǎ��I�����X(��n��b%�����yHt7f�#�E�n�.�e���sߡa����s�B���p{[��|�{!.vh|?�@}�_��Ȉ2��)f�/{DeS �j���"�cn��NOm����$)v�U�<�>��Z�J±7�|��w7�E1E���#�ֺ~�zAY��.�"��R
�E�*W���i��x�[J�;-�>�:�C��DXڍ�y�t(FP�ww��U�V�ٵV_���q/�c� ��C�ɕ�a��K�5La����}��&��_��/��)X�57��K&K�9�Z�z���\�O%Hf��X>9}�Q��mHI[̲�R"��u%�B���d7��i����+�Fղ/%�)(�ħSIc��d�-�Bh��4oQ|����o��H@�k�Q�#����Q��%X}(��fs���®�4���!~���*N���N�9���f��KXtxLŗA=���)a��R��&�8�al���RGx��WWΚ�J�\���:PRA����JC�{�����$R��_�^7�g?�~[�"�rt,M���X�\t� ѕ>s�g*RSlz���#�:� �A[I���%t}q�s����V���nm/+�A�����[�����O8�$U���oݳW̃�}��K�(���T��eA��zfm7��,����+��6�sa(M\�M�B���������8fc��5�����;�C���"9϶��PsW]���3�ɸ��b��3�uܼ"�:��ϳ5��0I�!���`�Q�X#KjP��v���U��na�M��6�N���������Y{��@�vUӃ�*��١6N��Hw5	gƸ����21�N���V���rD�3�u]� �����<��>�"$7����h�9xs]��"%�/��/.���7ș�/����OB�F����M�VD<je��7�Z<W���Q���vS�j��DްK�)��B�ŵ잵hB�Kܗ�ܾV�֒�0γb�h��Z��욭Þ�d�H7���F�ϰ���N8��kJ�W�p4�&=8��K�@7'��F��������s�R��3:�ře_��uD��V���:�I!Q `�}R}
^�*�d������+w̓��a���5��$���c��Z�w\�S��m��6kQ�0��j���m��+0�a��.}�2�}�I�f�ǬB��^�=X��<�@*8"ǳx���qۻf��bK�5�xv���=Y�YWat�B�G�8S��:�<o�}G�|?��sZ�G�Rkd��;��A�r����ӽR`�p_ƠL^��Vg?s��8����.�,w*"��M�tW,]�(gT�l�w��͚����qA����t)�5[u�G9�������/�uA�a�_N|�@̒�*�b���l�Τt�Af���T���õ(�`Dɸ�����Q\�m��,u}8�UR6���(��;M���$��"G]��Q�c��n��v�:�D��9��L����P�̿�����0y��me3���f�}�$47��/IԚ�g!Q�`��l��"�j���� >q�?_�n�m�M_�f6���풔��gR��{�`U�`Fw��86��6����H�Hzg019�x}51m��,.��P��ؔG`]Q?�Y�1��1��{�u"NY�xW���lv�#bL]�"�1�/��L.�mS7�E��a����O,η��w����D�Ue�'�7א<���DG�;��v��LUD�^*铌n�lE�m�D�_۳�5�7�WV�@D�څ�b�Y��Q�=���T˃2I.�ޕ��&������b���+Cp��=Ⱦ��5l��0y,���Řc�ϊ�w�>��RW�V3$�3���Ԋ?>f��,�����s	� ʔ�R'���d�gZ�Ӭ�V�m�m�@�J�W����0�ey�Z�:_ʬ_�7QX�&>�n��D���g��Yy�e��f}�K�P��I8�S�g�Tk�������;���M7uB`W�=&��S�Z���̥�;d��2-�JZnn �`U�W��@��SQu���Z����c�-AM�iR������Z�e�y����|�m[��l�kl��5�5�M�^�DY{饘L����̢Y�l��/��1$��p�ڍ�nfo�����	S�&I���`�2fN��gA%�A��n���S�Y���ٟ?&��nBi*����[X@�*\o��̶H�˅1� �j�T�����Zj�v�%�"���u%J�.K�Z�g��Cf�f8o�d�vZ�"n Ǉ5��4B�����|��v6(oc|Zt�e���F� ���I�x(
��?|^�i!1��5��8��֑�7���I�	�����iV����#�Z$�	�֥���cC��6��zq@0��$ў�#�ͱ����uj�%4@O�@j>C�0�nPUM�V�ST�!2����?�kŒn��bl���BY��Vzח<�Xu,�92��m����;;��*�C_��I�#�ܺ�()r�h��.�r�K�6��EdZvRmUR�>-���;ű�)��]���x����
�T�>�>)v#T��P4�^o$ĭ��n<9��ҋQSxε���5��de&�����W�����}�*�F������.YӅK�eY3�*��7
�@6���?������tQW�=�4�CB?L��m?,�?F+mD�
��9/Э@��|���mBL����B(�c���E�D�8r�0�JS�^���q�j[�L�W��d�&��$������5u�>�� U���ד���{x���E��>@a��{����� ��6%V	�vZt�}uZ�Y�;��n͖]x�sm|�ABО�^N��`�(��Z ʿ.?lbK����5��K4J��4���-;�(g8�Ⱦ��nB��6�$cAY�$fF���%�����o,;�?&��2KIS��8�7��[m����ѹ@�x:�W0�*wq4X����󻛁lM,,(�&7��g�'�}h�ǖ����?���wދ��4�\�UqJ�'��,]c�y^�ݸ�uFN7��s)4h��c���:�ǥ�6=�i<��}&
UmzF�t��\:�R]Z��B��܀�U��X7sj���:�W �!_�A�ۋ�`
n�-�U��]ॵV8��B�'s�(5lz� �ٚ�NB1�#<B����z9^�ށ��я���!B�1���T�"�M�+��V���������a�0 ��i� K*������A��.,R��T�XW�h}i��U�
�;�����b6C��D�����F�۪t�b0�'	�PiX�u�eCM�I���r�m��T�V��M,^�[�PWQ�uD�W�.(Aq���v
�L�a�����*���� ��I�x��;�|j�(� �[�����%�6��7���9I��*��	�ѰlS��_�y� ���2���Ou��^�S��&�яq � ��8�"fʫe���n^�qmC[p:[�sR8� �Y:�~��0W/o��@�(��1R��D��������JHQ���N��KT��%慄V�J��W}-�V��_�	X��ax0�w}��$�RX��w�l����6�y_!H�dP�����R�4(9����p�l��:�5��^�ݤ�8�{3.'���9�q�~	��_v��-���&�z�{'��L= �M�} HK�.} �J�%Ϙe4�x$'�	�F�.&� ^E�{��)nj�zk��[��큗����t��r���ۡH���z�#��U�@�m�&+�pv�e���w�z��������X�K\���b2iBԗ�y�6f�/aE��.� r���������iHsz��.0{H\G|:B;.� �r�@��[_��L�߄�)�}�{1�4 dn��?a֌�]U�7��9�I��̦�9�x�'Vy����^΅��GU�Qr��'ܮ&�^�/�]��w���TG�����3듇��<���]?M/D�4͏O�ϯ�%~s	i����<σ��Z��Qر��b�b������	���N��ۙ�Z;ƍ��� ���6�X{�e�����R����ϑ���#h�~5�u�߽�X�"w��x?��ڂ��u���p��a�&�eYj�lr�l��'�@b���~�A�|��pt�Z�ܲ͘��ӆ�΋�d/���A
��]��ؒ�4h�D�W��¢�b���%�H U(�/���9���d�0mT,H���K�6��(���M2\����5�H�%>cf$�K(��͎������_?XϓQ6P���vP熕W��l3ٓ�Y"��wʑϐ��ԭ��!��`�h ����6$�]��TT^|�b�g������!��Afv�j�I�r�Qb�������|A� Zi�n�Z߬�(���K��?����M$9n2��К��Q��y-�y��ho�bÂC8�s�B��<�����կ��K0��b��4��t���٦��޹��4!��"@4�
@ԉ�A-J1�ݼs��a��-N_�-FG
wS�����H��[��1��r�c&��d�8l��� {�(|�Gg�p��R�F�cw���f%�����t��=�&�~p\�p�a����yQ�a�T�&����a=Q��|W�Xm�����g��ge���=/�	�܌i�{�o$��>E���B>��ig������J0��D<$M�ɂM�7$���~b�"ߔ~�I�i6�q��M�KBl�:�/�i���~�֌cq ��篑o@��$y@��h�P��^���Tkե+�X�ހ��%��B�jR�3��2�P�#�$����jvYw���v�V\�[� q0q2����D���pY��ȭ����k�g��\V�
���aYh�rV~͌2��1�#�ɺ��R����G��YO|-�=c�+M�G�X�3� 4�r�@R�Q���毬,��@�̞�ǀ3� Ÿ�a��ZDq$��Nx�@���e�E9қ&(1|΢�=��{Ө3\:����S�Ve�ޘ�����hϸG��Ij��᫬g9�K�:+�g�hIC��#�5VX�k�����chP�+߮L�����Ə`��hؗɮ���9J����GP�\���*Go��R.�\��M��I��Ӭ�(��q׸2�0��ǼI���61	�%��N
 _�)qVJ��'��Cz]Q�(��K|,%L���
�a�m���?K/�)X���|3 K5R�Ὅ�w�\у�%8$|f	X%�U}�D���I⍣�fp��a%+��꒗��K��0���z ��(���HpIX�Ν'c,��ӌ-y�/��Q�)lQw����J��ɽ�reߊ�?�Y�Pf����G8�)kՆ`:�z豬�T����8i����B$D���Y�[pF�B%����oӈ��ZqƭS�>��r��[��\��T��?� ��:?D�h1R	׮�[� ���w�W�/l�=�5\�v�h���=A��J��YM'�V��5_6A�H_`�n2��G������'r%���?s��}Q-=���	#�a�������H�ǪHw�w���]#ܮq�&�8sv�_��+��鿸�.�-w�!#:�d���"����v��0[��C��[z�>�;�N{�qBÒ��H���ۤ=��f�ާ��м���YV,b�G}���*���"���|ub��o���n��wؖ�����*"?�j`<�Mۅ�u�|�	��.Bw���|�`���n��Q6N��q��^%)2.�����I��U�=?�j�Q�@s�B��#���{��++�,s)������0
��v��~8;ٯ�'+ąR�L��}>+�<tg�7|�F�_K8\��]��5��)-��D�s�"<
���Mb�b�i�#����`�?�����������C�����x�L�k����ŭ�1ތ�p
�����z�B쵨đvR~��[]��KF!T��,5P��Q��4�ċ0W(
����l��Yf�F���+Q�XҊFw����-A�r��eB_�?�ٕ�|%�mL�F���.�kp2���x2�]Z������nے�Km@�2���?Z�P>��GKJ�Ȗ�6��z@_�(Hsd�:��T�Ԅu�'G@�LLL�ٙ1���4�!a��g��T}Y�*�q��yi���\�պ�!���f�{-���rD�{�T���2�����U��o8p���Śf�HPB�vз�Y<�M���~+�уq�Z��/!-O�?�����	!Lb�h�C��{�t"��[��ߜ�\���,^Z0���bd�����t��(=��6��TV �	�6�B���@�WY��}ZJR�����/aO#"N��,-��8~.$W�[��������dա�[VR�HsQ��٤({V8�;L	� ��}rғ��}�U��1?BEy�Sv�
g��F�j}=��B��7OT��NDL>W	�����
S�oo��e��B�d�?*�d�zW��\ܹ����h'1����VGd��]	��	�Äը�+��L��I�1��v�S�
�n����#�` G�z�R��O���p��b���q��E�uuG��.]�������W�(&7!D5��=�d����	��prV�dS��
��j,���ζ�� �J�@���rF�9��k�nڣ#���̄�
� j�7��2 ��,�P/��T�]Z�1�.�(q�=^�L�=绳&
_�1�5�{���f�k�k���Zs���t��n&n�p6)�8SvtW y�f�q!)�sVæ�'�wł/�A��M�IU�9�������h��qвD�3��7��MH�	UW<Sh�G�'�P��ć����?0l��1�w��4��U�'�>w,�uWyz[�/�b��t�46|o��_W�V�	��%������,�q&�F�Q�x��R�͜�^��|���vFs��0����2�=+J���ۧb�`��-��n�����r�h��N��C���`�z����6h�BM�a#؛����[z��Ň�A���׏����Bd���B�T)��󹙗�3�`��:�����/��}GQ ��iߥ�*��Ĝ��Adށ.Hу��s�p��Wr�Ei��#����;�NT�E�SC8�D#������F~C~my��ďi>z��x�>�=4E�K����v\�zs�[Ŝ�퉬��ʚп|��z>c�4�H��z����]��uk�+����m�J�
ѧǂi����r��X�����b:/�ԟ�]y��f���E�j.�됏�����H����s��8�6 �{PM�|BTv.�Sl&�@��_��Q��`)��k{9$ l��G<�����U��A질��ЭA���(�y��f18�%�FU��I��t'�U�&���/�戰�!���ϝG�%P�� ����<���]G�/L��4����"��-RI	!�I�$߉<�:�����Yq���p�j�����	�k�N�?*ۡ]8ZC�������o�>'�{l2��F�Z�~���%������Ghw85À�m3��Ew��[h�|O����<F{�2�YJ�Nl+����Ԛ��oRF���֎�r%�@�6��J.�^M/\����8�|�+�󸭗�N��;|��
*�(�?#q�_a2���~�wIV
p6{{7H�����
_(�lqM�7��^/C1e�¿߃K���L?��A���}�e/�X�Xf����5K�r�8%�����\�%/�f�B�X���[�I�W Q��JE���91|�{���J�e�~Ni.�uY��D�.�D�<�5��P[�H��Nu�3"[�`��z�rM����I�D�WL ����1���Պu�|�w������Ֆ:ի7����q}��s��u	-:;,�G��rF-�COڗ�y��6g����Գ��\�r�}�.0O�~aT[���!��7�)sU��`�\1�`2��͟ ��J�N�)*�Unr��Z�zr�l�b�Bƶ������ȑLX�0���?����4]�� � Um�~g��{}Xډp7<�5 M��I�9^j�K�K�ݦ�8���O��[
���˷"8\`�j��Yό��|��(8|��v);�1�����꼁�=	��Hn���W�RհĘB9i��YV�o^5�7��S��&��p"�t�hck�J�=�k5��l�%��U�d�0�&O{]x����Kk�����ý�|��UE��߆�)�xV��(��
��i���'7�y�E�
@�T�2��Z���H�
�k�w?7u���w ���,f�|M��{$c�qx�&��Oz��s��_H�,p�E�x����,�7���	�NfK�D��>��P�*�4J�@�n�'�+�-��tk�i�|�ҷuj��gߤ�F)I�/əX-L�%4����ϭ6]���`����k��r�*�5S�:+��uBk�1�rjk���~
������)��:c���R}L������ņ��Z�M�ʾ0��@�K�%-}SaI�"Z�ʔ�)O9��,&����S�M�Owapaz���S�3Z�3F;��<ZB�b��Ú� �@!&Ho��J��;�����	��L�><�V��H�:�m�����\9�$h���B�U�y������`#��T���p�RQ�� ������n�So���m�}�������5A�϶�ݕ��w���ͦ�n���Q$��8kmy)HV�~#����1>����Y�o�1��H��Vv�;D�*h'�C^�`��w�_�"�9r���Jo���
>4��:��o��F{˨+痺X(��w������AZ�s���1�&�.Ť��m�!ҮҲ�A� �xi)2���p*�f�N�(�-m]\2E�?0�>��G���Ȭ2��^�T_AH��v\�P$aT��[u���G���Lb�9�4�`�,!����}�TSw����l�;���9��2�ukF.!�"f�Dl� �r���c���Ŗ����w���,��㙖��?���G���p�oV�M�Jz�v9�'n>���-�\��=��VbZ;C�{����(�ܧ�-;����y�0�;b:U�ǉY�t��S�����r��گ_�X�X2fˣ�@���I1Jh�b��	�a�DN�-���޲�w�k݉S��y[�ga��6c�9ad�֐2��wb�(���G��p�����cN����\�6��tsO�=d�~�D�p�Pq��ÓPb�a���ʽ���Y�Z=������o�"���Ԣט9Z�ʅ�/B����t}{��$�ĴE��U�!8��4i���1�(����$2���y4���|�K �~�/f��4��6�u�dT/Bc����\����~5�c���P\��ȺC�:�y7���?�P<��"�������~�p[����>�j)&�ɼ��2��c�����j�2(w���v�Y ��� (�!2A醗jn\Db��y2���W���ZB�߄���ѡ��B�Y�p��7�I`1~4Z��f�	�愚�GH.Y��"�ts+df��O~3�4id��h������=Zcv�@i���z3���O_�}oD�3sX̯N<��@߲e�k��r�13N͚�:M{J�����$Q]����!Gϔ�n�Hz�z�#=ǌ�u+�ۋ�s|���g���m�$W!bX�yԡi�9b�B}ԥ	Qyc�jf..�Ea�.��N�M�6�18�/�6s�������{��|��x.���{-@x�_�|����)���{�o�+R!R���c�IW 2�"hz\���ȳG�#S���<3l���)�e�n�t*��6?ziۛ�n�7���0�C�JǸ��֗瘊������4@�h*?U՝��,����BI��
5�Y`�f�1���j��eKl�+�MТ�Kү���ĕ��m$8�{�jdk5��4�|���}�ޥ�噾�����郎	}'%H��?�H�R=(�� �<i��V��5#��.�������<�c���⥭uk��l-�:���{�p07MO��cx(9��kv�d�F�｀�|��]E	��Y�x��@���W
 �ig��ҏGɳl��E�x
���7��"�V�rr1��7�7ݐ�����B�,Α	Mv(DY��$�ւq�̣�T=��%Ѻ�/�,؟�����V���97�c���;���)�>O��˒l�JR����c�ԓ;�'%�k'���0���!�σ���Z�ӗ'�X�w�%����x������V ��M�P)Yr	qDѝfH:�`+�ϟ��B�r��e|s�~r�����[���:�1��5�|LE���TrД-㴵¥Y�2չ����ٳN�څasS"�
�ny9��&�W�o����Oߦ=a���1��3�N�n�;��[<j���1�+ȣ ���H�H�v�]O;)�f�SM0�' L�y�͆V	�hHM7�m�}�ڂce9D����R����#��l� �cE�F�#�^�rp�Ѣ&�4�z̴"S�����9��\�{#��)A��*�Ec��0��,���ֱY��I��I�Wm�d�VJ'�wm�ɇ��av�a���������V�[�;�4�h������t�n��Q'd��*`(��%�"9���1�}���+�X�����UFeBl7ԡZ��
�J���}��Bw7@O�LN��,W0��S�
�-o6I�`�#��6d<6i��Z�W5'�\�j������ews1^���3�d�
D	�ǽ���<կ�O���/�1���vF�$qփ��xt#��g��aC����ЌƩ�lXf$<���F� w�]����������&������=""E�Ō�	��r=\�S�@`�ѓ>F4��Ty��;Y-2��Nh�@�ɫe�W�}�2�}t����M�� �l��Q^�C��S;vL�{׽����'.ҁ�s�0:Q�ó����<v �[���'8�P�Р��q�T��d_H ��e���m�)�c�5޹�������wb�^9���*L��7q�N��b%�0o-WnAw�_��۱9*td���O <�u�ۗU�� ̥��Xw���|�5o�LLrQ�x�����x)���GW���ާLN?�> Qg�S�T��#C��ު+���,��}�C�e��O�vnC�'8Xo��A��+���^F�}�8�<�	&YFD�8�<z]x/���D�)?��_�qs4L��I�_� ״T�ֵ��߫�`
�U�o';�dr��_�lC�e�=CB��߸z��.100�p�
��e�Fz�m��8��E~v*�]�M;Fs){���蹬�*�F�{����
:
���w�k�IF���+�}X���w�W�p�AV��7�.-C�+ϵ���m�l��Q��%�t��2i�:��-
��&�$��m��52
 �?�G�>�0GkȨ+��_=p�E���L;HT�%u���GxL^׋�����\��!3��yC8T�)l���������]���g�!b*�f��9�1o:r�)��ߊ���CӮ3g�s�E�A����d�'���f!�H�y�k?�M7S����գ����=��-�͚b�5�^b���C�W��F���$���,��<����0�g�b��}ǅ�0t�@O(�lX-����ۖ$�TϯG�o@���p��Jd��$ja��NidM-��oZ�>ws��Z��{�[Q>����>cy��d������s��(O�cG��Lp3���c��V��+��dmtoϏ=��_~��dp,�&�����?a�3�9�j�U��=$��1�덌��P<�5#���/>~f�_l�{���$,��E�M�w���iz�b�-/�D貾$�$�3I�uh���.�GA�~u����<��6�������B_�˂U�̾b�~�1c���̇ޯ�U%ؕ4�y3$u˻!EP8��������(����G�؋���	��j�k�ɸ�{2r��ߥq��j�Exw2!Gv���� $��2�9��f�ED������[C��˫��P��-`�,>�"Y;�L�p����1zn�d���m� c�G  pY"���p؊+���K}�3�L�4eI�$�������)_y�@}�b���3���p݅��QD�����N8�@[�9e�Yl�1/��P7{F~�/�������)�ދ;��B�+h��������yI�:�>K�����`~<�R�������91ux��������#��Lř��_�>!e4־N��o�hp����� �OL�����%��{?�N�h3�u`m�i���ԗ�IL�%��O Ū���)��6u6�*V����J��B�:�������fw~u\�x:GH�F�FO���P���S�g!�Ph���F9\
D8}8"IOa��T�I����஬&)�h��m�'\D#O��+�)o��/ʶgP�A��)}y�n%c�.�zt�=?���	�[�q����䥬��6��9t� �0���3�U ��q���yN�&J�5���7)l�j'�\K�����â8..����$es��/�8���j�tA�ch|��:�ĉL��:ٷZ,��.�	�+Hu��3=R�@AīȔi';&VpƳ5�h�C���p�����'p�c~��ߑk��l��+���0"8�O�x�P�%Ȉk�C��n����|�ojE􆎆_�gxi������
k�Li2�WҺ7#����E�
���D���w�l�=$�
#�7h�8��4����,y�M����$K#,q�v�����+����,��l��p�����_!��s4�AB���_>��7�=��J]'c�A9��^�m�RQk��i���`�(��z}������8�X`�;%�gt�5w���3�����h3�rt�L�hZ:�2t}�8D��%�z!��C��R�$ŉ�ƗۛȜQt���$)(d��q$h2�ɡ�TsI�:�6Ѿ:^m�[?�_��|q��8�(PCQ�UF�KI7:LU}������p��R/��%X<���u�K�w�N?d��O�\~r%�ʊfx�X��} d}�k
�IO,g�s�"��ǆ%x8������Z�]�&�W�̀:䕲��}�2�>K��c�*�I(�e�:�gp�ĝ=ǂ��"���N�S2�DD��)��&���]�RV��3`Zł�ъ�$��o��⟲_ 鲠R&����+d�k��B�T l�̇���4�ve��:0�c|y��:�UȬތ�Q���>�b����
g��fy�al���K8�ʨ�S�*
T��W�O�뱪�K'�7��`֭���IS>���c��Y�d�j)-��,n��`Ԋ7�cB!�/�Q�/|�YH؛s��- 6K�S���ں�H����@,���L��+'xk���(%5��Y�Q}�|Yz�ژ+���C`��q&��볺��Wׅ�#8ne���Rt��(*&�g�H�!2ſ˻���`^n��KS�b��h�H������di�_»��9@�kn�̕�����\ֿ������O.�Z���:ȝ"��,Tԕ��Z�(�gjc�f�oo��i"m�ʇ�4*Ӎ>|�6՝�c�o�U<t�f���kr ܷ5I���
ci&|�!������WpQ֐�U7�0In���:D���!�Q�#��l$�h֤��B���ԹHj0uq�����#����Euip�4�Qm����>��0C({U���i�!Qp3���wk�t�J�!­EZ��!i�a.�� ?X��+�8"��L��F��;�S�����X�[֓���)q �h��±�h�r=ު�2��nv���U&`>,�9��	{���������ƌNz��I���]�>(#3�~P�oô��ls�9�=m�Bq@��F����־�e忭�tn�"�\�x �*�5S���/����df�e��*(J*7��96;�?ă���s��W�fP�k#��Lr�m��Y?���D0&���Ќ9�b��ڇ�L����(��ޢ�d�6�7��~�	�^/���v��j��f�B��'Φ����ψ�`�h���� �
K�6´�#�xx��E�<c�@�:�+w5� r[%�&���#k��nEZ�n�;����U�ד{��fhT�ǋR�_�U)�'m��,�y�_�K����� G�4Ҳ-�j����/��&��!#{�5���F����ZR4(����8٨�mw�s"�֠�,u�ƚ���z�����Ch�`�͌-j���������5���e��~z=���R}�B�M�#�gⵑ�Zz�쮇��R������·�B��q��j�T����8���y���E�v��K�^��� ��"i{�J*˹��Ij�A�Q.�F9�����W�vXir����
�;t�
�a��C�>�D?v	�@�c�b��-�'��kP!c��-$�C!Ȱ�w�%�1T>��D�^�'�P�4u�r����sA)�h��U\�d��[�.��'���q�JR�x��X�4������R[�2!ϩ%�@����n��d@I�)��/��hI��e��1���T���Ek�u^��^h��V���G��E�M�C[�"�j���b^�0�C�Jp׆d�+6k��!�Yҹ��6kw0/]�P7ɼ��e������^���K݈��J r��o���z	�+A�<�J���W5�-VF�b_Lb��0�4w5ڿ$@G�ê l>������_��ZdQ��p�>��z�9��L�o4�l�9��Ǧ��E�\�w�3
I'��r9���~7g���J�=���><�7��3������Q  �e��-�����Pe� $�����,.��� �@�E������&��z#]�[u^��9�)�z�V�,��*Xǽ�\HYX�z�����?�%�+=LO�������2i�̎�Ĥ�X�	��mb�|7�O�RyM�fXHE�'E.oG��7�ѡBP/晵s2���IV{ ��|�.[_Tħ�@�Ƴ_Po����)kϞ{�3� #���J�W�U�\��I�=�w��Cp��>yL͑����՜�U�����J'�m& �/�V �g�3�v��GV���z�B�?�<mZ]��/�4�׸����ݓM	�5���L�<�^z�q���	AV��6��2��O�	h�ENl]��Q1�Z�/~�T�Dm��RA{�d����
W��^`�_�t�j�1hʜh5s\B�?��y�Q��ٓ�,�:�E���%���lJz��+��������,�k���C�M��z��5�J�ig��L\@���É�,`�ţ¬�5�p��z��(~��q~��2/D�.AUI��6+kt��w�5jB_��q�?Ŷ��eC�X��oI@K��L�����4�U-��/5FKX3�����K\�"��js�^�\���%߇"f��{X�l#}[����zI�QM�M�͓滌%үO�>����w�����R����}�x7��uoVc�2�\��-�s���bN�Q^�<���IٛR[���Fٹ�
_ힼf_}��f������4���a����*\6�(����1fe�K�Hxe&���h���Za�����C�8wV�M��`�>��+��(���[[���#R�w�_;��̓�������R��_j�^N^g�7��2���.��`	,�����t��n�L�Rg�8�l�t�q|���vA)�(4)Nt��>������μB�/9��AxU���a^P�𒸖}��q��H;�eD��w�E�ٺz(U<���#���uE�m�,�?���X	6�<(��M@Y��fGF��D��c��#����^K�Ǒ���0d�τP~	�D�d�׺�0<13����
�w�H0rρ��ԾR!��[`�NQ�&UQj�V��ĩ:�c?�n/RVM�l�6(#:�冩]���'g{/0��
΃_�e�2
6��
&\HEC�gT�Ð�	1�1H���y䑭���%�AaZ]��|�}�Jɦ��Ox"�iH��|��g6�G`@]Z�w"�Hl/)��.�ݡ7����?j3�O)�ˣ�3���<��󳥎�D������m<p��=��n�扣BNZ�K
�°V�}��<��.�FK�8�"Z]pԖ�׈7)7x��W�Cs,�����Wa3׬�eܑ֭ߣ��`
�g�+�\K��W��C�\��5_֜J߰������1(B�p�[x�]�Yz�ܠ���� ��~n�z]�xKFk����}������>}�zK�
2�-�����cnqF��+�LX�	w����w��AN�K�/��%^>�#IФBOm���(ˠ��[�l,�2a�����H��7��m�K2o�?�u:>���G��Ƞ6\�ҁ_5�=f��DTq9u��oG
|�LVZ��{˲�T�!+ ��q��T�G����#�z]�����m�_c!Z��f����)r�~���~����߮�k;�9�a�ד5���3��@%��c*�M/� �՛-��=5td-�W�Zy�y!b��&C}X�>��$ҧ�ܦ�c��O0�B8b�l�}b�t��xG�	�d������j��L"
?�@���h��J\�����aٮaNa�]-�RՑww�ԉ��s�[I����scqc�d�.��u��k��(G�MG��vp(ǐ2c� �kbkӏ��"����1k����^k>C��p~A㏲E��?"�Y�̫]!�0���7)��N���H�ƃ��u��^J'_�v��M^�K[0��;gJWGW���V��b_s������a�w��)$�&,�1�&l�؍5��_ 4+d��WY��XS9m�����/l�O�0*�=s6�c�z�¦'Vb�94$�~�|�%Ê�����*�,��8^���ثޖ���� g���-*��� ��#e�Ơ$�u/�P�.F %��E�#Ӳ���-,z
��[<�����P忓vU�qz���H`�z�n��ԛ}��<�+ĪTԄ)�����Y�̕6��/�Xt��:NHbqrZԶ7�y��Sf$�E҈e.V���P����� B�s����-S{'��|�!.Bػ�=/@I�_ג���~)��H{~� #����g�8�U+b��xI��
��8�.�i�ySs����Ü�UNk�2j'��v&��/���nD�]IG�S�!<��Ɣ�<�S�]>+�/#
�4��w�nC3���	x`�[�,<����	$�0gk��!N�~��� 	u?N�s&۸�Z:������FI�Օ�{��H�V�$Ǒ+��a����㑆hѵ�5Z�
�6ӽ ��X��.������Ja+mԾ�+�Ă�[X���)���ޗ}��|�J����#�\��Q�86 ��#����\���e�4�(E��q%l�2�Mi��{�IMK�6R��G�� _��q�k`�5=fCH
�¶'�K�D&L�:���
���D�Λ/�}�X}[��
(K�������E�\_>%�!�f-��X�$}a���� I���4�M��%y ��l��'���@���2��Ԗ�d��02�w>c/��8�-������QE��U���B��������Q�$�� �}�#f�o[Ǘ��٩k5�=۫G!	*���Cݴ���fL��K�o�x��1�V���d��a��]��kD8~E����'dr�[��hլS7ۯq!��K)a���۵���y�a�>���;"�J>[ӿ'�Ԝ|ƆP��kd��M�
�f���x�Ɓw~�Ӏ�X���%���Xɭ����&��i��r��Ѧ�3:��|&�#���r[�U%��~;M�����ԫ:��Q�~�L����zw���<�������������,�e=a�G�"K�є� 19ޖM&�����Ge�O(k�aKG����&3kk��7�;iz<s$���)��t�2 k�Q1��H�h(�{�=;>$�\]��P/�L��1�EV��H��,m°��k��9M�k�/�����{���V��\�����G�p(��O<G#R���\S`�h���YH{��d[��%�A 숀�Də�z������k����2�m�XlVs�ͷ�������2��
�	į����ޤ���V�;���h��x�k �T^Q�31�)�(����K໴0��}��;��W��e��� BU��c�q
��V��}M��B s�Od�NT��Wk��&+P
�oG��]��R�Jd�{~�tUVW{L\�;ԩ��!议�1Ǫ�`d���	�{����ո��!�ɟ�1�v�m�NY������p�l��g,�嵱�������5���3��%��)3�]��		j��g�z&G[�E;�=� 4��Dz	�8rf�$S\��VZ�zv��+l��տZ�d@��rV߄�''�~2#�V ̔S��#�G���B�;�P~P?D��d�\Zڛ�>��q��^�<I����dG`��}ӹF"FQ/f��.���7�ָ\y��5O�����v��x!�D�v5e���7���<�\��8�ȼ!���ҕΌDiR锂�֍���A������������V��=㻐�b�|��6��Eh���׃�HͰ�<��	C��kz��:���p��[=)#���\�������E��WȊo��$=R�ڷ3����d�X� �l�m*Ö�L���> �R����y�d�ү������n���a^5�������0��Zyn��: ���@T�QY9�>ߊ-��Gego�yu��'V`K{A1�JE�S��T�YP:��S�e-2�76Ld`8��'}KS ���-��D��d?#�-g��n/;[`6�|��#�Q�Y�������Y-����*���Q����>j�)l��sh3�Ә�xyk-N:�5�ٍ;�t���Yܦ���V,�V���@�e}��s"��7�T�n��.ϗ��$&
���7%2gB��TX��Bkn�	�Sd�؀Jx�� V��O<yi+#�����@�R���7���lR�����5���s�Z���\��"/�t�R��(�Zş�g̾hf�l�o�*����"�����4��ӯ�X|��E�w�o��It�|��� ~*Iyx@
��W|?�!2�u���y�/��a�70�oIP��\��J���P�#��-$ɦ���(��4@���;�!0��0џ�S#����+u˴W4�"���>��0��xUNߊ�t�!s���'�kFfZ�,������#	��6׸h�X��a������ޜ(x;����$��m�=�S��D�)�
�h�9��r_e�f���F��vsa�UHd�>�1�8�[�e��
p�Yt7�ӛ�+x�ڃ>��*#�/wP�P#o�?��bA9�v�$�d�B��6�c�x�Qe�0[���ɘ��)�^`*�G2����e����1e�ܕ*J�I7�(K6�&?���D�f���H����j�:��۴�G#՚����R��ݞ��@8}�΁_�{B2��tpYdwF*%c����o�zi��N����FSV��҆�[���\
og��S�� .#s?X]Mh�.�	�^�[e���}#��EYl���5���v�1�h!�!�Q�V�ޕ�Y$&����%��5�f��\��X �sx�]���*e('�g-Ԧ~�s�'&K�=
���paNK���*���]�\b%7�q#��^�!��v�W��?�f�S�f.��;���:�8��uy(�@vBl[�C�{ܶ�l��CyOJv��},�N�'�I{�b�Ԕ���7%$�Y꫌���H���-����f��OƒI���Ǽ'c&*�.��؈��� �����*��@��Ӆ$c&�������7,ǠOy��SBP��b�Ӗ��F�V���3�AD����7c��PA�m��!���`na�u�nj�M��Y1�R�Tn�A�M2VW6�B���(��=s�DP�{>�s;�.���2�6+�(tH�a�g�h!�+�$1���������OR��pw]��;�����YV��~]"�vӁK#�����˶n�]��J"خ�/8��.��7e&*��Ow��ČO������
�D�8�e��(7J4i<���w�Q������
�'nD;�[�p��߫9�@�䞒�Z��Y�
�VG��㍶�b�\���r�ה�������@��m/��bCř�v�Pcpq�=��T���\�#�H��x�-���Z���5VR���3�[Ŷ�犒�ߗ?f������{ �U(RZ�^���&d�#��w�����̀a$��ܤ*|U��'�0���y�;:�����Qk�<>1g��!���g���y�_y����KM��\��S1#T>�"%��e&�7��`
��9��Sr�uؿd)�#dQZ-�ʷn�~�`����c�JQH��L�'�-4��s���r��*��C���ȺEi ���_�Pk�u��Sj5�-��^�1�RY�Yj��c+�n��$7Z1G���%�����f{n�b�ϩ���� &�5�|��2y9�ڎ(��Bn� �Sv�����ܟ����!l4i=Mʻl?@~I%����Ih����A�s�|��E���ZݶT��fa"kd(��!�jZW�g�R]f�z}o9��I�j"���p�45���A�
|�2���}o��^t��1���5 ��dI�S�
*%|��!Dê$R��ki���l7B�I�'���x1�&�5t#���$[����9?����)7���0�0pѱ�~#p~���Du���4����3|>�10w��U`���ƹ&!�s����kX�$�~I��a֎���/����
eLXHc�lC9� Z�z�a;4X�������׏�܍=f)��h�����Vr�V2�8���X��v��NU�Μ>`��J9�������m��+Jid�}
��T>\#�x�P'��ow4���9��2�v��K�������e�5�(���V*!�,�>* >߉��<�7έ��oeL��*ܒ�7��6ʀ�?L����&��t�W�f�0bI��|�L�51mRG`?���D�"���+�@��{��;K�L�)6������2�2�k���e`=��^㙣���jnf��vZ�7ɦOD�G+����Aב�� :������WLxY4�E����v�nw�+´ �~x%i�����\�5oZ�,;I�͉h����c��դ��h����8(��VZSSW��:lU�Ci�,��˕�^�W�RDw��+X�[�#8A����9B��t���4Y���FX�1%�4���zo���2�Fƅ�S�t��J�<[���\�d��u���� r�~?��h߾�	��[�d���Vs�/X�l�2�54�!v�M_hext����"K>Y�}�.'��i�57�� B&�����˘�㋺�n7'J���9�s�K<U�=�.!\�r�	�a_l⠱̥� �5� 
�O���5�l�Iy̍�v�v�y���门�.�	��Q�:�e�ù>���r�v�D_[X2@������&�q�6�jn5HƘ���Գ�%�i��0�Д�K�1�b����a�*ҿ��]�Tm+b�t�o�8�n�#�w�����m�*����Bb<��j�]6=�T(��Ǐw��$|�W���n.�rQ����6#�)
���@�s���-�=?���Qm@%���#�4A�S��+h,K�r��P�����|��r�8���هa�+�	+�$��}�<L|,zF�
�84��]������f)o���u�sz�3����%��:���5)߱&`����?[�����e7�C����.'$d߾_��9�k��@]rd� ��$�gu��aJ���`
���Ӕ�MF�2+>{X_�w�+���ǓA1$�r!�Ȭ��&l}�iŠm٘�����8��O�%2�����6��z��3dm�2%��?'5�>u�mGX���Ck6��J/_� |��g�\T��u��uGM�[L��˙~�ط��!�H ��1TJ�����C��L�ŵ�������Α!�f�>��=r�Ǟ��M�\��ǖ��h��/�����@������%�+�M2���̸�^�����RI-�l�����l�b�)�8���B� ��:Z3�a�5m��ꫪ5=|D\J \�CS�ڑ�J��ʶ�/���T=�{V��$am�Ehv���_�hOi/������:X�S�g$�z��J4V����\8�~*j2�\���6SNO�?�B4�\�����Ӟ~f�c9Z̐���Y�L��E�y\f�0T]PM7 SG�����B�JK���+��� �jC��z�2����m�f$Oj>,wg�sv�]i�;k 9	�2r�g���TD�p��8V]��Cޭ��3ڼ��}P��X&�GgY0`&�����~1O�J�*h�Q�浚#GUN�Y����>+� λ3q�4z#���	��t����U&@�:����3� ��ۏ����D� �^N͔�@��`e��m�cn�1D��F{�;$&�ҨG"�c1�`���-h�A˚��^�S�4�/m�K��U�/��B�L�d����9�%[x�5���X#����C̆��eI	�N�Xd�������(i�����}l�ZoŜ��{N� 3j��`i��^֨	exI!c��c>e �g�y�x���uWǶ������8�ǻI:[G�*�����R�uQ!�:���GFߪFu�|OYQ��eٸ9}�g\��Eӝ�M�\?@f}�6Oֽ6T���i����)��[�m�\y�|�p��y�� %�D��$)r.�n�Y:�c�KzIx8���ڶ�e�*�����xO��d_��[T�Mr�	�E�m����U����lf����q�p�#�㻁KaM�2��t]T�g�X'�gE�-�����|?zn�dËA��4�j3UW�'[?�,Ç�y��ϸyK:��Y�N[�4@<��I!5��p��_a���E�c��E�F^b�ӂԳRC9������:�ە�sP������tJ3�G�r�'��1!_`p�;-�Xv�CH���vv�u�M�M�/ z+HE� "dBW��#"�k�zy8�n�������n|�GB�r�A�T����R��=�x��M��d������ �iiW�T���6�0��Ȃ�@E�*����  ���|�fI�KyY�x��ڗ3c����Ha�Ho��߃8�0��r��Ěȍ��Ό���?R��:��R����w�u�!���\�sx R��'_N��^�E�g������e3j,���J�t�����Hg���ll9_�U��rA�k�?�t����<�����H��Π��/�H�A\�ۆ�N4?��e�c�>p�,w��ɹ
�[(�=�(9g��@��s���5mi',����Q6W}(�SMg�ú�~�(m�(d�cF����Ѻ����uP�Ɣ3>�h��Pe�<�(���;�֔Jp3a����#��e��"z�!���`cT!�
"jBEkܨd���V�nV5M��U6��u(�ATU�y9�{����E�C)l����6��Z�e�H)=�g��� �1����&HZ�դ�z���I]�MZ��\��.pc���"�Yʁ i��K��˫��]>"w"�S/ϒ.�b7zN���z��3FVO�i���ʛ?n�Dn\�eGQ7_��<I*R�̙]�ç�x�1�\�rD�������]ȵ��I��5^��O-��V|�R�b�vb%E����nҞC�K�����f��Ϣ�m�7v�����eT�p&>�=P)f��'�ŸE��Y-�MN}�o6����	R�3�p��K���x��>�ڈ��Az R��R�R��r�d��"�R��]Ֆ���y�������/L?0���yU�I:�慬�:nQ��->F��tt3)Dgv��y\�2��Z�K"�r�їDSF��T�mwS<�Z�1i7�'`�M��f�S��
�t�Y�k�OdFx�-N��n��b`�#셌�h�x�NQ����=ԛWd-ɱ��Gi��lX�q���F,�p����&��V���[Gk������5B�3���X�Y�������1آ���/���5���b�n�)�Ϟ�����&�f�Q�2��i���{��\�nm�Skm�1A��;+���hi�����J@3ğ�p^�>d��S�֨�o��e��x~�Z�s���Ʊ"V���Hᕶ�5Z�3�gs��fFFoN�����"�������4ʴ��v"|��M���o�Qt\m�F)� �&I`
L&�|�f�!���9�G��y��ؾ���b ��{c�8ш�x�� 9b����(�l$�"�2q���]�xz����'�Fu9)�I~SUt&Ŋf��s���<l��J�Oؠr��!�K �%��6Btm���x:e��O$�c��	@.ۙI ZL�E�4��%�B�
z��5[�����E�����ȥ`�F3��Y�'Huj(z70a�)���?8+Y�Թ�M����΃�̪Z\`֭X�vޡ/v�b����0yyi��f�>SE��0.U%�SSء�4�-�s�
9�9�{��|�e.�HK�Ĭ@>�_lC�3�)�4{��� 8�7͓��sD]U �ۖzc��2���s yh���>��q UC'Z�l�'0)K&�#&/;�������i$Gr����[��<	Fo]d`/�]�4�m��#H��� o	mf)��^<#&\�G�Υ_ȭ�(J��ge�k�	��N��I���OZG��5O��Ԓ���d�{�RԨK�$�&S5�:޵�{z���h�F�5JF�[`�����1���s�肈ذ���AJ�O+L� s�;4�⻎_����	C��J^k�*X�\܃6���|��s�ſI����X�pp�V�D(�VMqP�2K����0�I"� 6Ǳ�����ǵ_�wq�t���dMC}$��:K?�aL%���=�PLR��a/QjX����ߍ>K��;�=����\�W�%{t�f�`�X(��}6R��a��I�Բ�:��%nx��5��NpI��N��MGm�����S����c�j����-�"��z���Q�c1�����7� ��C���&j�X��}�T�f]=���ٞR}��|� *x����r���&
ftzK1Q�x�����([��l�a�\l�Yj#8��V�q�|��P@�D���Y��BrR�ǀ�{�-����)ݍ+׭R�a_tJ^8�g��NC�E$��	z,�m���$t�?��h��g��gl$�^�N��*�Aŏ�P�ti��0+ZjW� ���X��/UX(A�^��y2��G��%����7��䧮��|�X���.�(�3����+e���g m!��,�X�����67�(7��M���d�=b�e���c����X/ºzw �-���L�� tPX������Ȕ�0�3�ܦv�d/B�����S!���`|��%Ij�:v�`i���n��M���6��J�-n����+�1g�{�s��������N�j68y�B��H��gpҐ���1�Dn�lQb ܤ�\��]�L]K������������"����"	���c�]� �"Ŝ/�[�.Ѩb72鍸[lS��n�Ol�r�Q����{�D&!	eѢ57t<T�����{"05<�8�Dȱ]��G֬h[��R>�����u��OeV4l���b����R6�D	���U�r������Z�J���r�ѝ����p��=2��uGM�p\�lG`���ȉ"�'�9�~��R�X_3d�R�L׊)������M���,� 
 Rg�G�T3dGsY�����ͭ�ϟ�6줗ck����0Ln�y^:�|����Q��o>�1,&���g.�Ny�O��(=K�c�ʉ�*S�JWT�I/t��W<�_�7�-�`�
kf��S?~��,��#/:d���-�n�+�`�D�D���0�vQ�qú�����	-�Pu��C���)������(��R���6�̬2�k�\mu�5���ZzV�"Y�����2�Z@I���y�2ڹ�������n�b��V�I&�<�	�,2�IA���@���]n��;S#����t���Ȯ�ij:���B@�5�����#A��;�`G�Ȕ���0Z�Z��p�[p�"���@@�n�sZD��g+Hkf�!Jo�d���"��u�4�ۃ�. u|DL1�o��2t1���y3 =�I| 
\|�SO!q$2��<�x�M��`�7�בI�L���G��i	�2s�#��$�T9��d���^t�vY��\06��޽�#��h�u��A�ɘ����d1�0�D/�#E���@���l�J�eH�5��a�V�NX[�-Ț�	Gw�2��0��ʬS[�l�����ch#dW�]�}�
&(�p�G�\�pM �ކ?c��[��mϵaQ�t�Qc=��~�#p[K�������a��������/�=����r'�����?/Řtsʰk/�>���>�{�~$[�2E������f�i)^������t�$�$�Ʉ�y��P~$y�ߖ�����6���;Bnqt�q��̍��~`Y_cs�B�;We���ěyBq�˪tP��M
��V(��mY����غ�r���j��bɇ�32��%lQ��g�j���wa�v��� �O �M2l*��HfD����"���������$_�`<��)��7�Y�W}ة0��[q1�7�O������G���Y�a`���d+/ɪZ�d3��44���ӎ��S���(�	�p�@��Z���3����w��Dz�C�N��V@�q[e����� �1�B��VZ{Փ�����b����Mޚ�t�1��hQ]:��~����٬���KEP �)�K����a<���9��xMC��7�|���{�=��\�#FeY�N��a�������u�~����Λԉ~�J!XN���3�Ux`�0I���]I[�$��2� ���s��W�u��A�yf��ɬ���:�)ʙ�0��s��F8u˜l:=��G@!�F�kO�����L3,
g�H�(��\9��}G�GOP@kT]�ˡc��=�S)5(�꼋�\sz��%3�}^͡씶���%)�7nt���]Fz��|.��� p�
���d0�Sc��2�T���E�^���U��� ��=6��Zey-<5�9�����;�/j�K�%L�hM���W~��n�3s��
�8^�Vj>�Z��|D��:�ĸ^�峒̷I`�����	W�mH�<�����R�' �ڙ0i62<V_��5�_�{4W̑A���v6�c�+��u�k�S�l�/�Ο"��n0��f"?�4��g�	)..MPX�N�(:�^��NVP�	}cv[��[͝Ɉ�}ç���{̠qظ���JEH���-��(�ɝ~%��42����u�&J,ba�{��5h*�Eo��i�5b�[�o��n|�nwE!�֦�*��b��o�<�����j���Bwj+�|���ɧ�sdQ#�pł���)���@�5���g�71?At`Q�s���@�#�ϢHy5+�Ⱥ,�8ޞ���}��FG6�83�9�|]y+1�аYg�}�x�<�j�$��F�jz8�2�]��Q�zT):�M����s�"������S�׏����{*�F P`�\�ʽ��(�z~	C5"���iϣ�S)I�Ұf1��pW�ֹ��zzu���Cu�~D]���F�8�y,C��2����R�]'v
u簓Q���f�+FR��+�EX��w�àZ�A��8���|(&�>��vm9�   G  I  ~"  �,  �6  B  �M  �X  Ec  9n  �x  �  R�  r�  h�  ��  ��  İ  �  O�  ��  �  ��  ��  6�  y�  ��  ��  A�  ��  � 	 Q � � " �( '0 k6 �< �B XI �O �V B^ �d �j Uq /x r~ �� ��  `� u�	����Zv)A�'ld\�0�Dz+4�D�/g�2T����OĴ�wFZ��?Yv�N��?�@`�X+��HH>S,a1���&���ghC� �=��2 ����2o˗~��.��t6��X&l0��I��@f������ھ}1�@�]CeFԝh�^�Y�fI�{b����m�5$�M��8�$c��=��ŕL^�9���pH�q3��6�����EIE�p�p��N���䧇00�j!lğ\�	��������I�T֒�a�
q��H�+�S�d��П��0��,l�_yr�'I�qj�'�>Q�� ����E�
� V���FS�kr~�����?)A�i�2�'��|f�'�RXZw�Vy��ˏ�@`r�p`�5h�	W��A��¤E���U���$�TF�<1e%jW��ڦo�W0�H	a��+[X�J�O�I\�v?�#EDFƾ� g�q>�R��B> �����)�B�n�O����O@���OL�n��0�	O�47��K�GKqx���	�*>�(ed�'��6֦�ߴt��I��M�eAI�ܛ6 P�E&�4�2��2��	hS<g�Lh�炆�!B듉?�,O"�R�B�l$d��L҉�^���C�O״.t����|����O�#$�|M��׫O�-�g)���KڴM\���O;�)��dם�:�[�O
3#l1�2�Շ{mmZr��c� �~�����-5��#'��fo��hش��gk�r�ID*�T���&Y;^���j���E��|1q�{o°o�>�M�a�iI��8P�Ϲ79ڵb%��]D�hQ�y�̰�t�֢i�V]:�׈K^��w�L)K�n	��Gu�,�n���M{q��w�0US��Q#��QR�� �#�=�tEy��J͠r�*�A��Mp�@.���9S.�G�5HD��?a��W�P���xG�.A�H�hf�)H(b���O�D�OʙnZ`��̄Q�qj0*`��h#�B#���D�<9��?��P@T�3��cc2\���H�%����BW�$�ӫ�s�X p�̛[|���C�i�'h�8��I��c���8��̓rq�(1� Ϻm��� D:� �V�M�Ą�cJV]�'�`�+OZ�'z�9񦂃RL�@� DP��Z|;���?����䓄?Q�����O �$�ʖ^Ycgg
�'��0��O��dL�	���E�>����4����	`�x�K�<p�1�#�6HR
�d�<��iٛ��'���]#)jy���6+��	q�@�>*���O:)�Ѯ��0m�K�$M8	���I]/�L�S�?U�r �  �0�A���.�Z��{~R�͈QFb��'��D{�\�N�	k� U����RM��i�'Gv���J�
K��L������MS���|"�#�����NU�T���
vGq�������(��_�O_�1�����a��`�L�B\ڈ���O�m���M�'�v1�>Qr2��:R#*���R�P�DL���s���D�<���B&�����?I����Dκ'�|V��<a�8s�`����FŜaU>��@a@�2�ܤ �h�|j��:\�� �Ux?y#AK���Ι4yt��a c�����0����l���k&G0F��|ա�_��I�/�Y��o�30l����@=d]`�l���䜼
��O��3���z��a��Λl�.=�ׇ@^�b��9�S�OӚ����s�<h `��Mt��V�'�b!a��n�Q�i>���vybΑ8b�0�[���5C���䃜"Dy8�/�>��?y(O�˧��4n��J��J�̀>v�pa�+1���?�O�5j�$Sl!v����v\@T�<
��'eCW����$LT�I"�>�xx������'1�T(�+R+M
��ю�џ�0۴cz��t�?��gR�(�C� �!a�"$��c���D �S�O��wԾ/rX{�!M�xT矀(ڴ�?q��i��6M�|:fK<(���'�$T>`t\����N�O�:�CI�xbRV���	̟�'q�����ߴ^"�mZ4(�&��
�3R<4H��K������q̜��V�O�'(<a�e�t�@���8xT*�1R!�=b!�A�t�:�K@Q7B�����dP�%���jΡsf�'�����a��gi�����lAi�	0d��m*c\��˓�M��'�ɧ����A�.����� k��г�]���'|�'��]>E�4Y�d��w��Q>l�u�х+�F�`ָie2c��hd��y5d�i҈�<��'=���O�fX#�MT7�,H#hT$2������'��JH/
�ź�Ѧ?�f�"�����}�U��73r`D���+�����=���� ?��z�ڟO� ��e���8�$��b�,D��m�Dm�(���73er�EU�!�ԉ����2��O�)lZ��ħ��O�����F��AK��h�b��z2t�L>������?����C� ���uf�TI�#,��t�FF~�`�Of7��O�5l��#�3e�����Z'C�H�b!M�M3��?	�.78X�/�&�?����?a���ygN
����E�˸E� ��`KR�'�~ X�m�YZ\Z���:��s)�f�I�m�E{�ةW�� @6)!�	�bCC�9&�K	0�����c�3p1�H�M�H�oɃ.���b'���p�s�%�⦕r�U�����Ob>���O��$B *(6�{qG1kYX���E�L_@�OR��$�IX�-RĀF���9A���剂�M�U�i��'V���O�剄��(�-�	�Х*&��'E���٢�W
�M+��?������͌���o@*m7`��T%Eۄ��
�k��<��4z!@���֡6����剅m�@�E,&	�n�D����� �[��V���ҦQ�Q�?o�,��Qld�ɾn�.a�uʒ�*-J$-��W��Xۄm�O����O���G�d@Q�ew��@�C�&}��q%
	��=�y����s�����@9�jY���|Y��'��	�j	Z��ڴ���H<j�T��5��9b�"5q�	�5R�b[�l�I柀�'|�����{m�k����A� f���䟇�6DJ����-�cd�Z�,;,ř��$���vFE�;(I���ަ��ł�v]V��E_�6�6L�d̻X1�"�cH�m],�'��:���O��oھ��]�Ĉ��RE�4S�\v. 1R�'��	S����"��LS�pR�Ź?�P�6V���'�ў�S�������t�8(�@��U��\���K��MS+O�Q��BŦ����$�O���Ò�'��Z��$� �Y�� �;+0�y��'�jZ�&��R��]�,�[��8?���'��iG�XIڶ�72���
V�l0�ɏ_������l��0yb �0p�� ��!	�]���F)`P��2�o~�A���?A��h�V��T�y%>�6cG=�bdƹx5bC�I&3y�����'N���j�8�8#<��Oh�Dz�Ĝ1a?h�+���8~f�9��ˢ8��7M�O@˓ �B�����?	��?�*O|�q�Dٛs�Fs��˅4+� ��<��/E �	ӓ"�vՒ`)] 6R� ���}�cQ�[�>��!p��V���tfņ17Nx�'�Z�[���4'�&�Kq 
>�ͻ��i���S����?�����lujR���5:lx��J��<����?+O
��.��M~r+�4U���"L-�h�9������d�̦���4�?iP�ig���?��O�2UM��5g����%����`��6��O����O�ʓ��a>	{�
Ԅ]�(L��`āk�z<���D$
c�B�Ii��l
�k)w��T��`�b��� p�.�f��D+o:��*�0�">�ՠ�/�J����ݠA�HbEΒ�yU�`�	4�M���v�'A�E�iU*���k�(���>�#���x��\2��G�jv�E�$����c�"u�t��4X�/O2��M*H��5��h�M ���"@"<s����O������O�d�O�9���Գ;���&O9
S�0ӧ
�%tIY�&/^?x\��^:G��!Q�2Q��) �L6g�ܙ��&u?F! `�.:ݳf�Y�G!�]YTj m~50���$�HO&�2��'�6�����I�vd ��Ĉ? �5$��(�z�'�L  �'~��~������&�A���$��≺qel�ىy��|��i&�`[���/R7|��1��o����D#k�h��NȦm@s��0�M�����D៸�	�O�����7F<���#��I�\P��f�OR�D�P�OP�d(��T�^dp���K,��2lYW[��'PD�k��U��f� ����5��>�b6ǒ�z���Ш\��1-?��Q����4ˑ>��'HZF`KA��p��Q���L{ґ%���Iҟ���t�O�&8�W�©ZR������ �i����ۦ���4��O�V�B�>J��9;׏�."��d�iZ"�'�r�Y������'r�'�9�Hԡ�S Ł�l}~à'�1�����\� ��ճ+{�b>�q�'�)�D�8 �}B��	3��D[B`�"\�T��ĕ=c��8Q0�
3"Z	����;NJ�'�T�i��Z��c���03�v��T��	2Q�$e��M��?��A��?A�'��$�OD�$�O��+��YN�����NF_@��o-D��Qb_�MdR��T�X�e�O���O�'2�7��O2� �r`ˀȘ0 ��U)t ��+:$-ae�
���	���Ioy�T>Yͧ+;z��D��y�T�I �^|��8uBR>P��E�ن2<��f�RaI�5:�C7�R�9*�瘚����	�P�N bh��^�FgRqS�X!�>���<�#Ρ��dG5pp����G(.� B�ӟ���4E���@Fxbc�	v��ApE&ɥLk8�+�l���6��Ϙ'��Q��&�"}�TSF�U�{�P�I>�1�i&�6��<�Q���7��F�'���S%N)ʲ엀%qbY!�W�]gR�'o�ay��'wb�'$ȕ���
��1��y��ݠ;j�]���r��D��kPN>���s��R&���l�&P;�ݝ�|c�Ȓ>]@@��`�$C���Pဍ�'��U���%j�2%aӦmZß�+���*n��R�k�;�"�����uy2�'��O��]~�e[)�H��u�Aj^$A�a��%ޘ'_ўʧ!O��a�vC }����%Q���0�/�86��<٦��9�}9����D�t��'H��xUb�*d��:à��u�fx�'D�l3	`�٦O��$9�SlvD�%NU�81�v��}Y�	5��k ������ˊ2�(=;'��8q��O�̔���G"m[��Zc�ո)3p4�O�[e�'�n6�S�OZ��	> �C
R`(�#�Ί �'n�'�s��D įϠt��J%�V0���?a��i�7*�S%�Hd���G�#�Deq�G��926PnZʟ��'�IbP�O(B�'��[�� ��Ւ1�z�1�ϥP����_ey2�'���z��'�� �B`��E��`H�&�/)�v�o�+�l+'lm^�b��Z���O*0}��OT%w���3��a��C�7-�ٚ�(u�Lٖ'��q��r͟�'��Mg��j�%�^b6ų�gZ��hO���íʞщ'�Д-���Ј��	
�M�2�iɧ���O��I�S��ԛc���KRF;>R�}���B�RmN|�I����ß�ZwSR�'���T1�5@A�q�ʝ�v��S�(=�T3��  �(�xU� ��,^8|ҍA��$>�� $�����H��D��Y&�U҅��?/CbС���YX3�׾m��@�1$ =��L&��CL$$)5 읹4�^�G%2{��$�æ�"���6z�2�խX�G6r���/7f2d�ȓfx�J>.���Ŝ|�dE%�<qٴ�?(O�x�bi�[���'N*5Y��k�pD#�s¡Hs'�ɟ��	0;h��	ɟ�'�r��`���1SNA)�!x'|4r)��'���KQN37�
uh�J�)��x0�l5�;��)2�H�(���	AL� �*�yǅ��L2jM�$ˀ�����M�:E2jx��e۔|�Ќ���xr��6�?�S�i���l`��)��)���	�c:n��M'����I'+��S��W t�t�������r��Ĉ؟���/�8S���F�]yN�Aѩ�O&�lVhX���?����i� 9�L�d651�!T��>�\t��,�>��Oz�N�!w�0��#M_.X�� a�'1�k��.`@>"��dhuM2�ta$�l~��!6d�đ�N֯kb�l�4�߁7�r-�ӠΏ.���'pgDab�r�m1O���B�R ��$�2��O��&�"|Rq�[�ת�ۦe�,R�N-,SO�<!Gc߆%%�P�ɪN]�'�_�'��	9�HO6�r�iD�]T�	����*�$�0�������	�����'
"<ĸ')�̟H�I՟<�I����.
��u�0C_����cqcD�c� 9�S��=Y�p	Z:6�h�|Z�/V�!Y��9	��qA��/8��q���B�,0� ��-i�e�P/Wz���'!�My�X��Oh�B!a�.h`�"�@�e8��!�fӔd�'Դ ��
ȟ�'ȁ���D�0���#+_�&
�P�"O��q��""⒁�R��4x8ԩ�>�`�i>Q�IPy���<O%�t�/ՕA@��*����o�����M�I���'h��'5Z�����	�|r�$0�������Rv|5����.�RY2�	��.��\J��ӗj� 4�������<��IŚ7�B�xe	pP�R3�RQ,"pJ��]�dVE����	�=9&: ��<9 .a�X���dY;[ ��J~0�q�	*�M3E�Im�'�F�1̅��۴P�d����'����_&4�@Ѧ���Rw'p�ɥ�M����4�2���O����H���+sϬH�:�W�\����O���D�Od��t>�R��Oc��X�FU� ���jO�+�\�C1O��y�	k~����[�gb���T%��� -,�B:��W9Zc�q�Qː9>����<{�!��Q�y���4
J�S8PH��@h�$5�S��&�Ot�j��9��-
W�ח*���1�|��_2)�7=�l�Ŀ|Zrk	�?Y ���;���.<�F������?��8��p������>qӀÜjgZ]��FI��Μ�ሜv~�#���O>��6����$/��,�2Bh�����^=8��2���7IM,�*�$OD�*u�N��G5�C�	�q��P���mY
�#ʊ
Y�#<Y�O�Dzr�͏!y��@��x�F�3 aI�#A�6/�D	�p^����O*���O��Ӻ��(�A�6�2!�9hL��4���<�`oY0
d�e��'�{@c>�&�p*�僿��*<D�D 㙾"�$Jr/��y��=[�JL6@c>�&��x��� h�z�@�j�$�R�0A�O:�CJd���ȟ ��N��*��X[dMN-Y����l�U�T��'Š�Q��3ٲ����{�(O�Dz�O��R��!3��
����C��� �D)Q�~�� �������I��4�	 �u��'x�8�t��@.  f�L���#�1��	�~��t�z����M�	�Tx�/��(O� 4j�!gв����#~0Q!lԔN�4��G0
Y$(;�D��/����l:�(O�s���p�%*��YI�n�Z�ϑV�2�2�O��U��$
���"��'-�(05�'��O�y��׆K���cj`�F��ב|��r���O�����H���Iɟ�"��18���#�!?��6���\�	'B���㟌Χ�����Y̓k�l��Qk��!}*���*޸X��|���m�#<����=�L���S�C�tu��e��\p��e��C����2�C�4��(Z"��!HfB�I#d�Ur��J� \T��'*�#"c��G{*����ɯ"������3/<1�G�K�O����Ӧ��ߟ��O�ty�'Lj��Wn�<��3B�/���6�'���G��T>�'���Ek�*H��� �gv���O�Mb��)§t����0��*X�t�BO.M���'�2�(���ɧ�l�X�e��>͈�/E�V��M� "O���G͖�C����2L��@���5�s}�")�jj�Dc�E҇v��8��`D=�ը��i���'��H�	U<@�v�'���'��>�J	)Q��1��)�M��aj��pa�Y�Waz��۰<��l� N?k�$l�$A���'���8�S�? R�ժ%=,�-���.���!�L7���.����ͪL���&�^+ }*��N��0#!��̱4H��3 i	���Ʈ�W!�I�HO�)8�����p���Y��JF�R�(̇ZM����Ox�$�O��;�?����4G+s�psSI̲{7dPr���g�&	�`,� �|��-O5Qru�I �����&��+��"lL	�4d�dd�/ML�[�0E�f�nO}�'�<1A�Ö�B˪L��+��dQ#�gO��?i��'����LS�3)�0\�%���c	�'d�=S��b��Y�v��� n���I>Q��i@�'��a�"qӔ�D�OJ�٤�A1>�~����9f3 KsG�O>�d@E\�D�O�瓠	��d!�� vuީ*pR�x��8��	��_<J�A�Ɗ�2�3�׺=��-�&�	�_>��B$K���yR�D����p+9>�~@뇪�� BRQ���`�:5�`剢�r��WZ�IK����k�)E4bD�1��q<\C�	)�H$*�Vh8D�H�,5�������q�
'n<"�Q怟�6l���dF,��I7m��oڟ���T�4��11i�E �3�<�%R��Ѓ�|}"�'A��!3�'<1O�3}�Ơp�Đ*4��!pbi�K�����"u��"|�AG��"�y�#킋}l��f@�n~R���?IU�|�𩋇7���Ş�*�T W@H�JT!�F&0�"����G)�4H�T��7;џ�q����y���0OU;Y��$��~�l6m�O���O��p��'��$�O4���O�݂q��9!��CվɐB�l/�`�$̈́S0��j*�)�ȅ�v/�S�� !���O(1���C	9�^�	�	W1h5� �[�┐�M�Ĕ�[P1�,V���~���~Qviq.�
r�ŀIS�)��'�Ű���Ϙ'��kC��5a��(�vmL�n�]��'���s��	@���l�IR!:��?a��i>a%�x+Ƥ7nQ��gܭh���f��_$�ڴ�?����?Q)O1�t�C�nd_8�r���c׾]b�/�Y�
	��gN3}� �%��?|���Dr䚅�D��(ԔV�+G�  ���W	ʄx�]@���K-���Q���)�5)�̏4o/��Ҥ'
^*-�q�O�oZ��HO�#<�W�Mk|V�s��Y�TiF�y��O�<��!�#a`3vjwJ�5)��GR�ɧ����<����HQ�OW�HA%�?���磎.sS�y�������O��d�ORQ�eɏ6C�2a��OЊG����"Ui]��!�JÅt�$ٛ�L���E�Q11~6)�i£C�Pˇ��>���t���5��,�����J��	�W��$����*,O�P-��;p�U�� N�N)���Ԗ|�'� ��
V&8l�ǎ�--:K
�[R�DB����+E�
_����IŃ�?�.O�4��k�w}ʟ(�'�?)d,�*��D(���0�6!�gƁ�?1��*u�\�`.�N \h�竗3
�l����ILwO����I��$t;�o�+���=I
�yu�R�ih���Dm4y��@�,x��J��&g�)���J~�@ 3�?�i�"}:�O`��u��
P��%0��,G�P	�'�b�@���]]�Y�U�� ;��)�����O�OGUXWD½X�p���46Ȁ�zwP���'�:�Z�O�R�'��]�����X����K�buP��6���Kzx9R�:^H$b�!H�XqH �|L>i�[�gxZ;�힞�,��%���"�C��1��q�쏂j��|K>1���>w�,�P���J� �DI��M��V�H��F�Oh��:&�xc��H<�ꬣ�!H0k�2q�e�f�<��D��`,9��&��d-�"s	�gy�,�S�T^���u.>'̨�1RQ$R���`��(t��sش�?����?�-O1�D����Ѭ�RS�ϥ %
�*˯8�
ik�.�8%A4�k�F�
ղLG�)D��$x	��W!ㄸ�"�0%���K?0~�-�l�&�d��KIw�'���Q�-�Z<�d:0��z� �(�lC��?��i��#=y���K�}�t�U�B�t�X��I����ۆO�����G������8���ly����Q^��� 1�\+,.���O&ث��'+�	��|����(,�?Y$���F��5���R���~<0q�� RV�å�DY���dQ^���YP��t�,8F.�0EʍE�1�D�U�^�y7.�H(1��s����I��M�EP�H�f��a��Hh�+r\ �%-��+�ON����7B��+�e
�ڽ[�'����ܱ��[�n��m���!$�ƀBrZ�ģ��[����?��OO2�_3N��;SLʦRΈ����_���'�.�cf�U3�B��׮P�0\,<�P�'���5��j�sZ�u`F��>&���f����<Nl��3�f�-r/��[�����1j��jD��9\�2� ����d��s�i�4uG��1�� օ�d Ōq�����,Ն:H��P"Oh�3�Ǚ|���kr
M7@XH����h�F��`�8�\!���Q�n��Y��o�>�.O�8�wo��6�d�O����<��b��8`�޷=���@��FHf�YS��� �ړL�7.���T�|��� 3���'"K�����^&,��p��EKZP{0�1'X
庉���|rhSL8H��D�x^�� ����<�r�Dן �e�L>�t��#�j��b`��_#�b�&�y�ֆ,H=P���(�r�����W�����<�"C;e�,�K���93����Â5j
+��i$r�'W�W�b>�y��U/Q�
���Qh��Q��2Һ�[��@��ƁM�*a�@���Q?fl���e��x���2��5 ����Fϑ�Mi��5�Աa.<��SI0��DE65ɠ�"@�$"�(F�nc�$J��C័�ڴ���Dx蒾)L�h�nG� �l�֠^��y��?Q��L��h��m����pe�	��:�ILy" ��+p6�"څ� ?gN����N:���I�T�'R�$Q�	�>Y�wFkɌ4� ��6N�� �2K)O��*%�	$E<��*��߲��9��I+�n��dT��,�$M(z�&��S��#wz-�B��4/!�D��0�<E����b���y��	Jv����O^�[b�H�7�z��V�%Y~��%�|2/Y�e�b��>%#V��?�I�G��������*?���]�{U�=(����X���0� ,ʧP�:*�	�;
xu��/�s.��'Q(�+��Q���L3���z��EG��`:_��ܰԈ�J���a!K���D�'��`ӮeD�45�~���M6Q�Zr�)�~�"O��#sl�*�`���Y�1�r�	�h��<�4�Q-R6^�j�Å�*�ʤ*S`n�0�d�<�F�����剏g����oP�D�B�J+ئo�c��3ƭ4LO&�m(l2=��A5�������azd߾.�V�ɝ :���"�>S�'=������Ϙ'q�,� ��
�\�{#Z<~�ڽx�'�H�� G�pT��y�&B05�	;.O<�Fz���O�l 6pJPEAS��%�#e����&`�z�$$9�ċ;,�i1��g85���OAPU0U���*�n�(R�B �
=��؊�I�8��R N���$�Ot��üe������$�xh��M�0M�S�/ܿBT� lZ8�j�q� D1h� XR'剱B�����!o��d�b(]���#4�ˣ��ăůKi�<+�? }��#��I�3�����٦	N~�XEA�lܞc*,1tnl��,O���dR��5�f랊XJ<��df0�}b��<9A��@�+S
)h�Ц�Qybj� M.N6mZ�b\��|�t��*�.M�-i%mA�aL�z +]���:��^���P�٣0� �{V
Ѥ*(�Xv��[}�s��4��[���H�+��S�2*e�\��yr�A@Ԯ�B�.�0hUhdDӊ`�P�$�
z�'W�z�9�C@8T|bz��T�B�0p�P9 ����M�wX���|�'BJ�mk��cB81�I�)@�VĆ�>��B�<M�]��ݤ;��1F{2g0�'U�ţu��+k��{A"�2���ϓ�?Q��ƈlJM9�?a��?���:��n�O��b��>sI I1"� U��\Z�"�4@Yhub��ܙ#�ZeLG�em8�')�DhG5}R��W��""!�>��DAS�7*����H�6'@��·�^`
ɟ�8�@aڇ��a�J�C�y>"����L���'f�����w�v�?�O�,���@�V�b�NTj #��@�C�	�u����-	l�2<���1����Vq�����'K�E�
i�1,�>^I���p(-g^�
��Z�j��	͟ �	��[w�B�'(�)θP�,��D��}����A�45�E@�L�b��A	� �oO�4�0$ӟT�v�Z��d�o��s&�"w{����c�
m��\��Â=c1��B��#9h< ye,A>yL�dB���&Tb�9oHk H� X�)��)�2L.7m�c�'�@�����K��99��/+���@�.D�@Ҳ��I.ҭ&�E'�Ф�Q�<�@�i-�S�8�j���)�O��S.�H	r��G�
�T����mdT��=*?n��O��DG���d��!˚�� ۶GA�X�����Ui�iV��MF>`q�}�Y)v�Us(�zUL] ��xrI�Hip�Xe&Q
@���Q�;j�(�3.ȴ
h� y���v�J���1)N~�u ��u�D�3��*:��m�b�Ey"�'��� ��I>8 � �	�?F$ �}��ɐ!��,����<LԄ0FEڑ�h�ߞ1 �i���'�70��������G�J��L�u+Qvz�kwR�������m�R-P���@�`���
�"1�Ҝ��Y�'o4�s7��
�����(34"��_�"����(�^�"���=�YZԋ��>�d�> �NߵX���AU	&|�`=k��t�@�UL�O hn����4�?� ��e�ӑ"`����4��y*�"Ob��0`	v���0R�P�{�F<ؠ�I5�ȟ��gϟ�^ɩ�j�����OR�t� ��Ժ����'��_��E3H��cB�Wo�*���%T@�07�ζS�tr�'R*2��Y#�:�lC9`��'L8�#�X�.~�}s�'>
u�	B���\�Y����I{���3A�
��Ʌ�U�$|�N�tZ�BX�Y��q 䊈F
�i���gy�	 �?��it�3��l�t��,1��L�s.��w��
��+D�H��!Q�n�5s�I� Nh�za��O�Gz�O�V���@�F�k9�u�E��� �n�:e�m�ґS��H�I���	��u��'�9�a��u��I���'V�8���ۛO��)5�B�|v�c�-�#yr���P��(O�)ȥMψ`(xu'ʚ$�@T�≷�Y:v̇�Ck��I��?[T�r�iV�TǬ�H'��A�	-}���D��r�F�;�	7}���Bd6Y�,�o��HO�#>Q'HN<i��ӳ%�����B�L�<a l�>�r����ɦy�^7��@y��u�4��<�!�#�?���?9�OΠ�gF�n�H��%�� ��h�#������?	��I�~�!� \�V �� ����g�-Q�ۿ78��a՗S~xu���('�Q��qH׿ _�@��Yi�́�%I3�u�+�w�����P�|����RӼ(DyBM���?�	�,9l��b��%w�HA�w�U��!�$��rꘜ8@��\>Ъ�a�%h�It����Ey"��'$�'S&)�����Y���O����Oz����#:�hV�x�NparF�9k]Z�[ሆR}R2O��D�<��_��>])��$��6����#c'�I:Zx�OD8s����I�L�1�u���vU8�/����l�柠�C��<�CB�� �I�?��I�<��)F��d�C=}ټy�B�ɶ�BT��4�?	�o���?��'���1��M��[��s����&�0(@�Qc̓(<+j �BBT�M���'�<�J�2OX�]ݟ��	�?��	�<����f�����%C���� �+����I��@Q���ҟ�j�g��D����_��y���H�A�2�)'��X����N����ڟ���-^�����O��D��H�+&X4
C��qnN)Kg%o�2 ���4t���O�P����OP�I-uo��s��΋���r'�'\|1IBl��n�8]k�HTЦ��#C�]�I⟴
��Ō�?iZwh"�'����;O-pВ&��;1hy�ؙ�r���2O�İ��'�(gݙ���<�����rش9�����ݘ ^<*F��ƌЃ_�����ybD��?)��j��O$��'�6T�U���!O��ʛ(R����� ~�����ji�`cU����] ݴ�"���y��G���4gD6H�89;��8ht�D�aO��V�ߤl�z6�Z]}2 ��b7�Q�?ŕ����Ht�H��A�`}T�`�=61!�D�U�y9���Pz��UO�%���'b2�'��T����͟��Iӟ�:�kЕN�0�p��3TmHsc@5�M���?	��?�N>I������A��:U�>�L0�*	�M�����d�OB���|����?��O�|�*pbP4SCI��O��T��4�?Q�����'�D�1tXآ��2]�AbUɅ�6�������9�؅b��R�0�NX���0g��6Ͱ<�N>�'��'�?�N�DRu��O�.t��ӓ�߸~j�I쟜��V��|z)Ox4%C7��0iB+M4w��	sp�<�D���o�.���X��ܠ(3�l�<ygǓ�]��K��	D�t���j�}�<���R�b��X��JT�E�v�r�/Cq�<1  �\��蠧BZ	FA�-�k�<1�n�4v�=���Y�VT�l�'��'���'�bK���YFF�2����@Y5�Q�4�?!��?)���?���?���?��L�RD7�W��
�r���X�0Y�i���'1B�'L��'(��'���'d&�V�	�R�n� F�H�Sp���Oq�f���Oz�D�OV���O���O,���O�<P��J�l�B��M� s\-��榡�IƟ���͟�Iϟ ����H�	ʟ���+ N�l�*s��Gv�-(fhі�MK��?���?1��?1���?)���?��I&IL��z�o�n�����jԊz����'�2�'H��'���'���'���$>�y�̳7'\|�Ф&��6��O����O��D�O��$�O��$�O��ơf�V���$8k.�1ۅN2^9��m��@�I���	͟@����	�����0^��!Å��k+�(�$A8joXkش�?���?I���?1���?A���?���d���r�˴f���ڗ��|܌)B�igR�'��'V2�'���'��'��0D�oX��a��8]P[��~�*���O��$�O\�$�O����OP���O.}�����J+N]�`�� B��֥D�u��� �	��x�	ȟt�I����֟��EȈ�>$z�b�/3v``����M#�'�r�'�ў�O��\��$ǽu���"i�Kd�0b��i�D���O6�����'�?�P�i��N�21����.Ը}X.�ZB��<�v7-^ئ�ϓ��$.�IҶN��0s�O�Q���B�Yr�dG�pB\�Q�'�,�3b#wv(�
���O�l�,nL���cef��מ�A�#�y�'e�7�F{>������ ��Ӳ�Oqzl��t
�9��'�I���O��mZ,�M#�'�ӰoZLX&�	=n!a�U;8zʓo$8���Ŝ�=iN��D�
;{��9�3O��x�������G��zj�!���N���3�lӾ<PХ,R�ܒ&&�O��m�&q���Iҟt:�4�?�,O�㟤�ȤM�}	�1(G$��ai�p�i�O�n���M���	Z��!#Sy~�E�3#;������$@ݪ���	C6E�3��L��?���hO&q�@�D7	���Y�L7K�y��<q�ifbP�OR�D��F˧�?)%C�`4F�R�!8���`@o֪	���'�M�e�i�$4�'J\ℳ���#t_Z��2e�0�Qt���8��'KƅY��|t���'\��'���'�8�"B��K��v�&�<��'0��'�r�']��;V���ڴC	���'2Hʴz�����q�[C�!����ڟ��ɏ���'� -A�I�>��^�t���u��� �t���(�a�
p���"� A�y�i"n@a�aM,V8.4Xv��>��ODh��A&��WN���rG�x�x��o�{Ʈ`��'�!2� U�b�t�aØ�&}����r�k�(��p(�v��4f���%� -nAA��xta�"E��@n��a�� �!��� N����u�!�ÌN)F�Bيv�\�C��P��L"I�Z��D���~��E���br��2(C'Z�29*Wh��Q��be�I�e��+�H]*eۮ�2�	k��b-9gQ�B䉓!��YaHY�u)��6_̜������R�Ĉ�Nܵ�� @��j���a�0�mk�KX�%ht�.Ѱu"���¢޽@��U[E��:]�gc�@�7NU�KMF-2a��6pu�}+@(�%��� ��)伣ڸ� �3��V�6�����<d]��k�,L��L���14xX�%Sbd�� ���=��u��'^�
�&��O��$�O`�O��!���w�0Q���z��)�qM�O�dB��h�d�O��D�O����O���O�� ��HS��1�0�@�ApE%�l�I���&�h�	����!�D�M`����))[�cQ+7#�@U��O��d�Ol���Ot���O����}.( �ӹT6x�@ {� � �`	%�˓�?������?���X�=��F�P-���F����G�>挵����?����?����?�������i�+8<qs�C&�f9y�%�����'��'���'����'HR�'k�m����+Ɋ��K�!4����iR��#eYQfmb4�\;^mK $�3@�q���#Lw^����
�� ��+L����%T�[ڶ�����OV�=�D�O����OD�O�`-�=�\P�Gi �J������<���?a�����?���?!7΅Ao`��%A��ڠ�c����M��i�����O������R���O�AmD	s�)E��Zn���� ��L�$��hՒM���)�6��H�Cﾡ��ߙvM6l��4���"��Q��(H��ѺU<v��GBͼĐx���y+R%�cA��u��q��bܲ.O`q�BT�>��ѧ�?�]2�w5l��B#�g���0`ٸ:g0��`S� ~,�s������N�|޵�!@�/S�(�R��">Ƙ�f^�*�D2���1�BQ�#�˒K�U*P�s��0�����F��T�1W�(�4�R�o���HB�x�`�1��OX���O��D뺣�4q�$�3I°K@�9QD�Q#�V=�CC2(��g�ߓC��52��N�S��`5�V���g�WZ�px�u��'h l	�ےIZ|�1WLʊd%�M�Ɩ�(kT���G@6��$]V"�p
�3,U@���kZ�%�'_����ӢǓ)��T3u�����)�"� ݰ]�ȓ+Ҥ��Go6���cMG)QKf����'D�#=ͧ��K���V��'/j[���
�|���"�)1p:�p���?Q���?�F�����O��tH��!0h�#7oשrQZ���EX(�0��'�'D��+Gb��8lq����(�����@{e��Rb�O��Y��@ғ!A
X��2�$����lm̙`��I/6m�$1k��¦ˈ7j��P�%��.+��'d�U!Ө�!�JdQ� �4��0	�'g����HJ�8*W���t�"H����4��td�!ꣷi��'ݛ�\�&�H���Ƌ"j��aJK�G���ðpi����Ot��2��{�d;z�f�c򌊌G�,���1I�ܠ�"��.�l0�؟E�F����:I���!N>Z�j�,�E����㖮��-"u�"��42vf�P�M�c�	5=���d�^ܧ,��|�#�C�4�J�ha�'mdB����A�r�zM���V��A&���I6�~�hBX1�.w!�$��L�M���͇�Mc��?�,�z����O26M��%����0!*z��e݊y���	�ς���^�.4�)��M����	�E�$>����U�!$d��̟�v�A�>Ӆ�g�t|g��-������ W8QR��I�8��0m�조��>��I B0p��^E�)ҧS�R��@�]���c
3�~L�ȓ,Pb�AΥ���xr(� 4��AF}��)�c�KGa�0+̶�`�ڠ0�:F�'32�'���EV�a��'���'��;uf��,��	�Cڕeu���jՁE`Q�1O � �a����%>c�D�C��n>�`0��I�uYB�3�b�T���'	F8��	!Cn���OVyj��Ԗf-`�� ��?K�=�rj���򤓃t��m���*���`� ZN��]�Eo�)����"O��㰍TN��g]/f����O�uGzR��>A(O4y�
� y����w�����>Z\�y�'�%��	�� �Iޟ �Yw��'��	�v�~�Ȅ(��SU��;PoL5>ݒ�ie���L}2v�T$3�az§�$f��u��	\<�rI��ݎ$�wJ˾	�*AbD�<�0=�e�Ŧ}q�(X)O�4�y���R|�#�՗=����
Vu�Iy!`�K�E ����!�dF�wN��qW�->>1sIɉi����O�� C�%�	ϟ\n��GB�q�H�SS��.LV�5k���?�MC��?����?y�	��ɷC0z;V�*d-ۅ|s�`�%��d����B&Z����+U�bk��Ey��P�Z�dK?l��Qd�8�3�-zD���`.8�RB^�yA�i#pf*ʓe��	��M�A�~�^��XBL ��ȱQG���x���?���ɍ�5�|���2vҵ��	�4U3qOV�=�'U���
tN�#:��I�nw����F"�by��v�7m�O��$�|�����?Q޴DRj�*�-Y�F��{���$&�	I$�'�<Q�7�	 !B�c���~S������v��8
��DD�X�Xz��G�bK"ؙ�%�)��$��-Z�2�gB(-�I�1�M���(eT�$?1w"���Qh���z�~%PT+�>aԎ埴�4i��F�';�>�[��>&Q �"��+%�mX��.}b�'da{��>s���ۡ����#����(O`��X#=y\w,la�P��;f&���@P��pc���O���O|�R�%^*;(z�D�O����O�tc�w_ܙԈԯ9f����]<�!�c��~��M�3�7*~ٕ���ħ������D�8>GF�Ɔۍb+V�C��3I~9ʐ�Z��M��n
�M3���_� "G@�Y�T��B�C"�d<;�G��Z�� c/�$E�.%Bi&OvM2�ҩd&�j�A'����U"O���L3r���z@��D��a��
_���؈��S�0^: ����*!�	��B{ ���D�,Z5���Iן��	�x�[w��'S�I�
4y*<Q�CP�*\t�吘z�ꀁ�.�lU�1z��'�⬒�U�?U���O�gv޼�PmL=a���×��0>����(�͏�� ��V �����'\��?�O>���?����LT�"�(\�`yDLcf9c���ȓj��0���,5Q�DB�kݳwd�O9�'>�ɕjŤ�z�O��Dq�<�����MX(��!T�}�t�2���ğ�)7 Ο�I����M�Do`X�"�\<M���:�S�[e
m�®�x`PXAvk�
oH�p���܋�F�<1.
N�pu�ؗ_:Ԡ��,�њ�l�*w��H&EA�|0�4��#��	��<�P���XR޴!��,�QcC
������
��L�O|��:lO��)�n��T�=8Ek�,D�Pk%��6��|Z!�O
�5�*�.�2�ҘH��(R��yy"��(M}~7�O4�D�|��l���?Y��$�t{����ǁQ�E{�$Ѱ	��f�z��GT)e+�����N�5��
�:P�O�,���Y�*:���D��/i\hK�O\���?q=ڙ��V*`�.X》��-?��SO~Z��Da @3HQ"y��#lN}r����?�$�|��)D4ְ"3�_/id�aEK#!�DO�ߌ�B��Q� ��Ia��\�Q�T���HO��#K�Q�<�*+|yd� 9��D�Ob����N[��У�O��$�Oj��S�y'O�z������6m ]�&�������)��˥��.\�R9�I|B�{�䞺rI� 
���Z�4eIF솠,"��:t��Ĳ6�^�R䰐;I|��{�P�� s��K�S����?�Q�':H)K���OG�Oׇ�'< ��R�
��W�e�l0��l����
JP�����g����#O����dЇj���5NؙH8��H�&5����!N�p��D�O���O��;�?A����#T�������6$������d2�%�OAc�$6
v
 G!e��ᕒkUL@x�g�1V�x���ݟ}k�����*�)��m���FI�f�}�؀�4�)N(��
O��K���3Q��C`Ƅ�Us�y��"O��↧I�3J�4��C7�����>�ǽi��'n�(��{Ө�d�O7m��K@`�J���h���0tnU=W���I!R7P��	ϟT���j2���6Q�^�<dmڢc��` ��%Q���� �cK�ax�'�A�.س�ÌD�'z(�ɗ �K'4�Q�Ǘ�Q��L�R%�8If�B�i� @���q1�֋\�^1�g�\r�'e�%��8���-%�t�ؿ@���a�ncrl�*A�K����O&⟢}��H��8�fH�%@ȱ?�i*��CMܓ�hO�)Jx?����Pξ�æB&�|p��%�#l�I�PEĴ��4�?������c����dӂlkR���"��@C�AԢ:� ���(���Pm-4t��2��2<�¤C� #�\�
@��b�S��r�H�!Y~
�2��ٛ�"�.��`��f��?�h�ϝiӞ��s
"?j���M�gjG�l(���֬ǋ.�T�*�P�xcч�O}%�"}��jK:������( aA �K~�<�F(��Z��H0⛿l]"`��NP�'���&��?}��EޓA����Lܦ6�����7�?���?!�/�#A��ls���?���?q��`�� �[q�Z��5���@89Lͪ�웥/Fr��i��ɴ�G+n3���O��*��U�2��˅&lD�kG�Cuʺ,��i[�Q�E�h��O���B��@������G���B-_����
S��Ci���g����,{�H�<Hq U�N�����`"O �#��Px�4B36��A+%�O�}Ezʟ0˓}��A���⢞q����V�F1L��1����?���?!Q��d�$�O��-���{�m�]�� ��d�utB�����j��<{&� )mnRT	�Z"i&����Ij�><�\s� ���I2=�)���=q�}y��>�����Y�)���I��7m�?G<>hZ1�G�h7J���
�:$���y�' `KA"O'���8��݀e�t��	���'��X�W��_�t�P�!�d�lU*H���4���z��i��')��`X��{U�^\M����F
���ƦzA(���O��d߉o�l�t��dd����NЙs�ƌ�p�xC�gIOk:My����'��)xt�Ip��;\���˰��"�h�8r?lB�N�q����O�8\��aY� =�(O�3��'���>q��Ĉ5s����fK*E玲Z�)D��Ja̜�9�DitJ������PB<��I���DN��@��҇f]((bӢv�)	 �9}� �[�6m�O"�ľ|
%`��?�ڴ)_2���'�3�dm����4HQ7��O�ض���4T����$?�O��O�$҆c��I��$`/���O�(1�NB�����"}���=����/:~�Ja*J}�E�?�ӓ|��I��iVp��a�L��!�"�ߥJ/!�Z.�0�H�F��U�3N�"vQ�0����HO�DS�B��� �x����gA"��O��$ġ2@��T�O
��Ob��Gĺ��4j����B�c��V��S x$� �*"lO���)�>�d��l@�.?�*��x�oԛ��=i3mߧ;%NG$�h�v\ ��z≣!����a8���T�۶+*��g()��y�9D�l�ĭq�����xD����Ǹ�p�����t����E��X�z)�c�0@�``C��Շ#L�	�d�	򟌚Yw��'��镰a�f��	�.:8�SA�'(�^��pkF��6P���8uC>�+1L�8ô���C��6��䓥@�4��D)NJ�)G�M
k��#�*L��9KW� B�
hЋ�D�=o�� ɰY��(IsM��)-�$����u	�����H�E�G�)M��Da\��u�'K�O������h�d��aæbR= T�>�0�i��'���S@l� ���OV7MRF6DZ�)B0V!r�M:5�$U�I��*(����$�I�eY�e��jκ0v��cq�ɶ���I��F�J�H��%�=f�𣠄����D⧈'ʓ]�ؐf��5Ovl�QB��/�dĊT�ܺl�QJf���AP��1@3�4A�����O��X8FOC5 �	+&��n�(q��'�t�4�,(�9Ka��i�ֈ��{��i>Q��'���R�ԉE�8��o�H�N�Dc��ـ�Ms��?/�B!���O�6M@pf��jw
��B��1�L�:5t�I+U��(t�Q�B��<2�@ăB4mC�,�v�
5'>�����K��8D��(�z����>��  �(���u���p��ح{1�$ng�S���b���,w�b� U�����|Jf���>��S�O�D�؀-�#r����QP�E��'� i�����a�I:��:���O��Dz�'`0`�B�^8W��J4���0��'^��'� ��G�5b;R�'v��i��0�;���36/��h���B?|\�%�<��"��0=	��:��٘���p����a
W0f-`4 `�io��c'��5�0&>�Ԉ�{�$I%���뤩�0H�Tk���+(Љ'� ���)Q�x�!ܰWT�yֈ�#6d �pV���y򏎉>u>t�!#̎)RI��0�~N4��|K>u��KĘ�:� S�J� #�A!4a��R-�?����?���D���O���b>�G�]�MnRx��� a
�E ��;,1
f�^'�6M�*:N�h�D��r��<n�����Z(�RX��AR*i��@+���q(�.Uδ��c_�1��TT���2��Dmz�T�@Э4N�^�b`�LU����5�����υ3xz,S�-VPN�bP�"\OXb�䱴eX00� =�qO�~BhѦe&}�a���O��@��Z¦��I��xoa�I� S"�X)rVB�uM�0���y�5���?Y�&�ےGR�>���JDd	�E"�XӀܶmzҍ��/a,y� BľG�"?�a�����؈�"".q�1`����|�UAZ���th�8>�\PK��&�]�P��IʸO�^����^8Fؒ$�A�}"
�'LQAq/Y >m��L2Te
�:��dR��L�QR��#���l��r w�i�R�'�������ʦ١k�+	&���DJ�^��gcʐ�?�L$+H�l��UDZ~�I�-�6:C�p2�ǝ��g�? ����k�s��4R@eY�;�. �fU���' �:��  �V,C�A�f�� {��Q���fV~leꄠî&E���ϳ���S&�6��Ӡ_�u��/�C�j�"Fh%O=B�	�!à�
��,?6D�5���j� �>���Ӈp�4����6*P&|�tk"H��}(��?��+P�̒�j��?���?1�G����-�����,�S��k.-7>]a�ǡ�M�m� 'N�����Bw⓵6/t�"�]���4��@�6��d����u�!/ĵv3�d{�4.�h4B�>iF|]$>EQ3��J��H�'�$��i�?}|t�2�R�=L�8�J<!�e���c�19��c�ȴ.W^��fNߜj5PX�ȓN�l�X���#��\qD��=W�A�Rj���S`�rF��@Q�E�WC��P$D��v�P��Ϡ.�T���ß,��ȟ�HYw�R�'+�I�	[R�#��w�6�U=[ܱ���@j���k�+��m:���0�M+� ��R��P .����Ρu��ݙ�m �l��];��A�}*���
R)��l��4_��<����¦]� B�F���4��
0fZ��ɕ"��DЮD��4EW&"�kehE�H_!�R�q�l��-��ء�ʫU[�����|�����l%r�'o�� ��h�] `�ЈT��,�"	1 ����-B�D�OR�$Y_զ�Q���f���q$�*|P�V%�
MƔ��%i˛I��@��'U$��O��S��{{~�3v�Η��E�CIɼ�X�Ѐ�1
@$��g��l�Hۋ�dE�	�n2�,iGr=�g�9G�J�s��ɑ.�C�I���ӕR�%�qKE'���$�G?�F�B�V^��kL^�,�8���p�$�"c�n]n�Ο�	G�T�q7��iߖ�2���#R�jEZ�'.
��U��m�O|t;&N[�sX�x�o�<9��)C�ǧ|�I|��h
�@��e��#{� ��Wf�l}rJ��o��Y{fo�/��0�C�y�O�l�0�/6�x�ذ�I�!	�l��Or�i��'�򟟒����v�(8�#��e���%�(kLd�p�"O6t�t/ &ZN�����)e�,����(�����0�(�d���%GL�!zB�+�O:���OV���G��]@n�d�O�d�O����M[��Ϝ_���`�ƛqI	�� ��f�X�.ǵ
���'eQ�~e9'>�aɄ87��I�d���s�?]�(�7�³T�$ u�ǹ���c&+�}V.2�J6���=!�~�y/O�у ��*c���+U:[�������ҮT��|���i/���t��B¿$b|dK���hu"�"O�d��F��2$V̸�KG�rJ*�0c�O iFz�Go�d�D�<��$J�Ai��Q��U R$J՚�F�(�l�
��T��?I���?	��Nh��O�$p>�ʶ-�Iܬ��)�w��!>���$)W�.�81t,DG%�E�pN�}�Q�<��[�U-���\�PY����ɓD҄ు\�9&uh��Qo���17��)uQ���R|Ӻ�b�7Mz���ƥW��RĩK��Px2GH��\�$�+]n���K��y���0!�H
cI (n��ðl�	��I��M3O>�b���A~���'�Ҷi�R�c
.{�p���#�}��c/�O(0cn�Ov���OR�j�3F��)��%X�Dy8�i�	�#�=P=���ED,?ḍI�i �<v6�qƒ62֢ �ʂ�L#j1����J�Z #�/b�Ҕ1*�%�����V��Ot�}����	JsP�����.�ܪ���u�<q C޹>�>�2�ѹ#;F9�ঘq��D��'�<�T�A�l�|Q�fM#��I�d�U������O��'b:T����M{�l�'Z�j��@���</Tp�֦��7���ܣ3�����	K���%񩉸|����L 
^��yz`�	#��ɼTp�@�/^
�q����.��$B�L�6V	���t#�,����:d�B�f��ݢ������7�ӊT���Cv��:�j�`���4�!��Ȫ]�^�A������x�TSa�	�h��E��gZ�I@�̢Pw~iv�R�P��'
2��]������'B�'��Ĳ?���-�O#Ĉ谋�x0�1�LA�+�,af�5��eh��d���O������)P��a�h[
c�ڹi���S(�h���%@�nߜL&�����T������'爭�Ȯke�S�[2�r��o�џ �D����w��,O���}Ӭ �E�T��X{,D1X�@z3�	h���ɒ���^f�H��X1,����Ms�iQ�'6���G�O*剌ys�D�Nh&F����%�,x)�J@�a/��Iϟ���ӟ�\wN�'��)]�1I�E�Q(H)#����Dg/`^�xFN�� \[!�R�^&�Y��b�W�V����3���z�*�,u<m����8]��c�E���9����6;IX#�⃦V(f���F�.���E��]C寍�6��}B$�0� mZ>���?������6�±D�� {�,�0�}1�.DD��(�>��_�H�:�N�Q��ĠíBC�DB���yyB�%c�7M�O��$jӼx�śg
B���dK4O=�h���[şL���ȟl��Ο@�
ȭ]?�	x�Ç/y=���Ri���CeH� P���Dc4쭲Vm��`�(�<1d�9P�P���㎌U4����8R�� ���c×���%�5I)@4��Y��<���韀���(��cav(OH�����I��y-͈C���&f@�s>૕�͸'ў�S��~�FˌjG����EЬ
��(���A���e���Y�4�?�����ɚ/w�
�j�`p
u�Yx\8�`n5�x@�
����58�Z����mľ6�]�+�d�7'Q��ħ'�8��.̍�4{K�7d���'&���)U�H�b��ȦU��;�4�B��^�Pi4�� :�8�ȢHQ$J��P�&�M���F��0�I���S�O�墔�ؓ6��9��e�{���'dЉ[ ����0K�����'ȋ�(O��D�b���"��`�N$@��$�Z�!w�(]+"�'� J�q5D���'�B�'�Ȋ輛�$z=^��D��zR��ۣNP+�x�Ӥ��z>���'DW/=�D�$>�(���4i�I<O��9�,�w]RL 1m�&7P�3�U ��pG�E��u&	�����O��2mW=+�� �֔pA�ŗa�~P�."�\O��P�'�4���� Q� �u�E�x6��[��[��!�$��l0���b���Y�\�;����ɬ�HO�;�$Y`f��MF,m�"}�D�t�а�%�6�f���O����OZ��;�?����4'�d�"Dq6h�Q�2����:!�Lͫ�aSw�ޅ3.C��y����pw��Dyc�E� �ppÝb���4�T�M���;���	W���]�x̖�����d��%Ey��^�M+�K�5����C���łF�ӻ2�B�I)C�H��ŗ�F`�<JuS/|���d1�	��lȃ N�N`fl���րu$��'c>7�>���>K�xn���L��Ӧ	�c�G���I/�+�\�S@���?�ȗ�?���?���+����yZwӺEY׭ű�X{�_	|�2�C����XI�ݱqÞ�*��t�ˑ�y�p|JW�%}�%�'a� ���KC�(D+�=�#I�Ɵ������d�v�ҷ�!{>����yrk
�v0yD��t�ܒ�D� �p?i��O��@�烊[��B
2���В>�4b	+3���'V>����
���lښ<T�@@��ߎC���I�D!�0���lv"U'�R������1h�q���y�p	@J|
�͂8b�j��j�u��#B}���O���0)�������+~ۆ7�_�7&��7Ű?�։�hZ���Sn�A�<���>��d_�Qܴ^���'ۑ>32�	� ������c
�)9�N&}�'�a{���)
�4��� U�������(O��DPV�'cL��4m޹��iՆFX�.M)'-ʩL�B�'.��
�Vx"��$�'���'�����V�{�]I�BF�NА{�ʎ�F�zm d痍Epys•G� �&>���yr�O�{�����P:j�YЍ_)�6t�P�+��Yk�V�7�&��K|�5��ש&��"d#�.RUb��P�1�|}�'[� ����?����w�F���j�=� ���j%p�!�'���1�.�&d4\AXP���g�$}1�'��"=ͧ�?!+OHy�m�/�(���.e�HI���r,�"��O����O��������?)�OW�
ߴK���`/B	-�X�BJ�(`�Vه�	�L��7[��E����`��2�N�a2�$�MseƩa��a������ĘpA!W�bB��!5�B�y�"Ǫ�q)7j�b�B�IR�V�3��� �B��C@�2�'�b�T�s�8�MC���?�4w�|8�uUJ�qc��qj�r��'�Hq��'<��'�6�Y`/AD�X��aX���)G&V� 0f�HTxI 	��f��i!���(O�  &	H4h�`S���4f�BeL H��Ȫ�,�U�F��ґ�<���nE��(OXd۷�'�B�>�J`��<N�`��h��y�n̛�G)D�pXR��P� <��X#i�L���h:�	u����j���@0g��o��Ń��?�\��Ub<}B�`�7��O��ļ|&���?ش7�HM/Y������_�� L{c�'����r�X�CS�ʹ'���k��/�Bm`����䓳l��CE�M������n]�����1
�ivG�A�B�j�KW�;����&'��LC�:Az(h
�-E���'��)��C�ɧH����*�"ƚ�B�a�#*��y�"O|S�^(x��1awAS�fݨ�I̟쨉��OF�,3�.�:MM A��ː.	t}
c�O(�d�O�s��B��d�O���OHy���!b͊��MX�*�+`lxx��D�������� u;����w<�����5L��䏋:<���f��"�e��C��Pq ���D\��q B�Ԧ)�"�iL�F=.T!+O$�pc�$A�+2N�29
]ZP�x"䜘�?)��'��5�+:;�z[����J�'�|ɢ!�n���F���$!�1Z�
�O||Gz�O��'��5A��L1%��U��ЗY����J�r� |r��',��'~�l�A��ɟ|̧	:!+�B�4b�5	Q�tQ7A�6aB$K3��I{�	��'^8}����+�V�2C=n�B��!#ߺI%� 1��6$#ў��P{�� A��qjD!v�ֺ��IÀP�PxN�<`�i��d[�j��I2r���y���7J���!M6.B���+:��I��M�K>Y�õ}&��'�"�i6�����ds(���'Z�{�!AgC�O���t��O��D�O�Գ7��b�I��u�r�j!h�k�n��rFӿs?:�[V��3��ak���0�<�[�6�K�G["��-t�!W>ni	�JQ"R�N0"P)ۀv����a̷-��%jV�	>5�n�%�8JVj�Oz��}�G�%i���Fb�b��(u�Q�<9E�.=w�Y)s��zL�s�Xe��hO�	N?w��*�\����&	.92�d�l�IP��䧦�JHQ,�c��Y4�<�R6��,t�DE���K&q;^����N��i)	2��I<�����ӟc�nI�Ԏ(%�f�@��
1y��ػ��$Ɔ�J�L*D���ЦL2'�|5 �BR
��)kç5D�H[b�7��I@lĥ���k#<D��BT��b\�urt�F<([�cA6D� �R�9;81��4\�t���H1D�,�R�+�BdJ�,�钆 8D��r��0^��i�� ��&��S-=D�lf��?Рa���A��$0R��>D��@�H�1X�T�����s2���&D��˂�èx#��c���O7�*c.D������$3�[��)>����"
*D����]�U�()�a^je�� +D����,E+V٪|�$��WDF�	��<D��ѤQ):�h��T�PV�x 'D��h��G�
�dPȎ9@_uh%D�@���@"dP�Fg�P���&D� ��-]3!��0� h+Hp��&D��0��0aְH��ɜ����E%D���Oӆ[�de2�A^2t�ة�GJ,D�`A�Y ���6�D�2��+D��#$��pFL j%�K0�&D�����a�x��(Y�e
�KS� D���r���{|B-�&읳�V%�P�4D�`x0@��:��xC`FJj�
��5D�x�F�vN���FN%ZK��;��3D��
������rm� '�`���M,D���� >��d�T-�V��C�9D�@Y H�=HR�tGg��13��"D���A�C�W�,#$�U0�`=z@:D�XC!ˎ�Yi:ls"	R�_',HJ�'D��Z�@�W}�0��V�^	2p�>D�dA�ꉮD*d���W3lA���G�9D���ƫp_\!��n��.����F)D��D�@�Z�l[���6��]���5D�,�d���i��ܛCQ��22D���6�&W��!$�0G�K��I�ȓx��,qN��z!AwA� �Z��ȓ5FLU����L���$)�.���XմqIᡒ�QB�0G��f�fl��M�H �o
6��qؠO	�{�fԅ�TØ`͊�e�Pe�3�p��e�|��`�eR�!�&,K,�Ʉȓ(�̍bӬV/z㲙6$�);���ȓ,t���EM4��S3H��O��h�ȓQo�0�ƈ*l�4*�kW&h�:���d��S �Bn�!��,��v���9g�]�Ԫ��u�|���A�q�ȓC"!HW
0K�ZE��II� Έ(�ȓ0�ؤ�AE�>X��+�KD)�^e��zx������N�Q���Ȋ&�%�ȓ�x�W�Ș���S-bl�q��n2�q��9�r1IS+M�1�$��ȓE�Na���:+*z��5Ҕp2D��S�? D�
��T�u��ju�W&,6��a"O�4�Ƃ���@����'r�|iCb"O\�3(L"x�0� 7�Èi"�)�"O�����L?���"��w{�q""OBI�O&m�*a��/��`�4*�"O�������rnԒyV^�[�"O`P{t�<�,}b�.O�CN�u�0"O�@��ɚ?����-U.��X"O8ɡf&�Y����띩��0"O���B*`x*u*֊`h��R�"O|���鈥I; �����#Ȳ�"O�qc�l���	ǩ6;�%�%"O�� ���c^,���-���"O��Bq!߷a���Ag��(��"O ���/�"���� �&��p"O��!"��`����T&F�Vs	�"O��S鎤`b�8�돵AK�`r�"O�isl��7����a� =QV �"O~�(���'+e,��G9�r�XA"Oȡc�(ka����EQ�/f��f"O.�9�;R�x-�2�@�>4!�"O����jT/+(�u`�Ұb� �C&"O81Aκ5�9�@K�Q�*��S"O:��3��*{�}etJ�pa�"O1�����U��y%�E%��y2"Ol5[���@)"�F$.�j�!f"O��ժ�6<�D�a�R�@D�p"ORi�AY4C�:�
�Hߺ'7j��C"O41��&L�T��P���,�!�"O`Q�3�������&�� ��z�"O����E�"	���ieŖZ��xCw"O�����(5QP�����?��`�@"O��i�cį.�<�IG�[�0����"Ol4��B^�f
}���T%�p�Z#"O�U��)\1�D�v���4Ҟ��E"O>�yr �60w�$�#	(,��"O�Y �"S<��IGAM=oaHd�e"O�) /�$����w��+���1�"O.}{vƈGJ(�萅_�$DR��V"OV�6J��4��v��,=7�t�`"O���MTk�n���OTa
�
�"O�\!��-l~~Hs�C�����"O2:
+��͑�N�D�|ȅ"Oz������F<KE-A5;2q�"O$m�re�9���h�f� %9�"O=��(S�b$Xd�ӧE"O�(ZV���2�{���	B �Uх"O6��c	�ㅌ z���F i*!��x:��0Wd�g҅!�dM���YrO��m�|�H�-*F�!�d�6�෌H�S���T��O:�� $�)�iI�#�~Ļ�@�+�l���C�!�$�2<���ĄW�G̈́�+�<1��D�	�(��	k T�٣��>{~y��d�;|�B䉬R���Sb	E9RaN1��"B�%�"�2U��8 �V�����`�q��J�}����`��I��z"��?�6-�'|�s���p�Ʃ�隐p�,��'�p�CGȼn~ ����@D���{���"�Zم�S=3 rQ�DV�<X�PSwG
#M�B�ɋ?>6ɛC�E	�ư�hH8Ec@���#3�	"3'Q>�ol��6&6h��Q�_����ȓ=����nR'[/p��c�V�G�yl��V�E��I�Il(���1~��Y	���1A?�����b�up��.װ]P� r5�]�QA�h��S�? h�8�Չ)@��U����@Г��@��(O1��a��oO�Xm�� �B�'�4H�D"O>l���̞r�~t�a Z3,�>�y��dP'8,�x��J�w<R#(Ђ˸x�ƂC��x����q2��!eN#P�u��CU�h��q�ƓD�v���
z~�E�a��(�  ���a)�㟀*�;="ݸ�IG'�8l���*D�(���ҢS����p��

7}2���O��B�
:n (��免$��Kg"O���� *h�<x	��F���$�G�����a�4U�C�U,Z�x��2 Sj!�$A`��Y�pO����1�f��.wj���$?4���f�_%5h0g��a>DJsJ(O@�0�!�	s(�CU�S1g�>]Ӥ�	t�fB���p74��`i%IўyB�	k���}�&�fe��&�42�Y�$�j��9!�Z��wd#D��; B:U�2tT	D�-і)��>}"�\[�5{@}̧]X�9c.�F�٢����-(��1�R�a�OB����L���U1�h*�(M�l1x���0!�<�1K��	K~�<����)*N��c�[���rB�Pr�DI1
N�	2!�8�'!�q�`՚Rd���i���)x�*W���(Da}"��0btt�G΄h��Dm��$O��O�}�%�=�0c�еH	�	ӑ\'r���)S�t�h�f���,~!�dݥi�q��h/]�a��X�=���4G7r��(J�@���)��Rt�	ЖI��˧Udb%�V)�7�X�pȝE�ܩ���Tgj5XE!
�E��1��*�"Ov�`у�(R�rd�[æ�C�	Η(p�PJ�~�>�oT2N����
�nap,iV��e��a�Ǎi��	%�V=@�I�V�C4�5\8���1\
	��IT8G���	
!,Y�#��Y�n� �G$�^�w���hO��P4I��|��QN��~�Hk�O�:Q���
�U׼hYa�'>N>l��'�V����l.���F')�FŚ�O�h[�A.-;$y��jמY�Xu�OQl|�2[>��/���8�$�4�M�a�,�|@�oT�|�|����P?�Z��ÒU?TI�w�&_ܛ��V(U bJ�i��Q�|4��ʀ9�0�f޻	G�x�@�8��"�`�PW��?Wj }zg�YANj �G�'��F��s`�9�7���GjZ8?���ćЌ^�.5%�D!t�/}�f�j��t���SF4pI��4��� �b*��h�Dߦt'�|1a"O����&�(��J�HO�.d%b�_�Zp���>Yz��5��#0�b>����?��U@]GF�\�q��4A*��e�?D�LA%#Z�B�
Pj^�!!���QH���QM�!�~�(�	�z"EL��$�DH�YU�]�R1���#���V�z��4���%U8��2!��!>�{�"O"0"|1%+.�� �C/�O8u�gM��W	hqr�͛ybp�sw�D>���[��pp�&���f�4=0ӨC�:�r���fd�!��<�n h"�B�^�h�pe\��1Oj�P%����O�,P���
�vVb߳-���'�X嫃@D2|��M)A
#F��
�'B�pp��!5" ��I߭;��
�'�4���M��� ���&x
�'1��@t�N�$�B\3 Wy�����'&.0�d<WA�p�!�h*���'�zɉ�HG�(�� ��@�Wl�� �'�|x����GE�$JAž]4���'ǚ������i�%�sM�$Rj�
�'���Ȗ�N-�̵�"�(#��*�'V������2�����(��k���[�'��4�rB�h�Z���A06��A�'w�2At����^��`a
�'�V��D\�������7f��]�	�'m���5<I�Pa��P�OT��	�'���K��, =��pB @q�D�'Ҵ}�rCA4��)[��(0��=�'�Q8���Ό��46"���'�(��E$�~�p��u��%2�����  jg��.{r4
�#W�P���"Od�z��D�^�G���:�p '"O$�ꅩ����a�"_����*u"O��*SL�8��\�&AO�D�i�"O,4��H����t@�l_ʸ0t"O~i��`�o!PnE������c�<q�
-���;�oG�/�z	�3Kw�<Y0�گ4��M�Q#�2��u�CJ�<�pKU�b�"��ဈ�F��r6.�K�<)�OX��*R�C&*�%�w�6D��"��UM��reߘ8�ޡ*��7D�t�2��7&`഻F�S�d��M� m)D����?*x�}i�JL(�Z!�0�'D�􋑆бFt0��vIQnik�
.D��rR)��D(Q�Q2��B1�:}�B� c%04�u�C6{Xp}��%���'O��2��ٽ<�PS��	�F��'�J�U�ĊY� ��fT|~n�:�' jl��� 
�h��G�ݩ�'��H�gьrF�L�bB� v�)�'����dd� VrV�J��ǖtq�'�0a�C���4	e�(�Ȍ�'�N���S�>Ⱥik%DS�^���'H� 1�̏,eT�9�t��0��	�
�'��As���jc ��"�L�,�.<�
�'L:�"���\�7�?)O@(Z
�'�`��F�-0l�	P	���8p�	�'St<#�N_\I9~Y��x	�'΢���^�&�êZ:w��]��'NB-8@cA�9V��cQ����2
�'�v�����-��}�|Y�'&�9 B l(jY��5����'����jF�*�3@B#-���i�'�`蒔ƙT��XA��se�r�<Qp�F]w��C�݅r$R�8��El�<!	�2K,��a�E�o����c�<��އy��eD �AAP`L`�<�@��Zp
 ���>O^x$��FHe�<є�Ʃ2� ��T�R�m��� a�Dc�<)��"/� �t/�|�p��$��b�<q���HN����?j����X]�<aa�_*`A�r,Ey�T��Մ�S�<�sN�!�T���kh!���
L�<Q�Č&4��)D��"?v�(��N�<I�m*���b�!N�By��k�L�<y!��3 ��0���S�<�����4cA��0O�㲂h�<��݁O���I��B*YlU�gCc�<���r�����
#3fp���_�<���E�H�����KLL�|ؓs�[�<Y�f�,xr�]��7iBb`&�A�<Ѡ$����8V�(p�%G{�<�׬C=u�:�  ��5�,@��R�<	t�L5R�Z��"��|����o�Q�<)`��N��aa�����ݟJȬ�ȓ7~����h9$�����^i8������z�h�H����������z�t���V��5�H@�d���	����#띪=@�'+�g`*M8t�6LJ�i �%
�?2�➐��	��+��S"`j���9+��H;%	
�5=��@㳮W�@պ�R	2�␓rB"}��9h���� �/n4��N��M#ϲ��EB���� �2��B��� k��Cw��Q����ˈ7L�v��ԥ�4��`�ޫO?�y��d7�ԟ��x������ȹ�"�-���n�@>92VT���mL;�"?����J�K#�$;T�h0ځ?^
�OT�j4*�)�	Je����j��(�jQ�1@S�w�%T��m8��AI� =v��{�? ��x��.c�MI��8eζ�*#�Ȩ��'��c?)q��?��uk�5L�:�Bcl��w�E��L���������"+*t����2��)�O銣�½	�V�; m�O��A���N?��j��xxA:�	�Y��O�PQF�̑Q�褻4-�9��XTF5%D�1�^�S���w�h��5�U.>�4��VQ�Z�q7���M��/�&^� (Q���`nF�a�/XK�'7�0�a�!
�z��^�d�z��q�Pi�'Q�����1_8D "D�X�p|��#W9/PX�	ǓPyb����_��y����bd��P�H�R�<���" �ē�hO��T� `���@
B���fO֣A�RL�u.S�*�=�?IT-J�'��q�Ŏ�J��$�LF����"�a�b��H���A@��eB�Ojn�a���T�6�E(@'�)ѪO��	N���� �/ݴ9E|e7�]�0aT��D�],"|�L�W�G���O���3_N%�F���|��#���}x�c҉dW�UӒ'�?!Dr��0��>	���R4o���R���M��hKT�#���~�j�p"�Ӛw@d���M�C�%��5�L�(]���䆤`N�jd�z޽蕭�3ݎ�b��!#�b��lىZ�J���~Jx���\W��"fӔ,y�#K�+t����0i�4��A���#<��V��I9�'T3!RXh(���n�d	qr܀��� ���r%�%*�F��*k�H
��i.BM�Rb�Ca%	�M[�Õ@�I?ED:��/l�p�j@+FcQl�QP)Q�#X���B׏F4b�2��F!�b�I�D��Ͱ�d���V�!E#-Idh��شYv�l�wĊu$he�%�U��`E~�L�;Xv���e41ٳ�Q�3x��=�A���~��O:��5��ٔo�p��)�+G�ىB�H6i_�L��7O[b/cY��]�rb�=��H����=9�rdk�&�a?��'t���'(P���+JqqL�!sF ��ӠV�X�YQ��[k�0�G��n��4��Q�0��d����+Do��U�R�ņ�fR���O^mn�=Hk��G�Z^F<���t����O~͘rᛈ`���� @/gz&���Ǭi���
2F=N  �p�o���O�\:V��09��Q5��0���;w$禽�4+�T�#u2y����He�'�>�nɧDYD���-��m�X8j���^�'��K4/[z�i�Y	Bm�	�4�B��I�pz��@���`Tv@��f9� �����yWd_�H�P�w��d���u')����'����R��TlO�\BA!��\�otڈ�Ę>{\ӌ"h�+!���FbQ�F_��+���ɗ%O�����>�,���QTOZ�D�O�����B֔��c��%P�T �&R�s�A�J��xy@O�5YPQ�a��G��������G���Z�%YџxPB�o���u�.t��pEf
2�M���4V#ι���.�MCb�R�'�x��$�4�Z�IV��##)>�0��o�'S�O~�a��	Qt鳤�Im(�bu��YV8���'�x����Ņ'���#+�t07�.���F(s�'���t2+���LռK�u�B���I��E;v*3j���;2��T�8��В� 9�ȉr�D,&T��OJ�`wKO�7)}��<|Y(G�D+67�%x�����?��ȇeܓVx���l8���8@�X8ch�;hn����ݦs����sV�ф��p<�эe:������C����ׄ�ڦ!��DW�\�r1�r���{��P7?�s�	+��/%�Vx�q�,z���1C�!�<۴
I�E�3G'/. K�'ݓ+�UY�T̜���$ž�y'oj�¼�"�I�P�c��H���>1�
��d��L�G%D19�ޕ��)����Sk���Ojp%�H�"�D�)A�CN��p{5�>�W�Re�Ȓ��(�:ɀm�c�'��)���rD eK�i4 dA��O�@�7G�@�0I�i:��$� @t�yq��Ls�՚�kٞ	�ax2hP�0p�h��D�*�鋏�BD�#7��JP��`���5��:-��E-�R��	a�WRD��O��e�G;Ď�A��I�s5�Y!!��v�hT��iϮ%�a|B�R��v,�!A��Z��@���ɐ{�`�1���Z�$L��^�j8�4�ӈu�⠀�G�� �GA;N8b<�m6�I�'��H�I]��=Q꟢6p�'� a��*I�n��Xd�I,�	9��D�!��y��]�� 0�VS�ɰ �u���6_a��@Ru8	FII7=�|m��O)de^Z��'�fm�b�Ό\��s�]��h�ش٬ԛu�_�δII���D~�M��f��0�� �i���ɀ�QX��a�ҝ��@�e�U�S��hX�B'�	1��xR_1&4�`s�7�a�7��-x�kE6��[�'�*��(�5a��!�D�(�:�q@��
1�P8p#/��>J�n�Ct��#N�nt��
(q�b�'v���O��b�����K�|��=	���Y0A;���#�I�	Y�qX�TV�Ii��Ի7&ʓm�F��6�%SXēBd^�;�=�2d�*�}S6�'�%𗯀�y�t���Z.�X�ߴD~��7G�\  �W�U1Kt�`E~���1Co�Ղ��	�/{$9P�+�|��ERNn��I�?�R��Y5�E���27H�����i��Q�'H�!�JT���N2������#0��g�(ۉ'�`ɧO8��O?�����-��7� �Y ����y(\uv隣2rh�b�D�,���Dh53sP��&����r��A���9L�6l�P��Ō��''�`��R�p3��L�б�I�M�&�SQ}����X�<`��G��0{@�k�&�B�9������I
���F��q��ɪ	"��lI�	��Y�#�!�>6-Q�v4�,k2i�k�` 1�ǧ������E�(v$Q��Ѣw1���0�VyX���W��A�t �_2!�ÉF|�x�` t8�,�H��N�\λx?b�kA��<O�=C*I>j�Bu��I�<TX���W�9�.3�a��G:���BV�b����R�=!Tl\"b��&9��k����3ժM��@O�A�@�
Kj6�JU�M�t�o����@Ğ��ѳ�O�!��2�l�v������ B�:R�-��A�+��"ؚ͸'mx<�O��NŹ�h�����b4�iu��:��-<��f�Q�9ˍ�D\a>x��Η�J��XU��	�Ą�{���d8��#m�+mnxq�'H?U�5J� Rv��
Ǔ" �RPM��ye��f��C�Ǜ�"��:P�Ӽ��>�q��9���d�D���p�+B�S���s����\��Oْ�#�
	,i�jG�'$���>q��O�abA�6&�=:�HHt�	d�'� ���/ڭp1�|j�>]�$%8�O|qh���j��x��O�Xh�a���Fٮ���gΫ�����A:�p<a�`�Mvh����C�K�X��C��Ӧ�����w8}�v� �0�h|zƆ1�)�x�PJ����4Ɇ�K�]�L��ƃ7�u���� ���(1�'��p��ϖ�Ib��N�XKt��y{l��$�z�b,�M~ޱ(Qk4G(����N�y�`�Y�g1���X�P��8Ojl�J?��5n	��J7̻F�\P(	L�z�̸��Iͱ8��O4�;/�7ʸ�T�XusQ�>�b)��2c�\'�)J�DË�R!mZ ��D��4L���f!"MNb�L8g���\�l¦�V�Zj�tRa%,��x��d�,�n��N_U�PQ�Fg��l�Q�l���N�J���Ӷ���D��R�$A�,ԩ���MJ`dA
U��#��R���Oj�e�M# l�4'2�^\2 �V ݨO6i�6ʦn3r!rc��u}�GJv��I����p�@,bP��!E��ebc(9O  ��Q��ݓ�a[Qa\I`�8��B;�8ʓQ����h�el ���.�+��!��얤&Zr�*��\2�(w�A�u؎�9��ˑv��fE.i9e U�H���J@zh+�b_;PĈ��,�fY����B�"�H�HY���Cc�%����i��E���|}�S�� �0bt�B��	A�83�)�=0�rm)V�jĚ�'���OfI	����v��]�L�A=J���j�..e�Ihu��5z�ү��;.&��Vw����#h�P�T�`ˡn[<A;1�R��'�<@95�'BVQ�IA6���3�瓅t*@E�0@Y�����2��P#$XJ�
D��p<�R��K�@���w+��Qg�u������ ;��iz�J�0[��F[N�!H��7k$�K|`O�\%��qĨ�yw/k��h
�����'a��A�D�#>c�P���NVV���H�xB�)��Z{p��e�O�9.��$��7$Z����6�M-C�d�؟p��a�W�Y�jȪO\�"!��/_�T�Ej���թ�ʅRr��!AŚ$�Ku I�
/�S���7nܐ�qkK�u��`M��vy��+ņL�6�X�l.jt�i��^����t��vN*��C��� ���c���e@B��%c#�ʢ�Y�TԨ%���Ϳ.qFB�xx�r���.�.�ۦ%ɶP*@B�	��ݻbKW��2S��
p�*B䉿W>@������L��hY�\iB,B�	t�T3��S
���'�>�B�IM���Ҡ"P0V%���lB䉣��I	�O@/H�1q�N'"�rB�I�wJQ��/b��� A�/��B�	�qbd�a����6��s֏@�n0B�I l�@����M�n�xVh!�$�9R%vI���I4��u`���+\\!�$
�@������Y�� pc�;Q!�ՐkU�H�Ն�p�P\HDM�-�!�՝���"#"!��A"�S
X3!��×@k -qR-�8�`���K�o !��-/���6�Wod$8�Bjк>!� d��Xpg-�.nJ�𧂂�B�!��L��m����u���� H1{�!�$Ǔ/ä���\++�`Y����{�!�[:b����!�L s�FL�r�-WS!�$�=o<.�kP>>�|P24=!�$VO��PXd'²1�`�rj�3Z;!�D��1}���v�zĲ��T	�|!���+-�d `�.�r�[��3ha!�� ��!�i��#��г �
�'aXy�""OR�!뗎5q�E�M]3B4ȋ�"O5* "�	tȭ7�ƾ]Q�{�"O�d��&J"�"�Q�%G+^[J\f"O�f�4j?�@@֫��A̡PE"O~�DBR�T�p�dĎq�v��"O�� �%8� �@g�20�"O<�ۑ�e.����P�z�Q�"O&����S�#w:��D�o�ʥ��"O 9�d!�v4�ǯ��{�nt��"O�%�CgF��l)�A/W�uQ�"O<Y:u�=��	��M:{{��"O�p�&�	o�d$�gk�AfN���"O�(j5ǋ�i�EK
P:8q1�"O����	�\@��� d!ֵ�e"ON$�1��B�d����ܦ��ڶ"O��4lI	5���q�Ӭe}"|��"O\�QG�H��B��#hvtЉ�"O�$CD�H�s� �5+��b��"O�ݫ�� |[�'ܻ^��-��"O���K
 ~�[����P���)�"O��1��	eX���N�D|(�0�"Oʭ��&���s�lG�Pjn�a�"O�I@���M(b����F%qc��1�"O~�s`_|܍�KD�+�d	)�"O���O#pw>9B�
��Y?��"O*�v��q� �w�!+ �Z�"O�es���an�SSJ �	%Q�C"O����Ͻ
�34I܇s�$  "O�1����9m�R���Bf�ika"O��j#��?ָL � ��xU"Oވ�&"��\H��ҸB�!�a"O2���ţB��ģ�B�4Z�֑ٲ"O:̘c��5��0�У�$r�=�q"O��(�U�_'r��(�,c�X�"O8D�'cb]�mD�G&K^��`"O����oJ�a�$`��ً@�H1�"O�ݑ �&�ΰ�� uк@�#"O~p��◪Ff"5Pd���q�`���"O�,�����hxv�d�	�2�k"O4���/�m�  ߡQ��0�q"O��{�	�w�r�
��8k��(3""O�i���� {]ƥ�3IKy���h�"O�
D87��h"T�N���I�D"O֩Ǌx��0�d �/ҴxA"O��5C�n�12/�W�Nu"�"O�\�C�t�ܰԋ�Y�PS�"Op��!O�
G�޸�d�ݸd���(�"O$I������D�ŉ��l����0"O�,#!.�n�ĩb�J(M�fШB"O��/�oj� Zv��7Y|�1"Of8b�Fg� ���S�(���j�"O�Qp�b���Q%�*�n�y�"O�<BpD�_�IX�0���js"OȬ��CS�I� ���R�eR����"O�B$OP*P$<!&���Ld�D"O�t�rKB�`AH�b��6����"O
��U�9��%ruG����6 !D�<�"��7�I�ah
Wʦ���4D��r�R.�|D����`s��j�0D����

-������/�x��2+"D�����,�|�*�΃_1�(�� D���	�*�4�*��/2L�� !D�(r�)��X����.��x�0��?D�� VYB'GU-V<~����	gxY3"Ox�p�l�yb��`���T���"O�pã�+�X�#NV.�j�{"O�D���	+�-��L.(�nV�t�<Y�(S,�E��j��,e�5��+H\�<ٱ��l�04�v`Y+t�@1BUK�q�<�C�h�Phv(V&x<d��n�<�0�K,�|�g�ˤ-�^���o��<�D-ǟے��@LA O`��
��G�<��cG6Ds��c��J�ctD�2��Ak�<aE�
tؔR0C�*q��p�u�^L�<ѥcی)%R-��Ƅ�h��i���VN�<I Z	�e:�LC�`R��ۅ
I�<��o�`��|)7��0Z�Uz�f	E�<�����9H�pr�O^��D�D�<O�>�h��fş�?U��"�V@�<ië_e��M(�W�o�Ha{�g�|�<�4��;����eC9%����A�z�<93��҄P�Q"�5L�8�C��x�<9@dH�K����iI3e 	��/Zv�<�GƆ{�L��ĺO:�a��A~�<�!Hr�#�AM8O��\��CX{�<��'�[z��Adi7qjL��-�k�<�T�;C�X�����6�"���b�<����+x��*"��|�&�i�w�<A�����D��*�o(p���g�<�����5�H1!�Ze���T�a�<QT+ǅ9e㳄�F=��:#�H�<�W%B�wfQ�͔�58J1jQ��i�<)L#�*�P%E�'t8|�C�c�<q��PVƉ��B�\ɴt�4oG�<��$�bA����Y�r#�D�<�H��
�ҁ�@8��= 2k�@�<A�#݈AKj����ݔ2DP0e��<�cG�Mɘ:�!�霜�C��f�<���H+batPt�SD���d�|�<���Q3�(����QѨ$P $�\�<!r{@t��2�:Ѫ@��)�n�<�Q�ߥ�x`��շFx�!`�C�<�1c��E�Lh
1�6El<�%�I@�<�JK�
!�=Ha-�0	�ޤ�"_c�<�5"�M�q�$��	% �9��Q`�<	�ʓ7=hLE�"�D�;㐐)�b�Y�<���
�U�g!F2�ԝx�q�<F�Hm�z��F�ؒY��4��Dm�<!t+Bxk�h�-d��j�<��j�TP2aeE�9jfQ�ƅXc�<�����A@���&Bώ<�*X:A�Pz�<!P�EuxN�zphQ�7ֶ,�楏L�<	fD��I{���"IJ�eH��ł�O�<���P�BQ���WD�9�H�<1��ȝcY��BqC�Uj�����i�<i���GX��0Q#�Q�ХA��Nh�<���'@["QЅ��~�D�d�<Q��Y/\$��*V� t.��@�]�<����(��ʁ�� ��h�Q�<���[�d�s(���k"�r�<��!)E.�-��e� MF�C&�m�<c-�o�T��Y�z�T��M�<�U��8d�BP�_�t�����p�<!�;����	�U�6y��eED�<ac	ԞPZ����aтrWG_A�<�׋f�$l���;,O������~�<�����x=9�K!If0��A�y�<� ���hT������[#�7"O���
��|p�ūL� ���"O���wg��f�T1ta^�<�P�'"O�Ł��S�
Y~ �q ǽU粕��"O�Yx���,uL�B6�#�b3"O0T��'�����4E@T��"O�����K��H���9F	�M��"O~�{��ЧI��3ì$��L�"O���RC�8�8	�E P]����"O"(�#�C59Gfu�'DT�3@��+�"O���޳p�*̠�"_�f?px��"O9¤�)$zr�h�NS�Z�"O�EH#���]���1�͢$2�ͱu"O
� �A� TvLmZ�eYs�p@"O���#K�ax�����W�L�r"O��@*��f��� �=E�b�c�"O^Y8�'^8a`��S!:�P��"O2 #`A��DT�P� 28�.H �"O�ۑ�_���\{5NP (�#2"O�=�c�^.e���`q�%\PU1�"O�@!2.M%/TLT3eD�	3��{"O܋�� �p|�#T*�v ��"OLT��&J�5�ܹ�e"&Dפ(9�"O�<ۂg��+�����Z?V"B4K�"O �ū�)&U�0�C7N�M�"Oj(�o�PDs�B� �r��"O��CB�.�,�y���
i�4��"O�Qy�JM ,��q*�B#��q"OTII'��F�SD��R�(�y�"O�x&��	e)�8��A��rI~�+�"OZ��B�'	�mA���|��a"Ob���["���T-\* ��x��"O�-C1��$k�����LN�j�0E3�"Oz�2�W?WR(�p
N<!~����"O�ْU#ǈJ�jUi`�g��B"O�,�"��+����N��E"Od���EZ��ᷦ�\�^]��'�qO �[�O$s}d��ԋ�<
n5K�"Od�"�EH�-� ��%N�֩8�"O���C�&���H���-��"Ol��)C<��(�C.ƵK��Y�"O��tꍺeY*Q�D��e�$tjP"O���� �,�d��3K�21rb9��"O�0���8%i��kQ�K�1"O&�R�����#�'YG6!�"OT%YǊ�OZ�"�:`�Ɋ�"O���e��z�b�qa��6!U:�"O @���H�ne��P
�(EA�!J%"O��X�FTz��Y�,��yLD��r"O����	�8X\�k�
��`��b�"O�=!���,�!u�#�Tz"O$PS�̗�&�a����T�h=bC"OZ�V�Yy�����:�2�S"O���J�11���HS?���I�"O�9Ӧ7hX�����+��	�p"O�9;R��+
�j��6��"��ݫ�"O�m)�"^�ch8`�@�
W�VEQ�"O���f�M"[��YT�p����$"O���˭4�P!�s!���6s�"O�M�B-K�-�^���Q( �l�q�"OJ��Rq��@�ԋ(����"O�w♭
�>��W�@w�%��"Ov�*��W�j+�Š�l��@Mp� �"O��a��XtC���ɇ�K2��+�"O� �a�"�\pQ����(!a�A�"O�����L��pVh��i�2"Oƨ(���}x������~��q"O8Y���-,�9�'C�����"Ođ�%h3s}�1�sȨ&M0R�"O�4!�(I�PnzDY���m��ٚP"O���e��!�(���6%Z�
7"O����02gT<�E��l��	�&"O�M�6���f��"�߼A�R��u"OJ4a�߂*�|q@������	Hb"O\uKtg�x���F&ē��}t"O�H!AO�[:&q��gןYŔ�cb"O�iO�*XP��3+�l�YR"Ot����]3A�`��_8!�����"O�bpL��kEH,�ڸ�-�u�4D���G"�7nlؠ[%�I�|�L��D�3D���C��)<>�T�R��*=�T19��,D�L�"¶?G�լ�	,a�4�V%D�D��eZvۊQh��I�%��l�Ё"D�@�Hҳ�F�q���+����e"D�L�F��z.2,��E��كp�+D��q��+xbi���'����+D���.��9�.�a�/(�䈠`/D�� 6NЉa-�VRE@��-D�l��d�2*��h��H�ܨ G!D����O%4��	H!i�'���+v�$D�����/��m��
	����+5m!T��QFՉ"Z�uP�%��6���"OH!ȡ�Őx�XV� �62x�"O �D�Z�?sܵY@�E-�t���"O8X�w�Y pԢ�1�(P3�D��"OP��"r�.�
ŦQ.~	"9�6"O6ٰ#��;.���8�@pp"O��	7a��lf�=[�'�5�P��"O�e
T�>,��E�2��7"8I��"O2���f��+���q.˜VFX C"O�t�'����8[d �N����"O���ɞ{��%��)�8r��U��"O�#���g�5�V�Q�Rwx��"O ��2n�0xؙ"�à
hL�J1"Ony�AA!��jE�-]��"O��J�j��c�ERܙ�"O@��3�фb�v� �$��_���=D��� ^��aR&��. BY�w�/D��W��u*�I�#I��~�a�h*D�P�����ʬ#���4\�z���(D��k�ZES�e�U��=7�L�`��(D�[�i��4ۂd)2L9�n'D��b�ă0��u�#!{�P���o)D�X�2H��\t�!�ɣBێ���'D�h&.@�I��[%	�
Qb�0f!D��I7�O ����s�`Yh���>D��y�G�C�b��C��:6zљ��=D��ǂ����q壆//b���d�.D�����Ř_�b=PPlQl��5��'D�L[�	&@� O�	�j�q�H'D�P�����c��	�!߰!�B�#D��BV�ӑ4��8@H0I���	�� D��
�*<e����	(~8ع��#D��ia�U�O�	
�E�	�N ��7D�HQC�	�q'H��p��h��(J�L6D��y �Z��,m�q�	:_�4a�`N2D��!�hS�'f�РNH�fRqP��$D�����Ls��P�m�.v�a4E#D�� 2e��7]�$xJF�Y�qg �W"O�5#s+����ɶ"�=��-�"O�D�1���L�dԺ�G�A}�q�"O�L�=i1Vyc�)��^f� ��"O�0b��P�6�����jB��`�7O��=E��I�#
[<��d�iC�!p��M1�y�#
�ޡ��:`����ʒ��ķ<)
�)e��qB�R�{�X�����Ks�,�ȓKيQ)b-U�1|hv���2p�'��~� 
1s�]�A��m�� ���>K��;���%APi�W��D�JC�>�~PA󦉨Wl���,T6�$��$&-Hpk0��i�L���W'MND�ȓ*�r�(�sM��p���'n�O?�1H�i�!QR!�ER>z���'�p"�L���UO�dĬ���5|> ���@�=�vU*N�Ԝ��Nr��$�H�H��$ء�r	��O*D�4�`�%Cbl��C�4xy��3D��Ғb� ���:a!� є�ק%D�p�)mv]�3��WzT�i�/D���!Mx���ԟBk$M�Є-D��JDYH�p��pm�"VB�bŏ/D���Эb撱���ÄTR٘�).D�����4v2X����¯e��<��!D��+��L�K�T� %��0Ո=D����5<8 ��^��`C<D��
�ߠ7�>���6��m�7�>D�S��اW 	[���W�ˣ�*D��Y��]�h�'۶H�D�R�*D��HwE"o�Lpk���-�DB�l6D��a�m4C�$�"�]?��`�3J���G{����k��yQ��,y��EW�4l!��?j�]0b(�G�� 2���"I!�$R�e��}�����Fa����0Q����	�NCJBj\6���[�D�JfB�	-[�Ap!헥qY�@�dgV=�B䉼U�p�S��]�0ӑ�ѾI�C�I,�^�"���:&ОDjw�S=@��C��Ob�E86o�,�2i"�̏<>@ZC䉊 �Z�����Rv\1���L�#�.˓�0?9�n�c�P�QN�/-��I���e�<2)J�<:�e֪�L�yƆ@b�<�����Z kh,!gv̻��WC�<�Va�/f~.h���)I�:1����y�'��?��Se�^^�z�N�nj��p�8D�ty�K�Yh ̈�gפcL� t�!D�����	Y) ���<`���$�?D�d�g �|2R!3��b߬���
=��7�S�'PîHA�M̜`0MB�k֨_"�I�ēRx1+a�/X�L+DH�.y��]���I_8��b�ԤtsH9jG�"p�k�+7D��å�:.��%��N"FT�Dm5D�,�f�.-�ޠKG��&!��G�=D�,Z�=m�@%��-P�Je�4`'D�@@&��}�y��H�G��z��$D���Wm]-.�*��բ	 !cT�6D�qGD]�q3r��D_����P�3D�dzS�Z����+R�9Sb���0�|ldF��U�a�u�3��C��㟸���#�88(R+�6<���$m�HT#?��i!)��D`
U\B1�4�ƨg�!�DD}~(�+�l+<!Q�V�*�ax2%�O�c��� Lܹ%��P�"B���6D�� f�{Ā�(-g|��a��%M�r]R�"O�a���ﺑR������C"O
���)3"�ZdSNC�%�,�p"O�AW���E>���U=7�y�Q"O~0��AP���@Bm'% �Q��"ON��FGU�)ք8�'M?|V�JU�I6�HOV�-�<��b��l�!6��WqNI������b���s:T�5�Z�q���ȓ�����䞹<-.� @���Ih��n���[%GC_i}�Ǩ^�c>>��ȓ  B����ޅ���DoV�w$Յ�z�8�7�M>5�ő���oǬ9��d>�X0��u�Ax$���=TY��	B���Ynmk"�[?.��8&����!�D^�Lx�p��&?~T89�I!~i��LyR�|����2�� �"G2֘8ɂ��#�!�$W�t�Фѱ�!y�(\���9�!�_�d�>�[vS�.ͼx��GZe�!���">a�h��D��<�@�d���2��,,OH���@te*���Ώ37:\B�"O���Di��=�Y�'Ȝ*_$�H"O����ύxg����;pp���-����"|�'^ `� ��4<����e�&��*�'�
(�7��_舀��!'+�Q��/<OT��%ſi��i�A��A<"�4O���[�S���T͙H� ��g\5��Q��j��y��	�X��	9�⅗=C΁e��hO�O��,��.��{Vj���<�JT/@F�<!�en��iCK�V���"R*�,��&�)�矼�r�aj S�O�5�pAٴ�4D�����[�q��a�M�"�PŊ�1D�<��nǪ'or�њ:.�Zq�)}��)��E�<%#�;T�6�zb�� A�6m0��/\O��;�']��I�g��Snؐ7�Of��Dй+��0� ҹ�~�+���_.!�d�)���`�ܕ� �آ+ê%"�C㉭)NHLi���2�>� �u&���r�h'�`�W!�iȽ+�j�45@P
U�!D�<9�fʝ+��=�WI[�&��X�=�ȟ�?�|���1
|l�*ঙ1aL$!@z�<��ޥ^.�5P��ԫ�!+Ъu����?�5G@�{��(�nyJ!Il�<���]����W�ڴ}���C�g�<�7�?`E(M
��M�P�]�g	c�<�cl˜k5�@�"l]�6���J��\�'��x���?n�HK$�ܿb�5�d'�ybo: vv�81�+0��˵nC��y�g+4ŋ�0t�H`��yҤ�5�8�S�. %��%��^>�y���6����38�cE^%�y�#�/��e��OP> hn�)PjW��y��&{�NX��jZ�v�t�Y$f��y�ڜK��@6��	?���b���yR�ۺo���p�J�0��q �Е�y���2h���!��c�͹�( �yҿ�dl ����h��Y�^knC�r����!&KD��s�I�\�\C�	�jm���Ldq�m(t��J6C�I?4 � 0cM���'""C�;��}"�#Z5�<�:0�جE:C�IA)܈��Aţf?V���k�C��B䉊(�VX�^1B��{�($��B�I��AG�@
_x��Iҟoq�C䉅4�9���8�>�8qe3#��C�)� `���O�����`-�l)2"O,I�0>3:��/D�cP���"O@Q�wjĺk���Pr��9K�xy"O�EXbD�Fy���M3:�ְ �"O�d��dN�^�l����d����"O���w�V�)+J,��K���* �"O�XpQL�;/�VԹ�+�����S�"OX����N� xի��%I�9�y�F\̅��h�1T��p�H.�ydI&:1��T,C�\�e��$��y�C>]��z�* z�:���F��yrm��Kg��y�*��xv�"Eh�!�y��3_��!#��'H����h���yr�L�!lld�'G]�$�P�3�!O�y�ޡ@�|�0��P��Qct�O��y��G�f� |{2�B�C10�Rs�P��y�cE�AC�V(�RE�Q��3E�Y�ȓ'�����
�+	��0�@%�iۄi�ȓ'o,0*�BUn���2V*Ћ'[����(�T�R�/2Zb6`��>q���ȓ{0�� 	��YV�%eD�O�X�ȓ�T}��߶k�<��t�zI�ȓNr`#( Ar<Q�a��x�,�ȓGʀ��뎂_��(����0"���ȓ12:P�.�.ؚ%���Ӥ\�bD�ȓ2Ak��S2�ڕs0Ҟ�^d��~��M�`��]�,���N��c��T�ȓ ��Rtk�F��p�!��@V��Q��T�5IX.=4�k@��$�B(��X�42�n��Ec�S��� v2��I�����F	4J(f
юX� �ȓ���Í�eh����P,t����?@y�d��B*@��I��@�ȓ-#��Yca�+t�x�� �K��p��G������+���A�n�S�xQ�ȓ ���䈖��v�R�*�?R)� ��"G,u�� X����d�;6���ȓO=:��pe��Y�v��4i�F������y0)V��0BΙnL�I�ȓ,h��p�����$0�
ؘT$�ȓz�"� 'cR!�ܥQ Oz̀����8:�O�)\E�و�"ݸtV<�ȓxJ�����(`N�A�P�пU�T��ȓ��|��m7]�2lh6w�D`��@$Hwj�_a6��$,P�%R�Ćȓr͚03�_�zq�H���1�l<��Y�H92�o�-08ap$�X� �0��0�ƨ���5s	n�H"i�]��؇�$�ꕓ&6~6�#��
F@�ȓ.v��󴎃2�*ƣ�)h�цȓqax�� �_#uNH�B���\��z�>���c��x �#a�A:��ȓN�r�ٔ�#���𥥓�+sܤ���`u�F���p����4~V0��W��@S& v��5*r̂h[|\��*��Ba�$9��$�Bb�<L�%�ȓF̌�+U@� ����!��A����ȓ'k¸1��W/c�$qSGMG�!Q�؅ȓg��svn݆8�xq85*��mM�ȓ_S�{�g$R��y͊�mzd��Y�r@�C��7�r���V$=+��ȓx��Z�*^�(���A�V�U����ȓ$����.Ocf�X�"
z3��ȓ0a���^a�qP-O=O@�m��S�? ���7���/�F��q@Q�d�ͨu"Od�Z %�=�Cb�Ⱦ'9HL�3"O�̣�%�%�m�Q�F�0�`�"O��Ë[sޔ����0
�ts�"O�1[G�=f�
�2`�v�<D��"Oeyb�F�Z����G1?����D*ON`�2���;d��_#vxC
�'�A�K�3���ҥ�@`�A��'��u��C�*r-��#� �>BXY�'��� tD߾}��9��E�5�ް�	�'�z��7d**]�Po���R�i�'h�Dꞩk�R���	F�@� �'	إ����4m�������'���
�'�h�J��2+�����"7\�S
�'^�{QM �y4�V8q�I��'�̕ᒦ����3�L&614%k	�'021D�Z��1���b,-��'�Z̈5 �	�@�H��p�^�Z�'C�r/�$h�J��@�.j���'J.٠R/˪�y�e�\:4g.�t�<�6Ǔ�}�$@��A�{��lieLBz�<��EM�p��r��RŜ-���O�<�A%L�A��a� �-�=k���b�<��#]?��˧�� }dI����Y�<�Մ�n]p��W���kb�zf�`�<qU���$t#�䌧*N��Ȗ�_�<1��� �����X,nӎ�C��[�<A���=���Vf�>��b�� q�<�R9 ����D��	v��9�j�<ATh� e�8�ш('�dH��Ae�<����?*�n�s�d@	ph�����a�<IW(��y�Nא�ƅ�g�c�<��-�Qݜ� c��~0��!�LE^�<����J�LوC��� w�PR�<�$CC�6�8�&Vh�����K�<1�)�t����܂S�h�{�@�R�<�� D�_������z����qi�O�<)�%�����e`�9�n��C�C�<1e���z��$��O�6����gg�<�FĀ�UL��@	ޘ&l�af��b�<�p��X'��;4)_�����f�<q�-�9�4�3���J�����[�<	FH�`��� "J�/3m�h��
�Z�<�3/�M�dah�m[*�X��T�<-��EQPǁ�J�\�ɑ��F2�Y���tP`�N z3v�Uk��~l��6aʠjT, 3s՜p�⨌�;��(�ȓ(`�� ������
"h�p ���ȓC>
���ۢn��R��t*L�ȓ�J @�̅1�Z�:�"]3۸��ȓe��({A�Z;I��U�JŰX�.m�ȓF��!,(G�����X�PՇȓ1�R؂� �j9�� 1�U�u��$��I/Z��6�U�&Yp�nݞ#/Ό�ȓr^N�q2��jP�tiw��]����pc��L-SAp�Ö��l�.=�ȓq����u���<4�z@&̷}�Dч�%��A��G9*t]�R3T���ȓg��2���hB��ЩW,F3�t�ȓ�V��[�ح�qd*%"8C��2m�lH�"*C�>;�,q���%KXC��/)&�[୔#uHypmQ($�C�I +bY3�	�"�:,ʇ���w#�C�ɽ6��z�.��]|8�v�͋9m�C�)� &�j��
;��pd �|�|4B�"O�dȂf��>E����9L��9B"Of}�݊T�I�,�F�z8�"Oz����L�$��X�@�H�&�	�"O��AG_��q���K��t�3"O>ܱ�L]{RjaK��~� �"On���&Ev:���:k��"O�SA���	{b�q3!"Oza9���>c�L��W��i3�"O�1��ƙ3�.p�EEJ ?'A��"O�٢�`رs�)�vdX�#m:hJ�"O9��"��j?���,�TVL�P"O������[ܬ�p�	L����"OVꦣ &7���
� +_���"O0PᥦԸ�,�T)T
m��t"O��u.��J�y�e׫'���T"O��#ER�d��
��v�H�B"O�l(F�:Fu2�K	(�pl�E"Oh� F��jkT��rL\?;.AK�"OJѻCC<4�bѠ���2���7"O"�
�5~�6�N���b��]K!��X�mv`����	�/�(�q��V�*:!�dTo:8y� ����lm��R-!�L��j�ю�'{�yI���o!�9m�@����X�z�a �!򄚹}IBlc'&BDH(�g �e�!�DW�5�"2¢ �1n��H�J`c"O:u���
�&#�T�%#��p�"O�A;��K�WU�e{�V�fP���"OX �S�Y"�� ��D\��S�"O� �ɜ� �|#��ʟ2�\�;�"O&�7@��L�qPŚ�4����"O�d�c�Y��Fa�F��bY���"O��6��R�*���.EW�̑s"Ob`�)YH�hb�m�K~�xG"O������!j �����q�%"O���ExW�GɁ�m!�mЄ"OX%D�һF�����I�?@���h�"On�����T0U(�y����"O�13MAF�(��Q�	�X8�"O���G	C�j�D��,�
�p�;"O< `slL�a`�)YrA�$bp""O�%g�(g� xsD)O;ڠڒ"OD8.V%36���� �zI�q"Ol qwm\	a^�-�@#3~`�"O|��Pk\'���"��AF$`��'"OX�j�C�d�9WA�#h���"O^@���V����b�bN�XX��"O
E�gP�=�l�j!�"چ]�t"O��#����15Q;���_�Z@��"OXX����(ٚ	%Mϙ8�1"O<1�a S������D���&"O��D�xU��Z�mÇN�\�!�"O~���ĕ���!�zv�0"O��4�]}@l�UfW#و0"O�m���سO4f�T���F+jx�7"O:(녏!�Q �
�<lP"O��:�B=�8��pi�0r$5*V"O��ZqdS�@�>ᘇ��D)~c"On�jT&3����78����&"O��s�>*鶹ae�U}h:�"OTS5@�'�qb�d*"O����$�*(���[n�ZX�W"O��(��0٨H1SFA%c�4H�"O� 8�@�MY}|�	�/�D� ISt"O~�z�d!P"�P� $K�j���"O��8P������R$�@ƶ�B""O� �B��>�n�7�L�,����"OJ�Qj�<�P�) �r�X-2�"O���"&ĦW���/�1�`T*@"Oi�s�قpb�,�iHG� �9"ORQ��(G#wR݂ե݅#��PФ"O.��%�!�8z���@���5"O���"Ț-6�!�� ��Q�c"O|;T��!w� Qz3I���Xu��"O
i��M2a��%Q��e@"O��{C�\'U���@1���rjR@c5"O4	��G�B�$����,B�$#�"O@\PĂͬ~״�Q��I�:9N��"OЉ8umOhX�!m�'=�h�v"OΉx���3{�x�ӌ$)�}"O<�XeiR#o�ldS
�`����"O`	V�X�+�~�q ���v��v"O���5�U�%x|H+�Ο2@HI��"O8�y�̊��hq�F	CVp4�t"O0��7.�[_Lيr��:G��F"O���1�!�h-�#M�%Q9��"O�@�D��(% ��n�2t)� �"Obtre��EМ���7T�4z"O	G�KF����$M�q����"O��Q!W�^��ɵ�L�`�J���"O �"t dJ����X�,Y�"Oࡠ�@��u�͑Q�J-Ԧ0a�"O�= bϩW�T|��#��b舖"O�T�"ψ�s�(���X�a���J#"O��ا%�;[#Fh�cDX����"O�Mr6ʌ�5�<����
~j1�"O�\ۗV'R���q��B��S"O�H��.ߎ;'��B�[�$��=�t"On�cWO[r�*Ai�oȵc�$@�&"O��s�)�NuH�#��Z8[�vD�"O���0���5�\QD-є	>�)�"O�y��Х|2x�$lX��!sp"Onlh$Ι���3K��\�)*�"O��h���:�գGJ PWp���"Oz0�vfX=���ʢ�ˡ��,a"OhI��ʟ~������.�L"�"OL��ъ��6�p(C3�2K)B�;�"OH�i��N�XYk�N�|?H�b�"OlQB!��?++�9�C�L4O$�q[w"O|yC�)P�ؼ�`b��p
� X'"O��9�.�i��Qb�2�1��"O�9����@���է �TD��"O`���C�Bb���W�!a����%"Ox0V͐>_Vt�+0�ʩq �T �"OH� !EF&0&�C�!�G<,x�"O2|a�Ť��P�@&"��"O*�q�M��2���M=L��"Oș��,���hcR�ת7g��"O���FL<#�4+V��Zʂ"O��mR�Mz]�� �|�@s�4D���e��:Fɨ�32F�"k�V�S�
4D�43b�n�J]��%״x-����0D�$���F�Щ)�	 g�mJ�*D���F�����R/�YͲ!���6D��26��	9�1j��`��ؘt�r�<i��-a��="狳4��x�Éu�<2h0ba�$��j���ȅ�׭ o�<� ��Y`�͟Qx����c�X�"ORab��ݘg��M8Ƕ+e�8#�"O�P�BnH��#��$P`$*F"O�(��C�|��|l+S�q9*!�6"O4M�"g8cM,ѠA,ґaѦ�9"O��g�΍S���� �*f��T��"O"��OW;Z�Ε���S<d�"O"0�u��7�H���D�1����1"Ob,Q�GԾ�г.��X���1�"O�$�)�5P�Ƞ*��̂(KD��y	�1Q�nQ7D*M0�H�*1�y�����Ġ�h#na�P៩�yR^�;�"=$˙�F�ЅN�y��	
�|03)�*
`�JFOE1�y�#���٣��P��G��yb� `�:-�$R~�^\yE��y �:�>IQeN�u\���_)�y�Mf���#�#�5
�j�	ɰ�yb�%Wx�� ԢI;�8U����y�Hڿ6=.	e醦~�
EZ0�	�yr
P��x��΀2tb���d!
�y��
�azǌ�|
�X�!��y�!A�9�E��;y��t��@��y�L��(��T�4�͕n��ݹ ��yr@��L�&Q�X3^�	��k��y2(�$"Vpk�,�da:����y"�:(��,[���'ܙ�2hğ�yR��'��MQ��ʦgf�ke
���y�O8}��m����b���b�k4�yrl�2B�j��U��mŎ�����y�'��9�mڀ�Ɂf�ܼӑ�>�yR�?>Uҙ��"ġ(��(�$�y2�ĎX��u�!�Ѱ(�D��Ŋ�y�M�а0Q�N l@eQ�G��y���:��L�p��yq�]ఄ̅�ybc�=Q�L�j�Yar�L���y%;��L!�/�S����g%���y�A�sb�<ٖ�LѼM�R��y�m�Fk0s�lY@����s*$�y2��	w�d���6A��k�����yB��&��Ȃ��f���a��0�y�C�+v�r��^�]ј=˧�H�y��+dҲL:� Z} ����yOW4Mdfp�&oO�)�``d�W��y�V|��!h`�R�l�(q�D*^��y�GW�W�� 	��e��ha��y�A� �5i��B�W� 4j
�'9*�a�#ߚK�ЭI3$[�^��PJ
�'�ހ0Q- r&2i��׻&P��'O�-x@#E&b�J�a�9��a��'�tồI�?��8:P�0M���k
�'VB� �&��t:��ըFk8	*
�'�0�*� N�O��pbk�1CԲPH�'�94���tBa�qk_�(�2���'����L������){��
�'�HulQ�|����4)t�	
�'�$��Y���|�^�'�z���'� ��oª�ܽQ5�^�%<@��	�'��� �Z�/w��dkފgP |r	�'D�gC�,˨�c�g7B��'P֍AAc�<|\~8
ZOz<|��'��؅e\�&��Q#-΁D�H ��'�p�[��\�#Z�X�ͽp��'�ް���ԧ<�T!��4�d1*��� z���O�(v� š�-Е_ =; "Oz�� &����X�9Z�u
�"O����
�!gZ�$�-C=Pi� @"O�؛a�*QD����G�{���&"O.a+���+?�4�dj�$u�8�a!"Or�B�@�.P�z�[D
A$~���"O���/'V(��� g��0�"O:5�0܃Yf�P�� A>m���Y�"O��Q�B<ag�U�A�[�K��(H�"O�zE.~hT�b�?Gv��p"O.��g�]�1٘u�ڮ]x�7"O� �mp�a�N3yjra "O4�ɒg������bֵL<���u"O��w[dd`�! ��K*���"OƅB )��t��(0d�W�F��[�"O�����9;���pbS�
Ix�"O��1&�C#Ƶ���Q5|pc�"Ol�y��V��(��J=vj,	��"Oh��j��2����G١Ly�"O8�����1q��(�fgb��`"O�� 
ܞ��0�d
�O|�Փ�"O���Y�z��x�0%O&Ks�m�B"O\�xr�D�"-��x�\����Q "OD<��M@+S� #K��)؃"O���A�/W̄Ő����E�H���"O��w�U`*�%��
�y��W"O|��`��eX@�V��Fw�͚�"O ـ��U%R1��Av���~lݰ�"O��%��z�� ZÆj��@`�"O�l	r@ͼ2�� ɠlD
� `"Oht����?���C���OQ{�"O�H5�S�b���@��ޑ�5"Oȴr *[
X�(����ݮ2�$
�"O����8$�*��ۅc��UK�"O�}) ]�Ay����!�05b����"Oz	�5!A5N"is���T��!;f"Ols��-����n�?$��5�"O�u S (4��$P�l�	?�����"O�͊&�L�~C�r���I���@"O��`1�U^�>�����a���CW"OzY@�`ײX ���� �	�:�R"O��*����T�@z)D%9A"OHS�A���y��Y3�T��"O�Kak�%R&����0us�Т�"O(uShT���ҩ��*�ޠ�"O�q��j	�5�UQ��@���%H�"O2���*�6IP�K`��@$mkU"O�|���֟t\
1B�L^�Z
�Qcw"O
��&ֱ2?�	� 얦�+"Ot$�׉4	'�E�1��
��
�"O"��R:O`eq���5'�^���"O(�����#�|���q��@"�"O�m��,A�.!���U�t�@\�u"O��3B�|�d�&�25�"O�ܸ4K�$'@j�ҧ�3�<���'�0��l޸|�	���ԗuc��K�'�B@�S���m\6A�v���'^N�#�Mǚǆ�Y���$M��'�U�܊!��}S� �KD���'�0M3�J�7yf�y�-�D|`�
�'�2CG�(p���A3Gݘ@�
�'�L��4h(	'>��s�Y!H
���'
Ti�s8YH���[,~��M	�'� ��`�&�^�1����eRzm���� xu��d��ez����>S�ؼJ�"O�M����,B�t�Ģ��M�"�"OZlY����I�"��0^�
����"Of�!2D� X�UauJ�'��Aq"O6`F	'P�<1�JF�p��C"OL�{�D_,("�PQ��@�1�8t��"O�tٰ�]8cJ^e�VϺ�Py"O��Ə% ��XW�_�l�"O`[�lN�w���5)�M�`%�C"O��S �F��@˥mGe��$:"O2��ag��Y��G�y�4��a"O(!�杤b���W��x�L좵"O��y�@�?Q��C˞����&"O"�C��­o�X�`��E�b�"ON=�'D�5J��Q{��ʧ:64�"O�ub�愙/��Q ޙ�2"O�A�J��JhV��P$	P"ґ"OX��@LWK���d֐`,�b"O2Q����铀��O�9)"O�99���;R�>�:��ڳG"L{�"OT]�e$ Rf4�i��*��""O��AB���z4�BD�>or���"O������SE�#�̆�n�"O���r��	���Ӈ��$�T)�"O�у̐1Mh�����,h��݊d"O� ���F�vpt�vEK)NV$�Af"O��y&NU(J"ND�f�Z�`B����"Ovq\
T�|�Á�C�|b�"O�<�n�*/� � ̓$�V��u"OF��`g�6,'�큳M�k���2"OR�!O�-{�!��:}B0�0"Of�iSAd��?jr�=` "Opdˡ�ނAc�s6��79Yvq+`"O `GaSC��%++ǆ;,p��"O�S� E�j��և�\'n��c"O8��r�'*�.�S��, BVM3�"OfQYa�pJ���E��#$|�Q"O�����w�xXc�:ap�ҥ�6D��4����BTo�雡�?D��+�΂5X�<U��,Bn��=D���[�eRm!��-`LI�G:D���r��2z��u��^V=I!�;D��w ���X�9b��s�XC��6D� �b�]�T#4�!q��8D�P��/��လ��kճ!���! 2D�t pM�J���G�0p�>T�v*/D��'N.�tq�G��t���-D��Zvҁ$r�q�4cH�^�eb��'D���F@�����qh+V<�{`(D�lzC㊽fQJ�r�φ�.nͩ"D��b�k�0i0rc�', Hj+D��2�F�%ȼ����j��H�q�,D���]��e���<LK�p�%D�<�vM %s�`DB��6]E8��ԥ=D�T�g
�(Q>��T��> ꠂU7D�$��K��n� 甆H��U�N8D�8�4��Z��q&k++�-��L)D�8!V -L����K5➭�t+D�,�CO@I0��Z��gQ2�7�;D�P�M�i�Y�&W��Juhh?D��k�ʀ1Gd��G׃tF8!�gh0D�,j�陁�]ˣ��3l��yC �:D�tC�
f6��Xd�ֺ^C���r.9D�,��KT#3T�i��C��MXP�q&7D�� "�a�&�%m�U��K�4!�K�"O(!�Q�(�E�4���2VQB"OV�3�� �������٦�6��e"O`Ɂ�L�],�Ƞo�,m��IQ"OP�b�@�V�\ �c���_�*�"O�%�¡^(��\x���y֔K�"O��2�Cޒ�4�:�J	�p�4-"T"O�9;ׂհj��L��i�#I���U"O���O�^y�$Ú/cB��@d"O��)�a	�Ss���"�5k/vE��"O�]c�e�8/�4�p�G#F��a"O� h�d�0#���! �1J!Z"Of�JQ��+c
ȡ�L�i�����"O �#�/)-�p��?T�����"O&����Q@9�ND�:S�苒"O��S�P/t��x2�׬ZD�ɀ�"O�����@59���!�A�6[T�l*�"Op�)"hJ��@��Ӗ؂4"O���d�Z^M�m�V��S"OzAkd��_��U�
�����"O @J�D�L$�4B�"� X���8s"OP�Iጌ���	�ToE�xh`R"O�!3�閣ܢe�s�ܷ#�Za�"OT�C�8pX["]�b	G"O����o��3��g�ȇa�Lz�"OD�`��m�>��ْ`z���0"O�Qh��B%]�D� �)�p����"O(���n�2K4��Pi�|߲4@C"O\D����!~��EnI�`�޸q�"O&�8��E�u��x���

�R�"O�*Pm�&bN!�X�n��V"O����@��D�hx��%�u����'"O ����Ľa�d`���A�l���c!D�:#'L��u��Q��Fe��L;D���ѣ
)�E��n�8zb訋3�<D���P�T(�.)zt�ʒ5��s��>D�,�v��6s�4�R�����|�#�<D���BV	���1���*���+u�<D�Ի �'b��m(6���HFYD�C䉻By2��@+(�� �g�.7��C�	�*&P��J!P�,{q���Si�C�W����CM#�t�k�fݱ�B䉡F�*�!ᤂ[���kݞ#*�B�I�,mf$!"i��rv��`�EL�B�I��,k�l#r&�A��כH��B�	�>\F�KF��?�z��4��MR�C�$dE�	F�k�p�rGV�O��C�I�.��1b��/�h���~Z�C�Ir<�!�CH'�-����Q�NC�I����+���X%c'D�� C�I�b�����X�[*%��� �&��B�I�|.�D�`���ZwȭccB]q�C��.��Kd�� �����(�;fC䉳hEj� ��%��!	�I�U1\C��E�(5NϮ4$8��&P/DC�	"������\���U����n�0C��|�Ě�
�\j��4���q1C�I:V��A�--��� 8�*C�I%92� �O�S����T�W�C�	)*��[&d����x���B�I�$�Z��f��:u�U�S�I�+��C�I���鐤I�r��5+��e��B�ɮg��Z�Nt:5�&F_�evB䉭*�v� �i ok.a�+1M�PB�)� ,8#Ŭ]8�F۷ud�`B0"O����a9C{��i.6@�!"O�!Aq��f�l�30�^^)X�B�"ON���cG�*�����*��%�1iG"O��{@nJ�nLM�Ѫ��#2�V"Ob�����P%f!H��߆|l(�B"O���ڦR�TS���C�( e"O&D��ܠ^���a&�	��Dh*�"O�"�g�
Kd-P��
�h�е"O6d�vi.�x|Q�T�D����"O@��5n��h![���,I�\��"O��H�,�v������"f�t��U"O�u�'�G�7=2y��Z����"O~И*�Ud��¶"�,(p5xr"O(��RNH� ��|��S�:�bd{V"OްH��1X��,�o۴�Xի�"OH��Pf��[mF`��K	&O'
�:r"O֥�
�<wS��r�aٱy{j��A"OX�2+@&W�P��r.J�N�x2"O�ˢ�p����Ďz�AKv"O̅ka�\6�0PE�Ze(9��"O���5��z���p�ᆡ<���ps"O�|��A[�(D`���Q� ���R"OV�Ԯ�4ց! �*p)��"O�Q[a��/��#��}f�5�"O�Y���AR���+�mNn)3�"OP�9��CT<5qp;*$��ڂ"O��W�ԁU��Pƨ��q�ѸE"O4y��/�"<$�h�l
�K^I��"OdL��j�) ��3!G�V{�h;G"O��r��j���t�Z ����"O^̊�X�,�U#�.CTU�S�"O$��q�@�z,�`�G�U��$�y�"Oz�����>"���v�ЕN�x��"ON����ՐA_F�"f�32��"O�#��רLF����⌸,�l*v"O��Q˓++"��3�&�(B,��"O|I����(~}�5�Ё ���P"O��0Tl�x�XeСd�.^�x\�1"O��H�x}굈0�g|Ԑ�"OF����������G4�@ '"O�}I.�<_����Fb5s!�D��"O`�����
�Bqgb�"rZ�Rf"O�d ���Ҭb6"͖B���0p"O�����6jA�A���'6B�Y�'�H�@�&
��9���]�)x���'�0زa(X�Ml�D�W�_.&���@�'ĸ�x�e�=���O�P8,��'f�=��Q#�2�ɐ��[n�H�'�jsBD܂Q|�؄�	*�	�'@P�	��H�N�uK\4S��+�'"�%HfB���35(^�Mi���'���I�
\!�$�*��L�F��'� �A0"ǄH��s�#PE����'`��Z6wA��G�G�)�	�'͆h4�ڸ� �V,��$�c	�'�:��F!�+g����U&�]�T	�'�A�c#K:P��9#$�οc*l���'E*<����9c�;Á�)�Ht�	�'��uL`>>EY���!{���H	�'��S�m��6�lq�u¦�1	�'�KB.��h������k!��+	�'S����)֏K��P7+�[�����'Ͼ�+�f*�ub�*�&QԀ�	��� ��T�D�;�`�Ƣ��7i\M� "O8�G��Ȩ �B-`^~�"O����$�<i�ļ��ߊJ�6"O��kDJۙ���!D�#+*�j�"O���0c�44�V�����&�``�"O�X[���)���D#s�j�k�"O�}���̋v��r+�>-�"4��"O���R&�h�`%�����3N�Kg"O�	�&��
�8�gX�u��0"O��8���^�rܛ��S��A�"O�]fÿp=`�s�]7(�Iie"Ot!�W��Fdad�M�EةK�"O� ��"'�b���MS�B��v"O���`Y\�B��h��l�"O
�z��ΊA��]�N��h���"O���Tt��������2�����"O|uCGP�}��(3"O�iOP|�%"O|%�
�2r�����J1!`l��"OR��e��)����fS���"O>�+�$K+d�H��ؔvwƕsw�4D�Db�\�uc��˰��!����0D��Еh��i���`��a�^<��&#D��*��9(��=��G�
w�0,u#D�<�6�=M�21cM��t�88�i<D��8t_"4������<墉rU%<D�(�gF��:����fφ${(�x�/:D�ؒG�6g������&�����8D��P�ŝ�>�Ը��H�s%����o5D���Gm�I��E�@�&(㐥���5D�<9�k��:�y�%�	zA�	4D��K0h[�h>��q�F�*�$���d5D���`T�sYFD�����:��0�5D���A�OIީ��N4,�21� �8D�ph�ɘ��$���_n杲�8D�4T��#�Z̓�g�Q?�U��*#D��s���:ai���f��?�|���+D���پ]��yDDѭv4d1`7D�P�V�*;���&�8̡'�7D���@�
w�t�����t$��!�
6D�,9� 2����P�F1`���"�J.D�8���#{+��s���h��KB% D�D��쎺 )4�P�&D
Ħ�X D�Ps$�@�[���7����>�O��N���{'���9�~���e
�2�~U�ȓ�ܨ��@��v�nH8�Ł�/`�4��Z渭S�|$dZ ��	4���:]h����^��k���Q�NP�ȓx�x�$N\��4�u��
O�j���f�N�����TcV�
�&���1�\Ui�$Xg�!�U��k����3���<I�`�r���=~���I�PI�aª*ި��`F�bzM��s��5�҇I��|��\2gD�0��@��2�CʭE༙
PA���R���-A"�Jv���AH$J���0|�na�ȓO�&@�r�ʉI&�l�p��b�|���<O���%+G�\��\��F
x�^���Yž]bP�X3�!�$Y���!$D��ᇖX$v�A6�� $@��$o6D�<����L�6�7�P�V�Ԅ�� 0D��.�=b�$���(����*"D�x���_-��ɬ�D!y%�*D��@woC*hp����ƌU��MB�)D�`�ɾa�u�2
F�X:8SEI)D�� N	�`�Hc4%I��Q���X�"O��yd��YYR��2+L�"�36"OƩ:T`��@�%R	�/R�Hu��"Ov�j!Z�M�(�0���dcR"Ox�!��L��Y��ʕ�`R,a�"Op���/d��e����j+~Q0"O(V�X�Θ��O�~@6@h�"O���!�E�0��!��X5F	�1"O�(�#� 5�	,��*�(L�,�!�$٤C\T؂K*?#��B�Hߏ!�Ĺx>1C�a��,�`D�(t!�D
)��q�b� E�>�i'`��!�$��W���@��K�6����,y�!�&R\�H
����A�b)G!�����<016�!)������g�!�F
r)���ӉG1`����Ԡ��D�!��]#,ł����\2]g��q���!���[�����0Wh8�4��r{!�^#S6�Y���s�	��*q!���X�dC��Q"���� 	�bT!��$�2��N�Мz�_�	!�$�)^��ga�X,���/�1�!�	F�ܩ��/�L
�EaP!�䇴A�t�y���q�@�K�G�!�dH�ޡx��P�se��X�>�!�D`F�`D�E� �4)qSKS�%�!�$�<4���GKE8W��i����!�U4`ZqS��A30�<���Z�u!�dܫ,��p#f:[
|��)Z!�XLJz�F��] "��*.�!�dշcZ�ϝ��@� A�B!�D�	nΠ�#rg�MpF���
W!�$�vD�JӨw�b���f[+n8!�d�vx�!@���ÐV%R��!�䐞;$��$�|���d
�:}!��!-��z���0,�P�9�ָk!�̪W���%��H%`{v �Y�!�$ќ�.�Y䒯-;r�{@�E�$�!�d�h���B+;>�݀ ��C�!�$N�Ajh��Č�5�,`��4G�!�ڻ3���5⛽`�>�""c )"�!�d��ԉ�օ�]��i�w�A/L�!��R��Є ȣY��l����0�!�D2-$qq��@�⸫��(6~!��	Ov=��"�"'}���!N&l!�䊕5� eID��5cf�P��=X!�� ��� +Z8Ic��j0��!L!���/*%�5��(\l�V�j8!�DʟQ��u�G�=A<d��j݉�!�$GoZ�̀���I"�@�-�!��eTn�p�hI�/ԝiwȜ{�!��@и���K3^D�贊
E�!��/M�`����J.M�)V�Ox!��9`�"d0b�8lh���F�!���h���[�Ү��CZL!�C"o�M��T�WZp���m��%I!�	ulb@Jwf�93���"�E�zT!�Dǋi�xX0�%V�a���x�j�k�!�d75�^Q&aE[�>�#fʘ�c�!�U1\�DD��C6:�(��T5J�!�$[+�����D��n'�yP��S�!�P�&� �gA�A 𡉌y�!�ۛ"5��Mߗ)'> ����[�!�  �0ֆ�$G *\ z�!�� ^RRf@3i��{�,hF���"O�aU/؍$��h�Ň�
I�S�"O����V�%}x��gd"�q��"O8q
�M�M���X2FA� ��"OD#���i紘:c�L>}�	9s"O��a� ��!�@L�]����"O�Dȑ��j�ZA͇$��p4"O̔!�i�q����F�A�t}��"OF�r�^�
�$�	W��#W���"O^����7r��V$�=,���� "O�l��"W+_��}ҁ�j;H�s"O�`GԿs�@U�7�Q�; 䝢W"OĄ��䇥I2��];Z�r7"O����!�%��@�#+�2T7*e��"O��+��Ɠ94���	ē3tQk�"O�z�ѳ\y��Ѱ�r���7�c�<�f� ���Q��HЩ6<�g"�s�<Y�DY.5\��sG�t��1��Mp�<)C�[�j)�4��P K��EJ��Q�<����(�F���no���IK�<��O;�(=h��N�Ρ� �bC�I����s�
*-
0�{UO3��C�	�G�۰��!TB�G��'[�C��B%�y���51f��wAJ2�B�	�0����@��5[c.N�FuC�I�>�8X��Z:<a��sj�%�B��9Fi�a!��E��H��D�Y�B�	�L��E�ӏD�EY���!"���B�>⬉z0&(x�4a1«QNDDC��?Ԍ�ƍ`���(
o�>C䉻k�t��0HP�+�G	
�<C�I�vt�[�g�kpsBf�&��C䉦U� p+]�F�:T��s�C�r: @��'X�71l0�6���C�?|Br5�G��;S�4\���U��0B䉥��I���;P�	j�F�"L�B䉦�,���^.kUܝ!���@B�I�,���`!�%g���2A�q��C�I���QK�)�6F�jgd�&w{�C�	]� �B0� �^U�g@'+0�C�I,G�t��dIT<m�"dn�>Z�tC�I�b�с��) % 
��N�rC�	��Y+��ݰ[��8��EK�T`C�I�Y�̰)��EBǖ����.B�C�I�4�<IӴ"1D��H�N�,i�C�	;Lo���'�;(/vaK��P�B��8^%��b�bڊ-�Tu���S�H �B�	�L�֝�2�Pi�AJ�l-��pBH��c׉X㬭��זME!�$�&VGTp����Du04+RjZ�y%!�$ӿ�RM�UB�0T����֗!�Ԋ{,�@�c*�.<�4��h�|�!�D��=�9[��ɮ4�֞'�!�$��)U�Er����*�ڤţ�&E�!�Ƭe��5�b�8s|�KA�޷P�!��PO4Vx!�HtT���W	Yt!�d�,\i*�@M�G�����Þp�!��"+�4DÒkK rH���ǋ�^�!�D h��ٷd�i���@K�Z�!�D7d�-BFEK)dŋp)X!�Q�r��Qa�20;�x����Z�!�䂀Z��Y�'A!}�p!ah�V�!�$
U�Խ��h��Ce�\`S(Z�8�!��<'���䒆TV��V)��1a!�� ��q���y}�Ċ���#}Dz�"OI8�*��{��C��
h���T"OJ����]3aj^�k7$�2\SHB"O-��fU<�%0�֣j�H`�"OXY6-S
[�D3�n�	"���r"OX`#�,ɱl���:��Zgx,���"O�9��վi*p����tf|y��"OF�8U��3E��	�ՠS7�Ds6"O��YQ�=ix��T�Ә����"O�H��ǉ(e��Ƀ}{Zl+ѣ�Y�<	�mY>u>x��J�$} ����\S�<! �ějѤ�@$�����oD�y��8eE�0fD�7�@Hg����y�Ӎ��ݱ��ɀ,�"��G��yB�:���@g�KA��C�(�yR`��g��phE�M�H5������y�/X�L�>u;5���K\�i���%�y���Z�B7蜮. $�'N�yIMg�:��R��)9�a�v����yb`�b�V�*B
�%<�m��鏹�yҮ��̞�+v*g�2CՇ��y2 ��&,��Ā��8��g�ۥ�y��	%�vQ1g�|nEP�	��y��E��tj�Ǉ Z�v-1󁟨�yBh�"q߾�xC��YM�p�iG�yR�B�0���+_Ef�i�f�?�y"JӜRx�����H��L�V@��y�LΌv���q�M�F�JL�����y���b.���aR��<i��@�yB(�	�����*���7	U>�y�i�/0��g��[�K��y�OA"7�.�0��A�WZ I��@��y�F,Z�Դ�c,Ryt�g�
)�y2׳
kR���6�∁�<��ȓI� x4�߹.���#��ĺh�ȓd�
�Ir`�i��MK�L����d veK3���A�D�1�2-��uu��b��D騡�W�]'d��E���1 1��^<t����$[��|�ȓi���Ŋޖy�0h���khl��f�������_~����B�e��(��h*Rj*'vz��B��s˂��ȓ)B�s� ׹6j1�Ң��BO�%��F{��nEj���6_hip� ϼ�y�f?Yf؈���5f�%ꁨ�y�:OgP�)� �{Z�0��+�yr �����F�9@`����B��yRE� ���+"���m^�9
��yrb ��r�"(v}2uO�$�y�L�jIJ���
����"R�Y	�yBA+Ax�r��uqtсn�
�yr����8�%^�p���r���;�y�o���ċ��
�a|�I;1C��yRH؇k̶@���\8�ȣ��^�y"���#�,��j�'N-3��Ѹ�y�^��2yB��>y$pj݌Y�!�[s�"t���E�$��kV.5�!�d�� �W�ӸO}^���  ?a�!�dA A58p����mj�P���J�!�;Gޮi+W��'`x5�ՎG�!�$g�r( 4�'t)��b�90!�I�j�}bK�'y}A�*أ�!�]�w�0)��B%S�"�3)I�>�!�dV�A�d�
��V )�8h	��Y/�Py
� �ȳ� �=�`F�Z?1J�)'"O�(�5���-2 #�H1��A�"O\�D��U�ĺQ��W+ 5q�"Od1�  �,�a��	՜& �hs�"Oح��,L(p)ĉ�Ԇȓ%�q�"OK�.% n쓳��xb�9�G��y����q!�ɶk'^|y�흟�y�%Ȧ=X�B@AS+dG qڴ��y"�Yf�fȹ$Ga�x�H
��y"L��k����� ٴZz�h*�e��y�ڬ)�4{�χ�=a�x�#���yr��>\0� �Ҍ@�x�  �A��yr��>��T[C��0f����lJ��y Us^�@b�ȪTU�\
�cT�y"�T��l� �j�=!����(ع�ybH7~\�͈9�.��V+���y�-�=+̾P�%B*cd1������y� *�P��!M9Uw�=a�����yB)]�w�d�rq�
�;�V4C�'��y���1*.e3 �}.�iJC"Y,�yR/�0,�<��퓿F��T����yR�C�*�d\�s�G�V��UX/�y�l�d�8���D�|�0���Y	�ORD���(��<{��ѦG�4A�H�<]��"O���`�oP��6+��@%�TB@�O�=E�D���V	;��T3B�Dn����'2�z��Q��Ҧ��8����ݱ��'�9�削%Pb}!��ٰX�4����k�B�I�1�­bS݁b���ï��â�
�'��~��B�-̼�5L@��N8�0>�޴�b�D��=(���
]RQ�cB*!��;$	�" �k�y����,+�O�U��J$����)��m�g'֡j�X=Yd�+uy�=E��'�1
�ᚷ`�x�l��w���k�/�S�$�g�h���\*F�As	��*���Qv�ƐY���$C\��u(���0ŀfm�����=�!���9���,	�{��ƅ��E#a|�|��HR�S'x����G�<QGG(d�"�3��5n�P`un@�<I�jX4J���*�� 2᫦ky�<���V�2x�ȓ-�=Z�#�CF`�<1%��j���V���4���Df�<A0&j��u�T��I��:6�][�<��m�+^��K��Պ��B��,���	2� �pRcJ�T��!�K �*��B��$���,ͶM�M���&-jB䉺Cw"A�J�*;`�㎀�(RC�	/-!�E�t
] >�3H_8NO����w8�=r�KA�U����nH!���{�l��A��Hɡ�,��z�!�䛴u⪸"�c��7P���f�ܖ$!���� ]|��f��<+��ҁ�C8!�Ė�4!^��I5%'pP{�BJ<!�Dŝ8Ih�� �O��C���Y�'��|R��
:buÒ�؎��g��+�MK�{B�O����(u��a���v�2����ۦP����;D�($`ׅ}���f��֩B֥.D�tӇő�a� a��=Z)p�:�+,Oh�<y ���	���$O`�Z7m�݂ͦr�Yc�S��M�F ��uݾ%�TN�f��!�c��N�<��n.?DlX�/�^����r�<�&ID�W�>4�s�C�F_
�f�D���'��O|���0O�f�E�%'�ȁ�"O"��Q/�q�1��]˺\�"O� ܥ����zJ*=x�O�r�� s����<�����B��R��7w��UqA(��Q�!��Faz�92�.�*�F�yU���O�p�O>E��4"��0�5�/K�U��"25!����T%!��+w��(5O��<E�=���$"�D]"$��-���=&f��Sn��y�!��J�v�s��F*h�� W�߽5��ON����i��#T �<c �}I%aW�`���ϓ�H��	�#CDl�:�0��g�Z��i��$_�0�����e�#/A�!���rI� �ÀE�i ��#V�	y!�B#<K��cr`��3�>�t�1:!��@)s�5 1�g�4|3T�H
!��Ѧ^�����Kj��V/ɪ�!�D����ـ���o�pK�M�g��|R��(�s��
	�e��T($���ֆ�93T���j����P-��'�� )Ŋ.��nZ��x�tC�58���j�i��E��HK�-L��Iv��h񏇇y�f1r"͑&?�����C/���r��7�=�9m�z��3(B� 2Ys�EԄ[�B��z8}���A���A0�+�ݰ�'�d��|�O,1�FB.p�A���$g�I�$Ǻ�yB� U&.�kd�	?]���1�OP}R�'W����U�v��t��FR��X�`�{_��&��I|��j�>B�y���U��I�<I��I!t��	��Aʲ|*
��-Yl�(F{r�CNg�h!��S=o�����Ə5�x���S$�Y��L�C��e����P�V���;ʓ*���i�CZ�kW���s �6����I���C�� Kt�����e�d���ȓf���٢�D�n�
��V���x��Y�JT�R*ԇ}�٨Ι�+�@���t��s�2�R�`��  
	�=IO����􄇼Tq@��,|*�ݙx�\��d�>G��'�B�1��$m����l���<1�����<��lM�'��uP�p���3_h*����'��'9��0H����˻�T�dݾk��&�)��)q�P���T�7C�^F�l�&.D�(�"%עT���Z�!�X�iC�<�	���5Y���O=D��T&��FR��'-�7��C�'6��X�]-�[b.A$r�a[ڴ�PxB�2D����uPWL3�(O0�$�h���������(�oX>v*X����$g��?�V�d�~2h�-�$�#@�T�ڈk�c�'2��$�<�'�>U��M��Z��Xc$ԟxFe���Mi?a��-�SG��&�;?�!�d 7��̘���1Pm�B�	)�D+C*�2)�剢K%rZ<��A?�O�q&?��~rOQ�1������ sYA,��yb(����4` ,_	q��4H�,ɻ�MK�?�Fx")I����[�]�z �0r��H+�Ox�=�O�8�f	�(n���$�R�	6 ��O<��)�S�K� �U��,|�b�o%,/�B�7q�aĆE�"��C�	T:+1�b���kW�=�wmæV����œk`�=�=a�β���Ot����f�j���ICZ%�C�'lOn�S��-����d�çJO�@���Zզ���4�����$hb��)
`�3�+~�b�����D��h�vtlsⓂ~iѷ��*[��1z�e��Vn�<y
�R�BhfCٍrv����)��]F؜�>�������'�����Gm��pJom(<�0,C�o||d�Ğ�|0���G�F��O�6�~�}Y�T�����ul�w����yB�G�F선�N�Jx�W�ފ�y�j�x_�Af�� iy7�S!�y
� �Ԡ���|;�,�g�s�&�1�"O�Zӄ�=+��YfG �w�:8��"O�����|<�$S�K_�R���"O�Tp�+?-x��$�ԁ,����V"O��-.:bd��o�D����p"Or[a-��p�(������ q���"O�T���[�4V��0G��&�K"OrŪT��6Z��󄦎;��9k�"O0�Xg�D'n�P̠�C�@�ؐ!�"O��&���=zg��-���D"Oyp�=���c!�5�&U9`"O̤2�L�k�n]2�͡�LI�"O�9i�H �"i�!P�T��y)c"OԀ�d�Tq4�����F�z�P"O�k&�!��]p]I���)gT�<yd��9`<Tp1�B�Vp-�g@�d�<�F睘]���@)�f)B��тJd�<q�f�c�r����F��Eq�z�<ACD�|�!�S�Á!pB� �M�<A�(�]�@sfO��y z i�/�@�<��%�ވ�d+�}��0��&FT�<q�n��l��+�B� d���bf�Xe�<�0�E4�e�w����� tωb�<� ��NF���(�)�&M��_�<�v/ɔB���C	?D4�9���W�<A���yw�r� �7Ɓ�t*�L�<I$AY�=�h2��Ü$
�\
�GN�<�@倉H}��fL�a z�Q�oA�<!Q#U�m��@���#�|�V+}�<#�&��1 ���kX�M�#�}�<y�.��L�I�@�+
��ł�u�<�ͤ>�jE��>er�����p�<af����ųEl\�t
�1)�Xk�<�j��C�M�ci�=�6*�L�<	���0nw�x����+�l]�wJ�C�<��L�OY����D��ce��`nB�<ɂjǁY�t@X�"G����ag"�x�<���cn��d��^Q�9�*�t�<�Ы2�JK��G�w�J�)�f�o�<Q�K�{ĕ�Q�,K��g�h�<��LM�d9  �.d���VĖn�<�d	�	E�b�˦�Զ XZ��b�<�%0U���BW�p�F�[S��g�<Y%�ץ4H�z2���&yC���I�<��]�h��-�J�����%*E�<���9�E���>yU^���PC�<��`X�Kt|	��A�#�2���|�<�"��
�*��!!\�i)���c�<)��G8����!���@<�p��ǘh�<��   �Fh�&�f���@�Ba�<�A�Y�r<�xr�ʛ�m貅�fFu�<������d�"dk� L4E� j�<)5e�<\��|B�HW E_���h�<q׬�s=4�8@VB|��ȗRa�<���-!����h�>~�l 8��v�<)r�d�ĵ��Ӻu~��¢Lv�<	�GҹC�>��'�:�΀���w�<��n�7L5#ĉ��X��t�WZ�<�tE�7>��Q�D��6A-��*�e�A�<�d.ɞc���@4o�P�'�Q�<iÅ�'��|�'�L��>�)C�{�<9��B��yV��9�j�yv�<I���6}R�#�?t� ZW�t�<q�,k�.P��
.f bg��n�<� �e���1g����$�H�yz���"O٨�gN-j��{�D�)[0��"O��FN\��E�_h�}x���C�<�#�/��LQԂG ��h�t�\t�<iu��yh��VE���@�a��r�<������$��,�c��u���z�<�	͌s2�pcP%YG9�wz�<�����'�<�I�(���g�_k�<�D7��R,�&��uC�A\\�<aT��8n�y�Ǐw�> �F �p�<Q� �/���S/�a�H[X_�!���o�^}j��%x9�ȱ&�1g�!򤝉nr�l��G�\(r�F]!�$`�f��T#��$���I�j!��#��K�@��z����ō�#	!�h:y� ��C��p�%]J!�ā�/2��T�4��c	�;3!�Ď�:W����
�no������/o<!�d�8cP�h���v[u�����!��ʠ=iI�)�*W� 8&��%9_!�DK�J��Q�ŋC�>����kCc!�䝹S�f�K�-W4��g��8[R!�:�p���??�z����_0Z�!�d��v*�2� G3$�%�E5e!�$�<��]�L#@	�GD ;J!�>-��C\�����7]<�8�G"OPɉElH�VL^-kV��pI�`h@"O��R! k��Y��*|�l�ɢ"O��y�O�x[@��SDX$}>�J�"O�%�� @�8.乵c��Z�6x4"OtY�\��l{@� 3����"O�x�� ��c<~Xʀ�B'l.���"Oؤ��H�.dJ	àU�G�L���"OehT�SRZ-� J)M��0��"OP%�b��5o����>_�䫕"O
�J�a��&��19#ɜ`�F��R"O��	��3Z&֭V.��˂"O���*�|��a�
����x*�"O���OG)?�D���� �m�A"O>���Q;n�L�� �\x�1�T"O�ȊJ�Rq�`-ym��`�"OTA��`ܹ(��Ёp��OD�Q�"O$��Z?j
pQO�T����"O�9�e���X.޽�5m~���"O���%ϕ(/��B�R4Y�v"O����ҌA���B0���B-�4B�!�N=B�u�u��4���� a�=,�!�䟫$Ƽ���MUr�K��-Ne!�D�+0[E�6���{\�0h��W!�d͔d�*�N��
R���'1#S!���/F�j� Q��.u�
T�a��/6��Fx����#ЇR��|�*��ǁ\�+��Ȅ�I:%���C��#Q���#)=v(B�	�Mh\Pa3���f<�Q#N�
�.C䉡KX(��+.��=G ˜mzC�V�V@�WM�',�z���7�PB��:&K��
��R��6%S&B�I�Q���;���'٠,�%K
�$B�	�}���h��%�xho��{;����bD�d��%kN�� 
C^��4���U�F�;>��� D�eptŅ�WO��k���4ݬ�QpE����ȓ3Bp]h7�S���Y��mQ�@�p,��Z��$���ԅ/[�-�@'S��X��S�? ��!��./9��H�!S�&� @!"O�!�D�$Ct����$�򱱇"O�9��%7��Q����;E�Rę"O�@3���Z��aT�����٨�"O��'��5)ytD���A&A�@���"O��:��Z�Ce(1���U�|����b"O� ��a������Y=�J�0�"O����@�e�~D�"��5yĦ�qc"O�T���{ֲM�Ub�����C"O`�9�闞}�6�ñ'$#�����"OvE*���1G0X#�X�^��"O�Er�U��0��W���k�"O�D�p�%`��2�zXK�"O�P�N�d���JV�LrP#�"O�p�7�3p-FP�W)˗#[���"O@���`@�OH�$a)�Fr�%�"O���ezi��	�(�K�����"O���Ϙ��T��g�*x2�"OT,���!S� y+�@ΐO�B"Ob pvJX0K�VU�$��8d���:�"O�Mk�E��� �$nI�e��u2!"O�r�/��|�*�f^	Y#�陦"O��� 쇡[�b�F�2�Șg"O�pXW
|�M1_:��	�@"O6ݡ�U8� ���5a���w"O��æ���e��L�|���4"OY����B Q�֣�=y$��"Ob�0�(�'=���8W��`o�m�|��)�j!��kP�3�~(����QCB䉹2��{�ʱR� ��ce͊8|�C�	a��p��Y�(�x��&�=}�C� w:�"6M[�K�� �4J��C�I�Ljm�eß3����h_�#�B�I9������P�Hy��c��\�MM�B䉙:vư���P�-J���XL)>B�I�q�����J 
D-R`b���B�(-v<j.��Vo؁P�ױ��B�I�^���0"��|kv9pŊ�1�C䉟&�,�RT���"rO���0C�	�/��v��6���3 �ʰ�C�I9m�x��� =*��;��U�za�B��;7c��Ӏ�P�!�� �E΀�]ܦC��2A�x�h��<v` �F���FC�I,0p�B��(h��2g�� Ct�B�� V�Ή�gE�	O�T"��!��*R�������D���\�!�$��f�"7�N+X�i���ʣ(�!���f�n0ucZS2�!3���!�%4�R��D�B���!r�P�_��'�ў�>s�BF'_�(41�m�.n�yv�7D�T��µ �n�*�+ɲ}�!0D���ab�v�jF�ũh�R܂�N#D��TMC�1��ԩ�������3D���C$' ��4���+c��AY �0D�d	����8]*A.�#~�E�1�/D�D4�,5y	{��
#�x5!#D��H�C���/���H�  D��%�L3RHڰHK� �'�!�ĝ�da��Cm�k��es�K��5!�L��iS��O�^q(QJF�Y�!�$�xpW��=��y�2��+D�!�dM�����JؾS��}r����!�d�y8ҹ�0H�mv�)w�	5�!�ӣx�Z����.k���e���J�!�� ��h6�����Wl]�`6��"O�D`����!i�����"O�Q���H�1���[��^�޹��"O~d��b�&:�Pu���^wv���E"Od4p��/+�&�@�]Il���"O�)�ᄝ�_l2�a�*3hPe��"O�h	N=t�j� �� v6;�"Od�;�K'!��t�I�ZT��e"O�1��x��J�2�B��u"OdXxB+ U�� �qg���N��F"OV���lB�Ö��Ԇ������"O�%�GA�"�!��;V(+2"O�5�,����2XA>y�"O. 'Ğ�e�*yqs'L�Q4A�p"OD�9�e��s�8,R%E=:B
""O� {���5t},����R$���&"O\��Ս5dWdM˅��rO��h�"O�=ƀ�);+�Y��ȔeB�#�"O	)�D�Ej Xq�%J�7��)b2"O�4J$��t���kO; ]�eif"OpMJTf��w�8�5#�#CX� �"O�mB�o5&H��kҏĈ:.9��"O�jԠ��J�,U�%�JH�v��"O ���.�G�@)�����.uh"OH%Њ&o��Y�L�ݦ���"O�)�VCH&Ol��1�L��#�x"#"O4]����Ͳ����{:�*"O�M�`
�)2�j@xDA�2Qfz�b�"O�q�V��tX|%)q�Ͽ57��g"O"(A�/P�N����/��x=B�"O4�!m�C����n��}�6!��"O���`�g�:�i嫍{@<��"O�]��Eϱ$�Z$R�-?F��
�"O��pdS���i��� ��G"O�I���8W(e�C57�v I�"O`�׆�2`��&B�ymX�"O�UC�4&�|���F�bk>�
�"O*��D��#VY��+�,7n��"O��qe
Y�0M�\1$P�S���X�"O����n�� ��9B����`@�"O �GA�m�rS�L�y��3�"O��x���!fى;�1�"OᐲM����Ed�5��"O@!��@�l�`�a7ɒ�8�`4"O 9��>`�1��,��6�B퓁"O��ȼ%��KE08тipe"O����d��x�����j̠��"O��q��Ԍ�8h�Ǆ�A沉�2"Or�iQ�A���@*E��,#NX�a"O���6Kr`��o)
�V���"O�Dr�U� f.��va�/�Ѩt�>��X?"�ۡ	EO���� F��fn��Bj�%�ޱȱA��J�0؄ȓultBb��I_�5��o��U6�ȓR�BL�BcJ�i#���F�G�r@��B$Z�; �0PRD�gJW{v]��C�
Q{ƥ�,�p�8@�� ����ȓkD�s���:V����E8
+"0�ȓoGĬ:��I>R�QHWF�5�F]��r �e���D5 X O��V���?	����*F�6X��"6�ɇ�8D��À�gY���W��=2p��I��:4鈌3�rFC�*x�ȓ j���aМ3 ��3� �=Q�,�ȓG$�&�!��CǋJ �zq��S�? ���� ŉ3���еm��fo�}JP"OE0�mXo�� �ek+tH*Ak"OTzFK2
�RD�W���NK�K"O�]��Dϡ,��-8�a�kȀU+A"OB�k�G�)1l!h�!�F���"ONu��m�<"�]`r)�/=� \�6"O�!*F�:}-� A
��;���r�"O`u�@!��H<�D�7j��p�V�e"O�%�F-��e%`ػv�!g�	z�"O��z�H̡G�2�y��vx�q3"O�%���[O�zDq�o�<j��"O,5K�@�*�)����y@|��v"O0}��J����d��P�,�"ON�E�n5FM�p��!_lpAq"On��FHU\�X����	��"O��r�V��hi6�C�X�H�h�"O�E
��&] �|��O��x�p��Q"ON= �̆�^< bcX \Ѫ�bd"Oz���H�Z̞�
�+�s&�p��"O"X����GȌu�֧�E,|qjw"O�R�L�;;�E䦐��P��"O��3%�\�8PHc��|�6�6"OU3F+�=���BB�-���"O���O)O���I��2X����"O�谖�ז�"���cGSy�H"Ov<�1��r"j�ȁ �d�Ĩڀ"O��@'f�i�.\R�I�9>.��ځ"O��3��)"eֱ�'۶(�$��"Ov����Ɩ�3�Ǆ',`�q{%"O�QRg�i�����&с'id1!�"O2��,X�{��,
�D[Q��ۄ"Ob@��u�r��c]�<Z�в"O ����(;��ԡ��欙x1"O���kX6^b��6�ڧ+؎�""O0h�rC�4if ���ɏFTv��"OFYݻ@�%���E s&㚝^�!�$S+��zł�~M(�����?�!��M�Df�` m���9BD�D a!�DS>7h\�����r�~}欏�`@!��*�RaCrG���ɥ�ޖ#/!�Z ^@K��j����b��X�	�'>�%s����M���c��=fp�L2�'���a3oP��6���Xf l��'\�%m��F�Ft0vJM[%���'p
@����y�V	��:@�~=�' j���S�|��\rK�B�b �'�����:8�^�8��=��@0�'g"�C�!�dp��Q�,����'��+l�"ԵA$��_�l!�'��48Al7�Zܻ6�O:3&P�	�'��(�#�l�Qxa�S�oPr	A	�'Z^ds+� "+F�hpe��)�$�	�'���"5�5.H3�闖p���'�p���A�Ҩ+EC�k�$q�'0�F����4��Z�^�{�'��4(`g	�R?Θ0A#�S�^թ
�'������G(K��D�L�d�r	�'9�Q��o�p�IR�`�6B�����'D��J'o�  f�[��;�:l�'�0���'������)�`�'~\Ue%�F�ܵ� N�+,�#�'�X��+�y�885jDu�0���'�`x!�sn�($�;`�jD��'�fp��hK�r�X]8'�G�V� ����� (PP�	�S>�q�÷X�,���"O��
0�ڹYö�Vl�	|���F"Or���ծGn� �":jS�%0S"OryА"�=��£�"FV���"O����ƅfy���Dؖ��Ar�"O��zF�)�L��V�ݹ	q��0 "O��@�OšC�Lj�$H�|�^��"OV�"�순Z���sDI�P/���B"O\A`��˶0&�D��gǀOd�s�"OЀ�j�<d�Z��3QY(�"O�L3�/��,����ҝPb
z�"OH�$a J����֤�^0tQU"O����Ýl]D�+"B;Y�ܵ[�"OL�KP�E;j���s\�]�"ȸ`"O1��@�E�!�j��
¬��"O��0���<j���g^5x�橳!"O*|�aE7Q�r��d�S��-QS"O���2f�$��@
RD =�2�K�"O�]9�C�	cĐ�R�D��)�f�"O���+*T0LD���v�)U"O1��G��Y[���%�
 p���p"OTP3�L�!%�H2U#� �"O����n-3�L4�U�
�@$�"Od����/L�D	��`m�J��"OzҖBLd�06`�*ؖ�H0"O�H��e��6�t�.�4��T"O��yE
V.s��qs�O�0���b�d�0>���bT�f�2��=�-L�Fd �Sv"O��Q U6mhb�Xu+KJUF�q7d�qOĬ#��Y�l�$�� *�n�2���*t��	L2D���+,N���S�6���ǧ �����4�O�Q��hZ�S����G�ݹ;49b�'g����O~b�$n�AjS"ڝ(�X��`���y�"B�+L�ꢨ�)3�xJ`�W3ȸ'b2�sK�d>]�������0k�E�#�/D�(� ��L3�D�Ofm�ajA�,�����<Q5��s��Upb�I�ovZ�Q�I�<qd��}�N5J��"Ft� E������Xi��̒�<	��`�@�"L�$��c:\O�,�=q'��f�c'�~�Q�7.Yp�<3��j]=�MX�'�uH�p�%��<�|���	<y�A;p�]�kcθ�S�p�<����%���� ��:�lY��x�-i:y���42If봭�.3p��	���W=�C�	�xh"�J* �L(F�	1n�z�OL�# /=ˈ��wN�u u���'��$;��
��3��0SbO�sV��� )��yB
���ȭ	b$�8sP�Q�.���	<#r�"<�*G�@-w�fT˂�ā�2Q'�Y�<��D�h�%�'eV�VdȅH���V�Vf̉hϓ���OW��=D��� �0!���B��|H���:�0�!��&��x�m*4��k�.�&Q��Mc���g2����9O6���:��&�2�HT�*\#@@��� �@C�I��>ѓC����7��d�Z�g6��}��Y��H�'���&L�^8�XaMV�8g��h�'0D�`s��K�h`��`�T�^��@�L0}��)\�
0��`̧]�<�)�Dݹ��^/��
kG�D� R�O@љR�G�IB^^�e����b�@�+�|��ĥ<a"�� p�4�I~�<i�N0.��=9�ML,E�!�*UQ�x�&NIp�	�7�|���~�R���$�)]Z��Ҥ���t��W�U	Na}�D�vr8uꃏ�I4r;Ѭ����D�V�dO����I<:�6��%l��;��I����T�fh��+ <��l2!�D�%97�=X�l�8O\�!լ@'��*eo�E8R��*a��
�\���Pȶ�g�? ,��a%W�<�ґ@
�kG,�PvO(��!E�^�qC�聂^�K"&��W jY�5�6���KރbA�lh1j�o���	��y�hǽI��hs��I�ax"��G>�HՆ-� �R?j��ĺ�/�R��Y�sm�*�:�˦��.o�I8��'e2ձ��ۭ\\x��(O�lw�Pk�O���@E1}r�*l�@�� 9���	r�e>�!!��8�88+P�D� �����N&D���q�rA��D��Z��r6�>B '^jpX�2���$7�� t�?�؀�j�$�Ͱ�h��c]�0>�x��,�Px�&BA �q��Y�\8��ueM�dnd�i��@I����u�A+�D�����~�>�2#�X���R����	K@�٢�LT8�`�+!}bf�6h3��V*,l���c�:>����ώ2�t��R�ȯ?�,�����mk���,ld���&�8H2�'����I�P�mE�����S�Z�Q�$�̧%��-p��GG8y}���JKa�<pk�`мtS3�W��l$1�D^y��]�lt��?~�
�������&��:K��I�hʵb䈻����y�վZ#��eCi��������R�b�^?�Eϐ.U+�Ѐ�*?��y"F�q�AY�I\�`
�ubŀO��p=��xc��yC�����n�A[�%�% �i�g�ڻ
�����'�\Ix�ݞX�ف5�L��Iȉ}Қ|�g�Euf�jSay�� �24��âۃ-�� ����y�I>T�G�[�~�p���d���'�r���D�Z�S�'%���pn��0"ҙC�f'`�l��'+H�
�ܫgB$FA�"{D��ȓcy�̩�@��n��R��H+(�HՄ�&u���`-J�^������:{�9�ȓX��J�`��y>T]�KӅ~��ȓr徥��@��YR�	��Y��l̈́��"�yF�¯�6P���i���U�6�f�A� @E�j:`N3��a0D^<30���:s̸�5�:9�ĵ���&�Ԉ�ȓVlU��N(;B��GDiD1�ȓc �<r�\l��S�,Ek��ȓo �� Pˑ +���+\*.9�Մ�qe �CSg�8��f��l0bՄȓ:�rS+L�f��|)�ʁ"^���ȓz��es��,,)�,��ka<���֕@M�Z؀�w����T ��H۠�`�	�	�0��4��>pԇ����j�K:���f��_�,�ȓ| �au�_� ]"� ���6v���EN�K!�P��D8�dQz����&|�	���V�R���L�/;���ȓ���ȇΜq�V$��D/}��E��{�¡���}�`9å��H�4��ȓ�Z��	�>�����#"q�"H�ȓ36�L�NF)sД�b�HL�}t 0�ȓ�\��@"؟\N�l�de;r�P��xB�q�*�:`n�V��13�X�ȓ7_t%b�$��u�~I�e��lI�5��]s���PL:R��dk�.H*b>y��'��	��\�2�>�Q��*�X0�ȓw���d�9]ơ;���&s�8�ȓB���D��,����hոm�.��ȓ�*��.�*W���
�؞ ��q{��s�a�*j��@a#yԄ�8�N1;S�Μ#.���)n�=��!u�Q��f��-	(���Ѩ�z��p��H^_Hpy����J)�ȓcd��a��%���f$Ί.�Յȓ;�\�S�+S�(��b�� D���nxsT� SB�`�b�8%���ȓقm0���,��D���F(j�ȓAK��!S-B�Xp܅@�.M1a$����S�? ����T�
�\��L7"��t�"O�����%0<�0����ZLHAf"O��A�Ѹ{�����"��W,80c`"OV���a_9�}kW`C,"H��B"O��zC)ŀO��	s��--�Ll�c"O��!��5�d���;&��B"O�� A�?XI�tRD��x���W"O�$k԰\��P�R"$�DYD"O�	���6'�����F�J�F�S"O��և�G֒A�a�YnrZPx"OD=�g"��̉%w����"O<�H�,F-~Dr�`̇!��Y�R"O�h�/��(*4�Μ�a"O� �j�3 4:&̓�8�K�"O�ܡ��2*��R�6A0��yF��Pl�8�V(ԅ{&�Dz���y�I�i�҃�E� "N�勛�yb
��s����e��{$>�#%ƛ��yrȡZ�X��E�m�v�Y#�y"�֜rs1�¬Y���Xd��y��PF$0��a.�(yx	�L���y��aqJ%���  ��ѥN��y�J��N�[e�sVB�A�l�yb��/,��0��%����gh��y�ċ���Bğ!CC�8����y щ@
<�y�n�T�P�Xg�5�y��ܯ:�vEP@5N���j��yB�,}�$Bp.�,O�<8�m<�yb�,,��P�%˸r�19SKߍ�y��Q�B��H�7n��B�O���y��C8$)d���Ɨ1�@��L���y`G$x�.UaOT�\ĸ��G
�y�?G�J�H��N89@�N'�yRɏ�gbZ좒+ƤN��T�&瓫�y�iF5��He��;��Х��y��6[yF���c�5�b��8�y�l�=�N��`��{y��4�ӭ�y2�v�@�;�)#:���WJR��y'H /m�8��"����PƆ���y��i$��:�eӯ�|��C	�ykMo���;�н	��x�%J�3�y�⊀_P��@�kx �5�uE��y��*c*M���+`����HS��y�.׭<A�i��)W�v�[u�>�yb
�,>P�ѕ��W�t��$�L;�y��=�EX�
	�D�ޤ�vnЫ�y�$[(O�0�!�C,2�4 {�JӇ�y2AX/1hr���Ƀ*�� 2��y���1?䅓��Q�3F)�"���yb�7'8�bPlS!�̬�!���yr�*.<��y��� �"����y)�S7f�H�nݜn_�I�I�>�y"�
l���ͪ
?�����ٖ�y"Dύd�^m)p@ʎ�PPP�Ŵ�yKЂ-A��Ʌ`�:dR`h�i���y�%C�d���	"��$SX�ܹ�b��ybe�l>�Aac�ü��-��y�X I0:�y���=�0m�N���y�����g��R�����.y�'s%�#�J�J��W�K5tK����'UN�Y�W�"�(�C� ž���@�' �ʕ��'`��)�s,�tp�'�ƀA�`P�t��٠�fY*Q�0eq�'�Lav�\�*�ҽ�iBaJ��	��� �xR9ؕ�&�%>�D��"Oj9�t
ҁW5L�(Ҧ�R�|���"Oj b�_�,�.1b�L�"��"O���0�C7Ȭ��ƢJyd,�"O|�p4��L��oۙda����"O�����ٽ#K�8����TUZ���"O�ݨ���HԚ�81�G a
̒b"O:DEg@�r(��d��1wP��"O��x�J54*F��2��Xb]��"O."�EU�2� ���藽}ĎLaG"Op�`�I7Oy�8A  ӴZ��(�B"OQȂn�1W$hԣ�oG7p����p"O�\�����!$�Q!�[�����#"O伈�V4@.�P��ز�>-9"Ox�1Яq%(\Y6M�,
r��E"O.9i���%o`����	�Z�!�"O�H��膸gD�b
Y"���"O�uI�f��Q~\1�a5�)B�"O�t�� ��4=1p&�v���Q"O�5跬�Jर(Fo�=	.�aY�"O~��ģ��3����QB}��"O<��v�5��Laظh���ׇ>D�����X�"!ȉ�2ڏO���3��>D���1�?W���#�U�����=D�X,e�t)��O�c�(�wŀ>�!�$�	]���g-ҷ.�<���(:�!�D�#b�@�o�%�����d�!���!�p��į<��� EʴG�!�䚢N�h�SP����	wӥ�!���h�j7�=#x�8[�W>q!�$M��:Y��EH!(������W�cL!�d#8~4u8���:pVa�Ì5'!�$L#�\�z�J�+�*�[7@�8m!�C�/}�$��L�8���s@z�!��(�(��]?wtL�Q��5^m!�$, -���,d�֠�Q`A!���"��D3�l��R��W 7B!���)v��-�%C�������'!�[�0**��ѣŭD"J@����+~!�dU�n�\) 4b�
rH�ʢ(!V�!�$�3E��X�p��!�8Q�'�+�!���Vb���"��-h����+!��-�����H�%=�"�hUi��=�!�D yЌ���H764�dc�� =�!�D7*:�C/
�Ϙ@�5"��8!�$�Ta�1B�Y��B��ܙL!!��Lo��36K'�4}�F�9#/!��S��aS�jY� ��T�d�,.�!�dD�Bș���]���G�U	�!��>��`��"�<��ظ&!͗Q�!�$�0W{=�5$�	�$qq���x`!��P�i[��cd�;���P��"5q!��τ8�Z5PQ͟`�ޤ��'OP!�ʏE&�;�NB=V�r���4Q3!�ͯR��%P���jT��k3��� %!���8z����G߰j"yB����!��ڸ`���pfNV�H
�0��Ӱ?�!�$ �dJDƛ�T�fM`PL�$�!���6r�	acA=`��Y�N���!�ϖ5��	���Y�W�D���T Ld!��	�Bo
��/�kzJ��*�5!�DO�\I����ʕ?R�unS"!�D�;i�$Aqc�YI��s��!�Z0n-����A�0|��2�!�� ��R���jȾ����A���b"O@��1	�F�88�~�:ēf"O`d��J&FW,{Ud9J`a��"Od5�!U��0�a�ۋun��d"OxhB�f�2hLʤa6���Y4�C"O�Ic1�_�]%��5��-H���v"OZQA �E��ebv��"5��5"O��ZdN�7 �(��
�{�r�P�"O�k#�_�q�VΙ�i�돍r�<�"�H������J�4`i0ARN`�<�d)2x`�P�NY2z�v�X3CV�<9�ߢ����.�`ɶy�v��i�<y+�e}����N_�Rp���� e�<�A�[]5H4��$m���4�
f�<Y"��^<h�3.K�(�ՏO�<aO�Dq�śC�0|�HР|�<�e�X&�� U�� �:@���L|�<�3E��_3d���^{ةk�,�d�<��h��q�B�\�G�<�SA�Kn�<����<-l�*��2)�R9s�c�e�<	7��P�
�䋇�Ut���~�<It'�bI�0�G	��+�
̒1CLz�<&g�(s����)���VF�_�<q���(]�� I�= ٠ġ� \�<a��˜x����;>�FH�K[�<QR��,5VTC14xI�s��h�<9-�:���gn�,��D�q�<!���2��dӇ�X�zn�ӱ��@�<Q���b����@.Ót�����G�<̙�|i�D���JŽ���G�<���� }�]��� 
��3�Zf�<�A)�1���"_K�� @
�HzB�	6���@Fe���X�'ٞt�DB䉜}k =�v,gx�����W�PB䉌F����eI7]Ӫl���_�"�C䉕-���!U�`У��۸W�`C�	3If�m�0�� l�"��e�Z.lYRC��'J��$��G�4�r@�]��C�<R��%	F����CF� H�C�Ɏ� C�䖪3�ֱ�uJǍod�C�I�H#�d��a\3ex���iB�e"B�	��L�*D�G�$�r!��6nvC�Iv�8i2��B%x�cï�""C�ɾu֢PZf�БOB<i�w��<FC�)m�x�C���8 W��8Da\C�	�%r�*���B"��質N�W�C��9\����ѵLu���6T�6C�ɟ	����nǋ �+ը�x\C䉌6� �b��C,L}]!�H���B�	�&9Bi̝3lĴ���[�M��B䉤�6���" )��eBs�?A1�B�ɀB��١iH�#�
#0���>fB�	�w�H��Ƙ�3zⱊ�i
�8�xB�-���EO���h2�Go�\B�	?tk H���*Qy����3�"B�	�2&N%�硙)}�\h��0((B�ɯa1�xÏK
i���*hF�a B�	�XN��J������C2ov�*C�ɉ!-2�*ܑ�:٘5�ԓ`��',NI����* ��B�D� F�H�C��A�p��C�(�+0#I�s���y�/e�����!W1�^ap�W1�?YFJX+pk�U�7[roZ��ا�ɗ$aN5��ɱJ����aO�.F�O|��P�+�)�i�P�A�� �V�g$�8�'A8�P���ċ���" �]	���W�x��I�9�H��?E�� ��2�`*C�:%�N!eE��SA�iG�Ku��ӏd��x���3.�5�
84�@����f>���j�10����?y���6O$��4Al���?%>�@��ߑ{� �%`X�m�@�R�
!�d�0Fڮ�b?��E`�PP���Љs7�H�Cɹ>i��Ĝ���H��`�s��.t6t̓ �A�2��x�il�ڕ��S+:dJ�51҄{ c��F�r��A�dn>]��*=5(��򫊛+�&YyǬ ��#IW�5�?%>!���0Q���BH�/mLHy�QN1��_ۚ�b?�k%���B^�e00O3D�8s�N�>�������(}2+��@�H���~�d�Ƀ�8�M�� �#���ȟ�1򖆑�9o��B�/G�Sa^Y
P'_���' ���	�������*�L��K-_r�OnD�B�7�)�W4Ir����&m��"C�!z��';��D���Rn��5�'���#�&�����c����	\~�?E��Lͯ@��-����L��|�PΉ�M�h�4���ȟ�d�s�H�_��=ZvI��L�J�!�=V�O�}l:�T���p���p�-ڴ�܈u>���$4��P�=�v8i�"�9Oe�%�ȓB�,<����@�����.�ȓ)��1���&���;2'֩;���ȓh,� �U \�o��%��E ^���ȓ^�pp0 ��X�(L�"��L��хȓf�N��-��r�S�>�ȓV�b@��:�:%8<T�݆�&���pƒ �<*�%�7x�l���|�\�ѐʞ�d!���z7*�ȓb	*�CbԞe�^|�7!�*�}��i�ڡx��S�hCa��$q��ȓ>Fl����E*�v	#�B�4)��n��P�i\I�D�7f�J��݆ȓi�T�B
�e�dj�;����ȓN2"�q���&mqԕ��BȌ;P\!�ȓig�]��@�12�� �2ad�ȓ}�"�[�I��b�y�*>S'xi�ȓox�`2�'��#x���B/2�Q�ȓ��òE[]T�!�ԁؠ*����G���i���%N��4#��� *:4�ȓ��E��L�E�\����F_P�h�ȓmXڸ�@/( �\�k�k�LҦ(��T2-*��N�V�$	��x�t�ȓ	<��$���ޡA��$+� ��"�P�·N۱.d��S	^HFi�ȓz��cB��I+&(��X�	�p�� j2�����W�4��ԠǏB����L�� �fG�E�xY� J�N8�� ԉ��fK�1�Lɩ�E(v�*h�ȓqm���*6��ɂs�۟M쨆�N��%�d+ �����e��G~�c��	�X�r-V�bU"ͅ�EȦ�8u�;c�А.�<r��)��q���Z ���R�e ��a\�M��@�b$�����Z����i�1>~$��s��ڲ�.T��d�g.E��Ć�qrz�/���Ca� c*��ȓU4��΋nf���"�B��ȓ`�|�9��K) �&�XŁW U��#'(=�S!�)݄(�F���!ra��_�~��F͈�<��옰���^U�ȓx���ЃJ�Bp���e��C��Q�ȓ[�"�be��0�f@@7�Tb�RX�ȓ����T�Q�*�*%HU��*;*�ȓb��=��Z+ �R�S�*��Dqޑ�ȓ$+&L�wY�z����p�`���S�? *�!��qR��Pf�v�]ْ"OΝi� ǂeW�H�'��R�Rd�S"O0L0L�  tz���\�\�����"Oap Ϗ�A	bA�8PU�r�"O696�J?mk����۳7�<��"OJL�d�:H�
8�憊hV�� '"O���:"<��5�$a�3�"O@)�UG���~����R<N�,�2"Ol�Z��O�<�@¢|���"O��J։V*Y����u �r�I�"ON��R��9��@ʐ"Ǵ�;4"O��C1
�6c��ؠ�GF�K�J���"On��@ѫ|��� mV��:I��"O� Z�D {����`��<���#"O�E a�ءgͮI����T1"OP��7?� pR��N��*�"O^��(��68�q��̄2��i�b"OĤ�Tj��a�~����[Ȱ��"O�̓�\D5|p���
����F"O�PHA+��d�=˓��8��0�"O�*/ 	>Ԇ�aU*$�Fi�u"O�}h!�B19��*BG�Y�4yJ2"O��CG�
�Wq4X��*}FL��"O�y�3S.-3��h'�������"O.m{����B�!vN��>��сs"O���l�"�ȴ�쌔8�Bt�7"O$,��0V)��ƃ.���B"O�E��J�z���
k��5�"O�0Д��=��6GN�!��<�b"O�!{w	�G�,@h�V>;�)+F"OT�Xƫ�=Y1r�I�,�I %i�"O�����"{�,R�Dɏ5��A�"O���N�.LIPع�a[�)�ּ�"O,�6�ƫ3�x3aңe�x���"O A��h�<lf�5#����y"O*�s��C�vY~,�p���8|��"O���Qo�K��M�a� Y{hɺ%"O�娑�F�)v��B� `��ȴ"O�1R�5<�$��N��y0�=�V"O�e��2`	��*UhJC��\�"O$H胎�w\Y��'M�:�:���"O�M�УL�����fJ���x�"O�a.�>z���*l=�iW"OJx����tl|�H֯3\(L�!�"O1���G<�@�1���8�"OA�`�
�ޙI���<h��z�"O*EC�(O�3�rY��Ml��%�7"O��ۤ��?׆�k��K�z��Q06"O�wf	�R�h�	�,D�"�2]�v"O��e��"9\�Ӣm�,z�čA�"O
)���T�Oڍ��p �"O&� ��)*X�Cp�3B��Bq"O�Y����[ʾM��@��0�l��A"Or�б�ӗZl$l�J���I�"O�9�(�,0��o&Vh�"O�$B��݄��ӱ%�H�	��"OZl±��S�l<0 �R���I�"O�-3r
�"#��!#�c�C`8���"O��k5�0g��Q�"�e���ɒ"O�9��Z5DWZ���aڞ+	H*V"O�\�q�\�/L�L�@T&(�W"OZ��'��# (s7�V
ACx���"O�`���'>[<`��4d�6���"O�� ��	`�8 &(�\���"O� �X��K�0j�ua/j�x�"O�e�dk�H� ����C�"���Q"O|@��c_;*<́cDǠF�9��"Of\
ǬŒ
)F`:���3.��"O�(�����&U��Z�f��hHst"O8�����s��e�vǏ�v�&�"OV���I.t��4G��ܰ�"O(���5!d`FU�44�t"ON��ejV�����@Ҍi���s"Oz�BwȞl.�p��WiY���C"Oš \�>�&�:e�ޝL�$Z�"Oj�r�G8F0`���Կ=��;`"O�`㑬�'>��b�iE�5�b��"O���Sh�.[�lUa���.��4J�"O<PQ�� �P�u'݇8F�$H�"O2�a���>U���dG�8+t�s�"Oh���,\б��>( ���"O��C�dS���,�<z�"OI��K/;���!,����v"OVԙ�̓�r\(�� y�����"O�4@���=cBvtH!H�?G��,�@"Op1�ޙwö�#�	M �:Eq�"O�Q
t��6�t1cw)Z�Atΰ��"O��#��,Z����&�mg`��r"OZ���a�>\�l�e�=#g ���"O� ��`�2뾡Ab�8In��C"O��pe��$�=S'C��FAD 8�"O��f��w��0��چR4t�v"O�U-�2h1 �i� �S&(�!�'����a�ݲ6��ySк�ЃFo*D�$�C;5���!#離�RB��$D�p����F��y���+Lkt�C�>D� ����p��J6�#[!�8 ��(D�� ��"g��A��A7d�jp���'D��Ҋƺg,�0*ǥ �4p����&D��t!B�tzn�9��@�	�(P�c�6D��w�W%1��l[qn��SҼ"�/3D�Ty�ɠ5����d6%����3D���V�*t�0E��<�0	Z�-0D������
c4�@`�� �T�{M;D��z5�D8�Z5ZSBS:1td��4D�@� S�H'��#��RLTS5�-D�4)aMʯ'���@��P=�W+D���q�P^uqGI	u��C��y��L=^�*}���)��컕�Ӿ�yҮ٤�TZ��ͥ>��ɕ��y��Rz%��V��uҗ���y�F�q�G� .���6D�y�+I~S(I`®͉�X����$�yª�O�X:���>P�2�MϾ�y���5U��� ��~��@�l��y"D�!$��⡮Ҳw�*��7
�&�y�� �|=��)4���\��Yx7�\��y�Os*�rV��Q��piW��yb�=,��E���Kf�( �5�yr��e������԰���U��yr&��8S����/�yRe 0J��y��
8=r�����2�A�R���yb)�}u���t+O"J�Q)%*Ў�yRK��N�|tbDRg0�� W�y����X�H��7��d�`�5�y��#>� �"a� sb(��Ï�y�K�FiT¡ rj��?�y⫘pj�J֨�=y�x� I­�y
� ���@�'���/~\萃"OVP���
�-D�_�	!t)�0"O��1�nQ�4��i��
���"O~@`���&>�0�n��Fu�H�"Ol��QD�+j^čr�fL�Dc���"O�I�!Wu��:Cf5
��#"OL��m�Su�A�D%S�0�X8!U"O��aK��-�1D�DєI� "O~�b��Q�p�N��� ��)*�"O��{t�We�̡Y�;,��{�!��U���m**�İٔk
�m�!�XD�2<
�h�s|��V.}�!�گ+j���Y�s^����N]�!�ܗ:�<� �?aV�ݠ�AƅJu!�D^�_-~�'l�!A`�`���s[!��u��[�`Vv2P�%��+z!��Z�E��5�$�������]��[]@��@��,��h��x���ȓ<H�9���R��u��b�4� �ȓ5�NQZ�+��-s^1z��\�^G4��ȓ�$�'��<h��v+F%W*A��Vg��J�&�<�u��:m��m��thb`�cC,i���F��Z
 ��'�0@;f��HJȝ+�9����<��*尥1�b��#}ZU�[�a:
$���L���Y��c}�$�O.��u��K���be�J����u��&\���T�O��������}}�U�R<h̅��}"
W�A,u���^F'��Q�#�K�H�	D P?�u�� ��9���V��ك�	���'�dE��.�� �~�E-ڎu'�}�p,�t���{$*޸Y��O<��<��oo�9#k^	���r�J|?y!�I�M�i��Ij�ղ��V�x :<�2�ZC��x�#�(LD�V�'�i>�|�Wٞ�Z�)��`�zD'M�kΞ�����q�x�/�5s�ej]�W�L@+ϟ�����y����)��X{0L�QǸ�qH��f|�ě�*�/5��c��c�LX��� �(�&?�a�w�<`�AON�(��I�%e�������?��i7�ʓ�DQD������-��|t�L��B�~�� �	y��hO�4�4D,��2���L���Ҹ'O�7�̦I�ɮ�M���J�'�M�6�\�!�p�Ҥ]!���Yd@@i?�U@	�)���'R����:���g��3�dA��3D�.̸M�VE���� b&�*D��p� ͇�a+�O�鋲K�
c�ڼ�BI�+�nѠvGU� ���%/�><�����
pm��Q�$�>�W�K�uN�+\Tn�DS�����q���O��o8�ē�?����Z\a�vF]b@�ac�g��L���?aC� �>bU��'ZUa�H��/6b*6�,���릕�SHyb�@�<�N7�tӆ	����uњ���G/Y;��i�˟���͟d.!�����O���Q��+�x�>@��l�0R�Mf�U)�}( ��#B�攛��S�aѣ,ʓ6T"�jÆ�f�k�X�bR�j3�F/�
T#�]_J�Qc�7S�x��
�tP���*��J�t'"�j��y��j��Y�����Ǻ[C��K�Q;'����<i����d=�'(��yƅ�!$���+ȁvf���p�`�µ�V,0�pE�� 3<�$ �!\KH7M�<a3f1H��.�Oz��=�Uhװ>)���T/w �q'̥����a�Äqӎi�����*�@oڙ4 ������?h��J�8�CI�;A�h	��)�	�.�e#���$Q(��f 8O&��Q��*u��]�H����qDH<p��c�W�c��Тa�O�`o+�M���ħ_�d؋�O�CY��CҤ��3�����Y���'���Y��v�^�	y���d*�U}�DSD/2lO�6M�ۦ�'F>Hf��'n�dh�On�1�`�<~!���pb�O ���O�!#L���O��a�,<���_
y��@�&��MSVI�9-��Xxc�O���"Q��,��HFQ���O��ϻ*�x���2?�o՛� �a��+.`�p��K�%��-h14�8 ���GZ��'i��.A$b�V4I��q�x�c��7}��I��M�2Y��[��3����|��L1f`�c�	�⦔���-��[�N���)�(V3����葛*
x��sdT���'�7��ͦ�&����?�oZ�VK�+b��	]܍*�܈q���'�a}"�+n   ���dc��Nɾ��V"O ӆ	�*��ՁC�Wa��h "O������F��a��gU��6��"O����(;G�0v'L��Z���"O}8��b��U�5�_��CB"O�A��2�8��¨��
;�MB�"O>�= �t��f�l+v5c�"O <[c�[r�uhF�N�D�\��"Ox�����?��D6f&w!���"O���ǱD�X�b*rn(��"O�@�s�I�
�@ w���y�"O��Q�%v#��r� 9G�4I �"O�$�qU=Ⱥ􋆩.۔ ��"O���\��<��*�_�$�"O��y3��<g$a���Ϋc/nr"O����Z6\�\�k��� $)��"O��w)^#<|R��N4Z���cd"O쐳*�SH*i�e�!w �W"O�X���"&��@�A�xՠYB"O�eű]�e�qI���8�pC"O@�P���^�����He�֙�"O� F�H�4iӋ
��Ѫ�"O8t#��h�p%��R������"O���@-�.g�ָ�� 4|����"O�PrD瓂,�V-x���0�����"O�$�&FN�u�@��3++LY"O8�(�/8
�h��«�I��L� "O����矆bp�Sʉ�.�t%l"OL�� c�?zr�kRJ_"0��AT"O��Y���7&9\a2��Ǻ.�F��"O>��uɗ��Q�@��dБ"Oڬ���	0i���&
��!�"O����j֪A�Ań�Xb���5"O8�V�q��W#��@y؍� "O.M#��W:5�8	���,a<YҠ"O�x:�M]3ƴ|�eB�gCb��u"Op@ZD�����+#�4��ٺ�"O��s6���T�:M����%�\��7"OF�H�"A�*dE�e��6Fm0�"O^P�SS:d<^U��k��'9���"O�H�f�G�F�F� ��%6��!&"O\��R >}�U`��Q�&"�]"�"O�˓SPNt(i[9��R"O��#[�xQl���'t��W"O�{&)�
�v���$K0gO���"O�|+#���,(H*u.W�,\�يg"Oޝ��ˑ��;AK�7 E� �"O����X��4�ۡ*�-{����w"O<�aV,L4w^�`��L3�� pv"Oq"�(��E9�3IS�t��]7"O�����U�:`]����W�����"O�ЀWo7{� -b��ӛS݊��"OF�@���kG�Jw(Hh"O� (@d�\�& ���,s�踩�"Or)hFb°2v�qX��>����"O����Cɐc���S���\ ��hu"OD�rE�c*��,�_9p�S7"O��2��M&[��JpeȢ'���"O�]���Z����c��߲Km�|��"OB<Ѧ���ZY��F�/�T��!"O���v��%H�,p�Fpz4Q��"O�s�@_,5P��b�\1"O�Us�K�"e6(�oU9dTya"O<<J�ɟ�>�Tppb���S>��0�"O�� QM4lh�l�`��r3ڜ"O�� �ğ&���&a,���"O���3*Ⱥ��]@eD#3nX"O^Q�e.��΀ te#<�(�"O�|�Q���2a��r�H�u,JĚ�"O �󱍙.q1Z��V���nB��`"O؈�3'�'��j�o �dF�
"O$Bw���t͸Q6a�fF�9J&"O�u;�N� |�<ڔ���K'XpT"O���� ��)s�ǳ�r� "O6�S��Bs�F� �Ή/�J��B����	�8�,4�ѵi�?�"2�H�Y��Uya�ȡ?��h�!������H(�]�Wn��;P��8p�S7`�Bɕ�Ђx��'D~���G�6Br)���.v��'����&:}2�����!�����AH&?��Eӥ�~b�h�4 b��	2��+2@y��d������H|�O|�Q�V�|7��(�8��DCtc[ܓ�?Y˓O�:�GN���+��;��X�Ԥ<�Bm�dr�rO����	�D0�x�_�QfʑaҤ�޴�?�.Ox9����"=� hUrp���V6�i"�!�#?�U �ńkg��p�U'h@��˟��[�y��$�w��U��)V'9�p�ʗ�H�[-�(���I���P�H�����M�Z��%?e��eC�y��v�\��� �� ���'�b��m������=:����?ߴzh:�s�߹����cH��l��w�d;�S�t�C�0;w�Y2BŃ�������1�M�i�e�������ɨ~�1��6IƠŸr��"d2�[�lRq5��{Ӝ����O�P�����Sj��HY.���A����d!&�s��9p∙�+��,���M�'��\����K��d��@�@�V�0� �$,Pt�5 ʉX%��2B�^��On�+�ʅ;e� 1'���tc!!/�"�b$rӸ�%� �Iß\�>�`�ғ'HDE@6��3AG��C���!��_8"'�q�J�.�����f�>t��'��Z۴[l�&Z����䍦�M���Mۅ��7Q�u*�F�?5���H��]�'N��r��'���'Ph�[����b�زRf|���C)��`�L���iV!*����!���7Mݳ@1Q�BWd^0v8>�h��C.yr��21��+��q�-IV"ӂ!L�	�B'�'Ը���N�;'�V���Φ�A�4�M;UoW�U�RU��%��,��G�S���۟L�'ӑ?�q
 �o��\����׌d�F$'$�`p�K/-f�5��(Y9-��������:���nWyΨ�L$9��'��O�\6�o��8�uF��e���x��v}�|C@�O\���$�Td�� �q*�k�$p�B�']:|�R��ח�0�R�h��R�i$�T�\��J��L�M�~)[Q�u���Y`ͮ~2�ꋢ(���8��Uz^Y	b!�B�	+4�n����0�4�?���aQ�\F`�����"2M����~"P� �I]yʟ�' dW�Ġ/�8)�鐴'�D����M됱i��'�Iڒ`W�u�ĸ��_Ċ�X���)M��?����?�@O�a�j4P���?���?1')��Z��@H�<}p��F ̞�b��#�ň8� :�CI�Y1<�q����䟸mZo����t߂ ���I�:+P4�#�@�/?hea4�"00H����8)�x���V�d�L�*�@�#��ۼC���|�y�� �^m|d�� �t�6��gy�c���?�}���mZ�w�L;Tb Z1dy����3)�JD�N>����Ă�'0e*ԓ��³O�D�POŲ���M�R�i/�'F�4�Of���S�<t�����&=����3a7���Q؟`(   ��:wP=�Ƨ��2T��дa׊������}�Ii�c(p�� @�?7�'�d�8��f�4�&>]n����l	V)��R�=�MA5'�F�
��������?J�,"f��+�(ѡ1(D������"�MS��iO�� 굢f�Vg&=�Ǆ�����>i���?O>��}b�F�| <  �	B���K��߱�dy�B�K5~�i��A���Oh������+.iZ��49;���3�4��<[s�Of��c�
��9�|�R��E�3(ʈ}�ˀ�0�rԨ�(�0zN8��M��� �٣O �X�!âͅC�*0�˞z�XP�"��.W���^˦�YO|���=� .�"�r�ÐB�9c�p 0.|��?E�d]����ڇn��dqP��2&�L{r�8\O�o��Mk�D-�Qrӥ�:^����� 0#ʰPh'i�|<6��ĸi��P�����?��>��f�{)ɒ�"�:=��L��DC:8l�م��79N��p��t$J���AG��)�()�w�����A�%G�^l��O֯|� �P�0v8�J��If�dy���$�H���&!���yG@��!.�����4K=b���Y-|��ă���*Ol�#���O秚�}E`�3�i̘9ޤa���ׂx~�d?��g�'�(}�Q�f�򴻢�7V=<���{�yӰ�l�d���?}�����IUn YHh���\���{����?)�b�.5�YX��?I���?qR��t�D�OP7ω ƞY+��H�4P2�s��,x?*$��*T16v����_	Ȕ̊����M�U CI�JʊdY�`]�r�$i!�˩H�M��N�$drakp���w��'l�ϺC ��L��HyaB���	����S�	�l�p߈U�š���A��oo��g�f�$�<i����a��eڣ(�9{�9�3���s0�	��"OEY�`	y��Qy�� a�m�r��MKI>)�j#�Z-O�|;�麓ڴ'��*!�K�U�H-�Dg��h�����L�7F��Sp��r�jD'3ǚL;�HڮM��2�ؿh�$�	gL香�F��f>��Fy2�ַK�|�92*UR\ikdG�3(�DE�V�6�����
&v|���	��SU��z���ʶU�2Kv�����*ݾH�����Vo�<G�A'���D�<���>�g�? ��h�*�7v�P�A	P����"O���G�Z_���i8z��ă� �>�|�0ݴ��d���խ��?����I�h�n�� �T�>[M�p�E>$;D��&��Oh���Oz�:�D��_��%�S[�>)�Iq�n�⺳�h��uBE�(^T�R���	� �ʑR���'䘬J�ED�!z�PO|K�X�G,�){Y
$yRF:D��f!�;.��F�;N�8jg�|��;�?��i&��$�'=�.�p�d�/�*e��s!0��=��O����?��	Wd5�bS4z���� a��I�z�ma�h|m�T}�fѩt�u�p'�N艠��_�~B�'p��|b�E���   �)	�<pnE[��N.���Iр��z��z��1�`�%�ɋ�����
���\{b��}�>�@ ���?�P�i�^7�O��?�/Oz6�P�3�:c
ͩ)7���åk�!�_�5�L�hۉl\�i拔�k�����4��(��������;A�0��;�M�SО_�Vd�ŀ �Z���0.e�����O8�d�*�����f�'�,	6OX��D�@�ܞj�2� r�L�J)�<�t�_5K(M9���,6���Q�d��C7#D��1L�5��V-� t��A�d��02�:�A��LX���Af��s.�+p	�E�I�r.>���ǦE�k�m�j���<_��H2�Ӥ0���?1������7��A(�
N�y��O<k?Ρ����?�@	��dg�� a�Ȣ(
�|�S����7��}&���	۟L'�pnZ*"M<P  ������{%b lӐ�mݟ��OY���N'e10mj�F�2j�xq�e�O������O�a�݅0/�e��ɋ�z�č���'
�&x�*6��+}xZ=Ì�,���Ũ� 8���x#f�df�Ob�D�|JTF��?���Mñ퍼0}�Jd,ܢJΉ�@�"�Pt�PP�T��3cb�� ��B�c�% ���q��O�k,�*H���v�Ђl�
���Le�v���j�h��K^��0��A/@�'��R�o;7����Z>��S���q%�5S,ժd��?��6M�=~���c��X�����i������J��AgHş#v��B�'22�|��H%37fW�d��K�-�U������M&�i�'V�����m��0� e�I��[�\؞�`W��
��)A9Z\� ��.�.�9�iŪ��&JMs����� �J�T@,a���g#N�*.�s�uh0�D����z�ރ$�NK��bӄ����'ӌ6�hy�������^�#".��"ޮx��h�,
4�~��'��'�ў�I=..�L������A�* �Q���ݴ��|��O��.�)@o��v��[�x�p��6R�'����I�d'�� �\P�#f�����P�
�@�N���i��	L�@B_w�Җ��	�&hz��YÇB�T��U�
�_��O������<#iC�	2�X%fdӘ1�!�I/|���7q�|z��Bq���Є���O����O� �@���iSu��x��ǃ��ҺZ0�z���Ȋ(C��D��y�B$a��Ml�Ο�%>)H2kP�ZV���2n�xPPAd���$�<9�S���G>��X 	e6Is�$B�a{ҾiS�7-�>9DK��B&�-:q��w}fy�e�_�C�๓d�^�S��'��O&�a�'�b�'��6FN_nX�pv-�)�$��R���q4@��ğ�S�zɐ�k��֜`4� �h Z˧�"P�q�)RFŇ&n�2���nLa�B�H&�Yt�ȫ��8��9E��	#A��cEG��\����Y>���w��k�JէZp�Rr����`����O�\n����$�v�>��w�P`"��FH���1LC-V�rAb��O�O�=�O�~�"�
-H`	 !�K���ډ{��k�քo�n�I�?�������`I6k��-�@(_�d�T�ؗ�2}��'/FT�@ ���$YY��U�,�`��C%	n�J�<qT�%o���pE"Y/� � #�W��u�����1y��� K��)���Y���(P
��Y���I5�M�g�~�)�%���[E��"+:�ٕ�Њ�B�'��O>�nZq+,[BO�@�������%����d�٦�{#�^m��b�0ќ��E�3yD�A$�����p%�\&���t/   �<+Q�@�i�R���	Iy��酌P
 � ����$����z�!����8Q�ME�z�mq�%F�qR�J-r*�oZvy�b�&Pz��ßX%>!sF a�N��q��l�`*�Iϟ���/8I�5�k2,mZ�b~| ���@�#����  z��!]���FyR�ֲ6Qʬ��%Һ T:�bh�o�8A�3"͞[�vM+�f�9��H�&J��  ��Ğc�m�ȹl��L�π ���ğU�2��ed�2L��	S䅁�,�'��)��0!�H>�z��Z�zl �+4E)�O&7� Ц%n��qQ�̖yX�t���Cvv�	>\�̃r�[͟��IK���Ǝl ��'Y���)��3���-*Ȥ��ě ����S�bx*��A�>������#�*������֘�dd����$�&(p��"�`�:d��7͆	�����B�i���
�!_�,̙�M	y5����|�1q�r������ �y�� ��#��uo.Q֞�����K/O�T�s��u"Q��i����'�"=���jt�O���+�$5��?�iC�Č��E�d�_�*�(�6ʓf$�f|�(�O*��m��7&�x��Pw�� xRy�C ���=y�k�   �c� {e�� ސ��I �	%?1ђ��ji`a&Y%.4�$��-�>IGK�֟0�ٴ����'�>͓�M;}�F	�5A���Ӭ>}B�'��@��Z$�-X��(�N�B��J�J}�'�L6����'�<�AnƵ'�Z<3�L�RB�S�L�2yf|�	ٟ��	�z���k�8��֟��	6y�N�2_�Н�^.',���Հ�E����	-
9c�ܪ_Tq:wן��	W�!��YsC\�� ����`�zL�xؔ��K��:��:oXU3�$�UbPU�Û�co�O�
433�ly��8Y�2Т�#�:PJ���OJ))j���'�D)��	�����'��i�(��P #!�H%��/P��r	�'�xA�G�f�d3��!$(���K�O��n���M�O>A+�r�Z"dr�d��k�z�H٬e���0�$F�����?����?�"�����O.��*;�j����Y5cM�r�NX��I����N�R��i8r@h��i72`�U�N]�'<p�͙�uXf�� I���ڕ�!e�!�c����7�,m�*�o�%�(OPrP�i1��3�)����s��n@�����e�L<����?1��'X��l�!C��b )��JT�4�@ͅ�/�jA�D��f���	ăh?"إODo2�M�+O|3��Dv}2�'כ�P� �'Ć�1�x�k�Η&3`����#CON���O��$��k�2;Bȉ��@�I��B�pV
߫Snf��!��+'����%'�C�I�_o�T�V�ͻF�y��ץ�X�J5�ɟ:u���6%ʝ%=�(�A���0JX� �	R�$ܟ�lZ�Ԭ;�B�R�K��ا��4N�`���?�������|P~��^�i(���UK&�|��'��6͘=(�D� A ��$;�H����7Lr��jG��<��	(q֛��'��_>�P�ώџ�nZ����)�c۝{m43�������rt	��F��W� �����&�B������A�:.���]�f�{6N�3}L�݊U��."��WvYb3)Z$3+j�XH׆��T`U"&����E�EӁ_��2��4#<����S�����O�m:�M����H�4��ⓒ)�U���J�3�@��>9����=aA��)=���(g��Aʰ�*�ў�PݴD�V�|B�� ���mʋth���xy��G	Bݟ�&�l��
I�v �   ���;S��A��[�`�s�2��5hĬj�����cM�7�#���d��G�*�y6&��Ȑ��HӘ��D��1�f�O6��O
#}�rAF�Z5 }K���Oپ��Eh�b�d�O$���*` 
@��iǣX��I�$�w�Q���ɕ�M���i��O��F�-gV!�U"D�/�Xt��s�j`�I䟰�	�D�JP�A/Fԟ��IƟ��	w����'1��`r������a�ׄƮ&�T���?}��.�IL#�؟2�i�G�h�ksV���I�f�.)��ǂ���
���L�H4`��2S ��P�� �6�d�y0���Ċ�9��#eL,\�KO�>���y۴�?I��K8�?	��3�Y���	��Y�����+��M��@K�LN\���#\O�c��ڄ�͉Of Q�`�)�]�pï����4�v�|��O����xh\� ஬��%��(�(�2Gbȝ/��C��g��    ��,���!�!�<8h��O��oڻ�M#O>Q��?i�OH�	$`@�?V$Dp���zL�����>�j�J`�O��d�O��$ۺ���?���.�8X��JP9
�6��6b�:l ��c痐��a�3�Ϸ^#���}�&D��(�(O�#��ڸ_�����[�8�,��4@�#ꍻ��V�O�b-� m^�M#���R���(O�5zv�T
��4a%�SQ^$[� ˸g���jӤ�n�՟h�'?�$�'� 0����N�� �qJ޿�Q��G{*�|8��Q%�����`�50�5����R�ɇ�Mヽi��'��������! 6  ����T:T��N����0t��1�M+ �x��'8�_� ��	�	<Tt��e�"]R�hF�)��o��Q�"�"!Z�I5C��9@	�b�i<X6�%�d�|z+O�]ȵ��B⎔��� �h(�"��O���f��O�$�Or���\��D�O@�U{�v P�h�Lz�}�0��-J�`����x���`�i}z�ƿib����|�'��eR���F��h��=�N�ѳ�D	��F ��Z�UZ��ʜ,�m��(OԵ�$�'����bJ�V;~a+g��7:5"�d79�O���O��ʧێ=2 F��3|ƍHr��)]�����h��P�Py�=�d*�<.���#���y��˓G�|pZ�Z����C���mUzb4��lC���j�Pm�����O���Od��& �*`6��C7��[1 �L6-˞�A��٭C��܁D�R�R���U -�~eGyb��zζ`�Rk��A1�"�9=���z7�B�r���3 @�v����!9��HDy"슄�?�C�'����'b��.H� $��H (�:����8������������#�#�ItA۰�*"Fy
ד�?�i��6�r�L��/J>U� �3�-���*�O(��Fݦ�����O�P"��'�¼i��l��d�$� ��A�h.z�Y�i�i��H�o��@�ք�dˇ!�����HS�&�'�R[c\@��E�v;f���Z��]��4%	�L�P�҆[�.u��m�9yj��0� 3�>�>�F���e�3�ʁYF(G-F�7m��b"NӞ`n��`F��4I�����7C^h#ЋZ�$�m���?Q	ߓ�MsĊG;��(	"��!�d���	|�'��6��ͦ�&�`�S����)\5�D(��b��i�O�\��'�a{��Ǫ   ���������4�?���dF��TɺT��-Ee)�)p!��"��'�r�'n��I���)����D)Q�^b
`�'�ўp��4H�Ƙx��e��`;E� :@��@���O�O~"?���
   �nZ�����e�To�H]Z}(�JM�JG�U�v(��
���'�b�'���s,�o1��IFL�)}P��C�ϟ���e����5+��45d�pшD�s��
1��!��T�_}��Js�[�t�$��)3j��DTJV�0�G0Y~����(G�On%�r�'�T7-�Ȧ�	n��Z�+���`Ǐ>���BA3�	П�'��'Ȥ�B�n�fh����19>`�f���w�0�1%$� 1�ߎ6��Y�ɒ�v�c �#��%h��'�2���f�0���'�R�� ���c�M�:����&X)șڵF��.nd �uO^�y:,���3Lj��`��L���O���;l�v��E���(�2(iW�n�Yz�
�M�z�+C�E��uٕ�W>l��$����,�M[�� ւ��kHES���(�4�?��if�7m�O����Y����͸&���GH��p��F/�?�(O �=%?��jՏ�Jm���ʜ/E�TX�?�	(�M[Ǻi��'r�Ԩ��O���^�P4tp�"�M=*�j���^D`�͈ ���j���O����O��N������?�ߴAþ	�*�u��4.)aB��p�=Z����M)m7ح��ɷ&����]�d�,�?T��[@�cEA/GX��H�@��rU^<����VP$3�cGi�\�;'h��(�m8�	
V���V��~�Yb�Gz`6�
64r�Ӧ�&��I���$�Xq�m��Pc��[t�>m��'�O��"F�Ct#�=*�[5e�79`r!�%t�d�O�q2�Or�ɺl����4�MC5z�c�D�b-�a������`�B��'s��'fP�;��'�"�',D�:6 �'��1c�4ev:�����abO��h�.��t�K��M����#0�<��$�/u����k H��!U8�F�j�Fc�(ui�(F
kR1��z��eEy®_�?iƺim<��v(W�!.٪��W�v@˶Ag�$�Of��<�)��h�j�p�G(4������o�!�$��8�3��k���ҭ�r��4ta�FQ���3 ٳ����OBʧXDqb@��'
.X�$�Y�4Tfm@2nB��?!��?���2����b��+c�$�U;�mࡈ�?�uKVm�j)&��7^�6Q:�����'���;'�7j5p52&}ߦ�e�̺>}�\�3_9�4����fhqrg' $Db�����Ol���ڦ���=U�#"�E�Gh��J���J�.�������	�`���RS=<d-ے`�~����O�l�>�M��O� 2�O>^��QQ���,;U��<Ps��!��ßp�i>�A�F��I�@lr'�Hh0�ݶz�@e��	M0At�O2*݊D��=�8�xQ�BHNb�a(������y�I݀^]�Y��	�L���j�@^�
����CX�R�ƽb��yb -τ�H�����n�9��ڧ�
�rVÐ�7��5������?�ԾiJR6-�O����Y��aJ�dQ�₦O���!��?����$ʨ&nP�x�T�5i\0a�KϤ�qOfEmژ�M3M>��'�Rٴ	��l���P_��p�(�N.��O���D)  (��Tt�pQ��\c�P��&�ĐX�'N�=�Lpݴv�$��	2�M`T���"�禵�7 ��o��<	�|�P5K�����X���ց�k�����]	Gq���d/4�	⟠��4C�&�|r\?��)�N���@O�� �yˢ�S�?i��V�v�����m�ڟ`�I�|`Xw]b�i� : �Z� fxhJ )>Y�0y�G�7@��00�Ŵ�`t�i**��5!h$V0-��'��i�b'�D���gي|*XZoӯv #��F�O4H5�F�ϼ���T��M���|Bf�Ԑ���u6�̸�����<&�BNf���%����Ɵ\�'M��ʔD�Æ�k�+)([�D�#"O�� v�_.GxP��)V�XJ �jc�϶�MǸit�'���O;�I:{?��@v�ӛ.��q�X�G��=���9f&��Iڟd��ן���џ���O��;5��>����M�/g�0|��"R�")H��������$]'�`|�'jE
h�dEEyr���FF\:�nثkr� RC^� �$5���Y=E�9#���v1:��i��-t@IFyb'�$�?a��5�����>\�9���"V;h7�o�*���<9�����'�]S@��E��C�gU�6C!�� ��X����B@9��gr^�*wCHΟ8�ٴx���\�P�I4�M���?���V�� �U�����h<+pR�Y�`��f���	؟D��o�)ivʑa�h����=R�qF�R�����NR�d���g�; �|̰��%ʓmk���^]����ᘻ�|L��&�6z��AXt@)�X��τ��(OHlK��'�6�B��y�Iy�dW�_�����"�#A���8�M̗i�,�)��d� �	0vV�)`�	"f��P�d=��C�'�6MCЦQl��[\��a�ۂNn �I�i��>���'���'��'��O�i��  ��HJƧǉ)2<5���ޡS�^1bB=Sz �!ɺ+ܴr�ƹ�?	��B�?���k6%��D-�� C��,��3�'�6��릕�	By��'!�'�R�Y�-[�g�(1rF���@��$9,O@Qk�ɲ8�
��;�eZw��McN>Y"����*O|�2
����޴Hm��h �.J�j��J�|�µ�t�'%��'u*p���'WB�'���ց�j�1('Îh	jD�G��@���s�@۲݂�ʮER
aǌT#�(O����)������,�V �D.ep�2�v.P(��{�u{5@�3�(O�1Cb�'nn6�1$Ā�-��}��i1V�D,	{z��O�������?%?Q����M��#9Xdp��*��ȟ&���-���u���4O �heҷ�M¿i.�ɥkI4E�ڴ�?I����i� \�X� WIX�0��V�0j$���O���OJ��BJ�D��A�i�
	���)
]�S+TȺ�����`�!��o�~�@���o�vD�d���&\((rĉfz���	[��u-��8�Y6g^>ig:!!em6&#Z�0���I�[2NyӢa'>��OH�܃�	
�f�b]���
\Z����2����"|�'}�Ÿ%��g����B
�R,��x�����t���N����@�If2��
C�n�n,�D��5��?���|z�䕧�?����?��4C�`-�1�<^�n���O��>.l�K��+6�Y���s��H`��:C����"U>���1��.Z
i��+�/$U+SĔ�r|m��B�"2L�Ѥ��2*�	�6AT�8>�>ْ�wL-zs+ƹ|p<�ړ���
��D���Or��	�Q�I�IQ�>�trA�b��P:��pl�8m��@��'�a��źА�0U#�7'�%��"����܁۴2������O��t�i}�i�c�$/�~)���
z.j�����O�m;���*�"�D�O�$�OB	���?����MS��rC�r��Qx��ZE��e{0<���S>�Xx�a�b�	lZ�P�^�3 ��]�u�v��b1j����Di�e:�j�!��;�4dT�h���L)s6釓��'���R��!!�f��� ,2p�7,�%����V�I ٴ�?�/O
�$�dA�8��Z�oL&}sNp%�)X�Q�xD�t�
� �n� �%�4���lߓuN	m�l���M��'���?�N�.�  ��G�%�`���[�k��ND�]���8ƄU�FO ��d��4�,QJ�H�~Y�T�-ʓgm�'�V/?���c�j,�~���cݥ)V���6\�z�l_�*X��ug���(OdAZE�'�^7�\|�S�mcU/Q)M.�Ӕ�'YbA
�Ѷ�?)����'��% �JF3}���N�S@bEA�*k��nj��7-T?#<@r��5iM���eF �4��DX5R�i�''�T>)�t�����Iæe1W&Ʊ�X�9� �<~�h�h�#X�{1��Rଉ1jJL{EmKT=@����˱)�80(����~��QA��>xc���`
B+r�5�rHs�L�$���aw�a�F�9ջ��F�D��Z��\c��� 6g��.�3c�@g���4��t�ɇ�?iٴ�?q���i/��$�=!<Ȁ��,Z �0�'�R�' ~M4��rP"��_�K`�P�{��'��7����'?u���[����SJpɢ�#,�΅Jr��U�2�'�]�e�&N��'vr�'��םП�nZ6Os� �D��)+���9��"S���w����	�,'� y�
�S|d���M�LHӑ�J�I9e��؊go\E��ٛ��R&τ�h�� 9UƑ�1jF9��i�~�%��2���O�Xh�� K�8-�z����G!ğP�tN͟@��4Z�(�gy"�'���eJ����I:�ҽ:��/����+ғ�.�*�n	>>y�=���T�Q�
��qBu�2m_���?��|���)qf   ��Q�X��i)	��M��J9���^>!�S�C��E�zA8��4i�!z`�@��ʦ�!���facf;}���"Uq�dpZ@���6P"P�Z�����.�	�iY[�^�&�b���0��E�!c��t�h��e� ���!��Ix���l�3x���a%��TBh�]�V��<�"�i �7-5�D���݄R�`�VlX���JG�M�M>�ۓ��� �  @�?�� ��'�6m٦	�I9�M���2���Mӳ���b^z�1%��D�vHH�-P5=%r��>�z@"D�'���'��$}ݡ�����l�1��Л�e�%O-�U"�bY��ɦjA�����^c��a�1�Bl
�bu�g�"�y�P�_�<g �6�CŮԛ:���f�&FT ��f�纛f ˚w�>�Q��d�&S�Q���O���&�6�Vq"u.�̟���4[��V�'��I�l&��1 %.hf��g	�=pw�ڔ�/ʓİ<�@G+Q$Вu��SA��{R.۞pd7�"�� �$����<� � ��o��!(�"L�쀣�b�)~ P�X���ȟ��	��L蕧�ϟ���󟄛$��j
�9� ѕ}$�⋉-x�B̈�J۴Trp�Tņ�r ��	��h�<A��)fR�m������ !�A�r�i���:b��D�5hX7�[�װ�<qP��ٴo� � D�z%�B l�Ԭ�%kU��ɇ�>9��?9�J~�SU}ácȲ1�`�k�X�'x�?�!�^�-� ���Tض�����Gg�&`}�B�O��d�OȓO�7��&' �  �^���`��mqXe�R�JY��Y�oW8R�d���?����䓒HO�����  �}��K �D*g�f A�eK�2���GX�c�8[%lF�C-��+s��0/]F9b�i���0�!g��kG�V�y����j�ڃÏg�V��O����O4⟒�6=���y< �Kt�25��T���>aN>I���O,4QЫ�=O����!]�^�*-�7aڦы�4�?�u�i��M� l�����<����uㆸԘ�  B��B_�p���.�����y��Hg��X����) ��WhE�9}PL�����Ѣ����@V̄�{�޹���&LΨ��B�ȗEyȠ� �T�!"Ib�Iڻ��@�όQxLh`���,d�1"c��[�b����	*�M��im�D�+ 3�X@���/��A�I�[d@�4�i>=EzB�H	)m���gE�;V������p=)��in�6ͪ>I�͐u�ft�4$Z tPL�  ��$HJ�plǦHN��'n�O�u���'��'Λ�\�;;�ГD(fs�e#Qȅ N�Ȱa�$Y����U�ҭ"1P�0 BU�ʧ�
Rm�jT��5F*�mp�*X'P�L� *L�~p��Z�eZ�C�L�zVN�)=�H�CGg�,qY�O��݆_��A��Q=;�j�*���V��mH�p�F/�<馟~z˟�Ʌ�d����(�E�?-�5���şT���ė��ɁP��O" ӏ�$GY҅(դűs(*��������޴�?�V�i5���?eoڈk�,TP-�u�6��Q #��� rE������?i���?���z��n�O ��zӞX��?Lt�X��)��T���@n����Äǆ1���J�ǁ>�\�B�إx��xk�
@N\����=|�~�wkܮ�
�����M�����F���>6h�6��e<ur4��������(h!S�3F�@�s	eӾ�x��'$47mX���� ��i�	?ty�B`N?0���hP�ϬIm#=����~2�nD�Y���LƸ3E�(z��'#f6�3��릡��ty��L#�N7M}ӲhT V�VL���68��+K͟L�I���u(R͟������2�N�2f��U��F�VG\t挫?���T�~}���i�A&�P�tj��<QU��I��À���AD��6��Qh���BR�ְ{ ��q�lh�faZ�0+�U���d�
~�"�aӈcTlF+>
��8�
̸d���k���
�`���<������'"��0�AB�i2�#aY&CǦ� "O�r���;O����Bk������Q�K�ިsܴ��2��n�OΓO�6ɪO� �  ���sl�=X�f�:�׆b6�(8���؍�0|Z �.T�:dYKJ�e�<�*�ϝSܓO�t������DnξT�����Մyv�Q�e�G���	��X����t
�*e$qH����qLvy�u�9���
E���3���]���C��H�'`�aR%"96mS8|	�"2C�4SD�b�@�rq�,SFß�3�1O����e>�E��>"�z��Q�@*[���0��OV��U�O.�+���
��9�@@��""
�:4�E6e���ϓ�~B(�����?1z\��L�7F�4�w΄�sb7��xk�''&��3���Pt�r;+d��b�J_2IΓ)�´�R�>�i�	X)8�ʧm:{��Br�| Ŧ��$���ȓX�H���hN�SM�_�&܅ȓ3,>�k���jH���󏃋\�=��M�`�cp#\Q�I�f�>�q��S2��0�O/qd>�R�IEeа�ȓ }B1����b�C�4&lb��F�<�1"2�0��O� uІ�@�<���|�ܙ	ׅ�(y-�Q�DEd�<ɖ�U>{���2�F"��m�D��b�<A��� a�E���C�O0T�U�<��k%~�C3�G�~����N�<I�R#.sHu�I'�:�u/^I�<��c�jU�Q'	�6@lhQ�aGZ�<�/�m[�՛��/ ������_�<�7(�8.@��Q�,";�5��N�Q�<�@ܟ,�r�h&�O%|�p�J�ɘO�<�7�]�p`Ԋ� �|�Y2�l�L�<AU%GL��ŻŌ�4@�B��t(c�<q��"G�9�1��4{�����f_�<��U�i��)���7p8ADIY�<�����D�l���/@<�\�7��@�<y��֤ ��:F'J� ��U�N{�<� �@;��F+Kgr�H!͟ju���V"O&,2U$�5"��I��mt�e0�"O�-�3B�q>F��EhC�(d����"Of ����3��l�a�P,Sb�u� "O�3*�]���jS���vH��Õ"O(U@�Q�o���jӏ��u4���"O�H1��T�Y�.��ŀ6uEt�q"O�� ��H6�b�pQ��?0N�#�"OJ<`�A:#P�բ���~��"O�-�0!�70j(���9�R��"O���#�қd���0�B=|z4�a"O��D��m0u�r����\�`1"OP�AVN;��JiB�8ߘ�Q"O���Ɇ���`�g2kÀ�s�"OT)ْnôM|����E�?�U��"O�����,90���]�w"Od�W��e��Aȶ?f,���"O~dʖW�N�f0��A�MO8���"O��;�
��p�,t�ê]�[DN���"O��h$(�q]p�P�J��2(^-�"Or���`�u�6)BCd��F�hA"O�;��"�4K#"Q�4X��"O��'ꞷS˞8㶯�s���E%D�x:'ԵJ�~4b�HA�B�Ρ��B0D�$2g�c��|5$�]�Q���/D�����^���ak-Bq�����-D����OQ���XQ*�)t�l�2w*(D�2�k�6`1&�´��3u렼"D4D��*�M�1c~E���D�\32�>D�@H��RGNt��ć�>t�>D�$`��vL���3~jU o8D�l�f`^  �6E�FO�+D8D�A��5D�`��(µ8�a,�;-�`�Bj6D�pB�	�S�TM;c֕WT]+�5D����>hA�m���#$qA.4D�@ �j؇<jV)�*,�X5شB0D� �i�p̢\��)�.d�V�#�.D� '�W���1�M���Ʉ�7D��ڱ��q�Q��¿\B�bT�6D��qW�����EΟ�'�`�6D����Q&N\\	+���Q��8�(D��zeh�K7&�3egP�2Lr���$D�(:�(�0T��f��b�T�B��%D��[#ƈ"���H�[�׌��./D�|i�-B�{�x	�F�;S�LI9��2D�����(>Y %�J�44LNq�(0D��;�)��Оd�3�_�Q�:��`@;D�QbLwx��1a��(!��9D��� %Q2��i!F'MR��2�8D�0C'غe+8��*�j�PK6�!D��	F��=����6b<"�<(�(3D�PX�k�2���JR�5r�h+D�P��Z*�����F2<�V�q�)D��RE��"�p�h����"-�5�-D��X�L۩#9��iB�ۑ��0AbK-D�yӪ	�*�rt�çە"��e��C/D����.�*lX�hmSpMa2ȞR�<Q �f��t	�,��qP`�r�<�vI�QeV�)B���X���p�<��P�)@\݀��2�9TBl��D{J�26@�҇fP(G�D5��J��y�G�*�ZU�+�iΤ��� Ò�y2��<�b5(��\V�ؠѬ3�y��9|��kšPL,��A���y
� �YA���b9́���
��"O���c�ٴ%g�ĩ ��!򀔉�"O�9����)��%���4��B�"O�Hc(��0,@cV¶Y�����"OĐC��D��-�cm�d�L!��"O&�і�2��P��KTq�)g"O��sV�S�k4��؆��++m��"OtM($�^6W�J�� ��/.e�!"Oʭ��ŕ"K� �a�b���:2"O<�d�!P2�x�1�I&[S@�ڃ"O�hh��ߐu�f,�W/�;!N���a"O❀VBFQz�@����7I>$�t"Otdg.Y�g�rv�|E�4�&"O���PɃ��@�Ti�;.Zt��"O��0��	?w{�N��dL y!�"O�x��ս�Vd`��ĖH�,���"O����n��,��$�s��

����"O��(��Q?��ICA�A�(����"O�����Z6t�F@��Jǅ΀uK�"OFD"�����ʩDi��}�!�"O�4K�ƓT)�]�E�ɂ$.�r""Ol1��O�� ���xd���"O�����]�+?�xX%��om��"O��8�m��q�4��jE�C� �1"ODacJ�:�̍��Rm�$,�"O�Ȱb�LOΘ�A��8�N00T"O6�	��U+D���rEg�x���"O������(!%�@�*�Zp�"O8ѓE��Wr�I F@�f�64:p"O�M��K�0@zV%s�d�N�d"OF�bU�ױW]bx���6���C�"O�\b����,r�F�.���"O��� /���b�D;gФ1"O �+P��$:�у�o
��qa"O��8���0f䐻<��9�"O��1�B�
R���{�`��T:��"O4Iɦ�3	Ly;����S'$��#"O3��Ȣ7|4���L?]�uxT"O&P'�b�b�Jv�ɫ/TU�a"O�DQrH��]7�T�E"=t�b�"O�	S�OJ=ߍk'��7��P#9D��� �بuJKa#
' "����%:D�da�ʵKs�ġv9R|21B!j3D��x6#�GM�D�.H$*E×�/D�؁�C52�a�e#��IK�"/D���S��,;?�"邌=��#u�,D�(U�ۃ8�\-٠A�t~�rv�%D�\Cv�J9#C@=I�dD�������!D�,��j� E$Z��4�ë�+`�2D���AU�y���2���|\(��6D� ���M-đh��������4D��I�iY"�`��"(���rP�1D��ꁣ�r1:�*Ç'g�qCB-:D�|Ó����ĥZ�j�.[b��D8D�`hu���&]��DP��Nŉ"
+D���i�.���8���Yh\e
�A-D�x�!f g���.�8W��ё% D�,��Ő54qXf�@��|��w�?D�$��"	eW�I��w�lL3�*>D��B�ѡ/���\�N�����;D��26�ʝJ�8ɒ`�6WT5�8D��	���'��-���H�B"���	3D���r�+B{�Y�A<4�Ti>D�x���',.]6N^�E�tҰ;D�� ĉ�*L<
�Aj�΃�e��a	�"O��0�h�'!�:�z�L�6\�lyr"O��QV&ۗU�&�R���	qZP�{#"Od,"dk�>B�l��7�4iQ��"OL]{�ɏ�y���K�dZ�;>LH5"O�*e�
f��5�ˍM2Д:`"O|]���@�;s�Q�f��R"�5T"O�lӡ͔4e�����̦�d#�"O~����D<Aać��'"O<}ӱ��0���;3�Z<>��=2P"O摡�B_�<�-b�D�s����"OT�q��M�Dj���^h[�"O.Q�ѯՆ@ZE�vCˏb�c7"O&��g�¬��V�ǹ$���2�"Ol-�$���������[��d�T"O*�AKB����a��!jcX�Q�"O�����sy���I UR��br"O���K
�(�u��?hX~Q�"O^�2�J� SXr�1u�AT����"OB�A���J����G���>  �"O�X��,��*\�@R�V����"O��
S�G�D�H�Ѡ���@hY�"OT,#��7`����Ň�7O��	8"O�0��E��̸�"A�6�����"O\��Q$Ôt��%��k�)*�0&"O��p��8�83�*} ��Z5"O:�J�l��� �7ʍ�
t�yQ"OZm0B�P�)X��I�I�� �H �3"OUY��G6`4d�S�����Xy�"O4�0E�gfr1c6g#(�>��!"O�$
6M��+e�yS�_�S"O����S"%b������"O��SP�Z�x��)�O��:�G"Oµb�h�!Vm�i�Ѓ����0��"O��0%��h�z�"��f��8D��Yo�銔;H&/�.��$	#D����B�l-��B��@�
��]�h=D�L���Y��p�I`_4Q�9�9D���Ǧ]�H>z��7i
��T��D5D�᧠��~*rTA4d�4n�rT��,8D�ؙ��Y��(m�a�?� ��/;D��S̞���`���:j۾HHT�-D��)@Ҽ��C� @�Tg�,1ա+D��$�Y�c��+�`�|X���-D���v�*[\`��\7f�}cu-D��ċEt��9ƃ��/2fu��l�<G��)��L�����R��*ŏ�W�T�ɝ]����Ÿi����l����'�/Q@R��FJѿR�>��>(J|�V"[����r'Ş[���r���DH| @�Ǿ'��$P䯅�S4����gI\�'>NP�sC˧7�6���&c]Hݙ��"����Q!h��t��ϝ},�H��=�Oհ��'(�7�
X?�QV��I��K���'^?Y��?yN>Q��ɂ�G��U1�",&Zdu���҆'ҡ��̢��g�	�H6�QB��!v\��lϦ�'��O��M����?y,�����&�I#��	&����L�]솘�o۟��ɸHK"�������`p�)T>4�]w1�jqV?53A%ʔԹ��`ƀW_|�xRf:�$��9�n\;����_Kv����2-��L�LG�"�j�DF�h���a��Z'>�H0�UgA k���*%�Ô6f�o�	g�<�dئ��+O�D����܇�.�C@I��I�C ׸'���$0�$��8m	�gA�����Q
v�"8E{�OR�6-ܦ��I�Mk�4B���z���$)�lqc��%B��1�zӐ���<�����Z����>6������^�t`jud5ZX��q`aг$!j��	�HAHKua/Z��L�^00o�]��Y�V����":��j�Bέ������n�X��a˨\*���}��X�!��
�$&%ݺD��P���^��;شp����'�$|�������e��#w�ʃHY�����L�33*q��.O��XD{��IM50���uj�PSR1iq ��-��-���-fӀ�O����韴�S�? T�2��L[ҲHc�C�%`�V�F���SC������	�����u��'���'/��a�K����d�`e�+�^8�p*��Xs�G>&3��,Ȼ1���M��(Or5R����25��[	ܱS�C,� Q�P�[&z�`}�d3U��Q+��8+^㟐�ٝ<ْI��чe��}ʰ\���$D��QP���!�IYӬ9AN�A�	�NïZ�6T����?!g�i�OH�=��B�"�x �c�4y�nI�� �\���`Ӥ�$릉�ش���+�~�n�ʟ(o�
��$ѠE�k��թ��
{�(��?����?����?�С��aA���>{d�p�S�X��$M����c/qb�qK�4n�GyBf�'w�	+���CBr��M|`lA0�ʨz��x�˓�E�� �M��I�!,j��'�@���OT@oژJ��$�C�`Ye�d�B�*�	f��$�O ��;�)��$j�p��!��R��9"g�	"���<r�	џ�(��A&��)�
�<.��FP�
іqXݴ��$W��ftl�ǟl��L�/�c����[|��Z1#ƻWa੓$��W�b��O@�:� �*��ƌ��z��Rr	�`a�D�p�~���A�vp
C ��gF�B�P�ɰl�f0� �ʐ��0�'L�yH����O4<�B��O��=����5Y�!"�o�8IҥiI<QT���X�46+���'�����{w�R5[��a�] �(A���O�ʓ�HOvi��K��P��CL�r����'�T6_̦I&���׎/<x���BA�&����8l�\�������O,�Z�
�  �	!�dVC��G�	���˄MՋ|�!�d�"\���[Gϙm�x�[��[!�!�� ��{AO��F�"(;�\3@,+P"O��R&9f�p��+�B@���""O��2��!u	��2�� #r�i3"O���P�>T/ ���X�gZP�"O� �S��h~��'IٹMsb���"O��׼j��be�"l�U��"O���c�/U�x�؜b�$QY�"O�Y�,a�DSG�C#1��̹6"O��d#O?=0��>OD��"O4a�V��)�x�j�N�w4��q$"O�m��C�F�Pu�� ��^ :���"O,-��EJ�-��q����7"��Q�e"O�� �����`TjԺ<��Ѡ"Orq�g%J�e3�i��_��M�7"O�Q{$iB�jxXm;��'t�ƴ�F"O�=���قO��l��̬GgF��w"O����_B4�gG�!;X�!�R"OX� 2c	�EXn����ŝ.<���"O�$��	�|�Q�e�҄2�̓�"O�mk�Y�Q��T�C	��2Q"O*��# Vo�V'9ji��9g"O�`:U��>��*�Ł_����"O�`^(�QC��zI@x��	
!�*_�
��DN�iL�t���t !�Y�h�N�{�&�5Tu�t	��5A!�$��G�"ׅ��А2	݇�!�L�Ab,��@G֡I!"�#�đQ}!��I�-:�лp�ƾT&�*"�ʹc!�$C�Ec�D����-'>�&=DJ!����U��I�%C�C��Ie��T�!�Dٔt��@3C\�p�G�@�[!���7M�z,�poʒG�%���E�7�!�D]�o���ˣ�R�@�<Q:��1�!�PŐy�F-	�1��>f�!�$^<?�L3�ЕR��X���P�!�Ğ98L��I���/�n��0�Lg!��j\��5Z�N��M�.~!��"�^�kf����;�.�6zh!��+4��Z�g�z����6NV�v�!��Z% �ti����W�V�� �K�n�!���s8`����6�T��"��a~��'�ɑ�bV.���S�E�?I�ZM /��5ZEm�x���	 +i�d����m�����̢i-��bG��HH��mʑ|���+[Ov�@rI)��^� �k.[��Pb.	�JY����Z�J��3wm���4�Wc�0+�jaç�f�'���ߴI��Qĭ]>���f�;B���dEr�.�$��Iǟp'���O�P���j��CX�%�l��\M�dh�'�T��A@��UI�"�a�hM��Rݴij��W����$�M����?�ٴzvY�H��a�,����ޤj�V)t��' ��k�cd�S$�&8��V8*�Y��� *N^�Q�G߂,=zUBW�ǝ=�����)A.F���A��P��C�˕���1��ob9q`�7�b���)]�(������9��Z�j��m��X�����-O��Ю�Mx֭���f:�H�Oo��	����?E�D-6n��g'(m*T��%?*��OX�=ͧٛ���z���XW�M�=R l��J��
���7�'��6��XXD�m�����'W���O��IG��q�M^�D���9�cUi�~�y���4	�g�CL���p���8#�S�~�`�Ͽ��� �2��(�08�=�e/�t}��Y-TfJA�7�ߴI�N)8�	X�����G�S���5���M!�Fu[���ib�o:��ɍ�Ms�i52��56V��F��	�@A�&��R��'$��'ў�'j���s�E�[�H��V�3ℙE}��|Ӓ9o�z�ɡy�aY��
s���9��#h"�޴�?!��?ѐ�J�x���?���?y�����Q�J:�^e���Y�q�%I�0�H�0k[&/F�R�阉w���쟰�2�ظx��=��=Q7H�j�`�����h���OӛB��!�կN�6��y���,�	S�D�a���&�Q�B�p����D�l�(%'W ��ɖA���Iܦm�����9y���Q$4��iDh%���Vb��?A(O��$�O޸&>���5áI��<=�2�A�&7U���챟`1�4b���'I�7��|:����IN� �-3�o�`��9��B��$FhEYAhQ��Y�I��|�IПTsXwZ��'>�ͺ��l���U�F��8�Iz�F�`E�>�!�w�Q7��� ��V�h\��̾�L����Жi�6쀅Z��P�-�Ge���f�U��X��	̑r��Ə����,yK<����C��N�Z��%� ��8X1�1ƛ��a��O���3���|�U�H�y��y[�L�G���P��xb�	v�'/���ऋ �����*�4��ORumڡ�M�-O����\զ�	�0n�0!����؞)h�)�`шX��q�������?��0rj0��i�2�Y�"S�Z�B�d����頢,ׅ�dܘwC��V�@(�CLU�'����S�ۍ>��`	tF2m����"k��O�F�9��IJ_F��s��?A��l�cp~b�0 �O��(��7��O�ם+q��ӤO�{m���E:F����l�?�|R�OZ���R�l!�B�?�Vi{C�'%�6���k��I�Fʌ `=��P���wpT�*O��F�sf���9�I �D�v� �  ���͈�	
�Cі�*��	X0d��;�Ld�+�UXJ\�>��U��Nc�4�� �7R5b8���U�N-�3���F�Ħ<Q�����P�ʑ�S(T���	"�ś4�luON(��R�_Z���7w e �Ċ-�*�x�4��[�.�OȓOj6M��9^ �  ���
  �y#���	>X"��׺i���uA���X��E�8v8>�%H^5nd�O�S��U�S&�dY��ig� �W$E5��mӂ�Ez���U�2�n�9}�V�9t�yiZ!�	⟨�ߴ��'���$ٵ��,�hPB�;M1���J�?As�i^r�j�(-n�H����J	�6��O�7� c��� H�~�`u��� >������X�WԟD�����b�FQ�:x�!�L��2�,1�6�����&>�f5�����c��dk�i�/��<y�ӻ��������s�"���.xj1�ef�L��0�K�h�G����
���d�On���'I�6M�/�yү��q��̣�%1b���GA��~��'����i�_���Y�X�t�j0��d�Q��#��D�O���lXU���0��C~���Nғʚ�m�@yR�8d܎6��O��d�|��ӱ�M[�%߇w�\���dw
>�hEDG�eWr�'[`P�gM�w$�8%#[@�\3��w~�8VT?���s�����O:POr�sv+�D�O�@|����D�P4j��$	�Qp��G�LΜ�̧؞5��OW�!s��B��
뤡%���ce�O
@o���M����OනY)R/� !Qc)��tT[�{��'*��`�'*��ҐJK7\2BL@�D��4*d}jǓRěVb`�JO^�#!n:f�,Y� �W����v�6�F��Iq�	z�'��	�� ����
��eO�'p��T�Wޟ�� 	�ٟL�	ȟ����;�P��vɎ=pw=�WE�MѶÏ3f�QrM�[���!��Q�YT �<�#��T<6�P3J^�K�}P�	]�o=���B�Y!�� K�?J�>������!,D-'s�O�m��'�6V��)�.�̈q�����e���}3���՟�?E�$
	0v"�w	�_�@���'��"=�e�v,}Ӭ�[t��1�P䀗s46Ѐ�<�@��$V���'b�[>-R&�ş@m�_�hU�pd08�h4�1#-1� `��������+GZa;@K�T���*��0ᶌ�)��ם86���r�L)O8D�N�0y���j
����'N�D�Zr���H3>�	�@X<4~�J�?�9��K�R���!��bR���À�>����柬�ڴ{(�F�'�>����z��qh&��~R~���:}�'��	Y��Z`d�k9��Ѷ��#o
Qqe�u�'��6�G�%�`��n9v�tin4Ar�L[pk��7���t�	tX� ��� 	  � �2�Bɷ*�pT(�8h��2�I�O����ʦ]k���y\i��8ny���֩�1r�j��?Q��?����O�PY����il\d��瑊���
Fa�TX�<ܴ&:������*U���@�=ڠ
v�
?=��R��0G�6��Op�$�O`��%v�d�O��t��PA1"��R�,���N�Q����� @"�K�ML�-:�!F�4iPĀ���o��O�z��;���{�,iD� ہ
�+h̥���6@��B
))�L���B�H�뎓)i0x��[?�*�w��rRE�G�m�R��%R:��r���OD�oZ0mZ��,��"|���� �|LY );L��Bb��A��������c�^X4\T(����\��@R� !���?�v�i��6M �D���i��`�'�`��ӉK*j�{k�џ�CW�_���	�������Y[w#R�'Y�vE���#�M��{:)`�↶)#���W�]�E�(d%�
A�h�qe�K�0"�����5��13��
k�ӲJX���b�ޠ}��q�� %-9~Ȁķ�R���.�&D\~��<y����ᖣS�+嶴)&�l�=pci�%�?�s�iݒ6��O���?�O<q��Ӽ1�<#�/^�x�l�E�'zay�e��V�j$0��\jTެ�6DE2[�l�L��2h>����ny��'�1̻9
�� @�?GF1�O��&iPw^v<J�o�O�.���I;f��iBda������St���2Rr2� �U�}��Ha��yr&L|9�}��S�u�>lP+�9�?ɧ�X�$�*99��H����	�#?8(L�`r���,ʼSXC�I4�pE���o���Dǯ4�T�aSN�O
�ۆA�+ZE`�c��|Fy2N!f�&M��B 9?G ؛�l �0?Y���!*x��@]���c��$���f'�����- �O�H�U��53W$�F��=rt������J%=ŀܢW�~j!B�:�x��d��)@��!PF]�<���şM��g�ҥ<`j])��g?aB���A�KW�XT�앧h�THS�\,U��ad��;te[T"O�<�N
;9�6Ṑ��+��`B').}ba�	V	��٤2��d�
\OjUi'n?�<���Q�|�!�D�
]M|���
^''RZ� Ȍ�� 8��	�Px�G�<�2i�oD2B\�%j5���y���� g�)!�E<DE��y���1�y
� ������ .:��BR�3�����"OҴa�`аj��'ܼ���p�"O�MCG�	�UAbaco�^��A2�"O���
|hh�֩�#�`aB�"O�م��cD<�H���Mo$��B"Od�3 Oʾ+欙#�H !C��""O��Q�Akr���Q2ZȩW"Od�����2* �$���_�$�94"O��� ʡ%�ZT�bҖ"<@AP#"O`��v�/n�q�!$�$O8��F"Ob��#M:<& �z�d
(9��,�"OPaW[-4�P��̩.*��"OHsӂ�/M�$� ȝ#���#�"OJ	g7u�@���g�/S�"O.�XC닾%ђ�&��1���c`"OdL�Q��*z 8Ղ7��'.Й��"OP�S�h �$W�H22��2BZ�ʖ"O��#�M�=#��bm��$z]�"OL@;�i�SX�Q��!��M��"O$�c�fk��Y��M�&��Y�"O�Y�IX�j�,*��ِy�l�"U"Ox�3����Z�x@�8	j1ٶ"O�Z5ǒj-�hF D{��]�"O���V���u�H�7/ޖ(��Ir�"O.�;����\���.0�R]3 "OLP[Eb�,��@�/�c��)�"ON�3�N�G�5INJ�I��� �"O�H2!��N ��#���Ybrq�`"ON��H�����aĝo����"O�!��G�%��E#�kτ���C"O����� `�����	�&��)��"OrRf�̞=�<�T��X��A; "Ohm	�dBn�(��A��n�zY:d"O�(�dI�8�f0��$p͊�h�"O�	ĥ�sd�8 ��"O��[��&F�`�)5,� }�(�"O^-��HN�?��xRc�ڶ��r�"Od\
Oŉ<�\PH��0Z�b�"O�hJ֮�	O>�m��	�gB�q�u"OJQ׌�,=���y���	ySԀ��"O��D��td2�c���zU\��"O���CfE-@������QV��`[&"O��RD*�b�*c�[�%�2���"O}���R&H���l��\��F"O�tcA�$�RQ��a�+��#"OX����C�p��Y!��is�U��"Ov�'�@�o��@���Ƈm$�@�"OtX�e`��0pj�`�M�"a�X���"O��;���=R�J����?��]�b"O�u�` :s����&�Ř3����!"O��d�@<+�F9A'퓣����"O<4 ��L�ưiq�I�n�z�Rt"O�i!�D�ZG4Rs���Z���"O p�BcR!H�����f�$lY"O$)%�٣N���dVi�њ�"O�,�A�DD<LI� (]BUꨳE"O
�A�D<����(�6TY�ػD"O 	*Rl�`��9pe�έ ���"O��D/�� qЈ�R:�"Oru��M��=:�`I<n�P�"O�H��Ս8#!'o�5_aX�I�"O�A�T)�3�*@�v�`g�%cE"Od�A�-ݠp�L4;���w�e�"O���$�9syPu��$ݳ����"O� � 	���{=T�c2�Lu��"O�5Q���2Xi�	�bW8'ޔ��'��$�qOb���Y�8����P�y,U�H!n�{�c<D���+�A���W����z�#���?y��u3dHIx��(:I�ȕ:vΙ��r�8��0<Oʝ.Y?�x�0�O�P2b)ϐ��PC6�φ���"O� �d	n6<�r�d�<v�2(zv�|��=r�& :�p�O04e�1FN3�q�l�,A����'	B��`�}r�D1�Y�n�콡V�Ź|��'��+���>��"�8r�-uuh��&Suh<�]\~p	�삗���(�޸�V$�[SfX1��"�O����07ʃ�w�|��-<O"u��A��}�h�O���E�P2N��eaBm��t84D�V"O��y7o�1<΀c�0�P$�|2�	4�xRDc�\�O�b�0"�4n)P���H)7@�œ�'�J��\�0�m1�-�Y��8IR�I-vk��'��A���>Q%mѯv,�c�
�OfB,AԾ��ȓ���JGa�0r���GF	i&(�q�J+v +�8^�V�^�.��|c�/�'o�M��00��Ԙ����	�h}d��uҘ�΄�(:D������~e�n�S�*��։�yR�V5ณ�)ՉJ��k�#݈O���ꆜ�(��������l��v(�R=��I�'<�A�DG[�+o `�� ͉�
��Hv�A����6��S�O��@��@ES�������p���"O�E�ѯ� X�8T�D�3F����Y��j�a�,#�%e�'܈L{&�	�Z~���1OL�*��=��u
���j�F%PcX$-�0Z��[�G�Hx��-44�p��Q?0�cEշT.�0�7ғ�
%إ�O*��?i�l.],ѫ`#
�аI2D��2#�YM�����k\X��#�qӠ)##��'l�AL�"~nڎR��Z���=<p�1�f�$utC�	7|D���L6%�.��6�����`����]7
s*��? �� ���I�q���P��%�E��MV<,���A��@iX�xs��U�d0�"ŀ.8f�k`mr4�RゞV+�#�:Ӽ 1��-1*��S�O�8�`A♶;4�ᐃ��}��Ҍ�ԧE�x�@Q����O�LQ0ā:p{�\�� э/�fY��K��?	��H�:�����DA�!�ߝ*�&C>d|���Cdp� X�q�X����j:Vm��L�J��i�&(�zcj�(H����X8)|:�p���#���1d�-[����җ|"$��Y��c?7-
x� %S�+26pV��E� (�����%��9[s�E>_1 �����}�8�˚�3{L��5�'
��6ip�A7y�ȉItc�}��d�8��$��"�hOn���[o�"Dj� [���r�̜ \x�%E�$�UJ�/A��!���Ad�����Y����>S$�#a�`-zSdA�:���e%n��I�Dm�<��g��g��H��$"���S>�Q��tU�L8d�H(DD�	�gg
p+���F8��rP`�V4��Ot(i�w'�q#hbuF��%����!�,O��!UC���
xS��3��h�]jq J�،��F	���!U&!���m�Mc�e9D]�fV�'�̤��Ɖy��d�p��6-�`���#�(���Br��$
�nʓA�~�kҊ,�,ē����h� JG=�?ɚwXH݊�KԨJ��������d�:�'�LIJ�4y��DR�˨^�:48#C�0?�bY� oO��3#B�5>��C�֤K�Hڦd +�~�؞��$H[�����p�6X̬�D���%0�B�c�H�D�f�y`P�7��S=�0.R��ÆOIU�8rr�F�Ge��*OV]c��I��clK>��[J�4:�7����CL8l�8���@8>8u��V�����? F��Є��Z>��I�iv�E��d'v�I�ol� A`dm��
Ӗ�O?7��V26�ёiT�^���0&.H�G��iM��!�
6���(������d�8sQ�-(���y���L����>O��"�'��Mq���RkΜ@�M�5n�нh�36|z�;����ks���eh��$��v�QVS,�n���l�?oN�h�"Oޝ��%ɸXoLP��U ~eڼi�(i\����>q�&1�gy�H"5t*�J�%��QtX}{6��,�y�J	�K��K��%jB3u%
�����jQ�Q�T]A
�bf�X��LZ�%Y�n�"?�h@���hNB�{d�ι��p�< s�X�~$��Z��@�4�� �Lx���%LO����O�xbp:�I�h �mI��d�ή���l���OŲ��,M�~�2��T�3��s�%��=�O� ̀ ���7[����&�X��5IF���a��>y�L����+�����ܼcQ*F�~Ep�Yf��H7%F��a�<��dС%��h!�\; ~��J�e�
I:b)�s�إ#��>	4R(�ؑ{O~
�˓�� �	�J
�vAdt�����p=��ݑ"HI|�<�a�P-@Q="�W/<��L�<y�h�Xm�|�TD:,O�1�1kO�ƴ��K!
�:����B�L�����&�S&L������8���H�>qa&m
G�(�*D�O��%��4�����U� ��r�#L�^0���=�aH-c����5}�3���R��.V8$�R�#���"O4�p�������:S��#,�H�1r�'z T���7s�4�O?�a�����r�	j�m��\�'qB��"�Y�U�.-��K�JЀ�&�t�'A*���UA�X���[Ȫ4��0�V�Q�/b(�Y�0�Q�j���S�Sc"	�`@�-�����%�tr� �腊i�Q�Ɠs9`����U	2`d*�C.8�^q;�C�[�Z� Ơv6��s�Uw���O����BU�} &[��	K�^0�ӓ ��h��a-��BU�וW�ʴH�oK����IS���J�:U(�K<�*A�={pb��֝����\��ځ��k�+��BԨа ,��|���&y2>�!��1�ؑ��i@�<I��nn&S�E�#��ْ��q��p��Ƃ1 -@Dkr�-���O؍���;P�䉨'�.���X�O��Sdh׫I��(��L��SF�n��T���#(r	�����>������!z L�yT�9*�d�����~~�yr'�8/�z��r�|x�4�����P��S兄\���C� ̰B>p[�O�H�J��>���R���P)���|r�R��H��M	� �X��C�Q�)T1�����+��>��,0�B�8����"OZtPU�JOH�r�cܑ�H�V��QC�|�����<�q��lO��x���)%t'ʱ8f@�)P����Ɠ3�n�8��}U���#%p�*$��IV
 ���w��;Y7�",O�P��)�c�OA�5�$��'`�!�� ΛE�	-9���R� �x5޽z嫏?)�8C䉔b?$�󡞨^k�R��^$m��㞬�Bo6W�a��'Z8�V�cak�6�Yy���,�y�j��yf
]9a�4QW@P32G���y��\�&�r��S2ICFq����y��V>2�cS�M?8�X��±�y����G��U5�T�gmD	�o��yR�
On��aʂ�b�jYX� �)�yD�V8<|Q�뚈e|`)АN���y�_��9j�*�3�P�'���yBH*O�l��C`�:]�v���yr��?#�3�� oŔA�F(�yRk�����p�֭]H쐠����y�!�-"=��jE�T�$<�	��yRFδ2��Cq&�yBz=w�P1�y�ʹ O"̫�Kդy�nt�F��,�y�s�}����pdc�-1�!�� �F 0$��6zS��P�A&{�	��Ei�Ñ��S�O�Fy�rᓣ8� ����2�R���'Yp��P��71: 8@�} ���E7? �@��JF���}NL�'��`y�H��Ȟ���!�̰?�i]�QH��2DnXLvF,���_3w:B�K�Θ�F�م�ɑx?��y�G�?(QCD��b�#?��2Ɓ��ic�ӯ3�65
�H9 �R�aBiC<[]>B��1.H�I3�k�?w�J��D�Y�^�\t����<P-���H����[�i��)��j[�]�0�D"O�E��(�g�"�˂�g�|L���D~2�WB������1��$+V�H|KW&
X���w��i���تU����앬=	����g�4.�Ld����Z��$��`l:q��1�|�A�W���4��OC0c�D�p��/�iF�S�b�T��D�'D����BO wE>PaM�����3�&T�h"6��@FR����7�2xat"OtB��C�bp01@=T�,@q�"O� 2���@����/�)"��
U"OFX���D�u��� �.��,r��"Ot��؛
*��� ,Y(x`P�"O؁���@�Τ�D��Zf�0�e"O����E�`޼���wed4��"OL�0"l��O̸ܲ��8({dT��"OܽY�l�%dP�Q���n� �2"On5zeL!>�̪g&J8Y8X}zg"O��v�D;N� 2�
;B��A[""O�|�hF>oj���"�tmA%"O�q��</�L����[��qX""OXI{�@0u$��0�b�8͒"O�RW!�w��
�hY�PL��"O$e+�遰*AF�b�&@�R�X)�"Ol1��*�9m��E{v�8X8���"O���V�?Qt�<ã�ޑZ*�p	"O�#��G�$��肀��py�3�"O�z�ʅ�D��Ti�j"I�!"O<|z�h�>�!�����3g"�@"O���M� �DȲ@'�uM���"Od���ʭg��&��<�B��f"Oe��%f�B	�`�#�V�X�"O�\y�Iߦ�ZUP O>)E΁��"O� (���� EnԀ��]�f"O�)2�E0���!���k3,Ls�"O*0k1/
�8�Y��#�"Q%F��3"O�IڲB�M�����NT$�YB"On:�OH�H���5!(5a�"O���`��A�9y\����"�PpVJɑDp����U�<�1�M�g��^���ú��T?)t�d�"�vS�dhGG�/ �H�RW�H��]��a��C��z�����4+j��'ɣj>V��M[� E�qIQ��ӟ�Ɓ�Gk�!�~��fɉ%mk�����u�ɇn��\�.O�>�p��
Rm��$�I;�Ь?5�:�qЎ�T��06a2?E���׃w=�""��J.��	1�����CEf���9����w;�@c`��!%n�)�� 8n�LC�CI���$O�@q�����O�&�S�!N�X�!*��/�V�3�O$PKD*I�_���w�O��5;pNH$\����QBN�S�:�)�'曖�5H��a�'*�a�e�� DlA��� /"������D<O6%�@lN�I/�����B~|�K3�a}`�?h�$�O���|D�B���z�ɉP�K��y�᧟�Kl���S	!�U2Q����E�ա�
* �����l���ty
�'Y��ԩٺU�,(��L?< �Ul�A���S-O�0��O$�E��� ���R�A�l �	SB4A�	����p,�&�f*U�rN!����А[4D�<1�Hvx�KSN�P>���l��ID,G,��A���p�$���D�p0�r]))#~2S	E O�2�B$h�1@�Фf�L���tS�D��=9 #��Mk�T����X>t�Q- 24|��/S�,�꧅0@��
2c��8��:�-~[���i�P�� ��I�CU�`��J(Ĥ�*I�P���1DM6Y�<���?9�bw�9j	��5�ԓsp�r�
M�v6B��� @�[�L91� W�w��PD��҂>&$�g� |CN�0�'�29�(��C�}'	�'�ČSx�(���O�8c�zg��x��^:a�̥���0d��g&��u�_>��e�5@.�a���b "��!"R,YQ�Y�'��Ύ�ɧ�O֘P��DEk�)#0��Hh��C,O
������S� �OQ>��S�|Uj��f�>���n4cx!�6>�qa�o�+�l)YD�Fb!���%�ʥ��-�9�lh��}�!򄙇8&��z�*٢^ƌ��A(E!򤇞!�d��g+�C�(uȑ?!�d�f��p�D$�A��,�&+Y��!�^WfY
ph����� "��>5|!�Էk��� �4�R�#�M�<r!�D
�
� �굀�4��@��8v�!򤊓�Zq�0!E�L7�d��V@B!�$�l���A4ʑص"�)P#!�� Ty!ԁ^�x�x�@A�z'0q�b"OND0��ԇ9J��w!L�`	6\�4"O��f��?e�:��/�P����"O�E�Pc_��$������$i�6"O\�r��^
f!�덥`�:�j�"O�!�B^1�L�X�($d���"O����G�0Bv�$%�1���X�"O,t�F�0�k4�%�¤Q"O���L��?����3"S1",��"OzY��!F���@	�bj,��"O�aȂ�J�7[0e�v���(l�ٺ�"O�cSK�-o�Dċ'�qL��%"OZ���V�5��Mb$H�9�|X�%"OBs�͡���Q�'��f�r���"O�E��ΐ�3�,�z��_QM:=Ys"O^8���n���Vc� "\�p"OjԳ�� =s��b�GW4|�f��a"O��p	��0 y�4ƛ'o�⸘�"OV�hbD1���E�� �H�`�"O *�FЌy����%��!��#�"O,�I�蒫/4 �¤_*\� "O�����~�@(�G��%��	�"OtD9�� <�� �C]�	`��R"O�E2���$(Wl��%%K�"O�,(��	+{2�IBN7B-��h�"O��e�K�6������K!^}��"Or�;RM] K>$`C �4#};�"O��Q��ҡ�j`za 7� ��"O�	hU䎭�<��7/A�^(P"O�`07$.ۅ���(x�2�� �!�ѝ~<�jK�M�����m��!�[�W�Td2��t��I����"�!���U��=��
���`�J6U�!�ę �3ŨA�3|��9 � �!��4c�f�:c�<q�����Y�y�!��n��V �Yd	@�$�+:�!�d�[0Tp��?�VܺFc�Ry!�$��B�S$�,H��,���{9!򤄬q"�RR�V^�X����ɀE!��_I�vts\�v,���:[
!�Ć�U�~�9��0���Zveă'�!�D��Wդы�nتeLH����%f!�\�<����će����5d!򤞔o hXX�"�K'��20mU?C�!��-��X���h&Ɲk���9�!򤏑H#�����b���M�Ne!��Z*(���Ò.Ԃl_ܴ;� #S!�$X�/-8����E@be�!H��8!�D�1_Tx��"���T���3T�ŀ!�ą"�fY��nܤ�N�ZCk]��!��
�I���G�5+n>|`L�pp!�d��ne�I� /�.5d�X��.I�!�$�F�� ��dC:^�Q�cТr�!��ȣL�4��Љ��)ox�s1�Ng�!�$pˀ@��ĕ<PK,�Ys*�{!��ߺ ��h�dȫ��i����yv!�$�'N��@gG,e�\����^�tk!�Q�����G�o��%	!g� _�!���{�l�KǥK�u �G�s�!�ċ��hAb��&x���#f��!��"~1���k��e�ծ�v�!�$Ȃu���8�`R
wn(�.2l�!�ĝ(5T�QD$H�ŢʥF|!�Dܝ*s&��Ə�dg�Ab��yT!�� 8��D�&8��\����X���"O��y�H��:Z@�CD�~�V�
E"OV�)Tb�a��\�?x�*6"O�����S�dM�"L�
p0�1�"O�i��a�ipx���ߥmZJ�Ab"O"��3C�"yu(-���i  ���"OL��A�n�Q���ɼP1zP"O���-�7˔�+`LA�	Yb��"O2�KVGB�r��<qKÎ.r���G"O�("�Đ�[8�A���K#rʔ��"O�)rDq�,���%޿@m�B�"Ob�����nCxx2��J�mF�P3"O�5����36��	�%Y]���"O�es�"xB���߃ ����"Ot��AMו/�L� �"ʾ'$ˑ"O$��DEL5T��|j��9T���"O�U��ċ4,&���Lۓ|H�q"O�t�bL�𕨕aX�phD�V"O*��aiҜ~FF�b���VT&�`�"O~��c��*3���Ȧ�A�rv"O@�j��ǖa�ʌ��׉X�P� "O��`��_��ɡ��ʒY
� T"O&5A�Ñ{1ru� A<+VɊ�"O�Ł�c�.����a�A��b�"OR��.�4Z_����`E�y82�"O�$r�A�11@�����3n���X7"Oعa3
��PW\a�a�D��H�9�"O:� �K�s�P���LS�-�SS"O�}���!����	�R"O,�Q6���j+2)+�B�*Z$�e"O�� $0C�Hԩ!'I.K��S6"O�����;vn:t��
1 V��G"O�|���ԚG��k���]�Q�"O�q��j��I����tJ�x�&��p"O(L ��4��XK�dC�玁9B"O�ts�X0
�\R�$�6N�ҍY$"O�tr�GΆ!�x��@�zܖiS'"O�pā�'�<��D  o%B�s�"O�J傽}	��T�X�)�W"O�0���#>$����&c��Y$"O�
$�΋%\\ ���0'6�L�'"O�=��^0w����H�~]"OLN*H�!�: �����"OL4�"���AB���paLU��"O����JF�iJ$�'9:�H��"OvIC�A�pT��� ��k��I`P"O"4��P�;�����`X�o��E;`"O|)����UA@8c�o߰ˠ�u"O|J��&nӜ	f._#�腀�"O�1q ������/�`G�lӴ"O�ycU��:*,P)S��)3��[�"Oԍ���G=.f����3�UY "Ov�i���6a��q��O�X(v�@�"O
Xqw��9zMQ�B: 68xU"O\ؚw��b�h�ꋣp*��[F"O����39g��"�)�F�x�y�"O�|"b�Ӝ�՘P�[�Orlt�t"O޽pw�QD�Dk�D��A��C6"O���eB5���c�D�\���W"O 	��ѯC ���G��B���"O0�R���7��1Po�?h�F��'"O�U3o
e����_�.�j�p"O9����*36�8c����8RG"OF��E�@6/`*� 7|��AF"O� �TS�OЁ8mz��b)W�e�<�"O��#�-��K��8{�摈M� ��"O��G��6��@�s�ب��8�"O�9��.fd���OJ�p��5"O|�1��~|���7��9c�>�x1"O����ҕv�r�w��*A��1�"O@�!���ƅ3��I"O*8J��9�BظP&��R�~3U"O��a҈�U�D�S�	��bD��"O�@��!X���Yv��#j�,yP�"O
`����@HfU�&��"4�^T&"O\���H��CL4��w��A�xY� "O~�"�ӢD{�=K��R�2g)rc"O�aS`٠(��S.�9Qx�	�"O�	���� �0T��ҌBP��iS*O���̅p���N��f±��'���"���x�\�S���QƠA�'���31I�SŤ(Y,��:(�'}zm����vt���e��:ԑ��'X�qT�!q�{�+��~}��'�>5�N,J�P���*��{�Q(�'O��GMbX+�|	�'�6��a��5Z�$��O˸��'lxurу�&c�1��IOJ��r�'�qt��u�H�4�@�JQ8��'N^�h��Uu��X���9@�1Y�'�"Y�� "�>�R��iZ8���"O������l�V��o�s�$��"O6TBニ%<P=��͚���b�"O�AXV�B�	5��1뚙p�^��"O����O.���?���"O�yH�MƲ��M����|�Ҁ
s"O��Z��G�M�t��F��_����"O�\ SlXW|�SKڦ��x+"O�"��n���ʖ�nD�V"O��Vb���jE�4�7a�-��"ODAҫQ4H,F9C��A�FL�t3�"OH4��]@j��D�"��$��"Ov8�ҮW�9+�q�gn��/�ZA� "OD�ᠩ�p��̠�'@�Q�����"O��%���bq�@fX���""O�\
d}�x2ф�I�0�i�"O��B�L�n�&d^la{�"O��#�]5AYI�3��VXyY�"O��'��L�^��Ç� Q\��#@"O��#�ʚ
f�b0i��^�T"O@�h�C�mE����PC,!d"O*�#'eP�`�QA�˴:���*�"O e���2�`��nZ����"OrT�u��x�,ѕ���G���Z�"O�Q6)�?�z-�TkL�	���A�"Oq�tk�l3-H%нL/��3"OvL�a�T<k^�Bp�
z(�e�"O�t �5<�F��tЅ/���"O�	���(E��� �*��Q��"O]bBF�o$����3��q��'`ԈA�M��R���ѝ;��!�
�'@Hq��"��ް!��7^j=�	�'�>��  ����	/5��8�r*:%���>��'�\����%rH|ʉ���A�X�ۃb�*z:�sciĺ���?�J>����?�+O�j�F�kݘ�ZP���~�bı$Ko�';���e�p���ئ5�	:JֱC�Xž %!B�&�(٨�4�?�(O��8������O���<i�LԊv( 	���.�n���P
��- �$�;ZJ��e��d@kQW>�j��c_�+R���`['UV�b��6wH<uy��ۡoEtq �0#��z��t�˰���L?hH���DC&$��hѣx��6��ey�`�?�����?Y�	(dig�#����g[��T��J>���IC�8��3�&
��e�@NIC��>�M��i��'��4�O��	�-X&��p@�
3�� �G8�!�f#H�M3���?a����d�|j�O���@�	b��ha�V�F�bq�i0.d^�ca�0��j$�'%�`� Z���=q���8rɂa¢O?R�]��՛P��E*�
U>9:�ۊ��ʼkxj�7N���7�Y�_!�?9��i�V#=���d�&Y8���6e��z���r U3V��|B�'E��im(�pF 5y�đ�Rs*Y`�'�6��Ot%m��M#.��QҦ����<�#dU8zn���,��5�>�+�������'���'��IĄl��t������E�q�b��� V ��ީ^�<�:��<I/.:��'��MK�X0v����1 H�x�T�"7�Ԓfo��h��@�]�|������DƖZ���bӈ��'#R�[S��d6J�c�k�%t8t(L>���D+��xm�,x���P�*1��&@�����Ǧ��JZ
k���ʧ�}S��22$J&�M�-O����n�Ѧa�IKyRS>U�	�cr��K�|a�M���;T����	�R%��)�:r��V$Qa�������f�;��Y+I���&M^-:ׄ@�b��xjP���lTp��!A��F�L��&鍫�Bc>�*��΀=p�c3�Y�_ߒ�:��8?��f���h�O�gĄv�����[�f0�K_)2�!���X�n%@�Z;T���L�.%�џ�@���E�Tlj� *��S
����1<��'��,�~��Iߟ��I؟��'m���!��iCL�8FO�'fHIBǄ�9�m��"Y��$ҲG�1����`ɋ�~�nPx�x��MI�Fk��q���-�FũT�"G�����N?A����c')(H����C_�4�kBiř6���'r�	2mb�d�O��=��HIƅi���F�fH+�G҄�yҤ� b�a��L3pF�4/ݵ����P����'��	�2O>x��ˣS��ԫ�Ǽ/���Y���{�������	ޟh�Xw�2�'��	߄5���ӰF�1��O�'&YT)�1�I��YPm�<�,�SBՊ��O��a��Q(Y*2a�/RR��h6Ą�SL�5�T��K����Ř`"��?!�L=0���4�V>${H�O��$�	�4�	s���rU��.(Z����4 ,P��"O$dZ���2��@�>X��*T�|kd�,���<QT�"�O��0)4�OC�����/�MK�����O�$�O��pd�0���ff_�ڀ��2���%M��ش|�ܙU6�l�?)�x�<	0�Y�G]���!��"�,lb��'M>����ȆZ6X1W"��T�ܳߴ%�n�DyF
�?�����޿kM��x��@.C����aDZ>%��'��'Bl��7c�� �.��'fa5��I���oβ~�9���ɠt�����D��?1/O ��v��Ҧ��I���Oo9��'�
�A�Kǲ	 DA�Ɖ%n�rE�'���"�j$Y�$J�q��!@G��O�I�d��i�r�$��x��1����Ā9	�е�Ԥʡ�еA�KV�P�\��#�)BK��T�K+8����� |��	�Tp����s�)�'*��X(�3�� �T��b}���a���5$C�!�L�jQFZ�RDbd(ڧv��h)�E�u��x4��cJ�Hiݴ��)�.|���?����?*O�L��F�< 8����Ó7.x)(G�K�/C�|b`%ߤX���q�%r�`b>} ��Z�E�����nA� �^g��9j��r|�=a3�[�4w0��e�ߣ��<Q5�iR��`� �'�Lj�*۷F�T�g�Y��"�p����$��\ b�'�ў�3�@�@}ji93O�>"�`��OQW�<�3�4\ʒ�j�K6H�r!E\y�E&��|����_�?`��q�63I�����z����$����	�����ty��$, .�l2���c-��*#�[0W�����=$�s�$���r���JT�����+�(�`iU#TG�)���#�$� F�+;ℭ�vdQ:[�>#>Y�a�$�4ͫ�눚~�R�
��#��O.�d�O�8D�d�AuJqB1�F>hd@S�CG��y��*q����ϛm�a�������'+剡J��@����$��������iD�� ��V
�4�$�O��Õ��OJ�Do>A��@%kiL!<�(��I"h�����*K�
����ф��?����$�m0��9D�C��6M(&�4S(�Av�U�z�(x�TĄrL`�+Td����To�O��D%?�5/`.j����؋C�^���,�n�	K�(a�����3%� I� ��3�O���	�4��`����.J��(��ŝl 
�d�<�Tb�Vv�F�'0�X>�&��������jgN8qjdK��џ���^� jD@R�gqȌ�$���?�O���/L1`�	��G
|�A�B�K��<�bǄҞu���F���h��!`� ��5̂ԋ�5!�`y!U����O���,�'�y�N�K��E�ĳ,'�""!^�yr��J�.�J#n�-�)��כ��O��D��n�N�Z�!��[	[���O�y���'2�'v���a���'rb�'��Nڬfk|�*�	D������hM� �r}�eY�9`����y���6��8�M_a�9���;l�]�$)�>��J�/wb�=�|�<���ۭJIZ���,C�Ȃ��ß�'^�8���?����V75�T��ЀI�a񢐋��3MZB�3_�}�����"|��0����<�q�i>��My�J^��r�3�0.mjݳ�'˯��u��U���'	�'����')�6�4��΁#n��Ԋ#�X	$�<���C=���G%CR�A'E2N�?���a�? �q�����Y��
r���x*�'_7����/�� gV��)a�@�%�ɥXR๘��.AȬ��C�[�
]�G�OJ�*��O2�9�FJ�f�j\em]8,_�Y�0"O�1�0��.fR�@ұC�tRbh2ŝ|B�|Ӧ���<q#�^I��'�2m�O �Fr�V���cߟ��'[)HG�'4��'N��q��g���0d��;Ը0�D�/�}P5�W�$�3ca��@ax�Hϲ#,B<�o��<�l!	A�Ǐ�XY���E82�Dէ݅ka*�q�L��>���Ey��?�Ƿi��6��O�ذeꌫf}� �f��[�BA���<���?IL>E��g	/��k0f�is�uc�/Z7Ԙ'rў�'U_�Fb�y��IB��Ƥq��5e���k�6��O"�l�8�+����Iџx���2
�Y�I9p��I��Q�\��u���W+�i��̟��gI�"j�@K��ԏ@�bq)�	U�f�\]��N�o�T�%6Yi�5��/g����e����d�e����"� *���'�ǡ��%��˚��S
I'�a1�I1iǚ=ZDʂ�jh�aю��	ɟD�t3O^�����8�^��,�2� � T"O�TAa(ôvRfE3�i[<<�x��I�h�R���� 	����� |���Uu����O��d>z���a�G�O6���O��$|ޭWDK�P�쁺d��5aW��j%eӿB)~Cvk�4E��k�C,a4vc>A&������xݤ��g��eր�z�
��;��$�4�2Ih ��( �pc>�%�`[��9
u�2R��H5&���r�ɁJ5*��"�3�X�fX{� 8��z�K2�ZB�	<%\���&-��h�IU�',�\g���B�	���͠�C�	W����'��]�(ER.0n"$�	��H�	ğ��_w���'2��rD4�)"�W�$^R��C0\,J��G�Ü]��ٰc؅z��bVDY3zP�p(��Ĝ4�Yq��֋RA���A�DI�c�`Ť=XBfo$L���!K�p���W�X��� �\�" ���r���`s�'w"�	|�'�Z=�ץE�+�ݠF/��1�&p��'��!qB�O�mp��)�'S���	K>�p�i�S���������Oج��&!eX�g�	��m�Ƌ�O:���I�v�$�O��Ӳ�h������UMӟ@;�K߼P�|IKS(�Qs��	��*O@	��W�R>�ڡ�@;c;n��	��&ܓ��X�lQ:����C�mFaxB����?����
2�����d]�� �mͫ	+�'H��'�$×D	%1���{A��k�6e2	��l�Bo�82���`�D�&���QGŕ3�?�)O�p1�B�O���ʧ�?)���3�p Ct?#Z�S��ԍ�?9�L7~!zqgذB��q�@F�4�����B�N��&�"^/p	�/���I�rȌ����'qG��Np�O��qq�/��IzbD��AK r:zX#�O�Ȉ�'�b���<) �&A��@i� �`\�"�@�<�5���� Y�/G�@E��:r`]q�'���}���c"�QY��N1_��(H����M����?��O*½P��ؾ�?����?y��y7��6f��� �%͉m� z�aS��z$J��A�B2L�e
=Cp�U�����'���*������ߤM+����9+]�1; ��$a�$�{'䎭�n$�#�	v��1c����H\C@l��Oh���1?��ޟ��	y�'�����-]�.���jA�<m�Ů�yb�����dD�=��!bdQ����Ln�����'�ɓ��K�'Ňo����uL\�=j@Q��@#Hl��ٟH�	៴C]w��'2R)1�*i
�IW?d��I�F(��;/H4:��`ˬq��W�Ό��-A�~�C�ֹ(��tjfi�5���o�&$��q�Q��q�W�c��">��$�4�� )���(�BaRD)�)|����	��MC��x��'����>oE�Pڡ%�0B�Љe�Ԏ&'p��D8�ɖ)����g 7_�v4h�,�V6^�O�yl�Mc+O ����Ǧ��	ݟ��VN���b(�@��}����Å�����zj���I���Χ?ӊ<�D�^�N�(a� �I�Z�)�/Ԣz1 +�`�!']�!pb\^����'�20�ҡ�ӫ�&�.����;@cɒf�� 1���I��߃7R��V4{���'��	$.������ C���'�[�}`�O���$?�5��Z>	h�ةS,�]p����O�ժ�"G�X�J���n�7�]a��'0�ɢ:�Z|��4�?A����)Ca���)WԪ��	}�����៧=:��$�O�Шl��)>"��r'���T>��ORL����[��2��Jm�xZ�O����,8�����R�O�U��Z�NIj���"V:���h�O���w�'(����<��m��`����
�7acH�S�<��X�E��|��)
�Mz�d�"fS�'��}���2�e`2�5Y��bWđ��M����?I�Z�*Œ�eW��?���?!��y�/��J��AZ+]Z�(H���2�W�
X|RD�� ��I ���yr���b$2�(W`*`Rj['��;� U��EbRA[�pZ��y
� �8X'�Ռ7��4x.ۅ\����bE(��ۄ\�r����5��Y�V���{���0�M�#8�!�d��6� � [1+���ڇ�K�P�剽�HO�)7���6�HtJ�W	F�νI�֕��}	�,�Z���O����OJ���OJ��r>=p��ɗv�)���;1ΐ�C&�� �����JE�	:CE��a���/�B��D�:i�6�H>-�t���)�v�S�A;`�!�<{�9���I2(�8�+��!`���@��xp
$�O:��;ړ�O�t9��	�L_6�P�쁨8ɸ5(�"O\��Լi�� oά56�)��/�DӦi�IYy�L�
��6�O`�-RN1�#gʈ ���m�y��퟼1gg�⟐���|Z��s����&[����w^��p����TC�� w���u�����OH!����ì9&H5�'�J$�Tl<GM�	�0k5��a��!����-$�G�D�J�X���!�~�ȓp���˒��69�%z�-�?	E�����?q�K'e���5)N�uа���A�{�	>
h���4�?����C8���5U��X -�#6V���1�.bg��D�O�y D�.�\t#�.c��()3+Z8Vz,��.(�7�Ӭ?��R ����T�@+A\~R@�=p$��C���>��g&�:��0cgRH��ځ5� (p�a�Eq����E8zk�	)�~��'��>�͓i#*8��>qe�Ak?�\T��C�ܱ�v��)+q��!�0�޼D2I%�'oP�%	��P�e0i�扔@�ti��4�?��?Q�̇=�~�����?���?��w0p�cSL�q.�9��B�R��H�gC���a�B���<���j�̘O���bV��\?�!�-��{��\f��Rլ6i1�s��M"U�pe1��+V����|B��Ŷb�
�I�g�΀ГL��y�@S%G���$>?�(A��IY�'gl}�C���d��i����L��"O*a5��9C#��Ѩ�?J���R�p��4��Ŀ<� ʗ�}K�#��Ҍ/`X\1��X��Xѧ����?����?��J��O��$~>�{#�.,9 HcS���Q�VT@P���;QFX���-&��z��\x�����pjE�7F�J�t#�"6j Yi�Bۭh+��3�.6�ؠf>�(�\lPG��bٜ���Ɋ%k�5`P���0���P�?ю�iCZE:�a�,A�ps���'&Ү!�!��B�+9��c�9I��Q.M^��'s67��O��Uh e���i���'	�b�lK�X7���&��+=8p���'�2�ޫoa�'��l�og u�7!(G8����7 �$��I�JE�8(�̨1��	�'�*���N6�aGf	p`��ӵ��W`���@��0	�Ӄ2�ta@�@�'V	0�)��֬c����اBV�s��:�U	�������?)���S�O<*��f�H�UN�Ug.}�T��yr�|��i�v4C��
��l���� � ��!g�����æ��ɽAM�}�	�@�Iڟ8�0"Zş�C��&	�ܹ�vʄ�'4YQ��ğ��	Aφ��Pǟ�!�@�E�i��[?]�O��@���.y��\Q�@_�����O�����Ț.��e
��N�#&��lR���G�U��Ԝ��×�
b��I���¹��	�f��̦�3O|����B�O.Q�j�3����N�"�<�O>���0=9#�e�����
9MelE���Cs�'���>)�����S�܉p�GQ�!5|u(�	�?TX�f�'�B�'��TK�*��v�B�'#�'��N�Qd�0�Ǽm@�u)��<R�㣈sO�zb��{Od-����6�D��+Y�K6��/T$x���}�`C�t�4�VF�Q�� �+�d�.>��A�M�%���L#��� (�)�O����ON��"��ĀI!��H���&`l���n�A�<����QYdE2�x���̙gy��.��|J����$�&r��c	�#Kג�p��4q(�I`�!�J�D�O8�d�O����?�����C�pl�$�f�əM�UqS�4`8H@G
Z��̠WGR�N!���ɔ,[��I�m��NJ��ha#�33��U+��b�h!��P�!b����k�'���5N7�eQ׌���"�M�?q���?�"�S!8G�h�&�R�)���i���C�	�k���3O�R�q�Vf�� ��O4�m�Ɵ<�'=��J�A�~���=0����48v�-�F���y��Y��?�c)���?�����Ī���ʙ�%���Hnzi��E��4D������<�<Q�W�B߂�D�B�&���'KZ�=N����e�N��b��[ ~Tx�E+���0��U�I�o����O��A8Vq�����@X�cA����L>��0=y!�!}�f8)�-^H����Bb��؁�w �i1��ĥK]��zC�4&�ҭ��Ay�R�`Ԛ6M�O*��|�Ɗ��?�b�C�N�8p1��T��0�ƠR1�?��Li0n�\jjE�FN�!~���R?Y�O��X��Dޯ9NN�"���dȐБ�O:��!q�\��A�{"H Z&A$�ӂI���z�̥;q"e"���H��Ht�@��џ`F�T�'|� V��p���6)������8"O�`3��D�@ͩ��R�r}^�'�	��h�i��U�N�P�����}����cpӈ���O��M�<�����O�$�O��dgޭ�pcE�7l����0�`��>[�ر��X�0��#�O�!w8b>=$�Lx D��")LMp��3��p'�5,�Vݑa`�|�� �1��D��t�|"�R.f@.	�c�{�r� _+Z2�'�z����Ϙ'@�B#��#r���7���N��y�',��S���7�`��@�2����/O�9Dz�O{�'��}`��M�z�lQ჌IR��x�� TB����W�'���'��mݥ�	����'q�Ut�^�`^і`R
"���Ƣ��P�&eK�M�Yg���d�%~�>s1��;R��="A��=�8i��+$��)*�*Q��p=��
I1 ���fbQ��4���Љ^Eְ����M�C�in�O���b��@1?Q.���+K�p	q��dg����?��#ɺ6{t�3��źN�d��7�c�	�MK���.e��m�h�$*6&���[�mț���6I��0<���c�'���'�]�z	��rq'�_�0��
Ó*�"EFxr�>T#� �Ո��
a�l�0�0<!1����<YVM��u����c�>�.P`u�t�<I�lV.BHZ�E��@���G������O8(�K���ir�}x �;"�Z$$��v����sl=?�(�2�i^�l��3�@�Djq�`_�dP���O �0Ǉی
!(MI��	�Z�5�)§*��)�Fnz��zS�����(�'�*p�`E�DY��xCcN���>U1 ��*�z�[b���Lq��x��>?������	q�O���3Q��E�'�Djr�� �ˍ�j�!���=cRZYI�%�#^,iSm<�џ�����͛ju��`P.E�H�0� ެ'���ղy���5C.���I�?��	ʟ�'u�y��f�*��X�B�@���eZ��[�j�O��hн%�1�1Ob(#χ����#��R�x�����2�qRi�O-VSA;���y���g������-^&���A��?��O�@"�'}��ɳ'ɘ��S+�h*|l�1+ �G#�Y�ȓ�vI�ua�-�j ��J
5��'I�#=�O�ɣW�*�SW��|�q�gļ?z���Ҹ|��$1@p{d48�aR�&�(�m�	 )��GG�F	���;//��W�I�@+8�A&��F3�=�� (����	ٟ(��@��I��s�H�+9�?�'[�u*a���$�V�V�/�fDE|b.�<zj�츐F��|��S>� ���@;���A$�ȸpDa=��Q�	��l�|�BI�)P4�����5����)�xy��'�r�V_HF�`�U�����y^�ɛTFdE��R���Z�^7$RP�I�P!���?q����i�@m����O��H�oڳn6�m*s���G�����O�}�%D�'`z5�̡b0I�i�Y6.�S��+��6#����H�%S)Z�JG�^�^�	�v�C�@ȵd�4�F(/#�m���ԿdGq�\�'��,A��	E�^�h��0:O���'b������>��{1�@�e�T�'�ݷ�r���.��xR f��j߾�� �CupZXF{�f4�O������/N���5�@'�������?I��?7r��Խ�?���?y�����e��ڱE^��8��L�1�:��F ŷ*<4��v�><n�b��׬��i;�I�[�V�c���f
����,gF�!�V�X$��"êz� Ys�`5��46�4��O~��e�0M���R��*\pq������OZ�$?��y�Ie���g&�&;���yЍW%�yB�\�Dtp����,3tp��=�?��i>��	Py� � ;�f���-�)J�fm����y�	���'�B�'��V�b>�զP5.��b!��!&��4A�΄��P���j�*���⚍O�M᥅P����Gy��U a%8Ub�A��J�p�x�"7g���q4I~�؃G���`MҤ�E,}� �Fy�h��?��S<)P�ӣDM3K��1�TJ��?��,�+IBlr7�S�AI�)"3�P �Fh�ȓ7@�l�FHϭH��b��#"��'H�6M�O(˓,�����IK
{������>�U@ 	Z�8˓�?���?aTdσWԢ��EC��}'��a0�V#}p�h���[l�r�؆ZxDe�+O��1Dy���og�m���h��cqc�6t�
�����m���ӴPx���A�
2JF�9Dy$��?i��ɘO��i�IƼ�j���$��4�-O2���	�X�i)Dkt������}�!�<	g&�(����S�18�Q#�őfy���z�R�'��Ij�T�'�2$�/q_�@7 �9%��4��@�<��dNj,$R�jG�H��Ԃ@ψ/G&z�Aw"��O�&����:��spJ�"/����'`�����Ʒ0�dۑ,�v�&��垶 {nD�}��� &��5�D�sf�EA5K��<Y�M\�x��X~J~��O� ,��bAz��u�&%�$?��6"O��z�	�..ʐ��T�7V`d$P!�I7�ȟ:�;���M�q�Z(
�8����OL˓x�4I���?9��?�(O�	�� �d�[���6���:V$B�0w�iC3��O����s*�tJ!�?#<Q���L�JS�eDj��b
���
���}3��%�1u�M��O&�1���+ɰ|���u��]{џ�|ᐯ�O8��9ړ�yB��=��i`6�B�.x`��)
��yB(_�lp�@0�G'wȭ���O �?1��i>���}y2��Eɔ��A�ӓ�X0��><I\tZu�'D��'��U�b>!�#R�<�Pa�ڧ_����6>�^�w�,&�8�2c]���<q�����xU2u/ږ�R	ʃ�}���0S#�&`�2���;��<	c#��0`Ǫ �΁q��9j� �����D{"�I��r(�E�Y^b=��nXV�C��yގK&��P/@�'����ʓɛ�'��	�x�L@����f>����K-5pȀkS�(�Bd!���OfTЧ�O`�$�O����B��7]6jҢ�0)�^��i>��#�]\���F���t_P��'�>�5C��l�d�RȆ����Z7�!)�f�xg��c�X/�D�!�O���*擟a����_j���4�țp�0ʓ�0?�s�tu1�=W��VH�Cx�)O �i���}�2��ƣ\�7�Y�rR�l��Ο���Z�'��DۼQ;��b�A���'ȹax���-5��$QRd����/M'⟰mZz��d
�O�Ҽ{姉4���3#�1&��9�}�Z���9"�d�ɽ�l��ON�)�O��	�v��5��J��?"��E�<H+����ܦ����6��E���<�U}nz�M�͟k����:5M��t���͝�H�K��?QG����y"��,�$�Or���Oz�I������
P��ZAO޶S�h� С�OT��/����v���
�?7��B������Y�@4@Q�J$fw��[��gL�	ԟHbǸ����O��$�����͊Ft����`�u�o�.`?ry���	�B�$�O��.�t�Dd�8H�k�?7�� ��;>W��Cc✤KZq�㟣%`�nZ�<�ԉ�۟���Zv�'�?������_�dҨ�2� Ρ��Уs�2=	�@�'�����?I�����h��r���?im�i,�A�G��%����33�&ii��ԟD�@���ID��/&���?��AbE�����2)t����%�BZ�v�H0k��DN44��'����'S�d�?)��}8���_T�� ��͚B�|6m͗]���Ĵ<���O~��D�����?��B����jY�bO]�::T|��)�*�y�M�|�ܐ�D��6s�1�c
�$�M+���?Y���?����?�+O��$�Ok씰�Ȱ V;HVL�8��K?�	H�	��'&�h�	� K�ɹ�A4(�b�X�!��W���'Ā}"`� AĔ��OB��%O�����!�pRׂ@�8@ "O6���催)��<�5a�1+$���"O����j�b}���R�|'���"O���E-�lJ��$ ʵB+L��t"O��l�"0d3�Z<�|yQ"O�}�w�,i�0����
k���	g"O������l8�)�m��G]��a"O��6�"v��U��K�j��њ�"O \"����s0K��L����I�T�Iß��I��Ԃ�l� �x|�F�@^h��0+��M��?����?	���?���?����?���mL���HV(Ci|��S ���&�'��'~��'���'�R�'V�	-u�r=�fV�L�T�'����6��O����O����O��$�O��$�O���].��x#�WY?��[5 J+0�jEo�Ο�����X�I��X�I����̟H�	*�IKF揠a ��Y��A�[�V��ݴ�?���?���?���?a��?i��X�0i����>po!:���01��Q�p�i9R�'�r�'!B�'���'\B�'����M 3�=ⵆɲZ4��bj�6�D�O����On���Oz�$�O��D�O�b��v&���h�@���JNҦ��	՟��I�$�I����	��x�	��N"Y4^�Z֍�%$�R�[��M���?���?���?����?����?�$+X$.R��ӺM���X:f��V�'��'1r�'��'%��'����,a�6F_-'h��S)�9��7��O���O ���O�$�Oz�d�OT����RN��v��PJAGG�)ioZ�� ��������P��ϟ|�	���ɤA�Jx�4���0�/=$���	޴����O��Ɉ�m��鉎~UiN F��0!'�v�Z=1P�D ���M�'R�(9����x� N^����7�'ۛ�0O�S�SMIjDl}?��b� 
dE"Ⱥl������OƟ��O �R"(�놌�o����1Ol0�o.�i:U�Q�c�l��'0�	m�I��M���h̓�� |� �?|
�V�j���Q���syb�'�8O�˓q�Ra���.	|��q%��Q_JY�'�$�jg��I�L�!�O�i�&�H���y��6g?�S'#T%$�<�1Î��d�<9���h����0[�t:�g�9� �t�����oӘ�cu�����4�������*��$mZT���bf�H�z���O�7�O��(
b���I]�,� d�]02�ݠjJ�Hy�ԇ\#*��FLZMF��=����"�
y�l��������C1�ةNzʓ͛�L���'��1ps�@8S��h���P�q�%ːEy��'k�V<O("}J"\�Z�P6(G��H�����'�&q��Zp~��7@b|���fNd��*%�X�M��ᓵ�+���%j8����E�<	�eD�f02\`���%W����aCJ�V���ӡ��$URX	��N����"�/5����|o�L���~������
�+,�`�gϱVRd @�+�>Y"v`��E�H��f�B�jY2e��2C�9!4a�+f%Jx1�bgm)�� �7�p`���?3���F �3�ΙH<<`�Q�����({s.�1��}0�d+"Gzࣵ�$a�@%+Ec+^��5�B/6D��H�m�P�VݣLG��XPw� ?�TcX���म��q���q!��H!@�D�R`0�����Y�D��L
B�F`V�+���r��_�I�g�ISp�5[ϖ6-�`A�4C��pr����f[��D9����Nq���CI�/$��	�&Ǜ��j��ƚ6�@#��#TX}�i�|XU��O2�PYݴ�?)��)��J�ሂ/��%f	BvXy1��?yJ>9���?��i��?�O��I3O��r+�K��F��?����?�-O��8�bNt��ßx�Ӣ#f�Żf,��~�l$�4l�&��%� ��؟�����$%���>���_�NP�=�dM�����ĳ<y��X�]śW>����?1.OT�� �6]���5��-,g�u"��'1��'m.��P�'�ɧ�O>�)w�� 3�1���N$-^|h��7��I�i�����S���$�O�ܚ]��M�Qoш(����qȠ\��d�.y�>���O���1�SПD�	�2�(#��1yͰpT)ˁVj֌1�4�?I���?�W���J����I�O牦f��eU2~}����	X�k����OH��O.T���|B���?a�����C$N�<�w ˑ�����O$�č#H�l�ş��O2Y�<�I�zC�|��L���ޟ)��+��ݟ��	����	����I����	V���'��i���ݯ8Nd�����Utu �j�O���O�O��$�O �p�eY�4�j�@`�G?I-����%��U��Ķ<���?�����$ʎQb���`ɒE/!��àB�=����?Q����?Y����b�%0(���N0=��PP��P�lk/O��$�On���<1C�[	q&�O����d�G,�,�E�� E��r�'G|b�'F��>P2���X#ϝ!Y�L#'�H0W�P4���O��$�O��$�O`d���@�u�	ҟ��	�?�&��	��k0��},�mx�GScy��'9��'��'	b�'�Ӳ2v�EXIT!
����%6�d���O@�D�S^�Un��L�������?��z�\�3mD�A� $��FR�vw����՟����P"5��ڟd��k��*.�)��T$l?Z�iQW�{<�t��UI�y�ói�Iԟ������O���9����d�+D��k���%kvl��S�cP��$�O���$�����Ɏ�Hq�� 1�}�����a� ���4�?i���?�'J�5�����'
�G�B��8���D
�a�֪D����'���'�,��f_>a�O��=O8��ō"m�0h4��	<�.iU�'I��A�����$�=P�f(��ݣH^���,�D,����OܲSc<��ϟ<�'�_���(ȱhڮG���"�-(�ԡA]��	����?���?Y��?5�4Rs A	W�:d�vH��4�LqFx��'F���t�� �|�Q�� |����O�n@����N֟��	ʟ��?I��?��+�F?I�E�X�D�@��� �@hAW��̟ȗ'eg���џ��4��t�{�,
� s,`ע�ҟ�?Q���?iV�J̓�@�Q,Q93,���C��z��	����?�*O��d�x5h�'�?���y���>a�h9�/^�l�$�FLI>���?���R���<�Οެ��a�F줸1�[e۶���'��e�֦��O"�OŶʓ.q ��ZШ�G��K����%������Ѓ�F�P&?u�o��'_s�t G$�?XL���2[r�W�uc��'�"�'��$V��'���U�<)j@!�ƍU����?�F�>���h�0�d�+��S��� �0FÖQ��n�ܟ���՟X�!O�9���|���?���$`;�Q�7N�S�0��ʑ�?i��?���>�4��+���'}Xq*sgQ�I�hM���Ù#$P��������&ԱC�&�A�c�1 "�s�iMm>ze�4�'��'��3Oz�:tDF�n�����[�R��Iۅ�|��'�2�'tB�'B�К'2�W=Xx����:_�.$��J"�'џ���ןx̓���֮S*wâ)f�0��G~R�'��$�O��d|>	9�E��k��� "ˑ��nl��c;��O�la��8*��)���O"������S�&-��D�s<��J�͜�C�I�:A�MaW囂�j9�F��V�Rc�pX�:V��$i��\iD#�A�odtу��M�lP"��4���;mz�R���(8F��ħǭG�ryX'�*O�f=�B�3s�,�������'��6>\H�G�|�� v*e�?��X�7�t���͂�]�f�#�k��O�d�wi�3��`+v��)<�*��HV-:���u���e�Չ��F&r����/J�I��T��?i���.؁��	H�L���PG��q(�?��O���:�F� ;r1"p�A7O�\Q'�+ .}�ޱJ �S�3ĝ�BFZ=\���\>��≟?2㤕� 
0&�!kT�.�D@`�2�nӼ�n�؟��~z�	��hLњB@Px)�q[��ߕ'��'42�'�P���	ԟ��� �t�g )i�0\�G�x�!|��LmZ�� ܴ�Mk���/,@HŸ���7����W�E?'A�7-�Oj���O�̉�b��hU��d�O0�$�O��X�n�P%�S������ nd���f"6f��Vȑ2F8�9�!��O~�6����?�G�V#��dy�	�DC h�_.h{�5x�	�
g�L� �Bǘ/D����D�i0(UϻH(��Q+��(ܐA�ꈓ4���Gz���'@��	��|����'�8�
�o���I�+�&Š�`
�'� �"�\ i�� �H� I�D�����զ���~}B�;g� �p�%j!4��0��]DBp��. <�Z���O6�$�O*�;�?)������K\��]�%c$�V��!*�>N����^�iE���K�-��!┆'�c��#.Ѳ{�(4��L�g��� .�88�t:[�����E0>����1&���Z��¢g2Ew���GH#T���-�O�Z	b�T����
�o�&E�� �y�!��<ṱB�*5���	��[�¸'c��PdV�M����Mk�C^.7�>�fb�: ���$��F{��'��*��'D��'��<hU��5)Bt����΂u:�[��Vap�l)9_��RҦ�TX��S�Ԑ{`8��F�9�R�*a��&!߮xi�
�z<f�7+�$�����v�Q��h���O�	nZ?�M��4LX��pp̄>!��!�3HR�K��$U�Drߴ��D+r��4֧tch���.h�Ѐ���x�*�l�F�+U��3!O�A�#�)�V����i�ªi����@I�Zg��$�O
����T�F~�ƼySO:mh�Mx��Ё*�@���iLٟ �� �ԍ�R�� O���蠩����3P?��O���Ѕ��) ҭc�m�h�t��K<a5��1l�X}[ aT(nD���Z,_��S�|I����?�P�9�O!�t�'2��O���t�fm�C�����U/�h��"O<ea��P�d�Z�ٳH�9R��=X��V���d�&ʓ|3$� mۙL�q5�W�)x�g#rӬ���O��OPЀ�O �d�O ��wc8�����i���R�"'$�H1�p �6����U�aӲh"��,t�t$?�CN������^����1�	89N���t��fa��MW�M�4��)-�6�`����i�k3�f8�"C=2�pd^6)��:�j���M�WW�X!`��O���=�����mڼs,������h܋a���u%�̫�'(�����)=�L��G�R�ԭ�~��'�X���?���h}bE�8��@)�%V�S�=b5��:6��6�%7T`�$�O&���O�D���?Y��������%Cw�T7�4x���� �@��n��`��`	�(�]���P%2��bw�S�b^��>\���k@N,LO��(���K�0���R��^������R���'L-2�l�;���Ƨ��B�Y��'y�E���S&R鐠��!��_
(�{b�,�	0 gr@"۴�?qߴt��Q6 �-���j�d��(�qJ��'�Z5 Ab�'��)U3B�"Fi q$�MY�S%A�P3��cw��0=�I��	:Ⱦ�:���-����� "i�ј�U ��h��19��Q�A"@Y��ß<�'�:,(Ї
��!޺�� ����~��'�2��I�,���R�I6���A?2����)F�<m3��T���K�2p����'���V�����4�?9�����&}�&7M�]��T�G,]�sw�� U�Bnz$��Iݟ�X%af��@��Od󄈀��P���	�~r�	��ZT�!i%F����  @�	���aHf��" �xeA�m�%$�ĸ�}P�
�NZ���"
%p�ȡ(Oy�!J���ަ�J|�K|*�*x�=�ѫ��MҼ�Ct�%�qO���6�d$���LTvE�ԏ��d��"��c(�����!��4��ah����R�bݢIq�!0�T��h�N�D�O&�$T�j�����O����Ob��w�H;���`2�qg�(���	��Ťz�D� ĉA
�(�o�b����']����D9��X�F��#7Yr�c!�T0:���؄Q�̐yg�J�ym^�>=�@Ê!�y'C��N`�&��8b��Q0L*N2��$Ty����?�}�I��n�B�@�KT��!a2�[D�8z���^eqO�X���P�	�T�D�1ෝ>��i�7�!��?��'��Ipr	�&�b�±kI�fb2�*�)ݺ�đ�O��d�O��ďݺ����?Y�t����%�/��C��DT&E�ÀȷB^jH��(6-���"C=,O&P9 oJ��p}����S�����2����-;����nPsX��Y��ҁ�j�k, ܅���^�X���O��n��� �'-���t��j��"t-A4�ʸH����	�$��R؞�K �̓i�N-"�[��&m��	>��s��&�w�˓"�u�%�iVұ� 8��wX�{��Qu�Ũ�՟����.!���	ϟ��I�Qm� ��ÖxL9�k��
����5K��	H��6G�#Y�����'^R�k���W�αh��#A��y#�ߢTB�W);9B�q��."�4�K���
�4��eh�P�oZѦ!Z��X�e#�%�rh�q��Xql
�����-�?���)�~���¡A�)tYd��7��$TC��d�J�=ZPk˙d�aȥ�uf&��'E�u�'�>6-�OP�$+�Y���t�^�Ix�����}�zA�SI$D�d�B��7ӒpH�,ԉK�rUҡO4�	�u�4ը���3�ʀ�fd�c�P�Ol� w��(y��]*rHH�7���8�"OFX����&ܺ�WFƽw�h�8"OHVeթ1�rR��B4}�&��"O��
����>M�.4e�8���'ے@B��?~�����P�Թ�	�'<��a0�O;1�tڰ�IP�
�'d��Yt�@%�R����Q�L�6xq
�'�H�p��<�8�)��޷E㚀0	�'���� �נ`7N�rW✔�j`	�'��|1���)ST�y��K����'`B�AAm����F�XF����'��lZN���,���N�~��	�'�HI�1�	�a��<�Iʼi;����'e.�#3B[�7�<B�E�k�����'��(E)(4���#��[c֎�;�'�Ν
�뇳GX����? f�Q#�'ְ=��K�*��V�%ނ���'r��*��w�x�e�3�6m#
�' R���l
2t1`&�y1��:�'�I1'g��O���Ce-<b��9�'�Rl��*��>��ܲBEb����'�x�EM�@���$�� �$�h�'��D��M)i\�Bg�����'{P��S���:��B�
���'�
�����0*��1�$J���v���'�1���*<��4i40�
�'��qj'B�}ޠ���F�yB�	�'�>50�C�!dm�m�S͕&Mo^�*	�'�BD��	^x�l ����o�-��':,Y�0�<D."���@��s�����'��h;��[yP��c�0L�	�'@�Ș֯���6H6R	�'������P�"�"в]ߨ�0�'��}J�HN;̎ PMJIW��
�'2�����_����7ǗY^h�
�'�&���
���H�;��Gn�.M*�'m�5�%D�q��X��'a�m��'ܡ�g+/	��\C#�"h�v�9�'��$X��Xj ���HX%k~��*�'����.��^�D����fh�a"�'(yZ�JP�#�8�"q.�S0X��'>��ҋ�6���)�C�7UH�
�'�HBd���Xֳ0�DdÜ�y���,�|e�R,]*��B%mڷ�yr��5|�`K��I$^ ��2���.�yB��X�&�CULӓM-*��#G&�y�IӖBG>�i&L��C�J	�d+�y$�9~j�V�(=��ȳE/˂M!�C�I��d��㋊]��@ZY��!�'SyY��_&�D4Pr���5��'Jܑ�Dճ?�Vā��8x��{�'kr���*��'}l4J�$�
LZ�x�'���R)�-&�:%
��k88��'�>H�e*�^j��įO2Kd��
�'9�%���ډ]��h��Ȯ)���
�'<DBcO�4)_� @�� >;�pq��� ���!oD�Y��)QM��k�=OD����2�p>����2f���p/M�*��}Y�X؞�q��<.�����'��L��O�.~��d@O8�� �'I�<�օ!6�;��S?:/T1:�y��ӿ;,\!�D�k_�F��!)�y!"C��$غBG �yZ(��a�]@7FT�*L�,ُ�!aa`D�?Y!�4����I�����H�i{t��S��C�It]P`h��*S�<$sSN�:EyX��E�o�
35Ⴌ��ɭ��l3���#��y��@Z�?�R��S+F~}��〶wT���➞c�H�4	ɺ)��q+�HƹB1�0�'����L��!D�&؝��aPI<�C�B�84��� ���=s@`$�ӈ
D��Vn?�a�$N(`:B�.���c@Y1'�α��mgV*�b !Y�=�	C���;.�0�@�#�SW�	�n���%c�-������H�
��$��{�B�r1҉q,�E�uf
�/�(�'�D�y6�x"ٶ^o�D�o*,O�ajt�R�8�@��sL�*Q7���'��h*�FN��^�0�㖺}��0V�E��lY�T,{Ԛ ����b�!��|���p��D P#n.��I;?�T��Rl-2�\���T�� t�ͩ焃4V�ޜ��$�
�y"dϣxeP����W��,�5�X�HI�����
dR��R�j
Z����L~r�J*�DIor�[�	쮙�d*�5�a��Z���TA���+%�	�di�/.�*%��~�
�M�#H�����/r��򄛉n��|�F�.+�Ͳ^�\]�����7lx�drCɖ�ru�#��'}�@`����I���N��9��	�J�B≓� 9�-k(�:��J8l���fbA�0��A]��Ã�
a�Q��6�S�Y[��Z-O�*�n��EJ��C�2�bX�5��
�0�g�s���`�+�7^��H��a��Pv�aw�*��C���Q���;��k�R""��>y���	�=r��z��)2�x�{ؑ�(E	]V�B@R�Q�'a��\�T��牐,W`��j7�n��0·�Y��">�e��OwH;#��{��h�˚�"_�0���D"���!���L���g�]O!�D@�i��뇪޹+q����X����޹|���g�MӘ	m�������=��OtBe��Ku8���,�m�P�+�'���y�ڧ~���Ũ-(	�	��PѸQ�G��=)@��"gS���>(BO�Y!���Ft�Z�EF'HIP�F�'��x O��h|q�惐$���""���C�<�rDpf#���b� /|R�8�2�P�<+�	�+����&!��P�D�-��	�� �!Tq�mä�$����'��4@�Q0E�b��N�R-&�2c W�� s�dP�z��!��d�D�6���dI!p��1�朶M��D��
K�J'܁{k�E���էA�&���	a�'T�:蒧lM�BlZ��Ư..~i�G�B�|�.��d�)��8���:C;8ı�1.y���@��'fP��c�OI�8�W>�A1�Qu�'eV�8d	)��(���ͨN��r��y�Ԁi�йhZ��pFP�li�1�K�&����&�H-m H�nV&��{�{�ӌ\�˧!�8L��h�jZ��*�+�lCRE}r�[��9���+Q�r!����#�>DQ�oJ�0�bAЃ��q�(��2N�%�?�`Fim�?���"1Rn\	�@ɠp��HB�JM}b�� N�k�'�)RdP����+4�"|
c����I��
�$jw�XطZD�<Q�&\KVX<�%啧\���j�l�7h�a�4%�"^QZy��˨tˎ $?}�<i���?.5��e�O>�J��p<a���$Y{H�*���R�d[6hܡE�����/snB
�/ְd����dȵ8zz}˄�:%�E/ay�)W"u$R2kJ� Z�II^��/��$|"Ү�:U�0B� JR�;'ײ{�2��Ճ"<q�CC���~�UCV�pcp��%"ʿ4�*�:D�|�<�bC�S�b|{��;6X�+S �G�<�=rYZ���Q�n�bpJ	K�<��ͦ#n$$@S�8B79s���N�<ɀO�3<J92G��2�4M0ČO�<a��<�~d;T�5\�]C5)�I�<a�kx�f=(a�ܲ%�vTSbE�F�<�D"�]�Ta���סq&pKA	JB�<qR'��BH0�)��6[�Z���d�B�<�v�Q,P�]�q�_�"@�kA'�~�<!�`�;?����G',0Ti�a�]A�<� �2d�LQva��HB2PA��"O�y��Es�@��D�&YJ�bR"Op�3$�C��U��%��Z�.Uh�"O@��$��C�Fщ�.M�$���""O`ِ��B�-$0�b-��P0L�u"Oxг��V4Sn��1��Ǩ-<fx��"O�� E������p�閍+ uQ2"O�� cg�j��Q(�(�>7�d��"O8���"�-̚�ز��[�*u{a"ON�֢�T��[�A֌����d"O�P'�]�����*��H)"O�e����9?�kV�� Q�j���"O���g�9KQL��7`�>H�Αi�"O@�a��F'H�tT���>˖ *�"O �b2 �6���M��i
\��u"O�DsD�S�	9���w�Kk����"O���#�F�c^
}RE�ӷc���"O����.���s�Ƣ}���5"O�-[S�b���z�lˠn�&��C"O�E�W�r?����KK$0���2"Ot��kU�@ư�he���`^ڲ"O0Ls&O��H�n�+x$���"ObT�jr���Y���& �I�"O@�w V����V,Ҥ7��kQ"O��9p�ø:�\y[ua�J(P���"O&`Z��_P�Qp�N���=)@"Oe13��*M�R��'/'x�0U"O�e8��m�<CR��9ep-k0"OB���摦m+@}P͗�lz�c�"O���#�\fؕ���I�q��(��"OD��!S�H�r�c ��Z��)�"O� 镅l6���;�pI�"Ob�uF �����ÇC�N\��"Oj�y��+*?�ѡ�!̬Ժ	 @"O��9ˊ0&Mk��_�U�2��w"O(ݫ��E('��GOP�`�ڼBQ"O�5j��D�=u�� �Oޕou��5"O�ܛG�ޢ)/�|��c�-8S�P�"O��i�i\�`\�P�3�Q8	B��P�"Oe�Ռ Fs iѫ�;���a"O@�Q�GׅpDf�Jb� &S_
A��"O0� ��F�.���$k3��"O����j�*D������o?���"O��`F@S�j�# k�m�ʰ"O�͢��[!**@ϊ5�#�"O"RцY�L�UZ���G:��2"O�ɔdZ  P�7&%L��1"O� x��ޯg�x1t�J=�Y�a"OĔ���G1jѬ� E����A"O�����g�TTQPᙩVT�ah�"O�]���b��,eQ�S����yB!�	�^�0�C��m��qDL�(�y�b�,p��v_/XfqR�
�y҈�&Yq���#�I���U E$Q�yn�,+2�%bļac�Tbn��yȑ0�8��GeL��Q�A�A?�yb# �:o�i�a!]O�Z�
���y�)�1+�i�	O��-z�j���y�dO$|Ҡ��9?�x�����y򬐊���0�ͼ$�5A)�:�y�GҳRv.�k�� UF��1!�M�<�F�9X ���֤"Z���Nd�<��J�xfn	�
O&S��e���Hk�<A��1����#vL�xC���<� h(��Kޗ����'N�M(,B"O��r-�MC��C�������"Ot}��F2S��ŉ$u0���"O`���eٗR2�s�OV�`�<��"O��2��0H�A�C��$Z6\K�"Ob�s�� h��sa�ǹW�ָ�"O��6�T�,bLC4@&����"O�|C�ơ?�B<ye`U�E��y��"O�PA1���0��PB���Bd��"Oz@x��x�
YSӊ&K���+C"O �)��ǅ|�>j���G��|p�"O�Xӂ2y��)q#A�V��ڇ�d�(@�bѻ�����#U�H��'��4�'jD�dr���E�Y-��9{	�'�ٙ��O�`´H��0{���c
�'(����(	Z�8�)���"~ ����'5�+d$����4�
}U���']�#�i
aJ����a��}�'�,܊!,�C��$@p+��`����'J"L-){
L1w�Ѻx3�Lsv#�y�<�v`_�U{Τ �'W�;�l�:���z�<	�#�gp�:���-�RV�Gb�<���3C�>�1��O<u3�q�Z�<���6خHQ
¡kL2pQsa�X�<� �6>4��nC�Jo
ݠ@��U�<a�D1s���#�{U�x`ӊ�k�<�1��1�6I��A1E�^��]�<��EB.m��k#��):4S6U�<�PbQg�&���(x��0���E�<9��N�Vx�,�lPv�.�:��}�<a���![Cqqp*��/h��"��E�<!RF 8���P`W�"�.�AG{�<�@�-Y&�kw�XUX<�F
O�<���*eH��(q�	����t�<!E	1I����5C�<O�v���DGm�<1t��)08͓� C�]�vQ�B[D�<�R�OfH�u����	b�L2С�K�<��J&jB`"և��t�q;��1T����(\�[��`�A錤&�A[c D��ʄ�˺x ��1�� �L<,X��=D��Х�%�ށ0��-��D���'D�$��剕)��Xj7��:~��
�1D�гB��0���Ţ�2��s�./D�U�&q'�٩��ȥb��)�8D�a�Ą�Pv���C��,D0�,��
K07�3S�RAG�4� '&(1��E����ݤb!�D�6q���͐
w�~,i�i��W�hQo�9`^�r��OT����Y��XG�]Pl�#'�R3[1T�˗�8D�D���G�8��d�wm��Q��%�W$\|5�FY�=W���/LO�C�nS�H��q�I�}�Hذ&�'��}��IR��1��wV���&������	�3�t�ȓ9dBb�� �oL� ��-@���=A�� ��#� L��#|rq���|�ɈN/��8�gIY�<Q��\*q�d���'8L:tY��/J7�̤�F�X���?Ѻ�|�'�J��D��sZ�2�`��@���!DpЉ�}��h�DzA�&�1�Drԁ�8F���j�L
z��\
��ɕU�P)2u�=}� j��5\OL�qK_?w��bq!�2f`.�����=���i��,�bi 
�'\�hE�J�Kɼ�	'�]TX�=Z�{�&
lt����P֊\D��"�t�$�&b�9}�\��%Lݪ�yB@@1a8<�� @�(i���A*X�h��˃�O�4���'A�EE�,O��"h�?q���H�+!">�s�"O6�ZŅJk��8�Ө:5�]0�i+�Q�g�1'��@��'U�ي$��p^�
�����#�x��P�V�p���FJ�*Qt�{�L!�i�QO>D�� t��Q��V�Z���@N�A1u�	4Wt��U��O*�3`O; �`�:`���]��HC��Cv�����x'$=�B�ֲ^҆�����Q*��sJ�3h�n">Y�C�0p���＼���Y!5A��Zހ[5K�:�y"���fՠ�n�_K2����1��'�2����<�Q�Κ9�~b>�(c?u��2��
P
�l<�O*D!̒�yR��*�}����H0�P�e@5$�>�S� ���J�AU����')��[�	:
�-����~u����OuY�e���M�&Z�-h6e?�gy���xU��c� �b�̠�wN��I+ZЊSM*�O��H%/�5,~P�#ң/\��c/�r\�������]~��O�q3����k�;��x:�H�����^o�����cr��֏�^ L�RrI�6lڂ!����~¨��y�NP�x(� �M;��$� C>��үG8=��`�'P�s�џ�6LZ�^a�U�c��� �� H ���.A�={d/�1Pt9���:k��lڒ'��'h�h�G�[p�'���	��'���W*��Bu0+O`�B�O� �h��ɜ"�BlcZ��O!����@ 9_vD�'Oڃƕ`Ĥ�){���I�0�0��`��}���`��h�h%w�*L��ۓW�(�)��>0<��G���oU%J������ēX�I���!�3��7@��C!^�,��\��J¦�����'��<Jq
d���Z/"��I&����1��(�4�wKW7T�?�2�׌{� �rH���Q3��T.�ΨZ��9p��8aP���laO>aT�������9����O~1�'��0 c�ƥ:��D)�h֩]�:�A�O&��VBɜ3{t��N�>F��ԺP?O�g?Y�$t�d��G'/��Q�a�?�#�����D�1Z|V��-�[�Ҵ:��L#IND�j��Ynt��%U�3��5��LT!F����^�?�$���1ϩ>�G�:*����&Y5<f0��);d����a����|�.��E{��@́:ސ$�'@�<q�2�[�#D�a{"�O&=Kv��W�]9i�D��.~��L3P,<O���PM0V��>�px>Z����藼B��Es��;�A��㧭	�h~�)�GIg�p�I�(dI�k�6ָ@�,PTH�e�R�49�$_0 �C�L��~��;+ܠ��j$�IT�KnP�r�G��բ�ꋄqd�ɷ;��j�%�$�!'�ׅJ�(#=A4��,l��	)%n�H�<�sd$3���4o��@8�)�3 s� �Ӓ~�<�h="�+V��5b�0TN�2Y���(R�"5Q��Y'�K e-� 5T��6��7s�>�"�ϣ|(�1QAMӸ}2��;<O�0SE	�9��:��\5�l��W�݁o�|�?9���9�qK�j�2ػ�Ћc�1+w�8�����#h�@5sd��"}�Y�c��>@���#����Ƃ<�|6-�,[�*�K�L��$�j��Ğ32Ͱq�Z�
��K$���&���6'�;W*�I�DЩd��h��Ծ��t!B� k����ݢ��H+S���0-�I� l���NJ�z��k�D�u��"=�e9�ʃ䟱4bٓ�

 M����+�~JQ$�n �O��I<[���jYV��&eW�0o��K���
&��E��mՊ(�v�����|�c��Jj֬S���*���ચ�AJx�����|��4cI+*�*�O:�IK��ߓY��tL�=r��Klf}�+�Ƶa�
���2�F�#����W�D" ������]P�x��K�C9$������Q^N�KW3���6�N�IS��d�A���ʔG����O��IҞm��`]/*��M{0A�� z�(�"�"�)[ч�K���E�<�H|��*#F�x��.qXT[�K̽X)B0@�i���>yT戦U\��Jb���`�"�"O�'�iY�iE�dV�y��^<bor���N"��ɣ(S��ٲ��f��U�K�#���dÓH�TiᠫN�K�����F����.zjź` ^��	�_���'h��2�$�V}�"ľ.�^���㙛VLV�!��� ��O:y�B����'��t{@H]"��y֯�([�zTb�$�ɦ��Gl-}R�ų�D~��	�[�� �nOԞ��'���ċm��Px��/}b��7��y��~�u(�_�D��sgB9{þ��c��pR��A4�O�- Q��H�hl`s�A1>�T5*A�>���@�B<^�kV��<i@�Ox�P�T�L�`�Y�_��lЩjL��+�L�f��M��|D�91�X����#<�L�Д�ೆ7Ox��L<��z��a@�lcP�.e>���g��}H8<�ȓ<V|@�C��. ��2T��8E �g�D��@���?�':�@�&�F6_�<8�.%H5i�'Q���n̥h������N�c8*�ہ'�|l�]����9��@D�QE:%��`I����DT��:$�H<��'D!Rt� �v�آR�hE���Y�<fŁ:h;0l�-������	z̓Co�豍��Ă�W�|�Q����j�*D��y�"�0�n$A�-?�P1��I�y�ě?���Ơ$y�(5q� �y
� �X��g�ε�b'�
?�����"O&$�U2T��U�`fS�Ĕ�+�"O�-� EϘ$��9��<B��̪�"O���t�"{n�y�RM�&�py1"O��C�BF�]TR�:E�K���"O��@��'E���@r�S�4��eX7"OZ7��͙��I���w"O��k�7`��`�w��'Ϻ��"O<�L�<��A�F&qm� �"O"�ϓ� E���ĦOi��Q�"Oz����'j�S�4M�فu"Oj@{����N]#f�0(� � "O=�����@�&M&�ɷ/n.!�
*��)3�fFT�Z�M^�]'!�䛪su�@E�F�q0�cW�$,!�� .��0TmM#z�ޠ��_�}�!����� �5�Ġ��K1�!򄒷 uH�9TjK*��l��D�T�!�$�k!2ujt�R>G�"h��C	�y�!��D��A2���s�,y&�Py�!���yX�ka�t�V������:�!�D�<�A��#۾��ѥ0�!�d
�mR�銊~�Yq���$�!��ҿ B�ծ[���%c�?+!�T5 �����ٱv؄�)��({*!�d0 4���ڃϐ�BՊݪ!�DI������m�.��\���_"!�\d�T�9$cB�7D�5�t�'�!�ċ�a�^H�S'���7��)d�!�$Ŧm~m�P�;��o�/h�!��W�$��q
��|	�H27�&^e!�dQ��	�!��{�ج�㉮l>!�$��k6U2��P>�L�Q�� i�!�SH���N_+sǞ�JZ�����'����}w�g���>r���'`L(�UI,�yq���@9Fl��'�l�9u����U�1lL1�p�
�'Ⱦx�aM[���Q�d*#h�h�'\�z���(�ǀ��%�\��"OB�B����<Fj�J�G�r���x"O���B���_l-�1��X�J "O�s�G��0Na�D��B�����"Oɒ�Z>s���+K/q��Y�2"O> 3�0��z�i��q� ��4"O��Q>���wB�3h��1b�"O
��5�3�e�eAQ�,�"�i�"Oр�ҜJOԳ$���($�3"O���f^8;��q�6��(f��z�"O��.��1RV�5S�A��"O�X�s����\2L	f#X���"O20ؖ�˗�)����"#02V"O0��������%i��8u�Έ�yr��1685HPM��2z��/U��y��E���ɨe��
f.�6B��yb���dyޜ	`��{]����y��z�NDBkAd�  ���M�y¬�VL��T�\!�P �y��N$Q�4(�&��Y���u�%�y��PM`	PeA k�)����y�`CWm�ٺ4��+�h��M�8�y��Ԥ$z6؃$�!2��P�;�y-L�1C�=��̂	���+���y�d ����%�L���6gX�y���#^|�e��.1:�T����y
�  
�W�or��Ĉ$>��"O�$�2_/�d%�z���g"O��+�`�0�C�Y��zc"OU�E*�L[4�(�Yl�F�xb"Oj���%��Y(�'K<j�~��"O.��`ʹ,�`K�EW� ��4�"O�,`Ǌ���7�O6��"OԩY@�B:YK<���ϰz��}A6"OrŹ���׊Brn�x����3"O��yp���?*4�1���Q���"O��	a�Z-���a��'�P<�"O�QD [��HAB {�� �P"O�A�kE9hQ���Wj�n\4(ȑ"Oj��
R�:j
����k���"O����,�F��8r'����ģ�"O~ [��s8%���Ԍj@p�(�"O>�8D�g��p;�A7[*.��w"O�8�s���g|�Gc�,>.��"O��0���	��D�S���%Ѥ"O&����E�4�J�``��*F%�ģ�"O��{"�-r��u��X4~B�ؠ"O4]�2��L�q�Ñ5�n3�"O& %9E���Bc�0�J�+�"Of����  ���ѩ{*�1��"OL�p ��U��؆�̩g7�X�"O��9& ��iHd�`�E� �����"OЉ��0l�n��ĎR5��9��"O���PV��e�#g�N,cU"OȁI�i�2�x���jvnp��"O���� ��1g�Q޸j&����)D����MX�3w��ߌ$����`;D�Y-�e�$|���"d��aV�%D�@�FE��]Z� zAf �;���z�"D��y�n�:a�e(h��e# D������a�Ш�"��?���	>D���Q�C":�@��'�tQ�E&D��)fh΄]��u
�Ď7x�����b#D��s�m�c���tD��d��%���?D�L�W�.<랑3�#4ٜ�i#c<D��A����Kva
mк9}��3�h6D�l���2K�$����oM�A�6D�0��
�qIf��H��~o�M��i3D��æ	��oڸ��v��c����1D�PS�IR�ը��`l�0�t=�Ҋ1D��$M2|�B��d�=XV�����/D�P	�c� 2G�¢Iɠ���5+D���C�(
h��#jG�9j��T�%D�lZ���J4t����}B1�+$D�$+���Q�<�SC�S�^i|y�>D�tRT�G��-���Y�1D�8U鉋	I@I�%P�e�Y��/D�p@���N!�:R�� (�̰Z2-D�@���< ](4��$��B�ɓ	�
9��&���K�掲H�B�	�vL��1&�B�HD�ArE�E5 B�	<D�D9�'���T�� $�B�	����]�R	T�⢌�:N`NB�ɑP� Xb�1B @�`�\Z2JB䉘yT�����I0d��-� n\0:H�C�I�^K��p��̱S��APMA��C�ɛI#6틷��<��'F�Zy�B��o�|*�BK�m�nX@�E�v��B�	�[ �m2��
�ud
����%ZjB䉽g�.ݙԪՁ�}���;g�LB�)� ��U�pˊ)X� �64!va*6"O uX#�C��E05N��G
�J�"O��2��א�(�*��FO*5"O��x�����ū�0NJ���b"O�=#S)N�f��cpØ.VBQ"OT=jc(λ.�ZL�q(
gCyCS"Oء�#.P%*�>m�SI�	^��p�"Ob,�'�ݔ%�v!�Ce�Db�0z"OB	#�CB�V������I�bx�P""O�(@b��j�2)�HU3Cv��B"O��1"��|Y�a[H�(WF�Q�"OZ��F(Y;����f�5۔�q�"O�\�Ή6B�	��&χa��p"Oz�j�����j���*:�RG"O�4ڳa��a,�*����n 
v"OB`I���T�H�"7+у<����B"O�:��Ȃ6�Z�r)�/G���0"O�GN��yx��kN ?X+�)+Q"O��Ãē�s�	&�+*��KR"O��F4l{t�jo569�"OL�Y��,��gor����ÿ�y�˓�9l�8'M �n�z�Æn˰�y�J)_Į�ƍ�a;y6-Һ�y@  ��Yj�G�D�N�s�����y��)��̛��Ŧ;�đʗH9�y�KY�S�N�I�IBt�0� ��y2">'`$�� ��f��E�gP��y��=R�����Q�ZA�Y� ���y�M��Jՠ�lO�	<�i#SE���yR+��)���� �{f�
3�D �y�c@4 ��pM͋x7*�S��(�y��*aX�I�hz����B� �yr�O�H�p��@�Ŧ�>�
sEA�<�rDl�t� (H:��8��Ef�<��*V_�	P���m��1�Śc�<��P�Rv���b�	^��r.�c�<���k[��ɡEE�w���qB�v�<�`J��z�=�$��@%���J�<a�`O+*p����1|$����NG�<���: ��G�zs���e�E�<�7OK�l��GF6pPx��#�V�<�$i��%�6��B��z�>}��^P�'�����*nz��a�k��Yf�`�Jպ![!��K2�كf��?Oj�ys(N;qX!�$�6k3��J�@On�fļU6!��M�{@d#���6l r�*aē�W�!�DA�{����^�4��1��8N�!�P�zD��:b�;LH1a��}�!��3���ZDnϭkSRa�E 	U�!򄈿�B�bʉ~��`��b�7i!��7��X)v� �V ��!Ϩ<�!�DLh���G��N�9�Fށ_!��\�8�ر�O�0:�j������b�!�38��a[��ռ !|с�9
!�dU����h�X�$Nuj�B^�!��Q���kb���i�P�a �ͨS!�$�@��(��P'о��G�N}.!��9z��c�E;z�8��e�.O!�$	�M^�@�蒩�2	��$�c1!�Ě8<�L��e�A�s��$�3�!�DV�U��՘D�!q�@�A�w�!�d�R����OU�DWtih�A��x�!�dZ�S�����Gv5�a�$<j!�.t��Hh!�ȉTֱЀ�\� K!�� �\3go�5V�4q�� ,a�nX5"O�1`���D�� ;,	��"Ot$ڥ�W_:��"�!k.84�s"O��cw�2P�6y�G�N�zL�P"O:�ش��6y�8�� ��p����U"O(鳥cĂ8�f��d/Ν��@�"O.Xe�_�K ec'͢Ag2{F"O ����8��Ѡ%ԉb�^, t"O�h�@dU����ADǑ7�Q
�"O���ntlE/dXM���G.&!�d).]�i�H��/��5rr'��z��VH�
VNאy_��U���y�i��b`\�#�\��T�;b/ݗr�*U�ȓZ�q�C	���Cf�s�p����dA��>����2<p�ȓ��"�� ]#p#F
����ȓ#��I����/yj��I.U�NɄ�E�	Ӆ`��fd�eC� -��8rEX� 
rږD��l
�?2���Z��Ԋ��zA��8��9(X<)��}���Z��]�{�4h0CP,L�NՇ�Li���5��/vXD�C!_��RԇȓV%�brmҩ%n�ͱ�H,xOJ��l0h�%ؙ3W�!P��$���ȓe�������r��%��B�=��(�N��U�\x|�k��$V��5��@��!��І���' ӻU�ʑ��A&q	�&̘ ;��3`(�r���ȓCI�)�s&Ŏ��LR��'uY��ȓ+~�k���?m�*I� @M)x�d���i�9rb��J1н�-�,c���j�c#�&\Mʼ�o�~4I��]1@xa5�@q��!g!8b�x��/劈�B�J�d�F 	8[[��ȓ|�D� ��'0]L�:u��6tC�Y��w�X�Af��.���P.�X}ʝ��q�x �lG��<����1t4������YI�
;`^$P&bU�Lv��ȓ]g.���5�n��0Z��0��ȓS+��ЕKνp��%Q�L�OC���6<�)2u\>fc��� �Ŋ����X��u��Qt%�ā1FJ���2�9s�
�*|��0KϬO�}�ȓ"�Ș��d�c���KDEc�� �'����`ʴ=�8AԌC� X��'wP%���B!B!@�cSl�)7͚��'U��A�{9�RB�,��8��'�2��LPRg�hY�g���Ɉ�'��i�m�6�n� r'� ��u��'5�z�Z�����S�
�NШ�'�D%C�.��k-�`h2��NH��
�'̪��n �ij��^����H
�'Z�)H�&�: ��\{�� ��-��'ax�a�4: �fn�*b�<P��'����C�9&Gt��@A��.6RՋ�'�N���h�N<�@���'OZș
�'8��і'ѫOb�����30ChI
�'z�$l�9ED�W],�d	:�'���Zb��:I��m���	W``���'6��6I�P2#��]D���'Հx��+"�DҒ�S
gd|��'|H-c%H%u�x!@Rb�&Z� ܚ�'w���v���Ҡ��(��a�'�<3@`�Y� ��V#n�
��� �6��^�`�jT����"O�yc���K�X���&�9���z�"O,H��#�	�e�<Gu���E"OȰ�G�	\�I�F��l
e�W"O���� �Hj�Ѳ%	�|��"O$Dr*jT�3�J�"�~�P"O����Ć �%�t
˾}Fq��"O���=l�:x�J�k��$�"O4�:��OӾ��Gd�ex�
�"O��s��S"�RyG$�D&�`�"O��*V֝M'���7d&K�"O��9P��h&�`B3��'%�h���"O��x��	l�����~��<�"O�	;���x.�Z ��6��	��"O��$޿-� �2��e��@A"OXͻ&
?.�Z��ªr��l��"Od�1�Y%�:�R��N7�T9 B"O&�w�����*�^�<hG"O�%S�Kҋ���q��X1�\H9�"OI�A�E!+�񡴋͋q�Z	3�"O����ӽ\�ѻqjI#3�܌�"O��ٰ.W�xr�x���\�4}1�"O���iB�9��U�L�D��9j�"O5�v"ѽ5���� ,�2D�()�"O���/N�]��$)'�Ġ���Q"O"d�¡ߜZHx8A�.�F�R9AW"O��"�O� ���s�ګ!�Ԕ�"OTQ0�$�Y��JF�u�8Is"O�����Ϫ+^hQ�C�I���"O@I�Q�Z>N��V%[�e��EbQ"O1��ǌ�Ak���Ɔ?>���"O� �a��%hn,�B�I"���"OƄ�`�$y8�ԙ���S9���A"O��)� P,D�x ��F;�Ƞ`�"O�z�(V�b��#�(S|�P0�"O�*@�P(n� ��%Z6!���2�"O��Y�G���BEʇw\�|�p"O�cङ�$p���	�m
�K�"O��`Ë[z�Y�����.���"O�iB`�	V�@�pBa�3�̀�3"O&�P�Ǉ1���
T7e
6%�2"O�K3
D���y��ɳ�FD"O�9�cW�h�բ��U C���E"Ob ���9=±�c�ل|"O`��G�I>`i���R���{#"O���@�;_�V
�l�1�T}H�"Ox0�0�2}����&!Ŵ���F"On��2�B##+|8(�H�E���2"OTH�gE
D��m�7�ԻR���R"O�LJ����J1lZ�ud�"OPEbRK�"tU��]�EEr Z�"O�(ǈ��l����j]<0���"O����)H�ęF
�>�Ԁ!c"Or�KC���"5�Qj���ҍa�"O80P�M381F�3�8�Π�s"O�̱S�A���JY$h�b��"O:��aHɽ:�xLb1�W6o�)�V"OliA�;��A���!n�Ό�A"O�Q�W%�GP�,�7Ş]���c"O�Dy3m��2�xM9���詁�"O��KǡC9{�|!3bE1h2��"O�as��U�()zƀ�H��$JU"O�yj�$C�`׮��&-��"O:�q���&��"ޠ#���( �'�1O� ����6�T�˙'k���Qg"OR8��jk����c���Gt �0�"OL�2��L�lQ����5xe����"O���v��4(�@qx�η0Z��z�"O�9��&K���#�=#=�lЂ"O�pq�����+ k,���q!�$��`bX|#Ć�<_�)!CŞ�_m�}2���Zccߚ1����c�w�R�E(/D�L���A�����,O�6�pU�g�+D���w���h"H��F���o+2YY��6D�8"�-�:F�źb&��@���c�5LO��d	�'�'%��W�V�9��c�!�]'E4nԙ�$�-Lٰ��дj���M��(��8S'"_�Q耕�6���M@�9D��:�O@(�Vd�w�\����v�5D������+�l���Kݽyj�\�7$5�O��I��|\QAAD�Q�I��L���`C�I�^�Z�#��[�Xj�FC�	5 z�˥�̪=`�az�S09NB��Q�ƼPG=�v�(�
E=4B�	0k�df�Տ.�AS����zNC�	�a���A-	 L�M(�B�	 J! �kT�=Onu�ը�@�B䉜i��YYg�кp�La���$~(C�		!�����@�8wB0�r ��`C��Eˮ���N�0�
��5@
;xR�C�I4��jUd֑=���;���P��C�Ɉ����f�UhA�� ƅW����'�	�>�vD
$%�1���Q�.�G,~B�I"*7����F��P��2��
�C��7P!@I�a�8)6Ԥ��.�4A�C�I*�<�p΋�M
b��M�%ɢC�I�!'����ܮ|:��Xp��6�8B��7D�6���۩Ma��*���JYJC��(3�H�HcO�o������YB��gsh��'�थ���+y�B�	#0o�� �A7WI�E�"���D��C�I(K�D�B��Q%g�ɀ�J�	g0��h��p(��եL�L��؀B��'0D����k��T�l#�%W�|��P�C;D��a�t>&T��e3�a��.5D�X"uc��?Q~��S�qw&��^p�<��T>u�f��X��m�K�	V*l0��1D��ӆ�R�
��B�!,B��1��hO?��&����F ��A.�!��Bi!�Əo����A�C;g�$4H�Ywh!��_P۶\�W��E��21?HS�|"�x(�EO.��%�
v+T�3�L�	ϸ'�<#=%?�H�ڶ#�,�spd�0 Ԏ̣ե.D������/g"�D˥n�e�v<�#�1D�hh�*@�M:�,����P�(#�g0D�8ڴ�%���ٶ�K:z�F�أ�1D��BA��P(����F�T)/D�X�F'��\{B��p���Bܙf3D�(�i��$�{g#M�l�
3D�,q�fC�>���Վth�]�6b-D�4:p�^�iY��7W{����)D�\ԭK�X�u+�i�\pt`0��3D�,�-
�K(ā����h=N�W�-D��m�<��T8T@q��VD)D�P8b*
~��B�-y�JJ�*"D���uI�ު�{g�I�3� �`�&"D��0��U�/�Ex"�ǈ{���Ж�>D��ʷ�1mY*؂wFح=n%��� D�� h-��`�=d����0#�PS6"O6����I2�M�+��A��"O��z�FN�@ �"�m�<tﮑ�F"O�`�n�4��H���ֹ� �RG"O*��c"^8�Qq,I�� �$"O\	JP���%!��j+W'��L�P"O2$��;Z���Ћ֓ ��P�"O�1&�M&*����@� 1!"O�U#"���j�	G.k�ș!�"O�d{%�R�w��8�sct�"O������4b��v�ŤnRn�""O�ɪ�.�_����m� GX] "O��k5+O�i_�P�e��4,��"O��q�eE%�����e�,ol�YC�"O
�g�LZ�𺆆<o�d��"Oб�Q��' u94��)O�9�A"O�p)CDU�q`������0;�"O�1��>Z� �����a6&Y
�"O~m�3C^%���dUtyF��V"O�[B"N��L��$��r�93�"O �Ӕc��+���c�
��5�"O�2@eN�#���`Ç7��L��"O��[�C��Es���Vl�g� i��"O�Kb��$y>1PT�+_����"O�,1�HV"*�ʸ���҈@��A�E"O^0�.��j�ˇk�lg�I��"O���DN�\(�I�JR�+Pe��"O��-(D��X�Q&{�-8�"O�]9u�B�0�����]<:����q"O�X��
	'�h�wH̴?L���"O*���hN�N.��Ð�`/��qT"O\y�8({��;�$X�"O"u�t�M�9#�űx�  p"O��9&+¼}�ԑX��Nވir"O�eiVlN�)��<��d������"Ob�p���h��r����M�g"O,�a��<B�<`�������B"O8Q Ԥ�(���bC6X�B)�7"O|�6l�--��p�D�ܶ)�}f"O
��t�تSI�R#�� ��!���>������C��	�.��%�!�$��/��賃m���v0�%K_�L�!�d�k���Cf'�^�h��S(H��!��'ot��@ ޘg�
��5'�a{!��	9*j �JP)�-_�Ε�@f%_!���<|�Ha�fȡ?¾D3$���MM!���!t|A��(�0�T,"ę+$,!�$B!�4�I��ѺU��@C���N!��8$�z�zq��,O渨���3!�$�)Q�x��&��k/J��p��=xj!�$K�G�I23C�����IV� �KV!�䖻z�ָ��L:N�x�k�%r�!�D�M��ⴍQg���-�Q�!��V�ƥ�n[=ae�u"��@�C�!�$��$�-��F��bF&���D�x�!��,B�^-a�: H�9p�+|H!�d�[�zA�^TcRQ���C4!��>vm�!�ա[Gx���/!���3uM\)���#м͸���;^!�$6.���5D2G��С��_!򄌍5��1L��^���@�+L!򄃺V����2
�1RH\���Q
�!��A���j�圶f�*�붭f�!�d�Y��h�2���n�Ҁ[w��# �!�� ��`���QӼ5���_B���*O�Q#�ėh�N�v),�3�'l
l���x���yU����PyJ�'�F�AUDV=�Ș��V�nʹ��'ނx:�J�'R��u9�-�$}����'�����rz��%�P���a�'�N�h��E8u2� �R/��C�]��'a��*�O�,M��X��B�Cc^���'D¨{�#U�AB��Q�-A�x0�	�'ռ��Т�A�jL�Qi�
JO����'���:GI^,7�np��6H�J�3�'W��XON�n,�������>�&ٹ�'l��C!e
�"v�`肯�.�v6"O�IZ �\&�Ne��C�9d q�r*O ���U�{;�Y�&L� ,Ո�S�'�����̄Hq��0�@�	W���p
�'�M�#�[���qb�8&|��'�l�w,� J,RD�q`(<��'`��A��~ڌ �C���L�b�'�Ȅ`�|֮�A���@��'}8����I/��U����^z��
�'����]>Z���c��U�&Y>��
�'��`#-Q����&�=��'� �X
��m°��)u*� �'�2$�S�O���j����4�'ڤ�a%�1!|h8�iVo��dr	�'ݒ-pl��
�d�Yr�N�c�FY �'趈�0�֑W5�JcZA��'�,<��-�r�1v	�U�:���']��2���a�T�U�`��4��'�h� CJ�U��!�@S���h
�'� �bO�Ѵ�`�K�L  
�'!9�����8(jK��ٓ�X��'�����]���ɢH���Xh�'�t�����Q�j(3�l��}���
�'vi�tBO*��M�bW���PQ�'�����	�x�Re�T�Z7j� �
�'�N�����,�X������p����
�'�fXKaZ�@4DEᓇn�~0��"OH�a�#Ģyhp<���P�B����"O�XsFS+.�� :���jOD��P"O�8Z�7�(���C�f1�"O������n�BP����%(�Q�"O: Fh_8" �{cb��3�,ʡ"O����g�P;���!B-lU�]x�"O4����92��c'�8<�P�Yr"O �
et������P1���S"O���!!P�J�А�#Ȇ H�{4"O&��$>挃s  ��)�"O`8PЋ_17�d�!t�׾�>eF"O��c%��]������_��q��"ODdӅb��9������N$�� "Ox�J��W�ОH�! PZ�a�"O�Q�A+��K���1dY�V"O��Ɓ�9tn����ƾO��m��"OI�v��!���FMzH��"Oj`X�D�	hY��FXNJ��s"O>|�d�P>�h�W%^�B=h�"O��%#�����1%�V�#y2�"O���M˾r2���C-8r�"O��S��*Y����B_�#' ��"O�K߀}V�QFL9,?>��"O�X:+��_pAf�'+6XF"O�D�T��B�SPE��@
��s�"O� �%�RČ�jW�4�!D�p�$�2�"O*0��Y%v���C�P/G�e�T"OZ��%B	P�B ص!Q��G*O�	!E�O^z\��E��C"� ��'�B�t�n!EZ�H����'�*A	��� 0�����#�1����'��q�NB�$��@	ՃY�0�|��'�j�
b�ʳMiX ���.�ը
�'����@�O���"o2!���'���Y	D�7��leD/&Â��'��8�p�\�!ʴQ4�R�
�P���'L�����X0De6��T�~����'^&��sF9Oe�3�% A&��'�V��_� ?p��'�5�X�'��RC��E'�eP�g�*�.��
�'w��k�[�F�LE �^�nzpI
�'Y�ɲR���x���8o�9P	�'L�(�LS�KĒ͊Ua��7
h0	�'IR�Bb�S)��C$��Y�p*	�'J�$a#��^?J`I��z2�	�',�`
Z&G���i�c�m�
��	�'��e���G�NVܙڕ�R�bxdP	�'�t%ѣ����V�`��/]��mJ�'�$��e��VFDx`Uʇ�B���'���w�P��@;V�� KN�ti�'֤��%�MuJL��5ݔ@��k
�'��-Z��Į?��Ju�^�14��	�'�\�ѩ܅%-���o�9%\ u��'�:q���
	" a�#�43Hmq�'2x�d�?-m2C�
9�`)�'���Y⫓��ܠb��2͈H+�'�:+ �1�����GŨ�$qK�'���7�҃.8���_�q�Ȋ�'��1�sP�����&b�+g (���'��9��ׅK䈁���Rd�Ѐ
�'�c"�!Gz�L�UlI�O����	�'�ڡ�k5�NY4k
I憤��'隘RB⏡o��,�D�Ƨ:���'�0�!���
�4I��5:D����'%F�3��"�J�!��4UtY��'�dE��ET�+D�T!�>jk	�'���5�;bF��0�M(3��	�'D� Y����C�Tp"-ז2�8�'��!�CJ�:!z�x��U)�fp�
�'��� Mt�t��֢Ũ �P�'N����)�3 �Jɣ��D��'-^iǧ�Q$�RF(� ���x�'��	G���y�������
��'���!��Z�~QS��v���'�xL��ҽQS����Q�jN���'�N1�a�V�t(qe��f4�x�	�'p����.�""����X������'hDA�6!��0��6�ԧ��p0�'-L�@���W����  ����'^�T*���j��b��d�'J�m(UD�.e����WX.Z�x	�'3�bu ��y�V�~�����'I�܉6��9� ���A9.�N���'��@(�׃M&�T ߗ(�6��' 
���LN����&O
x\�"�'�"��Ϟ�InVȩP� �����'�z	���c8������B��P�'�񠑧�u��C-��?Z�`
�'DԘ��U,
@LB�2fn�
��� R� '�g�>`��
�� ��"Ot�z�ϑ�G�V�Ѱ��S�^�"O��X�X,���	7�� �p�"Op9�)��a`�!ч	("����"O�̓с�\W�`���"jj$)
P"O���El�9��Ţql	4fF�z�"O���E*[?�����F39X�1"O�����2h¶Al:� bD"O�\��٦A�2 r�3�T��"Odc#&�"�(����	�I����"O��H�!�N��8%�!d't���"Ova��΃?w���8|2�"O�f�1j�NPc4J jt�q"O�\�m�7z�p�Qo�]��"O^X)r+L�p�Rq�&��8S��1�1"O��RDC��G�ԡz��̶�ł�"O�lyG/��7�Z�Mݹ"꜀K�"OR��r�J3B\yy��J?�M�@"O��*�k�%���i��<��"O209D��1����j3����"O�+��]��܈R6�ɬ* ��d"O>���Yj��,��$M�-���S"OP�V�ðZHn$�Q���Հ�"O� �f�ڃF�(p��ܝ_�x���"OF�S�~�>A���H����"O24K
�R��,��6�Ax6"O��Be(��pȩ�SMPId�$y�"O��EgD�5�����v?� AT"O��:�k�>f��@D�>pa�"Ot�B�(X*���yI�BR��Y"O9фb�B�~�9��h�xٛ4"OҵC�;F"�7n�{�*A'"O���\*#^�m�C�G/jt��1"Oy��x�Y�v�5Gh�h"O������EG�̀�jÜB`8�ڤ"O�drd� z�.\Y6�q5"O
ЙJn4<iR���>���"O؅��n�^A�Q0X�l�0a"O؂R��$��  �n\��ݠ"O��`@���8At4��l��(
�"O�`X0�8sf<Ys��~K<��6"O��b6�	�bW�p�0�^�"1�)�D"O"�r�B��DNإ�5���8(��"OP0B,Bj#��Y@��D"O�a)�>H���2��~��+"OI�үϊW�8�!$�4Y��)��"Ol�p���5H�D!Se�Zk~�9�"O��4L6&O~�񗊊�=�TG"O8�x�C�:�eℯL�gQb��@"O$��qE�)I��b�C�"OPA8wl(Z.�#�� 2f��\#u"OI�P�ų4%�%��<�8���"O�A�"�ō7o��u�E�0�ę��"O	�d���(Q�6���ݶD�S"O�@�&�@�f����%���?�*�k�"O��ӱ� (dm��,��E��"O¹��Dv���򦕦%�z��A"O\%�vF�(/��Ѐ7#E�u�z��!"O���N�m��1ip"�7)V�k�"Oʀ.��q1SM�>L!��$���U`��d��xv-�(!�-G��y�)Ϧs��u�C9|����cM���y2Z18��,	�b��t�$]�ӊM�yr�]焥��%ߒ{,@*�"�1�y
� �x��:�]Y1.�2�h�S"O�y���\��AZu♚_�2i�"Ob=�A��`��6!�z�|YkV"O(u ��@�<G$�X5��10�rՑ7"O�m������-ʶ/F�^؆�bS"O���t=�Y��nհt�>AZ�"OB� -�rX�b�G��
�E"O�=I ��R�P��gM4��i"O�TuE�!mo�\
�L	�wT|`"O���D�V
/1*�i0�
@�=�"OV౔Ș�AqZ��⅒K�0�""Ov�B��*Fy>L�u���E�\��"O<�U8It�i#�ۻ("�\�T"O�2؎�_��2`�-���"O:�wFA�PEb�H���.��u�%"O`$���
����R�t� ]H�"OT�����5L���H�� �0U"O�<���E�]SJP��h��T�$m� "O�B�8��QI!�i�θR"OTQ��/=�R���U	7�¬W"O6�kP�Ai��RQ�ʢj��u��"O~y�sm�
%�z��������J�"O�l:Q�G�<
ȼ�S�Y��(��"O8Q�Wf[�5��`�p��u����"O���9_�*)ࠫ'S�uy�"Or�!�Aϴkm��K�q���c"O�9�M�V��	B�k�	wn�u�"O��X�f�yv��U*Q*AP�[s"O�0p̄{�Ż葷tiF�5"O"m�Q�ɭ.�N��e��GW��b�"O@����x��̫@B$�u"O�S���Q�&1�%K�&P5��G"O~����&
ހ}q��΍�\H��"O����.Q�c�!�ǒ����W"O6�������c(�?r���A"OR��P�	 x�2zC�ʤ05����"O6�#�I%Z���;% �>  �l��"Ol 2Fn��L1� A�ao`%i�"O0�CA���^�N��o��m=�Q!"O���GF^V�6Hs��
LI�Dc7"O��@�+�RH=	�`�/72�l9�"O8dX���O�|�놡��uL�""O扛�!�]�rT1��7�l�I�"O��b�F�m�JZW �0~H��%"OPQ⣮Ȃz�P����Ԟ@���f"O>��ψxa>��4��4��` a"O��{���#'։���%l�� 2"O�̙��*:��*���&h}�"OHD)�Qe�� ���[�4�<jt"O�V�)mR�ᐥ�Q~4I!"O��CC�N�M
*E1P(U�|�8a��"O���mڇoN2$h�'*f�x��D"OR��1�E9R��'È;�yD"OF	�f��I�|�YS��
�J��G"O����h�:TT�:���t��A3b"O�Z�ߌ6��uX�KӁM��1"O�Xy��:��@7�޽=��a�"O.y���٫c�>��7o�%�����"O����g�0!idl��֣4��|�"O,��Eԭ����$ݧH�6uh"OƄ8��Ոa98�)�MͻgT��T"O�eP�n�	#�xC3��4O�-�"O�JR�U1K\�5aت�Ҕ"O q�&�[�
��2-ҳ\��\(�"O� j-8��Ԙf��$QE�	D�ޔ@p"O(1 ���)X5�G�\����"O�I Wj	8L@d�bΡmOpK"O�e���ٜi�|a��D��r��Q"OT�)��"�"���M�4���8�"O����ҭg��� l�^e!��"OT����>C�݂p \pcl5z "OH��2	� ��9��"jƨ*�"O � G��O����#C�z9�"O��0$� {QD�)bH�-�&�Q!"O6t��M]�E��3�`1�2"O���M�*�݈�ܩw� i�F8D�8��!=1�$M
 ̕�-�+&�5D�|�Ɛ�K�f���	XXĨ�g/D��9AKĮ3�z3(��-�ā�g+D��p���p>5c�C��=�!�Dȧ:<L�W+�$z��(V�
/!��H�9	��֖!z�!Æ�.)!�D�����&JEC�|��Κ-]!��P�Urc�Z�iDt�Sr'�7�!�$�BTT�Z���o=��Q���s�!�	
��4#���\�����-�!���c1�X7ď�XڬZ����)!� )�,;��F,HUkTAV�
�!�$)vVx8��f�_L:��d/L�Kg!�d�%n�ʡ9''Z���+�)g!�dB8�p�E�{�����/Z3!���eaD�[�J�@a$�(	̽-%!��#�p��D#�"%0䋴�֕F!!�$��P�ꑘ��8#�؈���9U�!�$N�o���S�HV����A�;!��
&���:��I�5�ڹK�嘈'!��ҹ0�� ��	�2XSCKL�!�d��Z�Ty�j�d�X�0 ���V�!�$�x�|�yA-��D���E�_{!�E� H4{g#��n�f�+Q�!�D��n�H���L�;}k�m�E����!�d�?UN�Pg��\M(����Y#!��ڗ"�����.�����s!��&ud����Ǝ�E����v�O�5�!���s*�`���R1Q8��b.�.�!�d�	U�E��JW���s-۔K�!�A6V4T}�dܦiBNԒ��Ysi!�D��/>8K� ٬r��y#A���fM!�d�*at2P� @�7?i|�ئHؽc�!�D��cC:����
Q8�d`D���!�̦]���S�B#2��P� Q�!�$��d-���5��<�5E�nX!�d��H[���c2�9*�N.W�!��N��@�����r4r�#߸�!��%2�.���I6z��l�vCb�!�r�,m�q�_=>��T��U�V�!�D�+{FPe!	Q+�t=�g�εu!�D�1O����J>���:�*�Lm!�$�$��H�6lZ' �>�a�H�r`!�D6ْ����>8���֘I!��N�fW��T���>�2<�VL��o5!�䚐l�^��nX<e�,���Jψ5!�D��v�R�3�b\�2a�@׋Fw!��;.ιJ�)Ǽ4�6H�Cf�c�!�ĝGk�����co��9��R�a�!�IY0�%�`KwӜ���� %DC䉉c'���M�,�x!�3G�<O��B�	)} �\{DG���L�z�m
�^TB�)� �%�M��*<�)�9DN�: "Oڜ`��]�{��ؓ�� 9<.��"O�cK˻ry�<�6�bE�);u"O�(F�5}��rQ�K�H&2��"O�)S	5�*=Z�d�F1��4"OTH��D�:8bL8����YD��0�"Or �V��U`ؙ	R/�xU���"O���$�J��d���ŮBXU2�"O�q��L�&Y=��ӄ@�*8ld�"O��pׄ������ԋM+��Y""O,���,�&��%:�.�5W�<5"O��(�f�/\L�W�ńW$�"OZ8)�ՠ|�`�a��h��\ �"O���R�8Ω� �@�s�Bŋ�"Oh�Q��P�x�`D�}�� �"O����ț�	��Z �	~�$�k�"O0�0pӜ6pЙ��<Rą�0"O�Le��"]��h4�	�_�0�"O
���j1��
�gE-2P�"O��â�5Qt�y���T��W"O
�@�o�$���h$�.��j�"OPɪ@��1G͂��4�ʄ��"O~�(g��!BѴ��
��p�ۀ"OE�%��61��Ɏ��@59�"O@9�	<C6��1G�\3S��蓔"O" 	�OU3q�TI�;����P"Oʉ7$Ry�,��U�D��"O~}z1lZ�"~����)43*�5"O��R0�߫oN9�0%߳*d���"OFt�שհ=����cѸb �#3"OYA��0/}����Z8I�R"O� ��T?0<*��Gˎ�8��0�"O�,�$Ī(Eje��ʂ�6@0r"O4R����?�^Ahr �����"O^������A�.މn�\��a"ODR�8:���-V��f%� "Oڵi��E�4z
r�	D�
4��"O0��c��mvʴB����jʌq`"O�q��N�>�0OH��jt�"O<�d�±+���)��(�����"O
|���$۾1��%�d�lE��"OY`q&��%k>��#�/N��8�T"O�K�(�8Ѿ�[7�Sd���"O��HG��*$eDk5J��*>X�"O�	��+�3s��[¨[�-60���"Oy#���g��p鶧���8��"O1��Z"��@B�aC�/"L��"OP%#�ځ1V��Y��=���K#"O$�S����Q�q�_�CV�p�"O���7�B����@F�C��X�"Ot�@F�B%�XU��T�oݒ�"O�  ��JW�x\1�qXĀP"Ot�Ro�$W�*da�ㄤB��%�w"Oڈp'�J�j��) %t�X`1�"OtY2թV*Wt�ș1BƖslli�"O0#*_�Osf�� ��O��J'"OjE�"a^�e����W�s�!��"O�٤/[36���%�`��2�"Oƨ�#ʂ�+Z��ٱ
�i/n�"O��w	3����ɺn!�"O��P
A!,�v�Р��6!�dp"O� � 	x0H���	$D�e"O�]�2kӶ:?*y9�O���Qc�"OT�X"��>��
G"wЄ��"O� ��;W�ڿ:T��s�HB;MЀAd"O���-q���J�Όfì���'�0H��Jr�3��!Y�l�C�'>v�q@�W�Jh���\���0�'Xٹ����r���A�B�)�r��'�n���+�R��q��L�N�P�'_�D��Q�WOx��#�Dd��y�'�Рk��N*�E�2�ȳ;���	�'�8\ط��	h ��P��/G�ꀢ�'�6<�����~đ񧛆F���'b@��H�@�Q����G�l|��'��0З`�6�����A�H@��'���@(�*b�)�B�ê,�Z���'ZM�� 5��}��C n���
�'�F��-�m: #A�ތk��4[
�'����D��ڲ%� ���d�r�{�'�A�!�ٺZd�uh��+A�p��'�Z�]dN��6B�"�)�'.�!���L�
L��&NS�l��l��'C$�`d�\a��؀��N��U3�'3���hL2�5@0�� |���
�'�z��� �
���,�)���ʓ������
U ��$��-9�ȓ8ZE[����T�*   �>.�̈́�z����I>��c$I6 #���e0�U�q(�R�z��w��$��(�j��R'[�_���1ӡK�$�ȓD�t�iv�
g�i���Ϳ�B��ȓ'��2�W�$��� �ȿ{<\q��&��0�S�ء5>�%�g��:"�HՇȓ`�H�����H����GS4_@LՅȓ(XQ����d`�۲�h]�ȓ~Z�&�"fx[RϜ-����ȓ�����H,��F'�t�����td&����<,B�dK�1��&5�b�K�}�0�H#���^h��ȓ��h��Ѡ�21�oG�N�p ��qdJL[�� �t�S�&��犸�ȓl(�#LOݼ,(l�.3Aj���=�����8 x����)IpЅ�[�l�7H���V�p��+4~5��*T�n�~����["o_,�ȓXx��_7�j ڕGW��=��#%|���#E�8���斎uఄȓ6��P1H��[���ɶ�U�2&�-�����ӧ�-R��ˠ�t	�%�ȓV}����ݛY��|s���f��X�ȓo�$��L�9l5c%��!1��ćȓK.�A0'�(5���0� �9`���ȓ"��l��9;��p8V
 0.�*%�ȓ�إ��Nٚ*UT顷░/��ȓ{N%�� �4/�ly� �9�r��$ޜ�7jnA(I��1O���D¤}���'��EP��.*��y�ȓl���@��_t0 �bN�"m�ȓD#l�� �qF���ŏ6h���ȓ\��l�ª�4IvP��Ā�]���LZ�s�/ķh�&挌I��܄�%�T(Ӄ�*RN*deB]rxԄ�+�ʐ5(�;k��!%N��f������э?C�D8CeG|_����&|��r��R5?s�a
�@	�I&|�ȓ[$�%F���p�Ɲ�4�
a�ȓS�8`�藞'X� ��Z5(l�P��S�? �i �«'㌕x&!ߙ!��Pj""Ov!V���Й�Ҁ 4q�\�B"OZًUdP/�b{����wh8kc"O�	J�ƙ&B"2l����)W⩊P"O���Pl�3���;�H*6$�F"O\AJ"��f�@���#�*���"ON 3A�X0B��+�bQlߠH��"O*H�Ib�f@B���$?�b�I�"O$�#�%ڱE�z��qK-��}r�"O��)g��&�v3ri�!�41�"O0-�Q��# � ��1�M�K���"O�X���-�dibGf����-=D���BLJ<��(a�i���1-=D�xᒟ/o��)P%&!���U�.D�d�3�K��*�J���|�l1�E.D�dQ�
��!MB��H@�k>f	�eE8D�@����.���61�i3+D����M�Y��]�0��K��%D�j�A,cX�S��ژT���u%D�����=��Qڒ��_��`a�&D���Bb��9Ϫ-�$ ��!Ph��h7D���P@������R��7<rx���8D�̣bFV.wF�h���	q �)��6D�ؘU"��I����(�[��,Cpc1D�d��� :��l�ċG.%$�fK-D��#G� (xHه��o4��,,D��P�{Q�d2f傝s�Tq��f+D�PX!�/q�q�U9_)H�:tg4D�9�����`L�w��O�N��g%D����B��ԙ�`-�dmdõ
$D�d6䕍SK��@ @3���A�"D��P�[�g���xL��_�0Q�<D�8z�� +�|�v�]
r"
1��G'D�0� )�#**����n/���h��&D��jGk{����R�1+@�5 ��(D�Lԇ�(�����&��PJ1G<D���o�4pW�(�u�X�
��8�#;D�42��Q�J��f֜U:��O7D�Ȓ��������A��,��1�8D�D�Q ~U��A��|k0@T`7D�8ѱ�l< hq�@��A�SE5D�!�G�-_�" ��&1'<�=��F'D�����V tԂ���>Ԥq��.0D�c$nM��,Ds���3fyx���0D���f�1���Tj߾O�f�+.D�D{���5f���'�A�Tm���+D��8�"Z�4p�HǸQP��`B7D��3e��<+��kN�SĈ��d5D��(�� �Tx,E"̎A�$H��G2D�Tc�
G�d�¥	���Sb�O;D��c�.�j�(�lؽ^b\�D%;D��㚵N��$�ӊ�Hkf��P$D�p:'��&�R8⑫��Z@z<�F� D�Hi�͉� ��	�1��\��y%�)D�8�F[�9��E�&e��0F(D�;"OX:^�����-�)>,����K&D�hI�n�9���kˎI����%D��k��G;����
 u��iBP�-D�`Jg�i�
�J��j�΄y�E-D���ǃC� }���	DO���E�+D��y��gF`q�w�@V~�)��6D�������%M��M�t4	��]z!��;�^� ��u���!ʼ^_!�DL�s�f4*���+tcP9�rmӨS!�� Ni�!�A. ��sT
w�z� �"OPY���ª�0
�bԚc�<�` "O���C�(%Uܸc�]�|��1j�"O��k���~���`�Ab?0�
�"O�pc��@�{G0�/]>3\(��"O����Ә
��EQ"E9F\�5"O �0���6M������O��҂"O�� 6 
2���t��\��ba"Ob[`��'p�RI�B��*S�8=��"O
ݺ�*�j��E��X�$��0ӕ"OP��p��^�Ū3��5r� �[0"O~P���O�?|���GU��J�ǒE�<A���z�x)l�z���f��<f�C�g	�	AfkĽ|ڜ`I�
�{�<1��@:t��AQ�94�T)�L�w�<�^.��d���f�꼳���q�<AT�:uY+�LFb����j�<Q��$��\��L%d�2�s�"Z�<��D��ej��٠Q>�hS��l�<�w�2�
 Nm��V�j�<�����-y�\ږd\_1�Y�lL[�<��솕<^,��m��%TaF�]K�<���	H�ȲaK��iKh�҂Ga�<���_�qìbt�F�j��񐥱�!��V'�&;�L�	4�Er#`J�o8!�D�8"�
I�E����0-_ ]"!�!n�:9���-l�`d�nK� !��7qD��'�+�*��0�K�Y�!�y��9DB ����7�A��!�dϝ?�v$+́�6����Al�&Y�!�)7�4hF �*�֌�ҪǬt!�$�[}b�Ĝ�G�&MaR�8�!�D�k	�T��
"�B��ɽtS!�D+o^�Q3#jK S�h�!�N.I!�Ĕ ���#7A����}�ƏE/O�!�I z~5`�"������\��!�$M5Qε���.�G	֞�!�D׺vI�@ �#R�>�ۡ�ϡ*�!�D��j�8���NJ�m�z��F��`�!�dR7Q��$q/D"p�k� ]{�!��^fLi���ܲF����2��p!�$��GWPyq��1[� 8�ƠS!�S�Iȕr�A��~�@5sQ-�>O!�d͋0t�M����I�\Ȣ�ʪ<!�ˊjD�easj��HpaC/�A?!�8������Ύ{e*'_3?!�$�(B(���c��l,!g�}�!���/�6���)]�H¦L�!���ky:��!�('�=�CѦ=
!�'P����́�bs���!:eN!�d� 7Z��;CB�L�f�����>!�0g� ���Ǔ�:\u�F��&!� uk��@�ՖR���3��_� �!�$�,�L@k&��D^H�͋�f�!�D��o���m�^aZи"A�S�!���.�U �!߲4(ȼ:b�ɇy!򤅆Q�0r�bY�8��`�&��+b!�7�ŨAaZ7S�РZ����N!��B�v ���F�%4�i�/�?(=!�D{�<y��I<"Ѻ��g�n!�䖉@/du  �mb�(J4��N!�Dٓ3��PV�ӵw]\I�е|���'�f�Ja�?\�N�[V#6TL��'���p���:RY��o3��0	��� p�K��ɒA�z�ENL��`(��"OE����*�h���SU���b"O�8�Ƃ	Ԡ=J�B�
o>,�"Oh �0K4?֍ِbσ-;� �b"O�c@a�Qߴh u�Q.G��11"OPU�'f�=;|r��T�j�`2"O|��N�Q��j�$�'9��e�"O���悟�<���B�@�_�<�{�"O`��SNU4KLJF�öo��$��"Oƕ
'�;^�8c�єx���&"O
��1HCk/�DX�-X�G���@�"O؝P��Z��у#��><`)�"O�x��%Ȧ1�d"t$H	hش �a"O ���!�|U�f�Y�y�\�w"O��"� #)=V��p�V(jhv�S"O��F-�7l\��H�=��ݘ�"O ��5.�%��B�%_�|}��A"O�i
3�߰q�ڤ�!d�9j��?�y�mXd	I"M����
S+��yR��<^�)�@�(=����y�9�L��Տ�?kr!⑆�(�y� H7B��HV�+CT
����  �y��Dh���{e��>b�i�sb$�y��"����Y�6T�+�%���y�H$\\��ui��y,�Y�g�-�yb%��w�^|��j�xY�=S`ႁ�y҂E�_l�ZB�D\�v0*p��*�y��ӍaV�#C�'�:쁔g���yb(�9B㚱 ��2&���rBW��y�ܹXr�P�A?��0Bh�7�y�"C'��Ȕ�~���s�?�yRֻT�n�d�@�z�F�k�n]��y�/�Q�\��R��G04��bZ�y"�	I�Y�2g%D�չ�nF1�yBo��c���+6��/ 4�b����ybOT�s��\�@��n$�y��Ug�����3��8����y�dYӶ����5�xY�e�*�y� �*ӂ��ǌ]&1���qF(��y"�Խq3-� �ځz�Y�Ę-�yR��1��<���SkΤ9 ছ+�y��'DJ��q#؏k�yzg̜��y"��9��	���2!V!tDV��y"��g�0�s��7�Zı�̃��y�.�|�(� �"�>Z�H� �T(�y����8k�TP@�g�n�K����yR��HxL��A;g�D3���yR�<	F֭��JƣK�@��"C��y&Գ?�h��kT#p.^�RB����y�<i��0`�gֽ|�R 9�䐺�y�ݖ޶�q"J>���(#F�8�y�\fw"UCA�'�������yB�aKf(�L,9vL��m�yb �;dl�R`� �|{�bM��yRJA�	Q�|��[�EJ��j��
��y�@�zڐA��ɚ$2��قѡ���y2ꐫW�9ASI�(�y1`&�yrk�'5b<Ѐ����%GX�PdԾ�yB�חM�ҵ�áy\HH3Ɋ��yR�O����.ԼC#r]����y���|[��!���-�N����<�yb-��� � �t�����h��y≟�'H��1�S�l\�p�Rg���y$
"|(�@om���/��y
� ^M���)G�x)0w͘����"Or`�@⺌��O�V����"O ����F)�`��G�g°��b"O
đF�	�Ng�����^)5Lj��6"O�´,��Zw��L=j�o|�<yQ�7P�ՐS+W$����`JN�<���
&1,ԫ�( V��G�G�<�L��m��%F�4Kg��<� T�V��|qV�6.l�+�b�z�<)��G�;�
�[ӥک °�9�c(D�Ļ�Io�H���:���` 'D�$�Vd�����To��X�~%i�j?D��jQ$̔����hΠ;�͐��9D��K�l�<D<�ʇe��D�6D�LZ�G��2�|��e�Z�W��� 3D��C4n:~h$}���˗|�Ƥp�O>D�� ��X�܀�S��7(�����<D��Ye��1����rh�Hx��&;D� �'N�K�ܐĊ��@�v��u4D�(æ�\;E=�	P�
�'FX=y3�7D�x�`�W2����cʉ>��*��'D��0��w�X��)>�ɲd%D�x��� \yz�"	6I��|��5D��dM� �UP�ҭ�L����
�y�%H, �"u��¾8����Ď�	�yR�\=~�ш��FZ ��	��y���I"��3��ݺB+x����5�y�Ʉ8u�ĵ��ʲ6YT�!Ņ�-�y��$p�� 6�G�+
��H�Q��yb��"}�5-��s�:����#�y��Z�vi>2�ʔ�p��ir�\'�y҃R�R�eM�#\fv��&�
5�y2G]1�tB��@3K��\���ƌ�y�MC#V��h�ʦ=?Ј������yB�U�z�8�KV�i�r�҉�y��͟t9�}��^�="��h�oV4�yb�Sxa��Q�� =1GD��T�Z��yBo�� 7�P��J�$f�ZUhҩ�yR��1!~�3�W��6,$���yr�ݺ,�6, � �&8{����y"h��]���Zt�ƣ�֬��Ë.�yr M�fg�I3P��2�3Ѓ���y�i[�r�0�oϻ<�^ 17�8�y�oho8�D���.a0R����y2�J�4��p�%�T(ʗN�1�y2lM4R��u��^'",v؁f��y�@�cM �`IΓL�	K$�y��@-X�s�g��+;H2u�D��y"m���T)�"B�Y�jdXt-[��yr��4�~5��PYj��c���y�iF'm!(�آ͚�@
���͚�y��Ҟw� ��cKS83����@���y�K�K>ֵ�G �99X�hv�]��yr�,L�2a��i�5/Fĸ����5�y�cL�W�AH��,,���ŮJ��y��P�p1jQ{`�[,*	f���NB��y�#<%���# ]�nR@�2�K�y�l7 V�)WÑ/(�|�/]��y"�ؼ�*�;Ca�\��+�����yr&�d��������Z����y��:��!X��(Bj�$r�M
3�y��C�;|.��%�l������y�f�6TGr��,G�yԬx�N�y��@��@���Ei��
d� �y
� >-bፒ��09�L��~v>�SG"O��HTO�;)H���d��Yy�Q��"O�A��CD�(К�8���Lr� "O|D�b��%z�����8� �+P"O�8sr�B<f(��x�g�{�L���"Oj�� MP�<��'��>6�8\� "O�<�c���xD��S"C��|y�@��"O�I�ϒ+Q�*\`'aN':_p-K"Ov9`��R�1]�,hQ���l��U "O�CB��kU$ٵ��.R��'"Oh�闊E�y�Ɂ�g�T���"Oư*5�0ᄼh��܂Y��+"OB���HF�2j�.Ak�|���"O�����:I�\�t�To��� "O$�'N/&�$8����BI�g"O�*2G�7W���r�j�=�0my�"O�M�p�[T����×%?����"O:�b֠�+}N�l
`HA�@�M�"On�J��C�B��5۴A�|�NP W"OH�a5�}D�`�K]�`����v"Ou��'��z�F@3R*ΛO�*��"O�8�%F@�l��t.
�/��uW"O��Q�ćF캗��>��q3"O�{��Z�1�@�E�C�αB�"O$Iy)�#%B�Hwˊ�b1kg"O�p�AƼ8:n0Jw*[�'��q�"O���&Ϣsΐsc�:�K#"O|��AW��bQlx5��"Od��N/3րz�A�c����"O�q��BN��k0O�5j`4Z�"O�Y��A�l�^�򤎖9dT�R�"OtQ���@��:� �[�1�E"O4\q�)p  ��!��,=V@	�"O�Ia��ЋdE�tdߎm�h�8�"O�a�BB˴ 1N qg�G�@��Q�"O��)釂6������gG�Y�"OH�a����ه%�3�F�m�,B䉴�P����ޓN�E��o�& B�'E{�����K�	�B,ܻA��C�ɈHm�$�9w�#Q��a��C�7��2e䁕ư�P�
V5g�C䉧�XA�tl ����a�q�C�	m�>��W0�����ԉu~<B�	�L��	��_� 8�1@T���B��C��0i�H����%�dX��D�
�C�I�
U�ˢD�/^�^X{�`�SR�C�I�RL0��O<V��eU.��p�\B�Ɏ+��k���j�6E@@bőg�B�I=g�"d��h��i"�QFOF0��B䉆t8�
E`�bw��He� �\�jC�I"
8`��υ7���ڠH��+�C�;hG,uy$	O�l���o�e�\C䉦4�EH�h^�A�AF:�B�ɐ������Vx��v��9?�C�I7����Q'>5�$1�#c@'u�B�	Dv� ��<-N��� �jY�C��(dS��o�K��y�/�t�C�	�q@��R��<0s����-g�C�ɧF��@��˓R���)UM�=��C䉱P�\��ѷ7�fM�-̑s��C��31��[*m���(�rC�I�[�1��c����Ce�,C�	>�F��S/U�i��!���&��C�	�$ox$�d�"lάHF�D�!��C�)� �10�`R�x��Q۶g���S"O�{�Ȉ8�J�Z�A��T��	�g"O��H�ӏcr��p���m޺���"OPHAq�WG�� w��Fي8��"O��#�)V.Aرo�B�x��"O(j.v�0-P����k��#7"OxU3�/�){dyc����)�b"O\�gBF1ݐ��� K���Ti"OPp�� ��<�@�[*�csz�:�"Oz�R�G�
m;|M���[2J��Ƀ"O@ȱ�J^�}��qq��/X�ȃ"O��:��[g����F�7)�ʠXS"O����*@"y�$'�'�m*�"O�ԡgG<IE��d%ԁY||�ٰ"OFm�C�#$m2<2ծ
:q&ȡ"O$��FKT.T-�J��ǰUp�p;R"O*��b��Y��վ<^� +b"O�1*���% `6��2-�""ON4�0ECq
u@B�W�!�>}B�"O����Lޠn��А"�����}Y�"O\(�GML�j�:���IтW�8���"OR���d1U���[�!FEZ"O����X=C��;A��S�y�"O��lE#fz��IR]��	zF"O�4!t���r������Q} �� "O�<`�%M���BD\D<y�"O���N�0NK��� ��/LUI�"O
$��BK���u��"�ͨ"O���f��lW���,O@����"O<�!7gV�B��!A�C?.�Z!��"O�9���Q/yz6�ص�V�4��	��"O&9sO�y3�x�qΌw��0D"O (��M/u�`R#��0q�AF"O�Q�SmI��q�L��?�^I�Q"OF��LEL�\�KT����	!"O�-R�J$���&�{EĹ��"O�q�`%כO�>�sR���>(&���"O��I�	ɳt� �Q��K�'zi	�"Oj��EbZ����v��	T�*!�"O������a��p4���h��T"O24C�σe����d��L\RA"O�a
6l�*�����Gn�H�2"O$��q�9  P������]}����"O����-|�hy� sjD���"O�7�I�m!L���hA�9��H�"O����ӨQ8EAF/|�4�;R"O6�8-�EE001�&҅ =��!$"O�� ��,R�x�zq�'h��0"O�]	�
�D�l!R'��x
Y��"O�, ��'�4	� !�*p�"O���3�Ѫ4 ��A��2X��z@"O<�Q��q��Yّ�ʝpnhD+�"ODU�C$O-$�b�U�օ4g���"O.u�Ǫ�:�fXďhZ���"O����T�%5Xt�q�� N��"OޘөF�.����!�;��J�"O���oQ�9�цkǠg���"O���J��V������	{U�M�"O�h��nжj�(��
Q�K:f�J6"O�"�I�p���C�ʗ�?��{�"O4�s�,�3����vv�"�"O�d1�W�,�z��/$u�"O�P[u-
T��*�`0 �"O@���@.
�� ����R"O�  �³�Fk��F��`���;6"O�8��'y����եT<k��P��"O�Ȗo�� ���k�䁅n�p��"Ob@��EJ�n���4�U�C�8�
�"Ox�b7��D�|8����"d����#"O|��B�$fr5��E	+z����"O���������N	�	��+�"O*]���������R:��څ"O�EdN"�D-9@�Ya�N̓�"Ojp�fN�D$�D��8W7� 1f"O���CW�z;�tr��C/��ZC"O4��S�ܱ]zZ�f��;"I<L%"O��s�H�Nq�K�M8�Y�O���7m�I�D�J��& �@^C�<Q��s��!�E��#{:1S@��e�<en�%6��i�'������J)|�<Ye���vn�I	ņ[�Z(��ץK��hO?�{;�0i�EJ�dgBQqf��rF�C�	�,�r���X	)x��S�T��RC�IG�~uj��=*9~�
`'��b�b���/��$��E�d� }	f5���0!򄆭�YQ7!�	<��|7:kYax��I'[�4<9E��g�ҙ煌R�\C�I�1�tdq�ʗT"��8`!O�"�^����Y�L�"�b52�ʃ9q.L@�"O��vNU$a��k�i��>XFᐧ"OޥTi��2���R�H_$oF�d�G"O `��@����7�Y�a�NIR"O�@ê[��d�1���S��u���	�0|Jb�	h�輐ш�D������s�<I&N˂A�q�T]�raD��V����>�G��2��9�n�IT�ARA��O�<�E� -_������Q8��2�r�d/�S��)�JUy��w�Yx橑�\�0��V��0���<:p�˰�e�ra�ȓ+t0�"���� �3g!�D��4�ȓF=���1��0W�vM��#�2v��-q�'/Э�jҠ;��4��N(_�t\����)�t���2S�A���	?N6H̹E���Px�iK��Xա�4kxcT
^�jD~�"�'_J�K6��6i
����G a~|��.���3U^F�J���>����U�C�I�Z�]��c$��REeQ(=�#>a���[J@��WeH+$��-���
K�!��O��	RU��:��9�ǆ��i��z��%�/�.ypvl�>2~��#�UN;tB�ɮ4f��2EG�K;L=�-��O�>x�ƓfU�䛒/�d�nY
��X�T���� �M��y��ӊ ' %��+�s�b�3�b̉�yR�*bQs7M�;6�\x��b�
�0<���$��H�TlK�a\fxT$��y~!�J�$���b���)$���5� �HaxB�ɵr(e��J�Y�x��ݖt�"C�I�aIQ!o��v�B�X���1;F C�8AV�b1���Mml���hs��B䉫{����@M/��H�Ն�+C-*�D�>y�Z��%>���~��˴A�z	����+ �|��n ߰?��'�*<0�Mnľ�ᇪ�4H��q����M�'�%,O5i��4i(�a�{��!q�ə&�Q?y�@,\�f���GLX��� �#�O��eX^xkQf�&HT�#�c$Lh�m���y?q��d�~څMV�%kv�' T�g��i�Vd�@�'�"�i�Q>���c�FXj�C��<}2ŠcM ��-�O8xPP��/*� 0h�M3^d�b�'W�������j� x��oخt�l*��D0t��F"O�u�IMJ/ք8q.��z5TQ��xB�{��hO"��1���zJ��y���M�M B"O�]�i̖E+`i�Ul,);�|�>Ƀ˄Xwp��)g��'Πl�Gi&;@���J6�v�ד!̶�O0��@bQ�p��dbU�S��+��. ���DǕ�C2A
L�fg��60F���O����#K�S;�ybf%�#^n4mK(<iu��a�6욵Q�}�@�s�
�M��8k�{��\�d�0��g�>�`��C�yBʚ�T���۷�`�C��=��'ў�Oܼ���,?fx�3c
]�:�r�#��HO8��dg�1`�����a˔���i��$���L�p��aF�+�넠*�!�Ě-G�z���7)�YIlms�C䉮lv-���!�8@H���v1�C�<�d���G=�$٥�Z$*�B�	�nL�s���4��$2p�2o��C�ɏH��U �p
��"��$xpC�Iv��h �7/&�<r6F`C��N��PR�׋ko|�Z���+l�8C䉇`Vީ0D��#2�Vt��$�OF:B�ɥ}O�[s��W��\��A!n�C�漴�K7_ζ��@K����C�I�N���'�Y�0���*�C��M=��� L*6-NAٕDF�x�C�I�p��ݙ��F, 	baä0I�B��4����� B ��"����dB�	���Uj� �U <1: _P~C�	���p��W,&� =`���) �xC�I?���$��\ �f��`;:C䉵s��4A͝x4���ŏknC�	IԪ����O��"l���C! �B��$@��mѮ5ȍ�����B�I�� ;%#L��Y�g ,]"B�	C�b��� ��(@]:  )(�BC䉗;��`�V
�H^y��@�%vB�I$ks@`��R�y`�(�ڋoC�C��,w3�u	��r�x�HvMV�(܊C�IJߎ��h�$f�\Hd��YVC�ə=j�4�f�
����$�ҭB�@C��5Qi�d�pC7u:�f���E�C�	�|�P��ҙe�9h��	"��C�IE�<���"V�,��0��A�>B�I�YC��p���"����p\x�B䉞O��nP0�F��S�D�B�ɻ8ĉ�e��h1Vp�B-i�C�
��yQ�F�/�j�*��x��C�	-}�<��j��P>$D�s�:"��C��6�dDUm�<M�d�6��2W^C䉯iT�l{1�׾RH o;yRC�ɛ;�B�0E��~�^e[SLÈw�C�ɛˠ)���$�PA�p*���B�	�mx�����s�6티� \�C�ɟC�B��𾐊wh�UW�!HW	0T���6��h�V��ĆAZ�t��"OFt��G�9:l�1�q�۰W�jA�G"O� �f��*���y��Y���bA"O�T���\!����#Js��"O�P�%��8�`�P�-k��)f"O�	QBG^���Q!�Y�Rr���1"O�!8�\�?��Q��\�)]b̢"O:�8�Ȏ:#[F
3��<JW��*�"O��3��2���K�,�� ��P"O� �-�#\-��(�F߀P�t<��"O��x��\+�8UJ�&��+�"�"O��I^'p�d�[�E\�Sp��ht"O�m��$��	����D�IV���"O�A�ԡ���<śdٞ7���Z�"OX��ѪڻTհ9�@+@�R�,I�`"Of�a�ĝ�)cR��q���!�h�%"O@����*N��)���3H�6 ڔ"O��
�KL�b�\\:@���~��X�"O�X����iC�в4�G�!��D�p"O]cNi��9[��ٴ{�1qc"O�4�Gk,�|H�eM"�B8��"O*� U�ð`��)�����#k����"O�(�gViȮ|����Ji�ԑ"O�	�� ��g�}�P�B9Kr�$"OV1��U�Y�	��`�k���@"O=�`�6B�,�F�-��=��"O� ��a)��1+�m��\�a"OVU8u˜\?܁�u��}�h��"O|!�1嗆ʦ���B��\p��"Oj}��CJ62@~�{�a@�T�p�"O�Tj�Ė���ړ���PDR"O�Q+6��?�|�2�#
�X�H��"O��9�*ݑ2I���!��B��9�S"OUf�{$�L���9��;�"O����*η'���aUKݾc�$U"O�ѳ�/k�=[��@�"�:ݠw"OX�RE�җB�t5��˙"2�]��"Ǒb#�ۢK�A��K:X~�Q�G"OR�낄Ƈ$2���ұn~T`��"O@0C�	�|b���i��hvU�"O�Q(T���}��X��Z�[��a�"O@ڵOG.~g,�yҰt�\x*a"Or�s�욁nz`�Q k��`��a%"O8HYb�۝KF՘��ظ;�,��"O4���lã�E�#��f���"O�:�ǋ�8���5u��r�"O0s��=,\h$��+��7�2#"O�ի%�!��ajS��=)lLp"O�x0�޺pAr��BO%o=��@�"O�a���E����'.�U��@�`"O88iA �$��\˳mS�F-$`�"O�!s���&T�u����t�C��+�x�u�C7n7<�(֎�C�I�y�"���Ņ:�.	�c��>X~C�8�|E��R�j�:��͏-C$C��q��8���ō&�{q��J�C䉊,�ĩ"$��[/�؉�-֓L
�B�I�z1�`��)�p�r���CE�C�ɵ]e���{���6�׾C�	�oo������T�P�4�Z(T8�C�	�"���+e/��1%�԰Gi�%D��C�ɝ�vP���C��-`df�uͬC��h �<!��M6�d��eŉBB�ɂE���C��Qиx(�%ЌYB�I���j�"=Xz��� ��C䉵m��Ѕʃ�Lj���0W�B��1�ʥ����g��$��>nRB�I��Z(�7�]�K��T�`��i��C��W�
%�b,�9��"f!�!V.B�ɦAh��@�(3_*�BQm� B�I�WZ-z���4�PP�WP�b��C䉬)��k2dP�6c�ka/�&I}nC�	:��e�ᅛ�L��a(�"͑d0�B�)� 2�!VB��,��ճ��إw�V�+�"O`iP�BV��(<��+���e"O:JCKK�?�8�b*U�}� t�"O�`1��'����c(]FH����"O�ɘ�-û:<����'I���Q8"O��@&��x$X�q-�=,q�KP"O4]�"*Xݠ��V�@�SY<�C"O���
K����I��nMx���"O.-Su�G*B+j=�P!D� I6��'"OT]B��40��U�G�P�k=�`aW"O} S�̪O>p�B+�Q.��"F"Or��2�D6E̺y��C����A�"O�|C�.�2#f<�`�E��rlw"OH�@gڛ<��d �
��zǮ�r"O�4cI���� �*]�F���"O����u�bA�j�g4��W"O6c�N_0�\�R�Ϯ:��M��"Or�E�,dH�ƈ/�� iP"O�Ѡd@��4�F�U Q"�#@"O��;p $eWJ@��+�H�Q8�"Oиc4�ÙcN�	r*�5R%�Y��"O��#H�6i�Z<���֩;C�$ؕ"OlT&��!�V�BiĹD,�Z7"O�D�C�//�l�*p��/��9�"O2}(��(TY�5j�ŉ��R�"OX��D�SA��B*lx۱�$;�$;�'/r��"��L�O����Xo��a�ȓ V��#��p.�����]wH��Rb���4�ɫ2i�H*��̈́ȓW���XR�`��Y���s��Ʉȓ��U�V��=x����Z�g�($�����.ҬH�����
m�Іȓp�Pd�C����D�Q���ȓ;��Tص�?�(�S ��ec ��ȓޔ3������G!�d��ȓ!��@�E�Y$?�Zm�K	 !o)�ȓq��q�S��$`<)"K�SkU��)��9X��@�&%��c���4C��Є�d� �X���;b���rۯ��@$����I����o���\��e�i� (�ȓ)��tK��2%�r��W�*	�����O���O���󒅑q9�Ԡd�|R�)�SJ�^QI�H�����
�%U�C�	�4E��A$��P'|T�"ON���
2���x�k��o
́��'sў�Z��: P ��OT�#�Qs�L5D����K9X��U�-����)7D��ǯU�SF܌0�Ǖ8��5�9D�p�E��l����#Hv��9D���d	�
����/ĕ������"D��Ӥǈ�^��{��]!�p�ٗ�>�	m��ħxy�`	�-c*��%��.x�.	��X���rD��D?���F�r�v���M9�#�_�h��uP����KRPF{r�O��� t�,bXQ� �^����'4t@R�R�?��xI��F E]� ��'�,p��R�)�l�qP�E�~l��'�و \ |H�	�GgY���0!K>1�'4qOq�n�[0��9uv�m����4ܜ�
p"O�)�Acb��ȍ�cl�2� D������cVi8"C��%�b4Ȥ!D�V�^���X�� �<�8�2�*,D�|c�A!U?����^�y9ق�k�����+��1�cD�J�����	��C�)� (���՗l�Q{wF�t�t�V"O�T�5#΅��@c�ꟹ�v�0�"O����y��D����u����R"Od��F��� �vhX����b)�S��?��iQ>[zL��ό/9�8��t�R�~"�'5`U3V�Q�z���0Sl��w���x�����ofyqm(2��z$���0>�K>1ԇӂJ�Xh�!G�3m�\T#ZJyr�'7�H�i�\6��q%�#<�1���hO�h�r�	�W�&��� +)�,p0�i-��dD%�[�H�(�Z�C�S=!��0�9� �a��E"կ.t��
O�-��@ωA��u��^�\�*uK�"ODX�ӁP
V8���$P��9�"O�`Y#�ͪ
4]�ǧH�� A�"OΕ����Bok�<UZ�I2"O\`�e�<!����%�+,���b�"O>\��nC��=R�V%���A�"O��2�M��Ā,��.a��홑"O��*6�A�[�D�r�^',�jH��'��O�(I�(
�}��]�6�]�sɼ�@"Onp�ņ��QA&����,Ģ�I`"O
M`��*)T�&��2"BM��"O��&l�*���	��Ѱ,ν˅"O�I��Ɯ�����dْ��A�E"O6l�P(�*d^��
F�O�� Q�"O���.	�BT�q;��ސ!�z�w"O�@ � 5e	@E9�� �H	8�*Od�0֤[n�L�W �>i��2�'�F���!� ܮ4���2f����'j(x��F�����4$8�C�'��2��Nh��Z�^��A��'Y�����&�r��(��^F��(�'�����'��'���BӌєL�Z%b
�'�t��1�CR�D�I�
98�'�`��c�W�,���DL�������'��eʄ���y%^-���zF ��'��I���,*JQ���Q�w��is�'q����\�n~����X�|�	�')v	��O�C*�T�DA�2M�0��'҄�bG� �0��9�+ɛ=��=��'^�Y�X ^~���Í�-��U�
�'��-��Oexv5��d��&�:]I
�'����U"�����lO`��'��
1Ņ\�l�bX�f�\��
�'61�c�\�UHn����.R},Q�'������}�aS��?B�Ra�	�'l%���UӴň$�V�:��-0	�'�:�Q(	a�t�sK� aDށ��']t	� �٤T���s�U\rԱ
�'N�|���"6	�o͜Xڸ,��'��i�݃=DY�b�C9X�h�'׸H�"��*Cfr�48���9	�'I>ܸqB��4 ���1��&����'��{N�#@����Ȓ ��h{�'C�}S#�ۖ�䫵υ'�@2�'����+�400�õA�Z(k�'r�L�`�C�bE��8ROZK����'@��G� ,��`a�E.@/�<��'^�"��S#NsHH�N�8p )��'�P!J�4b����D�$J�'�����´Y�l�ם?���'GX5�WƎ,.d&=P��4K���)�'*䌙�%6�&�Y�-�F����� �$�W��v8�P)��&R)�"Om��O�p�L���k�##O�})S"O`�����vmR����ÖCD���"O\�jW�O�tdL�h�"�%��qq"Or�&jͫl@I:�ɘ~ژS"OV��<})�4�,�1|��	&"OUJq�O�9x���M�=i�"���"O�Z�k��Jޖ@�eɜd����C"O�<�� S29uf���G�xD�B"O � �t*.$9�a�~.��V"O<������<$�Qf[�
_(��"O���"'�{ɘ�;s%�)R�V�'"OH	��V"�>e9�i )s�"l�w"O�m�T��Tf�kwȀ�W\�Cb"O���)�j�����gSB�y@�"O:tÃ��IiN1i���:}�&!Y�"Olx�"�(|�1��ҋ]]^�a�"OȽ�%]S��� �CI$��"O��p��ծ����1b�oFj��%"O84C�
��"���:3� 1�,}�"O�9î[�b�� -D0������yr��1$�z,��A���q��b�.�y�h�j�=ʧ���%#U-���y�gN����X�>��Hd�N��y�S�Zf�$��T&l014�
7�y ��N�rggY�@�� S�yB�Ш �4KP��wW$@"����y�O��k�����[5i1��
����y�L˾{�x̘�NT�:I����y�#/�Vh:��T��*Qc5����y��%qp�����/"ql�Y�+�yB-7s.��/�|^
G
�yY+�
86��J���5ߤ�y�m���\ 'Ö���\�4o��yr�� ]���jG�eTk�
��y���K�l p���{ TY���R�y���3%��i$�J�(D`,Q0�	�y��^�:��E��͜O��C�� �yr�>��ܸ���(:��zF�ݡ�y����9�ށɅ�b&��0���y�AŻd�L�3�M�Y,��8P��,�y�A� �|�p��AΊ�)��R�y�Ã�]Պ�`��*1��
��D$�y2����42!@ߧ>���W/��y�,���(*#g��5����(�yb�ԯSe$l��hB�:B ���G�y���8 6)sb&
�hyl��$A*�yb��;"��'�b��H2t�݌Ǹ'k:%B��t����8v,L>��^�O�(@h@��-X�d�A���I�<�@�%f�,���ue^(���Mi�<6S ,�mi@M@�IG��k�<���	�=e��ǃ;>����P�����V�HU�)#��<[����D�� ��"B >[��J� �|��n:� Q��3W������;O@.���ɀ��a�����HY2Y�B��ȓ�F��0��z��!�JȰ?X4�ȓ'oܕ#�*H�y,����'��g��m�ȓ\%)��'B#@ƖY!
A��ȓ)=6�*kǄl]�]��aC�
h�]�ȓ8�|Sਕ�;�5Ȑe،�� ���ŧ���uY�
"�*h�ȓRZ�p4m�%b ��O[g5D���O��&�I��>�6ǀA{�Յ�S�? �\�;�<�Q�F>-�y�'"O�53$�(�)f��4�y��UB��6�����i�% ��ȓ^��ٓ��q�p@����-�v���J�h,�E-�H���+Q;@��f��)�F-��jζ���χ�m�m��E�f�A� R��lzt��X�D���ڼ� t���4T2��ۺr:��K��!��:a��)���¶/=R��ȓ}vT|�b�I4g��AV	I�d���q����D�ɴD��b�B�*~���Q�Ik%�³:�|�h[>x���ȓ
V�f���06��` �-o�$؄����JG�I�E��e���Rm
~��ȓx�`�m^+6��pIdk�'i�@��3D�X�6^����"@�8�ч�q]��뵏�*��
`͟��(��ȓ_�|���ȁH�P��S$/=���k�u1���(�<#����X��/3�œ��a�XS'�b�� -�P��N^"5�*��cLX�k�`x�ȓnÎ� ��c�ȣbbK>��Ņȓf<43K�[���p�˅C:���eZ�;������ӡ'�	s��ȓ%rJma��:��1"�P�Zp��c��#6iO�6�Ƥ�.%��B�+�hA*�(߰W����3�?aynB䉲/��85ɕ>l%�\r�o�[JB䉙K�z���H/NΈ�Q�z^B�	xH�-�Ɵ�F;ɑ!�!dB䉳D��D��޾n��  ��M�n`B��!׮ep�Q�'������
�C�ɊYf�|:5�='���+�NơS�C�	&x� %e�6Y�(2��y��C�ɒ Ov��LW�O��e�ѭ ��C��%0�(�cC�#H�q��N���C�ɪ)f����9gW,a	v&�-n*C��6�6#���"���'`@-.��B䉂\a�|ꔃ�0o�f�y��O�C䉳7V�ӳh�z6R4�Eϛ�[MC䉞d��t1S��$*}�c�h����	�3�H���'�*�c3Ƒ�h���d��5��5`��(0��`��n\��Պ ��� =.�:����O�nZ!���;(��	��J1�X�����E=1OZ��䡄G9��2��0�(�ꔫ��,i>(�go���"OB(���Ɂ<��z��,I�y����#Yؔ�soˬV��DX�*.��6]Ry����)x¤��$Ȍ�6/��Ɠ�Q`7��hĜ�����
�"�ju��tR��&�L�	��5��1��{c Ь
��h���<]O`��I�X\�����|���tfP�2^�����F�p"��Űww���3O8d�Æ�-iȨS�u�zXд�x�Ԩ9��� )�r֨
�E�Y�'3'd�P����Y2��/=��]�ȓ"i�h�d�	$���q6(�>S��!b2�s@��x��Zf����`�'��MT&1�)D����E˚0O��*��$D&&v]J7@�*L��G�J�M�RL
���&q	�ؑ�A��<�2�
M񾸲FB�e� y���BS8���j�Yj���	��G�*�"կ8��a$F�Y9�FV�T���N�]�0�3��}��DQ(A����'+<�۲k��U�XŃ'	�N��Q��3��k�Z�9��(jD�M B䉂n���Csȍ�3�q2�S�J T��hO=2��[� �$I@���yJ<YW��8 ����00r�H� *Ma؟V� Q�=�r�H�wL��&Η>0A�)�葢.?�� 7G��o�n�3C�\2�<�w��y�$�y�٤!�\�m_�'�:ݹ'�R�Dx�mRҮ�[����L�@Y�6�gx�p��,mvn$�O� �8b%ǌ�Hla�Ǩ�'�l!W�O~Hb0˛�E%�@��Gi��fG���!�$�(X.pM���	� ����u"O�YB�H$jjp	��Ժ+A@��2̙%L�d��!�� ~@���$ը)��/��&����ʌ+oP�� ǩO�H��S
#�O~�	��P]�R�o��j�t�-J�x)
uX5�Z�0����jޮ0���0<O&��CG�!��T�E���#*~m���I�6y����,��� �$�hV�QB��N�_�]×n6E�Dr�h�c�m2	�'5*���� J_>C�W8^�i:�'�&���R34(`]�#Ŝ�e9<����H\<c?�zE%
 ��8���#���G-D����=�	B7P�(J�0��K�L��a"v�%��J�.���
!�J<A�`�v�<i҇��9d;�8I$��i��,
ԣ�v�b��[�`�H5e�;T͖ ���_�/��-Е��RX��C��ܸ'�νB��u}���*z6�s��U�2$�t�a�P6��O>�z/�!y�ā*���h?V ���*W�詨ш�]������
'��CSJ�Z��vo%�m)@�i�l@.m&����	`�\A�f�����#G��Q&N'k"T�)��@�l'q��0h�B�	A����ϟX�X�f��s&�0�egh�#���t�ʍ1�,��x�P4��W�'5bYz�m� �b��WMq��靵vm0'���գC�*!|@��0i~b+c�9�O��P6�<��F/1�����P�(��	{E�P�xi����L�
�R�=��&D�zH�-�V�9��RqJY�m��y���ɛB�8�؇�߫��5�O��*�\�!� nֱ��cڏ_�*����I�-�6�4�YF�'�1Xˈ�aq��p#D�lc��O����Ě#Nt+S(�&e�8�%��p�O0�S�"ېR��L��K��V�q�'�T�w�L�����(��G�4°�E�s"T�jH�}�v$0DH"��'��'C�i��}F���mߕ|[1����Q�wJ��n��:7�4PS���lY��k�D\(Z�Θ�3#����b?\O̕(��ݝ^PrVO͘FۘĚ��'&6����0��=�E���db@m�!q>��V圮&���A�a4D��S��E9#������U�=��"0�g\ B�*!�H����GR�<#�P�1��8-����KTB�p�N� X�B�$7��|�ȓa��c! ��*}
L��.
/L�6��ȓ]��,����6�TE�w�[/u+�ɄȓP���c�fߵ23�Ƞk�*3��̄�C�݊SN��d���ۜ-�>��ȓ2:-:�ER�;g Y2%�#)h䴄�U�ܩ#G͚3E�  dрB7 ���[/$����O����J��x��?�� �C�\4Ix�	a�:����ȓ1Sҁ��L�7��|Ab��x@�\�ȓ9��Q�Ƃ? |6���J<y��p���%��<ѻ0+��j�>��fبW/��\*�L�V��DS�ɇȓ`�� rb�jp���処I�Z���&%���T�d����H%LU�A�ȓ&����F]#k��T����-��ȓd�H!e ��r&@虂�ԍf�ph�����j0枠S+Y�ĉ�B�5�ȓu�x�t��
�@e��e�2�v��ȓf/�icpg� c�l�ː��j]fa�����E�ʹ�~�K&£uq�5��|oN�T�X�2��ࣂ��pGȓ~Hb͑U C0"C���W�B�K�A�ȓC���$Ύ������G�P̄�ڊE�t`�g�$s�c�7s�`ņȓi:�+1l�<�l}�#��	oP}�ȓm���eߝ7�8h�7H������ȓz*h|�Bfm��]���w(I�ȓ)obl��%֢$�"DH��a���ȓ@�č;d턗O_�ݓf�	%B�p��N���T+I���6&]&����'�h���I�+��l	�J�p��ub�'�Ġp�S).۶<�S�I?i�&�*�'���a�	�R�����̗=�M���� ��X�8z^8��d]��h�T"O��Q�@�7E<I��$��w!�"Onx�Q�ޅWs64�$I��'p�qc'"O�%"$�<B��=*u�1AZ��c�"OF�CW�D���)GBC�M�� "O �JQ6U9
�p��#v��"O�0��ǂ�o����t�Ȝp�V"O��Z��^'���7�G>�D��"O�AxƤ�u5�4�A��Z���2"O浂�hV
1�Α���%(d,�"O����"�*��[FF���xe�4"OL�
T(S�V�ic�GZt �Z�"O}���`�|y��@�+cl~ �v"Oְ���*z6���G/��B��f"O�l3�K����g��!�Dћ@"OX-⑁N�:�+EkI>}���S"O��!*+�t�*aE�)���"OHP8��۶W���g#ɥ�hЀ�"Ob�т��?/���:�Ǩ��A�"O"-i3���E���@��ʜ$����"O8� 2Ջ"��(���"ȐT �"O�8(�,G!q\�4� %úFZ�h8�"O��H��ң��i��'?{(�CS"O}X���R��q�#DRzu"O�����>qL�����)9v���"O���Fɼr��]��c�8la�E�"O����C�P��1�sa�0��"O�ܠ���\� �;«K@���9%"O�"�f�2_!b�(�`��L�"OJ(�Ū_)1ehh�͕�ޅ+�"O�y{2䀾��]��
+o���"O����ɖ����̕��"X��"O6���`���YQE#;%`�s"Ot %�^	$��YRE�,:b"O��)UD1�kG�j���"Oj�a7�L�W��p����.��y"ON���NM��=
5C�f��xC"OLY	��Eh���2FDL5t�2l�F"OX- G�B����LB�"�܈Zt"O���s$�N`ZH��ּe��=��"O^�W�P�5XD��M��e��u�"O��h��ùm���l
G�ԕ! "O��Q���*$���4L�(V���"O9�*
�>�"��ۣ �"�b�"OLHP&�Q�-~��Q�KN�V���"O�FK'/L� 0T
T�^>�]�';��Cl�k2j�";��U�	�'Rȡ���9P�E�SI��e&��	�'.-[��L�b��4+Ģ^^E̱j	�'jd��޼2u,p9c�S�Oo�xx	�' f�h��*u���˲jP����'�U��)�&-/pH򂔦Q���`�'���:�*ك08��s1��A�vD��'mPyJ����E^��Q�IFh(�X�'"��f�3{���2K3Iw���
�'x�၁CP0K�F�(5�e�
�'"��r#��"My�|�V�� {��٫�'�H��W�Z+8'�峥Țzư"�'z*��Qc�1���һbd��"D�$StǄ�i��P�2a���T�a� D�(�^�
� a`R�F�-"6��� D� ��bǲ���ô��Sd�-z�?D� r�	#xt9���¢r����Q#;D�P�U�#`͈U\?R�X���<D�� `��7�UK�!3w���`����B"O*Tg6N���d�&Bf�6D��&����|@tE�3�Bq+�7D���t	��\P�'�)��yC�5D����i��!v��C�N ��f�1D�0 ��(s�|�X�*L�U��X��=D� )E�_,6L!���1%���n;D�P�a�,q��mq���>b=�1:��<D�ؙ��4|��Zfς�)Α�d�!D�Pc6���O
)����(�� D��K��Dl|�j鍡*V����,D�x������@C
D$̨��6D�܀�($HB�|!0���x'�A� !D��p�*N"vEt����%��A[��8D�����,�%�1ͬu�&�!�C&g���bִkζ] 4*ûC�!�$�� Ğ=PM9��!PW#ÓP�!�I�4nȹ�c�ۍA��(c�#��!��i�DX���f���!ղue!��7F����Zz�lQ�II�Tp!���~�v`��`7B5#��S!�DG�$�0S�N<9
�����	 {�!�^�r�ҩ��N���1rƛ��!�$�S�*���ܵf�:�y �U�!���y�,a&P~В'�O��!�$�
_���$��x13�[�s�!��-"g��q�ŎPjf8��HOX!��B��r$����%�F��r�!�dA�f�ܽ�����`l��!�$�JK���"NE�\��\p�g�N!�D+E��%9�#��2��JtgY�4!�$��EM����R�wPM���	!�d�	����e�>X��\y���8~�!�18����qh�`x��(-^)<�!�$�'��!PwnI�R�Z��$�Q.d�!��"f��X�g�f|�x����&!�_�i|�� ��dV޴���P�!�d	�y�T��dR'y�F �F�	�!�I$���`�$=`Z���+�*�!��&=N�K�%�1l��@K�#a!�d_;[6��{�&�J#*	�lǋVb!�D�.^�T�0��L�y"PS��T!��[�
m�U	��C��HS�J:!���	���фIٝ3��MP�ޔ+!�Ā�;*ͱWmA�w�H�P��>\!� Z�Dq�3eQ�ϔȚs��e\!�$��-���'ه�h@S�/݈v�!�DB�h� Tؓ��.��`�.�2a�!�$ΆPꤘ�@�Ȏ\�.��" �)<�!���H�f��?����� �J�!���<���ƙ J�t��!�
P�!򤋿y�Z|��D�euT�)Ʈ�1
�!�ѭHR*)��V����nʔp�!��<<�FT9���<5�y�w�,<D!�$ܧ<��b������	�f,!�d��]�� ��0n9�mZ�G]�!�$��T�Y
Q 9���Ð�V	V�!�d�b����Ҍ�g�� J<P�!�$5�0LF+y����,��?�!�$tP�2d��tٚUhx�!�d��$}ܘ16�X�FQ�7�S/j�C�I/G�$�e�^Z���"5��
��C�I�fJ���[�t0���6��C�I�?��yG�;]
�W��x#@C�)� >�٣nͻ[�0Q���_'A���"O���*B6�-����weA��"O��y�J��4U^������p<�� 1"O`A��]+!Ϻ�I7��<�Q�"O2����9Z=$��A�g��� "O�b0�4Vyf��B�0l��a"O�@Ғ���Ud�,��L��PQd"O���p�P�E��h�DJ�>ud�m
�"OLQ���Ӯ@�r�
��W�h�"O8�Ƀ	g.��j6�B�B�`R�"Oh��퍓e��8c�KQ���3"O$�ӠGɢG��"n���J$��"O�	y��ڮ���@AB}eNܰ�"Or�8 ף<�`;Q��"=^� "OJPt�p����Jz 4�@"O�����/0O��r��Q�N����"O0$��d+�4,J2�L�v'~<2�"O����0B�l�Ǯ,�\ ��"O��;�FŬ�0�!�S9Oި�"Ov4*5.������Q�g�4��"O��G"Λuq��CWɓ'~��!��"ONe㡪�;#tբ`"�V��[�"O(��,�Rx�a�¢?M�0!ل"O�����"P�F0��kH�2���0�"O�u�o��"�ri��1U�%J�"Ox���K���.[u� �y�d@�A"Oj�-@5r�>�"��*v�R	�"O���(�:*��Z�*��l��Aa�"O�eҁ�H2,"Ш�4Aޙ���;D�`C"�3#�&H���E�RYY0�7D�TǣP!e�X�����a#�+'D���p�V�4���$� v04X�8D�ܙUEE�Z#+̈B\�)(��>o�!�S:t-�9Z��8"Sj[� -�!򤅙:R��4��8���.�C�!����e�Ǣ���X9ǕF]!�dr�.����͈]�"�iu�%D�!�d�%�8� ��Ur"�ʱe�
C�!��֐�R)J�i�:)��Z�!Y�!�^���PP4��#�q	�'d0����,l��x�&*'�A�'R-�6KFx���%��E����'��\p'�]�a��a;o�5?BA�'��0�Ǉ�G�����a�!.�H���'�|�	W̓,'�VX�O��Tp�'���1�/�(i( �C#�] �'�4Xqe�R�B�~��3�l��'Gb��
 (@��� U�,(�2`�
�' $�� �F(��Q��²*����	�'2�1�'��7B�������R�p
�'ξ�ic��J~�dq4�ϑ����	�'���P`���qk��#�	*�4u��'��+c$X);��h�-ӏ�8�!�'w8�J!�K�fњ�ȗᕽN8	�	�'3��� 8>{ʉ1�Ǐ8�b��	�'6|8G�KwP�ɜ' ��Y��'lx3f�H @p��W���8+	�'7J��C�׿ �2d���_8Dd�)��'(�ػ� M�89
��A"��C��@��'5v5�r�
is�<���%>@\���'�\(��)S�+��X� 4Q����'^V�����G$@|9�Kڹ!D�T�'�
x��؂)Ԩ4� $+���'8�\�d��2CF��\�a������� \��f�B��8����΂�Q�"O^�X�H�!;\��@ӊ=֘A�A"O�xp�E\#6����&��7�>D�DxF��;q�x3ag�-
��9�t(3D�h�2K��V~Y�U�؀�޷�$1D�`@��$N���;�M;����,D�`
�@�.x�c�Fɉ�@���o*D�HP�!�s*F�z�n��dvXq���<D�\#Ў[�.3$��2I�b�.-;D��!KE�X��d�]y�#�"D�SEM��
t������Y�ѡf�"D�d���O>MBFy����.'���%k>D�<mޣS;�����
|7�t�S�Re�<y+��4$�e�FB���dh;�M3D�$�.�:vn���Ñ �*�`�.D�t�k/.|<)�V���a,�§� D�@A��:�^��l˟NH����"D�Ġc�~b��x
�N߶-�b�?D�H�́�Q ���@�� ����:D�SRM��Nn�U*�m��<�52B';D�xh�I��eZh�5��+j��@�D4D�L�$�5� bDR�^dy��)D�4)�ᓦ��"�"ԒMyN�b8D�@���xC�tq��U�Km���,D�@g�����uÒ�r?�˲�*D��@!g@2Y����ïD*u��$���&D��t
ػP��%B�	3��P!ԧ>D���G��Sp�d8���%Fiلa=D����*P�87�a���#G�H�ˣA.D�8�׆�>��� R!�,'v�A�*D�\8��=�8���tRV0�Ɗ(D�X�VdT=fԚu�a a� ,��($D��b4�Ȃ
�F�3�ݒE��顫%D�D�VA�Pzޕ(@N5J5�!�ah5D�<�W�M"c4���G�;M�^�I��,D���%Q�4����b��:>��ٷ�&D��!�j�piܼ����(W�(!@G1D�,蔠	�)��!ɇ�C-6hI���5D��ae�V�6 b����Nшw(4D�p9V._<EX�A����$b4���`2D�l�U`�`徭����V|��E*D��g��%�Dq[�g��S��XCф>D��'��H�8��^1�x�Vk:D�h#�M
>�r�!���$Xx}��;D���-��j-<�z�_ q��`A��*D����g�]8ͳ�j�(F�*�1�B&D�P�J�M��xs-��!��"%D������.�V�X0o�<8&���+$D����O&k'�=�B(�Z x�D	$D�h�/�F�����
qP�i:gi'D��ʿ,��*rgS.6�\S�%D�tS���=Ϝ���B��PY�/%D�� ��=8�^a�U�� ]��f�#D�,J���m:|�RdJ��N!J(r��%D��9`�C���HE3�b !D�4��kCԑj��#11X�aF5�I#j�HSj�=Pc�`kBN� aw �!�B����2\$�\Фf��
�R�j�I��%�M>Y�JYi>QH�'J
]�L�l��?�&-*��QE��<?�$)"��1���S�ݠt4|�V��?n��LPB��l���L9�ZQ%�"|z@�K�NZ�(6��
�������<�%ϲ`�h���KJ��qP�c�O���h�ŤP�VUB�O׽A�����4Lإ��'�v���'���(F�(��|B�I+�����w��I{�G��t������X(am��p�}���:9V�����}z�[`	�4�6��sE� }.�L�	?��9I#Oc>	��M�s���A-)3&(Vg���JX;qk�8К"C����'9"~z�g�? YEKѢ�B��M�b��	I���X��(O�O��)�ǀ׷t5��!w5&��O<aF�#�S�'6��A�%̈́3p�<U1Pd= �jt�''��Gy��� M��[�k�O=r��$��ԛ��7��<�}篑�j������BZp���KĎ��|����џ@	�J�?D�j�·J<���ħ<X�31( �u'&a��ʕ��v�p��� �DR:�^M��N�O=Z�ې��?^��\#�锂.zZ\�qoJJ�k?�IA	�':D�����5YU����mי �豆ȓ"H.,����K3J\-aB�d���2=���Ώ!�Dd�!
�jp=�ȓ̎)r-��=��Cb���[V����oq0-rViL��DN� J��B�	��T����f�t
s��@��"?Ɉ����p��p�%H�EQ���4F�X!�J��`�X��ͭy<�$p��%�!�ǥO�`(�Q+�-A�h֊��$N!�ď$m̩3��è?����X�KC!�$	��H��fE0E�)�a�C>C!�$I�hD�
�o�$I�a��ްq)!���m�mcE$M�j �Ig^@!򄓵R�|�B7AٷJ�$tzD��?u�!�%A?LKr�� :H�<¦�."�!�D��0�2t(�Q�^B����Y�G�!�d1M M�u��m�J��%�,�!�E�%w:�[�[
뒤�W�T�e�!�Ď�n�lQ�'ID6T�,�!�Ȋs�!�$�
�\��ܩA����Y�!�$H�b{j�*E+�&!�A`ڪ�!��� ]���I!� X�!�߃U�!�8�]Ӗ@�&v�( ���ԗG�!�$�,iE�Dpf@ݘyb���
�!�$[�? I�PfÎ�~)��B�-�!��/!�Q��Fؐ��C��Ts!��^��v���D�K!`��$\Z!�1����V��#4	�=���)2�!��ާ��S4�Oe^5b�ډ
�!��P,v����H"7��q1Ѐ�L�!�dK0�QV��5�jɷa�Gs!�i�VA��mU'z� ���!^�2i!�dS�(	�-�C �cŞE9���f!򤛷�f��%+��i0�ƁY=!�ř9T`��Ğ�G�聛d`-</!��K vE6I��&T�QӪ�!�سPˡ�䂢��12��k&��C��y���=I�"�k��R��NX�&lф�yR�  
H�9V�C��>��� ���y��������<�n�� ���y�N�Q/��y��8N���TNG"�y�\�Va�$��&��)�HJ��yB-�v��H ��ϘpN��'L4�y҉�� ���A�y�jU��dД�yh�&s�������8C�mc�`�;�y��=�l�����m�(���K�y_(W�z����-j^p���I��y%ż8�����gU%g�l ����yB�˝`��[em�vWȵDGK�y�#H����ě�|�4�brL�%�y2�R�?�����mƉ��`M�y�\->���JaPr���Gթ�y�oR�$�XwG�m)Z�	F��yֱ҆H�6�+�Iە16	r���y��U�_7T�`e�� ����"�-�yr"��%�hB0��.n���t,-�yr!E�rS�T)�oɅa`z�� X��y
� ��Ju ճi>|�%K�9!F\17"O򽘕	Li�iH�gň,bR�"O�����=HH9�&��D�p���"O�0"� �)أ��F�!"Ob��2�\[�\���_N|̠�"O��q �rn s��Z+NVQ��"Of�sb�P|��:�⃾k��
�"O^hHa�W67�P��W�[�fS&Q"O� 2�c�!<%���û?�<�U"O�d��mD� )��P��G*�"O6թq��;��`S���)}"�)r"OI�TL�lL( ��J&W��S#"O
��ƤUnP`�����\��8"�"Oj�Kf��l�R���ύG�r���*O��0q" ;j�"�b`˜TŢ���'���R���
4˴�p���^ۦ�9�'�^U����)�؈z�l�U P��
�'6��ϟ8=�	Z�e�|�t��
�'����$)�2�z�����,� e�	�'����P���|u�(di�	�'����jZ�g�8�S�̿��y�'�@p��r�v`h��X�Mv��'R�� _7�|=S�ϟ��F��'x��5'2g��J�BT�)��Z�'`��ǌ�X9xA�L��n�r��	�'�)��e��<憐�7(O3��ܢ	�'���UmST�!�"U�2�d̚	�'�>�f���e�h��v�6�		�'���1�S
y���Ï^�s��k�'S���CMͯH}���HA1dv~��'�d�@�l��WK"ɹ��O�`vb�'z ���74r�"�o^6�s�'a�����Mi:����լ`î���'g�Ճ��>#�j0F�B��I2�'��}�:��L"J��Z&�܃WW!��X�ȝ+���w* ���ޛF�!򄀧l�~��߀@�y80��/G�!�"e3B�З.�?RM>ٺwa�4P^!�T�)��8�`�-I4|(d�ͷ�!�D�7J������J=.-�ABH&�!��l`*lp'��(G�������P�!�$A�\���:KY97@��Q���!�D�"M(�@��胎-���/\��!�΂P�@����#��ӭ
�!��;�����X��:��0� �}�!�݁�Jh��#	��x���~�!���yF��@5��<��ۧC@�[\!�$a�`���D)  �9	7@ʛq!��F��z�F�x�뢎�%V!�DE�%�X��s!����j�*t��"O����'�s4pA�B`��M�Q�v"ODxz�.BK�N4�Vn9)�"�C�"ONܙ
M�[~��؂�� +6���"O�8ۅ4B���K�#艊�"O���3fY'P��,��X�4 �P�"O䘢 o m����g� �i"OMٖ(�wt~�s��LM�$ہ"O�UXB�)� XKW�4Q�P1j�"O�a��"��z&|A���ʻG���"O�Z�&��U�ĵ��G�<� ]� "O�	o	3L���ƶ���AG"O(�Y�E�\O]��f^�]���"O>�`$MN�g'�H�!%f[��]�"O�Yʑ�β�$8zw
y�N��"O� ��R��8(�0ɦ���JwЩ��"O`�y��H�9�z��oP�G�n�
!"O4�!勆�*밑��N��{�Z��"O��;u���$)@e���}H"Oƍ2��N:>���#c�����pt"O9��$]-�\���4o "O�[�)��z#L4�䀀�Qh�!�"O�[�Q�s�1`��!��%�"O�=�r/�$,�n��훃z�ؼ��"O�0�+K!0��|	%�)(��!p"O�="t�J��}�1���&OtH��"Oh��c�#S�
���c֟o6�5�"O�����p3��	���yNՉ�"O��T�)c�1a#�Lܑ"O���I�Z��m�&E�o��]�'"O�hf/�=TأBIM�O�$�""O�\��⓴#�����'�)"�"O�A��
�X�vǜ��\�6"O h�� ��H�aWH^���y!"Ol�˔�H�3�t"6A$plbu��"O��R�9JP�	db��yU"O��">*r���%ƌ&Hj�b"O.q�sF�KD4�вD�n0�h��"O�x�!ë@}��e��\��q��"O���Sa�3wdm�F��1��6"O���A~�Jr$�ף/�J���"O�A�ɐ�"Ȏ	� G��y���"O�קۍg��E2���#|�H�"OZ�kS)���R���aBƨ�%"O�Q�W�À�:$NF.;��!�"O��B�F&} �JV�ض[:v�r�"Od�J�C�D� �ڥ��8�(��"O���2<�|����M%����"OR�C����A�%�TW��q"OESDK֟_�4����VJ��(��"O.�3�Ԕ^���Ru��)d.
!�"O �Cը�`Z��C��V&�)�`"Op@Q3A@�v�5�]�Bk�:�'l��D�O4F݃ f�,�h���'{T����� ��,�B#�)@���'���� ���VCJ-)�����'5��{�#�)c�#�,��1�h�:�'%@����_�9�x
[%-`Q��'-*�4n� �.�3��M3��MQ�')� #夗�i�d���L�|^�j�'&���-ƇA�(��ŏy�PX�'B�|�� dMp�����wb0%"
�'�ȁr���w&����,2<q��H�'���WݮI�p]�P�]�94	@�'?�l��mJ����``G�8W\�'/����(C!�4�8���t��',���D �C"6AzĲ
��%��'���0�l%C���q���I�',`-x3G�4$����Q@5h����'qĠ�TL�	r�TjRG،]����	�'~�2�`$��H"�_�ִ0	�'���z�Ǭoe��;���1�+�G�<��<���C�6��#�@]�<Q�&S4<�@Wl���0��\�<y'O9��K��>8��T�QoDW�<	��4~�|�1����]$(h:pg\�<�"`�-<Tu2�ؔ&�fJ��T�<�� ��f���#�G��r���J�<��*	�?�y��P�k�pe�JV|�<� 25��h0k��#���70ƺ��q"Ob�Ɩ��՘���i�T8��"O*|��h�8���Z(.j)�!"OJ����]=W��� <i.�j�"OT�1"�HPp�1��J p� �e"Op|ɐ�I_J���Ӎ>,��ڀ"O��1��<&�@iR�B���!���`>.}[@�7X��K4!�%J�!�W:�D16�V�rH�c�N$T]!��D8���(w�3S�()�.;{!�$Yv۸�S��O"��S�lE�JY!�d7;Ú`���'v���q�M�.�!��]��Rƽ�����.Y, !"OީjaǤt*x��/I�Z���"O��뒤 �}c|��b���+ۖ8�"O�Ԋw�\qKp�qlFe�~)rW"O0e��ˋ1E���������"Ox����{��H3uKW�QwX]"O�ܑ��φZ��]j0+�!*b�t�p"O4�d;�
e�"햼IL�+�"O�T�CϏv 0jVL��X�$�1�	ş���E��F�i z[�M�c�/����6�T��qOl��u�� �CK(���)@Z-q�p1i��N'ת���L�
?.aCj޿nࠌi��I1��m3���3Y��ЌS�n�D@�-T�`�����$a��x%ASe|(A0�剄Sx*�$��MI�4�?ᬟ������=_�:�*�O�!V -��ƚǟ �?�O��Oƴ	q��!�"�c�
g� ���'�Z6�զ�mڳ%��X�DkFP�AGIe	����k�dS��Οh���`m�pO��#��Ѫ0�x6�W�z����X;T��1��]�e��Q�jPfZ��7������_�!�F� �v=���iJ6-I�ĞA�u�7p" !���Ĕ{`	�T���"�
l �@V.`=�\{ҥ���Ca�Oz�m��M��䈟���џ���E�� )Ν	O�~2�'U��Z���ɗ~��Q����s:����*FhQ�\��4f�6�|b��"\wlĨǋiR`A��Ur�4�0!�<!P��Xe�&�'BT�pgU�B����1�@-S���A�ɑ��B�m�:`�pSV��&BV�I�2s�N,���|��v"ą*"��3�,{��+$<$"�&�`a��(eX-[��ؑ�&B̓+�6%�� ��d�ө �U
���'�8x��0�&�:��O��ķ>�%匱�hmc C���y�f�
E���3'�?�$�t���{���+ �^�h1��
C�"�g�d�mh�	�?���{y��Pj6�}�"�J@zR�IևK�(�h�S/��y��')���_��bT)�I=E�Y!Ӭع,g^x���BZL ⇇��T%�2�H��(Ox�B���{5���HΓJ٠�`��@3Lx@��D<
����*i����4�HOH�AC�')� ��I�BГ��ܘ2j@�i�H�8RQ�6��O�ʓ�?+O�b?�j�l[4|I���ՠ兏Bs�B��?	����i+Z��h��IРD���I	�MD�i�剞d�40۴�?�I|"���6x���Μ��ա��R��?���ML>��P��+w�aG�([�L�Yt�.Ba�Sj
%�v��@B&Rp5Ey2B�.��0l8$�6T�bL&Bڡx!�\��!\�B��C"J*j�����鉽.]�����xK|��4c�(z��	R�H\pE���Z�2��'�O?��KwR �#�l�1q�p��`���E��|��f�T$n��A3�lҐ.h�����66L�h�δ��+�ٞ�M���4����-�dN�@� ��R�я`�)(׮�<�� ���&6�uoa���@ܥ�@`�6�����	O�"�˓�5 D���@���M�3o\�J�]��m��l)1AS�+���]G��+�*X��SV���`�A�ܦ�b��O*�nZ������?7��'8�&���XS�Z+�g�6n�~r��`I0랸!ob�����>61�(S7.(ʓ
��ևrӐ�?!��u�pDA�(�	�0���Xg�|��'KTP�� ���   �  �    �  �*  �2  |=  �C  J  �P  �V  ]  Lc  �i  �o  v  V|  ��  ݈   �  b�  ��  �  '�  ��  �  G�  Z�  *�  l�  ��  ��  ��  ��  ��  �  �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d�O�=�:j_�[����q��Z�|Ӂ��H�<� ���.�:�$Β,�^���\D�<�$��
c�
�sa
��A
#nC����<)��7Q�D�u$8]h�����P}�<���� U��\+ OT�%2��ŋu�<���^ʤ��H�K��U��ASr�<�7.D�(�3��5o��Ձs�I�'�ax��ӊU�$c�H��xF���"��y�Ì�I�4 #1m%��u�������0>i�/.f��4�s��4D��`	�x���'��p;E,PS�U�B��D��<�'��8�I�)NX��a��u��y�`
�&F���4'�ZpbeaX,�y� ��"�f���S�iJ����y����h`h�v�L����D1�B�ȓt�V}*vL�TD@i̯t$h�q��~�	�:zxnt125��1�y� Y`)�щ�nl�5��ޗ�O���4H�Z�F��O$B�jv^��!�d�O2�HWJ�*9]x�ꁷ����@��y/�'(c�,����:�.��r-��yr�ǲl����"6$<z@�%�y"H�I�����V�����?���hOq�XX��g
-Ph@�ݱX&"\#W"OLl;�`B�dxh�o�1^#���i�����H�S�A�4�ę�#� �aL��I���� ���2���,�tlV��s1"O^�`�퐰l��H(2"�|S�"q�'�H#=E��-�>G] }ض�^"DZ0XR���!�$	 k���4��~]&u���y�e���Z�F�:&Q�sȓ���`�(.D�h���G2� %k0iΈX���6�7�Y�ayb�QI(���*پ#�\p������hOq��l���H2����,NRZ,(d"Or�i�P��r�ʣk��
S�D�Ӧ��D-�bO�J����S#��P���D/1XZTi�x��M�rX�'Ka|�m�(f�m�H�?�P���E�y"
BQ����-�gj5��(���0>!��9E���)]�M�ҙ���t�<Ic���X(LȆ�J���v��n�<�-E
Cl �X ,��%k�uې�q�'2����O�R�1w�>'�~A+��U�ghz��1%2D�,��%�.E���*�=t��!˴���'�F=O~��h�'D(�@��nY�	�eB�.�BB剕m��H�a	Nac(-�2f�1Z�,ʓIe���ͮ}�D@8�,�#M�j�!PiGb�����j�'v������Ï�9��`��`O"R�
˓�0?gH��NPr`Ƒ��0"V��\}B�'ӛ�W��E{�'k�m(����`�(TnX�>le��I�<�emaӼ\�'J)q�>��qbR�>+�Q"O��3FA=��)�s�	%6��x��I?�XD�ԩ2S������
[���v)����0>��1V��U�z�u�v2��O�7M<�&
�&X��$/6� ��w���e��� wȞ5��x"F-}����h�1�S�̐��ē�~�b�r~2�=��'�Iٓ%^N*V!�NC�%	�|��'�<I!��Q���%���ی{B�)�I���mIb�~fp��B��i�!��C�2���b7�̦T
\T�qL]K��<�c_i�"����q�s^�$���ȓ��́F��v	hiڱ����n�s(<)�@�1P߬9�5�ыe{ح�ʗc̓�ў����c�a��L��`A"h9�"O؁�7�\��i�b-���"O��@�ܿ_LhK�!��f+@�Y�"O|�K�r.PlΛY�0�s��'�y�C�Sn����� 	���CW	�y"���,�<��4p~���Nм�y"g(g��|2�AObA�AC5^-�yBb�"��L��ȂP������
��yrNٕ h@d����*N1R<b# T��y�ߧW�b���G^�HI�)$$�y�X�A���р�8E�-��L�y�bL�GG��H���B�d<�q����y��T+@����b�Q�(���y�ḽ3�|��t�ĚL#�(E�P��yB�R���C�́)/t��dM>�y"��,���`�����=����y�({Ɇq`�g�'����K��yGֲ4��=�EB��%|�U�q�P3�y��U�yW&�3�Y����O��y" m��eh���~���LY��yr��yf��:c���4����'�y�[�+T�8��K9�*U ��_��yB�V2�8|�҃�Ho@���jJ2�yN�h^��z�o�=�:	X�˅8�y���4KǮa!�돾-މ;��W5�y�� 0��2��Z�)�&tR�]<�y��
�e�������(4������	�y
� �4+�
��T�p�b �X�?3���"O��!ҥ;MN<\`�Œ�zJ��h�"O�5㱫�|l��!��)M��R�"O�i���7���TC	.�hl��"Ot���۶4<C��(�m�*O2�1d�F\X9�Ǥ�po~lK�'�^�#U�B�R)����t6���'� �I�kJ	Nr�a�M�]���[�'�R�VL�'ᐡZ��Ԑ]����	�'#���h=�m 6�5P��'y~�rPـ�BX���y�����'�|!�ȑ�Y���νb�X���'��I�%�^-:%��H1P���j�'xՁ�`���Z���O�C)�'�&3!�G ���YQE	P�(�2�'�*칣�b�4y(���V��Ś�'B��c� 9�h�#�N/Pu���'���p��4M�ZLi��U1L/��z	�'�e�s�� cap�R`BL�)�'�\0`��(mB�Y���F6�X�'8�(����;�\I���>,���k�'Jb4����r2FX�*�e��'`�0P#�L
t_⌰��,%+����'D����V�&��4$��&P�l�'�N18��A���A�B=���	�'پ���퐴C4�!�cgK�4���'�8l Å� �l����^E��'��0�.^7?_��k��֟{ᾡ��'�V��tD�_^&]Kq�K�l�����'�$|�&c�������ת]h20��'��)qiBQ���k��R�X�DXS�'��aA�Pq���S�yZ�'���I�].t)��p�N#�^���'8���Mˇ}�l=B ��&�xx�'���F�N�\�5��������
�'����Vi JJ��BF(\����'ݪED�rɖZ��I:|A���'=��i�ƕW70���#w�"���'H�Z�@�m-@y�Z�%�J<k
�' ��� /zZqp�+]�q5��j�'�X�re��c:	�r��q�� ��':�ЇeԊe�x�b�S��c�''�ᠤ�ǣ�vX2ѯ?Wv�[�'ڹ!tO�+��!;c"�0U�j���'��̊�oα\�؁�"��Jk(��'���� �YKt����G����'�6���Ş?�h�8a�[�3�\P	
�'�Π���S���b0��!{8��	�'���,=b���)\�נ�	�'^���G�I�/�:��g��H}�l��'� [d�R
9i�����܍T@<( 
�'�a!�ە3q�0(pLz �J	�'8�H��E�v-±�nY�H�<��'�`|)�	�D�N8�ש��A�����'`���uPx��ȒP�B�+�'�nH���q$|�c��7(��'�2�K0
���*����w��d �'1��ҕCK�Nor�C� ��Y�Q��'�F}z�>��y���*S1�#�'E�Yi�8>p �R Q5~\�Ԓ�'N-�r�U�7g�`��]�I�~��'�����b�~���A
@���h�'Vy"O&�hQ�ᆗ%*Uf�k�'<�|&.��h��h�p���.�|T���� .�U(
�7�l�+�K8Gj-� "O2L�Wt`��l��6���"OL�"䇸#�b�Z�+ƕR�L(��"OH�d�O�"!	�
��|i�I�"O�<H�IAc��i�C(Z�^Y���a�'���'���'V�'�2�'c�'���c#mʊ ���h��!MlE:��'���'�2�'���'���'T��'�H	B-Ȅ��KZ�B/�����'���'��'�"�'���'��'����+/!$�٘4�	�� �'�"�'���'���'*B�'��'�<8$U��q����+T�ܥc2�'#��'x��'���'���'���'!Ti�`�;YjDi�'S�	�0�'O��'gr�'���'$��'���'A��Z�RSV-�̓d�Vш��'0��'`r�'�R�''��'�b�'>��S�;H�j�( J�"4�'
��'��'���'��'��'*w�-N��Ã��
u/N��P�'�2�'���'���'���'%��'�:��	r'�y��[9."d��'���'���'�b�'1r�'$�'�L1�P�Q�n��dX��VI�t5c�'2�'$r�'���'���'���'��2o�>��K��� �0,{��'�R�'%��'���'��'�r�'��������OW���l\��줡�'��'��'�"�'��G|�j��O��bB��E�ĸ!5.J��H�3�&�oy��'��)�3?ag�i����e�s��"hE��9�*�����ͦ��?�g?��4pC���6R_P0�� ݼ��'�i�"�ݛ���h����-.2�y��~��aB�*�[���&	8�I�r��?	+Oh�}��	�j��}�e �4�&UawC�S��F�����'�񟠭lzޥʡ&@8Cؒ�R��
+S�� @*�?9ܴ�yBZ���jM�B�vӸ�	�$Z��IdHv�Kw�&Y��I�DT���M�v�`hF{�O�B�\
B�F� �&	�3޼5y�I���yr\�|'�TJ�4,Ih��<)Į�)����!E#��cb�&��'Htʓ�?�ش�y�S��4O�2Z���m�{1nm��-;?I� v�^�r5�]a̧\�R�S]w�@��	;�>��fR�yOv!�PO�.0w����d�O?�		D���T8F�1��Jܽ=��I�M��hu~��r�(��ӵxoН���[�\`r�m�h����П�nZ��"�G٦��'��9`Q�ڱ��qA��#�bx�ℝ�	;ʄ9,��9�p�C�o�+!�e��F]Z��L>��F�z�|��L>j�Z�Z6.�W�<�VjU�{P�����
L�w�ͨo�@����R�\���!£u���Z��V"krX1��L�� Z����Ȧs�0uJR
!z�X��O l�Sgɸ)X������X�P� A�65i���7)"D8*tJ*,<���e̶( C�TaȂ	� �B�I�T Z4�Y�N����%K��0,�	&j��U������	�?m �O6�F�a��p4*A�KW.4� �i���'NAXf�'ɧ�OwTPb����b�` ;T��
$0�(�۴F��`�i���'L�O�O���@�̴�~�\=y�)Ӑwв`m�9%��X�Ik�)§�?�Ң�:nJ�٤�O�N���yeI PM�V�'���'K�yp��)��OT���x��꘍��q�u�����W6{3���|�j�I�f�f���O���ձ;��A1S��4�
�.�f���l��0��E����D�O����O�Ok�
h�r|!3��7=�x��S����'�d���'d�'���'MRV�)�w��ǃ�6xaP�l�0|n���d�%�M���?a���?1,O.���O��$�3B�nrO�t-J���d�b�X{q��O��$�O��O4˧�?��վU՛�РM�L�׹��b�eV4�q�q�i#2�'��W�p���0��'dX��I7S���G���<���xc�{�Pmjܴ�?!��?Y��?a��NG�];Ɣ������.��vl�&JP���Lv��7M�O��O�d�O�5��)�O��'U��R�X�Fuqfhϥj���H�4�?����䖿v��%>Q���?�R��Q.��=�4�nUh�뵋Ԣ�ē�?���8�A����S�TiXq�����K�.0 )5���M�)O ��`��1J����������'����-R�>��PD�H�"e�ش�?���EA����S��(�T�(0��� ��%��l%�4<�4�?���?�������)@�,��]�#��+��,�E�f*lZ
Y�q��ٟ������O��'߮qPB��+�zIy����3�D{��~�"�d�OL�d��O�&�oğ�O*2�O&	�Al�``� /R.�,��i�r�'�a�$���?����?��O�r9�f��/u�^�A%5%��x �4�?��a(<>��ǟ<��ܟ�%��X�)IX�r�Bԍo�@\�T�E�v6-�O��C,�O����O��$�Ob�D�ON��X�2�414��� �f4�  t�l���S�Iş�����'b�'���hp�.g����Ñx3pɃ�	�^���I쟌�'bcפ��)�K��=���W0�HLA0�\�4���'����OL���:���3.���QRH�uI�	,��O��d�<����ă*�R�dB���;��GZ���i���4.��=m�q��?�@ �-�<1V�S�Zd �:C���sv��+.0��'K�	ş`��m���'���5����.�~p���#���u��9���?��#L�!�N>�O?� �-�uM5gQ L(�bX�{팸RFY�<�I�O��!�	����I��SryZw(r�Ҧ����X�
^�m1b�"�4�?q�!(�<Y�� �@�Vջ��#<4y#��b��V(�>}���'>R�'��4]��'@�B�cp�M�!����E/�8���ɱ�i��ɑ$�|�c!ҧ�?�pf�1�]��P� Ң�Q'8����'p2�'�|���?�4���D�O:� �>�,0�Nٳ@;(|��%M��5��ş,�I�|����.ʧ�?��'�j�S��U��a���w�.Upߴ�?��a\����{�T��GK��D	��_�+�\9`��Bd��o�۟���:�I۟�	ΟD�'�`����*;uk:Ԣ�2�%�<JO����O*��<����?a2�Ҙ-�r�Q�U!BT <
��M�IN������K6���x��%�ʓ��4&\f��D��̬#�O9�B�	�M����b��-�̔cT%ڌv����2F�[\�L��ϔE`v-9E�& �H�[d�!Wڴ��e ���"]��!I'
h� �Ǟ�Uhx�0�рa�4aKz����6��yu&Fr�$A���azl���;5P��{E��
�۔$�4�ؓ��N:\,�C�� u:�8�$��6TT2�a�<t�8t��O��ړ�8uT�ֆ��2[$�	qi�O��dW�\�+�aM���a��U Bpt���O�S�u�\���Q�#/ֈ�EA	;i5�'�0(B��V�����ќRP�S������O�B�b2�ؾn�pت�n���m�N��U��O�doZ��M�����OT����#:5�H#c"�(7LM���|��'r�'9�	Ο|�i�EjAh�u� ؇��db�;Z �������ߴ�?���i��a
D�<�j��ߧFnX�@OC( �6-�O(��OjiE�$#��D�O���O��0X���{B�7u�a�&Y�(n�����է@�����B�w����%��Ϧ�*��i�h#LA�ONܙI�Ɵ�Eh�(��Y-q����P.峵 AOS�>aoZ�{<��I4�N���Ei{�}aChߙ�$��4<��ɚC���4�j��)�	��+�#	�&��� NH�M*�B�	���%�s!O�`�`��(��i��k>����޴�?�.O�0	���:���i�N(x�*���_�Ƚ����OL�d�O�����c��?�O����
�3!�|" Ȓ9 O(S�h� O��0
cE˼0��!*ÃL.U��#?Yw \5H7�r��l�dT{�CY�F��łtᖻ,��u�,NTr�w�ɥ	��h�1�&Qr��3c^�vҮ�0d�O����NM�Pݨ�\Z�����:)!�)�����mт\�r��p/,r�1O�d�>aʒ? ��'�b��y��Y�7�?W�h͙2�ѥTT��'��I��'NB�'� �*X0j��]�b��mZ�7-�*-��T�ߋ]���ش��x����H�1�4Ô�W�N K�Γ5�TH%Ɔ)@�.	��G�Nr��G�e�PGyb�
5�?ᐷi�6��O��e�:������(_����'�<IW�i��Ib�T��Z�AZ���*� ��M����V��Ӱ�p-��i�(z6�W�f�ʰ��O�������MKQi�>mt����?���:�*�?���N�\&�Yҵ���un���Β�?��U���{�fW�{�"���	���M��~�,��:��J�3~�3�62	<�a�>����8m
��c��k�Z�l�o��nެg�� �c��W<�ȓ��]�<0�'�ph���z<ɧ�O	��qGY�3�8���ڡ!�T���'`�}@#e�	t �Qo�$�!�i>�"��@F������ʐ(C0�_rmZ՟��	ߟ��	.ir�|����������݀Z��8���^� �Se<�М���ZDD�oڟqNzx�v���'A"�'� i:]�����Oȥ�@At���f��j�故�M����������i�$IМ'���r$*�,j�ݰ!����i'.y�P!�'�������͟"�'��	��� i�����y��H�g����˒X�.�Y�^6RΨ{�ND>5����O��'#�)2����A
\��(*�hY4!� �D$;\���ɏ'���D�O��d�O�,���?����t�N?P
&�BՄ��l�0���Wtr�"���u��4ɴ�	L���"Dm�zں�-�B��g�O4q��d+&LO	s~�CS�г"���W	ڰg*�ȡ�'���!��;7&i�6Yâc���yb��	�@t0RAW�
R���d����'�Hc�t�ƪ�M3��?iC�S+6�t��&�)CN%Ӥ��"�?��������?��O���2�K\?����8ӛ6�,�v�+��U����%�p<Q��	'2��
ac�9#��M��40��pn�P����A9�a��	�<3B�d�O��a��z��^�U>B����O/ET|x��?��������̉�o�R>�Ċ`]+M�\m0�O1nں < p�ΐ9u�*�AүV���Yy��
�E�X7��O���|�@\<�?�D��,-f�����IV�ArR��?��eRZ�;�Ð�7d���g�Τ6|HX&W?=�O�Fm��'M�b�b���K@0>E��J��S0KӐYTp�s"��&l蕪Ww�'chH(�eMFȘ`�C1f��O�1C�'�"6MZ[�C��{����v��t浨S�V*Tvc����I��T�S�? >뇧[�T�������=��dۆ�'�<7�ʦ�%��Z�$G�dJ2�\�0�,��΄=�M���?i��&���a�.��?y���?��Ӽ�ŏ'h%���.��=��U���S�V���pᢌ�mT��	H~�<�&�ɧL̠P�f��]l�`4�]�p���NG=^��%�B���}B,ʸX f�	0%�����j��U̮�r���:j[H!������v`����?I��C*b�U=��9uD7qu���}�O�R���4{
��A�}oh�ӛ�|�4_�v�|ʟʓ]��J�c�\�:�
�=�
��@
���p��?!��?�պ��d�O��C�Q<YBD�w�]K ��`��d�l�%rdN)x	��3�2��˓m��R���F�*a;�^�B���� �W0%aa�w>:J5'�'K�B�@3T� �pn�,��5��nת�?q��
����'������?9d蝌��lSb`� �?��?)	ߓ{�A{�E�I�LU��UV
E�O>�Q�i��6��<���U�6����'������m���'N��bPl�t�b�'���"�'���'��s���cUk�k�%C�7�L5�Z\H%a¯P:� a��Z6S��x�Y;��qA�{��պP�O�0���`B�F�@��,E����퍴ȈOHb��'-J7����I�z�0d)r# �2mS^,�|�'\@6�1�	��O_��A�ޞ,&�P�ϊ*C���
�'�x7�O�}A��*�FS;�JP��T� W"n�z�	�@��[�'�@EXf[�f%����rUk�'].�q�肊_)'*��K���yB�BJ���������� ��yB�A�4@^��D�� by�� �y���GD�Ʌ�P;]䁓g�H��y�%�R����bӴ,
i�iCf�<�ʶ?��x� B� �ݳ�Nb�<��JT�t7B�	U���J��!u��a�<�$��h�)�&&a����LC�<��%	�`�dܡ���?,��0�|�<�UE�M_z�B��0W�  �DL�<��ʕ������J/ �9����F�<iD�ؖ&%:����ձ6N¤�%�F�<q�#čc@mH��_�B0����k�<f� � #�*:=��T��y"b�>XNz5�C!_.����p����yR`�##J�����<=Z<990g �y��Հ[,lI���3#�V�Q��L�y�`$�,��4�F��
�����y2��l�h�
�2z��N�y���,��3�A�\��d��y"/�Eʀy�
��Ѡ�[�N�"�y���v<���A��2}ĴAi�ٖ�y�c�od���c�"o��X�1��y��\�&r�(�S���B��y����	�H`R��чL?Ԝ{�o���yF�d�D����$DB�CCJ�'�yr�ڤ��E�g �9{�oϕ�y�g	�5�ba��O�]�^�u�P"�yR/R ��8����`Φ�*�ۄ�y�-ف����V��D�8q����y�*�%s�❓�hZ1m���;Dh�1��'�� ��4y,�9� |l�4�F�N5a*�ͻ��O�(!6B�	�R~�bqE�)�B��֪��2Q+��G
V�$����O�����3?1��³V��qb�6��Ъ�E�D�<�B�u���v�|e$ #��hT ��U��>-G(=�SN2\O����!��9�lJ3>��t�v�'V�k2�	?7�H��h��fr�{V���
�)s+ٰi�<d8
�'�\hx�'ַvۖd�AA��_�6���yBI��6��@���W�b|E������R�Ý����� ��y�- &� L�7obE�f*c[ 2e
��O@�}�pPE��O*�����V!���"���hI'"O����n8B/r\�w?l�|J����?o��!�*ץ<�p��
��~塤j�!�K��X�lY
�鉰@Ҥ�w�A�l�����#�&oN,�P���3��у�(��Z׺C�)� ��!��,&b��d���1wƴjV󄜇q�ƵhR�	;��Î�)áx��(�q���?�v��R ׅ?!�DA>z���q��ˡ�EIE�S���,�\!�v����
tO,�g~��LKaSC�,(�J}����y(� l 0�ڒ�[=�����4��Èmh��k>lO��84F�e�l2#�J.����'�r��DHE?�ME(1�nԳ��\t�ҁ� �Mu�<� ��Ci�萄/ͅ?����l�'�p��	�W�g?��,�Cېي�ύ�6��Q	ȞM���3�Ov��N<&�ܭ燊�~�P �Aca$�a�����c�Q��yg@�6�I��@ܧ1�:��շ�y�i�1/FE(��L,ʠ0l�	��lJ�2T�T��s�q��|��dU>;>d@h�͟�i��D9$�'~Lqb.�A?��Gڇ�^pq����#��E�������'S��UH!ϣ^��3�+�2��ɉ�?�l���"ފa���'��!���F�iaf�5������<��bK�E8 |��GR9cY���D��P���X��'$�1�D��"��"��A��2DJ#]�4��A �<)�����Tl�i�AB�D�k��,"�k�5��%z�0�O� ��֩�Nت$FI�zp��������vAi�㔭��Ħ�T��u��SV�<f�> c".�<�`�/�V-�T��&F�6���&�e�'�y��b�461���%v�,Aܴ���� �:�x��퉤.�j����/���3	�>�h7�ɸG���	�R��DU%S�Q�t�bt�#J��j�� �k̃*d􅔧�s�l�WmV1b(B�Ǻ��L��V�1Uf����r�=�%��a
��"2�K%�ܰ�$�"ތ�'P����D�A��	�<�$c�`R�-<ՠ�`
�H���#4�{ŁD,ty*􆜸Z�;C��W�H�ÆH'��K}��;2bj��P,	n�$��<�Dh፞�l�x%J���&Z���[�-R+/t�d��#A�]D1Ӗ�d��Ӓ/�?�H���$�T�"�0ěx��Y,h�$Eze�ǽ5���ORH�'�`hc�ƀ�L����fK׾0�*	�,O2D�sË{�� D�XZ�3��O��>ɀ��Wk�hZt�ם�
�ZQA\�<q�n����DƪJ"2eBem4�k�$l����؍�a,t?�p��C�Lϊ��C�͸A��@�Ǻ'�d��<���Ы.=dO�.rrĹ�E��j{����O �p>)�.�~o�	�%N&�^aȀ��ay�C�:x�ÒSf�
�z���<;l���4GR��ܘ��ƈ
%>���d��,�<�3#!�1U�|��c��0x~A��KS+sEN�+�E.\��'�
�SU��0|��` ��hPxhha��	5%�	���6"����<�"����-u��h�`�l���&r���Vo��V ���'��i:�}r��J�5ruk8:�-1gF��WN0�F%M7���"����v��
�ўP���ۂ_L|�r��ɁW,j�y�C���C/ax�G �*>��A�Í5�@���e͌JC��?{t��[u�l�'��ͪ0�^� a`��C��<8�r���"���K�.A2A,"?�����Ŗ��W�VUI�fi>\
 ��B�rƝ{Ć�`j����$��-C.- �ۦKI6�s�;.\�'�j�	��1�^Y4�+s
��z�O��#�lw�� Z�JVtB��5�b� saF�o��䈘^/���*�*f�=��B�鎉���?!��`b(�#!(*����4B���ئ��K2i�0]�+A3d�H��eJ �:%���%?p�5D{�e	5#ш"��#O	 �� Ɋ
dܖ�O ����*�(�����f8"��IK~(�a�yB!�`�B_ճ���"1��њ#�1"��8ò
$IȪ ��+T��&Л�@l��A�����TtI_�K2�_������
�Lm�pۮi�D�"��'��S�@�+@�*�0U O�%��l�J<y2��)@&�)��R�{�I
RӤ ���6ϦAӅ��6/���aZ�c4u� ��s#fm�!��d5NCK28�33������<5z��ʘ�A��S ��C���!U����0?���[oƑ���Za�p�TN�~Yp���n�zH�I%���<	��GyR�˩Y`BIa��[\l����ȵ��?�r���3�|H �z��ju���'�Hy{�Lʗ1 1�C&NJy����I�[��<�AR�DCFq�H�k�Ԥ��'��@�1C
N���I�MC���)$a��+����|�!548��@N� ��AS,*�џ�J�b�'v�J��0��@���C�m�>�SBŦ	���H�|`+O�V[ᗀ��� �	RC��p� 0>�(��DN�|~�òɢ`=ۓE�&c5�	���d�Qy�m��<ٗM�<Ѳ(�d�0(�q��h0+�i�N���Ҷ ��Q��Z�O�N��EZWn��%T�ѕ�ԉ�6OJ��K<�S��f�M�*���PM=�5��.2[��'�Q�PM�|�"�D�$\*d��{R*R2n��b?O|Pk�j+��A��D{�]qqO��� n�P/i��|�����X�se��KuR���Ž/��u��遺N��h%B	�ay��#5L�'�� U(͢b��Py� Ԭ1#��4�;D��C�ċBnD=2�^%p�u�@�8��N0����>�����%T�P��
I�XM��9�!D�pA�6:��j�<n����2D���Ф*����@�W�`���N2D���\�l#�8��LD
8����`�.D���a@'� ��֬� ,F���+D�0�k[�vsf�	�J�%m�B)�V�3D�@)U�ݻ|���C-ێO��[P�2D��)֍{5�	�En�0�~�j"2D��9��Dtvp�V"�BpS4�.D�d@��[4-؜��Q�I3S� ��g�(D��CU+�<1H1�VN��3��] Dk&D�4�rlI 5(��5�1�µ��#D�4X��M�b��AcnFeLU� �!D����M	B�@t[��+�ܨxe*!D����I����bG@���H%, D������tuVL�P��g��H1r�>D�tcaˉCe,}Q6�KI��S.'D����&�`�еqVa^'Crv�H2b$D�LѢiݎ^���LZ�)]N��k#D���ԃ�Aw��	"AZ.'�)���"D�\C�1^�
hH�#ͨF;�9aB�;D�xCgDdxI"H��<\A�vj:D��(Q��U�����e�-|�t�Y��9D��Zj���e�4>���� E��!�"�D�� �L���ْ!��>k�!�ĚR���Qw����Č/���Ұ"O����Q��B�#bC,��H��"On�	��Ū��i����j��	��"O���27�ᦀO8 ����"O��j�h\�X�8��M �SR��p"O�@:s�
</�@��k�,_D�r"O�XU��7��;S�ן�6�1�"Oح����c���B�v�.\��"Ov}��fm���R�?�)s"Ox�QBHˢ.��tP�����"O*���H[������)xx�<�"O��Ұ�_�r&�4���˂\��`"Oހ�n�+�� ��J*?D$ ��"O����<Sa���_.9� �"O@@%�L�3dl�A�"R�>��C"O� IbF��Z �L �MbFH��"O>�y� ����XS�_xX�1j"O*<zs%��,r��W�<F���ӷ"O$q���$P��1# �7�� $"O��eֆgZ�(q/S�*���X�"O�94��K���" lŚUZ<=z�"OvY1;�5��`I���A��y�f�\�@��R��g=�����R��y��T�`\�E��,�9��Ê�y��Q9W�4�r.�$"�労��y2��8H˸�@*��ȽУgܯ�y2h��B� t[�'�+� �(���'�y�Ċ�|<�ш@�&��dcR���yb��g�J�b��N�{b�ŋ�y⡘�d��aZ�6&t�qo_�y�+ko�8�愀Q_���E�W��yeGNv��׏�Mq(	[5���y��.�he�ܿK�ո���y¤��nVpٹc+��B�� �U��y��� ���d�n��2�H�6�y
� Nđ¯ۈ7��z��ՠw�}S�"Oޅ�j��[mR�(�$	vh��"Op��e"��A�H��a�K=cb�JP"O|�k�"�)!���i��Гp�`���"O���)�s����P/"�)9�"Oİ��?$�Hsԋݤ$X���%"O�<
0��i�$�	�J�&~:����"OPl��ď�*5�P��L�"*8���"O�c��ћ�0]3èG�	�ڱڥ"O0�1㒴bdP��M��P	�"OJ�Hf�l�,��2~ࠣW"O���(��l�z�n�Ã\k���"Ov4!��
B�c`�;<f��"O�%��a"t9Hu/ґW��M��"Of@�� U$�D�FV{:�X%"O��K�a��y��8�֭AUq���f"O>�{���u����,فa�� �a"O ��5OΕ7�Y�	�&WN$!	�"O�{B�
5h������!0�D���"O�e����	G��a�"���*�"O�h�wm�"s��t`BHƦP��"O��*�˕0��|w��(~�BT"O�����}��(��4J$ Ȋ�"O ec���B=��K�-z�,*�"Oܥ�6���w���Q͜�Co�PA"O�%�B��۬� լ�37���02"O�<P��\\�������)6~�aC"O�p�*TTMBPʡ*�vlD#"O�9Bf�ƿ.�P#rI18vFL��"OL�s��R���E)���u@�"O�� ��)�P�� Q��$q*�"O8�#�L�`jL�HegHz2�S�"O� �D���<�P���(N]�$;�"OF|!J?bu�I!G5S�Lx�"O*D �*�:Og����O�K�b�C�"O�hc'��?d�Ȉ���D/J�&�s�"O �j�G	;.�E���=V��@�"O��+�I��XQ.�sR�/<�%�p"O.��VÌ�F���a�̷���ʷ"O��� R��t��e׊U�$PC�"O,��a�72�0��jN�}��"O�a1@�DZ\ak'�X�H⬝*�"O�S G�@�@H
�E�v�<��"O2p�u�i��)B���"O�m�\�2�i���fm�d"Od� �;ގMS`��
��t"O�8U��>&��P��{����"O��aQ���[����hA){�1�6*O�T�c.�$8U�����$u+����'SH� �X �������a��'H~(��I�Dfv "SÞ����'l�!�gƟn�ѐ��MZ�px	�'_���g�Z�'�<a �`Z'���	�'�qp����O�d�W��6}B�Ъ�'"��Uk�;q8��7ƞ�*ld���'��Z#�ň)��ңE3u�
5�'vbDy��4=�����!� �i
�'9콣��ƝB��X�b�މ+�U�	�'l.�r����E��3	 ���'~���(Q
=݆�`Ҩٳ(�ʜA�'�����5EB���ʿIxZ�9	�'FX� ��O��bլR6=e�d��'��Ԑ�L�����I�"L��ة
�'�\U�QB1fH=�$�Ɨ=�H}�
��� ��-[�pԈ�h�H=�Ԙp"O�[�ƙ�v�j��e�* .9P'"OMr�hՉ><`�;!+utAC��'QqONL;0N��qX^q��*Цlp�F"O~4;��Ȕ�C�*\P��@"O䱸v�ñ>��� в]H(�ɳ"O �"R�JM�t�@�$\+�i.�!��g��ˢ��'q�� a'�B�FL!�$E�t�\��h�C�r���΋�!�$�"'Fxhkʷ�`����=z�a}R�>�T�o�6L�-Zuਢ�.�[�<��ȗ�N�h�*�P.���oH|�<���ܖ�\P��N@  ��%��@�<	g�H:'��C��ي*�X(�'�@yx�$Fxr�Z�o����i�
��Q�Q���y���zw����ۻ18~�r������"�S�Oq�@���_?i&��``�4�xC�'J�dp K�66�^�X�	�.�	�'�p�8�jM�*u�v���uD�	���~rkMp�Ƀ�H
g�&��V�ī�y2L LPfyه!�_�<pXF�Y��yR�2R��1��Z�����iY&�y��H�c\¨:���J�vq���F�yB놽2i�� ��E <G��8$F�J�<q��$c�<0z��ב&S�I� ��o�<�uN���Rӂ��qy��P��E�<ق�ӓc�.��
��f���i�!�C�<i���v�H�h��X,ku�y��W�<i����`����86E9@�O�<���
.fe�t�&}���$��M�<)c#[�zc�q�.Z7w宵`Ј�Kx��DxB
_�W��+��^_�T��n%�y�	0HET����Xn�|�`���y"�R�r#P����1V�,Ey@�N��y򥀣`�iBS���RlT�!���y2�Q�R�Aq�m�`���Wl	��y�M	�x-xU;-��^Ԅ�� ��y"ʌ)Vn�y���W4�����yB@ʳV�����OR�fU�E�ߵ�yB	כ&�V�ؖ&�D,j��H�y�'Y��"ܹ�b'C}Z0q�n	�?q�'�^ r�˗I�xd���ط&�Z�S�'@6$yF䂜t/�aK�IU"<m1	�'s�e����X�0=(D�^@'����'����_�]0$4Г�>��=ˎ�$>�S�$�<p�܂C�7e
�$���I��yR@:��{E�5c�bmS`i��+vў"~Γ/,F�+���	�:3�@�tF��ȓ+r� � �*U�P � ��:�PY��6�37�� 8y�k�M|,��I^�I��%z�"��R�L�M��bb��x��󩀎?<~�P�m7����N��?%!�d�8-��E:��:$���Ƥap!�F*t��ĳ��O��9u�!o!�Q�D'.[�O�>6@iF'˽cP!�D��3�6��ԏ�_%6�yf��:\!�dȩ0�v� l��T�9Z�!�X�}"��g�ؓNvh�	�	@�!򄌇1hH䧗�ewQ�('*�!��\Np ��ܛ^��*��C�b(!��9r��h��z[N��u�Ӭwj!�D:[e`��T�&%{�\���9"�!򄘾[X��aw�Y�ft����l��!�߁+��и�˅�>iQ�&ɌV�!�� H1�q�^^�LT�hʑ-�)�"O��K��(g�N���G�'�T �B"O�����Ť he F��!"Н�S"O"�XL�z�t49�E't��"O�c�E�0l��3�MV�|�l�3"O6��
�v2��MЦG��|�"O.�a�ؒEd��� -@�Q����!"O�`H�&�$=΅qū嘜�"O2�KŇ�,j����*P���T�P"O��!"�
��33�J$O��Ѳ�"O�q ��.
Z��r�5�ڵ��"OPh�b�߰Z�! ѶY��)@�F?D�tƣ�0"�2�ʶ���*�y�E<D��8�	ک ��1�% �@A%D�����;l� ir�A�=��l�cm?D����$�r� ��M�:Qc�*2D�X!���7T�B��s�NCB	S!1D����cƷq���P��]���P�1D���ܻ�`E[5��i��YP��2D��"�!;��ڶ�X�	���r�>D��!���9�H�bu����0D�̹D���.�+�
��δce	;D��3�Ȟ�pgX�`�&Z�%+T1jt�+D��a`��N�01�,�YL@;!4D�x!G+
5DM�QJڏO�R=
��<D�ܚ�ˌTTmR�Y0�j���-D�d�dCͳښ� UǗ!f�z��&>D�X! ?!\��C�F�m۴�KC+9D�,�E �++
r��$#�� ���J7D����"K�n�e��W�"$���3D������`�r&�W9���k1D��9�$�##���IRA��/R�B�"%D��! ��<*3���7��<��ȃ "D�`�� 9W�uq����se#D��k k� M��źTA��4����6�"D�|9Q�N���(��J�~2�!)E�>D��Ì�u@���Ћ�3���L=D�x  ��p��h�D˖%n���R�;D����j#9aƝ� �T�Np��)�B;D������~t�ff:{UXU�7-=D� 
u�	�=�1[S*ڴ2��x�1K=D��Q��q�<�8�f֑O � �e�;D���J�yw�u� ZwOڈb�:D�ȱ��>��{�v�t�#��9D�t ���:VWBq�a%�]�\���5D��1k��T()��T# $j1Ѳ'5D�$�F'8nR�9�Q�&����=D�+���u����"fU�$��+8D�@�"Y�O�TD�#�J7 f܂%�4D���NiÆuȥ#ʞS���ä1D�X�У��V�2	�g�ܐ,�$�!qk.D�$��LYgDd����t���
TC.D�h�bJ�u�+&J�>���RF?D��1�
U��X��%3^P�8��<D�;�ÿ;(�m�/C�J��K��&D�H�ځ02:���ʞ�Z� !�7D��S��i^ġ��"�,�k�`7D�D�b���p�H���=~�a2b'*D�X�Dm֞"UHă'ܚ^te�`a5D��I��Y� 0�Lڵ/q^�r��%D���0-�
	�`W�L�f�j�q�5D�T����9R iS��Sh8�3O5D�l�f�]�옉!���!� !D���`˞��24'ƹP���uc4D�� �E!g芌5�m3��U!u].Mkb"O<�"���f��p)YT=p=��"Ox��.��aٶ(��C�n5�b"O�����90fR�a�g˪3:��"O|���S�������%��j�"O6E�%IE}���cD]�s2"OJŊg+í���	m����ƫ	'�yr%�W���ʂ*�)iژ\���
��y2L0Y�f�1���hC��׈�y�I�XWy��^�]����`N��y��ɬwT�E�Wâcaj�b�R��yR��/d�\3 BAEa� c���y��J�L�r	�)K����b�V��y���*g=�0�F�L�~����E��y��ʉlm8�9uMĚ}� ���΀�y�̊���ʠ��	�Z�S�6�ybiwr���	���������y2�\0/�n�����>&���צ�yR�Y�H���%"�4����V+�yR��f�9uG"��I��L��y��u`�}��H��e�y��W�'��h��/�.+fP9fb֍�yb�B�m��@+R�v(x"�)�y�,F#�X[���2��<Be���yr
̎r�J�8gS�$T�<`"�˅�yb��0qXt��F2"���y2�L!�dɻ�ԧ���s���y���h�Xu�"g�%A�Y*����ye�61&����(w��kU%C�y�K�"kL�� f��P86����y���9%& /$؝蠀�T�L�	�'B���&��$�\X`1�M?J���'���
�'ӵ$ڡ���=�\I�'�ԙ�D��n���c!��/��!�'��E�T>Gp��3@����ph�'x��-D��"�0�bР����'��1%�S� �u�îU�rD,|p�'�L��d�H�A��`�e���%�v�<Q��ֆ1,Xغ�o�:u}���#��M�<�r��9,W���&fL�< �,A���@�<�%^C�x�XL/_��l0&M~�<yvoR�1�p��`U�3)hI�R�y�<�(Ο]����T�ϮQj���`Cu�<1�ꄛbށ��A�h��Ɋ2�7D����a�>l��X4��?�b13r"7D�h
E@�-3������*8\�2�#0D����/�
}9��b!�O�,%0��8D��*SK�6j��SW͒)4v�r0�4D��&����ĨZ��V<k�<s��3D�(3�ES7V
���g�*b�lH��3D�`���0�F� =�B�ǀ{�
C�	 >���{���`q�8�`F�N�B��} nM+���� �|���� ��B�I0�� 8c�$;`���[-�tB�	�w� �8Dhօ,Y2m�TC�)O�tB�IˎIS�$K�Z�B}P�	E�o|�C�ɫFu����A[�@z}1�X�0��C�I��I��a06�Z�`s��@�HC�I� ;�M-w�|X锆%vTC�-<�^Ԫ�k��]-�Tb�
�"g�@C�	� �����)TnD���n4C�
A����]'�>��#��y#�B��3h��ȘCB�O����D�P98�C䉡��� �I�#x�U���!X�.C�)� �[=)kj)�G�3k��(��"OX��Rt8jl�`�E8,)�"O��T&NE�PE�կN|IJ8��"O��ՀB�H���`���"OPy��S�eG�$�l�#]R<�f"O\R�S��jz��BVF̵�a"O<�B�"��7`�P��d��E+�"Oʝ����+N�,��co��'�p!� "O@P;,ٓ[���VoI�F�8��q"O�A���Dh ��A�,ǜa��"O>����/ZN�P��$D�|Lâ"O¬��� #��p������"O^� �A�;�|ͳwl�4uf5`�"O�@aF� �l<���Ń`��Q�"O��F�֑a���/T�|���w"O*L��-^�������S�bԲ�"O^�Ebw9�-�W��*6��M�@"O5����b��U�A��}z1"OH���,��@3TE+���I�"Oa ��ĳa�t���F�w����"O~L��"��>\�9����-0B  "O͛��	�BW��"B����RaI6"O�t��BC�,7Z�QQn���[R"O��ný���1���4���ZA"O`�ٶJQ�^8
m��b�[D��Ё"O�C!�	���x���R/-�D4jv"O<[�%��J��V@X�.�V�Zr"O�5L?lX� k'AO��
�h0"OY�r�� �h��v��F��x�"O:X3X�¦���`�HLu!�DR�X	FM�)6���se_$lb!�$�fk�@r3ϸglj��d��L\!�=$(`���@!	1Z,(p��2jK!�@0��7LR�t��{�c�(U@!�Y�n���d@[���uHS�\)!��?l�Q�b�G�����NH�!�$ׅ�,%�w�.~���Ҡ*Ҵ@�!��ȼ"(�ٷ�]z��8a�̉t1!�9S}#�ˏ�0�@��&�!�d>e��A�A��,�����U�!��%Q��E3W�]�K������j-!�d6�v�aa���8�N�aC2!���pX�L&��
N�8(�"]�O)!��w"V�#(���``�(
!�Dݐr1,U���k�t	���"�!��W��	�&ő�>S���;�!�Dǲ8�"�E≯R�6x��ʗ$]�!�$N�1����b�=2�\��� �-�!���"�h[�ڦ:h�C�b֓4�!��yZȘ��K�SHμ:e�ј{!���;�D�U��S�8I ���-0v!�[)-�&��0��7K��E� H t�!�$�3e����[<��d:3��j�!��7#���!�%� �FCҋ#�!�$D�q/ĭ�d�(�ذ�b��-N!򤊼/�(a��Ԫ�Ul�{0!���(�(�h���l+$��AL�/8�!�DZ-*PPx��,Y�(E����lΣo!�Z�^AҲ�3
,�8ȶ��k!�2@�t|���)+����-%�!�1EЉ)���*�h��On!�$�*k�Q�S#{�$�:��ىia!�U&�}����f�%���ЋU!�DH86��X���Y;���ѕk��+N!�� ��#��q�:��C*T#X	�t"O�����߅A�d��a( �&�)�v"O��@��z�>�: �R�U���"OKǈп(�rHh'�=�pe�p"O��Z���Q�֬8!k2(��{E"OD�9qR\ A��ɛ�1#T�� "O���Ĩy��c����R�z�"O$��:XX�Tر ��zɈ�"O�����}�H�he@̴8��0��"OJe9s��)�,�zB��'>�lՓE"OHS�畭����mO%
��!�"O�-�Slܴr�"܊��I��� ��"O�ԁ��)eR�J!*v|2�"O� �tC�%E>��r��ɠ@�*t��"O�5eG�H���)'nQ:Eg��"Oa�A�^l�˂ `. a"Op�W�+r1�Egj]m���"Oڕ�@d՝M�(�"�o���"O��PENƱz��9[t)��$� ���"O֙	�KG�H���R� �0,��"ODx!�*��Lv �� L�M���� "OV��6��
�����@�4�k�"O����BȤS�V��0ś\�����"O��[��,1��t	��LPu"O�{���Z��+�A n��5"O���c&�=��iQ�`��?ȮMjs"Ot��3�?�0�I�3Z6�[�"O�p�A�z�Fm�H�LA6Ո�"O"��N.������D7���1"OZ Ԁ�H�.� I�4��4"ON`!�
2'?0�Qs��:N-(t"O�x�WJ�j\x���OU�?�D�%"OT��Fmâ@���r��M(=�\�D"O���2@�=0eK���e>��"OĜ`�N�vdXrc�k�0�K�"O�բ���."�YPI��66M��"OQ��k[	r������x.�0�*OR��Tc�=5ΰ��B�B��Hu��'��vD޼58�s/� |M��'�j�RL���&�2&�fzؓ�'���� +ϥ$	����@D<m�d�{�'s�m@g��%\>Pd�'O��Th�$��'X��E�h�a��툲>�Je �'s� �@l�[�Dxh!�K</��0��'x�[�p�И�S�$�
���'F�<��ګ�$�0�&��d�P�9�'� |J3��vU�����)��j�'�z 0��V����htT.l�8qi�']�%)��D"I9�)(�L�r�,#�')��ȶm�d�|�bcY.��-h�'�l��3�^-f^-0�o��P
|�z�'��	9 C��,��!�M�V��
�'Ҍ�0�LŶ^��h���>> =`�'j���BԼI�l�P��9�6�s�'*Zxb�hؑ?����	NV�M*�'��<c��ɝA�b1x�#ȄӚd��'l̠���$l\�Ц��%b�*�[�'��@�Q�q$x�+G�R�"��	�'v>���'�@\[v��v�� �'�j���I����кb��<��'9�h	�+;,H��A�'Z���'#�3��Ӗ?�P�k�Â
MP8Y�'톙���کX�聸s�IБ9�'�v�� �]�1p��9FK�@���� T�s����:����ƈ�
�8�t"OR�sD���7����$ߘhlr�(d"O� "����T�0YbuDBR�$+r"OzȊ�GK������57.��1"Od)x��G�+H�Q��
�0,�~E"�"O �����3f�ph�����-p"O�p[�
	f�]H1��o�z"O~50��J�f���zcM�lr^ͨ""O�}��o6x���T�A6�1d"O �{��D��yw@��0�"O��"�ţ@ � &����x�1b"O�ХI 60�h����Z����B"O(t[��ܶ|*�3%���nq��E"O��`�W�B���E��Q[�t3`"O��x��A�c�B"Ӓ]U�  R"O�mqEb��r�X��Dk 2Ra��k"Oƥڄ�V/`:ƥH�I�V��)�"O�9n�c%��#d.�'^
 ��"O�x�d�ơ��!���Y��	�"O�� �"�||�S�׻:��Q�"O�ᐕiU:ZE��.�
r�8�v"OV�����>��1�8^�a) "Oȁ�H²r9��I��ҟw,$)�T"O�	��� 0�D�҂X7˂ �"O4� ���05��BE�=��}KQ"O��"���YU�衂!K�l�(���"OxD	�_�#������8~R�{g"O
QaD�Ño����><�&�y�G��M^��P���ub!�梃�y���!�^i�2˓*r��M ���y��C(j�6DXvHI_n�|����y�N.e_�8V�DP�P��퇜�y��J�C��$�@(M)�-��,̲�yb�D�J���A�87\DX�I@��y�d�!V^�M*FB)3l�Pu�H.�y���O�QS6l[�*-�1	U��y��,/�F�� 
Z��J^��y�)�J�c���
X����E��y���;�đ{ġ��	�H`�ȑ8�y"%Ϩ_��a��X�1�6���y˟%�>,��Z�.`F��U�\-�yRD��'�p9��٫%��9%�Q�y"+��n��<��H�
ٔ�:#F�3�y2���g;>���
�)���yҭ���yB�ޱ<`�����J�����d߼�y2�ʁ��Hƭm�d�b��/�y��&4��IC�ÒP��+'Û�yK
S;���Ǣ��!x�',��y��@:VH�@ � �|ܾt#�*���y�"��H�t� &u.�R��-�yҩ�'>��!���]	R@s�����y��9wK�<���0H�z�v���y�(���"�õ�F��P����y�6/��q��Ռ�R0([A�'��:&iU�KD��`��آ#,�8�'���� I ��tj��' ���'�nT���ݶwlN�@ڼ9N���"O�m�w��e���	g�+] �M�"OR�)v]>Ernd��	��P�`A"O�(gi��q֐��b�7Ԧ\y�"Om��H�I����aͪWi�"OʐkSm r�C� ���pq"O�᜙a?�\���	S���"O��s�
JxP8��'�4��a"O� :qq��L|�	����d���"O���5�r�b����G�i����"O�-���ʄR Iz&�Z/QP^1��"O�� Tk^�C�X���W�TI��"O���P�K�8�8�a%��!ڴq"O���@@(7����W�<��!�"O~�س*WF�p�	6��d��L�E"O~A��$��?�����!l��X��"O�|j!g��0�yc��g(� h�"O��
d��ke&)��`�<B}��"O��S �#����G`E-I�t"O�l�ӇW��d�ʍ?I�0m��"O(q�&�)q�Ԥ��)D�X�b���"Oz�jӦZ�9>DP�'X� ��d��"O�Y�qdn�R�8��ApT��@"O�AqC Z��cRu����1"O��)�3!0�̲� ��r֮�Kb"O���gG4��D��òu�Ո�"O8\Q�%�>(o�8ӑ�Tj�Y "O�I
����v��(�y�׍�!���hTkЍ�!j�:M9P ���!�´5�X �Ձ"�^1�@	
vD!�?h��c���;B*%���Q�!�d��>�9��Jؚ+%:��%m��!���.�����{!�q3E��4�!����|�P�Tl,�"�HT.�!�D�1�U�DƏ
LΨ��gLR����l��}1e^�s��A��B��h��|t�w�4T��5�
�i(j��ȓ ��bQ�z;8�d�$Ae ��ȓp_Ʃ��EL���ՙ�m	���	��pʐ���ۂ^�Q��jX*�����e������25���u�����lt�s��M070���V�D��؆ȓ~Є���a��!�(T�#炇��ȓD�<B�Al�B!�W5P�MV*,D�����V�zS���`kW�}�XA�*D�h����-���l�/K̤q�vk'D�0V�>,�d��q�H�%�@�R�b%D� �@J'o��᱔��<����� D���cgc��d���J�lj�>D�P�� �2�X�+R�n pЁ=D�,#t&�$��3@�M�m��:D�"���*1ZX�zi� /,�Z�g<D����&Fʽ07��>�"��F�;D� �J���(9�`oM� � L���:D���d,�"G�d�	�>����$D����MJ#.�Hd��*f�*I�$�'D��H�`�5�z�XbN�0)K�pj&D������-�$��l�����D:D���g�\'�t�8t���<�t�;D��J�j�
,�r���z7��j 9D���i6T�Q#H�U~z�a�	-D�Ȳ`�DZ��YQED�t|z�C>D��!�G�^�	&��s͔<�'m8D�P���������C�zT�1 +D��j��]��]�b U	7L��q�<D��·g��p5�8���!�DXQF�:D�@��_�	������ $�8Ԁ�%D��+b,+	GU�錍<��e��e$D�����HX����ǶN̖It�%D��bv�/D��I�i;n��9hơ#D�����V,zx���Vǁ�/T�%��!D��`��N�t�	��F��V\H�� ++D�� �yKP@�7Tal�8�o��k����3"Of��7��/�@dS�LD2|�T�("O�Y#��@Z�E�#b(d*�"O���W�CJ��J#�E[���"O���VE_#F<) +�� �["O��K���4f`9 1�C���I�#"O*1��/B�
����j\�L��'�|�b���.�x�J��\4Ut81{�'����
�A��=�!�*K+�}r�'ҵaѪպM���!i�w�B%��'�Aܢ<����@�7aԴ��
�'U�Q��n:�ȇAU�G�x1
�'g�h	1�¾1
|:d��E�($�	�'CN�2�.M��ïA�Йq	�'p��3��Fh5�b�Ԃ?첈3	�'�.���
�37V
%RC�2<Bl���'Oވ�Ebr$����LM�1D1��'�H����N]���Ѓ	�-���q�'�:�A��1�5�/&�*$��']�x�!-�R_���ↂ�-�N��
�'����H�E�� �`�y�ĸ	�'dU�w�2J���腡���`��	�'��h���ˠ�!5i�$�\9	�'��$�A)V�:d>tH���3�\P�'`�h"�Ŗ!ho�G�D�e"O�p@��,?�ZL�#N��?�� �"Oހ�%�ATp�# 
FXp7"O��A`E��F��@��'��HU��"O�l�4��:-�~���&J�Z4��1"O��2si���UB�8�dR"Or`�#U�;{�p��G��"��r"OL�f�C�mŨq�䖼h�hS"O��PE͑8�	;�,͛7�R���"O������a�.A��6 ۖ�y�"OF��0�̏V�.�paa �"�5"O���"��.}�T[� ܛ~��C�"O�����')�$�h��m���yT"O�����'��v��-�~���"O�rYu�Sv�F���9i"O�LȳB�5�R��2�O ǚ�[�"OP}�C�;]>D�b��I-��ዣ"O"�b"��vj����W͂ B"O(�����&�����B-�`�"O��@�(�r��CC�F>�E"O���5�խ G\ʃ�G!V��yQF"O�p�a��=��hF�,t
b"O�\�G��tk8�X��F�m�<��"Oؽb�O��n�X$kF�ܣm�U#�"O��X�׵d���G%ʸ&���R"O:����#^�@jq���:c��ad"O�RPA�8O�>��C86���c"O,��������c�#ġy*��"O����#�7�|�q��W!G���!s"O�U;��Ǆ,���f!S�	�d\�@"O�J��,�n�*�`��dtk"Ovܙ��b�qʰO�oSP�aC"OLH�b��Ď�8�]��"O �2��=�6���&��]#P��"O�\ō���1[S((D����"O�tcR@\",��S!�χ?H%��"O�j�Rhr���A֏�A�"OXd����w�^���i��F@�""OZY��kJ�RPq���:T�'"ORt
 �F�x�x��'T�[?� q�"O� <���o��1Jf$�Մ��{Ԡ��"Or�J�Ϡ6��`G�A|xN�� "OZ��� l�m�e��?Sd�QC"O���(?UpH���83J�R�"O蔡!���<)b�JY�2�U�Q"O����P��)q��'��Ӡ"O@f��S]^�wBJ�$��"Oΐy�ŏ�yX��o��`g0�ɂ"O�Y���$=�]���Ö/G�ȈU"O6@ W�I ;���� ��l��"O�+s���v��f��
$\�0"O�3˂ .@~0@��TW�T�@"O|��`�ƾvR8�����j��M�"Ony��ѾaG��R%B�*)�y�"O��`+��Uz$�
��l��`"O���oƭ&�vEuj7���	�"OP�� ��n&�ʃ)`�,�y�)D�4U��aI�J#�YO�h�E&D��Y���r (<�H/b<��Y'�%D�re#�	&,�A �&v�P�vn1D�da��63<I f�џODQ��3D��)p�V�w`�q�5�\'7_�c�-2D�\�g�"_�$�����6l�`8�&D� K��ȑ�X � FG�pB��:� D�L���ùq��ق-F�5�h��Q�(D��J2�Y��D�� �čc\h�i%D��Yw$�&Fɂ������c$�P�B?D�`#���M��y1b]�<���-<D��;t�W�_v�̪�J�#�"�G�8D����	˞`r�t �X� !b8D��#�HC�*�a�K�%�Ш�6D� ���H�!`"�⃯�C&��i%�2D�t�\-Xut���!��Ev��i�+D��i��F�P&,Z%�ϝ:(l-���'D���!���A2�-U�j�#b$D��x�HF�?�q8�.�8bch-�H/D�h��KŢX�ꁀ�e��?$r��'D�ܰ���4"�����o���;#k D�����)�v`��\.
�!3�>D�X⤤�/,!����7z�[�$>D��B�e��Uy'�	05D�yd-'D������>!1,0���_<���bm#D�H`gI�X@���V? ��Ao"D�T�1��u䞵��
*k�F���$D���fԡr�"T �9$�6�2��!D��	p+U;I����I*.�)�o?D��b��L�́�enܾV ���1D�0��\1��L�� U�^�yφc�<Qd!��TY�{�Y�elX�Y7�b�<q��DØd+�
�>�2-9��HG�<і���[�q!��G} &�8�ϓJ�<��)3~eåE;kU>��.G�<����%s�N�r����o�F��c��B�<� -s�`C�"G�h8��I���D�<���}���A��(!v0�&�h�<y��E*8 �a�Ŋ%:�d�)�#~�<9�d�V1����CƤb?��р�I@�<�s��}k2Y��E�q+�YYw�{�<A�.�2��M�A��
X�p�GkRl�<����d0��0-ˈG]&��e�d�<Q�ǔ00A8��@-�=d,��T^�<ia�]�g��22��*g0�j%��u�<���,�R�kF(B�jdH���Jo�<A���	���0�E�#Z.�s$Rk�<� *ȳ0	�(-�y�@��e�R��"Ofa�ҡ�����+�]8���"OH���M������/�zK�"OFum�h��qF�V��N�Z "O����A�q��B�J��3�"O�s$��9a���a/�<��Sb"Oh�e#�2n ��2t
���"OE���5a��}����4+�.���"Ol���I\
b���8�j�./�>�#�"O|8��g�H�Xe���
�@"O�L#��-$����F�0��"O`4q��֒sF�mC��[�H�ԭ��"OJ����Ů ifʎdG�D	�"O�u��`���"��2y!��)W"Ol)(E���39Ia�%�!:�@�"ON�2�!��=�I�0�
!���"O$]�k�dF�g/(�.�:�"O�]��+�?����dA�5*��*�"O��C0Nٕc�$q�C�t(���3"O�[$[7Db4�:p�O#�h�"Od5c�g�n����A`V��"O��P�� DL��F,Ԛ����E"O@��tL	h1��bfA�'Ϊa�e"O��K�B3���B�12�"Op��f�՗��AE!F�H�\]�@"OS /ьbҒ�ytO�o���"O����	LKl@�2�˂p�@�V"O�h��nʼ�4�߱k��Bd"O$,QuÊ�:��(b�޿glN�s�"O�����5��1�ʀ4����"On�C�� �j��u�O�^>���6"O8r�6l������ɩ6���(�"OH�kܧ�$���E�w0L��"OK�E�0p�E��\�Ac"O�1`����5]�k����C�����"OŁ�S�Y
������O�$4@�"O�5��M�
-5 ������-�^Y�"O"p��ҳ|�de#�.R�2��� "O�����X7^����2$V�)J���"O���G�lT ��$``jc"Oj%9�NÏr�����+���"Ox�x��V7�����gB�:��9�6"O��z!�h\D��E�j��,k�"O� Z�g��D������̊u{(xh�"OL���~MZ��A\w5s�"O�a;���u>�J��՘]�3"O(%pc�X?8�
a�&  &� 4;�"Oj��fh@�s�Dqb�	�A���B�"O��R`� [�� 'ψ\�� Z�"O ����Vh���5��RA�Q�D"Oj�G�(r�B�*�dS�J�z���"O���AO�f��b7���a%^UYs"OfE��	�!Y` t�W-�<:9��Q"O����N��I�[87#���C"O� 0%%˵q�<�:���	?*�h"O�=����@C��1�EQ�!�T"OFx����:&�D��'˃
�쑂"O��A�j�9A�\P�հx�`���"OnqKe�ݐc��Р��9�f@�F"O�0)�ʑ+t>L�1��;�|Q1�"O^ [�Iȅ�D3B�αqt�`V"O� �E�<���$-�0mjH`(�"O�����ǥo��ȸS��&��a8�"O��B�DR����	S����5"O� e��MX�J�LTQ��T����"O Q�d- 2�FD�e�D��ش�"OqrQD�	Y$])2I0!�:�Ã"OL����]�L֚�ҥ�M� ���"O�\; _�=�T�Ԧ,��'"O��8
_��Ud�)N FB�"O!�F��_�s�b��E	@�5"Oz���&N>�
���	��"O������(�-S2��*�j��f"O�D�d�K+K���P�ܩ�2Q��"O���JF�%o^=$�q�5�T��y��	�2:��	u�.���#5#à�yb��%K=���ԋW�7% c4���y"Ǔ�~��4�0���/7���i���ybF�!X�d��T��S~�Pc2���ybM_�SN���f��?<&u��&���yO�z�hP��%�+h��E���
��yr��o��zPAT�U�4�pO��y2�C*��*�@֊=њ�w.���y�*T�CPX�T��4�Y�I^��y򡓔zy�Lq��ׇ,J�;'�ߖ�y�
�#>C6�r���*�����
�y�˂	[,� (�#���t#�Y=�ybm��/X5i�$X�5�,m���ߧ�yrIWbɡ�IZ舁(Q��y�&�r����.Nx��%��yB�n��I��n�YUa���y��B�2�F۝�V�ڥi�(�y2(V?lfd(	@D��~i���㜔�yr��q�,:�!�q���`5&�,�yBi0<*��Ga%!���s&��y���d F,��$L�&����)�y�DS<�j-�WmN(}��E02E�"�y�� +q���7eW�E��ы!i�)�yd��
T*��
E�Ha�̀�y�{Kh`i��[ Sx:Td�<�y���	r.e��o��I�7�S6j�!�$L8!�l:@/޸;|�U�F���B1!�$� >��*ԬcqFm[2�ǟ;!�$S�4����v�\ ## B�R�!��ɶ���3��+d:��d��$�!�ǄG6���M�a��0A���!�Dşc�4� K�=1~��sD���!�dΧCp��Q���qL@z�`
.J!���-S]6�ڗc��; �X��Z�G>!���{J��c@��	&$mr�F�J+!�C�~a\����3  �S��!�D�4\H|(�M݇s�B�@r3u !��R�s�xJ7	=,Q�Sb��n�!��D,�qx�	�V@|)ag'C� ~!�S��d��W�E_VT%[���>v!�dH���xS@�׀s84�[��_�!�D� <l��hʞ=�	p�!�B�!�@��"K޶|Y�����!�D�
K۲@c�F��C��{�'V�3�!��1j�������4y�aD���!�DN�J����L�%E��!b�"Z�s�!�^>�d����$�R��Q���!��E�/�(�(>r=�A���H�!��	�y������'5�(� jP9�!�dT�u�
hjq��� ��J�!�ɸDO2!㇫
F�9�O�B�!�@��Hs�	EGR�K7��X!򤀤 P��hA�]묜��KC!�� �� �ک(,�ܪM��x���#"Op=�m�H�Ų���V��Ѓ"O<).�"L9`d
ݚ(��UP�"O�U���<|�
)��#�@�dY��"O����	@r2����M�|�g"O\m&<wz,��kF�r"O|h�%Җy��� h�| T�"O�D�Յؙ}i�H`(�4A�H"O>@0C� ��d+2턶=�	:�"Oj�b�H t�p��^�*v�j�"OL@�aDO�:��|cf��n>��iR"Oܵ"��<L�^@0s�пIL�D�"O.ȡ��L��8��B;oA�횲"O>��*����Z���=Àa"Oرa�Dm2$Q2��f��lc�"O��H)~� ��sI�
�RP�"O̬)�NY�@>�-�ȓ�d܌qʢ"Op�;��QF��B���~��"O�1c����s@p�G�]�8�Ɛ	�"O���r_��Q�-�;
�mcS"Ol��$@�  N��9Q-Ӱ	V�mف"O�pw��k�vx;�N+6�d��"O:��pR�`Q�e,�N��P"O~�c�&D&}M��!��5i�� �"O����Bf�ƐX,I�wr�,"�"Oy�։�7r�+�%oU��r�@Ku�<@���9C�=�t�ۦ�l�g�<���; j>���l@�Sy��*�.�y�<��H�!� S:e3�H�"�J�<� �P�Z�b�z1̃+';��kG��D�<`/~���d�ɱ�x�)��L@�<a�� �9Q��(��"A�ȓ'����X�!Ȝh��K�-@��͆ȓ.��$��B�6�J�ZE��.%�<Ԅ�mœeB*(�!�r��T�.��`�ά�f,��t
� ��G�]��ȓ*q�|�&k�Zʾ8��k��7,Єȓt>�r`l�h�ꠂC�ڨ�d�������RGP�b�0��GLO,��܅ȓ)���� n�w��pr��%"d
D�ȓtR,㵩K*,x��b��1m�`��:�݋�f׾|�������eĂم�.j0�x�&�/	��`��<z�ڬ�ȓ��US��'�j� ��y��E��A��|�2�:{|���(�3~��Q�ȓ��r^,S�n�Jᅔ�,��H�ȓ6m8����=�J92W/�: ��U�,��aZ5�@|�%��$����ȓր������7�r��#Y�\*%�ȓ^��Xۖ��2�v4�gB!~�A��Cc*�質A�_�Y� ������ȓY�F�K2��~�hrDC��J�\��u���靼S�ųw��_ݶ�ȓp�|��$U��1��D����ȓw����[-+���
bĸ1��cx|���_B�V�&oL,G��ȓ70��G�Vl:𣧮^K(���ȓS�BmCѣ
W�Ybe	m�v���Ff�=�5HԳ[*�T:Ĭ��N16���uaR`QD"ϚE���[!rE���:=�"��6H�AvZ�
,D�ȓ L&����?TŤ	iF��2��4��+n���ș�-8�X���Q!�$�/�F|z'���5��s&e�.O!�� Ru4�W�-2�q���T�sPzH�"O�y���ZHl�	T,�4>F��"O�h�A������0S�9G���"O��櫓�"kT!�rʝ���P"O�1 �LVC��#�"
���`�"O(43b�[T�`��@M=T8@� �"OB���@�a�ҵe��v.(���"OH�H��éc�)[焞4PMd}�e"O�4��Ě:{�\�� �(�r$�b"Of�zs��J�t	0EJ	
r�6�"O>i;�\�@����Vh�E�&Y+d"O� d�U����CV��]��)B"O&���7�&�/9ή9�%���y��D0���R�ό6Soh<sD@��y���6�P(Z�aT c�򡪣�1�y�nE�h 7�V]*#BͱQ��C䉝 S�)�B�4���qh�(q�bB�I�'b>�Z�7���wDH%]�C�ɡ��A�p!�.t���S���<k�C��t wF�6�>=y�(D�K�XC�I�-�������I,M%X�C�	�5� ������M�������%��C�)d���te��vfr���
�NB�I>�2���Zk>8��HM+C�C�I%ls�(`J-8W�Y5��
  C�I�F0C�Q�v�*&^��/D�� 
մI���R�J�p�ZȺ 9D��!FQ�B�v�J6�
�O���5D� �E55�ہIM�_3>�u�5D��ؕmơ��`ݛx�aD#?D��h�D�(2�D�iG��K��Q��=D�lgq�!�q�ʄ)D�U�Ӆ�~�<áG"� z"oX�-h��QW�}�<���9B]���:u �AE	Wq�<!��<-��[�m�A�q�Ҭ�C�<QNX;.��VlS�O�t�5��@�<�TjA�$��rr&�	��@����}�<�u�E�;.<�S.�<ETD�#u�O{�<9�c�/'Y��`œ1~�beG�s�<���]9�z3��l\B쉵k�k�<)V�bqI;r���*�0{���r�<I�(�+J؜�qeN[a�����c�<YL�
�x�N"��J7�]a�<��#_�<k(1�,��)���h�A�<I`�K�W�
��&i�?T��,a��UU�<��g@4�����	>4W�����G�<�e(z�.��t#X�=_J$�D�<���~x��%߫�^����y�<)ဇ/X�"��2L+GBx�Cu�<D��>� �Ώ���S"EY�<���ϨN�^|��" �ќ�[��}�<��8p�L��pKG�<�t,�E(�x�<��&Y	PL�e�
yE �(6H��<q��ۛ 
�Q�a�A��d�QnF�<��c�?�b���)��L16 �"m�L�<� ���`���*ΰe�p)��a�<�!O�)3lڱ"� �_
xU�G��`�<�D��3 �&��$(c���U��w�<�!��8j��Q� *
:_z��P��x�<y�DOD4d���8FQ��귣�K�<��� �Y#4LȌ@wh�X�D�<�R���{��3EJ�[��5�ǈ�@�<��)g�UA�
W8[������T�<��Ŧ	����	�������i�<� j��5�	�c+��K�KN�n�z��G"O�� v��<�1B5��*l�l�h�"O��B�f�;J��(;VF�f����"O�L�P!G�y`trs�Π����"O��F* �//�|[�TSo���B"O��)���q���᝕�0�!"OLPqGHT6u��o�~�h��"O��iT��M¦��-Y�J���9P"O1�'��������8*�4( 2"O��㜙	�(��-��h0��"O�`�2��P��MѦJ���"O�Ɉ$��X����MR|m@�S3"O ���-7(�ȱ�l�`v pc"O�)Z',���3"���y+,���"OT�2c�X&1@�2��6"F�KV"O�{�JW� oց�C�G
9���"Or�������XH�&I=0�t�X�"Ov�1�ԋY	*�+�nU*�(��B"O��'�K�X�8)6�J��49""OT�7'=���7*�Fv�x0�"O���C�	-�@s�脪l2I�'"O&��aE]%��`	@�E�Ĝ��"O�%@áY�9��������Lq�B"O�# &��n[��ۢ�٧g�|}	�"O��	
�|�*Tjǅ�6 !��:"Ofd�pBιH͈�kU��9	���r"OhU�eK�)S�P�D"T�Ӂ"O>u��%,Zu���Ͳ'�8��"O&�d���)�����!�JC��b�"O�yb���G&��AϞ+,\�|"O�z#��02�H�S�,�i� �e"O"� �C�;�v`b�H��M/jY(�"O�4x��,� )4h�?P8�Ԛ$"O��Aqo�!]M��H^43F�"O^��c�y�D̫$l���D01"O�ի�X���h��.پ�1�"OH���ցw��2E��H��!�"O�}�-Ɛ�FQP.B�A�"OҀ�%�2=��B�Td�"Oj%����E�DI���H=D��m#"O�)�F"	P�`T+���E p"O��c��:)�AQ�,�\)D"O������r�A��5%�	�V"O��
��&��lA�&@U��"O����>#���X9xAR�"O�@��*�,����j�) *]�"Olx:��)
�kVd"�:LZ�"ON�@#�*�Є��̞N���Q"OT�6"�YP��С�I�u��I�c"O~��bI
%`|`p@���.$,� "O�|�t��,E�ZuA��ϣo���kb"Ob\����M�ZUu/�ⶐ�"O�IJ��C0o2"�@��� ����#"O@�ӑ/Vzt��c6��9UhB1�$"Ox�ӱ�!����vi��]_`"�"O8\{�e֚*�|0#P)�4mc`"OF�3�k\�[���%�Z�8��$"O0HÃA
4�!�ׇѻe>�[e"OE��jՋ	+f���& �hpq"O�]h�� `�0�z���@��@V"O�X�bf�DU�|��,ȁ�P"O��:�(��5,��9��s�`���"Oȥ9d
ư��	�M�B�"O��@��B]�3�"D�Vʲ�P�"O� �]P5獷!jj%��b�Z��4��"O\�cf�	4/�䌈��-L�$|"O�-A�l8�P��jS]�����"OBd�D$(Iµ3F��?n��uBs"O��Q�lL��J4b�.�'Rt�H��"O"���≐.,��XmL�h Mѵ"ONi�!�W���C $%��;�"O�ceI� $	����Y^}��"O��f	ͷ" �Y�Ϝ�	�P{�"O|�Fj)?
�A�H�-r�Z�A�"OR��3�Y)>�Z�)��*r�dmzw"O����ϕJ�<4I~�j6���yB'J>G�
<ʅ�Y?A���j�C��yB)փd��	Rs��l ��LC,�yᝍiv��@%��c^��%�׬�yb��H"pT�vJ��s_�*u�I5�y�j�! 6�|�$A\�g$�Z�����y�J�<���@X�I�Qz�ݽ�y��F�0��
%I7��p��I9�y�D���t�� �!_^�(p�^��yr��ffnE�Sj%Q���qb��y�)[N����"�4Wب:�ܭ�yb!ߴk�⌓եB�&a�0k�\��ygO$��̫Ů��!�H����yR�V #�ƕ�ʅ:!�nԐ0�ѻ�y�ԪlBls�-X�@)�P'�9�y��8#d68�c[
$�tC@nY�y�	�/!�|�*��˭�����)2�y�̤h�bI�0�ϐ#�4-b��Z��y2�E�bEX�d	ǋ?܄Ӄ���y"�m؈ݹ�A� ��1���U�y,]�m�<� �r��-��A��ybÒ"~���V�Za�2�+'J��y�e��\��e�O;�@pQ��R��y�&�>J�ٸ&+
iBx� ��y�]e* As��҃3-�ć�;�y�fݞI\-z �n�#2
��zRR��ȓմIQ�E�;�J���b�<X��"L��Fc�hH��,U�r:~���S=���-�3R����d'��h�ȓ;�VM����t�*y!��r���ȓ1Dȳ�ǎ7SVɣfe�� XЄȓCn��:0����K-p�>h�ȓ0t�H֠H>(���%Î�Q�0���P��]�Rf�?%�,��2,[#���3��k� ЄGS0�dg� �jɅ�+K�ېdC�e��\*�H=Xt�	��sOH�7!G�޲�)���5w�>�����X�@n ���յHђa��c����Fg������8�
���3����5l�%Qv<Z�b٘0�E�ȓ3:���t$��*Ĵ| �eR;`���ȓ[��j�B5{S8�d�ضJҀІ������ZB[�M��)�6W-���ȓ�psF�C��J�
&�U9A����ZU�PJCz��A� 3 �~B�ɕm� �a"6F�����c�C�I�dׁ�s�h��)�ex�C�ɠj�(� �	�rh�E� \���lLb�i!Lo�ܸ[�O�
nq��])��A� Q��m��AI1(�ȓVPmJw��4~u��a�Ԁfn�� ̴�eA˻VS���<,	U��7Zx
т %*���+J1�]��S�? �=�e��pa��Bn9Y��x	�"O�w��2�<xƯ�/$�F�Y�"Of=Ac�J�!���o�u��4ؗ"O�a�tL^2,"��� C���;C"OR�/W�y�Ȼ���(I�Dp1�"OBAء�^�<���; χ�F	����"O�\�6��J�Ƞ�쐠 �!`�"O��F�؄R�f�B�kN�Q��,S�"O�i���+=~+�*_!n� m�"O2����tg�=J�¦w���z�"O��RDĘ
�z�����k)^!� "O�|�پ��v�?����"O|93cMR8�x���ՓA�
h��"O��S (V;*ط�θR�Z9��"O�4 Q�V1rƨ�5�����@"O��� �I'g;�)aD\�{�4�´"ORm#B L�7��m�"�N�x(`�"O|�I��+|��hX�G�Whp(�"OP4���Z�XZx$	U'I�{{R�ZE"O���2+�"zY�,�@�Thb.Q�5"O�ȱ��& �j�e�G3n��P�"O� I�iD�+F@	�#/�'��S"O
�QdL�B��1G�\�P�"Ox��?�lH����'G�V�@C"O���'0����َY���.��+ҧ2�"���H��*���1.:���ȓ9ߴ���,��P@A�Z�ʔ�ȓ/��b�>��A�Vb��5�ɇ�[d6�i�D։Mʅ
a��o����ȓKdhƽ/��}��mJbʂц�t�Zm��[���K�aOT(���u��"Z<7@1[��dT��ȓRM���L� U�U��Y�@��ȓ �IrVmI!L�Bu�BcB�<Uh�ȓ��ᙤ�5N���r�GN����ȓ(�r ���ϑ�PкR�.R����k<n��&@Ɖ5x�����6v���ȓT�.}{��'$	�@v���y!�O���'t&ʕ;~q.��V�^�`!�D˾<#�D��ƚ	X��p�B�~INB�xVQB�Kv f���L�5i�nO��=�~2#�]�h������&Jl�v�S�<���'p��a0�D	��be���V�<a�E�,�������C�\u떉Nz�'N?��jw���%�RҸ�᧣;D����
=�!��A�'m~M0�$9D����
��E�@�N�|<�ɒ"o4D��b��Y�nIJ8a�ʋ�x;ru$h-D���p۵=Aԩ(VbJ)�L����'D������dYfA�"
6킹1QC*�	F���'����o�M�\�֧�&^ �ȓ ����	�4fY2��JΆr~ ��C��+dm��ꄙ��~��DzR�~�`��- 4�5ƒ�[��#��o�<�a��A�Ā+�gU&"Zs��k�<��H�=�4���S�1͎���L�f�<1���S��,zW�B5Up}�
_�IY?��{������+.�*��L$y`���ybZ�Bi�!���z��W��y��:�B���B�~]�!�G�Q�yB`�;��Uj��Ćx��IJ�	��yR��!b� ��WD
�C�0��%�?�?��',|�:`"r�^UJc�P<���'�0aY"*�y�vZ)[9Nڲ���� �p�@{t�D�!a/~�����"O�]�d)B<)����b%@<=�Z"O��Z�'�X6%�q��=ZjԐA�IC�'�� �1��4���`�g��o��A�`�L���5+t�QILT'I�]�.ǖ��c���I�:1���c,T�>`�q�,��J����)扦/7N�Ǆ�_�񲳃� VV�ꓐp?��%#�Jt��¦p� �#�b\�'??UCefùw�x�BF�Q�3��Qp�I5�x�!�63Ҡ��D&�*��\�揄�yB'���i@Y+|	I@��tB��	2�މc��S%r~�!6 A )0B�I�!(,�3A 
vX��]�m��C�I�?�T�4���^�|�Zb�kʬC�ɚa~E�Q�� ��٪«O�{�FB�	�a����vFY7$x�Q��C)8�>B䉂k��	Zq�AH4u!!��&�>B�	�#� 髠@W�B�����V):B�I�mw�$��(]� �4��9{P:���2�ɮ����"�KU��� dh���fC�ɚD�zdY�H.C��1Z���
ZC�I�>.�"AM�5z�ƅjြV(�C���<Mk��E�ԥ�©�;4.\C�I�^I��%K
�zL+u��	:jB�		5F�1��N�;n�0X��:B�	A�+p)Z�{R콘'+��B�ɪ{+D���-V1Q���(���<PB�	�a`��4 B�j�u�#']+��B��[�ك �ğ9�����Ϡ&mZB�I:(F�H�&��<a}��2�N��6�@B�	�J:� fΗ^{$m�ӄͿ+�NC�#I���pT���LR"����U�hC�	�E&�(�T�ݒJ�����W�>C�I'j��@�ï�r�)b�%RO�C��6?�6��ԂH@<ÁF*;��C�3�*(j������J������B�	�RM�S
�Kn���ө!pSdB��JT�'��Vh�I( `Q(HyzC�I�0&��)
.l�a�g� `�RC�	
9�U���Y��p���� H0C�	5_ݨ��āG�(Q8��H�+`C�I�?�@ I����ɩ�F�fW�C䉟4[����ɓ[̐��È|�C䉢Z��D2�(<@�H�G��#n�B��1�Q�R��6U��PC�@,X�C�	�F|сGX6|����Ǉ�&d��ȓ�Dxe���jL�x�D�?�z9�ȓMO����{�8`%fε*|$I�� D�j�0���c���&a��%�ȓ�&!���'���h��G">Dj���sƾ���N�(_��

>,���h�mʦ ��%2�U�\"�`�ȓ�>�"�MZp�6�\�F���A<)����l|�8A��	]�>Y�ȓ}��͛�b�2c��8S'�!Gډ�ȓl�&�R���z �A(M��7p: �ȓil\������,���BW̗�L-:5�ȓa��yq�_"9��i�YO�&0�ȓM"xڣ�D	 {��p��Cx&��ȓ7��TC��-.�����H�}q$���j(�{Tc��|�\rS�ԏ�0��ȓ�r�Ô'	|�������\��ȓE�x��P*Q�
�,�p#e�-=J��ȓ'.~�����=��=PA�?;:���S�? FĒ��2���@��'�R4�c"Ov���nI�oJ(�d.	#7l)B"O�����$p�=�'��m��"O��B��Zu��a��-q.��"O������R�3 F�5��5
a"Otͨ0$G;|��ԸFeΏL �C"Op�X3�-X��U���5R�F�*�"O���*ؒ�!Eb)+��4"OP!HqKҤ1&�JP"�,=#꼋$"O���4d��#m���߃f�f0"O�h �KˣŮ��E���F�*]�2"O����,3`�L�g[���h�"O��`DI�d�n-�G�?|�ȭb`"O:L{��,6���ɑ�<	|�mre"O�2���� pD���Z-Qm�x��"O����||DA�CJc�� B"Ov5�Q�Ӆ���$�!���'"OPA2"+
�0�B�"��U�1��Q��"O�ёc n��(�k̸$�8�[�"O�LxW̞;y#z�+3��;��1H0"O�Z�i�'7Y��B�C%}'XȻ"OzUW���0ݞ%�EJ�]2A{�"OP�7,��(p*�d�%H�0Q@"ONE��M���ۢ�y₰��"O���T�J�f~���0t��9�"O@li���6�T@��X6>p��R�"O�!J`�/0�1�t�q]x�#"Or�fJ�G�T˒��+SΝx�"O�
��MR�*���IP���v"O�eX�G�c𭫇j�c4>�S�'�6yK�C�7_+�"�Z��ViH�'X��ʞ
�Hy�k�<X�����'�	bV�Ӹ 
�����' �8�'3ҙ:�-	�������}���'���Qb��J��x��_�p���'+$x��[�}�tl�1�܇�
�`
�'63Q�]0M����N���D��'��գ�.�`�9У�����'��\��d"uÕ?��u��'�����N-;���${Ì���'2,p��@�44�N
����'����X���`F	܌�� ��'cʩ�㢀!@ny�r
[x�$���']X@R�<�����E't"����'Q=���$թք�H�模���`�<�0�Y�y� @I�l@ +$��0��E�<��ጣG.��K�OA��b�HN�9����<-�Iv���<�AE`	J�����
^HAь��<)$A_j�� �T� �K�]O�<�G0X`,*7	CF����$D��k�덉o��P���&2�+��(D����@���=aí���:Y1W�$D��)�1�^0 ��j�\=��N/D� :�m��/�,8�žOZQ��-D�`v��%R�B���.�}I�+D���cF6l��dc����f�T��#�&D�����:}\
傣��b�<:A3D�$0ɞ}�.y�6��>C�m
��4D� T�28�fЈ&c+�Y�F0D��hVAC�H�ݫ��
3|���i$D�����\�-;`�G5���6�0D��Pf�P0v�@X�E���D"D�����X�(P�Y�y�n���d%D��1�\�-�clZ�B��$!D�� ,u�0!��,0���3)�& ��"OЭ��M��T����i��^7:��"O�m�!)�b���� %�)9T"O�A�Q�S�r��!����"OV��	�\Ԝa�g/�h|��#0"O���w�E��zh�䖲c�h�#"OF`QRS.�QsBđf�ب��"O�͘��%:\ [�B�=2�̸3�"O����Tx�f����xI��"O�a��D�@�80F-6i�T!�"Othy�A�l2���#{xE�"O�h�
���c7o��q["O(�����c7Թk��Jy�M�3"O�t1�����,�欇I�| ��"OL��0�.���C���J�"O��Sa �)8�diFo� �d��"O\��Q,�,5%N�Y��U(3�M�c"O��9�B���� (4͜;�ʅ�a"OrI2+˼z��ԌB�%�&|�"O��� cؗNJD�bW���, ��"O2%���أ_��8���2�pؙ�"O���(O�/(*�Y��K�"�vH��"O	�'�P%{:|��Y 2��"O�X��`Õ's�e����G.�P�"O�� R,��5�h�7m��x�"O� {@�@7C��	J�Z	V����"OV5�l%lP��V�	"A:��"O�(��@�*�)[�+
�:R�9XV"O�tK��X�5Ț��7 ȓZ�=��"Ov@���ܶ`� tɣ���Y��(D"O�@��" �F��d�G�)<h��
�"O`�a��@=b2�����/���9"O6E07(؃�|�Ao��k���hE"O�ň0i��6ز!�MH�v����"Opi*���rJ�S�+��!��QR'"O����	+�@C$)3>}BHb"O6�:b`B1$��ԙ��ǬRi��"O�$*Q�
�v�|�P`��m�("O�mHЌ�r �0�d�D���ȓ%��}*�~�N0r୞��ڄ��I�~�L4z�x2)O�{B��*���vqF��^�y�D�3lhcăvІ�Th�����!5�PvBa�$�Gy�M0��i���#���y��0Xsڙ0c��#p���#�� �^�ݴg�S#0p��3@#�`��Gz�����c+��:��9R�M���<�CkH;��	)r��C���A�h�.DH࢓+�0Y~a��==�l�j�d �;��M��ɬ�,!˃W� $�$!��+a��' J�Qr� S�P���\%f}��:c`D�'�6�
X:�N݇i��"(N�x��4�!�W�<�b	�JE���P� �b�D�b)K�r,���d
�0b�&��,��!�"Ix�DL	Q&q�w�>��+ �\��z���3z\��'�8��1�֭j�"`� ǖ�e��a�r�fp٢�NB�ud�x&�޷(��H;fV,i�,xڈ���p������*O�m0�eѾn�џ(h���p8��6��F��Q2�%��]t4��.]�6)��gM��)`%��H��=�u���=�tfq��p@A�Y����ӆ�Ty�a e��:P�ϙ"Z.�qQ�/-F ́���A%�����8-j,Hkq �C�:$j�"O�X۔b^~��	��Aߖ�������ٵτ>b�`�Po�R��}�f�'��I�|^�"�B��KRHM�-�����VbJ�IG�	n؟<����ِe�&M���jE�%j���ġ�ͺ�ti�,�P���!��"!(A0�×H� e�?I�2p�X"�קO~8�F\�'Nrl��KE�4�$E���7�8W$S7|�I$(��u��ȋ���Y��X�c�A�R�s�K�|����?�Ddz�D�*�f�1/�>Y���$�B]�գ�z�Q�V(��q($b	�];h��'����Ex������hC!r$@�R�"O��BQ�ب#v����3u��
,Κ�"`��	v�	3�A�:bT��Zq̸?A�-Y;
��1��w�HIX�#�N�A��I�P��S؟xc"/��� bmx���2l�r�D_�w-p�4"V�qP�	�Af�"H��BW"I)pE g��f��ð�S�z��I�\�b��6�Ew��ꦃ�eC,�@vb՚L��uh$gV!F�\�ÉF�.0��@Q�Q�v5"d/4>�`x���'���*]Red@�V����O@�
c� 4"��z��N��\PՎ��1<<8�b�C�N�Sc>�$�B��
,�)�p#�"U"O.@AV"�5�(=K )q}�!F(Cb.V�b�3�Ґ�f�(HI.��c�\�bK�%λ�h|چ��13��;A��3p�q��	�O͸�-�/R)����
��f2�@r�J�M��Bu���p�BV@C�%Ӥ��tM�,U&�"=�pK�d�5��eA,A�-��w�'Y�4�p��*x1��{j�u���I�M���2��\1t1ԏ�0�����
.R����$�L�ģg-B2���I���N7�I�j0�)�掰�\�J�'qC�ջ�CVc����(�JO����w��P nժ�"O�%��g��L?��SR.R�
�\*�I��Zs�����
>%�$�HѠ���OKqO��C���_���ZfN�
��@���'���ka/��-Ix=�b�)�Ƅ����:�tu�2�V�-���.`F���82aڠ�0@��CјHxTFƙ �џ�y�JL)e#��b�S&����Q�F<z](ə���_4$�%"OT\Y���B�d�C	P�r��Ԝ�x��'ȓ#�����iً)\�G�DȚ�?Wf��a�
�%]R���>�y(w�f�9�aU�&��s��
�x$X���B"jްv+�th���yҊ�3
�В�ٻH�ho��Px�ə	.��u#��֐���L�0�Da��`Ҩ_3���A-z�ԙƮ�߼ �X<(Z�Z�(9<O����)^�R�O����!�1�!�b�ӛ�F��"O�9p�G�yj���ԩ�D�x�@B�$�A�|$)
�'#�X�₃�)�
�2�"|v*��c� 3�7x̑z /�1��9�ȓ{	�IX�C�1@*��vhğK2����|���B�SL�E��IO�q��p��e\�]Q��ƺ}�f��� ��$v��ȓ	ѰyY�L��b�X�"��L�����c�x(�$O4N�2� �E�1����
���{D�7,dUC��@�7��݄�n*��C��N�D��c�5I�����38�Л�K�.Dn�!%�	>!5��X��R�\�L��ȱ#%�D20��ȓr��h
T^5/�偕 0}t��ȓ��ͫ�]7-���	�͕(=pp���$���:6qCƟ~}.���8b���G�9�@	9pf��N2r\��A��JZ��8|�`g;.�ȇ�g��"��ϫtdP#Q͝�%�ja��e���cɡ82���2 �-{����X*�x�̯i�n��7��0[ ��?$��A�A�<�Z䟲_�La�ȓ%}<���C�	C�ʌ��/-��)��N��⃈Ј")�5���[*��e��O����r��WF�X)T��e�֭�ȓT/4q�S�����e
͝Oݲ��ȓ/�Z��/�B�a !��nst݇����H�&�r A���z��9�ȓ$�=���Q'I�P9R��='�bلȓY�l2bJ(r�LU�(����)�� t޴ˇ���#ʔ���L�쥆�,, x;��A�e5�pK#�=�La�ȓ�fd��_L�^���B����ȓs�"%��PGޠ�wB�.ͅȓUb�K���DO�tr���
(Җ��ȓz��ե��8N(2d��d��Շ�="��JK~��YdA·SS�)��WƦ����t���(��� -�ȓni@cDE���Etޅ�ȓ�(��E)�!f���Y ��7T_X��ȓP�LB���@��b��Y��Xq��S�? ���$#�pi@Oߵ��G"O< 1��� S�	JR.ؓF����"O� ���"٣�͋�q�h|"�"Ob�i�i�`��͒��.F�ze1�"O��;Qj��I��!���R�n�E"ObQ�1lY�Ye����9V a�"O�t�!�9/�漣S-\��\�Q"O��c�*�7n"�J�G��ԉ�F"O�(:�֣���H����5��H�"O` Y�d�P�l��m�1�X�x"O��Hs��(Q.��eke��"�� N�<)]�P�&H8��q��J���ȓK?Z�"ȂiklM�W�(B��ȓ*x�`�ƛ5r$�k�-͒ ߴe�ȓ1��P�$��X�AS�ᏓN�\�ȓ�j!6Ӟ j��Y1����l��Gk�,)��5��2w��ȓCM(\Xpf�/Х�B&G/njԆ�ya6䱡�B�}D�d�()𮠆ȓ:��Z�Ꞣ�0���o�3J��a�ȓl��p �Q/�3H���P�ȓyv|�ء!����@2�؅{v�4��a>V��!U�a~@j�)�=.���|���3g��H��	�G�.Ʌȓl��XD�4g��R�ȃ6 �X�ȓ	5�)x�ʒ{U�}Zu捸ub�}��4Q����	(޾UkCd�����U��!y�LP8l�"O�.0|����.ld0t�T.�����X*e���Bْ���&�6c^����(k�ԅ�!�H��սFB�a�B�&{Q$��ȓD�4�a 
� �v�R�D�C�IV��T�D�]yؐh�֬H0EcC�	�xe�o��y��Ƚpt0B�	�.��a���U4o�4h8�Bƚ�B�I� J� ��_�e��!1؎C�I"h�t�ȳᒄ/���⭍r�C�PC\tzFUr�A��,E/�C�	�XxD���`$|��8���7R�C�	 2�Ȧf�U[��a�OP�^C�I-�.=����G��u��L&�B��Yta�'+*(����$$K7��B�	G��92JL�z��صDK�P��B��)7���c�!�鱤
�s5�B�ɼY�pɛ �,>r����� q9�B�@�Sg��8^�.���*AxB�MK@�3��Mee�e#�
	�6	
B�!z�ͳ�n��6�|��/�+�C�I-Dۊ՘Bw<r(KG��&(�C�	�V�ۓ��F0)���k>B䉢T�"e��NG�u���-J�u.B�Io�L8h}|�8�	H'o��C�ɫϒ�s�m�0c�H�Q��I	L1�C�	"z�F�k҃,4\ଡ�E5�C�	�!O�(U��@�!��
��Aa(B�	�P"hY�ב>h���T��C�	�uΎ�b�� T=s��5+��C�I*��Ur�˝OO�CuJ���C䉻��2�˴��u�Q,�_�C�I3{���q�۵	�	�(�M�C䉰)�&�"v�N0���ivvC�	>GB�� ���*���&��,C��28��3��k��i�6�1�C�I.c�xj�MLf�*\�V�U�6�B�)� Fi��,�7��8S��!E�6��"ON���o\6־� vO֊Q��\��"OP���_�P�Ƚ����C�u0A"O@��'[ w��A����j�c"OZY@֧\�/l �1� �g�!�"O0��gbې?:J�H�J�"��� "O��)��3Fl9 BB;m ��"O@8z��@\�����Ț�d	S"O-㍳m�lD���2����"O0�a�l
�:z8�����#J
��""O���3��X�@�'�E�VP�p"O�
Q������-ˈU	R"O���c��q�-	p%�kf�Jb"Oڽ��g�3荑$܉p�s"O@�#E]m���]�?DF�b�"O譛�Cz��ё! �z=��3�"O��
#��>b��/\9mN���"O�	�邰q5�8xP���u"8��"O�u[!
�K4�mp� {:�<"�"O��ciN����!-d/�9�B"Ox����P�Ro`�B���� ;Xh*�"OD�〬Ph@�3��]�u.&݉�"Oh0��E�33w��h�1X,X@;�"O�\Q�̋q�Qr&�.�8J�"O4�@`	�6\�ل�;+隙:r"O ix��PK��%��R���F"O���M�/��Q`�����1@"OA�$�J ����T�a���`"O Y��(H n:t�� ������"O�@R���M���)T)ML �"O���>>�f�#��]V*fi�S"O޸Q��M+yJ\q���<N
�2�"OƉ��h�H{
����"wr���"Oܥ�&�� ^q9�i�G��4"O4-�6JI e:%�1�� "O��#�D�5Q:���)�#&&^}"f"Oн�K@}UjE%��pl�"O��b	�\���J
�R�"OTaC���y����iF7f���C"O,��gFS�%�d,����2�`��"O�q@�*��C�H�r�T�"Op�R�JP��GD�M�F"O\x[b#]7!�5��P�H�D�:�"O0��"+�!���@��ˢ,�li��"OX�0�f �0Jt��KӓlJ��R"OH�0��;�8a)��PU��"Oҁ���߭LX̜Bh�]�<PQ�"O�lS%b`�j����]�@��t"O�#e&����	"$Ғn�ƴA�"Op���NKư��
c�:@�"O]@���b%�Ĺ�#F~B�5a"O!`���PX܀��֡T�(U�"OX��D�	�J�zUj �[F"O2)ٖH)8�p��$�KBj��g"O�����%>���$��TX���t"O<ѳ�@��~�Xg�Ѕ%��$��"O\|�d��=�8���<��$j#"O��*�A��a�)+�$�A�+P�y��PE��� ��"���)s�C��y� 
xi<A����S̶D�%A#�yMM�'��5��8�� P�H\"�y�ε�d���4��#��y��^�CVi�L�q8`v���yB�^��8dK�&h���ڟ�y
� ���%ͷr+agM^�E|���c"O���4gU,YD.DQE��3b��"�"O�ݹ��z�i*
�>A8@�"Or���7��d���C�1OflR�"O~m���̹'->l�i�"O�����ϕLK�hxŁ�|/rh��"OΈZf�[�=�zDY�j�4C��"O��ΐv)P�P��6M��<
q"OR��� �X�˅+��E	"O����lҋm��� C���n�<�R�"O�a����+���4L�[��ۤ"O�=��-�,�x0"'�Z )�L��"O6dYSdGz�r쁣�L�"��1"O���ƌ5������y�JP*�"O�1�"V�lQ�pI_���x"Op��3]0}θ��7	�@aЈQD"O�#�N��8��M�/׭=c�e�"O��"���/� �Z�cO%^X�"O`!�2g
P��1fAY
w"@��Q"Of���k������X$:P�$"O`EP�Yz&@B�	m#�la�"O�l�F˓�HH0ErUA	�#� b"OHUy����*2��hq��>%��[�"OD-����
3�X*��E��i�"Oha�@�׋<�.���.Pd8��"O8a�5�!RN,:��G�F�-�W"O:8�mݧf0����aY��8�"OTd���Ou�" �M�=��"Oʤ�� ʐ;��� �C*"��Aۂ"O���T@ �B�O4����6"O0�
�L3j����3,�:5P���@"ON)0�Gl*@��i57K�8�"OR��6f�.�h���=R|�1!"ODB�f�	L ���șE� �e"O�}�3(X#}2�pM�V�:QY�"Ou��/��<]Xe�06�9�"O !ZG�
�B�>m)�ɓl���jg"O6M�u��1_�X+��"(�.%X�"O��	��+�1a�7�8zV"Ol���Ɯ	<Z�H��J�X�20"OH�&NL�'�:�z�l�.D�"O����K�N�Pq�!�D"O>@1g�_bD����R�*���R"O������V||{f�ܯ�.�[�"OZ��U��~�n �#OV)�* +�"O<���	M��Xⶏ��>Dj"O  ��*�� ����	V�l�+	�'/�����V˂4x�痄#� y��' �����l�a
�+�Y�	�'�:�Ş�E�Z��f��O��Q	�'#؀H�l�R���fO�p��M��'o�=p�=�����5h�a�
�'M>P���#N�\8c'Ui�R�
�'Sxa��DZ����B��k����	�'�4 	TL��4� ��VY�H��	�'ݎ�a��b(R�#��U�258�'Q�{�D�<�V�s#�M�'6� ��'2��G��� [�p�B�ܜ|�q��'��L�B��8t-^��%"cF �
�'��L��J*~kR�`�,, �1�'����w̓4"ߦ'��2�X��'��Q�g���i��'��<��<s
�'�P�	��x��̱u�4�P
�'ʮ���-�6môTH��۽7����	��� ��W˒x�v ��é����"O��SrG\����� G� ���"O���UeL�p� ��EN_�@��"O^��#��.I4��'+L�O�nU�"O6%��E[��X��
_�=���;"O��aP�ݵ4/��;&h"w�L��"Ol����ר8���ϭt�P]��"O��K�S=(Hej��S*]�
�IF"Ol�g �*�0�WI�b0T@��"OHm�G/|nl�;���MY���"O��R���<�|e���"V" \)�"On@YQ�m���L�=#pl�"OP3m�>i<�sw�I�]��5�q"O���7!^
�q�J��oF 5�b"Ony8��U3tXj�Y�+�A��|[1"O��I՘nq�]*&�΃ZR��"O81ee���m�v��
�Fɻ`"O���!�/p*(x�-X1bƜ�(�"O�0;T� T,�z�fT"UX���"O�	��ո4&<(c��	�읻�"O*Y�g�h
q�9���P�<Q��"@60��mY�6����ARZ�<��n�dh�������*k.��QT�<��b�26�"����#Ƅ�G�U�<7�*Ȑ5��,�D؂���P�<Q�@�a9�4q1/�N󄵢t!�P�<�r�H�st�TӀL=A�zћ.�v�<��L�~*�岆�Ҹt���I�O�<1P/�y\t(2q(��*<�{5�F�<��.�3xQ�$�K�r\n�#��A�<Ic� � ��2�#Ǯղũ����<)��
fpT�s� <&z�qK�"Mt�<ڲX{���e�̾d�,tC7Ev�<���!)�~H:v勡G�d8��y�<�B!�5��M×E���Y�i�y�<Q�.��s�����̀Z��	Ū�R�<i�߹'��P�ɇ�(�n��V�<��χ.I��McJ���%H@z�<�j��M:�-��.%.l���w�<��9T�(��'AT�@��c�
^D�<�El�,e����rBΰ�J�BUG�<ѥ�ڌZ팭Aa
�$h�BFZ�<مaшZΘ�����2���N[�<�pG��)3؄��	�{,2P{�ARo�<i�V&#�,ak�B�9������i�<�1hZ�֐�Sɐ
�R�B�a�<A�
� ;�j<�F�؀&V:58��K�<�jX.�l�I:B�pʄ.�j�<�@�0"v��r���$�:M3�ώC�<)F�p�Z�Aq/N�7A���R��z�<ɒ?��K��ކ�E$�t�<a5Ň�,@��x�b���<`㉉w�<�f�S��0P�C��L��qRțK�<��L��l�H� W9r7������\�<a���|����h:M�b��'��A̓J�|���,^A�08��O�-N�8��'	��hK�+�Q���0IA��*� ᡒ|R�څ*a��S�e2F��ԅ�y� IS��F���y�"M[���0|r�ٜ����gJN8?�z4���Juy�Kߩ9������|��	�pU�D�f
ҹ)����U7B�m�"����'1\qxC!��������TlU>���"l��$����_M�T���'����6�'�x�S<Fi��}�"��j�����H�h ̀�k��~*�=�v/H�1���I���M��;Q 
ً3���m	�|X��ʄ.�����=8��d�UڮH�����������I��<<DXc��9N�`�a��:�f]���O�˓u+��}ʞO<RӅ ͘D2�q�F������{��@K���g�? �-�T��oT>�0��8m"�[��>�q�9�S��^��)0�Ӈ<qT{&��>���	�<�<E�TIQ�	ꜽ�R`� d[�4Z�W�[��%�\���O�8����?a*�I	nS�m�f��&c�`S��v�>-��?-��Hz�D�l���&>���D�	R<� 8���?E�`�����?)�c�O���CDM��TP���F�,����(K�:bb����3$���$B	qj��l���$�!��CE/{�&܀R"O��WC�)t/���p����ȕ1"O�ȱ2�Q3 ���U
;-XQ"O�t��g@�IO6EqF�J�s P�A"O��b1�M�bj~0iD
�/L�a"O�e��	(3���c��1���1a�	F�OƢM���,4D��q�<p���P	�'(�pe"��4�4y0	S@n���'b��g�S�'>=s���:��=k�'r�l��ݶD_vѡ4a��)y �S�'-h,
�#� OO���Ĉ��&�F%��'
��8'K�<� @۴jֵ�ReH�'��]#G��#'�,�`�:��D[
�'z֡z��d*�]��Ѩ.+��(�'�(����<�ʝ�ժU,)�0$��'ȦqU#��N����)#���'��A����VФk�ԧH�:4�'
hx,��_����瞯K���k�'%����Ò�,8�[��υLeĪ�'�m�KK91�]�����=��'�:����3���n�x����'���c%�AN�HK2��\p�Y�'��]R&���2���[" �Hh(�'�<���=1b^�#&c�#c���	�')x}�oM�?�У���*N6:���'bV��wk�Ht�4��h>H���'�ⅈu�ÃBz���$��3��+�'��8I ���!Aq�ȣ-�N ��'�� �nØm���Q��Ǥ����
�'e�
A��$W�
\�R,C�[>͈
�'�h�gI�"&ƅB��ǥ����'����W��p�j|P�hg�ё�'מ}� ���h�̈�ʁ�jP����'��	`A��:�H;珁�5���'�����.�w��%��e��1Gzm{�'�U!�$�wߚ�a�+!\����'p�AE���4TD�_��!��'9n����K)�2���1w��(�'����ĤʅT�R���g^��5��'`�,�U ��PH�M�6��V %��'5��
a)��%b�Cz���'�JI�&)��(��ٷ|�.Y�'�6\QF�H=e�$i&�P�_�B53�'��%�BO�O�ʨ�Ԯ�1%'^)��'8��s@��R�x�J͇'J ��'@��93��k*��R�CJ�Mu(�y�'� d�H���3�C� t� ��'��-��-�;������$4��uI�'��\�5��#N��K$�
1F���	�'��LPO�-`!�D���� 	�'Q0=J&�ޯ;1�L����ސ�:�'A�d
[!:�0y�RxI�L��'����� �C��I��fSe|��Q�'��H"�Bٛ+_� qF�"]3����'Y�)bڮ+!vYǦ��O�N�;
�''L4[S�]���p�3*:L�<���'|��0��~���1Fh�&&Y��&��� �n�&dg�-�GD�5ID�p��S�? p O[!q<���-��l��\[�"O�)#c��$p�@��C��V�V�QS"OH�X�	�$���8i�bui�"OJ�಩�<:-L�k - +��{�"O�܋������0�W�8��D�3"OBЫR��%pHQb�J��|S5"O&����-4Bh�l��a�T�2"O��'�&B��Į/eٸ9�"OH�@�V�(&��r��r��`��"OPMCd'Z#���yu���k���2�"O (
��)�`�a�R�|l��v"Od�t%˂.����[�y�8��"O�TK�Ń�\�l1�����: ���&"O�@`�/�0(��� ` �n�2Y��"O��Y���ek5rD�_�>,��"O@ՙ�&-zȾQ���U$|�f��"O�|sr&�O�ʠ:W��8Z%"Of䁢N�
& D#DF�f8	�"OtU!$0T� ��#�->Y!�"O�I����b�|����Q�D��`P�"O�@��eS�9����̐��"O������DH!j 2�0�%"O����%�h.�v�����f"Oj�j�=%r,tX�M0s��lb�"Onl&�p�@��z��-�D"Bc�!�H=u��(�V3o��Ɂ���t�!�DܿZ  �T䓽_<�A�ˢ�!�_�n� 	OY\Jբdk�J�!�d�J����,Z���@�!�!򄔬q"����̌S@0(f*J �!�$9�b@aݸF��{�)�0hU!�d�0	��e Tk8s�.���/^!�Dʌ�RM Ϛ4�:��E!�dƚA�rl�� �"S❡A�G�=!�d�(&ą��Z~.���cbT�3!�I�Q�$N�)�ɧ`ܻ_(!�$��Pn�����X)�a�68!�D]=,RI��X-�~Qx�Q�!���ya Ey!���,{�( �i�!��J%]L�&�O�4�j[v���w�!�d�,+���EQt�$� �B(r�!�:#���JI��3�0 V �n�!�� O��m���W�5&�`cR Q�}�!���L5<�y�ɛ�O!>y#¯L�%1!�d���p��5��f�S
 !��Гp�T(��[��@��C!�dT�[��h�a�\.$�����	X�!���p��pˤѷ'����O"6�!�zɮ�Y"��&>�����d۶q!���i���Y&f̘ܨ|"�B\;!��1^X<8��|ӎ(�=x��;@����*̄R��¥Ln�DQ�ȓqY���0dL,8������=��X��2������N���e;Gi�2@>І�L���鳍��@� �퍯V����Bx�cըi2��gK�- f��ȓ� )�D%
�g�P�*��_�Eؕ��x��L�5滑�b퇸�$��ȓF��1ū�1@��̛��U3L���CM����^=4܋�P�JlnU�ȓ ������ۚh^$E(3Ŷt�68��^���в�ަwE�H�5)X���]X�0Pu���\�|�X�e4y�	�ȓ`۴� �`ˠ{: �CDѴ.��%��S�? l,����mHA����3_����"O.4�a�P<+~�уCG�0Y�h�"O~q0b�|p��3�G'=tb"O�P�ԅ�"��Q�el�2Xr�5�b"O����J&VP�%�&�V�P�"O )�بD�1R'�@.��C"O�4��.F���i�&: �$��"OB�7��%k�EQe��<5�PAu"O��9�n\�M���拵&��XD"O�a��=���"���0}y0"O8!K���YV E�%&�"|��"O6���(	�ld�`J���x��5"O��R��I����m� /���Z�"Oj�c��ڸ0�ٳCl����e"O�c��˴H0���D��'�ir"O�P&h�'/"�t+��U�L�@"O�5�d%��P����dCҘr�}�2"Ol���HF�M+F�s��в2�|�V"O�TA�ԕ�f�h�j�4)��,��"O�E2u�5 ���nۊ�*�"OV ����W�Bu����0%ͬH"Oh�1��оe����"2)��ʲ"O2����#u��%�(�l��""OPq)�/��zD�k��W�$x�"O$Y�`��3��2��\�p�x�"OZ8����8T�$+Da�/��Ѹt"O���\li��d k�j�["O�HK��B5�����ݲlkB�Y�"O�Xz$�ޱB�=+���06g�DI�"O�,J��	Q{b|��%eLJ��2"O�=a�U�V�P����Z kI`TQ�"O�!�t�M=h��48��'7��Pe"OF�h���&LdF�B�G+.H�W"O ���[/�����y���1"O�-[T�J�-ku`���-��2T"O��+q�I&t��Tk��O:(��� "O�ٲ�?k��L��i��p�0�b�"OH!�bǡy(��I�߶G�^���"O��avH�8d4˵FH-{cޤ�"O����M�Q�H��Rd��	V"O||0&,oc.���=[�
"O8���-F�X�ڕ� �Є@4" y�"O:�S��!J~�aw	�J��9j!"O�j&�
��Pq�ш��=7"OvyBՎ#V�6���
Yu�!K�"O@����ժ2<>��Ǚ:N3�"O���n�"���GF��?<�$ӷ"O�|z$	�3<֘]{�d�8n�`�"OL5ƀ�8�"�a� �N)�"OR|��+Z��ĄO��"""O�P8w��u�:������L��iU"O|��`ߙ�ıaǂ�/	��r�"O@�k�ى9��0 �%G�@	Q"OX�����UkdsV�Q�c8,8�"ObT�H'`\,�P�̾�	c"O����*-����]���0"Op��6$	��̃��  �`	"O��񰩜�2|:�)C��7Bօ�U"O��@�>$�}�����h�^��6"O6@"I-=�,��`�3Q��\:�"O
`�!�F8�d��	69��AG"O$���%kg���A�֑R-z5�1"O
%��o���X���!5p���"O�58W*Y�5�xȖHH�eH �v"O� �A�1a���H��bi�3�E�G"O�3��R�6i�3�&N�`�#@"O�y��>���ڏ"j�`�V"Oh���#ƺ]���c��U!p����"O�@4n��2�� �5k�+�"O��T��D"��Q��Ӕ"Om)%��.��'��0lnx�"O���,�!�.HR��Ę�`r"O��STo�6l<XSG�J��Q*�"O��� ��]���fT6U��y�"O�}��H��qz��˕�Q!U��"O
D�Ңd�����@�t&�bG"Oδ�V)tu���&���5D*��u"Oj��A������d4@�A�"OX�b�m�"K.�0p�@�2q��0A"O����	;rkFDhC f^"3"O�tӶa��"���Ф��f1.�x�"O��
P�0cx�x�B�l�I�"O8�R�Q-e= �
d�X�'�Y�&"O�4[��X|G�� �`��{�H��"Oؑ[    ��   �  �  �  +  �*  !7  �B  �N  �Z  ef  zr  �}  ��  D�  ��  	�  �  '�  u�  ��  (�  i�  ��  p�  ��  @�  ��  �  x�  �   T �  �  [' �. �8 �? �F 7O lV �] �c j n  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��V�XD{��	A+Τ�)SĖZQ��A a4H��Đ�3��Q�#�e��u�0���r�P����p?q��W�Z���)$���:�a�'CAx�@�')���%�,沸I�Nѧ%W �"�'[P�w�O�7���JŌŜ�.x
�'�~Ez�6M�&�e�Җ"E{�y"�'����s��\��T��p}2�'fNj�����?N�X�!@�	�y2c�o�}q�eL�Pd~	�ץ-���~"�|z�o�"[����h!a�xl�6Hg�<)��1By���u��#XyL\;���M�<q(��L5�WMݜ(��YC� LL�'i���H��b��X����St/�[�	��'_����(7�����aV�Y[�	1qO�ʓ��I|̧+�6�)R
�$�(I��oʺ��I�8�u�ӭi�*	�����Xa9}R�b�$��d�'#K������'C�h�遼z�ay�󄇀�M�b��"��t��׃
����@
k}b�)ҧ
�H��4Ǒ\�Rd3�ڟd��F|��]3Q}�#}b�H��!�msT�[<O��)3#�v�^8���UG,H�hǌO|��3��:�O��	�.�����D� �gI5�^B�ɳ Wr�a��@���!�0�[(EZ�OV6�6\O��/J�U����u#�:B�Р#A�'B�I5T\p]B��s�zU"f�7"�l�F{��9O~(I7!K�FZ>�0K� ~��;6"O����/!2����s	�X�"O\���9ki�`a旬>�|���"O&A�v-J��x�)�e.���&"O؉!�
��MsX���8a��d)�S�)ñwJX��W�=����U�ߋUa|�|�Cښ,~�İ�%/d�`ua����)��<!$��*�1K�,O�dh�����s�<��e݃���*r�Į3�9��g�g�<a!�.> 4pA��p���"i]�<��[�?X6���B���h)��[�<�d��@��w��I����E�n�<�e�78�P O��e��A�N�b�<���«v�b��R�^�[l`�g��]�<� 8��%�U�(hTyxTP=Us҄)!"O��"%+n>IA�Vo��w"O@)�R�El���*;eN���"O�d��D�8O����*���0"O`�cO��p���!��)%�L9�c"O�J��ʝr��"��7rZ�`��"O��Z�D'e���Z.W_c,� "O�E*e�Ѻ6'�I�F�R-GGhy�"O����_(��J܎.X� 1"O<H�W��3�`�#�h�_Or0k"O�m
��Iv�^�A�g�;LI��"O���*[<;c�=����kO�5r�"O)A���'vN���%�O^e��"O�0`�%�e��k��������D�<�@̃O��$��f��4�d`�-Rk�<����n�֔���&P�Ã�d�<a�)����<���8F�By���{�<��J�
�1WF͍n���ȱƔa�<�N·dU>p:GΔ(��%ÈF�<����-��A����|H!/B�<9A�����2s�E	�*ȣ�NR�<A@I�9F!Y�hܬ+<�+R��J�<���})��K���{�Š��H�<��рF{x���"e�)�*E�<�cŔ
pc���q��4��5�sk�C�<9"�J���p����b�G�B����Ԃ��>�t�s��Z5U��C�I�V�DZ�*��J	���蒱��C�	����4b�s��]�Vݚ;��C�Ik�NhC��\� -Xr)ݰgC�C�	�54�}b��^6 ��@2���db�B��51� m��e]��8��i�L�B�	�C���z�E7	1�ub�k�3Z�.B䉜=t�Y�#�:~ጕ;#�Q38C�<U$��  �U�R�җ�M�,$�B����Z���}�P��Vh���B�(���;sII�w���R��C�	��fa2�'�=K�E��e�&D�C�	3���!�"C�zu~y�����2˨C䉖^#,� 4
1K~�D����e�XB��(?�p#!�D=X5G��I" B�	-2'�@`�̌Zt&řwCF!y,�C�ɬ�M�@*(�!��ϋ�4B�Ɍ |�Q�.T=��b��9WB�	�W�jQ�4�ם	�p�W�un�C�	
D��<c���OМy��L�3A0 B��zt�9IP+ж��= ���'�B�	/DR<`�r#��mΔ�� ��r�C�ɘO�PE3D�0HQ|��!/����B�ɭX�J����J�M���� A�B䉨<��Qa.@�b՞��bO"�B�	�&�0���9�h�(P%L�DO�C�I�G�n�j�O
r��I5md�B�	�D2���H�#1� �0Ʉ^��C�	"{�8Z���/���rU����C�ɞ>�x���@6$�Q6�J |C䉪%;���-Փ"��q��E�nP�B䉄A��1a^����ݜC�C䉂i�Z���-ñ�p���#6�B�6�^5��̑, �0���ƾ;�C�*i���Ҕ�M,A��u �"R�C��B��u:B��1����MN:b>B�I�� sE^�t�j����̋Vi:B�I<B�����'�=9�J��[�TC�)� rȁ�Z���}����G�)�"Otd�3j�� 3���ү�=6%T��U"O�䊵���D�<4��o܏n��$z�"O�S�W�I)���cL�/kdI�*O�q�c"��n]���.��9��?Q���?��?���?���?���3�F,���ѻ/H��V̂#Ee����?9��?A��?���?����?�� D�ᱪ��g��mLի�oԩ�?i��?a���?���?����?!��?�u�!xM`89��>dL�����?y��?���?	��?i���?���?�s�
*H.�<��"�1[��7�7�?y���?���?)��?1��?����? 
W�7Sl��B�P�d��&"��?I��?1���?9��?����?���?QC�ҳ.p-�6,&������^��?��?���?����?	��?����?a(D�-��ʕ�N\N�Zb����?!��?���?!���?y��?	���?Q�Ǒ
$�x
�
��Iq�ţ�?���?y���?!���?q��?����?aa�P� �`�	���#��q�gѵ�?1��?����?!��?���?Q���?�aE۳g�4�0�H�6�šc��?�?���?���?i��?����?Y��?�Rm ;LYR%��qd�zABQ��?a���?a���?���?���?���?��BĜ�^�B0 s��IK�����?����?���?���?���,����'��I-y?��)u��(GP�	��8����?.O1��I�M�_+*��*TgԨ;���c����'�l6�'�i>牱�M��_�WmfQ:��ɤ*0���2z~���'2]���i��	�66�	Sd�I�'�~Q�*�%#s�y"�*O�i�|�<)���$,�'z���Lĩǜ�sH�.kC$�9Ʋi`�Ҙ'���8mz� ��ή���QE��%7���I����M��il�>�|�gʶ�M��'����.�:q�d��b1�좜'��-i��=l�� �i>���>`6��R.�*`��J���o�"�IHyR�|"m�4� ��đ!%�Сfɛ�T��$9ǋ<~��O��m���Ms�' �I�9�hQѧ�:!X�h3�ab�`Bl�*�/	/)Ĭ�|�o1�u'�Ob��w���@a	�)��%݂Cd�<	-O���s���u�&U�%	M�R�@�I��b���شz�$��'|7-5�i>���U'@mj��qHːS�ȕ���r�t	ܴ<�f�'��`��i^�	�S�u�2ĝ�Z�9v&W�@;�A�gmI�E�O0bڢ=�'�� �	�8��rר�J-̸{B��8vO���M���u���OAX�(�&3���`��X�	�/�>9C�i��6Mq��&>����P���EA6��gGT�|��)����G���`�>&�I�J�(gݡ[I���O����ͅ����#��,��ɰ$��O�����9��VߦA�an��'`��X!]Q"���QI:���Bp����4�����'+D7M�ͦ��	(|b����:���W! '&\"6)@��Γ:�>dz��l��0hw�?��SѺ� J�=�n�Ik$=b���H�ĩ�@b����cy�^�"~:��2CK(5&舥�2�j�A@̓���A�����㦑$����&��= ��P�?� ���g��<q�OB�mZ��MϧDa~��ٴ�~2M΂*���/>m�h$��n�	BG莿U�B�FQ��ɟ��4����?Y���0�����*��`<zͱ���<K>)B�i;�s�yrW>������� 	[W���V��H	'  ?�c^�Hߴ2v��0O�c?�F��?]n��72�塴�_�h�F(`5⏽3���|�c*��uw�;��� uQR0x�*Dt�=�G*	 ����O��D�O���<i��i7�H˗$�)��bIC�E��i�	zM"�'��6�=�I����ܦ�9��G7p��#���-�4�V+�M�6�i��iK�iq�I�q�P��.�!�'� �yQ�Hn���
�85�(a�'�	ʟ��I័���(����� Fe�D�+ ��!��Ի\7́(�����O��d%���O��nz�M�w�\3Gy�\��l�7D��9���MkD�i�O1�,�3�v����`>�e	�ƅPeՎ]����	� 9v��!�7R��q%�З']2�'����G��!P���O�=u�Xy��'\2�'�^��ߴ'(�l�.O���Y<��Pa���^O��U@�4kH��<�O
Im��M듓xbȃ�l5rQ���ӤU9�N	���6/��#�J�8Q�����#�u��O<����(e�X4��*LɎ�I��O���OR���O^�}���9��#[+|yVi�¢�zrB�O�lo���"e�	ԟ8C޴���y�'@�ғi_W��%s�����y2`Ӳ�o�(�M3� �M[�O�˴A�;Xc�`��ޱ;e,0q�N5o��M�w�� 1�\�O�˓�?���?����?q�m��\�sb<)-�9�d�F�u��-S/O�\l�[F���I�����T���X�G���ʔ@���)Y�11�V��'e 6͜�=;O<�|��W�v�Py*���3s\$�C�%}�1�_���
��P�i��dݵ!N>a-O̤� iNe� �pPL�f��BG�O.��O���O�)�<��iV�C�'=��i�n��Z�Zlf�ǥ+�u���'Y�7m:�	����LΦ�"�4ś֧V�@#���X�����q �(-��ⅹim�I�\d��;�+_	3�<�$?��=� ���$k�2�*����ܠ
���2:O���OT�D�OJ���O��?���f"&�2���X��9Y�h�(���X�4?�X�O�7m ���m��T��� u<�k���M�~D�	E}��|�8�nz>��,��'$(�tJA45��9���^��g��N ���*(ZE�'�	џ��ϟp�I�^vq�Nbl���5h)7 &U����ȕ'��6-F	U���O��ĵ|�t�B�qC�JB_� ��k~R+�>��iW�6�����&>����;���'-�g��5	�(�6� 9��
�&>g^HB�F@y��O9�d�B��j0%�`×! �Zb�s.�~�.�*�Ǖ��$��P�	��b>�'�7���4ٌ}��I�f�r48�BM����M�O�������?��P�PR�4J7Ѫ�*��+�.�r�m�"Ъѡ�iV\7��"s�$7-/?��*)c�	C�m�"��$��T�˗I�L]!�f� cY�$�<9���?����?1���?*�
ei�+�2S��s��Ib�%j���ئu[���ן �����`��'_7=�JDzt��-Ξ�YG�HgM�y�V���yݴ&gBP��S�?%���	ǌ\m��<A���!׺�h�Lk�� Q5o�<�p���ԀJ ��䓖���O��E�G�����@�v7|0�ן�����O��D�O�˓��J��	ڟLK��D�'��P�a@=mC�}[ ��t�1�I�M�4�i����>c�ƈk�fP��?j��l�# �]~�%�s��Q"0��3B.�O���S�����p�<@���2Ș58����,���l��Ɵ,�IB�O�@��Y��� oԉ@�X�`��fo�(��ƨ�O���Ѧ��?ͻ8G�hI�� !�p��M!��ϓ{��#uӰ5mڤ=�(%oZj~�	N�:a�u'�-L�ѢԮ|�n�b6(�(;AQ��|bX� ��͟��I�`��Ɵx'']�v�b�Ԉe쎭���@y��n��(à��O�$�Or���DY�ѾB6�E�x����&B
�8K�`�'lj7� ��A9���H�Hy@ ����IЀ�ٴC��SG	75O�ȋ���<�NSwƨ�@[w{��O��(�xT+6��2Vp0ЭW. `%���?��?9��|j/O2�oڕ0�H�I�Y�b0Rs.�r������	p>��I��MÉH�>)��i��7�P�*ծ3A�e"[��a�6(�&<�94�n���mD�p�p�Y!e��
N~�;1�ڤS2̒&�.�C���)��qΓ�?q���?����?A���O����w�?-y4�f�M�l�,M���'AB�'9�6�ͥS��	�O�lZM�I-k����9T����gƺ't��:������⦭���|�f�0�MK�O&�ؓ��bɴ��'B�^�y��Ǒ( �p����)J���Oz��?���?���� �b*���֤��+�3Hn*P:��?i)OFQmړW�
0�'�"Y>���ܭtc^@�J��M�L��4`-?iwY��Xܴ5˛VK�O,c?��w�ҟl�]'k$�(�`M]�%B�]p��=���+�V��Sz��@��%�'i͠Á9u�9�W��v��r��'PR�'����OE剖�M��]
P��@%�1�X};DO�P6`���?Q�i��O.�'�>6M�!�ƀ��/Ҷ�2Tۖmۦ@$QnZ��M3[�ԑn�J~rd\�r1��P�aZ�l��	�J�,ĳ0�2:~&ieD�*V��I}y"�'�b�'���'i"Y>�A��þ �.�E��j�BȘ���M[����?)��?����c���i������D�@�񪙙L2Hao��M�#�x����Kt�<O~��h�!Z�q"a��%� �Xt1O���#V��`*)�d�<A*O��K�k�m�,a�d_�2� ��'�L7�&p����O���������dé`М`�؏���䑩Oj�oڶ�M[S�xR��Y��A��
�)%���G(
����q��d�P�-W��kN~*�+S��u���O��!�I�e��h#�Řc�*,)�"Oh�f��;�@��$�"<bӦ�O�tm�=� �	ğ$Zش���y��Њq0�R����aQ����ya�
=m�$�M�r✿�M#�ObY��i[/a�� �s�M7d�y(vo�?8�H�a��>�J�O���?1���?I��?y�9��!��)hkX��D�Z���)O�Em6hy����Ο��Iu�Ο�1�`ځu����1+S�+���aU����d�Ϧ5��41����O��l���[NG�{�+�	3.���d �K�ux�P�����Y��4��7F�'��I�.琔B2o� c)�sY3�]�I���	ڟ\�i>	�'[�6m\H�b�$�!I�,���6jg�,A�!`����Ѧ1�?��T����4<TB�i���X�MZ�}�h;�R�p{]�r�2����|t�Ʉ${&t��di�����R��k�e��''9n�	�Nv���	ޟp��ן���ԟd��QoG�	�u���_�'[@mp�#�<�?���?��iVx���O��n���O��Y0&a`�1N v ΍���^�8�M;U���	_5,������3.N�t�J�Eg�&X�T X7���[�|	窋 Y$&M'� �'���'��'m�	�"��0H����-D7y'��E�'��\�P�4��mi��?�����)K�X""#.s��������	���ă�e��4�����D�&�
����_�up�A2w����
(E�Bk�|�5�<�'B{���Yw��O a2�
��Wr��f`B>O�J�rq��O����O����O1�pʓQ��&%�}�D���R�eg�T��ݎ]6��p��'�2o��㟸��O�oں_Iڴ�W)D�7�l�H��ۏ03Z���47��f�Z��ƒ�4��g�2ޜ�x���]y
� .c#7 e�K���9;����q:O˓�?����?Q���?Y����i�4n��n�@rt��H ��m�A����Ο$��]��|t��w��,�S��=��q�@������i��1lZ��?a�O1�� �Ex���(&M
B�Z�{4��u`3K���I� Ԙ�QD\�^i�&��'���'�X�A���,���`���$d�2�'��'��T�+�4HY����?��r�$�2pnH֦|ҳ��(Zz-x���>1F�iP��=�^,y��b�<J�p��g�ӕ#�ɫy�`�H��(#�a&?]�%MպsW�'(��8�\*J֡h��m0�'��'qb�'�>����:�S��!;RsrI_�3º���2�M�6���?��O=�v�4�l%�Vc�.Lz��)���AɄ�B!>O�pn��M��D	 �2�4�y�
2�0��B��M�&<�F[�&D\r��,9U�Ǿex�:$.ʓ�?����?a��?��Z�����^�1�3���uSi�)OAo<Y���	͟h�	n�S͟h� T~���Q�K
��昃ug�9������Apش��S�'"~�`�T�K�x���ȐL���ГY�`#XI-O0�r��u�ם��dWꦱ�'�>��$��9Yy �+�&0zH@G�'�B�'�����Y�\۴2=���%pX4�I-)?����$n x[��v���D}�aa��mПĪ�EGK

��þ\��L��ٽ��m��<���AX2t;q���4<�.Oe��ڿ;W�9_�t��m��T�R���<���?���?���?A����D#1^��m�z�x݊E`���B�'���p�H-�`0�
��ݦM&�x�C�;3tyѧ� ��P��BU򉢆M�w�il����S��2Oz���f���`EU� ��z����$4z�E�(X����<���i��I꟔�Iܟ�	�?ܔ!�L��k4�ي�$S�u(�p��ߟ�'6�7��k����Ot���|:ׄ�#d�r�"*�8��a�hIl~���>���ig�6m8�4�X�)�g?: �
�$;:��!���8���<��Yာ�<Գ�Z���y�!�(OF��R�ft�|��M΀��5ٴ�Y>)��D�O��D�O��ɼ<!u�i���rЭL������B�m�b�c������'�66-�O��ODX�'�7m:B�p9p��;B��|�"���-/��oZ����%"�ͦE͓�?����!�L	*�!����d��$���d���P@s(� 30Tm�eyb�'���'���'j�\>Y(qˏ$#7���߁{&�c�@��MSbd���?)��?�H~"��=a��w�)) ��b���[�[%�(���Fx�D�l�f�i>������e�����G��%H�mX�V�NX)�d�Kv� ��l�f\�3RiGdy��{�v��?��x���g���$��U豌Zk�䈣��?����?A/O��n�Y� ��I����I;ҵ�D��6^���~���?�_����4a���|��/��c2O˓��&�y��''ְ��DP"1X�<KuX��P[w� ����Ry��{a�y�+�P�Эc�Fܔ`|p��֟|�	��<�	I�Ob,�,Z������s[����@L�X�2M{��A'.�O�dɦY�?�;^ɬ]�Mѩ<:�����xlΓݛ��fӂ�DF�'��7�l����5W�H��a��g�.�zԦ� _�ط�kKlQ����yy"B�&��?���?!��?���=2T��ԃI X,@���w�2�a+OJ�mZl����'�B����'�L�y�.<�I�tB�� ���ӱc�>���i�|6M=�4���	�O6�a!%�,=섫Q��8f�ea�	�6Ilѫ���O*�c`&]b'zYXu�9�K�0#�[�d�1�K+!=�Ktr�6Pw����	��������Sy��{�v���b�OV���3�Jy
w?*� ��D�OR5m���'�P �O�o��Mk��'Z�D��/ʏz���J���lz�`����Mc�'l�L�f٠tIc����I��u��wӚ��*�^a��
�5K%�ڝ'���'��'���'���b��F�G��U����(�L� k�Oh���O��m�Ifl�S͟��޴��FNt�$BĹ��X�Q�V�6\"�SL>�E�i�6=�䁹��j���TN��XsT�,Kd�fLP�l_D��6��:-|���䌝�����'���'���'U�I���_c �@�c�"�R}�&�'OW����4Q���j���?����I�-	�A��eܷl�:LYT�̖>������Ԧ���4���|Z�'j�e@�)IOt�h@�#:�����o�;I�B��ͱ��W��7�N?�uw��<��;e{}X�A�9KH��o�%ش����?���?��Ş��$_Ц��`Bɉ(+�h w�
M��X&�
U����Ɵ|�ܴ��'"4�h ���
:H*8=Z�=o�`�h&�޿v��6��Oh�H�
r�|��� ��͋�'�L-����fy�ĕAY.�kuhݾ7�P��%�	sB6M�<����?����?����?*�xI�Mً!���%��ERDyB�ަs�����ʟ�&?���'�M�;^H���MK�e��ʷI2L��i��7-?�4���)�O@|��y�n执���H��[xVV<7�ݨ	��	d���҇dJ�r6��'�7m�<����?I�"]�Ƽ��DĒS��R��-�?���?����d
��m�|yr�'��x�@O�yӘ��oK4m<�S�$�w}��mӦho�~�ɕ{]Z�i˔���=�����	ϟD��.�Q8d���Cy���I���׺;e�'�xQ��O�)S�H(h��>�V��d�'�2�'���'��>��InB`u#ބ
�V�"2mC�oC8����M�Ca�+�?A�fћv�4����j����⫚�L�(b8O��lZ��M��"���:ٴ��䞉d�5��/ȺC� rm·J߬r"P9c��\�x)��<!��i��I����	�L�	ߟ��	�|�Q� ��#�6cu�	7>j͖'��6M+bK��$�O��$0�	�O�#�j�0M������]�)�ƕ�� �s}B�m�ܼny�i>������q"v�D8����$H*���+��R�S�/�EyJ:vD����=�'��7ͣ<�U%�)lI���.#���fb�l�ԩ�4r&.����[�ܬr���"2,P�㊭\x�<���OV�6�D�V}��f���m-�M�q�L����r��W�G
X�����$���4��d�aVU;h$����r��\�cL^c���^���xa��A]���O����O$�d�Ot�$*���'�
;6	3��X[��ɉ��O���O DmZ�9E�����ش��W�0aT�ͻ�$�Z4��D"c%�x��n�`mZ�?Q�B	�Ҧ��?aB>��@4I
�
6���c��Fl\cתG��`J>Q/O����OT���OR���ŝ.��� *ֱe�u�F��O��<�u�ip��1�'+��'��/�Rݲ�` ��"�����6C���$��&�M�'�'����i�>��3k&/etTytJ7_�. �����x�aɮ<ͧrd�0�Zw�v�O��hB�n���1@�0�*�O�Llڣc���Y��̰:�����Ԛj�8�:6
ݟ���Mc��>�'�imF�಄�B��v?K�����dӒxoڂH ZYlZY~����, �D*K��	1h>�)S%(R�p��	�a�҇8�	sy2�'/��'���'�rS>-�qġD�PU��EE�G: ��Q.�M{��թ�?i��?qH~z�i?��whRt��D -C%ȿ05,���d����A�)�ә!���o��<��ן?�r�;����B֋��<�R/�=��a:a�A��䓘��O<��#���#�&���d)Ɍ�>��O�d�O:ʓi
����g��'�2=[d�{d�.�Z��%mu�O��'$�7�˦I������\� M�� ۬@T�`f,ԏ7��O��Z���q߀�Bl�<��U\��2^wČ�$GD��LS!aU�<^z�ѩ�+� ���O$��OH��"�缣D�խn�.�F��?�ؠ�O���?I_�G.թ�?�������4���S�Q*T{�hY�h�@ȸ�7O��n���?�ڴe�~L��4���K#ll�H1 _��X ��F˵hP 3��#-wl��5-,�$�<��d���ۢ�0;�� {0�R���	)�MÂl���?���?���4fݑ�<Pp!M^4�g�$R���m���s���$�b>	r��rY�ؚ��X?<�0��0�e��8���D�X��)�'�ug�6�D�<!uLĪ`�4`�	��8p��M �?��?����?�'��A��5�7�����E�L�Fݲu�$"�DՃ�̟���4��'S0�hB�V�r�bdl��Zq�Ꞑqfi���.昄�p���̓�?��Ł�8�UӶC�=��D������(�3��\�r�f=2�(�6~���OD�d�OZ��O���5���0F扑�]9B*��$��`��8�	؟�����M���|�,����|�e�t�(x�]�!���<[ �$�>���i�6=�^"�fyӒ�?@��Ҋ�J��,0�&�*BZ�)���N�~���������D)�	�N�K��ƪ1R]{�i	�}K�#<��iT��'���'��"ެY� H�������o���4>�	��M��ihO�Ӵvhd�SA�%$LZL����>Yi����Ʉ��q���Vy�O�0X��I$��xp��E�r �NY(]K��2l�ğ��I����b>-�'j6m�&�ցiBjũKN���� �R~��A-�OT�����?��Z���ߴ����A��������D�a���i�46��L!`7-#?�AЧO��q�֮���򄗼=/��bV�9�i����t��<����?q��?Q��?�*�>%�Fσ�j=�pV�	&�~�A��̦�Xy"�'��OL"@m��4��<`�GY+"J-p��3^	l���MC��'
�)擥}!Txm�<��F�KU�d��+Y�r@����<�U� H��ՠA�
����d�O��D�j�pep���	>8�Y�@���d�O����O��H#�&!ع�2�'����_>!�V��Ǹ�6��>��O�E�'�7�Φ�����¥8S�	�MF�a�$͑�Wf���OZ���jS���f�<Y��	bԭ�^wj,�d
'@ ��Ä��69���+�Ib�����O���O��$/�缻��N)���Z�k��4�����^2�?i�i;|]���'q��r�R���"%>� �%<�����	tZ�	�M+��i>�6mL�u� 6�m�\��>,:����!K>[Ek�nN�H���KL�!��dc��Ny��'��'"�'�2c۶dZ����ȁ:�dр�@I�� �M1X7�?����?�I~���U.�$�����g˺1�A�.�,�0R�<��4ya�fC�OD�����4�����P#&�H#�Q�	p̲H�`�~�{�<�0��<�E�Yw�$�O�ʓ!.�a�ّN�Lxӏ��!@����?����?A��|)O�o�x(�ɺhdP�S��BEb8�������ɔ�M���N�>1&�i�6-�������Z���B�O�� ;�͇jmR�m�<!�j��Si��l�.O�����V���EHZ}��;���hK(���<O����O����Of��O��?�P#�Ћv<�fc�7kbx�	�ȟ���џ���4�ұΧ�?�׽i��'���Ѐ韣>i��U� �09F�*�$�����|:��Ms�O�QQ�� 6�i�_Bz�yc�&Zg!p8�����y��M��G4���<���?	���?��o��I�*��%dF�=�l�j�ϑ��?9�����C��ۇ�Y។��ܟ��O��8�4h�|��j1�N��4��O<8�'>�6��ݦ�L<�O2�h  ��0Y���v;�p#s�O$Ko��3�N�i>�#�A�Á�|�p x�F�=�J�z�f����'�r�'r���Y��S�4SԌ<��7>����/`�r�@��"�?)�3��'�'�6�)ӛfÂ/D���cق,$�����ג�i�6-T�| �6i����%'\�
V!��*v�'�hp�ٮ#�j��Ă$�E�'������I��D��������ā�4��xEN�q�ŢAN�!/�6�R�6�����O��#���O�\lz�	x����w8�q)ʆ�c 0�FŘ�M�b�i_NO1��X���f�j��38ݳ'�9
��h�����T�4{����  ĎU��&���'��'nP�d �v�F�Kc���b��B��'w��'BR��ٴ�����O:L/x�0Ȑ�;5$L�r��%O�"�O2�d�f}R�`ӌ�oچ��5Q�` B.G_Pi(v��'{,N��'���B��� G-T�;$��ԣO({+���ڟ�K�"ݽ.7��0DL��3�Ѕ��ǚ���Ɵ��I���G���'��<�'�W�X�A�o�m���b��'w
7�7z���$�O�mZ\�Ӽ��!h8(�>
#���L]r��8|����O�7ɢ>jZ6�.?)�B�C�D�w��!"Q��(��Q�^Ѯ����7L]��IH>�)O�d�O����O����Ox9c�V�\ E݁b��$�sF�<�Ѳi�lb��'�b�'�O��b����2UȜ:#��`�H�9�l�bᛆ�mӊ%�b>�cC��,c �LI�↽5'X�zFƙ��`���Fy��#nrpC��zI%�L�'�"�rU �E�i�ƛ/{��T�V�'s��'Q"����S��!�4aR�Q��2hf��	G$c�j��T��9y,j�j��Q��6�|b�'2�.��&#g�ȬmZ��0E�TVڌK�
2�6\��M�����'�L��h�$@�PĞ��"e��4�ܒu��X(Y�S�L��5t�(��ϟ��ğ0�Iݟ ��^8��KBS+ɻ����?���?��i��`*�O{r.y�r�OtqF���2"�Y�  &	����wGПX�'�7M���?wF8�l�|~�A����$X%ˍ>N�Ԥ��Kϋ]�����̍i��P�$�|�V�L�������ԟ )&B�`4ah"۫�0鐊������Wy��d�n��Q��O����O��'hh 0��i���/F�8݈T9OP��U}�ef� �m�
��S�t���c�r���)�,}� �ä@t�9�v��1C�kPS��S��6��|�'u(5� �T*XQH�N�j@�S�'�r�'�����O���M�턓:0�h󧐑���6�9٨(���?!T�i�ɧ���>��i�P��0��l�L�!K�q
�%x�t��)lZ�v�tHmD~RL�6��4CB�F�qR削Hծ�cvBI$vWz,��o�	N��|y��'`"�'���'��S>�I@��qu�,01��gE*��bD��M�7.��?����?�K~���=Z��w�<c�ʝWon)��/]�W��3!*`�@e�	m�)�ӫˬYoZ�<q�ŝ�].PS���M|���&U�<���5]Ԃ����������O��$^�G����`恏����Y�&���D�O,�d�O�˓H���	��?����?��"��mـ��l�M���( i���'�>�ɛv!�OpOT�Pbº-v��A�\A\i�9O��R Z�u�p�7i����2�ɓ�u�f�O:Es��[��]P�`�D4:�K�O~�d�O����O�}����J�
4O�� �j��<D!K�I��f׃~��'�86M3�i��憂C��P�f�>{����d��ܴ{�6�d���4"���	ٟx;�A����1����k?x�zw!��^��pR�CM�L'�h�'���'h��'*R�'��P��c�z|�����U!��S�[�x:ش~�*��?1����'�?)D,�^E��1���u��������M�v�'������O��➴�.�,M�
d�ԥ�J�@�9$F�7���,O`���^�֝�䓈��>���aX�t�"|#��\�0�H�����?����?���|�,Od�mڒo����ɐB���Ǡ�)7�����J�%\�	��M;���>a�i�,��p�N�Ѕ81�ԫ!�U`3���}U�7m/?i��Xb��Pc� "��'����B�(��9:p��R X�a���<���?Q���?y���?A���+G-%�Գsm�sH�a�R���B�'���|��x92�?�q۴��#l0!���Q�l?��ѣ��U�5(�x�f�j}m�?5�e��֦�͓�?�Y�!txLR���dk�Q�A�W�p���G�:&9���L>�.O"���O���Od���!�g<uF��6j�<+���O���<qS�i<�����'�2�'W�S:������\�>�V���2��p�	��M5�i=��$.��*�*5��kE=Obm��↙c�5r��Q=d$���G�Ey�OPdhQ��h%�Ӂ��2|����+�j�Ӆ������ğL�I��b>5�'� 6�.M?~����ȇ7�1Z����l��r#c�O��Iড�?��X��hݴ6�̜Q�j��X�>q8! J;&L�iŹi�^7�U�~{D7M<?q�j���B�	A�G��d&_Z^Iz�㖙t*Q VO�D�<�	�/G`�ɒ�Ѵx)d\��,��c���hӷii2��V�'���'W���nz�x��ZV����d�.�ZQ���1�M˕�i�*�$�>�|j��Q4�M��� n�2 `N�j��)o�(-˃;O�PaT!��yR����);�d�<�.OT�{҅��M���:�a\�&'6`�B�'7�7���L��D�OF���,^晨�H��bF�7��:g���l2�Of�l���M��x��
�0Qƅ,0��U�̚���,r��#�G��T2�����s�z�Q��p�B�Yd��"q̕X�h8��y��Q
t�"���g�� %_
C�.r�4���O 0�r�'6�-�i����� ���q�*n����q��+ڴTꛆ�{ӎ�xw�t�,�Eޞ���=8֔{�y�R�x��3��ā�!������Od�$�O����O.�D��B�~������zW��!F��6oz˓_X�V��&0��'���t�'�Te�`N�<~�Ĝ�Q�Þ.R �J��>)��i�,6-J@�)��>>$k�ߠ�UG�Y���t)P�u,�'�2�P���<,�n�`�	sy�g�	X��	@�
��^����mE1*fR�'��'��O�� �MC�b��?A0�E ��t�^+v04� ����?�W�ii�O���',n6�TǦ%�ڴ�Zq17bM�.Ѥ�D��*W^�<�)��M��'��ˋ����"�Ď�	�?���r�fm���V%
�3� ����Ɵ$�I˟ ��؟�	`��iq�����7S:,����������?1��DC��f_��D�'Ҽ60���S@�pk$�U�<�̉۵�B�U޶\&��:�4*���OKb��w�iQ��KO��k����8�x C�^4Z���B��c��C�U�Zyb�'�"�'v2�6�ك'�`K<,���3GB�'h�	#�M/#&~ �I۟��n�D:iT�2� 
7U���׆��W}��w�H=n����|��';�9�OC!��UA��\HVDYS��1R�@&͖)����]�1�yݙJN>҅3hm�X�c��bhH��UeM$�?���?Q���?�|�.O�m�t��3&bI���m�V�ؗ$�A�������ɻ�M��"�>y�i�b��d�$��ƨ�7i�4#��f��eoZ�N#�lZz~b-�'-b�A[�h�#!�I/�z���B,u��M����
`#��IPy"�'6��'\R�'��S>��U��d!4��..���+o��MK��Y��?�ɦ���~��LA���TD�:s���D�	��a���� M�fBu�*&�b>"D�[妁�D��%�3ų�l��oW�)��̓(C�u$���e�H>1,O6���OPU�7!�>Y�*�bU�D�a���;ժ�O��O��$�<��i n�"�'��'Ʉ�􉊴z;��C5h�E)�����A}�Ej��oZ��ēU�lX·+�.NA"u*!�S6��'��dz�E6��834����
��ΐꟴa2�,7e|l�"{��*���ȟ��Iş0�����D���'������^H�xЖO��h}��c�'L7�Ȕ6�����O,lR�Ӽ��m����J��M�^up	�<���i�J6��ݦy�5���mΓ�?�t�K�K������{}L�bA�$�����W?SH��xM>�*O\��O����O��d�Od	��ܸe����>t͐�1p;<�5�i�mJ��'���'��6�	b�U_V.�H�j�=(�f����\}r�f�&�o���Şw m!cg�;�`����^*G��uK�ヱyp<p�+OVۅ�ۍ ��������_�ʚp��^����{t�
3L�`�d�Oh���O(�4��Wƛ�ٺ[�� �ؒ��W2<r���;%6ތZ��F���B}Ro`��l�M`��?4^l���M a/
���Ƅ	~���4���;W.q[u��qE����D�,H%4AO��"�{���y6��O���O.�$�O(�d+�Ӗ(����@0%M$�Ku�T�4�e���� �	��M+���|r�>G���|�d �L1�8��hұ>lt��1a�GMOX�n�4�Mϧ^%����4��d� ���&d��?�`=RDś�H�||�!��n:j�P�(=�Ļ<A��?���?�.�;t���j���5#��!2�ߢ�?������N��	�i���8��؟�O�p� �x>�	�H�`�ƍ��O�I�'(�7mG��O<ͧ�z
	"%���]�_�VH��'.o�0t��	zz�8/O���(֝����}�D�A�u�����ծ+FI���?!���?��Ş��D�𦉙vf���xb�@&>�p��e��i�Y��矴��4��'���?ڛ&�T4J �t���ݪM.BASU� g\7m Ҧ�q�-��e�'&�4!ա\�q(NR�P�T3��?��p�c�+lE��' s��'���'�r�'%�'���?mP}�v.Hp��L@�Ֆ�
1ߴa�(*O���?�I�O�ilz�Q3�_%*d4�" �H6+���c����M��i�O1�&�#D�m���I7+5F��+�H��	Qud�/I�扂^��|�$HV��'�p�'��'�d	SbZ13�F̚��תu��=P�'��'4b^��Hߴ#�]����?��,���yq �OЀ��f�[.������)�>y�i_�7MA��<[�Z�Nȭ&�Dcc�P�z�Z�I�����G?R�Ny[M~ZsD!�u�M�O�0cʌ65Ѓ�Ǝr��C�O����O����OԢ}��1J:�8��Y0��]y�-ޝ���p�?��g�:)�B�'ߎ6�.�i���FCV����
����# �e�4PݴH{���b�Tm�tEl���	���M���C.XnHl�8	t���'�0�'���'2�'k��' ���2MH�w��hR�!��@Q��ߴh>q��?���䧉?g���~ #�O`���gV�.��	��M�S�i��O1�@ �� �� ��$w�5H�c��*""d"���)1� �z�4I��u�8��<�BB�Jo^�Bz��E th\�?���?Y��?�'�����9�+�֟�@eL�$cA� ����.3���
1H�ȟ�X޴��'���=c�Ƈd�B�nډ�l-��&޽K���-kTt*Ċo�]��4��$A�6�l�嬁��~��J��ָ_�@�Z2��fBH�D�e��$�On���Ot�d�O�D0��0��x2e��>���s��;���	���	1�M[b���|��#��|���yx�M��/�W����ˊ��O@nZ��MϧZ@��3۴��:y�,��@�W��h!�@j���P�Ђap`�G.'��<���?!��?2cK�q��@��Y�<�Y��?����C��Q�����	ɟ��O�n����X-zD�
�U����OF1�'�6�̦�`M<�O�i��b�^-)�-E�Nƀ�P�ː�$�N�u���i>�hA�X캳��|�!�R�r��V�G�S�6����Ј=;�'���'����]��ݴS\�ȥ��3#���q"�1?J$�6N��?��C*�V�d�I}��jӬ���i�5z�`�hE- H�^ő��ަ!�޴QiP��ߴ��d�5�B����!`���h��S��Y�H�Z�-��͓���O��$�O��D�O��D�|jRfU�
nF�C��2-v�)�MN?_��M�t��'������' �7=�U`g�-U�<E,4~�x��SǦ��ݴ ����OfD�	R�i����@�M�e�I6Q�f@�M+U���մ.�M�Ŭ�L�B�O���?�d���1S��%{�\����L7^��-���?9���?a,O�<lڨG�ʭ�������{Y�t����ߴ��͙/�0�?Y7U�t(�4"�x�KT�Lg�M����4�Iր�<��DS�3�5�拒�K�ⓟ�LdLr����n�ఠM�-*Lx��BSVƅ���?����?����h�R���!��U9p�j�&O�Lކl�C��O��mG��9��П�Q�4���y���$�Z�"�Ϗ�t���{F�ҕ�yB�w�r����b"�M˦��'��i�&!Q����H��Ǟk�R��ii�Ի���>'5�'o�	͟���˟��������� ���;% J`<�96��A��ܗ'�7-��v�$�O���&�I�O�hH0)):(JC��*�ҝbb �E}�Es��X�	i�)�S�2�]�%�� Yb����
\�6�(�<_vz<�'5ڴ1���;�뮇@�	gy�'��Ɛ��  �U��Ќsa"�'��'��O��	��M�P�
:�?R�������;p��hA��6�?���i��O�'��6�]ƟXmZ�8�b�)%!D�\,H���Q��������I�'�Fԓv鍭$kF�	��4�w4P]YĂ� S� ��� R�U(�'@��':�'��'v��K�LwrEòA�s���	�O���OZ�m�3y]0�؟�޴��5x��+g,�Z���:��LbFmJ��xrJoӲ�mz>!�E�Ŧm�'I�Ȑ�!ɟV�Ty�(���Q8�L�5F�����L���'�������X�I1_mVu�plVs�~�Y��Ǟy���	���'H�7튯� ˓�?�+�����ɕ�^�`$��a�7��aU��4"�O��m��Mk��xʟ�LR嚙+~5��h[?��m���$QBf�p�ò1{&��|���u�G;��!�p��'F�1\����`�<~����O���Oh��<q�iu��� �W�^���3�~."L�ጩ�'�Z6�%����$Jئ]�s��;x��K�mPTu�1hA	ۅ�Mc�i��(D�i.�ɳxU�U�l�W%��'���x���G���3�'Y�xŸ�'"�Iߟ@�	����������K�T蔣n�A�ƌM'�	�Ut�:7̓3ݐ�$�O���1�i�O�Toz��S'�!p�Z g	��qc� z�o���M�%�x��4m�.*��6?O��a�g��&�=p%rh�?O`�+��B!/�1�>�d�<����?I���@ʮ�+$�R�3����ٔ�?����?��������=�O�՟L�	˟詐ē4�<c�����l �o;���j�O��m��?�J<�r)J�&�Y���7/����t~rd�-f����V�T��O��5��Bl��h�L�r�*�'}j��ڂ! ��	�,�Iٟx��G�O9r��(d���B�P�o�ԁ2�)Δ}��*|��'��O6�DI����?ͻ�ܸ�D ��BDD8(�ϓ����bӼmT| nq~��|� ���Î��4rM9�N݈.��`��E@��|R^�����H����d�	��л���N?�l��P�h�t)H�LZuy��a��D�s��O��D�O�����d�(_5�qrh�jY���P�];����'��6�Rɦ���H�е%Ƙ�zg`�Z6�&/K�`��H�Q�� �D��<	��D��:�z[w�b�Otʓ87�� FΟ�H���i /� �3��?���?	��|�.On�nZt����I9b���!�&�F���-�c[�����Mӌ��>���iȦ7���iy��J����A���\+tK1}l�n��<���f�NM�GG�-��d�)O��	��#�M	�=8G��8��qyE���<���?1��?���?���+�?��� �9I���֢X�2�'�	f��ЪV;���Vզ}&��x�-"�4�󁃕Y���j�����K���'}��I_	8��6�+?��� 5_��pa,�mBA�ee�H�,�W\�B�8J>�/O���\6��O��d��wp��Z�G C�$y�a��~����O*ʓoe2f��?����?!/��)��'�/�4�6B�F-���������Oz�lZ �?�M<�π �8�T'�8Mr�e*���3�%��&�zf�d�S�̧i ��|�w,E��u��+�d������a-��MN@�бH�\�$�O����OR��<ıi�<A����:!B���)����������"�'*�6M4�ɥ���Ǧ�zA�Ķ&l�!�
D�P,P0�@��;�?��4��h�ڴ���#��i����)$( ˓*�5g�t-2����et}zF#m���'�2�'x��'���'�������!�Έb��Q�e �Ӵq�4H;l�9���?����O�x6=�h0(��� 
���J�ޗ_����Ʀ�����Şd��Bڴ�y2AC��p������R�. �@�
�y�W�\����.i�'Z�	ڟ �I8O\$����-p���ʅ+�05�I˟l�	��'�7m �t�P�$�O����G�|{�*��UP��x�����O�!o��?�H<��i�P>&��2Fmd�Y#��g~�g��%�I2 ��6Q�O��1�C���p��.(�X��6O�2Y�6u��A�^]`M�IΟ��I�����h�O��a�#�$)y,�%B1`����	gR	u��dh�O��d���Q�?�;Fq�7�R|U �)��P�\���Γכ�#j��lZ҂�l�d~R*�q/ 	Ѧ��0���þb�nm�IC�|�U��|BY�D�I����������`O�	 �C���D����dZyRO~� ����O��$�O�����d��y��y���8+#���ϐ��l��'��7�	ۦ�I<�|�"o]�m2^���,24Q�kֹ_ٞ�bCC���d̯]�Z,k7Mm�Y�M>I)Oܑ�aX,'��D�	f��hIu��O����O*l�Q��O�i�<1��ji�%��O$�K�]����k�?Q�Rj�ORn`�J��ɔ�M��i�7�A#R�%)�<N�*�M�1D��L�v�i�8�ȟ2�]�'dT�{�MiyB�O���� �$=p(�8�c�M�y��'���':��'��'b.����4B�	R��I�w�:��x!��'�2BhӴ!9R?���
Ц���vyR�;�8��#JO#v6&�2cA$t�.O�]lZ8�M�'U� ��ش�yb�'�*�Ӱ�(ƈ]1���y�l
�dZ�k�0���_Ɛ1�F��&zQ�e	 �H�%��ID�!!�G�H����U%Q}�a�1���&���i�$ҕ0��s��� ?ɉ��Ѓ$�Y�1y2JUɃ�ב�l��O�a�n�rP (5��hE���tȜ�a�,@��W�pI�V�L+B��9�6O�L6x�5��ya�d��ə�uǦ40���(�B�I`nہ}y��a�Ge�b]#C��:�^�yT��P�V��&��2<���kЗQ!����B��0:^4t�c#��`�v �e� ���b�Bh��UK��b:�(Xrj�y-�V�'�B�'���E0M�0pF+u�2���F&:��O���O0���d�O��D�O���.�~��4��i��^((7if�<�D�Ox���Ot�d�O������d�Ok�J�z j�X3b�;SX��ᝂ*�F�'j���\�A��y����ȧ=ZrM!�!2��1)a ��M#��H*�?1���������O�ʓd{r]	�_�bdq"�E+2�I��i�jE��cSݘ��<�$$�l`U��$d	F�ٍ7�}l�ܟ��	ğ$�Y����o�$�'��DE+L���!#�	\f�YS�DI�I�<�q�
�6�OD��'K�I��%0 U
#/L+�(( JKwj6��O�Q�!�<q#P?}�IJ�IH�����o������L�"�
E��O�Dj��c��I䟈��ɟ�	ğ�҈�+Y6� J�+�%*������J�o����'��	ퟴ&���I�����&0.��3�ȩU�8�a��kA\���7?����?y��?1�Q��a�O*��^ؙ
����8��o��M����?������?��+�P�tM�ڟ��1cJ�?�@�Ӏ� v<(��FX�x��ӟ|�	ty2�0 ��!���s�T���%V�|���'�,�,�m۟�%�\�I۟�c5n=�	l��h"� Y�w�R��6m�O���<�e�'m����X�	�?r&I6U��� �(< ���ē�?q��	�����ן6���\�;鹕� �Ȱ '�i��ɮ��(��4�?���?9�'��i��C��ט!cB0R���*i� yx�%gӶ�D�O��0�?��Vܧ� ���VՖ�D T�;��l�{ �Iٴ�?!���?a��V*�Ihy����[d<;�@û,���k&��;(7M#(���� 2�MAE�/_��EB�D��<{�i���')�)
�o�����d�OH���xh���F\΢с�N#��ɒ�D�<P��O`��O��$����p��6YFU�H�.>�<l�ҟ��J`yb�'N��'�ɧ5v.C5B�=x�m�}048�(	����6�T�O����O����<Ig��
�d���" = ]���g���Z��'N�|�'O��Z!R�"D��,�Q`���>\|��v�|��'.��'A�M�PQ�Of	�`��	Ot��� ��n�bݴ����O�ON���O� yp%��8�'�T�7j�"w��8X�<(`��>���?Y����ƆQ����Oc2�T�m�l0w��H��F7��O��O����O�Ei�:�?�d|(ŮHi��yд��#��6��O��d�<qt%������O|�D���s��4��rG#{>*���a��ʟP�IF�X��?�O�~8�
G4m��찣DW�0�R�@۴����*�R�m��,�	��,�S����ƀ��b�Q$d�ae�Ɵ:K2��ŵiQ��'0�Ɂ�d4�4N��������R1Ӷ(��?��6MEMr5o��(�	�x�S���|�DN��OM�|A�_�%8��#VN�8I���E�9��'��	g�s���ɯ�� �a�f�C��.����0�|e�d�i���'V�/��d~JO���O���|i!�� ;)qJ�H#�M%|6��Oʓ0����P?��ܟ�Iɟ�1D˟��<����tr5���M��Zw�� ��x�O�r�|2k�l���h3*جJxn���Ri��1����d�O��D�O"ʓ>�d�A��C~����,��6�� �O�`"�'o��'��'n�I^�H��E�33ҵ	����l��)�&h\����' ��'��V�X£잘���̂�W�Dh��X�>eXE�=���O��D#�$�<W�˝�?��
>3���6�@?h���J-Vn�������ݟ��'`D�h��6��>>��)iff*^<���;�@m��@&���'� X��'u�'A��Z@�I/
�h�Z'!� �f�lZޟ��'�r ^�
N�럐���?��0_&�уm�/G�Hq���ǫDOd���O���H�1O�Ӓsw��2Ec��Z�eAbd�	y �듚?a����?q���?q���+O�NJ�U�u�b���dXKɻ}���'��	�"�)��^����J�q���*TJ�>=i�� K�62�'�"�'��$Q��^��Ր�b	;IT��Ac�<h��Q��U��Y��2�S�O�P4��F;C��P�+�$z3�`���}Ӹ�d�O~��X� ��S�d�>�.V�B\�#!�+#:�H�R]�/�1Oj�!��_��蟠�I՟D�u/�/^ ��q���J���JD�M���o��02f�x�O�R�|��VJ���o_
)���䋨���b-l<P���d�O��d�O��( ]��Ζ��Ic�&N]l�;���'�r�'9�'��I�e�^肖@ˢ,���s�<qN� ��ʂ埀�'���'�Z���(���A�2X��
&�5���Ƣ͵��D�O0��?�d�<QD`V��?�v�ld�FYbR��K׹Ub�'2�W���ɘעt�O��[)���.e�l"��7�&���i��O��d�O��Gm߬<#�'P��jpo_.Cﾄ����b� !�4�?Q���^98�8$>��I�?ט W.~-Z���ܚ����2^7�O�˓	 d����'���*�#>J��0��"��]B���=�Ms,O�����������Va���	z}Zw�2�`�p��֨�)�z�(�4�?q���<���D�OJ�>�I�ŦB�R����י=���3��w�4UT���}��������?�J�O�˓+(0� � kg��Sk��Dr��i����'d�Q�����o�ؓrj1FE�|SJG&u�,T�ƺiGB�'��E�"!^�����Od�	?	Pmj�*�:�����k}:7�!�DU��?�����	T�:d��'��04��%�MӢ��4�?�񤁂=���_yr�'h��ߟ��15ߺ(b�'B,R�`񰂄9mV�M�,ϓ����Of��OPʓsPly����^)F�9�K��\�Fǒ{���Cy�'��ß��	��tZ�!_1,^b���#J$�Y��Q0�@�	@y��'"��'�*{�>��O ��X�+�S^y�
8+J����4����O�˓�?���?A�m�<Q�
��	{�D�V`݀v>��� KE�f������	ʟ0��ğp�oB��M����?ɰǕ�l�J�n?JNd�[e���	����'�R�'T��ןh#�K{>Y�O��#��(hШݢ��H=	� �( �i���'��	:7[�@��:�d�O����"=`Cp��m^Rp��_U��8�'���'��͖�������Y)^m���< v�p���-���n�ky�Kެ<��6m�OL���O���^}Zw=��(���"g��u+�Nƣ&b�\�ܴ�?Q��A�Ș�o���˟x�}2(+=L��r�Z�!V��H���ͦ��F���M���?���Z�S���'�Xѻf��V��(�1"#2h|����q�t�x�=OV�D�O���,�����4#	b�h�V�%�0��Ʋ�M���?i�<ք��aX�h�'�O�7o�W�D4�tO�9%p��#�i��'�6	����	�O����O��C�J+��1�
i�� *F+�E�I�6/F�K�O���?/O����P�ٵ��k6��]!{����дi2�\�y��'"�'�b�'��ɛZ-vupwD���"x�POW480�#�cU���ĺ<Q�����O��d�O,�"%/�L�ywˬ/5r��T�--���O���OJ���O\ʓ"�:2���Ï�R�<K`P������w����?I*O����O�d�F
�I8&��(��c"	,�P&�I�D��?��?I,O�5QA%\E��'�ƼCFn�eT�$��nC.�[��r�
��<���?!�OAƤϓ��i���X��'&RE*��[=-ȴ���4�?���[[a���O�B�'h�4bM2}H�Q�"��H��:�	�r��ꓖ?I���?	E���<A)���?�J�� L/r-�P�ppwGj� ˓�\Ě��ih��'.��O�p�Ӻ+T!�8j�*�L��&nZЦ��	şHRD�k�h��z��%�"S1��`O#�nx1�W�l~6�� N��m���P�I۟��S*���<Q�o7Ow�q'	f̡���� X^���щ�yB�'���'�����Itm���D�H	sR璣#5z5m����I韌 U�D���<��~򊒲d{4ȥ��%]*&,(@��7�M��?���'�
�S���'u��'˒ӆL��8ʌ�:p&��A�.ٚfD{Ӓ��Y>��'N��ǟ0�'OZcY@�,�dȒP�_�W䂵ðe��$Y0i��D�O���O���O�˓~g� Fl E�ǚ.�ՠ�R+�4� &�.'�	y��'O�I��,�Iޟܳa4h�4�`iĞ�R��J/'�������֟�	���'�\�R�i>e�tf��	_�i&��Dgi����?�)O��D�O��$�q��ƤQ"aN.k�J�L�Z/ d`ֵi&2�'���'�r�'��ݰ�Ex�h���O^�cS�DY\��p��Z�����Oަ��ϟ��IyR�'^.�
�W����$��"� �;~~-�J�Jlv oZ�������I�5h���4�?���?	�'O����\L����dm��v>�BƱi rV���I12P��؟h����4|�*���&��4QT��S�R�oEyr���r�:6M�O8��O���G}Zw׾Zu�K�=���QNB:Sz6���4�?���o�i��?,O��>����*�]����Gj0}3�	`����A�㦍�I؟X���?�����P�	矨(��=|�)Jn�51Xhu�C,��M�tI������y��'��X)�-�&[x���$NT�I�Pq��z���$�O��Ć�,~`X'����՟��V����#I7:6���K͸�ޭo�W�ɽt�F�[O|����?��.}�p��B_ډ�w	�ߔ��Ѷi�"G�=	(O^�d�O2�Ok�� x-�L��D�,�D�9�F�?LU�	?b$(u��IyR�'������^/6l���?18R%��Lv	b�p�6�	ڟ|'�0�Iڟ,�H��A/"�"���M����o�=� ��QyB�'�r��Ԫ�=J�8_�N�+t��`�2X���<n���?�����?	��r�^���o�^4��Mf�`+t��zE &W�x�	��<�Iqyr�dm���@@fa])x�u��A?q����桏¦)�Iy�	ߟ,�i���ē|1N��r'��e�6���W��7��O���<�P�E�l$�O��O!N���M�	Ucj���$W�|8�Zb�;���Or��Թ����,��?��T%�/m�<0�e��I�\cdӨ�z�@�°iu@��?��'U���@��, �"R�B���E@G~6�OZ�DNq��� ��)�?m �±�1f���")�}��Ə
[��7m�O����O0�	�v����ic�G:`.|�W������N�0�M�5�� �?�I>A��D�'��R!G� 	V-��i��'�Le3ElӺ��O>��Ƨ|���%�h�	՟t��\�F��c�.18�z�#�:qc*-mZI��I��\ZJ|J���?���nL1ŋ[�+�r�x�	�$T��v�i�2�U�:c�H��y�i�MK�@�**��+�'��t� �>A&HD��?.O���O��$�<SAV
2�Dl8w�ؿ鶝8��	5�^��t�x"�'Ҙ|2�'
���-9�4	��1db���J7��!�'���������'��!p��y>�#�On"�B�,+�}4��>a���?�H>i��?�@�4�?��M����(�t��|�s��yY��ȟ��IПȗ'+��a�7�I��	t�҅���*��"�V����oP�'AR�Ƈ~�R�~.��Y:��������A	m�(�l���I֟0�I.C�䰗O\��'�����5X�0��	N�{,�����.O��$�O(@b�j�j�1O��q?@�#��5[!���U��[��7ͧ<�j*v��F�~����🟘���G*@=X��TL�5I�);�S�~���0�3�D �0'��ӆ�85�,8C�&���DҺ_Y"�'��	�?-��ܟ��'!N ��*��h�v֍�n�p��w�h��<��*
�^<1O>��I�0��Iq�	mQޱ��2��iPش�?i��?APdQ7��?��	F?��-�x*Z��3HB!�a:�Ӆ3'1O�H@��z�Sޟx��˟�aK�4��]�$ʑQ�B�zA)_��M���mp���x��'��|Zc/ȡ �I��1���"�r�3�Ori���O���O�����ۀf�.�b�hЭ	�̽{do��qk�'��'��'��'����Cƿq��;U���\`�J����'��'y�Q���ב��tŏ
?I.�2��,.��1�����O��D:���O���R� >��8d�I���F�L� �����um|�% ʍ����A;>	h�N�O�"}�pdM/fY�	xP!A>b�2�+�I�V�<�ƃ���X5��>�T�C���I?����{ ��!4��2�P<��v�b�Z�ÜH7�]A�8';�س���'�0z"ֆ��!�Ƒ:!͂(������c��Q�yr��9:���;�ۜ;��x�Ú,�2�ؤhX��:��7�L�k�r���ǈG��m@�`�6!*��� Q����7.��2��l;��Ο�	Ο(AE�*�$�����';*:EK���|k�;�N�',��ð��/I��h���0����|��$ �5��I�o�(-Y�hR8KnJ���$�ڨ��+��B�&=���0EB5����w��d��A�0z�dtCQ*.0�:�M��M8"�'��)��<���:3�!���q��J��v!�ČR0����;�a�dйp\�����4����[�;��ٲ�CO'W>P�#0S<���Ox�0�r=b���O2���O6P�;�?)�>������#���eSy J铀���Z,)Pb˿<v��$�d�6DE&4"c�l�H	��\���ʊ)b�%X0iB�R�bL�/�Y92�!d5�����I�l�r��Aja�R��՛D��dJT���mo�$P�B�'4ўܔ'�*HPB@�O�b�O/\�y�
�'��D�v��\R���Fh�M�.!�AG7��|2���ٵLo:�  D�a�S(tXN�amW~���G�Oh�d�OV���?F9���O��S�I�@�����JVBÜ߸��6+�9�
���AL3T%�PȡJU2_�
E�0�I�9��Ҧ��*Dh���0/,t�dѱp��2+�����'<�~]C��X<������	)���d�O��ϣOuaTMO'�1�wh9ړ��OJ	��ӑL ͡d,��l�֠�"O\���i��/10�a��ڽ/�^�;�>O��oZƟ0�'v6�����~2����[=w�i���?B�)��JA�d߲� d��O��$�O4�0�
�w��hg�P�B�����S�Zuy�)F� ��!�f�˟{8��y�̇2�Q�<Qp
���$����GK8*�/�����s�.�g�2U9�&Ѽ 2Fd"D/��Q��)���OV�d7�;
\��%�8�u�\�`?l�I@���`%l�q��!�G*_ �Q�"a5�OL�'��%HI���O�x�Д���u� @�bÏ�M�)O�ʧ+�N�k��?	�x����tP�P�0���G�$8���U"x��z�W���8�E#K�Xqj���=ИϿs��ҕoL��sT�^�{h�8GC7����5"D�ps������DS$���/��U%@�}��n�zl���O;*�~š��A'\�p��&��ޟ|��P~J~�K>���G"vy����iڮj+��;��s�<w��X���fަZ�2	3v�v�'90"=ͧ�?ٳe�UL����L4R���(7�?��A�F��Ϊ�?I��?���O5��O��$
,�
�%��#}]VI3a$�>f�TSlN"Q���7�- �Y�ݟ�1s�����'�&p��cK	\טּj�I�����ɎcM���ǫq���(��A+���A	�EV�5�<��H٦}���É!~���`�nJp?qg����3ۓ`�Xe�3k��&�x��8��_k�<��cѪrӤq�Y�M�\�(?w��y��$p��e��4b�(�)��,B����X 7QVHk���?!���?�7�ȷ�?����4�N*P�W��zT��Ê�&�aV�B�6ʔ����H$IO0x)©\,�LDy�B��He��B�|���Kt�8� �i��+;*�X���s@�0���\)�`Ey�B��?9��i�lebCK׫l{�yq�GM��8�E�v�j�$�<Q�����	�e��g`��4{����V-O�!�D��/�\�z���tVt(��i?^��d�Ѧ���oy")��PՎ6��O���|��BM����@�]�i�T#Ψ�j ��?a�Fr<<{�N���&|i󋟈.�c僰?����Tj�#Yu�����3��$rZO�Q�P�aO^)n�$���ŗ
S-�ω���1�N��p]�!\@\y����o~Q�0����O�XE�$��
*��O�I�<��
�#�ySxL�;v��r���EF�0>���x��ןU������l*8E���E��y2��-�.6��O4�$�|�@@��?!��?��m�z�@�:�fүe��t)��w�n	�Ď٤	f�+�.]�{��ԫ�@��u3���;�L�:t\-o�ح�'��i�|�B�O��rWU���8O�@E�ɇ1/ڐ(����v���y�.�R���jV-v���j�'Y�u������	ϟ`F��?��� �l�6��d��ʨ~,
Γ�?��Z~)ᑉ֍K҆p�M�Gy��Ex�0��|r��θ��K;�T��äÊH�����?Ic$�1 ������?���?�Ӵ�6��O6mk�.Ey��Y!��ce���O�t���Ra�$�C��˗�0<�­`/:��M��\�/�X?A�%"1I#E��N���$@���൩�KTx8��_��D�M��#lO`%`7*�06� �"��,{�(�kP"O
pт�v��Ѫ��ՓC�p�	�C�h����|�(���6�O�z��m)�ʁ3x�I`��9$-��D�O����O�D+2���df>Yi���+ ����-7z5Ô�̔~���3�+ܜv��|���7C>�	�Mx6�vG�)�����5R�����O���'&�mk�앱1O�m�ᆝ2�`=���'��T����B�S��ک%�|�80eOX�ū�	��y�$ǣ��ei+\�W�倂�#�yb�f�b�Ĥ<9c�5�&�'b�S>�y��G5e%�e���I�R��SH�qV`d�	�����L�p4B&Y@���	�0g|@cR��-=�L���޵,�Q�T��֟G��J���_RޙS� ѱA(T���@�v�Q��c'�Of�o�M����ёv�^�k�`ȩ>�|�c��16-D�d2�)��<�r�,lŎ���.�td��P���O<!��<$M�� SOY*�|Q����<�A�V�����d�O���"��'�B�'�rq�3̌�kL�0 GH�vo�0�!��*�\\ȕ�p"j(��0O�SS����c�U�z�m:�i�*������1����O�?Q�����!>�@�3�Y	N���>�OK�B�@���"�
���S�w�L�d��O�@lZ��M�������҅=���Y ��0`�jY�h��y�'i�}Bl:q�P�&H�P?t����O<�DzZ>	�K 	�X�¤Ʃ=�p��6*�����	6O�p����؟��	ٟ �	(�u��'=
� \XP,�v{�� S�9� i4�O��P�'C�����d������_� ��'@�`�C����`�F�A�WdAuҼ��'�%����=�R-���Vt��׫A^�\a�A�N�<AEh�7!>�%`U��?Vj���
ǿ+{����P�z� �*ܴܘ@W�ؘZ)h����V ���?I��?�ЇN��?�����tK�;}4�9[!���ſ��P��/0�j,��1�ON����J(V��r�Ý4%�<3�e�4P7,� Ș��p>!�D������r��� +�]�pܪ���z��B��=1+���'L��mi�티(ޣvpZB���K`�J���4n1�ђՌb�p��4��w2�p�i���'��SG� ��j�~���*h�tX���⟠������Mޟ(�<�OD9�e*�i�2@rR�`8��ĝ5|�?U��D�(۴�c3��|<�:p�+� c�D�	�H�z�	�nO7<�̚�#[=4�M�"O)b5C�c�ѣF�nVy� �'�O�@��[?Y��CqO��Q��hp<Oh�`@*P�����՟ԕO�R�ї�'f��'sTM���w����%;����5��o8�mXc�|҈��XJ�1:%@��H���C�;!&��ՠ�QP�I�I�+,��Ә���랺B��#ǂڤd�0�P�+I�๻`�'쪓O?���P�$� e≛ұJ���.!�̟>�p�h�	a�Ȝ'�P�>�챌�4����ơ����	38n��d��}����O�Qr0ܘnk���O���O���;�?�;D�H��N�z�&X�&EQ ��U��@��Ǌ	V4��v!�}тn�3��= bd��^��$�ɢl�cN[#00�C�jzEǀG�^b������kv�09�ǂ���ɓe��D���O����X:F���[�O 'q�$�`�ˡ*�!�ċA"dC"�zS����ƱL��AGz�O�'D��&�e�`,B�F\E�N�r�dA�y�zDpa �O��d�O6�$ �8t��O6�N��P밂J;t?��X�	�^8��	��<�J9(���2� �"ǉx�'	,X� ٳl6���K�B4`��A�=-�t����4,�ȼ��E:uџ��!l�O�o�*=9Jm��eM_�I#�g�i�pC�	BtDJӊ� $�$pH4�U�!��B�	�k��%�t�U ��Jd���y��扝�MH>2
E�8`���'�2U>12q/
E����A͕	�2y�ѡ�q���������8rRQG�O<e``G�>�ڽت�Rͨ��ٌY�|�@���PXb������T�I��x1��<�8��OH����MT��MY#�8�z}��D׶ALr,-ҧ/�P��pm@�e%\�iA�3�v�ȓ
�2 �ЉB�|��g
��Op9��	���P	�Г6@�#U7�T��CG�|��<�ߓf�PyR�#��11vm F�E�BP�ȓ3�J����N5B[^�z7�L$~�~1�ȓ{� ��
��.@R9S��<��-�ȓA*P2��u|��Ǝ�,�ܤ�ȓq�ȸ4���H,Br$Z�xX� �ȓV��AسI�bT�T+�f�2�"�ȓ@L�Ɖ�	./Ba���2MaE��e1���'�[�>�af�@,��`��N�8��� p�l�Ĥ*#�^-��;�~��@(�F��wD�(/\��ȓr[������	iv�rs�G>f�(�ȓ	�>p���N�*����"oҶn��-��WH����E�zCa�ba�J^a��w�8�@�ͅ-R�� ��� nZ�����Iڧ�J�!.�86��0��L��h
H�0�dL4u�Ιp5�ǯa[�d�ȓGgȭK�5 &��UB�*Z���3Hla��Ã2H��0���#A٘��#�dM0��ۻd��e �H̖E�D������J��"f\��%Q�B�ȓqU�Ld� � AHʷC��%zpC��1f��Y�($^t�kǔ�JC��8Z4�!A��"�*xQᡗ�;FC�I�?5��`w�ρ
}fY���ՍVi�B�)� �ɢSǞ�rCrz�j��x��|�1"On�Jp!X�w����i�g�d�"O.�(@NǯW�X0�bɕ�)�B���"OpD��L=fP�@֨K����`"On�C���	F���'
�vB���"O΍��'�d�谒�t���y2"O�����jՠE ��ͼ�Xp��"Ol���9#��PḊ/���U"O��`I�qN�c�蚶G���S"O��:a�I,a��Qa��5R�f�p�"OB�i��C #.�� �K׵e��ykf"O��J0�Q!ΐ��F��Fi�"O����*>80�!���5�Rmr�"O�6�\�n逕��d��P�J4"Oh�*`"M�s��$1�d7$���"O�h0!��H<��ł$Z���`"O��G���Y��:��I߬ "O�\�iK������>,�U{�"O`��!�`�t�3dc�8-�v"O�1��*��w�0PZ��!T���!3�Ɋt���ʊ��I�5�N�����-�X���� !�d֝q���!"Hpy�E��j��>��c�"~"�\�6��U�'[�њ��*�yr�-%|�A��)\#�������D�+�`���I� � 0�D�T�6��L
v���Dr��IڴLP�1����@��Hb�N�J{蝇ȓf���{V�p0��7]�X���|�'�����O�n����	1}%x���'Q,-�u@:,@*��@&cx�2�',%vC�,�D1��*&� �'��	[�j��2k�ZsoR
v7֤��'����;t���G	o��`��'����́#���
�8m�JL��'����v��9,U2��hQ!�';&�W ]$#�Ќ-arh�za�z�<�nT=Cޢ�B���<y`Y�@Cn�<鵅݋݂p�r���*�x��rO`�<�0�^�C%����5!�2i�QX�<TBG�Q�N9@҉F.SOR��Ձ�R�<!���&=H0��!d'5g��SF]R�<��Z*]�~$˄Eߨ�.�C	�N�<�T�T.t ��j�ύ�4}���-�e�<� ��?���RR,�"pO��3 Ob�<a��AL����s��d����d�5�D�2��qj�  �pt'��Y >Q��Ig̓Bj���;M�ޭ�S˞�c4j0��D���j��_������J�>*�=YU-!�S�Q��D�fd�38�^=������B䉰W����Kǜm�@��é�,cj#=W�'p%@2�&ed�D��FԶ!ۈ�
�'l�x�,@=<C$�z���!H( ��4'�%��}��}�!�5q~�d�S��OH���	���q�O�0�Da�'��5����Kxn�1"O6�����N�T�5!5o(�&�O�u����O��;ǉ�I�Ys�џrL
����`�9/�\���A��BH��Wu��rJZ=��ć�6K�(IE�,J�x�[��	�al�+�L���y�G�U˛v/�|�@Ezﮟdk$N^�Ux�9۶'�B��� �-7��ˊ{���O�镥(>=Y�͒�Aj�M1����Ѕc��Xp4@]�a��� �K��Q���'�M�~D��O,%rD��gF�z��=1'����|1��E���$�1g�$h�t[U�E$"��JVEق^�6M��g0�O&��Ք?�>�����@�R��N}�@�ɼt�8�[�E-1���gy�������i�B�4|CF�ä�R�_�N!�EA�ay�A�@?L�@�� ~
��gYŚ��͒z�Jh
�� t�PЬ�Z0��ORԤ���-�����0 �B��O��[3�F.uݰ�dH:GL~���x"��4�� %*?�V��!�
�
 c�x�౳n$� ��1�ƑM�@!�EOA[j�Iɥ�'��Ӡ�t%��<i9'�0� �6�녂E�Q�D8��Ɲ!�4 �g��H�X��P�75|�YBL��<遊U�TE:K~����X�j����>L���שP�+�����&�O��:��("��`5�X�%fR�YX : 3O*iA���BoS�Q��<Q�!Ĭh�<��a_�"䫧e�.z2D��)�0<�)Om{v8�g��~�^H�4��]rT`q�^���@���<��ᑥG���$����O�UO��1 � M�
��w���t�e$&�`MSA�@&5�TPh��>?�����V���L��
6$��BH��1� n��<��G�l�r1	B/u6y�Q� ��	#a e�Vo��Zup�e,r�>a��m=�`w*[2.���B[f.��Po�;o"ca��#_ �5�-��bs"Kç&6Д�" ߚ=Mz�k�+�>[�F�jf]m����4��@�7-M���=�b��?D(^}���}��d�1n���ܥD%��<w�B�R� ͙�]�4�H��i/m��c��0<�Bj\+xh��O;	8(�"F(2n
����G: ��9Y�.�,rB!ba�		hSh�'� `e�)(�h�t���eja�&/���� '��B�	#���G�+]���R�$U���:6�Q��@�S��v��u�g���<w	^nwe�M�	|����[���I�0_4���`ۺ?q���(=.��>!�iH1!)��Ö�TU��0�`-2�Q.N����a����a� ��ˆY�'u�D�)1a��7��I#2���dڮ�P�@D�R�f���w*p!�c�˿#�f`:��ߴ\kX	i"�y�k�'blm�7�����Y��EFQ!U8����A�!3�$��n��i�&�Q�T8��B��ʛ%�4��N�z�I!V�)�Z�
�၇%���:�,���D�T�',���T��yJT� ]����'�J�a� 6L��+3����l��O��SnT=a����5gN��8� %�2:�V�Sv;O���#j��v�IR�U$`3�ʴ��@��cǾd�\D 2�Ή���c�7̨O6�2T�O�F��rC��N`D��c�u�+ps�(̣�NՃh��O``���ap�d�OۘY�&�>U�as F�7��(���,�N���$S(a٣�@>^K�iX���~E�H 4��O
��L+�)��O��yG&T�XGtH��暋;�rӉ��0>��e����� "JcE��9��ՠv��,9�/H[��I%�,;�'X��H3R,�s�\hc!�?�h��O�p ����C͊[���B���
D*�r$ �K��KݪH���O���3�))nY
a %a0g;��c@L"���� &��q��
v��#?!�`�%+�V��%N˾���{}�*�>h�b�rl
l�}���r�&X�F�Ȃ�@�CJ��0���EIv�<�DEGz	�BH�O�h5�"���1Ġ�O�����F�<�@U>�z��<a*��EU�u�iASB�4'�Z��$D+9BU�iF�D��uh�΢&����O��?I� L�R���$J�B	<~qOtе �.35�E��ٛf�\�p$���Et���4O��gj�aJ3.��S2F��%��!k�=  L�@~�CL9k�֝��	%O�4r$��R�r� ���c	htr��On`Z��s�'&� ���� <�씑t-
�h˔T�"��F�X��C�x񢷢�/
�PL��AЬ24�-~#��դ ِ���=<x�YU��w��}�5g^�ԥQ�+G�S��+
�'���2�EB��\��Y����'2Lhf�6�OU��ၤ]�&t�6�N*z��v�'�����H��x�$U*a�d�	�%�)?����:D��(��K/F�u�a�4!، 17�X ��G�$��%%   Ꮣ~L3Db���y��LBJ����nN>�Y����?����z����0�b���}��9X�B$�p�Rs�"D�h��.'�p08ֈT���K$?!��'�<��df�|$�m��B�ZY	�'ⶕ�a�3z��@�P� ����'��]��oH�_����˕yp����'��
�oo��`�
8_StY��'��5�R�M�rBЧ͕�Sv���'F��҉�t����)Rzy�
�'
pI�mS�FQ�X�V�ŝZH8{
�'�~Iф/R,H�5�vc�)RDU

�'��mCcJ��G�DyX��I�w&��	�'F�� ���\����(�5k��Mj�'%X��$��4$�P���f�i�V�B�'N$Ā��R�(w�A:f�f���'���u�13<�$���~�< I�'RAx���o���R�I,i���'���wJ 7j��Gēc�
�8�']���f6���"��)�%���� �p����
�\�[W-[�D:�@�"O�xZ�ǌ X��qu+�?E)�@f"O�)J���㪙���O�V�E��"O\�Ů:-n"��t�ʛ'��2�"O���v⍕ED9@b)[��4���'��F��Q��B�?
D��'�D���<.��"��� 5l���'���2��5P����O�O�2$�
�'�h�rv��!�0���	 r�J]	�'T ���.@ Q���I��oy�A��'�X�c�����A1
^*y���)�'x��뷠W&9��U�SQ�v��l	�'n���d��:�*�����i�8�'	Bt�'�J��ls�j2ZŴJ�'���c����dؑR���H�'`Xx@�ש'R�I��F�^����'�J�� F�KaR���"�W�P��'Ǥ�@/�!'��� �O�Y��'?��nַh%PAi�#Ӥ"�Yk�'���+i�($�|U#g&�^H8P{	�'Hz� ��Ryc��Ni�X��'�]z��ٜ��jB�N ��'SD�e���qj���uG%u�q��'�!)�iF:@/n����\�5R@X�'���H��>{���Y��Ï)�( �
�'���S�m�f��j&�E�
�:�'׬0����P���6xU���'Cf�1���:�>\�o�\� r�'�:�9G��~��и�ɇ�SKD!�'�r�'F˔]�J�V�l���'X h��T6a�^1p���&P�2��'o|�*��ŝ^k�(Rǡ��@b:q��'�ε�r�U2yz��I�a�
FV$���'���splOd��x�%�K3ܵ��'�|��6kC�UZB ��
?��Ÿ�'K|4��ŕi��<C#)�1D�}��'Z�j��G�c#�]i*��^��	��'l9b##�A=k%e�"P� �'�@)1��K�2�����LQL(��'�D��� �1��� �SFP�l��'�n��Q��Y9�R7��
=:�X�'��-s��5�:���/;Mr�'����HZRf+)Ql��'!f�:��
2&��i�aۻmT��'f��7��*9svpC*!�l��'���`Z�$f�0���L��'`��jƋҮ�7��F�����'�z�"�c�8T2���̌/X��@�'腋 C."&x���`�$+HJp��'�*�*�b�	i��)kGM.#��r�'�	(�\�Rzŋ��O�B �;�' ���ųz��ᅇ��x����'6�C"���lD��/+�6"OpIBR�X%!��uk�7.L��s"OV(�2�5XA ��̗�z���S"O� �s��&`E���ԥ�;)�I�"O0A�Ʈ���n��/�'|N�{�"O��P�&a�IMHT�d	v"O�!�5$̐*?�` �>��"O�T��̠>%�M@�Jz{D��1"O�9!��K9)��ɢ��1Srn4j�"O2 (5�\�2��x�'���dT��+ "O���m׫fML��dj>�F�f"O�	H��Y
|12�+�OC�e���"O� �EY1�܆9xn�������z�"O�z7��H^Q�A�<��T*U"O�QbLO)8l��L��� ��"O�u٠��:[V�5�b��"Hk>�0G"O�M)��v�`x�V[�a"	8�"OZ8
�����R�~hx��F"O	���.�B B���8�l�B"O���%33NԛA�4#S��iu"O�i�iҕM����ծ�I�iJ�"O�E�梈� ��`2+K�=c�Q��"O���G��6]����(v[N �"O^��c��[�TT(0�,r52Mp"O�C��Ic�Fuz�	0*Ԅī�"O6��� �7ߴ! �e�r�"���"O��9��Ğ���фEK/}\�(h�"O���@�D2�4#���|�0�B�'51Ob��0m�}����b����d�"O��)1(Ѥk��ub���.���!"O�`q���T�N���1 ��""O@l0F�I������&!����"O�Iv`�XPT �����!�"O��j$���$x�	���ds��'u�OHxQr��{^����#p@\+F"O����,F�h�D���U�/P�I��"O,yA� =�&ȹ#c�Z7X���"O����ɇ ��=�Ӏ ��r�"�"OT��U"J��	��t��3�Ȃ��y��ŗ~,�8�D���&ajqp$Å�y�K�U�� +��"؞�G!�y���"� �A�MB>��iC��y�C(EM �`g%A),��+DI��y�l�W�R�;��AM��8ԋ��y2�&c����Rg��.��i��E���yR�vcj��pd�q�C!�-�y�섕:\�)�6+�%j ���M��y""�Mش���d��`��A#�k�5�yB摥Kq� �Ɖ�V�F1�'m�,�y"��7k���E���(,Ɔ�y�$��Ih�@�3z��9s�[��yR����t-jt��q�;��	�y�*^�J~�3!I���Q��Q��yBKK�)�l��T��d�c/�'�y����HE������"���yB���EX���k_�=�F�׫�9�yb�8@LL\���֘(.�A�Ȍ5�y"c�iʉ���wI�	��S)���/�S�O�.�K3%҇;���e�#j����'(蕫���?B�����b�n ;�'�蠋`��P<�UVN
�9�'+2AD�9=�
PK��Q��)�'!X�����5*��g��8Լ��'�y
���>xBU��*O1Ja1�'�� ��˴Q0!�Ʀ{��P �'��,ZՏ.-��)�a��s�*���'��Dа�D?+��1Y���p��0��'P��"N��|@�L��3�(-J�'� �s�LA�2g��pP���,����
�'�����`���\p@΄){�iZ�']4��Ar�t�G�ȸ��3
�'M�4D�2'2� ��Ώj�m 	�'1����5Ԯ������d��'TXQ�ǌ\+d�!�-��{��x8�'�@`U*Z'f ű�N�-H���z
�'�t��ㄊTʤ��Ɉ�G34����� B	�d�T r`t#pB<RytEz�"O�T ��G/1� e[4̌�^l�d��"O@��ǯ��d�fE�Tˀ�:�*t"O�`�.\�fq���Ƚ�LI"O����-�-�,�Z��
��"O�+���:��������05`ћ>I���)��Z��&���x����;�!�d@�#0i0s' @�(i��O)8!�	�]"���`dţh���g�I��!�U��)�c��$g[�1X8`v!�D�U] H�Vh�R�<�1A\�X!�D�:h��Wf�";��
q���!�Q2*u,1
W
(I�����Q�kt!�3� 	����	_.�^a���
�'�l+���%M:��ҍƶs`��G�?iGz��ΙI4C�ޏP�!��S�y�	=1k�͘�酓B�pQ���7�M3$�`������`�TM؞i�(%���U� �a~�]�pzw �K��)!�i(mA�,�C<D����$O�j�QsiІ#ق�f�8D�X9��JO��I$*Zl��$[��6D�褭˥$N͸��D�_�,<�&5�~=
���_�,9�5�_l�H!�!#`�a}"�>�W��
m�Tο]ߢ�)����<)b�'� I�7)��qm�l��+*J�H
�'���:�@]J�"���O6�����'K̐�Ug�"A�v�B��"_�����'C��%\$fb6���g�'Z��չ
�'H@�ӐM�k������I�Wi(��ϓ�O�m��왲t������_�j�pR"O��V���qli�B�R(.��"O�	���~^p��NJ�)A"O\IВ�ʐNk
=RCN�4n¦��"O<!yض.�C�̈́'P
�| �'yv�I�B <�%��J�Ur��I�c��C��M)8�[A���/-p����RN�4�=!�%]�ܺ&d <���eV(0���ȓ�t��#��f����cO/%��q��y��S���P=x���(�0�ȓM�d3�JQctB rG���w�4Y���0y����(=�L�e��"js��ȓ<L>+�*	�rxZL����Qd������4���)eF�qR#ӄ;���$���w�I�4+�ɡQH=X���%��rԮ�)7Dmi�K?I�����&"V!sp��(R1��d�L!B��`�ȓH�D�V��T�@�iŇ}���q?��*��W�ZV����gTJ��ȓ4���T�כ|h�೒�Q7d�δ��8��� I\b]B���܅��$�,X��6�|݁₌1w����ȓk�,����J�r�-�Գ�.��ko�\ⅣP�'�ՠ�J�m�0x�ȓO���w�G�GfD�Dɱfo���9�`p�N�&s��4�D�*b�4��ȓ�T�lS�-j�	0���y����ȓ,nL�p�
ߐ��Xs��<H�$��ȓ_^e�F���p�҅#��C�z��ȓr���H[�:�8-�� �h頰�ȓ/8��pާ)T���c�ѬseU��2X��[���!���h�a�^�Ʌ� ���#a'��n
�yp�_�0��9�ȓe@.}A⨑	�"A06�O-$�r4��z�b��dĀ�E�Ԕ[]<D%�<��)� �e���$	B���w�ƣM]��b�"ON���L�������?
Kƅ"O���`�D�P�|��A&7���"OH���ȧk�������o�t��t"O�fG���p�c����y�"O���d�ު����w�� �����"O~D�P+�&!�t�Y�(�+��y�G ?d�2 V� �R	r���y�"޷h�f�� �n�0Δ��yb���R���h4�� 0j��y�ᙎ.��׫�c+h�H&����y�K�^/޼�	��_���$���y����`Ȕ��
o[,�8��1�yH�&:L2p8��Y5kf���#Ҋ�y����%$��ɦ��4h�����杬�y���?�p����=g�B�-Y*R8�ȓ6���ǿjmJ��H�6|Ƚ�ȓUa���c�j��	+���@�8��cyA��aG R�(�rp,�f9(e�ȓ]�������\�j!cQ�s�u��2�y���:�@`TK u��!�ȓ��a�PhX!B�l�kt��	�݅ȓZPR��]nQ 4�C�.Յ�\tF �D�� Gϊ�C��
A�=�ȓQ��Jw3�L�*d��v����p+QiC��2D�̭���5o�JD�ȓ(��dIEd� 
"��:p�*�@�ȓ+:�3`FUm,Z9Z�N��v� �ȓ6�q�gl%�͂._�D�ȓ	t%9� �8���f=��U��O�����菽*���A�>���ȓm��H��I��	c�	���ȓzŰ�z�/�24����_�Z���F꘥�E�
w"l$yn�4��5�|�7�Yo�U�4��ti��ȓT&!��)^�;����f�&U��]�ȓ&ih������]�`8��bY#/AD8��D�r��p"W�H���c��
9c���I���̕ 0 h�@f��U��[�bBv��WE� \���<'6���6^ZN�c�)��G�Ɇȓ:,j��Ң �|�{�S����ȓ~�lQ���.�f��Wm_5OZ��ȓGRșH��Y2q�".B�t;���mh��B��2��{��ۼ1<�}�ȓqj�,�3(ř-d�X�R���6x���P+'N�n��a��0����ȓ*8a�SO���΍"`����ȓ/l.��5cE%U��(R�߅b�<��O�Q��hQ$MY�m�D��gJZ�<AC�ƱD�2��޶x�%��W�<��,F�S]���P��1H�(�kE$U�<)�%ې@dH�ň�w��P�#�C{�<QЍB'v��Qħ���̝����x�<�!��{� �	B$�0I�v�
�,�x�<!�C�4	�� ���(��^�<!�
&0�J�
Ūa��+ծ�X�<3���7R�%�W���K�H�\�<��®m �@ӈ"xh���3��U�<9�#����#��UG��g�
Y�<�T$G�
9��CG�8J�#�n�<�ì� l|QlБf�P,�,�g�<���ХMQ�%S�JJ�a�T��!h�<�oݞ3ͬ����O�,h�6%�_�<� �8ŨӜ	����T�H0-���C"O��6Gĭ\�&�23��.}:��"Oy·g����YVl˅d_�qA�"OfU�V�K�W0��P�Q�ZXM�F"O�`CƔ%�nlٶ��+�ND�A"O��2Ǩ�<>���B�T�8�"OjyY��Uc��*��;'�@!
"O�p�dA�+W���h1i�=;�|�P"OJI�*8t�X�Ǐ"V���"O�7c�%#������VR��o7D��˶aПO(�A�R�V8S�-��:D�|z�i��u� ����}��a��L8D��  �4*�P�[�&�c����6D� ��¡t���	��C.�ڗ�4D���d�K�t1Fh���!x�2D����-ݘ/ʴ����O�(m�isJ1D�!AK׵����?��Ⴗl�=g�B�2&I�iz�J��E\x�v��/z��B�	�8n�J��*z�F����U%r�fC�ɑ`'r����=e[ ��ƀ���B�	��rA��J$G�X�ɗV��C�	g2:qy&,97C�\����H`hC�<w^����	Ϛ���� [YTC��=Y�.5"bɳv�|pb��ȜlB�I.PH�)zhK��R�a��Ȩ!�B�	 z4����,��M��)(FE�ͦC�	?y �K� &x2�P�E γK�0B��8q�ͺ�GV:`Z��e#��7��C�	Y���
c �2$��L�YB�	�Мl�ÉƯ=
��E�߮T��B��4?Vȅ���7���+�+J�9�|B�	�mݒQZ��O:K)��k4!Ȇ
|�C�I�/a������(P�L}�"��'-�pC��4u+���pgj��C�A�,D8C�I�<�N��7�5fzȻ���C�C?�Բ�-ޔ9�x�)�-A�$C�	�/� �c��ހ	<�R�X�E_C�	0	�����3}&dA'L�&�B�I�Z]�i�ڳ
��]!`��9K�C�,8z<e:��L��%it�
/�C�I�/>`��V�R�q:�m����C�ɪ�j��ܒ=n�	��͇_�vC�	 0d�z�fM0'z�8���%D
DC�	:(��a�Y�n܁"h\�H0C�	�Z�\��S�\�W����d�[�~��C�I-5���WK�=��!c헋OYhC�I�p(r�{we_7]�j��(U�^�\C�	(G^D#s��#v0�aT��HC�	�>�B��K*}.�F��:W2C�I�6v\����L�Kq
���MQ(RC䉶y(�	�-K#ּ���؄zC�I_G2�rR��!̖ĳFk��<�C�I�(��p�J�nJbI�;l��C�	*&�����600$CÜ�;��C�	�D�Q\�.��=B0ď�}�C�ɂ	S�<s(X�m��튱%j�B�IZY��:D�šO͸Y�jU@!�B�	�"��\�V���\X�nճ0�pC��#6!+p��e4H�CΒ#F�"C�	�]�rM���E?!��h���C�}W�h�(����c�_-�B�"=Ԝh�A_)v��=x7�d[�B���U���|t����?�n�s	�'1l(�挌D��<��Ö>M�40	��� ���荾��`�P�.nx���"O.�R !ΤM��(a�K�;�p1��"O<�S��K�70�����dHr�3C"OJ��5��	��8B$,G�_b~]��"O��P��3��\9BJU���J�"O@���F:���޼ �dQb�"O�eH6'F�!@��$HC���В"O���𮚂7ƈ��Gmd�v"O8��Ɓ.*���N�<��Y@�"O���X�l���6��?�=�"O�Y*��m]8��	 (CFE�"O���գ[y�T���96h]��"O�Q ��'kƙ��#*�9�"O^imSCCP��AKZ��"O\|�t�߳~���W�\=XcPu�V"O�]�#-�Nu�i0'�1'���3u"O0L�TMH�~z���R�0��T"OH\`�Ȣ{V�i��G�a��и�"O���A�@.D�����v���R"On;&�֋<��9P�Y�j��$�"O�8�dA>s%R�0�!G :����"O�xA�O�'����F��Vh6���"O����#AT#'�~N4���"Of��2M���Fe��Th�,�y���`�B�"H�~o2�*ӣߕ�y)��1Yّ��B�Zh�b�Q9�y��B,WxU@f^&#3 �I����y2�	�G��]�	�EJ�Drq���yr�}���ӂ֫Et<qC$�y�e[	��	�Q
)T�0���=�y���	(�t���٨z�����:�y�o��p�D=b�G���p���y�n�����;J�/�����y"��Qz*8q6�^>��Sf	��y�#�rb�a�H*ONH5+�� �yb`�01,J���h��D;�鰢m�5�y���#�N{5�t�F�W䨆�.T�&�!�Ҭ�c�T3�Іȓ8��@�3OA)^�M�ScWv\ ��Whh�K���δ`5��4��2�Z=@���O3�10��o����ȓ��y�Ǣ6����c�Ɯ3�t��E��XH��LR'J���g�r���,�cTc��j ���1:%�ȓjޤ*�΋�{/�՛/�n�����9,	+e�E1my�d+$�PQ�M�ȓ$�z�Qf�V�C^�%C�)��7)�t�ȓQִᙀ �$ L��7/��M���ȓsY
��#����Y���-/r���C��s5��$����ޡ7w�݇�#ztE 6f�1%�������:hI��&�fL���n�*���&9�	�'O� H@+;3`(��g?@2��X
�'7V����U�(��,q$��;�$I
�'�M�v�>c zĩ �B���Ę����.��?��Q��_'!��ikF��6ƌ�f�&�D+�Oj9!�N��ΞkS��"�t�b"Oĩ[�O��H�X�Lb��ihf"ON��V��B�";iZ�e��
"O$���R�Zh3w�V�n(��"Oa��i��d!���e�3ĺya�"O�=�b$��F t�'CF������'(��'#�Y��'R1O�BSi�P;d����mA�"Oh�ѩܬ[~�Lb Ɓ���@;�"O� �|��-8P0*�%��^���V�'����#s��H(��\N��F�L�8B�	�N���s���\!�ͅ4=0B�I�Դ�Ai�5-뒠	"� ^4�?i���"&DD�QF�̿l��jD^� }��ʟ�?!���܊��{RAU?@�,%���,\!�$�)d
�Is�;'��I#2��4H!��X�lY�ujr@'e0Z�I��?@�{�D��z�le;n�(Sh}�(�@!�
���H�4�� Ó(@ %!��AB�I��"V�%.]��&% A!��Y$A����P���%ؠt=��)��f �UN��Wr=���^���U@�'9�U�ѿmk~H �����T��'��h�J��	���H�F�Pa����!?�P�>._�r`��&d����I�i�<1B��5�P,�e ȟ"5��.�i�<�7��P9,��k�6z�v]�V�Od������@a�旜y9���d�D><L�DҶ�8LO��xDǋ�-p�R�̓6`zQBu�'�b�'�ў��<IE�4���C�^���SDh�<��˿y�|p+�,�j����cx���Iٟ$�'��aͨA�Di�L_�l X�'и�T)R�u�t@�̵+�'A ����ֿ��HcϘ�	J8Dq��$�<Q���M*Ҽ!����`,�%�X�[�	���IZx�X������ ��3�L�̜����O�<yqJ�ܡ�E.9�ʐ+P%'�On�r��Y��U%�Q�җ9%�I���ԟ��<��O#�L�L6bZ�����a�<�0��`�\0`��2T)F%{e/S�<�3C��U���񪃧E����Ehw�'�?���i�6��`�t1�&�5~��v����sk
�~�4Q�	уg�pl��6D��p��;�$�B��/d�RPc�9|OH��/?Qcޭ;��E* ��0��]ІHY�<� �۝���0��k5�U`ŃVZ�<	�H2�M��M��9}dP�WGGR�<�䡈�V$p��78ʈ���IO�<�&m߷y�4�:򮅲�,e�A/�G���hO�'��(�?r	��EF��t��ȓ4;̍!�Hܷ\�,��E�9[�9��Iby��p����>;������31�fL1D�\�'���ev���;D�����\.��"��Fb��g:D�jU�E<R�5�G�C��|�@�-D���F������M=(��b�<q���S�1��	��C�Q�����b��<�B�I�U$���QnՉEy��4K�0�nC�	3
����	�'ZY�}�g��(+��C�3a�*=�fn�=0hh2J�G(6C����h�!AU@���^3Q~�B��/<��	���[�06����0lϖB�I�=R���.��R� �)�#B�C�I"0�<(��jߞoW�h��­B�DB�ɼ1�3��Xa����%E>)5*B�ɼm�(L�S�ՂU����꘷C�!�*��ȴ��>n��bʘ�Q9!�D�),��} ��i�
�ٲ/_�!��-2�m)6O��'�u+�m�>K�!�O�U] =�D��X���Q��O �=��>Ux�x���3P`֤K"O$�ڤ&*;.��!��Td��"O�Ġ�i�rr0Xe@�%S��8�"O� T	KAa�&�� Is�G�g;�U9�"Op�X�i�,����%�k����Q"O6��q�]mf�2TDµCh6���"O*��Dc��DK��;b�M���%"O�M��
a�+UH� ��P"OF1��KL7N�������zM����"OЄ�U�ì�����a�n�1"OU@���l,I􁆑7����"OFiC!�*��ıu �0H��X�1"O��jD��1Q� )�'N)�@D���'��I�A�h�S$�%:�����6Dd�B䉱n�������(9)��N	(��B�ɉw�X�@��]�W&����ƅ$��B䉤.yF�(g�<VO8�A��7�B�	B?�Up��
!'J�q���B��w*0Ї���N��B+e�B䉒|�U��G�F�,$����;tn��d-�Y��t��Ȑ�/�&X�a�
�i�C�	�:���نA��尠
U�F����x��ɤd���Jp�-6|���A�'�C�ɘ^���
�U��̻F�Y�f�B䉀RԚt�7(ކP��)�"�W(nb�B�	��x�"D�3��U��(�-}��C�I5}/�,#V�ήF x��.��tu���!k���bG�իu���S�&�#y.d�ȓF�z�1 G|�cP�&NXM�Iwy"X��F��'��@����ZDT�u��'C���'�( :��Z�bh$dg\�>�Rd��'Mf�qs��	8�.���o �:���Q�'E���� i�n�s&Q�CF���'�j�����uAT�Y%$��%�� �'F�q3��}E�Y⳦O�`���'�"PƖ�q���mSJ����+O�=E�T�#��c0o�@S\ ��$��y¥Q�	~�T(�@�
<[��&��3�yb�	�8��!˜�.� E#�6�yB-�Zx*���{LA�7���y��\�[L�u�&�J�i�L�b�B��y��K$I�|�x7���d^�����P�yS;u�2lB���dQ�P����y��;nV���oF�xq`�O���y"-�P��x�G�ϺS<b�`�F��y2$Y0�8Q���Q�6�rl���y�dR�y�%b ��0H�ne2��9�y���%�|���&�:@XtD[Qǆ�y¥�[��tˀ�A�1L��0�W7�y� �[J���U�
(;>4g	���y2n�>L{^��.��S���fHU��y���>5��(��*�X�>�V��y2��2�������6}�5ʵC�y2LҒJ%��)�H؍u�8�R�F���y���-pW�5k`�g%z�bĭ���y�"�Vv�z���bU�L!Qk��y-M��I�I�VN��0*�$�yȱ0Q�	[�-Dٓ�HT(�y�.A M�BXY��P=\9������=�N>i�È7Ft�4��ԇ[�>1�OJ��yr�N9�X�ő*T� B��M��y"�'��E����F��	*�Jԑ�y�iճ��0�͈-C�@ ����y�� �Xn(�C@[ ;�M�1#���y��"�nՙë�1[��Y�-^2�y��ȾFY�Ђ��)L�lz�^���xR/J�$�|�a�o�c:��i@Z�!�� �ia�P"b�H�h)K�HU3"ODX��R��d���M@ @􉰐"O$��3f��;E��H�!/��4"O�]�W��*xp��
�2�v4���'�ў"~�2�� "e����&Nk�\��̖�y�c�!Ģ�8ਇ�w����2�>��?��4�F� �P0(7b'i����'�(�a�o�S�~I�ƛ}N`d;�'/�C5e�#���R��cܶ�+�'�X�0���H�����&�D��L>	�-�T���H�!1�]P3�)��'�ў�|.��"����
:[��{�DL�<�s.�u D�@<P� p��s�<���G_`�QE�o���Su+i�<ɷb6Q\1�l�� ��p��!g�<Q�킸o�H�u�L\����cPyh<9O�<SƩJ�Ǝ�7���(u��y�ڪ8o�`Sᤁ*(��b���"�yr��L��(Q�@5�2��j���yBJJ00�\I�c����<itD=�y��Ao���Id����X���ϕ�yr'V�rS� -��@dS��y��Ϯ`���r��A*1ulK��y���WLx���l}��H���^��?Y���0?iEAL�J�`'V4kʜ�@��\�<���7\`�x0�`4]
)��m�\�<	�Ċ�\tt<[W��v`��}�<Q��5gv���$��8?mHI�a�x�<Q�*�`��+�������G�r�<�b�П\I Y�=E���j�˙V�<�aN�#\찬XcF%�\�JE@�T�<�1G��4R  5��?���ѡȘw�<�T$�w��8��mέ!$0�@m�u�<q��[}����4F�^��EA2��n�<1�͇�#h��� ��on�t2�Äi�<)�
1s+$�iaeɳ$�A�Jg�<�rB�?Sn
�p壕�l��\�рV}�<Y��<J���$�>K�X!v�qy��'>x`� lܶ�)�@�"6Xh�'��`�F��A�>�Z���Q:�8
�'p�8�Q�:Ah!�I�%e��
�'t����	���UJr��,3 ��	�'�r��e�Q�v�b��LW����'_*�����66�n�2���M*!��'�>�1qM�0jeh��n�NɻH>y��?�Ó�!�'�Y�X����ل�:�b�0�JѪ'EJ5��E�:b�����'N$9��h� ��NS&C�l��'�.`Z��NV{r��T�=�
���'���ĄD�@��PhaO��1��t��'5N�!��}?ޔ8�.(@|t��'&��p1��C ERФΙ>x�x(O����NT��R��(�嫃LH) џ�G�$�#B`���!oX9)�䊨�y'�.W��`ßn[��� �y�,�"b�4�T�[5w8QZB.��y�e[��	%F0h֠��fH��y�kЯPy�p�%�(k�MS�ӹ��xb�;J3^�x���f*t�AZ��!��l7���A�X��A��Fհ`!�Z<a���H́�V�$�q��?f!�3DJ.d��T�!o�H��G� m!��V}3�����F�SX�U��^O!���pꆵ���D�)��\����7!�� �D�p�	�ѳǞ D5 r"O���0i��Q�@���x��^����~�@��V;�����/^���(u	>D�4@e�ϻr/����6����T�8D�� ��M�p����7?a�<)7b$D����@�Tf-�5�IG�5�C�"D�D����F$>�s"fY�@	"D�����){}��!!Y9B$�'>D����(��B�}��f6�q(Ej�O����<���~2��5Eq��q�%5!K�D�Ow�<�t A�fܓ4�H�Gl��z�IEn�<����?{7B�����0<D���$�O�<Y�h��BNZ��%*��-�nhڗ�Or�<	��D2=x�`�Ah�o�D�1�e�<I�ʶ!���k��S����W`x���'��|����&8��b4d@.Zx��(O��D�O(�OQ>���	%d�e*4��4�y��B>D�<b��9%[��r��;A��풑�)D� ��/B�d�x��a��5�`	i��%D��@���>f6��
�-�:er''D�(��ٲT��Y�t�_2��h�2D��3�+L�"[��=�.&D�Ȑ��)^`�yrA)r8,`��!'D�\8W��#,���+�ֺ"\�(D���w���20�A@G�b�RD�Ԡ'D���6���(k�=��Bi|9�G$D�d�5�[9>�N!���_p���q''D�36�'��E	��/U��tz�K$D��I�p2m�q�B�5�� �!D�`S7+�!+�Z=��	�+l|"K��<D�(J���CfJBeԪn�P���%D��QHG /��٠��R-Ur�A�#D���Ċ�j���n�pf.D��(��X�-h֬)�Ƈ/�^(�a�+D�샣L����8C2�B�k>HB$#)D��b�dO�Rl�C�낼 ]ԤC`$'D�\���E�g�  ȷ�B38{���6b&D��R"B��g��`[���4�ȓc�$D��X�A�
q�&�����=P.nT��&D�`��H�e�f���E�k[��#D�L
#���D:�$zt+:��4��7D����3[�m�%��w�����8D� C�m������B]��#�+6|O�b�x�7�<�P���6Q�����(8D�H��AN7xm�0���T�Z��|��#$D�@"�>S��;���1\'�`p� .D��p4i��	���v	V�oA�8Z�j*D���c�I v�x�iW��V!H�
fL(D�X���^;
����
�iO �� D�� +N�Sj�}r&(�!a�*�D2D�0�UI�vE�����<cWL"D���p���S^ xIťB�9
(�" �,D� x�ނXO�  � ��o�Ȍy��4D�H+�[9Q���g�^�l����4�6D��bE �	X.�tт��_�.�`5�)D�`��Ͳ� Q��M(�+�&D�dH5�B�;���#��8��ez��%D������$�l�����r���#�6D��Á��G:�<�aJ�B�]�a(D�l�ņ���豶,�6-�Q�;D��!
C�ցCl�<q�pm+�M.D�  �L�#\��x7�<Av��3�!D���i���0X��"-#�:uR
+D�lKtj�:59R��VOڮc N5k�)D�� H�j�3b�H)��(, ��v"O��w�Z0>�©��C%3��b�"O�`abàK����ED�*�ܐ�"O2J4O� X�5�&���왠"O>�0�(�.<�0�TbQ�p]�mct"OW
s3�%�GI�vU�l!BcZc�<#��:�$��H
7HJ�E�`�<��|�l�C&��c6|S�v�<ن��Q����ǵ38`�c.f�<)��^�b�8�t�Ҳ2$���Lz�<�dR�|`&��`�0� :���J�<�E#�.��DH���	��qm�I�<	�)
��!
����X����筃m�<�2�S�D�䛖�t{b܋�(�B�<�S��;~� h�!� 
��w�<�c� =t �g�Ш.WġQc*�q�<9�_,cz�[DƊ�i���"�b�<)�F�1X���7��,�2��"�Z�<�u ѳui`��S덺�J})2��@�<��j6\wBݒ�M�5\�08Q7@y�<e�G�H�����<8�v��0I�<�0LG�8D�1�7�:bج�s�^C�<)\m�L�JP*�$�h���d��s�!��V:�ȘQ��U�5�D1��䊰(�!�ą#N¨��9V���c՜iy!��S`\,ӗ��?f
t���!�L�:M^YH��>������+�!�D������%J�?FUZc.�-.�!�$a�}y�ȍ%"'��±�����'��'�8Pz��;)�����C� ,�'� ��RgO<18�
Ă��ztR�'[��f��:>�����F:��9�'������+�l����i�^���'�xR���,P��t��p3�yy�'�l09���~*"hz��[�h�$��'~(�6�Z�_�*P�"ݼe!������?��)����a�3#�ѩ�o18p�ȓ�2�`��2~�fD� K-s�hi����s�$�7�ޘ*��?�|݇�N�J�"fφ1v.�ᱣ�	�[�^p��mbv�R��Ξ�P���al��ȓH����l��3%����oI���@ 0�h�B�g�(h�чΗe��h�'�b�'�Lh�JI�8�x��e딳Q�BmX�'�|a�� X�r�-^�Ek�Ȩ�'?fL FH��y`�Ƙ)?�\x�'��-4�lC��2�\��/���yro].����ԧ�4���)�y�$��}�d�P!��A44	����?��'{���ɷ,]��3�ɜE�By�����"�Ƙ'��!�K�;:�,=3I��5P���'}�	��I�f�ԭ�fBW$?F���
�'�������g��,�����5j��b�'҆��ǘ<z�j1NΉZ�.���'z��#'�+t���@QF i�����'���D4��r 4bb��'��A"�%Spò=�N_�>0k��xR�B�*Mi�W��r����Í�y���4b*f�h��½b�
V�y�o��!زMcBZ�u�4�ғ��yBLY3-�������eX���SdJ.�y��:e��1QH]f�pR󇘇�yr��2��8��Ħ ���1c���y2��
i�
���֮g/���m˻�y
� D��u�6f�8��)T�H�"O�p���B���vhBX @ �"O�A�]���$��vX�"O40��"��	��P\-@v<i�"O��˼QJ!�u%ѹu:�<[w"O6�����+�$ua�# H6>@	�"O
l �`��w�y�w#��AKm	�"O0|�4IR�g�-Z�  ���LZ�"O��q��Y�I��AS� �8+��m��"O�	Q��Ş���HU���R0S��D-LO&A��u����bdө`@.�rP"O1��	�&/��Ec�v=Pcw"O���ԄɬiZ��'B>F,`r�"O��@�:���Ja�)�"Od4��� `�h �o��^�*�"O�|� c�Zp��E�G�)�"OZE�
�T�h �w�E �^l�#�d�O,����7���AR�)�|AQj˯[�!�d��Y�Z�#ۺФ��g�R��!��[�u��Ex�؜[����ƅEo!�4v]x�xq�
�?�J�I���0#P!�$-�T��Q̑m ^���D̈F�!�бn����BW�%	�d�����y�!�$���*����%9�~�(�V�c�!�$����)��l����'K�!�dN�Mz�a��K�*X����b��G�!�	XEհCk<G��%�� A!�Ĉ�;���2��$t�б��MP�z$!�Ĕ8��K��:A���/dX`�w��<I�<X���(߂8�~Q�7iR,(�9�Iԟ�&��G��'��t�c%��W�\5�Ώ�I x��'��q�&�g�|��s�FxG���'�!�с�s����L�>դU��'_6d�g��P Q�39X$�Q�'�T$˄��)q��ӇS�g�f���'b��B��ҲV��ȶ��M�n��O>�
�w��@���[�;�YI�#�Z]�'��'��>�	�{0A�7!	-�� C�x��B䉢?��j�	ޒ,HjH A�PFqxC�	�H�|p��F�'u��푔�O.WTC�I��B��
�(s�a��'?FC�I�a^1I��1f5�ŀ��JC䉩(���$G'_J�����a�0�OT����+�na�#�ż[�L�zb�!`�r���O|�=	�^.p	��v��Xb����Ȏ��y�E�n��(�$D�U|l�ࡗ$�y�Ó�	?b)��MR�KH\j�j#�y�(��v�t<{��;�)�'돝�y�/3*0T����i�$�
�(�yrٜD!�\��K��+&�+�D���$�O���$=g�T�G!Y![��h�ֱ:�!��ʤL�`C6��4�R���ȋ#�!��R'�9xvFO cH���Ĉo�!�d�"6+ĵ�cܿ���%ߘh�!��L40i�e�˞m�؀�wI�!�dL��M���E�L8K2BH i�C�����(1�
�)����RW��0�'�a~�%�+ ,�UC$Hr�ф��y2��4��D�")��-��pp���y����ppv��ꈲXh�WHL��ybJ��5d$�s�g�<�<sw�P�y2-�n���kL��z�pG�D��y2ၜ#��D��`�	 <k&+@��y��-k����*�������y
� r+�	/o|t�$���m��"Od�*�e�J��hՀ�g#T�G"O��ru�m}5��@�L�q�E"O�u�b吝g&b�I�j��=��[�"O���MCi�4��f�QA��	�"Ov�eb	Zl*\ d%� *� PD"O`lC�P-^p���F�0i��"O��Y*}Z�sEDʾ\�R$yD��~�O����/�O�;�II�\�t��'�pA&[�6���! ��Y� ub�'�,��P�_��Y��GS�X'~�y�'�\��N��!T���P`:�uY�'�N(Uk��G��6Kio�}�'c��o�;�V�v��(R���P
�'���i$M5([��	���-s���؎�$�O<��8�'7�F}z��{)���E%M�c� �ȓO,�s��S#�b��e�
\����4zm��n�}5��Ƀ�W>��ȓD��f��9kn����Dx���ȓu�������.�KC*�h\���ȓH��
�z)���Y�L!�S3D��t�Ԛg�T�9%�0%��e�2|O�b�4�S����H�j�0aÀew 0D��X4�Z�LԒaq�ǈQ*
!zd�-D�XS���:[���3eEJ$:k��>D�4xń[�Y�!�EfZ�^]�q�<D�`ڤI o ) eڲ9� � ��,D�0 �Bo����a
w?�Z��0D�lÒFƗ7$�1�A��u����2D��C�׃)��;�"��c
���-/D�D�#��`���"B�!K�%���-D��X�Aƙ")rQb� F�%��**D��Jv�ȉV|�Ѱ%ɮ:&�|��D(D�L�a
�"V)����"�HƶP	�+�O��3e�Z�Z�.��� +�˺+=�C䉧pN�< �g�/L�T��A�dB��::rY��ί0�,P��/f\B�I�7,�r��|�&Ԩ��ʴbFB䉖_��yD��9I1�}s�ʛ�2B䉾9�LP)��X�U$$��`gʺ\nnC�	:J�!��&��5���Ȧd�C䉜hfZ�0�*3})���@G6F���7����_C�����"�' <z��&�:D�PRq@�&~�3g��n;t�8D�P	Vd�a�z�(�Y�~"Z�6�6D�t���.E�yd �	lz -J0	9D��R@�O
	�:���(7s��E�2D�dyp�Q�A�hxi�KE�@�G�$D��C�,��2,��R�/��	�b� �b$D���-��{�o�/��;�$D�Pcc�������5���$� D����!��|�����`����#D����"}�&�0A< ��Rl-D�8�L�3�����H�-߸���8D�l�"�.#���s�)z�0 :D����"@�Lg��"�
й�de�6�9D��f
ր%�$V�m�8őW�9D���֊9i�)P��^� ��!'6D���#�P�/�]@+�II���1D�d���Łtz�!�� \��	EN4D�$@�&�4+�L�R4 �3,����(D���玝:.���p�_PB��Q7�9D��ڶ�(8���/��RV��3Q�9D��z���|H�L2�[q@��t#D�� 25�'��7&��8Rn�'6���"OjA۠��$_ΐ�\)/V��"On�Ӵn�,$ݢ(y L]-{�i��"OQb&��
��p
�kۨb��aА"O��"4Ŏ?F��̐��!Y��P"O�)�h���$���DO;=��8pc"OhX8e�Ƕ��P��[�~��"O�U�� `h�%+z�ƴ[�"O�ŨGL,/h�J�'��'�V�kb"O5���P*�����7�p("O"��IHb�V���L
|�p�Е"O�|u$�?[X\�Å���2:�z$"O6�JA�P0d��E�/�!j�"O�p��3������e�t"O"�R##d�yj6�V�Q;�"OXIy2�G�
���@�
�vP$iY�"O��#7`�.Pg�H˃��g��"OP���,�`A��U�F�D�nP�"O���] 1�V�	B�L��]�"O�#a�N�h���1���ģ�*Op���&	�N��E��U=Y�*���'�mx��/<�(��`�db����'��YCn=������-j���	�'�K�C1X@Q��i�V!y��M�<�6��I�d�j��	�zlب  ��J�<)�˔8E���J�JH�8&�B[�<Q ��0,N��6D
2�b�a���S�<�f�[���ha*�-DD� h ��W�<IUL�%S�!k#��8H>0TcX�<����mR����X����%�y�<q�ҌK�65BuGI�DHp��b�l�<�6�S/0�W)XO�jR��^g�<�Y�<�NE��aI���y��d�<჋Q�\����&�725�!m�t�<i�I�O�n�hC_0 ����ǁh�<٧l�4Yy���k�"{f��8d)�K�<I�/�
Jh( Wǟ�{0���FG�<�s+[$`�� ��L��"�+�I\�<��nV�N�$X�̩��:�D\z�<YB��]c�a���ql�5`��Ly�<�ՏֳR�4�5�Ѝy��(E��w�<)�f 3o�R��t��! qAOK�<�%G<Q�HB ��
���E�A�<i6l�	{P��JO�U00Y���B�<y��$���ˠ�?R��R� �|�<Y�e]�?��4�R��H�µ+&-N�<���H���]!�p�0�,@@�<��P;0��XzdÚh�|8��y�<�%� �.+���<W����z�<ydC2_2��ō�B�H�[pN�z�<b畊���[D&�$o<���z�<A�QCL��b���D�9��u�<��N5]����^�Cv�yyg�As�<a��@�@i���$�� �͇n�<���\�Be��ˠ��5-;4tH�ğD�<�g+I?U8�X�U�3S��p`a@W�<��B^B�6��E��
�4\Ȧ��U�<a`�	cF��KeCMZA~�P��y�<	��B�q�Uc#�˗(?č�4Kv�<1GbS&>� ������f�s�<���(��5�tC�$�6�j���l�<!�����Rt�_�XQNQ�@.�S�<�W�84��cQ Ƭa$eBN�<�E��D�����L�?�ћb�I�<� ���-/$�
�JxF�8"O��F���4�{ɞPDށ��"O��q�7��(���%^D�Hb"O|]�3m�`TD ���Կ yli�"O������ɰ=3!J�inp�@3"O���Bֺ_��T���o\��"O8�qU��?;h��Pb�� ?�a3�"ON���ڌ5�4Kbd̿2��:�"O�Q*��8��ط"����Z�"O6��g*�K��0�G��̱��*Ol-��C? I��SR���j��Ր	�'Ӹ�Q쑖2�T� oaҲxZ
�'�%��6�&i@�)�U����	�'&�1k0�
	 �X��T/K�\��t��'��N^&,�$0y�F9V���#�'�!������	��H�V,H�'�Z���
�;���5*L
��Ț�'�]:� �7,��Ta#��|z�dY�'2�������N0m�X3�'�\%��Ţ$�}����ihz��'P��M�m�l�c�B�3�ొ	�',^�h�j�|�l�$�@�m!��x	�'Њ�!�j�<��}+�C�W��H	�'`V�3��V%�U� L]A
�'����G�Z�@_`��W�G<Nw�Pi
�'����W��	,j���Xhxs	�'���/e���kb�] '��H�<�A��/Mu
i@�:IN� ��B�<���ֆC�>8�(�JS�}�O�C�<QQ��94�8x�V&�ep5�� ~�<qp�����yg�֘\���KIy�<�nID� IfN�z�Vu�Ĭ�u�<���I� ��O��U����\g�<)�P��e�%� �ε`f��f�<��dމ:hN��6ńN�~�J��v�<)�ME.QT��s�E[�\%j1cr�_I�<��˙ 6d���
��i�ШH�<I��A�2�Tx�d_4}Z�ڣ._{�<���ܚ|�%���P,0� F
�p�<Q�`�4B>X�Q0�׊	`��q�<���?�@"w/
7��3��y�<iB��i�M����o/!jB�	����#�nG8zx1��	��B䉨~A��Y��>&4�{���;yŪC�	�IOxI(��z�pe��c�Y�JB�	�{��[�mU RªX �N�>�bC�ɞff���ʥZ~`�B� �LC��,���HW$ߺv�^�W)�;k"�C�	�Fi@$!���%�`��'����C�	�]�ݡ'�^�V7B��C	 5K�C�I�7��u� �kiR��@K\;�LB�ɍA� 5!����#�lp(��ܐ^�*B䉝*�p1�Lɱf�xP:G��nTB��%r�
�)�B6tȤ!:�o�"�C�I��&p�eםIh^`�f	�-k~B�lK����7�P�d��:q0C�#r�n�#�K�8t��K�67�$C�I&8ڼ�A ǅ�:�<A�]�<�4B䉐z����խat,�K�"���FB�I$~��A*��U>l�8��É]@jB�I64]"��5-���:��فs�HB�	)n���٢�N�#`�(Z3��UdB�;<��9puH�L���aԆ>�C�ɦ)����o�su�\r1�Щl5�C�)� �1��.����"�#��x��"O$��r+W�r�ʭ��.�� 
�"O�ԛVfY8>�l��k��Ic"Or�[��ؗ��
@ƒ�*�D�8�"O�W'B�
��X���E0��0Ig"O�(K0hH�fЪ-BF�
7�8e��"O�j���q���zhu�"O"](�I/u2H5�e�Y�7W"\ۦ"OXE���!�ZLZ�F��(Pr�q�"O����\8]�rlH��P�?$��'"Od��C��.o@H����hh�(R"Ov0��,�-*m���O�b�i�v"O�����.Z���'�Y�a�N�Qf"O�8�N��#�����%��Q1"O�5�AaЄ;�j�8�@ʻ47a!"Opt u,�%9�z����&��!��"O�y�#���gތ�`N1Q�����"O␹��grdr-�4�H�:"O^���%Ғ/�8p��ڥk��9�"O�x�O���P�	�1=���!"Op%@a&I�]����I�I�X]
�"O|�h�呍��� �;��#7"OVD
P� @��S�yp� "O�!�M#c��� n\�(̕�"Ob�ӏ���^Y�vg�~|{�"O6���A�iB �sa%T!1� {a"O�5� ��)9�|��⚃�2dI�"OJ�Qq�y�@���7z�l��"O^�T슋�,��j��j���qa"O��r�Ĳ3-,j�iS�X�6M�v"O�t·,]�e�֠�'\�J�8U�C"O�#�+�!��@�䑖	��5�'&��M�#7� �c@p=H�B�'[��s�g˶C�֝ ��C�ra�'���C6�Ql�k��Y�~e���'�z��oL�-���σ�r�r(�'DĘr�AL<F>J�KGΑi�����'f�U�P�u4&��vk[
h\ ��'Hp��KN��hmK5䂏s��Ux�'��t�����u���d1��
�'�A@�9��զΤc;�m��'�@=��MHE��Բ����G����'�z�����y�&e��e�K�0��	�'�(�d�$��B�@C�<��'�4X��F�g�`iH>�H-��'�������}k�3~�T�*
�'6^��P�{�8�`�Y(���	�'cBz3m�4R^XD9%ʑ�s&�|��'�����*_LE5¤b�9q`����'_�=��Ř>
��3�F����|��'޼�a�Ŗ�l��m��j�A��<@�'��] ���(Q	�ə&P� ��')�x"�Įyu�h��O�I%�lr�'A�DX�A#CT�$.|�æB���y��x00��1�ͱn�ș7#�8�yb�Qu`4	 ��F ����F��;�yR�*Rr%A�+
:�t*F�կ�y"�Wgy
��vL�b�b�N׹�y��*����RFHol�X��K��y��-A����n�P`hM��yB��oźMA��&n���v�5�y�웆/=�2�X�1��&�yr"�|�0`�G�7���+��yRa<D�j�!�l�d�)gd���y
� �@�t��mm����ՓF�\��c"O�-�!�ů^��
5k�7�NI��"OaxaH��.l�A��2[��a7D� ��M�{��3M ���&�"D�� 5��v�R����?ܔ�P�5D�P�⤛ ���Ɂ�'i�{�d7D�p@7Ã�c��dB�l+�pPS�4D�����8��0��(�p�HС6D���0'D(1����PN�,�`(��6D�����W�ֈ��E�ҙc��@���'D�x�Ϣx~ƍђ��h��Taw D�ؓEH��o��Y��Q'I���`�=D��k�ȑ6+�dՁϣZd��7G<D�4���I	{B�K#�I�~U@�Y�
:D�8��_&=�4*(�� >�hRAm=D���gA�4R��*��=I��;��<D��ڰ���Ex0hB�p|� c��/D�c������Љ^J7��"A'.D�T�!�֞�$-����m� 
2�*D�KY\(��2�5h����*D���L�:����	6*�z��B�'D�|�V�ߦ�8a3�fƖD168�V�2D�|"p�$R�(�p����L��1���0D� B���Xb��$�����i-D��\�1�D�*ÐM�sCJ��hC��(���Qd�X?-�x����*q2C�IZm���L��S�tRѠ׶1fB�	?l�H|�`bV+:$��B�/�UDB�Z,@dq�H�?�¥�F�^8&�:B�	�P��A�-�C��l�A�x�$B䉫(��3��y9�R���22B䉈X;�y9�ȻM~D���3u�C�	0;H2ك�LS	1o4�T�4�C䉮�a�i-}��$@��ئ�C䉯IS�lQBM W1��y3(��;����+�	��~h�+އj�V���)K��vC䉅.~8��ى-L���̬8fB�O�������O�HcH
-��ƌ���mӍ{rH�Q��d��%(^��xe�#He�e�4�0<�۴�BQ���¢VqpB®� L��Ն�V��p2��LI�4P�,вE��͆�m-�h���Y�Z	`�*�$��P��I�<�4)F x��|a x=*�b��]�<9Ƈ�5O��z�Ś�Dʀ<�d�X�'���E���c�H0Ғys���?6��h�ȓA�&MÅ��(o�s��\p��_����sI�+�ѭ�"�|�����r�̖�e�EМ[��ȓG���e�ՓiL�(��s�ĉ����<al�<B��5@dC	 g�:�Z�w��z����`%�'�a�\{Q�Td��d3"O��s�bq��5�'g[Vr���E"O
 �v\�(~��˶,�6"]j�!"OPu���Mn&MⰉȩ	V�h��"O!�jʈ|x	�r��6W��C�'|��'Kt���N�fl��DR�s�b`�	�'�,9��aӢ��9��Y�hd�`H�'=�a�s�:�i��Y�@��'�~}��D5f�xl郠��{Mt�9�'5��tnD�Bo`�#�Ѣ(HLp��'h���3�W9��s�� F�ى�'���)F(ԞE`�I�sG�2��
����9~���6�<)�!�ϩ}O!�䇹0�-�5㌫��yBA�=0�(���D�<� �#�&M�B�@���,
�D���"O�p�
L+5VT�!0�B&n�v� �#�K��DEb�v�]I�	�RЉ�D�(O^c���=�r@Q7�l�ѷ��8��סV��C��)[��Ų�!��@m��)�Cs��:Ǔg�x�ڎyr'�8��zw�G�H���%��yb��0��u*G�K�9��! W�����?ь�����(!�D��$�*�!����y�[!/����P�,2P}
��Y��y�h��h��Λ8�F�Xw�"�p=��}��/���#�L7lB̉����y�ϱs,�SA��$+p��eI��yR�;'�A�琥g2�p�Ý�y�$����ic!�Ev`a:�F
*�yR�s+��-��^+<��90��P�y2O3 ��s ��/��El��yr+J[���7J&7�iB",�%��<-�Mۋ{�.U(b�`�K͌�U8402�P4�yR
�+K!�� �HG�R74�:����'
�{�N�>���SA���ؓR��y�Ѡ~�DYK�'��a�7a���O�O�?P�ϔ�ȡh (G5,��Q[�'�O��'��t���ԙv	*1�3�� �*��$!O��Ƞm^�y�9��lՠC�B����r���)I�V��Y"��1F��L�/0dʎ�$)�	_y�fZ�k��i��(�0|1���B���'Vў� 8�G�&+N�+qO�=�ΐ �'�1O:H��䒄��@5� l>Hmʦ"Ofr"�N<s`��k��D*2)�g"O��ѓ(�c���c�4���\�D{��		�u�����[	W2���`�9d!�Ć?���H�!Y	?��o�v!���MH(��V$48H;Ck�s�b�)�&�<��3�Ǔ�p`�H2��	�'�� z�D��_�4Q@7��F�,�,O����2(FlZ�)����LوO�!�$ƉB�v���F\�}�*]q�L� #|!�$^'U�(A3��QA`�lS�Ҧjў̄�Ӊy�P}Q+^�(�
���Ur���$z��soS�EE����j�;-��\�'�Or@�'����ı�Ns�`հK��=����)�/��)Ӡ&R嚥Q7�m�X�FzR�?��%�S3����+�<*��E� 8��C�	�q���ʅC�:�Hi�k��/k���hO�>�ce,��	����`��4\��E�%?ً�ᓟ!XZ��"K�+�d�����HO67�7lO8��Ɓ�O��k˯b�h�#���&lOL��+;z$RD�G�Pn�8�,D�<B@�E�P�b��H�z1@`��.?D��e�ݺI]*sa�%N" �P��=D��6H��(Y/��i񈁆S}�C�I0�@�+"'ݶg�B�o�52������O����RX��c�ڮ&�M��"O$���c��l����VW�B��8ˆ"O��c`k�3~����].7�Di�G"O�E��i\n0��JRdG��{"O`��Q�V�m3i�96;6��"O��s���x����莝�	�P�d'�L��2[���
���(��q�)\;B' B�I��`��J { ��PQ	�ތ6��N<�v����Go�J<�a�K	�*�=I<i��De�\���8����k#�p ���yBȍx|��i�L�i�ȸ`����y��)�<�jd�ƂT��c%�?�fM�<qߴ�O1�� p�"���`�ƈ*7-��W����1O�7�r����f�^勒��*�t9�E� ������4�����,R��G��,�ލ��(Z܋�'�^�P� ^"!@�Ao�T���'���P��8�i(*nP Jg��zM�I�7�-�O@O��" �Q�`�}k���,�0JU5Of���RJ kQJT�WV:��GCL!�A.c�e���	5/\��9%'�M1!�D>V�ʉ�7JH�6��=�t,��!�!��ܝ �q0�,,J����C��!��>�IAbKH�y�����#J�!�N�>m��RE����.�y1\��!�_,:�:���H���Kd���kB!�$�*$]���@ؠUA�ޙ:&!�D��^��Y�dD�/�B	��g�!�DXq�)Æ��W�H��W*�d�!�D;h�ڈ:�m��F��y�7�
��!�
K7tu�U��(s��h���B��'oQ�\�?����*&�nԊD��y��gF�v؟4���JT@�I'����ʲs}֜�ȓX��*�C�P�&�A$ٯ{��t���x��>���%� ( F�[�-�ȓ��8u�ϲ-E܀"��Z#R���t�Xa���'Hr��0[hx�ȓ�v�хU�%Z���E�D*_8�ȓ9;��"�ӁQ`Z�Q"͋�]�(m�ȓ�r�!�_:k�Ԉ��Nަr^V���P� u����?�(�QM�>w���1�4�`4��*���0G���v2���$3�M�C?WF���eر6'*���u�teS�\�'ZV`�l*`�t\�ȓ+�B�)vo�2plipD�X
jpꀇ�*7aao;�r�{#GԇXĔ)�ȓ]�� ��#�64�)y$�;5d���ec�ـ��w��$�4f;d�� �ȓ4���g�\�z���K $�(i��L��Eu�f�,+F�ɘKw"d�ȓSG���#I%!zxr�E�1�6�ȓQ��!Y��+i8���m�<�6ȅȓ�LI���K�� G������� ���牋#�T`)��
����c���1F��B�p�*�k̑^~�)�ȓQ���pg�-�����
��U��YMĠ�Tb��6� �$I�����G�6�C *�"�p�"§��;ւ���jk�A�&���~l5���1`��E���TMC�	���Ѩ�)L�ń�Y�R%K���D����0����F����"Ֆ�I�d�ҫ	-�9�ȓ����G��iܵ�q-�>(�<0����u�0CC�M�JT�2	V;*�r��RD!���'��M�R+Z8T(d��.%��ZԢ�*h����4'(6,�ȓa���dkUg�3�L�r���Ia� PER2�pͱ4.7x�H8���Jy�� �t	�#��|ָ(��TI�� �撕R/��`���59�0Ԅȓo|0���	-�E��ױ8T�i��~�`M%�4vr��P�F�1��TB���D�^/pC�����i�����d1��+��(,ẍ�2���V�ȓ,؁c'��t�6��TBZ�e��C��M"G���zNCvH����ȓݾq��GF�"�ԥ���F��@ ��S�? �i�k��1
lP�dǨ!��x�"O��B&E�_�
Q���f^�R5"O\�C��ϝ(��ӶD��xU�qP"O0Ab�I�9s����Ĕ6	T`�
c>OʤK��Q:
ARU���(7�.}6�wzt�� ��3[QZep��`]�C�Ʌ/���2/=M�T
�VP64��'��|af�ü3���N��H���'�0���i�i��s��L�OGt���'t����ЖR!:9�e�/*RndH�'q���4�Kq>�)sE��'��<"�'F�����&2H�EA���F�I�'u<x��ۗcLIJeLA�{�Q��'вm��ʺɶ���F�,�(��ʓ{(P���g38��q�NUl���m�v�1�C�>pl�qa��5m���ȓ 1��bo�����Ȝz��ȓ8RtD	�oM.��xH5E�jb4��I.d�If
��:�J)H&OoF0���2�b��&%-�C��J
n����.�6dh���8i�"�۳(�\-b=��$@�%8$%˕f4�����nj�9�������P85����V�0*�&��ȓ%e>�&m.R��5k�(kP�����*�yw�_6`5�	�f,�&)�.`�ȓ;��� � ��"uSoP�2��l��Etjdг��20e,����(����h���l�9��9S�` 1%��M��H�)�dE��p���c갇�>��Ax�+��6�����_�ȓ?M�pi���R�LbBmH��ȓj44���#j�����ؖ{�5�ȓW_��Cu� :J�D�e!�H�Ny�ȓ;�L�r
˶����"R�8��مȓ@����b��9e�A�P�J;S�Z�ȓZ"p�ҦJ<G�L��al,~�E�ȓـ�e���G�Ab�̲c�8х�[��B�� 
��M�U��.	�݅ȓ:����ɢH��Q/^/Xv���J�ͻu�W�(�:��Q�&�;��
���=�A�Ȱ9�ȣ�4U���1	�$%����	��L�,��	K�*5�%�DZ/̼�;'m�q�Ԙ�Έ'a;��d��5>[�i�g��8����׆��/#�����V�+��@XR$IW+!�)�'-dx��I-|�� �׃Y*L��x�FWB�����iL`y���E.�f��cO\)E���؁ �I�F������'����$clmRL�n�0ܐ���N6J��vfD�X���D��]B�oژ*^�8�s"3!^��H�'!����D���=dgr�U���J�l��QP��q�GR��0<A&���g����qAM�(Q�����42:�� ��wf�0�#b�#V�LG�TO�5a��0m��G�)k�m���I��,��?�z�Q�X�z舤���s �c�b�6IU�)��M� 1�'��>���}����K����@�ϛ�/��C�ɉ<T���楕9?��ⳏ
�,���dډjVN��#��*=����$	~%�ò#ؕCj(h{��F	`��{��·$^d�8��I $�E��� Qj�2�� ��M{�"O��֌��M�L��b�<K4��B�Ɇ4Zb�U$�Q>�0�������!�%�*D?\�KW�8D��B��U�`�2 �RD&~4o۪$�nXH�IF���S��?Qw��FQ�"c�ۣ=��{V�_�<!�F�._��d�N~��Հ��_�<��N��X,P�h���auB��]�<�!$l������0`%�_�<A�i�G�L!i�6=6��cŀT�<i0�N�a4��C�kA3o�F����V�<i�
�"* 80"
֯M?�M�d`WZ�<� $�pB ���ƨɞ|�bM�1"O������HH�p�Gg��yD2��'��X���Nx��'h��z���23������ЂC�I��Hx3E��*O�ȋrL\�]V��'W�ĩgX9(�ɧ�O�@Ph��<b���3dؤ`)��*
�'C$��C�^��ä��*y���B�BY��	�_�������|B]�2܅Vg0)E];  !��ŵyI�L�vԯC@|4��G[%h3Nx��&llT�"�Vvz���@>#pʠ1��ÏD�2�ቕ�5���L�^�;z���^��5ʢ�"��x�ȓp���FC1*oa��d��3c��'P����	� l�ܧO>�J�Hߗg;z�a�	����z(�O��Z���HѲ`�ħت+v�Q�����m�6���N�{�P�4�e7�ln�:_l�y! �5w�JD�� 4�[����LK�+}����'���R��dw𰋢k�'?������M�mp��{�����Үn��l�"��^��4JT���p���^��J&g�K����<<���3�����$Zā"���i&Y��A^q�� \h<��ˎv�,`c'|Z�M�'��<|�����4œ⎋�.����;m���S<(����*�)92���Ό���<W�y�f�)�O��BdɃ,�x���+zp��҇$�<����+m��e�' -zvharM�J�`��&�]��)I���$��-��iP�'�q;��S�c	-j�Q�P��h��bp��hw��8��">mD��W�,Vx�}:!m�$H�Fz���B��X���E��� <k����ŋ́ɬz&e��W(�ɮ��`M�0/��"�Y�Mt��BȰ|�2JĂa`<ѹ��� R����Ep��[�/�2$i0`�SIa�C0g�s�Ҥw��J$�ڵ"5�c�'�.u��L֣Ү!�3�ĉp��=�p���Ӽ[uɨx}�A�*P6.jr<:�oCw���ˀ��'��dAw˝��0L  �ՠXv��A�K��r��%���F=�5g�1��xyݲ��gi������)�8�!Clϩ+s ">Q��0rx���p%S�<f��a񔉳�_,J�3W�� ε�ϙ:>���R�$�1r��0Y�])��#?�UhP�~R�3f�:.~��+s��Φ	5��*!|�$@�O6zg��?�c�A�-y����Y�
�ڴ�$h,c�@	�
�(H��CN��\�P�'Y����1,L�u���\�W�VaY�'�mA�SV�*�B�K�?I�A��&�8]`5.�F��ӮU�R,spb�4�V�g��6$.��_�b���W�r-:�0hͩ5(>�� ۯV���"e�S� ��$D(�z��l�)z�V�~�'�8ͩ�"�~�i@�ܙC��u*��S�L�Q��)D�0�����]܁	Jƴx���3.լ�y2o�(*1���5y�8[��م1񞝚�!�N�*|�g�3�?���O��@r_��m��N�#C�d�Q"O����iN�FUCQ��,�rQ1��'���!�Mշ��	�R�W�"�ax⢄�ay"ք'eX�	��7��=Aa&Ŝd�XD5��e/j!@!�C�"��I30�3!>�ȃ��xҪJ�`��E8�ƀ�5�D�����'@|(@ �TtΖ����̀NiB�(�?��&���SQضO�4� q$6D��A��H�~�2�wEȁस!D%�g����g��u]� �0�
�AS�Q�����O���+wuvx�%f�/%k�`rO���az�eW6P8�O޵Be䕵, ���
E����˜�QORI����L�F�xQ��O��t��t�'E��E���-R��Zҕ��1�	�PĽ���P_ܵ�F�Г-LzQXӠ��]|��o��������Q�7vq�����>�q�U犅9�Z.�Z�B�-@0V㞸�怏����x'�̠i��T�d�T�o
���LBp��dc	:b\�@q#h��	�B䉪��ƫ]�d�򴐵oB�!x��R��Ϙ`�ԩ{F��X�.� �ǉ*���9��)�O&�3 ր�:�3�M��!cG�'҅�V��F�DO�{��Y�	�6_�r�H��Р_;��Ή�$�X|�厇�&�	��ӟў��.��p	��&�x5PJt�L���';.5"B�$G�EE�81�ㇸ!A�T�a�B�hAD*k��-� O������;}�Ѕ�5HQ�L�N@��us�z��O��������6��hr�%ߌJĝ3th�y��!ln�-hB
7�dq���'��k��R�B�?E�2�@�d9SB K���p��/D�4h��|]ʼ�5�7)ΐ�XC��E�"p���{���c����G�G}��F�oE[b˔�=P�{BdA�$�H�'Cp�:�+��-�|IxB�ӗ[��l��4Y�z��-��	ߓ�<���!�,oxu�ʈ�����>9�(F1nm:P�,O|aҲJ��ʼ���'|f��AM�>;�ȭӄ�T����S�? �0H��� �r'L�efDA��-�w�)P�$Sj��ic�{��)��yW"����|���2Zn4h���yr���TS�`�0��V��tc�H 
�XxuL	���q�OT��fBʫ-j$\؏��Վ:\�]��g�@��-�B�E�p=����kǸ�IA�|��P�[�0�L��%���EX�Xv�}��i����t�E"�h��`��ꄶ
]<��ڈlvd��=a��4=��h�WE�>)��i$����'��`ЈDL�V���&��2<��8"O�,9�g��~�h%�@��@t�0�ϑUr���gZ�0��Ì$9OJ��}�1�r�ݢ�DM�`�,�&J��I��0D�|2���*�P����5����sO�'s�t��bMD���O�:����:�+B�щ��8Z�����S� >���I9y�h�¤���D���崝��*		�����O�B�!�$C�<�0(�ڭ+��,RF����O��bt���7�~� ���$� 5J�E�53�֜�JSi�<A���D	!��6H�pX�tE�=%�����>�g?�wa��ڼ����X��������~�<Ip!��.0�Rn�2&���h�q�<�c�o�!H�! -`6���s�<	%J�7C��s���*l}H�o�<��'��zǌ]o���ca�Gk�<!EG�$fI� ��>s��u�d�<�qăgyb�w��# _j���
�g�<abP��@0K��@����aIf�<a�D�O	J��@M�f@����a�<��G!W0�mI�G�2=Xs�"�a�<)E��GO��Q��& �\�ӥ�J�<9PE�0�-��a��eU*`e�D�<A��2UlC ��>nR��6HMF�<	�f� վ��/�CФiȰj A�<9dAC�2��k�X'v�Xe*a�<�פ�
�x���ŗ�,��&�\�<���='n���Ck�[���K1cB�<Y�ݥ]4�TR�悳O$���-DW�<Ƀ��̂A�P��j����a�N�<�E�[�M ƈ�q��+O�d��K�p�<i�c� ]��1�����L���`�<	p)2�x��ĎT*w@�d�1 a�<I1Ԃt��5+�S hp�Lc�<��`7"��1��s7j|ib�w�<٦�̥hH>���Ƙ3c��Hs�Ck�<1�(R�7��X�u�I�*���Цf�<�%N1_�Eb�bZ�7�t��"Lb�<9�(�ye~��B�).`�����A�<�lHX�6�`��$%���)�Y�<��,��� ��&!m��i�ag	m�<Q"i��u� �_�BY��Q�<)cIU"\#ÌQn�V�"Q��i�<Q�@(nb�s��g�����i�<RAN�~���`׭/�v)j��b�<)�\�m��A�c �,��(�T
�Q�<���5�ܩ�&ű��qf�L�<	�(m	�M7AѲz�jPI�C�<A2��z��Z�%R8�j�g�{�<��f#����&Ù$G�qr��B|�<q��ܬ;�N-B�,�/P��f�u�<�$��"���6�(}E8Ґ��u�<y���
;��):��jEt�E�X�<9u���:Z�jq��g0L!3  ^T�<q�
��q����3�_6:T�rw�R�<�b"X	JbIڵ����@O�<I� H�B��X���=3�~��GK�<q�L1	�1iS
<!X�8gIF�<�q��<Q\�YU3
e&� f#H�<	���a���t����.�Ȁ���<� ��ۥc6�fh�V�W�R,P�Ȑ"O�4�ƂS8\s^幤F8ޡ�"OV�@Ɇ)�X���%E�w�f81!"OR�)$&�&XE�}y�D���\a��"Ox�b5K�
��di�M�^��B"O]�s.	Ptʲ�E�M�"O�ɸ��@^���/��-&~���"OP��`ކl�r��g�^�A��(�"O�d�F��9�-�r�9rR�Y�"O����I�[~1zc�SnD^���"O$h�wƭ�,H�i,�+"O���Ǳi����T
otx 0"O����+*�E�e�F�,V��@"O	�v�4����$K�ac�+r"O�1�4��5c�&� *JLH�	R"O �!�F�/.ȱ�
�)?nik�"O����a�k��hfˆf�B��"O$Xq��A0W_��/�9��"O=� ����ӗH�\��i�S"O]K��C��H	��W�J��"OJyS��<��Q�v��`Fb�)b"O�I��E�%�ػD'�7;�ɂ"O��R�FJ.G�\ȑG&�24!� K�"O"��/a���	7&�mVi�"OB�7����.m!�ϋ�t?���*O�݂��F�����V�2"LZ�'��	(U�)\�Z�;v-R�|��D��'T��EʹU�J}B���\�Z�'�,��5�ɻ1��"D���N�8�'�J�hS%� `���˘�s�"y1�'����e�Q$`�c�l��h�Ht��'&��kv@R�|{��ٗJVgȠ̅�/G�Xy�JźK�Ȍk` �~r�H�ȓct�U��&��F��*���ȓ��s�B��4S��*����4����Nf��1N��B�` �ȓ����qe��@�;���HY&��FbU�עK�r
�#t	(qq�Ą�VHKEgT��63dɞ)Jn�Q�ȓywE�3�	=t���U!�?���c9�X��N�Ȫ C��J׆̅ȓ�&l��MV�S���z�.О3�ځ��2��T��G[|���+�����I
AU�H�������s������������$D�(i� �a�"�*'���SD/<���{�DIB<ʣ|:e�ׯt�.<��=l�ɸ� K{�<y���iǪL�eLO G�]�����f��|�L
5Y�� �����Dڕg�舥*˞M�|�2�� �!�DJ�pmbTXd,�&r�|�k�l4�ƄA̶Ar�@��az���@�@�`�N�T��Ɨ#��=�t���Lfd	�A	�A��j'kPG� b���8T7NE��'��rf
�> ��e��l��T�N���j&�"|�%�էB>��PhЉ���
d�Z�4���3D��b�݈QH��q�Z�"��{ׅڡ)<Ľ(�?���h��Ě;@h��w���)7����8�!�DL� ���y%'0&	ڰA�T�b^���Sx&(32��V�azrFȩ���g�p�j�J���8��=W�)�V���H).�h��)��;˺Q�	@�l.P�	�'��ibO���i�!�n��P{��h
�������(�� xqK����(t�E4��J�"O��r�Կ&��!��	T�ū �[-&BH�{r�_r�)�矸k�"��:��k�n�����r�>D��S�m /�;�N�;]!�)��?D��e�JL8Bd�N����6�:D�� ܉2��P�^��H�
U�:��]�0"OP�k�e�$�PQy��׈H�`��"O�|"e�˻?Hʀ���V���8#"O�LFeV9�`��.ًG�$Y��"O���bǒ	vQ`p@A�O1/И{"OF��CƲ��Ђ�̃8��Ç�WX�����f�'ԑˇ��7Ũ)pVϝ�Vl��a�'@8����zP0�@c�1@^\�!O��H�a�`���$��?�dݢ�����NA��)��N:D�x�GAQ���FŞZָ�p�E�{���Y�AHI�g�O�r�+S@��!��;�'�7H����N�f�s������K3��,5$��w�� �pM:1.�O�m���ܤ&ʊ��`+C�@1��i�'�()��\|�O��)@���+%neK���*3���9�"O,�J������$�BD�7Y�n|���Lq4eIl������>E��˔�'\lZ4�%A���f$���?i����ŲC�9/Ӝ�5�͆g��q��,:&��xi"�%̚*`�f�>� ?[	2 '@�3Ch��n�'8��b��ٹ?�	��O<8�̗H(��Kӭ!4g��{�K�\��h���^��p?yw�R�	�4�ǘ��d�妊g?��A�;�����K�5W>�	<,	`�)fe&7X��\�S�,8�$C��I�2M��gY�2����w���x�*�-q�d�	���5�Z����͉�.��'����T�͖)`R�p��~0�) H�L'�x�R�Eϼ�7-�(I�2�D�<�q3�&PJ���!��޷B(Q`�o�"}.��f��)�j��A&��1�ׂ[�ia"-�r���c<a A/Y�,哴[���)w\���g���9F�F2��>�"'�8�T�f
J`�h�'Ύd��o�Z\��E|�9�lH4%J|I����5�@�􀖚@ʂ"?6O�v1�q�0*u���K?��Ȁ�%4���)ڝ}Zʧ5����'mx<�iQ�4�M�.��
	i½i���� �X���d�5 �$*1�E���\��,�/w��Uq#�O^��F�7g�p���.�~�xb�Sk�U����y�.F2y�:E�6�^�Liǭ��p?�d:��Y"È�r���z�PeD�39��qz��q���Y7)�SL�9��O�1��%	�I�|����>q5�$"�j�	0�O��j]�U��u�'�$�KL#zP8F�?Ij���!r,�YvK���jq���5rg�Мg��@�\�͜�H���RX��e'R18��@%�W0V�@�H��02C,_�Z�O�b���?	$�D�v`����`��"@f�U�`)x����9�����]�$���l�VTP7M�7�1OT\pg��5���dB1}%��J%��пP���S��Q)�@�k�AāZ�!����AAq%I�\8�1� O	ou
y���O����Y� xHp���Y� �4�ݩ3��q��hX���aC�*D�ț�K��j������i�1�	+D��S*����bR}�言� ?D�����5,���! �As�`+�M!D��3�&]�^p[���1,~�}[�'>D�(�G WL�0�%=��2d*<D�X���
&"<@�DH��e��E�Uf:D�8 ��J�cf ��a@Z>U�����%D�hAB�h�TA"�BU�z��e9b�7D�P���ǆ^�^�W�V�<���y��4D���c�ݙK2���gH8�l�Vb)D��x��E aG6�[�F� 5z`�¡�8D�� )�ZZ,�(t��v�Fp�bH4D��;��i�@���?�Z,��%5D��te�X�q�
;I	!��6D�,:`I�0�dpH@i��MhƠ�1�;D��Z�vi�ؑ��A3;� СG3D�h)C�˘�Aj��	Wu��q��%D��1S%�>#��\Eŭ͢а�C"D��C-�<�FԢN+��k֯ D�h�.)3]h,`P,V�l���6�$D�@3���Y������DH&��� #�O�,R)�,�~�F1*3���Cȭ;�&�ô�9�y�E#{hp��h�0����p���'��N�G?����L�*�<���'٢Ԕ��:D�L��eA.W��,QR+VO%������LZ�Be��R�$�d���� 5z��
a1H�* !��F:h�`&�'f�{��M}��VV}���"#��x&�=(ad�
�M[�jO3Up��T�$|O�xpu`�Ta�m�s/�6;� ���NjB4���<�#�4=�)�D럜� ��S+m\�|`�Aǯքҥ"O^�!��_x�l�b������!E�&�W�  �L&#��8v�M��y������Λ�{�t ���%�y�N���I����Aw�P��F�'(��iPJڗi�F��O8UQ�M�TذX;��.�R5�1J1:�D9ueH��p=�l W�^u!�d��FX�h�� P I�~$F�0"�����0��0��L 4dT-:�P�#OD% ��=-O����H86�I}蕐���Ba��&��Nj��V`�'hX:��D$;�y���(H�$�ӆf�+Ƃ�J�H�0jS¸�$��>���"r¬qI*2��c��n
�Rk���d1�0̀�R!�dN�7��SE���z�Dtr5IзL��1C�P������7"8}�Q���F$�!gqJ�c��3�"�Rw�7\OZ4ڧ��4�ޕ�'5���kQ �xǩ�3o����'z�r5�� "������:QRaP�}��CV^a����PUb��T�D�K�₦}xC�I&q�P��4E��|� -RD�X��lJ�.͸'^�>��>@^틡ኩ���2d�Bf2B�	�YĨ��̒y��B.H�jx(B�	�3� �{D��3�����D#�C䉣J`L�h���j����G��`[B���I`�IK�+sB�z��)+�C�ɪb���+���0 ��mPrM̉&�jC�	�'򹈶O�1܊�Qn�ɰC��)G��ô�ր/vuH-{vNB�9&ؑr'˂t la��ŉ�$B�ɻB�v!�$#��v�E�f�^��C�I�7��5F��2g�$�b�$ ��C��N�*=`�	ǹ����f�M{�C�	 [��Ы��: ۠!Q�,G�B������mͯ1~%!������B�	
;��rpc�(m$UZ �C���C�I�&��`fW��bWZ9kӲC�	(�3��I	D^ԩ9g��#)�B�I�h`��QF�Jf�u�GF˾b*�C�	��0s�R$D ��zV̋�Q�B� 7/u�#��<vt%�d	-��C䉄V���d B�`���T	�u��C�	7��!h�* D�Ht�ƹTk�B�	�Vl���)I$��yb�%��X��B��$x�\���N�p��e��탢C8�B���
��7;pd��c߄TH�B�0�fa�H�[E ����KݰB䉆D�؝� &P?M����M��?�@B�	-P����U�`�:dҦ��w $B�ɐp�2�2�.���;�G	�v�B�I�VdBD�J�j���T���T�B�I��Dʁ���~5{E

�h��B�h)�U�Fc_�u�������_�,B�c,VD�S����@ٹ�eݝJ^B�ə�n�B�  YP�T��A�?x46B�*8�B$��*��p�����ۭ�B�ɶH�с��u��HZ ��<�TC�ɿ���+�9?N��q@eץy$LB��0'�]B��Y�u:z�H�ҹ>3fB�I#^������]�N��WK�hB䉑\O����l
|p��B�A� �C䉏�,i��m�)R�����
ÊB�IM����Y�L�]8��O%C�~B��%<��(�0b[*���%a�1YPB䉺xC�P`��d�Z�a׋�NB�I�Q�����eߓ>� 13 ��Td�B�)� :��A"�� ()K����N� �"ODu�!F34FE &ލ2����"O���1! .$r�����1b�"Of] %ʾ\*p�I��J����"OT�jDj�� q�)�> m D�$��BُDVک��ڷex^P��$9D�@	@l_�4\�ˢɗ'�:p�&6D�|�l�*`���Pl�2�$�@5D���Qnܱ$̔���׀rc]��`)D�x��e�+�`D�jյv��p�4(2D� �N�)j�-�7OS? ��xZ3F.D�hX`c�<�B��p��V;x��!{����̅�
x-Ec�?�U ��"�|�D�k��\���2�N()��I��k�,9�$��<(t����F�@ن��P���c["8g@i�ǋ5F��	�ȓW�F13@�)b*� ���m޸ȅ�q$����x:�����ȅȓ1de�¥.�TY�Dζ<<L���@h��@�}�$Tg�Q��$Յ�	D�' (��&F��@%L3��Q��2�Sb��d}r�t�T�
�V$���c� �B�� 8/�pY�	�9b�< ���(�U��~2C�>.Ζ���Iۣd!��g���93F���
��9BbX�䙒�(�~�p�eA�pr��7
�)X�ѫ&��_�r~�)��R5�ڻ	t���H��_T�iq�[�U⮹'�x;��$�Z��r���*U���;Sd����EH�Iw/��p'o5���3��P#2�oF7J$�{#��`@#�n�L�O<E�4-5\�����b6s��lA��y�8-�e;� ��~ʎ��W!^�Y�5Y<�p����H�~q��'n*]��C�>�~��ҟB��#`|����K�,M�!���$�/��]�t"��&�l�#��{��04 �~�4��19#x��)/�i>#<�eɰs�T��.^"02�B���>��T?�J�Ȋ8;"<h������h1�>D���L0�\������BD0D���͉�#4Ɖ�����+$����)-D�d��H�7;�$�S��I3>=>���>D��Ѱ�L b,B��%I6x V�jF.!D�LH�����p�D�k�>D�P�2D�����ۂAP$�{���5h8�s$&D��a6�_	��"B�P��8��#D�L��m�"����Qۋ����֋3D�DA�K�3o&]Y�׽YT(���1D�,9���A=H�.T(,��A�l0D����ӈ�yp�Q��$(b�(D��RdP'@�F�8 �!q�AD&D�t���P �N��,ݣ
��m"�"D�Db&
�.O<0����+=� a�?D�����j���9��_j}	!� D�T���p�� ����<hȞHZ��0D�����ي�2�B�?u�(��D�0D���W=p�܈���X�h�')D��R�%Z�i�(p�An��%N:a(�#D�� $�13Z}[ǤQ�d<��p4D�l:7IM�RnYPAQ78C��Y��0D�{��_�~�R�st<��@N2D���@+o{h�)s��0ZQ'`.D�|(h�~"B �0M! FE9�&(D�8�[�p�R�R�O� fD� �;D����f�(��DPS� *X2Ӥ�6D���1�æHE���F�̕�R3D��aM|�pGAP��a�7D�h�
� ;�fmp$`[ $��Re4D��0R��5�X��*!xv꘱�?D�����"����Ϙ�Q)��	1D�̓���OP��!F�ר��E0D�� h@�c�2x���Q)؎�JaBT"O�S�
�B�\av��GV�<Zg"Oq�
�N�h�(�-D=s����r"O�r�kAGC����ѽO��Ұ"O�ͩ�h�ꀰ"�.��O�s�"O��BpI�.Ն!A�M��e����"O,�1���P��v-ƙrȆ ��"O�x�b�=�.qSs��/Tl�"O�Jg���#�� *���.M��@s"OT�s�	���Ŕ#k�4�1�Pt�<1Q"_`'���A��4o>����z�<I�nW�-�¸(`� �lX0��%�DO�<aP `��0�A�S�?<88�:B��z=�B��%�����ڦ?�B�	xt,�۸5�a��g6U[�B�$J���U  uax�̔�N��B䉛<N,a qbQyV��('��R�~B䉲HҌm�䧜�nC�,{�N^'a�C�I}����d�+��t�$�۔e�B�ɍAa��Z��{�t�:��Z.	Y�B䉤LX8�� �<q%"ŋ���7F�B�	�!�@%1Ə�C���Hp�E%%�C䉦
	ڸ0�	�$�!Fd��~��C�	�Dh�9 W BǬݩ����B�0c�	�B!� n�9eV%B����XSU�U�D�*uD�7ڰB�ɺ+(^�C`'B7�Ѩը�(f�B�I�&&����ڌB� �ч&��vB�	�i�`��"��d��hQ��:hB�	p�����V��db�n\�K?�B�I����v`�5Fİ��2V_C�	w��B�Jϭ&�tۗcވ#w�B�	��pC%X&$:�QTl�=:C䉁Z��uCĦ�Mr�sT�Ӊ?d�B�g�l��O+U���,���p"O�죖��"�����<]JB"O�h�'�	g���mF2\���`"O��! N�j������>��`2"O6e���("�m�0�W
S�y��"OX�B"�C��	�֤R�x��"O�m&2d'L�:Ǆ��Tp}��"OX���k�/	���*���2_�uq�"O�!��.l3v$�� �+d���U"O�ɓ��T�����8ih*9�"O�zԫ� 3!���W��|S�#R"O�i�������D/HJ��{�"O`L�Ŧ "Y�T5Ҡ�Y���Hѵ"O�A BAմVebYk���Y����F"O*y���J�4�:T�J�D��y;`"O��J��~<*0Q3'\&7���H�"OL����A�v������e��5"O�Ъԉ2Er�Ї$Z3iB���"O�8
DC� .u�a!�.WW��Z"O� �Y->|4���UI�@��"O��c�_!i�Q�����d*�['"O692Vm�1�`8q��ϐg��"O��[6jV�]�
	�$fl���&"Op�(WL�&��h�r"�V:^��"Oy�g�B�Z:0��5�/1d�{&"O,��$��>]q���oX�u�E�"OH�r�L�'h�����ѧX��H��'���!�P?�@��"O�-J~�1 	�'Lmk��\"t���B�h�H���p�'*�-:wʋnV ��˓9�R�i
��� V�#3��,�Z`*b��pk� �"O�ٔ��q�p߄JRLXP"Oj��2j��j���_<-^$��"O|��R,�	:����bݟ� 
'"O @B���/x�JX��%g�� "O���e@�K�\�h�c[%~8�y�&"OZm�W�ҥ�@��vD�A�D��y�aW�I�ؘPO��B�pa��
�y�L�Sj����A�%� qn��y"FV=+p֠Z4�
�3�"�@ª�y"H��J����Ѫ���"�j�>�y�G���8�˕��f�iw�F��y�B�FQL��u��6&���a��$�y�) �q�~L��ğ5?ƙ�'2�y�E�<&�8��!.���P���yrlƛJ������!�9��%Q��y��U�>��`��f��	�p��y���"n�0��&�I ����+��y�kz�jUrS�B��b�˳����yBC�=\>$���ʑ.��&^'�y�'%�d�ʕm�z"ʡY���"�y��&b��`ʧ.�:th���j"�y�C�W����f�چu����� �y�.��n��T������K�H1�y2�EH�hH�H��x@}r�H��y�i�?s~�ċ$��\�=�HI��y"�>V���R7WQ�d*&IG��y�Ʈ3�L4Z���M@ !���y"/�,Q���	!�
*�r���y�B��h۠�ʫ	�(]
�MB�y�F�����Κ�t�� �9�yb��>f�T��d��L5$� 6���y��,/A�{��Z��Ţ[�:EJ�'� ۤ�ۍ���2o��@�"O�T�P�X�ȍ��h���[�"O�E�I� a��ěd�K�V�&�
6"Oʕzgo�^⺰�-�<s����"O�P�LR4���uC��,WԱ�"O�`pV��7��bl����@"O����$�t�vHރ��Q�"O�r@Õ6((D�H�f����r�"O~�H���[�8aŔ�|���!"O���dLB�F\�#£D�7���B4"O���S$�)	m�}Hr"�?T��"ON���+��n�Ny;w��i��!�""Oh�ӤȌ~�����@Y���`"O�!P2�XP6�EMUf,���"O��3��T:F����M��	F8�Z�"Or�2�½x�Bp,O�>��Z�"O�8HcIK�k ��6j��U9"UH�"O�X��/ЁG�� ���5���"O10�a�<5۸�A(ʵA�^�aQ"OLT���
7�����ˋFt��kq"O����Q%|RCBM:`��C"Oda9B��|�b��m�?K,��q"O�4 U��nԆ!�g,M�]=:	��"O4�Å�tZ6<k�M�;=7�"OR��(U�)7�=��l��&����`"OF�� �``�����;J|��"OdZ%��;pV�bE]�Řq"O�A;�휬[�f�p"'� x�Y��"Oj�95�?}��́g�Ll��)"O�M��ҿW�R[�f �c���)�"O������2\��E���
;Z��F"O� �X;��XaT4-���I/f9�"O�+�$E�H�zm�U�̛,�%3D"Or�mK��bl��>	��3�"O~�A�o�-u�� 0��+B�K"O���"�0d?�H�r!��?�l�ZP"O.�3PKK';e�Ȁ��`-x��"O&�!'M��f/`����"O��B�-V
H�B|y�hQ0�8H�c"O�Ek���+
�v����Q�#�����"O����c�7�\ɻ��@�&~��R�"O��I�oҩgzN�qT!N�taBX�g"O��rA�){�Ys%�-4���"O�L�%i�;/�n���C��.����"O�)2Mˬ�n�#s霔T�8�$"O�@��M>���cI�&���"O<��"Q�B��G̠�����"OdEYF��7�yb��Pt��"Oj	
�#��=�F���ƚa�(X"Ob����<<�0�p06K蚑ص"O�$�`�ޖ�!�m�5c�lZ"O  z�i���0�ˇ�K��{�"Oz]z ��;���J΁)�ٹ�"O�x�6(��e�� Fv	����"Ozac�`J#�n�k ��_�ԉ�"O������ToX�pc ��N���"O0��(&qvU�qB$L�"O�D��eH�&g��J��E�#Xn)T"O�\�D�1{����$҃D��j#"OB�p�i�)��S��� `4�]��"Ov|�ԉA��@�JQ
�20lQs0"O	�W���H�M)���"O
��&(E�0�0��H>�С&"O�K�-�<6t	p Ám(X�
U"O�����ޗy
����Hեg����"OxY�+��8������d�~��r"O$� �4�n�i�Сv�L4�c"O�-��50���A�&brH8w"O�@���Vrj]��ֲ*���"O��@P�5*� �@�����"O��#�iX)J��%Zg�V�VI&�y�"O�e�"���z�Xq��̘*D����"O�Ȑ�   ��     �  �  �  �+  8  -D  ZP  �[  g  ^r  t|  ��  ��  ��  u�  .�  r�   �  ��  ��  
�  L�  ��  ��  Z�  ��  �  ��  �  \ �	 � 1 � e# d, �; oG �O �^ k xr �x �~ Ӄ  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!%�G{���oόQv����V�k�ظZ��M:�yR�ч@.�`�f� h�Ji*�m����HO����c��;@D9���[�hMK"O0�h#ԌN͑��V�V��1�"O�P���)Fn1��/̸"���"OԨ�S��Z�\lK(���d�"OH� f|�9�	� �l
E�`8����! 0Z<0�ӕT�6�9D���婌�s��D�C�#\jܨ�d6D�p#��� �ô�O 1h41�!6D��t��]	XC%$Pp� S� ���p=Q�ѠT���gѕ8���`/'�T���π �@�5㆖/�pa6�nլ�s�"O~�k�ȅ&'L,�D _-�u�9�=�xN ������J��A�.�-�������?)�B	mj�L�#�B
�H)1�@$!�W�w�\��@/Ş��Q���F�ax���v��c}��$Oa�A�E��u��L��J��yrf�b��"�0Z�PL�Pg��hO���IL�v���: O/6|���� �h!�$�%�lZ�Nr]���D��sMay�F&g�z����֖X��R�xu�U��	l}2-SJ Pa��X0&�؅1�@��'���$9\5�e@�� D0���)P/��$ �k7�+2,B�@7��4�#�ZQ�i���5�O�}�W�_=�B��嘏$j�`1"O���N�w.��㗪.PX� "O>�o�6D����h�9�G�|��)��{�d��!k�8$d��+Аv�h���<����]d*娂߾~*��E@f�<�M��S�����B;Z$�d��l�<YGGU)#�N�p�)�9}��|8�B�A�<!�,�w���CK�1	�p���mR�<���o��h)��R�t�lU0w`Gw�<aA��{���T H�a �ɀj�G�<YF��-s#D�iw��<u��sA�o�<�ƜMJ�A2D��^g�{ *�d�<I�+��g�P�ʑ�v��ӭ�w<a�pl�`�"�$K��1��!O�nhT�ȓ:vT�j�S@Or�`�c��
a܍��!�ܰ%+�4TœWlS�1ܚa�ȓL�i"�m�;���m]�f�ƨ��o���XBc�|u�؃T182�ȓ	���I
�K���E.2�8����'��#}�'�<b&ŗ8+ E(#��Z!��'f:d�q@�;_� 	�2,ǙX4(��'-�UB�O�MW(�����"�dH��'`Y�A�F��-ӡlX9Iʬ��'
�}����w �q�@�?��� ���(Or��Ϗ�7��Ո0�аVxH`�"O��$AG�S�΁R�,[�-��l�&�i ���� �� ��m�?i���z 	՗Xa{��K;�<��a�[1��a"�I+4W!�	%��)��̗s�P�;�H�8iޱOʣ=%>� �j�
	�Ĳ�d�mP���$D���:~ ȡ��SCǪ��ЀN��HO^L��	�/��ct��rQ+C�D�<�B�ɥR��9P�ՅH2��)U��C�2
��ѓ�.T�D��r�
�	BB�	�E��Cu��*���b�MÃY*B��Lx�1�jFqf�[�A�`T�C�Ʉ����	ǿ%w ��q��Y��C�	&�R��)T1�VP)��S�m��C�	_k�u���Q�L��Uy�'�*�C��6F) tD���t�0�S�}:�B��o�(U�&�۝)ށ[%"��V!^B�/=�\`�E���Q��B��̑1b�B䉼C�:�#�ՆP��2�.%�B䉉���+��&B ����)d\B�I#��a`"|�xY�7+����C䉧]�N�hV��`E��H6�~��C�	(�ʬ!��%,l1�uϋ�x�B�	�E�غ�D��b�
�	�GF]��B�	�����	�*\��;��� ފB�I7-4���,M2E�����&�Y�*B�I�_����$��2�D�GkB�)� ��� C09lZQ0$o�8Tcth4"OH�y�̃01I��P���aWpa�'"O��+����V3��q-ϗqbN]Z"O,ՠ�dG�_��H�%�G�(r`"O��0�ł� �4�Ӕ
�iD3�"O6ik����͈���(ۘ|3z�JR"O��h'K��1[޹�rg��
��A�"O&i1�A
8g��S6F�4�T|h&"O�9�7g�,@.��d�Z���{E"OQ3JB2M.��p�N�����"O��☏\�n3��V����	B"Or�3���9r��L�I�� НQ�"OP�!B�;zf�����6�NP��"O�5r%d�g���Ǔ�pо9�"O�8B&G\�+C�x���&R.��Q"Ob�YWD�,S.�9�V�[�pQ�"O�B3'WC��53T`�)���"Ob�bT��9]����Oڼ|���s�"O*�I��̃��mys/��)T��&"O�ȠTA��B��� ^	@����"O-3�HP�9��}�����B�Š�"O$4ip��;*uyh O�(k��Qڥ"O>��d�I����d���b{�e�'"O�� sN�9N@�\��ƕ�|[x̒�"O��hU�Z��s��Ƀ#��88E"Ox��eψx�l�a*Y."���"O�m2&9{$V)c�Iޯ`�T���"Oh=B�<6t8
�o�r�F��"O2�5���p�y�oK�s�r���"O�ă�蓱O�X�r׎þX�~�1"O,��	7��@`CM�����"OF�KMZ�Pl cpB�&N�h���"O�]�Pψ=,�*����4�ޥk�"Or|X*O6�����Kã��u"O~\j�n�L���hQ�74�,��"O���G)Ʋb=n6`ө
0�I
4D�ȐI!W�ȡ���������.D��"�`�7M̙�O�s# �Պ,D�4� ��d4õAJ�v4�Yq�*D�0�gnʝj��Q�W��Z����A*D��C�D�j�Ik�(���\�u�3D�;���>Fy�[��с&���'D�4S��.0pe�'�ĵF����9D����O��da.mR`��R��qԨ3D�H���bk�[�	Ee�����=D�4Y��ŕx���G�`�� �O8D��6B��_����C�"ZM�vm(D��IUiY�H��%���;��)�'D��*4ƒZT4u���7t���B�)D�DĜ����'']܌Ġ��&D�@i0��ChM�BnǞj�X��c D���C&;sʵ	�E��"DU2@�#D�"T���-�Z��df�([	.����%D�0Kv���D����!����삄&7D����%�F�*�@��(�~8�34D���JM!ܴ�1�����L@��3D���g�Oz��um�`�v���2D��87"�N��p�A�'Vrx�a#>D�D��C�j��Ƀ��
7�6�" C6D�8�`�>0'
�3ѣ-�R�o3D�Xu���u^�I���(Fn�%�P &D��"�2�d`c��r:ʅ`�0D��o�d�j��D+�+uB2���s�<!�D��~%֠k3�֮�4%z�Nq�<� ���@aK�;�X�0���m��HC�"O,�;�_�?�r�C@(�.w|R5Ku"Of�;tiϨl�8���(VV Lp�"O�l��a"���G'״G�)&"O�\а�F�_�
���⇻G;|�s��'���'i��'�R�'�B�'12�'�(�@]55��[��])z��5�'b�'���'�B�'���'q��'p$Xc�D?=� ��)Z%��2��'�b�'��'M��'���'x��'� XPᓣ"=*�K�C�k�\��'~r�'W"�'gB�'2b�'u��'p��(fG��8N]����68���Y��'F�'��'
2�'��'�r�'�������V�L hV��7	]V�2��'t"�'qB�'x�'���'(R�'
����h+,l�,
ӡ��ڀi���'���'��'��';�'���'�ʝ �{,�	Y1�E':(9x��'���'�R�'���'sb�'b��'��8a�ؒ
S���JH�j��'���'b��'���'���'���' L���jΚ=�H��H��E;��'���'C��'8R�'��'�R�'��h3h՟F ��s��z����'���'jB�'&��'6r�'���'��pJ'��-�$\*f�s�ؕ�#�'=2�'z��'���'�r�'���'3����j�^�"�`$�؃7����g�'���'y��'�b�'Zҋx�Z���O"�z6��I��y)����� -���jy��'��)�3?�E�i��٧����Xr�BS�.kf�ja(\���N⦩�?��<1�iqP�m�%�j��ĩ����� pӔ��7��7�&?��Xj�ԥ�4�"�+�*
��;p�,��P�TBǰ��'�BR��G��DY�y�e�'J���ys���W�7-	�,�1O��?]����{�i�nY  !��$��Hu��w���k�h�p}���$()ś�5OhpעѨM/��#�)C��U4ON��"?�>��� ,��|��U������M$rZ��-؃XI���:����QCЊ8�	{nL�:Zy�(��E��o�R�����?F�Ƥb���G}b�(S��P�[�|egV�����9R�VH���B-xX1��`�ob�a9�u:6dۡ��e�2��/ь�JY/O���?E��'�<��F�0�t�y6��%ر �'@6M�r�����M��O�8� ���=�q�vE�
�ԥ@�'��7m��	�	�k�T}nZs~�F
�č��O�`�\<��X�&�R���� �+J�T�|�U����t��ğ�	�4���D8�$:7MؾL�L�eiy2�{�fa�t �OB���O
���$_.$E��8�ƅ��pk7��J`F��'�7�Y�5ϓ��'����]x2���P�5a�$Ӷʃ��:�b�!�C�Vx�w�,�zP� K.��^w��'���'�t�7ʑ0x�V��t�=v",;��'�B�'*�����^����45�	2�(�a nZ�(ٺYD��@S*��+���Ax}2`u��mZ՟�;��]�$��ͨFO�c
�Rп/�6%l��<��/MHT���� [�7��ۛ��U�� $kS5-�ҝ��qb��s�n>=X��O����O����OH�#�S7)����K9D��h)��2a�}������	�MSGfM������y$���f�J�+\IFܸ�I�t(��<��O��m��MϧN:*(aٴ�~b�Q��uR�R: ��X���?$���z�cJ�6c���	ғ4�ʓ+�ʀ�*O�d�O����O���te�*����m��t3"���d�O��d�<Yĵi{~P���'lr�'���5��- �ւ%C1�	B˸�,��)�M�Ʋi���%�Ӈ��H��&UF�4�cմ�h��*R
*8�FȕSy��e݉Q�E��suP��]�f��Baх~M�2%�	]�� ���h�	ȟ �)��Byr�~�ȁP׎Y�e;�����T]g��b�Up�˓xB���dUT}¢l�4��@��9"J���ԬmK�U��FȦm�I��64o��<���ޖ h'ń1lͲ,Q-OX����R?2��� c�/4�D��Y�'2B�'��'���'��ST�&�I��¥;i2P�ai�:w ��ܴ1��L���?1�����<�տ�y7�Y��&���:�ȑ���[7�7�Q�͓��4�|�)�O ��fnf�j�	q�j��RO�=o����B^!��i]5���~���R�@�ڴ���O���F�f�!TI����$��_�YyR���O����O��sS��f�
I.�'�b�Xʴu��,KH�x��~��O���'J�7MI٦����$T�jW�ĀE�M�IS P���v����O�X��P��x�.�<Ⴒ��Ys�eݭ�lK�t�"£>�cD�5,�fA���?)��?����h���d+&�n��@]Cx���Z�Ee~���Φ!�ˈOy��w�Z��82�PTzpiR~J�(��ᖃ�J�I�M��i<r,���V2Ob�d����	�$ʓ�(|m��H ��C�ҿG��b�<1 �i����T�	ʟd�I���ɩ?��`f�c����u�4�'2�7�]�j�$�O(������<��n�?j�v!��U�m��|���w��I��Mۂ�i��D?�I�����(�`���+�h|µ �8[�f9@"�0\��D�ʇ&ʨ�u�Ŵ<a4�i��I}��Y�f玞R0��(s�S@~��	�����ݟL�i>m�'l�6m :����k���!� ^��A�qb�����ߦ���z�I��DӦ�Q�44C����m��E ���Q��h��Oݬ��YY��ii���O�[�Ø!\�I�Df�<��'�C�� ���ŧ�wfa�2�-!��l��?OH�$�OL���O���O��?yye��0��=U�	�<a+��h�������4>oB �'U`7�'���# ��#Ǝ�H���:P�U�P*�1��x}rh�O7M��RPJr�c��I��<{j�92h��sA�1 ��܋6(��e��#C��9dԙ&���'�B�'Kb�'�vR'���瞸L����'FRT�t��4Q�=͓�?����IG)�����kN�L��ġʞ��I
����ڦ�)�4nnr��d�O>ݐ�\;_t��&I\�^�0���%3�,�nQ��'�`�釅N��3Xw�&ӧ5&-�`�T@�"�c�-��G+�2�'��')���R� ��4���d&����I29��QWN�X~҆e������OT�o�(��1d��,,Z�z���H����ڴ'��槍�Lϛ61O�$K!3��=QSMW62ʓ7jv �5c_�A�l����\a2�Γ����O���O��O��D�|��ѱ�~Q+���&쨄�e��&ʛ���yr�'�B�O0�s��+���+�G<?H%B�-�P����l͟bj���`�a��x}�OB�D�O�P(sôir�d�<r��Rr�>+
�� �F��D+u�c3e �6��O��?���P�� �u��hU1b�;uC�H����?Y���?�-O�qm�%&=��	���I:;��`ӄتu�]	��[���Iv� ��$⦭��4.b�R��#O=[mHpb0�@�1�,[Gc���I"� ���b�v�*$�'��dIX���B����d��Ux�0��,��@��MПh�	����	ٟ�$?��	�#"*���=e>$
�'�Ms^�j��O&Nຘ�I&�M��)Ŋ�� ˦M&�`�iޥ:�g���L}b$��¬���k�8���"ٴf!�v��ߛf3O��[���{C�U	;���.� N_*�@FQ+v��8�%��Oʓ���Op���Ot�d�O�v�d 3e-S�0�$S &<�ɂ�<�#�ii�� �ɓc��'o��O"�8�A��IG�a�����`��C*��O�Yo�;�M�ֳi�>�$������@��Q.~50�L��q,�����GkbE`6�<�WܲM�]w#|�d�<)Of��1C��< ����Y)�3��O����O���O�lz�L�<	g�iPX��O�)�v�#�ĥh�ܭP�'�z7�!�4�@��'Nd6�Q��-�ߴf����%L��,h��[�&��ě�?�M˜'�re�wi<fFШ�]���S��5V�E8���B/{ R`�A�m�2�'Y��'*��'�2�'ܬ�e��:�9z$��7#ԙ�C8y�VI2b^�bR̂�'L�
r�����1O�U��8�P�Ot�)�*Gse3��F	^���I�l�2�;��L��F�hӒHn��?0�oZ�<���)�L!�����*�(uhZ�hGV�8�,�j��P�ah��?�.O�˓�?	���?)�c\�T�=��k$m����� ڠ�{)OF�l��.Y����ʟt���?Y�S�FGj	�!I��L�z��VǛc�v����[�O||oZ�Mc6�i����I�-�x�ćB3+,�9�@��1��c�pQ��<I��q|�l Zw>�ON4�4�Z7Z�d�$y�: ��O����O(���O1�bʓv��Ǐ;J,�D�ֵ5�j���/8Jo����R��3�4�?qK>�U[���ڴyf֥b���0�hy��x�be�i��7M��X4�7�n����1u�t�2D�[o���'MP�rE��;<�F\i�c�6����'���ϟ��ǟ ����	a�da�p<PH���/l]��+d�"g�6��M7�d�O��d"�9O6�ozލ���f�(Ta�Y�)�h(��ո�M�r�i^��D�>ͧ�:�';�|M��4�y� ф
@����ٗ-KF��E�0�y�ƙ$Z��eѤ�\��'��I���I;�Љ�U<|��J�j�]f4�IΟD���l�'#�6-�K���D�O��dމ�V �q�+�b�biI�o)��D%�$�c}��c�*�l��?i�O��D�}]��U��n��첑2O����A��xǦX1Z$d����ֺ�uGb�O�P�aϤ���J!�1�n��r��O^���O����O�}���
�����B�n)���o��!���a$�F͉����	�	�?ͻX��02�$"{Fa��Qg�fQ�C��F+n�L1l0c�=l��<!�f^| ���[�����)�x���Q�_��M��[������Ob���O���O�����jYR���+�R@-Y�mA@�}#�ƀ�h�b�'�����'ix����<�������T1�>���i�&6�џ�&>���?�Y7υ&Z���[D�ԣvO��A0�D<"�P� �hyR�>n�L����'�P�'��:fT�\7�(���@�f�J����'vr�'����U�D��4 $BAH�s��	�e�N5s�p@d`��70z}Γq%��$�M}�c�^�l8�MC��.W5���[5�&�i��J.M���`�o����c?
D�x=�-i.�<��'ukkL�C� �*�47a�m8B,cy�$�O��d�Or�d�OT�4�S�+�H�И_<��b��5L�\�IΟ��ɩ�M#�i����$릭&���͂)s1���%���@T�0�?��OD�m�-�M���1�F�j�4�y��'��M���Ƞ>t�� K�\�%�� E�T��H=~��'���P���P�	.oJ�l	�Y�}���p��%y����	$�'��7-��R[��O`�$�|:S�[h�1��ҹ#��Y7DI[~���>Yq�i��7-%�4���)E�/��e�g�u҅f�32���ᘔ)In!Ir�<i��5L�Ĉ]w��O��1V�Se�f�HP�\`؀s�O��$�OZ��O1���dD��i��3RP���[��8�|A�aI'5V��'�46�"�ɡ��dKۦ�� Q�o�n)�����b�.8jR/V0�M#����J�4�y��'���qU.Z̆I��X�� �e�&�3M��{�+��W|��0O��?����?���?�����iM�O����j�T�`}��)����n�~�F���ퟤ�IZ�S������V ��1�֐�Sa�;2��l� ���%�6*r���O���\��E��*7�m���S� RyV���dA���sQ�j��!UOx�Y dE�y��Cyr�'t�ND Vg��Q�E�6t,p׊��w�r�'B�'��I�M�%m�?)��?y���&�T%*g���R\�c#�M���'6��f��V"x�H�Of��t�@�"@N�I���˾�Z�4O��I�ۛ"�Da�4��*Ab�i�ѯ�@	�Z������:�P�X���^���%�@�%r��	���	䟘�	r�O����;Y�`��@T(~I�5�ĩ�1@l�\!A1��L�ܴ�?yM>�;z��g$/
���"ah0��1�MÁ�i��7�ȵ^~�7Mj����l�6j�����y���j�F��(���afF

�B%b�r�M���d�O:�$�O����O0�DӾ(� ����Z5kD�)��1Kx˓f�f����$�O��?)�n�2s"Z��s!�c�A��$��DTߦ�[޴mA��4�O����	 ��c�/t�`gԠ)�@�22�n��,O� pgh^9��]8���򤐚:rأ,M6l��A�lB/�z�D�Op�$�O��4�fʓqW�&��r��鏋$x�99˘uNы ��y�B|�n�Љ�Oj�n��M#÷i}>PI��&�SwCä�ə��ۜYy�4O��� %�j���� AM�ʓ��ñƈb�JN?p����2�a�"�h�9O��$�O���O(�D�O �?u��G޼j ��񇏅*9��(�.�ן��	��<p۴|E���*OL�lC�ɯ�*�JP �B!��ˣ��Z[n�R����٦�Kݴ�� ���MC�'�2)��\H3����A�X���}4�-�  �Qva��|R���I�IƟ��Ѓx4�!$�V�cGEN˟���gyr�z��
T��O8���O����Ƽ����?^�آ��Q�	�Dف���(�O`8m��M��'��O5��I� � ���[?!�ؕ��g�����Z0�D�y2_����<|�FQ��'��'��X8��FKH�j��MDk6���'���'���O��I��M+��Q�MA1oɅ�]���	36��`(O�0n�䟴%����O�fӔ�p6�S �����*ÜU�hm�R�[����4e3=��4�y��'���a�g��_��i`g�%@�8С�U����r*n�P�'�2�'p��'2��'��S�!���R�K$��M������4LT^l���?q�����<���yg މVD��1É��:��|���aF�7�@ܦi�����4���������� rӞ�ɯM_�@X�ɓv��z�)Q�b�	�U�x�vO̾���'���'�B�'i`��PkC�?=65��镙i��I�d�'�"�'�RY���4A������?���#�8|x�����X'�@�vNؼb�r��>y��iFb7�\ԟx�'���5 �4��I��( ��\!�'QH��`	�	&C�T��I�?�B��ǺK�'~$EC ś�l*��#Ω
�V\5�'}�'B�'Q�>���7�(B�+�/�J �2c-��\����M���J~B�f�4���6�@M��
pF ٚ���'vBx�ɔ�M�־i��7m�&�7�u�@��%x����G���5�@)R�	X�Dj�8���#�~x6c�z�Ty��'��'"�'�B�D]����>m��Ka�t�Ay��qӊt�c2O ���O����� "%��������P�th�1Z�<@�'�b6M�צ�*����'�R��}��Y���F5�Tc�b�6l0�r��3n>Da/Ofذ�e_��h�]����$Γ:�:�`��H-i|����
�v���O����On�4���7x��폇Gs��ɮͰ���yJ\(�$!F��yB�r�X�88�O�l���M[Ŵis����Sx�R @���O�Uie��@��?O��$��6�v�P�Iиg��˓��ð��I�F�ʐf@t�.�#6��C;O��D�O�D�O��D�O4�?ݪ�HS0X�xY �$T��i�G� ��ԟ4��4-��-O`l�b�I�^L�%��O��  �F�|�������$���p�4��dNJ"�M�'(ҩ�t[� ����mz�H�	�=�r	�7h��X� �|2Y���������h��^�dȒ'g2@��q��ݟd��xyrO`�t��r?O��$�O�˧IXv�'l�8�I�c�_��8�'t��a�6i���I[���?�"��8�4�!_�jA��r�Y5"���2�L�:b著'��d�"ay�a�	��p�z��Λ{x����3(�0�	蟌���)�Siy�b�pp��ĕ�`��i%�G_�,đG+
�IX�5F�V�'P�'0��HA��'�,����c�Ҩ<y:�;3ḋS�6M���H�)	�͓�?)E�X���;0̙��H$nؼ���?⽠ ����<���?y���?���?�-��M��@#��� �8)� �ڦ�`���ݟ��	埴'?�����M�;x�
$ӑc�3��@�j��قa�i��6M#�4����OX��)h�v�	T:�` � 'Zf�R��)��<����f�1.�%���'F2�'88  �M_�i�̍7r�^����'O�'�b_�T�ڴр�j���?���pd�qB��B�����eʷ�����'�>�7�iE 7֦��O���3�����V����;O�������c�H�!\���zMO<�uGK�O��Kw�^Ij- ʐ�7Q�U{���O��$�OR���O��}�� m��bEa^�JF�a��N�(�b�X/�6iI*?���M���w��`@���
�2<#�Y ���'<6M@Φ�a�4i��y!ٴ���bR����YMH� ��:ӈ(l��PIgE�D�hQb#��<����?����?I���y2EנU��Ԃ B��#��6����DAƦ=p ��8���D$?�ɼ��DPT�c�H���)�ХҩO�ao���M��'9�O����O���`��)Y�̈C,ڞTT���X#���Q�����G	w����/X�''剐z`�8�A�K�a�0=�v"ĻH�P��͟��I��i>}�'��7-�!p���5-=Ӈ��=~v �r�_J]�d��-��N�I���D���ڴ՛��@<9��H g�#K��!���������i����Ory²�P�S��M�Dι<���&klըJ����3`��W��l@���*G}���O,���OT���OT��-�(~۬m�fg��Dě!f��	��@����M�5����H���&��� O�%��} �o��F���p���*�?A�O<�nZ,�M��'t�2�4�y2�'����Q�"��[pH.~�Fbsoݘ�L�vȎ���'���㟐�I����	�;���0��@�V���P�T���ܟx�'gb6Mѝlx����O���|���e�.�7lи1	L-���N~�
�>��iv6���L'>��S%N�B`�mw�T9t��t�i�$h����4��HNGyb�O�F@6���P%��;�N�?Vn�Ȑ�
Y6���c�����ğ���ϟb>��'�x6�8VZ��u�Y���P�D�ȯ(��c0�<yp�iD�O�P�'��7m�U�X;&IEv�E�q��"q�f�mZ��M�1C�
�M��O�T�n�F��u��<�E#�C���Q�hh��e���<!,O����O����O��D�O��'Il.Tbrg�(%H蘰�B2t�F�At�i\�d2��'B�'���y"kp��nI��Ҩв��b�E�'s	mZ��M��'��)�Ӷ7��n��<�c�.���iB#zbh���<Q�^^��(P��Ʃ�����O���TSt��P��#"q;�j�;w����O���O�ʓf�F����'��f�2������)r6H��4	��a�O�-�'r�6��ߦ�8���D��=$d4�1��Z�N�!�%���I �6��PH�S�z�&?��1�Ϻ�5�'�tQ(�oK���Y��JA�*�<���'���'���'��>E�I[�	8�g1OI�x�E��[�L����M#�i����L�a�?ͻJ�@<r/�t&�@�E
L�P-� כf�`�h�m�]�t-l��<I�b.,����u�D=��N�b��-S�EBM���$\�����D�O����OP���Oh���C5h{e���s�޵���%
�d������\U�	�8��R�W�!��	���<b��h�N(��/�M# �i=���"�i��I+\X����)� Up��0/�=e�!�a E	�˓Z��a�M �uW	9�ħ<	� �<�h�i��N90��8	N��?!���?����?ͧ����僤������foœr	��	jL�з�e�d�4��'C"�2 ��{��]o24�N<CE�
(D�D�s�>h�*�a��Ʀm��?�� E���e͌��d������2�:�J�(���p6L��}2���?���?����?1����O?�P ��v?�8��O�X��-���'�2�'�6�Ҿ ~ʓ2h���|Ɩ����]2o���DL� gj�d�>A��i��6Mh>X��Ӧ�I��4�%� 5D����#�cɆ)�[4a[�a0U�I�P�|%�p�'^��'�b�'�4�:��lj\�n��g�"0��'E�R��Rٴ�^ �'�R�O��4]-;b�3���,[t
��fA���$�o}b%p�f�o�?�M|���q� R0��*_F���BE79��ǟ�+�(�� �^)�����U��cݕ�N>�G�:M�Z��G��^i��OԻ�?���?���?�|�)OmڽY+L�c�B�;W�4�=}�ݑbyRr��㟼�OnAn�7�Ft��A�=��l���ߠ{ѼybڴV�vj�+)8�&?Of��V�H>])��\���˓r>��U��8-�9��9�B�͓����O��$�O0���OF�D�|ږ�H�R��󕥐�lp\�%˽`⛶kʶ|���'�r���'��6=�����'tՓ��6vD9�7�Ʀ���4^�Q���?5����l��<�s�ô{�ʬ14���B��9 -��<�ƨK&�ĥ��#�������O���L8
\�,C�T<[WR����8�V�d�O����O�ʓ$�/)�''��\�n��uH��#�j�)pa�7d�O���'�(7�XЦ�������܄n������'u�:���B��mH���OLx��
�%�b!�R��<Q��On:x^wE��$ͥjξ]�!���`;(Az�I7ʞ�d�O���O���$�'�?�ǍN!c���	���"�ʼim 9�?�6�i��\�aT��z�4���y�eE?[�N� q,7.�ɋ�D��y�FwӢmZ�M�gk�)�M۝'B���9�Di��[8�(�^"^���� �Q4����|BZ� ���������۟
���k���dX��ҧ�-�=�'��7MR,zj���O���6�9O9�&��;��t0cWL��Ö+Zg}"�a��4m���?�L|r�'�2�L��p�&\a��z��T��Ȟ�_�)�
�����#+�n%�%�h�iiH>�-O(-ँ�?)�h�6 �i��0Qq��O�$�O��d�O�ɶ<��i㘀�a�'F()�e�@����q�iȺ��t��'�.6�8��2��D�צm��4 ����U�f��}iRj��^EБ���5d"�i@�D�O(56�ҠCJ���֤�<���/�k��fR�y�%D.<	���ܓ��O����OP���O���"��	T��#6�,����Y���I������I�M��T6���Ȧ��IPy�I�1z����A�]�n���g���g�R���>��i�l7���N�アyӠ���R��:� 0ҷ��t���{'�íAڜ�0�F�*V�$QP�%��<a��?����?qU��-{�@R1��0Q�n�SAW��?�����˦��FI�ly��'t��qELH�dO�1U�b���.,<.�N��	"�M�i(�D7�	��b�	5�̈́}�������'��4ᅁۚL1\�	P�]����"��(�uG�%��I�j�G�]��~���СQ����O����ON��ɱ<���i��0.�/j�7�R�e��+�"A���I�M���>Y��i���s#�&1a ��'��sX��'d{���m�@3
�n��<��'������ƃ�N�'2\���]�N@��.�R"C�<�(O���Ob��On���Obʧ\�2]�2aK�F��A�d;H�:���i~�IS�'��'���y��v��_�Zd��q��	8F ��M��+�x�o��M�E�'��i>	�S�?��`�女�p���r�ț�"Ӯ*��W
+Q�lϓ"�� [W,¾?���I>y/On�$�O(� &�2Sq�P�TϞh%u��L�O��D�O~�ķ<�i�|YП'���'p�z����c�(\r�#�w��K��d�[}��m�NlZ�?q�O
`K�1l�� ��GЄ|��"38O8�d�mk�j�ܡ����ZViM6�u��O�4�&���^���@D�+�pa�O"���O��D�O΢}λ:�C�e�K����͔�Bn��?�%�ic�	i�O^8l�l�Ӽ��O�Q�y3��!l�vZu���<)��i�t6�����ۦ���?��hӥ �6�!��A?K1���߃[�����!ڂY�O>�-O��d�O����O�D�O�u26��M�0��ؾHtT��3�<��i|�m���'���'���y��ͩ?H ��VF �iSg�83��r�f�q��@��_�O���g�3,�Ȓ����J=���C��i�0��[�D0⭊?XM�P��*��'���e�fћr��k�(�K
k�5����Iȟ��i>��';|6��0Т�$��5��h��7B��� ���#��$E¦��?��Q�4R�4&Λv�`�
)�4�A�Z��`��	�h�P"SU�7-"?a��Ł&'�������C	k�hB`�L�!,����6k���OZ�d�O��D�O~�.�� ����G�ֲ`�D����l������ɛ�Mc�����$����%�t��&�7K�vxi�iE(@��"n̖�?��O��n��Mϧ�h$��4��$+C�]�ժϮh�5*���8s�q�@�q*���9��<a���?y��?Qv'��<���i A� :=8��]��?!���D����3�Yy��'���p�|����9���T� �_�^?�	�M�ӿi�p��'�S�|<���A؜Ox+���1irH�����6����)�by�O؆P��b'��Q 'g�����	�Y�8�p���������0���b>��'�06��]�B���֡*Ib@+�Ƽ�H�%l�<93�i3R�|��>)7�ij��b'��+c��0r��?i�����bӦ(nZ/4�o��<��.���Y�gM�,`�H�/OztquB��q����3P���7O��?)��?	���?�����i�l�� `��r���f�8i�lg�ڀp0��O���O��������]!<���Vʛ�_�H��qn�;=~��4��F��Ob��|����
���$�M��'��Iؖ*�!���`l���e
�'�2�c,:M������|B\���I��D�QG��vmY�ɛ�I6�[������Iş<�Iky�Fe�*�����OV�d�O�Q����O����W�+|���֍;��,�����E*۴1_�Z�\�fޘ;�:t�%EױD%z�YSOv�����[j0��A�
w~}�'���L��:������
#��v6�x!+��p�����	���	���G�D�'7L3�%I���i4��l2��'/f7�ϕ?�ʓ6���4�|@[�	�j�\��r�ϣ��S�>O�9lZ/�M{¸i}�u˅�i����O�0갣�3^h��J�	ReD]0'H�kb�QX�/׈=Ѳ�O���?A���?��?���8�
���C�*=,���/^:f�&Q�)O�\l��|��9��ϟx��]�s�'�.#��$��{ ���n·��d�覑��42���t�OU�t(RV�4B��K%1��� I�p��iK�\���	/EJ��8��	Ⱥ+��|�R��(`��.3�)�$ü�NY��)BƟl�	`�	���Ty"�f��́D�O��B���9aA^Ă�������:Ob�o�H��u��	��Mb�i]H7MQ(� �Q�C1
�k�F ����Fe���Iԟd� �Fn6����^UyR�O�Dט8k�H�b'C��PTď3~��I�	ß������	u�'!8�pz#���mp�$�!�Ɨ
�Pa��?������%��.B�I��MS������E��#+S.Q�XXGƍ6`�=��j}¦d���o�?��%Ȧ���?Y�d�,�����J*���&�� ��mB�^���N>�,O���O��d�O�<Ғ�@V�F���(Z�Q��!³��O����<y7�i�A���'���'��8���&���I$�Wϖ�f0������M�$�iǢ�d0���Z��gɍ�5O �q���.���1�W�g����r�6a���*dL�u&1��D-�b��dIۯ&5ĩY�)�d���O,���O ��	�<�!�iE����ɛ�3�I��-&�Wl�mr�	��Ms�"I�>)4�i�.�B��dT&�r脄*>�)F�f��pmڪ
�4�l�<Y��0\Ȩ���Z�|Y Uy*O~`���_ .f��DDۢ+����-Id*UBR�E�GX�}RoH�}��2%U*:)6��Fܬ7ٮ�x��']LR��K����A�HF�$�� �G������'���K8oq�K�+�(9��e
�X&������~�����,[�*��e�cI2{YHY�v(�&%ٚ�Jb�]�� �Q����؆laSɆ	lMj�Q���X��,�A��8�D�`&�3? 1(t�����!�ʁpu9�3��L��Ժ4j/ndbt�p:� �c��(!̢p�i��'���O��O�ר0�5��*�WԼ�ʡ
�-b�(o2m��A�'Q��'��T�|R�'�e c�F�`	My��ޛh���x����O>���9{T�'��S���I���A��ߌavޤ���8'�
�@�Od��Oyc��D�OJ�D�O� �t��%)��t����9&6�у�SЦ��ɸ/R�4#O<ͧ�?qN>!g)��h)����#�,i�1CC��ɐ7�Db����ܟ��	Oy�N]$o���(E�3h׀��0&� Z�xY��?��O���Oj˓�?���#*�tC h)e���s%�S
��&�}̓�?��?Y.O�%�6�G�|*�Ƌ�Z>i�f ��h1Rl�u}��'���'��I����=
y$�`��p���MH2��Aŭw-f��'��'"[��@��H<��'.\~dȕϕrR5;�D��E��dk�i���|�V��P�=�S�*���JD#Q+;Pv�����mE�6��O��$�<�M�>T�OZ���5ƭ�?e� -!��T�8�)���Q0����$�E�>	�'q�X5"p��zΦ�3F�-	Z��oZkyR�M�7Lh7�|���'9�D�6?a�!V/}��ˢ.��5����l����'�đ��O��Z�sӲ�{��
`a�bF���MʘPвiI� 9Al���O������%��S�e��e�bMp��҅�34c:��ٴX(F��'��v�s�L��%Q�A�
�DH��c.�q;,�ٴ�?����?��W#�����'�d��mw����NM.j$4��% B�o���\y�cU���'���'���*�l9��M�;$B��@
5YS�ɐC�D��'���'"b�d�^'��&AS�T� ��4��&s��IVEY���3?����?a*O��$�37��@IB�gl��{���QxJH���<	���?!���'�2�4k萸��R�p)��)���jp�k@i�6����O��ı<A��(m��O^�ĨanVV^��ÀJ꒧*�ɦ���ݟ�In��?Q��0[�B�nZ�J��U9�'��}	���6�W�8���?������O�%�C�|��IϜ���k��T�0�A�b�����i2��d�O�5�e��4v=�'j��1��^ v�PyW	><sj�Z۴�?)O�����w\�ʧ�?����:cn��J���`@�X����>��pOp}:!��C�S���U��)�Nf�4<よ؆��D�OΑ�P��On�D�O��d䟊�Ӻ���^����'a�02,���g�H}��'jZ�s���O���/h�us��(\g�شy~�Hs��?Y���?�����4�
���,Yo>�(��w�F���Nž`�~�o�7l�Y��/�)�'�?9E&�LY�����V(D,���jכV�'x��'^�}hQ\��Sğ��Iu?��/Ж#�v|"�.�$H�Bf"ϋc1O��b��t����x�	j?)�c�10zN���E�o�ȩ"Aj撚��9XB�'"�'r������`�E�S	���H���&2��	� ���C8?y��?�.O����[W��AI��\F1We��u#̅��e�<Q��?9����'���P�k�L�񭒮-�:�hU ��!B4������D�O����<	��Ph�0�OɲAq��Q4*pq�fڧhl�tܴ�?)���?y���'ތp!���MK7���F��8��Aǆ�C}��'�2\���I�F^֥�O���5f�^A��H�<Tէ��,S6��O|����/l����+�\2&H~큑�A"8 bri-t���'�IӟH��XS���'Ib�O\����De����N()y�@��"?�	ޟD��Ʊ'��b��;�̵�␶J��@�)��
kb��'�RL_Oyr�'���'9��V���1��롇ҌH�vl��
Q�듽?�7�O7gX�M�<�~�r��z H��I@`���0-æ�h��ȟ���(���?ɔ����'� T +�M�����&Nw@���r��x
�J1O>��	�PF��QcÛ�ON��{�e��vW�TB�4�?y���?�W ���4���d�O(�I�z���(B�ʠ�%�;T���DG�B�'l���D�O\�IzE:9��\�X,�:�EL�9�P7��O^�"㫧<)��?q����'  $�c�����̊%~���L<��f~b�'Z�Q���I;q��k%ʓL>��@�M]�R80�d�zy��'���'��O����
W0��&�ׂN��3G�&9���	�� ��	����Ihy��'s���ݟ4�2�茮W�=���iypI���iOr�'�2���O�:�̝�2U���݃(|0�G)ǬoLbx������d�O
��<q�&ؐ-��	�$˼l�f�JA	��)��ʖ\�v7M�O�⟬�I�:wv��I#�S1u."��n�6U�<��A�-����'�*�A�z�4�'�R�O�\��&�-0�N(x#`]�}��YH�M&������g�'#H>c��'{wl�HFh�#i܈�T#C�WP(��'*��[H"�'?��'��U��N�X�[���
t�s�6
��듮?�1%UtxJ��<�~r��";����BK�r����t7�N�x�����Odʓ��*O���O$!R4䃕7����-�4��%��ō����y%t#�y��	�OvX�U�3"v�w�E1wuDq�P�u��쟤���lr�D�����'w�O� M�p%"�lx��Ӯ=��x�p�[̓k4�j���$�'�b�O��qW�́Պ9��H�bJbUC�i��� d�I����	����=1VKM5�N�Y�j6U�z`,P��r,Тr�J^~R�'��Q�D���d[�U���H1R9P�مxp�(ǭAyr�'b�'�O����Q�,�*�E]�(�xՄ�~n�\��-�m���П���nyR�'�
�	#՟Șɀ�]7(���b@�AǼ�@üi"�'42���O�mb��ҌM��v)Y�N�� �X?*������$�O���<���yź=�/�R�I�0?�T!3�Brܐ'��)��7��O��|�I�
�z��կ#��L�v��� �a��5�qDA#����'��Iȟ��{�d�'(2�O����fʓ�FV^իuI�<~`P��3�Iϟ�@��T�0=�b��Y1fY"ᔍ��8�lq��m�Ly��W8�7��Ot���O���t}ZwV�$�g�NoN��r�	Y����4�?!��:�JY���ԸOSH�bB�.���ڳ4�N}���j��]�6m�O"��O����A}�Y�\br�?&���*�8f��4�$�ݞ�M �H�<)O>��$�'��02���8n��i���\� �rӪ���O"�$�h�\�'n�	��$��9��= ��2�p�*vԟ_SB%nZ��H��1.:�93�@m����?���ݼ-��8�R�S$}�H=��I4y���'#xa�$ �>+O��$�<	���T
S<*w������4!�~Ěb*�N}�#
3�y�S����şL��Ny�
G�WEr�s��W�,�3�
Ǥ����K�>�-O��ĵ<���?���D���R�P"g�4�)���:!�xF�N�<I.O��d�O���<	��[���iISMpH#�ʐ�=;,�k�+�&5��Z�h��oy��'���'�8�z�'��8�퓁'�2����<?�r%���oӰ���Oh���O˓E��d�s\?�i��:1�F�M���b̗���ƙ�M������On�d�O�!��6O���������%m��5"�(c�2Y�@|�|���O�˓k���W]?-�I��T� k*��"`K
G�� "�Š=6�OP��O�d)Gh�|�����k����	"�Ģ3)8�M*O�l"���ݦ���ҟ����?9��O�	+s{��V�h�t9CE��v�'�B+��y�|"�	O-D [�aےOƖTjU&T%�����!dl>6��OJ���O��G}�Z��!��ū0���6���Z�D!��>�MC��J�<�O>a���'�� �\\��F�Q}�V��C�X�Ms��?�K�$)K�\���'���O��E�%1��a,Q\P�2�i��'���J�����O��D�O@3T	ߍ;:tY�����X$/�����5xЊM<����?)M>���*؋�`�+&.4���#��J:�U�'�ba(�'��	ğ��	󟐗'�P&(K.�pM���=Ul8�fP�bz�O&�d�O֒O$�D�O�4�/�0LE����'#}��L�.ٸ��O:��O���O
˧@������5�bD�K���pA�'^���Z��Y$��D�O��5�d�O��D\�^��D֥=c���螸o�r�Bs����p�'�r�' T���weV4��'k����?��d	S	h	f!��i��|r�'�rG��yr�>�"��9� D���W$I{�nßD��oy���f�����$�����֒T��R�'�xJ��`�Z�i�l�ڟx+��v�p'����F�<�e���<�i�jX�KT�mZPyԓQ4$6�Q���'���,"?y��1Z��u�S ����ՃD�����������]���$�x�}:׍P�_�Æ�ˠu6h\�AC������"�M����?�����dP�4�@M���q+��=Dl �m�7)L:���v��c��]�X�I*}[|��T�U�6<3�×@�L1޴�?A��?Yr䓙UűOT�D���Z�甮Y�I�!/9/����u���Opej�:O�SƟ��[Z!g�yh0�i��ؽ8ܨ�N��a�	�YOL��O<����?yI>��1��8�OW��b�����?l���'�5y5�|��'�2�'��	08�� �F��!v��3af31�yQDD��ē�?������?��IfP����:A�Ъr`� � )�a�Q�?	(Ov�d�O���<�B1ju�IO ����&���&p�����;]����x�I@����|�	�9&�U[P��5�I2t>Q��Ǒ�x���'H��'�rP��[$nϝ�ħT2LӃ�Ԛ7�8�Z��
��01ְi�|r�'�Ӏ�y2�>	����t�,Ըs�{��Q�R�QǦ���՟\�'5��`"?��O��ɛ�2�n@A',0#�����S�:>d$���	���S͟'�x�'u7(  �K���Ii� )��-lZEy�"�*7�F6��B��'��4$?!��A3pL&lдƜ�T�E�k�A}"�'`�4���'��P�b?Q�3MW
\�hx��M*��!�g`��(
�a�O"�$�O�������O˧N�j��K�:$� %[�l=��I��iXȄ���$:�� ���� @��1���t�D�UH�M���?���) tP��?i*���D��d�iٟJ�Ȑ`&��N�\WL��'��ॣ.��O��d�O2-w�U�� �F��>��1j�������Xv 	ܴ�?A���?��0���>��I0F���фҕ|��qd�Y|}BC���'G��'�"�'�"k
���{ 
�Z�!����ĵ�a�'���'k�'�'j�'u�� �q�3�-t�*QOԚDj`YHa�܄B�,�O(4S#�է5�������YN6=; @6?N`�c΍'5�4��)�'�F���F^{�:b�ȨG˖��P�N�zX��`W��?�Q��(�-@)B	�Ү��/ޞ��  :�I�oM�l8p-Gdz1"�~O�,Y�é�Jd�f��(+�bh���f��
��S������U�"IA!���v �����2�������"`\�G�\�#��}S�������D�-X0�p�
�Jnɨ�I�VP�]q�DVF%~@ �� �\	��Bۊ2�Dk��
�]��d�/\�'�9K"��$�_�v���O2��g��=kΡ�tɋj@����� |C6T�S�|�C��r��ők͂%H��(�!r��?"Nܰ��O>@f�����[?B�9x��EO�ɜ�Ί���c�tI򰁔�8��<�@i���PG�T�'�^PłU�0L��ݺ�U��'�h(K�Z��~����]�ۘt8ÓA/����S��w
u�Rn�
u���Bͯ�M���?Y��'\�\�kW��?���?��Ӽ��������c��e���˥�w��xrMǨn\&���^;R�< ����#h��͓M���gA�/_Ed��T�̋r�~	��n�:Jx6��&Bv������Cܧb�0�Ml��z�%���~�*&��K��M����� �'�J}���|���3Y=Bx��&Nh�T� c�"c�!��V=\��� W��z������va�	��HO���O�ʓZ��}H��t�e�׏u���TO�1�U����?��?q����d�O��S�R~d��'��w�<u0��ތ	��9��+j1�q{&h%56Q� ��]�����剉j+�m qg���d)��M�j��r Y�9��i`�ڊi�k�60�x�Qr�ɜ$Wzh����,��Pf���G�H����O<�8ړ��'�8e�)]2�~�X�LGr�}#�'�p���@�^����^�qٶY�y2�aӰ�D�<��f@b����z4�U!y�����|�� ��%���T��.t��	ğl�'Qu@l��A
O�`���#�2p��)1�'P�<s�)N�	�D���
5*B�KF� ʓL�
C/��4) ���؞X�а�	A�X6^��V s�֤���V]�����%(ʓoZ�����l�'����K!�U*M ��y�yb�'c���#wd�{�/U�'l�,��'�t6-�- x�k^�;��u�j�9��$�<��F1Rg��OT2Z>=;�C��ě�N�sC��a��J݊�A]��d�I>� (�P�[8D�!��-@CB=H⮐�1p�ٖON�t֣@���A)eH��J6��:O�D��]�F����j����)�)��a��?eA�CrD"	Ш��1�TȚr�=}R�Q9�?���h����ŉGE�a,���Ε w��%��"O0peg09����-�+������'~"=1U� YK*M{h��j��}���1T4�6�'R�'�H�&������'�R��y׈��x���\bb�Q�l7p�(C���0+f������h���r��I\�.��'�>)1�!��`��Q���(^}��(��bq�}x�KU?:�ĵ:% Ѭ��O��9c�n��<!6*PMB@�1�oX?��ʑ+��F�<��Ȗȟ��?��?	�!������g��n�Z��e�<�*�-5`���"]�!&��H~��7�hb���'�剓	��hi���q�ը��;O�pa��Dp���	ß��	şPaZwrb�'�)M0a���fDB"I���$dJ'5����g�m+��ԎZl����y�\����lv�8�3��������9^,�`��?~r j���2i8��L;�����Ț�t8Z%���c۬xcFOհETJՒ��')��d��xв]I���w�ލ4��7&e!�$��{j~�kt��3��i��;O�1O�PnZ~�Ʉv���ش�?���Pu�'�(l;8�I�K'd؀���?!�o�?!����T.3@�X���
8"�-��wٰ3Kf�(��2	��j�X��!�����Ey�I�T��(�s��X��9��	^�:DaǞ>[���f�$�L���cøy}�TDy�J��?	J>y�I�;ht��� ̄�]z��Yr�HN�<aU(���%�f�K�Hua��U<���iq,)��]@)~ yc_�\2�1�y�J#J<�7M�OL�$�|r�iê�?Ѳ��`N�t	�j]�M�53���+�?	��h�E�d��S�P8�V�g)��8���)$�:,�"����B m�����۾{����3�>Qqܮ}��ݹ�@ؘ9�H�1�MTڭ��i;���E	���� 5F{�]�iVp��?j�"���NQ�6Lk� �/�j���P�!��ߘ ;X1l�� ����m͒Q�ax2m7ғF���Kf�nI[����>���Kp�iV����lZ:�����՟�����i��@pfO�v6�P��ډez%H��7Gl�S���0��M�Uxb>�O�)��9\�J̊�M��\�2m
��eN���O X��oӌ���v1>X�VJ��S�	c�CQ'a�.�s�y��Q'�?�}&�$�w�	�A�0T��I/ �0q� J0D����+8�� �� L���Â#?1��i>&�|Q����.��C%AZ�u�X[U���0m$@�Џ�����I���	�uW�'��<�L�#lKLl��&X
^��8Cb��J����J7N1q�#<O8��� j����ąu�6�UɎ�.HhA��'J�Y���Y���	o�0D�牸[���A��i�����LQ�?�����O��ɑp�(���4(�xi3�*�85�C�!d1��ڲ�E��-��WM��b����4��c@����iB��'�0-j���
V�tς�W�>����'��B	�L���'��	`L������F����d4-2�$Ճx{�zr	�",^�x�,��f(miFM%}r�:<wJ��q�ٮ.�r�:A��p<���؟��I<�֣�Xj�A�@N�Vt4|�6��l�<��H�I�D�8!&ڀVO�dc���h<	b�i�~�ab�-��K$��%k�4�ⳟ|�-U0Z�66-�O"���|��]�?i3�ֶ
��e�Ëמuuހ����?���6��]x��혧�ԓaM�:���)W�e��,��.}"J=�O�"���Mڌj�q(�',\E���Ֆ>��O埈�<�*��G�W�����Y� C�I2G��T�<i%G�X�A�j�}|���Gd�R��k���΂[ڀJ��S4O��Kgi�0EA�(n۟����$�,ɜu�����,�I֟��/3�1JԯV0���� ��<D0D3S�r��)��iD�X�Qߘ��?��"dɽ-�8����F�z����.\�qm�:��2�V4����7Cfj�j�U���p��	%�l���iUJ�_�H�i>���C�� �����`	8T�z8P@���J!N��ȓ�r���;{p��nТ5Xy�'�#=���ixP����)_> &�<j/F�|a�t��#8Uz�͹�d���T�����ɽ��	�O��S>	�8���B $L�)���u�ň�� _��8��'Ӭq��-̤<I���惄n-<4{`��#V�� s`b�L���T@�)�ӄ6OQ�Qu�=���bG�ҟ�	��X��hy�'�Ox=Rq�G
>�q���l��q"OL�c�BH ��բ&��w���R�D��m�	Uy"-X:6-�O �d[�K]dL`���0]:P!(Ӊ�!m4�D�Op(wc�Ol�D>Q#��BZ����i� MP��BX<~�Q��@�:A��ITKvRhQ�&�r�Q�LQ�)L
,~ �W�@r���Wai�	S��+)& �BHÂX�zu��`Ӫ�Q��
a��O($���,(nG��c`_�*	��8"0D�H�`Ǝ?@�J�C�g���b!��ߴ&=s�H֓�� ��	�I�x�#H>asd�NT���'��Q>��0�ß�KTJW5aZ�x E�B
M�A������3#?\A(�f��9MeZ��Z�<�O���D�L����(<x�k@�	
.B��'�@c�`�
VTʴe���h�Np�GU�xq(C�ی6cXI+G�>��P����<�
6i��x8���d78$a�e�B�<k�^ª!���> �mPA*w���d^�D?��{���k���jR���pI�an����������3n�d����l�����ݰV�V�i�	��|d$�	5�G7j���B�/���')��Q�!�|��W�`	J$�<4���M�sz�=2i�=p���[b�[�/�F5J�����^������R$��C��H׽Y&�-Z��D"��L>��КR<�����.r�e�c�<	1��Q�1�qi1v�xQ:$�J~b-��|jO>!C%3�J1���,8�re���R���BK_�?I��?��4q�.�O���q>�{��9|�f]8��I�/�^�	o+@��4�[�s(B���I�4�E2j�?~��!U���F���f��8��5����e�Z�w)�& ��p��?p@Mæ�.��e�B�ې��y*�o�O����ġsX�7��Zi�葏2�!���n]�|:D�@I�M���3]�1Ok�iO�'�Vr��eӊ���O��X���b1����!8�(����O^��Q `��d�O���6s�%`dW8(W8���l����bR�5Na���$ N�вL�P�'R�d�I��_Y�PA6��:]-hi�.7���zS�M�P��}�5i/vџ4�k�OL�O����*�FlN�ȁ8j��U"Otg��$+� �&�	��Dı O��n8R�P�O�(��JV(��%�:�'�4��� 1�M[��?�/��9*I�O{G$5,T�i��E$# މ� ��Or�DX_5�AR ���
D&�. F��O��(:��h�P1c�tJ�ƻ��'k�ȗL @Oh�h6�	3��#�����ޅ��� ����AW�N]�BP���f�S��3�viv$��*=����8h^��ȓ]��#�{��)��1p�$��I��HO8����U!CN�S�h��E�撚�	�4�� +d��7�P韴�	ӟH�iމ*q
J5P	�e��+|��YRb���!�g�DҦ��lڭ˵���ḩ��
 -�uk4KI�͙e�F�g�(��ԇo�*�3f��i]��Y�A�Zܧ��S�? .!kF�U��e���vD���9�IvL���|�N3NR���5�ޣs����˧�y�_7| �P�b^��(�I!��$�^�����|�%�������V�V) � �+��[ۢ��b�:���'���'������D���|�@�G�^cH�����[�r8�� �.�b%��}�E;�&�$h�q#3�I'A�� �5�Pm<�&��'��As	��}[�e�!˥m,��I���?A&gɃ�V%��h�2\��Y1G�v�<Y��оP�S���0��
g�y_�Ovxڀ����-�Iߟ�jQ�W	D� 1�q+=#.FY`�����	{�����ӟhΧg��Q���I�4ʉ�4��	��dRB���j���DjJ�Op�D�ֱVIR �fC_A<��*�'�R%i������B�N4?��l�$�$DA��Tu(��EA�8h�䩂�w��A���+��vc[	~�i(E��"6��A��S�'�0$�#�c�x���O�'[� ���z��	Y��O8h�n�b�&F�J�D�����?	[6�?��y*�����V�hE�$V"j%!���*�(�'�dk�����Z��{E�H88�໖l�y�spP�I���S��Ʌ�"_0�iPc�YDI��]�<1o��EZr!����f`�i�Kb��)��
=����1���x�#�\���m�ԟ���ߟ��Bm�Q:I�����	��5X]^!z�*��0�Z��E��-j���b9}�o͠i�D@���L>i��O�.�A�ϖ#|���"� =�O.�1bC�����$�L!K���Z(�lˇ;�*T
�ybK��?�}&�(��<7ir�+G�����cP�1D��+���0vk��#C�>ߠ��w�/?�u�)�'Ws��-�~4�"/��6���9U�C*�����?I���?q�����O�擝5��T��h\`�6��l�o��i&m�<~�
�L��I�.��կ�
R�">�h,l.����f��*�`������`��}.��2B��Ҳ�G�M��#>��`W$b]�A�eGB�2�s���#[s,��	�Ms��?1���?	��?Q���i½D?��Q����[����?p�!��Ćxv���v�τS/�2&��/v|1O 1�'���8A x�ߴ�?��}�5���/9�;%Gǿm%n4���?q���2�?�������4�?iM>I G�Y �S*Q�9j��_X8�t	�0������ōāS"0)s�ł}"����62�|�²m����S%V)z��t�1�ǜ�yr��-3x�+�f�
y���p����x�K|Ӧp�+�U�j�s$��,-���E�䝮���m��T�Id��L�T����>��9yeU,4h���H8<���'A�y#@�'�1O�3?���>E�l)0�%�,Dls7J@���-H��?���͎Tc �p*� #��)J>}aT��?y�y��T�
z՚��k��L+�y�h�?��a['��}c�=�0<)s鉍Q*�!+�Z�%��@�Z	��ٴ�?!��?� +	�p+��?���?�;_ mPA�@)
(,�bN�w"�C6֓"c�"r�\P8�QseZ�ߘOm�'�~��IE�J��C )��h�y�k����d�'>��t�ը� ��O�'�|���GߧP�Gᔈn�T�P�'��'J��&�����D�O�i��i�cC�A�b��r0�<2Am84�D�ʎ8�NQ��Z#�2H
��8?Y��I#)��ģ<)�(Ȗ(��Y#�ĵ:Tд��-`�V�#���?y���?���/7�.�OJ��w>�"&��!AL`�B�Ў%��@�>��B�	�v �PÃF�S��IR+O�R':P���&�L��
"u�1��,��Ԡp�(x[���$�O�ж�\5[�
�����?~l0�"O�����~��y�U�d�4�#���|�Co�0�2�i���'��i��k�-!���p,>M>@Q�'��ᑼr�'��T6=yґ|"�z��Y�V�u�LX���D�p<ɕ�R��m숋���!q�1�͒�;z��I�A����v�I�9�U8��[o�J���印��B�[�x���% �T���7ؚB�I��M�b%�P(R! Q,@�Tq��J�M�~f�%��ikr�'�5�t��	'.\�R�}n����_�� X����@#aП0�<����ǭ?��f����D��cNUx�BB�Gx���fO���X�*�.?F~��fj֜��_~���3�)�3� :��'�&-t�E0&f�>��P�"O�TjEb��(p��7F����t�'Ĳ"=�%ϊ.h�����'q�|:e(ɃXs���'���'e��3�F�[���'.R��y��Ȟ.v��ԉP%%�hyd��y}1O�'�'z��C%�.A+��@�L�m4h3�{r��-�0=)�Iߝ��ء�.�'�KGV̓$��)�3���<Ǧ@yᣝ�/�����@�*�!��ֱe4^(���{�H �� X00��	��HO>�z @J�5�q�V�՗^��aXD.�x|x�E_ǟ��	ԟP���ug�'g3��\8�JZ=~����G�Q�
���m�!��`�`�kE�/�.xM��Y��ؚ�On�``�J^���!B/�� EE)d��'�~tʐ�Ry����U�Y�ĽA�'�.����Z-��c�-G2N7��y2�8���%�r�8�4�?�� G�-�ƠϦqH i)D�L�j�`H��?�����?������D½�?yL>�w�\*���T�G�9*����_8�XK�F?��)8Q�����%r�A��})��� �7_�l$��Xp%Z�k�e�1�h�!/;,�!�DZA����U�ߛ,ݬ5�D�S>1�!�妱�6��~+��W�M�bO�5�R�7�	CF��޴�?a���)V$]����� m�ձ���?>Q����D0TN����O����C�OLb��g~���L0ȹV�u�(�r�����ɾ�"#<E���D b� YU�b"�̨S �I�D�,$�B���Lh����Z t�{r�Nv!�DХ]�p�R��^MQK Xaxr,*�W�����n��ܛ�C��M���iPR�'{���{���(�'2�'��wZ��!�ֵ�+�6��ɧAů��'�v��ϓk�6�q�lĶv�\�q�
CKy�=� ��xx�`�䂗�$��i @�ӆY�XXQ�T�Z�XH�)�3���f � �:Y5�l�@k!�"O�\ e��=���[bA�#d�&��'��̈���=Vq�,xc�݆-��c"�<J8�i!F
N�9�i�I����ҟp_w��'��i�2cv�����lFЛG��/a�B��vO�)�ELS�b0ReR�`�}�(q4�^:i�!�S�b�� w�1[�l%Z @'9Ǹ���'����D�{���QDQ�a��YҀL�-�!�$� v�RY��f]?<?�A�6a��^�1O~��>AČ����'�B�g���rGԃh�L ����	\b�'K�@���'��3��-���'��']�I��dՁV�<
Wl�w	+�B8��C�0�I x�p����]?=�|}�u�2J���Vw�B�7��40��iS9Y�1C �Z�w�!�a�� ����S�H�k��'!�D\�5)���'H;<���m��{�N-���#�	�� �ݴ�?�����	r��$P1���Ů�9`d�]p��{����Oجze��P���ɿ<i+��ʧk�
�#@]�J��1����8moL�O�}zAC��B�P��+�2�<
�Oܥ?r����l(�@�o��Y�F�o�\�A��>��nM����4���'� ���@�Y��"3#�>)�j��D�O�=�+O��z�#T�ܼ�SS!!��2�'^�6͈���&���ʜb�p�Xp+ �<Wb}�](A�4�?����?�s�Y�s��m���?����?��;&�=���\=bFf�c�H��4u:�y������<!u+�4vf+M�?�v���X�qO�1A�'Ì}��M˧x�l#w%Z>
�Xs���Z?
��L>9t���T�(W,ȸg����j�t�<�b���u)��۷%^М��	Dh~��,�S�O�0��T*ݧXK�5���\�e���b�/��Rz<����'r�'��
}��	��\��>Yֈ�R"�5"�����׼m΂x���6��Xbà|�u���\� �#a!F��Hё�E�d�(t��\��.y��!��Jp��Y�#�i�'��9��oQ�/ax�#�ˏ�U�7��?YG�iu�'�B�'��'��P3�����)Rl뤀��N���"�ɣ�yRÌ�_E���&F�o��!C�/�2%�Ot�'���=|	�ݴ�?���X�ĩyB��qxF �`�ړl8֭����?�֋O��?����4'�]��{c����ߥ[JLp�!J�9ZDL�3n�3��x���3?�``hB�
�*�$��
D�������eDD�P)��!�H[7JߗsASub;�	F�\�de��,6��V�9Ju�]��'�ZC�)� !��NK:k�vE�Ս�#k ���O��o�j|�	fh�Vڄ��G��,neNc� �4�B��M���?a.�^�A�J�OV��U��m��R�A�ک���O���Ҥ�>��=�|�'P`���o�"L�B�Z�t��KI����:�S�'c�r�A�9F:I�j��V2��O�|���',2������ L@4$kf��"��[��@���'���'��0�wD::#u����M�JH
�\���x [�cH��@v�B�8L�����M���?!��Tޒu�[��?����?��Ӽ�&J;N�uL8F8��&F���'�8 ϓb�:	�E�H7δ�CE�=�bm�=��oZx���B���� T	��t�.�Ǣ�e�w�.�)�3�d�/H�Q���(`���T���Q4!�D�
M���� ����X��,H�z����HO>�`WA��+e^P6��	Zv�� ��k����C��$���X�	>�u��'Cr?� �C� �"2.z��Ȟ]c���J'gi �#d�(=@FxH�`<<O�!BQ���HZr��	+���x��ڱW\pbI�S P$c$i"<OL��I9Wb�I��ȮC\�(M̻O�26�OZL�BnL�:�ԁ�A
9�B�qT"OրH��~�1��N�~n�=q�d�h�YBx+4�i�B�'#6���_$Oɪ����Z��-:��'<RR�zs��'=��?y�"�|2���6}z"r��[\�	�1F��p<���X��(����ōJ��P�CB�{�a���52 �ćI�I�V�δX3��_QxU���N�b��B�	�E�,1�&�Y�,�3/́4;lB��<�M3�
�M����ޮ$'r̓S�
<H �i�2�'���Z��1���F�Hii�-M(� ;�HӘ1n����Ο$�rd럈�<������.��4�S������H�%k��Pb2�Gx���%��|�0��୕)s�r��C���*Q����N�)�S�C�2b����gװԥ��v�!�d�$H� HXTL��1��
���>�ax�=ғ>�x=�%�$��������"옣�i���'�h�A����'Cr�'��w�f�#5��_o������j�`��D_\��y2���q��(k���"�XK�k���'Lr��ϓ)�f���;Vo6�0t"�?lM胚|���?�}&�0����_)�AT��Jl�2.D�X(1�+\M�I�mC�#�Dˤ�+?�e�)�'|>j�Jw 
9�!X®��:.ah��6�A��?���?��q��O��di>�(g	C�0�-A��8�sL��'(�41���v��t� �ɇ�8����tdQ��1��M�0�Y�Z��}ҧ^ Rr�Q�i8����S'~6(hzGJ�.vL�b�#V���@	Y&t#����)v�E b�Ola��	�0	$�y�A(Pd~H3�!�����:�D�`�Ȅ	U�0(1���3���B�y��hӠ�O�1kDBVѦi�I�a$�8b�Mc�-���ػ��Uǟ<�ɻD�(��	����'-JĎF�!�lLC�Q�q��b��ڟY���P%օ.�\�g0p�l-�O4ʓN��]�#���#��G��-�	58$ŀGGQ@�t!R�:��ʰD=�O���ɹ�ēE|&<�%�B�	e�c�%Ls�!�����TɋC ,i�UƊ�gS�Fx��i>�S�4k1��҃�>���A��9(.�����s����ҋ�U�g�6j��90�9D�x!�)͚o ��e�ɬ�j<���8D���A��VV�R���'.�64B��6D��9�y޲��7�����1�d3D�l��*�ޕcd`ML�4�!3D�z�F�-k~5���\�;,Ňȓ*� p�%���=�笄�.���ȓ�@S4��:)M�u
s�Q�7�J���G���͏l5��  ��Q0B���ҧJG0��!��U	h}�ȓ\�2̻1�?B�>��v�� �&x��X�@pa��4G$���,�����l��a���{Y�X)e�8:�0]��=n��V-�)D�h���-��r��%�ȓq���iu`ӳ6R)8!i�--zy�ȓF,�q�V��4Έ���Xsr����S�? ����'B&;2��ȕ�]
� 
"O�z�oC�S@�x��^��!&"O�su�K�{ਅa�BC��{V"O����> �J�qe�S�H�l� �"Oҹ �J�4�"�I�E8*\c"Oԉ�-�=X�P�P54
xڳ"O��S��0E�F0�#���@<�Zp"O�Q�'���ڡ!���R��2"O�u)*!K�d;7��~��*g"O(��@�I�mW�h�7��`�m
�"O�|RS`X=K���q+��;P�mq�"ORȧGAx�*���2D�u"V"OQX�a��$n�ɨsh�CR�"""O�d+�`��yTĂ����^��P"O|���̅O@�R3��8� <��"O��H���~G�����Ӥ�蹊$"O��Io���A�E(;��w"O��Sv�6t��D3Fa�43Rt "O�xE��gdɻ� ���q*�"O���F�
`I�p��X9'\Jy�u"O*ˇ(ډ]�����(4Q�� �Py"�<h[�0ٜW��x`���E�<i�(\	�ZQ'�^�<y���r�
M�<a�%^ �X� ׿<�4�PH�<֢ė
M�XG9l`4�U$QC�<1a÷Y_9&�G3����#@@�<�B��+�da�4�33��%
}ܓY���8U
�\G�T6H���0�G�2����y��<~���HI w�`�j�mO4o~�����.l�I�}QT#|�'$�!�B1ZBB�����Q����DhQJ�6�BEkC)'��}��&Z0~�t��g�y�8\)�ͧ��/Y(�v�����3f��v�X�%��x�a��^n�	�|�`��t!�<=�=vΜ!Yn�I?K2�o�?�����#'��@��� 55���ª-�O�՚�vnj���c@�J��AõcśH2�A �>�yb@�V���'X���cc@���a��O��@�z��P�۷;�
6ǎ�;O6��S�M�O��+����/��L!d�=c����<9��U�\P`�A�^f�ƴw�g�L�� �Z|�dbBg\�17p�;��E��Pa�E�Nd̓�j��4f!�e��N^�qS�Iۅ�v17��PC��Z#��؟�s�0J�$�1z���6Gk>y�qI	u�`�q�R?I����R��'\��S�O^?8�Ӥk*LO2Ő%��c>�3��X|��*�,�O��;�;O�ՂS�Q�FF"�Х�?1����\�ę�,�h������T��BO�R�a|���P�r��b�H�Ӧ���ɘ��RMq��B�2�)�e�)=�i� �4�y�-��ug�O�)	�D��l�4Wr R���76��,���4d妑����?v,B  �+�d[4b�k�4��gb�kq(�������&����&��Rr����f1� O��w9�x��O����<	��#���{�T7���.�0�
��;�9c�EUw���`��<��ߛ3�ZU�o�.J� �ΓY�,$���YꀀJ��hVX�!�R�ML�ᒡ�PVjp��I�7���W��&I�dpa�M
rab�x�iz�H�J[�b�.G�3��*��鯻�~��ޮ-�|t��
� ���p�T$�0>Y�M�-28:�g�4L�씀R�˸a��af������_+l����')6Y�[w~��T8?@f�A!�+�0��WJV7(�=id��9:%C4�Z�67�T��*�@9V�G�(uH�`r���"U�mo`�c����^� ��x]���r�B�� ����$Ŵ38�8GC]�1O�1yL�2h$|+5�����D�W@TaNӕ�8��� +:��D�R�4]k��
���'4O^�`��ƆQ/�Tp�ͣY;��x�Y��Z�F����L�2�az����`�L�(��:0�=!d��\x��'�� ���3NxX������ǳ#��΢�`��I�j&�!�LJ	���	I&�OJ1"g^:� �Cd��&�F�� �����S"Ŗ���bNV還���2Ib��pRiPF�4�&H�B���c ����-�'�:�;%
��z$Fx�)B�O����J2C��t�s(Z4�yr���l��X�	0�A�T��N(��f-�$H��:�u@�h�+a&pB�,��0Y�<�R���]�ܐ��HP C�(��& Z�i�͙�;X$0��B;/��$ϓiܑ��@@@̓,;�|Y�D֦c|l�Q$ǅ��˶kٷE�dl8
�x9��y��YP׾����FK܈�����<A��JXU�XF|�`�;�y�c_8`k�*�u-��`@/E��0>iED#:�r,�'�Z})���6VGj���J�&���E{b���Jh"��űZ�x�����~�
��a�Vi�U���]�08�
��OV@SǄ0C���D-;Act���� �%x��(�C�5w�`k2��JB�XP�����]q#�Vx�� �\Q,æh0�Ɲ�'���k!�إQE2m�(���z�`��V"ax��"}�V:�aѾ'?�)P��	��y��1/�d���Y�F��C��/�`1�'���03"�?z�|ΧW�2Q�"Aѭw�AX��)
���"�?�p>!BCL�`�IRp��)3r�+�H#f��=��Ϛ	C�p��6+G�a�5`���s������C+#2r�!�1Ö8�O�	�ą	�L@���L�#wZ����=Ò`[�,O�!�DS �Q�W�l�F݋P��Q� �EC3`��S�W�,&F܉P��֝�?��MH"��`ZL�q�灼Fk`C�	��� @QNX�)[Hm�7���R�xD� Te������6>�I(�)�<�}�;ةX�C@V�<��f���_~��9Vr}��"6��1b'!My�$ԋ��U"��+b�|��EW>�)f%	6��E��ER�ȸ'-4��2K��F�։�fڽE�|p ��D�?n`ZiJ�m�%M�w'ܔ;D��2On��q��YnQ3����.xN���FZ�HMÕ�C�M�דc�`h��C�T-8�Z$"T9 �F->�K�Θ�sю�A*R�#b�a��V��&�`�5�J7#��񘢨E�M��[�L	H�<Q���!u��$�W�נK��$e�8P5�E��?�F�0�ē?
�p��!� ���wY$L�&�\$��k`�O0�I:�C��3!D¡L�&Y8�� -�!2p�Q'<�(��%kԈS)���P0QCƈQ'R¥-S��4�=��n��B�d)C0�����8�p�a�'��!9b��2M4�Q�lV-M���s�����2��6��1��p�J-c@�,Ӑ�j��9s���ä�R��4;�DH�Tƶm�2m
�K�ę���L�c�E
�d�$�]X�<c&�3rM)�-��-ۤM����syZc�j��$đ�}�&	���Bp��0K�'�r�BL/����çLi��$�jd@�󵍈�y6�}yf̌���DT[���c�|��*'�bD� ͜?!�\��&A�4�0>��Fm:6���m�#L��Kpf�9(��
�nL8n�,��M�D�6�хJۍ`nƅ�
ϓl��4�M�k�h(Q��B�/e��Gx��7H���eP�T��S����f��a��]\]x�h���6�Գa� !��S�O��qwL<t��t��kŪ�8�k�eP/t� �aV�ls֭Y4��&ۆ�ssD4P1��.V�T�єeG��b�բ
n!�*R�Z�ڒ�� �,��kL3����Miށ�`Π?�Ƶ3��1��XNt;s-P�`��㠠�,$�̅�	7e%d��`O(/��8�Ι`M�u`%\ z�J����@�3���
��$��9j1�<}��R0k�Dxb�͠A��3Tb%|z�py���DG�C�&���n�>6����uQ	�y�GTxw8d�aF�;/xF�:%h��y�Bnd���oT����!�N�X@G*�v��ĥTPC�B� C�LD�C �%��)R�5���pC�����a����1!� =ĕj�D�A�� �Wa D����CL�l6p��B&8��,��>D�pb�Z�N^�		1,_=uϞ8R'D�����<yh����%�"���!"D�䰂��>f6,��E��=��?D�4 u�D�WM�0�e�:ȍi�H*D����GO���0#���~ʠ{�G(D��V��)@^��IV 
����㴦2D����ȒS咵��m��o����2D�`2�ŝ�?�¹�a���0xra/D�� �kF�Z��ԳAŭ#��)8�#+D�0�c[I���!�� irmR(5D�<�ADR%M�|�c�A��b�t�ʲg8D� kR �C����v�RI�]1� 6D�\��Ôkt��`2aۀ|�J�S��3D�x ���
v ���&.D�%G̥q�6D���E�#�������K�Yp��3D��3Ch� �̴�d���z�x�p �2D�hjZ A�]+�d�--Ӕ����/D�h(�*�����!�WF���q6+3D��p0L%;(��(d,BQ�p����$D�\�U�C0+t��F�)��B0D���4+f~��J��|���0D�@�ph]�s��&��4�,��/D���F����[p���\Q�i�U�/D����ܣ[ �y��ʚ mC�i)�`*D�� ��rB[?|`x�
ϵCǠ��"O2���A��X��r!C��A��AB�"OԐ�� z~@�z#�o� T��"O�D�%nW�}�l:�� �i�Qx�"O^�#��L-�(�!I�T60�q"Or�Z���Jg�<ّ"A7(H��s�"OT���לt��)��(9�C�"O�}+�	�#e�$Ls��8SyH)�6"O2����ڟy�mP�M:�$���"OLYBƎսvH�9Cː�\ܠ�2"OY�Z<%���1��E�i DQe"O���DM#L���D�Y�3���c�"O�逰��"v/���PjA<`�V��"OT�k��\ m�td���y�D�+�"O�����n%d��P��B�4��`"O&���bDh�����N�8��Uا"O9�)Ͻ���Z5ł8v�r�B'"O3c�B/S]X�5n�N��d��"O�@Rag��<�d�H�;#���"O� ��n$|s��9B�07"O�Y��.@�pqH!�)�Z�(m��"O2A�VU�h�r����	`�%�u"O6Ar��)w�-�mŽ;\�x�"Of,���':_������)N,h1�"O܌RU+O#H�TؓV`R8OH�A"O$���G~$��:HGV)�"O�,#�H!j�(��1�C-��p�"O�pd�E[0 ��AL�=S#�Xp"O���r��<a�䭑4�>U���XQ"O@�W)^��\���o�*A�
�zC"Op<n�q�8U;F�����"O����.�K�HY��ۘ����"Ot�	6D�
q���{`g���JG"O E��,QjX�A�g.�$Q�-1s"OX�!��*8x��IMS>�TY��"O�d��aR�+j�kAj��_�����"O�)�v�ɸk#^X����:�4��"OZ�P%��7P�['���w"O�|P'hY�Ha����@ڜr�\�X4"O�U���*l���Î�$��  "OJ�9a��e�4ص��&l~@ �"O���B#��Y��`��*H8�aB�"O�0C6�+�x����aYZ�j�"O*�2Nȴ\$
\bF`
�P=�)"#"OX�!�(��XR6u�oO)t��"Oܨx���m_�dP0�����gH&D�����E�rWrU뱧L�6H���%D��xCaďt�F� �cʹn�H]��>D��[4��
Z�qCa��@g(��?D� �0i˓m�^eh�#re� �'L<D����#�IG
�j�&�7g���h'D��	��_�|�u�gfX6K�8	F$D�����̨=��7��#D��
u�"D��sB"[�M����!��/[��@pG-D�xi��ðnl��Bb&�V��� +D�XJ����U��æ���dK ԉu@<D��i��ўT�^8K�b�B��Fe;D����ǘ�����-&ԡ��F;D��ȗ�֔]�n���.��s3�:D��qщ�M<@�3հ���-7D��{���̱�ϐS@�P!5G(D� �p�E�^��A�썂WR���d�*D�|�a�ƹ> ��C�	؇G�>$
&�*D�8���u�B�	 A�8a�s"*D�� 2dz%����j�h$c�J�w"O�P�dD
sI�ݛ�(V0��'"O0�h�-\�h�H�⇡�3���"OЙi"gǌkm�3"��M����&"O>x9�K+B���D��(�
��E"O�A���"rJȉR��ܖ?(�K�"Or��rJӇj��]�S��&�V��a"OP%s��O��4y�#�e�v�iU"O�("�p����b��8uݞ,;S"O�����Z
a�*�@�#�&�^�h�"O��¦AF;"U����#���B�"O��ɐ����8�ci7ܪ�HT"O>I��OU����G
7?8��cf"O��H�m۫/��JCݔR�t3�"O�tX���2 R�D)H
�"O:y�N -��&
��1�"O^�P6.9o�=��ä/��#�"O�8�F@/?���9橏*����V"O���W�R��T��	!h]t��R"O�E����pGz��І�<H<0 ��"O~[���;���&h@(^HTtaE"O���@J�+2R5k��ϙkEbM�a"O�1�*��|����(s,(�8c"O�(p$dG:V��oS���'"O����L�Z>�Z�nRJ���!�"O�Q��fO�xR%J׬�d��)I%"O����c��j��!�ضF�u�"O���Ώ�⾉@�i]"W���ʆ"O�Xs�W0D�S��Rr��]��"O��և�6� ��1(Sz���#�"O�p@�(,7����&Z5[��M*�"O�mPk�.@��kRf%����3"O� ��c�L�d�Zae��N���5"O�ڶ���_7���RB<q��h"Ol�8�O���BD�=��,x"O���5iQ�bl��i:ro� ap"O�@'n؅g�V��b[��q�"O�`��� z�!�"�#x��|y�"O��i��=`�A	U�L���"O ]��H_>8��ȓF�v�E�2�3|Ob7�H3��$�EKE#j ��S��'���9+�#��YB�G_������0D���a�ɑ� Aq�,�1��aY�J1�i�����	��S2��$�G�Yi���m�!�dW=�hɥ��2И@���aZ���fe�R�@�|�'u�t+G(�5�E��ȇ�I��'uҰ��&P,f��,p�	�L��x��M�4
�O�">I�Rnx*26�� ��
0'�Z�������$�?q�'ĄPr`:ULU1��)��y��'�ʷM��a����Q�7
��{���O���0�S�#L��Ō)����7!�(NB�	?|\�P¦�,I���b�	()�a���������+�P��A��JM���e�!�$�lTH�`�;`]ҠAA���o��F��|bEV �
m2�*̎�68�Х��p=�#)�ɍ+���V(װB|��)t^RC䉸Ce����D1	���V�/���d��#<y��	�� �c�h��}��"4hZB��?x-�Y�
%6Եa�Ь{�`�$ŌE;�"~��c$.�tE���(��Y�",��yR#�	ej�	y�j�M�B��
R5�7�&?9�:,�A�I|pI�MP�k�R��}3�A�ge�?dE6��E��LWdȅȓF�8���gB_��C2e�-�2U�>����� 2�ө¼{k��`J�x��S�"O�d��Cvن���K�Fln�i��OR���S��x��J�kȌq����N�Z��1*4�y�N�F_��`!���n9n�b�'ўb?QUoA�H5���2����� D�,Jf�Wm��Zӫ�*u�~��Q� D�mַJj�1��\(Y���$�<���v��%kۃP"T� I1z$"��ȓ>���@�[n׮�R�D��W�2���VNE!�ת �<���#R�(��C�}�Ձ[��5;w� [< ��@5�x���# ڠ ��F�W�)�ȓq����q 	>8I�X`Pa����ȓh���Ӧ�9�P�v˂�'@Zh��d]�+�8gb�ѓKȉ~|!����[s �6^|�1�6���{5x��'�ռ}r����T?&[L�ȓ)���2T(DP�#��g�bܗ'a~"@�7�6��³��I�S�V��y� �1�(��)k<x�K�%�yR��(#��!�C�^DݘM��y��n���c� ��Lsg�
�yRȔ6&l�,���Q�F�m#�/U�y���H��œ�k��.�B����y��#{��#�j�q`d��3C��y2
	����@�t��A����y�o
#g��U�u/�o�:�!3�!�y&�G*@-�FoN�[_(���C��yrf��PҎ�x�P�l]03A¯�y�a?Mc2,H�F[�<�1rR-ɣ�?��'l��s��{1�Ȳ#%�2�n�	�'t2�ѵ)ͮ��$1#�A4R�x���'m��p*�,��s�`D�G���c�}R�)�9S��1��ܿo�l�C'L�L !�$�p���A�p�|��L�d�!�$Z�-ĺ�h������#�.��0f!��ٮ�<@����,Tg���߫N!��G A*�#��B�u[b�����x�!��
δ/,T�2#�>Mihq3�`8D���2��Y�ژ�Ub��kB,7D���[3<H�4�6�mWƥ��3D���6�;(}�|�Pk��u҈�t�>�c��|�#��$�M�g��(�h��7�'D�(+�Ő<;S�@YP)J�ii��F�&D���sbU?s;($9#���@��l�p+#D��PW�L+���"��C2���;��#D��Jpμ:����� �"oh��W!D�A��I�ԁ`�ʝ\^�kg"$D� �L��e�%0EE�N�AcI'D�`��A�[5B��	�n��$8��0D�����
�s�t���(_8�H
/D�<c�/ǘg"8�$�gw��J9D�X8�J�|v�K#n�`�飡;D��ȵ�ȷZ��s��&.Ta�e�8D���wm�2?zuz�h�&�Je�X�Py��*H� 	��f��"�%�f�<�H�#Z��x!sK3�T�oCY�<q��WwR��p��J� ��`�<�D���ܔ��:�,�g�Y�<�f�a�p�1��~]�"��V�<��Bޘ���6F �&<����y�<Q%�C�P�"�h�GFz#HH7OM�<�1�4u��*���Cfa�g�~��$�<����(4l��b��^�<¡��v�<� Hh�GM�r!���V�_'�6(���Y���i�����	@��u�ڄo�!����<�j���O�����%۩^[!�dΰ"�Zذ�/�3�d	Ub�(Y�!��ӎu6Ģ]*�4�&�ħ�6m��'-h��Q)��J��Œ�C�R�N���'m֨���)f���`u/C�!�8�'0lrD���X?�1ɗ&�	Z���'�|�
��N1wۄ�)��)�����'v850�&St��@V4v�օ��'ڂ=�����,5LH`խL%v�6e��'��XPh�#$Hz���lO��2�'�
��D���]ĉ��k3"��'��вq�̵ x&�P��5� �
�'�4x(���q��x���Ņ9@f�9�'�d���,��`8�Ш̈�*.HL!�'���c�ɞ-�eɝX�X�Y�'䪴���U�$�@DST�޿~^���HH���̢2p"Y��hK�m0%��7�5�q�Ǖ}�as�
4�����.�Z�$D�vI�D�L>-ڲć�,T��+�v���ѭ�9@�	��9�X�7�Dq��H���5Ŗ���r&�����|����
�|Ѕȓ���!G#+L%�a��$�A�ȓ!V���cH��=N(�Q��ċ�f��yz�ujō$f3��;�ͶM�ȓb�5zF�O�����&�jZ���r�ظ@��3�H�pF���D�����?\0\�'F;r� �v���Up���ȓ@�hy��Y:��	U#��:�z���	zt��cOKW�|�E�O`�F��t��ߟ1����/ˀ;ZLȆȓ>��Q��M�@���2�_65�����#2�S���l�L�4���p��<�ȓ9�t�`X�6ܺ�p&�=i�&���sw���ш0��ThF�%T䈆ȓ@!TY[gd߭V�x��S ��K�Ҍ�ȓj"��R ���[����`��,'~1��dSv�2�M�)/=`�(��!b��`��$��T�4��"%���l��(%�ȓr���2%�:-y�E������T�ȓ5���,�&.R8�;tA�I���y�1�!�]2�^�ɤ�۸e�")�ȓb<��L��'� H���7����ȓTt�;W���T5��J�JѼQ�ȓ(!�t�Q��56��DeB&&�����\��HS�Q�#H5�7�����ȓ'G<��D�ީ��)
�{�n����&���%I+\�����(_H�)�ȓ$ ��X�(�M���X�lίFd,Ԇ��N�Б��GE��ȵV� �ц�8p4�i1��)�0�d�(5���ȓ,���lJ�S�^q� O��qXB��y��S-X�]J(���/фȓo����Z/NдaJS)�,SH������ ���s?IS�ʨ ���K���a�T]���"�'W���ȓ�ҙ�(�j]8С��K	t����D%���6 ���'ƈkol���H�<�H�+H�Z�m2JAqs|M�ȓc��	�пQ�r!!ٻ��-��k�}K�g��kkX�ȷ/̞+h������p�EޢEBp !)4�r��S�? �q�D���&���9c �Z����"O��(��;'jBpY�HM=�6+�"O<Y��Λ�P�ɇFB:sk
��g"O�h��
2ͪ�� � V���v"O�  r�	*l���Æ�2Fq>,�s"O���B�E`�� ��n�e�.(�"O�X�i�'L#������q�+�"O����gO�
=��Ç,��=et=�""O����`ƏD�ሕ(P�+e �p"O ��$��=ik�tKb��	V���"O ��b�͜��Rv̩�tj��#!�$�;O�8v�G�b ���hժO!��^
ƴxQe(:��yB�\�|!����"C`ْ=��p�5fX)un!�$�/5qv-)5�ؚ?�\U���_3w!���\j��`��Q�`
c2;�!�d�hp| x&�[�v�ޕ�硎�z�!�d�&�����&#H�`A�� ��	�!��3gj�)4�z�.���/�:Pv!�$;6L$�ACA,y�}y��D�Tq!�d\�1��C�Ǚz�����/�Qd!�$�������	������\!�dD@ƕ�e��|�L	����2�!��ԍ�����-pk�♫�!��׿�p��,��*��>"!��Z�vh�(��dۨkh�� ��ʑ!�ĉ�WHbQy�Ř�{W��;��]�!���bC�q��]�t^�@�u��2W!��)(m�Vɧjւ��-ڿ`Pİ��9&�yypH2f�X%;��y*"e�ȓil���3�7X{�ds��+�\!��Y�`���	�0}[0���D�7�D�ȓ{�^���@8� $
gj���ȓI�������>��򰢁��Č�ȓ`�`���#�&���b�6�=��o�(���iǶ	�|�q�:zi��{����W�c,�e��!��<�>�ȓC.F��K�:I�W��|�,�ȓct�lSބxe4����A�^J��$b��R.U�f��WOϔ;s݄ȓ 3�s��2:3T�{��4U�jt��|���,&(AR6P�:E��4��+��F�|c��G��9l����6��<҂&L	)��D���]b"���'Z�8Ӆ�ʲAM,P#�/*~��C����pꀩc� ��!��=jrzȆȓL �%���ϥ13��Rj��SP� ��;�6��m�;e�ց�(�D��p}j�Z5�T�N��HZ��0X�a��~���@m��n%(◡�;u�@��ȓ|HX�EaV��F%O�w�\܅ȓl6V�C��5M��1㤊\.}�r��J�Y*��;���v ަG�ެ��9ܵ@֪L��&�Z"
	�l5z��ȓ:1�� �"�_��� ��&s�Xy�ȓ.�x"�K�&��rRզs,v5�ȓuf�C�G;
�����i�F��i�ȓG6d�	�A�{	xE#G�¼Y�����B$e0C�)L@��a3/@9D万ȓ;<�,��IR�e:^Y���Y1T�لȓ�����ǘ�7F��' �?����ȓM�v�rŪ��bEwv��u��p�<�����2�B8l����h�<��N�(��#҆�	=�0��,^�<� 6A3r�]�{�Jh8�K���l��"O��J��^: 58��&ۦ���"O$z��*�r�y �%]�z� �"O��eʸ�f�`��ڻ��y�C"O�is�PV��w�ă����G"OTA����-y��i�傗��� "O�!#EM�a8�2��Ir*��W"O����ЕܖdSF�_�Iph13a"Od����Ǧ>2�!�R₻Cf��"Oh�aK�JaV�Yq��1+F��� "O*|�'�Z��6�:ro��!���"O�Ͳ��S&u�H9c�,V�R=�"O� �Ce�!b���P��v�"��"O�,#LM�=Ϫ�J��ޛL��15"O�0�%�_k�L�C��k���"O�(�POF2|�� ��b�6`{0�W"O�8kP��m����f�ʉ ˺5��"Oj #!�B�t&$�h=����!"O���p#��y"p�� gQ�o�8<;7"O*m�*�=G7�� G��Y�\�"O$��Ea��	�d�hסF�'̴��"O)�\����
� T1�"OXRUmąD�}K��_%Wl�"OP�rV"ڏQ��U��(W��*�"OX�;Ge5;�*x9$��t8��c"O|@ N�;4�K��+C:�t'"OV}&��"��I8�*>ͨ8��"O��T��3ޒ�c���J58"Oj��R2�;P�&}��ݰ�"O��ʊ��)b�a !7'~}��"OX0yp���g�I�����)~��ʶ"O*$k��1gI�ؙ 4Qb�-�"O$@�DI^�w��c��PH\��"O�a�C�����S��J�c;,)�""O��#v��s��x����)���"O���f̄n��a�*��� R"O�e�+��Xs'�� �0T�e"O��8
���2��Px�bu��"O1F��# �����N��x��"Ot�D"�^�r��J(����R"OL��R$=O� 
	�t�^YR�"Ot �����Y���:#���	0"O�ٲ��Y�9¸���;��!�2*O��3#�0q�H%*0�P�&옑
�'晲�+߀r��t�0H,�|93
�'@����*]dd��B,�=Y~��'ओ���+Y����
9�;	�' t	$m�k��U��&�}�	�'�&���0-l�0��ݭ%s�|��'��5�v)��(�ތ����%^�,3�'7~@*q��*O�l�` �>T�❠
�'Ҋ���Z;�0<xC��~��ȓJ�<�r���7��eC��W�LT�=��\xH�E*˕/Kxţ��y�V\�ȓ^�� s��>��L�&#
m�D5��K��(Sr�ПibPȨ�)bʌ����Y↮��J����,9��ȓOs��h�eS.9^]�V�	JO����Y>>ҰD��[B�\ f�?"%��\�I%�^�z����C���$�ȓU:�i�IƾD�6d��%�72Up��ȓn�6�G�ދB�(!���Ԭf�re�ȓhǒIyf勏V��	�$�*M�-�ȓQ�J�0	S/(�$"޼r����S�? dUQ�F2D'�!3�%g׊��"O���R�	�����f"T�I�R"O*���H��	��X�"O(,�:��s"O@%�A��I4�3d��|����"O���PTƔ��7*��ܘ1�"O,I� ��Z�R&)�!p(�"O��,?ބQTN�r����"O���6� ._H���@�c�B�"O$�#W��f�.�	�-P/e�-�y�(@y

����b��Q��)�y�ڒ4�.T�s/UBr]Y���y�'æL�``r�J�J{��̦֬�yt�hY #�FuZ��`��yҮM���[�b��B�rՀ�`���yҮ{md���ۄ1���ϑ��y�/�S5�p�"��R0La�jR<�y"*�^�b�[�E�Uk���A��y��U(XLV��0�Z�d��L�8�y�jG�y��в���?%�X:G���yrjڼ[C^��7L#�1�ǥ�y�D�;�Ӂ�ٝdd��*۬�y��\�p_�țG��>-R-��,��y�kŇ[�@�n��l��AB��y��2E)Z���e��,ؗiT��y�fƊ1d�]���(�dmӠ�H�y"(�OJt3�aP����-��yi+L���b��K�y�
Ì�y�aE0/mnQ��͚H{|A���Z��y2�,P���F��6x5����,�yr�R�%���@��>[�@!*٤�yM��vI|i(,ߓ/�R6H8�y"ᖩ炵QAC�0#�,���eR?�y�΃�����Uj��"��!��&N��y�ZK� x�#mL��z�����y��#j��G�ց��aQ&_�y���*�Pj�jM�O����	/�yR��rbz�R2�	)Hxt����)�y2͓0JW�1�R�IH�%��
Ϳ�yRXn,&�ХNR:D�8���M:�y�bޞeOZ��qb����Ȋ��yª�#kTⳌ�mI���e ��y.�8�`C���?S��屐F1�y�E-6�����vq�m(�	T��y2��G?��s��V)m6&AЦ	��y�CݍJ�,1��f[�A�m��yBbD/�w��]�~�:��&�y��ѮHK��Yo)U�(T0�l 1�y�N>_Dr�AE>`8�������y"�ѹS�,b�ŇDӆQ�Q�ۂ�yr�X$r��XB���pLf�YB.�y����
�9�N�_����͛�y2kD�6%ƴ�4#H:	8���։Z��y�"7m���,������y�K�t��=����O�> [6���<	@�X\dA�*�,�rv+�L�<��(��3�a����3��I2���<�ƭ^"���� C C>���"�g�<�vif�����|H����d�<%��an~`�6����~u�5$1D�l��(�+w���;��6�|!
�/D�8#T��8K�\i1����xRa�/D��˖IZ+{+N�)w�i�x<�A�-D�H �K���*��l���j���$�!򤘮bް*����3��q�����!�� 8��]$R��)�'U��:'"O�i�,Jd(�&��'�.�I�"O��$�#[le�5&�!��	��"O����1i(�pFĮ7��*A"O����~�*�Q S�&gl����]�<�aǺ)��A�K�U���k��AY�<��f	�:n�5U�a�[���N�<�C�=B�xc�a�HpVU�Q�KI�<��kA�5�Y�Y;*�	��H�<9��9�ȉ2��.#�ܽ��!�<�4�g��YZG�*{���C⨎z�<A�X�~�e����N挓��v�<�f�C*i$ ]����!bY����o�<9R PbVV���c�G>��C�l�<��m>�h����!F�S'BW���	\�Ik��~�,�%v��`��.d��#��y�S�\� "u��0�*�j�κ�y�H1~�91R�J1'V��х���y"/�;>��z#��	�L���fI��yrB�5o~�[0i!9�,���y�׫K��U�o�,���A�ʊ�yb"�Tʦma&"�1~�Q��W���4��#�g?���8/@��@b�8(n����E�<���@�XbKA�a���F�<ɑNM�Izn�BE�˖:r(Prs[Y�<A��;��e:7$��j�(q���Q�<	�gE8!���a� ��Ba������f���ϓe�Ȑ"�A̞m��%�U�A	T���ȓ<�P%�h�(�,�b��&]�����,'��E��'��)��l�o��9��`ەq ���'�HU�2&В�`���=����'eH���
k��L!��.��+�'������2F�lt���=U�~���'�jȁ�]�!��$`aDZU�hQ���O�u��ɴb|hMj!�����"O��*Ǚ	��4J4�ٟg�Ƚ��"O<E 3kR:u�h�6NR1X��t+"O��"C�W-u:��Q5�B�h� "OZ�-��:V>`�Ȅ�j�̕�&"O�`Qqi\)>b<�,.B�ر�"O�1���16x�=�K
(&���	k�O�D�A�L�����EDB�{X�IC�'���r��Դ1C��	e��*m���Aϓ�O��Ĭ�4.�n0�dbQ���Q�`"O�	�o����r��0&�����"O���U��bW���.�8m��"O����F��.���M�:�z�"t"O�лq!ZiY��ƁX�ht
3"O�-����?P����	A!tv���"O�x�#���%s�! �i��Uw8%£"O�Ċv��Z���z4(�A�D�B"O����X�����!D$q^@�u"Od�rc��%=�z�*���!X>e��"Ob�r��Y&0j�	�g �
C��cu"OVD2��%��$ɥπ�&�>��"O�)R��*Eƌ3�.�L�|(D"Oh�*�Ϳ+ɘ��3��K:�q��"O��1�O[��1�� 
0\�G"O��*J��U�(yp��'j�(�K�"Oz�s�ȟ{�tk���?|�vM��"O�,�2��7%έ���P�Z=!�d�>4��Y�k��pYTj˦r!�V�PV�JWNCW�m�g�JDY!�H/D��B�f�]�D��W��8Y!�� &�CņY
�x�ð��`,��"ORxף���8,�5��,r<�"Of|2��+���w	��W%4e!�"O���!�0�Qc��2��U"O�5��#�%=�9��H��@�"�y�"O���@$��
���B�:qx$Y�|��'^�Qe��*b}�	ͤ)�b1���O��`3��T��L�@DG�$j�ABg"O�l��S�A��{��4�^�J�"O��4��sn4q����v�f�C�"O�գf+B�e��!�æʟa��L*�"O�x�0�+{U�P:e^%)v�U"Oh����@.��@��&ߡXd~�h�"O�����'�li�g��W��"O��"��)Y�^�c�%_��q�t"Ot��W��+Hp��'$B��tu�4"O �I�;kq���P�8�21"O ��"-i�����M�.���"O�V��`�l�r�A]�m�RAC�x�<�EM�Q����s��=A���劜|�<	��n^i����6�N𰥭z�<����B������=)	LѨ� �v�<��DpaĵJ7���y�p`�Ϙt�<�o�9QR|A��Ԥ�I� �r�<����v%��q!a��T�FI��
x�<���ّb�K*#>�d��
�C�ɲ1��K��Q=m�( B�X2V�p��0?I��+�j,r���:hΨ�z�MJl�<U�T3`��e�h��]x�2qg�q�<Y0 7=�X]�����=���G�<1c!P�Kp�-�j	�c���!��JB�<9F
�_���Ӳ͐���a�8T��""�ڦNm��j�N��$R�ਇ;D�pèI2GM����M�(	���y�E8D�������W0Y9�d^B�1��:D�dB"���Q�����'�(x��L.D��Kd�>���v�۷pH����9D��0���b9�	��ڳK6�8zT,9D�0i��$X�6,�0k̴&BllCP�2D�cF�)a�ِȋ�~���@��6D����NsMҨ�	6�0�i5D��y1�H9E�Q�%�qe,�릮 D��21Kڈo�Y*�dEWN(�q�>D��C�E	S�X�℘�c�.|@�l9D� ��Aq�$��A��0X�{�6D�4�bIX6.@&'C1>��e�'J?D��� L�\����ꋩGx�e�0�<D�0��+ֲSܤ1�$c�S�n}��&<D��$�Â�(\�$�*���#�O2�pG��'�Hlٳ��v��-��✗^�B�I�00q��j��']Ĺ䨜�p�C�	�u�h(�ʮ5���H
G�C��-K>e��K�6�,I�Ò�3 �B�	v��p�B�O�I]:L�%��
��B�	0�ԲEgҩ_A4*�,��#��B�ɰk=R�v��,J���&� 옢=Y�⚟DЀ�˶9��(�g����1�i'D��p�c@��z�� �&S�-(D�x �e�S4�S�߻p�|�'D����ѭ�D!t��9J���2D��b^�3�|���kH�^>�C�A;D��pG�$9j���B/KB��.:D������}�Y[U�S�R�{�n�OH���O ��<�|Γ�y�H%�"!��-F�Ҭ�cmְ�y
� 2�G~,
�	J�JQ�p*O\�8��N�[� 18�Ǌ�B���'�uxa�Q��� �Ü	�|��'���1�ƣ��0P؈(�q(�'��i�@@�'� E��g���'N������-UAJ�8NR[�������?1���S�4�'��	4?Ί�0�̨O��ha���:'jC䉽3�5¢��2"+�PW/���2C�I-�X,zA`��R��Qް3C�	'�X̑���D�:揉JC䉮pc\d2�o�!�f  ���"2�ZB�	���uAj��>̡���1gC� *)��6��%���[3 A,94C�9����4ӌ!÷�g�B��.$/�ű�'+�>(�`�ނv��B�ɩe�F�*A��&�D��ڿr�B䉹2����PoȭN�����Ӈ[DC�	8U�&�Ł_�\��a�g#&��C�ɢR��|��ף5;f��JF�,��B䉍;��P@���*��x��.
C�pB�	�	$��K1/U5,g$o͌x�8B䉸C
���D@U�S��PoK3XZC��"���0��T��d�&cT	�B�ɗW�|ii�Ыn������
&�B�ɼk�=`V��'��$$�/��B�	1[,��Qϐ�is�U����m�vB�I19� �Wk�H.4xԣ�h�VB�	 /�� Q�q,��tm�%6B�	�%�^��	N�W��9C��K�by�B�	�d�x�C��
5���"��y
�B�I�wd@���J
� ļy�	�8�~B�I�,�H��z��D��ś	~JB��&F&̉��Np��RN�"�C�2�$4�����dlѡJ�"r�C� :{>݁��Z���,9%���hC�ɢZ���*�e�>P(Ё�!R�DC�ɗ��(���ҋS�`��E��0��B�I�o߸(���Y�o�.t�`��K�zC�	�)�h��&`��<Q��&ZPC䉶���"eJ�C�
���!)�HC�In�|���49�Jty�I޶���D#��
��.m�����͆@�U�U&1D�0!h�\�e��h��s���4d"D�$pS��:z�v M�w*�UcE�?D�\���XU��a
�ke� Ye�=D�@��oM�H�\�Bҡ��L䚹`�b'D�PKW M�>�����&Jhy���04����-�X�x��IT�'y�9�b#�۟�'�a|�1u�=C#�9(���� ��y"!��n�H!�I'@l�c��y�M��q#l��v��?)�ˠ���y��z�< Pi�	-N���7�,�y�E�}��D3� �\��d��y�%�J� �Z=d4����e֞��x�-Ř˶��E
�,�jS*�J���~���s#̻� e9��N/h��3D���c�3����K-��Z�F,D�l
UB� h�p3���	s�&�)s�+D��YW��sE�l�5�?vM�<�+D�Ԑ�C�,�:��^�<��<�4�(D�����
���iզZ�r��ԱrF1D���w�'od�b.ڿ"q�"�e"�D<�S�''����1c�o�0e� иG�*���>I�=��S�"�~s��1!���S�? @�1$��gY؜ScᅯL�����"Ov� �	�fM�b!�3���b"O25�q��6H]H��@J1(��铲"O��s2	�o���@`��R�"O������8�X,1��B�w��I�|r�'Gaz�Kñސ����аl9�8�fk��y"��JI@e����`����� ?�y�Z�b��X����#n�ı"% ю�y���?w�Ұ�\m'����+A��yBF�+eT��pAGl�C�b�;�y2������1�J`�a�EjA��yR��#5Ұ��WE���Z��G2��'���'�J��B%��^ ����q길�'^�$���_4V�疌m��'�PـqeF�є�����_��hK�'�v}{f��f��2��G	=��'�p�amŏz���۷"��\��'�\�qW?ʼ;R���B��'~�����7y���$�|X��'x�� �Ʋ_zt����Q>��8�'��XZDhΓ �܈SI�d�m
�'S��s*�3y \k󠁝.���	�'�♀'�	5$�N@PݤY<Ĕ
�':����O��_��C��F�z<��'����B����(� �=K
��'	����.E�7M���a�8.l	�'/N���C�L�@	^�y�L��'^H`%*H�wvYWK�<���Z�'�ȝ��OX�>m�«�	#��H�'�-�q&�vo���bS�f��p�'�@�%��^~1�͟�Vž\��'�PZ��G�t���@j�)�	�'�vʢf[��u��;����'o.1q��*l~:8�!O���
�'s*����9}��鑒�Q�C���'W7kӛ^krab�0uԓ�"O��#�;iHܘ��Z�bf�0�"O\][�%A�S>VH�0'��G޸�"O�M4��0�xb7J7ODJ�X�"O`�ԬF�|=PN�(HI���"O�dZn�b]�X��툋r�4E"O��0@�ٴP�����+h�^�j�"O�@�ȗFa����٨.�P�"O��y�F��R�ʀء�K�$�NP��"O����G
�l���`����v"O�����a͢�R`�oA@0`�"Oh<!!\�n[jm���CF�a�S"O�4�� �34�{AĄ25(�"O֭k��X��"h�aG=�=�!"O�rD���ڐ��R�1�"O��/,�G��u3 � "��)LO�L�^"3\	B�kЅR�i)�Z��D{��)����X���G�?��|��D�!�CS>@� 	4���a����p�!�DY�)�l��S���J�T��%ۑ�!�D�/Mo�=0g�ހ/bj� ���0B�!�5`  ��`�W�bW��y� ?"�!�ğ5Zx�|�� ӟ>#(�`���X��	\��(��!aAաRy��Iq!�v9��'^��D{��I��	
�U�S�Ř�2�#�垃2�!򄑫r���9B��-�tȋ��\#I�!��cK��wBH9}�>�p�Č,g&!��_�[�v�z�B��1q�=!�d��KG��+�1_DT�B��I�!�� ��� ��(�d�5�ͻ^#�]�"OvP����g�T����ˆ"O"��F&"
D�졗�ΔC��8���$LO qq��[�g������)g�xm��"O�]y��B'O<�TX�n�;�`q�"O&8҆�k�J��֏I`D4��"O� sӨZ�,h'HK�涀�e"OfPk"���>�dH�������e���|��)�Ӟ&(lr�ʏ.|Ϩ *��C��M �@y B�*��T��/lF�ʓ��$,LO�U9!gό1IPܹ$_AN�*O Sa��t&�:A�i(t4�
�'��y`��ۿ@�}h@G��SN~�;	�',2����2%�>���?by��(	�'�vX�ܳU�jt�j�T�x ���hO?�%�c�����Eܵ(\��	@H�<a6�ZU��tʖ0` Z J�<�eȾE�0�;6�$&2�9!&^P�<	V���߶X[�,��=V�9�K_g�<���/�b0+��2s��֨�g�<yI��KJI[��.4kbi8�C�[�<��M̫C6�(��?�i�D�˟��I`�S�O�z�X4Aޯ���2�h�uhZ!�r"O@�CԆ!Mt�I'%�;h�U`�"OR�s�ݯEt9pGdMsHб 2"OF�����s�	�jB(�"OR�t&mB��+U�lqs�"O^�Sh˩O��}���ٸ@d���"O�U��`�<Z����6l^L�9�"O�p��>h��,Ly����P��y�G,i� �$�O]�x�$Lޝ�yH�74��Bק��~�^}S����yR�D�(�T�[�IQ� �y���c$�����C�Za3⌛�y�O�(����L�9�
UӢ�'�y"�Q���8�'Ӗ-�WO��䓱0>Y��B�B�	��~��I���r�<Ae��Q����b��Qhb �ԏ�k�<��b�5D������0B�B��Wd�<�p��0 +d��Q55�,xb5G�`�<�)ǚ8͊L�b��4L.`
�A�g�<��
�T[!��$BQ�	�b�<�!E�+�fP"��_7䘕���HX�<qFd�kc^�R*ӳ�ؘy�f�T�<��T�x ��X��܈wR��k��O�<ɠ�V�T6�\��Μ	0�c�ZL�<ie�X�����`a�@�t��E�<����[�v0Eq!
 0����'wj]��d?]#J! ����zhR�h
�')(��$k]7v�b�XaA!n��Բ	�'�l���m B��5e��h_\��'2F�v�V�8^j5������q�
�'�j�*W)�/9��r�eҼG, ؉b�'B�ӏca<J1DƬ�頨���4B��9�,Ě5�H�v����'_�zO
B�8hs���R'��̤1�gA�[��C�	�.�`IӗL�+�����4�tC�ɱ^W�I�)+���鱃_�y�@#>�!U矔G��,�J�8!X�j
� c�G�E��y	�dN>�����sr��<��<ي��=}	���`�!3N�1-�+F!�;,���05��&�hx�Y�h(!򤕥nd@I�A��v�	��^$!��J�0�h�  ��ҦVoTp��S�? ԙ�	*n"�L+®+y8����"Ox��b�ل+�����Ƃ"�`�q"OV$ᶆ>Sw"8B�@ֻ �x�!"O�Aze�ݲ���ZP;q�8���"O� ��Z`��D�����n!@��%"O���d"]#���#'#��"O|Q�K<)�ҍ�aB�#|M��U*O���R�V'@���j����%�|�	�'��أc�Ѡn�����΍
L4���'0��&�[���5�ӶWΆ��
�'ٮ��n�%y��h[�*t�h̈́X�<q�dĩ8(�i���	(�u �F�V�<ɕ����a� �4v�փMP�<i%�\�/�����J��оqpTo�Ix�x���<Y �2$��P��CC�8Pp�BO�<�2	ؾfN\В��;���cE��r�<��&_r���I����(��vOl�<i�&A�}��({�@��yq��&�|�<�T��>:��t1q��v6�8�a�}�<qiA�_��ͪ"7����� |�<ɠ��t��႙n����F��@x���	�<IA�:G��x�a��p 2�Gy��'�$p����*ܐ� K�=T�<C�'GjHR%��FA�I;Ɣ?��D;�':}��E�%Ɔ5�P���'s
�YD凅^({�EQ W��Z�'�IbW�#�My �\�t_���'�r���M�zh8�0D�*.@��'���yG��<D�Eb�$j��
*OX�D�O<��䆥p,t@ .Q�9����f^2@!�dՆYz$����O��1��V2-�!�d�(<�vyZ2�Ðr1R�cׁZc�!�$E6~A��A4��:�<�1#��Z�!�^A��&�Z:C�<��#Bk�!򤁍Bc"�,
�&k�ıq,��G!�ޙ*ϰ ��l�.V
^H�e	O5�'_ў$�<�@�
f�,[�z���"��F��hO�'f׊D��cP
AZPIa3A�o5����i�:�Z��ͿP7v�pӄH�	��ͅ�(�޴I񣍳F44U�vb��<���Yl�y�ԏ��X��vD�4tN-�ȓ�@��R�#T	޴\5�)#	�'� H���ٯ5c&�. E�����"�'���՟�%?Q8s嘇m	��
��Бn�\�!�vyb�'�`�hP�?J/h�B$�Mݚ���'fL%I��_m6i�D�%pt�Q�'������H�3 ނa�4I�'|��K�ě�&�x Ӓ+�>?>ac�'�� �d�=��B�n��N��'���բI�_��% &��(��	�ϓ�O���Cߡop�t��I�L\Q��'��'İuK$��&"�l�ň��$�	�'����&��� �>���h�'w�I�й���y����r���'�pH�$�H2J�+�ō9(yZ�'^����oٔ+�*M�!a��D1S�'0 ���#ڏ͠-P&G�+($e���<َ��n_�`�~�;�a؁o�jAq�`[��y����r��A��(aSX��L�;�y�G�%L\V� m	�D�jP��.�y���+�֘�/��7
�8x7I�yB�V�_g ,qs�N[M�Q�� �7�y�k@�KvRݱp*	^f�0G���y���:#%%M�B�������OX"~� ���`��
�bQs!�T��(�"O����Hǖ�.,Z�*d��=�$�O�����BE��r4"�@{���!d	i�!�d��5F�ٲ$ΏLb܍꠩
X�!��/b���!Xt���I��!�$�"�����c�//>���u!�� �!�[�V�����H�g'ڡ �`�6�!�Dяw]���P��(y\U����4~!�$O�qu�I��Η�7_� a���Os�O��%����W@J�E�����:4�|�r"O8Tx��Ma�����ֹYKNl)�"O8��F�1f�V\p�Q��,�W"Ov��q��*5N�S�u����"O��B$B��-�*�x����X��$"O�0�v+�'P&���!e�Tػ�"Oj	Ja��+Kl� "#��/s���"O>�P�Q�|�`�@�K	WBH� "OP-Iv�2���+$"W%M*�01"O�Mk�A�"�V�XuE�0���P"O��1��O�{���oԉifZ��S"O��i�Z bla�9-d̼��"O|�ga�"("d�І�T\4��"O$�� bA�TU�����:R��6�	h>Qr� Sw��]G�${�<�� K*D��Y�l̹ ��%��bz>d�c*D���s�.�IE��%�J�膏&D��
`�L"���u.��xf��t�$D���F��0{|�������� �>D���2��tT8�bJ�`��=1Wh;D�i��$GR�pD��p�E�c�;D���GvK��3o��#Y�0j�C;D���g��
R�Y�N
-8-���N5D���1K��/�!sP��?3�8҃`.D���Q�&�ykDFKl�z�+D��� b�I�F��C:l��=D�|�VN�5�bi�CE�<]h49�e)D��0�Fw��T3����7�'D� �$FF�4?�A��!P6�{!D���j�;��JF�V	Jz���%=D�L#Ώ*�� ��J���DN;D��ʔ��#|r�/�fl��J;D�{���v��l]�o�F ҂�$D��8 .�<��<���E<N�"h� D�8
��V�<��y S*��*ʼ���#D����h�q=�L���\%_� CW�#D�hɖג(�
��:�JL �� D���0���e9��֫WZwH��O2D��07F��LU���P�!|)�/D�4���8Tn5���D����9D����@G�8�X��֌��x]���@�7D���0慺Bbd�![�cޮ�4�?D��R�E6_/���$�'S���SL<D���"FF0D�2J���)E!��5�-D���Â��yTm*���(w��(e6D��['ȃ
b@�u�%Q�g� kơ.D�H���<U0*QS�G Z��Y��8D�<ˠ�6L\$T[ff��y�$ȗ#,D���(u���Y�F�hw�H G~��ȓ,��I��A\y� ͫ�ϰ%�E��)?dxEj�9"��[0���9��e��>-�}3��ބP6d�Qe�s�U��
�P��H_"7�*���S�<�t��ȓ?ր���	p�D���[{
�P��5���Ѳe	�}���s`bƐrG�a��S�? d�
	O�>�<�����8���s"O*����Àc�qR���733ڜ�&"O��+Q)Q�4����T΁]����"OP%��)X�7lΩ��P�/{��[W"O�9�AR9>�����E	�$ ��"O���6��o�4u��DC�?�IZQ"Ox�&�Z u�X[w��
,�r�c6"O �{�+M�MႽ9p��&e͞��"O�s��49~���l�2dO����"O�}[U(A��Ru�ΰ9=C"O乃0�PM��#�i��>�J��E"Oj=�(U�>kҨ`G���8{v�s�"Oބ��kF,~�UA�=b��"O��R�ņ"=�nx3�+б_R�Q""O^K��	u���t�ڕJI�x+�"O�9�!�K_�x��ʺ���d"O6 8eo�7IQZ�2bJ��im��U"O��&A^�xETzw(2_x\)!U"OL��f�� 5t�� Ƅmm�a�D"OHHpC�1K�AHEFE�oj>���"O|����jɦLzD$	*'<��"O�h$+�'�"ɦ�5��MQ�*ODDb��U�ZݘxaQ4zD��)�'k�,@����.��a��$�+�'�h8s� �\�#�ǧ-���'�� YU	��]Bp<(F#C�XO���sad�i�՜G�44I���<�)��_]�U���̪���80��<���b�H�	�-(HHt��/|퀩��5��H*5ןlNB�"��n����\֩�$�3[�"�`�ɖ�B7�l�ȓ\2J(���ÞB
���,��!�px�ȓ/�t4��3HWX� �0>xb���.�"��.O[��B֡��R%v��G�0��U���Ke�Ŋ�ޥ V���ȓcDԲ���
� �X��P�<�n܇� � �"wkN6k��hԄY�i#Na�ȓ[�p���ȱ{ZL�8���a׼�ȓ^ۤ�R#��1���H҈��
���ȓ-�c���2��K R�m��y��z���	dɋ6�2U{B�BE����L��4)�Ƶ�"��4e�H��ȓ}����חe�:����/O甽��^�D�0�ŝo9�b��(��ȓ9y�f��#�\�Qf��L�jI��L��UrƯ�#�hH) ��k6���ȓ���q��=Y���UDIRC����	�N�B! �{��	F'ZЉ���f�����?h�B�إ&
��ȓs��§�ۈMy��9`��Ś8�ȓb�~(eȇ^z�����k�e�ȓ&�������Wgt����^�|�.��ȓo���(U-]�w�|�ǣ��;��܇ȓ�4,�f(�"t�2��,�+Rq��ȓrF���j�f� )�C 8���lov(����)��ݨ�M�����U���kseA�?�<� ����ԇ�#��5�oZ;Ȩ����6�`݄�((.�:ȁ1وe���2R	��z�,Z�'�$Z7���a@�:yPa��=x�1"���5VH�7�o
9���8�{4�oi��ȠE@����ȓ]���f��lLl� n��P��4k o��/�A�3�C	 ����S�? h��Z�'PF요�@qh�H�"O.�z ��7Bm�@q΂[��� B"OZ!�CC�4!�t�*2��L,�X�"O�h¯�< �+B��';��"O.4�'˕H��e\}3R��A"O��KTo�������
G��9"O�u�MB�M1~\؃���
8̸Q"O�d�vg
�zܞ!
�*�{�-�3"O^D �h?*@(��(9��V�d�<9S	ϦRH(��͌1���s6b�`�<I2��i����E���K�� f�<Qq)ŗvy����لy�K�%_z�<�s�W�W�Ҽ����h0^8��z�<	� �>�p��lq@nl�ll�<�f_��`Pm�
����HLk�<A���EFI���8E���*�i�<���Ɍ�p����2~ݎ�U i�<���lR�9pǉ�-J�n�;6(�a�<	0b��"Ir�Kpi��J���ER�<�h#�b���m�>^Kby�d�L�<��@D8)h��o�E�.���U@�<��gǛ�<��V�B����1��}�<���[�H���ڳ�x
�y�<��f�
�1�f�Q37�j����Kr�<����T�pPh&�:Zɤ�	B �o�<	G�U /38ٸ��I�P9�1i�<攈w��+e.H�8<���Wo�<	BҡXQf�����>K�\⒊�l�<Q5F#KW�0[�d�?��I�
Lg�<���Q��Ԣ7#*]+(�qeY`�<Q�nH�+L�(�ѧ�(s�4aqP��s�<��`N�G�d �$#� }�%1�iIK�<�m�	N~9�1`�5*�f�Ѳ�#D��is���<�PA���q���"D�쓐�� ����~�0����!D�laGY(#b��+��H� ���>D���Q&�6��(�m�,F��P�f*=D���%&�"=�Y2[��ZdH�;D�d�	� ?�~-���˹b�$�)T�7D�̻�/Jjk$����t�  i�3D�l ��ڸn{̳��{�hrկ#D�r���1#��z�8J�|{�n#D�@� �I�C�L����'pW��D�"D�<x�J��.CCA"��3�C�<�rœ3$0��Q7��M��|�<I���*��\��'�u�-֩D�<�u� 8����:\��j��@j�<s柣b��\8S:�`
�}�<��^i��!/��]����z�<��+�%D�NLc�I�vtC'��t�<�j����1d`Q[�j�^n�<YU/�(|�Z@� E3���"�g�<� ��@�H$Qwc#yє䑃�n�<�7d^� �,)@�͘�BuD�AGg�i�<��L��5Qĩ�E/�-�u��g�|�<!#f	�V{���
c~ٺ�� a�<)"��)j&�;��8C�A3��K`�<�a��&_����mT�)�9�� v�<�bm�>
�t��@�.�������Z�<��,��G����37��J�%�@�<��EV�Ш��V�N:���b�|�<�eK.a0��5N���<b�^z�<i&��l(8Xcǈ�7&8�ө�^�<�WQ��B%Q捞98G @�Q*�@�<� �=�"a�2xP]� %\�D Z�"O6��ꁪpt̰ɠ��>q����"O��q��!\�P��"b~� �V"O>mI��;%^�0�ƀ��T`�G"O��K�@*7�=c&��;����"O�|z%욄R�t��R���+�`1�e"O�Ei�L׶q��y�̘�=r\ 3�"O�i�w�UJ�l��� %W��I�"OЉ�6��1�ġ颎�I Ր�"OέHDJ�?L����,��=FFxhG"O���S�,M�Ke��0��*S"O$؄�J5T
mI�����T"Oʑ���G��h�z��`Ј�;7"OV)��bT5d�����_ɔY��"O���k�
5������S�4��"O�!	� ͳ�0 b�rpp5"O`m��WzEVb�iN��e�c"O��JA ��'�$0sHj�v�@"O8�B�Ǆlk0�P�&�'n\Έ3�"OZl#�ݿ}� D� �r)R)��"O8h�&�4��R���v+<-;�k��yb��.Mnb�0F�iF(\�ǯ/�yR�ܭP�6�*d�ɫa�ZUsw��+�y"��!��];���=`����Ϸ�y"�Ă\��zd(�\[(��G]��y���"6N%(�����@�G��yrNXUo��X�^0u�9*"�/�ybLǀ(]��R�K� �ܩ���;�y�̞�d�"-Z��5q<�@��
�y�낢X���s�nBy�Ι��E��y�V�������eV�i�H� �y2E�.k��-�&�K�[���bw���yB�]8"����Z�WLf�^���'�v9��b��ײ<a��P4,h�-!�'S"`�s��GA^ܰ'J"$�$���'ff��a�"�Ќ��GK8{ܔ��'�"��C�&�)A��f)9�'w�!�f �x+-��m�zx\$q
�'f�iQ��}��p�� H�n�BhK
�'�`�y #L$#ފ鈅��<��M1	�'��"�n�2T�$�Y�8�z+�'�x��� �8�"��7?���'��Ј�Ҩ|oT�q�/�'�2��	�'���s
�+K ^�S���<u��'���F��-c��Q�ȥˬ%��'�0���hW�%	��Y/߄W
I�'v����
]F!ba��!�x�'��`��-�?i�Ib�5��h�	�'
d�ӄHa�z��uN���0�@�'U����&B�~�Ia�*ɾ�dA��'�2�ڣ�؞6��Sd
�=,0�pۓø'��1��/h�>	�)P��p���'/t���)�Ow���L�3zP.�y�'.0*%�@�~������l������?��{�A��}E#g�^�a�f����$�y�X eR�RTe�1c�&�1�і�yRA�6
�}�3�C�`�܀2�Ǝ%�xb�'�~`�� ��/����+S�~(��(�'%�m����.�%�moZ��
�'m8}a�#�?*�&�[5خ`QX};
�'�D���ŻM�@�!���$`0����'H���UZ�#�JK*b�>���'T���תc����
g�Zl��'?�� ��D�����z��QKUg��y
� `zW��6��p7�ٵ�H��"O$���/<�أ0#؏�^�Y�� u ?��fHW>'m�u
W���],|u[1A*ʓ��<A�fҶL��a*�֣��h�tǗR�<)"e44�[p��#3v}1��E�'��y�U�~���#V5FE�QxU�N��y�OŻI<�pb�AW�8y���yHY䴓�e�06�>(3b,ל�yB�ƭ5�P�B�F�'K�H�FA��y���cN�ZFi �/����$���y��O1�q��f�q$��H��'pўb>�*��ӹt��wh�' ->�p <D��	p�n4*ۿj� ��@$D�����d���Ҧ�Ŷ+��pKS5D�P3p$���=x�C	,sgf��M3D�HC1�%����eɑz&V�p�?D��������I�3f���vT3��<D��Y��Y bǨ|�Ʈ��J�!�a}��>yN�.K�^)��A��S��J���I�<Q��l������s7�D�<��
��<Ʌ��<3=�!�,�k؟`��9�e�c.JXГ��-HU�ȓW�p��B^�! p�[t�ҫ%OJ��%��I�/_�"��E[�@�*Uc���)OT��䔏z^��1�K��|��r�w?��lE��"
!�D�
@�<_����Ð���:�O��2`��>��+1
P$\���"O�Ɉ�ɢH�d3�
Ћ(G"Y�"O��8�/�9m0��˅�sGLu���]�OZ�A"�Qd�x����$'AΝ��'�^ +F�9 ��9�V�
�iT:���'Ж�Q *ى/�a��g9B�@	��(O���VH�4>�]�����i�xqɀ"O ȉ���>"I���#3�
T)p"O$��2�H�SV�-�T���5{��'����O�ʔ��fv�{��ӈT�����i���>YH���b̓3���'&�=�~P �CX�-�04�ȓ60���TO�,����ҡ2�)��P�����L�Q�Ia��/}t͇�	~�$�Μ��f�	E�� ���/��匃�O�����5с�NL{\$��� �!��0a(��{C)B)�Ȁ��X��!�/U�R��f�U$|�Bh��Ȳ�!�A(Z�=A4M��2�<�ÇƉ�Q\!��o� �����c����J�_@�v
O���`�ٛA��&F�����c"On� �ŮEk
�;U�Lqx���"O"����#0t�F��L`�����G{��O�d��eCP��3KpAy��	�)'!��K�x�Xh�ҙI���G����1Oф퉈?PF�ڴQ"+��{#'L
{�,C��ݟ�@ӝ1PHa���	u���A2D��37��2;��ixv��+[U����1���$X�i��r�V�S�p߲�Pw��x����A���[��N�^�[,MuQ�B�8X�����;'�#�-ϊt\�B�	�zR0c��&�EX�Z:G��HD{Zwuў�&w�,)0c-	e/���]���D�*��}񥂴�^��gLT.=�!�dC7~��@p�˼Q���6��4HD!��'1�x@+�M��b�lu���ASP�'��|���B�Q��� D6�Ͱ���y��@�@!t"�G�<�X�:S'X�y��H���R&��A[<%��,վ�ē��D0��� �q%hĄc�S�)I�|�� �"Ox!��F�6�v �R�H�6����"Oʉ�6'�>&y�Щш͐�򬃐�';�	q~H�l�R�4�՜^x�0��Kj��C��T�u���^��8<O\������]�Z��EoV��X���d:|O�P
#㈱):�E��l�>y��=�"O�U��q�̠�楘�5�\��U7Op�)���6ړZ#���b�4h�2���"zA�ɅƓ7����EC�2�ޥ��
ׅ?��MS3�)��<�/�4e�,�bf�̸#�N��@S�'݉'�>�@Q�X�QAT��w�x��F@�O<C�	�K��(@�
%e0����f�#�OĄ�<	��Nc�0S���T�prg�F#xh���H D���AE�X<�go��#G4��%�+D�<��E
	-��\(�������L�<��[�G�l�߾h	"���[�<�I̞?ΖU�f.޽'�IS�WW�<y6��Y�P	!7��y�n(�b��<	���=ړQr���ۦ�FASU�ĩa��[w�ł�K�;)s��"���F�<)cg�9E�fXr+�-.8H�[V/C�<�#�H�W����O��O-R}�fQe�<�4�V8|r�鹔�Į~���(@�]_�'O�yb���JN0�Qg�
=f`� �p`��x"�8���W��	wú!�5k�:8�B�I��>4cA�y�x��p
$_8C�9�����P�;� �@�*]7` C�{^�s�S�;�U�IHnw�B� � qx�MQ {�u�ń*��C䉟Tf��r%AҥĢ��Ů�a�TB��@$A�E.y�F9`�m�Q8~B䉮xL�ոB���G�����n��h��	�]_T����${M`�[��Q�ŪC��"#� }���jF��1��gX�C�>#>�K�K�-x�6p�T��w��'�ўb?�ZƤ�t	<5q'�U���ӡ�:D�ȈfA�j�"H����Z�`��KxӘB�	�r�ݸ$��3VCx�(�KB5�.B�	��H!$��x�٨�k� �C�1n6&��F µY�la{�n�?\�C�	6w4�"$NU-(�>����P�B�I �Hr���*!U��;�B�	!��i�`�61�YQ�Wh�6C䉆#VZDAcAZ�EWv9��?�@B��8#���	@�`bE�e�_���B䉙�d���$�VI��&B�B��B䉁"�����L#d�<�!G� �pC�	�%��*���Yn1�&�7h_LC�S�~4Д��I��(��+�h��B�I��1kb�Li4��;�
�wB�B�I/?��� a=8�V#�)Y�@�C�	6|��lS �||�R�t�(B�H�����ލ= ]�6��O��C�I5$��<��΋,4� z��VD�B��Hƪ�*s 3w����7T�VU�B�	�D��"���+7�H��Aѓ:�B�o&B h�"qk���u	҄�8C�	o����i�9X8)���?9��B�	��&9Js��Q{����	l-�B�I+��0���
���{EoH5��B�	�VB��H����BLQCg�+Fz�B��<|�����<DjJ�J6ÓC䉻}b�(Cs�U�0N֔bW#�O��B��4��xTC��R���Hˠ~��C�)� �A"a��"'�01�C�yI.�K�"O�U�9�,5���0��d"OP1��
�(�`�'� -���"O��3���5c����:E�5��"O�	 @H�dC�LBeaT�͑�"O%�c(���Y�V�H���rW"O�\@D��<����B
�)�%"O�%����/�2�A"%L�Jm","�"O����A��g)�e��3dc��I�"O����,�)YP)�b%�W��U��"Oܠ��#���&mK�W���"O�ݒQ�����!�A��f��A�F�=������p`�L�w1O�yyuܢ�B�����+��b"Or-h�b+B"�GCÏy��Pq�"Oƨ��d�.�p�עZ�zI�9#�"OV8@g���7�Z(S��S>KRA0"Onp�vkړ����V@I>H�e�r"OD`Ȟ��`)���I��� "O6�Xv���K���-�
?F��A�"O�9V��!c�z�'�03"�sv"O��#9D�� �B-T;��"O�e�AkXS~�����*�Le�"O�٫�)����{��B�3b���"O�����їQ�\��'�f��1"O&m)�E:�Ni�%'_?�(�0t"O�Pj�%LJ�:�&�d���#�"O����U� (�4
�g�Ɖ�b"OV����-�L���v�b9�C"OTM��L���v�$�C8O�N�s�"O\T���&JW���b%X�wL|�"O�H��&��m�IS�k9tM�Q"Od�G��V�8d��Iϡ6�0��'�0�@��8H�(�LЂ�'B�<���[�(�0T�cE��r��'�N2WOlc��F�:�d�I�'+>\��D��TpL=�1.P 6����'Z�BТ�;0��mAvJT,#"� 
�'���R3�TH��µT���X�'Q(ЀE/0�r�PňIK�N�#	�'E��SI��*���k�"TjZdk	�'��R�QSB�k� ǻ~��ϓQRF�{� '��]'p��`*'bC�d�z�K����A!��>v>p�Q`�-j<"���v+^�`t��;(*��i�W	F��2���C1>�wHʳ{�џ ��K�T
��T��$�9q��h+��:fI��x�C�*3�V��]� 9c��+��b>c�i�l��~�x5z���*U�R\�巟���d�P��ڷ,��>�"��x֖���2�J�#���2}��p����Y�<0c�'��x�7��>~9�����E��cԋ�-B"�������?Yď�D��
t��?��!�A����-A%����}R&�{cAƻq��ģ�J�a�ʢ=!�$_H��T��N��P9 �$��PB��ߩx��TA�ep��H��W������g�
 d�Q��O�XQ���?
��0�E�Pb0x����vR�VA���<�E��7�ʡ}U!���0^��@� �E���\c&5QAd�I�M��]�<�<��Q@SA l��4|4�Ղ�R
��g�p��9:���Sƒ̊1��\���l�5F�H��*Y_?�ABRK]��:]�;5�>����z���gD9L��B�K�k���%%�/x������"��H規I�^P��x��\�C-D5�G�FeD���(�|=��6�93s��8愮�xV8Ú\�Q��<�|4"s�@0�����ȷ�ܡ�ɣ37�Ax�$��!�ru�:\��s��޼�%�Y�BF8ZW&h����2"<�u�Q(73r�yqJ��� ��u�,Cz��c���q�0��X���
�'���A!*E�'$͘u�5$
Y���(Uݨd��I�,٦YJf��	�VSځB6ؘ&ʈ]���F	_���H�)f��ͻ	v�X)NO��@ p�� �x����0���$Ȅ ��)ba�[�3��=�p�`g�*� \jP͊Bv�гk�|L,�R@�Ӣ�I���<�p�x@��/�h����At����V�8���N_� q���1x�8�1u��*�������T<�')B�U�8H�6��3��-��Q�O"� P� $in�d##�388��1DÏ9h�v&̷1����щE<�H�'f�q��)V�$��L-o��:�'?X���sB�N�4^�8	�	ɘ[ޢ5�%O�'$�XA3r�����җ!r���G"*k7�ڰ] a!R'Ƚr:x(B��'����2�3� b�����eTIcq��93�x��
Z��}	��T6><�oi�\�r1/���F�p`�%�X�y΃ 5C�d9���8��0�O:�4@#4Oh �S���蔘K?��闀�nJ�����"A�tAEiߦղ��03"@#��� �M��������	B$���W������H�^LC��_�y�a��^E� ����&j�QE�� -z`%1� �!|�`�#͎4�Мa׈A/����'��Jt��jA�={�x���
�¸	�A/�ڈz��`�-����$�� ��ቄ8��=�Z/�����?��'ȏgܪl�#���DZD��*�b�2%�
�o2�ma�K�"@I�2)G�Q��D��>!#�`�Q��y�S�L�M0�⋲P
B���e	�r70y���O��ꌎ)EҴ��&��d�i�D@�9�i��nְojε�`�����Mѷj�r=�VF]����	2e]�au �?!�LX��o�:G��T��Cb����K��d�!���b`Ǽ&/
�� ��'l��ف�#_7aAl�3R��?���?qF��ڊ��o�	�P�����ݛ%����{�������!�@�7y�vQ� �|��6*X�p�
_�k��l��w�'��a+Wm��.\��}�v$[���A 4�4L��/D�b�<"��ߒA=�Z���_�T�y��P��)�I�4�0D��$�j�Ĥ��j�1_l���żf�����n�l�0Å�ny��1k���"l�r����3F�T�1W�򰛂+
>Gը�����=U@�K�;)���{t�ʼLY|������?�G|B�0Ay�K�,jah<��GY�?�!�Qժ�˚�l�yF�C�|�hTE�.z�����,��dc2����+/�������+Aժu�vlU;v�Ơ�bkΎM�z�?��![0V�ȍ[���<8����z�X$	�kҺ����Ln����-E�q�"�S�K��t$��_�x�R0)��;����p���5�c�bbIx�߼_� ��d���'A�)�C�d)��UAA�~��S&|[a��,�=���J���KP ]��M��� �Te���z ��!���[\:�+�6L��壯OB� qG�z�L�)��T��3��~ ��`���D���>�@� !�Ӂ~�d��Ɍ��@����u|'���I�H�S��	I�|�q��rUx�t��>b��t�W!Vax⼠����%YTR1��/ȘNd5�ٴY}6	���J�eZ�	Sa�8���EG�M���2��_�0��B��Z~�A8P��t��LP��0!P����'h��i�f	v\N ��@ė t��sA��=x=�Ѕ_%� HAҧI9�N�Sq � ^��a�+�%~��#1.U�v�`%�#�4hb�?7C�������n��"��=D	�c�h��Q y��8���1��>��i�`o���<�#@ @���@3���jϓE> 8�� 8�����	T�AT���LA��'����Y������ \�T���d�	�I�����L����žlN$�*p �\��5�D��"Y�ÑfDS)�9�4���t�6�����&M6�X�ĂI�.�07��	N�P�R�$�>�dI�@L�|�@�(%���@���y
�!�׀E6����xgh �$<"��Ɖx�,�i ��u��	`�Mád��Yq�I� ����.&�@�'���1�ݎx���Fx2��^Kޡb��07,���M(s���&�@�E�����A�K�p��k� �p��,m��qdL�+w�����A�
K���v�;@��Bg]�l��0��ّ>j��B�$�?\�AHO�S��1��J�'z*����R����p�O?
O�}H!��8�$��	u��� Dބ1L���-A�/Hn�򀧏�D�Y��'�(��$֫��'i9@���R&9G��I��R/{��K4nީj8Mʳ$�p� 咧)�F���F�;A��q�l.{����+�fq�t8Mi�H�(k�\�s���'"x�����by�T q��M�I\AXH��8u�8 ˠ���dE�	⤄�3N �4� �^DPL��N�+?y�  K �
$����*7����_�&-�m�3�Ϫ�آR�;���:r�<F�2�}aϐ?��K�+K�j����p�ѿe��	�ƤG�F�~�
phJ:h
�sv��hC`{䭗�����ঐ=f��%��1F�t�b���:��m�����^�xM�EȪ@_ti�wj>�I�\���M�TEn���i�$�i��힫|���k����،;Vm�S�Y#i�=�0���M9cք(E�U���oځ񤵭;�M;u�дQ���+ ���8��v!�rL�)r"j�?$���p�@S�m�yg�"� ���ۏ6���!�wF�2Rʃ>%��ט�O_褳g*Y�XJ�\rV�C
�N�!�e�:x�����&f�8LmZ�8���-G��)�e�Χd�<O��b���.�q�A�l(pK������A܄.t�x��� ���j���,�7.�X��w�0�0.[�b����D"�T��t1��)���n^�H)�l5n�BN1O�d8e�FDظ��NڬJ)���s��<@8����˞�kF恲�B\�8�B���I���5�D��K(��o�Ȧ�x����uw��)J)���BBѸ&J@9!]�4t�( AȠ/%1Ov� @A��*.�������9z�W�� �"BP:^ T8�s�\��A��SЀ�u�E"K�`�0�4�>$��#ʙ0����R?Y=�yZ��%rXy�V�������;Aj�+{`�t��H�ޭ*��:����W�kE���!](v�x�k��Ȩ}k�T�V�H���k' ݽ�h�:f�1$��(gCT�`��Ø'iR(c "��M;#,@�x,�b���gD�Ov ���x;4���oU�?p�]c�bȪ��'cҍ�Z���'\�S�|8��i�`P�1!�Y~���fJ{'lقUS�d�bN�=*���.�"}�)X%���#+����⚱K��(�=yAm$rq̀�,@(-K��@n	��z���4d!��)й���x��1[���~����N�.�x7_<fj� :0�;���8�@p�Ag�4CZ�\9j����'V���#�]�Kw�`KA�G0���9D���1�i��)�hȹ�
�,��#.H3�0\�B(>4��Yвi����F�,YͰCg�~2$��7�&h����;��8g J�-��i��T�X"m���Mw�p�B�xӞ6��J��# \ +^���-�R�NВG�.u;��?�X��,�#� !Yd�S�T`�]1Q�Jj�d�0"�i�.}��*~��c���
�瘁na��0bb�*��-*���0x�	���؎%$@i�2�Y"b���'X�kj��0�-��rv��|t�yd�D4,K�� ��<n�'!G�F��x��X�S|�Ql߅~\Cj�;/�V�ɧ�_`��+ձ2�:��B�~�E�EaG:�@%c�JҸ)���!^f��C��00���R5��/oUPqRA����A,�O�I��dX�W����e�'�&�!ajޅ/L��r鍄6q0�S�Nrv��w�G �d �R; F�XA��GxC��@D�M�4t<�k��pr��gDKE%�dĜ$8~8K6`�i�|!s"W;!F�Y�cǲgX���Mײv$~Y�bŞ 0n${v �j�l3�"�8%@�I�� 0]���)>i���M�S"�U���Ӆ;h๢3Ƌ
�LQq�X6M���	�(Ƹ;��{�|1��IC<x�]�"�W�T�Go�n�*�#`g^�/̨;�ITz�|5����q�m�Ywj|٦��@X��Ai��Ƞ6ᇕi͊���I4t��;��{�ዥ�ԫx�H�F ���e�f�X�_�R���)��m07j�=k��ק�$@�7��u���?Z�D]��h�����AF�#r��d6;������*S*���L(C��=��/n����J�r%����Qܪt!�wKT�TP�1�ߝ�ܙJP`V0y�^��@�����+ `��)u˂�� d�fR��q��5@�8�J��X�I|$�e���qS�)B�sĘ�ꠄF eZ��1!6E�6�j׌X���R�~h��B�Þ�a�1[�9`2E��,A5��@�� ��=D{�g�3n����B�������J�{s����X=/����!O=k��ā''�1j�����hގ��ċ6�
}q�D	�@3f +uAF�DQ�u��U's�
�X��F1SџL���L5R���] �0#�м^������)o@���'�21���Z	Jq椚Fd� }� �O�����'�(lH��IPG^.Q��hj���::�`�s&�OR#<��CɫX�ݱdqb��T��4����*QvY��k�@��iBu���c�h�g�L�v�%�Fi��I�t\��#W 3`VYq0��g�f�@��d8Xp���١C��h�Lz��B�E6	��5j�K�r��UYq�ڭ`0HP��I� B��(wLp��"V�5x�P i����:��A�,��X���'h��BPh	�3�M�bX� �+|�@ E|����b�ƁPC�ç��a���֚~U�d{f��4D8Lr�i��v��Ŋ7d�ؽ �$����e�p+�y\�P֣ȀY��}ȵU�	f�xB��5I:��e*Z�p<Q�iA�n�*�VE��0�F�i��P�@=�Z!1�)	"[`��Ȧ��CAP�T�B�����̌h��`�D <�R7��%�5a���"$E�D��)I�hFzbw��$[�����6|��&S2!A���$
Fe9%A�+@�乒��͙b�^}�p`��QΕZ�M_(MAȴq�N��
Bi!u�ܩD���$�̛���D���!�Ƃ�4�n0�닪f�螲h/�AY�/F ���*�kD��%�'6��E�Y/ƘHt��'��rЎB��L����'�
L�@ �)�&�ip��X_Lp
�je��Y#�B^~ԅ�Fl�)w�Ș&�7.���g�8h��RG Oib����ßZu���L�+q�ذ�;'5"�g��L5Ee�dOH<Y��P)W���(,ܢ�	�+�$l��J����>�@4�rm˟U�e�Ƌ�)W� ��H���ħP�  u���m�p����;�\*�5<Or��֊:�X"�'}�5�Ƅ�*?)����
j�Z�F�Z�hF�	��P+��f�T-e��=���+<�,��� "
~A�u]�+���GE/�	��髲�O� �5��u�&���8�0DH�*-E�z @��v`JV
�5&���4��'|� q�z�T5��_k~=�� \+���'�,�Z6)[�B�^(�O��h������-d���)��2������K��"�D�Y`@]Bd��+�y"g�E���#�X!N��8i�c�
t,�H$(�9x�%��ό<�y�'�L����%(r��"1�pI��P})8��􈄲n!�`�'�vY#ԡ��u��4�qG\�}�NP������N΢s����0��#0���q��(Fz��نF� ��"��LZ�qa�e����O4<"d��JM�nK.�ъC삡<���nq�.���"7��P㘬l����Isw�����TN1�t��8,���ne2����ȥM-�E1�B�?�r����¨��|�L?�Q�4�����,bA�B�&*D�@��+R\��ap.
�{@b��6|�,������ 꾴�WA�7'I���I	�C�mM����<P�t��01�(������D�)�Q8`�;~R�ro��{\nYꗢ�&g���A'�/(����E�&{#ZtZր/�tq�͸Ư��)N�i��J�'��E~r��}�ha��ҎSj0}��(�8=�pb�O�OS����ѨM��( ��)�$�'Pȸ�n�`������C9](|��O���E�K�����*j���2KR����*�� H�C�,Q�S�2�R�3�$��y�c�גt)�֊"��t�rň)c5�Q�1��1dp�x��,]��bN|Rq��m]�0�'6�-�nZ#*���5	de9��b5�5�'�D,�T���H�N�}SPѺH(Z�Щ;X;�$���3����%�3��U�]�娦 ��o�FBH��;xa��c�r�Y�hL���їfg
!�AĢ9��������3��?��ظ:PJ����6D`���q~2oڅ�Ţ��J���X8;SL��7͂Y�'_B����Q���R�fKX��ȓ}��%�*ͅ
<�`����7�l ���X��㘀f��c3��@ܧ��I�xU��hW�zC �0��M�P�ч�*@ a��Ȝ-GHD��#��P� �zD�?����$ �R�����bb~��IalK�v�!�LG(�K���mj��҂K�!��o����d,Z�Z^Ĩժ�g�!�_u}��L�hO �IU�F)~�!� �0��	�iڥd)��(�'p�!�$�(](Pip���)=P��I!�D���q6(٩���	N�r�!�$՛A�~�(�P<xQ��
�}6!�D0j���,ЖI�pXU/!�� �lBchB%?�B|k����x�"O0}(pJ�(d��s����IP�"O�E+� Q�_n(�`�74HВW"O���2�R�vٚS��8$Dk�"O�01�D���[A#�8u�ƴq6"O�I1���~X,9�	��&�N0@"O&�+R�ε
A�(O�_�.$:g"O�9.���1'�V�1��b�$!�!�$��pXδ��Ku��e"���!��ˆ_V��!v$�&�px#�O5Z!�$G
�y
7�.|�̑�R�0�!�DG(a�r��g`��p��Qi�ME:3�!�D��|���"t���5"�i��	&�!�$ֈo�@����;'<��i�kd�!��-.����P_�D��`@oYb!�d�5j(Ń�HB�9�,+��?�!򤗧-EP�`��AM1%�I�!�%��q�'l��k�>�!��$��e�WE�rg6!��'!�pұRg�1Fּ��O�21�!��W�_&b%k�A�&;Vm�QMǞ2�!�d�6t�ļ0w`8(�R�G��5n!��@�H�n��+ }�,�O��!�D�	K�ix��k��Ux�N���!�$��9`�����O$\�yK1l��!�döC�M{b$��|M��A�m�!�ĝ:Uw�,s���.l������Ń4Z!�Ɠh�=����5�I���42!�ظ��0�!�G���2�H&C3!�ʏ
OT������f\@�h�{8!�d����I����@����!�$�;ؚ`Bܐr�9�W�E�K�!�$�	^���Èn�du��ʑ(�!�^$G���vJL�l�xH����6w|!�D��j���a@Hb� ��B�eb!�d�9�x)@d�]6Zvj�Xs ٬@!�����ec�̟9~6d03!��!�dҾjHzRH��fiH8���	d!�D�C}x�36&�2,�h�6�Ҹ!����J��K�6}��á$=!�dS#���F`��j��4��!�z-!�$N��$���
�Zj.�x1/�!�)a夠RC��=b��I���Py�gE�}i|�10Ε"F�~u���y�,�)m�(�h'@Q%wH��KO���<a7 �%vJO]SELn��1����:�d��"O����J<<a&-�����z��1�>QR�_���P�C:�М��%.cZBg+F�P������I����a%H-��O�`���g_>�mC��ˋ��У���?|�6.,�/.�3��&�𵱵/T�`q.�׆�h$�ɭ|�<	�C�87�nM3�퓢Lb�k��Ej`����"s�Q� ��UV�V� 8*z�yҀ�TTa/M8t��be��Q�0D��锝��܉�.T��1E��[�D��ӝ9p����W�6@���O�\�%��/�~´�K�?'VH!��)�&U`E����^�2��
(��!�R�J�@�I�"H���݀bJ�#2"ypDZ�",�`���؏,�@ip��҆E���������}SU�[=<v�����J�m�,9�ÿi�N|��g�Z�]9�=O�Q��J�~p�D�e�a��Ub��5�GƵ��=ؓ�Z�p�㖧\vv|+�M�ßt�E�:xI�M|�>�R@ǯ|ސ�h�E�/Jq\�Z7+����O[������]�p�@T��κ���G:.trM���;X1Q ��Y��� .SUP��1��9������]	L�*u�Ix	l�!E�-K��B�\(Zo�	���H�1ʆP����!t��F/��hz,�7I���J'��^f�%��
�3Ƙp���%r���ק$p,��jߤ-�Q�� k�����ҭJ@�D g��IYt�FkA;N$��u�].w�PR&ᕞ�P�rb��+]���"G%gJ�Q��)"��ʅ�'�DJ��͇+*4A�F�}�&@��I�V��p��BR�U'x؋wh�%;2��xE�/ ,us�<z�>h�c#��W��n�<N@PQ�Ӂ�5*}�i�Cm�35�"�d���?��7;݂3���}"(�����ú$�8�fX�h��%i1��)>�Kҍ8b�a�vH|�1&� �	���]2wǢ@3D��I�? ^�;5:-C��u�M� ���Zp�ĽV9B��bd��ݨO�h#�,߮�R�5C˛0�(�rP�/K�M2+_%oɰ�aj/6r��D@&&��y�&L
�2�*�J#�,K�}R��<!s*�e�j�*�H�:3j&�#�ꓫ7��tj�&Y"a�P�Z�D��vc�D8W�զUh�!��^��'e"T��X�R~o|E	AeZ�WZ�2�H
f'"=ȷ���?�W�#Uq���h�<֘kb�[!A"�a+
�C��=Qq�L�#�:�|�Di9C��2'(h�qW�]5A�L��^�y7��9t��� �<$v)`���5E�v=�S7O4�!�� �L|kL?㟼sR)d�� ֐ �(LC�N����#���!D{�z� ��M��iݙb�m�#>
t%Yp�C��ʠ3�H�2>^9�G�
�>5.M���+6��ys�T�x���Ge����`��P/��B␮K�)��Q�G��?�?)��	�hz��"Z+��CA% �`q��n��c��$���WHI�C��n	�╴]�ֱIA/�m�'+�y�UH��x�$ p�E���To-E>R�;C�\ AP���,e���	�)2��I	 �ſM|�:�]�4/j�2��CT�G���^��2(�Շ�Z��M�A(��U��j��[q|��,�d?��N���c�-a�&�'.��K��|QH�ۢ	Є>�HX��R�a�2��:.�}��*���ች�XD���&H>�u[���91�&�Ʉ,��E�D�ߵ]����g����O
.ٺ��:u�����!��`�@�S,9��?iRf�?Q�D��E�x^���7��X2�hĮH�Y���Uc��A��;�-2��|Z� �k�����)V*z�@4�t�'�Qs��B,i���}z ����X��7m��w�\�	t�	mF�x ��:|֨L+Ǭ�E��� T˟��'-
�v�^c>A��e�;O����5Gb��EIR�._���� (<U��Ď�: b�6�#2��I������$�9b�\&QѺ�C��&c|TC"m�#��u"e�<`��|��u�'z�
QH�PPy�5Hw�m���R��Qe��F�0\�d�9p�"AhՍV\QD�C4Hv�e�CW���Mj�T��a�һ�@�@ [�*�+�K�'� �3%6d|�;D\���	D,�3-B
'��YytŏiG�}�`�B3�(�`�,�GZ�Fݗ@"� C͂�$��MY$�ƞmB�͕w�P�7 F~ ڢ�dă��1I��Sj��b%h�~R��I2N��!r�ߨ[�'.�@ܾU�
��@5�V����ճp�'�X� dHƿR�"�+�N��
��u��]�,�cj�i�D��B�\�-������#:�D���)�)*l±���'<&(�#�Ռm�P���杫)���Pc�;�R���+�4s�:׍��=羐	T荛/��hs��³r�@��c���A�����]�nO�U0bW�nu��� �lX���I�Kt쪠m C�� �m
8yՊ`���gAuN�C��$�í�}ޘX����9H��B�(�6�r�I��"lO	Z���:��a��iPM�@i�#u���q昌o�<=�@��'Z�0Qa�8k���)��G�P�I�"v���ц�i�*�ई�}%۳L�=6L�%XB�O�Gfd��>��@Q]���N0Y��<� ��?���o�@ʈ=)S(S�"N���4�L>f�t,���2�4eBd��H���K��3[�	I�(Ҵ$C����{��.8���T�t�:���@�u)ͪ��B��Z{�ùs|S��Q�,�kq/��q��� �k�H<��!лK�8� �8>�҉�5��#����HB�����c�](���S#K*�b�2��'ǀ���o�1d�H��6�Dc�Ti�)O��:��Z�@�}#E)ǲa2&�sAٮl�y@!Ę5V�`�at���Pf`��@֖
�F=���b��� Ɔ>be����,-��:�GV�:�~	I�W�z�iR��6%��q�*�C��8`UH�'FFE+Ҭw�H1X���Q�t�A2��4!��Z	(��Iֶ��kގ{l��S��̀ z�?�bD�B�I�D����0y7�.N�Rt`�5S�n��t\�!�(!���Ԇ{������*Hx��s��S�h�Be��
ݱI�t��Dg��$�8�	�z��	�t�G(M��* ����F�#��}�l0�Z�����fK�P�g�1O��!z�^
�R�F$�~�b(�D����-��h����+���Wo���yr�X�_���	9q��5�V`�����|����� �
i��� ��Ǽ6İV�˸��d�V��~��C�gz���kJo��� �Ǽ3Аs֧
�B̬hk0Ɏ�o(=qthS5X��+Ԍ�7��L�F��C�<E����РM�t	çN0,�&��G	R#Q�T,q�"v�~]�'�~�>J���"<�A7�W�z|*���)�U�^0)A�ӟt�|I�����npgګ>�Ќ:a�n˘T���FW�'ft�qo��<�J�
f�1K!��W��q�D,NΠiu�Ľ	�u��	�*J��4��U6J؛��ЖZ�4�R�4Y��EZw'��ɐY� �: E�+�`�C0aV������\�bݱb��; r���X2k䐐�%/W)�l��aW�)�vn�^�`ݭ1�
y�G����T{���.��Y��P�/fЋ�*�5P�֝��4!� �Re��}<HM�v����E�`�vʃ�?l6��ǌ̽_�@�KA�o���g��V����ǫA.�`1���,}���20�z9hҵi�Qr��@�r�i �U?~��@�%v��i׌  �Nݣ�H�$��'�9�tN�؆�O�}�%"���'�}��M<l��h���P����y�(7jn��˖���n� :w�B\wi��ӆO�]��@9P��K�n�	��l��p��?I��/]T� ��[$j��E:��Y��¥EˍH������h�A�T
\4�ɰ��ܼ>`J�mZ�\"�B�k��M#'O�{$�S=R-z�H��S�v�ʠ���B���EVP�r�1ݴZ�ē���\����P
T�=���ቼ4T���O
�
�@���'Zr�J6��풐/[|�����W01���_-��e�7�iR�:V�:h4�ᛥ��w�ɤ/�x����@R+��镮bH@ꂬg�T� 
��S<����BK\��R,저���,f^P����|/��U�4���XU��q1���A?[��Tk�i��W��F|"�a�^4�F� G�.]8�d�0*I:сgkA�h�Zd��O��䓞x� �����C�$Q0޴`R�x��/��9T���<�$�	᭟�z�(!�֒��?9gj@?S�I� �T���-�%k���87%]��^1�p���^�$6햚$簀�v(#���O��,!�e�6
�4���Θ!E�ܲ��@=-O� z��H��0���d�#C����@�,M��'2j���=eu�8ⴢJ#|��3s �����#��	!J,�t)������b��|��O��uGZt����%�^'A��+KPt�iY��ۭ]t��QR$��P���e7����u�_"M�KK�
Rrni�tC ?$3�re,�+M��:jV�H5 ��	�!�Ȉ��{�? �=�Đ>eظQ�1kW#���Ui�jG �c�[�~)�q��_����ѽc��$��!���ɘ�hB�����HBܓ�I�*��4���I�?��I�n�&"�A�d啎`x���C�ߑg�t�����>z�Ρ@T��N*S,�;�,��	F�Pi;�DС0�r���i�y�ıXt�7L�'2	�ѥ��q�igC�.Kd���S �Y�p#��[t2r�$�<")�QE
�s�Q�C�,Ol���c`�0.`ZsG�6֞1;֯�(Ew��	��B'7�1�M�0e�>��'m�XˈOr0(C��3 ��Y�j]�M��Eq��6μK�������(�p�`�3��!�JݢL��a97O����T�͛���ңE�L���ؼM̜�ѫ�.��O��g2f���:vj��T� �I͘m�b� 	����熟N��Tl�*	5�Y��S�g�(a�ȐMx�M��kN���\���҈><�ѷI��O4���j��W:F9鰡T�lPRs�қN�`�ieÐ�{6��V�F����m�5'<��g�-k�Z�xt�K��XR#P�q �↊�B����M4#6��� �7�X�Bl�y ���.>;\\9 �� |���pd�Y4�J��ccD�
��G/��Ff�Mxs,,:<VL!  I�@J�ԧYU���@�˛(8+�$�d��Np��U���������JR�=�T�:���Pg�ͤ,U�����[�L�ؕكJ�tV�d����>L+�Y���?��� �%�.U�������z�-	<T��Ԉ�����˒8ф��鉍��O��C.�N���R�b��y�+]�q�Y�E�(=a&�.4��:h�!yT�R�c���'^힠�!ِA�<{��͛t����5"�90KL@�ŉ���<)dC�3�1aGKE�vk���&CF9��9�npi��eؒWb](�̩F]��;PN _�%��3�̘r�%�?��)�QEY�RpyxS��CT���n�O��b@1ǖD�s�Jj�@�4�A(R+4��,ȶ?_�l���"M9�Beb�0��U58P�d�E�N>�ZE��g��xq�$K;7�U�g�Ӱ8?�!(�o�B��CC�$z�,-˃�c����%l�o�01K���2[�́��F^��m�n�E�>��.I�.�~�����h�,	3��B2Z���BkZ�艺��9W
t��̃c5�٘��@)hx��S� O��@&Î���b���jo�KD��*�mۖ凘rKb%ɶ˰F�X�:!�4iTl�AgDV�n`�4+��Ī�eˆ�G�pNh1�$�"/�Va$�Y�g�Fqc1Ą�HO��I���E��*E�V1J��� 2�N�$+}Yâ�(	ְ�@$��6r�4ر�N3 h�� A9�I����p��Y��W�պ� �CX�0y��W�`!��;:uZ��	�!@+<yh�E�O���c�՟x��:4�R�x2������ϐ��2��G��4�B}:B��'�40�e�k~�y��&U�%	�H�K�"|Y��Ƨ�+max���;��`�'���M��+�/$V���ω~R�����_$<�<�Zre��?��H���� �i�#k/&SW�Ȇc�5R��R�d V]I�	]���x����}�X��nO Q3�iBӀJZ=��1�'�8�� Z��0���uCI� }�H��� P2�O���ܡ`T��t�B,6�Nm���YKx���T���7�He���O)���A����hG�]�rh��A0/ڊpdϘX�bh�5�F4l
,�2���C��?i��RkK$��� j�4	c��PܓM����i��(���m�a�,ULH����ح>�
�� "��u�(�*U0<�����>%��AG�'�ɻI�)z،����@2C�Ԡ �O�)�A f��Y1�6}�6}Y�o7�x6�Q���C�u�t�'#�k��A8D� #3]!�d��O#&a	�n���`A��S)|�B޹l�l��,O�X*�&��I�(�-��e��b�j˼u��#`�ͱ=C*��aO&�O`�BÊ�a�=��&�r�<�	Q:8vl�@v \1Jo����j1�$�83H,#0�Xe�'ƪ0��Z�%3t� �ӥ8A��b���I�j�lm�'Y.A�C��̼ ���k��]�u1���E�u�XP��@Q;�0?���\)���_7^�NI	@r}�h�$v��¶*˂^��]���@��uO[.h��DRH�
�G�&� �`�~�|�ȓFf��P�_��X��k�'~"D0Ħ�����.�z��e�G�+1���"s8�	�O,��0�NXTz����)~������H��h�.-6p��'�\pI��!ܾ\��ݲ��sz2����և^���E�8�$��	kSiQS�ؑ�R�� $�6�G~B/I����.M�_t
4�4	ܐz��a��8F2z̚u+H$a��*GJ��D���{4�'��t�6&e*PQ�vÑ p��O�${�[�����ƑZ]�IS�A���E��h �D']J��}�plݦ~�X�b$��'�y�ɐ�W6�t��� V�;�$�(�Q9U2�4�r�
g�j��pOS���'�"�H�f}�DTyO�i�R\:h�j��H��?���ԊzE�3�ti.T��I	"�ґ�O�4+r�a��B�K�*�"��1M�"?�Iɤ1�v��񍜨K&�� �H�r�'��Q"�q�"��CD� ��ezb��0(�6�#�'�X����@Q�<����H3�OX����K����/J���֚�<3��(�¥�E�U�_Q�BiS3S��c>!��nҀ �\��)[����
��6D���&2;��8XAmD�a`� a���<`j��dɃ�B�&fʒ7j��>	'�`:vH�>kӼH`!"��g���@�;4�,�rEP�K��-���;i�8��ޔ.U ����'1�q�2��r�Pu�#��
A v��'K�i�q�=M�@�*< h�'+r<�����J�^��G���Z�'�\`Ua�Tjͱ{R���	�'�`�SC�݆!&hyԢ˹u������� ⡀qm�Du\�!R��5�ȼ��"OѢ)�����ZD(�%;����"O\�c�KR5C�1;3���U�*p�"O�=8�W3A���
�P�$�u"O@�8a�]-eH-��n�e/f�G"Oz}:�`ůr���l��[VT�4"O$̚c!�<�DAQ#KU-�ʡ[�"O��*�;4|�\���C�]���k�"O,� �!��B���0E
�b��K�"O�բ��L��h��  "Êi��"O8JV�"#������Q&ǜĠ�"O����`�'5���В�	�x� �@"OT]��b�`�r��rFݮj���;$"Od��v��G=.I�ԘX� �b�"O�PV`,�\q8�mӫy���"OX4���?ךy���E	� �'"O��`�	R<5 �s�Б8���e"O4x�/;�(�Љ��9��"�"O.Xq�H[�G�d-�3��5���8e"O���Z{1�XJ�iF�V/�m�4�Q �Q�ĩ��;�	��#N&#�1O��W�S�.��4�"��f���"O��O�]H,� w�Q�'J((�����]<�p�^'�lIF�CW���y��C	&���e�i�Jp`�
������rRb��!��*�Z�S���8$^U�'훖��e/⬀K�"}Ҁ*�y�R`��ʌ�0��q0!���o�3��:3,}���|���'n���j�o�>fy�d3U!@"�:Y�6J�)�y���p��'w]�C,O�#78�"����Q{�'���=~�çc1u��jY�z� z!c�,k��;S��b��Ya��)�'5b���*,DB<�3iS?Hڸ�e�1y��	I� �I��E�(B���h��x��nW�`�1�̔���Ġ=�t!�G*ƞc�N牑*y>�O�1�C�eR@iK N߉��1�TmQ�c?v<Y6�'���`�OZ��0|ʃ�_=%X���ǃ�UV�t9$�<)�����	z>�Sue	C�Z��ᓅL8��XS��9P��	�E� %�b\��54�e�� [�XB&�vc�+�L��:�	�~Y�X�T@ǰv� ua�D�.c���ɕLa�D���.\��휌G�|I2��ڋ{Z�����~�k��<�3���@�5�ޡ0	0F$,�o 9�O�	��In $�����3IO�S��R8wc���D1�?SeZ4�EiT�WМ����C�IH�DX��ɇ$��X�A�?.BC�Ɂ6�T�;&�2Yj���Q嗊V.C�INѦ��bE��X]�$�S��%FbC�	 5���J򪀞V+x �6	S�\�|B�I�/[�	�`�}�L$Q��/U�B�I�B."M�n�(3���E&yg�C�	!�*Q:�ƽ�	����a46B��&4��\�����@�� ����-'B䉦������^�A$`���^:N�:C�	3ZT���b�"MH��!�"OC䉟y�0��'��ډ� )�e%C�f,Y�C�"8�Q`��U��&B�����vƁ1k�4��@�	{�RB�ɣ.�"���W:{9se����\B�3�J5��Θh���C�*,2B�ɷ��q�
���>�!¦��b��C�I�6I2�.S|^,- $�E�tQ�C䉛-�x���Ɍ`��x���Us`�C䉬
m��ֶ����Ǒ{�XC�	.y�f鈆o_�h�|4��D��RC��'#��)����v�A�JB5 �rB�	�QӪ9�ʐ�.�*X��j�D�4B�I8|*u��"WXHh�Ĉbi`B䉗M����aP�'@\�3�\�A^zC�r\j�y�,�8Z�H�+} C�	/|jI9�
��[E�U���[�E��B�)� �E��uȨ:�oW*Us�|k"O&�S�%�7Ea��1H��;p�sb"O��!���+�p�B+Wc�;�"O���I�"%1�H�ATC�nA"O�lB ��-u����/	0��'"O�J�È�&胰��7�x���*OUW���_�֠ 7��>��|�'���!�.����4n�x�'�HA�3Z��h��ň�:\~5��'�t� )kEԹ:�aИi�'F�����,�����ӂU{��	�'J~m1�̌�1�r�Zm6\�( #	�'i�,S�dRbqҡ�a-b0��'lL�4%�i���a�`@����'4ޜ�`bK=/�0|��Μ[��e��'Y�����ͅ?�����T#�R�;�'R�$�&�_5}�)��ċ�b�̽�'�8U��O�����W j�J1k
�'O`т@`�6ak�(��O^�u�t��' pY �·�M�P1�r��;D"�80	�'rU����?x|q!m&M�>1J�'��Q���+i|I{�Eޏ�l��'{�!�IN��T$x�͉<KT�+
�'
��
��_/]0&�zD�(;��(��'���S��҄e��$���.���p�'�NxC#�P�Y�rAda��^��*�'蔕!�nX�IL�!9��N�V��
�'�:X�G�D�d ���8�L{�'Z�@�]�QT@�3�Ԧ1����'�L��7eƕS#��'�Pe�'L�"j�0�Q8�gd��j�'��q���v�|Y �!Y��'(�TJp��JjE(`�>,5��'�>���BT'P���HG1	0�=�	�'��ءKѴmސq��F�8�t�y
�'�VP�U���<h�y��� �U9	�'�x x����$�ׂ�/D��B�'i�(!�����H�tI &k��I�'a~ ��!��5�|�2�f^,o���'w����U�z� �PF��b���'���P��؉u�F�ڷa��!b�'�LQ����'i���'J����'�P��A��L*��b7#0:���'�f�)�%vD��F��#+�(X�'��]J�ř�b�"��I��P�b�'�x�hȺ�=Ib��V}����'r�	�C�C�\XR�͏K���	�'���"��ԛv�`� J7-餽H�'����m��$]��(M��5SL\��'zH�d�Z4wJ"�b�?1k����'�ځc�
,c�PjV�����:�'PT���l\<Ђ��E ���'����Mۮws� ȢM�8Gd�h��'t4��U��9�uI���$4an,�
�'h�b�32���/B�%ܜB
�'nmA�M�3L❡�E�2nց�	�'���!\fp9�oG�$it�1�'�0�Z�n���>ˠ�C�@���'f)Hᯏ:xe��ϦX{*�'@����!B���żSn���'D8}��Ȁ+���d!M<F���1�' 4�b�ǌ�aƖ�*�V��t�'Ϊ���N��q£㏢�q�	�'B���˖	T�)pS#�'_|0���� ��Bu��z��$J&��H�j"O� �S�T8yV�����8��AA�"Ofa ��/�JQ�.o��"O���g�PA�����j��uԎ�	u"O&YK#N�7$�4!���]�x*X :�"Of�A��;d>, Ux@ʜ�F"O�`Z珟�V�[Ag;n�;�"O�Qi7��(.|��QG^+~\P1"O��0�K٨;���q�E"TU�%S"O|�*%�٘��� '�}Cf��"Ov��|y�+�lY�U��"O����������i�PSb���"O	�G�˝t;�x`ÂM�%�dm"OD���SY����#^�L�[F"O����K��t$��h���*��B"O$Ա㫌D���*t��ظ$"O|q�'���r��4� ���8X�"O"��cU��b���חX��Ȃ"O�����fsR��Ľ,fR�( "O����h �u�,]��M���<1�u"O=�7ː,&*�\�,����t"O`� ��::Y����Q�b:�"O ������nZ���ʸ}�0Xq"O��i��Nڤ���J�\ R�"O$��Ek��,���1mŬ���"O,�ڱ/��X^fm�6%@X�D(��"O�T��Q�*�ZN��QҌ޷t�!�d Q�XE�Y�/0�X��	;F�!�$�X�h(�SA;�"3 Ꜥ3�!�DI�,4p{�c	!{��mp�	E|!�$�T�>�:��ۮh���r5�Z=jJ!�$%3žp2U��V�P�xQ�/!��-�F�h�	��Jy��Q"]�!�d�9
���-soڴh� ��!�DϺ������ݾn<�*g)��!�ʘ`=Hi O�>�K�i[8J�!��Ȏo�����%�>a��'ꚋZ�!���'2����B�>vN��b���!� 6e(Ψ�#̊mz@BUɄ�>Z!򄍶t1N$�4(^������@!���=R@b��	8ԣ"�E!�d �Y�qEߛ3:|���I�!�D(v��[�ӈMw8m㇎�5�!�$ I��XTKE�� E�3>!�d¨�5�FB��
�)xDm��;B!��=sQ:y���3&D5���ͦ"D!�d_u�t�a.�|�`
�q*!��^9l�v��ЎfZj��AL/!�$\-NPxEq�(�v?�djF
M!�$A#9�X�v�[F�Qr�I�~�!�D��*�"P9�
�>2�,a! �!�D�5=
�N�s�(�sc��!��U<#�8����J��1��e!�D�0�(���.��"ёT!P�]!��f��@z��X7w���.��D!�.�p���U����ǭM�G�!��3v�4)D��'=��e;��ݏ[�!�Ė;;Q,P�,W�Co^�s�늍_�!�dQ�{^ҵ0�Q�DjJ�@ǀ	�!�.F�^�8ON<6i
Ѧ�D[�!�$�&��,�2�M�3SV���i�.�!���4C��áCH�5d�1IU903!�dߖ����'^��|#�I=.(!��
 `�&H6+4M�.�"��̬! !�� �<j�o�d~�qҐ"�#@�x9*�"Op0{��\<��	2Aܲ/�:�Ӳ"OrpR3Ǚ�ah3��/A
\(�"O`<�p$,'tE��0��D"O(�;�e�"��7�����"On4�b	�S�dXd �(~�:(S�"O�1��Jz2���O���BȘ0"O�d+��N��`=ѦNҀx�h�!�"OJp�3�R�x�d���m����V"O�bψ)j ��c�Í^��� �"O��ɁD[�5�؄���#�8X�p"O.<h�
ίq�ҕЇ�ݒi,�xC"OH1Y�I��\DCd�L
Fu�ld"O��a���t=���� �8�|SB"O>�x$ո#�$c+K�[vq"O2S���.� P#B(ǜ��2 Q!��[ $H�5
���$
�P�`%[P1!�d�(~���g��S���:�\�?!��]�F&�X�4����@9�Ȅ!�Ā�x]�$
bۺXU<���$��!�䗸Zq��V��{MH�b��N$H�!�D��Kv&�X��5lMLK��@�!򤊸eaJ��� ��m_XI0�O$8�!���(|;�*��	E�][�)��!��+����?�ɓ�J0D|!�Z5n�6$�C)�p4�!���7p�!��_(�ne�wlAm��T�F�!�d�%eȢ�j�$�,ugu 3I�Q)!��ӏG��Y��U� =��鐂AP!��\��x���(V�|#e�7�E�>!�ݠ^2�Q)�
�BoP<А
��!�Ė�'i��1b6�!T% �w�!�đ�"|C�(S�X^�@#+H$+�!���g�|�%.UWJ"��K��!�;	Jȃ���<<pE@Ë@�c�!�9?��̹ �֢q/�h)0����!򄎧�1��&Y�g����Uf�kt!��,8��@���.�v��%V�!��L)C��Ej��ۓOwt��R4J�!�f9�qK�l97t� ���|�!�D��lY%��o�� j���|�!�d	<��R��&�8���<s�!��^��f��'�T1o����qc�S�!�P8�(i�$dN44j��[p!q�!�)izp�iQ/l��֬��o�!��U6äa�QC�VR��A�=:�!����:�턌A���G�!��0&&�e�W���B(��ϓu���4p[���&$���� ����yBȇ�L @  �,�tZ�"O����bɻ@s�ђ+г � uy�"O�)����B�(�A*��I�<1T��� �l����y���1�C�<�w�D��(p�D�G�~���M�~�<���ەI�X)�R˄�"�"�`��Nw�<��b�<I2r�)�LV(:JF��Rh�<��'�U�r!�4%�*~����i�<Qc`��@����S��#?�
6�}�<a閼^� @+&����\�Iv�<���Z6`�Nܱ� �x^��aMT{�<�炍+���k���s�h�A��x�<�"�)(�����$@%/�P���w�<�b��9H��!q��8d<�	�nZu�<ِ��Xdn��tj/E/��ağn�<q�?udyr�A��j��#�Nm�<�O
0n^
[R�R{�'Fj�<1�E^�]���YP�QfV!�ǂk�<��k��t�lQ���!m���g�<��&�U�ɂIZg���^f�<1��_MJ���~<�(���VL�<!�'O�����i�)�|$+�GZs�<�F��%ݜ��ϼ\K�1�C�^q�<�g	̙G��J3>����@	��y�G��	��$�5��H����K���y"��"*����Z�@xZ��ШD��y��	��Ԡ�O^>�LY��M��yRf�
�:�)��	`�)�!�y�(3Ĕ��d� ZI�����y҅})iC
�x7�����}�j��ȓI�\�隩 \��{��_)��U�ȓ3� �ЇI�F�LA	U�9q̸��i�H�E���;缬Qt�82Td��ȓ
�`��)I:\� ��AՉM�U�ȓ�Z|�g
^I��`�5 ��a�4 ��Q���t*�x��M1!�@�
_�ȓO%��+�f�%?S�u���!J�؇ȓn�|x���&f� ��#Y�<:}�ȓ3�<�	v#WJ���`a^�-�f(��;��� !��pw��YmU$r5H��ȓ����l�d��x�����X��m��k�$�2a��QYw*��BY��v%Ve�EB)A<z	����L^X!��H�4|�U��9a��M���@#y��D�ȓWJv9�ҥ�_�]������Y�ȓD!"����Xr�9�!�( �ȓ(�b�Y�뒪%��őT�H�aVh�ȓ>v8A{���3<!�!K�l��хȓ7����g��*�E��'��p�ȓt0& ��|����#HV���1���Q���x��M"~bp ��#�nXⵌ܃8N&�	W� ����S�? aa��1R�؉���O�C�"O�<+����yzZ�HmW��)�"O�E��/�� Ҫ�����!�C"O*�Kg�_�~�إ�KΪ��"O�M��D�v�x!�N��9�"O�}PqH	��tĘ���S��<("O�-B� ��q�P�=8|��A"Or�Xq`�.g-�ar�+Ө))9�"O�T"���M�`��jV�S
�L�T"O���a��mW��hA� x`�	�'�j|��ț��� 	G9���`�'����$I2rA<�+�ǚ(dly�'�,YG�X�z��9! 'tZhC�'�䵂!-J9����\E��
�'T�ݙuK��1'�=H "X%[D�D�
�'v^�h3��2m�4URTZLy�
�'�pM+�œ�H�$�lZ�LZ@��Hɂ��`�*��q�FjQ�/j�0�ȓ]�F�G�*� ��t�#\Xlԅ�8U��A�-�X�@���"R�$���i��)��Pn@�h��Í��b��ȓa�XI��^=F�X!��E�F��ȓD��)����Q���`��[-6��YD�����L�~@b4`A�Z=�ȓ0f���I�v`z'��>�R؇�O$5����'3t��4%K�o��ȓV���;�N�(A��1��R�P��ȓ/Nr��ԦхL���WG^�( J���l+Bu��ɮ?�����j���QD(�Go�JJ2P�0Aۋ�v�ȓLA�9!����l�����ă{ANL��9���(܁f�����`�)&�P�ȓ6.2!{�ى!L��Q�G�$�ȓxwb!����6
p�@�(?V}��?�F�x��K��^��c�%k�|�ȓ$%�<��Z"�<�7DV�*d��=MY��X?e����v�����8#p�v�+r�R��͛�������($�&��4muh�q�e��G%D�px�&��H�x�j0���B�Lmi��?D�4h���1c��		��г7�$�§9D�ty�I��XB����&�� �'7D�T�m��L�@�Y��>6�2L�T�)D��1��Q�B��9A�J�
sR�$D����V�N�8R�F�V_�}�v�%D��āN7{�V�
�t��Ίq !�zy��k*N�Hs���5~!�×3S�=�E �4=��TXD���:`!�C�Z�8��!t��,kaA>G!�D�"f����2D��q��Z��W�@!��)w���EBF�"W�1���#9!��N�~���pM�Q��#�Kp�!�dp�fu�p�N�t�4e��!�$��T��ت�bZ�_,�Tk`��Oo!�$�0z�b��B��A/����ĥ>�!�$���٢3�ƵGu����:�!�D_I�8�b�Kt6DSBU<!!�U�H��4����q0��'��!�(�D���)�'V�������!��{��e3��>"k���GK��!��j��sᮛ���q榈��!��?"�� �q�׬R�
Y��.�!��*6��vK�6��� Bkc�!�ķhް��� ]?ܚ�Ij+!�� ~��%B��..��j����(��@"O���[�* �Z�	D���c"O��@�%��c��B�*S"y&�5��"O�@��9X���#ɵ>,��c�"O����\4�P�A���3���"O��Pr�[�J�&IC��:>�p���"O|h{c�\�h��rנ�7+��qkv"OD�#��?e�B<��
Ð[��l�"O��Rg9s5�<�s,� �|���"O�s�	=a�YQ�Sf�$M b"O�䂲Ni,�c��u���"O�)�l4/,˂��?e���%"OZۤC�*��Q2�MOXIW"O��1��C����s�I����&"O����C�r�*�sv(�yڲ1��"O�����Z�#�1�FB#2�^5�"Oց��E�h��T&�)�lQ�w"O�	j��ŷ3X�{�FZ=���U"O(,bo[���N+l[�X�WJ�=}q!�ӥ>	�I<6V������n�!�$ŀ=,4�wE��T�Y�(H.�!�D�3M��HgH�V�0�Y��N6i�!�74�B鉶�\�Py��H�_u�!�@�	l2e�	ג1�ĳ"	�o!�D
��2�C��S5tdp�4'�8?�!��"#����ܮ�\�S��o�!��Ʋ=D�|h��T*=� �(7D�ar!�~�-+t��ق�Jde�+U!�-Nq���ā^7K<�j,J
�'���A"Z���WI�	z�8�y�'b���0w�=�"�F�jnxe��'K&
�&�93Bm*^�8ݪ�'�`�C�P� smB�\˪\��'�p���V�~����]�&s��)�'��+���xՊ�<�8��'4�K��$?C"����Z�\} ���'Q�#����Xb���T��x�
�'.00@d�x�B� �?2��
�'W( �ǩE#'*��kbk�DS2�9�'�;��HL0�Bw���>��y��'��(�͌1]�L(`�C�=�nP��'�q���/��*���d0l �'�� ���8���%.�
Ybt��'j|l��C*<�$�S�J;X�$���'�6�bB�t#��I��8b:J=	�'�  �.%DUD����8*��4k�'����f�u(Q����m9�!��'��[�J�H��i`�A�l�*���'D�!�B �T���	BJ��v�(|��':�ٰ�Ύ�(�Fѵt��Q	�'��a"�(�c� 1J�H� B�~E��'R`�HE�ΑvxP����"��Q�']*%�h�0f�j�J���;~� E3	�'0�,��Ka@:���o�f�!�'����,w�l!+���2v�2\��'[�q�% J�L�jԂ��|����'J���Ԏ�K�f�8��N�m����'���C-�/�c0��^V���'�,���ߊn��Ġ�G�QxF�R�'phA���Bؠ�ŇC>~�!�'��=�4���
�o��;� �"�':vTk5Oz��� F���1���k�'����� Y�VN�y
�;'�ld��'
\`�����$�am���Ո��� PU�%���^ �e#���F$��y2"O����NA"	��1�g�HTZ���"OX�ط�6+����t�Y�[�\��"O�p�Q��B� 
�V
�L#r"O�0�Vp�L�k���
u���q"O�l��	L�}"dp��o�I�^x�g"O����G�6�@�T@��k��3C"O�|a�E��XzNE��.
�bab`"O�eS�ݕr��[�JM�:�����"O��å���'�tU���=b�X0Sp"O2��ݖ)�ĭX +��O�P,r"O�����dZ�Ăwj�<T㰘��"O^Tp)�%4������*��j�"O,x�d��?�<�@3�@�F��IP"O�$�ʃ'_�I���)fy:S"O�Z!��`Ifx ��;k+����"ON{hF�I$�A[�,7�dJa"O�,�W:�\�РƜCK�YBF"Ot����F	�.�2�O-G��!�"OTi��ŅhR@��҂qR�1"Ol`��	i%K�&��W �9C"O�\����A����%�_���A"O�q�D,(8���XqKƇW����"O�%�n�1��C�IS)���P�"O�j�����<kP(ک/�| xc"O��E��|;N-q�N �!@r"O܄��,�����
±x�"O$ٻ��
�)�M� �[vd��"OԸhc�!/�@��� 'e/�]�2"O����ߦ[��'�V�[�"O�3v�&z���7��:�h,�&"O:!���E���N�n�pt/�!�䓇_�L�R��K��7�Ɏf>!�D�HV�Z�H��@��	{�N1!�$O�Sw�}�v)�:UbV9k�-J%�!��ޔY�0��e��d^�U{���;I�!��]~>x����6k���k\�	!�!g:�sԣ��H�L�Rǜ	8!�d�H�� p�N�>��TE�,@q!��¬{���`���3����Y%!��_�W�"$�\���dӗgW!�D�4JrQ��aY�<��i�J7qr!�dW8}�@5i�K�$��:�ȱ�!�$D�Z�򰲡��'80ZdAu�ʋ\6!��v$�1b�gɛ[�X"�
^!��p�@�@�%�+�M���'�!��Y�;Ѡ�P��*6���h�!����E,�	]�(�P'3)!��·7r�D�tH�YA���p��[@!��G� 调c�y6
�BT�X<]*!�p��J�LϲO�A2҉��.�!�Ɩ��ׂX�:ƈ�Ńq!��Re�mr�M��m-�8�mƂA�!�Ā2X�4Ai4(JtQ�0OΏi;!�D�5U������@�D�Y̇1�!�D3L��Y� � �N�DD#�N�$W!�dS�j�`� �I��L����ʏu!�Ğ�n�x�#V@��i�_p���*O���G��5c���V��/E���'��,��cK�$�j�jV�P�<�֝Y�'�`�"FDBG����ɀ ^F:	�'7�1�s`�::@D�\xr:	*�'�̌����!���1Ԁ�y N$p�'ix����� �D@�<��:��� .$+'�tw�e��DvbV���"O� �@(LdBZ�Pc�F�]��"O��A,�-E�\� �� 	BB"O����덁0�8��@NHuV���"O8Ŋ#��P����OA�u�0s"OV�Kc  �R��Q/Dg��4"O��T��`�J���F�K��U"O� �j֘aD$�����U����"ON\�����<(�uAJ�,d�G"O֬{�֗�
��fJ�{f>x��"O��Bt++YbzDTD�
0[�(��"O<��WK��Qzu+��Sm9��'���t�\�^m؄2%�6[Uր��'�NĲ���pt2"�_A�D��';��Q&kZ�7��ˁE�J���'�X�CC7/q����
�p����	�'�$�`R�Q�>��i
3OfY^��'5�5hU	�[´Q�B� 0ZF���'��0c&*Z�P�Va��'��W}"��'Ԁ�r�NI$2��y"�`�D'ƅh�':�����אL�h,��B�<��#�m�<���߷��{�E��P�6�釦h�<a�k� tc8��ua�.- ���@k�<��A�o��X1D�(U����
\h�< ꏔ�J@8��\/��٢Jf�<��3�J�9R���~Y��ȗd�<Q OT���"!�ފG�`�Y�(x�<�W%U�!mJ��O���,�C�\]�<Yf�2z�P��fM��)	|��K�p�<�'/96p6�p��U�Rd{ʒq�<�3�̋?D��l)��aV��l�<�EA�@��l���O�=�J�Z��^�<�$o��Ċ�e��Hr*�2�BW�<��EJ2=��yd�ˊWe,�xŭ�S�<IV�&�Ls��Ձ�ؐ0�
�N�<�V��(}���>hB�pE�CM�<i1
�[@6]Ar�\,��Y��d�<1�+J�:s&����1��1�Wv�<�%'Ht̂"�\.D8�:��o�<��i�)QQ�=B�e�$==xH�a��k�<��@�&Dupq�@K�g�,�%Ug�<�5	�\��ѷ�] n2�b�]a�<�+:^�:!�� �<��L����v�<���	�Z���t���}�p@Z��B�I3P�7i �D�f訤�0�"C�	�Z��(�Ux1($�Tm]W��B�Ɏ,r��h�		x�Ѓ�Z��B�	"��!�f�#<��y��lʹڬB�ɐ5���;WGP���9YA'HcHC�II�� �D	����@Ś&��B��p���K3��C��mPq�BT�B�IL����vK֣�=*W-E�WƘB�ɴn����P�դ�\2�݈d~B��d�t٢f	%9Z��� �BB��M��X�c���,�{�Ż2Z<B�I$4�^���kZ�!�
!2�D�{�4B�	�F}4�84![�ke�RF�GqB�	1Z� ��NV�M�)�r-=�B䉸��#�F;�	��FB+5M�C䉏gl^@�"#�<o`��ih�?�B�I�rF�([@inQ���US��B��^���c��{�~I#Q�*�B�I9`:T�㨍� ٙ��R2t:4B䉞N�, �w�� '^ ��nSB�)� j0�e+��-J!jD�=	���"O��(a�\�$֨��ǜ"&���2�"O�-ىj��5�&
 h_d1�"O���eM�(O����Ɩ,qRp��U"O�P�O�~������:W&l�s�"O�=��.�x��C�cݪX j0P"O"�b
�5����v�B"4̀2"O��yBM�~o.����&�X�U"O�Q�bM�-4�Ri��պ;���"O.93Ê�,T��Hp�)E��[�"O�{։G�n� d�Ȩ%��b�"O°��h�%؊�j��26>ͪ&"O�K���%�f�JR*	�~T��"O~}iV�
~���A��Ը�H��"O2�+떐A���j�6"ֶ�{�"O����F�j'�fjR:�K5"OV=!%�̰-�d�熑�d�\�A"OZ�
�i�r<qG%�6@�T�"O�����=	�1���p"�x�"Ǫ�HߜZ~t�aa������"O�xڲ�ڢ3��W��`���	��ybH	7x"̻��S*��(�t#�-�y�BSLe�;e�ׇ~r*|R����ybg��P�V)���K�T$�X��y�G P8�xɂ�P&-��aBCK���yҤ�l�P�B�S�5��eV��y�τl�
D��
�7K􌤃�U�y�gS��*$AV�H4s��p3kĩ�yb�('I�8O _�6��"\��yB�M'CH��&D�28���Q��yH�z��A�vE�t�`
�nD�yR�T(t�P��E�܉#K�(I1�ǹ�y�b�4o�(��ҥP*2��z���;�y��K�+�b�CD$�?,ܺ�`"����yB�	5�
�cVBߪC�<��OD��yb%��,�4���`���a�C$�yb�áx|T]z!�� Q�|��^��y�#ѲA�$}�1����P`
��<�y#F�YZ(e���G�\�f��%��=�y"�*Kz*���ȁM�A�4�W�y�],\���T�֔@D�4'��yO���,���?g��C�E��yrʖ�YcP�;�ռ
0tI�B�^�y�`��9-��s�FT8	+&9���@�y�+�<z��D�1�2N�.axa�A>�y҂�̪��@�E��y� �N;�y��[�Jo8������<���5�y�/M�꒕��E�Q��MPw���y���o��a���ZC�����T��y�����:U��lҿ:��cჩ�y"�U�6a�rF�A,^��S�Y�<aҁG�x�Ȝ�f֘{�����F�<u�ї^��R^�x���ס�@�<q�$C�j�d)�JZ3��ő�UT�<�s�� 1��$�ь,�81���D�<�U��+ �BE�g�B�.��b� �D�<����g=`(�k�>m�ejF�<�C�*e��`S���*�Z�j�M�<�C��>�E0��\T�
L�G�Au�<q$C�.L�H�Y�#	�.V���
Y�<�`J�*�qc�H#������TJ�<�&e�Bg�@#k�En���$��<I���)#�ڄ�P!�n�ѳ"����m�%�u�Bz
d�z$
��i~����S�? �Lr@�*q�:��"�݇K�(��"O��,=}슥�Ǌ�x�E�"O~����T�~sdA`��L�"���G"O^)Y��,����v�A�I��"P"Oh\�JߖS>,��Չ7��a`"O�H��L�7B`�2T��0� (z"OuI�m<L��a�+�
0�5"O���5�1�r�@�X�����W"O�a(��C7�����+s��)"Oe)߷"�0J��x�� "O�<��>a�쩑�C�p�A"Oĝ&�����(�"ɏ����E"O�1�b�,z����!���}o�i��S�R�s#�FbŞ%��jJ�?����ȓ\�eJ�1k]�t@"!+M��ȓA��4���lO@�!PC��uQ�X�ȓqo&��PM!���c��I�(��b�b5�%�,9�ڽj���_:���F�ZUJ�F�s��2�� N^Fц�P\�Ÿ�OLn�A*�L�J�	��al2MA�ѪJ���E�:`8긄ȓE�
�ig���ZE�'��9>n ��ȓZ)�i;'"�2��Z,қG$�l���%i'�����'A.A�Ve�ȓR�m{%�^K�Y ��+	��H�ȓw���:g���\�Wl_�M5��ȓU�,!��E�4�TH��b�f����ȓO:1�ǐDЍq2.�������{�������J\$�/��K�(U�ȓh����m�%:m�c
Z�]����=h�$��+aЁA��,vL���G�6Ĩ 'T+h.��9���1.�����l�3C��>;��(��k�"o;F<�ȓ0��A�k�}A�y�oD�vպ��ȓaI0(���N���sEL� D�(�ȓU߄P�@AG�m.,u+��?<ո���T��9��΁5����O˹��ȓW��X� ���B�
ֱNgH]��{�0�{�;]L.�A���7r�ń���C�c^L&�H8`��^�(ՆȓQ%�m�P���T�l��@��ȓs%X�@��,wZqQP�����ȓ}�������!���
"��;DNՅȓnN���s�Q�..�d�ܶ3�<��c�I��L�	!j ��'��8�ȓ-�}8��T��N\{��߀S*¹��h�����j�"7�#�M��dm���1� ET�T4�A#߯_QP\�ȓ a-��j�@��S�JP����ȓH�v]K��MBv�-B�
�${�ʓh�2Ǥ�3b��=��*�Hm�B�I9j��)P#J'R�6p�`�D�R2�B�I����e�*]�4�P��ū��B䉧3��Є�3Tf ����B~c�C�I 
��q����	���8�-�w��B�	��@�r.�'�����O�<��B�ɿwu�|:@mM�7����I�I�B�ɭo
�l����+��l���Ê��B�	?��(Å�٫b
��ht(C�3D�B�ɣ����-܅kZ� 6,B�-#�C䉒mA�t���R�#n6�&�2>�C䉪K2�L3�D+P7�91��<<C�I�S�J�9���/9I�9q��
D�C�I�t�v�1��+?B�)�_?_�B�)� ��i6B�aѰx��΄���"O��{� U�w���;ы����"O�d�Q[<I	���7�.yi%"O����G7: B�k���)d�6 �V��5LO���BA(ǔ!�c��"�!N�<FW�S�@�HQ�s���2��K�<1@��_�h �шQ�#�z����]K�<���	g4�P횠Z��e�S�G�<!b䊬j���"#�
�E��Xj�DMX�<A��FFB��m+�,"��	M�<�e^�R��]8VB%/=Rܩ���G�<1���;G�\�%�Z 3��u��
�C�<Y���.~!����#�N�")���C�<�$i�"NF��5)�u�V�B�<��N�h7>A��L������Pw�<��E���@`���75N�)���g�<�u���m3 =�`����ƄS��_�<Q�M� w.QH'�ΚA��sS��Z�<��-N	������9K���@NM_�<�D�:
ǆ����\0ZL��[�<QcE�!�~ᙔ���v*��6�PX�<i�o��O��R^�0�T�����\�<���+QE,���ꙋ\In<2�c�<�1#<�æjB$T�)�gu�<�WC��]wҁ(E���P�"�"ɝJ�<�ai/P�J�áiي_b���G�D�<a!/\&x��RN�Ȟ�P�
D�<��bA!_F3V��=�BЩ�U�<	2�B!żx�@3�n�f+�h�<�%�S�\��ya�T-S킥�
Le�<��	a n9�m�&[�̤�a�_�<�3��$/�|۷�S�o�C�p�<������5��*�^� A�^t�<�4EKIb��(rT�B�\�GB�q�<�V!�8 ]�%:S�B�*�pcg�j�<)�tڀ�R�݇<�D�Rulh�<����@��A7om�ɻF�W��yR��>Ŝ�b4�� GM"�A��O?�yrI^q]L��a�C�;�|�fS$�y����0/ȘiY�ʅ�$,�|LE��k���	2FR� H�@a&��8�� �daA�c 6v��r���4�Ňȓ�	{"EN��Hɟ>�p8��J������Ԍ|G(��%^�qPv���}���f�]-G:q�A:-s�!�� �8�r���4"hpH�f���`'������(�B�	�HigA/qk���ȓ��ȗ��('��Ǖ<�d̈́ȓ14�U�\Ze���V�����,+(����d���@���6�0��ȓ��@S�O�0Ѳ���&B��ȇ�/xD��w�S�b��h�"¤nN���oc,�0˜�iu��'�^EX��Jq|�P�H@�8N�	ԦC;`w��ȓ]$����Ļ9;
����
d��!��3-�P`� 1�h�e$�4L\�ȓu��3a/��$��j#�D!S�@Q�ȓ�L���7'�Ҍ"sQ�	]����?���� �P5@U$E����ȓ.�����Ys8��U䞋YAV(�ȓ^+�!���0UX������	����ȓmtX�s6i�T�8�j��H[Q0���Z6꩛���h�X���B��p��(Ò��Ś�"@����q����S�? �y�G.O�	bP8�4�גb���"O���D�&@� wm�)W�$"OQ;a���~�U��EZ;Exv��"Or�3 �Ty2�dƷLM��b�"Oh�kg��	4�"�
7� ����"O�]���ɺB�6��w �$t�� �yR����Pːe�����)�y2l~Nv�
�LN 1���$�܆�y��D8rh^���n(�vX Dn�<�yR@MP��G錡��m)"hۃ�yҁD 7�&�pdB'�<0
�dS��y⚞D�l�%զ$s�A	��L(�yR�ְ5~jL1ŀ�L��u��� �y���0o�QsG�]�GP|�)(\��y�/6vX �V�P&O����A��y�&��h&�D�!k�5�r���!�yB��Vv�R��A4�@��t���yr�Hu�H(1O�b��;�m���y�X�)ŪA��*ͽ|� �
�HE�yr!�gA��Ee�")I�E�u���y�n�Hxz����%,Kv-��b[*�y�i]����+��ڱj,�.�~9�ȓ&����1؜cĸ�DGY�fg�e��@�D�ʦR�r]���!� x����(_0�+���dN.��eI�_���ȓ���XB�P�Y�x��π�K�����]V�1Q�b1T��A3Ԅ� `E�Y�ȓ5~4�f�BȮ۶	P1;��8�ȓXN�X9a��F֍:b�
,Y󴉄�e����>�᳅	�+���ȓEvm��#ʄc�s��(cD���ȓ/rx@R�a�)$��l��E({-X|���ژ�b�=228�韭G�D���y"��.=��	s��'yȜ̆ȓ���y��]4"E��J�&��ed��ȓzO\���
	j�>eaG.��`o�8��Q�t݉�#f��i��]P�х�#|��d�!~����
�S\�ȓC��2g-��fJ^h�)�\�(ц�2%~���L��`$Z��@��谆�;���.F�0��;CY�#�]�ȓd�H�ö́O����υ�3[J܄ȓ@#���!�F� �g��0�V0�ȓ}�P��KT;!�TP��)2��u��\A���T&k��S�g	+>@�ȓ��`��(\̢��cF�U*B�ȓ����B�&-��# G^�wh��Z��c�@�\�
勂.F�
�fh�ȓAęH��Z9<�|D�6�" ����ȓ.v�a��'�2��"P��s6E�ȓ4P�����=�D�T�RK����� `b�=`���G�dzB剒N�#���d�n:0I�߬C�	~4��Ď�.h]0�i�ㆢe+�C䉌4�ؘ����h(�X�0A�g`C��2ަ �vFW�,ʈI��1g �C�IJ�ĸ���	2��x+�C�7%vB�I9J@ cK�,�Vm8v��&z�fB�ɡX\��"��*Q2���"�bB�	�2x5��-Y{�|��DN?o]|C�	�j�hR_�i[ʌ�$���Q�JC��Z>΀IC�.����N*�C�	}�̬�!(ÃJ��2E�2�B䉕0S�m@��!S=����$pr�B�)� ���@�V�aT�0�΋!E��]�4"O�M! ��i2��sŨ^>���"O(93���a)�a#�hϣ`� ]05"O8Mj���,k���E��X� D"O0�R��#:D�0ud�WD�da�"O&��'�͇%�)H��_()nj�"Ot�@�/�1�N8�!�79��7"O���C揖�,�Q�і	��@�"O�D2e��.f�1��;h��}�"O�X E�P����c���&��D�6"O@I���SK�>x���_=U��9�"O�e�Eh?2�k4����X�"O �����Ke��)be��
�"Ol�P��W�/�tM{�툑1�V��"O(hs��1q�q��kʊ|e"O�qhr�ϒQ�$��KX*�b=�"O�<�֣��$���iPL	�Z	�""O
��r�L���0�i�a
��r"Ol8Yd9J��`H��(��u"O��۔#Y.t�RȢ���-C8<yS"Oa��Y�N@P���"J�.T���"O�]��j��f�@��Sf8���"O���'`�p��q��+*�%"OdM���0/�Z2I�Gʼ��"O����Ȉ6�p,�&ޯ<�Xk�"O���՗;D��@s��9��Y�"O�	�Ȇ�6�`F�b��W"OHY�� �lΚԩ �\.:���H"OY��`ҿE=�-:%��-0�8�#"O2-�P9��MiGaώet���"ON
t��7Ut�"r P�?l���p"Ob�J6�U.d�Аsn�!0n�4"O�`(A�R���!��V�f!"Q�%"O"A˳�Փ�J<��l�'OT�s#"O���w
;"�=c-ɫ�����"O�@�,[| dB�U.P�� �"O]!t��B!�_x`�"j!�䍻#;��iB�/Sr S��.1e!�dT�AG�u`7l��-A�y��D�S!�$8d- `Ad�^�Pf���Ԋ4n!�D��m��b�K܈pS�<����}y!�d̀ ��d� � �S8F��i�&}c!򄚠A����ޞ�҇�!򤐫K�P��P$@�4:�'F�-!�d�Pa�Jc!������K(N�!�DW't���ic��k�9��ƌ�8�!�D��R��fLEX��ˑ�՘$+!���[�Ȥ�$�)�ȑ%�8z!���3�P+�c̸ ���A0���!�B"�Lh��.�;6� ��c�)s!�䟍+А����J�[�-h!�dʉ5����� �>��0�ԫ�9M!�$
�(�����h` �K[w.!��\��h��kɌz~؜�꒣9!!��X?]u`� �v��ДC�q�!�M$k��@��*�
�|)e���!�đ�|�����Z:(ǂ��(Ϯ[!�$:wC���A���T�;R�@L!�Ē�b2����B�4U�A�,�!��5l����w���M������@ws!�$Lz���䠉�_�P�@��eR!�Ĕ 72ne�6`ڏ2WX����)=!򄒗t��J���%7VeSצ�[V!�d֌m�"yv$A���`�RJ!�� �D2u`Z�<`LY���A]���'"O�|�r��*8��� OE-M4�}�V"O����L'�*�S�#�<d��q�"O�+ ��H��4�q�I1��`*E"O�h��ËNg��g�ѐ5��� "O�}��ٙC��)d�Y�]~���"O܀z!�Y.W�J�HvB[�c]��"O����煊'�4]�Ł�&ΘZ�"O��9GAц�b,z�@�!%�X�"O����BQ&&�|�q��fe�	ˀ"Oҕ�@ �T�; ǁrJb���"O��Æ� J؂���΍;�h�f"OU� �Ol�ը2�ށB5���"O���g��Zq�xȄeL.|N��aS"O��#Z^t�ā*_��!�"O��B����D�&�*r�$>rH�"O,-Z ��u�`��aV#x��"OJL�רO
R���B@I�@�\X��"O�H;E����b�Z��l#�"O�IsԀW�hO8SD-���P��"O9K���6Y�Qa!m�w��yX�"OvXZ����Br��;+�hH� "OX 02�N1A��fٖ( �zS"O
�s��C.#�ihu� %P�a�"O^�rGN1���Z���O�r�"O�թ҅R*G��Y#U�E���Ĺ"�!�$F�f���mw���w]�!��<�%ił�69��`ϨS�!�)Ffֽ1 �C�����3Kz!����yQcV��mC ��!�$�(6�>��0*Z�.�:Xb���yk!��(R�e)RN���Ô�� �!�dW1*2\ñ��4 @��w�]�O�!��T�N%���%�C�k���R(�&�!��I��(Pa��9�rYARfύAv!���5x �h��_!>׊�Q���-�!�,Z���M�$hְ|�"o��n�!�DLC��ʵ煠"��l�����!�D�F2T��!f�*ª�Y��җ7�!�$<��H����4�$I��M՘c.!��2�xuJJ9\�x��B�A8!�Z�M��آP@	)zq�@�U�R!�̌<��x���'(��C�ݑ~"!� �F7�"��? ����N!�$O
R�~�ؗ�OI�+v!�d�4-���sM@�DD�
E�M#�!�$�/���0"� <ڐ�pJ�;�!�X�kX�-�'!Z]d���C����!�$	��Y�i,���U��=�!��\�n�F�c�I^�On����h���!�$G����%�IQ�J�(�8�!��6:���7��/*�ł��J�%�!��^����Pb��&m���jZ�!��0{ƺ�@6N�Skt����ߒs�!�$ۆqZt`��a�%q�e��Ė1|!�ͼyZ��f eiD�2���vs!��O�>5��,�wI��""�;l!�D� <P���.��!V ε[�!��=%��e�ȗI��8���G�!�ŀ� �y�Lr��0��N�#Y!��/��,@��S4K���hU�>e=!�d��#��UQ fǎ>+�Z����!��(ȍ�3���S爊�c�!�N:�.�s��
[��`h���^�!�� �XK�Lާ[�,L���R�F�A"O|Y7Ϊuќ �eHZc�Z� 7"O�Y@5�;3�, ���(�Ѳc"Ol�b�Yc)셃s�q�lτq�<ٰ��.X~��y�ǂ�G��l3#��W�<pd˗6�fXU�\���Q�gJV�<��N
i��l:�"ƥ��T�*\O�<I`E�&hi�@��$A�F@���q�TO�<���I�	�e�",�U���Q�<����?�qR���uaAK�<��I�9-���W�� ��gG�<)d>t�ay�EZUph3C�m�<�ց΢ǦM� �*J���BSP�<9W��>8�0�E�����%�WJ�<���Ƽ!� �X�ݷI�`e
�)a�<���2k�傣gK�Nj�Y'At�<�%��62(3aK��$���eXe�<����@?�HR����?�>Љ��a�<��ם~/��r'!@(�%�f��]�<��L������)Q�f�##Vd�<���	��9(P�W�,��P mb�<���B+�Zk��R��"�:Ji�<I�\'�T��v�
l+6\��b�<��[v�	@�u�@m3�TZ�<!WZ6����⛀d��t����W�<����]�j�9���vhA@�l�g�<�����A2��ۣ�R#X� X@�f�<�ѡ�=S��Bg��{=�+UOd�<�`�'M���W+�>4n"Q#S	Pg�<�RN�yw �$
��*��g�H�<��ɬ�L�����0:.�Ae��E�<17�M?Yl��hA�1Qq�����L�<)3Ӑ��9��M��S`"��0��_�<�"�3GU�yG���0T@�,�Z�<��H	�<�")KB���m#��LS�<���);F40v�z���R���Z�<��mA8V����X8HD�IX�<y��'���[��܅*�"����j�<a�O�X�����
�*h���Éd�<�C��Z��t�B�J�T�*y���_�<!c��{�V!0u$ݔ`�����B�[�<��n�=\���/�Ő�a�Y�<�BK�J�&�#���	{nHݚG
V�<���:3'�j����u2U{��M�<qs�T����q��V0f���c�E�<�A��[�2×�ԐZC��r�&�B�<Y��2h�Ĳ�`�TPr0��d�<�#�*[�10Y$t�҅bA� b�<��N�`�u�Ɍ#	ԑ��\c�<1@J�d�20h�m�y�ѫ�g�C�<�h�8��kj�"lGa�$�:D���$��`]� ��	����#D�`�Ŭ:L� |ŭ��ͺ��#D���rDCaC�d�+g.��z#�%D�@rgR,OlrB�Lʬ�Y17D�<p�J�-�̩��T�7�����I3D�lp3��#��q��R9XX�)��E-D���f����uyQnO�ZD��p� !D�4���O3T
�͊ Ŏ$���r��>D�4afӸ9�V�:���1pT�$�>D�H3C���[9gh96T���=D�l*5��7>���j�iI�^�Fp8��8���<�Ol\�q�O8Z�������֥H
�'~# �<&��Z��?�F8���� ($j�׆i����&�G$	)0�"O6u�a/��Rz*08��;��,�P�D&�Ş=
l���4Ri~���Z 4�ȓ7��dqc��<$@@�	���<<�ȓ4�Ja(.gkj	HS�W�n����&�z Y�[�9� ж����9��X����T�/�r���[a��d�������Y�X�t��9�<q���))e�\;n"D�`3�
W2PC6L��I\�P§�%D�P����Z@��M�"����$D����l�?<�B�r�]�g3L�ⅆ?D�l�EQ�*�<2��� ^�=J�i=D�䉀N>=<,��tgW�²�-D��cՋ�-՚u�FD�!�DH���)D���g�_ W�d| �<��`i)D����7I-Z�x&�%Va��f�3D���դJh{����(7���s�3D���Hҙ4�d�lm���3�0D�(�
��pD���I�oK�"�B䉁�V`:���f�v8y�	�;^C�I*k�AVT%�|E���j���d=}b@߯,ZPD���U�I�'�-�y\:
V�h�D�I�2�a/�=�HO�=�O��fE�(|d�1���1�y���XHH`�#��9;��a@����Py��9b�Q�5"#HfA�ׇ�^�<�C΃�|��XG�X�F.\��gOP~��'xPىDkE<..J�	C��n`�	�'��4K�Ҹ{�\۳|���Q#�>���d4�\�
�����M�@(�숹m.�~�Y��C�@2�`A1AK �J��3m8D��C�b�*��\��J�/�L��';D��XpF�R�*�;��G{�J��g�9D�X��J��j�FF�8<Ԩa�6D��2�G�-���Į??*,��'B,�hO?��N�NL�0�C�4$"�x�w`%�!�H�y`<4F!u��8�w%�i��vÉA��<��ꁷ�dIB��9 G
[!�d	5_�n1	5�֗!'��0���L!�$ą0/��U��N~�T��1�!�$�� 6  0��r�]��"I�5�!���'�2��`j�؊�E�h�!�D�RmΙ�+�UB�� �!򄉕p��b�7��2� F?`�!��t�����C�	B�6��5)�.!�O^�=��T���(i�.��O˱b�D,qT"O� �Z�CՌ�Xe�bw��$"O�e���O���ꌥi�����-�y��A�>��mH��#a� T��nZXQ�<���i�I�U�)Vxj�; .�'/\�!�pm2D��M��E���cK��rUISBv�����j7x$S�#�*3�d���m�V�hG{J?���k�R�Z����s=�}�d�s���'?�Or�=��#�.�s�܀J�=��n����q.�A���1��3En_
�%�'�ў"}r��x�J,�&���I4��3f+�m��hO1���	BE�4b��	%e[�t�`uB�"O<���Hv(b3�m�td�Ӟ>Y����%�0H���j�6t�D~2��5e�8��ҌO�(�"iJٌ:uBB�	�'�&t�sB@RF�Z�#?ZlC�I�g������32������NC�ɟ%%�IZ'�/k�Es��͈^@�D/?�M<E�$�^8}֔�1O��v�H�e�}"!��  �ŤP��E[��ȻZ�: ۲^���	R�D�����z)�u�[�&��dE{J?��
�^�Y�.�n�`Z' |ӾB�	�;��Xs�G�j����ׄaC����'=�O�qO 8��\Z�
�R��* MN]Sfc-�S��y���dy��`פ3�B��D���IxX��p�	NR��%�&8H���	�ON��$WB}҄��1s��B�͜�b��/���䓋hOq��,�Æ	0\�:tA��^�[p����IW�O2�l���_%��Lwn�	��)D���m
�X��܃rc�;��!��,�6�S�'9�Ӥ��=2���Ɇ�%|8���
4�X�Ӭ�i>�H˗-À�
y�>!�l���S�W�	:�B$'���'^a��Z�]J4L�V�X�U�3�ԁ�HO��'����䣒^�<��EW�`#n�!�y����:îQ�Q�##�'����<�}���3ZS}kŌU�0��"�AZ�<!$�W� ��2���>!{��V�`�azbܑ ŨH�̘3���C!̍�Px�ik2M��@�$EA�w׊7��)�
�'��1z!��'�V�Y�[�=j�j
�'
$b@�zZ^(��i�
��	�'��.ͮ�L�xq
N�R8Y	�'LX��$&�]���Y�
��9����~��ʔIK֤̑lE��2��%��	xX�H�ud��Dx�Hy`Ø==��E2�?�O:�e�dLR"IS�V蒥�EaS���1�ȓ/�x�@ɕ�X���a����	H�'x� ���C��3�#
_�A��'Tl�� AE�1�S(�5T�<h�'�~�a�� �	=�.E�J�Hd� o�<eH�~����(L�X�Dؑ��L�Qў"~�I�R�l�@�b˫`��А�>I&��$�$�?�u���D1A���<����l�<�2�ןO��@��%Ў [8HSh�5s$�<�O�����I4Y�}ّ��v7UXх��z3
C�INҶ�ӖV#H45��^$9z�����<����N�E��S�,�6Ȅ �0>�f! }��A�7j\
�E�X���ضDRN�zO��S�3�	:Y�2�S�F,,U`p���Wn #>y��i7a2]��l
]��R�ku�!�Đ�*}��+_�(��XRը�# g����	��y�Y�$�Ӻ��"܈v�"ayd�W���A�W�<It��^�PtL	 W�Ti-�m~�r���=���"! u���U
0ې��4�
<��2���H�iC�X'�
z�Z9�=!	ۓ%����g�1�����F�[Q���J�'�H��!�o56���C?���(Oz��DC0m��pC��
�8�6ϟB�V�)�	���I<f�Vx���Q&[�RQ�[sP�����>�Ğ�m���r�L�r�&�"��ZX�<�c�(2�$�)��+]�VX�U��h�<��+��-���$��#t���r0�:T�����	�S<��@�9>���3D���D��-k�9��Ȑ�6�:b>D��q4�ȑwjJ�'ڒV� Y�r�6D��� ����ݠ���(�H x�`4D�P��&!D�ɪuc�1�$t;��0D�챵턬aD���' �vE �;c�/D��j�@��K��}s��T	�Ѣ!�:D�(�������a"-E�
��7=D����΋�Eq*4�U�E�?ߌ��S�9D��Q�m���`�eH*�$1��l8D��  ��� /"�48���ШU�����"O|MnϢV��4+�d��1�:��q"Odl�wMT#�i��9Y�ș�"OZ��O�WJ��E`Kp_Th�V"Ov
��Q�{��d`r�D���d["O�u�T�]�z:M���"C�D�"O� �O�]H�1+a���W��mA�"O�T�T���c�K�*�\9q��y�,�i�BᲦb�"���z���y�D��p��Z6ԯY�����5�y�&�JG�,�A
T�����%�y�R	6S�����K�V��7�R��y��ȵM��=��o�>C)j��q���yl^�O��d�'͆��2@��&��y҇�'�.q�ҫ�/z�*�Y���y�'ӄ��e�#_	����D�y���ֈ��G�'8\p1�o��y$��j�z�[u��+&�r��BE?�y�D�=�x�b�eY��r)�����y�k\�h�4q��H���ѠGd;�y��2vv9a"�";��"�!���yr(�eӎ�z��,2��2����y�y	n���(�(�@u�˗�y�B��0�#%�7M��{D���y��:R8��b <F�*D`s�[��y�Ҡ����֫��C���"�J3�y����e<~�ZG�W�0��`b�P��y�N�w��iu-��>)ִ[���y��� uP��0�R�3�� ��,Λ�ybc�P��&K�$�����ѓ�y�� ȚL�fR�n�&@qڏ�ymA�^h�͓�E�u��y��Й�y�M��q�Ȕ��b:]hְ�`#	��yR���+ج��@�ՙ@5h`��yBA2r���􌛽w͘D�O��yҫH}����q��aA+�Y�����n3L��h'@��0=q�����TȀ3\ldE�dN�l�<�6j �Dz=˕��6R�$��!��k�<��
-]���fN�"��5��B�a�<i�d�L~|�12�S ���C�MG�<�"�H���@Ƃ�K�0!�#@�<�B�قz�!b�K5@|�Q}�<	����t�ҍ�Q�T?��t�T��A�<!���9)]^Xf���FElJ'
�J�<�uN�{@����-�����D�<qӠ�|�K�5����?�B�	�Y� �R��صU�9�L3)�C�I7$D[E��n�Y�κx�xC�Ie	\��iM�#^��t�X B�ɯz�zȣ �É,!R�2�� RN�C�	�%������X�><�5�J�i>@B�ɟn��KP�Ѯr�|xr�BWq&B�=�@���Xi�� �a��!�d�G�x���k��E�O�$�!��� r.l�v�'҈0#dΥ'�!�$W��F�bS�2T�ڨ�����!��	""�l�1�ͰY��P����1PT�z",�51V�y f\�<��],hD�ԃ�e۰E���Y�*D��b��-t/�uS�B�_�fq'e:�I�^�lYwŚ*'�Q?a�F#]�P���Y�Y5|ႰG9D�,#T�^��lƖg�ţE.�A�2��E��<q4/�8����BW���1���Lp���!�uD
C㉲|_���e�
�$���M�9'�h�e	-/Z�����Ro�p����+�	3�ǒ�@$Nt�R�4<O�'G��F(V\��t�� V��`M/�pa��HN����"O�x���=�d�C���O�\k�|b�J�B8�bH�S?�!`O3<Y>����̎ B=���!D���c MNZ��2)K�wEڷ�]�9�x)��<aD�_����	)'3ȸ��%�v.�ps����*�C�k_t����� ,H���QdAt��̒�E�*$��D�H��K��0@�UK�G5y��]��b6<O]cr-��z��E��Bv����\�^����Ũ@�$�$��+D�p7��8�p��f$CV����:�	W��� QA&p�Q?��k/P�� ��0����8D�\[6 Á>��!
���2
�܉��@�d4�K>�� �gy�.H�3�2|i�'p��-+2��:�y/�6�vAY¯I��8C����y���K��(8�k^�V&�3�Z5�yRgÊjFv��Q�	&_f�I�mJ��y2�G*=7D!0b��!*��ʅ�yR���{&��"�+N�!�L��o�&�yb':)�ԥJ��ɍ2���<�y����2�p��E�2�h��gW#�yRe�<>o �0�$��q ԁ�)Ǵ�yc�/ s����j7k=�Uz%Ǖ/�yR����3��l���T�M$�y�Ѕ8ߺy��i�e5�j�#�yB���fP�á�*���@��y���IQ�R��!��5)����y�oԺf?��I�*ٛ!�d�{6����y�J�@���k�g &�$j0���y⡝+!�z�l\�W�4�x0�#�y�#�%{5TL)���,8����)+�y�i[�X>`�1���2j�8T�vǕ3�yҌ��L�� $M�0S8�R��0�y��B�E�Hٗ��
q��1�b+�0�*�PL>�Bk����B����/��,�l�;�F�}a�B�I�B8���m�9p)�� �)�]�y���,�,���''*�Z��!T�Q�G�{	j��	Ǔ`�ZUS4E�`z�-��O��:��A�>�p`
mQ�`�j0:��)ECz����>6,�u4������D-<f��'X�3!/*_r�����ӂ��$��ٰC��m���ci�(�@��{��+T�>E��'?V����Y6��ǀK�w lͻ3�T���/��)��o/�3��K�>�:B��Y�T���WYQr���!Q��ͅ�q�x�3�P�y�o�*JU�U+�O��6�Ma��� ���t�kF�����*i0�h�C�9���`�ÿJ��a-ٳ=ax�&Ɗ}�e"DO�	j���"%J�"Sg��?
��%J�bM6c����@��I�$�h5KL8�񟬙u�Hn����c�)�����>�W;Y>`9q˓4��>Q.@y�+s>i@@@D?Xdb�{�A��-RV�zeEӇV����=4|���WT<�|�'��󁓂+����ѝ�b�Dٽ2:˓Gu@0����e��x��?if�W���R,Ovxi˗�ВrR�U`(� n&���4y�a� �ax"�V�\����V0lP�F�4$M-��K� *��p%��>h�MK�P2^��3¢_W3fL�&�7"B���]L��(!�����ڮ>E����|2�,&ƾ���Q�6�<�*�,8�t�R�Σv`}KCl�6�³쇨���&42�" yP
�r�+��tb�	��H5��-l���L	�x�n�(��'rvE�E���&����1�ݗ�.ɠ�'� ���ܳdDB�c�nPZr*py@���Ea�)Sf�'� ј�������dX"{��
W@Y/U��sa�޺/�ɲ_�r�f�[�pF0+��SU� �%J���'b�x�fo*zs8hb��@1gC�P v.�l�D�����2� k&�'�4ɇ$�"q�P��ԣ.ڀ8��ˑzDj r���|�Xꂭ���Sk�ҝ
4�Z�8\A�ώ��v%�2�]�=�nX+FM\&�輄��48)n`zeGW�r6��H�5]&p���P~`eP7!�,D�@l��ֳv��hEW�v*�R�'��ŀ��F)�uGE�v���O6\�ƙAUAF��O�hB♄8�h�z�敄;�`!1)��v�ta"�	�H%C��-J��(Gk�c'�Б�r?��G�X�:�|�'�8�5ٷ9f���D͐�I��Z-O�Yw�6E 25ã�� �lev-su$A#L|"����t��+�̙V�Ɲ�B��<X���; hʈI,�I�����V�d�}+3�~�V���D�fm!�61�Ĉ�K�*^Eʓ�ʐ�G��*_F�����%�c'J��`q�û.P���D�$��i��_�kE����*P��{CKĚ3W�dL
8��*��=5�B�*�B����π b�hG^�"�й'�-uZ�0��ɜ{�J����_�n��m�7���Y-��aЮ� u0~ŐӢA�an�I�������O�@8�B�5L���	�bd�\�'IN�`!FK$9���OQ>�XuI�2J��Y�ү]		3�M8��2D�0�Q��s:�%�p��i��hP)O���T�dY��_�3�I�.˾����u�sbI�6I���dI�-êٺ��>e��,H�e���f�t��@�?�?��16�v���!�_h��Bl@�'��P�Q"7BLx%>��M��y
����F�,�¥�D*D���"M�x�:Er'�D&-���vh%?��ΚN_�%
M>E��-K1@fh�. &
�z4"���y��1'#\�@��(K��r}�=�2@΋P����$4T��I�dDr� ��L�?j9!�$@��L��oT6-�|�5�τ(!�01��b��}�D��aM�=!��&�b ���Զ��/E�^!�$S�`�
$+�-�b�T�B�٣z�!�$ �C���"��{!T�{r��L�!�Dԁ VL���.ʥ&�������!����l�l���`P/�r��G�Y!��'2���v�;[��0�'��0!�d�U?�,t��?q  I���A�!��IT����+pC�igeF��!�13�\�sC�{�d�0qx!�D1(H�b� x�(�rS��i!�$�&P����T��E3`���!�Ā�wS$4C�ɞC�`�
� $B�!�D�@l��P���3�P	�D��[�!�<D���j�Nӧ+���[&N�S(!�$@6#XnX��i��X�ؠ��� S�ɧP�f�r��'q`�����F�D����7=^�0�{r�.�`����-�n��#�֧�ܵ��*D�F�bT�Y1B���lڻ�V���'꜄IGȪfeR���H-��dR�n	6u���O���]3n�IŬ
w�]k�eѐ�~�� /]�~�:T�БFW~y�f�W1��x�+S<Kj:@q���-}���cL�'"6٣�FB�Qp���ǋ<?�zCB�Hm4\I�V�,|�'z��X��	5'�R�N�q��Y��,%<O br�Ϩt��y��le��BJ���6���I�b�r5�&��(q��p�A��W!�\�nףkz�S�(Or��6�F��~���D<4�6{��|���=1�.!qgƼl!l�'ym\EB�O��U I�}��� %�/=���Ñ�R����@I��p>ac�@��� �3k�%F��1�ő1�;A�O�>��Ir���B01�+�O�(�c���#I��!1��ҼCC��!K� 9��� \搉�o�Hh<�E+���0 �C� �Q�����O� ]��9�̓!;��8����h8�ek�� �(0���R��ᡱ��s�& ks��;GZ�=،L��ȉ�>�R��DZ�>Иd�uH��8�\��FG߽l��b$�Q(3#�aa7�ː_�V�fh@�D2�
C"��t���emT<n��j�I�e-L�Y���	Ԝ1EJT�?j.�O�%��<`698v"� �� �yݕU@�I��0�mу=�ȴ��%�^�H�9
eK��ϸ1*B�J2�'�r�cV� �/��8��*��%�z�aȗ=`y����0���J��4�v�sv�`��J��^*f�����'m�]r�o��X�4]S�σ0zv*S�,D��ŏ03��}�W�15*���mS��L^}��Y��	a}����<�'ƍ�#��|���ιP����   ���ܫ�&�P��d���<Io��R��2�֛1�����`��v���5~x�)+�<����"��бM~�OL�XЊ��C��4��N��R0���I�Ez��`;
�ЅY��=��U�&�ZI&H��UIXГpHC�`$l Q�)ԓb���b��%�O��iE�K+(���T�N,�:��ܜW6���bL������O�S�}@*���kF�.�D!̓8�u˕�gA�jũ r����x�<��䖽,a,�Rf�Ϭ)�����Ct≟YR�ѳ���#n��Ȣ/Ob]��O߬���	2DI��dL	V�[�aڤT���2EK�) �֩B,����[9�pe�&"[ Sp�
�R������iq���D����r�,�g'�e6��Ɠ� U�V��7 uN�X���%��!"��4i� a;0������#_ǐ�pէ	1�T9��Z� �az�Äh�����@?iI�F4����=0%�fO�I�<�/�2l����e�d� �G�n�xP����ȟxDiC��	F��*�bC�ED 	""O� ��`��YDV0�E ��}���ز"O*�"��!Pt����H/��8��"OP�Aȏg�x���螌��"O��`�/X,j��VJѹ���B"O�t3kÓ7�vك�g��Ji�� �*O�}A�#����&"_��k�'Ҙ��mV�jJ�1�/D/�Ԡ��'�1��� C��=	v�y���	�'+^����L&�!��-A
'�:���'�
iB��8��|�C�����
�'LH����G&@�BdN]�4��'	
�D��\_ԩ��(�( r�@��'�Z���ꉼ�h�ZңC1}>��
�'�`��c�S� Ii��U�jl"�	�'u�]!�I�2}v�[Q��Xc��;	�'��p4�3�<𚁩���8���'N�  hά1d)��t�bA��'���b��R�/��q9�
�x7�i��' ���!˜ 7[�(0�J2Vؓ�'v6��.ռbh: !��C�z#|���'dj����6?��=2���O���;�'{F�S�
��Z�8<�q�-���'���FL�E7��ْ�]��t�C�'#��%e�!~lT��"��#{`>Y�'��}J�o�	0�ALނa��A
�'ㆸP�W9%#0�ۑb��^����	�'�bq�"�V
^EF�� ��?H	"���'όe)sK�2 ������@���'�8��ꚥt�����ͧ�4���'�H��0n��<�c��0E�x��'=��2�6 v��R�!8��'���Q�7x�IR��(  Ā��'�h����5g���aM�!sl��'���T�� ~��p��A�z���'|:��E ������:@����'֞��& 6����'���0��'�`��fʸnW��f�V8@���'� ����^.܄u��dC�csZ9�'m"����HA�!�7�ҕY.���'�p���&D�͐���1C�v�)�'���G̟	�ZU�E�?��\@�'�d����E�ܨb@ �:^�
��'^��a��6;Ɓ����c5��c�'����V(P	�¤��(�0B�9��'!a����d���@��FdA�
�' p��OY�;h��c�E�)��Z
�'d�1�s&���~���)C0=�&a��'^�E����Z���b��	??�q�'��A��;��A5A&�4��'�>�ˇ��(����Ć��A�$y��'�V��b�ڈqm+YV����'-�U���e��!�G�R�h%��':�*�\. �d��K�@��'��2$�|(tX����%:Ю���'�B��@��P4(l�V��X8F���' ����\F`L�2K]	D*`"�';D�u��9uP��"R�F�CJ��
�'GL�Y��Z x4u�!�
�4`��'�2B�ڪ9CJu"�˜�VH���'����ak��n��T�ءT@��"�'�J�ᰬ�� ("\�5��J[���UrEy��R����X�t!8u�BŒ+�v����/�!�~��A�@�B|4Y��r�1O~<y�FR�p� 8و�IG�# �0J�B֊�M	���`�!�� �I��Q�<`�o�pkJd�6Ꟙs���Y U��9��i�g��8�D�#U	�i��#ƀ���D݉9��
�L8t`~�4O�;h4�X�ڪu�p�sG�7�O�ѧ�(' l���ݻ�v�`��'%*p�Lܸ�b�H�8O���3A�)(l#��_$V���j1"Or��EAD� �VI���<��PG�|��ޑ9���(�`ƩZ?5ڐ�Վ0�"���� ސM�2'>D�xbE�<$�r6g\�+��1�$P8��{bl�<qևF�����6J"���$�>|9����3Jo"C�ɤ)����Ն�Z���v*O'�����	\g|h��%�_�LY�E��������$+�D-<O�� �(��<�dm�<�!��1ttYz� H�f�pb&D�(V�	�utD=3ҡ�ǪT�BM$�I�à@�Z��	�����J�J���H�&N�D�S0E؇`w!�$_�3����RK�]�쩱��o��(+[H�I�nQ>�f���cшT�:v�m��D��s!
��u��$����
Qj�c�G]�����p�Z [�(Ƙ,������}R,��ȓ,̮�*W�Q�eJ"�/��]��YT�<����4ۜ�����/ <���T�<Ar��9�h���Y�9nT<:SdJ�<��NêQ
��D���9�BEK�<)�ŕ�m��]h���6�
��'�S�<�Vl�(H���ڡ��n�xI�-UK�<�E�Lj� ��C�z�n82�a�A�<��T��|�w
L-M6f(9U�A�<9�$�r�`x��@Ţrhx��"��<�SLޙxf:1��G�E�r���\w�<y��~9(��`� �Y�h��n�<����Q��ds��7W����)Yo�<�U I�zU�Y:@
"�&`P ��C�<��E#^`u�2��'��̫��`�<I���+S󜹡��@s���fA�^�<���ͻI��P��;\�ń�Z�<�Q\ьD!fG�_-8�Z�NT�<A5!	�qYr���E�J��ёsJU�'�ԁS
�W�g�.^`���A�Ԉ9�Ԙb�ʓO!񤗘v��-;�B�X��isP'�8!�Ig��3(���7�~�S�M�;�D��q��(K�<��	)6D�+uB ٦(�'�6x��iE�4��E]�f2���'^8������)��w��XQO� �3*�*䶍��N�G�OK�\S�bӂ�	w��k1�u��'�`�C JMm�����J��	�f}X�W�����(��5�<�3�2GPT��]�^ɀ��)ۡ�D٢+A�����'b�<���#z��`ڵdʼ,!�PAr*�O,$[�L�<�j��`nF�n�ܬ*��'l���ŧ��ɮ�[�Z���g��}����{���W-�:�y�O�|�s3��%P1p����,��	�I�r���]HX�%?�X�XO��D6�0�撼5���xӌ�F!�$�!��0yT��Q����rJ�<f,"0�KSy�K��z����4� ����'���	�wG*�y�Əc�����ܡ��T{�'b��贅қ+��D��`�\V�1B�ˋNX,���K��8�0�E� �#�����%�)��@���d�m��urtF��RC�	�#䏾*�yb�SA��3�����Pv��|J�G��4p���Ί\�qP��M�qph���Ǚ��Dr�W�^�>���
��y�]2�p<��/��*�`D�F�	�p�n@��KW"	c�ԊqbF�r �L��U�9�PF�-��?���� G�V�{ �D)B�Rvb�I~� ���^�J�E���4ID(�(u����h%񩑸%'[��/#��5���8!�d�&����҆�-�8e"[�/�޹1�jJ�*a��J�O�U&�!�"���"N�P!�)�'�F�	7�b �h��U��~�K��E�J�YG�E(.�pL-��J�.ɣ2kN�������B@��B��$�i&�Ⱥ5��m#��sD�K��FK�?,��PvN�?+"�[R�
(�l�8'D�K4����#���aO�vE�e��	0:d"���g�-c���cR<1m�˓��U�c�	�L�Д)WL����	Ћٵ9��� �10H�-A��y��D�-�pq�r"O�8*��=ǔ�R#��O��4*OH�q�>���	-0F�$k���O7H�t+L`}��Q�w�t�OE�X���Iݣ��?i� Q�r�Ȱ��X?"���j�!�S�p���/���3�^,T���, h�џ(@D]9SX�RJA�*yNE�w�$�t�BI	��˫��1�^�AN޿j��` �O�
s�T|�bE�����'mJ��b�7�������0r�DmH+O|�"��ڠU�ơM��|*��۷G��J֮τW �@����T�<�0FU%v�6��BM
�@�J �rja���� �eU���g�VŮ��C�|
�) ���,Zq:����+Tþ��c��:�z��"�M�h|Xr���;�A��'nD�9��pK2}{�H��(����� t:�1�Mٿ�ħ㎅!Wn�1�>l����[����C�*$����9g��#�\:Z��'��+ЯF?�ɧ��i f_�(���a��\%@��� "O�@��E:;�@1�dԬ�
�yQ�DV�@��i:��ч�S:$�H���`�%�4��ȓ�R�I0`�8|#~���̓�h��,���e��7\����X�l�ȓ:~���T ŜZ���`��tG�T��'����q��C�(ڀF�\��|8bdpV�c�܅�P ��P��[���8��P�-��ݰ�@�*Q.�ȓ-�lҧ���D Q��á5�����)&J[� ����dʴ�Vt�ȓ#����g�N�z����[�~�х�/�~�㏟"`����
7�z���P![�
���M3���M\���5��Q�q�U-�
LC$Ň�f��CR�B7w�B���m�:3���0��-��^������� B�ȓm�tH%��  �����<s�"����V�u���B��P�WcZ'O���ȓd���h$�5n���	�z�1�'��|�1n\؞t@`c����)�R��U��݂��9��*W�j����CB̧V�f��,��kd� WbU���qLְi����u�i�N䒃J�Vx�D��#�O5T��fO�o��@$�L8()�D�>9�AH�K�tXB��ƪ3��Y���Ԁ"�p�;.^����E'C�T�Y�C�U����Q*���W����V��u-�Qc�%R �iehH9jT�`���6��M�"�T����N?i�$*�;@���*�7�R�HgB*Mk�y��L6�F��B�+Oi��/���n�*�2�BED���UL(�ح�r���$SN�`��_b��ɖg,^��W@�1l��&���xB�O�+�"��~NEA���H�� ���ɋ��]�w��5d������=%'<���oږ}kz@+a�'*�����L., 2-�c�#�W�Y� ���"bS09C��Q�@8��^ZDpb���N��)�?�"����P� ��B�%�1|���O��9��_")���sI� 9+�]���Ja��5��I�>�l��BاHd��)vI^!%����ơ;.�Mꄶ�U���H���E�A.�(qx�)��<	'A+�<Y���W�"m����h�����/~н"#LH�Je����-֫9��ẁ�]�2��,�����j�FyBĐ'9���G̟���r���������GKQ�3��<_t��iYw��Li��B��0Q+ט1�-�4.{�-���S��~�!���L��|��ևa�b��Ԉ�9J��k��<�dUx��+N�0����w�����V�`�`�#��3r��U��o�� A*��e� )PL������1D�H�bǝ) �p+�H-Q{f��れ�(tة����h�Z%W�;,�P�b��<����_b�0�O���J�@׊IXP�T��R����H����!�z���* /��#���[�"��Qa�����z�(�x2-~M�J܀���È��g���n�3�� w
M�3�?����G�ڂ~92�0�N P꒟:�@�$��x��Ј�	��59���"[�Azy�7�������40=�eY�˗3{����D�!�:H�ؖ��`��N�\��T?�낥͝?�hS���<����K>~��c�Ӯ���Q�k�<!sh�S� �pLإa�n��`3�Ę0K���E��%Nc��'�&K$�&��DƏc�yx@��wMhX��兴��?dNF�bh;C^�nƴ�Ƌ�a�����6,�u�.OR���΀����I(z���q`_Wl�B֣�j<�B�	�>��rF\�eV�se�L�=����(S�-`ʹk6Eq�� H�#OL(�q�b���?�N���'��Y�l#�}��p�|�c�iσgZ41��&Ch����G��(���R42tM��c5#���=�˚�Er1z��IEA8N�:�ᕡV=�p�	�P�!�C5��I �B�s��0��2�!�;B Ƹ	�� �?Ш��}q�'�HJ֏�e7j�s�lB4s����'f�|��!�Q��1A�a�u�
	�'��y�b,�h�M� |��r	�'� ���s����g��&����'Z`Rv P�[����S@��0�	�'��H���8�����^,E�l���'�(�+W x��#K�8V�x	�'>��Re ΰ �Ȉ�$3 8��'?��(��*x�HU����8��<��'�4!�!�/U'�%P`KnTI�'^J�"��=e��WԎ3|
D/D���Uh��B����Y66x䩐Ǧ-D�,���S�VЁ��f��e���C6D���LT�dh��G�M��	�a4D����P�%;5!f���m,�Ჳ�)D�X`RG�),��[�ĕ�v��M���'D���e�֏NKV���l] <܍�$-9D���v�ԯI�<�A��JLX�ro6D�$�D*�E�R�y�]����i4D�j���H��T�_��H����4D�����
j4��j"�N6m�>���5D�`4��wvrx C
$֥��7D���AE�
P$\� HG2}��$��2D�L�w��w���p�B"�~ɱ�i3D�,IA؏$�&��Pl�2*ULi�W/D�P�#�RF6(fa�'
(� ��*D�ĺVIZE8�ǉ
[Τia�(D�D2f�L�V�0`��I�����'D��P��a�� C��ؘ�2$�$D��1���/YP�����5A�HPbK&D�|+R��{,�I8�w�d�pa9D�p8���7;����E���%z@�6D�@����	X�m�p	^�H�d�X�4D��@LG�F\C��?2j(��!3D�8���Q44��X��UOFI�g�0D���c�˟D"�����9.�H�� +D�4ҥF�,��!�GIĐp���55D�d�1!P
4nΐ�e��V��pE΅�0&�
[h����>���ę0hV�JK>�;����,��<�|kF�  Apy��������	�+*έ��SCb��6��*gc����}��X���)!0�禁0��кV�~���"({6�R*i���	�<�wC�
���~�RH�DF0e�z�#�CX@P��f��7}"��P&2��=%>���?�r`+5/É(q�4��,=�DP�a�{���'ɂ��g
� ST�3a�1������'Ȁ#}�͙�)�P0:1BA�%���1�1ݞݑ�
ç p`��`E�(�����V@�y��WC����IH���G��t�R�F�ĭ�'�Z9��T?m%��:�k�d	�s#H�O���o�|�Gz����iH&`*����5z��d�H�RV�'{�	��0|:� �k%���e�W���f��|y��)ʧV'���aA�:D�]y'�ޣh!f��ȓ/>�)�� �I��A�`!��MF,�ȓW������ޝ_��e�W:�6��'ў"|24�Ҹ��A$���X����<I����M����3G���ǭ5}2��Z��OƸ�5*�E*���IV61���e̛^�hY�}���i���A %\����.p���.KN��I���)��0�dZU?>A*W�D<Eb���$"�S�� <įF7��=�7?��QӘ|"�)�X�~���eNĄP�6H��[� ���'#$�&�����i�?i�bn<.��g�I(���jΦȸ'Jmh%�Ok$�2"^�?�`|J���xl�O>A�#F.�z��>����\ `+6��G�؀1&�Q�<!�[�}�ڙ�cgD�Y* ���ʙq�<�4�� "Ȝ`��e����	Mb�<�աB7 ���e�,�t�a�<)�S��VQ�LJ=��t[�'�^�<��l�!�f=���ߵ,x����t�<�dK �S}D�A'���.ڴlP&$t�<��W�4�>�6�
7Y�^|�	F�<)�� 4r�B���mŴ{�����|�<Q �Rv��ԏQ3q�Pi6	��<	&ȭ)>��Z��[�fe����J|�<���	,���iզ%*`�@b��s�<��(��6B����*�z� ,�J�<����E_����F�	^UrԧSE�<a� ��:�d�Z�̎�i���
QX�<�����H8,	�Gr02�� El�<IT$�'UQ�u�A�ڽ��a��g�<�DG�v�2�;%H�iEȽ�W��d�<�s�c�X���ț8F�j�,�T�<y�lz� y��R^��q�f�<!&JT���[�B܄�n�`�<Y�
_-&c���oåq��D`�\�<�vG� U�R�jr ��C:6`�f��b�<)s��\/^����B�J����r�<�B�����WR�ĪD�4T��P��o�*�.��9�`A3D�3�!v���L�C�p%1`,,D��˧c�*(_*ٙr�\7eT2E2�j)D�P��KM; cl�jd�ܘk@��o)D��3R�F3%\��[�!n��&D��s�sv��V`̶}�mr��&D��$cY�h�b���o�2����%D�̉uiÅY!�APt�]�?��ri>D�`�҂�.�M��N@
a�� �t�8D���b�ͫU{Ray@�'_De F@8D���KϦv4>���L�:z�����4D�x`��b��Y�Y�|02�3D�Je��$+��H��V >�rp���1D�����t] ���V�F�xp��$D����NIi.|�H#���ah�� D��T�S4��1�$L�Sw�=D���ǡ_�t1����a�gb���.D��TM��hP� �$���d?D��ण��g��" P�H	�]С0D��zv��j��{ �"O�"D��C.D��Q�*\&;�`��OL�W%<���-D��2�jV5J�<9:��^��4g�,D�8b��*,<�ቧ/�roP�·f)D�4���ͺ"6X!B�L��B����+D������K����c�.+����%D�`{�%4.�X��jS�idP)R�%D�p �N7d�0.�*�~��b0D�ة�Η8�ab5�dV�-��B�ɬDaTY����t+�8�0���}��B�	�t:�I�AS�iQ�,b�HD8_��B�I�U��B��3���a��#tB�	7H��u� �Z�9���@Z'_8�C��,�:!�ɯnS$pR�@C�++�B��-F����JF��i��J�	��C�?f��8@&u��6��Li�B�)� 6љ%*�E�"5�7��\䔝�S"O��Ȗ�]�
P���P�}��բ"O~��Q�D-m���Ɛ��8a�"O$�y's2���aQ9=�Z02$"OZp�#�L'6��jsAN%c4}�"O�!�R�ݤh�Ax�@N�-��@�"O��
�͑�4ج����b��yV"O���NK�.�!� E,���w"O:��w�-���[��	G^5y�"Ox#%U:b��a��4w���"O�l�VȈ�n=����
^0δ��*O:}��@�c&��p�B!|p�b�'�N(�Jγ&����mxp�h�'~F��T���}�ܥ+��D�$\�B��;^�軖F�1`�9��f��0H^B�?.
�{Pb��!3`�[��\vC�0y�h�C�',���, �.B�	�ku�]��L�*)v�;��D	3P�B�	�w���j���S&U��a iԪC�IK�l�	�DI4v�&EJE�Y�c��C�ɢ7�V�!H�\� �3�؂U�C�	�<,�a��kU�,
�dh�'�G�B�	��ܻ1�I�V��j���>�"C�	-�P1P3=uu MI�n���:B�ɳk~������75�2I��RZ:B�	-a
jA;�)A��`�݃l�B��,���f�X}�NMA�� �B�	�8�#܏�
Uz!�ſ%��B�ɦYhY��'��=Zy��eޢ1��C�	�g���0�%|�M"��)e:^C�]䞜�e�3PB(�b#��2@C�/N�����o�֤�UJ�+ �C���mЦ�
�#$�|u���C�ɵW�dH�U�0e*������4��B�en���E�̜"���D�C�	�'�L����X|����8o��B�I3C1a+��:K0����J�$d�B�	'�.9C�	�C�����'\6'��B�ɶ/3�Tx��" �J�c�f��})RB�I&]萴X�f��*37���<D���ă�^��c4/JX�PA0D�4h�)�;�Ժ%.�,!�jS��-D�c���]�~-�E�Y5(� �'D�Dه�H�o����sŇpC\���#D�(�+^�T��|;6A��_;�]�V�6D����K�T��*��%*ֹӡ3D���d@�4W6 �Acém��us�3D�Ⱥ1-91�@�8��4���x��/D��s���:$����T��?��(�
!D�С��M\�� h�/,�q�Eb>D�(�W��'1�*mb�*>!ò�	�=D� �Ϙ�tV�e�v�E�3-���<D����].�0�!�NNru+tk;D���&�!BƞaKUm !&9 7h%D��5-�Z���F�,:���&'D���F�����)% 6��l2e�%D�DX�ԱWpp��7)�2Q��J	#D���W�K:�T����γ|�$��$� D��R�M���[î���W�)D�`�#�L!_\��P�˅v;��)(D�4���8sE�)ؐjD�wL�ya�'D��R-S��Y0��-[A.���N'D��Y%%�#2P��e"G":�D@�f�(D�T�v��>yʥ�ŮϜp��I�G�'D�� * ��H,=mz�(��1+T��C"O���5L��.��aPb��
�M`�"O|��@T�N/ƙ��O�&/˖0��"OB9r�H8�J�SF�;� ��"O��Ht�$~h�g������"O��I#`>Z5�Y���	Y�����"O�,���Q+5��b���$��|��"O���#X�f�H�9�!��b|t2"O�0�� P�.�p��@_� ��S"O�TÁ��(M:�P�	S�M&.\1Q"O��Хa��tD<��Th]3�T�:A"O��B$�Bt�)b�N9V�˴"Op2O�&�`�
g� ��Jb"O,E�4�U����^##�"Yc�"O��p�g3R�i�n�|눁Z�"O4]z�8P�d=�j�}6�l��"O������p�ܵؗ�C�b%`F"O����.0���G�($ !�"O�HqcƳT��<[4l�S&΅��"O��XȞ(yt�#U��/	<K�"O���3ڑbꮸ�1�H�B���r"O�	���	[�x��]f���U"O@�xenmx$�%w��I[�"O ��W��l"��IG��?� �� "O�I���a ����"O���P1<H~��OB%/����"O�d �ȼC&4��C��	���k�"O�qH6�]��S&Ic}.���"ONɺ��Y2Y�9�`ɰTc��Kd"O�xi��ʖi�� �-�i�:}��"O,��w&�/�L��f&�.s��]��"O^D�BfP�vU�52�#LK���q�"OH���m6���Fcۀb���)"O�X3�o�,̔H!��[�x��'�dD� G��]e����κzQt���'�~�2�*$�ʴs�D�m��h��'�=��fZ&dV�b�C֫k�Pܑ�'�a�,�d� ,R��H�qER��'�0�Y�aL�C��m���i&�Љ�'ET��ddצ��r$ȃ=c�xl�
�'��1"G�؉+��Hd�]-]f�1�'�,�(B��e����d!�|t��'n ����_���J�Ad`XY�'�r���@���
�&.��5��'�qР��*=B�s��4(�8�1�'k:Y��/<�PÈ��n���'���`�G@�|��Wg�w����'��,���*<L�������}9�� 	�'1������*�z�,�9"�t���'��3���AҦˉ�v-(�'�6,����x�6,�v$2�0�k�'�&U�5�/#�6=C�e,\5��'߄]Iř;&�^E�֧�%$��A	�'��q;�Ɍ&�
vn�5
¡��'v��Ӏ��?����oZqE��'���C�ϟ?	/L噖i�
���'��)��Ӓih՚��3M4��R�'0m�蘱ASh���,9�u�
�'��mŊ#ƺ`Y��*-��%P	�'��3FƢ��L�5�C�h�i�'[BL*2@Rj�|�gH^
5�ֱB
�'gFX���S�6�d��%g��3P^��	�'-|����N�t����"�-�d���')�	k�@ 7���,�\�2|���� ��������	��@�&K�Q"O~yBP�j�x��W��$A/6-��"O�񻅭S�4�����J�e^�C "O��h��:�3莢=$r�!"O��ǁ�h9d܁!��;%��S2"O��F�)ǈ��D�ת	���"O.�*n�5�@�Ȓ$E�ݡ"O�$8�E�c2p�c�\'�L�b"O(�s��X ̙�Cf±_�@�"O� `   �d     �  �"  �-  �8  �C  �N  �Y  [d  #o  z  ��  �  I�  ��  ߙ  #�  w�  ��  ��  A�  ��  1�  �   `� u�	����Zv)C�'ll\�0BKz+ �D������b�6�F�y����yb�҅w+~]�SO	"d��G�	�}<��2�"��3��M��1�cX:\'�N��r�ɞ=n���)H ���+ɀ>
�[`e�-��"6�	92��b��=CR�t
�i��d੭� 	��'�?9�g�x����mN+V��ea�.ĮOwRѺ��F����)5����t��6M#)S���O`���O���&c����g�6O��TȅN;B��OF���Ŧ�'��j[�gf*ꓚ?Q��_N0|�V�M ]�8�&���?���c����'���'��C�$�uW��5k�����&Էm�f �5�̩c�8I5dO=-`��F]��Op��&�	7`ڦ$(��

��Ȧ �b�X�yӫ]R}�<O��Of���T"��A/D-�iU�.MrY8��]�s;b�A��?R�"�'���'a2�'��'k���{�@��r(�MB�+�U�=�c����q޴Yڛ�r�^do��h�4)� y2�i�`5��Od^���K�x�q[�A�)>tj(��8�W��XI�+�	�W���a՜@���R�%3f���L�;P�	��J.P�h�'V�]����c�2�o��?=�'YNq��'��b�(ꥢ�7J<BQ�3c�yo�(E�N�r�㈲G�x��o�QDFE����rܴgΛ��{�N�����m3`�ZRj�\̾��B��+��T���(�%`cӎ�l�,�M;B�J�g���Z�a�W,T�P����wj��4�I�<V�Q4��/s�aJ�@�:ӠT��V��G|ӂ,lZi�6��q⏭	n`��S�9XxӇ��Im� ��3M�ar���M0��47b��e�1H��D���?A�"��2x"�� NJ&�,�(���3���D�O0���O*Ql_��`	kK�����	Ą��*ё�?9.O\���O���Z/4��ρpKt&ך%B���	JG �#I�&�<�&6G>8=ٗ�IO@�)k@O���^��dV/rK���1�U�#3ֽc��1?�b(h�*ҶQB��	$]|˓��I�p�pm�G��_�-c5ƣ	�H�D�O�D:���On�Ľ<Y�Lkj�El���<M�!�߉[q�����?9�!�_z`�M>���<ͧ7�I��c�<�{ԈI�[�,�.\�?A.OL2�K����q�'�yG�8w~�٪�oH;W�D�YZ�����y�bP2uM�x �� �q��i�L-i�d-rԦW.Jjq�ŗ7V(�;Pa���d�5X��u"̜TW<$�f.M�t/h@��-Ȍ����\��ikQ���V5��E x��9������M�w���|�6.҈-pR �0M� �K2�x�I⟰�����D�$)��y��G:5~p3t�M&�hO��D����"޴��وX�X@T����8>�\p��,�<h؛��'�	;t`9�Ɵ<�	ǟ��'��	�"E+��5����UF9�7	P2H���ӌ�	#�T�)%@��{����?e{����Qa2��8(@���=BǼ��B�7�rMj�GN�(t\eRwU�+�NTұ-3����R�O����`X*5�Me��:j�����xӴ)�'���1���ȟ�'
@���zFtH�R�@/AKr\��'Uў"~J2�Nl��Q���i6��7�?���b��gӎ�O�)៴�-Pڤ����+.e�<# �\� C���g/�I��`�IfyU>��'j��Ӷ|^J��2P�K�Npˆ�Z�Lz��S�ȀC@-�WK�*^�n��W3ʓXx�]�Q��.<jr)"�@� ]
W0R�"�p$��%�� ǆ��~X u�̖pQ�t� ߜ)\f���H�V�ļh���!��d�����D#�I�>h��+D�]�V�j�I�I��@�	ҟ���l�'�1O��Y�O �V�]�`%�_f,L8��|�Jo��ImAyr���6��O<�I�|��z �C�W^8E��o[�����<���?�O��0��ߏqq�Mj�4FϠL:����*F%O�1�\ �7��.AE�D�SV;.�<	��������`��v#����^X  yr�;
�e`�*.��͉'Φ�ם��&Ϧ���)�M;��iy�BǄH���	�y���$/E[�	æ�s�����?��}�b�Co���3a�C;��*���J����?A)�R�o�!;i�@�K32���Xg��-$��)�4�?i��ivx\�E�0<�t�s]����&�MC�'k�tͱB�_�x�n�C���B�������?'
��&���jo��.ѬM��SD���>ٸ�.��#	����_i�����H~b��#0��0 �$R5ч⍳;qp��k�9�,c�O�X��礗�ըm���_�"w|��O�Y�0�'�6-NR�Q�'J���3F^�e>�U)��A�2̈�&����M�	ɟ��Dy�F� Q���� W�a���A��"?�p�'��6�'�<6m�O@��e�[�k6J���f����'OڦQ����I�FL)c����	���ټ�QƜ�+��@˱TQ�̊��	" �ݱa��6R�R��*<�z�O>�d���"���'��35��Bm4#���.6�,?eB��+b)D����BE��UBFT>�C��%+��݊-�:80�族��{���Z���l���DX�^�"��'���'Gd����_��a�qC�<~h�p�|�).\��$2��
c�ěU����OB�nZ �MI>����+OV�
Th�#I^��Re�=
=9�b��w�^�l�˟�������'#��|�c(@d&p:�ɲ���.�SԘ�I�%B�)U����8i�(4��@4��<	���p��8E�V�W�\�mนj�~X��@/�8H�MõN�I�8pIdC���K�8@��	szL��,W�;��$�&�����+�4D���DFxR��������1���a&�Z��?AI>���?�)OʒOvX�Q���;�q2MO� �| ��C�O��m�؟��ߴ\l��]>m(���M���?I寉4r4��Ҧَ,n�}����?Q��u�ؐ��?��O5�y����ey@e�N�b� �aR��֒\��*F䁱<�Z%i�钽�����Ӓ]g�M+�"�����h�L'/~�qiV�6BW�|Ò���Tq��V1b�R���,uQ"� ��ؔx�V�!oT�	�8��-�!�d-#����
I�>8ʒ��'J���OnU��a̝e$���G>h��%�|.��&�6m�OF�d�|"t�M��?Y@��^E�(G�� 3��T����?���z��{�Go��1)U�ѡY"*�b�'�l1z��r���������x�'����v�G�hq&��1��7q�>� �!�(a�V�E��,��z��+?I�������E��5O��k���60w��9��܊f�4ػt"O,�C���<wjP��/J������h�D��۞;Ѽ�#�(Ļ6�͉7hdӪ�$�<�p!������?Y���$K�<��ف���<$�x� !�C$�mˢ�S �L@P �8;�L(�F�|��'6���1�GA?�ݢ&�Ax�(�9�
���.��;������B�(����L�Pc�P9��)F�s.h
�5�b!A�T�N���x�� !U�C�Jf�HŔ'�	���jɟ�'4!
p��zd� 5"�G1��'�'O�V�,��r����d��Y��EY"d2���:l���')�7����ɷ�M+.��i�|�s,��:����qe�X�uOO�W�8i��i3�?	���?���L;�n�O���>%��
�&>h�Hl�5a'N�^���c�a��$���r�$�Hx���F�	2 ��i���0dN�H���L� Q  D�F��j� �Wx�<I  @�s?^m��B�^��9�uU,����OL�=)���ܝ0\��#��a��|"��,N�!���	1L\c��j.}�6/��'��6M�Oʓhz����V?��	�g�V�P��2t@�Bp�Y�$�xH�	��8K��_�$���|��F�)#A�mss���I"4Wv1�C�u�����,bt�����(��b�4NN���'V`p�r�� Wu汁3	΢$(��3�@�$��П��'Vj���Hk�M2$NA� 0�`N>�F�F|q��R�d�A�
�}ڢ��<I��T>i���R���ِA�XGfȱ��Lvì���[y��& '�7�&�i�|���;��q���-�����I�\-v�8���?���D�(�<d��������B�0HFb+�F�c:K�T��PوJ'́���H�:��&%��{'Q�#L��t�R�h6�2R	��Dp���
�?E�c�M�Q��i��B:[RDx�,#?Y��Ɵ�ش ʑ>�'"��3��r��8��I�;��?����~R�`�
&@Z�*���/��u{�ŐG�'B-k�"8l�@��
0�VjTH!gZ�kcN�(>	�I���������P�LE�I����� �;;=.<
���0+�ѥ#B<7?�܀�A��'��!���G;�C� V�'uU�`
ŭ����a�%�TY����t�����S��ۣ߬%�,q�A�Rx�s�_|���I�5K�w�H�%kB�$�+ �T�Z��������h�"�'�ў�a#GT����q䀿bW��-Q�<�E�H�!����f�G�J�p�k��џ\����HO�	�O�˓I{�A�'�J|j��]U����:w����t��O��d�O����*�$�O��@�ni{w@�:?��E�5Iԭcx�"@�7wIj4��L�?k��7M�njJ���$ʓr�p1C��*N����19����l 08�8d��^�nZ?*H�c�⋜3\�aė|₋	����7�I�		�#��p��?a��D!��8�5���=ժ�3�*	?��Ԇ�I}�%=j��7��W�eز�֍g0�&��#�4�?�-O�=��]i�D�'~�}�@m�{�H0��oL�\>����'�#�8,���'��ỉAY�5��@�uk�U�n�6�Pb%���\b�J6�˩D�U�b�>VFh���򄜒Qo�`K�ǡmmX�[U��&l/�\`���S�8{����OX*��PJGv��Hf(s'T�O�H6�'_����k>�	Sկ:YJ�+�%��#�Oz���� �F�zl�!�)bꦕA���=��|'�'9�iC@(F��#ž7�ʀ����Dш"�����O��D�|dh\+�?�6�Y8J�Z'���'\%��kƠ�?���}B�I1AX��&,3 �O�^_J���?Q�OLެh��Y<���\�t�RA��O����e֢d�d%�У� !�p9+4D�y�'4 2��s �5bv��疶m��e�'��H	��?Y��Is�pzsfڥOb�寧X-:V����y#K̰=!Q��`H�(S�P/��O��D��BD�L��@G�T�`���zӋ�Q*�F�'�B�'YƤ)\�'���' ��,#����� �(�T�:3C�&O�R؁`��X��D��	Z���E��d�*�z�_�=�h��B�M�za耊K�e�>��,�A5�y���L�uA˓ak(� �=�n��̀�^��\��C~R`��?)���hOxD�'c��+��b��S�lI0�"�2D�L�Z3.�;���a�Rqj,�<Ʉ�i>5�IlyBjX\	x�(7\@�8i�R)HF}+vF�,40��'���'�z�]ȟ��	�|�+�8mX\����(1�&P�%ڊT-������;jPKϚ6ZHua6DӖZ6R�<)��KD�? &�z��O��D�����8[��'�ү��L����~A⌛'�M6�A{-C�)���O�M{��A�D�Z
�V$JH"Ѕ	&��'�ўLFx��F�9���Ü ���8�-$��=�yҍԾ%�p�&(Q(	R�x`/�>��W����'�ɤG�Z��ߴ�?a�4���!D�8����W(ÖxW@�����?��͘��?���?��39�hTj�EW����i�z}�W�V�l#�/��t�Zw��?@���Ey���/;x�R�)V���e[7��&P��x��޾MN��5X0Bm-� ��jS�M:(T�F�I)L�.�d�Ѧ��(O䄋U�ϫ0��g�S4Y+Rͫ��|�U��E{�Om���@B�,S�D�wj��(P��?In��Xd�99�B�P�h��D��CN����4��$V$�7-�O���|ru�?QR�ʣfFղ��&�妘"p����Iԟ�1� }ʑ3�0a:^H-ع��i1R`��4F� Xj��9�v���*Sr~��E\�m�0/Q3S}�|4N�{�h���O._]<l5��#J΅Yf��d�"J�O��5ڧ�?�q��5�|�Qkjp ��A��y"nZ�N�j��J�.��A��-�=��OĈE������0q��������4,@�Rm���'���'�:Qz3O�v��']R�'����9��A���9\晨U��%>�`�3��?6�u⠢�
S.�P�1�	T�cZ���'JM�(ާz�L�sÌ��(7�����z�>��d�;��R"���O��0�%�p?1���M��dـF�1!{8�ؤ����'E�p���?y���'Z��2�])%4�i�k�&p���"O�m o��Z�p��V�Z$��Z�����4���<!f�����u��L! Ly�N��L>8�@�ܙ�?����?I�R���O��k>����ـ#�4�A� �@�>�CC�`�\0�4B	a�-"tE��x�I��Q��0B��P��Rc�:$�����i�l���V9%�d-"�L�M����Lأg�Q� bV�Ҟs�������*P�Љ�9F:���O�=)��$��n�\�T·_��Q����!!���a���
�R�	cU� :q�'�6��O��S�f�Z�P?%�	3m�)E	۲5޸ bBP�jC� ����� QI�ϟD�	�|�����%��Da@Z/"����X�a�"
;<�:����8#����	�!%
]��(����I`TtHb�c�.j�~�R@�տg ���g�5Oў 頋�Op��??5 D$M2��5�px�� �V��X����J��8�Kb�ޔV�P�%*�O^a�	�\R�0���oc��3�Ѵc�D�$�<���Qқ6�'��Z>��������$m�WF�݌9;Ө7L<��'��ɘB+�#�����J4 ^�T>1�O��eP�Ѥl|e�1�|���O�Dk���<G4D�A�%8� Z�j3xB���t1�T+^�=i\��v"���������O��d4�'�y���>Bx9CA�Ƀ��5�֠�yR��=kn�8��?��r��Q��OQF�$l/Vvt��'N����&��}Û��' ��'��a��V�X)��'N�'���5&ݜ��ͅO�)q#����6�S�J6>n�Q��ے1�m��iW	v:���'] Ы$�_Uxpi��q.��Ӵ�,p ��A�=��w$ܫ��O�ށ8��Qp?q��K��t8�a�N��F��դɨ���F��	z�g̓7�DM�%��_J��;rC+��̇�lc�9cӭ�c���(���p��'#p"=ͧ��|<(i:D���-������Ɏ���#.�tz�=[���?a���?)P�����O��,���s��t���d���Z~�0�s
@%P�dA��x����I�g����� UU��2��ݡ$0�LeD��]+��QD
35��K�d��h/�}E{�׊s�Z�Z��U��4�c�=4�������?ٌ�3�f��zF�'q4����<IN��ȓt����U��k:��!��wc�e&�@�ߴ�?	,O��b&@�~��'��Y���L��28P��Q��VTğ���+��q��ß��'f�L�atu����$ڇ�?�Q���[�jQ����	��a�@��+���3�>�Q�@3�$I�	�@}q 3�G'_�d���'��/����dØA�'��I�N��(��_�t	��% 8
�O��� !cD]�a����ƣ��b����OL '��?�v8ʆ֭ר}�w�'���&n��|�޴�?�����iN�L�v�䛊%������+=���1B�U<��O
��pG�
.�XY�eߒ��X�l�2
zD��d&�4?rb0a�����ra�Bc~�b;�!ц��t�H��A	䄣!��ZB���)�,<�����|*���'pq��q�ɧ�@d9��F�Z�y׏�9|[�Kc"Opܑ0��w<������S<U���	��h�0��s��+�|]�3��$8�	V,s�l���O���x�V]Ke��O��d�O���h�=S����u|Y�n�@�h�H�F*uԨ������$(E4`�b>!r7����X��8`	� �X�bg�h+@��#I7�� 0"!k*��DD֜+���'yB|��!Ѽ� �񛣢ޅ"�z���+�%#�Q�'���*J�d�OR�=Q+L c5B�R�Q9f���y��k�^a�Ơ>d:���JP!�?����SΟ��'�FD���J�l�S�ѭ~ݬ�jW�G�X�2�1�':��'��O��'��ɍ�btp�%�2 ؐ]J�ƒ�W�F�B��L��C�+�>p �٦�Ij�':����%"i�%B�^�K�r[�%_.���Z��]��0��G*-Q3.#?��ւg�T�
Q���J)�w�(5%�P����D{b��*_g�A�-Y3"��$��y]�C�I�h�LĘHƒ��Q1��ԟt���O,�n�x�'Y@j�Au�P���O
��&��*H�oL�4Ѫf-�O��dL�R���d�O2��Y=�F�C�h�Ѣe�j[DIJ��
ئ��1= y)�T�T��m��剶ȍy�@(-��(6�ِf��1���2$\���.�5�@L��R�*��-;YΔ]H�i3��	���s���'�l � K��C^��	u��݈L>ٍ�d6�/[
�@"J�fit����߼Tw���G{�O,�6��6?��tjN��7EV�C��
`��uoqy�K��X�T6��O���|���8�?�R⎁d�nD ѡ[�v)�A�ӪF��?I�ZdUK�",
�*TDdÛc�n��g�L@��˟���/��%��U �G �1�Z-������ȃ \C�-[�h�>�R��_�=����@�r���A�2�G���q�S�����)d2�.�ᓪP����L�+O(c%/�G�&C�	_��H1�d&��Ju��:��?����_&PD�U�<`�s5(�Oym�Ɵh�����I7���X^�|�I蟌�Iܟ�;ɜ(P#��L�ɲ��\�р��͑�2�	*S� `0�*�3�5Gl�i�[8.�B���k8~�Z�cOT�M����F}�;D�+��A�I)% �I7Hn���Vb��^@��lڸ��$���"��'���'���S���>�PsC��H�`��$"O䠄*)&0��W-ӷ�ԒP�<{��Dퟨ�Ķ<�q��%#�dR��2H���R}2$}cd%�?I���?Q� ��N�OH��}>�97�E�sg�!��P�,R�8s�H܏E04����)q���p=Y&�L���t��d�S����.@Gl� ��C-V�`��E.3��T�����$k$�c�
@D��2�ԒS�'�6��F�ş,��_�
�2�B�$Y���j��!���'�:|�UG�$%
����f�Ҁ�H>!V�i��U����mݦ��	�OB1��cB�RQ����
�+ �MaG,�O�D�{�����O"�S2e%U��S2ML�hD�ϊiI�4��̎�)D���
��E$8�Ҥ���L��ɰ)^Vi����Ui�}
�dF��֨ɕ� oZ�g̊k@tZ�ςk����g �B0%�����O~�D"?I5OQ�HL����2jd�%@LC�Is��J`���A
�eZ&*C"�[��9��E����Oxu��+�X��t�tE�&D]�U���'��I�RRm!ߴ�?y���)�[�����	LX�a-}X��e�{�<���O��D�ZqT ��h??�Oz���K���pdР6�e�U�λK�*�bj��R�މA�Z��ᓼC�(Ie�#2=�!˂>,��D`�8�ɩ��S�OK��I�
���fCC<���'9��ңN�?�B��<m�Ha���PE�O
f\��䑨jE��k ��o��2��i��'8r�a��q�V�'���'�R8�2��� H[^p8��*��@��(l\`a��i�IK����F c>�:�'�'!(�D@8+<��u0���Ҿy ���ΠY��F��9�E��뉝��O[84ʇ�Ҵ�y����P�p�Aa�S������ذ�?��OB))S�'kr�I�&���`�*��`��X���y���h�+նĴ �T�E[]t�Iȟ����4�����<ɂ��
���f��u#�(KK�3����E���?����?q�������?��O�,D�#	���	Z�����!�nQ�M���'��q~��3R�[�ȭE~�*Չ��+SOs:.���]d�bwN9�İ�e��v6(��"�+�p�ȩ�4���[Bn\�ծ�C���Є������y�'��hzC�/J4TJr �?T֪d�H:D�̃e���0j�J�E�p�r%$�������INyrf��N��'�?yg
.5�$�B�ʼ#贴� 'D3�?��;^p����?Q�Oeh��Ê7�����I;1�P��=.�Z�S4�K?�ܤPq!J�WR#?A'��8~0����͗==ZM��S�N����t��TQ�`�-܈V�t�4��O>�q��'�R��X����.�Uh#
Ϝ0O|IpG�3�D/�OX���Ո�����C?]? LB��;��dG�aD��K��dp{EB�?i,O����Uɦ�	��̗O��)S�'�"����W�Ԙ�&◲s�M���'��JG2WK��:�O�<_��In�8	ڸ=@�ˊ�R�&�'*z�x�5�5����.ԇ%O:��'||X��P 8-�@c�ccӸ+UJ	-��z��Gz�f�)fS��*���$�@���x�ɏ,"���O��}򛧀 �lY�)ʤ�m�0* .kؽ�"O�uj'j�S�|�Y�Y좁[��I۟t��D��K��h"�m6J�����Q7U��l�ݟ���Ο����Țu�h���ǟD�I�\ͻ�,�ulF�bJ�1�$c����"�ܑ`���+6c^[jh 0��G�'l�'q^��b�=P6�	aPMX�Q7Cq�X��`�f㗐2���9vc�(��O�ZO
�[%�>[����RM�alHc�I(�?�3扶7w^�r�jE� ����>=��B��8��P
ʎ-�>8�^~@�ʓD����G�Ik��aR��!w� ��<<�l@Zvo�=E���	ğ�	��l��ğ ���|ڄ雼B ,�bG-�Bm��//G��Q��F7E�rx	�Y=X��Uw���Bh���O1A�° 3�	;=�Mh��O�N�J���@:���D���Oy�V��5l�4�dIȠ��cR7k��'wў�Ex2��/3椌�Ѫn/n	��N�y�a�{�H�S2��4#d�,�7k
���\��v�']�I-1�R�Ҭ� ���?Yp�v���t|��u�ܲ6���O��:�O��f>�U˅�uQ\|��Ñ����3����ktD�jE�V��d��իV>�j��ğ3;ت5��%�%z��H@��+:��qrb�F�(�҂���(� |�����cT��=�v��⟰�	p~r�ϛ )Z�r�M�&ri>�CGS����?iӓzz�s�o��p��}��a
:�]�<���T>�Q�|Î�� ���r�X,�rZ����IOyAH�`A2� ��I�|���2��l)�h�YL�Is��"��W�O��dF�$ `��eE�x��� c���"|��⊝N��h�F@�t��"��S~ҩ� R4x�"CD3[����퓥>�EA)C�FE ���Ø�r�7����	˟,D��3O��r6i�'	��I���3B
��"O
�p�d	6~4�I"�� �&Lx��	-�h��xZ�AQ�Phe{W�f�P�P$�'��x�W���Ҋ���8�Sܟ���Yy�� �55�4KÂH6pH'��ui�\�}���M?J;tuQf��I�t�ڒ��%A�p�$M9&���Ѷh4r�$� ,b���	���#��-����1r��TCBI�O`��"ړ
�PE	C��m���gA�w~� ��'����5�-v������v��Tk/OH%Fzʟ��U�,��a��bئ��5��h����޴30�,��[�ˮOҰ�r�͑�?!i��l�]��v�sȕ�o�84z�b�+:�T���FM�I�8�ɼ#ƞ��fP�\���sdD��?�'Znx�2fW͚�ە�زx��G|Bΐ[?l2a�]!J��*e�]����)gxm�@_�k(Z�3�ԥ�O�#��'FR�i̟wd��^�`Ls��˞e��x��L��Ǝ�b�Xxc�S;*16�b��7?��T>�K*O$�����,f̖�'�]c���Q���؈�M���?�,��9Y�l�O2�״h
ĹPTD�)P����h�4�D��r1��[f%���W%z���!��	w�I��t)�2D���
`�ߣK�hP�+�yrB74� ��R�3d�3/�/�" ��/Rxܧw�XF��'�CWǓ�?{��f����I������$����z��Za$ދ5!�H "t^�kp�߸*V�#�l^�ў�؍����z�{deV1Vj '��X�D�d�O��DS+S`��VH�Oj�d�O���F���+r�T��R���B �dǟk�������{���CBb���)��m���PL�l�&遇�xd1���(�����Y���)�M	���8�B*G�YQ��O	Ҹ�p懲��ဘw�p�G��(J��C�������O$4K��'���<���/F4TA���D?.�n��emAyh<��K�>E�l���� عç�?�?���i>q��Dy"/Q�@&��м���0R-�*]4�x���-P��'���'7$�]П����|R�d��~케�h��H �Sc	9bȤ��C��	+�F�RӪ�;5|H
ej�k��<9B�֓�xCR�C�uWY�#/_7X{0и��V*���P��	���V!o2��<�[�(We��\��,�#�֡���#Ο�F{���![����&BZ����
B��.C�	7�S��� y�<�#���d�"�|����'��	��$�鯟���z>���].~�6��<B8�%(���O��SL�O��D�OΘ�VnM&
��M�
V$tQȹ)�,�j�씈���$d��\�Sk�K� �SC?�Q�p� � ?S�8���ϛ}t�����2y�ڃsu��:#Kז{D���'

��I���v�ɋ�����Oc>�01�X<�y���֊/ǎ�"g�<Y�0��0�Ǭ��^y��b	��ł)�5��|B6^�l�"�L�2�|���M�!n$��e�<Y��W�ٛf�'�2T>���ɟ����V{
]� �(M�0I�a�T��q��'�4%�W��g<�I�ʔ<e{�����yt4�|ғ F�J�8��GOs?6D�բ�<)���V�H�a
iAȹ���J��Xe�BIQ���.�Ti�fʚI�����9�.̨06O��$�'y����@�S�? �h)QoˬXA�a��U�D���"O��(�c�A"���B㎏U~n�:V��O�Fz�O;J�CC �G�Y�����)bd�'�'&ґ�!˔�@v��''b�'��t�',����bђ8�T�P��ݯ`�)a��G�-!�铋Oc��z��*7w��> �. ��>��	{HFIA�MԽ61(��m�h1
)����j�[CH�Q�N��.��Ĳ�I����>'�nZ<�Ѩ׊��O� ��`�]j��ɔR�j���OУ=q�'��-+��@�(����gW�`DE��'�j�ç��rj��g�9@�m���'��"=ͧ�?A+Oh��q.F�o鼤��F5!�͹�	��3| U�B��O���O �������?i�O hv-V��D9�A	l	"��uO�~�� I� qVxӓ*�����nT�EӰ��e�1U;Jak�,B"˜��t�ғ0�򶣐&Q�b���փv�O�����'}Ȁ"A�E78]�be�1��1��'pў�E|2����^ت�!��;��S��%�y�@ӧ;L���7E��X�m1��A�������IZy���%�Z�'�?��O���s+�z���L�59��� ���4���?��h�t=���G+.��)�ʞ/>��%1�m��7T&��/_4fp��!��3�.�փ_d�'m&�SF�R� 0�3��ϊ�.i��E�k��] `�5Wp�<���:�ȃtmS^�'�0���?�����V*��+%�߄G�Z	6,_����4�O0�G'��,X�1	
:)�!�r�'�j�gSn�{c��5;��u�uDǌq;n��'�2�'b2Q�p�O2"7O���PH�*b	p�Y�▏JQ	2�U���?�*O%ԧ�O��#��Ԥ<H�`ؓ.L�y�ҳi��'0�%>�"�X�nm�Q��+�9fۼl��*�/�M�i�t%)�'3X����?����?ɚ' P���V��4�2IE�:D���7D�F�'u&��2�'����I-����u"0����ص�'�� lPjЯ�D��r�]�?i����UX�''���O������y�4k@�Q0fHX
"��<���S#		���D�O�����O���0eK��s��n��y,��RJ<�P�X�
��`jS�s5rA�#�?��e�8u WS?5�Iڟ�������PE��+O z)� %H�[rP���a��'���B�'��dީN����uǋ(;�{��U���\ tn��+a�܉�4a���S��?���8��X?��Пp��1G:6���KY=��Ȁ� �Q�|����<��L�4��,�u��'��d� ]��i.|�2��� ��1Z�n��+���Q"�P�#��6-u���@��Ҧ=��4DH����ug�O�T���	o� s�`�MU���b(.�X7-�g=�	�yWD�m���M#�'�?�R�'l^u��4@�L��+�<!�Ƚ�bC;;�z�y �i9~�*G�'W�$~Ӽ����	��'���O~��2����$D�;A��8��.D�` m�|�.4C$Ɏ��YR�	l�(�d�<���C`�S�X�����ɸ-�h�d�ո ]�t�&aP	~�	��OH˓�?q(O~�D�O2�d���Q3Ą��@�Cj� ��VCh��ʓ�?���|J?��Ɵ�]Ba�b"APM�P0���"O*ғc��Qk�m��$� -���B$U�؆�I�z?�91�@�p���R��8��OV��䏺�ęU�W�>2ͩ�&��!�$9������+!VxSD��!��6\F~���LZ|�V��"^:!�ϱG X�' n�bDڔ"]v)!�$�1%�
� �2�`7��/b
!�䆇4�(��2Fߚz3���[�Ș�"O���`F�
Q��X8"E�6P�C��5KT �J�&�/֘8s��eZ����Js
t'iN�3���"�˓���r�A�f���I���(Zd�3K��OL���m�6o8�)�}���n���ŬE��}k������'�9��ۅylH�!���4	����@�-x�Ƥ0#~�&$	2��r�@ϓ:���jrc)k^�PC�,mg,�Ȁ�7
m��k�B(.� p�5G���j\+�e�XRP�b� Lf�Gȅ摑���3~|"$'��D�eI2C��`k�����H�]80[�nH�v2l�޴Y:M@�xtG�
�!Ұ��E�'�"AKr���דza±;"��Bd���ǋ��ӻ76.urw�'A(�j�,E�m<�O�t�FNԑ*��I�A˾^�DIZG�	'a�HٰIC�\��+Ie���e���Pa��µ��X≌ ���d�ͦ�`��Im���S�xQT����߻fr.�Rc�&D��:���4yB4z�a[�e�x��J��hO�ɒa�'�b�� 7B8�����L$��V.���%�������'9HpG�[Ɵx�I��<���l؃X�$�%� a^0�9��BN�!+�)�>z�Z�o�$?-xh�|rCI߹B��d\=+�����9C$I�Q!��\:�i����'[rN�W�� �|���Q=� �-���i��ռ󦢜#����`U42�a�F�
or�7-`y"m��?�'���x�AO8wi�Z!�L�a^6�����y�kG=@�82��>\�.���f��~�'H"=�'�?��O|Q �+�$~4p�JçYk�	�t�W�,ot�AbIFǟ��	����	��u��'�8� ��=i\������m����4�ԥUV0��4cU�I/���єuE��S&"�&�(OB�� ��W�N1v�CwdG"O.����	C<|d$�q�¸q+6l�GՒ������}�4"L>�� ���@j��M)V��Se�>��5���M���h��ТuK�'xm�%��LùH� ��r�	�ӆ�j��&�Q�3��k���b޴�?	+O���Hc���i�$�fgT�kLiB$�I�q�~�����Of�D�6 �����O��S,��r�Mƀa�dI�NĩY���!��ȚL�b�UbI$)�"���Ov�[n�s����p�z]��@S��p��%���
%��`�;L����"j���'w��jش�:S&��Z�Ӗ��h��� ��	�p"^�B�ʙ�(@B���R(RCቇn������R��e`G#G�4��r�����'�6,��i������I�K�7�P~���;�.g^�z7%�= 1��I柠�f0@=�a2�K�F�K��R�Pk��~�v�O['�\�$�ֽq�f�&��J�9L�Dq�$�K���Y�L �6dˌ���YƉFH7v!�@D(��ēm�B��I�8G�D�i�L�K��ދ	Ğ���hX�B9jj�'�l�E��1�X5@�k�4�ʝ`�pcQ���(ϐk�!ۣ'٥oc��[ ��yϛf�'��'��:s�Y<'���'�B������ŏ|  <*-X-�~� "��(��|�U�͸�H}��N�*�������TU��rP`��/�T�GI�
A�eQ��%YpA�`�I%J⎩����O��Aa�f�Ua�㈝f��e�� ]Y����J
=�V��<�]ݟ�w�L<9�D��=D�Zb�=*>~E�m�R�<�%��8eE�;@|t!�EJ�$�u����'�I�.�8=�B�W�k^�zaEH�@�R��|n 9���?���?iB�����O��;e[��cD�f�����TD�1P��>�iǌ6WO�Wr/�d�`�I�>6�5SWg@�^E>(�W�/+bvr5�߲u;؜�4@��I~e�q��9`B�"T�I�C��L`�ŚQ"��b ��,��ɘ�H�O�m���HO�b��Ge��W�6XX�&�Vo���O7D���	�yr�ɲAL�tB��e�*�M������1	�4�.7��.΂�����5V���� 7*9��ܟ�i�'�����|
S�AR�#�E�[j��A���V:Dx@��C�-c���s�H�bw�0CFe��pD�<��� �q�p. �T�xj�#�=B,QBƹ�n�Fv%�Z�,�5�!�S� ���M���O�D�SlP
&�~<`��D�>��M�4��+lO��:s�D;p�tI %�!�Dہ
O�`:Uc_�@jԩw$�R�#·G5���<�b��������O�<���i>�D3UaJ]Ȃ���d�ڹx��Of���g� 0h�WxP�RV#h4 r���S���>��Tǔ�;w�4��]8+	&��wjΡG
���㌹g�Nc$ ��q��rDT>�r j�5��x@#D�L.n!� �.�d��j��DhӬ�F�Ա�r4���ސIf�/`��	$���Zl!�ę n@#�m�u�����HZ�x�b#��,�"���.N���"��B|�(P �bӰ�d�O���3n"��ё��O"�D�O\��w< �;p�P����P˓�{F��IU�\�֙��
��<��Q��D��ZR"�'���
S���	�<���QG�Z/B`(�ԅ_�/FX�K@�Q�G�BQ[���py��Z ���<� Y 4_>}�$�O
�y��g̴�R5��g�|q��!fQ|Hn���M��*]^�@�S�gy��i�嫵!�?*{�L�RHV���=B��O��=E�t*ԇJ�ЈZqaφYaʤ�"L@��~��'�6���!$��ٰ)�?=�'���S槜64b2�ɔD

Z���
[�8��r���O����O��d����ަ�����d�$�.7W~DJ�k�8����io+d|s�˸d�����6�P�E��8]}��Vm�b���R �[!f�6�'��;|��0!7m�u�'��ai@ ��-�v�C%m�����M�wX��d����4�?+O^���<Q�O8[�bU8�B%�ڥ\w��J�"O��K������B1B
0�L[ŏ�I�O�L�!�4��䖁mdx�;�?�4G�n<PwJ�&R�YJPf.N$vEs��'��/	i��'�b��;d��`	C��y^�i�P����:P�PT�ǧH&	� `h�Q�z��IC�vz��X��ޜW��w-)}8$ՙ�X$0z��nT8F�����!��O��D�W?i���=YJ"pzU&�*��(s�a?i��?1���'���'g���Ks/�a��Q�f�:�)��Px"ʉ�7�N��H��r5w'�C��{#�q�l˓=`B��iC��'���D�8mZ.Sz�b��$T�:1� �0,�����?��ɟg�����O;<$�8�0N��l�:��X �ʪ�DU��"�.(`��ī�2o5� AA�x"�ۛR��<9ᄎ=}h��Y�FO�x��uKK $\t,ۇ���^�n(�B��*e:���I1$;NOzH��'�R��ui��I�9Ov�C /�ZF@9��NX��xB�#<L)E,R�l���+��Dģ=ͧl�Q� `�F�~f2 �D @�����6��O���OJLӇ ��Z[����O@���Oǧ_Dz��@
�:t��h�.F(O\&�@�3��Ҕ,G�_�T��$�?�S�_��4���'rHz��ʔKn�TR�O�d@f�c��
�G\t���D�>L�րY��Wer�fM��`�n���=� *;'I��w�D�Gn�=G�tp�ß|�'�4�"��|���'#�a�6'��c�6�觮Xi�Py�'��@�ԠU�^\��G<���'��8��|������,��i3��";�����$38�;'��.	4R�	ǟ|�����c[w��'��V4M<`#��Îr����vEP�YHa�6%��l�뀓yG�L���td��"��$ĵs���ZR��z=�����+^���-�d`C�#7|�fqCV/l��a�F�[���&�|���JY��'�o�>iᖠFz\�$�O�3�	e�'A���@�%u.e (����A≧DK��遄��	b�&͛MMR�L��4�?�,O��S���A�I�kQ��KŎ ����>b��d���ӱ�?9�Fn��{��?i�O�P�B�敵P��,�f`],+|�b��O����#1pr$�����2�"QP��t�':��O��2l�2- ������)�Z�0�ތ�8�*���4]W"�1q(h�xҲf>�P�2<}ZR�Ȓ_'Gry�c(��p{����"ODctP�t�y��,q���v����bν%}��i@�d\���TΏ�:�FdX|��9
�D6��O@�d�|�q哑�M����#]=��*��V�J�����R�X���'���ȇ̚I6�����>f8L\�v�M�h�$'V�h�� Ё%�u*N��F�x��Ft���5G�(�kZ�=Rb�`T(�3O��i� :��b��JL���I�s�'����N�ɧ�O��)jt+� ����8��0��'���At��!Q�MYw�Ƃw8�ǓD�Q�X���'p����­W1��M1C���K����'h2�'���4B_�I���'���+F�^s��]+�ȇ)D>^X0�٩QEH��)ӵݶ0뇤��e�B�ZU�	MU��!+�#B�t��a�y�p*���:W�d� !�C�*n<�B�=h<��Eo��O�	$�i���g��C0���h�+yP�F��:E�'~P��S�g�ɤrn�	�2���4��#�.{�B�ɬV��T�����r ��5M�jͺ��ğ�k��4�hOp�q�c֬	��vA��!z>�h���>���HПD�IßH��.�u��'��6��D��7c/:m����G�̬d�U�`�uCdߎH���x�)A�{�E�B��,�(O�u��fO����9�;�eI���N}$@�c�ύ1�*�0��ъ�T���`ϟ�dQ�H.��� ��M2f+�0k�2P��
x�V4��'>���dQ&�de1.	�A
��h��	.��|R�x�*<���kM��ҭ�4����'�6�8��Q�<TmZ�l:d�P�Z&��-PZЃ��b���K���?1Gb��?y����Th�A$�����U�U�`qg)Z7�>]��`A�%
N�pR��7bPu���	2E^(Xv � >�@�1�JB*s�0�{%�.�6]r�i�w�6��ď-O�`���'3>�'�9�`�#7Q8��Ԁ��o����'\�D`��@Č� 2٠aB�'�� ��.A�{^�I������7(�~��'0Nay�k�����O�ʧ-�;�442�uZ�L�q�yP��Ϫ i�@��'�rHYc��s@P	]`�v�τK���YƎ�h���u��+�Ƀ�	�V`@��]5Np�OR�� �z�,��Ɔ¯G+�yXVfQ�<�-��5H�I��p�F���!��5R�d�x2)C�?�#�|�������
�1w���P�"��<.�Q�'�<���/�&�㐯��}�d�b��Q�`���i�87b4\��PS»(Л��'���'@ވô�T0���'���K�,ǘQ0�l�D��;/sD�'��\0V�ǖ\���E�1P��:���+$T|K�I$���f��
`�B��[�)�X�G���]�|	�K��w�a�"��.��O����Ċz���0�N�)�H���_vĠT��,J`�'èT��S�g�I�-�f�J�	����Po2H|BC�	�3*�4K���<��!��lǂg�b��˟��4�0O�d��(M�<@g��/.N�C2�O����v��ǟ��	�d�ɏ�u��'�:�����V�cjT�ŗ)zD�y�� �%��:�gJ2-�)�� <ILuD~���7"n�11���:�i�1��MШj��~�I��>=���T� �����'i�TzE��+W�
gZ�*��O��8ړ��'�KY�(�f�R�Ҕu(����n�<��_��D-���_�!#*h�&_�nꛆ�'��ɉ-�L0S���7M�j��YWc�)`\�l%��q�Q�	ܟLDm�⟨�	�|ڥ�w��3&��)8E���T�ˤ��V܂q���D�om�5Q��I�:jz�nn��C�Z(Hl	$�S5)��:���1Q��R*Q�z��E~B��!�?I����D_�x�������@ ƚ!�qO,���^y3�9�G,X��,��.��~-��DZ��ݚ���8p^Ɖ���C� ���%��O˓Af�	2�?���j�TN�w����j�vt:����,lʁJ�A�(�d�O�AB��+x|\�,��P�|�3��Ӕ��U?���皣rr���nO�%�����-/�$�&"���iW:�$��h�(U�|Rv�ͥ(݈Hxwk����BS�c�	�^!&���O�}*�t�? 4�iT$^ 	f�R\�s��J *O�Dx�(ƺ7�t�1a�@�Af�$�gQ�p�bG��9�X�JǶ��4B�m�1(w���'���'��P��N �}x�'}R���ӑ£f.p�p��_�5gty��
.���c%$J�TZ0���Nl�����1:���R&4|(�J������h҅[e�f@�"�VP�ËR�du�U'�
e&��a2��|��g[ |E󎈜~`x;�ᒸH�|l����4���I>�Ĩ���>O�q	��>?��\�J60mZ� "O��Qn��GIV�q��?7��w�O��dP\���ԟx�M�i��D�-�Ч���:eY�mPD͢=� �O����O&���޺��?�O^�=K'NN�Ӽ2�̓ lvL��ۨ�xR�C� N��� D.����$�=��%�
�'F���U�z�Ρ0 �<K�hi0.��?���'m� 7B� R����#%��	8Lj�'���`v拁J����ŠA��ي�{2�oӸ�O��IR$ZߦY�Iצ�
�G
]}R!��
ǆ"��%lڬ�?Q�g�|Y@���?�O:��P��3D���6ꗶ�x����&�y�7����Z���#���K�'8�Y�f� �Z�� �,��;���"_�ȡP��G)2	Zb@ڧjJt�S�l���|���?Aӕ>!�K�5`7P��"'�$���Eq�<����{��1�I[.md�j%Jt�'Wў��M~��B�R(>0��P'��hP��5��[� 6�
��ݴ�?���򩒲2�6MS�yd��⇉\!6`(%	*+J4�����T���K�R����F�6I6�ڄ)Ҹ>X��a��Aj�t%즄3P�V�3�Hz�(Aԉ'z����
\���}���Ga�D;���s��=#bO��?�ƱX�ߋqV��[�_a��4Z@I:�D�.�2�0��I �4�$�
8��sEՇ�!�����|Ct�M5��(4-��#{��D{�O �<yu$�Nd:�s�C�08�����	Y�qFp7��O ���O*��j_�L�����O���O�CV6WsҴ�`�Q�VZ!��X���r����� ��t�1�x#�Mj��0@㛫F�� ��]Lu�u�34L�B�����!���TgM5D1�ĎR��X�!�v(�Q����숻M>i��П�>O*i�%)F�.�Tp����&z(:��u"Oڔru���l@̄�G@��V�y��>��i>$�XD��8�vp�'�5s
�!ʄ��k@pt�W��?���?1������?��O�i��\Y;�t@TM^\�ځQ��^��x��k�Up�i7V���������p
�'l�-r+S2�^�[�a��}(wm�2�?a�'�69� �� �|��dPaN���'��ԠU�P�9�rms�@�@�4J�{ү}�ؒOe��������ݦ���K��h���?�*x�`X��?���XY�����?	�OB:y�����*����C�U�ZQH�y�bp~иs�͔^�J���d�A�#?�q@�20jt�Ǆ��H	RhX�i!����X;b(��@�!y����e���^���D�C�i��I����d�@�;���u"O~5��ʢd-�y+B��i՚`��
O䑊C�!D2. �Fm�"dpR$G�,�ȒO��xR�Ϧ��Iʟ|�O��|���i]��@���N�B��W 
��z����?����e �qa�[�SU����5(\�ЖD�����	�����$��A5PL��F�#-��'Ĵ���4p<@H&Q�V�pabnK�s�pz���	aT��(0@�7wj$ꂤķ�M���;��I�o1�'��i dnx��vɉ�#�{"V~a!�$-W����Ǜ/�x�Q2~_B�F{�O{��<�'a��F�Q�B�X�Z�a��j�6-�O��$�OX�2E�ՍX#��d�O����O7G7p{*ux$�G�'r�)g��xSv�
� >?ѡH]�!���|&��ҀY�Q�����$�4!�49aJ�7	aZ�0�O�|CL�~&�P��l'��Y��]�Y*�Մ�x��'-�3�S�g�X�nca�
�9��pu�N'w�C�	�?6��p���՘�a�M�u$�'�T"=ͧ�ē3d�{��g"(%�/~^�48���y�dQ6�'F��'���xݡ�	ӟļ}+��0�e'��uy��*���RUf�w[@i���H,�2+�0U$ 1D�-ʓ`[�Q��-��Q��i���@	&��~_�ɠH�n��b	�`�L��C!ʓI46dc -�3m��)�oe�d������Hr�������!�&��!���t- D�`�%���21��
Nה^��QbJ9��MkO>Q �ޚ!A�v�'���#��(p��&{~|9q'�]>t���O�#e��O�Dk>5	 �;dV��8��\�kWh ���?R,�xP��ݝC�<Y��Vy�hR��ǝRfQ��P�`ѝu6�XA��`>�Sf�ɜ{��3���m6d��B�3OS|T��M_�����B��_�����_[��/T�t�׶4�D=�����!�� �M��CI�T>���u�_�rX��B���j����
���8	)T���p�rw,��<�P�|c�'��6��OP�Ķ|� ��M;��H9B.08U�E�\nV�q@�
�s���'���`EZbP{�D�v �8�F'H+l�8 SS?�R�G�a�8እ^���\�CO;�ϧQRa��A�>{/�D֪'fЬ֝�T�m D�	4=�����K+��33��"~lT��0�x�^5�?���|����ˁe��D�!�2j��k�aˊ�y��(i�L�J�!_d��#���4Tq֣=ͧ\�Q��k1�1,h�b��Ҿj���XF�Φ��&�'P�'yX�鞰dSb�'������3-B#i���pf�Ӥ@+��glȲ/��
t��U������:H����#�I$}rJ[5�b��e�π@�:�`��C�M�j���X�jú ���݆Ac�丏��>�CJ̄��XT���6У<,�OV�����(��)����n#&�AAO�0 �l@��%���� �D�2�q�/W)}���O��Ez�O��'h�E��gY {�ԝ�"A��b�.-s�&��ps�Ѓcn�OZ�D�O�$����?��O=-�f�)���C��ȍZY�uz��ř�x+V�zP�AN�CH�d��*~��
�����n�J�*Q.>B���A�U��x���V��~BL�\��9�$�?5G\LS3����y2��85��̐Ə�,`�<�MT ��'�`7m4�$F�YU*��OޛƄL�w��xA��Har0�Cc�7L��D�O4y���O��$d>98Dc^�;L���"� �l��q��>"�i�*�,�^Y��M��*�Y����(mp��y�L���Fl�D�!��@�!:n��񂍐r@��!��[�'%�i���?��O~����L p��Q���%6� �"��2lO��@�Y�P�bs��/ �
O��u��B�@���˒�Ь��h�rW��Ġ<��n]:�?ͧ�?�(���y�r]r����-�{6HX�%�,DI .��X�I�O�l�"��Ə7��{W�>/-
=R�nT/��@�O�����%�M^�2#�Rn�b�N<���?�
y	3](f�f\�� E7k"�0kY�9���Rf�[4k���Z�!U <Y���H=*-�'��#���?��IzӦ0�,H��R�O8J��)P�"O0Z�i��f��p�B)y�m��ρb����C&��Vx�@�ڝy��e'IA�Nޘ�
��'E��'�B�<ڌX�P�'�"�'4�;6@�)Z�o\�kA���VN�X.D�b��*C�A�f�i�&��Cj�V�b>	�P�Hal�&G�}
��×��#B��9�(��lI���v��L�t7�F).f<1���@�0�ƬH,�r �����O�t��=�Q���3�a0)O�A�����`��O��;�Hv(<R��]8A A8 $�oj��ȓV1�D*�,V*<P2���L����?�V�i>���t}*��G�^����*ot1�f�N	���ˁ,Q�-N���O��d�OZ�;�?)�����J�8�e^0Z��+�O��lP��bH(]7�1��H lO�u*���?�T�I5�+��h���ُ3p�"��rr<��	�/���Xkk5�<�&	W+WI�`9�h�O��.���'�d��!�5o�.�s�bˍ�	�'�x�&�()mf�8ֆ�v(��{��x�t�d�<�M�N��̦���M�,{"�1rÊj��a�Ԝ�?1�I�}����?��O@��S��[�^L�"ٔ0��i2���w}��*�ÛX� D�朻C �t�D�t�'G؈R7E��o�@i�!��kO:�ks�02����Gq�Q�+\$�>���Ra�'�.���?��O�&�/9,�%�f%��K�h�`�d�OH���҂u�.`�&k\"eARL�q��=á��\M��f �&GXZy���R4f"�xԤ�Of�-D�����|B���ߛ@�6m�xu���o֫-���I�l^�G�����؟�Z +R���IGk��Hb4���X2� q�D���,�\�gl��_h���넻��3�8(HMD�lt����X�f��-��wШ���'r!H�M��q�,�I�*�
q����x�$U�?9��h�6-I� ��#�$k2��aID�?[!�$�>C��9y�	ǑQ�}�����sSb�G{�O� �<��%�x���3��?a�v��4�;/R@6��O��D�O�\|�
�$�O����O��S:]��E'
L�E:q`�P N��=�4��F�Z���k,��T�3�Ӂ0
����';Y*�o��zq�"�)c��4ʵ����i��nڮ0Z.:��
9]U�'?�K�lD��y�(��*��l�y�nȀdƊi�B�&�Ԡd�Oq��'r�x�l��H���:@\���%�o�<q�i�:�x�D7Iϼz�$�g��w����x�C5$�Mce�P5_6m8��F=��p` '�,�d�O����O����O��Dw>E�c�I�n��3�@�*SԾ���uä|��#SB�(S�+Va�E)$ʄ�Y�Q���f.�� ��;���V�&�a+W s���2�ƻDn�i
�VՖ�$	Q�4 `l:w`W�55s�q �š.� 8;%G4{l�U�2'�O8�$$���'!2��0C?N�R�[w�X����
���S�? �$C�еv��\�Tn��^��S����Ц��ITyb�4.Ɇ�'�M�ꗑ���wm�.>"��!�#ȍ�R�'c$Ȉ3�'*�>�R�@���(]^��d��+���F�@�E.r�"%f�Q��5�&�/[m֜X��1�(O ��A�v�AtK�2`
�t�P
�Հ�'�G邱q���)q~�����(OPe��'�_��X��cr*[�DF�p9��;�K4��|؞�pjW�),��G+�2�p��ì0��ò��#NaV���܊rL�����%*�(8��My�8��6��O��D�|ZbK��M�B��Nf)��oM�&f�iɣ��(���'�Xx	!���
�X��3)҉�~*���'*hl�[��qv��R��	Z��$����#ԁ~v�*B�ĵDg���
s�'9N>��N@@�V`D���0z�H$���H�O�	%�b?	b�H�� �(��u^n�90�:D��֪�IT��c�'��M�H\AQ�7OجFyҏ�H/��{���∓�J��4l�؟T�I̟�c��,<D��IɟD�I���V�dYp�_<;5�)%�܊�.0Yh5�(}�P�S�CC�� 2.�H�'q-=i��f�`�`�;SFR��(zTF5Bk�u,f(:���|��(�V�U� ��XO~���Y:��.+�4�y7�ґLk~���A�vj"*J>��ٟ�>O,S��N}������b�� F"O8��ɾu/�!aD&@<j�^-��>�5�i>�'��8s�Z8[v��(ň)m�$�j��=0����?���?1�_w��O��dh>)
g#�+Y��Q�0���a��;��Յ�$J�ej T�-C�	���+k3Q���խ�v�LI��$ 6!Җ-�CƁX�laː�K.B�Z��XP���ͷXd���!��lIm!888�e�*4H찑�'I�����D�l9�IJ�0~�p���!���>����ׅ�\)���4%qOP�mZw�7F/Z��۴�?Q�4?��TAp"�(��*u8�h�3�'�r+�3"�'�����b����"QWع�/Aܴ�ʑ愱^=$�YI�2uSa��_ɰtp�j:ʓ�~e�����!���Z�G1l� p�����Z!�T�RK�(5ء�栎�+Rȩ��D&ʓmJdL�	��	�c>m��/A=��yqf �}}�C�y�r�j�W#*���Á�G��C�I�9�:��A�\�G��JU�\0�)`�CY�$$�	hݴ�?�����6|�6�Ӊ
̒�
W�J�6f6t�0�lF:��I�4R��N���e�:�@�2T�>����gBW�� � �L��"��&ΎE�	Ε�ē%"D��$	ׇm��ä�
\N%I3��,|���')����Vn³��8�e�V�]Ѹ9%��Qv�O�<'�b?!�ӅA�{�E�����6���E�(D�<�! M��X���מ¤�0F9O�DyR�ΑU��ԡ��K�$���JעJ2��m�۟�������橜�-���I՟���������c.a�a>a_r������P�4�[�(zBY*��I�A���i�O�~�'s� A��OB���OZ�0���d�);��<x� ���4q��7J,A��K�
��>Ũ�b͛�y�"1J�-S�nҒL�<P襩�0,\'�Lȥi�Oq��'UnUYd+�&\P�r$�ɻY�V\
�'nܴzN_�%��2.�`2x�N�,���4�pO��XciŴq�����~.`%�B&���Ɯ�$� �H�I蟨��6�u��'X<����r%�; %xy�4�Ï| ���@S )G�s�D�m��L����
&{���1#� �(O�����é/��!�e��K�LE8K�Oxꐊ���~x��7+X)Ǝ��ǀò?�p��>����� Ӥk����:h�����{��`�I�p?ib-�2=�H 3�X� �����Ak�<��@I}����hGj�< ���^���|2�ʙL"�7M�Ol6�_�&P�bV�V�33�L���q����'�RkB-"XR�'��i�m�&�Q�˂q��I�%��h�+B0mM:�J��'C�����V���;�ꃧ|��d �C�.U�hcw��%F���i�I bUl�CACEj�'�$1���n��!"-�@��tq��0���
��`Э[)�h��[�`�2\�voW1~�2�h@ň�y�� 	7�Ε��1.�@H'�i�R�'E�S�+�@o�a(�P��i��y��B�i?n�K��?�쌄�n�P��5B}�!Qҥ�Z��|�`���鞦lƶ�3��X��n�Ys�Ƿ�'j6m����SV�f�,_�ִbU�E�,���r�O�|�g�	O�Tk2�.�0�1�IC�I"
\��d_W�)�S�䒭01��%�^�����*�C�I�+m��LB<b���@
t���4��XGyR� 0d��� y�z�#
:3dl�ğH�	ݟ(��
.6�8L����t��֟�.:*�mc��b��p���=o�"ң`�.���m{~���u�Kz̧L~"I�-�O�m+�k�e�������.�F�z���Q�,)���N�Bd����-3�pm�%M���IC�'��ϻ!P΅)��3DV�Q�ͽ{�9��>�dͼ{���L<!��фd��й����t���Fp�<��L6v�@<;P+Cs6��Q�\l?)�%摞��M�)� �1�U:
*`�8�� h��"3��u	ê�͟��	ßh�I��u��'��6�B S��¥cn�̚F��0�*����M�C��PJ`ŤC���BQLO�E��2��¾�(O�P�N��nR�+�4m�̍�0�۰m���!�ĳ;���ҷ+Q402f�EH�����@�%����SX�c)ȁ*�v�����M�v��O�Q��	�F�>UNU6w+`�Ç����c!�O�O�`�:"�v��c*L�4�T9R�D��Q%����ʦ	�O�ԐC��`G���+7A��:���&�'���Q?�T�aqŗ|�"��ȓZ{��`�Kj)�CO�F2��ȓ'3
���v}�5���ם�$�ȓ<U> �D��4�̑sa��6�ȓ���ȍbg0%�e;X�bE��>l��c��D�>	���#���j|��w8����-�c�,s�maR��ȓ"J��P���]�|!Q��!����> F��r�I	�#ؠS`~X�ȓG#͢c��8l��h��p:���@�f����h�j|HR��%96��>�^uYq	�	��9�0m��:���K@H`��/K�0���:^줵��-?��c�d�<0�h���;,�u�ȓ��ݸ2��J���/�4x����t-3GJ�(W˾�Z0��&��ȓ�"U#���~VY�&��'*Ϟ\��Op�h�����H��B�#}�Z��ȓV�XH�GIXl�da�a"2\}��6��=x���t��K�Ȓ`���ȓ ���#��< Lҝ��̚Tf���ȓ���BM=h\h�(�J�R�tɇȓX�@-�uO$I�2��%��.E
��ȓI�H����/@s�]���ˤ_�>���.00�
[QRћr+�"vs��ȓf��Yk@-&�yS�hX�y¤�ȓnt�����Mo���0�S?����ȓ0�>�qA��I�F�T�T��ȓ�z�sc��?+�m��N`�>)��IE
h�GۨFC�Ű�)�>pL�e�ȓ��Y3H�'6Z��� _>�>��ȓ~�b�!W)��I�F��,��:�����B.E�G,�?��Ũ�Ɨ�[����ȓb�v�h��O;8b�VM��TȒ��ȓi�*!��*��4;�*R�\�J��ȓ����e�����j�	K�e�b��ȓO�:��6�N''���B�OY#d�쁆�H>���֮2� U�n�u{d�ȓ���ڔ%��/ ��4�ΗV�5�ȓDʴD�)�ƨ������ȓe�"���E�{J��M��攅�,X�Jq��'|���Y��ӡ�4���1p��e�����'W#h�Z������Ä}�P�m�� �z��j\}C��
0�h�'%����d��3v(�͘�l&t�������V�<i�aK*� ��B>��۠��I�<��f��]x����ѽ�q;թ�m�<�C�P�#��@��W9~�~3�� j�<�Q�[�����������Nn�<��a���p�G��&r0��U!@�<7�,N����2Ժq�`�+�,�D�<�w�T�@�*$J�ϳ �X �%fHA�<�2�ĐO&����Z7c����/��<��J�c,�h�Rׇ4y2����T�<9�S�U�6�!�ʒ�����LR�<A�n�?<��	�5JY�j�E p�IM�<� �!�0�˃X�<����NX�1t"O�H�b��<_��(a�CP� t�ܱV"O�t���R	J��Л�(X4P6I�E"Or CB�-\V
['J�6خ$+R"O�<!�W�q����d�����"O��y��.�� �m �L�8"�"ON��f���}Ȗ��m�K����E"Ol�`5hN� *��l�h�ā�6"On0�b٣/3����>Iw� �"O�ة6�� �^�h�$޴aș�p"O���-vB���ʐ9[D�a�%"Ot���@L�_�L�T�ņ?`��r"O.�8��۟c�.�f�/A�F�� "O�L�l>CJ]��Ɋ3~Vy2"O���%d�!<���e�,?�rm�"Ó��&�3<ifqA�:[XD��"O�!�"�����E�n�C5"OF���,�n�����Y�@��
w"O8\"Ȝ/�8���*ϐ���"O`�i���%OT���ț�{���9�"O��A��U�FQ���[p
L+�"O"�r5U�GctE(����iX�R�"O88pl�#pR�J�LM�'�JQ�"O$��D�Vx
�EW-�b}*"O^Y)&(�/D�`W%ϦM��3�"O2t;3&��X{rd�N�:�:4�A"O��؁��y�I�bM7,�*�� "O����VЬ��]�2�*�"O�e�㣎��f5Crő]q�-�V"O\���Ҿ1������,
I,8��"O�m
��:u*>$�c�
7&.�t;�"O��W�
�W������̧r'���"O
`bt��[����*5��"O& �'�#|a6� �m��E`�"O�hzS*Kߢ���k�x(�"O�e�P��&���IfJ�G.�ʰ"O^E�F�H�~���Xhӛk�t%C"Oe�@CݖH�̫�'Ė*:&؈"OrQ�/U�,�(d�2L	�B�"O|�7P�gy$�f��r^��k"OrXj��
�>h�AA �[�� "OK�.�����M)P\��93`\�y�e�ͳcͨB嶤���;�y�	P"l�5��p
x}����y��� @S���{��E��A��y�Ѧ(���p@]6_ޘ9I�d��yB�J����a Є&�dBf �yb$�vq��p�<\��D�yb G�7#��e^73Rtk�T�y�R�8ҦxK�o�R���jBo��y�Ɗ@�Რf̎M��4E��yrBɼ.I(�"E�-��!lA��y�e�#m�R���ѳF�lΊ�y����F5
�D��F�Z0�F�y�DΖ�QӇ��R��s��;�y(�UY�w�:KѠp��Q��y�I��s@F	{�&B��!�#�y��]�X�0��h׎'��Y�7��:�y 4G���Y��Lmpᷡ���y����F)�e��V5J��)���y�L܏E�A �^�D�u׀>�ybB^*��,Y�ʞ�5%� [n	��y$�.U�ԸK���*0��('��y����G^�� ���p��tr��)�y
� 6M�r�8a���*g�L��hC"O$<�e�.2f� D�^I�6"OzQhQR<C�e*�	�X����"O�3�j¬"�vl�ʁi����"O�| ��[�T��� m-~XI"OB�ra��4A��8��D�:�R���"O�)�T'D�+;������|�UB1"O��c]��B��D�D'Id�!;�"O0A�7dM8r�����cɕ*P|�3�"O�Yj�
�qIN�a��@?0n���"O�M�w阜$���RW�	�2m�A�f"OL)����Fʠ�fľU�)r"O�r��uw����EI�@D��a"O8��+�-��Q�s�K�/��R"O�l��&�Q�`�Z��
2��0 �"O�ՠ�  ��$��舕r��9�"O�<"�ێuC�X0��H3w�x��"Oȱ3U��](���K@ܪ"OrG&G-4�x`#�e�U��\r�"Ot��GGɲFL1�<�<�`"O~A褮�4Z�49k�l�)��шC"O��c��A�,a U�K X�0�w"O�铅C�fl4�5dZ2	Ćp��"OV� �DKY�D��SD�J��A�7"O^u�pn��@��P���R�&��E"O�AmŊH0���s �r�2y9@"O����>4�KBL#b��,�"O���l�?C�� �N��e���"O����	>��)�3.��xM>ɰ�"O�ac�X�O�rГd��oFdp�2"O�-����G��i��E 
ۚ1"O�lZ�^�,,4�ӏ�5��hٓ"O�i�Eʫ�x j����I \@I�"O���a�ԨW�F��$�i�"OL�YRΉ 5��2bX�uy��8�"O�9�fL�7 �j|��͹
�Bv"OU�KwH@��@�	J��� "O܍����&<G��)���~�Z	�%"Oܙ�"ȕ�o�0�iO���85��"OQ�v�\��\L��$A�O݆q��"O�5��E?[@D3u��R��V"O�X���]�����Ċ�>�0��"OH�x���9���@� 
}��]ɓ"O�!C��B<U��d�⯊��P�q"O�с��H���"�9�"(��"O��
6�	{�,�i�L�#���Rq"O��oƅoC�mb�F�f��#�"O�xK�E$
Ȟę"E�"~�!"O@��3�"<�#5�m���"O�h�5�V�P��5HH#l�ʳ"O��J�
ŴPR�'�\�g��s�"OJ��w�Ū7,X=�u�;d��"O��15��J��A�a`P�DT�0��"O�$��,Кs�"������"OH$yס�h�Ȑ��0@��2�"Ozԫ%�!D,�}�l��JϤ"O䝰�\�c8�PbNӭ;%�Q2�"O�]���N��xz��E�%����"O���rHU�p����aӇGPPy@"O����
](�A�u B����"O���e��R�ŃT�L26��r"O| ��cU;HD�:5NP�qf����"O�q��P,v�ԩ��H�T���e"O ��	��=��-kgMD%!�􄙂"O� ���C�ۓ]!ؐ�#��fԞ�0v"O��Q�a����)�� Z>܂�"Or���cԙ;U�x��ɑ�+U�ia�"Ov��u�U�ws �Ւ��@�d"O����	^��;f�4I��U{""O��i������~�T�*�"O�z�]2$i橀�E˪:m���"O��Pk/MV���%�?	 ��"O�S�MM�~�aFg���X�"O�u�0��8���#Rl�*�h�"O�pl˗p�PBv	[84��"O^| �jG9a|e���A��q�'�m�C��`*��ƛ/��-�d"T7$Z�[�A�<3:�8d�#D���'��";¼��h��%d�G D����J��&
b��#�D�Qy(L#�$9D�l*UǞ�A�Tk�朑.J�c�+D��r���Kx�!����4Tʒ���c,D��xԧܸ;v%bve�ax��'=D����������a��1�d�x�7D�� 㨒�O��P����zX�uP.1D��kc�D6=䄵:q=Z�՘f�,D�T#��#~���a��ZgǦ��G�)D��S1AL�G-|ɛ���_&T��b(D�0�˔�8J��[%z�2�`3�9D���a�E�M�"$��Rvp��&D��¢e�d1r6!�~�n���O9D��A��A�2A��6!:XH%D��"Ҁա\��	����6h�d��J!D���C韗�Ta�QC��Pl$[�#D�P�k��cl�9�VB�4OD�(bQ("D�p 0@�� ��ZA�\��YŎ!D������"1� �$�I�-��P��+D�h6��	�!�H�-q���P�)D�!eG�����d�P��sXB�I�)CBP�bmW�\	��� fՠb��C�I7E� ����X3
��V�*<I�C�ImZ�a�Q�2d�ȳ�ߚ�B�I�F� 4j�#>���wl �S��C�IuZ�;P�W���j2��<4��C��4~ �U G
9�47ƚ�;6�ȓB:4x[�O��$���5n�����F�D��6c�#?����$W��*0��O�(��Ƌ/��@R��MBJ���� ����6��Q�J�C��ńȓ[~Nq�G p$�r��ޑ�ȓs)2��p'� `���+�Q�z���ȓ]�~ ��ޠL���sw#ښ_R��ȓ�ԭ�f��d����I�0�ȓA�5��$��صÆ�۷2� ���4$�rv ��������P��XF0i��εH�1�Ć&D�B�/-Q����;k��Q"�ߥUDC�Ɂ�>X1ɜ�GZ�)���\	
ҲB�	�0�4�c���Kچ=`� \�C�B䉳wx�����+}�rx�o_�(��B�I�O�Ȫ�&_f���sW��`�B�ɁFl�"&B��"|²E��WǐB�I�n�h1ڇ���=�L�t�P�~C�I,]���!b�>Ud� 9g��7O��C�ɖ	Fs'�� a�h�4A� df4B��!uB�;�Y
tM<!�D��$2:B�Zer=��
� uj����B䉳H�^�#q�.�a�E-̞u��B䉾0�*���` j��(���էkXC�)� �H�-������S���I�"OؼR�^9�pB�Ch��"OԴ��A@`.=�$k�W�ܘ�p"O�Hp�č��:�y�
?���%"O u��؛y �"J�-S`@��"O&D��j��b���*w��7n��HK"O��j�܁A2Np�1�\��u�"O2�s �-"^�%�H��5��"O,�s�ūs/R5�d+�>-a4p:2"OJ��ń�,=L!�K�Q��$*�"O�hH@�H.t�4=*�鎝-�	�"OjP§)�X3�Hh�'��J]�G"O� ��J� /*�0�S�dr��(F"O��)��D�4�l@hA�˴�a�"O �1�g||4�� ̦[�0���"Oi�R�FF� 5kf@��F��tb�"Od}�w?
��ˣf��F�`"O���F�
g��L�K�T*g"Ox ��@X��U@&CI%8���"O�����y �	��@Ͼ��m"O���B��J�Y���
��"O<�`�A�2P}8�RTņ�9��"O�'I3;Q�0I�D�6��"OvU����9�LY��^29�(�b"OƉz� �Ĉ�a�	����u"O,���:��p��
M�K���!�"O��:��T"Y���ٴ	M��0}HQ"OV�ɗ��Y�l�	�h�+�D"O��@�ڷT�U��%O�QB����"O���'�9]���7B�4 �h�"O�8�F쎷T�p��G�7W~��"O��!�Ά���R@�gb�@��"O��ؓ*��bRЛ�ACU��""O� 8�#�RA��Z�4 �"O$]�Q.�#�Уg#�,l����'"O��7O�+b�M&��$�X�3"O6�+s��\.Q�d�P%Q�ԱX�"O���D�o�R��1)֌�ZYH�"O1;��Ǹ`"�AT���Sքr�"O|�6�8"Qb(`�k����92"O�xZ�(�h����ϋR~~1k�"O<��u��5gA�9�CDLW� u"O��j�T�|}P�

�V��qP�"O^�˶JX�e����F���It�pq�"O���U���_���Ɛgt\@�"O����W<9��
D�\�30��"O0�5 	0��Te4>yz��"O4�A��]�0�����E�to� �"O&��u���	`(pF�Q�T<�%"OT�4G�9/вl�C�B2U����"O*$�c��q�
y·
]���+F"OҸ���7@�.A�FK@�3F���"OP���B\�s��86��A�]A�"O`�Ҁ�R<	"E��n^(:�JL�"O�pR�M���S��RN��Z�"Ox���ؾ	�|- �d��Z����r"OzX���! �����f�xyp�"O i�a��B�Zp�u���ص� "O��G�N�rV|H��%�(?f Q"O^l�Ʃp�&H�ӄ��JB`���"O���>�`��3)�)��Z�"O�X�TiĀ,�V��)����a*�"OrT�R%P?7�H���"m�ptH5"O�mp�&�
L���'�3d��H��"O� ���7� &
�i��C8�,I�"O���v�; Z�a��Gԟ5Hz��"O5��j	<P�9y�h	�"Oܕ��A����u蚩~٨���"O�|�Mf}�Ġ%�Md�V��1"O@XY��XCk��`�T�q朁 "O��`���'_�h����2W�BP��"O&�[7��-A삄Kgؿ_����"O��dL|0�H+f��p��"O��@U�M�c��4��� �585"O>L�th@�s����K�3y��Y�"O���Pnא\ltA �#L^|`��"O)#���J�~t*t�	�T����"O`�����zS��Y� FV���c4"O�PIХ�7ڭ0���X���t"Oȍq�n�~���c�!�����"O��"P@)t�$ɳ�B�-��-�$"O�ld�в|,��Zp�@�B6���"Ol���Qp�6ဃ&�)�"O`�5�_��8��V߂h�W"O�}u�ڌ6�\08 $�0U���3�"O\�z%�(&��습
�6z�V�;"O�iR�j�l!"ѐ�jҗz��Х"O(�7��J6�arHF<M�Liz"O<�#E�D� +��۸@& �ۥ"O>H�"�' "t`K�bFNu�lI "O�s����c d�$��D���yg"O��9�mb��T�_-�
�2A"On��D��@��b��S�R�<���"O�ŧX����G�:Ɔݚ�"O*��]WJ�BW�+'����"O��R�f��sF���J�W��Y�B"O���@K��rl���.dޜC�"O�E�Wh�|��U���C0�Ȃ�"O����#�!T�����)`�*�"OF(�1�R�q� ՠ���P$��"O�k�G��Z}�a�rH�@�"OHP�Wlݮ?�`i�@ì�""ON�S���W� 8)�m�3� �U"O��3� ���!ҌA�^Lx�"O$��W�Z��	 ��M�\=�"OP��vd�V��б�n�u��9�"O�u��b�v<��w���a��X#"O�M��N��^L��TW��v`��"O@�(�8��kC�2�4�3"O��*0���f"�����%�@ZE"O(`��]��1f���1��`�"O�ݰ1*��C������ñ_��t`"O��sA*L�*�6�s,�H���"O=��a�~DV����Ξ>&�P�e"O�TGÛ�f�BR�Z<5��"O�pZ#	�$?L@���%dv���"O�Y���э����!�T�@B"O�hK���3 pu ��IA�μ�"O���	@)Fv�x�˄e�f��7"Ov�rHN:���*�<�M3�"O�aF�PظI���!��$��"O� �'�Y���@c��&vv-��"O�����
ah�$���*f� *�"O"�2��� O��Xa�Ѕ2���"Ox)���$&�����m�zdq`"OR�yE�B����6�
��,q�"O�P����TD�4!I�r9�p�"ON5�w���m�C���c2�q�R"O� 4�b@o�>(İ�a�O�%<0ɩ�"O�xJcA^�z��K�%�>H�l��"O�a�/#�\�3�d8Z�L��@"OP� #��$t��۴��[����"O��+�"�+V+���2�9D� \K�"Of���+�n��D�Aܸ�ΙT"O ����}:*��Ƌײ8��@�4"OJ�p`�S��p�SLMz���7"O�$p��T�d���&�qՈU�w"O(q�Ê"�l�D�+�=�"Ol��0H�<�&����ձlP�)p"O@�M�#"��!T�$)�D���"O�8��oZF��D�'��9�`�"OL���S�Y] �2fý+���"O�� �.B�Js��"��O�JI��"OZ�An�LN[n֫����'�ց���4_�z,j��MpD�[�CW(J�"W̖1ID�4�ȓ|H%�7�Ėo6Y��M�Pxل�.�FY��"��[:�bR��&"�D,��#~���%�4j��� b���j���!�S�N�N���i�A�p�2ل�;�@9��ɹf��0��=���ȓ ,xR�VHZ�QjC�,�̇�M�*m1��B�<BH23k�,����ʓ ��b'#_�sAB�%�*V_�C�I3<䨰2eLD�ʼ���=U�C�I�9�`9�aD?
P�bCZ��C�	60�v5�!�>�`�
A�Y ��C�	���\c7l�0
����b�
rXB�I�Yֽq�KU�b��2b�^B�I,J4��u�G'��(C�R�B�	�6�^P��	WR�tAa�C�B�	N�"�:��L�����ρl B�	�p�#3Ȃ�T�D�ңc%j�C䉌p���4�[�'��(�J����B�	0�0�RVH�-������>	�B�+1,�PA@+�[32��G�{	�C��+�xkd�K>I�B���$]��rC�	a�:캃�߰DD�2��i�\C䉫:�^E�R�ӯAM�|#7�DI,C�ɀ\�A)�ٜvRV8S��X?[nC�ɔx��}2��M�g�-(*̉Y�LB�I1]ņ��'
�d�����VR�B�ɶP������HI�Ӧ�G�OB�I�L��F&�f~訉ՈC1yҔB��.<��RE��A=���2+�-�8B�I$VJ��!���Q	��醵6�NC�	�bx&$�ʖ8�ȠjTǤQ�B�I=iz �u��|��hK�JC�`B�I6y���s�U��
eH���!btTB�IS�ށ��	L[��de�A�RB䉺7��e����j��k�NF;Y�TC�Ij�(���zLL��Q!ʮd�vB䉊w�X�I#�M�%�F�{a�+�JB�	�2G��f&�9
�xe�4��.�*B�	CJ���ٙ:ܰx��-{�B䉖i����P�
Y���r�7;ZB��ipT4��	�+g���� ���L.B��A^�P�@��.�v�x6h� 	[ B�!Z3,�4*�.B�>����
{��C�	�j����'�h#�@U�V��C�	� �|���nשs���Q$/��C䉟4��9�)܍��!����I�C�I#&����H<��)J�����C�)� T�s$-�+�.\h�K�o���"�*OJ)BR���8:���u	�'(HAP�n�溈Iau����'��AC�䈅�,��nJ-��'`!�1��7�� [rH����J D�����зKTV䣖�ڋ{LI��<D�Hh�J�
���#�
W�3t*!�7$/D���s�2��I�J'Pi�����yA]�I�h���%E��Q�t+P��y2l8<�\a��GV�B-�h1���y�k��;C1�`� Ak�$o��yr+L�h��08��:8���TF�yr�ݛG#<tzqB؎Z�*�3 ۋ�y�m�&^ڍ�3a�<D^�T��S0�y��J2x[:���K�Q�6l����y�@@�[�zA0A`ق~r��d�ѫ�y�!X �H*W�B3���;�y�H�Tǐ1
����kr�Q�L��y�iX/e��p!�eR1�r�{�'&�i��<j�RT��N�A����'�`�(�"��N�|�Uiڞ	P�Q�'� �r����A�5C��\�Nx(�'�N-����[Ж�qw�� /v,z�'����?	��q�+� �l�
�'F�48 a�&6�����r�
	�
�'v��Ui˳��)�Ĕ
���r
�'��(��`�n���J�:c{�X
�'5q�S�C�E�	AU�8\�	�'L �eD63f*�#^���@�'(ejr�K�H���c�˭A����'��Xr�-�]��`�BU�w�V��'BD�X2�J����嘨g�����'
�fG�%�QI�W�����'+d�ⓦ��&)��J��<��:�'�hǥѮA8Fŋ� �wa��'1���ǪE�����D*��(�c�',�Q��
Y�Pl`�iٵ.�թ�'&P钵��3F�PK5��LP"�'J��� Ŗ$c�
����ޞh��'�Q�C���i��\�4mч|��d�'.D�@��Ǔ l�	��%ȺmΪq�'�r�á��B�d���.k�
���'R�8�����n[���'~RXx�k�I�҄�L̨M-���'Dv p1�H_^�Y��E�3��4y�'�ȴK�ⅥV����G��#��H)	�'E��pG�G�V�&��ꔺ�D�@�'`�PCgJD"o���f�������'!tp	&C�	X�lPQ���,C���2�'���I���8���2��qL�P
�'ӎ�z�_�+
�X�B/Wno<���'�B5UN�w�}P�5Y����'�)���>���FCگc�9�
�'��E�A&�8���x��Q	YԔ 
�'�C�H�3T�&t�B�Oc���	�'���1!�] z��d�R�}l���'�L��5�� E븍��$w(D���'�"8�'�2;-Z���aH=rKv���'��|�ф,M'f�x�D�h8z���'܂TCt,Kr B֋^"1zT���'S���Qm��ip�x+���+�4��'X���MM�|�; K��[3T�'�0�G
"Ft�!�-#��$	�'k]C��ȅQ � z��5���(��� L��� �utإ!w�O�x���"O0	�.�:b�@Ɇ�M��Z%  "O
��nϿ6f�M(�DE�H�X�"O���-L-Zi�ij`��(x�~$�"O�0�1��$@���V�%��"Ofp�aK�r�^��F�Vl���"O�l2h�L60p
�DI?7L�lhr"O8pzsB	_����U�E�i	u"O�-�����[Z��7dIE>�p��"Ol�Aadި7� �X��>-�$� "OL-j҂��X��$�B�u�A "O|q�7�F
"��رj(Jܐ�"O�3�L!&l�,� ��0"O�qBeGڱ@X���t�� �l\ӥ"O�<�r-�'�:)s�MQ� ň|�d"On���ьպ%kC�U�ڰ��"Oyx��ťo�*,����
jH��7"O<X@���*3|�k�� Dk�u�"O��a+P�8�8{�I�!j�Dx�"OP%�d�P0dd���G� 6dE"O����� ��	��Ξg+�왆"O�� F5<�
$�c��}��"O6�ʔ/4L'hũ�� �;�Z��@"Op���\���a��1i��D�"O���OD9\��ۄ��1!2z<PT"O�ĀP�C�P�Ӊ�]	j�hҘ>	
�u�HM��b��b����Հm+��ȓj=<,Z$��*L����a�#4?�=�ȓ	)�� �!x����1�̥8VR��ȓB� �6�T	.�yBCo�#~	 ���+���ɀ�߾�δcu % iq��A�sB�R�Ny����6����H�(�SP�mJ��Ԃ^8^�PԄ�n��+�F�9�ޑ�3��%�D��ȓ�ąX6�޼@B:�h��i�z!��u)֙�`菸)���B�� i�ք�ȓo�4BR[I+���P��! 7dI�ȓ>P,���� ����� `BЄȓ1^r�rb�3���ƩНT%P�ȓ;윀�&E�2�������:��T�ȓU�>0Y3f�^\L4"�L�P�ȓf�{�Ek��*��HǬ��I��ĨB^ʔ����3�����N�!���G!�|D��7��مȓ/�~D�c@0hY��"����A�D�ȓ\��a��8�\mZ���$y�ȓr � �B@H�$�bL�N܆Ʌȓ#�Ɯ��3t:�Ձ��ށ7�	���xyǐ<wK|a��EI%T5���ȓ&@���&^6�jаV�ܫc72̇�>6x}�֨�5/X��'#�@���X]�w���W����.KFȈ�ʓp�t�v��5 %��fj vvC�Ɉ{Gh�`��X�]��]����BC�	?i����F�o]`�j��L,9h$C�I�vZ�%�fEI�Hɒ0See�wʤC�I�5�~=��$^���`��ה*��C�ɋ(��|�Â�&}b��5�6��C䉶V���0Hۦ||B$;E!X�5jpC�	�d�LX� ��+dH[��
:#�B�	�h���$�эVpХKw��-U B�	�i��@¥��p�}��T�c�C�	�\\t0�#.\(�٢�W��C��#��8S�>�J=�!�W�(�C�)� F`���:pAb���K�v��B"O��cC`
9*"�
��&<���3*OVe*�.�R�"�2W��y�!(�'v��b�f�6�к&�H`��x��'
��рn	�Gmȕ���%fv��'�F(xAiB=hz�ɥ��H.�9
�'��`�5�H�pt\�pŉ�2X�'�I�J	�|�^$R�iɺD
�j�'���3��Y��p��8.�ݰ
�'50��cY<6�<��P��,9��
�'xZ�aro�4J��Tڗ%U�;�X�A	�'�����e�^%���B]Fݱ�'v�%�7,	�zSژ���/�U��'q�0V��u+�mfF-+p~)z�'�h�c�G@�}$H�mUcT��
�'6�4ʦ.��C���ƈH�!x
�'h��q�OċR8����?�f���'�f���� �!z5�u�Q<1�&��'~Zȃ��̈́.�6@i�n��!�0x��'�.� ���wӬ$P�H6�H��'�4�Q��Mo\��'H�@����'��Գ����Tr�����[}F�q�'�ݑa]C�
x)��D)4�
�'��F-kt����"�  @�'�t�4j�>I��5kgE7|�r��'���&<S@H`��ϐxJJ�[�'u���!�Q�5$ٲQfW�jk�;�'�=A�(Q�1��3V7_��<��'�����:7�hp���a4H���'��A�*��:M9U�ٝU!����'���򁞕+��zdeN┠��'��4���$`��,��c��F�x�:�'#֠�mW�]��8у�K�=�(��'mf�� cB�B��$J79,����'�Q:��(	O�� �c�(3�|a
	�'��8��d[~f����.�:\��'kr�У�.��Ei3�K�,����'A �d|�S���66���'6�����F�LMࢌ���,!j�'8 �0ӥ��2Y̒2�J�=M�	��'mV��@�*O��[�e����b�'�h���oD+$�$hRCN�|:�:	�'0�+�f�"Y���A`�]
2���'�`m�d�f�B�%����#�'�vx �cM�E�P�[��}��Er�'�zlb'��|��t @�{�����'�Nu�'��#(�Y�CJ[+m�� �'w� B���F�xcaS*a��|Q�'�И`��JLPB����!`�1�yR͟fR�s����E:T!�!��y҃�$�0xxCa�*�8��5*4�yR���+���*�V�dN	�y����f�VssɆ?(Vȝ8���y2"�0�����Т�ѦE��yRa:"�N�q!�S�/�8����y���?=�yY�H�(`엕�yb�� tmHT$��,�D=�H���y��B"_i�[��B88 9FF�4�yb��4-�4�a%�~xZ�!M��yҠ��n~�	F.
� ���h&���y��Ȑh�FE��K=v��HR��<�y��L�_oDM9��J�m`.�#��%�y� E�nԪ���ϔ�kΖ����yr�Y�
#L0��	�4/@�4�%җ�y
� ���7h�m�0q��M[1ZV��"O�e�MF;g\$Cu,дa�F�C"O������(�V�Aa�C���Q"O.���(U;!"�h ��i�n��!"O&���{�$�)G)[��q"O��xD-G�k�,Uɥ��+P��	�"O,ő&��Ve@�Gѷ��D"Ol�#�G��v0���sI��-�\��"Ode���!{S�!��0��ӕ�y���~��EǬ�*�1�R���yRQ�H��l'c�9��M��y2�ҭm��[
@ O�h"����y2$ʆw�)µf�	���"�B���y⯕�N����'�4��a7�8�y�K	w��bWl	�{7��Qp��ygQ([G,��Ɓt��$��Ǌ�y�MS�m�t�7akn\�j�F�&�y2 Ը]�|Y�e�f�1�`��y��o����dMY>���ɕ��y�K@�&^�t��n�)�݁w��7�y��̺B�|�����1�ݹFa��y�w�t� ��ќ|
x�F���yr�P;��c͘.{�>�H!�B��yr㜧8`��H��{-℡@#S$�y�	�8^[hyB��q>�Yeޕ�yr�NpO�(:3�_%aA`��*�y2eҢ!W6�!#k]�M�>�	C��0�y",D(bX���E��ӏʉ�y���u{���ï>
Ő=�dF�yB�U��LT;��E�	��rtM���y��ɸ�b�2�%� ���G�%�y�D�hi�xcdo�	�$��'���y�m~'����\�gLb����yr�b��$��4t���#���O#~*d��K�v@��]�p	A�c�|�<��脚D"iq!�&W��prACw~¯,�S�O�$@���'�Y3ϋ�$�(��'h�(�퓟%T�����+0�l҉{R�'�����cH-45��y �Ĝ1�\`�'`�z4)��(<��gƘWCʽ{�'	�e0�z��t��ΛHE���'a*<��ː0�
�I׫O>B�R���'k��h�Ĥlrf�z6��9�l�"�'v|���E�o�<��%	%��`c�'�x�1bO7�(�a���$�p�'~�Qa�+�,�d0���f�J�'ph8p�FW� @i`�k�D %)	�'KN���M>$��H��y�����'�@t�ɕ��ś�N�x�X0�'��ܻW��&��=�P5o�h�'U���gB����ȶ�Vfr���'!6�Z��<��Ʀ�u����'�8����{ܺ�[�"W�a�Hu�'�V�Z�-���� ��f�4a�����'#�i�WM�?#Ր���Ǔ�D���'"D10fD�>���R���;H*�*�'�� #d�);��0K�8r��a�'��R�G4b4���j�7��|�<)$'��.-�P���i���ha^v�<閎�$C쀓�mصip<����W�<qs��u&ȼ@��2��$(S�Y�<!�k^'�	��l�
�\!RD�Q�<9�n��K�:�s���N�����L\M�<��M[�
��4�$$EC�����"I�<� �q���
_����U��'B���"OV�CI��ݘI�@��#O-y2�"O:q�"/�"��;`Á�Mν�a�'���H�'�v��nR��0i��l��Rʐ�s�'P�=0���:c)&�� O�"��h��Ą�!�pE�D��G��`�O�
[`e����y"B��]Д4ɒg�=n�Q�J"�~� �� c��}j NQ�Ah�H�"���l��P^�<is�A�*��&�vBV���DFR~�!�+�N<���39���'�\���T�d]l��č1�M;SƓ�/���RC
�0;4���!l��X>B�I�V8 �˄iL��p1c~>L">�s�N�[t]!S�"�S$gkp@ql � B��#oϝPC0B�I�#t�H�F�ڷS#Mj7 б+S�����ۤ\ZɧH��R2�\��:��� �	�qb�"O`S��D�5e���3��4
��c�>b`���	�N�zyc�ل�f�Z$&�	Y�\q���3�y���q���*F'�V� �@�kA1�y�I-X���qAA�+9��ɷ�H<��Ox�V퓱B����隒}ժ��"/����C�I+|�ЀW H��Zi #ݡ6��əRj���?E��A�N��RH�YLi�Oղ�y���]��)��M�e'�|1�N��y� ��k�o��] �$���y�n���DЈs�۳� �7B��yrI�����ח4BɎ��y"NA�Hh�u��q�������yb�H�9�I�Wa
^F�C����y��7Ӱ��R�WX���q�Ͷ�yb#~����� �Tr�H�7�Pyb��-}.Q�Ԣ�YFn��D�{�<	�L�y[�h���&G8�"�Kw�<�����Ybd�ZVh6�z0Þr�<��n�5|��a ±t��4�e�Rc�<���+m܈I��j܇	؜�&�k�<1��P7Q��}�K�T/�`� �P�<�s�؟SL���a��;y�壅
�N�<����:G�Ba�Ï��2��Je(J�<��Ȍv���5$X#�	�SL�L�<�j�An�:`�|�\���c�<��;?��T%�$N~"x����^�<�#�Ĩ�$��cn�T���De�X�<ɤ�$���ڶ˞B�Vd��Q�<���p}�h�aC�"���YVI�<ѷF�*��i�Q�C�Q��)�5D}�<�"�4�H@X&���-r���pe�{�<Q%��6BT6�8�c��a��C���v�<9�
� r��`!&��h�t�W Eo�<�b�ŎV�&dKN̏4%� d�<ٗ	C�k��4��nĴ0��a�<��H�X ��Ґ�C&�����_�<�����%+�iP�����]�<�t�݁�:�{�&y�v����_p�<q&AT�2�b=�!��[��i3"�p�<��ÃLR&����^�����V�<	�IL�
w���G�O��PC�k'D������*W~��vD_�V9^�V�?D����¼X}��Q�Z�%Z��p�(D�,���T
v,�0�,��<˵�'D��	 (^;���&,x�)+3(9D�4��b�4*D��AѢ��|��8��6D�����5_P�z��R5Ҹ�(�&4D����R ����f\�_WlB�&0D����Ŗ�h�|u�#�gF��0D�� ����׈�r��+�HlaS"Oj��6LY�t������b�έ(p"Ov`"d��u���j	�/y�M"O�� "��vJX�2#�e����"Oꑱe���L�0`��ktBZ$"O�`Ґ^6]�j�����,det �"O���W�"O��� ֪�>Q����"O>���_�d��53�2A��%#"O�AA��P�P��@���):r���"O���EI�{n,u��̩b0R�C"O��ɑiDP�^�zV��*#����"O\L�e	�' �(b�
ҿ�<��"OF�)�)g��b�Đ;J�#r"O�,�G�ۃ{�Mҁi�d4}��"OD�c�1m�4��	]�&��E"O>��L�sРr�A@���Xt"O4bB�TР��Lc�J��P"O6xI�D;,�t������t"O��꣯ùl�"��G늬'qN5J�"O�]�EK4>��ن̎Hg�R�"O�<J�9�H�
�7oI@��"O� *H�o�	���DqA̸y�"OB}����'A�$	�J�G��!z"O���A�4{;�L�0jt�
��'f��\�l��!��'P�6��Ze��4A�zT�b"v}
���Ox`�1� �DJ����4�����SSf�r�ƒ�~�A�l�/�) 3嘷0Q�LB��K(�>�Hp@6r�r����U$8��E(��dKD�Jx�(C��(.+�"<	�e�ϟ�Ӗ�*l����%p^�h��'Z3!�p�1ߴ�?,O����<y���ҙ)X�����<��Cl�y����ⱦ]]5Vh7m�7M�U�.�VAwӮ������i���T,�un��w"S���=1��xR�i�џI�z�شJI�%Y�	*<�[S@�&��Pw��$l3ZH�+���(Ot0�cǌ�U$k�=|\��3���'9j�t���	N����ea"2z���M�$Zt|���dM$Z�Ҋh��I&>�m��hP��K�(X'C��a�2������������R. �2����1?��x�]z|�VE���9ٴX�ֻiH���	8 �l� �������dCϦm�����M{����D���0�4�S��F\��s���m��L��fåG|:�(�Z%>���%��'k�ݠ>�S�?��M�/�@L�S�M>k9 $B��5���AQ0�$,U��k�Iޭ:��$��(��z2D�|�1lw��9��?m(�,w��q�Rc`Ӏ�9��'�<6��Ey���������P=�`1`�G ^0�S��x8����O�OJ"?ya��U��d��c���*!�L�'�6�Hͦ	&������;A���S.��5-K�\[���w_�qr�'��| �̰y���'3��'E�����l��/hL�R"� q�<���ށJ���@�ƈ�ؓ'M1 $�	�����b�i�6XM>�&��T�\�ا��?ߪH��R�<��V	Cu���sMCf}:�h���d�0�X�ƃ%<��La'a�Ƽs�ޅH����'e!h�ԘWH�F}��?�?	�i��Or���O�s�� B�*�\���9�o��?ܤO~�=�|��4v�xT;bG�-:n�ٳ�S�p8JI`�-c�|5l�ϟ�ܴ�?���:(�r�ʥ.�j��,j&���}�"�:��L�q���+<O ��x}l����G�v�VM2�GՌp�p(;���:0���$�9ӵF%\�(�����c�W�'|��ө�$Z����C���gܝ�-B&l�@t(3W�� �ǝ����c͌o�'���2�cR��V�ְ,?İ�p+�f.���@|қ��'����<�?�O��L��I4} �$����&34�3��.$�D��cH��q+ǛR�x�hdį�0�e���M�)O:x��#�����?ɬ�΀��b�2=��s���I��cs�9@L������h&0j3%�P�r �G�z�����6/��x�	ݜ3�Đؗ�] 2��)�5 'ʓso�Q��P�#��V�;�Z�ڦ�
ֺ{b/ӓv�(�÷#�6IM�<�v�?��=��`�I1<�D�����~2ݴz���X�����q^�Bd&%��'��O?�$�%;?��V@��,M�U+�	����T�����
�M�"�i���\�HV��B�/d1�G���jf8��O����OF�O�b���ӯ
   ��     y  �  H  *  K3  c:  �@  �F  FM  �S  �Y  `  Sf  �l  �r  y  ^  ��  �  (�  k�  ��  �  ]�  ��  h�  @�  ��  ��  ��  �  ��  @�  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p͓��?����3&��H��� �R�ѧ�
R��%��	����J�7eBr�X�׶�yb���U�Lx[���l��}��ѝ�yś??_N3��F�s���; \��y�@_�-��L
͊q@�_+�`�G{��9O�qYAl_�|Ҁ:%E�g��PE�'��	؟��Ŗ��Pk�3a���ޞR�C�:W�4Zc�ćI:Thw���MQC�I<d�����C����oȔ�C�8�t�a�JU�`��Y`OZ~l�C�IpT>4h���z"����HX�ȴB�ɨ:ghU�k�[^KX�_�:���"O�6c	;���c�K�g��h���`�O��8�Ш% ��p�	���A
�'#�D@'Z��𤁤~l0 �'�`Da$L$RUˢ�̗q��=��'@���fbʁ���%��uJ�$�HO`�=�OO> 8&�ؚif���W�]���	�']d+&�A�x]u*�(P<����xr��"~Γ"�t�K�<D-B)�t�B$B/����IB�g�:�3����!���90h6j��	rv�d#LOD]�3IP�>�%�6�ö"B��Dgӄ}�O�b?� �`!wCU�*�I!c���h(�:"O.���b�L��Η�8!I��x2B@�O駧y�dP%1�jⅨ- �v� �!���y���8*љ�hW�x4��2��P��'��})ƀ�i8�� Tƀ'>`l%R+Ʉ,F�3q/$ғ�hO�ӿ$6l	�R ��y~�#��H�!��S�'��؆��I�0`0���'3�H��ד��'�
u�F�O&���0�)�ހ�`OXd�CЍ1�6��v!�(rlrC�$6�S���'p ���ӭ8�2���Kڹ!���
�'9~���KM>�qT�4���	�'�����Q `f�-��Э?�n���'i<��sJ�5Z�tA�fI[�<Ydޱe^D��/�%��a#2�z�'
�~rÁL������8	㞁:u�����I�o�Ad��7Q�~�R���d8�C䉯�ܼ d�|S8Ă�N�$t�B�ɘHr��C��#ߖLXB9	�	L��8hv�}F�$'ڧR���Q5�>D�(��O�@ D|��i�0'���;D�4�6�Ak� �i���]�~Y���:D��YOH�u.X��UC�5:���S;D�8k�&�&%�x�ɒ�ڪ-��4c��9D�r��:C^�D P��<�p�@�,D��q���"d���*�<K��pb)D�$X�'�|����j�#f,��%'D���b'Ú&.��#�� H#�1��!%D�����*y�7gS)��ٻ�-5D����D�:8$�ڠkQ ��"� 8D����O(H�ʽ���i$�j�)*D��H��1l���EM��i1S�(D��i�C�v����B�Ťgj��sh9D�ԩ�����D@W� �& z+4D��&E�"[�	А�Ի����	2D�p��g�Rt�T*�������Ñ�/D�����1M�
08�P�g,V@k�d/D�̸%��!Z�eYsd�(L�0�c.D�pX���
fp�#S�;+ل-�#)2T�4[0�Y�C��R���b�(�H0"Oh�Ц�V��z��I�" ��`"O�)��C̆K��%2R��:!��	"O6��t��1Y�6��I�t�*��5"O�Փ�-�2%�亥LO�r���"O�+%ِ+;�aF��#_�.h�R"O���ț>f2�aL܉{��ձ�"O���h�&=��JŬyz���"O�|��kK 4j�I0��S�Dx��""O$��@��"6�1���Zp�8;�"O�(+�U�P��	/ �	"O�����K G��]��i]�p�l�)�"O���wh��� ����5�$H"O=�� +�H�O�R̪M�"O�8�(�Θ��!��(��"O�!���E�,����=��$%"O6�q�E3�~ɩ��C/.�D5;�"O~���˻}T�S�-� �;"O�t �)T�f�BJ�g���"O�4ȵ�K��%8Q��f�j��"O�5�G��V5Th����)ή�J�"O@�k�,B=t������B��ؑW"O0�÷A'M�zKã�&F���"O� �$+ްc�: å�[�N9�A2�"O6�7#�"�<�3$�9_�:!�'"Oč�b�/�d��^',q�""O� L �FBS�JF�e�.#j�t+�"O�X�2Tq���*bCہ]���g"O�T@ 1U��D�L?L���"O���ጦE묈�� ؑ!��D��"Od�
��Wp�Fa�Do)
��,�r"O�����&jj�-`-ٜP��-q#"O�ee��[0�(rl�"ϰ9c"On��Ǐ�+o�T��J�	�>DxB"O(��f�1N�~�J�*�D�,�S�"O��*���Ӫ;�|�t"ORy�T��8�i�({��R"O�)��eZ(pNa��)�8Z8*&"O<��F�R�8chS�]��C"O`i�̉��(8Bq���]�Q9�"O��R�M@$lkJa�F���BsIBc"O��wc�3d�ЁBA�4�(�1"O��S�,��f�l����6.���"O �:S�T�&� PZ5�Ё%�ik�"O�'lX/��gH0�]"O�� �O�(�hY�A���x�v"Obu��K�&fb���O��s�Ҽ3w"O��Ac�a����୚�d�!��"Ob���,��z�t0�pX#9�pS�"O� ⃆�~������0E�&d)�"OveȦfY=*�*	b��L�<ʚa2�"ON�J�G\:x��� ��V� �#r"OLmFj�,Oz�<���X�P�zQ��"O�i[�c� &���ӫҩ�x�@�"O�`G�� u�2���>k}�R"O"��$��K�Zi�N��XO<�"O<T��كNed�a����0K�P��"O9Yw���&ա1��NG���"Op��
�/��"�@"A�2��p"OJ�a4eȵ6� �Q�)#���h�"O�� 
�D"���MO` "Oƥ(bgO sk�13�[-JNz-�"O��@��Q����M��J"��S"O6�1����I.�IQLH/ ��P"Or�J	֞@&�����R���"O�ijt�@�lcj�S�*I����1�"O����j�&�y�*��.��}�E"O���/V���Q�Ӳə�"O�|Q`v�y@CgT ���ȣ"O�Ԋ�nQ._��xf�-1���"Ov���!�"
P`�{AK�7 SF��e"O��@��;$hYaQ�W�jD>ic"O�cw��2�J�#	�<b���"O����Eכ	Z�Q�F�L>O49ِ"O�Qq�+�4𒩀�K�1D�0��"OX�%L�<04y���Fs�
m�t"O| 2��/07���i1�|"O�yx2�HN�Vr�J�p��D"O��S��fS"0���ܯF�!"O|4��j6-&�r�
�@`�d�e"O�l�`a�6J���E�ߙqY��pr"O�]n��f���rH� `��}��"Oވ��,�/�,�˲,N���9�"O� ӵʝ�o�� Ц�\1t�u#�"O���	^4������f�Łv"O���J3{��z�뒓/� X�q"O���V�J�H�.��"��"���`"O|%	w'[�?sF�f�+(�"O��z���KZ0��IU�7
ʁ*"OvɲAۊ*P@��3(�/�Ye"O� �X��ΐ���:�G7r�i�"OF��Ĵ,8a3��P�M����"O^�1���l<@�"�!��@�"O0��D�u&�|����!�v���"O�ՑEl��{�b����@.�Q2��'��'<�'
��'�r�'��'�z�`��1:��:u��_f�9��'�B�'8"�'2�'��'5b�'��͉��μ2'�(��c�Uv���'��'?��'22�'8R�'��'זd�g���I%�R%c�Ƣv���?���?����?A���?����?!��?��e��hZ�S᎑2q@x���^*�?���?	��?q��?a��?����?Ʉ�:lrJ�w[Ь)���?���?����?Y��?	��?���?�ŉIo�D��NAz^ {t'���?	���?���?a��?1��?)���?yǇ^�f�`�i� �Zh�UU`��?���?q��?����?����?I��?�6�՟y7ʤ���Ƕh�V�g��?a���?Q��?y���?q���?���?��ݸO�^�%V#�@l�h�!�?���?���?����?���?���?q�/C�Cg:D1��O	}:�,�����?����?	��?A���?���?����?�E��*L�*���� �{XP��)���?9���?a��?���?Q���?����?IT�ɲR�]B�EW7LP囔�L��?����?��?����?����6�'≌V�f)H�gP�PF�T�4%η4���?�*O1�����Mc��ýc�f1 b� ��A��	>����'�86-%�i>�	��M�����	Fp10�R$D�S`E�jz�f�'��p��i�	#�H�)�!Y�'SM���l�8�e�@hJ�"�^��<����;ڧ��܀HZ�!wؽ�BJ���)c�i ���y"�����ݶ�\��_%QGR t`
',V�mP�49B�8O�Ş�8Iڴ�yb,
����� F;6����yb���9vt�m��1B"�=ͧ�?����I��;�J�]�h@r�Q�<�,Ot�O�]o�W�<c�xB�&�8K���zՌ�?�$p��g� ����M#�i+�>!�OOӲ4��l�s���
 d~B�٘i>�8pHU��O*���������3q����%Z8�ɍ"��L�'}���"~Γ-Ϧ��QGЧ�$|��&Г[b��Γ>R�vC���D�����?ͧByD�rўY��[��f����g`�6G`�|��^�{��6�)?��
Z���g�c����d
�!����F�`+�T�����Y:��,%�tE����|�J�)��y��[/\`���mR��y�O��t��Á���aQ*����/��	�P�B�����A�����8�O3��m!�(�̀}!!���+��X9W�2I(��M�6>B��h��E	(�2t�9>��������n8���$]+xmC"O�*2I��^-UY
�Ѥ�	UF��pB�����s7�}0���M���?�����Ƒ���_�L�x�S�gU$5� 0�S j���D�O�hsD��O�O�)2��X}��0٣-Ǆ ��<q� ���M`�@�Hx�v�'NR�'^��f/���O~��Аa��xAs�ѽ,�`)��̄�j2��՟4&�"|��PCԥ�"gK�.����S�
z�49r�iEr�'���:!�(O~��O^�I��`�ڳ��Q�Ƅ �hM�\��?	�ΰ<[/Ot���O,����q !��"+d͸`g��Q8��av�6���R��.������<�̍�+P�ǥO�\��|L����v�w(7?����?���?���X����6bM�I���WS���)��?)���d�O��O^�D�Of!ZcI�_K	�6Eϋ$�=9���i��B��,��ßH�������{�,��'"��y�AN��x�����n���l�ٟ��I��x$���	�����'oպ7���5!X�S��؟t��:��Z����|�	ٟ���ڟ� ��z���'oB�9�lл씤sG �&�F�@2�d�\��?�D�O^�d_7k���!�x�@I.\ ��TE�*b�d��Ms��?�+O���T$�n�S��X�S*\\0y����H?z�p"�B��ذJ<����?m+|�����!M{��<�X�B(��<�&�'�r�[���'G��'c���',Zc$��H��yR�0:-���ش�?��9m���H�j�S�'-R�`ʐ.��zUFxS��\��l6�����ß��	ڟ���ʟ8��y��h�d��G�n�m����c��7��5u�%���䟌��H��E`g'O�b���x�+�M#��?��lw.�1)O ʧ�?��'P���7�S�	�2Q#�M�R=���6�IA��� J|B��?���:�<��D��Y��P�f��&�vq�R�i��
�(�O0���Op�Ok��.z�X�­�
p-p1,���'~���^������@��py��'X@Q �-�d�ab� ɬ���)C&��e��	����	���<�/O��鱏�7a��쒒�ոA�@��Sm�����(�I��T�	XyB�_:m;�S�qj�ԢCDΘ��)���#��ꓣ?a���?)/O����O �S�T?��&m݈�:��3���Æ�RUn�>i4��>��!�+6K����j�Q>�*fB� ~��7�[J�A�s/D��R�f�-'��N^�dR��)�m��̠��X6v���,Nie|����p����NR�'���D��&�t���M���K�>#���9�m�=	Nuғ)K�X�,<����.pPfY<���+H�$�0`xPh�Q�� d�Pe^A^��pfepC@��t�#AJl�W�ג]!�љTc��s�ĳ�
v*$�����O����O�ܳ4LX�.=�|A�b� Y�D�Q�ͮ|�JuR�e�G�	�޴�M� 	�([�dLɋ��;&��X��ApZ=@"`PS��`��˶p�t���7-w�t��几1Sq�G�O%�*qs���"V5�%���V~��P���'��6������r��?)  H�8t���Ϩo���Ђ��<Q���>iƄ���(�h�	��Rd�Ċz�'~#=�Ā:�?���J�T���Jܾ�H�D#��?Y�e΀��%I���?!���?����.�OR�X&E�|���\�:ɪtS���3<$ne�7������Q�F*?g��ӱԟ��D)Q�Ř'w&��l{�	���X�2=`�҆��	�2�1f��!+s�F�N�$��H`�RVY�$\���'p�DsD���w�~ܹ��I;'|124�'�<]yG�'�6M���<����]�]]�m��c�6kЬ{W��gR!�D�O���ж^UD=
$I%b6���s$�O�'x�I�b�',�	�x�@� ^w_p�Y�b�"�H��%.����'2�'yC��TR�'��fԸ$W�\�2�
B�l��i��-�]��_.
Ć���	�')�B�С�Pn�'���	5Ǝ��ɹqlPs���
"���t�&`�,�F�HD.��M����K=Xr�O�}���'DF7-�]RjT���"�ܡq�\k<pn�͟<�I�����ʟ��	A�S$�'��5向�Q�V�26�]��M,�L��8�1өUN4���I��|�(Tmt���4r^�\�hkF����M���?�)�Z���-�>���a DDR�� ,۸+����O��G:8�Z-�q��.-�tD`���b� ��4E8v-�Bʐ>T٪"EŕL��%IT�6�d7����G�.5��B�x�0%1w�؏Axx�Aǐ�9���F!��J��[��'��~d���M3a��4�'�欑p���}��X�F�`?F�j��'��O?�ɘ#��{嫏pO2Q�5@4Q�"<i�Ńj̓u��F�k���Ĕ3K��T��,�#��X��ɲ/�E�۴�?�����`�P���O��� ��й9Ƨ�m6́DZ�iw*���тs=h` B_�xdE�%!��8@%�)����*��h�:��ᄇ/^��pgď22k�=�G���@[�'��C#$�+�gۀ_�q�g�E3� ��U4��R�V�-6Z�0��'�Z7�������I��y�T���@�qM��[��˦d��<Q���>I n�Oq�I���$+Ԙ�[�MR_�'@"=��'�?��V�UH��zףQ�u��K���?a�\�PXɢ �?�?1���?A��t��OV���9?N8I���"���U*߰R�$QR�_*\��8"��J�8��ݟ�P���
�'��,���O!]U���@:F�������/n���[��_�.��Ս�����2@�5&�Y��IV,���F��"Y	A;�~��<5b��ĝʦ���4��'z��'�Hm!w
KN�6��M����'6���j�xB�%��!L�slƃ"#=y��i�"S��&dι�Mc4NF�?���)�F Q����?��?��Ƅx��?�O@�i[�f{�d��v��q��qq�_��!k�Q��lZ/	Ar�����'�(OD���N��;���k2��7�A�0�M)dL��ĭS7]����c�R�8s�8�A���͚v�2�DZ�R��r�����p�3ֈǔ?�(=�}���OP��?�ʟ���w�ʉ��옷hQf���cE�'Pў<JՇ�8���Γp0�
W���pܴ�?�)O��������	؟|�Oz���"�H? �0蘳灷(��p#f�)n��'B�B/[�Z}�pD?��X�P�7�|�*%*�vl	!"a킀j#*�4(Zbb���9_���� "E�@0#�̅�,��kO
�g���X��j��z�򤈪W�b�e��n��\�O��9����s�:EZ��քZ�@�Q%�'��O?�d��i��F])f�JQ&��B�(��dO�I�j4��&�g��Q��]�M����"kir�4�?�����Ů�>���O��d���� �i�
O��� &z0f���9�ů�� !V�1�߉3lv|YQO5���:	hk�s�:������Ҩ�SA�N8���M���|��� qޑA$�ƙD�:p�0l�f��;���0� ��ʈ ��'�iC�O��|3��2�)�矨��[�?�RH{r��D�$wM2D����T�p�t����'3?Z����/��LP��4���W�]l�i�P�P0ɢ4��-j_!�����)R�" S���Ʃ5-(!�ʺQ7��󂀺.�f�A���?G!��
�AH�1<�ڐ�0�"{!�d6��!'��1�n�ׄ"�!�$�8g�yCc%K;m� �(���	0�!�R�~D��Po;fz�u9���\!�
6lQ����GD1cp5 ]S!�߀`���Ia	3ObT* ��m!�:d��
��[}8�q+D��{!�$Þ Kͩr�[�t���E!�$�$.�v�[�J�F�r`´JND!�� �;�DC��f`4@L7n��	��"O�u �+����b���G����"O���S�[)�ȵc���wj���"O �+���I�\��`ҩ!r��"O�yR#�#:���)�,CI��u"O�p2�C?s��0���t9zm�t"O2iX���kމ����6_9�s"OnY� "�9;��țVd� X"��P�"O�A�T�^�N^tT�2$�6ED !�"O��xF+�)A6^Qن(}��<I�"O~�1gǾp�%�Ӈ�7 ̙"O�UW"
5	+ @�l��H+(T9e"Oȥ��fX(Q�����\�h��Tc�"OZ�`p�,_�h9`T�ʔqn`�"O�uAՋG�fx�蔭�	�h	�"O�u�6��^���:��vl@�A�"OJ��p�L%	�y��J
�d���"O���ѣ[�W���`C�y���V"O���1�,\�T �^��|Z��M�<IJ֛/��B'J\�E���h��^E�<�F�� Pa����pU�d����.t�	v	*?��	S�OP�}��]]� ��F��
[f�Aw��#z�.�ȓT��R�f�
��`3v������o<J��D��7,FN����U8��r`�](?�2w�̝W���f�<lO����"�;\,�y���8+�50t��!pEj)���4es�L��j-��I%�/o�@�P��p�e���8�	�.�f|"R.��S>��X�Sy�'Ζ����7�F����3] �0�ȓ3b<qy�K��b�&1+��d9'��~�ѳ����2�d\v����Q���8*�;k���0���Z�!�$R�!9�!BP�
+A�p�RM�,e��6,�
Pc! �ʠh���'�F��RGB�x;�f�?	iL<(�/�m�#)��G��ڳ��[�J��0���,z 8�5�ޛ9t0i�	�'j���ț�D1$��4 �(�ja�}2���©kd�/�Ēp��"S�T���Q)���ɄL�%tX!��&]ìŻDN(;���v�eÌa�1�J�D�����.g�@S2��T�I|��Ù�J �eh�l���9�z��K�u*� �Ҡf٦�	fdR�_	�lyAL�m��c�eZ� �&���޶Wt���$ō8�>���gP
bB$q�&��?
������W�|R&��)�0�S��vӨ5&Ζ<@8�e��.N�h�q�J�Pxj�m�Q+ �pJ��������J!���Q֤H4V�T1��L|��	�TX|������<�<]�bj�1[���3�"E4M�0��%3cFX�uf����Ҍ7��O��ɒ�L!`k��*@*Vg?Y�����H�'#,�bT	B�z���8d��MgF��4=*�2֡)Gj&p�O�R����IF:5!�@݄�����J[?��%̒I��K׋�=�BpQ�[V}fO�����
/X���nل�HO ��_>)��Lѕ'��S�[�H�d6$
�=K󌎢 �IF}"�B f��]��@�4VL�k�"�'�*`���,���>a��4�D��t���']��	��� ZdX2�A�=��=	�=�%jBbZ5s%��ɀ��4j����	Y?��Y��p�/	��2ҥ�:�����Oj��8z���x�'��CD��4u��Q� ��_���޴3@�YT��c��� iG��5�^��b�'Q��ɐ�ihF��oAc��<
�.��]��V���#Ё؝\r٘�Y���]2�)�>��֬'L��䂹���D��_�'��HQSF�9���Ag�W�,��,��u儙�W�.�~�����Xq�IG}�
!#��iFמL㊍��lȮ��05*�f�t��d_w��㦫C</��l��l�,;J���-�z����5|O"�㤯K,F#�] E��$- �d8�Ϟ`�.�D~��
8J\�i �"ˉH>��p��QM.�2A��[��p�Gɒ,:(�� 2*4�t�
d�C���!t�n��hҰ�ra��7��.U��@Q���ҭ�G��]�D���+Ĺ�r'`aP����~�.�W�BqV ϋD�+�a�����B�^E$M�M{Ƒa�J�!�����C�3a�z�kG)[�,ʰ��,}4=�ɀ�wy���S&ْl~����	8t�Ѳ�#�3��c��I�<=^�AS�K�=Qӓ>o@��f ǽmly��k$��Ukل&����@�٦��=i� ϭMTp8��V�=����c�	�3R��{e� :�fΞ<&P�3�X\N|���A��}N���u �++�M��\�'�L�q6��C��Y[�g�0}?�q��t�? �4¢kά!�h�*`Κ?.n�C5�XC��~�MǼ�h�QȌ?��3��O�u��܀\H���d�T,8/
e��V��@F��k&b�{U ˯v:d�Sf0�@br٘ �ҷ%�Z�� �'x��T�'�,sъ��G >���
 q9Q����`�<�r��+W����Y.�ɡU%���Or�sL<I +��<�4� /U��iEh��D�Pѳv >�O��ݿ
�@<�t(��
{���Lؾ���'��DȞT<�O��	�?�
����� �m3 Aξk_*�@�	y؟4#C�
4� Q�b���� �2"$�yQ��P�H2T*b��� �P,!F�w8��Q�N0(�(�i���ܼ��6���@�B	]�f�&�����E7�)n�4j��hT&�gTZ��$J�P�FIa�
O汱B��0�Zb�ňF-�t^��K"��2c�F�2v`�3s�Y�D���>��Q��0z�|@
'��|z� ���6D�P��<��(4�ӈ~DT�c!�ˎ�!5#A��BLŀ~�R��:��K<��έ:�h�S����E�Р�w+Zi�<�ۼEdD��e����N�*��[f�<��[�{���! DC'�p"�	B[�<i��Zj�Z���ۇe��8��o�<A�`�"c ��+ ��)��0�jm�<��̈�%B���K&#�+9�*C�I�]	�L���).T�yӣN�d�B�%C�,B�b[==nfM�P�s�B䉤p�BP�R��p�B	0.\+%:�B�,���CKոz:�m�U�ƈ$HB�I�[��3Ƌ��#(�]0a�U� B�IC�MY�N>5b�U�A�DCWB�ɱp�Fh��m�����<B$B䉀c�R7Nڒk1Di9�h�Gn�ȓ"
��͵IA,�%a�t�ȓ6Ԧ�KEV�I�ɶ݇ȓC�*|���=0���unL�vp��	�J���f�<x�ؑ����.b`P��ȓo��0��kĿsE>��&oхZ#�X�ȓ~�b  Ę��x�u��T��,��q5������x����1�X�YX��!ʩ���ž4B����� p�r��ȓ_�� �4�B*3	
E���9Gx����%p@�� �2?m��C�d��Yv�݆ȓ�>�y��^�LM��C�ϔ^>t��ȓ�f��q.��R�0# 2 ݇ȓ]�ʽ@�G�)rnp��L�y�f�ȓ!%|	{�)�4W�Xc��6���ȓ,�.!Ȕ�3g�!#�L�t�R=��EE1��iT;1n�cU�Q,h��B�?��U�pH�;AhP�k�ɷ{��C�	4��8�+z���@�
�b0xC�	
Ϭ�ௐ�:��h�FgŶ?:C�	|���!!/Z!H��چ�A+i��B��.Sp���`��pl��3��a��B�P�|�ɑ��B�t�˥���c�hC�	&!�x5�G�k�-���VC�ɐ�B�R�Ӻ7i�!�C�b�$C�ɲp��y"���w3���1��)9����1t�R�F�@t贈�(�9L�!�DE�O��b��3%�$YQ�Ŕ(7!�^�c�H��m]�Ad>$���"O�}��'.n@{�C� N�;�"O�<�%k�
�^!�b�3d�4�:�"O��m[��8� � +��"O� s�
����34@� �ޡi�"O��)�j̿,�D삠�O{�v�"�"O���F
�m��؀g�+��Q�"Ofԡ��Ý^�`��f��B�HK�"O�����J���	��O�@$��`"O�����?�>$s��Y�Ya"O� ��X�����,���σ,�Z�٧"O&�;�D�9o�A��i6���1"O��[B�\$$X�	�fP|�&@�5"OР���?S���a4��r}:7"O>�j ��A[r�z�M3W̅�"O@����ԿRg���:a���"O�	
B�� >q�t'Çw`@s"O���� Ű:6(�jv&�9dmp�8e"OZ���䒚��P#EL1M�����"O���ЊgI�'��$&#�Y����yR�P�zW�ĮQ�ڼ��Oȫ�y��R>)�Dl���4R<��hď��y����X7��0a��WvX1���yB�Y�BHbc!� z�$񑰄�y2�T�[(,���#)Z��$ �yR��Y`&A�)#@<�&��y�F9!�2�cɵ*�d��H	�y2���,��1�L�~24���Ȧ�yR��3M&l��#B�|�B�1�J���y2�۳/�����ı@J&��S�D�y�TN��]�7	W7-�
�BcZ��yR��9dPj���E��+.�]�!��y%ˡp�@Y�H*T�P(à7�yrF�(P�Y2�Ο�ww�)A�`�"�yRn^�#T�c"�5u��Re)���y��O�tys��:k��Ҵ����y�e�
zu�B5*ep��ԈI��y��Q
>��;G�����Z��y�.4gޱ0���D��X4���y��)MЊ	���L	5��yҩ;�y��B6O�P-Z�O�9yuΉ{��R��ycP$Z�9"�na�������yҩ�,'JL�p`��.ex%�����y�	�.�����Ɏ/P�p��ݍ�y�@��(�Y#�ן-�@@����y��*.x����&rN����yNE�|� I��_4y�\�DS��yb.�	>�^�i��,�`E�g��y�HVV��b��	�(<)����y2�ѾZ�4$���~�&����[1�y��غ2ôlj��N5AT@�83F�yb��'>��o(��e�ò�yBlI		n �P͖5�`��u�]�yAPJ�Di��/ͥc8�x���y"�܀1��\8���w[8�3�y@X,�$Cs'Q6s�xb���y���/K�T�y���S��c�	�y2�*k�XX��b
}�
8�Rd��yb	��b��`mĹpy���@�,�ylM�[����jpP�3��yrI�x�J@�s�R�d�`����y�͖"dN�@���:Wi ��j^*�ybM��N�@��$V��AQ@�/�y�(F�@w�9`& �=�>�P�#��yB��+'T�ˣa:'�.��,�y�$��x� q9�M'&�eRgo��y�&�(Ad��Q��ì%=�4kv-�9�yb ��:��7�F�[,����uB!��I
&��Xf〢g����G"�l6!�d�Q�R�)�|���R�[.j!�  o,e���=|�k0�B !�D��G;��M�n���B�S�}!򄂴yo��Q�ǎ{Z�4ҥbƗ0a!�S�����M:iBH�5K0S_!�� �hRŃ-J�n���NW�,�"O��3���Q�ȱ��A�yH��p"O����64vmɑ`�$�N��$"ONu��-k���ؑ��3jl��"O����Cˁ{֩�`��x&�L�a"O� AM�e��n	/�Pa�u"O0L�cZ�9���J ����4a��"O�y�1n2�8��Ԙm�F��R"O�q���85�L�+���s6�#*OI�p뛐i�С`�ߑ2� !�	�'^� I�\��mb���<z����'Hze�@�	mq��{�B�.u�ʕ`�'�X�k��Ȕe���"ǌ�k�y��'`2��V�HZ�		F*�f��	
�'r�%��a��\�F��`\�I:�'�pB�c_�Y]<��ă��<Q�'�訡$�J��@#���f��J�'0�é���!���f>��)�'�@U�6jn��i��Բ	������.D�R��.L�pS׀Q��fy���1D�؊���K��y�:j�J��.D���2��*R?��z�Bm�"a�T--D�pXR�]"FOȬ2���1��\#�(D��b艕p5q�G��7�����F'D�Ls�
Ս>���PbX�0t�3 8D�,a6ĕ#j 
�Y�dǬ]�ȝ���(D����"�v|�UEN�Z�-	��>���M�Ӥ�6G0Y����6	("�����?A�D )�И���uPpm���MD�<���ڐwՆ�k�O ĠX�tDj�<i��Ū�����GR	q�I@7'j�<�6�A"i��E��		�48agL}�<��mˊ�ס�����eLW|�<a�ԧn�h{�� '�H���w�<���	a�A��K�;��Pxvću�<ф�J,bW���V�Џc��)�&�w�<1(�(>�1�K����諶��H�<��y��%�@�½K����(-!�ψi�����A-�ёq�^R!�䔂!��Qi��`�Ҙ޸�D"O`��R�K���K� ��"�<��"O��)����]Px-R���6�T	�"O���t�3%���$�0�|��w"O�-3���XE�0�ӡH�iY�"O�F�\�ARS�ȋ*���r "O iB�a�'xӄZ����,�"�*@"Ov z��f��!�!i�=��Ě�"O��"�H�n¸��j�钇셑�yҥ��6$`X3�A˽K�d�
4��y�ϔl����._>|5���y��L�Y� ���ɷ7����m��y"��`��,�#�T�]��\���?�y��.f=�Ib'_�kU�2q�<d%��F{��T�Qr<��4k��{���ă��y�CZ�Ae#�m�:k�gT��y� ͝sT���!K�e����@*B�y���:#�6��AgN�\[�4(�GJ��y��+©s�C�Q��i
�d9�hO��	�6�qc�D�P�1ëU�2l!�DABϞ�@�?�f%飫�!5c�)�g"���-�$sd�IT�Ov����'���	��ēV��u23��3�*u�O~6�R��0>!5 �X��\�D�5d<%a��
m�<1$E�FR�[�k�5䈄��`t�<� ���s�ЕFFn�Y�L�ش��"O���!���qZ��ɨRȪ�2"O R��^.pC �`�#S�KB�'��'2&ͱA�"4�x��H�6&?�90	�'
`�G�o\X\�!���}�D��'u`�q J�$��%r�a�.
���	�'cƨB�b���Z9Q�z���'���d��7Db���ŏ9Pb��'��T�a��,P�0a�+�J~:�i�'� ��P��88Rt�P�C�@%i�'�z	8##�
ML���Dn�C�09[�'8%X%b�0��3���n�8Đ�'�@�C�?<�]�e�D�a��51�'MJ�y�o�]^:=q%ϟ�S�}��'~8}�/ �~�����2Tm��3�'9�,�`�̮Z@a�b�ά[^���'a�Q ��j��=����"f����'�U�����v��U[�f`r��i�'�p@�2-�E�hLp��ڨjF��
�'0����;S�Щ� �'r}��z�'������ u]��r��o�Ĳ�'` ��5`մ	n!9Ri�$2.j�I�'�=�u�.>�$x��W�&�D���'���R����3�Q9/";�'�T)k���ݒ��be��+&6 ��'����[�l�F�X%:�xs	�'����t(��<�L�wfUhw�p��'��mBth߬/��˗�]�im$���'� DR4B�Z`���Zyp����'@����l�a
Z<:0�qkH8��'��X��K�U����-[/v
����'B ��PŞ?o�E ���7YO�t��'ǒ\�_j8��(AL�P�1��'1l 8G5�B���8G���c�'��x�f�̹.��'���9����'�&����Ȣv��Z�I0$@i��'�����ͱQ�@�[��3gn�i�'�`|��jS&L�x�䤚+�����'�^0" �W�6�s$��%��C�'������&6�"�q��� �����'�B�6��H��@qE� �-��'BF!Pg�T�ePtI7L��	7B4�'�L����~�Bu�v��-�T��'뾈�KO�6�A�O�[0�0��'���Rf*���Q:5$^�
*4��'kFhaE��=2����P~�N��'F:��኎=�h�q��	j~�+�'���I���H��0��H�5Z�j���'�R�P�,��;p|M�`��Gq�4��'1���#��w=\�鷏��D�
8Y�'�J�|���+g��h�#��y�h��0���%��cda�cEO��y�ǚ����!�C�n/`�eY
�y�2}�b����&oe:0C���yBI�:T�6����P��܉q/"�y�!��a"���Cv���dT��y�FZ�9�=�A��1!���W"U��y"��$�Z��2�4vwr�� Е�y2I˳F6V%��$o�tÄi��y"�O�S���s	�0]��)!�K���yb�\�h�M	'��
�|Q8����yD�v&jQB�I[m ~eX�I��yr�͑Z�f)h���_���H���y�\�k��}�`�V�K�(a`Oӽ�y
� ���4�ʷh��
�Ȓ6h���"O e�`(��Haf>�,�1�"Oj0"$҆O@��[�e�;7t7"O9���]]}�a���v���"O�hK.X�5����� .Z|�j�"O4�(���<j�Yȃ��b�4���"O��IHN(~��bA��|nf�`U"O�8�V $b��!Ht��dq�b"Ovx����%�
A�5.L%H,R�"Ov��5*^�<��eD-V�W  �b"Oh 4[�+qz��j��]�ȅpD"OtR� ��"vurD�!}���u"O:}���D�O�F��t�C���1��"O��J��v)�F���V��j�"OT�I b�+Y�H:�锽+'(�C�"O
�Y�,�@�d�A���4���"O�[`hB�tq�i�p# p���"O\�sT�B�Wl��K�@�N]�5yS"OԀTCI�i�RH93gB�1���"Ol���dă_�h�� U�g��ɕ"O�A�s+ںS��\[�7wv���"O�����ʩ ؒ���c^?oZHT"O��a&�:do@QXF͓�DA)iQ"O�9���&,�<)чk�����"O"=���W�2������, ꕀ�"OBy�)	�=o��R0O�y"O2����H�8+�KC�]�j("O~�y��ay��@��:��B"O���p��0�lQ�@]=U�F�(u"Ot��G�(#`�����,e���"O.��i5+G�$
gˆ�*�� j@"O��&��P�����I�(�%b�"O���t��;D�H�sOτH���s"Oy��`g^�z�l�-}��LI "O�]ň܋9��T�Q�D+u&p<��"O�(�0!��gT
%yPʇ�?$��	"O���Ug/,��0�")6&��8"O����M�2��}`3��,�=�u"O� !Ga�mw�6�������,D�� ׫5T�������n����j)D�,!��slV��� �� !V�&D���N�A5���b��s�	we(D������j�����"e���3(D��pE�ٿR�H�RQ��4Gz��&D��W��t,\��P�I��@���8D�,K��S�P� ��+�t���7D�dP`╉8�l%#u��y>`¥J5D�p�&'�5\�V�s0(�^d�`�%M(D�L��cX]��B "�"�*0�8D����/���^�����[��(�q7D�H(p�պBAv,R��Y;���ӣ�:D��3��4!L�d�QELQ�hd�%
$D�hp�P�E��q�wgטn�:��M"D�@�ci;� au�3�؄�B�3D���dL��R�N���	�t`���u�&D� �G�J5:_�  �d�7�Z��f/%D��`��}YDI�A�G�#̰6�6D����`ܖ%�sbٖ\����"D���rm��f�hu��i�pb�&-D�<�e���q��q�i�?]w�ab0D���I:-g��[��X���2��3D����l������� �f:���1D�����[�8[���RA��sql�q��+D��B� �%d�,�����s�:𸗀+D�� f��喊z�r�%O�*y���v"O�	�e�,E��DHȣ>r�!Pd"O�Y2T-!g&T۰=!@��E"Oԁ9T�l�����Le�Tm"�"Op�(�/�\v�yWC��;�����"O�I9�Â{Q�]���w�Ȅ�#"ON�g�E��(��S��)U�de�"O<Lk���]v	�Ah�58]
t�"OB��HY3$���IV���I\(�C�"O�X�A�,�q;�&�J�s�"O�=��+J�Ll��C�O#l\��"O@\�B��)˸�z��C+f� T"O�p��cU-X?:IS��J� sA"O�`���������⇃aYju$"Odف��<\��e���B3m!����"O"��Fe�~���𒏆�f�uzf"ORmi�?R�6,%�ֈrY(���"ON)y�g�QR�A�(׫E���J"O����Ø1�.5�G'֘G$���"O��s�Ο�eS�D�NH�*�B�"O�s��Z"c�ʤ��&ٙ]�jȩ�"O�lpЗ6BuxD���\�*��"O��:�N�K��� �(��C+�CU"O���!�
�n�\�A""���"O���!7X��Vo��c��a�"OJ�;B�E�C�n$�t(�:&�m"g"OEqD�z�~`��H���pS"O�<�ҍ�&yyJ����Y���h��"OL<�u��6� ����9:���c"O���f��'��#� ˎ��D"O@�!���Zu��� ��uv�as"O�!��l^�U�FEʃQ^�u��"OD�{�+��b����3@GI:�"O��A#�y�puHe�:$U�l3"OUA��M#l���KS���"O�M�`��4�8���F�)E����"O�hyTG�:b��DR�Q)B9��
w"O|%a�OZ��1�!N���Z�"O
��*�
dؕGF�M�h�"O^!�0g?T�LMpV;`(	w"OJ��A��j#�S�z�>lPP"O:�:T�0�DX�ˑ9��3"O�-��٧ ����끀epxd��"OpĢ'j,#t!��ր}�xy�"OV術���(�����$٤W���+�"O${�	Ց	-�K���v���8"O�����Ŵh��0*D�+3�v1��"O�$�J ul���/��)M`�u"O��e�%-�AC$�3O3�Y��"O؀���_�+Rz�R��[�3d�R"OmztG�%?�t5�'�<���"O6Xhb5��v䀙-�� ڀ"O��r�[�5@���b i�Z��u"O��T�Ŕn�DaP+��m���c4"O��R��G6%@�h H �Z㴩Ȕ"O���4H�$�L�q�إ^��e2�"O� #�g�,��ݩ�![�|��1�"O�5�q�N���
�"�,L+�"O �sA	:נ�� �(�431"O�|�g	ޯG<%����.����"O�[�.WT.%��/\�@����"O,�(f�F&�RK�/�$����1"O�<�B�#
���*!]�oG��Y�"OB��DO!$_���F�i/J���"O� ��"��x���;}{6�1"OPM*��e�ĭ�r�^�}���c"O�,q�EK�0��疓W�>u��"OܑqBgG�U�p9�r�#U�D�K"O�J$K��ZYLT�`c�?K��	�"O:�KPP�{��Y"�-w���8�"OYk�)A�i�
���b���P�"O���ܛ���"Q4���z�"O�M
��55�"U9�(��1x�M�"O�%�ЂP6�13��8\I&��u"O>�v��b#���b&N0ʝ�r"OJ�C�� ��U�DGI�~;��9"O&�r��	S�t�s��;ƨ��"O�����Ie̼�{e��g ��3"OP}�RP-O���''��t"Oz�����ova��E\�r<J�"Om�̆*T�f���ש+̼��"O��#�G휵��M�'����"ON��LĮh�h{A9n�����"O�M:DN.Kj�aM�f ��"OȑCEDM;��@B��u��0�"O&���D�(BI����R8iׂ�� "O�I�5�N�z�����.[��-b5"Ot-�$��,8�C��V	f��"OʔJ���o�iKs��Y���Q"O�]S�)��w}H��-f�}�@"O� IsN�er�l��Ϳ�*�K�"O@���Ǆ�5|����j�c��:�"O�x�״IZl���5(��CV"O����K�);�"�5E�tP1�"O~T�b�H�G_~�Iu�Io��jR"O^:V��z���d��</wa!t"O���E�M���5�V�Zu���"Oj����\�Rxh��*cJ��"O��0�$G7w�𠦤(�X@%"O0u!5BAf�r�d��_(,ث�"OxT�3 �dCXrCH\�0�=�"O�(���Q�~tٷ�5���"OH����,V�
�⇩��5�8y"O�� $�E8P7�Q5J�l]��l'D��;��S�6=�fcП!�D��@�%D����C#=��i�$�ν6:`�ڧB"D����+|Ƣ4�7f�Q�V,��/ D���R�b\!:ԥ��$Fd�)��1D��B�C��x��5�"�=G`P� �=D���B��.s�2X;SfI��N�q��=D�l�S��HV(02h�%-G�t`:D���@@V�;�S2�Z>D�`s58�L-k�b�Kz  �,=D����Y�[��� !e� 	�����;D�ԸdþC"�}[��!XM �B%.;D�H�!��-�r	���U�s��$��e9D��B��&6�&d�!�Q E����6D�$�*x_���@�׮h�[�!�dh���;�J8Pg������!�S<R��dŚ�.,�(��Ux�!�݁7�=�P��O��:���cU!�d9�0�r��?���XǧվY!�DXj)$0��(Y��]�ȁJ!�DK5e��t��&Μ�]S�-G�\�!�D�\�E�����D�V���G�!�!� �R=�#�2,�p,�p�ϝ=|!�['ʤ��VJ�	v}��œ�jR!�dii�j��8��B�<!�� P�[���P�>�9�)�`����"OTd3E�A3D�`1#'9����"O���b�Y��BA�ä�� �"O�y��ċ?$�&��1*Z�'����"ORQ1c˳13�xw	X6�2)�2"Oށ3�lT;���0�÷pU��v"O2<��MdxZUs%��9��q�"O֥ �!�:��r�EO�O���Jg"O`��Q�!�P)f����Mx�"O���G�<Sl2��SeY�G�80�"OT����;K	����J*��\��"O�p�R��Y <(��S�|XD�P"OnӒk�3 �|��@��79dP��"OJ!)�' x�L�O�g� �A1"OdJ4F�5e2�d`sD؜=f([�"OB�0��0Ed�م!�3l��Y"�"OM���YxpҜ�J(:I"�3�"Ot�9W`Ù'p���たX�Mw"O��R $�VG�-�f#��I6���"O�Ӓ�KeR�r��s��u��"OJi��+ŻX. �(Q�Q�C���y�"O~��KߕxDq�gF�Hmд"O�L�'CO4]�V|!�/�6]�����"O�e)���n�ܽpn����ò"O�,��b�8T�,Kǆ",oL���"OP:��@//������%��}��']��4�
�[�Hٺ��L��ez�'�(�E+Q?azʰ96��+	� ��'��ۡ�՛ImNP�mڦ���'�jP��cT�gY�\���۩	�ҝ	�'��U(5�� Q�R�)��,[��x�'���+�B+n6b�ZF���2�T��'��=S�&�� �*����V"Ĭ���'�A0s-�3rǠ�
D��2ּ�B�'?�ABR(��a;�m*Ãͩ*V����'"l͢b��c@\��⍛/_L��'�@I�cOߕ;��Ջ�G�'&T�S
�'�x�x3�?.B`��$�q�}{�'w��\G4p�J�CEf`�DB�'���Q,E+�=�QDT��Z�'���94,ƕC�b�d�3�<e;�'�J�K���%M�r\�G%8���'9�����\;x�Qq��.{R���'mL��h��S��]J (ߘ{�iK�'������#.`x0y&d�q2���'�$٢��S�v5a쐌j����
�'��(���P�3�T�pGP\�)
�'?��HE�*?�E��������'�Xm���@��L�1���"	�'����m��j�X]f�͆ IH-��'��a��̈ ����5�C���9�'��5#�J��>`��KiAȐ��']N`&k >�d�B��t(҄@�'v�I ˄��dzm�,kH��	�' v<+��a-�l�F�cWހ��'Lm SN�<r$��h�ȅ�_H4W�<Af6t�ڠ��(M,��yją`�<Q�"�!d�:����=L*Y
�FZ_�<��2�ԁA��n�~���<�����3��x�`m��RYB�k	R�<�)Ιo�R����**�a0�[h�<ǆ*<�v�
���+&�]�<��)�q<)"H8k4&M�f�_�<9@LQ��E��T�C��}�Q�N^�<� �x�����hp�t��SR� �"O �8�J�`�Б��Î]؅8�"O6\@O6hb�z1l�9V�-t"O�pq��o�L� K��n9��"O��R���M�ʔJ�
Y��"O:肐�<th]Y"�(	ࠜ� "Or���a��nȮެ�S��)D�4��#]o8p��5�̏G�tE��%D�<ken�'8Đ|���<�|�wA/D�����'i�rL� m�yB$� /.D�x8Q�����`�D
�pQ2��6D��B��ӝA���¯���(l��G3D��F��%[76yA��Z� �(4D�t)c�" �鑁�0O��!:R�2D���m�8S�
7/���=���-D�,xS�Q4$������. �h� *D���sMƙ3�|�@Y�A������<D�x�3D�16״<भ�6��ԠI9D�����zl����G�5Nq�@��f#D����n�\:��k����#����&<D��*�DY��L����ʲP�,�'E7D��C�MԺI�=�e 	�ƦP��#D�h�G� z�N@X�%�"��0[ׇ!D�$�` �d t�@�⍮#����@!D�P�!`�!�X90��=s�`th6/>D�C!g]:���uM��W�j=z :D��I§ى,�F,�u"�.&�6�R�I8D�����څM0j���E�l�2%��b5D�\QC�J�U� �ib��2\�p�2D���AfS;\\[f�O�^fb�e$1D��3D��~�©@�����	�g/D�����C��0�ĉ��<���:-D�Ty�)��>:b�˲ɔ�.�� `��*D����I�9ym����Я@-6D�`knF=X�����f�&D�� ��2D���3��?�8���$���pS//D��b�C0�.���H��'u�|�ǭ1T�@[g"¸FT��%B��;	��"OR���g4,'M��'P�!�D�"ORmɀ��CC8)��Ɲ�?$���3"O
]�%�	�D\�q���U��i"O&�h�-s���
 e�{���2"O� 2�� ��$ꃁ^2���"O,�K�n-C")h�)ρ@bVّ"OV��'�)z>d����%}jH��"O^4��hʈeHt���;s\,��"OH����R��$"�Ҿ1BJ��"O�p�a�����͋����+�"O�1�r޷A���%bf�L ��"O yI[����d&V�3�FAA��(�ybj r�@%H��[�B����rB�)�y�� *�s�%:��c"�Y�y�ǟt���p)յ$q|��g�
�y��+� j�J	'�x��A.Q�y2+�+Xy0]qsh�?���b�8�0B�� 3@6l��W��\�-�5O�jC�	%:����c�4#�la�%Asa~C�I�V+����I�G�Q�Ȟ/+�B䉋 3���c�v��M��`�G�C�	4%�	�'-��e'`e�p�"�RC�IK�`���ą}�,�qEV34�$C�c�<\p�%F W�e�GhS���C�ɏz�n]��)��,�$��G.\UظC� �����$��SM�A;�ȕ�/��C�)� ��0���5X��AƉ!�ZI�#"OZU!dc-"�r}��V�PH�=sE"O���F�d��c�ק�c`"OhݹV*R_㰠�ga�^����"O4��o(H������1n�h��"Od��a�
�
�(�9���"y�*%��"O�qb@,�:s�t��eLr��S#"O��� U1
�@rq큧q��h��"O*TR�Ƅ*BW]Ç�]�
�<��"O(e����,y4�Y6H�GqJ�"O�9�U�^>R��8U�_"	>���"O���n��C�l��� ��-p"O��@��35ﰐ#��9�R�!"O�lH�b@-I��� ]�b?�`�6"OV]�QI�)�u� ��i��9U"O����'Q���(3I�eC��ӥ"O��"r��x� N��o=x,r�"OH�x4$	�6eB��� hI�$PW"Ob ��
�r����+8;0:]Xa"Ov�!�H
}�lL�p��j��a"O�1��.�3���9nŪ"O60jW
�'@�@i��*��#"O�����[ 5p�gуL��sB"O�1���δS'���DZ2R���`�"O���A�T[@]K�D�{�ҡ�p"Op�Q�JJ�U��0P�m�y�� �"O��9���at���gÂ1�X���"O]H')��G\�%@��$b�"O��g#I?dZ���,E,9��R3"O�}���ZkB�!*3f�t,�y�7e؞� �1O��x�R��yrCI6Y?�8���Ii�ɑ����y�H�V�m�T��0F٠�H�)��y�C_�_~�zC�J�M䤩j�+��yB�_�G���,�+}����yB�Y7ڜh���y0E)FA^/�yr�S�,��Ҟܾ�xUO�y�%�Q�h�� ��	���p楟�y�d��I���ad��X���D(��y2i@;8��"��ySH�&�y�J������Uk����R`ר�yR�ڟ!N�Is�ڪxEv��ҩU��y"��:]����>r,�ͺ�*���ymZ1K��� ��)>�V�����y�M��H���jf�!!FYǥ���yba0J�u� �҉�(ǂP3�yB���T���8�ğx�Iz�	��y�( ��|��LGܢ�!�W�y�-2P��#��$>0&ʱ���yb ��H
�	���9��$ʃ&1�yR�t���#�%K4؆)�֯��y��0B_�����(T���2���yb 'op("QNRS 	#�G+�y��0�8-��K?m�5��b٫�yҬ�%@)��#lC��@\)�`	�y���;��;0���"{pM�bW#�y��.�J�`�O��LJ�a�$N��yB"�Z�
 
��֤�酇�y����z��'�A�|�T���W�yRL�_����&�s���p�P��y"��:(�ȀҶ��<�2X�'g���yRQ"_�بd�Ȭ>܄�戁�yr:c*y�G �´�O���y�!��\�~�9��Q�}��I�D��y
� �����P/�`����R�@��L��"O��B0@B�%�b��%�� �����"O�dRW�=3nH�����?y�l��"O���E-8*pIA�W2?����"O���]#4f8!��#��p�r��S"O0�b�?z�L��C�	�Ȉ���"O,u�H@�7��$b�h�=���¥"O<p��f�c2���%D�P�(w"O�QgEؿ�R���G�Y�yq"O6�;��W~0wfV�K2P[p"O������f]�m���%G�脠�"O��#�!F_���o��}w��@�"O@MZǬ��/� ���(I�UfZ��"O�8���V�@����#@y4D�"O��$���Wu����,W�eG t
7"O�q��6|��4:TL±M=��a"OtlڃO�fȂtR�b$^1�"O��f���~�̱��GI�&ДI�"OZA��.�� хg�6i/m°"O�!L��Kc�$P��X�5�q��"O:E��9nmP�20��pڣ"O�Z���P�`'��2R�� �"O�e�B�{jp�`��1M�0�"O�t�V'L�+��0�B+kZ�у"O��W`WFnV��W˙4=�X9U"O���h�_�H���*���06"O�4G ӊLUmCM�l��"O�9�`#�y�����j
�U�P�"O�Lk�Á'����Q$�i���S"O�H3�o�1[Vd��2{��Ha�"O�;�ď�Ae�dP5NG�-���5"OF���oU3l���읗Q�T��y�e-����]�X%|e�I���yR���zx>Ř��T�@{�Ls�C �y�+�91>���B0�D�cZ<�ybOŚ:�еx�ȯ
ɸHA�3�y��	
>���+�1s�t�k��E��yb��9/@N0�� ȃn+���#�-�y2K�2(��tQ@$���� 0dL1�y��4���� }
�����yb�	�r���I�e�1�斗�yBD�R��(D���Za����o�;�y�F��� ��� Z2ze�$$\��y���!M�%y!˛U\he8$�Z��yB�O�2s0Lx���\M��z�-ˢ�yr��U��1�E�P�`d��F�y≊8�ةC�[<Q��ْ��y�@�$��wM��p{�a��y�
N~�deM�d�Ҥ�ąת�y��>&P�kG�[��%�dF�y%��L%B$�P���Y�(%�Ӣ���y�^�^�mg�"�~1����ym��)�llH��")>II2Ƀ�yB�Ez�� ޝ��E�M��yRO[��*5�`S�rqǇ��y��ٌ�$�����i�5�y��Og��A�ŊA��%�M�y��o��QV��!u�r�J�jА'�!�G�ph�U�F<o�YJriN�!�$�	�2���R������Ww!򤋸K�,�2��Y%t�<�@R�*?Y!򄒧� |�@��0*���ȇi[A !�	�\`�{Ć݉k_42��!�$#~�v=�'�{ 4�MJ��!�� �6�v�4�{�`�)U��5�D"Oܸ��MT�˸)�2�2.�n4B$"Oб�����{��ٶ��=�zZ�"OPXH�ǋl�y��놙n�h�C�"O& u�J_}��S`�
:H�����"O䁂�$�<fn��:7� �8��D"O�ēE�ȦE)D���͏:o|Hg"O�eѐ��F	A5�
� @��B"OHH*�)�\Ѣ9h$H�΅D�!���phB͚\g�Ģ�N�8�!�E�D��@D�8HvQ�E#Z��!�d��g�Ձ/�6l���HD��B�!�ą<b"����I!h�*ԩwA�!�ɚ�h��bV*�v�P��ԇ"~!򤗖���f扥FP<݈�茷c!�� �i��ŐF�A#$4��rv�զj&!���r#��(�3w�Ƞ��ǝ!��/vВ��f4$���*�f�'!�+ٌ�X��.%�\��R�E�7!�P*i�����gI(u�Q�5A�!��R�Vpe��fӾ����N�!�T&���#� Ud���8���5�!��F)j}�t	8kS:TB�ݸr�!���}���]��Y2͠%w!��{ɮtqn)M��2��<?!�$[�'St|��f_33Մ�b�N�>!�Ć�^5�m�%ET3d!�e�L�90!��'E�Uғ��,x/d�qKîa!�DǙTn
5F��O(�dx0�!�D�=<= A��rt���fE_�F!���N�>XJr��$Dh4�$&� �!��i�+Ş(n����fcN��x�ȓ:�L2Peڦp�	 �KN8�Tt��+�\Ԃ�ア��������b���1rΈ�U�� ��Wŗ�dy���]2@ c� ,hF�kVb[
L썇�#g<�B�ɣJ��qk`���FH��8ט�`�������"��j����ȓ��b����V��A�A�0�N�ȓS��T	��T��l�[gZ9
��#6�X�`�N��ǫ��N���ȓ`�N��c�?W�jH���ۮ��,�ȓ1�D$s"�)
fx!��� ˆ���Y�]��
-C��dA4Z;�Y��`mfi���*'J��䤕0�
�ȓgq�6a��X� N*8s�U�ȓ*��m0�%V f�:�J���)�Tx��~*t�)'�S\��!�*����ȓ+z���oE'9���2U�^ @�Tm��FP��B��~�b�"`
�N�����&�)��GY�d4��C\*I����OذQ@����"��� ��`�����G"��*��0N_����W�.�-�ȓmw�HyL6F�N�cJfd�ȓd'���A��2��򪗗4o���9"���d��6�$��+ݑ)���ȓ4J��C��>j8ʸ���Ҵq�ԅȓ%�xSX#�����i�ȓ%��(�<�����WRy�ȓ>Y�Pj[�r�	�q@S�t�ȓ;�Q1,��
�
k�nزP��ȓE�E���6N��l;�Kī\�����O�h��K��Nk�!�֤��h�:<�ȓXkf��g�;iP0ؒB(A,&�t��S�? ��3��\'}zvdxE
�e���Q"O8���EE$�x̱t�k���[�"OX#�C��H�b�@-˦��]pS"O��z�K�3��XT�U����w"O:�8���
:�ܨ���Y�c��"O�i����2�*Y)ዏW�t�"O�!kBݻH���̕	O��&"OD���Ea&��8��;E�°"Oڀ�Ƣ<>��X�U�]*b�t5P"Oʹ{2���`�����������x�"O\��� M����P�Y�\�R"O�}�$!pO���%׊�"On�ǩU?�䔣`�I�L��̡�"O��8�D��c�0Y�&B��~�.��w"Of�ؓD�B?$P0@ěI�NH�5"O2X�s�Rn~��n����f"O�\a�l�6> �<y#W"O���I�?���Ak�zӞQ��"O���pk� �x!`ʒ8Z��sd"O�\��dJ�6ބd�!Î]B���"OL���×s�|���u;X|�""O(���OD-���j��!�T{�"O�1iD��>�q���x)8t�R"O��أOQ��Ȕ�GeWw~� h�"O>4�A�� �����x�3lJ��y��S�>/hҒƝ; $�%�"��"�y¢���D���&?ƍY�ŋ�yrD�.>È�B�)V�^�hQfjE�yr$Q,�ɰ2� Y�DyL��y"��U(n���\�~P������yĒ�=  �8E� �C'@x���ܿ�y�ǅ5�]����80��6E��yR�� j+(ԨV�Y,�^a�$MZ�yҥ��uܽ��؇"o2���J���y�4��pP�Óm\���y�pl��2h���������y�)¹d4Ex��Y��X� SH���y��)K#}��\I���;�N��y�)�͜tA���@	:@b�%�y��6F����FM
9-���B��y�bȣ1~N��ӹ-;�,�G��y�$�"XJ�!sq�,�� ��E��yB��1�����*��"���H�#�y�.�y�������&��b�9�yb�Қ?;* ���`�\󂈛�yR������aD	u��d�R���y�EHT�����6@#��ٻ�y�◞[��S�K4hx"x"mS9�y���*	�1{Ga�f�������y�!L3?���Do@'X�ȌC�"�yb�}`"i��*U�P�<�����y%�ؼ�g�H	S�&u����?�y�ϭ(��h3���D?¸���y��Y�%\̓�g�5Q(ujSo��y���#l�BS!n2w��q�EC��y�fӻWC� ��3h9�(c�W��yB��r���ǆ�f�x�@%I9�y�g�#X܄`Q� ��haHM����y��8�D�pЃ��`5�B�B��y���<���2P0��`AmA#�y��2s|ec�<@��@���yJ��_K���E�.������>�y���^ P����3�"�p-��y2&KafZ��J�23�����֑�y
� 6X�H<8.ZQA����T���4"O��EN�M҈��v�֛R!�!H�"O,u���0HQ�q���;5B�#�"O����I��!JrN��@(�U��"Oqh!�$eB-�vL��h	�Ĭ[�<a3Y2-�o#c��xw���ybfG�����I0M��vm\��y2�֪!xJ��8{��� �@���y��A%Q����t��vE�qD J��yL��T�� �q	�4�S�K$�y��R� 9�4K�%d}��HBm7�y�℩R�	a#���H�V��a͉%�y�聧>Kԓ"���-��� !��y��"^�P u�ڂpj�Ѳ-��y�`��"���'�hSx䱒I���y�l�@|LP�U��3d�Zb`��yR�F�GU���V숇ae�,�����y�i?0B%2q�^��D$�ꁹ�y�`��,q���S��:�� ����y"�r-��(�BE��}�$��y�'N�P=^9Y"���V?L=�3�W6�y¡��U�h(�o^ Ѥ�a�O �y"[/72�9�b�	�:L�^*�y��4=����#�Z VҬ�'O��y��%
�����g Os�,֭��yL�"�|����_@s2豆œ�ybÓ�M�^���gɺc��9W 
�y�@
4G��3ХȵF~Y��͉�y��S �N�sӂE/y�䕢a�_"�yB�&
]r��U�ٗj�ܱ�NT:�y��5�2��ŏܓ_�"�$D�y���cՎ�I�/"�H!�bI�.�y��6�$	� 7��Q��ه�yB�1p����E֊dێ�s$���y�(�3'jK7��%�r}��e��y!T�h1@��#U�i������Ȇ�y'��0���P�O�x���!��yR�O�p�9�>q�����P��y�'�1="|bDG7lI&YC`�^��y�V������� /��ěG���yb�Zz�!P�l��ok�M)�$���y�A�0k��#D%��h��
�蜻�y��_Tp-����>c](1s�R�yBd�_���lU`!L�	�
��yɄLҘ �R��/)��a$��y"&L�E�v�IC�� Mi��a�AE�y�.^�v� C��t��*�K��yb�L�N�J�����e�2�&ϝ�y�^��� 6�c����S)�y��`h
b��]���o٣�y�%O<Jp�M�r�4kQ̏�y�&8�6d�#s�����К�yBn�3T%cO�e�*���C��y�g��V���%�*����H��y���,"�rDHD����)� ��y�O]VpI���2���g���yr G*B�~t
�KP��$��Z(�yΌ+�]�S�$6�r%��y�E�>.x���Ĝ�H�p!�Q���yR+Q�'�1���[3NRj=��J>�yRGնL����qKX�vK�����yhrQZ��I]�d���3F���y�ˤM{Q��RE5���5�˿�y��Z�}���j@��Ak�	π�y
� Tm�6$!ȱ�E���E�B�ڠ"O�u�tb�e��H�O�z��"OL�(@����yzvdG�
�Fm:�"O5R�UG�8�b�ɬ�Z�K�"OP�x���Q3���.4�E��"OZ%����Sd���]P��9�"O�a�0S�&$
�3Qw�u"O���`䊩����-	�@�w"O$���!���PeV�Q�JE"O�4d��M�@�Ɓ�=b��%��"OB��v��P��T*�6Y�be�w"OP��w.x���t�V @f�A�"O`�#3�P� CNL���U��16"O�h�ǌ�K}Z��2�;؁&"OV��"��hc�@��-��@f�y�"Ol㣔6m��p���Μ-%,���"O��!S�F��T��Ŏ�[�>M��"Or=��M�${��|��k;fm�"O,xHGGK�J]Ǡb9d�!"O@��"�r�dc� BC�E�"Ov)�c�C���D����-�4��"O�4�Ј\[�všf���N8�"O
ͣ�-K�
@���
#`�d�[t"O6���Cмc��Q��;	��pз"O$�C6�ʪ`B��e�,/ߠ��"O60{am9���S��n����"O�T#��A� xx0V��KA�X�"OTy[�I��O�йQ����y�"O�i�@�(�L#Yayc _��yR$͑gRExV,O�\ &��O���y�"�cԬ� ��2Q*=��e��y��D;V���	JO "`�Q��y2�R2RHh[-��W�(��	�y�Ǔ�V�>�!����JDm+g��)�y�hyaa�ΚU�}R1c�
3",H�
�'bA��
>(͒㠉�.�t��'M�	7��~|�bXw���'c��2mҧ���qk���y�A×�b�#A-�(�V(�pL��y"$�'k.�o@3VDA)��B/�y�ǂ�vMԵ�V�S+IR�u{"%ڳ�y�G�T�ęb��70�x����۲�y�,��w�8��g�֥&N�53�ӏ�y�e�/[���F���r7�@	����y"BE>L&��4�?���E��:�yb ���b��2͓E	���ꝡ�y2☂ÀIؖJO�6�,Y"����y�j�� �S5j��}&rr���y��%(��жB�q?B�+֠�5�y�O������=mA��2u�Z�yRI9G
1r����b�Z8����y��R(�kD�߰F��q�ra��y҅!"J���S�O8����ҏ�y��w�B�8�Ұz@�L����yr�І&>�݉�CT�y�n�U(�6�y�� 5Yu��k[?A` �^0�ybdY�W�j���<9{�h��m ��y�Qmbj���ɨ_4`�"���yE��	m� �h�QC�L��� �yRM��K*[�ҸI(x��B��y�	�C��T���a0�8�k���y��8P��h�bJ�|<�h���yr�Q���D�M$oyn	P᥅�yR�\�0\���� A�H`@����y
� @P�+��6�<���/ɥL��ͳ$"OU�2��2�,9F���T�Tp"O��jd�B�f~V��m�+_튕��"O^��bA�!o�����lN�?��t� "Oڬ�E�݃q�PIڌn���Z "O��95h����щM8x���X1"OL8�1Βm����qJ� z.X��"O�M�G�^�;Q�M붨M�^	�""O�H�d O=����4�	9X�^�B"O��`E�(�8�x1�?I>�P�"O ��鞀-�NY�c��� �6�ȵ"O�[�#�A�f�BV��#>{,ɢ�"O2���F؞
ܢ���B��gd]��"OB�ࢯ^��P���!��$U��$"Oy����
�J�M�y���yrm�R�h����A��P;բ��y��@
�(B�a�1�L�yBk>"� �P%Ըm�2ab��y���X�PfŜ[T��e�:�y��W�H��]�"%ԗ8��������yB*F8f���
D�2��! ME��y"$�.zK~|���K�(ܐ���ޔ�y�猗<:���h�,N�.Y��&��y��ɱ6y ]���F(D�N���W��yr�]�t�����,>�` �/K&�y�����"�gũ5l��D$Y��y��72� '��4 K��$�y��P�tmRM�-Z���˷i��y2%5UL�-���EZ��b����yA�?M�6|��dIu���Չ���yr,KY9�i+@ꚚoA� ��`�#�y��A�1<f�ǎ��b#�i�  ��y�+ν(�,�2���F}j�sP�'�y"��T�3�!?�L''J�y�F�,¼<Ғ"O�7<hTR3��4�y�+Ǔ"�R���)��Ed�s�"S��y� HZjV�*�G�9�Hg�T��y������%:�����,Mmad���';6	��(� FvX}�b�Qj�I	�'K�����݈[��ʤ�J1l��' �ܰ���V*�=��HX2Keta�'>8���!�N��,R;0e8���'�$e�E }�V�ɵ�20��d:�'���� �q�¼�H��+MXh�'�ʄ�X�cZ<I
�������J�'�͐���8"�h��9c�'����h٫ �h�b� |9�@
�'��(P�MX����E�5n�T��	�'�� ��,�v���m[_u�1��'�F�c5cK�=�LD��U����'Dt��ܔD8�qde��O�Q��')��f������:�P98�0�'�J��6$�-N�.=���԰,�P���'���Ȑ!�)p��"G\"��'�*1
�
ө2/�4゠�i�� �'�+�:L
h����� ?�2Ȃ�2D�1��M?X!a�ܝu�q*")$D�D��D$Dl���E�?�Mץ D��ǡ�&�:��D#��\�(�C>D�ty ��[f�(J#�~R���
0D�$��Mi���x����q,�A�E)D�����ߡ�bt���I+N)qL&D����a*{Z)�cE;|��l�D�0D�C�#X�]R����x3�0D�� ��BP��8-3hA#�a���p"O��9�#ħ^��$h�OI^Bʔ"OZ���
=�$�� �"L(��S�*O�,�E��@��K�b������'��%���J�&u���6�»��	�'��uC☰lyά����w��2	�'?D�[a���*!#$�]�pz4Y+�'!z�x�b� o��K�]�N<��'�Z�I���B5Y�[5HKlH��'��(��,GG�����l�����'o0�2�U�<���x�iǘsy�(��'�>�2�*J6yOH�@5%U�6b�q�'� �P�B��X�����&�T���'��jR�ߏ���3�]9U:5@�'��PA��S�MP��h&���"�3�'���0����8���&$8H��'��Xa������V��6]��'\vM�zN�Ivi�+�@��'��U c��uTCuF�A�\��'�H���̋�@�`�Kn5H�池�'P��� �I}lyঊ��Oè�z	�'�Z�ǁ�-�X�&�ϼDr��	�'� �R׮H��
��� >^%�	�'�����ge��"�I50���!�'7�Ջ��B�Gj��SoUm����'��u0d ��r!�ip���H�����'y<zR͑��f���?���B�'�,��gG�}��ѐn�D��	"�')�lK!��������KA4v>D*�'�<eI�������I!MԀͣ�'|���L
v�6E�f�D�m7� ��'y`�ǣ�AG������X�h�X�'}Fm	��FJ�{���<�H�3�'�ȕ⍗;��H�DHQ�<��U	�'|*3"Ã�!��h�d.D�<��	�'i�Pr"�]$����1�r
�'�Z,�qE��f� ���!�|$b�'�l���U4����e�I�n��'��8� �.Da�uLeM��'��b%�B�v�:�)tA�n��'�"-�`�KtT�qXC�T7W��8�'��iߚ�ނ=�"O�\< �'֜)knb�=�d�t��'V�]�I�lX�貅��`ɦ���'�䉴�T�e�)"�F!`l�	
�'��q���S�"����]c���	�'	�}H%k���'
�a�����'v!�Pe��"K7��S:�Ւ�'N��CV�P�b��)�f�E� �ȓ96PxA�^f���H�;����O�T1���#Sn��5B׶L�\Ѕ�#
<�16N�?⤈:4#��)�n܄ȓ%�5{�B�4pd���Bjϸ!���ȓy�hZ�mɬU~8#A�ʲ?����9�ԑRG�=H�* �3[�M�ȓc��������NspP�D�d?�x�ȓ]i, ��WŸ1̇�Z)�Յȓ�"�z������࣒G��V�ԅ�1� ��#׷~�`�EOp�u��'A�#S��@GR�;��V�/����<�>ᐦ؛7�ԣ���(ɒ��ȓ.���)�kH�_�`�k�+�"D}VU��C�ހ���R"�����Z�H�x�ȓĀ��I�?~T�"��c�a��S�? �U��A`����
ã@���"O�1�ܢe���� ۆ"�!j"O�a�׏S�T��L�ƮU-L��!"O�@1Rn6p�"yS�]��2�+"OB !�E�o@npbTc�,�� Ò"O���&46���#֡�8y���
�"O�БU���|�L5o�*	�:��+:D�`:b`�xf29�s�Z�bw��	e$.D�4x�+W��, �K��P�U�!D��"�"
L�ڀA��*�P�I5D���R*�����d��Z
��a�3D���f�0�l6��6�UZ��c�<rjQ;+��mrQ��+#��y�e�h�<�f*u�>	j4-*_T�l��
Dh�<AR@ޝS+Z��Щs�Zm�MLe�<���Z<N����&�`%�-y�<���3�����]��ȰtQ�<9jK�{�\2�$p�8A(�M}�<q7o�
]�pӐ�W�B�����Od�<�!�__|��K��w�㱀[�<��k�~�jP)��(��'�JV�<i�/�/)M:�X���$AfA��U�<��`w��iG�\�E)�C h�O�<�BJB#7�A�Ďم�L��R.UO�<I�A�$��qGA� 6ԋ���_�<	�+˿<����_�26D@MH_�<�U�H#"�6����eBz��7��O�<�S�B^�M�p�Җ9�ly�i�J�<��M�z�0��M�a�`Be��k�<餆X�T'�8;Pa�#T�����	h�<!�$��,�v!"Cm\�9d��ص�l�<)����b(e�ǘa�ڥ v��<17IX4U��x�M��{�hS�x�<Sm��UY܅���?(�,��E~�<iA�ڧ W2��1���4�0Y���O�<I�	�/���!�"-2aYR��O�<f+��c԰ ����	Z��a�L�<)j�V��M�C 	Pl�q��K�<�&3q���R��\� �O�q�<AҌ	#kb��!
�O[`%��cFm�< ��szz� RK��(��u��c�g�<1t��l�\0w��".p�{4�`�<)pE��f�(sH�1Ld����TZ�<�hK>xu�t����]m��r�_K�<х��j.��h�ɕI$��&˕F�<�*�*�TYD�ãK�L��,D�@�F,ϴ<��� �����&D�K�ޅ����cD�6�� �Q+!�Od��M�EϬj�^��L}�h����E�<)�яB'E�U��*+
M1`�3D�t�R�� i��%�d��	n1D��i�AQ�&%"D	�����׀-D�Hɑ(�Vۼ�h��ȭ'���#�i)D�t;��Y2;���6���$D�Ԩs,�\W�(qq��gM�]p�E"D�H�ѭ��x��)��Z�Y��#5D��##d�"$�Q�O�^	؈؁4D�@H%dȣpLt��ƈ#���7D�Y��J,V&~�I�I�V��B�`5D�\�@� �E�b�W��x� ��*6D��� �G�,P�F�̨(��]���4D��zR��y��i����y�y��4D��Q�6X���y�EL9 A�ux�j4D��R+�0&��·l)(� ���=D�� ��q7"R&_|����@�\�b"OŹ��K5�E��E�m�.��u�iJ�'A�)��|¤:Eg��ˢ!����B�����O�㞼�O\j�(D�|�@�� ��7���'Xr�!r%B=��5����+�NX�	�'����̔J>�b�����j���'�~����C� �h�!2��x�0�_|�<iǋ4%��������ޘ�6�T�<I@Ǌ6||Ը9�N3	��K�x�<��o�� �ӄs�:MI�C�[�<A�+ŵ^	 -�V��'}Ԉ���L��p=Q O�+�+'қ��Tj��EE�<A��[�5� �!gh�0:(�iF�<iѩ�2w�ȼҶ�+I�X�Q &IE���0=������U��Kǁf~�X�#cA�<��d�#.�iz� �s���r��V}��)�'��e�ЃL�mL�A��f"�ȓ%���r�];��E	ɳ(ϰC剰��WFM�������'xBB�;��1�'^$:��h`��$6�B�I!���BG�'$��1�&lSA$�y��I�7����UE)E��-��H#��C�	'��󔅒�+��z���r
B�	Yc����

\�q,�%W�C�	-F�`A�G�0g�b�	�@!n�B��n���%��Q�*
6�Z�p��B�	�B��%E�`� �?�R%��&/D�8��X� ����u�A-F]�])�e������'�����9"�H�c`L#�=
�#D� k%`M�'=Ba�ࠍ�Dx�cc�}��O��S�3�M�}�A,IrȀk���9;�!�䏏5�d�v�ȓl��R��X�!�`�<���aW	3k��A5�Y��!�ϳ	J|e��(AexD�X)q�!���7ѤmRě "N"Y9����C�ɈC58F�!4(����<^C�	fT�Hd/E=�D�@�I�+�dC�	�U�P!�A�n�p�������B�	�#�*��2HPVp(��?��B�ɴ0g����ˍ~�dl�BU�w$�B��<$Δmu�YI:,�%S�I�vB�IUe��(@��lS\<s@H\�z@&B��t
0K��\*�
���ٸC��B�	/1�bp�ҁ�����n�`��B�	�uI�q(�#��,��šَ/�NB� ,Z<r3*J�A����#��?�JB�I�eR��{a?~E��@=(�B�I�U��Pڤō D�`�g-y�B�I�j�|��7�O���Ц�\�DB�	��d�ڒh� ��Q��I�
B�<�>=����{L A�%@(w��B�	�� ��C�X ��P�����^C�	�:��A�8$���!gݢ`�2C�I�P&�p���@C�T3�<`�B�	�dXpm:�E�7/�r����	YtC�I�oZU�,O��T[�c�&5"�B䉦/����̟85��s7׺x	C�ɶl֦��7DS5� �U�E�C�jՈ��b�Z�^�K��Q$6�B�ɺ?�\�3��] '$Pm��J��jB䉸�my �V�h�0�{���ev�C�	u�FA�E̳o��Ъg�6S�<C�I$����:�v�St(��[� C��CS���N�;+��4�"�'�%"O� ^��vȘ�^�,QVcӟj)��Q"O�͂4���wX���hZ�Z�,y�"O��{VkھMB���D�u:����"O=!Q�gg�$�禀2I:�8�f"OL�3c��P�F
DTu��"Oz�P�H��I(�,C�IQ e\�Ы�"OL17�9p6p��Nu9D��"O"p�"�ӺT�]�lA�-`(�"O�!����c��A�Q�X7AH,D"O8��cnGR�V�h��=5��X�u"O���fԯ:��|��!�
 0P"O�h����<�8��M<AO���s"O�Dҁ��`�t� 4'�:�b݀a"O<!Ai�;	��A�s�h�W"O"L��@��D��
7���� ۣ"Of�%f ��r�k'A�8_4zp�b"O���hӍ�.%��P+H�t6"O�l@T�W�h3HU�&���9(��""O�����г>,�<`#%. D`�"O<�jTb�a`���C��H�j"O>�z��'|�Θ�`MH�]��@c"O� ��&/c-�y
s�8ax8h��"O9��i�EXcBn��H8B	�'�~�Q5e=�� ҧ�K�g�
�'�-���^�t�ʱ�扥,�Z@
�'��#�I��V�6��I�;k�ec	�'�6i8�W�h5Fd�iz�	�'�`��I>_=��` Z�u}b�@�'��DkR��"�� �V��>U@y�'�@q[ ����8��Ht�h�'��y�O^Y�y)�k �I��ȸ�'S��"S���h��СZ�6)�42�'��M�dL�5�H��D�G�x.t��'�0��\�3�$8�	��q�Z!��'��I�o�=B\��k�c�Ԁ��'Bl$4 �2 ��1�v�B.Y��I�'[�\9��r����L؀q�,QҎ8D�D��jT'I�Ĭ�GלA�<u!��6D�d���,!��-��U�&�� 0D�t�@	��
�A�U�(9!��/D��R���I6`�iь�~��7h3D� k�,�6/��IX$݇p2
��#B3D��*u�OR
lh6N� ��1D�p ��P:;��!dM֊ud,x�B4D��{Q�I51�z�3v�Sg<�q���%D��IF�M�)�h<�􍆗P�A�$.D������P��'�#g��H# D��q.�%|2�T��lĂm��eІ->D�䱲
D�z�,qqGFC��y7�7D�L��FP8e��T1fX5����(D��;��.y2�Q�ܣm��362D������4%SriM'%�(��f�5D�ȑ@���)�}!�dM�W�<�I1�3D�8�2-����pS�	L�OhdJ�j3D��qW�;k=��!!m	��4@���1D�`�sU++���"Ǧe���r"�-D��&��}3 Ʌ�m�Ʃ��&D��c-$9\�p�u�Ȭ~&�d�C�$D����ƒ5ɜ��:2�H:�EC�9!�$�y������f,xUAe%�!�S�S�����*v�h9;�c�v$!��R)c�������aM ��$�
l!�
�I��1��rE��{��h!�DK�hY�$Z�'���P\+�]�x�!�� ���U䐳a� �[��$r9l���"O,��N��N���J*/���"O�J��?���
W?~��l*7"O|�T�ʓj(X2�
�����"O4|� $O`f|P�/
��^�Y&"OFH�㊔G�q�����H:P��"O��	A�Id�R\ 2yc�"O"L��͚wj`@�����n.:��"O�a��IwX��p�(<2&���"OX������	g�$8�Q��"O�a ."Z�u� �6�9
$"O���&_�f��}D���a�
TS�"OHJ�� m����-�&f2fj'"OL�� SRîH6��5v�Q $"O"�Z�.7�N�pƪ[�l� �"O�l�r�R�;OҌ����7�ҕP�"Op<�F��%.$uhQ!ڐ��oKb#�'�
,����<7��̱�(��c�L��	�'I��OKCȊ����V�e�(,	�'3R���	��r�ܯT�<1)	�'��+��ݛ%�����2IHz���'
��(^�xƂ�c��VN��P�'�`Dڤ���_T�P	���K�bdp�'��D�u��2/��+/ĭ9�(�B�'�P4�%�Hf�R�H��ݾ6C,5i�'�KB9w0)@�5ϒ|!&�Y�<A�ʂ�UFB�ȠFF� >���,^]�<�0�C�{P�J&��2X���KG�<�0���}���WkH�~�k���|�<��mj�9e��;�as�*D��`�a����0��2�����+D����e[�&�nYSp�$]V�@t&D�L10�V(�ts�ͥvP4��s�)D����a6j(6�ѵ,�1n��0G�3D�� ��n���6'�	q��d�Q�0D� �n֛�La`Uf&�ظs��.D���C�}|N�rЉ�d��B��,D�\0�M��:s�ʉ'��;!�-D�%kU.~?�h!��˲�8kS�+D��;gB"a�
툷���,D�lIb℔sv��D�ĉk�l���-D�\��"sIke�ǆ)X��5�I=�!��Dj0���=~�E���)z!�ޔ7��J�EW8"�"�w��~!�$_-1��Q�%��h{���ie!�P�`�dY���^|b� �p�׽Y!�C7X�L�abH�.hX�!�D�Z!��u:Izbɉ�:Xf�AF���!�ܣ.����sDһrB�$�#Ǆ�!�D�$Z2�9b��:DnpB�C�!�D"�|�3�R�'F�@�a!��.�di���Ar/����L�J�!�L�g����i����4)�"��3�!���� �7LE�Z�$|�f�zE��dI���! $-T8P����ò�y��!F B#�88	Bt���yR�V�f;�8�M��i��@�H���=�$-���-P�� ��EL"?L��R��#�.�"�"Oܨ�G�ii�0�ό �-b��ď��!z��M*~'Zy ��1�!6�aS�f�ujt}�UJ��Tu��D�15�
�E�9
��[ҭK<9r2A8���r]"��j@x?���"��/����;�b�2R�q�Mj����2��م�	D��`��V��)����WlZ���T�\�|�W �"��Y�����djˮvR��@̑��(O��;�n����X���*���ӗ�	�g���3m#h?^6�ŕNP��k�l~�� �%����K�8\ʵ��Js
�����>U$u�DJ��]za|@M+}$ zvʐ��h䓂��Mc� �C�@����O�i�7�@U
�@\w��$p�cx^�]λ3O�T�1i >8���[�A^3d0�ȓP�0)� ڐ�KѠۏ3���A�]�b�b���xc�P�W���8�Hڴ�v��s�Q*��P�W���y��QM+�O 8A��Lo�4�r+Tdl�HR�J�7.dQ:��_�*�\� �Ə&��Y[�v���S��O����d�7j)VOA{�Lɿ�2�!�� /\����$���+f��F�bl���t���Z;e�|�#aj�i�:1��N'r�{p�׿����&CS����0bW}~�m��#���%�$����R��}QT�@%�4N|�>L��*T�)�d��u�ȡ+F+��^��X:9@ ��s�����t?b��s)��e��p	��yG�Q��O�$#�0I�$�3
ÓO�����fW�%H��!T!?S������bf�ʑ�?:J�CŚ�L���ش_7V��G©@}�HK��_�p�@����G�FQ}8��C�	�lP�4�To(�z+5�,���Dt�a#P�ͷ7��(�&Hg�>b^����F&��b�Al�3N����-�%7���ӌ��?9�T�w�6Q�ʝ
)b�8K�(Ե�8]0���\�O�
�Z�b�����A^&	��i�;.�xX�rj[� �
X�`M�2�pa�I%)��qX2A�K�t`����\�R*ۆ!� D�ĀL�7��I��|�{�G_T��8hE�E9#Q��ɿ&y��i�Y�@-:	*����D�J�E6�R��9FhP� I4a�.��6�1rԀ�lZk*u��PԶ@
�Zp�'�D)����k����GL��|��M<	 �ϙ���'���
Y�Mӣ �s���20��n���n�����H�^Ԫ�KM���=��k�i���("'T�/�����Tں�9��O�tY�E�n!��޴r��h�G)��<��M���ӖSEfEjpF�1V+����X�_�#?9���(��i�(\�����@�~$��i@0�ؑA��hx1�f��O5N�bPbѳ���	�g+ P�g��X�zm*o+/t�I|T�UZ�����Y
	U1�$��%g�	�1ٓD
�m��k]�YtH�c�ݒ�M`��%	h����+rK�K��$܀^�^����R$��A�Ǵ [�	��K�;-�,Q�Q���4zD�e\ \�J��̓$盆Æ�j	��C�
^BU�f�@��z4�t�D��f8�`��k��yb���h$�0��4|j���?�Q� G�j%�d`�V٦e�S'�"%/��'{z�YR�R�8��'X:�N�|��|���K�0cd�JU�؇6�����⌼Yu.�B��'�t�j���,���.E>**�Z�+�+.�f����-�P����R�������>X�����,$�b���*-�r��%(�>��L�>�y	��ˉ8*N)�hCǦ�+��1)-�i1�'�q�Pi�9uz(�;mYB��
�*F0|B���&�\�d��Fg2�#-�!$}� a�On�q4��8��z�!R���O��8e�-�� �O�R��Q��HH
P�R<�b*%�Ll15��M���E-D�.��-Hڴ,�h9�@�Q���=�2Lج�t2B^������*��Ɇ�!f0du
e�˱b����т�E�0kD�z�a�*ۮ%���@w�N,o��fJQ�Ճ� 5�6��-���wh ��M &z$�If$F�o������7e�� �<�0B�A�2�^@q#@ѤRv�����"< �����)e�ǟh�j�ガ�qO��Q6��Y�bT��RzQ��*ʹ7��, ���1J�/KaĨ��s�6�p��(�&��fnS�a�;$V	*V"\�<2�S�,Kf\�ȓ2@hJ��r֮�5�`@2P�a��'&$&�I4(�nYx�X~���O6�I��օ6K�	�p1��"5���l��K��<$��c�'D�!V�A�n��]>��^�&�8}'hFB7���!_8�=cZ0y g��@3��GyReD�F���G��IUvAۤgH�ް=3�J.i������x��ٹ�M�T�>0�ȗ	'�VA���'���PůCCX��`b+�&��(1�N�>n�@%(-D�p� �X�,�a�폍XM� ��g(D��%�V>��#-�5.x0�p!�)D�@(r�/I����jj�<]r �&D��1���0w~���DGA;GbF@Q��3D����b��. �<����
�d�,D�ܸ�(�� ��g�9
R2�S�*D���c,�%ؾy�$d˨Grz���=D���"e;��O�vH (a�=D�t�؈�ny�V��Q
�p�#�x�<���G1R�܌�w�C��.�I6��Q�<9� V�����A�V�a�I�E�<iCԀzB�LZ�.�6K�ޜ	��B�<Ap�Q.)��4.�K~x��/[~�<1�� ��t��Vg�R�� �f�`�<��L�a�e�`e��1�'��;���n��	Q�@Q�$����':L�sC�1DU����'���'(��`@3wD�S�T�� ���'�4�d��L�l}�"E*vN���'o��&OJv�Z���鍹�:`���� �!#�*�g�j\�M�G����"O�]��$���>�ӆ��}p��"O�`���K��W�C/B<��ّ"O�xʓ&�0>$D%�� Z (^���d"O��§X	c�d�!��:V��@"O�27��J��B6  �M�:E"O�����E�L�PBa#q8�ڶ"OxL����E�t�zT��J:��j3"O����+��eA�BT�ZD"O�!9�HyTN㴀O�wm[e"O� R���_�a�O��<�J�"OT�J��M�X��`�FU?74&���"O��Д0[��t�7��� �(D���#��=+ɞ����P���$D�Tkq�S�v(��,C��4kǅ>D���r`�;���E��+Ai�XP�':D��`��8���ܣZ �wJ:D��I�}��]@2��+�$�[։8D��x�iZ�੩2�VH�pp��G9D� SS$�::
��1X�9`Pa�	Z�!�$��^p]AQCD
k��tǟ?:!��3M�p"����AQ e����6>l!���R�+�<��� ,޹�^�*�''���&4J/&�s��J�p��}:�'>:��4X-���F/]$>�����'`�%�c@ջF|�5mO>.`�1��'\���7����-�Ua��$�T���'��CEUP0՛ahU� ���)	�'�r���\85�Z��Ļ 
*�S	�'���D�ʮw�:X��؈�ruP	�'�`�r6͜U��hqw���'��	Ŭ/?������L�X��'�q�sI�-������y��9��'L���FM�0K$������rI�e�'� �c��%lMH:�.}ঐ��'j�[Q�Q�Tj:I�G�Z5]M��:�'�@-a'@�q>���&D�KO�!s�'ZMx!���VI�dǫ��Ap��[�'�  B�P�Xب�Ȍ�(s��
�'�Й�lҬ;[ ��3N٭ŖD�	�'�&��n��]hD�m�]^�	�'�|�ݜ<��q�BF'IԆ�S	�'���&̒fB~e��*�D��`��'�)�DZ�*m�����ĉT�2�A�'�T��@@�k��K�h����'�.���,϶e�A��H�
�Z՚�'��h��ը4���� ���PZ�Y�'�bE�S!X�qqM2pb�yഄr�'� ��AjہkRE�wcF1hIL�
�'u`��Gfv�����(e�~�r�'�2�򕩂�l���p +V^$�@
�'��@��ݜ6R�����bز���'zHTʖ��*G�9��(��_qnm��'d*i����4n�h��łɝU&X`*�'p�� ��Ǽ �Y��!Y�֌�
�')��3�o�e���TI�	�m��'|b����R�m�ȠcU�ɶ����'�^�t�e>p��q�C3�<x�'�pEr���rs.y���R�blY�'�h�`$����*!������'Ů��t%P�l��M�У�?����'��@�e���(y`(�5
���j�'�(��6k��QѪ��T�T(��'��	P��4N\0{��K�xy��
��� b��d�N9P� ���͒�B���u"O
M��k\�K���(���=H�
�x�"O�Ÿu�ͰVvpYƭ�Q�z(h�"O,��s��5M�@eɳk��N��X"O#O[�-���J�*'o�4��"O&�r e��M�*��V�3`~��Ia"O��	U�ӑE�P� 0ǔ�����"Of��#�%p������\��.�"O串U��y�$�s��>F�D�Q�"O��ɷk�`�0P��� Hհi��"O�X�-ǃI ����h� �v� "O4i	$L��RD�s���sIf@��"O�Ð��L�"e�a2l�"OD�i��>-�R�)�]=A����"O(���m��8"sJNP�(	��"O�؉�%�澑)��͢0ʪE`�"O��{��G�d�ݪe��pT��@�"Of<�rF�zW
�w��4C
,�"OhMr(�99Pqk�Ό
]J��Sf"O��P��]�f�N�:P&�X1��c�"O�,qR�L�4�������9��R�'44�j⊇�]�aS�h��%�dp��'������Y��e��:'@ [�'^ę�7���d[�$]�l��Z�'��0z�b̚r��܃1�O��p�k�'	���3)F��:���MZ�swX���'��-�EA4"��b�&�{1H|��'������� T�BRf�ά!?\�Q�'ֲ<�0MFf~8�`��!1���
�'PP����%�^R��
8L��q�'���b�&�*�-W)7��ݩ�'��eY�#�������x���H
�'J��v@�0p��|��8	�'#�x���.<}5�<i� ��'7&����5_y����o��H��'�nU�T��/�ɓB/82A�e��'h52ՠ�^���y2m�9 6&��'�`��ba_���x�R�+����'�\ݚ��ȗ(�m���8��!��'w�]�s�H�e2�T�$#����'�)q��E�T�K��ޣ����'��@	X�Q��d
���'�X"@��+ar�0p�z.�QI	�'�T�E��s(��ep�ɋ�'xx˖�ς%�:-PW�� �����'z|�윻6��H��6!����'���M�h�j�K%�ټ�Hs�'!���	�|�Ԅ�$��+�$u:
�'�a�&G|��-�4D5/����'t0�CT��$3�94��+6_�-��'��E(�K�pSnu�C�ݼ|!�1a�'��uh��y���s�4�&�*
�'v�0ů�(F%�eZ�c̯{L0�
�'� � ��T%c����!a��P�nX�	�'���"@�c����0�YVG*��'��{�郧D�J�^H��(�'�CgO(��s�-K/9�61��'��ڠ"C�}к���GA�=�H9��'�n��u�X+P.z8`iB�2�6Q*�'�QKk�(9�����D.���A�'�A�NI.=,�E�V@���l�
�'i ��V�L�7��-I�K�A���b�'njl
���N-Y��X8(����'@��qU�T:v���)�F����� v}����1,�%qWF�kFB������(6�����ɞ%\$��cn��wϼ)�eFZ�"a~2mI�(�"�����b��	T��Pɑ/�j�5Q@H�!wZ��P��Oju�O�Q��AEH��K+�N�M	h(�E�>ړz}X�u`R��~�i�G���듺�Hl�Ɋ�&�A0%2;�ar����ta!�B"a|BX�P�Va,�%!�˲�Mc�C�+�$���Otq�o�15=�bYwAh��'h
Y��ϻ<R��[�G8"��8X&A֐�ņ�'�}��S�v�2��eH#��Xa"@�5j�,k�)B?tT�qR��"�u�;N��i��4+E��s��aQ�1P���qW�x�r���.�Op� �f7.8Rca�:D�|��!,��q2�A1X���W=7�����x�&)���O�8���B7]XO` �&/4�Z]�JF�th,z�I;J7�I�WA[a��;1��t�7y8�h#��nȼhA��X���<R��ͷ!�ȝ�&,�E��Q��ώc8�lK��h�J��a���B$i�o����-S*5:��i��%�ݹV�P�+�.ם1p����"�*Ex��q�6}�l�)BE�cZ�
&G!@[u�WO�=9b'�;~������=[j,@�ܒ ~��#g��Ne��%�g?�)'~���#���7|���s���&��*
�L��)Ix9l�Ђ;�Op�����7�a0��!�JM+�iٍAr�=��)ξ�2��4iH,���N��M����6�UM�&f1�A����fڲP��RG�Ǉ%�j�t�:�k ����ԅ�~�dT,��M0��DI��K�;5l��!ƪ'N��@�'�p�C�Α~v�"�Ͼ�ax/�z�1T��7��-�ƭ��yBhLBwN|�'2�9�c>]�1@_7>��(����N�<�{7�Ԍ#�q��F��!�$���+a��E횵°RdmQ�(���߸�^�z��i����8�K�=ܒ�H�K�5!�d�1㬘2��3��bh݂L����v�愑�H���)�'Nq"H�ᢏ��%	 
�`�fc3D�{FE;z�}20��C��r��2}B�P&:;�|���Se�,�'ݩ-.H|��댞v�~0��o�����D�
���3?Ʉ�Yg���=���)L��}�^��,��/� �Kp!߿5��,��'�0�0��C�r���B�nC\U-S�� ��	I-,U��ՠP�4�0�)�2E�t���������������8]�G�. ̠���]E�]�@��Z��l%z���-��@E����(4����S��13�i�n8��S)��еj��9c�<��Ó�M�}�N) ьR�fDz���D��ɉ��P���H&�+b��)4h�=|�*TR��@30y����^�b�*��'¤F�,+��C���"O"}�$늕�2T�୛H��]��i�nA��W�o�}��>I�4u��	�)'���l�`h/��J��U�UK�^�L,� �,bC>A4g��U�^	��'ì��b�߄ 9
X���1C��q�lʈ,��up�C�_4\#d�4Zɢ��"K� :ll�a�8�9�m`���-_r���t
�r�J�1��'���(�������O`��[Հ�Y=u���عh?���!E�J 5��Ϧ�� �����ݩ �b�&�P������p��aյi��`��7�|�$�Rb���Ep<���5Ez��gK�-!<T1���ӋC%�Qh��ȞKRʱ�#K�3
�.�X���a|�iՒP�)����7K�L��uO���MS2�ڣ&W�l�F��O�{s�+&��-ZZw_�A��J���܌λo{���J�V��p��M�1*��ȓ{J���բ_5qUD\@�G��ɹ��_*\(�A億VԐAD�]�xO���5pQRM�P�]�
N�D�rl°�t;��Ŵ�6��D�Yf\x"� ��c�/Q�\�����K���!`�0���%���Z�<'M�3���ұ-ȺN8��Z��Lr�<�c۽�txr'i0Q��  6
Zǟ��!'v�a} Ƭ{��L�e��\��C�H��y�΀�|j´`�fs֜�૆;�y"㍌I� �#�#R�Pȇ	�>�y2B� G�N�W�1IH������yп|�(Y5fG�E�8����'�y�*:xb����8SvE����y��ݽ�uԌ�6������y���idD]�"�M�/�^��b�:�y��m�.�Z��R�/���	䄎��y�Ɖ�>r��WK��1Mp��v��,�yb*�?w�zU���N#�d�`Q�ʸ�y�1nnP�ɲ'?"� ���y����D9e-�r	^@`�*��y���(5e��/�C4�y��B��y�O������L���p���yBk��D�X�3��5N��%�w�Q�yr�3X��h��N�VTӴ���y
� �,��jT 8�N�ir��b@M��"O^ �p*W�9�4)^6x ���"O�q�㊟4(��z���-��|�"O�`��o�N��-��fG�w�8<��"OxB�Ա�а�Ę�3"P��T"O� P#��+7����)E�Af̹""O�ț�D�#(d�5HM%�y�e"O���jA�~���ilv�9�"O�8�T�]�sY�!`��L��e�"On�7h[�_=b�Q��
�P{Z�Z�"O����S�LB(�ҊE�*i^\{�"O�@a'��J�΅��*/w7��)`"O�)� k_�J���sh�i%�Y�T"O�L°�� s$ܔ��J�n��Re"O�鱠�Ð �0�#肤[J�
r"O����L��n�	��Y[���r"O�l��瞒l��H$+��-�2��!"OLZ�(���ZH�7��@ ��1"O���V���"1�0�T�5�aX�"O����hZ.\�8+���I,T��"O��{#�/�]Z�d���$���"O�fg7d��ջ��>[��)a"OV�Gjs��BT�޶8h��"O�q��HK90�B���`؃y�>�x"O�9�v#��"tD۫ �2e �"O��Jܺf��ش�@�}��9�"O��y�Ie�D8�F�J|�0p"OfqsD�����`���:W"O�˥&�3[�LQ�R$C��P["O���%錞l!@5[��>x�@�a"O���V��F��Q%�J���"O�JU痊l65`A�zZlI�"O�I{3*L9p���I3�"��-��"O�a
qI�x
�Y��AY@�Z��"O��z椛>��%yi��M�*�B"O̊SHE==kW�Z�w�0��$"O��Ӏ'w�tuXu���]r��"OH�9�酕#Mj���X�`�1"OtT��غ!Lp<��
M����"ONT�3'�L{���C[�5(�3"O>��"��
�\��r�Ʈd(&��F"Oȡ@��կs��+v)زN���zP"O������s�F�`���P��<�'"O�K��ΝL�p�R�OE����C"O��!L��9xh�'�)�-��"O���iF�7?���Tf�$G�p��"Or�*�]�0�b �����Nd"Oxhˆ儜j˞���ANtx�
a"O0dx�d
�x̊��T t|xdY�"O~����ɽ�(�K�\O̥��"O�젧��#0wLs1�I&�u��"O.�V!�1{�b+	
l�0H�"O\,HԦ>> u�*�, �|��"O~�cDQR�b���Ȕ�5�"웠"O��4���ȉBF7q�*Q�"O,�`���}���e��^ĺM٠"O���a�W���RV�M5?\n��"O�!�R	�W��ҕb�:@;��ya"O��"��T���Z� R���"Oj���E/d����L��P�"O��j!�Z�{5�� �����N�"O��BI۶FBL��2��#S����"Ob�@�l����:V�Ҽ7��Y2�"O�����@f�HxfQ�B��5�a"O� N��*�-bX���%t�¼a�"OL�b].6I��!������"O��9��V�`!�b`�މ�1D�d��́�$��� �إ6!��C�.D��U`����� �.�}SA(&D����OH
��ě�ɕ�~d�TB�$D���>��(���4´�Q� &D�<d�כm0@�3da�����#D����
ɵ�x���@ξ2��E�S�=D���SK/Ob�pd�C*EѪ�VK?D���Qʓ=}��8�Ƅ�rE�Qɖ�;D��!���\�0أ2����< �;D�L����~� ի,�![��ڒ#8D�h�f`՞W8�ܨ�MN0,~д�P�%D�l��f�&/�������9&����"D�d�I�) .!à�+lh;��2D��J���j~^U!���A�|�C�1D�Ps� <,@�f+O�!�<�Z�a*D�Y�D�-z��S���W�{�F)D�4���5@HU9�(�:Dh#�(D�|k�L�;�j]�Dh�:dʴ`�`'D�T[ãI�.��R�P:A��,a"&(D��w#O�9^�`�ÚP���7a#D�$������2��O�1̂)��/D�����g�|9�Q��x'��dG�iü� �֣��t҄}�lQl�O�09���V^��2C-ɻ`�J�1*ӓyOlO� ��O�*�Qā�t��ݹReݩn~ȍ:!�"�:S���e�?1�g�*�SB�N�3
�Mn�P�q!G�{#f�.1B����fH%p���O1��&B�B�L�aQ#NsyL�rVf�\�&���u�@9�甫gdtb�"~��Ǎ�At4'�@�8+�E�T�.}ޜ�dC�S>�	����)�C�� �#�C�q�b��+�c0�>Yi#�C���R��.pmHe@C�ĉ�plJaHS�OL��"��D�H�\T�"AD�7��A`�O����e�n1O>9�E�J�X�%C�5¼�fL~��q�D� EY0b�"~�!��#����'��ŭ�J��� 坑�����O6T��O����X��З��!lDA�V-������0�"� ���bS�ԻGh!�DZ�_�͓�%ԑMv*B,S�L]!��~a%��!Eb0!ߥi�Pza"O��S�$��n��W�ȦK�s7"O��� �9dp������-m&��u�'�qO�t�����Q�iT_�I��"O��W�ɹ�Б�%�D�	�ʭʤ"O�=����N�0��%��0ED�"A*O��2��JC�.�SFi�h� �'�z�A"Į: �˖���6�QB�'�6<9�oӓ%�$P�ՠɊ.ԼA�'u��X��V�S�F̸6'�-)�Z�j�'��Ɇ�3`*Aqfꂇ��$h�'A� ���US�XI�b��]����'��̛�剌c�`����Q<QF9p�'j�u걉@�W	��A��,Vhf�{�'ذ��/�zt��� ��zZ�r�'PD���L9,��R�a,���'U�Qr2N�/c�"y������8��'�f}�w�	>q�M���M-�r�y�'0>�j�H/i������)~&���'�8�PHB��r���LS]��'��`�Β�T�ҽ���Q!(���'�)��5���4.D2M�vk
�'�nybt�ԃ^���e��Uoʝ��'"� x�� &Y��|��V-LU%��'z��PE��XSP�z�=k�l��'���^���-�	A�s������ � 3�i�'����F�v=$�U"O>H���̤%�e��A�*@�BP"O��R"��=&@�j�F�N$�X2�"O�tqt-L�)5,Y��J*�]�e"O�dB�޹��}!�E�:m4���"Oj��g!�%^��tyTD�O;�t��"O��ŀ�96�� �H\	,.qa�"Oܴ �&��+�H�q�HYw&t	�"O�:�m�W�T��&ѹX̘�"O��K5䌙*��z����)F!�d��,�$p���$�M�����&�!�č�[�H�q&�����/j�!�$�8 �Z&�K+&ьQ��!Ԭa�!���d[�,E��`P�n����պ�'E��a[�[;H�u���x�
�'@i[�#_2o=��9���u�L%�
�'-��K���!_���D��`�>��'��L0�`ƵbP������^e6��'I<�I�&�2��ǅQ�n&1�
�'�,�JUF�+a���iS�y�(1��'��h�.n�$XvDW�c��X�
�'�*ك��@:VJN ڹ\����'�tX��?-�dq%��("�h
�'*���4�N�enZ%6Ȉ�z�X��'2������ƢF ���yk�'Ơ	�S�ܩK��-W����s�'��D�Q�Z�Dj��F*oԘ��'G����H�~�BT@�嘿mΌ��'�����m��|��@�ct�"�'���Q�4n�P�@E�`h��[
�'��q�AEٞE;~H �	�K�F��	�'�hի���5�6�A!�)�F��	�'Ϙ)���"YD�лā���9	�'��AȖ-��N`]��݂�tز	�'v�����"V�>��vE���2��	�'N
�S"��.p��ٶ��l�j	�'+�I�w@��r�H�ФI ����'c2@�q�ÓF�l��b��&�s�'���B;���Yw�Հx	�'�
x�&�݅REo��|an���'�
�xt ʼ	^4�:Ǥ���T���'�|�5��9N8��# ��� ��'��l��ZvrȀ�`@�.�J�'Ǯ5R��[BGVPIĊ�hz��	�'-FD���/:�6$#s*�lr���'�~59�C�%G�<���DV�j����'N�;�+ډ\��X��µbȂdz�'����@�5��43��D����'����C�P����re�I��t��'�4@����t�,���W"s��-Z�'�J�Z���aѰ��A��Z��ɰ�'��]���c���i0�6�2��'w�}�0��PT�6n�/��p�'L�	xpH�Up�9E��lg�m#�'�ft�j��I�\Y��jY�.70Hy�'$<�� X�&}���F�'.�2�I�'��d��A�,<����64�"� �'�� BʩFY*��f�}}�UZ�'u�B֥��x{@��+~)K�'u�l9�Lo�N�д�{�<���'�����D�"XpB�#��A�(�Q�'\�k��^Ȩ݁2��*I����'f��3�A��y�`�:󄊔m�r�+�'�|��4a�C}����'fJR����� ��	�b�����c�>\�PȲ"O�|��F��@���ˁ`Rr�h�"Of��^��\���[#J����"O�@�"��B,��s&�d��$"O��y2jɚH�ɡ�d�B��@yS"O>x�bI
XanzVmȖzӸ� "O��B�h^%	L��b,L��r���"O���)4�|���Y;�-�"O�ɰ�a��|p6BÀ/t�pB"O�i�G��]A�,�B��VHp�"OH\d� m,���1���
8��D"OΥ�Sɱ|��m�'.��Y;�0��"O �ag	JR�Ect��F F��c"O>i8��(?�pQ4o�(4,8�"O���55���B��%$@�T"O� ��w�|�An�Ȇ=��"O��@�k�SS�k!�Ļ#O°2r"OBݑsA�3��%��*��o*��u"Om��*ؑB`��(�d�(#@�e"OuG�Ά:�n�+A�ĺx�]�t"OX�+�IO"LZ,�b��a� 8�"O��2�Al�]��A��LJ���"O��e����E���1FP��"OQ
��ۜfy|g�0	��"O��!ס�%kK��R�M�����')�B�&ھ���ɇP&��
�'��]҅LƗWZ�����Z��@�	�'B\�`PiF=,��僙�S��es�'��{E��� q��q%m������'!Z�"�-��-q5���!�V�+�'_��1�+�=����%���#�tx�'M���2�J%n�R�+�j͊;��
�'�P��d�Z��na��V�\Cf�a	�'���2F@�'yEl��	�<8��'�tu��IH}(�8zS����rD��'z��g�ܗe�$1�2�ˊm�LD��'Z8�M�9
�]`7ወZ<��'شI#さ�)UXT�k˺{����'�LR�T�eⒸ�1oNp�&���'Wh�S�O8K�p�̘	>=$m��'���[���	#��yw�&A�I�'s��b�>&����6�!�X�	�'��u�P�f�f5b��!}��`Q�'�P�zT�9cR�H�!J;{A�@��'����+D;;� |���J9|W��'�nm���7u��E���{��Q�	�'5f,����+������q=���'I �;Ǆ�(�\ٳC�'cv`�'�<�H2@� #��`�&�6K��q�'���߰[x�y�'�Y�J�Z$�'��Ж �.�#�Ꞌ�|+	�'V�3E�R)~]�z�m:w|XPa�'�����߈���Y�.HkU^��'2�qʓ�G�! l�E֚c�����'���B B�2Gi��u�0fʈ�'�0�rv�˨9�4�C�"�Xc�'?<hBE�O�p�d��AL�"�Z
�'����M�s�p@�[q)62
�'t��	���Xh
ض��'�
 g'�8o� HB�-D�;r(��'+HEJ�B!A�,�1"�.�6��'�TA	�(��p�X���E&v`u��'��}���onRL�� �-%u�E�
�'2�p2�cÕ-�e��'sܹ1
��� �����m��*�	[۶T0�"O�q�e��JP���^�D{"OD�1gI�Y�`��O
�4��8��"Obр����-�Cɘy�5S�"O|Ly�aQ��c�G��m��uX�"O��!%��5,�K�-^Ɏ��"O�����Au��Zt�������"O������7G�|�����"OF��A'ɻ;z���ͩI�M�B"O��T�E��[��V���-he"O�)CA��n���H�G�r����"OLiQ�F�K���C�G�e�&A��"O�@��O�s(0���%>i���"O�`t�Lx�\���Q�h���PC"O� Iab@%bq��(��ɫC��}�"O±{eLG�*���Ht���� ��"Ol��!�
^��h!̈,I{��:�"O��(��Z�J��P˟:irP4�D"OАst��]z�� ��"n@D��"OLȃa�M;�քk�.�E!��"Or�j�(I-KOT��El��>25" "O�l�c&T�*DKu�0]nZ�"O���V�B6+|]
Ã
�݋�"O����E�v��Q� b w4<��"Opi��,�f�ɕ@ҧ19TI�"OHP�#"��� JC8�C�"O�l��X
,5��!o׭x!H�sw"O�d�A$�E��1.yX�+p"O�%�"��/���ny�|�G"O���$ ��a-�2 ,���"O�Iac[�8�&��E�s =��"O�����v��(�Q��+X<!�"O��qp�ҹx��@q��lS�0PS"O�y�"�}LŐ�B�=Om�f"O|!��k�������%O�l[�"O�T
f�Ϻa���xb�Z�N�i�"O���6�I*nL�Qqj���D�"O|m!��+i��	jD�����M�D"O��Rk�-%�>yˤ�L`z���!"O ����q��šHJ�ZzX,�"O��zU摋d�ZY�DQ�AoH!#"O>`��
�a.z,!�	X�V]�w"O.�����3����	�WUz �u"O`�+�O��m�H݈W�!9��"OL!r���#�.�I �J�"�:�"O�!�v�I�q�9���#W"O�a�&��>Mv9#`�.�0��U"O����C�N��0�ɐ)T�h-Y�"O�u"$�����2J&6�L"""O�)E$W�:*5@�eBlz�q5"O4���%S$�0�e�Ԓ����"O!�夌�>�x��[�����"O"4PЯ��	�|$��U J�,1��"OL(�x����i�+B�2��"OVm�	   ��   F  1  #  �-   8  �B  }N  IZ   f  0r  �~  ��  0�  �  '�  ٫  7�  "�  ��  ��  :�  ��  ��  +�  ��  ��  *�  n�  � � 5 x � �% , W2 �8 �> hE 'L �R �X (_ oe �k �r �z � J� �� '� i� �� N� �  `� u�	����Zv)A�'ld\�0�Jz+�D��N�2T���ƕ#Ĵ���8�?Yv�N��?�@`�X+�c�
ㆄhש�~@�a;�#��X���ru*L�5�>�3g$�
%�.!w�R��ݮ<�����yyԳe���!���CL_����q.�$KZ��I�~�Jy3�a�9a.���p��f�sK����X�`�!H���B��3���-�La�A
�:���I�|��0;^L��jݦ���oΟ �	���Iҟ �$�-b0�J)$n.���j�ٟ�	��M#�����OP���<y�@��`�HJ9yQV� �*�`@��?��?����?i������;1��`��!H�-?^Hb����J;<�^c��Ƥ��8?y�Ǥ�(O�5
��� D��p�͍2V\H���A�<��y��|2�Oj�@Y]����No>a��,�3�4��b�$wp� �O���O>�$�OHen�䟔��@�?��І�Y&аkK �^��f�'�6͘ئE��4�����M�e�"
6�Fm�=l��ň!�[ 5�py[��%�ޝ��؋a}�#=�К\��)c�R
P����O��� ln���;�By�OƖ)����n��nՐ�&�2�'{�Lo�?}���R^wW����8��=��(�?a$��`�i���[y���Z�0�^̻R�_35����Y1�M3�i�6-ôeN>P��-�t�d�V�	�MK��R%h�<�QI�Ѧ���4ћ��R�l6��$Ĉ�
 f�@F6$V͐�! �tX\� ��ֆ2�f�*�M�i��H��0�l7̓��@�4t v�������q6�)$��E�2c�� ��ve�ǉ�@��� 1������ H�fZ��I8���:����r&�����w7>��)��Ɵ���ʟC۴��	��5�.�q�Ľb���[rfph�\����ٟ$���`^��+�iT��\���<<����?$.�HCb��*UB��ώ�?�ᱰ$/� . lI���&!�x��
��9`S�9=��(�?6P!w��+I���"ʓ�,��'l:ʓ*݌��ɋ�]�T ��h@�z��Y�	�����y�	��T��vy��'�Ȑyt�Q� -�G%đp����5�'���Բ��|"��y�O�6���q6>�!�$&!&����4[�S����0�M�����O�.�a���6���h������e"�'�,���`qRwŞ�5-Έ���ȭR���j��XD�4L�
{(tL����8�p4�k_"�I�".-�R*$*��#	��=9p,��rᔛ~
�EQ���a,V$y[���'�W~�FX��?)��i�*"}:�Of�� ��$�D���ׅw^�QM>����?a���?����@<���R�ߛK�m #f� Asў��ɷ�M�g�i��s���ӾQtE�0�Kg�@�k��Ob��o���'R�m1�O�R�'�2T��sG�Iר0*c�&{0l�"���p�w��7 L�������Hq�O���Ɋ;<�tS�'�MHWG	�;s"`At�E-~q�"c)V�GR����THPЪ��#��O%�l�eDx?�ւN�Q�N�����55ŉ��,�M��^���q��O���/&��9t���c�T���Q4D�nNh���I����v8�����%�)�CE׸8����fl�O��dO���	޴���|��'���O)d�x���̕N��q1��5+q�$���l}��'4�T���OU�	YTL����ƥA�P1�& |C4��p؟$����iB@J��(�D`1���9V�h��U�,D�����N�@�T9¦N�V�']|��r�B�j�|`�@�l��l���A��?)þi¶"=�����B��(�ɔ2g��L ⁃`��Ij����]2#�X�p`�$����&%���	��'��7M�OXoZ�M�-���S�MF�=���<�ψ"jnT�0����P&�W֟l�'b�'8�	S bPL��4F2q��i͹H3�f� 3siU��=��'D48P ����@��Q��C�Fn��5�� �/p�]�r`΀=h�����C��R��4i�WxX��`�W-/����V�ɛ-/ ��RצQ"ߴ�?���_i�6��/Z�S���j��b�&m�IL��&�>5��/4&��ŲaE 6��P�7%5�IP�	�� �O�L7͘$L��t�V�в:X�I��:9Un���޴D��mY�D9j�,�*O���
Φ���1�Z\��&�=Y��X{W��^`���͟�3w.ĬNU����ː1�����z�x��t��R���RO=f$R��ed�;��I1K��4�� Э�̒0z���n�1n׌����?mT�̉}��I���޹r�2���.?�×ܟ,�ߴ{��O�1����7ڰW��Pr�`R6-L�D���|��'~�'���'[�ɰN`،z��۴C�pX�g�DJ�e����� lZ�����4�?�D�]�6�� �2Ɋ�x�X�Z�j%�V�'[��'��xi�.խ^aZ��'��<��2b8����4�'��@CF4Cl�%rƇr�d����?U��?	�I>��%��?�QX���e ��C�FJ>C2�� `P�/]>Y�#��nd�|Rt�5}R�M�a%L���Ɍ
g��<Z��CWL�ւ�I}���#�?Q����?���LҢ��% ߮D�X�)uLȟo�M�L>	�>"���V��3Z���hI�!��e�'��7���'����?=�'�
��`�O��Ԩ�],0��l˞*R6M�O��O��Şg0���oLi�r͊D΂)m��r�F�k����+��z��H��@��p�AZ�'��l����g��S'�2�Vty��E�6�]@@�!9w���bIjӠ�ǆ"8��z�"�$F"8����L��g{�,�d� }���pb�'���'S�O>"|Zu���4�>��'!s0X���M���<ٔKO�i�İ�r�̲Fw^�b#`�L�	����쟨�'�� s�cn�|��|uXp(�\:���)ּ֕�	Cy��'�B0���{�,�u����gI��Ol��� QQO��Z�}��̅2��t���%��tَ򄆌[�H5�%*��7� �S��Ԧ��0��/�61�r �	�t\14���9}�l��j�n~%�x����O�m������RU�S�k/_�lBG��*g��'��Ip���ND�Q��s��h��Yi���'ў��Ǧmx
U�.*���-�q��d�<�M�-O֑)Ǧ��	Iy[>��I	 &����%\�2���ŋ�@����ٟZ�n�3L5����ǅ;H��ؒ��9��O����i	�(��i�wa�,��1�O�}BEiϳ7A���`��:��~�@P��(��	�s�R�"�O>H9��'���S쟜��$*F�p��t�J��Ep�<ABNψ;d^t��êq���7�u�'��}�$fD� ��k��2SF��U�B��M#���򄖉/Ej���O$���OJ�4��$aȅ�����/�x@֤�-Op��+9.���A@���ӤT�F���P�NW�o��( .9��huo�����W���$���4��T�$�>1��P�#)�4��DoZ:��$�Im��O`�3�$O�U(@�to9ªp{���^c����OV��?���d��8w�i-JH�F#H
/���Am�<a��i�6��O�lJ��O��SOd��&�$jݬQHF�ĕm���j��J��M����?�����|��O���6%�`�.��F,ql�!b�>�x ]�S��Y���f����ֈ��IA����HS�U�t
�+�1[�҈W�%�Oe*p
Q�f���.T�zz �3��Ŀt]҄q�R�Fz�I?d	F�9�H�*��rD\�W�l��5�\���ɻ���X��^�>ʸr��0�$�q+�4��D�
�.4o�����������d�:Q����M�v���';��' ��'�Vs)�1@FՄM��xa�],�y��
�Y/���Џ��j�.�0l�g�z���DO\Nzp��	��j���Њ��^�,4Մ�(1R=�����1Cj*cM�<DzR���?�c�i��˓9{��$A�E4�I��N�;,�l�I㟸�I^�S�O\z��O�y�fI?v�L"��M��,��r�%Z�*|}ndC7�'�?Q)O~��4��Ħa��ʟ�Of�(Ҕ�'��J5�w5�)��ϏW�� b6�'�R�V	O��@In�T&H�JL�MS,���)�`���F��,S�i�-?Ix<�CĂ�mf.�xJ`y�A����Q���W��u�T�Ô��,˄79 ��D+�uJ�1�O|hs�'���O>@�&��m�ZI�f����D�=D� x�k�n	R$�AnFRj"�8D(&ړ�?a1�ɴ"���!b�*L���@�=����'���'�����/R�+{R�'Q�'!�i�,�\@Ղ�b�dd� �Q�)m��Rh�D�ብ� 	�����/��>}�u��'�E��яY�t1w@�P�;s�.��1��)J1��1�ሹ��OT*D�Fb?��b9[��MڀE��LՎ�C4b���h�4�?Ɇ���?Q��,O��ߔxL�B%k� Ƙ)����� �R�'Vڸ��Ɵ�Pᨰ�&FE7wJ�i���?�"�i�6-=��V�!,��I�<��_�G�F�������%��x����T,j}R�'a�U���O �)?X���BGi��X΍��ϙ"@�";"�+C����g��V��g��+6C��ĉ�Nؾ9��9��X�d�.l�d��EW��s��~5D��L1L>t���W�1;��1A,D7C� XJB��[�����'tJ6-MQ�'s�H�/&j�$�f�0P%|���<���7�ɽF�i�#��"�l��D�K�k� �O��o�M,O�Tے�����˟��W����pڕ!BOEjh��.�ٟl�	.B*$����I;�*d+b�y$�ȗ'K����F:w%<��
�;�����'d=��/E�-"��@�j؃0��6-�l�d�gkԉ{FFA��h'}ax+���?���i:*˓^S���"`��'�X���Y�(��	 P��x��Z�S���0K�A�h��qbA�	/��|��e�O��{���̔'*���I7R�,8�6�ܴ!�0I�P,�D*��Ī<�2E϶:J�&�'�Oi�����
TJ�$Ĭ���� (u����?�Rhǧo���'���)ܚ|�.,ia�-OXYe^���z�� �a�§ �s��[��8橌���'/%��j�ʃib�Q@�P�E]b~2@M,�?AV�i��#}��O����c��5s�!$f��$PJ>i��?!�����:h�u�ȁ7�������2���`�	��MS��iD1�$A��b��An2Ht#5M�y�br�N���<��W��2���?�����d��]����B0H {�	E�I�*ʓ�?)!���0=y�^I8�2Y6�R��w�ltH��L/���M'!H|���"�S�:��Dƌ�2�W�cz	�hΤ!�d�S�4Y�	�Ds>��t�g��(hv�Y�E?{��k&��"]X��G{B�O�аhG�F�_ːY���K�-q
�)/Oj�l��M�J>�'�.Od�:K�!����-�/����ZѤ�0�K�O2���O��������?)�O���:�f�(�Hx���9v�����Rk���J]V�i 1AR����&��J�'R�|�
� Xd�u�	pI�����[iI�qJ6{�@VEA�P���.ӆ�S<�x&���)ǜ=��!R0�πؐ��OG�2���������$t�X����K�p^�Ic폊g�ćȓ[�t��VJ��M�@Pt(� �6i'����4�?A,O��a�O�t�'�`�s���K�����K�R ���'7B �R�'��
�qm�h;0&�h񊰳��
Q�	��D(Q. ��H�A��@c)<�=��d(
8�+D�boDYAB���#J�a�M�U��UJ� T-�C򭖝�v !6�V�f�h�%��BL�O(�nZ���D�&1��h���v 0���y��'a|B�X[c���#��l�bC'��?y��'nN�{1O�'$̆����[�^$�������7gtDo���D��B����F�"��U�BУAl�k��	�g'�O���'Ԁ,+�n�j.�Q�hOEޜR�~�˟P�2d�
c𼙹C�ݪ aܲ���4*P`��c!��$�ַ`�l �"+�l�']�tFY�l.�eM.y�0�'�Z���?!��)�O�c���jh\��kI�kd���7D�\��.RX��E���E�ML$�0@7���čb�'�ʭ�A�
l�ve�WئM�-yd�|�,�d�<هn3����?����DC:~^V���N0��YS,C*6�ʓ�?ypB�*�0=a�j�~̄غc�ؗ$km����\���s�k1�?� ���]�|�<1 /��x��,q2�Z�0�aV�	��Ms�Y�Ģ�	�O���)&�X�7��o2&�� EH���8V�Aӟ���syR�'F��}���c�t���h3et��ؔ'��7��Ц�$��S�?і' P��@mD�Y��m��J�$��P�%�J�d��e�'<"�'2��O�b�'��i��'��Б��-i�$H�3)?B�68t��~>TXҤi��������s3�`���d�ZVI��c֭o�J�Ȁ)/���OX�,Tr��t�E;`�Z�*��V��A��e�V�nH1D�Φ#�l�B+	/rI�@�ܟܻ�S:9(0��3H��<��'Y���ȓ�I"Qƒ
R!f����^9m�"�%�PS�4��(1��R(O��Ĕ �P�"�� �As�!?��OXY�3��Oh���OR�;6'�/bj�OP`I�Nҙ)h�؂�X!h�0U�t%*Oh@1b�ʞ�J��կ�<0\�(�D0ș(��_=S$R5��u3H�J���܉be��'
7�O<�����3"R�h`%���A���<�����'%R�'�B<O�Ex��&0d�W̖9C�j����'T���(Qꩲ�%����pr�-��7�<��h�
�:h���?+���:��O`2g�t]HL�J/����O�����1���9������8Z�[�"NV9е��%lؘ���TF~��R�}�x��u�S2�0|B��7xh`
 GqV=���k~�?�$�i>7��O:ʧ��iLJ
��!^�:"�p��B�T-�U�(�	vy�O1��8.D�D���A��ۜ#:8X�&�O@��*�$�O���O��	���h A���H��Q�WAܝ�2���3�P�	ɟ��ɸS�`|ɓ�K՟L�I������?y����u��%R�e§4T�-�r���	˺�Pt�йY̤[RݖD4�|r�#�-+����z���"c��8ZNەb�����[����+e��0&����ħd�����]弳��Zn�pp�ɋ<0@�j�`F��3D��I_�g̓ĥi����m@��I,�Yc4L,D��i���+�9s�Q&O5}3M�<���i>9&��B�(5K`Ę�$D�'*�
��G�j�8��ϟ����������u�'#28��@
ݼQ�d�۴���d>���/Q��q*��^%}��@e�'��w锇5H�has*޳*��d̞�L���Y����0���X��p��'�&b��(�&� ��5jv�ٟ���41囖�DOy��n�f컗僡	�T�ę�����r�8��?Nd�9�� L�q'�`b�Ob�y��10��i���T5��,X�,u9�pȚ+2vd�d�<9���?��O��2M>���U(v�1�A���I$ :l<�LJÓZgȀy��C*(q��1@ޡ%^�Tp���L,�<yW��%.�a�'�:M��0D|��E��?���i�@�&��!�_�af�q�Y=VX�a'���ɽ r��؂�7Y`�7��0z�ʓ��=郰ij`�p,��F�,0ٓg�"���BfnӴʓ:�i�B�i`��'��ӣE����3���yU�%в����o�����'2��5r� �m�3#�Djg�=E�����X7M��\qq.K(�j���)�>M��a\�e�D��2)DĚ�k�Z����.V"%�#�
���y��VV~R'���?y���h����׾0��0;Wj�d�h%�V��-u�B�	Y���+M	�.�l[���$0��"<��Ox-Dz2$Ā��db�&1	�ۅ��R@6��O���O� �'�//��D�O���O���A/>!P���)�(�`oFm�Z�FCK�	��,Ϗ
�\�ئJ(擖=��8�E�O,�f��J~�8s3m�oWz�Y`ͺB~	��b���P�d�"�1��Y�Cʇ�~
� 4 q�	; lۄ�@�7>�)��cӲ�' ������ȟ�'r0+�cA0��훤�S~и�"O��S�I*$���6f[(\���%�'�2f ��|���O�	y�I��6�ma�Q"��c��3����Ot�$�O�M�O���'��)�P�Ħbv��!�'U)Z���� P�rP�P����vD?0:p�f�.�(O>dk���'�<���_M���'�פ>�h�y�J��P�4�$�ES��� ,���Fp"V�dڄZ��J!Oۀnf�k`�GL8� A�'J"7͐�b���<)�i��O�d��i�DqhasR�B�k,�5k�I�O �O��$ �3}�(��A^ �b�f��[�`��?�@�iZ�%jӔ�m�d�J7 �6m�O��D�s����;��2�)|f����OF�b3��OL�$q>���FY0��3df
2JF��b �>|�~h�L��h'��#�,��T$�x��k�)�Q���mV�_b|"����b����ǯ[����ʏ�R�z�8f��v��h�6˒�Q�T����Oʡl$���B?Q�L��jS}����7"U�8�'�a|����T]sQ�ÀUY��(��F��'ў�Ӑ�?���ߣ\�
8S��&�}�s����t�''���n���2˧�?qd�� ,�,X��E�lX� �X��?���ab���EC�H�����(4�Ȉ��I�=����d�)5����7��E�	�b
=�B�p���󷅛 CR\�zv,�7q-�\ȷ� ��~��6NU~���?)��h����#N��1�+L�ze�@�S�,#�B�$)�� v�Ԥ*t���`U�$e
�?��S'X��-��F�veh|����!~/>qn����'�41�1�O��'T^��sS�ԴO���S(�:;�\ce����B�MK�R�jIY�E.`��=�|:I>	q�0ob�|������#7��J��ͳW��ݹѯ@=�M�|�J>��ȼ@�D��!�[�P\��C���'�ҡ���?1����'�仳E^�R#N�_�ҍ�1,��y�@I< ���5@�_AҰ;�K����	�����'\�9�����&�;o7𕚒j�
'��h����M��?Y�����i�Z]0(���Nm
 �Y��>_9�P�ި�2���L�oixERD�K�'�
c���'vv�*�׌9�p�H��_(F|IaC? �Y	 �Y�Dbџ �%��jSd��$j8N��u,��5Ҷ�D˦���d!]�t T��q��Ѱ��n�b��g8���ˑVG�K�뙻ID�!%�谩O�Ӻ]�հK~J1����d���%7>�C�����'Q�'�bIʽ-���ͅm�0��ȥ;���S���;h	^1�!jC�@Iv�&��a�r�1�oB�>���φ,��A�f+�r�`^�3UHy�t)<��O��h$�'��6�Rby�G<sh\�̍6M��A������0>���ʊ!�2�;���&"Ʊ��F_��r�N�����s4"��Y�0���my���21���S��X>���8c�X��*�a�J%�W�1=�4M�	��0T�Y�KǮ�� ʛ_����W���Ow��ua)�����.-̼-y�O��%�+L5T�{�聡B��|� �?�S�lgV	§@A��}ەʊ5!�����1����M#���|R�K�\�V�i����J�]��a�<i4d���j�!"E8���wD^�' �}�*��o��IRkY�HB8)���՗���<i�$)����?	���DWy�I	��ޘ_g.��0b��wt}���Wd�)X�Ⴃ8Jv��D�<�x�ɹ./����]��,ph�Щ^n�#ƀ�K~��is�B� ��9k�;�SV�ə$�@����R<���"؇_O��mZ��D�7���O��3��^�����
/�&�/��1��C�	�J��신}�j�%EFR�P}�����ЛGHBCs�Z�t��%pf끈g]݀#���i�I�����dy��$H�Vtm��jV�c<��X�߉V&Ha:�fZ�MêU��(M�f9�K���z���	j�����6/f!��N�S�����Ѧ�����E���OB�;��˲%Ɇ�rlni��L�:|~.M����/ғ�O���5��+�Z=+WF��}��t0�"O���࣏@8xB�¾[��Y@�|�%�>	(O�ـC�Jj��Q�&`�
�$�f�9q�½'L�D�<����?1�	~�BQnǺ(���(�n�!�0�Y�z/�Q�'�fly��]��џ�	�K�_HB���A��M��E�^,4��h¡�A>j`� ��* "�tG�i�2�?�5�ip�aJl��F�����0nQ�,%���I�/�8����σ&n�
�.jJ0�����Q��M�
�S�I�GȪ��� �Op�(��AҶV����O��U�[^bE�w�˗`ɚ��O|�$�INHؘ�NT��` �7'B�����#^�|j'�d1
��e&Xu~��G����8�H!XI���W-�C���(�֗!hI��YF�h����Ȓ��O�Hmڐ�H���3� \Lӥ�ک&j {$�Ӓ_��A�"O|p��lG-B�tX��N��	�*�Ӣ�	�h��耕'˄P�x� FNJ|`��hq,�>�/O
�æ����d�O���<��0�V���@�aÐD	s+B�W�����Kv�������� ��d�|b��-T�d��"טb�d�T	�f�\�k6�?uE�i(���p<t��t�|�#�5����w��#o�9����)�6�<�%�IΟ���Y�L>Ysg �n�zǓ�k� Xk�����y�СP�����ݴk n�� �

���_X���I�<A�T@s dE!^�e|4t� 
�5Y��|y4�i���'v2Z�b>ͪ6�ƽ+g�Dz��ܘ${J�A����Q���@8ć�.S�6�p��dO��2�#��:rv:8��Θ�&~��r�,-�(5��[�^���#��{0�$�]�`���h��f�^ ��7]���ߦ}ʉ�d2���������L&��ȓPt,�+M#c6h(3�F�P@'��ȫO
˓;@4б�i����pn�����HyJ$:d+�#Z�=a�' �J��I��2�f�Ja���3�T�.��faxB[�O:\��F\��\`Bd*$�ۣ�'1z������'²�J�-�	\> 
c�C[1
�'gڡ3�[��z��$͋N��)�	��c�b!Q+*�����I��>���s4�ʸ��5`.h
4��I�d:�萳%֒[�Y�Ъ�x�	���,"�C؀r:(��
I'Q>��U	<�][�,�:�����2?�tlT�`�@� <O��Iɤ,ʧjޝSR�Z����ڲ��9=��'<B9���7i���8ҧ���H��G�h1 ��H�pe��j���y�ŀrG ��1�$=�Di���J��O4�F��Ė�@𻓁L�/r>��g*̯eI���'"�I�c�`%��(O�){�g�+}�XAą���@��$M�!�az���	��� i���r�R<ؘ'�Y�	ӓNVء�������J&�,i��sL>qD&�ş��|�<�7Ǜ)R�:��Z�8��U�<1� �6Kn��gE�m����Ui�yyb�/�S�O��
եO�29p� �05��8s7���Q���4L��ǌ�t�L	 ތ�5��D��Ń�Ǳ1E�� ��w�x9�ְA��	c��[�8�� P�'��}:��'^��'eع�G�S�S�<�S�BV�
^1�3!�s�H�u֨&���!$�8ݎ=���E��(O�HY��[�6�4 "s��#�D�9�B�_���X)v�Q�4 �$YŒ��$�P�<�h-+�!1���<�dqӶ($?�)��Q���d]�k0\U�P�<��
\HE� jȰ�&�ӗaT��*Y'��G{�OZ���8�p�ۋ :4������'�k2-�B���O"˧<�ک���?�`,� ���f�N�5nP<�?�j]v\a���j��Es�&]1%�Ԅ8�5�O�P��D�y5����<�e���<�P��&-���s��2Vxz4#C#��d����!�S�W��!��o1�fi;@�V�S���ɳ�t�d����.O�O��STydT��L�=!o>M.N�dY��"O��k�eFxY�T� ��4����D�O�XFz�O[�A0с�1��<b�g�}9`��Ļlr2�'�f��ԠS'/���'�"�')�ם۟<�F�WED|Y$*¶;v�X�bD�_(\FZ���s'A�#� �Oۚ����Y���.�T%��V�bܸ l�eh�Z!��j���}7ldiU	J+��	E�l��d�I�q��Œz2� 8�h�u��Uӂ�$?9@��㟬�	S�'^�D�9Y3I�����Z4hA�f�!�L��f�ª&��0�!�/��|:���򤐼� yA�ψ<�`P#�
%bt�0���z�.q3T��O��D�O�x�;�?q�����&ͫq�}C���r#n�ׯ�5$	�"H�f� �DH#K�8a�����dDy�KF�?	�xg�� [�,Ԟ����4yL�y�h�1�MI��D��H� !ɇW��c�\P�A�O�D��ىv{�|��Oe��#"b�OH�=����$w0 ��i �t���!��L�h~ax��	KF�}�@�V5cU��[���֬ʓ%*���'���9�
Q۴J������D���-�f��c�޺5�~�� ʪ�?9&��8�?9��?BM� W=� �Z�Ԕ(�u&�7�f؛��4�Pˡ(�N���&�Lr��Fy"���0x@г�.�1)$̈` ҆x8��dU.D�l�c����8�''Ҍ/"�]CT,O��&OJ���'ar�iT�|��D&ֲ<-�Y�l��6-�]��D������%Z& �N��Tg"�Ot8�'�*x�c��L�N�P@h�*n޶1�-OR��v� �Ab����O���y�O�"ᛲb�Tb�"^ ���bB��s�"G�>l@<����'�nԋt+֪<�c��7��T�?%(Ū]�>a8�qiӴSH6��Lw�T�PAL�/���:�����!����	a���oӮi&䡱��8H`HU|�P���&�mȤ9OZY��'�r����:�S�? bX% �r:f�i���P�p�"O`����26�������Ƅٓ퉡�ȟ�P	��Y���q�(�N��l���O8�u�$<"��i3��'��_���:G$dy��#,t		O�"s�"���8�`Q�@�N�'���?�n�'��X�Aăb��8���A���p�k]�\z�虵�O��`�.������*NL�@J����)"��I#�>�ďyy����?9�i5�3��d���c	�d��ȣ���4���#D��1'G�1$�E���A�vN��"5��O�)Fz�O��U�|�K�(��)7K[�h�P�Б�;5�	8W��џ��Iܟ�����u��'�1�t(�w��9e%4��@�b�i�3	ʍs�h��_�(���*7k��jd1�.L��(Ob�aҹ8�\$27+��(z�I�e=|qa@D7g�&t��,�;]�΀X���1t��e��N�	4b���ӰJ��!�2L��C3m��*oڬ�HO@#>��Z�pf�£�әWG���Ϟ`�<�T��q�/K VHɇ�^�4���'��7m�O~�Bʪl!��iQR�'���@�S7�p�%lW�p?��d�K�(�2��_�"�'���	�d����k�GE���|Ґ����&����I���)��q�'\��1��<��)�����>p�����J�f�&`�L�=݈Ox�g�'�r6�l�(��'��)-�,!d���Q�|�a�S�9�2�'>�Ty��	q�|�s柺��I�B�o����.��O�.�����ɟ�x
���%����T:D�]&�ؓO�T"E��Oʓ�?q���?9�'�RВ��¶�H�`�d�'l.N䨭O��I۟H�'�N�S�'�<=p�N��R)�C,�15���?f��C≬Ub\?z`EL�$Q��@�3�bH����M���m�H��'�tH���?q���?��'��Y�BY�@���� m��V��d�N�'
���'�8$�'��D@�|~���u׈5�1d*����
x��EjSP�r Q&�O�dV.\�>�Iºs���?1�'�?�')��*�˵\bM���l�f�x�m\,�?�E�������y�Ƌ5������%P?Ÿ5�N4&�8U$J�[L���O�hY#�'PB��?n��맞?Y���R��#v,�ЀKS59�2�fC
s�nę&�'�$Uk���?�G�'�?�'� ����M��O��nI�fل��㢗� �4 ��HA�Q֛�<OH�
S�'
��Z�$϶��e�i�Iğ����l�<-��mSS�hW C8N��a��	��<Y�OA����I�u�'U�\�@��x��
�MroV��&!��eEd)G�f(���u�`3� �OX�M�tH�����I�&�|�Ad��m!�H��D�lN��ٴ1����'�ܔӸi<�6���b�
r���?yj�oۂ�ڠ��ʂ4�l��EcJۦ9s��Y��M�0]� 	���MSc�O��韶9`�l�\�7ˋ�8`����Y�<��I̼��&]��e�U�Sզ)��؟�����`�'d��'���'Kj Yӈ�6wH���r	�0�b�0�$�O����O�O��>��$oH��>}Ĝ�F+12�a����<��?/���$�OH���z��"^��a��/��x�B6M�O�d9��$��?Y��<c�b�:d@�[�43�Ɩ}�'��xB�Y�x�`C �F(f8di����M;(O��O�>���x�~�ٕ�)��)( �E�\�«O����O
��F��O�O�dHA�ڽ�(����֬u!�d�;�0���i��l,:��ȜL:!���;"֑Ȗ�J�cz)c�f��m)!�� z�>�z���F:a�BF���!�D��*�А�шà\VH=K񥈤u�!�DI0���p ˚3T�p��K9,�����	Ɵ����t�	c�\A��3r�,�KB�֋r�n��ܴ�?���?Y���?	���?����?���~(��''ӁP�Dy@�<"Ѻ�8f�i�"�'�'b"�'��'
r�'E���߇.ݸ�c�)H�J�Ӗ(g����Od���O$���O����O����O��{��J���b1J�s��8�Φ��I�T�Ip�����	ʟ��I�#Tˉ]�=X%ə�?m�ȉSҢ�Mc��?����?a��?9��?q��?����di��#f��WN��A%,���'�'�B�'��'�B�')�(M�El C�¿<p2]1�Iː	S�7��O ��O��d�O����OH��OZ�� "n�9�׬G�ʠ��훙e`9mZ�����ӟ\�I������4��ן@�	%��p7���h�fL8�Dq(�4�?���?����?I���?����?��?�p�eg��a�ⴊ��?Z���6�i���'�R�'���'�b�'+R�'��|�c��&l���ą^)��Ԩ��f�n���O��D�OX�d�O8���Of���Oj]��%$P��7aj�He��i<r�'X�'N�'�R�'K��4#���Qn�-P)pIC�;&B ��i��Iɟ��'�?����5&K#��,;i�� Ʋ�Mcs��S���O/*6��@	L0t�a�T�n�ph��@XԦ��۴�y�Q�$?���n����/�v�hs��R*n���#�c�j�$1�����"��;9ў���<�p��K�hl�S�IT�j� @���H�'L�'f�7m�H1O�� ͓"�9��@��ʚ|7�A{��$c}d�T�mZ�<q,��#W ��Xo(���
�>�@��]����W1kݔ�9�>ͧ^ܮ�h���	�Lۺ��P��/��	T�J�Z4������O�}�F�J�֣��^,���r"�?����	1�Ms׫�p~�.{ӊ��S�_�<
���(ܑx'Խo	ZX���M�W�i1�kЬ)zO6���ѵU��ܴZEԐ)VM�
%,����<2C��D{b�'e�IL�'C|>�A�.еS�Up�"F��M�'��7���Wp1O��?�Ӥ�y��f� �@��1CA�����Ʀ�
ش�yr�<%�#"��"_,p�f�l�` B�> �5;�����~F�,�2��Eأ��'#��b2H�-|�Yc���<iJ>�s�ik�0��',@`:vC �vpD20�����hb���4���]즑��4�y�ň!M��]@�	)�hyP]�l�N�b�]�|��D˅Hܬ����n��i���.����j�"�X(�qC��H#ĤP�*ǟ���ry�R��~"E!\��$�[��|�p!br�|�I�M���I~��g��b�(q��b��,[��֫��[r'y���'u\7�����ɿOLMH�Op�crǞ�BȐ�z�)EOk�ı� ҿUI,*W��"�^\x��-�8?ͧ��w�؊��ڒP��Ap�BO)YQ�(�*�O��O�mZ [ �c�X��|�1I�7\c�ݢ���.m&�٘�)py*�>�'�i j6my��&>��ӽ
�p�	�=r ���؟w^ �p�ư��r0R����BT�:v��ºKM��خ7�<��@�Z1c���X�'M{���'��S��'?�g+���ñP��]ql��Z2\!a�^�<X*�OH�o�U��|Γ���d���s%l�e��=×���
7��OR�b��|}��'��q	�kLY��y�O�m	b���"��=r�ቚhQF(g��O
��?q���?A��?����Y$P��0"iտ&"�tata��u�7C��O6�d8�9O8n�<iF��Cu��x�Ⴙ��#�.��M��i&X���>�H~��H̥F�In",yB��ڛIy�1pl�7#��D�'4�H��`�+���OLʓ�?y�J�f����zw>��'�%}g`���?Y���?.O�n�:;��e�	�p�I�1+\�çK*tȴ�V�[-8LX��?UR���ܴ4���&�OH�'��]���3u,��7�, �0����tSG�@)l��!0py�O^d��G`ݭ�u�1��N�Bݔq!�m��z㞩�	���	ǟ���r�O���ؽ5�:ّ�*��@W�M�v4��-{�zAsB��D�ܴ��'����"y|iyT��]����F�Kxk��~Ӫpl�)�Mg�*K͉'���{D��Dm��!d�+#l�B�G��)��.nc�'��؟��Iڟt������ɚ+rX�+Q�֩K��1R3Bo�b��'��7�՚'<���O��d4�9O�A8bE�Zh�ȑO��A�8 �GQ}Bk�D(o��?!��i��\dR���O�5J
ѡ�- mz�`'g@���ʓn�$��ď�s�n!���<Q�N�,Rq8�߅G�bK�o_�?����?���?I�����R�����k�� N¸M
�����:g�䠻�
ޟ�s�4��'�6�U������P��&�����dr����K��B�4����PZ�9-�Թ:b�ל6�@&?})�;$S"% ���G�ٳ|=��ã�ԟ��I�4���@�I֟�G�$c(U-.�����~�l��B�X��$�O�nZ2� �ݛ��D�ĩp
Ӻt��,r�D�l�b���>��iY�6m���d�$��f��%YX��y2�}8(e�F65J�%���	AЂ�^�iy��'�r�'�2`�oǬ��n6�ک@���)���'����M�3���?q���?�ɟ���󣊺k788lސ/%���uX��H�Oʵn��M�A�'H�O��$�-a�tL��d���5s0"�,B>����o��@\���1{�L
\w�1O,t�E��!E�89B��Z���\���IMy���O�Im]�e؅���<�f�ck�?�b<�:?Iu�i��|��y�lwӲ���J?2�<y
v��~F�%�«^��y���>��}s�Oܹ{�+M?b��YZ�
�*���OC���t�o8�m+CJC`�Q��L-����O������P"�ŭxa���
`�V�1Ѯe���0W��������mZ���@�N)mF�3��է���+�۩�M4�i��d�>9���r�8��X t^�i�a��{5���V�9yR��Ї��런�W)�h���7��N����:O��C�^�{����
�K�,BA�'E�w�I�MCF��g�"�\,!'�0`�l�s�S�uꤺ����~J�I��M�ie��|b&�C )���Ѡ�͊-k����ޟ���Z�b�N��n����g�*
��no� ���@,UQ��%�~>���<	*O��-�g?������p�^�,��}�#���� �4AL��'��7�O�O�	�j𜂓�
k<r`#RѪV�:����Hٴ�?y�j �|q�	˟�FN�Q��m�S�iόt!W,�|��@&?�aL>�(O�$�O��$�O^��O�
W���%l䱅� �Wz�0)���<�ѳi�����'���'�dP>�	\�>p	0lX5���Æ�Q]�yk�O9lZ�M�2�'�O��d�O$rb��p ��!̍K����T���p���" \�<WKX�K�2%[w��'�剪b���dL$,;D�����P�	ӟ���֟���ԕ'o�7m���d.� v�r2��.�B�$2fv��'m7-%����dQ���J۴:���?AN|]��+�1�􁠰fLDK�TK�T� �I�5�Ĩ�v�!$.E�'=�$!��B�H�"�"3���]<'7���r�')��'���'wR�'D>A
C��)��	ѦC�k�U���OH���O�l��j����'�.6�.�I�+,�m��h�~�P���7B"f��v}�'iӤ�n��?��sj�>����O�4�C�vf�}����Z]�졀"Ճ9L���a[�]AʒOH��?y��?A�M؜��
�1\�B���&�v���?�/Oo� �Y�I����IN��c�!z���+�E�,���t����dC}Bev��um���?i��m��d�0��sF�"G)Y�&�!,W&|���a,O��ê��Ů�����dA�%@�Z1,�c&��(2Vx�Z���?��?����'��I���h$�\�G�k�
*_'�q�0�w��Ozxn�G������M����g���[VȚ�g��f5.��fMrӨ�k�HYY�:IB�(�K^�0[t0�O�Aru�]�8dH��pgA
h�<|������O��$�On�$�O�0B4*�)��0�Rc֨��܊�$��M�P���<!���?)H~ΓP��0Oj0	�é"�v�9*���sG�o��Qm�9�?٨Oȓ�R1YEf�qy�C�5SR )���<Os�5@����?�2%M
�,�T'R��䓊��Ox����,���*�쒹!|9h�g{�N���O��$�O�ʓm�����:�y2�'�r.E�v��� ���F] DH�9A��O$��'�6MFѦ�����k���a�*2�8(`�*�	_�r�)�㊴;��%?:���u�1OL8��kG�i�H1��F18e(���'���'(B�'��>}ΓEAʠ���O���ڹ~Ǿ��5�M�ec�W~��{Ӹ�4�7Om���6O���v��� Q0>_�(�I��M˼��v�iX��c��>Q�dטP���F�z�@f�]9�D�J�&�� �R-�䓧���O2���O����O�����}A���4�+�(��ʝ�kq�1d ���)����O�Lm:�S�U��K'�����8�Dʃ�: ��Otm���M�F�'��O���O�j�2S��kff��""�`�X]��$��'�.P�!V_�ܚF�F�uw�|R[����l]S/D�)6�8�����՟������ؖ������˟��	>�u���q{��Z�5H�{(��b,Kr2�p�
��#��t}�~��l�?!��^�m!�����F�� �{�mȸc�%ȮO4��у	0=I��Z7BE�˓�S�wm�$S��Ǳh�����fݲ@Ϊ�Z���?����?a���?1�������'M0<��m>-0�A�'�R�'�7O6~մʓ-M���dڴ@�=�a @&b��v�9��ľ>aV�ig�7��.�jT�@�I�&�%�:zJ��p'W��]+㣃>>X�@�@�hO���<�'C&�x�����U��n�/,r��8���66�vc����'Y������4�
���!�i � 	�	��M��iW�d!�i��
�-�{n��Ԥ��8���r��ՠ �\� �������?Y��B
��uG� Z#Z�����8��bW��5	�I���'����G�Mhu&@��"�i@┌[C:�``�O�V6
����4���5�#׭)��"�ԉJ�����J��M{�OF�rY���	�)��@@��[�I��Q[I3�(Ө*[|`Y��S�2�,!�I>Q����0�'3�L����`�0i�g@�`�ٴ>�d�<��'��&i�63�V��S�,pm\��WN�K��<H2Ne�
�o�<�OF�iꟾ��J�G� ��'E�8$`��YR��oőD�����'(fi�b_3�ZXH4�i>}�)�(��VA�8Ex�������Oy�|� r��<����7C�F�*F��'��e���
�*mJ� I�O��n��MK�'�� \�.��E�6T�Խ��-ȚP�P��O^iC@�G��h��O���s9j�H[w��"-nI�
�Y)2�+pOK�X�2�'~B�'����<Y�/S!�8[VeN2�������ݟ�b�4'�r�y(O��nZl�������v����ܜ{]@��P��?!F�iSx6�[æY�F�J����us�5�Dּ
�0����i~��`��F*ġ���kOV��'���'��'*R�'銬���ɼL:=
���3y!�Ȋ�Q�8@޴F���?!�����<�&%�2�$�J Sیy ¡����M3�i��� ���N���f�@��`Gè	` /ul:�:�-
5\R�ɀ ��@Q�ܰ��H�;�����0Kn�X�cҲ2bqF!�$k����ޟ(��֟L�Iʟ��'n7m�5DPV�D��+�LD�MFVn���5�J5�B�����Q�����U�ݴc��W^�x!� &A S#����L��U�t�I�����AV*,ļ8�'U�ī��0�i�*փz�|��'��+Gv����'�R�'=R�'���'�>m���̙v(gM�)�2E����O��$�O�lZ����MR�f��s�Ɖ�Xtpɨ�@��2�lx1�'��I��M�нi����;�듒?Q ��.?d���_�g�\Uq�*P���yB���P�M>I)On��O����O�ls�ǟ?��!���(�ܕ���O<�D�<��i���ɛ'E��'���P��qr��Њ`��A9��4TʓH~�I��MS�i�>��/�)矖�1'�M0I����E�H��I��S����j��u`˓���ʵB��.9���({C���E
*ͣB�����d�O��$�O��D)�ɷ<�s�ij� �}�e��%�(%9#l�%a�F\1��,\��	7�M���l�>q�iֈ�A�HJ�xĪ�(j�^A���a�tlo�v{lU;�O0���6h�`e�uOՠ�R�	��ċU�L�%A�}���K�U�0������O���O$��Or�=���� F��aS�a�p�V�[A��7�M��H�;�?���?iO~�w~��>O��DK��l�t�96��&_�J�1�Bu���oZ��?q�O�������N�v��'���as"�?y�����E�,Ⱦ��s�'��h%��,y\�2�|2V�����@�A�[ -K��a���pk�����	��X�	\y�m�`�������I��P]�'�d�<D(�j�Pu�?QX�\��4*�����O˧o�!9��ܶI
@`�+��7�bm�'�f$�2OҐ21�t�5��$ Z�7�֝�<9���x"�m#Dr�A�����͟H�I֟�F��>O�A�#k�6s���U���f5I��'�~7��T��	9�M3�"�O�=��? �yǁT1j�<X*��'?7��ͦ�8�4@���X���I�S���¯ӺE�zY��X�$��(@�!H�e���v�Qy��'Lr�'o��'�B�+��1� ��\�J1ㆉ ��I��M�W��<���?qH~�ecxH��%@�g����ZC���fS�<ڴ���
�Oh�8�I���a4��F�.�ߞ FTh��hY�o����<��a�4Kj[f��,�OvʓϦ�X$�R�Z��� �ұ�����?����?	���?�,OfXnZ�J��	%^ ۷ӊ���tD��g/��6�M{��l�>)'�i7-��!�ǘ@�8�� �8!���6��I����'<�1�ե$OG�Pі�L�rd��Oa�`f�����a�I�<.B!����2j,5���'�r�'�2�'"�'f>�Q0O	:e.$	2�[26V�]���O����O�5n++�B������@�B䦜	<T����J�f�D�>�3�ig*7�"�aq(�y}��'�`�s3BS7S:��a��R-d�ٳ���Ͱ��ƣ�64�'��I͟��	ş��Ie���R�Ca?�q��+C&4�I�h�'i6��2b���O(�+b��!{�>5# L� ,�Q)ck�cy�-�>��iO6����@%>e�S-쪸(�c�	$��T�G�L��@B�S6V��KR`y"�Op���&bݩ'���)׺h:`�ɑ+�d��ҟ���ٟ �	ԟ�%?-�'[�6m͝5�(s@��1N��k�ɿGպ�9��<Y��iM�O���'�&6��@Rp�-�y�"��;H�m�M��ߏ(���˟x$�4n��X��O�Hy"�Q�$��`#>�2�B�)��;2U�D�I�$�	ҟ ���T�Ot���+i�dl�!IALi6X��i���'0�'��y�g�*�I{���Q @�d�D�[���14rTl��M��'��I�?����?)ȵ$ ���ğ�I�@�C5�P�"+L�#C��NJ���S90L���6D�`4��O�ʓ�?���k�H����-V%�*����5N$ys��?9���?)O<oڏ~�	ȟ�I6[2i�"	��N1����M���?��\�h��4L��V��O��' �2�C�_3@�pd$�%LU����ϟ��5��9�*H�T��Ayr�O�`�jCAs���fFZ�꘽8'"�׸ _j\�	�@�Iӟ��N�Ow�$S�',��R��A���J��FmB�b��0ȧ���y�0�$/�$�0�+��ŷWM��������O�Xn�9�M3�i�Q�,�>��� 2�-%���`ÎonD�WB^�T<���/5�d�<A���?���?����?���W�KWr\����&��p�-���Ѧ�8��Nǟ ���d��@��'�ڐ0��T>�1�t��"u��Лc�>�W�i'�6��ݟ�$>��?��b3z����)�_�������	]�����
_uyr�V�UޠM	�~��&�p�'��Y���C~�pЃ��լI:2e�v�'���'�R�'8BY��Kߴ�jL���I��(P�###�ɲ���a�r=���'W�'"��KH�6�~�E��	g�(,��"��χqf����f��듪?�3�ɃM�8�ЌT���韚��4|]$@�1i�	u�L�$,B�=nl�d�O����Op�$�Ot��!§Q`�d���ֽ|�n(Pf��	B׺���ǟ��	�M{Sh��$���<�c��?����߷%oT�
$��%�?ѩO>�lZ��M��'8c|c�U���I�<N���fd�=ya�L�pI=n}�����Z����GlN�'9R_�|�AE�)ȃNn^d[$�
^h�,��B�	�M�#��q̓���U�<fb�/�-�,m�FD6���9���VȦYaݴ�yb���O&ZdV_]l��r���" \�RեEfvtMH&.��������ߺ��y�,�lnX��O�i�L������O����g~�cq��}X7J�N=��"Y��V� @��]���7�MS����|�����_����.	����,	h�6M�O�����z}��'3�`ke�Y,5�ܱ�O2�9#52� �
�ǐ7���(1���O��Ȉ�����@�EJ�]p�F��/=I�R�q�|����0�ӊ�M�'?��Įڽ#�ּ($�
}�)�iP�7Mj���'����O��1���H��!Z�ʔ�#��SU$��<H��p��8����?3�eH��4����N��ܸ�lW��@H7������<yK>a3�i����y���=~n*	*��>yR"Y�ddT�et�O���'�(7�����򉋚N��|3Q&�#?����J�r6R�'	����D~B�`�OF����!��T���yb�O��䀀���}��L��?���?Q��?q���e�� x���ƙ-*(��0��y�❢��'X7M%e"ʓKi���$����&b��J5e@�QK�OZ�o��M�@�iu���d��>	�7�|��T3F:� :��=�3+,v�<�1qJ ������Od�$�OL���O���v��zBeM�1%�	���לC�ʓ/Q��hȦ9���'D����'Z�!�į��(�T��aU�N�P�J"����E{�4L)2����O����Jtq�x���
gF����}��L�a��>h��	'O�H��L	�u��|RV��±�=`�Y�%�1ZkМPc�ߟ��	�8�Iٟ���ny�~�:��R��O|���φ8XlH�@����k���OP�nɟ�%���OFqn���Mk��'��#"�B>�`� ~��Zj�\B�KL}�'ݲx7(�=^BhĪcQ���Ӟ����X�pdQ�ē$b�L��Nԟ��Iş@�I�H��ܟlD���ݺ���R._2Yp���U"���OYmZ��!�'J`7��O��?����!u���%�Ё��Ո����d��1��4�� .������,�p�!7�\�S��;T;��Ia�E,0Cv�"�Ś8�&���'���'���'�~@�GK����(��3I�h���'��[����4y?.����?����Z�O�X`X� �6a��SPjG3y��-O���'2�7M����ϓ�ħ�be+��b[><2�[�P���3���%P�d�(P��	\�h���l��YC_w��'��������+	l�!�mG�zG��a�'}��'�2�'��O��ɴ�M˔)"j��S��<i`�!1/�(l��5�'4x6$�������Q�T�����r�BĄKyPs��M�Ʊi{6�"��>���R�eP�d��
�R��+O2�� ̓"���D��>{�Źs��O�ʓ�?���?I���?Y�����d��ƪL6~ό(�d�� �6��,2��d�O��d4�9O��oZ�<)��A�j(dC�#	�<<Ψ��aU4�M�!�i�V�d�>��'���'R���cU��AF�F >Il�+���)B����1��՟���`��C1��t�s��@y��'��>=�Q����	m�t`�! Lr�'.r�'_���M3S��<����?�i^<�x�a�/U��Lࡲ#��'B������v���	[���H"N/a�wcˉc?����M��?)�~76��i�.�x��+O��Ʌ�|�P��;�y�1��U W� 	�z�%,\��?)��?���?���)~��c2f�,�\�F�M�K�DqC��O"�o�� ����'�B7�2���?]��!�P)����NEP8A:u����#޴v��V�f�٠�fn}B�'sn`��Y- �x�J�	Ϣz���3%1}I ���'0M��'H�I����Iş8��ϟlΓ��������0��мIΊQ�� �<�T�i~�Z�'���'���yb��D���GA�{0t��g,TΖ�*S�gnӾ��Ir��?���;�-iGkY�"�4�F�F�:�ۮt�ŗ'%|򧤜P���b�IRy�H�DF���;6dȻ���9N�R�'���',��'W��M�S%��<�BI؛F@�y�͊ 'oL��q�O" mJH�����!MޘG�ʘ�M;���~f�a@�0F�d�J���	5�fH[sP����nm�d�վ�ԕ'����<�d��]j9�o@�U�D�c�'�r�'��'���'>%p0K�7&��p��4x��l�D��Ov���O�]nڇM��J��&�$G�N�Ƹ��M'�^����d�t�$�>�f�i��7-�
l[g��[}��'�r46H�*\���E@F	_�p5"&jI�=|i��Z]}�'?�	ߟ|�	����	q�.\p�d�[� ;�`� Tؕ��֟|�'�
6��8g���O���4� R�A�rQ��Ե��z�$W\y"H�>��i��6����'>���}L8�a��ƈ �$��
U�=e��Gh��E�r�*���hy��Oa¹�k`�!'�����[ ?̔����=h�D���	ԟ$��؟��I֟X$?ݖ'"�6-�?-�|��\� %(����6C��Ӏ��8�ٴ��'���^���a��&��@�-R�xz*LZ�F�;`�7-ߦI�jӸ����Ox��+E�u��L���<���~���GF�7���xrC���?�(O����O���Ox�Ĥ<��d�p��v�߆5�ā�s���bTh�4a��ϓ�?y�����<���i!�$��U�8�R`��.�h,�RB 1[`7�]զ�;���d���)�����H}��ˤ(�h�lŗI�@�FV�p �m��!0����0`�'1�Iş(�I%q\�� �y1b��	�t�����P��ҟ��'ǎ7�ļ4�	���KՎ��^Eɻ�bܧ5��A���x�#����M��i�����|Je�_5f
x��G�W�D�z���	��!�Q(͍��ٖ'0��λ1���<�F�K�邠�X�f�`< �����	ɟ���П0F�d<O�i;�)��;&|�O��f&����'��6�T�Y���j����D��X�d��$�d��r �!=,T����OpHmZ�M�f�iq���F��>��W�d́� �$_@r����Q�DH�q"t�I�>�: �'k���䓿�D�O����Ov���O��d,	�h� �Y7O
�|�e��5�ʓ}�����u��'�����'�jH�.Q�䁘g�̤,'0�)1�>1a�i�6�D柄'>��S�?1�e�P�<H �B@�xiYr`�vN4!��^ybf�3�qDt�M$� �'������`[�T�q �Cxy���'p�'A��']�S�ԡڴ�d���,B��rO_��0k�D~!�0��#�����y}��w�xmZ��?��[��m��*��l����řK	|)��On��DK�*���MJ,5�bʓ�j#�w�*� ��R8#'fL����B�����?q���?a���?I���� :M�vj��(���[��--8��y�Y���ɬ�MK�����DT���	B~-�]H�k#$��=��`q���I��U��R޴hÛ&�O��@�'�>a��V����׈čsv��[�I��X'Ȱ��C?�l=	�;����$�O��d�O��d�!MJ��׏�(	���� 2x:�$�O��5ǛV�� kb�'���?�(���[D�Ă(a�l�ӄ�<�@T����4jH����O��R�iM�m��t�E W1Q�,�[�L& �DԚ�-۟Z>;���<��'*��p��.�OF(+�	S�
��Q҂�pd�S&�O��D�O����Op��&�F���Y��
-9��:i���KE�0n�����O:%l�P��E\��0�M[�C�$(^&���Ř�B��=Q�"Mhv���kӘ�{R��b}�'u�L�
+u�z"U�$a���hV:�1cE�+�ΰ�R)�ߟ,�'`b�'3�'���'a�S�a�H�#fd�/6Ŗ�ZF�I`��m�qІ�Iӟl�	T�s���4�y��?";�2 .�4L"\yp.W�q�F@n�>��	H}����ǥ-���^��	ă܄S3Zt����[-�$�	�@|r�+����)̼%����Ɵ���؟y�f �?���/��B˒h�E��|���T��Oy�ng���������	7sq�蹂&�+�ke�0YS�e-8�W�d&���شwg��O�7�l>}2Wm	`J��h���ԑ�ą�O��Ā	<ݤ�gK�c\X���O�3-f��O�$sgR�5L$��"�O�V9�d����O����Ol���O@c>M�榱ϓ!j=�EN�E�Pp!�-�&3�E���M��(Q�<����?�K>ͧ�yR�Zl���]�4-�Q:Q���?�3�i�B�e�D���q}�'bL\lJv�'f؆=b���;6��U�Ĉ7W^�+�ˑ�Yy�'U�	ޟ,��ʟ(�	������l����n��;2����H�dl�'�6�\=N����O@���^��<��B��z=��ZQ�*#ј���J�-Vz�ɺ�M3T�i�Z�d/��쟰�	� 1�xd ���|��"pl�dz�٠jO�@�~˓ �ȳ ��>�:�d�<��A�pe�l�v��D�L+R�
��?����?A��?y���S�� �#@۟���j���wn*;\�����ٟ(�4��'ܪ�4���j��p�I�d Q�
)s���v��	��ࢋ�F}2�'�^���H�(m
>*�S� �����f�øB����jG �2��d����ǟ����,����E��L�\0p���,3�1��H�:�?����?is�i��q�O��m[̓j� cp�L�J�ŉ��b	����d���9b�4�b���1����������.;J�aHޓ>���ZqX�)�|3#�T/#� ݠ@��\����51Q��aM�M�+�?�e%ԔB�@��vp�0!�Zk�<!��*��!�Lė~�Θ����'`��L�r/�D�X@iǭNl}�-�O̓$�*�!� �l� ��-tż����L8uy�ҟr��%�Q�߶W�	 \�me�-H�OU���=�E �($�ո��ى^�<	���=N5��q/���`D�J4&P Gb^ *�2؁A��+#�x�	ϿO�A���'�@�&�����O��V-ƌZ�jh����,�H����)�j��O>��XB(�D�OR��<ͧ�M�#@I�!3�ذ��3-�Y�V�J�<	��П���ϟ���ݟԕ�y��i�]!ƀ�!���U �$}yny�6/V�
a��D�OF�sp��!r��)�O,����L��� �E�����Շ���aC�b�Șh�9OD�D8�D�OF�d�<�O�d�� УL^�X��G['��l����埸�	꟬�	EyR�܈��O�����=Q]nH��?6��1ؓ"O���_,�Ek�U�@t���0<)�Ԧ6l�*&@[�] p<�Ti��8��8��Ǖ�x�lx��͹<��i�ȍ,WJ4���ō}���+C�,���f�T�9t���`xA�qς2eEL@��Cå��j�HC���q��G�q
\�
�cɧ|��)P� qml{tH�(Or,k�χ>���Κ��A�-B�H�d̃IW'�| �`����?���䓍?���W�6��uF�d] �L�;�����φ�?Q���?����?A���?��dƶ��ӿi���EK8r����KGqL`00'S���	��p%���I��@`��͟����$���Q��2+�Fыr�ǟ$��џ����t����K���'h���:@!Z(F�ƺx��Փ���?�L>���?T�ɋ�?1��?�Ju잵��D�q��y���?A��?��?�r��O���O�.��E	^�։��MI�s�����|��'������I����	០�'!���I��&�|��GE�N�A["�
�2 ��!I2nL��t�ұ-���H0�B�?m�;}8�:�=��K�NV"�Y�#̏#Q�GJ��O����O���=�$�O��D+`��rd-��6�
|2��ݍ�T���O���O& ��3Of�D�O`��O^�D�+i����ցQ�Ŝ����D�<����?!���?!���?A�����ݕ���d�^pf���ơ�M���}�b�'���'?�'�� �*K���A�_�X0)��X=�5��k: �0Q�NϺ@UA�T$8e����P�'��lb�jF1;,°�3卮(�� 3�Qg����D�?4���v`L�1+����O<���]${+�D����0�x��G�5(����[2`�$�(�s��.�V���h�0M��� �H� e�Hr��(�nX�e-Ϛ�]�>Yθ"��"�6�%�͟jبJ�d��1̎��b��<_B�R$��' J�B�s�������	��t�N����	�|r4��I�"`kg�y��xx�I,S|$�C�N�2U$T��Ԭ	E%z&a� �(�<1��+UK�Mi��-H�d��#?V��̋D`Q�;�E�$̢XW�(J/�!|kʣ<���\�(�D��� �jHi�����©[�!�� ��130��k���b����\��x��)� D<A�d�J�D+�P�h4��O�Qot�I=6����4�?	���I��x�,u��B�r.�f�^;�*tH�՟x����GŜ�B�d��@�.Br�$�e��lU�Ic����5����c)3d�hg�M�]:��<�Wŗ�5��؀aR�p�LQdi�2oTf��	�n,<���a����q��g4�<A� ៈ��N414��b�L)r�� ���W�+!���z�%�R��wH��^1��)����	2�(�ku��+07�\�`e�Q���I;�����4�?�����ې&�$�O6m��Z�� 4b��9�l��'�Vpþ8-�Q��80!J.ڼ��=4�D�|�1Z��\@6�Z�4�sЉ.G7�)oZ<��Q����dF�բv.K)eў�ɓ�^/[q�k�HO�e��㏕]�s�ʓ���`���?i��|���i� S�I�:d�U�g�f�q"�'��y7��v*<,�B�%e�xь�d�o���T�i�d� �L�T�9��^`��%��k�O�d�$������O��OV�$��������`�Q&�ʠSŢH�� B�Q;���B�L9]E���MԀ���P
9cQ"�d��T��y�F��g�����nڹ��0s�i��y���R��Q3]��ZB^?Yڄ��3ܘ'J�A&�R-ݜm���M�8V��Oda��'������B������ND$�x��_�!�[ 	a 9���<��a�ȍ�jи�k��4��Ox1���Ä0�:��0�M�;X];A�؀s�<5��O����O��D�m�8��O(�SD��p�խ��1��4�5M/>D� �ŞeJ�t26G�j���$�z�*��(5V尷`�8Fif��%KS�K��[r��Keaz�I�%�?��J�w6��� Ȑ�mZ�xū�.]�|�8�i�O� D��9�;��O��,-����"��ȓ8��ɇDC��M0Uc�86���[q�	Vy�O�2��7��O,���~2Wʞ81�$���M*<�q��s!���'�r�'Jr�Q�G�	�`N�	�T?=:���8s��(�c�^/���Ѳ�=�n�ƍR����jV$㉛Uⓘr	t�F�z����dH*n��#=��NL����򩕀3��p�O��HFQ��\78!��K�HZ���5DY"=s���-9�|#*}R"@��r�k%�
P1���լ��~R��/=FV6��Ol�d�|��N_��?���M�1&�#����b"@!"ø<��'�s�ܛA��2?tҰ�
�3-�Y0R��=�Z�q��Zx*�@�P�P�bGE�,���ȳ�ib�8!��"=+><��C�'F!�La� �}��N^ ��u���^� �sce5p���nZ�V���⦩-O���s�^8�GV�Mli[����p��T�O���<�O�j�U=Gs�Ī�H�tǆL)����OXiDz2�O����=E��Q�7A��{s�#��>.xZ��O��	@��O�\�$�O
���OШ�;�?!�4q��U��{Ԝ �q�M1$i�$�T��T�"�3��B"g}��$Z!zBa%�0�4A�.���C�,���Ѧ.}�և�{��xS�V�@W��O�RdBE'M@�	�Y��9����� ��(7_�
q��w��X	��d��f^a�,O����>�vG��!z0;���9v�쩃�L�Q(<��4.���bgφ�@�BAKW��c<9�§ ғ�����d�:틵�]%0�٩b�S�f(������!/���O��$�OB<����O���v>Ͳ4�ȃ;M�A�T7@B�-zQ%�/V��adaV����rg�Թ �i��QvxQ��D�Z81���T,���(aA�B��q�� K�U������ͦ���hd�^�<y&�E�<6�
S%�r�iLp�-��fǊx�!�ߡ���� � 7P��r�����x��	9W�� ��%�m�5Cl>^�ɗ��'��Q���T���O��&{����!�! z��+��N�6�jrMD�r�'x�@����q��86��~A��4(B�\�WK2N��h�c�'��A�m� �U�����
��B���1h��p����HOR�Q��'�b��T�i���:&#��c`$Yf"\�4r�!	Ci�O�"~�ɇF�̸+bɉ2~}H%�ʯJ�����J{�+6Xq@��
��%�b������n���'�Y>� �.���	�m����JG'߱g�X,P�ՆPsvi���ӥC��5�˛�m�V�V�6o>eC��\c�r��Aĺ7b����AG�\b<��4v�494@�!,y�<!�����u����:L�`��\c�<������ASH>8P�	ݴ9��$�	.�M��_�������>���9��y�3��4��YzvC�f�<i�HqHVe{'�Z���[_��?y�	��MC�4n���a�Dzm4��SkI"n�Q���''b�ހ9|L���'�b�'��Jiݑ�	馽��k۵4!ƉR��P�>�k���b��0@�+]�eP�n�&�j�'3��9[��.�d��2��8�r���hܴb�!OVt���=&���L�Rp���Q?y@#�[47�'[�X��eA1��ا �/*�!9�O�֐��,�
�]l�hy&�"'#�A
�g������M;�$һeY����	8��A�\�#��"=�'��ZL�=� n�iB׈o��j�I����]s�n�ݟ�����(��"(�n��	ݟl�'0�x�����T��@�	Q`�B%���׀o�v�J�OFC�P9A�X��O�K���$	2�}��o�YP���<%uZ��g8��:���7��?Q5�ܟ�H��N,-�D���	�-�:=bD���d����4��'��"}��E;��Po�"�f�(���2=�B�	�i�Tm��I�J�(��6��,2���	���<y�-�0���'��T?3��=¡�45W�ј���0-UXhx��?Q���¼�Q������_�?�(,��́ny���t�)؟[3p�j4f,�5ArN�M��1��COUAʕ�Q�é! ����M�)�HOBI���'�ȣ|�K��YP�q�IS�a���3d��|�<�ƨ�X=@A�wA�0�s�r8��CH����������5>*�ζ�Hҕ�ɺ�M��?Y,�����O~�DxӠ37/C
k7�&ˊ�;N��W�5R�� )5d�[�D\n�;�~� 5��.���3��\cTd�7Iȵ}V^-�C��}���ݴ�� ��ο��r@	ߒ8��(����k�p�>ט�v��%�a�L�S�������<!?�7Ҵd�r�t�L���:��i��ze��	d�P-McmC�';��'v�O��f`v�"A�)Ḡ�ˌ{��'�&"=Q���M��ǂ�r�2h�%ϝe���n	�y	B�'���ÄdO><�B�'���'������lچ��8�։©LZ�`Sr���MÞU�*�J '��u_�	���~ҶgY�n�O�_!yO��ʓ&��@�kS(/+̓愘*i���2�H� ��S-���1p�|�E(t�6�B��7wFe�!�J����l�`#\O>�c� O7_
�)y��E	b"u�V
O�7-N�z�sň�Rq�!À��i"���4��O���NH�~Z6��vʷG��D"�0�=��e�O����O��66Z4���O���j��򠇎�~���J�k�F�P���aSd~����3��a��:X[ ̑�T�iV�̠��u#�ŉ7y��`�d�D�\����'��9��F��]*��Y�o0a㕁H7 �����% ���4E~�
\�H.�2H��r����y�.$9�9+V�աq�	��%	��~�#�>�-O����g̦�������O)�s�' �+N80�w�.��B�,y���O ��.E���aŤ8N��90NH�B��`z��ö-B�Q��&.~ށ�Df�jF����I8@FQ�D ��0�'`	�^h�3$u�R�q��?Y4(������Ȳ�8ʓ8$���I��(�L�ص��XSDl�_�1�*"O6�bƎЖb�|Ez���J�r��'�>���4���O��R"�"�r��ѷ$�ء��O�t �j���U��ҟ��O9	aD�'|Ҽi�8� 'lS'Z8U����S� <c։��b��J�Ѷi��GBT�B�'��Q�x�����x��P6Y�����!�(�J����iȠ��%��(��,�QcQc�L	!J��M��\cjxɐ��>N���XW���b��Ipݴ�z(����S��Mp��`��ׯeu@E!��B�<9�,�4%N"�H�j�����9}��?�s�i>)o�s	B�b!D< �i��:l�x����?�"���w:l�����?a���?�����w���(����I($�#��	v��ڬO���'��R�j��'������� dX����B9P���O������Vd�����'�~�q��صS�2weЂ�0}�O�����'����A@y���Έ���da�a�<��$`�����H �S�V芀ژn%*��.��HO>�a��*\�@���N�=t� `��o�0Rq4A�t�؟���H�	w�@��I�Χq�!��ڦ���'+Vތq��S�83�����3�O�h��_��j6��f�`�COD����#�0�O8M���'�7m �X�dCW���z�(�� ��y��P�."�+w�Ե��BH8�y���	}t��'М|�`�sbCù�~"J'��@� ���4�?�������8z�@!01�� ���-_���+ "�ɟ(�	���ʧn�O��R��+���:%�m�b��"5B]����Q�u����g�<A���;5k���$�g�B=�D�%	���FE9Qj2��&�S��˅h�DM��<q��H��<���(X��*@��i�J�;3͏�-�!�$��N��6�E��-�&�����hO��J���5��ᣓC� T�v���H}��!�:dl�ܟ���S��Ws��'d���Y� w��3v)>��
fiX,�S�\�E��p��D_ D0�AK<8�AY��.�s����)K�l�Z`�rm��ktӴ�H�^�o+h423��)q�-���`��\c���ujZ��c'_ʎ09۴}�N]��+��S��M@ X�t/���/��Q�n0�jFT�<Y�ɇ����j��F-zi����VRܓ�?q��i>}n5Jcx耦	$4R;fD�	E,P��?y���23�����?����?�v��2���� ��!�S�5�P��L��d�q��υ*��H� �J���1C�Q�0`��|"�Ĩi�` ��qe�E*���(J�0�ա66���p`X�0v_?�І�*F�'�L��%NE�w	F�I��\-�D���O�Kp�'� ��Ă�v'�3E��!{J@��]�n(<aݴ1&-!�Q-(y�0�4�ք
JZȊ�-��|�H>�����0)@���L��$�Й�,�CU�!!��?9���?����?Q�������/!�1qشMJΝ��o�A#��T�!��M1�O���We9^9���T@�sM�h���A6��A���}P�0��f�>�:���5�TsP��	�6L���6��4UԔu�-�ud˓"O�����V�y�����,��g�U��"O��I5�S�%Լx1ׂ�F�p�O��n�K�	*T����4�?A������U}�a�����ȁ�T�2��)�v�������ğ$�
��op
���^ЦyRg�� \�a��J]&�p1,�����7"� `Gyr��x]�}q�Ұo�r1ۤ��	$n����E�?w��#���g�-8�E��e2���'E��'�e��o�Q>�CÈ��LT��L��=` �c�1D�\Q4�� ��P�o��Ni��Qi1}��i>��L� R�/ .\<R�:�Dۖ��嬰�� Z6�M��?-���@�A�Oj���Pa�00Rnu�Č	x�ڑ�c֯+z�cZ�V'H��T[\fA+F�k�t�Ɛy���.�Z�)���-/���Ժix q��e2+���E�H琡���w��5F�� H������.8�q�`��'�M#@i�ٟ��M>E��4~ʢ���F@ k�j��$�ܩ�ȓQ�
l3Є�7X]��U%�L@Gy�&;��|�޴u\M���D���l���PY��'��F�GjL����'V��'~bMj����K]���J��^�%,J�HRa�5'm|�y�
�&D��Q" @	�$S,�����3����90i����'r	�0 KD�Q���5�~}J�AƠݪ� SGK��-�6[�%�X��(KJ�DT�޳',dp�eA�>i�%៰i	דStq����2ٖ�3g�C�\�*)�ȓ$�p��%�5>>`�j�O4�IR�8��|�K>�֏�Z9\�&� 10�p�rT�8X7t�j�L��?���?��(������?1�Op�����Q�qwW�ۢ����b���y7�Lע���4o4��k��(O�]��hإ$��M��%@�rLYa3�A6�𬲂�Ʊ-)@ $�iꬹՄPb80m��}b�?A4 �=h���t
×K
�$	R�A�&jFC�	�3"XqG'  �@��O��
�"O��q���v�z���62��M ��O�MlPܓ�'�Ӹֺ�z&�Ǩu��i�Y29J���-�d�[��{U���|����7~�Q�p�A�_<P���0ǘ�[�^D���Oj)r� ��.f�!3�߸X߰)�g"O��!���8��)���.j���"O�(�G�ӎs��X����u6Z-�3"O^H r�=7ɢ�ɑf�-8-���"O|�0��33�|ˑ��8?\(�a"O΀�0ć�
�(䱷m��$�"O8�(�'uj5㕫W6S_��Yt"O&��@
6l`����&6Ԍ`�"O ��/�l�b1��!���"OZx�bj[�9u �2G!!:�bE"O�yj3C��R"��C���'0�@"O ���� ?d�<��Hu��pZ�"O�y���J�z�v���)��7�>��$"Ol���Hdr�tH��AX:��5"O�H� �(o�F�bG�1�2@�6"Oh��Q���[Px�R&�����bu"O���7cݺ
��C�
6 ��L�r"O�ت�ψ�yN����V��]��"O�b�	ȊL�u._22͈h23�!D��h�'9A���dٮi�^�2D�H�悔�UO ��C'!fx|P��5D�`*JG0(tpD2`8x���?D�LI1˻'��g$Q&T  tS�O(D����A�*-y޹1� �+nF6�[�%D�h�TΒ�9ZF�J�7|��)=D����H��ơ�P�\�A�&�(�a?D� �bIŀ<�H-Jw,0|q@$"&D��(R���S����w��J�����'D�� P�VN�}�)�����y#�"O����FP�t���#gc-Z���d"O�`�R��QyT0�P:��e��"OL��-Y�!p�z�6�����"On):�b�Iᄥ�v�R�o��U� "O�R������1�˚0���d"O�H�LD&7�T*�
�"rl1��"O���*TI1�B�H5�7"OJ��g(K�iq�9h�Ie��%�"O$�w���:٘�e2��Y�"O��� ̓Wbd�х�,S;��;�"O������\��xVB_�?EĜ�"O�9�C# $N٩��.wGBU!�"O%�����X�L�����o�d(�"O���"2Oͬ�Zg�ӸXi��S"O<Y{��%M�*�ț5%����"O���E� ;�n��p卿f�]�V"O�œ,K�i�ʬ"äC�IʮI"�"O��0T��<;�k1�ɏg� 1s"O�%-,�`;� ژ^��Ģ7
]%�!�dZ�'+2�J�O�.���wK�+)�!��T<jP�X����*9���-�!�H"K b��uj�2��Z��VE�!�dެKhy1I8&�:h���!��ޭj���2���I�ܴr�ėa!�đ0-L�YJ`�
�L�TJMj!�dGf�����+{P|p�j¿fT!�d�XH;�l��bo*Ґ��.CW!��t�� �۱m9�r�\3&T!��W��꠆(OK�՛��G"A!��K�rERĹÎ>ؐ�4ɁNI!�UY����C�R�X��$j�4-!�X���K֮�+�L��
�!!�6�$J4�H�O�)"��z�!�dל8K.��M�x��)p�	)�!򤏡^6b��q�B?;澤����o�!�X4`ق�#�D�IՎ�g	�B*!��8 =8FB
x�`<�"�uL!�䗁���D�T�#��i�BF��	=!�D\?��;��pb�f��Z�!�D�?����Ƒ�w`���H��!��:3��ѫTCإ/���L�)3�!�d�ڸ͐��2�d�Z	��.�!��d �)��iX9i[���7J�!�ݹz�@�h��2Zd` bG��*�!�d�d��1׏	9=�vYV甇K�!�A!� ��k��J}D��@�Nu�!���j'Nq�G̅�fg��Q����9s!�i�"�ؒ/�>[�M��ٿ�!��Ŵ�.����n7}��hD+z�!�DX�m�B1ꕊwC^�XS揓s�C�I�W$\dJ�	��-�X;��
�|W B��c���AË��=�@��1�B�R���+C��QI�r"��C䉇8ʀ��fɈ�z��<���\��C��o���	�#Z"�A0��۶C��C�It��I�l^�L���.XX'pC�	{�����9tƎm��Ri�JC�I';,XkI��V�L���a��]jC�Iwe,�Q�CϜ�B@E�:|C�ɤO���gmL>x<r=���T>t:zB�	=$-f<�"Cl�tq����&Gu,B�I��z��&FAa��P �B�G��hڤG�{�.�1���,BjB�)� "�R��(,����_2`$HA�"O6�#��� r���S툴jj@21"O�`Ve��l5~���7n ��"O"��q�Ky�U���^t���"O�Ib!���r��U�vހ���@f�<9�"W  ��-�~�p�/�{�<AFa^1[�b��6�U��ȴ��΂h�<�+��p>�`�R����Q�'�h�<�B�S�Z�ڱڢØ�}A4rf)�Q�<i�.H�EvP�ÇkX����v(�Fh<!��Ğ��(�q��U���qv��q8LB�I�%��X9-٘%�<	����0>���d�2N��X�f&\%L\���ǗS��ؠ�(9D��� ��q'&�
b_+
�:P�s�>1!	�8�Hq��x��iI<^H�l�2(4L��abߕV�!�d˟eF�t�@M�)��H�b��-��ɪTY�"�0\>����*�~�y �:�@�f�1��}rHS1	���蛟R �X��<`RR)�&���Z��EOڕ���#&�\�0E+JVT��6�I��B��`g�d����4d	8d�١�]>�Ρ�g��%�y��/�p0%�	�����G��M�����tA��<2���)��)9SC>9k���e�	��1��)D�Ԫ4�O�w�>a��P-y���j��-�?q���['��/|���R�$�?�=!w�շ��Y
���-r�J',c8�̩��2P��m9U�YG���s� �9�z	�Ί~{�U� ��L؟��1N?^�XD3b�ֳT���	��>ʓ!.䅪�.D�X�Nls@��ħ9�!��ݷt���� ŜU}xT�ʓ&�P��A*_�9sH	�A��]�uzR�U	��������]��S��?�BN�c�n�� ��ZQ+��B`�<$HN�Af��S�
��
��l�7d�#@�B�J�f�4t�@��zKX,�g�'�ޡ�dnC�A�h��OK�O�
y�-�4�k����q� iB�h+|\r �S�
� 	��$�<�Z	�TL4[e�6B"
�ƺ{9� Ey��
�V\��W2E(����Y�,|�X�F�6
w�xyGd�	�yb/�C�K�Z}��k��H4l��`nZ�B�d2��ηrJ���-�ȟ��O�x�bZ�G�m���a���y��6�U���,J=���b�Hø�i�-~�Zԃ	�10Y� 9��XV�����.)Diav������á�/\�}��]-YV�Ң�<E�:8���ʟ�n�a�Y"In�kD�X���D���0�РJ�57�j�Cf !?ў� �$íO' ����lAW�Y��i�95JZ�!Q,��,�R��D�/:;!��\/'u���6�u����5e %B��i��0whY<[[(z�<�:M��@��-Q�T���ӫ[��{�'Z>ɠ#�K�h�-ů�5"%�|�'�8����V�Y�S��hS�"H����	U���!,]w$�ku蕵S-����U5Q+�eY�e�z�^������+dQ�NҠI�����
;-�4�	�Q��q�� /oʽ��a" _�AF{") d�ViZ� ��t��h(Ÿ>�<"�!;$l�F��Ӧ��>:PC䉯qߌy&��X��T��e[#>���X�b���Ӆ��R���^/񨟌��V'�T2,�b�+X�O�d�Vh=D���wl�/)r���S��M�0TXV�	y¾��"g
:Ӵ����B�c���g�'_~E��'\��hh'�~��VBpx�H����+�6ERH�!h�M	6�K�=,�F��2$��)�F�a�a}bg�4E���B+j�2q���7�hOv�AS�|�`��Pj�=N�|�O� �x�O>{�|��N�~lB-�K>��4�p=�ŧ��VOn�����<
�u����<a�d�j$��Ӏ�6y>����ix���-^Bx� ���02t)��fٴ�yb
!x�����KB�k��P�Fi�'��ؠq$P?	���)����O>!�w�t(#���Jl4�zR�;(M��J ���,� 5j����P�e(@xQƇJ2[�x�&��
7-EH�	��"|�Fꍭ�$�J�V��y*���O�R�d�<�RP9N|rR�S�5���n]�Lv ���OhyB�'0��  LO��xd�W��Dc�ށv�(�b&����ֆ����c���&7͑���̉VJ��br��LҼKuF]��S�? 8m�VaN(J�Q�q�D�Ř@q��	E�Of�E���]��d0 g)��`� ��':�* �hT����o�)f&m��'��!� ��9nkF�C5� �+�&�A�'�45s�'4�@�bc�!�HDy�'J�5IuN�Ot�p�4G�")�YS�'��hPlN�%l���ɳ,۸�C�'�TS��%�V�)qǛALAp�'�lr����Hh���@�R4.���'�����"4��Ŏ7!K�\�'�b'�+c +T�R.5��d��'q���&�'Dl�$B�!ɼ%�h��'�8p�2��Y3��T�ܟ��J�'�	Z�`S����V���	��'�r��l_���ݓtj@��6���'2f��Qi���zW�gu���'d��x�!U-O��A�P�����'���ҒN�'��KOΆ:��l0�'�Љ��"�!#at�@o��qH�'A��F�����pА0����'$���Z'e��G�X�	N�I�'�(���KB����v�
	�4u�
�'�p|�ֈV�+����U��9j
�')l@Qc��(��1��BK�{`���'���"N�B�HeiJ������'��q���θ@B� ��(�U�p�3�'��x��M�0l�m�$b�6m�Qx�'�PXv"�;bAp�t�	^���
�'�n��t�@f���H�T��y2�'��RR~�`L1$�D�N��D�' h �9=>Պdɑ�I�H�I�'j�ԫ�������*R������C�<a'��!E"���A�*�\ zc��y�<٧.������@�d�VA��y�<�����6�
��ת��FبD�GęL�<�Q����<U��Çx��8�7(�J�<��D�#P1�D�h��� ���E�<��B�XBC.��Y��y���k�<q�!\�]~n̫�&)B�13O�i�<�a�ؿN%v9שϪ�����Ld�'������V v��r�O�Y��x��_G�!(���B�� 
�����J4�@��m<�	��]�RX���5���`�d��:2O��/"�)�ȓ2�5��C�~:���O/'t(��`7jP"����2K�}�v�0YN:D����ո$/D+q���푦���ȓGx���"By�~Y��dV�)#�ч�v�j �.ɜEI�l⡂64� ��'Ҥ`��кm�Y�E	ЙC����H-�ːe�6t[�h�2�֔!�Ԇ�uq�=�qV6D氁v�ÛU��؄ȓ{[��q��[�b��xaq�LD���i[DpҤ�D0c&<iA�*QO �� �R�#�@G�~1�uJ\3����N�¡٠O�#�\����Q�d�ȓk��`�L�0�l�S��;��i�ȓ-gvy��JN�i
�;�aղV^��Y���Q!^� ���ATeӹW{�̆�VV�0�ΫX��+��E3"ࡆ�2�}r .�0nQHl��茆,;����T��3�Ș=�&�b�6��ȓl�,�W��tN��f��2ojņȓJv"��	c%$ 1�������j)K��6����#3l����S�? X�1��s8*����(A���"Ot�gչ:F�( ��P���;�"OH���.�1�H��̐K�yi�"O��A��Ƅg�t �$��3� d��"O��c�@QBU�2���S#"O���6埀?���[F,\�w�r S�"OƼB,�9IL��V+��/����"OF!�gꁵ3��m�u�D�"T�8�"O
�yÈ���BMq#���l>��+�"OP��ghL H@PCT�P�;!�a0""O� ����I�6�bK��M�2�Se"O
��2/g�̀�ʁ���2 �Ym�<q�$�j�>@
4C�5���0GTu�<�历�jLă��ϦW2Bm°!y�<���V�@Ρ��J�8J�ǁ�P�<!�S9j���gX�/r@�p&�u�<��\;`���� �Ș3ցNw�<aG*�j�pH[�G�3}|�ى��o�<T�Y�:�b��t��,���I���g�[�{���B�>v����
+�:��H�B�ay�R�U֔t�s#�:FT��F̬3u��A����G�h�q!��^��O\�(g�'��
�������-�BΟ�A��b��ߧ<�ٓ-.��χ]�<�ۗ%ޒod�H�"�	f�ɧu��;uC8e����;�<� �A/al@�%���Q�R3�C ���7�#�$�]�B��� �%�48�VMA,Wڲ ��$D
� �[�C����S�=aE�X�g`D�[ra�{|T��St�zND�e�F����W��x ܣ=��0� �R/ژ;��
E��'$^�3s��)I�v�*�R��'0�|=�R%i�����	S�=���V(�L��61 P���1��Xi6�� i�M�tP��ˀ�Z�i���!HT��g�5J9�i�(�T����Z�
L>���$?�Z���T�sv�`TBL�Q'qP��``Zr�O8�t%��:ڴ~��E`�Mĩ��5@���v�x2+N���r2�ä`c�M�r�ς63�����g�:M2��T�'����`�I�[�J�Vu��
ڡ��:Ƽdﺤ��`Ei/���I Q7�H+����������j�"pG~R�Ӊ	���3aϛ	��#�ǃcb����/�,]g���^���^c��&҉ �xʁÄ!8�ZU��`�>	��i>�2e ޏ�� �Q��8>`��0'�CN0͘�aāS��I>��iԡSӚ��ƨL�r�,0��=1CI�,r�NEy6��5ohՀ���e��ШiG��(��AfȉhO���=�đ{'�����.l|!��K�%�H�s
(O�����o���O��I��L��� t��
�T�>��O� �D��p<1���D������XF�`�+��'PV� 3�O���#��)�f�A#�zL aE˄[|�e����[��x�4m�n�c����k, �1��%�q��%z��2���]f�[�'����Od����$�ON��D�w┌�4^
Z,k'�� %H��N8> B�&�$J��^~�B�ࡨՒv��hD "�	���1@p�4j缑��K/%�|a9�+�r�'���RF��C;�Bt�*缐�N<!!A��1�d��͓O|Z�1�*2R��(WGQp��=���%�	�P�]���~2Z���l��MK�X\�$h&EF�nӠ4H�Aܦ[�%���X�&�d��$��xOX�cqIػ|~�qY�c�WC�b�PcY?y�'o���T��/g�L��a�+<��0D �*	�_���%�S�]��Xc>���%c^�BKN`C�ߗ6��"��>Yv:O��'��5?�����P:<rȚc��.�����6I�΁�a�8��	4΀�e�>�����P.|�(`�=���R���Uݿd�|���Hb}�'h��fӈ%�����Qݟ$Y�'1~}�f�W���X;�F�'�i���')f~��瘕s��xD��OȐ6�"'�1�΀�c�����O8����0��)Cd&O����ԙ&����4۲=�����/���'�i��g$xs��$�TL�4$Z�/�����	�P5�°()����[�h����.���
P�� C� ��&S�t�?*���#��
u�ȢEH�"Z�y$(m�P td�{�&�P"pl�._��x$�ջw�`@���8�ɹ&���G��(p�@�@�T�~T<��?��B$b����L'S[��!�o"8��E&��q��U��T3$˂^a�*�,Qg��X��\2,���IJ?��C���q ��N��H�s�>~Z>��c'P����#)�.��
֦�A1�OI��R�g�1 t"?�2�er&O��<?B�z�cťRԼs��.'r�x2㝯UJ@R��A&>8kL�1&��a�*,n�K������'�T�bu�N�=����@��Nj�3��.T�����<N��-�p[�O"���J"pY�G/jan|Qn�NSqO� �e�VJĝL̪����8#�T�ިp�4���J	Q�20�&W��' 8Q��o�����_�
��!��0� ����a~�D��I18m�Q�R�O�B:dݘd�#4�׎h5��(�Kƭ	��q��nD���lU��҄@ƀ\Z���'���`T�B{�h�#fI�p��+O
�k����e�x����~���o��a��`	�IVi�2��b@�
��=�%�FT�iYEL�(9C��Bܼi��yA�A��$�C1�DkY "A�!~6C̜)u�6�3��0a�J�#�=��|����4{���T�Cl�J��t�E:_y���3��:5(Գ$`؅�j���KɄQ>џh�Tǂ�!�"驅��t�r���92�G�]~���T\)�y"�� i� �"�ؘQ�� �JJ9�	��Pro���I	*R.���$��{d>2��P�2<�p���l�L�Ɠx��E�V��R8p�l@��xi�3�I��p<���A"��=�2���*�k�ȝP$��[�\���'Ln|t	�L`z�P1%��x�����/R��T��c�b�z���ڠ@մ >�,p���?H<$��R[>�Ġ��cF�*��T@�$��H�PƇK_Mġ��kV�j9�U�'w���e�[1CJڕP�J�_#:h�wo
�ָ1��M)A���1�3,Od��]����1nd|�Q�L/p�d��Y��̙7Q�d}�U�\0vd�@�<�s�y�+,O2��S�@&/�\\��g�r<B�	�ٖĘwdة88�A�3�ξwn�@h�eYl?��
�i4v��S�Z;޸��wH��"����,��V�N�2���x6�u0��D����̙CӞ�i��U!]���Rȋ��O���VثH20�I��Z�֝x��	7e��Mȃ�R�Z)���Ю��O���C�#
¬��K�tuR�������ŗYO౻G�A�_:^�T&[�l��?t��3�\���<�qH^j&��3k����]�Q <\d��j�Zs�(�%Å\�������'��Hq��hL\9 ��>}�3��Ԑx�o�y�F�n�sۤ0�ňc9�љ�cT i!� 8�AI�؍;��OI	5�|��`�XwiێL�)��d\*�nY��Iz
�X��ιF����pǔ�9�>�BƋ-!/�kB��i7��C n��'�Lx�W��]�N�q8��t��/� �ўlqQ坣��BF�	}3�	"P?�1E^E���)v�J����Ya�1}R�ܵj�4;��'�*t��i�-��j�o�dg�T�p�iݼ�x�)3zLӅ���*�.T�2�'ݺ�Rg�')���㣓|~jI�vC���x���Hx�4��,�p��r/�`� ����C�>�i���*L7`	�z��)ɧ����/,��#���M&�	��q�l07�W`���O�e@D��%�i9�e�� ��mx�X H�y�L��/�2И��TI�� ��*�%j?"�	@�:�O��Ba���w�j �7�M8+�E�����P,Q��a����uL�&�(��sk�=:4E���<)���(�[�K�,�|pKu"��rZ<�'�ā|`�D���b(���O<���ʓ5U���i JۉR�|��*X�+-!��	Tr ���I>}�<����ԼUH0�B!�	Qi���y���X����DD��1Ok�Ѕ>+r�4d��]6���eB#D��}�mZ$�\뵮X�+��kS!@�3%�)UdOq�
Ժԥ���+�F9��H�J�b?	R5�J ���h�CTᐉ+��&�*FU*L�s��`j�"1���1Y��FӌI������!��'��9`M�"�ay�#\|p]ZWo�0��颠&���~��S���G%uٌm���Oz�b%4zZ�u��t�w�إi�!��ގn}�DAG��g8���I$:.����]�<It��y?�E��ʾ�����1��w����Ǌ0<��e���'D���'�������$T�EK	B��I�eX�<�n��"[C�Q�%��%���  ݊��Ț��Q��H=�f�;O2�'c"��� �@��/&8	J��ԏ)���P��(B&�rpB�^�L���*� �&lR
G����d�!G�H��K&�$�:UhD�����Hbq���&�>�9@�0i�}�?�4e�_���A�����EѐGQze��'��d(��Y�:A�ٙs���a��X�z�$�	$?���;ce|�)��:��	�g�����s�OQ"{:�TXC"O�1����P��e ֧�& �(�0��#��@ (�2��O�.�q�O& ��i$����Ѵ,yN�	w��M�8���,|O� ��e��
�έ�� 	1H�#��?z����UIQ������0�����{˓$��iѱ��1������_�p��?I���3�>�Ѧk�1p�x(c'��_��I.��t1q� l4 �I��j��E��z�����	7���1�-W*&��3F^K\Мr7E>c]r���h"��~b�w�(��L����D����R�e��'�b���E |�|ۄL���x�%F��0�̄9�<�|�
��_�/��O� ୉7I*8���Ba�,�*e��"O& �1�؉r��䘴:0m����"O���7o�J��ÁF�<'d���"O��1�I��p��$�ՄL�>���C�"O dↃR����/:�����"O�-Bnک{�fس G1�@D:Q"O�ċ3O�B��i�2"�7���"OL)�B�,R����a�Q�2��"O(���V�*@��n��}|f��"O��!4-�	�j��%�Ej��+w"OX��a!O0PG"T��杬d�0�"O��� U�D�,H�e�V��s$"Oм��� 
 -��cV�Z� m�"O��9c,H�7<؈�f�!sH|9�"O�$k'�)���qd_�hI#"O����!�� �r0��c� :QjT"O1"��K&*l
,�QHP� ��A:�"O�<���*-���p���c��-��"O�L*�J k��C��޿�fA��"Oja�hQ%-آ�� ߬nqB��"O�aY3�0E=�ؑEcC�M�~�bU"O� �BkY��#͏�f���RC"OD�V`�j��4��A�F���G"O�0 *[�vJ�ځa]8m��lۄ"O�i��2"��� ]2�n�<9g�Fn�NQ�%�U4L=�Ϝf�<aCm���(�@��/�P)e�a�<1��H=#d@��H�+s(\�`H�`�<atd�����Kq�Ͱ@]��k�*u�<!�1?�H�y�lQ(zҨ����r�<i""�_dBA��DפjR���)b�<qr�N�=��x��؟5P^�PV$	Z�<�4̔�p�xЈ���Phz�02LJ�<��.D�h�����!Q̑� bI�<!0���>s�1��VbB�4Hz�<Y6�Έ��`@���M�(��Z�<��ʚ��L���D�^>U���Y�<a�f�Ah�I�^{Ll�R�J�<���(~1�8�b�)��ZE��G�<a�j+B2�J�I+b������L�<�3�!3:"�ó�#R-@�!W�GH�<)� �	~�������3:�-j�'�D�<�B�$>�t����{VD�3�V�<��в%���ص�Mt�8��As�<��⑛ZƊ����&YH׈An�<�iA:~�(���j<ٸ,P�XU�<��F58�� Pwi���q�b�XP�<)�OY�0�,%��l0���@�<W�L�`��<�%�e5<���A~�<�����v�$ݘ���8uD����Xv�<AE�6@h
ЫϪNk�YJrp�<���8M>��d[?{T��G#�g�<��.+l�`����ו~����1�Hd�<�a���o��Ä�ޚ���a�U�<�s��)B��0��\�h���X�<1���/���m��,���c]K�<Y6St���ːN�q]Fxkt��_�<y�iE�����=Kv���fUX�<a&���g�>:���Pq�,k��AI�<q5(X623Z5hd'@V�|SfJ�}�<�+Tw�@��f��\R4b�e�<a��
���ZD�1��"��]I�<9�i�=;,D|!�c��}�Z�a��F�<q�MV�.���Ǔ!�� �P'��<� �q�F�t����E�9ބ�8e"O�3A�<bw�QP`%�2{zN`"O�3$�'u���x'�A���6"O�Pr@S9
����"�6�"OX�����09�Tl����:�.%at"O��Ɗ� 	��bTn�8a����"O𐳴�Mg������NP4D�t"O~)��n�5.Yj!��A��/?h�"O�Ȧ%�7�a����(+� �"O�q��G���$�Ωi��ͻ"O����e"ڵ������E"O���ASC����'s|��D"O2dZ�"��A���T�T���"O�0!�bW>h�H@�O�:0K�]I�"O�AI��N��a��WD<&ey�"O�mB祜+Dvԓ�@�.P�lȄ"O��[��L�%���âו`��<G"O�a�F�5���8�ύ
�(�9A"O���'H�*u�����2+�er�"O� ƫT%s `�բ�!{l�e"O�B����j�$ȫ��yЅH�"O$u��];o�`%�U��woh��T"O��1R��Q
Fѡ����.k��2"O�PP�,(L�1堒�,T�� U"O��z$S�_Pu�eV�~4ұ��"O�$�7�SR#����)�.�"O����CK�L��F�,�fy�"O�����	;eG�1]�}�`h��!�$��q�M+�_,roLp� �3�!�W�Y�$M����I��}J�nӺ6�!��Úx�B-"qfY�m�t� 2�	�p�!���∛�h«(��;�bT�D�!�<�5���9=�I;�&��!�d�.����g��ԩIgG�(�!��H�"Y�A�!��,Z�1�H�L'!�D�+�N�T.
�=�AHθr!�d�l�Xw�N��8Q�HO�C�!�D��7�t��� J���Ѣ�拕mj!�DD���A�k��=�dJ!�x�	
�'��$��B�<|���G.�t��	�'�����0y�j$a@hC0yi5�	�'�d�GjAd�f�gᘲ%��̱	�'nU�V�H����Pi��$E;�'X`  �g�4��7	��i�D���'��d�A���zA�WKQ�oI����'R,�Ã��+� �� /Nd2��		�'�0P@���D���n��]h���'2�u�C�!�e�BM�VI�'�xUj3g���a���B�t�S�'{����:>6�E��˧:��#�'O�<a��?C�̈$M25��d��'Ź�+�;\%6�yd��A_�l��'1D9���W����rkڈ?žd��'(^���JP�(5L��"�;R ��'���I��Q�	�rU�� �
f���c�'zM�����AV�$����'�R�3G��)oHyp&��xIz���',�!�'�-H�H�W�	9�����'�>�`#��/a��"W�Z�8r^�	�'e��JsB�j�;�+ƽbe��k�']�� "�&"�X��ҁD�_g��'���32.��0~���6���Z�܀@	�']��u��"@$n� ���x��'�p����&_�|	�&�O�J�S��� �T�W�%G�s3�%��8�"OB�#EL�19��%�5�xf"O�0�È
�^٥�T0p!X�1"O:���oTb��ƣl�h�"OX���Ϋ_�0�-^�Vb򱠄"O����b�*���X���5G�@��"O^qʐ)�i��,�"{]���0"Op�s��F({�v$��*ߝXV0�:P"OCL?/u�	g(������"O�ӡ�M�K�l�Iq���^�ЙP"O�8J7�
H �Y[�t����P"Ob�s��o�"�D���ѷ"On�RA�W�RFA�Gx���k�yb�֞@&�y�R�0�8U��¢�y�Ȋ�2As��Xhi���yr��5�
�x`��<\8�[�V��y�J  A�!"w���Ʊ��	G*�y�+�~�:DÃQ=S2HKgo�yR	Y@O�qcN�CR�l��̙�y� ��1����S�4B�6�{�o��y�A��/A�չG�R�8aZ�9�d]��y!_@�T+ �ճ3��9���2�y���{����M	1>\��RbȄ�_6��r��4CθzT!|�M�ȓ338���)��e<0�R�`_�>�$��C0i�D*+	��ebd��I�29��/�0 �fϙ���h��<�i�ȓOZ��	1�'S12�(0m�80䍄ȓ;3���uk��l��A�JC.!,���ȓy.��8��K�H��x��'jD��ȓBƀ$��l��`+X�P���=y\h��4P�(��iF�+�� U�7��ȓe���,�uN���+��u���(x[��U"q�3`kJT���\��}0��Z���ɻd�Y4\��+�����,�+B^�K�%�?PT��O��=�*���p���f��1�a���d�<�6���I؎�2�LQ�2���{�<i�
��M�&8k,�; (��JS��q�<I��X��5y l4mW8	�CI�<��60����@��0+��m�2��C�<1����>Lp
���-��R@�@�<y�CK\P��k���V!�D�<YRa\�1��Թ�� %2xt�"mJe�<�d��-�0�s那�<��"c�d�<�+�.( ����	�d�4d�(�^�<pS&	�ܘЭR�4��l�P�^A�<Q@�1����B��9�g�{�<�bh!U���a��Їڎ���z�<����~H�YM3Z-��k{�<11OH�t�k�˒"֪��g�A�<q#��%m̰�8%$� E�%�Wa��<��iR��}�+GX�Ȱ`Wx�<y�NգTsDMR%&Z8 ���v�<q��V�Z)豓k\z��Y���H�<��a4BC� $�,AU�E�x�ȓ7�H��g(?%��# G�k�d�ȓJ`�	A�˨j�|Q���&�R����t�6∹kqH�2���|y��HG@ĸQFL���bs�\�w�	�ȓ(��(W�58��xj�"��
�LQ�ȓn
����(��\o�H���[��\�ȓ}m@5P�7d�2���l�%!��<��"����A-ЩsF��QBf�#Hʕ��S�? ���7M�mcv}q�?7��i�"O`�5͒!��1X�e)�`��"O �TmT# ���K4�EU�Z�Æ"O�USO�ys�a��<:�dț�"O�M`C�mQ�!��Έ
:�����"Oh���ƴPg±��k�D��"O�� r��\Kv9��ˊi�"O�A4C�5nj��Tj�|��]��"OB��i	0Q��rC$�	
�luK�"O6���Bѿ:���ȖcT�>�
UB1"O6�q��U��t	 �	bT�I�"O�I����cvZ�2��D�Q��	�R"O|Yf/�'B�PX
Ԣ�k�&�*�"Ot��ī����k6Ǔ*N�A�g"O�ؠ��
tLN����Ev���S�"O�u��G�1g�l�U�L)%ǎكF"O���#��w�6};``ű]��Z3"O��E#�H���E� �4��"O�]���]&5�&䛠�� � �``"O脃��E��NC�T��"Ozذ��-E�H4�un(}�v�a"O�<C3�	X0Xu �M� 	�>�@E"O��6"E>N}&h�̓G����a"O�Ĺ��	�C�ꥊA��2@A �"Od�5;;B� vKYI6,��"O8`fh0H�1���x�X%P "O6H�Ȃ�i��E��<��y��"O�\���W�@��4���r�<�'q�i�.�T�13�N�?�
#�'�J@�s�V�&�b}R��mfT�`
�'�*�@X55+>��a�8�B�'�`�z4�>C�l,�@�_�OĜ�'D�){1�G	D1��@�H 9����'����%H�-bn�r'�qwQ��'�dL2#���?Ud-r�fI4W4MS�'LT��bS�uS���5K�:%�5��Z�1��lk칫���m�i�ȓ=��$kP	Y�Bjpvkś*Q(مȓRt���RC*U�У��?|vɅȓ	��v�J�,dz1��Rk��ąȓ�l��'��+/�^ ���^�v�=�ȓw�!e�S�H��+��]�(�ȓY4�x0��H~�Ltc��:�,��B�2�2GFX.�*�;�U
P�܄��<�8�[}�V,1�`��{����$Z��Q'/X�8���B7�q�ȓ�Z}��\�K0�8@m�h8�=��lX��s��_GD��AF�	�@��6j���Vhәx���"S9�<��#ᒸ����%�h��À#5f���3� =�$a�1q��w.��6�l)��w[ơhŇ��kJ���f�]9�ȓ0r>�q�K��9���@�"	�)�ȓ%X�ly��k�8���+BU�Մȓdl)�ܽ1N��2�N�%x��؄ȓ0�<lbA��2s\���@tk���ȓ�XH����P���0��*��ȓZG,���8C��S&�D(���I�qPi��sw���%�@�T��y�����̳wL��c�5�d���<f���.�����|:Ȅ�����3/D�C+��9��ʝ@��م�-M�0q�%R��9)�:����<>N�P�mՄA7HɰW�R�f�v���S�? �\:��3:`��iA�F�BK0E"O|C�� ,aZ�i��WC�q5"OzM�W)��.�Ⲡ �I&�9A�"O��%�
l�Ha������@�"O((9�AV����!�iY�����"O��I����$І�%4``\;"O�8P��Y� ƀ��b\�G^�(�`"O�U�4���X�8BG��2Z"���"O>]�% �._�(%D�W% i4)��"O`��+ǈA9lp���fha��"OXM��w<�T*��ޥB��ĳq"O
�hS
�;�X� �W�u�.��&"O����C�:~��
��u��X"O������eRHEqB� �� �"OpE���ZU�'c߸!�z�:�"OIذ�N�G�MX�AZ��0��"O����بd�, S�RM�2"OP���o ?g�eض/#���S"O�M{r�Q�K����#�
�i*s"O��IWD�]+@D���ߟ.��� �"Oz��S�ִo�2���L�u�8�:�"Op���e�u���@�]C�"O���$�դ��H��f%��"O���$���^0�i'���m�u�"O��B�T3�<�th�XZ�� "O�eH��P7X���RM�>MNdT��"O�a��E>]@�X�K65t��"O�|��d ?I�Nm+���E��Iڅ"OYY��	4H������[5[�n���"O.��4%�
q� j�MP�Y�qە�Il����T;d��A���w�0�Ϙ A!�ŀ.���{5#=P,�e�V'3����S��y�ĳ�J�s2d��|!R���cY��y&^���[C&�.n��������HOf��DW(i�p��3A� �����^9Aq!���AθH�2���9C*@��È9e��
O����f�@-!��9s:5�&�'~�1 >�Ui����kE��ԗh�<a�a��@�d��%^;���#�Qt̓�y���i�X�d1$�<E�f��GOK5#]!�d�'SG�5)�cǓ(>�t���1U!�DQ�?�A�FfC�R5lX���_�C��,�� 
���HV�EߐB䉁b�"���Q�&Bո�C�9��Q
$����A�/S�?I�B�ocYa�0��0�3��>d��B�ɘ$�0�@j�[�t���ӫ-�C�ɡ{V�q)fD_,J�xL"af�G��B�I�DH0�r�]�<D���T�q�B�	�!��u�Dd\*8�2 �"��?�B�	+��3F��;����/ڊ�C�	�^�I��kK.C�����aW7k�B�;���y�&ۂm�T�h�c;Gp�B�I*^� �҇�"O�����kEtB�	�:��<�3K�@�S�A� �B�!inΝ���7-3�r6�$��C䉢M�������"a�9 ��],"��<���T>E �@�!"�X���HΪ�6�?D�\��ĳq����ue�ʔ�"�b>D��{�Z�l9��P�!Ѷ.[J��3/}"�)�Ӵac��!%c�X{��zc����B�ɂ4Ң$� Nβ*�!�6Ĺ �B�x�Z|��A1@�y���8T��B��)g����MOj��eбEJ�B�)� �9	�[.#$d��jʜ	Gp�(�"O�!1�I���)h�KW"Xc��Q���q��(߯Xh�8�R�ՠ�N9[�6D��{3�HR���fһ}QN��"�4D�h�tm��<d^	b��c�8m���,D�܈L'E�Q� �M-_x�m��+�O��OH�i���f�P�b���ڵ #"O����1z�"H���j�`(`�"O<��R�M�촸�n\>J�l���"O04FA��.Ɇ�y$M�90Xh�w��X�O����d�3�����9�2���'7D�Vi[�#�P�R�F��Y�
��M<����;�Iv��;Eʁ�[�������+:�pC��QP �r���8��i�./�hC�Ɋup�e�nX�u&��A,Μ��B�	6�-{e��� �⃬�8�B�	9-z�9��	&�%�HV�~B�I OS,JRb	�m��͙ H�C�I
+�J��'aӂ���ʡ!�s.�B�I�:¦!C���3?2Fk�9IBC�><l��3��^n�Y*��\�z�'�a}�]�/T"W��*6>`���yR$-.T�jW���Y4J±�y P����fL�}1<�1�,��0?)��'�&�h,�E�5)t0�̬('vB�	�.���:eG0H�q˓�ҏ<-NB��)e�Ġ@�Ɖ�3h��K�"�%�C��>#�6-�3�B�g�l�˄kO!m�B�ɺ[l����_�8�1SK��SJC�	�Jx����٢{� �e�O�8�C�Ic�6�[��h\I9�N�c���D+�	s[�0�`~�8��'.V, ��B�Ƀ~v(Aɦm��"�����B�I�q,�����SQ�k�jQ�A(�B�Ir�2,��ӂlРse�A�=lRC�	>\5q�DQ}���1l�8T7|B�I�_�7��9u�҄��-	D��B�I\��A�qMJ��D��B�I�"��t9��ci�� K6E�C������'Xl;���1Az�#=a��T?��Ϝ$%�8"���`�p��B:D�!�[�}�ȑ��Ǚ�uX�g7D�4KB��?E����eG�n
�y�g�'D��I�9��=�v4м� K+}��)���bg����^C)���1F�B�Ʉ��Ȁ��ғv�)��
�6udC�I��Ԅ���S���H�k�cd�?���I�:DY�x�������.>�!�D^qԸ6��ƅг��!�d�G�`MۡɆ�ì�z��	���gӮYkD�.4��A�S����A"O�Dj'*��/�H:��'b �$"O���@��{�����e��V�J%3s�x��'T��cG؅iN�ycU�t��'S�E �!J�\K+cQ\���$�$D�P�1b���A�IζF� H��'0D��R�ݢu}��ڰ���R��QXu'-D����#�2&r\ A	�[ M���>����S�o�8�2�	�n�
UDۄ��B�	g�~�
��&�Ӄ�����C�	�g��p�ת��R]����:�C��-���ͅ+2:45�"�S4+��C��
Kfh1$�1�2I����!�C�6Kw�+�I��oX8��"��g��C�)� .��$�8�9ˑB�e�n$��"O��aƧn#�-���C�����OX�dS�,�R�[���'����A0;�!���PB��f����-�@Ҍ�!��ԷIV�q���ڷ}���:�@�!�DE�D��`t�+)�nT;���!�������w��9B��p����Py�"��IuD���@N�IO�Q����yr��
x�R�ĨI	
��1�ҥ���y��.�Q`[�ޜ\so֯�y�&��GON̈5�������y�O�"G� I9$ٱbE�
�y�F)?bQ ō_���ũ����y2�;�T9!�I�	ᆬ�'^��y� Ϛ]�Bh�&�����Â��y��J -�<A��Y.~،�����y"�F4M���y���2<�JD���yR�V4ܨ%�e�.(� ��cnZ�y��V�O�j�c�I�/:P�&�yb���H��4#�/io��x�X��y��٣x\\u�C�^��qptjȿ�y2�\~�4� GG$X������y� �>|�©QP���=ܐ1"`'���y�ᕍf�TH��l��>�(�w��y�jЖe�P,w��J?�G ���yR���bu�Ԋ���,y��G��y��Z�I��u�5b��UD���Ґ�yRF@�n> }��h<�f�%��y"�!	Ң`���ů3I��{t���yBL�4��x��[���������yRf��4��X`�*�	
��G�Y*�y�EL-7_��y�F�7JV��7��:�y��>B!�t	�� �
�+�쉖�y�	�(_dF�PC�z-J�� D�y�i�2��A$fJ5[<h��sm��yBJ�[�D�R@�(D��بRIL��y���(l\pJ�MQ61�!�䔀�y�e�6_���-��/~v��Ȏ�y�͋~�H)S����(O������-�yr�M��#�	�V ���1�y2� >\ �@AҁF�F}�����ߋ�y"��+d�=����6nD�jva���yf����BS,^Ĉ�R��Y"�y��X�O����Ϟ"\��`�����y��P�<�ac��^.Y{~D�5�U$�yR4 ��m�V|P���O��y���/��Bfœ�p���J$I��yZ)Y�`zpA��|���e�;y]�B�H�N%���تP6p�R!MʳY�xC�I�= Bأ�B\Jv�Ơ�2t/�C��!7�,`�s"��<ɲ�M�r>�C��6_Ex�2'��'�\qGB
�1W�B�I;P��� ���8�ڤ�f&۵w�B��4?�$ic'kֈT��l
�b�$-CfB䉲N�8Ų���'HO����`���C�	))���+c'�'_)�AR��+W��B�Ia���6�W�O�H(���	F��C�0�j��uiY�@�8܃�ɑfXHC�	
pT�6A�E�%�ŋ��C��|�`9(VH�����J�K���C�	{�J�*���k�ᤤV7\*�B�	�8XND��.ПRf�y�E��x�C�D	ʩ�A��
���3KW�o;>C�	`�����Z�ȹ��٢w�C�)� ��@�܁d���	��K����"O�5��LO_.�3(X#;�b!X!"O\1��)I �@��T�+�B,�"OB�������a���-�X�"O��2Ԋ�.��=���h��f"O���� 6/k���G\�.�f��a"O
ɂ�o-wP��*#'Z	#ipt�Q"O��kP�/,� )����>X����"O8Hjr
G�D�S�U2NBzIHC"ONyxG��3n�p���ʛ.\���R"O4	 ��dِfᔶ]l����"Oހ���R.4]�)��W�_x LZf"O�DgHB%��z2D�WT0�e"O���&�H�IM8)��Ñ2{�4A�S"O q�`Ӓl��$���S��D̂R"O�@AJ�%z;�}"�A��$FRpSG"O.��5�^&X�� ���C'|��"Oz����Ӽ�|y�E��u|��"O��#B_'61�E�"E��=��*�"O�M 6b(i������8 I�[g"O�}Q����ƕ2��`:����"O��Qd ��0,y`F�y7ތ)"O�4Õ��sטU0��L '�I�"OB�pk�9�h�r#X&���p�"O��4NK V����H�-�T�"OZT�2�ü%%���gAʊt�N|�"O2h8���LE�Q2ሀwm��Ȗ"O������/�8��O�69T4Hc�"O2��,�aOd�-�<>��X#"O�m���)9��"���H0k0"O:.���AW�j����3�X�[�!�$�6Z����4��"]�T9�k��V|!�d�;x����C㜓�PͫRO� Q!�$�) .ͱ���:�� �wm�b!�����ST�~��ɉ��[� ;!�DW�<���Pm	8u�P��,!�W#A040w�?+�NH�Ʈ[/!�U���h�s������DoM!�$�#��hP�С� a�VG'>!�31����`�6� `�0���!�H)��J���3X�����iT��!�
�{4����Ƥa��\�!)R�-�!�)��ms�o_&j�L%8��I%�!�$�tG\e"��� R��t��&R�4�!��<FUZ�YPC\��l�*qe��!�D�:ln��"�HE�yxJ<seU51�!��U%.�;��J5Y���4��
4�!��6`��(X���x��Y�r�!�$B�B6����_!وԐ��%�!�$	���$S	L#mt���2؆N�!�dZ�+��!�as@q���իh!�P)^T�&�B�CYn<�E+�='^!�¼=l����D�QOHp��N:6U!�d0+Ѐ��6��W���+�,�G!�Di�ta�f��4�� 5]	<!��AH��H2�.�&/Ѭ��嫗�#!��ύI�DkcM����8;ed��Z_!�D�&H|����^�"�
�*[~!�Y��0�an�S�Z͓PHx!�D�����Q�ߓ_����B��9Z!򄎳`��MY�k�:X������!�D*f��(� Ƒ$fT� 
���!�d�$���/W�8�H̱v!�d��$�(����80ahZ�8i!�� �ధ�!j��J�/\~px��"O =���!;ؔ@1�U�bh�9id"ON5)GFH�*<>��b�,v_�0�"O�|���Z�v;��17ZdiR"O�H��Ǭ^��	�+_9vw�e�"O40hժ��Cc� P�� ]g���"OVu��+�*�z��!�A�J��"O��VM�bV�q��5��@�"O�(����#H�1��_�XԈE�"O��
�-�:'7�"@䌝9(�q��"ON$�00%�L�3�D���"O�H��;Eq��튫Q��q �"O8��p�H! ��#���b���p0"O�@�5dH?���_�#��j�"O���W |)�l�v ]3}��"O�e{�Írt���O�yə"O�l)ַY�p�W(S�%s��"O|[4'�p�.���ނ$�(��b"O|(捍9�8����p�F��"Ov�H�IY�Kw.]"�lֹy׮��a"O�P��ӞX�az�KP�Ѧ��"O�"ĉ!G\P,A1�)C~:#"Ode��
�蜹E��N���c"O\P�gW�\P�*
�?�8m�T"O~�S��vCmQ&�	X�dja"O(�Ӈ��Z\��&Ƅ-5��Y�"O"���dR�&e�x8��ʶi�2l:�"O>c��OkĵR5�Ъ7Ҟ�c�"O���H#�BP��W�fi�re"O$M��`Ӟb�`�J�-�.:
"O<�3���-?�\(Ĭ'.6�Y�"O�$
��R�K�ޅӦ� n4�I"O���P���l5����żH@rlBE"Ot�GM��l*�ȫe��N�>�Zp"O�1�QFC7 Q t�3P�|��0"O���Ҙ7�x�BFK��a����R"O�q!cU\p��X�cȌ?@H�"OD�;e���F�6����2"O����'ɀ@�|�c"�5+���"O��kd#�غ�Ъ�Pr�9�%"O���fL�PKd�c�?�ݩ"ONd���]��a��,\8'�2P"Of�ଓ�#'@MZr%��B��Ii"OuP0�F�Ҡp�"F C�p�r�"O<]b���;��c�n�#i e�"O��i�&�� �!�n��Y`�tx!"O~�A�O��L⥋2�� )n�Q"O�=��gDh+�kF���S�"O�15b��j��;��.�l��"O����L-wwb4��&�7��q�"OIP���[NF��P��F�0�c�"Oh��3욷U�uy�`^*0��ݙ�"Op��Ə�6u��/�e}r�x�"O�Y�È�%/���:F�V�X��u;"O@EkJ� �|�����\j|�"O��Zu&UB�l0;ƌѧMf�	Ku"OB�H��!9����썈_Y�x��"O�x��dX0��I%��M>R�C�"O�DS�ŕ�Ё�"C�"E��k�"O~���OƳvAx��W���w8R�� "O���پ5�j�2���J*����"O�ԯ�y�c4�@$��%"O�u�6�)��U�-��
��(�B"Oj��'Ɔ)@�����H�ٶ�@$"O� R���_��i*j�d�&Dr�"O�t��f!��J��ϋɈ���"O�}�F�%dUr��5h�7Ô��"O����ެ �rY3��Э}���"O�(�c@�a!ȹX�M ;E����#"O*M��ɜ1�Ntʧ�^�~�p0��"O~�ʕ�B+;���Ѭʙ�2(� "OFmC*@�U���P�H3�6�j"O��k��߭PvR%��ʄ�a,e�G"OF������m2��^R~�H�"O������2`���+^�0f�H"�"O�}��-��L�X� N>AR$�rg"O�y�KŊfi� ��@K#(cp3�"Ot�I7�ѳ$a��xJ��wmx8؀"O��'��;H������RRp��E"O�j�J� V�n���M�([�\��"O����jB-���㐭ۀ(X�D�0"O�<��jO�Js$M�'�B�m�R��"O��b1�D�4�����W�E���a"O��a �ׯ8�Ĭ�΍-^���
$"O�s��x�j��ӵ��@��"O�)�!��JȄ������4�r��&"O����F5����(W�4�D�"O4}P��?�JlJ5�37��	)!"O��3���	x<�ah	=NB�Ó"O<��F;a;�����ԡGr,)�"O̕�ǎ&kʐ��E�/j���"O\�����:t iYR�?a�&I�b"O�P�%��,3���y�`�)��iQq"O�h:�*� `��!#b�Y�`���f"OBa�MR�`��;�e�y&��4"O�qg�Q7S���)��<<R�xp"Of1)��^0B�᱔цbNVԒs"O�qY�c�x�(�p��vC^�j@"ObzV�F8J���Y� 2P�C�"O̘�d�O�8n���D�S����`�"O�X�샂G����m��R�����"O�P"�ρ*�԰�ū��)�JP� "O	�̐�l�^�f ��p�*i��"O���� bQR(��M��~����0"O�ESs'P�
���y��R�vLI"O晀QC���4(p�e��:�"O���eGF�IdhM�v�ǍQG���"O@1
dٿ��zB�4*5�X@"O�,cs,���(���K�&��%ӑ"O�J��N�N>�P'�=fr�90"OXq�.��b�(�"v-a #5"O ����������sc�BX�=#b"O���2ˏY�h�!�F�QSr��"O��3P㊙# \��GU]���b�"O�8��u�Fl�%ŜjܲH�d"O"Y!�!*nhy�%��_�l�ۗ"Od���+�,�@���t��	�"O�!Ys%(e<d�f�
~�\!��"O~����� ��m�uKj��|�"ON� B��\g*lQ�K�g��qI�"O���F��u
D9I`)���yb���H^i����%Ǿi�h�ȓ=  PY�A�2Pp�	���W�ņ�F#d��iS8whB��j���Y�ȓ��1���!���iO�T򚕆�sF�!�ʹ.
���?�.8��*�x�9�gס�����B��<o�ȓe�8]���QZ|���U�15DM��S�? P<1A�S z}��0�[�h C�"Oj��b%��pr�C������"O�@X���?�8Kg�F�9��D��"O��8���O'2� AKC�`!�"O��"vW���\pPiX4��I*�"O��+��_��XQ�NA��A�"O��{�O�6O8�|"DX9%�L��%"O8@�uC1EE&I�"َIԀ��"O��+�
7KѼ���`(7<�9h3"O�cCa�%�!ӯ��-4�Uj�"O�pٰ�(8T8�٦i�_h��"O�iь�nY"��I�B�ޝh"O2t�g��Y!PɁ���5�^02�"O����v#E�9����4"O��Ȳ��d�~l���(O+�X�"O�<j�M�L�0uPCk�v�ې"O
��"Ӛ5�p�be���M%"O4<Q��P,/��D��Աev��"O(�a��qHR�M�$\��F"O��bd���4���#� n��P�u"O9���lx��r�L���cb"O}y�"�tm�u;/]�g�F|y�"O*�҆!=xBܸ����;��ّ"O��j	l��͈C�&����"O��SG!�����GWCtIC�N�<�ЇI5IT�H��-`�0�(�IJ�<	"��|m���
/�����H�I�<� �W9M*��B<xP�ZS�_m�<���!�B��/�2��e�C�<�U@2<	�A!U�A�s���"��y�<�$Z$drX��dH�Fn��"�t�<�ωUrɫPGT.�Xő�K�s�<���++2h[P��?\����q�<q�|�la`C��f�@TR�<yCÒ�h2�`#S���Q���;�#\K�<� ��,H$�h;��,p:�=9�#�}�<QVh�F���E��u�JdS2��S�<9D��I%�ј$mҰJ7u���SM�<AQ�K�k��
�f�B�P���DI�<ї��S���J#B(�)�5`�F�<1�LK{tD�@�,9zL-�V�C�<���]6��A�	�9���A+NW�<�@�'��=y�j� 2( ҆�HH�<qb\�\�<E�G��!Z�Ja���B|�<q�� Jp0���5L�^� ]��C�	�k���:�捉DbP�yEC�g��C�?u�|tc����xO0��dE�~�B�I��Bc���B �cە2�~B�4eC豲�>tbt����!h/"B�
�j��u/]�s'N	���	��B� M��xQ�
㌕ЖMP�T1�B�ɤ=�f��)��,�t]+2�Z<|B�	��h��E��0ܤ�pF;� B�	�G�9!C��f��x�����C�Z����MS?[t�R�E�T�C�	Q���(���;"nxq�d{�B�;|�9�	��V��,N�o��C�	/>��Q��n����i��F&hB�I�@�sęh��Xb*L/�NB�^XT�iQ X�}�`��tj�)^�C䉈愭��@��i�^m"�+�"L�C�"�V��C�ҹN�t ���C-- B��!LXnT�Џ��-�� � w1�B�I%4�X�p��?w�buqeh
�_/vB�)� b�#%`�.7�&�z�$X
D��"O>Qk5�A	A���qЁ[ u	"<�F"O��{'���OpF]H���v��I�"O�]�4v���H����<�|�h�"OhUQ�N�.�С���Fz��Q""O�u�c�tzT����T�T�5"O��A/9����A�e��T"�"O����.�	J��R2<D�|�"O�q�d'7F�
GK@��=`x��$���R膴LP\M��M�Ah�)��P��N{��I�p	�<�ȓNe.<2�JS	�irg�ڄw��e�ȓk����زYt&PU���?G\�ȓ0U`� v*ʍd�Z)¡�Y�$n��50�̩Sn�(Az�]�G	��~�t��ȓ0{�1�"G�Bʵd͉�� �ȓs����@ L`�̡���U�Ƙ݄ȓ{��͉"�� W�:��5�C�f�ȓk~�B��ڱb�0���T�2��`��@��4��e1$y��]�1X@�����)W턞T@���u�ܿ9~T��T���H�	�^��`[6�غ5���}m��̇�mZDW��1f��a�ȓx��|��G��
+Ï՘�E��|I�(���01'0p�ä�J�P��ȓI��:
���"fV>w�E�-�e�<Yw�-_:�b'_�&�h!���a�<���
���hAj��J],�B��B�<�@+E�R|̬{�%�Q)@��KZG�<! ��/�8��$��'q$\�'��J�<1$��|���1��V%+�T�b#�A�<�"E�+^�]�!`�M�
���iLz�<yn�'z��1�Veb����!Ɉs�<A���"��I��\�a�[X�<1Ё�hIƐK��3����i�U�<	��+}�|U؁'M�
JLXT�Ox�<1�Ǟ�}E�2tb[�F��s&i�w�<Q�'�m��x�Ġ�c��a��,m�<i��I���P!2Cƒ���e�<	�� \�欩2@K�s�t �0�^b�<�VO��^2U(f�O0_�l��*�[�<��,�
(����!ˈ!��x�e&S]�<����Z3�=3FjO�HW��B%��[�<����b"z�����5��T�6#�Y�<�pkͧ&T� j&���-�^Q�ǃn�<��)BI�ȉ��(HLb�T���Bl�<�rk=F1�:�P: A�I*#�Nh�<���ziN-�-ϳ"d�ѩġ�`�<�S�*,%������ �!���x�<�C�J#.K���uES�<�!��^vz��q$"Pdi� ��I�!��^pJ�	4&�$�˶�!!򤊗
�M3��q����V1	!���6lR.P�c ���,̆�Pyrȑi�h��A�:
� ������y�)ޅ�
�ڔj\y��2�ײ�y�BD�g���sB-�l��!�u˜=�yB���w���C�f�"��LT(�yr��^6��IPgנ[m�}r���y	
�AG����2~��3��W��y�e�<:}8y�a�ǐAL�y�ɓ�y2BȖ+�H�b�>c<T��I�'�y���ji�E�cDC�t��)WdA/�y�# t�.��"�ހ{@E�S���y
� ��a�G�p
P�q��Xj�؃C"Od�A"� [ y��)K�ء� "O��TJ� @j���)��)x�1��"O�R�J�'L�!�N�u����"O�p20Ƅ�_��bN�Z��s�"O�Hc`#ț^��T S�,)�X��a"O*�zZ����ƨ��a��8�v�˱�y"&T�6&��,[\_j�Xg��2�yB�[}�����Y�&(�F��(�y�e�uʁ��Á/�PL+#�>�y���q����/8`d��A ��y�'��g��y��4'~y�!��#�y�
�0��,Y��$#Er�4�X�y�F�xR�af'ġІ�)D�G��yR�3�h����}XL*��y%��u���k� �rѠ|;�
׃�yra٠!���!�Di�D�	%���y�ύ1=�F@[�(@&Z'�i3e�#�yoø-H"�3�ݶWR<L����y��)U�Сh��� B��f����yR#/?�8��(/8�*�`�.�y�E� J�b�M]��9Z�>�y�J�1��u�a,��'�2H��y��©r�*a-C0	��@A�A�yh�W!ԁ��(N��Z�e���y�%K�>�LcDU# �mz@�̡�y��{�N0�@*)|b�U�H�4�y�(��e��@C�'p�u9�(�y��ۢ�Nt��kֵ`G6H)F?�y�Ś UF��i0"GY,�ta`�+�y�R3#EX �c��=.��F��yҧK�VoXI�#��)e:���(_��y�;B��e����匀8I��y��&>�,����[�p����C��y"j���0qn[�:�����G�y�喎I������7g������yr�]�M�q��M8#�rL`�"��Py��ʸ.�����O	T�)q�Og�<�rL2M��P� �9,K�̰�b�<�
�
)a�m��ǆ�*��i�hx�<)�bB:� �%�G=�dPv@�w�<	��� u>ƙؓ���^P!U r�<a`�>x"0��Sj�`��o�<�ŒE��œ�,)���Lh�<9����j��@���,e����I�<)0���z�Y��R#��s2dSF�<�뚓X���`ѡ\�ge���#~�<9$�	� -2����$c�<���A%��8�ÅQ+CBA��^�<)�χ�/�<�u�T?-Y��6��X�<�o�zD��A��)�@����U�<�g#]�C���C��Um��0�A�P�<y�A�� p8�K�ů�dp 4��N�<yg�J��19"���|�}� ��H�<��&;;B����)z� 1��o�I�<q0��;xQ`�QA�"["t+�-�z�<�d�B꺀�3)H7x;*Ѩ��l�<�U���~���\��1b�fEg�<	S���,��D��4���y��j�<QC.� d����%�ҭI�fi�f�<!�D��0f�2jؔ;(��Ȥ!�f�<��烾L.��bF_�L٠�Cb�<!��wgp)�eqs�8G�b�<I�� �I��\I�jl�d�h0DZ�<� v���X�|\��Ѝ%��[�"O<����E�[I���/�5@� M� "O�	�T�&��M1� NS~� "O0�{��M�>�R��]�R�$�"O"H"��<4���Ȗ���m �"O�س�а�PHg�,8����v"O�����)_�<�4P;B�,�b�"O=� l0T��� t	C�Z�x�"O<���ǌ'-���B�7�Fcs"OD,"�
Ī:��H�щ]�h�~��6"O�����8M��H��4o����"O <�TKE(��(�gH�	�~�j2"O�� O��ot���`T)`dT��T"O�ab�cN�$�r������� ʇ"O��H&�9�B��1��s����"O& c2ıT��!�1s���g"O��s O 3�<�X�bt_�t�""O���b�����a��-s ѳ�"OF8j� �!��8C�+=��q�V"O:5����-�	�B~�a"O��K��Lp@T�!�W�qJ��"ON�8Vm�)(���Ys���J�K���y�B�_>X�gƄ�0��\ʓ)ʠ�y�O�>Wh�1��<y{�u���,�y
&[>~!�ߐC���B��-�y����p�*G��70��_ �y�8jf�{� �?�P�g��yl\O��p�-�d����5�N��yb�ۯ,r�0W�2R�ґ0��y�*�n[��3P�۟RZ����y�D��83�C��V+C*쳂����yRKF�Rv�A�A�ɖ=&�������y��G)d���;G�T7*!Z�`��O���OP����[�9 @���P��S�
\�'X�y�F�Fq6���!&�$�Ň���y2mY�Ռ�pa� z��P�C�y���+? �
�'�ŀT��L܈�y�CP��cB���{�ƼKC��y���=�ΰ�B�b��r�lO�y�Ĉ�7��$Z#��`q����D-��O`��7��|�g��.U��A/p�t��+��<1��� P�D(ȅ(��LLr�Q#Ǔ��B�I�Tm���WIش/��i{��{�lB䉖X��*�&�H�N�R2(Rg�hB�	B���1Ƈ��S�(��I�wBB�I�Rv����vS�	�ŁY�(2B�	NYl��5���3}�u9�G >�">q��h�$�שѨ �8�!�%6x�P�v"O*Ix�BD"*Ѱ�ϩ]p��"O~��$��AH	��F
g/FL $"OhU�� �;�Y	-ȟ.��S"O�)��;KK֡�P57.��'"O�<��"�;����' Ōg
a "O�@#�$Sg�I�e�ڵ)>�b�'r�O�QB
S�302�bb�Y:~b"O�kGaK�92�k�GA�E�H�)�"O����@����34 �,nʹx"OP���L���*�֮T��|�#"O]�" !"vvU���̈́*pV���"O*MҐ�6R��Q��I�^�0s"OdUx�Q����4
�pq+���y��'�O�b�I�_�(�`���;S2:��Ï�
�,�Iß��E�S�Ovx-3�±:1���s<#(���'��e��(��?�Ure���!��� �\��e^�4��1���P�Djš�"O>��i�@�:=��_>p{.I "O�����Z�J����%j\:�ȕ"O �۔Ó6ly�i��GI�5X�MA"O"h�P�S�A�jaǌ�U촫��$?�ŞYZ��"��&j�r�ږ�� �*����?iiI������3D���{�!G��$�Oh�S�g̓< �Ȳ��
->@Q(����.V"��ȓ9b 8�b>"�0��!��;P��ȓ*� �'�B"�(�e��n�e�ȓ2)�����I�5V	� �ˢ?�
����ş�?��� ����O2�H�̋H�<���īM�&$iG`Z6)G���[Y�<٦�e�R�xD�b����'JP�<I�LԏJ����k��iDw�d�<9���;7Z���^�N��4y�,Ya�<_iÊ�E-B4T����y{!�dJ� HP�h�;��형�,Tt���'��}�!EK�JƎ�
���?ql�2��O4�P%������R�n<�qF�:��P�.�`�I�oaj�)%	R9@��[r���ej���IOyRZ��E��\�H��Ijԍ� �偑�O/�y��\6:c@�j'H�^�!��_��y��M�:	�<13�։_`�w ���y�7!|���J�'[�,�7�(�0=1����*n���F ��]�hi����y�-r��` �ҳY��=����y���<���S��:D_4e���ؖ�y����z�!�F��Lf�@�0����yRfE@,�Ee�E�T��h�y���#	�$��Ǐ�f�^�Qt@���yR���4�\P��G/Z�~P+%P#�yfE&S2�`*^�MyD|���3�y2�������� �CH�)�2�x�'w���V�3Zȁ3OS"W"d��'��'���]y����\ߴ0��ɶQSX�3� �MN!�DS�y8�1Wb�D�61yя�-D!��G?�� ���^i4��%J3.)!�$W��P�7j@`�WJD;!�D� ��r��ͼs����
�>!�^�~>�p�J��ޘ�6��k\!��Z�u��	�G�V("�M�4*!�	g�J�!��ӣ�� Z�,];a9!��CQ�8!�v�����![Ƌ�n/!�D�� Na�(=��=��4I!��P�t��T�&�ѩxk����+4	��F��W�P�RpQ�a�>+��Q����O����Ch S�F�6;PE��aUl!�dY�GK���A��9F`
Ѯ�8`�$�O��d�<Y.O�I-�$��m�D��QV�p��5��+2�!�D���tj�ܳ8�N�C"̘RF!�d�2D����*�j�rЋ�;!�d�1�jѣb�H0V��WK�&az���[9o�h��D]���;poߙRB��vx��)����P7���'>���[F�z����I�O��I1�s��Ak���1�C�IV���h�D
$zl2�׆g�C�I�p����CfHI,p��w���iTC�.�zĲ�HӵG;��C=�RC�	M�6 � ߖ�,�1��UC�I�r�|H ��(�\ ѢI�7V��B�ɬk�\���.ЯE�r�� *�'z�C����8p��H�'N2�Gԛ �����q���	��?��h;� ��l�'��!C0���y
� �1p6�ÿM�&�rc�ʵ	y""O|\���y�u��fÍY���"O���fbb˞�{І�%��Mc 9OԢ=�O��'bq9�P�|7
�I��X۶��ۘ'�I���O���Y4��@�&����A�*���'����� y��8�
��	�M!�O0��'�)§S��`��HT�`�B�w�vE��y������sjZ`8�/��p���dL���RHV�^Uȗ!G5Q�$X�ȓI��t�\b^TTx�/
5	w��ȓk��0!$��!�xMh3�>l �ȓ���b�m��`���-ɇ� C��s`�U>7��-X���q�,�ȓw�6+`�*Zm�Dc��d����d�9�fM��tc�/˲X���ȓvJ8�3�:2�ܥ�W�Q�#kd���~9>Y�eC�1j�hV��/]mhi����s�|Ѣ�80J�`�t`ŤzӆH�1�6D�p�E���'B�`BX:�H5D�p(u�ئ$th%C�J�+$z�M'D��0���;"h=C�U?�9�U�/D��{�`�4=���0�RoK�!��J1D��@lZ�Y�TŰ�@["!`ݻ�k/D��@p�.
��-�3XK�f�!�#D����3w�E�ŇW�o3�A��$D��f�ƨ2�|ˁHԯ'b�BM=D��1J]�`����Sr:����E>D�H�'�܃�a;!��'c���0�(:D�lQ�<l*& YV�'X�R0n5D�1�dAQ��(�jQ_�-���4D��8����U����cKC�r�Qd,6�����(�΂3\,�;a$@0h�	9S�	mx�@�b�-�d 뱌P`u�1D�P!$a�hx`˃��r	���/�yR ��r�$9�ҏ\���1�u����y���`�� ��"�$�X�K��ybf�,>DY��_�������y"C0�Z$��1�.9��Z��$�Od��$��wNqfӧ#�H4L�*���D����䫴�T�$X�� T11���T"O�=��o��F�B&�ҵx
l��"Ofur�#�7��L��
�Sy4�
�"OdDspbևX�|�붦٦(ʲV"O�K�e[�up,!'`�8.�X)�"O
�*�范?�D蒤Kt�٣�������?�̍��ɛ�
��:�K�^Inc��D{��$�M*g�.�!��!`bᣠ��y�ʏ'ut
 K�<C��Т�MT�y"Ä2���Q�+�<<�th�ţ+�y��B�����Q���)�H�#�`��|I����c��:�(���	��f�u�ȓtan��������IÌ����ȓ{k�$Ƣ�?z��,<�H��<Q���銡k�����0^c*-�ʐ�%!��5 �Ib/-�,�W	B�,m!�:I����1��2+b��J˦ <!��Z�<+h� �F�r�l��ˉZ~!�$��<i�	�D��=���Kwe��{G!�M?*��Kda[�vE�s��x$!��=yHeX���ny�A�Uq4��D{ʟ�(	��C4 �T(��~�h��"Of��Iڨ[����BE����q�"Od)xFaW��<����
*]\� "O"���M��,������B!BH�Z"O� ��qa�Ȗ=�@�+�=n+�,["O��8��)Yzi���6w$��!a"Ov� �>w�hз��B�%k�"O�qRb����27�F#u���$"O�D�A�sz���_�`�,tj�"O~ 0&��bK��4+�Sc$�c3"O�l*G�F-i1�� � ��B"O��Um!X�5�̎>� 8`"O怱�+	z�X��QD�紹I�"O4HU�՜�����!N88A"O<�#G�N'J�Hf�N�
1�3"O�8���LA�9XtGqe���A"O*��hG9~2���&�)o�@Q�"O�Â�4Ϟ� P�9�2�Ȓ"Oz���\�rz�����X�*]@b"O��fL�:ufFu�0F�tnr�:�"OxH� ��8<�p�3r��g&H 0"O������9��$�EE �)K`�i�"O����L1ˢjԍ_:@��V"O���+`Iz,��X�J��F"OlI�#ĕ5�`X7��r���2"O�d��%H��频$�%.�5�#"O���b�n <ѳ0����i�"O�H�_�%��]aA@5�R�a5"O4XY�ݷt2��3���'q�(8+W"Ot *��e�$��ekA�Z�J ��"O�@�C%�1��8��Jʋ	g�(Q�"OpQ���sv��2
��\�8�e"O�ba��T��)�=:�٨"O�P �� �Pk次u���価��"O0��ЫF�Ls�	���UdҬb�"O�xX��2/f��t�_�tY�`#t"O��+a�ԞR��@��L�Yv�D"O4��Vyv ��iK!X���;�"Oʉ��Ӕ���"��X����"O�l�@ԋGO��s摒I�~�p"O��C�Mq�x��eX�Y����e"O��J��";|�|`�D�8C���x�"Oܡ[R��%&*���D�+V�<�#G"O�Ӗ�B�uZ< ���N��"O>��$G#G��5A0Fa�*,;`"O��p�ʧ.�~�5��C����1"O���%�'�<ITQ�:��%[C"O�1q�F��%�I8	��l��"O��b�ےe��l�'��'3����A"O��q%��	C@�iP蕣YИ%ٵ"O�i`��r�F\�FN�(�<h�2"O|`+�'O�'8T�e�Ń%�TdJ�"O�qP��0E��R�g�Հw"O������:��H��A����"O"���.@
\cr%3�^��!�s"OrlJL�Pa����/H�#"O�� D�*(�Tr��G2��c�"O2�+��?�d��t&��OwHQ�"O�(��I9OH���2Sg�x��"O�D⴦���j�IA+=`Z<R"O<�s�a�@��G@Y@(�`�"O����D��栍�w-lm"S"OTe�&�ׂkJ���O]	_3B�#6"O.�HT#̀Zq@H�VnAN����"OF��)�4�pU���7?Nd�%"Oj���nJ��L�`L����"O��Yf[J�h��7m׆uc2��P"Oٚ��&&����k;g[�x#�"O� Ę��jµ�Ed�<?[J�C�"O`�D��vu+#�wc���"OX�*@Ɔ�V:���͍+WN���"On1`&ץc�,�ꒄ�H"�)P"O�1a	/Ny�p�fiQ9���`"O>�c��Ǟ%0pH�7�
�@̼͒�"OLA��e�lMXbc
3`�l5�"O�����R������)��U��"O��J�N�0D���� P�y��%K!"O��/��0�0� �֣z�2�y#"O4Y�)W�#���!�&m�� �"OL82���|�(��jZ9=�x��"O���:2�d�wcϸ]�,A�"Ob�!�cW
c��P��l��k���"O��p"�U�**�4h�:�"ON��c��o7��)5��O�ĺ&"O��
���<����&�iNHd2"O����qG�P��&f@�	y"Ou��m��X�g�*3N}�"O�ȡc�1���Sd� �$pcw"O�	[�K(׼��uBл�F���"O�Avo��K��I[�'�,nW��2'"O�CV�;)U�0��U<!ې	��"O�Mw��	@ ]Q�@��
n����"OL�3��Dm�R�`g��$Z�Y�6"O�h�"ݴ"�ܹ�G%��":��x�"O�jD*Ʈ �U�T�IL|��*7"O�t��eA1u��ء��%lv����"O,�0��"&�� x4�Fv�f���"O,@�7�x�C�c�PU"�"O ���: j@d �(HP"O�<*��Ԡ5��(���/3�ə"O���C	�#]�h��7��%!A�P�G"Or������cn�1(�/S�Ai�"OB���ԯ:������M�<B~i�1"Or�Z�cV��1�%�|��Y�$"O l1'��:3LI�
���ТH7D����������Q�@r^��F6D��#�H�$`��p�`�<TI��!D����k�#hܝ�Ώ�3�`÷g*D�\!���s�P<ڥ	ьKk���j(D���F�I��*Y(1�1���oB�	*P�hr&�1�zy�O�+7�B��:J�f I��ԯL�p��mķW2�B�	Rh�2�.��&�V�5�*f�B�I;~ 8G�E:�x�l�:�B�	lxI�֍�Z.���`!�/ԬB��估���LZΈ�+�=�lB��:���m7���B
E�R��B䉭R	ga�<,���ejêx[�B�	�D��h� ASh7�\i��6��B�ɵ�.���� 弥#�B�9s�NC�ɂcؠm���
�
�̝S�$��
��C��n���I�/�/!}���%��!M��B�	,��=r�F���  ��N�PB��*r��	���5e����߄)�LB�I*u�\�k�/L$[&���.�,�BB�I�HU����Yvq�q[+R�B�� ~!�R+�}H93����5"OZ��eh��;�7�:kP�	a"Oj�2�b�70���i��^O��'"OL8b��3K:��
Z)c:H�	V"O� ����&%'��p$,N�!"`pK�"O4��a�K�>�b�K7��!}"���"O� �5R�+7|Ց7Ȍ1� �C"O���"ω(��R���/R��"O`h�oS���q���7�Z�"O�}CBH�n�q:� ̒Y�"O��#Q
��������.�P�R�"O�`��0JH� �f��oΚ=2W"O��$l�'*BujPIWm�h;"O���עZ?"�����,Sq��"O����dJ!8�!1A�ZUh��E"O�����7 �f!�Ě,Z�陦"O����(d�X�{�_�NldQG"ONL�2/ZP�x�A-BY:�x"O��1ad)����U=F�I�`"O��r�g^��J��s�̊+,�=�2"Ol��T�*'�Ѕ�ç���V�{"O��2㙗T2�(b�+A�	�"ORj�
�(��0&�-3*Х"O��6�յc�&=@p�H�!�m�"O�iY��iN���"Vu��]�"O-�T��23sLA���f� ���"O,��b��d�QC�[����"O��#��˦-."9�A"�3Rݸ$"OJ�@W�ə� ���-�S"OBy�a��x@��)/�f�XTp�"OtL�B�' �
���'м�)�"OL(�+�!7��|�s��Z%XC�"O�!@f��V� 7�U+^�Ĉc"O�4sg��?���ra�?��"O��{r�ҕ	#�9��o���� J�!�N��1��mֶz{���0��!���#��a�%ΜgruJ�̈́P�!�F�&;��P�d�d2,M#�D=�!��W'N���d&O�5��9�����!�Df�lQ�����*�N����ST!�ڜu&�P����q4����F��!�$�>r2]�6d�|�3'��!���x5H�@��g!�`�CB�
�!�DC6e���yr������V��
�!�d�!!P8�pVd��V� �k�n�?-�!�ǂdv��3��6?D�)Bv/U>O(!�$E s�m�k\�/�������=/!�J,���A�O�C��)HC�M�T!�3B?��+�Ĳ-{��� 
�!��P����d%ƚH�����ЋkL!�d��
���3eG�1U�L�Gn�W3!���t��֡	�d��QBO!�0ì8B��8>:N�S!��S�!��	�l�u3���X4eQ�a�9�!�-RӜ�0S�'DT�� \��!��$p�&�s�`��PdH�ϙ�`�!�ā�wiR�zP������H�!�d���Mс!�d+i���2#�!�Ǎ���9��\.f.�p{���x�!��TK@*�77!:�H M��!�)_ ��pc�(K�&� ��#v!�䗆jےA�㝳��b @4d!���Uqۂ(�-u��Ư؂`!��
�\:D��R $d���f�0+N!�d6 ��0��NH6E
\K��@@!��LT�Rd�cƖ)T�8Y�q��!�B:R�"�à��Y�`D�.MW�!��]�[}J�v(��bK<�k�-܍�!��U?dvT�pf^�=� 10�K�k�!���*�2�(%\�rc�eď�$D�!�� $�R�	�d6�qc���+R�>���"O �w���,���Fv_��xs"OA��-(���h "�
@Z��K�"OH FǔP!*���k\�7Tzp�p"O6d��gǰ ���!�)|:�lѷ"O�ŹW�	�\],�ا`)(��"OZ��N����s�;�"O,��@���w�^|��̰2����"O|�㧄������Ⱥg(����"OT���ު P�� �J���5"Oh����8F[9�ϊ?6��Dɇ"O. ������a�׵$�*4U"O�:@*��I_8u�wAw�^���"O^��&��:�Z� V��"�P�1�"O�$��B~����I��9i "Ov�XU	�9G��{Ư�r@�S"O(ś�j�3h=TX{[-d����"O� ��&D�Hv�p� �.]��zc"O,��e�<������YD���"O�`8��C0\��0"�B��8R"O�}c�dΝZ�|]I� S
B�2=�#"O0P�NSN�ړMN�5���"Oƍ%���(��T�܁\����"O Ec�jP�P���M��2���B5"Oh���%Zv�h��-��t��"O|Ђ�Ɋ�U%�a��Ҩ�"%"Op`��I�y�&���R.h����7"O�x�"L�%j��X�D�@3pQ��"O��w��	��){��5#艳b"Ox�S�g�A����m�,|��zP"OY�.T(5N�Y�+j�tAT"Of�
d� >v����i�9K 䋴"O$U�Q(V:0��o��l"�i"O�A���K4)v x��n�ad|Aq�"O���`Ej6Mm4/T���"O�-�3̃�gŶ�5L�R�6���"O��Q�*Ez�d*�)�_o�dТ"O�y��¿��q�dI\�@y��"O(����Egl-	f�41g��$"O�,׋����yh"f9��A"O(� �ӥFF�K�-ؠp/p1A�"O�qS�aZ�p�����=:���"Oڰ:���f��3�\<p�//D�8i�T�G���"��<&�r/D�P������m!��:D�:��W�-D�d�v&�I�:T1'^��,�z��(D��@`*�����n�8 sK2D����Êhێ��P�Y�.�0���1�O�����~�!� 5{��ȓ��il`93.�1�y���0�d��kE h�2��s�_��(O>�=�O��c�
�1{L��餍L�+1�Q�'$ў"}2�
���e���Щ1�M)b�__y��Wg��(���K�+2h����]p�H��"O��q�
ކ1#L]�`�Qf$G�Dt���	�L�}�u%S�$o���H[+˭C䉒\�vتת�-wh@����+�n&[a��R�d�����N!��8pe�W2��<���Oڹ*�K��z�M�' �U�@N�s�,I���*��~���OѤH�+Gh��	�Іp��҉{2�|��g�(#E�( ���ajX�
ȤO���Ȱ$�yR(]F��I'!�8+eb���K���$:�S�����2�A�#��q�d�J*\�Q"O��#�G �KԖ�P�n�s�j�Î*4�<����Q�4����[�#u�����=D�� A�i޹y̮�(�*V�ʐW"O�8�h�+n�����K�_].��b"O��bLJ�(D�h
�o*|�B`�"O*����T9c���A��-he��"O� -4������!�5j-qL!�D�Oܫ��P>n��Q�D�	���R5�i7��C� ���#�B;Sx��ȁ7K!�)	8��v(�y�2����D�x�!�DάJi�,����\�L���e�0��f�)����L��ؕ`��g���*.D� Q��c�X�s��N�H�`l��#+D�Ѐ�3!]L�#+�2&�mZ�.4D���V&�:E��4�uZ3�LJ�4D����$�&膐97���l��B�1D��x!c�3~$F�F�U�6眽{��k�"�=E�ܴ1����Ҧ�'32ܘ��U�;�L��'���!�)§�4i�b�4R��ՠ��M!<"��'("��$��R��)�� ��i0�y�D��d�!���Mj��A���
bfה`a2�OH�`�D�+KQ�e�1�+F���$�����@��ȇvҨ�����'<�x��"O$P;aj�*
�hUj�ӈ��I�C"O�PJ�̌��,�&+:u<E3�R�hF{���'m�h�bk��{���g"B�+e���M�|U�@`D��l�ů�%r���)c����>��I�w޼P����<��'�r�Т��n�
5��A5�V0�'���R �-W -p��}Lb�x�}"�OV|��)74/�(�b�.)ꔩ��ۧ�!�$�a.Y#Fϋ��u�!/ �V���&ړ�HO���a!�����G�aK�"O���T-O�FY���ZY~��\��E{��)Z�.�dՐ��$K�M1#��a|R3O�� �#
 BD���m��S����>דH@I�`kD�AT���H��kb>`�ȓ[� mP!��'P��%� Q8=0<��ȓ{,����=�eK��܍?��ȓ"s�5���F��KÍ2P�� ��Q�Fi��刞�<t��Z�70�ȓJ���q�FܴR�3r(X,k�j�ȓ"^��s��^�CD��b@bɧb�"�'��(��'9XD�DH�Z=���(H߄������ߔ��D(BU����ĺ��'��d9<O�hjqEA15���#Ln=�'��	˦�l'��%�E��#¨`����Q}ج��\��9�GL��U����g��u����=!�'��'�����TA��@N���)���
��(�?D�(ك' F�h���*=f��* ʓ��<��K�9c�#��ڗ):�Wc Q�<�P'9O�x<���̻\�̙�w�]�!�K9Q��8�J�� �Li�Q�&I:a~�V���d	R9sp r�X������0D��G� 2�i� �ָ&bt�3n/D� ��Iއ	>L�3j��l�&9�d�-D��:5o�pv��xRU9z$�"E�)D��9W�5Y�N 0� Ի/��Ѱ,)D�X*���Rb��3n�0�f9D�L(eC��=� &^8l��Ԙ�7�O�ݖ'�͹��:��"m�0 �X�'Ӕ�t���k]
)��+�m���yB�s&�y2�	g�K�G��ȓ+jv|[g�-�Q!G�
�y��#��|��Gѳ3����X�}ڙ�ȓ".�9�ゎSRr1C�ƶyR�ȅ�S�? (AH��RϘH���һ*���"ODY�)c|���0m_
y���Ce�*\O�d��Φ�T��-J�v�($���x��)擭Y�� !Ćm�����.S�|�m�'L�|:Oה6�� x!+�!qrH��yk2�I|�'V(���oR�P�ua�:|~�<8	�'@���n�_f�� �älf�8x	�'��G�F�X���b
;	�'t���և^#L��1ժ)W~n�1�'ϴ M�#�`=�@�Lr�A��yKء>׀�����& V� $���y�B�"x ���O��nB6U�c���O��G�4oܖ`hА�]�b#D�g�y�,�%"3�(���2X
�80���"��D�I��H�� X����'��w��}�e��"O6 [�FZ85�Dcd���`�"OF!P�Nږ��rb+�Y͎P	��	Y�����S���ʞ��Q�%A3w�!�O�0�X��a���1�NU;��]q��hO�xHq��:g��[E��`�А�"O�� ��fʨ��e£MM�Uj��$/\OpMHp�&�6G��К8�@
O�7Mˤj&�ihR˄�n[l����v�!�����ZD�rSώ%�!�d��I�̲�G,\��q���Y��!�C*'�0MjA��t&^`R$[�V�!��T�q��`��>7����R�!��!"&���c�
3-
�!�!�d�|b���Fɨ'
h\��رR�!��Є�$xw΀1_ �!I#(��u�!�$ȻX*��v��"� |�D-׌�!�$ZgI"�2!�ĕ�*��3쓐ul!��96@���ͨ~�9��}!���	#�8�JQ(ȟs
�( P>hR!�B j-Z��ÈC�]V(m	炅�73!��g� �1��""�]rda]�}�!��E��~���i�%|�D�Woȗ\k!�+6Pt��UEF�q![�9	!�Ց���I�)""e�P/�"=�!��O��l}���TQ"A���;�!��U&/D\rA��)ir�J�m�*!��	
���L�3ߢ�⢍@=o�!�G�E�lE���(��s-m�!�D�\$%0�L6p��Փ��#�Pyb �	]���`�ƙEt$q�MH��y��!/�D�a��G�����E�y2N�)���YӭΦC��w��$�yr�ױO%:$��L7cV�B��yB� iU�5�MB;> ��I���y��L�g��[�c>.캔�PB2�y�%P5��lҷ`�y�z� �э�y�)��cm�@p��X� ^���<�yRm޳B�@z���w	vه���y��Գ��y�( 	oL\��݆�yR X�csع9u|����#��y�`���qm����$c���yb��:?u��SaK�2�>l#��F�ybbK�@��Q�vB�	x�.u	����y��i��RcA�x��S1Q9�y�Mf{.$�U��D���%�λ�y��M)X|pyc�7;tp  �$ 2�y�HQ.�ڠ1� �|�d�T�:�y҆�1F��Ԃ�'�.]�Q�S퀿�y���RL���'6��Xb����y
� H%딇G�v/�iP�o�#~��%��"O�ಏ�)�$���,	Z�F"O�B�ဆS�0� �ًG��m��"O�xZ�"}�l����f�^Aj�"O��1�.�Sfb@I�A�[4N���"O��+���W�Ha��"�~p:#"O	 T��QpR�
��Ȥ�6��t"O�؂�.�����JZN�T���"O��` .�#s� ��W�����"O���˕�@�0:��%H����!"O�g���x�,�� &G�p��1�"O���*�:d���Ǫoknd�"O��٤hӹ!�;G���<?@�2�"O�I�2N
ܖ\�v�R�/<j�`F"O��xb)�-��-�m��O�&��"O�Ac� 
� �ؖ�Gzl���"O�����3�6�q�18��@��"O�m�G{�`L�ĕ	�1��"O4�ѥ���
�i c̓	��!�"O�*�̀>Nq�S&�?+�ɈF"O|�1!�Z�y�j��V�#f�C�"OP��B��&E.�zժɽ,�u�"OvM�ϐ�R%��b�f�1����"O0Q��"ޔ�hd�R���f�	�"O�]��Ȯ-�Hp`����Ri�w"O�$��+�Z-�2�Xs�q`�"O~U��JZV�D�@�
h���"O�E�r	I'fs�X�0�4}�|5�"O�A�j���Dq���-HiF�*�"O+� ���, �c�8ǐ)Jg"O>�c0 �Y0,y%�� �PUC"OЇo��f����
;��5xw"O�(�CM�	�4�f�N�Z��V"O�1$,�,Sq��j���2sD��"O��Ԭ\5l���f��0y��#�"O�e�o��:e��)E�]*tuX��6"O�4����=HRH5K����xv"Ov�7韌j�<PZ� ��	�!"O����KO�^�����
�L��D�"O���(�`��I���4{�<��"O�Y��#ͭ%�4H�v�'p���p"Ob�0M�3$W������`d0��q"O��R�&P�sl�֊�iH*�W"O���⬀�E�V��
��5H1"�"O�d��/�=[��j���s��q:"O6h)SLX���1gA� �vU��"Ob�����Z����u�fC�l�"O�����
,|xC�Ύ9��g"O��1��lɈ����Y�D��"O����9#2�Ly�(σB]x�C`"O:��tI�Od��Q���D�2`�"O��B按��V�C�$D0+���U"O�p	���|��	r�Wx:(�"O�P�v�S,�x��gi����m�"O�8fE��!���@$Q���"�"O ��-����Qw��+lz�i�"O��!��o[^�r(R�wd�;�"O���G�xnpB�.y/�A�"O���e�<��e�(�S�x��"O��7�O�<,K���jx�K�"O�P)Pe��y4f	���EsD�"O���՗O� �ؓN�Iv�Z�"O�9C�%��#��q�,J� �. ��"O�YB�K��a(�1$�ٴm�|<�"O� }"�R?]ނ<�iʨg��=�"O�l���(i ���ݯF���j�"O��{Ā
1&e���ç΀	�p�"O�)�D�e��hpt��)��g"Ot�$	 �a@�Ꮦ)�U*P"O��`ʞn��]3� �4I��˒"O6Q���V���1�5><����'+4e��,�t�؁��β�]j�'�앀�N@�7�ƹ0�nF8wn<@�'	�D��`ƌ33eƋ��,l����'��a�S�'s�$����"O�,��'�x�A/G$�,�ECThlh��f�)��<Q����d,�$3��	y�,!�q@�m�IS���O����kT<x�QҲ�Z<X̄�	�'� :7 L�J����g�$����'���!m� R��%��N�PA
�'�h)�qb��+eza��]�63�U�	�'��`�\�HU��~D��0	�'m��s �89L�97��6v���'�p	�-ʢi�4@i�dѽC����';�Y"3�_���Ƒ�:�*�0�'�<`S�N&ʬ	�W�+@l ��'��HF��G��ٙ�,�=)�*�"�'�8�U2A	���#�M9'`��;�'+�Ⱥ6`[�i"
|����2t�
�'�&�a�nѵt!ãV s,�S�'<6-���"�PXT�T�j0|���'r���6��g�Ty���ɗen: ��'>�@��䆬��C�Č�c��X�
�'<�@���p��8��[Z�T�*
�'�x-	�K�&��H���G�F�
�'�]��mR+*�l�AD��Ah�4p�'.��T�(y���[ѨS�=�Ʉʓq�I���:���F��(Y\ȅ�w��4Q��
+�����`��tԇȓ<l�t��ʚk�朊��R54d(e�ȓl���Y���$���K�ЉR�D��ȓN�v����W�� ��܁AD~I��t���IT�B�?�Е��H��[|�t��}�ث&�@�F	�E�
,�|�ȓ��9�,�1�P�I�lP
D+vx��7��� ��ȡ,�RQQBṅu^M��Y�QАF�#s�]Q�"]�V����}YБ����#O}b@	O]��=���Z���K����
Gj1����(*�)tkR�mЉ���ǉc�d`��Cf��#@NZn�*9�D+/�NT��Yc�9�Va�ju�����+�ꐆȓ|�X��ECW�OtM��ʦW�$m��3�&�0��qm�̉�B��72Ȇ�Ȑ�ju��
U@9v�]�#n��ȓO+Ԃ`�Y��8��@lJ��8��Na�l
Q�O B0�<)�k»+7`XER��N��0�1�G�w�`���-ZX8C�	���<Wɗ�h��@B��(C�	�%�`��P��7����G0c�
C�I7��#%Ê�;�H��Ɖ�f&C�	�'Mn�C�IQ���"!�4N��B�	�.�$*�LN���̀�DN�VA�B�I>k�X���ۼZV<1���
�AF\B�3;@��� fiE	�&��.B��JI�w!�	53�Jw"�� �B�I�p��t��c.�����"B�I-���J�bD�<}4�zp��)d{B�)� 0�c�ł$O@��&��#��D�V"O�4*sCU<`6�P1e��{��8ِ"OD9iФ��HLP� ���[���*�"O���)U�J&<�┄H��"Oh��=�z!F�G�w�t"OR-PA�����r0T�h�r!RB"O�Igc��8D�;rM��(��"O��:��&T��bB�NPR�"O�����M!p����5#0���s"O@ŻeE��i�x��#��w �8���J�OH�+QkVbYX}#�@������'O̠&��o�Bkw�	h   �'�0�0Cd��aFdM!7I͖{D����'4ĵ¶i�`�����9{����'� 9����!������(��=8�'8�5��R�1��(z�gN (�h�	�'���7D�x�( �-�8�`p	�'8�ȔA]LtrK�����	�'�F��O��{"�üx�4�:
�'�q��ܪp�t�wsݨyY�'aRi�)]+�<���c>���'NEI�#qV(��Ρ^:�e�'�"�C6�(z�d����� X����'����HO;\�2�R5��Wy i��'���T@�>�z���K8LV����'� ���'}� ����K[�8 �'�8�7"�>4~t���XIk9��'���ڠ/˶o���+!J�A�Fe��'�&}����,��Kp�B:pt��'�n��O�?J�V�`Lߑ4�^�:�'����ďlE�T!ǩ%Cj��'����ס܍d�u��b�"ƔH	�'7��K!`�}*�a(�BP�EZ1�'&X�kB5m���+���
�����'z.�*�k������E/����'>j�cf��hj��4�38�l��'��0Ë	�F |Qh��]��ց��'Mꨱ�e�(	�asS�Z�PI�
�'R�ps̟2V�
6�	|
��
�'ɂ�q$ߖZ�n��RIH{� ��'��D�	�*�B� ҥQ�|��H��'��ꆊȸ_��Q([>u�R��'&8�PB@�i�D�#�Ӌ#���
�'JZ�XA����1b�<q���
�'���i��J�a>&aI�d��r	�'�P�C���Y�J�K&�˥ݎ���'LX��,�p���RE��-'��A��'B���0Y� ���_�"��I��'��\넭;X����M�+r
Lxq�'�����o&0/lQ��AT�m�\	��'��,:P�SF�.tb0�P0�@0	�'0N�� ֹa
�-����!#�T|	�'TR�s0��9��� �	�����'0RU�G'_�=Ą	 �f�<u����'���"I\&%�$����}�8��'��h���t3��I$���t���I�'�(�wL�(8��A��G�  g�D��'�d�Y7�֐m�-Bv�Rz��y�'[���1�:-�
Y��.�	T�a�	�'���ӯF3D��ڷ���e�	�'Sȡ:
�r؉!"�*�0	�'�u�ʑ�YP����R���'�EoǮK���ܓ0��1i�'�H\ӵ�x��<�A�ل#a��p��� ��aM;eiZi8q�ގ�`г�"O��G�Z�S��YS��\�q�R�0"O֜S%D��i�L}��R'6����"O��*�*�$�[�I�"�:�6"O�a�փ�<l`Hj��F�i���"O
�S���N
�h��!�=k�����"O����};��d���~��"O�27����,	e�X��MU*Of���EЕ<n��¨��`�Mj�'�,�!�+e���`�S?�l��'���A�A�:?,��m�
�*ት"O��j�Mֆ��8E����q��I)a�zQ !�YT�����P� u���P?*�����Mv�n=��*��F!���L)e�2��/B��a��M�ne!�	�=��}��)˹��e��Ƀ9Rb!򄖑�Z��Ǒ�ɘ���ڗ5<!�DX5e�Լ�4���G�p��ɗ�!��u�
\r3@5W�j��BR�N	!��"p�)��n��Z��#���'W�!򄔨w�Ժ��O�:�iqoO�ur!�$��3��ZrJ��%��t8�H�
�'ݞlr���M�Y����Z,, �
�'�.騣�O?��2W��J�f0x
�'J�OZ#DbxaZ@�<9���1�'b�, ��յ�l�y����l�bpC�'�l1��=���`��)fV�x	�'>�@&���duه��1Q0)H	�'1:@�wH���bQ��τL}����'�*�9�?B����T/]?��0Q
�'Nl`C�S}Z�8Dg�gh29�	�'��͡t��h�:�Y�N\ :�z�'�Ĥ�$�������\M�pC�'� r#B$@��"��+#�
��'������E�m��	�bk;P�c�'��P`cb��P��2r�� �ղ�'j���&�1��a�9x:���'s���f+G6p���1�L����'��%�3bQ�$J��HT�A�y|�Y	�'���X1☤}Az<���F�w8\���'lV��n����z�@��]��Q�'@<4�a
X�P�.c����D�+�'L�	�E�jZ2�S�kݶ
��`�
�'�4���d�<XB� TaS��Ha
�'=�q1��V-0x�i�!0T��	�'���
���>SÔ�!p�ՙ� Ի�'�Z�FR��}���O�a��'n��"0	�e�XM�w`ө~�z�A
�'����bƌ6^���J�"զy�:��	�'�ly��]<g�Rp��,\����'��)�bɟe����ˉ�}���'�Ar�)�*O#\	a�Aq���k�'Ԝ��`G�<!t$����gF�{
�'�ĩJ��T!K( �!j�2o;Rd��'<,]0Ua�"r�&�Zi/�����'��ثC�N#=�"8rA�C&u͞���'?�i`�aԻw�Ҡ�q��3���
�'�T���
Vmz)R��B�؉
�'���0�bL�"��J"�>y�ꤺ�'�V�X��n)2��
���5�T�<�6$�.`��)#TJ��=ʕ P�<���Qx�x&F�.�}���L�<a@�+Ln4�b�+X�BJ���CD�<鲈J�L���L�� K���G�<)��X����Q��=���E�Ct�<� �5��c�v�D�HW�`�tI�"O��tHV�Z.�0�b��w/~x��"O��v�6$�8H'#J��@�$"O�8��[)AO"`�tN.6��1�"O��	V��$$��S��5=r�V"Ob����̸ u��2� L<�@"OH4�rlѪ)P���)D�,2��"O����!m^�7g\�6Ԣ ��"O64Sdϻ"�`1�Ǯ�8� �"O�O%���IF)_��9��"OfD��E
'g���"�
��D"O��E��5� Aq�Oǵj�h�I7"O�H+��s�dU ��%��<��"O���ef�fl���ԚPlx�5"O�Ԙ��71�E��B��nA�1"O*�JS���MOd$�r�/Hh:	c�"ObŠ ��#�&���J`f���!"O܈#4�U+5"�Y�
��)�4���"O���W��V�`�k�7�Θ�"O�q�d���k�!���#6�n�3�"Oz���.Ja��*V:+��93�"Ol�p�f�(9�@\�#�o���e"O���ǝ��r���@�I�h�8�"Ol8�� &}�T�F�^�G��UX�"O�,kt�"���#��<�(E3�"O� �	�r��Ԋ���$yZ��"Oؼj6��&��SS	�?��!��"Of!�\�%K4E)��7�^ye"OH�v��9�Ѐ��aJ:n��F"O���b�<殅	�@�>�Nt��"O�T
�π=d������#��90t"OD�:�.�#2TL2�a��v�(Us�"OT�)5�<R6�*��B�`��|��"O���&N�ܱE	��F}�0h"O6��w���yQ'��l��pA�"O�|K��=�2�:�.e�j�A'"O��e�a"$Q+g�M�"�'"OTju��jZJB�̋?P���Pu"O�|�Ơ?V�~��+�'_���y"On1�h�Lv`�"%�+h4ɣ�"O�}���oX�]�ŽS��+c"O
����S;V��i�B�ʉ�cG"O.��ĊK�� ֔ �����"O���%�ǯ3xn�[𥖧��I�"O��b� �%G��s�R�܉0$"Op�:ծ^OѮU8R��t����"Oxy��%�*m�D4Za�F%>y�h��"O�H!CR�y�Q�C�D3}^�� "O<��"�G6�=�r�_�l��م"O&ԩ�ŝ2=��t�$��#�BI�uO�ܻ5 �6*�ʘ( � ����hN=ېxB�I����!�قp����$˰<�2��'%J���1�6I�W&���
���'�qC��nH��І���ˬOjpS�-��@��l$�"}"sE�.��M{a2}C���$�\�<i���fHKqȀ�8�l����S~���\x���8�0<Ip��lr,5��E`�;i�Kx��+'��
rN�F��$t�Y �eE�cv�t{§ɋf��`��w:J5��@J?)4h�b��;�ʸFzB�U;��X`P�މ�M%?��j�**h q�f�(�P����'D����ԽK��D˗�*-�Y �y�Ĝ�	� Q�x��0%���~���i�|�z���-.����C�tRD��'U"@WFT�Ꝛ�d .��q�OF]�M�+=˔�	�������d+r`A����W|�fA�4B�|b&�2�. ���@H�? ��EI�.�ĉ��R*|R$P"]�����37d�Y��J')��P��Ä5o�<IÆ@23n�m����%-��@I|j���::^�E��h��a�����h�A�<!���X|�m�U��mf �q��b9(t�E�5^*`!��f@�5���'`ܤ�� � kp��h��l x�'��*�S�N�&�hV�R�ت���O4��$lCcX4  �������T�qZ`j�P�`$�dϑJ��|���<D:�k��N?�ᄪ�4+>A����9j�͠t��O�a�j�l���E0yv���G�*Q�H���J�@y;`��2}r�$>e����;SXPX��M)*�n\at�%D�|�2X�P���0wf���d0��vӂ+uJ�?��̋��Y���F��46:�m0E�4Z|Jm��]���ȓK�Y���7)Qj�����QJ��t �Ŧ��
�\���Aj����-�6��Պ�-q�Z�h�Kړ�h��dZ�b��HB�j��1I�'2e �cX�6oTd� h�������}��;Ԟ���Ӧ�=�T�=Y�_�%ĜhXG'@}��11R>!#��	
H`�å��J~�<[Q�5D��CBc�!l�.�k��E�z& �OT�V	��#Ң� �	�d&�G��
 "V	��脿^�9S�&��z�!�$$S�Zš� ��thz���O�Ntr]5�
dz��ֈX��ع�W>�<	��S�o���[�e\G�(��p�Gx��� ��G&�9QIO
(�Ь�U`�9?�
M���������]a}�<v;�}xb,�q������hO��Aa���l�$#�/�2g�H���Z-z0E7���b��}��q3B"Ohy{������y#耮09���A�'�=Y�lQ�1��R3^��n}G��a����i���*�r�r�bНX�!�d)"4F����Y�z�W3')��
#Ԛ8|(���9,h+R>�<9�"E� 1{��r��¤��lx����`�'!F���.>�l����AW����Q�L�E4��ClF�)a}��ȯfOTa���5`|xY�j��hOZ!9�kQz�G���Z���O����B��.E���ŪW�bל�0L>��4�p=)��67��{��#gfԊB���<yCi��$�Q{��,*0�e#��I{���6k��is����2\�����y"��9fE��� ���S&5F||�Rf���y2BL�eH�"=�^9��O�d$�<�;(��d��BB%=M���V�״t(Pm��I
UX��á�K/x:���� D��h���E@0x��"'#;��(�d�O>���I�31t��#B�P[�����[�'K���*N� MDi%>���� �p��c8��$��C�<1��M���'>BS ʨ[Ǻ=��BR;T�d���O�qsD�$v�1O�O�
hظ(ǅ�0#��B�9��p��M'6�"���	�Ģ?ً�iE=w0*E�aHɅ/<�M���?j}!�$�(!%2`9�I�= ƌ Z��K�Lg!�D�V�¹`Ĉ���PC���#[6!�$�12`��Vkԃ�R����
 N!�$\�\"�H�B�Gx6���숄`�!��){�t�ש��)|L��i�!�dï|��x��њbҙy6�΁8�!��˒oᲕ�1�EK�,SBZ1�!�dU�{3�V�S�y;Zl3$Y�!�$��-�r��  �k�R�k#���!�dp%Jy�J�4�p��s�),�!�$ŏV2� �T�B3y��,K#���!�$ٯ�z����Gsb�A�Y*r�!�W~�q��B�2LMv��@�Y�'���d�?6e�5�4��8J8
%c�ϡ�y� 
|��57Œ�A��N�;(!�X�oAҨ����"rz�ŉ��28L!�Y
o��U����/�\��QÓ�|6!��g4�����S=E���1`LW�1r!���>N����} h�V�!
�!��ȼ#��@(�a	�hh��2�Y;!�!�F2��yB�B���A聙�!���#Pt�x�Mļi�R�J�͘�"�!�� �D�3�Y̄2��C>B����"O̍�4��a��=��v�P��c"O|�&�Q!uc��1BX"y���3`"O�a�g�6��5@/R�`|
!"O�;׭�� 3V@�ʏwC0DbD"O�t���Ky��S�.�1x7l�Z"Ol!��ש $�i`��^.�E8"Ol����xÇ
��n����X��y"�ʔ0伲���\VRш����y��A�N�Zਦ'�Wpz�P�>�y"�+z02�2��۞HF(�[����y�(D>*P��j���[X(!�'��y"-	�	��da2nF�')0ݚg%R��y2�
}aB<�+�k�F��7M��yb��'��aq��5`��	 ր��yb��)3��˴�S�MJL�u���y�IG2#��Q.�9^� %��[��y� E�k%����O
�	*m�PD��y�A�'[nTـ"P�9�pјw F:�yB%[�4�Ι"`�R�4���g��/�y��Փt[����#7�N9�ǭW��y2�F�Q$��C@�L�V�h���I��yr��-M���'�=V5��b�b+�y���(a�"psw��N �hp�hѐ�y�Ȏ� �3���!tr�Q��:�yB�݈w�f����l�U@����y"�R���8��W�Y�>TJ�D�*�y�C,7 ��ч��2b�
��5����yB'Q8}�W*D<_^Q�% ҹ�yrK�$�r�&#VDE`��D���y�P�=��}�%��0h�H��h��yr��2#�Z�+��+.μ�C���yB�P�a K���H_��W�+�yo�4� �B܌KlX���y�a�uP����ǔ8o�uQ�Iſ�y�+�wa�H���n�& 8��+�yB���D�1��X'ʸQ�E�%�y2J�D�:��^�N|>58��G;�yRh��%7�Xb�.�:���q�+I?�yB�Y�.=ތ#%�о���0��y@C��L�B#! gİBl��y�N�WŴLk@N�x5��[����y"���ZY�y0`�Ӂ);��X��^�y��>^�Hkg��:)\�®��y2)��h� �aĩڇ=�
rrI�*�yRˈ�Jn �᢭��ec������y�b>��J�'ީ[��Gა�yr�C�5,�����d�nm��gϠ�yb��%l���ы��	z���y��7#�F� �ɧ^������y�B�\/@I� _;t������^
�y��G��-�G,�5\���ؘ�yr�����h���Mr�ҥgޙ�y��W�?��pb��1ת���+���y�@�DbD�Qm_�j1K @��y�"M�W �͵o��(r����y���qx���Bm_�o��[����y�D�7.ڠ"�mj�������yh��4���\o H Ǣ��yR`�D�֍���҂Z�.�����y�)��ł�rRȑ"J�r��N��yRN�>q���KS˙�bh[��D��y/�Lx��G	����������y�`B):V�1��O�%��aL���y
� �����Vwj䬹g��5~�ځ�1"O:$+��O�`86Dy��$K��`Y�"O��"��� @����G�te�;�"O̡��͢=]�dWe�'0T���"O��#M�)O�@����!$2I��"O8�"g�K9wG���pc�*k
:y�u"O�Y���x��E�5�V	��"O�|RDc�Nz�O���+s"O�-;��_�0�N�3�a�-s_D4�7"O���[+rтD��H8�`��"Oʡ���{�� av+' ��"O�q�0� �a�X�k���*��Q�"Oޕ��O�e�~)J
��
P5J3"O�s���7=�d�������a"On
q���E��A.V��=zP"O(��-ŉJ��97��.K�l��"Ol4�l[d�����U|�u"O����a���m9r��&2AJ�ZF"O���E`�')�<IB�DK
܊s"O�ܳ�nR�,�5(�T,s<�Y��"OZs#�%UCf�Q���*P�=Zw"O|M�&L�L2Q��@^�x�"O��s�e�C�.|��ύ>EW��C4"O̹�e��T1z8�V.K�L�@M��"O`��Ù�KFD�0�oO�6�
聅"O����g�S�,��p�QXg`_�y"CS �b�Ã	#YjP�V��yrbJ�|ݼ��պ{Zbe*wC��yN�4�����Ȇ-�T���
��y����	ނ��� p
I�#�S�y�%�U �!�4��$H��,�y��� VDd�$�>	�a�Q���y�҈~�^h{�c��&��LÉ�y�B\�z��р�d��(����G֮�y��sG��+�H�[�f�BU��y��Ā��4�v���\MPi��@8�y"#�0����
�S�h�*"A��y!�?5��e#U��z�lE�yR��#V��b���0B�-�) �yb`[�cش��a�ӈ>8<\R�`
�y�nZ�2v�U�IX<2~6DJ�.ċ�y���5"�x,���!��16Dڞ�y��E�G5��"�^�#��	�5���y�$ЅE������ h����EC�y2iĿcO^�2�s�6�2�+�y�MQ�0�0�+���������yҩ�k���k� ab�*�� ��y�� t�iK�^,VF��V@	'�y'ڐ;b�{��4���8f����yN���F�y3*�sԅ�2�E6�yR-I<($A��&hRx8�����yR 2X�J��ů^w��k�GS��y�搿s-`�%ㇾ/h)���Y��y+��f�Dq�	M �t��2�y"D�ώ�A���MVH�Rc�yBe@�<��� �NJM�B�U��y�*H�����G�x��/���y�䗿)��S�`5�� F�$�y��۪h~�#���]���Y��+�y��H!*���P$�A�^�x=� %&�y�`Y�,�EzE�5K�l���c��y���*�j1S�O4yS2J���yBB�rb���с@�,��q߲�y�*&"u
ǮF6:W�� ��ɵ�y
� t����".>�J����S�`���"O�pۄd[�U�:-�W%Ճ^�pC�"OBM:s	�	WPݫ�D�� �����"O2�i�D<��"��v�֜�"O��2Z9R�x}
�)Q�x�&��"O��J��V�y3lp��H> )`$�7"O���� '�ꑘ�hU�f2�L�"O�LxA��X�T��u��3>�"O�q�#B��A���(����j�d"Oj�8�'@�]	r�̓�"-��"OZ���,@�Xrx��+�P�ч"O@�	�#N�*@�y@dI4i��P��"O44R5)��b����"�o�ԉ�V"O��HRB��d��V�ʂ1�V��"O�P�b!,a�0�JD!�Kx�:$"O�I�"��;%W�J��1RQ�%"O6�QC�8}&`t@�F-&E��X�"O |��ݎ|���
�!;���"Oh�1�S=#�@�5��,�x*2"OBU���KY�(�@*P7W��x�"O��uh �9�e�k�s9nH�"O �#��33������Q�>ղ�"O����È���e)@���ᨖ"O��S� ��$zD���(���X���"Oh��A�+R<�#6���LplA�e"ON	kDI(g׮�B"��,-��"OE�a��R��=���8V��y�"O ��F�)Z����d'	@��1�"O>��',͏[�0` 00��"O@�pc�U>"�f� -�-�x��"OV� ��1�hpq�K\�䝹c"O@qjU,C�Z.������K�̜��"O�����"�D���JA�d�ā�R"O�9a1�@�9���&)�C�.	;�"O�Q@(��x�Fy������`��"O��Q㟕v�ҙ�W��-vԹX�"O��Q��U�fςPK��d"O�QJW�O8I�D�f���!��"O�Pz1iL�K/٘%��S��7"O��* ��
�􍨑
	�V��"O8�A��� /���D�T����y6"O��S`�>f�,�ǉ:$ڀQ&"O�I8��X2|O��ᴤ��[��Z�"O��ǦM�)!���7j:�J�"Or�0)�/?�V����6=�(ɣ"Onq�V�RY��+�Zfz��"ON��3��ݙӋ޲�֬��'�����$l�`�X�*�1Sv��',>�"��*8$Ʌ�V�J�N���'/�!���>D��D�4�Cx�'�J�(�� ���BD�A�8���i�'�j9wGޜv����s�7-�m��'8����P,X
��DFB9Sa6d�'R�Y�cd� Um"=z���21z5�	�'�Z�F�Ib�4�
#FJ/D�4��'����	@�X�<���!�!F����'CL�0�HX�u>ܙM�
&�'Ln�x͔Z�b��G��5m�y�'c�|z�͊�N��8VJ�#��I�'J�LJ�םW@> �PHɿ�H��'R�,릠�J|[ L�/v8k�'�T0kuE�\��p�V�+�1
�'� ��t�i���Q�JU_if|��'z���g��s�=r��0Fh����   ��!�8�� ��<e8��"O����N�������#^.U��*OvHK���S_��x�!��P�q�'>��r �UVt@؅H͕eQ��Y
�'Bl��I>n���2&"Q9H��1	�'*�986�U��r�c�,��R�ҁ �'��'-�U��p��Aʙ2~��
�'�����M�!:�	�#�Z�E�4�	�'	
��#�?HDd���!L��|r	�'���*����8��sm� :���'9���X�I
��Ycgʦ���	�'T=���۫"^4y��	�z��c	�'$�����c���S�^�vV�	�	�'���r�f�y[��bk�U[\ͨ	�'�b��U�q\�i*s`��W:
H�'BX�ڤ�m�@�2D��/J\a��'�d�� 8�$��H�v�d5��'h�ͨ�dR�s$�Y�2d��w%za�'��:AO]
1����aN��	�'Gz��7)�7o� ��ы�2X*V k��DV�{��@���Q���U��1AH�lƾ��� 
~�Ḵ$�����Q���ek
�R-V�K�AR,<��?�����9�x��3ꖔD�X�l���I$y�!QT��gD�L��C�#p����"j~<+����*A�N�ᆨ�%v�{q& L�6�щ:��O��$����!tC�d�����P��(A�|Hçgc,J�k��4�j=�C��h���>I5ڮ����'V��AqDň6�py���;5�'�����K�S�'tʐ��ƀ̀o5��d�:Q����'mx�a�铪Oc��ˤ�$^TT�VaZ!qk�7MLy���"RË޺�,x�Q��	"�l�PM�5��㟤�	�'EY"V���jAH��^�,Z��>��F���ħ,�=��,H�Db���!hy~�'�x��,;�ا�O-��z�䗎{�(���_	;��T�¢�찧��/����i��0|:b�lֈ�g���_��M�_ꦥ��Z1u�nz�K�=ia�Kç��q+3'�2�b�����	A]72r@Y(S� N��p짢��&$1��C��?S��;Ή�F'0mJ�O���B�i�,cd"3�LX
��I�m?�l�VJ��7H��r�1O��Γl�&�s��m}���ܙ��F���P�QN�	̷�a5�7�S����Ӹ^SVP��_'�Tj2��� B9n��J����>2��#��ӊALDQ�Ο^��e-�C B�!�%����;_���3 ��B_���AJξ  a�Ԅ�YJ����A&�-��!�L����d\�9&ti�@�O����'ev��EN�}b�X,�z�@���dt��U-	}c2�׊$h��}N|���O�>�v�ٱ�="�� C���!j��p���'АE��ŝP_ ��g��U,��
	�'=�e��kƘ����,F�M�8���'ȸŪ�B�@��ؙvID�?��x�'#��;#Gܿ:M(\�u��9?V�y�	�'��M�`���Q�h_5C��'x��1�K#v!������:�L!�'�RX�����x,f�Hec�7ꨐK�'��9�d%�z��㉤_�6x��'N����F�JI�ԁBҮT�j!	�'h6YЧaجc�Z�ڶ��I��h��'��$!'�E�%�`��3�$)�'�i1�B� �P��ָ%7^(Y�'%(�j�P�ƆɣP�� ,t���'��]	��8' �'�M�3�]R	�'�(,���˾2�:%��@�7af5��'�Xa3,��Fy��w��l���
�'d^`X�L�2��P���-b�F��
�'gvX�D	5����1�v �	�'J��a!
�}J�@U��"%ʦs�'�T� �8Ybjp���R���'��5`q)^�1��=�2����i	��� �p!3��	?B4�� j�VU9 "O���L�|��Lb���:!��%�b"OX ��D)2\Ԍz"���<KQ"O�P�i� f��šӥ((����"O@�{�a@#W�L�� r�XA�"O�%�f�<"�yj�?H�� "Of-:6�>ڞ�9ԨY����P"O��:a�[�_8Uj2��>J��w"OtRw�I�$�\y�ɚ�%�� �"O�H�7a�;MՊ(#Eߚ$4Q�0"Of��A�@)5#�z��#�$�Q"O�YBn+X���S��!S����@"O�D(b
�:X����P�)��C"O\�r��B�g �5R�Z�q�D��"O��?
���	ƩIZ�)"O�%rB�۰;���1#��_T��D"O�̓,Y���)v��p�p�b@"O@hcr�@1�|�ӥӫtP$L��"O`l�6��0IМ�ئ�um�9f"O�$S���"���-��_l��$"Of����@*0"RS�M]WSDM��"O�\nb�yv!���If(�t�<�ke0�yۡ�*/���0ץ�v�<Q`(�'%�zl��ŉ�6�pJ�^o�<!�����43U��xx��Om�<����9N(�Wj�.o���Au�[j�<�CN�$k��K2��-gP.�Q�SN�<a�*�\��%�צ+6=�a֮�R�<Q��D(,D=C������S�,	P�<�e�@"@N�p�,�G�R�0�I�<Y@eؽYm0M2&� L�8����A�<�1�Q�""R�x Ø	3L@ ��J~�<ɓ�!R�{�/}Nx��c̞y�<b��B(��Ύ�t���;�[L�<!�$�y�h�
e�}�@��I�<���ܜ��A�!�X@uH@�<ٗ�_���	17���x�z�Q0��q�<��՟i�.�Ҁ��rg���@j@q�<�q� #�<��/���ܙ�I�<)g�Ⱦ��a*���Tm�����n�<1B��A���@�Bؓ-dt���Lt�<q��X��	c�K>�@H񤌛p�<aBH.Z��}{2@	�@ :��r�Eo�<�$��jc� �!�A�ab�ֆ�R�<�	�s�v�x�j��U?�����f�<���
�2йc��+ia����l�<9���`2����ⅮQ�pt�Ѡs�<�"��+���c�J=�h㧡n�<�U/.=> ���#B6�9``h�<E
N�JO�E*/Sb3���g�<����a�`E��c@�yϛ��=�y2H�':���s� @+o�к4����y�'�a����CR�lz<� ��y�dN2X���D�AjT�h�#�ǎ�y�Ϥ��`z�G�eܜP��	�y��-r�n逅j�`�IiԈ��y���&x
a�WC�"+`hq��y�g�Y�R��vfP1$�R�(T�L>�yR@r¨-�7����lIBЮ��y"k�3���ZP-S|����ɟK�!�F9����愀�]S��
BZ�@�!�DC
���`�^�6C������J!!�D�;pL�	��J�l\��:.!�ܮ	�R��ѯM�8Fj<�t��k�!�� �)$-��,n
���B�(��$"O�cF��4s�X�t�
_+
�5"O��I�V�yE!���|���"O(���ë;9P��P��"[0�r"Ox��f�(�~X����)� ���"O�(A*�9Q���yF'�jv��"O�E��]Z�H$��pj�8xP"OP=�#�Q~�I�vC�9p��G"O¸�ǜ1P��D� �<X\̀�"O:�hB�|���ⱋ�(B�zB"OLԋE��)nM9�����7"Oʡ��鄡3�>qS�/��B��!z"O�,�f��3ts&D�hD�rc��U"O"eȷ��"U�ur���=~4r"O�a�ĖJ,�I�!�Юx�� T"O�y����
�v�w�Ӏ@&@i$"Oh��a��V{L(�u�L&q+��k�"O8� i�FD���@�Q� ��"O"0��eC�k�F��S�� ej�"O.��t(�-�P�"��mqQ"OT�N]�e6��*�#�&,�w"O!�E��p�n�:�O��JAce"O�1�jL�L��EKf��sn6!*U"O�tb$EK?.�N]�G熇�jyQ�"O�С��&ah^���Ji�
�G"O��Q1!/cOdX`N����1"O0�+@ D�v��!��ǱZ�"��"O���tbF:E�|����
L�n�+�"OdI"���̃G�sj���"O����͘�r�B�
�a��
"OT�����+=�l����+�@��A"OH-���U�wyJʦc�<uH���"O �VM�?�, ���: ��m3�"OR��Å��d�HE(6A�)��B"O:��VHQV�ł���rRYQ4*O��"�͋6&�0ɨo� $ɚ�'`�a`w�ܯ"�����$'C<�s�'���D�j�|�j4��$T$`��'ټ`b�䌕n�0)$K�,�h�'՚ĉS�D�~�4=`3�8� ���'T��肠�ʬ���(V4q �'6(0��/c�@´zD��v�ќ�yn�D�<Y���϶��AKf#]!�yB�Y�ik�hj¤��� I2&ω��y�O�� @3���j�V��J���yRh64������`���m���y���H(��6#�8	�d	U�B�y�N��|�VlQ;�����֦�y�ML��i�Ԡ׻j�zU	�%F�y2k� �H��"��h:�p�Ǡ�y��
���@�KT�^u��9�A����hOq��9�+��AmԜZr�Ԇd�Z���"O���kO:{~�ه(��xm� �a"O��
���J���	J,H�ڡP�"Ot�#��N�}�Bl�Ȟ�����W"O*U!%�ǅ��p0PE4���#��'���"/J�+���9�D�^�h���f7D�Љì��R�f�*��/]rd-C1�(D�d(��C�o���q4�F�R�#`�<D��G
<o��uG�1<
*�Y<D�0yU����@����lB�-D�Xx��^�*�y�6�X9,����c!D�2�KQ�z�ط�Y)L��X��?D�p�V�U�8v�0�KD�Pn���<D�� �KrF��`�>pk_�5. +�"O� 23.������L<�t�@"OX��j�/ј�3�-գB��5p"O�钄s�p�+��ь|��#"O�\����^��@�ь�o����"O�%pɌM32a� 
�QQ�(
"O�iʓ�ۓ;)��8BG�
F�d��b"O��P4ϙ�^��F�r�J�r""O�HŊ�8A&|S�%t�Xm��"O�q�W�v�-�&F�	�vu��"OPA��V�:L֡S&�#'�]K�"O>\�ƠLAN�$���+"@�}��"O*`���<9���y�❈gơ�F"O�d��@ƥ?�&�3G��?9�R,��"O��X''�/:��g�M'6̪���"O*�*�n4{��������A�F��s"O����ߍ+�L��Q�-�� 8 "OF���D��}�f4�R�·9��5�R"O��`!`	�?��p �L��Jj�!�"O��
�O�$�LP �L�)Pƽ"�"Ox�u�·uH���Í��|E�=*q"Ox���i�z�v�H��P!c(�\�"O$`g�]?E�I�
l!F�%�!򤈝{[V<9笌�G��2Q��[�!�䛻<�@#BlN�~�@��Oz!�D/l^��s�U>;����n��A�!�čXP>� %�N���2�φs�!��?e�l���յ]�~�B���wm!򤜾by��W땫^�P�s�%�*�!򄞀;�x1���	C�N�:w�@n�!���6�@8*'��;#X@���^�l�!�$�7��H�l�|��iA�g��/�!�$� 
������1��`��6�!��Q���t�FM�4�mj%�Är�!�dB JS���-I�0�LTX,�)�!�d]Z�Nq(��G�2������ T�!�dH/u(I9G
J���8���Ⱥ4�!�H�}S��� tP�9��S�u�!�N<����H�CX������1�!�$E9w^Y,m��Ř��	�D�q�	�'K�n�6,4��B�_�6�<���'��%1��2��U(��/b�Y!�'��u��I�8U�	 !)_�=���
�'u.P��??3LACbF<-hQ+�'�����]j�O;9�~��'�`ڵ��9 �t�tK%���'@�Y��iՂ?��cGNUVf@B�'ڌ�X!��+v&�����P�'/��-�,,t$�0�B�ؓ	Ó�?�ReW�T286ͨ>�a�]�P|z��c��G=�|3�eNo�'W�G��Q��x妆�q7.�ʂCQ�	��%r �6{�]�0n�o� �:C��9��ݲ��ӷ͑���U���1u��uj���/M�d)12�H,e��Z��Q�6>~`��LVN�'���j��&8��`���sT�	�ء��A�0{��A淟 ��Пt�?���O'�]b'�< �:�X� �E�'L�#?9Ї�KNh�0��E�'f�K%�'"P��i��,w�)��4�?yL~����Mk�њwd�K����?ς ��*�A?9�u��-PfJbt�$��!4U�u�ߟ](�l�OѮ-���p}B���-W�	|�;H<ѣ�4-=�X�$�׬U����C�+t)K��Ͷ�����9B,�y�b Ϊ<S$Q����w�=S������9�O|�L|"��A&�	3�m�����	Gܓ�?��2�x�H  �P԰V�^b�H�J�@E�p<	�iV6��O�\mZѦ}��"N�O�~�c�c��~N2p�_�$�v�'f��,(�����g�'�lôD�{5�0�
.4r��;��+z������:0�pR3��<d����?EAG`BM��JCzvd��d�nR�Q�`���q�T)8��@���Y�V�ՙR1���Ն����TB[qW�,�,��>��ϒKݖ7-[y�Ș��?�}��˟�m:� �@aW͛�8�m�eBR�+Ơ5���F���<�eIJ# �~U��-�6�b㯓~����AQܴ���������3 E��ꢢL�4f�٤)ƅb��a9�+� v�x�Iџ��	ҟ��ZwR�'�eE4O�^a���H�n�0�q�,@�p��݂��\-l-d$�UH��ɀ�`�+s�v=�f剰Y>-K�K�<iH���?/���0e�^&z��	���\�%�-�q�̛dq��tM�,K�$��
�����`����|�o��`�����榥9ݴ�?�(Oj�d�<��O�j� H�1p�j ��
*��"O�x�#T�`�<��Y
�Ȁ,�T�	�&6�H޴���v� �;�?�]I����	'un�t�ț4�¢>���+�@�äA�'�T���h���M��D	#�U�vD�{^�a�.�A�,�q��>�(O�M2��M~ �"��`yz� �A���`ȳS.���%Qc�*Dx��A�ƥ��ȰT �O�o�(�M�۴n����d.��׌�~�R��6_���	xy����zQ:��M�:��E"��í;�@C�I�^,�b���4Y�4�hB	өj��q�bA�5�'�
U�.��'��4`PhlZ���ѧ�,0:&�ؠ��~62�
���?�Ӈ��9s��q��6�uе�I�H��͜$0��'e"�}��	U�t�ք(o����$��r"ѦA�9@�J�[��k�NX� *,m�ے2�� ��`�=�\8@���bJĀ�ٿ�����Ɍ�M�f�����T�N�Mry�`�0�X���%��'��|B��<����u
p%Z�8��9M�x2.iӶ�n�I�	r�pqч�)R��m-p���1���?�H>���$ׅS� X  ��   ;    t  �  �+  �7  �C  
P  �Z  je  �n  �x  0�  t�  ܏  T�  ��  ע  �  ^�  ��  �  $�  ��  1�  ��  ��  �  Y�  ��  ��  ,�  x �
 g � � 1$ �+ �1 /8 U<  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}��za�@AIp '�`iF�'�ay��D�3������ ��4�%�x��'�za�(Nx�0�A��Y*�Jד��'08!��~��Y�O��Q��,�ۓ8�>�O�q�Axh0:Q)0W� P"O�H��/r8���H�<+�E����<������KO&�0�WK�qs���1b!�D��/�*lx��K_���R*Щ*?�i����>E�$Μ/2����@ΐjG^��w	�M0!�j��؈u��C�pT˔�M<���~�C�SQ���'�@��2j�?����Q	I�"�|(#���'�r�BB�]35Δĳ�$Q1OR�d$��>�Γ>�"䋥K�&\�B�� �c�(���	Y̓<���`G��5A������dV�C�=�S��?�e�}�6=��%W"R����r/DߟG{��I�6�R�T4e�㳊P�9��C䉺e�Z OK4g.���θY�JB�I�'�)�!�`�:�ѡ�BA�C�[��y���F24�$�d��'�B�I�[ǆ�IB����٘b�ȼz/�C�)� ~��NP�� QN�B "�x"O, ����)��U 6n�~��م�O8➨D��O԰��OP�:�����b�	�'�B��M���!@fGo����	�'$jE�*�6*���mO�g�f����HO�|�5�H�QD����mV�l�����"Op���1d@�@��y	>=X�"O�}ѣE�d#�0v@$S� l��"O2�:!��M@�q� M�2�x)�"O��E�[�+�� ��7/����"OTP��&
����n�|��+��'c���å�+|�Y�F��K��q���)|O��	m}�a�2P�-Y��L�Bg��	��HO����!���|�q0�ף��Div*O|r�'J).�P��Ob�X�	�'sV=���Z�\X�d��@�H�tt��7ړm�<@H�4[�,u�gN �d�D9��l�"X'ԅ��J����"*Ͼq�@iG�~M����l|֑ÅoH�1u�1�Ā�����g�]a�=��.�M<ҙ"�ҟ"�2�D{�'}�:��ơ^���箕/�J���'�T́�S���07.Gy�����'W�����0bN��!���iQV�Q�y":O���9`�A�B�X-��xB��5mf�~b�O��h�&�j�]B�"�X���jp�K���xb���@|��@JrHy��k��0=y��[�2�|��ҁW�ZxiR�V�y��')�x"P�ڳ��H!ܬ�iۓи'\���S�G�(<ĸa��5m��'o�t�wG�b�A0v�z�xR�|B0OluE{*�
k@�=.�P8`/X�|G�h�*O,e� ,�e��eHg��hg`��'H�ʂ��.24b@���2[�t� �'D�|f*C��̰�$�Y�ܡ��'w��"!�QxJ��E�$[\�
�'�Չ�E}����P��y�'�h�;1COs�<�ا�*y�^�8�{rmID���h��hF�4p���ɻw�L�	�'�l���K�	:�v�F�^=fͼ����	�z/b��|�"�L� �� #�N�ib�m�����y"!KD	ʈ0��Ķ.�~T�d(���M��OH��MJ?㟬;`D�	]��t
�L�,$A!1�&�O��	)6D�@���:j��1���A�� 
J<A�OD��D�7.��f5`ޞm�Ag��O�@D�d�ط	�������6e�R|ʂ#.�y"P> '�<8�7)�@�"mݳ�?AUX��&��g�+R^09DM�DD|(Jv"�J�B�IX����@�ɪL3��Y�ˋ�df�����ɳY�PS�
�1����P9�B�I!
o�%�%U$����S	N�N�B�(h���K�4����g��]�dB�	u�����*\x��
�+J��C�	di$�:��X��Rea�m̫C�ɓ%�hUA�E�^2x���D�RB�!���F�l�(�z���0�Fb��9�aKx���'=�Դac��_�ȓVӐ��eԗ�i��ÇT�4�Gz��'�`��0U��bC�2]��q��'��)H�L�+^\��R(�<?�^��'�P�!d��$�H����:�6B�'�����M��X��1iV�A�0�x�:�'�؜s�ҭ �(�Uሖ+# Aډ�D$�S��kUj�d�I��Na�H�����p>yL<����:��	����d�U���
��#=E��S�? ��r�C$NI�jؐ ��)����<3���O���e�Z�9uh�Y-R�v��9��'ua��G�D@%˝�Lc*P��c�yJZ�i�$DޡH�N�VI��y��
�W�h�0�#]B)|TJ��Q0�y��#�"�"A��6Bx����H���y�/�2�y{W���P=����C3�HO���D��М=��,#1�Z���,��q�!�к֍D8z���ҰM��A�֦�Px��h�=�`!@,�C̊��p=A2��4t,Vs��'Ą��eF�pU!��IQ��%�G��!,���+杋RT!��J�[uj13b
!(~��kDd^;s�5O>�ip�Y�g����B �0U8��W"O8y(vվ)��-a1��:*v�Z��'}�'��R�MZ�M*Qh��+A���'P@�G[�nC�͑�)F6�%k�N�'�ўʧC���sЯ��+@FӀ�E,y���ȓq�������X���Wa(���s�$;W��NK8A���3H������:D��q�.�7t6vDj'��1>��2E.D��j5�6;%N�)�LEY�A��J)D�)�L�!�P��L�
�Ա�3�'D�p21kT�|�@��SI6,\y��:D��h��&ahy�p �=&>I��9D�t鷌^� &�)���Q���qd8D��0*S��4���d�7H{�|ڤc5D��P��
�+A4�d�ԛV���fh0D���ƷsG�SWE^;dF��Y2�9D��r'�B�� �#���pxv���"8D��2�K!do|4($o��7��Dk3K!D�PYWm�V�P#œ�|Hd���?D�{f�P,x$��7mͰbN∫@�;D�L� ��s�,�p��M�|����N,D�X��$Y�,i9�C�,/��0D�&D�x1��N'R�ܳD�	oD�WH&D��(�"T�1ȝ�pe��[�, �H"D�p�K^Ɏ�8��=BP�(7�:D���C���.�Յ��%9@Ipŏ7D��!���f���"'RcN��Q�)D�$Z�(���1¨�?(����0N#D�pڤ/S9O��j��P�VLZQzס!D�L���@�C$e�Sg$0M�f!D���&��,+P}��n�� �g�9D� ���\$(q���V�$WΤ�P�8D����Q�s֝yU�ίl��S�A#D�L�d�]�R�� �� =PU� �?D�$2񏕍Fƥ���/Gԝ
��;D���b�^�9��
'O%ͨ}��H'D���0 (kkb������=�%�$D���U \�A,��G�g'�)*�!D�`�2�	6L��gD-m����;D�\9��� SY,������`��a8D��i�o��h�b��_���C��5D�0�"̙4l/�P�������2D� p��� H���8����MW�-te-D�, 1EP�Dʨ���ITP�|��),D�x ���k}����"!�Y
�A5D��&+ê �P���J�e�>�2�5D�x��6��M��>A�q鳌%D���G	 �bP�"_=CԬ��D8D����	�8u7���a�R�[>��j4D�����fzāC�/0�6��6�0D���g�lT0UJ�#�Wf��L0D�� ���;X�����%<qZC"O*����=4��]�����Y=̨c�"O�UA�a��!Z�%R�^����"OT(��#g�8R.S�gD]�"O��%C)�v�R�5*���6�'d�\��	����I֟���۟H�I�����$�7&�m��W**���ʟ��I���	���	ȟX����������")�.H� ā��кt-(���Ɵ��ҟ���Ο|�	���I����	H�zasuJU�|�gJ�:��p�������Ɵ��������X�I2���#�~�.�"$@��
�z��ǟ<�	���IПh�	��4�	��0�I�kVJ�`̉	�rx��2M��	ǟ|�	����t�����Iğ �I1��3n^�M<.1��j�$��<�I�p�I��������	˟���ݟ��I{$��u��%%���#�lR�0����I���I���Iџ��I�P���I''vx�e	��4,��/߂ߌ��	ğ���П�I��P��ٟ8�I���$)L"�p���3��x��@ ;�4i���P�	şL�I�����\�	ڟ��I0T��Ѡ���VA��1rO�S����Iџ@�	џL�I쟐��ߟD�	�,�I�8�[K�C*B��3* �
���	͟�Iޟ��Iʟ��̟��Iҟ��I�j��l`3�j��µ+ӈ4�6q�	ٟT�	���֟�����ݴ�?��S����EJ���1��[ae0���X���Izy���OB�mZ�U�H�	�h��_\"��h�dY�4?Y3�iu�O�9O2�n�.	@@f��6��u��X ^F�y��4�?��d5���'>�Y�5JG5I�b����I˧c�4a�nâ>���Z��D�O���h��9b2-��@�f�Z����,qKB��p�5�}�'5���w70U��m�"�ٺ��@v�\�!w/s�<ho��<9�O1��e�dO�=�� �C�p�ç��� �	������hsj�{��Ph�"�=�'�?9Ǟ<��Pss$�%Lh��Ţ��<�+O:�O� n��#x$c��ZT����VJQ�M���6�Vi����	5�M�%�i��$�>��.V"Ӹ|0�B�QC�͒��WP~,m�.��%�M�ӘO�:�iF�S�����P�ƹ*�% �5Fa�)F�&a�']��"~Γm�ͻ�ˎ�T��XȰ��-W0�Γ����P���Ц��?�'&���÷��K���q����@�Z��Mi�^���u�6������F$Ґz�)!e�"b*I�G �c���8�DƧ{=%F{�O��IO�� cd�M��O�EL�T��C�����VF��'��jD�Tm�/�b)��NN�:}f���&�q}gy�d1m��<!N|����?�C=[�4������;�040��׷;箅@�iI`}�u�=h�-��O��O>�'ij\B�a_t� S�A�[��с�'�Fy��|R�f�4���3O��4�Ŀ-`p�e�=��̊�8O��n�A��|Γ9���IvӔ���f�x�ː��bz8ti��ʯ3�$�2«����5;��:橔c�t�C�O,�Է� u�Yc��UeG)�,t����sبК'T�Y�ȕ����ĥQ�U��{��טG)v���$�צ)��)?Yu�i��P����l���+��E�!`n��T�<��O�	mږ�M�_^d�u
��<�3�(!r֐�!˃U�E��b�
U\\�B2�վ&���i�`P���	���4�V��?	����EBv�CХ܅;�[C���<QL>!��i�q1�y�V>m�0%M�`u���f�X7b����%?��R���شM��2OP���ɔ�n�d=�N��zp�*D�M�*1*�s(�3,��\"E�����bR�e�T�^n�5��ء�Ϗ��5!`�E�A �,��ڟ���ҟ(�)�@y��j�~�0�L&F�6����0����F�9��I'�Mێf�>���i�v%Sr�J�d�pȈ��B�l� �L~ӼTmZ%'M|]��`,?S%�?|�$���K����6OtF�X!�̨���ݑx~��<9��?q��?����?�.��y�E.T����-A��@@�ئ""�U�X��ޟ<'?�#�M�;]�s��U_��d��uCx-a��i�^7�����ק�4�O��dN��&��j�'�!��I�P"x����1b͠�'��4�n�'�y2��|�^�l�	៰Ѥ�	��[e��O�u�ū˟������IVy�ed�d�'3O���O����.!0�f�0(8J@H�=�I������a��4c�RT���)��0�v�u��F��R!?Q2�Įn��@��;��g,00 ����?�B�4fR��&f��F��[�A���?	��?)��?��	�O�d�F�q�`iiT��'�^�[�n�O<�n�-��і'�(7-#�i�E2!JD5l��$��cϤ��r"y�T�ݴ[�&�x�b��ŨR	Q����c�Q+�%Dx�毂 @^�5nM�
�n] 2�Y}�	iyB�'C��'�2�'����֒�9~�	`�.4�8��.O�}o��ksz�	����I~�s� wDR�U:�)�sA�t�������D�̦٩�4�R铮AW|ݻ���#섽�TCP7����6���tؗ'�0�[��S&Xj���|�U�t,���CO��q}�E�){`��O���OZ�4��˓/��։���y�%��j�� `�j�;��M��[6�yR�`�T�d��O
�n�;�M"�i�)Q����U�ٲCn؄� 2'˪.;��j�OX �Ӂ
32�-ѷ�/�ɔ�� (��p�G3XPܼ�7B�+1 �{v2O|�D�O����O��D�O^�?YK�ȂD�@��iA
�#6*��x��ҟl��4Ğq�.O~�l�W�ɼ�Nr�ꗅY�mh�G�N��c����d[¦���4�B$�X9l7�\��?y�������2����6,�2�Fv��|ꆌܠ/吩1����O���?Y"�#VT���@�?k�<�F���<iM>ɗ�i{D$S�yr�OJ�DL��V�Ρ���F�Á����DD}��j��l��<�H|��'c�b�`�kANP�
f(��:@F���*�T��h�$OR?�ֶT�P0��&(� �Ok��N�Y�5i@	ќ��䠈]�n��?y.O1��I��M[d�M*�>�I��I.]F���&]v~��'�6M�Ov�O�9O��mژ6֨�s�Z�'-x: ��"� %b�4�?Q��}ϓ�?&�ضnGN��`
I~BLZ�:�AS#�|c��cWGޙ��'bBW�LG��(������A1�ш�.R*��7͙>S1O��?�i���	�.��c	����j�Y(2J��ٴx��3O��|��'�?aA�8bf0�k��Xa���+�H�87�#\��l�S�؁p�ϕ�pE*1ʍ�4����]�n):1�ɳ X>L��甇X2�Ķ<�H>�t�i|�A��yRF�o���@Ră9�H�ʳB�T2�|r��>��i�>6m|���'�:�b㈃��"m�oS�@�P@�'��)�>O�"�	��I������m����
*�䋀ƶ}����Z��@Q��!5 ��D�O��D�O���!�'�?I�h5� �/�%]��"��?�ѼiY�ل[�T�޴�?�J>�;3�nAu�S�<sԸ��O)e��(͓1C���bӦ�oچ66�bv�n���I
t���h�Od -Ю��P����	����h�I]y�'��'j2�'�2�/7ʨ���I�4'�M��e�剬�M; �;�?a��?�L~Γ=5���e�Γ|�p!CX�O,;$V����4R�����O����	�>@r4 #��)q��=G��б�l��g%t����<�B�Ӥ	��t���䓈�$V�IT����62��0��ї*:���O���O��4��˓71�F�˕�R��4����+�'pl����y�'k�t� r�O��m��M�׼i;��r���:`&�NH/2=�(�+˷�*�3�'�r2-�*��%�`L���?��_c��9pf�u�P��e �'\�xH�'f��'G�'���'��:�@d��0ȱ�
�cN5r���Od��O*ToډFb
u�'�J6�"���78	詡���F��ЁE��ƚx��Z}�	b�<�lz>�h '�7���9�pYYcF@�Z�vX�p�9xv����+H ��Eϓ������O��d�O�d �@ �Ԉ��� �H��oG�����O^�
U��M��y��'�S>=K��І
 ��a��K�8��(;�k1?��S�(r޴G��&��Orb?a�$j�����f�	l��p �9J����p�+i:�}���d�K�G���ig�|���C�Y�j@���1�_7���'���'����Y����4Q=�ЃFÛ�kY���I��;����L|~y�����O��m�4B�@�i�4e�����;F��Lj޴뛶�%X�@��OF��fl��F��HQ��<�P�*�����֗�r�I�K��<�*OD���O��D�O����Or˧46�z��	5)�(�A�LH�ٖ�`��i'�h��'���'%��y��q��Έ�7X���(�E]�$����8-	�l���M��'�)��~fL�
��}�$�(��r4T�D�<��P�}�h� �<[��sKM[�IYy��'���	�X�Ɖk �7*�ʁkAfR9 L��'W�'#�	0�M�gY�<	��?!&k�fB��u��V�����׷��'n��F���k�h��W}�N��"����
-���	8�y��'� 8�K2DÒ���R����T��{Nԟ��ЈR�4�0��H�)����h���\��۟d��ǟ|�O����ʟ�.ߗy���@Ė���i� LɹA����Ħ�E�}yR a����n�����8>&8�$:�4�*�M���il7M@�y;�1OF��� E�$��"΋6��y��h� p٢4�VF�=Z��}�6�2��<����?��?	���?!A
@�r=4)���L�{�Dx�	�����O�����A!'S����O���Ħٗ�yb�W�H)x&HvF�!SU���o���$�fHp��IZ�S�?��E1�cc��T^��ύHk�|�֌3����'. ��q��nZ��跙|RR��؅�	�G�>|�Ff��!���f�ğ��I���ܟ�Hy�J`�v� ��O0]�� 
 ׁ�0��Ŏ�<��i��O��'ɨ6mTΦi��4v���`�\F@�2"���=^i��n�e��m�'G
�)fa�2?@�����.v�U��R-G�@L�4�ԄF�D�d����ty"Z�"~j�		��,��e�<A�P���̓\�V����3��d�¦�&�lY�4n���p��S5�	9��<�O�nZ$�M���j�V(KR�L�<��8kEyh�&萚Ԣ�;�:A� jX�K���Q�)�hO�ɮ<���S�]+��)��qBS4y�Ƹ���n��v�ӵ�'�哮tk��ڐf�~7�тO��7�P�}���/�MӃ�i��$5���@
$B�:�����x#���6, �-�H �]����?���ʞ�s�%$��)�g�y��H�&C�h 4 �fWYyB�'0�)�3?Y��i�`=��	ikP�D�G!j�ȝ�������ڦM��o�i>牟�MS!ڥ{�r|�ы͘q�r�����7~ӛ�'�@��p	^�y��'�4e�����衡�O� @٪���C��DO�:gi t�d�O ˓�h�����\����Fc�-&� �Y�����3��X�'>?��w�xH��)�<)iƵ9� �~�����gӲ l�<ѫO������D�-��5��7O�����t9��f �N��$!V9ON@Abc�
8aN(�$�<�'�?��
��a�N�L�P��i���?Y���?1����ɦ��។�����XU��Ȱ�qbܬ���qӄTL��G9�I��Mc�i���>�7(��"�Q�(�<���"%���<�!��O���B���=j��1��u7�������4@u���4].P����ƗXu؍x�\�N���I����ǟ0��{�O�®ޒ]�l�˴�҇��ղC���)��kq�FX���<� �i��O���B
����	L2g(�`x�iM��Aj�47��H�$��b�'�XC�'�F� �a	!�E�&��>c](A%�I*)124P��>Y�
�<Y���?����?���?1ǭT�i�6ْD J��b���]��WΦ���Fퟜ����\�A��'�UC��?w��i�&�><9��`�>	B�i��7͇�&>)�S�?�'"� C8���A'S�q$�]�A�C�#���	�Dy�B+!�Z�٣�x�'��ɩk�5���*.��#Ӄ�����۟�����L�i>��'��6mA� |� �Sf�e��R3��i��[�DE��y�?I�]�Tj�4NP���p� �I*Ǿ,v �V Ԏ<"�4V�̍=π��9O&�dH�@x���G�v�ʓ�
���l���G�Q��ͪ����1OV�D�OR���O����OZ�?0�J�1oua�,J��#%�t� �IԟxJ�4%�L��'��7�3���/b�f|:�C����2֧ٯ'����Ig}��|�|�oz�6�jb�]К'���!W$.��W{��	2�7 �I�c�
;B�v�7�|B]����۟�I��Jd揌k{HtC���XZ��R����|��fy2�f��!R ��O8�d�Oh˧<E�)�d�0^Ra	�cB�]�'@��f9��+dӸ)��V�S�?5�cR�!����e��VM�gJI&o���W�S�j`�'�����,bBe�1�|�iT2~�41�B�cnV5;J#���'}��'����T����4[c&�Z��Z sGb�
%��B�:(p7�_�������?IU��8شONP%��i��qP�(�<y��iQb6�B�l�1�;O���H �R<b" ��1Xtʓ	yJ�
B"Þ6���ѕOL�"�<����d�O��O���O��ġ|��(Ò���D)��]�&$heA�:���AT���$�Od�?E	���5�Ϝk�|���*�(t���	9p��v	����|}���"��`��4�'Ҝ�ĝ�f?\|�F(��e:�'uܩ��M-T��X6�|�\���ğ {Q�B �#,_�q̾hB����Iٟ��	vy��o�ʁ��?O���O`X%�ҪB��Ei�bB���T �I*���������4I=b[�d��YM(8YpT�9$�p�d���� G��ݒ�"�E0���'?�dN�x���'Q�%r���l�bp���̤��!P��'�2�'|��'�>M�Ip�|H ���u��q�N��U`��	��M���{~��v�z��ݩgJ��˟�&&�E0�lAp���ɟ�M�E�iF�6-$$�5S�;O���FFVꁒ!T2_KI��:|�bߵ(�@B�&�b%�')�	ɟ������Iȟ��	�9Y�T�SA��dx�ţ]P%�'��7��(���O2�$5�9O�F@�7sm"6��D�����A}}bLz�εnZ��?�O|����������S�ނ8�Ras�΅~r��C��B�yR�69�|$a �!G��TK��P�P�D��mR�jU��YS�@+a�Ο`�Iןp�	���Uy2�`�@�6O����|�8�;1�@�6YZL��4O^\lf��i@�I�Mk��i�7-ؕ	���Č|>4�Ɗ�:IabTπ�K���O>�A!ƅ<��:�ģ<��aUk�H,`���ЁA�8�@�'J��OZ�D�O���O���(�ӖJ�N1�T��rL,"�Ó&�pd��ß0�	��M{քP���ߦ�%��В�H8�^�3�DF쁓�dÏ�?��O��o��Mc��8R|�C,��<�� ZB`x���ǠԊD�vp��\�{KiH @�!������O\���O���Ƌ-�p����� W�:԰�kO"�����O>�*����ōf���'2W>i�f��#82� vj�k�n����3?)6Y����4M��f��O$��I�#�� ��N��h��확�X�yd�z��e�tŻ<��'V̤��!Ǖ��g�<(�"��f�H�����[�$�����?���?��Ş��$���
ө��e4�Cg��'�|�i�l��0���'�06�-�	����_��92�B���5E����A�m8ٴ$<��BFn��%
�'N��G43�\�g�SX�	����Yf�&'�s��]�!�\yr�'���'P��'�"X>�����?�܀���
�Cx������M�g��<����?�M~Γ+l��wh�p�$'K[���r��l��e��a��n��?q�O��8���3��P˄1O�GF�0H�J b5�z^�TBQ>O��V��2c�4!��"���<���?qSd_R6��1��,iDj�Բ�?���?������¦5`��v�|�Iʟ�[f��G�4@ȂE_� 3�0/Y���'����Ojo�M� �'��Ir�Vy���C��u�m��L^b��ΟX1��%',L���JZy��Oe�4qSe��+�(@�rD��
�ӂ�A?/�r�'1B�'ER�⟌�s�	(ev%˴�A�	�p����(j�4t�n�(O��l�㟤'���_B!#�-,
�xZU�)
Z�	�M�³i�T7�K0��r4O����N�h��T%�}�� bm��f��ceC�>�2��A;�$�<���?���?���?q���8k�$�2fhO�@Sܩ��*�<��$��%�"�������`��'٬����3��=1��֪J��y�V"�>�i:�7M��&>M���?Q��D�8U�QK�6"�p��M�=a���B�_yң��B��Ӕ�F!=�'�I9U��3�c�"'?Irt�M]I ��������i>9�'�f7�Ϯ�^�ҝ7���"���+0)8}i0�e}�d����?y2Z�p��4��&�n�4zҢ
�/렩� �8a��y�Cǔ6'd�y��<��T�b� ��[�)���-O(�I��KA��o.hD��G��+s�|�w���<������<E��	�b((���$KU�\���CO��'�&7��(��I,�ML>����d���#h$�B�AP+�y�^�@(�4�6�'DB�y"��)�y��'�rjL�'j�>�pפ�Br�%�BP�N�@Qb�)�wLў��\y��'],,R�mŋ-6X����=��a�'��'�~6��m�1O����^�����rP�"��V8x����O�=lڻ�M��'��O|�to֩,�*�A� �z�6Y����u�
�|�u�0�;?!�'�\��A7��{��u�0�;��ӥ�6Q(|(�/Or�d�<�|�'؎7�B��PJ��&����8v�L�i2���3ٴ�����'��6핫X����$+��
�!b�dˇ�H�n�ʴ�TE�R��۟{�WC(}s��)?�T@KF���۠A>4zٰ'iCw̓�?�/O�}���w,!�EH8"��x �+�4(-�F�Α��'~񟸰ozމ�C�"S�hP�'��H�<��Uj��M[r�i�d�>�'���t4e�ëT�<!0��2i'��8M��}�1���<a@-G�L(hl�4N�'����4������	r��.�|�q�Yr�XcG��O���O�ĩ<aQ�i|���'L��'r=�#B�e�DU*�t �4'�1��'aH�q���xӦl�II}R`\�`���O39�R#�O��y��'��hA�z�@��V����3���S���t�Ê�� lP'�b�L,��@�0�������|F���'�����"����BZ!w̎A�7�'��7M��7Q^ʓs��v�4�� R͊�U|��Pw�^��j���0O,�o��M���iQf��/��y2�'������;qJ����˲:?�� �U%A�:��IM� 6�'���͟���� �I����������J�&t�8��l�
X�Ѕ�'B�6�ޭR�P���O������<���BsV���T��!I�*ت�&�8b:����M���iw��d'���`�I�]0>��&A��Qp�1�&Q#��Q*Ѭ>��˓Z]���%V�G��ћL>��O"\�F�q�
��:��-���'f��'����DR�4�4X��H��+���+q��%�l<�$��(�̓h@���'��'-.�+��noӨnZ Csb@�ǌڄj�`�R��7>��+�aI ~�d�ݟ��3�ʞv�X�Z^y��O��X555�5A1,y��5��	ӟ��	�H�I� ���O��1�DED�6��1I������'Ur�'M�6�ߗy�˓Л��'��AgΕS�#X�Lh
��L����d���e�޴�?y2���6`��?�#��(p�"ٰ��p�IYƞe[��xǜ����W�Ay��'o��'@��=:��	7��xl%q����'��I%�M� b\�<9��?�-�:��_-�HŘ��0��8�՟�`1�ORnZ7�M+'�'d�O��N,"�4�;�k���FH��i���� �I5'-�y]���S��l� �j�ɦ^Kpi���B�,=ĝv��{�nM��ǟD������)��jyBp� �P��]�o#D �R��P�`�p�R?�I��MÉ�@�>���i�FTq��4#�ҩ�"�V,�CLmӤ�lڲv���@i�<�I��6�Hk[X��'��d�H�T>%"GGFP%�'�����0����	ğ���@�DH.�9�с�0
QlC�&�7��#M:��OP�d0�9O�Lnz����K�ox�XI��,��W���7��������4��I����4� �f����f8�qm8#�� R� Zz��䁓9�"�b�N�#�E�|2Q���	�xB��ecp�F�!�Ѐ� ��p������\y2�~��i�.�<�����+V��:Tl���յI��ˉ�&�>)�i��6-Z�P�'a�]���]�#>ԃ�ߘ2Od�(�'���@�G:c��֧q�	�?k�N6X:Ɓ�	�Q_�<j5��:ں�IBߺM���I���ϟ����
��2˰q��+��X���t
��d^��1�"�>?��i��O�[�������	�����~��ۦ�K�4^~�#�}Z�ʘ'�2ʏ�IH�\
����N��kͫHStv�;5���|B\�D����T�	�(�I�� R���>��([��Q-#*riIb�ryR�r���b;O����O�����E�R3�\�߼�x���<\���''p����NE�7�L���?���܂���	��N-�4٭��T1�Z�=8TI�'�z#�K�V���RՕ|\�Xa�&@�=]8��
˾�z�	ǟt�I����I���fyҤd�*=ST9O$���@`?���"ٳ|��D�8O�l�u�y�I"�M���il6�<+��C��!h��$=:�(�K�=��$�O�УA�,d�[A��<��'F�k�G*V�h�$R���q`N�/�$�O����O|�d�OJ��:��d�8@���dy�-!�H϶0�4X�I�����M�������禑%�lUG�^sZ���[.I�\�A�D��?�O�(mZ��M���~����yr�'�D�;� �t�!�-8.�p[#�ӻxVHq��֭Q�|Ū�B$�$�<��?a���?y��C��̡Dm�E�9�f�_��?	���$���A�d�p�Işl�O�l]J�@?E������!�ѡ�O��'Gj7M���E�����'���l�'�\q�',�D|�X".�3ϖ��J�7�RH�/O����8@6� �#1�DU4~��;�Q?KBך�(b����?9.O���	�<)��iB*�GE�;\�����,P��I1��R5����զ�?�P���޴~5�|���I���` aO�>d���ǷiH�6m�	xIس5Oz�d��yZ Ƅ��
ʓQ�ةB�%��u��;s��X��E͓����O��d�OF�d�OX�$�|Z���1?T��c�9�@-�%g�2���D ����O��?)����6$�׈����9{0��S�kH
���sӎ���M}�Oh��O�~]w��*�y��д'��)�e�j�X�&a�1�yr�"/�rHjՠ�!nk�'��ڟH�I��&!>@�hL`�k������Ο���ן��'�7 o9��D�O�D� &R]" Ȗ�^{.,����wW��0�O��o��M���'|�ɏR ]�sb>��PK���e5O�$�5*�8�"�B�
f�ʓ�jD��	�`����.�䁨�e	3tXL��r >x�ֹ����?a���?����h����F'�$���$ъ�,�KGdۺD8~�DW�X��Ey��k�z���)��!*a��s�U���4>�	��M3��i��6��Rsp8F0O��d�R\9t&�2�4�&D�9H	�)ro�&)�8�T!.�$�<���?)���?Y��?9ϳ_Q �e��E�2��t����d����ZT�D�4����&?�	blh A���!`��E��#��(v�`��O��nZ�M��'��O����O�k�Hդ5r�ʣgC ����5(\�htW��Y��Ր.�&�@5�G�IPy We������E.b�`]��Ɗ7H��'v"�'&�O��I��M�`E��?i�)�'�f�;�"�O�� 	D�<�ŽiF�|bd�>�B�i�J6����Y��\�a�,%�3_9i�6��@�;b��
n�`�I
n�* "��өb,��'��y����~�0�ZS;5��A8ЊI�<����?���?����?	��4"̊W츙�^ �ji٠�GT!��'FRqӄ��Qj�<�u�i��'�����]����^�,�����O��u��An�X�Iֵ0�p @1OX�d��e�p�3Ǚ|�`6 i"��)gC�=q�Q�Ҡ*�d�<���?���?�qn&��1���EX�`���?����D�ڦ�3��s����`�OK�$����"��8�� 'E�I��O��'*7mŦ�(����'����J9�<śV�a���PT�%�.�R���34!��-O��i��ܜ��j8�d�D�����Lj:i�DiѶEh����O��D�O���)�<a�i�ja��W�ܵ�L�Ut@��"�Ɣ���G˦��?�W�H��4W�Ċ�#�`��r +x�"�iH7�O�n�ȧ����-�PZ�\	��Zyr�8lA��;?m ŉ���y�Q�t�	��ϟ|�Iϟ��O[�@�@�F�6���c%S��0e#B�h���(��O��$�O�������$OV�mxׂD�kYPsdf�NWH�ߴm��v��O��|�����VI�8F���ϓu�!��HȔ�T�a�<OK P�4�1�6�R� $��O>�.O����Of�� �m3����lq�f�ia�O����O�D�<�Ҳi&�0Y�'���'���� 	�v�k��(](��i����E}�"f���oZ��?��O��JB�	3�x�1c�2|�v�k =OB����<nP�
�-��.6����n	���Л'7��2�D��B|�;��#w�����?����?����h�L�������a�A�69��h�	K�Zɸ�$Ӧ���!WSy��}ӄ�D=�4���p�L��%��>8���N��yb*r��m���M��(ʪ!�2�͓�?���
S�5s$��!:�F́aH��,�	�nև5�	�y��X��,
�-�<>��ِ�P/Oϰ`1��1D� 񳦞:�@a�M��B����iQ:`���3lB/�*ɋT�˯'�>uC��+�N�Q�/��V)�,�ckV&X�`Ӯ�4$�\�ej ,4bJDt�E����LX+j�.��c'G�O�t�!P��"��e�o& J�X��B��-1$� v�� V�Ql˪$���x6b��@C]��y�f�j�����O�$��U�'��L�q�Z�C+�][�m��lZ��4�?a�@nt)���?�����|�1A��a�M��}�Ͳŋ��{��lZ�(~�e��4�?)��?i��0։'���H�&��2�G�Yh6-l����O��d�B�'�?���[
܅{�#ďefT!:E*~M%2c���E����	=`� ʏ}R�'��	��T���싣���Q��̫����'4r�'x6*#�~����?����?�`��%oTQ�ㆂP�z�cH��q���'&��:�%=��џ %�֘-$9nUڔi��P �e���΢e� 6-�O�m��O�$�O�([��V�\���REn��}���ѦCJ�e��)ߍT�TX$ƽHT��c�`���4YQ�b�d܂����)�oWP��G}�jF�yK±S���n���	$�=k�N�j���>xT)���z�*!�-��X�JBŐ�eP� �*�E�jy+�� �I���N�����*��d������(��УPAԩ�6�5'�6Et؅�H6l�
��bg=5�
��rgX12��QѶ^�pAID#+��2U��+Z� !�ߨ5��`��?Q�Z�&=�R�D�6xp`K���#?d�FM�� \N$)����  v����,W#�1���b�'Z2��C�s�T�s�$~F岀ӺS4�r���Yjq���	�q֨��I_�'�,�Q�w[�>iJS���8��R�<�K�"D�� ``h��M����8plI��LE{�ONO,��þ�Z\�d�_F�{38OJ��Eh�Ŧ���ßL�O���p�')��'B\e���5-yV�	�_1 ���($%�=���s���4�>�J#�Ux$����.x1�'"(zԙs���6��yQ�bG>",���A"'��*O��AG��H@���%����A�d��ņ1P�L�"-�3<t͆��?�7�|���'�]VɝT�XL�a�ך�-�
�'�h�w�Ձ'�$�e���`}����S���T�'�,�눆	�r1s@�[��a��'����p��'������4;�N�O�.�n����5�<8�Y�E��K��^!�\Y#/_�Z!��ןM2�Θ'��)Rp�̸7@�#J��k�a<Sd&�Kv#��sjF��oU)Dy.d���L��5�I:s���c��W�K��� )V7Z,�ɲG��$@؞��3C6S�\��u��5}����c%D��,���@7�ނ`�tTz`eZ�7��y���4�|�O(ͺs��æ�Y��W\��Ȁ���1EĂٟH��ӟP�I5i$��	Ɵ�̧4nvŒ�CK�cP|�R�i��@��3��H�5�4���i�2"�V�DF�UJ���>ʓ"�0��k�+�V��Ė�]\^A�āD3@e�%s�l��7,lQ�ƅ�|y�4+鉸Ú�D�ۦ��ƍ!*�ar���^PE#g� D�t*��ʽq���A��u�p ��4D��X􄌘y��y��+�+
��pX1Eq�tbش���^I�P?!��@�4�[��$<k�D�*[úh!$ �B7ژ��'@2�'��YǥI�2��b#Ð�k��T>���I�@.���( ���W�.�\J2 �Q�E c[ أ�+ST�S44��#7(�¡ ���Q��<)!���8��4\
���l�%�e��R#̈́9.Q���4O��*�OΔ0�'^�/�n�Z�L8ShF�T�'�>O:@��̐�#��lq�+�V&5�2O֡R6�����I���O�v�µ�'���'1FmaǃϼV$2ك�!�u@�Dr4 a��iYo�b��U��<�O%1�r鑜0y���p����a����uhС��>Ԍ��)W�n���O���P�	�0p�`ՠe�����߼����UO�)����Џ dRd�që
=ju�p�/D�l�3e �EUF�Z�(F;XgF��*I���'~~.u��N�>�L �!�#J��8��?	��y��(����?����?��� �4���2�'
���%!��:��H'���J��^\���%��t2�)�?��L��y��T>~t�r�c��QI�DRd�ܯ>��Eʴ��*=Hi�A �w����O}�阢��`�qQl��f!͛$&��nW�����k�L�	��M�f�x��'�R^�p�w	��B(�.ͳa�(���	?�h�I�V��saFk����Am��
:�Y���$��@�$�<�6�ٳ{,�&�
A����a�I�ؖȫ�!0��'k��'�2) s�'��0�8L:�,ښk`$.��6�9�R���Bd�Q��+�8�jr呃� �!��:�(O�(�Q����5�ɉE�1���D4A�3J�JZ(qg�_;�MDn�8t�qDyR���?���i������R�$��$�i�h���d�<�������I;L�D)1�ɬ�R�"d�uIaxB��57P���@.K�!
&��j���	-�MC����d�r*�o���(��D�d�&�X��bЃ=j蹃(;ʒxA"�'%2�'�����*I��x*��\��������@�0�����J"�B�/��m��:�(OP���� =�"-c�iΙ�7��B�6M��M\�����Œ H�l��@���<1dȊ�����	 Z���y��ӂ#��fI:8!�l.(%��E�3lF�i��2'�	]����-7�$ȩ8�h��`�q	ؗ@Ű�X�'MruAРc�����O�ʧ_�r5��?	��8���O�s&xk�Q&�&q
��ڸ(s$Ǝ���T>��|�	$J�\�s�O�
 �J�2$N�@A��%��I#+Yv~���'~�X����qsd��$�P G� ����:���'���f"|�	�\�4ٻ7͜? ���\�2����H��I�B��4�dC"p�R��2�,C`#<�u�	X��"�"��X�W���
�*a�ŭeBb�']��� JO�[��'���'���՟���g�5��^񾑪�%� 2�Ixuo�.BlF�%/ҲY|L�)0�?� lF�N�1Odl�/Νp)�m̈4�4m��l��$iGC�P�R�Qf�����-�n<�yR�\�9���k�Ѐn,�Xh��~¥^��?�V�i `6;����iO�|q ��g��J3��j����!��OF�F�G�q�*}3�AB�[ׄC���n�'#�6��O�˓T*P]�A�i�~�S&ס5�xl��-eUl����'t�'��N��8���'����S���0�A�Ai��Ԯ�REY�<W��� @"�fz�E���Ud}��d<V��`1C@	TGN��`�FG� @�G��d1�Y�'b�����/Kp;��ѰS5y��Z`�>�f��4'�@h��30"O~��ֆ] ɦx���XԸE�'�ў� \Pr��(y�ӄ+I6^=t��?O4}mZ|�Ƀ�4�<�D�|��h/nR�B�-�ru�q���e���2���?1���n@"��&4F936d��Ǡ�H2\?���O�Y܊D pN�0'p��KD:�m7D}�2���j��qcH$ZLj���5�'�"6���䙕"5|���	�pl��$��1���Ԯ��5,X�[#��r�[��Y�y��')�}"�.HT
0�կ�d��rdؚ�0>�B�x§��4�x}�R�ۆ	�4�Q�/�y�i3K�7��O��D�|J�*��?���?�b�ߡr���s�f��h��@8��V'�"��k�������I�(�$�"�L`Ti�&\#źt�0�_� \���ػZ�(�H1�O
��}����;7XJ �b�ޥ8��;$
��F�4�r�%��?�@�|���'�f̹��M�8����ɪ6�ސ!�'�4��o¹1fJ���׼  �@��$�_���t�'�N<���Uغo���%xt�'����-{˾����'���'��Nj���i�Y��IP�V��qG�,�����1x��Má��
lHX��R��1��.$�}2@)���L�E
ԍ6��p��}�"P��,N�T�p2���?�)���?ųV̊>;1On�i��ND	䵊I[l.ms��Ol(J��':l6�Lt��ڟ4��My��/m+��i@E�19�F�[��̵�x��'K�0&�Ž}D��`OM�7��u EK$ғ�����DY�`�poZ�Aτ):t@K/Wg���iK�
Zr���퟈�I˟���������|�e�F�0o�H���T���j�2l"��f+ʁG\Fp��o�;J��^4[�~�<�gkʘG3��h��ֺ(�jqƀϷ7���;Ʃ�j��8���҄Uf�R ��&W�<Iuo�؟���4�d4���WlO�L��@:d�ȓt���j� -$j��h�d�Q���z�'X��P��_� �C�X�\�P�'*�7�+���1Rnhh�O��Z>	iE�G�U��5o�Z8� �� �}(r��I����	b�Y��%��f�,�&�`A�.��hI�D]	�*�R"G7�^�1S�
�|�ؒ��
��<��J���S4P�����,_���h��S$i�Ԣ<��M��,1ܴ����yi�儁n���($��24Z�s66OT��䌜8:z<�0�A<1rmj'C^�*ba|b�,�@q�bM���w���2��XK�d\b�mZן,�	O�4��t\�'e�0���"[�v=bY�A�bG����@QDX�nۀY2���)1�'��� ����8����L�)*�ʈY���#m��AJo��q��`��8�)����-!t��-Ehʼ���R>^��j�e@wv���k�)��ĺ�����4t�u�ʘ*��=��+D��/�i>j��H*rx�#o)���X؊�4� ��D��|�H'�P4^1`��fO7,4�D�O���uBR2CR����O����O\��;�?ͻZ�:䘀��}W��Ȑ�m�n�8���2���Y� 9����G�4���+k,b�Ĺ�-FA�8���ٸJ�bD@uaѦ����!(҆9��bx8� j"�I<>�Nd�3,�*y,L����x���	�c�������I�G����f���C|
ċP��7e��C���̑B̒6Qc�5��$ߋnt�ܘ�J ��HO�i;�O�?�Lm�'"�<R�䅦lF���!�:^x(��I��I�\A&ɟ,�I�|�r��dPnXq�@��@)�Ao�&T�uo��'����<L��<�&V�K�PM�ׇ�/v~j)C��TK<&u�7�;�O�H�q�'�"6�Å'}f���3�dE��"�s�!�ć�{@��H�A˗m�� �S�&R�ax��ɗ,�����g�.YV��Hƅ���2��'�l�aS-`�b���OX�'v���3ĀN�X��K�E��T�%@�
�?a��?�D�B�?�y*��Z��_#N��a�擯R6�}��	�V"�Z&��Y��L2�,
L{�;�L�K�'�L�x��?ё>�Б�J�MH��!�˾���>D�HqVɉ�;�lP2b�S��Pg�0�O�a%��ȁf�0��4(�n�;5D�P
o��b����M���?(�bų�/�O��$�OL��V�A�y�V�(����,��V�Y��T�Kљ��Ѱq/��4�]�E(?N�Tc>��X(Z�vҡ�_�����ޤ���f��*l~P�N�?�N�k2G1m۞��B��wYHEAE j�jT��
	D�Z�B�eTtU��&���Ove�v�<0��(�}�����"O��{��ҽۢ��q(*trZIۢ���O��Dz�O���`Ɇ�:BI�1�]H�/��U"�' T�z�B_�6�"�'��'������݉F��XE|�h	�OD�(�A��A�� ��π��`a��?�[ā>Jh1O~u+�kƦ ����"�]v��t�S�6�&�
���O����a݇~�����b�t���y��2�T�)R���DΖ��/�4�~�jN��?Q��'�(2L؃�z$��Mz)֔��'��2n�&�!��ܧ6���9w�B7n��"=ͧ��-��̂r�� �|����g[�mSƫ��F��IK�Of���O
�d�)���$�OL�Sq�~��33{lD�q�L�rY�ۀ�J��^5x��W�0�{Ģ��:�F ���ɱĖ5 �e��Dj�cY ]�x���J]~A@�=WMD��ԥ�,�r�X3剉73v��I����$�	8��]x�I�v�@��GK-D�4�W��]T�8�ԌF���8�d*OҢ=�`��#l�x�	��>|9[�K��<9��i �'�İ�e�T���O��'=�t�2E�_�2 v*[�tX�A0�	��?���?��!Q�(�A�y*���%���ta�H��<;��	"2~�V��/�*�HS���/�����ܺ���Ղci�W��#P� ��T�'�H@���
�>�:B��P3pொZjN�p��&D��㴇�H�B�	��`��	�"�O��'�P�%�+Bue����.P�驄�`��)��ڡ�Ms���?9.�J(�$��O����O�S�Q3	ҥ��C����ip`�V�Չ�FS�~R�7�[�g�sDb?	Π�|���"r9��ҊVZ�C��\�&ȉ�Ҥ��k�-x�C��X )AY���Z�t�ɂ������w��@�Ќ��m��hw@T�V��
���>���O�t���C�O�|D藃S2ʦp�"O��sDK�1ci�|8��D������O�mGz�O�҃�,,^�6��<d���D�\��'Y�lIe��H�r�'a��'��֝���ݐ(Y
`'�	u��\�V&B�||��"��c��QW��S b��TA�?�Fz���0�⟷/X�f�L�M�����?E����\rD��OAFHDx"��yA�Ê��p.\�e!P��~��?���'��*�(8qL�E#]*K@�Y��'
�Q�"ܦ$r�$���LZQO1��|BI>9'
�
t��u0�x� �;\�
�^"���'��'2MC��'A�:��yka%�<%�@qaC�p9Fh[�/�^P��!�{� ��,�ؙâ"�(O��a�Z~�0�W�NF 9�eVr�d g�!���E��$/�)b ��(O�QB�'?�7�]%i���y7��%x=�kG)\�4!�
1�
�ȕL�/�eQ�E�9b!�D�?)�,�Qo�D 
���tH�D��'���pC��M���?�*�J4��6��ر��ٙU�~���#Sr�N�$�O^��EoQ��U�
�,���(x�4e�K;(�T�Hv�Ba2�����Yz�G�2Q�p��%I2H���"3b��;�$7-	V�d�j�%����F�cu�URB���n�( :��D�-
��(�'�6��%@G�(R�����,!���4?�e��L�K����Q�]��9��yA��+��M�r�]��gS�3�~�̓E��Uk1�i���'��Ӆ�����ڟH��(2?�iv�̖,b ��OLc���d�v��(�$B�� H%Ɓ4��I�|B��ٿ��)�L�Ҙ"�jJ�h��� ��9ڼUS���0�~�)%�ȳ=�B��w�Ͽ#�l�W�A�'*��)P����ς����K���+B}�'����k؄5����x����ܧ&"�'��'�џ�B���):��ơ=���#j�6���*޴Z-���|�O��4�P+�έ� �E����,FE����L�t��&�p�
�낫O�!��.V�<y���b�ڴ	�*W��!�d�+-�qDL��o���HDiP�x�!�D��\��b���"<z�ÈL�!�䎪SOЪK؎Ȓ��h��\�!��X�"���%P�H��(IB��;i�!�d(<���%�]��D����!�D�gs�yZ"h�>4Hȕ�BN5!��8D�=i��ń,и��q랾`�!�d �����܀>�����)i�!�X:b�<+U,sb�@��V�!�$���R5r��T	����f\�!�!�䓑L� ��P5��E�D��X�!�d �2���I&�ժ��xa&/���!򤁲k���t�оb��B5F�;�!�d�: �$���16g[°���2!�DŕS�rY�V#�:Vt�`��q!�D�*���8.�:�|���M��y !�D����×��W�f��-�=�!�dX�A�L(%F_*Dt���J�9f!�d-yZ���c��X=x�(�Hp!��ݸ�U���U2��q����8j!�����ʞ�U�tؠE�Si!��  `8��,�V]p7]K� �"OT �G	�>��l�k�!Z�0qQ"O���"���{�0 '+��[��!a"OT�����.{�  1-GLȹ0"O4x���6u D��T��
 �l��"O�8�4�҆L���;�� ⶌ��"OHh����{
y�&צW�:��"O�8ab�@&C3�[ǎ��w@5�"On�Z�$��
��p����jd�RU"Ox�ځA(s=t1��Y4�Q�"O�I���YÒ��O�^J>�SB�A�yr��.<h�0('@t
������y�n�b
8#$N�� ^�UQ��O�y�&
��9u�6D^T1�)�y"�[�aQ�mM0]`�G���y���c�.u��,ש8�qc7� �y/�%?��2�X���'�y�M� T[N�%i�? 9ځ�����y�T#m�l�sg�4|�Ε������<hΔ����[I@4@Ԯ�z��L�O���U�6)�Ԯ�n�ar�8}n�[I�$B��0�����%�ԙ��=�ɺ#��c��Z9C�`QY�&�(��9��_fk��1����S�>�0O@*kQ%8�Q~L�/��Hs��A�0��#ɔ�p<��[���kl��p@�Ǧ���O�R�(�)��$x��xR�&^<�K��am�|��I=y��'�'L�����>5�`4+�k\�tv�9��nC�},I��{�)�C�'Ilj�ORj��դ\R���ŀG�j�"����Mr.O�DXc�]�]��I�]?�*U�|�'h������<�����ͺ}�P�"�|�ݚ=��Q��F���"5�mw�OrԲ�JM�c���`�"3^�0 Wk-�%9b&��y�V-$���<	�ipޅ{��^4U�U�
a.D+ҩ��(��]"$�&OP���M_�q�M+��֋?�h�鐤�{�']��~���ЏS��X���K������p<Y2j?7.<y��C�o�,�3�k�.���AE�k�0xU� :��?��|bd%�1F/jD�Ĩ�hp�7dĞ~��l!��,Gᄵ��($��i��A(z����'��mıOF�`��X�$���i՟)+z��w�>	���V�`���[�	�,��@�>�$��zԠ��ۚ��0k�!?@���ʎ�z�:����N3�-��$
T?��ȴ|�0}��h}����`�0HX�M��×/&҃IK+�p<��D��5��	[N@)3��
�=�dE}R��"g0,@�-�>���A7���/}�)��ɗ��HV͠?¾����I%Ll%��ؤa���u�š9�Y��'D��ƵW�abe�'��p�I�1� m��BϺ/�
i��]sZ�8JM<1�jC�Hf��s�b�M_T�[�MCAܓ+���i�
_$�� 
�	��<��+�b*���O�aoڸG�v��W�idQ@� T�ɶzh�0@�3}��Ia�����m٤�Ɲ@�8�#%�4��'��ђ�O~�	�B���kc��0�4a��NVr!�Id���\B�6m���V��i�����R\+��@�if���K#��A�mn
�I^?IM?��Of��``˨v�����T'�Ĩza�'#��"Nު���╙(2 ���	�R�>pQ"�]�z���8w+������?q��ݯDrz�'eR�4���٪7?���#q�t͑�	����7IT"�DO5�ug�����b Ɔ�yR> P��D,�콂a��~�&� ׇT%m�0�R ��+�?��2�HU�RE���e��~{&�&��R�X�]/�|3��&�fM��ou������S��c����<F&�oi� p���R$�h�q��~�R��� G�!+A*��Y��xZc���+�-����h'���`r�����"�O��'"����%��=d5B�o��dy2�#Ǔ6wp��� Q�Y^��� ���#��d��ɔ9��8H�-��JU�9{r�O��ɖD�*T�����QZ?���ٍg�j` i�)
��1bcL�H�θr�F�^�Z��s���}@"�8A�M�b�Գ�cŦZ�8p�EhVL�4)�����I͟�bv�Y�`��ҵjC�&�8�"0#3�$D=`Q��x1��W:�����*�B��X�WË�M�ƣ?�O�,hSL�1 8�ȅ�ɓ0P��k�٢vE���P��=�.OklR���M#�ݐ�I<)0NفĮ-꓌�'�ӹQ|dYR����]��p�E�#5��㉆:�u;"�E�V��2pn?2lКB��JP.�
��(D�D���'��Ol��Of���4"PX�ݴi���1�-��K}8	���
��PaN<��U�||���B�}&��t�G�v���0�J b�h����d�H�N���fӜ��$�cl�)��4j���/��Z�f�c�3�БT��?��	��gV��&�9���џ� #<�6��Q�	F[X8!�A;�e�7�xB��\����ɬ �$C�� o�yB��ʇ#��1C"O�a��,3zA�#���y�`�,O�����0V�l�H�咡rX��1I�Ct�!��5]���\��`Di]7v��1�e���C�������G@�[݈x�Ęx�A��r7��f���;Ⱥ8 S녓��'9B�Y6�
&C�LBf>G$ ��{2
�c��M��ޒ	�T1�m�� ~Xc@J�2T�����0a �%q��e+G�+Oa{�Ć9w&B��7)<}+S�ΨH�l�Auo4���z��×r%ay�,z��mbqM;/YNTIuY�y!�$2����aI�a��z��<N!�䕜l�`X��4Gc��˖!�-}�^�'��ؓ%Sz���O>((1P|�]�2��2��qc��'x��Vi 6�,P��&�7e��İ��_b��Q#g�.SV����6�ֲ���F,K��#�%b�fc�D���Ef�� P��w,zM��)���2��L��
Q4z���bf�Z.B���U�)��!�D˙+ � I�wM�5el~� e@ذ\=�� �9WT]Q��)���	�S��ء�[( y�0"�G��A1�	�}�:���r�p% �P�ڥ�K@��� �FBV��zf�8ɧ��o[�Ɠwr�t��N���у$搙L6,�{#cB��� Y¯-h"���=�S�QGLe�e��;Y�:t��_�e�la2%ȥQ�X�k�.,lO&�2f��T��R��@�D���d0z�-#�o)Y���=ѳ���%���!B��f��8�7f	Q�	�-��a�uA~Ҵr̀/!��c�@1�GT6 ���5q��H�B�C>��1Ca0�ܕc�"�9N���hª߄<Y�i�MF����p��f,�Lʗ�'HHA��ʍ(�Nؠ5���dh��邈�8k\��7�=:Cx�H��_��H@��[#N٢�y���=�I��Z�&-�1�5�@�L���Բ
�~,0���j�D���ӕ_1J,����2Z��@MR�(�8\��O��f�|Zc�t���NM����5��_V���'/|O���i͊Y�r����?a�8A7�^�X3�Ͱf����`�Ę�f6���1t��?���[�LʑEۙD�=�d)+�+�t�@ӡ�2fe����\+�'I���\���҇��%tX�c��|ɡL�"��IC����ж��2�a�3b��6��6�| ���ߕ&0�sBdF����~b�>9`��V	�:%���rf)֎_F����'x�$P��/j��(�K�Rur���_"e�L��̂�"{�)"Q/ׁ�~b�%��ӼCV�1N�R����Չ��H���n�Z����D"���(6�\'aJ�e;�i�/M�H���[��~�'˩��g:Q��t���a\A��/	>]�4Z�����'˼�c��	GC�%�ԯO2<��)k�t�T�
2��+$��
H��1+�f���DܻUtaR�=<O�UcBHI)*�t��� ����r�Lf���VD��x�����A��M���?����������y�8u�$�~h<�t'�u�j�Κ�����
��"6�^�mB�[�+�@��]���L>���hA+$Ԣr*�ٴR�����ɆM��� �E�4��Q흚P�t�'�H�m���#�S;PU��IyƊ�Oԅ���#��t8���qe\#{�D����n�&#=�1D\��ɺ6���"tLb�o�|��n�>yT���$H L줰�w��]��Y�@�HcC�'��%��(��yղ����Ia�$�۴t�30�Jr<=�'��� �B�?�	Ѻ˕e 8�x����g~�b�����x�Pt֨E�%�y{��z��A�{!�Cc�i=��&g_���8�s�O�D�{�i��R�G�=�J-�Q'L	l_ލ��,*�O�ai���Z��@�'��M�7d��l�x�%�9���a�'�m�����k� [��W�%6�}�e"��9�Q���u~�Yf�'�r�'s���7KLYZH��BO�4�.!�'��������x��y�l�q�(�"�G&����'����$���"DyaG��E���&��p����1	(`�qrC�v�nP�lgh<Q &U�I�v�k�#� {�H�;�A+E�RT��c��6�"Dy�';PH�9�I˼cH$�$�{��V���0I�J<aX>/2x���ᖴX���WWh��=�棝t	Hx���O7����J�X�I�;3��ڗ�

n븘C��@S��d7s�h!`ڢ�f}yc&��o�R�C�V'Z��!!O�w�B���&p�lt�!A;��<�5�]*GT�a��D��%Q$�v�'���E�$6)P�˖�r� $��B #��DP)��B�=�����^Hh<��6I�N��U�]66��ţD�
(a��ᄡ9a^D�ak��ɧ�S��yǍ�4J�T����)fM��	׺�y�gJY�0l���?"
��W�8���O
��S�,�u�IFL��x3�Ǔh��)��q����*��@1�Xn�����=T�f �Ý�]�xX��,�rx�G�7-�$�eQ�1L�`4!�'A��}ѶB���<iU�^7z�!���1�f ���w�$>u�Ң��.t(�A"%Da�Z̦O� ����N�x֤���:[���v"O�X�Q(@�RRm�᎘�G�*�`�"O}PB�S��́����x�f���"O~H����;T$�zp	ʬ/�>Ā�"O8�XҦ�1o�����
(���)�"O �S��hl�DJ�i��,Ѥ (�"OjX���]-������$�jAZU"O�-���_�>��ȣeEF.7s6�G"O>}j�%N�bgxu�%^�!BL) r"O�m��1Zv�=�%"
-#xj"O������C5 �T#�#r�23"ONI8&��!z�Hi �BD���CU"O�@QVnZ�%��1l��QX�"O��H�	�>z��"���y��` "O�y��^�xLʡ���E���J�"O�IJ�_T�X�EP ���9�"O����z��y%�54p-�3"O�8J�O�1��#��ź/�B"O���t� 5Wd�(snW+K�z�q"O����IL�e��$��-T�ZT"OjP��Ժr{4]���X�_h����"O�`i�.Ȫ<�R��¯��=blhX"O��� �@������>o\
���"O`��'H�;IH��"A�͹g=��rW"O�!���N�3�cU��]τy�"OV��Bwuh�A��J'$��U"O��x���h���*D����i�"O\8sF�K�|��ʒ��$T�tM��"O0<I�	Ń7�Ժ�e�n��yG"Oh�x���(ʹ��!�*9](�I"O��@��?*��)��F��!b�"OxK`ȁu~Uqq&� {�*�*""O����;W<�<[b+�3R�V �"OX|#�D^5Q;�ځ�+^)����"OZ����)%�����0[�D"O$p�3%��r����9]p��ӗ"O^�Xc�G�t�bf]�b[�œ"O:=2�C�nx�Cڎt��r�"O�t9t`��lH�#'Cve��!f"OL��� Ҏw����#\14�V�s�"O9z�/B�$>t�ԅ��N��E"O�y���L�S0�T�E���8�6"O� :�iCO8HM���߷c��i�"OH�"���؈�"A�P����"O&P�`�� �,�y��	"�^���"O�iӶმ{���UNǍ̀�b�"O,0Ag��5w�����(3[�!q#"O��(��D����`U&JSV!��"Oc%ɋs3���N޷XG��"O�m��M�,zL�q�� �X��� �"O����/���1�"'i��H�"O�dy2��=q���D�ϕR��,��"Od���dي-T����ٔ7�v���"O��HP��`� Uk�Sh��"�"OV�5Q�j)��A�)�==�Р��"O,��L��J��&I[Z�6��%"O8q*w琍3������L��<q�3"Ob(�E���4p����$�0-Q@"O�\I!f�Js�}�%,G}s����"O��
0%��'��@sF���Fb�@F"O�Yh��p-7*�2>��"O2Y�M)v(�Ԫ j�/$��:�"Oj]�/�U���F2����"O\����ҜA�v)ǰC�Nts�"O� ����J�aGV�#4
�G�ًT"O��#r
z��5R�6�Q�"O�`@+�aP�wD?;ؚT�2"Od`��Ĕd�XĊ@�T'��Ej�"O���'��}�蛴O`E`���"O�<e����d8sb�C81(�1�"O6%� �n5���5�[8s�%"Of$b� �X��@���&]r "O~�i�!E=j+�l��l�2k?���"O�u�L[�H�p��ꍾ^=6��"O��& Om��7�9U��0�"O��Z���o7JX�+N�U�
l�"O�j�%$7��Q��3a�P�"OXuA�oEX�a '�>L��8��"O�]���>�a���B�� �"OL2r�԰X₵0Ċ�->�0�"O$�{n�:�ʌ��L�;���`"O��M��b�@�n��e%��"O�t§��p�%2u��_<�@$"O*���^�Z��0�wjN!����"OH� ��P{@M3u��#����d"O�qI�(Զ^�^�y6�#_8 �:f"OJ���,P�tA���s*�	!�mx&"O�����Vc�g��\U��"O�ȃ���3I>���&P�U��!3"O�؃�N�\ȜAc�hI%x��%"O����k��a?�,������l����'�!���r�VI"w���%�4�H�!]��{�Z�4�v�2J	> c�l����4Fe���%�p;�N\(A���@��K)E��%��	`�����c̄�r��(���T'4��t��� ���μ]O<�;�E�-A�D�=1�����N@1C��8�CΛ
�X%�ϥ�y�
�h̪]x�'��%ŧ����d-�S�Ox>X[�O�a�0���J�D��(��'�Ьi��H�@Z8�I2.[?Wvq9�5Op��$�zm�%�3*յÌ����L4H?!��=%q��KZ�&E�ԑ�D^ 3,�'3ў�>������fq"<#���)'H�J�n(D�H�a�]7B�*,�!�,�Ա�a&D��I������4��ɝ/
�+��%D�����L(�u3fd��N��*u#D�$c0ɗ=�R�@%���ʙ�G��y���	�|e�g�eB�Y�㝌�y�Ǐ;&Q�����b@���;�y�cȮa3Np�� ɫ�>��WǍ,�y�ҳ3 � ɡ�[팴��Þ%�y�(��H;>�S�m÷K���f���y��؁2=$e��
ݰR1J�:f�A-�y�jJ�a0 2pn�+XsNݰro���y�J2*�QS�I�W�<�B�Ʀ�yr!@�2�`x��Bҟ�����)E�y�#��?K��v�i¬��	%�y�&A:8I�U���P���i�oY?�y��'��=��BH> |�C��+o�$DI�',4=0�S�r8�q���g�00��'T��G;l �!Q.T�u)�hҧ�yr�F�i�QW$��!�Q��$�yb-o�$�B�N����v���yr_$k�*ȺF*^�JcJ1j� ��yr�jPTY uMۀBt�͂"�y2��sD� �S��?��:a([�װ=��{�˃�wW��Ta�2#
����y���	�$�&H��)Sh����y
�  a��K.��J"dD�%b̻"O@h)QcD�!l��x�@1�!"O4�t��c��H �f��M0X���II������<�pX��[	-0�C=D��׆�+�|݂��4^��@��=D�P��$�y$�I��bM�wϴ 
�/>D�xID�f�a���<5�à ;�$%�OT�P���.Ve4-�AC��7��QS��IW�'G��L(抬RU��?�4���hL��yRÅ�3�:ĻD��%/QR�b�J��y�/��:p��FcS���ta��y��߅.�m��\��&� ����yR�>W�@�ĥB���1R���y"'�70ސ9�-�2�@;����yr
��]K��q��+�L$� ��.�y�C��-�X���e����7a\D�!�d,"� A�d��;E@ӛ��TF�T�B�
YՃ�P�6��ր���yR����d&nHN��6����y"$�.�U�Ɠ�G�4�bE��yR��?p�$5���-F�=��=�?a$�'��O?����K1aV��(�$�Kv��vLo��'��
4͗�/j�×_BO�m��4D��eD0W���2ek���1D�=D�	��7}�d���ͥ ����;D��z��͜�J���d�� �)a�;D�|�2�F<d�����	�d�,�eh;D��q�G�*}D��U�Db%|X�R�:�	S����P�Q�
5#-��;����04D�4P�	�?������[�p��D�2D������]%���_T���"D�А�m�9�8HsD�F�bv���k5D�,��&�4e�bX0D��)���`թ7D��Z��B=%�f�C�#�ĉ"L!D���5"�"��#�Όh`�D{�,4D�tR�ژ#�@��L�SpD��`'D��H3�H�vl��#'
-cvX�ITL�� ��I�/�s����u j�"�L�XHB�I���Cƀ�Fè�+�a��BfB��"�~i*M�M�Ȝ)po�yNB����8�s�ڈ甙�R��	
܈ء@h.D��JצM_���&ȑ,�(��+D���#C35� ��*�n�8�DG$�O���':RIs *�<�zABt��06$B��=S6��2 n`r����x0B�ɠ������7A�����2y�C�Ɇ��d,تLc���F����hO>Y��/7$Y�!!�E�@ C�`8D�@Ճ��)B�[�W�8 H,��ȟn�kG��><y����@)��	�"O`eCt�� L=��HK�$�,�u"OƙJ4/'G��(ٴ˝>I)��AB"O:�{wX�{�F쉳ɛ�;&x�"OL�0���T�z@��J9\氹;W�'��I�`t"e��ʆ�E#8�J�M�jB�	�($h��b 5lXR�!�&0�XB�I�@f�+d�V�/*����O-��B�I)��p1�O�fð�{檋�[�B�y�mbI4-��	pc�C�B�4"H
D�e!I�v,�e�I�]��B䉻l�58B�)��A
Cm.��B�I�?UE!dI]�d/�Z���;��C䉐@�*{�lҊc�~%��I��c����hOQ>����Q��L�S�T�*t#D�:D�� ���A)�
M�
Շ�9���U"O��K�B��qt��ځ��o����s"Obi)�a�a�h�5 ۦ#��]�"O,�eFO��t@0#@ިG�	 "Oʭ(q���u�Se�4k�(� �"O��i���v�2w�����с�"O�8ڣ�ݠ[��%ŧƄ}���"OL\�G��(�D�8�e����j1"OB�{���A��Ж%��a�>p��"O�5cc.[�L�P��J<����"O"aS��Y#
��aʃ�?���"OP��J ���pG��6X��S�"O��qM%9*HE�@�T�p Ȕ"OrT�CY����C%���y"O���6(�HJ,�j䥊%,%�r"O��j��K�K}�$1߳�̓B]��ȓn#�i����+.f*�Pa�(K�U�ȓ7[�H(P�ͭ`�R�V-��c�\��ȓV�J��# G�-4��x���z;.8�ȓQ�\]K$�:*SZ��2�vg���ȓz�*,+��ąp��[�#a� ��ȓJ��rf ���9��ȓ]ز�3�d�e�-z�C�1�ȓ&ꮄa��O�UrE��@��Ć�99�Ր� Ɏ�Z9��@T���ȓB��}0`[,�I�f�m=�h�ȓk^ sU�ݜ �5�
�䕆ȓ.D e뗢��5����	D��`�ȓr�*�h�R������Â5A��ȓ4�����ɫ�r���<���ȓe�� x��۴���B��86jP5��wUf�1�HRb@���	3;����ȓk�ݱ��ȸ|$��� ��.nq��?���k6̘�C<D��� ����.�(�$ځX��		'쏌<ME��Q��*֡أX�*�����	s���ȓlU,�q�@�8��Qa�x;^���H�(����]�w�Ll�u�	7T�(���d�Q�S��u[�`x!C@-�Z������ ���Yb��FB�H[^��ȓsv�t(�G�?���I�_����4�.Irwk�fmcE��Y��ȓA���1.ʃG��A+�(�4��̆�
��ks�R�a����L�B,y�ȓu�"�e��cB�X�&U ��R�X�Hr��Eb��P{Ʌȓr��QBd-�<q��q�G���r�b�ȓ84�����'��3��F35ȼu�����J�:vEXA��M�-��i��-�(����d(��O+U����3=X��s�L=^������)LHb%��5��	��\���9�Lڥ,5 Ԅȓ��a���L�?��\)A͕�S�<��#���+� ��!��f�#`���XJѮP'P��dq���@f���ȓ^d��a�*Ζ9�)������~�LURv�Mm}Ve�����ZQ�ȓ�-{�M�.m�~�!3C;{�:��������b��C���ma )��	Of8����� y���#�� &1B�	�	���mG)E^�g�\(0]B�� Kd������Vc�	<q>��ȓ $`d�Û/�f��'�J�m'��ȓ1J��H�R�.�T�91*�k
�P��S�? �-�!�9b�Vt�e���^�{�"OhZ%�ȣj�V`� �H�B���"Ox����Y$U��"�µz����"O���"(3�2-IU�U�F��d�Q"O��	I��K'������M2�c�"O��Js
���H�ڧΞ
%P�;�"O�l��	@���Xf��X;���P"O���5�·/�r�k�,F��T�"O<0�*P�mX�D��jIe�4yV"O�<�wm�MRtT$cL/I�ڝ��"O^܊Pȝ;^�-�@B
/�b��#"Ot�0�*$�6��@�C9_0���U"O����^(E!%��*!�)�G"O��k(Y(Z�����A����I�"O���	�2���r�OTn>�Ļ�"O�p;�	��@�(U.ϰ7(=�C"O�Q�#׷?N���Eh �9$"O�-:�F
�U����ik�X;s"O:��u�E�jpڄ���<R(zP"Olc'J��ugи�q�M�@>��"O>Xk�¨>Lt�̚�+8��h�"O�Ċ��Ol`6$b��6V�y�T"Ov�6�D�1��� ��!�� C"O����䓓3X�9�/��k���7"O�� ��J]��.��/��5�"O\�@�J�;���е-��3�̺g"ȎzDÖ�o��3���d���Jd"O����.#� KB�սx���؃*O��آ�KVn.�P%��Mz�y3�'��l��`�^�������JO�@H�'���b�84A\P� �9P��"�'�d2��KU�d �J�9�<���'����㖥j,mפ�/��<#�'�&@��B�z��%b�H�$��$!�'�����MU]u�E͗��,L�'.�)U(U���*��8����'�H0pdU95>�ࡂ�J���'�꘱B�;8�,���D�y�'��ȳ��U�27$�k��lj���'���Ã���)0�/�!pC��!�'�H�SfkZ�8�fʆ�'2� r�'_��a��޹b�| pL�<S	Z��
�'I:ݪ�o�Z��y�3aL:E�}I�'�F0X�MN� ����SD#Q}���'b���e ��pDy�Ƈ8{;���'dP����]��씀���<rf��Y�'*��#1d�u{��(��uN$Y3�'�|%�*_�d����ᮃ m�ȕ�'ۈ��TdO�a��	A�HJ!�'��̓��:l�4��2�ԀάA��'���VL��Ai��I��' �hc�' �ZT͂D	��r$�n �'x�@��Pgf��Q��Ƨ;x�x��'������-R�2�a�D92W,�+�'�:0�VG�/	+��	DHd���)D��c[1<�(�r�����LѰ.O�yB+Q�wL��D2 ,���9�yb#ܻW�|s�I$x���
�jͪ�y�$B�g6 �i ���kJ�p�'n�:�y2ɟ0�bs�_��X&�܃�y�Ğ�5H���%�Z*D.(G�\��y�b�S��+�͌�r���fe7�yr�ٻK�t�rg�c,i��K0�y��	6�.���kdC���y
� (��%�X��‛�a��*��1�$"OZ�K� W�:��Rp�۫2�Գ�"O��	 �!o����pFN�Y>4�c"O�1��c�/l�H��Ł<|��"O��Jb��92a�G�K�E� 鐂"O�p�B�|f�P�h�	0ʰ{1"O̠�t#�1j��s4)
!r�"mr7"O��cnA�i͞=�����yP ��'"O����cךtln��Ə
�u���"O�!�X/-j �en܍n͔�3�"O�����K>��Ɉ4h�!]����"O�C7�%
p��w�Q���Y�"OX4G��bN��	 �FH��"O��_X�	F'J�^�%+WM>V�!�d��sX�����%y�L�{dM,	!�d�>8�qQ���^���r�o��!�Ȅ?cȉgB�-�~�+.ژ[�!�䃌L�V���I����ߢ�!�F�	*��D�݁O������&x�!���UU�|"�K��<��� $7i!�WE�|�G.�`�E�,o�!��,oʌ[�%̲V����Ε��!�Dș)l�,z�9U��--Y�!��+:o@|���	n�d�2R�R5�!�d�v1��`0�K��\��K��!��Wr4��ʀ/5��,��K�y�!��7rx��BO�k/�ѫe�"'�!�Mo}����$�ޠ�d4p�!�$L.~���&LL�{w@t�6"�,U�!��:��XC�+7�8i�Ǐ�=�!��ոj�N�b���G���9����Py���xhQ�G3z��'�y�?{c�q�6���Aҡ��y�Bդ)�X�Q�"L�'�er�KC�y�̩w6��0e�^H��Y�� ��y��ּH�Ƽ��n�A8�12�iG��y�E�vA��ڇIF�7c2��)��y��Ž3�d�A�|��`��y�[�����ɲ>�Bi��e��yBG\	(������F�@)�%"���y"Ή��Q��t�̢�����y�k)d�V	���:j��P��yR
 �O�� f�Q 2o2�Z4g,�y�g��m>]�5�8'�Vl�cA��yBj�5r����!J%ЬT8d/��y�M�.�F)[��υ(��zB�y��@z��Y�l�7$�$y�I��y���L@x�࢛i�4ܣ�/#�yr�1ca0U����,<�1F-���y�G��pD �fV�o�*���y2r|h0�/y[�m������y��[9¹{ƨ�;w#J��4�]�y�A��y��L [!s�ޥ���G��y�0p�.��D��D������yr���{*�.��Hx���.[(�y���'�����=�4 �C.�y�S$y�dh����/)*�I&ܯ�y����A����y��Qt���y�aW�B�y��0@L�!�� 9�y�i$+y�z0�];#.<�Si��yf��j"`5��ϑj$X ڥ�Q��y2)����p�V fK�t� Ò�y�,�7~���I�M�NS�U�����y2)	.qص�ߙ9ʈ�x0E�"�y
� R5�6G� :�\h�P�F.b�J���"O�E�� �hf��z�g��Cx$A�g"O�d��m×/����)̝0����"Ol��X<"ʓ%�p[z���"Ox8����Y��ł�=F��"O XSS��/5ؼP!���,�y�"O{ъ��~ĐC�>�VL��"OĠ��bĒ�e#p�F�8�T}��"Od A�IY�.QX�u��/jrpXؔ"O�2�̚d\�9i1��	!]��zg"O�a�pdH�N����3!H��1"O��
�O:��"*���v���"Oh8(E0��I��OJ���	!"OF��$Ɛ'b�x��-���NX��"O��@�� �8�T×(�F��'"O���\T M#Ǣ�?�`�+4"O
<X�	�,�X/t���RC�,!!�䅈g���kGH�.<��3EÙ�L=!�d�� ���t��?H�V8VAϒD;!�Fy�z�j� �4T���h��Uh!�d��hhvlBR�LÔa���29�!�D׋R=Qr��ؐa������ݤ1�!�$��IF$�(���?��� ��!�Z�Zm�E��0)�N�q�ņ4)!��� i�F�H&M�0s�<��'��5�!�$H�]'��+�-ͲN:�z��ڴLC!�D �x����Ԩ'�:��D#6@!��b�������!w�I�DCJ;W#!�$\ꩊ���C�&��a�'gd!�ϛ����B�G�y�b��5"]�_!�$���>�`�����̑b�!���S��� �@^�/��#g��		!�$I�>�0����#.�˷&A�[�!�ы#FzS���Y���t��M!�2R�2�1�#I�<C0L��Ns�!�D,Q�Ȉ��Ӆ1"ɰ�+�!��%\i��i�"�R! q�g��O�!�dE)u=��P�mF
��PE\�B�!�D:Z���j���O	���Ճ�0j�!�$�� ��ڡmݺ=���xDW�)�!��@3H>@�(C#��=�)�q M�M�!���j�!�%����䟥N�!�$ز@Ү�z�fԙk��\���3Q�!�dӒF&<0j��F�3�n�r��0�!�ӷi���`��-�Rg�6�!򄐕g6�fiЄM�Р�7�at!�dQ�w,��+S&7� �qa��!�Q�g�l(�g`@�fI6P��oӽ�!�d�������L�Beȍ�W�Q�a�!�DɫjsL���4a�"1�bn�"�!��	�{���K�GY`��D1 `�~�!�䒂x��\��-��l��A�eo�H!�U/~����Ҝ�0j��bT!�DU;T����&aJ�8�9s���$:!���v��a6āWCt��0lV�#N!�V�0"�q���l1�ع��� -!�EJ��DH�e�r�j���t�!��%�P�c�Ե���	�!��F�<�<��0�A���$n!�]):�Ľ�'8�&0��j�4[!��B�� <��L��m�fhƨkM!� ���V��*{d���s��;{Q!�$�%>�h�It����҅�ԪL7!�$�37L��+@.߆H�zy�E�ܣ)!�� R��v��i��-���Ġ3Y�%
�"OB�b���)%���t�R0S��u"O���U�	P=�����?#>E2"O�"�HG��m{�灓O=r��"O��xW��dX�Q��#k0���"O��ZS�דe��@P �A��9�"O(\�E�#S��bN徜BR"O�|pgF�f���/m���"OH�!�+��!��oӿc��p:""O�XkՀP�19Z�kdҝL���5"O"���55�	� �C��91"O��c�$=F$c�[�0�� B"O�xj'��sj B�cZgO�@X�"O�8�Q���O��b "���j�C�"O����I��Ofp� 5+@>v��DZ "O��ٓҵ:��� 1C� nFR "O�uQC��)� �2A�wO��"O$D1̝"āe�'F�L>l�W"O�����<��X�DW�",D3�"Ot�h6�.s���w#���0L��"O�s"��n�����P�u�����"OZuZf�߆D�(���h��7դ%�R"Oޝ��#S�^�6pC�þS�@t�u"Oʅ� F�n������.�� "O>QH��Ԃg�;di�	E|pa��"O,A�M� F`�HW��	�^II�"O�xB��lB����jKjYZ�"O�8�b�''a
�XPh��!�Y��"O�-�Vԙ+���Sn�w�	��"Ob���(' ���lOM��[0"O��+������I�d["$��H��"O�m��] tȵ�ӣ1vD�4�"OҴ�'H�In�Q0�؏7p�0"O4�a�DS�������T�A�A:D�������:� ����!�rZ:D���GAQ�q�R��͞�V$n�s2+D�k�["<�)�G�ݨXkR�2&�'D��g���?=: �b�Z�$��[W�$D�@�r�F�@�l�IY�xJv�s,!D���ԊOO�J�A�m��BgdE32D��
��EP�l{'�$Z@�
� +D� �1cnHj&�%	�HS�*O�IQ�0p?����ui*}�"O�-����*B���F R�V��)�"O�p���!/N@��N&I��� "OĈX�I�T=s)U<p�8���"Oj!+ţV�T�����~b��w"O��H�@�5Q�]���ÅP��"O�D ���qP2T!�j��r����"O���ƻxR�@��鞔��"OV(#@-a�@�{����R���"OY�B	�X�B�⧪��N��p�"O\���M��DY:dg�03����"O �i`�I:�T�s6�ĳ!fr�Ҷ"O�����%xվ�a���5�LX�q"O&d�o�*<x�|R�չ��e��"O�YE
�1 �x��Dx�d��"O��z�;2��(S3B.VY  ��"O:ԚE
%�P�*�ƂKg��Y0"O�|���+����%�O�]�6"O� h.��ͪ��U�H�ҨHp"O�+QA�GQ��K3��(Q��I�%"OF�[G�Y�QG�uDXK�"O�����P�� cJ��Um|���"O� @�Ԧ�Yo���N@�x98X�0"Ol���%� Y"A��jsQ�]ku"O:U锌��j
A#�I��T����4"OJQ+4�A�V�I' ����"O6��-�%M��� &�6YJ��u"O��`LJ�W��+peXjL�\�T"O�=���X�H�`)��K�][b:�"OL���%[W
"���◖iG��3�"O4��f���6�"��,&�p"O%h�Aĩ@@Tm��a7xǄ9C�'���0�Ǵ.��Y�ES�Z�<���'�%[��c��QA�J�T)r8��'��ۤ 0.�H0�#ݴt~&��'��ᒤ�BU�Xi �`l����',Z���H����Y ߓn�dq��'�ha���C�&xX��FZ�����'k|Y�2�T4d�����˂Z��0(�'ȀP�(�>&D�dߋ)�r`��'(l&� �n�(l��\9�L��'ֆ�AW��3$��W�10h�+�l D�X���auNQ BE�K2:q��E?D��9�jW�.�y򣂂)}�0�4�>D� ��d�#0���q��7*YX�3e"D�`ّ �����Gb�'vNf}з�*D�����f>�괄�y!`�&+D���r�V�a�X|�\7+M,jwD)D�h�$��e�*(�Z+��*D��V"�&_%rl#����3�:����'D�,Y�T���U��&�x�Lq�f'D��1Pc�E������&}� ��#D�xW�՞_s�=s )ʏ��Q4�!D�s���1t��b4Ǆ+d�z��#>D�T�"�se����?����.D�d8�P/��3������y�k,D��3�m�5�J�1����@���A��/D��@p����U���4�Hqb'!#D�p&�X�H�ā"գ&��<�p�&D� ���A/h���q5jZ��:��?D��f�9;@�V��xq�=D����_�:��ă	ߑ?zl�[S�<D�T���Z�(�\�{C�;;�D��-8D�<�dO'ӪARr#�<OĄq��6D�,�����|�&��#?�� �!�4D���ꞸcHx�).%*��y��4D�d���ñ8�9a�'C�PV  E�/D�Dɧǔ���6�A�R�|ђ�M�W�<�F�@�
��%��h�z�D%��,�}�<)rn�/j"Pɲ���2����7FA�<���#)��E(�G[�\�~�"��g�<��ıOfVr�ψ�Pq��O	c�<af�U�5-H(�F��D�\9�5��[�<qN@(q�|��aE�{��	r�^�<�
>xaʜ�6ʍB�L��$X�<q1�o�� ����]c��b��QW�<��̅(8.�t2m��6�v���)�Z�<9׀��n�d��` �w>T���p�<Av�-֔��E�Ɛ�!V,Za�<I1K�/(Q�Ē�s�H��ek
`�<ه�N}��eʍ�Aݴ�z%�Y�<)�Ǘ�Vh�u�p�Q&���zPBK�<a7�H;��DÖ0u.%Pd�B�<&G�ip$��0`�����}�<���iIhp2�-x���y�<��쀊&������(p8ؐ�7n�~�<� bm�r#�58C�M3T�͌F��t["O�9 7J�8x�z��A�[�{$��'"O���i� Lv]X��(�:�"OJ�I��ā<T����Ұ5��%��"O��k�",���ag�G y�(���"O<W��& ��Q�|����"O"� 0�d-"��U��4��!��"On�1�J�l� �k��!�.Y"OP��J�'[�\ՈHM2Q��1{E"O^Uz�ؙb�`*��4?&� �"O�|�2j�z@�6�P�j��Ɇ�
A�<i4ȓ�}���(��g���� �F�<�b�K�t@F��Zܘ��A{�<�3"�<��b�!�S2 P�sc�Q�<�A��>6��aKQ�0Cș�%��O�<��M�FcݻI�1e����R�<��+��}�iAlW@��P�O�<!�d�y�*\��0�B���S�<�@ݥw��!S����E�ε���Ce�<��a��{y�dZ%	D54����K[�<AĎ�!P�2�;3�ȼP�"�ڂ��Z�<����k6��X��Ue@^hR��p�<!A��-zP�a���� ਖ਼l�<ᵧZ:Qj�K���-G�̀���h�<��e�w��&���F����Q��e�<��dCF��&��(W�re���{�<!A�(0��3�d�q4��s�<�W�$l���`o�J����$Qs�<�����V�@��߇>( pðnUk�<��΂� v4mȀuϾ�2G�߱�y��T Z�h\�皌<�J ��H�.�y�1b��葥݂0>|31aR��Py�,�7-��8��IL*��XGbE`�<	� ����u�\lg2�t�C�<A��|��A� ^���h
C�<��m��p�2�!�����!MY�<a1l���.���J�
�r	*W�J�<1F�
%V�AɔG�� �̡s�HG�<�t��\~�T�blP9��PA���M�<��O��H��k��R~�A�(WK�<9��d
h�Ѯ��Y�F�0�#�[�<��L�0r�f�Z�bؓG�H��E�YS�<q��Β xB��6B�|��Ȃ�Ay�<�4-ًu���#��9x�I��l�<q�
]>Kf9$EM�Y��:�ŐQ�<�#�ʏ( �2�@ŜK�6!B��K�<���ُ�P�r�N��,}h%SpnQH�<��fc�a�`�Q,7 tm�բU]�<醭�/~�Р��P�P�!�M�]�<9G̸j���C��4-~����N�<�A�f���B�Y19�h|�ǫ�E�<	���m��#m*E��p�7)G�<��ƌ�K1-�C%S{r�Q͈~�<A�V�(y%��k�	�����w�<9WGH�䆡����a����L�t�<A��Ť(r'I˄|,d!���Eq�<�@�ُPl�0s 	��2Ԇ���+y�<��f�%<�Ty�i� %@ɢćCw�<���ǯ)��x�f#��
�*��em�\�<���̛\{��)d�� sn�A( X�<��J�sܲX�v�D3 ��3��Z�<�F!�52=�*�+fLB�<a�i�0ѐ�!�L�x���2�|�<�s҄hݶ�A3���LX��@t��w�<� �"r�A�d�Ti�K�*�\��"OV���	̥I�\�j���}��9�"OJ�r�Ԉ#���rCM�lt��"O��1��0��D��Խ7��ɣ"O��zpśo�0pg!=�ܓ�"O�8����
�+7�^1o�"�""O�p�3��~���(��'�V5x�"O�Y�o�1;��r��I�0X��"OF�����^�hA�k{���G�m!�$'+���`T��A�+��!��X�A��c�䄟o��qۖ����!��&@�B͠�$AB�^�PgF~�!�$�aE� �1F
�(��J>$�!�D���SW$�9G���e1!�!�D� zⲤ�Um�u�2��C+{!�$��-��M��@��Z��`H�!�D_�9��$32k�Fv=�ffԦkn!��T�B/�r�7Jt|��q/{<!�$I0H&L��j�vT�7 ��P!����]H�%��@�U��C��. -!�dM"C���T�ݡBd���uKͼw!�䂉��-s��P%4R������/!�G!�~�[����u>|�K5K� !�!��P$b��y��d>v0���]�!��5��D��	 	��瓺V���ZA�%���blb8��+ϳK� ��Dj(U`�\��(OB(8�* �ȓ�V�S���cH���ě'�8�ȓ�ZyYfF�p���d�]�C��)���P�@^	G8�F�X�40Ԕ'ў�Dx�j� c�`A�F��6Eh ��*�=�y�/� 4�,�CP$!,���"'�(�yR�5mk��q ��&����q���y�"©r���5-Ͱ��4P��J?�y���o.���4�U�ߎ1��4�y�lW�}�|�KW�
>i��rf釶�y��/��y9e��W�B�S�ň�?Q���?�N>a��$�*� �a';���TBI?`�!�}Z��FK�<P:yc��Rl!�+�2�	�294��+���M!����������R. I�ա��}!�M�� �G�I"z��r��9�Py���E���3�;
z�Pq@.N��yr�Õi��@vJXL�0�:�Z����O���ĘW�z�"�c�t4T��"a�!�$˂1����Gn7��I��B�f�!�FJ��h%E?5�@ �Z�~y!�ҍ3�E��⎷��q�����,�!�҇7;�y�X<@F��5
P�3�!�d�Vz�%�4�.i�!��"�	W�!�;D�bi�B%��5�X P
� d/�O��d�p".�@� O#T芗��;s�!�d��Tb�y	fގ7��٧�?�!��N)��B�K��;���k�An!�$�����{�	�zˆ]�V�\�nk!��v����d��5�����LC�.X!�d�Bc�+G��]�6�p0�1V�}b�'-�d�na���-#m����t�ݷI�O ��-ڧ�?IR�ڵc��<�PiK�p(�ԫ��y��M�Vu���`��x�"U!Ɏ��y�$�-z<��)Ľ"b�yCk��y"�A������!@��T�2)+�yr���NK`����K�����R[��y�b�fԚ��˽���U+ۓ�y
� ��2�L�6B���`]/d�Ƅ�O��Za����-�&*��7��=pdN D��h�K�$�n����A6$�����E�<a��Q>Ŕ'��)�� ��u�1�Y�e�I�ƃL��!��:2�zm�g`����A��!򄇀,�ʄ�FJ�P�&�����}f!��<FD�#$��xtŃǁQ�;�!�D'S/䙋�M8o�Q8p텡l��'��'��͈E��4NI�x���9	�0�'~,�9��H1>@����$��QI
�'�-RG�I�K�d���' �(%z	�'�1��E?,B=  ��ܜ��'*,D�S��]�1���粌 �'9PQh��H�VU�e��5O�����'h����WY�j��e�˲uE8�*O2˓����'�(�YR��[a�� �ɋ&Ȝ��"Ov�;��U?��@�m�.df��9W���'&�O���	&# &�	S!3��C���ui!���\L�b6��6�n� �@ :!��̗@p�i�p�\�@�x�J.Y6!�7e�tbV�A�>y�Yi��К_�!�A�͉P�I�2m<-�G䝻\��O^���31��B�7bN�y�� ��N�!򤋻伄��$�{f������x�!�d�7+A�P�MŔ;�:��� ��p=!�_-��qy�-L�t8���,a�!�$7h	�{���?{ ~ݒ��Z8.!�H k�j���m[( �8㏓!��σ���@PH� +�pTK`[� -!�dRe!���e�q�Fe*�)��\�!��n�\�gK$9!j�Bto*�	Oy2[� �Og��|�����a��*M���e�A�<q�ɛ"J� ��I>X�()�Gi@�<�f�K�$l���φ$�~x*��@t�<)���,�`�p��E�U��!�w��e�<!�)ʳp-��X#�\�@�`q����_�<I%��T5`Di�ˇ�^lq��fX�<	P��C��5zƂ�+2�~ؚE�Z�<�&hQ+fW����)o��@ڃ�V�<I4o�"� ���@�-p�p�j`��M�<�Q&M�h���8�BT 9T���ZG�<Y��	.r\ �cR�GY�@��͞}�<iT"�:8�ȵ� �R|ذ�k�yy�{�'�������`���q��&o�p{�'{(��(C�Ht����%;��2P�l�'r�Ꟍ�1$R�o��\q�b�-*.�� Y�<)�� \�\X���+6���V�<a�j\��\��	�Xo��)��V�<1 g�:NRV|b�fC�`P�P�Q�<�q	�Q�t ��7�=��K��?��ԟx0�$�&u�N�j�K13�r��%"O(��qnN-%��J!B�u�9�"OX��
%]��1h9�и	`"O���IK?.�B�P'�!�PX�"O�RwғW�p���н-����"O�J`G?��i�r��2NȜ�`"O��ׅ/Jd�!��>��9��"OT-�b��v��[g��2Tp<"�"OJ�4���Ɣܹ��5PO2��V^�(�'�Ig�'��D��30sxآH��Ԙ1��y�*%̴�+M%SL�Z�υ�yb�B"JFd����eP`��޼�y�JW*1�qX�LL-1{�������>�Oj0WK	�H�ia#�-A$l�p����O�}Γ�� ��ВKW�rF
��Qb\=1��r "OJ��Q#Q�n���s�Ⅰ��'b*�-��U㘯XX�����փF�!�$�(̀ Ԥ�;9b�p8��0K�!��&1�4�	�X�[Z��G�̦H^!�d'&��-EN��9
q�PA!��������d`9��-Z<U%!�䛣%�� �8<���+���>!�dXj=z�#N@�ĉ��Kmd!�dI��0`Z��0� ��,�
]!���g�n(��P#Q��P����)V!���w���3d�؎;��8�ɂ�,I!�A�@�Jp�&��>vƱa�'P+�{��$]0N��K$��Cq�pk�I P(!�L�;��SN."WN���W0!���0{)�*�]v70�`$+�!�߳!��(�Ӈ���D� ��
&H�!��ߎe&:<:f邍1�2������='!�$��\�����ͤ
V�-�@nP<	6!�ًYG4@�`�!�u�v���!��Iv,I�#�9v�����2J�!�䀕d�~q@�9nlHr�ݷs!���:3)pm��% Pmp�C6J[�9�!�C?-ֱS�$X/7�ؼ��	&�!���(�*��늞	m��5�RS�!�$��v���g�
1�~��)��!�	�Hr� w�6r�vţQȋ��!��ɠ-PH1��>���*و q���hO�#<9�#�a��I�M"�,�p���R�<y��ӈ�̩B�Ѱ&��1�Te�<)���Z�9������ 	b�<����i�}b��*ĩ���u�<�P ��Xp��h٢?7��+�H�<A��.^�q�E�8@x�Qr��B�'���E`�	��@��rc������p�4�nX0=8�3
)1 ��dl*D� 2a�V2��r&CE�lK�i0h'D�<�P�H7d�"�H�4�Yr�*D��a�.-�Nis4b��]�4 0O+D��Zrß�_���`D4�8i
�M*D�|�����Cä��6f�8��Iz��,��0|2�F�9F��J�"
�3� �W)�[h<qc� <g��E/T:q�ؑ���y�G�F����^�i�8�y�gQ��y��ԝMA��cQ�x~�����&�yr��¨�C�4oL4�Cj�#�y�"�F�N=0��	?v��A�iS�y��:h����F1g�>�)�D��y≒�J�p��Zefb�y�D�%��x��B5+��� @c� �nģ��N$4!��_7h�b�OWt�j�1f��a�!�� �Uv`Z��ԅ9����!֐w�!�D.m^���G�~:H���W3!��=��\BGʎ,hj髐OV=`!򤆈6�Έ��.�26Aj�{�m̓WR!��՝����6�C�HZ�l��	7�!�D��#U�/@G�i��%f���x�d�Z/~�(Ё�oz )R�U��y�԰i]@���J8�0Q�ߣ�yM�Vf��
���H��!�ŗ�y���3Wqd5�a��9y�L���(�y�&�����.,>NMBb��y��H� ����C9}񡢏'�y2��\mP�j'��pj&d��y
� ��0 ϭh�
1�t>D��<@�"O�q��Ɂ?��%	q`���1��"O`��	�8dI�����vtԪ�"Oހ27�ڈ}����X�/a��p"O��a�l���#kP�eI��W�<I#���6@7KY#-� i�a^]�<!�B��	 L:�h�$n8�ؔ˔A�<�Os�4�&m�4oYʴ0q�Nz�<At��Q��\��/�G|X�S�+�M�<����.\`��cƇu��D�K�<Y��8�j�h�6}얰bt%�B�<)��Yp����J��ᘵ�Kj�<�3�T&�n�"l==K�,���b�<Y�,�?#sܑψ�`C���Շ�F�<�g]� �6�S�/L�H����
z�<!�#W�;GZ����ʝ<v����jE��X`��g�� �f-%,4���J>N!"���([���4��-?�i�ȓl7�daq�e<̀�,ԅP�����I0�9��R<=s�(Af�'�N�����A��)��A�LM��� f���ȓ\z�@)\���,A�<Ɂ� >D��J��{��4�@9�6qx��?D�d�f��
��ҫN���f�ӺrL�B�"Me�y�区��	B!�+3K�B��M3V������c��T$�B�ɜ��Aѕ��?K�-z�e.2��C�	�F�*���Oؾt��Mp��O2?�C�	:1�l9yQ��]6�@2Ɏ
$,B��>+T��@B�X$���W�H`�B䉢���l�<���0'Ñ>\��B�� V)��ؓ��.��):�L}ʲB�� I��JŊ�6J���dA�"<6�B䉹2�4SqJ_	��2&�ulB�ɪYW
�
Y�O:�e�����e�C�I�]�R��R���CQ��dk܆ �"C�I�4j�	 �g�2}1�ݽQ�B�	p:��m\����{"��B�B�	���
V��KW^i��C�>�B�OD�A�=6]4�BbBV%{�tB�ɲ,�.���kϚA���g���5�\B�əH%�4hPY����NW�8B䉏+/!q���1[���kQ�љelB䉉ꢹZ��4Hn�g���8�:B�ɲB�VP�FF�O6�A���#B��/C�Z4���ˮ=x�����*#��C䉞Mg����aR ��\õ(�0[C��;�$��N��"N�u�G�*_�C�ɿT���`��w��ct�K"-CC�7b�aed�+$l�A��'�@6B�	n��X��EN<�!���& �C�I��y
�L��3����&  FCC��8)��H�Oќe3����a��8��B䉩!��@�B�Y0?v4S�K&*ohC�	SwZ}@EKږ3�t�X��!9�C䉚8~|�����8�tȆ+m@B�|n�QKG$8�2�9$�D?Q>B�ɴu��ɸ���)$����b Ua
B�A�4�+Df<7�:�Cd�C�,�B�;LW�0q�����z	����
@nB�I��ҹ٠nY�����+��rB�	
M�����I�RX�ЅH(PB�	�S\�MI�bî��bP&svhŅ�F-��1Vx�p ��s$�8��S�? ��Q$��tzؘ��*D�"���"Op����*/�d9��/z�i�@"O~ �� ����6���_��|ڂ"OҔ:5K��%�Ñw5�ٺl,�ybM׌gdi{P�'l�b��yb�>4�;�˔�9
��Ɋ��y�IS
["��dY�D��x'$�<�y�Gճ*���[p�7RFU�N\��y�E2bX�(Z5���Kf8UPԈ��y�I̙x�fe�bB	�x�.��0��9�y�c�O6J���%՟mn�S3M��y�a�4f�c�O�M$�BS"T=�y�܀;<���'��y\���4�y�d |�j���U;|�����O��y�G9$�LPh��5y\Ԉ��V��y�A������Y�w̼,�5gز�yR���`��0hl0�z%o\��y�*Űq��)��^�I�~�d���y��)Ly5�0M�Y�����\��y�H�VFܕA�!R;>�^A ���0�yBjM�0�40��<a�-�E��y���`dC��	 Kȵ��h���y����+�a�0���{p=9���y�iB%r����*�.z��H �Ӿ�yBA�j��EZv�ϋ^�ҝP㋛�y��b=�pc��4�ψ��ybͯc�J�с!��}p*�:��
.�yrA���j8�)'}@�zt���yBJظs����f.X�w��Ȑ�&Q��yR'Q�3	<��d�]�Y�J��@�y���V�yXWa
�R�n��ME �yҁ�e#����F/$Hje)�y"���H ��
�s�T�냋���yb��'�B�B
i�A �@Q �y���?���j2�[�eB�`�Q�y2F�N&b���)�[q r�?�y�&�RKlT;Wˈ7Q�*	e�]=�y�JhM�4�F��� S>T�4���yr,�2 ̔|�`� C� �1%���y��8J@�1g4=�b�z�GD5�y(Ze~L\Xׇ-$MvE
�CO��y��N�i��x��G��ε!���y�+��p�p���Y30t�[㡑��yҦCu��Š��3M�<rB �y�ʒ�z
x٘壒��j(�$��y"M̗A��� �
��1EG��y��D�kӎp撆
�~�[W���yr�'�\=j�J�h`�(�N��yR�ɼ[��I�d���A�Vm��yf�@x:ۡ�W�i��}�gd���yr��T��ᨕ�C�1]�vd��y��O#4"�$���/'�ĕ&e��yB"U�%�i�j�Lش��#�yrC���@�DfB��R�A/��ybꗩ�A�7��
1�ru-�y"��&"��ab�"AL�:E��yBL=��1��/�a 2�M��yٰFb*��S�;&%�|�����y�*͐u��l�I��eh6H΍�y�F��Tl�T�B�ԎUT�YT!�y�*U���TE��Fa(ҫ��yR��-�d-h6�ưG$��BA�T8�y��j��i��I
(tc�-��Ǜ��y��Mh�$��D3��A;s�K��y
� (�!���*���C ar	��"O�1�Q���+��p�!%�3@eN�1�"O� ��Ñ(md�q��c`�"O~�`�&o�P�a�w^�1c�"O��H�4�]�� �'OK����"O������-���������"O �s�d֘k�\�b0L_#��%x�"O�� �l�}��	��K��� �2"OD<�f���% �6U�ȳ�y�!J��ؒEҭ|�|E8�ŀ��y�n��a�B� #A��G���A�ѯ�yBF��{\�dh�g�q�0�B���yשG���vH�&o�BQ���ӿ�y"a�����7GL7%�qȐ�y��]�yZj�{�Ã.g�48%�В�y��T�S�$�*/E�d�q�OB1�y�S�VЂ� 7@
E+�u��+���y����V�"�ᅁS?�lRoR��yRm�z<:`�0A8�u�ٟ�yrO'5,9�",�_�$�0̜��yb%�> �{ԌN<Z��e�0��y��ŀ^�9kEc�e�| Ѳ��0�yR,ܿx�0P�3J�L�".��y�-xu�0a�+��I��9r���y��Z<s/�l��4<:��@���y��>U���A9;Ǻ��W�;�y2�4wi�* �լ;!�)���8�y�g(8ɢ��'!N%33�[�� ��y��y�܄�`%��yjva�bA��y�i� �8۷DY�raTM;�`���y�C��p0d�pn�iY%� �y2FʬV(� �sb
?Y��`�ɏ�y��DJrH��PQv8(�����ybH��3���b@޷Wb |��"���y��ľK�xa!� #S"�J��#�y�I�|?NLb2�M�lD�90��y""X/	�F�����zd��T�y����(�R�`�7m�֡9��� �y�(9��cu�U�j���o��yB&�`8-A��/m�Z"L݌�y"�3h��C�~<4`)�Β�y��P�4H�S�L��'S.�@V Z;�y��B#��]zd*T�O���e�
��y��~�r�J��פ;� @�B�:�yr���2h �@�2D��(�B��5�y�JS�����f�#>�(l����y��ĘX~��{�	F�9���b��yr�5�
�t��C��-jTh��y���r�Y�aJ�1��Y1���yr���;���!	5n�=�rF��y")��m�����_���1�熓�y��QNdC6�_Ԓ�����y�C�mihh#�����狊�y"AܼY1.�3�� ��<�����y�g�\)*4�7eIrI9�n��yr��.ɠ�p0*ΣbJέ�c!,�yb���U��I�6C&]��:T���y��%bdҠ3��0[��,U*Q�y���@�p�̂�@�~1�Eˍ�y�I��9��$��L�N�4� 5g�y���Q��������Mr��Q3��y�"0�l=; h�	4D8�%bN�yr�S�*�x!����%*�ʈ�6F֨�yr���!�1�թB$�f�&�]��y
� �0(F@9l�$a��A�z����E"OV�5��7�Z�E�I7b�����"O,�j�H� N��y���WjL��3�"O�ms텮2P��"�A�Q�����"O���D�\�`�S��":�PxJ�"O�E^@ˠ�c�R& ����a"O���WI�?{�"x�ʢ!ϪEK�"O�,���\�"�n�C�5
f4�D"O
U`f�N�H@���	/<\�D��"O� g�ȇu�z�p���~M�a��"OZ}�p�+aF¼�7V�LxH:F"O�x�v��^'n��A�N�!xh�"O��q�Jƞj��q@��������"O��Y&��>c�bh�����L���"O��*t���rp�5nLo�N<��"O*���2y��G�'&iM[�"O�!ۖ�D�bd���=YF�b"O]��g#�\A��[�����"O�mNL���W$�"W}��J�"OL`Z�%�ETFdX��I:��3�"O��B���;x���dd�H#蹺b"O�@aACĲ->�ȋ���D���$"OF	3�Ip���DH?{���b"O�U�Ǫ�#e��b�`�8��a"O 03�D��&m���7`�&���"O݈�%	#-�t���$��
���"Onm�ՊZ�Z� 0 Ċ��h�"OnDq��]��4�:&�D/�ލ`"Oxq���Q�L+$��2᝭A}��!t"O�x� �f�$�Z'���N\��"OވU&ۉM^!B��Tg�=�f"O6���d �$[���D�a	��"O�zv.V�9�����\���y4"Odd�gN̘ l�=�@R�.�@Z5"O�MѰ/�[��i
�M}�љ�"Oz�����^d*��h�#f�4Z5"O�U�T��UH`�x�B .�8h`1"O ���	2+��o�:1J8iA"O�$�.B(���3�.�(Ib�S�"O���5)X<S�P�P�ƮgH�i(�"O��I�&Z�:~�:T���,̤ ��"O���W��zF���T<�.ܒu"O($�Ռ�e�\KqC�=�`�"O����e�Y`S�O�r�:i# "O�dj�j�/08�h�	i��1�g"O.�T�\��Hd��/:|i���"O��C*�!8 ��`��h1�	y�"O&Ȓ���Y`����F�Z �$��"O���HY0�d����_��8�`"O|@j(@<TĂuS��i�P{�"O�!Z��x,b��g .{a�Jd"O>�CDd�T-�AZC͒5G��u"O�akD�ݐv� h��m�^ ��g"O>\��d��e��EM�5��"O8́��݋���[���DB�"Oʅ��៺J��Ա�Q�g��x"O�P�(^ I��2�G��#r�DCE"O�];���>*7�I��Ө"a
T�#"Or5[��m��e{��/5q��� "O�V���ܡBSD�j�*	�!��}�R�	�`��dC����H�.�!��g���+3��7(jݢ��1W�!���<vl��Y%�L�m�}�͍��!�˞ps��F�E�&IT�@�L��M�!�� *��L��KL����cR9�0�"O�ht�ı@`�c2!�"�x�"O9�w"�k�t!� ��.��c"O�y#��.KL���	�<j��1��'61O�I!A�[�
*��&!�.WA��
O�6Ңr^J����v���κL�!�D�
IQ���_�)���x��>Jx!�^�y�X8i�#Ë`B�+!PCH!��&�=�g���Ks���¡��FB!�dJ�
�������sKLQ��]�\!�d<r�FQ8r�>4$��Щ]�<%!�d�5�(a2h28�Kq�ɵ4	!�Ċd/����Ǌ*����3P!�D�?��h�A�)�$�D��!�Đ�7�����R;j�,@���ԚC!�F$�йY���n@Hp��D(!���H��	ダ7خX"�]#!�ބV��������d�� g�*!��ƽTX$$��I)j�}�C ��!�$�:HAV��:�Z�ڐ��j�!�DH�d@BT9�/1�	�jZ�1�!��B�t�1��S�[��/�d�j	�'��f� ¢#��;׎<a�'g|\�q�Ӏ�� {r,�/]�"OpP�����<�����N�(J���U"O`��"R�N��Sć�k����"Oͻ�lS���X�4�;���c"O��
�;��u�\�r�p+`"OΔi,�h������I�;�J��%"O�x��E���tb����'"O�	�%��x��X�CdxJ�"O�Mp�*�.Z��X9��Z��$�W"O��y	ć%x�\p�ZT3F�C�"OP�ԉ�<:j$�`�e)�i��"OF�y�Ɩ�C�:@��)�>X(VHT"O��`� �0�@�P�i��L�"�"O|,��
Z+'�|�2iE	J���"O��QBuD�P�Ƒb��H��"Oly��ܶ<yh$�g	�Q�̤��"OZ�2Bg�3��32�ʬ:���B"O���W,F	�@�ALu~=K�"Op�a����1�  $g�X�"Ot\Y�U������l���"O���S�M��Z��<q�P�{�"O���]:w��<3�-]�Pd"O"��d%�e��T*R�@�a��!��x��'E
t��mB�u׶DA���7<��u��'��+1�QT�B����6�=
�'_�9�E�%F�x�{�X'0O���'�B�Bǭ6i�}s�i�9x��T�<�OP�D4`����S�$@x�A�<e��-�我TC��\Ы�B�}�<!�C��'�6$Q�L���2ȳ���y�<��� i��R!����I\�<	%.W�02 ��ğ@8�T�&�a�<W��6T)k"o�'vy���H�<�Ԇ
"�@ҠA�&���F}�<Y�	P�{�\E9�'ڋcl@�KAE�z�<)�og�,P��.) �S�˄l�<!3
��
�䡳rE֟	1� /n�<9C�[5dT){q�ϛ`p��@���@�<A%�:�~a�D��J!\X�I}�<)���)�l�k'���G����i�n�<!��޴�4\ ��ðg8����j�<� Z|C��8�PQ�A%ʝY|U[P"O6ѳAa[�"$�&Q
S"O���6�ȮH0�W�2����x��'J�!�d]�C�f����6�C�'܌��N�'����<S�4c�'��Pj�*�/��Q�"�"}� (��'�����ԑ%fUkr
"x���'Sd�e,���D�h��p��m�'_\h��ƔB�,5�#Q�{s:*�'x�\����6�6 K�c@�a���
�'���Bt
��'�8Y�EC�WJZ�s	�'��LhiU���tS�I���A�	�'�@5 c�� !�<C��� v��=�	�'�4�k�@�0צщ���/Y��
�'�-cdj�a& ��D�W�X
�'��]� n+S��ͳ���M�}��'ra�����=�L��UmRD{J��'�z9X��8t�)���4�Px��'0�� ʌO��@K��Ĺu���3�'�����I�rM dj��
a��
�'c�� �� �R�p��+��`J	�'l�  0��_%Z��6e�4x�Lq(�'�,���lۮF�.\�VEJ�z�lxK�'{~�c�d�*'D.�i��@�&ȭ��'Zp�1�HM���D�#��g��i��'�N�r��ob�!Ⲧ֫	_D- �'��lX��˜kV��c�Y6�-��'�P�d*C�]�!�E��H�*�'+��Rfi
�m� DZ�e�,z�Dz�'��!رm��Np
&MX8Z���'M~ps�I5
s ��5헱W ԍ��'<L����b�"��j��$�(�'t�s�-��+Ĥ %�0ځ��'0P���@�0�{���;�����H�6�x	p�ߛ�n��"6D���Ŭ$7��!�P��F�y�('D���4#	�"y��sd�9^J	��9D�0��"	���*�FٖTn18�I+D��0#�=)�>���*T�Nv���b(D���F��:kB��ܬXE
��G@�J�<��kT��y�O�
"q��s�LI�<�GI����({F"�q<H�cw"�G�<�d�F�Q��fo�^!�b�H�<�Bg۹++������;�t ��E�<��Z�9<�u��
R�y�����CA�<�F�� �$p��R&<�Hc���|�<	���v��&�ù���Bg�L�<i���H;, -	V���B1D���� �T�����RC�FA�'F:D��)�l^RO�y�2a� �v�P��6D�\�u�b�h����l q�Ʃ1D��#f�M/a2�sq"�-�
@@�1D��r�M�y_�0�T��� �"P��0D���X�R�����I
Lg�y�@0D����!5*x�snȐqY��ñ"D� ).��HN��e >G�f��P� D��"���=.abi
 K��p��=D���,ն�գE ���:%��:D�̺@��4k��r�
"��!��	$D�����+^ы�[
�����/D�4:셤TS�ik���( GB-D�0� FܐC�a��% `1$�� D�;U�2�f��A�Q����=D�h����}�����w�t�c;D�� ��Rbo�%b�h�㠍�*Eޜ�"O�5HqK>T�ڙ��n�����""O�X3���l}H��,�,s���v"O����l����ˑ91�P��"O�L��d�0x��ٶ��j��l���{B85�q�'��9�I?
J�f��D�����'��劑&�[-*��"�H�-j�t��'�6t@#�*x�\d���e����b=x�����	L��c&�Zu�l����xZ��H)w���X�X�ր�ȓ\P1� BĴ/	ܭr��	?.���ȓ��$˄�.	r$iПsm樅�D�D(�B$�j���p�St���o���+�u�DiA�@�>�ȓ\?�sA�5�h��$M�,]T���0�N�� (E�xڈ���д8e�m�ȓhA�Aj���5n��҅��0R���%k���A�B�h�5J �2l ⤅ȓS�$Hhg��l�B��/}�݄�!��} �GW�,Fj]�2EL-O��Y�ȓw�P�u�Y�r��'j� +|��ȓ(����UO�7q8�2�M�<ID�ȓ�nɀdK�+n9P�D�n�ȓO�R�I�&h�����(C8x�����*i;ᩕ� X�{��ڭ��9�ȓ
������{��h�bK(��,�ȓ7
��C�^-:͸m3ei�G�d�ȓ6�XD����me"	ӄ��|�E��\���:�2+�N�2U�˝:�R\��?�T�ê�^����hq��ȓ�R}�F� �
(���I-cҵ�ȓA,�!So�GT0�	R�g�\��Qi����+>Y�qsBЗ��݅�o���L&R����CE	K�`��X�]`�h�=I��C)�0�Ʌȓs0�CA�M�kT,e��#�ȅȓc��-�5	�!��g9D�)��;
�c-�_nE����!b��ȓ��!��#U4@`��O�^�氆ȓr�T92�Ϧ-:��A�Z)_�t؆�j��`�&$ڡ��
'�c�J1�ȓS%~䢒�Զ0����
 ��ȓ�:�[#,��t�A���E�ȓw�4��o��.l`���~��ȓc��2���f�����%�/+�4���h���{a�R�r̴�� ��}����d|����4r��
��Ǐf�dE�ȓ$��� �g�8T��$�O3�|�ȓ\|��!��ͬ'� )"��B;H~����-����-�V���I^e2���8$ $�<@�(����F��X��AIy˶jگ5�ޑ���%?�نȓx׼��<�|� Td��V1�Ex ̦!Oh�f�B6��ȓ-�&�B�ZvH�a��c['� ���'d�@��|�j!x��lM�Q��8�F�zх�5���c�IQ��1�ȓXӐaAƥ!
�E�$,K�ttv%��k�xSa.��x�nC�F�_݆1����I[������G'I9R�*=�ȓ#fֵ�2ǐ�G�X(U��;cD��� �:Y�����B�;cKF9mֹ��fw��Z����D�A�b3A�x�ȓMIҐ��b����2��(*1.��S�? t�i6ʨ8T�1A#_�
v��BB"O���V�J�ߴ��tcU7�0�� "O���E�6;���S�?l�li�2"OF� �~�|��C�
8��u"�"O>(J2��	:����� T�!"O4	�bF�N��0qb�@�l���"O�Z�CͅV�i�UH����8�&"O *��2<�4�2�GP�;_�$q�"O("턴u�$P��O}���%"O�9i ���t��fI�l�.�y "OXĠ�oº9�4���S�P���p!"O ����t��UcՁ
21zjm�V"Oxh;���$R��S�ˀm3D�"O�1z��U|h�Z�k��j0 ��"O�dz�f�lx�?-��f"O������P��QX�	�.����"O��Z���Y�t�(b�R
(�
� "O���%ƙ'*�\�f�	Z3�K�"O~�*��D5z��M)�� ���4��"O�\0$��M�T�Z��Zg��%["O}C#2z��Eyb`�>�d�YB"O�ɀ�M���ƄF69"Oʐɐ ҝK�8�e��$',���"O��*��I�E�8@��T)��c�."M�|J$̓4pYL���	�Sݒ��bܵ�f8S#n�?Vxd��$���b4KC�W{`H*�=Vq��˝b#^�0��U�LB�	�*	H���h��/�pO ��۪]����+�ʊ��B��<��p��%R�K����' �y"(]6�T�R��C�L^��&���q� �U*g�:��D���kJ���x��R�H��A���F]�E͂2�x���.IE��@5�
#[��	k��3I�J��DߌV6�(����1d�,����Y8�H��d�%�0�#	����se/�!�����%#ztxCs�O�>�4 92���������~`B��9@���	�'p����_a�Mc��JvЬ��O� Kt�:<^�H��U�;hnmx����G����K~����'�|b�#��m"�"�mQi�<YQ��z�N�)�К!r�Y�+���*��w���!����4$>JDC9-剳c�R��C"��$:(�+/'<���K	͆%{�
F�)fț0靟
}�����lT��F�>��݉�@P�2_���&�66���$\1/a��HWM�8(��E}r�	J�˒&݌q����#�Z�2>�Id%�8���
���T�DOF�I��'�D�#a�(B�D�It�ڪ/���'�@u"�# �DU�`�?u ��ٰ�� Q'�(*p��T��r,<�q	@�?3\�1#J��y"��~(�0l2D��쫠�X>o��\p ���[�.N>q�ͣN?�[���~�8�'F�+f�!\&� �G��L:	�/�Fp(aO<Tav�Y�H0at)���Gm
��֛#s�Pa�& 9ep<��& ���O���}4x"���[z�3���0@�ֈ�'@µ%I����a�?%��%[��VbY4�Ŕg8�ő � O�:�A�Ae؟p�#IћW�,�G�G1xix(��i���,6�M��,ߘdP� ͎�@e|p9�_$�����b%
�g��,дK��z*&4q"O��@4kG={W����iq�i14�C�j���E	��%�&g_FH�\JrF�����ڹ!���F�!�B`�D@�*7�~�*ǌi�\��Z��XmJ"� >1o�(����L��I�p-�%"�Cc�π�9؄�ɟG�D��4$̪�8�t	ޕJ�ƣ>i�D�MĚ��K@�L��m�T-]C�J��J1wS�@9`EXL���R���#��c����5*�B�gz4��À�g����<�-�é�M�`cN |���s�Z�?�B�iH|J��˗x���l@
4�
�>�ȓ6�h	C�V��`�����8��2{�U �*�&��\��nQL�ɔHu�&#�>��
!x��]�W�L-6�)���u���kf��J�jE���֛[�81���'���B#օQx��RN�n}KrkX�.6fYD~�cш�б�FC�EZ4��'Eɠ��OD$��7)�1�"��>-B)�Ѩ�+����Ƙ�n$�����`��	O��?�R섏�B�2��I$��j�O}�|��xB��T�r|"ǋh$L	��M�K�S�}b��#�+6 ���ڴ\׆C�I�\�4�܋P`�Ruȏ<�4���C�Ʃ EƐ*U���렎#�IP*T���S�? 8	AaH9����4��%ixl��O0q�1�J����L RM�&�	&�� ���<)r%�5j���i
�n��t��-X����!C�r���]06�@��6m�����5��e��S()O�%�B���%ѓ�vH<�B֝I�LCS��G� Q@��r�IE�|M���+g1Hآ�R�hi��-��L[- (؀gA_���{Q"O^���ͽ�<d�؆J������Տ}���c���pb
ˋn]��U,�(&*[�DF��R
*Q�.\�ȓjV&��tN����rD��T��Y�vERJ�����I�G�a{2��Z(��0!m�KW�����T7�y���}x����L�O6>�nD��y�@A%gd����9�0���yn��MPFW�2��]R'�@&�y�Ȣ:�rKp�^ �V=`t�%�y��
*�����/"6���yb��%oc����^�%���R�/��y2���	z��7�Y�&��l�g��(�y҃��W:=a�b�ԠS�À��y2�ԃbT�X"2"��d鑉M1�yr�O&1��pX���5�t�0��K��y"�աe�H*s��#Od�l��(��yfҸ"��
�:q,���D��y2��;:,D���E73q��%iD��O�6�"ҧd��5c���Kz�!��) �K�n؅�d�R����Q_Q8��K�U��e�'���)ҧC`؄ӠZ'z�<�i�*V')�I�ȓ,|�� �X:!��a���d����'�"�i ����>e@X벪��4Iʑ8�	�(ga}b�'ϛրO9xaDĞ}���0�O�F�]��m�t�P	�+�XЃEɞm��tEz��'}�F)"ʧv�l�B���"Q�����Ș5썄ȓ_|�!��`��j��Xp�ɲ�F}R�i��"}��a����HA2~�� 9&e�D�<	d�οk��5���Fo�R8�C�Sk��M8�xc �^\p�:&�P�6�vh��=D����c�8~�����#N�	6X�K7�=D��hS�Z�]!~�Y�捳<GN���;D� pa�%�����ab~h:@)6D�h�S%��#A8\��G(SLXh��5D�|�3�Ý<Ҋ9��*�P:L �PH3D�<J N�8	�,z�	��8H���<D�Hx��Շj�"!I ���T���g8D�P;��7QD��D�ѵ./�*��7D�t��ӽH
}(�
N+]���3ā D��'��#�<8!��	:>4$��4D�DYe#��6x�sBЁK����R�<D�`ڦ��H��i��M��`4��b<D�`Z�U�(��A�L�,���>D�X���?)g�����A!y�1��(D�����Mrz\!P�]?�m�&D�D�1g�<P6�Ń���dk�)&D�H�B��c��u�O�3s���1�&D��@���?��(�bfZ�u��p��+D�4�wY𲩹�+)7���3D�PbT�ӹ���D*Ϧ0+����	1D��"���4�����[�I,���./D�,��A���b��'D��/fi��-D��`4�9W��H`�49��r�+D�x��ّQ�2y�D:J
���)D���#-� qe��=+Р� 3D�����5?|��ͮ/+�MRC%7D�ز�K+�Ra�5�*`��Y�ե8D�ړ��.8Q ,!�HȸS��ڄ�:D��C�(%_�J�`���n^��R��5D�� �UB.R�%Gܥ*���S\�<�"On@��d����傀��Y2=z�"O���W�S�@��\j&�Ƞ���"O�)��fݥX�U귌��y�p��3"O�e1�E$}t��4�A�P�����"OȸӰ�ю^20��JQ%B�0��"O�1�M��*x�yI�J[�D�8�0"O��@����V��)ZQ|v�2�"O�d�k�%��i��Πp}|�) "O�)�( x�2PY��4Z�}�"O�h��W�0��!C@�gCք�t"O���e V�c�8W�>/M�@!"O��FG�
�^��qa� S6x��"O^���C0;E(��FF/5�%�r"O:���B�?��=�cE=I����"O��!s���j,��(��E���s�"O*4ШWg� `D�*@ܒ|��"O�e���$��H"nN#��q�"O��FP7G�R��7΄����"Ot,kf��㒤 �+�}����G"O��]U��9J3@��
<�m�A�<i @�	q�XQ;�
��`�������C�<Y��Zs��8Y��@v��ub҇�}�<�qN�+o��H/9�	WD�{�<Y2NG�\�^�S�ϒ��4`HGp�<15M�'.L�P*�=Glp�`�p�<�� ݈�h��.S:_x�ub�OLo�<����FB��pKǟ1�H��gCBA�<�4�t`�hI�`:D@��Kx�<�t�
4��r� ���Bb�y�<1�%�t8��n��7�Ȍe��p�<�����@�6��dE�p��q���l�<!LY�3�����.������`�<yqk��"| AS$�m�b�z�<r�'Ǭ�*"n8>�mK�Gi�<y��C>V�}ꔍW�U��d]i�<q�˳qN���G\��=�aTd�<1��A�}�uGP8���{4ƛ|�<ِ@E�S>n�jG��Rc<�p6�Qz�<I��;���� ��(��X���q�<Y���$�U1q��K:��Q�� E�<q��1Z�<�lH�L�T HQ�YC�<Y�̗�L�Dq�G	j�1`ch�f�<�4c+;�&�QA��)<�q�5�\�<�sKɲ]�P�y�Nή#�|�{]���m�j9�ũJt) �"B�,��9��q����8j�ѳ���i�xh��zP(�ȑ�Ǻ��� I� ��p�ȓ!y��k�FX�.��E3�i˴#%2���@:��qv��W.��6�W7[���ȓt��<����,r�P�A�P3d�Ґ�ȓn�x�P^��!��g[,1��I�ȓ%�B�JBn
<nVx�l+BR�T�ȓ,i\U���i1��Q��Fu̅�ȓ��YRC�:�D�����/:R܆ȓ8w`��'R"Ln�	�2��HZd�ȓx�ɛ'Ś4+cl�Ɓ�v��Ȇ�U��u��i��N�� E�֚p`���$nm���V��AWFU�q� ͇ȓ�|�fɽnj���&<~����U�p��&��10� �R�j
.J�����L`��X`�\B&��?4��ȓM����S�_4B�ph�`��bO�X��c ,��b��}���Au��'�tM��S�? DX��݂e]���	HI2�q�"O�����ɐ\�9��i,7C�|�d"O@�{���Zr��kJEQ/*H��"O�����Ћ[�4�P���6
���"O�lH�R�c��U��k�6y+�$�"O(l�P�3q�"�p�ʐR;lx�p"O���3�р �l�s3oŽ/L��S�"O���?,.��b�9���p"O��k !��)���Sƌu"O�X���Bc`�9�Ȥ,
��"O����u���˅K�Hv��"O�|��&=6Iqo�1k�Ġ�"O�p���� ��duL��6�28�"O��ٴm�I�\:���N�n� "O� [sGQ0s��0��ȠO�P�"Ob�4#�3^8Q	XB6#���yBᙿ7͌�ѧoO=(-���E_��yҊ��Ov�@��/q��Id��"�y�$��:�p�ɀ/��rtN��y�`�
6��LJ"��:vr��2�֟�y��H#�̀�oԯj�љ�kE��y@:��q��l�I0R)6�y2��8 4�=�E����x����y����╡����Vl:���y�e�2Q�)a�	�j�}k��C��y"�>k�4u�Vg	J!�XA�ם�yrm��7Dq�Qe\,V��P"sV0�y� ˡ>Y���f�]�KN�xa�L�'�y�[�.�v��Ȱ2E&}�T���y��_K^yI�GɣX��-HT���y�!��lb싃���	X �hdH��y�O����+J���(82iG�yrJ/ш��W��6J���L�&�y�/�W���A�-�B�P��Y��y��]�V�nj���*o�ٸ�� ��y"@�)y8����Q�Hvd|��`�;�y�W^nNY�b�ۖ?���i��8�y�e�T@�3"j��-��T�eL�ybj��P�B$������A��y��]�����$����>#�`��ybJ5�(E	VfM*8bՈf��y�):t������j���b���y
L�Z)	R�`֬ą�y��U3k�Lq$���z�p�6����y�Ö�z� s�$G��h��o@��y�k >}
�at�]%�F���K��y«}zh����� �"�D��y2(ϣ@���:�I�3aޮ%8�*��y�#+,�u��]�2��Ο�y��ߊj����5/ӑ]�jY��U(�yB@�3,���!K�^���bP�ݫ�y¦1C���qC� 9�ԋׂ��yh��$נ �D�0XH��&@$�yb�WP��ZV`S�6%�����y�O�;Kf	b��G!N�H䪢Ǆ��y�Gp�ӓ��(k�pu:R+M�y�.S�4w�m�g�ћh�|$s���y��K�|)F\��:6�\�hA(�yB1\��yCF��"C@�����y"
�_ݖ��A��qc�?�y���'L�Łэ�Μ`j
+�y��ʿx3j���b���ƸK�i��y�J�q<�E �̔���90/���y�.�/:�]*Sk	he�ak�ʵ�y
� Z�@�* P���9'BHд"O�* P3hy���E+��l�b"OȠHO�=L�2�H����x"\�R"O�A{�/��xY/��/�(��"O��j�NϭAVA��Nņnj­��"O4!����OX<q*g-�n�T�"O�Z�6�F9�4+�2,��}�q"Ov�:W��� �AR��Dw�8D��"OR}11H�2,��攰���u"OL�:��"1��h�"M6^����v"O�="�-�o��,����}k.aCP"O�\�t�_����)-GҤ�g"O|H`Ŧ�@|,��#�S�,�<]�"Od�D[,g����z,��"O��㔌�+aJAED*(~�`�"O���T� ���U��M����%"O�	�OM�0@�:Rn�3�t��"O ����«-�,����/�p��"OP�h2Kɓ3�j��a<����"O�a:Ӌ�����w�׭*i�"O���ծX� f�s�H;,r�˲"O���R/�Y�oZ�)Q��"O��y0',5�2���a��CSN�	�"O"�ӥ�P�Dƅ@��%I���"O��� A�D�$a�Cg4��k�"Ov�◤��.ƦX�F�]9�)��"O�l��I2C~2(��$\�Jr d�"Ov5�Q�N�%�\耍�puN؊f"O<�*�+�q*��x�̙e�0t��"O�J2/��£�T,��M�3"O�� Nׯerx�a ��[�(ٲc"O�L��ȇ22 -��Ɏx�,�7"O�rw$�'N��!�ʘ;3F���"O2�A&&S�ڵ��\��@u"O��c��cX�)I�V(Y����S"OĨ)u�&[Ĝ�A��ej���"O�H��Ɋ}�H����^�"�u"OL}Jw��2n83��"W�\�hR"OL@���69<T��p}����Y�<qAJ��:()V���*��Cq.�T�<)�*G�u�P�c!#�>9,�䳅��W�<�&B�=!��H+���8p6T��+�d�<Qbd�|�x��e�^34�Pi[[�<q�!�^6:��+*�
hYF+�^�<�"���o���!7'K!b=�L3/�]�<!�B� i�,I���(]��S�<i�@M��ɺ	Q���u#�J�<�����K0ZQHQ�\�o�Ey��C�<��#؊^�]x��Ќu:�લI
D�<���(wI�P"r( �+{Bx�dJ�B�<qə�%����*�ht�t	�G�P�<�q��p><���h���l���[g�<a�J��:��E�.�R �Q�R`�<m-�=N�Ai��G}���3#��_�<��B��;r� ��dZ�2��} �DZ�<iD��=ȺQ�ŏO�ANT�;S�s�<	`%�=6o&��vÛ<��-���Zd�<I��وa]LEXы��쐱K`�<�sjZ�ń,���#mMJa4@Oc�<i��ĉ#���ᦄ�~{@��c��D�<I�b[i��@V��V$��j�_�<�Q�T�<%�Bw�
4۾Y���JY�<ASf��_�uH�@Z�ʬ��)�T�<y�%s��uġ�D���z�<� J@�WbP�F���!'�l�0���"O�٢d%��{�DT��  q�ԥC�"Ot�Qb��-˴��6�A�R�X��"O>�s��ʪXĠ�0����P��0�1"O�� �[�L+�!�d�,�>�"�"Or(�`�0i<T�����|��)�"O�(�˘:�݀���&��h#1"O�j���̴�@�o��6稠�P"OViZw�W�s��qgT/1�����"O�	36O�>�͠�P�r"%�� "D�܁��ߎb)*�����=�iC�?D�4HǉV)Y�|����o��B�j'D�H���	c�"i �O /j�S��G�l?�H��3�O:���4~��k�G��<#P ҳ"O���m
�`Z�A9Ɯ��I�1&���i�?��+G-KxJ���u�H©'�ɺL&	�?%?��jK���.`M����$}"��<��O���� ��ܼ@0�&:P����1�O:��%"�)�'_o �:c�
-	�-���9wJ���&�.3��O�?q�p�ܽ��1��ʌ fR� ��[��'e�|��ӵm�h�1b�O*�%(��޵X���A�l�S��(����%���Sk\"r�'/��)R����{hՠ1�V�O[ppsL?E���F)� 㟢}�V*Kf��H��zv��4H\�h���h6����yڜ���ʾTT�l��>&J���$�	�bc��+�PU�}��ɀ&�lq:���W���� i�&z�lJ�>���V�I"4����
d�� ��ƛc0���%�߸7J�H�i��1��/\���S`�O�*J�aE�l"@�PdIE��*6=OT��6"�0
D�	q�O
�j!ND�b��Pb˂
�Vis�#��Fp(Q	(��d��<E�D#B,[m����$�
	�}�V'ȉF5 ���V�L��'@L0�}L|JS�X�^����� @̘�����D�=�֬I�K�L=��S��а���oN��1�W�6���(M�y������
�c xa�L3���	��]��peT�A������/Y����VDap�

�*����Ox�U���s�­��T#I����';ni9w	���N1��.�0|Z���7�`9��,�?t����@�%k�x�)�3k�`��PǛ �y���'X��1i�O>FX['�(?��͓	�'�iѦ��3ea�ve_�YpR	�'B֌8�D��nُEJ�2
�'��ehtnC"S�.�(e"��~ݰ]X�'��'+O�� lQ�c�>B���C�'vR�#� ѓVL`{bT�5؉@�'��$�3 �)!��D*�lتy��p�	�'����OVް�	�ʑ�c�&�Y	�'Z2=��E�#^���#"�	�f��'��=�'IK2hY��aJ&�]C�'sZ�� "Dpa�O��w�H4	�'3���3���&�8գ�*d�0��'\}iΛ�D>2����g�l��
�'���;`�T�Y,l�ȅ�@�\mk
�'>���B�Jnz�Y0O����!
�'2���Ra����Z[�B	�'z5��c�+&k-Cb��P@<%��'urd`r哛`%��ёO��H	�#�'�~c1iP�c��pҩ��H����	�'�����I��df���E�\���'A
)�E� ��J��B�$(C�';>䈃�D<m���C-�,H�R,��'oP0KD��9���d� J��Y��'ev���A�!.0���g�!<i^���'�(c� �t�N)Q�/gGp���'E$]��*ě+�Ш��˓��*�'d�� ���"Fu0P�vb��'�H�ᓟq¬�P�G��><�z�';r*�N+&5�򤘡c��(���� ���BNɫ)aꌢex�B5)�"Oxl��S�}���"�X�g�&��@"O� P!BEZ�V�P��3g�(�	�"Ob �+.��b���#U�I��"OH��a��v�~�Q��aIX��P"O��S�FR-Լ��UJ�;���"OT; ��B�,�9^Y�p�@�<1����"5���~�Z�Kd˒~�<	c�_50�2�+�N'~�`�dLx�<�EW/z.�X:��
=j�sP�TI�<YV$��3��P�R�f�[!�k�<)P�{�x�KӸx<��{�<1��G!8*	D�|ߚq�&�Cl�<ѵ��2P���0�٢��[A�<q��M�yX����rr;UɓX�<q�'ŀ4l���R�J�T�jDm�<6� ,u#T�Ȕ�H�*�d S�<�&�K+)��0��5"�X��1#�Q�<Q2/ь��т E4������P�<Y�m�(>N�z���(l�t��h�<�UbS�o���]'`���yC�M�<ɥ�=L��3�$�"qsA`�F�<��Ծ}�h�� �v%��kw�	D�<3"��q� ��g�$B���� }�<q�[�2V���IB84����Ѣ�O�<��#�>K�N��Pޱf��`G�	U�<�2]�v��=1t��a4i�jEU�<aă�oԜ) UHR2eѲT��˟H�<	J�
ߤ��6��C�D�R�E�<�I�'!3:}��C&>@�#�͊g�<��N�GFzR��"*"���[a�<٣o�����O�!Kth�:�k�\�<1��"���P�K?N\r��`�<�p�[�%Q�P��#ً_��
��W�<��D��Z�J�iț�K��w�l�<���8c��sƉ��ԡ���h�<9Ub�.R<(E� <�P�C�I�<�7i��<�"
 ��JR��D�<I4��#x��)�O�9b;hڑEQ[�<��&/|ɲ9�c�W��Y�6�\�<���S�����,��SU'	]�<Y���4,Lz��%hIq#���B�	L�����$��R�`�q�HϮ)bNB䉎j�6ar�ɑ6H�&�UJΙNB�ɮ??��j�!��;}83A� B6B䉯z1�Rc�B��"��UGB�I�jj�8 �T�Il�
5��n#�C�I�I:([1Ϟ>J�>�q�7$C�Iq��}�����j�*0�(Ǘ5�C��#�Nd�t��1��T1F�³)�*B��0�K4a���$I�i�j�R�"O���k��xQV��p�v�F٣"O4ȁԥ
<@ܪ7�,1�6PI�"O��z��ô8�Hm�f
��~�hf"O���rA׼�B_�d�g$�'Z�!�$>��p���;8�Rש�7j�!�D�>1�%1��#u"���B��[!�D&,���NQ�V�dّV!Y�!�D !KV8l���#���)�!*/!��Ǹ�@��ר�E��H+��L!�DΨ-|�x��D!Z$Ԉӡ�ʗ
!���T������'?�-�t�˲b�!�$u[z��6+��R�R��$��!��I�v��vK��b���k1& ��!��  �B#�p��|�!�"3V���"O�-A$MM�t@z
ҽ|ת��t"O����I$,�I���*�Ș�"O�h��Z�b0Bq��/�����"O�#�ρm&���Y=W�fh�"O��S׮�/�5����-��UiQ"O�(�V�ɶ\���Q�MřM�[2"O���W�i� �!E�_�t����"O���s�ѥI�X����L�u#�٨�"O�ĺ5�b:
��k�p��A��"Op��H	W~�����j�D�X�"O��0�Aߨ���ʜ�~~(�PP"O���v��99��R�K�j��3U"O"9�S�&m�f�ĉ�6hp*�"O������#G��H��!�bRP\c�"Ob�C�A=s�8dP��74�b$��"O,����b\4�&�� Y�����X>� �j��eQ�M��E� )Z-�Dg:D�@�D&B�d� �s�I��aev�14�,D� bÁ�Z/�,��J.��Q �+D��kX�s�	�ea	 / \�q�'D����C���
!�T�$�D�An3D�px@B�, @�p��(cL<�d�0D�X�&	-'\�Sf*��z�h�&!D��-�U%Zaj�
�`��aL9D����d�(T�t��df¥[q,�c��5D�pu㙰'��rqN�I>�� %� D��Ar�"٪$@Un��B/>D���tI�F���a�a�����#;D��(P��&4~�@���%Uz�ͨ�:D�� �'Z�L(!�N~̤XVM8D�\*��F�t����m^��x�#<D��;U���:��q�l@�6�
�m:D�����ð,{t)�W��7{���(�:D�H�^�O���8�(��cAt);�#9D�p��.8j���kԂ�jIt���!D����gқO�v8	AA0֔����?D������ QTg0�й�u�>D�p�w��+���ЮZ�����h;D��ⓥ\rex1[��Z-I������8D�x���ٍyȑa�*F!xER�M5D�9�I�U��E�5��y���Re6D�(�a˜ �.�+�C��^J����5D��+�Q�Q�DI�L�8D��4D�ha�3,��գY!H�vc�@!�$�&-LI��A�d�@�mǎh!!�D��0�th��U���ň!O!�d����ک�[wሳ{NP�� "O8u�e��9ff�sD/C4�`d"O�,0]�0+���,p0`!COj�!�D3Q��$��g:1J��\4{!�/b<�Mb��'?Z����z!���4�F���!\$y����q!��p��t�2�
�8�^D��oT�2�!򤟵QD���I�l�\�SE@G�;}!�[7VƭA���'�h��c�ܱ6j!��$q*�A�ʢ?�4�m�i�!��&G��#%��-na*U��e�!�D��g�Ht�Eņ�eZ�+�Ñ�w!��_�(�b�*!'�"�A�=t!��Z�(������Īqh��U���b!�$X��q��ӯ>f=J���!�F��@���p��S
O�!򄓥p��h��L� ��aq�\�!�� Ҵ. 6��� �H۠e�┡�"O�uBa��)t�ȼ�s�Q�g��08"OМ��m�A�$9:s�W&�R��5"O�e��T��Q#���Ը�`"OR�sF���豆�O��q�"O�qi���=gV0��G�VaI�"O����%��G�\|�/Ӥo+� �"O��EG�	D ��� ��%��`�"O�`{�.ٹ{�H����1�C(�C�<9�·
�ĳ��J�OI�1����@�<�@��g�(a۲kR���ِ�"�y�<I��; V����0aE�m��Am�<q�M^65v:���@�qcj��MUj�<��dR�9 ��k��X6)h���^`�<s��Y�8JFNߍb�0(i�AV�<�V��2�<�meC�S�i�#�y�/�k��0`ua���QCV��yRL��s�A ��މmB�"��.�yE��A��cĥ[�e�剁'�)�y��֍CbL]���� '��Ƞ�ˏ��yb�+1v�8�	k�Pxq iͥ�y"�@�O�8��ć\ S�%P@��#�y2f�����'��X�Z��;�y	�Y4Tlh�� 
5ڲ��yrf�*�0�X����XBs%E�yb#�]�`��Dϭx��5k�'�y"\�N��4��$��B���1�y�%�2pپ�������sUe�3�y2�� N,�j-�^,p��y/�;	V%�&f؀�t�0�گ�y���M#du���^�
x�p���y��ԏ}��y� /�H�����S"�yBG6'̑+r�J�9"��
0@���yB��-�����2����Ó��y2S- 5(��ϊzv��� 3�y��*���9���%R���`�.�yb�V�]�:���)��Ɯz��R�y҉� �D�!6��<N�`���N��y��!7(�P���>8�>\�Ь�yҢ�P�D��A�^ ,::U��"��yB/�>N'�@��R�[Zmy�h�	�y��^�((<��$�S����uBQ��y�
��    � _F���"O�	;���V�V���!2'�d�"OB���+�x�`7A�1���`B"O�X�
�w�8ِ��=b��P"O$@��(�Zm���%�n���"O|<C�L	@xps5#]�>�T�؅"OrQ�p����ƭd��:����'�l��E��\�<E	�D#4ҍ"
�'��]���U�wKΕ�$DM�a�r��	�'�~0�E �aH֭���/a��X*�'���D)��d���"�K�S����'�܅�T�f�1�.�dH�'��H)VIPH���K7GT%!�'q���g",$B��KK�*!�'^�a�� wѤ�E^4;a8I�'6�8 ��:�DҦ��hB(��'�$�0�D��-�s�2؀��'
��@��R����^6wzN-��M%b��F����;G`[�bH�-�ȓ8����5g�/�FP����)5YƜ��5� 0�B�.bDI�֊��B�
��ȓA,��cAJ�(@d�bE�%]��D�ȓyL��Iu�>O�Hk���c8±�ȓ;���!��.\qU��z���ȓ]* !�5	�<9���;����.�����J��y�2�P6��%L_$I�ȓgeJ����N�VӐ�����[54��`"	b�'�{��{��z,��ȓ�t� -�(�`��c�M�$�d܇ȓ@���Ԝf�j!8u읒��A��.\5�u��;d���Pሏ�`Y�ȓa�zL���2x�x��PN�	�.؆ȓ)\������,dvxK�"�*. ��%��#�)��r2i���`+v>���pO� ����.����!:*���?u�YT�ˤt��H���J�z��ȓ}u����+˄�dYq'KK���/��˳�@%���0����0��5dֈ�g�H�A���(ӃB4:�(���
SN���'C&��1�h׊;)�0��~0�j��R'
����������p�#�,�q����a
�-�ȓX���ɱ��)"t
5�@�=C�4���'TP�*'	{x�
&�Q8SC��ȓ����Ũ�腂�O޶n�ޥ��/"��̖/h�x"aJ	*�p��!ZġS�*�@F=(%Ǝ��hm����Q�@<�z�3�Z<T�y��om�hrŨ޻�@9�2�δ$����S�? ƹ��⎻/�d�0�(ѸDÌqsp"O�8(���#tŤ� g�8m��x�"O([W��5��cW%��
AɁ"O (d �3Pc~Q`�Dˑ;b��"O֠����Ӗe�fB��^9��"O`4���Q�*��( �1�<���"O|�S��m��1��
����{�"O�$c=��|�F�>o��P�D"O([D[�i��͓�ˈ}h	`"O���UG�KB#G�@�S���1�"O�ڳN�+("@�*�P=':���D"O.��E�
�1J�a!�L�r6�p��"O�U6LѲC��u	w߭]p�bP"Ot����Ԇniq��bb*T��"O�!�4׮Nj�����aC)�U"Ö�>"3�e����i)�Lh"O&�AFh4/�A`�F̿.Ğa)�"O��
`.�7r���u_���l��"O���1��S�L��T��<QT��"Op� 7�_y3�8@�B'h\(��"O��a�}� �
̡?VB��"O<,r�B�dǮ��®ߑyJ
�B7"OJA��	�-A���*GO�|=B�s "O��sf����Ap.��_6(�1a"O�m�"�'�@��^�K#����"Oh1h&F${n`��D!t���"O��Ab�ވo��l\�����"O(����-z(���v�K:�l��g"O���"�KRh�#n��7|� �"O����j+f�qY%k���y�"O\�s��Vk#�@Z2��4��q�"O$�rI��m\�����(���"O<��2�@"� �ZŔ�t5$ő�"O���D5>���hT.�l�Z@c�"O@�1��Ɔtl�m��"�Td�"OPl(r`ЛJ>h��G����"O��(�ϔ;	W��Q�#�+@�����"Od,0&j�_�n1��'�@��U��"O�)q�&^�Ć�`�+D��ra"O$|I�.�q*��H�)L�@s�t��"Oj<9�n��|��y�'�3rk����'�h�`�`�h��F	'��'�t(6Œ&
���U$�k^
�'h������L������[� ���'&��:�j���R⡌#X���:�'�j���& ��!W��R�'R�Y(��̂Ef�9�+�:x�5�
�'j�hH2j����i>\��̀
�'�,��)�3�<!:�kǈ^Rd@�
�'7�!���-�^ɫ���j��$
�'l$ [�)
2�����%m��
�'EX�Ӡ)�^�.�^����	�'��P�U�7G�ȁ�D�M��5@�'܂	�dI������oBH^��x�'���խݸ?�@�3!��::PY�'�P�Q�T�pl�-�'�W�7�8Q�'��f��)� �6@�'F.��K�'
���O݌^���f#�9@9���'�^$���J�r��;OV�D� y��'�A{�l�3]��RtL߁5�R�"�'Y�Q���Mh�
t���3:����'�r`*&�N�rv�$F��y.���'�F���@�3g�}�. 2���'����dP&uNE��ff^���� D���>���ywhS=z�P��P"O~���ÏOF��CC����^T�"O�@S��y�&��N��B�q�"O��t �*�1�M�"|��0t"OT���F+B��#�u�Z8:�"ODay��Z�Y!�=RW�[���T�"O
CU�7[�Պ�ŊO�JH��"O�ʧ*�)#�=���[-&´�#"O���b pZԎ� ^`}""O��c�7�\`�#Fds��;�"OHQC�žl�<��E�; i�iF"O��[t@@t�	��A�Np��[u"O��ᦗ.Fk�%�������"O8�-.-A�i�H�"O\}��)�q��p�߫b��4r7"O` a��,��uz���	^E|��Q"O�-!�N�/g2�˥� 5C�eҁ"O8��%�qרY� lЦ]F��q"O�}r��=E�K�H��/*�P5"O�DX���/ �zh�$���\*�"O�HE �Y��L��k���:�k'"O�}��(�t�\lSEjJ�5�,��"O@�@CaA�^7R�[��T�^b�\�"O 4��dF48��)�@��+\Rʅ�"O��9�LL
I|dU��-]�Pz=h�"O���r��){�|����C�P���g"O�(�4#̱t�v����7:�c4"OX�`�JξWm �h��t��%a�"Ob�9�M�P ̈H���u̵G"Od���R�m�Ղ�P�ML^�҄"O����ၞ!���%��:2H G"O� �r-Q�(�X�U@� �"O��;4�J�p�fc��>�17"O� r):}��i/ڥb�P)&"O�8�Z�*nX*wL��9��mjR"OJM��];~��e3!�|�Q�"OވX�O?z���1�	�*m%v%��"O�#�)L�X�[1GW�D�h2#"O:11���F����� O����"O �X�O&E��Tsa�X�I*��"O���`��%W�Q)�dhT]IT"O"���x�t��D��;h��@Q"O��ns�R����	|<y�"O޽ w���2:V��W��+&��=�T"Ol�3�N9Y^�E�5h��0��1"O�%�4�Β=j����&.�\�"�"O`���68��3t��&3h�X��"O�I�u��)a�b�Z�
�zY��"Ol)�1DQ2@÷��InQ��"O���']+'����gL�;E�Z"O4�hA����F����"Oh�C�h�^�!��QQ�z�`S"OЬ��&'X%p`��:w"O�!�B@�D2��� �Gv�"ON@�eOO?L���g�ʄ|;�"O<�j�ʬk�`�v@ Urf �"OJ��t'V6?��A�Ϝ�\�`�E"O��!��4?�\�a���X�AY�"O��Q�B�:�S�X�<(I�"O��/��I��O���� V"O�9kA�V��p �VQ����"O�{T�,7�4���H�&��b"O�i�he��C�40��)�a"O�)�p���1H1��D���s"O� �A�[/f8 `c�	 [dM��"O�����ł zU�U��lUtq��"O|ue��[��D$D��B'�2r"O�}��%� ���"c	,w !�d"O���P蔣˴<�#�d|]ZT"O�H9j��|s�"�]��l9b"O��[ ��+̴;6�ԙW:`3V�'���Su���w	P�J㌽���:يX�7$�!.�
����O�D�t#�������(F�,�H�ض`R
M�m*t-_&꺔��J�m��҄�<u�Q���S�dˣ�E�+��aH�'l�]��hK�^��S��-�$��Q��<@�P"<�'(��w�(~��s�#Ĭ"���M2L@�K<���?a�*�Z���cƱ��P�O�IĝHE�ODz��)=D,�����	� iwM�V��[�"ش���S1k�&Un��L&>�K���L���0ŏ=��H*� ��ǟ��f;uF>ē��>��V��_i������_����]�mt�D8p�ɓ3��<YQF�f4*1���P�}Ę��cN��U'ąl��{�ϙd����dO$r��Q�R����?��i����6��j� 	Y#DK4v�б�#U=�]�Io�S�O����ƈy9��H�pN�P�Hގ�p>q��iRh6�f�	�i�Qh5j���K5�lhQ��&�M'̇�P�F�'Q�I�?��SG�	�0T{֩84��3CB�/�ؑ��]�*�J@�>	R��B����)��T�EO�c�d�ϿS�
	4v�t8f���K*������A�@����� �E�8!z��)�%<L�C�8�s��Б�G�"D�M��@�F��]+W�}���� �'�>6m�Cy�'���V)W�uÄ9�戶6I�e�V��~��'�O#=1Q'�\F�s�螿ݒ�z�̕M�'2z7mڦ%���ݺ��R�Mr��qA�O�-̢D�+�b�'S0H�q��;H�2�'2�'3֝��Loھ�^A���M���X�K�t�|1�Q�[�~���߃O�,�Jf+�>��t�iVBI
K>ao��c
jyK$CGYM4�s�&�>��B6EZ�@�� �;_�F	�O�n�ӂ���6�e�O�m�o�*�AH�Ŝ�zv �3�J�����.�ٟ��ߴ�\�gy�'+�������ֵClI�@J�(=VMa�'KE��LL4?#z��B�KlB�#�4�M�i��'���I6�O2�I�z6�\���p�x릮

,�.$�hӼ`�~���Iʟ q�^�Z��x�4i�=Qr:���.�k��`�5ǌ�~�>MC^榕ؓ�S�8 Dy�'��͛���
�bW�`@I��J�5?8��*ĆJ�%�q��٭Z�J��Ӆs�'|�pX��=I�� &\����a�Y��@���I)DY���'=��ޟ��'�h��gF=M � ��̏"�ٙ�'�$r�jц-!� ۼ?=�'1B��6kӴ� ��@�����$�O:�'tF����S�-�+�Z�،B'���/�"�'�Rm3N
� ��	E�a~8-���l�<֝2��;3і0Y�t�wgˋm�
L�5�<�t�]:�5
t�A��[�
�B6+�#g�)Y��UaHQ��Y?,3P!RT�Ӌ5����N>Yt����޴1N�O!�Vb��l��(�a&C��6��s��q%��D)�)§��dL<T�V�!�LVd��C�	��|�a�HXm����[�s,�h��_����gM����I����oy�O��OXa���  �^8
��O
���O"���N0k@Ε&T�1�do\mh���'��'f�!�#b-������I?
s���c̏7>
f��0n�[xR���}��[��'c��':�ˏ"�0R�Ą�j�L�0Ӄ��6��6-�Oz5��LI�	Ɵp��ݟ𔧿�B��b�|����C>E��ݹ*�>Y��c��?9���?�-Op���C�B�$�SgAR,�bǉ54��>�������dN�����'ꏕȪ�+d-޵Y��(���O��O�ʓv�X	�3�8aF�6�X!��ǫɞ���R���I韀$���	��Z%�b�#a�D9��� ��b�(���-������O���O��~ƶ=qf��D�xu8�֪���fE�&6m�O�O&�D�O�|r��O��'=�Md�N&TD�� t��-��@�4�?9����ć;*��&>����?���r���rL?���pH����?���Q�� ����䓉���R?3�Дqq3?�lyBڨ�M�/Oʀ�BF릩�����$㟤��'�YI���]B�`�!I�Nx�%�ܴ�?I��-���̓�䓌�Oq\(�I-L�`98��C	2�Y��4)2ٰ�i!B�'���O�0O���I5L����1$Ԕ����I� �*En�~�0�	ryr�'��ry2�'P�Y���}�����M�7����$b�`���O��$E�"lI$�x�	ҟ��+AP���κg��F�d��mnk�I�Q���)J��?y��T� Y�կ�x�3�F��� ��i��Nt��b�h��s�i�yc�'�& "���&�� ` 
��.�>�D�?�?9)O����OT�Ĥ<��`��H�~�� +�����q�
��HS���O�OF���O�`[��	>�0���9G�D��!�b�d�ġ<!��?QM~r�oͅ��޷_؀[�/�>.�dS3���?9����?1��.�|��'#�.�DvH�`b�>�>���O����OB�ħ<�4�}�O��mqF	]�h_%R����=���}���ĩ<���?��d,hd�*������鲩����@�B� ��*YoZ͟���]y�%��`����D���itV�_˦!`��?F�9���s�I۟ �	cN���u�	m�'�
 M�����;]}�a �U���'0L���h���Ox�O���� ���AQD ���c@�L]oZğ,��
[d��c�I]ܧl\~�G��%e\T1D� y� o=X�V�۴�?����?��'"t�'n�㈳=��z����E��ā>7��6V���4�9��Ɵ��G@�l����#Eu8kR֪�M����?y�1�8��b�x��'2�O��p*��:z\1�WH��t�-9�i�'M6!雧�Ӿ�l��q ��t���5�ė%azND�)Ҋ,�!�d t�l��H����0�(I���z�D$v1F1rR�*4�=(5'>��<;!nL%RzDE�sg��D�B�ɼ֮��d�Q�/c�h�-*���{�kG3~"�%X�a��po8�AcQ+8d�� ��
@��AՁ
 ~e"���o�}�%J�B	 x`0T!,L�=�#.R�jRV��קN#d��CWǜ��(�9���M@,_��?���e.�]I��?ٝO��d՝3��m���j���E�,8���%$��$dU��p<�@f^|uԸ�S!�	eA�ћ�4�4�D ӏy�֙)����t����ɀM?������]�T2ю��#����,��i$Ցp*/�I\��8A�HZ�t��<*�-�cGL�':�ĺشIЬ	�&G�I'2�)!���>aϓ��$�:#2 �'*"\>�(������a�
�}KJ����F,���������ɽ�p��-��{�=�r�J�G2�.��ʧl�] r��:ef���/\�{?N��Ojp�"#ң|�� ��ͥ)&�D��%ܺ��H�N����%C@���gb��Oڢ}���ok��Q���)Yf�}���)h!��ȓ;�P�B(7t�ФA&lU���݇�	��HOD%Rv��#du�4ƔiU��Aw�UB}"�'�j�j���a�'�b�'���� �ea�%Z�Cv¥x�׮#k)�v`�2g�ӟ�C�\�f��c>�O؂�C�`Ġ��!o��u���4hv������P�ծ��9�q��'�Z0bI�)9J��V��:l�@�Z4�'��i-`#��|���dTA���uFKR�h����0Y!򤈐fĥRP
���xe��@�'V�ɏ�HO�Gy�#)	�) �%h�qj�	��j��b!R��'���'���П����|*3(D(�YI��^" �A���x$ ["gZ�g~Z
�#�Y��l�p�H>��X⨍,\�勔G_� XXl&%k�1���Bj��D���_���J&H�O��W'����D�O�=����� ,Ό�# 8z��M@��3�y���C�
�@bi��B���u5��y"%�>�*O�:q�Kp}��']��JF��7���O�%�u9��'T�8���'��ݗ�����-[���p0Ɩ*]*��0�3� �8 %V4C��i��ҁ9��I��$�>��9��Z<g�>�RPA� �00�,�k����iK0(rh�x���,�p� ���	 K��'@�8X*���G��<�\{�/¹Oec�P��If�5�o/1���
�#t:�"<Q��4���l��q8EF�#U��ȡI�i�,�	Ay�LU#k�7�O�D�|�r���?��!ˮk��PPWAl�d������?��}F�h�� �lY"���'�o���T���&\��-��X��"�xd��L%h��5yc�>Q�7y�.Uj#�F����L�P9���2"�ي �Xl��G2#^`[T��Y��[�dG2�yӊ���O�����P��9x& WB�T%��0=���Oz�d�O ���B���0�8`�T�1+)P%ax��7�!rj𫄢��G�x��c�L)e6�hz��i���'l���.u�><���'"�'�bem�}8cbFM�m���ʹWR��sAE�R���D\DDj4�޸#T4x�|Bף�%;��I�(氼���S��p�	�J�B �����"9$aЩ	+~�R�>���[�BG�$���:8�(kb^�*2!Y k*ȕ'��
2��Oq��'ϔ�"�HN1��9�gQgh���':��p�R(?G8؋%뎔8)��H�'��k<��|�M>y�P�g9�$J���<U�lh��G�<�`��1��p[ӌ4Ze<�qBEB�<AF�f
@4�!��~+�1@���|�<���&}�A	�셆r��Nv�<1@��� �Jٴ	�rPdY�y�"�N�H(6�.X�蓨��y2ǜ�6]���F��{���ѣ�Е�y ���ᎈ*nи���/�y����x�����k�=�����
�	�yb�8GvR�
2�:BD��G̒�yrA�;V���A$��$:�
�j��k?D�LA1/�X�9a� ;I�^��':D��(3$� �1�� vL
�7M#D��e*�b�B!��J��S�<D� ����qo�q�e�J�6��u8�F6D�̐ge �|�n4��%����1�B"D��� K�+�p	x�C�L�z	!��-D��B*�29cb}��,C5 o
���j'D��{�#9!x���ԙF��q�`$&D�����,d��=p�G 5o�U�$�"D�$Hժ@�7��a�A�C�$��E�K D�܊�"�O��	cŋ׼H6tE���<D��R@*�f���!��^2pѳ%J<D�� ��f�Q�g��aoRe���,D����!�K�l���RY&�� 0D�pȔ�R�]�� �*C8B���P�C/D����CG����_>��< @�7D�����$a�20�w!^�B��Y�6D�\*�X�`�ƜѦ�^�#l��O5D�dzB*�y2���L\�'@F؋v6D�ܹ�́0��1B�AJ\�*�2D� �� d�:��`��R:$�h��%|O�]#�KR�f�Z��u �5QC�?JXuz�":�FB䉜I\�X�R��5e��I����%~ixc��zr�O:�&p;g![�>V���&NH��X��M�L��%�A"OP�ʠ�.(n�}�CBR	I�DAt�L����Ϸ�$�� C�#}p3O� �1�@���X�V������15��)�"O��q�B;k��` H L����៴��!FT����!(8���hO���D	�$���hR��?3��:��'�
��c�������C�x������u�8j�ɐ�R9�x�sH+ZQ.]��I�Q;�"��]<`\��!!$7�c�hJG �-!}F�ZT��?6q@�s���O�<Bp�T ��ҥ\N:(S@I�6HC�I1O��H�`�7Rh����HM��Љ�� ��}!�.�.;.����S�O~��*&bTR��3j��s��ɠe�B䉾O�V���*`ز�9T�
m�����'���@%��ժ�R$mݍY�g �]	�G+Ԕ9�spL��$�����7��P�F�x: D��l�g��bRl �W�:�a�e�Ц~�F�*
�}R �����I�� AGeC_t�I�>�T�=5��hC�F��&0&(�u?���OK���'���l�y��99d�b
�'�p	�eofLJ Ӆ��+-\ �e�~Vq"¬H���ʵ������hg�A��O��j�82���N-��� ;D�L�AE�0����A��856�˓%����DZ�jm��/[�*W�8����>�#�FT�	*��S=��ѐ$��~؞t���FZ����!V
��B��-E�<��E�����d@�i�H��V��q\���	-W��3���%&VAW(С�0c�p`�4\�	rĀ&�Z%,}l	4?"j�kSʎ&����M�;�!��L�^.$q�S텥M��ɢ��P`��%��J�zU^Yؠa�J���O�O@$�?t�:�ځ�� .l)���,$�B�	l�T��-XE�6���f�s��!�J�l:'/�cfjT�;��}�$����'�TA�q��Wf�a�S��=v4�#	�,��4��Ȟ9�Ԩ��\?�|��J�VC>=�&�˞����'!�c1��3�p=�RGјw��QpR�g�4q7mR�p��L���[=����C�Y) �0�u7�;4h�P��
<�rYВ�H��y�N-F8�X�f��`��d�
@&n��`�+��+6��
�T�a �Sܧ��S:r� 0aA$\��t(��&Z�!��.g���#R50��򤓮Ya��q��Jb�0�S��a�:����	f��p@ˇ��d`tѣ�(��z𢬇�:tRN�5a�:r���4��©t�I��e�'k瘨HU��J���p�E0s�R�)5�ۉs3v�x�:�ɬ�^y��*�%WA̠H����Ņ�f�x г"d%�T�Z�w�R�r"O���6���TA�tZ�ˮ!���X ��/*IJ�]��:�Dƾ%�>-��~��X�ρVm��&��J�l���w�⸳t���dB6U�E!�Wx�p&��(�H"lC��}rc��?�>�4�[�{��If�Ñ=cԤ*�u؞|:�o��%�ᣢa���z(k�L��02��2E�~�`3���v�(P��	*:��e�׷{�:1&�ʓ+��\{v���t}i�7ta0@<�dN�.f�c�6i�,���y⁜�}ג��6��6����Qj��Ȉ�s%�.s�1k'A��|e6��O����NF��-�cj>O �s"E��!�=4e�%+	Y�i@a�E�'0��@U�H�2��Y�'� <��𙟌"��ǸK���jW���؄�"a'4��$��.3*%���6:]@XSUF4 ����4�J�H��h����ay)դ["�[rŘ��8�R#ˤ�<Y��!�<s��V�	A"��pC��@��y�!%T�AP*��5F9dDY�ēj��U�']6t8:�LJ K��'�t:3��`V�3Q��
�ɂ7��J|�`{E:5����<<CvC䉽FH�@��X'Ny�A�Q�����h2��94��t���	�]%H����0�3�dȅ_�Y:'�)�|I�k��
!��O5������([V4[g��6��S凕i騉A�mU�5f8:d�'7be6��<����߅����˓9Ѐ�'�K�K�Zx{3�V�,$�7�ܢi,�D����d��u"O�q�C&�1j1TIң�k;��C�|��,+�"�A�z�B���	pɂ�N_��ܸ3b�η� X��'��U��I���l�
"z�ܴ ��b6����S��M3s*��J
�y��GP�w�(���	Md�<�Ei[$e�鰑�C)q�1�q*�vy��VN%HŇ�!9��{�*�)�2�Pa�,��C�I�1�\�o�'fX"x*+��R�dC�	4e�:�e�f 6q��'�FC�I-�<)���D1��*��{pBC�)� T�X��-���j�p4�,�E"ON����o��� $Č���q�"O��hB'��E&���(��dZ�"O\�����7��#q(F�(��	y�"O%��)�Qܔ| �� ����h�"O�ES*+U�5�-�J��p�"O(���gHr��@���چ2*�Q"O`��iOUH�����綼I�"O���	az��
�J���=��"O�	"��5�lQ�D�׬\��V"O��(��h�h���+�,zQ"O��2&]�`��V�(ۈl�D"O�4�!.69�2|�0��2F��M v"OV`*GG�rD��c����J��u"O �2�f�+�
q�f�ݱ=�vd�"Onт�	y�,x��^_؈x�"O��s�N�}�>���I�����"O�q�.��{�4� T���y#���"O֕�FC�*CܔR"�)C<m"O����xt��
��l���T"O�h��Q�A(R���#�.���#"O4�战el4���&_��,ig"O�Y�V�]r�Xz���4n��tt"O|�� YS���u�2$�&�3�"O�e�ĩ݂��`3�*W�^a��"O�P�l� ee��
��� К4"Oz9hR���xwdXx!/S�2�z��"O`�ʹ-Fn���ݖJ��z�"O�R�J�6��Mc&�I�@�T�E"O����#j�m�b�Z/�r���"O�9��L�lmµ�T�(G�z�"O� KǠG�2��3��*4�H�Z@"O�лe%��J��xP���
!�(+�"O�q��I;6l(��?F�a��'#RS�KR�F��Coȯu�=�'W�B�X6J*(����%l���	�'� ��ѣA�����F�>c��Q+	�'	��z�-�~��ېǈ�i0�H�'
�*���Z���Ʌ&yߠ���'Ղ`�MY'"d�HpL�]Kȕ��'f*��GE�&(���F�"�X�'s&���d�j�<�G���DC�a
�'�.�J��B/ub Eඨ�ID�p��'�Թ��mϑ(L��ACC�A-!�'N��b$�K�o~����x 
�'�2D
�F(��4(!"Ⱥ�ؤ�	�'����m�8��J �Ѵ�@�)
�'r�9� �M3p��K�h�	�'x�(��i͢h�bE�W5v0�	�'2�ᡱ�_�G��ɨ�'^Rs����'�%;�N�*j"�����K�j�
�'�$��"�'��Yp��yl8�nT?H�f�S
�p��a�/O�) vj�<`��A:�N�4<xp9(r"Op墲L�iDق���v9���#�L�F����"P{��x�R�w��
���y��]4����/�p�>�r�<��e���s�d!���
"�PD� �
=͎T0��.D�4�qBҔO�p #�`C��*��ɖK�P��ɥr�X�-R*l"��з�Ʃn]�B�	l�H�(UFҸ'�v��&+C�pB䉤V�ڈ�@̜)��m��$@1K<B�ɷz�Z�XVfPB~eaTe^��C�Ɏ{�t�J3��y�cH�&��C�I.QҬH�g��h9P��p�A"w~C�)� n�(�.��Nw�́�IG.����0"O�rl��}렀�P(נ%��	�P"O�sO�$�*��UM]�&�4X�"O̼ztg�[
 �s̝ U� �"O�-��4_Cy��A�x�$<�"OnU2���X�`%�U�Cr�eb�"O�}(ᬍ�mR`�2�X�XT^�a�"Ob��r�A �-�@n_�QbŚr"Oʕ��C8Y��JӦ� WlѨ�"O�M�U��E�T�Ƥ<�Xmb�"O@e����}��l��Ňrߞ��"O
A���X�P�D��2&��h۴"O�	��g@M��ѻ5�R�ۅ"O��Ap��#$��鈖�S?V�~��Q"O��á�E�w�@��e/ �n3�Y��"O��j��/��zs�R�{!:\�"O:h3C(��#D2�9��X<x(��"O��A"_�Q�Z��5
��i�"O��*��FWr�\ZR�9n�0w"OZ�3g#��:��a	��M�0��"Ol(��a\�X��!�n�*m�Fu�t"O� �AX�imt��W�T9�С2"O�lQ0�(�K�Z
]7H��"O� ��]�H`-roͺR Iٔ"O��)��>���σe� @��"O��@T��i90�Y�U�7�(e{T"O��+�eM�@�h��P�W�Z��js"O$]�3�ބ/ �����,��<˱"O�0谆��8��1�	A�[��ٛ"O����&�k3�Bq!����0"O��1���2ET %&��^	�`"O���U⚽ �Bt)p%
-ָ$�"O��B2��*�H����ini��"O����蚀��YÃ�Qhj\5"Oz�9�l�)-������)BB�	�g"OV(�`M�es�I+ԩǢB
�pq�"O��s�X�@&��J?\aG"O.СF�_�ISh�5yM��+"O�E��HOZE�5�0c@hA5"O@��ԩW8���1�5v50��A"Ox�Pe.�~���⋤v�X��2"O����N_�R���@M�_p����"O�< F��%K~4��B�(�FP�"O���êP�Ml)arJO"c����"On���_�y�hL�u��7�n��Q"O �G�Rg��c�W-c�h�b"O��@J#������%`���a�"O ���C<h2B�����"O��S�e�(��đ/�dd�ya"O,��Q�Y$:1j��؀c�"O�8{dG f��P���	��Q@s"O��`���y,= *	����"Oب*t�E�(���V)����*�"O0��.�~d��H�Y�ֽp�"O�p�jT�"�Tj��ۗ=�lY� "O�����=KPL�P�'L �<q�w"O�a��*�e��8��ʱ?Yl�5"O�=ä��.n���Ī��)�q�e"O:��%$u�Hz��Y�!�Rqb7"O��{�d����H�I��p5�7"O╂�b��"��a���K�w/d�QA"OE
�̈́�oU��%nD7)��"O:5�
ˣ-�%��� �:~�s"O$���Mo��RS,ſ~��&"O� �H�#�<�B�t͎!x�<�"O��8�݃S��J�P�xp��Z�"O�P�L���1ɛ�0WҘx"OD��͙)}3���q3V0��"O$�3 �ؿv�^h(���La�Q"Oک(TG�V�Z(�M�!�)`"O"�C�.�'B�&��fA�m�H܊e"O�ɱ�mWp���UF�.��A�B"OD�s ��)c��u� ?����"OL�d��(L���֋�yjPhz1"OL�R ��;tRL+�ʘ�{^�1:g"OzA����:�\�Z�J�/@�\�"O��3�$��*����îO���a�"O�I�,��ejД����_�^�*�"OĽ�R'�|}�(��B���"O|� ��� �R��g��Ef24�%"Oԁ D�_{�C%�K�dN¸��"Oę@�萡M�ڝ`CN$T2:qkP"O,�YP�#L���ȋBA�09w"O"��LQ�W}t�;�FG�rP��"O�50WdU�x�ZX�`h�&m�(\S�"O^yy a��l�xd����s�����IAX�
��ۅ-��pc��T@���3�'D�`�C �!N�	#VI��{6I�'�8D��@���GmV��)܆S�]�4D��:Q�c���cR+ų�XZQ�>D�`Za��7	]V�8�����u��8D��� V0S���#�(ջ=w�]��2D��Y�'٩RGĀ����s^��'/D��q�ܢ#d��pA'�,
B`Z�,D�lb�P�n(�jfC� H�
<Y�5D�b i��cM8�Bc�ɤ""�p�m/D�(���P�^}	ԉF��ޤ��A:D���æX)�1�ↆ�t��a+D�,����~킭�6�(qW@�jb*D�Pq"�X/@:DO�� cDEK�&D��Z�dñX������R���k(D�p�DL�f����ڸ{�@���*!D�0��͎aN�|qt �D� Ƀ��;D�d#�Θ-� `�}0�[�	=D�\"t킍[Z©��W5`�(s���>	��Z3P@�m��Ι��@\����B~���+�ZZ��	�D?Dʢ���y�.
�|���S��;:�҄��Ý(�y"ʖ�2�
�� >�(����y�"2:D ���&=�l��aW�y�Zh6uҕ��"����U%��y�e���A#K�hv�xO	�y��Z�G�D)�LT���WhW�yB��FTLP�ee��* if�7�y���\�ʨ��)0g@�Rn��yrG��nK�MŌ)R��m��'���yB鐌(�,p�ЁY�B���8�J�y2-0�
��`%9a�H�%���y��'d�@�k]vX�Q�a�&��j
�'g��p�E��(��9�Qh��[�=B
�'CT���KɟD7����B���HI�	�'B�(#���!���
S��6b��	�'��I �q�Up�@>"ܜ\��'��q �(��Й4�1-F�i�'�ԅ[�d�'g2����3q��r
�'*��z0�ӳ�\*��<]��X
�'�0��7dՒ/��ݚs!ďJ1(y	�'�����	��L�Q#R�Z4���"O� ,�d,�	b��Q�3=���  "Oݘ�
��T��=�� ���%"O��@�'Hf�8 �@�����"O�ؑ�˙"?�����T�9�D�Xb"O���OR�����C�A q��D��"O�4��Cر-��};U��<~��<C5"O)�B�X�l��ZЂ����tq�"O�X�5m�TG���Ā�"O�1YT�ٞ��!�Y�T�C�A��yB��eL>�bTc@<`���-��y�*ğ?��, bHY�.��0m���y� )�Z����ff��r���y��F�.�@a��[	�0Wo��y�A	4K�����gL�[5��y�)V&M�B�d $ub��y�	X�A꜈�MR�OB:e��dL/�y�$[4.���j�<H��șB)���yBB[Up�ex�"��C.�PI�'���y�W�v��} J�6���i'�Z��y}�
lZ�˙%F��D�k��y��^�zU� ����?}n*���2�y���+p���Q��H0/9�a@�y��P�$� ��5/�5*4�ϙ�y"Ʉ�xR�R냩zq2��N���y���H����+u�mS&�yb�Α)!�V䖓\dx����y"�/e�ީ(��'U��(����yRm�"�Y�	X�D��-��'�*�yRA��*�X����K���ȃ��y2e�%�j�����*3�H�>ѴB��b�f�Ckύ-��sf�.�B�:V���u-ӟe��H�DB%
'�B��SmB�;2aT�hz\#DյepB��,}����C��}r4�"-ӆ*�:B䉄,J|�2��4E0d�h�;0B�I%R�	s��.3\�х��C䉏^VJ����%lRL+�V5%֦C�	�N�B�M=oTM�S�H��C�I�K��E����O@�� �.8C�IB��]{��{
x��B�ąS�^B�	8�.�K�'g�"}�"U�3bC�I�I"Ȥ���K�}3�Dd��#G�TC��,Bw�%d ,~�����ѕ`OBC�	�3|䝲Qc[�C����O�1�NC��0B@("3�
���P�¶q�PC�	8=��p�@��i��)�e@�K
���ȓ=�؍����:��,�wI��7K �'ў�|�K�9�v���$J�@��Ѐ L�v�<	Q��gFh�P�ɔ~@L�'ap�<ӆ6:R`
BBS:W�Nm�ȋR�<��� K@��r60OD�!f��%��x��C�!N.����<^��ӭ���y *�`�gI�U�ܹcÅ�y��G�KW`)�&��"�Ha�i���yB��aJx�������� �,�yb�8\~�H8�&\����B��S5�y�F"ʤ����Ƞ�-9�y��6{5��A��U�~��(C nR�y����30`v)�K^���J��y�M�w��Mxg�9Ԩ�S��]&�y2B8t��ك�\>���	�Y��yo�&D>��l
1<zRQȖ�C��y��8}�Ne��N̚<��lbƂ���yÄ�L՞��2&�-��Yɥ�:�y
� �t��M����Pf}��EAc"OqWf8/��Y����5\��H�v"O�x�tB������:��v"ON9+# ��'v��j H��H�zA�&"O����&>'�m
G'�
��8�"Oܬ���\<<�	�/O%�����"O�� �P�8�����oȺs���y�"O� `�0S��@�哺i���K"Oň�Ί�"¸$����t+��8C"O��Ś�W2H�;`�Q�m8X�"Ovȸ�aB�-��]	���?gt�q!"OVMc4O	2D"i����u]X�g"Oj� ���>�����cx���"O�sjٷ	^�;gŊ&E��3f"OqXv��K��i�a+^�&UεA�"O<�!@�\��L�p8�|�"O,{�M3d��{�
1Z���"OB� *J�1/�Q�T*�Bk�2V"OdJ�+��A
��y�Ɂ4\T���"O��'ID&Se����!R*�+�"O�Myg�Rq���s�P�]H�"OdD��Цl����gV>K���)"OhXcε�esv�ŏ � y�"O*�`�JM�!��&�t�2p"O�i{a�
,���A�$�I��JQ"O4��!�:�v$KE�:��I�"O
 	v��%W�4�ؠD�-�� A7"O,��W�ؠbi�����?�0@�"O������5��8uG�m��z@"O�Xc��T:_Ä�Q�L;8`�U:�"O8%�1h���tX�^<Vs��"O�<��c;�,u�r�@	jPR"O�d �	%�z���˟GS"�8�"O��@5dS5&˶! �B-wA�H�"O�����q}��	��$*R��D"O &�Y�k�4A�S.�N��p1"O���8��u�/
�H�"O"1�Rϑ�N�l80���/�i��"O�l�D��ZX�mN�Z ��@�"O��Bf�Խ���X���^ )�"O��(�*ԅ ��,U-���Y�"O����6p�Yː!exw"O����A��OA�gdF�����"O ��֠�#HZ�p@�7��Ũ"OA�Ä�-����H��z�Ȁ�1"OjH���'t�8����*6Lyq"O����[��	A�A��0��"O��TmV#�D9���]�<�z6"O�q����r��07�y�^ P"O��؂n�)��q#�U'"OT�����VE�!�'��fA�pj�"O��x�T)�T�,�4{0�@r�"O�i�#��6�n}`#D�--(�@"Ov���$o��z�#��(�Б+�"OJe��aB��݃�A
�����w"O�$Y���/��%��w%:@�w"ODؙ$	�*�tX��v��� "O��Y�a_��2)�٧+����"O��ɷ���Q��l�}�℈�"O�lBs��$y!�ԓ��7u"��u"OL|QE�"�E���� j��U"O�� е31�9�ԅ��k_��z"Op��Ck�:��D�#�R6(EH{�"O�a�Ǆ4��,S��>`2(�zr"O� ��#g"ڵ^�\��C4\�ő�"O<)�Q��'�v���AC ���Kw"O�4b��W$1'�0����*-��dC�"OP����|^����垽<4�P@�"O����ћ���T���}'����"O�)#�aJ�6T�(h�A�;)DH�b"O��Wf�K�d
t�ׇ>%.]��"O���ei�b�"ԓ�()
2| E"O�m�4ĈF	����(�9�굡�"O�����
Z�$`s�aZ�B���P�"O|t�DG	JmX�3� F�t��4�"O�$S �̻N�x��c.C�y��9�"OB�16��GB���K'^b�9�"O�����3eE�ha��Hd"O*%8��̂4(p�w�E�bU��"O��9�e����HJA�ߖj�8��"O��x�	stn���!�.��k"O�eC���F^�� ��U x��["O0y[��E6-2X�U��]�|	�"O�q(��F��a�Ä"IZ^���"Ot :b��U�
�?V�}��#Qo�<yc㔼t�$���;Z!��E�n�<���/Cg\��5�H4 �8�)1l[c�<	'�ˋ��`��3E?|��g��[�<���=<�r]�&f��c�B��ʈM�<	��@��Qh�DP�@|�)��NA�<#N��Zwi٩`����OU�<Q��߫
5v݈0��)gX{�-�P�<��
S���j�LG�
i��Bc��M�<�e�ԣ�`@��\�-�hl��/N~�<�r�J�!�z��2�M�kҖ|�R�Q�<����J�P�o٠>�P��M�<Y5m���׃��(p���m�<QS���(a�afԱse^�ۇ��S�<I��@V���甯oq��۷
�E�<i�ʜ?xX����� �i��@x�<���Z�m����揟1gn�q�2�p�<�1����}�Lͪ_]|�ygD�B�<IPL�;O�p2��.�|q�"X�<�$ �к��2��/�
ݚ-�|�<�V�J*;N�xT�[/`,Z)�eoS�<��*�
}��x�D� Ψ0R�)�F�<Y��
|B���"�t~�Y��LX�<��h�'h@!@��d&.l���KQ�<���K�fĎ��$d��F �K�`I�<��d��@Iژp���;sz"q��k�<�Ā� `���PRn�4` �m�0�L@�<!��*F��X�@��P��3��y�<��˛�j�6�����h����x�<�Ո;}�����R�q
^<z�ʕx�<��M�(���h�/X�I>�����v�<a�&��d�r��t%��8��*���u�<1� ��3WԲ�n����亰@�p�<�#!J�b�!�+�b�B�j�<��oķUi� r�'�>��QP�A�<� �ýL��� 2��S4��YӥT}�<a �53�zx�`�P�?ݢ��ƞ}�<i&�ǰCX�����l����Fe�<qc���Sm�K"*�� �.!�V��w�<�c&°q�*��N�!���i��t�<���";�>)5fG��	@��U�<�Dk���L�����euF���g�<���X�#�m`�*Փ	�t���z�<��ǆ<5�-���>p6�*#LSq�<� ��Pa�'�~����B�u��ٺt"O��0��Ԧ;��+Ae�-D>Rbq"OL§`S/uRX�eP�2����"O ���<u�*�c��_n�2��"O@qb�K�M�I��M�~q,��T"O���oҞr)�dx��).��Ra"OnM�b�7�T5Q�n+�vyx"O����,���	���yT"O����OUT�YL� E{�yXb"OXX!G)T�����+_h�Cp"OP �@��'�#W Y6A��"O����"�pғ̖6~�]�$"O�0�L��F*F�q�+�K�*�{"O��"���*��W�7��Tyg"O$}22f3k\�Q6LC�X���$"O쉐�i���2c�[�lP�"O�����F%v��#%.8�1X""O�̊�@�!sSl\�G*�/���s"O|�B�5l���q���{�i�"O�x3`�])N`�5���[;,�SC"O�X�l	8M��Ĩl�	8���YP"Of `D�>	
 !��Y>��4�"O�9���]24]�-����,��"O�� 
�!cXb��|���R"O6�G��7�L|��O �J0FѺ�"O��Q�H2�̝B��O�TN	ї"O��(���9XF�P�Ϳ[ۖ"O�I�X�s*����O�X�z1��"O:娚�;� ��D_��z3"O�}��F��&�A�dEܶzD=
"ODu� DB�C�	z"yԲ��"O\3w��*:k~4�4JS~ŀ�s'"O2�"�gK��&��2IH5x7"OfݪU�ѵy���h0�F�z�"OڍS���e�  ��A�z4�I�"O,�0��X2��P>��B"Ođ�Q6]�,��V�Ƙ
	^��"On@�"�4�,=is%��6�@`"O��îL�q���`t�6S�ā��"O:�!��+[6~�qR+8� �1"O�5�b�#u
1Q�Ȏ�o����"OhQj�/ڂaި��R���"O
l9PcS�S ��X�FB�wwP��T"O$x0�e��D:x��̏,s�$R�"O�x&�U��lX�Cʹ�P�:�"O�m��#�'p-�U�ĉ�7�8$��"Od�sBB ~Ѣ���P2�~9`F"O������0:jz$JD(��w�"O�ҨD�FHD�M.�9h�"ON�*�/��Svq�K�:W!�!r#"O~�h�gO�WBl���锉j���S"O���L��Q�ʡF>[㚸�6"O�E�@Y8������X$tј�"O| �0(�(#�м�� D�&�r I$"O-�C�/	ߜm�ŀ[>f��5�"O��01�7p�JT�_���0�"O>��k��'E�A!g.	�'�$ h�"O����nؙb� ���m[�% ���""O��!�c�#8�@IZ��M�g�]I�"O�}ZW���ֱE��
X=�q"O|������� )�e�#�
P�"O�x�ajJ.HI{d��D�"O���Ѥ��3HP�9��5��"Oʴ ��B�LDJq@V'�/cs��"O�  ic&��L���1��;(m���"O���$@�´�w䟨r�4��"O�a���tP:&-۽*R 	)�"O�A1�N�Jl��`QK
��(�"O���6KE��ۅ�Թ8�
�h�"Oh)��W�$�P;�N T����"O�Y���.\��kA���T��"O���E ɘ ���W��a�-j�'�1On�����C�PI��g|\+�Z���	_�Ț ��{�y�B���'Ѵ�:` (D��	��2D瘼!��5?��b��'�D'�Sܧx.X���%^�\�Z����8.�tńȓB�-s�F=#�zZLC��m�<�s��AvHI�)^�T�� ��N�c�<����K�DA�q��E�$�RR�cx��GxR�͋
 �`/��&�z����/��:�S�DmGTOt��Ӂ2(,܉��P^�<!E�Sj�\�{VDX�MO(�"��~�	��x��c����dĻ:�L�G�]�`�#��$c!��I��)��o�16� �ㅲP�!򄗸�Y#�%2"v�=�v�A�T�!�A+U�p+�&VV����L
3{!�	Q�l�zA�wPrC�둞m�Oj˓����pDB^�v�$����d��"O�˥��=g�����ս*$��'�Iş��?�}�r�^�1"*��a�dj�2DJ�L�<w���l���.،(����i�L�<a#`�/k�6�aE@Q�rJ��²��a�<���?f�̱V�Y&-@����`�<Q�n�GAvh��!� %o���t��R�'Ma�d(M�.��52��CP"5���ɭ�yB�:�d�zD�N�;�rqi�� �y�T�3���*v��,���ᦋ �y�
�r�ZQ��T*Ċ)�5H��yR�_()��IK�a˗�W��y�	ν}� Q�2	�	�t9��]	�yBʤ@'���a"
��@�Q�֗�y��W5���uR� uA����5�O���*�!``�D���#���"Oz��Ud�4��lA5�O�6�v���"O�M"��τC�R���N!"֚���"O<��'��;Bjt�q�C�nV� ��"O|�p��ӧl���ؗ͏3����"O�E�ޝL7���̔�4�~���"OtHQR�+?e|E����w��}I��':��p��B���+P���PG�ֲl���0'>D�ܚƭ_#^��p��dV]��T���:D�LH�NVp*bIG	g���0�`<D�Hx�[O�TrV�ĘM�2�%B9D�������u�@s�'�Ep�J
6D��{'@X$ 3������{���d�!4�0c�k�['�Y�GLםq�,D�"�Y�	Y����D%F�j<�e�߻ .�<IQ�)D���A��k��Y�G�]lN���(D�t���)k��� ހ�xD	%D��1��ҷ^�̅Q��ܲ
r����!D� *w��#l����!Ł1㬵S�.=D����J#S>�xA(��=w����9�O����n�ܹa��
<V:�P'i
=j$�d�<����	�S-�Ec�aB?P��e"��6-!�dѻb�jE�rDO�U�`�2a�H!��L�P� L�z�س��֒!���5\�R�ɐ�ɾc��蝷!��>Nh��rW�"J�Z���.9V!�� .�pbNp-f�����D���'���4��Ȅ.@�@��GBd*y���OTB�ɔ-[N]x�㛌q~P���ywB�	�u|��"���O�6P�鍄z|�C�9G�`L�b�2�ݪSC%x��C䉫m�h:�^�ĕ��∍d�B��*M���@�A�|߶�*T`��?o�B�5,���Q�
��=�'�E�B��B�I�-sHٲ��*��P��eW*\�C�I�y�6�;��5`״�s5�U�<C�I�A�\��a'\M�2��,mbB䉃"�J�A�Shl��>��B��\��#�D�@�H�*Z�s �C䉏L��x��JP	�@���X���C�I�|X��"ֶ�Zp��W�]`�B�9}	��Y���'�|-����fkC�I3!}����Q�pI��H�-�B�ɣA5��QAkЖD:���ŋO�B��;�y��C�|� �8��D���B�	6����X���id�U
[�B�	���� B��$�6�"+��C�	�^e��兊+�`�ĀԸ�"B�	�X�x�s�4W���bo�,��O��=�}�7d@�K�cѿ��]2P��X�<��^"L�|���aC�B�=rwG^S�<��/7���+�M��-��@��l�P�<�u-Ės	�(��2��d��J�H�<��-Q�MR¡2�,�*\=Z�7#DE�<1Ɓۂ?�I����5��)��@�<�E��Yt�8C܂0}�,��$��~�<Y��E��� pt*�s����|�<�2gQ�x��%�,ѥp<Ƥ#m�z�<!�
C>J����b��[b�<�b�3#��M����*�����T�<�#�@� ��Y?<�CRj�S�<A�mήD}�� ��m�\<����x�<!��>v��RET� �ԙ:{���]��k5GV�&�����g�R ���ȓ���xs��*{�t���9 ���l�]!&���a�α���J�[��X�ȓd�mׯ��[@�`y��5=*�������(��6S�T���+w���ȓH� �)l��H	���\ܾ����Je��`�4M�$��S�[�5	R��ȓ ʹ�h�މ	D��#aђU�	���l���a�X��ć�3z����ȓ;Z�I�$&Ȓ����_,&s:-�ȓOz�q��߾	(�	1��	�����m1���!�48���BR+
�1��C�ɲ-�85I�m�1�Z�+��74[rC�	�
H#�*�k�6��#GD-`S��$�2:�ȱ�#��>�U3Q@s�!��57�|�B�U�ڨQ����f�!�ǺC$�!��w�|�%c��W�!򄄊Mz.��u�9$R^�I�� �!����l<cQēG�r��b�J�!�ƖRis!� �M�"�[Ak�&j7!��ЁX��U'Gb�Z� W,��5!�d �N��^%j�T���3*�O~��d�'E�0�D�˔%�~�Z��ޤD�!�dR�%�ѳ���!y���c�_�!�d�F΅���.q������.�!��\p�8��9od���`���s�!�,#zthF�K������q�<� ��!/4��!�cP�R��:0"O�@�V�������>�p��|��)�Ӌw����]3'�9���A!6C�IXhը'#�.�p��g���}v�C�I/4����@	�c6�P�Ԉ2�C�	 U����"�:,$E0�i�3b�LC�	�!=t�� ȕ�\!�rsO�:snC�:C�yc��YE��y�hKD:�C䉿7���q��庐뉙a�����ɃZ(�;�\7H����+G(l�B�I"�m���7�y��GD�J��C�I<���"���B�u�Ъ��v�B�	�d)��*Z�r&���3)��C䉃K�"�1ц��m��	L'&�C�	=��s��6`���!�֕g�dC��6u�fxҎ$��(ҫ]��p�D(���ON�?�'^����6O��H��U�C@&$��'��8���JR�U�e螨,���P	�'�D��K�"�v����#J�	�	�'�>����@-!��A4@۹c��ȇ�3�ʥ�KJ�v�=��"X*Q�����?/��1�.8:��B����=��S`����O$�D����ޗ�$�|��I�b�@Y�G�� h8\@s��ׄ?>�C䉃'���Q1�H�3�٣0�U (C�9 ��i�5IX�U��R���)5C�B�(�.���T�r_���v�S�JS�B�f��vm��/�NeK�,�?_�B�ɜs�8%s1c�V}�R���VB�	�x�T8�7�G8&��)DX-H�C�I�	�B�����@�m���CL�C�I�X� pYъ�fȼ��!J�B�I� �z�b��C�m���i0�ވvB�B�00�T���&��Un��넭�8�^B�ɇ4��X0���"_B<�B��=�0B䉠|�pQ�5~��8*��\B�ɫ_'J�DK{b0q�0� i�B�	$l���L�}l���L^��C�	�&��2��ٍ$p@�\�,B�	�-n�i����~����([(&jB��?�و�H�)��Pɣ�Ʀ5�0C� ���Z�iA��T���I�C�)D�LP���G(e��jާ(��C�ɱ_!te� �L�I3��� [���B䉱t8Z��D�Nlqփ�80��B�	9����Ɨ�}�����;G�HC� �<Bg)��[�� �+�� w:C�	��%q1��7R9�TB��U=*�C�w�d<�EƝr	°SSbRP����-�p�D!��( U v�@͌�N���ȓ;zV�3����DɞI0�CFj�^�ȓ>��v ��UNi��0j�4Єȓd�$;rL�a���G��	���ȓ�d�[:[XYj�!�'3�d���		DL�2md���`��{;b|�ȓ:s�-��`�z���1��|�
��?I���� a�V�ZQ��KB���E�n|ў��ᓊa����&��\���5`C�\l
B�Ɇ	�*�B��$��|ң����C�/[x̠W���pG����KG"a��C䉭;^��'���r�IH��-|K�B�/V��u@S��PU��#F"M �B䉒O�4�Y��S�1x��J���O<�=�����U'��e)��	�p����K�,Y�!�� D��s-K���X7��%F��u�"O�(�h�(����e���Y�,"Oҽ1ϝ%v d9���/v��tR5"O�hq$$��* W�?�PYu"Oh	�e\�|��A@M^	
�� ��"O6-*c�A]L�yC�+O<R�(#'"Ox�@�M�.Մ��sQ���"O~�S7/\��@�$�AE����"O XӍ�5��y2���sD��D"O�,�'�\%Ӗ����X�,���"OޠiBo�:M��R푩)�R�"O:{��Q
�;�,�6uFLj"Od!R�K�_��l�q��6�PyR"O�Q�p��\�(E����4/�d�"O<Yɶ#�2~ �Q���'"O�p���i_ڑ�8u�R���"O����O"u�`	4̊&.��"O|�C�j�����+�R��2"O����UcWR�!�n�QȎ�1O�b�#�y�Bp�+�;bu�Mc��O~C�	�{iR�h�ꏫ�����g� >kFB�I��rTs�� c�*DxBc�C�	r��H�1*L9�oĆA�B�	/l����c�@��IY�I��f\XC�g���$��
I��[@@O�*C�I�(��cQ]K�Iv�ߚ(�B�		}��ɪ�D�P�J�y%�[=q."q��*!`�8S�Ã9�����'��/q@���=���像;y܌����}��Ѕ�I�&��d��:YR8�����
4�H��=���s�x�"��0���䥆�?hLtQ���64B�:�LY�p�t��ȓ�䨊�AG3>��E��W	�A�Ɠ@(���H3'b};��ڧ0
���xҋE�e��v�Ɨcr�	Q j��y�G5W:��!O^$G��9�GP��y��K����sH<�� �ڃ�yR��>=� ����44:$��C]��y�$W��|pǤ�>Czf�L4�y,ǉ%2(��-]g����Eć�y��߲>qR��iX)r��� �E� �y��I#Eu��{�Γ�hz��T���y���j��Gr������yjD�gO��q���cϨ=ʷ�O��y�DN�����nBJ�f��UDS�y2oW��z�����y��h���y��9I!J]Y%��p�X��V��ybC �|�Zdr�iP7g�n}�a���y�'��r$H�M@�W�}x� �y���i�1Z�-_�}θ`����y�NE�xԜ��7��^�V�<m4C�Ie��a���.d�q��Y*C䉏8F�%b����NuQ񅗹zy0C�����2	I$����2d7R���3?�s�^.(�R��w��V��mra
^M�<9`*�0HiBåT�E� ��O�]�<)mM�'2�iA�H�eD,�Q��]�<A�b��@������>OJ��t��T�<��Ùjd 
�d��B�(Ԙ珝T�<$��G&pA2���LH��`уE�<1�@���}�Q7|�)�F�	vx�̔'a½X����&U��(�-�1[v|
�"OKٲB&��тh�lV�$k�C�	�'[p���o��m�ve�΂Y�B�)� �� ��>Sx��e�N_x�("O$\�w \$2x\ջ��_��ʄ"O���#�&��\�v̜�U�>�җ"OT��EX�-��ۅ韤���PT�'�1O��s�NH�v�^Q���
B��:�"O
Dj�@�\�:6d��dO(��"O�YW�,���4��064�C"OF���.'m����CV�G��!@B"O��P j�1�.L �6���2�"O�)�$�&��]�f�e����"O�e`Z�k�~�`�n8l�P"O�Q��UCf���e��ai(`�"O �E��]���&db�5��"O0�Y5�ې|h:��!�9N�0XQ"O$Ę@����Qb�R�F����"O��j\�t�ʨ����0є��"O؁�D��+^S�@�v+�&�L�7"OP��.��Rk7�x�"OL��0D�rr�$Cp+\�h�"Ohؓ�
�Z�R�"װQ#l![$"Ox�P�%��%愡@�D>>t2q�v"O��`�b(y�� BVm���"Oj����!:��P��˴L�^�S"Ot-����2�����f/L����"Oh�[$�	m�%�)Zx$"W"O�2��	:6q04q��"Yӎ	+�"O$'#�­�$�=8�V�h�"O���P�	�[��l��^:�P�3�"O��dE
^�L"%D�G�<��"O"L�4-�j�*Y�$�a9�c"O&�2�ŵYfPpp%�D&K&Ӆ"O:L#"����*���S�!�6�	�"OZ�r�kZh�H�"���"On��(BP���*Q��Q@"ON�BebU�@�1qfƑ5��H�"O�I�d��Y�TI�%G�V*���"O��c���s����f�z��"OD�!#.Ж#�H�O^�ks��)�"O�}�E��=�(U���O:ٰ�"O��:w��(�z��V���
�
V�'R!�Ĝ-r��� w	��VD=!�M %!�
�k���ڷ	�0m�ΐqbmR!򄋽�V5J� u�ab�a
�
"!�$T�K���ұ+�+X�(�����!�DOk'��DK�7�$�б��Py"�Ĳ� �kVϔ0\����fӈ��x2@ۻ���W�= 
�'D�cJ��'qa~�_F��Q0�S�h2�QVDO=�y2��a�*��땨YɆ�U�	�y�������F2e��P�wb^�y�K�33��ir"]5j�@x	c���y2NӀ�r���I@
-D��Iu�%�y2'�"��`�,�)n�8�I��5�y��4)*�Y!M��<�����S;���"�O�趭�A7�Y��E�3���*U"O\��$��_!��vdݲ�(�ؒ"O����e�b�ˣ��2h}�q��"O��zF⟡3l� \�lq��kܡ�y"J�;ϰ}��V�HBa�F�T��yB�йQ��p�"�ogBI���8�y��Ll�`	�c#8� �^2�y"��E���
'��%`�"�yrIד+��i���i�^\�ĉ�"�y�nD�TΞ8+�M�26D�8t���y
� ��
�/�?O  #��NPJ�Y�"O��Y�)�����#�
��kg�T��O�Y����F�ʜ,h�p��o>��8�O�B���b ���aP�_� �u"Ob �a��ы6"��+���!d"O�;g�
	VI�#[�7��M�"O�a(wN�ep��'ㆋA�@�"O@�ZUG�OK�AA����af"Oʐ؂a+ Z4{0�(�h�c��Io�'��`�$���K�k�!i庵IY��!�$ؗ8`64�GdW�kT0�V�\j!�D�6zP�G"�rh�YȰ �i_����%,��9�׃�.SI�`�N>V���$�O����@�x�hyc��	,����&�!�Dك�� ��C�I�B�Y�ڱf�!�䚚(�\ZBY�����b횶K��O��=	��y���'�rp{��5t� �G���y��\*p��yv�ƍmKfɹ,��yҪ�2a�� ���Q��"դE-�y�a
�w��=���Jmp��q�� �?��',��*c�D�h6��Sa� -�Q�	�'E�\���<�4I��.�`�	�'��{RZ�[$⠪BZ�dg���'vɫG���,qcn�k�q�'��˲GD�k���%`C1�="�'�r���R�_;��6��'Xz��
�'خ���*��(=��mI�3^̜z	�'˼X�!k�AG<e(�0_��8K�'Æ� E��F�Rp�e��T�~���'S8�cC�1Tֈ��iİ��!�'�`�۶F^�3O�]�%I�&8������`T����j^Vs �3�y2�\D��BfEU���2L��y��	fs�8  � �^��� �'I�y�F9����1��k-$�p5����y"&	I���m#l}KV.��y�����t��D��%�R�#��x��zz$�����'~$	c���,Z�!�d�oJ�B"�΍Iؑ1�-|!�^r@�
^:F���r �X�e!�DO5'$Գ1��70����*Y�!�䊎y�@��Uk�3I�ŋ`�O* �!��
l�� ���0�,e "#N'I�!�D��M���`�i�;�H�Ѣ���!��=&
�0`�L8;ɤ�K��%�!�dj��e�D���ލ05o�/�!��)nj����K8p�l؁`N��G�!�dG�"�~|Z1.��c�VM	(F;�!���{ ����iVC�p% ևYR�!���7�D��lɸ51���F�g�!��^�@�Q-�)%��6Fy��O����F�#��9a4!�3p���R���%v!�\�N��l����6�@)r�BW)t_!�d^�$��7�c�.��p!�4v^!�D�C�L�jkB�{��|kEg�DP!�Q�/����劑9��H�o�%0�!�\�l%gfPA��-Ӣ� ��!�D�+�챣Vh�%��D��k�N�B�'��O?�g�{h"ar&�y���J��l�<)V�T; ڼ�w�_9X����hGk�<�ac2Nٮ0��#�2J�|!��,^�<YE��G/Ε��k�|���2��[�<	p�������6B���1c�l�<9q���_��a�E�1'�0P�bM�j�<� �%��S'>� (��ʂr�6h��_��G{��3Y��e�� 3|�1xq��6M!���ub�Ai�NN�Os��ФbO�P�!�dE�>�PU1��-B�Ƞ#'Ď�z��w��10�CP3 ����Fn�Y��4�h7m��yy~BG�8$���w���8F��5]φ�iV�Ƕk����D��YE�ģ?����PI�6Jm��E{�'��Ŗi�Bl�-��K��Ua�.�!�$ͅȓ��M�p�ӌ,
`9�R��x��=>���,E�=B��A�8�����23��&h#�Xۆ(�L_���m���׋�A�i���t�XЅ�=}�9�qFS���`�
�-�}��j��T�Hב�����f�%3��E��I^yr���q�0oGZ
�;e���7".D���R�ԣ�.=�7N	*���(-D��3��V-I�u�eS��4�W�7ړ�0<	�nK"^�ܨ��e�W�Ɣ���CN�<Ŋ�����Q ��-��q{@�K�<Y�O�8$��!&�3���R�_H�<�fG:e޵�ׂ_�^�>�:�˓^����}~2ŋ�fҠ���V�ƞ���☋�y�֙i���2�D�-_:�<YW�9�y��8|���(X'\~�\#2��y�������h���3��m�4�դ�yB�Ď��] 1�
J�m�ED��yBjH�\�4hX2J�Y4���cZ�yb
�@��M���>fX
c�#�6�yBL��(,����F��e�1����yr瞙Q��1���/�~��G"�y�B��k� �9�*U0~o��hR��y�'�]������ph�bG���y�ဟ"h����޲gf����3�y2ʃ�c�ވ��*��oKx\؆M��y��4l+�I�Y�n�з�Ƿ�yb���*�j+@��;X���@��y�(Y�gw�����*�p��@��y�����V�A1c?���I��y�߽�� g�^�Z�I��	��yrK\�YJ�!#b���SBL��i�+�yo�[�pP�ѽH����@��yR�L�jo&�A�1e��ۥ#C��ybX��N���յ+0JT��G���y�J��E �X$�#�f�z�@X��y�I2blP֮�&���	-�y�H��Q�a�c�P	�ԌQ]��y�E�::�T�W�SX��)ݜ�yb��8'� H�mT�I'�Q2Ŵ�yb؇m����b�'`�); ���y��!j�b�9�	գ�tșA���yr�_����Y��A z0��zf�]*�y�C��;L�����)q|� ���?�������8p �i� ��I�7��w�89�ȓp'�5`���J�b�a�jر ~��l����Ãʸ���w䛰$�D���Ib1�G�K�a��.y``�ȓ'�n ɓ��0�b��N�m�̇�fL���� 
	���q��#C�x�ȓbZAk�l��aMd�� hơ
F:�ȓ:s���V^��I���N�X�f���kx�dZ��֣R� h���jEZ���6�ԥ9E!$q' �2 �G8��@�$�#�,�h����a>RDU��S�? �(	d�^�"ʺE��m�&�hu"O�9vD5Y ��)�Q��	X�"O*}�D�.r��u��(S�NAI&"O����"�9.����*�&��!�%"O~!)���3�¹���۩v��b�"O�Y"�
[����%��(y����"O����)�C��i��GԪ:[�%�"OT�i&�ûm~YwG�n���H4"O�����м'�T�r��7i3HhH�"O -�h
�[,�����!�"O�2��J =�P��>8֡��2O>�A5gٓ�`�br(BLeB(��M< b��>8�~e�5a
33f�ȓ {aѱ@�v!����A�> ȮU�ȓ<?�����	o�搸�fӺ6{lY�ȓ����g�i��X�W�	�!��U��g�2�bB�5�F�8'\�7��`�ȓ�t1XQ#]��%!NX17����X���H�F�d#��1����r�ȓF�*9��m!!�ɜ+�Ɛ��`�P�)�2��1�cN�Q�\���\~�
-`�&�Ȃ�H�j�p��\
�y��M>	|�8%�ɑW�D-8����yҪ��z���SĂ�$���Ph���y�Ø�6㴥�$�A�"�T��'��y�ǂ%\^Z\�E��-Lu����-ӝ�y���Tڨ,�@���Zc�� �c4�y��?`a(E�7e�&C�rPQ�
����>I��?1�Eͫ3p�d�l�B�i���y2�-/��5�L6b�T�ER�yB҅I#lh!���?V��]�MP&�y�Q=vW��`�LЂM�>p҂��y"�GN���q���J�.IZ5`ږ�y����8�z��E;��hs���y�!�NK^��%iݐ2=0d�������>��O\���"^��a�jN�h��0�"O&l�Š�Q�D=hK��m)����"OD��feK�O��T#Ǫ�*?��2�"O� �����r��ܱ]��5"O��C�+��+_X�A�ŋ�@`���C"O�T��EC �T�򆥛AV�)��"O�uXciL�|�EZ�JS9�Y$"ON��ת�e�x���W;!��%"O
){�@�)(�n�ʔဣr���s"O����ʼ"!tx`�`�!^&���"Oh�J����"�x�cDoK>7%���"O� �6
ېY��!x%��#$ր�"Ory`�8x`d!�P/1�1�"Op�Sj]�zJtK �C3? ܀��"O����@�";��{ G�
�~�b�"Op�`��U'I�ń	%@fx��"O�����K]3:P�2�X�UU؍��"O�UҀ$��|T a1`"��Z*8�s"Of���L��O���qaCR��ؐq�"OH}(U�3{`P*V~\T��"O���c֗�h������K"O�TR���}�E#�oХ;�)�"O�-�b�вl�<����5֨��"O�	+���g��p�Ba�3"OP*�!�?<�f�1"h�(�h�H`"O,�"����e��,��8�(2�"OX;vcУv�JU�ˀt�>�i�"OT���ҩ[����w��'a����"OM�JVdx*��&��� ��\Ё"O� ��� �
\����(q]��"O\\�G$$r�9��ee~! 6"O�X�0JO�v�*�x �ǆ_W�f"OLl�C�<n�����Β#���b�"O��� �`���(���=�6}�"O�t��	��6-�"�!q�PMJ"O�83�#	�
�I��`:v( ��3"ObM3����mؖ��%���v+��!"O,��f��UY��Xt�P�Vn�0I�"O�S�-���|4hŮ=GC°�T"O6��Si�X�6M
��ȋN4�5�v"O�m12d���}�R'�Nd�g"O����n[7-�:,�,(M8�+P"OXTɐ�Xf�ib&`ͣ1�>�[�"O��R��J�@8��U�t��"OF�ɀbԐ �	�:.��A"O��Bȓ0�pT�&@�T�z�"O���	To,���n��`�y��"O4�(fhݕ_W�T�`�"6�pQ"O��t�q�T0�Ʀ��[R"O⌢��҅
��D��*���f��"O�D:��L	#L�!#�L׿r�}��"O���S��#'+��AdN�'�R�"O\� &k츀'N�M���Ȇ"O��3vAA �����n
4���"Ol5Y� �#z�����΄g��"O"���+�
d�L]�4IY�o�@ð"OȘP�
Ȣj�vd��H�/��0�"O��C"��5B� �n�p�"O$�����7C�mxC�"Om)c@�YT�b� 0>��3"O`l��B!$w���"ʑ��"O@�+�o�$%@<��R�4�u�"Od\�t	�b@td�B#Q�M���"OD��D��IN��hV�M�u�g�<�0������g�U"E���v.�F�<��fD3 B�Jr��#�N���W�<�����ja9���P1�`��T�<Y�#�Pf���G�o��1T@T�<Y�!Hj�D��,�
�V����Cz�<�s�D.%nMx�%Mwnܑ���n�<����(���.´0����`�j�<!E/U���9���4X�����!�h�<ٓ�")����gN/j�P�R|�<����:�0C�)/�J04Ex�<�ʾA�@J�喴9@��(�w�<Q��	H��U	c�X4�:0(�ew�<i�E�aD�=灏�p�&p��.�q�<y��<n���w##���@ �R�<�W�&�=2e�	��@�4�b�<y�e�)o�tX���!�P�|>B%�ȓ1���'Ȭ�R�����a�BɅȓ+^l���X�~ςp`��¤x�hp�ȓA�e�W��JrN}	�B� `c$m��U��0r����nD�ֆ�4O_ZX�ȓ�$�Qf �.BVDa�J�3qX}��Y2��j�;?B~Ey��I
�����鳴&͍D��T�Շ{Ip�� �Q@6�(&q�%:zu�ȓw6�<��J�f9vX��̒�&mDu�ȓrø�5,׆p�l�KǬH��a��$"�A�.�	��t��� _-�t��O����dS�3ߺ�ZV�:h\V��ȓ!��t`q]�"�*I�%�"t�n���S�? HHp-]#H�qqEO�k& qG"Odi��#�G`D�)IX�V�0��"Ob�G��	��	*�ϑ'El��&"Oʜsv,�p
-�4J�q7T}�$"O0�ن��\F�	�h˘d��a*Ox�VE�7���Z���E;�'.��PT(�9L�C�VG0% �'�" aӍ��"0��񂔭K�(���'�����R��0= `.F4��	�'������'�(�{�閸-yz�a�'S�(��	�Z��(��S$-$$��'��A��lG�S�T�eM� 1p���'Њ4�"�ΔP.z�A�#�R���'p���B���JW�s�-)�'���G��R��q�&m^Kmd�i�'�flZ�cΧ�*Q�e���@$b$��'�L��3�̻	zX��$Ӗ
���'����Қ\喕�X�q���	�'z�p�0�R�u�\�3��=���	�'H�l�c��(���7B6=x,8	�'��� bM5]�KN_�0o8�[�'���C�5!��v54� ���'&aL�6'�J��r�]44_H���'@�Ļ`�U"%��i��-+����'ZzlqJ_�8#	yan�<!|2���'�����j�~#8豢Z-�ІȓmFF!ё�(n�qh&C�
Yi��B�q	�ܩld�t��� !�Ԇ���5F�|�[�^������w̹���W�<$$+��1M�P5�ȓ0:����[�I��:��z$����c�`��Q}��aJ�Lڋ{o:���(d���b��|��U�s��"U����ȓk�\m;F'�D�L�
�&~��ȓH��	!K��9�W�F����ȓ��}H��׭A�fՉ�։F����
� p��̘'�ك$�����E�lCqfӲ�T��T��j��ȓ,#�y�@�N�%|�P�}|�t��xH�Xs�L�6�0��'
�H \H�ȓ-���x��ءq��h�(Y>V@���t���A��]�x��e\C|��ȓ�Ȱ�Ꝓ!�2��ˌ�z5����V���Y�"�3�IO3h�H��ȓ*���@��2�D�	#��'����ȓ'Adx�b���u����f���Ɩ��ȓg'��[%��j��D;�G%=�Ji��a� A�&]%� �2a'�!h�%��2<��A��Lx&lꧠS�v�ȓ-ϐ��#d�9:�)J����,8�ȓOv��s� <)��Cg�΂IB���U�\qeK~pn4�UhG�[|̹�ȓ%�*�3��"���J�Xe��ȓ!��4���%>�B�js��F� X�ȓ+<��8P�2TŚe��&M���ȓ0�;c��e�>��4 �!4	L|�ȓw��zs˓G��hB#�f�����6�P0dλ|�:�G�Jq:��/��ۆ��b]����I�LM朄ȓ@����!`�TPʸH��V������$P��A�#�"܄��+֍neҵ��Y���¦�T[�h�ҋԐ)�؇ȓG?�sH����ጐg�*��ȓ8U�TSm��0���Se瞋|@��S�? ���F�/Pޒ��D�Fe�ȑ�v"O���#��(_��y@P���T�!�"O�`���P�
T�:�HК|5��"OΰY��S#J������"�hم"O�aq�D��$�:��3f�~�]��"O�(����u[å[ lJ09v"Of�������d0Ս[�l��xC�"O*�i�iS�1�9�n�\!���"OLQ1�ӄv���0�@�J����u"O"ث6������b�'�ҍ��"O�s� �U���K�)<=����"O�lʔG@�CQ��҉�M'y�"O�8H��"�Q(	�ฒ�"Ol41Rj̱�̴k�[�!��s3"O
�{v��x���,�)�QE"O�����4X��<���Q8O��h[u"O��Z�� �Ca���T�=IH "O��9$lV�!�z%EӬL8��[7"O~�J�35(�&�Q2?#@m��"O��J��X�Dg��"��ܳ)L��F�'M��N�(Ͳ�!@p��w�O� 
C�I�-��X"��X�}�r����˖{�C�	0�̘���I1+���{�	��T\�C䉵T#̀�2���b�8��&����#=9��T?���W5s\�D��B9���ċ:D��b'�Y,1���DE+|�
g	:D��P(v�X�A4+�E��*�m6D�������B7�H�q/�	5�q�	�>�*Ov��I��'���'4�豯��5�rD��<W|VC�I(�L��D������
C*ZB�I�ٚ7a 21 ��3%ܶW�4�DG{J?-���U,
M*`�T	C�zм��e�-�:�OH�y�D�l:ر�Ag�F��\�w"O�i�A	�+v*1���
�3P� �U�'�1O��A�I�<.���%��J�%�"O���I����⁩(3:D��"O~����:tY����144�!"O��0gܛE~�Q��Q�w��h	��|�)�>#0�;V�3#�yFBC�a5 B�	8v��YP-�d��{����}���IW���	SŐ31����oQ!�<�#�/D�H�B�HP�½�'oEXf��ĉ.D��Z�T��x�+1��xX���c8D��I�"��
���aǢ�i�� 3�H���D{��IՈ];�x�,��!�"�*�!򄑦`/�����$I1�ՍN��OZ����#b�A�J�5s��[���/I�H�O,�S��y򫚀ڀR��/0��)��<�y"b_�.<���/}1@��Q-���'|ў�%��%�ŻlZ��XRMJ ��}�
&D�t�U�6Ԓ���ʆ�^1��+>D���h�5�Z�2c'E�~�F�ye
"�d&�S�'X ���̂S�p�P�(����R�M��A�A@ يd���d�Gyb�'�,q�ÎR�,���A���
0f[x�<�D �y�L�ā_�0�
��H���	\~�BV�<Z�L����(+0��C,���p=��]�|��'^\D�3%�4Tv�т����T`Pz�'�X�SE��8DtTK�$3n��{��)�i�$6D��OBc �Tb�"\����>�N��!���6�R�rA#�f�<i�#�c��	��A�)	�i���K<��XP8�G�;}"�!s�-7��uD~�7O#|�`�����Yd_�O�nU��E�<� �=�J�T�vL͛�+��`"O�ET���#���l�Z�,Ux""O����!ϒh���������C"O��!��i=Hd�q	��cbE�"O47ȓ6��HU�D2�nͳF(D���N60f�H���U�<hne�q�)D�|����TEh�0�/?���#LOޑ�>�CG�PU��h��N�hQYA���1�'�O?7��+^��Pa�d�1�#�	s�1O��Dz���P���bt"ôG���b���yb-�	}:B�S���)�mq�mA��(O����:ev����:t\�`��b�!�D�7,�ա"�Ü&Ju��K|����O@b� E{ ?$�ؑ���ϑ0v�x�#[�K$!�$)g���b:l��ہ$?Y!!�$J�zE�rl� `e����\�wi!��Z���W�� �A�ppՅ�˸H"2�ƓTX1�O-E����lU�A�Uđ��,Ń-I%8{X`��26,*�N�W����� )�~x��k%��0+�H#Dq�_{[Z1��4���g��$�¬Η'M��l�4�hR�J
IfN�"A�w&D�E|���\�PqCnD�ɦ�⊠�zB�	�M��QH�˵3 �	�lH�=)���d+�u������"9{��"u�!�ȓL���R'�3D�*	�w�_'�l��G���'��c1�ӵ]�H���K�:@��7*�00d��vE��R�E����u�P%�`ġ7]�Y��ϟS��B�I9H&A�
�5DP(����3Y�FB��10$AJ�$]5��Eq��N0-1�C�IxҊIs����n���˓�˱s|�B�I<jO������&�j9���.8�ڢ<1��T>��e��</�d��%&�P��D�*�O���F�����-�"��K��z݈6�6�4k?2_@�0��Z&2W���7*(D��l���@�(�b$��)#�%D��Rw풓T��eO�q�$"D�� D)��-��ax�H�>|����>����61��l�GQ"B����K[��C�Ɇ#����-N�n��}��	F�C�ɞ&�8tSĊ����I�@�H�<��C�IP����CbEe�f�
Vj�C�	=����C�Ͻ{0������
%�h�'�a}�dE�!�V��t� "��rm�<�x��'Ij���8?Ê���		؀`ߓ��'p�H�;39�t�g���=��'�"Ի��Ǿuؖ9���+�%��c�'ў�'l�@��CS��4��d#�*�'�ў"|���Zq�<�bRdʘj���e�AH�<��
#,�aZØ�>f��`��H�<�a�I� �8�k�*x�VX��FQB��0�OZl2��Ž:�h���O߯|����'��I����w�L��iRA��6_X�1�c7LO�7m~���'\X�i�J[ ��p��_оxx�'Ehp�3.D
ysl:�T>l��c�'V����a?'��Q�'$� �+K��E{����
1K�\�h�.d�@Mq�
�y"�H�U�~����"`��0I\��yR/G��]�E��X���"\��~2�'���Q R#M� z�kA}#ZhJ<9�yb�ĥ?1���Y2kh4�"/�y��%���(�OR��I����s�(��Nu&M��A[�XB�)� *�觥GCn��1�����)��'PўP�d��l��0��^a�dae�(D�t�H[�9�Ju�6o���V��E(|OFb� #q ��Gtdy8���j��A�3D�Ԣ$G�"szh�V�c��`���o�\�=Y���]?�D�d}���b�s�_Y'�B"O0�;��Y,+F��V  �����	MX�āfP>*NHA��΃x��`0�^��hO�O5�F��� &��)w�&����L�d���w>D�1 �T)PCn�RLx�����)D� ��]!cM��	S㞱T>����,��,�O�Y�T�ɑ$���RҭA�C�F9���i�@�=E�T�ձPV�8�Hƫy#n��F$B?!��,�� �F��h����ùN��9�OL1yt��z>�9Z'-�;� u�A\��F{���\
lJ5No�px�&hK�!�Dơ������%�\�a�X��!�ֵSd��H4�X>J�z-A�\!m��{R�'��	�9�����/v �Y����k4B䉱~�)@�>͂%:�@b��C�	< ��l� h�<y܀�j`�N�B�C�	Y�T�JT���)*ɚ�iQ [8B�
�r��#��h�F@K��O~� B�IQ�`*�ǂ�6��3֌�4F��C�	�X <��)<c�l�E��s�C䉈��� e!Dn��z0��C�CۊMk��W�oIVp��-�"J~C�]��R&��*��X��DY&O�dC��#��䛰m�3\��U��'6�B䉮S�>�r�?9�X��a��
$�B�2��ac��:�u�gO>|J�B�I�B�V@���!P޼����2o��B�	�)�����)�5i���둤xT"B�1{ۖ9#�8]��b`���9��C�	� ��(2č��;�a���C�Qg&J�#Ԛ|��E�i��Y&�C�	���Q�&\�1@�AN}�tB��/3 �D� �^��Ma���1�*B䉗p� �{1���0܆)�PXc�C�I�9���r���<7��M�G�+�C�	[����	�+t]�E�=6�C�	�w��d�/����_"f�C�I V�Z呒��7H��ݢBXC�	� �>��Vq�z0��!�:(C䉜f����bhѱZw�m	`LB�	�9r��fDyWti��I;}YfC�I�D��	��+�j59��IO_VC��Y�J]I��:�HG�"qG�B䉍	�mc��ڸ<��t�
_*5�.B�	6e�B��F�1(�����-x3�B����*P��d�
���}f�C�lt�e����
,d��s�D!fx�C��7E�p��tl�8#k��+c�z3�C�	+`@|�z�m��/FؑRN�e>rC�ɿm�$��E��\������
n��$H;'��0�U�E"a>z��%��0c!���Oބj�a��4�� zj޴s!򤟰Pfd�8Q��.9~V����D�!�B�gȰ�1���?Whp�ؕ��!��A��|�s5ːE^�-2���G!�d�@���B�O�t�7��9�!���b��0e:
�xA�.�!��Үb�<��5�\]�&�!���-L��5ρ0C�L%����(~!�� F%L��8(pT�5G�+��m��"O���7��s�����M�R9�"O����[�r��4��-؊F|�Y�"O�I�C˹1�0!�,G�#�`��"OДv	M�����1O*�Y��"O�\򠭟6!�b��ք�4�%"Onl����=&m��Y�B^nʬ�a"O�%��O�o&V@Xk�D逩�#"O��k�gʩ0`��z�_�ZƜ�I�"O~��QM	.2�X�
ĝL�`h�s"Ox� �[m���W�=Q��QZ�"Oح�͒&z:�!W�J�HHX� "O�l�Ak�~�Ȉkϊ8.���y�"O�����1`02�R���o���Q"OΕ0�O
U�&�A�NT/0���"OT�)��/%�H�a�O�
�:`�!"O��ʅnU/M��sp$Yp��
�"O"E�&��f����
$<�~��R"O�A�v��v�(镢�!��$R"O�99t��,?' �����%H0v�"O:5[� D.=D0HPÐ16�� �$"OX8�S!Q�_M9�F"�D�x0�"O�Š&�^�(�^����>��`�"O���R��0�tD� چ9���*2"Op�{LR�QV8���ŉ�^v��J�"O ��F��<�uaƊ�_w��*�"Od$��`ȅ:e�]��Ծ-WL�qG"OJ!K�l��X|����Z�0�"O4�*����Hl�1�!�7��\�"O��UK�,|H��`S)[y����"O�dKu�X9�ʥ0�iɽ\m�!�u"Oؕ�BV���ə���X&h��"O���c&�H��q�B8sj�P#"OX0)P,�g�e/eUz��צ	��y�
sLz���[�g��{rl�6�y�C[$vQ��"7, `��H�Tk�&�y����I��f�	S��ݒ����yb���	���嫔�Lt*��"�y"&P� ��*[P|B٘�)ٻ�y"��-�6z�a�,ST�$a��yR��|蘴�tOK7V��`�ҬT��y���b�^I95�\ _�\�B�P�y����)(d�K5��%���y"�G�L�lUj��:��l�CV��y�/E"�`�[���5$���@uL�!�x�"�vLX�D�k`�y0Q	��V�Qr�*G�4N ��'p����ĤORD���J�CmtUъ�$�6%"q�JT�z���?uY�BӪ%��@h�ȜN����B(D����-�<�&��D*�jŦ����?�x0r��W")5�����3��°��I�0�òC�ZVZB��,@�&��o�*gl]2��X/�t�"T���r�b�%1���R�'R�ҧ��>��Q�o��1Ś��Ŝ���>�5�\�y M��; 
����L*{h��t*0�\��c �X[Ĩ���&lO��r0G��M��ȴ�I�^���:�鉡]Jf)���Z�N�Fx��ݮFYXҥDփ9q�)�7E�P#\̚�N�TA�|��'ph�#��2m�����Iz�]�G�>��p �暾B�`����kvx�ʍ��Ͽ'�P�*Kl�s6%�����RD�<�v�N�"�p{'FҕFD�����n���ROɶwe*A���X5<<��yO��3s)*�I)�pij�O�0:�)jVH˸k����dѳCY�I�6΄�|����R'�@��L��F&Gh���m�.)|0�H��O�ubhb�� <O@ؘ��� 8�ѢƆIX�5���ɸG8���Q3Ey���͌�!��S�CY	��C'AQ�	��#�h��<�%J�ph<�2���*e;�cB+
i(=A��>(q�a�O��g72�� ��A`���Bg��,m3N~�;5C�l4Cߴ��Q�7��2xs����S�? �U�U��g���!V�C$(	<���͝^�<�h6�ޝc�,l�"@B,-���Be���֊"�d!H� y���n#,8��M�.{a|B�.n�x�#�ѦW�H�x��φ-�|Ԓ��3X�@D0�)	A&�@�bȆ,Z�!�5�'��uY"̚���8�U)QV䳊�� �~ST5�2d�lx�`S����Eճ,H��
F�DH�I�aE�@�T�r�$:4�� ��)�RQ�&o��C�>9�Ӯ�T�r-T'm��Jd.� Z�$��p�!+�TY&?�]sa��	�AZ���I�!���>bpB�I#9�~%IEn�DA�VD���: ���Q�Ba�qDѶhN� nb>-QΔ7Ce'�!!$��7Z4�)�	9c~�H�D%�OL�9���;&"��HR��+7�)r�Հ\Zp������3���%�N-���
x����$��Vz��(գ�#��鐯B�u��\�N?������FKB5Jsa�$�P�S�*"'` i�	Ҫ]^0��ǉF��(�ƓT� ���̈�
=�x�%@�=R�A�l��hςd�@�
�\�考�Z�P���֬'��缓3�\�*m #�X�J.ޙ8���L�<�.љ;���k���4yX2�14� ��3_�F�vDi�k� �*0�';���C����)\H��A鎓D��ň.��o�Ȇ�	,q�zl���*�PY��E�
'�e�!�Y�&䨁��'T�����bx�u+Nx�`�D*� d���P�B�>�N���#>�|=�q���g���rB�:�@����7L��X�`��5gHP��;U��ѳU�?D���� �h�P`em��p^Ru:�FO,?��殅7RѨ51�ŕ&m��ң�i�R�>�n,7�dѧ�$�H$�G�3{!��[�(�:��KW�.�ra螭Ȳ=�r<�tQ	 LB(��ł�\?���
@�++�l�.t�J�
c���F�p��ɜ D�`��B��5�4�󊟚��\����4��i�aΒ9��9�(K%+ a{r��H�p�`��$|p|�ؗ��;��Ol�bc�l恻ԯ�.��|b��柖��x��\��,�y��6"O�i���2[~�H�,p��K��~����e�R<	p�2ե�3��"~�§K�&�q�ě�6X``RG�H�<I��[�P�(IR�I��,�H�p��F!E�����O��Rʔ�Fn&>c��ӥQ0<	�@`ᅍ�~ $.��۵N�>g4�Z�%G75(�(�7lQ
+Q��cf��_pp��I�3���C2��,f��� GO�KbC�	�b{z��'�&�� A-A6^B��-1BX�PF���\�SF��8C�"�.+C���nF4����"{��C䉗D9$]�`S�H� t��;��C�	�pU�p�o�pg~I��Y &��C�	# �ޜ���yd����X�`B�I��ܨwǏ#z���c,߉+XB�	�a���T!Q�	9�)b$��A0B�I-D�R`�S#G�Y8F�*�(
hB�I�9�<���Ci�B���5J�B�	(f�@�R��Jv����A�?��B���F!��LI4��5��3h�DB�	��ڼH�F�K�E��N�pEB�ɘHr4���`K�F��p�`��Q�C�I;e}nت��I����O�	#�C�I-��yaD�޹=m�AxG��~�VB�>C�F`GmT0�P3-T���B�	8/.�Y�i�bQ����(X#S�fB�ɹh�����\'`�� HvC�	H]$Da�.Ĉ � ��@��B�C䉷2�5�v#�	�,uK�J%%��B�	�ed �+g �A'�ђ�"O��@���Kܺ��� $����"O~����-��]����3#�N�r�"O�5����~��0��fa�25lō�y���<ԩXA��!!H�$�ԧ&�yr <(�4}q�����px�D��y�� ��0ٛ�-��&aá�<�y�`����U,�'�IhSFމ�yBa�>K
�뒣[Jx��CG���yr��Y���/B;OؒT2#D�y����3��Se��Odn�BC����y
� 2r�۬T9�t�B�,aX6)Q "O�;GbI�R&�Hǁ[�"&��1�"O2����=L���fK<c�<C�"OP�b`G!c��t�f�Ѣ4q"�Ra"Ov�ِ@Y�>��pXW�
#e�,�C"OD���B�G� q�f)�"zA����"OV��Qv��!��G�D9pT
�"O������+3�Tk@&ֈB!tM�u"O�LQ.V�.�q3��M�2��T˷"O-��^.�R`S��(~��1�"O��0)P&uה�83�F�v���"O�E�4ʏ��1jbi�=�� AD"O��B`o�
Eo���gQv����A"O���q(B����I�&��s~Kb"O�D��+�0�(��Ѯu��1�r"O�ո7!�4c˲�`c*M#A�:�k�"O�ԃP#��H�I�`W�ѐA("O8Q%+�7����B�F�A�:�"�"OV��мc䢨S�m��+,�E�"O�@�B�(*&��s�-S�xixDJ�"O�7*�r���#nR0WE"!Y�"O��җ�������L�c��%"On�HuY�_�0��t�؍D����0"O��cp����i��5z.��"OF%�s/��y��Y�@e�8Yv"O���2�c!��!�0m�`��^�!�]-LA�C��5a�AJ�D��&5!���l~}ʶ�zW�쑡��>!��pJ`pFKȩ?5�xJ�(S�D!�N�%)V�uc�w70E�5�^3:!��L7`� ��e�8G9���g�3@!���'�FժULL�L CsƊ6b�!�12q��y͇�o>DZA�ǧOs!��(%#�mc�l�����Py!����~�T�"�oQ�{24Hd(	�I�!�7����lQp�����g7Q�!��"d�4��q� 麗&Ŋ:�!��"$�~y�/�1s��iA�Y#u�!�� \Q.dAS�2	��z5�*vp!�D��e!��A� �0U�(�2�l��n�!�DݔKJ��I�DF
&�ꜚ�kK/u�!�$1��e!����_Fl��� L�u�!�ߜQ����oLX&���M݀�!����;x8r&�_ ��%�@�+�!��ܖb�~���_
-{,�i��A)W�!�6j�~�[�
��Vi�i��0R�!��D�phJ�!��iQ��i���!���4��$4����u[�hS8b�!��]l��$	�C���Fq!LU�0�!�צ��U�[@�l�yԅU\ɊB�:mO%u#-$H���j�C�I�w��tf�W�.I���iXxC�I�(3��K ��v��ca�=�B�#���G	�!aH��(ʡGt*B�I�a
��J�ː>Q�R��֊��f��C�%K��}j#,b
�J�L^X�C�I-f�쁡mչ���;5L�#S�C�%:n���`��q�P���.�2�C��?wD0U1$�$=�t�I�Ǉ���C�ɒ`�N��G.K�Dd��X?AĺC��'z�<�(p�ɭc|3#
Y+Nl�C��.�	3&O[�~��%�iUx�
B�I�5�Й�3AK�r�J���4w�<C�	��:�:2(�a��(��.y-C�)� p�*��F%!�A���۱[���:"Oڠ�UG:`J=)�A^m/�02�"O*
E� ?����6yr�xb "O,Q��#�(�t��|fFq�"O��:�O9g�܀���Kw  ""O̤:�H��)��ݒ��@1 ���"Or5P'�+2H��â��I��
2"O�	���R`r�f ��Hy�
�"O�4!���_���*sN��ZW&��"Ox=Y�h
3{d����T]���"O�u����lG���R��m�@\�"O���իH�V)T�@��8>f�@�"O*a�#X�4�ʐ�	��|@��"O^���#�5�x��R�'��*�"O0�Z�X�64D;�ǖ�<��$
S"O�ē��9�H�����\����"O�Ջ�Ƣ�`���͂M�\�u"O�@�Eb�,�@�`vk�(L�Z%j "O�LbR�:Ո|C�)��v�a"O�����3��9�2�S(~.���"O�,��!H�I��13��Lr�!�"O�Q3�҄`W����K53h�)�"O�][�CL�����ܼ1���""O�����bgN�K!��4�d��"Od�K���:f�bYxC垚<��P�"O��`��A<>�j����ǩM��%J""O(���B�keʱ��1E�x:`"O*�����Z}t�'��6�$	T"O0q���^����G�5&W����"O�a0��Cu0.U���	�L_���"O`�8T Ԣ`��Ƅ����'"O��X�	�;���[4W��:�"O�����E�w;�쁢��F���"O���ڒ; �$�ތ.��l�"O�Y����:eXb�κN���q"O��Y*�8�ly:FF�)ݜ !�"O|�F-��J92Pez��N���y�Y<VV�@�&��A����y"==���ˣe�'ڦ�H�F�7�y��94G��K�QD�5BG���y�� ��g!�6G�>�����yBG��$�u���O��F�
5�y��#��h���G���t@
$�y�-�&nl܈`ȃ>F���To���yBg+p��e�R$^'���:2����'.�@����N��U�U3}l(P�'�T���ǁ1N*�����pU>��
�'��K�역%2զ�~N>��	�'�,L��J�R�),.q<���'�P!VH�!\��$O�\�*9�'-�*�ȃ*�I�%D����'����Y耊'�X)aX�Y��h�y"�[5Bt��IS�1^��x�@�yB��C��PvI�I4��Q����y�Z�'�-�B��^���3����y2�"S: � R<IzP(:�y2�Y�O�VHP�F��I��`:�AB�y�ʈ�+p����E�2�`]��yB��t7��q�N��b�.H��o¥�y�*�?\���� �J�VY�COC��y"�����A;���K�$#�ޅ�y��ѺC_�Y�P�_�1P��gD;�y�-�&-�R�k�kɌ��x��P$�y2c� L�3e'}8�@ voE�y
� �q��!4""e�%M�4�.��"OM9V�֥T���S
��p)P"O���)�1�*�8�B�s�"O$+�;�,�5�B9^m
���"O�;V��#$z��GZq^��"O��U�Ӏs	H�2E��L��h"O�<� ��)Al�P$ؼ6���1"OBMz�,�A.X�3'���h*�U"Oy�0�J�I�]�w�"��ͳT"OX*�O�1s|�a�1���RӚy�d"OP`�pE��L�08���T�R�uI""O�$�i���3�LD�qr�"O��S��I7'PP��=�l�Sw"OJ�B��~O
)��b�=����e"OZPهF%L���f�]&��@@�"OD`��+ѢS{ �X�σWA�\�"O���v*�]��g�*,T"O�x�.72 ��/U�ʌab"O���'�7�4E��S;P$YJ�"O� Z��9�8P�����$W���"O*x���w�Y��N��	��H'"O
����_��ٻ�O_�q��Q�"O��BTCS7O!c �?n�z���"O�H;�K��`�b��$�^�w��T�"O���W�^$I���	�S�j�1q"O"u@�ݥ+vҬ�R��S��Q
�"O4ݢ�`�����E��2  d"O����)A�r��ę�ۣ"�^��"O���XU��L"�,���6�Qt�<1�J��>U��3��_��B��i�<1��A
�������5�Gbd�<1Q�M�I��1�g\z�
'LXb�<�[$,[�y�Ƒq��Y�ve5T�8�P&B`L�sV�Ӗx��+e:D��a5-uN�2��_�;���1,&D�l��M,(1Sd����Y��$D�d��I�*����l�"Ppp �b,.D��RcUCa� ��mZ"}�HH��G*D����B�8�`�r���e�L*F�*D�4[��A�)�mP�tV<�K`
&D����(=�� �p��'K���	��'D���&֨KB.�#�	ͣ*�r����>D�̰��M�ESn�U�M�X�6�s`�(D�4+���]+�]�I�',�8#�%D���7�ދ��ɰR��B]��� D�dPA�R$�������	2���n5D��aKϞ9i	 7���"��P9��3D���->t���P�fľA
h\�RL,D����,,��٪�̼Sc���e-(D��+%D�9�����`�8`�� D&D��h!��D���sSbKN�ڑ �$D�\i�`��Y}"��c�6ܹ*%�%D�d
�i�3ei�	BB�h���0Gg<D��s��0oy���(]%s1��Y�&:D�DP��_J��Yxs
M'C�D�f@6D�L�sn�NS�a�Mޞ8,2D���.�=S�^� ���\���g*O �/K��H���-��RQ"O�Hj��N�{�"-b�\#nfq��"O�� ��Y>y"�@�`\�U"O�My���m:��#,Oz���"OJ�R&�;'�����*�xAB�"OVh
a-� � �;�C�P��l0�"Oi"�,Э>ߺT��X8|NH�A"O� vd�D"S�U��K��-�d�D"O`x��oּ]1 �ꄏ2�0@�b"O~ŉ��T3�J����ٜM��R�"Oh" ��:kB�	{�H��|{NH*�"O�D� E��j�r��qR���"O�,�1,�|6TYl\�f���p��&D��y��Y�VaXt,��9.��"&D�d8�O�MJH ���*��U`Dg&D�,;�i��hLT�1t	T$e��K6D�,��/�zð�j�$0��rb D�4��b�(;.���䏵,���o>D�����8&�����M4
0rgK<D��Rf꜖��bW
(���o�7�!�Cqu�͓�ԊC�.�iǅ��a!�d��!�&����!��U<!��>P��"�'�c�,I`�A��M<!�dh�d�PkU$�q�,��{׺�R	�'�2�8q�/;��#Q�ʳG�4�k
�'�Z�ɱ�G4L~.q(A�DE\��'&QA�;1$ļ����;5�tQ�'cҥC�	�CƁs�,̟)_��	�'���@����4Y��k��32.�A	�';^�[�a.(�D�á	
�{<� z	�'\��BC�B�7tJ�3$���b�$��'���G�9j0r$�@ƞ�XA@��'�(,ȧ"��@����?X���	�'~\0'��Hn���,N8H\��'k\Ő�*P6J��E��:���'zN(�5�=LX|j���*݈�'I�h�ҏC=D>�S� �_z�,	�'FI�k��<��L�W�T��M��'3�|�1m�9(�Jl[�e�N3DU��' r���G�)p��#�R:˴+�'̴I�S��9
 �|9B��G~���'�	���7	���A�I*:��Yi�' ���q�����[2�\�!�'��\H���&R��qx��S Q���
�'j2Ef6e��1w��J�Ě	�'��D��-͈�:tiF
Z=�REa
�'O�t� ꏲLd��̝7g�!Y	�'��e:��Fy���R����_*�I#�'�������
J�Z���㚌SM<�;�'����#uq�W��S���'����V�>|Ґ5I�d�[�$�K�'�����j�\$�=)F�^T�I��'�6`�S�y����W>��X�'�f��F¬tW���/N�X�11�'Z���
�QZR�a�N�5H�pc
�'�8 e��;H(���DL�?��DH�'6<9k ����l�F7���'�<�"Bc��?;нqDC�6j�)i�'��12�$�� �ެ8aE�f���	�'7�1�6��.&�o�6�@�x"OH�����vG2mQ�.�2N����"O�e��e�>�E��|���&"Oz؁��p4�1��y���3"Of�PP�P;,���ڀn� .tr�a"O0���g�k(��!���q� ��"O�`2�ဓ~�$��D�EMz9��"O8�S3���4� �7&["84"O�<���A4�\��K�#%�y4"OD 	�dI�zuH���Jۈ	�@esP"O��!���mYPGɕ�"��"O���A�p������ v���"O� ��R��zyLm2��E�*�ũO�)�I���?��tl3��M��p��Ǘ�@�)6���6���T�[�gy~x�'���*çc�rl���x����O��@��|3�����G�) ���O,���Ӧ��[<F������DX֢l?�!�Ϙv��tH��r>U��,A+	$\A���Jy�@:eix����`��T(���GO$S����IÝ��b�\1G7\A��%�2$�6��A`I!-g�{d�U�\^��O��e�&W�`���#��M�]�"��AoocrV��?q	_O>��Q�֊*_z�2K؈gD�p�(EDh�Ί�)J>mX�NH -PTMඊ��lvJP�AƘU��DB7Ula�C���2��s�q�������I�V��Pk"D�5a;񄖦F� %J�6���5��o��`���ɩ4~���_� ä�M�@IL��S�>E�$�ИB��ɡ��1-R%��G�;�?q1����J>E���K��(Y9�X<�!��$C�r� �p?�s'�:u���
�̔�����W��Q�<Aâ�>PNN�2�I�o{���EJ�<ɢ�U�f�(�S�K
W����c�k�<y`��'O|��d�
^�l����f�<����|�ehP��`[ڝz�cm�<	7@.�6%�6�|�&�XR�N�<����%e�pP��5Y�yX�F�< ����E�1/-M���B�<-]��e(�C�1f�!�&��q��C�"pԛ ߠ6_~��uႠd��_ �.�	ң��Kp���J�!�	7|=\��E�FF�m�� !�$F!|����&fP��쐬<,!��ùS��Z$d�[T|���s!��9�Ll)RjJ"ibF,� K�7XG!�� F����_�A^��q��8=!�ą"����R�{E��e��G~!��W
(�P|�+1D�dj�M�|{!�dNEZ���<:>M�kP�!�0g�*�;�GV�5�HI%Eի\!��\F�6l;�n��^�����b�?w�!�$1�R�5I2Mx/ۣ(�!�C�<X����AW:�9�k�!���@�T<�3,\����D
^,!� ,/H�b����eQ�!'[$!�Č�n� �����J8��:�!�_�8�N=`&��j��٠��JA!�D4L�� �ʪ9��D0T���!9!�d�74Բ���͕�E�.A�rL�'{"!�dH6� ���]�m�$��Ë�#-!�D�/����ʓ*����i�}C!�d����VCI���	G��2/V!���L�bA*�*Q,_��mC@'�{K!�$>s����T��E�$-E!�S�6��T�GGK�|���U
Q$a�!�D�}ylA �k��^_Ĝ#�HG�]�!�$�
���@�{]R@��(C��!��˾�@E��ՙe: �r�$I=|�!�$5�9�F+��C;��`CQ/io!�$��4�b��E�d�YV��-�!�d�y��B&�Bn��N.b�!�D_p)�xeP�u��eR5���q!�d��Ag�����;A��!���й0Z!��0*-���vŜ�J�D��ԣQ $!!�$;'�n�"4��r��R Õ.!�dğk4���G�W����ܔ�!�dQ�d�,���=g#<MX�%"X�!��KU��E F�	4�J���i�!��e�8��� �P�	c#S�!�D
�iphɗ�)�������!��%������#s�	3� ��a�!�� ��je&��(�,9�ƅ�e��<"OD}��f�ML>#�&��P"OX *e�Y3:�m:�N��g��9C"O �0�\�,�h��">�D�@""O�l�FÇ
����-�C��]��"O<�S�!��m��B�E�����"O2u+�J�9$�h�R"I	z��!js"O8�C0���/�}�(P�d����"O�I&�W	l�q`��I)a�8��2"O�E� Y4	>]�DD�1wAB�"O��ӓ-Ҩ`φ���E�t��hR"O|ф��7�l���L�-�6�e"O�q`��Y/��@Gl��ưHp"O�3��hE5K/�0g�p�V�\l�<Q�ؖ>z��xC�-l=(�2��C�<���p�D�1c�L�Wy�{a�@�<�1.�2��$X�%	�uv.���Q�<��=bq8C��(��ppL�<I�,��7If�
b��%w��$D�]�<ّ�m����Ƨ;"X�!���^�<�T,	�?�H͊E�[/�����X�<��-_�7�
$���6	BpA0a#�|�<a@C�v?vժ���VT��b�M{�<	"J�"9:���,U��A�w�<Y�a�33
��j��h0��oq�<! M8�:�*��
�Zh�Ah�<9�@��@Ҧ.��a�&�+�� d�<�� �S��ML=>��`�C�y�<є!J-2�4D3��=F����@c�x�<���I^rp�sH�q嬩�-Aw�<I�H�u��k��k���	Bmx�<!6��3T�eKeƏ<�5
���X�<Q#�7m������Z��l�$��S�<�lW�{N�8��ݫQ*q�@�U�<�U'ʭV�$Y!FU Q�n��3œO�<!R$0A�$��ת;sj ��XO�<AGC�yLp9��B�t��)�#&Eb�<)�hTz�Zm��.�& 	t� U�<�+fH�R�"Z!�%Ґ|��hO�O��c��#W���#A��l�q�'����ƈ����$���вs�\)�'L(2,��e ����Sp�"� �'�NE�bײ\�J�JL�/NP��`���pW�:��hjE��6sC�}���d�ԟy����숩hu��S�
:@F!�d	�#�QvhۯcϜ�fL�<#!�d�)z� �a��S��p�$+U�0!�)��pB�Ґ��`WIÄ*7!�D�9"��̪'G$s�����w!�^�Y�~D�Gk��YH,:��\��!�����j�N��q�GL!�Y7?��;�!ߴT 䍰�I�3h,!��̑1F�%{p�?G.!]�8l�'���@� ɍeLDU)���0�
���'�$d+2ř18�`A�qlű07�4q
�'��@`	A�c69���!�n���'���K �jh:q� �,	��(��'h��mV�drp�CE�0|HR�`�'!2L���_�Rh��0#,ш%�B�#	�'A��	��=1P�QrD�"��}c�'��9�� F�B��H1�� ��P
�'<�h�aڪ���ԅ�3H"��
�'�������lІh�-7�(�+
�'Z�4���̬o�8d+��Ț8pаS	��� �����5ل�Ӳ�ɮ�0t"O�p�
a�D�Pu��*adbD��"Ov=��*��{�
5���vTj\�R"O	���A���R��ipA"O�}�n�*S���
4���"O>!�ad6�4*2� ��� "Ox�.e�fz�C�:#�b�c2��
�yB���n(��2A��%��U��+���yrE�+V�n���φ�\љ�/��yRꜹG��i�r._�5�X�k'�=�yb-��`6�lX�R.��y26�!�ybb�1"�|�#6&A�^���%I	��y���:U�(���c��J��Lu�0�y� ��#1E�0,�j���k�0�y2EJbZ�m�P���"� �dJ�y�gH��l�r��nm��k�8�y2N�C}0��q�Lk'j)��ڻ�y���R� �d�:�� I�M��yBi�b�
�(�hX=(�4���ĝ��y���6^2��S�*,40p,��y��D�j(��X�阣� ��PC]��y"gw��(�E��tT0�����yiûU *��G䁝4��I�&��y*L&b�h���S3(�:��J�yR`�H\�ՉI	8���Pb��,�y�-ȕ=��m+�"?ю`��ݹ�y��P�<���@v�A�/�=av"�,�y�'_���9z���*1�� U�\��yR S.R�dLӴ�U�ҥ�ϐ��y����j��[�6N��	ch^��y� S|,]z��:(�Xm�⁎��y�,�L���1�8���%���yR!ӥOe��iE��S B!`�>�y�\�E�*�@7���_Z��i��yr�Q�iGb�ct�E�RQT�����y�Í7eȅ����7`����W;�y���q���Q�$j�y��Ƭ�y�р2�^q1&i��#�"9���yr�V�i�(A �h@��"�9$�֘�y�|�܈����y_N��db�2�y"��6V�j��k��!SQ#��y-�%+ڔ�BoH,14�ub'Ȗ�y�E4)��Zg���?BcS����yd�*�P�lήm���9�ѓ�yRG s���3�N8���r#h�(�y�e��x�p�M�5�-P�ŧ�y��� �*�B�(^&�@Ȫ��^��y"�A2@�  �P�>� ���/�y�m�%�Jxⷮ� �b�RF@��yb�ް_X���̶�I�&�&�y�J
6-���x'�¢'�����V��y��ݫg���)�
�J/I&#���y¯R*���cW��H�j���*�yR�S��<M���O�uv��C ʉ��y"��5Bި�J끂h�`�j�� �y"�ĞC�,�C�	%Y�x4�t��y�e�68��QJ��b�v��#�߅�y2M�;��j�E��T4T��j�4�y2OX�C_mb�H S�^�+�U�y������8R���D���rs��yB%�+�A`�O5��9�g��yR��H+F��0oM�:ά0#��yR<����b�?fg�	F-��y2#J�7,���`0�`����y
� `D��L�%;l�2�K#<R���"O�,K�̶	��Ca�i����"O9�� Pv7=�2� �C�Υ��"O��B���J� � 1�%җ"O���W0c�8)�N�;pyT�"O�"G�?NqB!��;zv`д"O���������rl�yS"OT�I��<4��R,�W�a�6"O*eSQ��=a�$�A�O�wLFyZ�"O�pRʃaخɐ��1٫A"O�=Yf�̏/� �S&�Ԝ/D0y�t"O^��U�ȣP���E�>�@
�"O�a�#��l)Uɐ��!"OftY�∈\4�D`�[;\��X�"O����)�\�T��7�S��� 6"OD�
׿qS4XťJ�=��)0"OV,ȖJ&��\�V���:.a95"OxI��H�~�zu��A>*QB�"OfD��(�%90u���A+�b���"O��A7�\w��s�͆Km~`��"O�L���ܜ�����6SJ�˒"O|�۷�ƭ6�p �C��G�z@A2"OT���`�)EԂ�p�Yr�($sC"O����r��v�͐=�V�C"Od4[�*�52 P�ₗ�0FH "OH1s �Չ4'N�Т��L��)2"ON�uJC�+�|�Y�ؖ�(`�"O�p����"	���d ���&�E"O�!���U�*R&,���
�@w"O�qS   ��   O  	  �  �   �+  l6  oA  J  uU  h_  �e   l  Xr  �x  �~  !�  c�  ��  �  '�  j�  ��  �  0�  r�  ��  q�  :�  ��  ��  ��  ��  ��  �  )�  � �  �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p G}")7�7�``5�:Q,L��R�H�2��#.O ������܅kW�� ���bk[�%��Q8�(O?����4�|�z�+*�Zɨ��;���d8�SbSf��boۀ��%��R�%��<A	˓ �R��V��2)��KE�`�@�Fx2����}ʙ'�i�|r��2E�0:��L0eO|��A�cR��IV�$<t����+���<�Om���!#j�$�N�A��;M����!�ybF�:l�����F1,*�:�+<����D<�~B��$Y?}�3	��7'�<HB�K�K�v� &	.lOL�x�b�\�C�P� ��f"�!�V�7�y>Y�O4����-F�@���� 	���nW/Ĳ��i� �>a����IƄ���C��r!v�����J��p��I�u���c������Q�^�I�[�xR�|��tp��U��d@h"��?Q�'x�ə� �(C؁���lᓏy���wܓ��'K�qF��F�n��0��	��l���k��F��/��!Bz���V;7v�D�w��y�aפDB�PJ�D��`چg�1�y
� ٱ�d��X'��P�^�@��R�5O�b�`@��<qs��Se�|	��|�2¦��P}�)�'6&)�Յ�7`���貂��DoD(<I�K!	}��*� �m�㪑F��L�>Igc�{9�KnM�9~P�kP�@�'��?��ӡ��J�"�>V4��ˑ�?ғ�hO�Ӭ_����UJ�Hi�)e�;]��	u��h����dg�'�r����fG��"g"O��2oR�T���F�:R�� ��C�d�cbR�M	�����"f�A"�>�Odӧ� �n
���c�jRP�'"O2��
�H���0P'�m���IA�Oy:i��*]���xp&<Df�Ui�'=����&�(-�&�ڧAg�}�'�@�z3Ɏ�`�����B�3~4��
�'7�l�w�_l�lȒ�ͬ&��y�'�ў"~$�P>/�̉�� P������O�<A��mO o12�*���L�lt��D��,D{�'kDL�&��J���4��Mh�U���gyB�˙q&P�h���*�|�� ʛJ�"<iϓ+�~�*�ȕi�x �� ]5ڰDy�X>�pѦ2+ˤ�!#JJ�Y��]�#;D�4����>弈�,
�=� `Q�&}"�|������|b���@�$`�!�A�$R�)B)�yR���v��呠O�l�J�iFdM*���0>�`aɰ2Z�
C�^#Z SQ��I�<a�h�x�6��#��T���CD�C�<i�� ]PΡ��F�*p��P��c�<��撚�ܽ�aA�U>\ ���X�<Y�1&U���F׿HZ�|���HY�<QE�	o)5{w.�&b�qQ��V�<�v�F]|I4�ˉ%#rM*6S�<1e`��~�H�8�F�O�&�ВΆg�<y��F%����b(:18v�n�<�����8 d�Уk?&�Q�	c�<�B�Pm[��a�bל�.��.^a�<Q'���2HY �YϾ��BfE�Iy���O�q��EZ�w��M�{�\h��'Ј� �Ċ�g��Sa� �y��љ�{r�'��x��d�@�P��2o�DЁ��~��:N�LL���ˌ\l0ECfJ�!nB�I"�i�0���P���Y�j�*MW�C�	O`"�І!�?N���b�Q�u�C�I���S���r�\$�1Fx� �OZ�=�}:��#t�MKC�	
���@`��a�<�f�M�Y����G)l��U�Z�$����I�m��a�g����0�#F�MۂB�	=J�x��� �]h� �&+%'�(C�	|��������(�p�	}�6C�ɥZ	ta���.9�N� @��fB�C�	0O�,��#�47?j\4A,{�C�	�a�213����=J�o�o�C�	�q��ۦ@�Kh"a{# �C�	>5������5\�0�"��Z>XB�	!��-��'�([��ɸA!G�*B�	�w��\iS��c'(A������C䉨���Cr���%��(�&syHC�	$�Z�A`Ua��`�'��S�Lb�@�����9ҡ�?^�����Cq��	�'D�X�3jT�~,
��G�t�<<q�d� ��5�I00��EO��!PF�߳-�B�ɀb<�Y�/D�'�-Z%��6>B(C�:�ܣ�&I�2UaWE_|\��	u����(����C伉 * I�\�u�|Ƨ� �D[3ߺ
���1��%f��<`4�$;LO����P�$M�B�	A��Y�S�'��ɠ:���9E�I#!+�Qj��w]NC�I�6S$�z���0:wB�遂��k#�<�?���$A�Dj\�z�n�Z���c�T�yR���� �*OO���t�ߠ��'uў�Ohdİ�,�+d�d�;$㍘D�����)��<1�G�T�x ��DПGx�a¤��]�'{�y�Z4:]�·PiB�uxdi�'��HP#I	�^L��1��?rnQѲ젟x�P��wX���/EJJ�B�K"V����$lO�j6b���*�Yg�oy %�aC�!�hO?�Ү"^x�V�2@��l��g�[#铕y���	Ɖnm|��QHF/'�5�F�#��Y��4�u�0M/�0�G����c<D�x�ӉV��q�掇 �>���&D�4��%����55mF;�8Y�*�>)�;��철-D�{����:f(8��4&)be'lF�9"sʃ�rhh��ȓ-��]��
 &�,�aK
Q�M�'�ў"|ڶ%ɭn��I(ā<<������t�<	�ʒ �.	(ơb0��KTg�n�e8�ZT+0)NP�h���r
����6�O��I�1�bU����洛�jl0ȆȓI\Ҵ!Be����d͙�'���G}��ӭu�R0p�"Sߘ�ؗ�Q���C�I�)��a��[;�8$y'O8*��'�ў�?j��	)�
����E��� �6D��As���$D	�R�2�Z�F3D�	�����ӱj�+�!��/D��qG� �쁈C�N	���AU�/D� 2��GD�>h�&��y0�lKQ-D�([�j�W醼�`Å�C
���)D���G��lߎ�35b3cǶ�5)D��I���q��ҴkS>�P��%&D��
�h�h�H��
ѹU�0e:�!D���M�{%�@*5�MF�n03�E*D��!���~�n�ps�M?DM6,Y�(D� �I��O���F��\
J �uF&D�h�,
8DA�*�8X�s�#D�l	Cے��)��0�dp6D��#�P�Y#jUkf�J�걒��3D�x��T�
| �8��ݷK`z1b��/D����爛,�Ri���3Tb͓��.D�<��"��[~N	˰��!2�%8s�&D�h�Q��|ƚ��Ei�Ј	�@2D��(g@{HEd�\<&;|7/�Y�<A���.W[�=j�H\�e�||z���W�<Q���j��\@AE��{�EZ2RW�<ٱ&چ*���r�ͼ2���Q@c^G�<Q�l�X��S�COq�	)�Əz�<�B
�b�Vl
�G��i�PH���w�<�.%nTƥ�E�F�z��pQ��^�<��*}���v�V�=�`P@k�Y�<9�7EJͩ��M>]VA����T�<1���%L��hБ�9+��y�E_h�<W��"!������Z��`ܫ�Nc�<1�]	pThA�#Άz��\&�]�<�vᐷ\bx�����z�l����P�<�i=O�m�E!	?b����P�<ɀ�) �0[�
J�s�� !�M�<�TCQ�F1�R���(%���C��E�<��ȏ����*�N"7���+�M@�<Q�Nܧs��Q�q�ϙd�H��0Tz�<� E��GuҶ%zDG��s;��c�"O��T��gU���oZ%i�Z�I�"O�Qq c�9\Ђ)h�eD�1�^|ڤ"OJ�r� .Zzb Cʄ�SszՑ`"O>A�W�3 .@�#���H7� �s�'b�'�B�'dR�'r�'2�'d��,�Xޤ���H#lo�����'���'���'��'o��'g�w�.e)ԉ�>'���0�B��l ���'��'��'�'r�'�R�'�>�A9���aąS6r��-���'iR�'7"�'�r�'�b�'�b�'P��:�(�9
R40�m�;ٺ)1��'���'�2�'���'Z��'���'�� ��Ωho�͙`N��@�^����'��'���'��' ��'�b�'�+E� E{��]������I����I؟`�����ޟ��I�\"�JY_ Kb��r��0�����I�����ʟ���ǟL��ɟ��I�T���e��=�1�L���$mɟ��ܟ4�	쟌�	���	����˟<�S��3�̺r�� ]�*Kf�Aߟ ���d�����Iӟ��	ş ��ݟ�u��
V������XO>5k4����T��ß��	�@�	ğ��Ο�I��l��G�Q<��o4+d���'����I��,��ܟ���ϟH��������8��<Z>�cD3{����Q�0�����Iޟh�I�@�ɜ�M���?qb�A�=�8��G�%3
���}���ƟȔ����T֦͒䌃�e���2t
���d� I�0�`�v�'�ɧ��'C&7X�DYJ�92M�,s$�t  ��H� `m����Φ��'����A;.k6T���1���b~ �C��ֺ%��xV���O�ʓ�h�f��e���=p#���	�:�X������S�&'�l��>F��w#��c���!]��L`�N�0�Z1�{Ӱ�l��<��O1��d��$k�z��Ȱ�	?�~E�@�"	��手�0�C��5�L$F{�Ok�GA�u���6`�	�JE�e%�y�_��&��zش#hX�<q��\�`/���bC�&w�T9bw����'�8� .�v�f���g}2˄%V��)g��0E�*�	Am����%1�^H�d@Q�a1��`��q݅��g�����!�r`ұ�P�/�p�y.O���?E��'��q�ѹ>��t2% ^�nѼ�؝'�7mm��I��M���O<B�a��	�U!,U�7�d����v�h�4~F���'����V�i����7Rzi�sƙ��j(���7[��}˴h��_ߴ�!��G�G��"v��{�>�X�̙,$D���� t�p&mU�K��ya�B�[�5���)Zi&O��h�V�O,2hL�'K�P���:�KG�v��R 82A�x4Kz�H<9�̊Z��iS��i0���W��X�U�,G�ԑ�"�i�U-��J9D�]�$qԈ��ٰ����>��)EG�m�>]p ��r�D(	@O��j ���Um� �(��ȇ�
�\I��B�A��0�f����L�!Zi�^HК�G�<�R�c��ˤ`h�H�O27�1��n�����I��h���?M��ޟf�p�dz"�=a��vD� ���O,��Q��O
�ĭ<ͧ�?���6᪴
����ɗ(�~�@̪�i6�5{C�rӾ���O��D�����O���Ov�����h�.����R�g��R����-�������O���|�H~���p �7o�;��D颌�+�j�` �i���'U�k���6��O���O����O뮔�zJPD��
y$D����H��	`y�a���4���d�On�D��S���P��J�Co����*o�mZޟ蚦,�M#���?����?eZ?9��q�T��_�I<䨪�A�i��'���0�'�"�';��'WBY>9��˯L���0a|Y�<�s���/����4�?q��?���+��STyb�'�����lڛ�L$Y
��?iXAr�ɡ�yY�@������I䟄�I90;��pڴf���b�̺<� �;F�`�5�iz�'q��'�RX���	J�S�(^����M2:�Y#ɗ�ndM�O+���O�D�O��DW+T�(�m��h�	�9�Vh��눈�����y���Iߴ�?����?�/O��$�r\�I�O�����M�R�qRB i�0�ࢇ�9ff�#��O��$�O��^�%��m�ޟD�I�d�S1�X0����e:��S!��q:^e*ݴ�?�,O���bP�I�O���|n�/^k���%��t��R����Y�7M�<A�FX1F֛v�'b2�'��D��>���8lS���^���+�X�\N�mZǟ���\��h�qܧb��,�2nV�.h�:plz��m��r1�Up޴�?��?��v���Zy2dQ�z��R$�T?~Li��OޤAĂ6�T i��d#��1�S���Z�aAh�fa���[�H��i8���M���?��{��EC4U�`�'���O�;F�L�w�H�t�	g,b%⡱i��'�.H*�����O��d�?�s6mֆ-�̵AA9��}���cӶ�" 'xm�埰����D�	���i����A+Q�NАh��
}m��ۆA�>���M�<I��?i��?���?�����I�jR�+C~8k� Y0��(&�x��f�';��'��~".OJ�d̼',`��ݽeǂLH��/4´MR!1O���O��d�ON�D�|��@3��v˺$��|�a��*�T�x��
�1��6M�O���OV�$�O�˓�?�a/��|�1Nn��1�C����0O�!Is�	ܦ��I6i������4�����z6�L㦡�Iџ�an�fa��v�Or��Y�R%�)�Mk��?������O���E6��˓i2R�H�e���j�r[���eX@ʊ��?9��?��_�vd�i6��'"�O��Ļ�Ϝ�5�݊r`�`~�{r�r����<��W�~<�'���|n:� ����l�!j�$)�B�;�L�`�i?R�'}��|�`���O�������)�O�1����'�Μ��憈�.��DS~}b�'D��e�'��I& &�e�I�5F�Y� �k��7ʘ+t��7��'iR<lZ�<�	㟨�S�?a�IΟ�ɂ�P|�A�.j�l�8� ̂f�ikݴk�����?Q(O�i7�i�O��xB>dp�S�g�&�n@������	ן���6__���ܴ�?Q��?���?�;f����݊T �Q��5C \l�Ny�P%` �u꘧�)����Od����,6�D�7*&8�@�3����=�ɢ�XE�ܴ�?���?Q�� ��K?-_�&xq%��mfL���U4}��6�J�Γ�?i��?	���?�,���a�ʙ,wR*�J��T/�� 3I��l�n�@��џ�������<A��?�NY	Q��'7&��	"
�`�����<i��?��?��������=ΧF�[R�_���\*T�Ձ?i�'���'��'��	Y�P�J�����|����G[�D]�'_b�'2Z��PI��ħ<b^��IU�S)���V)]0����ir�|2V���m$��2~�����'֓o�����h۟[}�6m�O����<97�Լ&�O���O��H��B+��=#�"�;ƨ�+�3�D�<���_���	�8T�&��$B���u���Z�Ls``��M�Y?���?	K�O�̃�)�+�l��"���2Z@�շi��	 L�@"<�~���#6	��LT4'(�!�2�	٦M���E��M���?I����'�x��'��<����(�( ��X�p��[��w���q�)§�?��B�j5��Da�y�-��ҦP��6�'��'��壔�4�D�ON�$���	�.ۼsg����f� 4
V �5�-���YMc�,�Iɟ��ɺl ~��t��xPċ����Y۴�?��R�O��$#��Ƣ@���.Wn(59E$� nRn��EP�c�,��ڟ����t�'����C��R�P��)j�4��*�9<�O���O8�O�ʓm��i�#�24B�:�'�??Zt�+CB̓�?���?I+O��"I��|rAcݦ)S.8q@�
����Zd}B�'�r�|RQ�T:Bn�>!��J�L�+&��7u�,� �/_}"�'���'��i�C�� w�Ӆ1�Y�5��5�`�7&�� �:�4�?�I>q-O�����ǡW���V@�p��B�=y?���'eX���Q1��'�?���W���E��(!׃�u!��p�xR^�|2�"�S�ĭ��!�@���Æ����kʻ�M[+O�h�Ǧ]+��F�����q�'�~�PҎ+-��T�׉	���ݴ��+{4�b?Aڣ�/(
�&1t��	rBu�ै������Iݟ��	�?�(H<1�&e<�H�'_�98��x7��-a�T-iD�i3������� �cgϞ:��P!�J�UV�ء�͸�M����?��w��Y��x�'���O 8�)���T��i	9T| bt�D>�1Ot�$�O���æZ�\,�'�4X�nHs��3k���n˟����ݿ�ē�?������3�b�PQ�0�����M�f}R����'���'2�T�\X�Ϝ
3����J��XKĠ�G�҉+K<����?N>�.O��r�ٜRb
y���G_g�\Q&lC1O��d�O*���<Y��
L��	_�):�ԲP"���`�ܙ<`��ğ0��H��Dy�.��DW�'�\U��fܘ`��\ sI� #^��� ��͟�'��8b��5���(#-�Y)���^�ԅ��l�A���n�ҟ�&�ؗ'Fn��}�&�{}v������.U��M����?	+O��` }���@��{`&M'nօqD�S6I��^T�L<�/O�P��~bt��=I@D�a�G�O�x@Pբ妽�'OL�{wib�P�O!2�O_ ��vu�+ݗ
PB�� �܃U��Po�ny�G	�O��d�h�Y��jD1d�7��� `�i���R�kӆ���O
�����>�����@��A�N><�aa̷x�����O>�����e�٢\�>Y���3<1����U���8��<-+��#�}"�'���Y��X��� �1n�8JA숒��O�����O��d�O����?>�h%yt�_7���ڤ���	�	)�0��I<9��?�����P�ũ�>;��LA�/[�����X���,�IꟌ��˟x�'����Y�^�K2����8Q"�¶s�O��D�O��$�<A.O�� RlW*r�6�ʅ�О8�3��ކ�1O���O��D�<��oI%�J�9.�B%#�M̢�z��~����l��[��jy�����$B6fZ�۳��4TYm��'0t��	ٟ���矤�' ��D+��Yz�(�S�@�H*������DE��mZ���$�З'fh�9�}�L��&��i3W�ѯ��WC̖�M#��?�-OP 1�ŐS�����&�P�;��Pz� ���8z�6��L<	*O��j��~zt  �jp��BF�c�00�!ۦ��'A<�Z0�a�ڰ�O6��O{�H㮐Jq��9@3�,q�N�91��l�UyR���O��bЂ��v?`�P͌�
�@��A�ic�`�@�g�@���Ob���8�$���Ƀ?>.=*�hZ&O�J@�e۷F������?)U� ��(��D xjN}�g��ElhhA6�i��'�r�N�* �OF���O@�I�n�$���5�y�#���h����OD���O�����D	�, 5t>-r2����M��^:@9ఒxr�'=|ZcZ��c�u��Q-�u� �����O����O�ʓ@7
��A� jyS"�.l�T���/j�'�r�'��'�剂w34<p��%��E*���8}|�y�(�����˟�'�@���m>�ڒ$�?}#�E�3��{"V@�FC/�d�O�OD�J���'�u��n�3o<��A��\��X�O����O����<�.ʓA�O�"0��eX�G�D���Ο�tP�Q��sӺ�1�$�<!��C^�m��i��F;7݊틶��7�ZPn��\�	qyd�1������	��޻<�LE��;(<@�Bd�]yё�O�ӫ6x&����d�p<���ķiy�ɥ"�d!�4X|�˟l�S�����x>��r�U5\pI3�U�6	�_�(c�.�S�{�.����O�@Fds�&_#_Y�l�#����4�?���?��'4ٱOlġE/��g=�A�H�''؉U�JҦ�9��.�S�Ov͟?*�yI�C�8�Mۢ%�U�7�O�D�O,y�B��r�I��X��y?��i�P�,�R�':�� ao�8W}�<����?��5P�C��/X��r�ʝhd��3d�iv"�	Z�hO��D�Op�Ok̜s7�Qd�/?�A����:�ɵ,�c��I����dy�
��.�eg�
~��B�G�f-�lA�2�D�OZ��"�d�<yN{��ecPb����Qb���yj�Y�<A��?�����@ (�6��'H�䠖�Q.nJ�Y�E�cm�M�'���'
�'��I�8������A"��i몉x���`Wܼ�':r�'�V�T)�\���'G��@bao�s��bp�0g:A��i�r�|�Q� ��>��7�^M@�n�}F�P�U	'.��6��O���<A�dG;��O�B�O�^yf�Z�Zמٓ�	4o�����n*��<)�%Og����ܕQ��yTN�0I8�@�N�1�&Z��{�·�M�QQ?1�I�?�Z�O��k��.�>X�Ģ�
�4R��i���#y�#<�~��&��oQ�HI��x�����¦9k#�ˮ�M#��?����#�x��'���	$��"��$�!/��cO:�� (c�8�
��)§�?QGM���"��ꞁ#�D%�F�'���'��(�b�$��O�ļ��s#.1[9�
�#U��)�w�'�	�4�c����֟`���<���b�'�l� ����
�/=T�ܴ�?!��'>�'�R�'�P��؝�ٳr
�<a�2jI�
�d�8����<����?����$��pCn��f��O�Z��@�֍s�0�{��{�	��������'���'�Z0���ƉF_���t��7D�J�X��Й��'���'��U� 9�T<��� � T=�yb�fԞA�"�J�������?1�����O6�DK�tC���j#�)��᜘+)��y�,`t���?����?�+O�c�%�[��
cҀX�FD�1q�@{�M��k�<ѫݴ�?i�����O��d\=J��>��\ �(�ٔ@�.��P�p�⦭��ԟ�'`ny�d���'$�t/�X�< �@ ͆���a�K8uD�O�˓^~=z���x{2���*��D�����eK��W�iN�;a�A�4mU��ԟ��S�����P�"���M:E���H�#�h���'B�V�yr�|��t"[�E��`8P!�bDT�b��D��MccCTi���'�b�'x��� ��O2,���N�|�%�����1������-��+����&�"|�����0W���
�e(���i���'W�R Z�ZO����O��	 �����7w�;RHއ%[�6�0���7U^��%>��	˟L�� *�ٹ��ڴN��)5� _�R۴�?9�IDL��'wb�'�ɧ5��3|�PŊ	C��*��_��$�"qV�<A���?Y���W��H���0�Z���K�0�)#@�I�������Z������y����R�ľG�})�
Z";�f��¥k���'��'��_�<"�1���	a>��ʳ���v}
D�����O���1���O����~�0:s���@đz���꒠�L���'$��'��_�����"�ħy��)1�G�L(�s����愂ոi'��|�'&b��"e,"�>��dՅg�x��`�2J��2�����IӟH�'�L22�"���O��i�4��9�e�B4i�TpQ��%��'���I��4�e����X$��'ST�9p�h΍'mpUQfE�� v�moZ|y�됩,I"7��v��'��K2?I�`�Xh��K�������	��D1�>�S�'Lozd��.�;��1����%X�r�o�e��1��4�?y���?��'z�'8�'C&6�H�"�Ιe����O*rj7�#�֓O��F�T�'�HH�a�J:)G �'_�\�Εc��uӒ���O����DCd�&��������1�Zti��C=�B�����>?�p�nZJ�	�y���(M|2��?��]��g�0�]�����v�DIG�i�BB8,�O����On�Ok�����8e�X�DRV�#g'�f��I�D��(�	xy��'�R�'��I��� 6p� (�f|!
��"���`��$v��'CB�'��'BR�' �	K���)0�w
[�k�.a0����2o�W�����8��^y"�DC��ӧ*&�����8�������G�r꓆?������?���*�Γ�N@�E�ho6��4F"+}�Y�UR��.��R�υ�_��)�')�����C2�����L����(8R�+��Q5H�5�fjF�q��t��J��M�oQ4W:����d���Y�_�)hw��._�q�cF�D͙d$W	o�R v��,th��יCRZ%�U��[#&=�FN�lO�-X�#XS���Z���66u��7�܏o
�Ѡ��0x�%sQ��t���$"0
r�RA��/w&T�BǊ�sX�q�@�˫7���1�O�D�O�����:<{��1Ц_�Sp� �fƊ�%V�|���: $MoZ�6�&�p�Ak��w�L	*AE� 25�����A�\�����=&8l�P��6��#J�cG�
6
q��m��/0�:�NÈ'�X!�G�~�� ���'#r���	%��,����!#^M�&"˜Wv"��ik�D�ISx�t"W ��@SN�[�j��c��l�R�*�	П�K��4�8��_3
��$������v	2�'�>jK��O��@�_?zX��O"�D�OD�;�?)��1pP^
�n|�Ч؍P���+¦W1�&�ؓh˟=��6�u2���DbPb��2Z�Y�VÓ�k�v�����d����g�x���ݟ�"=�7JI�Ov`t��L�&k8����Wq?�3��ݟ���4��F�$Db����Us�Sg<[ϒ�ɞ��y��G9dNP h�De�����"6�#=�O�剰<��4E��1��śZ^
 ��N~,�����?����?�5!��?y���$J5h|>1(7�[w ���:l����V M-��y���FL�yR��yB:t��A�y�P8��SB(fȑ�.Bd�x���Dm�y�NB��?��`��1�� �Bq���<X����d>��m�� �G��4���e$ʐ�
D�ȓ-�.)C�t����(وa�$ΓN�	cy�n͇���?/����޺89H���wtZY�-��B�����O����$h��m���Q�(o�]E.Ń�M�O�䅈 �/n�$	wA١C��{��d� S�6M����'E�̐h�Ǘ��O�X�@��'֩)Ĕ�Aǁ�Q��k�O�lzI�~Jt�� Ma��٠��*l����1J��<��u[L���@�DF�`���Q�]fR|��	��ēaJ�D��K�h�r�	5%��̓O�Y��^����d�d�ĮB��'�RD�>�v)��g�,on #���
U�Q�S��L�I�� ޫ53CP�5Ȥ�����w���ѕ��-` ��Վ#7���N�g�&�����{5�]q�%��B��x�թҾ��Ͽ�B̟bq��*.Y��0�J�8P(�����?q�O�O_�'�M�g6_�ܭ��Dl�'P�=�+ǆ �*�Q�Ń!8m��y��'��"=ͧ�?ɂ�����T��k�`���*U��?Y�6�҈�ʊ	�?a��?���g��N�O��$�}�8	0�DD�	a��A=&�R���	_NI�}9o�� 
�Pb�ݟ��C��*Ϙ'R��"5E�m�fy�fJ=F`�p�c�0d7r%��W4o���j7'Z�����Įb�|��<	�T�t��ы�mFL	a�OJ��?)�k��?�i���'�B�'Y���yW,�pD�qC
T`�����y2e�9Y��) `��I@���y�h"=9"�irY�T A#��Ms �7ĥ�#�RX%ag�S��?����?��4���x��?əO��p��6�貁�ڜ(|��!ꍀ
 dJ�I�)n}H
�.�
��.�� br�3a�H�a�%��\ �@�D9v ���	�L.>��Ț�+��աUz���Z)���@��,�M[��J#��<9�m� ^���Ǡ]��a|�<AC��\-N��wZ�d�� 0�!�<1"^��'"���e�>�����I��6m,0y�^;B�x	l�l`Y�F�O��D�O>E�e+�3I�x��Ңp����|�F �rNd�u`�	QX
����x�'oH�����E($�y�	f7�O�yZ�+l DU��Mǖ{+�ɏ򄏑|B�'D��R�� ڠ�p)��x�T谠=O��$/�OLঀI^� !5�H=঵�g�'�<O�@����>y�S/IŊx�T<On�)`�����ϟ��Ok�u���'��'��q�i�����@��X�Z��A��)P�-�f]��W�uh��D���v�P�m��NKB��6�NS:=Q�t��^����w�_
#�4�B�\��p�	V�F�%qk�!'N�����w��M���C"��"�kXzX��	Z�ai��`�"d��*���'<�dB5�Ґ/!qb��ãm�B���'["�$)ړT����ߝv~�(qf��k�l��<����*s�6�O�	��DXX�.�8�<5��YlT�S��O�đA�h����O(�$z>�$�S���'��MJGkˈg��A
�3L�C�'�����i�z��c��\AR���'jDt�CnE�H�4���3R��PG�KOazR���S%�Y���,Y1��Ӣ�<G�b�%n��zӆ�n�?��?�/O��"���|<����ˀl�*m8r"O� �����?X%(�y�j�T� �&�g�'f�S[y��R�R�6��'u�Ȍ����-W��U����rf��D�O��D�Ob�$��O��dc>M�ĦK�Q2f���蕊�2 ��"/p�N���ϙ���|��&Q�N��d��A��S$���8��t:hBq�.)��ɠQ
���զ����71mr��G��sx>�0nŒ���?q������iI�'k��3�A*y�Ĝ�'��x!�d�X�42xT
�K�z�7OHa�'�'�"}�CoO�>�Ωx��+bIt�`n�[�<c-˴��ŧto>��Co�~�<agE�%eo�daQ�H+/�B���.�}�<	�@CJR5IBC��%�(Q��C}�<���3}'UY#?{t��~�<YG(T�VP�Q��E�B��e��}�<��cR�?�ܸIb�>A^�3��s�<	���m<(���ᅴm#jyXa��v�<B�'x��qy��U0ܰ�����u�<�֠7�V5ѵF˩�H��KPq�<�&J��D���e�K��,��K�i�<9bhL�'�10�f�!?���"�]z�<�� '#�
�t#N�ty mc�u�<y��P�.k`�����k(�;��V�<��c_gF�1�ɕ�qw�9K�q=�'@��0+�3`�$��@� %+����'�`�䎰f���G	]�ۮ���'��jS-̀@�B 9�i��R���'�Qb�_�i<����(Z&
���	�'���I��f���5� Ќ��'#Z()�q�>h�5��a���'S<�k��(B���D �G���'|�,@ee
"#n�[�Y6�K	�'R�6��=,�Y8�<�c	�'�T���@�?]z�S��\*Iу�'�9�V���lo�Y�L��Q5�	�'0�Ujfc(2� X�$�"P{\(!�'Vm�]�<{�8�.ҍ(�@��,$�C���	"-ΐg����!~�CQnQ�#�A��H�T	N��� ���ɓ�N/kbfy������ȓ: �Bh#\)&� �$��I��Ԗ'p����� �&��W�O�ر"L-V�*p␌�/r9Z��]���`�NIh��,O?�8/öqtAB'O�e�d-��AU�#p2m�'�*,� cA'N*���OL�z��ؼ]���3�5TږřuŤ��H�h��/��в$ތk�Q���ų�v c�a �Fx���DK�%d2��a&��h��ٽ4�\@J>��e�:��1��!�=[b���� �h-�Uo�(�b�<���b����<@h,�Q7�h��WG�	�b%`񥏈�<����&}��[?Q�x���-6y�Ƀ0	H��?%?�a��Q?u���˳"K�r��8�>q/L�U٪����X��1C�Z�'����Q��&����5H�%�K��$��D���U��OP���1@�et剬;�x�4�r�H�w�f%AC'�^�̣,�O��ؓj�;1f�M���9;�X���})6�g.�4 ��GiN�e`��<�s��Ra�K�Q;��@�C�F�[�%F��0��a��K���Z:�`��F�?` a�ٜ�(O���	�X�*�b��V��!�;b0�-��ۃn��"��ȵ���bW*F��4Lѩ4ɇ��1�C��Q:�:�P��Z��	=F刭�u`�	E&�U��K��j�l�n~r�"g��� ��$Gv2�إ��5�(O�\�v�'M�����2�ڡP�$���B�	<��ĭ'\�4�w�FZX*�˔�C:�~�оo>ax��αB6���AD�8����(����)`럨
�D劗Aʭ �iz���k���#6�9a���2JLb1�3kOzP�x�?��⥡��T�����-�zi�&���JFy��z����%mvzh�"�`����f۬\� ��_XS��2�I�o,���?��o
�Q��}��m�5Lɶ3`������Ɍ!ʶ��cԝE�0���	Ҟt6��i�5nbT�c ,(��8k'�ap]�?�$~�q��#�`@sQ�I�x��	R3���#�zK�PmR l�!���"1kϙxr�V5�)�'���',�'��r!뉎D����� �=B�y��	W2��J���(O���A��!��I�,38ѩ�P���O
q�Wi/�)�3� f\���'�4�r�-2/�Yci֕ �<��F��5��,�^7@�ż2�� ]�	��6�j����D�05]z��Ot&��X�>X&ܢ�I�R�1��;P���*(��1�ɬp�؀ &J?l�nP�?��ob��׈W���HTa����"d��C՟<�A: V�Z @�!���iL',k�O��eܾLa�0~�E�u���dP�@�m�x.DRD�
�\��J�	�-_&��*Q����aA���]�2��GFݾq���#R����=cX��C�,��<�'/UB���J�
WP��p�
7.����V-��(O��B�*����t�n���:6����.�)vŒ੒M�K��c��ON�)�O�|�\�s-(�	_u��ݑ|�`�����P�	e ٶwqV�'�X�:�*\CH����*H�E�0�h�5�ԟ֥eJK֬9��m��1���[�bM
&�˓��gj��ʊG��pyi���
�sWG�/�L�X`�ϰH*D��7����N>�O�ݔ�yg� /p�4��H�*<E1`�t���o_q��E�f�C4C �Hc���ˋ�,��1A���wf2����,���*^h�1�Ix���I6=b�.��q�O�"Y���Ѓa	̩�q��/:Δ �%j;����GC�QQ�N�}�t�+!�w��`j�Z�o�F!�ҊU�āg�ªZ��Ńc�&��T��f2@� ���t#�K'8U�����@�3�6ys$Y������N������	⺐�ŭ|����'7V��i�rJ_�w^y1D�Ӌ�p��z�]��z^E��D�Ot剞y�z�j��֫9�Ar�^A���S�ǈ69h��'i�;dw�(O�I�~P�nލ� X�I��hqC�Z�M,p����(,��d����6w���I���/��">ͻǺ�iU��X����	Q���O.�a%$�)�ӛ#*�m��"J��p�����#M}��;��'4�;��3��`��J�Y
葪2	�k�(�!�{�E�?��cC����PD�D����O��+ #�����w@�$�dYP�	,'d
�
��T� �\� �������Ñ�L�{x�!�d۪P~xq���O�e���	"�����)�����	�z�p��	��MFfeX'LXK6�"n6�Ҵ�،Lk�id�P#u�'�K��1	�OW����o��2��ճ�A
�x$�s	�Z�r�zFÛ�u:�s@�V�8h���Q%��'��d/�S�������뎦C ����o�Y�j��S^X�����|Qt��0��P/BD�� �2E����,����'X����BE��(�+���$��9C�K�'n�*-ѫO8i;Q��"\+�HOZ0ѡ��5���/��](ly�O��r0�A"�Y��F��]	���!�����ҝtZ�HD,/	�f8�wE3ړn���Y�,�'P�"m�'G+Qg$�nڛz��D� �I�mzd�j!✄]��g�'��=�ǤZ��̙��DB�TQ�|P%��38̪h��'I���$���P>2��a��d����_�����	>a�Q��2���;F�~�����]��M�ЧB�J���ēo>��eaƥs�d�h�%}��'�i�@��4��;2j�b �|b��	ƾM˶�&(j�J��<ɲ�?�)h �Z"vB-� U��)�ԭA�@��9@���M�"�E�4*�Ѱv�az BsPr���%y��k
�HO�a ����~bA��<c�ŖO��iR)P�/m�m37L�~p�M��'-�4$�3e�r@Ȗ�34�&�ri���R9Q2�O���'t^&諞w����3,��O�µP����u�^Q�'{���ɏ�Yʩ�-Z�\�kVi2ғ
�y��O�Ce����)�$��U��M f�^-D_b1��ω�:�ў��%k�0����S���(�q&��O�N_�]	�h�bIQ�#���E
�!1��d��n�8F�^?ڤK_���dv�Zk��}���`�r���D`�.]	eE��O�b��DO.Q�	�2�O�#<1���� d�6�,�H%9�B�C��|"�P6��>Q��=��](�Ǎ�.4H9����8u�:�a�O�=�Ok8��;
D�X`��8R��Q��Q%+P�}��	�
֠=�&K��]�jYk�٩=:z�P��P�	�)��'��������ا��0K� S��	)��S92}��e9HG~���N�>�HO���Eȕ�\��ö��c?\�x#�OL�"u�8?qLh����z�<| rF����gJÞP�������s"\�8P,ړ\�x�R)[���t�ԭɛb:$%l�c�*d�IǵN�4{WD��D9p�I~�'����%�Լ}X@.�1/��\���-J̙��'�7cV8�c��lt��h��1�f4��>x�Q��'I:M�;]�n<���ķA�H��g
�=t���ɢ^:L�q�ɦ��d�/l�� ��ָFt㞐PBcL:�!J2��3�yc�N�?a�?�^1!M�,A���
ܱ>�xa�'3P;��[0G�����ߟW�LI�}�'`�����6���8�%E��B�D��8`�1�~�j���c���'^<	��P�v�"I���X3Fz��S�@��jc#��8�(Q�1k�<�|�i�uceh�Ւ�X�8ɣ���0!R��0��֯*�v.[�P��C�0i]Q���wp��%�lB$�рZ�x~����]M?1*ɯFTb����ǟ�ӄV��y�F!_>��F�ل@��םL\`������N�7BY�A��ǽ���	� 4�A�a҇h��L���1k��ja�
+<�heA?$�&|��c�j���4 �+�*\t`�0��Ԁn�ԸZ���!4&u��֝��܋�fκ�O�S/!��IhS$ÿ$���A�Ƒg�&b�d�d�)��	��v�2�I��[=�u']����J�I�>�(��$;ZkӣS�\��u���C��2I>�OqO��˚:���F� q���xf��`a����K[
+ĀӆM�'v��<���p��&cz�XkP����#_��pd�Q-l�8��'���%d'�y�X
�uxEm��{������SAQ��ɛ�^�tzAe��;*����S��$�aO�u�*0�d "`^Ь�K<aB� @��[��D��|2 -,aSح`�H��<e�A�ç�Q����'�|�+�=~�����o��ilV�Cش���|r�MԡЬ�#�5��ܪPM�wYD�O�7����:�j�5�d9�N͚���9��JDB(~�R�b�O���:�5N��$�����Ƀ5fؘ��SL�R��}p�G��^<Xa��I�zEy#Q#�'G�dI�Q�3��?�n�� �M�%������L�s�\(����)*Mہ�Qp8y󥦕K	�AÔ��*Lم�A-^�8x񡮅!�yg�y$)� �/F��=��aF���'@�a�4�ԟZ-2�띜:����M��j�ʁ�/@�a���'�T�QĦ8�����]=�����'������:w�:Y�f�v$ �sD����u�$�DָQ��k ���'Z�ݺ��	L����P��zM���ύ+�ؐ�b?�)ڧ66��J�i�	3�2�X��G��B jcK��D�27"ӨUl��%��(O���m�g�#�"��9X�(�ODT9�)��؟L�Eۣ���Z���/[�Q^~,
lL�]:��Ey��G2Z���'K��~-d\��M�Ԥ�<:} ��5 KR����"�m�#�jyP���d��̆�!�H784k#'Ϣb̾�[�$�t����a�::(��gY�I����N���C�oA&_�"=Qc�D˚�
�����A�'�<I��A�@jhi�D�:ȂB�5<@,iV#�*z�Z=���<��̏�ez�H�8����1*K�IY��A�$ha}�͙�up8b�#�/[�={E( |����T��2��ClÃ7D�Aá�	�y'��/T(�s�nE�o+�U��^���>	��V�GBZ�C�ᆃD�Ӱ�/cB�q�:l��9KB剓dD�Ѵ�
"o�B�u�,]�6D'a~)Ae�XI������9&@��0  ������Ш��H��X��3`��9�/��� Y1Հ�/6����w�*��Ě�F|~����U�#�T����ߣ ���XL��<�oZ�r h��f� ����7$Qrm"BoU -T���8l��x �)�F4��,Oʕ2D�L�h`�2-�p,i:W�L	�̵l�FX�8�󏔩GBN ���@(�Rǘ~H�x ��<0h�B2m�O�8FyR�p�ѠRhU�N���K�j#S/h��s!)���#?yC��+	�ph6N��jꌈF���rQ��
�����6ʓJQj��B���2�P��*AA��mZ2FF䙧��Z��j���A$D%�OV���PȉI���X;DXCSg����'�)2��&����-�y�h�'Ծ1�0�O.9p̙#H�.Fj��t�O�����.Ț�pIg�X�$���@%[-���B���H𭑿��O�>�4q�VC���h!�C�	ք,@�� ��~BQ�]BN9�"l1��$�+TB�M��(X��`����	��xY�D!�0O��ۓ�ɾd.P����VD�s�Ȁ%2t�9j�@���|1jqHTZx�8h�L��ok|0�%TI@�Ik4N@gt(��Ri,��D���`���
���-
�l��'Y�IZ@]�ȓ�5�ӇW�qC������r�ąȓ!���@i͸w�0��5!�*�vȄȓ1���9%NW� (��� M#5�R܅ȓ9=�����*6�����f,N�ȓ"�,����+T��&�<`��Q�ȓ3>�A2���LU@�!R�L"��ȓN�y�D�91<�ɡ�R��v��u
�I)�@\��I�lo&ՄȓNș��ͻ%=`jp$V�{���ȓ\�ֽ���.����%�DH��M�8��d��.y�Z �����v�T��pl��)Jd(��%�a��H�ȓ2^���<V^���+_�����ȓW���b_Qz����:,�`��ȓ3v�AŮ��`p�0���X ^�N��ȓK��Q��7O:�2@E��}���ȓ5��9!�Y��-#�v�n@s	�'��`��RQ��{���b��	�'�v��@͍i �����>"V���')��Y&�ۧ�xp��.I�qZ�(S�'� �� � ��<�� ǡZ��� ��� �p�/ŚA����Ī�`���"O���FS V-�\�v��'�� J"O�Tf�' �Y��h��r��[!"O�8p���j���h���{��	�r"O���H�=$�P4�î(�����"O��
7HX�[V����kF��*��
�'��6b�?��5Y
M*g����'��yۀ�Ln��DK�,K��5 �'�U�4	���8�%(>6|2�'m	Q���hmQ��]?&���	�'ܚX��DJ��%�4@�)&��9�'�d�S����iVı��G���h�'��y�� ьz ����
��I�'���@E��0�~��h���
�'�V���#�PJ�آѥ0(؈B
�'c��c� �Q��̚��/����	�'mz�K�/��w_���qNV�
����'�
鲆�>c6�A�W�nn�3�'��P��M�q�iS1��1;����'��d@����|I.�J��/�L���'�B�X���4qԽ+ǀٻ+y�u��'�P;�D$Dv���>&T^q@�'�^a�v�J��مk�8!|��R�'�	���nۨ8r�C�vHa	�'��p tO
�H�|a�a�j|��i�'g�8��ј�T��*�d��Q�'���5=Tq�wHd��8H�'
�d��f֛6M ���	?�:���'d|�	����Jyfآ�[;V)c�'�,��%�Tі���|��z�'U4�Âh ���W�y`���'^䌢4��/+�=�@�q�
-p�'���* N@x�Gd�zЬȲ�'�)2�W~WL��w�G z��(�'�Vh�҃��<��8"�s.(�x�'j
M��ڏy��@7L��_����'�>��cϒ�w7���7��9(6����'�Ȥ�U��x
"qG��i1tȲ�'�Ȱ����x��HVDa�@�j�'��Š�GM�E&XR�ԄZ�'j��AB#�)�@h1EjW�Oe,�K�'���ц
@���-X��B��a��'\4-�Q��R�s��?x`���'Ol$8h��	����͎'9o��j�'?tm�e(]6eǴ4�"I�(1�pa��'�2Bdl�_Jl�A���$�8B�'%N�x���y�f�q�^����'Q���,��~�&�2D%_4�%3�'�2��n�16%�hT��a�^[�'� x��e�/v���4��k�dq��'#l�赇џ4�F�z���-9XC	�'���pEZ`1D�G �.��'Ȯ�h lҬ6���0K�v4�	�'6�b̖�&`x��N�w��
�'+�0��$��\���@�I�-��'~��W)������$��'�� `��Q"9�ı�2޾w�>�z�'zqj�o�/3!��##Y t����	�'��<�K>d�:a�E��6똝�	�'���9T)\�#��`*�#X�i�'=����O}T8ऌ�"�Bp��'hT!��Y9�C�lV66���'� sъ�?�|����8t��}J�'
JMZ!�>9��s�i��sDNia	��� <QB�-�z�����U�9��<:A"O�%����
a�dH.O8����"Oh̸@����؋W�6F���"O���R�P�L�DІ� 7� $ґ"O�,��*S��={�)Ֆ��\��"O��׉��z���i.�i�	^�����)M�5�b�A��[�B�#O�!�d]�u����&Z��H� �'�!�d"l����cN�\��}�o��Q]!�D�<h* Y(%�ǥ8��!w	GF�!��>y�DHlC�9 [�+�!�$ y�0��ê��)� �X�wZ!�$��{-^��7HY�n& �E(�xR!��2<��g �a�8D�V�_7!��`�l�x���=ʾ��S��)s3!�"t|$"V�ҩ/��}�U12�!��Tx��-E�F���i7Cşao!���X��ݥ5�r 8�BT�!��]�C����p0�/\={�ay"�#k�� �J�z^Q��	��p4C�<2^��Ac �f,XyAwg��O��=�}�Wmύ6��f"S%@{J<9�%�`�<a!g5"WH�ڤ�^"<,"Iɠ��f�<��̓KjJ�1�K��nlsM�z�<a�I�<q�r�a�H�J	K!��P�<I�e�C�.���.�^<��7c�M�<�+��e����*�H!B����<�¡K�8͖	� ��i!z��Cs�<��؁O���� q���	pi�Z�<Il�-LAq@�P>S���W�<� �"�ȓ�@հhܱ��i�V�<Q���Od�p�B��L9l��ue�z�<aƤ*x��� ��1��!�r�<���L&R�8�AV��X7�I��m�<')��*���M�0p��]�<I����ٳ��67~a���\�<�un�'rE��c�N
;b� 	[�<�CbKoJ��cC!�o��:���[�<qVØuB|��V. �0s"�*`�r�<��ʗ�,�c�䐟bԼ�0Ŋz�<���۷S�D��i%�0q��t�<����&I@�@yר{9t��n�<����eę���<0S�$`�<���M(E��k�E
9P  ��[�<�#��+<��դ�Q��D��{�<�RfX���2VL�g��]ʢϑ}�<)���f$�^�J��|�<���#6��D��Q������Zd�<A�j���;#��t��J%Ȉ]�<�t&F4=@��B���-�H\����U�<9�@p�DI�B\9�6��I\�<�5��L��=��I��g��%$%�_�<�E#��?!XH"qGB42l�@��� C�<���"�,�aOI�ZP}	$�N�<��gտ~��=@� r�i�ɆP�<�ΐ�ggvIY��
t�b��
�@���͓�TY�G�d�J���l�K����ȓ�����]d\@�JF��Lun�G{��Oo"a2�k�4�,Ɉ���$m�M�'���G�+x��Xd��{.��k�'�b���M�,88�K�F�&^S�!I�'d:�OL�p�ɲs�

K���'�2|A��Y3&pq�jH0u�N��
�'w���r�	8ޒx�F�V9aƾ4�
��� P��vC��zt����
;�ڄ3e"O��	�W>>|F�p�X%8�)A"O��2b��
N���叿X@���"O�6���P&�ȡ�Y�\c�"OZ�� N�/�lx��"Z���Ѱ%"O�8K!�۫�s��6v� ��a"O�MYWEˉ�h�H#�.�d �"O�U��t���s @�Cu$,�"O�9��#�@���aR�tbj-`�"ORHlI����f��s�e��"O��@��u��j�(R�Ba��"O��P�`�B���+��_�Rn�[��)�S⓶O�@lB��Úx�݈�cƎFی��hOQ>�1��Wo<|�����tXRh�$�7?��ᓿ)�h@cC,Y� �bj�:I`C�I4����R�D��I�Y.G�B�ɉ{ڜ��	@�%��%*u�֓HPC�Ɏ3�=BkM�O��E`�e�t	B��+(d�����h��9FaR4�C�I�\j���҅ɄDg^`��Q;<�C�ɝS�F��\<`A%�v�
Q��B�4z6�1�N�(&�sD���UiB�	/	�M�o,a)��a%F�$V��C�	3]o51@LՇV�v���1�=�ç,��B�J���xS��*��}��|�����876���늷9R���'��\9a@jl�lz��	�"�Z�'�f�I�k�`��3�h��'�( �����=%��
�%I�~*���j,�S��?�6���u撈�3G�q��T��ʏX�<���?pq��$O�h?�ؙ0�U�<�&ݻ<�r�!3�/ny������G�<��-���𥠢H�=[f�\k�-D��h�c֌x�\Z��TOv��jPD0D�|"WJ6N��Vu�����*0D��#��Pz�
���j��n-Jk��0D��j�D�)��ƓpS9Z0� D�4�� a�yƆؼG8��sp�Ƕ�y�G��VҀy���R\ Eq�-X�y�̓
E��l��hG)P��1�E�yre�(\{h�Ο*Z�� ��&�yrH��&E]cR'I���\B�)ҝ�y¢��n�^l�u�|����	���3CI<4���spR
�M��y��ͥ^-6L�d�Y*f;����J�y�-A#�l��5bn�l�rfg���ybŅ,Nέh�ei.���
�y��~����ƙ7\������y��͹r=��RB
]��q���yr`.v�虗��l���#�"�yB�^IF���"h���ʢL��yb��2j���b%��[&f��a���y�∅I� ���1S��PсE��y2��f}��^��8�=�y�mD�~w5Y4��c����sL"�y"'_�H7�����	��`cG��y�����;���-v�)�SJ��yB��>4��$���V ���&����y���%ع�M��N�l=*���1�y��/��B%��Dܠ0gÔ��y"���m����E�ΠM�\�ZfB��y�)�!g�ȨZ4���v-��3)�.�y2����qE���" ��GZ��y��V>ϐ]��ŀ�x�"��Q�+�y
� "U(�
���hL���1�򰛖"O�!	�@,O�R)"�	�JT�Ё�"OP�[7N�6ς�x�%T�-�A"OBU����,����#�кd,t9[�"O&�p@���/�L�c�����"O�T�m�Z����xv��`Q"O���v���A�0�N�ygV��q"O��PC�9{��	�m�&k\����"ON��n$$��(C���0F��"O�\���ׯs�2����)_�Bd[�"O�0C�Z:R��sIG�y�敩w"O�}0t��43ѤHQ���?���9P"O�M9�M�<9
#)ߤOK��%"O�x�����5^����'!�6��g"O�Й5�_1GL�0�jؿn ,d"OV-���h>�]�*�@U� �"O&�zc˞CIQ $���ZC,���"Of`#b��u��R"�	p�8�K"O,����3�De��#�P�"O�Uc&��'�ēÀ޺X~X("OH� `ł0�x%�q͓k=�	�"Or9ҁL�F+��hl�[!��x�"O�!�ucө5��X��j�>m��ٶ"O^dQ�b[#f����"�.n�@��!"O*q��.܉e4b��&���'��q�"O6��(Ψ zZ�� �9����a"Oz*EFM�:��i��������CW"O��ГaD� ����L���3d"O
u����2`TJ3��'|<�"O\����XpĲ�Wc� y�\�u"OUb��īz&���$&CZ�m�"OҠk�@���e� C��
�"O�Y���#�%�V�=�.�!t�S8�y��.�����\�*�ܩ�skU�y�&�<aE�T�c�;��b3D��y� ��H�N䂀 ���0�CԾ�yR�1�~i�D�1��]��,�ybO�>z`,z�OZkp�5i�cQ/�y�GW�Db<q�7���j�aS����yr��86P�j��C�[L���B$�yK��;���b�@��(q��S�eE�y�	D:x���s�N׫l�=�`��y��O?%�e
�M�8w�=���y��Cc|@x.4�AS�H�gf]�'�D����8��M�M�Y�r���' R�J�i�	\0$�p)�>�
�'����#O�?s�E��_�ԍ;�' d�$I�)_<��C�V�X��� �'|�IB+�+H�t$J3�Ɂ"²���'�@�1�2H��؀񥖇8t�
�'Ty�L��*B��7v�̱��'Nv)ȓ�G�|l��q�)(�'V IG��9zy��HP�X����'B�(C�-P�j�aˊ!L��8��'g�}��E��'HL�"QGDHQ2�C�'8�@����r�V�� ,U:P!ze�
�'qd-�MV�&����͛H���	�'$(,Y�nU�4?����qRV�	�'�н3�����MR� ;�ѣ�'�:��Ũ�V9hTk�̄w�����'��`V�ۃu������P�k𪥳�'�D�G��A��`E�_��	�'ߴ��P/P�ؤ�����c&y�'9ީ[&f��3���(2���T������� �({ ���'M&i�TcO�K�b��V"O0m�R�t(D���n��$"O `��,�	 ��h���>����A"O(���<6�֌�pF|.(��"O��c��ɓlL��a�D4T�D�r"O�}��N�*��L��W�h��p�"O����� t`0J�`��!"Oz%��m8jŻ��)�q1p"Onٓ��Ǆ6J`-��m��Z�lMXD"O\�)NO
Ѐ�+棃�=6���"OΠ�f.�F^I��a-?/lE[d"O$<c�c�!e�p@Q�elİq"O%@Ҡ"�"��c��7�,�g"O��b�jT�b`��=�xtð"O���F��2W�D��A��9����"O<���Dܽp���� �T�u#�"Of@)׋��f�>m[W/�$U��m�S"OD��D���bLpT%�B�6�x�"O���
�W�
{0�	(P��mX�"O~�
��Y1@��Bː=���!�"O:���Q�p�������!	���"O��ˤͅ�5^tc��^�j\��u"OP�ȅG��[N��q��D�z�#�"OuZ�Ϟw#B�+ЪS�Q��� �"O&�a���]{�k
d�n�b"OyEb�0CJ��RW:��lh�"O4E�� & ����7?8�E�g"O�a�1�X E��|У-W>|2��#"O��ek�\�"<i��&u��R"Oԋ"��/`�^Q�)C}24Z�"O�brS+�I�e��7���U1D��BD]�Zd�9�T%R��`�C0D��;4�p��!׬L�ML��)$D�T��#K'oVa!����lx�&0D��Ⓞ	�W��D�6�B'G���!�@2D��N)8����K��5=�X�6�+D����Ɉ+V�@Dj���::�)��I(D���ʃ��8��,�+�����3D���E�C
[O<�	�/�77�Α
�3D�P3̏7Q��P4�J�U�5;m1D��I$�Ԍ0޲�idCӴj(�q�aj1D��JP��1AAz�H&�9C�Xa��&%D� A�)o�X�!3-��=�@ZǪ=D��1��A�w�������`�&��$:D���EB�(*v�P�]�6���8D����l�+�D<���(�o�$B�	�+��� Dàc�� [��B(8?�C�I�2̮��(�2�z����$b~B�:lm4�j2��%���cl�9^��B��5~�0)���c�+�#��X)�N:D���aLڳ2Ln����]����I9D���bi�$5FQҶL��s��AG`8D�ܠ��c�\Zvd�@��+�/6D�T� C9Q/�WOYi^�@���/D��S�@�A��t�P� ��!��B�	�F�8�6�Y%�&�Qg�͘a%�B�	+]��3�̀�HKYH%�J#�LB䉲�8ˤH�+���p�� Q�B�	�)B$�A'�w��+�j_{�JB��,B�t�A�K��움#ܠ��C�I�=g�������I�>�bB�I9���0pg�>rP��'܃�$B�ɹ�z%ە�����b�>��C�I! �݃�l�k�5r�dY+ ��C�)� ����k՘�p��"�ry8d"O�A�G �+�:أW�x�M �"O@Q!�I��i����-("O�K�f#�:���AN�:>��A"O���A�6�h�`@C*����"O��)#g�0u?-J�=?-���"O�xE ��c*U���'<�BU�r"O|�T!�������9u��e��"O�=R�lJ�Q6]��P�`�R��"O4|�qи3L�X3�.ǒ�$�1"O��� T<OX�4��Y+#�2�"O�i�d�-N��+t��$��"O��)��KX�y��.��\��"Oz� �k 3y��
H����q3�"O�p��.^<���G?!MJEJp"O���P�\=3L��rT0�pW"O�(�6n�#���FT#5�j�1""O��J���&���A���j�iE"O��R�
@�h)�dG��,<�5{�"O޹��GƳ!^*$@�C�H2��"O��p��X9g<q��z!� #�"O̥�f$�L�4p���.���#"Oʄ*��+=�]�$�.4ppj�"O�`I��ȚI82X����34"O�d���5��9�֬@!,���f"Ol�0�U�S�z� �
�j�h�"Op(�a�2}I��` ��uy"O0�q1�׃9Hlv,��`(9��"O�50�)Ъ;`ye��.jLy�"ON�0D��de��WX��� ��y�i�$nh �[��:$�@I&�y�'�;O4V �S��6�T������y2���*��H���@�2d�/F��y�d�)*��
��눩����y��wq�XK�	}�����HD��y2Ϗ�u�^���Ǟ�����#0�y���t���mیl@� �S�I��y2@�_f\���O�j�-Q��\��yң �-��IP������ O
�yR�_�n(
��󌜞5\��ܸ�y"���Z:��jtjH�c(��.�ybDR	[i �PA����"����y�A�WF����$۫S�Ƥb0͞�y��Z���9s�ޥF'�!�Ȑ�y�@#Z�,Q�W��Xb���y�\�(ĳ&M�$$*�2 �y�c$=T�����=|�D��pfC��y��B/	x��g��oP��P1@Q��yRm�}�R�Zq��bfRd��B���yB�
�l��U��.ڦS.�d�4�y�LV a��c��e����W��yoR"����S"��Y���ֺ�yb�6#����)�!k���e��yrM�?o�y tI\1I�U��֍�y�c�,b��#Q�3�B�ρ�y�aG�	+��;樝���%�C�ِ�ye87��,S3H@�׼�a"����y��3A��RqEK'kv����H4�y�c��i����-�#�����ؽ�y$R;)�&���,�
!�,�! ͖�y�WgK�Pr�j��F9�t+т�y��J�n�\ �����h㐍�y"I��_D��W���:�e�!�yr��3p�2	B���QV�Kef�&�y
� dSc�D�>��u��40�Z���"O�h5��x�8]�$�-0t�\Iu"O�-��	�욥dQ�3�|U:r"O���J�;�mR�Z�L:P�"O,щ���7<�`H��6qiE�w"O���֦��9�ТCD�*
Z؝�@"OP����Q;�X
�3AL�a"O�)÷��~��U�qA7"6���t"O:��îR#`Gp ��Ư&)���W"OX��-Ip���c��G�5	���"O���ϜV�^�Ȱ.M�O����"OrI��_z�P����g��X�!���=�.u�G�L
�!��L,i|!�D�=�H4+�B��R���H"��R�!��IK�j�c���ZG��8AF^�;�!�$�"V�=3f�I#
nP���4U�!��
Y��ytɇ�9�8)b�dm!�d�q��˶�5Sn��ڐ�x4j�'����!�e�И�lτtT�ػ�'7�(BQ㓫.�qh��\��`�
�'�`+PGʭ���m�V�Y�'��mҐ$ԋK�|A6��[ұ�
�'�}�F.3���E�IY��J
�'�(����;��B�ۙQ3h���'E�[k�4�DA�VM�NBn��'��l�Q��h7�ʐ�I"R
Y��'5�(��;9��i��E0}oHLh�'�Hd+�L2Ʉx0�Ǆ!;�Eh�'��Ա��\�̍Х�ї����	�'��Peۓd��!A���~��'�8q`�.J����jzkA��'|t��׉ȍ#�]J���3�԰�'O4��ǐ�^0��FL�b�̤Z�'���j��U#``�	p��X�\�j�'�veȒ/ĩhĐ"�Q�>�f�
�'u�U���%'�bi%��=.���'��0�g��h p�!-�0h#�'!�P[���_#�8�v�P!+���K�'�d���ݑ�I�����%F%��'ؾ3�K �2HB-^W��9�'��E;P�7/�`I@-ЃN����
�'^RIzBO�8EY����`����
�'d�y#�'�cG���/7��x�� [��cf^�m�t��Q^�+�"}��&Ŝ5�6��3�\,���ʋ@�F���e ���됮\�Q�%�, X��>��h�qc
;��di��P !�2$�ȓ3��I��[w�y�*ޖӜ��/�`dh�|���pc�_J�:d��7�����O�����v���B�����e	9,A䱈2����u��[�.!B�kP��:ă���,�^ͅ�c��[� X�J"�l˄bέ�T�ȓB����o�g�2Y�Ceϥ$���ȓ7q&�A]L���Y-2&b@�r1D��Cp��Z��Z��ØV�2xRp�;D����ҍR�MsCL*Hk�+<D�|
2.�)[ܒ8
�a��Dm����M/D��W�K��+�cJI�$S�2D���@CD� 1�"hF�SwV�� �&D��`W�Z�X�R�#CAZ敩J$D�|���S ������M�Ԉ)�զ&D� A��1�,�K�(M'=Ѥ��b(D��QR�84�P�'Xnל��U�%D�� \	1�h�� �zU�c��2����p*O��!shߟB^�iC �7�l��'��R��[��1��mݵC��5	�'�0� W�I<r�R�z'�1>މ9�'�pq��I�!P�=���  �`��'�>M�&a�ZO�	�&�
�'Q��#�܄=���ha�h&�#
�'�Th�ү��<܈�ph#�7"O�	���ޫ	�&,�G��"^�+4"O��kF*��X�))Ď ���F"O���A�'9R�cB�F�1����"O�HQ��?>�����J�Y:�"O��R�ɳf=����BI-Ѱ"O
	�E	A��>|��+̦X,,
�"O9g��G���"*�.=��	�6"O*R�*�.!U9��&��<|�X*%"O�R�����j�N�"Co��v"O��"���J�r�P��%q:�h�"O�<QWõ[��P�D�'i9М"�"O\��� <%>�a�ǁC�$��w"O�,BE�GVp�K�G�r�pZ'"Oj KDD�=��u��C�G�~5�v"O:�)`͹S� ��Rh�"��U"O@eh��R�N\��Ӗ�v��5A�"O���b��w
13C��1���ȇ"Ox}0� ���c�գY�\|��"Oĺ��Q�J'Z<9�l� }2�s�"OHh0�E�P[T��@�t���"OæNX*�^@Q�-is:	�u"O�`�p���M�v��k�(Hg���
�'�8�����$40�=+���&3L ��'\���)U���y�\l�'L����F�8�k��D%��
�'o���Ĩ� R"�x��
C��@�	�'h�#d�3(�ʹ4�Xc�X�'�*(:7IE�Cb���6K]�U�p�C�'��p,	!!��e$­Tܭ��'zx��+`R�ӳ��1!�)��'��]a @�N&�X��=p��l��'�LĚWe	�5��c��ʞiJp$�
�'D��)�o��$D�,Fe�i��()	�'4�e�t�k�Ћ�K^Y 98�'����fɯ`�6(��R1]_�|h�'a�� �˲&���0�/C-Z ���'�~����R,҈��D�R�  �
�'7:�j�Ι-�tY�F�z�uh
�'�^��t܂9<�H��@�
�V�
�'�)R��6JZiz�U�U�"�0	�'\��Y��8�V���.��c�����'��Xq���	pG�#X;g�07"O���$Q�p7�=�E�����"O�	�&������V�\���"Oإ*���0�U��!� %"O>$�F�ޘ|C�9�J��1`�"O�l &�+z\��7*�0<���!E"OvQ	qZ �!�ɘ7�`�@"O�P�`�+i½[p&�b��Qp"O���0��do��0�
XJ�Ce"OV��97��ӄ/L��$�[@"O>t�6�T;$0qkG�f�#d�Jx�<���y��-P�a�?�9tN�g�< C�O<�r�B��*�ʤ�FVc�<�g�͞#!t�"V��\�P�X�\a�<�RX�I!�ä*�r�3P�s�<� ��r�a��0lL`�m�O�T��"O�Y��w�z|��+�:�Ł�"O�	���<�h���j�$6��ݒ�"OfH�,܋oo��yW��5&& hh"O�����$B��J��Όl
��A"OT�B�i�G�-�����L����"OJ`�CƣM��� �x��A	"OT��튣@^����J;	 *�1"O0�X��5$�������mNA�'"O�E��f��{�lp����=(5"O6�B�#'�Y����4{�\���"O�I�p�Z�D��]�%.Ef���KB"Oh�$dڅJaE���r(K�"O���CM<�AS�����i3�"OU
�D��~v�r䮙"d���!�"O�t����B�d\ C���lx�"O�5�e$.�eh�ϟ�x|�	�"OɃ������A��	��"O�T�s�Z8="8�Jc�їX�V$�q"O����\2��Ɂ��+Q���p��-D�xᵮS�!���T���Ń D��҇�X�ʉ�GG=�\��B?D��@�\�?����f�'�x4!�<D���w!��J��fL���3=�C�	]i�-[��K+C(�is*�q|B�I��h2f��9h�J)Zq���k�$C�	 3�ˡŋ�}�j%�U��"O������&/�d��_�4�N��!"O���E�+��ĲT�+��*�"O��A���1j^Zma���4����"O��k�ED0V����Пf�HEx�"O�pv遤B,��~�F��"O����F�D)I��A�+�DL{�"O
;"# D`ҵ�Fd�ŹE"O��#��ʺ>�|�{�b@B�nqx�"O0y�`f��V�,�9B�] u����"O,d�"倂6�>��/G�M�Y�"O�I��S }�����PO�ذ8�"Oސ*��>|m�}�f�Q�4��Q��"O椢�^J@�i�

]�zU��"Oj	3@Q�*]�i
�	�H�|��"O&�8F��l"��C�)?m��0 "O��B56�e�Ite�ܒT"O��9w��W�L��N`�`C�"O8�$��R�
Pm�:B"O��Pm�b�"�����nƄ��"O2��D�*`N�I�����"O6}�EF�	@�W�P���!�"O�åŖ�1��]2$��N'V��T"O ��~���f��b5��"O�Թd	�	����tKњI*���"Oj��q΁%��2 �vF���"O�e�%�Ů�����L��u<��z6"O8�b��H�\Ũ�lS3(M�"O�����>ֽQ��V4[$�8h5"O♪c���B�dh��;Jq[�"O$̘�� #2��x�K������"O81�b		� ��1ZFI9%�643�"Oբ����~m�$o�)����"O�fHͤ-�ФR� !!{: /�!�$�itH��,G�B�k"���k�!��ϤS�+	Ad�J {��8~�B��ȓv����X���!,EV�܄�2�,�p%k�2
�n`j2KJ�x�Ą�S�? �x��j�;A��+Ũ�LK40�7"O`���-�o�v��h@�~B��@3"Oȫ5�ܘjy�@c�՗?=L�"Oh���M� �L�9r)��	+:"O�s��:m�� 	�8�E)�"O*yp0��;�<-ɃBD 6��@�"O>��D�ڻS�^�QcC�qfb�J�"O���̧6F�X� �.�E3�"O�|�Do�7D7���e�[��c4"O�O�%^�%�� ��0%"O�XT�U�,�����-�m�V(ڲ"O>��$�&g`}�E�P�6�ڽ�'"OFE
!@TV��0�M'P�����"O�9t�"r�U���+|��hZ2"Or(�Q��".'�������3"O��S.CWX�ѱ,طD��)Qp"O��0�/�7k�	 �lN������"O�XJQ��%7����H�V~5��"O @�g���F�&�*Y:89 �� "Od袷�L}�(��(��;���"O��J�|��:�B���rv"O����ו@�*��ɋ	�6���"O�8apĞ ���Ke�ƅit�Z "O��a�h�`��ꍨKt�۰"O>|�����n��̋ �|��"O�ݨ��B�9�s*S +Pݲ�"O` ��`��q~5q���!t�l�U"O�EPj��0"�@�ZM��"O0�4E����r�\;aF b"O��%TsE����D�OG���"O.!H���;=A}ذ�� v0�l��"OV��
T'���(�_�:)|��"O���Ē#6\��P!M�)�'"OH�{�/(YL����@�
O��"O&�X4��P�<tiS��A
���4"O��I'��.�4�v�U�p�"O ���`�lk���1��v�[�"O�,����`G�<SuG�> �j�"O2�cv&$-��I�T�tLY"OJ�@Jf�h��r)QZ��,�"O�h�ꖂFtS&�޸�z���"OP���І`���c܆j (��"O�u���n�b��g���B�"O�e�B�մf@(��7����F"O
q�A6�������^RvE��"Or�"tE�6	�+K�:|̺�"O��+a�	d��rC��+%��[�"O9����/��g�Q:IĒ��"OX�`�4Jn���!2�d�Bc"O���0B4i��Y�/�X�b,G"O���ο/���HZ�l��"OnM�B�K#�.ac!G�$Q?^��"OB��$D�@T�W��7��q�"OvYY
=�� 'LܠwB�"V"O2�Jdɕ(����bh��P_r���"O>�1wiڿ#�)���!bLƠ�w"O�As��ë/�}�񨖚%5���"O�Чa/uZ,$��̛{�Fu�"O�E ���9c2�k@"iE�0i�"O2E��H�薕�!hLe����P"O���EL��S�$��C�Ux��x0"O��đ7����5ʒrt"}�"O�����f�vL{�$�=;^��@D"O&|��MY)�(�zQcF�Pt��"O� ��y׎$ �X����1���6"OB��檃6s��� U!N+.;"O��b��� �;�&�-)����"O�]���J�M,���;7�����"O��!�L�m��HVi^�K����"O���e@�c���sH��z��h"O�8�藮l�`�qwf7��Y"O����F�	�b��:pxI�"O� j��"\V�`-Đ*�`%"O,�<,��m��O��*�F��0KH\�<�D��l{6�떒o�NłAN�Y�<�$�S�y�
�8�ń<GB�KvdX�<��$֤C uai�D�YbA��R�<a䣓�W/ڴГh^�xPZ���M�<Q��9,�1L�Q��:�Ur�<��*`.���0�DB,����XH�<����=%�8C�A.y��QA�C�<��jN�oK>�l®6e�� f�A�<qfG�X�T�B���0K��kF�b�<��[<{��B���u�@�4��Y�<�k�9|D�E��x򸨂Bi�^�<���	�6U �Μ�hBpN�\�<Q%H
W���SA挎>1v���B�<q����V���1���>⨨�%&�A�<a� U>X��$�g��,a�IA�<)�T8S�tę`[,�L�(m�D�<	�� �adI�d� Tx�b+@�<�b�¥5�ڌJg��?�~�����z�<�����BC�5r���'%� "��Nu�<YB���c 3�"��[L�s��o�<qկ8O�F� a�R�@��7Ȉo�<AU�H��fA�p@[ _���э�m�<Y!*�uo&a$EN���Xp�0D�#�H]�h���²�f����5�,D�ܒ֧5r��L�dA\�;��p0�C,D��#���aI2�U�!�zX�B�(D�,2��#G�,	2G&Y�R��E��i%D�4�[?�lPi`-a�l��"D������ W��y��존.D��XTƇ�}�H�H�"P$a�4��+,D��B���)�v%��Nn���+#o(D��A�.'��)�`�gK�0c�`9D���;\�~M§��\OB4"�7D�����w���'ZE��)��6D�@*(@l�6���W��%���3D�r�k�U����I��]�J1� +0D��Ki�/1��4^�[1^<"W.,D��(RC��9�*��ƩZk�x�AE<D���DJ/X��L�RpZd�u;D���K8�F�X�lU�\���;D�T#�	,N�9#SN,>,���-D��2�9H���H�� T8x=�0D�Xq^�k&0���&~�D��� D���ʫj�z����BE��?D�4�7�)�(�P�!
�'���i��"D����"����ì�0T��n"D��J�	�v�"�I���~�.��>D������%?-�������� U�`
>D��`�/\�� 9e�	�v�@�U�!D�pp�A¨*�-�J��	3�(��2D���ӡ:! ����DFX�A��2D�0��B"�5��%�g����0D�8���P�����E�\�
Ov���,D�d:���!�<���\kAJ(D�� ��j�m�r���1�"ޮ��e�"O�Y��Ѱu~L�vB�Gl���G"O哧˺nˢ�D�D¾�z�"O���îpZP n����zd"OV�+� ߡRG,pq�l��8�2r"O�h�`�-L. �V�b������v�<�rb	߼=i�f���t���ŗv�<��֣P*�혧�\!<5$ԙ�	U}�<A3�	u2z ���9ɖ�11�B�<��퓞,R��I$Ƃ�v<M9��{�<a��̞^w!�p�#���6�N�<q�L� U� �:�-����8у�J�<)�g��?m>��VC#\��lP�_k�<�hGRa�����5P�]0�h�<�`CT�	 �\��`N�c"��bBc�<I@����	�̛�`����Cg�<	ыB�Q�����@�ܝ�w�XJ�<�C�ɠ �bx�@�c�<k h`�<AgU�n� �22a�Ld �PÂ_�<9Z#�<�1�#N� ᆉZ��f�<�3N�o�2�	�ǐ'.�ȵ��_�<Y�I�?��iG�uV��aV@`�<AbJ+�dl��N�o&�`��EV�<���G	Pl� 1�R�)%p����U�<����� !FӏJ^1��/�H�<qwj ����6#ևD� ��%z�<!!�� s��J��L�R �Y��oIx�<���̮S�ƙ2��<J�t���t�<���A-lx"��θfp��9�*u�<���U"\9�dP�AF~ʀA+Qf�<T"�3n��)�F�v�&PA�N�<��hH;b� ���K�o-�1����u�<���['<�����!m=����W�<���Z�/��|��I�V�eY���x�<�QN	1.@�L0W��	\5MY�c�M�<�3���X����,ݝy��YA��_J�<��Ԓn
,ʳ�(T�0%�p�<!!L15ލ�����	fY�M_o�<�2G4C�pZ�'�$U�(�7�Lh�<Y�ܗ'�����t\y��c�<��(�4"^�s����MP2i�c�<���86ٺ�1�JY<�\U@�u�<Ap��,�L}j��Ț��$DEL�<!G�G/_���F`�LU =d��N�<�A4q�����J+V��� �]d�<iP�l2x�q�C_�$m��͌_�<!�IL�U���f�pa���[�<��P�C*$q#eo�l	4!zE�KO�<����N�Ȫ���*H86@�ǫYO�<�"��,1�a���I=h� ���C�<�#dX4J��Lр��xN��ؠ,�C�<Y$��)���`��m�rL2�iQU�<�BD�(,�X��G�K��YՠBP�<�s�%EǤ}����q=�P���a�<!ԃ�.�v@`�-���i"�\�<	�+ɢ<���Rg��	��Y�OXt�<���N��J���f�q�Ze�<��Ø�UH$��.��A
Yj�<�A���lɔl�d#��9�𘙠�[�<�S��oD��Q�>($����Q�<�t�Гs�hY@��ڔ�l�d�<���������Rh��8�q`Be�<aѭ�� �t5 1m���)uy�<9$@A�J�[lܮ.���Ώs�<�  Y �WN�3 �+H�P�"O�l��ȗ6*s�)��6)�$�"OHP4	��Bj@�]�^
�1"OF�R�Ǆ% �{OӃ:���!"ON�����Q1�`8!�x�+pI���yR��	ͬ��G�Üv���EW�y��0.U��6�	tQZ��D_��yRo�e�V����3`T<���M6�y"���rʣ��)-����e^��yҁعm�XK&)~`hم�T'�y⩎�>��	��6�:����y2i�KX����/�$	���+�b	 �y2�THEr"j��y��Q��C��y2�Կs���C��@{���O���y���	8��1��[@]��qF��yR@S�u,dx(����D�tUy4l�0�y�a�"��@�ԏ����# ��y��P�,<���vb�|�C�:�yrA7$�I�큓醬k�-�y�`�$Y��y���5`���F��y��#~�ʵ�S���!ɔ�	�/�v�<�D��K\���
xt(4��_s�<	����r``eq�"�	k:���̈S�<�2Ec��qm�2"���N>!�DR�Ֆ ��^ �\ʷ�R��!��*�40:�'ڍt���yL�W�!�P�802U���L�)�rXd�ю�!���yƦyHQkH�\�>��i�9�!�ͺ|�F��t	���@��(��C�!�d�-�]��d�'�P�btIĻG�!�D-�|(#�E?l`�b �!��7��R#��?c`�� A�?�!�h�lѻp�ژ&D|}y2OZ��!�dM�d���(�H���T�!��D ��m0Ԯ�(sj�7LI�!���vh^(�2�ɒo��*���
2�!��zk|Mz]>~iX�y�<V�!�_�V�)듪�0� �S��8Mw!��O <���0�f�0�b��=g!�$ǲ7	����Dk颩K��cb"O����HІ.��� ��n�"���"OΤ�OI�����b]�Z�j%��"O��a�I[t�� H��ʾ7�ѐ"O���#� Z��uX��E '
��y"O`��.�1k�)��Ud�$�d"O��92�O�JF�p'$��Z�Hҁ"OT�@�����Qr	I� (P"O�9q&�0*�X���"p_�4[�"O�1茻( :�dXL홢"O��Q�¨&ê塤bڠ
�)��"O�`���8]|U��(��k8�Ez�"O�i�V$��!فGү '�Ibv"O$5@�%�*K�!�'�V%#�` g"ON]�G�].X
�x�̡��c�"O��E_�mg�`A��I��lS�"O�P�"�Vf�cV�U�%��"O|��p�u%�ڐu��9���O�<�paXc�"}���0��\���s�<����2����ꊬO~�Dhx�<�`��/V�8�
�B�,����Y�<A6�͙RԚ q�K<���E�X�<9�hO$������,6��B#�Q�<��'��j�Ss�C'?�,Q�e�@K�<��-�~�2C7C��=Z��9��\�<� |L 5bE��,���EV.u�<��"O"1a�c+,�hSg%ɽ8�9
"O����g��ܡxA��PV8"O@!�P	��V��(SeE!-V@�F"O�)ru�-Q�̽[F$F:�ڑA'"O�ٔ��l��s��?��(yD"O B��s�HM+��[�=��Y1"O�U��h�ua��� +�vD� "O�D�uL�1&(� ��/sXV��6"O��
���;�z�$)�8H����"O�\��o�^�2QE�� �!�"O@�����NάT
��y}r@�s"O�Y��E�	s3T����ח)�ڕ2"Oڥ[��P�|�Uم��.��<"R"O���#c�5�J����H�1X  "Ov�����1*|(p��x��h�"O��BU.DR1���4 ��>� "O~,����5u�xH��)-�,Aj�"OZ,��� ��x�E���`�HQz�"O��S�f�n�(��!ʙ:,��aY�"Od�0g ��g�L��W]�L�C�"O����`B�h�*�����Ye�p�g"O.�i��3c�T4�#( �_K�;�"O�)��HD:~��q���"h3� �C"O4�����]S�x@$#K�n��T"O�yq�u�����4\�l""O�Bf�S8<��Ht��b��L�Q"O,<�6��'$�*�/S)����"Op��6(O)]l�c�6��;F"OX�a�CF�Q��ߊ��(�"ODa�B����T�z�.ˤ;���B"O\��b��4���`�M�^gN̋%"O��;EğR�t(#M�rE\`h�"Ovԩ,P	ciRX�T+юl�6e��"Ot�'�
>�q�E��7@��2u"O`���	Y�v	�$�ώ����"O4�[����:�*���H�#f�^X�"OؑX�#G�W�Q�D�q�z	��"OL�E��d�� Y V�Eִ$��"Otp�EA�  \u٦� %N1�,-$!�D��h��ѹ ��T�
�aϦ3!���z��X�'�Gxht�`��4�!�D�� ���8Z�u\ö�K>%p!��#�h@�D�� _���QaJ�pR!�D,x����ts��	VE�yG!��%v���Ic�%:k�DR��ݻjA!�D�|r����^0}^�(c����!�d��{)x<��
�B��ʁ�P%�!�$�W�@�JV��*˞Ȁ�ĂIf!��߿si01���: ��S2�2uf!�D!g�J�����D���0e!�N#D��u�PA	lc:��'�$(U!�$��n�Q"�&M ͩ�A�!U!��͛�mMh�m>��	S��4[!��()!BC�:t�D&E
xS!򤙥�Е����+l�Ƽ����e�!����x<P'�z�(�l��!���c���lҥf:������!��7y��:@�%  qFc�!m�!�D�f`5�� oR�@P�fo!��	�K�>YPTKJ�2$[��ߛ�!�Ěb�2a'�֛3�d8+��<7u!��u��	U#�\�b���H�;h�!��+!:��S㐚W�j��Bg�%WX!�� j�R�ǘ!�dP2f�h>�S!"O~H��Kվf?F=q�N �
zF��"O�}�Fa�����1N%vJ![�"O��Б
RAh|��,љ�� 0"O�����H����Ʈ�Y]:͂`"O���n� [���sE�ғD�$�3�"O��
�J� `Yf8�� $i�͡2"O�y���]3����&[q�@R�"OV����$?hF�3�Tu�@�w"O����O�p�%��9f�"�"O��8W�.{ʐ�xӪ_�d1d��"Op=[T��!ud0
0��/Dr%�"O�M�#g�i:��Bև��q08`v"O(}�
Q�R����`MҺ~搳�"O������20�&��P��3x���q�"O�ݻ�� 3Mɐz�v *3��!��Q$S]����Z�����4~!�ĉI�7NX=h�&ޏ�!�$�^���qB�����#�%h!򤂺d>"���D/T�rf���[�!��4gB����Xi��f��h2!��A�y��P�B��f��a�1�!�^B0��n��@�a�G�v.!��
�PS�J�W��0 �<`#!�$�Zt����� w�|c&�Y l!�DߜS�H��ܧsZ�ѳ�`A�W!�D�Ws���hʹ@�,P`�P�S�!���l,���,�XE�G�hT!�$U�bhl�E�Z?F�3��oJ!�^�<�qbe&�vtz<B��-!򄁃�H��D�b�(&l�".!�d��[_���D�ßKH�4j�K�&M !��3�4�) �ז;&X� �O
!�$ޙU��C�ل���´��r�!�ā�t��6/��r�p	�%+H�q�!�dT$����$��(q���>\!�]W�}��G�2���	�Z"q>!��C+Z�a�FZ$$��`A��7f+!��=`C� ��B�	�$�W�U�H�!�CiO�Z����-w�I���x!��O�v(X6)Ȝd`��!� |!��V��"aP@O�QJn��SJY18�!�ĝ:U�
��ck�s̼\��H��!�$�E�L�Pt^+"x��afP>i!�$C�|��%a�a7V��ѹ���V!��?�^����	ܼe��ʾU�!�Dí�IKf�Ǆ>8�<�&�8�!��يG!�ћ5E���d�a��T.x}!��O�����ͪY�D���X%?m!�E,bԹ��Bн./zܲ!k�+W?!���w�"!�P���!����K�*�!�W!)�`�1��R$�U���R�'�(���O���{��F�v�L��'�܅J��ӆ[5ґDw((��	�'��K��±kJ>x b��n��}
�'b*�@��x�,�
�틩lL�y 	�'�j[P�I9��r�ꔛ]�ԡ�'�hY���d���8@�¢6.�(	�'�p聢�� u p���V��z�s�'���	���h��@����+Y�u!�'�u�P��#c�Qrj�[��UJ�'j��y�˔�5��bO)YX�| �'���)a�է.e�鐄�w�N1�g"OF�z GŬ�.2�h'>�(i"O� @mҴf-n� E�B�ЄxA"O ��1���_w^ej5�O��u"O����A ��s���#�)1"O�Y� �K����I��D�s"O�)�A�-��P�,@a~~q�7"O64+*26����L3XY�k�"O�T�� �ƽ[�Z�Q�nP{D"O��i�!|�x�oQ�Dd��"O`����6�T����!:1NȲ�"O:�b�a\�!�����,�w����"Of�h�C�1L.��t��"O�x��f̳�8DS�m.,�t��"O�mP�O�"���5l�lr� ��"O��cr�G#Lԛ��܍bI��PP"O�0bG��5w��ĘS�U
z����"O�yt�B)8f�A���Dp��h@"O^uc6\���q��3}��<(3"O���&L��H��6��w��A"O|yQ���'X���%靅��)yC"O���)P��Dh�n��C�"O��ʔ���ur<yR倆=��x��"O��P�b�s��c�PyT� �"O����.$쎭��M��t��@g"O���N�v�Nɡ�c6��A"Oz�!T�����EL��|`p"O�-��wTf�1��S��〘�y�͕�b/�	A���@�����y"��>9���j�09��@���T��y��ĮV�� H�6ߒ�03�ǣ�y��������@�3[��S�Ǆ��y��c&�e�AE_/1ݤ`
�y�����a�c�H. �B�:�+���y� ��cބ5b�CF���yRO��`h����<���G���ybCC��%�fJ��T������y"]�t^U��җQ����yBJ�q *u�VO��F� ���yҌݸ����v�'n.Q3��ك�y���{V!Ehc�q��֞�yR�qr��SS �6f?6����/�y̀?��ѣ��^�hR&�%�y�P<L�k�߽h��!�ř�yR�Ǻ5���igN�7z��r� ��yr��6T��ը�y:�J]!�yB��\t0#��E���bQC�&�y"�6u��0�˚-n����ʸ�y"�Z��ر��X�h�d���I��y�:8�:���/PxX�=c��A �y�W8��� Ŷ����c.ח�yb��x8a���ڂ���*ȉ�y��"^�tQ� V/�dqq`��'�yr㝰&�`�G�9u�By�Fڏ�y���<N9V�r�nكhxqw�1�y(J.\��ist'݀n���J�ޯ�y�6R�dj�N��#cE��y�o��%f8x�JK�6�S���(�y`��QS�$����J IfHЋ�y�gX�kl��	�n�\c���<�y�Bҙ?p�%3 ��l~~(3���y"eגu��jW��6km�9�E��yB�>�b������t[��9�yBDݤ:楩�mA27�2�h���y�ؽ����V 4�4��)����'�ўb>1���9@M퉱�K�Tt�S��;D�� ~aHrb0^W�$�Pg�<ֶ,y`*On��'/�'vQ����W]�|���'�D�91N��4Pxd+�
Q)nl"�}�',.�)�ǋݺ��t��E��A�'5b@;��O��� �cP9�d�'�~e�5M�~�J�:j��D���1���ɪ5��Z�'��T2� ؐO΃/+�7��<�R�-|Or���� +�h�
ϭe4�Rv"Oj��qHW�Ƅ�X�Ɍ#eh���"O~ؚ&+O9����'V1)w�|��I`�O��� AD�V��x��`A�5qf��ȓ ��j�'�v�
u/2r��A�ȓV;�M�k�"�R0	�93�`��'�ў�|�ɂ
��H+���$7�T�1' f�<Q�
�0V�.]�Bw�m9r��G�<�sIY�t��<� �ZX�`5Q!gZJ�<��j�=+E�4u)��� r!Jy��'���r��wBZM㝮e�H��Ó�hO����ń7?�B�)��/W��I�"O�u+ֆ\�`�=��۪G�(	�G"O�E���9JV�ix�g��Bp<Y�"Ox�Ja��	x�&��*J�h��"O�j�iS)3�-q���+!����a�cH<��*�U��!����?g]�Y8C�EX���O��{��..7��9f	_8bk�}BO���Q{(2��W+'%��L��ޘ-��	Vx�@h�큮# n�Z���f<n����6D����^8z#(Y��@��$6B6?I��d#�I���D�$ ���cD%Z�`C�ɴ���k�\�Umd���"S�LC�I�0]�4���@�����o��km4��p?��D�5u���!@��t����w���'u�PY1�E�Vs��@�I���ȁ�'�p$���1q��0!�B��5���1��d�ƈ�����G@�qĺq[���3
y@�|2�)�'�T��ű�>d��mu_���&��$a��S=M�탄/\�Z t,��J���C䉝!Ldև��K�>��󨜸f4\�'�ў@�>�-�l��a"�� �r�n�_�<��I�;"��H�Q�&<m�`�Q�<����F�^�(���'Nr���q�'ў�' 86`a7YrGz�{ŀ���y��N�@�>�
ְ�鷣��2�,���Ζ�����ȓ>7��Q���j�����Y�L�ȓE�������MH�n[_Ά}���<,��hƒG:�p���� v�q��<ڪ�Cf���,���gF�
4ą�"j��"�ÔS�Pta��^�� ��ȓy�x�9"�1((��Ȱ�p��a��oLp(xS _(+����fb
8�u��"}b���f_�� R<"��`�5���O+�	=�0?�3�=o:	BP�5,14��I~�'&�O�X�"���~ND3m_�?~j0Y��'?��3Q$��Č�,KWn�ɢ��7B2vB�	%��HF���U�B}��`� O��p���OD�(N2E�gt����;Oz��w#�2gs��Z�c�o����"O���W.���N��㞄J��S"O����r<X�ٔ�ٵ|�|����A�O7j)#��:x��'׶o*�й�'(04
�=,�&��P�	b�tm��'���aS�k�<���	\;EQ���'.���ո����bfB;P�:���'�6�����Gu@���*��O%������ *��dfƭ'vh�#5E�.��B"O��Q` W	9���W Nʀ�X��	Hx�x��$�q43��&�X�c3e#D�,��QaJ�Te�c,�����hO?����2��i�R��
3��9XqI3va{���y���q�K���p���JN�'�|�o��18���Cže8���2��;�ybbӵ�����N'\��L��o��y���D3�0f��|&�TgH6�y����� �lD��q�J��y�ė|Gt��/�2VU�����Ƙ�yB�¡=�=�P�\+@K��`3"��ybc�R4V�A�ԏ?'v�㉁���'a{OO�My����kM1e�A×���'��	r�O��ذ��η?�JAB���H��=��'�X8r�ӢiH@�H��X�qH�'�4-Q&��)'���
�?�4��'��Ё2�S%[K@���N9���' �%�e�oJ�=�`/�z9�7�Y���)�f<j�#"�rȴ1r�%H�!�$�&��]�rJ�#X��I{���h!��Ft�`����H̽0�`> �!�U>a�Ri���}^2�SeO�s��z��d�������L# 	{���6z�!�d3\�buPԩL-����'Iy��xD{ʟ��cv`��Y|�哠�&���5��$$�S�O��<3 n[5�by��GL\(�'eVLp�a�6!�p��!�#����{��'��]���K�H�
�/(5m���'��B��0{0�`WĂ�^-�M	�y��z�`�DO�*~z
�Ĝ�p=��}�bت#>�XC����{  ����X �y�	��4�.0;a���n#���D�/�����:�)��I"�Pk�G����a�*Jx�Iæ�ϓ��S�OyRhxV��~c���Ӡ�B)��1	�'�Z��J�k	�9@�	Z4��@k�';VśǍ�.��	d'�V}��H�'a��!j0E���W7E��`�d���yB�\
K��~�;KZ��p<Q���l��KŨ�;r5��f�K^a{��Dۦ��aK�28��PFkQ�A	�O��IP��~��3l��M�ҥ�k۶8�С��'�#=���D�E?6�@Z��WZ��`"O|K��,��� ���*Bo~�*�f*�S��y�JW�8g�p�I��F���D7�yB���#� aC��R�rA�B����/�S�O,�|z焐�s�a4�Ѯ2�`l����~��4c(���O M.����2mcqO��=%>�9$�_�g]�����B�`q�:�O��v�(x��ӉK��|X�Ο9�XM���M#�� m��L��>Dp����l~��i��"|Z��H2>���P��W����ħ�i�<�U��)��A��S�>@�ኂh؞,�=��.\�'ylx�2�D�L=�uHA+�f�'�?!����H|J��(jL��"���c�<)�>L�>��DQL�@�@�J8��Fz�O[�F����Ģ'�"H��͘��y��ZC�A��� &���r&)5�M��'�:�w�ݾU�Q[�N�\S`�
�'��<�aI�f��D�s��2A���
�'F����&l�T(���ĨA���(O�$�)ʧo vm��	Vk[��S`�@�wZ2���Dx�UƄ�j�{�I��6Z�чȓЪ��τlм)�"���n)��S�? ���"y�Tiˈ*?yʙ"4"OJ�TF�m`��I�#`�|��"O<�q6��J�X�GJ `O�@0"O�����Q|is�<^���A"O��)�*s���x�ͯV^nXa�"O8�:��Z�e9a �gSޥ��"O�Ճ� /i���ܺ[s�u�v"O��+㩞,9�x���K�pI���5"O� �q��Be�+�?2$عR"Oҝ `e�'*p`H@�_�.���S"O�4��l��Ka���k�/y�N ��"O`E`'O�#L�8�P��ʷ���#"O�-ʤD����Yj���:L�<��"O쑈X�L�>��j[r�@�S"Ozx�e̛���o�-���""O�aJu�3a�nU���9~E��"O���3
��i� ����٣L(¨�d"O<e�DW�B�FEKd�7/<��E"OdQ�J�!��E2Em¸;�0}+�"O0�SfKҦFP*�Tk
���X"Oe˱B�z��aP�	��|P�"ObHQ���?,�Dq�+":Dȗ"O� �� e��;�_7O/��5"O0Ma���&�b<sw)��L(�E	"O�P���ðtEr(:���YF�̨1"O<(!Aʙ!Y@*��dx�)׌М�y"����� 1h��!-�)�y�#@%���c��>X��1(��y���`xD�!�3�[�f�
�y�L<�aX �j8�1�ٜ�y�n���|=�Kߎ[ԣ�,
��y��"J���3�\	���3��
�ybI�]*�� E�MΜ#_hM��'�x%c�)͞�% I���1娚l�<�'a�0߾���������6�H�:�X�� mf!֟24<��Q�(Y��קVh�9���V�\��ȓ��""吇iuIVF�v����'���T�Ct�����	�輆�?�j',��+��t���{?~P��Ϻ�B���u��M�6`�9c�BͅȓU:��ǝ*���b��2>� e�ȓ;҂<�t��I�7�,m�	�ȓQ;$=�t��(�>���aTF�ȓ��0%�χC\��iql$IU����q<�0`�A$��<�rC
�<��u�ȓM���(��?5����C�/V�����6�ԣz��,f��-a>4��9�z��w�C��5馎ܗMl�\�ȓN��up��	�I2&� ��ר�,��ȓ~zx�+X-{X��"�^*Sd	��,������GD ���f���V�<�T�Ņx�`�F�|L�k�B�d�<��nXDo���P��76M�H���k�<��@�0Gt�`�AG��U�u&�a�<9�2|����S@��M
�+��X�<�����;X�
��.>�l����l�<�U(X�!߼͡�IMn4�qE��k�<���Y!.�!�����9��_f�<Y�fÁ4��&��!t�zM�6� b�<�W���@�"i����6��Y���JA�<ه慶iS�0��I0��C�Jd�<y'�ƺ~BpsT(�	�� Cb�z�<)�(T>X{�L�������Gv�<�3��,�*�ۋ֠��$z�<� ��x�IƝcQ�)�.�L��`�#"O��x�#T*0K�yhB�Z(�"O�)�kW�H�,X�E��3��HE"O`h��w#�T��+�1f�Z ��"O2ػ�)("�$ajπ_�ޙ��"O�`a�����IS���t�D�0"O��صM�9/MJ z��I\��y�"O����?��m�TbI�|5��"O�(h��A?D )�a��'����"O=8�!a�]�[�@�p1��5EM!��CP�z�iҦ0{�e���ͦ$!�$J*�@k�΍ W-f�D�D!�D�2%��PA��(|����nׇ;!�$ϵ`�>\�a�%(g���U6r:!�D׊_\�·��6kAb`W�`�!��֙u	n�*�K\Mv8��v.ݨQ�!�$�;�j�+�EߏNB.%�E+Zn�!�$�iT�5�6��8�����v�!�$J����b����i� �Ub��B���<�xA��28
�q�Ua(iH`B�ɕq �Ő��B+w?���aH�;�$B��"|XHM��bX=>��5����2Z�6B�
@�< ���#	���@<B�9d���g��SL>��D+ e�C�ɩoz,d{���DLJ0��ީ4~�C�	?kDX�B�̎S�@��O��~��C�əw�Ɖ2a畜(��t�$�C�LC�	�54�TP!(�/[o��a���.v4C��'y�����&�%*VV�� fܯ
�PB�	??���F\(w $Rcڝ#��B�ɞm�"��*�If>�XR��P�B䉐my��+���H2��v��O7�C��4&Y��%*Q쑚�G�1-^dC�I�h'�� K	" !yp��vZJC�I*e��p�����w˻>TC�IZ��K4#�(7�Vub3g8c�C�ɉ0
��
@��x����J�6m�B�	���j0*Z.d2ة��E|���,ռ$�SW>�^93b�ڂC�!��X��ik��ĔB���5�!�D %6�Ҙ�r�,9�x	U�	�f�!�$BE������,q�la2�r�!���$_��嚕�K��y�W'ί!�]w�\#�E	Gh��2���F�!�Q Y��%����1��	��#@0!��L�i@2�E/Q"^���eM�5!�$ё���a����H�i� ��?y!!������'�̩R���8S�O!�W%bW��iU�F���c�"N_!���n4�)b�͖*C��H���!�DC<�$�b)	�;�b,�p/S�&�!���>r%ik���-txD{���p�<9��ڤ	���n� S��s�<�2MU9e	��;�m��.��h�<Q�"��~v��㷨��I"��2F&YB�<-�|f�W�2G՜�mG�<��Ǟ�zrɠ�A�����b`��u�<����f1����.$Y���#��n�<a�J�@	��m�.z<�����a�<)�Q�:A�	$H'$(�@iSB�t�<�ADƤi:�\�r��j�H�P'l�<��ɘ�]���� ݜ,V�� ���l�<�!F��b�}*%����@�Čk�<!���-+�cS!=� aE�b�<� H\h'�N�[܌5r���G=l]��"O��k��\(N�Рj����aI�H(g"OF����,F�0�Z�C�K����"O�})���/����E�-�&�K�"O�T{�@H)p��9�Ȏ�'����e"OV!܍��98��K�R�
Չs"O4�x�
�������fI3���1"O�pH��"~����W�J.j0�"OJ�J)�r��i�e�;�M��"OJT+�#��]	x������E6$�"O H�@аg��!��0y%���t"Or�A��V��y�VL6��;�"O�x!R�M�T�a�CP�<���	"O�k�ϑ""�1L��� ��"O�|@p��k2d�c�>t6���"O�hksD�%O���w"ѺHQ>48�"O
���G��29<�ppLV�"T2�i�"On`P��D%4%���&G�V��R!"O�@	a�I�	L�� �畷.�����"O��1��H�e�;�k̂v*H��'vr� X%Od��Z�Mʂ3�l
�'� ���!Hb��ȜNX���'Zj\hu��5�l1���G�� ��'����J,4���U`ٍ"9��a�'����߿�`��e/ԥZ�p��'Jz�k���b8�$GӦ�,h�'N�h�ǯ��5A��a���~n%p�'���r*�_�<�;��B�R �
�'z��CcJ��BA��1�>G����'z����T�kFȌb�b���L�"�'��3�A,,�����ܠuP~E�'��x:4�,hɐ��R^�c�B- �'p�b����;t��q'��U��a��'O�!�����a����A��D��'Qp9C�!J�g[�+AmB*?/	�'` -��g=#xFI�Я���`�J�'N-@uB�z�Ҍ��6M��P��'��4����&�4@�A�m��'�H��%*Z?>��-kt�ғDJ���'�1���M0�J��D1�
��'�ޱ�Ӫ%ڞ�ڷ ��.��xB�'���R��A��Q#�-��!���'��Ւ6�ۮ9{&$�f�.$����']��n��W�|13a�	�$�
|��'��A���"P�g�6c����'z���m�1s��!',��+=���
�'+�fo����V A	���N>�F@����$�U(���v�]& �
�Z�.'��~���:-7P��`�ʺ\ö0 t�O(`��1��΍4d�����Zi#���Hj-Є
6s6XG|r��+o�ZlR���D�Oذ(���T�el*R�iX8����'���� ��d��-'zwbxI��&�1�7+�a�W��"~Ұ�<3�d��N�%���Pf%���y�C�~��P��*K���piEl�!*�<���V]� �4�J)f� A��HOLt"':yy�s�?'��98
�~LnIK��K���f-W"�vP�BϬE�DH�"��l�z�(
�C��ASIJ?�f� �j��M4
HDzB  V�2����W;d�i%�~�OUt�0b�(RC�}�5�i�<ɖ�V�:�Thx�eT+#$6q�3�]�ٲG������Ťw@�K���i���"�
0&)�0B���.*��`k�'���`�LREXn���$�<"v�Pu�ȟ<I��D��K�����鉯L��P�%
�:���)Ð)�&��D�#T�e�E�����)5�TT����@�Κ��-��P�N��䐉jz]a�5�: �%�a��0#D�9��9�E��Wx��� ��B��7GNd٦#�5|v[�"OP�`��˃:l�:3��)b��̂�im�dQ @�/Sm2|y5,��X��#nZ�)4�ʗ��9k\ldZ�N�~S�C�I�q�D�$w&�8p+ĻYb�9��'� ��@�ƃ_)��"S]>�<I ,9,�x��	s�:0���kx�4��hժ����ŃD�x@�ԅ�BA�T-�
_T0X��'<��j��O���$)��4q������X���ÀQ%�֓�8�m8\d␰��\��H�$"O�YI G��JҞ�!fE���t�OF]���،0(��N��}�Ǭ�<D�m)�F��F�e��v�<ّ�5�0�[�o�=	cL	��v�	aH��'��}��F�uR|�a��&e�=��'.��3�Y�2Ӗ��J:D%T�*	�'68�k&��/�4M�!F1#�ey	�'�N��$��^0A!,1�����'f�� ����PA�*�7�@�q�'�~�qH�:����6%�v��
�'��q(�cJ)(zTP!b�opּ2	�'��h�[yH�<+�#��,
�-A�#D�T������HӈsV�� � "D�����0J�:��1O!x\T����?D�xK��4`�=svE�=>�N�R�;D�tQj�?+-2�B�H�1N�Ð/:D�����ye���I�	=�&�8D�Ȋ���-�V�� �~�!r��:D�����?�����ΛH���;`�6D��k�$S��	yq�؋K�~@c��:D���1��$B�H*@CV�b�B�d4D������?.�v"�� U�Ҝ�@0D���U%�mC(��!��]�vC��5D�P�Ҭ�6x D��8_�<=!a�3D���W`ĴZ:�8!N�7�M�.D�i���<{ΘD(0JC�"�Ɛ��M1D�$f6+ ����C�*yD��	� D���N
�z^D���(��<j��=D����ა3�$
��B�>qZ"�8D��X-E�oP-@iJ�~4Z�I;D�X�L�j�`h��gB �#�8D�L"���9�bs�\^s��A&b4D�p�(�*Dd��XGmɷY�.�[�(<D�Db�o�$^\`0y�"I���ɀ�y"g\; $���F�&k7.�W���y�HҢK4��䧇)a���2�ݵ�y���:����(�.b��3�I��y��J�ME"]�s�R�Q���WT��y�-"Y��3 É�~j�͝�yEN�vj0)Ԃ��?S��ر"��y�n-@�w�^���a� �ҷ�y�)`���I�x�X��ᅆ�y��
*��$�uH�6fZJěVi!�yBH�'gk�	r'_�޺ye��yB�Q	~����`ǳL��d���y2��$��ᓐ շ[���iTŗ�y�H����i���:X�	�k�y�nD�}?�Ђ��K��H�+���y��تp��ٱ6FJ�N4@�2�φ�y���y#q�V�Q�L	AB�6�y"�K�F?ɀ��֪e�8�s3O��yV�4<�S�ސX�A�ܤ�y"��~��!HԂl:v���E���y�ɓ�=�\X���B�X�j�����)�y"#@��D�*E�Q�BEz���g��y�+ݥieZ�cԇ��:5`�{�n���y��Q*q,��&��?b��F�σ�y
� �����F�$�r0�^Z;�p#"OFl֭(�){3(g^Y��"OPĨ�G���:fD�4	���"O�U
�7a��x���W��5("O�8���|4R����2M�0\hV"O܈{%�:*M��'J�^�Z\�1"OL9	��Ѳw�t�Iթ�5�v@`q"O�l�Dgb-Z�cC.L
T����"O4 5�X���5�̓J$aV"O��� vts#���q>��PR"O��җ'�?J��H���2���"Ov�P�L�]�X���A�M���F"O���#�t:��� MA�^�(�"Oi�� H�U$��ZV��+�:M�b"O�hs�)�;tA���5�9�N�h""O���Fl����˴�&k��Yg"Op��b��ɦ��Q
Q	I��}:�"O�)�GvɌ-c�!���11"O&i�d�;}o��k���
fs����"O�E9��GH�I��`x�K`"O���=!�p�s�E�>����A"O��[��R�U�Z�b�� "O�]+d�ݜ湸� �6[��$"O\��.�b��sl��,0�}H�"O
�d�L�o��8:fK);L�:f"O �ab�3<0���/) B���"O<�𧨒�P�4��'Ė7qL�\#"O@��cd��')B��Qa�?#����"O:y@t��4p�z%��;�S�"O�r��>AL\��&�""�Ph�3"Oʸ�%KW�r��U�r��C6"OZ��гW:
��@�,U� �"O�RDl��3�ဈ@�<�SW"O,�1�İ^�0��m�B��aB�"O\�P��_kБ�jǿ(�<1�"O�5��X��������r(�	"O
0҆�M"zJ��'M�x��"O8�ؓ�W(9Ep9)�;Q�d�0"O��,�	��L@p([�]\Jh��"O���
�8H��LE;]\��'M�E#��X�FW�,h'LR���I�'A�Lp0K�dy���i�%N�Z��' ��D Ly0u����Vg��x�'��1�͚D�2�c�A�\Z���'����.�!	��eH�CT���'N��J�]l�xp���V����'T�А(V�{LJ8�&�KC�(P�'Q��8�):&$��Q�jJ4CC����'AШ�@h]'zB~��R䄤>,���'�q!�V+!����À_�`�0u@�'Wj�aTb_*Q`�Ș��T�_A���'7��".
�} `���M$I����'��ǔ2~�`XH�O�Gp0�q�' (١�,t��e3F�RbX��'�.l���pUnЅ_$H�j���'�Șs֥ĸ���U�ݝN��%*	�'�l���'].{>	�)�6���	�'ƬT���y�I8!&��b��x	�'X�i'�\/i�>��@��t��1�'�@H���X�TmbE��k���
�'�*�R"k��*���t�ۤae��2	�'�B���)�4{�D�@j��hf��'�xQ�l�9��@�7��
�'�%��a�I�I�QW2lX	��� � �rb_��D�Y�p�E+�"O����	���
�A��ۢ"O��f�W�w�y��Z��\0�p"O6�c��
z�$-	��ϯ_���y�"O`$��$L+�0�ee�X��#w"O&Řb�åY�t1$�k#Č��"Od���$��jθ`��Ňp)��"O�P2�J��tE4H����b����"O0�SP�I�~���Q�! �)"O^] �D��{���F�#<�Tڃ"O`L1�j�6H���`. �r-�&"O�����9
$ܘ��YP "Or�NT�&��ԘiP�1�!�䐆<Z���d�)7��:�#�4j�!�ď�Z��m���0 �%�R�ۣH�!�Dޖ3L�JWMOpy[gS�7�!�Ğ�!�>Q�Ȍ6�,h�/��-�!�)pF�b-N'+�q��m 	g!��X!�H�3����g!�ė�8�:5`Ă��!xp��Zm!�^)1�m���$����vLYFX!�DL�! �Q7c1Q�B98f�wD!�DеM��ّ�̻A1��Y̘�;H!�ā*3d��ʇ�o��F]!�dA ip�f�2B<�Q$ �%�!�4��آ�CQ9$�%��E� �!�S�!|vY�0g8�����!�!�$�5@�MȔn�%�<a#��K?w�!�H�`@��E\&=�X2��5]�!�$�Gg�X#Aq$Rxڦb��i!�dF`�����Ù�e KfAL�Q!�D�����D�"<�� -P�)\!���s=I����*^a�!m��s�!��FR�!���p4yX�n�4w!�$R�A�r��`��!���6�Fi!�זD��+�jےC�f����$}r!򄄀^�b��7g]W'�2�F�i!�Đ�����S�B�*ÓC{9�|��E~�x��ɢ
t����OAWl�]�ȓ%h��W�ɠR��G�؅�M+�݉��ɮ!�<طۍ
����ȓV����hL��!�x��ȓ ��s�U�vuT�9�T�X�xنȓ~�J1A3��3\�������;m��0�ȓJ�D�&˓�i�H��s��6:~zY��'���x���F������
D�d��ȓq��U�_MnT�6Μ�_�ڽ�ȓ,���[��^:sd�{RޱF�|��ȓp�k��V�A#��k����4��c0��� �T�N�q��n[i��P�ȓz���*2�U��D��$cn�d��ȓZ�|��7��#-���� �j(��ȓ���a�4?
�X��2\@�ȓꍡA�C5����`EK�Ꙇ�q�D�cg��F��EV��0��}(�M[Ao��>@��sgW�d����O�@�M�x!<�Y����$�zɆ�f¦m9���?�P�9�����ȓ~}�Y��O>xD1�Dn)Z�цȓh����F웲Q9�e��o)D����aM�U�T\s6QT�0uӤ�+D����.�	
����Q<m��ŀ4E)D�PaĬ4Y�5�c
O	)j�x��!%D�(+�:J�.M{�d̚GK�K�""D�� ���Ԍ�P���@�X?4,�1"O0|���I�n�^��+�
^�� 2T"O|I�gA�/I󴙪�
LM���"O���Qa���|@PSIH��ڑ��"O(E9����1f��J�"O�|3&�ɳK��mJ��FQ�t"O�e��!��	��t�#�L�	�����"O���p����1ʒc�04*��hW"Oؘ�r��>G����CI4_���1P"O��n�~��!"�L�L�"O m���0SG���\I����l�!��[	J����Q�>�Q�E܄�!�dTDD� 0���s� ��ń�V�!��e�^��w� =���K��Jg�!� !t�`���ʢ\��m;u�Y]!�$� k����5'�?S��9P �@�;!�����7g��0�G5ZD!���,w�-1U�܄n`�-S��Z<%D!�d�h�@���K>\�8��` !�d�4	5\�v	[9���X�A*g&!��{/���vǆ6��L�&gc�!�DP����R�3���� ��/4v!�6o6^�[�䌨1R���D̑i�!�d� ���*M�\F��Z�a�"`!�䊥0J�@f�ܬ7kp�0�mi!�F�\�Q�EDڲAZ��j�`b!��Q�ea���Q_�+�"�9~!��1X�]�FM�Y�f��,T!�D��y�����aT5ol���	4!�d��K�8k�m����"�!�$Ҿl=���+��~L,{����R�!�B�<)�*���Y���ؕ�ݍ�!�d�#)'~�Mϝ���!i]-lO!�ĕ�}�b�����@k��3	��!��/H��5d֛KS����&^�!�DX2|����+st�񠥒'P�!�$KAF(X-/i¤KдĨ��'��p��H@&p��9"���4�5��']VD���*!����$jA��t5��'�l����	�)����`Ұ�,Hc	�'U.�Y1f]X��q �	=iq	�'�Z�"�jB�@O���$/
&S��J�'��]	5$ɸ���H�&�Ҏ����,�ޙ�@G�*;�I�[�:]�⬂)C4����I9"�8��'�y�(L�"d�ͦ5!W����M#g��ק�)#�$�E�%%Ɓ-zt�9&� �䓎hOq�N�!ҦW�8_�tk�ϑ�)!����]�xE{��	Ȕ(6���e�:$#��^V���M����DH0GD��P�Z��D~9�E��"Ota��B;ju2�t�T<n"6R7"Op�� !	-*� �%_�B@�$4ʓ��)��XX�d����H��-3�0�a���>/O��O�>��c�)d\��f#O5x����AN`��J��D:�h6&�*�)���!��4U�vCB(�剛Fj�<XD�O��Y�e��y2�r�C1(�ޤ!��<qw$��Ģ s�j$�K�<�pvʞ)(�Ha�DB�B�0+���T|��b2�P#��]	��$�Ĕ~2���2���$��|��I��E����)C
�	@8���kZ���Od\�1@�O �a��K��f��P敝�� ��L�<��"����Ba�-3U
��	Vc#�H˥O؈,�ܖ'@���2�~�S�3z������z�b��V�,��c����I�8h�`��=�>|S����Ob�c�xGy��)ȇY}HH�֧�	j5-&h���O��=E�tB�P�� ����4�^���L��y��H
I;4���7+,
�(���?�'���� V�\$rkT	Ĺ;2V�z�b�)�� 䀊�G��5������<D��YK�|��)�(��I��R�x��f��4m����hO��lX6��{�]�A"T��Q��8mҸdl�;+>��Iܴs�~��2n;�)U��O��t���_^�NL���XjLH�'����F�>8����
N 7����'���
协�*C\��c��#�x"�'�p\q$��N'Đ���Fܻ�'hn�Y�ӹ`�k7c�$��|��'�ͩ�,S�v�)ˆ$�/o�m��'�`�Q�	��82`��M>cRX���'�ȕ����&Ĳ���&.�x��'���9B�^�Zh"��A�0%���
�'"�ئ+��P�[Q)��}m�1��'2��q�Bx`��h ��K]�q`
�'�N����D	^�Q�օ  J��	�'{T�	e(U !8Ii��o�Rlp�'⎱!�Ҫ� T8V,3}�(;	�'-4К��2t �A�ՙq"��	�'���kC!�"V�0 W U�q1<U3	�'6y"5�׮k�1w��2|ƪ2
�'.���c�A���=6�w��{	�'�n<
���5,$`��d�>y61[
�'�U�iM�m�����	r��<
�'�U�τ��|�i�%�f�&-�	�'?�p�Q��F���4	�='���
�'_^5������l��S�
�.rV	�
�'���آ��= �����Q���'�,��#%Ę8��Y!0��Ѕ 
�'�N-8wn�2�p�9׮�H��x
�'~ֵ��ɖ�G�� s��.v%��9
�'^��0���@W��+Dłr��"
�'��q�5mRO��3Cd �h��P�'��2%_�źB��'Y{,Y�'�,�u�\�-ެ�j�%N�V��'��tR�4S��b��>�LD��'$�rc�Q�.��1�L�6i2 0
�'�"l+� �!���{P�Ue���
�':�Qx�V<,6]��G,'�fp�'�8k���	F��hVL@� ��S�'5m���^"-�@2��Q#�Ṿ�'I�T�f�
[O�p�MQ)�x��'��`*�F�%�f��4���|b����'�Dp��b�z�����60*�'�	�c�#s�v=2�C����'�����ݥ{'r5H`)y�ݠ�'�"4�B�bP����Qk�F0j�'�]YY�ĝK��
XI�iar'3D�8����:+HX�vg����V�<D���6G7l�"�_�M
.m�'�<D�pED�r`!�,�" ���փ:D�D�0��$\�\�j���,�j�9��7D��d�=Y!�-2׉ѳ��s�)D���u�	���Ĳ"��<D�Bi*��"D�ĸ���	����-��+�R�sR�"D��S��:4�B@��/Tm�� D� �Γ	rJb�"a�,�挚��>D�\7�
zr$@�3`@9zv�c��'D�����N= )�qjX�]r� H�9D��:�W;f�����Ip�p�D6D�Lr�&(̢}�҂G
�ʵ���4D��`/��;�L	4�P���}�ec'D����m�'��]�`O�����'D�XP��\�@g=H�@�:�:`�VC'D��`Gg]<KCTC���C�2l{�$D�� �e��l\/3ꢁ���M�
�J�"O�<���6'��%�KoZ�Mcw"O����\fe|M:6��b���"O�)��d��ue�x�Eb�5��U"O�|�"I�G�Ԍ�tb�&=��`�D"Oh�
`��*d=�t�@ֶ1��]y�"O��	��:6D��!؝Ju�y��"O恑w ��* ��ٟl_d�"O�$�gE�iY�)�!��1�~q��"OҨ�"^�'�$�d���-�,��"O���.]4�r���-ڌ�\|0a"O�D�u�ͲA��)��-�$�#�"O��Bbo��	y�JCH���ѳ�"Oj����\W���d�2; ��"O��1w�'F�$��蜒"O�Š�KN�.48��0#��c6"O�a2�	�e�\�I��V E��[P"OT�('�ɝNm� 80gF�8ݪ�ӑ"O��	#	D���Qh��2��a�A"O���-\�pF����'�6�"O6��7���e����
��a"OH�Q�
)��X7)[3�ԩ;�"ONqb
0w����n��u���C@"O�1	��/�ĭX�/�(�^�X"O�-� �^;,kV��įZ3L�zA� "O�� r-�$� p.У.y�e�g"O���#oL}���i׮T0Zvj�Ñ"O��#ǡ%�݀ ��e���"O���a�X�!�#�SjW���"O$iBӆ�-=����E��F#��`"OR�KO�g3x���A�@�q!!"Ov���3U��A� �9`mB��"OZ̛����-��	�A)!34Pq�"O6�Ѐ�4�R��f F�\RV��"O�E����Dd����[�v.�Ӧ"Or��EFlC�-�����zr�B�"O��AD�Q�k��h�#�	}nD@�"O���̪��u�"!˽KZJ�"O��
��	J�D-^�F��"O���a��
��Q�l��_?̐�"O��kem�Scj�;�ː�zZS"O
|{򣑛'���g�°��U�t"O�+ ��f=�� !�g�l��r"O�L���f��`Q`Z�7��0Q"O,�Q!�?�U�rD�ir���"ON�k��.B��� �S�xg<tȢ"O�h@�bW2��M߷H^8:q"O�M�bŮH�b�c�!\�4�Zm�#"Oz�;$ĕi!0#�1w�a�G"O�	��j�v�Q�"ț��L�D"O�4�B��oj�	%���,d��"O�cJ�.$y��~^�xz�"O�$��� 	Nfj؃�@�:��3�"O�u��]� �����1:�a��"O6���FiQ��1��f�̤�u"O.�*�ڪM�T�6��=���8�"O>U��(�0�>|�%�*w�� "O̹H��A?_F���O-l�x�"O~�b��=	����.'�P���"O&���Ɨ?.�z�& �O�PՊ�"O�Ī�C�k���Ё�R �"O��-u����� Hrr�6IĄ�yr \p;����5`�C���yB��"gj��a�$.Hz���^��y
� �!��ɍ�;�@H�d��bmfe&"O:��CB;w��)��I�8J��Rs"O$��A&B�f��y�o�8у�"O���1B�+4"�pm'3v�I#�"O��Ѷ��L�̥0V�/v8�Mڗ"O��8cAPbqJ�w34�""O��WO's4AZG*=w(�\;p"O�d��fÅ'�����Q
Pw:�)�"Of� ��Y|~��4gS�&`�9��"O�(�Ҩ`I#*J<0�BT���B��y��Ǭ |��Ƣ�1-}>�)C�.�y�L��[���a0$�S�a��γ�yR��>M�:���6R���y���3�y���;QJ��)@焉M���M�9�yb��S�z��`a��F������y�AVkEt}��I�<!9S$�y���2�^A@s�^3��iZb���yR`O�p�h˰G�|��1�*W��y��XUQ��O	
���R6�]�y��E
Q�$�0�!K�~�$ E��3�y��<~u:A�2��5y���:"	?�y��Ɗ,��a+i��Iΐ�4IL��y��N8[8|�sgA=	�^�P�D�,�y�i�C#6�����-|\4rC�,�ybh�y_��2c떄b�0Jf���y��)?��a�DޮTOF�bei��yR��2��x�f"O��	r��V�yB�	_�	1Í�H��K�"���yblJ>:Hˆ�K�?�A�D��yr�B�2�0��ȁ@�l�v����y��?�x���$C�o���%��y�o�,!�Z�!�L<:�"����"�y"�4?��d�򬎾H�u"��]��y���>Z���ҧ kZ�T�	U��y�?	�t���Q0fnpU��*�y�CK�3���b*B�[Ь�y�ח�y��ݺ9��I�_h�bEg�&��p��'�t��ai��_dɣT�X��A�'�e��ɘ+U�جq�o�xU�}��'B�͒3�,b~�I�*�g�h��'�RQ��F�,�>�#&�K�d����'�@l�V6�BY�����U��	P�'�0���1HK~�`��_Q����'R�K�D�%j{�`j���$F02h��'9�^+H���@�Q9>��b�'-��L�<L�e:p&ϧJ����'��$� �߮D�b@�W�
�P�<݋�'�T�ѭB���+'�
�V�z���'[����	��"�x���G�D��ȓF�Y�� <
ڵc�$O�
��h�ȓQY���������$V�"U�؆�pnr�صf��H�i���T�B��ȓ6��Q����y�8��Z
-�,=�ȓ����ȟu�r�c"��2�����m\:Q�Ā�/]��CRD�_�����u�	Q�#� %F��d�Ӧ;g&1�ȓo{��A �A8.�2���;S�0��ȓV4�5�(�&crM��(��A��X��R�t� A�)#
V�X��."4@I�ȓ{ I���V�&��R��A`.u�ȓ�I7�V�5fpP`�,ˀQ��ՇȓH=V)�C	x�v��aEϱM8�p��G t�8rk��"W& �6��,D�l4�ȓ)�>�"�mZ�p���'i����S�? �@�FdGYqa��H1�9� "O`[��E�+��ɣ7���:oD�s3"O�)I��|Ip��!��~^ !�"O\P����9=��\�� 2/S\Uq""O*a	�'�S�
����^��"O���7�
�}-��Zvd]�cg��"O�pkŌ;�~��ը�y p�"O��A��������6�2�B"O23� 
  ��     �  ]     <,  �8  �C  �O  [  f  �o  qy  ��  *�  9�  ��  *�  ��  ��  C�  ��  ��  �  P�  ��  ��  �  ��  �  Q�  ��  � � � � A) �7 @ �M �\ &d ij �p �u  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�aʵ)�Y�!��-'���ɤ� ���r����=�B�	�b-��I4�كH�@�
BlC���B�I27�p)�$��<6>0@G-��f�C������+�1�bD�`������0�d�os�\�� Ŷ��H0e�QD!�0x�*f+�0j��ۗHӭ|��F��F�6�\"��E4F�!4@��yrHJ�R"d)���Ƨf[vD��+��͘'��{ү�=@�,
�KZ($D0�.� �y�bŋB'�U�g�O���Pm����:�Or���h]&E�8$��Cj�n���'��ɯ|�&�ɥ!R�>NH\iFW6<�"B��	�Y*�H�(c<�!���4d���=�
�'W	*�S��/9����D��`�ȓa��i�F�0�81{@a~�L�'�#=E��/�A����$ͤ_'BY�"�W$�y�㐚H̔5�V��'�RUJ�
��'qح�§<����Ǣ
z��JTJյH� 9�l�$'!򄇔O��H��ڥ64JQi���k�x؅�G�n�+�����A�A�����S�? ��wN.P\�Q�b��;(M��"OB��'�->0u�3hT����"O�$���n�б��'�l��l�T/�zH<��Q�h/�iQ��[{z� ��x�L�az�f�\�[ФN,�2��m��y��
p Qs��`���	,�y�/��D�f�K�VJj�3*.�hO8��酔3���B���pa�dK�#�!�Q�zY����W(`���qG_��!��v��+'��h�e�?!���,j���J�z��-"��� ,��O��P�HL�����E�.V7\Ջs�%D�`ѐ�	�fRA���ː
�l���(!D��6MG!7"�FI�:���#� D��x�*f���+ *�%:d��{R�9D�`����'�<I��	�,}�\3e(6D���WmJ(=w��q�ɓ�l-\� wA!�O���<.�.P�kћ>�h��Ȑ�vX���p?qCj>\�L-���Z�dS`h���w�'@���O��(qA��S\���+�@�6,��"O<�cK�i���Y��*�q[�p�ObҧH���)'I�p�鲢�����;%"OMa�%���h��n��J��q0�Iv���i� oi�;�i�Ҳ�8�'�5X�!����\1 �b^: ����B'ϕ/ԛ��)�禑�f	an�
S,V	B+Ƭ�A+D��K�	vܺ�*A#�>eЮ���i��u"������O��Xq��3�ҝ8��<+a��2r"OF����6D��ͺU�@D�R"7O��=E�$�.]�PŊ��"� 1R"���yr(�/"��K�B4����abW#N�*X��m��L���ı0���9ҧ��'�^��N0|OrbK<yqԀ\H���c�)]-V�Ҁa�<��
6q��	0#�"��I�� ^�'oў�':�\`�`{a��Q�SF�H�q�^Y�<y�+DhnLsp���|�J��@�T�<y�䕏y�4i�2�k_��j�B�<��'�qO?��J��n�1CnC�a-�֨1D�K�k���`�t�	vK�d��+�Hy�/�П���	<��A��*)�LQa�	�~������<�VnF�]6�!�ճF����	U�<�Vi�=]��,)��2�^�@7oHT�<�2bM%2/���3����v�(v"VP�<�VǑ�x̘���(T}�C�NP?A���'����$�#N�M����t:<B�ɂL� �p ��� V���K�nb���=��ƴ,��P�k9�VL�'�%[/!�ĂK������	� �f��c��@�'��|���р��ʩ���0cM��d&�S�O�:��HӠr��-R�nL!p���{��D.O:<�s�@Zej!t�`�Ne�4�'�B#=E�t�N��2� _���@�� ǨE	rO�80�Pf��A����&Z�PAV��$E~����}�+���Be�H&�a�!�$��3\",0a\�E�)V�N�Oh�=%>��bȽUq�
v�H9isҩ1�E;}2�)�S�t�����8\P�%���!�c���뉗&�X`�S��g�<������p���k�X-�&��{�t`��G9G�^C�Vq�I����&y�g	�aa\5O������m��A�dHɮ$�Q;��'�ў�xf��B�PaȒj��l;�[!�,D�T�J4 �&aA���fp���h*D�(�`Ē�C���e�/l�R��+�t�z��� f�0�Eņ)%�PK�'�\Z�l�"O9@f��zh����H>0wv�����?q &޴);��RP�SM4��9B�ʾM�!򄈭@�z� � �	�©yg��x�!�D۷O�D$��
ےk�R\ �_�-!�d
)jj�p�ĕC���[q�9:�!��g'�\ȇ�U�E�64�f�F�/�!��>6ƨX�R
NBZ��BL!�"K���u�C�Z�,����M\!�dI/Y��R��	DI0�N:DRazn>�� 03QdC8s����	5D[�B�I�8EL����Bg����H�L�N�O�\1���	�X4�w,�1C�tz�B\�S�!����<#�3@h�`�LW��!��Eخ4Q�/
�NOh�ŊM-=�!�$4�^� ��A�>���4h!�D=*�x�X&Eܟ&�䈊�
�zK�LF{ʟ�ǋ`�� G,G�~a�YӢ"O���`�R�ecV��X8��i�,ϟ��?E���
�5��gA�${����ƛ�W���ȓF�^xȇI��}r��q"�I�<
ʈ�O �����تr�N:bj�+vh� v�2C䉕+7"�ӄ�$�ʘ���ܰg+0C��K{�s,����@at��*n�B�I�
]��
PI�;}��(��Y�zB�	6n|P
 �G�����ʑ�{�jB�	�,�α��ń�|
��҃(�372!�䙨l���ggĭCdY Hw/!�DD6[��3C�P�Lz���I�!�_�|]�5��'�w�9"'����!�Ɏ5< �nZ4R�c�Y'Z�!�DM�Jf �E-�{�T�3U�U{E!��-b:*��AMP"W�B �R�q1!��4D�"���L�P���*!��S�m;́9�%5X�.Ja�	J%!��Q"]l��4k�7�2�9#E�!�dE=0���7LY?5/��C!d��7�!򤛂[ˆq)����|!p�^�!�$��m�l*ČQ�a�ZU!�"l!�D&��0HP��3eφ��1���v#!�dE�}��Q��P�x���04��X�!��$Av��V�&z�>!����q�!��EC���Cg�kŖH0�I�z�!���X�D[�,K��C٨4%�C��$N픙�b�ާ~�&�`5���L�C�ɚo����� ;n`�)�Z;[��C�	�z�N�[�=f�X�J�O�C�	//�$�s5e��m���աU) ��C�i���HF�`4xY��_�C�	 z¢i���A���q�G�JҊC�I�`�x��цÇ�;Ä�R�!�˨id ��D'��FaЈX�!�$O��Q�ߪ
��S�#�!�DS+���#��-���B! ̓#�!�����0��=j�~�����`�!�D�n�8��殄9;�(�㪀3y�!�$�C��*BI���p��	R�/!�0Z��աp�`��,j��L�Y�!�߷%�@�@�ܨi���g�T�!���/��x��F�4_���:^�!� v�h⭁YR4J�&ߺ)e!��O%6�Xi����3;��8&E�V!�A;wt��`iP�}
4ĺ�[�m�!�E�j���[<2���qeOS�!�� n����3O���M�W =��"O�ر�
�����g+GjO� �"O���'�r,ikF��?�P@�"O�d��q� e+��Rx�}+�"O�L�dj��]��q[�Ĳ��'�B�'�2�'�r�'1��'D"�'�
��sDܪ�bT��[�.�rM@�'r��'a��'e��'���'h��']�Dkw'�Rc��(\7x6�����'2B�';��'��'R��'���'|赣$��57t��Ӵ.ߟx��b��'��'���'���'g�'�2�'t�[���%fa1*�+

���'l��'���'�R�'82�'j��'obi)�"c�EYЊ��D���' ��'���'�B�'�r�'~b�'I�]���Ԣ
���Cdߌ8�*m�E�'2�'��'XR�'[R�'���'q�����ի�`�g"�-U�|���'��';�'���'���'m�'�l��1��*;>()���?��$0�'0��'�b�'2�'�B�'Br�'��q*T�F> �@���?1���1��'Z��'��'���'6��'�B�'Tr!z�EI� ^R�R�N�R��t�'`2�'�r�' R�'h��'X��'n")i���/C,�l�*1e���J�O����Oh���O����O��$�O��O���eՀQ����cV? �l�`�O����O����OX�D�O�����!����T�2퉥f����r�� �� w ض���O��S�g~�s��X�*I%N�����U�d���ӋV�U��ɴ�MC���yBfӶ\��?N ؙ ΂����rh�Ŧ��	�a�an�r~r�x�d��X��
�?,U�fY�j�L�[F�]�RW1ON��<�����q�l�2v&�$�2�!�!�)��o��QF�b��b��y��F�;��L�GdD�1m$PN�;Hj6m�ѦE͓���IVlW�6-f��h���/�\����{��\:Gl�4�2*�+4C���'��e���T�'y�L�l�3x�и��G�2,�pL�'��^�I4�M��Ɲ^̓��������.�#-P=7(���2��>�Źi�x7Mm�0�'���d"@i �2񢅣P"��(�O� 2��
�k�h�)#󩅧n�dם�?q�#'��� c�v���Z�k]���$�<Q�S��y�)8+�DK�"ȞM������
�y�c�6ٗ��� ߴ���� ��	���"�)x|�t�p�I�y��k�ımZڟ R"�L�Q�'C������,,����5�0	�O��k�H�� a2��'��i>��	����֟�	�(�����HI|���ˍ�$�i�'d�7��gj���Ov��.�)�O�%�K�[��0!�%AT���{}�kb���nڙ�?aO|B�'���˪p�8B���u�"�ra	p��4h &[2�~�)� K�^��C�ܺK��>A��<)0M!�0��RN�K�	�E���?a���?y��?ͧ����y�v���T�DG�-�ʌ9���
šu�՟P�۴��'���Z5��uӦtoڨ`0��p!Q#@Y
ъ��*v�)!�Ԧ9��?��N֩�N|2��M���$��@	��G�^��dH65��aJ�g a�^D̓�?����?����?i���O@`��ReY��2 ��/�0�XH�7�'S�'�47�Q"��)�O��ly�I?<�̌�f��yJ�=K2iݾ�������I�%X��|��W�1��'��D��/>DhP��E�r�\#�h�kZ�(���U�aM�'X�	ӟ�I��I�t�F`�?+�h{r��&Ā���̟P�'Q6m:K'b�d�O��d����
�Sʈ�@ϐ�n�0� ��>����ĦY�ܴ1�r���4���cΛ¢�L�"G�\�B6C5V�XI�bN�s�053.O��	\�2�]���1���(�G���<�RAh� ���?���?��S�'��$��mA�l�
�8��VdT���-Q�B�̟��	��M{����;��0�M{ף���5X`gN����r�̔|!���c����i����럘���E�1Afi�5GFyb.Ó�� � ��.�RXh�`�3�y�_���Iϟ����|����OT��# I0:����dΞ�c��b�Ж	8��x�S@���'��6=��� 򥙓k}��#��K�C��5x۴u�rV���?9�S/ ��m��<A�+N�T�f���iҩ�� �ˀ�<)�m�)���x�O��䓩��O��	�� �h�#M�@���P�"���O`�D�O�˓Jv���Ir�'�BA�?���@�x�4��kݰN/�O�5�'��7�Xæ��������-�hD�$N��`�T5@�����D�On	���/*&�Ȣ��<��'#��p�\w�(���Uw�IS ��(���@�ʔ6�.���Op��O��$,ڧ�?��� �����-��ʂm�,�?�иi���R��'X2�j�4��4�4�e��]�:$͉$��97j�Ly�0OP�l�%�M�G�i-:$bði�D�O��`ǚ�r�}���
_�*�Ɲ�5��إ�ſ~Q�O�˓�?����?i��?�P�T �*�Ѹ�;����-�:��$����֬�����	埤$?���@��%K "��P֚�3T�5��0�OD�nZ��M��'��O����O��x"W䂭Dc��ҤgE�]�� ����_���p�R�̰��HI<p�;gb�'S�Ir�)0t�ԉ~FdA�L�6�dx�I۟���ٟ��i>��'}�6Mv6��$� ���f_�<��h{fGY�Z4��d����?1"\�<��4�gt���r��-r#��!�Xgτӳa�Y�h�"G6O��$1!9h·�23#
˓���� �,���]z�8Dh�D��}�1O��d�O�D�O`��O��?U�₌�A@�N���=�Ģ��4�Iӟ�S۴��$�'�?��i��'�b�j �y���+钦$"���O�O��h���nӦ�)�03��6Mx���A/2P���Z�Đ��Ӭ`4� juC��jn�u�!�"�$�<���?)���?Ӯ�&��Erci�Fc �_���	ϟܔ'�6J�E�~���O ���|� #�9
�b�)��O81�\H`!��h~�-�>aG�i�H6m�('>���+/�N<��N�v�.��#��@�|��o�(��,[_P]�'��D`H����Q�Ɏ Ԥh���=N+��M���'�'R�OF�I�M;��Һ0`,!���I�M1�Y�������?��i��O$�'�D7�L6@lH�d��%^�ʥ4�b+�o���M+��M>�M#�'�� �3N"2!g割V&tDX%G<X�h}ോG�L���Dy��'/��'!"�',�T>1��5&�b��P���Δx�,%n�9&�j�	�����c��u��w^�Ax��K4B�N�y���������z� m3�?1�O������	IV���3O�p@'��lm��I�m o� `6O�Q
��֓O[�x�r!5��<A���?	3&I�VE,1#CN�VpD�3��?����?)����æ�(G�������Ο�����u��mB�O
^�����o��b����M��iC|���>��`�nC"<rn�����N��<���.�9��!Z�	��QA)O��Iւq�*���?��̓0��"AN�&J���� �|���O��d�Ov���OD�D�-Y��Sן�x�Jȿe�����I��[U$�ϟ�ܴu������?y��i���|�wFxqSg�2i�5 �U*Z��1��'1&7M��Mh�4}e≓ҋ[�<���?����"�G* �^)�!G�2c��T�biB�@��[�ʉ������O��d�OX�$�O�J=R��ݡ�E#E� ����N�� Ǜ�W4?-2�'�b����(��}Q��B+�v���_�5�� �'T�6mO̦�����'����<��l��l��r��`�*)�L�� �F5�B�p+O���D��1�(4A�$��<���e�:��¦^ �ީ��'�-�?����?i���?�'����%��jV��z�ŗ7z~��2�(��,�. (C��޴��'���K{��h�|�nZ	L�~QB�� vȺtd�6�.�W'��4��{ 2�jWku4�PK~:�����)#�I�}��!��r��1O��d�Ov���Or��O��?�Q��ڮ��u��耈L����0G۟��I���޴x�'�?'�i8�'J8�	�#9�F�s�Z-:1�����Of����u�����9�2�:O����[@��Hsk@4@��mT�Z[` ��~�(�C ��䓉��O(�$�OH��W�إ�	�q#���@��H���r��'rW��b�47��I���?�����J� ȐQ;�-Nm�8�g�'|o�	.��d�]��4g���T�O_f=�2CD�
�Ę����!8���d֍8~eI�)1���?M�����1��%����5~hJ����8i[�C�`̟h�I�d�I�b>]�'47�� LX��텇) Y�����R�*a�B��O\�$�Y�	e�	#���
��zc�[�n�� 
�~#vX�Vnՙ�McQ�i2��S�i|��OD��T�U{� 
�ó<i@��4�l��j� @"2��$�<)���?����?���?�/�~�9%�~����&̘�ZfH1#�Tͦ�K���������&?	���M�;61&hap��%?x*�Z���GcV�aѲiL�6�ޟ�ԧ�O� 4�H̪�y78� ����+Ĳ��G�B�y�	��K��鉦�	z��'��	����0Q� �T�G)r/>�kV�& �@�I�?����	��<�'���ݓr92����p���)�N���?]f:���I�?8�0�?!�U��
�4^��F�O��*IzPYƌ͛7����n�|e�P��?��P���vbDL#*OR�	F06Hԑ�2��O�*S!J�W	D-�E	��g�\��g�O���O��$�Oh�}��2#�b���:s�N����J�_�H��i@�f/��3���'
6�:�i�yj�)@B��x��""4�`�*~��3�4n-��h���d��MF���O�рK] ~v�M�`�oJ�%	 )ǰ�[�(o鄒O�ʓ�?���?i���?���b1��լ0k��r��&�Ji*O��l��o8Q�'="����'G`�!L�`|Va�W�\ F�x��>ᕸi�7����$>9�S�?́����|s���o���E	D�j8"�c�eyV4�L=���Vx'���'�r$��ȕq#�<�e�P,�
UQ��'��'G�����[�ta޴-�H�z��L���_���´� �JTXZ��z��'��'p��l�6Dm�plھ4\L(�r�ї)FF������E��pȲ��,��	ӟ�[$��"
B�8Q��Ey��O���Vx\ŉD�э��ar�F�D��	ܟ\�Iϟt�Iٟ@��[�'t����	œqY̓@��D�T�Y��?y�� /�,���t�'��6M!��^?R���z3�U-K�F�,��&w����o}2n{��m��?-��
ߦ�Γ�?�֏�#p��UHU�5��C7�A,�p�X�Ο�W� �M>Q*Ol�D�O���OJ=�1��
���Kc;Ƽ9g��O���<�[dL0{F�\��x��ݟ��O�t� �U�g5J�2�,�#� �)�O��'v86�ɦqY���'�j1)�6n���b�Z��@g
��"�#�Y*vm+O.���y�h��&��!l$�l0t�9:�)��X�����?Q��?!�Ş��$�ɦ�a���mR���
�qKȥ@��H�V�$x�����+޴��'�����6(+�6�Q�iP-Q1��Ã��C�7��y�� ӈ-�~�y�����j\�'$���)O� .���]����R�A�>���{�0O���?����?���?����L&���oɯeJ�rQ�%H��Ho��Co�%��韐���?��O�Rv���1B�$ 'lͧ4aaQD��"M�@l���Mk��'[�i>���?-@6��E�Z牦%�"tC�'t��kuM ��I<dŊt#b
�iU$�%�x�'t��'��a&H%\��kR�Z�C	��sC�'�B�'��U��J�4j��-���?A�'�N�#aDԞX�0��
 �<^&ݱ�B �>!�i�<7����'H�@��/�Ġ2!I�0x�F5�'��L4� !����2
��?�r#�S˺+��'��ՙ���?�.��a	@=)���'���'r��S�X�%X+H1��Bf���H9������޴HC*� ��?Y��i��O��XWQ���2͓ 6�33��pe�DA�yݴ(��vi��0�и��O����[�p]`�M'9�d�1���"����(�J�O��?���?���?���'f�(����'�>I)�'�L�^��(O��nZ7?�8l��Ɵ��IS�Ɵ��#dŎa�n�:4j��h�K"X�������(�4}j���}���PwťK5�!��SLh�P�J��|�'�N� �m���E������$B�ØYr�H85`�����.L�H���O����OF�4��˓��6hW�y��D\F��d�7!�΁��`B
)ҢpӸ�@�O$o���M{ѵi8"��s��?O��@A�L�;�,}kabߌ:����OY:� ���� �I���1�(��]��+��]Q�O��<����?���?��?��Df8����*�+�,��#�+.f��'��af�v���5�R�$��]$���P��*==Ta�6��siz(RƊ�?ɫO,�o�2�MϧY���m�A~��Bc��@aT_�L���C�8(�B��+��$�|2R�L��ß��Iş$;1%�%\AVC�$�$���i柄��dy��@�Qd�O*�d�O��'b㚠д)(s�"=�u�,�I�'�6�>�F��8a�	f���?E�Ä��F��5�W6GR4���K�6=t��#*ʭN�E�'����
=k�1���|�։<���ňւt�t)�I\Ar�'���'����]����4TȒ,z�@5����dJĚ-�X��ǣ�?Y�q��6��i}�z�6l�R�U;�|�u�[�`�]�&��9�4Tx��ƭ��<���Bbd�$�,P�~��-O�	xS�Ip�NHSS��6��Rq?O���?9���?���?I����	�0��Ƞ�@޴��P� ഑m����'����D�'��6=�F��[��x��T����jlc�6-Ʀ}�����4�������� �(��$	6	�����#8hRc	g��JH��@	�g5D�OLʓ�?���l��Y��.�dT�NR�7��$K��?a���?�)O��n�YC"%��ϟ�� �9'BQ�j��;u,F3��9�?� T��ߴz���O��)��r�!E�=���2�фX��,ϓ�?�s��&`"�s6�#����0��V#'�V�d��T{���a.'F�@I�&߹J�v�D�O��D�O���8ڧ�?�p Ш){��;w
�*Վ��#�?Y�iGN%b�'��&dӒ��
S���
%�5M_|�W��K	��	��MS@�i��7�	m�7�f�X��V�f����
�r��(�BA���������3�ĥ<����?���?)���?��M!��� ��� �6�`��%�����A��f�˟\��Ο�SP�d�'�2u���ۄ� 1�*�y����>)��i��7m���&>���?YCwʋ�%|����O:=������!����69�'E�L{��/.�b@��ĳ���1'�Br�E����²���e:�P���+Qc:�j")�$:�@��f�@�� ^��j�0���QRT���5m�U��/�>��[`LV;P� H���o� �K�*
��X��e+C�h�r9)�	P�^�����>X�.X�oUo�(�kɾ�u�Ë� z��8��ͺHd�d�'�U�4� ]@'
��y���뇠@@���@��N��9��¤t"�ᤫX� uft��H�`~65y� �mh�<��C����&�P�]=�U�3Y(�����ĽR��8F^�-g  ��4Qh��ChO�Q�<�kd+\7JB�a��x��'��'���'�*ĩ�;O
!�h� �ց��|J$0lq��d�On���O����O0����O����OMX��� Ґ2G		�,`�n�⦝�I^�ڟ���2��l,�d�88�Q%�*8H;�Ɩj}���'�R�'&�(Ѽs��'P���?�9n� .���J(:n�|huO����?��pK�8k��Z�S�D�'R�2��V,�4�3`����M����?qêU�?���?	�����?�1.��IڧJY��@::�*Qm�L�IH�B���H.�)��u� T�`E�VO������,=HL7����d�O����O��i�<I.�"A�E"o@L!P �
Vj&�@��Mᦅ:��7V��c�"|���0(�Fǎ3\d�h�^�Z��i�"V�@Cф\ybV���	X?3#�{=��o��r{�u��	�5N�1Ov����WJ�۟T�I��@{�W�E%|��u,Y�D�lyQ��M��`FN[/OTD�O���|BcQ¨麶��4�DMxV��t��l�`ЅL~��'���'T剁� �O^'�\T��Z�|���G���?��?�,O��$�O���cGG;O����r�F�)�0Y��D[1Od��O$���<鲢Z�)Y�3m���&�H��]�����|s����@�	ԟ��'�'9���������<��Ԩshݷ�Xi�1W�L��ӟ���My�k����$3�,̘e1jؕiRa X�4fN֦���͟H�'r�'�V�X���ܰ~��p�������Q��Mk��?�,O�@j�n���x�s�� d(�*ӽwpʙPW��+����2�i���������^�P"|���!�0I�y%��ّ
�k?� �}��#a�i��말?�����);�_#:��	��l��Lit7��O���,30��S����ē�z��<���
.ŬQT��n�ݼP�ߴ�?A���?��'>��d)0kG ��V��(\�T�F4Cƚ6�$�h˓�?9����<i����:S�����V>��!R#��M���?��r��x�x�O���'^
T��]=>�����B��TH���>��?�W�n��?9��?���$z��N��W��qg��R��v�'<&h�w�4�4�����O�˓z��kd�K�F���J���*����i�Bh݋�'���'bQ�$Y�*B j��XB��F�,_�Ua�#_�m�<��N<���?Y������O:�.�%/Y�x�&��5r&t�)D��'2�'AbZ����c^��� �/mh��E�Y���Q���А��D�O����O�ʓ�?	��*S���O7B���-.�l��l�0"�vU{�O<���O����<�JU��Od�Q����D�q�
�|�XyQ�t��d7���<Y�aPW�~���%N��`9�$�<9�$nZ矸�	\y�N'U%����d�k�[�oŴ���X[xr�#ʱ���]�$��ßX�?§�n�A�đ#!�%O���R`�D97�<��jX%����~���Bf����G�Ī��I��('�,@ �Dm�*˓5@~<��	;��iw��ӄ�'\3�l g��F���4g����iI��'���O�pO�雦UДu�F!S
~Φ��b.^?��nڐ��`�'���'���yr�'�:��G�����-0�H��{��՛��s�d���O�$�J� }&��S֟�|伙�,T�D6�}��Ϝ�J*���'���
��b����П��p��������jy��ϻ{B��C�i��g0��	ݟ�IƟ8�=tD��N�i)��C f��A ��EU}���"W��̈�O���O�˓�?�Lʯg4Щ�̘�xxT<��ᑨj:f�r(O����Oh��#�I���&��$	]�z�O12oN��@���Tʵi'*??y��?�+O����"R������"�
Ǌ(�\XAj��s��7��OP�D�Oh�L�Ifg��)p�z����d	Lqd�jC$���6�yP���I՟̔'�BôVl��xP��ZG�$�jE`N�@���M����'u剤t��OZ}�7�·:���ȡ�L�z��B5�i�RU����_� �O02�'���nD�P| �R��L6��&��6#��c�̔'�� ����p$8�fY�-ĥI��UF��0�&^�h��&k�d��I��8�I֟��oyZwDX�0s�̬q<P���W�S���Od�D�F�D�c�����&|+��.�i�H"�nȵǛ&�8'���'2�'���Y��ȟ\[��hɈ�LP+ ĐÃ�P�o�2�n�h�(����?�)§�?�c �F!���s��X�r`�w�Z']�6�'|2�',��r�U���4��S?�`��E�|}����<�(u��HW/u	1O�P$��P�������\?!�R[d��k�ESɺYi���צA�	"O,���'�R�'�2�d#~wܱ��@�#�B�`�ʝ�M�ɩa�����9?����?,O��g���}���B�Bui���<���?A����'�rD_.9�j� Ί5>8�����P	Cuv4�QAY5����Ov���<��:Ɉ$��O�h�JtB�Td���=9�h��4�?���?1�R�'�$��RF���M�2C�;BJPh��O���(����d}��',"U�,�I�,���O"蝷O��})�Hߵ��IZ�G�&�J6m�O<㟈����@І*��?O��ʂb?򴽉q@�.���'c�	̟�cm�g�T�'52�O��qfm�)z:�H�*\�6�,Qs�I?�I��x���Z
fYb�����Y�(�
�l���e��P�.�'���Q-+��'���'x�P��]�e̴([�fG�;��rC�Fur��?��'Hg�8��<�~j� %3�&Y��*��q�����/˦M�v���ITy��O��i>A��;J0���`��*p��B�Hރ1h�$j�4 Ah���aMa�S�O�B�%~��	[��"|�E��?r� 6m�O(��<��.O��O��d��() �V�F��8����7U�u�2BU-��'/��B��*�i�Ob�ĳ��K�bN-k**� �[4^.�`��!i�J�ğ�0b��?a���?	�{�gA1iE���ק��A�U���D�S���������ڟ��'���&�u���H,N��u�f�?a.<�냦SyB�'���'\�O0�$P�a<p�p�� $1f��Q�R-��}	Q昳(�����cy�'l�%!�ޟ��DK]Y�A�H��]0�i��'!���O�!b���{��&�*������bZ��r�,,��$�O��ľ<Q���m)�r�ĕ`���D'}��Ъ1�G�J��i����O�pR��ẻ'�j9�g���_�����l� BB�� �4�?+O��דi���'�?9���B��� R��Nc��;�a($�O��O&n�Ƀ��T?1#'�M�'��$ f
���& X��>)�+�	`��?Y��?A�����F�J̑"z���ԍ�?#�c�^���I�uRF�6�'�)��e$xp�ǅ>�0!�
@�0�7�^�?!���OL�D�O��)�<�'�?Q@� �hc�":&Աx�3,[| �u�i")x�([�阧�<��
-�z�17�R9<? `s�݄0z<o�ܟp�I��� Ky�O��'<���?�^iz��r��1AC6�|�<Q�U�<ɉO"�')��j� Q�+K��bҭV3_��6�'~T9uX���I��|��eܓ�|J�g4��%)�醯S�Ԡ�'�j0��>����O\��<Y�Ӛ0�"Ͷ�Ȍ�WG�3rp\I�E��C%�ʓ�?����?A���'��Eh�,���f͚�wݲ� �K�N{1�O��$�OZʓ�?	A����4��X�qR#�r�i��"�M����?����'t�@%w�p��41� !e��7X�ӣ�7X"Y�'C��'��Iß@j� BK���'�����-	)R鸳R�?4��i��|�6�$'��Ɵ\`���7� Ox��� 2q���be��TpI�жi��[����#]J��O���'Z�$�׾'NI���HY,���˄��c���	
t������!�~�ck��Q�4�J
�d���+�v}"�'�x���'���'K��O0�iݕ8�#Z�>!Hh�Q
����0�+�>��E�倣"_~��|R���?��ф !��@Te��^k@\YS*�-A��)�.�B�'bR�'�D[������	�/�<��1�@ ,B�B��8�Mk�'��y��]�<E���')�(hQ�ڑČ�2�$�(g��v�kӘ���O����,��|b���?1�'��a�I�e��<�"c���:�y��%�:1�p8�O|��?��'zd �' �V�P4sÎ�0ot	xش�?�Щ�	��d�O���O���TO��'��<��9�4ʡ>�6�F="WN0�'�B�'sB�'��&U#TVT8�f�r��կɧ|��H�
e����O����Ox��O�� Kp��rw��b�&�������/���H�I���I�����ğ���ꚩ�M�A�U�'������
�1�\��Ʃ�=JD���'Y"�'�R�'F�����8R$w>		�G�5y �s'H�IB���3���$�OH���O����O�Ѳ�$䦁��ԟx�'�,Z$MABˑ<��EacgF��M����?y����O��W8�T�����[b]�=2�eA.g⮸s2Jd�<���On�d�O
��D����	ϟ��I�?�X�o_ eH���ƱmN8TX#֍�M����Odi�;����<�禩Y���Y��Q��%E�v�qQu�<�{�虠U�ib�'�"�OL��Ӻ��j�U� ���0��H�Џ �	�I؟䲡#u�$�T�}*�JO�2���!�/,�IqO�]�B@��M���?����wW�\�'B:@�KQ,5>d�wn�O󘔓TJm����A1O��D�<ٍ���'���`�]SfR�I ���'t�	�t�k�T���O��90�^t�'f�I����v�V���H�C$��� �%�$im�ȟ��I�m��af�v���r���?Q1�
�4I+��((����:����'���z���>�+O �d�<����d��pd��r�@�x&�ʂG�f}���y�'�B�'�b�'�S�΄��ʁ�E��d�d)Y\J�+��3�M����?i���?��Q?A�'�b��+<Æѧ��7e��8���.9��y�yb�'�B�'{B�'��l�yӄCQ���lP2*Û���f�馹��۟���Ɵ��ITy��'�j�Û�M�kT=%ɱA��p�.�h�
A��	���I�$�	�t �����M����?AU�-��;�C����B��#=ݛ��'w��'��Ο��'r>���^?!�#�wʰ�qk�	�,�;�m���i��ԟ(�'~<��~���?Q��L<�Ѱ�W�w:�b�B�o޺Z\����Пx�	�+Yx��z��'����U�r�9W���~p��s����4�?1�(�ʑzF�i�"�'�B�O7���'T�1�c�/�x�mK�-DzI�p�>��� �(��?!/O�(�ā�7%��2 �tt�!��&,�M�$C�6�O�d�O
��������Ob����?��!����!3��g�KZQm�:D��q��(���ę�t�'�l:5�Ӯ2�q���5^��R�g���$�O���	E^���'2�	�x�h��T��N�j�j����Ɣ]�(n�ٟ����d�K�-r��'���?yS��3�ZpO.Wي�s���"l���'�Te�eE�>�)O<���<�����N���q��;'���s�`	l}����y"�'I��'+"�'s��'�MP��^�}�[�I��z��1���b��7��O���O���}�Y���	34HR����F9y*�Eo�py�ok��	矠��ן���џt�I�	�n��4���w�Y�<%Q�r�_<�N]��i�'0��'�^���	o��s�}��)��I��X�uڌ�ر��>1�Ų�?��?���e��U�i�"�'��9���L�r𴡨 Gʶe�pHBvFl�4��O����<��]�P�'�?)�'��5.Z�	:T(�	a*�M+��?I���?I����h�F�'���'=�To&3�<�ې��7�<�"4L���7m�O���?9ҁ��|z��?�Q���|n� ?�]�OO�����6��6jx�6M�O���I�m���m֟������S�?e�	�k�<���E��7Nb���N�5�l˭O^����"G��D�OF�
�XN�i/��G�#�d��ڥ^��(�rƜ��M1C�l��f�'��'���O�B�'�b�_�;v6ŉ��+7�0I��d�3BJ7MҚ��$:�4��������&�������_T,Lr`�ף	�r�oZџ���ǟ "'\��M#��?����?��Ӻf ߫?�ȹ�D�,x��W �����I��|�o��B66�)��'�?���|�tx��:Z_ʭ�����h� ^+�M[� ��P��i;��'b�'���'�~
� ��I-\&#g���f�*^x��+#\���&
���	ٟL�	�x�	n�TK[�=��@#��^x%�d[�͌�#���S�h����O����O��O/�	�8�5��8r4mIV�S `��D߀J�.�Iן\�	П��	�p�'�����r>ciZc6v��a�۩*9X��,0���OP�On���O�ih7O.M[uO\�l�j�� �(c 
ٱ�c�X}�'	B�'Z�I�^u�M|2��7�f�Ə��O6��[V��U����'��'���'�d����'��X7>�J O����"v[4@oZ���^y2d
4w �F������T�&���f�D�.��`GY���X�ɭ>|�^�~B&�v���b�E��/b�p��Ӧ��'���h��k�0�OP��OC��1 y�/D��^h��bJZ;�4mZ����ɸ B���_�Kܧdڊ�+���
]A֭c�F,~�l6�NpH�4�?Y��?�'r*�O��;�+�94��!���ϴ`S2��0"[ʦ�3�B~��%������V��٢���!cO�a[�-�<Y��0�i�r�'HRD�F�O����O����:]J`Y%�)p�ʼK�H_,J6�+�$�X�Z�$>Y�	͟��	�<���Fo�-�K����:��ߦ��	f��݂J<����?9M>�1H6�����NA\�5��'��@J4u�'��db��'��H�I��',�@��l�Ja�y	A�#`x�Eb$�^5c��	I�Iޟ�I�Ba�[U<xge�d��A�*C?l��'���������CyR�2��ӦUbz-a���-3@�2q�Ɖ0nꓟ?1����?9��= �2��M�d���B������z+���Q���˟��	Ey��ʌu��2����iARm�#.�\��%E�e�In�Iʟ`�IH��	j�I�Fͼ`*�(�imD��瞧Q����'�2]�$�B@��'�?)��N��u ��P����r��Z�2uR\��x��'db��)&��|��L̹R��Yo� ��S�/~�
԰iV�	���4��4g�����S��D�2eze�?�=ӅG�s�F�'���K�s�2�|��)�}���\�O��3Y'a?�8W�T7m�O���O�i@j�i>5�u&�S�J��7�*k�Ȱ�&kU)�M�ԉ��?�-OHQE���',L���Cu4��R�V<)�����h�����O���۷rZʓ���O|�ɶ}��L�@BK_6�P@.����b�����)�Iޟ��������N1LhVHhT+IuZ�h�����M3�/�Y���?��T?��	^�	1L�|$�v�L9*��az���v��e��OY
���OL���OR��O���!f��Z�jMQ$+oo���B�,m����O�˓�?�J>��?QM��y4 c�a�l�JrT�%1���a��O~�'M�'剞N�2)O���jB5{�^T:ġ��
�H��O����O(�d>�I%,�|�"Tيv�_�ؑ
Twt
��'_��'�B�'�"��7o��S���� &O�Uu�У?��gE��M������?���tzh����}��8�h{B��=�5�ؔaB"6��O��$�<q@j�ze�O�"�O��R"��+�$�&ډDN�4*�+-�$�O��dܤ7����r7���;� �sꟓP�nZpy¢NT!�6m�`�4�'@���)?���Pպ��Ӓ�f�ÃTӦ��I���B�:�S�'0K,� �g�	�P�gkE�C�<5m�6I���ٴ�?Q���?���*:�O�� D��D<8���x�X�.�ꦝ��+��OA����d@��I��g��,�Af�7Ad6��O<���O��#WL쓴?Q�'��1�⏵ؒY�RȌ$5���B�}�Y*ј'2�'��ǈ�?�xI�O-;�x�k� �H6-�O$]��g�O�������Z�i����n�s�v�Ň�2����ǡ>��m�v��?9��?!.O�Y(�Z!��\��чJ��@��e���\�>�����?���ö�z���㒁��=R� �Bw̓�?Y���?�/O�!Jf���|�@�X&r�  r��L7���'���I]������W�|�,�򰃴�ޏR��Q�V��+�˿>���?�����D��b�\&>�al?%���6�9�|!A��M�����?���S+���>Y�؏&�KS,�Д�0h߲6,�6��O����<#l�1<�O���O�~xh�ƈs@�H�IR셚G�.�d�O��d?1K��yt��i`���ǚL+�-�qH�oty�L1i9
6�^}���'m�� ?�G�4?�Ԉ��E�0O(Г��-��ڟ�;��$�S�'kW~Y*�C�,��)IvȊ�e�9oڼE` �ڴ�?����?��'<T�'��ϒ�e,��s�E-A�l�CdŚ-�f7�3E"�"|���1�G�T�iE<Z��~�9��i�"�'�	��&?0O���O^���&���6��dm�a�GM#<#�c�<Ȃ")�I˟���ݟh3���K>L���ՙx]�8�
΀�M��IR��$�x�'��|Zc� L��f�Qu�r����k#��R�Oz�����ON��O�ʓs��! ��,;�0�p�N���M�#g~��'-"�'��U����ğ$�M�Iz���&�6BIx,��D;����3lPq"�܃Bw�h�RK	(h��s&�֠;╉�lT��:LX��E�q�(�xk�������.���)� >�&�"�=I I�8K~���S���%>Q�왆��0�!�P�Aa�BS�̙g����j�)[�N��#ˌ.����CF�}���uiG>"��H��
kP��y�o�3o�4Bb%Ē�B��FK�I�^lS�(E�&$uR"��	9~��P�E�P�z��CӠ+.$�����>Һ!�&-	�]��k�ǝ1R�q�c��%o��ό0`@B���(?�-`&FJ��'h�5*aPv����耫TN���#K�5V>	�T�� zo� �e�ʘ{��Q�k0}�.�"����ӲS�|j3�M��#i#�����rFb�C�Hϗ�VB�j6��I.9��$�O�}���N�p�d�$Q>l4Av�ӥp֨�ȓ�.Q�Є6�@�`�ͫH�Y��I��HO<M�Ъ.J2]@G ��D��j&G�Ԧ)��矈�I�c)\������,�I�d�i�9kqJ�
j���GG�mmlY7��s�N����]�p� +R�6��t
0��B�,�a1c*<O���\�.�I1� V'GKʹ:Vb8�&EK����|�+$&���5eӢ{�Z����yB�ή!P~1�#u���)����F���hD�c�Y3N�4�p"��}Y�|�c�S0d�%�o�O���O�d���?y�Or �7�ԻIWR%�eL�YK�}@���v�L��E��z=�T�"��$�4(Yb�'�L��� ף+��="`�ʞD4Y�����M;t'S�~b&�x �=+3�!�����(OLK��ٌJB�� Ν��:���(2� �O��: �Ԅ*'d堒/T}>\�b�'��'�нca/�<i�`�W�����y�Dh��O�s%�p���'�ݲ�N�2I�'e��0q���'	�&G�C�'��	��8���֢��&d���*�-Q5�%S�@HJ�l0���{�ԭ�D%Q� �ܸ����GE#�1Gc�_����]�:
���i	x��(1nГr�BY���@�(�-1��3X�'��	n*^-�6 �I"d�Qv���;�(c����I4nǖ��&
�q�*Y��FܾB����M�oN�F�Έ	Ǥ����rDJ-�?�,Oh�k¼@nҟ��I~�$�P\I�C֚.�(��G�B47��US��R1b�'Ħ� �Y.%?�@2�e����a��
̯�PU# U>5R�O/۔�paȺV��<Ӈg1}rϋG����	�r*�B"AV�It�(��O�t��@�48�!�[PaK�L�5��<���r�)��< Y��� O�zT�q2��:1B�	�y�*��p�'.=H��d�$,���D�z�'�X)����5r�N1�q%�8�K>p��F�'�"�'�bɃ�,MMu��'7B��y'-ZڐLp��څJhm1���1������']d���Ò�8�� 3�i5L^eq�'� �HX!_�� #Q�[8� Sk�>Q�\��d���(����"̋��O�TH� H�<�� �3�@�y�){�VHّ+��S��OXX�������Y=v��5�O.mz�bĠ��Zpĸ�ȓY�4DBG��,
"h��v,�U�"��'�#=ͧ��z��s�A �	�F��%��X!��2t�TA���?����?!c�����O���]�J98$������شV&J�����P���[p���_R�j5e6Z��xv�	]�H���͊5���Vg�&Q76��Ɔ�?"UY#�E1QuJ�%�]!]�\Z��ɤ;0h�@;�^e�WEI�c8�=�6��O���>�d�O���:�ɕs�lS,Q.o*@M�'O+KB�I"]e^�
�+��5N�cK#�qO:lҟ�'�BM�!K`ӄ��OT5�ç�<!�R�3�*ɨU*d�So�Oz����l�����Of�S�$�[���sf$����������
�ů�]��ıth�#u�Hd�B/^n�Q���]`̨v�H�y�<�D-�:��P�E�
�fEj�-��j�M����2?��C�	�;�n�d`��F�0�G�PD�&�%$hB�I#	gll2�iP#�ґ�3-���RB����M�	�$'��б��L20����U�[� (�CE�i���'!��):ư��.a��ܲ�^ I�X�B O��?4������@�M�0�Z1j EJ1a����Й{ۚEӉ�x�ԠL:@���F�	���G6��IW���g�W���%{�n�`�@�,}�l�˟:�Z��XqŮ}Id�I�d��m��>�Șܟ��޴F��V�'��ug��q;4��f�;������$�O���hO�Ec�`A'���a�h�b��<h&�'�7�Nܦ�$����f�b��$[�&�;�r� ��9ir�����T�im���B'���'l��'���ݰ&�b����g�����kW�F4��
c��%a��	h�42�N8�3�D�fiTp�#�H�ZPap�V�{êYjGB��cZ�d]����L>q�+�0G�p�"DY�����P6f��'�����S�g�Ɂ��LjE!�dH	�֊ؒ,!TB�I2��tAq���)�JE�p��l��0����t�ɕ"O��Ӣ��8B��䓼9�<�hp���v� ��������ϟ��Zw"��'���	�h���F��sA����:M|��8w
УU���)���CE���d8cɖ�����_��W�G�E��[����0`��B�H;����Ԕ��`�[M��U����0�僀�'ü7m���!�	`y��'��O� !���4��)�Ӥ��>0 �B�"O(�q��Y���m��Vc*��4�d�0w(�$�<9p,L"����Or�䉦k=�@���b��q�� ��_����O�dд��O���m>9Q�G��8��H� �Պ��&�p��� t�-��:O���'�ɇf�D�OL./K"�T�,�8b���p<�dP��0�L<1G�/FJ�$��?�P�0�@Dv�<E��_:�8�*�A��x��^<鲵i6�8*7&Ad�B�rO����8Jv�|rb�<��6��O����|B�+1�?Af���)d����c �D@�
	�?���\rM�����򙟄��+�U~�Q��}_�Sb.!}����O���{���'c�a�L�H�tPv�>1��͟L�H>���� �J��v.]/l�쨊V��E�<a��Z�pgehTJ��v�>lrߤ�0<���_I@ ��i�.>;@����P3:�`���4�?���?1V��{,�X��?q��?�;J��؋5��:�he" f�#���ɍ(j/�l��
x�J��#�*p�1��'y6��� �u���Z��JDjg���d�$�TG��:2�ŀ~�q��'p����Z0vL��cN��U�
i۰󤁿U���L>Y��̮TqDɑ�ɍ1>v���Z�<��ƺVr�KB��,9�z ��+M~bk5��|�K>Q��S�v ��
�K@�^Ob)CF��d�8�F,,�?����?���q�n�O$��}>�"#ʋ�?����F+�8�&,Q��U�ut��* Q��|�0J{|�S'\�ؘ�e���ag�����&���Hó�0=ჲi�$걮^	9���R�S�YS�{��,�aD��*���+��8A_�kU�yb�������AM %>-p�+���'��6�7��/{H�mퟄ�ɾU��9�C.l^xt�!�ۓ<�������� �ş���|����`�����
��!r�.\���g@�)�f����׸0D ���MC ڢ<y'@�)��	��̗�(`��u�7'&de��%D���lI4�N�Y�Dt9��<yף�� �L<Y�$��Bx6��� V�$��!A�g�<�#�$y�ڵXGl�SlyHsKN<)ԺiDb���T��{SE�4|�S�|�C	"�66��O���|B�X�?I��v�x���٣c�H�c���?a��$�F�5j�V��t0�)�y*�˧h�!��I3Wh�9$�V�-|HO^lXXL��ۣ��	Z�t����iB�"�|g隧I_� !Ғ��L�� ����S��tk�ġ�cK&hAD�`-]�Q^$P��:��`MŤ^���V�Z�L��y����HO^Ba͗�o�� �2D���h�%����	ӟ��ɍ,��Lrgퟸ������i�yZ��\�#<U�&�^���A�:W{L�*O�����	�1��'�$:c*�5i�4%$�Τ4^K4�ľ ���5�^�s`�d�@�H��O0�́�BT�<	�ǀ?�����A�����ɀ(/�'�����S�g�ɀ�pQCM�"*Xb!�o̹|��B�	�y+n�D��)�l����|���K����v�	�t�����fF�%A��
�نP�H�Fɚ�3|��I柘���Ȑ_w�2�'�I�>]X @k�H.=��"���X�@����f/Bdr�_6b�B Ƌ9��+�B� �f�1cP���2KӍ���#$�^B֤����t�bU!��OX����N�L�1­޸#ֺ૔�#j���4�O6��HK�(`z��'��g^`9:A"O�,��W'`,m��C�Z�d 8���Ԧ�$��I"kº����O��y�JʤLo��90bV�2���r���O��[ 5.~���O��0}n�3� ڗ"����	M�ƀ!��ݽ�X��c�'�f�!RBA�'��̓@��:�A(F�u16jW2`�Lj���#2�טZ�џ�+��OZho��d
0��a���֫J�x�����'\r�'�@�� (��B>8�q��R���Y
�'�7m7W�qz1n�;=��K�h��b��D�<����R���'��U>}���B�����E�u���{�ơn<L!Fc�ܟ��8tO�����
Q�tx0C%B����ʧb�jp���(s�z̐��%BX:��O|I�b	�.[�|���J��B�v�2�E�|삤���Pl2����.(��'��d ��:]ɧ�O�^,�T` 1[�I�@�܉@3N�!�'j4u{w��9a[�l�%O�%1��}[�4j���0`�F+�z�@j��Z�� ��*I��M����?i��PnVT�0,I�?I��?��ӼC%�ЃTr���`� ~|�ՠ�̞�Ԙ';$e�ϓ�Ȣ�+�\y��B,�l���=�mPx��#@5���� 8s* p"�����p*0�)�3���(V).���7��Y�QQ!�� �:`K�'��
0Q,���*������ᓞ�	���5v3jl��C�	�)h�\�RF�Y�Iß ��Ɵ4[w�r�'`�I��D��y�F�[�@yÐ��3C�4Ofa�%��c�/ϗ�4������Xr!���%#h] �J�^ |\p҂��d-2v�'?�r�Xr��UqE�*�D��]#�y(Y�6�� ����U��7�ʰ՘'#b�,q��Ћ�M���?�����Q �ɲG*V.�S�隨�?���ΐ����?ɛOr$q�IE1?:.�R�.����IR�ۈtk� �I�tO�y#���uџ���P� H �lڒ@(�J��J=�>`�%G�G,$�2��j��0���Dǔ'Ҥk�v]�'���s-��	����_T/�X�'���'3�O>�z�i��Y;��	���6*qȕi=�@��4�p ñ�$>�2ba��s���;���X07��oZß<��^�$l�u���q2��A3�OL��d��4�"�'sp���'�2=�QkH��'���]�R���H=��}�#cU�_�2��$%7iv��i��!�!0��c�H�sB U*]�=�ځ�I��S��� ,Q�#I��Ӭ�'R�B9��"O��y�

	M�8+�K��'h�̊��'��#=ٕ�9e:V`�k��$�z����Z8��'�r�'ڰ�0w��t�r�')���y�M �SJ�)�$[� H<|�v��;��,�F�5>Z1h�$�Zs��|���/�=`�k�������ۋ���I��ܗaϾ��2�W�Ly�Y��L>iJ�2� %��b�
a[x:SO�f��'\p�����ظ\�an��rAD��Ǜd�����|q 5'��V�6��XP#��'R"=E��FE�T~V 9@�J<����62D����% ��'���'rT�����|���߉G��:4 +�Gѵݦ��:c�h��P(2�D�r��R���a
X<QPE)�׍�8z�-Aa��cZ�I���?�A	�x԰��Z-Ts> b�A^�<I0
�W�x@��%])�8�����̓~*�OhX(�k�ʦ���џ�R���� � ]#`�՗J���J��]���ɺ`)DQ�����'��=
vD��y�h;��O��r-�p��t�a�۟d6��q�'����-��X��� ȡ�dغ�ò9�*�����.rp(�C#�J�:���L�h�b��"Sm�O��%�8)4'K
HIp����kH,�9��4D�ܪ&g��0���R-C}�uo0� Qٴ_����hV���@B՜ ��M>9qf���F�'�B^>���N퟈�3h���T21��ES���f�ڟ8�I�0|����|�S��O�X�2e
�X�rh���VG�jX27�>��iRt���O]����ܠj���dIՒX鄙{J�P;�I�O>'��?m�-2v�Є��ҭRB���I(D�T:��غA�T��$դ4Hf�P�E9O(�Gz��F�Ykt�{��=N�~Ě�u�j6�O����ON� P�T<K�����On���O�Y^ā�$��"�xx�VF��5��S�F��I�1�ƽ.5d%ps�ԃ�OY�'�r!���=n��pX����lA�4-�"��e⧍��و��Ȗ���O��'-鱄L��P`����Xd��'�d��X`��L>y�̕|F�A��ŗ��U�6 �w�<I�I;n�$YcE#�{����IX~2e9�S�O|D�Y"\:��@SB�D����T��Q`�'�'��&�~�����4�*!��� �@0*]2�b	F W'.��Qe�6�蔆�XF��C$��W��U���fh��u�E T��%�&�'�RŊ�'�{��ds�I8�6T��jՕ�?y�i��6M�O���?��2%�ښ<�6)ƅC�]r�M���y�I�'��E3��!a>�J�,ՙ'������A.xI$�m��4��\�	@�M�:3:P�2*[���\��ğ ���ן\���|zP�۟x%��b�ˊ,<;|ݣ扜PX�=�5b.O~P�6�$ƌNKRaa��٢���fT1a��x�	.�?	�xB`�b��H����U����R,��y� ���n��̟�N����3@�x�s�v�ϛK�$*��'v&1�A� >m�8�	P��
�'��E/a!D�"Z�_��e��l��JP�'�.ٙ��'�1O�3?��OO	4ҰPaЈMZ��Z6+\b�Dـ>���?� �χK���͞�lgp�B�)/}ҥ�=�?���|���/ŏt� P1�̏'n5L�����yBcP�[¤��\�A!J����I��HO� ����@\EF�`����>hP(�H������	͟��	8% �١H ��������iޅ+b��]����ջ�X�x�'�Zȅ�IKfBA�*ܗ1�X�l��2z�=��_@x��9���	��{3쒻j��qC����i��a�)�3�$
"g��!�h]�����kW,�!�$�]{z�;�͘�<e���``��V��I��HO>�f��"�dă��ܸ-�=�2��M��X������	�`��
�u��'��?���:����K���mU��c6�Ƀ@Du���e�.�ࠏU��M3Tc�-b\����R<���UC��D%�1^�J1I�h�'���	�Ȱ?YdC��Y��V�@r����P�<�pM�"��i�6�D�7�8𲅪N�H �Ou[0�SȦ��Iӟܐc8��u��cI�:��a����۟��Ic������<̧�\��z�ɾN����/�1|K@у��Z�V%X��D��&��O0pp�(\�'�l�*H˩|��Eqg�'��$����1��ڔ�Y�@\h��I��r̈́ȓQ�&JG�1%&x� �Rt��._���I�&�P�#� �/>����qA;��'�@�a~�D�D�Oxʧ7f-�
$�a�E,!��l���im����?��O��?��y*���2����ϞLN���)S%V��'�B Ҋ��)U�m�$� ���V�B∊�d6��|��l�S�'z�r�[C�^��I A�ܗ����ȓo���#�h0��S���;������HO���.�{v�I��8+��m�se^�i���p�I?/�˓J�������iީ�w��'��Q�E�
�b�D�	�ςR��s�O�!jn@�:w��$���|��Ɇ�<��,vdI0&�� Ɩ�#�O
�E?��H���2c"1!��'c����8�ӨJ>�,��:O�� ��"P���c�#��T)���!Yl�I�V)����|����k�a8�/ )`����0���y2�ܔ������2R:60�f�U��y��'��"=ͧ��^��r& ¹*A�����6�x%p!I�>qƞ����?���?�6�����Oz�S�n�PD��ϳN�����+]蕣R�)�X�ń5��A�r����c#�A��ᢶ��6�
�:�����<�����"%�4��28) �(�kJ�a�I�Ͱ?iT�]�`��X�/'j�	�F�q�<9Ǫ�wh��Q��U�섡�*�n�*�V�|�/��xX�6��O���� 4$R���V��@�0d^<L���$�O��S��O�v�z�� ځ:P�ΰ7&8u����9Q�� v�%2!�M�R읤=�h���,�W&&�[��	.2#rMAQ�-�u��J��cIL0:u�ӚGa��b�4�*��G	#d����	r�đt�	5D&p��R;pp)*rCP�q�C䉂'�d)7��F`i���[iB#<q��4���nڄ!���zO˛I�� �O{�I$�<�0�@��M����?�*�:��7(c���F'R��	�ڸv�|����O��d]
Wh�c�Di�䕪vF�>':-x���"1��'#f{��\�r�5��HؠŦO�Y�bl�	;�|��7�̷T�v`�Lߵ)֔��ɟX�(ݬy\��R�"F�����5}�BE��?9��|����ț�Ȥ��x+N��!�ybW
{w���-Qo���8�Њ�0<A��	b��xB���5^�<����%B�fq(�4�?����?p�T6�5���?y��?�;N�������-�PT��ߧ4���z���$�MS����f���g�?_�1��D��@U$�y�J� )�QB'ܡ�V�5Vh�p�+1C\ 5���O��Y`9�f��}��'v��݁u�v�e�q��b(��s��"0��{u*X��3���)�3�DO�
�#�ō�]c �A�-@�p�!�d[w���s�@�6bL�$��.~h���O��Fz�O0�'� @��WB�r B���kt�1	�'M­QR��7��˰͔�f0�`�
�'�F 膩g{D��`%�8g��Q�
�'-<��F��.[Ř�iHA�Z�6-�'�d��$ �0�`�"����d��'�X��	,q���9�>{@m��'%�Ę��ڏ�h�����rȸ�8�'����E��U�
tKG��5l)<d��'О�bf��{Q@�R�e(T"�U��'(�(à�<�%�Ǉ�1\RD���'t]8��."�H�`Ɠ\TTI
�'���ǫӓ/t�M���Y�D�(ex��� Vp��[�"���&OX��= "O�����#86*�孍�)�|��"OhxQG��;9�h�B�T$�0�z�"O�mJJ�;745;�͛Jp��&"O���E��mi*��5/.�؅K�/�y������(ۊ1ypp�eN�?�y�Ñ(At݊R�L�#���`eN��y��9:۪I�%ٝ��Pe�X��y��-r���J�ەq�(y�Q�y��^Jc�����ٯTE qi"�	,�y�jV�Xt$�
�� 	�!z��މ�yb��0�`-k0�	�U�t�P.�y"��/ނ�ڣ&�A:PA#p�J��y�c�1r�`r��Ɇ'�"�Ҋ���y P�^�p�悛0*�zŨ$�@��y2��B}|�3��+�B��!��y�jR���=8�DMr/�x��E��yR�׿>�l0S��Ʒ4yd��U�G��y��e�� �9�0�U�߻�yblА�ʄ
�"�{�p{�aބ�y�	�""���"���
&��5�����y��� ]���($J"Ѳ��R���y� �7��6�&�2���W��y""O�;#p��vJ��!~h���D��~����t�G�(N���/�}�gy�̀6,����5-�
mC:Q2�e��`]i�f��=S2��
�2�x�3h�*%������Y .Q>a(� F�P.~ܞ��f���w;��ڳC�4/�j�ReAX�?���A�?��!��E�>k.��JC`��zX�����F����J�O�D"e����O��ة�,��'l����RgQ2?b��(�Qd&$E|�E����-H�W� �$x%�ܤdX�D��XF(�8��L�NՎ J�Ɏ�Z�~�a�®c��5�P��$�y�ɟ���
�ٿ 4��c���*�8:�f��	F�^V�y�6g���h� ��_�3?9@`ݴ2o�X*��������NôC��L)����)H�;ߓmԀ����k$�����%E�Ȕ�B؞0�h�F
H�<]\PPP�\Y���w����g��Jǰm�'f��|���1�	U�3�NW�?��*G��"At��&傺4V`!��I\M�D�%5��@�O��,�I���'\(�{m^9vVd����A3KV|F|�U� ���)�ƚ,w9jb�Z�8�$�3	�|<y"�
�l���ϞpR�0���׳g®��2D��az�˟��,p��,\��V'J�:6jm"S�~�@ɶ��)��u�g��r��,t�T�3?�Pꛞ݀$3���h��ӁjC�N%���X_਋
ߓ ��b�ȃ84}�Ӌ�lm��K
vϊ=��I÷=X��_P���w-���U�K�b��)��/M(��T��h'�2�B�E
�Wg��!��#Vb<�%+NA�DN���Oؤ�zqnN1��d-��|��\�[�����C�o>@96UK�'<b�IVk��W�}����'hG��h��O�	�.ź[o�����,rn1r�'���x���/L��a�w��8_��X����'`����H��C ��8p���K�'(D���"ƀѡ�L*p	DP�����q�:a�@���#�x�𦤔%D��6&KL���wL�O���� E+��O�����Fyt��(�nڵ]�` 8�,ؘNnŒC�˩rl�\��sH�)�s�7-�ْ���B����.�O�<p�|a��X����G,M2I�v� ������r�9D��g�X�)��+���D"�L�����]�(��f�D�V�9a�>�O! ���);vF��ugϽ��I���I����ЀW�m����e�4/L�UAIj��h��|���w��'x�hY��ѥ$4����#E���Gx�@@0p�а�'��Hi�c�Ƿ4A��i�T,�hR�����҅7[,�(�C�"��w�,�*���x��J#Ԉ�B��j�0#�.U<X��3�	Q�(�٫�"mRā�[3g����\�u��%�������b��4Q5�ΐV��S֣Y{��4p��U64�a�P��/\�$����D#)\�!ÃԦ����~��Χr��g���t8ָɀ��j*�hz�X�*=a|�O�o@�T��U\�(�y���Y��	��CH�*�r�$���w�^X��卲K0�V�E���%`	�K?	H�ϓ�,-���_�/F�p!m�� �`a�}2}�4ʕ+)%��A>�O$��`�� @>ҁ�xi̻DJ9�,8�͹��L>�0�Ԁ6���#DE�;�앃�D�NCLj�JB��a�?iG�'���)��y�/M�G�ޤ� �.^V�1��_<z҅yP�'A��q�w�*��W�]AP��r�ڏm���pM>q7O��r���?�����
�Ԭ���ֽz�ح;��l� [e�����ٸS�5��U"�%�?� :���$V7F��49��˞-d6�`E0ObtaT���L>A�씚n���OU���2A�.b{hM`i�=T��$8�'�d� ���$V�AaG[�#����6�?ӧu�MK.����` �._�v`�p��G[����Ǻ<مI�!��>�O*�7kY#k2���[�y�0	r �� ?3�4�.	O�ěs�|�&�<� ���<Y'-��E������Ŕ8o҉���5R�Y��
,�^���^4p&�.��*�Ɇ�R!
̎����$��L>ar\���PH5�$N����<*C��wlx��K�f�P��n0�������U� `�Ҥ0
��x��n� �n\�V,{���`U4��h6a�'ހT�0����~����%�4��^53'���@Q4��եȨ\B��Z�7Oz�M݊��!lόe�^41#�7&�La4��78Yl��#,Z:Y�	s�\�/�� æ���E0LcH|�<yc�ϝ1����gD�V�<�S�w������\�F�jq�`�Ӻ��.
0�3�N[ �Y�%�N��T�ڧ$@��3W㔑ER��Y��$O����6x��Jf�88!��ͻ'��J<q�4voj�Z�ۢ���~�O�L����|9 �um���蘔�	�Iy>݃�'# 7�L��>]�擣1��h�'M{�d:RJ�D�.�D	�F�R��'�4���Xu�L��`�%���* ��lD;%̍�}?���'8~�*b+�	!���5�>�~��g�?����u"��S8���h�:F@�3��d	�z�@�1���-��x9��ʳP/��0�ɜutܘ�We��l�1Oܙ�Sm��,D�=	�`��[C����'�pD�> ��I�"O�	&�l<�U��H����t8���Cʓ+R�����
�e+r���n��X��=�&m�(��AY�*w��>��O�	�o�$��}2@`Ip
�='�BB�Ue<A�F;�h̛��Y
�	�M��O=�I#{Sh͙��+�
�RQnP�I�r����KzZ��U��!-y��:���������	0A@����FxB��cNn�!����Ԥ��ї��D�,E��"�.E=X�%C�g����h�	�M���5��T�r�c�V�����@����]��&�>Yp���rt���kvN��R'�%g�(�r!7lO�̻6�X;Q�S2'�c"K^	��i�őUyR��Ly��)ѐz��`���h���$��`�#����O�"Akǧg���P<i=xE
��i�:��*X��,Rw)*ئ���'?T��'԰L�ɽG��	��j.��'���V?W�	
qi@?�p9B"B�"0��$��T�aD�d�T( ��FSײuaPߟ泟��5MԀ�'W9bx\1���8QZ�4p|��(C��K��5���Ǻk���,�P��8[e���RdU�H3���!I�����fY(�?�di�<�Χ<�Oz�1��Ӫ!8m��AqJ����:c��{��E;wj�X<����E߻F�i�B���4��A�<9��Od7��A+m�d�1�O}��P0�Z�~gR������c$����W�xI��\��R1�q�T#��q1��֞B��DY@j�.O�	� KW�y�l�+�_�E$���8�)�&��`�����'W����Զ
�
�S�T���'�\L�D���5zT��s-/�Ll��P>�o�8R��D+�t��/��sK��رƋ�cEz�B��\%Hq�hz��ݯ]�џи6B٨z3�����<D�ʭ����+����3K|cH��̚
�n�}���p>M����
a�j� ���%������?��`�e��+��{� �zט"(lA� �_�,E�U	Mˬ (��.�<�S-ԦE������A�]n����i�
Ҫ���(�#��#3��#$���zش1:i�r�փT��aq ��Ԧ!��@%iR*��݃f+�T)����a�4��۴aV�9TlĖ.�2����UӪ���ȶ|nZ0s��9��"Q��
dA'�VI�1s���:�t�T�P�P�rPk��>%?�i���5��9T��xFj�   ݲ��H?aSD��PB����(TF�?Y�fN�jtԽyC��*?H%*p�P?����;2_�Q�G&I�G�O�%��g�Ɯ��@�(Ӝ�K�m�}t2��T�:t��6�9<O���D�X�t��0��Q�Dkc%L�2yj���y*��"G7b�m�R�[����&?�(�lz���т��ژ,���$E�4��W(�,^4h亥7�� 7�^��D�ȝ)�xs6`��D�6M˫<�0��-9/N��꧈��&��c0�P�,X�2Rm����tr���7
,�)%��V?E��'�EXf�]8,�`�Uw��4�O�E��iї@K֩��̀��O��t�Z���箈8v��	��?O,Tw�9&�`�!�0��'�4�B%O�=�P`�G(�V��k�47(�A�%V�p���Wߨ�A	 6Y�(�bh2$�J���دp��ٓ
�LF�OR Q���$�蔐��S���9Ìt�5�Ĥ@S�$�JH7�N(Gx�K�9�8�Vg��)A&��}b�BӲhs����4��\CǏS�iXe�6}�x�����+h��s�H58DD�g�eJ�Lk���p�L�#���3�@H�4�JE�����1f�"���&�7��DZ�mh��a�\2>Д��D	a剅2I�AQ�J1,�����4Z3N����.�,}�a����M�1�,8/`����+�&Hh�Bo>�	�J3�\�m��r'�6m։H�ҙ�^����d�!r��Q�#B��p=�t��!�D�˖-�)h�*iᲊ�-��L��d�vo��� ��4n+(x�]Dv�(s�H*H������T�3�R@@SA�&�:���O(F�0��UI6�#<�`��:*E�UJ�E�0�`����?�	(��8Qbפ4(Tz��F�Zn�¦g��W�fL�D�R�G���	,���x�b6�Y�� �1�5e991�j��ER.챳$�æ�b�'G�Xm0��D6��>)�DV&�9O&4�d��2_�\��I�����b�i��Z��[�+@<=�t育x��x��7Wh�qa�6Jo�J!
�VY`c����&����8)���O_\���EE�ɔ1��S1
F��V�͚
��|B�[�3c:pSEڂs@��$�?AM朁$`�6-�z�Y�����R���|����L
VI�Bʢ31H��R�I�5�3a��=Pέӌ�$+Q�<�$AΔƸ'���Pg/1��D	����.��2!-M�&�PG�\�p���N�I�hh�3��Z�>y�l�D�\2t��=O�j)�5H��<��D�'G�8���	�d��O6xe�Ӽ3�Na&�ʼ"6lq��i ,y�s.�)cLY�S̖mx��*e
^���[��=( �)�I�z()�O~�HsLя}�,Dh��Q�L���mXc��5���m.4�dp�"�9I�>��f��!?�8���6�ɯn�l����]�Lf$8�T�I�51zR���C�h"�����
T�!�M6w*Xq)E<	�u:�"�;f$�eq��СUR5詟0!��Y�(�e�RV 
���o��(��<D���t�K9U�:����N�\��Y*��uӮx+��H�S�K�#��<9FOLO�t�k�"P��!1�Qo؞LSZp�f5�q���x��t�L݌Y��h�Q�*�Ƚ�O���G��x<�K᭑EH���� }@�����kpx#|:��ǵAX�᤟�3x�Y�rH�M�<A�iT�&��|�$FMk��0���I�<)e�]9X�(� � Jq�8��H�<1��v� �p#��1S[�4��BXF�<��K�v�"Mx� �I 6��3�
B�<��/�<x��q�T�Dfp���UW�<�$)�b�$+硕>K�*q0���n�<!�!#fe��J� o���۶�QS�<	e.�;�zxyWb��W��#�!���pT
��A(�*�+�m�6�!���o��`�C�q�.���M�*_e!����z��֎H����P_!�S�g�d�r���+���c+��<H!�d.�N�y�E܅m�8|c�I��.!��
UO��Pa��N�2uR��-x?!�d�o�0����N��h)c'�*I�!�D�$V�
�9s¸ �BYbŢ0�!�d�\܌!���?�Z}h��*d�!�$ n���SU�	/MUf��Aj�5�!�$�_�X���.M&R���RIB*�!�ܷ>R��J��Z�cOr���!I+!=!��s�0C���7P�!�(F"!���!K��$��@�˶�Y1+�!��~6��y�#S���I��Zb!�D��;�R��@=�\\���-!�dȏ%�
|q�m	$�1 C�UQ�!�$D�7)������΄ [���1T�!�dкgL�0s!fK�P#X�V�_W�!��
eE*5��C%6|������^!�	d~�����$'S�  $C_!�䆭7rn����'LHX�dߺq�!�Ą�L��*�a�HG]
�bG6c�!�dC5<��͒w]u�Bp�!�
&l!�d��W"�����U��<R����&Y!�����ed��ʐ*2�^L!���.G�F���ծ9dJ�:�GW�TE!�d�
y����*[�)�aǑ�9!��NjR���eIZ��2�TW!�֐^Q�d	�pJ���iǿ)b!�D@B"�;G ��ɫ�'�>v�!��J x��C֒GN��M�-�!��/V�͋t�B�1��p�4c�!�=�~u�ċʌ�z؈��1d!���kG�\균��<��Bēs�!�$�) 4 ѷꝯ9�����=mc!�� (�y���#[���
W3�lM�"OT����i�-Y���+R�A4"O����C�x"���D�1:���#"O�����\>tP3���Rl��"O��ˁ��>�����X�L&=�"OD (���R��ܲ�Ϗ4[L��"O���Eܱs�2� X�F��AA�l�<٤��v���mW����ʵj�o�<�e�|n��������r!�n�<9R�
lx�A@R.��u�n�<Y��je�(�H@�,7(�r�H�S�!���$a���a��?A�^� ���7'�!�DQ�B:�ucǛ�3��E����!�Ă�v����&��&#���%���|j!��s;�S��ۦkUT,:�
";+!�4�H�( %3o�	�(�3,!�d��K옠c�
U*�#TJ_+!�d3R庉��%�>N���O�#!�ě�{���J� މ%����dQ4<!�DD�j�~��)�8;��S!��D	|n�<���5>�KP�Q 
!��u���z�J�c��"C�!�D�Z�>����_m�h��Fk�2�!�D)m.0=���M�D:�!�
��!��U����1�F��Ԥ���!��;3`��� ����ώ�!�dM?�	8����@��j���$�!��W�<G��9�-��C&@M1@���!��"�*�� ��9!D��E��$J�!�ę%�"@�c�*w�	rL�K��x�& ��:!P�<��x�gY1d)���Y��)�cś	7�lx5��N��ȓ"�@hJ�oA/*���#w�]�� ,��&��@"�.b"����ٵ�F{�'�~�F�ֽq���g�H/S�:����d�3+)U���[�P���b�k��5�!�dڝU��@Ԝ]>�us�J�0e��{��Ov�-�Պ�j��G���ЁmߧC�J�ȓ8gx����o/��y���.7� ��ȓ.)fM�G�T>�:��/Y�fR��ȓf��!��ɵOs�\�6��6N8�ȓ� �0�Y�gtna��?X�\�ȓ�����<m�|�C��¨2(>���L�f� ��E]
���f�>l���	P����\@q��/�P�F������d0D��ڥfb���a�Er ��+0D�(J�FYK�%��B�V��%��C/�O��VI�����F�hЛ�#@�p��8ܺ�*��kɊe�E ŐY�B���1�B\"&�E'r�2���̑r�H�ȓLd�I��Y�p6�9�T��IşD�?E�D�����M!��\�d�z8qb�t�!�#	�Z�2��]�c��<a�@ N��IC?�	�HA�<;CF�F��丵��;bhT���M�5��&-����`��>15�t땅�Y�<!�F�1#W�Eit!S�=^�qZ*D��Aw`� o��m��P�f��S�N&��<�㯖$�(aŬ��I7�L�IG���O0�*R��n�"��W ��=l�)�'Eʘ���0{Pp'I�j��,��'����
��<�)�h�*
���-�%�ƨ7UT�cT+�4Q!��#7.���oH8	:<�Q���PJ!�$�5I�t�8�"ڀִع�.F8X+!�� �e��γOf���1g�(+�<5`"Oz=x�'��3�����6*�l�W"Oz��"��YǦޑ3଀w�O,��d�7#�t)�BG�%W��Q��e�!��T8W"�,z��r�����%�0C�	WQU{3L�Oܒ�2��ת,�C�I��H��A��@gP��@׶DE:B�I�3]��w
��m"Ƣ�^`�O�����' k��"�Q�x��Jv�٢^!���Or�gB8K����cԝ0�1�D"OưRd�
I��U���˼^|�j�Ig~R�i�����BA@n<�E�F�Q�lC�I�����Ć+	P�����
0��B�I4$��HPK$&8ܸ���X7VB�	Q�d���e��\���M�b���=�Ó}��+����/Ƅ1'ʅ.��1��f �9�lK�|�6uK����6��,�ID�����4ӡ�!;��(�tǺ@�t�Z�"D�$U��Z����h�8��8w�2��hO��I�$���*.�{�f�ڥB�}��C�ɏ�Ih�l�8nD�p�q#f��#=	�T�������^����gg�Z��ȓy}�A����w.�1[��������?��iK�M�t��u�<dK@
4D�0��g0xhQ9�+��j��B�f2D��SvFR� � 41��s@A+��hO�S= 4�|K���2�.���>d�4C�ɢ.�d�[B��U�B�Q>@XG{��9O��A��B4@�Ւ�/�&����"OZ��QJU9
ǖ �$�����"O��P$K��E��h	�g�>�4QR"O�a�hC�-��AU�H�d��6"O\=�X�BVNm#��3@�H�"Od	��,a�r}��%�'8 ��1"O"5�D#Cx���D�*#�BYg"O�!�7���H�| B���4���F"O&�2L��6LY��AG�O�j� �"O� �@�\u90"�[)d�b�\�8͓��'&Q��' 2
���@�n�rT���7D��*R	�4~)`�c:9IT�"�7D���DJ(�����ˢ*� Hb�h1⓳��8W�Ւ �\m��d\�`�h��"OH���ޤy�N1:c�I��qu"O�P�H)=��c��ߒA���sd"OdeԯUh|�4'�m�h��U�����t�d�Q����t�A�n3#�C�I�y�h����"��q�b^����O£=�}�㠆d�@�*�CU�R�AL
H�<�g���t��q�e���� 0"WL�<���<V���ի�-K�(��w�AG�<�Pgn�^��tƐ}�Yؒ�EB�<����W�Fy,��"�����m�f�<yaO>G���DݞO/h&�y�<!ǈ��L�a�o��:X�YGRu�<�6hC��U�� y{��A� �e�<��B 9P���
�(����тy�'Nay2,�{�0����ȬLu���"C�>�yr.�r��!�fH'O� �O�&L���ę?�"��`��k:er�mA�j��z��ė/d���8���2R[~]���J�ay"�	$js ����^���q��>C�	9?{����'D��z�A�ۈ^eC�	�<�5C������҆��cLB��;v�`�"�3>ډ�*f~C�)� l�P��-�8a�&nP�GB6$���VsH<y#)\V��ɰ	m�!�� Ii��X�?�ųjDQ�F���B�IWD�4�!��l�N�%F]�.9�$I8M0!�Ӑ0�d� Q@K�>�93(Ӫ9!������ ֣4���)/�!���
�v����ƫ�H��e�H77�!�dK�I�``����XaɦӧVs!�dO�.�j�ZD�$u�4}�D�=�!�$̝cY����)K�8�rS��%d�!�-&���d���8�L�
~7!�d@�(��"�L��(�J!�$�?Z1��b��Xg�>����3�!�DL#BL6R�!y�����<���9O����^�Vp��AamȺ*٠X�"O*t���`$�={�,������"O��8LN+Wf����%��P�"O�ز�h�q4�*𭗧!Ӗ=��"O6�Pס�!9�-[����/��H�"O\�	�
��.�@Y���1B=��`"ON4�&A2{�^\p�@	 6T��0"OU8Ǧ��B���#��`,�t"O�}{͌�SL�p�m],�|�"O҉�W�C��!�9�.��"O�y��͍(�A�ạx��ar"O9�ǜv;0Ih"!�_46u(A"O�d�E��:�D�C��)iD"O�a`4�T9�����N�.lJ,��"O��8��K�<���T)Vd"O�a[�`�9s�6P���s�j r�"O�b��zK��!ĬQ�A�d�"O�ZP�^�|�nR�)�,c���d"OD�C��E��H��G�&w<-�"O��:r�W9�,T�Z�Oqz���"On���ȞYFx[P��+n�Zs"Ob�� f%K �5˖�U |?<h!�"OzyʗH��d_6%��,,^݀S"Ot
7jj'�U����G8��ˠ"O��P91������.��=�v"O.��F,�f�<pb��"6�ذ�B"O ��qiƢp0�)֮�5SJZ�xu"O���q��mm(������.����C"O҄�r+@�B?�1Y���:v��t�'"O�a1��'�\(I��	�N<h�ad"Ox؀� �!_j�+��Ǚ%ܱ�r"O^Qr�jĠ,hΉKD!�#Vf(�"O�� ���\�`��9K
��B�"O�ꢌ�)��l"g��"� �`�"O��RFѧRu>��AΞ"��4"O�1��Q<^���ʉ9"F�!c"O2YC���?Ӏ����W�PS"O���,*���!�͝'��W"Olb�	m��+G�;w<�a�"O�u;ү�(�x�w��Ua�D��"O�PCOH�d���XeB#6Gnȋ�"O���G��Qi�9X�!��j.p�!�"O�Ujq(��\9��a�<ЀB�"Op�@Ů�<B?8��0ӵN�r"O2 ��͋�L0�I�B�~�"O��H�F��@u�F8]����"O�)Cu�֥A�q�O�iO��D"O�a!5��#}Ѿ��5eKD8��S�"O�P0�H�%0vx0V��=D0���"OfX�fa&G`�`��
�B"O� P�SS��7L͸�����b[��J�"O�4	V��29#j�1O�,%Y���"Ol�k抟J.:0�v��m����"Oj-�-O���ja��Jb���"O���b[�Y�<�FgS�#V��	�"Oȱ8�A�-`B%E�5S��z�"O�|�����2��F��EPl��a"O�Qϊ_a��H�+J-e:��J�"O��sNV,<��2��*\��G"O��r&��#�t-1RI��pf@�"O��re��%���:�A@�r��)�D"Op<X���q��@���޸L���n"D����G_<N���
g��D��m�r0D�����	"���P�T�4lr��&�+D��Z�j�*nV�(5��;4t���>D�����ag�i�K�>U�<���:D��q��Ci�
!v���
�"-��4D� Q#��#��"���6z	4%3 �-D�$c��W'?�H���@ ��Kw-D�L�C\(b�`��,Իj��PYWA0D�ਓD2��eJ0"T��82�1D���$�("�"�����,jj�G�/D����%��@R��2�6��0D��H���&I~%� A`�X�� /D���Q�H�n�2����_X ����0D����V�g�!2h��]B�0��0D��hڴ9����@��N٢\�F%/D�(�Dhh<�� ���_td��@+D�0`c�6x� �����+�~$ �n6D���R�T�,����� `=����b8D��(���%��5���'g�\u�3#8D��QD"̏(��A*ЭR)I2<��5D��h���)f	����Sb�4t#-D�h�B�3yo���sѺ�и�/D��0�Xt7b}�(P#LF���E;D�$����O<�U͛7.�(��$D����(� o�ԥk��b'���A�"D��.����Qx�i6�Ј�i&D�A��R=H��٥ ��n�Y�h?D�<�0&�M��E�P	l���r��/D��s�$�5�<]f��v*����+D���t��
Sˤ%�p���<,I�+D��*��"���Vːu��逋+D��g	%'�講�$ʺ`��$-D�\�'ߘ>�D�ơ�ޚ<�ҏ=D��X�
ܲ~5����p�6��:D���t��Q��%{�"��c��� 6D���`F�,tD�` �5!)��I�I9D�p��)0�A���k�M(��;D�$;1ǉ3w�P��rVR����$&D�H��Ί�G�^���?Ų�r�J%D��a�нM4��I����鐤�(D��8���<�㢄V ����*D�XB��U�j-����6_�N1�6D��R�К�����̔� 8�h�C'D����ZN!3P�N%Dh��j%D�����Δ>j�!�3t���=D�ܺ�iW�;����1�E@��Z"�8D�����,V9�يD��>50bO3D�x�Bɐ�?��L�c΂t�����<D�Hj7ol�"]�ui��+'f4�w�?D��%�Կj�ԴQ�%�0xC`�k$a"D�Lj#*�jT�cb��)s�^��S�$D�$�(�h ȝ�`��4lU�-D�� ��"o:��a�ԉ��,\"�*�"O��	B�I=-R-	7��(>~� "O���@� 0�L��V���C'
�Ap"O��! �Xjp,�r�]��c3"O�i�b��Pܕ�p�
�S���"O�d{D(U?vE���̏% �Hę�"Oڭ
��>�z��� \�\�����"O��a�F�]��OЗX��ĨU"O �Ac��&�P��+ΧrF��"OxQ��F�|�j�8f+*z^�d�R"O��� cR5&8NiS�I5<A�8��"O�pJ����1�l�Sc�ХhB�Xs"O�i���!Y�4eTE��'(*i�"Oj1�k�6�x�C��,<�A; "O��*4Eʭ<�ix��_Bb��"O�(���N�l��a-p�jQS"Oԑ�����cD��he�ؖU0��"O*t���?��p�s��'���"O.E�����A%��!�@W��]�&"O�hK�M�,��[U/�T�Be�$"O����GP���SÇڜ�*0�B"O@�ad�S\2��d_')�ԀIp"O�#̋�1P�!s�M$�4�"OP���	_.S��C7 ݮV� �r"O��֡PMw�񂶏�;����"O��-ʉ@�6%����*� �"On݂W�F#[��YC�M�~�l-"O�i��`��I����G�#�0���"O2��n��>�$�Q�E��,��"O|Y����#S��!K��m�xp�"O�HV��r�U�0DV�qy�qPc"O}
&똈t�b	��W�b-ʄ"O �Y��Y�pc�Р��|����"O�I`�퐍�"����>c�|�"O��S�٤t,�����B���"O�H�B!]�Cu�m*.T#
F���"O��;en�:"H�yQnU�LP�S"O�}�W� wE�Y�g�YHl �"Ojb� $th;�e޽|L�y�"OL�M �G��1�L%� ���"Ot�0��]+6�4�@��X$"Ob�*"��"�(�R�P7]#�9
�"O���Ԋb��)+�5Q���e"O���⧊�*S���D%�gd!�v"Op�+�޶
X��C$�F�ʀ"O𐠠�O0P�Ӕ�	�v��"O<5��Q�<��3q�Y_�Hx��"O �(��2�Xq��_�hr��"O���'���N&T|��e�{jnIaS"O.�1 ��#��Ī���e��("O��)G�E�sl5A�M���"S"O�x�� ���R̃�9�,l[�"OB}��)P�d�|�`B��'G��1�"OT�Z`LH�G10ey�j�h5 ��"O� )�H�.W����+F�c$���"O�$�F�4��<1�`����8xr"Oe�H�(�D�t�R�v��m�b"OHű&OYl��Y��@s�"OJ�q�BaE��[�&�]�нЄ"O^�`��
�t )E��$�bq��"O��{$��"4���A.��%�b��"O��r&�0&�MIP�-}T���u"O ��Y�o��k�!Wx��"O<�C�-a<0�T`ϧE��h7"O� |E��ɀ�Wbx�/��~Ҩ!�"O�`B�#��"�T#%�i�s"O��� ��<w|,�D��o��d"O�x1P��Q �JQmY�;���$"O4�B����b���iC�#�2�	'"O@c��!�`U��i^�,Q����"O�AZ�%�3m����5u4�ɀ�"OR����N&Ʊ��_!Wx�(ӷ"O�}(����dBpbfۭY?���2"O��NۨH�,q����FS*x˄"O �9��ֲ]f�$ꝇ-�t0q""Ot̒5�Ѧ:F,p�6�/�h�ڕ"O���Fh@*�^0��G�+O�:�Ѡ"O�D�E�w���iP�1@����"O���' �@*|;g?eDU�a"O�tJ�e�^2�A��I�WU
ͨb"O<[�) �1�44y�H<F�"5"O�P�2��	lW��B
 �1�t1"O�§�P2Xμȱ�8���r�"O"y�tGI�\�ji����Z�r�"O�ah&肜n�V��B�&���hP"O�a
B�]�#�V0�KJ}��-�3"O�!����"�`b�@�FK0�!e"O���R�ʖ9Z}�wr���s"O�%��h��JzR��E�В�DPS'"O�鐂�T�Md�3�(Ѷ,K�� "O�E#�U�M;,��Da*t+l��U"OB��E�߭@B�)a*թI��"O�ճ��F�Q㤼r�g�!y
�ir"O<x�`AjJy;Q ;�����"OvH�gI+��K��|�0�r�"O�Yq��'�x8���o�x�"Ox�CA"��X�9âAM<E�l�"O���dN��PRqaH�3�Q��"O��re�6~���9��31ؔ�1"O2R���9W�,@��/y���A"O�肅i��j��D�H"&�RUk "O
�1��߭j����� ��}�"O9*'�л`�x��H<貵��"O",H7
�=|^���)�ܬ`!"OtUsQJ>i~�<�P�-o�0���"O��قO��&5�bɩ��p"OVYv���.�X��ЏJ��)9%"O@�"#DG(���b.�v��8aS"O��j/���Z�M	&(>l��"ON��8'P1�
?Pn%��"O�Iq�Rlƌ`3U��)w�z��s"O�A��d_?{m`�b�+@��!�"OP�Ѥ	���y�g ��Y�"O�pp���F�t�%�0<�u��"O�=�i7D�,��gH[6E ı;�"O4���ٌ7`��NV�s�"Od�i6���Ң�xŬ�!���"O����H�a?�(��mħ��`��"O��P�M5RL�p�&�n<Z�"O���ȅEA��SfПG��Eja"O��"d@�\j*,�b����T"OfủEX'c����+q�0�g"O�}�%E�.O4
��<:�4�B�"OHi���9Z�Q Q�bx 9)�"O�!8t�;Z�>��O��* �"Op9�)N�e�x�  �̨f���#"O̅R���"O���ʲl	��P���"O
��!��0:@��ʢ�O�f���"O� &4�ਟ��Řw菗@� �b"O��W��>19��(1��>�=A@"O��gn�av�����;6�Z�"O C�L��U�.��o�"@ |�Q"O2�iQi��k5�E��`V4C��"�"O�)��#� �	�e .���%*O\x�"�޷J�̄� AD!a����'i�eA�N��2#�I8Ѝ&%"	a�'�TԘ3!-hHBǥ���L� �'V��`ڸ�8�A7�< ��8�
�'j��C��
L-�f�Ս&H���'�N��gIP<��M"'��:l�^I�
�'�ͨ1
��Y�b��рL�yʼ�0�'(��$�J.>x�Q`図����'��H�#I�;}�&m	��*��'b(��T�w>��/�@be�<�yb���,���A��N668����yR˅_��mP��E��r��y2�B�,�д���Ϫ��(�N��yB��';�RdZ�-֢z��$/X�y����@Lr�	Xj\�� ���yr���n��b�㏥M���cs����y�!7Y�X�`�$>�v�3��y�"_�0���:���0/,�x�B,�-�y�.��c�R��*�,����BFM7�y�鍑<M�L�d
 %���k��y�)��^O||HV^�G �	1�ҙ�y�a@*&Ϯ��.8f�ө��y"دo�*�$׌P��j���y¡@�=ڶ�9��O��|�"�%G�yR̵K��1	`J�7�F!@$&�y��Z�&\蠇�5~PD����y"���F%	T C�uʠ$���ķ�yZYy��l�D�ҝ���A�UR�B�I�3>�cSR�+���Ò�ɸu6nB䉑�f���(L6g����0TwjB�ɨ6�NAQ̉�^'H�{u�`�:B�ɇ"j����7}lj�uHK�4(B�Iy�xA��8�r��D��NB�ɨ]�P]���X1���M@B�IKi~y9&�
˺��ƆKB�	�d��̛�͜d��\�5�ڻp��C�	���q�m�9E��{b�B�[��C�I& ��!q%]*�@ �@/D�C�I5vV~ ��g�0�;�k-~|�C�	�Pz����;�mY�ᛷ[�@C��g�zQX���Re�A������C�ɬ��E �� r��y� ���C䉢-��Q��S6W������ÔfdB�	�sk�� u��i���#DA�F>vB��cW����J������n�"C�ɟ6xT�:�l�{ݤ�[���N��C�ɸ>��jC_�s�X@Cbd�.j]�C�I6\��i�I�cd"�S5��0<�C��=/*	�g���jS�˱_�C䉩mx�0 ���B��P(D`�pB�Ɇy����a�3a(TP�v��#�DB䉁g�<�!4�ή-*&TT*Z�B�ɠ��P�$��V�ը�R5�B�I]{n�U��x�:M"�hQ�;�~B䉶�p�"BDGN&�A��/=Q�B�+�� ���E<������"�B��8��hfI�&`�\���/��B�I��P��K�l��l�6���mC�)� �-���:P�ղ�+V��s�"O��83���,�1PǍ߾
��
p"O����F�Zj�dҋ΃�:��"O�aK�M� �Y�����T�fDs1"O�H�GK�P��䮐+2�@p�2"O4��r#�1$ P2-�3]���3"O>����nP�ԛqJ�"���"O�A�P� ?Ν8!$U�B����0"O��+�O0W2��{Ƭ�	��%"O���LȿTL���Ga�r��"O��&aW���-t	�>`�N5ɀ"O����
Z�_}"�+YR�dh�CJ��yR��e(�Ԛ��A� �ؕ.�yh�kXXHHA��~X��(���/�yb`ψ�"��!f�+r|�I�(W�y�#���(�.A e�He2��T�y��Y�rE�� vE��\�䐊�O��y�L�)N���Q&LP� �^m��-8�yҮS�z����f�*�8`�@���yb� ������ς��Z��X��y�#ړ5�
�� �]�jb����B�yr��#L�*X�V�E:[�t�7Ć��y�$J�8t�M����$G84�v�Y��y���]�����"%|Q �#ڝ�y����4�E] p��-p�H���yr�KPFh�J�@�B黶AӐ�y���R���c�
���d-Ʃ�ybȜ�t�,�R��f��L��y��E�p��M�/4��W��:�y�������q��y&%0B�R�y"�]�3����W���V���H��y��-	��sE@� �&S�ɗ�y���?zе�խ�6$gh�A�$�yL�3�* #ρ�.��C 8�y�`�Q�q�	&T��P�c�ʗ�y¦>~�UH�c��FBH�©��y"HU$x�v���/�?�� S��^��yR��D � J�6O�!����yl�#�������MN�����y�*��I�9R'�OI��Q��4�y�&iZ7���Au�|r�ٴ�yr4��X*e떈:vz<Rō�%�y2`� 2�;�IՁ9-�)���y��ĴQ����%�_*8h�]��ȣ�yr��&q��K1f��4^�u+�H��y��LB@��p��9()vQC�쉨�y2��m���҃�8���#���y��>p�>x��ʖsP�2��O��yR(Q�W�����_�q��0�VIȁ�yK^�:�V(Avo�=v_�X���ɣ�yҀ��{]�# ��q� �1�Ȋ�y����7B���'^t�2�ju��yR͞�@�r��ѪȢo��	H5�¹�y�M3�Fl�q͑�S0Н�����y���*��ERA�ָ!�&P����yB$��i�����F�e6��k��y�KF�]Nz�8CL�Z�L�ă��y����v ��D"Y�(B�GT�H��'7�Ðc?�l%14��W�pQ�'�^9�!��I�ȡbd��G TYH�'~a�7!��(oZ�$�G"@m�'�T��@3:¼4���0��IH�y�嗗Dh��	�ʩ ~��B���yA�7p�U{����˷c��y
� �h+���1��mj�8"�T�K�"O�93r��9:�23s�E�F�A�"O�\Z���g���p�U�%$P�'"OX�!#��xw~�B�D	�Z�*ڂ"O�'�O8t��2� �>a�b0�U"O
�y X�@("��Q��"f��"Op��b+�j�>8�C��u� Qpr"Of�3͉�L�P `�l��{iLZ7"O$p���ʗ(G���d��7C\J�"O�X���X��HQ �?U��Ö"O6D�cI�2.�,QeN�H8��)�"O������^�xe�f
�89R�"Od=��Շ�Hy�aE I�q��"O䭒
�8i)�Dz�	�5���:�"O��q �#]>�q�C�2uQ�(�F"O�1�����I��1�GܯD!,l��"O4��� :�<�8�L�"L���U"O��"%�ƻ<|�a�m�\�t*�"O�	���e聡flG�#���"OH��n�'9T�j5��#8: �"OF2W�קe���&͏F$]�@"O\ݘRˍ7%`����b��~hC�"Ob���7G7FS��D�o�♻�"O44�L���Azt�G,���;�"OV9"�z��E��A�����"O|��a-:ҵ��L�:p��}sp"OȼѶO��nRDmX2��W�����"O�*�Y �E��j�5�p�z�"Otk�	b����	>Np^<��"Oy���#Jv��o�4wMp�	%"OD�3*M�Z��h$K%SK<���"O�lIg�RT�:E2�-�;r��"O�����DVpx���5o塖"O�`[T��+Pe@��!j[�`ؠ"O������7q4��3����\aT"O�e����P����p��3 ��s"On3u�A�"TZ6C�7�B��"Ojm*3�C!B�z	!�61v\�1�"O�$��m��mZ�!2��P��N�i$"O��$Y�s,vL��&��qb�"O��ca��}�"� f)��a�"O�p`E����:��2���A�"O
 ��FY>I�Up��m�Xt��"O6Uȶ��5P�,�@��;���ʂ"OFlV&	���؃����6p�q"Oz<�%`J�
`�;A��lހ:"O<}h���,mg��B��^>S�Z��"O�A����'{(�Ac��)k�,8)�"Olt�/��m�8�b�*�~	R"O�@鶃�:�P�F�ίY���8�"OI���5�4xb��@I8��F"O�A3�!Nb8�'�R3�h "O�`�Ο�q�h�C`�0,���"Oҁxh}�:����7)"��"O�}��L �.�S��W�w䌩$"O}yv�� R`P�(���F"O:��Ǉ�yv�@�M�(�ȑ6"O�z��Ͻ)�ȅJ"��|?j��"Ob���ƨ�`���<f�ܪ�"O�2�b�4#�>!{�!>J|�X��"O��!U��0^�E3��z��;5"O�PN�R�*qQF&�n}���"O���f�Wےt�b�O�w�� ��"O��*Dh�@�Ѕ�!ǖ,�(���"O� � �&H�r���9t��8�2`p�"O��y��ؘ.A�h����рj�"O氹��e�H@뛪�X�J�"O�-��c�!D1X�
;n�~=Ї"O^�i�G[�z��{�bA��	�"O�I��'/��U�S�x��h��"O���eL�)I�H;s��'@��"OLц��RD���!�0@U��"O�xs4��
U"��@�'Z-ֵ�"O�]� Iy&�B���h���p"O�@�3`ρ8������3W���C�"O���ԠD-m�|��0i&3{�;�"O$B2 �-k�b0v掯:��"OD(Ӥ�=c:(�y�D�bje��"O�DS ��7u����%�Jֶ�6"O��p6M�#Pp-*�E'�N���ymт6��
���#ވ���֩�y� �"U�wʑ�".~�(妇�yB��=F����.�-"�tr��&�y�)��̎Y�Pċ��d���y򂏚t��)��Q8�]��B�ɦ<g�qrT��PFL:�T;�C�I�'�>"a��j���`�����C�	c���s���.�2�H>��C�I@Ԃ��2EYSW������E��C�Ɂf��\��K�)5����H�,�B�ID*�9ÃD5xf����k�,r�C�6'l�(�k�?GK��2�����B���D!�
��b����00�C�	� ��1���Q�� �]�/�B�I�!'����R��I��l:vB䉥L���Z�M/�%R�\�TLB�2;�0��^-涴Q�T�n�B䉹s|��bO���zr�͞ �LB��<�$����M:i�n��'�
YB�	�8o|����A^JD9$��7��C䉩sў*��]0.p{�^�J��B�I62ݨ���bI�/�Z,3� �:c� C��!��$�a��,l�
�F>K��B�I&	{��u#!cH�UAC�N�D݊C�I�j�ޥ��d]�O�Ρ��Gڽ:��C��6C�^Ĺ����f�bR��;\RB�ɪK�@)U�N7�B!�/w$B䉮&�l�Y0�G�X6�|�PR2B��C��*,��@�
�FVi�[��C�I���-#�� M�r��L��P%�C�6+<��E� �x�Aۀ��C�	���hV皡y�����ܜB�C�I"����w�F$����[ m�NC�4kA�Hzq�!Fi�@�-�� C䉞|#NhR����މQ�3lZC�ɘ���Ȱ�� pl "�UN'C�I5Z3F ��+�*Z�3G�	lR�C�I/F����w㋥�.�����}L0C��4Ъ���>i���	���+�0C�	t:$  �ڵ��b�ٖe��B�Is�0��V3Y�|�i`�	�<2�B䉓U3Ȁ��OԳF|: ��i��#�tB䉀򾅱��������҆C�~{����5)I$Pj�〘�B��]�X�pȆ�F␃v꘏H��B�(B��m �,��XA�.?�B�4%v
�(��W*��|
`�	% ^zB�.7���
��>e�r����ۖ.�JB�)� ~A��+ɮ<B�Iց�4����g"O���u���Ӑ Сk�z�0���"O�ib�ɝA��d�E��:��q"%"O��@ϔ8#x!`�)A���d��"O�Ej�b�^/��v��(�d���"O�xB�ն"7�� '�΋hCh�Y�"Oc�Y�R�@��錙Y��s5"O��q4�Ę ��=a,��H��"O�L{� �d`l�
v��3$�B���"O� �E3��}#�P9?����"O�(��^?V\����z���"OB��,���h�ӯJ�^�!V"OTD�PE�@�fi�+Ĥ+���j�"O���g��#��02��)#�D�"Op�@J�L�<�JE' (Ҿ�q�'1O.��"�F#Z�R0�W_r�� +q"ORE��n�2b\��D�,Aې��"Oƭx��5d�������ؾ��"O���pb	;'{�<Sc��Q�Y�"Oh<Z�"΀��� Oy�4��"O�}���;F���/�'!�� �"OV5:��q����e�w;��j"O�l�gv���ȹ���"ON��%�Ì"��iju���f��9�'�pq��.Td���L�m�l�{�'���S�eY-g��tb������m�<yǬ]�~����3��13sG�A�<�Z=K��X 4C�,�f�j#�H|�<���A�2C"�S���>��}bl�}�<9�&�3o������ =���_�<�W���$�*qG*+*Q[ĥB�<9Ǥ��!ۈ�:Q̋�Z��dpf��H�<��+"�s���7�0��bF]�<�&Ě�Pu�K�&z��{���X�<TV�����`-�I�qK�*�I�<1���_�J��'�+!}H�z�%�J�<%@��>A��KN�$��b�%�F�<���\�T���(�(DvR&Ǜn�<Q�ƶ7B�Lۃ�&��dQ��v�<A1���2y�q��<�u�Cs�<ɴN�r[�H wǓ�.������W�<�CǙ[ ��e��G���`��BU�<�\#Yʆ�c�G�-�ɢ�P{�<�0�	+]�/�>A_�eJ���l�<���^�̙w��>ZF�4���l�<IЧߛD�\)ڒ�P�R �TE�i�<�ᬊ�%�f`�$E�.+Ae�i�<�@.� q=�IB�^�D���E]�<�U� �!��8a��4+�`t�&�Z�<�휕eVzL+��O.��&B�<�b��"Q��ՓW�P�����@c�<�t���+8�!Q/��R� ]��<T�L���Y?,0��@��U�>�`���.D���4M�7/�1�4k�=SHA2%8D�X��j�� �J�HU�dO"���,1D�f̅�.�9*�$/	�p��i.D��� �'5#��{�C�8V���',D�|p�`�njd�[�̂ ک�!�-D��j�=��QWO�8G��9P�*D�h�1o
�l����Cy�ԓv�:D����Mےu����#���b��s�7D��Y`V�0�4C�� >�y�W7D��VO��4���@��<ؗn ��R���S5l���6�I�1�1���I|B�)� �m��&��r��d��+i
����"O9"C�U0<�����Y:��"O�(��G+� �窊7�M "O�-��+�f���cS*�1i�(��"OF��R�@,z�)i1Ď�/��x��"O�qvꉂk)6��A��^�|I��"O�Lx��M�U�� Ǝ96� ф"Ox ��4l��!� ��7&<�""O��e%ʴ~=�|��/��M�,��"O>���A�vq1#L®y@�{�"O�xX���)W̠A3��Ҿ*m�h��"O�:ca��Yr�Ve���"OV������#�*ً ���iU"O�pxt���-�f�({��!"OH�P�}K
���ē'���"OD�P�B �}~ � ��/^����"O4ARb�# �d�T��+fJ�Q1�"O�!�:i�A�׃��N 8[�"O�Q&E�%!��UÂ�7e�0�'"O�Ș�	6�4��;S�ty�"OL�Ap G�j����A�P���1�"O��F
[�X�b�B낪��$��"O*)���&P:�"���bx"�Q""O�(�/?N�8a�i�cj&�
�"O8�Ȁګiͺ�q0�݂0OLH� "O�,3�I$3-깑CG�
\/����"O"��Y�ZT����s~U��P���	C���Oh�yjG�G�hxHP��*ɑ���3�'tՑR�^�{k����Ɓog������ѡ/Z4E1$�>3fh ��Y5�y�!sB��큉? ٧�yr�AP�d�0�S10�0ˠFұ�y��0�Z���l݊-J�s���y�%�>l�Dx��:l�$�B,��?���?�H>�+O1����@ ^T��`�ʼ6.<��J-D�4���ZZ)h�a	+�`�U?D���l-�$����~W~�ʗ);D�x��Y�kQ]y0�����D%D�4����/{�|-���C&������7D���o��Y�N�iB��d�2 � D�c�!L4#-z�R����$�:V�O���)�ID�O6��3	RtP¨�5܆1��"OƔ5l�$�0�C"��_eQ"O@��3`�&w�"!!�Ǳ1W� P�"O�1���շ|����q9
 "Or� `��i���b3!ЄJ�Z51Q"O��# /e�<����W��
PO�P����"E��n�$�"�` &�<)����(���
��ā}�@��N]�Qg�<��"O�3S�:~�ي�c[[E*tp"Oj�(d��d�~���C ����:"O��J�ώ~٢�C�Aܘpb�`�"Oz���hL�����jS�Ţ	�'���b�Yg�z�k���1�괪�'T�ti ��8i�v� ��S $���-OJ���<����O�9�v�\�2�ءX'(�2`f"OJ9s� �9|��(��'Y8%p1j�"O0P�3�'��H�DǺ�ba"O�E*ǩ�)�d�	 �/W�
���"O� �PJ� 5�R�y"�'A�T(��	Nyb�'
1���Pt(_3� %@�Ly��F�' ��'�=ڦ�[N���G�>K�VE/������E{R�$�%u� J��N��,ˌ]�!�8e�hX�O�5��;l�!�� �41���%��ф
� κ\��"O�8�%� ���i�>L�P�y�"O���5��5��|���<8q�I�5"OX�i� P�Y����+UlP�$a`"Ozu��1��AJͲ @X��g"OR�J��@ �x��񨐒L����"Op�RQA�Z���rM��W�0�`"O
�F�[#%>��"�B�Rz&8�"O6y�d6UF�VQ,q�୹A b�<A׊R�bt0��֨".��7(�s�<qP�H%;b9�ᛦ7~HCe�th<Q�ȁyZ.I���V��>H����?����>��-`R��-�nx8'f� 1T����b�B�-�2�� a��?j����\܈�d̝3LH�+k=s����ȓw��4F�%-p��Ӗԍ"i��bZ*	K��ޱ��K2�ϋ{�2%�ȓ'Ѣ�DD�[&2�**��u���d~���w(� Ӓ#t	a�j��?y���?y-O4��$�`��8hJA�O�ޡ���>&!�$?w~�����S�b[%e[8h�!��ٌMj��%�ƘP�4UÔ�Y9a�!�$�p�tA�A)�9J�VT4��6T�!��`�S�]�P��43"��s�!򤜭����dOm�Es�C?�'�a|RÒ�~�����;���j�
�8�yR�6W`��a�W�0[`�C&��y��:Z�|���$�NTZ�gE�yR����4�&@�O�Н�'�y����}���Rwh�1Ī��	���y�T|5���E�(�V@ェ����x���)BȚ�y�ւ&jj��!0��	X��`�B
�-v����#6�H��/D����ʞ["�`SSI��:� D���&��)��xSC�ǉ'C(�ԩ=D�H�Qm�,��eO�@)�A*�=D�t��N\"�ru� %"��ŉ��?D�<��f�/��D���:>�^��g� D��֥=`�j�	��K�P�� Q�OL�$>�O^ܻ%��#Y�q�C�O�#�=�B"O ���8$���,Nq?J��U"O8�ɇBO�S��bG�՞%T�
'"O��+@	�5l�r<�J��baN��7"Oԝ夗?i�$-�bJ�0��}�"O��f�߂:Nh�YJU�ʉbO �����=YŘ���ɟP�$�d��O��d1�O.!�a��45�<�2���Fv\aCQ�|��'�A� ��.�t�3��&9t�8�	�'@a2�*N���0�F�/Y$;	�'�P�Ռ�:OD��C*`���'��qT�)�@{��j2�iP�'���Zc.�h���@Ǆ^g;�'kʄ�0;$߂��w�j�Bx��'֑�ܒ.8� ��W�jQ
u��'�F��%��n`bi���<e��'J�#�#�?�BT�[�{nd��'�܁oH~�������vθ���'�<xQ"�l4�ȃak_�b��m�
�'M<�x�(ޒF�dtZDDR�Y��J	�'�8Q��Dj��Æ˙M�Fe��'�
��IϬ|�PMJs 
A��z�'fLHdAO�?�����>����'���1'Oҏ&R��á!Ϊ2����
�'ծ����9���¡�) �jHZ
��� �����XU��x�Ò��4�{V"O�iӶ���I�r�������E"O ��#���T36@B�One	�"O��q��À>����UN^ d�(�"O�4HrHC i*��G@$0��S�"Op���-�^<�ˡL9>րE1t"O�I�H2�0'IF�+�x��t"O���i��/��(P�(߁%)�xЃ"O8 �c��'<��5��� �M�V"O�P�1�1޼�sяY���i��"O����0Kjа#3�Ɋ�ڀ��"O�Y"��X�.���a q�� �y���צ��r�?j����3��y2^Y���Q�Z�e�Q#�-�y��3$���ش�T
Y�ra��c�)�yBE�n��U+���I���1/�!�y�L�#� 8b��1B�p��Fِ�y���$� �i��^�,�� ����<�yr�">�L���\�VhA['�ĳ�y�gϰw�hI*r�ǬUd:�ӪL��y� ��/F��a�
pz(2�ɹ�y�cU:]*�	S�� "x�Fe���y��=?�ث��˧i����ъ���y"BX�`������R���y�*�
�y�'U q[>���4g�Hb%����y�	�2TQ��R�B��uz�(%E���y �l��x�	('4��d7�y2\�C!����}��%/�yo��1�b q��1��y����yBMҼ)���hč]�$d��a
�y.�0�d��m��M�!l@$�!�$���h�8fgJ'q�H���K�
�!�$������O�J ����}!�Εh�� �8<)D�b(��
!�d��r���D�"�pp�'�!��*7N�k����/�\�!�6Gila�TK"z�xp$E�f�!��Y�\�th�e�8�y��@�wl���آ5)АpS�Ws��ӱi���y2G u��uS���k��Z�EN�yrh�9j.���\�:����s���y�
�h���t��>h��H˳�ɠ�y҄�k�X��r�ִUQ���BS�y�����*=� %x���0'��ybn��pd�\�T�v,,Tc0�"�y�䍬5��X�P��u�<tA�N�)�y2A
yN.��Hٱn�����y��k���ĉ6>��, �����y�k;G��̋��5�&|
��3�y҉�ppR�2ǌ 5P�rB��y��3S�Z�ZTF[-rB��!�C��y�̆Y��Q�`B�ѐ�,�y���$Bʮ�h���u��.���yG��_8�'�ĭ�@�8���y�(RL��X�tb@��I!��y� |5���a��T�:��ԯ���y2뛕1b,����Eġ��W��yB��_��H���
Z'"���yb��u�tX�e�[�	�Ө_��y�aʺ��Y�T ݓy�V4����4�yB�
$I[bP�$.�#kZԝ�s�P�y��ʔQ"2�@����67�	��.�y��-���̏�9��	T��y2Gƅh��E���0XFM�R�3�y
� Z���/�z^�j7�V�@�`��"O�p�ҍ<�h����t_�DY"O^� 7�� 8j �f�
�zL��`�"O.@�UeES�v\B��7YHj�
�"O���V��z�ٛ�O6?�U0"Op���-�6XBb��.,3ꐰt"O���EE�>�ޕ���.�#"O E��̔�
�8�k��!��}�"O�mذ ��W�	F	�5]�L�2F"O|�F�/3dA�ņТQ���5"O&e#'�:y�	K@#8F�(��C"O6y�b�T�Vu��!زd��k�"Oʘ�W��)nŮm����c�8���"O��[�%�Fin͓S�9NfTS6"O���1m9�Fm�R�u$JTk"O�K%--������B/K}�-�0"O@�
sd@+B�<��,�Pec�"O��xb�210kױCGVY��"O���eDRo�n�`��B8-����"O�d��㚗?~��kS#�&;��X�w"O6�����.?���! (���:�"O$��`�G��%h� ��t�l\`"OT�ٷ/��Qg"�ɑ%�>C���3t"O��q!٫r�xY�CP�`"O����D/����$)��H���"O����6��u�ՇC�D�Z���"O
	��%Ï�p2"F�0�&�`�"O`%�v��\�8��$L'L���Q3"O�@�JBX��Б"��4VFP) �"O��۲��=�͂!���T&R�� "Ot���#V%@�6�� �ۃf'X=ȅ"O�5�^9K���.I:I���B�"O�� ��;x�u1�M��dC "Oj`��@�;~�y�F3C�*���"O򭣄�A�q���ñ+��C��� �"O ���T�
�D��$ Zy�zm{�"O>�0��I�|��e�W{�Yq"O�0%�׮��1K���*)Y�ѣ"OT�"�H:fT�Er/�P����"Oޜ�#e_�]=l}������:�"O���g��'-�@���C�5"p�"O��@u�/8<D5�P��H0���P"O�)³%_�U��`�Pχd{0P��"Ol��Go}%�Vo@0�6`q"O,x�"`��)��b�.��i�n��"O���JN#5�Z[�LT���<K�"ON�dN�\��CmJ9�Ĉ9�"O����Ņ���*$�]�!�~!�T"O��Y�EЍ$��ѓ��&|�XD"O� � g�%��<�0KV^P2ds4*OC�D� \(�9U �f>t`�'��\x�A +A��$hL7���!�'���u���Y�L�XdO�9U�z\��'���MT/[D����#��K�bё�'a0ը����=�@�LBFfȣ�'������$^w�<	���7p/�p�	�'`qP'��Ul
׬B�d�0(�	�'H8g�",��!x��1X����	�'��-��nԥM8(ahsA�L�qH�'��"P��I���L�xa"j�'����FJ�V��x�A$r`n�k
�'%�%Ja�J��0�PM��m��e0������¹=�M��oːu� ��	�'�*R0�Sl��g�	sܤI��� �Q����@Z`m* l�d��"O���&
Z�	�-�ѫήk��jU"O\|��#΋9��m���
�Aw"O  ��Z�y˷(^�����"O��hp/f����7��YZ��e"O��O!_�LXƅ�>Sp��"O&��Q��~*dy�E�"I����"O���j��y#���&`����"OJ]��X�����W�<W�a��"O|�x`m��s�@��Z����j�-�y�'�ߒ �&*��M�n�b��#�yr�K�]����5�P�6]�AJ_��y��µ1&؊TB�w)Be����yb㎸z�5R��Кwu�G���yf��������|���rdH��y2��WQ&`RS"1y��l��O��y����L�ҵa�8 ��d�9�y�܄hx��Ł^����ȝ��y2�
���;����T��ت�g��yg��sg�l��Wф�r�B&�y'@�D�SeM�>�������yb�"f(ܘ"���:�M��	�#�y���
d���A��0:�v�H'��y�a��Z��u:%�7.p�iϝ�yҏ°;�x���Z��d0P*B��yb�9j��|�ǦF!<e��?�y��O�,�hu�M�N��8�A��y�� �k���b���I�j!c�"�y"݁fD�i�#ڊA�80;��'�y�!�!z���&*�6��۲$� �y�#��=*tT��̒*w����Շ�y�VW��@IP/�*���cw����yb@�����I��M�.o���q����y�
RD�!R��5.PHm[�#�)�y".ϣO��l:���N�۱��(�yr�J�r�@h�CɄ�d$a:�J��y�$$� 5rQ*�U  �PA��y�'R�u|��KV���5Ӱ`" (M��y�
�8)�֍��kW�	�)���8�y� W�a(��`c�C�d��F�<�y�ȳ!X�B�O[&sX=+&�)�y�@��a"�{Ɓ�#�8@�EH\��y"�ƍm�1k���fx���ԧ^�y�#D�A������adɈG_�y��\*���0_�Hbq����yr��D����R��,�a�H�yR��a�<���i�)�Ҡ���y�%##�}�&D�)$�D�fM\.��U}�����eL���ʃ�'e�9A���}&���g�IqCBɚ ]�	1q�FdTC䉏' �Q��i����EB7{X�B��h��U@oA�JʮI���;a���<����S�OI��@M�y�r�T�wu:��')D$HU�BY�H���DU�@�Ρɏ�d0<O���f��`6������C��U�&O�����	{VtX2N=v�Q�3(x�H��	�~f̠�(�eY䵑C�Y T�d�'X��$�i�})S�M&KV�Y�"\1ptk�a(D��s1�r�r��]bV�D�u�VB�	-ZX����W�.����-ǈ-�<B��2W7@ر�G�4 8P�H�A\C�Ɏa�v`)1�	�_�@
%E@G2"C�I�aB�$!�+S�,�'�ތPH�B�I��*�N$���oV�u�p)R�"O� $�) �7W&��96%S/ߊ%�"O.�ّ���S���	7D�f4p��1"O`(�G	�"���Q�ѬR&�Lz�"Oz\�妐��$���ѪGg�!Y�"Or��AD�uD��A�[J��8��ɇ�M3���G2\�h�Zc�S%R�>i��Lܦ���D��I
ba p���87_��⥉�;�R��GlQ�"~��/.Д�GN�<��];7l�E�<ٕ���gAp�S���&S펑1��\�'?�y�K�Q��اB�J� )�yBGR>? ��iW?#���)^=�y¯f��iډ��	�`
B�yRG=]|}!f�Z5�@኱��y���4H7� ��@��2�1�N�y�h�^ �bc�o�a�U��y¯�F�b���G�W��,#ê��yr�P��GR�PР|Pr%�.'\>!*�'��8�1툦o�e��'��+���@
�'�x8J��P��q !� h��}��)���':"�dEރt�&}$��m�����I$FҞƃ�jxEp���|� B��$Jj0m�aCB��xm߈q����<��h֕�4i��B��c(���"�^؞��=i%��.H,�!�Z�Eř��]�<��!��<1EI�x� �Q4(IW�<4�� ݚ���L=&.�	��{؟\�]#�̃�G� A�lcf◠^up�>IדK�
T eL" �$s㏞gR	��=�\��˟��΅KC� �h���IZy��Ѵ2�FI�lE)it��
���y�eZ4@�iB�bT�La�N��y"��IT��� T�Kɐ����1�yR��	U��s�ܶB�l�:%�ñ�>)N��!���H�t$k0AY��.��A�&D���U�S)C�p�7d���:��7���<Y˓6���1G_7�M�pm�-c������x��L��lI��_�Y�V��ȓU��ԩ�d�?+���s�� ��UU��� �U?$0`�:�F�1��ȓ"֨!:Ҥ��v����I���m�D"�����J���2���Ɯ�ȓ=-�� ��,���-x�2��PB�s8�(Dz��׃-}��
��׹e��4��gۺ�yb�P��娠�?H�d���lƽN����)�Sa��59��кA��c����6�z5vC�ɢ��X����Gy�L�/�?]�X�X��	z�t�=|v��3��)U�"�Ö-Ӱ<ш�$�]�\Xc��4X��}�1���$�P������ēm���Ä�:BUc�Њ�PȆ�L8x�!�1MN<1��fO�I
z��x�� '��p�Ń�/ߪ<��Y�g�>|��`,�I�-2���|2Յ�xht[f�0$ �y'�AT�<y�m�(�r��ڦ�Tu�րMN�<���C�H��<�0hE��F�:OEj�ybڟP<Q�*��O�Z��"��4>-Ѳ��x�S����ɅB&:�y�	#lf,4��
Ĵ0N��Ma���	]�%;����oN#&a�"�B�{!�0X��$ۡ/,"�X5i2�]�';r�Ii̓Jr�1��#�8�
pz3�_�T"��G��S�3ж�`j�?�w!��?��B�	&M�T!!�N����q��9��B����ʥlٞq�*�h��A��;�A(D�ذ+�����HF��8*�K6�$D�Dif-G>0��q��L�.t�ƅ*�-$�0�	� f�������HK��$0��
b"O�h�A߷x-�(SG�)�"���"O�l�iqןnb�J�J��W0�O~�=�Z�
_�8�tLD�H���ŕg�<�B�EfazE*شdq�,��e c�<	��!�����
R�n��X��a�<Y�+,Is���F*��.M��ʧ��H�<I���(t����������q�
L�<�$�$Hbl�jaEI�m�T�Z%��E�<!W���UCvK�/����p�[C�<	��V?l�(��i̢��	1��{����?�T�W)Z�-�Ю�/JH@a��y���$6O�l��7H8��!��*(��a�"O�i6���~.���'�3�^ C�"O�xyq���8�
�b�e��Q���Be�[~�P�P�J|J@�~�	2j�
a����X�J0JO7i�p����<aQ`�rd>L9Q��WQq�c��hO�'+���≕5��`��Y=��E~���Y�*��rcȘ(5�M��b��Rn�"<��h�x��������,�%�X��)��"j����R��Q��h� ąh{vB�I��M!w�՝�PL-q-:���i��=y�i�>���ȼ9�j�@���U�e�t$�1O6���E�3�B�X$�͊Z������(@�	R8���`�QI��u�IB:��G,(|O�;�4���UD��nQv�ꙫ1��h8!��U@��@J��(�*�ɱkS+O"�	ɟV�-�Sܧ68�{�ȓ2���S$ ��@�ēs��
���Р����>]��:�b��`�OL������s���n$Lw`��BӠ�8 ҫ!D�P����4l%���F(]�(_Ȩ��'A >	b�'9yنN,�rLs ~��P㓙�N�0����R}Dp���>�P�ȓ9:��X�@�Q�舷��&SPD��7�J�"Š{���P�$XWRXQ��-�b���CO9{�ZDd�
Lulm��du�E��O@1�F�,v�Q�6Z���pp"Oz�riY1r�9���F��Q�!"O��C��Ur�8���1�V4�t�3�X7?�I9v}H����Ƈh6���D!Q/s>B�	��e��D��m(�HJ�΍:#�U�'f���O?I��TR��6���@�\ECe2B��&�0�#�%2%f�ȳ"J�JeB����r�K0<:YRQ M5�JB�"� :Ĩ�2N&\RE�J�o^vC�	:�օ3���0U�iS���==1$C䉶|��)�Ɔ�W�~�J�P
bC��<O���g��Zx=x��C�NC�ɗUy���2�_	%y"m`��6NV�B�Ik`�YW�ހ@^�����n��B�I�n�L)E<
R.tІ�!��B�ɰq$��� ��OB*l�"��NC�I�Z:8咲��0u��i�̹n B�	�;�H�5�w�)aT��0�C䉫�V��*'�ft��E=
��C�	�#�e�� R�(� t�b�B�I o�����&�zj��p�?��C�ɖE0�xB�/Θ7�̭k�#D2�C�I��F`��e�	#&D��i2C�%&
5���R7`c>,���cנB䉹)��[Q�X5���HB�S�8C䉗L�l��g��R��(X7$[C�	�9��CM�Z�T`2⌗]OB�I�}0��1����n8�t��&�*B�)� ���Ƒ=x�E2��\O�)�"OL�¦�Ep�����@!j��S"O:=�b�$��l��o_�Z ��"O��)�gP3|�8�Ǝ�8CL�Q"OH�2�۾,P� +@�I�I��1�U"O�u%o�'R�5�:ۊ"�"O��D#�|k��p�ޘJ"OE��ڄ~��Q� �RE��"O���?eQ�+'��Io���`"O�9�Q��)Z��D��bH���"O��Q.�)��=��E�'���@"OL<�%%�&p<�X��|�@8I'"OJPI��gTLB���C�D;"OPA�H�*b�:�A%b�+A�DA{�"O���v�W2]��9"☔b���!�"O�0�$�:24�3�&^���{�"O�$��)W�Pp��'��+x��`�"OPCG�,DDt!I5@�?KZ��+�"O"��D��A2�e�ځ`��9�"O��E��FM�Q�aM�F��m�"O��bA�\k�I���ig��W"O�Q�d�O�M�$���Oͦuζ%��"O�Ⱥ��5Hf���72��]��"O��@�*'z(�=��� �� ���"O�`�&��@��}�mD�4���U"O�x��6e�
*Ьեw�lj�"O�[#��
�2�+��E���:�"O|I�&� /2��"·�%m���"O�Ѳ# T;:
:�R���z\�U��"O���aM4���BIHyn�;R"O���f)�is�FQ8fA���r"OL�%��F������=X�xi��"O�x(�#L�n8p{5nAT����"O0a)"0b�ґ.�B��"O����S?Or��*H��8�"O��T��=%H)�B*Ͼ��(("Of��2�!l��Q���3"i�"Oi��ҳtqZ�QQ��N``��� %�����"L^2���!��Nv1� J�X�\Ց!a�	�~�� S���퉶1kԽ� `��~0=F~$!��Y60hе�H�LR�M3mbҠc�a �6�d�:ӈO�$��&�:�4��HW��Q�s��&���ē��=
�/��!�"�K�6x�@��ɟ���+��3�Nxk��4;��9�ӹ"�&	K|ZD�_�B+�$zE%�eC
��!%ʆ"����ĕ!g� B*�T˛'B�y	�@Ӌ"�\��!"�p5d��	>�b`ϥxT��W�� # �L�g�:�D&2
iѳ@�DӇϚLD�m��<&�1����t��~�gD��M���4D$6"���X��2�>�h��-� tH��A��,ۜ�ca��xX���'Fˬn�@!�63���C��k���̟h+��ș:;P�WF��d � Q���0���s�ԍ~e� �Ec�'0�"Jي#+�h{�f�[5�~Ҁ�j[��rl�3E8�HSH	!-�Ĭ�V��&���1s$R�0��0���(oYĠrb,_�4H2�PC8����6%�"�$�Q'�IgH�q#�ŕI!��M`�x�͘g!��B��,�?���T�7����Ù�Y��X�#�+\R	
�:8���%L�	6����%4���#�\� �'��Pq!�ٞ<�@�4�?�A��O8��wh��y��r���(- ��s�mIS/B�CZ��ei(��нB�>D��OP��`f� XY�C�KB�T� �'N^����A%k��Yg��&r8�m:7DT�~r@���$� L�"�{�.�K�v��t�H)u�Ͳ����B�b��6L�^�J���n,�p?�6+>�� 0�MB�O�>\Bc�;t�����荃r�(����§1̨{7�=?��  ��I�6PJ�'u����Ch̀cw��y�<Tj\��f N�$��u��3k�s*O5x�9�%�����c�j��TŒ�Ylm�%I۪bO.�:6O�MY2=����$X����䓫f�p���ӂ\�=8�[�S����AӉ��2���O���F%[+t|q�!Ǉ�y�ް:`(Y��"G0jP�Z7*��!I��:��V��([��mQ����4Y냋�cVn����:�l�,]�4�#d��� ��T,y!H�V�O��5Γ[B݊�b�i�>}�Dj�"g���0��i�F���$
�h����P"#�$aqh�Q�����ꆍ
-:
��ɋA"�+W�<,����_��̐1X<)��ii<zH�U)�O����+T�0�1n�G#D�r6���7F˟����J�$����dK�
Ò��"
���� 0�AI#���%"H.Oh&|��'�,�LQ�\"�����6�
0� �	"���u���Nk t��@�a��N� 4�b0%�r����w�8�I�\HD�q�x"ep����'Cؖ\�БӀ�A��F(�Pi�~���@�J;�:AJ�"�2���K�������(O�=�3���q��% T��K�h��D� �~�c�'ƵØO�|�S�g�E�P0g�̆u͐ɒ�L��XD��$Lw��|H��'���3�ً]}H`��[S,3�-�?"���Ѝ{��_B�NȺ�"�1��ĲB@�Ok�\,r�$s�	�$S�T�E
�V!򤛾10��� �V�0VZ�k�*�}���	�D��b* S2�+X�¢~j����
��%v
:1ф(: o�A�I�1Ӏ 20����0���BlQ#?�v$�e��<>p�J�iܿ�?��͇�Zv��3���})�Y)��iG%B�,b�(��IOw����M��A%S'�q����;J�������J�I'탖U�)Q �@1*�`lD	v�:"?yW	p�Uq5�S�S}�����w��\����~��g���:��=�gD{�~�C��Z�iE��?�2��J4�r%�+�
��7�	�ۦ���=*�`�f��T?���]?Q82�Ϻ\��Y$+K�p���rV�>� ��ZQ����D�1	� ����8g�@\ktφSh~@;t.@6"���[F��4D�j� ���G�x�ϙx�OE��]u��u���|��%���ei����~��-6|�H���{���#T�N$"�;p��.��6�.(r���"U�+A���v�8��C�U�D<�<1ÏC"W�f���U,��"��D
k����F=Ɋa@�b8ړ`� ���Ø3s�Y��d�;�b%#�����Q
�c�u��sMװ6��U1��D؛a��h�/R�Zʓ/U
1���נ'����"�����<���;��-��	n%"�Ξ�D#����?������!�&o[+f#f��7@:}�^6W�@��/�t>A؂��L̮J�	�o۶[�))��d�K#G��	�F�Z31��U���)N��N .0�Q���,�A����8���=�e������	/�\< 6j�hʒ0���w�U�2Ʌ�d��%�l�: �n��.�RP��ɊYj�8;gͲH}^���n%��$�$<(�YSe�F�Cd&bߤ)S�N�Yr��D	!v�MBF�01�����&i9f��8��<h��C�f�x��<y�n��b�n����g�D���L2�2�H���?��H<
��\�S���l�,��`&=D�4�! W5aC��yN��[RN��b6�
��G!h�\�ka�<!�R�p��I��W(���ڀ�@��6���YSE�/!�$�!A����a�\�#Ĳj�.J�m� �j�����a�,�!﮸�F`M�C���Gz� �Q�D�#dkގw����e읒�0=��:ap�J&�ȁΪ�B�&��!�H���� �w��I�6Aº7k��϶���	ҵICo<�aȂ�"G�@�jp ��M�����<���M	��sVL�-v� �f�0z�Ќ�O���ĈG<M��0h:�!Ss�@�~�����tX�$a�X�pd��bFB�)ID�	��\�e��S�f܃.c"����!����qf��2�
+LL��1O�m��AB$��C"�	!\��	;��	#X��);O�h�(�!�h��� �<>�q�M@�D�,�Bb�׺/4��s ���X��.%�|��B�S�> <�a�-�E��,1q� (��)� �
��@PM	�U�E�@�8�[�I�4����jl�+A!x*���xJP� �7#����8������l|+ &�3��N�|��wm������iL��[�hj*zHK>Q�(υk.pP(��ZXnQ�.����a�̚j|d]��U)8��**I�i�~TG�ߴ*fF�Pc�S��l���$p��A�BF�+ 1��Ej	7i�zXw��XA��m��Y��`�[��PB�ޔV{�t�&I_�y��� '��Ua���i��y� ��^��-@B/�U}ȼ���@�[qr� �C:d_��{�+]  �%g�P�6�v���3g���@ ʓ_
 ) ���.?�������聃�� �����H	M�,��._�~��9XG7��X��R�;��G�ާsE8BY�@;>�k���w�xB'-J;n.�qH�C��7��`J�ƛ<�|�`�Zw����d��`���.���C�L4\��+V�ȧ^��R�J>V��u�A��`��L�u!�/���5,�6Z�nJ��u�B�� �8V�3�� ��O�!+�i��m��I��
	���O6��Ã$*YRa����U�?OLX�kuJ%
��[���^=ճ�9P�}
� ^<�䵃��MKH�;�
P'�MKa�NP� +��sU�a�Fh
�}�`@� 0�?1g��'h���a��V�8K���7u]�]¶�k���������Ӗ��'�؃��:/��D���J=n���*�B�;ǂ��B�̕	��b�X+#��j>�hI��Slelh�u/��{ۺ �v#��18����4Z��0�'��m1�'���7��i8ި�e	NB�P9�ĥR�5�m�r�pu�ÆѨVJ,u�=q�Ȕ*!��`��(�j,Ԝ+��4,��S��.0\�6ϣ�^�C���>�j7-�8���I�C�wl4x�Ǜ.(Tz��#,A2��H��c�-c�(E�� @ɶ��'VP� T�=?���K�� b�ȉ�aK�0'�р)����(�HN�;bhĂJ޾$�RoM�1gΝ�Bb��;�r%��˲(�� S��]:(!����nցL۲8�2�M20eȉ��"K=�h	���f���<�I���M�:
dY0�i��k �Y��5;kր�@W�c���Q��:�v�MQ~����ӜG8�aP ^�Y�]��b9R��K���6	�)���4^!�X��%�B3�MS� �b�B1�Y
�2���w���y��0��
R��e�0�J�{������-��l�zpqC��b�q��^�� I[�=�H!��jݼ	+��_�p��A��. FP���{2`" ��|�fM���������
��aV"q� ����K�FT�%��`��g�`82w+�x^��t��3��QG�w�$���e��FU��C9w�E�3���%9 ڒ
��!o��f�>	�E�Eд!m�3
r�qdFD\Xт �M�Dݘ1��'#^4��#mӗ_�nH�
I���5�%�ܡ:�2m�%ɇ4��x��#]5��'PƠj2�>o�~�0� j���-�-�p�0��K;��,Ӵ�>;�H��PIF
$���1(	3O�`��D��z�8��~b��7��t��B�adm�`%�l���)�I!|VA�W���V�H���ȴ�F#cbe�?a� ]�W	������N�g`��
��`� �m�Ș�g)�~��`�V
�ن�LȦ�P����4�۱j�e�@�5���]���#�L	�e6�@^�����\���3����Qs�g9����(�V�ּge�řv�� 	Yhx��!o7b�CF��j72��%��8<��cW<fd�ٹF�� 	^�"�@4����*�r�BQM\{�'��]@1��W�~�����>j��F�iT��I#��R��ؒCc�qx$�0b�\�q1b[-F
�5df�TG<��ş'��ZL?af,S?-��k�J��K���C��B	i�LP���L�w�����	8�:�Цi�5�M���\�21�S��<�����l���@�ԇ�9S~�PQ%a <b��1��`n�ա��U'\DiX�o2t�<���\�R�x��5��'��u��V�j���d�����}aWǖ<�"5��)[�Lzq+vxv��f�]�6��hI�@�!�\�#��z��+�H�a��0r΀e�'��B�d�!��R�e�&@�ܔ
�Lґt�`��'Æ�vw�i��M)0�&aghW�z>d${gg[%F�°ZSL��s�f���1r�q2��ѧf�V�8��̗Tu�!�Ä1��Op�PA��K�r�h_-��Zw$Z�mZ%c��� ��˱J�`Ls�g�4r%�+� ؈|�(�$�G7sqVdC�b
3T��`@�
0H�f@k�'��r'�e Y�v00Kխ�,�FQ��D��,����C2W�(�2�Jb\F$�A�O�4<c��R. �Xey6Ņ�&���i�3T�T5��3h�&��ԊC�?d���E�1I�	��-��O�&�xQ.P^-A��1n��|���{s��+�ř�w���4dkӀY�"�yİ ��.����t���ش(�����l˳k�N%�qI�iV�q[���(&3��� j�`�b���`FF�
������Ez"��
i�qٲ��2&+R����ٹ|W�Q�G�{�bH���i@������$/v�u�7F�g꤭�&��:y]�q���4z�d<8f�ۙjH���瀌�
(.�BY�[t�9�4#���gK&�� �^�4v>�� j�xzb���	��G&:Â��U*ݫGd��gM  tp�L�� B�Y=l
8�PҜeH��z��0ی��&@��	7"Ű��ʗ@P�0Wf�j�\�j�,� �PaԥɁumx=��'��Š�BJ�F\� h����n�J�2l\-�d�r���l�=q`��F��,�T񉶮X���XH��d�jq��i�Q��w`/�^���M�3�����w�@H��_[�8��#&�#1S��b2��� _����l8c�
C%�,%���Z!HP�r+0��GN��MH��!� ��2�"#����+�G�W:f`�c�2�^Y W��g�&Гug �sU0[�	�v��mq���?[q����1�Fq@')_g�8�Ӆ�A�vR );1�@	r@�G�_�V���J�m	)/H�O�!�剃�,��N���ɔ'^�����9L��Z�OϓCo$�Af��1�"���DY�e��0Q$�Rd�5�P�:D��2��Fg*�Y6H�3�r�GsN +��A
;,F-#v�U��~DiQ�3q?��B�O\��p��U?��E��%�4
L�_;��0ƌ�[h���1)G��r�ނ`�
y�5�ΏȨ���ʯ�%��0�/���۶���4�5��K�N���4u�0<9��3'@xpY1�+S�e'B�?y�DF��ح���q�H�yQ�\1"�8�c�@�#�\�u-����O���D,Π���kE5Qp^W�)�`B���"Z����B�t~�I�r��$A��0�ը�˟�a���.v�tz���#Y���ؗBpw�e��$
�;�ސz�Nb��)yTLMQ���7�|�k�H ��L�e��S���H�9'���b�Y��P�ю]�_K6 I�(�1$�ZHASIM%��yådC3�nS�ȅ�6��t�A�ܴZA"	ӈ�p�d	)0�.iӥ�ԗW~�`�U��B#-��\(NyAe�0ʱ!��I(3�>M�b�^j0�� �Z��s�К��	�Э��jX�ƒ�ON
�� ��^P�aꗂ!n&����i�Y�GM1i�1�D�H�@�p{BOԐyS�Y�M[��sT	� ��X�m��(; i��s�8 �6d�7��	^zت��U�<N��tq�.^�u���	52�F �g	�+�@���)_�}����Qm�LBg�ݻ?�5�����]�=+��'u�ʕ�������͟�;G�i@z�
��{���H�bN�f��rBR5�p����E-�����399�1��Y���C�nI("x(��ͧe� �%�0}a��;C��*IT@*��� X%��7f�=1�N�n�
I��X�녶e���G�x>����� ZF��>�� �� ���a�N"f�ny�c� ,T��k����42�+;�� ���
���΅�*�`��w�>�[v��'s��U��>3��)�I�>c�8\
�K�E�'T$���Р)̹ؐ��8TE��Ȱ��,Yob�"\
3��*Ъ��У ґ�.��՘O��	#Ę/:X,Zufǚ	�2�2�1@ў)�˄��@��F�O�D�w���*�8�9#�Ǟ|l�Ó�2#����-��6�d��ga�:tj	{�*�Do.�?Ƥ�3_�EH���O�� ǘ&$K�-R`��Q~��OO�8�׹'n>��〉� �0�DH3A~�cR&��9��];�-ެg�p�p�@�$>`i�������	B�X���'��}��-d�z�h�`�~ΓM�h�6I�%��Ҧ'�6m0њ�G�b��U��(�npQ��!-N�z�I�	X������жl&����P8�x��¯~@|��&�1t�X}��$�҇�uf�8{w	U���O�xj�	X���
"+�T�9�D+TئĲ��Y�X�|�RT�G�F�j���NǊ����V#)�P��|�s�^�|\b�"��|h��H�;s�E~#p�� ��S9E�&�y��}�CnS4;����щ����Ș�>�:Q���������^o��1�~�/{��aK���h���9�Mj갈���^�	k趄�������ěb��������i�d�a�lY�of�3��B�xY5��Q��!�07�y���T�,�yƢ|nڒq1xDȲ+����5�Ȋf
j%	��<yo�#(�!�����R��_����l������,�HX�5ȑ� �����syr�V�F�P0RNNX��(%��E
@P�Y� �򥈷�S��mX�@�d��q�xZ*��IeGF�ؤ� �K*� �](N�!���$Y�XR�%�,5��ԣ6X!�ĔM������T" ���;nC!�$����ɠ�;($	Ӕ�ʚy!�$D>1�2�p@B�*x����!�� �l9����!վ)(�H9m����"O$Űu)�9f���
@�:[�zHx�"O�*�
97��Rd]�"v���"O�ha��H<T��K�E�:e� %"Oz��"�	����"#��e%�"O6(���̟`�����&�t��"O� �l�.~�2�f�ND0��"O�Z%�G
`��і��Y5�` "Oju�c(KO����B�s?P�:�"O��R�Ӟ#�b���ɽ��}��"O�zD�.It[��8j͞d��"O �U�þU,� �!� f�4m��"ORQ�sΏ4f�r� ��7 �h�J"Oʉ��K�H��5a�@�@��`"O����*8p����)F���pS"O@��d��_t2ͺ�ㇷ[t����"O��@ :t"`<����Q&y��"O�36���N��m�%o׮[ ��"O ��4G�7n84�1HCQ�x��"O&�g �f�PC�U��:�)�"Or��qI�a��際���"O�]�6�1�Zl�4�?`�j�b�"O�83����8�)�G�
UVYI5"Oؼ���!q519�F�&�(��"O-��� � ��=#Ή6W�س�"OQ�BGE���p �(<>��"O|(�`m��`��dΐ����P"Ou��!� ���(P0>���"Of�@Ҍ��?㤈������"O�bB7n(�REÅ�7��a�"O�����J#�&� \�	6`(A"O"���/:o��}H�nD=kRB4"O!dǃ�BQ���+E���T��"O�كPD�4|�6��CJ�Bx�\2C"O�Q���Ł�F�p��^~����"O�T�#��/_���tҙL�x��"O��խ�q�Ś��ҼCyb=��"OZ�@�,]�`�
u�GyzpT�#"OxP�fJ�SS�y�Ӧ�n}�[q"O��x���[R�U:�ŒnH)Hc"O�9�e+���v�1'���7���"O���Omi2I+%jگP�ʵX�����BMv�O����f�zT(�����5�d��kX#mʤ����4�4lOh�E'�1�P��ܽM4��a��Yv�}�OjX+r�A����@�+\^����F5�
$�N�`AyEi�,�rHHE�RLC��-Y�^`K����_�|qXa(5
��1�J7�6���(��\���J1�\���\�xu$>�����/ơ���?}fQH���50A�x��[�,U��5�U��� ͓Lv��p����
�,W�=μ�����$P��j�b�|�L��?��P����:��x����0��`�P�R4ѕ#,ɋZ�'�����@Y�1�p�"�X�ǘ��1@0��$!�"Eu1�����;s����aG�Q/Zhpwɭ)6��	��<�ЫT�@x�X�E�C+��%�mD#�X�2���?��N�38�X ��KT*Dr�p��	�)���3D��D�j���(�h�r� ݿal��
�d[����:*$&t�ЅL/k�,����2N��-�2�ä^������
1h	���ۓ/n"|��E�/j�6����w>%�rf�V&5����"jf�ن�Q���X˶�'E� i���Z�X�$74�bnܬoͶ,����U����ON/������yNM9%IV���r.�-mʦ�7��P����O�0�ȗw	a���0m�(U���0ڲ�Nd�m�� �����ݩ�Z"L�R1�#!0����$B��4��dI�&G4YGua�+N%�+3�	�"abX�Ed1O@�AK��&��@䓷h�
q"T�U���PB+�I�YVLa�&mܞ�$��*;<f`#L�k��=HQioBDaVɐ�7��~2�M1vX�M��Ð=p���I(r*����\8 �נ����Q(Z�U�у�w����Op,���]������M=&m����-:	�n�%Q�
e�L�1h��?�p�t7ؼ�F��:p?z�`�o��!��Bw�o�d�kwÖ���|�@�˯p=Έ���V�t5n�'p�`�u�$>Z����T@�N��ZC�99��P͎�-��䇫6�lŁ� ������7P�x�X�FJ8u�L5��i�&YS>i3e释Fl���͕�8�@a���v䧀 .�y����0k:�[�NT�hubA����t,�u�6OFY�6GV7p:�1B_63l6�{��զ͒��O8�T�� O�N�T���ؽ
0�B	_��U�Tk%�O�-@�­*�P��E��	#O��6�"� S�w/��yD�^�?!P�O&�`�O�� �YV�t�$"�,O=�-CWbD�)��,1ϓO?�![g��(���H��,-$�pzP�d����=O������Ya&N�j�:I�W��"�lB0k�e�������M�1�E�sb�C��Ō}y�5����k�<О��T�5��E|}�!��)ު�Z\2bc�*u��#�,�6��`���'0��r'���r���
Qh :rӟQ���,Ѳ��Q��aO�1� ��:��A0L7l٢d$1�4H3W�Y �>���̐�7A���1)_o�� � ��)<��Y3D,�Oj�WLk�V|BdA&'�T)I"�� }�9���d�>c��x����' ��*	ҟ֘�$�2Q�'�|�����%A��C�I�U�$�i����iA'��<�^�L��a�-J�52͙��*���V0��G_�Lx:4L��)����|"l�+���=�}:���"40��K^,;�r��ǿ��1jC@�O�ɚ#@#Q�f�'>c�Z�I=x�����%9�W

�$���'v8r��T�g?!��LD��j�����8@+DV${t +3��)P�> �`)ô��O$ɃCyLJ�4�
�]�$0r�]!"���/Q� v�$�E��#&]qO��
�P�+�=����z���S�IB��%)�g@.��b���#��w3�A
��,K̴ ;A؄3��O-F&�Z
�0ؙGd�
F }(�O�X��!ξ&�B�x�	�!�~����OD!�#E֒t.���R�_�(Y:Mє��<Vh1	g��+b�������y'.L(iV�E�Y,��`�ƚ$�̬��&������\8�%?�()�Ɇk����UG�'j$15��V�l�v�
�Zs. S��V��)!�n�i�1O�!9���4�:���ȼDR8���ĽJ��U�@MC}Ȇ�C��DQ�r��%�5�m���5Q!(��G0xh�%B0o$j���Mܑ����a��H�D����aC�/�˓p��@�挀����P`C`~��<�p��cl�Z��&j�p���&�)֡�?ep�%	yOL���:��ȸ�3}§��w���Q�_f>�8�ַ,Є�!ԩ�t|�%(G�zM�� L
KV��솄]�p� $��C�C?�.^���"�a������(�[�!�=I�#-����I4��i� U��ˆ]�Xa�KQF�ei `P�@�u,Դ��9A�I2)�T�	WZB�����*�����!g�nP���w�UA4j� �ޅ�W��@�L�S�J�&j�|h ���p�	�(f�h7�4J�|�j�%_�F��h�<yօ��B��\�P׊r��i넍�(bV�!JT��?Y:iI)�F��"��G~�l*�e&D�� Ѐ����Y�3c�L�!��5&�f48p��00�C��&J�I{R�A�'vՒ��;Z��1Vb����E9� 6���[*���o����cgJ+&��:5IAJg���V雿8|��J�@�(P�`�DZj�'*HÒ�T9/��33��+j1�\�ӓr���YcdT6H��� ��%��x��$E%@��pe��,�r�ch��zLTLY�ON���d����O�a1� ��gK$��� t�2�w��v�"-���Z��eS�$�>HR�\>!P1Aߙ�n�S��{m�|Jb�+�ѡ�;T�a}҅�U�
<����
�(q�Cn	~U�@	��A��H`˒�9�$���U�4��o���"e�cN	�<Q%H�d��(3�k�w�������7��w����׷�0<A@�R�������3>�je2�֚f"ᱰ���E���c�'p�l�iPfR���@�̱=�bm:�OVe$�s�9j�9Yb띩p�I��Ƒ9$�����	-v�����.@ꀬ�D�H�"�B)�!�c�LF�����H%*�,�:�a]3;1��YD��F�X�r(�!�cE���wz<�i��X+�L�Ed)7�J��I>�e$٩6�@���'�T��Ɂ-��3��L{T-b��] l�����G�ֽ�\Rp.Q�0T�x�G]�`�P}�#�� �(eM�mw�9:��';#�D���\����̂c���n +�~��jŬ~��$0��`� ��1/���L��w���f�
�[F�+�v�� ��wۄh�HA1E�2��͸8�~A�툧p�c$-R�Y���˳.Ǒu�Q�I�-��]o<��$�P8 ��uJ�*�J�⥦�J������Y�^����+\k6��$�P9%��E�ī�X��%��
������. ,��P�$������H>jݺ"<�w-ۖ7TxA�K&�I>B����/��ð�K*�I!c�\h���(���FY�6P8�U�W,)��� ՗G0��*���B%�G�Q�м��(U�0�"�A�'\%F[�Z%U����:N��t1t(i�ّ�� Z8l�C��/�V@�}�j<
���8-� �2��5
����Lơ%R6x�B΢+�B5@�@z�~1�d�H��j�Iq�J!GF�}�j�K����Ѝ�O�Z$�u�t-��		�r��@K�@I�Ah�4�퀧i��z�h��x��,���B�89�A��bI�}�����i��2t�c�%()�b���7�
�;��I�!
�R��u��'p�`�c�&��y���r�PRg��<��'s�l:w�l!�+]H������S̎!x �G,�Z��1]-*� *���֕\�
�� 5"|i�J͍ �<!�u��4|L���H������R�_ �]#�4I_�iq&��>r�iz���7l4��Ee��kg�Ч�5&ƀ�|3B���3?��"�P���dey(p��^#y�����Z��Ui���z��wh40��#��n��BC��"����f4m2����aȪ2]0X��i�h�ƃ,m��bsER%�ى0�N�h8��B#�K:	�lZrc�8Y��!*�	�22����@��''2��E�#f�{�ꊹ�D�aӪ�S��ҠamHQ�����Þ����L�i*�y`EEz'F�ᐭ�9{����@F�\F��'D_�^N�AGl?��Rw-1k�ԉ3 �(mb��C
�s�$)�v(��6�n�"�`h�Eۥe��G�S ��h
� �=��Oܻx�N�sB�#b�xj�#�0?�ޑۧԽf"qO��sf
^1
1+@ӊє��ǆ�*E9h����>m��Bf"L�bd��u�T,�q�7[���t&B�*C
 WL�0y��lݑ� -J>�49�Bd[�H)��2b�?>���'�Vt��'|{����'��#S�D#���6[D`�g'[vjA���Xg4�Ҥޱu'��'��([L��e��/H�q/ ���f�([B��O�ґh�._�|S�x�&ݎ ���F�29� <:2��W��� ��]0b��J�!'g�!Q�#������9���H�vKV�B�C+uxB�a"��1b�a����th�T!w�Ś'�X+&�&i�	'FN�w}H�Ib�q�1�>�@V�[�~�j�A�%~�5��ejܰl�(r`|�ǂF�R�:�Xf�F�[�v�n�O�Xܐe�V�̔Q�w߂C*>�mP�'\P��JX'y-�	x�BÐ�Q��1-Љ&_L�'��~ T0"�P6�CF�^.l3��{D��Vwyp��dg���F#>D�JJ%�І5�8�_-m0��CɄ!Vw���e�-�h�Z�k�0|d0ɂ�ɖEP}�k�o?L�����5mUѮx�%j[�e�"��u� �"@R��&[��eh&�_� �!�¥F�4h�U�[d� �O��O�Z��9@��&I��%0���'2��@s��m�D�T�����TCǂw6M�;�*�b���9�p�x��k �y�pJR�ڥ>W�H������Ɂ&'`�H�/z:n��Sl�ۤ S�'���`���-l�J�R�_<X��si�6������ ��ɓ5������6^�^9Q�_�	Q�����r!�Ã�6z�p���3��!
�`�0>5��� �N�'�> ��(ŀ]�.����\r��v�I�-�h�r��R/{k�P�5gޯh#����/�u'+�$�f��WK['���аO��ᇡ�0v�9U�U�b��uä�h�'��m����^sB�P����iJ�=	>�3P�K<!�va;�ŀ$id��8�־ Ը�{B���$PhFZ�d�`�sЍJ�"�pm#�� �ie�����ެ����R��TtIC{h��C�r��1%�C���V���W��hx�	 �@~b��"Һ8[8�������&�$���� �|C�Ey� ˼c�"�.�) ������"<�k���Р�%�q�<���O�<���~Q��jg��N��|�t����܈�e�u���N5N�� 9� �)bGH\��͐%DDy�ub� ��J���'z�
Q��I3����̨����r+��`�.i�
K�d9ڬ��j�>.�.=b�����jF����ћ�� a�(e�@*J�`>k,�)~>.��@�@�[��i��U�a~�j�ZAZ٣�` 51�@J�!��3���(��)@@;cI�a?�W+NN5*��ۚN��0��y�T�bq�" 	��Qщ�!.�pT*�mYF�r ��$�K�'� �R�F�$тi!Do�E&��) �a�֔���.as�l��Dوm���p���NG"�B�
�F���v+Kc�ư�Dd"ʓu#X �FM��A��#�֑*`��k'�=h�VO��t��C�9'x�v� #�b���K��
=d�KA⁒Q��pQ��/^�8fR
R\<)%N�F���Z��'W�C��z�ZL��VM�4��ѿr"���Ť^xEफ �[�+B��y�TL���W�J��wA&\�'I�R�R\c��_�B����=� $���>M����(s�FU��OZ�F��4��o`�
�K𬁕n�<H���� �G�u�R�{��Z�B�OX���p���u�A!,ް�	�&Z3W�h��=A��~7���f�.P
A�Fm��2܊���_�~�nLY@�[oռaPQ��#o�>�w�G (�����-(���}���8 'R&^4��2g���F��+%��M����Q�I�!pM�Lz��O&H�` ��4]� i�K��h�d�#=�,����.��Ɓ��x9F�J�$U9$��pN�?a�d�m�)��O�y�9 A)V&gᄈ�Af[i��t�Wa݂�|��	a��V��y�!8�)W$c銨��ڑ~o�q� M��4s�I���7t^��'h��t/[�m�<�M��ECW���c��i��ݖ'@ꙑ7 ��4U�AJ�_C�0��.ٙ��Zs���#���$�J锍ё`߫0\,Sb�[D� �O�	r�W�)��|	���++�W���%�p���j��!��M��bءvH�)��,��PYr�_,$�%�D��ғ$�\!�|x�i�=��]"��_�H���E��C�`���-�'������~� G&SGx��&��G����i�7r�TR�d�'	`\�d��@2�mܦ�r����5'� B��K��e���1�0����*�LJ�bF�:�� �f��(��ހO��$ ��Xer ��@�,�����LU��D�$[�-h��*"-�< �I�7O�![ɟ$�i�i�:���l�W��Ѯ�~(�{�/@�`�j�!���<B��_�ʖ��� >ܝ����Wd^˞����&7��0M���y��\�
�Zԓ5�Id�̭�`��'��a�����=�l�q8��S�8p糟DAՉR�H��!A�&h�<`[cȆ�R�<�4���S�E�V�B76�bde)N��1y�a�$l�$hC#��U�(Q����6^Rx�ip �c.�ܫ1$���d�ue����XV��?FTPG{b��/��!5�B�U攪��]�t=�x��ޜQ�"ae ϫm��3ǃ� .��a�/ÒP	耲���͚�ֈ��%s�&��a�xբ���#4g0$z�];L��d(�`�5i"Hh�ʐ'mz��;2�[�4���x󃛁7�m�v�K�'��q"���	32��OJZE���enlspfԢI:�x���M�z�J�X6�IJz��'���j�l����:E�G5�yՏޫ���H�i�-R�b��@�[TE��c�!fY�EP��^5C_�h1Q�3�%26���%�]ZY���ڠg[���<Y�h%U<V���d�nKv�Ӑ�N���Lb�U�O�<�$�;T��apH�'P6B��Q�̃lLz�ˠ����scB�"fz��c)ÙbBPC	��?��\j�x��& ܞQb��-��x�t���'�(m��I2GB����逤J��x�+ӥMł[t$�-�d�4IM $�"��,)�JH:��6#�<��$h6��5W�¡���3���10�2y���޴HI8��S���m���r�9B��4a�[<q �馁�.*�n�$/�Dָ�OW����DԾ��3G��{�̰��\y�"��	��#��O �ƹ��P��~��;'�5
C�ib�hH�f��Q3.�oM�4K@��!�dA��)_�:y��d2f�m� �Vy�S��M�!��njl�0BI�2��Lpv���XD�'��xr�Y1�?q1IB.�@�ߟ��1�w�(�T����!��
��5�-OfP�2��z+��˓t�>Ӏ-M��j���\�3 �Y'�S0���� �֡xX��Q>K`B�"$�0��O"&
���$�&D�� X]��b�<�X���`��9#"O�|x�S�W��J�X��v�;�"O��B%ܢj��%`�jn�4�c""O��KC�iX؉̢ �4"O�5��B�f�l�GM-�xP�"O P�U�G:[��5�Ѝ660p 0�"ONaB����)������&j�,y�"O����i�B ��aW�2lzث"OΜ����OQ
�0�&%Sе"O��w�]	\B 	���gz� B"O��E\-�𹐳�-�%a�"O�=���3�r$f�P*����@"O8��e�4Ff�H`�:nL�mK�"O.�����/5�(�F$� _�ryc�"O*����8A��äB�#�f�"�"O��2c-��gS��A�#8��a�"O�!�C| ��Ţ>dW~��"O�k��ƟO��	���fY��@r"O|�E�� H�� �
S%v �Qq�"O��!��ޤ;���X�*�0+$����"OZ飰�W*�����(N�,�d��g"O���5j	9�q#�(��]-��q�"Od��fD*y� ��F�>Uv���"O,|�G!\(W���� �P|�}��"O��y��[*\�����!p�i�����n,�t9�oĦ���	�!���e�K8W�i�NwT��r��y2����y/�����SoSX3A�	j�(xڦ���������u��'m��)�'L)JlZ7 Q�V� �8\�@�ʄ�d���J5?Q��Ib�B�� ���/+K�d�
�`T��:P�.��'ȶ����O�IުG�P��@ǝ�R���sǫ����r�{����2�JՇ:��%�UH�ENR$Q�Z�L�B�Or�lih�:q+p�O��!�EHڷ6��)�d�N�L�}�b�U����:XX4��E��W���[r���: xD�-�?]h0�I� �ݡ��<���OQ>�[蘾n��YQMX�g���t,Y&5����V��Ԇqp�O0��c?�
k"���$�U"T�G�Y0��'}�g&�H���P�o���0��Ґ.I23O�',X�t�ԟ`��	�{�TT��r3l�����3t<Od�X#L�����O�JeMӸ!L:캀"K�W���Y�O�	i�A����'��3�I�G��GGSY)ڠp���&]�ڥr��!}u6�"}b��O�"�,��V_�����R�a�j���R���aٛV�qӑ?�WLR��±��)sT�Ap�w�0���2�ȟ<����E+J�2XI��	}�4qp��i2��`UY���wnS�<E��(V:@�Ph��'G*���7K�%�`��'�:=Z1]�����  y�!�|���q�L���$�����	��>�M~�0�e��&=�l�iƎ8ʈ���]w|�	;��S���	-ϸ�#�G�?b�y��8*�"��ڴ2a��`O<��ɧr�KQ�f�N}�'i�VTLb�2P�c��|r�Y��0|�bjOj0
�8$L�$7$�r�����7%�b��n>��b�&����e�(3C����3D�H�G!�\ D���l��p�4A$D���#$M3iGZ؊BV�!��c�!D�dpq�	'Z�:�r�� @��a� D��rE�Rs_ry3Ce����I D��B��� @�����՜bG��)�"D���f��2$
	s�Th����>D��y�(�=N�x{$�S�yU�)�G<D�h�5D+{�4ġ�ßw�V��1�<D�D�a��.|�ak���1#��(=D�Xp&E�E�$,�Q�N�W):VJ-D��)_%~Ĭ�����^�(�t.D��b��؅8G��W
J�4p؇�(D�Ԋ���Vy�&��EFu��C��4u�p�6��&|*u�$遰TC䉧!'ԤH�j��Sy-HP�A�fC�)� Ȱ ����$h�� pi�)�-i�"O(ѥ�B M��sN�N��mˡ"OI�O�y�B�@W��yC���"O��#�"eP\#����v'؁Cg"OR�xUy�%�D.L�qS"O4���\��GҘ��i)�"O������$mN��5F�F��-{Q"O8���D6ip���ǃ.>L.�"O�5�c� �>��e2���k�؅��"O��
��D���R����Lm*�"OXܒe�P�Sw�D����&��A"O��xC�X������6o����"O�I��jO�~���V��HQ"Oʠ��he����p��9u�����"O�H�a�[� o0,�����>�2���"O.�C�+ƿY�� S
Fw�Ёy�"O�]:�)�?y"tp�$L�)�V"O8��BD��fi�Y�� {;P��c"O��U��)�UK��ς#4H}K�"O��R���p�~,ɳ�#z%>��a"O��D�J$'�f̺��R�1�Q*�"O�<� F�[k����.�z�<�T"O`yr� 	���q-]��%��"OhURЄV�Z�JE���"�V�"O����ȭ�X��+��,��"OhE1Pđsq�H�P�ܹ���"Or�pa'@h���a0�̾@�̭sQ"O�x21f��d�D1�1E�DZ�X�"O:�uᄪZ�>��2j��e��c"O~���<>�x��$hPtG��h�6D�����O�2�re&λ��s��&D�d!�NJ99�n���c.(����i%D���Wh�(ViH1���Q%D�����]x6LA�DS�A�r�QAK%D���qh"@�L�!-Л8]N��f>D�T���ʟsDv��rgH�d,(\K�;D���(a8L�	��E6@��h��:D��@D���`J܈!���]|�,�tI$D�h�K&v���h��X���5�%D� �t%T?7G��0�J.o>�j�O%D�ċ���@��$���U K��"@d6D��I��p���L.D=��IM5'�4C�I]!�\#�)+=�I��YC�I5v�D-�OU�H���-�>VcBB�I�DȆ��%�-xv�4qvMԻ��B�	�]�T�z�#@�@�XtC0 �'tC� @��9��kŲaaY�AN�c�B����$�Uן튭ॠ�7|��B�ɱ`�Z$���]�_�|a2BO5HβB��+(~�*R۹?\⽳�i�8�`B�ɔѴmB5�7Onّ I��)�bC�ɇi�p�ht���_�Fݛ��À9d`C��GS( ��#L���3A�&�JC䉷2A�9��ۥ"�I)���ofC�	�r�J=3$�ԋg*�(H�� BU6C�	�?\(��a�S~X��@A.C�	*��!�@V0d���`���B�I�U�)@Ň��	Lp�vȓ�9�B�I1@uz�'��"Q4���2%5�B�	�@'6i�@I�x��D�3	~bC��+�A"Wk��r���Rf*>o��C䉢)_���5��"Z�
=S6`N�)!"C�I .<)��8d^�<���+`B�IZ+�p꧊�8Zk�)�%ЩX�B�)� �#�_t���@�k^�[T����"OT*b����ʉ0?,|"�"OP��ÒGV�d�Q�Q#�`�"OPQsc!ߗD��-�4�
�H��"OƁ���_��`۵�V�k2zL�"O��J!�ƛL��б4-؆Q��qJ�"O�Tp���q9|z��"�$$��"Odd(p@�C��	�!��aI����"O|����Y�w��E��JK�_2���"OV�XE�ЧleP�k��L��"Of��Č�� �4>ؖ"O��:B,l��aEQn�!��"OH 9��P�L>�s��Ǟi�Ya"O�	�2A����b$_�+�A4"O�豦�S�f��F�߈�0�""Oj@�0��--��A�ĝ�]*xQ�C"O
�Bwa�8���Fd�� >:�	�"O�C@,�Vǰd0f�ת>^ȫR"O�xS�ϊ��0�Gʅ�Q4�1�"O�ի�-�E(<z�iL���`�"Oj�2D�P5�X�(��,	|�Ya"O�LK6Bڢ��%��f�7xfd��"OV�)Ac�p8n�! M(G_�=&"O�A�	1ypQ�0�"L�u�V"O8�+6��2K�����B+<�:`"O֐i�H�[�艇�F/@�k"O
L�$K!y���4NT.~��Ô"O2�O�
+l����MQ�?E�W8�y�oߙ���#�FPXXs�L߇�y��B�s�.E�뙞|��IJ �T�y����o"0c��R�g�qx�*ͦ�y2_�\"�t �$6)��A;�*-�y�QI�����
x�j��)@��y"D����`�`L�Q3��U��y��d¬Z��X����ͩ�y"�H[m�ZAB�)Q=ԝ��F�yB(ͲN� �cԂ�zp5iɂ��y2�[#��b�]�s�:�)����y���3j("���@�m`-�q���yҀ�O@\[U�B!k�8�ҡgE��yB��%��q�Coj�)�h��y�ᛢFU��"�Q	z�t��\1�y��u�n p&�L6jf|hxt�Q��y�O�
��qE*F#^<(1�g��y����s���c��=]P���t(�1�yr�ߜY�$L�aGE t�;�g��y���rPl%Ҧ��o- � �D�yr
�e��y�"C��֞Y�gf ��y/Uشl*d\1\[�����y��G�]�y��S�TT�ATJѕ�y"ʎo�����ϤE0�a��(�y�'Ȭ}OU��-�Al�` O��y�MQ��1�HSҐ��$�2�y���L5���ꒂG
�I��ջ�y��7c�F�k�g�9ʾ�8s�O��y���03��[%��?;,��I��yr���/�D�wf�����,���y����Ytxpa�E�j��z�l�!�y���z��M��o��iP���y��L7q�:8� f�4w�$I@�Ï�y���^���P��7o��tG��y"e� �� "EC�`���D�ʩ�y�ʎ�s��4K!��]��ݪS�N��y"��i)�z�K��%@t�r�0�y
� �Tf�<U�8����/��"O�1Q�暡nz4,���4�rT��"O^r���]�x<�wN����t"O���wؓM�:Q�HI����"O(����#�t����	�&"O��Vk�ъ�ÆBB�E�h���"O���Ĭm�ʕRR�T�sxZ���"Od�KQ��nV��4ʁ�"ָ��"O��x`o����i�\e�"O`���3SP5��햄!8�	�u"O�h�$� e@	4��,�4yg"O�Qc�5;�Y[W��dъ�"Of�sQ���2��ū�".|M��"O<���
D>~�� b �^�6(��Ӕ"OB��7-�;s��5� �H(��"Oy���Z�$��yE瀯U`0�"O6Pւ�`L��_�F�ؗ"O�@3ƌ�(D �#r�j��jp"O
Q`G������hXq��"O�QPUE	ܐȳF�_h���"OR8h'�Gޢ�aClӌF^Hc�"O~���%׫mJ����u�0q�T"O��r���|K.͈�DQ(]@���"O^�ǋmS�-x�#�-YK�T��"OR�s���P�"���HJ|E��"O�X����F�&�@:|���2F"Olm�L�5P����I�_�
eX1"O�0x ݳyhB����![j���"Oи�QU�q|���a�~z��"O\��ϳx�,��թ��>n�h��"O�(��N�9�R��o�*
F��9�"O4�p�I
W����G�I����"O�(���Ϙ�T)vA�Si�P�"Of���m��G����

ajeX"O�X���~Dh���zR����"O�ŚԍD6v��{�D�%f��yR�Z�d�����gA�"�UiB�I��y�DD�m��`�Ű��1!I�yR ��~��SeK7*K���0"Ͽ�y��U��9�3E�>V�(��d��y�`�x���8!J�갑t�Z �y�(�w!�ڂ��V� r�F�'�yi6/�8A�*L���OR��yE�#�1��>�~����Py2ŌO� �!��5Wpd�Ҧ�D�<Q�kO "�<Ѱ�D�6N�uhd��B�I.oj�0�g��&�|=鐠׷�C��3Ơ�j�K&%� 8��ˬi�!�d��Doܒ`�5���C�@��!�:{'P5����$
L\��vg��O�!�$Z.S1�4���,a/�Ȳ�˖�!���:���j��S2�ƕ���u�!�DC�W[d<`7l�j����aۦ�!�DXt�   ��   �  �  B  �  ,  �7  xB  8M  �W  �b  �j  �u  �  �  h�  ��  ?�  ��  ӥ  *�  s�  ��  ��  D�  ��  ��  �  K�  ��  ��  ��   �  $ � � ! n$ �+ �2 	9 K? �@  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
  yG�O�,�!�Oz��dI0v[>��˄,` ��
�Z!��\�, ��:��+Q��*�h�~2!���
U�>$�H܀��� �T�Q� D�4�"Zpx��:���{�:�y��C~v��g�M�+ג�7h��y猬g�<����!](�!D���y"��)[Y����Ʌ1B�����e���y2L� ����M9�,��0�Ƌ�yR�[�)� 3���91�80�g�Q��yM�c�!·( 2=rݙ�F6�p<A��N�]��l�7�
9Lr:��͊]F!�d�S�@Ɂ��D�.7��H�!� Y!�� �2S�7o(̡1�aכER�@R"O줳uHq_h��e��	g�|���'��(0��S<$°�dw�8��(�$���^	��m���%��I��?��6�6�`� �r�yX��[�P�dJ*D�XzP�J ,�RF״i�$�q�$D�y���x�4}�6���(B�F!D�TC����2��T�أQ\���3D�@����&޸��4/U3X�%�F�1D��"K�U�����9X_t���2�O��d��C]2qҌ��B2���8_l͖'ў�|B�E�%;��� @�k�N���e��t�?q��=$��\F�_I��㴎K�<�"��#%�g��Q���IK����?��L��6���B�X���h���A�<�d��"S�ԩ�l˒'ԭ���s�<��$�=�`1�Ч5-䰚t��kh<�և� `Q�,�hG'�ص[�L	(c������7_p��cqN/}�*<��{�l������y"��H �C܅t"�4
3$J�D	<QH�NV�~��
����+�iB�.ɐ(kb�����OY�E���~T.�X�$P�PЖ�x���t�<��	��؈���)��P;�L�<t�R�HRm8A��k�Jk�C�<�4�SF���:��ݾY����U�J@~R�MC���6�[R��,P���2�nϻ+�hl��"Oz�C��$o��<JvH�!,i�"O�Dz���0+�2u�v�<KO.�����G{��d�'�`�4�"�\}�p5���'����C��8|6��+wm�-�l���'���2j��Je\p�3c�)1� s�'��US嫍9V��X4�L!<\0�
�'g1iBI��-��){ ���iP�{�'�h�����Y���ʗ�Vg|�h�'6p=�&��8���a��Z,.���'i,���%*����G�WRH\�ȓ-Z>����6�6��FjP*x��ȓnM�dj� �
�vlR�J�(��ȓ>Ј|p�G���	�D盂9��y�ȓoh�$��GS�)]}�ŢXl����`m�:�)V�L��MP0�x��ȓ`���t��^~Xyv�n3}�ȓ~zB�Cc�^�m(h��bQ�o�Ɛ�ȓ0����uL��.�FK��m��Y���M��k[!�lB�o�!-�$�p�&ST�<f,�1D\�r�b[7s������0=a���pY�X�N^e̩ ,
�y2�}r@X�#@��|A(�.���y¨Ԣ5��%9���>�R�Q��y��3"�B��u���>���ؠ�yr��YL�3̬��!jfH��yN\:i>@��� v���� �yB.M�r�1�s	X�y_Z��/H�y�"�m0E�T�J,jqf-��y�O�##��(���\)��4f��y���V��m)���ai�d����y��*'Ơ�s�Y�
x�uり����0�O�1��%O�fj����\!	j*ܛ�"O��B���0�����R� h��g"O*|�5�S�;±��K��R(��0�S�Ix�h���'e��\SLG$q�!��Շe�L���U���q�3Ø}H�OR���OR]u˕ǂ=��}�Z�IՐ>i����Db�4Y���;ӜD��"��\>�*�:D�� �7��(x8�H��AS_� �"�	T�'���PI '�V�7� R��=6�FC��$vZ�B�i	�i�A`?Rn�MP�'h��O>�$�R���iѷ1��0+�#V�\t^��s�W��Q���>�S��� �
#�Z�PL����1��%ACeZ��LG{��)�H�H2Ec��'��k@�Ѱz��O���:�ɦ��O�
����N-�B�0 ͞?uK2���'�*�f�ۅ<�f)J΂�7%�+!�n�Jc�D8Q�<��ĔP-
1
B���k�P�.�l�<�%M�����pт �cO�ğ�	ɦY��&0<X{ �;�YZ�I��Fy �?�����Z))T,�7�2�c0gT �!��W�i��:��˿$���!'��O�1O.�O�}r�f��P���`�!�l�f`�t�<!��K� �ĸ����:��,��ry�̂��O�"<)���]�@A�q�׀t�|9����p����']�M��3]4�����/0��'lў�}*'of��{�_U�DyX&@�b�<��V�+�dI@�T�e�\1�$�X�<q4)O�pa8đcOK�0$��Q�<邦zQ�6c֌>�f(w��K�<!�&_ʘ�����1 ]b�<�R�H4po�%#p�M�-��3�oE`�<�׃��=����Ӻ)h<�j4f�[�'@ў�'z�P���`�U��F��N�py�ȓjs`�2���zbv�gXG���zKd�	�n-�f��"О�.dE��iQ>��(��쐸�&��� �)(D���ի�6q�J�5ꀋD�v@�'?!���S:c�<�#��&J����LT�PC��5|��HF%Q�8&C�3X&&C�	������H�>t��	S�̔�C�I2E&�)
bNA5m�t���hD�}!�T�%	X��*G�� �_&���"OF���\�5�b�n)~0aSf"O +f$�%�ȁ� _c.���"O�L 4�R�74�5���PHD�<j�"O�9�f��dT��F-�V%��b�"O(L"2f��Kt��R׌�g�y� "O��Kշ`��QcS�aO襁�"ON���@�'�l�a�8	B��)�"OV�
d�N�.`�4CfU1?f�5"O�];�J�8���+�=2l+�"O��".���Y��13)��ð"O�9#�V�U��ŉ�
ۀy	P#�"O4�1&׉"�V<�GiG�i�|%��"OD5�t��V����i �S/\Őg"O���G7c�ݫ�
���"OB%�vEQ�@q<aÆ�F�
��d"O���B��}$��@�dБ��K�"O�@�`aE�1�Dx�B�H
Ɓ�"O�,i�hD�@���ōF<�x��"O9C�#̣Uf2�"� w����"Oj�S���~���D<�ic"O��t�H��t,�1�P�IR"O�T '�3x@v��Ŗ�.�n�R�"Oj� � Sl���j�Y�D��mk�"O&Y��ѻ>@`rC��;���2�"O ��Dۺ*.�wՐ|��"OȽ8#˝�}\�X;u�ߺ#N�I1e"O�����E7 nܝ� �Ң`�@m�p"O��21�úf3�غpMw <��"O8�R���y�dD�C�äM@�`�"Ot5�'�G�7�$�"="�,��"O� |�C�E�*c�|��P5l
�2�"O6D�b�[!�����W"c�uj�"Op�Sƫ�H|.,(�$} �X�#"O<]S���;g���G�Ӌ���T"O܈%�2)b����&�.u �(���'�'"��'�B�'IB�'b�'e��c��y��I�gV�H4 �#�'
��'x"�'�"�'���'��'V�@JE�+5S:�x��
�cRҌل�'�R�'<�'"�'Z��'J�'��{Bj�	@  m�C��&r� �A��'���'N�'d"�':��'���'�JU��jӨk���Z���#|�[G�'��'��'�b�'�B�' ��'���qj��I��)R��;#킾�?����?���?���?����?���?)7�"oD�A:0>>�S��<�?����?Q���?y��?����?���?)ѢY�cLR�+��\����?����?����?���?���?���?��i�	1�>i��v��(#�@&�?���?���?i��?����?y��?���"�ЀF�$ZNp�቉0�?i��?y���?���?���?���?q |�*T��	kČ` �4�?9��?I���?��?Y��?A��?I�L��	��Y*�&^%P��8s!E�#�?a��?����?Y���?���?!��?�m��`5�X��gI�q2�u�����?���?����?Y���?	�.3�F�'M�gE�~��2�Q�nܦ�Å�B���?�.O1��ɪ�M�� �:[�D�Y׏R2O��`�v�ڥa��'*&7m:�i>�ɀ�M#a��HL��Gˆo�:���$rכV�'�hX�R�i!��+&�%��C6h��'(^&�:�K�(.�NБ�	�U�H��<�����8�'H�"7M�%���aË u}Vɀ��i�F䨋y��KѦ�]`LչE��-*J�RF&�]yR��ٴZ���6O��S�'la앃ٴ�ybk�9��L{�_�.�^��^�va�TH怨!�V�[�H}���4�n��L�7�Z�! �R.r �el]�e��<iH>aĶi�rՂ�y���U֨]�ٽk�@I5G��U��O�i�'�7-B�����߅F��Q�T���Lo�y��	�R���-o9��y#�"5��c>(�W㺃��'��hh�O?�:�KS�X�a����_�h�'���9O,�3뜁q�౱ �U�J�K�2O�El06G����v�4��	)b�1zԾe��EX!M�B�?Oo��M��u�-{ش���_!Ѳ�J��j!��*�a@�l��N˺���	�O<�d�<�'�?Q��?���?iGlX;"=�Q+�nD�+�&��΁��P����/�����	ҟ�&?��f:n��!y{�j�LOf���Ox�n���M+��'��O����O*�#�<�� [L��x3E�t��F\fy��4ξ��W�<q��'�"�'�l%��#��Azܪ��Ͷe⼢��'�'{b����P�l��4q���J���$GG�,*�����W����i���ɼ�Ms�i,t7�@{<vPa��)q2��$�΍uO9��Gv����O$ܘ��Z@DzHì�<9��7k�9wܜ��;#x����P���O���O����O��d-��N[$��G�Ҟ2b��BjΈV���ɷ�M��M_�6�"�y�V>m&�,"7�2o���ī��?��Yh@�ȡ�Mc�Q�Xzڴ0=���O:�}
#��yb�'��-�焆�ׂ���=K~Eb���� ��N��'������I��!'�QX�F�IB�uYe�N�I�l��ȟ��'a7mړ9�@���O��$�|ҐH��*/t�G솸5I��rW��f~b��>q�iښ7��˟�'>A�Ӑ(4��� 8ugre�-Lh刂�V=<�Ƞjg�TPy��O��jݙRX�'s���L�,!.P$�������'�2�'�����O����M�7BF���p�)=Q�q����"���Qo�F�';џ8I۴|��X1�f�,,���J��/P�I�D�i��6m� �X�2�2Or��כM��r���*0h�z%,e�� S7{nv̂2���+rEΓ�?����?����?���?������ >��!EH�=��UX��R�c-܁m1�牘�M�����'��9�<%[ū�H�P�SF�Jq�������U8�4R��&em��4���)�~�Xd.D/==�d^��$HѤhW	X(42�(
���Q���!��"U�t�O��D�Ov���O�	���P�A(DDarH) �����OV�D�O����<Y$�i2����'՚6��O>�[��	$q%��a�E�?Z�\3B�#�G؛�i�D(m�����ʡ3�~p	�Mښj�Q[�DP�d1��O��i',EN=>I(҂�<��'~��D!Y��y���D#��
N�p4\���?����?����?a��9��S̏�]֌U3C�,��XpU�O�to��j ��I3�M�'�hO��3�/')�lpjc�G!T�20&>O�Uoڕ�M�`�i��ئ��	�yb�Z[Aڧ�,MHƩ�&�<0kL􋇭�*y@:IPE`ŁZ
�Q��ʓ�?����?����?���(��H�Q�	1�x�k��ԛ
z�dB*O �nZ+l��\��ҟ��IJ�s��Dh\3h[�|CB�]�x�� ɵ�F���Sݦ�a�4(������Ov�TDW�s���x�U/I��#\ 1�)v�IK ��ѽ,;��%���'�`k@��}P9BM�=Ww�)�'U2�'������T�l+۴B ���I�΍!&�il9[aNks���>
����L}�&{�,1mڢ�M�l�]Q���$Y� �nU!V�ӌX�2	aş�<�*W`Ud̉c��^W޸r���_8����� �욑�n*������ Op�覡�O��d�O����O��$�O��?��T(���te
���6�@�v�a���ش�?	��i�����|b�����MS���,QR)Z�
��7��w}r�d�,�o��?���-od�I՟L⦃�_��E��+^'�<�:�2� �WХy7��'��'��'T�'Ȭ���!�X�Zd���V�j����G�'YrX��:�4*ր�����?����	%m�\���L�1�޽8QnQ	@�����dĦ��4x����OCL����G$p����6k���2�T0:D�{旯`���?�6P7��z�1����U��)�O����bgI/m����O����O���<)иi�Y��l !+r���`;1C�c)��yb�g��D(�h����&r����a�*C>��Z1��6����SG����I����c��� ��My"�ɁL����l�h��g <�y��')R�'HB�'|��'��V>Y��I�E�	 6��W������M��H��<Ig�isb���U>��~p؉�'�[�@3��C�mG�F�]��41��Jp��ק�4�O��4$��8�#�'ԾY�'� �4hrTI��eY��'E��(��;{�8�X&�|�U���	���0ՂƳHmH��eg�J��d
f̟��	ڟ<��ay��p�@���O���O����}���Ï�}�V%r���O��O>��'�6m��q����D�>��+��B:a𼰁���>J��$�O�s+ſV���+�K�<�'eɖ���ү�?)`a�LiBM; ,��41��߬�?����?���?!����On1g��T.$�)�Cga$GNN�r�DPƦ�
3hf�k��|����oz(�C���_���ī~������!��4u���LǚI��|3�'�ҏ�$��-B'��=�^���Y�c*��Q�L.IW�aD�|B\�T�Iן\�I៨�	���2�L��4`=Pe��w9���cy�w�ƽ�3��O���O���Lb���3��%�l�P�� /Ţ��'ժ7͞ئy���ħ��'��u#���6\�D�8&���X�JǱ_C)O�GI�ü� ��
%��c�B;BԫqM�|� 8����t�`��K��| ��gk��2�5E�0⪠bE�0<O�b��_�f�F��qF�=A��Ka�d�5u*Du;���?ƪ����΂i����W�M�(]�� ϹkZ7�͇ &p�f��>^&��� �~O�,�"��\��=B&%£_v��@��^�j��$jN
�(��C8(8�ehȓwM\�Qu�_��� ����V��l�GXb���g�>��Yw-�
�D$2����#PK_�\��'#	�v�޿�ē�?�N>)��?�Th���?��<;���CMP�]�q�L�4^���'�'���'bo ,���'�Ǒ�R;@)��-��5G�۲,� �6M�O��O�d�ODD׽	��'Dj=b��X�j�t��D�D�D��4�?���?��=p��j,�������
�}[�;vjI�H�2yB�T�c��'��'p��B�Լ����I��L�Z�f��&�I��\�P����'P�Q�5g"�'�"�'3�TW���1J��a���&Ƥ���ɝ.�X7��O�d�/�<�B$���6xFb®V'Q� �stDI��vhCD`�'��'[�$�'��X>���p�j� c�%S'줋1��!�M���a���<E��'��5�b��r���g� Y�V���z���$�O����@��D�OJ˧�?I�'X�	8�O���΁�_���{7EĒS
1Ol��m�S֟d�	�8��7L2]�ԨG+r�:��T/�M���%�����?�EZ?���k�I7L�x��!5V" 0
B��h�O�}	�_/��	՟`����X�'
l�C�ߩ4�bt:&aB���H��`ў��Ov���O.�Ot�f��%�d!W2q����T(;i�=�RG�x̓�?)���?/O�4�#Ė�|�%�A?/\��Jf��+����HX}��'��'D�	��0���Vx�O�|(%*��.�p���� ,�'"�'�P�1�M��ħ�-���K���Am�fB�K�i�R�|�R���5b3�Ӣaot�B�]��hѪPf���~7�Oh�d�<q�	��C��Oa���5�C�*yq�1���=LĄ��0�MS-O^��O������?7m�5UG���ˉ4u"i�WaS(���Z�؈"�R�M�Y?I���?���O��r�N-u�T ��ơ;�j�ˠ�i��'V��gW��'�&�܁�� �*�I�Dg�!3���Au�H�������I���	�?a�O<ͧXޜ�n��.��uIS�9��L�i��=�#P���	ȟ�3�IڟPkgI��P� �)w)�?:��8��F��M����?��7���ȧ�x�O/��'�BI
����B��]@�jY�/�V����>���?��a�}̓�?i���?AVh�k*�m�D�Ɂ!���
�/
(ӛF�'� =SX���|:���?+O��0	�6S��u`�O��8�����������h؆c����؟P�����	Z�$ɐ�Z8J2�kU�D�z$,��f�I,�M��?!��?	�Q?5�'Q�fбF��:�,-iA]�P�t5�'��Iʟx�Iq���'�
�`E$w��1�R�����y9�\$9g��#+Ʀ�������֟ �IAy�'��МOF�H�M��~Z��0d
��Qu�;�
�>���?����?��w�@-r2�it2�'��0��m�@�z&�	kJ��ps�o�X���O����<i�f�Χ��ɿi3"M
!#��mj&O��v|�6��Ox��O��$��>޶Inğ ������ӈH�L��b,�L��5C&�N�-��e�ڴ�?�(O(�d�:AO�)�O���|nZ�bKj}��#\˾��E�r\~6M�O���,�B�lܟ��՟H�S�?��	�ڀ J�Y0dP�8�(�3U��9v*-YsS�����I�����۟$���$�~:7�R�?M+��2%
�	��^ަeP�5�M����?����bq\��'�Ja�5 !V�&U{$�յ}���8�ok�"5Q�8O���<���'@"� ��RC�)�gS/2mr4�Km�.�d�O��$��'����'C�	��@��{.H�� 2��q�նBp��oZD�:��)Z���?y���Ii��D&V�e�'IbPM�d�i��	B
'K����$�O���?�1"�ջ�B,;j����VW�}�'�~�c�'2��'�R�'�2S���ā�7oOdX(���"���aG�0n�2��O��?�)O���OF�$[E������Y�}�����L����R8O��$�O|���O0�d�<��Gà ��I�9C�B�Q%ɖ�P����EUt���X� �	[y��'��'��ۙ'��E��%[n�-1��:8��%�f�Z�UZ9�d�OʓRlи�[?-�	rPQ��i�0&�d}��C�a�,ٴ�?�.Oh�D�O��ā�G���&}b�P�ax���W՗~8l�iI^��M���?�*OX𡵨p�d�'r��O����w���a��xȑ ��3Ԛ���>q��?���9�d@Γ�?Q(O���0vp6	A!.ĔTS�R��xx�6-�<�v��\��V�'y2�'
���>�;~)Z͡4KWU�i���C�D�]o�������	a�Ipܧr���j��O�[I<rD����Mo�i/���4�?1��?���-���Cy� L�t�E&�
 ����N�7A����O@ʓ��OK"��;7�t�q�ӹ�:�`e�hŀ8ߴ�?����?��7l�'�2�'���P��Ӓq	H��ǍI/m盆�|BB��yʟN���O��d�a����B�+Xm�F���Lo��Q%����'�^�,�i�1��m�,w�cM޻Cz��p4�sӴ�w;��O��$�O:�d�<�`��!٠ˠ /C�4Ҡ�ڙZ��)��x��'��|��'���w�H5B��מzA�	[�L�X��� t�'?��ͦ���Oy��W�^J�擼6*��PH�m=�a��7q5���?�����?���I�r����0D@�$�&�,D�D�X�y���s�T������kyN%q��� �� ��:NN� ��"�Z,���NѦA��M�ݟD�	�K�p�	J��O5t�p�N�dF�؉$f��F�'C�\�������'�?A�'�`����=b�,��dƼ_�ԪҞx�'�B��O�S�2ȅ��OO�^�^���v7�7�<١ǧj¹~����j���ز�.2.��؂gA�/؂���!|�����O0�*�2O4�O��>];��D<<�t��S�|N<xyc�~�t��S�Ѧ���ӟ����?(J<���7$�X�D"
7v|���J6$���i#P��'ɧ�l�d	\d����:e[��XZ��iR��tӘ���O���J5G�&�0��͟��9���M�Unj9sD�C�#���mB�	�jWp!�K|���?!�Oh��"ad��N9��cekJ�c)���۴�?qvh��	��'���'ɧ5/G��� ��<�n(A��S��d�P��d�<���?�J~b@�LȌ�����
xp6܊"��1\�����xb�'��|r�'�B�>ON����GQr���X4�3uQ"���'z�I͟��Iǟ�'g�99�Kr>�J�
�%��cb�&%���)��>Y���?QO>Q��?��F���~2O@	9���'�&���b�N�����O|�d�OH�
Ϡ�s��4BNB�ڍCtNk.��tb�KC6-�O�O���O �)�D�OB�'e�ڱ�5:������H^d<ɀ޴�?����$ȹs��$>��I�?�ڱ��Go9G�pF��U�@����?	�-n,|���S�c�Zu��2��R3e�Q���M�(O|e8W��a���d�D��
l�'�<Q)шL'Q���(n��[�T�Aڴ�?��JtP*���S�'h�
�9ЬR�Q�̈��aN�d���l�=$�����4�?���?�'b��O��e埆2�=y�N�e@����#D����%��G�d���B`T��ƍ�J8ּ )[P�$�{5!�$cw��E�� :�������M'�RW�sJ4|y�V�d�� BV���Rn�{b kn�A��zڰ�U�'�j�AN	�lt��97ޢI_lu$�O�
:^�)�K�yϸ���FP:[.��K�`ӐxL���٬Uw<�S��J�b���@�Ē�ۇB��F8���e�I�Y��a� ��w�h	� ��C*�z�)���0��Z���L,S�,-C� ��x0�stn��rɪ�@�2z���?A��?)�h�R`���?!�OZ
���Ovp�ԏ��(�P�(�@2H�,�w$�,q����Q�$̫�9a���<�d���Z�Ԩ^�u8��C��_gF��y���pe����"U2��e#�E:4�Ez��M8�?Y���:�:���&F��l�w��4h�����&�yO����@�l��5i�Y-f����+��q"S�L$9,��w��4
�\d̓MZ�6�'��I/b�]Ү����|��H�bv�Z%��E��83�n9|��a����?Y��eR$G�p� ��6VŰ��g�E�
1B��	k6�`1�8pj�EX ��&�<��琓\XZUQ2�� G�Y!Նځ&$M��eOoz ��+�
1M��H��wg���#3��O��$#��%��;"%ڤb�z�h��Q�7*���|�� @B��T�����CC�+Sڤ��,�O��&��z�mL� �Bh�#���]9W�~���E��M+��?�,�l��5��O����O� *0�
&Q(̴��ID��5��� �$��c� ��?�Z�!w.��hM�A��B�fF�b>�΅�(��!K���/5fz@ G�="+\h�a/ש3^�eS�K78E"�˫�H�2��w����_K\�]q���($��ЫL���'*�)�i#�$īS��MA"�ߺnM��yj���!��]I�e$�G>*-��'��b���d�����'&8�w9`�x��E�D�ĥ���'!�q��`T�'.r�'�REgݑ��ϟ|�gM�{*��y�F k2H(�f�J�_p> XVdߚ$.���%!�XǨ�ө"�>���ʨ[�4�ɴH�!`'�]B�B��_Gr��l�{�� 
�FU<aF �vԟF��7#����'���6^7Z���+$�b�'O����?���Ģ<q�,��j©�!k�����B�<QW�O)|%$���MM9}�tD��
����S��(�'�jTp%�`�6�;a�T�D\����)H��	��H�O�d�O���-�"���O����F�R��O�۲\�-�J=j��*]�^TZ�G�@� ��"l��!���I!]��T*��ʧP�\cՏš�z@cƎ��bx+#M�f����QhI��"R�	* �j�$��٣��8��CW�@:�F}�Ɖ7D��{F��	��5��*=>z<y��	4D��"v��&2�`-�f�A):���2Me����4��rp᣹i���'��6�ZU-��U���@(�_*��3��@�����#���$�<�O֍Ж/a¬�!j�7w�}���,,e�?����<��5:���+V{�taA�#ʓ�:��ɡ�H���0��Q��(i��g��P�"O:m�@�z;�颵�=mvxKw�' O�E��H �R��M"���Te�5p3O��E�����ߦi�If����C��'����:L��-��ƥ>�hy�rf�=*��K]�a �܂�Mۏ-5|�q�eD�|��j���w�ؑ�o�v�� �EV0G�����IO�����ƃ$?���A[�d�Diϋ��Ͽsp��.P�48�2� ��(��5�"��z�ɧ���T>WY��t���t�HY�0��5�y���w��9��T6Ā<�7�\)��'��K#��|Z�C�!�b%�4c5�ܙr��1a������?q!o�|�l��?���?!b���4��푱	 �@H��*����iG�,��Td��R��jSk]�vd�i�;?~)��y�̠z�Y���J�iV5�g�`���׬�%j��v#�6T�:�jA۟0���ʊ���'*��d��#F�\����B�K-L���'�1z��a{�K�2I�3��$'���G�U�xr�'rҕr��c*5@�*)j�pJ��"��|�I>1�5�&a_�]��YFŌ�ܭ(�"��'z�'@�1	��'0�1�RI@�ia�tjaE�KT���C�O�Nt��6D>�̱Ge�d�0�i�
vYQ��T#q�<��`-�&AT�[׎��:}.${`�ĒN;�PzB"A��h�@!����HWe�>�����	��M�i�'T�uP���t\��0 G�I�<1e� 'n��"2�W
z�L9#Y�D��)�lp- t,�%-�ȁHB���kt�(̓?8���|Rj!hr6-�O����|:6�P�O�F���� 1SJ�jq��=����?��p���p@V(}���bH�)<�㲅G�nb��vCɐ-v\ఒ��	aRˍ^�'�X�u�D�=�D�Q'�H�d	i��M��Mk�)�XH^� ����T*�N�(O*����'�Z#}:�_� z����ZW�@X@ZJ�<�E�͛W�x����B�h�c��a~��i>E�H<��#�5�(���9�,Y[v�[�<��1r>���'��[>=YrKޟ���(ianP�a�J��b�Z�t��7�5��U�Ik�S���d��5E�����@�l��,h�JZ���4"��4�S��?A ��5'(���P�^�8k�`v�(��XS�Wɧ����Z�j� z��O��X�@Ǣ�y�%�0R@t�%Dݠ2<�]/W��OEzʟTHxGȕ�3�x��A�Yh|����O���ЃHGr]H���ON���O(����t�4���BӰED9:��-44��3
ˉx[�ՃQD�"4�uk��v���&H^HV��'=������I$<�f���;=^�%� �$x��3fVv}��#����tǗ�+T���̞,C�Ʉ䠈p��J�*��W�Aa.���,�����O�'����꟬�'��-�����:A�	��(�'d�O�eGz"�O�,�x���c���((ě1�!�)aӜ�nZ� �ٴ�?q����/� ���	�ŦUr2d� Dmj�aVmE���@s�����Iן��	}�d}��̟��'3� �>j�:�p����}n�9����	(W>Z�"@�����#Sk�%�1���(ObJ�$�w�rh��`��/�%��.Ɯ.�у�?mmv��� R�9θp�L�&�(O}�@�'Zt6m��G��@�m�x+>�c�4�ȓL��Ѱ��2A��ᠵ�#^R>݆�	l�'�P����h���!A[�rdX�X�'�@6->��ϋe��l�����	J�D�� 	&���{B�16��>e���'���'�����g�-89�a!(�I�1�Um\�l���� ٱr�',Vބ3E	�3�"��@��.8�����$*&Č�bE���|��9�r�H�|HI�1�]h�X��U�>�Y1�)�I$�H�$5h��:����V�D;y��Eئ"O� ��@�P��`����A.��D,��|җ�x"$�'�h�ّĺh�\�鳁8�yb ���6��O
���|�s�K5�?���?Wi�.%����cK�	J�*��ȃy�H\s+V�.�<���	��\!��6�Tm���;A?���ƌ��d���ٖ6�Jh���Y��h�R'J9nR�pP�Iv?0E��lU����Y�K�<�U!�a�+,fD̉u�A&���	���S��?���@�$��-z6����Kj
B�)J�t�óo�'i4ը��½_c���	�HO���O4��Df�).�tS�F̩v���&�O����!sz�I����O �d�O
������Ӽ�%ϞIX4!��� �Z{Z��$@Л(?&8(�gS��|L:��͑�M{�O���+J̓o<�����*��R��P�ȘU�V�KBF����B2�x�!�Db�Z�4��s�H ��$��g����[,T�H��c��n���%�B�'R�ʧ���A@E��|�a�'B$'Vv�"LX	Z9�� K���#=ͧ��!|ᘂ�i��"NP�=Zl�� (/�J��$�'���'�B&J�K���'m�)�3 �dӖ�\�(����X�\ D%
������iu���E�Ń<�@�R��9l��֠��T�mb��~����- >#����`ƔI�dˏ�e���kB�6{dZ�%��KB��O��m�X��D� ��%f��t2��8i��B�I�%���)�7Qq����$[���d(ړI�d)�O�&t��EZ��p��A�V�|2g
�6��O����|�`��<i�<��֞l��m@�//R������?����A&h�=|��8h7�֖u��q��Z7h�P`B�C�/^���dV�cW����l�'mpc����z�֣R#&`h�b�7S8*����!?Ř�1E��?p�Z�y��j�'�Р���,đ>YA�P�:��ǒ�xC��q�$3D����K2ky�tk�>�~�qç1?َ�4�	&�0#�Dz0�ۗn>tsz`x�p�b��>�M���?�,�|�u��O*���Of97͏�Cn�T��&�,y�e��l�B�"xY�Dǌ
%~U��ǖ�,����OU1���@�~���2��1a#��G�� Z�hy�͗<�$�[�DF:� �h-��߅��kF3�ĭ肊[�8��`�U��f0��ӟ��䧃?�,O�� 3J�)���Q
��o[:q"O���?b��gݼV��`A���HO��l��̸S �!C����&)8��SWџ<��mR��8!Ɲ�����ݟ<�I��u��'o�*�*n��h��� J��b͗h��`C��� �X�Q��#l>>Ĉ�OL���2�N����G���n�8���a�Rqr��h�s�g��(�Q@�g�?�Dz���"݀]9���0���:���~rl��?q5�'��N��J�ԁ�B�5!�x5�
�'>�ٻ�a�6X�m��(݂ ��D�L%��|�H>���E�ԛ&�W��M��k�Y��2������'���'�b�ڀ�'�b?��@S/��ư%�������z����j>1n�91���y��M��y���
�(OP!Wh�"!�2Pق�N"J�v�{�`:l?K�;��~�(m���J蚢e��Xv���E��%bFb�{�,�1���!��<�!�$��9����mٴ#eR`�RBΫp�!�$������G�Ҵ;�f�:�-��@�Q&�J0���M����?,��!5�&\�	(�K�:��59�L7��D�O��d�d��q�tA?�Y�IӋ�T��O�<x�HԴZrb��cP7B�Ў��[�<�	�ؼp�L���+#w��.��p�SϜ�_�����ծ	�%Gy�OP��?�F��$�Nib�A#f}��Kǯ@xY~C䉰v+��p��"S��|�t!5>v��TX�I�&�ȱ�CϞ1�r�H^?{�t�� Z��۴�?	���I�"R���O��Oe[Ń��z�Đa�Β3C`W�6㲍�`_�qi�L1R�D��x꧶�Ͽ����nArG�ۀr@�X��o����,Sf�)vƘ�p�I�匟&$ԥ�}�ݍO>�������e2��Q-0����C���<E���f۷����捛  ¹b
��ȓA���k%��3Q&��0��8((�Fx��:��|�֬Ѳᢋ�A-���^�8_8�J���?ae��E,\E���?���?������4�9P�K�@,�亦��7.�X�� *S\��x$A�]*d��kH�=��)-ғ7�r�����>�^Ոpĉ�o�����h"<'b(��hX?!�h�%�GcZ����
@w�t��	EN�r�ÑT��D�<N,r�5lO��+�����Af��>�E�
�'��X�d,ڹ\�P���C�(y�H�*c$7��|:N>��`�PG��l*o�D0b��M06��ykwaՕT���'22�'��5hu�'�"5�d�
��[�F�� R	�В8�',ܫ54��(��B �����B��?��%�@@���-� 4Ă$��jR,5��:"Pz9:$��1j�8e�^h�'�@��ě�bO3n����6�P��|��r���y½����N�og���s�����1��5*f%@�E45�B��!W�]���Γ[���|2A�6-�O��d�|�&k�s4�0���ͬvF�C'�)6ƒ0b���?i��93<)C`�+AR���c��qfFI)��1�L����@d�Xt�N
(����7�^O�'D0E��mM�S�T��Gͮjd&S��L8dI�2'��9 �;f�l��q��I�'`v���q&�>A�2�͵D*<���	�<-�1B D���i2�PE�z�[dm<�O�($�������ĘK5F���TX�Jn����I�?�M���?�)��t�a��O>��OJ�@���ʑ��o�:F�,�V��sV� 1i���le���m�1�I�"��c>�N�)LK�5�CF75���cG��Le���w�S	D��R"�%@MB=���0{*���@,����B��]�9�^�!r>\8�J��w}�=��=��S��?�eAJ�<z��6s���[�O�R�<���M�AG��Dd�/*`|ţ���P�'d"=ͧ�?A�hԖ?_�,�t��*P!f-�׊ʅ�?���.Ԋ�Z@%��?���?i��[ ��O󮔪E�|���)]�`(�b��>hA�=�CFhCN4�5�80�X�֟��1��Θ'�h`s�B��&����69⹲,�,�j@@�J�(}���ä�0���O�n��Q�<��>�fX)���rv(�&��Y?�v�J؟D�ۓC��5 ��N�tw ��'���t�%����(S��:J$HD�a�F��	��i>-'��3"@:�M#&J��t�8ej�6��M)����?���?���<tzXq���?q�O�4�����?q����0QE��/�����%�R8�@�@ž<)aJJ�%��� �f��6�্�V8�8�$�OP�n�5�����9we�|x�/.�B�I�+��
5.[�"���5耚9��B�I��ĩDlܛ)�����]�d�#��'�=�aim�����O��'s�"�(�[!x������P�4��Q�roI	�?����?ɣ��Hy",�O̰k����:�q�Ē  �)P1���KҶ����:tbL}GyR"٬2 N�Q 	�?y��up�Ɩ'O������2�H���V�3W�(�ɘ9,d.�Dy2f��?	��S@Q���ߒL�B���Z%W�LB�IX&.����j[�Īe)t��hO�E�	�)�H,`��װ]��"��V$^�ɪn�rQ�ݴ�?������3hsH�d�O���W��5y� ��aq�5�)�AIZI��(W0j�E�R�]��eH�c�9�R� #&(���iQ'��N�*�[��J��L�&�Q�B^�ᓷ�F(a`�C#�P�_WX�(�E�Oq��c3:���5�P�:�"�����>(P0��'��O?���%c�����eX>푁 R!�N<�*��O
.Sd����[��1O��$�i���T�'f���t*RᲣNVi0c�'��͇;������'l�'/b��i�i!"m'�Z��5mªe��)�u���(`
Ti�6,�DkѻkG��S�g�"��U�$�	��}��g��Q�)P��!1� ��i\~}�6m ?=�����?a�$�#fm1O�07$X�JQ2�A����O&���'����D��Y��a�"��j	�Px7��u�!���O� �wA˲?�,u��h��~��]#�g�m�����|ŗ=-K�6M�?��Q���O�Ɇ�J4.����Of�$�Oԕ2��O��dj>	�E�Q)9�D���*z���5�8P^�4��g���(�k���cK+�Q���M�=GH���H�)7��!��ǃx���q�Ӑ;�J̫!%F�fԤ<r�ӿ)�Q�໒j�O:�o��kҨ����>�����{"C�	����I� �#$�:��j0���-�u&Xz3�$j� s�,ե0 ̡�H�V�|ҭ�X�6��O��D�|���G�MH(�N˪P��� �ܯA�ʤ����?	��M;�K�q5̩�شE���馧�"o��)8�͛�Fjp#�o 9TQ)E�N��(Ob���t>�̚Ս� D=ֵP����Q���?h��X��lڿ7�6�y$mG	l��D��&��Gl���&�'+$>��#��(}jr���'&�ꑄ�n�2ӈ[�c��j��[!%?`��'�ў���n7�US�.]�bBL���4ȼ(Γu)nlP1�i���'��S {.I�	˟��	! ��I2�@�rը��t��OU$P:��=SlH�Tz/hA���e�D��'�@�jR@��m��=a�'�=X@6�0��aTI���@�|"�B^������F�������ьe� Y�kҀ6�d4�p�'�O?�D�+
�j�=T�B,:&*(X9!�d�pZp�$�R�����@��쳍��?�3�#OWĠc �J9D�ji+q�[�������8�)�����	��8����u��yw�ʼ[DʅY��F�ʡ���~"����>Ir�C	v��A���sV�q��z?y��Ix�� ���E@} �
1E5-���O���C�'%���D�Bn$e#Q� ��z� � G�u�!����X�h$H�GD��* tEB�s��Dz����l�2�o� [�&�`�	SH|5�q��3f��	����I����U�[ ���|���\�������(iDx$��*�ƨ���*t�1+eF��v��(��L�����<��H�*��f�J�H�������(=�F�S�s�~)0��U~����ޮ]��<��O^ӟ� �4r�,#R���4��Y����8��L�� �0�y*L�Z�p�HI=pС��IR�'X�{� ��,���̛�y_JLA�'��6->��HSJ�Ym������[�$�M)H�i��"�������TjN2��0�'"��'Y�Y��"$<b ��u�̋���BؕZ:�@�#J�978`�0�?j���ߞ��(O�(�1��\p�d�J4�Ѐ>�D1�I4^�z����iy�+ZU���<i�	\��`ʎ�)��;r� ���N"��+�m	@�!�ā=#��HS��`�n0K��##���m����l&��R W�@����v�xK[�Y��$�-��HmZ̟���i�섚b0�'���h�d!A�\/Qf"��k[Av���H�	' l%;6�ϡ+�|��r#�X���0��w����!�*xߊԘ�J�8�P�k�wx�����p���!X{hTlʁ��ܦy�}�#�E�5NHM����A}�4� Y՟��<E���u|)C�\�"r�Aᔅ�x#�Ʌ�QzY� &�-&u]���V�r��<��b����XC�f��*�!�eΟ"�a:�����T�m����a�Z�p����`�I��u'��y��؃!\��hw-�k8&�pe���D�����p�P\ȅȑe�HHj�O����u̓=D��ŭS�
*t�3f��6x�0��f�j�:Y��"��T�������s�$/WN�c��KRF0M=��e��:0zN�u���t�1�O����	� 1�3F)�mGia��SZ>C����,�`o ���E�D:�Z4'�HO�)0�ę�t�8Yl��")2%˰

�s� ��K��G��������	�h�W����I�|�@͏�}��*�ƞ�X�������b�
D�Ո�n��m�W}6��
�2���Gy��'^0Ј2��2v� �ұx�$Р%�I7��DQ��g��*dm��iH�1@+ "�'@��4�6�� :��4e��'Vl��vꖓ�y�l�-x���˞Up|��
ѻ�0<���d�.�x���I6%{f�8�o��d����&�끈��M���?�*���p�ƈ�k�:�ꡭA)Nk�8� k�*l����O���H9�>H��Ō]��7M�`�<�X3'ڃ;p���Bٲ,����
}�`!� �(�)�T���R�j�8�ʖ�MǸ!ٓ�.-��c�G	iW��LT)�Y P�F F��M>�F�0����T7�=���L��U�5)W�K!��aך�3�ع��`sv���K9�Ip���D�$�ջP����KY3q���x)'J�Dз]к1oZٟ���a�d'.Gd��'�� ¼bD�E�r-��g��C���<�pJ"��D�P�Ɲ.�B�aІN'R0P��a��w�-� d J�na� Խ2�����?$�����X�Xm�Q�p��5:�ʑ��i�q��G���,9h$L�=Q��e�/~
�Ƞ�'v6�O?��ͩ5�0#r��1��'ĚkG!�D�~�������Y�,�y���'61O ��A���4�'MLq�jM�O�|u��O.
��k�'����|������'@��'1� o݁�i����O^0��S�+E�!��G���d�h��%v`ŐQDS�	}T�N�����d��TPz���
 W����h-fPx�c
[���	�n%����@��M%6��c������	��P�&�,k8v�{��
˟��P.�����؟��<I����O^K4��Oݒ4:�
Z7_E!�$�O�'%>�2-(G��=�"��e#A�����'��ɈK��D�ߴi���`�O��i��GOR`���?���?��c��?q����ԍ��+;H�Q�O�FL`���U2�-� ��N̥�ߴPcxc �;d��A��r�@b���k��L�ү��n���j�rvƽj�O;��� �+5=����R02�>�O���'\<6-O{�4��MB;rg.��D&݀	Q!��@�x��jK]Ib�уB�FHax��IPt`�ˈ�v"�����z�6扸�M[H>��c̜z2��'O�T>m�˘�vǐ��Z"():���e3���������	|7�8��Q'B��pn�]5����͆�	�R�L�.Hc��heIՕG��5X��Z�'� p��ǳqC2a&��a��Y!��v�vt+W&X Q��}#��,)=re��iU�F^�aV�|��U��?!D�ӗK$��A���J vy�qeM4:b~C�ɯ`�Y��7�ZA�e�12(��hO��`�I�!��DR� ޭ&A,�p�ȥkJ��ɰ^�F�bڴ�?I���iA� ���O��dE�H��$��0@_�o8(�36`�'�v�,�|Fx�K�+�&p�B��#�P��Q�܏s�ڠ�i��p�3oK%)�(���O\���E����b�`Y�ʅ���PH�)��� ��f��:SK")c��)}��a�"O��@���]��5AІ	�(� �R��ɟ�HO�i�OV�q4L��j, "����a�$�O���E#Q�Y�m�OB�D�Oz�DM̺C�Ӽ�  U�*� ��̠1�ސ���M(!g�!ȃ�N3w��4�����M�Om2�Ҥ��h�l�b ����-V)�eY1 ���%��:�P���T�z2T�*�A�fjt����b�$R�ڵ(H�X�P�4@�+��X�@��O28��I�A��k��P�4R��;[tC����u���N���B���pՒj�a���HO�i>���("�ԄnZ�v:̡�ވL1�š	8z#��	ߟt�	��0�Ǒ����Iϟ4��a	W��GKlMU**@2��P&�� ��L�cZ�`ɪ�a��:`�x���� �� �����j��B8c;\ӗ��8n�������H� ��)K��0b@$� Dd����MK ��B!��/�p��J	P��yb��iZ��'���'Vb�'�O{
Wc%bA	T"1 �F��C��0<���C�UD�9��o	=3?�$Rq@^�I���X��ߴ��'���'k�'N��`F�Nj�	�1@@�dxp��'�֐�7H@a��^�Z �a
K�<�R�0d�>��#ꎊ+��b6�~�<A��2Y5*P�y#��bTJ"O.e�6�o!�0Ђ%��ݲQ"O�I	�R�T���T@�Nz��B�"O(�)���Q
R��w�ɯ7l��3"O�E(�o�`�X�6	��|�ҝ�"O<IKF�ݿ &�sG�nD!�"O�#���Xw���P�h�t�
�"O�E�#��<${�I߶w���q"O��`G�IF���r�U�F��Q��"O�!yf��,��M������E�3"O��	�ՎI��)�V�R�:�.}P�"O�h���k���$(��L��#"O��c�%#hH\���E$)B"O\ĈҮ�� =�t��P�$���"O�2Ҭ�(������/�LxZ1"O�Lxb��;��)����i�J-�"OV`h���:[dbP���8��x�!"O�p���I�H�Tܩ��^����
"O�]y!�I�T���w� ����"OB;���YN�	闥�zuH�"O��L͵�4���/mQb8�"Ot�VN��P��-xi��#K�1a$"O�Y��FM�Mq�hCT��i���"OT���)&	�T1�i�W���"Ox�s�/���5yG��Hv0� D"O|�8Q��P���5�.+g��C"O��wj�4�,����7II��[A"O�X�C��#��h��7><�1�"O|�h#�R(n�ά��J-�FL�����h���H�6*c@�� � 7�"=yD"O�EХ� %m|0�$ǃ\��8�WZ����)ʧ@v����$݀���A�ȓMa���2`���G�`�FQ�O�(�'6lO��Q�,QB2$qg/]6Jk&����'��lP�	�M�a\�_|���_�Q���i�L��Ɠ7� ij6I�
���2��@�N!��Fz�.�9H�4�"�5��O�V�[�,�tȸ�V�)�<���'Ri��V#w6�CWѯ`r
���4	���)g��6(
!�)O?7�+M����@J�E�@��,�&`t!���Du^L�Dʓ|���° ��cD��$V������e ��I�?	��c�b_#bӜٻVo.\W
����2p>��+�����@�¾+z���!C�2뺄��O�Pp"@�#W�U��lO������I*x�Qr$
X�C��T�~
5hI�"_�Yx���H��uZ$�v�<�4OV�2女AB�	{Ix��acW�
sd�*�f(DT쐲+O�O6���7}��X2W�'gZ��4�տ��xB.�(V0��*J8����E!TB��hp련��I�j/\@!,<�I�*��3� ^�����_�MA�k��FN`�Q�'��ݙ��� +�� Ыܛ5��Q �t���1�)D`���%P�X!B�>rMI���D۾&0���f�T�CF� �wd^"�'�}Cr�؜z���)�%&�P��d��=�r���B��rX`�%|ζ�ڧ�'RNm"W�	�8���[�nU�#���ēe6�ܨt�~j�Ծ���'�lREei��m�P�%˂a(<Y�A�~�~�����"C6X
��ԃA%Q�c�:�*�\'(u0����'������\ ��X��^�0*\\��	�7߬� �E�vw"6���<qe��U��!C%(A�~N2��c`�=WѦ�Y��
R���H���2Iv�)��^W �倓��*'��j. m�/�1�*u["��p�>)��.q��y7fH5E��hT/�{����ٰ7���č�����=L����,�={ ��rd�Ak`��mZ�S�$�c4n��Y�{�>	H��+�U6)�blz�(0�y�N~��H��޷Dᆥ�vȞ�`��%���4��|Ifh��QD���֝��r������!���G���;1,C^8������2N�T���ԐL�����W. �x�z�g:Y�4�t�ɻ#��(������X!�O(�#g��S�A��b�p#*_�k0�+W�>�0ND�TW4a�S���;*<��RD�s}J?aP���$͌����L[' Y�#M�<1&�V2r�l��`ɞ��y�(YS�'y����F�E��\����;<�z���P�m-l5Y��ۥ���~&��]�F��L·\BH���\��yұf��9A$}��(4LO�Ζ���i�M�Kt�'曇S���a�Е� I�A�)�'ze`��B*-�$�js���qP�R�U^�hs"AG�#􍙄��z,�1�t)ŏl��DjS�l:ΌZd�-q���VYt���b�dZ� $6�����e´5bx��bW> ��9Ua7fXЉ�'�@Iw��.L����RO�R��K>�'Q(�P�@��_���A5�� ͒y#�'���(Af�y��k���h@)C�􄊸m����Z+4�q!�d�d����Ԏ�o`��@'�4�����ʞ*a�!P�(�/r��#�[--�(��"��=������B'.���Qnĝ\��6M�RX��9��s��Ie���T�{�N�At�ʥ�:�O��"��*�R)P��=83���)��~͹$�&��O���%��A84��c�I84 +��i�EJ$I��5���Q���~���0N�dY�Fk�����H�%j]�<鰻i���t02�C!���OST����F"z�y�t}��:Ov1�KX�Fz�)�#)Ѥ�{�A�H��kED��<�EJ�g����H<y��4pl6p�\�wI
>br�I�K(g@�`sG�u؞��4g @�U�"/��Ѓg�8|�6�}�@�Yw�$��p:)S-�xy6Jƻqf��k�ΈW*�x�e�YoƘ���'�^��PL[���t�L��Lk�}C��L>��'Z2�c�>Yï� ���'3�0�:d"�O��e��rҘ�"^�Z�nܣV�>1�U�05*ܺ�'��@�$�ğ(��J�F��i���%a�6^�*��9O4Ț�_��~R����P$a����):���^�j�����.�p%�T�d� -V�bp�O�,�i�9� C�����.�x�J䉣B�#L�����(0�O�NVQQ,�q��`~��j�%T����s��=���4��/2ʉ�V+�5A
5��DS4{>e���V�0<Q��	�g�����M6z�Ί�GǢ�b�:f7
%��h�v]{(O��*�P�\yt$
k6`��i1���ra��\h��ƌvE\��R�IcތŠ�4?�󭞳\F���4��<�5���	�~���54@�xV�� ��� i����-P����[�yH
�{=|]E}�e ���(��g[T!P!,��#�&�6t�mAʦm�<9�'R�ʓ�y�&ƚ7��w�ˢ��}0u͘mb�{��@���=A��w� xjkO9L����I������OL�ϓ6����f1���H>�Gp�vЀR��d�tt�� ��'+����	��P$Ѣ�ÔE1�=[%� �h�]��K�� Y�S�)�6���g܊qP�i��C�������O�EM�Pd�v�4x�s+��w���O汁���̽m /�L�Tls>�"n�^�M�0W��p`2L��Q��`k��_~�l(��:8@\9��	�]�fH��I�:tQ�%Sd�J�=p�6�,	>:P��iIXϓ|�v�ķ>��}��\c,��VF�
g� ���H�'d(:��'��r��Xx����B�*`JYA��O�d Y�f������U�nb��+1�O�<���OTP9�'���:al�'@0�!��l�uu�,��䔑 �����O��o�8ml��ӄS!c�xhFM+e,D-{��ɜ�M����2��nڶ{�8$�X�V��YZՉ�
elνS4
�cO�H�7k�\y�F�hH�<�'�|����4%@Æ\
q�s�ҿi�<pb�GC2@�l�áX�L�ɟ������wv��Zt&S��Bh�S�5��\�4����ெK���iHI�dհ����(U{$(ӣ#�&A��Zv<����",OJ�V���u0�͓� �@�P6l老nL%��ˍ{�O�b: Yh���1��*S�ԺXW��*�A)䀹tQZ�'%�ĸ��FW��I�$<� ��yS��/A�N�t��'XUH�a5O��P��E�<�Q�?F���{_w�eէ�'(�|H�A�q��a�㕐Ep��'�ԉm��^[��*h��}J˟h�P6 N�0L��	��-��)��(`�E�$-��OC47m�٦y�`"
80�(HIa�Ob&�݂��'π�kXGx�ii$.���bB&O��i\G��hk &�Z�dC$G�6�~ZL|�&�S�d�F��1�ߵz�X���G�,�:4K�g8]��\�#�'���J�2���L?k�p��U�!���(�+�?���'zP��H>�3?9�!ȦaB�E8�W�<`�	_;_E��V$ҙ-�(��	S8x��(�Op��'Evxذ�d
8o���O(����e˖�i`��`�z���këg�F8�.�6P�l��U˚���ę4��� c���Vd���œ���}�Փ?t�a��Q�~I�:�yB?O�;���$N0�A�ų��`���	U��)�h�u8�<Bc�-6��R���"��R���C�'jq���E#I5�T#CC����"H�~/Z5�ش*�`i�	�Ӽ�U��8ǬE�����p�Y�l�y������zSV�r �Y!R�@A��DL�Ą㉴'H� EL	S�0�����5��ǌ�\� �ĩQ�h}���D@1Od����D�w��B
U�g΁=J��]���6�x���e��
�'��:�����8�CA� 8x�}��=P�:��A�C6 7���������,�n�1��Q�aBr��A���l�a�m_�u9�+��/&�u���Z� ��I�3<��f��<�I�!N99P@�;v6�����i���ꄳC��ac�'x�N\	@y�b�yb�Ha��0]�ax��#� 1�$�SC�3i(!(����^ �TEM{�'��KGQ���4��
I�j���ݴ`Q��h�� 	�F��X�ɬ�MC(�b̓M4�Γ}@�9a�	��A�)�E� ��$��C�,k^�U�/��$�]�dX�֠��2gx���! ���)Dr��b��;�`K���<��'�v-ÒNM�y Z9!� Pn�'����e@�P�jq��9$Y��[���`��s5,O�Q1�2O�)�ҧ�7�p`��Be�tQH���2j��|ad G!6�ay�$g�I� Q�|�Њ���=I88�����>�RB�'��G1 ���ǈ�\o�W�]7R� R���<�xwH�
o���ӫh���V��p��=X��9[�@��5O=��oڷ�M��'-�uO��m hm�!U�9�q�S��Pà��r)<Z�Ot� ҆�:F�\�I%�a��8�u�?�ɢ�y�-��v�8��N��v���B�OtZbhjf��y�
xd B�u|X��,�BW3�qP�U�oj��I���'�X	�O>q�"��<٧�R-E�q���F
c�´��=�.Ԅ�	�}�V�]�k��ԀsØ�N�h��NY:2�R�I-x��(�H<is�Av~NX%i��I�'Z��ZdD2�h���I܃o�d%���d��@�n���d�����"��,6 `�7GT2q�f5@�
�O<� e�>i�*"|ф�	$l�H"��L~��ӺDf4�Y7B,N����Jմ�0<1��ݚQB`�r��/*�<S�aM�Cp=�!��|G~"��.Xxri;`	�#Y���b��쀁/�V�h;u��EH�*3 R�@x �#?�Qn f$��D �'-'�a�@i}��~ҍ���4�����`L����� 72]����]cDd�i�� �n'l
���%F�Ć����P}��~�Ӻ�f,��	�y�d�C%�1����p)ì)'�C�	�9tdQ2�M��P;-�#ժTi���O�h
����}���HP�j-���`+?A��|ҏC-L荪S/ �!)e*��0<qDgD��re��&��Zчs�칉�`%n�\��KП?�z��ˎ��6P���'�B���9kM~�0˝]�y8M�� �';�$�th�<e�'&�a�O?���!��=P��H��?�TY�UC4D�<��I"Qwrh[Ao�;�b�iBI2D�h�b^��$"�k�uzˑ�1D�����ѢN��) �л�,ш7�$D�����2ME6�۶�=���AF!D��GoѬ@��2 �=D��ta)D�|`1ƿx֐�s��]�$D�'�(T�L�eV0
՘��&zܨ�'"O~�a�WsW�#sb�C�L�2S"OP��K�TB��H5ǌ�b_�;�"OƝ�Î�c��c��A�8U���"O�+D1i��g.��3H�"O��sM,�B��j�H��`"O�HaW��/W,}´���j�"L9`"O�,@�#E�\z!���ي'����P"OL�k�%�."��as�.<xu"OX9s�LY�X �\%G;&[�"On�3w��G�r���PZ�N� �"O� VD ��֠R�R����"�䤓�"O"��D��j��x'���o�A�"O~Ց�*��d���f� 'r@$(�"Op���ӊ8��I�7��,��"O��S�)Gt�A��҄?�i�"O.�󫘹'�q#r �'8,�h�"Ozh@w��P��dѳ��(q�J�Jw"O�\Æ�� K?�0�e/�J��@&"O����U)�6��V�9@	���"O�|(�ڑ6o6$	Ŏ�h�\ H"O.�{��̶t�h�nZ�1���a"Oְ�G@�%��">+,Ѐ�"OJ0ja�2����РfD��"Ol��e�W8eP�����"O�T���(�=؃ ��\�8���"O�0���I&(�L8�Po3
=��"O D��b�Y��q�L�j	�c"OjUsd�28�
��!䋐v��l�D"O��it�ԪJ�.m1v� q��Y"O0��WDe��v�ӶI�R��s"O�a�CC�>[b����ڲݺ��g"O���'Ӳw���E"Ӽu>��T"O�eq��Pk�He�ס�#ne�]�'"O�[��ǰ�DIHAW	kW�l��"O��2A�H�jE��� �-h��7"O~���J\�;sl{�hZ2�r�p�"O,�b�I�S�d��>ڂ�"�"O<рb-�XҲ�Ʌ$�g����"O2H�c�db�"Ǣ|K��j�"O:��f���f��#'؛ ����"O��h̑�;&J8�q&���H�V"OD��#-	>b�|�F��M�@���"O�@���ȣ<�
��Se+�2Պr"O���%`����B�a���!"O��`G t�����a�.pT"O�(��F�1�=
&l��>�����"O�����oy���t�G 5��a��"Or����e������H"P�y7"O~���@��^�̙#d�������"O.!Iek�;�R a�,N���C"O�*��R*1����&�$ ��{6"O���:He@��$#Rq�i+"O�*�*]������ITt �"O(���O�4����!X�$B��q�"Oh<r �L&([T@gW0h�\I��"O� q7��L����@�SXP�4�y"���j���G�T���C��y"J��+��UБ�,!�"\(�y��_�{k�U ����3�4�R�(�y҆U$J�t����-*����ϔ�y��ia���j��aRM1L��ͱ�'{v�+��# r01�d��/�U�'r@=���9*��$��# G��B
�'w<���Ə��61c
X�j�"��	�'S��02��0�𬨁BX�L��	�'�1j�\XaM��ܜA��c	�'%&�k$� �|9�-B��A3(	��'������b���`�
u�:��'I8is���-6&��q�Xhخ���'�v@���K�nz���WSm�x�'~���$I�%k̰TAލ�`�
�'�z�&��i�Vm[�'S�G6���'��IRc��%N���C9N�!�'��H�H��6J�`	��u�E��� ,	�Af�V8���V��2�"O��BJٔ�vpXGm@�|4��3"O���΁3��Xwk]�8��"O Đ�L�< =^�bO'hl���|��'�.	��W���'��,�Z
�'�AKF ��*�IUN��*p�R�'E(�@�KR~ۂx�K±5�ܢ�{"�2�S�S%(icQ/�$�0���,X�@7fB��a�x|�又�up��u�ӱ`B�ɑ��i��읈6K.�3�`Ԛ�4B�	,��u	�$�2�" 1�o�v��C�~�p��+
��1��u��C�I�W���˗&�$N,ڕ���R#B��C�I=f��p�oO�]���P�Q3-"�C�IB$�G�A��~T���T�;	&C�I FlUk��O��^D3����IB�)���3���t��:�노X��$z�@.D�d���C����`b��M�t�R�!D� q���<�1�g�(����!>�Oh�	R?��葃,� $�3霂b\�<��g��G{���i����0F�=E��|+ �ǜKB:@b
�'$$���&���O��r��i��'O0H('�@�x��A+����A���{�'�@19C�\�cՄ�!�\>( ��'=�h�E�թ��\���ȈQ�݁�' �Y2aT36�.�[�LU#��*�'L�D��N>j�.���'; ��'��1��?9�R��Q�φaP��
�'��-a.I�i���
!c��Zk4��	�'�H�Ǒ!�%"C�P/���+�S��:��)
�Ɣ�$A/:��@��iA@B�:$���6hȀ'm&����P5rB�I�8��d"�ą� �
1+�8���<��c�a��p;w%��Q������b��!�O��{��B�l��BA"c[��ڱ�'���/u�QPѦW"f �Q��2u�!�d[����
�: +F:Y��Oʓ�Mۏ��
0�#NC�`���Y&��<}�j�a"O��w�J�g�ɨqn�"Ө ��
Vy��O�)�3}r*Nt�$�����S��JGe���y�ϑv�L҃l�&]����(�y���8& ��Q��O"y����Kڰ�y2�Z�8�L,E�,
���y���C#�U�R������I��0>�L>��F��y�.�z5iM�N�T���p�<�`�O�}a����1>f����Ak�<I��8��*�E�k��Ԫ�lIi�<��IȾS=4����
�?՜��Cʈz�<�B��R��@z M�(�r�[�l�\쓣hO�OQ�y�E��I���2T핑b� ��
�'v,�95iNl� �k�dk	 I;
�'�}c�+��CP�U3pJ�����
�'��H��#��tQ����%A=аy
�'2D���#�?�F8��̂�.�A
�'[�܁�M�;#o����Ɓ �E	�'1�Y���)Y(	Ĝ��E��' ����{:����f�1(
�'=T�� A$uXٱ�"$�V 2	�����2�$)�@�GI˂���#D��� X�*�V�q�X� ?V�K i<D��[��@�H�H�$A�i,��&D��r�˝%Gn0Q��I5d�`t��!#��蟮�B��%�v��r.���"ON��4�K.�$I �<#$2�2�"O� �2P�\�,��iC�
��;\�A�"OVx��BW�{��Sw�ц?����"O8�YO-�-�W`M6U� �"O�Za���!�z�!šE��M��"O|�"b��Mv�|IP�Y�c��4S"O��"t��0aM`�C���(u����"Oܸ+#JY=^�q"�+����"Or�C��Y�j���Q��X��"O��B�9NX��B'hA�S`�
"OJ��tk��ef�U�#�S�����"ONu��ȍ&px���%ˣ:% �3s"O
�0��7Fb8)6o��(�Z"O�A�Yp����@�]�Q���'�L�	Yn��W�Q�s��͸�J�#6FC��^&� �nA�%Ƥ�Q�O�-[L*7�*�S���<��O��G��$�f��M�QUby��"OР�Y�/~B��Wl�MA�)���O�"<ɍ��M�YYBA�s&O$y�2�G9^!�d@� B����Ș"x#��M�x0�������;��?�&��a�L�-2���Th�i�h�Q�7򓯨�֙�2������0����3���P�"O�xh�U��=�S�}d2)�$��>��	��1��`p�(�
N<IT��8Q�
O��C�/V�~����CNTp"�x��'%jٲӧ�L�Հ	{����y"Maܱ��M�cn���+9И'�{�1tP���R�C�g��D(c�шO��IL�O�4PR� Q�D�Y�@�� �Lh��'?�0��L5o8�!��.J*�РH<�����7EF��RW�v���f@=+!�D[v����6��;*�1R�2$yT7-3��;�ҧ(�e#��ȿ���z� D�iD�:f��<��a�'N8��r��?D���(���Q����@�E,>�	Y���O����=D���S&aW�2��q�'�  Rf\�o3,Y� .&�	�N<����IϫYl����;����"�!�$��w�� �MɢB�
�q/�!�T�,���Ϙ��d����f�!�$׳M 씁�c[�#d�����ۤf�!�9'�]�� �^��Ѐ�$!�D�j�~��$߆`���8�/�r�qO������KXiȠ�<���� �Z��!�dL������{�R]�4K/P�9�	�'A�9kЂ[�%b�L��c�/�`��'�d�H4��4&�`�$aS�D���K
�'�q���R&��@@�Q�7D�����xB�L-��}Xcaō,`pT@�,��yR��J��a;���W�HɫD��yr�X���+�=M�H	�G�1�y�'�(��L�#��s�й*1,Y�y��E�;$Ƞ���0@���y���_�
�G���I�C��yg��(����؉}�
�c���yR�%	v���u\����́�y��*e"�z� �'[�L8C ���y�@:���W�բ�FA@R��y� Q�-Ф����٪�{��ˠ�yE0sc ��t�ޕ
gJ�(1d�"�y��8�>���Q��+p%S(�y�b5nې��dA�E�f|�VN�+�y�	>5��� Q�/f�B��ۊ�y�ő�~�5IB&ŀ+����E	�yR�H-;�Q�g���"Ypqf͗�y
� ��X��>5��d�T�ƍ.�=��"O��s�1Vcb�6b�?-�ܘ��"O� �c\�_��} 듶 9�Q��"O �EL�5��a�ȡ"�`a"Oa#@iZ:.�ތ�!����{�"O�Pt���v�i�l���-�T"O�����'�Ԭy�"$W�ܹ�"O(��0K�5PB�I$g�I�b$��"O6L���+?%~e���	�V�H\�q"O�5!T�W=<;�D�=O ���"O 0#B�5�=2�hQ�B3&�R "O�C!�A-SBi��63����r"O$)��̇((8�y3K��]FTY��"O�X�r'U'D���AGg�p�0"O������2OH8�����0kД��"OJ����J� ���U��3Ob)P�"O�� �k�4v|��󬝴`;��P"O��K��1B����T0�tq�"O@s�Ćj�� ��'�h��0�"Oʩ4%[�f:BE�E�/-ی�ҳ"O(��AD�d�h�� ��9&��3�"O�!!�`S�z&P(�"�Ξ�Z�!�"OjI�(Ҿ^Jr��$ʮ\x�xt"O��
D5":tqq�I�Ug� �"OF�9��	����L�0V`1�r"O���;9�X���YegJy0�"O�\��\�:Om�@�_>`�-)�"OV	S�j�#� !a(��!wX���"O!�N��q���Y#h�l�9r`"O���KB���L�e@U'V0�2"Ob��#D�4Q~Tx�P�	>��Y� "O�����P�@pnd8g�F715�t�f"Ox`ʳ/Y�y�|�(EA8	�{�"O<9����l���TA���*�h"O$H���)GR�X)�a\�8-��"O�0��FY�l`�S���D\��hA"O�6��y�Ô���d �f"O<l�燖�v�p��eÎ�'�@9�t"O�(�L�=/�R���Şn��m2�"O��� Ѵ��q�� �0�ԅ�"O�@`���n_\���IRwl��"O��85I�8sD�ݸA�,rn.���"O�J%l�_�$əp&OP�Ҵ��"O��B��Ǎ5ܨ�B�H�3ǨLhb"O���(E�D��CڥX_DQ��"O� G��m��t�!ʴ�  �"O���'� �r02��!��9�d"OxEI�ۍgѲ�#q�+R��	k�"O�����;5u�]RAl0�2���"O�Ta�.ڀG-���E"}��l�b"O:J���b%���O�:L̀�"O��I�/E�g&@�`�TӜP� "O~Y���0�91#��q�T]�"O���/ߐx�P/Y��)�@�y�$ �:�l)�@l��S[�m�V��yr�ЬAB����	�_jɪ�K���y�ց6�4�r���0X"�Xp
(�yb��>N ���CY�H���3c��%�y�	��y�7 ,2s,�h�d��y2 �'Njb 0��[0*�XÄ���y��*�d�pq��%,Įm�o�+�y"��5�����2���X�d�/�y��E�B����۪2�2E�3�Ӆ�yR>0�q�WhC
,��i��E��y
� �X���TH@����(��s#"O�Y���:[.��W�ʆM���"Olx#�C���1�*A�tn�1'"O��
6�=P���ۊ-�̈��"O�e�u�`���W��~����"O�r�O�b�"��B�OM�l���"OLX""R�R�Q&H^�Y��@`"O����$>��[��Yu��$��"O�PS�5���:e<Ҽ���"OD���Ʌ_f��PF:&��#"O~���J�-Q�Z`ĂƜV��S"O��aT)@��7ˍ�T�H-D���!�?�l �V.Mh�H%�"
-D��� A�E��zF����� D��q���4H��Ae��Hi0�� C=D��
dm(^Z��G�T�0��uf'D���PÉ�@}��#�XP <b�;D�L�`�=q*,L�T�-Rg���1M3D��"�z��HH�9��Z"�/D��SԠ��[�E��'J� ��]H+:D�h+RI[����=�X���"D���t P�6�$���]�<i�H D��`s �Rf��RG[��͉��?D�$��/�'��Q������I#D��)q�3��m�h �pf�5D�t�r�W�6	0O'I�����3D�D"��Q<h����*T� �G 0D�pk� ���xm���$����9D��kf�8%�����cK�\�X��u+6D�L����9� I�. ���1D���qO�bA���B�]E"���#/D�@õg��'v^AFF�AϪX�3�*D����N/6CV��5��&@~б`��)D�Ȉ����!:��\�|��{��%D���ǽ,H|14�ۍZ��xw"D��{#�9 Hp�H�c��bN��J#F>D��	�k�'5�豘`D�
A)���<D�P �'P�g�%9���#S���z�D4D��@���  �����9^f)Z��1D�d�"��"\cJeˇ;���Ӕ�9D���`��89,p��A䒸U��K��6D�p��OF�4�}�����4p��[3h3D�\@d�� P�	R��ɨ��,D�\�f�-��I1.ΎNv��!�,D��*e� 3|є`��/�+L`�8PA�)D��`�E�2�����j�2a��`&D�,�҂�!7k$@� �>�"��YC�	
o�ň4#��H�0LRc�
'|^B��/wt����"b��%���\�kCjC�7��t�ѥ�1AŖMcT$H�4C�4��x�&I*A��`�Ve EC�	�j���;�gU�l�l����c�B�I?{��\�g!]=.%:|�c�B'�6C�	@L�I3GԿrҥ�N�X=TC�	�t,:�J�BB�Ct�k1�!�|B�I=Р�q�Z�s����!��!D^B�I>Z�l��ŕ.?��d`�3��C��#d�<�Q��)B�ԁ��)$B�	:���Tf�	F7Ĝ"(�!j�!��U>	��f �<���X�K�!��e��sĬ���1@
kF!�$���"��Q��hۄ��!��!q]�u�sJ��@����FN_�~�!�D_+b����"O�zw�ȢW-��!�� ��Zsh�?Y" ��cN�]�`̓�"Os���Y����@L$p����A"O���!�	`�H`�e�9� uZS"O4dj���2I�D32�8�2h�"O���P���Bx�vZs�8�"O2"0�V9,���bЀÊ\�=�"O�����8I"� �D޹V��P"O�q�J@:(�Y`��!A:4B�"O@����L\<訇�ɗQ�bp�"OtpSAH��c�V��Ԯ�M'�1�d"O �b�b�VP 0@ϿTt5ʡ"O��ak�;]�p�V/<D%�P�"O��`�]�x ��UF?�1D"Of�EK>}�Nu�#��|���"O�}B�m���*q�� h�L=��"O��M�6:�8�֥�?��xU"O�e���'��5�Q�S��}��"O�e,�Q�l��#R���j"O�kt��uS<D"QcM4Ae�8b�"O`YP	%E_"�5蒙W:���"Ou���H��Na���G�=@�!K�"O̬�U�N�;*@���L-tdRv"O�=Ɖ�o*����y78���"O�QC‿�\�b����p
�"O|�Z%
G�k��h�W݇�`�"O�<�ō�O��y�լ�-
��,��"O6���*Ʊ[Z�T�p��f��� D"O�,r�$ˑu�P�Qs�
 �P��"O��aC	o�4��bE�e4��t"OJU��JN*۔��D�"tN(B�'���$�ec4x���!K�q‪O��!�C�Yi*���ʁ7b-��g��"2�!�H :�`%�ݺMu�$�%��z�!�X�X^ԽJ��B�-�1O���!��@��.�*Qx��Ӂ;�!���@�!�����ecr�j�'R�
�!�$ŁK0P��O�7FƕBs��*	~�y"�']1O*�"$A^j����H�(u ��I�"Oxp�����r�ؤ�H��D�{�"O$шA�2m �uBSg0�ܡ3"Ou����{�)b掆���5"O ̘3�B�E�:,Ӳg"�V���"Ort(�!��-g�S
�gz>��5"O�AHs*�$fw�@Yc*��H�(��"O��A�o�Ov=i2������"OM(�d"Kk��pg-*ɢ}�@"O����+�^@����XKJx{�"O�蘡����EKI�I��r�"OԴ �U�ei��Sd��C�\K�"OP�J1�@?[M��qa��k��L��"O�H˰H�"S҈�2'M"e�0�4�'L1O�A�w������8%��< ``�P"OX�r##� 5f������q@�M�t"O��%��mN<��So�>%V��a"O�BׄC�(�܄�l9y),�!�TF�\qhWkɱm�Hp%S,o�!�$�<\K�C�'h�<dS��OQ!�ɝkTVͲ�"K:$�.�q��	M!��H�-��0hU ��~-
V@��85!�A��,�����z�x2o�L!��׻[�Iڥ�Z15�<%�D A!�Ę+f���!�J,��Kȥo�!��F
d�V�a%E�H���2�QI!�d�4��
�<?�*i���;!�� �9QV���(t��"G�	�<�E"Oh�=$�sh�,r&\D�5"O���B�""�1�G&B"�܅B�"Oĕ�S+S�\�d�ҥ��i��b�"OPY�a�iqn�CU�%L��
�"O�f��.[u("��82(�
0"OȁK��.�*<8���@��僢"Or}`�X&u9�Йv���S��I�"OV�9	?v��HT������c"O�QkV��1��a�)�X�6��"O�M0�n�! ���裋H��लu"O�9Q䎋L� ���pR%�e"O���#��$�q�E�O]�����"O��ӥD:W���P� <��U:�"O�Aӥ�.$�p�-��b������'^��	Hb���║!:�b��<9!��$oƔ10���\�BF�\'N!��2^W�ݑ�!ڕiK����w!��64u�����(���H�C@!�d��j'	2m60aZ	 ��>!�׊-]���#Bts�� �k��}�!�dov��S'OIxL��i��~��B�k��иAc�:L" �e�(L
B�I?X����ˣl� ջ���%%dDB�I27�R�Ғ%�-'��xR�eʰ-�B��U�.׸:�􉄈"v�B�	�jI�9��AB1�v`:��SU�FB�ɓ�r�V��8V;8Ā��R]B�ɚ;*Q�q(�$?@dUhQl���eO��&*XA/x��(�+�ȋqC�OJC���p������7F���kʳtJ�C�I:�~���n�Z"����&�C�6���h&�܌{���;��+�B�	�t�0�x'm�>RҀy)C$W�B��?bh>�NP�A&�1����C�Ɍy'������N���Q�LҲ|[�C�I5(�\p+Ub�j
�!�1&��z]�B�ɍ1���; B�UZ�0�k�D�pB�	>h��BU�@<.̊��שR�YJB�I�gkl�C�N>��kS�L3!B�	�A�y��� k�u���߹_��C�ɋRD��+b�ܭ'��رC��:z�C��<� Yj��J���.�~�ȣ=IçKG\�%��.�Ɓ�T#E�#u�i�ȓe3>�;#b�cC�m��H*B��-��*3�|�&��+�v���,یd*4�ȓ �Δ���-R�])/�`M�ȓ*��L#�R"y�a��GȘ`m�X��J��1 ��$C�1��G/
� �ȓm�4�����"n<9��F(CE�Q�ȓ[�vq�C

.�6�P��}�ȓR�2�H'�%N�����a�;�4�ȓ؊YY��
�c��e�r�	P~�1������'�ɨP�, #�S�����lHNp��1	��� �X��h�����I���%�H�c���V���ȓx>�&��=�B�J�'>8j\��'�ў�|�J!�Zu�b!�:P5t�Sm�s�<�'�	jE2M���P:)<�ͣ��r�<	�*_q�T�
P4 �hCW��w�<y�n_�RYh̚Ve�.m��b �	]�<�� ��T*L�Q��^�U�z�B��]a�< `O���$h5B^�L��H�u�<�!hJ�2��IB��\�0V1��BDmy"�)�g�? b�a�CD�A��Q�%� <%J&��C"O�ɐ�� {v2��g�Y$��1S"O�I�s$:�"��e��F����"O��K�(�:M���@��Y-%ܖ���"O�R��!=�j`A���>��:�"OU t)�o5�,9���Ֆ��f"O����+���Ie&��wp$����'u�Od�҂���hh���$9G�-I� ��y#}�$�B��$�4�ҵ�.�yb&N�j��%-��e��y'���,t���ڨ�k�EY�y��MK	t��@S) g�%�ȓgElUqv��϶�LH�'�,�.,����<� ��jЙ�DRJx숡Üf�<�e
���X���8'���a�a�<��(��q�씺��Ͳ{��E���Y�<�c�!B�)�C��IB����T�<I'���@�A��Q�d�ŀ�S�<ifo� 5t�z��:C־1��M�<�S� �L��ك��9T��-����U�����;`4P�E*��l'���ȓ(�� '-L)70!w��:�u��U�<ؠՇG�"����b	�~���ȓe��Y�q"ׅ?f�C�͊kT�����Ұ�߭dy�kf<@�Bj)D��g�.��I�*dִ�eD(D��j�ЀQ,|���e�
�s�&D��bԔ��M�al9[�yQԎ(D�F��'9�hy)Uϔ9,��I(D��@v�3�����S2TY���S*&D�02�˄v��{��K|�3�(#D��`%��<�mb��_-D�N* �#D��"�_�tS��A߷XD��P�"D��{�C^	���a�'�-]�p
�� D��YAIQ������)��	
��3D�(��ɗ[�K��j<��o6D��J�JˡN��K�"*��-��4D��a�&�2������߶?[�=��� D���&�)��l�0M�,��AD�*D�(���;�&��'��9߰��(D����$v� 
�c��9���f'D�4��l�4�26�z�P�AւI�<�a�-b����d)�
0���!�}�<��"�Xrpx��@�?��S3�w�<I�L��C\1ir�ʽSo�9)a
�K�<����;}��́*TKYх��D�<���l�Z�곏C�"~������A�<A�� _����Ň�+4q��eG@�<�2�˜&��󀑃r..���ˉ|�<q�Λ�P\xC� If|�䧕b�<T���4�ȼ UC��~�� �Vd�<��,S8�r���G �|�S+�f�<�	���UK�;a�c���X�<��!1B0j�*��KxJnL���n�<D�����a�O�v^$9��ld�<��8 L�u �Ȉ� &�Y���L`�<�6��N�	�w�P>r��#a�@�<��(ԿG#���nֶ�k�]z�<��Ő
!�m4oS=3rj<rGi<D��s'ʍ�{4����C/zW:� ;D���w%@�@�s3�E�|��ą,D�P�w����d���%��d b)D��k� �w�TcF*h�N�I�H&D���"!��V�����h��ĉ9D��  �����+��(�_�]�
���"O<��6'S�V��:TK� ��"O�;�ݧ&��`�R+>�i�"O���֤��s(d�׫8$����"O4U����;M��:C��0c�<�4"Oz`2�,;�ȰJݢ`>*L r"O"�bcݎ9m8�Ӈ��wnr�"O�$�TIK�GÖ��g��rd�I�"O�5���$?��8#�Y��x	+r"O<�e���Pl�)s�^7	%v��"O�T1v�_v]��@�
;B���j�"O�+���5�r�� ��e�6��6"O8CRk,�H�[��O�6TAt"On�Z�)18��ypfoP:Zu��"Or!x�O�]M���+
�p�I
T"O8���cC"R6"D��	�+VPZ�K "O Ր�R&e4����)�)z�M�"OZE���3Ul�#�)�8v~\M��"OH�)u�Ih�D���&^B*"O� ����V�ȻR(�v!d�d"Op2�(ڃV���X�"�ٲ�"O��1g.qC�I p��._�PW"O\YB���\8���㋒wJ�T�R"O�Ivaã*���W�EP��Y�"OF	���i�PH���;dP�"OX- ��>l������6 ��!v"O���]�Y�l�q�T-�ЅA�"O�TU�K�6�uaƗ�[�p	��"OޔA�-í4��#Q%ҹvx�T�"O��H2cڭ��	�ÅI9-t�x;�"Ov��6.ū@2�z����4^XtH�"O	��/(/2��ta�Y$8��"O$��QEݜ=�(i֎�:	G��A�"O��J��G�$�M�	O���w"O����e�\d�"bmϾVk���"Ov�����������3NFY��"O"�*��W�0��iK+|�C�"OZ�k2E�w(P9�gL�r���"Ohh�!�L�s(8�����P	&��"O�ŚuGC['N��,� ��U;�"O�j�+��;��`�AJ%l�j�"OV����6��	`bԞ%삑�A"O���'��o�
(:����t��,`�"O��ZU����9fڦV�du!G"Ov�XVaR@�+�:7e4M�"O��㡪yBP��W?pP1"O�-C���`�@���ŀ�(j�"O8�#�ހMj�E�7ȃ�����p"O��߫jͶl��G˾���@"O���C!$؜�cd���a��"O�mї�	fv�C.V�8r�"O��y�J�I��X������5�d"Oҝ�!d�Sˠ���×��L�"O�XP�$�)r�8Ԩ��G78ِ��"OfEh��+Q���P˜���yr"O,a�T�H�_���ԈMI�� "O��Ef�>p�����:	�0"Oj(c5!	'��9%�̶v�Fu�A"O�y�D��4'���#��+*�؜KB"ON`�J �$~���3F�%�����"OP�9�FQ(D���Z�,�����"O�X���2mW�$X��R�Cq�u��"O�H�K	(4�Z��B%|p� �2"O��HPE�
�:�J��
�-U��2"O� �����A&G��Swڂ��T"O��!-��G�N�"�ꃻ"� y�"O�����c�V�+�o�/LLn��"On�#C�A�I~�:Ci�'׾��g"Od�˕M�Z��Ix�g� (��0"O�9���Ԛ�H< �!{0"O��AZ�z��eC DX�M���V"ÓF�X=/�j�ɒ�DȈQ��"O�]�̅�v4�w(^���,h"O�s�EY]��U�����"O�q�R	�Vy��#�^,QX.q)�"O��J �,��H�4;TI��g"O� a�ܽ>nj����|Ц)��"O�8P䦚�=m�RfHcNH;C"O�	�4�I�A� ��يH��I�"O���Pb̜n�jy��e�%�D*�"O̓!�Ĭ4tP@���ձ�:�q�"OF�AT�JP dqD�c.Ld"O �"i΁h�>5���܇��zR"O�I b����H�8D�\�X�b�!�"O�� �&�-#�d�R���I�6"O@9(�AY�+��	J�Lܡ~��4Y"OБ�!iIF<�8��G.(���"O*��j0<D�������G"Ol� 7iB U���.H�|�両6"O�5+U(�.�k��G<xp2�"O���A� *��@qM�*N��R"O5�C��vzJv��b4��i�"O��ZFA�2�ʡ��4)ȅY�"Od,���
_eȶ�K�2	�R�"O��č�q?�r�:PQԱ%"O����3��`�&Lॳ�"O���fO���)�7'��wD�-a@"Ohs�nW�4x�&AJ��"O,�)��5!���	�-l:����"O����0Ҙ�r��M1134��"O$�2C�̮?Ʊ�����3+����"Of���"o�+�$AФ�E���y�K� $c~�C��$�^IV���y��BVH�$��E�����#�yb�Q��L�	��W �yBf16��haH4Z��5������yrK^�� �d)�L.�R�%�y�%���l�J��a�w.T�y�]�{:f���2S_R����y���)8\\��дQX~��׭�y�́�[��h�#C�H��P�w� �y��;r��5�.T�3� }��ҁ�yr��= �E����+JT��%���y��9n�>8ib�! m�Ӆm��yB\��TU�F0��I����y��̷\a�81���8+���V
	��yD�,6 8%	k"1v��r���y�P9{��Y{��Ӌ0�:��s���yR"%p� ����[0n�
p'C��y2�͢W3�;�,CZ8���Ě��y�a�fkfK��H��j'/5�yr��|�����
�E��Px����y2�ƇA�ʍɗ��
�.y��&�y�7d��!��C9z���:�MO��y��/q���Z"
	�h��ܒ'Iе�y�J�76�않q#T�6T�S��)��<I���ܛ��qP�N�\���%���!��K�K6j Z�k�46�@���Fj�!�� ���%&�2����o 6)|,p "OR� C�ѽI�{ǮU�&TI�"OT�ö�_"҄�ʱ�ǈ,�1X"O�H`�Q��Q���2q�t�b�"O~mb�L�	oVܤ5J��;ؾ|���'�T��e;ZM����!�C��q&n/D��C&0N-2�Hv,�h���+D��kx�A bO�Lx�l(D���0KpX����.�j}cR�"D�X�7��	8b"$�/}���� D�Ѐ��ғt��D��4i�|�b?D��ӦיY\=c���n�XK%�8D��⠆�%R^h�hQ�O�hz�e�8D��[6cܲm�R]R�(7 �a���8D��V�A*f����k4ۤ*D� ٤�$Iq��{��M��� /&D�( T0'W�i�Ο�_���g�1D�dSe���q��c�(����,D����Ї?�HQjV+Ȫ$�����?D��YGh�e�1����8 �8A�;D��{@��&	�����E�lQ��Rw�:D�$��.ظo����k�N��ÀD9D�x(f�[�+NX�	e��<�:�Z��7D�P��r�x��惍_Wҹ"D�9D��ڶ��/�#w��-�Z�p�8D�$��C�1!d���)�8O�"y
�H4D���p�|K���(� Q.���%D��ۅ���\��`K56f$l��h"D��#�'�x�^0BF�!�dO�aNz�x��3�
��"ĵ
�!򤝧� ;qa���t�� 8�!��V6?����I5�@y�5�^�ne!��^=�Ի'.�?H��"U�{+!���R1Z$RWOV.TD2y[� J�!�dG����D3:��,I�"9:�' �\bc 	��a�AI�;�$�P�'<ؽ#r�îD��0�n�5\J��'fl���H�B�!�C$Mn���'?�5���q�<P�B����'�<�BE�
�:p��� O���'���3 ��
���qaU�z�̚�'��mj�'3A� ����z1ڨj�'ݦ��炖�N8|���ϴzBx��
�'��i���r�z�&� w*T p
�'�lP$	i��yT�R�����	�'$�@�E�bl�m��Ɩ�s�>=`
�'�J 92�ظa��-�b��,]�>Q��'��]0o���P>��A�'�Rբ��� 6����P�Щ18Y��'�Fm"2Ȗ
4�P�q��T�! �	�'	h�r��}`� ���fHa�'<��3&nR�	�%��lMb�'���sC�O���k��5��(8�'6�;u'�&r�m��	:|�Xuy�' � 1c���
*B#"lZM�
�'!(�[��0@�P8�v�ϼ&zU�	�'Z1y!!DZ�Vɳ���Ft��'����$CT,����i�� =TMA�'/��S�h�Fw�M15��)h4t�p�'����'�K�s	��t��2��C
�'~q`Bƅ�95Vl@���5,bTY�	�'-jl���x�jr�F���)[�'�jQC�e��Nς�Q�"��F\�
�'t�,��@��p�z�$`��&D�� )��ICΩ�ŝ��vm�C"O�@��T�L��=�@d_��<��"O������B6>��q�Q�n'���"O����f	X�� �/3P�:ɛ6"OĥP#��(e���b�5k���"Of5Ö��f�5yq�B���""O,���D�<;8��w���Č��t"O�C4�Ɇ7��ɳ�$��� "O����G"KkʰP��>v���"O���#oʁ2�xd��o�,`��j7"Ob���� ���+S.��
���!"O�ݪ��ژa�vH�&H�8�F"Oh,KE[=#\��u�P��H0�"O�Kf�ɽs�(-���V�إb"*Ox���"H�QJj��F=�R�"�'��x�#�-"��H���ז0%��
�'����ܱz t�[dcN�.1,���' �1�ǬR�X��,�T ���W��y"�)`đ����(/.�]`�\��yR@F�1|����H"%C4�����y�k�8,cV8Y!m�H�R��!�Z��yȕ�
(�j����;Uh�� $�;�y��Ւb� ��Љf��8Õ�ξ�yDҩD��t��'/L���/T��yr��$��� w��<+�9"l��y�"�8��)	�|`|P��%Ɲ6�B�IT�4�#G�B�z���r�� S��C�I���FO�ByzV�&hD�C�I,I�-���f��!B��C��K��Y���<����A��/_8�C�I�xQ�Q�tɅ�Rݦ�(����
��C�I
2�xX�W	�d�<��(r��C䉑i.�W ��zpB���j:pC�4v�0�0�I1?��b�n¤C��b;��H����X[�i�7�!�D.8���'�ֳ��)�`���7�!�$�7:\�LR�m[��Ԫ����!�@("��T�傸L �Eƨ9p!�űc�U��c��-P&P�GS!�d��'����e�>|�B������qO!�D����ly$�
<��!ܔw�!�������<�
���o���H�H ����K�g/�ط��y �>�"[q���Y�49r⇇�y���6<L.� h��Y�&]J�+�;�y҃zÂ�ӓ
]�Y�.]����yR
Y
(`lg��h3�a���y�	ţRʲ��W�K��u����y�M,~�4hD�Z�I3�Y�ᆒ�y��Y�$e�ŠA�6� $���7�y�'(X�А��F�6)���B��y"G.�<z'�-)�Ԙ�U�Q�yB��x��&��/��maU`��yb@�UkF�p<5�8����0�y�/�W-��)���*ƅ�¬�yҍ� ?���鱡ʭ]?�ma��y��\�dx,��	(P�Dha]��y�'�$J�����͂W�
�Tf�4�yb�W�<�}�B��r���y2��:�H�%�&����ӡ�yb"6� ����&'i����#�yRM�F�(�TE%�B�3d$^�yB*�A�a邬�#�0Tƀ�y�ȗGꐍ���ПC �*tF�y
� ĺ���Fĩ��ݒu�`}d"Oh��H�7�(e�NT�%M>q�#"O>	i�Jվ�R]����GF�Hk�"O
�Rbbg�� @օ�,g���Q"O�9E��#qJ���6ł�-��2u"O��Y6��|4�E�؆"�@�"O�@H��x�4<9L�w�^$�e"O�M �)����I�G�^v"OT�`e��$��y�JƜ6��	;�"O ,`1����T9�i��$x�"Od0����*�d��ݶR��`S"O�IkL�"����w��(`�Lz�"OFlz�7-�D@����$E�4Q"O0�$�@#7��U��c^�W�] �"O<Q���z��cbԬY/���e"O�̊���(�<��!�yH=8b"OBX�:J�b1�L��	a"O����#��	���B�' a��"OI�����\�n�i�`�p��9g"OL5�C�J.���"Af��E"O�@r%̓�k�D��$j�EHd"O2(C���!o�`���@�B͏��y�(Z�7'
�A��	�s�,��"`ǅ�yB��=`�䐨&.
�}�0��EH��y�jڻ.��%s��Czu�p��h���y���xMֽ�s��j�L��#�4�y��^c���[W-~�SBӺ�y��[��T��R`��(꒬M��y�cv};�j@�^d*�rI�.�y���v���!bl�#|��ǮY��yr�/5��)����Q�m-�y2 �)D`<��w$�VJ��b@^��y"�[��~aB��@�J�+�̌��v���h�&��� `"�ԆGO���ȓ���1D�^�y�u�p�\??��y���   ��P�2v��d�3��9��j<����� lX<�R�(���W,�X��C��yt�$^�n����J�aA��n%[b���w3%�ȓQr�y��
�;�	�4ɶ��7���w��aQ�Ģ5`U�=���ȓt��BW�J���y2`[,g����)�X	s@��T��5j�"P2%z�ȓ|��# �?�
�jSO�$Au�ȓ"���8֪Xt���{�EMY��]��SN�hs�F�3 mc����u�ȓ-NQ�B�0Q]H ��hH�*"~���)��C`Z��N�ʲ(Ա}x"��ȓB�HPb�Gԩ����ùu�(��H�$d�P�I�q��X�%�Ͼ��ȓl���i	�	<kt	��d��UP��U"�#1P�p����fZ���P�ȓA�h���cU���Tǎk�>���B� �6��=eGrM��ꈊFb���+��D���9�ؙ����<G�e�ȓ1Ɍ�1 �K�q�rĻ!��6FhA�ȓ_ʐ]+Bb	
�}��ω�_��L�ȓ_P�\	�CG^�4d�QKW�ITཆȓG��p�+O�&H��Abb�$�Za���2	[%�_�:钕�+X��5��
ƀ�*��W/[,������v��y��Y�f��8R�1BW����t�ȓs�l�fnS[���r��o��ąȓ*0(0ٰc��b��	� I��	$���S�? �Eh0�Ĉ>�H�9V,Y!(��i�"OD��CM�r�x�q�*0zn�+�"O@=)��C3ob����֡F�D�"O�E����n���w�Ɯd�Ɂ"O����+0D�A۵�Y�D�� C�"Of�ʥ���c&�{�e��Htnp{"O ��K��,�L�u��5wj6)��"O�%Q%Lc�-�r�E�VjXӓ"O:�j�%8 Y�l���ȋA���2#"OF��S���
��4iw%�#��yQ�"Ot)�b���L�Ĳ?���"Ob`E��/t�%s�	)�����"OhUp$_�:� �(�₭s�١�"O��bN�cf��ƠT�* 3�"OpyIիf��p�"��&z���d,D� ��7I6h�Y��&+D�`��P:�@Q	E��#r�U6*O����� ���yGϵ(Ժ�8"O*�@2�:�>�BeA>^���
w"O)�"P�#1��{2BK��<,��"O& �&R�5�6���4W��`b"O�|�S�e��t` H�9��"O�xx���:B}cd@U�ov��7"OVm�1E�N�$�׼[ �F"O�Y�0Z�.D�%bb)�6=��p�"O@ �A-�u��!x懘���a"O��e���hI
��͵1�t��"O���J_386ũqfY9A\��A�"O�qG�p�2��X�@J���D"O"p���9Z\ (�p�N�nG>E"OƽbOڐK��0���E8���5"O{'�%I��&^"w	v1�5"O:U*�	_�r0##ʆ ����g"O���2C�<��U���[�
��""OF����cH�iP�@ ��ı�0"OH����D�j� ����7�T�S`"OZ�Y���=N���nW���QAV"O -[���=]�9)R,عZ�n��1"O�)��H&c�����D�!}�⠊a"O�����6:��ؔb�!�

W"OB0c�K S�*���"�,b�Ȓ@"Oe��� !ٖ�"��e�č��"O��;j	<��qW.eQ���"O�XR��\�6 [ÎD�p2W"O `X���l�L�+��Ĩt>dH1s"O���������i����.Z$��"O�(�d� @,�/	�zd� �"O���_hEx�,-�ҙ2 L�_�!�X�Z����=#��v��
"!�$͋9��*�z$b Dҏ!��O{�.��u����f�
�i�A�!�Ă�p�W�"�J���TvR��ok���K	p�$��&��l���ȓLm�� س9�!�W��h��e�ȓ(�:mHT��K�
u��.�S����ȓeE���Lւw2� �4חB_������5ڒm� W�X"�k���p-�ȓ�.l�O�q>r�`��Xˠ��ȓs�,1eXAh���Da�Ąȓ~�TI@)A�Rj<�#@^yTȇȓpX��bG˗
m*D���$�TE��J�bq�Ά�WJ�H���8���ȓ"�ҨPV�fP�a#�AC�^ah��hV���B+r#R�Ȓ�Ѝs@���S�? ���M������s�zy�<�S"OF����b�T[�E�����@w"O~8��g����ᰂđ�WV�H��"O"dx!$�O:�I���V'V��h0"O�t&"?]�0���șE7���S"O�����%k��ƦJ���"OvU������@͔� �Dr"O��!"�{Z��Tj�9=�1��"Oy���\�����װ���*O�Ⱥ#��y�i�3A�h�|t��'B4z1IP�/�~X��e��e��Ai�'CRA� �- ؑ��Y�c�$p�
�'{�p��)cWde���	�S�F�)
�'�*}�5 �U[�P�/Q�$�	�'�8 ��P+|�z��V\N�>@��'z ���n�eL&�fm�M*|��'�Bi���;�ؓ& ��|qze��'Y�`��ĴJ�ʍB1��	n��]�'ݺ�
ca�	�����J}a�' D��0�B9g��`DO�H��H�'�&aj����`QX! d���m�0X��'Dh�s�+�~�H��&b�`)I	�'��+�/�(�{�UaU����'���wI�7u^,+�O1�(�h�'�� �)XЎ}Z/����Y��'6��0w�B�{#*�)�'��<�0Ř�_�L��FV)M���'�6H�7�@�*��,:�"��E�^(9�'/��YR�޺uv]��e�ğ=�'�@@�(Ի8�lL7��63��H�'fvEa5N�8Vء����#=�(\K�'�2l �f�r�5�Ǿ4���'�!�vCμ.`�j"�ĻyR�M1	�'�q:g'��X����`I�B�l�a�'����E+9�ha@EkӸ7�&Q�'��4��M����
���c�� �'ɚ�zpeִl, i@o[2��
�'y���Q��x��_"�*I��'��I���*y�-h�`ߗ�.���'L�(�E A�𸢤z6���'B��Q��c�F�[�	_�L��'�N�RB`�}3��9��;W��]��'�� ����"ܸA3�5T+ h�':8x��&�0�^��FR���
�'�]r�M�",iD���ҏ~A�}(�'�� +�� m��Y��c�}b�X �'�(��@�~�)��@�0*nl�"
�'�Фؔl^&4�2�G�����	�'� $��ѡ8�3���0�t���'�H��T�͞!�Z2�lF�Q�fՒ�':��)�IҪ8�I���F;���'���4��~��P�� �I9���'xYJկͭ���9���r�.���'K�c�]����ۓǛ�m�rT�
�'�=���� ."�� J�
r����'i0� �g�8w1� �'�
ɶѓ�'�@�( �Јy<!"ā�5,�,�
�'�0�Z�F��^�@��ڼ#�@	�
�'���"7+S	d/�ѳ��*�b��	�'�H��BGZ!��2�D>-��b	�'�٫tJ	�:�"|��a��O�a��'�N܊�����(�Si��t�X(
�'��]��K�I�$a@���Tq	�'�z��6�*k�4���J�}�u���� `��e�/��9BEщ/ȶE�W"O�hZ"�Yl�@��ݺJ��A��"Oz�YR��>�a�wl��d<^���"O.��G�YRTXs�lF�P�8�ڷ"O�芲�����C+��r�0��"Oҥڅ�U!�\m` *�7U��%��"O�d[-�E�`hW��
2|!(�"O�m��C�U䧓DH�e�ҮQ�<�S�
�c�����BB]x��¡N�U�<�ѡ֢s�����#�SK���h�k�<	A��*퐕{"��0V"��@g�<���e���jw�����S�j�<Y��#��)v�Y,BT��W�Ad�<��둥I���ꗋI���N]�<Q���g�`�`S�����*6�W�<�g�W-g���s�<u���Rb�PX�<Y��Ϭ((4A`e�b���u�SP�<qWCW1L�"�;�❉������T�<)�
�ByE!d�dzE��O�<q����D�v@�7�.LV�C���M�<� �21N��7��nWV�6$W_�<4L�$	TJ�ʄ�2K�+A`D�<����P��K�� ~��K�*W@�<�!��=N���!n����B��c�<�E�wr��tܭb@<�O�^�<��Ѷh`��S�E��z���CX�<���O�p]B���'��&�T�I�<� �6 �6�B�����3���O�<a")�2P�D,ᥣ��d���21��d�<1�Iv>�Y�#&ˀvp\ڶ��w�<	P�б�,p�޺[\
�� v�<�d�i�@��f��p�T��j�<)�Ub�.pB��¸,�9�1ŝO�<�To8?��/Ƚ ^�� ���A�<� F>z�1I͋�$��FFe�<�G Y�;MD��1�c
� �S,f�<I�hV�U��E&��nT $c�<�D�V�qV����1@��#��I^�<Yè�,	���}.~a��9�B�ɡ���
�-ˇc�V�!B�"5��B�I`�� ��皆&H@0�ALhP�B��`�	P��|�~�c���*O�!� �:F*0j�o�Ф,`�
_�D�!�d�{u6��f������U�w�!�&`T~a���� u�((񤬄(�!���#����lE��
� h!�dǅ�V�LF;8�l���zR!��S�&���P��s�����W�k�!��+M����O��KMn�e߾S�!��'}���j�NR7"��$�3h�!��
=Z芑��#>}I���t�!�
�o�X���E���B��r!���H���Q#
7���c%ܥvR!�D�O�R��$
�h�b�B��k?!�dw����bK�zo&<�G�0!�Ĉ�r�~���B?��颱���H!�dͶkm��q1�p��<R�4Z�!��I>k(H� ��M�4����a.��W�!��E��$������4��|KpC䉴��u���̍K��kq(�>q=�B�I�8�x xEW.1���M�fB�		�!@�W<-�H!+a�` B�/jB`��D�P�!�D%x𮃯�B�ɻr�(�E�%@�K��\�C�)� "e´��&+Д���E��w����"OLњ<C����5�܈V0v��"O�MAs��z(�����qw���E"O��zqCA�i�}"R�c
�r7"OT��eY�|���o,�P�"O�a�ׅ��t�H�"�*�+	�8��"OV�`�Of���镨�E��"Oys��� �#�$:G�H*#"O�D��UZjH]1�`�,4F^��0"OXi*��A
$oD �h�mC��E"OD�F�ܨ/R�dyҧ�9>�`�B"O��E��|��Q��fI��詓�"O�A
@����J����T"O�X�w)Υ͐y{ ��'g��[1�>Q�d�h�cÜ=�ֵ� ��G��)����t�2�L�]Vl��oQ�m�ȓ��	��i�:Ť�cc��M6�m�=�����Tj�p!��ͮ8�4t��$�%�y��\�zFn�Ʉɜ�_�0�Iڰ�ē�hO���U�fĊX��5ivH|�a��"OLxk�܊A+nБK'q�d�"O 	b3�Qp�D	�AGG=sX��(�"O�dYFLݳϬY#T�[E��"O�<s�K�
#�qZ�*2�{R"O޽ZF�چ4s 0��H&Cɂ�""O�����3*�ޙʑ���J��,˔"O� �Y�h��VMF�{��urs"O2%`��bB�@�N�W�(�a"O�(
͟%�Q���'zΊp��'�D�fO��X@�7|��ae�0*v!�ʠn_�	c��8@B�袾�B�ɋ7vp���Ã��H�6Ś��ZB�	w��Ii�_�h����Ӂz�hB�ɟ6AR��s��1*f���7����`B�	��$�H��]�}4�����a�JB�	-r���b�[�#$�8�P�FNB��J�n�eN�Bn(�3� ؟0`^C�ɝ$�M�ƅ�Q�6���b�N�D?�xq���D�Ib�ƒ7�rl1�K7D��k��ӽ|o@5*�W.w���E9ړ�0<q&j»1��p䇣,�h�Bc�J�<�n�[Y��� 
%S�|�l^I�<.L����Oωw��LkGm�kܓ�hO�OO-�Fd��ةP@��9W�,P�'M\yRT�^,*�����K�K����'���SQ��@� �m�,A�j���'޸8
�ǍC�v�P�Í�H���Jߴ�Px¯�.q�������
l�}`����y�N�#6�d�Ib���̀ЙAJ$�y��փc�jx�"�	7Ԓ�ՋW�y�͜�$����(/)�y�L�y���J�!a�q�ڸ+�+׹��>�M�$b���+�,:a�91R��#�$D�L�S�EN��M�0�3N��E��
&�Dh���:�L�B�L��d��9R��Zu :�O����'1��ٲK%h�!i�!<`4�i�'�*��Tn�@h@��XQ� }��'̒�!&�g�tI걃2Fr��'rb����H��D���?��}�H>9����� `�%�U��*w��
� A�W!�䉤L|Q��6���%��&�!�D��V^���f o��k�d�4L�!��"0ل��g��fh� �W�i!�d�8O��8S����1E"C�G�Y�!�� \����T$7���b�5t�H\I�"O����d�d��a�G &X"O�j&�#tz�"�F͆;|���"O$]So^�,K�H��	%��8W�'�ў"~����*,2��aQ-�09,�ǈP�yR!�X���D�
�+�R�ڶ�L������>��B�'=����nߒjN�Z���s�<Ar���TW��Ƣ�F�n�Ra��m�<1�]�*4�L��I��I����q�<��ڤS4�	�)�=[����HG�<q�� F�����!�?11��a҆�g�<��@1m�-�%A׃wiµ!b��K�<A׏�;ٚ�k�m�<0�@��d	ON�<� nڒrGj�0�ݰ#�� ��2D��"�H��4��O�2FTnD��4D�p�u�	4o�A:���g4�H��3D���-G�5~P��IBR�,�$�&D�p���W�T�"X*%���P3N�R�A#D�p�Qm��i�1@ȵGb0�L%D�4cp̊�3y��c�E�e��% ��#D�h�pi=[s��[]�RE��1|XC�	/޸h�G���{���ܜu)����>c[6Y�E��ʍ:ܔ��T%|�<�g�
ts:R�!���왣���z�<A�o�>3���h���ViJ��\O�!�D�,p��5��E�8��gH$y�!�D��mX�,��(�[ъ�F���!��d���\�kX���r�L�;�!���,��Ѻ2L�u@�
�l�7@!�d�2NK��!�V%"j@�d�Ĳ<2!�$�Y��-�� ��yB<bg�S�9-a}�>���`�0��Ǹ����ŖJ�<��ݫIj����$�=4f��a6b�@�<�,������%�ĸ(��=c�%��<���]��Hd��
_4 #
��	�P�'�Q?���� :c����غZTY��-&D����d41��M�M�l���M%ꓺȟ(l��R=�faB���FP��"O��"%`��&����gCC�Vp�t1F��$�S�iΆh�|E#@JʈX0|�a4�<e�a{��>���X2%���ͽS��œb�C�r"=y�E�b�CT ��L<�Hk� Y������{�'�88�m�/rl�B&�̏c��J
�'U~ ��%ѦY�J}��`��S��!��OΣ=E��AU�'�<I�Y
�]a� V$:�������?�Tް)��$��D��FU�RZ��=� �E�a[U����%"^d�Dh�TX�t�?A�̜8V`���ꏪ;q��2`)@�A!�̿l�l�����Je*w�V��!�$��3��]�hxIڔ���k�@x�'���E>t�`��E-LN���Q��yr�T$���ҋ��E��"��y"O,4���	��T����,��Od��D��!�<��`ƀ�j<�ծ�v�xb�Il)p�Z�ˌl,�=k���B�	/$y-JrKȴ��!{!�0/��#<��0?ш�)%\g�(Z���2<6��cӅ�!�!���q�Nd@'��#�����A�ly�$2�g?��-�Рp�aʨ ��	bN{h<9"���C����uD]��05�!f���?���0?q��SC>���R�Z�i�^�<y��
��qcP- pʹr�Y�<���<�	>l=: &�@�<!�D�N��Pᓧ	2- j��M{�<� ƀ����p�ARNX�$1H�"O���!	F����@�
�(��U�w"O��E�7m`���t�%k�"OnMX��Ox��p�ŏ��5�R"O��SG	�Ab���-ءI��A��"O����:�x�s�ԗuI����"O�!��㕂~���(�c�@|M��"OlP�%�˦X�",h�&�h���"O�$�#%˯|�9B��!�*$h�"Ot���KA�I�,�ɐ��"C��"O�l��j)p�	��[�>�Ih�"O�@�	I�kf��b��P��`"O蜪�/" �eK�A��	��S�"OΙY� A�CF�ـA�1R�1:5"O��AS�^'$1�˒�ܬ"�x�d"OɁ��K��\:�eO�o'�И�"O�Z�3��ѣ�?{!*�X7"O<���?V�\$�B⁗(ģ�"Obukd��H��`����1`)����"O�����3�F��w�
%y��"O�交"8F�%�t����Pc"O���C��@��LL:ܝȰ"O�{Dm��֝@uaC#�%�w"Ox�	�dӾ^B�����0(���PG"O�q�tkɴe%�}�Q�]:)�y��"OZ4�.�4Qh&LГ̈́�N?d%�c"O:Da��<�<Z#��H�p92�"O+�H�m�����f
\��	(^U�<�A�̾/`�UC�K�1wS@,!N�<Y�N7p�P {Q�Q-W-b����Qp�<Y��(p^���� >�钠\w�<��aY0'��XӀ���� ��TK�<9/�7��ڣ�[$3��JD��Q�<q��kC� $#�'o~j@���N�<�pnL�vm���o#g�D�z3��Q�<�e�\�f<�C���~Y�m�M�<)@��C�HX�UHY�ղL(u�K�<�/
=@��Ё��'��#2.�F�<憉8P���@�Y�A��t�V,�A�<�'#� \D��HF� wИ:�A�<I�����叨[%�ͫ�-�g�<���|a��D(x��S��h�',H�ARa���tx��� tEBAh�'����P���+sέz�C�'6��z�'{�͈�͛�.� s�f��P;�'+BH!dڥ!Rt��LV�Tg�E��'ʼ��pI)�@�R1�Z"O����'gh�yJM�&�PɨUɂ:�ҹ��'B�j��Rd l��U���5$�J�'s�9��8!XV��P�Г%��� 	�'�~e[���QI �����r�G�<q�j��7�<�02��Uْ	�4�U�<)D%�䚲l˔k�<�LO�<!�HγE~�qAg���?|�ԭ�I�<�IT�t7�	��$�~PtݺR(ES�<Y�釄D�x�"R% v�^�zV�O�<	�ܲx�<�y�.�=I:8�Z��q�<A�O�l^^�S��F;c�R���U�<Q6�)B�5bĆ��
2��B_�<��B��*2�Y���0U�0�)3E�s�<I���)�d�b�D�':Ȭ��э�i�<��%ѩq;��y�쁹��1ه��a�<�&�ؠjj�	�!�E�5)q�ÅZ��e��k���FmL�z��9�[Ab�����s�<�f�s���jã�?i���R��]eN '�x��/���)� �9Hp-�_��A���?�0�p�O�Šr�]K(��hćZ�F�񰢭�(��=���OG~�|����]��/�]Z<����İ<��%�!��d�̈́�e��dH86��HҐ �(>��l�2��%F!�Y�,G
���l��^��,[7`�xF���R�:]����q
�����ٸ.D���Y���Ͽ;d�_	JX��C�$ w�s�YW�<�Ǖ$�X�$�_�w�H����E�fp"J� M��K���!tt����%�^��߹v�N�'d�u��ć, ����À�?9���ۓ\~@ٳ�G�_��X�f)Y�]tl��G�K�hm>%��L�p����g�+y|�4��&�+M̰1ǹ���s��u�E^�Xh Y��4���76x��=�������4��dB��v(`	I/o �����'L"XXe�P���qCnGg��y�HV0x�6�xhH&�8LOF�kq��Gւ%e�ϐpC�D���/\�1�X�S�(Q�D?T�#�╚Cߐ#a�u��T�T��A�Y�Wց�p��`R*x��ZM�<A�$j��l��>dR F���y�F��6�$m��� a�xtIa�'n��T�@-s����v?�����n����P�<�#�"Ӣ��$��v¥�����l�x(���	�H#��+z��x��K�qߎ���.3W����g�̤.���Q�-X�V=KO٨|�1O�Y���(?��)%��C�Ѝ{b(Ġ	�Z�7o�c�H�q����_�Z,��E-q�2��dӽ3i$`qE2^���B� C�fG �㦂T 4ۅkY*�0=k�<�����E��!�j���,E�u���{A�I�~[~�"�͇;�B�b�N�����we�+%�d�����켻t.ٰ1m�:5Ԍ|<Z<��W�<	�g\�Z�|Y�s/M	#bH@�
)fp�u��N:�ڀ�FE'I�f�2�眔^�jmأO�'eBXʔjW�a�IQp��f�Nu�D�����Cf��p���@�s�̱QU��PZlH)s�wy�bi�<2 .�8W�VQ���g���-�(�[� �t�payE�
����(OR`��kӢM��0�/��XP��[4�	�JQ�OP�4����ӵG=��#�W0�y!Q�í5��Q��)RUn��WCW�R�j� ��ئ�0�`��[z�|�B�̣xn"h�1���JK�P��Y�*\��g���b���ʇ}(�Q��!~a<T��h�OB�L�w���u�ш�{�8kR뙱U�`�8"�6D�$3�mI����VÈ� �f`y6k
0'Ԃ�(�J�k>�<{�ǔa���m	���6c�0�nxA�KK�#ݐ$H�NMp�ee�	�JL���-lO�5��y��Q�"]�E�ݣ5FP�C8�A�tj\*���� �>]c����N�Љ��[�G���E��8��'�RȠą�Q{�� T�S9�࣎rj��}ׂ��a�K�R��]A���,IF�MSbG'=xVaj��Y�vt �J�l�b	�S��%q�j��լG��=ɔ!^�i(>��J�%�P���H�L�͉����<A"��$�ԡ�j/0<�Q��"�|��aH��u��v9X�Pӫ��~1l��WC�!���
�&y����a"$I��mMF���`*'Z$e(�"�'}��L,A�	�.u���~��Hy�]��V�����M�1��9)�*5D��b�\�SԳ@/T	I+zx���Q����Q���	�B��Ģ�ez0��2I>�Gb�SǖYJ��3a��qx`O�\��ȉ�\�ds�Hqw�G6�0��g�^�{Y�1��kqC�H|�@�����<����vB��q�
+G�� r%Q��"oN�R�B�$eЩ, � l��TC��t���ai�v`��4A��Px�$��%o����C��\ @F(��!��E��`�V5�( �LV�9��$c�.w�넘F��c+���yrE5>`^�xĊJ xh-b�/`X:d��F�A�� 8�GV#e�`�i��d�1}2Ja��XB�D�;����W<`U�B�	2<ľ�U��WQ� `�.�'�4(J��:U8P�%́�x�9r����p<!�((���4��D0�k	@8�,*T�[�a�n@;�!-"Z$�V
W-*��
!oՖ�>�[�aݽ&�|��
�'�\�򶫞�70~Yk��{�䍛O����LK��l�c�OV(Y�l�{���.�O��hւkV��cTL��v;��r�'���ؕ�	�i?*`��`�hh&��ZV���&�C4-��U0���O�.�'c<Ið,¥ъ���Oӫ[(���'��yH��WԤ���ͽE`�0P$��:G4֠�����Y���3��F���d�$ FX�db[��y�� ���xr�n�6�c4-J�Y���)A�w�Ĥ�WkN+NY��	ͽ�f-K�,�����Sp��5��=sj͂�.1}���x�8��Տ��?\�M
Q@�z�B�>)�(W�' �sr�r+tyA�8D� !
��A�J�·�L"Z����ؠ�>�`T�*y��0�e@��IǞ�>�:H�ppt�P5U�p�CVd� 0�p���;�<"6��$��B�CѠQ*���q"�,g���2-Q�49zBɽ���p<	Q�)��,��NZ`t���憂N8����h��l1�����Z�0�s�Y�� �(���)($8�F�#�-�ēt���#A�W�r�qPm�+%�&��O��
��8QEZqZG��$w�10���V?����<w�Vt���?|�!�� Ȅ'�E�޽C"nE�g��*��Kw��d)ݺ%�VlX֮�,'�q��'����(��n*��� '�2iK
�'����N��XX�+�<XI ��«j�f��aD>t���d�p��(k��0�r௘n���s�����OLq!��ǿd��!���G��=s��39��S����!��#=:�P�'>�)7g^ p���T�=d��:�O����O��\�Y���숳0ʧ0lF��s�>4r˕d���ȓ)�Z'�N
Z�8� �^-FL�T���Щs)���a�U��*T	F��BX�#M�y�d`]�WN��#�,\�m��I�y��W��T���ST�O�?��D_�>�|Au���B����I��p=9�L�6k�X�b���I?.Mh2�Ud�'ɼu���6-�`m� XJY
��6)�������,�j�D"^%�ȓG��dg�K�U�lЀu��H�&�"X^���#�/dp|*�a� IQ����S/0�@�x��:q�T䪴�(p�C�	<#���A%:N�9Gʃ"]�<��"̼)*H��@w�&�5*�dG)�	�'�5(�*M>w&-�A
�n���B�X������ŬS��`�L�;ne�w�H�2@�RU�I�+�r傓a�f��HR@$I�g��2 *)Z��=9��8�@��1f�������F#�]JP$�z��l��E�M��\�a 8j͒C�1v��ceR�6Hld�&零i%\���*�L���J�OԦicq�9�轀����*��D1cOZ�}��p�Ι�r5!�2;ڤM:����m��C�[�5�ӭ� �<xq�Ο�L2~��%�~�}"�_�+:����ՍmGr��!��p?���B�{︄�$�	E*�ɳ�j��ZyZ����Oy��i���i�����ɆHH1��G;q�,L���-�>���2+�h�['�i����'~>���X�V]r����A���!7�*D��P����J�ғ�X�-��|0�n�>Ag�W��q��&�0w)P�����;�%�5%ܯx�BIp�ڐ!�DiM4q�cmV�)��d[���)�M��OT=��ΕqU���qO�9o��(�*�@EI�w�D��O�K0z.ʵSE���pĤ�<+u���"\�T�,��D��6}��+�J��R�({S�x⡞�
�Lp"I>1������&�ܘa@PÍJ�<	���*dp��m�Z8ȼ��F�<���e� %yB��6j9�(�`$T�|@2� ;> ,2�e�R|$��#?D�d��kl�b(��藾^�!*�:D�pIt'��4HPC�.��.��� q
7D��BSa�X��{Qo�A�d�qӎ4D��x��Q-�v�胆�!3jPq7�4D�T#W�W��V�>f�Lب�<D�$��&�|������E���9W�4D��a�F�Ж����^r~ܠ��5D�LSv͍�p���ٔn�(G��MK�3D��x�G�1�B�Ғ�Hi��0t�3D���W��L�&\8S���~9��'�8~�x1�?�|���W�䨃!j�xh��Mc�<����+&�Z��݁7�*����Z�qO�hk�,�3}R,@�4�����(sR���I���x�fB�c�҅�roY� ǎ�kF��F3(�c�Νh؟4���M�>,Hi���Ty���Bg <O@u�@���ē!@�QS�"#�V4Ca���s����\\�];!d��K��H�GG=G,r$�D��'��D/qOq�.`����4�u� O?"�
L�F"O���'ۑ3���c���M��`;��(<r�Oz���>�3}"�2#����MɧjF&l�.���y����FǤ��@<
8�s.Hn�Q�8c���d��&q�
Ίn���
b��$1�azB�Ͷ^LJ)a��X?��C*i���e�*$-���Tp�<����B�����/4pP���v�. \(R%4+�~� ���,4���.No��S��Tq�<ɡ!ρ)�񂃜<�&���U4� p�� }rI)�����@�6d:dɆ@��������vK�C�I�f4���͛�m����2O�o$��P����?ۢ5�&Χ� F�#�
U(>�y�Q�̡M���u�'�2���P�@_��H(�c�K�k8$���
�v�ІȓyH\�s�D���aӇ�ŦCψ��<��g'@ʆ�� �'*�P���癬g*(�"P(�%_�^Y�ȓB�6 ��L�e�reHvꏉaE�2T�a��'G�F�,O4	��]�qa��pm9�Mx0"OvMIw �H��@�bKϸ`��|c�"O�D���+5aу��v�^�H�"Oy�4oD.<�����k�3U�9;"O��B.]�,F�$�DϸIs�"O��6�[Kn�	&�e�b���"OFif�&����#^�L��;�"O��� o:)y&�S�̐!�����"O0PcJΪe�Ր�	?f%�푕"O��pD�	*6@1�-+T���"O�� !�%��`�VoA
���#"O~�H@/؟w�k�OIC��Ě6"O���#O�2A_���.�����@�"O���'��B�R����B��4��"O�����	{� baF�3O�u�"O��A�Q.J%���/��Jt"OdX�ٞ� �5jӻZ8� �4"Ox��rJ���p�Z�Jָb��s"O��Ë+jzɨ�� S��`�b"O��i�ZoS��3P��H�5�g"O�ճ���dH2��A�NW�(tb�"O��+p#ֈP�$bԱL����"O"�1�k�(���/�#F�p`��"O�ģ��U�hb~�!�oM0���Z"O�)jdM_9$t<��ԤE�<�F���"O~�SF�i?8Ĳ �ɧK���aC"O�`E�̵eT,�����v�b5"O��ץ�?i�r\����t�h�H�"O�x�֎�/z��ڱ�ٝR�^0B"OJt� 杮Pr�@0ԇ��3�|��A"O��#�ˀ�="�A�'�D��1�"O�;rE�������(K�J�c�"O$=����PFO��� ��"O��A��I=X� ibI�'_a\��"O>q�TE�f��m�p	W%-�� [a"O��d,�)� �(�IĲe!P"O�Yht��'��������*\*E"O��!�]q��&-��p�����"O���2�u@�A�A�DOzX�"O�xIU�+&$��Ri�5u9,�Ye"O�P�,�<M�˷�	��U�"OA2D%G�5{��#�FI2y��q�A"O�I�Eg��}2����[)e���x�"OD@�E"V�K7�m�Ӣ��_�0���"O��W���֕�g����P�%"O��T��'re�b�D��X��"O�D�a��Y�
�8���x��ȳ�"O�<XQ
��02�2�(١x�$C�"OD3�R�N���y�H���0�!"O��Rr�@
��@Z1J)V��Q"O8H@�MI�ބ��f�pA�Ae"O�0�OC�,��4��>i@���"Obh�𤐊0�bɊ��3XQ�	k�"O4pj��2,,`���JPNళ�"O�Zw�U,I��E"�
���R�"O��bA�iKԜ-I`Ȭ�o�y�Kɮ88
���Ρ|c 9x�,��yR��+e5� �@�j�U	4NY�yrcĩ �b���ě�;Lh�vH��y
� q��-�.r�A���="�0P"O��0	�RJF�[p�V8_/�40��ܯH����S�9����Ox@,%���2h� C�	4U��'�ʧ"�R��Ռ�$s�P3^��H?�LE��O���e�:�1r���"?v1`�O�X��*e�|�g�Z-�\��%�R%9+��2Fʦx��|�
�8\�@�p��&sE�穞.��<�&a�:N�4�SS�\V�D_�� ӥg�,�ج⁍ 	XD!�d�- ���L�7g�($0��M%$(�o͈Ip�FNA@p��a� ;�A���ɜ�AS؈Rw�ǽ��Ъ�c�?W!�$U�w��P�.�O����L�#DI!�)��'��un�0/��i��	؇��ޑZ6)�ʖ�u	���!��DС��.bv���:E�0p��1X��8vF��xTZ��6s��` ���beџԹ��R�$���pD�Кo����5O�Ԋ��ЏEd�I�b��Wr`��D��)a�U(s�E�`|a�e�5\�p�26�1�O��1�F�� ��%Y�߃��AsE�>Y���>:5�6�U?O�L�d� lL�c �~���ٮ"�,Qd�F�pdL�iwl�d�<y��Hv	��H�]��P�*�%pO���DVZ��=����2e�}�v�F�S�6�I�L�XA�P,]C��`���8B��B�ɦJ�J�2�L�OT�B�dC7gs�E㕆��T��,r1��2E,@懝�ZnD�j5�,�?Ѷ�*���#G�~�G �����H����ݺb�b3#�7*��ի�I!��b��!�vi�"��?� ��T"YX�<�u��K������]1?���� }r�:awhٳ�^ ��I�I��QʔcfW�>3������W��'��5@Vb��s��C�I	$B��Paޞ#��@C�7I�9����A�![�0��A�j�%�Oj �۶)����-,�n��`��	b�I"cq��D"X�BTc�+��V�d�H�^tq+�n�5s��1��LI�8C1�V44�Pxw�QM�'Kj�:pOQ.&��sBܛ	4J`
�D��h2OD�wb<�@Q����b��� X�Q���,����-���BY)�@4v\���W#6�l�ÃGމ!:�@���*��@8h!�#_��2t&Y�uw��C�����	�%�?��CN1Z(�E�l��X\����m>D�,���".�4���ѼC�l�	��|hrB��+�[���Fs��@��E�d���6��DϻڨY� ���ԸI4�5}X�<��+@�-��m�)S/�H���5�
8ʄ� )�:�:łI�+�H|+��� K��5��P(��x4��0Є�`5��Q\��g 7<O��@e��RZ����E���9Gh�W�+�N��`ے��u�t	U �?A�I�	������J�1����'�,1W�c���
-3S�y�KɈo�xrc�<z���*�&	��D�ǡ��:a�m�'�>-� 	&'*D���.�Ja��V���L�p-
/@�5� T�=�~Y�Q.�
۰�*��ؒN�O�M�;j"\�����u"耮b�<x��"OLp8քI2��P��HA�|�aq�#�eF�x��K�_�0�7.ٔ5�O�%$�T�v�S9b��8⁤�:P��C�>�O�Y�
ScU�0b�ǌ�3�-%�V?��x�EΠAq� c�S�f�#	�!u��pǟ*}7�u��3L����:�X���,\�En��%} ��C�ٜU�l������}��T8d��>G�C�ɤm�t,�¬��1����V�� .�L�'av��S�W�FS���Y T����7�%3�L�3�[*,a�ϝ�12C�I<W��iqg��%�x�#K�:o6�ȸ���z������<�����#*�S��'yDA�Ν�},��r�cI;-��B�	�>�x��#ՆT��-#%M�9�m�cJ<LQ0��7]Ș�����p<Y���64,P�+&^q�=��dK8��`�O}H�eJ�Z#L�����-x�pq`�cɖ1`��S�ʝ�`͒�',-K"N�>ݘ@�a ����L�8��#@6,p�c�C&bF�큤gɸOD"v�P�unH�3� 2 �.�	�'h�B���(��e���;L�
�qۣ��B�>��Ď=��O��'���7$�*`��ՂQ+=�*��'����s<��r�cN`+�mJ��ƻ>��𛱋@� 3��h��Wl��d��'w���%UC�NhP@'C?H��x�We9cq���>�s���{�����?W��IH���F��̉��<�h�%�p{�����9�ѹ�B3}��	t0����D�j���0�N��~�>]Æ�9%0�2�K��-��5yC�/D����hޜ}���Z&�ƖN�܀;G��	Y�����`jdx�$N�9p�z�>qO��8�N�~o�yc'0j!�5��`'ӌx?.t)a� �] T�����e�<��G�	Ժ!Ayl �Q�S�? $Y*�4s/h|�Sf%6p��`q�'�ĥ�a!O���f�D;M�Ƶ@�H��%K0i���2�V�u�!�W?>�}��V,�-��eY3��-\2���
1=i���pǆ�L~�����Z=8��S����^��#%V~�<�R��ڸT��U�U���8��C#*ʖ����-nZ-Y*I�. �}&�P��T�U.ܢ%h�z�T8��H/�X�G�#�@8bN �@Sǩ/@yr�E�A�08!�5w��z���
x��8���(�$!c�a!��O.�g#��W��T�؅8��9�֫B?�Ҵ�&W�C�:ŀpG��aќC�	i!���d˫='�P��T��%XV�1��0b���K6` ��TlJ��)�q	4��b�U*e+T�\=!�d�>X��Aa���'_L��h�@���/ݖrk`i�%A ]��8�ה~���� g��i.�720	�FW�M�~BI���c�� _ƴA��<T�@�ڤL�S�����"��sM4\O����
ߡ9��(C�ѥh�n�Ӓ�	*(��9³�
4�a�J�)�̸���I~��ԑ���us~1�����!�L!F<&0��Ʈx�L ArC^Q'��є+3d�����D�B��Q�UE�$�û�6�S:���rC[��y�MI����r,� �h�p!ϠeҊ�" ���D�^%!p M��0"N?�Z�{��;6�ɀ&��~��Y1�k΋�p?��"V�2�� z��8%F�hq�Oa|�"'��!0�6��
��)�4�'�&<����4&L�|���S*������$I��a2��h�*�Z�	��O� 8���9#vH��ҌU������9�yc�!+ .���aF_���ѡ�R��~R֎:t�rVlO�Y�p��1'j�|zI�=;�V���/. �U  ��\�<!!%��o�Ȑ.�!H���jåU��a��� ���Di��.p���c�P{�(f
<,��N��l���.�O�6f�)C�	as�[�Z$�'[vW@C�FP�3͚��%o3cy���$�
Z�U�QN�����sNyVQ����H�4��-`�޸?��]�G5��5��.�u� cakؼ+�܁�"OT���%T�\��k��J`|�ST��`�_�^t*I�`cۜ#(r�F�d�����҄�R�M��\� @J��yd��W�T̻�B�)Sh�������D�A�'���#e�
&�ϸ'D�Jd�ڬ9��	oB|�<���O:�Ո$>��Is�b�+p�❣�/ 0P��t؟��p햂A�p̹��кx��p ��?O-����B��'�9���CL��c��j���'��:S���i�ȩ���}�m��'��ZČ1m��[���^LV�0�'��1� i��PtLM�T���	
�'�P��k�<&EY��.�M��$y�'��ɓ��ӟ[A.H��A�}W�L��'��hق���as���%G�iH���'���K��U�q��1¤� 0l&��'�|���C�� h�u�5�F01��!�'!�@bm�t�̭3ƭ�:�L	��'��a�#��	j?��&��In���'��kM�?Z�5�� nA�@q�'ּQ2�����E��8�H�'��l��C)��%��iN�}4H8�'Lu{��DD��GCh(�%�'rF,� �4Ύ��߾b8Xr�'���ƎC�u}K���>g�� ��'k�@��BH�T���PH)�
�'p��)Q�ys|�*@�^>A?�p�
�'��0RlI
rx2��.�C���)
�'l8�� j���].:t\qP
�'��@H�g.�\˅����P	�';����j�&	���@�ֆ�J����/�qOP�F��O�M@0I�8�T�鑊>x��q�"O�ܩ3�_�%CsQ�K�rn��)J84�ybB�qX�pʐB�?{�I8EKm��4���4LO ����	�Cc�Z�'�:D ��K�	�hdq#�޺.�6$�'�F,�ƆP�#cJ�$* az�yR��!%]"��b�π ��c�R8=*�pq��<W>d�`"O����K;*���a0�F/9f��f�,)����J��H��-�g~bR6k�ˤ� �R���V㛣�yb�U\�ـK[.eHv!�e���6BR�pY�_�����6ʔB�Fշw�l�Ԏ!b����l��Q:w@E��~�m��*�f��Sh��Qݪxӧa[�yR�^'˸���Ö�MgV`�G�٘'e\X���ZB�}E����c��T�fD�NPZ��eˮ�yR�?�8�jԚ;����l@2�d��S�#�$�2�(��	�l-*�Z ��?�Q3Te��tQ&B䉑Fq�eȳ�D�Q��%X$�ڂ�|C��2=�z9�d	�0��Q��9wpB��2#n0�$Lh���d�:��C�I%IʐY$�V4St쁔�P�)�zC�	>�����M�)W�r���-JC�ɭ_Du�_! �ꐚ�R-�C�	�ze6���E�h	�᤬��K�B�,O����o�>��m���B0��C�	4�`i8Ul*������J��C�I�UI}�7#�6�YZ�q'�D9D��Q��)��h�է���*�M+D�XKAh �D��<Y��-\�!j�,D��0���;��eO�*l�UK�&?D��T+��ҁ��� p�`q�-8D��ȷV=0��9q�m\�@�ge7D���T�&e2�!�e,�� thPV/0D��	"���>��%�TGB+� �Фc1D�dH&�9G�d�����nh09���*D�$9Ah�>?����(�:p����"�'D��ȤA��q�V��0�&xκ��o!D��qPFF"v���󭑨=�h�
:D� �&J�D���R	��2F���Q@;D�8�����0s�͞Q��05�8D�ha��@*a�����K
)W��4Se�"D�����P�!c�-����c�(V�/D�8���S�H�ɓ��(&�4|jQ!D��1��0�"��*)+�y&�>D���C۶m�>% ��MqѬ��է?D����)��jPACO�#f�Ԩo=D�X�l����m��Oz9��@bD$D�\C���
�n��֤�u9� �c6D�4a��{���[@���jԜ�C�&&D����BK�|�YjQ"4Ef&D�d�0o�+5/���Qk�U�T�y"�%D���%҃r�2�Z�
M;� \�5D��yҩHf{F�z!
ȇ��uFh7D��x1�7\�<}�C��]���õ�!D�P�W��!�@�pB#I[�|�(>D��i�h� �5A%=,����2D��R$K�Ǫ��0*�s�J���3�^�z5:��6X���.��>�DΓ_e,3@	�%^�3gF�+��U�����#<E��L8g|I��-Au&�Ժ7
h�c���������dL�W�$S�Q�oշgd`Г|O�7gf $>=��?�d��m��H!��jVbE�=��'.�f(��}+�O�����O�D�(�E�*qĭ���	'E^2qAW_�t$����Ʃ���$�)q�P��񬕛%,Z���ԝқ6.U
t0��������V��&NA��p�Wo�]8�����y��;�i�m�S�'./�9:����� Y�H��l�GF���!�)�'L��*���>G���(�ś�9�(D�t�)��'�*@��S�@{1Y1��\�wŅs%�����d��̑�/��"|���ǲ�\}�(�b,0�x7	Ʀ��'��I(�"�	�~��n�?9���S�d� @@���W�"<cR�|���P&I�E�*��>�ϓ}�De�f��#�����6/���j6l׌9�X�}m���|B��O�����D�:�T�Qj^�*e��L<�~�Z�<)F	�t���F�g�? �a���Z�H�`�p��L9�<HZ�_6z���i>�}8�V�ʧa�|���N���>I�&�ۅ�d��`O.w]�@
D\�o�zp��J>�Vܧ)��P
E
�$8�k��_$2��	韠��a	�ا(��T3!Ŕ��=c�hKn��ݙ��'SRH1�I�s�SnZs�'>x��q�'	B�i�$>#8��g�_�da�D����R��1G��j�F;�y��>��b͸v�a�Tŋ93�v�
6͟�5�4Yy��Ͳ?T�vV�|R�m����O��I���ty��aS�H�BD�� ���P��,���_�5�ƙ)Td�B��J-�s�����E�'�Dd�n�Qs- ��IX {�HI��O T(q�Sɺ��'%��!�OS� ,��1�<M�h[B�1�6����8s(P�D��2Z�^�+��:�C䉵Z���8B�xof��"��d�^C�	� �FP�OW���	�<~�BC�ɜ,H��»������!i��C�	�in�dx�g����%;�.��4C�I�q�F�ku��B���@f��)*C�*Q�.yB%�C7<���)c��B��>���@�:<��!Ƅq�B�	3/Ύ�c��ȑC��Q�q�ǌ\|�B��2I��o�}c�U�C�Q&�B䉐A ������wE���GDN�
�"O��s��Hi��z$�Z�ZZhӣ"O��@f�"�B!�K�j ���"OL��m��{v9h �ԑ8���"O�3!�H�@0�&�P�=}.��a"O����ҹ7<�� v�ه`�)G"O�9�F�*yRm@7r�� �"O0��U��z���w,_�:��4�e"O� `ro�_��D:c�M�K���A�"O�ձ��Ң�֬�O�1G����"O���*�
#(�R� �[�T��"O�p:U���B��7J�ӔѨ�"OT�G/HЀD�-2��R#"O��9f� i��Q��=k���T"O�y�W��$p1�1o� x
�!�"O��� ��X��}�v$	T(��"O i��!U�9���A�i	o4JX��"OX�q@��"l������0�� 5"O� ����z��Q"�R0�Q�"O���tJ�'a#zH� [�SꞙI!"OHMy2��4& ݻ��	1y�H�q"O�Pq!#Yh�1ዓ�7����"O�)!��3��YC��"����"OZ�92���f8�I[�kS!��Mx�"O��w%ɩK���0�T�6���S"O,(��?Y(��Qׄ�V���"O�Q�Q��<m����Y2unF(S�"Oc7@��4�B�r��N�ȪH�T"ONL�G*�cBd=Q�bş.g�isB"OD:�j��S��݋0�
'q+iUm�<	F'�O|`B���~sbd���l�<q�I��*#r������?-fL�b�h�<�R�V�v������a�D�"�c�<�tO1u:�]��D� =����(�H�<�w��%t8R�+3hO�s<Z��D�	A�<��L2#�=AeB[�Z���%.Z�<��c�5u��5�WL�\��B�<��Z�"��ձ�(J�Fަa��e�<y�,ɭ0[.\�Vk��>������c�<!��@U���i�B�-@l�[�<I6$��LlH9���f&aV�K}�<��D�{�]��!��X�d�
Vx�<I�ܐ1��%+�&4}n�I@���l�<�� �;aJ��$��09B��5!Ij�<� �e!F�iT*y��E
`��� "OFu��.M�D[D��B2'�<A��"O4 qF��:`�^(�sl_��X"O�=Y�)C�]�>�r��ſM�6� �"O���V+%x@��#��m��"O��Ku�C�g~& ��M����<�y�c	�n��}sw��2lh�h��fF��y\` ԘC�f��R*m�2B�?�y��T�m��$��`
�XW� ���
��yR��#�N���R�C�(��y�.�����IR0 Ӈ�!�y�A��x<b�Ⱦu�,U���F,�yaF'e���hc`�ne�R�	ĭ�yR�s*�  �h��(S�k;�y��{�d�yv"ηr�\���HM�y�%,`#��&p[0,�	J��yr�ĺp�тDG@�n�R��a��	�yc΢e����lSd_�hH򠈋�y��;֐M��H��O:0Ai� /�y�B�c'��"�Ó<A6�0�1+أ�yㅕ2H(# Q+'���ԝ�y�4\A>P��C�2�\��Ǫ���y�*K+�`��~�����y�"ԮP.橻���x����gF��ybm�%H�s�oL"u�.��#L��yR�/����F[�����ӎ�&�y�LV;-��%ْ�60Ʊ��)�y�IL�r��ISh!u8��.X�y��ȮbCY��풓D�du��"�yR��4n�
�(�!BӘ�ف�/�y��	9�̘����	��i6�V��yZ�����J�V���륧�+1�6B�I[
�a����>x���뒶^�B�I(�`���� h�0����vB䉊-^�@�aއ>[j$ �	xG$B�əN�l�y�!DK|`���
-�B�	1hQ�T�U@�7(<�c*Z�t�NB�	,+�@$JG�ϗ/�P�@�⊶i�LB�I�g1�a�W����A�<��C"O��!�	I�RA�|�5�$���"O�x[FF�,���]�v�Yj"O ��������JsE�+��r�"O�xhdl�.D��P��� 7�x]	�"Oƌ��a�� 
�]���F�4�e��"O<Sà �p��X:P#G�X��x�"O�I�Ď�d�2��H���-�c"O(3��U"n�h��G�8)��1p"O"�y��N �$q��jŸ 8&$(f"O+�$]��� "ǧw��u��'@y�<��f�x�<�
O�X<��A��J�<�3����'��M�f%�hI�<!*U�53$���GN^|�e�a�<��h{��1
�I�\
B��U�Z�<�BX�PN)�D�K�6����\�<�ao޴��a���4x3
x��I�V�<1��ĝWH�Љ�#�q��BW�<a� L�)0���
�#��p���w�<欍86F6� EB����X�i)���ȓi�4m��%2Ќ ����<ѐ��ȓB��I��T
0C�PD��<gAС��AN
��j\/ �y���2�d,��Y�б�̒ %�`�T�/ ��-�ȓ �|@"�D�mʪ�B�k-���t�0�ᙾ1 L0�ۧ.Eℇ�S�? ��Y3��z��X�
��T���"OԄ"��� S�5�5OH5���@�"O����H6�J3b�6��"O��`
9*ˆ��!C	5���"O A���,6{�|���+��}p"O0�C��7�<�1��H�2��"O�A��/gؘ��>�P�c"O2Š6���/>y��N�v�|`E"O$�R���k�a��n	���Y""O�e�$�7nja �A�,��"Olul�0ݤ<�1��)����M!D� [��Zp�z�������I3D���1/� <<@@)��A(j�偄	?D��h�㏥A��i��	_�(b�D���1D��H�$q��Cc�HR��p+�j2D�`�qHF�_( ��
#|�h��g0D�$!"%�, :� ��F��%�3D�<���B5T������n1�0D������)��#�لTW�t��"D��a��őꬒ!���\NĨ�c!D� �$�%nn�H�eA�4V��P� ;D�����s@��N���e
�gϦ�y�f@�Y�r��si�=r�����<�y"`�Y�`���d`ųsʞ��yb�E�d���A�)Ʈ'�����)�y�oɐ	�4�b#�\)N,� !�y�/I,i�����!�A4�+�$��yOĮB�橛��D12H&��%���y��$\���`J�%&����׫Ҿ�y�"�3M}�X�2$���%Β5�y��Q�u���a�ǟ1d���d�*�yr�� ֊<;C D>�5�ӆ���y�����+R�W B:Ιʒ�W'�y�S�&�����(h�PAgM���y�B�
ll�P���	V
Ux���y2EC�:��ux ���DP��e�y�iD5&"f:v�ۇA�� F��y"
؝)�T�!S7H�{��6�yr��E��0C�"M�2哧�о�y��ޭ!�t|�'�Y�.�B|r6�P<�y��
���kBiVwΖa��j��2bh�1Aiȥ�@[�zj(��m��}���
�4���C�� YU�d�ȓ$���� *ӚC\��"���&Q��ȓZQR<y��� <qtKO�r�=��X	f�Q4�Ŕ&�n��*W��(M�ȓ:�Z�Q�yF�qr�۔#�<��1uLIH�ń	#�2T!6�7P�	�ȓ=I��ѥQ�b�����@Pd��b��D��N�:R-�a�ĺ"7����N�iSi��K!�!�ҲiCht��7���� ��D�vj�2b�9��P|ظ�����!��aʯ����(��T��fU�

�(Z���/O�`�ȓo
�\��"����l�Ӡ�b]�5�ȓ�<ݫ#���r18��=d�8ń�ReT�M�C���۰�Z: 2>��=>��!�4p��a���7Gpv\�ȓk��;G��;8�R�˲[N �=����a�Y�c;کI�ج$�i�ȓ���6������`�,�H��vȲ�{�d or,X!�>Hu<�ȓv������� �,�3�9kV���3��Z4�=TX2e3��X3H�D��S�? V<`���No���d[,K���!�"O>��@�u`�L��É�~4��A�"O���@�Y8L��; C�@Qv!�@"O�"�lڼ2��ɡ�b�(tFԹ��"O�0($���^g����
?X,}0"O@��Q�
+��PtG�|i<D�"O.�8�`/i��95��
�D��t"O̭����c���àg[��p��"Or� ��!L�ܰ10��*^~��Q�"O~4��/H.�%�@���kx�Q�"O����h	5�X�Hz�`�1"Ou�S-M�ǆ@"�ߘ#�f-��"O�pi����7f�2�Ι{�"O�-�@�d����Ό-8(�"OP��!�d2R�Z� 1 �z$Aq"O��{B 
  �X   �  �  �!  ",  t6  qA  �L  �S  Z  b`  �f  �l  Bs  �y  �  !�  b�  ��  
�  �  ��   `� u�	����Zv)C�'ll\�0"Kz+�D��|���b�f ��yr�N��yB`�X+֜��$��y�"T"!��Fc"�(D��vk��I�iFQi�x�T&5D/뎇qC���bF<��	Nx��Qc�:�(����i� �sf�%��]�!Ў$"���>�୻��X;�'�?	Q F�h�*e����7=K��g���>���paX�	vB��V%���וr�7-� ��d�O��D�Od�Ğ�T�
�H$��)�V�[�cH�m.���O<�l�M3(O0�Đ�&�	�O��F.[�PD2ҧ�'�,�R��Xd���OunZdyb�H�=L��9�u��;���e�ty`4xf�A�Qݜ"�1'���IG�<!�OL�[��/�B�� i���[���P@�L.��%�F���$|� '���1{61!a�D.��%N��Ģ���WXՠ$�T<K���O���O���������O-��L�x�׈(yT��ՌM�h��f���o��MkuW�L��4c� ԋg�iG�Ɇ���t�q�@ã<�Z�R� xQ*F�=ғ
�μC���p�x�enF���t��X��BD_T8 VG�S0Pt�C�U�)�D� qf�b�&u�.e�x�n7�M[�'��T)Va��ЭҔtR�����G��e�%�,�M��.Jj4�̀�ٿH�6Uò�^��b� U��$����vӀhlڽ*OA���d�R�K�E�.7 ^A��$���B�Hf���M�i8�6mG!0 ���A�%ꔽ��
.	��9�J��)��H"><pQJIY'��m��"W0 B�o��M1�i��8x�����Y���I^¬j%)�
Hpœ̓#W ��J8W�P6m.��x(5d��P�]�U��"�	0^L�9Q*� ?�x�"B�@����{���?q��?	e�iT��f�X�0��ۤ�� b�O�*�����<����?���k���5M��% ��c�)[c
ז�&��ʂ
yc��(8I0�
>����"/��"�� ���(3����tirz�A����*j��5	��_s��qhT�7ʓD~�'u�˓}���ʖ��C�(��\L4J\�I��Ik�I���Idy��'�N�(iP�r��= & �63��;e�'�bA��0m�T�|���y�Oٰ���&��y�AHD�P}��
b��H'�Y�|�-��MS����O+�΅50�q�2�q��1r��n�"�'2�šc�K�H��5L�5 ���QQd��=ht@ɟ�����'Ҧ�c#�J�Wwf��R�(?�aA�2L�Wc݈)Ұ�r��G���t�����p�P��(:�I���L;[+��Pl�٦����If>E�U�\�*i����3m!F��l!�d�OJ���OL�$1§f �)0e�`NU q'�D{r�'f<6-�̓�Mk�O;��i��O�z8�0�gզ@�_<� ��AyH��	�����ߴ�?�,O����A�6~8i	�e��s4`�c�Id|>����ُ)ȴ 7 A�:n�ʧ���đ�>�4 � }r�c@�93t:��� �(����aɤTc�8J��C!$�lp���Q̧`�qq$���p��;%����N�B����B.Φ9+-O����'��t�?�O<С��X&m���aw���Q ��O��=E�d��iFZpJ���> ZL�u"�,|��'w&7�æ�$��S�?��'n����"����`��f��>1&���ۆ-1���?�����|��O���j�^r2���<F����A͞��$Q�$ڎ\�G�����z���]��L��gK�h�dr�l�MJ��tN��OP�=q�+��`,!'O��9�ՁS�[rP��	<�Ms�	u�vSB�H�IKv�*�r�)�z��O��=E�$[�u�d���!�D�b�qM��?Yѻi=��z�t�o�L��j�Q��7�OR牿/Ӑ�	��� I�-H��T�:��$�<)���?I�O?�|����[+֐��4Z6�0�k�E��4jN�q�
�*�5cR�@���%�(O��[M�8C&z����\,s>>��Q��)k}`٤H�H�Z�R�c:�8å�@~�<eȗ	-�� ~���mӾ�l�ΟP�1m���d�R�N,�l�{!c�IyR�iu"��3��Ouq�:���+l�|P�ր>��t�$ �$�Oʧ
6�6����%z�f�i������(267��OZ0l��[�zM��.
32e��' �Ԅg�|��@�u��:�!4-`�a������O �q���<�uslL�C��3b����O�2M��OEj��D�,̉.�n�Q�� ��(U'<T] !�_���Bo�Z�n9X��� ���� �N��$��>}(�$?L>��=m�ɶ�M����i��OY�l��dQ�X�J
:��'�2�|��'�b[�d[�m�2~fQ��NO1Jp�0����Or��	����M���d�l�M~� 7KL=b� 	��i���'��D�w��|�$�'��'Z�>�qė{�za�¨G{��
�+�	'���t�\�-�zXwa̸V����?]�J>�u�%UX��D�AWr�I�.Hq�<�{�X�[
��Vc�H��|�;}"L�-�<���R��$C�j҈eۛF��g}�N��?y�����?�� h"�2 G�C��yÃ(ˁ}R>0�L>��RL5R�M�,L����aɻWS���'��6��ߦ�'�����?��'�P�v�4$����Z+[�>q�a�M��6�O��D�O��Ş;%�����JY����Y�
7��3$"C��Ha��cˋ�B���<xG�k3o�]�'�P��\�t�v��W��#>\ɪ��Y��yrǨN z�@�˂�z���CE �|��m@�	2����|�,�X���&qp�/�p�
���?=�����4��'>�j&�)�b��ӑ��e�uD%|O<c�L��#�=C�ܩ��h��q���`#�6��P�����{y��a��7�="�f�E0>��C�����`!
ǟX�'sr�'}�	[�8J�`�!�����)QA��50� 9��!,����U�W=���94g�42������!-�����	[��XT���Q֦���M,VW�أ6��8A�p}��F́?�z�*c� ]J�&��2��On����ҥ�T�u��F���̂Dd�'��^�����>t�hp⨜�VSܽ	�F*��'�ў�S��A1�I�s5x ��퍩^/$@Ra.���M,O2 B�ʦ���ʟ,�Ǫ���'��fߣ^�"e��hު^.RT[�'BN�.r�>��I�_�ਗ਼ЅR�d��맗�Iա]�.9��P^����r+T����5!�]�۱e�uK��>�V��
�m�@���<��Di�e_I~�KJ��?����h�`�䂕O��t�`V������ҠK:(B�I[0��ŝ�@J�ģR	R�f"<)�O�aEz��W�u�~���hY�;e���!)�h'x7m�O(˓,i���'�?����?A*O]��C����BH
�z�btp�D�<	��)�8]�
ӓL02 {V�]���I��D	<�����8P��:��]gB� ���_�']#��'W���	q���j��y��D�iqL˓gch��	�?����p�YxB �l-Ȝ�@��,����?�.O.��/�SI~�Q�H��**X4x?64r�!������A�ش�?) �i��S�?]�O�>�jr%a����M��(��$�9Ep6��O��d�O&���It>yjDD��XsV��0G�Y3�'�7J�C��&1sR`�`F Jl�[�)[0�~�q"�{g&�1W ] A�n�)P�	���#>�Q��0�,kF)�Z%z�[#~p��I
�M���	s�'rT�d-��d��  �ɱ:��)���x�oA�hv�07f]���AV�گ��n���m��2��Y(OB�DU���QD�z*�A���Q���d�O�{��O��d�O��0�V+`\@A���g砤 �ԇq�P���\�X�Ku�O'��i4g@/uQ���b`:��y�$�}qh`N72�<Ip�g�}+ 	�F��!��
P���HO�ѣ�'B�7-��U����*�%�w~F�ժ�$'Ū��'<���'�r�~����;bX��N��:
�0�Ä���'ў�'�ƪ�koD!�ʎ{l��dU5t�6��O�<m�Ѯ�Qݴ�?�+O��I쟫�ipP�B!eA�x�6���dA��*��'3�*Y�x-�'2��IF%=:J��n�Z7�%y���!X�@ID��q��3�`˕�h�x�$K0.�,{"�Ƕm�tȲ��A���O48lڨ�H���SFU�m��6<��,[��O�x�O����On��=�'F@e9tC�:'ly)GhThV�Fb�s��mZT�'����f��֐{�b����4�?���?�"-Ī!)�=����?!��?y�w7r�+�#�	�,t{��
�o�H-jq!�!U@%)��\��`kh����O�F�ʅ�y?���1p�P�ʃ��&Yv����O��(�b̘�<1mz�fީX���( -Y���)��N�by� 5��l@�@���� �b�G.x�� � �n����OD����OX���<����?���	��]¥-%E1"�J�Z��o�<�R˂>,��h�*��AtL�J@�����I	�HO��l�󟠔'�}bO!h��j�k�� =[�<^������4�?�.O�˧��d�S�Ah�c��,Q���PlK�glD��g�E� �B���c"�b0ɕ���F��Dy⣅��0�'�:wFغ�-�k���A(��Ot�m�R��4
�`���C�\�Dyr�Y�iS7�X>>rbiX�M�L��}+�-w�f�$��O���,F���I�%S�ʨ<���$6�I�%u��+!J	�Z��$8ďԬ+:|�OZylZ-�M{-Oc��Ǧ��	ßY���+J!�gP���NIԟ��	I<���������
k�q���@�(p:!Cش�yg���fP�Q���H+lׄ\c7��0<��j�/s"��#V"H�2��Tk�/=~l�*#,�J��@L̟,0t �UÎ�<A%�H��شg���')n��l�-{ؠӑ떟6zVQ��W�X�	e�S�D���xQ܇`�Lə�n�ulbe.�Iz���Qɦ��\�ad��k
���o��MS-O���6t��������$��y�'&0��3X#��AY.n�~�3�'"b��%t^5�OF��"��CSfiZ6c��Udr=H0��|��1�'�0��
�]�,�"3nζ������0z�Oyjt�M�Cz��y�&�k2R<Z�O��#�'fl6m�v�O�i])�T�� �0Tp �됊xf�'Z��'h�Ӣ+0�0wc�����n�h`@'�ə�MC��i\1�6q'`��r5#D�H0/l�0FCs����<�I>�r��?�����d�4nTT�Ě$"�<]�NL�7.ʓ�?�T䓣�0=i�b��L��}�P�� lz�}�¨ҳoA���V<;���C'gY ���|�4!�|~���*�j��ʹ6jwi��֢�<��P����SI�L>�1CBkBXX����U���A#j]5�hO���)�2A�̲�A�q��� �\�'U剄�M[��i�ɧ�4�OY�I�0G��)BɒFn�i9���%I�l�Q�A�y���ڟ����)XwJb�'��)��=��k�b��sdd��2��y��AJ�Dڸ	�5=Q�1�K��+mvj��dM�-� *a�ٌ���Xf��j�F<B�`R�W���)0�_�u$iu�H�x��	�Մ5�$%����:�* x�̕����s��������������>�0��MH'��j#��kq�[�"n�,��Aغ2r�_�8&��`"�sY,�$�t�ݴ�?+O�}�C-�|���'��!!NK�gb&IZ�͌�	0�qQ'�'�⯌����'�I��]��z���*HV�P䓈x�N0��@�Z��<{�� HAj�$C��y�pЎ�d�W�\�z*�k4����7�8��U� T	�`G_2t�6���a[��	�B��:(�&�6%�O�Xn���=hH~� A�s]8'��mc�'a|��[�"�C��,,>d)��o���?q�'^eC���錐�eN� �����D�9Es��d�O����|�W��?�?�L�Q��l����ba�������?� �&Y &E�('��#�/�V�����O�XT�ɟ&u5n�2H�I4,!Νc2��4aQ�T:>�:F���X�[V�ٛ�n��$Ģ��Ɏ�Ӛ�W"��f�y)@��9~`��[����Qm�)�'g�aЫ�$u�ѓ�l�6����ȓX�
m�!I�.,���+��5�%�*����r�'[����]�L�1"��6q���"6�u�����O ��:/�.�W	�O��D�OX�dd�Zu �;n��h�2D\��P���EAh��,ǟ&�@��^�U�b>ո�&b���Q`@҅�$BZ�y�.��0��7�ҕ0T�P�ZpnM1�H)��q�鈲2zIy�'�5�g�f����B�X�6&���i�H˓9�Z0���?����yO�4�҈lS��@˂�w,�	��"O��Rp��<u�i���)���>Q4�i>���^y"�]�z_�d�!����^!���$>��9�/H�"B�'��'O ��̟����|:J��9�be�uK��k��ݫc�Ȯ�|�3퟽l�����Z)|d4CC��*�"�<a2��'"�x�ėb|�Ӣ
�\�P�I�j�A�Ԭ���f)��cD�<aF�;�F�p �ld��F�KQ�����Mˡ�J�'��w#e6��x�e\1<|ӓ��'��x�����(kBl�T&��?��4CL>y��i~�]��DB؟������e��0a@O
2
� �q�PƟ��	)~����۟�ͧ/����p̓w>�����A1v&�Q�v��Tj���ɜaB#<!4�Y %i��j�A^갚W-D�4i�O`�&���%Х4u�j���:!�R� ��!D�$jaf��:!: R�WB��6n=�	r���ݟ�z�� �̈9`-K� �f���'��X�K�ZoZ͟H�	I��H�44�*O�Q(�a!r.׍QA�i�U�T':%��'��ayV�'D1O�3}R���fъ0c#�^`�A�_����5pN�"|�$
�(ܚ5����|>����L~��1�?��|���D�$,@�qdJ� j����+!��0Z�ɔ
�>F�!�'K=
��'Ϥ"=��FKݎ0�"y��І��Yn�6�2�D�2���I�O����O�ʓKK�-�Ra�+ ��z�M/i�bޗbʬ1�$3G���Q����O��'�J�%MW $�"w��W�E�3� �]&d���Bhp	�]��O�'5|��Ԏ�1`F���)7n%����D�
n���'����:,���ϛ�7x��r�	M�C�	04Ů@�a�l�J�Ip#�'���Jo�����'����6�)7��ʳ�C#?v�IdH?Y���S��'���'F��sݕ�	���ͧ���y���t��Z��L!p��8pf(Z3��ap$�	�3C�\+d��U�`y�1�$���!�ǈ!P�%�w/$A���:�c
�v��0)G�J��;WHC1!Td� �#ʓA�:(fn�8?Z~��0Lɇ:S�Ȳv�����i��]<>#��K�.��A�r���e�k��X9�7E��!	��ؔom(�&����4��g��mK��iX2�'��$$[�I%���S
������'R��G�<���'��ɓ����`i� ����W�X��	ax�㍜�O`0CD��7�>` ��v����'������D�'�B�(�+Űx	�-Pk�a|&�S�'&���ŗ�(	FLP7'5[zz	��y"�|Z��'NB���O.swI����'*���J>�eÚ+%����'�BZ>�����ҟ��敢&�|�2� ��f��0YG˟��I� c���IS�S�L�|:t�	U��+�E��J����0�6?���k���� r�;���V�^�s�ND��8m�O �$�"|�mQo�:u����GI
dh�<� &�L9�!��.��!u�(��a�'���HO`�����hP��2Q�¢��N�H7��O����O���+D�o����O����O:�]�<�r�:�l��B�	I�]Y�3�ɘ1%@��d��2���2�'P:�`�Єcb1O�=q#��� �T����&��6פl&�,x&)��ץl �����,O�`�����O~�ؤjF�M@!���,}�S׉��") A�V�#-剘�HO�i3�$��ƌ:2P�a�n�S-	ZT"��r���'���O.�$�O҈�;�?q�����Ǻ�zY�,��sg�� �E�ZT)�`/���RyA��:1�ب��I,_�� �#	4r�E� �E5D��%� ^L�ra���=�������g�'pE a�F#@���B啙0�@�%�5�?A`�'�@�B��FR�q1w*	��fݑ�'�±B#W�K�)KT��I�`��M>���i��'���Fg}�2�$�Op����%�P�h��� �I:o�O.��kol���O���0���������[-R�y�⍀EL%)9��F�00��L�o0,��q��.); ��E� v����ZE�|"Ï�+`ֆp ፕ wx�M �+�>�`{��I�U����DD�	�$�n0ȃ���.������L��0B�	�~E���X��Ux�J��D����K��I;J�̲�-�&u�;��!���t0�o�����IP��R/r�א{���r����=�PQzc��	T��'�u���'1O�3}↛:PKRhSA,(a���^�*�'�<13���?%T�`��{�tM����$Q @��.��I?��S�OĪ�)tH�]�`1`�'�6dȕ�	�'4��lu�|a$�#=3����O�OmD �r f�Ġ�R�w���3öi[r�'���~�2�!��'���'9�7�V�k�h��/�"h�V�NYu,X�	O$�>Y�ÈV#��U揀Q�1�f�m�B��~b�^�+B�9�D��v#�x��cHV �1r$�)���`˄5U��`��D���<X\��'��
2(����J�h��-U��J>q�h��8�|�<9tl�!fjθABi�P.,���u�<�f�D�~n��*Y$���Y$,��<����HO�	2�$�)0�91lڲieb�ڗ(:qhq�S��̦y�	���Iiy��T+�o��h��pz1֎����L��*V)E���Q�Z�� �*/��iqB��ر�@a�	TDZ#"U��X�U23 :�yR�����O�X�v�Y0�Eഅ�0��X/Yw�KxӾ}Dz2ቘ?�t�ˀ=������$&�B�	���W)���r<�Gb6x��O���'*�I9)%�M~�3*�/�W�g�@9��H�B.���<i���?���/�`���9ahb ��u�a��B�w�,T��?��I2��@џ,���A6 t�gm:I1֤0#�]#MF��[iߙdP����� �ƅG�]��?I2�i���0u��+�V�Jjl��HG
(�'� ��ɅFv5�Џ�)R׺��%c�6S���D��,�ĆU��\!��+B@�3d��O��|�y�Z��'��i�OZ1K��~��m�q��
a�:u����O�����(���Kޞ/���@��D��������T`�	'�	�2���jqiZn~B�	bI����%n�xă��#��\(�k�Q��TYp�|��Y'��@��`�O��m���H�\�S�8�0��r^3vWZ-�Mu|tB�I��|U��,K'��ڨ�iDD%ڧ9n,9��%F-KZ�tkǏY�D��O��L�����?	���?I,O�J%�ÇRl��X"�Ι2� �D��QC&��dr������3Z��b>1'�|R B���(����R>�Bݸ�Q%&�B� ���%v��c>y%��e�D2�P�x��?��ȧ-Nʦ��.O�� �'��Ē?�ON�9f_���aaU�ﾉ��K!D��a��'����b�:��Z�G�<T�)�-O~�1t�E)^h��h�?vxQ���B�<=F�oZ�h�	�����O�T���I�T<��q"	�;K�q����F�N�K4EE��񑐃a�Ģ?3	�
h��c��ݺW�L��-EBb@�EmE!R9�6oȌ+$J�2���׵�L@u:QR��Ͽ|��h��'�F7��n�'��̠Qn�^N�)S�
,#p@݊��)D���)4}~&�� W�W\Ш��&�Ĉ\}V����A��'o{���3#2|��� `�>LW��	zy��'���'�~|�+�0qPĘ��	܈4nn=���M MZ�!�6�F%Z'�DHe�� �?�E�ֺ.�(!��ݤR���ISo��(�B�=�4���M9ue(؃��D�9l�B~���'N�+Ԁ�=8��G&����QN>��Pv���B#1���Q�yE�̆�	��?�R%G�2R&e���3g�t"���P�'FZ�`!��>�OY�S� ڢ�(o|�:�"M�X�"B��� �I$1A ��6*;���n��[FEZ��� S�6�p+���)Ҵ$K�lP+��ā9*v�Hg�ըt��#F)��R�N�?5��J/"8�)$#��alj4ɄI0?bHF۟���4��>9�g�? ���g�?L�> aсΌp����"O�Pj���YQ-��b�!T�������h��������$�~9�C�Ԋ5�H9���>A/OL81��L�$�O���<Ye�L*���C�>[G�@���� 'P���L��M���fCTvH�
��$�|"�=V����B�T�a�#�H��Jl�%wA��A�I\� �1���t�|� B�;�6�elڍK�����^�h��O�<�n���d��^�L>�c�ˢ=���`��B;C�4�*�d�yr(���f�j�ޥ70���ږ��Dd�����<Q#�p=,!!0,�3-�~�KSk��h8q׷i	��'	�R�b>�h��%L�4r#�����(�ZK�~(��NG;2�%:��UF�R�я����)����C�Ժz�-j-ܟ_L���i�5-[�-����?$�-0��'�Դ�I5 � HN���ߙ4���&V柈��4!�� Dxß6��<#���>$,A	�A[��yN�3���33x�Ƙp��0��~�I|y©�( �6�<�e$T|�Z �!΃7L-,eS��h�'��䗴 d>�A�[29JPd`V��53�1Kec0Ou0������t

�o���#)G���_�SV"&�$�.0�Ms�#e�J��O�g!�[�Wf�Z%�ء=|tY�Aˎ( ��O�O8u`�WN ����PO�Pq�|�l��s��c��>��V�4?����.J8@�`�<?�#P-i�0<)CC� M����%�(ʧDB�ĩ ��O�4���O�B� 8�'���{&���*�>Yφ�|0D�DиO���84��)A$��q��"���D	w��`� �F�D9��4X�"�(�fm�ä��Dsn�qc"O^���8z�&�j��h���ɰ�h����t	�x���1t�#2|��Z��x����<A���剶4��Bm�4���1��	*wNb��H!c%LO����I���P���̊n~���5��Xaz�!�H3
���O2���@a ˡR
�'���p����Ϙ'�M�B���Xܬ�� �0<B���'v�r0GƧ7Y�������9\�)�-O �Fz��I�I�H���ӿh<pAk��K�<�Đ�WB>ūbA�mA���s���so��yP5s! �6&k�!�w�b�&G����c4o�PWJ|���'�v� �'�r�'Z�L�����dLSf��@e��R����Q��a���\3*P�\��"P-D�5���э�(O�a)p�(:?Rܛ��]6.�#�d]ZҸ���̳{�T��TH�8cQR�@0�(O���'�P7�@�C��𸥯K/^����6��"��0?	�&�\{��z��B/z�l�Z��'��wtd�� t�\���.?$��'�|ѣug�r�$�O:˧:x��H��?��h�Qf|]����)k	��@JO�?�e#ڸLU��7*ΔAf!�t� ��)]�|Z�dC�6�X�E���g���d�<�*ϯoZ*uKe�W"f)q7�� �؈ʶe;�S�V�i��
& �|����7b7P�g����\����.O�O����R�'c����H�U��B�	4D$Dy* *W	�,1��ɕPӪ�=Q��Ө4�(�Q�b/	ƪh	�
�g�	�	ğ����AV�Ӈ����	�����u7�'9�$Qf#ЬvvjA+˕3����F	ud�e/h E��ɋ�7\ZT2��?��ݍ�V%���0�)T"l�ǐ�[l��	�d�9<I�i9S��zp�5���@�$`G9�>��OB���:_L�K㮃�l��yӁk�<	/���ߴ���|>O.A蠭M�H��C*Ǻ0�V�P�"O(D���\�]���`u��|ʲ�3��'�0"=ͧ�?�.O,�0�ȅ<P�X���F�
�dl��g֓!��� A��Oz���OF��ߺ+���?��OX����?(�#S�D�{�
��`"�-woJ�ʕ�F�Y��)��75CnY�d@Is�'VJ�fCK"?�ҍ��ʃ$�d�K�k��T}V��q-Y3�r���ˠ�
��F��Q�'���ͬh�S��<)n:�C&��?b"��x�i7n#=!���6��a;�3K��aL��/!�,iƖ�[�/S0a��� +F�u�	 �Mk����Әf� ��O��0���C�Sz^�A���8���'ҽ�W�'��'&��Ph;�#�F�-:�P��Ԫ||�b6�T�O[�U<l�%���(Oj|[���&y�3��V���;F�7/U�$�n\/Vf���e���c����(Ot����'b7�Xk� i�nV�9�j)H�NU9�6��0?�$M1ݶ��D+G3a$�Ka�\x�<�.OD�S�)�SZ���e�7&␃�P���a��M��?�.��	��O���_�0�t����"AVYY"d�8���DE�������5�1�Ѝ �θ�ҁH��?/Tc>Q�Cf�B��0vh��j��X#+g�Y	T���Ǩ_���ě��u�zxI����d��pc��\�+�t�ǦM����7&�
g�h���䧿�� ��� ,Y��حJs�5!���b"O.����،R��*�'�?$�	b���%�ȟ�Su��+NsX���`��)a�L(��Oz�D2�Y2�ie��'L�Y����i��;W$<rq*phS��$�t8��#G�F0.+G�6�1@��)�� �9��'K�1`��!�f|S�$@Iv�وq"?DT�!H��M ������UcH��H�p�򯇗kX48�r�b0�Gy�@��?����3��g����o�Y3�VW*d3G�I8L(!��[1W-���Q
+4@ğ�G&"M0��|"����g�B���
�P`�N'�H����~���OJ���O����?�����dJ��vǜ�8��6�� ���!�NM��eP3;
�y�B�@ymx��.�<6؍Fybf���0ɗ�n9:#�_�+���)w@���d���䓤29�]�aT@i�ȓ���(;��[��xRG��?��n�FM�c2A0e7���"z�v�:�OD�PQ��*z�M�s�"�ʌ��"O ��c@	���i���>#�PJT��!ش�?�+O9��O����O�S>2x��&	�O3tHI"��=Gp����o���O ���<R��:򄅚_a���A�3��[wk�*4D�A�� ��(��!(!�\r�'E�
7�I	v��H��
��M��a�&q�[B�j�htr�g 
:�A���+�Q����O(Y�j��8\:Ft�V�^9:Xc3�H�<�`�	`��5;�N��i����.�E~b�|�&\����k�?)�T�2Κ�tH�kት<Y��?�����|*͟j��PX�����)R��p:R\����?�,O�<֧�O�Dy�Sg�.E��%M�%C�z}�2��/��I�`��~*b'T8'�jH�B+I�D��*��&Dr���'\h!I�8O0��t�'@��O�0O�
GJS����!��J�J$)����f6�OR]֨�O���=��s��.�h�\c�~Q��f׎K�����@�䶌4�̟��I�Oz�4��u��'5��Or6O0=�p"�K��i���(E���e�"��'��t@��'���d �����u���<	�h��>J)����Z��%x�N$�?ٗÔ۟����7��X���"���O&�I�O���ą�?Ԋ��b,�|퀗d���0�CM�O��d�|���v���?7��*���-X���L>XD|���eֈ q�!o��<���֟��	?dQ  ��uW�'���O�A�u�ؐ8���ғB�N�9G,�(3��z�"�'�B�ϟ��JC!��'�M�qLG�q�H�[F��K��P��	�4~lPc���yª�?I��q�R0�O�"�'���� lуs  �t��b:����hӞ%
@�n�ȒC�উ��4�����y��L'<	��)L'V$@��*�yN���,VF��eJ�C�V7��ß o�%���4^���P?]���)_\�!�b����� ���_6 �'7�9�b�-�`���R�l5<� �4�?���?�����O����Ov�d�E��݈T��rt��Sp�� .Čo���0�	����	Z�	u�'[H,)Q'b +	�� Ũp!�l�\�' B�'��S��	Q�V�I��C6l]�^�1ڲd�Ŧ��	�� '�$�?��'}����M�3���1kڭ6���و�$/O�PS���Y��-�G��d�T���i,�	a�i>y&?��I�*2,���"�(�;�H#%�N�p}��'���4���'x� pf�&OYB���.�!p��J�'���I���.�����X�����'��q!�ȅָ�J�IH�Z.XH�'b�Z��N3Gݾ$
6a��vR��'�p##Pe~��{ �I�y\�p
�'� 1�ȓ�l�~"w$�aSֈ����8xZ�K_
z��� 4�Y>F6� )&}!E΅7ui��C�S?��ԩ��B񀡸4����?������ڬ8�OM�5c#�V_�_��Ā��'GB�c"�4|	X�MO	VdX	B0E�.sb�8�w%�)3P�ekN�vo�\�gG�rKJ�CD^�@��9��A�8G
L���#�3(<���I�B<�Ӕ�Ј��p���&'M���5����+ �!���2b�Q�q�ĈB�P;��|�1��!;�³K�:�mZ�r$ �
�w�\xZ�T�^�B���?�ר	;m��&�U�CS�(����O��o��b[�a��}���Ǘ=|�إ��5��x�D�rM�X���2ת�-8�y���$N���q�GL ?�U�#S���~��IԟhE�t�i� �C�'K(R���lZ-@�Լ�#� $�����������V;���,O�yEyB�p�L��	���ٰ̑�C� �D�O���O~�B�ߞ]�����O����O�
H�|(���%��Gp�,�O=�\,���h�@�mZ�mlԽ�w#XP��-ڶ	��pI�l�5�����b�1!p���MC��s�M$ZI�f N����~�seK=[T��=]�Wh^8SC�UQTWX=�Im~����?�'�HO��A���$u*�uR0�K�}S�uY�"O��ń�% l�8!Ğ�Qba�>a��i>��	c}R�ߕ1؄@�X���,��� �9�V����-p��d�OB�d�O�����?q����d��zu���W��]t��; d�HӔ���K#8�6 �+/r�9������ �ձS���!��a��=Fɫ2f�)H+a�[�h1��ڤ��O:�(�Ě+u�t��@�L�!f@�RJ��'�b��8��+"�˄(X+%n �{�OB�S[B�	�\T�YYcJ�Q^>���Wk��p2ߴ�?-O��0U��i�T�i�||�mκ^A���Ղ�2����H�O��ę;s)��O���.i5NB�`��"�:�ҺQ��1��E�t�H��5<���#��.+3�4I)�h�|@���' �rB�Y���M@�4���0���"N��̻d�-y��`5ʓ�Pe��4�M[U�O2�蚗k�,���<Rr�S��d<lO` 0��ZRJ1C��b��G
O�eA��ӐE�g��fe�W)\*��D�<q��.wp���'�"[>���ަţ����-�`}ȧgC��$��$S��?��t*���bKL&��s�4-i�iS��Cݦ��"�~��珮8�Zĳ$�D'S�P��$�M≘x�>!v.�3�4,��L��,��L
a�T�˲�]����  �f�<Lq����J��H<��b���h��4&\�O��OW�#�. `u�@�)Vi��J����ş�&���>� �C^��U�ç	�8%�4�$
�ў�Ӡ�M;Ŵi,�'!�12@�	=)~�Hj���E����J�9�Iϟd�	�o�B���П<�	ߟ��	��	-K\LI�m;,�JM� 䊐I�\Q6'K�4�hyb!IY�����5-v���� �
�dx��4(0 ���bCO<`U A��b�F�
J$3��}j�&
-󎐍~P�0H�f����$����	q~R(��?ͧ�?!�}���Fq*�͙�C?�U���	��y�m�)E�-0ʁR� ��7R����'l��+��|����.\�!	�.B9�$�L;
�0���-W�*t�I˟ �	��`�ӟ��	�|���)g�"���L�Z�H�'�K�tG2�B���b�X@�c���M��4<�B���$^:mr�+.����Ξ`X��`����9����/�.6�>orX���$��
�j�p��N(覩����Y6:D� �'8��v�g��ڢ�P/t%�%iɀv�m��=d��ct.�-'܈�K�-�;5f �=9a�i4�W�1	R��M���M�W��44�L�Y�HZ	��8�Q1}DB�'��x���',R�'��8�=� �9�+K$�v�1��5����t'X�;b	�<�P!�%O��49$���D!�0���=�0tK�LNI��HQ�c�
e��L��hO*p�8�<���ؘ�4+���M�x!��6 ��#Yrމ+�'�'��O�~��E@Ѧd��Q���X��T��R��)B ��[�>�'߆w��:��5�Y��4���� �<m�ş���V���-f��芚uh�8k���G0�H�A+g�����O��G&ޔC?((s�L��CH��:�-T�pq�U1g�~Z� �[U*�y���)S �u���o�I�dҒH��Nm���u� <��Av�
%Y_�0;� J�eY�2�D� &D��*O����'7�HN�O�.��|6�:�
�.09ڴ��a�y�!�DQ'p��At�L�h$ ���!I�Ns�xb�.�\~���E�Nk85�fAS�~xL'R�'Wr�$\������')b�'��'!�"1���W"M�����,dc�+_J��ӕEP$r���1�1�
`R��*�?�5��?&��wnE99@��a��[&M,BѪ��φo��<:`�L�<��a���� s���]�b��9:׬ۡ6��!�%�'(�.��$�i������Sܟ�}�L<�D��.�ʄJ��4PB`�W�B�<i��%6}�U%H�w�(Q��~�D�o���d�'���7;�`j��G�0�*��;(�|;�DyU�q���?y���?q��
���O���:n<Y�&V'{\xD��)ǚ5�V����	{"��!K�F���`nE3xm�<���	{�<Q*�%�	iP�M!�ѽ8��$Ӥ�Q?l\�Ga�
�y*pL�)z��Q���ɤYh�1uJT�7�psa�w]l�Ɇ&�OTh���#�>�B�b�$�zl��%Z�/V�C�	�^���� �N�6�x4��M+~�㞄ٴ��.�~}8R?�oڎukJف��A����ϞG��h���?�H�0�?�������K�X����ˋ90Vm�G�Z	*SƼa��J�`�����+�bE��c�lplGyeK*2f<��ݾ+��)%B���m�q��Ӣ�E&.��@BI��'.T(Ey�"��?Q���d�~j�����^�e��1Fݩ1�qO��4,O��qO��ЁS6��#�~0�!
Or�wl�p�5{��3��!+e#?G�4���<�WÆ�?ͧ�?	(�j̢6lq��)��A5o�6E���M��2��.�Ɵ��I�7@4��.כK�r��B ̶�M#[wRy	w�~�R` _��KpDs�(���[�	)�ʭ!g�S�'�cw������e�?5��S��z�s��(h�P$:7��;��O<�Ht�'D��ʦ鸀�/�F% ��]�?����m,D���%���<	��!!{�
��U�>O�Gy"��W�(�R�l��oex|�d�A
Y,�o�ǟ��ߟ)Yw�>����'1��'SJ��-����U��c9�%�u�A�v���Ν�d�� ����cUp`qM�/��O0����
��4{�a�,+�Ь��
X�Q{����$H; x��q��2R�T���%Ș ���}��B��$/�� �{�#B�$ax��� ��e��[`�����f���)�3񤐷�^�IMF���h�����!�$Zv�|s�%�o9�%b��\1v��r!���b≕Qz��L
Vo`4bI��z�zY16����r����?���?���Z���Ol��/Q� sE�׺)črr,�<{(��5b)a$�5�ä5�pR�s�'�B���D�Rؠ5�f()(h�؃��c��P�^�[�np`��X`џ�Q�� �!ZBP�cC$'k�!�C�m
�$�O���;��t�'#�؀�eL�"����X��ȓb��*����R�Bڿ����=�ֲi�BT�49�����<�	ɦ�@���fs� ���@��A�S`I�?���`��qP���?a�O4J�(��r�	���ǐ$ψ9�`�b 	�'���f(*r�=�26-�;�(Ol $I�%�����G&��F���<���8��ܹ*Y�P2���[�F�l�/�Q�ؒL�O�ťOzH��f�)�2�#3�%~�x�3�"O���0b�.��#�F�*y�
O,���I�����,�&�E�Qc�����=qO~����2�jɫ"@N�?B�c��'�ўd�2�U|�ɨc	�3V�d���4D�Ě����iiX0+���
�N?D��ٲ�˝���a�E��"���?D�$h�S�,O�mp��2m�t`X��=D��{�֎Jg���d���d z�;D����	�|(��'�K�)����&8D�p{4NA�A���!�D�$5�}J7D����Q�6D2��-;.u3��?D�`;�d�n�ֱ�w���=����*D� aҀ &g�H�R�	M�F �2#'D�huB_�	|�z�o�^	\Z�9D��I��4xpv	�����ٺ�E<D� �W��:e����5�w�6y�&0D�؋S�3<*��Jq���#C/D�4���]-h�r� ���.����O"D��CQ-�b�e	� �(!~����%D�����L�.�JeBl90��$m7D�41c������(@4.�
q5�)D�����	��^������	~�0�k;D�<�Rφ.��<�h�$�n��Cj:D����㉙T#���+ؿ�D���K7D�LR5n�b��|�����6�D�e�5D�Ԑ��Qs`T2��+�2q���1D�,��%R>�$�;���:^�$��6�+D�1���i�h�a��u��'�6D���b�W�x���<+��X�/D���(�:��aV��*����B D���k~ �`ֆz�4��V=D���V�
�ݫJ 5}�`��o:D����%�c�X��`���r�|��7D�phr��/���3��=��$p�8D���v�~p��k��Z�*�@�F6D��1&V�v�ع���?V�)S1D�)���6{�R����qW8;�a,D�hyG#Ͷ?A.�+3/T�
}��� j(D��ԩ�,�T�ri�7�P!� 'D�����~d���&��YD~Py�M(D�H�sb�7*�6]���2
Vp���"D���%e�6$y8=ö�Ͻ9,蹃!�!D��!�(Lud�s�l�6+���2r�>D�x3��?j�� zA*X�	Ę�`O=D����NT-/�0��-�~	2F<D��#!AWsO�� ��� Z������:D�tb�%�+]�2 ��:d�N���.D�\kK�13(\��cbJo�:%�dH:D�8�C���jJlk�C=v�,��§7D���)ʀj!*9�vB2z�$� B�3D��#�V=I���r�FA ����E
>D�� ���pn��!,H h�	�.}�����"O�D�ښoϲ�` 抭�����"Oְ�r��d���cD��z�����"O�Eh�m~�T��K���C"O�,�ZQ1��A@̀),���Qk�S�<)5��$�D��͘�kv�=p,�X�<-���Z�d�2I�y���tZ	��)�ج��CD� 	�b�0��Յ�f�hh`��Z��`n�4=�2��ȓ)ς܊��F�mh� �:��\�ȓ_��@,�r�T�ꘑ2�\�ȓrE����a@=U�@d�Ꮘ#'��!��u&|��&N�34�"pܐ݇�`�d�`�����4ʵ�&��Ї��2��  1h \�r��=�8���)�J��͚�O�X9��g��=�< ��.ژ=S![d�d�[�E޽7�̆ȓ�P�5�O�9,[f�R�w=�Ԇȓ �Ta(2�ځSj:���bQ�xA꤆ȓ��)8儔�+����G�Q��`��y��J���R�*i��J���܇�gF`}�S�LI��x����-�H��%?.�A#����2�$
!D�@��ȓ6c ����9�~Pڅ�ʖ ;X �ȓ2�^�ؓF�/Zr�s�
6�BĆȓE�\�)���0`�J�$�lw�`�ȓw�~As�j��/G
(+�!��i�4���jJ�̢4��q�0C$(@Av$Ȇȓ[�
)b A�75���E� �bu��f���f��,!�5��G㢙�ȓv^���0Ewv�X��K�`�t��ȓv�4�r�v`�
���.��%��&����n�Q�T��B��%�!�ȓs��M�p�,��{W�́6����\�U#��@��]��Xs`��YB�`+��	a֕K�BU��ȓ74����%D�`=Cs�^�[��}�ȓ>�p	w�۴8d,����Z,��ȓE6�4i�S��Jcl	M7
 �ȓ]yY3e� �z0�J&bЇ�3L6���͐��,Y����5��n��Y��$J9��|�u�HD�݅ȓf}��B2��+T�p��Ĩ+��5���y��Fѹ@�1��nX�^&��ȓhTy#AV;,d�������_EĜ�ȓ:���0�뀵�T��
b�< ���� �g�!;���,OyX1��S���)�����⍪S��Q��f����w�&�pʖOŤC7j]��J��p���I9)�0��A��id���ȓd}D���9��� �ؖv����T�a��,<Q��`k&�y���ȓl�J��+[�@��U%�R���x-;ҪQ2G{:=C��O<"�f=�ȓy�tU@gn&E���°��!5h]�ȓK3� �<��2�D���a.��`��B1�y�����O'!�ȓ�����N~.Ԓt��!>1ƭ��;�z8���N�Qۆ�z�c�9ƲD�ȓ���W��
$
 ���ǙPK�l�ȓe∩04
Ո;o&�`��,]�����im��e � ;. ��@�"eN���ȓE�Q9�I�X�L�
�� W���ȓ}��1��j���d�a�2sh����S�? lL!u�)5�т�,����j�"O���"+9����EK�9�T��"O|i�Sd<gIj��GD�2�٩""OX����K4Q�4*���$i���"O:�c�j����pv��D��"Oڌr��!�V4)�	�=/��q��"O��Zӫ:P�p�ȖD0�)��"O<̑�gڥx�ZҨ\�K�x! "O��B�G�b�C�H�^k�͹�"O��'�jw6�3P'ĒY�)�7"Oj����9�2Q�ԀQ� &j�h�"Oh�� �W��)IT��*\8a�"OZ9�b�CTl����3O ta4"O� JԬ��s4T�#kL�.즷�"O�]���0�nE���O�X���E�<1��G�+c�i`���6��fd�|�<y�*��bU�,��A�@<�c  �z�<ɂ��%p�ڼ�V�P,�j����~�<����p�H���+n����K{�<q2��>�
\QѨȩj���)�&Vw�<�W2��8
B��8r<I�'��o�<YȒ�T�<�h�J�k�^�s҃�P�<�3ȓ�X$�@A�@Wh�T��n�`�<�B�G�mq����bDg�X���U�<���26Ҹ�*�h��9R��*�$�M�<��%Y�v��|��Kk:����E�<�hý5(�������0sץ�~�<�� ֵ|�@�)�A���ATX{�<�G��T�it �@�L����n�<�@�,8.����C��ِ,V�<�UkV$~7 Q�gn�I[D䑲-QM�<�WO���"1��(�� �T�J�<aBE�-}�6]��hA�H|ڢȆ{�<!v@�
�����JE2R!#F�y�<!��*S_F9+B�ҕs+�
��n�<7Eو�̰
䄂�{��!U�N`�<aƪ]l�au�B&l�t�yb��w�<Qb���fC��K���(�����I�<I��'^w e ���� �CB�<�q��(P�p�v���vN���A}�<�E�Zr aS,D�����p�U�<IQgX�Pbĩ%c�?g
�M��N�|�<a@˚�"&�(A�ޡJ�����I[~�<I�h��(�b@��r�(�K#�w�<Y2���W:�"T�;}�C`��r�<Iˇ #,&���Ǘ_W��g�To�<�c+�(/'@�EB
�Z��l+dg�g�<�C` �x��X0a�WK�v�R�a�<�E
�8���F���t��F�<qS��&"ndK��W�'Y�t�z�<A����(�xdA�vf)B4,�s�<Q%n[�`�Yi���q�j�0 Jj�<ɅĆ5#Thр �m~e��Jb�<�%c\�(\9���V\���h^`�<!��%��p��M���+`�<QT��pE���Q��2��v�<�tcҋ{����H�D��Cs�<q�oO5�<!2&N�'{͘thֆ�U�<���-d����1� �L50q�l�<I�Ò=}#��S0��j$LQ�7�Hr�<!'�~zX��R�_��MI&�Qo�<Q��C�f�:���K����T�n�<�tͶ�1)3��t����#�g�<iŧKSU�@��HB>Tl�����z�<� �� ��"P���(T@��,���"O�$����Uޤ����#j�,���"O�D�N�DX��R-E��!��"O�}�OA���˓�T-k����"O�,�C��A0(Y��
��N@B"OX�Ȑ��5X����'/oT��"O�4�]>^�� �oA'fSp؊G"OV8[�RvR���D����H,�yR[�3��͸T�!�#�%���yO�m�V��F)�:
~$�����y�Ti ����Ԩ`�`��'?�=ifїa1� ȇ! �u��i��'R�C*I�L���Ѕ�J�kn8u�
�'���+! ���������s��I�'�T���FG%l�vl�Qm�m��X�'�^h��Â6?�b��D��d/�t��'� ]��,� B HjD�U$cF�M��'��5K��F�JN�lST�GIQ��'�@	ʅY� }8����@w�1r
�'��]9U��
�z|��!��g$�k�'�dPs��0Na��.�w}�9�{�ɫ�R�"�#��k�h܁s�7��.\�i�bb\�p�$�y��$����Z"}Q%���"Y (�5`�=R����ȓ
K8�r� �_ ��2K�cZ��ȓS�Y�Vb(5�zp�&�4i�u��;8Ȝ{E`L�J1f�y$Ο�,I���ȓNp�b�䌞l� 5
�m�0u��k "��@��{��t䪌�H�̆ȓCo)�P�/>�ԙ�χ�����ȓ_���WGƂW��]��qoԼ�ȓGfa����$�  ��H.*yΩ��T�*u��Ė%����&��*0��ȓH-��#�i\�G�t=8�n��O�`	�ȓ�AZF�Q�А;�ı<ln���]^��³F˹  ����7�(��u� !����k�@;$�P�f�<(��D���@�/bڂA�!%�Lk��{������$,���E뛀M�5�ȓx��q�ص>�L�@3( _|���0�`�����BK0a袊��wv���@Kp��Q�E�`�F� �jԔW'D��w\��2/�kyا)�-ݬU�ȓ!	�Y	��E�Q�~�r��.|��݆ȓZB��%����9�q G�(��4�ȓP���%��E��oP�7�tC�	�#� ��W�56쎔K@�@��C�	J�@u��B�|%�n�"v�C�ɨ`P�qBh_ku��Q�kP�C�I���4���eH��b�c��لC䉀1�.��a֝KD�B�U;T�BB䉊r�$A��35��|zS@_=.B�	 )�j�02�ɉ'<��B�	J*��l�?��Xj��S��C��2.�P$C���0:��"��/BԎC䉪|� �XW��<Q�1JT-�B��(!;����h̹q��M"_ԊB�I�2a����F������4�zC�IZ d�p��;H��OU�C4B�	�o�j���d�l���C� ��8B�Ʌ��8����0�0˚
N5,B�	�O�P��?t��p���Ǥ��C�ɌH��j�G�`��w�ǦX�C�I��:���*@=ٵ�,%C�C�t2�`G6D4�b��C�P�C�)� 0)pDK�1:,(�2���A8���"O ��	��UBj|q6(��q"O��!ëܲx�i	�,��TU���"Ol���¼�ؼ����1�<�"O��aFM*Q��B��N?%"d��7"O���g""�:Q2C"�'uk.��C"OH!cc՗H�LeA���5,�>���"OȘ9������@f��e�2��"O.��$�ƶ-d-!Ģ�� ���E"O� j�.��j99�DϟM���"OZMpVD��_��ݲ���%��U"O��R�AXeah�P �O�m�"O��ڂF�*zYr�j
�'�ER�"O��"�:.�������Sp~��"O2p����,7t��2���Bg�D�F"Of�!��[.,b�h�èޢ�
e(�"OJ01	�h�#S�V���"OrM��m�<M��a���E�G�Zyj�"O����!�d��K5e�� 
� �"OX�"���{�6���	��!s<�"O����5b�2���o�
oO���e"O�B��J�̖*5�C�EF�y��"O�HR��Xj �@kV&n���a`"Om�pC��$�}�f
��;SQ"O�x��ڼ]�<�2�	+���bQ"Ox)Q)��G���7ʣ9��̠�"O�`��Lв(��y�G�\�9��"O�)�Ă�+��� J;}uJ�8�"O�ĺ5�ڶI*69as�L�\Z��C�"O�< &J }��Q���P3{6Fe�g"O@9���� �~d�d+ w-�� u"OJe�o�/	*A���J-��@"O�Q�%/�8#��L-i8*JAl���y⮜�M�|A�ǫN�j�TAQ�ߟ�y��R$_�ar�
S��p�iF/�y��^��-�F��`��s����y��K�!��1�B�,�� ���G"�yRG��znxs@.� �B�U��yBNS) J$Q��Q
�:U��h �y��ڪ�j�ٱbW�&����y��g��H
���SV�pP��ȴ�y�ˎ�|�X�c�֢F4�p�E��yKZ9V�N= �	Q�|���PP�I8�yRoԠ.~r�[��8
`B	S�y�h�}rn��C�x�p����yREW"?!,:T�	;obޠ��`��y�oO��=��Ƈ�g��x��nV)�yr"Ѿ%�U�A�f�� �E��%�y2M^T��z�EN�a^�pI$�y��C;/��0Xpm�H�82��y��]"�eX����ڡ ��)�y�˙�2�¤����	Dض�y2��4���@
Bp5���qg��y��`���H��/~�|0 ։V0�yr!7s�\�#�L۝o�\t:�]��yBH�Bli��֛nuvTyWbȃ�y�F��>��A)rQ�̞�yr���IȔ	�Q3�8�ʄȕ��y��-���"B�^� 5�ߘ�y2(�R�����Y�&O
�QWL,�y��� �4RQ�L�2�f��.�y�M�"���6Ԃ	�<3#�y�H؈q��dc�Nܚ��:����y2H�<��5;'��jcX����y
� �R�m7n�h��N˟
7`�"O]�G��?	:9sP��J��ST"O�A�$�G5:�+�"�5A���Q�"O��b�C��CyH��bbH��H�D"OҠ�2�A9,f��F�@�?�s"OB1�6��7��1Q�	P�2DkF"O��3�
�<� a�	�[���"Ohx��	��M@��ӯ��="���"O`���L?L*QI�#I(c���B"O���A%ى �X�0��#�01�"O�EA�ϑ�tx$��S!�@媐��"O�03�Nߦ /�Y���K ͪ�i"O��d�>�Va3tmҗa/�r�"Oȁ���;[�y�#^g�D��"OR��m[6m�����>xJ�"Ox5���2�Tyq��	q�zh(�"OnY8���<�>I��3%�H���"O0�`��	��9�7�ې���+�"O>�ɕ�<M�V��e��+EՈ�"O���م���v�c�,ѻb"O�1� ˕�>� T˨Nμc�*Of��% ��(���4�2d��'�"��0LEy��e���2�R�`�';�S��m|Z��rLJ�+�N b�'ϪybA��m\9e�܋T� i
�'qVLA�����y��+��_CxUK	�'T��zÂ�(\5�)�\�P�X���'[0�r��>���N�[�T���'�f��V��|H9�VOKX}����'}�`�4�Ӭ{�r9k&G٦��C�'8e�n�M��%AH��MOpS
�'Lᐡ��z�
���=3D�`c�'?��!��.̌� wdԠ:��'8fb��5_&>�`��H�"�RqJ�'$*��T �/(F�;��J$!��'(,�n�"�p��)Χ7��C
�'F��1��4}L1!��>Xt:  
�'���D��N��4�p�����'����EGC�����eT�ä�h	�'�T��ℇf� (��T>P���	�'�b��C���k�� p\�]k�y��'��Q"�iK.	
�Ҁ޿Y@<X+�'+�=��eA��(�Yb�W�S����
�')@��˟g(����᜴`�̽ 
�'�� �Û{��
4��b�^���'-B� ]s���Bm^�'Ր,i�'Ζ�����9@<pH%M\X�PP��'C�i�ӯ�(��80��,T��tS�':�t� ��-�|9�S�Y�E�J�Q�'�J���/�>9T�����qA����'�D8A
��v�┻�#M�}�$��'����I�>O�F�{ )�=|���'n85xqFǠ߰H�Bo<���'v�t!��#��Ak�	�k�t�#	�'/(mQ��5qr�+�v��	�'�<]:���z��eR-%�t�)�'X6l� @��NaS�N�*GlRt��'�,Uhj�6I+�Ps4"܆z�{�'���I��)n�P�w'XpҚ��'�NX` Z�Z*R}�&E�7�\�yҏ����^�ov��+�c���y@	1�p�Z�f��a�� �GW��y�B� D�p)yT�ϰ����*Q%�y��(lZ�k44)ܞ}"`蝥�y
� <��X1�Z����Ժ2� �br"O�}�u�T;"@�� ��z��iR2"O�q�u�E�`��l�Q�Ťr�]��"O<�ҏN�	� ��آ�E̫�yB� �#���&�� jƉj�ų�y���Qژ���6��9{�A	��y�cs�y��Ԥ-����� ��y�վg�ⳋ�Q����K �y���r�`��*	��{����y�g�_�\���O$iT�B!˓�yr�N��2b�Co3(h)1���y2$�1j�m�0Lױ`�l��Gc���yFQIIt4A�߻'���pW#�y�-�?dt	��*!L�Sh��ȓ7��T�K?;��5
�eB2�Xh�ȓP�@�H�h��WF�c�MW�0c�؆ȓI�,y�uH �!*���h�dPE�ȓ�x����X $�3��w���ȓU¼%Å��RC�|�GQ+F�نȓhVٱ��.vtr���oʧ5B}��Im��ӏ�2��ȪpFܛ�l�ȓu�<���� �v��G
���@��ȓ��T��JO:U������Ҟ]���ȓw�b%k԰q�2pB'��0G��)�'� ��j~^�a�h��4��{2�NJ������p���[%��=�6(����	T�0��ăoUL��Hi�I"%F�"Y4h�h�A2"���ȓ3Tl(�E/(��]�t�W+uL���}<����@1TP�� ��\<��9t�*���,�<�a�ᐛQ�����}�D=QwJ�*Hf�E	�Ϛ�l�΄�ȓVS�L���;@�6|�(D��c�����U+?*�ðJQ/F����)B�ࢂ�;$�¥S&�ɧD�V܅�T�؁$�>dn`Ӵ�)���ȓ����"�	3:�N	��ʍ�����-!�z5R�S��A"p�$0�H��8'����;.��H���WVVY�ȓ@�!��C�3�D�Q">E�ZI����ճ�_�x�N���SP�������!��>��UӅ�T�0Alh�� �
M�.�h�H��Сe��5��<n`���(a�5S����|q�ȓ]��݈G��N͂�@F�2خ-��{lX��'Ϳ|u\���{�B䉷N�V�!��:$Z�is4jF<��B�I/1�4Ȋ��  V�HlY)$ޖB��3Rᬙ�$�[
lg�t��$ zB�I�a���{��-87�5����%6/�C��:y�h��cn��{_.�i"�M�:��C�	�|Ne�e���v�P��lʷS�rC�I9?،�I���8vI�hjC䉁D1�k�Ė?\R�e�r��|�,C�I>D� �I�1�!�l�W��C�(���v��NB��+D�;��C�l��5����l�$�+�,ņX	�C�	�?B�7���*�Y��'_ߠB��+���:d�T�$p�a���d�B�I=��k�i�krt�$n;_�DC�ɛ8Hm�G@�.AV ����~��C�	�v9q���H.$Phs*IHv�C䉧=�!˖��%"���H��B�	4�����DA4���qL�>(�B�s"��P6b��IK�ɝ<��C�)� la��e�3'2�����X�p5�"OB�YщJ/����=f�� `"O%	F�]`��i����7'rHj�"O��	���@�fB�4+&��Ƀ"ORV��5#���BH=n��)��"O��AI�&��,qS�T1K���"O"�
���-��aB�X
�d�"O���\{c��`oT;Z\�:b"O��[2���QkBe���1'�2�ؤ"O	�k˱
6PȈ�l�$DY��j�"OR�qse��T�F�)�� H�Ρ��"O���� �N�d<q�$�G���"Ore;�f!�}8��˹S�H�� "O���t(@
]g(1hA��t��s"OD���o]�I��4��"'yӌhXP"O�	uG��5ӄ�ys��e�r}�`"Oa ̊L�ؐ��78H���"O��B�A�6� �v��){�Jš�"O�i8UЁmD��2�T�Y��hu"Odz�e�6Z��	��^�0=�"O�b���G���	D�7Qޘ���"O>0{��ob����d�|���s"O\tA��W�B�HU�#J9�\eR&"O:�p�Q�b!��+��A��Ř�"O>�a�+�V
�ѓ�@��4�0�"O�� 6��&fh�b��Hp����P"O� �dLU�i�����m	����J�"O������)�^�!�G��^��e��"OY�W�B�F`�h%�%�rs"OP!Ю̊5'f��@��r��Q�"O&1�m���4�󣂗m&ґ��"O�в���5f4� �B�e&�}{�"O҄�N�K���ǁ�:���"Ol�A�F=�tF ��v��	�"O���&�'��5�c�ޱprnL1�"O`��1�T!�0�%I�' ̄r"O"Q��kJH�3h�Ǣ���"O~��� M����蕁T��	A!"Ohe9�S�TB9C�GO
b̚�KD"O�%���76�T<���_�b��!"OF�C�o<4N\���
��81��"Ỏq�iK�Bԁ�����"\�"O$`i�F�^	���ˍ(Il���"Ov1�w!ũ����LH=(;��!"O�<�/ }�8�+��q��"O�h8q# �H��+��8�;"O6T��,C'1 ���E��r�S�"Oи�p"��3I�x���0�.a�Q"O����C��H��-�#|�8��"O��wl��M���S�bL�rY��[`"O����NxBR��8Y�M�a"O�!�f�
T�|�s�Y�dIA�"O^U�E�$)L�ېl@�7���x"OB�$ ��A3c��jmz��"O���	��H���֭S*^O��"O~�!v�16����L�=��x�"OR�P���'�z�A���q�p:1"Ol�3��G (��-kAFW� ���B"O>xz��ȏ�&5���� zz�	a"O2�J�ϻw�Q��bӗm���g"Oh)��a�^%��`�Y�"O�E�EH�~#�ɓ㇐m��0�"Oj݉v �8w��e){�Rě"O�Hʶ���J����mE"O� �I���q��5#򂂥6�
�'"Oxxc�c�)uVT���� ��ؠA"OV��q�_6D�țfL�7B�~�@�"O�*Qm��:^v�X�kK�0�9�"O�ĂV��/M���cc�\[���"O@m8��e��HAlʴb�|�"O6ICО:� `�#L�^�"5	�"O�qz�E�N���g)U'���)�"Ot�Y�I-QA$��
xɹ�%[��yRK;R�ԈH$˅�K�|��K�y���`��e橆$=�\�HL]#�y��ya'�r5(�#���`F�M8�'�@����	k�H����\՞	��'��N�s�L�c�����q�B���y��I���PΨ	0M���K(�y����7�$���-S�k�A4'��y��
)ee����H+愑���y�̺9���R�.<:���^$�y�;"�.����]��@A�Q)�
�yrƓ,°��WK6tHP��K��y��ШY00k��
K�C|���"�u�� __.`1+���K���
0"��C��ؽ"Q�U�RL�ȓ+&0�ďY�/@h���ԍ }:9��(g���E�J�8Z|i�Ny�:܇�m���ҩ0id��q��4��B�ɽ�|���m��H����E�B�I/C�&`�  ��I(�(�
B䉗>^!��ꏽdrb�3��� w��C��'6�TJT�MB��&C�.��C�	?r�ԉ��@�&�t%3�C��C�I�b-*�v㔓!���ѐ�kʼC�	�<"���si� ��S��{ �C�	'!E2(1��~B|�ĠI�P3TB�	�;�q���Ή$���G_x��D@���僇��wbBS莫|!��h.h��?��ц@Űd&!�ݡl�����M��1s��-d�]�W"O4,�b��%q�Ɏ5y�x3�"O�ѩ�d�5F�١�S�*���"O�y�A�X4zT���L�� yG"O˲�ړl�~����Й�0"O����,�
BzD��#bν9����"On�Q��@65N�h�v���(LʘX�"O�+��_M� �+�h_
o4
��"O�Ъ�(	9d��٩��Z-���C"O�!P�F4��E�gD=?��Q
"O޴�Sf��*]�!E�P�("O����AND��%c�"��(Jg"O8Űp�.�~�cU`C�}`����"O�YA<;'�)��] eI��"O�x��΅+i:,j��ݲO���"O4������N?�0p6�%}���s�"O�9PaZ�F��2K�;m��X��"O�@���4�� �l�	��(a�"OXT+K��yN!��J��F��s"O@���3e�R�C�JP5|dy6"O��e0�d  #*�)"v�dB�"O���g��%��)7�}A�"O�l�«�* l���'V *�rC"Oh@�$T�|��(Ƿ6�R!��"Ov�h��N,��AeG�����@"O��8B*֭����c	%S�I
S"Of�e��{(��Hт�9S=B�ˡ"O� ��7��d���a�`Ǽ~.p��"Oک���<(V=����"��xp"O�\Y�DҎ-3���F�A(���T"O&M��,�
-e,�#��	��`��"O\��w��4O~�)GgJ7U�� "O�5�U�)���(6�l��l�"O��ȥ*W�Q��{e`��j�x-Y�"O�� 6O������;��H�"OD�.�:�j�ͪ
H-�'�S,�!��'2v@���ϗW��7L�:`!�d�8NXቅ�F�uk�`C�J��f�!�kV� �J+\��cQj@ <�!�L&=�ڔ
CH��mR��\f!��4,<�	J13ObX ѩO�(Z!�d�.@\��)U��F�P�*��$�!�N,N��ZGd؝s�T�S����l�!�$�}��Mq5��&KL��Ek�.���DT!(���6���D��ʆ'�y�CZ�P@Ѝp�d { ԈbEa�<�e��?u2@{��?�.�5N�Z�<���2Ua�T�p���h�(��m�R�<�Dʈ9|�A�C��
1��}B`�s�<i*W�1ˤ�
0���WeYF�<�F`�!	�Ca��v� ��e�C�<a��M:T9�U&V�!{��)'�BF�<ٖ!I#�f�S#�`����A�<1�M�9q�ƙ�qˊ�U�|�[bHH�<��I>[f
�n�5!ײAK��I�<�qE_��P�5�HU4�AhGG�<لe��H�/O�t��r�D�<���[�)r�,	�	S��a���T�<q��	�%��e���N��q��ZN�<�Q*Q�X�m"4��[7J�� hXA�<)�K�/��8!f�K�Hr� (�b�<a�j�4�
�#�Y�,d�ƈw�<	�o�:�z�	1�" ��K�o�<�E��fo�h�%�x�차3`�Q�<ɤ�^9r���e� �T�҅�EL�<�s Ѭb�B1CAk'���6�G�<��$�?'�40RH���θ��y�<y*�'i6(�s�M*�v��t�C@�<�`��;f���da�
;�=���G�<����!Lr��`E���l@�1��]G�<YG
M�8P!�џ0<�Q�@CG�<�w፼V.��"�A��)����N�<AdA;:��l��YQ���@V-�M�<��i/̶Y�@�,���z���H�<����	W��q�FT�����O�<��@�|��8�Rz�����~�<�1-�?[ģ"*�ODA�+�y�<�q�۟x������w�`��mw�<2d�"@���ƒ�i=D09��q�<EIE4Mˌ���Ǝ�"U��S��k�<�A�גPD`L����8#/��3V@]�<0��"=	\���D�:]�h�g �D�<ƀ٣9�R!*��Ug�0��M��<�2OVn'ޙ��l�yD"� �Βx�<�kӄ[��3���r�9D#�q�<��]�v�4aH�q$ 5)Zh�<qE�*S,Z3��ؽ�@� �e�<9��U��K-�ȑ�@��,C�I/P5��1���@�ڸက�x�C�I�Zt@�� �v�m�4;�C�ɀV��B@XM�P�b�ځ0�B�)� x�	4��o��L䤀P��#�"OJt2OF#�^tNH+u��|2R"O���jăF( y�E��~�h�"O�ѩ �R'q���gjE�Y� �I7"O�Z��F/>�����n�>qq����"O�����ո=]�*�	'U��2w"O����I�V(�Y��K�sRz-�#"O�eJ�!ȑF�MH�����Xe�g"O�I��O�x��Ԡ��E�Ns�"O`�9�CH	:�̪y�:5�"OF0�ߣjK�	�GjJK�"O����K�1�\���qf�	�"O���jD�k����g�8��Ad"O\1j���n���zS&����b�"O�)��BBVeABeG�{��	K�"O
�ӥ�3��`�⒒���A�"Ot*�d�#��ARC��>@.�=z�"O��iv�Շ}�~d�G�5~7�5D�Pbs�Q��������" c5D����@��
^������W�
���>D����,�#U�z�a+m�����=D��c����t�ۿy����H>D����B$X��$Y��D$�� �<D�����9Pj�J5�Ԥ+tj5D�TR�œy���;3���������4D�����1|�&$��ұH�tXQ�&D� ��Ε!Z��d+���0 3��AF�#D��*"'HE�l�*Nv��P�Q4D��r����%K�i{�K����a%3D�\ C	�)%�\����&I���� 0D�tB���%f 0�k�ũ?���R�,-D���T�T7��ib�E41��§n'D��Y���-W���dk��\%:q���&D�h	���7ؒ5��E`i��@)D��Ԥ<�j�ACLI��M�$D���*߸�����)˝�@����!D�@�E@�6?��m�����Mj5D�@���:�F�������jh��L'D��@��:�<��W"��U�.�K��!D����&<��7螱n(��qW�=D���� \�*h����1?�y9�:D����iF2P���x�ɐm=��3@,D���Ti�S~l�dk���5��m$D�xQ%B�1�i��>5,d2r�#D��%��وQ��4��)�և D�+�fP,|�L䋀#ȋ�r�`gD D�s�G��f���jT�
�V�v�Kg
*D���2���B���H� ���s)D��;��с� �f�\s��d8!�1D�4A��/}8�,A5�1�B��m�Y�<i�%�A�q)4Mʳ �(i&��S�<I��I+8mo��b��aQ"�֩�y�Ė�g���)�0n2�X��Ԉ�y�A@4#�xI�3'H	2��� M��y��ӓLt �2���\�R4�Ńڻ�y�A �h�����%["@�QU@T�y����1Ӿu�%�.WVia�Ko�<�D�s�Е��L�O���Q�i�t�<I�G�?Z�����O�SE��1��y�<��-<����V�5�ɐ��w�<�Я�)|���Fe8KT �pTq�<����1�>IS�ƕ�Ja��i�oMn�<閨A g�֍R���<EP9��j�<Y7��ch�CEύ h�2t��g�<� �X��HB(T�v���눊��Y��"O��*��E>F��;���-x�ؚ�"O�u��\@�{���))[�Ei�"OH������\���I�\N��P"O�D�w���\$�H�C�mD&l�"Or��7~R�]+�� `���"O�5:�&��J�u��0�����(�b�<���:^0ɂc)''u:u�v�_�<��>C
�b�cY(��=�@SD�<�ucؽfh�U#�N��F�x�Z$/MZ؟$�2��A G�?|,(3��XbF*D�\��)�r<�QJI+i"eY"5��҈��P���C,^�c�9�4-��"OT`J��z��Cя7�B`�U�8F{��iD.f�l���.F�8Y��k��#�!�@�0'��	'*����8A��,��?�� �V�q��]=O�N�ҵ�R�a&8��Y���ffՍ�"DRO�tX 1��O|��̈́��;��(C��p��'��>i '%:䬑�hɟJ���x�<q�+�+ׂ�#"��&��(GƂq}�i��OE�O�>�:w( �W<�C��:�6�[� 5D�L�Q@�� �L�����L?0�8G�3���<��+�YFĜ*�G�	4��	�h
J�<A�Z�X����1cG�9��Y�7�!�$��c�P�9�nǎ�TYl��o�B� Wh�!0GŞ/�p9�R��42�C�I%E4q��/��3�J�1T�{\�C�	��HLP���8u���)��ΰH�C��
M�J���d
�4J�X��nѷ,��C�ɶp�p賢�>4S��q�
L�`W|C�	�_ulT��/ 9�N���Ȉ\NC�	�1N|�rAÍ~o� [�`H�,�6C䉆g>����F�� ���Z7��I�C䉕qY���1�>���E�{��B�)��cd)H�S��M+ �m�B��1B���[�Y3%�։Xc� 4UlB�ɭC��P�S�A<E]ik�H�3B6VB�Ip�����G4ud�4�Ѯ�2L*B�I�u����V7 ��}��N9mB�I" (:��S&mΐ1E�Qj�0B�2uz���J;y��J���91�4C�I�>�\X!�3>=4���݈D�B�ɃS�E�,N�4b�����B�	�):�YiH�."��L��B��_`4D�EfO�[����(ߴ3߂B�I X�� �N[������!g	.C�Ʌ2��A,���ʽ��%�4n�C�i�N=����k�Vu	�FH$r,B�	!~�x�!ǧ�<AJFm��c�?�B�k]自�7 }2v�#i�C�	�mf��6iF�`�ɮ'A�B�ITT�������$\�S@M)'�TB�HLj8����m���[A��31_ B�I�q�v�[d�رo�!�q"��C�	�� D+��
bص��,����B�-AR�p7��t��bG�ËulB��&Y-~@��%�v������U�W�B�	�_L �#��8<%ޔ;h�L��B��53�T	'�˦(���Y@Ğ�P�B�	!u�ZP����$)�L��ЊK;�C��a�����.��&$޸�B^��C��+m�*s� �5GԤTP���I��C�1U|i�v��8n��� ��:	�C�)� B��vňI��P�HY�:���"O���vC:vwc"G̅[��X�'"O���᭞�N�-��/�� ��"U"O�Pq&c kaf@0�ǍO�>�Q�"O�TP���=��Q��i�G.��"O��0�^�M�@���M;.]lRq"On���)����(V�PXN�Z�"OP����,���r&�י9(��e"OZ�b
�*,$]��X<p
)B�"O�-��	 E�`�@���,T���%"O6T�Sj�:�ֵ���׸��EC�"O,`�cD���޵a%ʃ.���!T"O<��-ԞM�H� S)A�r�f� D"O~��'1����g�ju���7"O��)���:��҂W]"c�"O�jťC�U�
T)���\��5"O%�$�<=�2L3�ś�?jl=�"On]�î֧Y�rm8��=��Ѡ�"ORpSB��d�py$�2�"X"�"O��BE̬nj<m*��s���u�V�<��^�LeB�D��<�Z�	G��R�<A�"_�T��� ��m��I��J�<��K��|%��G
	�0L���a�<�ҩ^�3I$8����6Z����e�<y���)NJ2�Di�YKH�	�^�<�A��+vP$�1HM��zЃ��Z�<�e��Z��X�����&t�v��{�<ٶ��)_ݲuh�!]1�l�@D�L�<a�F�+�L�CеPa�кt��P��N~�5S�J �7XL0�Bg�;�Z��ȓ0�ĠHF�N�>b�J�� @v���ȓ+S��Q�H#1~�e��+��^��ȓᆍ��H :��v�Z�K1�0Ex�'L�u�EӦ��~Z��ĒūөR�5������Lܓ�?i��/K� ظ
�x���gc��b�,SD�<�` 2˛0m�d� $E�k�\xEy��ȍ���xQ͟-Y�Ĵ�S�ɣk������K��c!�יl2HУc,ǣrBby(��d�,qMo��h%>�oڴn�&@�kɛ@R6��u��Xj�L����������9>(�Y�~(Kc�X���ɣ��O�Uo�M�ߴ|OL9��c�~�"�K��N�vU����a��Ô�i��Q���?e&���q�
6��c�ւY����`OV��x�H��D����%�Ţ<�duڂh�6�O���h2�� ��9eE̘�f�DE��	l�)/�Ĕ"��Ńa���®�!5�$,�R��B�@T$?�ؙQF�� ��mr�p��F0E7�H ?i�D`�L�����i��I��(���@ѓ�i� ���(�'.��� �1ct�4շ	�Ipw��a� �EyR�vӆlZ��D9�4�?q�'�u	��DH����.\<:iÄW�4��˓9x\�$�i�ayB��z��E�*\j|��e��5�W��oK�(� E�Kٶ�y�����E��249*H%�|�ׂ�\��$��ƹ&�J�z4��~LTqP��	�v4����JH7w�$� P�q�J�ɎWH�t��)e��%�p���1<�">Lq�I:�M��x��'�_��Ӕ눣AgD<���/V�T�J��1}B�'=�a���G4<,���Y%�H�j�C�Ҧ��4�����'��dF6k�A���X�;�`9{4'�kpT;A�G(.Z����O���O60��O���OrdB��;!?`���C�x�tu(U��k��9CJ{	p<�N�k�in��S<�<Q�F����� n���O.��|�EA���(��3J�ޠ�����K`���m��Ja�`�	�,$�`UM�U���я�2AP\���J���MC����O����O�v��ɜ> dL��v���w6�9C�'�L�h���+vR�PS�Y iL��+�'ʠ@�R�bӞ�{<~,Q����8�)�% �=ʄ�O��@�0��!UqO���А��)Q�];V�J�JW�d����#��Koj���� '�@����91�	Wc+�V\^�
C�(���0��D!�v���)=�Yp� ��=
a����
IP.���QY�'r�<���L`�P���~:�bRJ �)�jU������Ǡ3 RR�薧�����	�d@BRס��{�L��>Aشr^���i��#�C9�T���ݧ+v0؂�'�<(p�
v���'��<t����៼���t�z�W..���d\�~FrpU,Y:H�©#2GC�2H"A�E�J��uW��W���?	��&� �{�dےS�8���ϑj��l�0M-f���LP>n�ܰx�뒌/M�{�ž��vjC�\� 
���f��� ۗ�]�,-� hG�i�ڬ���-�<�S��MkT'͙W�ڶ*�R�ri��f u?Y���䓠hO���,e^�F�V�f�Dy��G�(On�n%�MSM>y�'�u���N3��UIW5N�ٛ��@�;r�O�����$g� 8  ��J ��cȂxh�ݻ4�7�y��F,<L���o�Zt$�N�ē	�Ex���Y#YxHa6�L���Z��,�yB.K�]���0�F���H�m],�ē�~�+0,OX��I˃4d��"EϐS�|���'&���9tXM���#�Fbg�֑f�!�D�*�t�{�M��O�أL�!D
!�D�0�X��*��q����g+[@�!��H~
�Is쉳T�ڨ˅��8~!��*�f�����
�fQ����U!�D�?��ܺ
T�(����m�+or!�DЊ@����↑9Pul����\�"�!�ĝP�A�A��+%
��r�&�!��D<G�8t*��?�^�*��MFl!�$C�j��-Q�h�% �@�B��T�!�DC�'J*��b@��_nP�E=9�!�dT�90B\�*��l��T�U�,!�!�DF2�z��"�
l���}�!�Ē?^l����\�=�u劚Fd!���2{6,��CXZ����tJ ,6!�$(pZM�B���2TK�I�.�!�� D�p�� ��l�b�Yk�^�R�"O���,ޢ��Vˏ�r_B@�p"O�$2`�U1e�t%�E
-N]����"O�]�@�X�
A&��5���;,h�{�"O�0���2flx&��+s&�@�"O�����@�N�څ�+Ϋ:W\a3W"O^J�ʞ<!�:t�`�CYtM��"O:i�b�Y+5��g�ͯ.:��"O4�X#@Θ(�"U�
��
%�)��"O��B��ڲd�i�:#�����"Oҡ聎��,�I]�B���"O  �&i=�,(�f��b_����"O��b$� �w��D���'�qE"O^U�n�����KR%
�,[5"OFM����3�Z �&�USȹ{F"O d�e�ے}s"5�TB�26���(q"O:b@Oқz�U�D�#���PD"O #�f�'k\�5��T4z�:�"O��@֝�&X�p�z+��"Op\7#�1U�mc��J!�r�"OzU�8�"=!�F�!
�`�� "O��3$���N�0�ĥv���"O�܈�/�f����c	R{�$�"O�l��O/o����QLR!`J�l�p"O�<�Kξ,�����kA��X"g"O
=���JgFu>>V�Ad�W�yd�)r�\h��+غv�B1P2@#�y�J� C� D�#��'u�6����A��y�D�,  �A��� �A���'�yBe%X��p�gJsDe1���
�y�f�=X����"�� �d�q���yb-�����g�!uR�3@�Ŭ�yr
��.������r���Zw�P��y҃�2-��<�3S�� �"��y2�E=J����0��>Y>zM�f��y�M�zJ��J�W�\�����ƽ�y�I�+�0��"���:0��,��yR% 0c�6e��˿L��rsc�y��6S��%����Y�-�y)��g�e��l`Nՠ����y�+ȰO-���*�0{*�h�MW��y��ۉG�ȳŮح}Ҕ3��ɾ�y#1@��*$G�m]��!nؓ�y� ��5#��� & 0N�̵�2�H�y��NVz����f����[��W�y�C(W�����֓�� �(K�yrS�&u��*�"A=}��0a#6�yB$N^8@��_�dD���y��j,��Fg��M�T����y"$)I�8���F�K
��"RB�yr��~&$t1g���@� ��1OI��y�kڽ#:��-�)aDUZ���yr)�f*�}���U�,�*8f
� �yr�<h�<@@J\�nw�$���[&�y��� ���A؆jI�L�a���0>y��|J :J�J�h}����M؜��jP%�����'���kv8�����ooN����JoT ��R �-�5`X+9�bDP���i���p��D��~\��ĦT#s�^�i�� x,|=@t��5�  �$LY�2����Ӟp0V[#�*bk��ć�&���d��ruD9��NM:Y9���Mw�	ޟ(�IT�S���) �c�X&�d��4���~�D1�S�OS��g+܄d:hr�H�a1�'N6Y�%�'/��	�`Ә�� �ϣ|��� CA�ʌ��N�^qOD���	�e���J Ll��yǠ�-wΊa��g$g�� ّ�ߴ5�jx��E�?���)��	�r�ؠ��.�����C���D�j-��]���%#�~ӓN

.�\��Y��s#b��	��M������� ��JՄJyk!�
%P_�0�§�ޟ��?E�Ժi�T}Q�B�/(�t�r�/3�~<�O���	h�P7�:(��e���*��<�v%,D� ��ߴ� L�ӵi�_����?9$���w�Qf�\ps�[��$�`�y�ġ��A�f���gl�}Є\\܂��O����@������^h�s���1ܮ�nZ�e���2�S'��5���b���C6�ȗ�6b>�X�#��$�B� 
� �NW
ii7��#���bӜ���:��i`0P���{{�ű�AO۾�K�'���9ғ4�n��K�*� �s\�AܱGy���Ęl�m�	�?��;j-� ��5@�H���M�b0a�6�'8�g��Z�	��'~��'l��l�u��ۦA[�(��D]~��e�7a�"�҅��)5ɖ\:7�h�E�5��3MF@S�'D�V���M>��ϘP��I�e��^$Dy�Nؔ|�<�G�7b�;�Η�"E�O(����?P|`a'�O\bSX�L�0h�'W�<�)��U�H�eAٟ�i�4O&<�gyR�'��I$2��cU7s�����NEB
�'L(�j�,�#dH���.P]�,��4�MC�i��'�FE`��O+�I+��(Z�"�0�~����)ՠ�h�#�g�ͅ��ş��bş�/GFI��솳zh�e�cg#et�@����su����b���*WJ�=.A��Ey� W��ōE���0�ޞ ��q�(�h�~�`�*
c��� ����V]0�M���O�mт�'(RAs!刘f���(	p"��G��6��O˓�?A/Ojc?�x%��8��I���F41$ɑ��3D�$�2�ݽvT*�۷�B���1�
���[u
��M-O��n������?���X� 6%ܩ'�Hi�������b��V����ҟ��ɝ
y��!Ʀ�ɂ���$8�:d Ywt��IF��1*��ٔ�?2�6h�Nݼ�(Op*։ŎCV]��������4d�Xp DA"r�0��'LÅ"�|�d�;vq��i-��I�����ئ�PK|��4�F��\p��c̥bQ��!�'��O>��'��tr�#Z�t�k��/Gbnl"�LA���{��6�I3X�
%�X>�\`�&ȓ([��?������'ڸ$� ��(   q  g  �  �%  (,  �2  �8  L?  �E   Ĵ���	����Zv)���P��@_zX�B�W4T���9Q ʍ;A0X��O����66�L�w��Tx��������/�`�	�'3 �H���,.���: "7!G	�C���B�bh�+;6:!�e��.�H��$<��mR� =5oN�� @��kڜaW�7U>��C��
�=~� Qr!�L�0�2&��!>˄�8#F/
􈥮� yf �
r��)V����"�P?ȩ��f_2xC"��ǧ�4��L,��=�(#o�DТE?gt>��O��d�Oʧn��9��*f7�ذG'.,��d��+4��t�! �����s��N矚�yF��F�':,�+�!�|9�� Ӳ(L����F�Q� P3-��:~�:�'���遭f� �%�(��b�*ZZ� �`ʍF�~��b�V�Ċ" ���/!
���d���+s帐螨�DԺ%�V;N�l�2ռi:����; 	���b7t}@���"��F�g�:%o����zݴ�?�'��-���@�$�2`%	�"I/@,��Ì&l�"��)�Oh�d�O����к���?�O�n�c��/;����%���e���s�㜯>�"8 Q�\8b�"hȤ+�&,Z}K@�X�'�"Ph�Q�U���!��*���Ղp�Ψ��	;r�����6y���$q�'���p�e�`�D�o����ѤI�;�H�S�iW�"=!�����h�F]>w�p�+����k�D��'�:�+��\�B���S/W>W����O��m�����'�1;�g�~����d��j�`�
��
�+ �E���˃�McD	-�?A���?�� ��r�<Q�v�K�;�d�-Ȋ4>��ׯ�2P`n�X��0!VF����	�s;�Fy���d� �D�:�t9��D�H^������9|���g>o".���_����Gyb	?�?�i�@b>���b�1a�V8�!㌟	e,'��>i��t1������S�Q�"Q�	F�������ja���߯jxd��Z�Ms�	�Z��ٴ�?�����)Lw���$�Oj���c��n~�qӀ^�`B�����BզM�'�� Zh�� '*T���I�a��,`L}�'S�2<S�B�2�)~t���x��A�*c�D3"A�/���*�+_#3-��>�z/��pq��`�K�,�:\&�ӟg�O��lZ�����?	1�^	E8P��$
��p8��,P�<I�E��:��A�O�e���xf�SJ�'`�#jQ�Q�x:5�A`kphYt�!H���'��K��/�L��'�r�'���`ݵ�ɨ�����si��{�@�Lo���h��|�&Ȓ�ʽ4����$P���閁� @(I<�&�U�4:~�x2�է&q&�R`��[���$�'feb�4 �|�Os@�9oDT�I�PŖu��*޼��U���, �g��I��MC"��V?�'g�!b��-���J�SFd̻�m�B�<�� �!TaS� �f�r]��	妹���4�V�Ī<� ��K�tQ�ML#eyZ%R�j��(�0�K�?	��?	�T��n�O���y>��G/X'6}��rW�� �t%�+r��ȓ�Ug����rL��}"�-S�OæN0Q�,�G$�
P�X�B"�
�� ��ß
� !C���=b(�ʃ�FLMM�S�^�S�Q��"E��O��� Ǉ(�|�&n�5h�zf�������,�E�Z�ԊhLN� ���8H��B2��W�*+â�`�����'h�6�OH�JL4�sQ?1��I�ÂR�5�6I�Q�tV����U����wß⟠�I����K�OY����aX&��L��$�20�P���p�>�(R�ߢy�4l�#�<#���<���EG�~uQ)��O�t$��K���v0@d���8ı��(��|�6AR�'X�o�Ƣ<��k�ğ���4W�1�
�+��tNV�k��%OZ��7]����;{(d��$G�a����a�ÐmeR��$�x~�E�e��(�!	#i(�Z�M\����R�)��Or�$�|���?��D%
i��AhiN��ޟʅ�շiҍ��@2-�@��fO� �0�{C���  �P�)�"Y�/˼7<a�T�@5.�"�dZ�G�ltz2e�i������<!T���D���O��sׇ�%�@��d��;\���P�'z^Y��at��«<%?��O}
��gϸN,( c2�Q�zAJ�і"O�U��K�8~x��G�C\>Pz�	��ȟ��°�PAۑ.�d����,���o��`���5�,C ٟ��	�|���uW�'�4���`�T�H�:�#D=:
�g�]>\,X�-�*&N0�Qe�3SS �':ŦHq2B+�O�vNp��%�֦=�2`�Ьʯ*1 ���B�2fgj92��9����U>	��NB�;8�'~�M8$N�|�:�[�S'Ns�,Q*O�)���'�<7 R�'���G���b��#*"�S��<|2!�d��v+rR�FU�r<\�C.��0�&�:��|Z����=<��8�/m���y&��� I[4E�.���D�O6��O(��;�?A����T���?�ë-G@���#BQ&&ժ�2U�}�M�)�~�m� x���I��1g���o�!��>)�o��(�0((t���_Ͳd��S	�yR�[�1AgK .DC L��y�k�Y�b��3I�-�����,��$�⦽%�0S��'�M+��?��O�)b�S4O�H��ė�KQ�1��4{7xh���?���"����혧�d�Z��{Ph�]�<YtI�hOeBA�3� 8\�����sn�P)�AWh�S�1����M_�O``����75<pI��L�78>��'����4O �F$#pL�=+n��
������Խ���<z^�	i�(u�n�dr�i��'��89$
m���R�oT�tT�7E��{��T�ɹ�M+�j���?y�y*��O�=Ä��^x*���A��z]���'϶�����"y�.`�K˙<&��*��;<\5������i�)�',��h$�lx�H�f����ɑ�'�{��I�X��Z�Ye0z��dD�O�^�z���!@Z�p(�(߿0�����zӸ�d�O����w���$�Ot��O����Ok�X�p�j1aN��y��M�ԡ�e��I�2�.��$[���)��ڃd�`R"�F�n��I�\cZ��dX+}�(f�R0����FF�E��IH����]�����%K% �aX��C<T͜���8D�d�A(+��I����l�s��c�ܵEz�O��'w�<��` 2�2q�f�U���u(�ϗ�i3�'{��'���t�a�Iܟ�ϧ|iܠ�I�Lr5�kL�je$�Q�Yy�rkd���9<�qӎ��v�9��$ۊm��؄�	�o����� g\�0��]pԴ� 0tְ���o/� 	���g< ��w�Y�[�:���S��S�= J��hj�L�'6�8���N�& lZ���IYb ���0*u@ٴB#��#�"A�q�W'�՟ �	�d�6���\�<�'�t *g���~� ��b�շaEpF{�7���z��I�ql��렭8%��M�E�ɘ\���d�_�OՀ�YӏJ�@��5�	b�	�'*P
!�+��$z�L�v\�`��-��-kX�Y0ƆNCz@]�V�\�:���o��"�i���'�1j�y�I�����Y;��8T��[���6J��M3B���?�y*��O���C���@lۻ_��2��'��Tx���/W`�I�� ĝL�~�*�ĕ({��e�I�\L��j�)�'I.�is��Nlt���؈}��j
�'J�=�b/[4�-����0������d�s�O��PVh��.�t`cf�!@b٠�v�z���O���W56P@��O����O4��;�?�1D��2f@�E}�!�1E��x�ȸoZП��Q®Kt���ނ�0<��ϑ�B�r��b�S��Sp��A�oJ"���i��'<|���O�d�4A�O�I���مˑ�gNT����"�6��O|1��A�O`}l���Y�t��]?a�'ٸ:�R��΃&�8p��_�'��xR�V5��$Գ�~����Y?.�"Dn���M���i5�'� $�O��ɣy��-���5.�~@a ����cwB�2-q�M�Iٟ�������^w���'��O������,7<m���4%�PY�d-̔ˣ矌�p=9�D#�*lX�投L~BE�K��&����6@O�&�����X�L�Ʃk2�2]l(�<�冂Οx	%��4&"��"��$*��t�M�M��x2�'��T?�r��X2��NR&�4O���H�!&�{4[B�[�B�V�I7�M�A�iH�	2�!��4�?����T�I $�-��'G����aQ#��M�ţ�5�?����?A�M��l<��sU�Ki�jS$$�9IVEڂ5v��"A�g��p pk
Biz�Ey�BZ�vH��$EU�J���FB�����Y�Q����� � U�~m�Em��O�@�Fy��Ԯ�?���E��dQB*�%�M���Y"#D!�W�R|Z���Ćt�L+�@|1a}��=?	��"z�R]3�&��s�ڝ��  H}b!M,N7��O|�Ĥ|*�����?a���><��U4�ݡ׫L=m/N�5�i�5r M�+��	UK2���a��~���h_����ݹi���$dV116r||��
*w5����%Q,x�>Q���m|�� ��S�&*�VOϟ���'�O���+?%?�II?a�CQ��6���bŖB
��ۃ��I�<�����b�HũG*�j�\u���E�'/�#"�Ƃ��\A��S�8���*fC�m�&�'�"J �r����' ��'�2�f�]�I�GI����	���.�X$�^�>���u��>�8mЀ��s.�y�`���.lt�1�����Z`��&<e�i��B(��a2n�3�`��Pk���	�?�d�����	\���:�ǈ�xc �%pI�����In����TbN�w�n���M�RO��1rL�"�y���a�0��(�T���/�MK��i>�INyBmO��=˒��z��A��UW�,B$I�.���'�r�'Ψ��P�	�|"�N_(����<�ԩׅO~OD��sV��py H�F/�����!aF����"��z��QQe�I����1��(�t9
%n�EVB,Ȃ�1���������� B9!��8qF�A����a��c��i���D=�����W7.���`�l>���&�2D���a�,���NE�i��>w�iY�Q�̳D�D:����O����a�LP�ՄA<U��T��YU��6�������O��D�p���hz�&�?m"v��1j��I�iF�D0&,��R�����yc2�	(([�qi��#â��GͶ\�Z|Χx+l�*�g�-DB�)��R�n�V1E{�Dފ�?�����O���ED�u&\��'�ۋo�\iI�O�$>�Ox��"��G���ف	�?Ϥ���'�`�'9Z���I��Tmd�;sY���'����Bs�����O��'{嶉���?i2�H�k�ƽ�* �d[�4�V�^&n�vL�.͎�!u���L�$a�e$@�N�Z�sbM�u�1����5���^Җ����ʤo��i@��O>�y��TX�f�Zd����V\H&�n�DI����,M�S��d@R��0?T,�JCˈ�]>r�J��?���������'��DI�v�Jx�'���OB�
D��N.!�3`YC;�����W��@��)�z�Lр&⃗2|m�e7D0�m�d���8 f�(CH����ߟ��I��u'�'�hLCfᄻ9�J�%2b�B�T/tF�p:�Ѫ7=� Ҡ�)k��'�O tC�C!6UzQ�&�ĺ�:۳�O?L���k�G>^��,�s�W$
��D�'9$d��/��a�l0���)O��c.O�����'�����I:ʬ�ㇹ4[<��I w_!�$<��<� �T�~�����!ء(@�v("��|�H>i��ט:nب1�,D,�T|*��P�YxjI#Ć��?)��?�5��O�h>���KJ�����@!1>�<Z7�
-'��� ��y�Ƽ���G8EWxl�468�<Y.�^1HĨ�5R6v�:B����]���@�.�r6���8�`��i[��Ey�Ŏ�?��M {��X���5gH���%}!�$�=r�ti��]<&rl�Sw���e\!�d�gIZ5 ��F<uc�1Q�d��u��6�M[O>y�'Y�lW��'��֟R�S�@�4H>v��D�p�����iv�೶�'��'�1$��%{��l�G1h�����I͑E(p��*ܹR��y�K$;gP@�ݼ�(O^q��,\�
=tLI��F?+5��f�Q'o�y�E���kЦ�#nG8;(  c�F�(Of��&�'X�"|ʃ�@�%>Jx&��T?��
�H�<���%Dڜ̡`�
�EV!qf��AX�P��O8t�Ū�uD��K��]�	��h��^� beQ9�M����?�/����	�O���+`�X����~��,�b�L7]=$Uo�PΈI�I��vw��e�
?Y�`)�,������|27'�)@��q����rPLF�N��?�����e��8Q�:\�6��.8S@��D$�ORӑnS�=���4̓k��&�'�>����ɧ��҉갨B�a>���J[黆�6D�(16,�4}<���Ԙ��s�)�\��?	����(\$ ��I���gƵ�MC��?��[;7�T����?A���?������Ƙ!@�/Q���g�H�,��}+�FD	9m�-��6NJT���"u��Q�'����(7A*}J���:m"hڃ��i�V3��9��/^�1�O=�@�t�R���8�� `Қ-���<q���h�����?1�O��=��ʘ���PB�kƝ'kA�	�'q�\�����t��JR�\>0��!��44쑞��㟀�'�pٱAٔl���n%��	=*��@�'"�'�b��a��˟��'��d�D�-hd��.���)�	��nr�K�Ĝ�q�2��L�*�ȃ�*ʓbJT*G�X�B[�b�*C��J��h�-p�\��ʲ}�r䓒,�5����!'ʓrX�ɀ}Ԏ�#��ڋR�i�ȃ%u�;�4�?A�R�s�4mh�&�3|�ܛgҧ08��e�'Q���g��X�H	X���BX���,�>I��i2T�������M����?��OBrazbKK�+�vТ��ViZ0Q�4^��y)���?Q��.\`Cv�ل>��p�4y����˦��aS |vX=H���mQt�2�S�+�Q�X�qO�K����َ_Q�M{"����� �b�5�Gg\��EK��5zo�	PuI�J��5{o.�D�Φ�QN|�& D�)�� 1�gN�<��]a�e�sΛ��'��'��#nB|~�p��h�6[�J�L-�On�=ͧ��f�|��� *��(�@��_�Z� A�%�Xw}�Ըh���k�=9�:OB��HOB�k���\B�Y����zP"O�Q���
:�LHW�1{p�"Oȝ0��G��T�3eF�l��ZC"O=2ą�6S/>41��
�!,A�"OdXc����'θ��J�tb����"O�1�tn�iS���D�~4BX0A"Op��N<֢�R�/ۆ��[!"O�U��(\��y&�H0�n���"OR��T�Y�$,|��Q�N�Y �F"O� 	+o�6�Ȃf� er�x�"O�p�+�Ǵ��E��g�@��"O��Æ��S����)#g�G"O��t�O!-��)EDV�TP�"O�D�v��n�l�3�.K4���f"O�]+�^	^{x%��H�^�|��v"OL� cN�G	�@1�����"O�c���"�������v�"u
�"O:d�2ȏ�_>r<(�b�=6�4"O���� �̅AL��mz�j"On�+0n�$o�TL�磓>�"OLa�b�Z�=������Z�}��"O���!�W.y�Μ����L��8k�"O�Y2u��5iaR�fU.9<4�ʗ"O.@���I9|t�cc��``=bR"O �@4���IC�
�/���"O�Ye��'����H��tJ��yBG�PТp�2aԽL��0d-�)�y�/։i8���bNVG4�!�����yJ12�~�7�)B�``�B��yR��>1��]hA/��*�>0(����y�Bڊit����L�-іK�F��y�i� ��8S�l��5�T�d<�y9a�x�9U�Z52Cd ����y2�*�@�D�͞0"*�@7l�s�<��j�;*q*���_�n��hucQ�<%*��M�d��g�!O���m�<qD#�G\��cFCv�����]�<��
�%�H)�����D�\(����Z�<)W��+R���R��ر>�5�D�GT�<I%���JI�m �MҢ�P�s�o�<9Rd����)�g�N�d@�&��a�<I�	)�X�H���@0*�c��a�<�w�"�R�H �_�FT��@� &T�L	!S�J�<M��&ݦ7��5���3D��"O�b��D9!�U�Z<�Lzt�=D��jvK��W_^q[g��5c���9D��p��ϝ$��B �ҽ~ 0���'D�� ��J�%2��������8*O��¤�E�2 �U�ȇd���)s"O��re�8YF�J!�"��� �"O�%s�D��*�v����>I�x���"O~y��� P�2�S`�$���:Q"O��;��S�~ll%�	o�aJ�"Ol����G�i�jpцF8=���Q"Ot�B�ĸv�Hm�� ey6"OP�1��0����Ȓ�8nN�Q�"Oʡ�$�Ȃ.H�F/C�>�r�Y"O����e̸}�@9r�,^�f,��'"O^:�Ƿ}�,�vl��	����G*O``TA^�69JE�⒎�B!�	�'R,TI��&�"}H��**�8��'�y�%9�1"F��&&V��{�'M��s�+��`�|�p�Q<����'n�(�6�N[n�Ђ�/O��t��'$�y3F)� 2���Q&�D[�$��'���� ��g���`�,ɢl�9�'.��RɮZ6�#�Lk�����'��ݛ���A?D9�J¥c3�
	�'��B��Y��`��
ĮLlI �'rVjbƑ5j�}�bL�t� 	�'���37cP�k�:�H�96&0��'� u�A*ʨE�L�"�0�~@��'x��͠ �hl �KA!'��I)��� �hJV�A) ���1	ޛte��"O�\+�%�h�����������Zr"O<�"� ��)O���7$"�p�3�"OjI��������Fj!y�t�B�"O���־0u�#$h*�z�0�"OR�������X$��E�F)9�"O& ���u@v�w�ƺp�8!��"O�,ر��a �䁥�.5tM��"Oj0[��@�n%�E�c��s@��"Of���A�Cw�ԡN;,r���"O�� Ǜ?t}ᴂ��l�8��"O�}	w"	�lt��w���oNn�H�"O�
%���EJx�l�M����"OT}R3N�&^��,�ʔ3"Oh��:� -+ (X{V ��"O�0�6��lYO;Y>e��"O���@JM; �\H�7�Тs����"O����O�O_�-RaLf��"O(A��P~+h1��pZ���"ON�	3˘ cL��"Ď�M�E�"O��;��۴��h��7BR�p"O Q
�n]�2�D��)�"b���"O�y��ź:*���
F�3s��J"O���G[���7j#Cq�\�"O�u���>�� �ר!���"O���ʑsn�)0R�ڷQ� @�"O�x@A��m�j�ʓm�##�� "O�����Ř{j���U�C�DD��"O��
@�#���HP\���"O�kb�����jAk�����"O~ix�	� ��:CG�{lQ�W"O�X�' Qv4S�\�F��TK6"O ��!�"M��*�h̰B���"O,�wI@�5n ��w�ˊ!�8=�E"OL�3�A)��@�Q�9�֕0"O6��s��;e~�8P��}KhŃ�"O�A���ֲ�k���t�L���"Oj=��E#K<$3b	B�y�"O���a�_�����c�D7[��r�"O`I��D�yP�A]F���@"O�}ۆ"��W0t��˒�x��a"O����'���b	��`g*0MS�"O
X� d��^�8`�%K �`"Ol�V�:6i�@C&Б s<��"O�ՙ��^4x��z��?&Sd��"ObQ�5�ţ�&eY���jP�l9�"O��ʖl�9*��;��)3��9�w"OެӤl�%.g$�iC��`���"OHy{�S�#@a,T���gB	��y��	*�q��h�:�C�⥆�_Q!0��$�T}���y ���X��CRb PZ<ԣ���=j�8�ȓ^����p!�>��\����T�<��M�huH
%'�&�
�l�@�����)8d�g��� �2Bޗr
6��ȓ9%�w�8�漪�ܕ&7�`��!f�0���%�V��t,�.�)����X���S���R�#N�ueb���b�҈�"�[��N���L�ȓp�]��@�6G!�Yj��Y��JU�ȓ{��d���ϣ]N�E.�%1�&̆ȓg��pa�ʅ����?	�Z$��B	L��OX�:@ A��=��t�ȓs,&���ᚗ[��b���.؆�S�? �0����H�:G*�$J���x"OQa�-�{è���N3��@��"O�`Zv���NBIĎ��w�ZX��"O�-�)��J�x��Z��t�@"O�uc�U�
��T*#G�U�����"O!R����(�b�h�C˄��*O��r0�"A��E�����yZ�'��	#d��]���z6̅2o�1Z�'�
P[6b*z`H�qF<F,�	�'j�;�n�k�l��bX)��8�'� �#e\(5��x��KG�^Y��'�Vy�rG�-�.q����T6y�
�'>ʈy�+L�
U��H��X!:1y��'��*�
R'\%N������1�(� �'��	���R�=�6�z�^�\�<�K�'cP�k�� ��"�>Tq4`��'o�L�D´4&ةc̎!Sʤ�	�'N���vo-U�X��R%�(D
�0��'��ёR`
�Ѐ�����~;4�2�'�d�B	L�6�s��L�w�2P�
�'$\�C���W��0K���p:�-"
�'�0��FϚ�o�d�*Go�8c�fy�'G��3�Ư>S8I9��ٻ�((�'�F<Y�U/�n8!�%شk4��'�,��HYe�Xx��Ϻ��)�
�'x��DD	B@�
m��9
�'ܺd ���k.� GB=<��� �'|�yJGIG�f�,!Pi'-�Rԩ�'���	1⍥9e��H�/X>sښ���]�T)��C2`��xv��pz��ȓ|�p����.���·$8���'��q����)U�F��u�Y�d�ȓIg*�H���P�|�����#����}v�t��l��Y�<�G0I��ȓP�\�c�	$I����w��
2b���I���0�ӣ-T�y`l��7����|���L�6�$T;/���JԄȓyǠ�(𮑆.��Qd�,�bP��&��a�,�z�~�R���.}�܅ȓ@�UBUe�J玩���b	��ȓ� )P�QL�X"0ěy4��ȓk�v0�"囧G
�f�\�Rۖp�ȓJҮLKT� �Qg��e&�-�$����Q'�<5aB�N	�T�Fd�ȓ`���AN�6
���8���ȓ��g�A*Q��Ue��r���<c�u��@'���c����:���D]i��2C�e�� ��W)޹aGO�b�(L���L;[�F�<1�h2R��4���B
Թ3�T�<Gj�.�n��`�L\-QK�d�<�ń�_(�LI�,�9�Z�yC(�`�<�`�� x�Hz�'ܵIW�w�<���C��9�0Ӽ]�X�4�Xk�<W,O)a��-A��Z5c��{dEm�<�EJ@IJ�� ��0�����q�<�tD��9�<[�B ؜�����I�<I�7: ���FثG�nA��b�l�<1����EN���
X,�q�H�]}rN�,h0�`퇛e�l���@��HO�����F�
�PC�-?1���u"O���c'��A�� ���]!���u"Op`�TA܅Ԓ�≇E�4kw"O��傎�,��\K��_�\br�"O6ԛ3�M0�XLPU �'[��"O� �%��GC�q|�,�[f����$"O��'�V�]�N�����`q�"O�)pu�� w+ԁ G�4�ΤiV"O�|q�!��O��ď�-!�بzT"O� 4�U�d$"�ئi��Z'�p��"O&@�O�?9���7��@l���"Oް�A���
����F�J��G"O�*t-I'���-��s:	8T"O*TK��ڗ��x挂�3r�@��"O$()g��>|�H�S���.�� �"O�1�EV
�L̉� %o䉒�"O���iA�%U��1J��;[|��5"O*�9�ȗj#��iZ8�3"O �q�b]
u]���1�K�ND4ir"O��r4��,p���I) "Ob�2ӏ�f�f�A�b�/d��B"O6�Q�)!Q����7L����"O���bc.8$���#�/O�3�"O$��bU��|:�
�JPX!d"O�:D�W�uS|Y�6˥TQF�w"O� �̆	1��p#�C�\9nr`"O����הu���ɑ�p4.�+�"O���b�ɔ&t���nG!31��"�"O���N�/�r�[G��<;�"5�"O����O�^�j�ZC�8c�`D�'"O�0FM5L�� �u�� jn!��"Ot��ӄ�|�0�����+1 ��"Ob�31�׉+a���G㓭"~Ł�"O
��0�:}|�+'C���]�G"O���
]6o���Hp��DP��s'"Oj��̍4�T|H3�I6�Py"O��a��贪t �(5=
!"Ox`��S�+0���[<j�	�"O��5I�;��2`	�(p�V"Ob��,�(a���&��a����r"O�)��؊@_� �2�׾=m|��"OX�GW��@�	[::��ݡ�"Oh�R�oކMwR��g�0b"Oآ5C͗#�Hb4��'�ƐZ5"O�aI�Ɋ�ZE~�A�+ɾe�B�J"O��QM�%r��ѡ�*˾%��A@4"O6P�f"O1$����F8�R��B"O܍sCĞ�`�iC��9l%�"O�4��4U��I����P��k"O.ԑ���&�}
�Ky��H@�"O��SD  1?�M&�ߠ���"OvE)"+*Z���Pf��j�&k�"OP���럻
fl�hΈ�a�t][W"O����\�UJ��&�$w�dt�v"OvE�` ]��dQ���)��]I�"O�1�� ^�y�E�˧���)3"O���jL<���dʭd���S""O�5c�̘�$6�caQ�8��ʁ"O|�F۰ mj0@u�ƴP�Ҁ�7"O,�R�ȟ�hR�[2Y�6�)�"Of��¡J�;ȀU���	�5G�r�"O�¶a=!>����B�v'�"O��� ��a��dPP�ȰR��"Oڌ�@�{C8�)У�+�Z8p�"O�8gB�.x$�sCS�,g�m{�"O�9*��΋>@ꖢF�%���yR)L,x���3ԣʺ�J�BŘ2�y2i\�V��A�'�ܳ~�P�
�JD0�yr��4���1n&p�:!� �.�y
� ��pCe�1wV���D�L$s��l��"O��y�ʫz���b��w���J"O$E��8 J R)�pwj�Ie"O�h ��"DVe�Eh�.Z4�S�"Od�(a��8��w!]
T2���"O�D@�W�t01 @F9}1��9"O���!'I!�iyR@W�$v���"Oܥ:W�)n.u�>���2�"O�` ���R�<�
�'�%���2"O�tR�"�?|A� +D:޺���"O>��҅Ϫ1�
�R�
i�Ĩb�"O�XU�іy�&�o�>$S�"O��v�;5����O�t��"O`x+Fa�e��h$��({�qU"O�B�]�-�ax�烁wn�tkC"O����d�'4NPP���X�Ck~Q�5"Oy�C	
b�L1FN@6;� g"O����iq� �H�U3�-)�"O"8"��ҡX�>,�B�8���f"O�a�gŘ
INJ훶и�f"O�Mxp��U���iᬃ18FE26"Ol�!&�KVD�C��pQ�"O���"Ǟ2MȂA�g��=����"OH�* ��W`�8!L�Jj�y��"O�q�G-2&`dQÏ��rKPQ��"O�%P���&)���blYcޞyC!"OĈ7N�	^W�`�4��Z�F�C3"O.��)E�d~�	� lɪ�C`"Ot�YǢ^6u��s�)��\�L��2"O2Y
��	�T�n<kBc�N9�F"O�љwiJg2䡹g쨥��"O�}�r�<�(@�S_.�&15"O|�� �m*�����Ĵbɬ P�"O��zt7i��i2�gV��9�"O��W.F�>Kf=� ���H֥��y�O�}�P A�ĥYQde�r(�$�y���1e��T� d1֐�V�W�y��5��@c�l؟[f���v ���y⤌���A����"$<L�U��yB̋�_�e�m?�X���=ٍy��P��v�pe�:_\ZS��y�)B�W� ��"�S��)��>��'e��EyJ|B�@F2n����^(7o�<9�a�T�<YgK^>Px��� )J(9�8Yd���(OF�F��O�M��OθU<��O��h|�G"O@��"lҰ_�(	�ăA��w!����t�څ#��ֹK�e�a_1]����	�M֒O����^/T��І��� �d�u"O�x�� �B>�@9�K
H��!�ċ8M[�n�\�O��5+7��C�ܑ���J����' |h�,��GN�+p��J�Y��ȉ}�Zc�"~�F��E��E�]�4�s�CT$M� ���&�	�N&Y���2ݢ)_E�'�dek�|}�8���RL}�o�oz2Y���}?�0�O2��`m��Y��1���)1�dp�e"OPPǮkJE���4[�2lV��<�S���rGFY $S�L�R�R]�!�	u*j����Jd�Cf�7!��ĴsȈA��bͅ�R,���J�7P!�D��R�F��SiJ�&�T|!s"I&:5!�dY��2Qd¶d��@&+�NB䉰o	�s@�Ew���DDN�&B�	9_ Se�Y'�����o�B��m�45�QF��<�~�iaQ�3_�C�)� ��B%��_ۮ��S�^�io���t"O0}RE��d���c�`�|j��r�"O������%_�Ԓq/��rW�t�t"O<$;�M3Ը�!��i����"OR!�(W� ��-L� ��8��"OB��r�˰'����GU�UI��C"O䭢RB�!�d�[$f�%E�*1�f"O�ueeθ=B  ���Z�^�s�"O�����n�B9;��=�,���"O�-!�C�3G�<(����JĶ��"OLpCRW�xةC/E<?���B"O~%��^�Hr\�c�%<�@�!"O�����9& �!�/G���I�"ODP�d�PA�,�3��A�V���"O�$
 ����u^�R�T"O�H��Xk8&q�ciĖFT��� "Oj4�7K$U�r%���֪	j���"O��@��'V?��)G��keΌ�r"O�-J�&ΙWQ��r�Μq8ĉ �"O.P�T0^��CgE�|����"O��ȡ0x.ֵI��+{�u�!"O���+ |;셃AY+Ps �8�"OVdh��^=~���MĒu�ti@"O�]��-�"����ǌ,g���kt"O�5e��=�H�k3l�:/� �:"O4�VMy�!P�̶G-�����^E�<�/��8�Pc����wƙ~�<�t�$jg��`�V
3s&	���v�<I�l�O��q��茛7�`�( ��I�<� ��/msY�M̓Jv�\�D�IF�<���#c�&TzdaÓB¤P(��B�<I���+Ij&m+�E�S��]��VA�<!5�V���H���^�Ȥ8 ��@�<!@-�%x�h5+P*V�qV��(��~�<��e��`a𘃂��#]�P�1��|�<Q�Ĕ��&d���ؘ!��y�<!���G5:�	4Ď D�r�r�Ku�<����Lz�P��N8zV�@��JWp�<�����TQ个�IJ�{�4B�F�n�<٢KȪb�2���NǴz\�@�o�<	���>�@-�PD�g��L{��g�<����Wj�0 �.7�Z�+� i�<1� �k�ً���/� ��'�b�<QQ��7���RF$J�Mȼ�%�a�<qrN�pl���-)�����h�Y�<��V�n� � ��V�`܃��o�<�&F��H}^�$�S&�.0��]A�<	���8����� 8�`~�<��ݤ��6��	,G��Sth�d�<�f��>$I�a��rkB�"��_�<��<{��i���ЬUb֑�bG^�<��	A�(fJ�����'=@�#��C�<�p���U��)��nѦp`��m�}�<�P�
"Ȁ�#�,F�n��0l�y�<��"��q�h� ��:6��3֬�J�<I��Z庵�T�I!�s���G�<� Ά0��	�-����z�a}�<�f�>8�~�KaDӞ����B�b�<��+@>)�H*0&�e8���H�<Y�.Ć?7V�K�S�f��׭�m�<�E�Z�'<��CC�>��cU��d�<�eIW�U��i6�˿�d�ң�^�<�5ՙp~F�h��\?N{(Mg@�X�<!�   �l����i���⑄>D���#۝	�X���.Q�z�Ba1D��ЋѺ'�f`c$K^�Q��jUh!D���WN-jŶ��g\wf�pB�C>D��aB��es.�� �� E��\j��7D�lڤJߦD�-��C�M��h�)D� ���M%��YZF&C�B2İ�co*D��j��E2H<\�KR�E����q�J6D�|�u��<u�����6'�r���1D��  ��LM�q� q��u6���"O|�q-�"#�YBՏ�vGLdB�"O:B��!F�ҵ�q���x�Q��"O��z�,�$Z6��So���L "O�(2p%�=�v��FIߴQ��)�7"O
����  ��]+V�.	��jEJ�<��$��zd��螧~J��aT-�l�<)3����ѳ��V�(�9��@k�<�U�߅��=�g)��Ulr��Q�<��N����i2t)�8 �Ѐ1V�<	#�ޝ8����F�}���D�G}�'�F�*S���_�&�S���K�s�'T�%e�+,��9 �뎌@���Z�'�:�a��������%�h)Q�'g�M"�B*L�k��	��qk	�'$���-�=e���+bm����'�N8bnE(~z�T�W6(Ǥ���'�H�P��qb(I��	�&U�*�'Hڨ�ӳ +0��B/ݞ#bN$k�':J���Zz�-�L��$���''>0�C+V���h*��M�����'����	Ò�^���`�.8����'�^�I#��)x|B�dE�{$�s�'��A!���	tRj�q��0gJ59�'[�0�fۍ
���*]6_���b
�'���¶N�9Z$����C(\���	�'��)��Д>BL]���նC6�1J	�'�d4k�oR;_C��Y����'�p���'�X}��- ��J>o>� �.�y���x��#�`���$(Fn���yri[�BS��o�)�% ވ�y"]9
�qF_&��VK��y�ɓ�g�A�!�+0������y��A
���)���'�T�� �y�ɥv�8(���Mh�Ă��$�y2@��[��AF�E@�A����yBj]��&0�6!��:��I �̖��y"�e9K�h�$<�T�&	ف�4C�	�¨�+j�^đ��b�l���E&D�����ߴry2 @�Ø"P�b�ۢ�%D�ܹq���b����*p�8��&D�(�r.�bה
#f��	(D���#��&�����m�B�c8D��3F�14q`�1B.H<JV �kF�7D��Bϖ}�<�y��D:}c��B6D�(��L�)pB!���^#r��m���?D���iM9W��5f��>O�I��<D�T���B�#�� ��.3�	�Ī7D�� ���!d��kfA�
�CN���"O<k�dS��4��o�1i>��"OP��A
/6�����%8]05'"O����݅��i�p�l�:�k�"OЀ���U�b�00�߀@�x�{"Oq{��� n���b�
`�p]�"O���Ҹ!܈���"^�B���S"O����-�bA*�O��Dj��@"Ov����ɵ��I��2tS���f"O���vi�0��E�B��(-PX�"OH}�V��??#����W9j8��"O
�Ʉ�%�r�r�nҟ?�A��"O� ��Q7z�����F�0����"O��!k��u�.�ƃ�#C�b"O�,���=Pl�4�+:u��"O�PaF?3nh��v ^!=�N� "O\� ��0T��� �Aөp�حҶ"O�,[�K�,[!�>"����V"Ox=��ƞ�oĺ�򡝗h����"O�	I�M�,��� ��,.x�U�"O6d�P����� �86���`"O��Y���	�2`�B���!�l��q"O6����V����1��A) -q�"O�Ȑ ,����]3�o[����0"O(�Ks�O�tH|(��.��AX�"OfD��ؒ0'O�? $<��"O��ig�Y,Uo�����q��"O��������YR
4���b"O^�
W��������K��	(V"O-X�D�+U��yWKɧ_�ؤ�"OH���@Y=P8��g�XsJE�f"O�`��C�[�-������0"Od4�G����c��=UON��"O���/He���C��M��h"O��y��;�l�"����9Ժ��U"O��P���J���䞰O�f�K�"OΈ��e�}�1q�dV	Kt
��!"OD`�FZw�Ɛ2�"�/	SD�ӑ"O L� !��H���#'a�5G�Q2�"O62&͂�j-q���Z"��P "O�`Cb�Z�sL��Ac�';:�q0"O�D�F��'X(�j� �""����"On�*�O@��J]��R�tj��d"O�L�+|-�"`@˳_pZ�"O���jL8�Du �Ηhaji�g"O��ȁS�lP��ζ4Y��"OF@��W�1�E0n�iV"O贫S��/�6<x�#��bS�ّ`"O8��Ȭ=qh����	4J�!ɑ"Ot]���3o�"�s�^�*1�P9Q"O�p�R���?�����%Q�B�"O�蒈=l�}ze��9X:,�*"O&	J4h�+��p��Y�D�1) "Ony) "�+\�N����.FPQ�"O"9����U:M[�� �<��"Oн ť�:PU`�bͩ(���y�"O��R�d����]Z#Ӕ$˜�{�"O\|�I8Ԯ�����D��d��"O��8e������+�G���$I�"O�-��	�t�l�t�W�q���I6"OD�&	�<l��PD�B9�Y�'"O>ະ%ױ �L����ݳT0�hF"OU����:�ڵ�Ra�~:�m��"O
�!�	�N�8��!
��3�"O� z��Ыn�|�ׇ�h�0"O���#�"Q�"���/R�����"ORUiЌP�j) ق��p���r�"O��A��<����+�<��"O�y3�Z{ ��*�Iw���b"O��0�(�I~h�5��4~j5:�"O�X�M��N�	��� }���"O����hG,$m��I1O�i|b̑@"O��K#�]�]�z��-�*`��p��"O XsO>- �� � �|����#"O�h��fU�zd���³���Z�"O�U���Џ]���X�+I�dT)C"Oj��5�9M�`�)=@c�P;"O����̂G��,�(O�CfP""O�x�N�;�HHɂ)M�q3�m�"O5
c�Y36�L%��L�P# ���"O�H�5�3Y]�ݛ$Ȏ,^
����"O���P�1��!���?sb��$"O���o��;�H�C���<]�H�(S"O,���B&N�8�ň�:��L��"O|��W#���sE�ܧB�2Th�"Oh����Nd�[���%�ZXK�'fjqRC)�9X%���C�,]>$X��'->�C����'����韦}��p�'h���
�1��	�qc	!	N���'��0 �@iU�T���7e����'r��pc�$GofI������(�'j�4����AQ� h�����'Rp|�թ݂8y�Y!��	� �{�'[�%GM�3!�R��!��j����
�'�����ٟ��-�U*Z�*
�'Y�J��k�E�eK"ep�	
�'72��]�g���% Z���C	�')�X۴�	�*�����rςT�'n��@���V��D�� 8Z�'���e<5wVP�d�_/]�k�'x�<	��68��	�$j�-^�V�	�'ad`��Ȩs��fP�%Ɯ[�'좄@	�{PĊ��١#�� a�'�8P�d�C>�hdC� kR���'f<5)Q)�]c����L����)�'�bT(�ϗ!u Bm�d���=���'��`�,1Y���Ѻ<�0I��'c�l1�m՟K$����P��f;�'2�}�F�>���&��`<`�'Šq[.��*���b��~��<��'n�]���$th���E,p�|�k	�'����gƣn������<n�J�:	�'��A�a)�!wmZ���G�0gR�Q	�'����D�� Δ���HN�'��|q�'&�6��D�LK��[?���[1"O�m遦9�)�H��o�`m��"O�)�B�)z���+%���� "OV����U!�>�P�iY J����"O* �7~��Gn����j�"O��� �9����"W����"O\�# �L��`��)�yE"O�)2d.�%�E��(3v�R"OvL0��Y"C� ��W Y��l�V"O�д%�0�0�����F�lAP"O.1����ƄI���X3�"On�0���Jy����'O�g��b�"O،��ƌ�#�լ=�\ 2�"Oԡ+2��'ep}�C�0<���j�"O� N���1O:��k�D_�p5"O�8�6l��x0�A�$ �ZA>q9�"Oڹ��G�g��p�U�_�%�Xy"O�$B�L�?e.��#�!�  �\�$"O��)3�ss*L� �J�62�"O^4� b:���6B�"s���
"O��@�U�O�LT3r��8v� ��"OnP�mَ��PBc$�¨��"ON���֩V9�X��� ,~D٩b"OF����ίw�0�����p|�HF"O~A�b�!�ܑy�A��~��a"OؼpS�ݟy�lX{U >|v9��"OTQ�sK�m@2�zR�V�P]HAkV"O.�D��6t��N�	P�lȱ"O�yHpJ�xs�l�d�ֈ9�"O.{�jͻ(�bE#'�4vB�"O�Ea��@7cp���T&�nU�2�"O�9�����'Vd�`үԈ 7:�"O��.�)�L�[CiU�$v\)F"O�x��L"[;~����]�	FYR&"O��Cq�������Y��LY"O�0�!�Satz��	�S��""O%	'-��Nz��⣅��*��&"OF=H��I��}閤���U�"O�0�7+����ꃭ�4�`D�u"Oи��H�&�8s#g�,X�K�"Oj 
!��x��s4f�T�,9��"O�#gZ�_�hYg��m�4\;q"O<�"�\)o�X@�e��=%�|c"O�m����0T�qۥ����`(r�"O�5k��ß`����|�4���"OR����E7I�}��ɰR�Փ�"O�J1`�_z�ٛ�J
)-ef�f"O���� ����+��)��E��"O��@#�[+,��j��Nn����"O2���,�]F`�"'��6:Y�E"O���a��*:�=���Ȯ3��l�"O��#a��F�4�Se[$_��Ȃ0"ODL˥BҜ¸y@��?Qfix"O*�ithP�MM yi�"�G*0:2"O��K@M�sl�R`Ź!�n�I�"Op�{S���$^�[��J-,��S�"O�p�b膡$�l�*��
+!���"O,X�u-�=a�`zt-�.��l9C"O�x�G���pxR��0��q#�"O"`�wP0 0�[`�E�Z� "O���ƃ5VW��	�Ԏ0����T"O�����`�"���B{$^}R6"OT��Ҧ�=3���)�H� ��"OV%�'C��i���S�.q��"OΠk�`ל\P�{���
���Q"O��B�ȟ/W�Є��� ��<2�"O��2nY9���H࣎;.f����"O�pd#��/1�<��֮/(��R"O��Zu�N�J�Y���A���ʣ"Ol�:���}�h��,�b>�j�"O��J�*n{H�c�LN�Р�"O<aAT*Go���%���!��U"OxY�w�k
�\+q �-'}�#"O2�D��)\Ǫ���N�]Jٰ�"Oz���*E0up�b��F�3�<�"OJ�ye.��3~�"�����<�U"OIyG΃n��أ0�\'l;nD
�"O21��l�V�����v\(�"O� ��²���9��T �	6��@"Oz9��d �e��Di��H�U*tE0"O6-��"׸7������]�@�bř�"ON�Ӷ�E������F~T¡"O*8Z���`��5�!� {h�8 "O�۳�{��I�#KF�]q�
�"OJ b�W:h�=���;��u�g"O�U@cG#AT򼪢��&/��@�"OraDSθ�ä��� �p"OP�� W�L�D��7|�ԡ3 "O5�&��Ol�ѱeB�Z���"O~����G1� M[��R�:\��"OXj���/�D���$	x�8�
%"O��iW�D�(��v�C� K��P"O�<:����z�p�іC�P)����"Oz%��� �k$���p"6��"Ox��G��%'4xhJ�l��%
�5�E"O(Q��g��N�I"��Ş�Q��"O|ٚb�D	�p@�a_��L�#"O�M8�'ޗU� R��J�X~l\B�"O��(��7o�"��'J�ojB�"O����b n	���yg��J�"O��:$�PA�썊T��-(]��H@"Ox1�w�V<oK`]��EKL�}�V"O��aY�@3�ԉ��� -�I3�"O�Y�c�ǨP��Ţ�{�=��"O����)[�WѦ}+��̓G�U��"O�a� H�W����ǆ������"O ��`I���er&kY�\I���"Ov�k�n�d���`ιqD��W"Odm����0EbI@o�'=�q��"O4u�b[ �Q�W�<@��"O>��f\�&_�uIG7]%�D9�"OJ�u���hZ�S&�>hl9�"O�����дv|T���ބs�E:4"O�#@S�V6��U䚪\�!��"O^(�e��, $�lڇ"]�Elّc"O�)q���ˆ�㖡I/��<�#"O�ʖ��1w��E���n���C"O8����'��*U&^��L�f"O�X�e��w~�{��x~�q"O�������0iQE*͐|��X�"O��	�N�'��9�G�El�li4"O���D�R�Pq�� WRZ��4"O�<[&Q0 �X���:���a"O0y���5mz���eZ�9C8��"O�$�F��-�Zdj����o2��"O�pKP+x��Y���:K�=�"O䠀�K'9�x�3��'-<�1�"O~ 3�j�-iPؐ��גV&b�H�"Oґ��h5So�M Cm��` "O�p'I=	��hS�G 1�ڰ��"OL�S��0�N�;�DZ�K��dR"O&A
s�/n(q��C���A�"O�PRgj�6%��ش�]-Q�<}p�"O�J�c^5~�ha;� @9(�����"O��dJ�=-"���N�c��[e"O�QZ��� z�*s�Ĝd�9j""O��C�L��+�xPBlCLe� �"O�-"4�ڋ?��]���ܒSb2]��"O�jE��m8i���kM��0"O�A��Ǘd�J�e���hAK&"Od��D�B��>aQ։ƨ)À�e"O�T)�ݗVJh��*$&�d�u"O� t(���/s�}���	@F]��"Of�;�D�sl�ᚅ盔;X����"O�!u���y�\�+s�u<���"O��at��85 ���qM��!�"Opx3���GN���g%\�_�qb"OT��H7ڬP�'�M�K��"O�U#j� �"ɩ�lY2l8�!�R"ON�	 i�!k�v�yҋ�.l/��"O0v�̕9�v�j��9�PJ"O��I� �5Vs�(��J��nI8`"O��A��$d��!�**D@H�"O��
sg��!�H������[�"O�c��9��
�O\�X��"Oxx����(��1�ۂ=��"O��0#��B�8Ŭ�4^�dL��"O(L� ���8���@���07�|Ź"O|`I��۪GLX	��AI���q"O6lQ�))PM��l��AA�l��"O�и��P5{�������K!f���"O���!� �g����ۚy��y��"O`T��`ˆ��pcg��mк"O��:�!S��zM�s��ΰhKR"OL�)Ц�"�8����M���;�"O������ 4�\��� .���ä"O�d{���\N�qU��Txn�� "OT�"�JN��(x`��	�2��"O����ϞiO��a)YXP��&"O�DЃݞξ��Ei�Yf"Oles̈�z
"�Zp�MV�E"O��C����Kgɒ�<��"O�u)�\;����!M�8su"OT%�@�ߌx"�u�eO�WE�ų�"OX��@�8��l�L�1���"O�8��*�E�e@�)2��"O�I��I�C������ਈ:@"Oʰ!!��(/x��J7-��0�"O�=祔����
�#$�[�"O��eJ<t�p�*2G�0N�@!r"O�����\��CF�<[k �h�"O�����_Y��Щ�d>(j~8��"O� �o�xV1a��+z�}A�"Oԑ:e㈅Y�XE�P��zm��*d"Om����(â%�)Q����T"O��P7UǊ0�V'�G����"OXт��Hv<e!0A�?BY��q"O�u@�)�3� i[�F_(vL���"Oq�mݚG	���u�(1����"O�m���KsK��:�B�"{��X�"OlA���t���a�'����"O��B��XU(ယ���K�"O��A����(�����a�4-h�d"O�(�/�7��YH��Uq�"O`�v���!.HiR���T�R���"O����̹GX���j�#+�nx��"O��
��p6��z�ǂ�! ��ZC"O�`"��X�+���Q5���s��	�"ORE{G�=�pbB�'�p�p"O~��i�7Yβ�8mW-.�ƕi�"OFģW�1�ñˈ/OV|5"O8��r��c-4|�"�	Tn-ڤ"O��
s��}�r��	 `pl�U"O,$c�ܵ'�H ğ�EF���"O��f�Џ[f�sfB�iP�P"O\H�'��j	��JNX�Tb$"O� �Q���^��e@�h��L���e"O��p$�C�#G��y8����"O�x�#Ӈ7X����I@U1��"O(f-��<��!��l�Lr5x2"O����6�^�9W���g=|�!�"OT��ꀂ*t#�K	�8�<���"O�y��pa
�0rē�N�
MS�"O��i-?	�X���(@2�!��"O���5������u�� ����"Or�a�畜�:<�֊�6��x��"OTd*B�Z >���hO?"��r "Ot��RA�8�p������L�v"O�A3ck�*x0T�� ��`�
��"O�Q(��'
��u:��"S�-��"O�����@�H��f#Ə|:�]z�"OT�(BB�a�r9xf�� E��C"O,��F�6h]�$
�24$�9�"O2�[ӥ��?1��H  �H�0Zv"Ov-I{dqJ�EUX�tG"O���o2w�H�95���3"OH`f�D�	 3�$Y���"O)� βk?H�r�BA#���2"O�EC�ō�I��4�#dT���L�c"ObE���U&gvAR���<��|�"O��Y��?=pt94&�U�4:T"O>��E4�@��7��A��I	�"OБ92䈳B)�U�f��'��"O�Ձ�=c��3��6���a�"O܍0�$L�Nn��i7�y�(��"Oڹ��Lٸu���1NE�r�:,QW"O�0
���1�|����S�u�"O:E�3FR.G�i�T�W��!��"OlM��)ǁx��q�A�3߶1б"O�H �P�d~��ǅ[8Q:��@"O4�X�j�-\\��Rd�q�juk"O�"�_'b�$�S�#�,v��]k�"O�P�dJ�N'�xQ��	�
X��"O2��U���h�ׂׂ;8�@	Q"O���T�_�b�l|�r�p{���u"O��#&韼~)I 皛dQԬ��"Ot����<>48x�7#�xX��"O��ժ@:Ϟ9K�$��m���jC"O�`��%�X�
�#̷Sqҕ+�"O�9*sCߞ�>�+�"֘�d�
"O1zs��E��X6'�[�`��2"O|5(��%7��H�a���[�0"7"O�$`��T�U��'fɪ"'��b�"OL��@O߬pR�E�0 �v"O��+�ȅj���`p$�,<��s"O���AewC����>���A"O`\;�� "#�͙�/�;��X��"Ot��Ǩ�q�������,��"Od�����L.ƭ�&J��D���"O�T�%I̴j,�%+&��i���A"O4�R0�ɰV�cf䀦	�B��"O�	`��3��R$�&*����"O����k¢Z�@���ωH�"O���L�)8][��A ��tJf"On@�r-�=3�i�_���=�R"O"�;V��0_3.�زDK%)��� �"O��Q󉉮7[�yC^_@����t�<�Va��L3�T0s�I_ep�P��n�<p%"C������x85zWp�<)଒�L��8���XFp�Q,Oh�<� �k��9~_���޹+�&��"Oz��ĢD+:���Aޫ#�*��"O���p�r�ju
N�����"O�hj�aY�n�� ��GV��y�"O�$Z��R���2��	�/�V4�S"O,ث2JL91Pvs�F=:�ZA��"Ov�]G��ǋF1P��d�c"OQ�t�G�o�|���Dxڼ�e"O�с$M-w~�|���@C���Q"O*�[#��B�.�3�m�&2Ȱ��"Oҁ8EQ+ �6}`B����B"Ov�@%�m4��C��3IP�P"O~��e�V�	P)�eH�z�α)�"O���t� �Wg�������ְc"O�9b�KS!7���UZ?!�N�Q�"O��k� ��X��K�*��Z���B�"Or�� ����Dj�	 ��u"O���Bώ)K��4	ύ$,��"O���0�ڕg.̀�(
���,h�"O�-l��p��HК����D�d�<Y̚ ��0�쇎#D��,�c�<�"e@b�95�G�\�d�3��`�<q��	EF2\��S�Şd�<q���b^
ݲd�ŝ;T�[Udb�<au� 0=��=�֥Y<�4슑g�d�<���N��̙��Tl^6,SF�E�<�׫��V�$���Z�6�,	�Dg�B�<��DF P2@�˖Gk��Z�e�s�<��m��ki�t�C�P7.wҝB�IH�<�+�,L�cw0G�F��ƌL�<I0���@R�)4��#��H�<�4MI���<��HN!X�N�B�J�<���T e���&Op�\�/I�<AA
ʰ>Ev=P���O�u	�*�E�<	���v
Rx�,$({4)Y�)�j�<��3jZ��P�Q��䡳^�<1��I�	���!B��aU9;�\�<�(��iPC�O�:�*���Z�<�$�ؓ]�\�p�B��#[Pջ�ņ[�<�b��}u,�bc�L�D����d̓U�<4�;�(�pr�LiF^hs��
M�<IE�*�0����J
�ۗ�q�<iR ^/Tfjh�@�D�z!i�o�l�<���5XM򝱃KȉoԀ�`�j�<�C��l��1�#	e�I@��Lf�<!��"�:�R�(��MX) �Eb�<ׂ���!mJ����k�C]`�<ɤ�K�8�@[e kb���^�<IG��%���c@ f��Yk��Z�<!7m2PD���C�;��P���m�<Qц@1�R)�)U�Dpz�r��O�<Q�aU@G��s��I�q@�	%D�0xs�W8���so�TW��b#!D�xV�ҢA��!FɦcQd��/�y�k�G�XD��+��u�Ȩ�yB@�DT�k�"E� �p��G"�y��ɗQ.�C�݄G�f�a���y₄�,��h`�ٞO��Ӆ*��y�I\�L+l�x`��N"iS5�Q��y��ν���K���C�H�a��X
�y�m��7�|azԢБn4)��`
��y�c�>�Lu)%�N)5�4Dbq��y�MN�@UB��/�6+�@�"���yR�@  ���4`^�*�RԨ��Þ�y
� ^����J#�Ñ�A<Y�6E��"O��s �Ο+��؈���B����U"O�٣�"ͤ ɠ`�6Dؐhju"O2���ʖ ���OLŬ	�*O
Qi �W7�<����`8�m1�'X�C�AF��S�ذ.�~��'"O��@V�q�L�*��]E�<�F"O*Q���T26�ԸF�áf>"X�"O@��3FY�l\�u���>3]+0"O@%pU��b�^<	�1(��&"O�0�� ��8_�t9A�	
%>0y`"O����4�@����~	�(�"O.� ��K
#�����P�^��"O�\8���c����Dj	b��SU"O�1�,P*U(%�'�?o�,�T"O`8o��:���k��j�"O�d�� ���R���ϔ_���B�"O*��MV/\��e�EDR��>�jF"O�y���/*�P�B&G:Lg ��"O��p�G�~��ő	E���`"Oj [����Bf��"�%W�@5�)H�"O�z�.�=u�"�8kI�:v��"O��;�k��A	��Hd@�"O$���ͪCJ�m8FlW� p�y�"O�s�m�<z�ȣ�L�Z��#"O��zlC��@���G�{�iC�"O�06��U�.H;Qh^&��t�"O��&�	X�w`�MQ�v"O�\7L� ����i��CW
$�"OְX7f]�NBJXq�J˥l$�9�"Oh�qTÇ����ƈ�V储` "OV��A� �,�e" �u�2H�S"O�s �kG�i� (	.!��!�"OPP+�O�'f����g(G�ƠC�"O�!$���U3��c��ϯ���"OZU��gƳT�R�2��L�vnr��"O��eȜP4��A��6^�P� "O�YI��g+�jc�9�l��P"OE�3�Wx�z)��d��mF��q"O&+f@Θ:�B@k�B�f�v��"O��8��,C���fH�^���pe"Od�B8� 4���6�u:@"O�i`&����N��]�h��"O�dr�--wf|���C	.��$"O��ztO�a*"h�eKĸ/��(�"OTpag�;+����`L"�Dm�6"O�Ir�o��,��lJ�X���#$"O�,���Cj2-�� i�UAW"O�4��P#~��L��ST��){4"O��1E�6� ���B�|����U"ORв�Ӡdo�T�'䖪.���aw"O�`q6�Qɖ�c#�J�-I�"O�Qq��Y,h�(1�p�]�c󼬈"O��q��s�t��DZ@=	�"O�Xr^�XIJ��BRl��,��"O����jU��r���f���hAq"O*��)�BG�<z�FA�uԖ<�'"O��)殁��.��օF�g����"O��ɲ��.B�Ge�&T�
��U"O"���L# `>Zdb�B� �9$"O��v���cQ���/�lb���"O��`e	R1:�h�-���@�W"O����WKY��bt�M~��"O$ar��ѱIO�qi�.#@��J�"O� x���'�lD�P�B%���"ON]X�A��k_�u���8t���"O�buAY�P_�90�V�4���B"O��9��'-0H�����`���"O�1�󉐆B�̀�pO�ZwZ�! "OЗ�Dd `��.Y���L�ó�y�)��\pB�IGm�#�(���R�yb(�4&��-��7)ZH"v�)�y��Z0;�8
�i�!ò雴B��yb"M��DhrQ�G3H9 ����Ǩ�y��^ ����W�8�@���y2dGF�vMJ�[ZFY��P��y�#C�U�<�9f�7P�BURs��.�y"�ĔE/,}��3An@[!����y�c �����;�>��CV�y�����>��O8ز���&�yR�B�]j*X�eI�4(-���yB��bɸ��BG"2R�E:R$�$�y�%��D�¬0è�0W
	�q�1�yb B2C�1$y��Ј9� ��ȓi� ��B�6u�t�@ԩ^\&���ȓo��C�&�Ak69FӠ�p��{�N�+����|M��]V���Y�F�*q��> XК�Π
����ȓ1������m�p���o����ȓ@<��rIM0��gψ�l���Y����.K/l4Pc�
�.uNT�ȓ)G�A2@��0RtzL�RC^Pm�ȓ9�x聐"���,;�͒�Y�@�ȓ�B����o�aȐ*ʊ8��$�TeaS�]1�Jh�5�S��ȓm����E^�2��D34�ʕ�U�ȓR��*�l��T���vn�
Q�ȓ%�����X���y����Oa�هȓ.z܋t
�V�0�72�������ثK�����6?\=�ȓ!��" [�-h|��G�S2�|���&2��p1d&0Y8�qGgI2#������L�A2N%1 r���)_T��k� (������$ �AC��ȓ3

����U4��l�ºӂa�ȓl����
J�y����-.e�̈́�)�ȁ����zcd��i��Gct��ȓ%�v���A��A��qX�}�ȓf� e{��ڣ7u>���n5l�ry��hPs�%M�k�Nl�Q��6V\����vrv����8 �h|h���g�ąȓ{U.�B� ��L0H�����3I���X�� �F��0ܢs� �E ���>x���F؁0huJ��͊(��m��c�����u��Ub�DM!
�м��xoL4�@����-2v��}��a�ȓ4� �r�[z�fZEO�o�� ߮�kpND�|}{ᧇ-^�Hp��SV5�Qg�qfN�x��t�y�<a`�̺0�H��	�%K����z�<ᗋL�I���E�E.1d�D��B�<��4W�b�(�Dk�8�s-HF�<Q2b<����f�*q�m�<�$E�B�@��C�ջX�Q�2B�<�iV�t"8����=d���r�Xv�<���)"(1�Ю�;32�A�r�<��i��Q���ʴ9�JV�Lo�<y��	}�p�;�.[��m��i�k�<� �ȲEO3,a��l� �*2"OجH$�P8xa"���Q$d�j�i�"O��kWd]�dZ�9����3E�Zt"O\1xE�]��;��6d��<�"O $���/7�U3'�ř)E�y*r"O)Rv(F�(��%���	 PC�؁�"O���Т	8M�F\ ����1�<P��"O�	�)E���zg��� ���"O��	Gj�Y���i�/DV���"Oje��)U+Z*� 9��Dܒ��"O�PV ,!�|���F�-9 ʀZ�"O$�C���K0�jҦ��$��"O<y+���uK��/�#��Ac""OL��R/ɼs�M"s/9#���3A"O��cJL�:_�����[B�[ "O�캓��x��k��Ɵ7�yp"Od,FN�c��1A��{��e"O�3���#�F�3�ǘW��1 g"Oڭ`̗�\x�M�����`�,��"OF��3˵4?������|�&���"On��T�Q-M�$c'!U?Az��� "OZ����,aVQ��!�uq��"O޴QP��!M.�p�N¾+��r�"O�58��8=��|P`NT}�e�"O��bpl��<6�\sG�07Xޜ{�"O��Sց�!X��u��M�r'��"O���f�˾1((%+P,���I�"Or�;5�N�m.�I�J �;��"O��:C��v~��`VD\6 �5�D"OҼz�'I=%�h3�V+Q��t""O��-Q6\t���!E�C��P"O>�֯3ԅz`*�b�z�hF"O<���'���iEIW08վL["O�����T~�̂���L谭�"O�ؙ �V�<O04��ȟ��@5Z"O0�c�¨��X��)%�bT��"O�f�:m�0C�P b
��"O���M��� �sLL�5��<#�"O������ed�qXA&E-(����"O�]CH�$W��:�䁌HD���"O�p�D�������Cχ~ 
-��"O�e����hHe�.���0�"O�%��V'xx��Ɨ�l�7"O��It��4�P�V�HL��"O�5xFn޳G�UP�$��.
�.�!�d��3�D�H�Z=3,D���+,�!�+4�r$r3g�
B� {'뚙Z!��t����O�gv����q.!򄂣Xa
�k��s��ɴ��.%!�䍠-�D��V�z��h�%(�&!!�����X��{3V���ޝq�!��VQRVѫ�ݵ.+^xI���N�!���F2�ek����NwF�б��A�!��; ����,O",v��#WI�!���]�vH�c��
B��:u!���a��) ��Q9A���"G�R�!�$�G�`Ej�jɝ9��X�'Z�v!��הe��
�ΐ�=�B��FömL!�DJ;��a��M�8��b�[%5K!��
/]��{b�	yr�w�U�c�!��O�D�0�\4�B� ����!�$]s�0=`�DFV�bw�,M�!�ā0)�4{4G&@�$���u�!���"�Xdkċ?0�5��/�9t�!�� ���`� �fԒQ�TP I�"O4� E*M� �D�0��^T�E��"O>�a��[�*��ț5M�%vP�5Xw"Ob��膢G�\��q��Z �Tp"OZ����^	"f,��a�_� ���"O<�c2�G�J ��@ƙ�x
,0��"O�%s�J�X� <�U۳{"�"O8�0Un�`_�$MүB|��"OR��"/��o�`P��
��pr""O�A󀭎:S��Mn�/��e�"Ol<��N��B8#vǎ)�~=Q0"O�Y� ���,��Dl�-3^�R4"O2Dp2ѰS�xE��>:+��@"O�<�VIE;P8��j��S7)p]�"O�Ԫ0Ĕ�|8n�ҴO��ou�@"O�u���̜:��<��I�:��C"OБEE�G������ELr�z�"O>��MpW�$���Տv�Ʊ�"O]Ƅ٨9��b!^�_lE�"O��s�����C��.]Pl�6"O<p��K�0+q��[sab���"O� �a��7p�<��U\ *0"O�	�Х8^3�X�@�߲l�^��"O 0���� @�2R&˝+ E�F"OP)�M̡!��yF�TX*�I"O��3q�B��p�p#d'C�`S"OZ� 1��]C ]y���z���s"O�iH��V,/8j`+�@�n�0���"Ol���bЀЧD���&eڥ"O� I(��_�����S�=2��"O~y�P�Ȅ&xj���bʡ~�d#C"O�`ea��X�H����|mL��"OP99��&�]�!O?X�g"O�Í��N���
��jF��2"O��\iz"�Z��)(i΀+r"O�a����\�i 'N*uQ���"O�<;W#�
���sgfӓ�!ч"Oz��g�}�V�SW���Z�"OX��g̀�Po�;a$_:�>�Z�"O�Qس.R��z�)�9L�ʜA�"O�B�K��H"@�x�	��ꘪ�"O�`����iܤJ��^�a^���d"O�t(.�,u,�AF�At@ {f"Op���yI��@�� +o~�؆"O iӰau�~$[&��	XwD�
"O�H���E���[ k٠A	��̥w�!�L79Y�h�%#ƨB�zxУGʧT6!�$�uL�MJg.�$?��ᒰ�C&/!�$�u�0\X�J�?z�i�M�
=�!�$�,��(�n���*��ސp~!�D�:!�ڥRD�� $�  X �A$u�!�$�& ���+�^U0��&c�A�!�93��]a��TI��e��gQ!�R=UۜͰ�#OR,��Z�(E!�I_�9�󋘘Q%�p`���,!�d�,4{��x�'�8i	���.�!�dѡ2�@I���ǔd���á��!��A�z��b��L�q��
nB!�Ӯe����I	�"�Ɗ�H>!��4nQ��s�!S?��-h���h�!�I�l�eH�@E*�1O�8�!���.)���Sƃ*E�h)Tn�+"�!�dA'7"��X/?(Le{խ)d�!���)��la�"{�|!rgH��!�� �h�初�^�&<���]lL�W"O���Ƭ��P�<�1G��/bFq�p"O��k a�/�n�!�f�Ld�Pr"O��+�c�Vi`50�e΍l��y��"O��R��[�V�H�5�ȫ(��1�"Oh�0��@c��#`BYY���	F"OVHf��@����j\����"O�3'�Q��V�{�c%��t�5"O@(Ҧ(�gD`����(L����"O�Bw��;06�h���� �t�C�"O��!Ѭ�&:��ʔkV�'g�@7"O����"�-� 놝nG4��"O�m II0T5pԻ��QC*�`"O��`�Y&���sp+�6x.z�!�$_:,4��5펄@��$�`�p�!�dø5��S%*���P�OF�Z�!�$�]�
��!�D5)��5���
�!�D�_�
$qg�����,	5�!�DҪf,գ�	�L��=R�+�)F!��wL��X!��z�$5bӨ[)3!򄄥Μ�@"� O�ZqԇP��!�D�(LPa�j��2D�ci�.(�!򄕤g��(��C^f�A���S !���l8�������$t�!��>bDzГ�L�f�uJV
�/b�!�Dŗft�Q6i�<8L�h/s�!�D����ٰR�R�G��N�!�$̓#�H3CA+o �m��B�!�d OvI�%���$�RdD�u�!�$ɵ&�|�K�87�j	��R��!��KW�V5["��p�H��"�O�!�λ}��i�%7v��ϡ�!�d�5��<y6�H/c
Hдm��-�!�d 9P����]���Ʀ�k�!� �yK�DëG����[�!�$	-4|�|���	�Ȕ|����<,�!�G�-O��s�_�K��h�3@̗y�!�$�*]�4�郋��eɂ�E2B�!��Z�D�9�tK=7�)�0kL�x�!�dA�.u��B�^�HJ��p!���hآd
@$�7>Š)��e�I�!�DP�o~�Y$�G����	�+U�!�d�9G�� � 	8���1U�D�@!��\�VX��G��(,I�b	~�!�D?��`����|����ٕ!�T��p�TD�?d�]�.X<a)!�$� |sE�M�8����g��!��t��v�� ��	�H�3 �!��̑bA���P`����xM�!!���'^0��D��
��E�"?�!�E�{
pdr�ԇ�����L�!�dK�b���S�(	���C�a�!�Ć$294yP�κ�"�
��B�!򄄪>�Z��(N;B��!P3&N���'@nKvA���ؓ��U�/Tbԇ���%0��F�b1�pb�@XX���9�����J�'��Պ9[�����:����&���F�C?\5.ф�50.=o�
^��{�Nθv�P��'ٞYQpmKU�xp�]6g�@q{�'x�!؇gF2Z>��P#�\�<��'\ �R�NA)�I�0` �v�'��$S荥oj�@p�!~� `"�'�芷�2H�����R~�ry���� � B�ĲP݂�H�Ԩy��`��"O,�sCl)�d!s�h�\��٦"O�mq�ל>JX�u��4-F��:v"Otx���R�z��,S�&�3b�qI�"OjwI�-o�X�c�J�����"O4�SvC�@TQ�%�t'�!��"OK�RR��!�::~j�� ��y�9&f,�
�H�>b�h�ZP/��yg�&,$�D�T����`G��y2=}�} �΋9`�����K��yC�A.|����Y�p�կ�y��'E�V�8�ƀ�;�҈��m��y��Y%,�V��bF'�h�J�y�l0^����VD(\֬��N��y�Q�U��zN|�Y����yBE�/^x��Q�\��Ґ��'Ĩ�yRK�8g����pk�hѲ�y�ę��y�5m�z,H#ǩ1����%�'�y��%��1���I� (CR2�y҉�3i��u��$ [6��V-ސ�y2�\A+�gޤz��4J��Y
�y��ªg�h��쌌nSIz�A�"�y�f��t�$|#G�X&�q�U,.�y��J9ni��*4Dau�ě�+L��y"AI+gj�%� �\̦��1���yR#9��I'�V�L1�aj?�yb�8> qc2�I�^~P���l��ybhQ0'�����[�W�S����y2M�]�^�����('D� c��=�y��%F�#өT�F��5gP3K9!�$x����a�D�}Ĩ�n!�D�xv��a��H�^	J\21H��S!��vM�`%J�m0����F;p�!�
4AD�˖"2�P���FVX!�\9:mH�����f|SR�82l!��0�.��w �8���3ņ,$]!�$�,{g�N��\��c�{P!�D>Yߌ��#/1��q��#F!�دW`"�GS/b/j�ꣃӐ0!��	�N&�3gV-�m��P��!��#0�0��X�_�����i�
�!�$��.\ђB��L���$��G�!�$7mh����a�4\݉2��I�!�$�rOHa��#n�I!K�\�!�DU�'�"L��Ç�d2@y!�d]�'�yu��=(�Tq�!�X+!���#5��!�"T#~�R�+g��+�!�	�v&Jd�p/ڙ)�p��f��!�D�4X�aб��s�(d'؉\!�d//T�0&��6?6\)U��/b�!�d��x��5�j��E��`Z�FN*P!����[�+ܝfn����Ee0!�dĴ9��t{��	`��s��U!�߄?Ò��� ?z١�LT ~�!�䋢NS�q��/t&DEZ�,S:�!��'1�xlq�W.���,
`�!�I�.Dh�2��Y��Q"v-�
%�!����-�&�67���pMe!�$ҵE��H�#��&�\sS4=�!�'~�e(�W�x�[���Q�!�D��7<��V� uq�=��(W3r!��d���H�$Pjb����E� `!�;	�� ��X�d\�iX�#,(iџ,G�D��7s<��q���,�P����y
� 
���.�"Bab��S�Q�S"O�؁��Z;�NT�#4�Y5"O��
���q����
ݠbf"O&�;��- 8��E9ª�0�"O�aꓭ��V�BA�r#?D̙�F"O�� ��T�tLc�B�d*��"O���S/�=T��e)�+��A	�@z`"O��s��9�	J#+�M�=i��D8|O�q1l�(B�ܵ��)�L���"On	�Ɖ��[�D���-�+��E�E"O|�#ef�x���d�Z8��U@�"�c������D f4$��Q#}�$�Z �O0#+!��J�� �G�
�J( �m̮!��M��M��NP|�����	ؼ>����D"�D$ �R �ѯ�`܉��Y�V�!�Q�,���-�|�Ö;G�'��L�S�'�*����.Hm���!B)d=�ȓ� ��=8�|��Νd�=��It�42�D��Ō�h�B� a�'W�C�>�0�b�͉�i������m���<���T>�k�.��X*��FməA�J]��:D�@�Ë���@
�)	�wj%s5+D��� h�����V��"�-D�@�)��m���)ڭp����$d�O�B�	
9X�-ȴP�l~4�bu�Q?[�B䉷��)�D�|���*�B.jB��h����ܐ(��:B�I5)����U��"�=�W�ZB�I�;��P�D����z�O,3Y ꓡp?��K4"^,�I3%�2F[v�10�E�<�@��U�"�h�-B	f�
2�Z�<ѕ'�5<����U*H�L���Y�<����@�΁��&@05��;Q��[؟�2�'JN� 1ϭO�����̌�p(J�"+Oң=q��D
PCN���k�$��@af���Q�QN>�M?1:'�I�v��j�n�>̖(9�9D�8�W$�x��;$ �X���;��#D��q`�Ц+[F C��D2�M��$D��b� �?Y;�)��A�*u���0$"D�T� �I�yD����N:��c�#D���kD�[� �ˣ��d��!�4H#D�,�Q�� a�Ւ�����y��&#D����L6ͦ��'eU�m���;��6D��`�
Tk�8�D�n�Y��8D�hӕ��O>�A
!c&Zf���6D��
V瓄,��I��(��B�$4D�(p��)�"U~��g�0D�L�C$24��+�4���V/D����܇�����ODF��!vA!D��1d`�8rW�<Xg&�,z��0�A?D����M�/r��@g�<^���s��;D��Nѕ\58��	�v�N��CH8D�Ԩ�!Ǜe=R�!$���8�Z�4�3D��*��m�jE�Dd�.����n�<y,�/=����T.U���k�F[��ў"~�	�W�~�k��P�RxJ�q�lXj/B���0ړA�H��K7+����c�������hIb�	�\��ZSs/ X�<�ȓL���g�&Zǰ��3���*��ȓ@H�%H�� C�l�A��)�����H��ͪ��2cfi���;���ȓn��y�R�6R��4��8����w���P�A�8�ر5q��E~��S`h�YQ��O�~x�0O^��C�)� ���2���@��m �aŢ��"O�Es2�	(=���M��S�6'"O�(�b�X���쇖3��YS�x�',9 w�Ԓ���P�E��\k*u"�'��Hi1B�M�|�а�-O>&`�ٴ-��<E��4]��b�@?@�̥��gK#1xZ��	t��^��)��V5�5E��l��?v���D=hQbsU�[��Yr���Nx�$�'�
��O��B���� cքq��1�	�'#�Q�*��>f��d��{������6,O69q��I���(� S�J��%��'��~,F@B�@�F��\��B/���'dҰGy��遨-�a�H�$��=f+��<��x��ɺv��	�֡�35Le{$�,\�H�O����?(�t���GS�6�����`ٛd""B�ɝ�#˞�1\�	���"<�
�Z`��i��׶zX��9f�� d��'��}�®'�j�`��-Wfi)a��y�m��`nt9f@-`0�Y����yl�8d)�K��F1 v (�b��y�/E�V[�x��A�;��0A+���yB'P�6n�#D�
��ɪp��6�y��)z�6 C�l�tĘ�J�/��D2�O�к��Da4M��M­A��W"O��Gc��,)	���=9�2A""O��鳆A��6(��� v�L�ʁ"O��@��l5�1h�aˍ=�JU�D"O"��ąA�q�Y�AA��/5ޙ*"O�8H�H��A��%O�b4���"OX�ĥ�|SЉ GY*���Ȕ"ORX��	�U���̕�B�*p�"O�\
� �b�H�1g
�hל=H"OF=Q�k�<!�̰
��8�B}1QcTF?��Mc �{�<E~2$`�p�����<� ���G�Px�A�',�� �at��aD�4�j-x�O> �E�P�V��9��K�+<3(!�b�|"�D�O�b?qRd�S�0dlL ��љ�N�{ֈ)D��9�N%w!P�;�L�!�6D��&D��q�����B�6͈&7�T�E$D����+�Ls������
�M !D�h�2���VF��HFO�@�C#9D��c!�R8:���qs.��c�7D����Ņ66�L(P��]���k7�II����;��]Iw��x�h��W�BC��1O��!�7�]=U*���$�x�&C��=�D0ZR�
�l�n���ټ/��B�ɠ:����(��W,D����$u�C�$ȁӀ�m��:��(C��C�	.<��Uk�
٨���i0g�2B��&�&u�����R���`B�I�(k.I*�ϕ'WI�;���8��C䉐"�l�֤ՠ�	&W=*�C�']#,���C�p��ÚL�zC�5���CX�<�sa	�<C�	�+�~5`�LKY��ɔ�pB���%�G�֍��Ig4�B�"O�M�e��E�[T�3j� �B�"ON5��R'����N�2�"O�|�W. M\h͡T�ϭ6D����"O�U�D�Gyt���ϓx��J�"O �K0(-I&ƴ�T~���Ȱ"O9�n�,M��`� �� 7_ܳ�"ON�h�F�0y_:��fX9{���7"O@���ݥXdb��&r����6"O� ^5����U�)���ӔB��;�"O���4/�bHUc�YҨ-��"O�;�L���ED�4Ĥyr"Oέ!�&�zP$X�s`H�H�r�0v"Oݰ�e�9�d�u.�.A��	3"ON5��ā�NL�R�H/�PI�"O��qJ�]�6I� P/M�L͂V"O =�D��2l��-kR�&�T��"O�ͪPg���䉉W�˴:�,��"O�)���I'@4�fi���<���"O��GVM����sM�4Ќȑ"O��*�ĉ�4�`��˂�,�8[`"Ov�Je,�aޤX� X�$��1"O֕"�h��)�6q�F���Y��"OP��nME'<@�]7mv ,{�"O�]P�k�*"��� �
O 7�T<c"O"�hRf�%w����J��p����"O���a���[�bL1!�(=��!s"O"�P��	�3��A�I)Yr4"O"=C'��=I�xjeʣ�P��"O� �PdS�m:F�rV � �DX�f"Ol� QD�+:Q��h��+�D�S"On|�-@�Z�^<!�f�%V���H"OZi:��ůd�*sU3)$X�Z��䔰.+F�"AT%D�26N��1Oٹ#4&HtS�	Wtpu�b"O(=�0���UM>�8��b��D
P"Obʁ˄�e똀�0I�6�$�"On�zk�0�x34GH�>A�"O�պc�֞L>���%�?��E;�"OԵ�1nE�yD���c�;�F��S"O���ӂ�5���0��(L��l!Q"O���OC�L��%�6`�y�0t��"OȨ;��A |����R�U���q"O�D�Q	�̹���*��L�"O��N��_�z�ٕ�F��X�g"O��3�N��#�,$&	ԫ�0m�t"O^0`Cl֗1��<S3�Lr؄��"O�a��4��0����KRP���"O4�ٓ�9���rm>(\�0A�"O�t;P�P4|L���f+^G�*p"O�d�˚�:G�`����9��KB"O豺���9 A�˅W�N �B"On��'M8X��a�)2'�B�A"O�K��ĕ3��q��b�N��"Ot�P剋RȢ��'	8��(R'"O0�6e�B�p�J��j����"O�6(5y����[/1�^S"O�xKq�:"�v%+t��W��u�"Of�i��6:�6�1!cۗL��aٖ"O��j��=��a($j�"O���L	5<PҠg��B�Q"O<4bECQ��İ�O=����"O��篁�V�@0����:���q"O�{���z>H����5��8"O���Pn_�8����1[�^躥"O�`�A��70���{��L�e�n��b"O>��&�K9B(h�HE���h�����"OH�sf��>s�X*��.q\�%{�"O���f'�Q��K5?Ox\�'"O�ҶfƊes�t�F�J�<#BUi3"O(M�`�Ń@?��Y`*''X=��"O���WDA4�b��'i�,+XH" "O��+�%#+��N��9/���'r\�K7��Qsn",)~@��@X����S�? �Ms��L�o��x��L�Ea����"O�sdk�9��Y)��J-��:Q"ONE��ɏ�J@
Yʐ���t���S"OV�c�˄u0�eZ�"Whm�`'"O^��E5ܔ��a Ğ{0`�B"On��B摮�"��"��M����"ON�����t4����� ���sU"O@5��%T>n�f����`���3�S�O���a���X0�d�"Sv&B�I8I^�i�Ɋ"�rPД��7��<q�j}�x��f�\����҉��*���ȓA2H�$�Ҕ������ٵ#�`OB 2%J�!dQ�=`�jũ=�B8� �'�b�;CD��:�b�fI�nXBQ�%&D�4 uböds���!��#(B����g3�#�HO1��e����S	�U�v���)P��"O�݋0Ƒ�|�b�2"��3+���AW����K�<��>���I�Kc��xVᎃIc�u�`��!
��B�I�r�����;�q�e��"�H}y�OF-��+����<�w�.P���"e_�~"P����h����O����֯t�d�A��-�ZQ%J5b}ȕR�'ڥ4 �
�J,C�m]w���y�=?iW˃5J�?U@bD �;Z��y�ˤuH���Ю1D��Q�F?t���?]�!� �>	�#�}[��DI|~J|�'��Q�rM̮��� �拈gl��
�'�\h�2M�%:����׻~�B�K��%?) #�.t�T��)Nւ����5\��aN�-fQaz�+}2��OԲ�Q( �XHP!a��ܠ��'"O��aP(J�=I�ؓ!�[�_�" �����Y���O�QG��4�����"�:��'�t\� �6;�m	���vo��8����pX�0�` U=(��j0#�"7}b�h�l3D��[�@��7 ���
%�cԉ>��C�	�i��a���J�����1x���2��$y`�\�D�2�j�P�o�&w|!��	.�����D5�D��!c�qO��=%?=��&�3^�2�ա��&�"aK2D�0B�/\�v�*�ψ�I:|P$7D���ӵ4��SU�	�Y�����><O
�Cu��� [��'|���@�4����%	�o�P���'�>�3�N�=!~�����!o
`E�N<�5���A�ЪTMRg�O�]�R�?m���#jS�eD�	�'���	�)ަnװ�kPG�.�X��0���*�>��K�?U�>�>�OTe��.T�v���٦��o��9'OPi��N�>
n�'�,n��DC�OI]��� ցy5B����'���AW�U�6 �&�o��I��$��Q<Z���YK�a�g-��?qiD%T�9�F�pM̹��H=D��y�&3z�J\�FNC6x�Q���<!A��8	[�����ޠrgе���>ҧ$쪑��! ���G	�6Q�
M��>�4MہN iY���j�0 @�̈C�6�����m�,[��O�3�	D��ٺ��,ڌ����ց_ ��DG����bo�3*v��2�e�-O����R��(��۲��.6Q���T�'e�����Bk;�����+�J���FN��@�D�A2��!d���}mnj�Hܭ%��yR1̘)�4�@&�`}���`�`D	�ř3�q����l�>�O��X9��sG�6�*��_\y"OݝMB,��J�x~&�ە�Vv�1�8ዥI�v*Y0��&F�z�����PPw��<qR���E��|�1����O�$R�/�W�ֱ�#h�4 �J���务B��59����9�"X;���}Q��O��U�ک�c�B�"�\��W��#F�0ՊQ	C�}3�a�GB�I�qT�Ӭ�:���'D:݊A�d8��I�)l�\�e�bhHTF �]�&����%Z"f�2��D�c,-�u	��X�e�k��J�_g8�X��	���1e�E��0<)��F<F|�PdnX�]#ʹUȁ�
���JA��;h�<A a#Ϋ$%�4� H^� Ԩ�6�R�8�B�"K 	���Ba�M;i�:Q#�) ,��`�i�Y�,�*"�p�І�	X�(�N�T��a�*��%(���3`��a5D��/ܠAK ��	�_D��a7�XI�5J�lW����!d�ːtՀ���`�!1�`y�P힙A�Ez�	�\��CR��7
,@��)�1w�z-�u�]�!LJ,1� ��I�R�ɖ _ ��#�$��2"P���㕈6� LY�C٣*�����E�HcUf�C5���(�@8��H�a�  Ӆ�	Z�D3�C&�(qNC�_��h�E�c:\9�C��$�;'h��M_Zl� ��4�F�5�Щ
(���I�j2�y"�(	<0��#l?�, #J�_�l� �W���풂yt�����
�h%�;�&1�W��.X�HCp ^^���GSf�nZ2���R�	�;}����.���O�����χ�k���R����S�ȉ<��px ���M3�cF�n�P"I�4㼌	��K*=��	���(�0�.
V%��JA�ڜBΑ��8�@F�
F|q����Y��+p��
7~HӐ$֤~�	�E`H>�~�P#�4�~���,��k =.�g����%js�A'*֘)iI��u���kbX��'�Mo�r��%+Ӥy%�	�1mГ����NW�[�6E�g��	Γ���R1�V'J�X�c�[""�,�a��
n��(���[�DԘECS!�\ܓjͦ���c.}��$G܌i�AƟ13��T`L	0�����U�wxL�B�Ƈ٦�a�'s
�걮O�X���@��k-I���(�U�̌5��IQ�}��\�W�Ƙ=@Q����ʷ	�<	u���-3tT��%6������V^ݙB�ǤB�詫pmLF<�8�b,@��THGn8��4CM .�����p�J�Ӏ�-ғlnT���0	#��r �0^y��%��!Z(>5��BX/ �F=�E�[<WL9��2(��ΓYv��o)F�H���ᘉl�^@��� �✨����ж�ɶD,4��stFX{>O���B��]�v��$�P����{rX�a���i`@�4k]2��'�P`ʖ��"�l�BA��F��F�|aA�%�a����.}��K�(��i�+=ڀ�OU�
���?v>�yu�&N����_�%��u,�$38 X�O�= ���d�*�qa���l̘5��p�Z.Obe	Wk�=�j��b�X'+
,��a�t��}�Ë�O�}��A��^du9'kߔ8�pċ�#�.0����w�����[�&(<�4A�|�q�a [���Ұb�J*�����D�=pf�1\h�)���d�0��Ύ���T�&\�o@�E8f��m���@(��_n�9�Ƥ�f�(0�f��@}�N�S��b�ég�ơ�8S�� 5K@i�'����X }�]��.?y+�3XyQPAA& �ȲfU�w���cT�92��
-h^EbǬ_>BI	��&��Ɣ&�y������)܌����T'���8 ��%�êH��ɰA1�ӧ}\�l�0�E����a$i�?��� LD#l!R��@�D��M�k���^��"����ԉ�8����\��C�g�Uy�X�pA��,;p!CY�"t2h�g
�� ��c 9��)�V~�t���̓*1l9aټ#p8�У��[=< �.+��Ѳ$�:�he�U������i.Od�D{�Î,Yz�\�VG�X�J��#kS� ��ݚ%gO�my)��Ȕ�b�R�p��CG
5;�
��
�]�$`��:|�p���ȇbT�zv@ʼVJ$(�s��([�tD|"��Q�l�w
�w�du�'?�L�0*�Mi�f��{u��{&C�'��ĳd���n���G�X�b9�T�P�>Om �VL@�x}���w�~4�q�5D�X�v闏u��M�� -.��Yk���5>m� �^.����o[�~��aj�F/K�,�%BZ�(�@��Q`�جL�:<�E�Z�*�����(�%��W�p�N�G�1Y"��2.��Je�@�Z�д��!L��XAm����2�f"ҊQR$X�\�r�`J�J���� iU��W�H�P$!�a��zڈ �v%
yg����ɑF/z��W��K �ɐchњ�u��"G�~ ���D�<������:+`����H�N�7�#7<�'&�@�a�).N�BS���]�R8��I(,H�Zc��\��	��\]fC�k�,���-��r�Ni+l�e?|tҶ��ل�B�mT��ZMF�O�"��MI*w�@�x��I*v���j.��z��)7Q42���ԛ)��L��R�¨5S�NĦ|�����jF Q	5)`�G�]���ݡ-�v0ՠ>h�"a��J���R
�A�'�r�6]lX]8����ER�{��
�,%n�#�L�ufP}��+Y�2�� Lav�A�TR(s�nIz7�@����Y�G��N�$���G><&mzlR3}�.��r9:[d��#�il�e2OUr[@�gJ�B0��%e�RQh�'ps��<Y���G*@�S��L�4!2�`B�%r|�	�hB8ۜ"tLQ�,�P:��X��,��!C�A�"M��S��ĺ˶� `���bq0�QG�լb`�0��B��k��뉘&K��8��'���D��5�&M�SL�64&��Wd5Y�|�H�>Oдy�xA~\�e�'=VT�a�H�z�r�HjP�x�}"b��U8�O��jG�)��@ӠÜ/���REfNR��V�58B�I8]X�q��9�Z�Ʌ.Z=}�^C�ɇ2b�q�Ǽ[�2��͚�E��C䉶/,Fz�O���P�MU� ��C�i�Lq�:��ؒ�	
?���)�'���*�Lӆy|�����)��
�'��	&� �4��\�"]�a��'ژ%���[/c�X��Ed��M��Q
�'�� ��"�� k�#K=�F�`
�'4����iA��@ �Ǉ{�Z�']0ya� �k��\)G�N������'m
a��0j��(��PzÔY�'�6�K5�ˮg���2 N+��\��'�$H'C� I����mJ(	�i
�'�<�1Cj̠D���$N��L�R�'ꬕ��-V�pZ|���	�rŠ�'}ԩ��a(\��J4*Ê?J�Q�
��� ${DA�~`��e�R�d�<°"O�L�oΝV\0�A�'/����`"O��:6GE�.�P�qd�;k�&�ʃ"O�,r�G�E;L�`잸+��Ŋ"O��8"���D����v�N�;�и"Or)cd���^�FA�@&��v�$�P&"O��b�?�P�b�O� Tl�f"Ob�2s���Fr¯�|NZ���"O���!͔��֡���9<^���"O�x�IB1�dX��'3"��"O�����up2�@�LW�o�(Q�"O6�[u����⃊ͅn�t �"OF������)��j_N7
ɈP"O"��BH�*l��p�'�?��"O���b�A�6�Q��<i:ʨ@�"O� zb�S�ޜI�5�ɏ��� "O�X����;s�zh8�bܸ�:���"O�	��׀{���c��G�ܐ��"O��ҷ�2�JغaN
�B}�p"O�ec'�S�3t(aYFtp�-�d"Or�k��
0�`�d=s�m#�"O��y�EC�+ӢEBh��o��)�"O��vF�j ����VgD��PP"O����D[�=Pb�Xn�t�"O��se��L�AƘ�ؑ��"Oޤ�FŖTm��I�nP;�JA��"O�K�bW�s��x��j�
����"O��ӳO4K+ٱؔO�2���"O�T��k�A�b��!���`q"O@`��PIPe�rl;����"O��p�"�/>*�:��[J���"O
0#�H��)��Myi��3�8ѓ"O�)�6J��5;L1����/1��A"O�m��߹FKr�A�UF��I�"O�)r�F�h����R��I �hF"O�"��Q�!��0����0mL��w"O"��͘�(�U5}�T��5"O�������ÇG��Vu��"O|u��`ˆ"����K4P0�"OF؆����B��ˠgX��"O֔���x����A���6P�5)�"O.yC�F>3J�� ƽ3�r�q�"Or�0���:Gg|�J�����\q"O.9��[
tv�Eͅ�#"���"O�Ii��[8k�~��q&Q)W�"OhˢiOV���kĥ�~���F"OZ��t#�:�y��DA�5�}"Ob�Y���5N�q3��a� 8�u"O�᧧
�眘ʧ��ߜ��"O�cc熢.���+��É Xe٣"O|�q����"�>���O�
4�q��"O, ѓe�6<�8]�3B��!"*��"O�)�/ÑZB�aZdc�^��
�"O�T�pa�,wV1�b�
�6@d)""O( ��)Q;w��*��zCZ��q"O����V�$e���AL1Q�|��q"O����mH�E[� �.{����p"O�`(�k��	h��_l�!"O��3��&�ޘ8�n^>:��"O"4�T�O�A2��HG,] k�J��"O�%�'L^�1�h�k�j�a�"O�RqΖ9�Ji ��-k�@�#�"O���t.D���d��'Pe+2"O���㘮0Q��t�
�BL�0
�"O� �X#pB��.Q��W�j0���"O}*k��j�N�ɢN�
#���t"O�%3�cS(^�м���Z��6"O����Y�7v*a�W-ϼ>�)�"O��` E9y(JG��*�"O������Ts���$Bp\���(�yR�E�N߰�iFm o,�;�
���yR�L��Cvg�&"����F)�y2�`+<�5+�'�P�`lU�y�e�>�0dC: �l,Ƞ��4�y�&��T�Ґ��o�����:0⟙�y��jL�J�+�(����͓��y��O<>�A)�xъf��T�<y�7[ ����T2 ����̓u�<i�ȀM/p�	@�ȭ(E
��g�v�<�t��^$���[�:�0T��z�<��I����ZSn[&����\�<��b�+z� kPQ�"0�� �Ȇp�<�N�MS {�AG�C�QP��z�<�����.\�� h��ᦃ�<��ȑ7o}����)Ze��( iPz�<Y4���N��Z��O`T Tu�<�qQ�m]$�р��#b��Y��\d�<�S�Ԟ��y)#!�R�S�Ȁy�<Q�C�5d�B�A5
Ԛ�Xu3�(�{�<�����i����s�J����R&�S�<��-ӿ#Xɪ����ET($hu��M�<���W�$�(��[vO� Y�n�N�<�S)7n]	�����z����EW�<p�ʾT�P��1B��<Nx��V�<	��R[����CT}(���AUW�<$L�:�z=¶"j�n��DDX�<�@ʫ19*R��n� �C�#q�<IJ����"�H��"TԨ���{�<�#°_��K����7�콓5�Oo�<�1�FI�����4�Xā��d�<��ߏ]���(�AF��Gl�e�<��b�Ny>M���*q���Ir�e�<	�����i����$:0�(jCg�<Ɂ+��u�rX)#,U��	&P\�<�	��~
~}3��	�B��!1F�Z�<�x(�e�Ժ.����uŕQ�<)D�A>7֐yif���'1`��#�Lx�|aF� �&3d�(O���GBS�H�����6��U3r"O�5)�ݸ��������_.���f�x�g�11�T0!A�P��ȟ��P/rp\��V�͒Q�"Oj��!	�S��.Ja h��@�5�H��Or]*S������}��ɰq�=E���� ��Ȕt��|����Bމ}��x�&K��'����GnB.m&��gKH�k�����Y���5��
HY�k\�R/N�?CLV�"JA�DĬuF� �O��]sWb��i��=��Ξ=���{�'ޜ����0t���{�X)	8=�,O�U˃�.f�2<�D蒵d�.p���	�x���Bs�����BB��,�!�P8 �[R��
d�z�ԠC�O����O;&��H*�C,�����{2�ɂrr�j��6S:��������?yv!	���A��?5���{]pD���[���9fM�0���C%�t��a�iʃSa
��CIT8~����%#4��(B�a�ΦV����S@p�b�����BdĔ>j�9C��%��ɐ"!��Aӭ�<�t,�}��L����nϮ��v��<���j��Q&�IY��i���(b�X��U��h4��|���۲q�mI����B��T�ּ?���c`�Ui���	5h��Ӊ�u��>9C�	�@�zi{�fR�������;4[��`t��4dn�y1ʙ>�|���
A�pqK��Q���P��91R�����U;uo|�^`�X�/Z�iz��ʠjݻ5=���$ح��]:S��M!�`�%NغK^LS���'7>p̹ĂH�^k�d�5V=�qR��H)�H��J^HC���0����
����C)D�"���'�ND���O�J�	�.]RPc
� �pK��ݕ }�����D,H�4�H�.�M)��عY�N�BĢT�Nφx[��]���ӕ�կ@%Z�۴�������C�Ua�}`�)��3� ���#}��S
`�%S�q�.X ���<�07��lP��wo�����x�����W�7�L�y��;J:ո��ьk�h�"��rd򤻴�9_.2 IT��	+���A�ηv������C���2	P��xkwJ
8\(< ���-���(�4q��N�
||�Y�L&rIx}1s.ʑ ��a�g�S�K��&��|R*�ZMv]*1$)]a6���Q��e�5��Fx��u�Ӭ����^�\OvY:��p��T���E{H���E{(t���M����u䍸hR����1L����ń�;o]����X��(+�`��T:�剓���t5^̓��1���E+����W�I����Ҧ�Y��F��q��z
���!
_.�MK�_�I�j���J�h���[P�I�K�d��s����%\�~���_<�Ժ�DX릵�ǁ/Gp�x�E(<�V����H:;z�Z� QTڼ���D+o����ӧ���HO�T��M�`<�A�O�>
*�lk7�_#��p6��r����0�
5rȤ`�5�L?�7G�O��SEî6^��5#�-JG��0䬗s`d�Y���X9RĊD$.�O���0	ۅߦU���ϩg= ���@[���E8�-�
���b��r�扴	%��I��1������JV q%���-J��e��hדe�bE��c�} dqp$�8&��d[�cUqF��&�_�q!�7T��?9bN�5[�
�;�9vAZ�f�)%�t�լ�<@�X�s��Z�ͪg0r�Ƶ��Z>x�\��=�V���g������%ߞ�#��T�j���;��.s�x�@���q�r��F��5�ᰆ�A���mc�Fj+ЕC�#_o��8`.=�%tJ��-y�X3���f�!x"G��g�W:j����NG�5�٣�A/wSvŰ�'�p�H�4#yR!P����[�	K7_�:;d�ȶq�,]�Q!�O����1R�|�qaP1T�F	�Fk��d=sŨF��oZ(`�l�V�b��,�R�X5���w�6|H;N����*y��p҅�'�V�#�DS/ ��bDdрo�48r��[Ԡͣ$I�@�O�Ȃ�_'NQ:DXB��{ �7I�l��e�,O�!X��$ �6D����=��L"T剤B�1h��ڦ%�,p�JU���pZ�@�RW����#�;-
&��!� Pl��j~6���r���0\i��ר}���?�Pc�l��p�
R�XZ��5F��<نNށT�4��u�@�Yl��蠃�k��9u*S9[S��'�6����2O��u�ݧ�����8	�������pK��{�a�;v���#�f�-ddJEpG�80h��/?dn��b��vF��ƹt��VFL�bkT�]�fM��˒-4�J���M|���$��J'�ڲgY;��e��Ӥ1������כ,~��Cn]�i�0Y"�蘊Ab��b�����Y��i'6����)O�c�_�l₁�G�%h0P���	|��S��_�Q��m���OD�ޤ�H��~Q���tn��x��8�p�V�Iz� w&]|hM���D�nSL�[�΀�?M����-��	�C���
F��&��c��ȈK�D�x�x	 kù*1�Q)#/�<Q@�!�p��;l��\2q+��1�	�'���K��i!TAp7H
�1�v�c�N���m���p���z3�F9S����q�k%RIxȊ*2�d��w�.A 3BJ����,S���'�(Q+v��7K�e2C�i�j�3�-�E��|CD��T>z�����t�K�2@�Ij�#�o�tO�5�G쓻(2�9KȤn*~A����1M��0D��%�����)y�-˦��yFAkg�/G���
j�Bҗ��w4X�b�>��<AF۫IB�sρ�@���Q�O}2�~0):�o!�r�KM'	.���ߴD
��)�탵Ș-g��q�'��K����"O,Q` �����z爽UF����� ����٪`z��kU$��Kh.�O��4�G��3���]C�4|���oIظZ�i���$ ?��A �oS�u��E�`a�Z�-�(�Rћ��}Q��!�/Q�EP@ˬW� �F|2��{����J;U��XQ��V���O��FB�;�j�*<��%LM�����w �%>��&h�8~
X!�IOU�	�Δ��@�I��$�)��
��)�'N���!�;=̦X�u,�dMnA���
I���K|j��D�;�0�;���*�.\IĀ_�<iP�Ex��h�K��6qx�"�ږ�M��ϑK~���f�/\A�D�J|·O��]���B1f��A^�Ct R�/+m$��ɒC5`���2Z)�e�ׂ��6r�#�	�%ϓ.>H�!���2��Ʉ�	�jL�L�%��>���
^����Ǘ-�9q�M�(E >��׫��G��e`Ql��?�6��n�ca��C�*̉CA@	��T�ȓ ������V�Xbl���9/���ȓiR=`Ŗ0��9� I�	��q� (�ᛯb����k��% ���2�`�`�I�mq����=m�B5�ȓx9�5[�L�40��	�&�[�:U6-�ȓc��=��¡+d�b���~e�ɄȓJ�T�AG��z<z�i6$�0G��	��U`\�2Q`@�H��e�5"�*e���ȓK
<�EN֊�����E��Te�a��P�0�����r/
@���nP	pd�8s��T�7]v]��S�? Z�JP���i��bO׮Ȕ��"OH�S	̜��]��.�9A����D"O,��*�f���C5���i�"ON5ڄ��*��p����^e�(ӳ"O*�kRI��$���N? f`$�"OX]�cЎ"�����[�"ք�b"O�Qs�I�+ER�KF�m&�y�B"O���� X086P�+��F|ڸ�$"OԹ�#ąw�d��l�Of���"O쐒�kD�+ZL����yF �C�"O~y��)
�V��1Bj�hK��b�"O��z��F ^�Q=NȀ�P"O�{�k��EPp	�3��*Q*>��"O����NZ#�$���b,>��"O,��C�	 \B�9W���\	ڸ�#"O�����ؓ)�R�@�m
ڬ���"O�F ��~`�����U�r�U"O�1fyk����e��ѩ��^�!��Mh�̈�GA�JT�I	ui�!��!��d�7�Ԇ{_�9�dgK!kR!��3�N��ㆫع�g�5$!�H� @m�3D�>%�Z@����	�!�ș5��U �.�m����K m�!������3I�^���q4
S3�!򄑉= Pi����a*�(�\�!��IL}���<ml^�+@�R�:!�$�6.��K���
I���ńB�Y�!�MSf�Y'ΏR��`F�%K�!�Dɤ
K�8��d��!㄀��k�-Qv!��6r�A� 
5��ғ`
�f~!���/\V�K��S4�2���Н|�!�dЁ�29������9��K	��c��&��
�5B�A��@���3õ>Y���O��jWAӱ����fD��P:���Ԏ������<�����. �d�ы>}0x ����۲�'������?�WM���Y���ԟ@�X���or�T�#G�;.r��3.�����'8 �y��W��Ov�'d88�Ze�r.x�0	�"��I�S��{у�!XI�o.�矌ap�	�j���נdiȄ�ql���0�V>�z	B��>��M�|�w�E�Hr2Ŋ!���@��uA�h�x�X��4�c��O�?�3Q�ފC��!#�	\ޜ�s�ź�0��9��%���p$l��|�Pà�'\���a���	�O���#�p {��ĢXE�j[4+���Ě>��g�6hW�9�xJ|j�'���1ҏ[,	�J�2�K�y_�E��O`MxD
թ^k���|n:�ӈ<�b�I���y�a���]@7�,=�01�>	�'i�*}(e��!�&�0��|�a���RwŤO6ʬ��O����\#����bР���H�8�<���y�hU78�>��=%>�R�՝M��t��S<��pw/0�$I&x38)�{*���(쀥&�Zc�UB�V�6��'�����RJ�S�Ow�D9A�K����Ӯ��[u}��4(&jq�3�1�)�'T>���f��E�<�3��'!IPK�c:Z`�'C���'05�9x��ٚx��b�/�N�8,	K<�զ��uPJ~�)�	U�w�ȩ�n�~��x9q���S��d�w�j�Sv�	���S�O���2���}�b�R-Q\����4S'ބ��o�Pˢ!��Oeh6�y��Z�+O��;G�./X2tٖHT.U��@Rp��0s�N���m�F��i�&
㞄�b���z�6̣����4h� �'�ܣ�K���O� �B�L�0"�����7u#���'ʆ+2���~�ͅ��$����Y� z����Pu@C�,{Htk��_`�<i�M�B����B�
�Ā��nD]�<i��F��\���b�x�}Ĉ�c�<��l�0\�rB�W���q2�	[�<Y����Z��U���-��5q`�S�<I���0p2�+Gf] �"��	�L�<�G��L����ղ["x"4��}�<�劌�|��1!͈50��X�FPw�<)fP4� ʰL��B�6 �$Yt�<� ���`'�)6ݱ"7���C�"O����h9zغ�9�!J30�`T�u"O�!����dn2EӃb6(�&��0"O�أG��i�l32�Jg�y��"O�(B���%X�=YƠݹx}*��"O\hkG�L�����Yl�A�"O,����2f�W*m3��Z3"O���0!ܛA��;���=5\x!S"O$�sRϐ�/��)F�̉):���"O��H�mJTqd0Bj�J�*Oi���A-����Ҥ�6�0��'�z8�@A>�:Yx%�[Z��
�'����p�6_�z����8f5
��	�'j��i#C^�"�$`	�'I�[����' �8��8}�� ʀ� d�a�'��˓/.er�����%�FS�<�R M�4��0���.��a��N�<)e��#C�<��Uj
<j���`�GJ�<�R)I�i�m����P��b��I�<�叙��q�"�5u�u��@~�<�Ӄ�I}n����%z`��Op�<1�ն�B�(����l�lȡBMp�<� $ p�8s�.B�r�NdᒅZU�<���]T�N����^�=��IMQ�<����u��A3���s��� IQ�<I�C�3m\ɂ!i�9*lpR�P�<�HW]�C�a�"���NJ�<���<}9kC��g�j��U~�<� /�9BIQ �?{7�5��ƕD�<��Ѝ>'8�p���T�9� �J�<YPP�ߺ�����7H�M�ȓ(P��UNW��z{P��F�^Q��9T�'L�'��z�C�	?�I�ȓ]�2��!B�MS	�����QMtl�RE�0j=�e�To�E��X�ȓV=��p���s�"�R�2���ȓqI�XZS��  &*aj׃ٓIj ��ȓ?p�1�Ń�%�2e��AD�]��{�� ��H֫`�4���FbBL��tuę�퉮Vg���D��

�d͇ȓ:whER�hY.~n6�`�M�b����5�r}q��6XS����F&r��ȓKa|���BF?@��*#�?�8؄��ne����-WԠz���?k�8D�ȓ6�a��D�L��!��.1Z ����ͪԙ!�	7zo,�I��߬Ax�%�ȓst ��D�t*^�����mTH��"��Z�MB�r��RQ(����ȇ�6h�i��#=�}뛎k�\��~�tb��D	-�5�@撥��ȓҰh37͓�x�
�CaU�����ȓhđ($�_3�QB��GE����JD��Y�&س������%�hd���l����]�j�b�k%ѕ/�N�ȓ����t$B�84��1"C͏.����; b�zA�S΄!�I}P܄��B�-�B@�*1���G��Gb�}�ȓl�	;�Nf�yL^��Gm�<9�]�^sR��&��%N�Ȩ�	�l�<)�H4N݆�8�` b���d�r�<yu�_������W2`��-�U�<YǊd����	ljX�� T�/SrB�	"2��RC�	:b7����ꑫ[�B��bu�s��G�N|jU	s��y��C�)� \|�C��&U|��SD�8ξ�"OXQ����C��0	��ǟ�t�#"Oh�uB�/��8��$5�
�÷"O�	�AN;G�r��hΫ?X���"O�Ĉ`@܁E����e�16"RA��"O� ��Y�ؽ�0N˪l�fy��"O8�S�
<��"� �L�hy��"OB*�'��dFJL��ʛ�O�b��"ONe�7��<0>>�g������b"O��ȒKU-�͑�e�:��"Oe���R�2����/�ei�"O�u��F��f���s���Z��+"O��*čƄ4�#`G�B���D"O���ɞ.>]���!�<A� ���"OP��q��bd�yz�@B:O����C"O( ��Ǔ�0�<S1������3"O�@�&���c���_��u �"OV��H��4'@A�`d
�ܾTA�"O���r�[�N�2T��
����25"O��I�R��A���"Or�z�쁄o\�- ��*��� �"O�Y���f�M�c���9pА"Oب��IPWH]�ԃ�� 	�""O�X�Fa��S�d8y$#׷u�d%��"OZ� D��)v�֕H�bP8pꤔ�R"O0ݹ��τX�h������K�"O���@�:��12�m� x��*"ODsŎG&?����w� ��Y
6"OJ��U�ȫV�X�t��24�6���"O��k���~V�1i�@!I��*�"OF8W�B�tMԙp"��
�j�[�"On��%��/J�YpnJ�����"O��9��)HRE�a������"O�d fl�/s���;#D#�J "O>�A���D�I�g��3�RUk"O��'J��ƀ�4������	�"O��;�)�"a�>�ym�[�����"O��[%D�.hV��k�>��q�"O �ф��.2��H�6�P�!�Pã"OJ����:������ZQڜ��"O��5eͯ1�j�1�m�$}A H�D"O���`�[#^�v�q���6;Q��R"Oέ���"F��R�F(D�rT"O�U[P�(�M��W1t��"O,T8��^?W��⑯�&!.��"O��;1j�P ��S�>1�L+"O�]��F�A��9���.��\��"O�ya��DN$q0j�Q �P"O���W�譛���2>�$��"O�8�#*�#l:�8&��֔J6"OĘ��!g<�Q��8�Q��"O�y�'�Y&��H��k߹h����c"O"��uj�aʙ�Ԥʡ$��|��"Ot����<L��0�D�I�f�j&"O"�kեߟ<�Z4 B��$�F���"O�*�e�v�%������I�"O"�y@��#R�@� `Ã �jј "OD��A ˵Tz�	�5%�c���be"O�T���@(9Kd���[�*!�ն���BbO#u���ʥ,C�s�!��[>1��0�ubU-�*)B!�R�&�!����B ��b�����*�2�� "O0�2�eC�'���УJ�&({���r"ON�����kK�'뜮ix,P�!"O� |X�G��~�-�sǏ�P`��p"O�qa`F�ec�T���ܗ�d�"OB`�a
Nk����L��l��C"OXyx�+�S!�ȃE�$�\�BU"O�|$ ۶ U�i�qgāpN��q"O��vbȼq�n���OJ#�ج"O�QH�L�+t$�D�'�vdC�"O��R�P�f%
"T�$W�(8�"O`��ƤR�Z�6�s8�)#�"O���@�p��&&{j-6"�kD!�.*�6��� 
-P���f*W�~8!��O^�8���n�ͻ`j�jP!�d��N�LbGl<|�8����hc!��&�T�r@OȳH�Z��R�ʥg�!���m��Ā���AR2�����"<{!���(W�U�4	�Y<�\��7?r!�ԻF���u��>e/�Mi%��BR!�D�w6���R{@8�y6$͡h�!�D/2*��gI�!"|{�K�N�!�D�q��TPҨ���jӂ(T	!���L�&�8��ӓf<���ԏc�!�"9�<�u�C�oh,�%��1�!��6��}��4u�Lh�7M&�!�$B/�(#�)�%��bTi.}!�d�e���㑏S���'h!�9(*}��ℎ+�6��0�=/S!�ċ�Lb1ZC��	
��	 �L�iO!���z�:���F�]�ؑ�7,�5HC!�F�X��81��B<	|^4����-!��,s�8q����zi�4;ቝ��!��u�H���d��{����h7�!�$0K�\֍Ky��A���#!�dT�A�%��t��K��n�!��<�쌓��C'P�Z<z�A�;�!򄝝f�����)�j�b���~�!�)� ���ӰA�$�ȆK*S�!�ٳu����@R�Qs��K�J�F?!��ӑsH�q�C _XI)�N=-:!���9xU6ݣ��y~V�ZBmX&u0!�d	�X��H��R=R|�T;��
�D!�$�|`L�*h��H=0�r�lM2:!���m 0���]�4�Ċ	�p�!�$͜|
2�2a��sb�,kh�6�!�K��A����OH�ܺ歇�w�!��z�l<�CSGa~��*�)P�!�$�5.�j����@n�P��2T!�DN����f�P��(3�&�!�U!aRx{,��k��HP�*0 !�->�L��&B�t�K�)�r!�F�s���q�����X!�DE!?.�{�ҵ	MZ(U�ɟr�!�� b�ucE��#LE�1Y0a��u!���AH�`i#gR�V�7�	:	t!�Dʈ{���eL�m��a��#N�jr!�䙿"�$�������Ë)`!���q�3� E�ے]���^5[!�Dָ!�4��ᙈ`zRH�����D!�� @��	�DcE�)Rrh���3fS!�DM�5爥��A��:PUc�㎲,O!�Z��F%�7!Z����@�-�!���:� ����:=�|����^�!�D�b �  ��   �  �  �     ,  �6  cA  �K  AV  y_  �i  �u  �|  N�  �  _�  ��  �  '�  k�  ��  �  7�  x�  ��  �  D�  ��  ��  _�  ��  ��  @  � �  + �2 69 x? �C  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��	h}�LO��dFug�	E�-�y"�_�9MN��փP�A��F0�y�SJ��|@@*f���� N�y�bO>1�$���Y������yϥ�n��,[)H4S���y��v*"U`3��'C����al��y��հe^����ǿ9&X����yB������0� ��Ѵ�y��̠^��=14'@%�>����^��yr���:�$0S���5*@ū1`��y�o˹g��S4DLa�9��S��yb�\S��!������KdW��y��M��j'�Y������bR��y� 
�N���Z����gZ��y"Ζ�=���	p@ٖ
K*��`�,�y"�I��R���F_|�PH0�¼�y��^�`Y,���G��fL�TaH9�yb���\q:T��H�	��i4Ɓ�y�*�)`6���2Q�i�5�yR��: ZD�I*M����=�y��+T�P�
�@�#L�u��I�y"�P6C�������*㺠�ƅ��y�G�#>^p�ȕ6b�B�������y��Y>NSh�!㎬m�DM��^�y��%	M��6L�m�����EȺ�y�k�I���j�F%h�Ny�%e���y�L�`��;��N�(ޠPz�Ն�Py"�^�p��x*��Z�"$�֮SS�<�#c՛o/�=K6/ߏ�y�A�I�<)$OA>a�d�(��z+�sϑG�<� ��u��7L�Jɱ�!����"O�0a�&�`��{�!ܭR�\��"O���A��=#�,�Rd`Ө~��y�G�'��K�jH�A�K"0h"�c`���/t��ȓI�� S�
��]��cD ]�9��Ix�'v���E蕬p�Z���/r#&=��'�~5��&ȦJ�]
��#[{���'�J��C���>��FӵSf<���'�
�i���=�؃�ǀK�V���'_V��u�ǒ@�d����)6�l��'u"��"�p�h5iP* �=�Oܥ����$�"}����::�n�h`N'��ҖmI_�<Y�&��4H1��8yA���F K^̓��=Y��!J�9�&$Q�,l�!jC!�U�<a���1Kc���X��5�a��}�<�a)ˡ���V�m���X� �S8��'�"U����콓7�Ä-BX�æO%D����Gh���4��3F"l!��(D��A,�t���y�i�b/�@��f"D���s�y����Q��,k�x���>D���W�dN��9BE�9���� >D�@��C�8�><�FL^&f����7D�h�L@�FlP2![� �K��1�I� ���)�q�Q��~6����(޲C䉼`d��	��RG�ۂ��&F���w}ҒxR���>���ܦc�Є�N]�I=��X��;D����
#l	����_��q f;D���,��6�EA�Kg�t��"	;�In���D^����K�$��eȦZ |�21`d#8D��Zg���p � p��	-,����1���\(�6h@&W`�v�T:USt"O�!��$W�?8�is�ȏKD��#.4����>gl�Aa%\&dйp�'ړ�0|�A�I:;k������BN$4j�v�ɢ��F�'|��2FY$iR�Mjǋԋ	������hO>y�+z,,:�$�i���4'�T����?E��1��M�����;=�$Dx��z��D�,|��V@͎�"�УK�M��~"�'��v �#&A���.g�#V��y���+����(���J��2���hO���D��y���8[�f!١	W)�u��A'�yr�W�;�lY��7��I��I���~�<OJb��}R��><)��t)K`r��!���t�<��(\�`bpucGF���Bg��ǟ����'y�'����#M8�y�mϔEl@5���G�<B�8t�T�`�!bH@h.j3d�{"Oڈ�H��D�l���N�2%���I�<a���\�P>,��ʽx��2�a��1瑞���I3R�� ��C9�0�Ӏ�9f�OF�'��?}*q�z� �eʊ6VbȌ�F-7D�`"t#�� �Z#��7.K�ī�*6ғ��D�>�I>q�-F�Bs��9��I���)���A�<�G�#O�����I	�SY��H�NNd�<q�F/27r�`�n
��P'i�Z��$�'����y����`l��aE8�j�'Zў�}�(��J|�!�:[t0���Sx�<�!g�TWd��D�;6�� ���p�	��0>Y�L�y�@QQ���hv���c'�<����4@����o=h�P�"8�.B��3i���)�s�j!z5�T�]R0b�,��	�C��tK���,l����ҵ(B�	���;����AFQp�̢D�Rŉ/�>��铊=��S�kM�<�@(���PC�I�{����l�"-}���4��3Wm:��?a
�S�? @u!��ypl	�2��/+tT$#��'ў"~�ק�$h�Eh�0N��sŌ��y��G�]�[��Z7�6AR�nЛ�~�	~�TӨP)�ʈ�a�V���WLч�U�R�0&�:M?��Q�
�.�`�'�$F{���%�d��!�1z��#��ׂ�hOh��	�$��Ͱ&��5ؤ�`F���铇y���5g��q��|��#\	j���u�jc��ק���
�U�t���
)�N%��NS>6����(�|Z�N�_|"%�G:�j�r�I9W���<��Q�mr� ݷ(߸1�Ej	-]n�̆�	O�w�Py���`���ݓr�0��'{�~�n� ,Uq��@�Px�A�N&���s~r�>��؟,�'�~�@�"F@�T��;j�e�A˂���ɱ�p>���U����.S�(��_��x͓�n�[���e^P`2#��(�����M����M9
p��쑤OofD� �ן��<��O�=Y�G�8�h�8�ǝ�A�^��!���O��]�O�6�R�V���F]/K�L��}�ϒlx��iVꖻ[������%e����D<�O�牗R�l�QV���6�����ʜT����	�>��� K�r�~��6���s�B��ş�(BY�`��4�@��0rM� �#m#D�cVh�x��d�!d�V$����L�'�1O�>q�񁁍{��0 66Ln9�##D��*B�Ж���H7-Œ��E������0>1eoC�kQN,����0X<���{�<Q��:OV��fƟ>��P�h�w���=��`H
Q���Qk�3k��"���Z�<Y��7EQ�Z3�H�;���$��X�<	��3�(ꅏ�� ��i���h�<�e��@qT�;_5 �M��$b�<�R	�%�6!�C�p�tAƋ�`�<I$��C�|�z�e��\��Y�Ch�T�<���1< ����W�|	I��O�<�W�P��)�1�b��w�Gt�<��D��� ��ܠ"��ŘӃLI�<��h��$����,��P�=��gJP�<���N�dQ��#EC�-:�m!�]L�<�T��~��۷�&�0 (K�<i��bm�����,.��Ѵ��E�<y�d�s
z�y���L����U*MC�<�#.�#eB(��jΟw���tJg�<	�c�[����)C�^Hcm�c�<���"+��1��˟o�4T!%Kt�<�a�<F�PY�bF����b �Wm�<Qbc_#e�^��OO�a+��Q�<9�n3Z��=�ĢկL�T:�RV�<Q䬙�/�rAcO�y��h�mX�<Rꊠ+�n��b��-D�2�[��R�<���,c�%���.bM�"-Tw�<Y���!Ju� q/�-B_��V�r�<a���&ED�	�''�����p�<�@����X�F&[�Q�wLB�<i���?��p�B�+R�,�HF%�}�<9�D��$��Y�юW)T��wn�<�d��tJ��	��C���)���h�<QF�q�q�pӜ�5�Ci�<��)9���R)ӱZ�����ʁ|�<���Y%����"�9}\��k�#T��K�,��M�6d�G�H�"�) !�=D��*�l��$i�4_v�	/D�@sR��``>Q�6��+��4��.D���d���ضI֧haFT6�y
� r*Պ@49�f�x�M#��e��"Or䳦�'VP�" /�1&S�x�"O�ً���&<ݾ��A�Ĉ$߲E��"O"�c�8L���C��*X�*qA#"O~�eK;/t��W�K�b�0A�c�'��'�������'+"�'���'�>�9�,��#�H(X�h�8Rz6	bu�'���'��'���'���'��'����*�S����ν|{vp���'�B�'12�'��'L"�'�'ּ��BJ�.��i�H!b5p���'Z��'���'���'O�']r�'wq@A�,���w�E"k�DY�W�'���'���'�"�'���'���'��qH�ዛ]�JE	L2@)��'hb�'���'H�'[��'�'F@�ԯ�_Hyt$<:@�<|B�'2�'"��'���'Kb�'0��#��1;�`�2j���4�UB�'(��'6��'�2�'��'���T0R�Z4NN�|T.M�6i@6{���'��'���'�R�'���'�,�e����䥖^�6�QF]" ��'Cr�'`R�'���'���'��	�?�ؔ.��D���ϼQF�.�?a���?���?i���?!��?���?$뗵7�bI'� �`-H"/5�?���?���?y���?���?�Ӽ�C䏣.q�̍@"����j��?���?����?����?A��#�f�'�N�Ri��I���f9���.G6?��˓�?Y,O1��	:�MC�J�X>`(X�Ht��m�n]��	�' 7�/�i>�	��M��F�k��# &���[�=EDHX�4�?�Uʄ��M��O��D��ktYzO?EI���=��st$Ĺ2�:pb$�7���t�'9�>���=GzarB�ÐK�:)0bV��M{��Bn���O�l6=�,h��0($�r��[�5���#�¦=�4�y�Q�b>�(n�Ʀ�ϓy���1b'xp�lx�(�'h��<�#vLB��Θt�p}���4���B�M����-C�8�Q���)]�<�H>1q�i�n]#�y�*��,�T� ��؆0�0�S��#��O���',V6�G����D¥_�B�3�iL�d��e�4'���I�ri���u���6m@b>a�Ո�1�'��\�q�F	DM0E��Mܞ1||ɑ[�0�'}��9Ot,�R��p�T�!a� �
$bh1Onl�9ud�c8�f�4����[AF� 5(�< 8�@�&?O>0mژ�M#�
t�t�4��đ<P7F`���8xNM���_�Ϟ�R�揖E(4���4��|�/O���D����",n`�O�O��m����tX�4$�	�<���d�ޢ\�ΰ�ŉ%�ACC,�<ڊ�.śVӢ��q���?���_mp]h%�� J8ЬrB�"_��l�vg��U���FD��Bf��>��]���	���d�?Z2R�iQ-������g(�t��<	+Ov�O�dn�8��I�u�kX�
e��["�׫;��I��MÉ��y�Ci��hlٟp
 ��JG�mXr�[2/��h�(S�z��Xl�<QP�ē'�XX"� ]<�,���?���M��}<J �!m�5X�+�cl4�I��D�'A�)�'	�)!懆�Ry�,�cK^�|�<���i�����O�(m�M�	�<|ҡ#4��=y��ܱ����n+�������ݦ5�޴�?�Ce�!�Ms�'����#%7s�4�����W�~��2ƀZ�h��3�ȱ���y�>i����Dy"�'}�ų�m��s���a��X2nx��'��'6��4P�1Ofʧu;Lp�W�5)��Ԉ()l`��'�T�Im��Bg���	J��?�r�#"��934J��G	D��a�!!���4 �(@���"R)A<�u��4�D��p9�1un� j�n�ЏE�*�����On���O&�4�UʂA�O�81�ލ�ܘ��Eu�8��lÛlA�UR�'_��bӐ�O���G}@}Ӵ��NN/U�,]�-�,���r�����ݴL�r���4�y"�i���p���m^.���>	gÐ!�R�
�JY��Y1�ܭ�y�]�t�	���I�����ȟ��Oݨ5�Td�2����I��8w�|�:�2��O ��O����̦睱v(LH@��A�����K��B�`޴i(�L�O���|����j4�ȅ�Ms�'���k�ʓ,Q��F�3^�Dr޴}�y2�`��2 R�SF�r���P���ef ��C��;k� ��窝S����W-<Ų1A '�� ��Qj 4�T*'J�pl�� $׹0I&� a�<a�fC�^��8ـCE�I�ֵRk^Q{T	�o��,|$�E�X /�� d�oQJ�D�˲6X��H�Hq��#�1z�V����̞ojxX���S)�IC��ƨ&{漙g�d���g�>[��:b�$@_�M��-]�z�tdӆ���W� ���S	Q�&YJ��H�ٴ�?!��K�p��c�̙ZPD�Ty���iR�|R]��$g9�jf��:�D�7ɲ%PFf�{, 6m�O���<٥�6Gś�_>����?�X�WZmb������ٓv/9]�7ͪ<���?���M�O_��4@8������
)���$��-'r�o�ryRȇ�j7�y���'����6?YD
�p��t�'��0R��=ɇc�����I۟x3��_vyʟ��x�o59���R��ٻ-��4ѡKA��M���	�V�'L��'��dO!�4�<�ᕪR�|��ׅ7x�� �q���)��H�Oyr�'lr�Ϙ''���A|r�p�%ʸ$�@�CW!n/(7��O���OFA)0��e�i>��I�ȥOɱc�.b!��c{�P��T���D�O��d9s�1O��$�OB���q�? \�s�i���=��J��R|P��i/� �P����O�˓�?��a�^`�Tf��v�Y�U�Zt�'S����'���'�"�'��\�L��B
�Z��bM�,W�.m� d��"?4d��Ot˓�?Q,Ov�D�Ot�d�s0p�M�;�R��� ��5C$5��4O��d�O��d�O���<� c=�Ƀ�1�8����!/�f�p��ϑ���V���IOy��'���'f�h�'b.��r��{�6�QEGܶ	�щ�fg�,��@U����O��Ch�^?��i�1 0�B'N�t����N�d$�m��f���D�<)���?���o4�5̓��i�x���!�(i�1�sn_�?�Ei�4�?y����bm̀W?�	� �
9.���N\�}�IH@��m���I�O(�d�O���	��$�|����E�k�`b%㒲s7peLN�M�+OE�u����	ܟd���?�O��ϰ.�mkDg�x� ��!uʛ��'�r��y��'^�IF�';W�2��F�AE+܄|z��n�Gf�\�۴�?I���?���Wp�Ixy+�<(nIpbA \���1<kL7�ؑ?���O�˓��OR�c�-Rd,��G��J��7M�O����O`1�7�b}b\�D��U?I@�5�H,S�ǋ<���t$Ԧ��IIy�ʜ��yʟ����O��d,6��9�#-�.0��k Ö�[ض�l���t
��G��M����?���?��^?I��q�Bm�@8kS��B�aX�bĆ1�'v�T(�'��'�2�'0r\�tk�,��* �d�R^}h󁘁QN����OXʓ�?�-OZ���O���	���У&[�4��	Ęh�5Z�?O����O2��O\���O���K�Fg^8n�:s*�2���3In�PTڬ@��=Yܴ�?1���?��?�-O��N&e��i������a8څp�f�16�5S�4�?��?�f���[��%k۴�?9�0�$$"p�<q4e�P�^ VCr-Ӣ�ie��'2U���I&��՟`��0)���o���j�C{�дl���Uy�b�"vp�'�?Y���B��ШW���1Q��_y>�(f �;0��ɟ��	���n|���	oy2֟��Z�	_Fx<a�f�,B̲�`��i���'I����yӤ�D�O
���B�i�O�d�Īa(L����˝s;Jt;�bMg}r�'nZy�B�'cr�'�41��O$���2�ϋ���b��P�KΈ�n�K��
�4�?i��?Y�'�����?)�%����f׭$�ms0�Q��^�o�i�x I��'RQ��R�ܟ\R�� vӐ���L��*O�]�gN� �M����?�����۳�i2�'k��'kZwp�4c�.ي_J�9�G�]����4�?Q)O��C0=O��ޟ$��֟0c�BJ�|>��@m��x���2 &��MK�)�S%�i�"�'`2�'��맞~�" �\p#���xf��R A���$˽�yRZ�d��ȟ$�	iy�Y�g]phڰ���5�z�I�Rz�Vj'��O6��6���O4�$�]4����`��)c�9i��7Od��?q��?�)Ov�kP�L�|Zs�7
*��  G��2�A�FIO�I֟ $�P�	֟쫁*l���6��>c�R���#ݨ/�:�H�������O���O�˓���[��Ϙ�^7>9�¨_�!b������u��6��O8�O����O�)i�0OV�'�`Q���Q�|�,�A��v���޴�?�����$�o���$>	�I�?�1�<29J<�$�%�XH�E���ē�?�� �,̊������D�,SX�|�Nvhke� #�M�-Ox�K� �릅���2�꟢��'`��.S�H
��f<����4�?!��c'p����S�~���r�F�p8�AE���It��lZ?8�~�3ش�?����?��'�'�Z<��a�2H%@IҠ�[;B����1�ik^h�'ɧ�z�Āo�J�I@�V�<3�h�AE_t� n�Ο��	ݟX�tIݮ���?����~��W�gM�Ţ��
eD� )X �M�L>�Ɨ�<�OkB�'B陔c�I�a�4'^J�;���y�6��Ot�jĔI�؟l��m�i�%
��E}��I�)�:ܠ}��'�>����<�.O����O���<) �.WF�QS�X
a4�����ţ� ݒF�xr�'\"�|b�']b%ڈv�V	j��<Ep>P+&��e�\=��'|��p�����'���"֣u>����դmɄm9G��9#�"�I �1��O��O����O�ъd3O\���g�1Q�4���l��9����o�`}��'Y�'R�!. �M�K|za�cn�y��� +8ObL���/A��f�'��'�r:Ot(&�'�E؍���՜q��P҇�T�PZ��m��l��^y��%@�@�d����r %Ղ���R�&��XP��`a�	쟴�	(JZ���~"dK�4���R���&�jH�f��Ħ��'���)z�I�O���Od��#�ʘ�D1bsr%��S)5R�oٟl���K˄u��jy��I�K�~�J�Vn8r0+X����$P�6��O���O��	�Z�I�@2�#M:��8T��j�`D�'�M;���<K>E���',4�h��w���D�Lm�8u�tӢ���O��$��<�^�&���	ԟ���lI�2B�$[�bu@�O��@��>AbKI�}m*��oD��� +�H������^�\sJtK��@X�v`��Ȍ5��it$B�B�R4 ���w�~8�CΓ�h��R֌L��~� K�AJ�H�r�I�{�(ay�dZ�p=1 �-H]R1�ǒ *����+Tv��T��&���5�D�Xi���4W��m�6T�6	���!@^����
�������p��e2Oǧ�q���D�H���`�Y-i���A+�R&0����R��r�M­�J�ۂI(f^n��s�'[��� *�02(۠��@YS� E��a��O����q��OH�1%�@�� �͚w��6͊�/,�����X9(e�� �!N�y�N����fE?ʓO9,���b��+� x�� 
$�E�����X��"L;@� ��TdV�h�
q�#��8H����ēy'@�"����ےT��(�;�>��>�l�&IF�'�Ĵ��d��c!0�Gx�i>��42��"��B�"A��ѫI	C��0+K>�1jPD����'>�W>阷�۟��U!颽;���B�"�3��۟0��?fd����S��O��pGN 0,����_8�b��U�>�ѫ�p�2E�$X�[c, ���);^���AiKz �e�E��)(���	��S��SZ(�xCյ7��q&!V8�\��Lh(�3�/
��X"�@7v��I"�HO�P��j�A��TX�B��9yPa��%��)�I՟��ɷf�:\��柤����<�i�YK���Zf�$�ص��!sg�Wq0��fg�xR`��^�2v
]�|�R�R��	�P��]��\$F*\����e�:�j��	���[�b ��=`��7�Sw����3=Oq(�G[������i��
{�:c��O��(���i>qG{Bj��8�8�k ���@����#�˛�yb@;~�poN�-��I��h�����c�����'��	�H�I@�M�4������Gߊ����O%cN�����P�	ݟ�I\w���'4�I19xl[�!_�9z@��a"NB�AB��Bq>U��!�t���I+P��Z��d��Oh� 3C��LUb����*+��H�T@\�9�2��!���zq�!��"�����Oǌ*�zpD�v(`���'����g��m��b"#L+ri�m��k����"O����JdC\����	��+��$���Y�	yy��9&���?YE�RFT~@+@��+@����?����F�1��?�O��Bb�&V%h���Q��i�Dd�� *0���=V������о{0�{�āx�'�X�`+�a���� �ܾk|8�Bn����v'��!D��=����ᡅ8Iᔣ<�$NYǟD�	GyB¶�F�a��]?T���F���'9�{�l�7-gZo�H�ҠP*T��(:�'56-Ē&\*���NrP���s�"�@���<!��ܿ=���'?2V>	B�A�ʟ�8�� =I+M�M/V%��J+|+2�'����d�ly��eU��>�(��]�}[����Z>����=�����R�u\��o*}��Ѿj��˶a�,��u0�d_j<�+&hp��Vp�6��p�ئD9�e�h����ɰO�z�$[L�)�SMt`I�N�F����稟�\�pC�Ia���y`-��"�J�]�d��D|�'���+��o��� �0!��%��.jӂ��O0�DM$;��X�O(���O��4��թ��(w�Nhr����pD>ԫ�Cӄ�<8{�+iq駉�$8Q�S�)�#{����'1
E
�nߣw ��p�)�5�֍��e\,V�*�{� ��&9�I�8��O�P`����<a�Y�W/V�
���/f$�*U�M�'a,�"�S�g�Ig4�q* a,�qaF�<�B��(J���ٷ��g��](Qʏ.���r1���E�ɪ��̸���r1�1�œ=oV�0��&q�u��ן��	ן��[w�R�'��	CW(�B�OÁQ%ە�+U��w��) ޜ�yM�jL�T)Q�J3(%s��d�)��5Q���,Z� �*4C˺!Ɛ�C��Pa��]�vn]�uVR�a���ډ`��D�	VP����ЂKB�5��#��r c��'���B�Mu x�֬�P�FG�A�!��F�ap�ƷĂ�R7⃭�1O|@�>�����Q�F�']��N�&0�B��_�����a�/g��'ݶD���'�>��5#�k��f��pfӴS�"��!�C_���a���(�VիeE]������(Oq������Cfm*�Pugp$r�#ɷW,JQ{�h��f��(c'�9�(O����'��'܀L$�̚H�X` 3zG"�`�'�DT���n�D�g�$lr���'d�7m��]�AC�N&t�n�ɐ�ӦV�t�OpKaK�����,�O���[e�'��p"S�T�hR5h�_�m���'R@���v�Ĩܞ?�Ѓ���[��x�d�O%K��x82H�r���������I�(�����锌Z>h�'�8 >�sE��W�����kE�t�ZMp��4}Ri�
�?)��h�����"GL�rǞ*&b�B�'CD��B㉉W�<q��i�axxi{E(H�1�6��d�C�'�`IS.��b�4�"�� �^  (v�����O���	):~Z����O����O��4���Q�_P!F&��5N�ĩ��.�I7""��d��A0�!L|T"�2���B_qO��3 �'���g��5c�w-�I�� �*���O�Y�����J?v�7KGw_�ѻQ�Ŵ��<��\D}��KG�$}��33A���'�#=E�DΟ�Gd|�
á��/�B��	�lI�2�'��'w~֝şl���|b֊=� B�[�@�*,)X���mơu�6 K�/����c�$	4���M�s���#��	����NN.4p��ӑ.��L�0L�!p��A7FNW��������9�̼{��	�E��
�K�)E���F��=�����g�O ����J�Er�ϔ61�����Gܕb���?�])Lv��@\�[Vͣs�G�k1O�0lO�ɄJ���i�4�?i��\�*�,C�� x9�#�5.�6�I���?�uK��zl�՟$�'Ev:M�IS�	 �iz3̕�wT�I���+o-���+aB�O��
wK�L�|mQ��V0y��aiR�'8���W��'NI��hV/?�`!�Th�p����	�'j��q��*� ���#c��d��'�6�ِc�bY�V�7���jg@P	�1On��C%Ҧ���ܕO>z �w�'�U�w�Z�Y�4�WR�w�>C��'wү[:M���T>�g0G�K�X�lԣ�A�?U�O�e��)�S,0�q�Q�D��9��%*��'����1=ɧ�OV���eꃷ=_Tp0����5iЕ;�'��T��K�SǈAH�W6�Bт
Ó ���hڦ,�<9|+�I\�:OzLhW�Tҟ �	��8��1Ze^�Y�^�0�I�\�i�1;�AP�-��9�oۊw�t JF��PYs�׍}�8����1d8"��p�9�I�(SY�%ۓ:O��#��#t�`Q��<Fx�R��W:�A%J#����S��=[�q�8X���S��y"��n�Ay�.S�U�|���,uZ2(x����ԯ}~���Y���	*�v��%�î^��`���
�p��̟���I����uD�i�X��"F�; <���4aٴK���|��O���V�H��8;3ĵ�#E#)��	�N=w$��J��ȟ��Iџ��	��u��'�R2�z��F�y�
T�T\99l�B�ۜ0�fH�mL�n�Y�@`��~�zu �KK��(OxՋ�6)�:hhr�J2 ��S��B�Pd�h��[j�B!��'u�eP'�-�(O^Ԓ�CU3Rz�R���2�%ssh�=b�g�0�o�M�G���~u���S轀���4�\���'��'�2�BqjE >� 2H:4� � �y�Au��d�<	�É��&�'���;Mh,��,\r��"KQM��'�Q��'���'i�����72�1�NQC �{w�
�Q1, ��P?p�l�C��ݘ�b�V���(Of0`j^�Y��qr�(P�ּ;)_�h��cCcȹ`Y~ �`���%��+�(O|���'�D6m������^%f�P�cڲl2�����z'H��I̟D�I�|��N��I7��r���.+衒�'�?SH��Ihx�P�޴A���H�jW��*�#ã��̶�c�i��I5$*�5��4�?q����W�@n���x��EKP�&�v�� $wJ:�D�O$��훩s 2��� x���J��Ҟ=��&�|2&L��#�z�̆=.�D�+&'P��PM8Y���B�`�8C�4��e�$cQ����X�-&x��
	fuP�HL3J�����`�S��~�d�q�N��쁉��`����ȓ&�r�1Ԧ�*�� �*�@-Z��4��HFz�)�gk�$�1,��\O�ѹ�Y� 7-�O��$�O��kv�D9���$�O^��O��E�KzXP�"٬[���ܞc�t�Va{�l��͛�Zz���o�K�'94���o�*�
�2�|��A��'�r$H�,��c�~aPȃ�/��I8ck��T���W,���)��*mR�"�w�@���Z?Ɖ�c�+����H!���+���L>�t�H�>�`.̕(La�σ_�<�p-ʸ{:�J�aƒG�R�+����<��;摞�c�1�|��S���W��������1�4��ٶ����ԟ��Iן��[wy��'K�I� R_
XZg����VI;��F�6��M6d�((�1�i't��ϖ�/ v�e剐l�ܳ�%8�-����M%��0v��=hSns��;�ș�$ڐW����E�-�`�%���E㝝'6�� �߳g���Bt�����O؟�h��$���&t�����(�0>�K>�S�[�L� �CH:m.�HP��^��B�i�'VeZ�z����O�Px�胳D!��HwO�W^�ё�`�O���Y���OV�S"sMB!�6퇗G
~��bϞ�^m1j\2�Re���8BvMHt��M�'���k����S�X�F��OX(T{��	�Y���X<X�0�`�lW'�џ`(gE�O��&��y�T�#��p��DX�D��M��(%D��ǯ��]�8��E	���q�`!��B�4q����a��a�)Kp�[JΰɻI>�����Aϛ��'��X>��%�ϟHA\=l�nկW�ja��F֟T��5r�������KKLݨ� X�[��z��2ʧ�xp
qGY�k5�c��'2d�O�H�$� 6!��h$'�^q0�a++�#��A����!D�؊���O���'D�(����ɧ�O�<EHcIwVx��؁%�D�9	�'4�����2�B��c��C��s�w0���t-�OF^0�gJH-�:d�a�+�M���?1�uV
I;0�Q��?1���?��Ӽ�A�Y��Q���͒�!@_�vdl�6FUMƺ�b��k�M����D�,,��S�? ʥ���ѻ���p�@C&�1	�H���a�b섦8c�hH��\	�q��S"�I��yR�U:[�=#�'O'	�(H��(U.P�\�O&X������f�B���Nĩ@e�A��pTP�ȓD��TQu.�Iw� z�X�;�q�'m#=�'��L*���-�+9�!ꦭ��P(x�8va�����?����?iԽ����O��>_p�i�m� $Ƙ��qʅlJ��U��p�ȐC#i�(���P���@�'+Q
�CQ]��Y�&�K�ĸx�&U�"9̅�V��0XEr106�gџ�&P<��l㦮^Z&`�X5�ŷ�
��v؟��u!�66j���B<+�N�u�6D���	���X#�cA�^�$�K��5��M+O>!b��8C���'x���	v
�}�K�
$;�O�1W���'�X<��'��9��cS�E�bƤr��*G�&�FVr�}ꆎ�<~��r&�'O��D~r	^,F������	��j��"Yhb�Y�h 7b���HBvХ�f�*�E���	��ēZ�(D�tl׵8���t	�i�@Ą�{��t'L]���#�Ļ�,����6�ƃ`���ЉY�|T ���H"�'_�@4-|�P�D�OJ˧0�2PJ�J���0���<������՛f%Ġ���?I�.V�y�=5D�}�bLA��H��`QZaX ��iU/�,tmE���0�S/:3�\@�)�f��mT�8�&�="Ju!Х�l:�'a�z�Ѐܒ|휰"� �B�ꍤO�)a�'�P�O񟴖(XT�%P[*+g���y�E�G��r4��)F(MA�M��0<�`�	�E7BE"��՘%�<�3��V�1m@�Sܴ�?����?���:&�ڔ����?Q��?ͻ"N!\h�Р�9{B����ݾ(\9��(��(h>I�D:Tg��"����	"n m� fjt��DP
��av��aK& x��&& ܵ0�kS+[E"�&B�S�'�L�Z�d�|S��#c���C�V9w� �pL���t�0�)�3��śz䆥x`��j��<H��:u
!�D�5\J�yDF@i���0����P�I?�HO�	-��6�P�J�F�Z�� ��;Ob����@��l���O&���Ox����?������O� Vb�������1uQK��]�`M�'n̐�c��x��1'M�db�EyRb͂F׼��G�A����ēCM�,���8KB^|)���W+�퀇��t�`9Fy���4(�	�Y�
��de���V`h��a�ыr80*����@��lRD�j)�ȓ9&�C�Ӭl�	` 
�T��q�<�i��'���j��F�$�Ot���EAn(`�����%���O4��D�Q�P���O��TI���	$�� ���]^yPp�7A��<+�8��)�2�܉��	�r8���A"4�ܜ�����|��e�|2�St�U�Jp�IX��N�M2�@��'^ r>�	'�H����Olo���ɟe����'Cam��CPB��i����	t�I��I]�x�ɪ2|}�F�]3dX8���L�k�L#<y��4��hn�;b{��K솦<-��`��"/@���\y�b�4)�6��OT�D�|��)�?���Ȍ4�1X#T3� ���皯�?I��mv�e0M�F���"ń,a���U?�O�A��1"��qq�ա �m�K�ؚ!@�bN�ۧ�M-"�ŲRg�'$y���CE���Y�#h_�uy��O8ճr�'��O��@�A��&hR�P5FU��^=�g"O�1�b/IaV�NH���9zw�'\�"=glK�r8����G����97)�vǛ��'�B�'
�q�EV�N+R�'U��y��ˆg �X�M��][4T�`�.	�b��J�t�3G1LA�c>�ORYp5o��a� `���V�g?rMAE�[n��M��t���*�3��W���*�-jnp�%J�,�p�%�l�%��Oq��'C��g��/Y� �r!�4�Jlj�')B�S��;� 3�n.�ެ��O��Gz���J��L붫��0]�ks.�[fs����C��$�O�d�O�H���?���$(��U�i�bLaB�i�۞+	�l�S[��4P��[�\ R��'!���@�n��hA*E;E����nC f����'�&ʔ F{��Q%H�>��@�� B�DD�Ԅcy2ɢ���?yKC�I"�`BG�#z��p�`�b�<�0n��8�J���O�J^ ��DlCc�5��O�%���u��֟�1⤎�C���J3GY�[���ss��i��C
g��':�	�e:lq�&�BX!4Eƍ:�� 2�K��N�<�Y�N�V��Ǔz������U]���� �1�щ.��G)8a�B���4]T�%O����'�|O ـ��	"�}�R���3��1�"Ox} �"SN��Q��9o}v�A�O��l���|�#�$��� I�� -�c�ܚĠO-�M����?�.�<ԸÏ�ON	G��+�>P	�Ƴ9���$��O����W����0�|�'NMpa��"u�VA�.L4~�(L�X��+.�S�g�? R�J`�_>^FD	�Fƫ�&l �>!R��͟��H>�r�/1�0�f֞7a�VZ�<i��ܷJ`B��Y�89$��bMy��	��D��8��h:���\��\*���:T�Z�lџ�����򦫘-+��	��I��1q1I�!tl�QAↈ"�X��<y �Nx�,�eAJv�"�2��U8�E��2�	�+����dО�0�~u �J"��%[�0�%��j"+�Oq��'�x @�n�$���]�P�dmQ�'P(���J
�]���+0k��F�����O^ Dz��	�&'2pZ�dB�L
���珴$�0�TaU�hM$���O����O.t���?�����^�$�6�� ��������^>{g�1h!�6>Z���J��X.=�ÓJhi�#*@��ms`��+� ���(�6R"3G�׭7[��`�Np���!L�Z��(AF�bӞ���eSZ���R؟ĸ�k�5T��j�T*F,?D�p��6�X��`k�>扦��'e8ZGIxӦ�d�ON���B��8B��ɵ
��%H��ڰd�O$�dO�q�����O��S.>T����5,�sB �w)j�:�
)Fn�e�	T�-X�tR	˓q���0�׳K{�H��7`~���b  �z8�͊�֙x4�����%O��hv�'	�O@<:�@O8T� ��?cJ�"OH��L^*�=ac)O*����#O�1m)6���K�KZ"i��B_��b��8q,���M{���?I*�:�����Ohؑ5�7���:7Fz�r�����O<�$>D���$�	�h�5�I	�niK$��M�p�'ZeFq��B
�"c��I�� 3O��`�OH�(��U�X��-�(���h7���Π͟��*g��j�<H!Ǘ=��	�R�>1�B��H>��4�Lׂ���U4j4饥
_�<��+�pn�r�疾o�N�p$�[��hO��~�'�
�@�喴H����t+���^ {��pӴ���O���7A�2A�B�O����O�4��V��0�v�;2�D�v�x�6�F8[��qT`�eh�W�g��#�v
��	>�Q�ݷZ��� (X�2����P)2�Z�`"�3���/+�Y��On�5��FB>Y΄m����I>7l�����?i��~
�r�GZZ�X컠F]-Z)��'�
{i��y��d�G'�3��b�O�XFz��Ou�[�4Т�E�O�q3Vʝ9YDZ��E'`��Rb�����	П4������O@���$Bm֍A�O�.<�jL�&.��{a(EGޘi�p�b��i����DAf)��I�e���3�N��m���S`Nş!:���c�d�8�/�'?�T,�A��2MR*Q2e�I�S�T	ٗ��<$���G�J$@�L��%E�OL�����]�IHy��'��O��1���)��[�k+}�X�s:|OʒO (S�OO�p|x��#*O�z\�AB�"�$�9q\ynYy2�݀f������d�I�����Hҍ7$f%Zr��4M@����l����I�|"Μ�'.�kq̀�},������i�S�ٹ���J�[�:3>٘�l�@�<AR��#:��u{�
_�a����30���C
T3j��]+#Ō�zb$�S��8˜�<���Y����	Jy���ŨqS�W�XM`��O�+ؘ'N�{b�	�5���F*�MeZ�*�'��O��=ͧd������5��iC��|����p�/D	�_�40��H��M��?Q(��I1�H�OlDa�
�8t�{d�ْ�U� ��O`�DU+p�P-�cgW�*?�6͑�F�p{�.J�$�O���p�M
X�`ݨW��8��PO��Ò)�]��b�I�+*.:p���7/�9(e���&����;[��E��Œn�j��t
��yp� �O�p��'��O񟔑	Ꮛ�.u���
oe�K�"O�iC��S5Q��:gL�_nB���->��|
�鉣 >��5)�2`h9�"E��!�R�4�?����?��^8�lj��?q���?�;R��)����;z���ϧHU��j��Ã@�vD���04�H
ăբҘOi$̫WeX�<�Ȉtr��p$��g.u�Ǉ�I��Lhr�8$P�ҵ���s|��dNņ'�=��4��y⃈nޥ�e�L��y�S	T�U�1�?���E�)�3��۪ �ě�`p��)p �:l!��!�v b�f[����bǌa��OH8Gz�OW�'j�����s�\��7�X��7��1�F��������!�u��'?�8�R�r�&V�O���v X8b�B�L��*bE;b�Lbҁ�f�:<O��Zp��*�t��fe �:��8l�*�D��`NU�_0F��CV9�$��1��"8���@{�ğH�Lœ����t����!A#D���|؟�jׅ��:Z,\��o8��Y�!/D��`�j� ZU8���b`����+.���MI>���=;���'~�E�1�*��b��e�5�#��#9 ��'���zv�'6��4���'��'4h02�)H�%Ɖ+�b��+L�ex��N��?Y5�?u{ܙ���� HM)��X8��Qg��O�$�� ��8W�V8�Ha�φ�?E���"O��yT��&������%9V�ÑO=n��r�8@�u'В#���a�F��v��c�|q4$L3�M���?Q(��dB���O�i�S�\�(����jZ���$�O������6F�
,(ٸS��9]L ���mk�ʧ\�>�Ӡc��pl�5�]�\����O�\�m�7�V)j��ԇoH�D���}��:˟�]�3�  �c�BK��ݲe�>y�ǐğ �M>��A�;�h�3���C�6�����v�<)]y�����=Rl�|���ܳA�F�=ͧM��x*#j����1O�S��	b,Z#�M���?��^��ߣ�?����?i�Ӽ3�ܞ
-40ӳ�^IԌ��'���'
<�
�kF�����]�b�HLr���gِ
����'!R40���f�g�Ɉ<��8�hL�:9�e���R�7�Hu�K>��R���>�O�Q0�ׅZ�d|C�ǣxe�`��"OܡJ7k	�{��aP�k�9I�y!���(8��4�t�O�	�bk
^�H���됯"-F�"- �Ȁ;��Ob��O�Hۺc��v��0�6��Eę�(gtA�^�
����lX���pC/*t���8
�^�#\,N%������D�Qr�U*WH��)�&D�TI�YfiIw�!�ւY�H�\K���
R��P��	5��@��nOu��ɩ&J>��#w�'��6��q��ʟL�In��|�p] �R.Z.֌ chŘQSx���Y��
բ���f&�f��6��ox�c�41�4�?q)OZ��6��ɦ��՟tp0c\�]�`Y(�)B�IjRM���Uԟ����X�*8�IƟ��'~��9�u��;`�����ј5Y,�!B':���8��۩,>��MӀ p��,'���89�?�! w��*sެ�Ð;0�YF�Z�>:�Q�HS�aT���<ʓ3|���	�ēgY�5H�퓿S�$@����{K�|��!2(��ѻk $SS��;�plDx�i>��4��a)�'oǶ�
D�#E��xI>!&IE�L؛V�'wr_>�h�" ɟ �$�لPsx�K ���!8@�����<'_�鉐Hݞ��nZ��2$#��K>5xb�K(�ziY�	B����s�R�􊲜>Y�aQ �h���W�-�q{2��#ai �̖�d?DM��'�=;��T20�VYZ � �h�'gȭ��cɧ�O�l]9���f�0 ŏ�S��Q`�'�00C$B
��X�a�9�.h*��i>�r��W�~ 9(ѡ��E#�m��L�V�l������� r��,�l��ß��Iğ�2X�� ��ƅ9pm��Id���f��9 3gJ�6�6#
K��O�Ꙃ����<�7�D�x�ny"���<���W�C�E��T��K���(�ˣY��2�tl	�O���P�0�>��1��C�&=2��5�!� 	@�-Es�I �(���|iބ..��a�F�2Bl���;�y`���G@�%{,|��	��yb�'��"=�'����e��BØ����hm2ٲD&]��8��?���?���X�D�O��Ӂr���17n��!�$`��4d@J�l��D�4]ya�l��|[# �z�T]�;�(Ox$6�.J�@��T��49*Ĭ�"�- �D3��7O
�ݒsf��(.}�t��¡���,��F���d��"LGbNԫ����z����e�5]����KΠr||��	f�)e�	�fX�d�hb���c��b����4�hO��![�eБ�J=t�X1U�B�I =l�a���t��0�BR�B�*	�BD�!LNS��er��ΨB�I8jR���H�< @i�?k�B�ɠ}d&���̓�=��[Yp�i
�'C�كci��3�����%N�2��l�	�'Wd��-@F�q���ӵri��s�'tʴh�+�H�E '��7h7\�{�'�"�{���9[ԡr�B�c���	�'��1h!�L3T5��X*`�	�'��	�`.̖-��Yt�@}��@�'�ht�S��k�������n�B���'���jc�]e4��b�ǍX�k	�'Lx�P�5�4jui�/'�0�#	�'(U�3ȝ�|��(Q��NVD���'] ��@+�cL8Q�ӥy!�'�T9R@J��F���s�˃6>�J���'�t���ȕ'd�*�HȽ�����'�\�"�i6�d̪F-5^p��'ʪ�z�@P>@h��BF�д�n�:�'��ī7�[	�bTȤ��[.1
��� D8�o��\���!#�����"O ظ��:��s���q^�Ts�"Ob��f��)>\�g���<Sp�jB"O�x���)3[ʝ��DV {6�ɣ�"O�}8��)SB�9S���g4���"O��*��R2[��pE�� �Yz"O@&��+�,h�V*�R��h��"O�9�&��b$�X@G�	��ʒ"OB�n�GF��ap�ϯ�ju�""O���*PS,�e��`�*��]�"OD��D�ؿpL�r`�!�T�s�'̐p۴~�t���O�(��H�s�f�ů��Xyz���"O��s���@[t���B׶4�x��NM�lk"Ν8μ#~
aD׶Zo���� �p=Pc5HW�<!bIގ>����.M/���Fb���'C�X}�HX��Zc?O7@ڧ]yj�q��A���f"O @�&�"�fH�gU��&<�D
�Q�2�)d��=�a|�'G �R]WO˗[�J=[�����<SG۷J<Y����y���kn"5x�B5y�-Ze���y�Ϩs�¹C�KY�g�p��,K��ēVOt�X'$I�x�z����ݓ�� �gëq�Dċ5
�"d�!�d	&o���)��zT�i��)y'��b�N�+!��۴r�FBn�֝K�$����λIT��TiŗM�����Pt���ɦ8N�� ��W�d�^��R�ԡ!+\ܩ����wRL���0?�W��x  [��r��dR�'�<��P)�4��LҺaH�HX3لhϖx��B"u�i�3��1ˀl��dɡwv�ؚ4k��*����V�xc��	3y���"�OV�c2�[=29�A'�&F�0�úi�f`�g�WG��%ۀȘ0�X��Cd��اy��:pb�����,aV\�2 ��1�y�a�a���3��%X��#)�:��\��M3:+⟘+�oT�kʰ�	�OB�E���3��qt�ڍh�� ��H(I�a}���ذ{B��z�P�D�<����媌0D���'�ԁ1�E9!P QG�9*轐����IF̤�C�4��AK�j�O;��x�U	�c�R���)O:;x�$P�b��Y��6��~2�ت�#W&�Q䎂��n`�#뛍*�r�#um�x؞<�!�:)4mJAY���q1�p�d|B#M���")I��c�&x���2�`��K�B�eB��9`�lL��"O�i��%�ۆ���j3R�0� �[�QD}2HQ�-��X�2+E*��n�&>���@���,�_$�}�O'W��h�E��D�Zph M�F�nM�0�.X�1OnL�4�.�H`��FR��h����2L�ł%vP��ǵܨO,��#�i1Xѡ���=|����v�ԫ�(�_P�9ja�E":z4�qLBݦ������J IW��yR!�ZJ�X�q�S��ҍ������ϓY�:��Ɉ0P�e��ʚY���G)�➬K��Т��ɑ�kMB׆ٚ�?�%*�O����$�K�ZI��6c<5e��k��|�ۓ#L��8"ū��X�(��G-W8�����.p	�W@<v�y0e<+T~y#�JC2	E~�ݣic�X���R�p�A �M33��5m*t�*�xZ�Jd�k�'��07��-�t�"�08�Z�J(OH��4�߁.� ���H��Y%�Ou3 N�x�A�4��
Y$RD���I�9,�+@�b�{�"*�4�'�R�BD��+�oϐ�?�޴¸'��0�VDc>�Zg��6$�n�hS��w�ƴj�ތ5��lA�F���>��b�g�n�`D�ژ�T� ���ݟ<rJ���E�׻{�T&?�~b�Ki� H6Ğ9
ȴ��R̧fa{B	�6�*����#Jx��f���$S�Ɛj&��hܠ
�֑iԥ=��~J���a��M�-����u�B�s�@*���?� X��R�{��1C�ĩKq�T5��n��O(��$
ƶ�F���@��V�,c����V#ê5p
��S �!�P qA�)�Q�h
�����[sC�+�țO�� ��e)J�u7���'p�h�O~�s�m�5=[�)�� <�B0�4��/M���n��6�R�`'1{؀ՌPX��9B���Y[���d�;�EnSY��B�Ќm�p��B�&Eѥ��3n�"�*!��an:Ջ�E�69rk� �����nL^؞�"��yY،�'�3wфX(!m�,gbVXsթO�(�� ��M���6�0�n���-l��aI��Ra�J�cBe֤_Lx| ��Y)ji���2�I����� ��~0����> �d�v��g�f�0�7��qԍS�`��a�@��s��õ&��5B�`��MD�@:��D�2{�4�B�OK5�i�3�Ѵ<C�(��@�D}�U��b��~L�7�?7�S���- �%�=B� P(ڳCD�Y�D0H�s�+D�i�L�5�DQ��X��X��'N�9���r1�W*T�}⧅���&^�yo��s3�gӸ̻DO
O��䉶��X&��Jµ��).� �=�#��!|6��>lk�=r�'|t���e��@y�O�K[�����|`tY��l(|�4�L!�a��H�!`H1��t�tZ<t�*-Cǂ�.r��Y؆��br�KY
c��S�!I�%<�O�lJi�O�\��&0$���FɆ ��+���;���)A)�t���v�Y!U�d�b?����H�RRa�E��(:��kr�^+Y��I$�$L/]2�!B��!9����B��B����!�'���g�H8�$�$M-9���"D��].����J��F��Ր���
�(�w;I�[5�C�V(ܝ�T���4���@i���p=ɡ�A�ya��o� ���b�ߦA���9Kj��3��1�@L�K
�=�>���/wV ����@��a*v��U�$��z`t�fn����=��	V�-f6hi�4lX��b�_$��E��I�w&�����
*���fGK��41�d�z��O>d��e�E�3Ǧ��3��(n@�i�Nܧ5rQAqc�;9�H�Y ��)|����ׂ���堆�~n�\mX�YugچXtxUcw�XUTXS�j��M����.d�Q ���(/"BL��ߖI9��Dx�	� r[�MpM����4��"0	"��̤ W�p�T ���M�F�Od6���j� P�aC;+L @R�_")�)I������髅�L��ЖƋ� 1X�	��'��@���*M�X��g�xR���4V��pY��9L�N(U1&0  �Q�6����Ӧ�.����SR��[dI�� ���<,��}��)2`�lQ��c4��2����M�v�Y����[<�kӌ�/�D6�OX��rE�	��E�2��x��	֛-E�5�1hRjd�p�����'�~��M��;��ր�?yO<��� �/vh�z�Do���,��v��]'��f�C�^ʐ�BU�#$���ډ�>��R���@�ɀ!W<2!J��#�e���R%D���C�|"J�v� ���.E+9�d���G #v�L���j�2x8��w%(M� ��Ŭ|-���D�"$��$�G�I�=���1)��-@N>q�)� �	L�z<����٦����$�y�-B\u�A���0��d�%-/lO�Pr���,1����K$&m~���7^��pq���mR�#R��Q�5�Ϩ������$˓.<V"��3[�8ì�/~L����
kd4�C�+5u�d���}BEM�`2��W0G����D���]�<���OH�j�ӓ$��gѸ�U�i�����H�=�Rt$$:5;����OlT�V!4�4���GSk�=p��V�Q�l@�B��~52��#���nr1�!�|uY�)˒ )Z�Ў�/v�r�9v�D�0ƢK��-Ee��`��'���h�̈́Z($I5�ZiyT$�P��l?ю���w��bp�1}:`���[8�I��'P6}	C��`i�1)��^�]IRLS�c��L�u&�
!=ВO�c�KVDC�#s�L�q.�*a���y�m1I(��Dƫ<�,a$�q�c���n�!3��%S� �3Y/���=�Dץc�A#��K7P��؁�V�//�. Z�ϓX�^�p(�tx�{���'>��j�-�nQ��(��\Z\��c�KH�VX�M�-�"��$���J_8��SŲ�B�pCe�6/�>��pBkӪ�Z��OR����'�Ni+��ɌG��A��,YK��/@&u��:t�>���$9@~�[��K*E�-�b��r��},�jaޡ�e����:Y1R�,��R��=�O�(�� �<����S�~Nl�	T�Ř^���W�'"�q޴ E^�{�-�= ��x��i�la��b�#\g���6�:y,dz��ɀ'hl`��j����2�9�d���`1��ڮd��MAEÎ�Mj`�';��	-{�5���x،x�ڴj��̓��$D�F0��kڠL�|�P���r%�f��(&^zL�፯_����G�T���O� S6	��y��A ���>��P	% �9��\=D�Ji�Ǥ�A�ӧu�y⭘4|����(B�[&rp���l^�H��h*�O�@ '����d 3�߱9沱�'$2R1O��<�g&+92�n�0% u��q�*�F�QQ��K�y�B a�h7-�!�<U@��3"�$��) �?֦]���I%D/nc�\���?�b�J��>"����|Γ d*s��>Ix�T+�+ReJ��hQF�I�lJ��i�'��0қ'�v���7�H�`A��N�R8�%�2d����Ċ*x�J�Ғ$ڰy�3,L\�0�]�l)*���!;6�i��4?QP4Ov�'�t4�YwY��'���p.�c�,����O�H�P0e0LO��[D��$z)�1\�x���Ƴo��J��O�v,`����]�u�OV���/�>�eȒ�&�	g�S1kp�}s�f+{�d��>����f��i@,��E�����Ez�	�]_��2�D\��h]�6�F0��b�\�2�VT���-c����&�I
i(� �
������X�3�T����R?@�Ψ"5c_:Xl�48˓zY��d��-"�L!;�g�����i��A�	$'`���O�20�k�$??.HQ�%h_�a��'��c��benKU9�<JLV�d%��RąM؞�(���
�1����6$z�􀧉�78D8a�_2�*��>��<�(glp�dG�����NΫt�6T�Q@�e,��[	��O�!�����=�T�W!	�����f�>y��J��Bq�ȁ89�,�ց7:j�EjM>�҉�M�Xw�B��A�P�\�O(�P��%{k����S�s���g�R*5YnY���>}�:9�%щ�?Q���[g��~r:O�O�5H�� D9�Z���ѬAR���UK�(�@���	^0̄剿*XLD�ը�	{�R�q�e� C4��޴(0�3eGK
|��䧈�>���NJW�tb�@BH��8�[��<��i�N��Xcl� 9:5i�:o����F�+��V�D�f�[!�5�S8��)�I����(��ԯ�Ƙ����0����b+�d�)1�J��䮁N'��*��V�-�z�����<n��'��gk>5��ᔟ�0�(O<��R�<:�X� Ȉ 0�t��,XU?ѕ]���I<�O���Fؒ հ}�P���t�\Dɳ'18~� 1G��p�8�K��U�|�2��o03Լ��$�BP��NX\��}�� �O,��d��չt�@/?k�T��$χ��0-��&����,�Q!�t>مȓ3�P%0F ��t��5���J	�@Y9WE"#��HSO�_˪u���uy���w}�|bf ��Ƒ�sN3�
��
�'���(��&_���.MK��q�4T��	�
84,���u� Јf��b�P	���5-��	�S
FEc6�5�O[$4OB� ��=J�csaV�(���p��~
�	�K3�D��
����@�<溱��J@�c
���97��PãB�rB$ ��OS�[$�y�ȓd���#�H	�4|�j5�Ջ"��ԅ�1�u�@C:T"������ȓi���I�*G\t�$i��X	�ȓHR���0cY����� ��$7�̆ȓWR�q�L]�!���$����ȓE�Pd�4aJ�'`-��K�R潅ȓU骳�	xm腺!ы򺡅ȓp�d��ՠ$�����?{�Ѕȓ"'����A����y�gֹ�p�ȓ%NB�h�-R�r���)L:)����<i"��'2���K�jTQ�T�ȓf����Q�����.N��ȓ��Q_Xe9���<�,ԈPC�p�<�a�v�� ����L-���n�p�<���Uג��h�Xpj��@eJC�I�2�Z�x���Q_��f)�'2C�ɹ	��9�!��)�0� �5�$C��$KE2�*�oڤ������ޢVbC䉢ut���+@�4�HɹT(�� D�C�6g���")j<eSWH�]�C�	�&���Vc��-w�8��C5!L@B�I�%#�L3�i@\���'M#H�C�	+[Ύ}:�ɁSlR�y�,ɰ'ͺC�I�fd,t�A��E:	��$S/v۔C�*M�J�ɡ-��$��K"PxC�	/	�P-�f�3s��;'�ٓ6<�C�� �����o����V,
,W<LB䉅MC ���B�-x#$isglZ�.3�B䉣p��bׁC�!������ZQfB�!>X�����> �"���!B�!�FB�	1w�tiC�fP�I��(#B�{l,B�	�`���q�X���ɜ�,�BB��$i�!�S$J.0� M��8�6B�	- ���EdU&p��H�%:D"B�	5UslٹD˕4X��D����6C�I�7�z� &.� 1�&�kc��I[�C�	�X-b�zGB���Jl�bԇw|�C�I��@�S�"R(����L!:�B�Z�BD@��#w�X;�`�=CHbB�	��(�b`�2<Ѝҵ�S�6B�	�6��#��%-�؀�ĿNC�	\�:B�D}�H��£iw�C�	4+��1�a�6-dA����#w��C�	,4��Q�%��]%0��=u�C�	3y{f4�6$ʶnB�h����n��C�Ɋ"S�ݻ2$B�X����g#~�pC�I�"^���D��:V�ч�U�3�RC䉏w ���H�Z�xhfnT	�@C�	7 T��C	�zN�PG��(�^C�I�c�T�֎ØkQPl���C�)� �T���M�k�t-y`���<;fUK�"O��)�i�(�~����-b�d "O�蕊D|�<\S���y�vq�2"O�|+�cE3K������)3�E"O�\R��M�=��#��`�S"O2�`�D�k@�Cti�H��P"O�QE�S�O����q��V�h��"O�8&�N����DI@9���B"O�|v��7lX<dqsg��I+�T;�"OjMB��\�ygۧw���`�"O�(ZDg�,ǘ��f��s��@(�"Op,!�b	a�I�S@[t�p��"Or�p@Y�~6~�rƮEi�[�"O�L��[�k���'��":<T�b"O�Qi�.6��ň��J}�"O�Ly���(#͊P��Ds����T"O6��`�9c`M2�eƬ2ݠq"��[�O~;���P�(��R�i����	�'����I�t=$x�t&��<�ܴ�hO?7��*漌������%�=vV&9��j><\P�����M���E����'��@����1\*}�iX{8<-��'QR騕o�7'p�h��Uu�&Ļ�'��8�1MD7q':���F�t��j�'�&)�B������q�ܴ	���'��d�-�j��<����*7�0R�'�xJ���>P�-�P������'�jS�a[�}�(7iĮea�'9N	2s�֛~H�8T�P\#�Lh
�'��H���H�\J����iR_Ҩ��'m1�ۓI+��C�+�-Q��'�� ���ȻYYP�!�ȇ	<�4�!�'a����h�9�%°�S�8���{	�'��9�'2��8� ��.-n�(	�'^�P1FH+h*�D"�nβz�'�yj�a !+��})J[�=|�t�
�'Q����U2gt�i���,8ʉQ�'XZ=jmL�n�xT{��ʠ+Ƭ`x�'_��*DMLк���g���'�𔘷E���l�T������'|�e�B�k�T�@$���_6�i�'GJy���>j��It�M�_L<�
�'#���P�_��bY��HˇYSfh�'���@,�b���'�A�CPvpQ�'�$t���	�S[�Q��� ;G�)�'�b����IRr�yv�<�LH�'����G�F��TzBA/ ��8c�'���E�gNNMpr�N)Jf�h�'"頒��&6�`���I�5 ��I�'�"ܪ/�3j���)�bO��Ǔ�HO4�&�Vq��[`n����T�"Oh�P�M
m�H��A �7B�,�)��O��=E��!� O�4�e�G.T6�@r��y����n8Ѓ��3���&�(O����T1eD>�"���b>��@�Y �!�Ď3F����%J���$kV�T��ɟ��?E�T�0E] �J0#��E��SUiC&�yM��WF��I�K� wnYZ4���yRCڥu".����rjГ+���?�06O���!G+qP�A����	E��!c"O��GQ�1P�=x��լ$ ��`�'�ў,��@6;��E�vi�Q���7D����"��k��B�4$���6o9D��ʳ�M=�ܹQ�[6�H�Q�7D��  ��S(�y���:t/H,W���g
�h�����F�&�� E��l�\8�n��y�%�̊e�P��|�����yҭY	,�����k��$"�IB2OG��y23=6jT)e�ev��B�]!�y��Vn�DRn	:U���d��~b�I]��uCE	%�������b4ba"a�Π�y���
0>��� ]4CG���u���y��&I��˔��s���)�\��y�ֹH؜�C��6Aq����y�f]�tE\�cgˢ`�z���I��y�C,������l�NL���܍�y" �5�$�p�F>��z�΋��~r�)�'4-�E�E��3r�^��5g
:�vلȓB@�����G�I�>$'�V�*���c��bK�)�.���%n�<�ēF�Թ��w�Ф�������i�"O�i����F@��a���Ra�a+e�'�ў���L�(lH�Ĩ�s�L5	��#D�Xc�N��r �;"�/U� ��"D�t�B)�i\M: AՑl���r� D���"���Y�Yő�Ilt:g
=D��Q1�B?Ny�q+���V���D�z�,Γ�ا��xԃ!N�!2����S���స:�"Ox(`1��qG�"C̟�(���b�"O�9��ʊ^�l��Lǅu0���
O�6ǖ4g�9�!�w�z��`^2L��'���2� ��v9����.@�d
p���8�'K����@9>�$* ��+<"���ո'��"}�'A
5�r��4jT�0Eܳp�)�J��D{�����	?5�o�BrN-�Q =�y�ړ]8��c��7bv�0Ue���'�铄HO��`:_F�isCŎ�3�0�hq"O\bU` 4%�,����--F\��"��E{��� Bi��ؖ �"R���$�8�!���<L�ړI�<�2J"�F�.�!��M�~Č]�ơ�1l���X!HA7!�D_d�0a"B�C�lPuE�!�䒬Iɺk� �' �ּ`� ūc�D$�Sܧ{Ǯ�IF_n��q@�5䨩
W��fA�C�&-8�@�

7)ҀHPJY8Y�"C�ɖ4�dM����,g���T�UE8C�	a�z%�B�
����P%9v��hOQ>պ��83ڡ�4��u����`<D�L�p�W��T��AB B��}�;D�`
cHS#N�$�Qw�e��8?ɍ����9O�azf)רe��q*4@��>��X�"O�� ���	�ڭ0�d&��S�Y������:�*��ϓ�SCl4�s剚`]`B�.3� 0Q�C�t٨���S�(X�'�ў�?U��d9���+p�]#)�P�q�.ʓ�hO�Ӟs�`]��J�^'��8�H,%���t��Ƀ}����灛S}4�$�W4.,��D��sC%��k>����G�47��[��1D�$�Ӈ�q��q�0 Ly*VYSs�/D�(1���=�"���"]�2���C,|O
�d<?	!eL������R�l�v�S�}�<�2EP(|�C��
��8M{�"Yx~2�)�';N0!!�!�Y
����-�0M�=�ۓ-0! 6#��2^���H_�i��'cў��������>�Cb,I9ĩbĞ�YC��
�h������
���c� i"B"<Q�'jў��ysl�
5hD#f'�]�ԙYddB�IK!z���K ����b5�C�)�  �fX�R�<PqE-L[�5�x�)��,c��kE���M"�{�IU:��B��(1��t۷�m�|���% 1~r���v����{R��-%bLxcKO,
��� +�y�h�=��%�
�:H��"Q����%������` *��T���&�)[��Q�"O*�QG
ĶS, �dN3�*��"Ob1C2�9δ��COE�SDz\X�"Ȏ�Ï�d'z�qS�`Z���"O(����CM��=��݊ �jYYF"O�8 Wυ�}�:xY�	�HyN��"O�,s5ĸ
������Q�Yq�"O ���s0����&ʾ`�`q "O�)5dΈ�H��t��&o����"O6H���	u(4���Î=3BQ��"O�X���ߏ,�YQ���j,�y��"Oz]jEhH�Y�ZUcfcϾb��)�f"O�9�M+V:4����E$|y�@�"O���&�
���@W���@5"O�a*b�R�v�`ф�ې��$Ȃ"Oh��
���]9w�U�$w:�B"Ohc�׮CeJA�P���i�rQ��"Op�K@��&>���PV�7kɆ8��"O2��˞�:�R�i��+O ��!"O��{���$y<ݓA��gD\M��"OZA(0�O+
�T�Ak
�^,��"O�ِeϠ�b�ٓ�W�b%n�K!"O�!�A@-MJjк�aN�7jA�"O85"�D��l����� nT"O��K �O�Sz��A0"� L�I�"O�Y��Qr�D�x�B/۠�`2"O��a��H<p���?�6}0"O:�#�D)��19��KhQ�q��"O*P:��))�XI�D��J.|�"O�����:$�^L�7D��6:T���"O(��W�?v��
�.1U�c"O����S&D��x�� �rG"O�=����<�4�wD�+]�!�"O�-����~ ��Z�ѱ��I�"O|�����6H�A���S�>���6"OP3�m�.b�Z�"�(-����a"O�鑶L�"}�E"c�4sw0��' zqZ2���T�D��e��:��'��t"J!H�n�Gd�,�����'Ɇ�aC�2� �[6
�&9��'��c�aڗ�@�򔨝4�y��'��@�� ��G���Ʉ��:~8�x�'.4�!�[t���4�P� ��)�'M��#�ǔ,�(�Ȏ��|��	�'i�Y!u.VӞ���,�p��'8���<��}���Z�*���'JH4��+a+��X�M ����'�d�6��:3x��{wk��7]�]�
�'�t��d^�p���)1G"z
�'�EC"�G<�tr�F,C��	�'���X�Ȓi��6�ͅ#f|1
�'���Pq#�5�@q)���G��x �'���îխ;�	b[�m4��	�'~:�S�
C�:��G�i�@���'� t���У&���3�"W>i����'m�
/ʙS��@����+�L��'xȘ�&̄0YĀy�C��BA��'zQ��Aʰ%,��Pס��7Ѹ�K�'�dc��TX���k��',yj ��� �i���2h��y;��P�s��|1�"O*岢d����"�Ծ|�����"O��䈞�
�0r��)JYr�"OB�0�K�7Qu	�|Pۥ"O�����5*ip ���K����E"Oz� F��q��K��] p�J4�"O@���Ӂo���X���3i:�"O����Z� UT/Nz���"O��'m�1z��ir��8Mȅ�'"O�z�!��_� ���֊'�`��g"O��S��F�<3r�7��ɰ�"OfXrjP.��i�F�,!'t��"OH���] ,�x����3J/���'"O�H��=7)��۳�*o-D4""Oa�wo�5Q+<IN8ႧG�)�y�l\Z���T�Z��Ӧ�݇�y"'ܗI,)2�(�EǴ-���0�y��&��4jQ�[>)T|Y�u���y2�fN��U��>8Q�\;eL�	�y�囝y��ڱ����FM�sm��y�a�'m4���H�~ژ�уd ��y��	$G�B��Yb*��!��I	�yB�HkBАr�
�ҝA�J�y""�9U�y�"+�"��S�nE��y2�г-D¡�#b�0>��J�É��y�!ܚ\�p[t��h���1vꃟ�y�#�=Z#�AxW-Q�[�&�ZgU��y҅���t�D�T<Pgv�;��A��y�n�	ר	�S��K�(�� ���y�J[��j)PA�.D*������y�ia�=[g%�<8�d�1a�J��yR�E�8���[5�?5��)ʰ�/�yba׿	XRpm5��m�����yr�F�FQT�(�\H�ّ����y���j��4��	�#\�PQ�K��yª	�^K:��
VPN�
/��y���n�0ij"鈹�X��b�y"_9|3Ь
C'&i�}�f�ک�y2�b"$�p�
)x�sW�#�y��X;
($�[�D/*02N��yf����CO	�)�ddjF�_�yb�N"wj~$�B.O1l�L��`A��y�A�e6$B7��cZ03AJI?�y"E��)�ظ�c��F/R͙�����yr��4|!���E�*����>�y�5T3��8��
	�$U��ś��y���s*�ɣ�MI�C�,S��y��ث ����E�@����)�'�yRn�{8�(�<�z	��E��y�B��b$�L�.�bE_.�yB�-�V#��,ev��)��y��щ}ղ�A6FW�z�=i�*��y�)9 fb|����l��3 �Ѓ�y2/�y@rz�U q�``��G��ybJ �@���jL(m��4�ed��yҬG�� u�
ƛmE(\H���y�+?+�)�V,�3�2� �g��yRn�	f�S�(�q��k���y�M�J^h$��i�0TȨÕ���y���4s楉�dV�y�����3�yb���6֑���&�z�۔�S,�y"b�*\G� p�Ȍ�ۢ��9�y�O�a�Ƭ1$��gW�F�~L�ȓ�8���1@��ܣ6�|:��S�? 2!h��$W��H�v`�囁"O�PZ�AD;N8�V͊7sIP%f"O���TE�xR���Fզp�F"O���ǃH8{�:к���C���"Op��/<@���X��@���"O��&dZ??�F� �@���R�"O��+�̍'nbI��I�1�bee"Oܥ���60�D<��H0 ��h��"O�$��%̮o�.l����(gfm)C"O�*e��2�B�"� {\���"Or ;s���z�8ʵ���[�1"O�Ѹ�
�Dt.}�r�� 	&p{A"OJ�ұf�	x��ݣ���2螁�"Odq��%T�vA��QE�Y�.��Q"O�t�ߎ(�@Q �B1P�m��"O4����vS�Q[D,�j��d�"O�; /ʄ+��(�l\���W"Ox�iV*��0R�BaC�of4z0"O�]��H�����@A�Dc�|��"O�,Zp`~��zT/�i���c"OP�ەJD�dg�����	g��EA�"O�:��3	���!�n�R���7"O��@��gB�	�uN��.L�x�"O>�%įt�T�kG-W&b��	�"O��s0T!\8�%��4 ��;F"O^d��@,r(VL��+��<�"O�� u����D �k��ᡤ"Oz�����
*Ⱦ�5���8(ڂ"OB)�t�L�u��8�En�(L�6�!D��S�]�\̔H�R�ߥ&$��aS�?D��)��.b.���w��=���W�"D�T9�Xb<��xcB�=g������?D���CC�,n*� �b�p��u��;D�l{N3��u�H܄^5�e!��6D��I� ���`��@�R��T3D��{��#d��#��#��ԫ��0D�����=%���=88���e�<Y���.60��d\�7D.�2�O|�<q�`/5 �e �"�Ҩ�`�<��K�2Cf�[�'�� +xPH���Y�<��EX�g' 9[�o�?v�bHBe�R�<�R�U�ҽ�`Eξ.�9"��L�<af�E�S�����
 $mz%&_d!��7� �VݝGV�!K��&�!�dڻ>��]���I�v���d'�?j�!�d��p0,\�����d1Pe(��e�!��@�Ĭ��+`L h�,р�!�$D�i�Q)��49]ԼKRK�,=u!�$߇����{Z6�8M�ni!�${^r9cE,E�8jD���(`�!�DZ�s�`|�v�ܽlp\�F*��!��:6�Y�KH!E\�r�H�3�!�d��;�b�Y6��s>L�h��^�!�ĉ" V�C1o):��P��(f!�ځP�)7�ܻUp| !�ӀQ�!�DĒY}�U҆Nn^i�R�&!򄝟릍%��{�dٷĜb�!�D� �" ��_'p|l� Uf�o�!�D�N�B�� ��
=�$)X!��T�!�D]�5cƅ#4��E������\!�Ԫh��9˧�ސ�����
%	!�ϛ����G��On��㞨�!��ɱ ����G
��i29+�!4�!�d*3����ʑ�DΔ�!��ݢI�!�� ���"�	@B֭�B�ĠT� x�f"O��Vo'D�T���ɘ�S6��"O����Ƅ4mdLl��O�q=:�	�"OH�����71o&��0k��@':�Å"O���� R-I��TJ#Z���*"O<p�r�ߙ`���#� e��}Ц"OH��w ٬U�����Ȑ��(�Q"O�9�ō0DRk���Ky��f"O��-sUbh�B��f��0JT"O4|!��ʵ6Ȅp�0c���$�"ORU�B����\�w��^�ĚD"O����8�B`I�
�0U#"O�9#�¸>N<�#k;�H�"O�ó��-˪9qᬇ
�v���"O�%�b�7q�6��g,W#��$1`"OR�g
�=v�v O�W�(��0"O
���.Q�;��$x/A�r��9q�"O��R�9hQ�ecl��Aa�"O�2 �4	���a��7d��12"OHTN�
7ObXQuc�,>�b�"O�	r�@5��}hF �tw��	P"O��:u���D �/�Vs%b�"O�يElK�_�`��(Ӓt?Qc�"O���qfV��Jܻ�dI~��r"O�8�f�?�^�Y��	:� %q1"O\�9�$�����Ӏe��u�䑹�"O��S'#<k2���dC�8���P"Ox�ѓ�A�&������;��i�v"O��kc�_�Ӑa�� )}XU�"O*@��Po�JH������P�"�"O�e�̙
';��1�X8JC(]H"O�q���I�	�&���p��eB"O�ӱ��T|6�Qr*������S"OJ�@!A��?�<,aA�F���DJ�"OR�;1�L�R�<����E9��c�"O�@�%��{ώł�mƽ	�&�x1"OZ5���0�Z�X���E�J�T"O ����s"@��$꜡R4�Z�"O���%�Z@W^�K�֙
�d�`"OJ@�'ՀW��أe��JuQ�"OD )��E*aI�S斊SEt@�S"O\�S&Օ2Ԭ����4{5��I�"O�IؐK�H�d���ӅV)T= �"O����
7M x��2��F ���"O0�I����
5��C�J��hg"OtlCq
�K"�dX�eS�Ry�5i�"O�Ht����QV ��('ű7e[e�<yÎگ~��eI�-< �)��]�<9�"�6[F��B�A}�ٻ��^R�<�Q-�Hݰ���B[a���D�<�6
N�z�r���E�:�Q� C�A�<�ć4��}�Aʝ U�,5�%z�<S*�!	��Aq��n���S�Oy�<)U�׳/� �����|t��A�Gt�<1��]-
)i�C_.J-�mJi�l�<��w!Ps��Ho�^����f�<1���Z�|��	Ȏ*J�2B�w�<��fK�zɪG��}J�]B�i�r�<���R~��4b1��7_!���w�<I��;�,���7��Ё�N�z�<i�� ]?$�0��D4[O$ e�\�<DmP�R���u�-
�d	�'s�<Iv�\7��U��B!�9ٕΎF�<��.=[��2�؇.��� �F�<� (!��9�� �a�W?u��E�w"O�$�`J�1���W�I[n��"OJ��J�)Q��p+�gqܼ�R"O�0sC僓4�`�t��S� "O ��G
��B@����n�	W8Rg"O�@�1Z�� �BP�k?~i#�"O��S/ɰ$�� I��˘SZ9j�"O\a�	�4PJ����҃ �R��`"O���F� 0H�Hq�����:B"Oh��#�Vb��\�R�@�2�ȥ�%"ONY����x-�qc�D�*ư���"OT�§H�%Ȧ��C/�?V��q"O<��NLX hhqS�Ĝ:�*P"O�@#� ^�st�гU��I���:�"ODzA�E1]��"mڅ\�T���"O���𭍷RK��(��T)f���"O�����4Kjes��C�(O��4"O�8���D'*ڜ�c¸1=h��A"O��! �/e0<h&L\+
(���"O��K��;R|bё��\�" �"OH����ق} �x���ߪX�X�h�"OV���B>�B�h�	j���sG"O%�biߠ�p��%߿	���"O(AV��
�^��ӄ�=��4�p"O�th� F'�t=����7m~���"O(:`c��F0�Y�!B�Rl��j�"ON�f��$5��!rnڪ?�l��5"On1�C�4|�4D)W�Z1BX���"Oƅ3��W�p�R�akK'Y" u%"O,�c�j�1wC��H�IF�ihdI�"O���۫GiZ�9�iϣ&��Z�"O�]#� ȥ'Q��3�����c�"O2�[Dʲ�cp- ���`"OF��_�[*�%�3]?D�N-�E"O���C�ru��Nv�UBE"On�:����������X
��eSb"O��"�B��,p	E
Z�����"O�2�ص����&��%��"O���o�,6��2��<���"O�X�t��r�~�I䢘_���Q"O�6���hl�+@�NY���"O��S����v����MkL�@�R"O�y6�z�\�!n�v��0Z�"OXDPQn�u �
Ķ��P6^p�<	vN�5�����Κo�ȸ�v�<��"�v���)�[ja0�UZ�<�RM�_�|�Zć]%b���sXM�<����h���B��"2|��Ӱ��E�<��%��Z��v���u�����m�~�<I�"E�	a���+֜X�� @�'�~�<�2��-���Q雕|����c_B�<�&0x���kד_v^P#�B�V�<�r�J�j�w�Q4��apN�O�<� �"Npp�r����~�$9y���I�<�q�S��B�J��� ��,�5��G�<9�L2H�d�(gH�$#�&t�4Ǝ}�<��Ð�\rpp����:�xFWu�<iw��4��lAFkÜG[$�[�q�<��+U:��Q�D�#J�ԥ;#+HC�<����. Nj����:J�`P��If�<i�%�������.%�����`�<F��(XM~�����Iq�ͻ�DW\�< �-|����0D@��^�z�/�[�<Q%nZX��b�Ѷ=�TM�3O�a�<� �xGjǓPH��K.��xi�"O��9O��� ��F�]�As"OҤ�`H��"c�|[��	
�Ĉ�c"O*�J���3�p#��'s��1�"ODxu��7:��;%j�	,�${�"O����H�8XTMb��.	�FP��"O`�#�l_�S}и��h�0���[�"O�QQf-  (~"�Y�� ��y8�"O��Äʋ&\iL�����J���c"O�u�b�%����Ú�f�tRp"O��s�� fO(���g]EQP���"O�Ű�Ä:���H�&T�|��9��"O�Ap�,���C�k�=��Ai0"O���1�<TH�{�F?t��q�"O&��a�ª��[�م[�"OȀ���	5~ZQZ ��F�h��"O.T��m��|�xGg��Z8��1!"O���޷,e��R�惀f7���6"ON@��J�� �uC�G\FQ�2"O�§� u/&M���1h��"OZ,��Q0h�Y�GO0((�"O(����S+y�.XRAG�R�xhT"O��s� �/�����_�����"Ob-(4薱T ���I:	�^�6"O��Z�!E�=��� #\,���D"O]q�n@�D�����̢t?2y��"O��QM:�=��o�+Np���"O8Q:3b=UB��!��3W�T��"O�l
���-xJ6@���D>l ���b"O~����R�J�x��k������"O�pR��ʫ]	�0x⯘<n�f5S�"O���g]�@����{�,д"O����	�7<'��I�a7&���!"O��;��  �AF�{�ڵb$"Ob|�S�T7:��9r��Mj��H �"O�X���A��d�C�C�P��"O�*�삅F"(r�R�>l�%��"O�,j�d��w�\eIp��Zz�d"O6Ƀ���1�p�AT\�vlz0"Od��1B��d� uSQ�z��ѩ�"O�YQSCG���DY5��$혴8W"O:�Z�D�?��0��I��0�¤/D��b���wĔ�a�e�,�昡A.D� �!C�����Y�坶W)����'D�P�gg�3?�bL�vJO� F(�;�n"D���ǅT���6Utd�1O"D�(�į��\�X4���R�.���@d!D�l�E�V�H6h0�œ�a����6�2D����_�6��άKE��@"E1D�̐�B]�M�4�r��md8ys�)D�t�3�c�r!'FSkl�� <D�t1�h�+�1t��lP���E�;D��b��˗iJTR�,'^���Dn?D���"��O���)`�?|����'k?D��:ȏ8F�$3q�\?/��|D�>D�!Da�	n�@ 
�"zBp���k1D�(�b�]cVd���쐠�w�*D�$�e��v�0�N�D�"�	A")D�(����rx��1�B�� �H���)D��KFm�H�<)0���_Ph��o'D�����=�Ε��Ɍ�;r]I0&D���@k��i�|��텯\�C�d9D�죃H����܁S��o�$��bD8D�x9�@թ,m�)��%�K���1�5D�� @� lX�ZL����e/��=s�"O���lN9eb�
��$>���"OҴ��F�>jI�eeڷǲ�у"O~���MM���&E�I"O@�q#NE`�A��6Tv�ˆ"OL�'��@t�pl�/^6���"O��8�a��B�>!�t�[(ZT�1�"O���rCɄ|)�T� �L17��zA"O��SCn�_����s�" l�K�"OHȪF�G�\��a��^��0"O�`��c��8����nͮ]�<:"O�m��d� ���;�#�v�a�"O��cP��(
h��I �*̙S"O�9�Ê�$5�x�ˑN¼%��p��"O&�!����K\>	1�� �Iwx��"O@��6@O-
�&0����9R�b-!�\F<�:�m�>*�īӄ�4�!�d�B�\��H\���ػq���!��X��uAt�	Y��0����!�$»05| ;��Es���Ю��l|!�DT5K�� �W�r	�3�6rp!�D��!��Er�g�yC�����7c!�d�&'Z��@��W���5�J�/5!�.� ��Tf�D}��RЬ?�!�D�je� 3%k� J],�u,�V�!򄙇<���A�ۋE�0h�H�!��ժB�[��B�DrD��!�<bZ!�䛯_/�u@GJ�*EF�Rf�5f!�D�=|�XB`�@0Y:� ���-|G!��:[!Bu[v�ŭ,Xz5@��X<a!���-k�[�A*?Ƒ3�Tu�!�dҷN�,#���J<�Չ1�!��Z�e���F�3'X���FnZ\�!��'�!��D�1p/� r��F��!򤋠��ݹ��!&�EɠFA�t�!�$Z�B�ˡK�%^�0���EgIp�'����,�le(���E��yV��'2�e
�d�8zln��g�=���'D�4����X3��)hwf���''>鈃��i8�j��dU�A��'��SǊ@�� ciB<`����'[fa���q>����Z�T�l|�
�'��4x#G�+Հ 0��6P�le��'ؐ�#��K�F�urP�[�����' 2 ɓ�ǨO���5�>R�j�x�'�|}��ΉL��$�i@,�A�'�J�a� �g�X1�tʖ7&�'ՖX�!�+6b��y�`7~�n�!�'p���@�G�N�)���y�Vi�'���h(cp���_:pU@��'�����gK�GT�[&@�pY�3�'ɶ��!&�Bk�o�����'S&ԫw��$���+@�] �	�'x���'AT8[(}󡉌-V& ��'��M"d��D��uq�ԓJ�@��'�<�H޲]$����7IB)��'m�%��� �f�����?M|��'o:�Q���P��%�$;��Ȱ�'���j/�!|r�;� J�l��'Ӓ� ��_� j'M_NLv��'����q*˷Ԅ���G!D��'h�ёGoXld�f���}����'����䉧/	na�bl��t��	�'�xӱ)A
)Ҽ���! �9���� ���Rk��P;AGU�h���D"O� �*�Vn�b���g`��c"O|��!�15D�!1'��\aΩ��"O� HC�7-�`�S�E�+Y�Ӏ"O�U�#�Gvp�ʔKJM p�"Op���*AV�rP��oߟl.��#�"O�\��5pظ�
T��n5*h�F"O~�@� ɪyx=�dOB9>�ش�"O��+#G�^�eyu�A7x�BDK$"Oΰ�e�)&�蒋ќ���C"O�]���	4��� �j��6�̠*u"O)9fGB�(v�̚���;1����R"O�;�TQ"���hԬ=�R�P�"O�e�U	�Y������H+h��D�U"O\1���_�HfJ��TTJ�Z"O.�8w���w�.�S�K_�o7jI��"Ot�f���v�����bMYs"O4��G� �+���'`Ċ1"O!��ԯ��}:�M�>!�8D[S"O����Y�<�B5�E�׶��u2�"O������$X�˗�Sdu���V"O
l1���2~E�����J:<�l#g"OF�2�̔]�0ĩr�� ��p"O�W*�8� �-ϫ"���ʇ"ON�e��{u��p��2���X"O,Y�3�-Re���,6�^-��"OL���!�J�h٩dK=,����"O����Z�P��As�I>� Mc"O�d���ڌ=_�mȡ�W�'t:���"O��;C��.W�� C��cY|@C�"OVu�gi �B)!�bT:r���"O��C�J�VZ��SC��F���F%D��b��cU�=�W*8���j��8D�bT`c���HW?I�6	Rt.6D�1ǎ4+�QH��3�R]�p�?D�ܹ�f�p�N�D�Ij}���>D��S�Ɂ` X�� �Ĥ*�~��Re1D�LÕD
q*JE�4c�?Wb�)��,D�@� #<ݜ����@�=�x��/D�P Ҍ�g�m�BȝYfD�cC`:D�Ds�҂EW�0���
+���=D�|8Rj�i6|; ��Z,Ёd�7D� xw#�Ƞ:�gU&B徕��2D��k�@@�;�B�凂j�~=�q�/D�x+��3o�$ҵȂ�i�Re��(+D�<�#(ѐW� ș��^�Q��,�to$D��"�9u�����ۀP�����5D�� �<�8��]�P���2��0|"��:RlY��)q0XiX`�X�<��^k�N�I�$�ԉ+$�V�<Iu�@�*��ݙ�"�=.l�|�<ї�P<m�! (�&0{>���B�<A���c��!�cڥӰ��y�<i�h�Y�q�`R=
,z�����u�<�J�	�\0��8C�čBBe�o�<�'�*E ��ȃe��ͳ`��y@��O�Fiz�B(C��9f�Х�yr�1W��x��	��Ҡ"ՏN �y�lr��)��7A� T"#��y�[�G���s�Lע/8�m#�'����lK�s5ZU��.+��'��	��$S3��q�(S'�\�:�'�Y�$��L��`б�,mjΙ)�'��� �o�:X�"Բ,0� ��� ~�:u�F9��̐a�r��cc"Ovp�׋J#|��7����s"Ol<�0=�����?�RD#�"O.PQ��	0ܩ;�\�V����"O��.��F����DM�Xj�X""O��X0L�-Jc6���6L�Tx�"O�%rn�mZY �ʑ5p�Hc"O�9ҡ�m˒��^k�U�'"OJ��wj	7߄���Jɉ lp� �"O��X0%N�
!(ޏP��"O.XjbbY,� \����.�}�<ɤ��:?�eZU�ϋ.`)��n�<1�M=(��`h�g��$� �Gm�<�V�'|����@�0FLQɒ�A�<�3jK�K26��Y2[&����z�<�G�/B���@�* �B�VH��(��{��n�Ma)2/�w�!�ȓU� �؉Q��HY � �(wH��ȓI��AĎ�#sM��c��{�����c�\	�hȩ9���&"�.ц�|Ŏ�z����9��p���AZ6m���|���,ϟ1ʆ ��M�����ȓH��@W �I5�-Եi~V`��J��a!����V@�~����W�V�Ip�Ѫ^��r��!%�Y�ȓ ᦼ�/3)¥0�D־מP����Pv��hyt�S�D��.��d��-��[B���Z`
�3t)�i��}�ȓE�� ��"��n)�p�e%֍c�L���
� ��R�A�{GS=�(�ȓO+�X��C8�A`��M�'�(���u� L�g��Fz$���l�&Q����D\��s,�@�K�D�+ F���nÊ�3d��Ӻ�#���hp=��8I�x�ɉqW6 �RfW�a��d��7�P��aʘ d���Aăh�~���JQ�-���
f>pY��'�38��85 0qTƍ4	T��"��ޛ@���JTc����H�L�+��Z�k4C�I?_���Vk�6\�����ӮZ��C䉂Dlp5ӆ��==.����O�9c�C�	�+'�=@k�>��$z�	Y�K�C�	EZ���K/�@�4X�Eu�B�	�Y������E�|��Pd۝B�bB�(yM�-H��@Ԛ�j�>B&B�ɝa�p`�SaU?�������.�C�IjlyS�,Xȭ5Y�5{hC��t��EH0��7D�T|i�˚5�ZC�ɱ2ז���	ti�]�w��N:C�	�d�^M� 0^�.�TJۣKC2C�b)�z��i�Q'6t\�����>D���	��A6���B��R"`EȆ�=D�D9�&А���iҚG�*MT";D�����x����Qb���b��m:D��"�#mR�1� jͨY�*�6�8D�����QʆtAB_�u����Q�5D��`@*8Bh�Ib�&�N�e�6�4D�ȐQ�+4p����XK2���ւ2D���A�J>)�M��Ӝod^QZ��.D� ��.�z%�с6!�*SSNY�`"D��Y�K8TC ̓RMV�}:�@q�@.D��q'��'�\$@(�8y�(���0D�AЭ��A6zhR��S}|�B�-D�ȹƋ�����0qbS/p�DX��,D�� �E%'���`qA)�4����"Of̀R�� �(%K�ş�AN$$�"O� [�_�/��РJ.5j��V"OL���l�r��*��\�vD�R"O�DɱI�3$W�����A%rB���"O��b�G&N��0�	#/� w"Op�3�Ώ:	�������!&�|�"O$���M�?�ȃ3�I�z2E��"O\��q�3+�����hH%*�9a"O:xpM��x��d�����|��"O�"gʅM��4�r���C�R����'�� ;T��"g*��D�	�_�(��%D�´N�B�T �1G�V,H2�5D��K�G{�ะ.��#��Q$D5D�+#n_�d�*�RP�ήy=��ѥ�1D�2P
˗i�@{�"��

'Mv!�ĎY�"m���O% ����œCk!��Rnȡ�ۮZ�f}ã�r��ȓ	@�Q���	?���I�Ȃ�!z��ȓ��VC�.gL9�oP�5�	��eT~e�F�O?q�P,����ZZ��ȓW���I�L|HZ���-�����i�ʝ�/^5��a-�=�@�ȓ<� Б��9V���GE��Xe�ȓ��
GC��EF o�Yc@!2	�'���4/@�O��;ÁǵP�v�[	�' ���A�	���r�[�0-t8*	�'-t� uMq2�rqa�<wҀ��'��	��C'�B�Q���oJ�D1�'i������<JF�cUA h��,��'V�U��f�n*(x����J�"�'V����K��Zض��Ꙇ7�u�'�ju�66����3���R�'ِ��NZvj�	%&��F�a��'�-@�+����SAS�}96p2�'�,�������R�z)��K�'�Թ����V2t�+"��*�U�'����Ϛۀh�.V5 ����'�"���h"�(�P䖝r��'nHSP�"9<Ѡp������'��!�GO�T	���9���'/�!�D!�e�z�I*�yH.PJ�'��AQ���0b
]Y�=xm�r�'��@��aҖ��Z�&��`�
�'�P�sF
 j��b�Ƚ`�@���'�.؃�ůK=�x:q)�0n�����'IV�!U���b5�-��g�	dh����'s��١DUJP!�֤2�L1�'���0�L$@�{a�ס bP���'���Y�ō3W�H��`�x��E1�'�((	���	SY��p��rtZ�"�'(��sզ�&kL�T��K �2ݎ���'�B)T�Q�`r��wܧ1���'!��% A;�H���卾%���
�'z8<)@ �~�X�rbH�G��	a
�'���+eD��= Ⅹ4c�/jn8	�'�� +�5� �匂�gp�1��'6T��z	�j�H�0��A��'�6�����^s�ɱ# --0f�+�'М��჏4&8��S�J#+C���'�t��N&M|��*��T� Z�'#،�N8fH����G�MD��
�'a�����=��t;udQK�f��	�'��Y���87����!Cb�{��� �-�����8pt�{�dI+�,��a"O�5gQ>-�̐���m�.� "OR�H.N�9�B�Q���@�"O�#�	������������"O*��t.�"	0 M{�m�h�~Y�r"O��DD�,�����kհn{��"O��p�g��(��d`y����"O� ɦ��6h{��Ү~{��؆"ON�O��z	�� 2�X�'���e"O"U ��K�JA����ג8�.A T"OڭjV	P�	�:ؐ蟺��
r"O
!`��\@`h%��;0�̸P�"O���#G��6���F����["O2��Qi��FӀ�q%
�&�b"O�A��N�5Y�(usօC,I
^E�d"O>�����$��%�'O�<�1"O0X�'[q 8t�Qc>e��2�"O(�J7��2"�VYs"��z�\�Q�"Oz��ǎ��>�=���H���"O� `��Ҷ4UӠ"G<X��"O��!!I�N�(��F�G�<����T"O |�1�	!0:���j�]��9�"O|A3I#}(�Ai��0:r-�c"O8��E�$K�6��"g�6:(��U"OTKs�ƌX�A�Ǥ@�f?\�"O9;���'3M(2$ML4���d"O֭���u�6 ��P�<��K0"O�����G�:d� $(8L��"ODqI�(%|�>l�W�(N�u�E"O�QV�ۙE�^�cW���F�4�"OR�㩇�k��y��eV���1"OH��A*Va��ʣ��0o��h�"O@D��h�Wj@0h�f��O�:4��"O�) !aݮȦ���jٯ#�Ҥ�Q"O� ���8Zy�ՉV���X��"O�[��p=�Y;�a��|�FE��"O�ܪ��ټc�<Ĺ�*��s�ܸx�"O<�8Њ�' �2�k`���$����W"O^���j�0@������%x&� �"O�q���J[+�15J,J���2"Or,ӗ�S�@kXL��� x��LK�"O�M Ѥ��ثE�����p�!"OF1���#_�T�+�9�2 %"O��'%�ۘ����߭YKB��"O��[!��!�t��$���#lEq"O\��J=S��ɵf˴H�	1"O�A�E��p�,�bg�t~��"O�0"Ⅲy���p�Xa��y�"OD���/��1�J\��A�>�vtkc"O��J��A3wqT����"����"O���+�!h�~��4$��p� ���"O�ɑ�FL��������`�"O܌{�oB�S>� ��&>���{b"O��86�M�`��Kg(пp���a�"OL���n�b���Ň eޢ��"O�h0���u��A*`C���b�r�"O�|�M�8vZ���b˽^����"O@Q�LY�'���*7+	���Au"O��2R)�TE<=�� &"�����"O&丰gZ''E����$t�L�[e"O��#ׅG>Ej��� %̫l܄�"Oz�J�Ă�<5�$���L\$iHG"O����<�DN���=yt"O�I)'甝V��Mz!���@�"O� ���T�7����E��l3d"O��׍�7Q�ր����)�� �"O��YqC�%^x2q����|�P �"O-B�&�
4B��R�Y�u���%"ON}(�n�����)�ݒ'Ϗ��y�+E3�H(� Fc"�X3���yb#U/�F!���G2��c�ݻ�y2�LT�`��6�}�(X7F���y"/N1(?�eo�E	�����yB�9J��X�BN���s�i^��y��Ѵ�h�H
a& 6���yb�G慂�qx��q��O�ɒm�'���0��SA�@l��"8P���'�^%���F9`�=I���j}p�'X�!��eU��c%oН��%��'B2�bB�W���u�4ΓX���K�'�Z���	��'�I$-܅R�4��'��Z��N 8=���p�Q�B�<d�'nn���.˶D��M�5i|���'�VtSw�?���7�@0rXh��'R�W ��>��q�7��� y��'�@��g�a�
��F�8�(��
�'Ѿ�a�g	�$@Gf��w�Ѹ�'��@��0�<�C�ȝ�s�"ma�'�H��6��/\j�sq&�<o��1��'o|X�$�20�����
pF\��'�v�qD��@_h�0Ƃ�t����';���tƌ�MX�0���g��!�
�'��(&��6 n$1�N:XS��j�'�����O����J
N�j@�
�'��h%�G�B]p\�'��96(n�X
�'�F�����З�:���	�'��$��*X|tRw R48h4�
�'W��E�͠K�����)�����'��'*Jx�5�3c&M�
�'3d����#BR��!A-N*�"90
�'��Qi��=7G�h�	qnF��'��TɄ�R�F��=(��]�k�L#�'N�m��i��{&��;�/�9e���
�'�`�E�Q�SM�q���%��Z	�'몭���,I���r�B�$�%8	�'lL跊�9(��C��n��d��'�bX�BC��g����g�1c�� 
�'N�cʄ+-�P ����kwp���'uH����ϰyvl���^�hG��S�'��U�2��ZK���U���Q���+�'žH� �]�+6$)1Kٯ8��X�'�8��ǜ5Qc,�h���&�F��
�'�B,Y���p��I2"E�߄ ��'V
��O�.h��J��H�ި3�'� �++���ARb?����'D�������0(�C,:,�e>D�Ъ7�՞2j6�)�I��e���)D��.�<o��, 䠞17�XY��:D��u+}DU�5OA�f��=�G7D����0ez|�9Q�J*Z��P4D������G�H'��p���%D�PФÖAI��
�1���z�!D�@h�e�:��G�Xd�Qpbm:D�<9�$½/)j9Q@L;�NE�rM9D�x1vܨI�`��#�>�����8D��� �^�F�2u!��T���sd�6D��J�nu�\�g�U��R%5D����@�<"��
tn��h�f=D�� ��hcZ4[��p� HZ�3�"O���V�đ;I���bDʫ}�( g"OD-ZǓ/�2�X��=%��y��"O
E�SΏ6<.���Bؑy���c"O0�����z�: �H?%x�q�"OPH 呍��5a_;d"�s"O�ăăA�Nc�8P�7]�2Ƀ2"OT�(��υXa��R���y��m��"O,U���G"(��(s�B!�΀�"OB�z�c� �җ�>w���#@�y��8wv����ף4(b��e�C�y"	���5 �b��<�mR�!'�y2��aD���s��]�my��E��y2a�+_�i��	O0k/6	��X�y�$?+ԮE�wk�>07ąH�G
��yR*�nD�@��%A�|@ŅM��y��O�t�eS� U��0�R��	��y"�7����Ai!$��YS����y�郞mE����+�Z�Z�B
��yr��7R�%�6�P�d��ǃ�yl[w�YYwKQ,@24�s�ë�y�*�3�x��Ս3 �X#�
�yR�9<]���ţ ;P%1�ǔ�yZ�'V=1��wl��XT���yR��W�ihbÈ� �VX1h�y�H�(�`��c�)���aS��yB/ȗ�

���������',F�!�D �d�8p�X	�DB�'_��;de���Z���X
�'j��5ʜ�Eƌ�qsK�D���	�'�����,<��c��Oi*���'��8��2`��`����RЈaJ�'��UB��5
��Qz�B"�-*�'e(��H�l�ȝ������9�
�'�D�)%$
�x@���]�d��j	�'�p0 ��T�ReqV�B1X��y�'nV��r	CC��ʢL]�R�zhq�'Hh] CH�g��y+���Q�,e�	�'u��bi�>zbC�EL�l���'��J��(�*���IN�h�*�'ƈd�(�>�)Ċשּׁ�'3�d��o�	�����`�BL�'r���ăT`��Cn�6!
�'AP�5o�BH^A��H�a��x�ʓ&�4]s)�	08hy����L�لȓ�4!K�-�]��[Wݸ,@ܑ��G�8)��\'Ssĕ�%� f�`d�ȓp̄�	g �=Y�r����<v܇ȓ8H|��	�Є��b/�5Z�p��>��02%O3J2��:2-���ȓG�BA��Â�H@HI�"ɟ�U�T��D�
(V�ud�.�mP��>.Ѝ��B�x���a�'�
a�ȓ��\�$�	32�{�N ."W�E��9����![�Q� `#$Y�a���],���R��&<M�UC��]+` P���ޅ@��Z8X���M+'���ȓS'�Xk��5Y2h�p�]�Sm`���M��A��z�h�"���1Li�ȓ�ܑP�5;V8񠂂K�$��e�ȓ/T���析;�xm��#l���ȓ '�� ��NL�ʤÀH��}�lɇ�f�ƅ�G���r���C��_���ȓ u��`�+Z�h�jR��'s|̄�S�? 4��a��	�b�I��<���4"O>������ZŨv�ب	�-�f"O~����ݵ!L^�:C^iв`C�"O e�'���16�(�(e�lZ "O�pʷý5��8��CO
w�
��"O�B�ܩgf:���қ�X�`"O��0Ơ�$��jF*'X0���"O�0�uo��v�,D�Q��H+ڤ�5"O����`�-l 4Q�Q&N�b��32"Oڡ��iF�k�jV���k�^ ҅"O�t��!�3^��p�r��@�.%�"O�hc'�ۜ��w�V��`��"O�\Hg�P�Y@&u�F"ۖ���S#"OR� ���"5��K#Q�X���T"O.���#
R��\�7G�~pYB"O���'a,& i��8i�Z�zs"O��B����%0���56��%qP"O�\r�/�)��87�n�~$�v"O��#߼g�lU�g�_���pQ�"O�҅e�?�FT
�Ν�b��[3"Op��H-�}��O٘1|0L("O����1;!qՎ̰obț�"OH͑d�F&Wi�<���=,����a"O̡k���D�\�Ѧ�
K���W"O��ȹ*�\ћ4�I�h3:���"OBQ���'n½d\=l#��i�"O�`st �h_� 
5�@,�0t"O��2@�чL���ʮ5�B�[�"O�@z�.դi��`�a��/�d(�"O���I�(�b�b��Ĳ*�x}�%"O����3"Ѧ��V#�Qn�`{f"O0L�R ��;����a�;\�r�hb"O�y*r䚷:�hh�Qk�'w��e�"O(9�@�6��u"'��u��zQ"O�X����*m��8k�HA�@��a9$"O����ED�G��3�>�bQ�&"O�XӦ	�eoD�uF�94�d\`�"O����ù7�\�����]����5"O�}1�ᅓ6��4�ƤJ|�-�"O�5B�ł�4Q�%C�W���v"O����-�1`�^I8L�8Fkv}�^����i领�OA�nY��w�j���"OJ�#$R�R��"j�!Ҿ��"O��s�*iF��`�XR���C2"O�R�	�9-�p���6�6M1�"O�%R��X Bg�_;F����0"Ov�	aN]�x �$�E*�*�X�i�"Oz`P��9q?fт2gJ>,�Vaq�"Oz��)C�p���Bb�Q>f)�'Z�'���� F¡d�t��!�0�~ I�'O�e����#K�0*r�p�}b�)�	�>@&����LR"��C�In?!�F�dڨ��xN��*�m�6	D!�d�fL`�lޱQ�ٻᎉ)�!򤘗V��!c�6mj��P4�+T�!��V7q��R`��15�`�R�,ۨ)G!�DQf�����\2�*U����� .��0�O����CH�q*�%Y�ߙd�xD&�Q̓I	H�O1xX��ȏ�w�p����Y~�ȹ�')J�ʄj�SV�8!dS�J���{�'^>��i�p�pA�� H�Ε��'J&�!�F�YL�2�*.� ��'�X�l�&l�Q��� *����n�h9؁/�}���D��:!.L!��S�? ���,F�8���r"��l�t8���2�Ş"]DYsG*6���@H�^+xX��e��X��S�bR4��"ź�.e�?a���~J�c�	r��-�FC�$PD�#�r�<����� \�0�Oy�CRm�<1��� %�nmr��7	g����I�f�<Ѱ�^�.ECk�1l��=	hl�<�g똨�0�ѱ�0=�܈A�O�<	A�P�9����^*B���(F$�q�<��� �*s^� �O�);�;��ʅ���0��s�x[��H�*���CS� vIC�!D�d1�+�;S�~ ����q��dk�,D��(t���
J�1��)/ؐ@Q��4D�XÁ'�hz��a���kڞ��7%4D�$�5�J*{f�c��),��1�
%T��;��T�.�B����&U��iQ1�>�
�Ath5K �g0�5��#A�P.Ԇ���c��[�6�ZzC��	!�������.W���<On\�3�-u�tx�w�[2E��-5"O��S�1���k�?OЁK�"OZ1�^XՋ5M]<-�D��d��.�!�D�D	�T�R���`��ӥ�Y��!�Z�6O"�5�K���2
W$0�!��L�m�h��n�Ve�J��*X�!�!te������8���'G�Py����9nY��	�>��풖���y�	�h�x%��0Ԑȓ��T��yΓm���	q�G*d���5Q9�y���EL}X��s�V��u���y�F�g;Z1:%�� �%���N��y�	�R�QxC!V�ҳ�N�yBL���G\�I�Hqt�"�yR�{�|� !F�=�Թ����y�қUH�����˪/xLUh� ܊�p=��yr`�V�����I�3{�yB�P�VL8B�I^����R�_Qj���$�0�$��D$�	1x^�X���/L��IyeG�D�0B�I�0�Z�jq� ����f[�Nt^����>�Viӂ!�S�ܵf�\U�v$^h�<�1�����9sdi��c���ia,�f�<顃M�k�t��W�٧+cHL�S�Kc�<q�靋�Q��
$�z�Ҫ�^�<Q
�܍ڰl�%U���J�U�<�á��a��hT"I)p��;�AM�<��0!%�Ӧh�37��~~��'=�ͻ�G^ZBt%��g6���b�'���AO���>�j��7B4	�'�bD(4,��E�����L}�j|j
�'E\�3w̔6=t��҅��r��S�'��Qba[���EPv�!����'r�Y��a������M�hj�'8\m�b1{��8QFFe�5��'��o^{~*�bӬ��"x"��c"O�� d�7p�z�c�
'`�|��"O����Ȼ JY�d��s��#r�I�����"]:t!���A%(��DE�>!�L��D�Ԋ�c�<�4��Y��|��x�E';�^�*A�;7�2x1a�Ŧ�yr���V}(8PT12 oֺ�~$����O����b�OB��2���(�,u�"Oꬺa*��L$ ��8��t\�0����&��D� ۠��`���x�pC�k�B!�%C�u� �{�@\#⟐F{J?�ᗦŸb���E�E��u��#\O�b�� >����G�-��-�g����!`G"OPT���K�"�&)�4�J`_|H�����n���1ɲ��(ǲu_�l{U.���|�ȓ=V<eB0�Q")�P�%A�(GyR�'��و��.c���S��\�C�B���'� (�����u�Z��co��=Щ����9O� r�V�����fF�pdP����J���	�
t���� �j-���A�K�Py��A%N���I�n��<N�[E����yr��B|p�aG4	��ʴ�N��y�향J��жd�$�xP�Ԭ�-�yR	�����Z�˒r���ꋋ�y�"W
f�X� �U�b�!F� ��y�aڌyd���KY���Ɗ��yr
P�j�80GO�M �L�+ӥ�ybb޽MRac�):oV�g���y��&\�|p�d�W�7��<9V�Ö�ybK@��@��欁�=R��
�-�y�A�#�۬b8ԡ�EZ;�yl��!�,0@��/I`T����y��3� �+�I�'UB���BF!�y��V�f�Y2�"S�2h#p%��'��z�G_��
�8� D�M���J$�J��y���*���z��/Qx`�
�L��y�"�<�A�	W�Y�0�z�Ô0��'�ў�����@'��7#|)�r� G���Q"O�-[bo�% M�!rc� �hF��5"OVh����:�n�B��S�f���JC"O&` ���3!��Ի��@�w��l�B"O�04#L10$(�hT��,@�"O0� �#&6d��&�D�\ɑ�"O�P�2�P���1��%��Y�|Q3�"OpQ�҃_!Bo ���o�N�8 q"O���e�G5� �ؐL�8��i�&"O4��"+��9�.����xyl��u"O������	%���qBc�Ը�`�"O��2��˩Tm�阂$��S"�I�"Or�A��E��������5"O������ �Ĉ��A�Pt��#"O­����>	����0��&qiw"ODhC�Y�.P~d�5O��R�nER"O�-:�-ˆQ��paK�I����G"O�Hʵ��*E 8���KԦU�v���"O�a�,Q<l�8��$Z�)�p�"O��ԣ�5H���8@�_���3d"O@0`��M,,I��I�JAa2"OZ� ��*��!���~x���"OV\�Tà\5X��A�F)t�v!bR"O6<+�d�.>�{3M>2cJz�"O����Q��c���lR	k�"O��p�`�~�n���ڻpE~,*�"O�8s�؟qB:�����Y/
1��"O���B������ȓ.G� �"OU�h3]f����ǈ ,^lT�"O�٠�AK,|�)y� `��Ys�"O ��b�ڄT�%��G���`�"O����.�����,��͑�"O�YW^�zQ���5�ڭ	W"O@HA�ܸ3̲	Q�����5"OF�0֯:�dڵ%'3�ܠP�"O  ��A5O�|�Zf��3E{����"Ov��@2r�2ĪD�HU�[1"O���$X A�Z�:���5a����D"OJIb�=t�A�튇@�mPg"O� 0��E��2����k��+�0�)�"O��"Ą�G�ظ�B*S�?<�Z�"O���5蝋����F�R
+CZ�� "OP�ad��d��D��f7x\�"Od��"X<B`5�腧|0�q"R"O2�!ւ_*�hLB#G��K 1x�"O�� C� 0�2���%Ǳ1Z�`1�'@��b�
"L��OǛ%�)�bވ$U�Ӈ]��\��'r�!�#� vz� r�֋6�jT�	�'ɔ�[bM���Tk�E,� q��'�x���J@�ad��|;v�x�'��Xz5/B�]$ fKזe˜S
�'x�	�&Kԙro�1C��\6 ��
�'<�l��K�n�p��*^�V8
�'��<��ㅣps�Q�a⊤#(���	�'gU���ـ�<X&��au��p	�'$�!��p�6���*K�VR���'s���@�)��9IrJ$BԚ��	�'�`���6邑���E5o����'+���Wd&t��@�'�!U�.���'�޵	0*_�kOLUb�mY�Gtܱ��'���Q���.	zBt���`��T��'����6�&�A�D�f`z�{�'^,�i��+7
t�x�%V�R���B�'4�,��(��.4C#�]:2d�K�'��ɂ�`��p�~,��EK�+�� ��'��i�	�8y0Q�ƫ	�']��'�|d
��`��y��ܛ*�5��'iJ�3,�e�H����_�i��'���ih
-(}����WJx9 �'c�}qӯVs"�c��_�<m^��'�p���L-1jj��'�45#�TY�'d4e��" #�����V'�`��'�*q�B�G���R�i��  E��'��4�K��J��EbN8
:�	z
�'PX�Q�D} �̡ee���
�'�:��3ϐ?V|�Pb�-S&�(2�'(�)�D6o�ȫ&���P��A�O i�����O�0�`&%d7*M���ߐB� �1�"OFq�dC���r}����,����1O5#!��&{N�ņ�?
��8y��W4����B�iD������)���&D�����D�[�K��Za�P4늅��,D�(�r/��걢f���>A&��-��H�
]Hӈ
<z ���i�[�5�4$�']��+v�\	#U!�D�"An�� �N� $�)S^_�!2�	�&h�����w˖-�d�XP�g�ɏ��)å$�^����o�fB�I��1��R Af`��n�D��\��^&R�fG�%�B�x�ux����98��A��}��h*dI ��z��(�2�Y�Pm�Bs	���d����^-� hH�Uè��Ua��x��$[R���[TRg���ѕ*�%��I"c��$�TMN/W.��gMD�j��5
&�i^:��1��R)v�Ȍx�
MN�!򤎃w�e���63�9�U˃f<� ���;J�I3CY�_�.�(V�~
��r�I�e��u
�,��Z􎕉2����
�d�7��8�lU�C!�1ta��k $\�<��a���>�ex`�X���$ӭ#�pI
ל~�A��%	7�ўp�4+�&XҰ���k�"A12��5H��d*�Oku���t��x�^I�ȭ��xBA?��媡eϕi�LDH����?��I��P�p�.�#u��ӱ�D�������IFe4"1���Jwf͛4�5/LHB�I�6�𵆓�s��-Z�D�O�VI�R�Xf*M1�J��#D-����|�%�*o��'��D����DЈ4�4
�K$�݉�J ���`j��:鼅[�E�,d��c+�B���d.;#S��*6���;����),O��ZC�F�m�Ȁ%B���x��I�>��t���Z%=�u�f��##Fр���C
� �ʔtݨ�R�� �>������o�DY���l�� �%U0D����mT�P��ؘ�a�OVsTI~����J��.���n�(e�4�kE�ک|���qk
��� ��b�F]"f%��`C�Μl�M�`"O<|���=r3�s1-\�$�V�ː*��d�K�Û3����O8�0d+��=r1�K�M?#�H��`:�h�Ѣ�Hy�V8*f+�.��@�'��9���+7^��1+��h{����2���*����Viiፁ51�P�`�k-�D���U�T�{�B��D��x��ˇsΦi*� Q��hO,��/P73�vݪQ�]1o��0$	C�\� %���:ٸp@h�*ժ�R ��+�����
����2a�*LOB�E?
bdۢk��2 �1Z�M��߄;�A� ��$��	�=#�}`����aB � u¨�o�];�t�g�ǡ]ZȀ�"OjA�u�-�=���;:�|mSWW�\��=� B!�д�'�zy[gC�g�:�*.�Y���ͻ�)0�M�uɂ�SC�5F�V����5D�X�!�Y"�<�դ�v� �33��3GW����'	��k��^[��T�m �"�ʸu��c���͝q�:��$(�02X�LI��3ړOBz� �ǝ7I|$5r�l�.\̓���17�y�%��3z�<0��b�~K;�"�jؾS�JQ���cG@��ޕ���Nɲ���O@�0!Μ�?�PA�1�ЯW�-�����ġ��H���?���0u @������EA���׍�?����!�� ����˟_~��r3%ސp��pX�h�v��ș���/5W�97�%���+K\w��
��v���:X�Vpc@ʼZ�,8��ö+��}�#C7(�֝��b��7�-elQ�&eԐ��m��Px�.�f��h^P!aA(�M�C>O�~Xz�c�JÉ]�u��YHTAj�`���7ړ_��l"��li��[�4�I���L�p��	�Q��� (^�|��%S
ڳ��a�X��]��I�e��:A���P� gC
\��Pf��Z��+@}(��u��b��B�T�d��'B�_��H^cwd��BH�,K^�r��P�d2yq�'��c@orцx�PX�{�\m�ԯι�\0y�-	��������N���Cp/�pԌl� �(~�FQ��wN�!8���2�1+�AE�@����R�!4폾RH�p'AE�D��xAG�$����G̐PP\h���Rj��"K:	s�0q��C��! ����&)pބ;�kV�c �m�� �R��O,�"
IZ�1�.p�<�`�!*�P����&ܒD�uh��LF��)];��2͈�_�-�D@q��$c��3������ZL�N��ЄU�t�,�

:J�Y�������q�"+񪊻B�I�����JT-���\���0+�ڎEp�9Y|B�	)��x1d�Z2j%��ܝ>����m�D��##I[��)��H���d!�D�_>|�D%1�֘5:�X�� C|s�u�.jL���
ۓO��ق��h�R��'��`J��Zm���obH, �$荦��Q�&G^�W�Iv$�H��\2AI��jp�Oڰ��,�/��Q�N��3�r�ٕ��L:ffM
BN�~d� [���:	Д��Ɩ$3'��kD�3��F�6)R���t��	�X�Ac,�e�q�
ߓ pd��D�?J���e���
R� �0&�㖂 Q|�Z��|iA��E��a{�F�*�j-X�̸p F�Oz��L�͹3��/����ȓT�Pҡ�GĹ�>�.|35�T"q ��Qā��A��6P�^	�����L
��!O��0@��T��"F*[	M#*�	���)>�\���'��(�GЩr8����3V!���J� J�t���A�XYa�#��qr��[��h�hT�<H�A*�Q����q�,��o�8U` ����' l�!T�'
>�����=H�#� �D8P)`p`©|2d���$�EE2����ޟ6�l���[ ��)�Ă�Q��Y�`+|O�!��w\����/B�X츽#�C�2~E|=AW�؛~�2T�e.�%2�����pS��͓]⮡�C��,� IוJ���VG[�ݼ�e�'��E�ҿ8�<�@��Z�q��(���X�o�r��*��b���QW����y"�W=;�4�P�)�r���FL�h�l���(.��8�ՍB,I����Tg��F��"?a�� -kj�ɦ;Y�-:G$U�Sw�h��Z�<�
9[�F�s- �i�DG�`�ʔ��N k\�i H 6cv,)�?���I6 �`�CE�	�p�0o]\}��� |@�'s� HmAF=��(a�C�[�2�#�GK� քa���эѶ���C�g��D�����`�M��+; ���N����G����|�w�,O}��ښyM^-3A��}M��$G��x���ٷdU��r�/	�Z����]�
]
��uM\7��7�� Y_���$��^pPq�ˡ!<�		�l�����bI�x� b2#_u��L��4TX8��B��ug�@�Ka�T���ėD�n"|�Z�(G�^���d�"ԎFNX��h�����mD<�b͈'��
^tpk��~�N<��i���򘈕�2`��_4F�x�ݰ��'{�z�_ |�i j�=,� ��d��|~�:qm��
b��
�)�,�g"n�ܠt��35$\�GNQ��Y�S&�O�k#B��0>I4KH����!��[pP�ӉS�E������A�x�աF�9�*a�k	� �@ �6_~H���S�CԈ�
��)��!�:Q�"G@�g�<YWJR��� ��Z>�%�ã�p�6��𬌃nѶ�Q�� 84�A@wJ9������2��3�ߑ�O�1�!�W�Q 2��Y!K�� 8�)�'Z�H��:[�#���9g�H��b�&�4���^�#�|��FO�'�-Q�<=T�){��d�4)L ���!
\8s��h��OjB`��o+H�(�D� �FG��2���D�:z����d����%ǇW� ��cǠM?���� :(�\ۂ$�;�.z U}	�����6*G<��K" }Ni�G ��/	�p�2D��?�$r�O��T�^��P��A3�(��X��!�� m��6�3�!�:0c���-|�����<b4�3��J7��$k�� �K��7l��a�']�p1ň�1���A�ľS!��I�5eF�se�ё^P�DY��U�Gl��yF��?�N�3��͏ �H�4��`����C��T���0@�y�'��&�"9��B�ez���{�$�3>�P���F�36� �1��'EZ���U�}k�v.��c�h����_�b��`�ӳv�� f�[�� �j	�|a�E�0w��O��`��`/V�^}|%W���x�f=��֟�~��:R����;�v���'޸"��=��Q�0���@�O���#�gĜL� 2>���(
2�qA�I��~	Q4�Xm�anʱgB�A����U��'���̈���k��F�J�B�4 "(	W�B�'�Ω8u�4[$,��a�(���y���H�ĳǈ��]��J�P�ոp$���4ɍ��ǉ#S����#"���ˣ�i��I�t���J.ΐ5���	"���,#NH[g�ț��	=/��jO�cB
	h��T���r9��~B��䈅�Eg0wC� R�m��0
�a�n[xP%3���!�^�9�� ?Y�ΈG/�� �6ﶜ�5�uuĸj�fQY����'��!��W��"�i&`D3Q��y9 -�.��;���g �K�k<jP��g�
J�� {�BX�Nۦ(�FCF�	{�$�F(� ���S�_>�1�0\�W�����ȅ�cײe"CkF�!x�Sʚ	,�N�&�T��"@@0`���"��Scw$�ҬĊ-8{�k\�(�6'�X�'
�����6X��i^�%%>�
���6�ᣄ=Y��y1�B.��Q
�9F��剟��d�r��(CAnE��b�z��Ơ^�n�j�/���a&��Ɣc��HJK�*tl�{n|m��:A����$[�A��Y�ǆw�ڹIgh���Pc��M��n͹7Vj�KU��(�v���(F�'��}���7$�����:_$5�"�=c�v�ȁ�R4MiT����R�n&Z����p<i�$&T�R:	���D�d�l̐1�<����>"�Di���ut���X�xE{�Eڏ1�0kUiړ1���i��)0Q��h3ϋ�g��!xf���K}��c�@^D�,1�,\ c��D�
�=^ ��u�*��=K�|=8䓯Z�p�.�J��nP�R,]�n�G�����Xq)G0�U�/u�D�a��۵!Cj$�s�L�	��ۄ��'1T&D;�&�p8�NL�I�iy`�Ǚ9��
�hC5�Ҍ!�\�)f���/U� h��̻O�iQ0�?��b�b�Y�3�^uLx��!�Q	��E��<�O�U���]'?��ٙ�
;!�~�v"��o3�����kb)�g*����;A����jع$�j�[����ē)�F���PN���%�o4�G{R�$�2�c� �$T�1%��D*�
W�G�NI��o��Y�4|�ƥE~�vk����p�eCm]X��$��!�b���X�-�4p�u�38�"Nְkʜђ�h%X@ -�C��"�n	��8��8jj��
"J5=(U���M��v�<��žC6��"�Ǒ]}���ӧ��Z�\�dც-�pᥧ��9zְ�O_"��y�B>��A�AҊs`R`�a%�p?3X
b�4��V�Y���|�E��$'t�h�.�ma���'7^F�UHb�'Kxܹe�+x�D��@#��I��4����:�P���0IZ.�j��Aܶ=����B�qr�Q�"OjeA���3k{�q��KĿ��}��V����MN.�<b��|��X9�V��2�^$Y��vKc�<��eB�y�XY�dK[;T(�}d`�Z�<�`"�z+@h�pCU0�Ơ� ��Y�<�Ҩ�/v�����/Q.l���H�<P�r-	�D,��IG�<iA@�Wl|���K�|���s�HB�<q$���6��I�Bͷ<���	�A�@�<ᑇ�&�dX[�
ŭn�D�!D��w�<q�G�.	���_s�Z�ր �!��W��qBa.РOp�\*䚣f�!�4[ˌ��͏�lc� ���]�I�!�/(� �y�N�] Jl�Cӆ�!��<�8 [��B6kr4yK%?:s!�D�6�t�J��M�Fx��Zd=|�!�D� /�:Y�a�X�5��ё�bҎk�!�D��\��mK���/��P�ǀG��!�Đ�{��ZgKK�@�I�a�R�B�!�[3U��xSCȅd2�	�M+�!�ē-e����➂:&�� c��XR!�4j7��[u�ׁN���&�P�NK!�d�20Z��&��<!,��9��1}%!�DK%U <���I7�� 
��!�Ȯ@@�}�b)�6�IG ы�!�DN�!�<��A�q��=ˣ�_8�!�E�Y����k�/�~����@/0\!�� @�Q�b��f:�`�V�#�d�:r"OVx
"�W�8P��A$
��B�"O�d�7@�6�$��p@�)(��yI�"O"j�[�
C\1q�eE�3,Ƅ�#"O8��rG̺�J(1��(Lت�"O��a��ZK�	r��V"O��Qs�Z�iH��;ᎊ������"OP`��CI��` �����p��""O�9����xM��8��IH@��"Of�(���'K�L���>Ll��"O��� k�D\p�2o�2\��T�c"O�)ˑ��,����� u8"OXƂ3y�}�V�d���pw"Ot��"��,�.���悇3�R-2e"OD- � ,6�2�jM�d��iW"O�iY��[�����e��b�@%c�"O*�`�"	�<���H�u�2�I M0D��J���K�N9�$!�D����.D�l�)�>m���h��W�\�u�f�.D��򦇆3R%��#Ӭ@����(D����J����	�.Z�63��y��*D�l�P���d���O����Հ(D���V�B�#�d�ch���P��+D���E�٢oLH�𧋓w�Qa4k(D��yA�+L��a�N�[nT�@�+D�p����/Q���t��7]�*e�"D��X�␤7 ΑbaC�+!Ԉx��>D��Y���9U|����N(z���'8D���F�k,@:���x�#D��j��X-�R�Q&�E�_�v�� c>D��t�ǯCü��
�2v��{�L6D�@�b�˜ZJ=xG&�� m� D5D�xc$�ŖKLh��eB_56�lx�E0D��y�hO�x�(��$[�@�f���b0D�P93@W6DV�y� k�\64 @�#D�0ic��v��՚�IوU��%�>D�S���LDU�a@T�bb�y� 6D���T�E *���b�߆8F,�e4D��2C�=6�4���]�[y4x�B�5D��@ ��F�*��Z�7(U�*7D�8En��N�H�*YQ:B%;�9D�X�I�%)���xA�>"jM�盕9�T��/^I�S��?iįA�;E�Go�p��8�%�TZ�<٣�SV�ntZ�ŏzQ��k�<qu�F�w\�4�7�'gP���z�.����	$�l�ߓxI�tqR�rcV���d�C�t�p�&�!p�Fer��F��y��"t�����X�G��b�� ���'��p���t�ށ3��?�'l��T�`׺1�H��磅2�� �ȓ��E�ÔN<�%�鎩{��Aj���/U�.lѤc��`����Q�}&��q�˺N�n��VFG�5&�٦�1��	AA�-w:���],rQN��`�ӳ���R��N^��z��E

�:9�牍`��MA���%i
�"�g�/�`�?A�It1����	�o�:���1wd:T!�)�R+L�!w�
,	
�YfOL� �
L� h~��� �Q�d�Z�X���'N�*S�N����6=�`i��
�~Uq�Ώ�RJ��"O �� u���l�>�ҥ�D'��d�=h��K�o�����H}�']ي�'��xS�[�Ckl���O$����8�OPC�ř?Ԉ��PGS�T�b�*�_X�����~"�a�P�М���5<O��R�'u��l��W�$�:����I�g�X�ɔ&ܠ4�"��Ŋ,	6f�+�:
�+�`I���R7�qT���'��x��$�n �aIB Ie����7k�]���"�:8꤆ۙܵƃL�d�0��~z�ǋ"LS*�صLZ�eX�h�4
C��y��	�<��%�$IY��*�vL�0 ��~U`L��L�C?.��*��q�QiSr�	 O�����V�V&�x�ˊ�#'������  �,��N?� ��Б�W�0 ^�� �4�h2��t`a�B��m��x CPMX��z���Wv�z��A5��ka�.ړ:���)�K�Z�@�	@�L!a�@h�#�5�]YC�6'�E�v�Y$D�Fd�B�P�t3�eP��0>�f��HM����`�3\"&H��Vӟ����H:��ՂC��v	��a�MG������2^&.X�Q��c��O	S���	*l�~���)R�<v(��( 
W	Z!:�mH�Y�g�<|�,át��-��0I��0��((*7��7�Q0�D�μc�˜���L��DT�4�A8�m�fx�H����#�֍����9+|����{��}����)��������g�Z� �� o@	?&b�a0)�	�L��y�c��>u�rD�
�=!�L�nuH� ����F�y��E��慉�c"�i3pF��Ԉ�� �bW�r��۴n��c!Ȟ�0=!R��4��za��4< X����R�A��<�y��P�� [�h�)2��"�O��96ЩT]
�g�0�j��C�,U��p�'B���"�p�A�R�N�M�d/)=֌����-3��}�����l�� �'ҰGX�]* ��tK�b�?�d�Q&�_��,���_��>�j�IH� �ny0�l٘����&қ!���	�f��А%��6��0�vO��A�"�1F��KS1O =3�j�$$a��2eט2�
�p�I=J�B�鈛b�p��FM+E5>��,�(
sD�@� f��,٧�������Zty� ש\̚u��ɐ!V�ź�P�WP")�0�:"|��$[�8����S�~T�K�&Y����IQ]8��$w�)"%�&k��*Į:uh�ە� (r\�C��R|h�J��
�H��h7����q����a@����ɡ�N�	�B`@�*���d��^�o:���HqH��C�6i��sWN�*5�������ٌN|Rlq��S+���i�*n���(hח�2հ��$����&�G�`Q	� ��jB�(�	�M�v�9�!��$�D��΍�Znh�=�u�S�Yg�I���Ⱥ�d�Lט\	,]�%����e��������Q�ڼ�h@�Xx$P@�X[�� s0�L"��겪K�j���"�O]�D"�)*�� Q�N..�ЖK-⅒BJ
a���A��2�5�ԝUްݹ��n$\aÈ	�y �W���K��) UH)2f�P�����>c]�J�e�#a I����U��$��(#RXj�B���y�MJi�h��Za0иr����p?�չ�����u�IB�!��Mp�����Oz,��0'ڦQ���'�)��=�T'Ӌ
z�u:�D0P��9ʒ]&)r�A�%�3둟�*5�@�(u�s�9)6x�!W�٫T�ܹC�A�&BAVmǑ"���w�<[p���Df��{rMʬjD(����Sc�^��ю3���7Lr��Q��y�`��Kے��P��'�*�h�ۧ�@�?�*�g�VGL��t�&.g^p���2D�@D��$zHeK�_r�ls҂C[1Rg�5C���i�0(5x$�S��/��g?���9���5AO-	.$��� d"�p�B�'^��;�K��8�����9!Ѵ��w#��TE���CϚ.�V�k��Z)z:�U1��K>���z �z�}
5��Ĝzt��t�Ov��D}"�Pi7@6�N���<)ϗ�68b�՜dǠmr�����	I�'���D�1�웥"a4�H��'����V��2,���,�R!`�'�8󒮜�xʈ�R��؁����ƎI0*��1�ǌ-W˞9@��O`�MC�����`'E�ѐ
�'��֑�~�8u��w�h+��Ѩ/Ar-iPMV
V2�)[��� 
����p�%ԏh��YˁLi��D�QX�%K% T�-Z�1��
3�O�=��
��E��Cv��6��`�p�Hh���6�K:e��% chN�	j�}�4�߽hܠ�+�j�1��\�?q�A�z�)0��^Dy��C�o�'��|hU��}���g��@�r�8"k�SA��xq	��@��q0�	)��\!Q�
	��a��� ����0\@�=aV��;B��(K�W=4�"$]�e<��[D�L1#�f�;C�����2L��yBDU-yn~)��"V�Љ@&B��a���r6XC�I <��Z�D�	� yRT�]7
�N9��!�)bD����ɐ&�y�m�?����j�)Q�C
�I�0u�i0؍u����#H2}�Iӎ'�O�Y*��F�\��Ӧ��wR8��ˆ�/1��cR�d�PI`n˅2_|���yC4�(W� �L8��nV�[{���%OF�[�D�8b	�hO0��%��o)n���װV3P� 2�B8^�pM�%�ҡu�N���V*�p��� �]]0!"��E�:h-��	��H��� �;�f�h�!����z���W|�8q�>�t�wG��M�@��-���;i�^�)�|8�#&�-=!~+!1D��H�憄<�5�FD�y�"i�dpt�1㛱DcHD��4 �
֕74&��d�ج��/��&���;\ܸQ��"̚	4L�hŦ�Nل�I
L���1Z�,�8\y��%=zȪp�#.�|��C�y�cG�/�z��j���&`0 ��;w�O
���A��
�A�f3.KP"s剠3� �A���9Q�ֱ+@F-z���N�6+_�Y}��@��L�
%T<8��Uk��ۥ�ی5Ja|��́W�
]�D��6�T�P��:^I�HUH�NޞEkq�T.YX��%��S�y�ԭٴ�D�*�D:�y��|���S��v��ap�̤�y�d]�;�H`�n׳/rt�d
�AF�1��.�!�t�7BƵN��!i�$];�@XRN�1{$j@Ӕ꜓Ŀ�3FU��bv@O�q��hx4����=��N�C�\��7��|��dP�<k<H�ł�7�� ���ZD����aR8(C��l��H�e�)� ��V�ɢO�Ճ��(?G���d��H�8�~̓��C�x���جVs���ci�ݸ���JO�T- I�SA�.e�r��)��TR�B2�Or��0gF�%�F�a'D�x�X�@$���zpp ŝqM.��m��C�l���Ǉ �P�!W����?�X\�,����!׮�l��"O�T��N�(s3��rl��\P��&�B�rWJ(!ŀ́q�D7)�����p:��z��	��Fd��'�~m�s�Ι-��2�+�k����AE~=8��Sd�ɲ�'��y�仲��5W�xp۔�_�O��|�稁=,�`%m�4J�乳t��&��Ob�bь�Ik:|��g����Q��D�]X܈��#�aiacA�:�n0��L�Z>V7�ı;�D�	�J]$]R>]�JQ�+�P0��D��p?�E��9
8Z�kC턓+�^�r��N+^���PCT=0�\�IĪa����� �7�$IL-L1Cguޙ�T)���>��0"����34����ՅH	ZQ	�ĞsA,�AB��{�N}�� Օ����-�ૄ
B& ��0���:%���R�OޕI�ΐ& %����$K7%D����'BLQ�+�kA��q��87�ܱ�7H���N�����M�.Ѱ ��x���1	�~V�]��S���������xV���B�qӾq�ѭU�g�ʓ1=�Aۦ!F5R�=��_���XSC]6jvHe X��yB	�S���i�"��i(�)4�T�'Ɇ�J[^���s��<F����a$��1�F�qQ���Y�4���`�B�b��OV)1LD�]=2�̻]��3cN3m�3oK��܆�ɾ�|��R��J@�D8��,>ͳ����> ���D?���޼;�Xh%��'&b8 ��G���S�@?	@K��&�B�3��|���Y��Ja�'n�!��	tA���r��:��`Q�`W�V��yӡև@���5��1��� �0tApT�\<�,Hl.L��E}bLH�k��rE����h�c�8�?��n��T�5!PH� 7��K���l� �
����8�O�p+��ŭF�l[��<$]PA��6lR�r��'Q$DH5�H<�d�`�)g�j���R���J��F�BVh��z\>6͓�~&J������W��z�?�"�.Y9D����D,|pe)��D��>9�H���X��K��F�.C�ŏ=�@�r��� Y$i�0��|��+]x,)���@�0 +0�:�l��U����Ѽ�U�AKL�4j�9��%ړ��+��ƸaZ|�jcŌ�\yԝ�kA�B���8�BW�J���2��<�"�cr�� fq�diܭ7I����'�џ ��b%>)�����I�fST��d��OB@���	,	���ƥT:I�-�4��; ��h�9eTZ��сI)Hl!%��1ڲ�����-F1V%B�NP��B�I0
��M��D͘j�����К�0�@�YBưɖ.�
nD�!,�1	��U���h���&������FD�2B�ă��ݴP�����ݵS�����6�,%HL�	  Z('LL��/�3��Qx�o��*�Ƀk7�u F>�Z��xePg6vH���/Ah���U<�hO�H1��Ѐ�v+���Ce��B�Y�o��6�|��0� f_����m�t���z����p�Śhx�XW�A&+��h�!p����BH���$-�� � w��SQd$s��I��OK��2I9��*Q(l�9ql�[�y�'�Z�cBoZ�5	����a���Jh��$��{󠟉
H�)a�_���i��1O��7�L
@�����9+�#��'��I��^!/*��7JU�CX,��̐�Ze����ѽ�\�!t�E�^���$X��;W�!g�*,#��&Lߑ��`�`߸�5��Ӆd����O�hD��Foy�� �.���|�	�'��[ď��Q����C�$b��+ODQ`�'ˏY�1OQ>���f�C�\x�l��$�R��U�*D�P��/����vb�	�| A�&D�Q�jY2-�Pxp���.a9-'D���p�W�n=�C��B$9C'&6D���2�ў;_<	��a�	<�Ȉ!�D#D���	�$B@�2UƄ�7��M�� D�|�g�ŵ1�N�� �NY!)(D��ˑ� ��x�i@��'C�ĉb�:D�4����0�Ɛ�1�G!Y`�]P27D���0
�E�5��Ł?��m��e+D���k�	O�\��G�t��-@��*D���RI4a��m
��^�uߨ��fg2D�LxV��12�:A:��߸r^�����1D�x�v�M)r�YS@��71��\�1D��)1e�f�(0�[nצ�QAk;D�ت�$J36�&Xh��U"#,b���E8D��!߾ ��d�J��
Z:�d�3D�(�׏�%�xu����SLl3�1D�0r��L��x9�)w�*B�5D��A$�	��L���V�鹢�6D�Ԣ`��!]�2�A��JyTe1S�4D�� �}[��׺fM�,��n�ޝi�"OdL���PK
��mKT�0�	�"O�,�Q@Ԯ8�0����W
6��]��"O.	�f��g�D)ʧ˞F�^-�V"Ov��eI/p�q 	�q���"Oj�cd��@�(	���˘��Q�"Oе'N�7�P��2!������"O.A�CE�*G���A�`h!r�"O�֪-p�|X�O�w=d41"O�`�Ga��z�����(} �H�R"OFL��˟�0�6h!��H�C�Jy�a"OX�Y!�M.�Ƅг-S�3����"O�Y� ��#����	�4x����"O|����T\�Q�#�-�F�"O�(����p�lUKA܉f�=�4�'���X��0l��PjV���t �Zb��(��A^by`-M<Y���<����<�~`�F�xG�a�L�`�Pz�J}��H3d�S/O��`�(��,S)�i�:d��`�nѳB�4��Ƈ?c!ͩSfݏF�=0�Lo~�;����ul���%�;!6|A�%�&m��X��V8i^ �r��$]�l���D�~��3F�.�{@+��v�D��JGA��5kD�B=��b�m�v@$>��}r�-u>qC��8�Ly�IɗQl��B�i)��&ι$R\|Z�?�)�S�c:t�R%�'7�8�Gh}���'Ol<y�MC��P�O�dzp�0k,$��e�ɯtU����L���_�b�"|:���(���ʐ�š��$���G�c����V�0L<�����Mc�L��ɣ�,ْA�v��af��6�ʐ�k�|��N�O;���3f2��M�#L1�T`�U�A�3s�;Aa����������3T)ٟ/��'�(�w�2?>\p��'9>�8��+�(\(=1��#^�p��'�A�R��}nO�>q�Ŭ܅�����$���۲�xӚ�����P9��&�"�bؔ+�J�S`�Q<F�)S�G�1*�I�Ҍ�|�I�0|�a׷s_hT�R��8.^0���Ity3O�dlZ4y���ԟ��P�1EuBT�`Q�|�Z�´��XܓR�Re�Yw�o]�OH�����'ÒUSG���,d9pѠD��d]�`�l�K����Ev��t�7:7z�b��'��5H����&7���O��O���=pL� V-�t"���D��r�1O��

m�y�v�N8`Jҙ���R��¥�=ad�)�b9;q��2� �x�,��> ^�Q6�a��A$�3v�F�|�$�|��M X�N���J��'�����&X�� �Ȕ
�yb�ގq��i�O��5��J/N��M�aoLhz�C�����d�=1M�5�ٴ��g�xQĉ�ф��b�^Xa�>\����b���� E՝z���3sc.�܇�_��Xx�T�>���s��o8�Շȓ4�x� Ua� j�:h��K�"������u�F�1,�`',�����ȓ!'6�3�� 5B�����`d.����mĊ�[%,ҽs�ƭ��^I8���ȓXa�y�#�ɤ
�h!��Ŏ�w����T+vQ4c�!Xorœ���GÐ8�ȓT�)c1�^.x�q�K�'�|��R����W.�_�i�
� ~	:1�ȓв%!��鬜��>fb���V".)�eBh퀉)t��qy�̄�A�z�A�#E�K����t�5(g���ȓ54�m���ED�b5�l��M7F�ȓ$�����J�_��J��,qS`��ȓt0<��@_{�^���
=p+݄�P���AG�|ì��E��5uD�����Fa �*��J�j�k�����l؆�j'� ��E2E�T���HǪ",���k�~U���("
�����*c��ȓ���aS� o���(?��i��.[����ѳ2H���3��ۂ�R|�<Qwa���Yk-Y��w�<��c�N�ܸ���Z.^�~�L�o�<� B�uGڵ"���*D�[�s6�y "OQ����2�8�Q$)��#5<��"OL�i���0\�����Ȓf1~H�"O����]?�B���'�s	�Pd"O8!�3�s�T݉���@�"�"O���RΜ sКG�3��*�"O��b�!]�D��	��=�B�3�"O�˒�Ch$@��J�Y�R�b�"O�e*Lg�-IWn��N�X,
7'�V�<���D�b���" ��} @"�Y�<y�B=EU�Qc6ŏ�f�y���MY�<I���a0�c��,	f��3H�Y�<�t��~�2\Y`�G�X��0#*S�<�&-�) \�e��䈼=4B���B�O�<	ĥϪ;����2� �H�D��L�<�GL#l#�Qw�U|~X��T�<)�P�$T"3���{����[P�<����*G[��UI����5I�<��4x��l@�I�FuP4���[�<AcmT�G�츒p���j�lБ$�X�<��o�6�$�B�n]�J�IP7@@Y�<��*\4B1���K�@9�x��]�<	�LȡI<�-R�:��#��B�<�&ݼ�9K���^d`���T�<����2������N�J%9�#�@�<�G�.c��3��A}��7�{�<�g�B���Xk������%Uz�<�b�U�W��]�F��	G@���v��u�<�-��*���1��*"��GBo�<��M��YՐ}�we��w��-�4Oo�<��<J�Ľ �L@�BO�Q�GgG�<Y��(O�4�d�_r$9s����<�7H�*}Ю��% X=m{�$D��x�<��S�_ƺ�g�R9��tз��t�<�Љ(r����J��k}u���UH�<��ə� d\���ܹ+p$��#lPO�<gS�,X�9w�U��.�Bās�<)D�ȹY��P�̓?zc�=*�Eo�<Ʌ��
.�����<<O�Ui`��i�<qS�ǿ|x�A/?�0Y�ɛg�<)���\HzD�@o��C	z�pB��c�<��gA� �t�@�D%�V�@���f�<��o�'�x pɇ�C�*�pr�	f�<aS#z��̐�dT�?Dʔ(�͏^�<����:Dmr�_�Q��v�b�<��L�yP�1E��(M2ɣƏD�<9�"�"P��|5N]�}�Ī@@�<)��� �D�z� �k�4d�x�<GFܻ��h ����|���u�<�cH�'�䴉�琀(��y�h�s�<�� ��wc��Q揚�Y<�I� �Kn�<A�$M�� �/D2ǲ!qFcn�<�"����S�(^��f�p'�CR�<�`�U�v`����8�`�W�<i�,�K�Q�cٱJ�yv$Ck�<i��(\	#�_+c�����@�<Iퟆ$� ��І2&���{���<I��ھ"�Z�����-.s���(�_�<)�,JN(9��C��&�;�A[�<YU�+��+ք��_��I֨[�<ya�L05������Wdr���Z�<�gךW%R�e �PiR��U�<Yǡ�z��$2 Սn|��p�!�P�<y��nH����
GT�[�J�<� 0̰��G��-� �6W�!�"O�E�$� �)���x�,:8ǘ1��"O���ᇣ|s|q�6��bj��"OJb�%�b��P3D���Hi��"O(���DR����_T<�"O�P���
��Tz��@
AF��r�"O�)��Q#M�ڵ-e�]�V-�y,ȽB��m����Je(�K.�y���+��Q�R�߰_x����C_��y���TI��HW�� ̹�ĝ�y��9	-��`4�W�ޱ@����y��OJ�a��C�mu6 #B-���yR�ǐG�p�X��s@� b�"�y�+&��Y��Di�"��p��$�y"@Z::���r��]\h� H�\�y�X�9N\��«r�ͱp��4�y��?����r�O8Zb� �V;�y2bS'zHeZ��ܜT��hZ����yB�غ
KD8Q!��t[fa�y䌫A|���[���}�����y��R���u��P!+��8ym�ȓ*8xqu��e/P�DdY98S�q��#&7�,БR��$#��ȓT��� �I�,6�,(����>��������d��J��dQp��4o��@�ȓ���HS�"0����6;L�ȓ@[ܴb�˄���X�e�2�H�ȓb��!�Q��<`e�:f*<t�ȓ*�|����׳L�+���~;�y��"O�{ծ�5v��a��v��E"O�	���&(�ё�!'�ʨ�"O�<�P��>g���ț\�z�S�"Oɋ�"�ș��DT��X*�"O�����p]�����8p�"OMzf(Qr�x�F�߉S���j�"O����ɷ
M�EK��H!�6��"O�@���T4=�K�H?#s!1�"OV)�֨���	@F�a�b�2g"O�1b�����5���FǨ�c�"OHt;���'O~T�a���1���bd"O�!��Kǜ��Y��ŋ�rM:�"O�9a�ihY�|����"O��A�P`5	�-}����C"O�qPi�'o���xqm�t���("O�Aѵ`��>��6l�2g���"O������
7�q"�Z@H\pe"O�r%�Y5B��c��>*|Ő"O��R�j̚9~�h�HJ�DrQʲ"O�1�����j�a���=e�%qt"O���Yq��� �w4l@`"O�;��ҭga��)*�`�"O6�`d�ݢX�PtFE�͈"O�$:Aa�%y�4;��G:u�,̚�"O=�Ć����k�(׀h�4�t"O�`�s�_�>Ջ򇂍A�|���"Ov��H�9�.�a�%*H�(|( "O������gxlx��" �|1�"O4y"��#�F]� " Cdm &"O�-0�Á��Й�V�4*��[�"O(e�fśl�*�:��Ѷp���Kc"Ob����W�6�V�#�APB���t"O6ْ�^&o�~A����2����@"Or��fc�
� 6��=]��8�"O�R�E��2����a!��J!�R"O� ��K�� -.��A���Q�����"O��rkS:9����a�/�*)�a"O.\[Vɏ&$�i�cm�^��, g"O���E�*VZ�m 6L�0|�p"O�T;FÌ�d�E��
 i��"O��{�n�	�0S0
�5o ځ"O(j�(�=�l�f��M��1�"On�v�ш	�H�r�M�X�1�"O
uY�e��0Ad�0��T`R"O�Y���<��i*�#9?���"O��J�^r�����j��"O�����I�i��x���m�(�z�"O���w� 9b8B�C�/�/�F��U"O� 0�2���s�¤fdD���"O0��Gd��@���'B�7aX��A�"O�Ic��EYc�E�L3Cr`��B"O!2�J�@��h��/whR"O�zRcV�4ȲQ!�!�� �TE�b"O�(A�M K|�!H�`�j��XQ"Ol4��D�I�HP �ϗd�,��"O�#7�ZSJ�h3�m�4W�R1��"O��[���K{V�!g�<��xb�"O�a{�ѼQ�l��H�:LN�ؠ�'~$M�C��\Hy���!9li�'�x�g�~"X�xC��HL��9�'͊�S�G�&.o�,�"
��A�]��'�l�@��
|�V�����%��`2�'hh����:�@������'۶1G([�w��yf+в�R��'
P�H�a�,9;\HsAL���r�'w�`�Q�P�d��E��H��'3~��ȑc�}��*�?�~-P�'�2��e'�8������Z����'���ad��
EF���ƌ�(�.���'}������Sn�
�D��!~<aq�'7�i;��*&q|�� hڱ��}b�'�4!K���1{�aӇ��I:�Ȱ�'D!	� ��.�
isb(�':Y ��'�z��^'H��`����{R���	�'9���䖼=��Pb�ݸ(@(@	�'�t,�G��DH�y�����V���' nA��L �R��ؘ��^y��J�'3�p����3KF {�ŉfP����'�ȕ� � x�$�b��YP�d��'�.m�  ���   K    �  N   �+  �6  �A  �L  �W  Lb  Rl  �v  ��  ��  ��  ��  T�  ��  ܩ  �  a�  ��  ��  ,�  l�  ��  ��  +�  o�  ��  ��  *�   � � , � %& f- �3 �9 @?  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,��	�<���� Wnb���,;0�iG�L�<!��2TZ�,�!ÓK?n(J!i�p�<�v�a������ObT�Yi�<i�#M!>\��	��vD��&�e~R�)�'+�����9V��ɫ%�$��,�ȓ ���,�@��1�n=�4�=������� ��2C��
n�����-�y�띯2T��Ga�kU88�^��y�m���`'MZ%i�h��O
�O�7��O8�?片r+ �)tN4T����҈eO��l�`(<I-�4*ڕQA�H���pе��H�<�f���vFP���Ӥ;�ȍ���H�<��K��]P����� )�à�D?��'ea|"�šX?����-,[�pq�ƭ�y�+���j*f�J4���`���(O����6,�x&����E(0���!�X%�F�A6�X��ѱ�
:b!�G���m�hٷ35�-��O��d9}�>%>Op-���K����ڰL�\O.	h�"O����"M�N\�a�M:���g����Ip���O��ؙFj��l��}zp��$K�������Z�ɻh.�b��$@��x��|�4�=��4�M�~&�Z#V�i,���b�Äw=����+ғ��OH�$6Q��p���e� 	�1 �!�$��>AQ�)�� �2x
7I
�ui!�Dʌ~��l��DZ�i0p����\�_]џ�͓�?ٷ��$�A�*�� A!���Rj!+%�X.��'�ў�O�<)*�,C�
�h��l��AŪI-On�'w�S��4e� ��V.���v�˧n��5#���Z��� ��>�X� ���("$[D.
\�I~J~�'���I?��a��V<.R��P�u;ZB�ɑyx(��A�Q����Fo�y�P�D9ғ-��	[�'!"��YЃ;=��(�c�0U����In�7�*̙��X�Qz! ��O2kg,��'�ў"}�1����R$��y�N��7E�j�<A#bWj�D��g�"%:)`�_�<�#J��0t𘅈NZ4N�C�B�<��.R�R�>��蘕 �R(:E�A�<a�XNA��p�� ����Xx�8�OHE�� �7I�]Jd��x������'�'7]��Y� ����)B����WfmDyB�|���م@�&A�vD][@���C�<AFk,W�Dc���;Ã[���0=��BB��v�Ki��Ni������'21O$�>ҁ�����y��6WL�L�ψl�<1eNΊ�(}��i�7Q4\��C�i����<i%#�������NU;���ҫ�e�<��.�b1A�](�(��dP_�<��MD�0�RD+�Nł1��a�s�<�r�[rZ��%��;�%zs�Px�'�ax���Lh0Ze�.)�f-�Vd�y�x&����Z"<t@�V!��CC��$�"T�U���6�d\���Y�tt!�8D
�C�+�I�p�HC�<!�d]�y����A%,p�أ�a��	��'��f�)�Sd)�9�@�'�؄Tm�<!�B�ɰs��£B1v�X�ޥ;n
�G{��9O�3GE,Jֆ��W�ON��y�"O6E��O>s�p0�kʾi¸��"O���pR��$���@�hxJ��'�1Ojl�!��� �pi@�K�(�i�"O�IIcD4<O���6�J�"4R���L����޿D � �'K!D`�Q�
�xU!�ĕ&l]��# Jp�q�.�5ў����''��$#7A�t �ؓkT�B䉃v�IIŅב8'V�Ӑ�W�(��B䉺1��JF�#S(�����(E�B��*s�9HBD��y4���©W�B�I1N���봈�6
�!�$c����c�DD{J|R�Y;����բ��wǢ��F�v�<�q%�T�@D����1 2@��
��hO?牠K|H��Neb��+�$L)�B������lI]��EC �X���ٍа?�¦�) K����Y������aZI�<��-�3k�n�j����N�ea�H�'L?}���a6L,�3�s)��aVK!D�`�
4�0 ��#M`��}�5�3��ȟ"�R�+��tI��K����U�Ʃ+d&Ra������^2; X���ႠԐA�/ي��?A�'�R1�S��S��:"	�e���P�'�a}��'?�@f���OPTqQ�GP9c������W��y2�'Z�O�}�vOL�Ѕn؄-�̑��d-�@�8�[�jA,x*�Z����Pq�'(�"=E���C i�Uꌻw�ĨSf��y��E�=WԠ�eS�rz�A�%�T�ў"~��c
I�@�%C�!�l��۫�yb/N/}�x��b�X�O�H���J��y�'��	���Ii��-@�^T)�%H�,I`����O�p�ܣE��#ب|�5K�Qgxd�ȓX�
�c�J/VG��ׯQ�.8
M��|B8��Bn�>6�.��oT.�R-��e}�T�V�%aO��3���EKt]��S�? �u����C��3Djb�*�i��	U̓��O��q׉ȢsU��P�bK�Q���'���U^t~L�3�ƎP�X� NŶ?SZ�mZW�`�>AD��q`����$>8%;���z�x$���^�$pT�Q�#Aq��K:�ɈG�Q���Ip���0�������$wR`T"Opi���M8��sǨDxO��V"Ox\{�S�<�ۓ�I@�XIVO|�D�s���0&oxy��)�D+4w!�ۇP3������1��PW�</b�'�O�Fy��
3������3�*��E��?��'���Bc̕�x0r��%,V�t�SL��D{��tCC!c0\�J .TeVQ@����O�"~��'ƦK�;��>��L+�T���=�ҍ��Y��(��M�,�J�J���R<���0I��r�g2?�:L�0�ȩb@�ń�d���q�Y,E)��I�W��
���$��3��@��l	�0�
���G�ӈs����b6*��]yt/�i��C�ɳT������Ɖ&m�i���R)��C䉤S��u�u�2ur�k�D9.},C�BF�p���>vȦh8��Ĩ+�FB䉇)��|�%AO4*o� �"CDgxB�IP��A3��P�&1`�:@��!YRB�	/]�R�@��լ�(ؠ��"
xNB�'-1X�Y�����`�b3FB�I����'T `Cë�<SOB�ɤp�J]���V�ah�Yゎ� �B�	�{�V ��L����@�qYB�	*J�T�I�.*	�v�R���l�>B�ɔ3��]R����feh�����*p0B�I7A&�=�1�޵7hl�3FT�I�4C�	%dt�q���''Ȅ���LAC�	�:2j�j�O�6B0(RS���ߘC�	��� ���.	�0q�2�l����M�W�d�`���=�ą W*��!�@���B�.Y�`�����e�!򤂈��ṕ,�,H%���u�+l�!�d��pcZ,(��c���st*S�])!��@�6��A@A�B���QU#[1�!�߹Lڔ�{�C(G����Aũ�!��.zvL �+�.)�fmb��I�!���2'޹�q'�)���[Ǧ�,t�!�L;xQR#��y����wDՃd�!�dE��^��Ղ���B�Cf�.V�!�$����Q��!~r�D�gB�Yz!��a	�9�a+_96�,��Vg�\!�� � �8sk�%z�EдJ� 
!��a���5m�ka�%�X=]�!�ì6�h��Fn}/�Lq�\>y�!�ъ��`�Gm �~%������!�D�t����B�{�ʼ��!��P�!�مZ�@�91�>�dxjs�G5�!���?po�����Պ}����PK@ [�!�DX��Q)���X������!@�!�$I�*���ӯ����fN��!�D&N��OP.q�>�*��!��s\ ���@$�D�4.S�b�!�ڲ~8�*0b� R
�=˵�a!�$#�.E�$Ɲ.`ඥi �¸_�!�d��5VeQ�eG�j�$|�F
��L!��YQRѰ�1��u��i�)B�!�D�N��b`�֋n�������
�!�D��OL�as����
\`h�@�!�� d=y����]^���I�pm��ۡ"O�5�W�X�z_X���ZZh�s"O��rdA�k����3�ONj��"O*X[�C]O�J��0�˸�6T2G"O*\SFB��F�D�y�bC�3�,�pv�'"��'I2�'R�'��'�23�֑���W�M�J�I�}�!5�'ob�'?��'��'���'��'mܭ�3�O)�j�y'�ˇEҪa��'2�'(2�'=��'���'�"�'
��%.C�)���1g(�B�1W�'���'���'�B�'���'���'����E���)�=�E���Y��'�"�'���'�r�'���'�B�'��Z�$��x"h��F:h"d����'d2�'���'rb�'�'~��'�$�dՌ��O�V}�1��'3��'���'��'�b�'��'.� �p��A�F�ms���"�G�?A���?��?Y���?q���?���?1�D q��z�T�_����䎾�?���?!��?���?����?I���?��剠$��芒G}d�JAc��?���?Y��?����?9��?���?��NȌ���5
��hߘ���n՞�?����?Q���?Q���?q���?����?��f9��HH�i��`����H�?��?���?	��?����?���?i���CwɦD�� Ɬ$0y����?����?a��?����?)�i�"�'U�����_RD�r@�#Ht�8�q��<����󙟀��4\�!��Lطw6��3c�P��NpA�S~�s�T��s� ߴ���uh��D�2�W2��0	��i��&@�f��r�OZ1A�.��zO?!���ʊv?���L�P�B�ёo&�ݟ�'*�>�X�DݼIuDU⁊[�@x�TK���
�M6��i���OB6=�%�U)��Z]�(3F�
�4��5Ah���fӌ�	J}���+R	w��Ȣ�'�U1Wʘ�o�P�`�MJd�P�'��ـ�Mިp@��i>��I<�2؂"�'[T��bjVm���IAyҒ|�Ah�\�*��D��_O��X�I�#l���� C&�V�<��O�l�"�M��'s���Wv( ��+ٍM�����s���x�$l��z�Z��|z�,��y���8�{?����dY�H����U�ޔ�/O���?E��'ʚЩL�\�H�P�ʫ<�'ܶ6M�4�I��M��O0V='��fT�xQîG<I$�9�'B7��զ��I*	lFpS��(?��#ܝ�|��ʋ8p�KRɚ2���P,Y�N�Hs��#�N�Ñ=Ѻ�����>c�h��l��;Ԭ�8�.\�Z9��򤎭4D���e��J�̸a�#4�Y��������Z
� �n֔m�܉p�Ȇ=hs^\�t����6~�T3��J=z�b��T*ަ{z��#C'O�EF��+��^�*wh�*���iS;Ѣ� �V�l��Is�� �ީ��ս'p��J��"M���Ѵ`��s����AR�X�qr�C	���ޫ(L��A�(YϨP�5c��o�؉+CN�*X]�}��Ə�.y�#�	�fA[�W�@*�{ֲi�"�'���O\�\Q�S%m ����R�9bB�lZ]y"A]��O�2}/�($!��R���;Z��a&R�MC �KZ���'���'<��,+��Ox!���ܡ�����HXA�hH�NAܦ��ua_s��|�<���e�P��hY.4��q�b��9Ô숔�i�V��q���`y�V�$��d?�#$)��:f�M�v�:Ԉ$e#�1O����m��ܟ��I� ����yo0���
�`Du�j���M��*Jn`!$�xr�'�B�|Zc�
ES*���|�8��Pl�&D��O�$�5��O����O@ʓ��P�Ǐ$�r|Kp�M0^�n���ǖ��O���"���<��P�3����瑎!�����	GHny�<y���?1���?�Pv���3�r]¦�N�9�>��0ȉ /�I��i��	ܟ@%���Iܟ��$�]1 F�6M&���@2G�.A*��L,"��IЯO����O �d�<i�&<��O|��ah��}Й��([�!%Az��$$�d�<��M�[�m�ͨ@ㆠ��y��,۲x4�n��T����`�I�=Y.���͟�������S�;�0�d���a�.��"��5;��N<���?�qkЀ`���<�O��2F#N� �I��� >SJe{ߴ��J���m����I�Ob�)_~RG�1e&�i��E>����ǿ�M3.Oj)�%�)��LC����I�(',���P�*�6,r:n�$�O �$�O����O���|�Ч�!p����ϔ�O0���$޼Nϛ����
d�y����O@��RL�L�Ƭ;gm\?T���m]ڦi��ڟ���H�MP۴�?���?y���?�;0�4Ճ1�"�Zq'X��>Qm�dy��5D��p���	埐���O6�+7g�
	��I�sEB% ������Ԧ����s갨�ܴ�?���?��}��a?)gꚿ;Z4�:#�*_��5�"A3��7����� ������	j��'�=s�Ӡ}��8B�j�²��3"��7?>7��O��d�O����g�dZ��I)&�&Y��$׾ c�0�� � (\ʀcz����͟���� �I~���N.46��*L�����i�AD�7Qt�\l���0�����ߟp�'��"]����a�4&~r|+S�G�e��)�T���>��?����?I���?	��
�;��F�'�r'G#��`��ş�[��:���v7��O����O���?�G�W�|�K����=.xbٹҗT��Iٴ$j�d�d�O`���Ol���!�Ҧ��	�����?�C2"��oE�J�U)>f�Ey�(��M{����O�E� ̽<!-O�� ����k�t$� �R��^���i:b�'��А)v�d�D�O������i�O�AÃ·'L��y�ɉ	Kn�p���b}R�'�P�`�'ɧ�d�~J5ʁR���PĎ
�� ]�'�Hɦ��A�^<�M���?9���J�S�@�'h�Rb�
�kZ��D��5�,�6fb�^m�25O8���O8��R�*���?	�/��p�
 �`/ �����M��?���� ��i���'���'�Zw������ͤ��+%��R�D9�ٴ�?�,O�8�>O����I����!Af��M.�rCǕ�d)��	ӟ��a	��M{��?)��?a�V?��R���قj��1Tt�(g 3Fܐ�'@
pқ'��IҟX�	d���'��|����d��s���m�\	I���u�4�?���?��\�xy�'���1���.��Tx�.�#�F�y �K�y�[������O���: h�6M\-\|\��� �>LըY��fV&��m�����Iퟌ������'�R��-��tB�$hd���'@_�J8�,�F�\6M�O��d�O����O��d-L�`�l��	Y!��҅��=<����p�գ$Wt�3޴�?1���?�+O���Џ��	�<IQĜ)�Vdy�)�L�&EP���h�2�s��?����?a!�>]����'�2�'��$$�!f��%�%F�vp��κXuT7�O^˓�?������$�<��i(1�^,7'HiѦ�C+��RGms�����ON�����ڦ-��ޟ����?����0��@A�`�H-��n�/�x�)�!K���D�O���`��O�O��-���޴a����h��rp�}��
��Msa�A�yݛF�'�B�'����O��'M�nX H<aɴFZJ�r��v��7En7m3L����3��՟��"B����Ui�=�0 Ά�M+��?���U*$�Ǿi��'��'�Zw?���#J�m~lS�O��/ �ͦ�'� #�"f��'�?��?�'��T�6��`D��+<,���F1W��'����g����OP��O~��O��D�O� [GΌ;N�4P�L�ɉ|���?9��?�����I�|��@���ź0��BEH 4�t�lZ�����ş������)�<�
�@91U�E�2�aՊ��K��	wa�<	+O\�D�O���OD�d
&=�Plکrj>H F�[������&L�F��4�?���?Y��?�(O��d�3 �)1��œFe���@4bb
��j�m����h�	-����Q��9nZԟ��I�xd"�͢k��,@ah �@���c�4�?���?�*O���^�T���O���S�\�8%+�l�2
0����m��G�n�2�O����OD�DI�k�(o������ʟ���d�� �!k�� @��cwU#�4�?�+OR��X�"|�I/�4���U7)g��{@	�v�n��쏨�M����?i�������'���'��4�O�"B
>Z�ܹ��D
�4�����C�I&���?i1�T��?	���4�~�OIȈ´lG�)��T�*R-��9
�4*-�Ѐ �i���'���O����'K��'�01���G�2�ЉMR&:�d���0&�O���<ͧ��'�?��C!׶��'o��!��0V�CH:���'���'d�0�&gӸ�$�O����O���� �d����=�'�L^J��PѸi��I�f�t�0�ig������?�dȗf���;eǈZ�$�SQ��.m���'Ӵ�b�G2��O���+�����sc�#���M��1��P06S���6�	ҟ���韈�'����Q�FW� ��M"�J��=�.Or�$�OZ�Op˓>i���##���
�����"�M̓�?Y��?9*O� 
��|ZEJֲ����(�ӎ�����Y}��'�r�|�\�,��>A��φcqt��ǌT�%����W}"�'/B�'��x�A�I|ڳ�7� �d`�ez�[��B�jH���'��'��5]Nb����$
Xn����{�|ኀ�q�����O��T��T����'L����<M�׬	�N��T�uA�#-O�˓4�Dx����	Sf���[�<�v 7�i`�I�^��Y:�4ms�ȟ������ |=����e�m3� ��r��_�`��:�S�s���:0�;(~-�N��E��TmZ&�ء;ڴ�?���?i�'D�'l�Fծ��y9��Zfq�����gb�6��P�"|"��B̰�R�F��b���G��	e	�ꀹiB�'��P�U�6O����O��	�'68��hМ7�0�����b��b�)�M>�	�D�������в[�P��1�E�K*�5��MK��(����D�x��'�R�|Zc6���s��*DE���RM�(kv
,��Odk0�$�O8���OD�tP\3ǣ{����4�
�fIQW����}B�'�'���u��Y�į�S%�e��	��'t, ��J3��ߟ���ß��'֎,� �r>�z4m�����Cg.K!,��v1���OV�O>�:?���'��L#6��y0 !�rF�5@�x��$�O2���OJ�P��|���$��6nA`�1d�GWєp��/L�Vl�7-�O��O��t����>��	�okq� MF nF��P�����̔']����,#�I�O��	��&�S�E�[�$qRl�
>P}$� �'g�!���T?iK2A�(K��i��F=E�49��g�$�b"���iT~��?��'o���3��ъc��'�X䪡I�H�h6ʹ<�'�G���Ox��z�u�Ƀ?4�(I#�4��,���i	��'�"�O�c��zFºA��	���@���R�C6�M[�Կ�����yr�'�� �9��֨Q��YPg�FP��z��i�"�'�S�O�$�ON��.P0y��FY�n.�Q��ؓS�x,�>ɕM�w��?����?����fӀ,	Y
Ff$�4�I�F؛��'u��Rí(��O����O<��� $[�{tL\��E0�l�(G}"�Ӿ9�'0r�'3��'T�S����8&Mɔ5%*�9r�c,� ����=�ē�?A���?�*O8ʓ �m�цF,�D	���,1�T̓�?A���?))O&AJ�L�|��]c��R+	/|=`�~}2�'I��'��xy����)��` 5���w���f�������<�I��8�'6	�q`"�%-����d�]!8�h�B�M�U�0�m�ڟ8'�d�' ��:�}BH	;`��qf��u��A�7	Q�M{��?Y+O��Y�Y]������S;�Бx'�&lZ�s�[�%��D�I<1(OX����~2�瘜HH4C�]�e�ElFΦ�'K�;Gs����O'��O�2�{d��80�إm���r�F�6���l�ty�B���O��x�r�)׍"�.Qq�a_�:�ȢĻiz Ñ�q�����O ���B4&�T��3L�VI��a�bn ��gοKP%Bݴo��Fx��)�Oa(��L�/��Pu�׵=�����������	,Qj�H<���?��'��XA&�*t�4�vj��X"�ٹ�}�)��'m��'cr-�8��`��!��#5V4��*�]��6��OT����J�����Iw�i��󴏇5^db8�s�31�~��r$�>��BK��?y��?i.O>���ݤq���2K̴	��Qa��. L@�>q�����DT�L���e�!?p�Q� Kk ��'��O��d�Olʓ^)R=؀6�Z�qAcI,��D�ٍ4SxY��x�'I�'Y�I�|��s_t�]+9[t(�B�vM�%�'���'��^�0�׀���ħ݊5c�$V� �LQ���](L[�!h��i�|�\��rEJ5���N0�Hh��)LJ5*�E���6��O ���<��#�$lj�O_��O�T�0���`��hGdҪq���P#�?�<�G�OA�����fY�|�䙱����ׄW%3���\�܋���MR_?����?�k�Or  K�oXƠ1�G2.J�d0��i�	(4P#<�~��ɑO�ð�քU�y����!�����M���?���R��x��'l�l���]���s�d_)��|�Tv����3�)§�?if(��-��4R�����q�ĿDv���'�B�'j�|��.���O��$��4Z�D
w��+�$�Ag/��$��b���I��(�	$�ض�W8PW�4��R�0f⑲�4�?)�"��'R�'eɧ5F��5>�������:\`��$��$R)8%1O����O"�Ģ<���[�2�pU�q��/��2(I�b�@kŚx2�'EҘ|"T���v�#t訩�╾-:�A3�̡v>�b��������Zy2�84o���l�,�ȑ�W�"۾%A�d�b3���?���?�)O��d�O��x�^?��e�6^�c��ڹ�6,bB�>���?���D[�"CP'>�8�%[;j �0&�Q�Д�n���M���?)*O���O�IIb�?�.�T���Ä\�т��W�~tl����By�/��zB\�����t�:�g�<њ-��b��f��:��ڦ��'��'���ɟ�i>7�M�n8� �#\�Nn��r�F�fK��]� G#;�Ms�T?��	�?Q8�O���
$�
���t���c��m7m�O� =�I�?Ox�R!�ߪn�:�0�ݥ8u�,���i�°!�'P�'��O��'�GB }\y
f�^��t1���9�6-݅ �P�"|��$���@ׂ�&p�����EN"XzA�i���'����L׮Ot���O���5�\	� í_�MXШR�o̪6�&��#U%>����|���T���7a����C�*��l런Ru�M'�ē�?i�����3�έO����`F�_Y�Բ1I�`}b��'22�W�����P�I^yB́�<�|��fRmK�t%�*P��"Al/���O.��:���O,�D�"W�Hl*��j`T��R�!h<�!�8O˓�?Y���?),O������|�&���( ��ޥ>)8�i���X}2�'�|"�'�Bm���y�I� �H��J�C�����r���?����?�(O���hE`�S� �y�V'�-KJ}�#%҂&�-�۴�?9M>Q��?9�ǘ*�?iH������'"�Y{�"Q�0��Iz�mlӰ���O^ʓ4��������'�����7u��Ѷ�&F��*�X�H��O2���O`Ӥ��O4�O�4��TH�@A�i.�XBր��l2�7�<�t�ñPǛ�»~Z����B����a��Y\�8�,A�N-SC�y�N���O�\1���OD�O��>5����*
N�)����/yӖъ�%ɦ��������?�8I<��?T������`�C�tZ.Q�@�iP��!�'Eɧ�>�d�&,J��@���8�l	���U�\&ԵnZ�T�	��A#��ē�?���~"ϒ��)AdH�Im������M#I>Q�!��<�O��'�2�Ŕ읚&')-wZ��䍪�N6��OܸZQ�k�	��<��g�i�A�`���p�Ac�S�,��<��M�.�dT�#���d�<����?���DM\�? ��S'"=p�`}	��
Jd�(FDM?	!�'�B�'�'�R�'W�� �[j@�ʢ�K�F]���/��rT�l�	��\��Qy��>6T�S9i��DT2N�z�!t!O��� ���O���ۉ.���Pl�Ex�e[�oLd9A�ݑ.�<�'���'��P�ܢ�e���ħ`���E	�>\_`��僓�?G\�%�i���|��'�"!��y��>Yg-��<.-8�K�\��KF�4Q`_I�R(���.*Cf���$Jإ1DN4D.4C�A_�fIJ�r��)9SRs�e�@,\�^�Iũ6�O�%���E,(�<��eBXＱZ®\�MP���R�Y(��կټ/��EK�F�&��D �J��=C�Y�e$�[��H\�51�T08�ԋeɟ�_�`�!�gW)\����M�R��YK�qj U�_&̸t���Z�K�I���) �d��g	Gs��UQ%�,,)�L����G�TؤO��j*�|!Т�O��d�O��̺[a*��E`�eiCiB"�z�B"��R�`P���đw��$I(&TQ��$�<sA����h ���Oc0E��fߤF��9��ɕ1\Z؊G ��X�"���Rܧ�Α��O ��+
�q2Ѡc-O75�*�PD�O��mi���i>]E{"A��9�X�8�HZ?_�<Hc�8�ybd�;�8)�K]�$$\U�ŏ��HE���T�'��R��ܸ�$B>m�p�� Q�����a5*��IΟ��	��Zw���'������2���C�S��cg�S�x�p���ïz/�tYb�W�BH�e!�ɇ,/��@ی��įw���D�1Ц#ŀOH���&�Fx�t9��_[�����"gn���L�'V̨#��<2:��+ՙZ�X��DU��?����hO��<Yc�N�5J>(��	̑4$�h���&D�0�b���v��IJG�^0'��	��%扏�MS���B�>�H��O��N���;���?La:�1'E�'��mY0�'�R2��h���׍]��
��-%.dk�+�=t��H��D��yeR���'45�ʣ?I��	C��)x���t�lt�ӆPf��#%�2��-�	�l�i���L�@�gcӠ��'�j�R4M�"�جX�p! Y�y��'%�yBi��،AC҇��(�pC�(H �x��`��p���J�Q�L��Ĝ�Sk�=��N�Oʓc`0�8��i`��'��S7f؅��/b���Hi��!؝C(��`����ԟ8#�� 4�NܓIU4T�� `��.lM
���u��D��K�r9A6��`�-�����I�]Dk�O�/�J��N۵�J1�.r����S�XI@��Y�?DJ�U\\�Od�(q4O*�O��Ui�Y�W�ά����}��D�"O,�r NаJ� Q��(o	H���"��|���I�]��Y���2u����`J�T<��4�?��?�
Ǒ������?��?ͻ_�����}5��p���*�b��W<���@�@<��
1D#��O�������<!�l	�*����-��E.���!�~4�)_�$�v<
rƂ3!�8<�}��hs���WGȵ*6�>.����4>��zM>�W�����>�OJ�X�	���rI�nj@p"O.����7^1�)[�c�8
\Z�X�8O��$@M�����|�8x�9c�� <�-��ao�)�%t���'/"�'b�ם������|j�"�.9��-)��<K$�P��Jx����ݐR�S8@��ŤD�/�) �T<���i7�k��e���\�D v|�	���?y�	��]뒢�A1RC\p��QE�b ��� ǅ)Eq4��<���Č2@�1nZ�����2.��� �؄	Mp@ĩ�3,�����͟�:s!�ş�	�|��Bղ����m���������|wO
C$%)��2D�����[�C�2ty��?�T �(��-<|�ބ��ń��6q�K�BI�fl0�����A!��]f�'v�ej��0n�'���[�) �>M� �ԥ:"���a�'�p4�A`ߛY��ͺ���?�"َ��4��|"r�iplxџ0Д�r(� ����Ր|bC��0��7��O8�ĩ|������,7�.�W�u��h� 6U�����OP�!d�fhu2&�5 �,D�[�B��a&�|+�n��吐��1�^��R��h���0Z����c���y�d�v�a�.�'O>�`#�=��ݹ`#��D)�ONM�3�'!ГO�ȳ�J��D1�rH\�f�e��"OP��	!��@bgPI�z	q�%��|���I�M�ޠ���������ZL�$��4�?����y�B�r�\���?����?ͻ.�h�A*V��,�6I
�D�Q���`y�pk�k��U���
�B��O�z@�B���<I��ƾe��!g#Q�7K��aaE�T9�x2���AZ��$̑9&����
H���'n����G):��d/Ɍ�6�z��:��ɍ���L>	u�\�h[ސ��.Z��>���A�<I5�A#i��X�AI�_��c@��<�
摞"|��M�
���r �?��"o0k���UF��?���?������O��m>�����k�	 A�6)��ksh��6��C�I�2���Di�D��RD�m|�Ո�I4���D� j`Ȗ��;9i ���\F�h'/�O����4	E�m[�+�� �D�ʒG߫@j�C�I*d���
�Tt4 tęI_�c����}��1l��6-�O�d �J0r5!�J�!��9��]�-�D�$�O|��c	�O��Dh>)XL˼	�u��@P�-� �W�D�=�-[&I���H�W�ŀw��`�¥�(R�Q��[�,�kEɛw�����������-G(~�y��@ɲ�1n^!aQ�Bf�O��%�4X��
kn��@���y�XX�!D�P�$`��7lQᧀ�'���@G"��hO�iۦ��Y�4��yp�I̖;~�ys�$Sy�ɧ0 ${ڴ�?�����I��	���D�B;P�����v�n�� m� J)���O���l�*:��EǤ�B4��/A�Aņ��K�|@�ץC�xʡ�1k��Ke!�6aP�B������!-�)i��e8f��;L\X �+�*꒴ڗ(ѝ!�BI�O�5i��'���O��Xjr��|7��(�
�, Ŝ1��"O�e󖈚&.!{C��-Q�ꑡ�a?��|ZQ�ɿUN}�ʦ!KrL3��{�ʔ3ٴ�?I��?���Յ!S�����?���?ͻ9��e�"hS�n�f}�sN0h|���P�X"����l���4V���O�*����C�<�#���
��YФ�%� �A!ʔ�D\��s���b�45� �!�vܧE�0��v��1��9Euޤ�_�j6ֵڱf���i2֥�)�3�Ă�.�zA�vl��h�`A�ElS��!�d�=����W@�ґ� L����D�O��Gz�O��'�$4���^6^��1��_�h�
���g�r�e�'���'o�~ݵ�I����')5¡�<qO<�!c	�3D��'D7vL��c��`uj�f�0C삤
��*�r��͈$hg�H���]�gH�I�g�:p���u�ĝR-���~y.��,ʓs�̬��i���i��t�������۟p�����P�< ��Q�$öhG����	{�}��� u	�.mǀ���!O��b�C�4��Y�"Tɖ�i�r�'¾5b�#���p���c�:S�'(�+E�"�'����5��X'�� T՛䔮s���2Ef�5[�<� ���N|����7d���6�I>[�����O�;d�ȑ@��Wm�!x�	w�xQd ؐb��p��@�S��`9�Ȅ
ro^�$�|�H�O��$�T�coB�I�X%��g�e"w�!D�L��H�_���xr�M�r鮉У,��hO�M�=;gce6r�X��
�c�p��s�I��q���|����I�0+�����X~�:���<$FvH%Aް`6����O��ZA�ښb28�
'':|h[�/�%'��1�g�|J�F;4�zS�iT�V�U��'&�������͊1$&ʣ!X7mC�� ���ۢ1��֝%}�.��4&&Y$T$��
��A� �'�N�@�[���k?�'�R��\4o^�ۄHZ-5���q�E;��x�#�3F!���<�*�`�19:ў�S��HO��*Ր���ǅӍM�S覍�	���ɯVt�P���t��V�'���'h�"T�w�؄)��&n|h8 ��6ܜ�zj�Ŧ]R���6%ba�G�\�O@��a�f��<�p����"Q�#aƵ %V�;�Z������{���à?۞=�3kѹ;��"��l3�2���E�_�x���Ρ>/�m�`��N�	�</����|��	�l��@ ��G�Y:�3a���yr�,T�`"��%�ص 1���y"�'m�#=�'��]����@��'%�� v��o�Z�+�H_�^�.q���?����?	P�����O��ӳJ)
+A���-��HGd|���t.ܱ$�`�Sh��C�}Ѕ��G�'�L��w)��\�R�ʳTߴ�y�n�3O��}���� Bp��U '�џ@
�F�q,�`��d��c���%� �h�d�f؟`9%j�$0JĹ���G�H-<�ʶ�7D�4)�=TJ�h�EV�41Ju�D�Ԧ5&����D,�M;��?��mò5��l�T�̠q�X�Ī���?����xB���?ٞO�B�8H�)C��l�'���E�������W<Pq�"��/v�1z�A�%K�џ�9G��`L`@ �E�e����v :^�Q��ҪM��#Q��]w�F2�2�?I �xȲ,��%�1FΝ2)l�{s ʻ�yr&_Z;|E��`��%`V�pS���x��`Ә���o�y7 \�iǒ}@�(X�)�Dރba�,l�џ��	L��O,=F�)�$n��K��T��=�&ڄ9���'��d+&�]�}�l����|}*��˧D+�2�`� ����]~�$i��,}���5l�1�j�
tE2��F�1��E	�B��%�Da�Ab�2Q��,A�c���	�g�.��B�)���^�| "���H��a��u�<B�	�Z�xI°�]����#�F�(���y�'.Ψ��O�4G�l9ʣFI�zΖ G�l���$�O��D�e��͂%O�O"�D�OT�4�<U�f��(���R��E�(.�;Fb<Z������S*�$3��)�<�Si�	{����B�06��H���\0��-�F��b�n�J5�(�S/u���1]�H� G	[�K��&gѮD�F8��4���'��YT�����$�O� ^	� �#�=)Ņ/B���<4�D�fc��Kc�u9�V�"��u8?��	�?1�	Ty2.G�5R&o��Wq�<���Q��H�.�5g���'o��']��������|Zы�']e(4�%.�M���Qh�(M���UĊ�b���`��+�������
�JQU��J�
\�d/L��F�x��t:6l�LN>Z�\Z��)�Q`��8է�<hɄ����-#�ؘ��̟T�����iE(���^S����'+D���DC�70�q���6G�h`�'�I�M�H>a������'h�	5w���#�M �h(�����'`�hsq�'��;�ZtBA��-館��ꏆ鞘�T*��5
���c����!@X��j�S �]��(OV��s�:U@Ӧ֚��@�ˬ;��y� S�z�FdK	r�@�!ʓp������GL<iĬ�1�2��EY�H�ȓ6��ֆ�����&Ֆ�Dm�� ɛ�ר�ꝓ#��,���"��&J~�'4�|���i���d�Oʧf8�A��Z��m��aL�N^�L���%N�|����?i���M�%ϟ� ���"N�@�d���)V4���E� h�: �a�2s�"���9@�N�u��P���]%-�lr��4BN�E�,aa�G܊XBe�'8��'9꼂�Arɧ�Ok�������X���A�ɉR�hQQ�'�
�Y��
$�p-����8FZ~�cÓ/�����7ؾx���@�Kú|I�|��Fڙ�M���?q����&(1�?����?�Ӽ�V��%I2L�Ҥxb��h�2[��i����%T��c�Ωˎ�T�x�B�;O��8
�l��	����G�)A�9�	»`�6�CΕ�}�	�����xR��$�t-�J��{�FC7��5-}~�OHCw�����W����j�	Ħ��'�F3x�⌆ȓR/��ѩ�"&v���\,P��u�'��#=�'��u�z�#ռOb��"?�ҭ�C4K�����?���?����&��O���(H�Fբe���,�d�^�� �	Bj�ZX����j��|�6����܁Ŏ��f剼ZZ̵:B�ԥ3����1�Ūg�q��1#
��;��(��0{�^>��JA剪d8��ej܏(-^l�����Y�$5��O����I.Ժq ��+s��KVLP4|m�B䉢72F˴�&=���j�m̂d�b�(��4���ވ�2�ir�'=j��Ĉ�0��!�-@�d�����l G�p�I០̧o[��'C �q(���I�i����"KU
جXI GG[�,0�"ܖ��s'�߮��#�b_`�����-�|���A�-8$ÄnY1h�\�jҤ^q�@�"DN2z��O����'��6m�٦]�	+Pf��W�B8t�|����.ϸA�'����+C�T q�27���I �PFB�I��M#D��*<����	u�ıq����?).Oб ��m��$�O�ʧXR �K�f��U�E�+ ����,  �A
���?�Bh�a�R�ps�5Z�h�x��6��	)fʜ���Ǉm�ĸ��#�Xjͪ㄀ ����;^B�$ ",ɜ[�`,���on�i� �?�0AW1?^�0��3u��g�+}"@Z��?���?!����Os��t��>9� ���I��<1��yb�'��y�%�V`0� �T"�!]?�0<IA��>R�h�gd�<�d����=z\�+ݴ�?��?���/���h��?����?�;1` �Z ��	�֤S6ȇ��N�� D�6>R����4N�T�HB��3c1��EA��y�IB�AF�{�eG�!Q�Qp*Ӟ3�da�g�#w3�fㄾ
AfA�擟�ħO{@���`�e8a,¸qu�]�#�E2�ִ!0�J2�M�A�i�r���5��,Or�$I�,k0���V=ay�gI�IA�B㉎\r�цP~�2@8��Qp�T�_����W/Cğ�'~�P��K�rt<�	�
M3V���x�)Gr�V�W�'���'�"�k����柴�'?
%
�H�qdm�B�ӟ8����,C&t��)tC��X�E����2����,�c�|!�8s��zVbщq9�TK!Fӓt��s"1WI�%!���(&�� �J
S�O�����޻o�i�&F��b#�Ż N^�z^�8�O�I��į<'��s��P�q�"On�a֍N�7"%��Y00�����D�Ϧ-$�HzE������O촩�3)R��Z�a�)���;�J�O
�� 2H~���O��ӧ Ԑ�#0�t	R�L�:X��MV]�iS3G8VL}��c��h@1l&ʓ=����e`J'C�����_xa�Iۏq<���u&�v�>�Q4l�٦�Z�h
`��sf�B�}��!�'~ZpygKȶKt.Hz�LF��	Y�y��'��y�Γ�c�b��[$JKH1��B��Oܢ=�'
a��cۼ8I��ZDÄ;A`��v�#2:�R�,��W�Mϧ�?I(�V<���O*ȚA%�,r^T��ɀ��O��䇑���A�Lx�L�L� ��R�*<y�j.�J��鉙j�h��",�$Ԓ	�f�>����-$�"Yޠ�"��ā]������ލ���dR4�
�T����ꙭ0<�'�NM� ��!�'�jg�! ���B �tU����)��x
� ��$O�6�R-X��ۦo<�)�G ��|���ɭf�r$�s��*�R����O�<�ߴ�?����?���������?9��?�%��,���N	Oh��A�3��Y���2�$<Y�a\�dv�8��֟#.b>I�4p���~R
�;���	���aJ�rd��$犣vZx��FR�
��(hT�'�M#� j��Ӑ��\֍ၧ�����dl�������)�3���@�����D�F�P�1l!��G2�`����EC!��x$��H��I4�HO��>�K��#��LF<hb�$,�n��P"����d�O0���O� ���?	���4�N�g����f��?�8"�! �X�Z���_ L�"�E�>Uِ���.x��]1�������rE��C����������͒7c���Jw�'P\dP��ަ`��\Y��ʬ��2 !�?q��'
�H�,	�f�)�L7_��X��'"B��l��^���mXhؘ�0�y2�'�	�L����ٴ�?y�d$�Xt�Sx��i�
�,<L����?�RGC��?������/��x��H7�eY��H���Q%&�a��&�@��	x�	��W�.��4���!B���6ޙ8Jdl:GhC�&�
��Х7^ 9�@�	�$���˦m�۴�?��Y	:�(,�c�7W�>)�^9���O�"|Z!cʊHT�3Mܘ�$�q�'Ux<�ּixTMr���t�aX¬S.@cV�C��'��I#e-ڥQY.��D�O�˧e_1��j��閧ri@U
��Q�]Y�����?���Y��uI�R08}j �b��:J@ѫ '�����H���Z3�34� �� ��;��D��[�	�,���"eE��9A���'P4���%�n==R�^I@��Otz��'���O�`m"2BT![C�0R�g5�:���"O��+��1R&MУ�ϓ�f���0��|r��	���u�MF8(�� ���~�fX@ش�?!���?��+�X}�Q����?A���?�;٬��e+ڈX�MH���
��O�g�FY��'~Q�3@H��������C�}}���`ű�]�D@��S]0@�@ϫ;��À��[kq� ��O<�s4A˘M��]�3t�-HQ�{�it����|�bOU�d�K�E vD>lcpC���yL�@�"���5u�r����d�i����[e��xNda'�!N�H�Dݛ7���P��Ot���O��D�������?�O,:�J�m�z *%KAE��Yf�PW���/I9`���Fō^֑��Z�'}�H��Û3�>�2�a�iH֬�C�Hv�9�͞� :����c�#*9f��g�C@�'r8`F"#sv$�{B�/V���g���?q�����?�����'~LX�0��A&���pOv�Z�)�A��'��j��Jr� c�$�U��И'�p7��O$�O� \k��i�R�'z丘��֡`�t���Ʃe+���'��	�]��'`�I�V?���v��4WDά�%�cI0��A�W�L�s����DX����",��L ��DV�L B��,���xgE9,�^��*�n��LɤL�
hX��SHȅ΂�����ȹY��j=�d��G��р��K19,�%�!&!�d¥M����&3�:8;1.U�vj��F{�O��6͘-L(��(`)ޗki�����c?��OЄ���BΦ5�	��H�O��t���'�����gNG�pz"f8Y��ja�'R�ɼvP��.K3$�j����}���saA�#n��S XG�#N���p�N!)�$�'B�8 a�u4P�!"'�0�z�c$���d�OcȈ�ˋ0s�����'F���H� ��O��'��?�BP�\Ì��N@<a�N;D�ԚBg� ֺHF�H<F���S���l���T�?��T=j��0D����
:�r1��i�B�'b^�,�h�[d�'k2�'0�we�@�����Y0֠H�F��`ሔiΛ6I�!<2@��Aa�b>թ��Vu�6X-����@O#-��i0��T#2�i��e�h,,�뱯�p�J���+oD*i�O]��ռ�Ro�x��a`D���H�����Ó	$��'�����S�g�I1Q��X�ЉQ/C)�[���8�BB�#4�d`���;E�<@3��z�h��ǟD���4��O\�R�k��%�mja"U%tp�#J�\�ʜ{"�On���O��$�亓���?��O>��3!߫s�����.]O���C��+xl12D�8�M"DE�B�Q!"B6�(O��r�%�Z+XmzE/D�B���D�2&Zr�:_)U�d0*�W�KH��#�1`X-V�*���0`���`���|G�P���-~�����'R"���E�F��zǤN4o�8ds��V	a|��|b��A  u��O�Ar(�[B����'��7�.��n�.�o�ߟ����#0�ૄ�œ~��#��J�#a��	����CB�������|�ve���'�XZ6[,�(P#��6*����"N*O�D��d�:6+8�q�Ă�8�jӅ@(K�xrFA�?�Úx�ϝ,%-z�#U��6Y 5sq菔�y�hl���Rg�6l$���AZ�xn!���� ƈJƋ_�8hx�I��Y�(�@q��H*�Dlڟ��IF����yi�ڱu-kb���3tšpU���'ƐPYP�'V1O�3?��	F5w�,��6��ք�;���d��ʶ���?ѠB����B���#�"/����B0}�#G �?�Ɨ|�����	�x0bV0��������y�͑If�@�ۣ&@)�Z��0<���I3��4M!��T�LMhh|9�4�?����?��D܎~p%���?����?ͻs�J@��#�?v�BMYa�&C��T1�/JZP�|��h��.T�Y���C�O1>�_w3�-|ǌD���IW�T���a�:���*D�v�z��'cϯ9�|�c��I�A��x�XRKP�`�`���~-�d�*/��})�t�)�3�$�2A��99�탠i�VY�W�'l!�d^� �pub@��5g<��$ލl	���OT�Dz�Op�'0���JZ$#���)TD�\�xYTME7N-�'(��'�kz�m��ȟtΧ6����Xǒ���ʽ,�΄�cíT�0�v�P)lج���M�5�6�.ʓC�4�BC� J�"B�A�R�k@�5X�� �6eAd�9���'�Ą�E(ʓ,^�L�Q�� q,��#G wgص����՟���� ��!fC�4�Hp�U��z��ȓ!��x�/ @>���>`3� �<�q�i��'�N��A�|Ӗ��O��s�G�Z$��� ���p���O���E'u	f��O
��'66�t*�F<��q��&�iR���IÆ8A'�ߢVM­���?�,���	�I�N89D��>d?9�T�$%�٣@�J>�]�SdОNXl��ަ��t��P��dS^�8�&��¯\j�a@��:X�C�	�T�dŁ�N�4IX `x�m@;�"<Q��4�&Ym�M�8�-����a����\َ�%��ʑ+�M����?	(�44��OM��j�(|��YNA7�$ű�%�O��$
r�����o�?����(�1I�Nh(�� �&�'�d��ղw:��!%蔦O`�iA�C:%�P��2j#��>��ɟ� ��H�B�h	i5��}#h�
d�>)�j�̟�M>�RoT�A����U���w}��J!-�U�<٠ß����=qY(�s����hO�	�Q�'�� i�8��"��?��˳�l�6���O��dȴo~�@�BJ�O(���O��4�v*�-�la��6|�<�@!�3HȜ6-�fTiїo��-�<�|�tI����	�\�h���
�+�'Ò�Z�ٗƀ�|~��$�n4(�*Q��fh0Љ/�du����y�/\�� ���+S���w�	[���O�7���S���B"R<���ҕ��2i%b�ȓN9>���ȱ� ��)
��5��?)��i>Y$�XvÏn�����<`8Ѡ�݆8DxdB�
���$�	��,�I	�u��'B6�l�����HR��e��Y��y0�UG�}�5�E�Q�6I�+:3�5[��)X�Q���K7t{�i�/�@�x���� �qs�Ƙ#�,�x��"A��m�r�J$Kxp�O�r`�H	�bq��ON{��⃯ԔRb26�O�d��]�;L�11�L%|_�p���'`�'�ެÐ��@�F���2{��0�ya���OR8��IB���'(��c�Ȉr�L�Fk�5R֝� �'!򧁭b�"�'b�	�F�+���=pw&M�Aץ
�L�	�L�'Kbl���m1R�	:�j� �F�Ï���H�U��9pv@��M��x=K����G��ؘ2��PYʰ��A��#�J<A'����OD0Ag�'�6-�]}���+"d	��ŋ#�XT���['��{b֚����/>�ڇ Q/�O�=�'o���*�mU8��Gd1^�`{�b���P�tk3�X�M{���?�(�������ON	�!�f8�����V9݈��O�Or���ݶŐ≄%h����c]�SMfiёl����':RZ5[ ����:���6��Y�O�q��L��LK¥3�2Th�\�Dd�<Ģ͟���b�8OXB1�/̍q̰�S�>	BH�Ο��t�SY��/WD8x�2
m��"�E��zc�4�	mx�bhƔC��Y s��w�X���Tq����
/ғJsb�	F�E%A���+�-�0EQ����?���6����(��4yB�¯C�`��V�|�
�S���(wf�^B�I� *���a�	w�@������B�Iv�m{g	K5:���C��x|�B�I;2�>P��H�MDp(�'��T��C�IOJvX@�ˑdS4��c��;H�C�I�$�V�RE�'�l��p��nN<B�ɢ0^�-*���&��2q4B�I�P�pK�CC5'��1�V�<��C��SG�h5)L�}[ą�c)�H�C�ɸQ�L�f/���nH����m@4B�)� ���+K�D]i�Bҥi��@�"O�i���3I'�4*ġH�a�(��d"OB@8�FƆ��8!C�fs*yk�"Odٙ����|� �!s`�+����U"O�As�ǔ;>����R Z�	:�b�"Ov�j���|C4�	$�U�=!V���"OF�) "I���pCݬ����"OekR!�	b���E8�L�F"O|-�U��'�Hٹ��G�y$AQ�"O��2`���f��e�_�n�"O�(X4L �*f ���m��Wd���"Ov�u�n��! ���5��
6D������� ��҉��t2��Z�N2D��p��X=b�r��i�#6���/D�(����;W"]����q����%0D�$�ШT�{4�jݦ'�����#.D�08tgЇV����ۃD��Z�F*D� 	���M���JFت'
XQ��C+D��T�I742i����h�zU�3�&D���d��z���a<#Ziq�>D��𵇔E�y���)|��t�CL��*�����SƠC"�^��GB6}��Q�~D���ɳ`$kQH�*}s-�0�QgX<لV�V���dD#ZbN�{�	?�t�E/�X*�X	C`P�?Q �!N��Ztx&��%F�Aܓh���дd@-;R��5�����@0�B#=�f�>Vh<j@쒨=���8)!��"B^
u�$��k��r�h���D� #R]�X;qOR��I�]�$��B��e2�%�'���*�L�n޴��C�P�8y�4��3�ԩ��@���O$\sQ�*W�ܽk�k�Z��p:�2Ofi)p�^1!�\P�]�*���B��O"����o�U����~3�:q�	�}~� �"̦1�p���c5 �`��	2i�@L[�ޘNw�qB �=�֓O�p@$n�ؠ�!W35�a$��tD~8J�Ɛ-z�r4QW�Iq8��g$@)'~x\�wgHi�bM�ă
�.X
Uǔ|?D��'�$��<�E������D��c�,��aC�(A�Mb�������HOD��\�0/  (���?yH\�\Pe�3�ʛfr ��d�L@�걎Z����e.bܓ���d+4a�bD�5T
��I�<��;�f�	 }�&HΒ;~�6mQ+�N�r��/��Z��x���s��>S���D��e���ϓaN�� 0�T�K��%�.V����	'2��(lv�0e�g`\F{R�!$�)�vn���e�K:-�B*��N�����E�}�.��P�?��=.�	���'��F0��hT�
�EA@�4Đ^�rj�K��$
�e�"'�:�
�2����ӊ\�{��h� ��s��+�|�(�S�V-rf�J Bի��N[�雦kF=N�#=q4�dizt+��M>t�>gc.Q B �j*:u8L��-v�ųJѭR�VEU���',��5ƶ�3�7
I���23P�͔w���KC���+F�YmZ��z��tC��8��s]�1T�ݴ7P��IG���k��X�%�i��-��� f���2"׶Lm���H<q�mT�-�i�ɂ�%A��=9Gj�9Z&��" �P���Χ�y�mL`R�C�%x_j|;Cb����1
p��5͔�%h + ��U%4��Z�D�� Ǔx�PY��fE#��lYv���d�m���_�G�DP(aĆ�M3��,�Ҩ��'�J�d�s�����Ō[�謘pCP�;Fz�h��/xp�dʐ�#�VM�% Ρ�y�ϻu�>�Cŗ*(c�͂w�Βlu��>Y��S��|��6�8G�-�Ro�۟�h� C9G9~}p��Z����q�k�e*� ןoN�]�Tc?W�n}���O~|r���O��Bg�Y�+���P��mL��@�yH�����,,�q��
�s^�-G{�%g��8D��x�&ٚF�/��0s�1�w���Tg
�^yphb�N-0#tH���]�����a&�x"ɋhv���"-�����*�u�7^8Eb�$"�S�'P�b�$$��1KQ��=O��� ٧ �H#=�Bb��>	���҉ƾg	��x��Cp}a�.�nE3�^#4�������D<��8Oܘ܈$f���4r�M�7F�"��Ƌ%G��¡���bQ�ǉB5\����X���'\�|Ġ ��*80�z�{�� �oN�!�E�V��`ЌBBl���� �R��)�n2"kZ��3/0�T^�1:"bS=N�\�A�G�N�B���c�qOd�=��<N�u,^�\�@����Ɨ[� ���0@;�ĩ��'�n� t:�ܱA���$Z��u� ��!.�>����i�^"=�"GO��u����weʐB�ዲM�М�aK�$�HO$`�R�˛r�H���MɆ��ܲ�U���%�>\ڈ�8����u��r��>�B,5�m�����L�T���/��P��$ٰ���h@.+'�j�X�m��WԛV��3S���`�G�U+���S��M�ס�.l��X�q��9U��S'�?�����'�(ͫ�9T���O&-H2��	flu�`�7F� �31d¢d�ȝ�'��00A�����3ʧf�jP�%-S w����CH�j���R2p˓\��Z��� ���b�~��\�d��i
���c�8<�V���B�Uy�n>Abr�@N:�0��O2h�*�$�*�)� 0�f�]טy��/	�p\�'�j�ʵ];ء����0:�u�`����дa%�z�Sܧ!�t�����Oh+ѩܫJl�qc/�,3^9�Ʒi�:�yQ�]�{��$�aΛ'V�� *O�,tH�b@K��y�7e��"ЊQ���O�YpQ��iK��R�R�.�:�@5�ɔQB@��	|��*򧘾|�dM[-4��ؿ"z�L�	ç��Xz��������P1�r(�堚�g�J)IǓW���ɥ0��	@�)	�Q=: `t��=8�T]�&� 4�Qѫ`yr)x>az
ǆ���7d�9�����o+�?�0<	�kS�	
\����<a���'B�؊4>b����#W�"��&L����q%N۟y�rT֧�O�^�64��0�B�D�a@ݨ�/K���+S�iܨ�*7(�[u�dPKW?E�ܴ0WzA��@^o)D:�.�4<�Xw���~"���7�h��2��$����r&��uk@pK���*���Q�8�Y�K��Q����~���̐�Ъ�$S	E9��� '�J��TI�
��x���,�J���V=��%@=A���x܀;��%�fkɊ�(O�i[�:ڀ1� \���I�;wF��'�R�i(���X����� ��{�@؉�
F���O����⃇�!L���v�K��1�,O�1�go˵+�,8(�A�O�YÃ��~(�k��5=O����4+��4�?�)��M葡�d�PS�׶&z�P��	ʤ^��Q�=� �>��BTU�A8�OЃ
^lp��[l}2ҙ>U�]Hf�+�o�2N �`*7��K��tӐ��S�ψ�p<���Z�',�d�	V�P*!/�O�ѳD�c�a{b�:�ؕ'9�!�� m(>u���Dd"Lڌ�d\���)ӓ\Ҝ��%�P�����*�#A��O����@����t=��D�9n������-9���{�i��)3�ły�S��MD��=�r�c7�"GA.�S�?� ُ{B�/�g}R��U=4�ڢ �� �z�0�Y��d�6E���Ы��pO��E{���7|+��ʑ�
�����
3�tXZ@�
�\)���eh8O�-�eażk5n��J};��?qR C0�]�c��؍��O'J|9��U�R!A,��(��ܱB�uis$�"mR��h��Iu�Cf�H�8��;����U_
&����M�<C�����͖F>��j��	
^x��Ӎ����h�J���U�r���j�=��V(����Q��@rV��S��M+�)�)!*��a�\4SP�Pukʿ�ћ�'d��x�J������O���B!F
E��a�Q# ]�gl��m�b��'8���
��I!�'"6l]�d��e:eq5�J%o��"f�ƅƬ�R
Ǔk��X2�Ha�4e���,���k�/+G�H`�0m�$A=⬖',����M���sI�z�hX*A��	��"=a����� �Q:�,����d}���rl�������ռE���u!�Y�<,���<�}r���9~��Q�?tR�{f�\�h'!�V�,*���^�2O����TSj`y�M����)�;E3�%0a@��~�&y��:J��$�)CrD��0�S�8�PГ΍�Ykў[�lF�C�\�rFԙ3�R�9�nG�Nf�:(O��I!���0|��ã{��5��c��R, t��, �8=��'M�p<I����3�Γ�w��|"�V�{4U�d�?�<hy �Rx`��'|ḧ́�Ӎ`��ɺ���fb֥W�#
�H#=�@�V�(d\��AqkR��Łe}2�θW���⣟'t�(4�!LT�^�yQ�K�o��x@�RS}��K��`=󎃊J<%�ٮs���Io�1��V���=�!�q��|i�,�S��MӶ��$k��ؒ��68t��G�\-;�Lp�'���7��"gB��O��;6/J7k���k��&PX9	vcY�#s�u�<	rk)�S��	@Q<u*!�P/�,�6"�6O �S�C�R��xRkȨ`[<�,6JL�بv͈u��E4����4�S�'t"�� d��I�1b��M�9!L�YQ�S�&�r"=q�˓�@d�s�ͼP��*�!Ds}2��Q�%8bH[�O�v�0͝���8�I�G���ItĀ�zp��e�{,f��S5;�,��9U`���Aw��n�E�\�!�"]�0	 ���ָ'��5[ąq��Ւf��FBU$}R���7/�5�T/R*"葆ϊ�Ab£=��t��c��o�(�c%�V�i@�m"D�$*�SZ��
� �v*_�V����鐌5]ЩbU ��p<	 Ξ����n�� ���ܦ��Y�6���)�S�v/���� �2�*l"�k��9����B �� �_��6��1�Ѯܕ���6as�y�-O�aV��%�D��V�-B���@[�fC
�P�[(s���I-���
tN�*�,���G#S5�7M��Έ�P�%ð�j`���qOx�Iܴ<���L*�p)P&+�f���,�FeP�[�rIY�2�.ڞqF{B�=~y~�a��. aZ� v��,����'ړtȜ��}҇ìE�n�!�`���ܭ�b.�)I�8�X@�:2��x����p'$��9��X�oV�H� q �ۢ{�� <3�e�@�A?Dc�<�O����L{�? T���ʱ�2�ٰiQ��Z@P��*dJt��/�mڰ0O �=�4Q�H�ED��rE���z��o�
>�_�\���y�bRp�`���%y`����e�`XQՌ�K:��a�َ1�7�,k*�p�iY'1��8ٍ�d�����*"�1�խ ==�@qC�M�#�`�:������R���XA2�'�`���,1�0iD�i58mq�'��O��&$^��ɨVSj�h��It��B��m� A*�~��"C�g�|"�y(���3�z�����9�
�9!+@v;Ĵڦ�O ��H>Q�6�I��?��B_.�.��_� '�I�[�T����H�'��� s�'@�SAҥ�>�
I�,���Q�n��X��Ɯ��$�F���K��]~���E�C�b�2@P���&sgcr�Έ�MC`
�T�`�\2����A�&�*�'�z���իl�@hϋ*����'.^��  �^U;�e��=tl���d��?��k�E�t��0�DM�y�V��HPܓ>����I>A�.���ɍWP��W�/(T}��֦c��z�Y�?��x�C����4*��
޷Y�� �'�-,\��ϰ!/��O\�K�g̓m���ϦK�PZK�a��"��%c�"=ѓh�7�(,���Q�pe|���Q}�92�$)�#�0`���# �?!�C�"��',��Dq���lO�X� Yb��PVr9�G$��v2����NC(�,�lZz�e��F�|��h��'!������<Ʌ$[-H
2�j!'ºI��*��C{?Q�9O��J&�F9%���@��D�'�H�1'��^���Ǩ� �蕙�'���@H�m�I0
t���dF&]�'�V?pL�l)��
�i�l�Jbl�<Bj��k�䱥3���J��i����U
�b�q%�'+���|"*M�?c��s��A+��	F%�6��D����HՐ��	<;��P��]Ѥ �y���%�@��\`E"ǯW�#F�,I��i�΀��)a�	�~Zw���Q昱i��e�`��2Fo��e�H�xt�<���r��!��Kz��ONTE�X��c�,C��L�ȼxC%�
>�XL�ȓ^���B��C�"�T� !	V�\�Z��Y(	[b��q$N��Q���!b;D�8P����sD�a3ƨ�	A �*O��lI��\i���X-��`V"ONXaSA�,����a

�W��z�"O@���ΰpϰ��P�@�<��lC0"O���C/�XhEcՕϮ0��"OpP�E�^�2�:���� �����"O���ȍ%�\�;�/�1H�!"�"OƔ�vDB<#��`1a�_�z��H�"O�rq��\��� #������"O��Ef�qﶴ�d���^�.��b"O�ty�m��^��t����8����"O��Z���
 ���r@)��"�"OЭ�`H�c���b�U�U��0�"O~$s�	��%`�%X%�,� "O��ī�%U]\IZ�EE$�Bq�"O� �B��10��5�$�ӄ�d�҅"O�²	A*N4�ط�_�G�`�Yp"O���@Jç`D�h��  g�.i9�"O`ɠw	�N�⤀��W�M����q"O�����C(���ׁ��J��1�`"O��2�H	���2 Ù���"OL�i�O+��ᴯ�$mx�5"O��Z�I�Rc�|����d˸��"O�)��m��%yD�e�ޙ� "O�Ő`J��>m�E �VR֌�"O��v̣a&���c
�6ɴ8Ѣ"O^e*��>c�,,X!��!-^��S�"Oča�8z�H���(0+h��'"OJ(�v�!8��$�ѧ�_�D���"O�ѳ��s��ƨ-ؤ�12"O݋V�h��1!R�	%B^, *�"O�A�C�0Y
��ύ(B� �"O����Gɖ�V<�&�I�^;dle"O.��]��r�'O?{��t8�"O����¿).��;��̰]����"OBdr�$�99��VAEv:�л`"O� J$�; �I%��Q#���"O�ݒ�è>$��@�M:Fz��@"O 51�*,���%��X��"O�u���-=F�T��݀S"O����FM��,蓠i���X�"O���"�4Sf$PU`�24/8qC�"O��C`�F�X�8�˔N_���f��C�<��&�m^x� D�:*��A��d�<y�ό��x	4�I�|�J1��d�<a�A�GX���>JW���L�]�<1�ˠ���3mL3*��(�V�<�U��J��@2��V�oKxт2**D�<�bEU�9v�ٹ��Ԕ�����*D��-`z1����$sQ,�)7!�IoS�
�e�3H!n���(Je!�$ħgɫ"-� {���P�!�dS"j��z� �_֍�����S�!�7X��`�$��h4��r`U�!���4(���?����Яc�!�f�Aap��ꩱ��!D�!�dR=66�[6�ڂh������x�!�58p�*�'Ì9nRP��M�o�!�D6`����Z$GPz	��A�L2!�DO�*�\EkPb��f1�=�F �7�!���lM��([=X���-:m�!��+A$�TP2c��|�� �)�!�D�
~�@֥�/}�V����~E!�Ev�d`VnZ�>ɴP ֏�-!�dē0�p�@�G	�~A"0�1qO"��$������aV��:\a����a{��xb�i��j��ܽN�<��M��nB}��'�����ɡe����&	B&�@J�'�찡�W�js���EM��n3<|��'��#��ϖe�$Q!E�+n����'��A�#��ҭP$�ȱkqa��'W����֙	Z�Q�%�JP��8���'\�؛�K�l��)3�D�)(&V��'��2+_�Hi^d#ae�*�^��'zܱ��8of�{�B^��2AI��d�O|�Gz�eA<7P$�"���.F�be�V0e]!�ZR5��	F�'H���Q3B��Y!�d_�N�܀��"Qn�"��zW!��ԛS6�I�倦g��5�`�DV�'�a|�6W:��F�܉:�������p<����[{��� *8B�y��!�^Ą��&uR�/�,r�e�g��=B�D{b�Om���7	[�V۞1S�F�3K e��'�L��ãȝɦx҉��,	�Q�ד��'�&�iR,�;i�����c\34.��ߓ��'c�����"c�P�q��D^�e��O���9�)�'[x,\!ba$B��Ah�gL�,����	^}�k�r�r�cE+K*�H�̀(\�"�O��S�g�I k�n�z�EY%�>���*�.E7�C�IA:��+v�D�ykGP�pp��	�b��~R�̀��Ӊ�!b�E�3&��~��=�O��[P��N`�!���W���i��I�<1�'F�O�09 !! >U�Й�V�A��L�'$
�e�ӳ:_0F�$y"�5i�O���S�O���[!�"q�5�.'wK�U;H>!�V(5a�A����y�֜��m�ȓC`p�Q��i[taIA��1�"��m*�$���<>�|�iπ&�D}rd�I�Oa�Ys�>������. 4��'�������+6V��G̏ �<�:��� Ɉ0Y��)�@V�<*�`��"OzE�t�ߴy9�Ui��#�p�!�"O��C��X�G�`)k1��Y�(YP#"O��w�Þ��`�tN�}���p"O�Çl�89��=������E{c"O�u�C�\/�ţV,�/��Xu"Ox(��eC$O��;�%^��4ѻ�"O�I�#�O�:�$�d��PTM"D"Or�JТ�>����$OW���;�"OX��ɮTuD�'DN�?�|�h�"O������nF:�yCM�n
�"O�,��/����}
a�]eD�B�"O^�a'.�/N�8����p,*r"O���m$W�Ѹ��Y� T�"OZՙC�D'"r쩳��L��9�"OF����*M���(wN.��"Op��6�ۖ7��  ��������mX��H(�p���
�"U�,�����B'D���fB@�4aP$o��C��A)'D�\pQ-Ń 5��Q �C�N���b�/D�����n�X�cC�;��	��/D��3�����AGX�jE�+D��;r"D��7��XzP��V�$D��
Ң҅K�훇gg�}A��<D�LIQ�jC�p��!Z�VD򐫢�;D�D���N�y�D���@��E�g�;�O�OD *�o�!���'lN*;`~��`"O8-� �Ռ?�.�'Nڐ~H�j7�d�\���ӋJ׶Ё"Gtq.L���#�;Q�b�)�-ߘ�
��E�w���/-�>hH�'~��hQ��2a�]g�+�4I�'~νpk�"Ln�1��H"��`��'�I@�(�:�&D�``�!�B���'ݘ$PQ�,6�Y�'S+����'��x�Q*\�T���;p��1�ꔚ�'�j��f �8hm;g"΢/�DHx�'�`uCB��n�4���ü7�\����9Opl���18�ȳ���Fk�!:�O��4*��GP�="�E�4:U��P0�2D��[f�T�[���FDڞ!�v���m1D�|`B哺|Xu�sC�_��bF,D�*��}h�0 ��1����(D����}�u;��"�����1D��@�G�5Eg�p�	$0��"P�0��Gy���Ň�az5��'[�+�z4�u� ���I$kz(U.(�X ٩
�Q�3D�dH�͕�'��m�B�\�7(�ձD#2�I]쓖�O3�p�bg��^\<��)Ԫe�-��'��d�AJ�)Z�p�R9L��)��'���	�M^�(7�qZ���Fs��+�'by��a�(c��xq
Y�ҩk�'�<���J�80xPD�=��hR�'��Aɴ*{�N���.J9'�J!�'�R���S�zY*b	%��b�'n�q��� �it��Ej���':`�fM�-�*�A �� ]w����&C ��@,�!V�%`"<`�'zў�|Z7Տ1n(\����.� ��x�<�eP	$Kе0!.
v�f|`����E{���D�]wR��Q]�{�v )T���9,�C�I���-�"!�d�B�͜�n�̅y
�'(�FP�K�J����S�j�%��'R��WI�z
,[S*��XGR���'�"|���Xx@J�J�c��	��� 
��b��]I
UA��,V��$ �"OFD�䫞9�T�+V��7TJ��5
OV6-�-v��+Tm��(�a4�&z�!���Yy��8�l�[~M���X'0�!�Q4J�tEއ9��s�\:6�!�D�O=�"U8��0�D�	�j:�t�㜟D{��I�~���[�%��cq6,�h�_�aR�O���#��&w������/1�^��"O"qK"���5d���&��%j?� �xb�'|�d(N(��J�vTpFB��_�!�U�v�&q���(x �Xt`�"!�D��T`���&ʈw�I  ��7!��к^]>e��5�
#��2!��!��g
�( �" KN�)�!�d
!H�$�#K��%Y�W��!��x�j���H��AD��Kx!�$HAtY�c��?
,5��C۲.c!��XѼ�ya�*y��󏐑u!�5a:��b��R�p�
�/�/e!���z0
e�SB�^jp��dnB
	�!�E7��ӏ��he"�2�8r}!�d<��\aѨ�!J�!�v�-z!�$\29I�����
0>Ω�E+
�y�!�]<���;�;������>{!�$������. &ȕ�(�q!�لj��C��?u]�R���!�<�ƴ���)���J�
6$�!�D�QF�F�@;a�L$�%��^Z!�dN6.�u�T�B�-|�X{e�Q�Y!�d�n~�b%J�|:��#o�16>!�00!����	�ʐ�n�3K�!�D�$̝H�,[�f�dKs�S��!�ɯ3Q����O>`�����F&~!�¨t9��3���2���k�!�D�A�<�s�W,��U�Ѡ��!�D�]��i�����8 ��$O!�dܨv����g�ÏW����w�T�(t!�DR�EGt�RiǕ&�p��0�@"b!�d����G#Z�Z\�R��Ua!�ҟ{�b�{d"��Z�"�8��)cE!�dK?d�2T�U#O>�<� ӄ"=!���o����'��j��e;�$��I1!���mI�\�7m$R�v��֣��$!�D�D`� �� �fh.����Ԋ�!�ĝ����� �h ؙ�� ��!�ʂ(��iCSoX�!
#��6k�!򤐙At\tۤ̀%
�p���W-!����~��n	!!W��#Ӯ֨Qv!򄙂G˪�DU8E`���?>e!�DF�R��*�=�fH���k�!��,|�A!e�
C`h%�ϛ]�!�Xm��|�q Lb��m��Di!��B�5�U �q(���ۺ^O!�Ĩ*z�(��B4@Lek��!�D��4S@�!�?M��zsT/�!�D�}��*�G)f��%�󃅶�!��M�>,a(�D�}h������!�D�#\z���$͆RHvqy��L�|�!�DN�^�0���-O=ଈ��O�!�,+�m�	 0% Pj� !�$H,g.L4jq[�	7%`bh�/�!�䟍](.t�뜂i�*%�#�˙�!�D�6ޘR�a� B�Ta��S�!�D�G7�hra�ۿi�XA���/�!�� �U)�H�((��k"�B�|,P��U"O�]CG�Z�Q��+TAK �=�"O�-�ġI�2hd5�F�O<n�v%;�"O��'�U������4@z�"Oґ��)^�j&�	1pe��;�"O ��
��|mv Q�#ݱa80)!"O�\#�W�<�L��7��m)��A�"Oz�hյg��9BOE$~PD��"O�I��.H�k3:��
6bt$��"O2�0al��s�m�㋄)"sl��f"O��цM�.>Ɣ%B��+o8(�z�"O��-_�'�A�#�D�,*Ԑ�1"OPܠj��u�" DJ��NҤ��"O��r��U�y���1uKN.8@)��"O8$AĆ){��C	=F�����"O�;�.e,p2�<�Y��"O�,� �,��\'D�cxXT�"O���0��	��@!$��j�,P�"O�ܒ2-�7�DX���;K�vZT"OP�Y3�ޠK+��!���@:�"Oв�1p!��H� �|N��1`"O�������J�`1#ʑ*iM�Q�4"O��1�	[��us$H��aԤH�"O�YR���OA�����߲K�P3"O�i���A�o]�� ��(�0��a"O�䙥�!�Ȑ�H�{�(	23"OV�#�@(g�>-kउ�x4�A�"OxXbe؎8M��%;!��З"O��8ӨH�|�u�&�Ƕ'n�ؘe"O(|x0�I�B�F�B�aA�Hp"O�R%+�U�}I�^!l�*�5"O��2��S3>@��)`���"O���Ā�\B��cg4"��A`"O��@p�^�:�f���&�/�04a�"Of�1EI K^x睫>���xb"O&T�͉�F�Z�[�哢M�Q�c"OVY�N�n�j��0���zp8Z�"O�� qL�x����� 2K���5"O�5��.�m���Ru��i��8��"O�Ha3�L�rt�3gW�~�`�"O�]�	��~Nf�X�L�|��H 1"OhmK4��/>�}�#l��&q.�9�"O�z �3	�
����:1� �"Oh�B�Y,&�����>�ڡ"O�`A�&� ��t�LS�t���"OH�!͙p-h\�'j>
9��'"Od�i@�}.���;*NYC�"O|)��� ���s�ꄵtd]��"OT���(���(�	Y;Es�,T!�d�"%v�JD\�p��\at&�R�!��y]���gQI��)�dٔ�!��.@2P��d�;gu�D�W·^�!�$;U��@R%9V���Ԯ�%[�!�Dx� y�E.��Vz�i�n�;9�!�$�:E2���#1Y��K��ǭ_�!�D���,���%X��H��KC�!��ަw�&��R��	W��qX+Ԇ�!�d�
��� T�N����V�]�QS!�D@�a
�M/�$!{�(�(]E!�$�=t�f���"'d���a�1D<!�dE������N�oyZ}�ύ6m!�D<M-V��eY���ċF�\Pi!���$� �@9C��9��[�R�!�d�=G*��'��֭±J��~�!�� ^ �U�-'L��Q�JH e��X(�"O���Bf�{��p�)��%����"Ovȓ��՜Po����h̺�`<چ"O��#�C�C�,c�ĵ'�����"O��$H�J5,E����[���{�"O��w�2z(e�Uf^�"uܼ��"OV��]!nM�maR�Y�r��9""O\��҂_0/��q A��[]�)2�"O�ec*hzR`0�\���"O`�K/X��8�m��L�𥩖"O�0E枃P���1a셥����"O�q���m2��z���x��6"O*�ڄhY� d���jH1!:��"O ����:C�M�<Pܽ �"OȄ�p0U~T�[RJ�� �:1%"O��JF��0��$�iS�i��
#"O��3FE�*W�zeƗ+X䲤�e"O���C$ɫ�2��+T�ҝ�W"O�I��-�"i�l]KӉ�$��h�"O�#�G������^t��"O�LpFC�pH�)���$`���"O���SÆ�v}T���&��5�lDs"O2(�p M���ó&�����"O$�p��l  K�+W�_\�d`""O��E��e��$ҥ��V(�م"O�B�gLQ�d��ţR`�d��"Ohɺ�/@0"����P$P���B"Oj�`� �?nŮ���J$l��"O�S`��=��a�N����v"O"��ȕ)
��$�B���m��"Ot���GƞNE��	8�B(Rq"O�Tz��V�[Lċr�.3��	 "O� %A�/�$P�@ʔ5%r �r"O��[WAQ�HV\�9��@:!d�:B"O�e"�#�">(�c#!x	Zi�g"O���ň����iN����"OP]��\�l"0MCv�y�
9��"O����	$�"�Ύr�\4�v"O�5�(��2�ˡiǦ\�z,�v"O8��M�f.������!S9�dU"O��Ï�bM�xyaN1+�0ӵ"O�]�N�l��(����x��=!P"O�X�$l��V�t�����&!��+�"O�#Qt�(2�۩|gr9���i!�L�{QԠ� .�k�l\���'�!�S�ƴ�f����r��`�!�$D	b{2]+P(\�.̀���i��!�dӪh�R&�7obrYWC�(d�!�d�^�l�����ȱ�B��B�!�� ��4�7䁄T��f��{�!�D��^xS�k��/�2i��昔
Z!�d�j)ް���Xu��
惓�oO!��j�5���hgB�B���UF!򄟵liN��b�j�5�&�E�pQ!�D$s�z�sS��R�hI8Q��jO!��6e�veѡˊ.H D��`�xF!�$��P礰��
^s�m���12!��"a������F�I�Ȼ��4�!�ɣw�M�E�E"�ȥ�X?q�!���e�l�7�8M
�rg*$�!�Y!6rx�c7�$+��%]�!�!�D 5#@�EcY"��� �H�;z!�$!t�5��c�a$��,g!�L�;-64��,%(��K�kҡJ�!�� l�H�ƋD�>8[� 1nR���Q"Ov�1�M��KO�����ZBFQz�"O�i�N;D2�;E��p<$���"O*\���ձo��PS���)+#إ�"O���#&OU��P��'�1,R\�b"O6��F	��U�ȥ�t
""O��`#ϓ&˾�b�d�:�R�"O<�Ӧ+��׆4"�G�?�<L�V"Or�s��݅X���˖���_&`��f"O�qz§�?��49ëgn��u"O����Ɖ(�Ɲ����s)j���"O��l�/K\��e*>�*�"O8P&$^�P	�L�)#>��v"O�m��Ý�xf��(7�̖{���R"O��a�&A��Ւ����|�"O2��P%M?_�%�3E[}�M!"OP �G�	)�vm�w��64�N�I&"O<Q����M�(���NEI���#"O�6�;�&|�c�Z�.����B�:D����ȕ&M><�i�
91W�7D�� �ȹ79���'�U2v]�4� �9D��A�疵"��t����%�Բ�#D�\8���7��,"vDP=j�4�� D����5����N�ߦ�� "D��Vj�D���b��<O�|(� -D��S�+��p�,�:�p\�w�+D�x��RC��%gK�3>\\���%D�\���I�P���C 
�w�"<kef7D���C�8�=�K%�$lr�:D���V,��H�C'3��ų��"D�<C���;�2��U��*f�|!tC D�̻W�NW�b�&D
\T��6>D��Z��Ѵ=<�s���#��܃�1D�Xj#��	g+tA0!�E�:�h	"��3D��r�n�'7�5zt*ߣ<�Jヮ,D��	#��H
�� qO��Ea2'/D�@��+jqhPr����T���З�,D�(�IL*Z�Nh8D�ݾSRx���*D�İ1�A��x:�mN	!HQ�'%)D���QݼH/�a�AI"a�l�uc9D�8���u���s	D8}v�,3@�5D�����d���2���H���Xq�-D�p�U�3U��U�6�1 �fL�c�+D�܂�i�<�FU��	`XZ<��h/D��i�;no�i@�J5�8��9D���'h}�"֤����d�9D�|:�l�4dl# �P�	XH��j9D���.��Q��d +?���'�<D�`����Y�H��*	,)1�Ű��;D��33�Z�0��$�F	;�|-+"7D��PGϿN{RS��=pL���m:D�Xp��Կ��)��4s� :�5D�8�U\�>VW����Kn���'Xl�+Q�UD��Ō��FdU��'�zh E��2� a+#��kX֡��'�Ȍ��Z�Z��C��Ɂj�(��'����C-0q\uXB�Ef�l5;�'1Pd4��_Q��B�Y�Ұh�'^-��
�}L��[+LM2�
�'�TE{r%=��))�υ�AV!��'/�X��ǚJV�0�u��)�~P��'t8���IY5],����(q<T��'z�Tͭ`���E�T����'�buz�̭c�(��u��Pj��� Zmb ��`qb�i�I�3�6U�"Oz���/��k����V2wԺe��"O�����ǯv�%)A�V��I� "OV���)B�̀1�Jˤ+�Xh$"O��PtC�Ƙ(��
�x�a�t"O�}A
ӈq>�Q�)�!A��"�"O����/�J�����F��-�B"O���ƥH�  �1s%܈"�~HR�"O5)THS��ɐeB�"]�) �"O��є��,DJ��*�8bj�,�1"O�i�)�]�}ؐ�] ���Qt"O��)ք�V��!Z�-�4m�"O����3,���6�M28�*r"O�hP�;0��Y��@��|��4"Oͻ'bJ�l���{�E+f):�q"O������7�� ȳ,���|IA "O0sWg��1a�
5V�v�z�"O�A�0"�:xe�t�^0>Ϣٙ�"O*�ic��U�`�5\�r�JQj�"ON(�(�S~��Q䣔�7�����"O0�GID'xǬ�hr#�b8
-P�"O�(����d�6�C`C܋Gz*�R"O���K%n��u(qԔjC�]�"O�� ���H~������&G1��	�"O��ɳh��/��@Fǣm"�8�#"O4�Xā�����''�,�x� "O
�II�_\B���)��ț�"OJe��EV�	8�E��"���"O��*����N�*��c�G�Z�p�"OR���=X�$�Kb��^Ԣ���"OЀ��J��O�.8#�fO9̬�[�"O2��� ܥ ��M;���A"O�, Q�1G2	␭���Q5"O�I����j*�M�U�I����J�"O�TQソ"]��@:��i��"O�A�(��&�a%�B�B�p��"O0��AcN�Ryp=ibC�>D���$"O�i�&/��P�h�!Ä���(�G�<Q���*z��ɛHl�,���G�<!шˈ��͓Sm��&������J�<ٵC�:M����O�uSLxq"BC�<	RkӇ'���)3�SP�i5 XE�<��ÜoQ�4��o""Ir�nNw�<Qba�Mt\���Nh�݁GXH�<�1�
�J�JE�#��*v:\9�Pm�<!���%"(�)ӄͨ3����Lg�<� ��A>$x�-L�*ðLcum�e�<�S
�&t쒰�87rh���Cd�<���M�H-�̠pk��c:�����R^�<����b,�%H���CDܨ �M�b�<-��/J�P�&�!��.Y�"������ �"��qz���7Fٯn\�ͅȓR�n�����iH���Z&)��-�D@��a��_�p�"�Ӣf�)��/� ��a«B�P񡂯�#Fq^��ȓ`���WOG��N����O#3�
݅ȓrF��䩌U�xl�!oH.tQ��Nah���i��G+��J�B�t���0r���o�@Y���"����ȓ<��E����_��9"h�բ��ȓc�V�13���ej�)�>͇ȓ;�4�(c�D�5��d�лDM�0�0D�Xao�;AP)i����xw���f�:D� ��OF�Z�+ө���ܱ�d�7D�� 0`C T�3\}��É�T�J���"O��Rt��*��K�r��]��"O�K��Ȗg$@�G�Ū5�v��"O,�be���D�NX�傒4[�� "O�5�V�@[�d�U�3E��%7"OX�sv �� ���ZR���D�DA��"O����C�~���N�%Ip�(w"O�|0��W1}��Pa��i�qR"O�0�o��X>�hP���F�Z�"ON:�o�!Od��Ю]�|5�"O���.��cn��{e�:����"Oȅ���4tr�Y��C�|���q�"O�<i'圇*m�y0/��}��QE"OZ5���ڂ2�-bGO�~�C"O�D�F�R�α�I�:}�0(�"O�a��v��3�U (����"O����O��u:�%��o �f�u"O�u��К2�^�RO��z�|��"Ohy%�3�X�c�0\X�s"O �֥�]E��ؒ/��W �F"O��c��ru�qf��z9�|��"O���4���5��y��R0��f"O����Ҫ��������0u"OЌ�g��$��Um�(֠;�"OX���!M�L��{����h�{P"O�xx�C����G��vH�!"O\�r�^6���B�H�vTH�"O�ԠԀ��N��;��. ��Ӏ"O1!Ƅl� �%��?ު9C"O��z3�L9C�)@�A|8,BE"O8�1����1`o�ckҤq�"OF�!�ŔP�t	CP���?i��3�"O�M����2�naZs�E�G�l!c"O�	� �;'2���J�9�y�""O�D�$� 9��^�d�ҡ� 5l�!���,0^iq�Xm�X{���vY!��3Uo>����:i�C�R;-!�D���N�"�O�<{�����J!�+�
���铯t�r����V�!�d��gp��[D���u�9(�#�!�Q0\���S�>W���
�!�D�]|�Q��K���0x��Y3&`!��)O�q#��U�U���z#n,�!��ӱ%H�u�ܟ7e�lXPM�&0�!��͍d�ډ�W�	�Y��5�0=�!�D�o7,(0�V���� L¿K(!�DѮ5�F��ӮD�\����g�V�|!��
�/dT�J��QGs���BBE1�!�ć�]���ӵ`������c�!��Ͽ<�1Y��>Q�f�����8,!���3��)���&u��1h�V�t�!�$�H�R9��T�#�pu�AoB�Z�!򤑀OS�	�ҠV�����0��k�!򄄩h�ڈ�P'
��ۖ�A�6�!����D��[�o�ڐDC�|!�d�K.>�0����q���P@g!��Y��R�I�n�?E���&��"x<!��n���Q�
�^����BlRa;!�Ǫ	��}��ݗ[��k`�&!��R,Tۄ���'xf��CB!����H ���~�����ӥ�!�B)  �!r�J3k�`�r"��;�!��R�z���E� �2A"��9�!��l�t���Máʆ�p5�LQi!�� �U�""���R��ۍ?d�x�"O�YBF�^�6Gh<�!=(&8��"OPQp4���fgl��^�]�<DH�"O��ȕ��8�X���3�4鈂"O���W�M3�P���^�9Cx�a�"OT4�"�Z�2DmZ��M~`pW"O�9�B�ƋQ,|���R�(B,5��"O���Z4Y�N��l)D.d�`"O.���	��:hP��@�>M�p"O����ʔ(=�R�������y"O�5+�S�b B4���ۤT(&"O.I��MRf��@إ4.��v"O����:�a�́�"��2�"OP�!�	�Q��@�+L�f7"ٸ�"O��;��T�@�$(�� �y;١@"O�X����9v�jQj��)mC֑8�"OBl2S�0���!�Hk�@�a"O�	p!�J3�`���/�V���"O� 8&��54�H�`H�&�:�"O�$�#��+����G(L��h��"O�E���6��7)�1���+�"O��iCk�:H8�2򨅯^y��r�"O,��VGe6��@�e��tk�R�"O0Հ�HUkH�phEeq>�ra"OJԸ�i ��PЉ��`\�a"Od1��*��d�D�<͂�K"O�e��[&��H�S�����"O>���(Y5;�@�r���0[��Pz$"O\���C|9ug��9y���!"Or �$�..v402ĕ3V�m��"O8-h��WT_z�X�"T�V��'"O�@Z,P#_oJi㖄�O+x(�"O�n��o���>b8����%D�� m-��� �;k��aF$D�\Q@�Z:t��/C�hZ�%n?D�tY�d�T�vmx%�F�9jPѠR<D�@6#M�V>dܹ�ĘYaN�0�@>D�P�X�zz�#1+9^:.�0�A7D�𓓠)Z��G�@�m�bL!7�3D� ɐ^$�.Q��B'o����f5D����Ɗg<e:�� �x�z\�#4D�h@���bօYF���~�2-�V'0D�{�M�h���8�cu�f�Gj D����\bXU��&��%�bݒWL;D�@��&�@A3Am^�+�f,D���EЉQ�p�� #9wJJ�P#0D���s� �@����I1]���(D��r/ݓL�<�A����y �i�צ&D�(��͕=
;@tJ2%PT�,aj�)D��C&��?��\j�#�N4@�	'�&D���)�J�J�K�Ê)y�4I��1D�d�L�;&(�����ONpQ��-D���e�6�6�h�g(2��(jBF>D�0���!�(�8G(��kP��i�>D��9� ʸ��e�;~�H��d<D��H�Iĩd[�4
�+�Ld���3a D�X�-�7�JX��<Z��I�#D�8xע����  aمMRd�
�&D����A9�̴9V��3H��e�A`#D�p��(��r-(8�@#K<4h��?D����h�:<iɡF�n�^4�'#>D���� PGbL��W$[�}�P�S,=D���`��zU��`1A�"s�����:D����-�xrfS��4b��k��*D�� 0�ׯ's�
����֩s�"=k&"O�<S�&��i�,D�B�SҔ$��"On��R���$�@0D��t��驄"O�sQ N?��YJ1����ȹ[�"OL�#kbİi�"m=�np��"O2-�G
P0H�2ȋ�B��?�a�"O�����(��}�egF�]O�Th�"OjT������K�],&��"O�!��'I�����T�6�aX�"O�����n4�đ7�\�"����"O��2���:������u�����"O�Л$B����-�𯜀~�j���"O���W�M�0�Q�T@O�~�Y�W"O��b&��_�d-:��S(3�<��B"O��y%�޹p��S ǳ|��HK�"Oh�@b��uZL@Sw�#Nq���"O���.���b��O��u��"O aBeFƅ/d�1�F�G�*�H�"O�l�&�O�����V#�c����"O�u��إ+�x8�c�V8�X��"Oj�9��;x�h�$*�#�p���"O��@gQ�&�� ;∟�F�0��"ORL	�		q=�;�m�i��a��"O\�����1e4:�/U�(�;"O���g��GG�*`�x�|�Qq"OL�bV�ȶq�)��b^�Z�XYS"OB�
4aQ�L�^D�F�>a. �X�"O��0��\�2 QcK(F�iJ"O6���X�p�$��#{"�,#"O���dI�.y��M��L͈�n$� "O@�i�# �><�U��.�J1�"O�Y�ūC�"�	�*'���A"O�q�M���9&h��hb{�"O��Ѥ�Raw���Ɖ	U}�*�!�DS�W�#�L�l;"H�sF9m�!�$ۼm�d0s�.�X>��%���!��	� �a5&¨�N=��	�)>�!�d֝��Ոda�&x����3�E�|K!�Dc��|3rL�'9��i��F��L<!��	�\��}�Ĭ�s]�#pHʕbB!��y�2�i�䚉3,y%g�.1!�D	�fYvezC�ۺP���=O�!�DX�ȁ���S)}�8���ԑ2�!��pH\�;�ƌ�U����F�c�!�<;L�`95�R[:H�Ufݵ!��Z�"i�n֪[+�b%�&h�!�Ϭ2�$R�A�u��Yb򉆶F�!��ߘm��\�E��M����$��?�!�dG2;L�ѓ&^�,�.�v*Ӝ�!�dL�o�(�����$�#�!�䒉\�<�F�%��X���&M�!�0@�z)�kW(��iQǟ9w!�$ ��5���)pz�� ��W!�$�3X���O�s��}�V.C�
!���5`�\�qSZ�����_�?�!�΢U-��`1o1cjd�7� �!�ğ�FWv��� �� �s�Х4�!�dX9~�J�D�.,�5�������'���"�`�n�{f���!��'t�YƆ��wD��;Ag�%<�����'�@�����'\��� ��5% �9	�'�8D3����O��(`p,3��!*
�'�4AQw��z�Lȷ䞆#c����'�e�59#�1�ǏDGX ��� 2��n��w��XD�&xv���"O��P(�m8�$3�*ߛծ�i0"O� ��l�wN�]"�@ԑ
, ��P"O\�Y�;N�D��bm�^J-�A"O�!؄�ˆ4B܍�q��{-T��"O�,��Z �y��U)Ql髱"O��ȡ�A�:Ql���a�$���"Or�[���&$�xq��3j��"c"O�eֳQȔ�%W�P{��R�"O&q�#�R�jS�H[�$Ui$�"O��
���7�\��b�
�SLсP"OF��"�Q�1��h����3\��"O�4S�`������"��CJ��"O:�!cmۣa���D�M�q)
 �#"O��WiJ	w����I�:t��1�"O��XѦ(D2\(SbŰ�(��':�Ӵ��+{w,�+��_�6�:Y:�'!��;r09�*5�%\�-����'���c���GR:!����z����'j��s��1�歃�%�b� �'0���F!3�A��\8L/�T��'�@Pq5
�I8 �e�R�G^�ȋ
�'_Ȑ�!fQb��g��tQj��ȓ{���ʤ/?x�6����F��=��=�|U��i�.�4���O�\ʘP��u����!� x�U D�-*E���ȓ3�X�B��??��|kp�A=����ȓ�<���H_{B�!�O�D*P0�ȓ7���	�&���9V�
z��+����1�I68�	Al����x��/D���o/%7J��ׄ8�	�ȓt�D��>}�(��/]��
�����)s��'f�ҝ�q��tȓd���1��!YP���L��S�m��c9�1�G�ӄmg�����>+����ȓ���#6)H�/���	;H�F���,H�8�gߍ2w"�*�J�G�p�ȓ��( &�53FXi�F�6g��h�ȓ0g���!��Q�j�sc�D�"]<��W`��J���g}����AW�����sE�p"3!݀n�e��K�g��ȓo$�
�6o�
��6
��,x��0"�����6V����'5����	��a⁈��e�0ȃ㕣}�Q��qH|�IG,�1Ij��!lىs�}��*�`��CB
: q��lիl�d�ȓP`,(��*�4s���ɋ����ȓa�2U��� ,#��G ���0D���Q�_)*Q"%L� }����e.D���Q�P�9��0K�iv���H/D�8�w*9z|����|8x�E:D�PJ�OH�J����k�F��W-D���6�#8(V�06�Ҿk(��Q�>D��RvU���l?fQ�/ǂ�yr �?�&��cfԊl�,���$�y�<1��iV:5��#e�9W�e�<���ӻYd\k���!�&P2ӫ�l�<�R�_#UJRp�ٻQ8�d�#�Hh�<	7l�+~��� �?�L(ɣ*�c�<�7g�!8V�X�t���~fp$qL�W�<Id���uId}h#�pH�X��U�<���)��ЂmV�P�x���Vg�<y$TI^$	���o�|����I�<�&N?Ed ��׬Ic(�:$D�k�<� ��J���9PhI�4��*H�ֱ#�"OB�	#�J�_��y2��c�ZL�"O��XC'(\�aU`�i��qXv"OT��.�w�����{D)��"O>�2��)M1aS� /=_��"O$$k�,��*� ����ƦKTމ�"O�%b	��C��9�gR�'R�i�"O�HJF�U-��T�򅍊f�HE"OD�F��&�qE�ȉu�$�""On�X �A&E�N���ϭu�vUxg"O��!B��/!vLl���PB��R�"O�!؊iC�-K5)T7A\ ���"O�@���ȘT �"#ÜOC<�3"OthRq+�T5b���,��"O�0�r�F6�f�r�AԹ"�X��"O�Yi�&GN����8�=�E"O���ĎV4r�@��S��]1�"O���`͕2bl�XՁAJO�=�C"Oʼ��
ܔ7�Zm{A �'6:!rG"Oީ�F�T?\B��2�M J�";S"O�]q#X���qa�nյy����"On�٦�Z:4N�Ր���:{��"O�|B"F�.�jx���[�r��Zv"O֙9�ʕ�2h�o�1|_���"O��3��P�0ͮ豰���\�Js"O��RP�QT��Y������(�"O�z�S32��c��	01u\�I�"OB�Z`�$X"�Y�BfD=��!d"O�Y���04&��pt.޼ⶀ��"ONQ��g� V`��1E��M��;�*O�<����{R���6MTI��<��'B�QS�ť}����cǿs����'�(!9�E��6����P��fz�]k�'�}y�I��U ����CG�K��q�'>�9�
ɺFM U��jJ�=�8-�'K����H�2��%6HE&�\��'"J�S ��>O�\�R���Db�H��'���������2L �D[u��'�� �Ҭ��f�2k\�OF� +�'V��p��^��(��
(ynݠ�'��PK��3]��h@�&���'�­���0|5��7C�3W�M�
�'sFAç�SUU�S7�*�PM

�'ע-ہ
�.V�r@�_%
=���	�'l$��t�N�3��h���6v�J�b�'-z�f��;;"j��f'ʦr1�p��'Ԡ��F,�5�Nq�( ��'3
����R�X%��s��U~��:�'�����;��y��JQ0t�LT��'�l��K�y̔�Z�eF�2
�'*���"E�<��S`��ɀ�I�'���惖C4���B΍[�^u��'��%r`j$\�`�S#C�a���'���Z�HB��lejkߍt��}�
�'��\h$�*0�T����3s1���'ɦp5Y�����=?����'�P�$	f���7��.�j�'UP�1EM^d�t)+G���
�����'���׌�QAh �6���H��'ؐ�@Ć!Ѳ�x#��~\B��'8�XG�[�"�� ە��=vx�i�'�P�x$�B�&┩��F#^p����'�~)Ib����X���H-\R��K�'����C7p��q$b��U5�hH	��� yz��� /�� �i@���c@"OJ�� �Z�+�0Ek@�ι&��mj�"O �*�(ܴl��e��{|��2"O��8��-R��(�+����`"O~	!�ڹJ����8y�� "Ox��s
����ht䋂h�L�"Oj��5�I�8�0���_%	`�l`0"O����K_��HE�7S��y"O��#� �	*ȱؑ!�6S`�4  *O(i���0uRС��#�X!H	�'�l�+��g��@D����-X�'����%�@�6D�I�$ ��^=i�'2�ܘ"Q6��f@
,�&h �'��@ ɚP���Csn��y�$!:
�'_�A���W�EՀh"�n�����'a�6O2)���vߣ ,�y�Q"O�iu�$9��8� t��Պf"O ah�a�'
�E��	�x�0R�"Oҕ�LH�p�0�1u!�8j���"O|dj@K/3:����	@>�I�"O�BA�D'�0Ѣ����E�D�Ӕ"O���5��&49���`��*���C�"O�|p4�:8��z�i�<-����q"O6m��W$�ݙf��#���A�"OH1��5=��a�h]�~ЛC"O���0���[�J8gN�1e�9��"O ���N#(�����7N��"O4q�Cʧdh�J�,��;(	82"O�؋g�#�pÃ�Öl�1 "O�P#��[�G�4��c��-!!�9��"O�!�Q��p�aѳC|�i�"O��Ah 5bx��ӬR4q�"O a	b��n\H0��]=4-zb"O4 s�A��깡�� �^�FC"O�)�G�<P�,D�d	�8�P�Rd"OX`#�J�V� c�U0hp-"Oz�U��e ���CFB�"O�@�O'��	 ���"D���2�"O:P[3fN&�rD�5H�D��c"O�{Q�Q(}c ����B�
ºe{�"O��iX/؆��Ro�VO�"OB�çȿ
��m�4>���e$D�P��	���H���W
�<��?D�$z��ǜ~/~��E� ������8D�p!F�Ņ��Ď�}������9D��1A\	{���q&j�Q�|�ѵi;D��[�Ěg�z��5'��O3�pz�8D�H���O�C�����J��p�7�1D��Ip֣�Q
����V���{�2D����M�g�!L�1/�|ԙ�#D�,0��T�Z�x���Vz� yҭ?D��P��C5EG�PTD|6���C?D��k�h+��x��hQ30\�D	?D�d{�@#yQ�DE�4��}��*OX���OI�*(fЪ� �
v�V���"O5�B�K�E>"���ʃ#\�ig"OڬT�E�9�<�
���9��pH"O�$(��X�ed���$ι:��-{!"On�!�	� *�c��A.8)&*O���@�IXXܻ꒩06ɻ�'�&���R�H�fZ��ԕΊ�!�'�إ�"#$�^4q���bw00�'츠�pO�2x���`H�)SZ]��'% 8�7g��*�N<�	:(�� ��� �1��U���k��׉A�5��"OxQ
6`�P�P(�صI�"O�񪥥�8��0��.�Yn>́�"O�૶*�rd�ʦ�T*/\*`Z�"On��2g�����y�l[�F�A��"O>�١��1��C#ϲgB���"O��I�R�'!VٲwhN'4(5"O�P��K�nB�Y�DH�-��Y��'�}�D�Q�6�^��&G;YPL"�'{d��SG�FE �h��PU��;
�'0Z cW�ҷ����uD�H���'��	�M-/�~!� �F|b|K�'��`��)K�_a�)�$j1����'v�!�g#'��4�]�^��'n�M
5@��dR����^�^e��h�'ƨx�c�~+,�
h�V-�
�'x��Z�L�5�(��˶AO,�Y
�'F�q&f\,7I�A���jO��s	�'�D���L���Ƞ�)�>6i�)��'�l�4O�0}T8<p����< p���'��U��cE۞�F�� f ���'f,�"�ʉ�R�I?���'��X���H�@a
p҂��w�X1�'�2݂�ʔf�F�c�I�o2��b�'&����N������F[:b�zA��'F�d�C�zc!��fA�*�����'4�lE�
{
�z�"ȔB䉎O6��Ï�/W %����%��C�& �:��a�Vk�dq����"Od��cD�-cy��'��W�չt"O���`H=k�+z�2����!�dۉmD��S1�ۋn?��ya$ ;s!�D�"��4� ��>��@� �%"�!���1A��II��A�~���'!V�Z�!򄁶Y)R��h��;������[.Bm!�dƵC�$����79��q�ஔZM!�X</�&<�Kؚ7�2��6��d�!�ɘ{jt`$B��!B�;T�C�1]!�2'�kVƇ+:�PQ� �)1!�����y�@���	!�)�2�!�I4��`m��<�
�Ȉ0N�!���a�8�s�ˌ%�R��N]�!�C&�zL�@ӥ ���H�샽J�!�Փ5��h��J�*R���b�9xi!��ө#v̰J�����Jᄧ 5X���*n 6�R���Ŋ���u#"Oځг�L!JeʠraJ@$2`��k`"O$A9�C�s��=���D�����$"O�|c�͈�htj�+�>,BRu"Oj�P���;�t�	�+Q^�>�K�"OX�!cK�	I��	BjX�.�]s�"O,\aG-S�0�Ę���?74��ٕ"O �z��G|��=@���?cMX9z�"O.��S��! �R�O��G`٫3"O�T����_ƨR`��@D���c"On�H1�[�Etqb�$�3%&ވ:�"O4][�oΧ>�ƥ��eǔ��#�"O�51���h�-�D;���2"OPI��@1"�x�[qn�3蚬s5"Oظ{�c�i	ܨ�6	�G9nܛv"O�ܰua�QF�
�旤B���*�"O��`��_AR�x��%W�DLS�"O�!xB_&+$���Sm�@l�c"O�5	6o�	�XAZ$�݇$���""O� �e�Ak	:ek��K�iѿR��TZ"On�R���D�+Ù�z�*p�"O8H�6�·&�^�x�"ހ��ے"O�}�G �	 ��(󠆳z���aE"ON�D^��qe�F5C<>*�"Op��w!ŶtC����I$���E"O� {������Z� T30�U"Op�s�DªNe�D�
�G ���"O��� �Q?<�a�i#	�r4*�"O4�G��I/؄I��� qT��!"O�����4�,�b�рa�|Z�"O$A����3T:�1Ӊ�}V����"ON�)���|�Dx�T��<0=*R"O��aM��>
�4�����D)C"O�0�g]"Y��H���M�Oab4R"O�%1��A����ѥ@�bn���f"OƁQD�ī?~@�R��? "Oda�`��Q��*��(t�@Cs"O�$����)���k��S�V��8"O �9�"^�U�"�b ��g�F�p"OVT��&Q+2@��`I�kxD���"On�a���}��)�"n��n*���"OvL�&�;����#*wV�59'"O���/^/؋�哰S�r�y�"O�x���±/fh��p�ЄJ���"O����W�A�m���e�Ak&"Oj���唧/	>4� �ڝi��h8C"O�0�DaN3�8�P�h	�6]���"Ox�6H�yp��*P�>Z h�A"O��E���r]�xq�o7L`�0"O|uza�	~�b�D�nOn���"O$��!>�v,�6K�.�*�0q"Oȝ`t��b��,�� �a�P�"O�}zgN�+'%��cS�G�g��Æ"O>d����%o6@s��R�O��PD"O6ȉϖ
{:�go��l&&y)"O�Dӄ��'#�����
8��uk�"OX��
�,3}�I����k�F�"Ob,'FMb��� ��X9w�~xrF"O���с�=�V=k7'� @�vx�"O��g�5H����6�S�|��;D"O:iwK�8q H*�!�0�
���"O��)7+ǅ2��AA^y@��h�"O|�K7��
� �#p�Ћ?*~-�b"O�8�Tb$k��Q�P"(�1�"O ����>␙#��1T�"U"O�Ѻd�" ��t���oW�9��"OB��ŧʪ{�	0@�77@�D�g"OԘ����n˜�3V��l�\�Q�"Oxp�6�L2���S@@�p���("O�:���vhP �%W�a�d(ѷ"O��уA�2�y�e����P "O�Qb�d�s���C2��f���"Oਲ਼�Аb��YȆ��=���q"O���gP9B^��`�����l�"OFy#!�L=4�Z����� F�.=X�"O,��P�S\���V�F�Y�"OФ��iN�`�`P��Zla�"O��i���ptA��X�`Ml=�"O8��"ȑjpS�n�u0���"O�P�r�����0�+�=#*�A"�"O�}�tk�pS���A
��Y{�"O���j��w�Jh0щˢ&����"Of@HV�O�4z�j��L)�d24"O� �m����3l\��G�=r��"ORT; Ѓf������{�Hz"O쩰V��WV\�K�ʔ�A�,=�"Ol�q�1Z�����\'8�h�s&"O<����!+� ���j
�Q*��"O�4B0̄,Ϯ4���5T��"Or�S�@M�.�d��%��e�I�2"O`yz5$�p���	E��@O ]��"O�U��V�e����lf�,�"O8�Q5V�~Ȳ��$�U�@�"O�5��i
K&:��CCY:P��4c"O:d���]xxQ�o�.z\�r�"O�Ls5
�7s�<}�D�llvTQ�"O��V�1��!�0�ò
�(˃"Ox�c ��m���(t���r�4PV"O�lR����4Ɇ�iH%�Rb.T��;��Q1�Z ���ʁk�F�Ӆ"O�غf�W�:`�>E����"OĴb�_3(v�t�w,��m-)�"O�)*� ��n�����$N�u���"OB�P�)��f (��@#�-b�q�@"Ohx`�J~�8w�-��Ż"O�B6�S�v�vT��J�>~�6��d"O�� 8>��u���e݀lA�"O�ꕁYQ��İ���G��,��"O"$�
 t����T(�d�"O�1���M���e�3V�y"O��T/_�*����`U����S"O�3잝RB�P2`��s�n�Q�"Od��Q`m�X��8W@���y⦂#"�H��VQ��A�CO�yr���u8xJ���ʕ4���_��B�	�5� F��/5>A0��L[pB䉗�PŁv��(y]Y��бJ�B�ɓo����*� 5�@����C"O�uSW�U���i�ǧυ~����"O���� G�vP�dX�%ŽmP��"O�Y�B�,%j�zVج����v"OX���m̌~+t����5V`��Q"O�a�1�K0��a(�
��X���1�"O*�y�R;�n�Iؐ��uC"O�x��Ty:�B��?�T�@"O`���?|�b" �	�����"O���֥ݔ~�za�i1,�DL#v"O�Юˣ � Q� $��0�:��v���A1WK�	�йt̭c��ȓ
y 1�V�^.*HE�a�^�y�ȓ�(hH)ם}9\��$L=�����7�F�pԪ����`
T�Ƥe1\s��O��=E��	�z�R9 C(׺?��x��]�yR��v���)ZB����j[`�=E��J<�����&����וX��9��t�'���F�֡Y��t�ǌB-S�>��'f�@�F�'qh9)�S۠yyM� G{����Ǿ,o���r �i���S̀��Px�i�"0�V� MB,�@�4��E���)��<1d���Eˠ��wF�*9���z&��Ih<��Ć(n��iQ䞬Q�����m ?��D�=s%�1�)�"N�>���K�r	�O��<yI~���}B�5��I\�<�i�䑽:�!��Y.#��@�åY'e����J� Gx!��ǹbvx��/��>V6카�8G�!���fTxс��[I\Y��P==�Od��dV*}���3/��jD+���.�!�D�O� �,Pf�#:�4�BI˒]g2u�h�v�'�����3AZ1y��ѻcCw�r �W�9�\��>��#���^9u��o��&��w���v�'�vE������H��A�X�OB6-,�S�O�L��G�, �,� ���<,i��'������jz�p����"q�$����'�S���_v�K'ɍ=D��z�).�0<�r�Db�T�c�/F�S�ݷn���;��9D�\��-�<;"�A�/**̨�3�¬<��O0c��Gx��ٙK5K�ca9����
0�xR�'n�C&�.'J�m�6W�dkZ�H>1%��X�[�j���ƓHI�9r�`�)F76e����<)Ɖ�>�\c"�t�����<1
��OR8���r$��ū2.���	�SRQ���1��5zh�B���Z�>�j��t�Bበ3� }YեĲ1Ď���P�6%D�	`����6�$5��6��S��xV��p�!��B�.�5��X�Id�|AM�y!�đ> I����J��_1� 0�� ,n!��<f6a��-�"d�ZL���^!�$C#iT�;�
�#V �8#��2_!�d� �T͋i�!O�
�m��/�!�ݸFBH؋s�8�I#����!��֊B��ȳ$
!|��t�;r�IEx����G^.*�
((&��4�,�;��>QÛ�̡�a��R������5|la�6*��0|��LġF+��тըNG�UH�K�<�¬ �s�ȹB���z�o�@�<���7��ص*�Oq�DK�/T�`D{���N>E$��6��:PĜ��$<&�<�$M����ܓw|8�d�-d���7��D]�'P�~�+A�޵�S��3"H@�5�yҀ�d_Nh���
�5r� :�y�O�}�� �����[�B�y���p4(�1
K� �P	D�ēB̢<�~����8j$�J�?an�Q���_�<����y�����y��	��]�<�@�{ �d���3o���Y�L�W�<ɕ�B#KDd��q��;��<�gNS�<i�ch��T�!�*��gA[C�<	A�	�"���"�'/���H"��@�'�ў�'Xo2�Ycn���Ա�+
�W ��ȓH<<T�"��	t��I��� J�\l��vV���Y���qa`�ݓ�:�ȓ/6�M{�Cޟ+f0y�bD���ȓt$\��eH�&���9���)	�XX��*Q���-��w>Y(�a(m`�D|���<���@���94�20d�#c)
B�%eБy%�̱b��t���	7�B䉖i�zuH#�-sFX9�����C��"?0f9p�"
�S�
\����iK�C�	�YT���$��i���Fm�`��'���mۥM��t�w�dݔ�`�'
6��p�� <�x;�]#E! ��ӓ��'3򨙓���a�.���@ſ5g���'��qG�2/�422`��<�Ѻ�'4�Dp���qT���./5ΪQ�
�'X��"�R8k2���NW�`��5"�'�`a"i�}[T�x��+@3ta��	>D���se2M&�h��%�	$wZ倳�/LOP�P�&��"�� �W���F�I��+�O��I�|5\�����
W�.��E�Z�^����O4�A"��z_�#I�Cs�D��"O��l0J�
Փ7�W1���Z""O� d�ȦD�:(�b)#�X g!�� S�	]ܓ��'Y6xR&�Hn���K�J'GP3�4�Pxƃ� ����ލW�p��ʐ<��'D�'z>���mG�@�[񫓶$�\@�� ��0|b��/r�^�
�
4�l��[x�<�uD7 f&�ڃh�T�J��p
S_�<����kV\��A����`���<Qsj7,���H�,B>F��3!X{�'=Q?��F 
o��y�杮pȸ��>4��c�iʆ_��X8t�I��Ȍ9a LQ�<�tH�+�A�Q��47��pp�	G�<a�I2:�n]2��ع^r8�q��B�<ق�[�=�쐥)�4 ��@�'�Q?i��_�b)�1�q��$1�����>D�4��C�D�1CW��d�d�B�뽟�sp�)�S|?�vc�3&�ңd�:Z���!�J�o�<�fb=^jjM���� e�_h~r��xD{*�]�a�!P8����	P�9����1�'��'��	����TOM+Z/4!��W��B��C��k���&3X�Ff'w�C�d�<Dp%�Q�h�$�� |��b���	�V�s��д\]1e�_XC�I+?5XzЧȽ�Z4q��73	C��5}e��za��Md���w�L�)�����9�$�XD�h�܅K�r���O.Sw!��Y�Re�} ��Y)lfH��7vj!��9lȢ��#���d���E��t[!�dʛ��壵.��=�
��Y�q�!�d��:	�2mN(l�
d�U$��R��!��'{�)§\L
h3uB��:36��u*J�!p��Uі���W�h�t1���0-�x�ȓ_���+=�����Ɣ��a��f"b(�C�F�WR:��Ы��j�H��ȓ/� <�a�@�n��|�`�JUդ��	Z�'�R�XӉ�(�XX�f���}�J�0�'!.�y��PmB��� Pt�F��	�'�l��f ��ؽ;b�ɭV�<�q	�'�"1q���&�@́�	Ê]�h���'7�AgW�;B�t�E	]�Z�P��$.�',����ƺ%Wx)�')Vw���ȓ2�  ��G�l09s�_�_�ń�od29���ʒ����3���YN�h�ȓ,�Ih�38%#��W/(.y��o= �s�!;��*�*����@14�)6˚�� 1Eh���ȓRPmw��?RߦE �(�XI��Bz�9&̚&����P���k�E�ȓ ;8 R��[�h0xWO�'D+��ȓg�P-2b��2%$L�+��PJRY��jv���f����4�#_�/��C�ɏ���!�`�<5��j��ؾC�	0s,��H�C!!U�%���lLB�	�����!J];3�ݨ�(ٙR�DB�	�W�R��0G�uWj�JtB��H?�B�I9,t9���AHz8��6��qpB�5\�V��� _6i���L�VB�	#-�b��$k
>�����+\5�B�� CH"�bT�]��=qe�G�N.
B�ɈA��}*1H��$�2e>Q�BC�I���-�#F�5} �4��+�2C��K���Y%�*"�^����j��ȓS-�x����<u����הN�|��'�*� ���%���֯O�A��݇ȓ}D�!�!>���c��[�9��S�? �	B�"66^؂��9f)`H�"O�d6F�;�4)��ÍuΡ#!"O��QR*L�
=����"rh���"O�p�R"�		���R%�� jT�"O.�J�K�U�Q	!M4V��2"O`M�&�N�Qȕ%I.4SL:�"Ozz�׎Pע��E�%6�:1R"OT�K����G\^e�-��y˔"OH�0v�C.�V1�����|�F� f"O�`�ҀO�g��d�*N��b"Oj�ԉJ�F�v@��(9�UX�"ODث��Ҧ%r$)�f��>Z�K5"O�Dj�T^�����߫()�tAG"O⬒�2��-Z��
'0�e�"O�E0c�U0�&XL�[��O|�<y �Sj��葫܈*��4�C�Fd�<��e�%k�`��+��!��){7j�oR�`
@�̥^��d`�	Xq����1��,İ���b�(76|��+&D�0���P��:��5�)���ɢ�!�Ĕ��]3sݐ��
A�|�!��I�Px�녡�J�����!�N�'Q�Q0+�@`5RP�K�!�d!��
q��&�t�	�@�!�R(����ڹ4�<��!F�?�!�6Z�P���<J�^h��e�=�!�\�TD�y��p�p�˵�Ď �!��̿Y-����� n���Ǌ��p�!��Y�0���3̋$U��B�h��[�!�[�;��=��
jظ�����l�!�D�qS�X�@�_ø5�a-�+H�!�D�^�L�t'��w�X`�kZ�j�H����=��z��!�$0f(�g��ۗ��+b�Bp��u�j��SK�.d �X���&x�r}A���;�"�Z6�O�����W����^ T��Dc#�c@���H��~�!�d�:apm	���n��I�����x�V��AQL���蝵�
����'!jP[��U�DΌP���	 V�Yӓ"eB��#�х.�8#ګ��+�UpZ�2�H˼JL�R���;�y"�/B�����4OH��� ȕ�r�y@��5���v�|R�����&C+8�Hq�G�,\���k4N���@�*4��+�� �;�V�q1n6Q=�)�R�/�O,	�鈜}r ���R�J��`�fA���������:� ��hK�m<)�i��t��� J��l�&1���d�ޢ}守���D>s���c
Oxu�@D{X�I�0��@Ƒ}4Ll���U�1�,s@:�n�w�D�}T0cO�3�� ��P?!p�@�
��u"�c[�bTDY{8�t8���2�q��Pa���� ���)p�ǜ,?�4��6/�-vs���HYF}a~E���4��鉴iU����_���dShТx�w��Xn�̪Ā��z:%�f-
�|��'91"�  �N-H���S7�՘H��Y�ȓq%��;ѥ�2N,�����S�j�R�X�_�W�dB-�6�����')�:�V�ȼ��U	Fx\a۠�C,BC6�v,�K<��U�gf�J�G"ss^<�`�$}��x���.@t�	j�����l ǈeh�
���F	f��`�	D1e�G��<D�ax���O%f�1ph�G��J�Å�-,x�Bg��$$XY"��8B���BF�C&(q>	�`�'�"Ѓ�!R1!GD���싥tD�x��O��h�Y�H᚜���|](tr�ĉ
Y�i��Ψ|B6E�w���9֌�-��Y&�Uh�<)`��>�0�P�(R�&�	�Wȁ%l������3�4]��B�|�t:H~�Q�߱�x�;#Z�%�e��RH}��F�v�����"Y�1�r�Ïlj�|��޻O?z����B)�<Аf�$a���4�F�(e X�J��hOt-i�lS<a�Z�ˤN�&޶A�'��#��'q3"��f������&�^(`��Q��N|r�����k��:�J�d�DEz�AÔo����d��re^mk�BM���	.7�Ƥ�V�&$\�"��3;Ҏ�j3n��o�\�'<���I�lь~����- ��4�ȓD͢�CC$��hR���HN�4$ `tl[;2H�y��E����Jcb����
��b#� Լ�e�iX,�����$�d�!��YM<�2�v6�r`�ˍ`\��te�fx�hG����Pv��?GZ��ft0�2���ˊ�24z䡖.�$��b�%�ax��#�~� �	�< )T儌ր ���b@�6B)]�q.T�&�5P��()�y;��0�OHB��Xy"5���}dxR��@z�K޼^�԰��I+%I�|��N&e���ە��L��F\�rq�I�kDpYjd1��O1�yra�B�ZӠ^/o�����Dxmh��1�ղvA	hl�s���$54��=Γ[��1���5$�A�6t���by�AEl̴s<��$*ƽll�{$�W��Tk@g�)I�h��6 �8E��a��O2��T�&�?TT 8X��]nPx�rr��5%����G�)ߨ��$ԐhM�q��JJ,�6����v��(����X���C�iy�6Ҕ%�@�@�'�&}ن��13��h�FB� �(�@O>����"�h�R�n�b�lL&`k&�]�*�1�T��,��݉l
u���cAz����|I���a� �#�Ҹ(����D��BkR�Q�:�*��P�}N�4Y�ԝ��	�O���L L%�7h����m�#*�)!�$u�ʭ����=Iz 5��Υ_鲴@giܫL�����P��T�>OΡ��K�<K~�Op�5W�@;�<�%�~r���'����/�w_t��#+a��hSB�Ǯ��,����d���Op)x�'؁NaX����p���ɐ��a��%J��Y�o�8�¡M/�`�˃{y�̋0�F���C^4.����KJ�0("��8��(�EaW�8#����)� �\Ei���N)m���f�$�Sp�@�g����p];�ɭl��C�I*�v�̵\>|)���f��I�c��t�E#Wb�)�'s���$&$��s�-�)�pЄȓz�����,V;X��l�2�B�D�O&��b�H�,�yB�^����b�WƥIS�ڏ��?�sa��d~h��CR	r�rG�-���'�4��B�@R�1!���X�'��i���"M?h0��-F��U��'߈\��l@�QĀ�˅#�(2����'���	S����quF]�-+����'s$X��],Mʸ��t� �z`�'���&�$I���{5�h3�'�&8�c`��b	*��T��mb�	�'�b�9�i]� -Z��ݽ\ ��'Z��%�
�|����]��ݩ�'��8P�E}-�!ːA/Q�xĠ�'��J� ��)�M*P,խC�A�'���
��;Z��1�>3V`���'�Ha��&'I�C�ڤ+o����'��I�#��BSx�:��+z��'X6Mr��K�4�N���D�
�����'J(��q�|ı���x�d�3�'�`���5�f4��0s��\z�'�tpG@��p�p����##V���'�l��q�]8�B�b��I'+g����'�y��,�U���3pLT{��@�'�t��n�h>��`p��W���;�'�`��m�~� 3�'V�yҺ���'��F�C�p���j̙�X���'��� @�?[ed�3t��Ȣ
�'���I�n8�$m�HԛP�6$8
�'� �C�

G}�|8��\�MLT�y
�'5.*��пI�P�p���G�0�	�'����a\�À)��\f�P1��'g�j��ܵUjHA�bjJ7#�ak�',�	�0	�8���˕Z��
�'="Y�G�<�.�;DE�Hi]�	�'�����iJ1K�x�jC/��@؈�x�'@�T�C�]
���R�G��T��'&���G�
 �,���ۄK��I��'J�%
�C�0ˎ��KF���'m������^0�dȱ��
n����'�h��щ�YI������Ha��	�'����Ǫ5*"�b@�^�|��i	�'"0$��ۦ�@���#��Q�'.f�c���t����&<� ��� ptY�O��ъ��Q�	`��as"O2���\B^���\��*Q��"O
��CF�.Y�
m���Ʒg7��D"O��B���B�e��;t��p3"OVX���2����&5f�Ph("OlY(Dl�KT�:ǜ�;�@�A"O�<��	ċ�8�����9BI:22"ON��G��<Vv�͓��M�0=\s"O��R�`Ɔ\�}��A�*��G"O���G�K����:��SY�"OB��6GL>�=�s
�I�B���"O��A ����gѿr�r�x "O�S3��,������N����"O<�7�ۙI<�La ��H�T��s"O�I�6e��aG&	�lЛe�����"O��Yf$�M�T<��`�8""Od�!���?uq���F<6�d��"O�8i��v�KP6��i�W"OR��F��'��j�i�8)�$�0"O�qf��'W�S���%T���{"O>�+�ǔ�_��,�4�ҥ:�H C"O��#�b�/sFđz�&oPZC�"O���g��?`H����
b�E W"OX$)�dߺ&����4��!��"Ov��F�Fݖ�`���5�� 0"O�]I磐44F<0 痬Ȕ��v"O�Т/�`8F$�ռa-I�"O��Y��ɨ!4Ld���ƛ+���C"OD9c�!����'�͠7f�E��"OnDyE��?d2����>����"Or�9�!�G��ͫ��Ɓo�j�9"O��(&h��GK�1!����Ԝ��"OHq��.Ƒ��S��8^�b���"O�Q��K�8Z(Y�&��?�h0�"OfA���Du&�'��!~��3�"O�Q��l°=�&�#6B�� "O����o:%f�L�#O��Q�Z)��"O��k��	�.y��CDI��L�^m��"ONq�`��#�$�#��n����"O�Yyb�?qV	"���"_�"d�$"OĲç��}j�䂳̓�\ ��c�"O��j����GC�xT�>/�����"O���WG	�|�Z�;"�Z�_�:!r�"OfD+�&,PT@�*� e�|�Ca"O��w���D�|J��,2���f"O�4rD�ݓ>�3UΕ�F�RE s"Oڝ����T=�5(b�
�.9��x�"O�\pv��>@<�lз \�;��cD"O�� �Jև8(�=��� 7�q�P"Ov�1��L�Y0�ˑ57kPj "O�1:2���4��1��PK`D�a"O�\&D3Ě�eP�q�b�"Ol �bD���9�1'K��ĉȂ"Oz�!����e�B&�({B"O�y�c"��/Fq�aE�C�%�"O���L�lJ��� P��p�"OpĚ$Z�_�$U � ?ް8`�"O���'�U���
EÜ(Gƀ�)5"O�I���C��X�1"�t��ea2"O(��E$�aSg�(V�x��"O:ɺ�L����S�(�L(��"OB�;�.Qn#���1�E6m�x	�"O���r�I�a[��y�b�i�h���"O Q��&�Z ��c!O<S�����"O� r\�p��P},��Ւg�(bR"OdQ���
�/F sԄ[�[1C�"OD����d���H'�5 *�ʔ"O���RI�}��@q��]N4`��"O�@����P�L�Pa�;�>Ћ�"OLlBŀqd2��Z@��H�"O�a�ҧ�)J�|%*` �l>�l@0"O��a�JӗW �f�[�f��yW"O��ؐ�F�w�0�B��U,t�01�"Or�K�m˂s�@�q�I7mV�lk�"O��ڔ,��O#�CF��zN�1 "O�d9�L�j���9Wc2"1�P"OЃǩaq|9)��W)A/L�r"Or1���qp�,�4 ����"O�@�i�s�ZH9l[;�lap�"O����ҵW��k�j[$&�KG"ODp����$�\y�ĊԽe�*"OH���O6]l��4nlAXY�"O�)��L:��l1'����$�Z�"O�d����0m�x�D(�b1�"O�����N;K/Y��m��Xd&���"O���`��?*����TAo��u"Ol8!��+cp|@�BRMC��f"OxSu��LԘIS1���!!P���"O�G�ћO�||X����j�Ұ"Ov�J���^Ԉ�L�'.���2B"On���M�����J�~�B0�"Oށt#�,T�,Ct�D�B~*h�"O�Ѐ'��&M��X��$�v�� "O2\+�eQ3svу0�U!4��d��"O\ICe�T-2XÖ�T���A0"Ob���OY�/؈� �0!�4�p@"O������̘��/��Y���p�"O$��-�0F�;ҭ�1Lu-�4"O��h��!7��|��R�bv�,�P"OVLz'�N�?��1xG�՟er�Ѕ"Ols�o@�~8X�GK1BhJ,з"O.0�Q�I>EIB��qƐ�"O0�p$閧p�(����?�Ҁ!�"O��@��Wjʦ `-ܱ2���9�"OR����BE���<O2�9�"O6th��ēP��l�V�H�^�B"OҩU!K��q�*2HA"O:D��f�(S�J(�r�a*N02�'}8J�X��Ќ�2�� 9{�]��'̜V�6��mt(Ȫ;���1�7D�pbR�v� ����3��p��L7D���p�S�JÜ�SA��30�2D)D��
�/� 9�L4+�A�:d�P��%D��1*��H�T)mB�&���g�#D���c	��JN ǭ�2Z[�!�Ī!D�(��!I�8`(��%�{φ�� �?D�p��IY�!�����?b��9��*O��Q#O� ����Ƙ�}䆬�"O*��ťV?�LΖR}����^�<��%��A:�eqa�Or�Q˔�Kv�<A��^Lf6]
c�N�'Ï�o�<avgC$��	�CaQ�0+�:���l�<!��'m@�c�J���d�Ȅl�<���M�<EΘ�tmT!/��]��#k�<���: �*�i.Ks���`�<���m�^���#�5d2�D�{�<�(�0/4�Ţc�έ?�D�ȓ3���6l�>&PA�QoO)u�܆�S�? r�d�Fg@��d膰)�nd!�"O�Hb���W�p�+D��:sn�mr�"O<��'�øK��T>H�����"O
5�e�a���q�f�����"O�����L3S�ɉ5�ڏPD9��"O≱� \�x�e�.{�"�v"O����_�k�f���# \~襑�"O� ��I�+d���ႃN�Lm��5"Or�����3ӌu��c43M:x"O
I3��:J���ȃ�"OHP5�_��j�C�F�S�O�\�8VB�2sfUp�%k���'��D�' ��>&��C�+�r>��L���� ���x���C�����%��[���P�a~r�ȩWbF42��2��� /|��"�玞���=J��Q��ĕ1Oɚx��N������Է-=���Jt�� bU&����W�n��ū�JQl�<i���$6�Zf�V,��#� �<i�) j­qM>E�D˔�L
V8�.M#Π�c�kI �y2��L\�S���j�����O/����4�)pk7<OнpQT=��=q��Q.@9P��'�(5�	aȐ����?+����!M	y���O@�EV2xp8�#%��i�$��I�k���2��F��_��['�=g����C�-P�y��U��`kǎ��+�jD9`!��	� e̓w������S�O^¨�R��;KF���=�X�'���aw�6H�j��O/qHa)I�$ ���]#���$�+� p�;@:�C�o�"��2O)�=�!M�/���#AK\�E3"O=3V�^��2�.Ċ/����G"O�y��Y�B"�ٹ��GY��j�"OZh��!�X<w�4fK���'�ܘ�G쐐_�d�����&
���'M�<kc*��F3�X��l�4� ��'�Y���K�im2�b�+�	~P�'Nn���a�BVx���/rj�u��'Z��{�G�b ��[�p�����'.��C�&������g#Du�b�'���l�.b@L�����0�<e��'#V�Q���"#N�8���~�
�'�ҡ�RjG&��$S-m?�]�
�'��� !��+�Z�� ՠ7�а��'�����M�*�=�$�=/Ebq��'>���%w�>,S�!�8T�Q��' D,���Ĺq��A��=A�i�
�'�b��CGی.�l��R��<?<�	�'Ò1�RnP��M��j*h�	�'n���w��26�ɃN��r^�a��'%���j�(U�S�_�u�ΐ�'_��"��=/�Riz���o�2m�	�'ވ$�r/�Mxđb�ƷX$�ȋ�'(�h�u�s��
�O�*E��'W,ĀI V����OU�$$%i�'DR�aE�I&
��A�8�)�'���-܀^�����  b���'����tݯd�0�@k�Us�̘�'�h �ۖ=t��9ߦ���'���a�@�");(a��J4ݢ]��'�z��ʋ7D�$�oϤ9?2ap
�'�rXZ3��0eRpY9Uf�n�L���'�F�8"�9��{�/˘s�:���'-tii�!L�H�GKU�	�'|%�4��?�����
�I�']r�@�S61^I��`� ���
�'I�1�/L�m�� B�����]���� X��
�pM�H*��K�&Xp�{�"Or��	�9�J���JS*W�&���"O*��Q���0)>�iƆ.Z��<z�"OX��q��<vߖd�"ˏ�_��i!3"O H33*�V���5��/<�В"O*`��l�Wڠi'��
#	�B2"O��@6�Lhu>��U�O;Z�Qѧ"O\Y)� �WGĢ4��"Oh��p"� >V������lxB"OMIc߄0�����	�^XF�j"O��Ǎ�UP~�s�%�E�
�*1��" Z��RU"����6._?Pp��m��\R� �	�L�#��1�x����e���5k_.I�&�9w&�@�ȓ>l��EfL�n���aB�Q�lh<��}n��K���@:E1�D�P�A�ȓT�,����e�H��P��.,j^��t�nl��+�� 8!'�)�~̆ȓ6.>0B
Ĉ?��1�&�['9^%�ʓr
�(LZ33�Ĩ𢅏9#�C�ɧ6������9��-���qSvC�ɷD��aۇ��I�SBL�V�LC�	�l`,M�W闞i�������I�8C�I	$���h��8Ann�X��I�i}C�J�jT:�m�J�t�	fD.,��B��
-�^�zC��I��z"�;��B�	�&��PM�e�;AF�A��C��>�@����K�]-�Lq��L;95C�	(P����R�Ŕ�12G
�4��B�ɸEU��0���z9�Kp ȭt�lC�	��X����-��ƸU/xC�ɣ8�F�*�G�#&ߒ�t*X C�kT�dz��@�T�Z����uF�B�I�C����I&{��[e˛�d��B�	�+6�@WMXc��8(M$B�I2r3�S�MN�^�]�eR�J8�C䉏x�P$���=�j�aV�G�iQBB�ɿ}<Ĭ0���cG���,�k�FB�	�b�L=�pˇ��i�J3>�C�&{.Qsd��|��p��l�l�dC䉦=�
D�B��+��l�G�~�hC��R��b'�'��t�c��X��C�IP<0y!��IJ���Х�\�C�t$]�1�a6�Ts�N�\:C䉙zR*�)C&�0,��CP摽{	ZB�	�8B֐K^YW,a�p䄤=�LE��'}^]r �
<3ܢ�I��:��9��'K�;$��~����VA`�f�(	�'�� �کf��*[�:,�"�K�<��.H�=_2q��'F��	��A�<��eî*ўࣂ��Ix�����t�<��"�.X�@uҖ�P3+��Qz��x�<ї.F=h,�Z��ѦK�Ղ3��v�<�	U?TuN�(���b]��j@�<�h�4yZp {��+lW =�CiK~�<�ףg0I�I�9/�H]�C	�P�<���ĄMт2��L�
��x2!EN�<A���i���E��( ��6�n�<���Y�A�& ����L4���@j�<���	m��9:"�ȉ&�`�j֡Ue�<%e�V���d �-�e�<��JN8 r,�zV\!A�i�w�\�<q��Y+u��tr2�T�Z���&X^�<y�Iŕe_���M�mw����X�<� ��H��3����|v@�2"ON j�SSW��J��\�����"Ol�RfH�y����I�('f��3b"O ��ŋS*q�T�k�ŴZ�J�"O�1r/ߐg���3hTE�����"Oʱ��O^�%b��B�	�@��+�yȖQa�Ӄ�ġ;1p��n(�y��'~n԰��ǑE���R W,�yC�J�Dp���9f$ G��9�y�._:_F���F�7~���ק�'�y�o5TF$	#��,`(GU�y��/:O��Y!�C�m�D(DnW��y�
�%jɰ+�`Q!Y�F�hDbݻ�y�H�U	P� .I�-�"�R��yb�ל:�F0"P����.D�*���y�0б5@�<W�`��Y�y�Å�yK�͉�&�3>��acR��ybn���}1w�\!(���QK�?�y���	/���2'��%M��BB��0�y�� 6d��{��#C�4)
����y�&T/Ldt�s쀨i�Α�1��/�y���,"zII����x�"!Ԕ�y�� @�xa��|P|�e��y�==K���c�>xm��B� �y��WO�@���9s�\�R��hf�t�>)�C7*R_�I���y�R��Ou.�5�� 1�M@玍�x��M�0���][�S�')��,��*����I�<�.Q��O��<X����H6"�V(ۀҘ@ z���+Εl��`+�N�r�S�O��P��)�i �IX���"�,1��<X�a��&՞xL���� 9tI~�{U�׿�'�ҹ������Ɏ���qѲ�El�b�Z�����	&�P��?���J�9)��qI�Dֵi��d�â�B?qG�"���h��$# �S�T��L��� +(��c��<��ɣ,��y�A/������5��B�	�^��`�f�ڝ8�)1�e�-y�"=���T?e8@F�2M��r�MU)%y<�J���OFD#�^n?����Nw?a�So V�۱��\�.�Ҁ�5��P�@�y?e�׆�~����Z�t`S�����)	G�t�`J6��^8NHj<�ɧRh��ᓣ-����^
��pSՂ�4[�"<�ϓ,��4�#ś8>��Xrh8 �"Ox;�H�=�L�QIJ�3p�����'~A��x�lC-X�0 �aV�?���T#���~�!ـ��O�>��gi���Dc٭ n��7�W�Il-x���ɏ~��p�#H�0p���['��{��\�?If�3��5yQ�s�2��T���fc��U�d31�㟒��d3��D>�"x*a�[�_�`��>�D�7����O�j�����	<��`־&G���'���@p��S��� !vT�	I� ��j��1�Y�����&D�!$3�M+�E�v�Xq�F�~��i������ (�
ʤ��;H�I�u�QJ]I�t�#e�A�s�B�I�^�ht��eގ���kg�@�*tB䉷\b��	5N̔,%�M��*YRB�	4`�B�aU�ܙ��F�H�vC�I�VkA�a�_`_�uX��
p��C��+l�^Az�狤2r�"�K�?�C䉼7�ܡS���1M���fm9�B�I'=PP��2@�y)H�ti�C��B�ɃFt�8X�p0�,[�OS%YVC�I�,X����:j~p0R�ː�a�*C�I+^)�a1#�	�i�P"���@�B�I�<�L��	S
c޽�^�w^B�ɔ4�8|a�E��04��K��u�ȓ+V|�Q`\W�u��	ΝU|`�ȓ�,����>y�\lV(�e�����S�? Z,�d�W�lڠ	��� ,�b}" "OTT����$E4�&��(:��Y��"ON�P�bI�@�0{���"O�%�dK�y?��#�
�89o�\�D"O�`�ȓ�T�F�	�g�#0��R�"O�]K�!3p�L�9C��+�^a{C"O�}Ȗ���R�$r�U�����y�˝ M�(���KZ&��J3n�=�yB�s�0��ӫ�����Ab���yE_+M.�m����{<-q��C��y�[/!���!�*��}���(�y���KA��pĈqP�Y��cæ�yb,ƧT��M��(�=' �a�؏�yR�U1��0Br��J7���&�\�ybaV�+.N����@�D��L�u�2�yb�4-j�8�@f��n��R%@��yB�Z�v�X�`��]�2��!hO��yR��6$g�����F*P���K�eʊ�yB"��Z�V1R��6D��	�D�6�y��Q>s( �����!���ycP�A A�  �5zc���T���y�G��?�8�Au�I�[� ��Cn��yr�
W�De��/V�V4!��]-�y ʯM_\ ��Yv���R���y��о��{���?~���h��N����p>!��Q�4�$����< Y�{gi�R�<ٓ�	1F�Z�L�#a���x�<yG�Q�q�Ժ��98�ب��#�t�<�7�Y�m���f4ao\��R*�l�<A�mǿC�0�Y���X!��(�d�<����*�`Y�f�t���ʀ@@`�<�eI�BRU�qD,$����AT�<�G�M�!�U'(d�5*�D]O�<!!���� �ʦ\
���d�P�<�����'[~����O�h=~ ہ�T�<��	��Q� Єd�0=�`����\Z�<Y$
�VlVb�Ȩ\�Ԭ
���Y�<�#�1�����]y�*!nVS�<yf�T�K�zT�5�[=@�zI¥Y�<�wMC�6�xD��7p��:4'@W�<	�m��`.��  2~�IAm�Z�<A�r8������gа�j�/͓R]!�d8*L|٣m\<_皸�eN�9xK!򤗑fq�Ah�d��ܠŪ���0�!�d��xx��qK�0(�)3D�=!�$���T3w�
;t�E��i\�-�!�_/b�~� .�<n���2hR
q|!�dJ&�>ݨ��9�\hU�R�!�ă�d����õ+/�QJQ��!��ɈXi��Z���Re�c�!�F�!�k�5U̅�D�\�!�Ԩ�Vb,��P�:�� w!�@�uF�(">xR���DT\�!�"O�D�$e^"L�REOI�4d,M3Q"OZ�(w"U�1~͙���^K6���"O<x��.Y%x	��P ��Z��a�"O�����޺M��YI����,��"ORe+�$ �i�����=w�8�a1"O�u���V)D��H��ׁP����"O�=��@S�Gd�P6,YL�!	�"O�@���D�F����A�W�|	�"O����p�����G�`)�P"Ot� B��#&0)�Zi�J��@�Hv�<a�mV���l�	*��f�XI�<� 0�%�N�A@��˥W$	�""O"|T��>��`gN�K��Q8R"O����k�"�J��o@�RT"OT����<zjr�+!��<y���"ObU#"�!�(�&l�O�~d؁"Ohrv�$#$�A K�4�"O0p�4�B#��*�l
�^��}C""O$۳O�#Ծ��w��G� �r"OjD��b݃Ø���
H$S��Q��"Opy�/�(�$�{C�|M`y�"O��1����@��\&F�/�8:Q"O�uHr�#Q��AG�E?W.bX*�"O y�˔Cu���2%N`^�Je"OP��Ň��&�2�;�#��^
ja�"OL�3.ܨ&�;���-c��a��"O.�B�
��[�츋�M��s��@S"OP�{tc��9��ڇ쓧%�h�"O�D��
8,�z����ѐH��iu"O@x
��W�a$�9j3��&�xP�"O�t�u.@�p���h��(��X "Ol�$MZ���d���D�u�~A8@"ON}��b�<{y*a��H@�pK0��"O>}�beƓ`h�Q�fU Rㄨ��"O� HSmN	R#Ȥ�Kɋ}ז��U"OD�6�A �Ra�0�@- �* #q"O2�Jcl�ڜ�h�o�:ݪ�"O�:p��z �E����!^���""On���ø/�MI�+A|�c"Oz��\26��R�o��9�����"Oj��%� �:e� ��O�!Q�"O� ���	�A|��"�UO�\2"Ozucf�"�`D*uL�H~�DW"O�E
4ON�"�4h�K�n"DJ"O�8@����e5��� h
vE�x�r"O�(K`hT�b�0�"��M�I�6P�"Oq	C�b�e���H�4B�"O@q�+�7k�R�;.��I�"Ob��T�T/��i�D�8�Eٴ"O�tʗ��E�:l�L�V� A"O@������+ۂ�Iǂ*#��Ap"O�ْ��9�8 �뉺+�~-0"O�T���J��a@�	��9�T�yR"O��C���G��4x��X�t�hC"Oj��MB�2���B�)��ܞ`s�"O4A��'RR�dP�wITv�����"O�X�W�^t2{�+TL�"OXZ��:
��AN&&{Z�@�"O�Ո6H��PcZ5C�4�^��7"O����N�d8����.�">�fA6"O.H�꒼:c�\����_:"�"O�lC��H�����T$?���"O<��H�H��bB�V��h��"O�x�#mD���	�ʌ�S��U�D"O,��Gَm��ͻ���K��"O���o�O�N�YF��=~�"OH���d�7~Rĩ���'M{(��S"O�����º=l��ti�d��S"O�T�U�S�zM��s��O5����"O�EAg�ɛ{a�WI�c����"OJ�Q�_��b��VGýH��,&"OZtA���U�J�x@]��Yq"O!�`P�Y�p*r������V"OX5Y�h�,34,�Po�p6}C�"O�#"�
V���H��w��;A"O� Z�rv�S�j�� k@"�6�>MS"O$�&O
15����@ۦӠ�d"O�-��	������@��<<A`"O"<$Ұp���"5��BG>K�"Oj4��E�nB�(�3��+T�0c"O�8�EX�Z~Ac���M�b���"O�p�kH!MX��a��H�Jm`B"O����N�h�b�>gwX�u"O���Jè���\�{$xc"O������4P�^ѱe
-PH@"O,�Z���_[x�@��\��.؃u"O��@,�6|�~qhV@�*�څ�C"On��A:�%��9(������yB��
-���;׏_��	#L���y���b F��p&�!�������y��1��\�%%Ҧ����բ�y���9K�ɠ���|�T�G�Ρ�y��ձ6prl��eV_~���[��y���tszE��5!R��唸�y&	1u= y���R�(A��y�$�2{�:iWb	�zt%���U�y�*F,���#C:y�>E�����y�$�;�VT@G�/o�U!��G)�yB�K����ԉ�h���g���y�'@
#`��ψ�o6洢����y�HU���x�P"t��%���y�`�hD��dF�'L:,U�k���ya	�^� P�@�A��%BC�֩�y��aF��! C�;px�ҫ_��y"(@�	0��a Q�9\0�����yBM�j%\@�ʁ	+.� ����y��M,�
)9BfXu�q��M��y���$@���q�`��`�6�y��t�6 �)͎;��q��¾�yB��]�NM넩GF���P���y
ږdAR�as_+O�Y	�&��y���#٨�I�蜏B�~�Р�ʗ�y�$�0D�0�H]8[�1Z%N��y����K9<ԑ��^6)��Q�C��7�y2�_=��4���X<6�`d�[�y2�=5zf��1a��d<DC
�4�yB��	�څ;�����B*�k\3�y��^J��-#�G\5�C�� �B�ɢaK�!�ժ�<#A>�Q�F�h�B�Ib)��Y�E�zqlYqN�Y��B�I�9���f�1e��� ��Z�5��B�ɈP>�3"$4����ڀCe�B�I�j�M��D8=d�	�c�>��B�ɐr/���i�iB�Kv�Z8p�B�Ij�I���6*�"�������C�=������8q3&�&�C�I�kwd#E@�x5n�b�E1M<C�1{�r�7D7
�!Pƃ �TC�	&p�a�`�_ �9@���k�C�I�!�x �   ��)�m�2��B�r�`B�I�@Ί�
6H��>��J����B�	�� C�#4s�M�5�?`��C�ɺ(��0Pq��D���g����B�8>�Z&˂C��q[u���2*������ ���n̼����{:� �3D�4�7�\'	�>!�p`̈́/6h�B�.��ȟꀁ�U�o��Y�eظ)X���"O����?u�C*��,w��c"O�"��I��,ɣK���I&"O��xQ��66��K��[ ^�Hd"O�1H��_1/r�!�	��(�i"O�i3U#	'(&�u��I>sp9��"O����g9�R����#�"O�=Y�'v5�e ���=k��$"Oj�釡K�J"dト��f�Z�;V?Od�:��+��� ˦C�%3�H� j�6s�݅ȓ5�$��B��'��i��u��U��dK�#ЧU�r̻ ��y\Np�ȓ��M�%��+m=4|#r�S�0+ ��ȓ��y�3GP<����i^�R^`��8}��X����u!�y u�[�od~P��-�f�qA�P	X:�2����M��?hc��C�L�puBB'�@~����?9Q�p�b���"̃����ȓ"�=�7�^ܘ\ֆW� �Y�ȓ(�TDJq�H��x̹R�Żh���S�? ���S����l��+Q.a�~�S"O���tL�)���r *�+�����	l�O�|�b`�'1�r���Gh����'R`(0&���l���y-�IOЕ��'�r0�Q3cT��2d��?rzP��'eE�3j͢GZ��!�4�&5��'�B�sWC�	r�4@��6&�.Y�'ۨ���K�@�&�{�l]��4�X�OB�=E�	��/T��)�
�~���&�y�!�=S0�K�#��}OR�	6�yrcɦQA�#t��w�n��!H��yr ��Rtji�;uhv8�/�=�y�H�0��Q��	4g��a����y2�,6�8����^���C���y�, E6dD�Tf�=mWl�Z���2��'Xў�����s)�!M�H�r3�\�/��St��{�O^����N�S'��i��Q�
�'C$$��N�)���xT�ݫ:�b�����Q���*r��:^px�vf�4"�C�	�d�@@4l
�Z%�6Lɓ��C��<v/| �@Z�5o�}X����z��C䉯@V\4#��0f�.�qE@���C�	�=��Sie4�wM^(+�C�ə&TU�΋-�ܬ����"	�^C��=m6�0��t��P�'�*JC�{�ĐE�+[�]�c�>m��C�I�*qș����P���J�qe�C�ɐO0���ˎP9F�TKš̸C��,`>�� P� �*��ǫya��<)˓8[pMH@S�_����J���ȓK�L�#��-��i��E�3��X��2�Q�����(ԯ�-�DɅ�z��
�遟D��L�0�

_�$�ȓx]��0F
N�K�� y�L���M�ȓ(f�R�*_�Vm���ԹE
(�ȓ$�n*��),�r��`�!=b���ȓ=�x�d�8Ta��	%q�ȓrx&�p���x��xCUr�����{Ԫ�H��F� ث`�I�f�u�<��a�%�`�DƷ>����'Ɍb���=1���'G4Q�So�P]��1�Bb�<a�O��0sů\��X�p	�a�<Q�́+p�ڱ�0]�Z��@(�^�<)�
�o��MPʝWj�zn�F�<�B�:	��u����9�(TC�<i���� �,��4��a6���ևS�<@���E �1���f�%��q�<1V��IJ�p��$$j �hE�<��P�B�z]�u� s
E��L^~�<��@�=�h�`�бļ�&��N�<��Z�~�Pp�WG$��0p�b�_�<��`�
 �F�R��N�>ކ�Sv�_�<��L-[f�x͛t�z��`*LX�<��kI����S��6oA&]S��R�<�;^��Tb�d��6���A�\P�<9&`N,7��yBE��%R޵B���w�<����&s�:�ǌ��t���ckHr�<�1)P%Z24��#7�h�� �S�<y�@Le��j��P6��Bm�D�<1�璡&���H���3#v�I bZ}�<1�ϖ=�� 
��Y->V�����y�<Yi�j��)�KR&=Y模C@[a�<y֩W
m�Ը6F£v<m�3j�^�<!s�0����)��)�Z�Ad�Z^�<� P���
�c�"=K��kd���"O�͛vb]�ĝ8�aҘ4aL�	A"O \��B㨴��`�062�1"O�i�S�c��(SeRrI���+�D�<�����u�P�J����=/���� �x�<)�NH(\ �a�"c� ���p��w�<�4A�T��)ֈ�%)(���ƅZ�<1�G��#�L��k����`�[�<i o�" Ĩ=�p�"@� q�BY�<Ѷˎ��aTlM j~�c�IQM�<�f�.�hի$Ĝ�&7��A5��G�<٧ ]4R�p9�5N�GH,��"�n�<q�l8mZ�Q��
�0l���Wg�<�Sb�-+���	������IK�<�0�X�x��+�����'GL�<��gb'��S!S!s}d����K�<q���p���cR�O<�Xы��MD�<�t��1t�X��X$9��UU�< �5$Җ`:��^P�֍X�#N�<$M7���%J�F�V�BNH�<�#j�$)����	��H�@|��c[�<�d	�{k~�n�<Ǧ�Q�iS�<��D�Q���3�CA�
����L�<C�R Q7Bȓ��\\���H�<��4{SФ��f�;-o*-�w��F�<a��ތT�xRm�5S�!�uhXF�<���X_�8ؠ���$(:��F�<��>s�h�� 9P�vT]�<����%���U	^�@Ī���\�<��㙐g�h���� �>��m�Z�<	��B�a�D� ��bA`R�Y�<y"�_x� +�OL�$^.8@��U�<���EҴ�!�C'�քa�S�<��bK�~�̭B��y
�|[Ҧ�N�<A��@u�Q�!/Ɨ�,��ԢL�<�&��gu �5n�3�|�
��N�<Q�ӗ6I����ЊC�l���`I�<a�nFwC�d�&m#t�xuO�A�<�0	�6�p���N��HA��p'��C�<��+o�@�jB/b�n�H`,@g�<Q��^�o�>��ݬ(�IX`Me�<4於��tI��\*f��`���`�<�B�(dm��L��*R��ɷEKg�<�'eڎ�*�9s��-FIx��"Gz�<Y �A7C����N��x]�W��z�<�w�P��M����M�f�9'�o�<�#�x��x (?���C�l�<Ywl�$c��T��;EDЭ�C�_r�<�B�g�(���4:�,���Mp�<��K��V>ԩ��A��w�0$ـp�<its�N�"�dE�W9�!�7 C�<q���"r�]�&�hta�҈�T�<�C�M:���r@F�3-a*��P�<��Æ5r&i[u-&*p�1�4�KT�<ٲ+Y�(��t1����5)BnPL�<�P� <Q�1�Ʊ3���� J�<)i������d��L4;!�DA�4^��[�bR�$��ذ%"[6<S!�J3�M�ŏ��=}zm�U��-;!���7�6��桗�%d!# �ϐ]9!�Ĕ�,����)���d�)!�_�x�R�w&���,�� ��!�$g*P���֘\�a��띙cN!���< ��cFɓ�p���2����!�� �p��U�r@��h@�Z��p�"O:(�T#��@ �+��H���2�"O�XȒj�5Sl(��'̃c���"O�$��q0�{Gh��H�0�ұ"OF����f�J9�@9k�"O���"/~�UE�y�  �"O���*��x_F�C!�B&/䪨в"O���)�����g��?��mRq"O��ґb�<j��\8h��{C"O.���J�;-L"���l�AT�H"OP��bo9k,jŻ �L�&�J8Ic"O�u���1:t�m��%�'���a6"O�����?-���h��X�@.��"O�ɨ%�ƳI�0� ���8v��"�"O���Q)5������R�G�N�e"O岆&^h�hp�N×d�P1�"O��F��@#�{SطD%��1�"O<��HՀD���UV�Y��Kp"O�(cv'Δe��t:�� �c2֬��"O��{�◱h�:dsc��V$�I�"O��ha����͛W/À��A`"O&�)��קV]hࢦ�\T�!�e"O�5�G�^� l%�I֫H�� ��"Od����}�1��#��
�"O�jfF]1d�Ĩ�b�5@&u�"O¼���N�u= U��=?zh�f"OxzR�q. �q�@�1�a�"ODZ��*�y��ȕ5���a "O��N.$���A`G���r0J�"Ob("��;��8C���$RpP��"O��I�LD�D�����%�Q=8��"O P�2nC���Dc�$ƐwJ�Lʶ"OhȪ��X4��B��J�,@����"O�y���$T^��z�ك)>6�s"O$Xi����B��D�`n ����"O$!�ӏ�E�V�0��ڪ�x�6"Ohv�і"�ĵ����q��	�E"O:a��H� $݋�E��\�� �"O���!��P��b�#�Nٌ��%"O q���$Q��
�s�b�U"Oh�3g��_�j�	���I�.԰�"O�PõC����H:O{̌A&"O�)T�	x[���3OAB��%�D"O~ hD�Y��i1��Ɛ=�:D�v"O@|��G" �X,lIȁsG"O���	��F��U4y�z���"O��SN�>���1i�{���
�"O�i"ř��r�@�Q� yF@��"Oh�r���9XM9�Hǧ1r8(8�"OF��ʓ�`�(����f$5�'"O�Y"f��!s� ���h�fd����"OpH� Bi�՛F��x�X �"O`�4��iwVX�=ؚd""OFY��ߑ��)��, �����"O�#!��X=hu�UJŦ��ܻt"Oԝ �)��'x����ьU�����"ONi��� 2Yi,���'F�,�J(�"OH�[FF6~|4��&�$�
���"Oz\�^0tE4щb���v�4���"ODHB���,/L��=~��ES"OI)�G2}l�DKȼ~��:7"O��� <O��<ȃJ�bS�5��"O�����S	t[R��i�d�8�"OiH�k@?8�4��E�>JU"�"O� F	;$/�6V֡R��lY,�J""O�V�:j���
�Gx��q"O@`CT�N�(���ʒ�?R 0�x�"O&��#�h�4E��&��R�|C�"O�i��^�0�S�&�+2*Z���"O my�V �l��ň*�	H`"O�ݐ�

ά�ic�Y�t����"O|xK��
2JJ���"���ų�"O"��b)ȩ!2J�3��	�"O��W��lf���)���b0"Od��Q��X^F5���V-4�����"OhqH���S��pY��8��̉�"O:H��`ɭY`С�R�@:Q�����"O69�h@Ԩ�Dʽs�p��p"Ox�����Q޸��	�K��8�7"O���a* ~�:pF�0���s "O����'ZU�Fy����:��1��"O��;FM� rP��b@$��"OԈsmԆsɠi�W��-=�8�G"Oꤸ2�R�ST���"&��I�"O�1�^�-�J	�$ԂV��}1�"O�ٲj�9D�|���F�y�$) �"Otxj�/�t	&x�'�ڀ2����""O�x0����k(��ZCP�nԼD�w"O����J�|Q��b�*j�	�P"O� ��/��!���!ŅQ�&� �"O�J��CW��ay�/�@�@�p1"O����DrW�U��N��e���Q"ObP�k�!��1@��#��`�q"OJeрa-I�D�cY�R����D"O�8�*��ua��S" �2c��� �"O�82D��7�̪w�8�ԥr�"O2eY�'�!#
�H҈׋L��p"O���� g�]Z�hY2���a"O�1@wH�#)�<�8�m��!t�z�"O�MiW'��Rٛ�G2"X�|K"OV�k�h��z��EE��&�`���"O0�f�	,��@��x� �"O*����M�#^� T$Q�:.qk�"O�p"ɛ�8�AXGJ2e�6-I�"O�T�@�"C`�d)�$:h��"O�p�V�F��u�RBE"|�� "O���H�j���96�ыt��#�"O�)z����>��0x@�L�?�~TV"O�EqB��Yq��1����a,��"O|�����'G�������'���"O�� u�D�/w�r��Y8�x�q"O�pv�ǈ�p}:gUZ� 	S"O6�� 
��i�e#teA)I�\��"OL�C���0}�����6��r"O�-)F7D��X'.�%:�Zq"O�ti0N��8^e�r� �i
p�RV"O4�X�ӈ[j�� EC":P.��"O6(B��Oo�Dar�	=&�����"Ofmq��J+o�X��P#ޫ �\��"O\��$����	Yg *S�� w"OJY��� V<�׀�����"O�q�՜X�*4C��8,�^�5"O �r����,�$��-� <+��9�"O�@��'_�P��,U�"���a"O��`+	[,uƋ�4L�:�"O��KK+@cD�FK\�#��e"O@��	%��XP,>8�W"O��hv/���}v��5B,a�"O� �	1�(�
U9��n�[a�d"O���M��80��,�%�(�"O�X��EG�^I�G&��`"O�ܒ�[6$�����T�v����"ON�Z��҂vD�t�K�i�p�"O��01ǚ�/T��׏<"u�"O� ����Bm�� ."9�"O�Py�HΥqu��f��d"�$�"O $�/�g����)�%����s"Od1Y��P�u��#CѾ��"ON@���u���3F@����ju"O����+P\ZC��[�Bu�@"O�q{����M2��3dL x�"O�}��坏"��cǂh&d��"O�31D���R���N-!�8i�@"O��8�L�?^ �Q`�!�M����"O>�x�F��P\Qe�� &Nqa"O≀���Sv�D���VN��"O��bdDJ  ��m�7)BH��dA�"O6����QIL�� �ަ,xH��"O�P�ċ�H���i�oʾCs�!#""O�;A�՛V����NR=wv�"O�]��� �@��f'>
ޅ�!"O��{d�����2f�@� �|�"O8Ȑ 2KS8���Cߒ:�Ht"O��C&�U8`K��֫�/
i��"O�	c1��A���f��ԩ�"O���mԏ�"�`�
�k�B���"O���!���p]f,@V�*&�{�"O�)2 ��Ep�q���%
DP�f"O�)q�H�;hNNt�H�-qҥq"Oڡ��+�y>M��'�#6X2"OH�b�E��1�6D���$K�Q3�"O�ͫrʗw�����ʤkK	�"Op��v'� ��cDa�7
|�"Ob�Y�!Ր���Kc�ѱ| T�"O�����\&�|\;�����&%0""O�m��@�9X��Q�Z���Q"O����t�h�UFj�FH��"O���-�d�ν1��\=#����"O �J��8R^���W� 
	��4"O���FD�"� �9G��T��4"�"O�q��I�b�X�A�..�{"OT b@@��Y.d�q�gG�~�&A�"O��q��Q��AhS'�����!�E$D��B`'S�؁
f���]^\�0a�%D�Ի�s����E��	S-����%D�8�Cƙ_SΥ�e�*"�d�.$D�L���=U��lm�?Q�"I��Y�<'aĽa�R��d�4�:Q�aHS�<�3iL�/j�c�4P����A�	Q�<�fkU+R�Vihv�ߊO�(	[�k�F�<q6��%�Fy@R
V�C�N��Ǣ��<�C�$g�	�gN�y}Y��AC�<1������t2�E�%ff�2�z�<�QUV���"��aQ{�iv�<�Bh�`5�t"`Y (��8�t�n�<aƯǢI܈��+�2Ę �#JOB�<��#P��M8B��8�,�2B��y�ɛ�/����d�^��msrBC��y"�̣Fh^����W�P����P��y� ­Z�F}3pe%C�.��⥅��y��9z;��
_�g���Ҏ�7�y�C�:e]�I�IW�Jt\L�RIH��y
� 9��!�./ ɰa�/_@:Q�B"Ol���a�3d?ր� �?\Qx2�"ORP&@Ӗ�|���	'xE���5"O���C��hv�p�+qCT�0"O}:��Q�]�n!�/%����"ODԈ�g��,Ҥ�@b�U�6&\E��"O8}�!�M�`��hR��_h� P"O�4���nE�����KR%�a"O-��������E΀"O������*`�<�ф�)B~}*�"O����iӓd����'��V"�� �"O�!ky���pЃ�+��"O�p��	.q��y�����)�"OJh��<8%H�R�.�7<mZ�"O,dx��4������{ZIp�"OH\Z�/U�G�+����fhb"O�EsCזX�c�]�l�Y�"O���f����"���a���Rx{�"O�u��]f���Da������"O&��k��_��� 7��)q�"O�9%o��pU�G�;	�Ip�"O䨀�On��= q%�.��F"O$�-��V��*�T��hb "O���m
488�`�闝�����"O��k�!bvtܑ�\�2sj���y��ҨNnl���Y)>~�å'�y�H�jSX���'�$/d�%�5��y2
�g�>�� a��#���ꔧT��y"E�D�0�s��� �T�݁�yrH	�3����Z�`���3�yB�T0k�{�n�55EsD'F6�y�j�gfH1u���}5�أ��/�y��V�Vd��2�d_�$<��s�Q5�y���mb�������Q�$�RnS��ybϔ�R���M�4��=�@��y䖥~��P���%��j�,G!�y�E�"k{^�!���g���*�A��y�:Pɲ��c�˶�F��yB��.�`sJΈ%sDh�թ��yR�0s���@�\�?t5�����yb��?w�4x�J��J���Ϙ��y§w9^��E	��A�'A6�y�D?``�C�H�ZD��`�ď�yi�?.@��n�Q
~�+�)���yR	b�ҥ��M�@5嘼�y҅ ��Bȣ��I���0@���yR�\SW��!3W�H�m�w;�y�H�%���dm��A�����Ǝ��y2ɛA�����=�(��3�B:�y�f�#Њ�3M92��j�l�'�y2D�+���
�,�*�f��@
N�yRښ?0:a��Ǎ9H&�cm];�y�� �o�|Ţ !��Am�؉�G�<�yR	�����Y����8ubhAcÇ6�y�޷�ĥ1�͜�7`�#3B�y��S>�T����3��3���y���ŘC�q`�P�a�ȓ@�H1��(Z�O5q�����Sg<����ſ'Ǻ����y�0�ȓj��ģB����h5@�'Y���ȓH��L���9H���ck�&Wa>T��Q0���v�@4�1�ǈ[�E���ȓfb@��V��]O��u��>S���ȓ��W`�"}hH��F��l,��S�? d��C��j����V�@��a"O�4hwc�!?���H$W��I�"O�����:,ٴ���C!R��D"Ot����͵5 �W�0P�����*O
Л��]�hlZ%���T����'�DK�	��q8�g{�yi�'���E��#��$���7zЌpk�'<hQ�o�B�biy�æk2A���Z�I !	�T>J`� �3l�����{���ΝX�B��v�ٲ~�|�ȓi�e�$��:�L�R�ܤ��P��3��Ȑ/���%I�ȗ%he`�ȓ�:$��mȧIbN�P��,C��d��o�R� �ěR���x�F\�y4le��C3p��3G-��Y��$A+?�p]�ȓ8������UOXyRe[=>����ȓKٜɹ�J.���5l�7H��܄�u�i�7*��in�ѩ�lX��z���ּA�'acԸ	ug�'P4��ȓSʘ��w�=X����`�'lzԅȓi�X�Yv����dE�l�F��ȓK�D ��MջH�x ���8�"���m4�y!��Y(E�1�_�y߈݄���\��ŪY5������,���fF�q�4FN)�Xq�'Fخ>�N�ȓ+1ZTۇ#L��E��+�,Xk0��ȓ>z�u�'-Ήe؞�B�,It�-�ȓn>��ѕE�2Kΰ]��Y�X^Նȓ6;�x���%a_��"0�0E~Նȓ7p�7G$lu�vd̢^-z��W�L,P��1�D���߉(<�!��N��9�-�3K��1�5C�G6Їȓ,�Px�PD)�~�� �O�$�x���fH��2E�r�^�@3��"@Y�ȓ@�bi"�,�/�|}�����v%�ȓx��M0�fCT7칢�χ�`M�ȓ8*�4aט`*���eW<c>i�ȓ��u ާT��@fb�:Zh�Ň�eA������ r�6I��������ʓw�:�Y�o�.��y����C�I�
�Np06K�8C�q�#*4��C�-:�r�N�"��QIJ���C䉑�&�;S�]�P(�Y��[B|C�	�s���,ǡT���J�K� �XC�	=!j���EƁ1�P���S$+��B�I&D3���%LY ($�Ċ��CB�B�ɗW� tDi�=��D�D~bC�I�5B����+��{��O�XC�	?�6����^�0)��̩g�C�I	e���ؔ�7�{g��sR�C�G]r���L@)��
`�J�zH�C�I�&�D�GLjB�[	�C�	��"�)��Щ(��G��w�nC�	:h22ɹ�&U�`wZd2��H-FC�	)ኩp�`�+�:�C��Y#f.B�I�-Q���5@՞��25o�58��C䉭Ҩ��K�7�&1�R(ڂ�lC�	'B�z����=V�=a�]+y�dC�I�b��	��%T<!�*�'+Lx�B�	�v!�pc@f^�O.�T�Viث��B�I�0|T����?�`�3�e%nA�B�	J���J;|vVh/�%�nC�Z�|T�U#\�$�H�ص
c�jC�	�����`)���DP���=9C�)� B�`#��o|��ja��VR�T"O�@y�B��*ԁaN"g4~<�f"O���V�`��v7"����"O1��k��'��U�aW;��Zg"O6�񒄙�"�
�f/E�N1�c"OpQ8`8&.�3(G1���� "OT$���(團v!��Q:q��"O�����q����oJ/.H U�F"O�H[�+N�sTĥ��hG
X/ ��"O~q�q �&(��ɇG��.,�"""O�Ax@��,CN��'��l+�Q�W"O"-������m��F�0%��c�"Oք	��]4�����gS&e�V<�"O<`���'z���b�S�Y�4��"O����$��t���a��-�p�h�"ORh��E��M��	J�Ĉ�#�"�q�"OR����-P7|�WB�j� )��"O��q��G.�i��@�F����E"O��q��1:q���P��fuV���y�+Ȟ�CN�~ �iق�׍�y�ǐ,?ܵ�Mܨ_6tZ�����y"�<\?�D���1)��Pҗ"[	�y�A�˚�PG��k�F���*���y�Ǒ&b^�Z��0e}<Yk`�
��y"*�B$"��,`�T)C#���yn�[_J�p�fP�X�vȳ2�A+�y"CD�A�B$#v��XA0��BF�!�y҉��o|f����]��ibE�ՠ�y"H��T�R�!���]z�Q�̀$�y"O��Z�I�cT!XN���jǱ�y2J&~�p(C�Weʒ�����yb��]� �6�>-�2�V���y2�|��9d �D���c/�y���H� ��@��V�"�O���y2gN<�@X��?/f ����yr�E�cenpׁ̜	JE����1�y�ГF�zQ���Hk�lq����"�yri�93�ֹY�b�Qf�Cӌ���y�� +�� o��HP�(;֠��y���!h�Щ�D(��@U#M)�y�Ŋ6u��Aq	��d��k<�yȁ�}d�p3��~����$!��yR�\������MH�Pŉ��>�y�M� �^Țw�M8Q� �9�=�y2�&*>����\}%rm�����y�l�l3�DْG�v�T�+����?ٌ��S6 m"D���N�Х�A��X�ޅ��}��=IwKE�'w<Q��ڿq Ʉ�D�eL�	��5Kt�'3q>��L��)��+��$����J�+�,��c*�A�4�A�U� `��/�\�U�ȓ:<�5���)��1�ʖ:(2�m��"������I�Y�cI�sQ�y��P��yi҄��`�΁����؅ȓ��z�f]�2zHuHa@ն�D!����H:SJO�.��'�B��}�ȓ,u�3HF�g�n1!")�#>®ԅ�ON��KF-�2g�|Ѹ�ᑝ}�|��ȓpt�x9q-W����� ��b�ְ����(X#း-Ήȧh����pp�����^�n-�#�F=kI ݇ȓ��BS)X"x��}���0O5Z���A��`��8ҙ�u���6�����8@�JR~�L�kE�4ZQ��S�? EaCoŮˠ-�POV�a�͡�"O��Y'��\'�)�R��a�"O|�b���gM�$�2�"O�]b6����!*[���0��"O�x����8P����g�(q����"O*��VN߯�����J =�Б�"O����'��\:Z� ���^��A"OT�*R�J >hy�'�e"O�ek5���m��MJf��U�@�"�"O�9��f�@���ɦiH�W�\��!"O4�q�)V�L�����S!DZe "OZ@g#�� �\$ࢭ"O�5����1)<�0�;9�b��"Ol���Y7Kg�}�d&�%�^M1"OB�eA�%%T���9}���;�"O�8�'M9z� ɡ�"%�.��"O��bW
��BDT�5J){t�M�"O2AcQG�N��舄ȃ�C?,+P"OP=��pu%����[����"O,%kv��dD2i󒄌Q��� "O�٧d�'1�B�B �·{X�=R%"O:%υ](|��@�ҹWߠ�SS"O��!֤a���i�l�  �"O�9�"ίG����q��(�#�"O@p��G|��|)0-��L��A"Of�(�K^7v��	86�©h�"���"O.40�H�|�����N�<�b��"O��Cv
g#��s O�g���A"OF,r�v�CC�&߲P��ѭEN!���(
)�����k��j��@�!��C�q>�a���
`�h9%$�+@�!��ڃt���;�͓3HB|��bל�!�^'�a�R�ܩ ,��KbG�;�!�$���-��U�|���˪d!��c�}�5�?j�3�@�gv!�dG"Ŏ�q�\��D0
G.�(j!�$�,�JUE8sI��@�k�.Q0!��m�X��G	S�>���gs!��4� �*x��� "��9Z:!�đ�av ��i��$���3�H{!��34�5JW�E p쉶�#!�D	ކ-s3�7O��I��4AS!����<ıQ�Fwx��!�$��54D=�`'Kt:��ҋ�7!�$̲n%9S���Je����EZ�|�!�Һjނ§��5N�и�Ù�V�!�$��+4\�&�P�Qh��	�C���!�d)k'*|��ϝ ?�@�"��y��'�f#�,P�c�,���A?5P%��'Z@Zu�PE�㇇+�Ƥ�
�'��$��R�}W&xJQ��>xY��'iTD�.��Q��t;bl��l3�� 
�'�	Ri�.WR|0��g�и`�'0j�`U��6*���j҇F5e���
�'�Lp�R�]�20�0V��R
�'�
�T
P�zj���� �5�
�'ڢ%[�
�>ov�HpC�Ʌ+	�'�v+�	O�*��l�B
6c�X�	�')84�ՠ�K�p�ұ≀X�BP3�'@�|1ӌ��DT�j1j�/Fj����'}���'p���� �ͻR���'����՜9Z��2�)L$� J�'˺�xb��|���gX�h��'C��1F��Z�0I��.�R6	���� ����F�n�a�H�#�2y"O��I�#� �&�?T����s"O��ـ�,jL�Q`���p)�"O �� ���i���AB��#Uq���s"OH����ܵv��]QdW5M>ep2"OH��%P�n<չ��GP֩�w"O�L1�ܪt� �p���5(��5"O�Բ��B �����BG��0"O�4�D
6U��C���A/����"O���靸-�.5��jL�f�Ta0"O�"�n�{�\Aqρ�U��� "O�Y2�`�~�@ Un�7�b�"O�Z�#]�/�*�#cL�\����4"OlQ@�lĹ>� �J�b�=��Q�"O�j�'bp�����1fl�w"O���ϖ#<\}C�@T�CT�"O��TD�H�j��۬M4~)�"O�U��En��r/	�O�X 5"O���@
/6�$���O�<�xr"O���k�����޺pN��#�"O��#��!�4TP�-�$m�"OL��D�Ž}�I�s��S(�xP"O�A:�+R/�<t2A@�-��3G"O~x�p�J#Ap��ギD�fB+1"O,1�'W.l9��#2��.&Y
�Y�"O~��I���(����!SQ2�"O��i@@�3r��b�6l���"O��#g�,���pк2�\E��"O��)��ˊ�ʔ�T�Xg�,��"OV�h��ہzY�v�@����B"Oء��k�$S�zHH��1H�H�C@"O��x"J�2��b`��|��-��"O d�D 8)���y5�ض^��"O$DA�k�(Q�ƴ@�`Y�=�"O>�Bd�
� ��.�)�(�(P"O�qA��W��)�.S�5�܌�"O �qL��K�"��QD�[�P��"O�QM5>־��s�طCҀ �#"O���L�r#�LP�a�m�<�"O 㳫و.n�jR�'
����"Od5��W�uk���Sc�6E�2p��"O���e-:��0#"xޮ��"OJ����L*OV���W8h�V�*q"O�E����37*�y2�_n�N�x�"O"�y�ΐnf�-SF-ϲ���"OHX{��=b�����<;���;�"O�(����,s���IA�`�0HJa"O�����pG������Up2���"O>JS`[w4��r`��Ec�J�"O�m�G��~,��X�tUL���"O�-��'���j�lٴaG�d �"O��H�/Z� �b��׊V�
% �P�"O��p�e�)��a`�HE�e	B��c"Ov	�t�X(��Ҵ�
�+��x�"ODL���*@~ [W���Zߨ�9�"O�d��ֳ��a#�q:��b%"O
��qEޞy�ڡbc�R	 �9"B"O� ���>n3@أGi�����v"OT����Ϳb�h�Ċ�W�("""OԀ�C,N:!���Q�IF�{�&]2�"O"`@pM�}�v\�EIG-5����p"O��J�@D���b�gR(x��i@"O\���΄d&\�EB �t�%"O��鲆S�b�TlA��W�@��"O� p��q"�)��eJTȕ�^�����"O(�E�#u�ԍ*Ԭ@�3�@Z�"O�5ied���x�P��N�<�+�"O�c@@12��l��mU3H~��""Ouq�Κ�034@�%�ܚU��*R"O����+�&qXt���M�9�P$��"O����k�?�H�{fMN
l��	"O�� d�=���Jr��fj*��"Op�
ы-|�A ���c,�}Se"O�]���s�f�h����r!�"O��I&���J争:ai�?1O� ��"OF�Ya�Ӱ	��a`�ԇojHPY�"O��S,O�>'�x �K��W����a"O��B�BJ�kB�I�k�7I���"O�P�6e�9;�0y�	Y�-���"O�whU.�8ɖ�ҴC\V��"OdQ�ݑ�v��!�XN���s"O�)��6S���A
<��0Ҳ"O�x��d�0J��!&�j�����"OFT�f.�<����ғ<��Mx�"O�����,dP(d����:J`�a�"OFM�S�מr�t�&��;��Q"O��aRhɳo^����Z�_V(�$"O��hA�:]�Na�Ԁ$=@���"O�5j֚i8r���>m*���w"O�eӱ�3T�x�aV�"<�a2"O��CB+�ޡ(!jBqr���"O�D�u�ܮy�Ωx�K-2�Y`3"ONE��B^�?z����#n���P�"O��2boI	=���k$���:&"OԹ�dO:�| ��en��< �"O6$c���3��h �B� �,k&"OB�0��L\�wAI��Dx6"O�-������*0k���X�@4Z�"O�\�&�0\$@#_
c��H"O�l�Ã�;K�n�cDB�r��9�"O� H���f	yFc�4iv<B�"O\9Pbk��=HvP��'$\2�*g"O��kۛD;nph����Iĕ9"O��eܑb���J�,->}��"Ov� ̛�o��UҊ«]�\Hz�"OT-���m��:f�	/.�d��"Ob�v`�!+�Dy��:{0Ta1"O��q�C�n��3т�t��"OбsjS�g��l��K�g~�"�"O��I��]�+�T�����)tH A�%�'�!�J=����M�z
�����O s	!�Y�C�z�9��K>uv8SL�*8�!�$N�K�)1`䊔L��a�݄f�!�D�96��#�"��� �A%	��>�!�dJ�!�t0��ǘ??��(:��ηN�!�d3q>�ͳB�T?4�H�(K�b�!�dR�i�fpy�z�,d�GϮ�!����P#^1?���{���;l!�$8Md�	�B�W,{�)0�O�!��U8@����\mpAJ�j�!��&Ts̅�G�QE�,�&*G0#�!�� 0.��u�v�����ᶯ֛F!�d��=F.Xp,M���'�T�	l!�Ĝa2�X�r��<*|����ڟsY!�V��h���>Sy�Jr���QY!�d��R���HR���x�q���ƹ h!��sݰ� ��ڤd@�P�U�NR!�䎂iRJ8Qn"y�(�cS	I�W�!�� � �`D�}�$��늗?[���"Ob���*/iP�JGcM=	W�	ʑ"O,Д`��#>L�E��TB�E��"O�Q�3O'L<�]���)!�hrw"Oz�X��E�VU"㡜	S��X��"O�	�2�ʃ+�Z��� ��\i�"O��j�(��F�Y�gǯm�
���"O6�H��El8hm�EW�C��u��"OЈ@�i �i���� g�hЛ"O�頄�:�p%�E`�9"4@��"Oܼs��T7rM�u	���O��"O��)�m\��VՀfKZ3�,H;�"O�@��H-4��5�V��7)�mJ�"Ol�kVI�M� m*67	Z0"OD�I�j����`ƈ�82��$�"O�X�� �4pMj�H�<hc@"OX8Ke�T)!��hW�\b��r�"OP�P��U63�P�'%ӑGT�$�u"O��{��j`��ɲ���j��"Oxɡï@�������Ƣ:-��"O��K���J� =��K�$!h"O�y����9����#**{4P}�"O�[r�اe@���[�3B���f"O��!�:lJ�p��B��"O�hp���@��L�u�N�rǄ
�"O�Z	�&t�nE�����3"O���F.��=����B�,��"O|��aS?9V��a^"v( <J�"O�q�%-�k~�hȰ F�?a��"O�*2���񷯓3���"O��hd�}�DL����7 ���"OP�ɢ\)_���Q�"_?8�J=w"O2�S1� "��brJ��R�ZC"O@� �]�z(iT�Vs�t9"O��rddød�P�sCK����"OY�UIʣF`�M��b�;d�v�q"O:�Bs(��z�sB�ms�X��"O\�6��aҠ B�T0dÒtK�"O��R"&`H��3����<$�"O`Ū��!��Y�C�Y.�p(S!"O`�Q*�!V|�I�㞗	R��"O������KZa;'�:UY�4�T"O �#���3�Xm`c��bXfQyP"Od�Q�N�O���5G� qJJ�;�"O�Г��J�C,��@��e��[�"O��b��v���� C�{jAI"Ot�����xґ��OƗ}�f� �"O�͡�J�<J�!��U�~�aˑ"O����F��n` �EA�4����2"O��`�O�7l�����fh"(�"OΙ0��m��y�ʆ�@4b䑔"OL 0u� p���S)T��fY�"O0��Mb`� #֧����{�"OJ�����aO�ī ���D��v"O�8jf�6H�Х�J�y~��
�"O�|y��ض3X���.�"^r���"O�8�S�U6j��`"�<_V&�K�"Oc�˞uq��x��S�g;$5��"Oj�k&�!9�d��Cʖ>5�$s�"O��!Gʏ4�reZ��D�4�a�@"O��&�3S�LZP��(.�Rm�v"OPۇ
���
,J'+��Z��) �"O�4q��O�V��:������3"O�(��Ɨ�P��9P�ƍ�.8�0��"O� nԉP�R�HW��ՏGv��"Ol�c�٣D��ӡL8p���"O�#�dկ,��+,����	�"O
H�j��8<d�JB�)p�b5"O�!����-|^�h�DM�g�q��"Oh��+'N�X�Ӳ��L�5"Op)���Dkh5��CN#s�����"O��6�٧&��ɦB��0�.A p"O�Q��kѨ�����~0\��"O�(ز��T��h�]`@)�"O�ID��D�
��%IҬq]h C�"O ���)V9XE��zNF��"O�ș����V2�*�͉�v��"O�L��D��)�41�,�s�"O���ƒ�Y����Ǽ[�F��"O����h�>�^!{Qʭs���`A"O�s�+� Db���a���g�\{s"O�E�.5i�9R�N7}�"Op�P��	��y#f>Y�<5�s"Oԥ�4��&,}hQ
�/�*���"O�=�0�\�I���"iQ*mF.��E"O=����2�6�5J�0]��"O"� D�k�Z��aɖ�/��U��"O���J�UF��bS�ЬO��5"O���"μ2�sV�'y�:�ڇ"O�tA�k�F���լ��+���$"O&���jӷx����I����T"O�"G�ߩg���Z���چ"O�AB���p�+fS�FV9b�I�<)&k� 6��4fF�9z����Z[�<�aL� ��H��c4-5���A,�M�<a��&\�N%�0&c{ZL`P��M�<I�A
�[�4T"B)@�o�ؘ�G�<1����;���r�ញSÒI	"��y�<��'V��P�ȅ�Ԉ$n~%����u�<	�㊅NǢUB�J�Y�V��6̞}�<���SDR1Ѡ��Y�"���#�q�<��R���F�C,e�t��!�j�<Y4�&F~��v$��l*Y��)�b�<�B���|���i�k��]K�K"D��2�@ҥm�XU0� G#~r�!�u  D�8q���/��=I�j�B2�1��:D����߄.y��g+04�	)� ;D��:���A����jЫX}~�2��#D�����8H���7FOmh�Ӄ�!D�h�!b�+r�5#r�N(�e#0�=D���bE_�f�RT�)�0O���g:D��xbb��RY.Ȫ'�6,@�c�i<D�@�$�-
6����jN�'�As��-D�H��H3#����7��.Z����P>D��cR��'����� `���Q��0D��CR�X0�j�p���7�y��h-D�<I�`ݺ<XM:D.U�aR���Bb/D��g�O�P�P2�'p͌�r��+D�����.��)35�C7:(��#�)D�đ�/S�<�>�C3� Nd|� 	=D�ܻ���x�:�b'��^���%g0D�0�%l]&3�L����c`r�)e�!D�Ppt�!/��� �,@��݉��>D��A�E�G�e��$�<h���qQ.>D���V�
��!�d
�;c��͓@,1D��Rm	��\�����)�L9D�����J|�2VËL�XH9R$5D��k"���p�0�HHL'D�� � �d�S��4����of�ɠ"OFh��O7-��E)A �Vyx��"O� S&�9j9,�R�N8}j��"O�	���2/-�8Bc ؁4k���"O���R�W�`�:����+��1W"O4��.14ݤ<����+����`"OL����Jw�(��Xwm�x�T"Oν���+��pZ#!ҙhV��2""O�(I�)ћ{Ͷ�Qf��|�H��"O�m�!`� �؈c@�:�꽛D"O���Ò�A��q׎H2g�%+E"O�q��C��XYޙ�C�yw�%��"O�q�EN1'��3�W�aT��e"O��I�eڪ�h|yv�F����"O4,����"⨋�eY45��ب7"O�t�t�ߩG���v��?��cD"OpL��Ǔ/7�*�����@"O�8�T���X�ԁ��1.���"O��r�D�C�L�:�cZ�f�\1�A"O���ê%8��XcrA2�lEHt"O6��'�کS����Oݫ2:M�F"O2�@�J��^��m	�.��|K�"O
HP�N�R�����ѡv��,"O�+�JK�#�TM&" 'w,^��"OP� (����	���8s�j��"OT�J㈤\��1�0e�0��q�"O�4�PfG������C�{�Y�6"O�h��&lq��.ۭmrr��"OZ豖��F���y��E�Ra�q�"O�A2Gg���!� �hC�Q�"O d"K�[p2�Za��%�Ty�"O��K��ۜ`�@�U��	T�R"O����n P)�t2Sk��VZ0��3"OJ�;�nnaJCq	[�Q����"O�5�BN�5�D�˰���b�x�(�"O�u��Jm�����O�i��d!�"O�C�kH*'X�<Rb�� �µ��"O$US�0B� I�r�<���q�"O�)	���{���3���v�axC"OL5#�&\Z̱��=b��Q�"O:\c1�Zw�dx�,�����C"O�:�(Ϣ�(Y���`;0"O���1�T�Ai��q�KN�bQZ]9q"Oh�k �MbR�@�&�׊Jf��"O@�/K�
!;EF�"FE.��D"On�j��%I��p��./���"O�r�EG�X]�؈)*��ab"O�l{A��Z��t�6�
2�)�"Or|�bgC�Ɗ��EH^��m�"OLi��Ĥ����!��?rશ"O�m���N>E咅����l�Y�"Ot<��ʙ�9���*���KYN���"O� H���I��iT��79v8""O���f�j�|����c��"O�Hr���WŪͩ�֌'O�D��"O���RF9C=kG I2L;bL��"O�a0Ӏg�$`�t�(��)CD"Oj0��ᎈ4��q�2A�J��H�"O�Ų��B�UX2a�?s�d��"O�#&���;SR�"�bC:O� H 2"O���Ð�\�k��P.F����"O^-�턍��� t ����I�0"O|D�@P�?��k�%) �C"O���0)��q�\8`d�8=�(c$"O� \(i�UX����"ɪ �>���"O��R!��t��(!�	�h��}3"O~4A@��:�~�pQ��?�Z}��"O�#w�ϡ#Q�P�GJK�/O��i�"O.�Z�NF�k{�u��I��x1��"O��*�BNh(f!��I�d��:#"O�Tk��� ~���*A�T�`x&�rc"O�qR͘xR=�G�!di��sG"O� 	����`�dAqY��"O�l��"ӝa�2A�@�O� Y�u�"O@a���W b2�鄨C�ͳ�"O�� Q�/n���@HS�'(6I#6"Odus#⃫����f�&}� �U"O�9��Z�2�4S�[�M[B�b"O$�CC�ݬpT�4Y�N'-g\(`3"O&e�U���y�6��g�̴`b<9�"O��)��LV@��s�.^�|���"O$و�n�)js�����<���G"O��!��a�.�����	���8T"OH� S'���1�%��
� ��2"O��#%�d��%Sb�Ġ#Bx�"O쵳+H� z�	B��9z
����X��2&/K�	St��mǱ5��B��$D�L�Af0jdEʬ�8	IGC�훦��f�'0��3�
GJX��{�E�<t�i��,LO,���a�	3;�Ȍ��QZG��:cC4A�B�F�~���7o���r���Ig�OZ�	Ӹ����Ol��x2tњV��x�P�t`\�[!�ֿODp�'
�B*
d��5�0�>)���	/<�H���ۃI}�8$�ۘ%��$�-xi� �ق]z���m�>�<B�ɞ;e�0�UY0S��TH%�ө� B�I�J�K6-[-^�h9v�Q9B�{Z�<�qG;��zD��i�
B䉌��9y�n��[��OY+d/�C�	�Ki�A#c)T����I5�#V/У<y���񳣅�������&qSX��t�Z��5'ʃA���3�M�mFp���X�h��	4P.:�+`��R��t���)/�J�Z�	?�h���v �[��T3I�ij���<�Ȅ��	�<���m�B�-q4M�r�+/��B�	�P��@����[��T�ec�ԥO�eDzZw0��A�Z=J��8AvC�O����'����K�C�P�sPd�IPi�,O��=E��`���0 J�=�A%�՝�yb+ϕ)��P[+Q d�8�㎷�yr�W�(k�0+�替|ܜͺ�FL����hOq�^�Y�J$&M>�K���7g�xUh�"O�@)�8����«��k�ƌY#"OFA"r��8\�Jѹ��U�B�"Aju"O\�BOʷO�m�� ���a"O��ƍF���� �H	k�F�I�"O����ӸT0����K|��X!@"O�	��#��Dp"���1dYP"O��SHP�,��*��A�0q(Q""O~�(Dd��4ND� �v܀s���y��<�\$�W�	�c��QÏY��y�d����H���>�@�pc	��y��={n� C��3��8��KŠ�y2B�6"f��Ԯ@*1�~8jF��yr-)ֶ��$�"^��� ��yb��u�u��+E���&��y�aO�[d��4D+k�����/���y
� ��Q�3Pz�a`��x#�4�"O�-�U�ˈs�$H��N#��X�e"O��f��e�j�ZDk�$*��e��"O��d @V�� ������V"O��	�F;�u�@G�z�:H�"O�����?~*�S2M�2O�I�"ON0���V�C�M9�KT�TD��'o)�S��yb	��`�܁�6N��&	��bag��p=��}R�ӧ$��z@ܰu�1`J\��y���~!�J̀C
p!P�5�ybJőF�x|��C0���
Х�8�y��NJX!�U�|�1�"'I��y��\�18UK��+�<�2� ��y��_�/��0���L>q����ď��y��!E0XI�$M�hC��ɧ����yr��">&��"�"_kd���F��yR�Y%@<�Q5f��^H��b'E �y�J��ԅC��Z>�)Z$(��y爨61L�1�iT�M�vd+dE��y��R6u8�`��?C�$p3�dƴ�yktb!�5��}h1�a/�y�+&/U�[��9��(S�`H��y �
��q��G�&6�2� �^��yR���N�K$h49��8�o�y�%��*��1%��b��;�y�jD�Q��`�c��+~��FE��y2̛���ƙ*�bQfȒ��y��W#@�L��V)�%�Q�!ܙ�y2$Y�EԄ�Ei
5A�B�M��yR瓁?���e��C�~�c����y��OO�ȊCC[�pNQ� ^
�y���R$B%�Ĥ6����b��y�@�2mUL�3A&K7}(`���y��Z�l��2���t��H����?��'���@��ВC����q�I,;���j
�'TЈ�,]4��y!dH6{څ�	�'��Z�L0:D�J����1%����)��<q��k  ��w��9)0P	BGD	D�<QV�S� *�嫕��1*X�̑w��~�<�3��@���)�A�-@��Ԙb� t쓘p=�6�/#h ��%=.����Do�<yf ��bjDı�DP�|��!�k�<!�G��H��U_�	'l]��fO�<!@'��t ���+Y� �
�ӁNJ�<yթ�Y�b ZDkG������C�<�s>�������|�@�f�<��@�U+�H��D*��P�Kb�'h��B�OH
����X+=I6�Qp�ϊS�M2	�'�h�c#͊!di����b��\X�	��H��	�(DhFA�O��8Rl�,[4B�	�_@�V%v���D�	p䈐�#�a�fB�I�v�xi� gJ/-MP����%A���D;��5m�(Ёg��Yh^D���A� �C���)����X� P��ԙ�y��'���x7j��"��'E£�y���Tܴ��@�
9��Z����y"nޗ,��y`�&�v���ǩ�yB,�<v��4	B�ҾW��x��-�$�y��!-#"�PC/O�W�^h�孟�y�(��i�F��e,.%p�d�`DN��y��ۡVY$��6�ŷ%����X3�y�)K�d8�����T-#���d"�y�/�.{�4k����\�g��y�)^��
��J�����W+�y
� �	��KT�W�,��g&�J@��"O���U�Y5�ċQ�C�'�Ȓ"OD������LI����r�m�"O�(Yp�X�@��r�̄M�йC"O���	�]�n�	4�#5>�[!"O�iR#L��n~<��v,��ufz��"O���a�ͫG�$0x+J<@>���"OF;�n�6rK\ ru)�<t&�E !"Ox���ӑP���Ӧ�!$ƥB�"O�4�ЎTEjveQT�̀x�+P"O: ��fΤ]؆�ܡ
���ç"O�fh/F�`;v,�J��a
P"O�l� F��viH�S3�գ"��ݱ#"OE��)ݿZ����b���\�z]�"O�]R�� DP͐�� gw�p!R"Od$�+�({,�9iB�'fW�U�'"O*D�l�z��i��X3I�- �"O�p��j��9�f��S�L�&����"O�B�mX�t��SG�+U�H�"O��c���&K����,;���"O�A�`�ڢ=��ʇ�5�n���"O�I`��o0qp#�)m��(��"O�!��S	��m1l^��ȹQ�"O"�# �4E��i�Vk��4��"O�ipևkQ��`�JM=Jwbu+w"O�	(ejˑ]�����ǹ bF�p�"O4��ؔ,2XТ��%Xi�"O*��lJ�z�ʴj���,G���4"O���k�8WL@i�D͐#7�l*!"OJ�@�h�/;���t#�e4Ȱ�"O�I��$\�,��z�a=��]�v"O��3�@�h=��*�C�,D|��"O޸REbZ�[�4ق5�8H�p�!�"O�A�D��3�2�K��Y�uEt�BA"O00�'�˱nX܈"�=i_v@c�"O�52� �V�� z��>m�<���"O��R�ΉT���i�8�-x�"O@�	�	��d��W��Z*p��!"O |9�GL_i��)��B���3 "O�]��nř�#]�g�F�F/�O�<�AG�-'���B#_*`�@��ETK�<�����_渥�a�#(s�0hq�<� ��J����	@'c�$�I(p�<i�Å5[�p��f�%q]rP�g�Al�<�ٞa�����k�	�>8:&��}�<	�JR&*��!$IT�i7�Hy�<�l�_*<�Fϛ|�.8�Q�Jw�<Y���*Xo �K�$߽mt^�z�Άq�<�b
ԍ�:|�"B;4���A��Φ.�^�aH4+M>�;�(�\��0a��A�rO|����{�� y��=D��:��9d�����ި :n��&�!D�(�"�Yg��mJ��T�x��!*D�l���*7
5³�δ�p�1�#-D�6��=|[h�)�-W8�X�X5�|�<��U#Xf`9�Ӛ �⠨V+�p�<����d-^	3"睔yJuЀ-As�<�C��� ڵ�4���`Mn�<����#�T [;`�P�kCp�<a�I�'8q҄��L��L}k���p�<q�J�,]��Ԣ��@?V':��Ţs�<���E1�$� ��;'�zk�Of�<�soп"
D�qD\�
\�Z���g�<Qe��
�¬�V��*��Z�<��Mt0�c�6ib:�i��|�<� ���V���X#�q��2�"Od�1!�O�tQZ%O�>-�0!�"O��	3�P'N6��щ�5f�d�k "O�5�0.�H����i��N��A"O�%������N	9�(�m"(�qL�(y�������(��JW���@hi��@�����yRaY:*u�L���؆k��C��?�BI�m�a��N�;��hÓ;B펎P�N�a��w�xЅ�	>.�����8%~( CQ�1��p��
<�xy�CQ�3-
��'2��97d?{�>�x&GG�6�b�'�� �KH>65е�����M��'1t!��h�,S�Z���B�OZ(�،�D&�S��͘8�@\�6+XN��+�����x�ւ
~����+X,d��[uÐ�~�v�/�S��M%ː�'2,�2�MO67/>a�U`RNX�\���ۛ�(E����H����O�1t�I~��}�Ӫ��D��ЪW��ȋ�D�'��U����S�iO�	hh|�f�>{�Feq���$|�B�IHSHp;�F�:!�������K�������i��܉��T?��u�H=� 8U��IYP%hAi*����g����`�H��T�g�R�A����ڼ�O?7��;�U	�A�5ʺ��)�*v<�xB�/*�0�@+E�Nv�b��B&wp��X*vp����I�X (O�4;T �L�#/�>�����F\��>��)�'i�:b�̱A���.{�^B䉭<K܉y���% �52Z{�"=����^�O(^tc#�*��N�
i�^��
�'��2�ςCy�p�Xdn9A�4_U��Ex���i��l��
p~�:S�O?]� YK
�'�\|�W3�r�ХK�P]�DˮOz���'�Q��cX�5o��begǱO��@{�a��]�'�LŁ&�O�g������O+�իߓJ��,���>��#էo5��M�#S>N�qfM�'n`l���}Z��%N"@�	Z�e�"�qO��%Q�X���ۊ�陆}Ԇ�iT��63ryEÕQ�����O?7M�]�t��I
�j*�$�AD6��u�A&>��ʓ�v�F��O
kE`öBS�9��G�L� X��^��r�1�O
��!�js�p�w���6�c���>:(X�F��tǋL�'�0�k�O�`@�[��E��Hޔ���	p�'��U��Hߖ{���90͉ƦE�'�ʕ	 nD��E�g�����=ғ��G��`&e��B����(�L��آ�ēKS���)��@�����_��(�b0 ¸
�HH`��X�<�j�!�i'�EDy���i��;F��i�!�E�@NB���c���j��=�	�(�!��L<�!RzM4 ���al��E\t}��AY8�L�o�Dz@}�O��)��Di��R�w��i���V�`�ҏ�T�'Q�*�H�B�%P�R`� �  ]�1�則K�������G��[)�r1ڣ)���N �a� �.���Í�d?�S�dg���@�c���i�|)�F�
���8�����Y�(8�D�Ģ��(�<��-�.�$0�"A�m�p"O�-�2oT$JN�A�%�9��I�E� +�Ra℄�$�?)�K%Z���'y^�:B�˸~<�C%AMH����'���@�c�/h�ˡ�� ��x�G�V=� P�׹� q���v�1O2��hT��`���Ip�M�#�'V��P���Mx�Q�c@S�QCR���N�t;�@�2r������Su}�[�y���G��v��O�$3O<�hP%%���.�"f��C0 �`�I�#e��s@�!B�YB�?!���@�C����zR��+� �/5�!����l�Q��;�OZ�B�-�����}�r�����$���n�<��'uH��'�96Ǫ����`۞w���ad�$g5�AS�M�%q�8�*�'Y:�4��!
��O�<�"��Cw@�@!Q������� _Y8����ȟ�D�2;�n�`t����0�ΎN��{�Lq���'��k�B�8������t��ԍ �gc�����|&x� kV��b&�/"}	4�&n ����	_s����Z�x��i��Q�$4���C�ʢ�̷�����3T���aa$hx�����"@�h�ʥ��ph@�T�8��*��5�e��C�D�*E�ؓ4���*�� Ұ؇J;m�P�gc4T�]#�"O�1�Tw(%U���%x��!���bV�	wa�Vz02g�0��|�1�Fp��L '! Q)�I�$#n܀"6"O�Ab���,��9HW��ZA��.��&�F���kY r����䎚��Y",/��0�����0.�@|���r#��k����D����f���OޘM�Bӏ$~\:����f��hv�V�E�*�����@]s� Z�d�fyA��'��#O2K�<�8G�[{i$�M>)w-۔xa  ��aJ�}>�˔.�vݴM�צ�Z��'�<*��(��ᜓpĔYBnE}�ٻb�'<�mk'H̏����]v�l�bc4s�����ρ�h��] 놡-:�qSW���ц�݆w�`�w;�L�� �
�U��b��K
�'���%�z�܁*�k�6wK��iÏY�|���o�`�zuCǄ�2�\x�U�F��ƵBv��pD��s寧��0�݁}~F5��9[�4��%O��1�,��1�v�#"�Z��<�G����q&�߬)r29xRm����r���%e���GR"ޢ����h�'�n�1r/��q���QIC�A�Б�O�uC��N�[A.=I�y9�n�U<0]h�hT���³��&Y�����D1�\��¥<��D�E�I�p?�[�
��d�F�M���Ƨ�,}N��A�JQ�JYt��Da̿jwH��d�F��	*H���g�yE��]�n�2-i�'��`V��v	��C�ɷ�YH���k�$��ce̘
qX1T.�+:��9O���ԡF�}a"�-l�:쩓�~Fz�'��!���"S��%��+\�=k��s�n�@Y�'��,w��і/�&sG�Zֈ�6[B��JH�7���W ^#`�&U�@�|��h �L�z�-"&�I�]kF�[7�%JB4#�HV"7���'(��P�H�/Ca@���8��T��a��"T�\�<��29��<R�F\�B@�1 4��J*�O�48e"ӗ;����n���Ǌ� T),A�#۬+g6���|��`�2O�݊�Ə�m�攳:���h��n�@t�4���/T�Q
OJ$y�D�Gb�*��X�Q�Z"M�RDxpQ�֯�yr�Ѡ!�B�S�d�H|�RS�V�)"ҭ�|?��À_ �@T_�W2���HJo8�� 3��y�@����_�.��� �>mq(�Sv�H�mO`�Y��&*�TȻ�g��b����&��tD�Ҋ���O.�BB�̔�8��#C9��q��>a2	�(yr���YG6��b��!�bX��g�:%�牜:&i�7+̳1" (�K��5u���c�~��~R��'T�8�[ׇ�,<d9WA՘��E:5l8sqEQP"v\���\��MGn����%��Qh`杶*m�� Ã��kʤe��*Dl�v��DG�(k��A�:z��y"X�:�4 `d#EB���l|�F��4
� �'ц��s�f���� �N?i��Y�J4p�����;B �*�R�'�,���W�=  K�G �;��� d��q�7��#Sv�4b�*ǉ$�,(f�߄yLPj�ǈ�Q�h��1�ʃ�O� 8a���\ĩSf�,a�.t��S��RqGH���� m<P�Q��|���ԫ�(���̓	l �0�E�(�z���N	#`6X�@��	�\����V�H��([��9���r��m�-F��g��'^X'�Xuϋ�1B�� c�Yc� �Hy����/G�|YȈQ:�O�IS� O�c'&(���0�.$�	�Yt�5+N<Y������b}��i���>��k����+R+*��1�ʪ*�tˢi!��I�L�@�gѷ-��`#�J%���tLP��J�s���/"�`m�h�|�q0�O�0���ZB��x� %����G�'�:p�F�T����2��H=e���)Ot���Ŭ$����fG>	���H偁�,�R�Zڴڛ�b�Ќ2ZZ~0��/\;	����XeP=Yrk��*�ƽ�@�'���rf�^'�r�A���6Gu¼�wϬa��I�@����HCgL��6M]��Y�!�#7��AC^"�5ft��t2o������Ӡ���?1'M�p�L�����U��-�f�$E�9Y���);O&E`5/}�H�$��#��b��&��#�-�N�$�B��*U}��� ��2�����~������I�VzX��C�/���Gҡ|��	���J�.���<CH��Fߙ��	�ď�N��M��dU�k恱�m]L�6<�T�\T̓K�L$���ӚC�Z�JԘL:V��'iyR��
�Vl,�05gӮ��ͩ��$SM��J�&RVw8�Ja�C�I�i���ǍL�Hٵ�J��&��n�oSn��$hD�_h���䂣
�d�F�@�R��E���ݨyZ0� ��hqUi�?Iޙ��"	�r%��'�O�q೤�z]>$���
-�2H���
y਻�㜷 ը���ڕX'8��C�К`
���R���:�4phs�Z(=8�A&��)*g�4���3#P�d��ʂ&�<�"T ��*9?�W��+F�6���;>�h�9�*���oS�,��������|�!�� ?ĒE�ȅ=C� �z�H�P�D9�S'�B�KԩA,�j�yE�U�=a�H>it�#b�9�'`٥^X0p�w~B/��H��H���ʫi��I4�M�a��kJ�m���fH{�&q��#ic�}:TNT�Q)�!cō�z<h�Ʀ$E�V�(�B�rX� ���R>h��̒ ��>��8jز	�2��&��=�1��O�U���Ь�<����ܦ�xE*X2�$u��E��H�`bAؿ��uzRd@Z��%;@|��K��"(AB���X���k$gX�c����'Nf7�\";��-�'���>0|���=�p�R �3o$�Ai\�8��4(��'m"�11i<��pA�@(��*��~������Sʰ1��[�-ؒ�T3X�� 2��X�`]�AS��*�Z�=�6�m~�)ħgV�s@`Ρ|o*(z���'m,8Jf`[�p�RT���� �'�� d�9����0_�j]!q�0r��P���o�1��N�X5K�j��,Y��S�? �]ɢj�L��$���E����YBKZ�/�ZQ�Hm�Hp��j�� ��M��:O��FM7���9��)������Q/Ek��M�$5���`�X�x�!���_���#I��d��A�A72�V��%k�<��F�r�i�(�Y��=��)�5a��y!X�5�k�W-�h�B�J)u%�����)��1|O�,�'�A����6C�)����;����HA&X����@�R�
��C�)�DZE	���Cu
�
9����q�!?�Ї�*v80��JҎ�h a�J�'�|r���'E�F}�1�\�&��	&Vqh%:�®V�̜s���O�}.U�y�!��Vmؕ���%	�8���	 ��}�����*+TEG Q����~אL��a�#/1��� ɀ�M��/��&�e�U�I@(ܺ���{�hK�1��B����%�]�Jl!�$HR��`T	솁��K�M�dE�@��?��iWr�c�+��Rn�)4�#3�� ?��}�H��ѻ"9�а7`�%-I����7��AUS �Ж���:w�\J)�X% �o�:Q�Q!s�͹�⁊VT�ȶ؟�[R�tR�Mv���ґ�#3�����,6qҭ�"�#~����T��T��_�`�:��[�gYH�ΓL~��%��QM�yj�{�`9�*�)(tN�
�/�P/�%��8%*_3:�X�3�����Q-���/֣M��� s,Hn5��Ąiv���ȓk���"��R�#�j9:�� ��k?�I���O�(&7��V�K:N��"Oұ+��M(.��I:��ӰBTv��r"On)�p�Z������X�/�=b�"O<��v� 2[�4�c��+t!���"O,u�@�W�(��x��*&��$"O��+�Ξq'�E�&ېB����"O�͹p�� �4��D���t���"O����i�P�~�ґ�ԇI��|�"OB����X^=��#�M��2��"O�HJB�>]���Nèjo����"O��sE/T ~�`-Q�HHW���"O"�qQ,��%�V� ���YA �x1"O��EҀW�V��S�	'T1��`�"O��a#�����l+!���A"O#Q��\i8�"p�ʗBz5+�"OZ�P��RUَp`C�2��"O�ԸS���$)3!�Hd)#"O�,��nP�y�TF�(�МhU"O��J��G\�)�d��?�D�x�"O,XCck	4_��]�G催7f�DR"O�d��E� XObyrEE�=EЁ:3"O@��0	�OuD-���Y�f�� "O4s��%��`z�F��xށ�'"O���"�O��B� n�Ne��"O�d���F7�4@C n�C�D�2"O� �@&�2�r�� �Y��-P�"O��BOI�Z:�d ��̋M�
!"O�� E��*��YǬ��Q#n!�b"Od�`��v|~	�f�V-6)��"O8�)��8FC@䈤�$%�p��"O>Ɋae� >��!ʚ=!���"Ov��šJ�]������Ż��yE"OP(CF_Ht����J�*^���r"O
XA�#� oں��!J�jL�x"O�ᢩ	����o܆1?��ʁ"O���E�^	�Ջ����z�A"O�� (�(��婀��
$��q;�"O� 
P���r	���M	�@YRt"O�M3E[�+k\)�oD (�Q7"O�pR�dU�=�fh9T�$qc*���"OԑI&�_*���7�%Kd��"O,Q{��I�j��(a‮}p��"OvUɰA'�4A�G�ߔ��\�"O�!h$
�8l�^a��O��4Kʤ��"O8,Y"�fxS�OΕK�x4"Od�H1��m~�!����~:4�Qf"O�	T7� �CЪN��,4["O� ��9����Io���4H�qD���"OV�X6�ؑj̘T�c�@c"Ov�!��ŝpG��cc�)	[���1"O��@*ޏofr|X�]�]��4�"O����G�6d��B,Y��̘�"O���hׅ<��@J�?)�&(I1"O��9��Bb�8�@�ʅh����"O�\rC�^;$l-��ׂ�d���"O
\��J��x�!�
Td9�"Of�"$ �9�0��� 4$Ѐ"O�l���S<s���@�&�5+�ؓ"O������e a�Q}���3"O�q�R��:Z9.P��Ϊ-0����"O$�����K�(B3�i2�"OΤ�B��J>V�@�HK1W� �"O`��D�C�Pq"C�ђW�`$K�"Oȩ����T��	�y�.<�d"O������z��"��Y�$��|�"O�XhŤ�>s���⅕��*�xG"O��嫜�,���Ғ�������"O�yZ�b�@�e�!b JqvE�"ObYS�`���h��h
�s�XD2"O�<��H	!)��Ѐ�̞]��A��"O����s��@֥X�M$80"O^�D�0T:\Ѷ��F�nՁ�"O~�S�%U�>��Z$��%=����A"O3���
n���	D�������"O����(�������.Y���"O�m@&Iޮka�dc���7���"OR 
�)U�c�������T"O$��/�\,3D�ڞi��"Ol�Q�C�H�e��Pa+�X;�"O�PQ�k��偲�J"6���"O.��V!�q���ڑGa�"�rg"O a�!ET�h�1��ác�E9�"O��A���f/���A�J,>P�1"O���PE�VX��JG�
0�ܗ�y�/�)
`���փ�"pD��ք�yb���\�T ���%�@N���y",/_��FA#u��3F�y�b��=�����M e'z��e��y��#P�r�h|c6�{tF�Z"!�d�"]]��Y����]�����;!�$	�$~҈�����hr�ʓ�,!���P�7�K���yC�I)z!�d*C��򁏞���\���ʅ�!�䅦�Ɗֆx��I���~�!�Fa�����¼f��$j�o�-5�!��A�P��� �Q�61K��<�!�DL4�8IR�5�s�jV��!��#��b�%�1IVXz�#Zu!�DC=g�pMh�!]6O܎��Z��/D�xX �B�n����%��L�� ,D���A20�R�j��(�҄ 0�-D�X�r�܋�	z2/O;Q���0�M+D��9�eʈb�:d1��U��I"%@-D��KU�[G�R��#��=.�����)D��y���$��n&)���UY}��߼t�4�X�V��Ȣ?�h��@s�@�Э�x񥧚lX��2��O4[��1`���z��yWk\�T6d���$J��P��;�O@��	����+��~E
�YS�I4�J����M	|��)ԫJ���* ����,Ǡ9�Vc�.�]��C�ɪo*X�Bʇ-MSc��yJ����B��-�r4���67໗D:��<�nW�D��@p	�&}Ɛ��U	^q�<� ����FQ,.�D��hD!T&С�Ɥho��B	�H�T0
�"\����&1ړyf"�U`Z�b}�D���I��謆�	�Hi�t�a�(|m4< %&�1'Dp����Ԭ��b�Wi�032$�7��>��@Ňd�T�0� ��FI���z�h�����		��	�2��-*䕲�Q>�b��:J[ SZ�VK$IvB䉴N$����	�n��$���Y�$aC:���`�vE$�1��t�O����7y�xX�aI
 �|����eC�ɫ�8�jͺ ڵh�h������@���s �q���bѭΫ��J8pĉg�>�cmV?�h@���rB���Te�V����L��"�@a�§ʞl���bv.����s�/=]�$�&!��a��� �ν�����ҙ`�����&�9��UP��B��%��'R���2�͝!��"(PD��0���)���y�M��%��=a2"�	�����C�*$���4*�$ f��D]9A0Ad�\�*(���!�u���;�dR�F����r˒~x$Y��ݸF>])��),�����v��5B[RHR��6J�T�C��K�\{���ڡ/�$pb���w+�jd�R�{м(�C�vSv�Y��I�E�&e�� L��*P*G��q&�0�m�'|Ɛ��+�P���mM�h�� S/�o�(=���64��}��b>_�������cR��6?r�1۔@C&+u�F�<#~�A��'�H"H8"Е:n�;���� �"����"�>�`���lv�@�aBq�V�d���(󀛇(���Ĝ$�b�j&MO�3�)`��L�#UN b�d��w䏁sH@���'�H�#A�N /X�+�GR P�1j���8�r�95u>)Z0��0�\�K�'U �Ç�!B�Y�wȽ:Yڄ]0��ؕA��u�6�U(<1�*D`�H̯hՄ���GVfD��?c���	�]th����z�k��,oښāe���i��Y�*D
ף� 3:�2D	
�x2��	���+Ѧs;6$���5^$P2����q�x�f�7$|�ɫ��æT�6�S���0g�@+rg_�Y:�>)ׄ4�lI��i��A���!S�c���7x��)�F�=@�l�pFS�n�"Q��(�3i���'門
Q��'P��($!�:{؈�BCH*��u��Ii\@#�*��ygm�5"��Z��(�g&ķ��U㇆�Z(�x���	�zbF��5|nu�U�K^����R]��I+t��$2�${lB�	E��`���M��A{Ɔ�&i�:�Ō�)�
!�t:OLx���R	F^�D��	�0J��}6fE��#)�c?�S��`���ӊ˭1� ��g+�P8�p����+��L{��^.+L��o�H�N蹁B�0�n��m��QH�L�EW:xPSלX��dP��ʅϨO��+��վ+�v@���Rު	A#�>�F/ݧ"��ikr���~J����E�n��]�*�$c^�!\ic0���W5���X�$y4���"7!�~�/
8F�IBs��*�*h�@���8�l����ܧ2��e�rIä�B�cOv�oZ�3��&�n8Q��"߼sЅ�+QX�)��<�����a�n���j�EL�Y��	ƥ�!�`�D��Q��U��%IaX�m�m����.k�.@!���5I~��Smғ�P��'GP��J��H�*#�w�>Xi����_R�z�
�;�邐E��Qcdt�L�0g������O	ZHau�E�1��[*dV�Ճd@ėSn>Yzd�	�
C���@��"�;���]�6�B)-Hl�SLݜ�(+A�V+�^����D=���	�n�ڡy����1��٠�Q�Κ7unVl��I�p�K`,��B�|�C�ǁ�M�q�o�3�<5QDkF�Pq��L<y�H�v��hg�Aü+cM�`��΂<>�d`�BG�B��$�G�J��RF�r��5ғ�O��򕋄�x��_�.P�S��1L��p�n�?Au��т��}?w�P��@Pu�_1H��P�\S�'OT��!�y~� XEo��uBޡB$��>�!�e�)9zv�%L�n�>��3��!_h��S��8W�Δ��-���Oԙ�`��%�	 �lQ�g/J�5V�$F��1@@��@�D�r�:��)�d #$�i*�6���i��쌥
��9B��V(f����M��@��#U(h���ə,���Z���.-X�b˓�VN��2��-#���""Գ*�0x@���M�e�i2��He�K�ItYAfk��k�����8{�@Vpx��'.�O��[ӂI�0S�E���>���B*NZ�E�5vѠٴ7�T�
Ui�8j���� �9AciD�S��$�ÆK<f6��3��b1
 ��*+/��G�N9q��Q4���L���7/؎x�Ȩ�q�?#- �0�-���%�܀�Ѯ�&!�`%MV
�|�.͙��Sb"�W�1O~�y��78��T.ߡe��cR���2d;y����C.�Y`���̌(N>�����>�֠�eH�Gf�"bc�6�x�/�$@���TA�.%+�y�N�$�:D
ϓft="�oD�9o�� ��#W�,�v��D�PX�C&��$G8bUJ�ezz���?QRd #W� �(�����"��M�p�@�4��gݠE 	�'*�eρ�T"2�1��J�cay�f�W����PN��
�'m�PA�W$"�iud-nQ!bF��S�
�"E��oXڡP��K�zh��E���O�mI碕�B4a�Q��r- u��'L.��U�\��B�>7��H�d�I�@%��͎�
'J�C��"G8��n�_��0&�$���9r b�0G-��� �c'.?�QڡB'&=�'�c҂�K���1rD� s���i�N}a�f�s^�`��V���Ђ	��Pc<qI��C؎�HE9,O���eK�yZB(�mIu�~(��^(X�.M�w�E�-ވ�0��V2����+�D}b�f�l5 ���*]�����7g�2�����7��a�b0��?��fB%:GIz�e�>P�����ϟ�:4`҃d�1^4�~�����"� ��b��B��`�/��	&�y
� N��Χx��I����H�qR7�'���yƅ�"L�U
�IŨ<
X�OL=��� 惝;��I�� 妁�gc���b�S�Gñ5�!�� �;Pu�a,�}6�S<�& ��jx�H7��%����<Y�+&�Ή	�A !i	��V�rH��jҋ��<y�G�(M�pzp�ҁvH�1%��3rv�����$ (0) G$A�P��4��g2T�ICjH�b��)���&�|@F�E7���`fi_0>~�]z � e1\手d����'Z��T�cD?o�e���)�1�DVW������1����	&��0���-OZ-�E�X���t�q��O�1�բ^��-� I���<�h�HH��y�}j��هdZ�U⤛�L��|
%���=��M�QQ���`��d�T�Fm���[�F
=a�oL�M��]1dF@�E���C$�����X��l��Ek��J�>���ǆwL&�2�gU<2w����չ'������Z���Fρ4>Z���'��dL�9Q�ī��hBEǘ�K���S��K�E�l<�1�L�Vw���d��&�����G���0�T��$�L5�\x�O�����
�̦���iFA�ɑ�#ҞP�D��!�5���KƗK7\s�c��b8�H�QOr���O3W8�<P�"$�C��p9���� ڴ6���b��W.F�(K�
$@�K�I_�5����%Q  i(7`�*r>V4i�KN�!�%S���$O8$�"��yx�2��I�����!C�$��Z��W.",���T��>,�g�$�0>���@"G-x9!��U�Y�xBcۃg��е@2��R}%�x�M�)q����놺`��d�6��2��P�j��dU.-�����\�A}~��&���	�'���"��d��>�����R�ڢ�w�謋fo�:9h�!�!��/L��|	
\G�NQJt��d��ʌyb���f��ܴ����B%]���f��kH���z��I )<T��@���\��ȓuߠ��[�ND��aC��n�T�ȓV�l<r&O�.e�A�q��*uX*���F.�C ��2�LL�W�B�B&0�ȓ.<��a�Ig�Qy���#=�\��2��!򲇑8��1��5;�y�ȓ ��|�i�!U�:K��PU��m�ȓy��!9�f�<|+�]�cl�<I�,Y��JB!�0���f����艿Ob
���F��q �; :����S�8v~y�ȓ'BRx��ؚ4%�i��˛�"ȅȓ�}�'��J���#�RM{���ȓ3\d���Μ
K��I��k�@�4�ȓe��KcGC�1�^	���:p���
��x���] ܴ�$�/(=��'>ڑ�3@Y�Z� �*S?	����r� 
7K�K��YZ�	۸J�.x��bv�`&ӄM.52g$W�,�ć�dS4��6LHo*�P�ӿg,\��ȓw����F��`B5h�c��-��H��h��;�@�"��Q�U�*� ���g�|�� ��d��]آ�?����ȓ���I�
�}�4�P#W0�фȓ�,�ׂ�+?��Ӓɓ�k��Y���7䚞D0&$ �LZ�:�$"�"O�0a����$ْ�(_�<Q���"O���FT�xPΜj#&A;��и3"O�A�̑/=l��{���p"O�= E�Ձx�}���J-m�����"O���@LO7��7 �-
l���"O>��Q�xt�T�D�9A�mBe"O" x�E���`�ҹM6���"O����C�}K���B�	w�����"O=x2d�-"��ko�ƀ��"O����U7Z�"Ժ��t�^ À��
w@Iۅȃ.\���0��'��C�.2J%�uEB�i�*�y�{2�t~�O�2K!�e�O�*�q�'?^��CA�X��M�3�^%Y�TY�Õ�@<��ň�4<��Q����g}�
 �����kڀ�k�����,yj/޽���-�>!v�+x��A���Td2���j�� �ř�ꑰ#eڥA�OV XT��V��!��O�N!*"�C�h :mH���5:��Ѱ1\�@�I�ǮՑ��x���Ⱥ|����M�:K�0�"�T �d�:ݶ���dLC�~n:�ӿl�4�[bk͋l��+V��4y<�öo����N<E���π X���Όf��ݸga?��'�u���'���ظ��$��h��?=c���ds$`�ǃTN��n}�nQ̓�M�0%��ƹSO?�&>9��
I�$�F��O{Ԑ�F<ufR�(�'%��IϚr�ʥ���<E��`��X�t2/50>01���M[KۮC'����C~��� 
`��t"SLE�r�m�'du���O�2�V�O���)�=g68���T����q`�b,@�{v�SX≦V�Z���^�/�E��fi,�3��b"�!&�\@1F ��F�'�b>e�W�O���Ј>(��U��g!?�g�Q�|Q��'��E��'�7.`@�OYHoz�d����M��E )�-��x��)ʑ+��B�j��G~z1�VQ��R��d�D�'��O���M~2�I�"�l!AsJ�`@P���Þ�3!��"�V��~�B���c?����ᣂ+ؓ^��AɅj܊<`���u�[�*��9��T�T�	�m�.���We�OQر�!�7m��X�a�-P���]+s}o��:zP�E�1�a�$*�g���4�N>/��Y� � �P�ϓN����2��5��8)�:�Y��s�F@J��9UHd����e"O�Q!�o�e�thC�@�a���u"OB�Jb쎈f/������p�6�3s"O�ŀ���WގH��%޶@LH�E"O`lۗ"GV��rEޑuz��"O9��F�($T�( Í� �C"O���L��u�n����߁e��Ձa"O�xre�*h�����ӹ�� ""O�����0"詵O��=�=�e"O0U�NӋ��HU��5z���"OT\�"CIl,9� U�g(�=x�"O�ѣ�)�h��!���%�$	 "ON����{Ef0RF�Q�^FD �"O�8pG���̎lꆇD�j���B"O�@�뉳6������u���"O:���uT�c�K"H��̓"O�}�T"�	,�a� L�Rgn�"O\mXD �Z��Ӧ�O�3V��cG"OU����f�=��	6ߢ��"O����!T"Q�����9s�:�I"Ox!A�H�4 P��L���p�"O¡�1��<W�ʝ�S�f�~�#&"O�u����F�����y]j9aw"O�Г�j	t2B��֯�WGep�"O���f��k��8b�0U"��6"O�ȋ�AL#��LX�g̓3Z�e"O6͛�G�/�xeB,�pH�G"O(-1���z�H�CF
�X�j"O����ۉq0���oU*V�D�ca"O�5q���w���0�O��os��A"O4�����3�
8�OI."c�("O
�ɤM#L}�M7n�\�\�E"Or�c=A��)��K)*B�0P"OX,��F;s��9&�<F0��"O� YAI��=b����-N9d�� "O��c"/�Щ�*��`;�J"O��r�G�N���85)��y%��"O@ec�ĚF��0c(�	pP���"O\��w��U�M�d�A���;d,&D��pX�M�~5�0�˥}*X8�D%D�Ă���}�F�r%@�3_�p�a$D��ɑ̟�r�ܼ��5$�(��B'/D����暤)zr��UGK ��-D�p9d�D?C���4.��>	q@*D�8ʶ��l%�ȑ�.̒W�h��E(<D�|����I�)�$J�q�Z�z��9D�����7�@A�Do�"'4A0UO7D�6'�����(��Y�E*�no�<I�kD1�R�r�lҺ&�|90!TF�<�����y�(�	v��6h.�t��@�D�<� ���$�|�aCRl�5sd)�"OH�(�j�[�Ը�.�L`�h8�"O�q4�R�cW���-�;Nܵ��"OV��$��jt
�X/H��0"O�p���4%<�`@g9n �)��"O��Ĭs�T��b��v�H�
c"O4D�ׅ\74�	(�Fsu�5�G"O��a�� ��4y$EW _��|x�"OJ��,��t;����*˻1W�$Z "O�I�ë�|s�KL�BPfe��"O �(7��&Z|�@�b=�#%"O�H#�* r�
�jE4X�X�ٰ"O\� kŭ�8XBf�ӱ?]��;3"OpŸeg� 7̎�Xf�r>��r"O
`��-]�:�L��f��N� xK�"O���� �u�(0��E�X�R��"OR �'&�v;�Q8�NG�����"O�@s���T�Z4�͒s`��2"Oht;Tٝ|�V�u�O�[��h��"O��䯝3%j�Փ�bGM��5�"O�SgM6��� Q��)���+�"O�����W�}ZbAN\����yrʊ� (�a�2��:�1��-��y�#Ǯ*����!��w�q��§�yb�F"D]������6ip	�@�ۃ�y�B�8e�˖��p�S�ď>�y�m�i���X�&:|���(0�@�y��<MSV�
��?\LPvb��6D��B��tќ0�+	`Xxd�A�6D��1�i��z(�v!��3�p$�n6D����P��E3Df��\d�`S�5D��'��% '4dвOO�W�2��k5D���R$"76	�D"��%�\��4D��/�n�Rts
�.Y\���2D�H+�ND(�.	K�aヅXK�!��;��5;Qc�#I�|��ē�K!�$S�Tg&�B���(`����G�!�D��bP��M�v=R�����:La!��3�J�L:*1�0���H�N&!��[$(�����v�����}!�;}���AA�B������Fz!��:x��A��x��01� S�K^!�$Tm�
�+�ɶduDq4�T�HK!�$I!QF�4�4U�kx�#@��
L.!��^5T�R!�6mN�0v��<!�Ė,F؋)�j�4cj�c\!�$AB����f#��}ghq���ȁ`J!����aGE�Ya���3C��]h!��Y|��,��l�b��=Wg!�	�-y���!b�Sjܸ�`A�z�!�D �(<p�0���1>49�T`�#�!�d�&
�ɈCc'���Pϒk!�D�)H)�Ä�-wVAQ�׃	!�	�Ac�l�v`ȟ�t�`Շ�1!�>U
X� k�"RҌ\��X��!�ֆb�n!��L+�������!�D�X���c^�W:�S՗�!�䟐I�$�ȁb�)�t�w��X�!��ʚ1	��e�
x����!��Y�!�$	t�J�ҧ�i��
�o�6*(!��_4�B��VET�	Ӫ�hp`A�.!�$Z�1�굡g��=}j3�eP�#Q!�$O�(��
�����'*�!���P���(	}9�Ò|!�� ������	 2�o!�T(0"O�"�ZI=µ`�k٬��]��"O�ɻ4�Ԋ]�Ƭ#�l^M}V�k"OXI��<WvTL����^�0U"O�$P��խEX��:�Mpl���"Of�c�D�ӵ�+f���"O�)�ET�+�*��ТҪ	���u"O����\�>0f�@��7t�d��s"O<��2�5W� �s�MI��>t)�"O�4�@E��O͘��C퓡��ɛ�"OH�s��Ɖ`n�ܸ�&�VԲ��"OJ�Ђ��#8b坈�4�H&"O6�۶��.<X�{QDL/D�L��a"OhQ�1��[�z,�#�8�:lʗ"Oz$B�k�5WT��D"�t��(�4"O,�ӂ��,m���PdB�~&j1��"O\��.�0��Aa�6`u�4 D"O�ɨ`�	,�N�۶�V
a$�"OV9  fV�5��� J��DG�$h!"OL%#F�1.�l�p�I�5@�$"O���'-�8!�ͦ_����"O���WKI�S�*�8�,p"O0|2U鐝{�aY�n ���X��"O����#���̸J6N��C�"�3S"O��H6i��L�`"� y�r�C#"O�b%�
{��PrAX�m6.yX�"O�Y��,3=0� B�/,X/�\B"O�<9�	XW�T�qF�BS��m�s"O8<�c���B�ɔ�ڴa�� a"O��X�g�����o">O�!�"O�`�vE�R���?o�,��3�y�l�	X"D1�gDL�4?��8A���y�\�m��%�IH�����]<�y��J='�$��� >�i��Ź�y��@	}���ɒ
��8��#��yB�K%��3��<�v�
d-��yB��	L���DmM#m�����Ǆ�y2�^(`4�]�EM	J	>�����y��N�|܅i䆒4m�9 wo�8�yr@3�T� GAD�����A�yB �Lufi�0�ǐ�T=cqF�=�y2 �c��$Ra�E�x�*\H`���y��j�x���v,��i'#F�y� ��f�Q�J�o�Ѝ���Щ�yk0���čk��)R��Ԅ�y�I�\�"X���Z7c�8Q)fAI2�yr&R>a;����>O,���UoӴ�y�ņ0j�̬!��)AF�E�4�$�y�-(P�I!��=C��`R���y`�"D	��B9qz�К "�yA3*b�:h�	q��e�Ǘ��y�+NC���4�5f5&����1�y�Ε�%^�u͕*[_*a�Vc��yB�:&�^������u(��y!�^�r�P5O�%L�-bX��y2-G�oO��	�,B�ı���Z��yrf*u���se�J�b�B��.���y�n� ~'�����'W��Ȳ(�5�y����)��DS���"	���2�я�y�ךN6 5H�Ȉ6K��l���H,�y�`�P�Ba�È�n�9�B@��y�@!9}�����D�3.
�1B@���y��]�w��R�݋0�~�k�ƛ��y�IC1[A(Yz�N%�̘KDB�y
� Vi;�Lʿl-r1��ӡJn�r"O���V�&�$�1`��?4���s"O� i3(�:���Q,ݢ-�=j�"O��Ig�R+]�vlB�+�2��b"O4�ЫPx|r�Pu儩E9� U"O���̈́kh�QÒ�R��@�"O`y� ^ gB}�1A�X�21"O~z�J��?���ul^�[��(K�"OPt����Z��$X����("O�u D��9�p���ŞmB�3�"O�])��\�58�"�!��,�A"O�T�%��u�9cg���s�[�"OQ�LU�o�l��A�rBX���"O.�K���&���P�C R*���"Oʸ[f��d�z�gŅ�2��4��"O�����KQN鳇Ô(�^]s�"O����Qg-�9q�bE=����"O>�y�蝙3��-�PA	
�B�0g"O�Y��~`� ��4,���a"O�YzѨA3Ab,Ԋ0�/���J"Oq`#�6�LP�#TP�Hh�"O!�$%[�i��=�2(2?��"OLy��   ��   �  y  �    	'  11  t7  �=  D  HJ  �P  �V  ]  Sc  �i  �o  v  `|  ��  �  (�  i�  ��  �  `�  ��  Y�  ��  ��  ?�  ��  S�  <�  �  ��  �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6�F{��'O��V���&�;�+0:��x	�'%��"J�[�]�R�K2r��"
�'Oe#W烹�R}aC��z��
�'��;��7�������L	�'�:<*b&K"4����M����9	�'نx!c̓>�D �,ݻ2zX�R�'��@ �F�9<�m�7I�"+�a�'ր����>��Y�
�%&���'��0��3L�r5��M/� HJ�'U����J08fx����I$p:<���'6�D�)n�N]	0��K'~8K�㊵�yŬJ�Da3gǋD|H����פ�y"*@-0NPI�-@�=�D@f���y2-ݘ;������H����u�O���ޗd���)�S0L!��҇���Y�� 9b����2?qEԁ#�]1Ѕ�'?/�tzV��J̓��=iWɋ'Z��(���Z�:H�p��P�'a��G�ԧ��/:9��ƌM.��s�B<tK&��ƓK��8�NG�&�����!x8��2.�L	�I�ǐ�+��F�A����ȓGs(��4��>Z��$��\�~�<	�����.&̕Q�/B��nͺ6��bC!�˦Yҡ�'��h�T��^�!�J�8q,M	Q��d���Z6�D-!!�d���6�K��2Ĵta D@"-!�$�jU��j�����c6L!�� ���h�#]�3�l�.x�2xP"O`����3Xwr� c˔�=�(�"OLx�W�D�B|�̭5S�8*1"O� ��Ɇ����v 
=>�{�"O0��5��9)����C-<�#�"Oڤ�[�Y�Ȕ�A!͖yq�q��i���W�+�P� t�H-�<5��˅6s�a{��d�@�t���Og~�rt�ď{!��2\|���H%9���CT
O�<��!�O�@�7�=��4k�� �d���"O�=���_+L�(�Pd�͸L��uip"OR�8�Q�c��-(�%�
#!��"���[���)	>Y��t���M/L��`jV@ h��$<�O4����Ǆ[�PmA����q�詚v�')1O-Kq���q�g ��LL�"O�Q�(P<l���dK�iذ��"OzY���)}G��
�%V�$���{s�'Z�d�<�Tl��X 2dX
I�>P[��t�<����
	��0���	R� �BF��ph<�Rg�f�mz)A��L��I>�y�I	F����pI�}ܤ5��V:�0>�K>Qq ʽJS& � �۹)ך5GeUh�<�M�4�T �,\�h�~D�a�UN�Z���O�Z\�@���<�dnN�(�ZX�'�*�f��:m��`3�l�&Mp�8���=<O�9�d��>�\9�V�;o<�|�O�8hEj�#q0�)p�Z�D�P��6aEkh<!C�W�#����U����b�a�\�<���)��ӬY�L��u��T�<�3�[�u(��xRB��Z�� G%Q���'��O0Mj7
��I9N%c�@���(8� "O�I(&,�'��1��L�6{�
����$�OL��DO�K��ra��zP�|��fΩ^�Q�E{*�8�#T �h'�=
T���O��)b�"O� zD��9IQȤJיL�G�':qO�(�ӫM�P�4�
pJL�D�^ ��"O�Q����R��D�?��R�"OD��'A8w��F�\,���Rf"O4��
�(j��u��I�w����f7Od��$W��qf#:l�z��� :!���."=���3"�8v�\0�ڎ2!�䋜&��ԋ��܏	�(*0 .1!���M!.�۲�I6nd�)�AB�|!��:ʉ�p�TH� �@���!�$Aq�, ga.900qw/�<�!�_�X�2��D^$wI.������~�!��F'���y��鄈B��ǐi�!�dͻr�Xw���3�|�(��X��!���P�j�r���%��5�����!��G7o���J���je�KJ?m�!�$U,�0,�Qc��F!���L	{�!�d��C��U�"v��ra�9h~!�d־h�h���T����Ko!�Ƶ�Px�WbA�ry�勇Ìt�!�䖺a����?c|�ژ4o!��P��x��&JX3�t��A��r!�d@�����R�1p14�&!Q�F!�Ւz�$r��X�|�;�
�1�!�S5�֐WMƓy��䋵�T�!�!�]$U�Z�j���2I�p�5�ɻI!��W�Z�0@��j	d���S�!�:{|Dd�Q�0�֜��ǔ>A�!�-d䨔�`�Ś� �#��a�!���?�}�v�U�l���ibdM1|�!�� :��k	,nE��j���B�&��"OZ�Qj&t)2�b��0=��a2"Ox��%�N�=dIs��	�|>D���"OԵ��Jȋ�L	3����Q�|��P"O|�Hfߡm$�3sg��/"XA"Or�Ш�	&_���ү�l���"O����L���2��:F��|QD"O�l3V+2���TaV5'�
��"O��$L�hb<D���Ûo˺ �"Op�:�E[�"�0 ��(TN}�7"O���Ю2o��b�	�~��u0�"O�h�Pa^�z��UJ��	3_��AS"O�-e���
����R��=x��#�y2 G�9��+V�mpv��7�yR!�\�8!��͉���V�`�j�'�������#GM\�uSe�'����.�	�>���B��hXpU��'g�d�5.O�V�,���`�	sf���	�'1T}S#�H\�Nsw+Q�<d���	�'�.�(�	�8r�Ll���T�J�JM	�'�\�YV..�ܰ����YRM��',�ā�Ȉ���:��?{vT�	�'-����H=6���L"dJH	�'�`�gF7J{���L�p���'����T�����񱫍�?SD
	�'�n��i�Oa�aZa�Z5�l͊�'��Ue���"�PlJ�.�j}Z�'�$]8�I"��1���)^`h
�'�xmt���	����������-D�$GK�,��*u�H�H^�[4 <D��Kä���ҍ�����P�A5D���lR�_�:|j�a��1�I�ï=D��jQ*Z%0��з��4^A.|�G#9D��B�% 0OΨ�JC윎]�R%s�I:D���!�(Y���G��;,��[�i8D�Ps���-V`(LԦ�&@�T�z��5D���p"��=�j}@'/X�R+P� �!)T�܁ԦߌG \$8#k���:싥"O���J͙n�E{���C�~�"O��ʀ��-�(H�6�F���	�"O�Ԡ� ߂qk�,K�j՞_���ӡ"OP	a`�ì;$*��&I��RDBk�"OƘ�T!E�s� }p&�/5��0R"O��Hcǔ@�����#���"O* ''F�m�ȥ	�M���	cg"O\�95�T~+�= fLH%<G� C"O�S kC{��fK6D�%Q"Or0�����Z2��
�l
&G+V��b"O Ɂ�mG�[/,,#�#0&��3�"O���'�B?�թ�B��Z�"O$���Vd��˔��&G�f��"O�d;��X�~����s��4W����"O���%��EYFd���� 8(�"O�\)u_�P�4Q���l4��r�"O�-��.ԓ;��}{���%�	X�"O�Q�'D
^1Qsc��V�S"Od�c$Rf��rd�',���T"OT����j�p�� A&����"O�@��?qj�=	!`��Z��9��"O,hP@��$E�Y��	!H��\v*O��W@ׂ[+�Ո��&@48���'�� �Mĸ[/���mU8 d��'>^Y��NdCZ�u��?}����'�x�1$Ŗ�����1d.j�.@���  A��䕃 _�Ȅ"�L����"O��P�n*@5E�ۉ$���ic"O���e�_ n��O�;}AL��v"Or` ��I�|�MV60$Ґ"O�:aG�\����U��
5�d��'p�I���IƟ@�	�����̟X�ɝu�5�!�G*L���dl�t�zm���l����h�	�������0�	ǟL�	�cҠ󡫚B�FXB��ԀaH�a����\���������џ���ƟH�	6"{�@���0&;^�P��څMخ ���|�	̟H���(�	����Iǟ(�I M�"���gK�8�X����ȗH�&�������şh�I��\����l�I՟��	���@3�D� [�PH�	�<����x�IҟT����(�Iş��֟��I0!x�b F�� ��ҠVM��	���	ß�����ޟ�I�8��"��̩����C�(�K$����4A�	۟��I���������	���	�h������Pd��moJ�1���*=����՟h��㟼����L�I���	���	�>�@����?3�&)����m/���ڟ��I�H�	П��	��p�Iǟ4�Igo ��ŷ#Z�\��v܌������	۟��	ٟ��I�����ʟ��	<y;0�wbʗLp�I�1f<��	ޟ�	Ɵ�	����IҟT������%�\��D�g%: X��R�p1���	ʟ���ޟ`���������Rش�?��u��W
#�j��d�^%�4�3^����My���O��m�:>�4��RR&�I�=z�h�%.?q��i���|��y��o��Ჰ�E"!{�x4��7�	���F���	�B��8B??��H�

-� .�ԅ����̞�b�����)؎��'��Y�xD���X(P�~�S�fE���� �,<9�4R���<i���ce���3"(��	��^�%Le�dAX�J,4oZ%�M�'��)�4i|8AW)|�t���'J����fW-"���#c�Ԣ�KK4<g�9A�'Z�����'�(�
���#)�2�1`�՝O�);�'���i�	��MC�	�@̓+xt#�l�������d�=#,%��R�>!�i�P7Mh�(�'z�mY�� %u+>������wZD�s�O|@�'�8M���85�)E:H®��7d�O�h��Z;GPL�Ɂ6a��)"�<I)O���s����!Ф'��i2N��q��T�to��z۴;MH�'@�66�i>�sЉ\�Q,l�"NТ(�$e��lk�D�4;����'挸��A����V�'��d96�f�$��GY>X�h�H�4�\X���+Ϛ|��O�P0T�M�����8�.�P�*ܦr���q1�K!B̅�`�
�Xq�Z
%�����#���I��A	���r�·$�6P�B��n�4dPP�^�7�@�����7��a�7�F�un!�u���LM�r�g��FVt��`�`��B�/j�i	��F�"�Ah����`\2`e��n�Hc*I(A&�-{��Pc�i���}zå�.�)[t��#�P�o�������L���D
]:
�薦ʺF�X]�1/��/��	������VM��Γ�?٥#��+a��Z%�^��h1 '���.\ Zh6��O����O��	�@�i>	#-[O�\���I?Lx�5sd��5�M���C���'8��y"�'<���o��<����zt��#�eӪ��O���Lˊ�$��S�T�	y�x� ��r.�,@���)a����4�?����?qg�	U �SܟH�������G��������_	�PH�$��[.�i�ݴ�?��e�vJ�'mr�'�ɧ5v�äsp�a���4��K��M���>8���?���?�������O��q��](x|�Ӥ����1
ϊR�P5%�0�IƟ��IO�	Ɵ$�a�B	z=ĕ�-�(���ء �y�b���	��,�	Yy�I�s���E�Q��8�\����D�vw�O��5���O��L��I�Gj6 ��#��2�A ��;\�듵?���?�*O��x"b�f�Ӛ�������G @�&4�J���4�?1�����?�T��C����%<b\����5g8��Y6%r�����O��kv(�������'*��$�"�\��4nH�Q��cňF, O8���O5��C�O���O��Oô]����v�h������@�3�4�?1�<��9�iŌ��?���=���_���q�VD !F)E�5���?�#�^���'E�L<��̙/U[�0���ޟ9-X`�Φ�� ����Ms���?���RÔx�O�|v����"�rd
��T�:�07����҇��O���O������˧��)XJ&�����S�0t�3k�:US2mlڟ���|J�fyʟ��'�d�P����l��N�*���O<���(������'��d	:E7�]��nXA�V�iF��*���'��R2X�8٨�v�,���ȼ�P�#��Xn��#���M���BX���K>���?�����ă%LvTYDD���ڬ�C�M�%-ҙ��G�Q�ڟ��	�l�'k��'�p,c�ęv�]����%+�L�����S� ��ߟ4��Oy�N[����S,�졠�ɚa6ڌ��9���?���?�)O����O$�Q��OZ��ɽt����r���Z^}��'�R�'���s[�\�I|br/��
x��J��G|�I�Ȏ&n���'�bR�0��ߟ H��U��O|���b
�0K� ���#&��@���l�>���O��_°���T�'�\c��uɢ��6�b�Q��.�aJ<q/O$�3o�O�����3� Xt����>p �f�O�|��|R!��p=�m0O��(�Tr��f�<Y6�Ծr���(�m�hn�0r$�(`�P�S�O�+�>�!&�$I�dТ6�P6cΌm�h�|F��2��&|� 5�$�!Z���7؁M��̰�iY ?�����NW�Mx��e��e�0!�7v��I�݋Y��l�gj^�-�5�܋�6�y�jܜ(�Ѝ�acIu�8Q���\�fZň����?)���?i��&���tY��2��d34f̵�������`��!0@yS�Ǭ�p<�����K_�1�v%	`�]��`�Q?a�k��i�y0jƽ1��xr��XGp�q�<R�<�R!��u$�G:��'m���D�O�����;����x�yg,ɖh�@h�ȓ+���k A4!��W�T:4E��@�IQ��Q����Ȓ�M�%3%�b|Pʒ:�����	�?���?A�ct,����?�O�N:u@̀<��RĢ2�BL���ޮ��񹷡J��0>ѕ(��P�b��u���K�Y>f\P�)]'Ap$�I�`0�O<���'s.6m�ID��d,#��a���\���%�������?�O[P��+<).�{w� *`44��'NXpR���--f�w�5n�YK�'���^Px(n˟T�I]�t��O������<�0�1�Q�W[�D�$�'�B�'��i��B�]���vUf}*����� %s_شJ7��K����	5�2l�Y����`b�'Z����%-���(f�8D3�aDy"���?����?!���i�%89uY�'�5< �!����!�r��4�)��<���z�@D�P�Ź(���Qօ|���I<�slփ)�$蛵Α�M��H D&Lz~"�'�r�'���x �;���
��8/8(��'�L��P�G����Gܾ6�]��'���b���A(u`���an����'%��h"��}�н�P��+�H��'����3ȏ�bu1��Q�9GJ��
�'E8�'���x�.����H:*��1��'�h��s���B�Ħ��/���
�'� i��6Lzz���� �d�
�'��Uj�T95��x:��ԵnK`W@�<�w��\�B,i<x�RĠ��R�XC�#kF�cq�QK~T�#��6�HC�ɻ�t�І�8�H�;m�+tB�ɒD�l� �Z�1�,������T�"C�I+'�.pˑ��7��a��F��B�I��t�Z���	9���"�߮�dC�I6"��󱥇�L,�2�B]wzB�I�F���
R�E|f��ӑv$�C�I�t5z�jE���sr8Y֭��C�I80Efx�QdD/h�`d�6��
�VC�	�.]1cm��n��)/?@C�I�E�y�w�">4v��ԁ
��B�ɖ3�h G_�8?�P˷�;4�.C�4!�xp��)E����ys�C䉣�pȣ�c�e�DDp&�O�@�C�I�[�>%c!��\�`�O,xTC�I�DĖ@!�~-�H � PC�	&\6P�#fi[1
�H�P�
�/C�B�ɭ_p�YrC,	�C����Z�,C�ɰP�:���Y'6����dڬ2��B�	�w�j�0"����Ac.��{y�B�I�n[�᣶��0����Ö	��B�D��a2n��x���ԣW�~B�I��=B�E��C3iL��W [��y��E��J�I�$\�W�XMө�y�a�-?�����ۓU��(Ӄb��p?d�\��Mc�E(	c���!���$��|�<) "B7�:���X�%����k�y�'�@Eꢈ@g�OMH � �\bҜ��Oս0�2�P�'P9æBֱe�l����V���'�dyU��V�S�O`6��Ѡ�<	����O)@#HtP
�'>�pѲ��|���3!	P�2�O
�
� :�p=���G;�\0Bq�P!�F\�c'_J8��p� ����uɞ������ N��,T0NQ`���	��Q�m�1��NB�YX�p�a��hv.������zޭI��#?!Q[;-u(�Y�D�'.��yB��E�?��f�F8!���`��u�����=D���$�Wd��M#0H
\f��F˩R~�B`�bD�O�'T8�1�������5E	����nؤP�󕁇X<��ܕ>ɮ����-/��a鐦� 5�4�'����-U3A� j�/ɕP��Fy ֡:.mQ��L�3&����.���0<�ua��5�3�Dԧ!��cV�Ȋ0�J<��h�&vKS��'nFD��3m�Qj�i7�O���RLƜT�
܃��>aF<�r�����=�z6��V�
ț��4��<ڷ�Ѻ��!a4�[V|�p"O�t�VA'NvU؆�� N���Wk['-�q�mO������� >�� S3�:uq��:��ʶ�ք1��O:tu
ݟt}d�X�/��TP�a0�O�!L��Iwi ]�fʟ������Z�Q�,p�G�!�&D�$�C*$0��"O�+3)�q�R0�� �	5Ֆ;�c��JY�Â�] ��a�ְ\[���D���x���	� m�Tۄ������O�$[����'�$���珔	68+�խ
[P��=�'N�d#"��9 :=�&Q� U�H��WA�<#q�P�w�ԥ$h����s��3r7��zB%�) `��U����;�|d���\%�����*Dg2�8��GM|e����5e�bip�B��6�#��l~�b�*w�l9$O֜����OL�'s��E���)㪙8�bI�O�ɳ�*=DLS�ԁV˛�Lcu�B��5��c�@�4 ��py���0a��P7F�6�L&�'��WT	b��`�D���G/��ե#?������
�:���)�^�P��?��u���z��ɸ�h��A����b%D�pf���,Ө ;�����:uk�)��d�@�,��rӡK��91TL]v���	�,[�d�R�NX�	�u�P��%.a���6�䑁��%sA�:0��b�(�QIA>��Y0L��C#ɧ����֥Ӓ���[�s����B� ���O.ܚ����OY�4�E���D�^}�� #���O�%���ÿ/���䗂y���1'Ӵ��2sO��	�y��#��?�;�/��4?ͩ�_;J
|Y@��k-��b)��yR�4eܮE�ԞY�Ddp�	A4�?Q��J$1^@�I&wD�Q ��<�ӾD�?)kp�
+Pr��ef�D�pC�k؟�q���5h���q�O�"g�c��*, M�"ځ[���	�6T`�`�O�)]�s҂�$j2dk��u `�Ӽ�xM�U�.�aS�Yy!� �&�Ǥu�%h�4��%�D��9|���zgKc&���j�H�1���ol��dۊ%W�̈Q�q픜)�I�*w�I���i��\��P��eղk�f�I{?y�'Wf,3��R*&��5M��8~�@x "O|]�'H�zb`jva�u�̘���Ǖ=� �#nF?��'���OM.�#�F�9p0�ݐ��$b��� 4���%��Z�$�����a��У�o��K�8MSD΋mN2M��OG?�'��8�0�](�b�8ST ��{r"�!}&��C*KAL	�0����O��7��>j�PXfJX�y-�:��it���QaGx��+�/�	5�@*@�ʨ�vE��cJ�}�x��	<Q*`��:-P^��Ţ���(��h��J�V����B��I(���~��O<) ���$�\�S�e�+3D�Y M0D�H����p���hќ"�ȴ�S��P���#=�	��?�3O�i��bh����߼�@�ǴE�V���O�8R�xh���\<�D��W4�]��t�|�S����Y�`9sAۥ	0rŗU�����O��	���'�t��D�yxꁑ�dC7;jD��'�+�:��-�ԅԮZ(ŀ��fP����Y�8�2`@�?GN�b���P�-�A����=	�F��H������W5�&�d~"���K.j5:5D�	�ީ�� :ḧ�v������(� �S�c�_�<in�t�>��V��Y]	�Df_�VamB�瓎.�n��=�O2�1P�ܞ�yw(-H N[�.�=+���2� �xr .��C�Gt1b��q��cȘyM��bW�̍yF(�3��<�𩀇&6��<.tL�Q��#
0D����H�J
��d�
'P�%��-m�jTP4�>W�dɢ$ۑ�&E���KZ¥[�G�j��[$fB�Y�P��d��9(�	MH
A��� ��%[���TČ1��O&x��j� ��4<m���} ��qg��[��Tӷ�X~��ȓ6a ���h!�Q�%����I�<��X�S06��0�t9��. ���>��R (� M�z��s�C ��9D�d�@ T&6[8-�BF� {��$%?Y6ƕ�J����D����0ãE�
���n�3@�~��&]���Ƌ')W�q	��W�*#`M����3�y
� �dS/�ޕ+EB"T�V�qq"O�=q��;.b�(*]>�t��"O��H��/7��%��K�ߌ�B�"O�\pǌ�j\��e��3.���"O�u��K/G�$�q��ј����6"O����لUm���t�?��3a"OBQ��\�]�����G�V-j��D"O88�U��,b�\@�OF�JL`�"O�Ժ���[� 4r�A�5fH)U"O,,[sm͖.�� �k���͛"O.�9WE՞$3V�;C�Y?�4@��"On��c�"b�,�@E�۞-��� "OD�R���p��� �D�8;�P貣"O��v��� j�����K����b"O. �� ���`qB��J�`"O�d�3,Z
|J��5dr��R�"O�,��C*-\�$��dB�LL�೧"OJ4�6R\��B��-�@��"O�Ĉ���3W��<2!�ϙ��=��"O�u�Z�.�js!U�乐�"O ��W��2i#� {4[7��Eq"O|��f��&���J@C݅M�VT�u"O@X��S�R��t��+X�xӊ\��"OhP��#�A(�.bzE�"O���a x��H�M]�6R�D��'&��vJL
d>�=2W"J3(і 	
�'������!
�0r�dH�4wl�'0�B�Hܶ*>��C7��2��R�'#�tj�N�z�jl�3+P�$D�-k�'s�(�����bM>X�B#�5-�*@j�'��dC7&�3b�4t��I��8��x�'b�Pa5�L�D����=�%C�'�W`\ $P�I�QB]9Ė�c�'߰�s �5T0-���'z�d��'Nh�;c�Ǐ���7Ѧ���	�'G�-[�$�
�>I�r�|�a	�'F�iCЃ��8p}	�J����q�!D�l��k�X� dC�E!n�e�g�?D�Ts��J�l��*fAC�[���K+D�R�A��d�x�I�))��qk-D��Т�u�J2 � �o��`,D���e��C�N=q�,�-9��!/(D�䚀��w�L(ӷ+S!z{�`�Sh3D��K�a�RHFY�kͺ,߂t�D3D�l
��O>%��Y��"�Dԃ��0D� ��90=�����Z�p�A�0D� Y�Ξ�^��b�Țg䕃�.D��#po^���U �X"=>D`�m8D� )ä�h}�s6HQ�X8a�E6D��׈�61���aQ#I�QX�;v�3D���s� YL:̪w�3|x���0D������'`��HQ?��i�h,D�d��cZ�Q�YY7� *�Iw�'D�P$��*��L@���LR��벡$D�Ī�kpҼi	fOUT�F��n%D���6L�!������"�4��B@"D����/|�bUs���sX�	�#�3D�9%E����>4���d/D�JP/	A<\�O��̍��$/D��QTd8{�|��h*��y�`�+D�h��F.]]�eR��K�b�Ӑ�(D��)���L'@�8$�?��bAl%D��8TLۏK�>��r�F Ё���(D��:�M�p��}!���%`�ı��*D�� �0[6�*k����q�S�_2(��"O���2��ElT�Kį_��=Z"O��b�A!	��S���W����"O�m �d_nN��q`��ל��7"Ob���IW
P���vȓ�\%��9�"O����'�v�R���M
�B�"O�y����L+̚QQ&Q��"O���F�	@n���b�8[�}��"O(Љ@�\3��r��}C��3�"O>�ac	҂;W0$ �ߠ!����"O����'�B��g��3lҍ�a"O��B���<Z}B��e�'c8I�"O�U*���k�����ͽ)�d�C"O������0����]�n�Xs"O�u�V��\O,�E�_�}�"O�L	Y&	 �T��9J�F��"OFL���� :~q���O4g�$4�"O��(��F�@�`�a�#=
:DE"O:�i���2#�|�Y��K,L	0-��"Oޡ���)>jy� �85�
""O�I����:x�@�Զ;TS"O�S�]Q��agn� g�xm�"OԌ+dGi��Ò'���ڒ"O�����,m�s���^��"Op�*'��������Pd"Ot����!z���	E���q!"O�ua� Z�[��40�ȕ�y�ȉ�"O|L� (C�z)�g!�5>o�M9�"O���Z���o��i����"O(����ni*��ț!��As!"Ov(�s͡�7g�c�@(a�"O"�%D�c6pi0d��X�B1ȳ"O�I:����Ui5H@�V�dP"O�6KÊ��`�M�3z�]q"O�5���
�z�Jd�A������"O\d�F�6���ӧ�$�����"O�8i��J�?��M)#!ԋ'�@@��"O��� ���U�(�����~�6qs�"O���r��]t�`vɓ"~f�9�"O&�Y�)���iT�ƈ t\)C"O�m��B�>p',BU(кur�4�"O �c'����haG1(f�S�"O�`�&
�'�|h2@�OUap�"O���ܵ$�n�A��
�3�p��"O:��b�Y�p�v9	�.\=TLQ� "O�|�1�� xk49+D=�����"O�(�Ë߯1׀����K��v���"Od�ī��v��t���ĵ;�px""O�𳕅J5t��E)��T�C�}�"O~�j��w�l��H���u"OF]���Y�+�����'tt�u7"O�I��ƾ��u�R枻F���"O����&,��kQ �5��{�"O�!"�ڲ*n�Ђ�oC�a\��
�"O�S)��q|.i��EI7MEh9Q�"On5pV
�>Q����J�%,:`	�3"O�+�J �2�l �U�Y�$�@p"Oֈ��3Tܶh25��=�A;b"O�1#���A|�q�N׍p��"O�1c Dc�U@��6E���""O���� Ҡng�M� ���<N��"O>80�$�RKF�;B�T��Q"Oz�F�5F��]��nB�,Bt�R��`�O����P'k��1�Gl&~� ��� t0S�D
�[[̈����C�I�""O����ðzâU2�˜�J��  "O��(�JP
�����T��"O�i �$�c*�Lᖀ�2K�
*E"O�hQ�D�b�AQ�-Q�fV��6"O ��ѧҕ��
q״�95+ID�!��z�p�(�op�uJ]�?�!��7�����1Bl�p�QJ�Lk!�DJ7��Q�<Yġ�v�A!�V�{i��Z��^�yQL1��'_�'��|bnD9<�\�K%�(&N
�{�"ի�y�AG�J�y�w�8�ޡ�C���y�
�e�D�RF��7V-`F+Y��yr+[�+���t�U�D�hu茗�y�	K',4H���m� UB��t#I��yR�8Tjz)`�N8� �1
���y�ȓZ����(��v��y�O���M
�'J\#��*I�
�a�o�847����'��!�"�� K���W恈]�4Ej	�'fv�9����
�|��º � ���'��`�GP�S�nQ�#�J�z�'Ҝ\*׈��t�I�ςRi�	�'��y��C�-�t�ɑ�=\�&��	�'�n����&nJ�8�-�l���	�'�JI ���
�� �`M;Dt�'t�|���T���q0 Ht���'HF��с����g�[${>��j�'Wli�#"T�H��M
�I)�'j����F�<J����ڸo��Y�'U0 �!��Z���aZ�i3
,X�'�l@�4�D VH-bdL�9�zlJ�'��p�dh[�>��,d�- t5 �'�����H��>^>5s�8,
A��'�X�rCʔ�`�T��W�A�$�'�`�XS��D{\�BϚ��,p��'[h�1a+�� �
�Y��'�(HVfT
3�z���nF=�Z�s�'�`)��+	<j���*P#|�z@B�'%||!�a��B]���#ԍ`CF	�'&�=#W	7^mhI&�^�&D ���'�iS��L�^���aA�|�*�'?�R����J� u�4-������'�P�U뙪u7*y�`�R7f9�'=�����R�∁�n��(�"�'�����ϒ�5��8�[Л�'�@,I�O�N���Н.�m��'�X�
��M	B�v� r��Fm ��'�J4âm�c���a���Lz��	�'9���3 �����3 04s�'�F�!$��2e��T�q�R80qtl�
�'���fJ�2 �9��Ċ<��l�'�820FUQ�
x°m�b���'�*��s�֢z�"��Po��b�vaa�'��T�5���X����L �@�[�'!���`�@y"	j�o[{��)��'�J�����{��#��PW��#�!D�BbϏ1�4@�UD�k^�8i��3D�Xc��Y'cʰZ���5l �Qp�$D��bf�P�
m	R�-h�,�ô�-D���g֧S���0���� � �>D�@jV�.)�����Y*A��{�%)D�l !�K8+���rn��S/�)�U�<D�|q'���:�[t��	H������.D�h�'�²5M��t�@�1��-���+D�� �8XA�վN�.b��Ͻ���p�"O� j�m0G�X��END'�0���"O�Xp6bAl�l���������"O(� �)Η#C��#�3�$�5"O���%����˷b�6�pl�"ON��r�S�F�0=�E�ET�8%"O�1p6�'m���
D�?M<���"Ov�� Ę[4"a5ˊ CRB"O\083f��*����oH�a�D|1�"OX񢔨	�	eL ��%��2��iq0"OD�S���i7�EY���.k�P�A�"O��q&��}��Ԁ`����F\ѕ"OV���K]�,\<�6��q'��C�"O�ᰣ��)
�kDõ��̙a"O��a!PѲ���$V]ʠ��"O��R%�Qe��a�U)Y�3w"O�DJ���H�\�X��ѽ6�T�c"O��A�77t��G	�hxe"Op8��)�'R<CB-�7$��A"Oj�����c�ԡ1D���LM�"O<E���
�vx(q����f=""O�\��)P�H���ڿro�L��"O��ӧ�R��X���6LzA�!"O�}� �ev�AG pC�	�A"O�s��W�1�����%4�\�S"O�y��ӥ���'�� � PR"O0�+6%�O�.���0�F��"O��d�&*������w�&� �"O�ajQh�A�P�yǎ�vM�W"O�lT�P��>���Ǆ"h|���"Ou ���pT� *fƓqiN�(!"O��s �E�a�����$*`��Ku"O$�1#$�:k��:rj�< Q8蓗"O0��Ǡ>N���n�9>K���"O2%AC◨JF�,G��"MF�ap"O��s�B�h��<��N�t�T�Ȓ"O�q�@��O�8����ƿ,���#"Op���j*c����R�����"O�ݱ��ұ#y��&�&�L��""O:9RN zE�9�OE�!^�Xp�"Of�sb��h�I?AH4��0"O�{P�?�������%?-�$C�"O���eC
)'��� rڧ'ͻ6"O����N�8u`<!F'ٕQ%�d�"O|l[��c��I�.{>���"O�(�C��-d&��Nc�Q9�"O��#'�r�r �`�� ��d"O>w+X/��t{6H�4`���P!"OZ=�3�V�i�D@ae��:�6�3�"O���g�!����Qd�;v��I��"O�%I���%��ҵ ́#��*a!�$ʆT��
�} *�(p�Kh!�!�j(KFkPM�x`򫇣{M!��T)��H��-OJ�����NM!��>x�쑰Δ0&&�����!�Ĝ6w�[��'A����C�$�!���k�y�m8D�,e��*(a1!�_3�t��$8�~p)���s&!�dU�3I�u���9�x����Ӑ�!�$J�7���N	!��e����#A�!�^1Pz��	�2�݈��V+0!�$�+:�LY@��	�p�=��Q�2!���
����R�C��L*��V�h!򄀅� =���Z�t��I���I$P�!�� �ŀ���ҡZ�V�u�Tا"O:ő��ȨW>`Ȋt go<e��"O"Ѫ�]i����߻O}��9�"O���΀Do��9`��,�>�$"Ol|�oP���Ð��\0��"O���%��h*x��s �4���IE"O��*�J��I�,�B�ĉz�ڈ�'"O�E��!�R;�!B@,�x����"O<P�D;�Pp�-N��2�"O�Crj![��	����> �֩c�"O�M�q��2u��#ч�!Q��DI�"OH�2�F��
%D�;�eT��zX��"O�q3d���c��#s�.)[T"OZ�**א��`�,G&|C����"O�����[����KA=��=k�"O�T�Ў
����C��Ѓ5Ƹ��"O�u��C��^ Rm�hǑ@1�Q2"O^@��%�o.���%H��i���"O�����ݖx\(�,ݒ@:��`a"O�� �/ʀ����iS%$���"O  ����g�68C6���8��"O�����B�<a���w�Y9S����"O"����Qa%/?G�I�%"O(���)�dI�J0&2� S "O"����C���4TB*r!�`"O^��6.��W.Bq��՝E���i "O�%��F�Q��8�C[/OrZ)Z�"O��	v��EL	��Ť0ł81"O�ps�.�1'���6�
�j��c"Oj��1��T������܌]���"O�Ka�
@��AJ�E��˲"O ZA%K" 4`q�E]�Na�"OP"�@L�G�<�9SL؛o���%"O�f�I�ѡ@*�V��c"O.MqIÖ?J3G�
�N��"OT�h枦`��)Y��5h�H�Q"O$=`P�Kv)��t��+U. ���"O�`��@[�0m�����(Y����"O&���U��5
僗$FwN��D"Oi�F	��(��@���v_ ���"O����A������3R��D"Ot0���LB5v԰��G�eE��{�"OFp�e�Ԭ>�l��i�?�j�"ORP`�癔AMڍ �ЍW,��w"O.�Ы�D= r���4|��S"OZ0;CI	Xz\P����>$��Y"O�A�o�$j �8)���0#�B�"O�`���2&�]b5iWSl1�V"O�lRCLP0B ���BR�*��7"O�uЇ�Ʈ�z��U�o��"O"��c��<iZ�T
�R8���Z�"O�)��
�E�!$˯o�M�3"O1Z4P�W�2a�1)�7MBTu�"O]�D�������]�6y�t"O���%O<v���G�c�����"O���4��ƴ뱅V�M�E��"O�qy���>]z����Å>y\�c'"O B�M�J��� 'Z��"O\��eS��]���.i��"O�ʂ��>k���P�N�҂���"O(�CO�;�`����Q$-�|[0"O����	e�Y!D���lz$�`"O��p(�=���' �^�B�S�"O\t�<B~l�E3:�:�!�"O� �U���V:]S�$Ѧe��W�P� �"O����IƗ],�jU�ҾI���V"O�!�M�_�^�bH%4��a��"O�}�`	.��3p� - �)�"OndJ�ˈ�\�y$�Ǭ,	����"O^��"�U n���!�ֿ�,I��"O� c��[��@`邰F�N�w"O�S��˔f!���b�Ö��"O��XPA�H� P�"�́e�p��5"O��#��V� lN�"�K)iR.pR�"O�����\	m�L��W�רGؘ�"O�!y%�Ϡ%&�RҊ�N&T8�"O��D��"e�lj@[6_�AZQ"O\���)�0�3�!ԆX�����"O�U:
F"��Ig���
��R"O�����7����da�g�<%�"O�T� ��P����/�2�T=9�"O���̈́o�.9E�Q��D�i�"O�!�"e	R�����'Ā"O0� Ђ��K���x�����\�e�!�$��G0���`/նg*�ɚ2�09�!�иb�N���7@$�0���!�dW8>oR\�1&�#ʽ�&J���!��	C���w�D2x�Z�(!�!�D&�.�q�lQ����P��%�!������d���*�ft[�� �!��NA��xW.��s��`�H!��5,v䕩�N��y�d�0i�!�>=�"m 0.p���I�	$�!�DQ�m�>��nW�/sx4����h�!�Q�;������,��aÇE:o�!�ok*B�K+�j�3F�U !�D�D�����)=1��X[ƊNm�!�D�����zצ�O�f�c#J4�!�D�3{h�EH�/^��C�ƕBg!�$�=N�Du w�(Fc$�D�nP!�D¬h���t���M �3e�=@!�D����Da���*b�H�Qa
2A!�$��P��(m�:���j�@!�d��{x�(���#�<h���QG3!�Ė�L�|Mb�C׉^{e�l&!�d�
0�9u�gm �����
!�Ʈ#}��p �
Xh��`�D�!�$�������!�D��j��#�!�d�$l����2�ƃ/�x�ЊӲ-�!��Z_v��E)v۴]X�2w!�䙞Hd��C�ȓ=�l����&X!�dަ=I�J�K���, @�̋p�!�$�	I��ECAVE�&!� ��I!�P�^]6ܒ$
��P���-C �!�$��/+��p3�]�Lr�(����<�!��T3��4�a
b��`w�!�H;sԶe��*y��ۣN] i�!��@�E`(!#-��Uffm��D%yZ!��Q(��=��T�Y����l�lJ!�D�2_�ը��Z�.�rq��%O"4C!��iʅKg&^�f���;��C�94!�dX��(�D�%�8 8��	�2�!��(NA�<b�eP>=��B�\�!�dƤ��ᣤR�6Dܢ��W�T�!�$V�KD��"q|*] �k�0rF!��x*I3�f9��%#c��;s2!���RRI22�w�-R��"*"!�D�9�$���T~Ptr���'h!�� r,�$Ӗ^�@ :���@yf�÷"O�PbȌ(t��i%��K�h��a"O��R��'�� dU���r "O��x&C��|�������q�(�[�"OD0�Oֿ,WZ����6Fc.�b�"O.,�Z3����#��r����"OB�x ��\!0��qAD��~[�"O�Jq�آ.���q�-á��s"Oļ0a�!*B-�$�R-Z�U�"O�-k&�Av?�Q���5N��C"O����2���DO��03�%�"O\�[���nm6��d�L�z�:���"Of�HЯFKH$�P �3aqv��1"On���OI�{�@!#F��X��"Ov�u��p�֑ Ū̫,��x"O!p��E�FdD�2�I����[S"OR��嬝<R>���"��"O&�+銒|?�X)�K�7Y����"O愉�$=
6�{��%I��e��"O@�t�C��&h#eC�pޙ��"O�(�&N4�Rӧ푲Mk��#�"Ol�y�]#s�l�@PC<6&4B�"O��R�P7p��$;!�Ju5��v"O`гQ�L-���U	��9�aI�"Oz�Q#l��jDS�G��"�*I�6"O�tZd�dab��	tL��']R�!�D "��q�ĳyf@�qGM*J�!��w��ܢtK��S�� AR�:�!򤁁zV���+��U>��K�`Ԣ!��3<�42�}:�}�"��Ac!�D�^��'���;��y���S!�D�!Y4t�ycB�j�ր:�Q7& !�$�}�f�Pu�ҳa����J�1k!�$F�
���	p@��Z=bkEi�}!�؄'��a�nM�R4���e�!�䆓\��yB�Q�k�R�3���:&�!��{�p۵ჱd����CƴUM!򤄻R��	�Ư���@3b�3i!���վy`c�-8��5S�*�&%3!�$M$Y|�(t�؞i����ڻ3-!�$^�nު�r�3]~r���2!�$�*�rMc׋ɿS*P����1f�!�D��{��-1&�1yL��bFN"@!�dĵ9�8Y�L��20�����rE!�5a40�4��,��pH��!�ē�Dن�#`��v���#�!��	�A(�0b���1���D'xa!�$��?�aBs ȟ�����cNS!�X�_[@A�mCd
�I���3bV!�@	;�4X�W�|����U�&K!��).�:�hĬ�̔��M�I+!�䅀nPкv	޼��P���A4!�dG]=	��Q"xm[�P�>T!�d�N 5iD�̡�X2�.y�!�S��B���B -�~���!�D�5\p�!���+�"\�5�݊WX!��Z���Z��NޜZr���wG!�x���F�ҳ2ɾ5R��?_�!���#���ek�(D���Bu�.+�!�$]��avI��~nĚ�����'� @�NU�N�����)5N2\��'z^� ���u��j�b!��ȓz�$��líY�Qðe��-W�8�ȓ�5��܋�$L{f��cP�x��S�? |I��ΖGV�H��ׯ}�D�a"O.�x#"�2e:���"��)dp��"O�Q��䕙]F��+e�,�LB�"O��hT`�
��T#"wt�K3"O�uq�nc��Pp��/X�Z�"O���!}��� &o �"�"O�ly�śH����.A#v�:��"ORh�Č0$L�Kp���NXغ�"O� Ӷf�P⤜���ߑ&F����"OH�b�OK"8�G
X�R$�#�yR��L@�����D��8�����y���dX�C�ŀ4R�!��F���y�h �]�ʔ�$+�L�bv���yb#�8Q:؂���$���Fo�)�y���fΠ��e`�7 ���R2�)�y�IH�9�����Mٳc����O ��yB�KFl�ؘ�ꃇqg��C�?�y�*� Yd�\{	��@��ea"ꞿ�y�$�z[ܹ�ͅ;�`����ժ�yr._�4�~��P�O?/��-x6����y���O�⬁eQ�r?����D��y����E<�Hk�nB�p�5�4�M�y2gϢ2W� A˕�b�h��d�ޔ�yҊ�l?v���d�U�@h��E��y�C
	�T�3U�_�"X.]��ܜ�yRG�� �ȹ�p�����8����y���L����5�,a'�R��y�덒$���k�-X�ZPH�'N�yb��06PA�!�@ ���&˿�y����|g~iwcɔ��ѲV#��y��E�*0P��X+ ��l��DO0�yb����h$옎�%�ٜ2&��ȓ1m�q��<\�}R��]�B<T�ȓL�� D��"���ӱ��?�D4�ȓr�4��&�(c�)R��Zo�q�ȓ##(�	��@ jWYX�*߯|����m�X����R���'�6�)�ȓ,�,��G��Onř3�D�3&��ȓr�����cb�j�4�+B&���g��A�B� ZG�W#QN�)P�"OB�5틀WC���v����<��"O�#��߂������o8j�"OΉy�����ȊwP�z
L��"O:�8gf#9#��IAm�>[��4�0"O�]�fJ{��R%�С:��Xy"O֔�p��I/l�Y'f	X�@�H0"O�xɧ �t6н`Q�M #����"O�Ɂ�iQ�N��+F�Ӷ=侸Z�"O����+fx]�㈋$�豰�"O���d�==5�yX�a�k)�d�q"O|u�6(�5v�:���73�T��"O!�h�'b�zX1�%�-k���D"Ob�Q��lT�-�!ƞ���� "OB�"cE½W���1!Eǻ-����"O��.mŠ
R-L5@��F#�y2�b����!g�B-Б�&�$�y�BJ��RUO^/2;|�1�.ɗ�y�n�* �<�rb��-�<�!'���yR���)�Ű�CJ�wd`��_�yb��TO�sj��m���3���y�K@9N����*�Gx\���]��yrm�gf`,�/�Wo*�ӂ	��y��N1O4��A��1R˚}`�A��y"o�	O������_!{���h���y
� �`0B!sP���Y"?�@��$"OF:��Fm"L�6�R!#Ϣu�"O�;PԬl��ic#�&�x� ""O-:)�M�vE#�/�����"OL����DP�2���� ��8@T"ObAbG$X�Z�:"�.�A"O�UᑣBl�4s�L
��d��E"O�\P�n_�b� ��
Y){����"O�4(�%�u��1����Ow�9P�"O�Q�c ˓K��|0�'�fa��""O�2�iͳi��2�Fük�|��"O$�qs��+���+��/Z2��i"O��c��x��XIB��=9#0���"OV��ʚ�(� �&�F�;,0��"O�=�rŪDb�i`H�{_�H�"O~�`��{Xz%sW�z+-��"O�� �&�.:M�(���H$�kG"O�E9"�	)7��ip>���"O��xd��~��U3ץX�c^e�"O���!�[9Ly�$R3\8��"Obe9UBE�-B=�C�ّA��D9�"O~\��G�p��� �A�N��"O8��LZ�p#b��Җ}�����"O�8��Nl4`�0���W����4"O�$����o����LJGn��S�"O}�s�;`&�F%Z4TNε�"O���VO�E�bۧ䉣Gת|��"OnH2�L�&�! F(T��۠"OlE�[����;q�����+�yr�տ|t�`�5"�1�vZc�Q��y���e�\0�s�ՉS<�Q��_��y�#xڌ��)O�1�2��y����bC�,q�ve"J��y���j@G坁g�h�[� �,�y�.�j7����Y��5 T���y��؅\>��[��W�r0JVM>�y�؏>�i�@��
Q����ej���y2&�D5*EC���S-f�R��y��.�R��(� !X�@˔�y�u�dY'H	^V�����y2̈́�j&ht˧�9W~p�R2�y&��x7�,0�C�"{�i'&��yB�ȰGR�\�ӈ�^Ϣ���@��y��U6i�D)!-H�)�봀�yaG���d��*!�m���\(�y"��A���Q�S4���Pʈ��y���*HO8���̤�b����y���8$����m�{?�X 5#���y�D1\٤�!��ߝ���d���y�^�h�T0 ����Dp��M�9�y�F�Y줜P�.5�|� ��yB�"z��u(,ws���a���y��r��Ws�hPka���y"Zn��a�ÈqB8((!���y❼.��$*r-�kb*I�@����y�^"\����Qg$/�x��	L��yr�;*e�ʧ1Hh����yrn�g��M����$x���f�۲�yr�]�x*֭h��U1W���3��,�y�̑71�yX����X"�����PyBÊ;��5�r�޼F�e!B��q�<A�g۳9�|����Ҿp�U�Wj�<�Ѝ��D���BD 	�_��"!�Kd�<As��)D �E@��� F��I�C�y�<� U�EnƝV�F�i��oP�q�"O$H���i�T��U� �m���"OԠ#�!� �ӥS!��]K#"OR�2 &QA�nV/U�l�9T"O�҄������@5W\iA�"O&r���O�����8Q���kG"Ox,[R�2Y�:,�a����I�F"O�`�u ���SGBUk�j�s"O�C��� >5�zD�N�k��Lb&"O
��mH�{|�e��'&Q��"OLqHf˹E�81"Dӎ*�m�u"Oe)�a5�L:N~�x���"O����&Q_��:�j� %f��U"O�=(��Kz;Ă�� �$�d`�"O���FI�'=�<�Z7	�<g9����"O|Ayak��Rm.����֧)�}�"O��pMM>#�pDaF�����t"O�٠Ӥ�jպɡ�J�@'lu�"O����x9��K�M1�0`"OT{Ӕ\���M'l�q�"O�e���݄{FPYqF�H����P"O��ʴ����Τ`�Z��ͣ�"O�\�#��"iV�i�@Ҝ^��A�"O�P�2D�
԰��C�|����"O` 2q�:LP�p��ŏEj�	"O��bL ��eXr�������"OZ��0��q|��v
�
�d@+"O,� 0
̵+ތ@��K���p�"O��aץ �x�&�:�h����'"O���e)	 ꔡ�&�Q�$y
%"O���Å�p��D��掃#�� �"O�qz��K�[Ԑ4O���"O荓шX�,v�O|�Y w"O�W�ۻ|�,�Y0l�^v�� �"O�!j�EB�1@�e
�T���@"O�u��c�2m���A�)��I�
��"O6謨Xf(4K�샏6�T��1'�Y�<�5���~o8P4�Ge��P��W�<IQF�9;�����ʛT@ ���8T�lpwπ���h�%�M�:��$D�Zd	�t���Scѯ7oF���!D� ��+׿[q��@�(��2(y f#D�t��o��t��=��i3.�9��!D�РqJ�9&q֡���"w/fA�Pd4D��W�� �
�k��I1}@����0D�Y���${�i��D/��Y��*D��a��(�rè�ƙK N%D� ��ģX\��j
��|����.D�����~B�\</�HU���,D��(mߪs^�[�W2?���rpg*D�@��ĚxL`��C���t:�C(D��'ƕ*L��(�RCU3iP��&.1D�|�.�#|�1�C���h@�2D����k�{&�����
���IVd0D��J�N�x�Ε u��
AC��0�(D��2g��?j"4i6��P�|U w�(D�@���$M��Hk!ZdZ�!&D�����M�b΅��O�4o��E#7D����Vl�~P�� |��H��i4D��J֊�3_L����ˎ�I4���c�0D��H�_�PS��%��E"I1D����ƭ2��87���	��Mz+*D��P�F��2�I!"v���*D� A�[^����-]�$�䱑 *D�� ��Bc�%��Q��G�"X$��"OV����C��P<�4�EQ��u"O��z���G�L(�\�J��Y�$"O6���-M(y���@5nM�p�a�u"O�Yƥ��{���ق�//f���u"OqB�@�P�|�Cv��,N���"OzeqSj�&���C��Цt�� R�"Ol�A6�C��0�[��[3W�
AQ�"O��9��z�8]��݉Di�0�"O��s4�L�H��]�X�2�"O�@XV�q��Y!1��$�e�2"On��疔�Dm
������$@�"O:����.(};�� d��b�"O|���/�7Oh�2��)[q,`0�"O�=	F�<>{��P���K�03�"O��!dG 9;R�gCBR<�K�"O���0����0�u�@�x<���"O쌸�e�1��BhQ�5�q�!"O<	�-P�0@R�+4H6>1*!Q"O�x�	�l}nޜDcB<�W�2D�|ٴe��E��L�e�΢|B�P�O2D�@q�*���H&�˸_�x@p&m/D��kqh͓L��Ы����/m0�a�*D��wK$
�԰��"Z�nР@�)D���g��#y�!����P�0����1D�ԓc�,|�A`��/Ta+�F2D��`a�Fu@�y�"�3(�`�Q��3D�����
kπ�	t%��4`Y$m3D��'�.�l�˙/;���Y �3D��`gC$�~��3��q�j A1D�I�5>��x�rB� baH�j.D���b)q�`�GMڛ_0�U;�>D���[[f��pE��W��-;D�D��"Ĩ%�ԔkAa=%���f�9D�dX0�}������PmF��L;D����$V���Q��A3K�j��3/?D�`�V��)���q,�#};�lc��9D�p
�g:l�A�_>0^�T&3D��D`�a�x�"�NX�M`J��� 1D�<�#ͦk�p����#�.���/D��h�훩W�d�f@,p\��{��+D��Q@�Z�9�����޶���,D�������$�h�Sƛ�e�I�1i%D�T§���o������*��b�j$D��:E�	��P�2���MQ�	)5� D�0�0G�45c�HP'��  F��F�0D���e 2cl>`R��ܸ+
���,D��� ˢ|}��It�T��H��E*D�@�n��F�%�,�FL�	e�(D�\���[�����E�E:9 �*S+:D�`��FХ'z�5J�@�z���5�6D�@��쇩i���g��x�p��w`6D��&��$J!6,97��1X\�ӡ�5D�\��ON}&f	�6�\7*V8e��'5D�hH��(� =Q��l�@���(D����!�Gp���7��%T�t=��('D���㟃5fx��D�+O����I1D������XI�1󆝤m+H!�Wd.D����'�@-xZ4�Y
y V0�g"-D�T� hؠ ���Y5�ݛmG�R¯?D�I�ҟ$#�����/�T!��*D�Xف��2z��av�s6�R�2D��*sf�<c��*�O� 1� #D�Ȃ���@��� �,�J���C�*?D�� ����ݽ)j}YTJ�u\���4"O@�Xl��Q�8���B�l>�P��"O~u�cA.|l��;gB%|0��2"O�a�f���R+�
|�Ћ�"O|�B���"r�98�*@�s�B��"Ozm��`0�AҒN��1ʦ"OXEz�a >j�� z"%]s���6"Ob5W��9ov��箍;qXlR"O����e�3������8]rQ�4"O~�2�I�k��) ,�;:T ِ"O�t�v"��ŰDi�%E�V")�d"OL8&�8:s���vZ�9EҤc"OpUA��GX�Be�n��f�d�d"O�x���1	$�a�g]�-&,tP"O�T���Ծ�>4@��PKb ��"O�D��%W�M�rL��-k���"O8��
1���E�7.>]�R"O
�#*���%Q1˒"t�h"O��r�KyFQ�`�-���"O�I"ˋ�Q\|c��%\<�ȱ"O����#lEЀs1��%����"O�4I��~W�ٗR�5�p�2b"Oܠj�,@)Zx�ˤ��R��8@�"O\,I7@�8<ۊ����/�p�٥"O`�bFC�Q�Z,K�YC�!�q"O���GLF�귅Z�%�pH�"O�c�+�7�aDC�9j��Y�"O"��3�ѓFr�Tr`�?>�h�e"O�� $ʏ�CNiS%�$>�Jq�"O�@귫��cIԵZ��n��Ը�"O��Csj\"�@���H!��M+3"Od}H�O�<Ug }	5�Z��~m�U"On-W��/`~�"�P4aƚ,�d"O��w�=[�䒳H@,��[�"Ott�"�
�0�����åV���2"OX	�F)ŠF���$��LK�u��"O|�R�)ߟ*T��@*/��8ct"O�!@��G�o������8.���v"O�9P�GR� ��y`�^�4q�"O8	��L�D%��_
Q�mp�"O
:�"8Dޜ��#ܢm���"OD%*�)S X8x���P�7Pu�@"Oԁ!�G��>M�ѤB!��p�"O��D��y��#Qc��8��u"O޹ ��QAB��A�!|��P`"O<�;aKD� ff�	�b�G`Eb@"O���׋@�a��Ç"�4+4Ja��"ON���!A
�}��<r.b q"O����ʤ)0���# < "O��+�j�	��X
-�	����"O����+� ����L_"#��U�D"O�|Q1�T%,�X�Q�\\jvUs�"O���!�S�GA���H���V}�C�IN�~��$�A���5��*@vC�I,a�f�c��?���@q��D�C�I�5p��a�b��g��+:�PB�I�~�^d�sN�-U.�����W��B�ɒA��i�M�0y�4�����VB�I�pDY"�D� �.�Ұ`_D��B�	�Z������>w<,!q�(��'�B�l��J�=g��Ȁ��XX�B�I�I�� `e�Q�h�ؔ�Fƕh�dB��(�fH0s):Xu�`��ƅ�(��B�	w��6%�;�j��soŢQw^B�)� .�c�bY��
4�"�|��m��"O��;��!|M�����|�Q�"O�th��ġM��2��\�����b"O�m�r(�4d;(���~)�p"O
��4�`��9S��Ge���"O��4���Y���@L4)hŐ�"O�8xc�I&Ll�E�%�V>b��8�"O�ă3�ިRx.�PR[^# �q "O԰*bk�;/�p-q�K Lpe"OF� 2�'��T35���4�(9kF"O>�q�B6hk�0�b���L�@�"O�g -+�����ɳ_��$k0"O��AG�Pu���@G8}�Y��"O�m���N$Q4�`��S� a�"O.�j�A�@�B���ԿQ���7"O8Qpt���Y����aE�<[2�:�"O���G��.6\�$$@8*P���""O�4F P�tNܠ�����<7d�"O��JQ��7k`A�G��~� ��"O�K�̑�Nϰ��cE�n��X��"O�<	@���ˮu��a�@�Z|	�"O(��r���~Qs�@ZF��UP�"O,��C�ד�ޅ�UO;,W��"O����n�8i�X
�N��
#��x�"O����ńgi:-��M�+s0�ja"O�-��(ј}2�٨��h�Ȋ�"Oin�x��ez L����RE"O�@+S�����(X��ͣw:���"O̰:�jG� �.�c�6�
 �"Oj-C��#���!C@J�H�"Orq��D8�4�P'G�欰%"O(�r����6�!��Q�G�nl�%"O�A�H� PQ�#Y�����'"O���R$�4g�H���M�=��IH�"O�(9ԣƪnE�Uy��	�[�"O9)�&ƱX��a�m_�S�j!�F"Oz�ZEG.-=���l�̂�k"O���EZ%0�ҋ��"8z!"O(h����
9�LrF�
0%�ּЦ"O�uH֋��{��IzH.���@�"O��+���6&Vq`
F� �lH"O��{)�b�������)� Ӷ"O�@��もG��0����#0��9J4"O�p����6 xj���x|2<��"O�5s��J�`�i�u-�d��q"O�KC��.9x��ۨ3Fb�J�"Od��D��DvRa�%����t"O�Y���ܻTQA�����	6"O8d��aR�h��-��E��!U"O������p��ؐ+�[�fM�W"OxaA�9@�� �ԫ�>n�Ա"O�b�(A
(�5��
�A
��"O���խ�2[�Mb���|��H8�"O�����I<�0�` J�-X��a�@"O���!���k��h��/L�vy�@�c"O�e�/
m"q��ݷ:X*)z�"O����;`��B�Aat|�;Q"O2H+�jŖ	qLHzqLY�j���"O"�@֌�:}����J�i�,�a'"O|T!%	l��MӲfԄ����,D�l �/ȍ"1�ĠnY����>D�КA�$3,�3��B�]�U�@�(D��3�f�'�P�8��E�9cO(D�$���e��D��4AQ�1"ad(D�� X�1�_ [�,��ѫ��L� X��"O�]X� 7�~0MM�M���"OfE���-]��}@�����Q��"OBAr�,��9�2�ݦĄ�3�"O�i�b��8X�p�-~S�Y��"OB}r�)
������¯n���@"O&��5k
��租�Wy�P��"OX���f�P�΍�c�9r9jf"OP�׉L��0��3	ه(0�(�"O8-QC˝�B��T����u�>�i"OV�E��|[���H��0@�q"O��XgđWR��p��S�M���HS"O���"�y3nDI�J��/N�ܻ"O�-�FF��Y��࣯�3+����"O*��Łՠ� �{�gX�a0(���"O����^=x�JYд]-a��"O�UQ'l���b�d��dl	�A"OL�A�-�9�:��4$+X�F�0"OčRàE��^U1���:t����"O�I�f�
r�J��EA��߮���"O����i�X��E/�)!�8�"OR�+��"kVD�!.�?89��R"O���C{R\��E I�Y u"O�8� 1X�.��R�Of��"O�ɤ��<]�x�q�M�=UhT��"O���!B�0I�A�| �q*S�y�R�B-p�PT3]*��0a���y2���q-ʕ����P�\YR�3�y�ᔏZ�saB��Q%ڴv��y��D�B�������\}�"�'*H�1`�<g��0�5EViq�'[(��@J�yj�Ё֟'r���'�ne�ŊZDBP�#u��%~��'��-*�\
�m0��M+$r�8�
�'1�D�� P�s��ӧ(ǣg� ���'��=�D �]����f�I���'��m�Ee��hI*=	F��Jrڑ0�'/ ܻ�F�-�f9�r0�LC?�C�I>�<���Fs�~p�4ˀY�B�I�+y<�"�G�/�<|�	��h�C�	B[j��G�Y�V5T@ƁAA�B�I��d����9�1ٗE}/"B�ɂ5Pf��7IXӖ���ոX��B�	7&t�yq2I��� ��g��H��C�	�eFe��
E�&�m��Q�B�C��X]Hm���,"z���"R���B�ɏW��P�$,ӳ��z"��K �B�6w5Hu ���7 ?8I2q� �2k�C�I�l<�Xbn�����(3h�#C&ZB� /� 0��E���p�ƀsFhC�I�D�RL`�,X��) =s�ZC�g��Y@Bf	�/��#/�~�C�	XT�nS�cΚ@��0R��B�	6S�-�$m��`?�%���)/��B�I5$�p3��0xR�=���ǹ8�BC�ɟȖ%ړ��4�إ4�Ʒs"C�3U�5A%�. ��`E��1H�B�I/`3�	��L�'u���	8Wd�B�5<HԌӆ��+p�Tl:2$½K��B�I�R�Qf����"t�ҩ���B�ɗLm�p�
)g�Q�S�5s%pB�I�Tن��$ll��s@�� B�ɔ*��ª�3�! Ը3��C�I�jd&X� E�:�V=[��S�FW�C�)� ��k���1cO�|4\�JW"ON�5G�����F�(�#"O��3��[=pI��z��BBЍAp"O��'I���Li��)a#��;�"O��A��*FH)I�
#���"Oli� L.C���S EB���"O��
`G,.`P�w�V�<��D"O̅�6���j�T��s(�;Ҧ)�#"O�LѶ`���쨥����b�"O��1bY
?�����D.'�ґ�D"OحJ���^G�� uE�'T�zH�a"O~y9F�D��փ�%X�
墠"OP���*\�H$:�cȈl���"O8�8�"�$c���ĔAb��"O ���+*� �C��eS`}��"O�(�d^�m�|$�3HDu7�H�"Op��� �:���U.����*O����Z� �hJ4��v��'�f��&A�] Z�!����ʉ�
�'�|�b�Dnz�`�"/I�~��	�'���RB�p�2ݠ�ʶ{�PP	�'�z�H�h
0>�ұ$�*v�l��	�'����g3-�j����g�Zq"�'O"���ޚI|l��Ы��[�-��'
��� ݵ�vL� A�U<%3�'���8W�w ��@�,�wu��k	�'���v�^�m��婅d�h�	��'��T<Bz�h�D��J+ܝ!�'�����ΌS�}�amΤo����'���z@���:"�u��4aFj�a	�'����a	�1��U̅�[����'՜�I懚L� �l�-[Jn,��'\�ܡो�X7����*LEd���'x*y���+�*Fˋ�{�̍�
�'n��Z���&sn]��	�m"��	�'i���*Ui`Dȡ��)V>E��'�x���f[�a�v�0�c��?��!�
�'��8�iH�H@5i��0����'m���f�0�pi��*̌-�r�'�t�X�p#�uc� �nl.P��'D(\�� �=[�\V�i��� �'�����2���hfkL2Xe����':�2"..X�vlїLv�q�'ʢ���$r���(@(��GI���
�'�A�䇖�`�� fǺ9��=a
�'RP��� '.j��^�.R�Y
�'�Z�HǮY!d����M�,��X�
�'k�x�̉
?��5Ȧ�̤$#��A�'��Hة/� �[����ZBd��'p�fa�����''R5 7�՛�'�\e�3��`e�l!G�
gH�D��'BZ���`ɏ]Y����K^�d<���'.���X}�mh�%Nb�"�K
�'�:A�5E�Ta�ӞV���	�'̚!hA�l|u$��$+b���'`ڴ�5G@�U�$u���S#�<���'ʰ�S�. ��b6�W/�l�8
�'�Dl2&�`\+�	S�!�D\X�<��!��B��cT)�?��\Y���}�<�*�}:�aƆ��y��� �v�<��ꟶ*d4m���:�
Qs�s�<s��F�������� #������r�<�F�r��@���$e<��A�v�<��i�<6;Xm��-�$	 d���M�<� 0YlR.H��ܻP��&�|:V"Oд6C[�/K��ا,�*�,�G"O�ieLㄋ�Wf���"O�U����5nC��� �H� (["O���Rɐl�\8�I�.߾գ	�'�4P��G�8�`Ek'��X	�'�
�ȇM�:qF����O������'����M�!T���r.S����'����шr���)b�Э-�Ĝ��' ���aa��HfE˱:Μ�R�'�8��Ve��dղq�ڿ �ꙉ
�'��H��e�A%~d�ʊ�)�R,h�'vH!AV�7e����� �e��	�'	P���fĬi�dƆH��]B�'���V�����\�E�\�{�',�[p��&l��;ӆ��7y����'�lY;��R�jl��(�.�(�'l �k�!��&�ԣu��V�а3�'OT�� K(l�v��$��q�ī�'��8�7��t�:DkA�%E\��'In�)��t�D��p�Yd��3�'���s3M]��d�7�Kr�X�'��`�&@�#�T$V=Rh��'�� "�Ǩvd�ڳ��5Ӭ�"�'� �"Q�V��H���/rh���'0�� ��2$Drq@�	�8�C
�'���1���J~��e@Z(YpeX	�')�%�vmF�3Q|���o�}��'��d���BX�䬍��&(�al�b�<�5�B�M����K��.=�.s�<#l�K�:5 �+�em,;s'r�<Q�Uh��J	7/�H ���KH�<	�߻"�j�c�AL>v����\�<I!�)zS�A��(K�> �;���X�<�TMԔ��l@c� N��T�NS�<�� ¡%��� saZ1�b���e�<�����M��S�,D�q�x0��m�X�<�`@%i9��2��!qHԘ3S�^�<)B�	�$������U�{�b���W�<���5~�1�МY�������Q�<��㌄L��Q@c�^��T3�EBY�<�W��x�[�P�0�ZȚvNa�<�b^�8��̂`�R��1�Մ�Y�<񔂉�$p@�!�Y��%R�<��h�m jV�Y�ؔ1�a�5�!�d_�C���w��iݢ�c�ɲ)�!�DjK�T��Q���'n(b�[�!���΄2��z1�,��Eۢ7�!��×:
�d�2�W�g0b@+�Z-H"!�$ m�(̚��ɓA,�dP��L�!�#�0ai3�U�:{�ũq���Lv!��Q���q�!O	
�D��cҌt!����@d{�KĔ!�J��6o�!�~t��d�F��#7�/l!�D��:�|��� �I�
�![�wa!򤟨J1~b�\�0�x�H��՛0�!��L9N$����ňM� �f�(N!�ɍ4W��*@��T��(��)Y�t;!��� #��r��)mw�� �gP�,K!���9�Pp�A@<ZV,�镥�);!�D�4�$�i�/�\9Xã�<%.!�䇨o��(G�%}H|�c�"�$l,!���_�T�@���j>D`�C�Ǆr!�ɰ{�a�ʐ?&���M�j!�� ���P��	p� �m0(�2e"O��Je놏mp$�p֎��.x�A"O�ka�0I{`|��g��L)H�"O��:��� jP��b�^�Z��J�"O�x�
��3��ʱ�	;�L[�"O��#WF��5ѳ��3R)S"Ot9�!Z�^@쌻w"�;!.P�{s"O%�Q �"�d!���F�d�� 3�"O�kE�M���H�*ȗmL$�:w"O%B�fR�<�P+w�Z�+�@�"O��@R
�� ���*��Ӽ�x�"OPL�4�O�7%%JK�V�P@�0"O�k6拜J�����@���"O,���Y��� 1R����A"OtԐ2�B�~�V�� �?i<�!�"O������]�pD�!�V�#nD( "O�)���(p���2G��v�Υp�"Of�C���`�C�"qxw"O�ԸB`
�f.���P�&Q d�"O��SJ��I4������7"O����o�Ϩ�H3A��"���z5"O ��/*B�F�9֯�&\����$"OB��`NK�K'�S�!��aO^��3"O�XSe�Q�J���M�B*P�"O̹�P��GU������ghՃ"Ot�0��D� ��r��8a��"O@Q	%�ؔe^e�ۮ/���%"O�Q��O�R)X�ʿv�x��"O�l������-��ZM[�<�4"O$�FϦV�$I8��V�M���"O��YTj���-���������"Od�����ei2MX�o�D"Ol�bA�C'<�鬘�����Nl�<9�kS83�"�T/N&
h�KQ�<q���'icF\�%�� j����b�_b�<�4-A�I�&�{r&E	 A[�<y�������B������U�#>!�$�6����+8NU6�H"f�2y8!�Ď%z�L"UJID�m[��Q4!��M�w
zpD�I�K�l`�����,�!��O��2ԍ�����褢�%w!򤞒 �dl���$>�X��T�%zi!��׷C��WEC�b� @g���Y!�Đ+T{�ɢ�J>J
BdKr�۔�PybJ�"^K(T3�'�<z5��0	ƿ�yRǄ6��=;7$K�vL��ᜎ�y�A\��a���L6�����מ�y��T�H'�#�f\~�`�:	4�yZ�E��'XZ�b��'�,!��4p�'Ѭ=ɕiU"A�I�0lӰ`U�
�'�tи�!�b'Be���o
dH
�'�x����:[j֥��lp���	�'G@�Q"�Fn��v��8�@��'&�YƧ͖:r���Sa��a�'eHxQh�K��I�$gH$_*´��'���S#��x�����.Z&��
�'M��1��
C�B��@�e
1
�'�ژ*���sD�q��@���k	�'!$Qq�M�?oI� ��3�:ݛ�'��XRD�ҏG>2�����	�'��u1�]�v�2�w�����[�'��E���~��p2�lвrJ�9��'èh�F�Rw9����jX$�!
�' �b�'�{�t%#1H
�7�bً��� >ū��0_&Bp�G:&j��Z�"O��zŊ�W��ys��
?9�h�"O&@�gǋf�!P�d6|%�z"O�51B�Y�2䈍�2� Px�9D�DQ-�Ar�D9�+.��J��;D�$1c�ʄXH%I�)��jU����:D����!A�8����Ҕ�M��3D�Ȱ�Bb
 ���R��,#%C/D�H���֕v�p I�Ȕ~ٌ�c&m"D�$��膲lP �!��ŃI�0���?D��'L�(M[�Nª��r&�;D�p)BBL&�0��߸�{��:D�X(��_����B U o9t�4D����+�7X{<�S�$=5�� b3D���C��
}��!�J�Cԝڔ�0D��hsa��������
��-r�-2D�|j�G/:�H��օAmP�Q�h+D�$���˚)dnL� j�N���)D���CDi���7m�!i���B7L(D��Ҷ
��%�䐸!O�vr���!$4D�\���\&B���حkb�-D�4A'i�P1HX�t��Hs�u��H,D�(���֡j���J��\�^|d�	&5D��0�dj-*��6��7t��Da�0D��x'f�9l�&)�sh�:*B`�"u�.D�d9D�]���B�h�byb,�J,D��@�U�z?��:VH[w
��0�'D���2j��nwf���H�:S��y���<!��哈o̥�p$ϜR<pe�#J٧�hB䉫�8a3v�W1)�Lmit�ԩXA0B�I�F�����T;[��	K�d��y>�C�	�"�p26#
�gøII�M]�?�C�I�?AJ����hVZE(�n�/S����?����%ڗ�f2n��$[Z�xV��y��8ܸe��C^�~�u��(T��y�&Q:�b1��%�0`F��fA.�yҊ^
l:=��.���*��I��y�ș,���# �d�4�p��O�y�!��1t8$�g� s 䝩�B-�yZ�N�iG�͊X�r-��L�m�2C�	 JH�IS���G�lUh��	��B�S�t��rCA�^�P�AG�ܸE�B�(�n��A�v�D����B�zB��h��0����]ܱ�SF�j�\B�	$Wt�S�/V?a٢�ҷI�B&���f���Gb�?t��4��D�=Δ���+D�����?*T��U�ŧ2HlQ��@5D��qEM�KZ,��ˁ?#`U:Fl6D��h7��&a�z���M�(�:�y�2D�L��C�+RQ��`0b !j�n�)r�5D�p �ޓ���p(�$J�^L��C2D�yP�� {�Xhd

���Q�1O�=Qt䍄{��Ta�ǒF��Ё ͊\���=�p-AM�r� �)T�ɵ�W�<��O� � )`�
S�������J�<�g�(W�llsEї��)�1��l�<��F�c]4(p'��;<feB�i�<!��E����&��zw����_e�<Q׉�G����&�H����%��^�'NG�D&� �4K#��/h��-�W�C���Q�F��d��j�l�5O:���(H�`�O^�=%>��GY�Rt�%h��.xkԍ*D���u�ӱf�8|�� �m�`lz厵�زe�>�&�5�g}�`
�l��b2�=�"�`�B�:�y
� ����Q��;gA�#�L�cqȏr�������B9rlaB��*����y��_�M��㵋U
���E�W��y��C�?�	�h�gX�s�J�y��c}
�9���&؁x����y2�Hx4���Q�*� ��y�cR�}�b����U>s��pUmY0�y"m�e5���$�ע4~��	�y"UcU�ԇ��9��A���y��ζtØLP��r.m����yBc�.fi�v��z�J��  H��yb
�->����r�~�3��
�yB��Z�Г�b۷}����ݵ�y�؁m����͕#z_>��f�>�y#-%^�P�p��3p�8AT	�y�N�m=J�AÃĸTi�"�K
�y��N���A��)�`�'�W�y��W�>s�U��`	$F����P �y��F�����hOɉw�U��y[1[|N��q/0e\�C���y"m�1(�)2��Uyk.<�Ҁʤ�y��M�6���!p��*��y���yb��r�<<��
ri"Q�[��yO��JM�j��"|A˰ Ƹ�y��N50|��V�|"��g����yrÀ�:t���q-��|�V����R��y�ΓC���6�\ ��$��.�$��ȓ:ĪiP�!BG{J\Pd��襆�[�,� �D!E%���&�\8���gS\8K� R�4(*�����u�y��oA p"��vY��R�D�z74��,r>�P�h�
(N��p�?���ȓK?���r�ȅ`h��ò��;à�����5���lo�T���7�(�ȓ))X�@�&�lQ����ͅ�(-�ɒu��W� ��sFbOjx��Ql�M�F��5^�@�s��}����ȓ#d]!eh�d�j%���G7;kJ)��ph�� G�[��]9QE�	N�=�ȓMA�}��nT"]��S� I�ȓ���aԯ)|�a�b�K�I������d��-+l� +�5l^�0�ȓB��ن��PH�\B�֚p�@�ȓ<���K!�?)�l�#e�"�ȓ4������*�(Cv₼OflB�Ic���u��\z$E�ר�sR�C�}|F��~����,%jB�ɺQ�*l2�Az�� J���/dB��H��9Af����C	DZ�+"O��;$M�3O�B8�3.�&Rl5*�"O�Y7">�nD�FnY���i*"O�y�Ё�<m)~�8���y��-�"O0 A�f���͹����� "O�� �j�J&������-g�ޤhv"O걇�T� �@�E�.9r�c�"OvE�'E�B��}���t9��	�"OT�K 	 ��$qgnę"%��V"O2�+	"�����ߘ=��pE"O�D���5�x���l�Pp���"O&�s"c��q�t��^��Œ�"O�� ��� �8jR��P+�ib"O�u!��ȅ7~>l;��K.(t�T"O��b�!�~��	Z0 ��5�$"O�=��ʜ4Yd u���F��pi��"O� |��@Xsv���g��B���a�"O���i�n�
����I�yL,3e"O��p����o.ΌH�
�D
F�"O�Dq��߫#�v�ق,ӆ>K��)�"O� �E���D���ڒ�44�+�"Oڴ�4��-Q�"`3�)0��%"O�}���֝a�B�&�[H�1��"O��{1͋�S �0�e�'\A�0��"O���CH���`䋚8%f��f"O��{"m�X�8p�T���Q"O�+`�J$8�R�"L����qp"OĹ Яٓ�����B�����y�"OH�xRcJ:+�4X1�R�����"O��!ef	�-$ UӲ�@5^�B��"OJ���5� )��+�3᪐�"O6������ �x���6�"���y�$Ӥ#�J� ��C�'�*d��N��y�a�.
|�*��G�pBu��y"��	(ly(��U�)_���^��yr���YC.�2��� |���2MA��y��#W�6@ GB��ˎܢrcё�yҭٟY`f��/� oRJ�
2����y�(�6�>�	��R�o٪�a$\��y����ܡ�aN��OZ��.�y��2s���2���o�*P9�ꄷ�y�N4H��΀aјL�t�]��yR͡���j�aPaGrX۔��9�yR� /Z"T����UY�����y�A#_D|���J�$.<t��J���y�e� �X��錅i��÷)�y�Ȋ2?����oN;a��9�Eð�y��O*��zf�Z\�uy�j���y�� ��U��X�Pa����y"�ڇS%�({��4bx�m�3�C�yb�U���2�lN9^R����ս�yb��[�>q�'ƄDf輪$��y�dk]�X8��
�B݀q[
���yR >mZ�
%�A8j�2���F�y��͕"���Rc�Зg�@�r@Ǐ"�yr�Ё��1Au��$/���Dd��yR�N�F4٠��X�0�k��y���-]�H�k���I���H��y� �-ǔl���::��%�yR����}��'8�P1+��Z�yRaJ(Nv��E`%.�S�7�yb��0>.䑰ρ;� �ʁ�L:�y(Q P�G.�N��!�ظ�yb'S
E@D́�By���"�y�KV+�,�{��ӕ�((�u���yb���d�*�ꆃn�Y�hˮ�y¨G-U�p�v�Q�\���O���Oi��"�wCe��L��Ȁp"ODH�ըIq)��	G��i��)�7"O�u)s��l�N�k�Ku�l��"OPP��ӢU�����\5C� U�"O�y�Ň0j=2S-]#X�`$�G"O��)p�4#>��u��2�b(��"O�*�#������ѢT��<��"O��銖Gd�i�׊�usN���"O�,���M'a�2�	�����&"O ����A,�&���N�"O��s�ǅPZԠ"��3�8�ە"O�Z@�ÕC�6�"��w$��3�"O�L��	�k����Fh=�	�"O��Xqd��Ae~�@���r�z!h1"O� ��P�nȆH (B̓�bǐ]�"Ond�6F˒/��y`�c��yQ"Oh1�B�eךD;S�	��D��!"OPM���E9c�zDqC	�k�z��"O$�"#K�z(�p胫���h�"O�U� N�
XH@�����T�f"O�����M��9�NF�	ވ�k&"O,��&��3<�[�(��5�И!e"O�:kL����ĢE'�袕�RB�<�5��_b)�����C��hB��x�<�Va!�h�Je'Ղ
�݉��w�<aUd�j���"u/�w�����VX�<�ⅉ*'|t�1�9Cl\	e.�O�<!���$����E^�{�.q�b`I�<��	p�(�0i�3ZF앋q��s�<! B�	� 9��(;��m���y�G�/\D��/;�&���ύ�y2�^a(�����L9�q*��J3Rh�5��/N��(��<E���:��M���Ԫ,c<\����-�!��B?��+��Ae��E���_%����I:r��IV����] �X�(�(�n�|3&B9S,�S��1lOF 0G�"{�6(r֥��Jhz���2ţT VG�M�Ė ��?�'NE:����� 4ݦ<���Le�nQ�B0&R�s/�9�@�^���N|WnWu(��#������R�Yg�<����6L0~�#��I~@�Ѡ\�|�d#׾2�@I��dǄ:F�tG�b?�����xd�VU�F�
��^h<遫Ę9~B�s��T8<�D�cM��J����<4,B9����?�>1�����O�)�re�w@`hR5C�$Lv�] ��'�����ƧJ����p$�&U�X�V��w�=�1i����D�E��|��I�O���d߮@��hq�I-I�:U��f�3\�'�y��/M�d��̛�)Ɯ=�EIQ�H�ܨ�O�z�M

Xlȹ0@ǬH���'�Z�SÆ�$E8J�d�%F<�#L�91e��¤B� B��pZ�$�c�%�IZ$E(ӛw�P��ѭf��Eh�+��$
ԙ!�')N�pC��F{���S�]Y��3D�7�<hI$ǟ9��M�1��9K��QHC�Es��H���ӹޡaď2-��=�V�*O``�&��ϤzWě.�b���V�$�����'��|(��#�n�Y5�B+@	��+F���p�K'd�c ��:J�'ʨ9
��F4x2`�(���jI��[�a	nD�����|ʳeC�je�� (�6<|q�ԡ�@�<1�&���ł'�����c���8d漋�J�~_���Q�
�'�ȹkp��9����7�\=���K�m���1�
�1A�![�kt6<e�0�Bzx�`����p�P�������(R��R𪐀\-�M� ߼vxq
�W�[ ����� (��K�'Ч-rO����ߍ;�v��Gm��&�)��ɲ.��Ӱlߌ9�|��7m̨#��R��3	ĤC9�08��O>@`�`��47��/z���!3|���i�z�����-:�����ú
�x�ȇ�M-�ȊӮ���0��@5o�f��TB/?� �˱L;	�l�f���'���$ո��Żv��`I؏��?Q��x	��a�@	���@��!�j��g@�2#�� @��'�r��� 6
��X�jϱ��!�;)�Ҥ���E3��A�@�6x� ��	u
�y��k-�¸���/�,�2�AB�$+�m�˦�ृ�_(0���`-�AA#��\<6�	p偀 ���b�>��J&/�"�Q�J� ��ikF�A�lΠ���r&QA��N#V,ba�ڱ/��Q�eҢw��"��`���-#�\*� 
�0j<@���{ip�.:*�G~����mJ��e��B���:�` '�a�P���W��`���Pd)��	g^��@e]�A��5@��#�Q��#�tЪ���_�b?�@�,A2<�i7�ZL��0JD�Z�4�iprE�fΐ]����"GM��)�͐�&U\P16��l��D[0�
i`�eaĄy��Ip�����}��@X��&��i:���԰=i�D��N/FY�GJ�&����0$޹�-Xc#L�l�����O�N��3QH��75�D���
y���`�^8��#M�h����'��á̗�O��݃ i|	�pM[�B H�C�Ѹg6��C�1x*��a�:k�#�c;�xa��)S�O�ڴ#�D.�t��W�~�&	��N�8d���x������O>9��"�5羈RQ��/ְ�;�dӲz#�9�.�+�|�2�ۺI2!���6ᴜr��,ޤ�S $�0 P�XĂ΂w-���̙�$od� �C�	F)� p�[��rMˋ_S �b�c\��2��n)Դ����ì"5�Q��(C�_�$���J�_Q:�""#�Ղ�C�3RD�����I��Ć,�����F&`�a{�ŗ^���\�����(�o��06J[-�t`B1CҳP����V��d��ͨ��&2*9�+Z	l��v��/�~tbq�3�~��4+� �i��{�)��h����'9���h��lBz�$S�!�hJ�#�?��ɢVa�ոmJ�@ACJqɓ���wx���ڷO,�h�(�++p"H����O� ����0I�`2BAK�b�A�$(�]AD$'���`EO���ޔ1K�h:R�� n�Td�*ze��i׉"�ؼ���٤�h��c��r���� K����&�?!�M�&�Z�t�p��o�zg��S"Xnt�%sW�H����7f�>#�U��4d�B�̻A�yt��iV���O[9U�|��}�̹�C����H�D	{�mp߬̕ö��J���g�7�������P�IA��<�U�ݪ�@���e[�%��@�j�'�R��eBݫ�H���EP̧(����eUO��]q�H�5?���3��t�l��G&�� �0O�$�Gm��B�ލ����C��$05�'�$0D�HL�O1�`]YP
�%�����L^$qZz�P���9��
Q	���xR+	�@��)�GN �=�H����\��L*���O��C�4�~�$�|Ė��=�]�@8}"��C<=�@�Ԇ� 4�`C�35�dJ׎�-%�h�!p�D��(��&v�6�z��'���c�
ӣlm:�)�ɉP=�q�wOZ���(���(��)x�r��g��[����4D�p�VGٙg/��8V@#�E*�N0J��5�V-.�;Pn���8�ȸ���8s@�I�ȓ>x��`ꑪ2��ca
՚�����=��"~ΓFr��"e�ݚr���clN�6L��:޴��+�=�2-�bL��A�)͓����Sm3�O�|�)�1��4r���rb5��'�]��P�(��DH�vj�jƤ��^���p-4D�̫gě�(j]��OY��h[#I!D��0�GE$y�|q�a�˙4�ԓ6A(D����I J���8��	�F`���-D���pf�j��T,J9j�F�F�4D�DD/ӆa�h`�C'J�p���V�3D�,j��T&s�V��§=X��}b�*+D�4�A)ڔ@�Te�v�ݦ}K����'*D���a�jƌ@�&�2�@@���,D��*�VfT��LS��2���,D� �Q�ד~#��C�r�U�h$D���$�	0x����ƄɅR�f���d$D������c�bx����R�n�(��0D�4ѣ#Ƞ-FQ�$�JE����C2D��9�Ά%�4��p$�&p���,D��6朤"
`3�MZ�	s�ZÊ+D�XPM1\^,Y�yE�	��V��y�`�	a��4{T@5InX���!�yB��3���s�����0&ߜ�y�E{߆��F��j*0��a\�y�鎫�F;�R�xRDi�o^��yB���8~�(��Q),*�*f���yc�
y.���q�C�*��8�B���y���s��#�̞N�iZ���y�?<tl���I�L	L�Х�G��y�-ʅz ���,�
���*5��y��ڕ'T�h��ӡ�Ҵ�j��y��
Jˆm�CC��p��U��kܙ�y"�$og�B�&ܾv��sS�^��y�bD�&�B��ML^�6���ђ�y���)��Q0)Z"TҪ@�q�S��y����:���2P�1;y ��6��y���zƺ����;2�*q�5�y��9?uP<�#�@�(�(��Pi��y�k9%�.��'H�_�t��f��y�J��k�h���a��U��Tn�y�/w�,�[1L�?M�1�����yR�J?��{�V8|���P��!�y���-1b�3�EY`mƉ��\*�y¡[�Bq�Q��i@5f7�L�4'F<�y�@��bH��N�'[zl4De��yr�� f� ]& ��y"DV�x�2�3��(V �����M��y"���N����ę�J�!)B)D0�y
� r@�S�#��P	���,X D�@b"O�ɰ�f�	x����I�)�u�"O�9���Γ{;�1��ň�f��!"O���Ć̡W�D��E��z�J-�b"O�p%�ƳD�&�P���qD����"O���#�ޒfn��G�
\-�JQ"OF��#EQ�80�J�)c�>��"O�\a�l�v�Z�b��. Fe�"O�����;p���䂩B�f�F"O��1�� !L�}6��'R��!��"O�XX�Ɗ}14�"��K(E�"B�"OP�G��!5�����̸d���"O�⤫�?4{x0r�� @`� �"O1�GIg�����Q�WO4��"Om�&�	G�P�eB�$챃�"O ���W�4�F}C��S��U�"O��*���cu�D"�)6�N�#�"O�A��B�TsN��Q��1�x���"O(��* $X���{�4a*�ш�"OLIèL�W�t���0{����"O��j����m�4@+2c	�.X�Y� "O�X[#�v��y3�C��I���;"O��(v�E%_��}�e@�(�TD��"O�=��@�J?� �!���"O�!�ë�:bg�IIV��K��4p�"O�	R�f�-;�@�5mZvNE"O� �'�$ӄ,:�쀀U6a�Q"OB����x�y�ՋE�ET���g"Oݪ�fX_�N,Y /�;c5���c"Ot(%�_�k|��{!G�G� �he"O0!8v�׬2���je��9h��7"O����Y�8	��K6�#0��9Y�"O��R���B�̨�`@V6?�F�ʖ"ORI�C�҃ulZmȆO�t���b$"O���#�Z�Kv��u��"O�XRrB\�x��������l	��"OjU�AS�W��(��R#�&dk�"O�	���1=��MR�g�j�$���"O:��5�ؚ2ò䂷��$3�>� �"O����+#4�����π	�b5��"O-��:9l YRe>e��E"O$QS"���V�*�"4��̜��s"O�H1��(c|R�	� Μ<�S�"ON�[Ѓ�:$�6���͡�(�;R"O�`:�[�T"�`�DcU� ��@�"O����RM��(�c�9c����"O���>;��j7���̑"Ob�qӈ�
J��y���G�fd�"O��h�aJ�N�0��GX���YB�"Op��d�B��89�SI�5֕3"O��-��m����pͪ9( |�"O�A��ʍ������ôT����"Oȴ˷IF�l������B�j`�z3"O��� Λ��P���đd9y"O� p���L���F̘%~���k�"O4�0��_%I�x��N���� ��"O�����D�D�Y0}3�=��"O
�A@�Ҫs��30��W ��r"O 쁷&����*��<D��"O�;KY�{q��H�);@��"O���7�͘I���@'�7��)�"OyʷE���](�'Q1?��P�"O�x���'{ϊ萔'@/7�X�"O�@r�ɘ�q���}�v(�"O� �M����0�u�ȒXҒ��"O�\r�D�J��LKg�Ov�-�u"O�}�b���7ܪ���S�[I�t��"O$�#1�Q.rV�*���g&l��f"O�m��"�+�iPRC�05�X�"OH����^؄�ӂ�J�z�pt�V*O���AIQ��� 0ƈz� \(�'=6D�b��y�4А ȏ#{1`U�'$��x���]� ! A�M-�pe �'�P�R�^���� �Q��e!�'�L)$*d��,�G$�*��z
�'LH!��Q�����G�->�	�'�%�b�Dn��	�]1JL	�'u2�I��U��J}+�*�/^�`	�'m\}����Y�$i�&��>��'
�QQ��y��t �&	p�n���'QZ����5l0h(�f��b�'}����+�<N���;�%�L�0�P�<rƃ���� E�E�`!D�Jx�<����;z/�������I
�*�)[z�<���_��%L�8P����O^�<a7	֌?���\�G �bӧY�<q�IZ9<t,�RhǳBb���P�<���F�Bɰ���9���!&�V�<�և��w��pI����gE�W�<����'3�^�	'��/M`�w��L�<��d�$`QT�Ya� qR����D�<�*ٹaM�M�c-^,���xTI�N�<1�.0����AN�'��	p �B�<�@ĀZ��0�e�G�u��#0�}�<I�i��)Ȏ	�M�u��p�$k�v�<)q�>J��B�ܮ}��e�q�<���p��t�B�E� �����U�<QgM�i���'�H 27,U�GeP�<�ɿOR� q�"]�d�A1�v�<�f���{LQ�Թ3��Vh�<�f��F�ڦ��<MjD �@e�e�<�� �4e���8M�~!����h�<��'X�nK~	!$f�1NIdx��F�@�<IPǕ�X�������8�Zݸ��x�<�u�މu�$0�IQ�!^:��gǆt�<3��7gFH$a�'M�Y�d��l�<A�-]�v�d����'4h  �m�<��cՐTM̨�jҙ`CH�S��P�<q$n��@�T�� J��-/�`�@cL�<�AC;u�����/׺UGCp�<i����a�r�-y.)s��h�<q�O��P8>9�d��~�ȺPJGe�<��4uώi	��&��eKU]�<0��s��%�h�ZHY�<�p�	Su��P%.#.���'W�<g�Ǉ"nv19�>l���AS�<�ŭ̖'��1�sKD!�|���JI�<y$M�Ѩ�#)�8Sb6�p�̗~�<I��3G�uh;d��(*a#Tr�<HF�y0�� V���+���цLs�<�b�M�8��ֿ[�z�i �j�<	2CW',zι�<����Cg�<��׆G�Щ d�Ȓp�����V�<Q'�*m ����ߌs��i�$�Q�<ITm�L�l�e�[�R��+f-�Z�<�Ԇ\�:|r�����P��W�<A��ݐ(`�T�d,N5���Q�<�AQ���y�
��Z�"��N�<� ����aڣ%`j%z��ZE���@V"Onaz�A>4�<�h�ǌ`m"OL#A��&}AJ�BAE�v���"O�u ��N�"Y�}A0 �1%+`a��"O� �q�^�>�ӑNB�
0���"O��NCE؊���X!b%9�P"O2͢c�X�g0�\3�D���
�2"O�H3H]TX�EA�u�\9�"O���i-���x� ӱ/괼��"O��Ӡ*^�?�l\��/�8o1�8�"O&�
��aI���$�/6~��F"O쵪Tc�m��
u�� R'~���"Oj�x2�.c����ӆ�H/RIg"On]*�ŝ81 )%�Z�a1A"O��᪋!~����あ5�Le�"O`�	������I#���z�"On�`6/ɤd}P�x������!;�"O��i �)q <]xEhT�n�%"O���%d�
�n���.���}"O�l�f�Y';� ��,�P�d�0#"O0��7c՛pf��7���%���"O��R���T}�BfؑJ���Y�"Ot��d	ω.�P�q2x����"OZq"�f*	�Z�R'��#���z�"O�Eq�	ˠ'�dM��H�=�<	��"O&$B��Z' M�a;�lR���s"O��iU�X�e�A�J^v�>�s3"O�qe�]>< ��ĊD���b�"O�� ���1;&��!�*��k�$�2�"O�ȸ�C�<2蔘���P�x�ԭ��"OT�����1~4}`�υ�5��\K0"Oޠ&훯YT1 �i��~���2"OP!��(������,2���("OXm����f8R����&�&e� "O
 ;�@�0
��S ѝ%�vIpg"Ox���(�a-���Na�*�3R"O8 �5D�"�! �b�!U��"O��A�� �J�2aX�@ �7"O�0{�iE�7e���t`�$s�t�b&"O6���뇲@?b�	%��6��eؤ"O���6Cߣ~��ت6���p@Ӓ"O�0�m�� TSw�t��\�B"Ot���B�y�4	G�䕓s"OJ`hd��#3�9  �Q;=�li0�"O�9�1�_�|~���gF�0�؊�"O"�y�N֮ ����&3$,x�"O`�zbk�=K��� �F�g�,��"O�rGc^'*����ǟ
�6�y�"O������%'���I(Z0lb�"O�T�(C%t���ad,~�ppu"O���	3PHQ3&�_	)k�Y��"O0	��67�@ �Kֽ}]z�F"Ol�B#b���頄�53��X�"OR�BE4ry���cY�5�M2�"O:��&Z�1�`T����MK:!�'"O-��f0���a� %�B);"O��	вO�(,��B�)��ś�"Oe��R09o��넠�V����%"O�I�&�@�d��q������Qp"O�q+���t@����Jp*1"OH@�+O�i�h�Z��
�-�p�a "O� (ܽU<}K��C�N}�� "O�9������ n�/�:����b�<��T�t�v-�&G\n��-��� `�<� xX ��5Z 6Q���#{�tqD"O <�1E��wa��2p�G�Ljl5"OVܢ%��lL�3eŃt��%��"O�Ti��� ���9��P��蘷"O�9yb)��<ȸ��h�3$�Lӓ"Oz���G1,��is51?�Q(s"OܕǢ�6.�}��Ȓ�$��
�"OH0�2��Mh6)�*؃i��a"O�����}
�xJh�!
�d� "O��9�6��Q�Ǖ�8�Ա�"O�� 6k٦<�#��W�i�ڄ�V"O$@�^v<�aGY�l��2�"O��g�:b���c�.��͋�"O"�Zb)[M�\��M)a���A"O�2��=�zU�a�S65z	�P"O�idf�E�u��u�x=�`"O�D�@J�1=v�T����X�����"OX�����MN��I�W�@��$І"O&q�a�9>���2D�4*�ق�"Oș@�c�7'J|�j�ťz��l��"OZ�b�`�!i��Y+	��M�d"Oh�H��_;x<кWͷdT1��"O�yP2j�K׎A CL *�0�"O� AA�4w�M2q�
1E\A�"O����K�c�����wŵ�t�e�<q&@ hmz4L�<Ŏ�`*a�<�/�=of�;��	+��Љ�f�@�<����<O��RA�[
�z����W�<��	�c\�l�6�ؘv�V!U�x�<I�G#D]����X]3^����n�<ѣ��L��@!�i�O�4P��m�s�<YV��2�ND!�D@�+�Y�3eWi�<���6h�6Ų�o9cj�Pb��f�<���Պ�z C�&�r��r�C\�<��*#�P�š+�$����\�<�`�Y�:�+EҫT4:�d�W|�<�)[�g8��YR���o�z���'Wc�<��͔������T>,���K�@]�<�	G9G�ٓ�M]8֤32lX�<��B�-f�,�t#S;���6KW�<I��?W�<�tIOF�9�	�Q�<1��`���N�2x�Θ!"'�O�<���LHh��eB�o�`X�DSG�<i�B��g>����g)*�Z|�!���<�S'l���C��I+y���	�	�n�<����=�p����A�MA|���n�n�<��D�Ia5�B�&F@������s�<�Aݱ�q�*�&v嬑��΃P�<���#mL々�"EN�Q��l�Q�<��JH�!&8}b�f&>r.�Dn�V�<ф�y�A�D� 6�T|i�.P�<	�N�nC�|X�@���X��VM�<y`�O @Q��1c�� _�hRs�<G�YQR0ٔ�_�R(��`�ij�<6C��,��Թ�H���6�P�!f�<��
�'R�H|C�C��f��)[�E�^�<biM2 ��<��K���ڂE�Z�<�a*Y���� `����H���Y�<��N��h��K'.��)��ʘr�'� l����� �lI
�8Z,Or� (�)�'c�(���דі9��'I�&���;v�hP|9�M٣y�J�x>Q��E2E��EK��N�&_�\b`bZ�~X [�i4�?a⅍�'���i�,"�^9(��A�/\���2���M�d�*��ßp�҅
-�8��D�O��@P��7έ�� �q�.ɻ�O�O
�pC��:�)���<�0|�휞;t,��@��q��TȚ�A���S�½?��7 �1K��&�ӵ��� ��
 ���H�t�쐲vY�ۃ�o�P��|��03��E��dF�  �&B���тd#�=�7D��� �a� ԫ`�)@&��}BFQ -0������ C$�{��ݜQ�4�KR)I�ldX!d�<w����n�8$�a�40kА-JE��M�L0�C$�.b��-�"T5�,ؤ�D3<E U�
çY�D��#�A�^����I�0і��oԈ>� ���!)�@ My��?�Bu�kizh�-�*%�ȓ��K�T�ĸ��6߰�Z½i��t���N~����ʇ�<�Ӣ��d��)��Q�.,�xp �icX0��W�|n:ҧ\�,���~t\����g��u�?����?�0<Iԧ��K�������P��OUr�<)�c�5N0t��nB�.�$���Ηi�<9 �Ԕ�`�Åjz(����Y�<�S �)AK�AI�jX�e�T����V�<��ƜM˄%A1Ɖ^E�����i�<��c�sx��f�Gu] ���̞P�<�6"�!��X!
���I�<!U	 6,�#���g��:u��E�<I lQ8����@�a�t8r�A�~�<Q���P�tɃ�_.d���LQq�<�Îy5�(�
��a������U�<�c	�$1�-��e3 ��(ȥjAP�<)�N��CaNP�I,7�bxX���g�<!�'��Z�F�yr/&�L%H�`�<���&R��Z�#��=l�U©`�<��b�5$����K#(��u�ht�<�"��U�5�W���XJ�lE�<a��~��2�
E�aߒP���X�<� , 4g��8��V=4����MSl�<�A��,HU��@��:%��K�f�<i�ɩ��D�ѧ�*����Y�<I��{��=%���`��q�<YF54]�u�6L�89��!�@�w�<��K�,%����7&M�`e⡚fbOl�<��F�3Ut��a�,�vE~(z�͎g�<y �&F�u	s@�� ^4����`�<��M��T��xt@��a׺M��!Td�<a6��&(�6��%�Z�2%i燃Y�<q�/�T�Ȑ��Z�i	����_R�<1&�J		0ԛQ�A�%�P�A�K�<	���61
M�¬G�;���q��H�<IƈV�m� �G�̢mTJu��JG�<��Bºh[@�R7{Jt��F�<�v��+d�J�Bδ&����V*D�<�Ĩ�^%�)I�%]��i�B�<���׊x�l0Y�oR�A�n=���B�<q	
�h�l�B��_�&ʬX�! }�<�3mT�sA�\<
r��y�<Y�H��R���
8_�.� %��r�<�rd�9e�F5p��ʉ/ƈՈ��^k�<����3O���SE�v�ұ.Hg�<!EB˃����&��4��ق@��n�<A��+C+ȕ9��_�E��6�m�<�u��1qX��C�N	��z�ESP�<Y ��rb����T���K�<��L�N�&p*D�Ѭ�(�bkE�<�\�+ˎ!V�
%���h�!�dBr�ޝ�b�3:D�%�s��q�!�Ban#�&G����bI$;�!�DL�C��ӂ�('~`�r�D2k<!��1�tP���6����z!�67m�u��y�BH㲡��0!��EE��"�H�&��7o�Y�!�d��)!8�tF;��Q��M�0�!��T�����H(��P�Q>h�!�$�/�p��� j�l��@$J�_�!�� �xk0 �Bޘ��*��[Cr�!�"O ��;�<�ҕ��<ʵr�"O�S�.!n��ԃt�ρ@8���$"O�5������B%@E5T1�,�	�'���ۺ���G`͊ej<���'��
�B�><�"	��/
*bv@i�'��s"�7�м"�3�­�
�'���*`/�-\k���� 'KHDz�'1��Á�$u*5	�#'!(P!Y�'���aܭ}q@ع���� ⌽8�'%@��r&��9�����Z	ָy���y��P�}��;2����YPhA<�y�f� P����A� ����*�yr�J�(��I�E�,�� R@�Ҽ�y�.Ŕ���6D�)ZV����@/�yRfD�b3����.s|�8$ �0�y����13�@R�N!"`zd���y��F
k��␯� �����y�BD�_����ʇ��r=HP,K�y�՞U��a{F��t6RP1�M��y�!�1l�C�(x��ܑ�)G�i !�ă�4k��
X�<� d�W�2!���3"�!���P��=��.��rg!��W<��1�$��b���PpB%I!�� �J���gǦT�B��G '*!���88���2ǃ�:Mz5���2,!�$\�e1�O��i�a�&�Ɠp!���;�`1UE5T��)���^�!��R�&���9Aza2�K��D�!��_�>�r-s��<(��`�k� M�!�D�i�䡋](`BW$$��$"Or5�%�y�P�[��@�u�a�*O�< ��P�r0r�����i��'+�D��U�LB�1��D�-�*S�'#J��r�\�P|�,�CG	w�"Y��'L�q��mDY��@�*��Պ�"�'g�$�BaO/9h��K�
)��ѱ
�'^����c��E���B60ޑc	�'�<5I&�_�P��%p�!Q%+	�'�f]�m	 "��`��BO��t�'��1P�ē3d�����aɞ 0b���'� E�S�d�ൺ�M�Eb�ț
�'�\��&�ڀa�,��?��$;	�'��\adL]>T	yc��8ô���'��I���-x���#Cc*��Z�'$���L�&r�|aRG	�0:0��'9r�a���"�X��&��$i�'�����/��	 at��B���h�'
��Y���?g�8���.٬k�9r�'3`������b���鄌�M��	[�'b�qcU�׸f��J1�A���*�'1���X�~��0U�d�I�'. y�`Aڒ �I����H0D�'�v����*���&����2�'sД�0�<��<�ckû"5����'Έ��g$��/@\d3,ھ��q��'����Ç)
,tɑ�'O��R�H�'�V�sT�)r*erD��8����'
�D���?��8�b��(�|L3�'�����W7	�B���lh���'��=��A��f�����$7�-�'7z]�d*�-ꜼÓA\+Hi|�	�'���CD!����A��M�l�	�'t���¬�^R��͜ ���	��� P`�@-��fly7��#�*y2d"O��� jE��Ԩsp���>�l��"O(9�rnU�8���P�Ú
[���i�"OT�b',ݵ6z�<��ѩ.�ha�"O�����>)�������-�����"O��{qFR%~��+�c9�6�1"OZ�Yש\�&`*`�Ƨ/05�"�7D��B�ᓔ~�j�"�fq�;&*!D�����N )ީ��fex��`M$D�< T��I��i�ةWf:
��?D�<r�b0C���nַi�^���;D�0+C	�+�x!�)� w�zrƎ<D��ZU��x���j�y�f��&%D�0x�D[2`��Pc���bA<m��$%D���&�3���\6&(D\�#�0D�����8C�|u�q�Vh�f*Ox`RW)�8[���Q�ƅ!2��"O̬�@у~���2'�*=Zՙ�"O�d�͈'L�J���%��|Y��"OұC!�ڱMۘ���Y�9_��"Od�{�@g�hL��M�M]UPg"OJ�	&A�U,��"c�\<��H�c"OЉ�2�2z��|KV��;|�Ȣ�"O䭻��6v�M��JY�)<8�%"O��3o^�{z��Am����"O�<�Un9P�}��K-nؓ"O�M8���^9�e�@�f�МP"O�SM˨H<��@�@�5�N��3"ON}�b��n��I0�Ə*Â��b"O�3U(ݏx�ܵk��V�Z�xLS"O��;a�/�ґPG"ĨI�� �G"Oh��qBD�o+ĕ����0�!�"O�1;�j0�VD��`F�z��a`�"O�xG�E-D���)yv]`"O��i��
D�j#���2Z@^��"O��FM�.�6��W�c.��""O�9�VE�.������cz�%�C"O>�φ�bA��K�f��6e�(c�"O�iRF�=���]��衶"O��W�'VU�����i�(8"O�|�7#̰q�`  �ϊwtN1pt"Ođ+5� Q
�S��TZp�s"O��[��=[�|!!�F�+Cl�;P"O��s�N(q�s��}���P"OZ�;Â�o��I�@�Q��L#�"O"I��%J�������g����"O��8�K�3�taz$��:�2�#F"O�䮇d����փb�!���9�y<'M.�	�C������$ԫ�y���$Z�.p�v/�vu�4��O���y���C��+fH�y�t�A&T�yI�|� �u��&y�4T9��	%�yr�e�,�m����B�y2*_G�Q�tb�6^�����yBc�7$���1O���Ī���yMߡy�����`ܗ�2(��)N�yr��Z	�p�&Մ���c����y�
(*��|r�+U�v@%���@��y���,�&pPwO$u�x�R����y�N��'�����M�$}���ӐC��y�E:db�:tͲ���K.�y#��x��u�fK$�43m7�y�%�O��!jQBݷ��]���ە�y���{��z���1:�#���y
� �*��$V�|a��)�![`"O4l{� wʔ�r��փV�dh��"O���@Íl�ъE�Oކy��"OF ;�O�/�̤��ϝN΂��d"Oȵ��a 0�̌�OM(|���"O��b��:|t�!c�T;)��\b"O4���/��s�H5�`n��'�Z9+'"OTTr˘����Iu��$p��i�"Od��1�
kq"� D�+B�6�;u"O���4J�:�̥�ӂE�A�=;b"O��­H�|X t!u!\���p؄"O�mi@R�	��b��Đ7|%�P"O�-#�P.{b��
A���t�:e��"O��P��Y	���s�N�8RƱ�c"O�Er!c�*GGF܈7�1�*t��"O�q��	D�(���:]s>��"O�-�ь�[p=)lQ7&���"OB�'�L &^�S� #A�x8h�"O��S �@|�2αt� �G"Op$a���?Q��
D6}J`+�"O� �D.4|� a` ��Ii2"O�q��ÝT5�Ѭ�@R09�"Oա��ҾhP��K�>[\b(��'u��{  ���   �  N  �  )  p+  �7  �C  �O  �[  'h  Ws    M�  ��  �  �  -�  x�  ��  ��  A�  ��  2�  ��  �  ��  
�  W�  ��  ��  " � [ � z e- �8 C �P �\ d bj �p �t  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�:Qު(�&� \O@�C�h�6u�=YN����X0"O�5e�-���$@ق !E"Oh�G��&l�<����es��i�"O�MZ2$	7fy|�1痮hlƀ;�"O������'v�:]q�D�`Zq��"O:���(]1��RR-Jv�x�"Ot�t�P9��|���Bxv�p"O\0�`�h��0p�L�m^"u��"O����e��rD6�h�	E?j���"O�����D�> yJ�ƀI!�p��"O�� '����e�qLL%��� "O�%ڣ�%+U��d)�#�ĨR�d,�Ş!��͒�s�i!���m�ȓ>2�|���P:w��q (�"����>��`��ꗍWa$�(��-'Z�t��ȓub0�!�wf.� �͙�,��T)�'3��x5J�.x0i1��=��5��'c�����	�$��e�.�M �'[DT���J��A�3��o�>���'�.X��'9'�P�c$�(otTy��'l��B��΋g��p9�Ǖ�2���h�r�'{<S��:udb1�ΏV��١�'���"g�	L>��۳�̈́?�zX	�'���H0�K�O>t�/�4/⑹�'�H �C�T�`��{bd	'�:��'��!qQh�@��[���"&���K<9���iN0�`=�эpv�AqaC�jV!����x�M��v�s� Zp�!��2|\��"N�RX�a ��)@����J�6��B��y)��Жlی�y�Q"��P[�eʁ[L!���y�K��I�|���
�\Z��)�B�yҦ��]���l��A���1f��y��r��Փ��U0j��k $��y�W������K%aɔ���G4�y
� ���@�ԝ]T����I�� ��G"O����D�sO� ;�Cb�T* "O*q�2JB�s��K��7~��ܨG"O�)��*j\0b�eؕ�x�A�"O��ӓ�S�H�~�`�37�Є��	�p���S�*h��iV�S�9�6�2'�?�C�I3��ZC�IB�%B�혈w�>B�I;� �� �	�1��ұe�NB�	8$~�����C�@ݐő�&�# Y�B�	��X�p�ʵWft�!����v�B�q�MK�.�b�"ȍ��B�ɸ(�ꀈd���&Đ\fg��ҘB�I��p���"NH�q��2�*B�ɍ*|�Y�gڿ��E�bL͆H��B�	"^N&�b��&{Ѭy���ʷ��B�I3f۲��r�'��mB+��"��C䉛#T�𒂀ْn*bp*@�O�M�C�	$:/5�7��>�t0�l�2Q��C��D�^T �͂34�x�e%W�HE�C�I"/8$�9���k&�y W"�B䉍:����`m��G��Zg�ȿ2B䉕Bb���Ř%�����'l� C�I�E�FL�b��gkd��V��,L��B�I�f�zTy�H�0j����9U��C��$��×2(���i>^�C��j�dM+q�T'|����`KvC� `��#�-J�z� 7�^nZC�P-���E����Y�WpHC�	�� �I҃��cT�Ks	�{@C�	4�İ�R���s��K���C�I�k! ��T�^�_!��Ёˑ�G��B�	.uPű�	�NU�ٙ��OH�VC�f�e(5�G?��!7ğ8 �LC䉟S�j�y��G](�R%�E0C�	�,��{'/�:�\��ש� C�1w;��Rg̍���!Y��T�W
�B䉁�H³H�S�����ކS��B�IJ�,��
6TT�Ph�!ޟ+�B�I��-�`� i&�pѕi�9�C�1�,5R�l���@7� 5�C䉼Yi�H����4r*��'�C䉏8��H�%l]5'.ll��ퟋCB�I�hnTS��]�H<�r-�.f�C��+n�t�`�cQ��|���H�x�C�Ɏ5�)�`쑾9ɂm�G�|6B��z��D;#����pcJ#*N^C�	�Zm��Ѳ�,�^����\�i�C�	E5x���*	�jĚ$�_l!�Ås���p���Dn�U����*\v!���@��4�G�A�7T3l��Bq!�d�84�,)�M� q̈́M��aC�h!���+qq����kF\�%�``Ն:!�dG$"{T�[��X �)s����C䉖4�����@�#�j��	ۜۊC�ɚ>���U#H/['�h���ٻ9�`C�I
D.Q�D؄(�4��a턜!,C�ɔi����ްe,��smՑ��B�"#)&ٺ�J�I0���� D�C�ɡOw���aDѰ�.�)�~C��.(�X��A��>18u/��LC�h��Tv$��W�ƈ9v�.<��C�Ɉo�^$���Z=gy�4!@���a��C�ɠ Ҧ\X�i�b�,�HA�S��zB�Iz5��RBح8f&��"�7$��B�)� �yv G��`��D�<nI@�"O��;�A
*n��R��/
�P:a"O&�@��ȃc� a���	T"Ox1�i��$�x8Ɇٰ`�Tɰ"Ov�)���i@|�)����%���!�'��֟@��ɟ���ҟ\������	�<RV��4݆P��D��\�dMT��I���ҟ���ٟ��Iß��럨���E�LU��C)?B��#eԸ?�R5��ҟ���ş���ҟ8����h�I���I|sV�A�☒~�ɨqɝ�+p�U��ݟ\�Iʟ��ԟ�	ן|��̟��	�M�.H;AX�^V��PU���u��4�I�0��ԟ�����џ|�	��ɨ?Մl��^!�|I�g
w�r�	����	џ��Iʟ���$��ȟ4���m�HE� 	�1UT��h�N�v* ��˟�������I����(�	Q���I��&�&D������I�|����8��ɟ�	�(�	�x� ��퓴���W��]�����	�4����`�	џ��	����Ʉ. �+ ELb��������
����	ޟp�����������Iğ���������Ԍ],����j�?R��@c3(���0�����I����Id�I�h�	�� w�4��-��J��k�:yЌ��<��ş��	џ����t�	��,����+`�I�t�X`+n�*L � �D��ٟ��I�@�I�������	��M��?a�c��@��Y:�A٪
-���X�C:��Ɵ`���������	 �R��sHM�^�~� 7�� �,�2����4��D^Ц�K����:��H��>l�Z�2p��M[�l&^ȡ�4��$L�.KT�t������� �����Փq�����1H"b����[y�S�7JD��I J�I�4��eR:�۴P48)�<��T�y��N�4D��&��~۬���I��9m�8�Mӛ'��)�әN>�]nZ�<Y$��xV&0����/8ˢ���<��Y�\ir�&���=�'�?��璙�r ��M
1J
�<�%�<1(O*�Op�o��oҌc���g��8&O
���ȚC�εc��X�Jf�Ɉ�M�i~�>d���*e�𪁐&��f�\~��U�&M�D�� ��O5�['���	�K,F@4�\��Ԍ��W�Z$�'\���"~����%��v�  %k��t̓CS�V��������?ͧ���j$͛�k�����'c�̓&ӛvaw�R����w�6�0?��Ik���0J�/|�
="���*�vq������!?�d�<ͧ�?i��?!���?)�oG�9DE�DO�6Z�J�
��_�Y�dLʟ���ޟ'?��I'1��3tE� �D��0'MDlZ�"�O�Xlڙ�M��x�Ov��O2��3�
'K�p�*3k�F��C���}��k��O�4�ÙF�@�]w��'�<�'��! �Y�fB��;g��V:mzp�'���'lB���]�H��4����?����3���a�#��l����!���<�R�i��O�L�'��7-O¦A��45��,2 �>-6F���^�I��5��L���M�'ޘ�Kҁj�`���|��O�����q�歌14� 02'NҘ��v���ʟ��I���	����zt�*U�ƌ{���V�{���1�?i��?6�i��d�O�b�xӀ�O�Z�kUk=�4P�/V�
Ϣ$�Te�a�I��M������Ѽ>)��O6t��ЀR�^Mka�H�N��t��7�)!T�*P�(�D�>Ybb�<���?���?9���+�0ȑ�N)�b�)�ҽ�?1���d��uSQ�@ٟX��֟�O$��Z�`�%)k q#�D-;"�Y�O�X�'�06�\Ц=@L<�O���W�u�V�34��P���q�ЀP� �镩Ũ^��i>Q�ԥ���%�|�Mԩw�"�D���O���8� ��B�'���'����[����4$E̙"F-�&	���9ԩ�k�� WdP*�?���Y����DQg}bjӸ�JFˇ�4e�����<�|E2�B�!hߴ���4�y��'����W00�A%_��	��+%T"���$
)*���h���'���'r��'�R�'���2d���B6{�\|!7�Œ\�rĨ�4�2�'Br�I���
�ƨ�kT��F�T��YE>@3�4p���O��|��'�R��\��M#�'D��B&O6za��sɓ�d�
�)�'5�4�MΓ�0�H�|�]��Iܟ :��Іr00������(x�M�柸��՟��I`y�v�|�p�1O�d�O�0��؅#J:����A�5=�I1�ɯ���@Ʀus۴�X�Ԛ�-j�8���T8�D0[�r�`�I�:�`��aJ��v�Vї'����$��n�L���� �(#Ɠ\��xGJ�������(�I��<G�d�'(J�t�ǈl�
���M8W����'h�6mJ+l�I��MK��w<�%�FW�$�� �3	�R}ў'�j7m�ܦ�S�4j�č*۴�y�'���j��WQ:�����������B�(���W=!�'��	ȟ��IşX�������`q~�{(�xw�T�v� �9N���'f@7�ל:��O��D럨��<y���fX����|x�c�e6�v�v�b�bd�IB��?%���EE\xC���/&D� �Y;O��@w� g��Ԕ'�PlK��_�W��J]�	gy"�=�Z�ѷ��WP&���nW0g���'���'��O��	�M��a��<񱴰K2��h/�0AQ��ru͓<%�6�'a�'@F�P���v�j$mZ��X6�L��려�y���X�֦y͓�?�4/L��5D�@3e�ʓ�b���� t�)!�\��000 f��c浠P<O��D�OT�$�O����O��?��ңH��q�L	�	���8�{�4��ӟ8�4*ø4�'~6�(����E���kL�dE �N�D'�a�	}}��h��ym��?����
Ϧ���?��郸�}C5b�ǜq�!Ǹd��\ ���)W%�yJ>	*O����O�D�O��s&h�P+�* |ʆ�@��O����<駷i�:Q��'h��'��S	z���Y.Ys�@����*�@��	4�M�ֱi���6�)䟠��E�}:4fH"f[��JTa�/q6bba�R&zX扮B���S%$���i�]���֌,�D%s%���C,��A�c�ҟ��I��\�	̟b>]�'i�7�G?:���l{φ��ᣒ�d�D⒐��sٴ��'�P�c����L�!��a"c�����UE�7�ᦕ:&A��	��?!G�˺Q�|�z�oY��$EYh��KS��8M�dQ�gǒ"���<��?Q��?����?�(� 4��`��`z�Y�I&iօ ��Ǧ�xš��0����\��j���'�N6=�q�����*�/_�{�H��Yٴ �����>�'���'1[�8�4�y�.�4�H Eg$��h!���yB���^�:Y�#L���'������I:(ITD����<6�D1!GD5�	ҟ0������'v 7��@V���O���_#{
>h�p�FV\�4���P�s����#���J}�i��l�M�R�8#1B�4r�Q�s$�&�p��v�H�I�<?�M9�$At�9�'��t/��8O��� �u T+$Nܙ�b��%��p��LQğ���Iџ�D���'���!#g�:�|� o�6�@����'O�6M�/h��D�O@ymӟ�%�杊{��,��h��i��ظq�_$�ɲ�MSP�il6m2,n�6�j����/�Q{e�x����Ƴ���jd�V{z��n@Q�IMyB�'��',��']b�(� ���ȽY�����ğ�q��	�Ms���6�?��?�����'B;��q�w~BL��B�
Xx��S��Z�4E��!k�x�$>)�S�?}@�nF�2tf�	R�+8� �iV��U2���Hyb�Y
<�Qq���%���'��:QhI>!Q��i�h�s���k��'�r�'�2����Y���ܴE��!��q�0�YU��<%�~d�a�)KZ`�A��6�dWi}"�a�&dm;�M��C6ȼ��ǔ�QӺ��	��$�����4�yR�'w0A;5����W�	�?]�Ycr���	{=xi1q���eZ�苚'�r�'��'*��'�� ʇ��$(�lz� H&DŒ���C�O��D�O� oZ�_�r�)���|R�&i��5@C�͡2�8*��͆�6͝x}��b�P�m��?]�a�̦y��?f�2Dâ\��A� P�v<��΅ M�PMHQ��	O>A)O����Oh���O�`c��0{
��FfW-9	n09��OD�D�<Iбix��Z�'�"�'5��O����O.z�$�c�*uܝ��O$�'��7�ߦ�����'�Z0��03��%�U=���.��#P+����zY�\Q/Op��Y^�����	e��xU
�$#������X9�mI���?����?��S�'��ͦ�d%͋J�v8J-X-	�d��eM�2A3̬�	��ش�?QN>�%Q�(�ܴ�ђv��	�����~ ENنW�6�hӔ����j���I���#R�?E�ݘ{yR���@�!���])x1�v`�
�yRT����ǟ�	ןl�I̟��O��5�׉�Q� ���>Z�b,�q�w�
T(���Ox���O@���|��y7��wP6 �nܕ}:v�z4� 4eU:�!a�B�o�?9�O�����)�d6Mo��؃�S5�n�C���<J�5�e�d���ʕi�Փ�'P��Vy�'2"[�	�X
�ć:B� ifEX�U��'j��'s�	��M�����k���d*�O�>���b�l=;�:�ɣ��$�Ѧ}��4Q|�\����N�gZ��n�
Nʆ-�QJo��	#q���3�X�˂��'���ӧ_��.��,��BL.2������R�g̟���ӟ�	�XD���'��}��e���0��p���MM�y8��'g�7�KC���O^MoX�Ӽ��튾�҅A+OX}2H*����<��ipL7͞ߦ����ݦ��?��'��RQ�--�>{7��bd�W�k��A ­K!Y� H�M>1*Ot���O<���O��$�O��d���Bs�z �0�<��ir��0�'@��'���y¤T��p���yl.��T�-u��wD���`���%���?%��=2{VA�u��Wf��)3���Qu���O7[��]�'�Fuj�jJ0 �뮟F��jy�)�G8qX�F�g�v�G�}���'�2�'M�O$�I?�MKQ��?�?�u�F+o��8s
�i+���G��<q��i`2�|r-�>���i9�6�Ŧ�p��1��$��$WNK�U�S͚rEd�m��<Y��|z8SH�#Ye��)*Ox�I����䌬L� �E�1�1�S<O��D�O��d�O����O��?����H�J� a�̍?@� J�N�\yB�'��7m]�sO��O�op�I4d����4j3Tnh�$"O�]�X���D��K��|7�6�Mc�O�!� f�6V��8cWL��G�x���C��U�8Ds���O�����<�(O��OR�$�O�D��L֩	�Ҹ��� �)��I3l�Of�D�<A#�iC��C�'KB�'T�Ӯq�~,��O_�`I���s�r�IX��O��o�>�M3��iW|���Ô)��]�%�˙G�{7-<��LY��۩*�j����<��'<�&(�Yw|���<Q��
gAblj�oҘ�HE����?a��?����?�'�?i����Ҧ��Fڨј6��8��x���{��)H��'a��y�L�O�	�r}�����6D-��y��ِ#��!8��Φ	�޴��ݴ�y��'������I�yʊ� �[�� ������x����E�2EhA3O���?����?���?����)ʩG+�W�F 	B-�K��X*��oڍ;����	���IU�d�'��Dd��N�j=IQ#�*\���`��lZ=�M�i���|��'�"E
�M{�'�
��B$6Z��탓	�H���'cҁj#Y/�|aА�|2S� �I��D�J�U��q���������Z����	�D��`y"d� ���@�O
�$�OԜB� �+X�VU��i�i� Bv,�	��$ 覭��4�y�X� � ��_$�k�/�/r�` #p���_�v_�Qҁ�-�v�Ӻ�]w���Av��
�93�a(��2Mz����gJ���z��?9���?����h����Oo5ΰK>d��;���,}���0��'E�6-�O �O�Ձi�e�B�I\�;eΎ���$W¦��4�?��-�;�M��'��|�rJ�x��us�* (�R��;���O�1l�,�"D�>	�<ͧ�?��?����?�q��_��eqe� ~����lW��
���jUݟ@��쟐%?E��.z��Uc���$�(��i��V���Om���M��'��O���'[�J�.�������X�h��ᒦ"�~��O���Q'\=>�]�����K�y,�i� ����R朖����O��O��4�X�?훦JˎD\���r����n�30�J�	Rh�<�ry����q�O��lZ�M;���nm�b��@����7�]�k�f-�v��M��'�"�؄n��U�����J��1f�,�C��5"�DdA���>��Γ�?Q��?���?����O�B��͆f�8��([�$�Lu��'�2�'�7��)`��i�O�!l�m�I�@�4�Q���#~�p�J�x�L<�g�i�87m�h�	!d����8	�F���2Xa��D:o+f;��.:B�؁+5L�&���'�"�'�b�'��|��-K3~\\a�:����'�W���ܴ8dtxQ��?���B��S��@��@30a~q��b�'��P�'Y��Gśv�c����Y�S�?����U�3�X���%K&D<d��-:�jA�ө\�_2�Ԕ'��D�̨N�N^�G��JӃ�_7�t�j�z`X�	埰������i>��	�'X�7M���CE�;&@��`�N��={F��1,�O����O��D�<����D\ڦ�����"?�9�c#���ve��Mѯ�M#C�i\�xX �i��$�O�9���8Q@t��+�<!�\?\V9� O�5(
]�A��<�-O��D�O(���O����Oʧ<I��d�-g���X�N�E�H�:��iQ�X��\����?�%?Ɋ����w��8g ��[��5:W퀱Q���*y��$���?Q���u"AnZ�<i����Pm�@�U�5:��A�D��<� ḛC�
UiÃP������O`���|���@�BU�Qz��0
̾���O�$�OX˓1����(���'��cĢq3�)
&��'#�����	s<�O��'s�7M�Ŧ����Dӟ+�8�sGK-I�,��C��D�ON�r��o�P�����S���m�"G@e]�T�,��a9���N��'i��'���Sܟ�/ټm0Q��	W�*�9��	ܟ8cڴ8܊���?!r�i��|�w�`��*Q#`���I��\*Hm�p�'m67M���)ߴn�J��޴�yb�'Z��J�L�K�زD��	^Ę�Rt�M![��Y�tKLi��'��	���	���	����88�\B�>0I��T��'X6M�n/��D�O�d%�	�O~�!��ӱ@�.-�HI�W��x�Ð\}r-{�lڞ�?�K|r�'�r���3���˖��x� �����(yg��؀���y2�éj��Ǌ��uG;}�c�Ty$��/=��V�T���Pr+D�z��'��'��O�ɫ�M3��?J�)�����O�1�"K<�?93�i�O��'�*6��Φ��4-�y��<
�&���]
.V]Ӄ�ͳ�MK�'7���.g�h�2EÄ9yX���?}q]c�,�hՇR�*�>�A��ɬ'+��[�'|��'�r�'��'��*`�����x �(�1�L��d�(�O��$�O��l����ן�aش�� ��}�6@ʅX���)��@�'���M�5�i?��F�?u��?O���ĩon5K3�X�*m� �Č�!{|xh6�µ+����ц(��<)��?q���?���7�Б��"��6d�Q$����?Y���������
ҟ��I؟<���?M���()]�<°�H�ʔ�+3?��Q���ݴ	��F:O8� ��	bb��b�7ݚŉ�˻e�P�!����"?���`��8��1Zg���;s��'ࢨh���cH��f�T<:�*�bT�'�b�'�����O��7�M��J��r�f�˓,R,��+�E̔U�PL1/O*�o�H�����M#Q�F�Y��;vm�C.@�Skz��'�ظ郿i{��O$�Z��˷pK ����8h��/A�6�XRF�T�fX�d-i���'��' ��'2�'���7i��6��
X�4���� 8���4�u��O����O�����d���睼3-�A��gW�u��9r#L0�j�`�4H���7O��|��'�?Y�H��Ms�'�ڐ"� ^!�<�3�ؽi�y��'6�R�+O;u����|�[�����"@�(�tMZD舶g3t���	��I���IQy��k�
(r$��O���Op�{1o��@�#��E���qE'����dUܦ���4�yB_�(c���9}y�����;���1�c���	{Y\��Q�?�F��g�(�u7b�OZQ{@�T	q8��*�!��}8�@�O�d�O����O�}z�l�����Z�����ㅞ b����|������'��7�?�i���.֝9���7.�0T7��rf���۴_��V�'-���ֻi���8T���0F�h�b� *��D��>���(H@�3V�-Y�"��<�'�?Q���?����?�C��Gʂp�E��l{d	ID������P����s�I�|�����&?u�	�V!N�c�!�>/:�IBf����X�Otm���M�f�'��O����O����1W�l�����@z(��h M_\�j�Q���%H�|��e��V�'(�	C�����D=r�H�)#��2Ќ�����t�IΟ��i>��'h6�C�Z����و(�J8KB��-(��� X���$���IE�	
���Z˦xٴg ��˛0=���	q��Q ����(�
�{Ѱi�$�O��q��C1~u�b�<���\�k�[��T��ɚG��@�#PcF�d�O����O~���O(��?�*,}� 11��+2ȕ,6$CF���ӟ����M���|r�#"�֓|�K��l�g߄MָQ�� 
��b���>���i��6�H"4Ln�@�I�d�]J~dq�݃L+���]��*�╀�8��%��b1��<Q��?����?yD���4!X�������!���?������d�B���®<	�j��OO��!����?��-i ��\~~���Of��'>Z7����͓��'��Kݍ6�����#3N|r�5�V|��� &A��7;���'���(i��^g�	�V:�T�S�*�.UXb�
@P�����L�I���)�Ky���DՃ���	,t��N0Wz�1�@R�q�����O�o�o�2����M�b����q�M����1IֆD9���uӚ��q�cӒ�	��$p���0L˴prT@^y�΀�a��L�f͉�N.%j��F �y�[�<�	埸�	�L��ԟ4�O�ĸ��3nz�(P���"ݱ�of�P=2�-�<�����'�?q��y�&	)v[P�8r��|��e��DZ*;,�6mΦ�ϓ���i�&J�:7�i�X�a��� �a��-�f�`�p�a�Rt��� '�R�Yy�O��h�&ߜYp�咵LH�+�'t�R�'b�'�ɾ�M�s�������O�;g ���(��P�M`�,�	������ٴ�yrQ��KpΗ�D5� ���5�m�`�;?1#'��u�6ē�y̧9�r$�^w�����V�L�l�x���j��h���O����O��=ڧ�?�@i��	�XxJ �&%"�
s�X��?Q��ia i��T���ܴ���ywȑ�c¢�����Z���tg�y"�kӘ)m蟬h���զ��'��@��n� ��9&/AB�\y8ԭͱO$���K9&��''�i>�����������I�.1�	�"�.o8YGK$���'l6��=_��d�O�+�9O �&C�8%�&-��ɘ�t���K�S}2-k��mZ�<a��i�	:y
��;D�"��\P�z4qr�
&y��I�( x�:��Ժ�Ş|bZ� ʁ��p����Ԭk�E����	۟$��ӟ�Fyr�pӜ]Z�n�O�%XSɐ�4x`�j�28PZ�z�?Of�mG�En��8�Mkúi��D��?Dd<#�ƚ6J	��J�ꟾ%y���i���O~��҅��Z���E��d���5v����:��A�׭��0�cH��y2�'E��'��'�"�iʱ9YH}����># ���sM����O��$ڦa�Fi>��I?�M�I>���O�^`n�#D�W8Kt����>Y��+�>��i�7M�4DӰ
a�d�IԟP�B����dXEʇ�k�\i�g$/0�l�@�ÇV�|L'�|�'�r�'���'gҹ��U0rQ�'�J�	(d��'�"W��(ڴl�z���?��������bO�T��&$M5w���'���Ux�v�|��lZ$��'���ݻ3��ЃHʔwv�٤�N/g�*�C2�J�x�x�y-O���]y���?�,Oi��!m��)��e��}c���O����O���O�	�O����<���iyvPV�Q�v?��sU+��&�5x%�cg��'�n7m!���OJ��'^6-� �tpj�O��5�=)@C͔lxQnڀ�M��cN�M{�'�"�S�qC관#/�*�I�	�V��
)��U�G��$�6�yB�'��'���'~�^>���4'	�`���{/r]�q����M��M��?9��?M~*�3��w���� ��Be�|�qJ�'٢y��7�i���̟(֧��O��$I�g���<OX�T��UF
 
giY�S��5P4Od�����oJ��2���<���?���9E�e�0�B ɚ�Ʉ��?��?Q���֦QǑ˟���� H���$9�����D�:a8u��@������M!�iN��>��Eڡ3��8U��6�p�h��J�<Q��[�l�ԌK�^pH�)O"���51u:֝��?�7�N��B����=�8��U��?9���?	���?i����O�:���:&	����7hXj��!J�O<m�?�����͟��ݴ���y7��vx�������2��qJć�y�cj�>Yl3�M�7/Z(�M��'��́9r��W��vH4\2���	� �!��~�B�V�|rW������IןX��˟�5�M��
G+���y`�E�Hyr	v�$<�O�OB�$�OF��D�$��)C�Tx��]l��CNF�"�PP�'��6MR٦������'�
�'3�>pإ���#U"����//���R�P��ԐY(O�Pc/߿]yR�����E��P�I�M�e�S�ؑ^�d�O��D�O��4�J�jț�ψ�(�OԏlT��k��T?x�����-�6%�Fx�T�d!�O��o���M��iŀ���`��:�A<b9|lҴ�ȟ:��qnZ�<9�F�})�mK����S(OT��X��b-*k��T0�E"� h�'%��<����?I��?���?y����oK�X�Ɉ=D���'��y��'��Ob�ֵ�ҝ���4�?Q/O�Pb!�چ^LL���Ԃ�,s4Ì�h�'g26�[��q��Y��n�<I�%�p� ��!�n#n/|��B`E,?Ѷْ�a
	�:(z��?��<���?q���?���>$f8��E�:/A��UM��?������ᦁ[A�ݟ\��ԟ��O�R|@3�׵8 ��sva[%#�*Ћ�Or��'�<6-�Ȧ��ħ���)�
x��s�D�e�P��{����U�ְG�d�'��t�O�];�.�H�t�6�0MP��aJE*�������h�����)�iyw���O-�:�u��'k/f8�f�*$�����O�dn�N��,��ɝ�M�q*�!��o�7|zE��[!�&�'G�C��i*�D�O�ĳ�Ƚ���q����C6��޸3�Sw+h�L�'���'W��'u��'��JI���j�&�"3�R#X=hP)�4=���:��?	����<�e��y��BK�R�ᣆQ31�Y����6c�46�N馵͓��4��i�O��d%c��牘SR��rB��"�S3�±xnj�I$'D� ��;60('������'4zB�I83yp�Æ���o)����'^"�'BP����4s8Hq��?1� p,���JC�jn�M��1B$p1��>�d�i�6�J�I����păA�t=�4�1���IϟZ@N�+��	#�
HiyR�O4$�E��ɥ8P��`�|�j�Z��I����	�\��n�O�����$ ��ٽ-pR��Q�B%3��gӄ������4���y�#&��0�� �&0�}`K��yb�k�($n��M;F����M��'N��Ѣ��+���&<(�
*>y9"Z�/�s�'��	ɟ���՟,��՟�	ٟ��I-j���V_�7������/h������T
V�#�\p�I����I*�Ma��<��!�P�PŇ��TPanl���n���<Qf��q�v�'T��j���O"&7�/_�iz��(jmPM����'3��J�/	�0��˓U�� C蝠�u�2�D�<q6K��;������<B����P�ߕ�?i��?���?ͧ���U���+jJ��#�b	-��}A@mZPhX���"j�P��4��'-����VKe��oZ�dr�ih�k��G^�=�,D�`R�(��[����?Y�_,iǰ��d�2�������Ȫ���H�h�2]�G�T�K���OH�D�O0���O��'���Zv�=ŗ %�f��H�l������,�I��Ms���9��dӦ]'��C�l<*e9�BU��V 1�/^��ē�%}ӎ��62��7-r� �I51lL��!�x]FP �S��8xhd�[�h:x�'`DV�^y��' r�'G�KՁp�r����%s֖!;��э^���'�� �M�����?I��?�)��}����&[,�����=h期�J�O`l/�M��'+�O��DC�4��-����|�>�*�ϓ�r'd��#N�@M�O�i�(�֝0��(Z~ �����HH��be�#?�fh���?��?Y�S�'����¦��rF�E�����k�Bܒ�$X�.:L��	��@�޴�?AM>Iw]��A�4zj������:G�H�$R9J�N���i�P7퍪:6�{���I%TF�U8��B!#��a�'C�a	eb�"�l��uh٦R�R��'%�៘��ܟ��쟈��|�4/�8��y�ĕ;J� FI[�9� 7S2���d�O0��?�I�OZqoz�ճ�;i���A�C��l��FHQ�Mc�i��$�>�'���U�(h�۴�y��ǏOdl�*��?Ҭ!S��y�F�e1��9@�.%P�'2�i>)�ɾ\C�)!u�ʜ3%�����>&q
%�Iڟ�	�,�'W�7-ܙ���$�O��D��o���nF�'����ɒ&iz⟼�O��n�<�M{�'��i��T�/��X��@z��i 1Oz�d��H�fpB/�9)�I�?���$�ٺKa�'^�d)7�O3yV��۹����'�"�'���'m�>i�I�(UrW@��Xe�<�s@��B\4$�I��MS���?Y�>���4�@1��:Q8�]j2�
v_,��!;O~�o��M��X\��
�4�y��'-P0IҨTe��	�ʈ �Ե���6�z}[c	?��'��i>i����t������Y;%�Әa�f�&끫OO��']$7�B4\
Z�$�O���,�	�O2��R�&5���A���D�YFDx}��zӄxlZ�<O|����?���O ��diI1/z�H�%�1ґg`~2�8w�^��ǳ� m&�x�'��@5+�*,0�4�0�;ki^���'�2�'������Y���4%�T� ��"��U�2�E�3���OڰGzP��0E�v�$�P}Ro~Ӟ�m�П��CP�z���"��\�y�<�a�ģUZ�n��<i�9�@�p�������'T�d/t��0Q�ԡX*$U�+Y��6B#lc���ß��	���I�D�2��ɋc���ʛ�l���s�
L��?1��?q׸ifR��c\��Kݴ��y�,U;g�Nb���S,9� ���'���,�M3'����:	�晟P�fcXO�*]B'�-�$�{wh�R��t�]�""�%������y��Z"e�j��ӧ��;����g ��O�Hm�jԜ��'��W>1�יpg� ��� \�.m��b3?��S�l��4J�FF<�4����M�nz)p&LZ�hu(�S�H
�s_�$�!��L��r��<���zf��[wN*�O�Ѫ3��!W�8Ĺ�.�x:�@$�O4��O"�$�O1���m�Ƃ�/L;<	��fK=h��K@k�PDH��S�4�4��'��B��Ʈ�C�b��g^^���G]\,D6�O]Qr����Fh��ˁ-,�6�O��ѓѧ]�#qF�R�`3o��)�'�IB��\B��ݛU��`���ɡ.vRE �#[��M���՛���O,�?�����@&��(����$ĒF$���f��jr��v�r<%���?!��)	��oZ�<� РHp�D~�@����A�,X&��A;Od�`ϗ2<1��;�d�<�.O�� �o:X�J�"sa�,F�~e�F�'5r7�B� ����O���5"��U�"��p��f�����O 4oZ.�Mc��'U�	�Nn��F����	a�柮de����|@PN]�VDdQx��my��O+n�Q&�����	�#����+5 ޭ�􀋽Z��B�%X�N$ �$ �@���Z�̨4|�|����M#H]�������?�;��i�Ƃ"0'����A�Q�8̓d��e�(�oZ+Zn��<�9�ȅ�ቄ�Fq�̈!���j��æye�Y�u������D�Oh�d�O���Ox�D��,{�y{&��= ����˓o���A�$E�I���'?���7P c�D�/I��jgo\9�q@�O�n��M3�x�O��D�O��Za�ӆ.N���D�B�=N<�	cޞu:61#P���)�~Q&�;3O�'�剋lR���M[� �L�,3Z���ڟ���՟��i>ѕ'i7MZ7�Z��0fA���F�]�t�� Au����'� 7�$�4���'��7MMҦ޴vImaC��	W��e;��>E��Y/��<9�4�yr�'�qpf�H�jĩ9!^�,���u�uk�$nRR��b�ޓ,�|�B��v�H�	�D��������:�g�l�
,�'Ꚓv:P q`��?����?���i9�O���tӦ�O��Dc����BH)X��� ����,�'f7�QަE�si#e�*�	���w�#�~���IC	q��B��^0T� �Ȯh�4P$���'�'���'�� ��!E�aC��Z�O_�B!E{p�'>�U�|�޴[vJ����?����)�6O�̽��/���Da�("g��O�Q�'I87-��c���ħ��K�(mH��䃪g�P��
���.!�R���$N���d���9�@%�ErN>'��xU� E�"��� &���?����?A��?�|B(O��mگ&�(&�B���L�DG�4�`=j2�Nҟ8�	�MkO>�'-���3�M3�$��J�
)R�%���3�
'(\�V
~Ӭ�xӣ|ӄ���Ă�&��-��4�e)Oy"�� /��|)�M�-��
$FN�yB[���Iߟ������̟�O�԰�TFӺ_ʲM�F��	mzY��lgӪh.a�b�'`r����'Gv7=�������h���N
�^X�)��Ǧ���4@�_�b>�؆Gʦ)�$��A�رy��a'ґe���ΓĮy��@I u��1L>�*O���O���I���to�5 ����H�O����OF���<�°i����w�'W��'�bt��*eٸW�Y��Eң�|��'���4ڛV�s�x��	~}DN��ܥ�`1�(�'`u��X~M WAҏ�6�H~2�Ց�u���O��B`M�dX���T�z4�����OJ���O0�d�O��}:��PW��#`�Z/~�<������N$A�'���ې18�	��MӉ�w�Dq���cC���6X*�'87���	�4`����ٴ�yb�'��Ѥ��Hyp�#�"R�h�N]�%����Qc̡kr�'���ܟ@�I��������A�H�������0kCnɜd��і'��6�\O��$�ON�8�9Ob}���?
WI�W)����ʗD��I�M{��i1RO����i��oà,����"!�HLR�E�wZ���r�\#&@ʓ�Qf�+�u�)��<!��]J~HJB+ԒCE�a��IX��?���?���?ͧ��DŦa��)�џph�@M#��yD�;w�l��b�x����4��'���W��ևi�>�oڝ?0�u1jC=� )�%���t�-�%ĕ릁�'��E��.�IH�ې��T�w,��U��%���3�z9z�'4��'s2�'l��'S�^|�wB�$f�j��T&������<���A��넯�����}$�h�R�-1��sU'
Xp
E�G&�����v��鄅g5�6M-?鵥�~;r�>�:�d�W�Ze�խ® Q� �I>�-O`�d�O����O�aPpCP1o��̪��F�y�|ɗ�O\�D�<��i 0\���')��'l���O�(0�D�{H��PO��\�TR�O� �'rH7M��;I<ͧ�"�(C��(0 o2E�:���Bʾ��%�D�UX��3.O��"Cil�ݼ���n�P�%ީp#�3����0)��?����?��S�'����Ha�	-Iq�!�o]#��BGƖ����Iџ��ݴ��'Et�"���z6���JŅ4~�#�&
#PX7�Bܦ�XSK��͓�?�'՘$zD�����������[��m�>1��M�[���<����?q��?����?�(��x��ؚ���dǮi�>h�5�Gئ!S�������ş$?�	�MϻSװ�c⟈I����,%Z�A;�i<^6�C�i>���?E* "�즭ϓ�Dt�!h�Fy�rP��8��l̓��!�p��>ô]�I>�(Ox���Ob�� *T�� �u��=lA.y� �O�d�O>�d�<�E�i'�����'���'�����2+��Fjώ(����'h�'.����v�{�N�%���g��D4��iH!w��@ccgs���I�Ju��0O�5)@��'.��MC6%h�ɟ �� �3G�LX`�,G�K% ���ٟ<��Ο����$D���'�nQ8���M�,���"Pʘ���'Z6-�W��$�O�nE�Ӽ�p���3f̲��B�{� ����<9հi�6�ަ��a
�馅��?Y�'�'!���a��K�,`uGJ�Q낁�_�\��N>�*O��$�O��D�O����O Ru�̔Y�4y�Q�ڸ8vB����<!��i�ı�#�'J��'��t]>�	�bؖ(�R �@�|�e��#�nt�O8Un��M�P�x�O����O��R� RE��
�z�[�@0}r�Hզ7��ʓj����cP��u)"�D�<�ХAp����N�=o����B��?Y��?����?ͧ���Ϧp��؟��S�ʝk�PVK;q��\��a��ٴ�?aO>�3S��ZߴK՛V�n�$|�ԉ��1�	��.�XaF����>7m~����	"�$�@��h<�)�'��w&B�vL�'|���jŗ'?���'���'���'db�'>�9�eg\ %�v���KU5\Lڄ���O��D�O,nZ���u�'^6�2��޶qd�rw�C�E����mQ��a'�`@�4 �v���d��F9O6�dڶ|����aT5\�l��*�Bs8�IӮʭ(fJ���!��<q��?���?��-� E���aM^�\<�Iڶ
�>�?�����������ǟ��	�d�Of�P(V �/n���D:#zT`�O�-�'cV6̈́٦N<�'�
pa��4MDd3qB��M1¨�-f�S%T�N!
�+OZ��ݖE�6����51\��%��k |IVo�<j�����?)��?��S�'��
ئ�A��[	4�p��DL�	q�E+p��44����ڟ\ �4�?iK>q!^���۴(
h}��]k�t�(BN��{�Hr��i}7-J%W�7�h�D��A�4)��q-��'+�$�AF�9l��b�/�V���'f�Iʟ���۟<��ן ��t�TD͢	m��P��V�R��!�ɬ|{v6�
:3���D�O��)�i�Ov(mz�u*`���qQ�1�W�гD�29��Q�M�ľi�O���@��K"��6mv�0U'WA� H8�j�>��A��Es�����$��؃I]g�Iby��'<��"a4��uꈙ7������C�b�'��'&�	��M�rd��?)���?9�g��h�̬����3ކ�9��E���'��כ&o��t'� �c �#N$�QE#�5'�@��o����U��\Xp9W���'@��@0���H⟨���"
U���.]�Kq���)�Ɵ0�	쟴�����E���'~y R�h�x�r�Z!Ybq���'��7[{���OV�n�~�Ӽ� �H��qc�K�.��|��FL�<���i�(7m��i�w��n��<q��<�V`gI4$���MW�`�������1���䓓��O`�d�O�d�O��DL�n�2��'L�&[�^�H�E��j�N�fʛ���/��	ğ���k�ӓ@	�q� h>RB�C ⋠*u�9�Op�n�Md�x�O����O��PA'��L(jmzfϳ��mʂ�(fEV�L�6'Hl6P��;Q)�'#��\~�BrG�0������+R�������i>9�'4R6-�!��Ăr��6��(�S��%L��$�ަ��?��W�Py�4w��V!f�̥���I2O,�m�Ԁ@>D�U����%[7�b�l�	�j�2�9c��g�X|�'��D�wX�P��=w� ��-���� �'���'�B�'^�'1�p���S?lP�4��=e��(���O>�D�O.�n��>�'�&�|B�	;~�u�p��:,���`�сM7�Oءoڝ�M���moj��4�yb�'� 7��5��!�d
�J7� �Dj��7Ƙ��h�5k�'�	ßd������I�ɠPNj1�!�D�5���	ǟĔ'6t6�A�>�d�O�d�|/�15�J<�W,^�(P�`P~~l�>QV�i �7-My�i>���~������v�@�s���4����We� � R�k�kyB�O	�D�c��6�'�@"v�Ωj{(���lT�}cܕ���蟀�	��$��؟b>-�'�*7-&_{�8��ُ2 �'<g��d���O������IS�I�����e�dJ���$�4F p�|K���M�d�i�\�� �i`�$�O:���G��$j$y�e�<!@m�{g��b�Y���"��<�/Of���O����O(�D�O�ʧ�v��4�F�/�D h��U��E��ix��	��'�"�'��y")|��N���Ґ;f		i�@���M�K�oZ��M[q�x�OK��O%h���ip���+�XP3�էP�\a��3M�$�AkhDZĨ@?FГOlʓ�?���?}�(B�
&����-��~��(����?)��?�-O��lZ�c?u�	���	�9��q�@Lܧ{jܨJ'l�)
n`�IW��'������}ߴT�'�vQ��ͦ"� 8j#�&TU��@�'�b��:���q�	��i��I�?�0V�^纛��'
9	�JT� � ����V��^8�U�'�b�'"�'V�>u�	�z�����<_z8e�2�R��E�	 �M���&�?A��P3�v�4�`�c��+9~��a��L����1O�nZ��MS��i7���P�i�$�OB큳(L�hg�x2a?(1���Q
E���*@�Ѹq&(*Q��<G�9��į� ���性Q�|5�ڜi�0j��ԲYV���G��ڠ��'
&_x6|�Bnݵ]�:�+�
z����D�1ؠ��)�,)�T��C�v�e�(���<���Ƅ��t �a�yRi'4������z�͂�1����bn��~d�Y
���}�t���#����K��ۙa���3�lvB��h����d͹��?����g%�0� ���Гu��!s!njz����F"E�1!� Y�����E���ě&�,u����Jݦ1�	Пt�I�?���O.�Q*�.3o�P[��H�p ���M����?I�L%�?)���?��"O?-����;~������*u:�e�4�kb��ܦ��	ݟD���?ـK<�'#���	��Ԯ2pP,[�g�D�S4�i-8�!�O�����<�5���A, \,���9N�ظ�4�i?�'A��z�O�	�O���?t-x�I��*1P ��[�H듷�$8{�1O|�d�OD��/.�ı(���N[~�D��ʀn�����h�5���|Z���q,�x���Xz�x\��%�jS����V�����7���l����P�'$�X0w��������]�@�P����	{_�O`���O��Ob�k(� �I�%II5^�Ԑ2gn�	3�� d$ZQ̓�?���?�-O��(rM�|Z'�)z$����ܷ���Zw��f}��'�b�|�_�8�vȾ>�R��:jTs�N\6$���2S��b}��'��'^�I�c��)�N|�oՋY�B%R��!��M��i��L"�6�'��'��I:z\b?�%�o�^�#��q�l�X�tӄ�$�ObʓK�"��s���'�\c0�d���A���,�R��&v�t��4��D�O6��Q�?>}�s� l�D�À c�yB�����ҽi��I.[Ơ��4������ ��d�: P�����#Q�6E�SO7 T�({`�-?�O���M�u
ՐL-�%�M��^���I��y�����M���?���ږ�x�O������Hjl����H�E��"�bs�@��d��D�'/��yb�'�$�KJ�
�$""��XC
m�P�d�O���R�{j��|B���?)�'�>� )��m0��Y�ǎ�\��<�I�O�zJ|���?��'���j �9yT��<=4�!��4�?�C�.��$�Oh�d�Ol����D�Z�ƴA"e���`��`�> I�V�f@�'�B�'��	h�o���tP���p�<sQ���5�f�'{��'�D�OV����L�7;�24{UF@�'�B����Ҳ#?��˟���my��'�nm�ҟ�,�C��	l^|�rlʪ^xMAԷis�'9���O���P� V��&�S> LC��A�`��ɘǂ������O���<���;��t�+��䟁m8fEx3��2}�2n�?��o����?��&6��1JG��%r2H�_1wH�����!�\7M�O���?Q6�����)�O������d*d�,zv`�T�O6-u�1���c��?q��S�L�<�OjuX��[�=�8X���"c��EӫO���^�$~���O(�D�O��ɵ<�;2�,,�u#�{M@�	E�7�h��'�O�w�FEj�y����
�^��EDۙb/
}p�菈�M�fj�2�?i��?	��j*O�i�Omء�<���h�"bu�m�ӦQ�'��?l�b�"|��}�e�3�	x��S��&q��E
��i[�_�X��/Ty�Oqr�'@�$,U��\�� ǉ%"�#�.,M�=�<Ѩ�2�Oe�'K�J��Z��v��rXj�RKK�	;5�Dї'��'�B���Ah�*�-���.��B]5N���5?fvx[�(?y���?�/O:�䄨]��yR�A)����m=(�P�+u��	����	ݟ��?��> �R'�Ӂfk��ၟ�5�-��!�*t�����I埴�'���<f���N�KAv��#-M1u�Lp�LЎE����'{r�'��O����S|��I$�iS$5��N�,�]���X]@��OF���O��?Y%	�>����O����J9]n=(6��c^��滴7��O>������l�
�=�dU4��5�F�
�XЌp����e����'��ܟQ�NZ���'tr�Oxt�YҌĳf�(�dL(uSڈ���4��ԟ(��L��m0db��'�~���fӀ7 �x�?\�0T�'�bb��(m��'6��'��W�֝ Y����ď�tډ�g�[�C�들?y&m��!Ty�<�~�F��!v1&1�W║\�k���yg.ꟴ��Qy��O��i>��ɲC�� xC�4r�P\ڑ�-Z�dxӭOZlXq�)���xxSIӋ/����fŏ?z�ͺ0m��M[����*c�|��|���?q�'�8�SK�5��E�@MݲF��9�`,^��O��'���]8i���#dĜ�(�\i��l�m�v�'���ST�H����D�	T�z�>�8�eٌ�n��A�B�U��'�	��Z���d�O8�D�<���]�L�����93��#rW:���Z&I����O��D�Ob㟬���$�$9�7�H2y�TI!��2�2B+ϡgq���O&�D�Ovʓ�?A�/����t#��v��
��X�Lohٓ��1�M{���?a���'��/� 8:!3۴}�6�i�◪&c�,Bg	��V��'���'�Ɵ�avd�V�$�'��!\,R1�@iv�3�D%SB�t�`�$$�I̟X�,T1�O���
^+�V�A�IZ��|;�i��U���	K����O;�'���Ε�F ��٤a��j	zCh0	�b��	&.�}�Ԉ,�~z�Iո,��䋚�|�B��S��T}��'\�+�'�2�'���O�iݍR�,�/�@pn�e��tZ�\���	�yx:�y%�*�)��)ɐ��R�G� S��h��L�	�7mV=0H<�d�O���O��<ͧ�?1��WkĈ�Ag�)�<��EX�6`T(D��؏y��	�O譩�/d*6!�CfW(.��U�aa�ئ��dy��	��i>��I֟��*�Jd�= ����Q��]�W󄉻3T�%>��	ԟ��*���"��K�>�Q���e"Xoҟ��@��cyR�'N��'�qO��{!�]�s�,��
D��v��]�@H��X�+���?Y������OaI2mO:��?#̝Z"Eִ.ô��?!���?Q�"�'��lb�*E$@��H�$�}%N�C�X�AQ����O���O��?	�&������_�-�h�JҊ>��T�K-�M���?�����'�2�ҶJB�
شP����.H
=ޕ��ń�Kך�'x�'g�T���W������O③��tʈ�Yv�KS�JRmA̦���Uy��'
b�'�^���'��s�� ���-\�RNT=�p-�)	
��9ưipr�'2�'J��#c-{�H���O6���\h�dET�s�)���y̺���%�����	^y��'�H���O}ɧ�ܴBw.�` ���jH�8Zt�R�kLao��p�I�,����޴�?���?����b�4<�ؙf�����c֧�],��PC]���5A�2���؟H�	U���~B���D��B"������4NV�������!�Mc���?��������?����?����A��(pa~q	4b�W`<۴p�l!(O��|��d�'M��Hk�4P�tEꆦ�{��4 i���d�O��F��)m�����IڟD����֝ 
 �:!OY�eV���k���6�$���pq�?��Iş��Iy.R ��I� :�V�Y��4�?�E$8���Gyr�'c��ǟ��6ƔTqN@�r��#dIȺm�7-�O�q��9O<˓�?���?���?��ɂ�ng��õ�ڈ f��yԂ�	%��)A�i�r�'���'5��'��D�O�,��N��^ݎ$0t�@y����H+�1O���O0���O��d\� Z�n�w��@�7a�$J̬����Ry�[�4�?���?i���?�.O���H�	>5Դi�)`iT��K;[���'��'t�P���-������Oִ�SI�.�ȩ�H�17,L�*FA��ITyr�'"�'�Ҭ��}2�ʴ=o��k��Y�����Mc��?Q(O�HaWd^��'��O��Т��ʎM�PIBV�\�8�!��>����?���E�̓��9OB��o�N\s�T�J<.��C�mz7��<�D3s��F�'���'e��A�>�;�F1���D�����Æ#aJ(�n��T�� �����9O��>��	ȸJ�pxq��!��p��*w�$\�WH�Φe��㟬���?�©O˓S@�G�$Ne��J6B�iQ��i��ј'xRX������wpP(�ׅ�-"�"F�O�,�1ƴi�"�'K�O�1>�6-�OH�D�OT���O��]�h�\�����yX�Xݴ�?)O`��:O��k��'<��Nͼ�BVĂ��l��VM��8�&7��O"�L�Q��ڟ0�	������*���e.�0�C�,UC�H���]�k��7m�OV����OL��?!��?�*O^k���t�Aq�T[�T��BC9*�1oZ�L��ȟ��	:����<����
�j̚{w��r��ٌ��"c�g��?����?���?!p/K�^1���58�8
���%{묠��ˁ�<6-�OD�D�O��Oʓ�?�D#H�|z�LTİEi&mR�(B�� d7g���'�B�'�\��(�(T�����OV�0�%WJ`-@��5���C¦���hy��'���'�"4�'�� � �{d�3��� �%�TDL�oZ�@�	ty�j�mh��'�?������L=e�x+��B�;� m��	ٟ���ٟ@�r����͟��	v�Y2T�(���m�?4ԕ3���%�'6��!a�|�p�$�O*�D����קu���V1Hy14*�)D���X��_��M����?yQ&���;���4�*@�B��?9�}�O��7��_8��mȟ������S
��d�<J@�>�1ل'�:e� ��`����f��%�yҜ|��I�O����@4�b��6��a�d�'��}�I�t��2���k�Ob˓�?��'GH�P̒�R�JH�5���?Ur�O�ʓ^�������'���'*��ʆf�t�11h��ap�P��Io1�-�'�I˟�'ZcdB�X�X6OQ��k��B��^���Oj���2O.��?���?�,O ���;;t�����V3V�f1�U�ц!���'��I����'�"�'���<d���r�<(I�m	&%�E��'(b�'�2�'l�R���tHC����n�4 R���1v��A�Ƴ�M�.Oj�ļ<���?���/B��͓l��[U������"���p�i���'@��'�%`d��sO|jU���s�:0s�C�%�l])��@c�f�'��'�r�'�~yi��'��B�T�{����%��Ir�Lm�͟��	vyb/ѧ�z�H�D�(�R����e���Bs�ƫ"�&��f�T�I͟H�	�rN��p�F��F �������eJ�E��bE��ݔ'&�DӢDj�4��O���O���R�ZA*�B�����u#����n�,�	�Q�"<�~��j�|�dt1,BQ�\��,㦩�2.?�M����?���"����wQҌa��� { �1p�%V\Yҽm��F#<A����'^��Q�m�&G������ 1R�r�An�*�D�O��$�<^���%�8�	���b�>����W�v]z ��O&�mg�I0u���)R��?��O��Ă@
N�l!��jX�H�Y�7�i����b��x�'�ґ|Zc��+a�¸=(��$�Б ��my�O �KP���Op�d�O�ʓ��1����MH:!97'J�(-F�9�$�f(�O��;��O�� {3��Qw`�-X���sIM�T�s3O���?A���?y+OL���KX�|�$�R;`R6�y�
N�G`��	\}��'B�|��'2 �.�yB�]O5�%�f�&A�> %�D�M"���?����?)O�|p$IG�~�	I��qkE�0)أuڴ�?�*O���OD��&/���D�<�;a�.ș��A�`b���Xc<unZ̟��	TyR*�5w�����$���A�AX=�y�)L�kx�$AK�	؟(�I�l�t��\��x��)�H`5oSC�D�b�A�𦱖'��M"G�wӢ	�O%��O~�f�y���*����T�A��n�n�����2��1�IM�I[�g�? 
�9a�E�dR.�j��/�N�i�i��� j�����O����I%���Ic|t	&��>�ԉ�seK�-����4'��Li������O�2$��'�x:$�	{غT�@H7 ��7��O��d�O !I��O����ĺ�����=)3p#ԋ��lŪ����'����E>�)�O���Ot�u�$ ���B'TDD�����]�I�A\�d1�}�'Iɧ5f*I�~��r��:a#�"�����Q�1Op�D�O���<Ith�7�%��":H|P؈�Aί�
<s��xB�'^ҟ|R�'_B V�/N�u�l��z��4��̱8(&�R�yr�'7��'��`�� ��O8N��˺e�\��`�5r:�-@�O����O��O����O
`�0^��z@'�
Z�Xes3�'g�)I�>9��?���?��a���.����N�uH�����иyԕ���E�,!��l�Ɵ\&���ƟI�@A��O^����U.j%��+Ѩ_���9�iB�'�ɓ^U۩��d�Ov�����-�F�C�"�M"6�EJ�&QlZz�*�����5f@
���!����>�yIF�4�MK���?i��W��?i��?Y���*��?��~��@Q��*(�ds�I��"��o�ߟ��I�j�����;�)�ӂ:�,ؘ�a�)��]SV�2�f7�Ӭ�$�On���O4���<�)��Y����7a��z��/5�@�(��ݓE�+����9*�j�Y�d�
�A�> ��'�4��B�I�,U����S� r��;���d��hR�@OA�����F��j�dkwN
F�<t��
ڣx���7CL�hیp��MF���m*Ǩ�~/��+�Lj��z�k�=(|	`
"G�XA�E �<��q�C�����@8(`"i�!頑�S�ᩔ��3+����q.AD��g���1!J�Ѧ���b�'�'���9a�'��6��Tp�m���޴ vA�"!zP���Z��!8�ʓ�"r��[A� d�d��C�ܙ�(On!�,�2Z�DN�\���$Vqre0�+&��@.x0�1��[_�'�������?	�jКq.��U��.�}�!�hO&�?9�O�"yÖfZ(�|1@�mI~�<�7�ȦCv��)��A��ڄssJ��<���i�RQ���cK������O��'>��ȇ?
+,]cլ���cp,^��?!��?)�V�2�>���ì2E�]��U�)�hQ���ӓo]�d�M�1<B���MN�v>�uGy�U*[2t�h�KP3R����K�M[Z�ZEcǝ8�%keY� ��F��Z|�0Gy��3�?�����O�,����?,���s�N�M��z�'��b�ݰp�h�F%P�:!�P�d.�0>��x�ㅫ"\��;ӭ0:,\��F\%�y"$V���6��Oh�d�|
�S��?����?!�l�=EL�*DK1e��Z�%�:��hr�GI�&�0"ŨA�1����%�l#���;k?
�"��!	���Ì�r�^%��GM2 �H��ӌT<�rqP��PZ��b�z���u� JƷ	�۷���rb�T��T��dl��3��S��?�R�JFi�GB�R���"n�x�<���
6���`J�U��= 5ɐ[�'[�"=�'�?Q���:	�Y&��5��!�ҁ�P�<Y$�<�Tȳ��0ef�8��jK�<�!�ȋ)�̠p�Eh��Q��Ip�<�#|��CA��n JqRӌ�q�<1!�$?�dIk@�ʭt'~���E�<�� ��<{�E�w��-|dY2@�J�<QPE��( �PK��wҢLJ�F^�<�rO9B4 "��db��Y�<�7Ԥg�jd�Jè\��_p�<i�"E&�]Q�Y"MO�e����e�<���,`} �RNB�/�!'�d�<��-������4��`��	c�<ٰO��Bf�Fʕ�5~d50V/[D�<�F�ݭa>���3�E���#��SY�<����I����$~���+_V�<A��=(}�2������z!z�<��D%¦��OK�,�!����t�<�HT!
Yۃ���� ��#r�<aA��#�Yy
�G+,���j�w�<�b�"�@����q\��u�<�B��)����NX9o�h�`w�H�<�HςW����D���<XчRE�<�D��(t� R�D~־�+T@�<��,�^�ܫ'DA,oԑ�$Y�<Q���j����NGf�h�#�Sv�<�d��<:�Ե� ���Z׈�(�ÞF�<� >�!�U�U,P��%�+G%�T1�"O$�@ Ԙ|�̍�c��,n6�H"O ���K0�h�I���]a>���"O�ș�K�xM���dėj�>�AV"OflѦ�� 6�T���Î0+ҹ��"O�m���&2��Ò"I�$E����"O�,p��w��h� 'l?BM�&"O��ru�\���P�W/PCdU�"O���GX�*@mZ� Y2��U�@"O�����*�����o����"O6�ɒC��K����3��J�qz�"O(��$+���3��7\ٱg"O$$ ������"�! u-�H "OR�!��ŠJh��p!����C"O�TA�7(�>�H �Z���"O�rkV�w|��'���D�jY�"O��2엾W���g�̟!�`��"O��)��@��Z��C�a���K5"O�yHG��H2u�0韹M�p�'"O�U��Īk�	�R�9i�Ե�"O�H�rf߶$�N�����!���P�'&��fmXw(U�&�9y]��ز`U�9^d�Ŝ�q�L����d���F+.-�i�ҫHU�<��<�֣X7?<��A�k�`����d�?�l�y�E�)p\�˓a@��O",��2v���s�S)6f�4�Q�`W��-��pdkF s �-Ɵ�٦a0�g~"��}`F����S(�\A&�G�2��	��f�:l,�"�O?�	�I�0�Rraϯ[�J1�e$''T��� �e����Q���bq��	�����)0��r��Rw�#�Qڂ��,�,c�P؆��Cy,p+q�%C���2��-CI�Tbpd@
�ыN���0� ��������Rs&�@�/�%P�Ёc5�MtT�c��a1�]80��T�5o.|�\�r�� �u�@�H��y�d�`E@�'��H`&~ㄡ���ď|�ְs��ٝe�Lt�E�ʂlsZ݊3dwؘ�[r��O�-�2�3?�f�3T9k`$u!tDӳxϔX��7	D+�$�o~��9O��IBm�.�h��� b;vk�➿dT� �ej�6Z �k'<O4�b�g7`����=5	��)�6O��0��;�L���_\�Q�H˼"�5�f�[�p@1�E�Q�d �`�R����D 	F]a�J��iW�4<K��'T�
��bC1O@ԩ������kS�|˦�?mDl�3`خ p�K��ol�} �x�'X�Z2A�aǐA���	=�L�Ck¤=�6y"�ڀ~���TIݔ|4&M�g`�O���3?��K.^�����\!l�n��@#�eP�Ģe����5槈��D�>!\PcS�Ύ:̢�̖�5=����v�����:Ol��7y�^U��B�l��������iF��Tt�<t��l̜;�qO:DI2n޽3�.L1��� ���J�b�+w+��@�̃	�_a�@�eh̠��LT�Y�<P� ����P�UJ�'�j�He��H�O�<��g�B�9�4��2C 6a�p��'h}�k�A&���Q�	0N<�2s��;v��=E��'S�EZW�@80��p��5b2�'h0�UF�y�d���Ǉ{t�'�dY�3�]v8� b{C<�2ƍ_6x��1��!�O��a�����~�O�$	�<"-�}MB��*��y�N��1�ؙ���r��rJ��ON����$���J��q#YD�	�W�2<��&"O����j�z�()Y�؀u#�bR8*����{��9O4��	��+�Dx4p���e�<a�&��v zeK�$�հfƓ�<i�G�4q���G'k�ܤ1��բ�u @E,sa|�� j*`��k���j���5P����e�V&B^�0��vk&e�"���p��#d���Fx�� ?��1D�4d� 1d�:"�z��ɓ��I�<�aDG3Y�F�:6��Ѡ�Q]�t5q$�!�)��<!G�3g/\"���Jl��򣁗R�<��*�1BvT��/B�]�����<a$lW�{z"����4d�$caN6o�@�d��9a|"Rc0����L�@1���M��8���m�*��S�? �XK�/ǒ22`uH��7�XCD�	1+�e���Sg�h8#!���y�S��&A�C�I�\���B/@{	�Epc%܉?��Dk�M��jtqO?�	j�*`
V�@��iⲀT�C�(+w�����Tʲ�Hc��̪�ɜѼ`H��'�fT�V���a���r���X����b�P�f�H��Ӳ %n�+���`2T!��:D�Pk����۠g�&M����F�h�'Y��A�Y9T��>�)�lB��&�Ӂ���5�3D�4�Kd!�E@S1e�%��^�Q9T�bHB�)��<9�)���Q���Z�읉s��P�<���\�G��@���w�\�e��<�u�)L�Z�i��bHC���H��+Ĩ܎c��Շ�Iev!����[�#ʚp[��@Fߝd-j �vf)D�K .ʾh�z ��`/
:�� �&P����HL��h��(��h;S�­[��^��3�"O����CU�Fuj�d� R�銖�9o�T�hP�6��s���#�B��������@5�=D��y��0�Θ�́�\9��:
|�`�眩!\i�R�:�Qa��1��%چ�i����C�-�|2f�O^ä,����h�����%^���G�@4'}̄��z�
u��aI�ߊL(���0_1\��g�Q��Tq���<��:>fT�K>�OM\T�G���P���ٍ[8\�
�} \D�ǯ�\͓_�v������DD�IbjB*?�&T-�v��������S��y����'в�ɗ����$�ݴ��'������ܶ
r�9��I�4mJ̹�iA�g�p1pU��*�ČUx�'|O`|��\=I��E8�PY�<�rSQ�h��O,�2��%����O��Hcᄹ�y2j�9r9=A�kD�z:�0 ��0=��"A���'a"T���j���J���j��a*�&C�/�� ꦫJ��y�'�B��O�S52w^���WSg�EenXk*�b�dZ�nY�ē*�ެ�'"��	�O�F�Q0J�g����$E^� �Pg�|�S��yr	I�4= ���Y�P<K �/"��O<�8P����� �-�y�,ɕnn�E��U����B���y��K�ka�}cǞu<�-��
m@ Jǥ�����z~B���f�f�kԇ�~j
@j��4�1cN$�D=��Mֲ:���sW��%i$���I�Y���kL<E䘶mM�����PN� �˞UL�H�R,N�%ưI͓H��[�쉴iE��[.O��3i����`ů^�$�4F�6{�đj�y�F�4��O�9Y��*�'�z!�ӂ�w�����se6p����?y�iP�m�����|j�/ʓ#�d�!Ӱx5 ��&2G�%yB�xZ<� �'s"�]Z�C�ٛ`�8�� �C�`
�k�	 �6����4�y2���v�x���	 }$h���:<t*h wFT�<�ARG����@�6y����&iu �I%M`��'� 1G�� �p"ҔA_�XZ� �0�0<!pɄ��'X�� d��	��M�� H�?3H�I�m۟@��I�V���<�7����~�J��HJ�O�d��;�� r E��n�C�Rlz��<�àShr�O1��l�#푆Hpڕ�@"�k��=�H�����2��ʃ_ Tm�%ၦ�ڔ�F.���'̪�����4 �	P=�xc��)�I.�����H���z�,�`lFg{0�� F�6>*,0B���2��q��;H�m��hh8"�)�<��O��	 �A�@��n�Tt��u�d�4����q��� Z��x��Lm���I�_�)I �_�b��l	��X<�bu�f��Sa�h�<�O,��� ]��M�flH6Q�3FH� �~ �C�Ǥ�?am�(G�� �"\�l��d����0@4�Ԙ�W�̧�Z4�P�C!^$�e`e"O ��qσ�.T�X�Y 9�a���:����F��1�%�I6]>���wÚ�L���[�A��'�Y��� �]!�H��|`T��	�6J.�"�BT���#v��3�D��	̄\@�r��4��  4�Z�mjEU,��l�3� ��O�͙ԭ�"���r�-�:Q��5���$�
1r��Ĭ��{C��p�%�D���ܞM�����f䑺��\�x�6 �nA���$�/6�j8�-U
-�"��I�}'��!E���QҤӴ#�>�Dِ�&�-2�z[#-D(i3"��E�-��N�J0�0�%R�?�"��Wd�<{�!�<}��B�)\�"r�YC�`ϵ�@���P3PR�h���pA�|ۀ �1_A�%D�B�hX@�lߕ���N�kUF�����:ڥ��a�yO�y��Z�Z���m�<�lu�RmD�FsV]�h�	Җ6}���5"X�y+��
0�F� a �����џ �էވ{�J�i�$B5�#�I�	J�%A3��q@�|��靘WѨ�"�P P�* X���iIa2� Q�T��<a2@^!l" �LF���rwl$r�^���}S���qC6A!��M<?��a�3��=>?��0�l
&v�N峃�?��w{�� D�!e�ҟ" �u���F�*�ƅ�d"O���b�
0T�� �&�X薠p�L?|h�A��TTe���n	*����n�:p�\��.�(h��W;@L��o�0W��,I�*�xF���P�"P���7(�s�M�>�`��0/�0J� ;j�sP���G��L{"�?�CBB'�Ġ���+*+l�;C�px�����j�|�y�K����T�թ�~)�4��I9(�X"�0�H�h��'�O����
��:rbG�c+�i�D��Ȫ;Z6p�Oo�bm��L٫��a�R���Ks�(�iȏ�����[,4u��W�@`0�I��`c���.�� ��b(L&�!��h����-q�R�����gt���N�6!�� Yg��I#D�N����(@)!�(�v�����)��ܢ�.�$!�d��X�*�!L�#V��1�ˍZl!�d�4]�{�a)I�y
��c!���r�0�uB.]l���'O�d�!�YnI���Â<�T��#�ץN�!�DV�+��L��� �9�6�;p(�	!�$�� m�`�g+�
��ܛ��̔r!�dQ�!7�`z�l�?e�� ��C�;=T!�:B�z���I:\���s��қ$�!�d0�%�D%�(,2��C�!������.Q��"Γ�M�!�Q�q�HmI���89���3�LV�!�dڳ ��b�h��6����F�V�!�dN�r��l*���wu��*��F�C�!�D����y��fɢ���O<x�!���:���x1a$G'}X�LV��!�D�8T��A
�J\=0���<}'!�$�� 4�{�c�+m���8�$�<M�!�d�$13R��%-�X����e�H!�d��,����MY5F���{d#�P�!��:`r�u�`Í�YF�)�0�!�dT&�p�A��%b\��r��|!�@t�� 6�A)GH8i��<w!�D�7f�`�(f���E J�{f�״o`!�D!�$%k�L�>;b�Ҏ��4K!�G�dԸ��҄Ƌj0x�"S��"�!�U�;rZ�xP�
�-���˃l!�55����HS$A^�s�jWH!�d�"5��H7���d�I_�!�d �n�s�Cϝl?@�P���r�!�$A�y˒"s�Ҙ/"�����<~�!���;�t!i$�GL�u{��ݡT�!�$7� �#%7,�.��!�;m)�S�%�2,bə��/b!��L:r��,��c�>V��,�$�!�D��	 �0y��N�E�@��*���PyRI��y�Lq�s.��m��P�Վɿ�y�fG20z)�Ɠ�g��0Ø1�y�댨ZѾ��WB� Q�;4�0�ybo9-��ԫ�C*�8�CB���y2i��fg���T��{��٨�y�DβF>f��.4l}�]jB����yb	�aԒ�c�ED#qz�,{�/��y��/Ez��h��e���g �y��Fh����oo���2@_�y�J�c�6UQ`�rW��dFI�y�!��Y�퀰i��v�B9�&*�yԮO�i��I��s�h�a�.T��y��J��:d8Uü8�H� ط�y��Z$��X�pk�}������8�y�$��8�
�*1
�'�d�) ��yb,�����!��h9���3�y��� S�T����|�`g5�y
� �Q�%�"n��0�D�7?�TK�"ON)�$
fi��S%��	�s"O�l�)�2h������&DJ�"O2����ُM���
4�סbʦ�a""O���$�C�ml�:5�Y�F�<�S�"O���ĉ�`Vy ���	X�L\X�"O5
F
�$	6�m�	
's��4"OR�SS�g�(�%�5S�HT"O��R'���q]�぀4}DT�B"O��{�gJ�����	,µ˧"O<|��ğ;	�9�,�Q
�"O�<��P�M�t5Z�a���b`"OL��q�� �����*A�)�`"O�)�c̢y>��+�
�tD�E�r"O^@��h�>F�ZP��9{���;V"O%��OB�< m�0@���8�C"O��1���8��y�ىch���5"O��igH�-k�( ���m.$BU"O�)i�k^(.���''�.$>h�a"O��I��j:��s��y�ȑ{P"Opl:40�4��,�"��p"O"�E�*t$�d]�g i�F"O.���,$����dʀ=� �"O�u����C&���p�ݟ2�h�"O���G ��M���:U!^4;�"Oڰ!l�1+,Tq�bۙ&�ay�"O���f8:�8����
b��Yr�"O��7�S(L��0F_ejl��"Or�S�j���u�2 ���l�q"O&�
B�4�����NI�u{���""OZ���m%�ģ�9w@�(f"O�fl�Qi��S��&7�"�3�"O�AI��4c������+�d�r"O�kPmAy�̸�4��*�Y2"O�`�C�������v�ĵ&��"O>��E���H���J��T�'X��3P"O~���96��	���
l?N�� "O��r�	t�H�ɈW0���"Ol�E�l�܋UjF�K�
��0"O�]�d�Ʌ�ԝ�BKJ+��M��"O��HV�X�fȎ�Q��4wҎEȦ"O�9+��8�tz׈G�1���["O�|/YP0Ap�@��>��P��Ċ�y�H���Ba�;����D*�y�	�%�Rڵ�Y4@�0��l�0�yr���	PD��d�#ʰ�"���
�y����'�fd�#D[��=��J��y���i/�¦����kse %�y�Ǐ�z��p�M��l^���/�y�k��Zj1�&�5�
�1�J��y��
u�H��Q�I!dp1ș��'�ў���U�e�A9d2`0��E	}I\��"O�$#T@�e�ʜ��bC'EL���"O��B��v�����]�D@.}��"O��	���-L����!�	�B�c"O�<��	f��H��IXɸ�a�"OZH#�k>�H�D�x�H�Yb"O���S�+2����Ν'S��"O���1@��vE�����ⶦ"O@1�d]�O�0! fL�@f|�z�"OL�Ha�Y	t�@�X0텏r4qag"O�db\(�څF���E��eǷ !��-����ኄ%�� k�cH!�$�?!2�Z�$�+"�F�+3�G6!�� ���e��1 X����ΰ)@�q"OH]baÁ ����4�<`��HS"O���J�4h����&&�dqkR"O@�*Q�Ձ:,�"�!J? ���"OԸX!S��p�!
��у�"On�X�#K1FV:$Ȑ@���2�ˆ"O��@�n��1�dO�,f��ŉ�"O��7kF=)��Q
%-��,�*��r"O�=�b�.B�dha,Jh����$"O�I�#,��~�V�ȲD��<�����"O:	�DG�7#`���yp��"O�)	�[g8mrUE�"]o��E"O���fkҥ<���Qg\�J�Ӵ"OR�h�
F<mZ��%V�is,Qz�"O-�AO�&��Y�R%j�U�"O�zF)�?sEP͡d��=_� ��"O��@�o����(�ׂ��iG �i"O�ؙ���9<� x�gG"^b,*"O6 0ц fJ�z��Ո0�䊢"Ob��.�2f���! ':��c"O�<�f%�9U강Q�����,�"O�d�g]E�ݓ��[R��\Z�"OD)�&��NڄU��A.�xa�q"O��v�a'霽rx6Px "O,b��!E�BIR�G:8dj���"O�D+�.��c�FXq�f �-J@�C�"Ov1��H�^�|\�E��8��P8�"O$)Ig@2�tXg�7c��|�&"OFp����/��t�䇎E*2�{�"O���EJ�+"��}pWf��m,��"On�j�R:&w�7�ʞ~�
�"O��C��ٔ?���JV�<����'"O��8�"S\�0�*U��\�Dm "O:��gۧ[U`D2��/{6�"O:[�U�NxԸ婀 -n�\���o����	�<I���B/G_~�3C�Q��yr�V=�i:WH'2dӨ�5�y�KP� �r�
����r]j��y� mH�����W7�\�]h�'ap�Z�̘$ �7+��K
�'0&=©WE|���B�O&.�l��'"H}څ��:�\��H�%v����'�qѡĤ9��(��cA�_j||����&�2����hXD%��	]-Od�ȓ;���b�@���`y�a�%c����f,8�S4�X	y�]qf�
�{����ȓ2�����DZX���e��C�6T����軠�Z�a`pi���#�FD��S1"�+��@���� ��9�p͆�S0��"��
���A�Ty�4aS"O�f@�6uŰk���t,v"O�����Q�V6�|@,8_�y4"O�A{�̹>����rXd��"O�ݩE	G��h�"�䕜@�!�"O��6J�t��\��nË��)R"OlaC�H�+da,��ҀK ��KV"O6iɱa�Dɠ��J�-m�L�"O�J�V�j���#Bm�P�v"O�
�	�v��) 7�߂H�n��"Ox"�CʪE�$��vmH�"O�`�6�A	��9��CJx���"O��ɴHՁB������*JT�@"O�@�ņ�m�d�:&Ř,(6�TC3"O���b�IS�����m(n��"O� *[��G7v7�@�=F��Q�"O��D��Qg0��F��:#��@ "O�)����S	P2fX(8��X�"Oz����\ �0���aE`̈%"O^��GG A�!�޺Q)nh8R"O�KtK�$g�ּ���R��ɉw"OXɚ�%����y���n.����"O���!Q5�n�+v����2�!�$�#a�ؘP )V7��A�
�?4�!�D�C���q�S'�D1�h�P�!�S�I�P4b����R?	h!�݋����Ę�+YjXh�Y59�!�$4_&1��fǳk�b��ʘ�
�!�dLV��Y0�#cjJ3`��,t�!��^ɸ�ir"�23p���tУ1�!�Ո,�]��U�C_ڝ���,�!�d�4X.}!���Q>�`�l��!�d��~���Sa$]�NK�]f"�9�'a4�*#�W�X#d�� �>Y���k�'-�D��B�&��@%W#V���H�'�*i�fF�e��$W���B�K	�'���ؑ+!]��1��ލ-�p��'��5���#!t�)�	4I��r�'v�L�m��t]D�h�gM�j*��h�'Fȑ2#F�`MM:兓c""	��'}�������&4ruD�T5\�p
�'6~�kq�\�O��)�D(��[��U!	�'���aC)��C���G+bV�p��'�����!X82X��$B1
e�I�'Bj�h`%�l�b�FgK� 6��
�'�v���fO.Rì����
�r�v�A	�'�t`c���U.���T�ϗ �����'R�A��Y�$�V� �ˉ �p�	�'�`̠7��D�!0G,_�f���'�Xy���&J �H1��� L$���'M���b�Ŋߖ�
!`4q/�=��'_&=�Q��#/]�(R�'e�"�'���A�M[�6��y
'M>j�щ�''�т����ȌQvD֫]?���'f�ˤ@��L>y�d^�q�U��'�yCq�Fc�����ě�(��!S�'��	�鈢z_����x��b
�'����G��/��ۂH�tNpz�'�,Ԁ�$
3yp<��ŠI�sA�P �'q G��0"�x�b�T1�r��'�{�FJ�pM���,R��9�'�)�jH�"2.S����U��'���f�
kr��� �ĜN4���';�|�0CPA\�H���ƸyW�]�
�'hJXaʏ�C��ʑH���
�'>rP�5N��~�`��и(3´
�'>�u�G�&��Q+܆i�Ţ	�'�pѣ�� z=)R@�����'��XRg.��M��Mn�R���'�=j��� ܘѶ�PQ��j�'�µL�hž�#����N�rDj�'���	߽-�q��GRP�>��
�'�X���*�"1T�E�u��Ez�]�	�'������� nt#թ�)h��:�'����b���|T�|��m��y��ߧb��ٚehխt�hA�p�
��y"�V8*J`��.�?o�t�1 ��%�y�"
�?���%� \�2� UΟ�y�˖3�A �G Ph�D%�3�y
� ��b#M��PC�ϔ[0f �"O@����8������\�*>� �"OT��p��E5���Ռ�p�@�"O$�b�˺�����jΨ��"O�k�W2�\Hk���lJ�2F"OB�3��1#A DZ)̄4<r�xe"O�"5p���$O
d6���"O�� �������!˜̡D"O�9�0PݣTdP�?��|��"On�3G�2lb�L��<am0�"O�QHG��	}�A��.%��*�"O\(�9䮜 �=6\��E"O���W"�(Zs��CP0?ɘl��"O��ŬLc �s�oG�d�H�9�"O�u3�I[l��������b"O\x&��'n�}�G��2w��� "O-�BJ�c��(X��;�����"O(xA6/�u���Q� �J���!4"O6�b�-�Kz�8P�S�S0�m{"O�(rG��
O!��$�$|�x��"O�hc@+��{�H	���\��Ha"O�}�ԮG=~�=�V$8X[B�{�"O��(d�G�������C���"O��h4dޒ`��	�TCX�c$�)��"O��yK�?���A��.�N-C�"O�8	a��=,�\��%B�FܤY�"O"A���+�� �(�vp[�"OĈ8h�9?�5qkL�Ba\p@"O4	:��ɇKk�Ӣ�ܒ\Z(i�$"O��afD��Po�\Zb)H�Glx��"OVt{B#kJ�ty��Ͽ0�n�;�"O0�8���Xq��b�Q�^y�Pb�"O΍8̉��(�C֒�6�J"O��'��7(�|��7�=�����"O�¯���f(P20t�<��"O}��8RQ�͈�`�5�!Q�"O���F	,QJz�� ��j�"5p�"O������~�^`���FI�r)
�"OPqq�ۀv�|��/N�'-@�"O����ڋ{���A���hB�"O���)F�I�>��DJ�^p��"O�i���J�t�<UK��7s�ёs"O��%(�"1��B�+=1iQ"O�� t���]*b)�V�I4k#x�"O���J^60�j$���4���2"O�X����$���3S�2��Az�"O����iب�>L㣮�)q��@�"O� `W��Zfp�n�8���x�"O\	��%����ȣ��U2a<�-�@"O��1��8�\e D�g�[E"O0-�c��?]�5{� 1z�R-�"O 0˥GV&!2�y��;\}�x[�"OZ}�����Jp���
ptj�"O|xc_�a�:%q��X�id�P�"O�|��`���J=qĤÀ@'0�J%"O�,@�e��,�\��E��D�¶"O���T(��t\|���X2�B��D"Ob��Ĉ}�f}�*�56��5XA"O ���Kv�hY�
��/zX� "OMɲ@�".����D�#� ��"O��w�\"d2a@cS�:�^xS�"O�!T.ǡ9�����8)�:m"e"OV���d 0�:`�+g����"O�����fX�B�� �V"O� �0�M m�.l�7�;���@"O`M���A�V��A�=M|��A"On;W�F��`/�Ѡ�Z�"OV< �OQ9ժ� ���	�dR"O�tؑhCX>�!�@5~�<5�"O��b�
���C�e�� ��i�"O�%:���U¢�"R����dK�"Opȡ7�^�=ں�cT@���)��"O���׀��҄`S]��Y�"O��ՎR�s�X���e֘o� ���"O�E��J[�_h�)pN?:j܍�"O�ѣ���m�2�sCT�5cJ)��"O����
)~�zi�"b�WD�M� "O� i�,� 6�6�ɣ� HX�9�3"O
x��-ɏL���s`(�)LU !1"O�,��/@m�R��L�k<� �"O"}Y�شi� �M[L�l��"O,���/4$���P~�4���"O�-���!/�i�Ŏ��Q�����"Ol�Ip�Iyb:d����Z�1Q"O��T��8%0MZ�D֊��b"O�u���ڂ0=������!l�t�e"Ot�t�̆x��y㬊�PT���""O�Pb�o�;G�o���(�"O(�9��Y�y�xQc�i�'*��� B"O֨��JΞf���r�W)I����"O�c4��XМ́�&9*�h�c"O��T���GW~��DY�4�hb"O<-���� �&   ��
���"O�dYt$��@���g�Q(� Q��"Ot���@��rHB X{�XR�"O ��� ݠ	�ܲ剒K�R��"ON�J4�L6S5>�c�=t�v@҆"O���(�4��$"�!V6t~6�(�"O8��gT�\���� ��Wy�\�`"O����
ƾb>@���NSDf!!�"OP̲b�!#[��D��]����"O1a���)"ڥ�P�ơ7A� #�"O@����R�M�
�!�/��qG^̺E"O��K�.�[����&#<p]��"O����Α�A�p �N�K�Ps�"OL$�� N�y�
&�*LB,L��"OI*c<^񂑋"m�+=��(p"Ox��T��"=M��r2ś�>*���"O�p��AV�i�BL���@�R���u"O����~E
�lAE��)"O0����7"��ȡH*~����"O��k��E��Y�G�3>�T�"O*h0��w�U)��<�.L��"O���!֦{,���gf���e"O�!�[�x%n@�e�E���e"Ol����� ��B�dj��;"O�-1��I"%ḥc#��6BlD�a"O�1���F�6��>n729q�"OhL3Rl��]���p��e$��P�"OqQ��_�ŋ$�+:��"O�+�/Gd�*���gT�]� 0�C"O^� \�J�;$�՚_���jF₌�yb�U?'��h5�T�Z9���g[)�y�9"����!K �񆧞+�yb)��Khi�0�ȍ?"��cc�Ҧ�y�d��P%H�"vŕ72�dU�QlȽ�y��ZDEb�cݐ(��14���y"���4PF"In��yb����y
� bBD��4_��4jq�ޗꆑX�"O�e�e�NI�} @̌&]���j�"O��@&�B�&�
���6��Q�"O�a��;[�Щ�_����"O�5�wҽ�h,��+��H��%!�"O��q5&�H���K�0�IRb"O&\RIF�Wj`{BkʭW0�8�Q"O �1Go�>jn��5�����1��"O�( lQ�;"��A��J�g�p"O�}:�.���4����40L"O�	 �f�4T�����^9��d��"O8�z�I�Xe�Ң%F���k�"O��"Y���Cv�� �"O�uib�;y�LPU��MX���B"O���#��`pI�B��D��"O���N�j9vA�"��n���'"O�5{��G�'>�  F㙢��<�"O���aI�'mGz�r#�]/6$%9�"O�y3� Ȉ)���@T6,r�"O�� d��t&�0#��W=I�zٲ�"O
�90��!ZUΤX$��%�"|�"O
�*&��>��$���%�\�Y�"O|��$�2mz.��A�A+!����"O$d0����L�6t:��A���p�w"O��s�ŝ"(��HKc+ʝ?�`y��"O�l���$��Bri�t��L�"Oj��AK.W�$E��Y4�`Q�v"O��r��b�j@�w	��w!�e��"O��>Z�V�p)�+:'\ly�"O����˦:�>�����y*d�"O$��5�ΥWD��E�]�8��"O�I+�H*�5�S�H�g�y��I{yr�	�K�����OV�6�� J�b^���߽-:�Dˤv/�5���YP�B�I�+3� [&�0�����7�C�	(�*TG�i�ta��k�0��C�2l�9���1u���:]jC䉤mD5 ��Æ�:�S�Z.>DC䉴|�>��w�.1�J	I��Y.�F��d�O�c�d���R <r(`�&T�g�l�r��1�D5ړ��Dt��b�_;(�8��r	��`^@�Vd$D�0)�ʋ&q!��R�,�'|akU� D�|��<�����\�NaYa�
2D�B�)L�b�  �ն<���s�*0D��!gfD-*�R�i��,��x#��9D����"o{�I���ap���Q@6|O@c��I�Q<B)�<0�E?(Ԃ�y��8��r�'��ɭu�<�ȑ���b��C@H\C�	�]��HZs��DxP詀�#�FC䉀]��|�`DI4�<D�cǌT�6C��*7l�� �H�@] TC�Y�-�C�	3N�X�d�^��}��M؝"��B�"��A�b�ZV̵� #U)y�C�	Z���E�=SXX�j�"G6�=����f��%lѣQ�<l�(0*��(��!D��t#&l�@�AV+7�0$a�<D���jL�R���%˔u_F�Ȧ7D�����&I��ɓ�n�tQ�l3D�0�7�V  �]���U�h�E�0D��2`!P���`�F�4d�l-$�-D�@����J�˘v$hq �%+�OP�}�<U�7�@';�T$ɐ����Hi��DǦ�rQ��]��F�X��ȓ��IB-X<sB��UAPOX��S�? ,Ԡ�K�#�ꁘ���s��"O�us�)C}����A��-8U"O )��Hͬ� �Ф��"-���'�B�'a|��QӖ�����1~��t�
ͳ�y�.H/U�1棞�t�Թ�%�$�y�B��B[½��dO�k��p���E��y�%<W�A���5���D"�y�̚[��uѱ�Ц3A�I��U��y�DO�g!�ũ� �W�2|�&�'�y2���@�<+�,=z��1�Q��7���0>%OKYC�}#�`�\��֦�T����<�d^�8i�Q�W";�A GO�<���	���c��aVW�Pp�<�%ω_�t�&蘓:B~ɚ�Hb�<IU�ۿ�N��Ҵ"5�T�eC�\�<Y��N(/����Ό3E�> ��LXU�<tkL��pF���Dq�X����Пp��ٟ$��	�,�	��"[�H���1��C䉎Y� �!7"Y�V�T>T��C�	bӤ�9E��tu�C$�?2StC䉁e��=2�Ċ/;~�ԱG��B{8C�ɋr.��U��d�R�7�E�"�
C�	�8�d�0 ��\q��ҕ�B2U¸B䉙d nD��K���y&�'NjC�I5w�܅���^��r�тT�F�B�	�pH�i�GE'yj4QcT�8B�I"ޜ�Y�`�� �Z����W�1�.C��s�LAqA$�0Vu���E�7FB䉊v��h+թ��B:Hd���$B�I�S�B͘ì	�g�^Q������C䉓cf)q$I�58N"��t�G;qTB�	/M����#O9Xq)WAp �B�	��:m�0���N#2)١M\��,��I�x�Y�.E�U�az����h|�B�e+�P��(ҚU�4h�#)�B�I0���'!	�r�b�US�JC��}x���ؐ�<���iV�$\��:;�Ѝ����BY:@��'�>������yT&M:G©���D����,�<��db��mF�v#�$�D�*O(˓�0=Q�+�;�`Z�M^(�VeTV�<A��9v��قnW�Mܪ�(7�Yv�<���"�|!�E���	�̬���f�<)$&��.���t,�c6�!m�_x�XGx��\�c����,�����2'�/�y2l�6`>��%��`w2u{#�:��?�'�Ɣ�v,�;itʴ��&�X�u�����0=�
I/�����ŝV�  'Ln�<i�l�2q�I� q�\��Z^�<�Ca�B�qS�ו�9B�T�<&��e�����fhRea�LQ���<�gi$��M�%���3�)�F��f�<�,�	*�jH�t�T�٘�៼D{����� a��"w��AN�*�H ��4D�Уqj<�ix���(0�
h5D��@3��)D�$�����<�l�s�3D�Xٳ)�5�h���K&
(;�7D�̻ăG8ʼL��N��Af�6<O��d�O����iIg�D-�~\4��&DTy��X�F�:D������#�=:~���I�b(rE�4kFl�X�.�� �f�%���Ia���3f�R4(`�)E>�ܒ$� D�< �Eόu�Ȑ��;x'�h���=D��[!��"w��l�'@�]ҍ��	 D�� ���aK�:pN�*�d�O�^U�7�'er��ـ�
k"ԈDB8��yBቪ"
�3AS�KD<�#H&!B��=Aq����&:@E v&��2[�O���D��� 8����J���p��˩0�!���Sx 3�X�j��ݫ`Ƌ�Y�!�(W�"�ȅ��;u��l
���Ry!��(�"y�P�
��������a!�$6 m��
&���"1�LI{"�{���>ղ#m�T���#��@�V!�.B�ʨ(C���(<�sꎇ;��'7a| H�
E�Q8!, /�⛌�y$�%?"�Y'�"x���P ���y�̃�ʴT#`aW'C�	�u̺�yr�$64[u���>C��(pʟ �yB"D�N��p"�=E2D\���˜��>��O"�aE�
vT�+�HI4V�8I�"O�5	��+p4i��p�4���|��'�5IM�0x��rs���|䘙��'�0��tk\W�&���&{����'kx$�#��:b`!��C�;o��	�'f���E���R�����q  �"�'��r�T�'��:���0k
�5��'iL�e,1~XP�A3_�.TC�'���3l�0e�8���QOj�Q(OZ����w�lH�S�.���u��!�D�,w$��&A��\�b�4�Pyr�!8[��
��W�	���K��yR�.=�����@�`�A� 銠��<a���'��y��$O��T`Pg^5s�F z�'�>�p��-B�y��+�&C��(���hO1�~�=46u�#!�+}Z�j"�� 
$|�ȓI:���f�ɪvwFᢇ��tk΁�ȓ|bf<icNF��Z����Q�����ȓp�
9�_��'h�-��i��r}$:��'P۠���	k��8�ȓ?Vd�����q9搙HЙD��!�ȓc)���A�݁@4 ����E_���ȓkVt��P�(���ǝ����p�d-2��m֠M����`P�ȓhj"��7������a+���ȓu1.��t�X� �\��m
�M/`���̎YqD	�-��I���+3 ��ȓP�h���iͪO���:��H�[�6}��Iz~�ҠX8��:`D[�I�>L�g�/�y�V+:d�E�υ?D��J���y�j�	 &��R�ػ�'�*�y�bˈ ���K�H����S����y�-p�Z4�͟�}N��[�[>�yb΃�D�����h)Nh���(	�y�yj�`������,@����'�R���ޭ"&M��*�N,�`JD3B�()�?)��85��Ò�p+���M@0)V��ȓ)x��#L�-�~����O/Q�z0�ȓ<L:i3#��*�>�@C��1J*x$�ȓ�\���uN��!+����ȓ[pi�BþPh�-ӲL$n���hK桃�\6`��S���.��]%�ؗ'ca���m��ur4� )����m��y�`
�]�hs#��"s0��"�ҽ�y�%Ⱥy��E�b���qD<��qi��y�(�87'r�(	�{�h08� ݐ�y����4�Y����n�~PAe�9�y��4���B�a�^ȁ��烌�y
� �������h��T	Gb���PW�xF{��i(%%R���9,����Ζ�-�!��SA�Q:�'�*�~���Kr!�D��B��	���8t��L9&�ċo!�ׂ��@ҫ^$J�J��P�ËE�!�d��
ve��j� ������I��!�đu��!]	Xy���w��@����J,����C'R�,�������D%�S�O�����(4ǚ�aB�%l��}q�'�$����d� )ۆf8��s�'/�v���(P��ZO�52�'z��#C�ظo/�D��- M�xUA�'��k�)w�F=��
�l�(�
�'��,Xd�ɀY����'������'I��#!��"����]�צ�h���hO?���*�=$<Ap(*:y�a9`�F{�<9F�_�� �M�Bu�h��s�<Yv��(��k$gh���`�`��ȓ�Ș��U�pQBw�[�*4��V��yV��]_(���.@�/�لȓ�4��	k)D]�&��v��-�ȓ_��x`�X�d��,��m�V��'Eў��0�'dps��.��U��Jْn�཈N>��Ȃ:���9 K����k�2oi^��ȓ����%�K�&H���g����n����(;W*D�>�d۰n�#@��ȓ <���F�%�(�"1,\0'f�܄�\�|�tQ�V��lP�����&`��G����Cϙ%f��3��-��m��U,0���4plė2J�bUQf74�[�E�+nJ��CaI{hf�9��Af�<�$�[�?�8\i0'��;�����H�l�<i�N5@���7�L�����f�Ks�<9$e�#&�T��'�e�����p�<�HǴ{��<0���{��i�<I#%ǐ<�4��nڬ��%����p�<iw!^�
<�Z!	&w�m��L�A�<���N����!g�j&�ö'U���Io����KK�_3�ř5eU�؀�"O�L3�� ���?h��%jN7Q�!��ϡq��ҥȉ"���AFݓ*�!�H-0��d"��33�$�HPV�!��S0r��I���L�H�X��]�!���|���b��b`�L���!�dޝ{.�Ѻ,�]�D��%TY!�X�o@`��mI�
V��j��A�HX!��K؁q�0Ut�fI�|C!�$�$7�;"��@���AG`P=!���6X���Х �>3�8d���4K/!������Ė��J�����V!�$�4N�k�M�)0�� !�G!򄉫 4�H���T�L�����Y b!�$�5N����8S�$��I)_�!�Ɂ%b8���GW�[�0��qÓ�f�!��P�x���N4v�D���5=�!����ڧ�^;����c�!���t��Qۇ�[�o�<QBP�Eu!��^<��R�Ĉ8p���򢜻Zg!��-i4Y��5xh��ք}l!�$6/m�y1�LJ�i�0�g���M!��_94-nES��r�0��4O��7U!�$I	Y�8�A��^�%�R93�j!���@�}��θA�J�3�:vP!���@1�Py�^�P���aPE@�+E!�� ^��I_�3"��BL�'D��S�"O����)
ed@�*ڌ4�0��"O�9@Ѣ]��QR疼i�X��'"O��Zo�	��3�cV+T�:8�0"OLi����	K��"u��2��L{2"O0h�FH�@�Dj J�Y�JX�"Oعb�$%~�	��ڽ*�p-h�"O Y�D1�P㶈 ^I��aP"O0#4KUz�P���<4B\s�"O|Hx5kY�w���p,�Tn �"OZ$�ٴlhtMc'	�'y#>y�@
>D��򢩀t�����תKw��[��:D�$Д/�V�
�@�F6
����9D�XK��80�`P �N ML-W`9D� �*�"i���*I�E��1�*O���Y�y�)�ƃ®Ѹ�J�"O.�Ж�,L�*�i������ �"O�p�&F�"~°�2��Z4�"3"O��fb,?�"�n.-�Ą��"O�a4FU�TPЈ�#m܍� \"Oڐx�
��'�|x� X��4�u"O�����xO�< ��F�O�`�{T�'�!�ğ��<��4��?G�n�kF�F�7�!�$]9������,<��z#hK3S1!򄌮H�ʠʶ�Ǒh$tᨗH�7%!�$ڬ"E�h����$�0I&�@�!��Z�7y���!� ^��m+�ף>�!�B )�Z����bVX%�&'��L�!�$M>`�nqfC�}ke�0�ݟ`�!��73Ӱ�X�	MX�)���7�!�DD�/�LP{5��R��d�����U�!��_�C�l�³ψ�H3d!��!���4�R�
ҏV�L`�郰/ȥ.!�D
�
2@0������Q����b4!�D�-Q��U
�' *J���ে7g�!�D��*�έZ�E�v�89f�K2�!���P(�1`W�X�����ГP"O��b6d90+nU�M)�"O.�{	Z7p�p4��Q*Fp��"O@��0�L� ��|�����o4�"O��(�L���2#cSB[=Hs�'���`oT<PHPh4��Ω�q?D��f!� �(1�D��\wf�k��O.�O��D7�3}2�~����M4Z���e��yre*lZ��p�ͦ~hA�ebH�y��/C\�]c4�G,	�d]��1�y��;��T��M�}$�(��K�y���%<��{1A� H��X9�AƟ��=�����$�0wQ"���DS�;'E!��y|=O�)� 
�sO���Q�[(\L&y(V�'gў"~r�iǽ�4Eڄd�l�|������y2��M����J�D=03��&�yB#M�B@�����3R�𲫓�yRś,e�N����N]��)��:�y���RɁ�!�}�n!{�l)��=�/O���nP���N�Q	�j����j���O�ʓ�?A�*�;/�>�
%�� D���+Y�y¯
LL �V��'c>���b���y���
-U�mq�O�8��}x7��y��K�b<B9:gY�t�����z�<�᠔ L��,P#F9hA�����S�<!p�'�J����s����R��K�<�S��$̡�kÏ;�i���m��D�<�kY�3�������k�~�9W�O��L�� �IH
��G��ȉ����pK0"O��P��19�P�G���(B"O�Tc���-�$ ���������v"Oa*C�A�wW�l�1�	g��Ƞw"O�ڒi�%��
#ND�B�@H�"Oj HEH��Bx��L���� �OE�E���( ب7��S ړ�0<� �[Z�,�J��,v7����j
}�<��0c�,Q@�..�kf(�_�<qE�
�Y���kĮ�(��8�6�Za�<���np�b�@���%�&?�B�	*pE`��!V�L���	�=Ir��$�O@�w�PrT���m3��4lTh0�ѐ�$<O>#<a�`I��l�G
��FF�`DD�I�؄�I�'/��3
�!	zBAUHFs�B�ɕ6���#�N��]���$x'B䉤{��I����X_�%�S���F�C��
~S���Q(5��-3bDA�F��C��3$K2��`І.��E����`ؾ��D�<�'2��Ie�Ǿ4ʚm���<~cj��
�����?\f����'[�����hT>X!�Զ���DJ��va	�P!�d��	lR`)�O
<�p�s�h��t!�dG#7buS΀#P{\�(D��'�!�$Q�2��`6,�>x�4H�+�!��%>D�AJFj2U�v1����k�{�'��?O�Щ�AǬ>��1�]5e�ث��'�'n �A�l��N���^�/HL(��'�!�����QJe��P-N�	�&V!��
��1��ʹ9�ԭD�R!�D��-C�*�-�b��1I-�2 �!򄛮�x�u犈Mlf�za�N%X�!�Z�[�z��C��WžT�� �.r*!�$�]^9����<0X�ܫN�!�J�p�����!&O2�a����
k��)�Y^rȄK��_�@Ɂ�֕Y�q�
�';�`ƪ��b|@f�1=6���
�'��}p$K�G��сB��$U����xa&5b4�A�!�d��'lî0�p�����b����� ��M�tP@�ȓzh�|�dƲ#9<xjD�,HxT�<��+�@�Il�'"��ʥ" �{[�p�oMct���'�(HZ�OF9`?��QCǕz@,�̓e��a�"m~�=����X\nC�ɩ]�`<�b��=/��eh ��Ri.C�I��\�r@�ӣ�jy�5��?-C��G���ǲ
@<��H�!�B�	,�u�/G#W�Q3$����P'����-��ā��˗e*^)XG�)~l����\�'������?5��j$GM�Qw��"#7D�,`�(.4G��CEMO�]1X�a D�$��a��cPTm�aAӨ7�℡d=D�\����R��|����	iNİ��'D��+ ��?oK��ҥ�Y��@��8D�d؅K�1p
qa�D�8Lؐ��5D��ZbAց��p����-���e�2D�DD��`�`�Sl�&�Ɣ2 �.D�H�Œ��|��+s��TBt�-D�0AfM�U�`	b��.�b0�4�7D��+d��:�F)Y���Li
Ṡ�5D�8�DS''��g͟c���� a0D��0'��
#?8�E%Ie��`D&.D��c&mırmZ@@ �Ha��У�7D�,���J�!�o�1w�9[��6D�� �U�BL O|r��5%Y�P`12"O|`��A|�hQn��',ɀC"O�i��v+�5�bC�M(�g"O�`�N�d���@Ac��q�"O�:�¯^��e!Pǂ-bBiCe"O`9v�'�le3V�޼R��@Z'"O�M�R��E*,��r&ٚb�q�"O(`	"�ψe�r$�������"O�u��иJ����aM�)�ܺ�"O��Vm\�A�|����^�1��ijQ"O�4��ԙtȦ1������f�|b�)���nQ���(0
�t3���=�jC�2@��A���c���6%VI�C䉋0�H cc�t�����ȑN!jC�I�4��)�E	�A�f�U.8�dC�I�7k�񓒠]�@�T�bf*NiTC䉿2Rk���!m�N�¶�M0TC�	�o����ǅg�*$[ "��>�.C�I�m��E��J4 �";2i �4�2C��\P�(Q ��41l�ׄ�.3C�I�-�r�8I K�P���׉ǸC�>DXڡ(����!1�����Ӊs�C�	�\ĺ$	��N�h���$�Ɗ/"B�ɴ(~L;PnҎx�ha����1S�C�	�G���5k?VL<�㧊ۓ%� �O��=�}����#&Ӓ Z@�� h3t�G�<!u��!n��p
_vD���k�w�<I���%�:M�7+D23�"��d�w�<��LLou�!W#@�&������j�<���/\2�Iq�)�*�i�c�<1E�H?'��k�G����"���c�<��_<-�L[�E1�d k@��Ih<Yb&�y���,Y)���[%�A�y��,��x�Ȟ�ny豀�2�y"-�Qj�ѱ@�X��@�AgA��y�/Q�����@ձl�F�R�H��y���y�hc���7a�x��C΂��y"�U������lX�6h� �y���-r�2d�c�0C�(`fᒱ�y�D��y�z:�)V�H+:� ����y���-}m�݃�b��NV��č�8�y���,t��,z� ��{�*3���yb�N0=ŦA�#���>���G��y��]"��3����:Ț6-X��ybeF�N�� ��zɢl��g��yBl�\�Ƹt9t������yBh1}�&�OV�����@�yb�؊[��ap��<AJ~����;�y�)�`� bd�i�@0�-O��yjP�B�ص��o���ZQ`ʕ�yR���bL�$�tg�	"Vꆟ�y�,d�^�0�(h'���tAK��yb`�Ig���+�?Z�|!1�m
�y�*�7gj��Э�)Xh�9���˫�y�,z�8	�� P�@��/š�y"��@��	��-�[�n��RLK��y"��BEFӆU�PD��YH"O�ųeAS���9�1da��"O������#[�䍳Q�
�`a#�"OTm{��I�;���aW@U4C�<���"O�p���{�!��ѢK��E�R"On�SV� �p��0مA�+m���0"O�Y)���� �����:�V`��"OxIɕ�\+W'2�K%/��N�c"O� d�AN]@���nXoT칤"OJ��� Wڥ1c��"v3�ܢ�"O�P˖�a9lٙؘ
P���"O�Pc��G-:�҄��,c�u�"O*}5��7,\����h}d��T��%LO6�ECΨ*�M@�K�ڹA�"O��S�L38w�����2V��"O�p#(��0�Έ����\�pС"O`�(V'F�%������ٳ��C�"O�<sSݹDn�����R{>IB"O��xVB�
�0Q�U%�
We�p:�"O�Xx'��&D�i梛5gT��`"O��&�0-����Ё��?����"O��[�O�4o�T�G Y ���bg"O$�isl�K��Wd�L�"O~ �G�X:8n�L0N��+},�"OJ�i6�ޜ&T�d�qf�,qb�Yb"O��@��@=~� �k¬$�u9�"O����a��#ͤP�QjR)��0�p"O.9�6��?C!�@����k�Jh�v"O4��SGP kD X��ށ�.�q�"O����y�����tѳ�"O��j�
�(xo(I���R�M��""OȽjFW�2���P"
�jа "O"Y��J=9|�%��%E�h	��"O
T��BT:�(0�o
�'�v��"O���wb�j��І�%=:�2B"O�!�A�!�IPF�&K/�!"OL]��e�/k���T�^>p-�m(c"O�-�� P>���jǄ��:(By��"O�س2�:�DM��0w��	g"ONERn� �(�U�ͼ=�4xu"OP�xP�ɰjNX���1���"Oh��4�Q��H�BٟG����"O�)@�G�0t����$�� ���:�"OJ�@(�pD��JAA�z$���*O��hW�N �h�P��¥��[�';��Ҁ ��`za���}>ԛ
�'7I
'@t"�x:#͊�L~�q�'ʶ��!���^�,+��H,���'����Y��rF�5;qhl�"On�XՊQ%.�Xi��ٶ�Y�'�ŋƎ)*P�Y����)5�>8��';��ӨAab�9�	5$T�J�'/`�ĩ��$g�ih�M��1l�:�'�ڔ[�A���D�@�X�.��-s�'\VT����G.��i&Fţ&@��Z
�'s�� �(.�h��ʀ/wft�	�'>~�"#
�k=(=�׮ŷ����'���0�3n��k�iXH��'FZ4��=&&�)V��cXq�
�'G��t��TtZvj�p���;	�'L��qi�?@XM1�!�h��i
�'e�����h��`���*�c�'�b��X&dRl��Z(�p�8�'�`�Hr��_���������{�'�pA��̈�?H)C!�����'��d�uFنC�����ؠw����'�A3��Z��*��GB:X��'��x8��H*��<P4C	+I����'<��	C�R�4i�A#5��J�]��'�>��Q��0|H�4�� ;�r�	�'Ϧ�!�gٵN'0A���-�r�'EV"���m�TkB�	*|x���� �u�fƐ;�l�Z���A�X�"O*� �J�/G�YY�b0`"8  $"OJkaʂ1h[v��#k��.��"O�`q�Q�]�0��AILe���G"O�=���Ȍ"��,B3B�Q�"O��чg	y|�x�6�)T}p�D"O�$�aZ�?>��B�Ƌ0��"O��hF�����P�
/�%�#"O�q2�͈ �p�ا�
�G"O����=,Әݐd	07}ds�"O���ä[�v����ƜX�j��""O�a`EG�B��#D���n��"OpȻ� ��fP�cBR�(@g"OBm+ׁ�x�i����
 �)�"OHHcf�
p�Mc��̘Jt4�0"O@M8Oa`]y�-_�Op��"O\�s�O�9.�T!f�0n�@�: "O����o�%!z���p1��"O�l#D��(Ur4�1L�tr��*�"O��cg�/J��Ă/m�ł�"O����P�(�D�YU�1�r`�2"O����&h�,	ImN�fB20s�"O������TX|!�����)`�0S"O��a$hަm�,=�㍒=]�,��"O�E�#���F=�3s��[J-#"On�*!$�.:վ�rBG=d�eqv"O,�� �!E�������}�.��E"O
%�%KF�[? �;��Z�;i2	Y!"O�{Q��3,� )R�Ϯ4�!+�"O1���C��%(�cW�-	�CB"OB]H����Z�Bt3R��?�X��!"O���ĝ�y�$e�� +R����q"O�i�p�Z-L���.�	K�Ɓ[�"OR���W>r��@��l˼$���&"O`%{��T�x09Fɒ�`��X��"O��U!Q�
�#��  ����"O�� "� ~�8����W'8���"O`�j`�!D�r,�(U'�>��"O�5q�L�*Q����F�A�tM�"O͢�K�.����d��%��8��"Ov�R��K�@�{�"E#DQ����"Od��GJ\C���n:�jC"OD �%!P�
�<�z�܀
Fp"O��9�dQ͊�A40�b�"Ov8���=fI�5��I�H18a"O9��Ę�)���M���"O�dn� SX��!��	dxE"O\��TH�B�!�J�!�F��E"O��D��+)��{)�'�,��"O�jGb�:E�ГML����"Ot�#*��#��k�-*���!"Ov�ŀ[00ܼq�q��w�<��"O����	��HP(8ېH�73�`�i$"OH�H��
�V��ELD=ѓ"O�U�Q�8��P�R��Z�"O��+q���q9F�H�%- Bj&"OnDˢ�3}洓QNKb���2�"O��
���XSP��­\�9�"O��qML1n���B�	3T3"O<��1��F*�#�$߼
�J�"O�T��b�W�t�1�Þ-P�:10"O,�X6��V���`ōǽfӐ ;�"O^��A&5���� �\�u��0(�"O>}��DK�%��ӈ�t�$T�"O� �H���R�$��������E"O����� bT\��A���\�"OqBr��;C��� t��?S� ��B"O���@#Аe�b� R�^��-�"O`�9E�J f4��%ƒdS�"OJ���h].m��XeE!�v@�"O���%C$R�J���P
/�̨�#"O�4K�H���Ub���t��l��"O� �2���&D�A�m��
�\��"Oԙ�� ˣt,�1��/���A!"ORݱ�O�z����D�%�(d�@"Oz���琳E��i�Q�ͤJĲ��"O2�*�&�/��}{��M:H�1R�"Od(���\�T�pgE�#���3"O��A�oȬM���$d�rf�)"Ov\�Tl�2)R`���8��(�"OQk�>�R9����<}�L-��"O	�&���2� �;��ds�"O�+��8�A�Q��h:�"OX�Ja��"[Th�w���Vp�r"O��Sa�ɯ]b(�衁�(�@c"Ot1��їi�Y6&U�	���C�"O𠒃.��$Rj�Y��̍j�
5��"Oz�H:0*vXn�u��$is"O�|�P�M�E,Ո�B�c��]�"O��cRaƗ�<`�T�<���2"O�T�"������k�^""O�܃��,^�ny��$[i!�"O��"E B+�V�매��1M��k1"O�U���d"
� '��,:�tA+�"OB�c�G�EҼ��r��'�.�'"O`A�u�ԲV��P	4ᔱ\��M��"O���(�7h��(QB��E� ��"O`!f+T��ؑ����D,�
�'��JS�� ���Tj|
�'c���G�ղ! D ;Fk�d}$I�'����n�J��0a�X*0���'��e��f�"��嘮8�ؠ0�'1���2LY�f\.@���<�J2�':������b��U�2]�9��'���B�ٰh�zAb޼QZ����'���d�ܼ{Vic1�0O*&0�''����)E�w�]��D�89v���'l"a�łqNvU�VÊ, �y��'m�P3T抭*�fAF���sDe�V�<I祒>j����.ݗU5H3��P�<y�폄.�T�PFC�^�*&a�I�<a�^��:�i�rmH����JL�<�2C�. }ڍ���E�t���f�S�<�A$��G:�Sg�>t~��	O�<�T�/x(�B��V8!�` �3�	A�<�� �
d�K��\)An�4�d��u�<����9ʠ�pa����0��Ln�<��_�;�d��hF*�p@nO�<�Qȅ8b�p�S1�	�N�|����N�<��h��l�վq�� ��D�<��I���ҕ͗&z���1�DG�<!��ijD駦O `��ѩW�D�<	B��~p8�xū�G��x ��}�<)�=�ļxc��~�aF�^|�<t�)p �ADB<
d� #��P�<�s�_�+�6lB�މQ�2��N�<	�ꈂ��A�a��#HY���G�<I��G�F���! �W02�z���A�<� E���.9U�U�#�&�` �"O�	%"�%�PD٠�b���{�"O�d�G�9>��e��6��d0�"OB�1�-޼F�ڀ�#�>cZ,���"O���OG-N�f���@T�K̅�R"O@ A!�@;0,����/�(FD��"O�MC���]�Pqp�.�0@�|x�"OF�BE%�T�.�kw���diC�"O�Z'm4N�؅�C�Kl
��"O0����	r�0�h˔W��z�"O4��qNC��px��pO�8�w"O�i��)^3}a�x��%�!��"Ob)�!G@#y���T M� �J�"O� aG�+Nc�H�@�80�y��"OE�B���SR)À����"O����I ��1�(����8�"O��HTN^�|�� �W��M���#7"O`����Jv��"� �7~F�!"O0b�f�XR�/1<�B�iބ�y����	#����4#��:򬉠�y�傁?�rm �N'�~� ,���y"kW9m�R�8wDN(���yUA��y�DN5u,B�jT'Лh�l�9��Ȇ�y"EʫJ��ZV$ЮgD������y��%�TT��+�>�4���!�y"���J&���EG�5��	��kY,�yB��3+����DO/5`HvM�F�-D��[e��D�Ę��P+ ��H��.D��B�M��#�����g��.�Q�A8D������]CL����<�(ݓ��6D�x���v�$���<���.D��Y ��T�L�!TcҺo�`��`+D��Ѥ��Z�0�gJP (l��HK(D�p`���v,� �5"K�hӔe*���IP� U*�+�#' a�݁g�jB�������$.R����{�VB�	>3�͑TM�6,X�JE% (�B�	������/\�MVnt�
׬*�΢=�çF�
��TG�AR(��v��'y�`������׈	�hT��K�mG&���y�~9t�D���6�������T�]ԛ�k��f�A�#@>�� `©�ybH�v/X@���i=(-�qC���O^�P��,�'LER�� �K�>9�(S5Hބ *�\�ȓJV���DL�D+���BЉdC<�',ў"}�ɔ#l�Ȁ+��űA�vt8e�A�<�2��*>�j�+��
,/�����X{�<iDn$Q� Z$Tgk�1i�L�<Y�ǻv� �\e��Z��ãmx!�Q	B���Q�M]�N�$C�(y�b��T�OB�TxŉNp��흑Z���@�"O`p�s�!O=�Ĭ�3nfd@"O"5rd]4ؤ-��T�=|��!��'N��o�xEI���q|�9#Ɓ�z���W®Œ��߅H)~%[�ȝ?}��l��g2�l9Q�75�@3W�ķSx�$�����'�1O��ɴ�ٍ:f�!���?9:�BW�'Xў"~Z#��Z����NX�J��y�����yb�1e�,8cE��>��{r���'O��i�>�� (:�Ɖ%-�������|��w�,���� R��'(�a��m�ҵ��.�=q�D��e^�`�����?J4I����)p0����x�<y�e��(��(%��l˾)����<� �$Z����!B�*DT�x={�"O~="U�S56|,�*`d�&��Pk�"O�mhQ�}}V�㷤׿��DB�"OpU�!�N�9�A���2�T�p�"O�����I�������@8�q���*D���U�D~�Z��EP#Y\�p�������'�l�[�&lF�$�VΈ�p�q	ߓ�M�M�4Ó��+�3&�g�����$&D��IG!Ȳ*��<�!��Mb�2.c���Ob�IIܧ����<��5*�F�GI0��4��|�@B�I;4{�4����6(��4C�>vZB�	�r:����I�N�0U���e�����)}R˗{��4p'�	>�b����M	�'~F��FI�c�a�1��^`��
�'�l��e�4xs�� $YZ4d��'.^t���ņn�*��w<�Xm
O<�����ۏ��-�b+�Lms��T?!�I'I��`�`3n�ȝ���>!!��E��]ƌZ �R��%��=
ar�Op@�Fօ;*B�H�K��.��"r"O@#%Тj�3AE�����x�C���O��sV*�3퐐!4̢�O��V0[��р�@�7Cz�p���6��XD{����pA�4g|*�	�㖘u����"Ob�pH�5v�*�gS�Xe��\�O;��!t���w��x��8�ʓ��3��J#'�����3BeL0���2�:"J� PP�ʖN	�F�zm�ȓ6�޴
���=h���S��2fN=��
��ph�E�H!BKʲ:}अȓpظ�����|IU�+�h��Y�1K'ˬ*��H�ǝ�ai֩�ȓ,�>�����2.^t-�u-N�@^��� U�p1�ҵ;��A�f�!7Ȕ�[���s��K��T(J��Ѐ��F'�TY5n:D� ���S�Jd�Ԑ ��Z��T�F$D�02��>?>��0���4[�k�#�O��	�mnR<0''�p~�{v��Z�B�I ��i�_�`�f�����=�ç�8�6#�<ez �(�"l���6D���
��3J&г�k.���j6'v���^�S��M�c��7�<��ˆJah���HRh�<����%"����`gнIZ���by��'�<�fU�v��`���� �=y���I��x�T���d����T��)t�B�	�j����'v~�	�)��qv:�6����.�=6����B���S!K*D�$��e�0T����D
HU�9��=D�L����O�,(�ǉ#q�uf9D�ҷLZ/|�)��+ńo��=�� �<�9�O�a�a�*u)��� �`�BQSQ�����Ӹ���&�p~j�.� V	K������y�&��\�@$χ�*,+b��(O�`Dz*���j�
g�t�e�B�,�v�	n��uG�'���zfV�R�fh���4iU���+!�S��?頥H7'�0MKҫ5���b�F�'5axB�<��W��L��P0"�&�y"
	�%�.MhC�.=����G�ƣ��$&�d4�'u��C�"�����ڴ/���HN}�Մ�7{�*,ٗi11݂�ȓ84J���čX�#��?7�<�ȓ- ��8a�L���X󉜸k��:�'(ʅ���$1�ZI3�JA�g"�� �'M�`c��X�hL*�NΘn ����� ����2a�63���l��Y��i��I�</O�㞤��N�y���
�=#"m���&�C��iҡ�DY�nNA����o܀��E�M��V�|bX�b>OV�r��E�[��x�/g*4,���r�O�0��픿
p<X�u������'$�A1D_��]�C!Yp*�'&��i�@��Ka�&U ,�'�e@��^�L Q�Y0H|s��D$�'A�����a^s�ܝI��(]T�)��$�\e��:Rt���E�,�܆��,��&K����D@2VC�$'�TF{�����g<q�%�^���B?��'v�6�	J�ď FN�Z7S�Xd<����M��'��z�:���cVj,²L�`���y���+��`B��{7�=8 B"ў"~�%���3���{�xӔhT*y���ȓw2�f�'O����]78���i9���*�d�хl���@�Fx��)e/C|�<��-��O5މq5#�i�<�S!(I�$	�� �V�;c�Rj�<��`�%z�qT�H*4OB!I��i�<��e׉4Y�v��'vj��d�b~b�)§8I(�w�M�v�1�n�.P��,��W<���&*�xI���x��Q�7G�j�<1&L�S�H�g�ߍ|[�43�LB�<Q&&�#8��q��O��{��0T�~���hO�'z���Ņ�$��Dޏ> ���+V���PbۃLf8;�#D'�
݆ȓN~����L��f�r2IX:P����ȓ<�ti�kӰaE i�$�u��ȓj�.E��q��kv"R�d[����w�
�+�iʥMKN�B�F�P���ȓ%@�At�ݽ>�f}"�-܇#�|��e�,�CV��z�LRB&�W�^X��}�f��!��ʚ�[fj8I�y�ȓi6p ���;&�@��69�����*���V N8I�5�`��&@��̇ȓf���	TOȃ�IQ"����ȓD�-q��/Fl��3/��;	�����
�@��N�&�Na�B[<`9>h�ȓm��*��O��H��Q9_��ц�<=�8�-��x� �$J�4/y$���{����� v���ώD��!�ȓd��ŋ^?Y���sFY}��U��i�*��%  �Z��-J�B\)�ȓU�Bc�D�iy�b1�^�_�8��ȓ\�L����&N����S�7:�0X��2_��K�ɝ�dI8�+���_�8\��t_��"���KQT��2�
�|rf���*i�IP �Ά|Ӗ�2�nb� ���t�I¥P,l��B��\6)L��0�D�(�1tRR����YU� �����y���w��E�Be��N@�q�ȓ<Q��aS�Jf�4��U�"���k���3{&5,!��x��(D��ʇ�U A���B�"A�c/� ��*D�l��� d�
������8nq���<D� ��銣30~p�'�#+��D�9D�@YE;^��k��HS��/5D�P@��&,��y���1,���WA(D���	�S�� 󥄵y1�U�`9D�dC�h�`قLݡ�9x�	=D��DM�+'�T�Y�$ �|L�z�*OD�'�&bѠ�ρ-l|�,�d"O� ��P��t�D�G͇!"O��J3�>&�����Y*����"O��hVfT-y#|(�U�  d
�b�ajX����'w�H��Z�\�<-��2Yn�{	�'�&њ'ˍ~��<��m[^�0�X�'�<��Z�!��lۤLH�S�v�{�'�hBR�\��ݣ�nѐKL�p9	�'�F-�a�F�9V5��ˇ�:�@�	�'�J\��$��%4���*�1!��2	�'��`²�
�%?6pxIN<hl[�'Bz���%��6oZM�Z�/[��K�'�����g�D�&��E��Q��$��'r�a�,ԂW>���g��A��pr�'N�eK����P�6<ԣ (K|�
�'�y�d��-E�T�S$ �-H�.���'�.%�d�ȟ�ܸ����r��u�
�'���:W��3]� � �k����K
�'AT�K���l�"  R]�\ۢ�B�'��cU�	�n����юD� �Z���'b+�@W��!T��4i�&G�-D� �3)�?/�,Ii � �^��x��<D����Q����c��qL��#e$D�|�ǚ&g�� �B���Љ+��1T�p�U,�i,D�z'��+޸y��'�:��	1Q0����VR���`�H��U[Z���G}B�Õ�'�PЄA� ��E{҆�Q�v�d��I�'�~=p�#Ċ��tX�Kr���?4��a4-��{�����
��_Pԁnڱ:��q9 o\R�R%�+
:Q|jG�\cʨ�H�'̉0V ��4"�.XNt�#�'��M9��N��2�[a�L��2i��*R��T�!��8���ÀO���d����'8�S�	d�\���Иy=2ٍ�d�2U&�y��B`����dE�Z�H��L�"�
�X�Z�Bq���T�\�D�	@+�}#�O8�9���/ih�Z/
<9����?�|E�p��yS��Qwm^&���s�V�0f9�g�^w��u�Qϙ�y�ε�g#�#Vz)
Bf�1t��C�	$:L��)D�|��h86�]�RE���f�VP�w��bs�MKU�&>K��1&�}��|f'�P�7FD؈	��6w�-Ѡ�Z�A=����$@9i[4d�=��YqF =P��E���E�4�t���"m�sUo�J��N�?��QiR� ?U��c��#�]�<Z��偛A�\|z�#��@\Y�-��da��$P���4� /Es%�a����a��18k�9p�
���<�I�oU��=���C����g#�����R+&!˞Ʀ��BC�3
��D��	U�f��`�^v%$d(�@�O���Uk?	���G+����9���^(|h@T�!�yr�ʚB]�ə���O,r�q��ٙkr��T\�Md�����6�gK�FZ����&.K&d�)C�؛�y�k��F�����ן<�$Ma�/����>��&��l{f�[�Y��P�ί@PT��I7Һ��N[���ځDħhH�PI��ڎ]��(  �-J1OZ�F��8�HBMX���I0��P(�!s�ȟ	x�vL	OۆXU�a�P��b��	'�	"�9G\���U�*��u��bX")-j�{�y�B�"(/h��O��d`Z�j�~���0/gtY(�i�
Xs���>LLQf̯
�:	�) 5G�@�Ba��dT����(� �� a�D!|l�pנ�'O�R!ċO����N��):�W�3�	�r(
����v�t9J �٬G;"�2�‟8z�s��֡ ��r���v/�ӇP�u�f��X�C1(��@�N!<k�@N�6$XU)���>0i��T�A3�p<iu%\�ʸIPJҋ¶�Xǫ�$������Kܕ0ଚ�t�Ќz�`X]�%����	ʢ�P�M(&���%r?Y6-��T��C�k�0�ʤw
-JKFP�>�d+R�\YKЬq�Ҭê�(N�,)aI55¾yYV�'{o^�#G�Q�C�B��K�g�$i�Ǧ�=t�� Ԫĺ�~)�<5*����&�)�q�>�b�@���怒�,]�3��Hg�B/%
�T�𫎩:�ܭcJ�p�6�R��J���L��3���N �x\@�x1�{�L}�bkT�b�����'�T`��˕%/�R�hZ>�<�'��Pc
�bl��?����EO$
q�4ՆA+#�H�.9HLA�g�<J�J� e�V�)T�.t"U���"�=s���)3� Ū�IA�cP�1���[�e��#?�U��K4���ڜ4��D�|�t��4h�kr.H X�Z���n��C�m˶�Y;"�����~�4h��7m���Z�� �z(k����q{7mQ)��'��Q����^����@�[h��V�\5F�@=ء(��VO�@��ʹ&&��U�T<�@0U�ɖK+�`[���*Y�X�k!O�O�`��b�t�禑[�JIg��1 ����(�����@��@&�Y�C�t�0 S+>���ܴ�V���(X2eu������3y6�ʠ�R�x����g`�..S~�$S.=8m��)�xF�g�'�(�0��:_�b|8�Q#B|Us��F 2��%���2��V7q�(� �һ\�nh(!)��FnyK���D��y�Ø�6���"����E�n��#>�b��� 2?<Z7I�8gy�� >�QN!kL,X�n�$H�%ᆥ�=�1�E 0���R�kS.����!iH @nM D"�ҝ�����90ʡ16FۈQ�� ��f�����*tp���M��́��G2T�3Ս�C�0�`�����K�kB�Vך(��%�Z��I=5��Q�B�z�?}cƫ��OPV�����m�DD�-�<Q���;-~��B�aV6_׌�B IҖP�Ԉ���*�S�	`h�sBn�h�lL��Ń L�x��O�H�$�ڝ.
y��?#<�N��}Z�Qp��0Ph�agP1-��7��^� SG=z=�OdT�L��H�I��
�c�Na  � �P ��̆{J�MT 8�牆z촙R�-ԇ���S�o�b�+�#�`9*F�Q��2���a���)sR�֢`"�!�h��j�<:K�On%"���JӐ$��T����h������>��2��	#o��١�Ѱ" (��K@�e�x�T�S�`i(9�T�R�I�@a3N�MD<�0�&��Iw.�4<O�a�d��ah1���N�~���)b\ 7�@��R����8�7J�a'�R��T),��iS�0{���V✠6�D����y׫[)Q3f���K�D�����>�M#
ƍG`��3����DS�9�&Pp��u��!�+8K� ��� *��	�'�A�H��d�O� ` ��~��)$��;K�:���M�(�>d�n�;CP&|�`���Ue���䐔:8+B,ԛ3	���I
���1���J2H �q#'ɕ,����A�[�4�|a����4t�x�R	���P�'O
�a3W?�*֪/�0Z�ȉ�8`��G4�I��&�Y�Y(�V����!"�d����C�U������R�^�ȨŢE�X���˃T�8ṅaJ�_%J��1��O�0`��<)�+͕��`U�G	X�:�3�%@��tP@�S�n��e�B�;nrhrt���hM?Ѹ�w"RcV���?Y�ZP��~��DI#b�d��q�C�Q( ߨ���(,ON���RG�����[�>ѳ\��ҁF�J��b`��_�4��$��l���ED!�`"���K�&�h�*�0��Y uM9p�=xd�H� <P�s�'�(
�d��%V���.�L��@K$ˋ�~T.4�BiVh}$$�4�H�A��̫7�5.�n��v'�H��L[�+
��?�bI6����;��L-%|ղ6cT��b�� e)���I�G��*�T���ێU]d�J0iKaTh�:���P&иA��&Xx�h�'��F����e���M��(��	�E�P�;!��=L�zw����s�ԿH��#`D,v�B�yP�?G�V�3��$��R%C;E�^��b�D�A�N(X�� R:�k�Ȕ�(�^� �oŰ<�c��=Q=�-��kXyh�Y)>� �#�Ø�7�!�F�����S�P9�9H0�YjZI0��X*?�"�{�"��.��TA6��9G;���N̥��=1���Ε���E�&r�2F�$P�:x2֬��`���bD�-b��E�̓'b�`q1�I�.E#~�&螤P�>p:�����Q]$y8��I��ł�G�'�O� ����X��X�Pk�&��7K֟��iB�7vx�w�.`�bL�`�l�64:c��B��"�j$���)2�d�/Nд��&�B�h������4k���$-K�m�.\�f�>E����j��|;�"��-~�#T� 8R�`a,��f%&m��'�A��P�cEN8� kg�:� ��A�'�8�O�<��<�BO��1G%�'	s$��V�Q�|����2�L*Y����͞g���;�M
�J8Ĩ"�'�H�!#h^H��- ��^�c0�*�OБs0
�?Q�z�s��R�:n�kr�ݸ�1��y��!W�P�
��!����"O����9{�8��ʋ�x�P94�P<@ڰ��AX����WK��En1����G��Xj��9<�\¢� /s���'�Pr�	�LI�� Q��!���!��9ZЙ$$M�~ޠ(��<⵱��%O<�vm�?�Q�����HxP� A��M+�Ǘ!R5@@݉�據czt1�`a�±�P���־}Cd�Ý~rYy�i_��!�-�F5:���э0~��œ�C�N؉�����lxd�"\40��D�;�l�` NB?b�K%�G�@؁����``TC�>"ZďU�_�*�s����艋b�<s �lZ?W�r���/�.L%JT�����s�[g�=i���2��t�(9��0�ݐ t��Y`�ÎH����#K���|rP�#?�����\�����	ʖez4ɍ8_�4 ���
I`<� ,ؤB��`���J �P�Р$ 
Ϟij4��9]�4豉5%A����K=Z�1�TMkb������E�#�(Є�I�\<�dn�Zw�eY3@M�R�����!N�����G��BMX���eAC�M�����5�`�PeɸX$Ђd�������dm� @����JU£?�7����	b�w� IY�kA� 	!�ݕ_�Z}rA��&_��@$!E�y���T���U�嫐�C�5
Z�NY2��$Z��h�f�"S�I��Ҥ\�:��!�Ȥ��]�2�����m#Q�U�&#ӧZ�.���I&%`` zu�(5D�*͝7Sf�Vg"%�^�:�aT�e��a%���iJ��+Wa8�*5�Z���Y�1��+f|@��� Cֲ�����V�
�"���=��)b�-�+<�8aO��`wTřSn�"F߸����i�)�3� 7mu��r@ "_�h�XZl�6;�P!���Y�r$)��Dҁ}�zp22��. Lz�k���!�����$""*�*�$�:2�0*���}�nTb�",Ej�C�.��� ���.��r��d�`!V�J��tS�I��uMJ<8gOɖ��� ��kA.=��H��!��O�
ߨ���a�/cB�@X��]�x�*�@�mJr�Z��ʆP����٦��1A�-dL�d �4\��}z�my�	�s�N�~���q��������1UD��" q��g_0:����'�ؘUI� B Rhp�BL^�]0 H@��G��Z�iwύ#��i�% v�rP� �w����Y6
DH����	�6��X�`�;N*Z�т/��D ���<^����.���0��0��t�3 9K#J�ᒏ_	�y�i��49䐚&���96f$K���8��hR�c)i@���3�4�(��O>���B$u�Nd�s�,f:��P�77�*@B���?�Y��&���}+ө&p�VH��7/`2��O�V�r�'O 1����.6����n,3r�<�A0�'2*Zp͂;Vx\Q�I�Zbhh��"��rIr�)��.,!cƆ6y$t$y7FGf:�A�S1c�O��P�C"��!b���f�$� T�	��
ؠ��wE-{���A�|RcE,||����%Teb�9�Эʙ}>D��Ǜ_L�Y挫tE^<Ą�>-�ғ%[�$�ܤj7�E3DGnģ`B#;S���Jͪv@T,䤧~�֒VoP�rW���@��XQ�HL�A�+``]�� 	�Q�y95kĖm�R�F��� �AX�P�LD�qFѪgr}���X�!��T�J]BfAեY��𡵀�@�"�E
��bNi�%��Y�)Gy���9g�r ݝe�� A�_�3�k�!���&��a�����9e�42�M�a��&�?�"KI/;�"��#�#yӚM�g䖪D�������.:�����+��l�<�[�T \B��2m�Wt��aQ
Q%S��$r`��;&�
��'	�U:uKΣ��'1)^�V�Dde[�$�s�,͓�%�.,F����� t�<�HA� �X���C�)�/�~y���ƖsN�����8p���h��O��x�����A��͏G��ŉd�O�P��Ptq��X�lޝL��l�����1w��D��Ca �?o$���*�=Z��Q�#a^2Jh/�Ј��üY��q�ӡ_�X��f�x�"��%�[�8�{� ̲x��]����>r����3Ț%}�� ��
�&iZf�w�Ⱦ;��q�WM�}��}���D*-�@1�p	��;�pԱ��+h�8����U ��`�3OF�]Wb��&R9(�D1�)J;�~Щ��+��	O5�Z��B��\ش�c�ؿ&���C�Ĩ,��H���DԖO]�tвF͝G��I�`�R��$�C�{@Za B��GER���(ԭL�"ذ7��&������Z��>&�"(Y� N�#�r�2�j��i�85"҉�94��p�GܦL�2-�O�5��o�I�TE���BC6�+��'�����ɔ�d�Xyr$-�d�xX�!�DWޔ�Ԍ�TۈM(O�TX	��(I��Xim`�bl���E�Tд�,�Rלm�9q��D�1n�&Mi"xhtoV[��S7���`FE�0�)%���u7�92� ��P��HiBQ��ݩd
�(ck�c���8��%��z��5��Y(V��a.�"�+b�<x�<�I�c��3�g!I�~��務�pL䄑�пVr4%���<]���+g$��/��+��S�O�~�uK�uFꐉ�P?Uv 1Z�&��U$˳]ä�aw'3r
!�TC�YM�(�%�D�
[J� ��웟s}���He��bj��j��(�l	�p0��:զ�.'��]�.�!Ƅ8Q��Y-Ta��r*�&h��xB,Ht4��j�wD4����a� �e�I�Mj�y�O�8�˙�|�ʠ���I��6�|�'HO'W�0�(3NII�4��vS=��|zeN�7� ����j�6���O'U�"�x�nH�J�<��R?{��`J%��3E����5F�
�:8��,�|s@�hɚ^`���C�����W>�	� ��>K׋�W�	�p&ϼ|���+Q��a�b}˕���
k���W�ؼ$�I ��ֵY��� ������<�0f�<3�	$�
�\�4�JP�&¾aa�#�F)�d�E!΃m��ZR�?�,y��KZ�,�V*�.�u���3@�#��W3k�� �� J1}ތ�c��4�d�6oK�~1Of�f�Kz�<�g-<t+��dP7̈́�b6��>����.Y�X�a;�숪g�^u������Oς�Z���58���QX���3ྙC���91�L��-Q|��ra�M�T�Z�
��y�DF<�e5�}�-��K��B&�t�ލSVC_� �m�4�3*h�8+��\:f1�}�I6J���S0t�څ[F���-����Su��:4�XXؕ@�sld�!Q�O֩�bB/��'clҡ	�B�>��(H";�,A!�LL]�CӇ�j���Ӯ�ԟ�ɥ.z;v2e$?�O�,GI��H�,=c�X�nq���Q�q�N���iҲw�����J!�#�/1���ӌx��kÄ�4��\��Ñ�"�<�<"u$S'�x��V�lbd�t�"q��i������:�Z�ѳD�ΥD�`�kF�6����O��x�ҳ0B�ޜC�*�)��'n̩R5�TD>��"D�`�nH$�?B3:5ˀO!?��ȑ|�vT*�{^��~�$O	%�,�0��;��ع��|�<9�	�F`B9zV�0��y�b;`�jPp$�����Ŏ���c>c�4(RGʠ<T틂B�K&����6��E�Z��p�Wf�^'�5�#d��$���ՊI�}f�I��	 p���ߏl�.4"BjƔ7`��$^��>rGLŐ*O��:2�5�T�i� $���V"O
�����cs��Qo�,�-�d�D�,�)��{��ԋP�U�`��㜧Z`��d��y�!�d�y �H�=k�䔓'nʸ�y2+�x-l\˒�ѣ�`h�o�y�J��T�1!��e ���1	K0�y�[�МD�#o��\��R�Έ��y���|Ȳ���ʐo�8R׆�yb�J�8"0`J/Y_R3���0�y��O�.O��(u�įgs�Ic�`��y�	�\��
)]�tIB#����y���!z�i#���%��B)ؚ�y2�M�<�
&�32�]k��_��yRoǰ��y�ꁺ���V���y��J0fB�|0�!EjD��^��y$H���`��I�U����,S��ybN��m����@͖9�1\�y��>p	�1k�-��Pp�9d�R�y2�E'.�^P�Q��&Hr� X$����y�M��-�xQ;��E�ޠA�A���y�H4�:�[����?�H��,E!�y"eP�&)r�х%�0~�ܱ�K�y
� �qS�R���X"��ܲ��8R�"O�!i#m[��|�d�	Us<`2"Or`)F Z�X
g�5dd!Q�"Oj�q�!�k�>(�@C�/+��q�c"O\q!]=�r��B�S���(�"O�lcaN��9(�%�Fa	�
 �"O�p���sUB��FŎ�j%3�"O��;'(]�}� #C�F
4���"O��i��4UR��3G�խ�n�"OBaC�_�|1^�!�8r�(�"O�b�䁕�$X�K(�ч"O��@&T��xG��"$�*"O�5���E��p&ʏ�W�9��"O�H�&m�*i�*��D�"O��c��!},8�ߔ`�"�$"O�D�uD�J�}!fmG;,A�	�"O4�(�&�c�lX��*�`q�A"OV��L2A��s0�Q�'�he�R"O,Ѣ�ֿ}�JLZ����4��"OP��B���X�w�m��%��"OH(Z��� MT��u��> 2"��"Ol���*L�<���9@����"OtH�A]��A#S�ۖZt�|��"O��=y�u��^ P���T"Ov�:P�^�<���jF��(��`� "O�pC��X�0��L��cmU��"O���mC }����jYl��2"Ob���M��:	ՊG���4JfIz3�'��D�5���[��$1%��� 5��h���ȓ.xH�c�K�(�����{1}F{��˄Q��2i��'G�j����'mf�e��%��2�XY��'$qrWh �b�� ���%��l�!O�� ����Մ%��`R�0���@��Zz =X�@��<�dЕ�QF�<�Ά�/��a�O�'S�h�+Q�j₏^{�hd
����4��Y��}����?���<xU��'Ė"?���+1.JZ�'��]��o�П���o�,ax��so�]F��Q!@��}z� ��>j���U��������Q؞���#ڣSM�i�w�O�H:��P���z�,K=R||�P�!�hUL`���P+"ú��׈'�`�FE���M��E9g� d����2K�B$"O� �e�S�6u�R���՘G��0Z J�a���5R0y�]|^� �"�R�4}���ŀg5�H��v͈3j��CuE7^&��8��''���ED�l��$�dNɌ{3�̪��\)�Q[G�M1O���7�L/N@ԡP��4wc�0�T	y4�����T�
�A��e�ܠ�ң�p�ў<��U��Rph����6+��(#��K�Ja3%k��?��!�'�Ң?��&�"W��	����zh:��A��Q�C�
@��(��ú`h*CIc�~@sQHZ�a��UW�LOf"uX�Ʒ�����مp6���Ɠ"oz@c�.��N��ͥe��Bq�KZ�<�A�D���iQr�c�$:1ݕ�@8 j��!4�+V!��V�y��E��myB�f�j�\Լ�Ѵ���D�}��E�&��4�`��X9k��dҚy�fPѲ�؊O2҄�&FG�o(5��Ά�2��ħc�HC3#�
5�
��c�$�\`�f-�Ʌsˀi1��x��ԋp��!�#=IpO�aʬ�r!�پ]E�I �,P��>�v�	�bq�3b��lI�+M8�������:/�AM��U�1O��a���r2��CB�B�`�d�2�%�qX7F�}Oxu�¬ЯZ̬x:��+�h���D��.�ղ���$$���ƜR0
��҅�/��0)` ո=��� M�`qr��*px4�KI|�>�篋���yEh�6��A��]���q�7�ܟT����C��r�܅
!Ϟ~���a�*<��w��*��a��한t�N�H��C���y��������i8���bGU�zY\���� �\`3���&����!��Z�ajpɅ�RY�xa"��az�8����Td;�eM$����1��� ���[)>�P�C�)D��%���e�c�<r�s���z�D�TT�sǤ��Y�yg
ϯ4�A���]2m֪�b��ג�M+,��
�ХC���P��b�AԞ�~�N�oӠ�z��7�iF�H��4��:R���� ��j4��-L1n���O�in����!I�� 3��;Q����6`�d�n�M���td��1LZ��� Z;H����'FB�2��ĩO���P>�<�NΞ)�ت��S%�$�+�$.����B�ʯ_� a�qAq��e�.�*���E��88W�ؤ.���Qw)Sp��|H��ͦY�����k�p� �1'*�G�'l<����5[�Z��TIM�]�F������r���Y�湹emU���|�q�)#��	�/��[�B�Ӂ��� ���O���%-�(w3R�sV,Ɨg~��CV�V�7C�b�܀%��=���`�oٰV��a�O�^��,��\̶�L\�L�(��ݰJ}"��
��­��Ù('�%뤇�8�?���M���~� D�)5鐪^f܉�W�Q)�MS@�D�W���%��	3dypE"6XJ�a�4P�֌{�",	�Tx�� j��#�O�I~q�nQ5y�^���$T�����E�}�'K�?j@R�g�'~��Q�@Ѝ!��hp��$>Y~�J1g��x".̄@�~d򳅖�|��A��"��|`�KF�:Pl�rq���-#�!W�@`!6ںn���PN�08�y���X4j�5��j��o�HpiB�F1%�"ekRK'b_ni˃��� <r(�-S�#��EJFE�5:��Q£0$�&msb�fVv�Ğ#9t��v��;"t�8���P1Fe0��?�$�#!͆;vA��9�lN�(�p����P��v�;TbA6��]{��_�p^�;��E.�1c��$p��Y ��C����F��S�'$1��Q�ۍ6~���@� R]��x��˯*���4 ;�,���Z�3t���������i_�#&IAT�@��l�`U=l;��
�
:�S���q��O� I�.^�uHԉeD�I���2U��ɲ@�I�T�P�8V$�7=��ӗ!FE�ِn���RS�%�T��g����%�pHJ�s�|����U y�yb�
r�z���U�V�L�6)�2�64s�.N?è�7�L�l�0 3L�12���F��|S�\ۆið� +��<b������F�c7BK�W[�M5��T!�YFx�j�8I�����Dw��䣤J:�T��T��*x������$?Y�i���5Ғ͡���L{RP�ӅK[�	͓*�ʁ��Ed�g?�$F��R�h�2�
�B��0cIa�\�P�I�/��	���7����&�
U�|����C��e�e
��jy�xS���
|� `�0��O<h���p@���<ie��7+��E����^":T9���S�TA�R��Zd��uB1�X��S�*��Y�5� X#8dQc�T=U�Dy��NT�u!�Ӳ�RF�bQq��N �p=��'[\��(K�R�x$�O*x���Ɠ|���'I�E���Rg�8Jp$�'� \q�L��.q���	��O#��6h�o��+!
x�ډ�>��޼rk��h����Yj��[�,Ż/a��;��O	B�D�i�"��^5���eL;y[RLhA��2'T���CK�]�����F#|�'�x�1��Ƀ�X��U$�'w:`æl�G�0�ԋX@�\"g�5k�l�q�ɂ��'m��1Y7Z�Y%�\bz�`�F:�(�%C՚Py֑Ig��5�f|���EK��"Q�R/��P��	�_�teTDI+�6]�����nI��iv�%	rjD+N���-Ƨ]nI��A�"b��#� Ė���U�bQB)LOd��\�M�2�R#�ݐ���`��C�]=(�d"A�u��Q�Q�ٌ"r*|�UcR�L'�`Wh٧���x�G��X7RbN�Dņq���aI��|X��B$��'� ������Бr�G%#j���m�z� �S�a���Yʶ��00}^�VF�z0�� X�j h)C�GE0�?6'�gyBǔ�LZ���L�7h��!��pF�t���DA�(S�FJ4Phr!g�.MXc>uJ�;Lo1��)��){���עu��f�#����g�
+�t9*q�!,O����N�A�F��Pd��[N�ش�H.�H9�O��M�U��]����w��J�$�&�.�3G�ta� # �DHb'ݕ*^�8�A�$+a{�+":��E=D�w_'X���`V!EUή��4C_�ze�y���Z	fZPa��I5���7Ɵ&X���pF�Յg��ݪ����<
����; �8�P�D*	���e!��-��S*G� )�F�R�#ܦ��)JK;!�z �T�w9�yҧ�"5��+r�&��Z�	<  � i�枙S����c�ϧ���" �wn�)�I9}��)�^�үџj����j�0�96$��-}r��P�A�ւ��ɦ�n@1�N1<��`�$�<�0�:���㓉3�$J	}r��!w��%\��aRf1�P�Ѯ���T��%� 5��3�!̵�Px�E�"׸�2%�4)b%Q��7��$��>nB�r Jj������[�F��Ӄ��{��`Xs!� xF
p�.^�v�!��L�A��(��g
�i �U�NI}��@yd/ v�H҆B�$3��󉚥2��I� Ivػ��ޫ3"<�[�@��C��6Lx,�T!�jl	3�	�;
��K1�؀L��v���ڍ�pY=����dS�s`���J_�
ӄ�s�
�.k�2m2�4VV��BAڰ~�^��E�v>�p��<*�9�W��Z�vY��n�.�YE����T�!	b6-��8�Ov� �G�^���GnB.����K|�=�%���~�&��"jJ����T��Z����B�.�� 	���3J�5�� �Z�&�1���B(e[���>��'�<U�G�A榍����Q�`��-�)��,�/�=r�,E��/�p`t�e� "���K�i�����k�F��Z��bKɼp�&Q��oN�|�U�,?i��)n�2��hܴs��d1��Wkf��fj���mk���f� (I���m�>ٱ��p��h!�̂�Vid��1٭v@���˼<-� A�F����Rw�]����c���jL��	!6C4E+JNA� 9��
*��%"sd��3M����$���0��!6@<QC��NG�9��J)��9"�Ē
-R�͚�E.�����r$`���1��kA�0j�t��A�����C��L���I���{7Ϗ�N�e��L6L P8��J�<r��"AD�%=��T��bđH���#��ΩG�M�L̷N�"�iS��$ �4�C�E�*61�I>s@�"&���4f�QR�ɒ
7H�!B���4�!��"SϜH�����1~�	�Y<��	Z%쉔_�Lq)s��ߦ=�gb�;C���r�����Y�4���ؒQ�J��Y���1%ǆ� �6�c&d�" 9�	�W|v�sPh��eF\z�P_���5ƾ�yW�
/^GL�+�nP�Yp��u����yb�ļ0�
I�u'ȾRd��F���\H�UK'�ʳKz�4r�	?~��UD�5t"�(��'! ێ��1^B�}�K1Or� b`-�>|��E�޸I<HD#dG����x��n>Njl�����O��`b��*����gIL,r�x��e�|����cҌF6���/�?Y)$��w��U60� ���>����"����IUcS�A9��l�y�Fh�#�[.By$����U&���+�ēM!<�s����P=�U�5�Oq�0��d��6�y"���Y��yZM%�P�k��.�F,�dY�3Z�	�	��4e�b��#IĒ�D!�Z�c��	H�9�<p7�ѱ^�(qs��P/�� �S���tf���6D�
)��I�?� ��P�[�8eC��y� �9���0-u�)����<~408���2)Y��B皑�`�� ��3�ɕ,
���hÄ-Aԁ���2�@<��`Q�O�4L�B��5@�rCl�3K��T�(Kơ��-����@��d�CєE-u)���B�.J4m�7B:EExRG#*�J��l��"�}��z� @rWO̙X&���!8(Y��m��r�иٕ�C�z����"1�i <�$�c���"�!�j� �hs5�?:c X�Æ�^�;g,D�C��d��!�1Nv�
���n}�؈�T�E�\�8$� }��G.W���� )��@��,���Z�t�d+��� �V�t,� |���`~��ꅠK��go��KF�L��<\�� 0��}�ꄁ��nƤ��#�A����O�!HN�6��=_���� |
���M\©`��W;A><]pqaæ��l�%�4f�K4c��&p�(�Bw
Fjӕ#<n��a��5.Z`I�� #e�2M�C���2AÀ���Bu:�Jҗ'6~��ٴ��IO�k�jA'�� MC>����0M�0�F+�u5 ���D�&#\�X���#||��nF�Nz�0� V�6��ԩuɑ��h��D�5 p�{+�[�1�I?�bw��=�,��|Z�@R/+\pg�ި/Фu�q
�K�iѰ�x%K���bq�"9P�TU��͊W�P8zp)W�^�����;cʔ}�򅝃Z��U�[D|�kfl�*U�1���3^��2_��3�[e��-H�[+D�R�H.�^��
\;G��� �U�$]��2 $�҉�!*B�B՟�y%N]#
�JI��MX��}����_k��X�G4I�N���K�b}z�f���ll�T
\��c�@�Lb�0�逪L���A�ģY�������
���4j�.�D$���~�(�	@+L��ɲ!\>}`�`�1�*��OM�=} @��M�S�Q@s�S
#��➤)��|l4�A��j�<�20� )pNx�H�}��@���,�!/��:! (Sw��=Ts��j������S8$�佪��: ���'Ta��#%�>4���2�S�E�\t�Oh]��F�v���*͜D~�ȧ�'cj`��Q�O��t��!�\a!֌̠Q�����;{Z� ��`��B%�A s���Gԋ��)(T�#�/�޼��+��8�m��7���2a�4�̘���P!�Ѐzé�0-�X	���k��ӛ`Y6 �r��R��Ac�!*�2��m��Z�=���ڵD��4�rOÝO�,5���/��u������'��a;��&s���m�%O��y2	��ǮLz�/����H�$I@�?�a�
$w���1͌'H��AbiұŠ\*�!�}9�2A�&Rda�!�Я	��'c,B�a*�yQ�J�MB�&�4
 �p!{X�h�ǃ�D(L����
k6���O�(b1
�%/�|3	�.U6����#�P����7��y̧?�p�E�n�jBA�A �h��'��� 2���wgX�7b�>��`��)@��b���4��	��L��ϨD*ؠ P 	�I쁁Pά|"B��"�2-�w��9Bd)˞W��H�B�4K%R��wiY!A���1Q�')�]��b����d�b���B�.3L|�@�)9a I�2�G�K-z�b@�D'	�䔺c(�`��t��7Jb���$bQ�Pe�a���Aܘ���� <�X�lT%:�*$��i�	%2�t�(���nڢ����U-�&Ӛ���ָsY2�9��O�_�X4ߎ̲��Vx̓ ݆؊ �׺vS ��`��?�%�5"D�e��G߶n_�\Q�B�R��l޸ࡒL��?�v$����ܳ�J�/�ZDA�O!�\�e�X0`W�7޶P����N��Xl8�M�I�'�P���IߘXpb	��щ.�R�y˽Z����g�Dha7ꏀT����ό,��'Y�݊�w�x�C֠g1v�A�[����D!L %=bW��t���ÞV�q��'K&h+#̈�J�ter��ާ}b��d�6ņ���&(�a*qGǉ��g�ɶ3��e����I��D��o�Q�0ɉsKX�e�4�	T�����M�} ��2KTw�8������Q�d�� 
�V�VU@��Y�
�fq 3��=d���_*^�x�M�>
4E9�g�-n�GR�	�WU����Q�i��EK$<��i
Q��}�uk)���qU��t����q>��GsVe��`�X���ݶ}}D�@�&�ʣ��i�����-/�'b��q��u�b��3󲼆ȓQP���	}*�\���c�	"e��:B���--�kը0�3扄7���&C�Vn�&
J&"�LBቛP�-)P�T�@�P���;6Z
}i�B� �F�(�HU_X��#p��-*� ��F �`�x�T�%,O$I(�퀼Q�
(�(O8\�ǧ�᥆Fx�@����y�Y�}�4�Z��L4�~�q�����'�|�Q��j�S�'w�zl��ʌ�[��GB�.�\�� |b`B�iܶ-zչ�dC��ȓ(��Z���hѩnÌ>�j��ȓc���р�	1�8��T�C�6fDt�ȓ"�!+ )�8w���`�H_Hf\��bֆI����9^����#G�7b ��ȓ�葖!\�$ ��-x\��ȓ.
�����Bq��z��ҭ!��0�ȓ/���;\K(1��,$�,͇ȓ!�2%s5�����y �޷2���w_��xu�P���"֪z:>X��)�����ǝ\g�`�b��" w�����1k'5�h�8 j��d����m�Ɯ�#���ғE�!>"�І�L4��P[�P��!���E����j�^5�eڟ$+P���D�&��%��S�? Q)��Q"t�:LI)	��P�""O�́��U�At�шԡH�i�"O"IXW 0L�(r�J�26~\�"O�	ҭ��5��d �	�V̴R"O�]µe�Z1dEf
�M�8CG"O��{c#�e\)�E�Ig�P-�C"OTY���X�> �D�A��
�"O� ��
�5�e
��ķ{���"O̭��fT�8
��b�$��A4"O��Q��Z'��`�!L�T���"O�2��T�a��@ �=�,�C�I�4WV�a��'kve1BK��t\�4�γw~�U��'�V�!!�dc> �'�̧s�D���'����q	M�?i�H!"�f�D����0�FȔ"É�����BG�P�^������]�{�թ�CL�t�
Q�%..�'�'��ĀT:H�t-p�(�%R�B�@\�J��T�|R,*�0|sI�v�dh�zvf���^�K>qfF��\ń�S�=�x�@�R���
@��]�$�".�1��ƍ��S�O+𴰇L�];n(
�Eѝ
����'�ƴХ�&�)�'� *0AA�*@� ��G*��)��`I �O�?YJc��)Cz��W�ͤh��U����%��'��0��S�N,�E����:?��LR@�\�~�~�,(w�SJ�'k�-��*��,��	�Ah��q�|eI�H����ا�Ok �P��FHHyab�aH�\h�'�21�Pb*�)�'T'th�c����a\�v��Ceb�697"c����C-3��솾w8h!�nE�=b��SA�O#�V�jزjT�,��Y�T��=�@�G	+�O�Y��B��S}U������'�b��R�O<�G�i�8�>E��J�'>�^��oX)�̛qk�@wȜ�#�E�Q��1���<��	d��i>�w���J����t�n��7R�y"��a�T����:f6T�����	�8��s��B�<9�H�Ozҙ9�Ú�7���(��C�V���O�����&h,\4��Z$2��U��
,Ln`E���#+ �A*���0|�7+�ը�CÌ�cc�7J��d!
`�Z�tcj��e�'��@(	ç]��yH�,Ƣ #6@��h�9QW8�E��D�`( BC����S�O� kh�0���a��7.2�Z��H2f�d+��k��s�,���$:��4�bd�1z��9+��6D�(+��6[�`rR�|�8��c-:D�d�VJ un���%.E�8��(J�:D���0�_�F���p%K�s�� ��6D���A(˯]"�XIUfD?UG����5D��B&�.s�\�x� ���]z�I4D�h��铢o�Q#UG�#~j1ʗ"3D� C6#�!V�D��↊�$�>I��c/D��j��S��L�i�:�� `#.D��]��-��K�f�Տ(�rB䉮%\(��W��K͖�b��� �HB��"6�VLJ�d�$>y&�*s'=a�C�IU�ej���x��ra
9{0C�I�jI������-W}�4:�Z�w�C�@�����U�]Y� �� ��1��C�%4�����d �K"�4	�.�
;)C䉅5ռq���A����qmG�>J8B�I�f%�Őf���me6pK!:�jB���x@x ��s�pR3�#9�@B�n70�鍎Z��825��%hh&B�ɜB�ůׁF-�5�ύ�.����-[:|��G�ňM�t#�;�!�$��_`����Aڕt�|�ā�E�!�B�y��ƕ[�p堓A�7�!򴔹2�ɜ�"� �vd��P�'B��00m�4x}�M��Q�v�2h�	�'r�*Qد#z�5	w�WixV`z	�'�^%y�NJ�[R��Yƕ�^�\E�	�'[p�
A��n�~��D�,OW�xa	��� H�)�NW�o�М����81;�#�"O�S���/%v�Y�əp1Nl�a"O��s�bʈK�P�w��bI�8k�"O"��ގp�@e���ξV<�m��"O�E���"+�Uz Eá1Ƙ�"O0�z����x�tр���T�(���"O�q��KBi���	��D�>��MPr"OL�ڵ��=b���� ~��)[`"O�XV��'B��f��XNr�"Oh��c�B�3�Y+r��-BU�#p"O|	����B��I��P�1��RE"O4%�ȁ(S�d�k�ڠ�:���"Oj9�c����A7_�Y�a"O�$ ��ݍJ�E���ߣ�.��"OX8�&ףe�J��Wχ�uײh" "O�$�G`U�t��0��3Y�D`Q�"O0yZ���Yi�D�s"�!�����"O��xS匃$��M�Հ�fep�A"O:9*��_U$��#Ʌ%�<p1"O��ȵD	�؊A���)xF,H�"Oh�k�L�)0�0� ɀw�H�"O�	#�J,���s��:Z�ؽ@�"O��R��V@�D!��0i�-��"O��$$ϊD���TO
 �r�Z�"OX8��M8%1x� ��ѭ"�lHF"O�EY��/
<ҥJ @#;$��إ"O��A��z�zx�#���A)��6"O���&Đ�B�Z4�e��'M	f��q"OT,P��&�9�񪁅T��q"O�a v�5��aCȞ K�$��"O�Űr��X�ڝY �0j^��"O�<�����cԕL�`9��"O  �"	Ĥy��W��);�v��"On��B��{N�0
f��n�B]�"O̘*P�1��s�*
�Y��"OR�sTlÆ;�>TXt�
�zu`S"O|�q�*c��`	���1l�]��"Ot8���
�-	F*� M2W��p"Ovu�����J��OVD���"O�(1�A3.%���V���P�0"Od�sD��b����L�w���"O����g;�a��ʛY��H�"O�x��'��H���/$�����W�#�!�
M�����ۼB�:��F�< �!�M�gw�,��#>R^� �nJ�g�!�$SJ&z�kB&A.@�l �P�W�!�$�]�j��N�,:�)���U�!��Ŧv�z���R$Y���t�!�� Z5�Iٶf�V�4p��r�!��($�,�R%źmy�	��E	9,!�dC� ���/�p�2���$D!�3ۨ�Z`H�g�x�pC��!`_!�DܧE�^)�W�G��Rb�(-!�$K)O�q�*�
�(��`�
$!�D֯8��ඏ�1U���c�.�@!�d����H@'�	~���RT�!��ߒ��"�՚tb�l��m	�!�$4n6.Չ���(\�^ݫ�13�!�dܲ�x�a��X���Uk ��!����%f��&h��`�DI7�!򄄩�B3w(�:NzL�B�N�!�B�*{�Lp�� p���
�!�D8ў�KA���<��o�!���,}� b���8&A�K�վmt!�� �莿A�9
Cm�@���$"Ov���d�*j��N��N`R"O޸�Q��t0�q�w��O�l�""O���+�]�X!�*Uy�*���"O<����� c:�C��;�:�	�"O$�� E��(��ӱ͕:r�,���"O��sIí8ɰ�Ȅ��a���x�"O�uCW�Z�m|�C�͉x�}�g"Onax�C�g�>-�k@,Q�l� "O�<��`K�ޒ幁�!P�*�"O����C�d�ƹ��*�"=�Ԝ2V"O���/5"�Q�0�(��p��"O��r�f5JF��&�=kkdA�"O�x��Dɀ�ӓ��kn�z�"OL!jg_P�d�	5�Ta�YRD"O��K�E"�>��ߊnR�Y�a"Oh��@��	#vK35#⼣v"O8옧�H�Tܼ��OH�D���"O��F N��Z�6L�|�B��"O𙻂�8@b��eKI�d�=i�"O��Z�O�U���R����k݆ ��"O�h���L�������%d��*V"O��J�h/V�!E+��*���"O�m�F�?%xl4�)��>+�dz "O^���Y��V�
�ԁy�"OL����*#� &@�O��4�v"OP�0G�I��ia#-�(8O�A٦"O��I�<�\���V:\M���s"O�m��GU�s�D���(N���"O� C��s�t͒!�C�[��͐"O�m�W-�P�>����΋r��"O�P���� d���r�F�[�"O�p�D�k�.����؈U���z�"O8�h��$z�@iֳn �G"O���"��'�
�2��2�\+D"O"��DL] 0�E�@-&x��w"O�J����m�<��l��r���"OE"���'Dd����R� ��3�"O9��J�'y]:�����74��1
�"O(}R�KщrZ~�S�f�*5����C"Ob���ͥw6������oE"�
�"ON���/XPv��
g8���"O��"/A2O��������m$��R"O�%;��X9"����噼T%i�"OP�(��[5s�N���]�@#�� w"O�����v�x-Rbjă;�`��"O���Ŧ�)LH��T��	U�R�Y`"O� A��<�>��%�L/#�rȉ�"Oa�P�-4���1f��7�4ʠ"OF]��
$��`0��>q!BƐ@�<!@�R�<�a�"藨]�&11!�Q�<�_3\�)���R;��]k�
p�<9��B�̠o�<��!h�Q�<�C���7�z�� �ʹk���x��L�<ѧd��ި%��M;n�*��&�O�<)�G�
-{N����ʡt����t�GH�<�0 ����
bcRn��yi7��[�<�0�S0\��Z��ڗ!��ܻd`�n�<�0ƍ�(�jya�QB���u�<I��V1{�i�'�ۚF�l�V*�G�<����v�i���(��J��N�<���	2�pS�Ìj��FE�<Ѳ��0�� �)���B́E�OA�<��g����K$�p�֙q�n�@�<� ����L�mcN�x��V�5� ̐�"Oq�e';}�zX�d��q����"O-Jc镡i��#U-G�A~ڸ��"O�� d.���#!�W8Ctx��"Of(�TI� N�a��k�&15pM�5"O���L&�4�aT����y"O�Az�E�<p�R*^���c�"O$ԋ���=���r�A�v}����"O�19f��9�\����\/"mL�v"O���a���<��9wf�&d:=`�"O�aH0���6|]�ʆ"O
��� 08\���ڹus��h�"O�M�6Dذ �Z��K�17>�"�"O�X�F�:.�*%����4��"O`��3�T	%�"�P!�ʎj�P�0g"O2�b%J*RX\�rǯ҅'��p�"On�k�c K���#�o��AR "OE���׳V�F�Ԅ^7Z7č�"O�0ҥ��L� 2�N݄D7$!H�"OГW�	7#�2r�k@/]%!i�"O��b��QN��qÌ�%KB1�yr�e�z�q�mԮc��1IG��y�eJ9)���ԏUB��y���yɞ"P�,�QWj�*H��`(U.ҽ�y�fuPI��V�>T���U�԰�y"��h��ZD#.5�4��u	� �yrEJ?3��g	Q�*�0�5d���y��U�[܍`a��|*��yr.Z��Ȉs�a�l�'hF��yB��EE`k�L�-y�y�&�6�y���B����l\� �0��O*�y&G�*<�1D� ƾ]�&���yb^�
0����͙��D�9�a�y�+�y�Ny�q�E�yt=bū�-�y�"�0^]Nȫ�%��z�\�1%�R��yb�m�z���rׂ1��G��y��*x���So�%l.�h��=�yR׍R�XHsG�G2\�8���)�'�U��W��0z�L�/yK��
�'��	�ح?Ȫ��$(�8x�ZqZ	�')&Qs   ��(��KT�c	�}�ǭ�y2��/�N���*�&EY⍈W(Ċ�yRiW�$_B͘7EZ?� }�v�R�yB� 5��#�HI6,ؽx�Mӂ�ybG�D�<Ҩ+�8�`A䂶�y��sY�L�c,6xD�I���y2��e*����̪~�j�����y
� Z���B��s*(   c  W  �  "  G(  �.  5  S;  s<   Ĵ���	����Zv)���P��@_zX�B�W4S���y��ƕ	#�e�H<!����іS�E�aYҋ�k�<�%�
I��Br""�.ٺ�C$Z�h�����,5���m��e��
��Y�@<j�Y2�~y�
F*F�y���J!G�}[�璛ynơK!F5�V��1�Ҭ��9���~\�q�Gv.*όl3�X�%��a�4��.���0p.(�j�.�4�Q���>�x����$u���(3�'���'�BS>I���cr���+M���f��fn��C�rZ��	��j6�E[Zw��Pf���3M<)Т�+ vkUF��f!B�ö댯0dİ3gY�Tr���f@�E�0�O��Y0��7�$�0'����C���CpY�RΛ��'/�|h`�'�l���|�'�l�]���p��Y&&gv�@���Q��Ȁ��F��M��'W����͞�0�V!��hJ	r�Z��4?�&j�,�����=�I�?-�S_�$n tj�,q��D�bw#�Ta|�p$^�a�"�'�'�����	�|r����%ܙ3���T���&߷3T��#Cѧ$>p� K%C���e�]ȣ<y"�=P0@u�ģ,�d�	(w0����^� ���Jҥ]��X[䥄�{�2�<�g*����q��U;�I��LB�iX\j����M���@�'�4�	 L��İ�*Ųj����'��1Cť�� �Ș �ϭg~�QQ�OZPo�̟��'2J��7��~b�����:I�!AuHڭ���Ƿ�M㖊��?	���?y���Z��j�E�
�H4�퀒\���C썚Y֦,�4i�$�P�R~	*� ʓzo�h��cݿz3�q���`���̱_��)�Cm�-<�b�qFB{��(B�1�!����;�M[��)6|^b��BZ�4_ZBC�8��Q��\ҕ͍?_�X��lJ�/�d�(�$�O`4�'��(b`I
�F����C]'YKb8ٯO��[���q�	ȟ8�Od�x9��'��Ak���&yQ�-R��S�!��7��h�V\�"퇪U�̫1��	����F�+��b>}�c��T�){���]��"��	����bV�`n��ڤn�:D�8$�0H�)5\��iǖB� �0��X�Dcl�Kp)Ĕ/����sZ��vӞ����'��	 �K����F�x����V���8&"OV}���3cg���������Ð��9�ȟ��ʷF� ^͖��D���4I�����)��ß��#�9L���	����I��iXw�O�+`��[���?h�:�*ł�E�@	W(�*oyr�+VlìuC�hF��|��T,9�
ObQU�W)����CR$n��l�ժ�x���!��7&}���K�f��ӪI��x��xRdZ�zJ՚qnR�>�@���fV$���IDbӴ�Fz��ODY���JV"0�2�Jw�L�y�"O��.V�62����Ȕ������"��|b����$N?X`���	�L�d�h'�O�Z�!Aj�GѼ�$�O��d�O�L���?I�����@5��!��>|���* 슀m��\jP%
-���jkӧ+�z�i�Ʌ�<<�Ey�&���Vpg���i>�æ���6!�t��@th!1%E�9E�iAB�^:qNaEy���?���`N��P�X�S|�I�% -���G,���Ov�Cgŏ9��sm��$|;e"O^<(�/K��a�ꄚT���A�V���۴�?�/O!��f�O�4�'J������k1��7Y� ��@oՉ �*M�x<"�'vE����&�܅L���F"R0)'.�R� �`7���1�
�Q��W�£^�p�x���m^|=��c�r��qv$N9dҺ$q6W�O*�a%��*ڒ�Ĭڴ��$+�M������MÒ�)ۓv������xA�D)O_$�FS���I�[���z��Y���d
�;�����k~"�;w���b���Ef�q	am�&������O��d�|�����?��!v>l#�B�U��#RTs�8Z�i��� �Өm*�1�NWY�q%�	��0��T�iŴf�)Jf*P�Y����¬>���Q�^���4�� >j�|�*L.\�r�C%���O�0�b����TƏ�*����'���fg��@�<%?�O�
�t@�d
qk�+MZp��c"O�iR�`פ{ט�����:_Ό+���ȟ9Ѐ��42P�_�b�k�L���1���0��S�pL�OL��|>�$D��[VXUyG�O���4�Ї�4%��|:vX�^�( ���{jq*�JK6Y;�= ��H�&�x�*�#T�H�ZC>U��AC<6�����[>���!$��|9�(�2|
��J��ēG�&X��J�,YRT!�NݓNI~	�'y�dA�YM�F0ғ�~��4qR0��L(o�Y�*���y��>�"$J���~)<�Xa)���M#��i>!��Yy�B��N�q��Q�|�H#'ȉo�2p+�H�102�'Pb�'���Ο$�	�|�2+��(J�}Ւ0��#���uQ�\��4"Ƣ�`
�Ӷ.�Ȱgp�(�J;�O�	(��'�]*���pðD	����6��G�8D����ݶ0n��+A.ƆtN�]Bu�6D���7.O�Ra�GB=M���Tb�>�g�i�'��`P��z���D�O��ӭ?������/.?��U)W.7m ������O���4lw��d.�?eX��� w��=���ރ$�2Y�4�2ړivNmD�� (�9��:sr�E�GL_�#�Ę�3�	9B��MX�O@80�dO�7E�4pH�l�C-,(�'}^��&�0�sU��8=/4a������o�+������9��nΖ	�d�M�h!�$�i�"�'��-�:��	�@K�.�L�y��Û10<m��M���P8�?q�y*��O�(���<~�����.�9�]�M˔�f�����Z��E�5�(u�E(L�D�Sу�ORX��'�O?� c醞p��C�B�.����\O�<��hA��ecM�TY�U�P�SC�'b�#R K��qJr�B�]،��ˏ�E��'2E�)y����'���'C2�O�Zc�xر��2ủ9�>�2�/ODhPd�'DkY!(�r��j��'�n�Z,O.���'H�,��*�8CƄ�s���<�(,O	��'����dW 3nZ���Y��l�qT�ɲe!���gW�`V �[�h�	�D�W�5��|jN>�t! hV�ʴu�ѫJ6a��0����?����?��a;�N�O��$l>�� ��O��b���:���ZPF��ј���Ix���c"��t�p��'8��(�sK���j�@"�"�Od�@B�'L��4@\)f�,�� ��+(��Y#�?D�ї!��3V����ĀN'<H�eE=D��� �^8��G^/�$@)��>��i�'p�Da�.z�����O��Ӈ�����#a��㟷 ��7��!.�f�d�O��Ē,8U��D&�?yKb	;���˳.��J!�p���(ړ �J�G�D`I<8B�,(����b��8Ⴏ���hO�Xr�'�,"|*��$���֥W/``I��r�<�A����|��G�/u3X� iX�L!�O�@�E$��w�Ya�%E�6DP�r�Y�p��芄�M;���?�/�`|����O��m:�e���k���:�o�@r1nZ5/y L��x�S��}�$�&Mg�\���O��YK�(��?醠�l����4]� X�1Z�4+S��&�` ,�O�%��';�O?cU��I�Qs�͆f�N�+�i�<!��C��l�a��ŀT �qv'Mb�'��"�Ъ�/q���yr�ƫ*�4���e�5����'pr���б)S�'���'���kݥ�i��Sf�Μ5P��d�Ζ芄 �h~Ӯ�$��n��h@��� ����cnx%Ղ�]�� �3�P�8�`iy@Z�b_��x�
O����l�|r���f�O
|���%8{�<��a�t�����iAb'��z������O��	'R~~�+�*��vEd���Y�q�#=�Ǔr<X#�̀3x�LQ���7��MmZ��M���i��'�1@v�O+�ɟ[V ��h�Y�A��U�-B`�V*W�����֟@��柔Zw�r�'1��� l	�x�@�
�:n��0'%yF�����<B|��2"2�p=��D��r���K�L�x�!�Q�I5��l�e[����/۸>S���%�&e���<I֪��T'oH5D�v쳧ݴ+��u��Ν�MCՔx2�'-"�T?��e�ܔB���jք��C-@I`�/�d/�O���W��#K��K��6.��4�P�T��40��Q��Kaa̰����Oh��O�%Ze�NV�"�56m�r���d�O��ă�<�HAd��$��عRG¿RF���'�ލ��EC�_^ bf�F�y�z�G{"��)@O���3� �D)�/P(n��T�C@�0cwF�|���1��'�ў`;���OH��:�-
�xi�L�����
���?Y
�X�D���ꘘr����te��:ZQ��	����-��D�QOI�[��{�ꋤq��I�%�V���4�?9����i>L����O���R/Ga�q���8OL�� ���r�n 9�E1�cCop��&�J����'�S�|��p��l�$b����� �) >x�ɳ+��a(!�D�9��,��I�E�p�G��)���y���'����O #��H��?9�������'A���-J:sT.$�
�#�U�)�!�_(jւ��X/Y_`�pƌ��/*���������z��q��I�[�=ӁƨM?z�l��0��*�(�bO̟��	ʟ��-�u��'���!a�?Y��lK�
�<��
��J�002F�
�}�r�	0eЦ:"B�'�O�)�땤a�Y��J+kx)˥	A�:Ժ����[}r4jҰ�Yk/��#<I��P_��س쟅=Z��fZby��2�?���?��џZpC�
D\�؀��Vw�ɰr"O���a�����)��_�W�%x1�i�#=ͧ�?�,O�8�uh�9�A�5
A�yʲ�+��W�K#�T*C�Ov���O^�dNݺ#��?�O&�EᐁLE6<�!�&T9�� �����aH0S��������џl��i ��p.me��
'��L1PR'ω��]�U�·9`�E� I�?qp� ��q�lW�U�Z�Z#Lڎ'v��C�i��� ���b�N":d #`��,[�*]Z��?D�p:4jX7�,q����p{� ��,�>q��iV���I��\faa�'���!J��x�R���/�06c�0�bE�6��x�"Oh�Y�'׆96v��rD�T��E�"O6P���b�$:wj҆_����S"Ob��b�M)'�>���ߍ_�8��R"O`�H��z��
D/Z�;``b�"O]AU��Y���G�^�vx��"OQ�sH	�rV�c5iO?|0��"O���6���p��WO��"+)h"O��P�E0.)��r�B�H}�e"OZ�Z��Ͼ-�^��J܁;��h��"Oh�4*d��D��)ۯq���JQ"O�� �i̳oT�Pb�m΢X$i��"O~yQ���f�
�l��`$��	"O �i�K�(�N�8��JV1("O��⧫���zV�J�8*�ы�"O��R�ʉ@U�ᳵ'��n��s�"O����	�@Q��Y<t�ȹ�"O8xXя� q�IbaE�F@F9��"O�\��b���΅ڇ��6����"Op �rB��1��E��)J�m���;3"O�8��l@
s�(ي����' �(�"O0y ���g��A /X@&b�"O��n�	�Fi��@,�|�!�"O�� A�V��1�\T�^�"O���e��GYv-�D�3f?���"O�,h�'N
4LXc�C>]R��s�"O0��ś2�z%�6�^�c�6p��"O6�q�˴8h�c�5�!�"O(�� m��m�P�\�6�� �"O:��cL�5p��aZ�7H�r��"O�)c%�(1�%;� f�:�r�"O(�5i�
vE8�M�И��f"O2�cviD0N���BMS��|L�g"Oܠ3S��z6���,58���"O:��#H�op ���I�B!6��A"O�Dh�*0ƙ谉�.' �4"O�a�0+Mo>�m��=We�|�T"O�ܒN�9?���3
߭&Z:��q"O��Сν&�<2�:=A�0kF"OʤP5IۊЦ�SAN?(�XHH "Oܘ�l�)p$Q`�*l��͓�"Ox=p�@<4^Ya�g�8/��"O(U:��׭�m��fS>_e�&"O"H�B�[�	����Ao�=gl��91*O"T�3eN?Pe����5irQ;�'���`����}Դ=c�)'��$�'�m�P�OGb��9r�מ"��@�'F4CD1^[l�
C�ؑTs����'^����6:q^�2��#!��
�'�lYD�ղE��=�r�����	�'���S�V�Nri�֟6� ��	�'��sm��)|:H p֭(���	�'l���-�&AnƩ:t�'[�t�0�'�lA"$�@�<�0�J�#A�، �'&n!�a��<8锹ʦ���eh	�'���{�M;^f��!�1
�$B	�'r4����){���c�o�8 ���(�'H����,Ӏ(�d�b�|�'��ى�*Y�b^���Fm�;���	�'^�2���4k�bU��D)X �"�'��(�P�C4�p�QEVH�"��	��� zQ�RN6 h�������t$"O���(Q�!�J�R�νS��=��"O�I��C?~�]���^6vv�۶"O��b���a4(L�CNȕ�`"O�;�^54�8eK#�'�X�"O�iؠJ�䅑&^`F���{N!��
�Ph���uƕX|:�qa�6 �!��Qk�$����[�����Ed!�D]�T�td�3�T��÷iG$NR!�9#�Lj�JN����6��0D��ǿ@���1�lI�A$�	ۄ���y�!��Nk�[�Oyl� �����yb�.\��4�`Q"�,�y���+�@�6M�`p��͔<�ya�:hz����D$�t����y�&�<x8|0��7"'d�����yRcۦo57
!��yR򡌀!�!��5L������W�����H�!�$�2 ϶\���k�DQ#��
�!�d(����-��Q�gW�<�!���(`^����jE�A�4�j>!��Z5�H�0Td��2�R�b�EX7F!��U�uS�N�u�*��ܖy�!�C��԰ V�^=�K�5n�!��3e���B�*
"��Ԋ�/�!�D�������8v1�Q�h�!򄊔��Y�"�/\z�|p��
�d�!���L�
S��1h�t�W��/1!�D��'h.d���'�N���B� �!��ҡM%R�`S�ϣ]�$����	�!�H/Ƞ���#Z̺1�ǋ�9-s!�>BpH��V	'!/���Ŋ;�!�d�*|��� �I d�d	�F�[Y!�DG?M�8����!l�X#���7W!��y5nP��m�pC�yȇ��4K!�d��Aɜu�I]�:�;���!�ϲ`�Ӥ_�t�ꨉ1�	�.�!�dE-cx��vaˠ�$)3�+@��!�$
(C�\H��;��i v�\�B)!��	)��]��j˘-v2�Q5��$}!����18c�.-7�ɸ�mM(X!��B�Ve�ʶH[�z>�!���eS!�ht+%c�zy�G��H�!�?zP��B�J�#4�E�c�gC!���+R�ٴbE�# &�c�$8�!�D߆�`} G�7x�y�˝>/�!�أi�� ��)��K��V	!����	נ�?�V �)ɩ)�!�_�s.����I����r�Fm�!��(HH���&�j�e�İO?!�$��zϚu*c�Ы0�@��D
�s�!���9]_.i�S&�-xL����f��F1!�DY+��䒑mE�>��x��F��Lr!�Ď.E��`J��ʋx�j�2��˨;!�R?��Q��d���20c��Ukn!��� w"d�Q��@FY
����	�!�$B�ףׁ��mBcm�_�!�䀨�
VC��5���P�H �!��;X�&�`#)\�o�x%�,[Z�!�Dٺ|$`�E��2��"@�#-!��H�v=ȱ
0=fd9�a	�!�đ@��9;"ڜF_�t���":!�O�$2���%�O�d����x!�dǟi�Xۤ�2O���IAi!�� r�P'�ܔU������/;Y��
�"O*؂� ^-c>�u@g
֏}P�q �"Oi�A��� m8�O*
��Yx�"O&5:6�ܙB�b���'ݐU�81�w"Op�X��Zb�KqV#��a�"O�͸�"��|���f�=3�xX"Od ���	 �Y�b�
}R"O�-s��m��T�R�Q�d6ָS6"O�0�P���T��5�um����	`"O�%�Wh�K��x$��*[0��	"O|�0���A�<�ń�5Z�H "O�C�8>زő�*
vw���"Op�E� T}�\1r�!3��"�"OF�x�h�L��`�ï�:.��i�"O-a�':����MA�_3�ŠB"O��*Ǭ\�n���q�a�N]�b"Ob	�c��r�����D�ĸc�"O� )#�?i��P!����Jq"O�e���=���C��P�rD1�"Op�*'��WCX=����8�Ru��"O��"�Gɷ�2U��eS#
4�P� "Ox!�P�Մ ���FD dD��"O�إ��i)(H�UE����}�B"OZ����Δ8�����$N��lSA"O�H�`���S��hK#虓5HT"�"Ox��K� 1ԸrF1�`<�"OB��s�Л �(����2I�x��u"OR�X���d4((�dN0'?�i��"O�-ұ�ʙ(]$qA�)�<o-�h�"OLQɦ!�&h��t��߃s�I9@"O�x�V�i�Y��խڞ4Ye"OIe�Q���4�Be�)>ʢ ��"Oze��!�3dY���"Q=�1b6"O����B�;}S�liRb��82$�"O��5@�=�|��c�M!�)1�'�`�d)$ �
@�e��_N����'0j1�5J��$�RQ1����'
(p��M1Y�K�J[�C떡��'�,�� &ܭ!��Y�rn]COP��
�'�N��b ��
��fϏ~��Q
�'v�KSP�Ta��	�-&��	�'��5��EL�HA`e��dŭh����'��x�W%���6�8��*�:e#�'s�95�����WC$[�����'ȕ ��4(.N���h�WFE
	�';X���Ȝ� u�ͫ<C�Q�'�N���9�͐RD  ~UH�[�'����g^�!�ß�^���S�'hX�Pg�G��X��8 Z~���'��ia�n�1��2`H�?�b���'EL,j�a�j������F>2D�X�'�
Ha��P�Q��S�$/hXe�
�'L"9�ae�S��Qe��^zт
�'�|% qo�D���i�Y\��Q
�'n��B皝:�d%��h�V��h	
�'~��*�S�9�0�ǍME�M�'���R�¡=��hb�J�B��|�	�'-p���"B!`c͋���.��m��'Z"��R�׳���r�H&,2*Q�	�'�x����N�38@�z"#�7n�*A	�'�����
, �uAA &��r�'��Q��4���A�0:���'A�������0 Kq�ՀzZU�ȓ|�[R�G?��I��ņ�}Dm��S�? p=
s	� ��%���4&��:$"Ob�U'B�����QgH<S�"O��T�J�`�Ȉ��=c�xQ�"O�=�O�s+��K��E�d��"O6�����V��D��jً�
��"O0X*�΄"_�<<�1����`Q"OH��4�Y:����M�r�	�i�R�q��&( h#�΀3dv6�'C$y��C/1E�i���*TS!򄌦	���۠J��&��Dn�3P!��Wc�։2�QM�|@;�JQ�tM!����:u(���t�|�ɵ`_�Z�!�d�nq~�uk��Hf�[�ϑ4?!�d�n��@#B3?7r��d�V�90!�(xl��m۠04���E� ++!�@},�:�P.$��I�ȋ��!򤒗kP����!1���	ͩ-�!�Z�P�2�ʊ1���
*r�!�dV�
�~��4��؅C��h!�$?�Ҕ�%�ؙ"݌��ȗ%�!�D׉w�LX
7ᇕ e�U��hޓUv!��7f&���6(��[d�J�E�@!�!��B�q<~9��mH�W�!�d+c�v�3f �*���!�()�!�$R*io8�hf�٨|�����ו�!�i���BLP&e����Ga�!�Ă}��kd��u�湃��Ҩ\�!�䛌[�Bm�ဟ�']�|"	#D�!��J4>���
lܻ
[vء���/M�!�$N�B\�H�eɤ QP�� �>j�!�$qA���ʅ�j3�)�	#Sl!�dVw��6��5{)l�bHіBy!���{/XىD��9B�X��W�F�!�]6�[@��*t�Pã�_)h�!��S
|��	��p����%��L��򄇌<nu�#�)i����0�yb(�F|��&��/�p5P�A���y2�Ɍaz-3��%tB�a�jc!�d�]� m�S(½)&ǉ�b�!��Z�:a&-0���		NC!��̢���#M<HB���%-Y!�M3�8�8�Ʌ X5���4��AQ!�ď'}�*QS�!R�ʢ̺�B��;�!� U�z]�ʖ�6� �B�E0�!�DEpҘ%��BGLJ�3��D!�DғI�0�Q5t\�tk���d(!�[<T�ڍs3�2rH�<�'�M�D!�dO3�6��SMI�aJR����"�!�d�D�n���F��F������1L�!��:4�k�̄2Tۘu��ϔ��!�$-"y�5�I�{s�Y�(o�!���w+N\27�-v�jT[�-���!��?E������_��z�R�+ڳ-�!�Ę�7=6��CȜm�`ۥ�� ?�!�9 ��u����P�6YK"K� �!�֞,h�����9`�����
&A�!�d�4�����\y4dȕ,�!�D�^�7%%S���c�Oh!�d_�$��I�Jd��!��%$d!��z���0��=��A�wf�l!��z��=�g�Z��m��><!��q�JԱQ�5_�^�	wEU&-!�г@���p��&� X�GCA�k�!��M�(��{���hvH�:A�r!��B�pr\A��7���!�/<T!�� ~�p�o"���+2�P�p$tmB"O�|�"g�+m%�1.>Ω:�"Of�ɔ�^�&��C��1�FT��"O�M1��6Ḩ�bc�7f�2M�A"OjA 䔱��tR��ʹx;"Onpr�׌	6�����.�(�Kt"O<�$�1(Z J�i�U��Uۃ"OĹ�Ġ�'gN���)ݚUҌc"Ol�Sd��>`�8tqHX�\ ��V"OЙ�M�{�a��!�"�Q0"O�ep�Ut�b
=>���(�"O��[��֐pq�P��
_�j��B"O5�@���	b����Y��"O^pD�Lr6��p	:Kղ4�"O��%��h<↏V4d.<��"O!�������G����"O8i0�L>�
I�ѨW�6�U"O������H�^1y�F��qpu�q"Oflr'����4�SM�MV�]�A"O��c#� ��!!�N��EG���*O6���(�`�v�r��J:
���
�'?�� b�Ä2|~ɶ��/Kw�a�'?�5J���M�t��Xw/����'Z>�$c[�U�{P�[�iw�}I�'{�����K�-<=2Pe�8��*�'!|3��L�b����Vb���'���h�g��&fBD�ä�8F$�q�'�l���U��A#/��*?j58�'?"e��L�-�̝�%lֹ4� Xi�'?�	�w͍ |��!�O�}�	�'Q��1u�U�W�� b%R/"ά��	�'w4l3 ��"ldj���>ݣ	�'n�T����-	i(uy�oŭp����'��C�0V~l��k !4��'� ӭ��Pxq12J
:E��R
�'Nay�C	LE��Qτ��`A	�'�t�+W�:l0p1V@jP�#�'�h�(��C�>3|��_+ ^��8�'ĥa���/_��å`;A�a�'(��q���"w�0���� ���'�"�jp�ԳN[Bq*.I{��P�'`��z�
��~9���;q��H��'�di9m@���d��Lo�\01�'�(�C����za�m���;] �Mh�'' �+A�߭D��H[�'
N�U�
�'��m�0ͪxej���o��qԌ2�'o��{��(`;��*�E�0yf\aK
�'����.Q�"� !�t��9rO��	�'ql���a $��ؠ�MP)e5ԌA	�'�Z�MX[f��ů�`��)��'�L bu$#{i*���;\��A�'�JЪ"�%c�uD�U,IDd��'p������ IH�!Ԑla����'I��k��_�`��&��leh
���'J,���'��{o�0Vc���L��'t�4;�@LU��ke'E�t�x�
�}�/t��ħ(~�lX�U�]���+�c�;k�z̈́�'����<O��#��!�$����D��(��ɩ&kn��qm����� �T�;�FB�If�M�2��m��-���O-�5�������%N��S��b-p)��ΏK�6��d֗d˼٪E�>I�!��9��Yc�,+:>�� ���<)ӄZ ����&��Sl�94L�'�p��� $�Gb8�@)�4��(��
k9t)��S�? ѹ���Z�Xh�3"�0T�V�h�"OpA+��Ŭ-44؃a�&n �"O��5D* X�!a���٘�"O�<h����f��l��$�"O���Ȃ1ju�`E�~oPTb�"OЈ�bP�i�4���ҹ1�Θ1$"O�m���bfx�*��F�1���E"O*Y1EZ�.E��8U�U0u�4�T"O���1q�0���F�ADH���"O���ʖ7����G��?��0"O��{�L]��ً�!�1( L�8�"O����ޏ9�R)��62ց��"O\-�Uh�x|Y���6�h�f"Oɢqi�ft�a饋�P�lP�U"OvL���2	vMڷ�M��za"O�iz6�؟/L�UR�)�<
�D|(�"O����)��%adΔk���s�"O(�ɴ,�6"��P���Ҁ8�"O��(��/ޒ�"``�B���"O�����Y s1��-�� ��M�#"O�< �ݘE?�4���#�h(d"O�I{�8�Zx�#MM#y���s�"O��{&F��ƑHL�i�m�a"O]y�&'2������R>Ru�W"O��AJ�[T��䋋 7P��"O����Hƒ
]�c�N�u�:@"Op5��$��"�����Ȃ�
�Z�"O~9��΁e#�z'��<(,�3"O"}��Q�o���� �Z�<��"O���@��qPRt�R	ֈl"r(p"O�i�uhV�8��0�B�܀Y𠒳"O,�1흟0�K'GK'�*�1"O�,*��2s� �#��c�� �"O��R&ʊ�Zy��C�~�<#�"Oh@���.c�l�C�S5(�!"Oxbī��H�P ��K
�<5x�"O8���i�a'8QW$^*s�ڑ�%"O�s�L �M*��/~�yR�"OڰZ���r���`M�^zZ���"O�DP�e� IՖ)AT�1pE|AQ�"O���e�р4�h�4NS�r�0,(�"O���U�΀a8(��Fz��pq"ODlHS֤��Y5�]i�N�J�"Oh)spj��s�v,Pu$S.�r�B"OVa8"���*X���ȨL��۳"ON�A�����*�H�E��b��`�"O�e"5���~�P�#�O������"O&p:b�ѨY������T��`"Ox��EB�jH��2k�M~�k"O�p��O3A�
aE���Y]��"O�� 'ƙ��RY@a�ǅ>X��"O@p2��D9<��bO�*$�U��"OPd�S��*h��(��*wp\;"OZ��i�O�<��홱j��%p"O0��ƊF4"�z�I�BT%?�q� "O8�T@�$N��ݫ� ��	���"O�Xb�a�X�\5��)F��s'"O��� T9��$��o���"O~����
�H�
C�4OҪP�f"O
��DD�?{z�]��^P1�](�"O@�p�i�q�g_*01�"O��P�M+��4&K�E?\��r"OF9#0�
�Ȣ)GE�-G�b��"O8 J#��f޸"e#,��@�"O� ��@�$àd��ᏽLqR��p"O�0"G�҇Y|<��A�_�J^$��"OH���j�B���񤄳� ��"OHq@�ȇ�$�pA��ż]���"O����Ew�֙C��� %�0���"O���'��Az���g�pK��hF"O��p�.E�DM��,=8T�"ODّ���[W�m#4�]�#<<�BB"O�!��(�'�t$K@DY�bZ�]"OD��ef�/P�0Hx���"q<���c"Olx���/Q��(��CW0��ųw"O��	��
  �      Ĵ���	��ZpC$��8<���dC}"�ײK*<ac�ʄ��iZ�Fm��x� �^6�	�^j�P��'�P���# h�E��$�0Pn��M�Bhǆ�.
�!�4\��'g�P��ß��'��10@5��jݧ���A��4��5��P�p�]���}�N�(gY��R��d-ޯ\����U�A���uA���Iv�1�G�B�>5�I#Tk����� 
/�剎xR2�����<���y0�)�r��5��~X$���v�B 6#ұ$>�		�3����P�l*PL!��.��r��_��4'&���p#�a��ěA�,H+��Ꟁ� �	��	���N�͊�Ȧ�LCE34t�hJ���Q����J�L��á
���22�ئV�P�M^�f�}��yy��OZiY�P�:����<YbA	h���Q ��)b����p���2Q�����<	���O�̹SiOT����O����zE��O#He����v66�A���(7���ô��O �!*˙
��'Ψ�B�O�:$��8�'��,@BΓ8��YP��X�]��JB����S�SyRD	�: ���'�X�I)5=�M*��'lz��� �z�,�� F�X�Z��O0X	�i��'K����)��Ƀб�䂖>M�Y����<_�=�4�S�F���'��j% �a�j�O>u[Zl�ȁ�9y"��+e$T}L1��$�I�I&+��!��� ��.p/��0OnQр�Y<"��ȸDW�]oZ�#aP���N����O�q��B���'�n}Q�_�y���:5�(�,��K�~R7�y�4��f���(#�?y7O�!��%ƙY�� �\�^~Q��@����E�@�w��E���=9�HӤ�	��y'>�Z鋓@�?��A)r�'�t��`hŦM�j�F��v�
���O���R(�#�(O\<�N�؋�n�K�bE[�N�%�͐@F�>��%4�"<���U����ٹ#l�"A5�!�ʊ# �  �i���]�pU��:uG��i�Ȩ�`�2*T��'St�S����3&��yFD�(��H�;FY��9g
9��?�{BL&EH)��@���$��u��7>q���qO���b�3��?����2�� ����H4`��Ȁ��I!^��R��7$T&��I��ܐT���B`,>��,��#��r԰�ad�����ÂO�S0t��?Q��������LC0!�]��	@KFQ���� A��   
  �  5  �  q+  +7  �B  eN  iY  �c  �l  �u  }  M�  �  H�  ؠ  E�  ��  ˳  �  P�  ��  ��  -�  ��  ��  #�  e�  ��  ��  ��  � � � �) �1 I> IN �W �^ �d 1k �l  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H����<�۴#��M  N�2��e�wH� Cs�e��2 mj`Ni������	�<��ȓLu�8�5��%*���D����l����f�$'�VDc����8�ȓ��E$����"'����5p�d@�aY�V�*��g�Pt�ȓ=U҄h��p7��u�ޅ=��$�m#ᡃ�J�^�*d�+�"OD0Jć�;U��*R�V_��S�'ў�"�9:��au��qM�̋t�<D�h ��Z� &����#G���ǹ<���2�S�Oq,(��Ֆ @QJC��38Y�'�`��N��e�~��S�·0ra(O>�*lO�����@+����J<�J��"Ob������ D���X��>���"OL�`c�	 ?���6�'�B�Hq"OX�Z���e��� @�8���"O��@�eJ�FH] ��W��ơ�U"O�����F�v ��Kͭ?�
�j�"OV�&��P��Xb5$$D�"O�u�S��,\#�	Ѥh1�|+g"Ota��Ğ�E"!3"�֥"u��a�"O�q�	��0�R����J rGn�A@"O�I1�G�S������?H��,� "O� I%+*%��L�� ��qrP"O� ��jC�,LZ+�O�Y�(��f"O1�a'H����1a폰8�f�f"O\��Q�)V�i��ez��"O|��@U��AHt��L$l��"O�|r�	e�l��N�s�R�"O6��r�q�Ɂ�I�#�P�iB�N�<Y�!��~��V��q�l��[�TB䉅u��˕��,�ƽ2϶��B�	������ɸ�8!LN)n��O�q �'��)��Ej��(c!�.5l����?�ݴ*�uRtK?�ԋ�aV�m|P���|�ɰ-�$�B�Շ~��ex�I�/>B�I��N���U���c��:��B�	^$�-�1�v�hqJ��L3RV�O"�=�}�+D�eR�](Z3z<Q�lSI�<���ϩ/b���آo��p ���Dܓ��=y׋�r@���B�U��N���d(<��H
�@ؘ0aa�ѥm��� ��(@�<���8��O 4��I�(L1%�Y2F�29.��4��4�(�<��scI3{�<12�LX�".$�#���Q������%����F��52��)��A��p!�ڽG� p��*�Lȳf!�?��c���3�g?9s��w�� 1R1m�9ps%�e�<Y5mE,*�:�B��D�8�v$�1���H���'�O`M�P���!{<�
�Ò�0e�	|ӎ�AK�8F{>ia��"~����VM������Y8��&��#􀟂`�{a*͉���w�8�b� �F���E "Za��`I�,������W%�y��7:���p/
23�\,C�*��Mی��s�X� T���	�,���E�3ɰ�K�"O�ܱťT�zGq�0�;d�!�9O���:	�$aR���'0�-h�ϘT�!��\��Xi d .DА��%!� Yu�E,�u˴9ِ��x!�I�.v���2ۚp�\���^�!�D
�>�S��ݒ*N�4Y���ZƉ'�X��D�?)����Q�{���5��;�!�Z�o���ҘV�X���ο_G!�$�x��	ؕK��� ��V�M�!�d�b���2QD �P�Z���A=z�!�$Ģ7=*H �Y�������5t!�D�_^hP�A�1+q�p �C�CoayB�	�
>A���/.��Kq G^���͂*�~<bfI)��#߬
6�H����?}&bU�;� ĨU�4�Vt�b&D���Z�A��QY��@!WX����%��<A㇞<N���v�G�V!�i[��R}�<!2cS��) @�:w�:Ű�&�d�<9���EK���GIW�09H�P��	c�<a#�ׇ	�,!9q�I�܂D��Zj�<�TEϜu��A �D���k�j�<�lۜWS(��GF�J�ҵ[��	c�<���"5x4��G��6 -��&��y�<�FK�) M��z��=��@+��w�<�5�:G.)�ǁQ�`��Yd��	E����/��ʓ{��#?��ؖ�ʰ+�&��B���}��x�'�<��=D���[-Vp8��P�$����K؟(��$�P�xu. &X  �b<��6�Q����ғͤe�^L�"��,���w"O<ݹ�h��&�)Is�H6x���&ў"~ΓkV ��EǏ�Mt�`��GM�BT��N\P]��5���E��<r�x��	]<9�FC��1Q�̆9����APB�<�3G]��z�$��9��5LD�<� 2��K�z��S�n����LX�"O����Ց�U�n��� �"O2� K�
$0�p�?vi�00�"OPaʠ�Ы�:dZ"��r��E#%"O�j���5R��و��A�F
�%�`"Ov)j �47,���)�"O����E�q�0�bL3ή���"OB�SW��h�Bw�0#���4"O�qd)�!>ȼ��V/���"O�q� �(��1�j�2'Z��"O�E��	9@t`�i'�x�y�"Od���#&�l-��-J��L�[#"O�A����7� ���Y�#�=*�"O�KAN�@�0�$e�:'^Q�"O��xA�#3����j�<.���"O aSQ��-x�����D^���"OhDX�f�8q{AMH�H)�.�y��~#�e�юfr��7�҄�yl� -�T�&a�1^��9�͛�;�ў"~�K�h݊䥒 !��M
(��e鈄�ȓ#�܌P�ʎ"@02%( ._Q���I8��?��A�J ��#s�!ҵk�n�%�pK�e�#{[�m���-6P��G5D�LvL�j��DPUa׷aox$)R�%�HO~�'O$%��� �=�g�`�d�ȓ,��}�ՌS&N:�9"�<4ep�Dz��~24�B�?���E,��lcB0�ai�D�<!� �<(�5`FjQaY�+�e��<����S�	O�Lc@ܻ0D�1��F�B�ɿa�΁����)$��!RN���ʓ�0?����`�q���3�Zq�Ҧ�S���hO�u|�	�!ǔH� p �^�p��1�ȓ~��飋�P0H���,��  ��ȓT�s��<B>�� dɐ>�p��1����K���A#�A�(޲�����5��)�~q�D�	����v(�Ժ����A��9�K�=e�V��ȓi������ �<���FV���ȓ5��9q���A��ѪVHl��1��d����?q�l�`Ǐ.e�Z�ȓm���RS��̍���ؤN\�Y��SF��1��Z抅K���{|���ȓ���`���=�@�Je�Ȟ]�����/� 5�$�(i�`�.B�%�l��ȓ%7>Hc i��5N�@R����p�ȓ%������e��Pf�ٻ}-�ȓS�>L��(S!J����7��8"1���ȓ��ڢe��jiHGm�"���ȓK
��R��e���S�,� 6<�0�����h� �Q<z��ɐ~<�܅�q�h���$\�
�0�aq�A�R#�مȓ&�܌he�
:t�,���|i���J��HheN	,>V��!�J��!j����	���X*e��Ś2�I'>N���yz��.η8�|��Ph:/B��ȓc0u���!L���t�:K쨥��Y���#�_>�б���N�T�@�ȓB��m��*��e������E?NT(��ȓSnx��ْh��x�e��\cHm���\[6��(-���C%/�!f��m�ȓ*-^шr�T;��$��Lq�8�ȓ]u��ه�ޘH��,kF�Aj�&Ѕ�6O΅��"�ޚ�҃�C�b�ȓ8G��Q��R�J��9����LW����S�? �Ũ&L]9x<�#d�]{��m��岶��d��P��h�d���F9EH�NU�X�[�,`��[��t9�ޏ0�����
t����I��Y`���<�G,Ə{%X��	̟��	����I؟��I̟��I͟����^�t��4g�%]|�B��n(^���˟(�I�@�	h�	����П,�I�D.�ɩ�+�CNm�F
Y�Z(�����ʟ����|�	����IƟt�	�~���D�џa��]XT��9����D��ɟ���ퟐ�Iğ���՟8�	8Y�(�鰢&lB��T�ծEM�E�	ʟ���쟰�I���Iɟ����@�I�?vX@�⫓�t6�-I��[�!��Y�������(�����	ǟt�I��h�ɥ|��a��ه��E0Ã=fvp�	ܟ����	� ��˟��	П����+l��G�N�o�B	q�oA� ����ӟ�Iǟ��	ܟd�Iҟp�	��T��� *Q]��PGřz����T�I��I�x��ן �I۟ �I�22�E�'hԞ!��%�|*H���ӟ����T���,�I۟���֟��	�jڸ� ���:F	�ԫޯK��Iß��I���I� ��؟��Iퟐ�� +;H!BAj8/��S�
�� �����	����ӟH����T��ӟ�I�l���P��Gf� �� �!��֟t���4���|��ǟ���zoZҟ`S%	|E���+��S�� �H����OL�S�g~�n�|L��b߬n���WD�T	`����:-�	��M����y�Lz�� )�d�%W����
"8��`WЦ9�		gj��n�R~B�#,{j���Q��κ6�������,#If#�c�$��Ly���L�����"	�Bx�&��/���ݴ+2R��<Q���h����M[x��viA�^��nQ,��o�M�'C�)�Ә3�oZ�<�`,�-'�6L� ���}�Ti����<!Sj�7
��Wo���hO�i�O�]R��	M'040�+B�Lr̴
�0O���#�����ݘ'DT�I�gN%p�@�a%c�.� ��P��WF}�Kn�Ąl��<٨O92/BZ�j�j��׳yd��V��|�ՂҚ1Kpd(R(3�ӄ4A�|��L�2-@| 5hdύ����)�%��K���}y������$�cT��� �N�������	>X�dQঝ���7?� �i��O�I�B��]�!.��R����ƧM6k��D����8۴�?��1�M��O���3�B4n�H��)��,Ȝ�ұE�KN�H���L� �=ͧ��D.�Ɂ(@|X4(M�7O��*V5q����M;6�Cj���O�X��@�zi;sϫ�m�q��>���i��6-r��&>��S�P� �\lhѪS�نH�x=� *�];�0�v�>�ƫ�OV��QBa��M� p�OF�9@jù|��l�A���B�O4���d4��ʦ�!�e�dȤ�%8V<�*T�=kR��i
b��J�4�����'6�7m�1�ɞ��	 ��
₴�'�B,$�L�!h�Ӧ��6�p]�����" $�?����3��`�19�n�&]�t	�f�4}���8�N�h��Py2S�"~C@�`�0n\����Q�O̓>��F�����e���K>�U��`&^�x�PL�J��
�yBR�(�ڴt1��O�vU�"�i�dF��j8���O��l���.!���!e�N�;���ؓ�M��Ft�i>��'�2�U�%���#�X�Z��yR�|b�~�f�
��|�NU�߸u3&Jŉ6�(�
�\~�o�>���i��7�`���~�g�]]�h�Ġ��Sn����j6�H����o
���T��!\���i�3���1Z`�p�ѕdBdxЧß4�����ȟb>y�'�6�� b���&	�0 �K
$p��ӆ�<�Q�i��O0�'��7���/'���K�*Tf�	�=�Xn�џ�"i�֦iΓ�?���t0�{0E�5���X:d� �j4��
^�����?~��<9���?���?A��?I,��=Y�B$�ޙkUDǻm��a���ڦ		SC[�����⟴'?�	��MϻEK�4�`�e� iL�� X�i�46�y�L֧��O��ĝ�ț�4O���� II��
F�UxT8#?O��C(8	#R�'���<���?Q%K�1D!�uo���� �&g���?���?�����$Oئٺ�"�_y��'n��bA��l� �3֯Z�UXLH���MM}B(i�T�n�<��OFdh�h>3P$l9�mր7	x��1O�����[��`f�8u]B��2�B���u�E�O�]3���I%"	JG��+f�&�O�D�O���O��}��c��Q�*R.w-R0(ꌀ��4p���^ި8+O�Qo@�Ӽ����"�ȅ�c�A�lD��Q(��<���i��6��O	���iӎ���#"#X%D$pFf��t�4|RdcK4Ԟ���gX%9��&��'���'S��'�"�'��Za��7��A	�D2|G[�k�46�0���?q���,��$
�p���-��E�:h�AV����'	D6�������'�
��?�F�0oT%�^�
`�4����ŉ�)u��@*O�ŭ�$���]�����$��X��D�˂n��A�B��%�����O>���O��4��˓z�����J#�˵6 d�[�i��U���[��K��y"cu�6��4��l}rnz�v�mZ��X��d߇n�����ݶA�x����RAH-m�<!���x�M��[�q	/O �iZ�� �}ٖC@4D��/�O��@��=O2���Of�d�OX���O��?I�a��f-���ްsA
}��	�\���8޴;��]�,O0-nZb�I6 Z��Jb����,O(y؂q���D�֟@o���<���֦}̓�?����b~ �A��N�9�$���'�R�x�L>�+O<���O���O��p�CJ4":8��BG^!��ݹ���O6�$�<�%�i-ZL���'Z��'���@ұ�ς�j�� b���,h�:��	��M��ii��9����]ɇ�V�[�da`�G�)���&Aݕi��ǟ':0`�.l�]��d׸R������i��Bf� ��H�@�4PХ�̹Cð���̟T������)�Py�}Ӿ����50p�s���-RJ��R�]#N�ʓn��&���m}�h�,�@�3zȠi�>V��ڑ/�Ǧ	�I^�n��<��
Δmɱ���t�XA.OƀPFb��"���Ӛ3H�"s>OL��?I���?I���?���򉔹Wx>�br��J|�$CAF�[��o�[1pY�':"�O�O7=�xx0f����:&��-�r��!��Ϧ�P�4�yR���?��ɱE�o��<�k�H* ��$� :z���F�<٥N�̂�p��������O���W�v@NIn� zDKD&�('-��d�Op���O@˓P���KP�:G"�'�"A�7 W~Eʓ,�1AS��*�L�b�|o�>� �i��6�j���'���RF%	-�t�$�d�h�P�	�8mxU��m�&l�';�D�K�gR������;M�0@"�/\ޚ�P�F۟�����Iݟ�E���'�TU* Q�6I�耣�C�\� g�'AP7S�#��b��f�'�ɧyeы[��� �[;3�E�s ��y"&x�,o��Թu��¦���?�E(ܗY��XX���-M� Տ� �$�j॓m>9�L>I(O0�$�O��D�O��d�O8M2�9}��<�媗 f�(<�u�<ѡ�i�I�v�'�2�'r��[>��������V�F,?J�Ekf@�9cBb��O�mZ��Mw�'�O����O��X���.�d;�HF~�x�8����(#r,c�Y������	R��;6��'J�ɧ4�V$�d�u��IĮu!f�O����ٟD�	՟�fy��u�8�:�g�O�(��%-�.�1����
ph�g�O�Um�D��xL�I5�M+�irr�G-(�|�2�-�L�p)fA�1O�У�iJ�I�M��1�-"|'?U�ݤQ��yi��zH,�s�_p��ןH��韸���$�Iz�'X���(V��v���
�"~���-O��d�¦Q�ǩg>�ɵ�M[L>i�΍�������#J.b`5̒��*
���|�����=�6mx���I9t⮴�!�O��a�L�6���8��t���$��F�Py��D���)�dR3|?��d/X.��,B�4A���c���?����	�)�����Npa���n�����MƦa�ߴG�����ٿ!{��2���%{�}��ℤE����F9����p�<�'|�t��Zw7ԓOHE	P��jm�����<*(hq�O��m1{�^LzP��k��p�W�:�Vѳ�n���ɍ�MC����>��id���j
$K"�H��5eF�)Ey�ZAmڇwh��o�a~�
��4���"e
�	�.LH�`뛥{*��F$B�O���	Ty�'���'F��'��_>mɂ�Or[�x�)���$�![�M�EN����$�O���r�dЦ� wJ�@����4�|a��ʇI@�Q�4H4���|�O��$�'��!�C�i��ę(��aؖ΂GJ�ҧd� ���+�t�1�c�>J�Or˓��DƇRbT��w�,��l���*I�ax{ӌqir��<���6sV�Z7�,XM�ڳ�
6��+�b�>Y��ip�6ON�	�("H�1#e�BxN�B�LI C���P�:���,��K~�K��uǪ�O<H����Fk �Z�6���(�Op���O����Od�}���5=��3�$Z�d���c)��4Z��n��.�zHR�'QH6��OғO��
o�D� '�Q��F�s��Y Po�D�Ǧ�ܴ�?�W�O��M;�'L� �`>Y�0�E�E����$�5$3�t2��=7�T�[�|�_����ڟ(�	��T���X  )HzAq$Ӻ;�z<�s@Jy��`Ӧّ���O^���O2���DۙE3�m PO5`� M�@�;*����'Z�7
���cO<ͧ�z�''U:}`��9
�d�(�ʃ��ʍ�Q����b*OT8�e�ԛN0�ݪ����$�x����ס�uph 2�
6���O|�d�O��4��ʓ4����J�F�!�r�"%��ZF:��V-*c2tӲ��ʭO�l�
�M��lQ�5�qm�"KpT2텰bJ�Jǈ̰�M;�'�rM@�Xv��g#�E����?i�׼tB ��SH�0˧�,oe�	�D����H�������R��%%��qO�4ٲ���O^|ZJ���?9��ܛ���@K�	�M�H>ag�<;<�V�w
Z$H$�ϐw�'.6���e��B�\m�<I��d�h��1ꕉ���B�(��m����T
����J��I>-O`�d�OF�d�O��B��Th���B%).����DC�O���<��i�juJF�'X��'��S5*;��i恉>�Q(�Qo��,e��=�M���ip�O��V4�Gʋ���8s��7F�lG�R��k`���0�� o�+�u)8�dI8z���z`�qs���- �����OL���O��<	@�i�\��e��B��a��%~	�ѣ�@28\�	��M{�b��>QA�i"h%�C�g;>���Zo�ؑ��tӘ�n3V,�l��<��m�]�4a�+�Txc,O� Zexa��(|d�-	�Ѣ�j�8�?O�˓�?���?!��?q���Iޢ"��!#���F<��Z�̚�
�p�nZvn���П|��~�s������ˁjҀ��ّs��9�T)pq'ô|���-~��&���?!�S��z�n��<���ߗ^��3�5֌I�D��<�[;p�9`m�����$�O��
a,�3W��]������ҝr�
���O��D�O��cǛv �2x~B�'�bE��J���[��Y�E2Hq�F�S�O\��'y�6����$���2GK�zb�H��r�\�!,l�x�I$F�[�,EZ�'������*��ϟ��/�-s06���0zIx1�� /D�����/x�֔�s��?T%<�� Oޟ��޴jt���/O� m�}�Ӽ#d&OxF�8r�2x��"���<�Ŵi:6m��-��G˦��'��ňD�����#��W�t�u���T�&��p J������`��<(6�� �`A��g�� j��͎x�v��^��)��8:��d����[�d)������yB0�B b��f̔'Ua6Q���"�r���{��d�W�����H�H 0�LO�wkv����w��рQ@����;���>�x��W�)�����mC&@K��k��1@�CĿ��I���}�4�8Ai�VC��b�)N�8�z7ϑ��Na�uEɥ:�8)BE�i�d9x�k�J{��
Ca�/NB�J7ҁS��0hWGѣ aj!rc�JN�Qj��0�M����?	���ў��z��?��1�5OR25�	�)s�����Od�2�)�ӗL��u`��08���ـDи6�E����o�ɟ@�������/���|���B�F��#֬��X-��1�ȄB�Έ�|��	͟����?c�|�I)k���2S��/�&CbK�XP���4�?1��?9eB	.9���d�'���ƞy9�7Bd(���ɟ����?�nj��<I��?1��cϺ�x��s�``h'c@�Ov�1R�i��g�bO�i�O��<qņ�&m��0��:IDX�	 ����'��T�y2�'�B�'J�	�?��(X���o�F�ç`'Q���b0�8���?9��?�-O2���O֘H�	�\����K�%?.a��\(1Oz�$�O���<Q�(����IE7EtPlaƭG`#�I��Ǎ�v@��� ��~��sy2J����D�*9���S,R'"�kՠ\$U=��ҟ��I䟬�'���b�/�	*%2@�Y���iw�8"��վt�l���'�d�'�������ϗ�� 8� �r<��k��MK��?i.O�����H�����s�]i�-fy�DJ1�Y�pϤ�C��~Ӏ��?q�-�0�G����M÷��; T:��U�m?qj�Cæ��'ZV%{��sӰ4�O.b�O�8�g�^���щn�d�b@���&��$l��0�ɶ����	���'<����L�vڐ���CE�x�޴����i	�'�R�Ow�O�,`��9��c_�|~�q��J`T���	\m�IBy����'R�Q)w�֡���Q� %Z�O/�47�O6���O����Bf�i>q��ğ�[W$�2���#�w:�]7� 3��D�O�^6*1OZ�D�O<���\�V�q�M�*`z Q�l@H�eo��vN����|����?Q,OT�iC�LA !���m�J��C����ɱ��c�l�I���	IyZZ��i� ]�j�� 1V����iL[��'>��'�'?�"d"E��,[j	j��Q��6�m?����I⟐�'Y:4Z� p>������E�>II��]kH=�sg�>���?AK>�.OlK�Q��g�Y�1�$#w�F,$�<�T��>����?�,O���D�c���'�?�֌ɦ@��z�*�)�#��7���'?�O���F�?V��^�6�؍�������#�G`7-�O�ʓ�?	q���)�O������C� �k�\�5���'�]h쓄?��,��_�P��<�O�`H#�UM��miiաF�l��O �^.O�����O"��O(���<�;<*�+�e��$g�;�f�'�hȓ<"��y��D�J잍�ċ#�A[_�vPl��!�q��ԟd�'n��T��Ο<�����Y���#q㘕�E/K��M����+N~��<E�$�'�f�zć[��rF�ߘ}`��"#�g����<!����4�j���O�ɓR��m���$!����Z�)Ԥ�Ҋy�+V�?+Z�|�D�O�	>V>�=�g�԰Q�eR [ZT6�Od��6��<����?�����'-�q �@Z��HH"-�?K��\h�OFM�������̟��Iqyb�'.]���7ro��4&Ӂ#d1ۂ�_���ڟ��I��`�?A��	Y�)��O�?�J�H�A��f���B��	m$��'���'��	��d�Tb��m�l؈�c��&�|����¦I�I���k��?y1#J3 �
�l���ȴ8�*C�}!���a�]����?y����Ov9���|��ad.�#���;\�[n]0t�k��ir���O<����
�'�Ȕ�tLU'\��Ժgh�/ Z��ڴ�?�-OR��
"Yt��'�?����)Z,Ug�$g��/n����ee�O~���;��`�e�T?u��G٤MB�6iȵJ��Р͸>q������?���?��������R-
���s�eˮ!T�HKEV���ɑ2�"�Zu�%�)�S�6�5�5"O<����ʱd= 6͛��l���O����OT��<�'�?Y�64�pl��_3z���Ѐ$؄~��	�'d"<�|����A�ԃZ�!���h�BƤ��оi���';F�i>��	��`�S�? :�Z�hW9-w������+*X��K�V�'������O��ɰi^���2(Z?pΈ�2�����7-�O�1��.�<9���?�����'�&�IB�\)Vd���!��!6�婭O�M�A�Ӱnq��ҟ4��ky��'{�=KV�	@^��'��:Jͨd�akR�l���Ο<������?���gD!��F��uY��C^�k����U�WW�Z�'�B�'���̟C"M�o�5%2��Y$Dm�MjT
Y女�I����	r��?�k�B��np�r�X���� tJ���*�|듢?�����$�O�}�c�|j�V��i{enG_P��Ї�Hg`f|:��i�����O�	�3���\��'����?Q���S��	�=>^��ܴ�?I.O���Bf]��'�?q�����Y�q]H�X�/��ȡ¦F�5xh�O��D���8����T?}���U(Y.�����w�Y3��	���#b�ӟ �����I�?}��u�n�99J�zq��@A
�I� ����O�H�f2-1O����;'(ШE�*(!0,șCk��6�iL�<���'2��'���O��i>M�I2A0�]Ð��q�:����ΪC�z<�ݴ=�t���!�X�S�O��Ce������Or����%�6��O����O(�� ��<�'�?���~�E�?p�p|z�˘30��c����c�<��g[?��'�?����~��D5Tx���  �|8��U�M��M	0]�,O(���O��D0�	 y�@ J#Y���O�~��I���HC�������Ey��'uJ��5�!/�L��G����!I;PB�I��|����H�?���SV��3�Π<� Y�����٩S)�A,��'��'��I��]�g^Fy��%��i����g�2��'nb�'��O���R H����i!p�wb��x�Z`��N��1��Ti�Or���O�˓�?�P�S����O���\�V=�}YcE�65�V4ǅ����q��?�%M˚$*I%��Є��%i�c[ ,冈r�y�z�d�<!��Ox(�(�`�D�O��	0}xe�c�2yU"8��HU�����>Y�~nmb�Qb�S�4$A�/�N�d@ˈX�|�b�������OV�Q�J�O���O����&�Ӻ%C��g(R��F�<���A}��'��L���/����O=�u
�h0x�NMrTႌ2���q޴SV����?���?��'��4���DV��8�x�H+�����"S8%oZ0>�����M,�)�'�?A����a U1�~)!�Ɩ�s��4�?a���?�B��4���d�O��I�i�J��b��8CW�0봨��ib�yB�'�X����ON��	.%k"`ݍ\�vd�%E��7�O��ȑ�<)��?���۸'���D�D�*	Q�M(s�OJ�h�W���	�<��|y��'������=����@��.(ETh!��ԩc|�I��	꟰�?I�l��%�c>=*��RJH�9,����B�@	�'7��'���՟4p��]"#Q1rT)2T��+A�Xk& \զ���P�IZ���?Q��Y�6uo�zy����G�*�H�Cs&�	M6듨?������O�Ԃ@�|"��=T�������tϢ hD7;��8�i^����O )ZU��n"�'8��c�
���)�D�3~+�Hb޴�?�+O��$� @ʧ�?1�����'�]S�1 ��w���S!��nc�OV��@�
��J0�T?��#X<`�Τ�Sj�֔��>��AN�`���?���?I�����Ra𵡆�ۂ-� t-Q�R� �I�+u\�g%�)�S�V�b`���F.%V&̱��&=��7M+k�$���O0���O��i�<�'�?9ÜrX��0�2Xm@Vk	�c$����5��<��y��I�O\a)�$NxV����>3r2��tK^ܦ��IAyRդS��i>9�	�����3c� :���S�p�{F#�uR������ޡKeth%>��I��@� 
F�� Aϸ��V,
�A}v�s�4�?��A3N؉'���'�ɧ5Fh�%�)�B
�$e)�Q��Խ�MS�g�� j��?Y���?	��?i��?�N���腪�M�%h��E'N�8�:98w��O�Oh�$�O��@��-�
lz6	�+#,5��Fٕ ,��O��d�O���O"ʓJ��A5���Z��:��Tr���Ki���Ŷi���۟�'�B�'n""��y��U�1{�u����rg���P��,*�6-�O@���O �d�<)�_�Gx��ȟ�AG��?����7B+ �4Pq�H��M������O���O@�0�?O���Q��"O4,!�exFΑ�1 �"E�i�,���O��a
�W?���ğ��S�<�x�DB-o�<�+O1oxF	(�Oh�D�O��$��c.��6�$�?z��	�9C^j����a��uj1�g�˓,�tLs�i@�'BR�O���ӺK�>2ި\��0r�I˥�%�I՟T8`�z������d.�S�_L���	=Y���Q�G��7M�24"<m����I����S:��$�<9b�������@�qB
�n��뇧�y�'L�	@�'�?�2@ܰl`l ��ރ�<0�GȎ�+a���'O�'�T�q�J�>!*O�����@�.�d�ll�R�ͷ3��|���f�ԓOp-��3O�ß����˷�u�D��6�݋�����M�4�?�޳R��Fy"�'�Ɵ�ض40ak��,X8�V �$�7-�O���7O��?q��?i(O���`8b�8` ��L�j�����G	6p��'m��ʟ��'l��'*"e/� FA"�$	�^������8؀��l��<�-Ov�D�Of�d�O6��_<>�v,oZ$���	c�3?�͒' B5��([�4�?���?����?�+O���Me�	O8̲Y�!�ߚ-�z(
5HJ�K��l����ݟ��	���I��%��%n�ԟ�I4+x� ��d͉+��b���d�p޴�?���?�/O@�d\�u�<m��sz��c	3z(���K���'BR�'�"��$-��6m�Oz�D�O����e������S�c+Qsa�ޏ8���l�����'�o�����'�Y>7���vapg�$
�4x*g��h �v�'���GGj6��O~���O�������$Y3&Y���Fɸ	�xٲ2)G���'I�c��Mp�|�Op�'p�(%�&L�Y*� �"5<!oZ0c�����4�?A��?�������?��*4���_�.@Ā��3x�Uɖ�i�t����'r_��B�����%�σk�T���ؓe�ʸ
`���M����?q��EY���'S2�O.��h�4p+�4����-?�&Ma��iC"^����Ce��?����ṫ]3��@G��0����aU�M���W轘5V�ĕ'�Z���i���ɶCQl�sv�\2*=�bn�>!�d��<�)O��$�O0�Ħ<�_:=?ҝA�Lp�'۷-v���S���':Y���I�����9O3r1q��4�V0����4��X��`�P����h��ߟ��IUy�СHÐ�ӍEQ��Qd��r���xg$�?%d7-�<Q�����O��d�OJ�S4O��y�m�P�!�E�$D��K��WΦ%�I��$��̟��	��33���M���?�A�0��	S�
e����0��O+��'r��'��I�� �$Gd>��O�Mj��4N���e�F�QǾ�G�i�B�'�"�';��T��:���OT������#�H�&G���!MX�̀!m������hyr�'N"1��O��V��s�$yr�JoцQê�*&P�(��iN��'l)�nj�����O���0�I�O`]�!�Xx�xjBǌ!hARxnEc}�'M��1��'*r\��J��V��̑Y}w )%Mm}�֢S>: �6��O\�$�O��	��x�d�O��¬-�R���Ι�[�8dY�Zv�RxmZ;U}d=��ƟH�������'4����@�ep�����ʒgs&���h���O\���q���'p�� �p��%�q�|�h'��.	��qm؟�''�X����Ov�D�O�;��8O�6m�f*ъ^�,Q1d�Rʦ��ɱZ�l�A�O>��?+O<�����9���,|�`ZD��������_�xa@�}������x��Пp��Ky��N�6{�q�	�vd�0��<���3Ȯ>�/O���<���?a��x�F�j�c���=�����I����Gc~R�'���'+�Q��Q�T�����I�A��eĎ{G`ّv*�6�M�)O����<����?���U�ʬ���$ ])p��uh֠�Ĳ�贃�榩�����ߟ4�'�u�Pc�~*��u�.y!��3J���dO$/#�y�iBrX�|����	B��՟0�I	q�(�h�@P�0�
`�#�~�b�4�?y��?y��7���iH��'�2�O#�K�!�(���$��^h<�r�}�:�D�<I��i���'�?Q*O�i���$oQJQfT�n�q3�4��Ǽ?��xoZ>��	�O���Vw~���<�q
�Lǘ[�*�8o��M����?q�K�<�J>����@�m�F�`Ư�W��US6���M��،bϛ��'�B�'�ԃ9�$�O�l˱�P?H@p�V�_%k���jG�J����doFȟ�'�����H�$8�k�42���r�	B&$%1дi���'Z���,��O��$�O��ɔD����5ď3Q�L���!Ż	d�6-7��.e���<	��?���k�� D���t�T 
����ͦ1��1��qL<I��?iJ>�1�.L���{����%�K�b �'�����'��ğ@�IԟX�'�<!�
|{X�����	4�`DD]z	�b���	F�����IFu �� �\���a��} 0�X�i��'j"�'�2P��Q3���k�3�Vk�:&F,�D�C���d�O�D#�D�O�$��^>x�d�vNl�j�g���RJ�-NZ��'���'��R�<���Y%�ħ�Ax���$xq�5	�	}y�r��i���|��'��Ño�ҟ>��e@Z�����U��,�Ĉ����̟T�'.:�b�N*�	�O��iB�<W�	.A8=Ƽ�#�ܻ3o�8&�|�	��Ă�)J��0$��&ex�A� {���bC��5M[h)nZOyM
h�7m�b��'4��:?I�hU/De�4i��VD��;B��OT�d�O�`Q��O��On�>�B��#�$���̝1XJ|��m�Vቴ�QѦ��I֟���?�1�}b�·p:���>n��s�nŽXb7�@�i���� �d'�ßh�&��J�Щ� j���.�����M����?��$r�r�xr�'(��O��C��^�T�)�FS�[�D�9v�i��'G�3`�:�	�O����O)�Q�ʫ+O����� LY����]�IcDXxI<�'�(O�11���>�)Dc ]Թ�\�L(t�䟈����L�������Hy"�rpa�g�0R^|B­�" juA�i7��O¢=����q+b�R�wӒ9Xc/G֢u��)�(�?���?���?�����iЃgMt�䌵_�&�@���hW�0c��NEnZ�h��؟�%�l��؟��d-�>�p(�N�lx�r�հ,0D*V��a}r�'��'G�'Z�19�Z>	��+�PXj%�Œ+�4kb'�O��,A(��d+���O���W\6d�J�x
� �q��@��3�x��`꓇jq$M�i��'�I0t��kH|����r�_4(����-@����PK�6P�v��ڙ�?7�@nD����<����  ʩX���'�r`��{��'�b�'�4Q��&.'�p��$ӟ|ZV�k�(1�7��O��䃀y�,}����)��:K��!eO�:+�Z@qR'��}��c�2:V�7M�O���O��ɕ}����X�CHWP�S��FG{�m�pB
��M�6��`������
j�J&��H0z�L,BAX�o������Ɵ0� (
��ē�?i��~�l�9#��]jDC7I����4K�#��'�TaÉy��?����Ԭ�h�ؖcL5O�б�uC$8`��yEl�t��c�$A�ԣ0 �x��I���.z�����g6	X� ]�)P�|9R(�
��z2I�/[�2v�ô:@,�)wȜ
(�^�[�m�'��P;P��d��y #iB�;�]Г-
�1(���ʙ <�3h��J0����P�t�� B!H�����ʔ 'lJ!JB�J �H�E��f�$�($),p�t �G�_��� ��	1�YA��;��\���nn<��i	^�vA#�K/�?a�&Zؤ���?�O)̌@�@�l�6
�'2$���,��$����y�,���X��џ�P&���8�E)�>T1��C�O����d��>.@����[>TF�J��?�A�x2�S��ԑ�0���-R&"���yb�޼:H2A�ݟs��
&�]&�x�la�:���4PB9��L��XLh�*�3���N|�n�埜�Io����n�REH9 ���X#J�+]�,�#�h�f_��'���vϒ��0�`�BH�4�l��@��m��=R�X>#��֊?$�qp A>H�2���8}���1N�@�AЮ��Yd�y+���,5k�,c�/�]�dN��&��
�*L_2Z1bp�S����l�Ėg�)�S��
������ПT�<��r"O��2��ܚ������
9j0�'(#=A��i��<���Ȼ7Ϊ�1��B���6�'�r�'����B�
+���'r��yW���}�%�#9�A�׾A�6h���W�%/�9:0'�.�r�kF�
��U�'�D $b��j��%���4e����MfGT��Rr��T�J	�Ovp`�C��<0Ό!j�k�G'*��9��Á&�?��O<�s����ɢ8G���q��_Q�h���0�(C��(�rф��a5���X���vԑ��ߟH�'o�m2�#�,h�*�Z��ȳK,(1�� ڱ]T���'�2�'�#jݡ�	���'@��=�e@�'��tj�bWE��9b�m�[��A!�>FB�Mi7)�T�����F1ʓG�уW��.x�0")��qya��[:{dfM��Α�`�!�47����iAw�'�t��9X'�؈W	H*W$��Y'���?��hO��d8"�g>Ƙ��V�,����ġ/D���cK�Ү�ec6@�0�ۤL.�ɉ�M�����d��2�Z�m�����IN�fP�!�/� �����4�	��
W��8�I�|�Ӊɹp�z�)���*'�z�g�H�X�Ղ䇙'$# 2�H�	8ܸm��U�|D�<��Ǚ>$M@��J���j՛H["2~v%+�LW�C��A!BJU�4N�� A[/���<Y0�Z��`)J<��I�PO�tp��I?܄QF�Ss�<A#�ƜYKhG;4��Q�ěr<�Եi(j(ӧ �>!��Ig��;L�]ٖ�|�
�p�7m�O"��|��5�?��l_-t@rH�`$||�	�O�4�?A���0�j�Gڗg�Th����1s/r��3(ӫ�E -�,�c��P������/MlI��>)��T�_����n
H�� :ꗟ�R��VO �u�0�ꑣǀ�I�Rd)סSC�db���#���
�x�����$E"��)�DŷY�!�d�(T0�$��h �����M�axRm.�c>.\K��Q* �5H��
xg��b��i��'4���{��!�&�' ��'��w�:\2��U�<u��{F,�4tP��x�kϭ5��A��'vx��'�;���B'PH!��ȿ\���w��5IX��B�^p�p�8�`O&�3��K��|�"'�(E�XR�s'~�&�Dr��Oq��'����Щ'| �J�+½T�\���'(PY�	�?JB�x`@KHx�%�O�yEz�O�'t��2��ݪVi�=P��+3853w�ԅ{�R���'���'W2�}ݍ�	꟠�'px6���胫[��4��QG��ᧁA�(�.8G/*JA��G���Lt�$�!./ʓ?�*��H�T�h�3\��亷��zC����n�3�jY>�$UJ3���(O��0����]l�[�IK�\c�4���ک.�20�Ob��%`���ە���$"g"O�}�*^�IT�Q5ޚv��P�e��e�*���(PY�����6���Ib�N$.�R �P��T�Q�O���/\$�d�O0擆b�A�F@]�4�:̛r�����H�K�&.���4=E��)���'O�4ٰ�����E�η&E�6m�="��a�S�3.n�x�kV*`M�xB$��?�����߳t~�-[�N*���k\�FR1O���><OJ���!?W涡K�*��\�|@�aO�<mZ��ِ�&ٴ �81zѥ����ZyRI@�?86��O,��|�����?� 89�$�Ȏ/V]�V���D��,�%��OJ�d_	:��@J'k	�/#���E �3s��ʧ=~��ª�� �D��87",`�O|���	�`�ب����Y1��:v��2�p̟D��a�
-x6�KE>����>1pl�֟�H>�
�c.�����)w�|��[�<�t+ �y�hL��O�Bf�i� Y�0��䇑
�
YC��K:B\��"�:6rjm���	ßؙ6�ˀAJ�9��՟��ٟ��yt`3�E�4�8� Ї�&+�2@��@G+e6tuhp/�|�(��OC̧#`��b�n�PSaC�;c�t&m���Hr�W�'DhRUM��S��hA0H�	Iz�>�i7aJ��d��0޼YJ��8�D�J��'
c��j�Oq��'C*�b�]3H�Ȍ�k�_��ع	�'].���"=�( r�["lA�i�O��Fz�O��'����dfR8,���rK�35��M��iY�NP���2�'���'��Fr�!�I�`�'Fb�;3���(�\���֨ZU�����٨3(�K�' ��95K>M��@��A�`4�Y��AëazdkR�3�O(��F��V#����;K��2���&�b -�O���㟅w��'�R�@<�u��"O��HcnHr�\��� Tz|S@��ߦ�$�lC�K��M����?��C+2��s�c>E�ص#�(�?�Y�����?a�Oub<����<�
��ӿ<�f�s!D]�P��x�:�LIr��572ũ�XC~̙��;O���T�'�Op�ҡՀb�*�ÉOG&�}�$"O�q;�̎5f�\�G�R��`��O~�lڄ}� 8ƃ��\1b����̈I$�\��jL�M����?�,��0��,�O���7�.E�J]2�����FA�O����D�@Qz�B !Sz�S�U>��$F�/uu қb��	��C-}r����I���A>�A���!lX�Zpl��=��0�'}�`��?9q�|���*R��h��S�"�\���֗�y�鑑g�2�re��	q8%)D&Ϲ�0<�c鉕v̽䡙�7t,����Np�ٴ�?A���?�3��5�R�#��?Y���?ͻE���1(@�>ߘ�8B��o���7�|r���]�<P��L>	0LE|����gE	F���Ă�4_��`ǅģ�y��1{,��}&�|�@�i���PP��hAJ0;�,ˏ��kEJ �)�3�$�2�Q3��L�+�����1+�!�Dvo<��r�+�+e�B>|�ɨ�HO�i)�$��4���l��v���3�ő���K�.V����O��d�O��;�?����t`�5=�F�q'n�Lo@�"@�h��l��Yg����`/�0=6J�)]d9��fL�8�˞��ZQ�u���q1Äռ���Bj��L�u��B�	 ���0S�ȼ�6�'�86�����?�!���W�<��A#�8g��pW�l�!��U�PX�t���N�<cX�y�>�,O��B"��⦝������E#�D@��0թG9_���qi�˟<��(Z�`���<ͧo!��K�m�����o\�n^X`�Aʖ�Y&a!䄏T@�t�bJ��,ʮ91c�?ʓW�A3B�f2����L�D=����P;|	���2D��!��^>Yu��IF:�dU����$�M�`�i�bB/-�R�
�KQ  �&d�q*��p�����?E�t-Q�	���3�ˎ}$j5�a��x��n��<C5-
�Ȉ��K��(�բv��O�˓:��	XG�i2�'U�S78����	�9 �,-x��Da+p���E�O��$C�yx���da�|������|j��>yt.��V�C�(DxH�4��y�DH�05�h�a��@ȼ���I�%���qS�����K��84{u�G�	��6 ^�8��y����S�'R�p��LL�x�pP!��Y�5��$�ȓX��T�P	یb-�\@�GS?�8���I;�HO"I+��	��p��	���a�����]�	ȟ��I3x�L������0��˟t�i�v�/vl�4�_�t�|rQ��*S��8dòy�AV��>��|rM<�&F�n �`'ǥC�0]9��XD 1'( ��3��ގa�RA�}M<�P�ٟ&��Q
Be'�hh� \�~t�'�hH�S�g��5	����E��z�y�Ɵ&ZB�	*{R`�"�I	0M5�[�߫o��e���S�@�$�@`�;/N�U�$��#�����܏k[���	����	���Xw���'Z�)׏E�8���M���igBT�WYh�S��8bԉBj^�fv�]چc-��m�:�C�/�(��a��|���i�#1x^d@�`A�bwv9x�Jٲ��O��y���#�l��%�!H�,�@�kY��&�O.��ҪY�;���j�0�XЀ�"O�l�-�)X�[��Ӷ4����D��6�O"D���E�I՟8�4C�	eH ��W@�-0���8b�����	Z��	˟�ϧF'��񡧚���5Iq�E'|3�� l�3�X*�vl*�G�p���X%@b�؁��*��l*����rĲ����<3JѰ���k�`ԙ $Q^�d=�3�Z�I�\ԙ��Dέe4b.��9+�His�'k&���#�=q�!�d�"|����I�+c��sgӀ2�!��Dݦq��.Z|*�0a��G�Ґ8B�PW��*@@��0ڴ�?����	��E���DUo��K"X�/��)�d�9�@���O�)�A��'hZi��-O�I�SVh�$\>yk׈�-N�6�4��d}h�c@/}R���#�"P����X��q;7/؛n�����X�*?_<i�u�=(F!�q�>����IJ>��Q"����h�tN֪=�"�tkX�<yrcq��������`��	{�t��S'q�(X�D��*OX��Ł�7�$qn�ğ��	ş�0���a����0�I���SH�a���dx���^ς��<a@8�<Q5G,lCZ8�S�:ق���b�M-&�	˓/h���ɖU��p���dt�����M1�����?��`;(4y�rܱ����sݪ(��'�=�2曧fP�� qbљ<e�A�O^�Fzʟ��b�P���lh!�p��=��m���Ŏc%����?���?٧��,�d�Oz擟!W�؅�Ë�|�	�D�:�k��-���F����*�#����:u��}��C������ �2����aH�=��!8VG�O���I'�.)(�O,s�I+���Y�C�)�&S�N�1EjZ�δU�\c�p��}� H7%V*7�O����*[Wd�����r]�-@�  �T�D�O�4���O,�Di>��C��O��Ox�U�{��$aY (Т%JP�'R0���˜2�0��q�L�R�8V�ϖ�p<�TN���AI<��%��rbV��5@� M��M�H�X�<����'{�����O�S�J�BAlRT<I6�i���9��٣b�4�[׉��W��-S�y��|��7-�O����|���ԑ�?�cLT�*�:���-���p2p���?��1���b��38H��O��A�dl�!�v����Q�`R䫔`Z ��I�W��4�f��y a��'�Kj�r��H<`�i�@����Ix�H���U�4�?���T����QI7"��4`A��'��'���2��5du����;�J��Vߑ����bڞTE�����R4SF���M���?���'t-�W펷�?���?	���`�?�|U�"r�;7͇���'K�P��b}����1�ڀ�3 ��
%X��=!��O\�����+	�A� DI�` �q��x� `(���|Rl\�.�pʀ�4H�0��y�d���
$��NK�BE`�I�`����Bi���]�Q�;<�	槕�(7���CI<'~��J��O$�$�O��$Nۺs��?ɘO�BH8fU>	S�W�]��.��'b_��x�X�Q���Ӄ��Cp�h9r�	N���8�'���[V�T*�<}��\Z��rS�@��?	��'��SF,IYr�±�JY�P�
�'���5�Lz�:P��XQ��J�yK'�I���ٴ�?��󮘰��\6L�2��2�
G�����?!���?!����(Q-�?�J>���2XF�A6@��
�f�H8�C�5�I��J��~%@P�ƽZ�B���'~\��a��'�Y��\$j �n�, ��*�'Πɂ҇	R"���M�f&�l)�'1^6������(sf�i@��.?qO0qrv"f�<�$�O�˧�����x�ۂm�$!���Q�C��^紽0���?�ҭV�?�y*��Iu�8)"��y�rة�炑g�"�'�>U�����;x08l+�L�M3�8��|Y�u�f0�i�'��?��SL-i�qHvE��� ��&D�$S&
�&k�vm[P
N�beƥ  e9OʤDzrV� F�aq���)VZ�H6 ��SMb7��O��D�O�ZkO��d�Ol�$�O�n�?Nt�93�C��iيm.E���I"�ۃR�azb^$��y3�O5��d�!�Qܓi%�y��I{7��h�&RN�S^���O>1^͟�>�O�[bI��$1�2"{�<��"OJ��B�z�^�@�@�fJH4��@����Ӟju�0�N3_���D�����ֹil�0�I�	͟l�Xw�2�'e�iWn��}2(F��ZI�5`���<B�Op�S� �t(!��zSΔ�pLF�R*�`��%�h!`O �n�'�t�! .�?qQ��$�Q؟�MK8n�6yf�&u��C�'D���`@�2'���KO�jp��)���'s�Ģ�$}���$�O.��P!��)[� цE�:�I��-�OR��K�BU��d�O��S7t4JW灉*�ȕ�/��3aX�H ���~�@�(�dX�H��i�'�T�']$u"B"Vb�#Պ��N?�Ѐ�d�+�̄�ሴ:y���(˗( џ���O��%��� $\1����4X�r̺r#*D�ذ!D�J��4+�Gc�+W#�6C!����Ahbڐ.y3wH/}:T|#�'(�I"sJpT+ܴ�?����i\L4��`�=���:�(�� �R�(�4���O\�ذ�O*c��g~�)&��8[/�=g�́! ���L�@#<��b��p�f9f� �v��G�A]���9`E«<���T99��Bㄅ,R��hZ��	�bg!��W0��QA�!���"��C}�axrF:ғ+J*���5��R�N��/�0벴i�"�'N�zkEY��'0��'��w�����۸P�v4R%jЁ}���7��K��y"�J�]��;a������G��'K�y�ϓ_h4�N<i��P�L��w#�*�y�̝��?�}&��I�DC�c�:�E�)�Y�5D�|�mX�eA�l�' �G�t�+`J4?!��)�'<R�d�����ȍ�a��(���9����TNR���?!���?����~�D�O��Q����!��
��	�2J��XS� �����UT�dx�I� &��Q�a`U�7#�C��V��T�p�4
+N���F�-r��\I�@�OE���1+ q��G<#��� �F�,
~�C�I\o���p���?�j��"��b�<�}���G�7��O��ٓ�� �,���ֱxs郎} ��D�O:Ls#�O*�Dq>��*�OO@�v��.M��8���j�QJs�'��=��R.ؓz�X7*D�P���ݐ�p<ic���iH<��Ec����L�*��%XDMZ�<�W@�n���p�8z��ћ��
V<I��i��*�N�y����vC�yDXz�y��?]F6��O��d�|�q.���?��&�8+�>���̝	r^�c�DK��?���y�l���Ƙ�򙟠�
7�|ic�K�([�����A;}�Ț��O�ʅ)����r�).ϫ&��d8��>Q&\ߟ�H>���L��$������W�-`�IBU�<����B�2��1jL��lYS�L��&l�6E[����v��M3�Ȇsen�������!+�.��E������	��])fT�r�ڪ2�r�s"ײB�TP�<����kx��!"IŽ�S0M�y\ZA���"�	�����D˕}|�;�&^�n� Y"��� b�X%�D�`�Oq��'���aN<^Il�@Ԧ�{���'�v�y��i���r'�-n�@��O2�Fz���ʓgx[�o#%l��@JU�B�r}��a9a��$�O��$�O�����?������F`mI��+'P�g+\!� �'*���6�:r�������x����n��xB"�B2��(D%i��(aB��+�"�	���?y�-3���K
�x0�`Ӑ"�[�<���ӎyװ5X����0S��2D�a�O��O*D)q	S�5��؟̱&m+
�T���lیzJ�sn�ȟ���$����	��ͧ)����IN�<!L�m�Q)��(�^!`��ōN���Ď�&��O��PVt����FL�,<2�W��p<Q�"GڟعH<�"�9E��(�W�#gG�Й�)�\�<�֡LVi�\q�&�S ��V�A<A!�i�D@84�A<_nL��A6/��aj�y2䙨&��7��Oh�D�|���8�?I!d@#LN�{4�G��1����?���O�6�Q�������@�LfL���ʂ_�VY��*}r�V��O�Ƽ���/���듉�k�fh1F�>�'����<�R �>a���N�a����CXL�<�!HH�{����70�(�UB�a� ���$�)�&`*5*�p_�L��+؇&$�oƟx��ޟ� �	N� �e��П���ɟ�ݱ{��IA4��Fk�5�7�����<��mHx�@�EU����z|�����?�ɬ	���� 8��1�E3��X3L�8jT!+e	�_�:j\���|r��=��%7�� |A�")�yO�h�����Գ|���S�#���dNV�����:��ƞk^��� o��*U��cW�� � �B4��O��d�O����޺c���?ٟO^`4��o�^�C�5i�&A���xB@0j�x�s2nX�5s���'(v󪔁�'�p��mJ�o[�`a�͒z�ez�kB��?���'�̀@��P�Bؒ�@��A�B�\��
�'!h��rh��x�;��I��´Ҍy2O6��i����4�?���pX�M�"�:y0b1P��g1�,r���?qV�]��?)���T��!�?K>��m̞��3��>c�~�[���^8�`"��"�� `Ό%�W�Y�0
���d�83��|B)���2-���.bajp��㈥�yB�G�\���ڠ�ύ^�t�I��چ�x�.x�����!X��r��8�.L�&"Oࡪ��_>w�l�K�ǅ���Z�"O��IfR�x"��fW�F�L(�"O8���AZU8��ѕo��"O�в1ÃV_��0�J�Jo E��"O3L�%�ij����EV�r5"O������r�(���]m6(��V"OHu"�@�
/4Ia�#��n3�|Y�"O>�SB��t=@i����P)���"OX�0!.Պ���!.�9E8@3�"O �R��
 �V�IQ�֕�D�V"O�� �'�J�XA�OS��0"O �K��1qY�8ڥ���An0s&"O�$iB%���cɚG=�}�Q"Oԙ�f�a��Cf@�l�h2"O8�B�Ƶ^���WmƤ@ތ@p"O�	��h�+��*���G�ň�"O���U�X5��t`\�d^�� "OP;b%C?���*�(]Y,*e"O���A�ïs/�1B��	)PHj�Qr"O$�`��]�K# �y4��i%� "OD #��Ǟx�A�r ��4R<A*u"O4Dh��U�R"n�BDE&?
U��"O��Ad�.&�;��+y�)��"O�Q�3k,}�9�f�	����"O������kS��S�A�R��x�"O�D0#�͸
��ɲ@cX804c�"On-��G=�������Q�Ɋ�"OzQ�g�]�U�$����?����%"O�@�v��85���PV/�z�ĥ�w"O��� aŬe@(N��؝�"O������	 �^L�ɘ�W���"O��EDǺ]K	
3h��=�H���"O`+���T\;`�q�����"O��YD�ǀ#���ӷ��$b����"O���Cn�F��`Þ�~�(�T�'�b���B�(������9|8�{A�.��Y�$4|*��ŏ�Z��l�!f]�_t�)�EgF�]�B=k@��VKܚv?�Q�ެp��p�.��as�.�&3�Ft���ƩIe��0�"OPA�H6Mf����Xa��h�Q��e��l�+K(�	�� :�}�;UF�!��#+˦�r#�V�Z2�H��["��1Պ��p���pq&��=(�8�!jH:S-�	
!�.W��؇
��|2��W��͂ݶ+p�Ce+ǊY�����
�F�,s0r|r�IB��"FLD,U�����N�21@�E#��� "D�}���,�8�إ�M�f����Oޜ�L��FP��C6N6���|*u�O�-� �6G�&�*19�,�P�<�%A�!:R����:߶tjbQ3Y��Y&+�#\���e[��4���9�-��B�l$4��̇,��� �"O(a��Ü�!\�9��ź-�d�q�6y���f���N�٦#Q�Y���,ړ]D�Ā�n�I��Ye˒N;|���
dQ�e#�f�b� b�
w�5\��T(�FE2I�Q+F�0g�Y��;�O ���&׫}}r�e�ЃH�䲷ቢvV �sG\�{����F�G�(�O!:�D¡(	��;FO�t��#�'� �)]m�P���A��:L�wcO҄�R*�dYإ˔�97�>�ݟsҺ0����\��d�D�2x�O�e��	��X��N	�h��5��&@�H�ii��"L�}��Q��~>Y�';Z�l���!ӳe�8u0R��@1,�8I9��ʑ�0>Y�Aڑ>֎u�6�<z6�I�mv�Y��1<6�g�[��%�2C:?4�BC�4�>�O��Uʛ6FzŬg�>�Í����=8Q)1��)��:����U�m���xcϘ�C��؛���M�ڴؐFȭw6X�O?��8
���QU,�/�Hɣb���5N���Y9E�� T��jv��s�|0Uϝ� ���RP��(��u�5.�O\�
��EΝ�4�'��H#BW�!�Y��7��<8�'�tTyjͰ��3��c�ɀu%��0��Ł7*�KSޥH������w�v9SQ���0>��É����h��C6Q0�E�DY��}����� 	!m0����|x�b�a�9��!�(Q��ȅS?AS��\�� �d([?	t���$�a2�����љX�:2� ��q��-`&���Mm�9rG�&m��!��0�J���n�G�dm����1B�Z�;.x�������nO�I�4��䊗�ah�<��&Z1\l��`ESܦ#}λB�!c�F|�)
���
�u(�����F���T
�\��Xκ����(O��%H�/��!IB��G�2Xz1�P� 	�d���{0'��W#�I��?	���c��x;��Y<B$�PB�6�P�Y%��Pf�"�A�8%��i�T���O<�aN�6���Q�F�`8�=r`Q�PU�)(td�v�l�
�K�G������p*��N�@x=sZw�BU{��������iʕJ&��n����ԝ�|�<���'-�ڴ"�$D\n�������aR!��c�EG\�a��ЊC�h�S�-2i�F�[r�>&m�: �-!��D�λso�ػ�ɭj���"q� {]0]̓_ֈ��'�R���å3��ٹ��vN��hN�c�؉aJ۬)^���E:X�f�:�⓭xf�̘�mn��y�FR�'�Jٻ�M0[�%��LЁj9�������K��E7�[�KC��K����iڗd��	{R)�"����qI��� ѓ�KӜIk�e�=��QQ#(Rt$��0o"O �`�M���h�Q����a�5H����Ħ � A`	�|��Xa��t�4����,$��O��7ݟ�� ,V�ED�4��`s�����I�F���H��؁]�@d�P�Ф+�I�o~����'m��)83_�7��?|�a�%�E�b b��_��}�1`�Lۧ!��LCtt�"M
�e<�iϓ9�b)��LW�hR��Z�� ��M٣)7ʧ%Q�fP�:gpx��HѦ0��ʅ�A25���w��/
l��_L���ڑ$'���
3ȶ�2]��d�T�X�S��	C�����d黗!#B@7����BWm	�'�NL�J�er��pc4U��{��Ԕ�p<������#]�BA��N;�� $D�Q^X1�q"����u�m�	�|Q� a"��ސI�J	q�ءvO�i��9B��6�O�c��9���� ]Q$Ox�ܳ�\�\=��u��7Y�������]��`j�랭Ȩ�%�lI���d!�X_�>(A�4O�Ee�X�PҌ���2�$��O�^��'K��S��
:~LP`C��|��1�#XpEqO��}�F�P����3�8�Ke���m�<�R�j狷�ĤO���$o��P]�(u��w$��p�.�(:�j���k�;~P�ٴW��AoB��<D,��5���a�.�!$��U{@����߸�� +�V��+�3~c��1�kH��*����U�*����[t���A�|`�퉁9N��4��/,*x�C��+���]4�Y���7<��r1i���\�A�'��@y�JWɧ�'7C4�Q�]
QǸղ�)��P!���>Ib-D(">�Ӑ�V)6�D�R�RF?�'' Z�����І����5^�αp���4�2���]���Pr���j�C�&"D�m:7�G�"�&]���˦jx�D(F�̆3C~�)fgZ޼m���O��O��'��c5n�!I32i1�EҠN��
$��c��0+�6c�$��ğ3�D�c�cӴ���0� � ��8a�'�6L�T#M��O��yZc~0���()qL*_�(�����'��A����&&��y���J>�y�C�� $4��g�:}B�9A�Hi�'��Q�%ǳ|����tO�E�W&բ\�]���)��)C��	�hzʥX���k����&-�%H�	�/P�U���;�dKע�r��@�`Z��Ja��B��0�z�c���@�RaU���'l��6�@�D��qO[�P��J�'C
(EL�-Qw�	!!Q�d�l���?ђ$�Ɩ�}�Z*Zh	bC됀@䭃%B�.nP��"��r<(J�H�Z��4��'۫Y��X���K�ܜ�b`Q�M���x�4P�:O#牃A�&ًr�@a�FU�g��<3o���w��a���@�mpAT�`���`�3�X4B�eŭ���*V鎘hOt�n�B ���QIY�:�Q��_,��	۪�P�O�l��ªW�T
g*�@,���,2&�f">���
aL$����>w��C¬�?���.�n����OЖ�2"���b@�Ύ*kqM9�  /':��ݛ\�����D_#F*�����;[)\Q!ya�2O������\P%iQC��C���e	�Q �"$��"� �㈏4T�����KQ�]2��`B�~�iAa�+|O����Q�+� 9��ζ�ġ�
iP�nZ2`Gz�Н'<2����_6C����$����� ���`�+
=�h�WK
�]
��'a.�{1��G��Q���V!_S�����'\�vI��4.>$�h`c�v�+�,-�d�Ӎ>��OR,�`B�Fg�
y�gE
�bR��R��g�$#>���@|�I�SD��`�d��<)S ��-�4�g�v�$��Iݜ60����L�=�Q(�K����;f�Q2W`?�I�0�@d�<�Lj�̆=cn��	!�<��G�T�&Ml�1�[�p���	�<)�ß33U¥ g�{�\A�# �V�.]�􂀻AY�����>
 Yb��"|O��37IE�!��A�$�ΝR�3T�6�O�版jHع�$"ג�� �$�0�^��w� �0�C���``��$���Gf��� �C�Rej�P�Q��=R�ܸ=pnZ�B!(�"D�",�Y3O �j�)�#Rdy���1��$"p�G�_v�����!o�\�7U)v$q��dW�x�@��.�59cP�`C�Q07��C�]�t�He�Ǥt|�(R ���cv(���M�njl
Gg� J8�{�C�Wt�
�����W�t`5�]"3���JB֖��	�m�3��GP2���A�'�:�$q�A�kJ_|<�b���AQ�I¦��:��X�0HZ�xyZ�E�&h��AU�'��f�"K�n�2A�_jqV|ː&����˦�͓k�¥{�j�A�B�2�ѝf\�����C����ܱ���;Mv`!�OP�c7�ʈG5�y!�К#�����yYu�ׁx�t1�B�%�R}Bn��j=���O�8�)�%$l�X�
ٴxr�ѸiN8dQ(�p��� �<�u¼0H�Q���O\ �'��1
FG��:%@�fĥ]��+�N�d������R PbV|�%+�F`0H�G*��P�����P+z��5)�3E4OV�(�cB�{�i��v�����'��q�D�
@Bc'�|x����Mv����f#0~h�tȖ%+O>��	�3��Bf¤1V���c�o���9��k�L(�i���<2o�]k��M-r�BG��..�����lP��D�M���#�Y"�>\��ɧ�-�d�$4�T�ڌ^�aA@���M�b���?�:p۱�h�85����?.~H�'o`�!�PL +w���_��8�v�Y_�1�C�A��"?�̑�KN�1�N�̩�4ϼL"W�G�UPf���헟c��e�p��&v�j��m��H�n�yJZNϼM S�V���'��Yh��M0i�� �u��O"aA�F�'���s� X�o�3$��y(&:J��a3	R�R����n�ib��@�9r0�)��'i,�%�E�Fe��:�Ə�7�e�'�"4$�DA��Z�Ne(�n܎c�x;�,qݥ���6������/<�
�P�������:_0���NV�mV� �\C`X�1'�R�y[�e
��i0��� )9�|(�gڿH�č�K|��hζ;B�Y�O�+p �0lr0�@7-��MK�9Ex�a�g���e*�jd`��V>�I�hG2]��]	qG<�z�څ?d�����'�ʵP��B������$%��p���2��O�����8r������b��7c �
��(.^�n���$�O�x��H.[wv,"��,QMx��+۴G���kF��80��RU�F�%2�l9��]��, ���X)�UH�%K
-L�aA���Hե2}�Ah�wm�PU:�-�	�����W6SD���4j��q��p�<1��(`����@E1.��K�S���@���\$1��nѾ�)qU���O��]���U�P;V�H�tC�I�e)����K��,�B���0E	�t"�~��!Y���-`��-�ݥ���=��OLP�U(ϐg%^sPH�.%�4�C��'�
H�!��$0@���6 �(�)�ɟbN2���S,"�AC��S�&Y��k�,�q�����ON,m](�4n�=*�*�i.�	�
 D\ط��}9�T��(I~��@Ňy���*�C'�H��V$SM
%�y�At�"�ɳE:"��C�����&C�x�@���)�{��I�a�P94aq���λVs&�KD���}2�4p�Y�nP�ȓ%�Lq!J�>��$����YE�h�TZ��q��_�Z^f����Ms%B���'���z��f��T�( )M���ۓj|�$���yn|��H�~_�X��ǌ>8 ��#��	T$Q���X��遗�'�əqdN {�UQI�%:�`��T�Y��p�7�ؼ@v>�4���~�O�<ᙗG�&�f��'S���S�'��ܪ���+aV�i�CN���
�'�>d{Ab�3Ȋ�����-I�h9!�'ڂTAF&��kVG�.Xu���'�< ���P&k�p� v�ȀP�L�
�'*��@GL3mR��"��]A����
�'��\�d��=v�e�BΫ?�x8�
�':i��H�����5"�;�h��'ef9PĨ[���P��!8�8a��'Ȏs�dR�rt~��g�R�G&�-*�'���8%� �h���/�j�R���'z���G҂a�
�q���i��	A�'��� WO@�E=$��v�+N0]��$2
��&���ar��K*0K:��ȓa��C�G�e:5����#W ,���S�? P�	&k.D��M���I�c�P��"O���O\#�
��f�#n_R"O�� v�׻Hܞ����/��(�"O�Iu��~�"Щ�矮K.XS6"OΜse�� �I4`�y��h��"OVq���ڽc�d����5�(�Җ"O�C�G�=�P(9EK���$"O<u�NҸc6�(�	�N��P�"ODa��NE��DvhΞVi1Qt"O0�9�D�R�4� ; n�AYf"OP���gE0HIl��(&�D���"O�i�A̓I�P����D��`�"O$�!͔���Pr�Z38'�y��"O��Ѓ�ݾmU�D�۔$����7D�,�*b�0lW��#�N���8D���R�<���1O�O5(<��	1D�Ԓ�m�K��L0��S5U�й�4�*D�p��,�>N�yI&AV5:��*'�(D�tRf�	�[��zW�յ	��di��%D�T2F
c|`S�Scn�4�E0D��-��*�dAؓ$����q�.D��3�bH�l`䄣%Ɔ�!`��2t.D��J3!�EEЍc�gP:R�\��� D��b6�
r����O�h�f�1 $D��@�HN�Z  @E(M�$�J)�U'$D��
�E܁b�5�5f�)@�
q�7D���PV /�Q�(ɹuc�8j�5D�r����yXR��*-��L��4D��X��PA*;����=��P��5D���R�@+�)��]0G|fX���(D��@���"R�촁Ẇ�'�4$�)(D���6+�-\�v�
Pd �xv��&D�H�R�gq���q�-q24�
�|�<�LY�#��5�+=AJx��	�A�<fň:�܌W$\�e%�5�rO�G�<�T�I�?�H���(+����jWG�<���K#���C��
$oT��$ȃA�<i�!��^W����
5�J�h!l�X�<��$���V��O�� ���	Z�<ɱ�	,T�2�pB�O�h�Ke�H{�<a@j���yI� �=`�i4.�v�<1�#�l �p;��6m�L]��AM�<�W�� {����L�mnZ����F�<D��Z�.�PSƈ4�N�b��A�<ɣ� 	��2���Q����{�<�Ť�m�t[tB�´qr��Hv�<���E��$��腍y���1� Po�<)0撼*b�$���Ӊ|���fh�l�<�EG������ܟ	o�yɇ�k�<���	5p(J�g��8 ��+D}�<!�Δf9L,Cc�>��u�Qs�<�SLL�I6�@34M��6dC�Øp�<)Ԡ����D�`�J'�;��m�<QRf�:Os�%@RJ�L�(x%
Ge�<9�C�� &��(C��"�1�5!e�<9%�ݲ���+B?Xv=�a�b�<A�T/�l]Y!�Z;jj�(����]�<�" ��#T*8BH��-����S�<ٳ���D��"!R40�Ƥ���R�<�%�ܿq����<.���K�I�<y�,Ft�F]8��%D�{6j_G�<yr	�4c���0dI?T�q���D�<�WG�{��ͨ��ȃ����c�@�<����0�́
�	��h�1�@�<� u)G�$,h��eS�v�8U"O�iӨ�SAB�Q�"�����"O�Hr��ɵW��5�r"ղ# �`S��D6lO�U2 ��	���*"��S\�3g�'���I�u�H���H�i�V��A��U}�B�I�C��je�ـe�p����r#?����A�'�vM#S��G�bhC��*�!��J��u�d¥�xh�0�A� �IM��(�Ll���P�lP��M�'�\y��"OR�;Q��=`|(��L؋,�tx"O�Q��H�~��!2u��@ʶ�:�"O���f�ԯus��E؟OW��"O�i�c��/F��`P�Z=X�˅"O]���+K4|�4���x,2�(�"O���U`U���p��ߒQ�$ِ"O�$�b↓K�JHSr�M�P�n��"ON�������
0Kؾ��q�"O����@�<d�v'س\�|��"O��B�A77(9���7'6	�"Oh�	E��
c-��H`��@�`�V"O*���$��(�|P�Ʈ��i"O<���+PW.�f��|�hEi�"OZ� aZ�V�Aط�B��dR�"O@pfm�&Z,����E��0�"OZ��c�ȡ"R���Dߘ�D��#"Ol�����.) 6<X��غHi�ʕ"O���@g���\bs*�2;4�����[�O�j�ɢc�r�8b�	�lq� �';�M��L8X4��E
r�D1c�'&�Ey��I�]�pH#S��3�r�"w͜�RF!�
y����fS�Zî}�SC
�
5���>q�$T>A.d����*B�u �ȁK�<q&�8+�����K�#>@�"���x�lG<7���q�2<;"ݨ�(�ְ<A��Dĉky�$����b�!%OE�Jr!�dG�cv
<S�L�&�0X�M�n�	��H������CI��4S�
SҎ913"O
��"�P3w��!CB�-Hж�A��+ʓ��'e0�kr�5l�>�W�V�S=����4�?��'���R��k�.�����(�9	����(�"Т��\+| �@IB>9]:���h���'z�yɑFH�G�>���2��6"O��x���BH�9��ŞJ�~æ*O��b5��"�eA��BZY��'|�5�Fn"w���Q��H���'�*]s��o�v�9PN	J�R���'!L!��	��h	"S∢;���B�Qx듥�<�K��(P�.3!>$Ӱ�ܶJ���#�B7D��в�ƭ8 e�UPqmԙ��5D�d�Q�Đ�@P��oW�Mh3N2D���ǥ�Ĕ ��GF.#�t����3D��ʳe?
d�)����b�@�[�%D���[�0��+��((��v�Ѿ�T�E�� j IG�s���s�j�50$��f��x�����Ĝ9z�1��Q��|��cڸ,!�DԦ:���r3�ż"VN\H�!T��!��نs�6��- >�ɑ��L�!�S$7v��gK�V�\�Ё�
2y!�Z�q�0��)���z�PV,�7�!���%5��TAˀKV�)sJ��!��I8k�:PHba�_?*��i�$�!�D��l�.�x#�����{�'^�b�!��{Ӣ��ȑ�Xl�åY�C(����/"D�P%��(<>�QuX5D����aE D�� �`Ǌ�#v��){���(R�+�"O�Qb�ʝ�o�Xp�� e.e;U"O��d��{�쩣��!t_Z c"O�9��N�d�~-��IB���"O�H{vd��L����Ǿ"(钠"O�`���I��A�3z?���"O���A��Z�ّb�	6l@�"O`�Z�GW�m���	��N�`���;2O�����#z��t��/P�+n �E���Q�������:\��H�X�Y��8u��f�!��X�R�11T5)Ò���K,k��	Q̓�h��C1C^XS��41�v��a��:�!�DݬY�b$C���h�$�+�!�d$U\ �AO�2֠����P�az2`�ߦ5%�h��4D�9�CE�fq³E!D�\i����s�rL1&-7y�Y�Sk=ʓ�hO��4R���c�VW�a�T&�Ť��D�<�Gk�f�J�@�Ӑl��x2a��k�<��`�r���!�Hi�R!�j�<Ы�%$qҩ9�C�n �\��f�<�F[��a��Q�%�>�)%�`�<AD!�&`��Xc�������XW�<Ae��5A�(|c̡>����c�|�<Y� H'	W��#u�O���%jСw�<A���H
�����4_CFH�Ul�<1���NR�Y[�U�K
y۲�_S�<�-V�H) �b�+S!ʙX��\f�<I�Gs����ChJ�C`�Y�
�_�<i�J�t#�dH�C��TAb ]�<qЌ��3:��a�Ŋ�g��1b��C�<1� �,$��Kp�in|�V��U�<�E�˨3X� P!�D:E���0/�R�<!"f<|z��e��@P0�C�O�<�E��hM�0���ƇM�r�JMLb�<��H� W�!���X���'kZu�<y�C���M��S,*�pHB0*�n�<�tOI�h+֤ؒg��Q���a�v�<Ir���[�pd̝�qҘ�x4ŉz�<!��[�Zi��I#P-�̂�cq�<���	&�B=җ�ga���m�<	�I��;����#��=�tN`�'�a�t@�����P� �DH
�3ꊭ�yB�N
yK�m[a��9p������?���'��#G�I�6��"GI�S���'���K*��R��#�*Q{��'�� ���G&x�0IN��6��
���=S6r���fH,��P�
�Z^B�	N�v�Ҕ�K�e���t�F ?�D">1����4P��*B�^�>��� �a^;:}!�L�������b|��A*w!��L1tx&(1�%��_@p1W��k�!�P9Ra�����/Y*�"�b�A�!��W�ZC�r#gV��L�j��A�*�!��Ԙ 2���޽	�
y�c�F�4�!�$� s���c2ő>ǼԈ��*2<!��/LE�F�#p@(Z�TD!�d�����)�& a2�E�2!�@ 3V.L��W~
n�!���{!�H�!V��#��s�qHc�Z;kX!���3�y�(�;"�����hV2Q!����ɶX� ���H�TC!�7mK�l�(�2c�<E���:
-!�$E7��C���>��ei�D��i!�d	U�x�1�]��=�a�Z�<�!�� P�cd(U<n��Aa�Hټ�����"Oj1�c��A)��!�N�(r˰�Z�"O&���%��L&�Ւ��\�n��"Oб�
Q�#��9����9�6M�$"O��Jb�e2h0�mL4�@��"O�izc�Ґi����į�$��U"O��Z�p:�Cܛh���i�ɋR�!�X����eC$;����'��S�!��S�>��HҦG�& �Z�\�!�d�4W
#O� �p�����!�d־�*�H@ؖM?�@r�ō�o�!�d;|6R�ID�6�2Q
7$�!�d܇(�>��v�N.�P"ģ�q�!�
�_�N��ऎ�;�V����D�!�DȚP�x��*Ҍ�q�̵#!�d�f��p(Ƈ>����
�4�!�$T#����s*��w�EqB��p�!�D�61�ұ'Zu��h%HZ-K�!�҂c���Q����5E�<!�DX-"܀����C_�ĉuF�*!���wJfā� Ǚ�P�r�E҆H;!�0�0��Bβ}��B"��t�!�F�H�l@E���(
���"O�=�!�dݺ�ֈ�E$�h@�� ǎ��!�;7��9�̙3X\Q�V�Ƌ2!��ԋ�<pA3+UE8,�	r���ZA!�č�J� �S��+v)@��+N8{�!�D��u"LX�edƙx��(���
�!��ƅw��=�&j�\�xL*�R�k!�dٵC�P���J�@v5cM�F2!�d�8%��5˧.R;c#X��E�	2!��_�Og�TH�LJ�X� i�E6!�19�V+S#uL�'��6/!�D�5s׬Hk�D4`r�1(~!���N����HY������
E/#~!�D�"=F" �gϐ�Gʰ����#%d!�C;o��{�
�r$�y
��<S!���+�*�ԫ�n�<�X�!�"O����E�J@�L��Ð[�@� �"ON� f.��C��0���,I�x���"O�H8�ã��!+�
�+ra6��"O�A��M�8�``0��:��d��"OhDyrnHhR�-��N*W�Y�"O��4EO�l�D�ʧhX*f����"O=I�BH�1N������=_���"O�9L�@�.5ZFDۆ*r:�c"O��8� ň"A	�Þ�\��H"O` +�.M"�l�@@��-s��%�w"O��H捌�{�D$�7��1�Y�"O��E"#H���Eg�}E�=��"O���5�ϞB�P��bE��66SA"O�k@��k�P�G%m'�ib "O��c�X�Ox�˲&H j�rœ�"Ov)���
�e����&�|i�1"O�̋V�[�r���%%ʺd��x�"O�� ���& ���$@�p�D�"O ���D�}�ʵ+g�[�*�jt"O���e�=S�`Q0��1.�H��"OL}xc��w+htA�QH��ٲ"OT�c��W,BP[��y� H"O�˅�V���<kr�ؘ"Қ�Ӓ"O�M�A�*7�,tR��B�L��"O�j�i�e�����'Y�d0��"O� p�	�(�b�O�7����"O� ^Q�R�W)FH�x��'�Ba`�"O�؈�o�&&��� K� ~Xt[�"O��+��=y�}��f�.^�,Q!"O�aȁ H,Fz(A�D7T�J��"O$�I�mY0�&̲s�� >���: "O�@������3�[Mc^�;u"O��W�R�]�ʽ@��G�d�W"O@�`EH�SL��K���<RГP"OP���?L�#�R��ԃ�"OP���.�bv�`׀��g�����"OX�yƯƲb��4�q����"O�5K���!:��eQ,Y�.�"O21�Ǐ�H8b�#S�ԭQ`"Oɀ��?]�PȤj�`�d�K�"OH�G*��H�D	�!�X�ڦ"O���a�g�a�	� e@T"Or��AE�'�5x2	R�a�"O$����n�raLR~���"O�A���ZD�"���J�eI2��"O�	��̗,���"n��rCT��"O���o5�y㓌[,Y׾��"O�̚#��4u�����
ϳg&@A#E"Oh��%��#U�<�e+I�j��@�"O~�HW�V�S�6�A� `,�`B�"O���@i�9\P�Z�K@�=�*W"O�d�T
߀LPpPA�^<�:]��"O��sF��U��p�4� KuP���"O�ոנ['����G�P�|���#&"O}(`�J���b�DӠ�$��t"O��sɐ�{+V�:�h�d"O\pdkˆv���F��++�:Yq "ORD+�nIM{@��3�M��xi�"O4yK��^�8R+̏r92��"O��`�֟T1��0�B*|�-��"OH���	lαY���M����"OI��oC��h�J�&~����"O�E���?J�����n�v�g"O��� 'S�e_��2��������y�m�5+�����Yzݪ!
�Y��y���4px4��K){=�D �!��y�G��J"�p感�x}��#���y��Q�"������پtS|y����yBƒ(s�P���B�m1�೧/�
�y҉�)���%����)&ԑ��'���	p�+iP(j��> ���'��8Qa^?���H ��h��4�
�'�ԃC�M�bB1;`��cJ�I�
�'F��x3���#L^UC��\�@�'�j\�AN�?xsV����\�Ze�xr�'�@e�m�$ 	��*��86�%P�'�z��@L�4*���P��:x 	�'L0��c&Ǣg��
�:QnI��' b�4"ҡZZ��G ט���'sx��ɓ�ZGb�S%���ZfdQ�'������?C��x�K�1~	���
�'�PHb`�/bXP	��s��E�	�'�ZC@`�97����n¿pF(\��'�.Hq��ײo.��4�B�쌹Y�'o��h�����%���	
Jv(c�'=��t�]t��y��A�M����'�: xPBϦ����FU�F`d�)�')T���F�m��C���0;6����'��"�����I�e��4[=B�'Q�g�����!Vb�lS����y
� 2|�2,$(uSuI1T�a��"O��1E��H{51�� �l��!`B"O��Ce��d](�A#iR�/p�X�"O�4�F���b��T
ãm.�Ö"O
A į��L��À�Cc"���"Ohx5�8i�6{��.=R�@�G"OHU��Ņbs��A��N->�tu��"O&�vmF�
_4�!jc�����"O���ccT1e�$|ٵf�$Ȗ�K�"O��b2!A����:@��p�V�q"OYc����d��J%U$u("O����PD�X�(D�ô	N�p{6"O����NH�L݂=���+N�E*W"O�p��$��I�U�&�:({u"O�Թd�V�-Ŕݒ!�>|�J��"OP,j�'@/&M�0� +R�*��("O�� C�[�4�9�P���Y1�"O�k��C����T���z���{�!�d�	�P�֭T�~�����8b�!�߬ +F�;�������y7"��V�!�d�dYl��a��y�Tmx�G�#,�!�DB�FȌ�@4Tm������-�!�B'+|<$J�<=j:�À��(�!���3`��[�HV�pY�ty3��92�!�_�R�\�+�%|���cD'�!��?��sԆ�7-�V��RCɫ!'!�d��M�~m�FmI,
��%�Vk�/�!�d�9o�XR�̰q����pIQ�Z!򄛙E�±pjZ7|��邑M�4(!򤇔H����$`X���V��K!�����ڟ`[����	Ԃg�!�O��`ѲP���0��l���]�`�!��"�� ��ЈTa"��0"4]�!��)MpIIB��`WE�#`��6�!�]�7�~` �ҺyM2�P�i]$*�!�dG |n���dMϞ'�~�(aj7C�!���k�~m�4��'^�QB'�C3+
!��Q0c��̑�-C�I-L�*��ĄZ�!�G�:.����I0*��6�B�T~!�D�0���eG�`|�`�ߍw!�D_�je]J!�H'U쮄#�j�x[!�.ޜ@�!'~(�G���x<!�N>a>(����)EG�x6jE�r�!���d��b�GL(ǩ_ p�!��J�r\���+I8��jQ�Z1q�!�O!#����D�h��"�1�!�Û �<|���Ж2U�% dc�8w!�$�F���.S�Q10�����(Zu!�	<�~�#tFA4w�V�R�!<]�!�d�:f8v�`3�Ջe��㧁ҐV!�DѳRJ��ȟp�8ɃO�< !�$�?6��
Pʋ�{�
��5�!�Ә2\�x��$�f�L`+Ǉ��}�!���-m�2��R�� �t�بN�!�¢mv�hr�M+^d��P�%+"p!�� �*�	u�
�yF�d�Ǉ�SZ!�ĕ�L$��:gjP?!6�1�Zqy���z�O��D�14�~܅�`�����N�n��"wJ+\�"��ȓ~��ň�{弬RuB���f��ȓ'�ڈ�bA>~	�ѻ�-�#'4����A�
�R��R,��M�eEZ���E���b) p�F6c��Ʀ6*~�|��S�4[��O�n�D-�g�^�\
���S�?  <�%�C�8����0H�`�"O�`5-Z�7dP@N�q�=y�"ON��'w�~:'��m\�l��"O�p���4q6�!�gbN3M0)��"O��c��"$��}@��D0��x�"O� ����"�]��S�T�`�"O(=�E�
�S\�t���N�慪�"O�T�V�R��	� �%9�V0S�"O�D��� ���֍t��1�"OV܂�9'V�B �bT+\��Py!�>��9�fW<H'�@Y�Ro�<v�]+M������6[�����VD�<�g��rl
X�`牳;wx�Zv#V�<�v�L?bHִ���R�<����#@z�<��Qp��G��ef��٧�p�<�𥄔�:����\;-S⥩E��k�<�7�V��+V;s�.��g�_�<�4�L,�Q@2)E�V�U	g�W]�<���4!���K��$,���%Z�<ɖ�Y����Z2I��i;�L�W�<�˗9��e�)	�8��U�<	ǇRC9$�ȓlƦd���:u��M�<iUO
3i(�J4U�{;@�R���F�<�"��%G~]R��P�v�����z�<��ª_��۔��3H]3�k�<9��5S'$���X�s��MC@Mh�<�GŔP��p��GM�D:&����H�<�CC���k����>�x�s�F�<��B���V�)�hK���a*2�h�<aK8(�Q��$���%�#�b�<��������t���Xm�ʀ�D�<�AbD!V��`Q�g�Ta���g�<�T�a����ׇ��H8a����\�<��LM|�����u�`S�	U�<ٕOƇ%��a4hW�*�2$�d�Q�<��g�Nx��ED��U�t��u�A�<�7��u/΀��ʿ.e6tJ7Hf�<y�"-��9��X����
_�<�@���t8��!�Y.�dq��%�P�<�F�˟/�HQ�%@��fPD�<y�(@�F���V��������e�<��B��[����=X*D-�b�<	6�z/D�q�ҖjS�A���[�<a��	!��i É��F�fh���X�<0-�:��5����fH�U�<���^jtr"�H'8y��Z�<�+H!,��L��W��1����V�<��	�Hv����c{��q�&�]�<�`�.��Ӆc�� Y�%Bt�F@�<�p�5�,�p4�܄DhP����c�<Q�l�)a�:8�o��:�5���`�<q�&�Mʐ$�ЀEPبAu �^�<�`m�c�D��%F���ڲ�U�<�s-�1wg~�ÐkZ�yh%3�KBU�<aF�F3[{0P�f�F��M����y2���>��"M \,���r�ʝ�y����c�L�GzN�@b��y�'�1����uR�<m�e`�I�yb`J�A
�Y#���� �PV`]>�y��O�P������~؊�B㌀��y�a_�aJ�8�\�c��Qx�I�y"K�	F�����-�O��q�S㏂�ybV��-�pIK�H��b*ő�yR�CM�.�#��:�hh2�ޤ�y
� 0��$���P�%�O�v2R�I�"O�*�N� � ��"��#4�y�"O�x�$焟����&hn�qa"O` ˢ&��M/�03Û�r��I�"O��"V煏Fφ�HG?N�����"O�ţ��n��)(�%G
O�,�A"Ot�cEE,4x@5���	6�z���"O���w��=���:##�9h�}X�"OBܓעV1�V5���Y���p��"O�aY���!"�̰�׍�1��%h�"OH3fR���c�썎Y�~�2"O�l��JL�=��ĸ�����j��`"O�(�AK)7k�L3�I�5-�ҡ�W"OZ���Z�P����G��-�1b�"O@���f\���q-٢X��E� *O�� ��@�Rz�P[6�M�ju1�'��0�S'����\�.��C
�'b�	1J��;�4ܺd��[hԲ	�'�ظ��f�s>�P[d*I��s	�'|Z���ЪPn�jc��&?�4a	�'�����% *$4��Z!i@�X�'΁P�E��xlr�?/�:MC�'�<Xz�i��:�F\#���z%I�'¦��b��?�ҠBP��g8�P�'w��yGޯn�8��ƉXc�'+�QH�+v��Bc1z�1�'��*PI����v��t��'
*͡7����9!�֮W� �9�'����5hq��te��LE����'�F�i*��,�^m�$&�?�Ji�	�'T�y#�BL#FF�X�+��>f0	�'J��;��8a]�5��AP�9 >i��'tr��Ҹ��G&B�/]���'� ���֘[�(�Ae�!,z(��'p�0X#�C�Da��{��-o��9�'�|2��� �8��	�] *�
�'3vmc ���6����.�R�baR�'<,�
dDL��as��J�(L �'bX5����eA�Ђg%;��q{�'@�aI&��1�r�2B@�%_ ,��'��x��҄Sƨ���X'J< �R�';� !"ՂT���1A�a��'�(��e2KC(xI4K�;,a*�P
�'��y��mArl �h��*�&l3�'�49��a�
�D��G�K$�8Ph�'�@�l���"aW��Ji��'��xG�����6�O>%����'a2y8�'q��0`Ƣ)�
�'X(���@�z���d�Z���*
�'+���0�σ!�Z���@�[aD$��'�F���[0;��axV��!T�<! �'�U ��J���˚(#��8��'�Z48�!V<�VI�e� ���#�'� 5 ��Ⱥ�xɺG��@<
�'k|)`� ��FL�șDO�!�����''F`��ꞧVJ
I��`�]\����'y܌"�@R���CX<RL�@9�'�%���ֻs�2����~/�Ћ	�'��:�%�+��1:!ʌ�s2ͣ	�'�1�W�%ve����r�|a	�'q���S �9;��wj�*d�(u��'Ř��сȂ[Xr��M�'^��d��'�$�E��%h�����M��\�.� �'u�x�4����q��㟈M�:k��� �|:�I�a�z �W�	�-(%��"Ob�A�δ�X�(�7�yb"O�<���H$h�1˧GǓm�VdJ�"OrXCq�Gb-�
�'�C0�V"Ozq#���-r�H���JXZ"l���'��e!��&ƊNr�2�$˜g9!��=Pd	��̎X�P�b�(.!�$� 22�9�B�}x`�4�V.h!���ZjN��ƫ�|Z�G��D
!�]�O�	��IF�=�DQT(	� !����i�E�0#���򨒱b�!�$�A�� S/t�0�H#�ϝddf����埘2��	���T��,@��	� �o�<y�GL!Q��4+խ�+rKqc�L_U�<��J_����caC�{��"��R�<�q!Z�$= �%�?}]�����c�<y�!A�a���1�#z��@���i�<�F�Y�Q]����3X��r��\�<�c�� 4�X��NC�b�Tu�M�� �=����akB�/��Xea�T)*D�ȓ��XB��+Y�
]0#H�c�*h�ȓp`~<i�k��\�rUg�8
�ȓC�6%
�E�b�֭�710�ȓQjD\�5��O@$9�$�E-���ȓfe� ���
YƊQ��-#����d�V��AJH*=��Ђ]�S�|�ȓ �N�2%d<���DKЗ>����,�(@��+�� <��鐩I{s����P�y"���P�m�DF��I�`8��)=H�ɠi�<X]�a�V�/3RԆȓ(v\����͢	| Q%*�Qr��/��̋P��F�Ф�63�,�ȓCn��F��Ђ����ȓ{�n݂`�� �83� ��Q�%��q����+I[}h=ɷ�] ?(VU��<�F]�U�eKHa	Ҧ�=j�de�ȓsL��Yp� �V̓GN@�=�����N�(L%oض ]���B%S�]6��ȓH��T����@���hec�84���ȓ^�du�r�]��u0��S��}��cY�=J��+!iP�C��"���R��pC��?�+m@� ��[�<y���>>ݐ��FA��:�� �&T�P�qɖ:[G� Х�33>,BF�9D�43�bƐ0`����g�����c8D�̃��҇u��Ց�ߴ'��d�;T����E>V8v�J�φiȃ!"O��RW��(0ܰ5���Dh�mW"O���M��q�̡�2�G���H�!"Ox�qB�
<(��IFܔ&�	*@"O��jå92��LB���I����"O�%`��X��ac�,��	�"O�Q[q�K����Ξw���"O|8r���&=��0oD�P[�p�"O�I0D*͊vU�P�%7)���"O��@��U�%ѧ�<Z	+�"O4d"�G�ʪS���##"O�$-}sV}a���B�H��H��yb���q8�����@�ơ�C�ȸ�yBn��xr��U�4�j( 3��#�ybc��C8@�(0�ݷ8.�I2b(Z��y��?>"�X� ?%.~8� ����y��
��E�J%Cx�i�BF�y�D�R���CFA>$F���a%=D�� ��*P�VB�Q�!NɸG�V�hq"O����K�4�����M�N��H8�"O���V�
|h%�r	[��8�)s"O
����Zf����ȭo��y�"O��:ħ�yU��{lҴ��"Or\���B�1q���b�� "O~��o�r��'��"*�N���"Ol|[�gt�Txare��i�Ƒ�"O�8A��:�49P�c���^+�"OT5��E�G(�<�_�R N�b�"Oj��a��^zZ���@a�P�P"O�����L�*�
&.p��"�"O.�"ƣQ�`g��}�z���"O��A�!0��yL�,x�L��#"O2T҇�#u`�3��P1�J��P"On��0,ă*�zb�)�0g���"O��*-��/�̫���)��4+�"OT��[��$Y&f
rm��"O�l��L��0��G�%R�A��"O�9�p�J<;��H��\'~�V"O�3sNG*_�Fq� �+x�3"Or�h�W�h��U�a
.$�E;D"O�uC �K9a�����խl�i0u"O dB!�K/G�J�.�Y\��s"O�!�(���"�\0N��)P"O��3�9u�x8B�E�M
Y��"Or�z�/�"D��A�N���l ��"O�T���l���M`7��;�"OL�Ȳ��)|�x�K��m8�S"O���$ゞ|��q��Rs2��"Oȴ��A�N��9`ܐp���k�"O
9{�'A�e�2(�.\�)c2}J�"Ob%��� ��>����,
K A�t"O�m"m�G��� t�u?d��w"O������Hv�� G;%��Ab"O�-���6N}-0G�
*z�)��"O�%�@-S؜��e6g:�JB"Ol�b��I�tB�b�6!��"Ob����H�hk��;V*I(�r��p"OZy�­ gۂ�A�(�1>�X�����XF�D��48+ y0��.f�$�y�Ձ�yr朂J �p��읠'��0n���y�
���8��-�V�:�� A��y��ڍ<p�`T�?U���G���y�ڒNM" ��
w��!w�@��y�)��E0����o�9�F��-�y"�79�Z�#���Q���X��]��hO���A%:G���b�ƩX�� �7-!�߫ue`
E͂�:'K��$!�d�!TX�q&#�.
n�٘f��;�!��.�H�X�H�.Wx�Ha
�g�!���icZ�j`�|NNd(Ƶ-!�DG+0�@F�i1�|�1F�#z@!�dݴ0�^�:'�dsd4��s�Oz�=�������^�&9���ij�Dӵ"O(�Ч�6"��*P��� ��9�d"O:4P`®n�~����Ð�J�c"O���G�((�`��!���)c�"O�P��ʋ'��mj�!?%��l� "O4�Qf�A%'�F�ʶJ�}z���"O^D�N(5��y"C�C�%uY�A"O�I�&�;�<� 5�
-�̔��"O�l�#l��a�-���%�B��"O.E��DG
��ay�@I�N*$=�F"O� �;d�3!T��	'6y�"O��hv�-;���妏�C�Z�@"O���#�/E��<�ӧ�~���4"Oz��l��k��B �>=@�zV"Oh��&/оt)��B��v����"O:	�Qj�86.b(�qa	�Zj�A�"O����	�.p� ����&5����Q�L�Iٟ�'��|j#�ϑq�l� ��@5���3*�H�<Y�I)J�<��5�ʉ[K졁7c�`�<�f&..>�i`n6}xQ��r�<9i�?�|���s���Pd�Ex�(Fx�H5&xl��ګ�R����;�y2�V
 c���`���%�%�C��"�y�`H�=��d#S��%fp�l��aT���'��]�'{8e��B��P��R�D)<�4���"O�1��S'X����'���S"O�]��̘
�꘨g��	M�4�Y�"O�mb��  ^i���SvR<bT"O�#0��u��8	�Dݓv��"O>��剏5t�J�cs���gD���"O�:�a��}^�Q ��,���"O����j�S��F�`CօqD"Od��)A--\PHA �=3�L��"Oz�s�bב���h���7�@$з"O�)S��=-��8�r��!`�$�"O
�I��0FB�xY�bϰ[cp�p�"ON��@H�o$���a�~X��	�"O|{��ʃv��  ��9z%r�"O �  *iT��P�aƴ"�9J�"Oj�b��N����
j�"""O����^�@�낃_7����"O�D��ݽj�8�M(r
|���"O��p� :H���{�i��$�r"O^�b�R�]��!qO,T��"�"O��j��_�N�h� ȓ/�P�!�*O��0GK�k�60	a�C
X�V�S�'v��3� [�P�P|��`�Q�6�"�'�R�"f'R�F����a�G
�M�
�'54�'���y�����\�20�\#	�'}t���+[-����O�(�����'�P��4CÓG�h��T��&z��r�'���S�F�+`�z�I�eM$oJ�j-O��?1�y�g,V�r��&:h����J-�yr#�W�̐�u
P�8X̠��ď��y�&+�ր`���;|�LP��%�y��)%�Q��E���2O���y�Z�)�8yd���/9��Z2�y"�ɸ0.�� 4�^2{x���!Y��yra�5$����J��Љ���I��C��'����/L�CJ.�B�%��C��HL���SEG��K��_�]f C䉴yh�I��,EU|����O��B�	�G���WB"_�DEr�oQ���B䉺$��9C�/W�"��%�K�Or�B�ɓ/_$dCV��T��� ��S�@��C�l�b�8��Ӊz�����D+	P~C�ɐ>�f�*��8P뺸Xt���8��B�I�Zȁ��X�c�4��(�+M��B��1b����&�j�hPW #)@�B�/���3�Ƃ�0�,h6�A=Y�C䉐�p�a���/�����f�C�	�h��{�	G/X�,B�"�>R�C��0#/����+�)p �,���O�"z�C��.j����Cv��Dk�&(��B�)� ��1ɟ�?�p� ��L�\��"O�I���=H�#GH>,� c"O��'�L�|�i7#N�k)聠�"O��V�$ qB����CvYh�"O� Y5�W'y�롉J�r픴�"Ozx�1dN�$��`3)��K�A��\��F"��@�H� @C�(|�a���_�}�!�D�W�n�Z �4@��t��0�!�䅊g�X�X�'��Q�^K�&���!��F7|>̺�#V�.-���1FD9�!��Y�����&���e!n�!�B`2�<P"�@'|�ĩ��85�!�$a��� �/O�^����$)~!��A p���K���!Ժ!��>n!򄞙�T4��Gܢ(��F�ʄ=`!�̶ v0�"����z�a�_!�$�tmj�;Q��0]�Zň֋Ppn!�)����a�±E����/��5�!�Dރ]�y�G�H1L��Dy㨃41�!��
C�~�"��%�t8�d���p�!�d'A�,i�&,T�/$9�1�O'lL!�$	�w��-ADi j�rPep�!�$�S�\H�"%1_ �D�ݡ'*!�dJ�	c�9�q Z�c�dX�ET%.(!�䌦���R�鎳k��#f⛊g!���1*<�� V�5�~�It"#!!�d-TaN�Ղ A<4�P��3,!�DƓ&��[�LGM�5 �Fk
!�ՠ3G��Ä�[���ӳ�=O&!�DN�z@ܱSC �?I�����L.G!��&C=X��	��y��P�QA�J�!�;�~�i5�@ jX�����,�!�əOX��Oˤ����Y�v�!�D�	@��j�MEBNH��3��	�!�*�&����)��%	�eɶ,!�A�N��1��l� N�>�b�F�|'!�P�9�2���l��\��I�G�G�d)!���u�%�tB�5KS�* ��>o�!� /��K��OG�s�bʽ|!�$�$-��S����UCC�Z�f�!��?kG�,y"h2Y�jX ��ߡ<!�L.��B�E�0i��5 ��	�1(!��W�u�����584n�3V!���]�r	�㇘"q2鑄L8!�DϽ^�Ƒ��̛4��P#fA:I�!�$׻F9p@p!�|�Tk^hu��"OP�zS��2O^z\EDH�l�9�"O�!��N�|��HA��DJ�"O�,��n��&�b������	���g"O����JɎ+"8}J6fIF!��y�"OJ��d��-S��5EԨ:z�a�u"OH�K�'\�K
�u��ӧ0L���"O��K�-��3��|:��YKE�"O����F��<��҂M<`;>�r�"OƘ�s^j0�i�B�K|`�"O"�57#rt@2���j�X�`"O�` `�[>#��s  �z)ڡ"O|`�7N��7ґ��g�*P�5���'��LQ����.ձ^|�	`��t�!��2Sx�PC¥N�Tf�-�I	y!�I�:�X12���4Tp��(��	!�D�2��p�6���'N�)��ϘR�!�$^>t(H�J�� �U�!1��7L�!�
���S㖡�@`J�@�v�!�� � �Tn�"$�"��J�7���i�"O�[#�u�~���	��y����"O�r���6�h$���ֵj�~P"O@�d
ƹH�l9��0@�ɩ!"O�Ax�jLa4 �Ң�H<"�x��"O��P�.����А�¨R���S"O���O�������7!>��"O��L҆3F�q��C��c2�L��"O�,إH|V(�hU�� 09��"O���a�7i��af���+�PT@�"O��! �+-�X26�� �6���"O��9Q'Чt��xC�{hE��|b�)�VA�L߾V}��lɤ$�^C�	7�t�G�P+0: 2��d5*C�ɯ2��<��c��x�,z	���yByS b>�v�8�#@�eؽO>Y��,4)�Lڮ|�j��eI| �e��cS��G��6{	2��ᮑ�+C�Y�ȓG�xt��/,�dh�&�(T����]��� �!@l�H���d�Ѕ�*)�#���@�0 �Ua7{ a�ȓSrx�+A@i��5[m�5�ȓc+"��*���a�%eD)O����ȓ� Ta�[ >ر��L�`�fT�ȓZ���s�V�$Ƙ�p�H�ml����D@d�Ȥ�H� ��U�J� ��ȓ��hpS�L���gߑ2�
X����<��DT+�$1V��)L�q�ȓC�l�EAY�Z�LD���S���ȓn_@5����'��U� ����]��RdR9����|Ԁ$���� 0X�ȓAᖱ�RKѥc�)�\@��ЅȓC$:���B;(��H)�[���E{�'�ў�҇f�#f�zԫ���-EB�Q�<I�i-b��%2M�E�Ux�<�Ş=ci��!G�<��$�{�<q�(�+M A��g8A��4���B�<��#4uMP=�3d�:(�BψZ�<��a�I�Ug��-�.���U�<���
��0�A����ܘ�C�I-<�0q��J���J0XT$�B�I�|AV�R0��G��qK�I!��B�	����(߾:�|ٳ���0N��B�	��v �g�B1SZ��JGBʞ(�C�I �����=���CǆȖ[�C䉝	j��Pƀ8_nM�T�S��C�ɂ<GpHYh� c�+���f�nC�	5w��i�w���l��dj�!׻D� C�I�"p��脘g�<cC��!?�B�ɩ gh{�(ɦC��i�)	H�`C�	&��͐ JO�XvJ��a��)O%2C�ID��-r�VT1!I��&C䉄Y�����.�]�
�0�XC䉚+�j3�Ͽ:��bG��~&PC�I�)tDz��F�hY؜[7���.�C�I�Y�u[�� ��9�B	*�B�I���s�&wi���$nD&Ww�B��,~7�9�Q�N�@�Z���/e�:B��26:��I�a�#L2a���BN>JC�	(����f�� �Z���B<�BC䉽=.�tr�%�M���D<IBC��,x¢�X@e֑?��#ӄő-�C�Ʉ?9b���J��a�,7�B��1z�2 �����,�%D4B�)� �q�2�q��� r��D�(�H�"O� ���x�#�e���&"Ob�U	=^���7��QR"O
x�2�*u��I��^� "O�x�ā<
��0!���E��""O��$'P?�[w��;���k�"O(��b'���AVH�+8�+"Of)@�nI������t���iA"O��z`�J j����� ;ډ�g"O���BNϬ=ˆ�q�%��1"O�s!]�,��)᎗*}�Z���"O.��7�T�\��!c�Q�>PC"O.�s�\�|	�|CgA�!��r�"O�<��jT�,��)���=>qj "O` yr"&n�pm�p�Z	��c"O"��$`�-q�d��yܾU�"O�isaQ#����å�:A*�'8Đ�Pb
�-"�-I �	Mq��R�'�ځȣʁ>H�p�3�ֺGUf��'<���gJ/b�N����9>�8�J�'݀Q񷩝6��!��(�k,8
�'�P���:It���n,^ٶ�	�'2����hұ�����X��ܘ�'�xL�4�C�Q(n��d͘�^]�@�'dl`�Dξt��hj��f�H��
�'���C.ǖU�\H�cY���'b�]�Ɣ�f�]�)`�sg��r�<��=���r�6�N��T.Ys�<��MI'X�L�:ecB<	�V�JWHH�<��� �i�	��C��^X��J�<Y�J4h�Jw�ڥ<~x���C�<�b���εR"�!�YzegT�<I4��SDd=Xr��hJ���(�w�<���=/�%Kr�G%m(|h�T�Aq�<�	�0��"fIB"}ĨiRcIKm�<�s#�&0��P�Lr94�zDPc�<����7��0���cxZ]�sQW�<�d�po��`���&a(0�V�JZ�<с�ŭ.�L��'Z�v�P:�VM�<�5&�}������)@J��E�b�<	�-})�T4�(���G8%c�B�&s��`��^���g�ʎ@��B�?����< ޸��nŖn�C�I�O�<2%Q�:nԈ��%�-̈C䉍a�5��'s���r���*J�pC䉆F�!�F�~���nQ5C�B�Ɏ2�ЄK���E�uP�ʟ:��B��w�T�s�B��g���2��K8
 �B��h�ЈKU�_�G+~�a�ǁ	��B�sjR����Z����3kB�I8H$������.`�`��
V��C�ɡ ��@s`�Z�.Hq�o�5:tC�I�ritt���ɖC��M	��-�:C�� �@zUctWʱ�b!�/s �B䉅9�� eM۲ݔI`ƚY��B䉋0ޔU�!�8a���4��r@�B��4^�ZP�$�l�w��;�jB�	��������b��Pr��� >�,B��
����Ö	>�� ��.+WLC�	�j��P2�-՝s���a�i�&[1C� gx(��O>fC��s�b��z1�B�ɻy8�	��m[�F�<�D��'|�B��>2ˊ�)׋ �P��G½~C��d�>$���4D��a�SNNC�)� ��X@�^E��DN��e���"O�%��`�D+��p�FQ�-ܰ�y!"OZ0:v��hq���G�
k���"O�@���0>���dI�^�N�A�"O$a��扇l�$���*Y���#�"Ovp���S��,�pa�)y�8t��"O�-e���P�is� C�[p�ur"O��AqK�3��@9��\"{n]�Q"O M�b�� �0��a�H�k�"O̔�P�X� �ɱ��A6m�b�r�"Ot���K�o�6���N�"{2�H�"O|=���ۤ}<m"1�gf.��"O��z����u{
�B0%
���p"Of!����\�h�R�״?T�)��"Oڭ؂��t��i��G�$TN�`"O$��uDU+Qޭ	��� v@���"O@@0�&�ıP�N�{A���T"O.�cU�TM��=����//�9�"O��8$�I�:ɩ �)�@�""O�UQ0�S�6��� ��28q"O�]�(ް&�em�$%�����"O���ƀ�2|�����J8�4"OV�y�EX~R�r��B�2p��U"O.�֠�����i��v�0$�"O���eϾ]��*Ҽ+����C"O�P�o� �&�;!�*���"�"O>��0MM�>0�ǭ[�lslh8T"O%ڣ�A�\�p�#L[l�%"OLL�P#ݺx��1A�D�F����"OLmT�M���y�� �&�*g"O�t��Ŧ�:A�P�U�y�
�3�"Ol����_�*xN0��o�?�6�8#"O��R�I<X<z�׭F0H�8��q"O�rgaM 3+@)��ky�y�E"OZ@)�� L^�q�����-^�m��"O朋a���F0��K�݃6hꄹ�"O�����^J��[�-v�x�"Or}82mRN|����B#R��%�P"O�	�$��{n�ԩ�N��@��"OPɗ�U�rj���L��YҰ�2�"O�)C���?R&01i�" ;�T�å"O�PȟIC2�"!��?��i��"O���ԓ+������!o*lq"OfX�$k�%��x��^���JS"O6x�Æ�8-'�0 d��g�4q[7"O��q����c+��T����$�\B�I� }:��F� �fJt�_�4�8B�Ɏ���P�ᇾ�\�����x�"B�I$`�ѵN�oP. $)�4B����-k��An�j�ǈG.6��U�n؈DG�%���3�Ei�!�DQ���3i��.�:�ȃ*҉a�!�D��
���/ÔN��p����b !�$AZ�5���,o���D�	!�DG,2�|m*��\,@OT��s��1�!�d�S��(��e�I�0�נG�
�!��@d���ޛ.5T�0���93�!�D��*[��D�h�C�W$�!�D�OnrX�#�'8VȻ��M��!� U�|�o�!��R�$�){�!��k���a��@�Y:a�;�!��=?�V�����Zt�09�d*O�!򄇼.)$���.�dYNf�߸_�!�䒼e��8J�� �H�1S���,�!�� ��F�)�&9!b�M-��M�'"O�4�1DY�d���*WH��pl��)�"O6��"߹v���Cf 7c|���"O޼1R��#�J����Q��v���"Oj�rfD���\�Q��<E<�xT"O~�X�g�;m���pPBW����"O����{�l�;#��*��tQ"O>�s��P�*j��h�敹���7"O ��bd^�U|h=��c�U�<��"O
hC�@[n��I�̄�pnI��"OBbI�'Ũ@Z+�>\�R���"O�0`R×"`Z�f���T�d�@6"OV�gZ09f��Jc�X%3R2�"O�q�1͒|�` �%:#Zya�"OZ�y�.G4OԤl
a΀"����"O��@gmN$a���벭���l�)G"Ob]X�R�0q��LK�|�p�Y�"Ol��%�Z#'p��ړK�=����"ONMc&J#m}B���S�y��2P"O2���M	�#���*�l�`y[�"O��Lό����ªR���w"O��@#h6��u�Uup���"O])6n%QT"t��N�tb�T{P"O:�X��C�1t�@C(��}d0��R"O��BÄa$�����kNj-ۆ"O��b�����9��.t< ��4"Od̑�T�$X�4�@<0�|�f"O����(@2&��ti�L �Q�"O�e���� }`�h@j.�pW"O�Rh�	]�@!3c��{���q"ON�P�ѥ>N�a�q��8es�QD"O�I����tt�"պX�.�j"O�T`��:QB�c�!X� |��"O�D�(�j�t�S��z�B�P�"OY�ǎ4m�h�I��H��y�"O��u�^�:��q%�� 6R@�"O��S ,U��arjL�Ǯ�c"O�8T�K�aC�[p��4�z�{r"OT͹Qe�c������2�")�2"OxE��$ҺC����:� Q�d"OuI���YU�h�G���5�d��"Oƽ�oB%6J��4�Pa�݊"O�e1��L���yw4�����"O�E@��y{�(�!ӵi���"�"O�Ą�a�e���s��Mش"Oh�ā*-$����u�ȉ�"O�=�d!�&R9���ۨv�$�Å"Or���%(`�Hd���EJ�<	u����\h�OA�3VP躂D�M�<9íI0&	b�ɗI!�f�ʕ [q�<ɱO�>N- �-!%[B`Ӳ�Cb�<�э���Ӑ`��\�"Q�4�Os�<���P�}�@G�PX�1�P Cn�<iU�N<e�8�c��?>x(�+�l�<i%���g�VMhK#['��*p�g�<����x���2k,�d�18�썆ȓs3B���I9Srܝ;R�^- �^���q� ���W0p�8�SmD�J t��ȓ.I�@ Q��&q�ՠSX4���:5� ��@���Ы@.#o*���8.N�A��@� �1�& B�
p�ȓ	�B2�� *��!�i��3
,��ȓ�"X��� �@f!��,���ȓUI�!�@�i�n8���ΞW��H��S�?  ���M56��8��-z�,"Oh&H\�:w 8Z%�W�@�"O���֌l-���򋊶)k��`�"O|�A*�'b������s~,�P�"O� �@n�5��X[�G7��գ�"O���hz�xA�F��/R���Z"O�$�V-@,=�8���kr��P"O
��$%L2j�C�ʉzoڔ�V"O\4ڥ���Dc�=K�L�"O"��aj�1d��BԳ_�]@&"OT|�PM�.�b�遄��.�2a"OZ�iЌ	�v�2�ʫ,�&Ċ�"Od�"p�ZW�� �"��K�m��"O`II�����X	 ��n�,����tE{��i�5A���*Ă�5(�Jpłp]!���PJثh�S���4čK*1O�,��ɏRnhH`��U�,��d���G�R���:�$M�(���{sf
";-␪��D�u�d9�O�HY�*O�	=��p$�]�94�̛u"OD�s(�<:X!x��|L��"ONt�m�hQ����N�Y@a�*ʓ�?牝K(���R���)��Z���B䉃OB��U�])���#�2Ś�O���$G�`��2eÍ��`q�Q�M�!�^�t/^̋F�W�O� XYb��=(�!�$�#+�Xy�lP#�$ԙ�&��!�DEP�Y�х�k��ȡ!%K�j�!�d_�a�64Z3-�J��YA���Qc!�~���s�h�E�` X�b�5pD��
O�,� cJB���H��368�x�"O�a��	\��krX�
��q�"O��iR.�%	�AFl����qc�xr�)�ӫ_DK��.N��a���,�B�	=䴽 �aض<�v]yC�ݟ5BB�l�)�G�:N|�5�[!YMl�H������?Y��0;�iC�+��=��)�%[s!�R��H�פ$���JCHO�\[�yR�I4Sc~�ת
c�"�0kZ�=�<B�I������*�;�`�%y(�O��=�}���M/^��p1��h�H����~�<)`�)0��^�G?���.���]�=�۴��hʓi$�G�f�����O5,9� �'y��'6����u���^1Vb�Pf�;[~2�B�Q��?i�O�)�3�$�
9� ja�b�����I�PO1O����J����
�h9��%��&O0SX��>�O��M�*9�ȂP)�[`��H5�'9Q��po�*���`e�;e����e4���"~�Rʃ���LaOE=.q�re�<i��m4�	Q�%�}T�;懞 �hO?�I�9�+U!�&���U���b���	� �=bbJ�����R�B�	4#fb¤R=��Er�Ѽ2����$��D��H���f�F.O((��2�g,,O�<��
� kb�SG@g���#��K�<�Cd�%u� Iƈ¥d��1'W_�<�A��gҹY��� A����ma~R�D>�G*�i!�ς{_$���H�
����QCz��kS�kI����+֪9|1��I~�`�r�JЁ_��Ƞ	s�G�RF�	���>��R�xs�T<^�^Qqc'I��%���T�I�}��qKS۬]8��c�NFH"<�y�	�p�'(�9cJ��[)�B��Ӂp��FxR�)��M��u�! �2R�	hU�_��hO?牽N
q��Q.Y������$l7mF�(O?7� b�Z�_��`TBTb�ڠ|���x��'c�z�gL�?�V��r�/��-[#a#�yR/��1��X!�@��Ox8k�I���~�2O�c�8Ez䄈 ����"̂f�#��]�yR)
�t�=�cH��"�>�8����y"�D�3�0���I�o����׵�y��'N�*�RZ�:�V��b�0FF��T�Oӧ����A -��-4i�I�W�{x�~"���<���ߟQ�#B� xIF��t�W�<��W�EذI��k��Dr$F�<K<y�O��GzZw0޹��nƉO��4�"���I鞔
�'+Lus��S*H?�H]�R�F䳙'T�2�T�D�MðČ�_�(�Ku��y2��1	S|�Zc��I BC%jW'���&�S�OO襋W�޶Wxi�3f0Kl���'�iɀ�"|���2F
#B6"O�1�eуjer���	ĝNwva����(O�8�1��7N�p	�ux��ěEQ:��t
�u��ɓ�bފ�e��Z~����e�
]h�HƼl�
�B	�4N��D|��Fp�����zp.Ĩ�TA�C��4; B&�f��1A�gn*C�	� ��hwH�}7̀��\���B�I����9@�(��e��f�k�X%��'��'��y��Q"<ApL�r�ڶn�8�L���y"��%]�ҥ�ٸk�^u��-���y��ܙh|�"��]<0H�τ�y��ט1�����L�S�2T��MS��yB��!t��Q1�\?Ff$���iϗ�y"�Q�Yd��چ,P>~�,9���y�E�,1W��ȢD��9����o��yR�+
~�|õ�F	46�X�#I$�hO>��铀&��t2�լ6��	s�84�!�� aOzhSG��7C�,�я��]�!��PQ Z��Q7ҠÒ�j�bO�U�Ɓ�|D��P� hN�b��'o.�O�8p�c�'��$ɍ��=��"OJA�@�$U�f�	ޚ����'S�'��)��x��0�<�}QÒ�b,���'�H��FH�g�\��V�H�Q�N,k�'���)�8ol��SشJ��:#�)��<�#JF=c^<L����=}�U(�b�J���0=�@�]	��8�!I*?Kb�* I[I��p=��k�(�&�3�&�M~8x�-T`�4'�xҰ�]�l��	U1d9��3�).?ى�ᓣjx�CW�׀akT	�� '�C�I���<�I�a�*�{�ř\�B����dPU�L�'�\��5��j��"?A��埪�� ��3:t��	ē�h��iK�'j�zB�S<P�Yf@D'>X�c����y��A
�H-Q�h�7tI;���y��K����ʤB
>e 7�3��'|"�	�<!�D�63R�@e��6V�-�2�PO�'a�tOކ?l��k� Ll6p���.�yb�$�H'D�o��3P �y�I�m�树7c:w=�h���I��M�y��'�Ի��Ǐ��"�j6w��
��(O�,��ON0��P�m�I
�M*"O ]�6i[�����5��`�w"O�ܰ��	�<��!�@F˪�A�D"O�1�Ԇ�0	&詳PN�c�UP2"O�=���D,�M��m��.����"OB�w`%U�=�RF�����D"O�� �GFGhԣT�7.���)U"O� ��5�R?_�֔HG#ͿO����"O�p*�f	�\	\D�#e��z��5���'�t�?��
J�Y L`��ƉS�H��Cl�<!Go���,����Æn�v-9Rl�d�<�|&�e8�m�(8bE!�]�<�Q16�l�`Dθb���LZ�<I��)�Y�.�PQ�#W؟|�g��1���
"__rK�]t������e:o8x�d����f@8A��o~��nī/�pX��N�����j����I7o�T=f��5D|
��ȓ���T)�	2H:4�bV"Ot�jE �l[�U@\DD5A�"O����ˑNj���mN%A�h �W"O�4@c��d�Hͫ�̝%q*��!E"O8�( ��&F�\E*�l��" `�c�"O�����u6�p�e;4r�q"O�����:,u�n�l�P�"O�]��B��vA�7cY=2�:�b#"OV$��%�9�F!@$!����� "O�t��dT�g�$S�R��AB�"On���e��g*3p�����Y&"Oza�h[�2	a�H�4�\��"O2iR��N)	܄m9 �� 1�,{%"O0��Bˌ�~hh` �(��p@`"OD�p`��2K�	I�շ���q�"O���kY`w�<3�	{rA�"O>�!F�Уm��ŪQ���p��"O� 
F�)=l�<ۖC�3�D�ˁ"OH]y��I-ܲ9:1�ʝPy�m��"Ov��Vi٩>���;A*W�S9�P�"O����X����r� C�<X�%"O���,��q�
-�Q�M����Y�"O`�¢�� B׮P�jn, �"O�X�V�ײ%�� ̓W`h�S�"OR����ǼP{A� �.MS����"O�(�jPE�ي
�!~)
�q"O�AkV�=ap@�tg� ���"OD�b��X�\HyA)C��B"O�a��H7Lv�Q��A�:��"O�0�#a"ݞ���D%-�Hp"O
��O�%�8K�%�>��ܡ`"O��s*��	��m���(4���d�3�-�sI�";�����5x�1OQ�Oݴ|Nʽ�G-)�^��"O T2�Q4R�����ԃ�"O�����mWΠx�@B � ���"Ot�S@�Of�ږ��5z�V@)�"Or�s+ZT�LrЮ2C� 0u"O���a��L�^A��	�2$�%"O.�����5r���s.�T�~Q2�"O|$��`�!_��UB�X)����"O8҆ I�&�	�NI�L*���E"O~�Q J�@#� CM�/[ ���"O��OC�	���:LŮs$����"O2Y`���?P;�xULZ�:o"O�E{.
�t�(��+�62�2�`@"O&Y��٭�ހ��c�q�0�K�"O^y�5&�����K���x9V"O��,AѠ��`��P�ͳd"O�8�(P�j�6D��:�,,�g"O���B��Œ�j�S�X}��"O ݐ��*PZ:�;�荟2���w"O �bdD�`��hy �р>� U(q"O�y!�^� ��'b�(q��"O� <�V��6��V���pl2�"O�$����dP��g�βg��"0"O �����<%(y{%ս!,���"OpI#��=��<,fl�b�\/�y��	yB�(��_*L"���$P��yR�B�a��e�=ndEj�`�>�y��\
8� %p�Y���3!��p=�׃�ch�� ���ZU'�0;eā	&KP�PnVT�ȓck萣�i9��A7!*8�$��QAЪ9�(���&^��,��DC�w����$��Vz�C�I�nj6H�2c��p7ʀ�h��`����1p��(骅Ӌ�L<����
7��A���="�`�! _(<Q���

�\J	Y��	���H)i����� $76����H?�O��g؂7,������;GJ��`�'	ؠHC`��� uf�<���ц ��e���'R���Rh@n�<��咚O�Ex���	dK��pnIw~�*�φJA���jT�LB���^���##�NQ�`d���Y��B�	�@�v,����OS`�cB�tPtH�[���ɁW:*$�Q 6�3�D��5��rǄ�+
��q2Q):Y��}K����>馆�g@Ბ���`�"i!d�o�F�Q�fU���@I��R���'��HQ��6@rt�'|<�p,��R��쩂O�mO��
Óa���*���cu�E;��?�5IōJ��S�̆�I���E]y2o��f,�#2l��wf��J�*>Hu�VbArd���v~"̈́1����'i7L]B��SY�l,p�f?M����L�/@���5�F��?�4�^�/��Q�r8�����m�.	"F�K�lq��Łm��ዖҡcF��QT踎��'U��
�<nb�����(]N�dbF◂��y��Fڊ	yT����,lO�DsAA͇@�"��̞�r����Ow��TP\�,�Q�_6p��D`,8���ٌf����0��~�����e�2� �C8��)��[�dG�$��I�?́0.�*��G����EP>"����%GZc~(!S�m�O ��I��[z��i&瓰!�����[@t�c���>�P<{GQ�'P�E�'|��P��[�IE����ȁou�>��0���~=;7c�8��a�JF����Ipq4��K߄�~�z����>!D,����bB ,ӂ�a�F��tH`�^?�6���
ZV�>E�/F�)#=k!���җK$ ���°�U�PJ( i�"x��L�*)
�ɀIY����dI H�0`�V�-ن,����z��m�w���f���H��?�G,��|�0X�)֚c$���y��u��a�E�5$#hR��pa��db�%�W�|E6�5*�H� �ʲ��5(�X�P,�33��ݣ�!�6�:V�H�c,����u�*`�P�� !{ݤ��Gn�\A<�*v�H c ��}ꨐ�%�S*`��a���E����1�@Z��S�9i�'�� @���=8k��I�D����A�I�f�4ً�6��A$"�Pa"��ؖR�0����ْG%���&5g�QQQ�yD�ۘQ
}b3��T�&��ռ[`��)c>�	�'���~uX���T����?ܬ�t��0#Ɏ4��4�ɗgH�%	�%�I[��`(N�S������N9� �D�`��)�
4�`Z��Ǜ%�� 8#!�����Y��xb�XF�ȡP��uPZ񠵡wQ��,��M�\(él�X���A!H���A��](m(�awE\`=�D陚C���Õ�R�h;΅H E�Q�4A2�_=^�&I�&�݊[�,1U�S~����\qZw_�(	��^�M0�PҤdY#S�����2y�<�㉧IE�eA2e�$f`4���!E3�L��Dٕ#S��"��0|�R�&Ju>h8�J˸A����"�v�J�bcǣ<a'C
2M�]1+͜D��b�P�s;X�`�6�����h�0����i�X@6��	[��L� �^0�Z�G[�'��3fbW*'*�ic�C�qq�m(��a!f�*�w��e��
�`�`�:s�6o�DIPq�[4^���3vȆ-0ONU�����q�՟?�ʦmک&4M��C�5:n��!�C�W�@H�s+4�S�׽�<����M�2�t�zעC49d�Á�;Z�l�'f��aK��3	a1FS,��H�VF��!� ;���6i ��H�mmP�rkA�7  Ii�FR���p�vfT�"�8S��.r����"��d���2�����g��*?�-y�&K)p��S��L�/	1R�`�NLYj���͟(N��ː��0� M�v�րE����R�Y;�vY �(Ro�d-�ʍ�(H���P(ք3�2e���WA���ɀ!F�}B �2Ԧ�,0d��Z:�	!7X @ё�I��Y��C�=$h*C����a0m��?�z�oD�RO �w�@���;1L�%�H�juDќw*ػ�`I?˲�*2OE)QJ�O?Aϻ���Wo@60]�p¾���
.x�ٰ��A56W�P���ԙEV� �|�'&���K�k�@S1�a�����I�欈��14:A@s�_�{~M�T���N��0�u������䍃O~9pԊJ8YD�@g�ɺMr�րA����e q܊����;�n(*�\�H8Op��ӎWD�r	y�V�2�tL�����I�@�3w�C��1O�nY�/�<����,9��lW7���	`@�����
SS�Aȃ�O�5�r\��X�,"�E�Y�=Z�LQ�'\�����W[�e���7�xH+�e�/$���M-HB��cTE�)��,ӀD@X~��$T4�	AȂ4����		3q���p%�d�S��Z�t�Z� H=LpU��;Y��}1۴]H����m2� 2W��,aL����z���#� ���h�@%@ӭBg�9�g˝>�T%�C��P$�.�
��eΟ
I��A�G��f*��n�۷�R�v��ȡj@�Ͼ�35BE*4�a*��Q"�r<�`��?V*\�Rs!�$Ge]ir�G"κ�#%"+7��D�a�4�Ш�t�"�Q�W�~9ZI_J��
�/u�mE��!����J�+�`�rg�ЦP�n:!i_O��*uǗ�V@�����ɟ����e�X<Vr-R�Dɸm���A�)M���dՒ'�qz �1td1Q�o��Z����'�#��@�	_d��i��[��Q�g>��eV?;��]��o�r�A�VSz��C)��[��� ���)��ԑ+�L6L��R�n�<AwP�6�&a��(�8n�\"#��"p����S'.�����&ϧb<d(s-�9#�E��� I�a3���"0�ܠS�їh��raę4f2vrs�;'�a��
!L�}���H�
$�p&�#VK���-��+���t-��je��*�9��)Y�M���&A�TN��b�� *��	�$m #/��1�d�p%�U+"�&M�$|��IПO�� ����7'�|�$�b�wɑB��@�"^���D�Eu ��4+�.�����
�D�x��u�ӛI������j��d��[�*��T��(����kʣG�r���(N���0щ_:x!�d��`��̍j�^�����"�?FP顎�<�Ο�$� x���w��Qۇ�&|Ap<YƑ/4>0$hRLD�Z9� �7D�i�r���$�@X��γ|@x!�Ƒ�05>4XB̤��kR���T��Fk��\�cIW�N�vӨO*P#���O�]R$�Y�N����7dk$���$G��A�*f�b)c�Ǉ�'b�<)*�C��xF�׳e~p�S��%�t
�݁f�bvF�!i�b*�#F��5 ��9v`�Q��
j�!Q�� p��#���k��� ��wOZ 7MO;pk�-	��;b�	dĂq��SwL�l�D�Xc�.mV�x"�DM�����-č7�����E�%7M�(:�;j�Z�8�hȭj[�Pb�O�]����
1�l���<	�Ԝ���	�MSQᇘKܔ�w�X�80P1*��|��\w��7�	�8A_	O0e23˟:�-����<�����S$6�杋@@X�h�� ���<���܄�P& E�C��b��ҚH��G�28�ay�e׍� LX  E	y���3���f]x�p���X���-L�>�ey�E��"\@Xu%��`t���I{�Q�gO2 7��ӱ���G��	�<ˆ�H.�p7����!GR�����&�zx�C�>6S��'�9�n߄T�$X#��@.i� s��y8�/bӦ�A���+��8t�,����A,v8�	Te�5�����\�#���4�Xe��)r�qAi@9���	R	Qn��a�ƚ�|�cO��8=�� ��!���D�ĺݚDd]��M�t$@�Fq a�F�m�.	a��[�d��0P��1`��O�l(AO %gޔ���(6y�Tӑ.��x:vؚ>nv�3�M7�p q�%fܘ��3��6{�\Á����M�%Z�K��;�&L�>hM�{T���0��85d��(� C 7��Ol(���>l��P�/��Zq�Ja�����΄Uäa�r��*̼8q��^�x��d��[�)����g����w��VƠ���Ճ^���قn��x�%e��LJ^c�L	��S�SnIz�f
85X�q#��U�4�<5A%R�f�l�fص-�V��!L56i2u&Ȕub+P�H*pa�pf1��)۠�;2�Zw�$���F�&o�\Q�pk��c� p�&г����׵ih���A�B�,2b������ע� |I@�L#b#0ݹ����ߝ�r��8�q9�ܝ3k���'\9.��IP�N��)�6O�b�@9�u)�D�3k�EX��x���J6𖫍�&��x3TEHaw�ͩ�Ēi��dc2M7F]��p��[�M&-�F�4#�ʼK���B�]Q��ܖ��XJ����<!�ܔ��qq���$U
��܉���Z��
�۶EuF-1��4W�`�)D�]	K^�e�UT�i;Ĕ�@�Ե�dEZ�CxXQ�'7���Ŧ)תR���y�,,9_F	Kd�K	.�#<9�!6&Z�r ��]y��z&��T��"V�y��B2q��ЮGJj@
Ph� �13���T�pkȀS��H��>�O�:��u�ټlo
�!CH��� P��;^Ґ�V��7�F��'���*��M�ml�	�E}��P�s���Ъ"0�Mb'�ʭ ���x��~�$J \�v�qO�>{������Sf��.f�Ex���s�j#�_:cl���ڇq'��RWJW������*l�m0�_�v�~5�U�B�b��( ��a�A!o+ayb� t�`�f�*T,��¡]�w�Bu� #�Q4!8W%�8͸��'?^�Ha�ӂrT�ȓ�LKt�RU��#T<c�x���+h�VlZd��{Ӑ���K<}���%�=��m�9�EAu��N�FI����[�|�� 
Q�D':�q��ӱ�&$�Jĩ\uTe[4Cs�(5{�j��y�B��E���[����Y��ӝ/�^��ώ����� -�O0��R��0��,{�I�8���A�d�+�N�z���Sज़�)4��e�u�	�7Ú�\���R�'�lK�  .�R!��.+s�a
�H�DH�!@�v��n9Nj
�p(��-^*�u"�^W��4�2	� �bH�ok��
2�U�M���R�a+ax�M����0"�66�C�E�40�"æ�-d�	�D�BA�}�cO*5cf�"��٣2H�t��&0�*��-f��2A#��CC�iR0���p��Z��H;._�6Z�A9�=?�F���:g�D뢆�9j�T�����q�%�0�i�bԪJtH8i5HP0h9 I�*�j�Ƹ�t煑S�1�6Ck����ˌ�Ip^)ŨQs�$T��h��S��h	���<Dy��O��p��H��?�sц)�p�( �Ϧ�B�W�?s���e�"�!�R-lDP���p���W�M�r�Rh��kU<D0�jȠ���S/hL^�0@a<�	'\����e��f��j��
 #S�IB�Ϗ)]&f��=z�� T�mv�|�H�/�X�	Y?=�T���_P�I��φ�yY�M@�<�%���8�b��!���	�(��׃���f��П�2�*�&=Kp"2�P�Ylh)aA,'��X��A&!��ץ��*�J�'>CXz�Q�BGպk�ˉ**f��%�"
���L�1n���� �P?a�E�c���#���B�WB�GY�g&ʈ���.%{.d�K2\g���Ї��2X�`�BN>�0��+p2�q��ĳ
*h�4���[g����'	N,����J9��'kѐp�)�	�7l���.��x�a0�O��C�f�=� ���P�{� yu%H�7m��3�N
�{�"�I�E!`��� � k�u�S��`^.ڐ�GJ8d��'�:�1fŃ#j��̟�q #l
�
B&���&�{&h0;��}��i�0dhx���b0S���7�݅@(���f�/vkEO�|��}�$CR��5!�g�;�&8)A	O�b�d�� x��ۡ������k����mI���t,�g��m�4�T��R�ʔUDfUY�ѕ�HX뀮T��OQEDV�f�M����X�����QMxyqV͑�^d�`C�>e�4��5��-H�r@cv�<	1��C�'�hM���z���w�;}���-�M�F̛�|p��WI�)�f���芛?i����#Y�������(y����3F��?�h ���ɨ*�l��W�ʘ:aB�F!\������������3�Ejs�E���rG��`yR�'���t��?��i�l�8%�갓ϐ�O�e����^_&-�GS��|���QZ񼄃%e� DpDh��OI�u�
:]Y.!L?��B�t�z��V)�zM��@J	_2"t��)5�b�`�V�n�����C�A�b�C+�*�jQ����]6:T.Ǩl��(��=����'@"��ɏ��]���J� XBdR^�U�*nE
�O�;f��
�jaՏ��S�r]�F��0b���j�R���8Չ�i��o���J��
�8ٮ�eОEh��X�V���
��jI"A��'V�0��	$)t�ȸ��Pa�� |2"�ͻa���@��o�a
��W�!Cޤ#V�O�1�h5Q@��$U�x:��:b�����O�EJ�)�  G*H	�Õ_6 �ҌΟB��k��
PF��0��M�$��'�Ԍ�e�8pތ�iăS�-�q铂W0�Hwm�F::�R��<-PaU�'ւ�I��*�m�ÒxҬ�>N�jy�I	�%3�12��]8��$$C��x���"v�|9�o��^ֺajb�	t�B*��V1q�0́ ��8� ��C6ta��8�a �yb���9�<h[7�Hx�����J�n�*��`I�Veq1��O�<�F�/����7�З������j� ��p���])���.�j���얒J�ifO0r_$��6A
��yrD��-�(p��&�z�ۆ��SBh����S�b@�ah�8o}�d(͟8(��c���i�"�J�O_�JkJ��v��&�R���ɰU-�y��b�
e�i�j[8��ա9)2Ȳ f������ ܳS����I�l1��]}��p&��1h��?9�h#u�}����A2ܜ�Vnځ@Ҹ�@�ջs��7$F<{T��v�N(<P.	�?@p�ru�;U(	7
Eq�KEȑ�:"9�(��j���O�l}YV�J�eǒȡ^"*��!L�o�<q�VZ��
��,�@J��%xz�б!�-సP@�OV�F��O,}����)<�.8�GY�Q��e"O\�UC�-s����IA�T��8�i�n��P��.��� &�x�dQ;\�r�z0�J.O�y���	���=�d@
�� �R��:^F�Ԋ %�(6jr�j��J��nԋR$.$�����u��ucS��!c��!�a�%�	9%>��xQ�ݱ
�>A���)�4gl�2��>;y�pX�(!򤅸D��\�5��.m��I���e`X�S4���]�����<E��'׶Q ���IYR�
AW�l�i�
�'q��Y$+n]x!c�g�<})�'�&!@A���0<���$��#&H7���m@-sT���D -rV�I�ٴ�aX���x@��F�a�}��J���95O�7��kGL�\	���ȓ4��X�e� �w���b�Z�)�xu�ȓ��X�!'�� �(1Ùs�Ņ�l]�ui�*7��(��愸c�����Uvl� �9v��샤�P4����n�nm�6BN�A�̊� �n���X�6��� 9ײ%�n��pVJ=�ȓ-�f��O��x�F5x�dڂG�J �ȓ>A�$�ъ��2�JU1ŇѼ(_���w�r�V�T(jK"͐�	�yB<���hl������E:$�P�Y>9�ȓ>a��i��ެ���1�@!,��ȓ1�<��%P�(;j@y#@�<0����(���ӆ��Ȏl��mCa;�)��;D4�;�
�3s����!n�Xԇ�S�hBf�����'��"I�]�ȓSAX���]6�RT���ͦG�n��122M[��*+J�ˆ��?pЕ���@�aS�ÅM@l���:l0$�����P��
`�lu�l�1f���pXL��clV�~�1�#�d�T��"2
�/��^$rs�� r����	���	�NV�lE�$Js�O�`$L�ȓ3�D�u�ZTo�E��`��4� ȇ�aoN1�ūͯ"�aX!��EΎ��B��{�F�ccX*P�\XDهȓp����IF)V��K�Z��)�ȓ_�Su��u��h+%mT�{�L�� ~���bE��j�#���s� y��\S֨�0�	�*c�8 lI�4���ȓ=��;D��?K�u��LG�f�Ʉ�#�H���l�(�*$&�� lnl��Cb&�s�矼t&�R�/��D��ȓ���B��C�<��IZń�E�*��[�X��'�(���N%e̽�ȓ9�j�f��9_t>�h�8&s�ȓb��lhQaR��>��1G��1�x��9Ld	���/lӺ Rm�+��Ԅ�S�? DP���[�&i:���[k�q�"O����R?��5��)ə@"źp"O�Ar��Q�ѓ�"�z�2�PU"Op��Ff�7����E�m��"OC�D��},�m��Oߦl6*�"O��K�,*o�X�AN=oleҰ"O;$��REC�GH�FP�l��"OtI����nL���LX@�i�2"Oܳ3��ao�i0k#E0tA0"O�z��D�p���k�IP-;q"O��P��U� �j��ʅ�xr��'�ؤ�R�G~ ͘=�ђ,E(p||�G!��yBk�%mU�U�e���"k����@���"i������}�D#"��ρHS��R�� +�@21�EG�<aV��`a\X���U�E���F@��d�@�6�<Qw��c���'�@,�1mP�:���V4�fD��'!��d¥W<���k�������/Λ,N*@" ����-��	 ��y2wÌ�4|���޸#\���1lx�p	ұx�|i�'�&�'ƍ���,�sB|��R	�'�, ��J0z�*�B6�ŇZ���	�O<]�Ռ�	�������B�^�}������&�(ޘ�w�`�<��㕈I:�3R��=~�-Z7�OJ6J��ăP��?�ӧ]�q���|&��(���UR���&<��p�-I.2z*�#��'f�@(G�+���nA�8=d$a3�S�
��`"Om� ����l�,��ƒ���@�'�����?!�X��ÓE�r�0��8��!!��ަ�?�F�R҉���ȘU��x� �{y2�S�#g\=R�CE�5�D�2օ�ܖ1��j�_t�;���v~rŕ�,�Ġ��hδ�9��SYd�Ā��R�	�nru-�t���Fˌ�?���F�V�1y��8��b&�gr�P��e��MM�SV�]i��*�Ii]ҡ��9Mte����'Lpi�5��*d/���1��'d.fQ��lH 3�2��r��˴eb�"6lOJ�a��g@���2Ɏ��+�L�1*k���D�I�}T2�i��p}R�]$`H����	cJ�5z�F����Mq|d�%��Q��4*�ϟ��0<�+ �(�x����y�����<q��؆�Ӎ`�2ŀ3�T�C����lL4�H�,=�R)jT��>r�"~ʡŒ7JJ����BȐf��-�b�-��d�#�^��EE�_��L�fi)�'g���R�AɅZ�*�&���)fK	�'�T AE*va�)��^���	�l�*�8��Q)"�3D�4�����MR�a.��I�	&�����܄����"O�7O�*�oA+���K�̜�8���Ӓ����HJ~������$��v�AF-Y7s8 "�C��`�B�W�fўm�p烠�?�MF�!�r�)�m�5	|$<BP��b� rȗ�gz��R�l9(Q���i¸0�'��PѦ�ҥK��d'�T��c�$I��p�&`�˟�B�\-t|�-��@�8��*�����r��1W_�aD��~��X���\,vx�13%e�@�>����
���b��Zn�x@��AM%Q�e��J���Q�i�"��������x�L*���7,���P�O����bn��b)C�Ȳ'�� �g�O)�b���V�0x��*�!z���2�l	��1!����wb��T$~������ێ%�������~���U�f��N$2�I&>�@�)
�Oh�%�$�G�:*��!��d���ЮҞ	`�o�X0�ɣ�L�|�E���v}H��#=(�pO�TX���7-��� pB����r%_��i��ۍ�M��Y^����N��M�t�G ��[f�W�'�"8����(f��!֠�f
�)a�fT���Ū"�f~�96`[�iB��'��2#̀7�u'J]s�dA!c'�4zQA��}b�ï��v~��	3A���&��;�b�xׇ�2|YI���~e%�s/G�sw��1��8����V_+uG֐a3g�?�L˓|��q#fF`��u�A�s3���g�3o��a4���?�!�$?J��)�@�G�jƞ H��sL����]��dh�f�I 2��Э9�8���8ӤCb�M'�y��J�6(
��lؗ#H�D��C��P�B�nǊi���j�d��1$
	7*��)�x�Zw��h��i=�(p��	��$BO��	�&��L���+ (.��뀁X�i>�0C�K}��]�����u���dK�9`!�W�_E���A˴A��Cװz������@��D�4!4h�Z�o�9���eǟ�?���+t�N�%p�ɢO��[q��#�<D���b[}��z��	:5G�
7�T�g��;��KF.E�%{p4��%�,ٲ=#��^9a�D|"���I^P�I�s�CF��'h ��%�.Ҫsw�߸c8�\v�[0"�:��gV�2|�a�C�>I�I�<�����`��U�=�`�XF��uړ�I��E�?	���U�3��R�e�O��dɒ�f��B��Y��XJB��.^b�@�Щ2`�)ҵ����CSA
�Sm ���mH��h���<2��X����h�vdJ�E��[s�?����ɖ��*}����%Oe�h����[�R$���̳.�T���l#t �˥~�0DR�6,�W�y�˂'AQ��@l�P��S��@�6�9���L��͕�;���84�Ü!Ly�'�Z�9&�#_�4)e�V5z4D�L^�`dj�&��W~`A�����衐�Hfym~���P���v@Ra&���5�*Q�t~0 P� ݊��1MA���j���w�	p��h�B�J.sw $H�眂ـ��a� ��j�f�{
4-jf��-/�u�u�U����^�_Pp�ƫK)N��L�� $A�������5o�����M]���RF�����N�]�ryB�i(Ƹ[`!1=��M�%��MF�Ţ̻4=��&]��s�ى�o���09��;W� @��(���X8��nBf���S%� 5*��̡��Ű�4 ��b�^�0m� :r$�S	���E���DA��ͫ�:u0�`��L���ME��Ơ�1y9�f��D���EB��Ţ�1y9�f��@س@�4��V~���6��/޵�0�K�;��Yp���9��'ն�2�O�8��\t���8��'ҷ�<�B�4���a���{�K��cSD�rw����f���q�B��fWF�rw����g���y�H��m]O�x{����UX�pv;�ỉِ�D�UU�~y4�bǊ|ؖ�C�TZ�~y;�ġs֟�L�W^N i���u����R{
��o���O i���u����Us ��b���Ee���y˜��T~��f���Fn�ֲ�+yԳ��g��u�0�ն�(y۽��i��y�=�߼�&yٹ��o��q�6�ұ�	������UTt��4�h�x������XYy��=�h�|�����]Rq��0�e������m��̩��]%6�U�C���|�i��ɭ��R(=�R�F���{�e��ġ��U->�R�F���{�`�z	)�ZžLT��z$u��Vw
.�ZùKS��p,~��Z	/�_ɱGQ��|!p��[{!{��E?��]��W�M�"��b,��M6��P��\�J�!��b,��M7��V��V�A�+��o!t��@�\r�zo@��t�?.B=�?��^y�rjF��|�;-@>�<��X~�toL��s�9/F>�<��QvsL�@��;�m�*7�:���qM�@��:�i�->�0���{F�K�� 1�e�/?�1���zG�J�=�H<�B��nq�UQ��	�0�O:�E��a~�XR��	�2�G3�M��dy�RY���:Ǝ����=A�~�UJT�Άw����7K�w�QKU�̅s����7H�x�_D_�φy�� W!�� �Nzֲ�:l���T&��$�Fq޻�=i���
[,��,�Awڸ�=i���Yc͘�j�����`>�ņc͙�g�����b1�ˋm�j��� ��c=�Ώl�,j��[�%����z�Dx�+`��V�/����r�Fy�+`��T�+��w�A~�,g5�C���\����ˎ7����E;�O���R����ɋ0����D9�K���R����ˉ6����A8�Nʊ����g��:�����ew2�����g��:����ft6�����b��9������bp:�����|�t2�����>��d�A�9�}�v1�����=��i�C�9�|�s5�����:��a�I�3�w�~xpN�Vt�/��u�<}��C�(zrL�Uw�+��p�9y��E�"pxF�_~�#���0w��D�/|sM���9`����� u��G�2��9`�����u�D�4��1h�����}��D�4��1h�F/>b��9!�a�{����N&4h��3+�n�v����A*=`��?'�c�{��� �C+=��^+��s�6��s�#������Z.��t�=��~�)������Z.��t�=��~�)� �����R&N2��L�t}9}��G+l�B�I8��B�|s2v��K&a�K�C0��A�}p0t��J+m�E�M?�┒5��mL^���wc(%|$֒�6��mL^���wc(%|%Ԗ�1��gFW���}h%(q/ܚ�1���=*�2��`ʳy�Elee�����5%�<�kϴ{�Dnfd�����<-�6��mɴ{�Eldg�����6'�﮴�&΍H}����<����ﯷ� ƄCv񯋺7����⢾�!ˋAv����4����﮴��'�?�kF�����\}�w��#�5�bL�
����\}�v��%�=�jD�����\}�v��%J�v@�x�AX{nKDC����XMG�{M�u�HU{cDHF����[NM�rB�x�B]|fAON����RFJ�v@���ꩰ#�q3O�u厖`�"���ꨲ �t5H�s���b�"���ꨲ �t5H�s≐e�(�����[�# j쥉�|�a9����P�(.dஃ�z�e?����W�,-fஃ�{�f;����Tsq�.�s�ޯ�����n�p�rq�.�s�ޯ�����n�p�uy�%�~�ե�����e�z�wu�d!D��R��Cs�	i1�7ˊ`$B��T��@q�i1�7ʈb'A��V��@q�i1�7ˊ`$B]2UYOc�P���K���0G|_0T\Ij�[���B�ʏ=MtT:]_Ka�T���N�Ł4B}_3Uָ7ݘ�k��e3mv�;'lgָ7ݙ�i��d3mv�;'lgָ7ݘ�k��e3mv�;'lgָ7��{�R��\�����z��6`�r�Y��[�����t��9n�}�R��^������p��>i�x�!)'3زxIj�9�swy��!)'3زxIj�9�swy��!)'3سz Mo�<�wt}��)!/;�A�˳Tl+�߁O�kd2~���N�˳Tc%�چJ�ie0}���F�û\d#�لK�ie0}���F�Ö��%�Uz�;��$��@�����%�Uz�:�� ��G����� �	R}�>��#��E�����$"/u�<1����-�j�S�0� *r�5;����(�i�Q�0� *r�5;����(�i�Q�0� *r�k��r�o^�����x��*r��c��t�k[�󛙛��(��h��s�n]�𖕕p��'s��n���&_y0�J&��u��W�Jo�b�$]{1�J&��u��W�Jo�b�$]{1�J&��u��W�Jo�b�&Y~-uHد.�_��9:3�`��f)~BѦ'�T��9<7�i��h'vKڢ#�R��9;2�c��e*}AҺ��_�a�՞Z4��	�����򺄘_�a�՞Z4��	�����򺄘_�b�ӖS>�������񻆚]�ޚ�;�G�K��+;�T {��Ӗ�4�N�F��*=�R!��ߛ�9�D�N��/8�V$~��ޚ�,�ݛ���^%&��ֹ�~�p,�ݛ���^'#�	�ݴ�s�z$�ؘ���^%&��Ҽ�y�w*�٘��Z�VOu��\J�(�D��Y�^Bx� �VC�/�A��^�_@z� �VC�/�C��]�dB�sZ\60P�{�h
��hE7kO�yR[33R�{�j	��fO=lJ�{R[05U�}�c��hC1hI�z�Z/zր/6&�d�f�6tr�P$vԃ.0!�f�f�6tr�R'rц+5$�d�f�6tr�W �ަQ� �+ZV���+l�ѪV�!�)^S���
� d�ަQ�!�$S]����+n�ԭ/k��wUc�����Xj�=���/k��vW`����_l��>���/k��tTe�����Pa��6���-k��GYy_d�_{Ȃ�g�F��@QpTi�Z}ɂ�c�D��BZy\a�UpÊ�k�I��OQZĐ΁���0>�`��-��Em�O��́���0<�e��'��H`�EȔɂ���0>�b��*��N`�B˙ŋe�w�+SQ:�K������,d�v�.VV2�@��ʋ��&g�t�$\Q7�B��ˉ��!o�~�h��[<�<��qm��.�#d��S:�?��qm�� #q�"d��W6�7��{d��.|�%g��u]��GN���<4���g)�fzT��GE���42���g)�gyR��MI���<4���g)�gxV�[m����l�ߨ�
���oGYb����h�ӧ����hCTo����n�Ӡ
� ���lD\e�����v�r^$���`�/>m�� �q�xU)���j�*=o�� �r�~R!���b�.>m�腘5�d�	��߮�v��jo����2�i���ߨ�v��lj���6�a���Ԣ���oj����9���9����_/�fIZTY���:����_.�bL\S^	���8����_/�bL]\P���1�E�u�pkP-�㸐�W�/�}@�y�tnW%�鲛�^� � C�p�fP �벛�\�%�w
H�.�K��Y!�&X[��93�&f+�O��X!�&X[��93�%d&�C��S*�-RS��?6�+i%	�F�	�4t�qY�J �:Hbn��4u�|Qw�L�;Hbo��<|�w]}�J �:Hbo��= � X�n�~5���

?>����J 6�L��CٽmK���c�ɫ=M� ���x:���f�J==����d� 4ꨅ2b
H+:�
dj�1��1'�'�����#�E��<SAr��V�\Mi��"?��dV�V����t��t��䜦LO`YK��,I���( @�=:M�}ℴi��uەIZزg��*]Bk�-HU<�R3>F�,�#����ɚt�'�2xئ�Q�,E��f��V��H6�U�Ǟ$����.vmN�bU���gsX����H!y�\�r�FԫW��pVG�R��,uhH�B���&�����@r\Z��))ў����ғ�p���jχ!;,%Z��W�X�<�Ԯ@�,��%���I5�)``KݟE�J�
��B^ ^��^�B�$V]�U=*�$�� ��ы3��dy�c�x^ֵ�m�<����@��uI��׶X0�xXt�#,Q�8t�v�hM۵c�DtA���B>	E�@q4�҇~B,�� w���p$ȔF�*u���'(��(�̞H�2ya3D�"a$�0�b��y���S�5�H"r��!��x&�_�J�6}��������
>8�u��ƅ1u��� ��zGr���>D�L#��<u�`h���&CWf��f�5iJ�WhGIDa4�֊#m��-���4H*}2���_M��2@�NDu*�C��p?�pg��xa��c�0>N�Q�dM;[]
ah���M?`�0c�U�#A̘�UEPwI�x��ހ0��T��iAs�D+1'ǚ��O�0#s��&w�E*���d�����aŬ� Q/݂^�a�� )H)pUv
O�٠�h�$#2Xs`�H��hQ���dūX�.EB�#�  ����P�!���<tY1�Ǻ{��iBt!�;nZB䉃j�X�����=��4C�
,���U�xPCA2r� �g}��UJz��g��X�n��f+�y�C�-e�I"T�b�r�(2�ӗ�M��,�JH����,U@.}�
�+3ڄ�(.����Ë����	�`%2�(�a�8/4֔���M@8�s�۩ok�h �H�4�!�$:�*�� �Xΐa$���z��O&���֏w%tM`�!ȋ��O�d{��޿�l�#&�
Z���'W��@���0/Z]iu�:{4�)�`���ے!�W�)��<1W*E�\�#��P�b��I�y�<a�Dмf��4x���MgDYӦu?A����d*�:LOE�$Eٛh�8Hv��ǠQ���'ƢY��FĦ�(Q�ū({�S��Cܖ�ZB(D��J��U���B�$Z�j�a�*3D�h���(O���qA�X�t�XS�.D�����?#�̑�w�4�D�5�.D�@a֌N4C>�V��Tz0NĪL��B�u,��&
�_�n�jq̒u��B䉘
��=(�D��=�Q�1n/l8�B䉨1�b%X�jۏ��a�@�E4�HB��43���Q��:n۲��P����C䉼a9|�*���0�ܹ+�o�l$�C�Ip/��q1b�/V����J4�B�	"�{U��>����-_�T��C�I+&�nm�E
��6h�G�����C�ɪM؈�tF�(25�rتK��C�5%�>��#̋<�\��O˄H�C�5&��hu�ŵ8��D@�8�\B�	%!��X���\� �цļ"�\B䉰D5��w������i�n�zB�I�-^���C��]��Ţ� BvU B�<]^�r���wȴ�p���8D�$B�ɱ�\ySd��h��q'�W7s�B䉳Q��4@���4zܓ#!�b����S1&�
c�ˈ��6�1�A&�	a*ĈHT8{r�){��,y�U�'��<[�(�%Y�.���S1�PAc�!�)X��>0���Ɋr� �l����S�O.&�zg�A�F��\��� :^����BR(wG�b�)��`�)�'8�<��r�y���C�J,���;'�'2R�=�◟H�g��6��� �u���Sy��`�%M��I+�O*�K����t��y�i}���j�'�*dqd�
���O��I.e�,m��G1�s���[�������{�(d�qC�J�����l���O(%����¡R8p<$�Ǎ&/A�$YK�ق�x�	���%`α�l�&A)��:��4*E>�SJ<�eV��𩃔B@�IY�2M�
���f}����]4f|�'d�ȭ�8Lm� F�HQb�a�~�K@���
R	o�;�RqQ!(��v M�q���� ������'��l�7wa�OQ?�r�c�0'��R���
	r00�O��Mk���ē��Ӫ��π ��36ʒ�8��.�}�����۾c�.͘�O@I�t�dᓱY�ra�.Z n��I�!)��Q���	�Q}�n�Φy��=��$���4�v��Ӆ�$	w�AT��v=��yVZ�L�S/ *�����3R:�~j�%@w��kg"!�L���ԟ�d�\<v'`���k��I��3pzd[��_�
����=��<�g0Eq~�	}}�O� �zrL��TN`��,�m��kQ)B/�y�$��h�e��|2����"��	P� �F���pҫ �\8(����@y��	/�py��Ss�A��ĩ�@�aq��yy������%�gZ>A�P
�������umȄZA(��$�(�F�^�ϓBH"U ���m�T�w=M��c��|k��&�i���[;Լ��FN8k�i9��L>���腣��U���ڄ	��lp��E+/�\<"��;��I���Oa���+"�$�֋�e�d`@�H��yBO��FޙB��	 b΀Zs���y�`�%�0:W��|�"���y���9�z8�C�M�����X��ygתT�6]
�ǖ�e|~q)�b��y2TC¨!#(XZz���IЇ�y��٘5�p� �SP!�%���R�y�Z�v��*qA\.E���8�y�CC�@ꂄ�f�P�9Nx�����y2�¼g�|X�*	EF��!5��6�yZ��s�]Jv��+���� �ȓ	Fy��'�
}��I�3KZ/7߂���X� �Pc��p������*e�^ �ȓz�A�����d����ѯ��/�؄ȓ��H	���O�*9���Y�.��ȓ]��C���eO�i�%.����ȓw�p##�?@�l���SUB���.L�)Çh�4o�E3cX6lӖ0��!9�!'̝W���A�2��ЄȓF���8���%
��3���ȓ~�����A2Y�-�� �K��܆ȓ�&�����Y?<���S���d��J�z$aH�.5�@�5��58�5��z$|�{f��K��\I����7}�Y�ȓ-�H�2G���\M��)$K&�ja�ȓ/��Ջ'���F�B���ņ/�4�ȓ����̶�x��+̪#~�$�ȓ-��u �˚�n�`��L"�!�ȓ8Qb�����5\k�S^�L�ȓu�Tq1`*L%>Y����O|����ȓ"t�((W�Bs�`����].z)��k�� �[� �(4˗/�G�(���蝺b�P**�2��O3~S�q�ȓ@�p`K�)TWl���Ы�-I3�X��*�X��`Q k|>1(�i�(w���ȓu�b]�a-[��	��Β9)p 0�ȓG��d��h!?%�"�R ���6���d�z���=9���B��X���]�9��@K��F��>���J�v�G���?e&-�+P�9��1�ȓ ��|�TF�=YD�}:��B�;xʠ��e��9 憱������{3h��ȓjV���"��]�ȴ������ȓh�8�N�.]��1P�I<R��)��Enfܛ���l&�vOǴ:��������
�1{���k3��1U����Z2�ҠG�'1�%�&0~4����xR�$
�v�ơR.�<(���fR*�!&��v`��@�G<ر��=� 8�]�%�2�s�h
 I���@F(���:kb�1���I^���p]N��e��-3�)����6=��ȓj1������kO�AgǡD�x��S�? n�C�Np��Q:�b�%?�d쓦"O���Ug[�!k���hB(g�T5�"O>��rE��vn�mK3	X����"OT� �J>m��Z��c}�m17"O����*AP�1��C&4iV!cS"O�p[�J�2��5gU�YoF4��"O�Y4��g��X��O�b���"O��
� ��3�qi�#P�M��� 7"O���U��o���ՍU�] �e�W"O��;��߃|@n��PmM(�xu� "O��#��K�%c�+V�`�"O�	��"4�,�����1p�����"OT�Q㋂>�X���H��<�F�ٰ"OJIj�͂aWpM��Q*΄2"O�}I���B2^�"d�!�8��"OX��T36�X�Hqg� �e"O���gĉn����Euj9 "O�u��m۶W{B!�b�/y�lj�"O�qq�	n�*5�d�	\p0�2"Of-��C��hv��֥��@V��3"O��2��-�M0BD�:h|�P"O���+˭x �q�Q$@�D�"O@] %b\�Z]V�		^�$^��P"Ot[���P�`u�ǅͺ`"py��"O.�)�(�)�yr$�%i>4�p"ONd*5k�'oQR����E�p�+�"O� �v&P.����Co�2,�D"OLQrr���F,ItN��Z��Lx�"O�E�A�N��`�����2�"O��K6��3J!�Թ#oօ;�T���"O�=���P�;�"��Į���1$"O�\ٰ���@I����킞wodq�U"O��;c��5����GLV�@^��"Oq�b暦��1!�N�5�p{�"O�L�������-pR���3"O��(�fB:qD><K7j]T,�X�"OFT0E�Y�u
�
�*(|H�"O��a �-�dQ��P)v0`l�W"O�#���,U���*#��=DFh��"O`�$�
b����ŋ��Rhv"O ����f, �լP��y��"O�]S�-D,P��"b��ƲX�G"O�ԂA��\Mɧ�a���%"O�\��F� B2R�����>���"Or5��̚c�l0!G^J�pc�"O,�s��b|[����4�N�q�"O@\aP��*�"�� ��"�:2�"O�U���J�h���j�3#�����"Or�s��14+`(��iýd�J%9F"O�Lʂh�:O���0��� R� ��'"O�(b�L�>�0�����S1�Ɂ"O��� �߱BȑI"��Ob}��"O\0��E�8c���7�^0aY�m �"O��a#G��1UH�R���k�x��"O��p�D؞\#��S����}<X�"OFhiBcG�N��A'�/mD�`�"O��R���]��e�&�#<=���"O���4��*d$��jDȞs#D,��"O�i��Ǒ�,��y*�:/ xٓ�"O�}�#AB1I`hj�刨���"O@ڃ/��<�f�АCտ6�` 2"O�e�fO�\����������	�"OH�A4KV�0���դG�B���"O$`����6(�a�[ި$w"O� �MB��(E"�%k���&ev�Z�"Oe�q��%]�5
�c��KW�\�"O��r�D
�mlIh���H!�""O PI��bX��1�ܒ<���R"O��!�!�'��7φ$����%"O0IR��pX|�eՃ [Xl[�"O�,Cׁ�{� �ó#�%EbD4��"OTI"a��F���x��ɜDS"O��X�H��A��D�`��qNF�C�"O�qh�s���zRkʹF���)b"O��8�)(��yE
�*gԄ���"O�ݸ�Ȓ�9���k�h),T,ڶ"O�p&��'_Lf}S��R�O^�"O�A��B�>~���p��W���d"OZ��L[1����Jp��Ȳ,Bz�<���� G�����.H<����R��~�<qSb�8�<����|�pHwhY~�<�K�.�����Z+j읰!dI}�<��˧~?:�KCL(����� u�<�T� G�T��S+O�,?,:��r�<�I��+հ�*K_'.'�ؙ�BJk�<т!Ív[Nځ(c!7F�*��\��#��z$k̴p���Ǡ��l��������H0�ڨ"�@�}�ny��UՂt��� ���#,Iq����ȓw���{S��1��	s�1h����L����EK�bI{�O�T���ȓo�����	�F�����F߮��x��e�H\���UZqRcM�V9$���7z������`Dτ��I�ȓ-��p)�-�8T�I� X�q��M��53��˧��@�����f�]��ȓ 6�ɛW�ĩƊ��!����}�ȓ901 BОR��!�#��y��j�Pt���O2>l�1Mo����uEZ!�F	G:-RY�m���� �(� *O�*��eI�f�^B2̅�|�� ��)ӔAm��䟅TN��ȓ[�*I��s�8����7)Έ��P{�A���2qV�k�@����x��"���E�
f�8��.#qV���ȓ%������[��
f���p�p�ȓ�ЕR�ߞq|Ґ�#��=k���D:Ho��I��ʏ_\��ȓrΦLX��5t�Dʱ�E�En�Ȇ�L>�����_���t�j?P��ȓe�ܘ�p���px���̛�U����v����R��&c扫�(ρi� ���42��E�D����G�2���@���1R1��3���b ���ȓ$:�Eّz��rգZ9dژT�ȓJ?ZP��$��@�b���û�D=��W �fj#����CAϳl����ȓ���1ɝ&zv~8ٰ�L�"�D�ȓS�̍3�ŗ|'Nq`��,Q���ȓzF�ⱪ ��<���#Y�x.t��ȓrY�Dz��w�0Mp6hʼh6q��;��yl̖3��qY􅟾%ւP�ȓc"�Ṙ:z����%�}�؇�(.}�!*T(;9.LafB,?��K@�u�v�R%��m;���{��B��1+&'ȷ�t+Ge� �t��o�b4�E��B�F!�F.C=kr�ՆȓOL�W%�-��i���κ�H��S�? >e�7��NL��@-u�Ġ �"O�\��VP����j�z��"O����a˔@��Ķo�>h��"O"�c�.c5l��@��d�#�"O�$��@�x��j����-��"O��Õ�ž ^�H�a�At�"OB��p쇽*�N!X!bP%(�hw"O(�`vL��]��p�3��M�iP"O�,z� �Z<�h�FD�;c9��ӗ"Oָ+�c�
c���Q�R�JRbT"O��Sg䜠L@:�Jᇒ3k
qH�"O��I���6�a�(X0t��"O�����#A2��+5����"O��w-�dF���/����E83"O�t��@¡�`���퓌;���0S"O��S$B�`�4�:�-D f����"OX�IC   �(   c  W  �  "  G(  �.  5  S;  s<   Ĵ���	����Zv)���P��@_zX�B�W4S���y��ƕ	#�e�H<!����іS�E�aYҋ�k�<�%�
I��Br""�.ٺ�C$Z�h�����,5���m��e��
��Y�@<j�Y2�~y�
F*F�y���J!G�}[�璛ynơK!F5�V��1�Ҭ��9���~\�q�Gv.*όl3�X�%��a�4��.���0p.(�j�.�4�Q���>�x����$u���(3�'���'�BS>I���cr���+M���f��fn��C�rZ��	��j6�E[Zw��Pf���3M<)Т�+ vkUF��f!B�ö댯0dİ3gY�Tr���f@�E�0�O��Y0��7�$�0'����C���CpY�RΛ��'/�|h`�'�l���|�'�l�]���p��Y&&gv�@���Q��Ȁ��F��M��'W����͞�0�V!��hJ	r�Z��4?�&j�,�����=�I�?-�S_�$n tj�,q��D�bw#�Ta|�p$^�a�"�'�'�����	�|r����%ܙ3���T���&߷3T��#Cѧ$>p� K%C���e�]ȣ<y"�=P0@u�ģ,�d�	(w0����^� ���Jҥ]��X[䥄�{�2�<�g*����q��U;�I��LB�iX\j����M���@�'�4�	 L��İ�*Ųj����'��1Cť�� �Ș �ϭg~�QQ�OZPo�̟��'2J��7��~b�����:I�!AuHڭ���Ƿ�M㖊��?	���?y���Z��j�E�
�H4�퀒\���C썚Y֦,�4i�$�P�R~	*� ʓzo�h��cݿz3�q���`���̱_��)�Cm�-<�b�qFB{��(B�1�!����;�M[��)6|^b��BZ�4_ZBC�8��Q��\ҕ͍?_�X��lJ�/�d�(�$�O`4�'��(b`I
�F����C]'YKb8ٯO��[���q�	ȟ8�Od�x9��'��Ak���&yQ�-R��S�!��7��h�V\�"퇪U�̫1��	����F�+��b>}�c��T�){���]��"��	����bV�`n��ڤn�:D�8$�0H�)5\��iǖB� �0��X�Dcl�Kp)Ĕ/����sZ��vӞ����'��	 �K����F�x����V���8&"OV}���3cg���������Ð��9�ȟ��ʷF� ^͖��D���4I�����)��ß��#�9L���	����I��iXw�O�+`��[���?h�:�*ł�E�@	W(�*oyr�+VlìuC�hF��|��T,9�
ObQU�W)����CR$n��l�ժ�x���!��7&}���K�f��ӪI��x��xRdZ�zJ՚qnR�>�@���fV$���IDbӴ�Fz��ODY���JV"0�2�Jw�L�y�"O��.V�62����Ȕ������"��|b����$N?X`���	�L�d�h'�O�Z�!Aj�GѼ�$�O��d�O�L���?I�����@5��!��>|���* 슀m��\jP%
-���jkӧ+�z�i�Ʌ�<<�Ey�&���Vpg���i>�æ���6!�t��@th!1%E�9E�iAB�^:qNaEy���?���`N��P�X�S|�I�% -���G,���Ov�Cgŏ9��sm��$|;e"O^<(�/K��a�ꄚT���A�V���۴�?�/O!��f�O�4�'J������k1��7Y� ��@oՉ �*M�x<"�'vE����&�܅L���F"R0)'.�R� �`7���1�
�Q��W�£^�p�x���m^|=��c�r��qv$N9dҺ$q6W�O*�a%��*ڒ�Ĭڴ��$+�M������MÒ�)ۓv������xA�D)O_$�FS���I�[���z��Y���d
�;�����k~"�;w���b���Ef�q	am�&������O��d�|�����?��!v>l#�B�U��#RTs�8Z�i��� �Өm*�1�NWY�q%�	��0��T�iŴf�)Jf*P�Y����¬>���Q�^���4�� >j�|�*L.\�r�C%���O�0�b����TƏ�*����'���fg��@�<%?�O�
�t@�d
qk�+MZp��c"O�iR�`פ{ט�����:_Ό+���ȟ9Ѐ��42P�_�b�k�L���1���0��S�pL�OL��|>�$D��[VXUyG�O���4�Ї�4%��|:vX�^�( ���{jq*�JK6Y;�= ��H�&�x�*�#T�H�ZC>U��AC<6�����[>���!$��|9�(�2|
��J��ēG�&X��J�,YRT!�NݓNI~	�'y�dA�YM�F0ғ�~��4qR0��L(o�Y�*���y��>�"$J���~)<�Xa)���M#��i>!��Yy�B��N�q��Q�|�H#'ȉo�2p+�H�102�'Pb�'���Ο$�	�|�2+��(J�}Ւ0��#���uQ�\��4"Ƣ�`
�Ӷ.�Ȱgp�(�J;�O�	(��'�]*���pðD	����6��G�8D����ݶ0n��+A.ƆtN�]Bu�6D���7.O�Ra�GB=M���Tb�>�g�i�'��`P��z���D�O��ӭ?������/.?��U)W.7m ������O���4lw��d.�?eX��� w��=���ރ$�2Y�4�2ړivNmD�� (�9��:sr�E�GL_�#�Ę�3�	9B��MX�O@80�dO�7E�4pH�l�C-,(�'}^��&�0�sU��8=/4a������o�+������9��nΖ	�d�M�h!�$�i�"�'��-�:��	�@K�.�L�y��Û10<m��M���P8�?q�y*��O�(���<~�����.�9�]�M˔�f�����Z��E�5�(u�E(L�D�Sу�ORX��'�O?� c醞p��C�B�.����\O�<��hA��ecM�TY�U�P�SC�'b�#R K��qJr�B�]،��ˏ�E��'2E�)y����'���'C2�O�Zc�xر��2ủ9�>�2�/ODhPd�'DkY!(�r��j��'�n�Z,O.���'H�,��*�8CƄ�s���<�(,O	��'����dW 3nZ���Y��l�qT�ɲe!���gW�`V �[�h�	�D�W�5��|jN>�t! hV�ʴu�ѫJ6a��0����?����?��a;�N�O��$l>�� ��O��b���:���ZPF��ј���Ix���c"��t�p��'8��(�sK���j�@"�"�Od�@B�'L��4@\)f�,�� ��+(��Y#�?D�ї!��3V����ĀN'<H�eE=D��� �^8��G^/�$@)��>��i�'p�Da�.z�����O��Ӈ�����#a��㟷 ��7��!.�f�d�O��Ē,8U��D&�?yKb	;���˳.��J!�p���(ړ �J�G�D`I<8B�,(����b��8Ⴏ���hO�Xr�'�,"|*��$���֥W/``I��r�<�A����|��G�/u3X� iX�L!�O�@�E$��w�Ya�%E�6DP�r�Y�p��芄�M;���?�/�`|����O��m:�e���k���:�o�@r1nZ5/y L��x�S��}�$�&Mg�\���O��YK�(��?醠�l����4]� X�1Z�4+S��&�` ,�O�%��';�O?cU��I�Qs�͆f�N�+�i�<!��C��l�a��ŀT �qv'Mb�'��"�Ъ�/q���yr�ƫ*�4���e�5����'pr���б)S�'���'���kݥ�i��Sf�Μ5P��d�Ζ芄 �h~Ӯ�$��n��h@��� ����cnx%Ղ�]�� �3�P�8�`iy@Z�b_��x�
O����l�|r���f�O
|���%8{�<��a�t�����iAb'��z������O��	'R~~�+�*��vEd���Y�q�#=�Ǔr<X#�̀3x�LQ���7��MmZ��M���i��'�1@v�O+�ɟ[V ��h�Y�A��U�-B`�V*W�����֟@��柔Zw�r�'1��� l	�x�@�
�:n��0'%yF�����<B|��2"2�p=��D��r���K�L�x�!�Q�I5��l�e[����/۸>S���%�&e���<I֪��T'oH5D�v쳧ݴ+��u��Ν�MCՔx2�'-"�T?��e�ܔB���jք��C-@I`�/�d/�O���W��#K��K��6.��4�P�T��40��Q��Kaa̰����Oh��O�%Ze�NV�"�56m�r���d�O��ă�<�HAd��$��عRG¿RF���'�ލ��EC�_^ bf�F�y�z�G{"��)@O���3� �D)�/P(n��T�C@�0cwF�|���1��'�ў`;���OH��:�-
�xi�L�����
���?Y
�X�D���ꘘr����te��:ZQ��	����-��D�QOI�[��{�ꋤq��I�%�V���4�?9����i>L����O���R/Ga�q���8OL�� ���r�n 9�E1�cCop��&�J����'�S�|��p��l�$b����� �) >x�ɳ+��a(!�D�9��,��I�E�p�G��)���y���'����O #��H��?9�������'A���-J:sT.$�
�#�U�)�!�_(jւ��X/Y_`�pƌ��/*���������z��q��I�[�=ӁƨM?z�l��0��*�(�bO̟��	ʟ��-�u��'���!a�?Y��lK�
�<��
��J�002F�
�}�r�	0eЦ:"B�'�O�)�땤a�Y��J+kx)˥	A�:Ժ����[}r4jҰ�Yk/��#<I��P_��س쟅=Z��fZby��2�?���?��џZpC�
D\�؀��Vw�ɰr"O���a�����)��_�W�%x1�i�#=ͧ�?�,O�8�uh�9�A�5
A�yʲ�+��W�K#�T*C�Ov���O^�dNݺ#��?�O&�EᐁLE6<�!�&T9�� �����aH0S��������џl��i ��p.me��
'��L1PR'ω��]�U�·9`�E� I�?qp� ��q�lW�U�Z�Z#Lڎ'v��C�i��� ���b�N":d #`��,[�*]Z��?D�p:4jX7�,q����p{� ��,�>q��iV���I��\faa�'���!J��x�R���/�06c�0�bE�6��x�"Oh�Y�'׆96v��rD�T��E�"O6P���b�$:wj҆_����S"Ob��b�M)'�>���ߍ_�8��R"O`�H��z��
D/Z�;``b�"O]AU��Y���G�^�vx��"OQ�sH	�rV�c5iO?|0��"O���6���p��WO��"+)h"O��P�E0.)��r�B�H}�e"OZ�Z��Ͼ-�^��J܁;��h��"Oh�4*d��D��)ۯq���JQ"O�� �i̳oT�Pb�m΢X$i��"O~yQ���f�
�l��`$��	"O �i�K�(�N�8��JV1("O��⧫���zV�J�8*�ы�"O��R�ʉ@U�ᳵ'��n��s�"O����	�@Q��Y<t�ȹ�"O8xXя� q�IbaE�F@F9��"O�\��b���΅ڇ��6����"Op �rB��1��E��)J�m���;3"O�8��l@
s�(ي����' �(�"O0y ���g��A /X@&b�"O��n�	�Fi��@,�|�!�"O�� A�V��1�\T�^�"O���e��GYv-�D�3f?���"O�,h�'N
4LXc�C>]R��s�"O0��ś2�z%�6�^�c�6p��"O6�q�˴8h�c�5�!�"O(�� m��m�P�\�6�� �"O:��cL�5p��aZ�7H�r��"O�)c%�(1�%;� f�:�r�"O(�5i�
vE8�M�И��f"O2�cviD0N���BMS��|L�g"Oܠ3S��z6���,58���"O:��#H�op ���I�B!6��A"O�Dh�*0ƙ谉�.' �4"O�a�0+Mo>�m��=We�|�T"O�ܒN�9?���3
߭&Z:��q"O��Сν&�<2�:=A�0kF"OʤP5IۊЦ�SAN?(�XHH "Oܘ�l�)p$Q`�*l��͓�"Ox=p�@<4^Ya�g�8/��"O(U:��׭�m��fS>_e�&"O"H�B�[�	����Ao�=gl��91*O"T�3eN?Pe����5irQ;�'���`����}Դ=c�)'��$�'�m�P�OGb��9r�מ"��@�'F4CD1^[l�
C�ؑTs����'^����6:q^�2��#!��
�'�lYD�ղE��=�r�����	�'���S�V�Nri�֟6� ��	�'��sm��)|:H p֭(���	�'l���-�&AnƩ:t�'[�t�0�'�lA"$�@�<�0�J�#A�، �'&n!�a��<8锹ʦ���eh	�'���{�M;^f��!�1
�$B	�'r4����){���c�o�8 ���(�'H����,Ӏ(�d�b�|�'��ى�*Y�b^���Fm�;���	�'^�2���4k�bU��D)X �"�'��(�P�C4�p�QEVH�"��	��� zQ�RN6 h�������t$"O���(Q�!�J�R�νS��=��"O�I��C?~�]���^6vv�۶"O��b���a4(L�CNȕ�`"O�;�^54�8eK#�'�X�"O�iؠJ�䅑&^`F���{N!��
�Ph���uƕX|:�qa�6 �!��Qk�$����[�����Ed!�D]�T�td�3�T��÷iG$NR!�9#�Lj�JN����6��0D��ǿ@���1�lI�A$�	ۄ���y�!��Nk�[�Oyl� �����yb�.\��4�`Q"�,�y���+�@�6M�`p��͔<�ya�:hz����D$�t����y�&�<x8|0��7"'d�����yRcۦo57
!��yR򡌀!�!��5L������W�����H�!�$�2 ϶\���k�DQ#��
�!�d(����-��Q�gW�<�!���(`^����jE�A�4�j>!��Z5�H�0Td��2�R�b�EX7F!��U�uS�N�u�*��ܖy�!�C��԰ V�^=�K�5n�!��3e���B�*
"��Ԋ�/�!�D�������8v1�Q�h�!򄊔��Y�"�/\z�|p��
�d�!���L�
S��1h�t�W��/1!�D��'h.d���'�N���B� �!��ҡM%R�`S�ϣ]�$����	�!�H/Ƞ���#Z̺1�ǋ�9-s!�>BpH��V	'!/���Ŋ;�!�d�*|��� �I d�d	�F�[Y!�DG?M�8����!l�X#���7W!��y5nP��m�pC�yȇ��4K!�d��Aɜu�I]�:�;���!�ϲ`�Ӥ_�t�ꨉ1�	�.�!�dE-cx��vaˠ�$)3�+@��!�$
(C�\H��;��i v�\�B)!��	)��]��j˘-v2�Q5��$}!����18c�.-7�ɸ�mM(X!��B�Ve�ʶH[�z>�!���eS!�ht+%c�zy�G��H�!�?zP��B�J�#4�E�c�gC!���+R�ٴbE�# &�c�$8�!�D߆�`} G�7x�y�˝>/�!�أi�� ��)��K��V	!����	נ�?�V �)ɩ)�!�_�s.����I����r�Fm�!��(HH���&�j�e�İO?!�$��zϚu*c�Ы0�@��D
�s�!���9]_.i�S&�-xL����f��F1!�DY+��䒑mE�>��x��F��Lr!�Ď.E��`J��ʋx�j�2��˨;!�R?��Q��d���20c��Ukn!��� w"d�Q��@FY
����	�!�$B�ףׁ��mBcm�_�!�䀨�
VC��5���P�H �!��;X�&�`#)\�o�x%�,[Z�!�Dٺ|$`�E��2��"@�#-!��H�v=ȱ
0=fd9�a	�!�đ@��9;"ڜF_�t���":!�O�$2���%�O�d����x!�dǟi�Xۤ�2O���IAi!�� r�P'�ܔU������/;Y��
�"O*؂� ^-c>�u@g
֏}P�q �"Oi�A��� m8�O*
��Yx�"O&5:6�ܙB�b���'ݐU�81�w"Op�X��Zb�KqV#��a�"O�͸�"��|���f�=3�xX"Od ���	 �Y�b�
}R"O�-s��m��T�R�Q�d6ָS6"O�0�P���T��5�um����	`"O�%�Wh�K��x$��*[0��	"O|�0���A�<�ń�5Z�H "O�C�8>زő�*
vw���"Op�E� T}�\1r�!3��"�"OF�x�h�L��`�ï�:.��i�"O-a�':����MA�_3�ŠB"O��*Ǭ\�n���q�a�N]�b"Ob	�c��r�����D�ĸc�"O� )#�?i��P!����Jq"O�e���=���C��P�rD1�"Op�*'��WCX=����8�Ru��"O��"�Gɷ�2U��eS#
4�P� "Ox!�P�Մ ���FD dD��"O�إ��i)(H�UE����}�B"OZ����Δ8�����$N��lSA"O�H�`���S��hK#虓5HT"�"Ox��K� 1ԸrF1�`<�"OB��s�Л �(����2I�x��u"OR�X���d4((�dN0'?�i��"O�-ұ�ʙ(]$qA�)�<o-�h�"OLQɦ!�&h��t��߃s�I9@"O�x�V�i�Y��խڞ4Ye"OIe�Q���4�Be�)>ʢ ��"Oze��!�3dY���"Q=�1b6"O����B�;}S�liRb��82$�"O��5@�=�|��c�M!�)1�'�`�d)$ �
@�e��_N����'0j1�5J��$�RQ1����'
(p��M1Y�K�J[�C떡��'�,�� &ܭ!��Y�rn]COP��
�'�N��b ��
��fϏ~��Q
�'v�KSP�Ta��	�-&��	�'��5��EL�HA`e��dŭh����'��x�W%���6�8��*�:e#�'s�95�����WC$[�����'ȕ ��4(.N���h�WFE
	�';X���Ȝ� u�ͫ<C�Q�'�N���9�͐RD  ~UH�[�'����g^�!�ß�^���S�'hX�Pg�G��X��8 Z~���'��ia�n�1��2`H�?�b���'EL,j�a�j������F>2D�X�'�
Ha��P�Q��S�$/hXe�
�'L"9�ae�S��Qe��^zт
�'�|% qo�D���i�Y\��Q
�'n��B皝:�d%��h�V��h	
�'~��*�S�9�0�ǍME�M�'���R�¡=��hb�J�B��|�	�'-p���"B!`c͋���.��m��'Z"��R�׳���r�H&,2*Q�	�'�x����N�38@�z"#�7n�*A	�'�����
, �uAA &��r�'��Q��4���A�0:���'A�������0 Kq�ՀzZU�ȓ|�[R�G?��I��ņ�}Dm��S�? p=
s	� ��%���4&��:$"Ob�U'B�����QgH<S�"O��T�J�`�Ȉ��=c�xQ�"O�=�O�s+��K��E�d��"O6�����V��D��jً�
��"O0X*�΄"_�<<�1����`Q"OH��4�Y:����M�r�	�i�R�q��&( h#�΀3dv6�'C$y��C/1E�i���*TS!򄌦	���۠J��&��Dn�3P!��Wc�։2�QM�|@;�JQ�tM!����:u(���t�|�ɵ`_�Z�!�d�nq~�uk��Hf�[�ϑ4?!�d�n��@#B3?7r��d�V�90!�(xl��m۠04���E� ++!�@},�:�P.$��I�ȋ��!򤒗kP����!1���	ͩ-�!�Z�P�2�ʊ1���
*r�!�dV�
�~��4��؅C��h!�$?�Ҕ�%�ؙ"݌��ȗ%�!�D׉w�LX
7ᇕ e�U��hޓUv!��7f&���6(��[d�J�E�@!�!��B�q<~9��mH�W�!�d+c�v�3f �*���!�()�!�$R*io8�hf�٨|�����ו�!�i���BLP&e����Ga�!�Ă}��kd��u�湃��Ҩ\�!�䛌[�Bm�ဟ�']�|"	#D�!��J4>���
lܻ
[vء���/M�!�$N�B\�H�eɤ QP�� �>j�!�$qA���ʅ�j3�)�	#Sl!�dVw��6��5{)l�bHіBy!���{/XىD��9B�X��W�F�!�]6�[@��*t�Pã�_)h�!��S
|��	��p����%��L��򄇌<nu�#�)i����0�yb(�F|��&��/�p5P�A���y2�Ɍaz-3��%tB�a�jc!�d�]� m�S(½)&ǉ�b�!��Z�:a&-0���		NC!��̢���#M<HB���%-Y!�M3�8�8�Ʌ X5���4��AQ!�ď'}�*QS�!R�ʢ̺�B��;�!� U�z]�ʖ�6� �B�E0�!�DEpҘ%��BGLJ�3��D!�DғI�0�Q5t\�tk���d(!�[<T�ڍs3�2rH�<�'�M�D!�dO3�6��SMI�aJR����"�!�d�D�n���F��F������1L�!��:4�k�̄2Tۘu��ϔ��!�$-"y�5�I�{s�Y�(o�!���w+N\27�-v�jT[�-���!��?E������_��z�R�+ڳ-�!�Ę�7=6��CȜm�`ۥ�� ?�!�9 ��u����P�6YK"K� �!�֞,h�����9`�����
&A�!�d�4�����\y4dȕ,�!�D�^�7%%S���c�Oh!�d_�$��I�Jd��!��%$d!��z���0��=��A�wf�l!��z��=�g�Z��m��><!��q�JԱQ�5_�^�	wEU&-!�г@���p��&� X�GCA�k�!��M�(��{���hvH�:A�r!��B�pr\A��7���!�/<T!�� ~�p�o"���+2�P�p$tmB"O�|�"g�+m%�1.>Ω:�"Of�ɔ�^�&��C��1�FT��"O�M1��6Ḩ�bc�7f�2M�A"OjA 䔱��tR��ʹx;"Onpr�׌	6�����.�(�Kt"O<�$�1(Z J�i�U��Uۃ"OĹ�Ġ�'gN���)ݚUҌc"Ol�Sd��>`�8tqHX�\ ��V"OЙ�M�{�a��!�"�Q0"O�ep�Ut�b
=>���(�"O��[��֐pq�P��
_�j��B"O5�@���	b����Y��"O^pD�Lr6��p	:Kղ4�"O��%��h<↏V4d.<��"O!�������G����"O8i0�L>�
I�ѨW�6�U"O������H�^1y�F��qpu�q"Oflr'����4�SM�MV�]�A"O��c#� ��!!�N��EG���*O6���(�`�v�r��J:
���
�'?�� b�Ä2|~ɶ��/Kw�a�'?�5J���M�t��Xw/����'Z>�$c[�U�{P�[�iw�}I�'{�����K�-<=2Pe�8��*�'!|3��L�b����Vb���'���h�g��&fBD�ä�8F$�q�'�l���U��A#/��*?j58�'?"e��L�-�̝�%lֹ4� Xi�'?�	�w͍ |��!�O�}�	�'Q��1u�U�W�� b%R/"ά��	�'w4l3 ��"ldj���>ݣ	�'n�T����-	i(uy�oŭp����'��C�0V~l��k !4��'� ӭ��Pxq12J
:E��R
�'Nay�C	LE��Qτ��`A	�'�t�+W�:l0p1V@jP�#�'�h�(��C�>3|��_+ ^��8�'ĥa���/_��å`;A�a�'(��q���"w�0���� ���'�"�jp�ԳN[Bq*.I{��P�'`��z�
��~9���;q��H��'�di9m@���d��Lo�\01�'�(�C����za�m���;] �Mh�'' �+A�߭D��H[�'
N�U�
�'��m�0ͪxej���o��qԌ2�'o��{��(`;��*�E�0yf\aK
�'����.Q�"� !�t��9rO��	�'ql���a $��ؠ�MP)e5ԌA	�'�Z�MX[f��ů�`��)��'�L bu$#{i*���;\��A�'�JЪ"�%c�uD�U,IDd��'p������ IH�!Ԑla����'I��k��_�`��&��leh
���'J,���'��{o�0Vc���L��'t�4;�@LU��ke'E�t�x�
�}�/t��ħ(~�lX�U�]���+�c�;k�z̈́�'����<O��#��!�$����D��(��ɩ&kn��qm����� �T�;�FB�If�M�2��m��-���O-�5�������%N��S��b-p)��ΏK�6��d֗d˼٪E�>I�!��9��Yc�,+:>�� ���<)ӄZ ����&��Sl�94L�'�p��� $�Gb8�@)�4��(��
k9t)��S�? ѹ���Z�Xh�3"�0T�V�h�"OpA+��Ŭ-44؃a�&n �"O��5D* X�!a���٘�"O�<h����f��l��$�"O���Ȃ1ju�`E�~oPTb�"OЈ�bP�i�4���ҹ1�Θ1$"O�m���bfx�*��F�1���E"O*Y1EZ�.E��8U�U0u�4�T"O���1q�0���F�ADH���"O���ʖ7����G��?��0"O��{�L]��ً�!�1( L�8�"O����ޏ9�R)��62ց��"O\-�Uh�x|Y���6�h�f"Oɢqi�ft�a饋�P�lP�U"OvL���2	vMڷ�M��za"O�iz6�؟/L�UR�)�<
�D|(�"O����)��%adΔk���s�"O(�ɴ,�6"��P���Ҁ8�"O��(��/ޒ�"``�B���"O�����Y s1��-�� ��M�#"O�< �ݘE?�4���#�h(d"O�I{�8�Zx�#MM#y���s�"O��{&F��ƑHL�i�m�a"O]y�&'2������R>Ru�W"O��AJ�[T��䋋 7P��"O����Hƒ
]�c�N�u�:@"Op5��$��"�����Ȃ�
�Z�"O~9��΁e#�z'��<(,�3"O"}��Q�o���� �Z�<��"O���@��qPRt�R	ֈl"r(p"O�i�uhV�8��0�B�܀Y𠒳"O,�1흟0�K'GK'�*�1"O�,*��2s� �#��c�� �"O��R&ʊ�Zy��C�~�<#�"Oh@���.c�l�C�S5(�!"Oxbī��H�P ��K
�<5x�"O8���i�a'8QW$^*s�ڑ�%"O�s�L �M*��/~�yR�"OڰZ���r���`M�^zZ���"O�DP�e� IՖ)AT�1pE|AQ�"O���e�р4�h�4NS�r�0,(�"O���U�΀a8(��Fz��pq"ODlHS֤��Y5�]i�N�J�"Oh)spj��s�v,Pu$S.�r�B"OVa8"���*X���ȨL��۳"ON�A�����*�H�E��b��`�"O�e"5���~�P�#�O������"O&p:b�ѨY������T��`"Ox��EB�jH��2k�M~�k"O�p��O3A�
aE���Y]��"O�� 'ƙ��RY@a�ǅ>X��"O@p2��D9<��bO�*$�U��"OPd�S��*h��(��*wp\;"OZ��i�O�<��홱j��%p"O0��ƊF4"�z�I�BT%?�q� "O8�T@�$N��ݫ� ��	���"O�Xb�a�X�\5��)F��s'"O��� T9��$��o���"O~����
�H�
C�4OҪP�f"O
��DD�?{z�]��^P1�](�"O@�p�i�q�g_*01�"O��P�M+��4&K�E?\��r"OF9#0�
�Ȣ)GE�-G�b��"O8 J#��f޸"e#,��@�"O� ��@�$àd��ᏽLqR��p"O�0"G�҇Y|<��A�_�J^$��"OH���j�B���񤄳� ��"OHq@�ȇ�$�pA��ż]���"O����Ew�֙C��� %�0���"O���'��Az���g�pK��hF"O��p�.E�DM��,=8T�"ODّ���[W�m#4�]�#<<�BB"O�!��(�'�t$K@DY�bZ�]"OD��ef�/P�0Hx���"q<���c"Olx���/Q��(��CW0��ųw"O��	��
  ��   
  �  5  �  o+  ,7  �B  _N  dY  �c  �l  �u   }  	�  �  R�  �  h�  ��  �  2�  v�  ��  �  Y�  ��  ��  Q�  ��  ��  �  �  � � 2 2) �2 u= uM �W x_ �e �k �n  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H����<�۴#��M  N�2��e�wH� Cs�e��2 mj`Ni������	�<��ȓLu�8�5��%*���D����l����f�$'�VDc����8�ȓ��E$����"'����5p�d@�aY�V�*��g�Pt�ȓ=U҄h��p7��u�ޅ=��$�m#ᡃ�J�^�*d�+�"OD0Jć�;U��*R�V_��S�'ў�"�9:��au��qM�̋t�<D�h ��Z� &����#G���ǹ<���2�S�Oq,(��Ֆ @QJC��38Y�'�`��N��e�~��S�·0ra(O>�*lO�����@+����J<�J��"Ob������ D���X��>���"OL�`c�	 ?���6�'�B�Hq"OX�Z���e��� @�8���"O��@�eJ�FH] ��W��ơ�U"O�����F�v ��Kͭ?�
�j�"OV�&��P��Xb5$$D�"O�u�S��,\#�	Ѥh1�|+g"Ota��Ğ�E"!3"�֥"u��a�"O�q�	��0�R����J rGn�A@"O�I1�G�S������?H��,� "O� I%+*%��L�� ��qrP"O� ��jC�,LZ+�O�Y�(��f"O1�a'H����1a폰8�f�f"O\��Q�)V�i��ez��"O|��@U��AHt��L$l��"O�|r�	e�l��N�s�R�"O6��r�q�Ɂ�I�#�P�iB�N�<Y�!��~��V��q�l��[�TB䉅u��˕��,�ƽ2϶��B�	������ɸ�8!LN)n��O�q �'��)��Ej��(c!�.5l����?�ݴ*�uRtK?�ԋ�aV�m|P���|�ɰ-�$�B�Շ~��ex�I�/>B�I��N���U���c��:��B�	^$�-�1�v�hqJ��L3RV�O"�=�}�+D�eR�](Z3z<Q�lSI�<���ϩ/b���آo��p ���Dܓ��=y׋�r@���B�U��N���d(<��H
�@ؘ0aa�ѥm��� ��(@�<���8��O 4��I�(L1%�Y2F�29.��4��4�(�<��scI3{�<12�LX�".$�#���Q������%����F��52��)��A��p!�ڽG� p��*�Lȳf!�?��c���3�g?9s��w�� 1R1m�9ps%�e�<Y5mE,*�:�B��D�8�v$�1���H���'�O`M�P���!{<�
�Ò�0e�	|ӎ�AK�8F{>ia��"~����VM������Y8��&��#􀟂`�{a*͉���w�8�b� �F���E "Za��`I�,������W%�y��7:���p/
23�\,C�*��Mی��s�X� T���	�,���E�3ɰ�K�"O�ܱťT�zGq�0�;d�!�9O���:	�$aR���'0�-h�ϘT�!��\��Xi d .DА��%!� Yu�E,�u˴9ِ��x!�I�.v���2ۚp�\���^�!�D
�>�S��ݒ*N�4Y���ZƉ'�X��D�?)����Q�{���5��;�!�Z�o���ҘV�X���ο_G!�$�x��	ؕK��� ��V�M�!�d�b���2QD �P�Z���A=z�!�$Ģ7=*H �Y�������5t!�D�_^hP�A�1+q�p �C�CoayB�	�
>A���/.��Kq G^���͂*�~<bfI)��#߬
6�H����?}&bU�;� ĨU�4�Vt�b&D���Z�A��QY��@!WX����%��<A㇞<N���v�G�V!�i[��R}�<!2cS��) @�:w�:Ű�&�d�<9���EK���GIW�09H�P��	c�<a#�ׇ	�,!9q�I�܂D��Zj�<�TEϜu��A �D���k�j�<�lۜWS(��GF�J�ҵ[��	c�<���"5x4��G��6 -��&��y�<�FK�) M��z��=��@+��w�<�5�:G.)�ǁQ�`��Yd��	E����/��ʓ{��#?��ؖ�ʰ+�&��B���}��x�'�<��=D���[-Vp8��P�$����K؟(��$�P�xu. &X  �b<��6�Q����ғͤe�^L�"��,���w"O<ݹ�h��&�)Is�H6x���&ў"~ΓkV ��EǏ�Mt�`��GM�BT��N\P]��5���E��<r�x��	]<9�FC��1Q�̆9����APB�<�3G]��z�$��9��5LD�<� 2��K�z��S�n����LX�"O����Ց�U�n��� �"O2� K�
$0�p�?vi�00�"OPaʠ�Ы�:dZ"��r��E#%"O�j���5R��و��A�F
�%�`"Ov)j �47,���)�"O����E�q�0�bL3ή���"OB�SW��h�Bw�0#���4"O�qd)�!>ȼ��V/���"O�q� �(��1�j�2'Z��"O�E��	9@t`�i'�x�y�"Od���#&�l-��-J��L�[#"O�A����7� ���Y�#�=*�"O�KAN�@�0�$e�:'^Q�"O��xA�#3����j�<.���"O aSQ��-x�����D^���"OhDX�f�8q{AMH�H)�.�y��~#�e�юfr��7�҄�yl� -�T�&a�1^��9�͛�;�ў"~�K�h݊䥒 !��M
(��e鈄�ȓ#�܌P�ʎ"@02%( ._Q���I8��?��A�J ��#s�!ҵk�n�%�pK�e�#{[�m���-6P��G5D�LvL�j��DPUa׷aox$)R�%�HO~�'O$%��� �=�g�`�d�ȓ,��}�ՌS&N:�9"�<4ep�Dz��~24�B�?���E,��lcB0�ai�D�<!� �<(�5`FjQaY�+�e��<����S�	O�Lc@ܻ0D�1��F�B�ɿa�΁����)$��!RN���ʓ�0?����`�q���3�Zq�Ҧ�S���hO�u|�	�!ǔH� p �^�p��1�ȓ~��飋�P0H���,��  ��ȓT�s��<B>�� dɐ>�p��1����K���A#�A�(޲�����5��)�~q�D�	����v(�Ժ����A��9�K�=e�V��ȓi������ �<���FV���ȓ5��9q���A��ѪVHl��1��d����?q�l�`Ǐ.e�Z�ȓm���RS��̍���ؤN\�Y��SF��1��Z抅K���{|���ȓ���`���=�@�Je�Ȟ]�����/� 5�$�(i�`�.B�%�l��ȓ%7>Hc i��5N�@R����p�ȓ%������e��Pf�ٻ}-�ȓS�>L��(S!J����7��8"1���ȓ��ڢe��jiHGm�"���ȓK
��R��e���S�,� 6<�0�����h� �Q<z��ɐ~<�܅�q�h���$\�
�0�aq�A�R#�مȓ&�܌he�
:t�,���|i���J��HheN	,>V��!�J��!j����	���X*e��Ś2�I'>N���yz��.η8�|��Ph:/B��ȓc0u���!L���t�:K쨥��Y���#�_>�б���N�T�@�ȓB��m��*��e������E?NT(��ȓSnx��ْh��x�e��\cHm���\[6��(-���C%/�!f��m�ȓ*-^шr�T;��$��Lq�8�ȓ]u��ه�ޘH��,kF�Aj�&Ѕ�6O΅��"�ޚ�҃�C�b�ȓ8G��Q��R�J��9����LW����S�? �Ũ&L]9x<�#d�]{��m��岶��d��P��h�d���F9EH�NU�X�[�,`��[��t9�ޏ0�����
t����I��Y`����<�G,Ə{%X��	̟��	����I؟��I̟��I͟�����Mk�hƞ�5�eI^!/?��	���ş������	ğ��	����$#�Ѐ	G+�\X �Pi�9%�IƟ��I̟t�	��4��ǟ���؟H��ek�ȏ N'T�#'(Q10 ��꟰�	������T�	��`�	����I�E���R�W�s���jF�'1��IΟT�	���Iԟ��	⟘��۟�	�{mFl���7�����։.]��	�����Ο�����0��ǟ���ܟ8�	�F��"��C� S�P�A������	Ɵ�I�����ğ���ܟl�I<:w��ڰ	��L�� 1a�v[Y�I�X�	џ���ҟ�����L�	ߟ(���AD�FbZ1uE�Jf�������	��ݟ�����������I�{��y��%��M��,�=m�>��I؟�Ŧ!������	ٟ0�I����ݟ��b,V�ΰ�ˤ
��3����8�Iԟ��	�p��ҟh�I�<�I�� ����<P�$,��M��k�\�Id���������	՟d���d۶�D E�PaP����F����C����Iٟt�	��l��ޟ��I6�M����?�u�DNE�Jˇiۆ%E],)&�	�h�����d��= &�ڂ3�$��E�$hbp����b���!ɛ��4���_�-*V)��X�a���js4�ql��M���1?��[ٴ��$C,'	xrO�4��S� �����
� �ã�T#�b���Ipy��S�,��s$���5��\����39�D��4{�$X�<���4�o���:>z�U�c%J�%p�Z�d�Z��o��M#�'��)�S�B+T,nZ�<��Y
:��U�$D�V��ؐb��<�K��pH�P寅��hO�i�OPi�4�_q��(8&$�g*ұie3O����]l�D���'lpY�v��z�B�!�x�}���Up}r�z��n��<�O�@(� �!}Hx�Hc���<.aiT��X�,�'��`��M.��"�tx�;9K���KW�ňA{k���!��;/��	Ly2�����$Þ);Ĝ��À3 ���/]�AA��Ӧ�p>?I&�i&�O�	�L4�y��=ظ0��W'�DWئ��ٴ�?q֎
�M�O�0��R_|AHFW�(N�#$�� ��|X`mSpr�=�'���,�I��P<��1�"�8��I2�̒�i��I��M�'��r���O���wДH/�e:�۪X\�4(s�>yG�i��7-i�h&>q�S۟��!G�8�峰/�8u��śf�&�D��i�>iem�4O�h�%u���O�Xz�Oܼ�@�&(ȡ���*w�daW��Oz˓���-�$Y�1���n�h{�E�4&�ؑ�
��8ǭl��ڴ�����'8 6M���=�I�h�h��LսUaZ��n�.4<h�h��ͦu�\ȭ���ӎP�,1��?�������m����46�
�kT��#^8p��'i�]�|����Aa͆�(��9��g�2m@B$94�����EHr 6?�p�i��'����Aݡ-��q*dƅC�Myd;O��S/������^9�7M�����(�;pp���eFԸ:7�hǒv��B�D?ZH�#q�>}��0?�'����O�Q*�Aƭ%�������S��08Of�O",o�0J4b�P�O��TK6f�{��Y;��E*��� �O
��'G�6�ަ�͓��OzL���A�a콐�ꛤ�.��ń�/��|������4��y�nkݕKM>�5�b�T *l�B#�?���?9��?�|�(O��m�JѮU�&�H�z�̫1%F#�h���Ey��e���쫩O4�nJ�����a�
]e��a$K�0آ��ݴ�?q4Mߗ�Mk�' b�;E�n���G�2}��84���'ذS����-`V�My"�'5��'y��'�rT>E*7�Q�|���PǡQ=LI�q��E5�M�/	�?���?�L~�Jכ�w0��ڗAϲ/�a���u�r�J�~Ӳ�mZ�<9�O�i�n�Ď�f7�{�����$
 ]i��Ap�hCp���.����H��WO��xy��')���YLNl���Ȃ9<*Aൄ�p��Ɵ��IKy��a�T|����<a�Jϐ��`H�0T�~�S��@C����E�>��ih�7�m�d�'&�	�$ʭ�z}h�+����B�'n®�;f��la��ݱ$���?!9����w�'*��k���P��EHFH\5|��x�'�"�'���'�>���7O*R����µyq�dQF'I>9`^]�I��M�3ٕ����ᦡ�?�;r|��`�T�F�Y�瞉P��`ΓoA��-lӔ�d��P�l7Mn����=T蕀�?}
��*���||bĆ۾K@����{�y��'��'�b�'�BH�C�D���b�	j89��CQ�*��I�M3��V=�?����?I����9O�yh�E������>_�T{Q%�]}�m�Љo�<�K|��'�?����.s<!��,3�І_K��y��޿��$XN�թv��N>)Or�@߈x赳LM:i=�������p��럀��˟�GyBn�^M"g�O����D�V�8P%�45ntK�7O��nZʟ@&� X�O�-mڝ�M��<�̡�NC6��� Uj�d
0�y6i�-�MS�'��M�&�Ё�a���n�I�?�1_� ��*�IR�%}��*g���z��6O&���O.�$�O\���OT�?�{d�iF�p ϔ�qW�����	��T��4u�؜H/Oxhl�E�5�~T�r�!	��؇�ɩ�~����dN���l�՟tPui����͓�?�f��B;�HҮ$%<j�._�n�5�Q�غ)k:@*I>�)OH���O���O�,�+ͼ1b�1X@Ll#Ұ	�o�O@���<iQ�i��i�%�'���'o�S�v�y�gŐ��@C����Y�I��M�ղi[�!��,GeJ,j��i*s�Ё}�%�.@�	u�eDA�`牂|�TZ��%c�����i���6�(�I�U�w2��H3hLԟ��	ȟL�	؟b>U�'A�7�\�tؾ��f��4�|�Y��	�Xv��r��<1s�iN�Ol��':7����A⑄x,\Y�P���lZܟ�СdCЦ���?9�X���bm�3��$�3=�����A�:��X83�?P��$�<i��?	��?���?�*����ޤr!\jpE�<�^�	G������Kyr�'I�t���go���[� L<(+&�ʛT�|��J��1<�m���M��'��i>��Sڟ�a	���ϓR�hu!G'f��t������̓gt���L�@1�	�I>�+Ov�$�O�Qiӣ�:b��@�+g�̋d��OR�$�O��Ģ<i'�i	��Z��'R�'
�Q���0���o����ə��'��'E��@
��p���w}�&�� �Ty6�T�Q� �gU��y��'6Jtm�u\�ҴV�t���v���;Mh��Q�D�>�#F�S�zΠ�#��ĞK���'���'���py秕0��ڀ�2t{�i w(՟@H�42�A.O�o�ğ�%��]"w�P��}f(�1�!�&:>�I��M3a�iH�n�Eӛ�=O4��u�\�3dy(:)��k��->�0`��6[��а��3��<���?1���?q��?�#�!.h4Xb�c��)� @���Q¦9�W�Xş��	ԟ<��q���'Ka(�"DČ]򩑣g)N�����>!`�i_:7ͅɟ|&>��S�?��-�1̡ ��A*^�r��$ۗ<�
�!$Xy�Ɩ>`�����"�$���'��닫;�6);Q�O9`���Ѓ�'�R�'#�����Z����4az�����<��];V̖�MBtU82�.s&�9ϓܛ���Yq}r(b�Llޟ`
'��~�k��?]X�"G���mR~���7��R���_��O����h��H f�!T�|��і�y��'t�'6"�'����ܞf�HI�i�0q��H�@�����O���Ŧ�Sp�c>��ɬ�MKN>�#O��_�n�X�i�$L� �2���,��&�rӀ��G�w%,6�l� ��yvm���\�"�R�*1���T�LDN>#�n�	]y��$�P��d�(#�r����.f�,+ٴ(B�PA���?�����V���KCB��Cyt�AA��	22�������˦ك�4E뉧�)�@PtE�B�$]����PO �$*�2�7 T"U*w%�<�'�T��\wWؒO��v��������!#�,�O�Ln� �����$m�
 o�%h��A
 
���I�M���(�>�f�i�}zG��+=��q�ʯOތ� �p���lZ���l�~~"m�"��Q�i
��I6@�)i��[�r�P�L@u@��	Ry��'R�'^��'-�R>�rτ�Q��e9W�ȼc�����α�M�2�Ӳ�?���?!L~��Y���wO�A��</�ܡ@�i�3MD d��@o�^�m�t�i>������ ���Ϧ�Wx��1�#$=��)6�U;���g>j%�fa݄a�V��H>�.O8�h����3�Ë^LX p6��T�8��I�Mk�X��$�Or%P�E�"l��1���fuL5�j7�����٦!��4L�'��1x�욘ay��	��H��O~4r�"ַ}T9b9��D�rt֝��?�d�	�K+����?6(�%��`���?����?���?э�	�O��{D��j��-�GWz�B�8��O��mZ7%���'��7m�O��O�9Z���rGݎ>�Fܐ&��7'��AЦ��ش�?q�j�(�MK�'*����M3��A%��-���.]���cu�#2zP�ќ|BQ�0���X��͟�����W�x�~Dy����,Ӥ�oyR�|��`�&�Op���O����S<U��m���ѧS�X��'������'N(7���)K<ͧ����q�xe��ۛ2� ��͢h�Reb��(ma�*O�a�����j���&�䓪�d���y�o��q0���$�-�����O����O��4��ʓe���A@��ʒ��6d[f�r�L���͓?w����[}�N}��Ln��&O%)�5���'�|�JC ��g��oZ�<���[i��č�IT4�{*O>����N�2� L
D<�|�`۹hP�B;O��D�O���O:��O��?��nA�$F��*�#�9+��5Ò��h�	ퟬ��4g��m/O��m�h�	�u�@d�%#L��zT ��E1�JO<)s�i7��&��`$c�B�ԟtZ���^�d�)ˋ���pZ��[���J��Q弼&���'���'��'��z��O0�U��X�9$Ȁs��'��[��i�4$	����?�������TmN���KN0$0��y��=\��(����ʦ]��4l���d�OH:����ގ�t��6/��,��-���C�T��4�����I�?�3�ús!�|�B4��ؠ$_4� ���	8��'W��'���DR����408.�����Q萈��.\og�y�#ɸ������Y�?��^��R�4z�����(-Q�T��"�6KE ����i�6���6�e���I��r�벧]�Ҷy��� &��e,W��0�6�X8v��]��<Ot˓�?���?����?1����)�)O˔���T.F�*a���P�*9n��{��������t�s�������g/�'rN�����-K�9K�[����oo��%����?=��+N���o��<�/~"���3v;F���B��<i�')Z��R���������O��dP�c��1 `��/�V�8�O����On�$�OZʓQ%�v	O5��'�E�Is8U�V��5XT�Q�5��O��O��'�z7��ӦU%�t�0Ŕ����l�k�bT�amq�����hA9˧�H�Q�|�'��$�#G��|���\�u�T��ΪWx�t�E�-D��xD���'�1]`�)�V�ʟPXش{��(.O�Yn�E�Ӽ{�K��8Bh�o:��G�	�<�3�i(7Dۦ����٦��'�4����ɲ5�үJ?�<	奊')��Uh�K�9�F0Q��<i1v��+^�L���a�݀}�W��1���(5I�3�6Б��38'6YR�+<��l
'�S%6���b0�8<d �Ѝϣz�%�3�)�9s6�C;���ꖎ+*���E�y�plk�ݻ�.��AmB�qT �g�������i�8�D��i�4�KA
��~x��oG�mlp�0�LYE��`*gLe{`5�R)P
�l��7��D��q���T�&�:��`JTi�@ ��I
qS0���+U �E0�D[2	j��.-tf A��)�
"=X=� �!v������M���?9���"C��0��.��׍��Fmciq����O8M��)�S6�> ��b]`j�qD���?	�6mNMK�o�џ����������|r���:dlqu!���Yd��'jA��d�9"���T���?c���	�	�4���/#٨����ŃR#�\�ܴ�?����?�t+F�����$�'�"
֠6x�]i�lݏl6����`��[���?��o�8)�<���?Y��<�}r�Ý!.�T E��<���ҹiJ��L�O���O��$�<y��8}��X2�eLJeAQ�@�㛆�'"�y�'B��')�	o�T�+�͋9�AH�K�
:���I�ē�?��?9/O\�D�O2!�A�����q�q��vq<�%��1C1Oh�d�O
���</����)�nH�s7lP�,�ИG�$�	����	|�I{y��������'TY�d�4K(��ND2l+�I���	��d�'BBa �+#�IU�(�Ҥk���O��옻w�T@lZʟ�&���'�z$����k<����iQM���VM�$�MK���?�)O�b��Zu������s�9ш��c��2UC�'$hv!'{���?I��a��E���M+�$2�xhz�ǍT��e�� ���y�'�J�B�A{��I�O8b�O���z�@J���5�T���OC{��nџt��0]\�m���	���'�� �0�$Se��F�.���ݴ���Q�iW��'���O�LO�i݄H��pp�BU�-��F��r���oZ�C������9�9O��D��5�IH 䔵�:$��g�?d�"8n�Ꟙ�IƟ\b��\����|����?Q%���[�R�`C��.S��&�5jf�I۟���6o>�c�0�I���-J��a8���'ɲ��͚V�nl0޴�?�&-����$�'X�V�d8 .��l�l�A�MQ&���S��M���x��<���?1������21��ai1��\T�%�B�E����(�V�˟h��L��Ky"�!T�Z�B�<X��t�jt�J�y��':��'*��R,ʝOO��+�큍rs�����s�
T�Oh�d�O��Ojʓ�~��'��Y��l�
z�4��g�w�IJ�O��$�O ˓�?Y�����i�O�\×��`i�h��f�f
Aۅ�����Z���?�N�N�d�'�l�T/��E�"�svK�hn�:#�o����<q�h�,$�/�|���O���\�*J����H+�J�K,S����>��u���\�S���[�K^��F�8LrUi�,������O0�����O0��O������Ӻk�Ț�<�^��f����p7j
h}��'b�PbIY����O�
�X� -��� ¢�9����4d� Z���?y��?!�'��4�r����s9�Lr�PUЦ��e钀i��<oںTʪ��z�y��I�O�L��Y��(4�6Fj�h�8�n��IǟP�	�'�	���4�'�"Q�$��F��z���*!v<�[�ʙm̓rD]�B����'�"�O�����˥f����E�قC�izk 4=��Iޟ��	����=�b�ǝx��49� R# Z^i���L}2O>o��+�O"���O���?�玆�T�b�-��*m\�扑)r�c(O��$�O���#��ן\R�&P2S���KO=4�: �g�"���Ī#?1��?�,O����8���S=Y�䗒�޽7F�SϬ����i�2�'�b�$�OnD���9M��ɾ_`zŲ��T� �R�k��V%����O���<���>O��b*�8���/_�q 2Fŕ6�� xE�M���n����?���ayĈt�k�	�Nժū��ٖsj���I	[$�[��?9.O �Ę�6��˧�?���*V-J)�"-��r�X|��S��O��$K�{0Z�qC�T?ɂ�	�U�ʽ�7H�-qĩ�"�>y�<�l,a��?���?a�����R9I�j��0J�rt� ��u`�\�����,T�0A<�)��>\��(s��:�,��[
Rϔ7�]�u����ON���O��i�<�'�?��#aJ��m� �1��Ȟig��$�"<�|��MJf̈6�ێnᢝ�dA�3��T�t�i�B]�L;E�by�O�"�'��� X�q��ɖd��:�`�9 ���#�oe�'����D�O��	d�`9)$��76��iց;
�7��O�У��<��?9����'�`��BM5������;�B5
�OT�G� ;���֟t��{y��'�X`���i�~��h��s���(� nh�	��������?Q��!ʠ�hg��?c�u�Q%��p�� X��	y���'��'&��̟���j"0��
��Ҁ �]�XB�N�ܦ�������I^���?1S˂�6���oZ8<��8)Y�w���G�x&���?�������OQ��O�|z�'�7e�>h����&JBq��4�?Q�r�'�x��Y��ēT�:�� �߂+�H8 ���EϾ�nZ֟,�'�B�بZ�S՟p�	�?5�! ��{�ԄX�w���YsO���'ib"��c�̃�y���91�ת� ���M[e��AX����\�b��	ş���Οl��YyZw����e�qI�����J�$��èO��$�L�Z����Ӱ�4�a�H��)
d���ig�fN�Jkb�'���'R��W�����`�
	�O>��iჅ}i���R���Mcr��
E҂M�<E���'�>�K��ɘ*8t�׋���D	�Ric�L�$�Or���&E��|���?��'C�X��+��6*�P�Th_,ih��«3扜H.��M|����?�'V���DK�!.��jDeבDnHl��4�?��6��D�Ot�$�OX�Ћ&hQ+�U���ЭH���#�>� fT?0x���'���'\�	ϟXi�S�n$�aQ���.�a3	�f1q�'5��'�����O��f�N�V �dS�$�_��E����d����ؖ'��ÖV/�����es"�R�nx  � E���'G2�'�O���5Y� �3�i��xbEGB3w�� !����Ol���O���?iF���ɬ���a)F� �L%Rs*F8J���r3Bh���d;�����Z��
g�O���(�.Ř$�2�L#$�́���i6�W�$��1[��I�O_��'��4 	's� � ��+G���	� a�rc�`�I$
��0Jt�<�~��鋉\ �:g�ˏ:4��k�f}�'oD]ذ�'#b�'V2�O:�i�Yu��.�x���R�h�W.�>a����hu��B�S�(��|{0n[�j�8��Љ'R�8n�!#�9�������ڟ���wy�On��$L�����Th:��0�c�6-B��Deq���Sӟ`I󮄓o����B쐥� D��M��?���"��ȓ+O��OH�D���3���yl�lö%�!`�h�a%��ܘ'�9��.'��O��$���b��ԣ�v�s�n@?T����f��䌈z��˓�?Q��?i�{��-#�|""��?�b������>TQ�K㔟`��۟<�'��շ?�����N>:��q��#:�>H{Z����ԟ��	l��?!�&��QZ��C�����������[�k�I��8��dy��'�I�0ߟT*vH�J� c��Jb�$���i���'B���O�4�c�Yxj���	5�ԁ�!�\/o�~i�B�#����O����<)�v����-�
����(숉,����h]���Dn�ş��?��$�1:I�_��-d8�(VK��b��PXToQ�{��6�O���?	�����i�O�����P��H���T{�����\��?������p�<�O�ic�'�z�� �NY77n��O��r��$�O���O�ɲ<��Nj8�dGW6}��C�e	r���'��KR�	�fm؊y���H���y��%Z2�d�Q'��M��ݾ�?���?�����)O���Odh`�G��� �tWO�<�lYͦ]�E�۠{`0b�"|*�p����}F0��F	h`�ғ�iK2�'BA�%Xk�i>}�Iݟ��/W8�� Z6~��ua�E\�(	��D�b���&>���ڟ��� g�*���l�'��Ĩ ^rh���۴�?����d6�'�2�'�ɧ5��B��ک#�Gk9��I	�M�7�fYX��?��?	��?����?I��^+�@P,����7��w۞M!����O��O����O^���O�i���U��+0�){�F�7m�����O����O����O:˓i�����=��A!��Tg(���邂>��MB�i���ߟ��'���'~��Ν�yrY�i70d�3��(�I��>~Ԇ7��O���O
���<1teC��S����)�U� �����!=�~x�wd��M�������OB���O�K70O��禉;b O�l�sO�����	q�>���O��N���AP?��I�� ���0��钁�t)@2�в1� ��O�d�O��d� 
~� �d�?Ғ�6����/�y^��Ah��ʓ;�ƍsƲi��'�2�O6^�ӺKVn
�d阝�r���,���*�ϦI�I�`������'�Ӽ~D8��P�׵u�*�!ɩ]�d6-ْ0�nϟ@���t�����<�ÉM)-1~Y��;J�|zc��A�&���y��'m�IV���?a�K�WQ�ܸf��{�4�k0�V�����'�b�'Q:�
S-�>�.O`�ĸ�
%�K"�|�""�]���"Bc�N�O�]�0O��Ɵ��������ˆ(G�ƹ�f
ˣm��܃�V��M�]r!��]�d�'�BV�`�i��1� ?L:�Q���cV�ї�j����8~��D�<���?y�����4w�U����N$��¤6�Lňw��U}�R���Yy��'b�'�� @���N�tLІM2�09A���<�)O��$�O��d�O��Z�C^�$mڼw�n�iDI�(F�(�qM38�m��4�?Q���?���?i+OH�$GO���M�.�m`�oȝ$ǌ�PQВz�JIo����	���	)���(+�\�lZ����ɣ��\��)���Rz������4�?q��?.O��DϛND�i�<�4e��V<mX���_Q�L����H֛��'S��'��! %Ϫ6M�Ol�$�O���s-���O����1?��nZ󟴗')����T�'p�T>7m�)A�9Q� _40	�r��=r��6�'+��&i�(7M�O��d�Or�	៦��U�q�V��2�Bċ��ݞ+�PY0��>���4�}����|N?�5�n�P�+<TԛՈV�R���$T:a�l6��Ov���O4������OH�d�p�ك$�U�4*n尗,��FJ�Hl�:����I�`���Ě��'���P_��}*��"'�
�$B���M���?Y��KHz��[�|�'���O<�
O�6!���3� �m�i�T��Ed��?������!W"���GS��*�2��nZ��"1FQ��D�<����d�Ok��Rn �ˆ�P�&��ip�����	�!�H��Zy��'Y"�'j�	�\����@lӅ[7�1�r���r8��T�^�����<!����O����O@�R��*lK���!��:�ek�jD":���O��D�O��D�O�˓��Z�8��0�*Y�����;>�`8+d�i��	Ο��'���'9�i�y��
y�>���J��y7$J��7m�O��$�O��D�O��d�+��o�ȟ��I�O�t�Pt�yȸx��#M�-�t�ߴ�?���?,O��D�}U�i0}�͙�cvԑ"��<x�'.؅�Mk���?����?�$��7C�F�'{��'N��� �|ߐ܁��>Y����Ɩ�r7��O���?a���|����4����F,�,-C�MA�m�B��u���M���?�U�R�g���'��'��t�Oq��F�8<�c�&H[��qi�l�!C,ꓶ?	a���?���4���O��@"�N!W�x��S�o�B1��4Kj�ixѺi��'G��O����'���'������X�p�:��PQ�pp�kӒ%��n�Op�d�<ͧ��'�?���H�(QBA���	�4�с��
)LX�f�'5��'d�,�f�>�)O
�d����
D�j`
F� r�ˁ�h�P��<A���<�O>B�'��
�	k�����hɬ>���jʟ^�6M�O��a�G}RU����yB��5Fg�*Fz�n6��dX�"P���D��b����O��d�O|���O>���c�C&+vp ��$�X�15��4j8�	Jyr�'��Iʟ����2��5'��h3@��+o�ݺ�B����?q��?�����d ��N=̧��2���!@)��Brʆ�ZzZ�o�wy��'%������	러3vb��*s��a���1z�� �C��q��7-�O�d�O2�d�<ac����`r'�H\,�!Pu)U�D9ȕ��C���M������ON�$�O��H;O����O.�� �8H�T�&ϛ!�4\G ����	ܟ���Ɵ:1 ��M����?����.ۻK#
��cb��R����3�*%��f�'��Iܟ82�k|>��iy��MKaBߥm�DrVb�a2�*!'���':|dApӨ��O�b�O�+�L-J���(k)60�Dv�fm����`Ő�	L�Fܧ=d�3�ܒ�Jd!�.~H��l��!f�M@�4�?���?Q��uK�'H� �1|��i�4FN	)������<X6�#>���4��9��şdK'�i�����*X�@�{�/��Mc��?q�5����x��'M��O����&��" ��K$���i�'�쀀&�'�I��T�	��=P�m�5}k��F��H�26m�O"Iq�n�p�ߟ���`�i�9�!�} �L� ��	���r�>AQ�5�?y(O>���O��ġ<�5n����,�1oԸ|Ml��%CΑM 2����D�O��O~�d�Ov���kGx%�d�4��#Vg�#���<)��?q����oef5Χ*�
�a�B�)��T �i]�\��'?��'��'>��'�98��'���׃ׇxN�q!���u�n`����>A��?a���D�)�2$>�����b���c�}ժt���M������?��)�ѩ���	;L��K�[�<x"�P"f��(6�O��$�<�4L"K�Od��O��7/ʦXsP=�!��'z��( � �d�O����)����.�T?E 6#߾4��H�rE;7���qE�`�dʓ"���Y �i+
�'�?����'a&���!�9e���	T�ǖ h:��ߴ�?9�'������䓹�O˶x��MH�j> �"����nN�D*޴25�I�g�i�r�'���O�O �K.SI|�6�ư?��}��kM�|��m�pJ���	q�)§�?Q��#dU��qɋ�����+�?���?��S ��r��xb�'���O�j�H&�Z���.W�	b��r�i/�'���qv�*��O����OX�0ń�e�ʽ�ІϵD��k��KӦ��I�O�P�N<�'�(O� A�Ȫu�2�AL^�N2ܸ[%T�X���͟����������oy�#�jmP���:*\�E3r�H�q�@���6���O��=9��m��tXa�р&�X̀%+�MG�8ȶA��?����?���?������8"��$�5Z��� r�&(�N�{�jS�@��Ql������џ &����џt:�%�>q��%FVq�M�w����BFM}��'u��'���'���x�V>��T�y�q��hꤰ")H� oZ���%��	��*2d�"k��O� 0����U�b�HpcG׻s��R`�i���'o�I��h��N|�����-ڇ@�6\aF��>I�*&�ؼt���D
�?7 �"��q�F�C�.[���$؛F�'o�ʌ�i2�'A��'��R�֘(N��qG��m�l-�1l�\��6-�O*��Ӈ'-x0"u��)�#<�{Մ
v���j�@�c�� �x]�6�O����O���TS����0f��k'�����[K�17���M�ŀDy������ȵr�bt*���q�T�D+�[��,m�ǟ��Iß4��Q$�ē�?a���~B.K�,�:��d�&J��=Z���/��'x��k�yBo�!YBL���V��V�aGC�#5�`��"H�?5k��l��o\��2��2�X,�$N�z}D��8 ��=�Q��&��f6��C�(�*3Ѿ�iK
�iR섆�'/~�Ѻ����?�������.'�݊�h��.M6�QF�ք�AH3!ߢ�.HH��Us�2���:�}�Qj����ĩݞ!l$�	��H�N�*�j�A�b�]��S�rB�J��ħH#����#�.O���L�Z�t,*d�!
f~){��^=B d�c����l�4��lVR�h$�V�l�����O��2�E�O|��p>q���@)u{�Eie)��[ʬN�^�g��	yj�p�Fm����^�AD�M�h��\ѲD�~y��ǐ(W"�h���x��I�	G&�y���v����Bd≠(0����nY�A�tI!GBJ�-��C�I�+C�XZ��8vB��ɀS�C�i!�4m�:�)
 jj�� Wk����v�	�y��h;ߴ�?Y����	���]oD4�ek��T��P7C����D�O60V��BTf�Q��RY-��5�͈c�
�)�e�|*��	ui%!���f�ΐ@��y��6��%�j\C�qyB��#���	����i]4>�j0�F��lMy�n���$����,��S��%�.���؉T���q�5Lf��ȓ�49H���K-X=��)ԭmK�ት�HOv�!���(`��e0V��0�n�+%�����	������8�\���H՟P���X�i��k�P�sr|u2�̖\S�3�ȦUњa1��ڼ@Ά1i$�<32��|B���]��	��=��b��$�;~˼1��K=Y�:���FQ�tĴ�Kg[��O�!K��<! M/)"�m��$O8�[���?�O |����54�ҍ�:f�ػc��/J�B�ɎS�<��mX,���o�C9��'ϑ��Sʟ��'�f@!�	.^u��G��D#d��q��r@s.Vٟ��	۟����uG�';�0�ȌiV.՚A����d�B���cU횳4�^�i���ksbQa'���l�d�B��X��(O,��F��
�&;EaL;+�.�B&F&Cy,��򪎹wq��nӈT�w��5Q��YP�Q=�<9�JA�M.Ft�k�<_�\���Ov�=����q�r�R�}�� @�R
���'���x��8+r噴��]�6}�yBk|���d�<11A&_�F�'�"+Y�wC4L�� WRx�"��2�'7��IE�'�:����6��Dj�|Z�Ǐ�9�\���VA��T�� T�$	��*Ƥ��GE��(O���D�ΤI���1�j��4�F����/x�84�G㓴~��i�.�(Ol@aD�'�:O��E�C09��%{"�5�ЃT"O� �A�%^��%j�u h�On�l���6�*�O�&cTp�f\��N�%�Ly�j�2�M���?!,�������OL:��˓	���J6f������O|����`�$/i���

�|B ��M�Q��˧c2L��G�^�nl����5���OHa��͗(t�Q���0�6���P}ή�2͟2!����`�����Y2�f$�Ԝ>�q���XL>�2�B�
5u2��L�"}��mn�<aeH\�tH*<8f��D����P�X���D��Z�pɷ��-˼ ��G�10�m�̟���П@�,��W�v���ϟ��	���7�Z������lI���S�	�$`@ ܇���Iu\�� '�.�3��ޛ3�����;n��l����2%��G��|z���.+��y��L>	���+{�ES�)�<� �h�dG�'��H�S�g�I�6d�q⦇L�o���3Å��B�	�OeLEɖ(P7s�p��!�j�����SW�	 ����ķp$�00vME	B�:<	�J��8�Vx��Ɵx��ן��]w��'>���0�sg�7S�T)�΋�>�h�caS8CQ�RF(X��Zr`*�b�9B��V8B��� �� ��FY�H$ e�4�R*�Ƶ��l�}r�G��~w����$�0;\ȑ{"C׬r��1a�e��a�i��'�v����'_��=� FF�*a�@�^=4�!�$�2쬕a�*�,JՖ9�J�:?�1Oh��>	Wl�40��؟�#CbI���C�J\��0rƌ��0�	>T��d�I��<ϧ`�"\"֭�o�J�C��I��M3�U�&��x[��Y2���&�@p8������P[��1��Mo�0�z,�J�)D4��t��"1 <��Đ*���'���)",�!�u,���n�6O.b����sx��@��S� �mj�]�M����c"���4
��Z7,��.ES(���
�����d
�`�&�n�ǟ,�IO�T"��z
� $�'ғwӖi�Z����%�O��d['6�d���¸I_�����w�Z�jJ9���'C;hQ��@�{>���G�,Х�O� ئ-�Iu� #q�J#D��hKk� ��Ο\�AD���l���`�<�.Ѣ��>y�����M>�zvf�iy�BH}cV��f�w�<� �	!���e�߇6-�(���M�'�v\���
7Tt�S���bY�)��Mg�.�D�OP��Z�j���Cd��O����O��4��*p�ш�.<(��@3l$�4,Դ;W�=�����W	�˖b�vc>)���AA��D�<IR���+�.f"�3�"�:6�n�Y��[�I�愹1�L�#"b��	W�!E�5��'����Ím]r��#�\�CW�����L>Y��+b��|��aY�ɜa��r�<�!������;�KW*y@��¥O�p~��(��|�O>f���z���{�� 8JL�7I|�<��'S8�?��?A�����O���{>9��A�7���ڲ�S�
u����*q��Y`/�1��>AF�h�S�Ӂb���񗨘�>"����B� a}R��(�X|�ϐ_8�<����s�����|�ah	&-d(T�pd�9v��$�C�ڴ�y"k�(���1	V)j@^�*t�'��7�(��œI�jEoӟ���;u"a��F�-�VA�&�Y"���	P��������	�|�c��h'��h���Y�V���8;!�Y��+O�;2��Y66��}�MO�+�&@���А)T�x�%W4�?!�x�E��B��� ����kT���ŋ�y��C�?�d��c~���X6F��xB |Ӑ �CJǟ��E��Ȟ	!�K�.)��S0`E6��П���y����pBR��w�N%��n�zg�Yp'��l���'��e�4 G"P�M�ʧ����M�xH,��9�
*g�
4�V���ܣs���铏CZڵ+T�^�.,��!5-���M�	���S�'$R�"Ҡ��`�����H��P��[W����F�����C	C��%��	'�HO�)s��ϔ4�n��b�9\�T[�����I�D����{ݟ������i��h�c�6���Ȣ�X�S�d9waו��4<�8�E�O�g��?<� �� _���k�#T�oȠY���߀~����uR�%�V(6�3�䇑{��M���wX@��ǫ�=A��%����+�Oq��'D�rk�CW�$���L�E���'��[�F�5i���H*@����O��Gz�O��'�\���̜�\��v��!�c�,� K�tp@�'#��'�r�l�a��˟,̧m���思�4�: QlAN�J@}az��Md��A��	.�2Ћ⁍�/T89�Gj/n�� �M5x�аa"�L�>��dZ<�E���;o�T� ���~`͚V�'�.7MKʦa�?���ހ\�q{��R�x��8���b�!�$I5��r�=��P�Ōv�1O2��'$剐|M�MR�4�?���C4�9�%5:f���Z[���b���?Ag��<�?����� �)dN~y±@Tg� T���UmNĊ�&X��fG�-���� 	��xDyR� T�$�5AI�H(z�fD)^0�P��l���|�*UB.SVE=c�ȱEy2��?�$�i�6��O�E@g�v�N`�c)�����<��������s���{.l	+B��A5pqZ�O�	l�*y���4,J+`��[S�E�]����	Qy�KM6;t7�O����|j��]��?�������č�
kB]��%2�?��G����F�� 9)��U�ʧ��.P�q���T�"�j��B1��<��A�n�P\�A�FM;9�t	��P�`���'8{�E[$ ��%SH1� �C����O��b��'��O�z�[�BQ.I[CkP�<�B�C`"O4yp�n��oA�i��/N��!��'tR#=a0��(ܘ1w��)Y� �0�)r���'�r�'�(,C��W��'3b��yw�@Bd��p@�HI �Eif�)*yƴ�����R�1����XF�"�Sb�I6,���@��_$��6���[BR����P���8q΀�u)��"!��a��^�bI���+"��C�-�&�`�M>y�-�П�>�O�}`#O�-U�ps��LNj�� &"ON�BF�@�!۴���@Ux\����������4�V�Oj-jW�Y}���à�;M� ��0��*��O��$�On�dѺs��?��O�p�QnZ&~bm��D�	�J���+�6.�~�'�#,=H�3�
^�џ��V효](=�DfO�Vے�ӂ�Ų&f��c_�\0(��/� l��FRj"���35*��l����L ���o�a��	�D#�憘q��x)R���y�˱Rt�Y�0L�A���TI��'�,6�2�ğ�4��]l��\��>.��3b�O�l w�:P�	ş,��ğ����|���ӛ-pL�ĥ� gn¤��>� $�q��٭\y���w�X�n<R��\`�ty�v�I�\{D��V ��1Ĭ�[�E�`�|L���0d~U`��H.t�<`��É-O��(���@ 2��7�W?�0�Bv���l{�y�w��t"!�׋��d����oh��P�(!�d���f0^���Ɋ0N���%�P�ɣI~���4�?a����,���'oo(!1�|L��Z�Jg����O�jcH˄]�p��5c�:XOh��Bj�t]>���&Y�NP8kq��M�DA��*5}��
�|	���Q�!� � /�WA��2hѕ�	��11Q$N�1��8B#�>Y"�HݟzL>����V�-#RT�&�$(
�VO�<y��� |]��۳&��~9���J���DDc��.�0�<:%FP�mZ���̟�
M�/cg��	ӟ�����9L6�� #P�m�|ͫ���R� ��<�sEI�<��+�9�d	%K�I�ʴXp%�z�b	���	�}J�V+�-���X4l����D��������?��ǒ\ȥ��'U- �2!L �	@�Q�'�(��E�1sN��P�	b ��OaGzʟHʓ ���F
�f�MJb�K %Xd�4
X��c���?a���?����$�O��Wq�(��f��*��J�#W*d��"��Q�
�c�8	�Y��)��j�q�C�Ia�$�`n�P���F@'z\1c��OtL��	��Ƞ����>�����߅=.�B�ɮP+\��'iɵs�Hp�T�����c��{�}�œ��6��O���-��)V3BH�D����$�Oq��C�O��d|>Ÿ�/�OV�O�9���0��015a]9#p����'��pb�2���?�B #Ũ
0~�F�+�&�4�p<1A��xM<�ʍChhTP�R�,�l���MP�<��`r ��]���!@t<�B�i���+��j��I���@�U�X{�ybO�~�6��O4���|�c��?Y�.S���p��0�(L:r���?1�mızC��h>��O�Q����)~sĨp�ׄ]�=�����0�ԐzEbŵxa��'	��Tcwk^� �;`�Y���<jf���YZڴ�?ٍ��"��^��@�Y�{��0�-�'��'�h�&M��ꩀ�� o�b\�Ó���ܒB�Č/-P$3fF�.R3��+TEB��M���?����ui���?����?���ϿâD
N"� X��_��T�`ɋ���'�h�ϓn�eP���$��£B�Wr�=٣��rx�pƊT4C���:�g
6�Q�H_���|2�A�)�3����V�H��N�J�(@�B�G�!�d��p{�,:�<�0��܀W�����HO>��a�^���l�l�c�XJ�x��Nʟ��I������u'�'�R8���y� �"�Q��g��z�
 t��
mk!��A1���̕��潐&_0,��BO���G�͔����b׀t��@@׋�?I �)�O���7�A�~Kj�+�\4�����"OD9�gL�[����#��Xg��A�D�W�Rp���i���'٠Y��@�4�!y�����y���'�"�a���'��XLR�|�d^'�؝��hجK:�b�9�p<Y��z�+�"a[q8�T��E�2�z\J��'�2��7W�'�p�9!���(��y E��O7$���'j��a!$��<�ҧ$LO$���'�7��56 �)�.�@4dXu�K�	�qO��hV�~Ө��O�ʧ10�T���b�~ �%�;w��;�#��W�Yz���?�G%��?�y*��	6J�p�dc���P�o>��'�܌k���	�<���6�ѶG����4O�n�<=�	-��S��+
.az�c¦"ތ�V�TCP���ȓb�4O�Q�P��#��܄���HO�Y� �S�$"q�ք˺}�@��զY���`�	U-N��$���l�	ϟ`�iލ�` �B�����R+�n����h̓8��5��/!��c6��#(Jy6�9
� b2N,<O��*��${��x����pٶ�h��Cn�	rپ���|iŚ	M֡CC�#�����"�yR�خ|;�k��������nۦ����V����@`�&�^
>�Q�'˺0�@�%�C�TSvYw��O.��O���ĺ����?A�O~���&��H��^�4�C�%��xR L�? ���s�ٽ�(!�#���� ���s؞}�h�AE��DL���%����F؟���]�n��!�a��f38�q�f"D���voN5g��"i�pt�в�� ����'8�u���c�~���O�� �"��.�,5r�璺z�xH���Or�D�t8���O�S.��!�CE�jѲ���KYn�ӆJ�{��4b�̈́���b�e�'�0�����u
x�@͆5C�Pqӡ�8ZhVdK�ʕVt��	^�-Fџ�y���On\%�����kx����4[������-D�4���.2�sa'����9��z�49x0�$&�]�\i���\�<Iq	�� ���'�"^>ݘ�@ޟ�9a�D�W���'��=܍R�Vڟ�I�#ʜ��h�S��O�i
�/_p񸍘�*r�n�Cp�>!�CC���O%6��b�R_V�����,�H���i�O�-$��?�	D�W�? �|�cP'� ���<D�<�䎚�4[��rfe؟j��@�WK<O�YFz���5EV<���e���|�`�BR�6��O���OhE	�,D�����OX���O�)=`u�
 �a��В�@�	�
c��Qc,<O��+���R����C�ĹD��� �y"�F=e��I�R�E���2��5q81O�2����9W�k�Ea�9s�	r!˓�!�ӴJ��DR��@�zXDu��!��	>�HO>Ҭ�4ej���
L)\��q)�)пa��j��Ο��Iڟ��� �u�'��0��8�C��n���4.R<8���fX!�[�:��(�Ahҥ$1�kL?f�J���O�8���JuP���ƀ e��
!�,%�O��2����]��ƞ?���A�"O^�`B� Q���� J
8�PxB���G�d�Dm:�i#��'-5hw͎/�8�htn�!P�j��'��*�@���'o�)F�Ҟ|����e�@�;j�� ���p<�e��^�ja$����+��K���t⩅�I3Rv��d[C�`T0!�ҭ޴3mP)J �*rB�	�d��b���{
�BG�LS8B��'�MC����h��mR<09��@�F̓lsF%ʒ�ii��'�哘f],���%��$i#�H�x��2L�W�`�Iʟ��П0�<������S$6���Q�P�6�ic�@���g���Gx�����]�f�K�>� �P&�7��	�}@���J�)��6@�kG
���qF���SZ
C�	 :R�	a�H# 2�`R��� ����L�'��) ��F�;���Sc�X�����{ӆ��O��$N�	N�i��B�O���O��4���S��C-ns@���Ԇ(���B�-�	�F��d�q�����ˉ�XJ�ģCM)3`qOlm@��'g��J7A]����5r�����rI��O|��R�����5=^��#"��c )�c�$�:��O��k�L
�T���J�8E0�'��"=E�4�~f��)'(ʵ�e��2�P����dq"�'u��'`�֝ޟ`�I�|zG�^�h1��Ҕ$^�6J�qW�H�3����K^j��AE�"ڊ���
�&@iT C��Mc<�EL5M�:m�r��h3>���mN:
��D��b��d���2�%˂���4-,D�(@����rq�d��;U��� **�	���'b���d�j�����Oh�V(N�}l��@�F�S���	�F�O��$�[�z��Od�J *��'�dS�:��a���*k�@��4��#
Q�xrcؠ��'|2�+�/���\Ls�O$��ő�zr8�ɜ��Bf��d*)	-V�Y�mZ�+D�5�ȓyޠPW���r��t邈	��(���{��v+�:}�w
=:�R}��g���'QА;�Gj�x�d�O(˧"����nY;�Kz�y�o�E� �2���?!E���?Y�y*��� �ԝ�q�[�X0����)Ƃ8���'��Ը����մC���ኺO��`qA �RI�v'�@��s�S�'C��q�|S6X�"���&\��0b��f��2@� �F�
�ZR�Ņ�Ɉ�hOT���cW
$^� )�ܙ��be�h�d�O���K�8>�CU��O\�$�O��4�V��E��S�%�W3I1\T�DO%扢~]����	bR|��ˊ;T~����@:$6qO@�%��� ByI�o�{�����fx���b��W�ɪdx����|bg]?:�1$H'5H�M;�M:�yBH�(E���A!�(<��˒����\I�����)T�Y*^!@ܲ���;�@���&q���"�O����O����S��?)�O���
�'/����,�PRv�hnO��xb�˼oD|:��4p+�%��dtT@��'L|"�ک\���
��A�'^�y3Qo�!�?���'��1[�.�nm���m��	 ��'� ��o�4������ܛ�y2�<�	?��$0�4�?����5�e��'3���9��|��?	!�ǻ�?A���쒦�?aM>��� 2S�����7}1��� �P8�3S�*���(8��hP��h�Ą�$1�t���4��|��6v���X�9-�Y!уC-�PybgN�N�*0�E�Z�l�h��D<���i3j���/�0����ˎTp��	�y�C!Xz�7��O��$�|��B�?���+F���p��Q:	��p�(���?a�O��)ʣ�;����pȥ�Km�p�.��5#��0}RE�,hZ��=��b*̺I���eK��EH��n�W��8_��'M�O��OAzh�G��$T�݃�#�&U*��yB�':�y2����⌚�E�V� �c�o���0<y��Ɉ%TT��P�P2$0Y�N�%��P�O���O.��t�Ī'��d�OX���O�n���	�!�]�x��d��0���j9+@���zĐpk B&�3�$�'�"�G/`/��j�lƕ5��#p�_$CƌM�	>���8���|"CbCN��WK�}�����<Vr��4��#�O��OB�t���׌��-�&�@!�6$b5�2D�xh��Ь$>i:-٫�ӳB0?)��&��d�<-@e8�X�/`���7怷'>�C�ɇJ}�1��\�?��H�O '$B�ɂO-6dq����H���^?o~�C�I�Cmj�ȁ�{�~�zfNY�eКC��b�@���_�Xp�(���S�u$dC�Ɇ/�r͡���8^f�b�	ānȄB�I�<p�;祄%d{���6Q-rB�!,��B��Q;=}"J�E/�>B�I�f��} %P<C7lW���|��v�l ��اy�Lk6Gf*�]�ȓ_�,��R�W� }8����c
J��ȓY��A��D����;�N�758HH�ȓX.4�r�  ]V>HZ�$´yK�X�ȓM�
�����'dd��"�*^�����%b��Y�o�P�����g�6Y�ȓJXr�Rc;%~��Ϙv�чȓp��z�b&6�n!��MAR�r��_���pc���dK��R1N^�I�f=�ȓvZ�Y۲�УkC��H�Ň�{i��ȓY��-he���tYp$'�@�!�ȓX�,e�����{ɴY�S,։<��ȓB� �3qD�K[&��� ����ȓqL�$��Y0_a|a�s�m$1�ȓ4��[����R	���w�Z)���5��̀Y�$=@2���~���ȓ�2�Y+�<���C�Ц���Rz8�蒅I�Z����b�Ev��ȓ%gPU�ګz$ A�`(7ॄ�4�XP�������L�Y���ȓHG��{�� �>c�M
�i�(����`g�-XZx�"�B"NQ�ȓ3�a��Ń�G�P`J�^�XBZ1��2��t�l�Q۲m;b/AM�ȓ�B	�7�B�E���+5�N&O����lWr�j@��U�^�`��#�^a��+�(r�%�!g���(Q,>6Y��Ң�W��pb̫REB�a��z��?�EIS�D� �cT�4�`�cs�DS�<1хZ.�t@x� #K�r9y�ň0Sݨ� D�W�20�0"��ی	�'�hO� @%zC�q8
q�a��>b��8r�'>�Ar&бk ��UA� S���'�W�^� ��u��#x�t0��?B�}bi�3 ��Uc%��)�x	�e���OlpB��'�\���BW�r��æ|ʓ�R�{<M�J�"���v�<�!�Ƶz�z��C�	8C�qr$`=X�h]�c���J�ԝ�7��VЁ��9#ף�7Gr8	s����HἱC�"Ot���A����(�(� fOp pCE׺y`t� K�& �(`� w���1ړ��$r m�+B��4b��(:�݆�ɆQ�td����)���G'R�2Cf܎.%B���ϰN0�sp*�Nx���&͏6H��"�L�4�v����0?6x�E�[�)��M��j�T�)��Y��U���eƈ�<�Ҙ�@"Od�h�'�94����87`.`��FƩV����� z�H�q�&l�d�}λ�T]c����
�r� 2� ����ȓF8@C%䟃
0�Z�'�0ST��e�T��8�D	B�A�B4MU�|B���ߴdP�A����k����lT�PHa|bƟ<&#r�@�gJh�lq���0 \�1C,�(�$����Z��O4A�D,QG��O�O�dDsm^�~� ]+�b
���!a��@d&Ȋ"�ʜH}� �RL�4L�
ʧC�@���DO�8��Y�8�d�~Ne���>���0�gyeZT�4�q$[S�`H��F1:Ц�B!�QYǲ�2���T�n����'(@P�vA���41v�C"B��{V@Q�rI	8G.�M�i��p=IE@X�f�Pe�b�h y����<i�E�i������^i|�S�d"K=�F
BB"��$]� ∕�P�^	6=��QH2�OJ��U��|�3�Q��^bF�M�|�Z��H���-Od��5cQ�W� 48\wy^`��)��.���8�Էu��tJ�";a#�d`#dT�J,[���/kq�F9ˣ�.IҾ`+Q$�?،�7i��|:`�Ѡ���?����0���'A�FA��4��°�O-߄`����/��)I��OHs���S��M;��Q�8XCŅҀz��e#��F,��A���,�q@IonU�2�^8YEzB��'_b4xJ#C��6N2��6B��y"N��t��8hg,B:,��}�'�R�䬍�H)0��qE?^|��qeX�MFf�`AK�*��`�#�Q�^׆T�`lV)V4Q� ����{���.H��pz�gò11�$�'��\_�`c�7�6-V"r�!����<l�FP��X��������m޸~ ��k�`�&�F�C�F
�O�I��˜1} U�ӈѾ��8����tD�_�6�"!nD�z-RH�D��V�d��CgZv*Fu��*��l�@)wLm�,D@	+�wG���)y��m[�N�(vt�qr�,)2��CBɖ��E�fO�=�?E�\c�$��J��D[��6�Z�9Q�֎<�0�pB�Q�EPi����SUh�ʇS.gtQ���À,&9�a�vmU�Di;0�U
y�H�lZ(W�,`&B�-�&��'f9rA�tiu��i:2�]�?i��ϸ ��clS�yC>l�U� J��)���~F�x2aF@����C(F�����)�@<��	f��9�j��l�V�m(����ch�����X"�ʼ?۴a	ݮ�`���/��P��7�&&-����5Y,��y�폝A�T�(�a�0��j��^�L�['�x�<�AE��������5b8�E�
pl���8 �A��[7�!���Wh�=$�ա����<A5�9��A��I=���X3�
P�?Q ��
&�@�K�I�F���+0�ܮ�.0a�	L�TX��k"�^�B���X��3F��Dy��0$ v�0a��Q�j����1�Ah�+S�lQ�G	
��`��ޙsrc��_��QsB�?��T:R8�t��ƆJN:]���*N�!��]��x�m�4H���2	�x��jҥ*�j!��Ӿ'��)���<.&\�ƫ"���w� �I1�0�uڟ\it⏔rNL���:�l\���d^��Vƙ)a� ��W���K�>�
���qB0��B�.��&c�F�!a,��y��Q�)2�l�b`�1��O��m�fhc�A��ֈi�C.�/�t�2w�a�@�c���{d����B�3wA� w�"|�#鈏)'n��f�D�6�z="s��<���p�^Oy��R��I9�oҹ�(O� �Aɕ)���fBe�P0F�^��]���O�)��� ������)��PL����%�'��v׎��y���dʄ�v��O0H� ��uI� �T>L�my�����H�''�`0�dۋet��n��5�H�$�O��W}"�C�fXrA
h��!H��O���d �,�"IC��?^��bS6O.��ŋԌ9B-�����"��«<H̚',���?��HrO.��M>%>ͱ��|���K�h؀F1� ��欟���O�C5���-w��Y�wir�$�O�I�,��K��6k�z��2$V1�iR�J_���qG�>�[[�l�0)�9&��i����JB��ƶs�.MHc�Y�"|�1�L�)��y�%ć O4B��6tvf��J���M�虆�5�
�.ł����6V��!���۫&���V�O��x1��v^�f�>%>��Ƃ����%<Z����)1�4:*؀��I��hФJ;p�2��@lW��Νfb�2Ґ�Bٌw���OXIAU'���̩ �-�Oox�խ��k���0���8�VL��!¶z�F�D�Rg�(yW ��e��qڬ�F�s��Aw���� �4 b��q(O�9N���t�[w��	���@�bj|�AF���}`� ;�K˷\�N��$�����s��}��D-"�|���O��P�~~QR �T N����C�K���s�E0L��)� �,[a��,vp�i��ĩ��bْU6��@%a�`����*$���P�fPHi��ԉ���Z��6a��0pМ����)G4����'l|Y��ߗI�6���F�M><�0$��u�ɲ�n�8ct1�T�ґK2X���.�&�I��>=�O2,�ٴ�(yȝkT�1�4�;rG41o#>a*�3*|3�+��7��	�"^?��`T�$�YgE��IјQ�Sj�&� EI��1�D(ؔ��?���]��PP� �$,W>���EO�4e����ïNQ������IW.�1X�>��-��9OpA�t�B�X�Lٸ�!��.a,y��6 ��v�̍/�9��΃%E��l�|ȼ�A�O�up�C�� ;+
y�K9Ty�Q��D��%8@��O�1��) �"?#��;U��{B��g <h#K<wwP؅���{��x�,�'E3ŉ��^-:�;��6��7�	f�(�RS�T�r؁�+�8K6�d�/1=Z˧j<�*F�ތQ�Ũw�]��8Y)�G�Kq�ؙ5�Xu�	��ke������ �w��J������95XP}��F2x��ᴊ �+���%b��=&�8� �Rf�:/Z��`� �e��dx��y��Z)� YR�^�W pAiV�~ΓH'��V�ͮqV
-u-��l��Y�M0f-؝;�ѠU�R����uXT���DX�M���U\^�9��͎YH��B��
����<��E\�m��D%R�N�{ ���?��,�V��҄�L�(x���>Nra~�Cy`�ÈO�40��3�M"I��ڢE��M���8���ALӤɁ���?��c.N��$��M�L��N��O)���O�0A�,��@���3�!�:{��h�
�#f��D��i��)�.Ѭo
�U�F�Gba2$�
�f�&�O�j<��Q�$$Gʸ�+�&��/��u�?�H� r$���傗Q����	�<%O+�.yc��a���@�`?њ's-P�I<D�@:��w����g�X������W� �0�)[=ƈ4��	=Y�ZA���˭FԲ,�u��g��БQ�zL����y�.?]�Ja�C�ʯ\������.1�:u�����l�*��̜R��������t�Af�?�6ذgB4�����Tۦmg/�$_~�`�n͞
�(G��Rl�e�O����!���v��M[ga�|yh�B%!鞤�g�؆��O� ��]+�K�,��?����R)�Ȏ�A���b4Y�� A'�&��ɐ��3M%�`�un�
|R)����LI���б�Yv!�e�8S�ܽ�vd.�Dێ1&ĸyC�ؼ�?�'�^�~���9nO��1防Y���[�* .8+���"&�uJ�q��!��+AP�� c��-a�(���9C8n(�g�~����^q�����t×�~���ϝ?�����(��÷w��yô.�R���2 O�e�.M�T
,�x���.%�W��æ��B�P'�|�%L�?P�Z8:X��I�T/��L�=TsJx$�M�>�� @q眡r����uΌ�{� ����ս3�L1�K�s���	�a�P�p!*�1H�}����Z��a��K
S�9Pd��Q�E�4J�Ār!"�!q��\�?�ѬĕpZu�!Ks�<�2��l}Ң�.� �y��>	3�'��d�o����Q��)*F���- ��9թ��22�"��&�HH���̽��=�S#�~��-�@D9����!�Oo~�'�O�扝�z%�T��a���'^�4T���O�0� ML�"k���U-��L�:p��.�2�c���}���1�Z'X�!ҕ��Ya�6��'�Vy��+ 2�|{�+M�(@�OT��s匌p�p��ڊ>A��A�${��x�-���(O�X)�ʪK�>@��I���9ObptυN��2M��)F�|H�+�C�L8��a�n�����υp�brpǕ1
��+��=|S"lAPȗU&�`"g��2�Z��3-�6D|�Um���3�ۆ[���r�E����k4�O�1m\8Ґ���F(�
ڿk��YWΕ��=9��̝U�Jɒ-W� 	H�搱�?Y��p��#g�@��3BNdѢD�fj&��' 8�=�3,@�Xg8%{QL_)�����ɫ"z�I#�� \u���@N�r���3c��<�����s��I�&á:vv����Z�Q����+_0��=���j�U�r��;�x�te�?"6N���D��T�v��9{Jx�H?���.Wb�갠�*�)��-9�q��%Ǭ
����ۓfC����� �n�b�4�*�I�~F��7 S������:}����$�=^�H�#g�,�̗)�l�A�<(;,0CT ,h�\نf۴[�N��ߓk����u�-��$�a��9$\��>!r)S���(����""��@��1y��+^W��  �� b���h����A2�y��F5:T�!BG�.дc��ؿJXlu�H:f��Ͳ� L���Wz�q��T̻��$kRcRp
��/?40������#�@�`��l�-qL?t0��@$�$lB��r����CW�l����U,+x.���A�@���9lOr�'��<,u,�e�I8b�T�^<Zh�3J��Z��\c��2] ЪA����=ْiI�u���&�(8uڶ�Bp����d[�e}b��Ro��������2G�}�tDi"��h�l�<u�Q	�:&�½$pPH�W���@�%B@�Kw��C%�NU}���u�q�Cek��9)U������%'D��G��7:�x��r� �k���0T�$��K��\��ب ������,y蒩ncV���G���A�:D�����&��0BQ�f�$	�gH5D�ĠB��a�j$0��-ko�Z6�2D�� ��&$�.���wA����$�S"O���'h�=L�R�B���r]q�"O,�9���9},�
Ŭ�/d� �3�"O����  u�5�T%�	�0�a"O>ܛD��#�I8R�ƇL�� z "O�b�&ϗ b� �l�>d��!g"O���G�!��H
'%����v"O�͒�K͂6�ع ��c����"Op��S�[?(��yŮ
<u�tm�"O�02�"Tc-�upNH,R6>\�#"O�D	U�;&۔Dx�64 !r"O�����<b�h�Z�+݂z�3!"O6J�FD���)K�'���1"O\�RH�-
R��!��R�lp#D"O�ep�.�;��U����Qy��I"O�4"�� �n8��LN ��f"O���JFlX ��M�m�@"O`8���Р{R�З��TrP�c"O|)�D3x�����/�1R���I"OP�kL^�O1�Q���iЀ 3�"O��PH��+�h��B�˛U��0�"O�LC���w�
uZ�N��A�P"O�!1�� ,�" �i��|J'"OX��`��c^x�2B�p�^m��"ONX�a�7!ܥP"����|���"O,H�%CC����Q0�D��"O�80�!\2��<�@ឃd��a��"O�����HP�&A�9i���
�"O�9㠦���])�J+{j@���"O2�!�
A!P��x����%?.���Q"Ony��V�(m�t�11>���"O��B��u1:-�l� F4�1�"O��Y�K�?E=T�b�.�+�x�"OnP�ёv�4����eBf�:4"Ol�zB�L44�H���N��:ޑ��"O�I�EbI�	u ��9'�鐀"O|	n�:'�Q����>�p�%E)D�0����Jh0`��:x�^��M%D�)#��:�|��f9(M���� D���h�� Q~)C&`�� J`\�`F>D�x8�f�4~�Ja@��a� l�v=D��2�2f�ޡY�KJ�F�f�?D��ˆ�,%�n��ELX��u�<D���Q�߿WV|�g�H���`��N:D�����'~�%Ҥf�Сi�j;D�X Qk��go�ՠ���|\��.D��Y`�Z�����oֽx8���.D�Dc��q�s� و6��9�$/D�j��t(:LqckU /�䁋�-D��ʄk3B�l�E�0I[��I�D-D�$���N�=?pi!���O`���`�+D���S΍h'NxRCM�\��`c4i)D�\�F�C �D��1kG X�ۓ/4D������k�jX��h�B�681C�>D�l��� Ob��p�aT�n���	�g<D�Du�� zʑ����;4�EҠ�:D�L���Z<M��3� ��6$�a0�7D�(8Ϟ�1� L��k�3C	���4D�bTJY�j4D���׮�e0��-D�0	%$t�H�"	�[�`�qN/D�`a$'J6i�����nTH�B��Q�.D�p!�K���Ч!Tj���;cJ/D��
�%1Ip���Ї^+q�����+D��g�Q�7��=iD��:?%�tY�>D�� �ࢀ�����w�pL���#"O�Qb���W�&QR��A9�MhG"O6F	��!�$`ّALr��"O�)�֍�mY��x�.J�O�)�A"O.�`G@n��N
  �Rt��"O�=����8[p�#�G�	F�(T�e"O��#�N'{Md�a��x+�Xf�<�D�ζt�tq�h��#��)�~�<�dťl?��s���/�v�wE�x�<��*�G�b`Ђʄ|� TQ���H�<C��H�#�'�#��h�O�<�h���r�}�ix��`�<!�k@&	�p-kwcO�UZ]�ukB�<Q��=̨@P׊ߝL1f���jYC8��Fz�!U�L#��ش��̪��Hf!���+߬,p����H�2��W��'aL����HO�>Q`ca�>2-:��WED�\�ti'D���gQ�R�牏'7HP��%�!�OL���[�Z��VC�*
B�'_��,�v����'�����\�1!��H_ڨt�.����A�\ !�DB?O||E�"�1��9���p�!�d��>�P�1����E����%�!�DV?���0$ȫ`������!���'�Dip5��^�y��τ'�!�DQ�n��q�@�=�4YP�ńV�!��ۇ�.(J#H՝���hK�!���6QW���!Z�Y��,р-0�!�ą"�tLZ��J��kB�Q�!��H����72�lTAL2H�!�A�'et�����b��H�e�ư-���5�O�4s��U}&�4�q�ӏ:�4 ��'k�Ip}�A�Ԭڬ��I׬�.eF&B�Ɉ(��h�&�kڬ��hJr��C��~i�P��X�R�n�`P/�9��B��/x�1��(i�d�)5N_���B�I*�����Ia�R��TA9<�B��;<1�(���[Y:@��Ճ�f�~B�I.]ь��B��7n6A*���)LO6��$V�M�d˦� ��Pj�ȕ�&��~b��<�VČ8 ��1˗�ЬUb�Q��C�<Q��$t�4�`�>S?f�I�#�y�'ɑ?%�f(Z�j�l���B q�-��:D���Xd�F�PȂ�Aa�z�H7�IS���O��E2ᇄ:��q�ڊ��yq�'p|��@E��x3��Q�u�d�}r�'��a��Pa�*e$�q�|���~����3A���B�I5xrfNّ�y��(���t&W	I�6��)ŷ�0<y��$�1�:T���S��Q���DD�O���D�O��	��_m"RR�X�/�B��C��
<!��9M�8Y1���+~���jA"
&3��&�)����	Ɵ)_�@h��v3��V�M����|}��-�g}��:5d8 ��@V�"��X�y
;ܮ���a<4�$�zq�;�y�ᙼF\Y�G�-�X�R"N\:�yn9}>�:�J@$L}�� �(O��' x��'iM�g���-��!�l�Fz��~�`.�i�HC�DA�t #�⦩F{���i#"L�O[/��KeGȃ'{���'53�h�pŊ���Ϙ�]]@�'tޭ &�!4��I��~��ъ
�'O�Q+���"{r��Y��;!N�D�<�S)��&�d�k�	]
P�D��
j�'�ў�g�? �Y���=������֬M�
es��'��'`��b�c�
h|-c����v�5�'Q�͹qlD:gFb�!�'׆G�	�'䊵2g�W��� �w!73���'�����#�Pɧh���)p�'�8XH[�%�εK��Ý$d}��'}���l	�q]�8r�*��T:�'r�z�d:�Ӵ�>�4q	�'�^T�w�I%Oc2(� ���=��	�'C��H��"�fP$
/8�OX74�S�Oz�%�*ĵk�[o �!�j��'>`�:�mA%]�NA"��E�!��'C��r�F"Fp��NN�?�Hq��'k�h����x�l@`�S�&O^�Y�'��́�Γl3��Y*�#zhP�'�r���&�b�NM��/���c�'�R�S�(+f���DaS�e͜QQ�'�����\�6rl8[���8^C �3
�'t����cɺ\*dE�lK2��x��7�S����7H�Lt��[/Un�AJV��y, �l'$��&���֬ѷ�Y��I��p>����Ɣ�c-�V�l�s�͘E����'����vb �c�CLTE�m�b!��kf�<��"�W�`�����k�!�D}�5�3
�$K���d�[/(�!��A����MڄO��Y��ře����>!r�Ua�����ax����-�f\��CԓWq!�ď15(Ќ#!bY&E.�AB�S�Cq�d1�O����D8 jA[��B=
�²3O��=E�4�T�b�`���"�D����$ΐ/�y��ޑ4+�8��	Z+���3��L��y��%Eg|�" �Q3�h�d�ú�y�� \b��)��E5V������;�y�l�/\|�p,�/\�\�K�焛�yҠ�"O���'@�>�~e��f���y�B�:G���rAγ4?&��塖5�yB��$ ��	�Ԃ��/`r|(�B\�y�#>3]�@yfEB4�1k7��y�+g�`��ၦs��Zr!�;�yr���J\�TrT>�qQ�I��y2a�
'~Lb0$W�hP �	Ӳ�y	T6m	!�E�^�|	3�'ĸ�y�g��@��i�n�^s��ܰ�yr���w\��E���Tu��J��yZ�&�e!V	��_�ջ�����y��+Y��$pf��'80jC@ѿ�yB�̕Z`�CP�G� �0�8"���y�?nu�6e�s�=!���y2�
"^@x���f(9I����F���y�7a0�jA�)�^U�҉��yBoBxz�����:o}�xQ!��yB�-O �x�Y2Ŋ�х��!�y���x�8G� )Ŗ���I����7�O�=9�f��C��Z��17���Z��A�����Kp�;C�8{��Z��̳=38C�	7-�D�RfI����*��ly�C�:RN��:�%�$$(�@W�P8 ��C䉴8b�q�a��J
��NM��7�,�S��M�A�\+�4�I��>4��( ��v�<Q���@E���EC�.5��[5OYu~R�'H�ucC
�6 �,�ͳD4`��'���YF� 4KZa	�+>��`�'I�/t�:%ƉY��iįJ�y��+�0@�j
7S3>���\��y
� ^H��ꋠ[t��
�Vu$@V"O����U�k��K�js�-��"OFx`��U��i g��yb�4S�"O��A�U�P��*C*lJ*a��"O�  !DJ#xT)�O�?qS`��"O>�
��V#�X�#/^f5���$"O�Y���Ʀ5gd]�c��5P�C"O�]��#\�,
�ذ`�=. m	�"O��!�I'M���QF ,,��S"O|��G�L�� B+�:Eʔ"O��3����|�1+[���'"O����);;Q�-j�`�x_�HY�"O�U(��ʓu�4(�e@��O���"O����ԉ��X���3fƺ�)p"OEq�V6w���q)S��hm"O��D�b<��"j�w���g"Oni:��c���4��qo���"O�ep���%��l[e�Z#"hY�"OV}*qG	�X�WʪE��`6"O�xX�Örͬܲ�̃�^�$�"2"On�Jg$^�|F:4�g�P�����"O���k��b�BY�A]�0*�0˃"O���v,�� U��*gg�)}�$�je"O����b���0�T9=։ʷ"O䨡���4�ƨ�w��?A� ��A"O4І�_D���`�ȷ"v�E�a"O�a��B�\�� ��Ā
Pd��C�"O"m���50��r��4O,,�v"O2� �!P�t��R�[I��PD"O�A�'$ܴ�킡���j�Nhɐ"O�� @�$\L��#j���V"O�,��$�:�l]Rb�	44��b�"Oޤ�#�ӓnA���ƀDO��a"O}B�L�)��Ի��Щa����f"O*1�8��%cSh�/���d"Oh٣c�;a3d��sfܣ|܄�@�"O��b�]�I﮴�T�;��`""ODC��5fح��˻WNR�KD"O����%N�P���!�m��Rh�I"O���<f��
`L?6,*�"O�Huo��x`@�#숤^��(�"O���dOπO��X����b�"O`�Z�e�>vv�)·�M�Fq�5"p"Ob�ɱ�`����ViqT��(p"O@�x�*�6m��Sꃴa_d"O���
;��`;�G�+q�!�"O"<���	-�6=+2��;S� ("O�S`aC�1��kco��y�ԅ�A"O���d&��R��LzQ�JCz<�"O=A�̆����M�	?�!��"O�x� �[�#�\	��YM�{�"O��>/�=���4.����"OdQ���@�p����8��S�"O�)ȧ�}��p����9i�"O�� �S�O�ʉ0䐻w�6�"ON��v&K9EL��5��v�$у�"Ot���0���q ��O�.|�"OL�9�!��n(&�R�y�9�"On)S��@�fL�0����?Zp�"O�=Ʌlئ*�`;���3R�J��W"O92��`E� MF��Ȃ"O8��Ge��s���AŮ�,U���"O�]���R-k�z<�����,�͂�"O��
��V�B�H�@]�,L*�F"O� ڡ� ��3�y#��
C±;B"O��ji��8���N��/I"Oh��d���W��13.�P��;T"O������,nvYR���tb�q�"O���%rL�R`�Ć�v�"OT熍�5��ꆧ�<q8�)�v"O
Т� �$�59կ�üyp "O���%ބ!�Ĥ+�m�W>�S�"OTi�7JA�V�=:���5vj�"�"O�q��AP�(��г$k�'�xq"O*pH̶s���Ȑi��+ܢ-�"O��"�Z�Cz�`�U�DdhH��"O����y�(qRM�!gF !��"OV"`�.<�hU��JQ�4DZ��"O.�{S�I�<,�jު*H���"O���qO�rC��kp/�=&�e��"OX�7I�2Y�*F��Sd�ġH�!��@(r��)M=&`z����!��´6l#�,��	��M�GX��!�$V��ڤ�B��To��#bƄ%�!�D֡K���C�]� �p�"��ʠ+�!�L�i�,Z"!�*İ�E%� �!�$_;>�04�WHQ�
��1"�DԺpk!�̋ted-)�(�;v��q�L�O�!���4\�Au�X��X��@�7gP!�DQ�"`��x��@�i{b/��SE!��O�
�Fɀ���z��dR5��?k
!��\������!uy B�M��!�AzQ�%���
{u�ݣm�!��>
�ĤY�O�(+rr{h7�!�DV'90�+��$8f�)밧�+#g!�D�29�����K�=Q�Q�Y�Q!���3f�i�ꛀ-3b�� ��<!�D��dH0P���>��mcG�ՔM!�R0h�����G��ġ��M>q�!�$��(G�� U蕇~�
�t��	Y�!�dT�P	vpP ��h�Z��&��U�!�^x~~ ��S�M�b���G2)�!�h��HIC�\)�<ؐ�A��!�$��
����K�)e
���4�@h!�d3#I���@�Ӗ Ni
.�./d!�$�Jyj񡵉Q�TH�)En� M`!�!�h�pR���Y� y��n�/�!�ēv��e�T�J�`�B#l��&�!�D¯}R�M��
�Z��d��G�}}!�$� \����^�RpP\C��]�}�!�Ğ?/:� �N!1�If��2nW!�ɯ� ����ϔ:�@���Œ[M!�$.W��<��?/�jt1uhɑEC!�$Β0�b�� ,��t��D%Z�~A!�d�%����/N�4C���"^
!�$�nTxX���/�$Р�.Z)�!�$��`ʨl���I%���D�?�!�^/#�2�AG�B^�4M]�!�$��q 4��N۷��c���!�͎r{ y�r�D�h�b��[�;!�D�I���������)5��	C(!�Q6=Z| �#޸?̦�Kjݢh�!򤗈j�P �Pq�`��c�!�d�6ʒӧI�9p]K"�H�!������%�R�p���
1�!�4eQ����N��="�AZ��!�̊99F�D@�?�P��D���!���)^P�rEМyp�Z�ĵ�!�� Rt��@F����c�FB�05�8�"O�Ĺ�%T�5ٞ�#0��3�xpr�"O8�����@�GFT"]j��rd"O�� ř�!���f�Y*lPf��"O���c盚?���q5��'SA(�xd"O��!�g�i����c�=/t<��"O^�C�E�<��_�kg��!�Ҍa���S�M�f�[g��<r!�d��Is���F͋"fQ�T�KY!�$E0l�����o�>H�v�M-�!�$/񶌻4�\�g�<i���!���[,4��1�D�4p���A��!�/@A�"I8}�n���B��!�dI9x4�i���*�`�0��Ԩ�!�d��c���`roE3���΄��!��(|�u1d�
����-��k�!�D�V(�y�A�n����"dF̆�<I��x��?���ԫ�5ɒ<�ȓWB����=�Xh`��B�U�di�ȓnI\�7H�e ڀ����h���ȓgk�pA�8N��H�X��Єȓ*�@!ЅR*��E`���MШ�ȓD�� I���2G7p\�e�=������ 4��&X
f�[�	�L��͆ȓ(�~����m��dӦ��&��}���`X�����Rk�(��d��%�橩uɈsL-�3e��\�r�ȓ	?�q�oC:t�2P�6 ԝ�(-��1 ���JW!pD@����_^�͇��U�d �[�`r�FB�Dć�7&@j�*[mzAr�&�H m�ȓ~`�U�$N��PV��9!�h���u���Dl�9��i0���-w� \��\ѠIA�*��CL��R��4<�\܄ȓA�)8��.T@�ꡆ4 ~vh�ȓ��Т�蜡k���cCM�~��d�ȓy���`j�
o.��6��$����CLV��W� -�.��#��CE�,��B��|���Zi~q��}�����6}�@�G��	�lҧ�@�y���ȓY:p�@�M� �fX1,�7�@�ȓy�� ��2#f���kÓQ�2Іȓ6��Xkg�J5���B��t�>H��jj��CKYus�͚E#�"--�ȓb�(وգ��[]�XJ��E�� �ȓ%��y3&B*2p�@7��M:��ȓhu�%9�n�D��Sg��Mz������S�� .�R8�rGH�9X���V �ĪG��>Jj�§a�78F<P����\I�H��x�8qj��V���ȓG2��Xc�d��!z�k�V ��n�4!��}vX�	@'_r@��ȓ}�>�J��֬b�@�ögL�O^����I�x��K�aK�u[���b�����{�
Ms���pc �V��@�ȓ���7h� ng|-kˏ '?0h�ȓ?/��K2��S��*7L�8M� }�����ckI�RQ�4�� �)6J�1��>�*X�!UeR��ҵ��a�����p�u��C��~`ciِ���2&R\�2*D�ڮ+�o�O~�ȓ<Z\���d��%E&�j�HXEW�̇�.t TJ Ɛ?sX��SH�f%L��ȓ~�¼Ȳ�ȠXM�=�WBT��S�? ��aq�ٞ#N�`���2g��c�"O�	�v$��HF:�{���I��	��"O�����[���B,p��I�"Ov�s�ɱf�2�Q0N@�(�"O=(g�׶[Ȃ qB��&�ps"O~ ����+[��"��۾Sd �8`"O~-���ؾv���!��� k��:1"O X�M�HG`�Ҡ���m�E³"O��s0�Z�S��@O9/ ��c�"O��%�Z��}�S��|�T:�"OZ�q��&:�� $`�9W�@�9 "O�*"�S�l�\�p$/�1[� �!�"OPd��͹dm�V�A�E$:�"O�w�ʙ\-b��c��$z���S"O��,��x��e\�oX�	� �#[�!�Y���<�$ᜅl��{%��H�!�:PJ�)B�$up�ٚ�M�4�!���$��2�U�\�|u�B�\��!�D
7Q��|A􄚐k���q�6[�!�)t�YB/���\���Y
!�d�'0��3#Ĵ2���'	*;�!�$X)h�H��%�,;��xD��$!�
�
�Fh��j�'b��}�@��!��ebq��[�rg��(�"^4N�!��Z��@Q	�dd>ݛ�b]=p�!��
Ӯ� @]l� �+0=!򤌶@#(eX���"C>hp[�	�D"!�I=%~Ό�s�BVZ���K�	I
!��%`�:zr��2T]P�_�+!�d�w�����D��`�`ˎ1!�2K��1i����U�N� �!�Đ�Ob��r' ��ɋ�)�=2!�$8�a0&F���&M����B!��'P��UҲ,ȭg� �9�#M.!��#od+�FA(|���G#S3�!�J<�.���ɒ(�x�0cA^�'�!�d�@'��AUL�X��{[�z|!򤋧(*-�U��++��1���.^!�dٛ9�Ii2(� )��qQĐ/ B!�d^jY`��/d���;5�\�u!�Ě�G,�Րb�O+H�"��3 !�$��Z��H�H��\�v	HիMu!�d��Ly�b,�Hh�Xx�O'&!��\�������-�Ԍ�N�!�K:#=�$�T�ׁljI��P�!��,Z����`Y'P���JdB�X!�$]�9����cǰ
(�d�O�5�!��ߔ\��Z�ÝK��]��-A(�!�D����׌o��;��L?;@!����N���
�g�u��(t��'!���*x���ch��m^%����8�!�D�`5N�3"
�6\,�`��C;�!��	t��q���fB����˿Y�!�d�dA��S`�ףD��W#K=y!�D��:�|�i�g�1&Hyt�Id!�;5���"`��Hz0�2��%T!��F1l܂@ ��F!�GF!�K�12xR�#�sGH��� I�!��361\9"(C*B1�v��ox!�d�2�>ժ��.}����(�!�DR�=ݔ����6���P#��%B�!��9N��E[I^�As��#�A�7w!�d��hv�`CǞT��12ˑ+hr!��կ]�dE�&I[$�0h�=i!�� $u��H�%D$��G٩i[^�(�"OX����D����FB�N���"O�1� ǩ%�|@&��Ab�V"O�p#���<:xY�V֢�B"O�$���)� Se	+Q1�U"OzT����-��Re��
X

�t"OF���%E��aU	�U�CW"OZ�8�ME"W��cI�H�@L�"OVX���8��U�a�ٞ\� �k0"O:dk��9q\0��([� ���z�"O��`��ҁx��h�#����j\	�"Od8i�U�;/�0��FM�{lj`� "O����h�)��8�����)���"O��T�4D|��'�����"O��ʅBЍf��(m�����"O�0c�L�+n`K7�H/%i:Q�"O~�j�m�`%��&�Z8f`$=9�"OJC![\�� ��i��a 2"O�Ð�{��=S�!FjIr"O>�ѯ� #��ӰkH?7B��*�"O �s@$Ʈz�����E�9͋p"O���G P����
�t�����"O���ًzw���S�q�p�{ "O���w�ܮv�-��+�=U�b�d"O��� 
�S��806�@�>��-�3"O*!��+�-C0!2�2QS���A"O�H�b�D,-+�Y��B"t34a�"O8�����4~*�)�������Q�!�:)� 8��-#Z&Y+�D�,w!���+e��RmF�E���*��E!���H���2 	��5���ۼT�!�d�*ox}{rFܶR�"�� ���!򄚝[=|t[�a�!*��p��Pi�!�$��N�����O�3�N�r�M�6$!�[N�|��`Ă�t���얍 !�ś16l�sh٭6��ae
C�!�D3�3��h�
h�`!�d�&�tл��&��]KQ�%Ek!�d��2.�Ccj��}�0%�Pk�:(^!�$�<* �� ��	 ��5��X�!����ꕋf�l��}k�F�!���'y�@Cc.A�$�@�R�IV��!��Ŧ��S�nIniQi��!�Ę;,��B&���&�,9�F�Z�!��=eK��qDĒ%] �8q@���!��!y?8�e���� ��5�!��T�7�D�+�mF� Q��)<�!�D�"8���l^�GN��#�JY!�$\�{B@��DΞO������K!�$�.~a�Ŭf(� �n&^S!��U�=���
d� `���H#i5!��\�"li��	`�~L�r��-!��(�����
2����&��?�!��
c�>q�R�n���Q�D�'k|!򤛔l�(P����NX�cٸ0�!�.?ށ���ۙl�.)�'%E�}�!�䇆_\�0�K�!p��9�!$�q!�Z�,|� u��� ��!�	&���Y���N�t�rr`B;{�!���/a�:Ĳ�E؃?�:D`5O�X!��&/&6�;��Q�	�>%��2xB!�+c($ b��
�D��͛�N�!��C�H�81-Z$�B�wl7�!�DӾnmI5�_��XD��}!�� *�� O�� a�>T�n��"OTq.H�[��e+A�*�����"OJ؛S��#��e �唧,� `��"O� �k��E8��h�Ǝ�d,�I�"O�k�F�(�1c�@�~H��"O<���%�/�Z���G( D���"O��@�&Z� ��x��Z�R��v"O��c�`� �0mN�p�j�1"O�MAp��&�̠���b���"O,��ue+t��s�L-
ϬXA"OTu��S�f{Q�$ߝ�Z��s"OL�0T��	;2�Ԣ��M�C�Z�!"O6�Ҩ��k�����,�!��HH�"O6�3�W�Hڔh�R铙T��a"O��Q�j2Y���U�A��z�"O��P7��#|<v�J����Yu���"O( �k�*w��Ζ=#]*3@Q���t�S�OΤi"%�'|b�T��%5�H��'�v����>+����U"4���'�l3�![�d��r��� �T�!�'�~]�d?!�a1�$�-Lb�8�'��7�-K��@2R�Z�>,��'?�ٔ �Ȣ�31�D�3�>@ �'�n��AeO� !���]1Ψ��*OF�)�)�'p}h�7Iǜ|�`y�+0~r��ȓs�X4��g�$=�|�1f�*hu>���qQKbI�8'�"���N)t���g���b��<r�t���,y�d��ȓo�.�y�m�ZJp9��#&�\���K��jg�1^�Xe9`�зD�.a��x(�/���ؐ�
F�#�@$�'ў�|�@��Li���W��5c�]L�<�BU#S���Z����%\Tp�IN`�<1�Ι*qM��Łǵ4$�3�Z�<iM :b��ꄦH�o"�Yw�Y�<���g�b�F������R�<	aQ� ��0�g*s���qS�DX�<!c�_,��T� (�%S����d[S�<��̄!n��ц���L-���4)MZ�<ig�?bA���f$
Wg�X�<��C�`�[����AJ��*B�_�<�nA)o�j�i��Nw���!
DU�<����"�&��&]Q�d2U�YJ�<1J��4�0Eј8�>AZAKH�<� 䒒l�sC�b����!
EG�<iV�ň���0	2�9ƀA�<�� � ꍢ�*_��c@��e�<�T*8�^�b���@d����ʀe�<�1��#;�@]�Db"'D�1P�j�g�<Q�k�q�0�(cZ�]�<�ҳJ\J�<�e� �V=ؖBQGd��vEH�<��D�o���0b���]�f�{�L�<1��]FRZ��#OI�BH0U�^�<As�υ%�|�"B��{c��K"�t�<��hZ���݂�G�F��x��u�<�2�Gu󬭈2)R�y����Dr�<)�k݇	S�p�/�(?zS�Sk�<��&��La�� �i%8)
�fS�<� .N9 +p�����"\(Z��R�<�v��	��#,�Wd��	K�J�<��#DgR�Z�ɿH�4ȹt&D^�<��@ؑ`� �1���m��d�^�<I�EӬ_��W�����C{a!��l����ڶ�@� c��!3_!�� ~�ҭ8��*�ʀ� �5"Of�6Äy�,����kĦP��"O44 �	8
����<1�@u("O�=���,0(V�bc"��5��m*"Od�6b�!#9te����p�z��#"Ox�J�&�� �I����6U��Z"OH8�W�?"X��D$INE>���"O�ّ�	H9U>��iA�".8�d�G"O�pR�ڹ6x�C�b��F>x��"O������:_Ƅi�ʅ:� )�"O���#�N)���dB�_1�x�"O��a!#�"�~aړ��0&����"Oީ�'�߉�Ь"��;3��4�"O�YA��E��$
QmNJ�L\��"O4���-TG���%[P���p"O�qqg�d�fF��$$�W"O��Iu�IR�|�r�Ű9���"Oµ(P��)7�|I�&��;�z��"OH��IŋE�xK�/Ƅ��F"Oj�1��t~$Ī�兪>L��"R"Ov!�AN�7�������z/�z"O�1���Y�>��p�	ǰ�I�"Oʤ���A7��5�T$Uf�M�V"O��[�cO�'��5ҀY	g�]sv"OL����.'�
�⧂]>,T���"O��CRB�w�\�Y�C-"O�ѳpo��]�&͘Tn�
^@��3"O>\K�2H��-�)F10\C�"O�I�R���e�aK!�ȵu�2"O�!ZTi	3vF�a���H�	ڒ"O.��K/j���P%� �R�Y2"Of�����A�d, ���=z��R�"O�8�F���>8��B��<b��A�*Of�Zq	ӧqkBqcG�^�x���
�'52q��}xN��U@��!P	�'��}H�=��,�dw"���',XА�YWs^�iq��0^���H�'Ȅ����2��a��ߦY!�8��'���B��Y dH��[*;�hxj�'q�}B"�H/�\\�C�"2JT��'�\zu�F T1�#H �<��'r�����"h��!S㕁 �}2�'�\��׬O9���	��� �����'Nvq�ƌԅXG�䰇���,��'x<{ ���y�i��͋t�����'�M�4��.�v�!�� �`(~���'���,l�r�m˟Q �"L�y�M�-��=q�١M��!���*6D�����R]�eIP�Ӡ\�zH��4D���˅�P�=j��Q0�rLH��0D��2��YU�H�0���Z��(�-D�$�&h� �N��4�8׸Dæ�>�D�O"��d�b~(�䢈 `�P�k���e
!�p @ݰ"-�Y��+Z<cu���"O
t�aFT��b5�L
EԌ��"O�:�*��z�b���n]0�x"O�ա������0`CS�*H�"O���/�w��3c����r"O�=)Ā�F��L#��l��8��T�܆��!"|�L�ț	�N��(�#:C�=P�2�[�ѓ+\�T* �,.yC�IM�d����-_���3OZ�(��B�I38�ҝsa��O҄�8��Ҩ|�\B�I$:�S���n("="��[�z�nC�)� ip� [�H0�a�%ɇ_"}�"Oh��V��j� ,��.�G��kg�'�!��C	O�I���ëe�r�(3  p_!�J�"��|Q`f��d0ld��Ş@D!�d"K����&ǖ/P4h�PHS&D2���҈Q8T@��-p��T
�	�y2��՚!"�l��)·DH1�y��˫\Ol`���_1V��	'c��y�gn�114�C�6����u$B�I��d�2N�m^B0���z��C�	(WXd{�F����A�R#enB�����yU)K8]�� �5�lB�ɮD��}(t唻*��Уm�"H�|B�I�^+�@"���T7�)�R�Խ{C䉡:�}��)��]��qaV��.@B�	(D�r���O"J!�&��B�?yA��Z��׷!� ��^�7�C䉉YN i.\�L�L���/5
 ��$�OZ�&mѨI�p$�!�,z������O C�I�H�"eΒ������`]6~B�6�`��N� �d%���F�y��C�	d�"�z� 	�y@�Yr���+5�C�I1)#��$m,d1Q�2f5�㟈��	K֢Ȼ�ԐK�x��N?�C�		%�0�s��V���a�ˎ.����>i�8Iz����-	��[ �M2*�L$�����f�x�B�_�z�*��F�s�C䉨76 �p��E+b3,8�f�B�-20�ʅ�ǃ2�
����@�<B�	�P;�\FN�0�\٧ L�F��C�ɖI�[0�2<���%�):E�C��9wp���&�V���%�;| �C䉊pENQ�� 5�����!*�,B�	&XpЬ��a�pʂ���.��C�	�C��e�jܚ_�x���+��rC�	 Qֹ�A��!��"� �7ge8C�ɜh�Ι�w�Nts��w��?��C䉠|OT���ڂ+���î¡-��C䉎`��
���� ��
i�C䉔!�JUbf�#M-�4�q�O�lq�C�B�0X`���!�s&�W0Ob�C��X��2�+�N�J� =x��C�	�(���ĀD>B�z�۬\�C�&���Da]>}�֘��͘q�LC�I	4H~E;���w��VMIS3C䉔�:�qe�-|�� ���75�B䉥/x4�kǄFaݾx۶�R�E��B�I)������,��D�lOJV�B�	�ys�0'�LD�(i��� B�C�I:F��(�m[;Zd@�gE�oE�C�I#jU�p�N3 �8��M�4��C�ɜTY���	D�&�u��e HC�	
�ƨyU�VB��6Ɖ: k(�=�ç]4��hD�ÌU32(@��<ӆ(F{R�',l%"w
۔=��,b��D���� �'=����"2BJBTC��� ���*�'d2��FiĸK��,w��)R	�'� %�ah�`Le#�ǲgP^)	�'Y�M�nӃ`�*�Sq�
$b?^\�	�'m��+�K[�y� H�Xb��l��'-�,	�
�s�U�e�_�T.!�'4��dk�2@Ps%��L|�'�p�Q�L�z�H���3�r�
�'��$z �"0�.�z$鏂ci���	��� �@��"�< �2}��b��n�,"OrI�Ua�B���P`6Q}��2"O
Z�@]'������{g$]
""OX��ъEz���U��&3�$|��"O�43�-NY�U��Z��"O�!�s�=.��+ċA�~�{�"O��IB�Y�,�~�鴠 �.�NxA�"OV�5�>��ZbN�� Q���"Ox�`h�8E��o
hM�a)�"O~cp��QuDȣ%O�DL�	U"Oh��q��f*�\z��`:"��C"OY�����[r�\B�#W"OH�`)G�J���p��ͣx=:L�q"O� ��cP��uOVb��]�t"OΤ9�d(C�� C�Z<��Щ�"O%��'D9��LQ;vx�Y��"O�m[É���a�F
�+k��� �	D>y��oB���KK�BM�(ˤ+ړ�0<a�匩�V%�fN{�tY1�nZO�<��;k�v�@P�Ɍ!� �6
NK�<�)\EB����#2`idhNF�<yC�ǳ'�♃P��"<r,�H2�ID�<	t��$4�Ȏ�k.jx"���<�cH�<D,�0�����5����t�<i6D�_�U�f�H�'IH-�I�<�!+3	Ȣ8x�k�:�,Y�A�j�<a�H@�E���ݞC�P�UM�<I�e�
xzq�璦8,��P�%�J�<�0Ί�QOx�5ѩ:���j�BI�<Ywo�4/X�˔��_S�� H�<)w'M[H��k%ᘸ�:�
j�<I��V<p��r�Q�b&-!Bf�d�<��oT� W�A�W1D�9�G�J�<G��*P�!Vl�=SVA���NF�<Y%oBXb����ٞH�lH��A�<)�̈]�,̡�
�pܞ�����z�<�B$�:R"<1��r
� �шUM�<i���;Z(�c
�}�ฉ���K�<Ae�ܜa����t���8�`��@�<A���]�bhz�H�x��x���<	`��p��ɂH���湰AKy�<�4ʃ�K(R%r��Mm�U�U�x�<A��KL�j-���^�wDh:���t�<�#�Q�<reZ�a	
h�l��v�h�<YƋ�.�4�EM�m9.��UNKj�<��ٹ/�B�	Ac�$<��A3��j�<)��O� dpT���$7B=��h�<y��۳[��\�S�K�9;�4yf��P�<�Ƙ3ۢ�0$�m��gn�@�<q�dD�'S��z��ǥA)pX�2�s�<ISdS2r�DB����h:���6Hy�<�����K�\���"� 	ǉBi�<qV��3�0)PaNH�@���Y�<�u�Y~@:�&Z���zw��W�<��@��9Il�[taހ$M��
�E�J�<� ��W�P��ؾ,@����B�<	�לϚ;sNZ�?��ER1�X�<�&f�7�Ę¦ϭ/(J<*��Q�<��I0x_�0�5��(J����IEP�<q�n\�cVx��`B$3.^੓�b�<�o��AJ#��?�U���_�<y#��j3h0�A%O�T��Ip�r�<���2�)K�ܽ"d}� R�<�u�[L����8)� �:F�Q�<� �a)�٩1#*q�bK0B�(�E"O��9�&�u��#Cmz ��"O�m��`B@�bXh4+]X��"Oz�B���tk.�Z�jR���j0"O��PW-23a�Vi�%s��Ax"O�H �)D�g��irfA)�qɠ_� F{��ɖ%Iq�]iQF O��YuA�Y�!�dD�,b� 0K	:�`�3o�j�!� hp[(Ӛ+�v�H�n�!��˞�α9N�p��6MH �!�D֋�~;C�C�x��r��|c!�+w
�@���6"�)fǽx�!��L�CPd������v�`d�j��!�D��A]���eb?%�J��(Ⱦ�!��]�}�*���h� v�� Pl��8�!��o�ʼ��i����4��S�!�$��iH�x	cF�m�x��� �!�$VrbL�"�P�\��C�W#c�!�S$$ZCcy|xB	d�!�dܕd�����JE�������)r8!�$��?6;F���r���#�V!�$	�2���!cU)/�^�K�gQ��!��],wV~�R �>�Ɣ�אK���(a�H ���;fHq����!&TC�	��>��&gׂF��ār��3+80C�I	�}�r�U�)����I�C�I�z�8�b�rkH;Z��آ?Q�����F)����{���9p!��r<�0�ס5�zȋ�f��e\!�$�4+ ��W��o��mY�+�!�[�i*}·�T���@7�L�n=!�D_}V ���N�G��ɵ *!�٬����F�� J��#!�F?�!��Е5D�v�͋YuΔ�t�_(v�!�$�B�p���Y
R]D֦٘��~�!���7�޹����=XT٣e�!���1-���GM�D(F�*�cC�_%!��=m!`1(�jW�:!:Ea��!q!��gH.���عx5x%��@ž`!�$M�����I�87�@�@&:K!�$_#WN�)Q��*�Z���,B'D!��L�q����5�����RD�#o=!�D�#@��!���g������68!򤒠^�mB��?Ti�������)�{�󤞆}�l�+1,���!!��}��'�a|�I�:&Z�Ykg�xܜ���y�J'�4XH��R�w|f`)�iV��y�d(&_.Yba���o� ��5Cœ�y2;~�ʀi0�	:��=I��M��y�8�hdU�0;`,1r�\��y��۠�x���5��遤���yb��2�^��Q@�<-H��E]��y�H�b��eϋB�:��w�6�y2��I��u�B�Q
l� "��+�y���0�	�)�3X��� ݩ�y�c
 T"`��JT��(�e���y2�؁����d��a4"p!���y�[��ZPr��2lMحQn���y���F�p���ŭt��h�`�$�yh
u.�re�Ge ��@��yb@ ��\����X�W�bDz@ᝰ�y��=�h'C�Esj=�PD��yBf�,q��#^�7�^{�eX��y��G���ס0��4r��׋�y
� �Q0'LV�BoPM�#�מb����w"Od0�u0]�2U�u��&p���i�"Ojq��Ɲ,4e.!���?}�I�"OH���-��fl��1hX/�ȍH0"O`�iUi�=*'���W��4T�0�Ju"Oys!I(�<5˔"E X/>�H"O��ʏ�q�i��J� ^T0�"O�^��iI"L�W���kdG�&�!�dQ=�"D�5�ŪE��-�����"OV�q�Ɔ1��чA�)P��G"O�ai`�9W�z�A p����"O^\�f�'��\9R�M�.
�3"O!#w@WI8qSE"\�&>l��"O>�{�տp\�� @( �4H"Or����3�� N^8Sv�x�"O�Y���
<ec�Q�E��t�"O�p��(��t�1eP� �4�r"O��UҭvA�������Cǰ97"O�ʠ��T����e�P�]�s"OB�J��i&-{���S���U"O��C�[�:�b�-F��B�9`"O����5SH��-�p<�Y�r"O
���Őlʆ)���BP<�:�"O4$`W/ݹH�jA,��yL�
c"O�Y�&���(J�L�T 0���
"O`�l���<SR�B�:1!�B�(5�`�A*m��̨�)&6!�d�`��`�b�rq}���a4!��E�w5�M*��MM�%!O�]{!�� C�"��«B!2��"oG�P!�d_�P�aA�*�P"t�Y$o!���-3�\{C"X����r��9|U!�d�/#���&@6k�,+�ۑ�!�O�j7y�R��;�2�;�`] v�!��G->�p����J�B@"`EȗyU!�dϵ:AK�ŝ��Fu�Sc��H<!����<�D>��A���X�!�$W [�Y� �U��Q`�Z�C�!��I=d�Ӕ%�%@>q��l��VL!��WC���W�5y�d!&�m!��O=,$M�
�D?R�"PF��R!�$W�Pg�8�@4c!B�$�q!�� �l҄���7��}�w$+!!�di�dr�̎��p����؁t!��C1o�*9��KG=�J<�ՏOw	!���t���ai�3�l��b����!�J�av����-��T�V�H#!�]9L>�� !:p$�P���T�!�d�
y �	�4#�gcL���
+!��X\���QC�
4"�+2�x!�۝b0�P.'�d�j�
1h!򤀢cC�@�D��ؚ�+�,R6�!���??Euh��V?>�t�"Kظ,�!��&VD����&�F��4�ٮ7!�d�uuL��)������cԁy�!� uP J��b�f�+�$S��!�dX�jN��G�1��h�SF!��2U��26�Y�d�E����P�!���9!y�U��C�9Nb2X�B�O!�$֟y[�5�
5hO$|c��G:!��ǪS��[���V�0�v`� !�dѷ �H0Ã�6l��Z'OH, �!��� ���2��	�i��#�� m!�$اX� �y��*���)$��r"O� �̡�K��� �KZ�I���I!"O����e��,�x��cH����yqW"O���B�37�,\�G¶�F�a�"O���'@AtE��2�g$K��Sw"O�ycV��Z8�eF+�T\I�"O�R���1��KQ�&^�|�qe"O���AC��e�hi��"V}���"OD|��F> {T5p��ޥK�ѳ!"O.����ϥ,9��sv�C�zFB��@"O�EA��L�|ņx	!�RV�"'"O�U1�Fz���V����"O"|b�X��^�	�]�!4źd"O&���$�1/���-N�j8�UJ "O���Ϩ	�Nqm�4'>�A"O�ey%��6 ܹs��6i%�Ia�"Od-ѐeS2u��x��R ��a"Or�J!�����s&-T�lI�"OJ5��E�++W֬��o]ࡡ�"Oܩ�S�U�\9��p �N���jc"OvHk�g�JP�����r�ܭ� "O�)��؉��x���=Kj��J!"O�1�3��/bD��(2���Z�&�j"O^�y�&ۈ0޲5�Z�]�n	�4"O������+Ä��:{<H8r"O�9��\SV��r�-5Ͷ!H�"O����BA1E�����F4m����d"O0x�wEOZ3�e�y��#"OMh�T NC"��傄.���Q@"O*��І�8p��H����W��q@"O"�C��M>��]yq�T�fV�I"O���K�S��y��V [�L�z�"O^E���� o����")�7Mj��a"O���W���xT��3����?@��1"OrXs�C0���jј1�)�2"O�SP�22��	Cl��US�"O�%����~d9(ň@�}nx�'"O���C&��\��r�=^^� T"O*z���:s�\��� �L���"O� ��ȧc2�	"I�8n�j�i1"O��r��H>��1׈a�2e1�"ON�)�ܟ!�4)�
V�+~��"Of񂢏ήl�NT*���*Jx�"O~Y�m�8y\���]@L�p�"O:ыr�R�D�#��-�3�"OH��g'�N���]'R�2�"O��X�F�U"`�$�>EqCM|�<�@IZ��=��N��Q���@���v�<1WL#`�fp�V�ҔByܜ�Wg	r�<iTȌNI�b�
�|F���J\m�<᲋bn�l:%K���@����o�<at/��$]��s�F�[\��7h�<Q�d�f��-K�l�4�8��]�<��J/~��C�.�;eθ���aVc�<��l:D�x�R�$���W��a�<a���?kؘ�Ł��~���1'W�<�r��$
8���ԕf��s���z�<i�͟<5��S�D%�՛��^�<13b�	��/�mP���kK\\�ȓug�XP �ߥH�@@u��6Ұ��_X��Aa�Qx�������O&�Їȓ�z�!��7X#*��#\�rju��r��8�*C��[DdM\n�%��jwn�s!eS)r�Jйr$Hp{Έ�� J�H�������J�u�Bf�<� ��SR������bR�n'�@��"O��P�I�&r4,�pbG�* �mӦ"O�iR�*� \6����i���U"O�I�Їֆ@�A�+G8i���"O251b ݦ*Ԑ���M�$�+C"O"��f�V�J4�TU�:5j"O�����=�\�"��:�M�'"O �Ki͏,h)�➚A|ܜ�C"O�y˦�I0c�P���6L�8�1�"O� ��Yhu�.-�����"OLQb��LA�]��� 4,|�T�"O�A t �d����V&�Hϸܱt"O�)q7�J�$ ��e�;ļ��"OTPAD8�P�(aă��J�"OZcC�_�zk h�e��9c�
��"O�`�1H�8Q:<I�Vd�6~����"O=i����P�r9��ߕ^�b��"Of��"�/�^����2$܌��"Oh�S"Y�l1���d��z&�A;%"O�dy�fW��܃�*J�K�=sa"O��薭��ȁ��*-\ZX+�"OڠV�S �a�k�)1<�C�"OV!�ů�M/:p�@� G1Ф�0"OH�h@��5��l�c���3Ґ[�"O��p�HB��|	�oG�-��1a�"O����
wv�e�ׯǓPR(��"Ov<�`@
�GŎ�#ro��==��9�"O.1��D��.?%ڦ�ɋ)6�ݰ"O�aA� Ιgs"@R��q	"O��0�N!Z�f�j���tX>�
@"OF���,e�^�QelG5N �ڰ"O�!*&-W
/������,���YR"O��B����]��ً��Х%�$9��"OF� 2#��=��?a�9�"O1���4E�������+",}�"O��r)�"G|D�JB�#W^�@�"O�@��ŗk�8����4B�tz�"O\hD�_&=�ip�F� �谺�"O���Fט7
�%���M@n�Y�"O���'N���q���m�p�
6"O�=)$·N# �2e.Ī2ZH0"O:�4�?.i4-L�;8�p�"O,�Ĭ�1m�v8�'�6g��09�"O���>���"�L.w����"O~����ENP�CP�+)b.��"O���6� /�$�������U"O����P�v8d�a�m�#	�T`Ҕ"O(��h�b�=�,]����"O:ٛD"Ll�, Y ����9F"O���c�Ê5��H%��"{�&p9v"On����Ĉe"��a�N@?�f"O��R`S�d�r�F�/64(a"OF(�PW�^i|�P��%D��*�"O�|��bU�iZ/S<[%P<�"O�t:��=|��M�1$��W"O���`��b�a���RE�"O:��$��2xW^=���Ka"zc "O�0:v�Z��͠�O\�E�$"O< `��!��X�EI�7�^"O��y����]�T��H�Ӯ˱"O&���(Jn�;���;f��Z�"Ol�(%�G�N�k��I�;r:=r%"OnU��k��;�u �;e��q"OҨIFIȞ$��%�0�Z�LX0��"O� �i���	A��l���^A�T��"O&D��8\'���
R=�PK�"ObBRpr�y2� �y��`�"O �`���5G�Tp�e�#.g�Q��"O� ːH�
%�� �`b��a���s"O��X�L�,��}j�2[KR�K""O�h0��2��� ��UH��`�"O08i� �f/�|h��V"�%7"O8YB�4)l�����!:� �"Op 7�Y<h8���π^:$I5@'D� �@
�-�<Ź�N$t[��1'D�x�^�mS>�2���3����T %D��y��ŸN*�jb +y�����>D������9 J�����1�T���:D�\E���xŸ��̔-N�qX��7D���h�?Q"a)��ʓ�� �H)D� �!��4���@�J<c��x�&l"D�$zAK�,����W��)84��� D��X3AQ2<�z9p,��,����=D�ؚq�S6"nx1r&�c�Zx���9D����c2ȸ̊V-G<.�p h6D���c1e.���!,D��e�s�5D���a�3�� ��M0a�4D���d�-FX�P a��3f|���� 4D�lJ6�,���G_7?���&�/���I�h0�ykU�Ǯt�v���=��B�9v!4����ި�~� dQ� ����d�Y�'� �r# �|��dy� 
�65X��'X"�@A%��:�&�R0"�mb�����O?�	fÊɨWb��_8̐�r`R�s�B�I�0֬�z�A  ��<�vB�#��B�ɱ s�tz-ɝi����I�5?���� �D� Y��*u`P�XY�l���	b����p��0sV�Q7,�[��IȦ#6�눟nQ�U'W�:֕A�"� '����e"O�k��V&!@bd��4}���2�"O�a��Q;��@�
�,}�R5��"O�$��_)C�`�zWJ�;J����"O
y�qkϞ-��qaG_3(���"O�-Uŉ�>k��v&ߓ^0�H���9�S�ӂ�|ݻ�葝'U�p�Si�m��B�	�8��8V�ڀ7�h�e$��D��B��%X�b#N_�\K��p$A�4��B��.��H�ANK�y��Dñb�8gά�
�'�4�)�$�sEb��(D�zU;
�'�6�8�Lڦ�2 �_#C7��:
��MC�O�3_�2�JT?�z��"O"pP�$I�8�45����P|�B"O���k��_B��z�g��������;LO�(���)���vl�7G����6OQ� ��j�@��V�	,Q�t�/D�؁������$N"y�p`(LOn7-a�z�'q`ի�g�<�Sa�I/JRI�'�a}�.N�Q� �ؙD`ɦ��-2"�R��n�$�'�O���<�?9�O<5����m0���7����'�ў�� �!z�Z�k���pQ�!c�h1ʓ�hO�S�6е��O�L�:�s�gU�e��B�	Ou �ɂ 5[p��#ʑ�'3�b�8��ɔxi�i�S��2zPH��^0��'Gt���	'.PLm��hO�TP�	C�ҵTW���%�D@<{Pዕ�Wv6�%>�ay��	�S/@9{��1�TpD���B��
>(V!���O�iȡ��%�LC�*6ΚM�gnE�X��Q��W"���hO�>� ��!���
i`���j�����7\Ox)��"�!d=���ņ��p�ʄ"O^MyA�S�Z�Hd�2%�K�t�vOb���.3�^�1R��CP�5i6I���'��|2A�i��*��n[�9�e*�yB X',���I�j��K��ɭA,�O��m:��<�(܏5#�+�͊W��WA�G~��)§X�2�1�G��1!
�:s��4�D`���s�� � �>zoJa�� ;���Ӄ�n�|�<ႋ+OT���<~c�����s/����:O���D)��)���Ì՟?0��q�`��a}2�AIy�*�89ݰuʀB/�� HPd����O�$?�'!����-ǋ|[*pP�U�z�RM��"���
!a�;4���F)��0uZ�G~��~�S������J �]�z+N}�2L~�<if�ҰbD�aN�9rq�c{�<i��ƌ������&��� ���K�<����nb��B��i�u)Ej@S�'�� }�k�I�Q���4�J�fػ�ę5 !�Ė�m�9�2 <���sR�����Y�(O�>%13�0x2r7��B�!�J%�ē����c�C�/
pT�HԈ��"�dl���x��9�O���	
V�,*ck�<F�V�r1�`����T76p�TZ%�q��d�e �*@!�$D��x�Ko����D<=�6OB��C�H�m{v`De�1F�mt"O��KPe 5�p�b#P�A06m�"O�A���*��$�S��yz�"'�$1�1��'��T�7d�&e{P�ɜ<�jX��'��t!c��
+ ���Gy:Tб�'z�xXs��O�dr�
H�wϚ�
�'�Ɛ�	�66Ċ����"�J$�O>��D�*��T[gH�)|&�
t�F e�!��>��T���H�DyV@�܎�6"!�D���:,�,����Z)�'�	Z��A�'/�J�jC/\�K�bXy$(�4��ć�$�l	,�P��,D��	�� |Pm��f�	Zv|3��F�t�z��ȓL��Q�aբI(P�j��zt���<�
��s�u��2���&vP��~�\)"��pՈ��͓k����<����$(�^�PĈ�JHe" �ȓaQ@�����*��C	�T�ȓ�hqa�!�:��	�\���'a~������7��s8�=*RMǃ�y2(M�jd���؁rjH�#���'	ў�O� ��^���y'*��N����'ֈ�SD'UY3��Q�-ony���	a��~��H���a�H,;��0� "ך��>Y�O,��.�U�<@pL�.�L���'�!����R��	P�O�4����)_!��}�޵��h�@���F�ɫa||�UZ�` z��ٺH��T�����<��䚬k�jx��(A�x����)Oay��I�*��L�2�/c����۱4��B��(?^�yA�������gح,y(�G{����O�@㏞i|�h��-�^�"O��Y���>%�j��Ŧ_���Q�"O��	v�&?��)ZD�L�#q@��6"Of��k� 1�����o
.iP�`��D"W�'�'�T��j�<r��%v�$�3�傳EZ!��I0��1Fe	�.�D��8c!���%>�� ���5hi�U�FH-axR�'��ON� �I8rn���f�,�8d\��D{��� ̡z�,G�k�t�1H_�B�:a��Z�d��ɳ+B�u�B�{���W���!`�B�"trj���Pȣs�vb`Ԫ�}��d5�'?�����D�*?�@���X6"�x�ȓJ<M:�
D�ұ���I�r/��>	דoT2��薉�r�t��Z��ȓOJ��0`"X4�pElQ�p����mD8pH��Q"x�,h�k;QZd(��
�����O�v" ��B׶rv�1����S/8C�( ��,Ɏ�v��Bu`�K�nE��M�h�0{��ȓ[���Rd���*t���ȓDȅ��az/Rx��D�u����ȓt��m���������ި�>	��(<O�5I�j��zq���;b��y�"O����c�/h�x{!��T+�*�"O�0���C�
m 0���*"L��T"O> ��h��_�@�!� �#v~X a3"O6q*�RcO�c���E]��E{��	���Cs�A��zТ�Em!�DD��Y����F�ā����`R!��ǵ(p��/��D,��4aE!��#ᒽ�W�A+N
]:$�[�(!�$ΣQ��� �ٟRG��Eǽ�!����|����mJ�(�߯VQ!�D"���A���� m�t��}!�����cGGJ��ּ�È�~"!����@���iUO�)"r��`G��_!!��Vt�`�&ED����󲧇�	!�d��`M�����Z�t8�bh��!�$9���j��P����Ѥww!�Țk���ǭF5A �Z1珷g�!��E�a�PY�B\7��Q5FWC�!�ŵ��}��ȍ"Q	 ,1#˄�k�!��y�ؐ�ʌ�6�U��
�!�$ۓPe��4&L��Q���
�!��Ȼ
%�ui�'�V�z�*`��G�!��-uT�Mi�ˆa�R�H5Ñ�X�!�ʞ?(�<���Gx����8'�!�䁇b�@�	����T�b8B�"F�E�!���IrL#ׯ˼]��kE��$�!�D�9>�6���k��"����	B�!�$�|5r�Cv�W�Z� ������!�u��@rP�� a��9UnȆ�!�D�6�D��CC�0	����5m�)�!�DN��l\3�.;V����6;!��2t�83��V0p�@��CX(!�d�60
`�H�(ǦN!��?:rBM����0��Ͱ��N�\!�$F"k��T(@�i�����%��V!�$J�%ֶŢfeЫ�����*�!�d�F��?&�T�0gI)VT!��,jń<�Ɉ�b��1b�jQ�b�!�$��{
:]�� J"X|1�ȅ~!��yeP��^*���d]�|\�t�ȓc��X+�̅&���k��a�L��ȓA�8���2|>����� Ბ�ȓD��k�-�*�"X��(�t"��ȓ,<���F�+���c����'��\��ua\5ӳJřTL�%��K�4c>l�ȓ\~A8�J�4$U&Y����:y��|�x#��@.Y�h��GA]��8��ȓ��Œ8~�0{��.,
!��_�<�DmP>|�)�O�sJ^ij��[�<� 0�xN'�:�K�+��섐"Oڌr�/@7(`3��P P0(�"O$�Xgl5�D��ę�\��2"OЁ�VM�>����DݽU��9��"O�D��ȏ�/�L0;� 4rƜ��"O�M	�I+cІI)��*W�-��"O"䫐���w�ŉ��X�nY���"O���i�<}���$�<�h�"O�ՠ�)I;B4Bb'G�L�8��w"O��r��%�ؙ�`��M����"O �2��.܊ �� H�X��S"Oz�*F.E�� �3m�k�zs"O��[PI(#3��g�*O�R�Ƞ"O^$хbȹERy9ӌˢ���q"OF��j�G��#+�7Q�D�'"O:�kw�8g�x�k �9�*�b"O�L���`�1�"��$�z��t"O�	Rn� iZ����J9J�8�Q"O4��1D�a�L�k'�I�vZ[2�(2qO�)	��Y�@I��-�v�k�G�Ri|ZGK:4����Τ��*��ē<6S���l��@��.��c�a}rɚ}80Ax ����kV�L���<��d@�.^���̜�~�o�u����E����u�B�<���9|k�a��F�p����b%��d�H�QU%ʋ}1t�1���ּLu�����:���H�ww!�$�6����U�IAy-	t�	�`��+C�݌^��$��1J�@��L>��k�.>�Y���r�<���C�I_|��':Ra�DA���xR�y���Ax�4�s�&��Fش,��/�H�"�D%Md� u��:�����ؗ!�9��ī��a�d�O\lT���@1H�G,�v q�|��-�t�=�}����$D�sd�@;:0B���@~¨Z ~6XT��;>�;��S�X�.�:��/9�$����ٚ��"}��	7���}&�8�j����h�*CbE�N�5�����)M៤*t&P�D�c>�cʴ:򨚀	����bӄE<�h�mނg���`K	*�{�h����	w�K�@��� м�l�r'�v*�Z䯘�0�	�>�RL���f
��#�B���ڨ6F����i��0��7#I �0<!�DI�,���־N�X�=u�!Z&�ٶs|8� ��m�@|�e�}�GSu����Ħ<w�?�jq�irK��Qq`ym��	����zB���R,8�R!��H�O�rXa1K�	kX�x�� �r�4�Q�+F��𝸦�+� �jw����ɠ-3fd���[�/����a�DȔ=��CG?����9.�I	$,8��O�E)D�آ);t��jI	KE ٳcH�d�*SL�{������A<:�z���"������3 bTK�˟2f1�p�U�h��C��F�u���S�hk�`kԅ��99���EO�2y<��~�,s'삡w�z����S#P�H��]�	��a�c�L�H=2�'��0
��ލ|�Z�i���E��J�#P����Ḡ#��9�*W��<�͞���͢XpD��Ѩ-B9)������R&�"45\��Or	F̓Fod��%H��?��OW�`C�(A���~J3,�JZ��v
��� ��1�⠉���-m���˛�vaQLKX�'>�ښw�����H�-S"�XV��0��Bg�YIo��	�dF��1��t ��$?��K^�s����� O�Č���(in0�2�@�=B~!��̍n0����F�)"0
d���J�֬�F�˨��J=ޡ�b��EɆҶl_����p�C];,�,�I�L�O���Q��
5:ԍ��S�B��8�&L����X��}���q�*e���Q'C�D�9X�v�(�c�3dx�s,��D �b��Sl D!�d�����G*��tC�D��Hި���k]Y`�z��ܓ<��ڷ�E�6�R%k �^*v����/��n����%(3����p�%E��]�$��_&-��O��Y)�>MY�Y��4'^h]���ĕ>�6	���˽����ߜp8�)�����3P�[��â;�����Y#]=x�@�X�#W&�ɞ�t?�1�c�7Z�%e�˖`��R�S�+Ԅ=�t�Z��n�Pqj�<$�HU�-V/BP�Љ���$����?��-�L��- nV%��F�<QKx5
	_�,���1�T�`�S5d�"B�࡚�̀�j^=�0F�<��

�WLT��O/s�t��BV	ei�d9$�&(l��G��}/j� &揕TNP���/r�@�wB֊be�t$�G5|�r�e�/Fs�d�t��+F��1$cW)sPp�
�'ȴM�r�*O�M�Eː�$�&���KJ�/t ����#g>�$m��R0T�A�E��H1Q�B�H�b�UC ��N�XAI�!b2���=�M��#�/2�Z��E.�6 R�G*Hͨ0Q�Ɋ�r:X|�'#TQB6��(H\���a��Q 1ѣB�&`Y�����.��IdT�}#�E�N�ā����>�Bi�E�5'SL��j]�*�6���0�K;lA��j�	T�rR�% g7��9�K۟��P(7G�qKRD����f���!��qu��`g�ŔO���k�|�r�\�X*	G�p�Ma�"ĕ^=B�2��"oa,�zW�U*��KƋ&P�2$m��\�:��ʄ�.�t�@2Ż>Y_�����F%<������ur�|�E>�f|R1��9�TXW��UP�Ch�&2�����D�vy�@a�ET��l�8w^�\ ]yfM5Y�]a�(U�v��q�@%Q�rk�t���P����ӆ(���;�F�z��)T*�9\����0�83�u��W�ޭ3�ǚ��8�0;�q��R�ՠ>�̐��2�=4���R�٥;�ϒ��;����Qu.��Z&�%�+jv����Qu,��].�.�&a|����Wp*��]!�#�/ hw��I�_����2���l�\E�W����?���a�QN�Z����2���d�WI�B�:�u�OB�!&э�{D�O9N�0�r�GJ�)!֊�xI�@6A�8�t�OB�!&Ў�|N�G3C�>�#��Wb/`}��	�~:��./��Xn"cy���s6��)+��]	k'gz���s6��))��,�a=�F��Q�W�~,�{(�i4�L� �Z
�]�v+�{(�h5�L��P�U�q.�r �fr���;r�6��3u_��8y��	�=u��0�0w~_��8y��	�>q�8��8yW��3u�� |�?�*T�_e�Y�9'��]v�>�-R�^c�X�<!��Yq�2�#[�Pi�Z�3.��[r�9�'�2��	���\
�Ƽc��E�'�2��	���X�εi��M�-�?����Z�Ÿe��B�"�1ۮ�S�D��Bb���/�tm�ܪ�U�E��L
o���+�pa�ӥ�Y�E��D e���,�wh�ٯ�Q���?��5�f��Y�p�
���6��8�j��R�s����7��1�d��\�~����������{	xu�|���e"�������tuv�x���m*��������~}p�{���m*���������~�Eg�O�^Ex�9ZeBi����{�Bf�L�UMq�7UjLi��z�Oi�A�TOr�3TiLf����tj#��#sT�6��hD���o$��.~_�>��kF���o$��&tS�1��aM���b)m4��Գ�M���|[t�p1�)`6��ڹ�N���pUt�}<�+n6��ٲ�B���~Xp�z9�&n9��������G-�`H>��+������G.�jC3�� ����J'�g@4��&���d |����4~v�������hr����1tx�������os����9s}��������b�u���
��~�"�����~�����s�+�����x��� ��v�
)�����}��(s��_;����O������*q��_;����G������ z��S0����E������!x�ꌴ��:�L��>����|�>�:�����;�H��?����x�3�8�����:�B��?����{�?�?�����G~�y��f5w�� +ĦBy�r��m?~��)ŦBy�r��k8v�		�
#ϬKs�/��K�� M�(�Ё�u�� ��E��#N�$�І�q��*�
�B��/A�)�ׅ�r��.��Oj#�=',/�(5a�uİ��Kh#�=',.�+1d�r÷��C`+�5/$(�,1d�}ͺ��Ae.p�!6e�ih���?��h�p� 4o�mi�����2��o�v�!4k�gg�����:��b�}�+>3��>����-��I��׍��6��;����*��O�z�׍��;��6����!��A�v�܁��4��8k+�
�H�_ ʲx��ތ��i-��M�^ɾt��ۊ��c!��A�T��q��ۊ��c!��nKH-" ����*V�������kOL)&,����"Y�������jNN*%!���%Z�������jM?x�ge�Xb���5��;}�mo�So���0��;}�mo�Rn ���3��>x��O,�jD3���I�0�!�G��@"�dE>���E�=�"�E��C �dD=���F�2� �@��G"דy$�E��JH�FM2��g�zz&�E��JH�FM2��f�y~#�B��LM�ND8��o�sp,/��- GE^����69�@qY"��%+MIS����0?�BpV/��- AD\����4:�Ew^%�� 귗U+w
@m���i2-N[dF귗W(sGe���a5%FRnM漝\#He���f>'F\aE跖Wa;�h&�L_Cd� ��rɝf"g:�e*�DQLh�#��qȟe&b?�m#�HZFa�%��pȟe&b?�m燹T���Q���WO�-C퍲Y���Q���VH�(@W���U���^G�&H䅻U�24��Ú/����m��g���36��
Ɲ'����d��c���36��
Ɲ'����d��e���8:�����Q�������褷�����X��r�����⯼�����]��r�����祵��������eJ��dK!�"�E��es����eJ��dK!�"�E��es���oA��i@+�)�H��h~���`F�j�ϜȨ�-8����.�A�c�ŕ���/9����-�D�d�ÐĬ�/9����.�A�c;�Qc0'��"��uN&�>.};�Rf7/��-��D*�1#q0�Xk6"��*��}F!�:-;�Q$��շ6Ƹt����P��$��Ѳ3ýp����P��$��շ6Ƹt����P��$�ɻ�/ҫ�A��� �0X����"١�J���)�;T����-Ъ�B���*�=S����/�8�D7�n�f���f%�,���8�D7�n�d���e&�. ���8�D7�n�d���g$�-���2�H<
��u�D���?�_,�6�q��{�K���9�\.�2�t ��~�O���9�\.�3�v��O�Y85��yl��	��O�Y85��yl��
��K�^0<��qd����K�[9����;W��6w�
@���ߖ���=P��3s�A���ߖ���=P��3s�A���ߖ���Sd@�=�8�g������WgD�:� 0�o������WgB�=�<�`������R_��r�q�r<r�`���X�5�_��r�q�r<r�`���X�5�_��r�q�r<r�`���X�5�^���3�JS���D�8��ǮK�1�KQ���B�<��ǠD�?�JQ���B�>����N�6�M$녠�p����*���k�'$녠�p����*���k�'$녠�s����"���m��#!���8ς������KȘ��
���1��������Hʛ�����=ʇ������Jș�����=j�+��0d�(�����F�j�+��0d� ,�����L�m�/��3g� *�����E�i�)�qo4�Й��<G|���vj=�
ݔ��
;Ay���th<�
ݔ��
;Ay���th<��!���*&w}�`l6~�ө�(���+$u�dk<u�ܠ�$���)#pu�he3{�Э�&jh@u�[.����)QM8WlmEp�^/����)QM8WlmEp�_-����)QM8Wnn@w�F���؊�X���˶���U�O���҆�V�~��α����Y�G��߈�W�}��β���T�L��6���n�ev�;v����h6���l�fu�8u����h6���k�ly�7x����k4��6� ��g�Y�$�VM!g�=�(��k�[�$
�[O!k�6�#��`�Q�, �WM"j�2��삯�<Á[t�z�60L!�킯�<��^s�q�;=G+�ꇬ�<ÁZv�}�?:F+�全�Y"�ļ� �gu��
�ŉ;��V#�ȷ�*�lx���́2��X#�˳�.�mx���̃1��^$��2�<Euӑ"���1y�D�?�6BpГ"����<u�@�9�7L}ۙ*�x
��1y�D�?�6K�A�,���m�rif/�97�)C�I�!���`�tob,�97�)A�M�&���h�sif/�97�)C�H�p��a�-�\���۴`5l/}��f�-�[���Ҽg3i+p��a�-�\�	��ӳe6l,x��l�fi�b����2�
�a�7�fh�f����8��d�6�fh�e����4��l�5�fh���F�8��gj�8��Q]��7���B�5��dj�?��T[� �9���E�?��kg�4��]^� �2���M ��r�)��p���!܁J�D�o۫V���o�=`�&z���J�	�?a�@@ i8����)K������;]�}����	�r���I��������m�@,��}����Q	�Z�
]����h�g	���ii�\�\U���	�T� �K�U7�y��'M�J(H�Yᬘ��.--	�m)�D�*B��ܫʩ*Ȝk ���9�rQf�Ԥn^�-�������IF�f�LE�I�/а;���ف��?7���w���Rp$ԝR����!�"Mջ�4R��ڣ�ٜP9~H)£x�4�Su@I�>����cǅF�:(�W�S�Q��a��̍1d}jR"ѯ8�j�ɐ�'��Ȑ�% (���NF��Ɍ� i(��u1�l��!�����B�%0H�x���	%� �X"��
+6pCR#�vZ�p"�A ����Ba��!8X� W%P�'��@�J�	�R]�AAF�d� dp���\�'�o�,�LT�E�^:��OV�^�?���d��$GD,�"'��(�Bd&��dy*$B�r�la�!(Bh�dhA�$FI4�'�I��?)�f�ni2tB��5��9xM֕8eV8Q��·^%�]R�y¥B�]"�Mr�
���t}�3�E�DX X����&3G"`��KP9F���P���E󢀣�%K��3��Q�"R�'L6@��ː9G���`�@a�dZ;x`֥H"�P�
���������'�
%A ���@�8~8�Q��:|i(��������-���'&^	&�lc6��=��Av�0y���䖰g�d���b3N	�Ǔ&eL�qd�����M����1v�(sr�DE�t�P�޶}�J�Gβ%bB�A4*(��E����u�	x�\����g/
�R�*�5�%cAm�e��TCi��W9�Xbv��T�L%�$%�!ٜ�y��$c�.��ϔ"HXR�P�-��uw�Y�sT��h��<A���#�f9�h�Xl�Ux�F�LG�Y���'~b�!v��ڟm�/���y�� !�ΜKD O�1�4����T�Z�i��A������l���Mb�j �/�I�B�>�Dd
7�\D��
�-S�$#>As٦y���h��PJ�N���JR�1��e��Ǟ'>O��A�КR{^]�6//����LNU\���<t�P� D���t�ª@�Un橃���!V����Ƅ�.��R���%E�t�8�B"aZ4�B����,�y��v��=z��I�+��HZ�J*�p0�H ���RˈТ��L~��T�d^>_L@�9���2`V5�w�	�O�!��F�p�DĐ�QߦS���E�� ��I�-��aa&(Æ��x�
��C������gb� ����=����F�Q�r�T475l�bA�ҥj� q��iC�wM��b���Px�%�J'zUR�,�D�<}y��F��'^ڸ�!A��%<��%���}�q�B�K��X���yJ�g�E3Bف"O���b�:%I��@rݼ_E��$%LC+V�$�'S����h���0մ���ۢ\��)с�.O!�DX5T6�]�G�#�Hx:��
 7r��u� �QJĦ"^���I�8(�(�U�et�H��D�U F����"d#й*a�T�s�\��L���\kB/_*2��1��*4����E��{�� ��L%h�{�D9�wI����%J�z�#|Z5�'K�d k�(O�6P�l�o�m�<i�)>p�qCD@ַ$"��5 �ş��#��DqO?���҅��}s���2y�.4J�"CC�<q���$`\��Q�#����� ~�<a	W;$*"$�#�0q�e��Tx�<��D(6��-��� Mzh�e�{�<q��ِU'\�Q�N	7�l���p�<��g��i�����O�,l�bf�r�<y��71�$�{*�n ܚ�r�<9���]DJd�Ыs�PR���h�<�C����I!�%;ݢ�J�Λb�<���/l�p��Lݣ�U
e$[V�<�t�U��H��P�6��E��DV�<�2"W�p��;��2D�f���M�<�p�H�fx�H2�Y/HDx�J
p�<�Ŏ:M�B�Cᅕ�U�H��!��l�<�a��)�%J� �6e&$Z�S9LC�	��F�2"���S�I�2�[��3D��*`J?}.��8��O�$܃G>D�j CL_*�5
�*�ʤ
3D��a��^�M�н#��K�/��x�d$D��;m��/EpI
��Z9�����&"D�\�Ԭ*+]�l9f��Q�"f2D���N,��SE��Zs�Y$m%D� r2��U���`�ƯI�F�b�#D����d�"|Z���񁅭X�][ D�|�"�m�vY��@(T��)�m?D�`h�@Y�
�@C9`�e�a P13�!�D�<]N5�� �.��U����Q�!�� �ٗK	�$��G^�'��V"O��r0-I5I�P�C��5;�^��"O���y��#�/��"O"� �l��E�q!�G�0�a�"O�s%�^-A�X�
۲�
l)t"O�H�BovV)9n)w�T �q"O��iЬ
�,0�
u��!8p�0"ONXjAjAU|���"�;aI��:�"OV��v	 �+�h�"�tD�a)0"O����,M7|������ֹp����"O��3�4P�ō/J�4	`"O`a�3aT7d���aeBz|X�E"Ov�P)^�8;�\!����s�B��u"Oܭ0��V�:JL�aB�Dq`���"O|����	G&p�Sf޿|F�IA"O��[QìSWd ��5'�\c�"Oh$[ O����	�'R�*�"On��v�C�,�jl[��B%T��ؐ�"OB�QB �&%,�S���S��)�"O:�R��mŬ���IT+St����"O(|�p��?N5�G�S��Ј��"O�03,��t�9Q¤��T��"O� �ѡP<"�|�BF��'j��4!PE�"qO����Y��)�ꘓO����9~��.)4�˦$���<ȱB!QtuRmba��mHd���*a}"F��.3���PMO6N�@k���<���n�:t�nV��~�eM;&BXQ��-@�`�u��+�yB��]��eIՇ ��<��Fn@���I?8m��m�=���0����ys$��n��<��k��  .B䉤.�����f%�,H'Ae�h��*^�C">�ɺ��h���|��I�!�՘1�S0"�@Ip��x��I#�����<���yr�Q# �ji�Qa��;{.�S��H�&��{��Y,N�
���-"��	2&�?�0<ae茜j�̜p!-�5w�p�ᘍ��,�3���)�,Q�b$��!�lь�qOq�:�x�n��C�d����$!T�����0��@oBX�@�HZ%�ԥE�� ;]ߨt�!�=��  1�	�+
T��M�6��'S��>�O�T��C��K���O�:� 4Cqd&?7�����OP�3�1J1��ɒ6����81���C�F�8H�1�Q�̵k����S�	���=�f��D@fB�qp�BOL~\�|� H�b+�Z�G,��$�P�[�΂[�꙱㯫~"��Ӫ3p����1���1���m�<���9�������U�h��-�& R�ђ���Z��YG7O��j�;�
��5 ��vp�`E�DM�6#db�r%Ǝ�d�8�D����L�;΀!(�)�S͸U�V�,ڧ#���������ѩ�t���r/."h���K��D� ���o���ņ�P�u�V�n�>�2
�^�H@��0Yh��S�A'�d�E��'%�t�5
Ą��qB������ƕf�Ĺ
��<b��]"o��dPaד~���+B�� �p�A5��; ��l�U�Y!L:�X0+F�Wv��'��I�I��\;��Z`�OB8���ܟ6Y��%���'ǝ�E��
��'FX(���s��cK��<���4v�S�#X2>�+ǉ��_�Ќs#�; 6��A3 Ҿt�0�%k�5t ��O���d@��Xi�9�@*W�o02�"�E@�j���BC }RjK�
��s�FPeL��	&Y���X���J���(�uͅ;n�I0eX�b���!��]�V�#ц]'Z�!@�	��U��$�E����I66����r,J$ R8 ��<c�5}e�D�"�� s�	3D�6I�W�ȵs-�O�:Iˇ	6t#PP�+M8\X !��d��0yUb�O�>ͱ�Ⴥ��[)NW%d`��K��I4H@0*�d�!id6Ps��)]��`L�k!^���4پ����?
���VbE�ko$p`mJ�X�֩�ӠL
h%T�^c^�1R2 '"���p�c �<�N���#$ d��Y
$=ٓ��
%?
��'�1a��CP
Y ��Ň;s"%�3�!�.mP��FX�'S�=�rJ@�E]QXw�Աܴm75 %i��,������9	Z�h�03�P$��b�d�`'`̱��iv<Հ�S$���V,č9���֯w"�F�\@*��fP�9�f�bwA��dT��D�2f���W-s,��a���XI>8�1f��yg�A6q���㭛Ua<��a&V�<�p3�i�>ܼ�a��i|���	�p��'�R�Ǔ�h��\8S���)w�(�����~)J���%4������1:8\-���)J]�@�.(u�8�ӣ�rya�<	��};7OK�#z�[�	GהU��ȟ4t� ��<?�0�-X
��u37o�"z�k��QA،A���4rH���,�I�(	��= �i�@�=ǆ���/S�u�\�#P��'ӾH����Oj� G���P�OJ�n��v��[�4�x��ЈR�,����`���u����P��1h��9C� [�]� �@�j֖^���w�0^'���dO�v�`e�'������$~��[�kʭ[�~���
�-VBD�/A:`��4 S�3 5�����ɤi'���M{D���"�&%je!�6&��h���%@lRi�!P�E#�.�\���^�����U��)���ٞk��R�����Y��/���Ԛi��V�����U��)���ߖb��_���"M�_���F[fZ ��B��+D�T���IUiV/��J��#M�_���ASjW/��J�� H�>��>�:Ĩ�P}v3 �<��6�7ˤ�Wxq;	�6��3�6ˤ�U{t<�=�ۘ4t��6FV3��gz��}В<s��>O\	9��b~	��}В<s��;HT5��nt��qܘ;v֭����+RCR���N~�XЪ����,TGQ���N~�Zխ����
!XMY��Iv�P׬������ta���6�	�a2�	������ta���5��k9�������~i���3��f4�������"/M�F�Ctx����þ�2-l�"/O�C�K~s����ɶ�7)i�%(J�C�@vy����þ�2-l�"/M�4�%	S�Q�x�x3��y��?�,T�Y��3��u��6�'R�Q�x�{7��r��4�%Y@cȤ?9M rBUar}�O�\Ef͡8?I*yNXnq�G�Y@cȤ=:J(xNXnq�G�XDf���w�ɔ�MPt��ܽNM����~�ß�G[��յHK��������EY~��׶LA�������M�:��|�\{LJ�pH����J�<��{�YxNK�pH����J�
?��|�QpFL�yB����CgN�����y+��]�[��mK�����,��X�[��jN�����u&��^�Q��iL��f�=�����h��hl\vqU�f�=�����j��oeV|{\�n�0�����o��khYpvR�`�>T�J�X��'_�z�8w�8U	�M�Z��*R�v	�?}�1\ �N�Y�� X��:u�;V
��)F�u�xgK�l�=�ؑЊ"uO��ukA�g�>�՝܎!wN�r�zeH�i�3�ٓӁ/{E6�0�`��>� $F�;�=�p>�o��:�,N�=�5�z5�e��9�,N�=�7�2�(�i�k���)ow2��Xf�'�l�j���!fy=��Xi�(�m�e���#e}<��Wg�%�c�Yw�9�i�\}�B?\	�YQ�\r�1�b�Qv�E:_�YQ�\r�3�g�[z�H6U �T\�Q�� �vn�ϯ�H�͂7�8�6�!�	|m�̬�F�Â9�5�4� �
w`����D�Ά<�0�9�-�q�r��%���Jr�$&Jy�s�r��%���Mx�)+Gr��}��*���Mu�.-Gt�x�z̤K#;�R~�]A3ц����G/6�P~�YD=ߋ����@-4�]q�RL8ێ����M&>E1�{-�~θ8�PP��e�I;�v �uõ2�]Q��g�I	>�q%�v
ɾ>�_Z��b�O6��˳� o��{������q
q�ͳ� o��r�񿤮�wx�����+e��w�󾤮�wx��Ž�J�`
a�4���0�j�Ohg�E�`f�0���0��f�Njj�O�a
c�:���7�k�Kml�H�m��
��I�Cn�����T����� ��D�Hd���ĸW����� ��G�Nc���̰^�����
[ZR
@&�����B��%�FTZ\J%�����E��"�D^_ZL&�����F��%�FZZR	"�E뼨5
���*�D��E�&�G뼨5
���.�B��B�.�O㴠=���.�C��O�,�J�uO��@��O�����{[h�wC��D��M�����|]h�wB��N��G�����qPe�}�e�=��^��؈� y}��,��`�;��Y��ߏ�%||��/��m�7��Q��Ҁ�(pw��!�
�`�Pf��I�L_���܄��r��Rd��O�MZ���߈��u��Xo��E�FV���׎��t��Xo���p����o/!��@R���w����`!)��O\���u����m".��L\���z�_C^:��ЮrѺԒ���[DV0��ڥܱޚ���[DV0��ڤ}޳ܘ���^ASz�w��cJ'1Z>d��' [js�y��nF,:V1i��$Yfw
�y��oA+?U?f��&\nr���|"���9�v>6@Ɠ<�	��~"���9�v>6@Ɠ<���{$���?�s81H̙	5��t���=�xU�!g��i�s���5�t [�!g��k�|���=�
yZ� e��l�t���0��䝷�KZo��%��dg�E�x��䟴�M]g��-�co�L�s���CRg��(�hm�B�{���7���'�3n���8��}`1~���)�=a�
�;��~d4{���"�6k���:��~d4{��zK��j����y���J
c��7�p@��g����y���Kg��4�}N��j����}���Ci��=�xI�6�Ta8�x
K���M��Tr,O6�Vc;�B��D��Qv.N6�Vc;�B��D��Tp&G<�ZhKg��tS�A��dZ7�*Me��~Z�L��l^<� @l��y_�L��n
Z6�)If拻��@(1���9�^�]��"����@(1���9�^�]��!����K%<���3�S�P��(����ԁ͖��CL��ư���J��<ӉĜ��JD��²���K��8֏Û�O@��ò���J��<ӉĜ'���-���OB�c�ڈ4'���*��	@O�i�Յ8+���+���GJ�k�ދ6'���V��2�*��B��$r���`�W��6�/��G��&s���`�V��2�*��B��$r���`�V��Pl|�"�°���K2ߔ]aq�(������@8әTo~�"�Ƿ���F?ԞPl|��y���d�⟻�#S'Իs���y���f�᜸� Q%ջs���y���f�����"P&н{���u�[f��7�hY���EVW�+Ӗ�wTj��9�gP���BPS�)В�rQo��<�cS���BPS�)ѓ�pSn��V�*}���w���R����zV�*}���w���P����xR�-u���~���X����R�(|���s�r�:&o��]��t���w�t�=!k��]��t���w�t�=!k��]��t���w����K�$s&���&?��]����O�#{.��� 5��P����I�$q%���/5��^��������ҙS�����h��5_������ҙS�����h��5_������ҙS�����h��5_������� ��z}�0�	x�9���F#�����x~�7�|�=���H/�����x~�7�|�?���@&������3ܒ1�oؔ��z���"��3ܒ1�oؔ��z���"��3ܒ1�lޓ��r���&��6ٗ��}�8�A�a��;vz�U����r�6�L�g��9ux �Q����y�=�D�b��:wz�P����y��bC��6V7���^���[�bC��6V5��W���S�fA��5U5���]���X�`A��A�*����7�f�~�� �G��D� ����<�n�y��$�D��F� ����<�n�y��$�D��F�s��`��c*Y|�%�́���F+��i��f)X~�'�΅���O$v��e��`(Zy�-�É���F({��g�%moz�r��'h�cds�=��.� hj~�s��&i�cds�=��.� hj�q��'h�cds�=��.�#mm]�L-}�4�}\�����(�-W�C%v�9�]�����#�!X�M*z�6�}^�����)�,U�G Rz� �1O��j����v�F�'Rz� �0M��i����t�F�'Rz��5J��e����~�A�$Pz��c(��h��|�7�4k�m-�i&��d��~�7�:f�o-�a*��n��t�?�0m�m. �f)koui[���
�+;Vnk�inui[����!0[c`�aipjY����.<^ga�`frn!�6���8>I�Ƞ[3ꨀq�/�7���24C�ŭV8ࠈx�#�7���67A�ŭV8ࡊ{�&�0�6��J���G$�=1?=0N��9��@���D$�?2;9=B��<��A���O,�8:220N��9��@ 	9���T�t]����U' =��M��G�,J��'r��DK�'��,Z@gP�a�(�'?9bO�O�`�R"�� U2�91��T��,���&�=eat`�a͟=ZD��; ��X�*�A���I?�l0c�6-vY���'���ˑ��6<E��
��>��t#�6
#lQ����O�� �JMo������((��� f��������O)+|
6�?�x# R���A�厂V\0���45	2i�6�Y.4̉$��5}��X��k ��ɨ@ƐE��o�`��l�F�H�lZ?}B4�
������	�/�ڽ�GD�~�<��9)��!��\�zI��w���򕻲� (�ā���'�*8� o�;-�K�ag� Q�ek�~��f�1Ok�)���~҃׿1�}J�@L�6a����7D:p�sӯX�7	� ���j\~-K�72�"a��̏��XD��E�0E��]#N���P�qoEoUn5;4k?n���y���D��Ш�͟�p�F(��i~ ,�@�ܤ�[��݊ A�͛G�	����ѭ�=7� P$�-y0�W�	��s��;iX�M���O����*��r����&eo��V������+�.p�'I, 
s�M�d��5��&�&z���B�3�ؼ"6�_na��,|J( Cj�)g���e���{���'�C�5]�48S�[�Y�p�`m�'v������Ѵa��9�F_��f�������7lÑ.��×A��4i��4�,0��:~���਒5f2�M�C(��ç�ߟ\sf5|�$<����5M�:�01j]��B�Kw�ſ�X�<AG�E>�H㴪�ƹ�1M�?v�Nܣ N�6V��!�'�34b����CQ�1�N�(�Assd���<]>�ϓS��	�G�5a����1}�)z��"��+hbD �g璡A��O��.�Р�V��#r(���~�������)kgB,�7G� ���=!�:��uG'�E�â�8?�|��Zevd�A@�59*0��K!O����K�>��U�7R�^)�1,Ma���Г
Z7KYA3������ ��<��Y�4eQ�Q�\ם�7:�-
go	�]m���Pש4�����ݧq��~�)\=$�Xe���_|-ν���ߢ#�l(������a�w��Y��z� �Z�ݿ~S��(����z��d�WZ>���[1  ���)Z(=�v�"��^8���0�K'h�"˜�p~�mʦ"�#_�Iʡ/���H|���(]�,���%�tE�1��6Ȉ�'�.����L�W�2�Ȅ��~�����̓Z��D|�*���$���҃W�1��B��DE���9N �VIV2�� �g�ޝ#����36�` �G�e.�I���>i8 ��9<6 k!/I��]#@A�^�cÃ��q��i;f��)N�6�"�怣 �A�"O�웁��4V;��������bT53��T�G�D�*��I:\�O�N�:I�4��'� :'���,#�%$D�	!	D*���8�d�01��8q�b� �`ß�XK��є%-&��$����ʖd�7^��*�ŜP�a{���[ͬ���jۜ<
����njl���oU83��Aˡ�!JY��D�4��)����pxKV4ZM�a��}�V�s_tM����8A�l��	H��΀6T=#fG�jUnd��'�z�Q�ID�-:�`�+\���i�(��v�Θ��Y�1B��S��~rd��u�r���=m&8���1�yңM��1eK��44ݚ��#�?�!��Q�
tq#��,8�n��D�o�t�� �_�JoJ�`�Q�.a|B��+:�aq� 7X���U>e�Jq�b S�mp@1�O���`�zk��E͒P�	TB��� Z>��u�7$ZY@��Sf�v5�P�-D��0��HE��M��N�@2 ��O��A��˸����({��3�X(4n�RUH���@:D��k(O�<��x˥��,s��xU�4D�0�B �	}0Zk�hn���0D���5)��������ɪY�j<p�G1D��xf�ߨѪ�9t�F"�����+D��he��-�48�С��6���Hb�&D�܀�������'.D��rU>D���r�(e�6�2��^9�����*T��� $ۃ2j̗21�2`��yb��mB"a��A1���1�����y"�] wĴ�Ą�� �ͩdHM��y�� �3l���FD� ��֭I�y�n
?N�)s�͌�d�N��yB�əvP�5P*W�XKR|K����y��;O�E�t,é$��	IE&V�y�#P�U$i[�
��i6lqr5#;�yRl� DfPx�̥C������y��˪z��Oݳ	�:��!���y�]�INԍ����_ NQ�ȓ0f,0R��x�F  �c�>GIz͇ȓ#�sc)!3ZA����*2d)��b�<4)1��*Z"�@p1NZ07|XD}R�b̩�5bH���v��T�g�F*9ț� I�i���b�H�x'l�*�Od�i�g�? >�𡦓�O}�M�c#��9����Èk8�[rl�!�)6�<!�Td)p�$&&q�\�ٓ�3?A4lP�L�D���5����3�M0	�x��aǘ~�L�0B�O�MX�ON�S�OS�D`A��@,x0�FҴ@��h3+�d-?��>��O�gZ2p>Z�HՁ�V�`�o؎f�'rZU������O]���H�r��m�T㙨.󄬡�O���'αO>]��)�N=��ͅ
b�<�01�a����'�^b�"~B�D@P.�!����l�4���D���_�S�O <؇��/@�H��+�;>���b!�>	�����
ç*��rd"?N���T�Ɔ5x�t�B`ɩG'p��'74�ɋ�ԟ�NS�==҉���G�6!���Vƚ�FL�' ��oڵ)��lF��	޾ZR�� M�5��qc暛��D´�Mv`̛3���S�O�K��:�z����nyYҍ�Da�i��i` �����dˋR��V�e��9��ڲz����]�N l��@ƙSx�F/�>��'F	P),Z�c����ݕU�j��@՟�3!j�XQ��k>e��	[;[����b��V�z����O�A��5O�`Պ��p�(�)�s���B�G�`��E�ኜ�*���1�O  �UW���9�ȟ|���ؗ2'R�D�E� �<����'N�y!c�MX ��Myʟ���) b��
����7�
*l��m�4-ۂ wX�H���x򨤖�蟂�e���FfP�i�#�T�΁��\wjbt&�_y�n>��ǽp\ Bv%�	���z��!Z��#΋Dɬ��/g�n���I0[2.\8��D������)��N.� �5ÂE?	e�O@�p��ӹ�r��� J�@���q֘���OT��`_�b�6h���?#<�Gn�6��Ѝ��m(���+Jk�<a�	^��52զU�7�&��v@�c�<��Lɼg�R����=\\ͱ��\{�<�p�F� ?�ĠW��!+`�e�s�<��O:y|$;@�Yr2pUlPG�<IƇ�)�\В��,C.�����^F�<6I;�.5����v��h���K�<�$���< i��� ���!�R�<������v�_����@�Ǟz�<��+���x5	�ijD<J��ML�<e��`p���B�9[�Nu��]�<a�`��Z~1�n[�d��`���\�<�Po�#Jͨ��ɝ8�ހ �^\�<�`��B5>`���\}�`�R/Y�<IOE='���k�F�-ቂoT�<A�`p���F�,�bkAR�<)�fܲ��Ĺ�2]yĽ�FÃX�<�%>�Υy@��+�!�HR�<��]�g	��B�*W8:���E�<����U��m�3#�88t+�D�<a#���R����M� 
�k�<�7⎰s}�؊qn��NJ�K%/d�<Q��´RP8B�A�l��hC壀v�<�f�,�=S�eض��d��K�<���X޶�BrI���
�kQc�O�<CC�E��3�+N�#T� [��N�<�PLō@"��u鈺|��rU�M�<aP��&B�=���7s�4�A@~�<�B:i��Y�
3~H���E�}�<�Ń[��iJ�G��-K`͢��a�<ɂ��0(%n<��̋Q�H�҇G�<9�I�8�V��$܏s �Q�͋@�<���F�&���۴��vǘT���z�<Q���%?,���j�g�d��Nq�<�eL۞1
�I��%�3<�BĘ� �l�<�Am�8!��Aa�ݱ��L�DCP�<yo�"4 �a���\nౘ��Dt�<��D8A�DTz�lI�]��8xv��q�<�@� +�����}8}�-@V�<ᖠ��҅{4mS4jH�"��]O�<9�æ��p�"L�) ����taD�<� �,��@��Us~���Iѹb|Pl�"O�'�9�����?:yH�"Ovx�.Rc��:7��aB���"O~��u�(J.̭х�6нE"O*�����yHƌ8��Es�����"O֌ӣg���@<pRdB�#�!Q�"Oܘ
��\�����CC/5�N�j@"OX�馊h��@Pg�دd�.���"O��"pG,b��}��F^0W�"�P"O�u$ܸ
1���ԠA���b4"OH�:5�2���ؤNۨz�L��"O<��H̟Ѱ�K��z�Y�1"O����`2��v�]�#g�H8"O� ���Ӹ(��a�A(�
P���"O`�����
L��AV� �l�\d��"OnMz��^XYi�
7T!F���"O��'�D�L9�N\�W!(�{�"O2UZ�O@�H`���ߣd����"O���ϜhA64S��zh�)"O�@�բ��x�ة"�kA��2"O6<� K�{:�얎M,�P""O�zQ�ߟ)���Z�,�I"�q�"O�!1cJ�z,��ySKO�:X��"O�|P,�j��:5�R�>��kt"O<H����Xx2]�� R�12bl�"O����[ /�n�����(�T��"O�к�GT�4?�49E���bƸܙ7"Ob=�PDQ?����'�?,Z�8c�"Oȸ��fݽ��]���Y�(Zz�P"Oܠ�'Ȣ��D���p⼛�"OƱ�Ů�)<��c��ޝ+M�t��"O�P��h�VV��A�{����"Ox����t��c��&+���"O,\y�$��P�@�\#3l�Q"O4�rB���~�������r�V��a"O�`�E��0-�4���-_�ze�r"O�r'^Ac�UP��ՓU�����"O�A�T"� $(�b8H�F�+c"O���v�I����`I���p6"O4�S���)��h��8A�X��"O>}곥O qFA�۲Pj��YV"O��Ɗ��2w�����1b3^la�"O�9fe�0�Iy+�E��]҇"OP�q ��)kq�׽�z�{�"O�Xk�M�6n
�M �܂g��@�"O�,�U��E@,e�3��M�P��T"O�L��&�l����S�\��<��"O��3a/и(ؐ��֣�+7�^�+#"O,j�[�g$�arFm_��H[�"Op�Kw#�S>m��+_�,�4��"O���,K^��s� 5 ҄�@q"O���T�4Y�-�JT�}����"O���3�i:g��88�`=�""Ot	�2P;�r�Ic���dI�3"O�y	C&��
R��`@KB��� "O�m)�Î{ �����KEn(Iq�"O]f8&��E�M�(?�(0"O�1b��c�"x�$k@<r���2"O���g�Y��yKc�Ӈ[�4���"O�Q`->���BHG�RU���4"ON��D��ir�t�Cj�-�#"O�y!苋���A���@Pa%"O�@[��J?Z_t�aa�<
L6!��"O �a�ìc�>��a�>5�6"O� dLrW��
j�^P(��M#v�a"Ot��KV�R�Y�c�0r��qC"O&�b�G��9J8�vK�~���A"O�œQ-�K���k�;N>�P`"O
U��6R-�
��.����"O��F!�!Xc&l��Ǆ\x�P�"Otxi�^�os�ћ��_�[D"=�'"O�})��H�y1��TP�|ѹ�"O�y/�>3�64�GU${�r�A "ONu�n�u��t�!n���g"O��!B�B0*d`�@�,}b5��"O���NV�r�#`��5U�` �b"OZ��E2g�XCS�ѷ�P(�"OP���YJ�n	�΀+3�N�0Q"O��içK<`46Eڣ-��� �"O�C��� [F�h%f�4o^@�j�"O6�p楈�.�L��5E�x�"O�����9-b��҅���� 0"O9�^�>Nԭ2�#ՑhV��b`"Ol� "�2nl��x2�F�vX���G"O�983-���N��5�U�%>\�j%"O��,�1oa�ٱ)	
&M��8�"O�dkwd�
i �l+'�׉N3�-��"O���&q~��
��#S�*9`�"ONX�J@�ra��ޡP�5�"O|���� Z,e�e쉥Q;j�Z�"O�hJ����u��
�6()�-�"OP��(�|��	h(@'Sr���"OP�5G^)H �Ф'o:�"O�p3B`4qp�����1
dP��"O��8v*��8�i����I� � "O�u:���g����P��U���S"O��	;O���z�e� �A�r"OΉ "��iF-d��`0Á"O"��$�?h��B1e���DѶ"O�u�ɑ0#��=7�A�#�2��"Oބ��Pr���	jj �
D"O(Z5�'$��ԳT�\�Isx�"O*=H��_ l��a�LG� `����"O���!ǟ�0X�0HC�K�a!6)��"O�kaIG�w��KK �PB�H�"Of��R��+�hҕ�ޑ[��p"Ob���.[Ta�Y���/q�t��"OLձ��'ºu�DVg]`�R�"O�Y�
?��)�ul0����"O8� �!Qq��8цk�)��Y;0"OL!+$X�2��$���C$&(�D�4"O��� O�Z��u;e���0 C"O�횤��O�)0���uj���"O���y��A��:v K`�2�y�
�!����%o_�~d�"��;�yb�P�y��(����6�`�n�)�y�k �(pb0�0�"z<��(ؤ�yBH��vJ��e�]=w�T!�W����� ����i�-yߐh��a�Ux�މf�)%��F����ȓT��)��#u���0������A�6�۽�6E��K�i�6���*n���W(�
h��T�+;n!4Մ�@��U ��qZ��J�MG�b�h�ȓZ(�`r��'4�$�
�̰C]�p��X *�X%oP�;2���4N�a�$Ԅ�%�:Y����+G�D<��!�&l���� "]򂀖�5*t����!A���S�? T���e�`��uK��_4`m~Yː"O.գ"F�,�JXW�f���!"O�1в�
����kG�wb�8��"OZ�b�06�Ή���I�Y�DlA�"O�%Z�cJ���{3`�b���"O,9ʳ#\%�Jc��:�	��"O�3�m#l�Y�"*�6 ��S�"O�Y�&,�.'zhĊ�i;7`��b"Ov���-ϒ]Qn,A�*V�*	rP"O��')U2�.AXfJ�6@�4"O搚�ɐ&f��J��:��e��"O����A1~����t�^�6�h�1"OL�"@�;:�ȍ���[>�yPC"OڀKj_!/�|�bH��(�00"OL �fK @.PD�y�r�b"O��c�RL��gŀt��LK�"O�R�)�(�0�b�рv�@�"O�x��׻k���#c^�D�6��"O�@@I��r�
�J�K�~R>�"OD�!�X8d���㉊L�̛"O�X�&ֲ7�I8o��NgN��U"O�ꁊ�� e��_8}�0�(�"O� �P�ՑDR*9R��Z�+ຑP�"OPL��/gvz�1dR��t���"O1��MA�6��2ď���k�"O�|��	68w��H��*�� P"O����P��@��	�/�Ȼp"O&���   �   2   Ĵ���	��Zl���5Y���dC}"�ײK*<ac�ʄ��iZ�Fm��x"�I�
=�6�K;F�Hi2q��\q��X$��=D.,$Kd��-T"lZ�M[�O�	��.H-^ 9�ɻJ�z������W�H� �^�Kӯ�
����vN^6�p�_��s�-]�~��!8J����l�-gf��[pE�(B���A�ixA�Aѳ0?�	%F�|�r��C�]�I.?���A.�"��	"[��Ԣ��G!A���f��?A:j4��/��OJ�&��9+���%>�k%�:|y�x�E�FU ��3񋅭O0*1��NG��2X���]�D�_Z�]9��Ob��0̈́*4�1��kF�plj�:����L
�q&fx�]�D���x�#J~2���r�!���2�@�K4�G�-h��!���(�A��!�eq�Q�Y� I.t��S��9fh<�:��H|-%�80�N����&��Җ�ͣ-^4L�O}в�O�/e������� B��|�Є��\�H/�I�'s捙�K�?e$�d�<q��/Bo�a�d��A���u�D��rO^�H�q���j�y��Jx�D��a֦���n�5_b����e��Y�0�9'�:?	�������S��ly�	�X�"L��P%��>�i"�1O꼸.����� V`�'���r�<��8h�H�.�~s�27FD T�l$�PЄ��PJ8yˠ��Q�IA����x�4z'c�lF�I�♐)�"�ʴ>AtiX>��$�4�!�@���O��E
[�3+էQS�u�'��k�l��<�%�'�*Zq�L+�~�Cw�l ��2dfyy�ŁC���$�8���Tm�ϖ��S+�@��+���J��IQ��X���4d]�����Fh�O�0B$��)3���k�>i�U[��v�2#�O���r�'o�(
ɼA�j)�$b�]?����n�L���N>����3Z�,��<���9\X��0�dK�Ha�	�$e�+O��l��'�8��@ ����,�yN�.�@��MXp�i�e���y�j�Wvi��H�A�D#bќ�ymĂ�2|�I�55(ٛҦ�y"�v�l�F�V���b��)�y2�[:� �:���<}zH���N �y�
$7
�D��f�w�ډ �eڥ�y��IX��{�D'g�]���G��y⬙Q�4I�r�J�M����1j�3�y"+;˸�R��N>L��     ~  �    /*  �1  �;  �A  H  �N  �T  [  Da  �g  �m  t  Qz  ��  ҆  �  Y�  ��  ߟ  #�  ��  Ӳ  �  b�  �  W�  ��  ��  9�  ��  ��  �  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6�F{��'O��V���&�;�+0:��x	�'%��"J�[�]�R�K2r��"
�'Oe#W烹�R}aC��z��
�'��;��7�������L	�'�:<*b&K"4����M����9	�'نx!c̓>�D �,ݻ2zX�R�'��@ �F�9<�m�7I�"+�a�'ր����>��Y�
�%&���'��0��3L�r5��M/� HJ�'U����J08fx����I$p:<���"�����" 2�����bh.�O�l�<�#	L�|X��:M��u�F��d�<I���1;~�jd� "�� +�_�<���\�r������2!�ځk]y�'���O�#<QT	��L�`T*�.@��q@�W�<�#ǘvʈyt�ƫ�>ii�C�x���=q�$�?z������X'�d���d�p8���?I�4P�n�q���2.�p1�N��<!��ȓN��vg�L�i2(
� ��ņȓ9!�T�p�"�R8��@�p�t��Yİ�]�8 ��u+Њd v �'"�6�HF��O�]+4�s}�)T�5)�P�"O��6�X�rR�z5/2��ȵ�D�R؞L�!n��N�������[�L��vd?D��t�ɽ:��C�%_�6��@�/D�X���[vd@ȢiX�K����)D�� B� �i	Q���Yu���wѬ�%"O\����ۘL��h��H�c�
`�"O&�i���2�� )�(7}N|��"Oj=ȥ�Қw�L|�v�ؽW/�m˥"O�52���w!��JĦ;�ܱ����s���IR�8w���1*�Z����h�� �$هēm���׀v=x9j��F�(B����OܓM><�iV�B+1NF��b��.1�ȓpo�m�3�S���1F`Ԡ���?a5훦���ÎF-<z��"`�c�<I%I�r�
����'��t�Q��X�<Y2�6K^���r�����,y�D�ȓm(�{�%��s|������V��M��_<�'��0v�#��":��3&�g���#��x2d�(C4�4�g=/������P��yb���H����&\��|3 ��+�yR�0��i���	$Q�z�����'\OP��E��z�!򤗴-f�d[�Q�C0�r�X�i�!�DG0E��h�Rkۭo8:]�Ɇo�!�dA2�$x��ɁK���脊h�!�7y� ��#9��٪%�O G��|B�x��U�Gx���֝pȺ<s���yB�{F��X��f��105.���'�ў��M���t�N�W�0 �ॹ��'���|pa�!Vs�VE;q'X�x�(�Dzr�'����j�h�1�C��W�2	�'Cn��#�I6Uu�q�6e��}�xY��'>2)S�87L�e*!oT,|����'k0PC$�*�D1�JˡF�(�h�'��x��Ȇ�]�<�:�'Ӿ,X��9���'u�)��4��Iv��^x"�'G`�����^;l@�� ݾD
�'j�%��%a9��~Z����d%�S�T!A&J���i�K�8J���r���y�+Y� ��7,z�X�-�=��{�	O+:�I�o�f�D�R#Z��y��Ar�кQK0W
^�h1���y��B/q0aص�/I���j�����yr��06���@��GR�z��I��~��'�D�C'oI�Gz1�O�+G�����'�丸�#)u����G��E$`	2�'��̀j�!�,d!�'��6<l���'4��KA�7�|��� �5��'�5��K�P�h�NڂI�`�q�'g�0+��0WSpm���D9��R�'�`4��L0i� �0���K�'��$P��M�uJU��,a���'/���1��H;��1��?�HlP�'�n�q���7gOn�U�fQxe��'����9sf�X��̄J�}�'YЬٕ���Q:�]��a�BFP��' ��d
9H"P�2!�>|q�	�'�^]jk#^ӂ0h)rԘ
�'��� �A�HXb  �ӭZ��
�'�,�/e�6�AE�8]'J���s�<�' ̐d��yӥI�N�"h:,Dl�<Q�i�K�$2��B$X�X��	P�<�Q�۷|�j$sfHA�1a���-�R�<��?%��	@��N,v�
�I@S�<��-�[��,S�mװ/�-�2kP�<I�n�/�ƴ;�I��7��9��a�<��!)���g��r-ѓ�]�<���^�[�R��a��c(9�"n s�<�D'C69����J޴D��"�̏o�<� �3O"h�
 �s��A�6"O�= �gN5,v�X�t	���Y�V"O�U��i�6J
�j���{a.�ȗ"O����d�<C��i�R�*M���*""Oj%�$ǃ6's�$Ǎ��v�$8�"O ���ݏѲ�j�Y�݊Exw"O %aRhԌx�g��E(����"OH�@�v�� Q�Z.	"$��"O�x`ïI�]^v,� ��Ece"Oz���Ow��zC��X�hԨ"O�ᵆ�`}Ҵ�aoK��bu�F"Oʕ!�K�� E��Mک4��A�"Ol� ��]+5h�%���a��x�T"O"�i'=/���Q�9y�|ʦ"O��q�	��3\Py�'鉶+kအ"Oxx����$���(Ѻ3���V"Otp�"ɺ�$A��H�1% �ir"O��h1	H�U5��G_�k@�G"O��ҭX�kf�` ������"O�,���,��x2dEƹ�J�Xs"O��zWB\��8��sm��Th!"OF�[`h�G7.ܚ���}���� "OJe V�[*L������0h��	��"Oj�����x���(4��4� �(f"OT(�B��$�Z�S�{��Á"Op�P7|���!F 9){��"O0�!4��H +�dߒUz�p"O��@rcÒF����݄7�P�9"O�a�n����As�()hf "O:PK�+ݚ_�ب�� �kH��q�"OnEʔ�i��d�2(� �� 0!"O$�˦G�=4����	swpE� "O��� �Zl����V�X�\�[t"O<�gZF�p���.ߵ��Q�"O��4)��8*�� ��< Xl "O��z �[-=��か�3_�T��S"O$-���E+Oru�$�>g��Л""O ����}�0��B3RK��;s"O��9A��P�FX:�$~��S�"O�r��ǩ"R��w)4/�Rl��"O��X�e� ? �#"ɑ�e 歡c"O�A�c�E(����׮r��"Oƙ#e��
m�f,9��6�d��A"OFe+�ۜS�ݓ7�L$H�LY�"O�]�h���T���S
�d��"O����*	冘Y�ט���"O����+ �i��N<τ��g"O� h���.�(I�a��!�b�{�"OJ��`�דO��J�-�3J�e�"O��@D��2&}�t���� o��6"O:Ѹ�o�6 �Q��j.}�"O��ɋ�, +��Y�;�pS�"O��r��%�ֈZ5�Y9�8�"O����ߓr����,��"O>�7L�&v�裧⑆�� q�"OD��ClX�V�38�����"O���FX�i[֍2� joƝY�"O���gR��м�g�ٓ�Z�"O`y�1�ճ'�͈W%(�\#�"O�e��(V�H-f�kq��G�x��T"O�����
�c�JY�!��� ��"O�1{��	�0�Wǘ(���!f"O�93�-1^x@�EW[0��r"O"�b�e!t�8�0�DN�i4��"O� ���`
_<]�g�F�!��T��"O���&�ػe$��r��f��5I�"O^� ��/f�Y��į��T"O>L���A�z�i3�˓A��)JD"OF-���81Ƕ�е[�G�z%�F�'��'���'���'���'��',�-`�e܁,��(��V-H�p��'z��'�R�'e��'��'3�'|j8YDҴR���{��ڻu,:�0��'K2�'�R�'{��'�R�';b�'x%z��E<�� Ў�}����e�'���'��'�2�'���'���'�!ddl���2��X���'=�'���'���'R�'��'3�}*cv�¤:�� T{DP��'/��'��'���'�r�'q2�'!��{2h��M����ċ�
��;s�'�b�'t��'���'���'���'�`�t�&=y�	]򬁙'�b�'���'���'���'��'�Z��E�+Pt����ʍA�4�X0�'���'tr�'4"�'���'���'����W��a�H�@�F$������'*r�'s�'���'���'�r�'$��RC�%0���mӭ�Ԩxe�'K��'���'���'��'���'E���Qf��4N�,�S�6OJ�'�'z2�'�������'X2�'E��'t `ʐh��a�����K�3
�i��'���'���'2�'�R�kӔ�$�Oh���,G܊ :1� @��%�Jñ����O�S�g~��~�d�8��I�{�
�(5A׵i��T��K@?�	�M;���y"�e��آ��*pB�@V�r�C�ͦ!��%)�Fl	��:?c�ޟl�"�e�?��c�:Sڮ�[p��,F�J�3�d���'��T�lG�4CJ?_*Q:�_�:���ȁ䝊[�6�M�b�1Od�?	����c��D�9�y�k��L�H2ď&i��g�
�	v}���Ǌ�]���'��tġ�L�<��T�5�B�ћ'6�����=w3����i>��	!�LĲ0�6.ę�A�;���	lyr�|2�f��qb�Dά)�����ןU݂e0"�O�a*��܂�Ov�l��M��'���AB��`��ώI��q�Go�����|;�B͸S)*��|� ̦P/��x��z��=��@�!k4-�4�	tLm�/Oʓ�?E��'-Z}`A!Z�C�12f��uz���'6�7�Ǿn���9�M���O"��i5��b��%N˘nB��'�x7�̦��	�Q��9�G�>?�e�4?���#A�D�\T�0��	]�"��{�HxsF�[�J��Y�Ր1���4�3�d����G%������b���!�4I��Ra���G�<0�Ā��2ikPDJ��� �H�G��Q����i�DJ 
	T�l��E���B���ǝ�2��I��bƦD'8,��d�: $	�0ː9EB��+7�'GS�������T)3egͰhh��uf�04&T��(�$������؟k��r!�òef(��Nե%vr8���na�f�'?��'��TB,?�D��TX=����8Bn��!M}��'�l�c�����'�!B��8�b��ɂ�B�,�)�4\��["�i%��'x��O��O��^�$����![`@�Ys��'���mZ40�L��?)�g̓�?9��[��$�2y
�(K�aG�R�6�'��'m8풰-*�4��d�O$��ě�I]�P�c��in�tbC&EԦU�	ڟ���I��������d>�d�O���i"q<��&�,b=�NŦ9������M<Q���?�M>�19�IR�ҩ��yw��4�4l�;�#�џ���ğP�	����ORf�-,\�l0� \*F�t��"�*y��ܸBJ)�d�O����O�O���� �媘�='b0i�o�!@�H���O��$�O�˓�=�5�r�M��C�0�R�E�K�T�#�d�On�O�D�O�T�P�$���"w��(1��)_\����>A��?������?%.��$>�9�	����D��L��rCk��M����?�N>���;Ҫ��|nZ3B��Q�Ip�"�g�ߝe8�6��O���<��I�UX�O��OS�0�3�	�'����P+���qp�)��OP��R
/���O@�D4�$nל&�0� *��/�<���U0�M���?1�mD$a�探~j���1��\�6��#���C�YvM0�e�>��-#�L��R��ē_�t�ەB�
X�ϖ�D��o�&�Ld�۴�?���?���x����c��6�$��F�v�}�����6Վk���d�Ov�$�O*��|�-���s���]��Z��	fM�x�Ƌ�˦����x�	�[�fU���)4}���<~�TU8c\`���
�N� ���?q�J-��'���O����K>Xx��e`�i�����i�.Ɛ��I���)4�I0tD��:��H�IZڕp4G�LƖy:�4�?a��� ���?���?a.OĥB$�ĮOC���Sc��~����ҹ{m��&������4��qy��'�Rd�rcP���dI�m?���F��
4�
l*��'��ݟ�I؟�')Q9��`>��� � �RQ2P��;nbRp��>y���?	K>q-O�p�Tf�O( ��֖e�$�iR/V1zκ�0���z}�'��'�c2�e1N|����Z�J\27%N'���P�ΪE/�F�'��T�(�I��LI��؟��O�H��Ӿ�.5KVk	!KO�)��HX7�M����?),OI��a�ӟ|�s��� �C
��P5%M�If�(��g� ��?9��e:Mx�����O����� �0�� ��1�|m�&(I�YV.D;�e�!}��~5�c�&$��g�/eZUk�FU�hl��tl>�t���u�v��è�Lq�ł֋7�ԍ
�̆�>�X�Y0b2U0P͘��߭z�4��
S�^ѳD�Ӂ#֤m�ρh�.��5�<��}r��P��ak\&fO������"}�4���H\��������2�U��dp��h[��^՘��N�V��� \Oz1S��ړNL���ak����?A��?���d���O�E����-�$��d.5L���Ӄ����P:0N��H����e�ҧ��)^Av��3�y���%W�E���C��;��K�f`�Y��E�U�Bq95L8e�f k�OK�<E'�3��X�$�`H>�q��Un�I&CX���K؞4�j�l�l�a��~��H:��1D���#ҽ\;֭z�Mà<���H@�/�HO��>��A^��Pn5"��ѱ��א,��)�v*�FU�I՟���Ɵ #���|�	�|���;1���.F�TYr6鄎(
v�Q0k��OE6uk7n�T��0�AF��1�ڢ<!1+��O+v�Z4�皤'�8��Ή�=F��q��:o�l�3Qh�
#���� ����(Od��2�'�h7��v�v��7O\	Cf�Ĉ��R	U�!��0(X<�#��+B�"d��cI.1!���<���	ؿHx��C�)ߊj�$Ц'���d[���$�O��'lYp�p�*�"���J;`bp4 �HL�?���?�VB	�2����Sl���Q��
&S���C���F_*%$�Z+2�iA&g�2l�uDy��r;��r'���#@r�9Ea�\������\�`��%Pp$%^ ��
�Z��eN���'X����`\��jK ��R>i� �?���ĦϠ=N%ˤA��M��i+������	�I����A|��A��̈́�	�Mñ�i7RӉBc����ǉ!��͊׌ܥDmD7M�����l���Iџ��� |��	�4������K������]�6��lY�遅o���)s��3�<9�@���i"��OX�0 �{�$9h�/�*c���҆��2����ĭ�&��uim�=3j_�L�q����0%8]�#CEb�}�I���C�'�B6mayJ~2�'��TvH�Hf*Ը��m��K��!�:F��a)����#w�A8��._��L*���z}Bk�%T��K��/�Z�s�CM�R�'��E�bJ�.e5"�'d��'�X�]Ο|��!��ب&#Z� ���[�	�S���	��F�qQF�jC�ʦv��Hfi�?Fz�O��K�����33=�Dc��$�r���C]�-�kˈ��~1H&��?=���3�ɓ9���3��#y�������;d�j�I8]���K��e[޴��'ϖ�'3Gh�Ja9Q��! � &�0��ȓ|��)P�k�$k�B8����iph`2��I>�M[���D���n��k9x=���GTMa�������ݟ���П������	�|Z"f�����u�J���,_��pڳE��������
�Tp"E-E	o�K�'�������ݞ0���b��<鄈�,d"�� ��B�ll��"O��� *��B0yaf��RS��L�<�'Q�t����kL)>`pJ����<�p�dӊsdm�ş��	Z����@줲�B)*�D���X���'"b�'�0�DjH�,jJt�q�):4ԠK'M��O�T�]�T��5J5�˅Qo�I�0?�(OM�W��c�X�;F��bO^��3�Ԥz/��5DA Ȳ��
-O��8���U��(OT�Y��'��>})�ML0.p8QIT#) �iԯ1D��[��K�I���e�2�:�x �0?��4��i&�T����o��&x�j�l�Bk�6�M���?�/���	ua�O(���O�A`@�#��,a`O�]�0�zV���3j<8��	�0��d��(O�g06�0s���:��b>�� �8b:�Z��֮KH)%H�'q],�� .2�(�����f�V�o���m}���ي��X �X�d
�A���K�-[��%����S��?��)v?�̻�N��O]b�i�]�<	0OP�',E��:_�������V��?A�i>��(~������RP�p������Iڟ�AoX:�V��	�\��ş�Xwv�wE��rv��P(x�S��W��@"��]�����7?e��Xf�͊���bA�<a���������,v�#A�Ҕf��� 4x���(ό5����wҟh����8�'m�M偖#pF��[�*�$x�j��'���d�a{B�Hv�&�(�+�*N�]zv�<�x"�'On�� �|4�Y���Ac��� 9�S�O� ��2�f��9�bĴ8̞]�W��������Ov�$�O~���-2�����O��S4�:�P-�9U!���DL����$��y��-<�O8�F�����	#3�%(��ꕇ(&	��/�x�a|R�?�?1�i`	C���8I��A�)��Q{gO7�$�O���4�)��	�AöJI�X��$u�<iB���R���.]p�U	U�<�U��'
��@�,j�B���O˧2��
@服o�f���"��':bY
V�A��?����?�b�>S����C�T��MT�ɼ;)�|�W��u�CB �/x��$��h��u�d�򄈝w���Ja'�Oʛ6�#Z����G&� �ᩐ�ט@�Ċ�,|n�k��1FA��٦i3ڴ�?.��\���PE�|���L�H�����Ot�"~�6֮�R�
�-oLU���x�D�']ў擁�ēcM��{a�!"���a�؎V�8�Y2���/��?9�����inN���ON�D��'{�0�4��?RJ`@��!�4MY��qa�O�b��g�'�� ��%�-*熅��eժZB�(HRƻO<�"~�I>8��l�rώ83�V�qv�RZ���s�ǟd"K>E��/��*&j�8�t�ɴ��(���ȓ4���!�%�ZY�ͻ���^���Dx"�)�S��E�C<���K	O����%@��'`��&�@�C�'\�'�֝���ݑ! ~�j���=ݢa4&PU0�F�w��X�P@Хcd�T `�?)*�@�5�1Od(�B�+�M���j�JX0E̋�y�R@�*�~-
��S��i2���8�yE�O]���ӷB-:�h�υ1�~؜�?���'����."2�\"�-��Z^�(��'RnM =i��� #��3v��b�"�W(#=�'�hO��䍚�O�u#�d��zp��"OR	�#��?xY�r�H�jTT�"O��R�6����ǘ5I"��2"O��a�I3�*"�W�=�8Ȁ"O�u2E�ЈR5�`
L�j%nx�"O�Y������A�ѧ%X��&"O��"�)��[�(qW�/�,QT"O���7��'/m����ٴO��HCu"O(�d���*R  �,�+�R�$"O����I]�\h�
�� O���2"O4y� ���+����IH��ĥ6"O֍1s	Qf�0p��H����"O����� �:�$4#�ŗ ��݁&"Oqrt'�9ƨ��pܰ�X6"O�Ԑ�����aIZa��4@�ym� Zh���f��l�� P��y��ĺn�t��'��&r��r��>�y҈�)*mѐ�n�Yv @���yk VHl�b��H\)�푰�y�G������ǋ�
@��9�K���yb��U[�ذ�L��:�<e�t̚�y��;.v�c�o 0�� ��Q#�y�l�7����#��yf��'�^��yB� 4\�jQ)B�_/� �xw+���y��X9 ����&�t방熑��yb�O/E��A!�#�=p�����a"�y���)-�<�f�W�SzW��yr�F; I ��#џ?h�U�C)�.�y�H�&5XJQ�3�Ɖ6�dܓCgL �yB���a[m"e�A�AM��p3��5�y�̔�����̳g,�����.�yR`��o��C�%�?w���Uï�yb �(��PCS�$��ी���y��	�WB�x`��tƂ��y�L�6��FС	��<i�D��y��W�< �H��D�D(�ǧ�#�~@U�,��O�>�{�X�_�,�R�&�:dFf�h��"D�șю�2��铀�ڻEtD��M!?�#	�7����3^� �3 ρD@�L$"G/ia~����AE���IA6h��y�p`��J?������	�yb�Ъw��mC3!XE_���GA���OLX����(��P��Po�iB2�˨���y�"O|- �%�� *��qcm@�]�Q8d��"@�b����;wVӧ�^���t�b�5�Q-:��JX�r���1�&�4�U �6y�|�C莆�-�R鈼Z;\˓{��0i�`[�crj�r1�]>q��DyRMN|*��1�<%ʴ+�Ç�0<�W�ŭ��(�T�M�Xܾ�� +���@a[�ì��TCJ�(2i��H��E�0����=�O�a�#ϪRD
`M�t�$$���"���Wh
HJR%�L���ZS�4�V�5�U$@F!���Z][
��2"O� �D�"%�0L8�C"ċ~���v�X�iRB�ňK����)ԫ>P��r:��x�ԏ݈|�Z	BA���ar0�$O�y�ЧD9TZ��� �l=����#ы��	
]�I8qiG�W��*�R+x�Q�<�BP�{����#HPK �1*-O:�i���<
�Z ��1��q" ��U�@	� ���x��ɢ�&;WaY���K�����-,Z�B��	�q	�@�o_zB��'c���Ϟht�#��]�<hX=�=�'X�������x*du���d`ńȓx:��;�&E9e_�u؀�ڧIh���k˿S�ҕP��*�)ڄ�ʇ	�λ(9Z��T�IP���V�{�4���D�(8HV����!�d��_�}Ru�S~B��8������gIj��3*�A�'f�z���3�6lkg�*I�T�9	Ó]���Z�iK[HTH���9S1�<�s!�=J���Q8)`���Fϫx��aۧ�
=A���Ֆ}Ft��Ƙ,.�Usr�P'/����\ͩ��ԁ�&�ٴÐ�qO�鄀x��A��
�	 q��r!AW$!�Ğ�#�9jeJ�*G(q�@��/��hm�'m̨!P�E�d6�D�C'rt }s�wT�LJ�N�5�TI�����Z�P���'ԬMH���=�VU�$�Y1r��y�W$�����eE�N� ���gy���lK��R�F��h����5/b(���%�MX����Pz�jC�[&��0�F�X'b�M�$ �_}2��1�d��2��H `e�/[�0�HN�Q�'�~���I�S�gx��#OB�f�� y��օX�t�b��)W̄C�/*p��ǐ�|5��g׊��Oj���U;Bl�A�<��O�S)A�>-9�NI�E U;��ÿCZ���D�p|lE�F92�hk�	db� �#�U��h�+�v1��O?7�6(LT�#�`���P� �c��@c�*�D�ɢX,���i��#��Qe�Q$��)��ɐ�a�tS�1BꙄ��b `@���[U���&Ȉ@��5ܨF�����P�X�����Ob�K�@��;��R`�Y'�D�*�n>D��b��/�N�ǅ�!; e���lӒ���	>v�B֟�`����=�M���|��1�N�FY@'D�A��(��%�O���!j<28��a��\�>�k/������~���h�3,ih�1C-����'6T�5ʈ}�e*��]�2��]x����Ɯ!�'C1f{���[*���^t�-�t�A�]��Y��bW[0,0�E/ɒ���A��E��d�HX=�$Y%�d�X�10%�>�e/�*h�!A�B��iɲs�L?��'��Hc��`�A"�E9�X�uH֕V�rB䉅=��i�SM� *�����¦l�nY��Ŏ�xU���'��d���)̛��Uڐ��ͼ��"L�F�,�����1:�-��G؟`�t	U����q�J�~�"&�8	k�"�$�~b�O��� �A� P� Fo�%+]�����M:!��,��`P$ n�.H�\џ��ޣ\�n��6�����.�0#�@��0[�8 tH�-bm�4��DѦb#�@ ����g�����5|��%�%�3IX4�+x��I J�O�iz�$ˡ��P�韴�q"���ɇ0F��M��fŻpk&d{��C�<���D'�P(K�'��\��ݜ{L%s�h� �5�=�O�<H�&P��y'��������K3rh���L��x"���S>��g�4Šl0��q����N�@�d��]bdtCuŗ�<Q⍃��(�I9]�|�r��!�� ��]����$�S�~	K�o�0�頰���)��Za��*���c�˱8�(�À�UV��d}f���DXq��dN\�HH�p�k߃,����e1�ǞGX�J#�a����@�2#�!K '�#G�)P�,d!��?��i�ӨǏ*0N�1��B�b}��GA��xz���T>��gDY�E��5~���uč���`HP�C�	'u����ǭ_�t��$g&�.��a#\�:��$K�Đ��Pb6U�p�'��'��m��,	�3x�B�WMH�Ǔdx��O���1���M=zЕg�N�pf���<�R]��Qx��@��ɩJCڅ��b�wrvk�J7�_�t9;Q��6����6J�g�P=¥ճ;�C�IUf��3@��?z0M�N�\���!J���?E�ԢG f:L�V� #B߂�*C(�yZ5t)� �_���Z7B�?:(�C��3ߜ1�c-[�
An�j�;��C�I�9W���U�ל>I^EP���;2nDB䉟p���XfE��O�&ՋUC�:�RC�ɢq~���/\����Z�C�	�L��{����J�<����I`�C�)� ~�ӑ�9?����
0��`�p"OpX��� )�xV !�Zˣ"Of	�5�L0���D� �g��I��"O�,R֦ ��M�WH�?}���"O^���D,8����P'xF4���"O��bƚk
�!U�O�'ڠݘ�"O��9�/M`3:��gES2�(��"O8}z���3���Ig�=v "��q"O���!k�X%v��c��L �Q��"OBC�H]"�3!�P�d�5��"O�d��b�4Ę��&�R.��tSS"O������-z��3���k%4a�C"O�<ڵ@I���s�Y],}�a"OR�e&��x����	41a��s�"O���1ၗo��5�rO�WY�}z!"O�d�t�Q�t��T��.����"O��1I��t� wχ5a�v}{"O�!���S�U���L�3�2�f"O����?4+65�����8�"O���q$ަQ���Z%N8i��`"O� y�" 1�d���6&�Ę��"O�`;�^64�Ș���8�TQ��"OX�7
���> @dǃ|�b�zR"O����M�^a�,df�Q��h��"O�*"�?,D��D�y6���"O䑹���?��BP�˭9Pt)�"O�����Z�����@J�� ��Dڦ"Ob�� K�@���p�)ވd�Ԣ�"O~U!�����l��oƧ?�x���"O��X���}$�����.��"Oj�p�dG�T��D*'���Dº��"Oz,����Հ��ڲ@�
8B�"OX!�# ���R��-��)b"O���J�6�E���
D��I�"O0�bC��=�Z�vƁ�~�9B4"OB����ȝ\q:�E&^*Q��]B�"O��ᣀG-���`o�Lk�lH�"O�}[���u��J%ܑ~-�1�"O�BÖ�)�b �� p��r"O�<�ŗ�7,Pغ`��2g� �k$"O���{�Z�1"`[4wʺ�!"O�� �`ɐ���b�A�p��I"O*ՠȒQrV,��ߘ8�D�z�"O
=�O')̬Kw�"sdy��"Ox@"AaK/p����֧t�8X��"O�KB�ʟi,6����t��|��"O�`���+��X[�4���@"O�-�/F��<a(rC�Az:��&"O�Ұ�Q�@�u"@6L���"OhIj��&z�(��c�R�*���9P"O�SC�ے����f�D��ٺ�"O�T�c㌙|�1 ��(�B�IV"O�ܛ�@ަ+mF�����8�H���"O<��,AP�T����9@i!�"O��"�:(B�`0�.��-��TR"Oʘk�i��ƹ�2��X��ჳ"OI�F�/t@p�k��xi4q)!"O��d���)��� �
ݜ>�V���"O������79K�=5)�%}$A�e"O�1Ң� d_ڜccj
7N�BU"O$�0�T�ɋgf̂Y��� "O��p�i�2E�j�P@@!X��PB"O��UN �ְNG	R�mj�"O<Ax"�9|�xX���)�8�v"O� &��ǤE���3�oP�X�q3"O\���"t�"�#�mțl*���"O����Ƿy^��l���h�"O|IS��(l�|���
Vk�,ѡ"O��*����I��iJ�@����"O��;��M�sh��+2iQ�:����c"O|}s��τ69|x�3J+�\���"O���G�(CFh�F0#�Ѹ"O`=�E»;t��*��W =h$=��"O��QĂ�6���I��,��ر�"O���4' �A��B��M�M �s�"O��zQ-:-���3B]#p�"O��Rg ,ir")�A��!�T��"OM�WEC"If�A[��<R�|�"O��`Pg)&�I��;9���1"OJŠ�f\&_��53!/�-�f\	0"OIC׆�x���6��9�B(��"O
�!Il.��PpK�+�s"Ov�����=���0j�	����&"O�Ѱ�-�N0d;1/�m����'"Of�M4}���#��zAB}��"O u���_�NL�qP!E{,PM��"O����OcB��N �h�"O���#�J:�U�тR�[ʴ�A�"O*=Vf�&ڀ����,��"O6d����{~&�*���/H�֌�q*OV��qFf���2 �Wi�=0�'���Kg/ԏ5�b\�t��O�a*�'�F�3����;U�	�+d7�P
�'Qr�9�BM�K����-2A|��'qb�ۖc֚V�2�c����,�t��'�J0�ש��m�Mz� Y�(p�'�v15��/��b7(*W��H�'c4٢���q��<s+�6B���j�'+���Μ/���"����Y
�'�F�ZTl�7�����J2\��@
�'َ��£&���Qm{mF��	�'����nQ 6��@n��r�:���'�g�0{��E8#��n�TaP�'���!�oB�`�b�!s�${<�Q�'x�����;��� ��s��`��'z����A�t �2b�8(x���'q��s1j�1F
*"D�*�8Պ�'��0���6���ِh� ><$2�'��4K���;p��Vs2y��±�yj�4�̩��c�i^ ��O��y��� ;��6L�m�v&�]��y�H��B��&&ǫy-0
�NɎ�yB)̓=���Cn�d  ��G]��y�i�26��i�Ą!Y�)IDʎ��yr C�G��ȑ1E
ba:|�6%�7�yB�ɶk�Хj�(@4-
6��U�M��yBb�-
lp�eH�!%�:}��Ϙ��yr�Я��x�PL��Nu���4����yb��u�����8C[d������y2 c�:��7 �I,l}�#d��y�O
�Ac��	�
�Iߜ|�%&��Ҙ'�a|��K:�� �c""Y��r���f�<��(�q�<���cB��@M�"j�_�<90�ф|2*�pҠ`HP�/�_�<��(R0��K��D;kt��LX^�<�ǅ���!Z�`�VP��E�]�<�v�#g�xH��A����dK]�<Y��1E.�ġ�Ɔ'�R@���Z�<� 9��)�N��M��Ϝ2�T w"O|e�ׄ{�<͚t�ȡ�M��(5D�X��Ӌ<�֑y6 4�PX�&D��S�'\b�l�� ޼lD@p�&D���+�c�����fF�rl4-?D��BG�*��|h�
H��z�KBn=D��P#M:������)8��M>D�d��O�G�e�T�ć6����;lO�����̏�pT.�k���  Ь$D�QĈ1 ��,���{0vC�)0|Oc���� nr���0QlL!�	1D�xY�.�3����5����`��;D����հ�\�:㈟�95 @���,D��3�LӻTi����K��=���!a��$s�Q��G�`�!XJ$x{�bڿ74P��gO���=Y��D�ZjM��&Ե4�湉r��D0�9�O�e�2!�	{�Q!�_���A��"O"���EW%P1�C���SeD�I�"O2 �w�-K��B����u�0�zD"O���-�p���!����S�"O<hs��[EͶ*0ǋ�m�B��"O���7 �_G̕��&��G�n�v�'���8Wk
�	�4cڝ�''7�y"�Ř&�(����*NY��f�M��0?Y(OȤ�'���C���ʃFI6X�,9�"O�\:v�U�/�����.:W���w�	L�OSx\��@��q0%��#q�IB�'����ʎ�"p2Xb�'mڂQ�
�'����S9u��]� D@:$S�'D����N�"a�0�ˇ"�xtvhq	�'�@[P��;MN�3�⚢H^���'�6��'��02<��ӡf�3L�8��
�'�`���؟`�ei(� -�� ��'f^��BX��0�5�$�nx��'��r��!d�-:�C?R���'��feZ$x��;D���T��y��+2�>eb�!�7(9a��7�y��?{�d���7,"9��G��yR��n��i�	+>�s� ��y��}��]��&	&"Sؤ�5#���y�Hѩ_��ht�Ú�6Ԫw ��y2�
)#��4��E�L�FK��y�� 8 �:�kѽ�:�zEk[��y�e�A�r�)3�B���"4�"�y`�	/���z�
ϸ>e< ��8�y�OΈT,��peƋ;7檬����y"��`��4��ʐ/}�(H���M��y�%q�V���m�r��0)��Y
�yr��	�.�i���A3j�aAM��y���D�@$Y�[25`�Xi�F��y���	4���d�Q�.��)�eޫ�y��G�	�:���Eב$�������#�y2��%?� %J!��p�]k��[��y"Ɲ�P������*Y����%Ν��y¬/?�^������^��T-J��y�LޱJ�.H����C&0!MB���$5�S�OOnY؁Ǔ�7��̀�P��\�
�'*bx�Ć��Ήz���x	�'=�ȗ�؁=��5�D�FR@�Ǔ�HO,]����d�䙛t)F��|"Od�ʒ@�6�l���8_��"O��!�D���-�g\ LV�tH�"O̕@t��i*� @��8��QP"O��Kɶ.@6|�%K$5��A(�"O� *$X�h�	m���`K�r�P�"O�5CP�#s^A3�X Q��y�"Ot�H5�E�v��
"��5~�1��"O�m2��Ҫ_��փ	�e[�\��"O0�$�j������)7E�ተ"O��$�V ���pB�0K6��Se"Oh����7�I��gİ�yf"O<�n`����c�"�h���"OLɃ�ʸ&h����0<���"O��6�_#4���+�[�XD��"O�Y �,��g�&� �h���}�!�Ԯ(��`1�X�\�y�E�!򤞟vHH�Ks	��~i��&�7�!�$�.W�e��8VE��K6u_!�dQ�=�@ݸ�cԒ0��h�E�4P�!�ؙN;8%�fMվ&���j��6�!��)dJ��h�H�;H���
)�>�!�d�^N0���Y�KXQ2����c�!��Ūk�����L�P@�h���!��(qd<��$[6H8���\7�!�d�V� �f�P������u�!�d� vgF%��\=s�(x�!�ݯa-�!��aR30#��1o��c�!�D��<m\q(�C!!,ɒ�K#=!�]�\PBA@�ʉ%t84��͆#G�!�dΰ4�褑� ��Y~�
�ˈ�V�!�U
AԸ��B���[ia���!��بm4�b��V0T���c��j!�$� Zyv�s�a2oD7*�!�$�nR�*flα�Z`Y��նO�!�ד#���(@.Ѷ\b�	�c�u�!�A%\xJ1�P���\ �|ѤX?j�!��F�����H	��I��c�@�!�dQ�६(1�ހ;�E��i$<YS�'�F�g��L�T�W�_;uZ�x��2�l B2C��?&|(n�8�ʔ�ȓv0:pj� ��Sg�v���Y0���Ҫ1��=�d��z�ꁅȓg`�c�鐈it���E��.�Ҽ�ȓ.�<%���|�R7"��M�ȓ �tu��X�\�h�
�|14���?l�)�	Q�[��5��c�"_���ȓW��j�L4���AO��`��	�ȓ��X��	u���r/ה!�PՇȓ���@f�9S�6�1f�8l*��ȓU�^=a�	J�QJM��V7a&l���t �&��<V�ѠAĞ5<���6C��@)�s�q���N�^=�!��;,�l ��@�z��4�Ёk�[��4�r�ZF(C�vqT�q��V;\�(���+
� �A�Y9Nz�=���
�9��X��K�x������uC$�O�3"OHI ��=�~��t�v�X �"O����F�)}��krȅ!>'b��!"O��7�I���r-J�Im� �B"Oz��6G�%5HMsa/H�8�"O��ɇ�ȓQ���풢<�Z��"O������މ�U�C���@A�"O�m�fA�>k�깪���)H�<��"O�r�IY$R�<5Ag�2b�	a"O�1)���o�+���o�rU�waH�<ɅH��oq�M���R�-����D�|�<�W�V�z/��p&�T �r *(P|�<0E�	&�&%����N�F)�уMz�<� :����0N��c�$		��K�"O6��W$�TW
mᓉ�67�9B"O�|u`��=Ei"3�Gg�0 "O�Y�ed�6
blӧY�=���(F"OFEx �l�2����!qg^���"O*�2,B���e�¾Tgd(�"O-v���<�Dge���
�y��L�C�ะ�ۖD���Cw�ї�y⅙4C��y��,��5ᬌs�<�!�[�)��=)$$&4���0��ܩ&!��Ψ@��7K�%A��)z���*}!�D5|�XT�O�XY4�a2���%n!��+g�Qa�Q�`�>=����
V!��#&�x��w�	�U����Y<FJ!�d�AC�a���R�:=@d���'[,!��<#&¢	�Щ���!�D��%odM��f�.H���`)�!�m6�yJ�)H/6�4 �Q
�U�!�$��<�
専g	:yX���D1o�!�$*�L諒EǎK��p�2h�+uB!�$U�m�Z�3r������瑎R:!�$kad�pK8���_�:%"O,Db�*�]&v���'�N���cU"On�*taLw@@y��S�;��-i�"O@�+�H؋C5�qY�D�O���B�"Oΰ��L%E_P��ℼs�I1�"O0͉�,��N�����Nh��	2"O֍�$C?��iS���p��"O���ʉ_����OI Jt��h "O��Y�d�	V�8K��\���"O:�i2d
����ס���B �"O$<zU�żJBN)[4a,r��X�F"O�Ej@k��P�DXU��(��1q�"O��y�ȚS�4͚�R!#��
�"OVpXA��ĨF�T�re��U"O�[6,�m�ⴸJԼUY�"Oθq�M����Y���wA�H�"O�-h��1yz�1V��Z]�js"OL��P45|�y�	^�AEp�2"O(���$���B�ʪ=,���"O�(�Ź-����ˈ%
�~��U"O|���ݢ[���+���x�`i�"ON��Cl��V�hb��Z�p��)0G"O�U�^�viܙ�.� ���F"O8 �B
,^�s��?=O���`"O���G�RWC�ay�`��,%��1 "O�]��/B�e�p8c��2���"O���5�W2�4��� >2�@д"O�-���8����bM-*�R��"O\mӥ�ӼQ��}9�!��a\���"OjgDW?
b�`C��S<A��|B�"OHm���5/�,�
����z��-B�"O�ɕ.���
�MF�v0�Z�"O��۰C~����pO�&#a��)B"O�Ѓ�ś#~ܴ3�D�gb�I  "OȚ��5z�������2
D �j�"O��B2+VB�9� �ܦl�v"OXQ{@!I�|9B�9��� x�r"O�Y��(^f�����,O���C"O(��%��O���E��0+�]�"O:�*Ӭܱ'���zE��1��;"O>�L�>S X�tȾf*~���"OZX2�˄�u5<C3��>d�,��"O����L�.��� L#2Yt"O� �P�&OCT	s������"Ov�H�JP�.�=�AO�?�f�Bp"O�aq�j�=KP��Í+Gv=1�"OҀ�d�3mPI	�f
�$6�|5"O� p���R |�T�ن!�(x;G"O|$��ѽ�a{W�C����"O@ �-A�J���R�U+Hӄ"OH|�0��7�Ҍa�Dɚ!�j�i�"OXX��nމ�J���
��aո�6"O������5��t�FC��H�1�s"OL��S�N�(��<��g��~��Da�"OTՀeg\V����ĭF�
�|Y:�"O�A���+�|d�&JH���y�"O4k� m�v@��V	 �F��3"OT���
T�²%�\�&�ZV"OΉ{��u�Z���&=O.��"O䨔kі:�`YB*&>1,T�G"OdPs�E\.s�>=��A���	V�c�<��ǐ�<�|	�pã�ܥ)e�[�<�	�	9J�Z��J%oPi��AT�<� (qz����O:o�v�i*D��b��҉4�F����ˬl&�y�'D��`d��D�B�#5+�t���[�#D�@d���X��%��n�c�=D�PR���3��xb�E�#��}3�0D�@Qd��9����F����.D��9Ω6E��xU�ť]�jl8D�D�uB�6%�i�dKE�b���"D���Iۦ��Ə��`< 
CM5D���B�.)��$a͝�D���2D��y�i˦o�@U����B�����#D�4Q�gʅ>Y�E�w�|��2��"D��P��;d��a��w��Y��?D��b1�I�8���`�.ޮe���c�#D�`Kc�F�8���1pb�A4�"D����5d5p���`�/
.�q�/6D�������X���M��ʶ+6D�hpU'����q����h�)��3D� �gP�2a��	�W++\ VC3D�0���X�*Q�A�1ˊ�Ni�!k&D�T�U�V�7O2%:�c�) ���#�(D�D�èǩn+��+r̟�Nn�Uk�&D��CPh	�G	����m,�]��*O,�P��,�����$<��`�d"OYk �б1��3UιG](v"Ol�;�@�>Ӛ1��ݍ3Ev�!�"O�2P5x�RL�m�J4fJ$"O^�1`!�&Ո����'/,�â"O��H���F���͏�1&z�z�"O�P¤86�dm��m�2&���"O�T{��l`F`H�l�,`z�"O��q� �BZD4��F���� "N�<�'���t�8�a��*<�eh0cK�<�`HT�(���)/�<V�Z��fLP�<i��ɺ��8�I�2���22�Ys�<ŀ	�t���C�A�[5n���Wm�<�b���(�����:k6�4�t(@�<�  ��B��F�8XD�Ճ�,��g��Q��M�8#�iI�`�`�ȓ � ��7 �:x�~�s�K�[r)��C�z�$���;��u�ټ-r�d�ȓn��@΁4����P-�8z�.H���Ģ�G���`�@�E�f�����"P����]-p�`\�so�:����S�? ��	�I�ZxJ��6 �
@^�Y��"O�(���4{b�H�CA\~Ժ3"Oa(�A�+17ll��D�vD({q"O&x�3�u8hqD�Bn�� �"O���u���LJ�I3q̋� `�r"O��� ��9}5Zʣ��A����"OD�Q�C��;����#�R���"O��c��,T,�jQ/�/7ƾT��"O�H�w��JVԀ��� 9H,mYR"Ol]�g�Ӌ>��8Pg(\[@T"O�aʥN�"T���@F�B`�x2"O4���"`��x���M��P�"O��剃c�h�H,��5;V�ؓ"O��jf�=8�e+���#��1�"O�P!Ī �6�	G�}P.��D"Ox �S$����%*4��v�Y�"O��ۂ�@�8@�f�:��
�"OE��ܜJ�92�d�����3"O6�s��۳E��A�rd�`��C"Ou�W@W�<����Q�u�B��"O~T�u/N�;��c��$Q�b�Q"On�P���S��ݳ��3�w"O�U2�
�(a�HH���#6&
�8F"O��c�⃇q��� v��V	�`�7"OT	Wj�+<����I�^&�-U"O��s��1wF�� 7�O$#��Z"O��1&��vR�$R��A(��Z�"O�z�C enTВ�B�
Bڍ��"O�ٲ�)*V~�1��-� �T"O�q�M��h%HM�uJ��cB�#"O�ᅎE�S��|�`	P'�����"Oֽ��Ȍa�BM�!
�%w�p8�"O�����"Qz�M3�oK�tTV��"O���O)Ey�Ġ�izhP�"O8���K2G��|��)����"O�Xf�X�UT�M��X�@Sl]""O.�`�
1���kHJ0"O�p�+�,1G�p��kV`��(�"OP%0e�'�$��V��"xA6��"O����J�rP��c	�c8 �B�"OV�j��Je)�A�",DrF"O�I���-:x���@��#��`"Od���ψP�(�R�D+��2�"O��wl^$(nL�` �lvi��"Ohq�gGճRZ��
4�� CO\�ӡ"O���s,��l�0� ��]�"5B�
q"O�I#b�V�H`�iiP�K,��V"Oh��e�v���V,��p�1"O�	+�mM�H�ƈ�1����H�"OX!���Ӫ�V��l��I&�B䉕R�X��1fܓ~A e���mu�B�	(@�pqb�n����Cߨ&�R�����r	ճ:�FIQ�&УK� ܇ȓB�8ER���vx�)�k Z�l��ȓ~�hhq�,NAݞ͡q��X�&���^��t&�q&�5y�Jڗ|E���ȓ����I�rZl�@T��U��i4�qD�_�h
`FG{�$���<H�Xa�NKD��cR�b��~��б�>nn��*�Oׅ{N���ȓ`���1t���3�=�*ټ]. Շȓq?�8q��"���#��1K���|����J�'=w�u+� B���ȓ'���b��Ask��Q���k@� ��S�? ��{����o	I8'C�NI�#�"O�,z@$Ÿd�����Ъ ��m<D��;��A^�bƬ4&R��%D�d��2�vtRe��=&�֨?D��Qď�?
F�ٳ�]��"Yy�c?D�D��'Y���@N��\ZIB# D�x��$�9R��4zp��|XU��=D����/Q�>�����F�w�\�� B9D��aa(ѾT(�hD>w�B(S�B<D��C�
��;�r���+�.T[VZ1F%D�ؑ��6�B\�r��A2`!�b#D�xc5�+,� r��^:@�y��"'D��P
�	?Ąz'B:4K�� �)?D�����n��0I���0�r�;G�=D��!���PJ/\�|�|��V
;D�P����-� ��M��K�!:��:D����k	?}�q�U��jJn��f$D��3�	�;a�B-�BK��8�!��%D�DX"�?u��1(3#��T��P'D�`��m3D�N]Ⓣ�	�И���%D�: `�p�t�E���g���@�"D�pH�h�%�Xtq�nL�p��H<D�h�3.	<bj��Q�
�>rRਸ਼5D�tqv�I�bl�蓞,���[��4D��4f [�*�Іֹ	,����& D�0D	�`�����;�h�3C<D�4�qms�����Č�d�!�>D�ȋC�X�ä�� i�K1�ip�H/D����КqZ�ث��:g��q�p�(D���W$T\�)6J�-K&�U���1D��A�D �X
|���\�5킉!�/D�h��Q#@*���[�4�~u;/D� ��ƍO�N}@�IV3�@uɖ�8D�|1��VFr!*�!Ԏ�*I��6D��KTAO� +��Su��>~���i��6D�|�DdO�4`<�b�O�j����h6D� �Z	 �9BO?-/�)ɴ�)D���Sg:Kx}3Ǉϰh�BIJ��:D��4���H�mq�Ͷ�� {�@:D�LJE�
`�X��HK�A�ްX�H8D���e�
��0�+	�.��[b�5D� �g�.|�������?H�ڷ�.D�H��@�����S^7���.D���!�80p���̈́�fΈ��,D��`cg��'v�\Q�e��7*��C� D��1�#z��Fλ>K8� �C>D��!t��4l�b0)Y*+2���:D��C%£j�0qaa�0 ���Y�6D����,X�(�$Aj���y�#�6D�<���߂�&���M[�Tᐦ4D���&�"n?
����ِ<�(���1D�LC� u��}*�#�95����-D�pb�D�?jy��B�%�1:�-'D� �*2*d�������ސ��3D�4�Bl���e�ߥS�Ha�-D�����D9S8��:k��PK����F?D�P1a _��0�{�����j7D���&\����×�<�����O6D��3�� Z���ǡ�'�H�vK6D�ಡʑ[p�$qT�E*�.)3$M7D��Z���l��k�U�e`�G7D����i���(Q�(���h�*6D�l�N9��d��P)}�x��D�5D�4����2p��Y�s&L�%cD�g�1D�� P��Dg[)ɜH��%{�i�"O�q����g�~���)C�}x���"O�](g�ٶZ
����i2HP�k�"OZPcDɓ�8@���-��b�"Oi �i=Q���R�3O��F"Oj|G�'9N�j�'�l���S�"Oڹ+��|�4��#^��p8$"Od�;��7�ԓ���c�R���"O��#Z�A��F�<5� "O����F *$���Z�M���#�"O�+���N9iԆ.L�����"O�š�%Ңe8�E�GF��uh��#"O2�" G�s�҂k�$s�*xX%"O��c�$/K�	3$
�?@�uQ�"O�$8��9��5�����Y�&"O��B����%�):��T"O\+�K�!�jIi��սn���"O.�$aػ��l�9}Y$x�"O��IfrX(r%íZ3$���"O-��J/�p���ņ�.@	R�"Obtz���z��(᧥D�?H���"OFl��C�R'�H0��	rl���"O:d@�i #5�� i�� Xؘ�e"O~qa���'-�\�c�ۛ	�H�#"O���eFZ�#rN�s��l����"O:�k��ƐV�j���_��h�7"OЌ��kU�U���.Ҷ$��l��"OHA��cM*2���J�� 9��Y�q"O�p�Dd�)��h 1=�6tҦ"O�֦5`��`���{�T)�"O��[a͵B���sD��<��b"OXr#�.yJ ��LfhJ���"O��㧌E|\���E<<�""O@,[��3�|���)�nT��"O(��%��2����S�BTk�"O"Z�E��a�b9CI�\;БP�"O!q�D�'���1+%N ��"O��zrH�\�h���԰i���E"Oh,���TU�d�Ч�3d�.�Cv"O1�׊�m1��[���bq��0U"O,ȉ���p�(`)r�H&Ia�X�v"O,eS�j�`9���Bf�7QL2(��"O�e��)�Yqh�Q��;,@�m
�"O�ܛ�� <n�P0{�H[�MMn��F"OE��W�pj �:���a=�dK$"O,��ԉ�7(�L��%C�h���)�"On\z0�A6�̹yB�X�ndVl�"O��p�@�1S���%L��jE~���"ORLHq��	9�6��!��v���"O���~��8H��J�~d�+B"O�@��H�'��UBJ��=�g"O ���+���f螀X�nu{�"O��sgdD,x�:��Aȃ�.��@"O ��l*vqk'K28s��U"O,�kgf������d��W~�)W"O���F��i��Yx'׈q��4Ae"O�}s��
]�d��.6 ����B"O\9!s��(����E{����"O*ٵ�=.D���10T���S"O �𱉙�'����'Ga(��"O�\�gGl^X(�k�0H����"O�fg�>{h�ShːfB�U�"OD�%�N�=�1R�߈0%8���"Oh(�����T�8$��l�."�T+D"O� �h'�
�]#�匪O*
��"O�|�ƀ3rZ�����k���"O����U��|�����R���Q"O���M�3<��;��Y$DZ�b"O��C�f�,l@a��	 Bt�"O�a@gM
]�1�㇘�3"v���"Ox��b��+�fa�S�)�E��"OJ�U�Y��ȁ�쎨/�%�q"O��bw%\A1P��6l�iո�)�"O��j$b|N���

E0^$z�"O�@�BȤ4��	��&�+V0�"O�t2��F�c:�ED�.h3f"O��UǏ�Zl8��dV.>-2qP"Oʬ�3E�/]M�ȣ!W�&0a�E"O$�hV ��hCAʍV�Ru��"OP��7瀎hl�ԯ�5@�8 
�"O�����3 ���[��(^��y!�"O�����07>U�P�#� �9A"OD|�Ā
1Ymx8�fH-����"OV��B�&)vF�ӓ�ħ~t����"O�������VL� ��l����W"O�����_
+� Z�%��"�x�"Ol�;��DL�Re�E�����"ORL:`�8h_VJ�C�)
Ҵ��"Ofm�m�0m>01�L�8.Xl��"O>�p5
_�}�8��c�ʢ- �h"O(�����\�h�R�� ̄P�"O,���E�Ċ�������2"O��2@�הa��|㕌S.~
"}�"O�0�cM�L���s�#L��= �"OR=c�F���$�qc.��0.Ɵ}�!��6�ꑋ`lZ�KD0Q�nR�k�!�$U�mjx�ٰ�Ќ���5k $!��9�Bщ���٢�g��#c�!�B�a���i��,Y7,�"Ї֌h�!�������0�.+:���ɞM!�DG�%.l��@_	[0<8�q��1!!��",<�d'^�o!x�C�ԭx�!򤟘㔑"���lm� ����4c�!�D�>s�����9h�d�'���_�!�ĝ;5m2)�ug�:��Hq�O6K!�Ɛ[6��HUd�)�؝��f�D!��Z�
�� §�ˀnU�=G���!�ܺTf��-4K�Y���@f!��G�J2R	�LE�sr���_6?;!��g�4�ī֙赁�oK�w�!�D�Z �@�l�f��cn��w)!�Č�$C�"�J��}� m��s!�dQ0J%�Q��#n{��[v��8< !�dڰ �|�S�/��Vp�88d,��D�!��Z���a �vi���W�!��ɢv� �����-��H��!���3�vu`��AP�Z��+QO!�D;<rf�D�ȱ6P�}�)�pH!�D��oMrd�"�]�-0���H�h!�$T�>)R`c��3;=vqyWn_b�!�$ڤas5���G�Ы�+�<�!�$S${�@\� ć�x��x�j� �!�$ȯ]�ٔ�	$�^���kWJ�!���6�* KֆϩUs�=ɣH�=�!�䙑}��+7C��rZ Ԙѧ`�!�D�� `b0�J=I���CM�+U�!�D�P9P� �3@��}[�.�*�!�-1Ѭ!��`��q���W'O.!�� \��Bc�0���*őJ��Aa"O�`k)�/.�֡�v)ڈj����'"O�Hٗ��"8V�=�@NK�����"O �(�-�;x�>��!c%cZ̷4"On��Q��@��A2 ��	;?��c"O�Õ�	{MM���ZU���y�]��p�t'T�x�� ��`��y��	KB:yY�O�c4��!U���y(@�8�*��PiT���!R�y�N� -��Hz�h٘R�����Ǆ�y��=ZClH�ΐ'31���  ��y"f�?6����2(0#u�I�b��y�v���b���,0t�}�B�I�_/(h�X�F��5z6*����C�I?N�9�� �'N۠��%��Y��C�/DТՒ���:qr|`��
��C��Mw��Q��x3����̅�6��C�	>-[�ˠ@?gF��i��,�B�	
 �<uۡ�ֱ��x�2��+1��C�	�ZL��q��r�` 	B	ȷL\�C��	�yCVn:ߘ-��j��hC�		,�.�s�	,0�]j�\�#mB� 9R�p�KO;G���X#��"��C�4���gYy� ��oS1��C�-r��5�@Y�i��ȣc#��C�	�Aն`�a^#*�	�V�<�C�I)hH8Q���_(ı9�`�-#�XB�	���G��ALl���
rB�I�v�"Ĥ?f�Q!�!r �C�Ic� {��^�g`d��mЪEbC䉥,Af1c��!Bg��H'dG2&C�	l��Jg������e��.
6C�	�	h�P���X��r,�Ug
�)(RB�1�8����67����#$ɆC䉹;��M�� �E�`��u��=`EB�#��t`�>mL��ՊA�(B�ɭ!�l�u`�%9K*��ֆ���C�	,z����q��/��dd�G�C䉍��<!�WYm.-i&!@�g�>B䉏8����W�ռb^"�A�-^=�B��JD 4r  �5m���%9Y�C�ɫS��	��U�H1�l�!b�;�C�td�hv���}��h�$\�8h�C�ɦL,`�R���9@����X�g.|C䉔XFލ��˞�DS���`RC�!R�Bhs�'�!3@��ś%�PC䉽q��Ṗ���0�H� �7W[C�I��б+�GB�}�X�C� ۱��B�I�6`��ED�˖ȕ��B�ɴ0zA�1�55K�S9p�B�I/e&ȸ�(G��	W���dB䉷_����g�G�p`�t�)<��C�ɠ}����GϐA�x�s�֋L�6B�-vf%�bX�ᳵ	V�</<B�I��P{�`8�ȵD��2@2 B�I�}ȌIi�HA�p�
 hE:q��C�	*.��A\�xY�Y0�.�bC䉎b 
fN@Iǔ͈1��=08C�ɱd���	ӏ(ܢe�d&��$�jC䉊�ɀ�E�@��Ȇ�U��C䉙�6�r���Ҥjt
��`��C��x�|9��A*R|��&-	�B�bC�I5YB0��
+�`���%D�AtnC�� %DHKV�N�� ��`,=0<C�)� �����>g^%ð�~Q�"O�M+��Q��I�E�r���"O^�����:�]�|�uY�"O��Ҁ��>"Q�ӋL(gn5U"Ov�c$ߍ^N��'*�0R;V4b"Od�1dO�hY�[$�A2@%�PQ"O��q7(]g"�=Cd�Z�Ԅ��"O��@�kZ��V٣FhY���b�'��AAI{kX�1�K�NX�	�'��9(�G��z�IH��A�4�;�'0V��dO�(b4HXvj 4��E�'���R�a�S�u٢��'bj��'�4�$���#lk��+E���'I�ٚ1�>@�n�H�/���N���'C�y#d��p� L钭];h�hep�'ߠq��]�A�t�El�q��r�'ap��̪���H��Z�v��41�'v�q��gOMD`K���~�V���'�z�ag ���
7� �gt&}��'������$6J�X�"��W�rd2�'D �����v`D�U�f\��''��{7�����1��QW��
�'�����A�|��� [5�A�	�'/�Eр�}�0$�Ё�
1;��	�'�xaQ�������/Ū2��a��'Ӓ|����:����`����*��
�'E:��G��DU��E�*�F�b�'�p���$xJQ��91�6� �'\���N(�	$fG0�9{�'�X���Ɣt�9�Pk�z���'fa�F�*h$�&�]��X
�'A���@�q�yq��P� (�	�'�X�r�� mzdhq�Ɏ�L�*!�'���ȣ�ҕ�<�� �V4<ڄS�'�6��$f{9ZD��!_2�q�'��u2F��c��m����"FF��'�8���?=ax���Ђ?�1b�'X8��� !rL�Wc�6B2��'+�X8������6��a��'2���-lh�Q��)�0:�'��,#`%�<i�\"�&�']���
�'(� 5�֤laA��%l����'�%��=�V�ii�-�I;D��`�Ú9:�gbBx��還N;D���s��4vlL����Ֆ(6��aS�6T��ȲmöA����wI��@	Kb"O�踑ez,��A�G��Hnr���"O�1YT��CBX���itԊ$"O�����_�}t��R�I�1��{�"O�m��G0iF:3T͌�o�|"�"O� 󧁃�s���@�����@"O�a�Bd�\�<�Q����j��U"O��*��$>� I���V�̄�"O� ���~R�D��DXb�jF"O���Ε)����FNG�O���̓/�*����y��(S�X�{�����!]��8�@�AƒP��5�h�ȓ�@(ħЮPL�@��'��1���y�|� ���)֩r ��&'r��ȓ<"�܃��1H�� "�n&<��	Ŧ��&ύcH@�HF -�Q�ȓ@Fn������. K�B8rL��?Q�<�U��^���b f	9�N���%��K�о:��!�ݍ����S�? ���k��
�t����˰["�X�G"O��TL�O�MhN�,	B@�5"O�i��G�6|��E2Pd}C5"O-*D�Q6S��ig�;]~1(E"O��RbE&ʺ͉v���Pތ��"OЙP0�3c`�1C�D�&6��`"O�)��1[�nu!T�u���"O��ڑ��ߴTR��T.Zq�9�"O�,� e�b�>;�<\er���"O��f���b��؂��mj`q�"O��)�D��^���)2a��k^LA"O���@ŭ@|(�ԏ�3^�͘Q"O�D��㇜*X�c$��dBV ("O�]�1"gɞ�I�ě8�c�"OF��b�2]8i@�d3Pc���G"O�i0c)�d�ҥb*9X�f"O�Y��.hm����8d�c"O�p��ʊ��\թ$�K%,q��"O�M�H��Iu,H�ՈL�
�y��"OJ}��ЪX�����
�% ��"O:��v���Y=�	a��Cx�"Of�J�(�9^p @��k<și�"O��+$,�!0$��N	>7�u:�"Or�R@�[3I�I�/C�vJ��v"O���!\�4Xe���:D�%"O|�+c��+TD��ac��Kc���r"Ofh8VB�}w i!�F".7jŀ�"O��i��������^�1�"O�e��A̗e+~�A#JĪe��Ų�"O*L����)�D����$v)t�0�"O�J��Z�d��q�I�QNlq&"Oу�G�j����F]�fFL#w"Oܸ1� �j0d��� -&��"O�$IѧI	3�Ѝ[��O�.$�"O���$�0�� ��ዮ�l�З"OR�Eˈ~m�tx���3H�����"O�����(	�.� �͎r�Z8`"O��K6n1s����mQ1���"O�A#��v�h��ƙ�I�<�I�"OUx�בd�;����mͦ\��"O�i���(z�U*Wl�H���7"O�h���Ȧ� ��ʮ6�d""Ob]��/�E�N�g���^�P!D"O�I�TˍUR=�C �	DL(QP"O��bnX�f�5�TH�#�(�u"O~�i�cD7[��Kf� 9TŒ��"O��X"$&V��|Z�G�>���J"OX�����!g�,d�C�v�	�"O�9$�B/|w�!	��Y3d4�ܨ!"OL����E'm+��Պ�5%,��"OnŚ�[/F �q%�C#Ό�"O�Ш1�؀u��D��FׂR��U"O&�c��2{�H�a�t���Q"Opx�R�M`�<��r/�
[����V"O<XsG$I�5��i����Q�6��y��>k�)�铁hനZs�ɞ�y� 2M�tP@I�5*(��Rg'�y�r�V� �B����+#S��yr��;�X�7��q�Hc&��y�#H�V[,!��K�����PBC��y��/PW�p�i��~y�d�A�>�y��V���@�V
s�Qh�O�y��!/rP�2G�Y��� �僼�y��Pq��	� W�4�2$�y
� ݋���0dbn4�.j�Z �"O���ސv<��'Nۄg�p�0�"O�H2�8TA^���O3iO�;�"O��k���5 ���v��Ӏ �h�<ç�^�;U,]@a������}�<ё&�:r-P��K+����DQv�<����,3�*��ҭR%��=`�G�p�<a`��edy�W�G�8
ε)Sm�<��aZNi��4d[6c�@Tdk�<�4IÁp�:�
",��'Ʀ�3D/_�<�r	C�;\+��R4�A�%�!���T�v�`D�@ONNh�Qi�!��*@��$
׮�:h5����+�!���]u��`�2]X���H��V�!�Ąs��$�r��"�N�  �(w!�d��<u2l;4���O0VM!���\7*�0ԋ2:����.Ǘ)2!���5zԙ ��P� �ڣo6!�DLr�X���M�1y� �	����3!��"L�0� W�P��R��(,4
!�$@&ט��&�>l�p��[?0�!�*tH�)�aM�.^.�F�E94�!�d\�&�
� �CG8C�"���!�$T��HjBB]
e(b	��aM-�!�$�;Zr��&ݦ\��#����1h!����W�Z�`2��S��b�$�<-!�7'�
|� 	�+�8p`eC�By!�d�!���%G1;��}JW��D}!�$O�"��D���v�ص�ǳv?!��5�i��%ޘ2��h�vh�3!�$ħn�Đ ��6�(�6�@-!��=����h^����*S-!�$A<�(�H���:"�&5�өS?%!���8�aԃ^-z������ �!�:E��<�dM#6��5c�Ϭ�!����%cՠ�o�✈��8Sp!��!���`�	��b�ˆ�A��!�A�FQt-	�Y ��� B"�(~!�Z	=�����%�<E��x`���m!�$��S��rbƝ~�-Rc���$!��ߜhr��c��T=��ʠ&�"�!�ğ)�B���ŕ)#��GG�!�D^=.;N9���
� �¬z�h�t!�N4 Ц�ڠȘ�;����gCo!�dįME��y����D�0�Z�GH�=W!�d�)T0���B3����E���JV!�$<��)S���atܘ�ֆ��74!�d�v&���t`G�#��(x��+!�D�6!C�mK��#KȺY*�dΠQo!�A�;�b�q�.(ض��tA!�$�N�F|�Q��j��[5j�	T�!�d�;}��!s�42�@]) �&�!�$��~�%a4�F�^���c��.V�!�d�%v_��Ѵ�V�&�lʆ�X�On!�d�$��P�F �6Ց�`S�:n!�Ċ�
y���s�	�n�4�(f!�Ă�wh2[qB�<D�p��W#`�!���?N��|����:M~��0��˯Z>!�É"16��$	��G��0yF���H�!�d"*�>,s1����YSO˅�!�d�=N��S�ɯiw�	p���w�!�d\�a���Y�	��5a<H#��ó:k!�D&SϦ��Ĩ�67F �*�GI�|d!�]�x������W!����h��!�� \�8$D�,M|���&��B��L�""O<Ly���Gy܀z�ߤI����"O<�1��Z&k�(�!Li��`3�"On	���J7th�h� N.R��"@"O��)яXڜ�y�ƌ^���1"O�A�R�ܤ�Y��LC�n�ȧ"O��z#�Y�B�Hk5nA�n��Sc"OL-+��5W�d}�7�y�l5�"O衚�Nժ茭! �߄&�fY�D"O�0� ���u�fЛ��^��&m�"O���W��8	xE3�@(��1p"ONA��%��-�J鶁Ӱ!��%;r"O��B�kӼ ��"[����i�"O�e#��$E���2����J	��"Or�kR��g
V��MK�Ԣͨ�"O�8x�EK).�HL�+́���YG"O��[a�Ùp��	K��7�PH�"OvI{�$ؽ\c�|+���`x@��g"O@a�ϻV� �"@V#I�<�"OiF��6]T��`L�A1�բq"O��0���T�N��v/1+���D"O��x�o���bIP0P$�t��"O\��%ꇡ�����H�T��ܺ"O40����D)�q�Ea�+���;E"O�1*���)�v��5AS�����"Ol$����&0������Cn��p"ON���, �fBB8��Iy��+�"Ox�#�0�t���:<CH�{3"O�t���½��){�_�T�t"O�`����#��$R֌&c�ȡ�u"O���F���F
8�M�'�.4q�"O~qڔ�8,�Hu��`+�@(�"O��� C�UK�W>9���"O$Ț ��9U����E�78�H��"O@�Bd��fd0�J��L��U�a"Oʡk�
�"�8y��I՘u��"OJ��%Z&A�T�P���q�
-{�"O�`��K�c����F�$�"O �ʷ�ت7�<qSHTݨ@�B"OPp��Y�N>
���h��(��"O@ �(�Z��a��-h��|�"O6e� +K(H��E�����"O�,qӥ,jyj=���'
�6h
u"OV`Ö`TA��d1�I'(���Q"O T3d�%�쌋��n�M��"Ov\Iяμ���#!��LÎ8*�"Oy�7e�P��0�1 �c��x�"O�1h�~ղ�XgN�#�R�(�"O���͛�p�ڭ	%��4f�����"O��`	�b#��f샛j�,���"O��9���	]⥊��	$v�fp��"OZ �Lߜ	Ȅ�
��~o*���"O�� �J)��!�D�>o����"ODj2 [�o;�P�"Ob���%�����rhJ�C�ڬ�5"OU��f�2;��Л�h��;b"O,�����{ ���U�@jq�	�"O4}���$|�(MK��Ӓnd�$aA"O�� T���+L�#��B�"�!�d�).4�X�ĪK5���pg�L��!�$CEk������*4��iA'��_!��B�[<�95N��WP�:�d��!�d�4!̑)R���,�����Z�!�dڏn�r)9C���S8~1��"��!�� V�$��,�\���R�l4ٻ5"O��� ��f�bE�`�@�@�h��"O�IY�dB�V�L1ą�2"U��9�"O��7L���m3�� na@a��"O^5:���K��y�2I�!����"Ov9QNZ�*�9�jA�B옒l]!��8��������7��W�!��n~�:�S[�(,r���b�!�ϹU @�E�� �$��� [�l�!򤇠�� �d�V�o����`ǅv�!�S��G���}�&�;��پ�!�d�7$�*����&\�,�0N
�9u!�$� cF��5��h+YW�'
�!�Fa��A��;V�m��	"�!���d-$mK�׭x��%���׏
-!�$}eA�� 
�N#��r���ȓ�h�
ʄ=����ě@(n��ȓV_R�{%	C� ��� j����D��Q�^)�q��B7��k��(����	R���ׯ,Il�S�o5�d�ȓC�|A�c�� 9 �$��T�VW�-��H���V�XԺ�R%��)b����ȓp���ɞaBlX'Ͽ=S8х��@��aY��*x���H6�̅ȓ�F����d�*�&T/)rȈ��+f��钆�6�dl����H�L�ȓK\��3�U��r����G-�H���w��X+R�O�G��kM�T)2I��ge�ų��_�O@q`&cn�м�ʓs�<�&�G���J�m+�@C�	&w�6�iP��6{�1���ݞ��C�	���6%�a��AC�B��C�I#3��%3���/T�!�#ؼX�dB䉂9ti�ģ6�5�r+J�PsC�)v��("!7G�ZM���72B�	<��H�Ϙ8�P�b�;MB�	�cHVd��cRw�z,���Í�&C�	^B��S��T �8t1!��!s�C�2YoU�v�q����fI�+��B�	#|�r��7��5�h2�H5ϮB�*>�1��R�Q��`�f��q��B�	(��y$R6�$�E�D$$�hB䉢{�j6�F$��yd��bHB䉹v�^y�&���i��Զm�B�?Jx։��QasVLy��z��C�	\��T˱.E��>x�瞴�C�ɊF:0iL�|{8�4�]��B��2�V�if��I�$fJƉ��' D��A��ا<�Eh2HJ�B�����=D�<Q3�,p���DK�d�0)V�:D��bU�_�=j٘GK (�q9D��[sf�%t����L�f"�X���7D��	� ��5�dya���/�n(M5D�ǆ�6u����> �D0�J5D��x���,�H�Ia 6�ڜQA'D��D-�h!tA2�-��W�ru3�-0D�83�aI�kEa��Č,��p*U+D� �@՟�&���!�^���I(D�$@�m�0*:l�bǈqt~ջUd)D��P%D�ts��EBh���%D�aՌ�*4��D��<-"�H!D����N�x��T"��c~ ���I+D�@��ȇ	�8��$�9��#��*D��z�ǆ30�\�3s�Nw��]�7 &D�� (�i��6X�D�@�����@"Op���<���S�]h�l�""Oh H�F�&M3�M�eJM(
�"O�Ԑ�N�2R���JI.=���@"OZ181d�&:�l���T��x�"O��"R$ԛSW���R�Y�uFijf"O���%��z㔩X�m
 �~���"O|��q�ۯ.�bt��3z�5�B"O� �1�G醍�FJɽ0{�"O�ejc&)oޕ��)������"O>� ���/�F����D<�0"O��	F)W275°�է�,Rr�-��"O�1��I(R��a�s Zp"��r"OV{�ƠVQ�q����gH
̓�"O`���4��)�t���'�(:�"O�T8Ŭؚ�zI�#AV�}��
�"O`X�n��u��)@G�DiQ�"O.m��m+c�d�袥Ώ;�T�x�"O t�1#�Hr�¥�ByBm��"O� ���H�V��ۤ��)D$�w"O�iYbC��L$��o߆�̨s@"O��H䍔�q��l$ц@�4"OQ��ӟI��0�.�"O$̣V��U�U2��m�P�Q"O���2��%K:J(3vK
�O�n�"ON��bٰOaVES�jC�z<���"O�!��g�-R r�\:\�Ρ�&"Oh)i���Y�JD�gȅ-w��Hy'"Or���X�d�ЩI�Ɠ�mV�A"O��3ӫR�O����F�r	&���"O\u��ݺ/��X����;��! �"OB=�'L�	T�\,�GCݮL�YC"O�� ��98� �|.�ҡ"O�,Rg�.c�ä�͡Ch|8Ȑ"O���Lۘ.l2$�r��d\|� "Oht���">:�wO�lM���"OF!2����$܂!�~6��V"O,0��ЅM�U"��_�n%�k�"O���v����l�%��0bdX@"OFu���M>G�ޤ��gů�P��"O�t��J�Mb�I��W-};"�s�"O�y�q)��x�x���& -����"O�!�iZ�	^�І#ƗW�U�"Otp�W���PK�d �	*`����"O�)cuN��
|��*�� D� "O`�Q����+���M6�|E�t"O֬2���C�5@��ھ4zt��2"O��*'�F0�=��Dfu<P�"O�,ҷ�V<�e����,R����"Oܔ�󥓇?T0�%�X� �I�"O��`SI�nn��C� ΦV@4L�"O"Xa�Γ�����4bсx]�ib"O�3��z�:H�4�J�e��"OX��#.UL+ ��.@@��"O8�"�+Bi�X����,6^�ap"O���l�]~�aX�k��y)�5G"O4Ah�E_����+i��i�"OH���F�m�j��L� k�\���"O��p��
��lZs!�di32"O�`����9c�b���4Ln�e"O�Xi�Uvh
Ǩ'jvŒ4"O4�Jpj���݃A��D\�qh�"OTp�GCM�{�|I�X$so�B�"OP���'�'*tq(�a�<?��}@�"O� Z0�rA�7V�0�*÷WLy�"O:�򋛩Kք���JH�:dv��1"Oz���(>�	�´�^�A�"O���f�0a�!DC�O��HYq"OHH��D+���E�(4�L�[F"O�[b�0,�pY+ԃ"\�L(Y�"O��r I�f"��%��$]���Z0"O.m�s�\�v/̑�DQ�.{�yI�"O��ද�=	���a�ԈRr,
�"O�pSb	�Evb�@���>u
��D"O��w��jPcF�շjjRT	�"O<9��cb .����(?za:�"O
����8P�4 @�x�a�"O�@q��Ѻf<Eb�EM�'
�k1"O8��q(�}�R숗�|؈�"OpQ �!oreÃ䛵`
��"Od\zg�_�`���cD�L�R�"O���B�*B%�hH���H"O�srC�.�q�`�#�΍R"O���r�t��b����B�M�m)!�Z7/����(B�҉A�,��
��7O�a�sɏ	�Ƚ�Q��%���%"Od�!��Er,]3%JE�c6�-�v"O�������J ��C;j��"O^�s�^�H�s! �pJ���#"O*ɷ���	|J�9��W�y7�M��"O6%���L�j�����{'�\���'��OD���,k�: K�*T,�TJ� �B�!�Ă%>6T\C��u��1
ϥ@�!�D�6S��� g�6w�E� �J�!�d��d$
�r���1b��!I�G&!�䒙
��!�/ɶ��:J!򤙷#��mI򦆎S�܋r�!�!�d���hѠ��kG���G:w�!�$霼�ddR:?x�H$�!򄃦_� �3'Q]K�`�s�ǕE!�$�<�����[�:���J3���~�!�
6q��S$��r��(6g�0"v!�$sv��B�mJ�Jy�Ī@�Q�	i��(��y�0��)�V�T�?e�@�k�"O���2BM�26v�PEV3�^l	�"O���2F� t��x�c�7wI�q"O�a���S��0zf�_�)B"O�yQ�Hw�����J;#�H "O�t��?��%��� "Od�c�V�hp��I�Z>�\�P��4�8ړr�pt*�M��~l�p��լ��ͅ�g6�� ��G�E'��4-�h4(��Lv(���P8r�P%`�N@�{����Y���B���#m��J�.�Q�x���)n5s�
�H�.փUh�,�ȓ4S�mdآ}Ǝ90�\�i^n��ȓu�)�B\�!wƱZ4鑯�	$�`[�>�Q�+� �dE�BI��p��0���H��,��'�
@�R
�0r
"��5l�*=`�9�۴�Px��b"��+�!�(��&� ��=A�O�p��'�́Zq)
֊q 1�iΨ�R�'(ar�[�0y8��U|��ZVf��p>�I<��jӇK>�pCr
��g���b��G�<i�� =�X�H>eڤt��@�<�D�]2T�x���ռV��� �r�<���[�Xq2���T: �ɣ#t�<	�'�fF�iEW�m�b�Y�Fm�<���gа �7`�%qgg�A�<� L�s����;� �і%[�.�L\S"O���̀�9
���0�ƞ���ȓl��@а��;{�b$:�jԍq���ȓaB�%���`Uv@�#IU	w	���+W،zb��`#��)�`��h"����H��%[�^ [aL�1䙪,̤x�ȓs��8c��V͎����*,�&��ȓg� �rBEN4�ЙA �$]]E��i�r�S�4o$,�bd�6.z%����alÃ��R�4F{P�ȓ@��T�2�	_2q8f�/X��H��N[@u��7�p�s�$�0��T�ȓE��0��FHo����+}C 	��| $����R.xX\���͖�w���Fe�E�o�6��Q�,rڦ��ȓ�|@�0�Xh=�5ԧ?=�Ʌ�$S���ĊP�C��5�AՆ�{�py+���-�쩐g�"d�p�ȓ:�r�)ţـ]�l�R6�U��B��ȓG�y�"Ȱ&�ppbu��%s���ȓ1��B����8M�#�ʉbq��ȓ����m�"Kq�l�`�P�H%+9D��1� �j����M�k\�(n*D�t�E�$���@�7rЉ�h�+M!�O5��I�"IV�\��QE�"&�!��+�L@��l�_ݜ�j��V
qġ�� �6�q�ѧM��<��F-9�y.]67N�U��F[*���@�aN��yҏI>mR���!ʈ�C�"i��yB���98-ȧA�,*�i�q���y2ڠ����%)��e�d����y�D������3,�)4,�5�y2
�p�����]�l�b���y/��#(�Ѫ���Y&\�؀�yb&G68�r���@Y%<ئ8�����y�΍7��2�#�#)�^������y�@-%�&��@��Z�X�3�C�y'�$��3�
 0��ѫ#ច�y�%C�a��C�7�	ateD��y��I0-�t�"�FS�~���
��y��4�4�� �1%:��0�y�Z��ywg��c48���y�%" �����"�py ��:�y҄R��v�3G�8�,�dD��yb��6~hC�OA�(���3�0�y�'	Ĭ��W*����W�fP�`��f|ҡ�$��@�Xq00 H+YV��!61�d�	�)?4�c��ag:%�ȓJt|t�0Cd���艄ȓ|��@C�2�Ec��2�l�ȓ
�4<�kǼ2��᪡)k_V��ȓq��L�r�T�z	Z���@Z�H���ȓ �� ��MJ�R-,\nm��7�p�����Y��dj���KYX���8 �5��rQ�� �m��\���iod��&ř@�Jݚ�V�Pyf�� ��G�ڻC�(z�B��A���}��t��"ؐN^ �6�ч4m�ȓ�̰��X�Y:0�ae	a�p��w���h �B�*Ϛ��䆌���Ї�&�����9(���υ�)>l9�ȓ*ժ��JZ�zE�M�g�L&d3Fq�ȓhj���cb
�j�@�x���$b-"ȇ�z�TZ�nX�l��0���(`�&"O� �Ha��:
�B�[`gܱZy���"O�Y�R떻h���ѥ��_�0` �"O�����8�~LцĔ�z�B]SE"O�P��9e<�Z�cS3���p"Ohi'�׍8b�L+�#�(<'8�{6"O=b�ׂo�0�0� e��d��"O8���d�@�F�yr���F�кr"Oҕ�Di���a�W&P=��¡�&T�| ���l�*a���'�d��)<D�HJ���:2��Ӭ��M�*�`�7D�H��D͹b&?/����!�0� q�#+�;}2���@�j�!�D�:&�y3�I�]G�ts��	'r!���:�1�L*D��F�V!�d֨��*��F�4��hБ���!�$B�c*!��B^3 ��#���!�$�3m6x
a��/̪�)�ló4�!�$Y?�\�E	�?�"��NG�+|��ė�c��� 0&�U�\I�����y��i�R���)�>����B��yRn�^޲Ta�%P]S�ȡe��yb!X�iܖ��S��XRX83����y�F��� X!�!R��);�(��y�i��f����ц�,4߶�3 !�>�y�!!��{Qc\�/�r���� �yb�@8N+��h�FJ9'c����^�y�������k��$�v-�;�y�!��Ę�~���k���y�)@%�8�Jb��x���jI��yrJ͙<��3eD�o�@a�ѩ)�yrLTe�<�X�h�cz�X�b���y�g��J�b����(Pyy����y���m[3C	�b�$"��yr.�9t��5#R�R4ϘP$O\�yҡ�4~���V��.|0��I� � �y"f��+KT��5�
6o��E 4����y��Nь�9�J�a�Z*sH,�yB%�N8�"mŔSN�aR6�y�6&봱`�J�Z�M��N���y�فI�ν�&���Nİ=���՝�y�\8��$A�J(pJ�"��y��k�����6��;% ��y��F�B!��^6l�q��-�0?�ײ;���d�>��( U ��{>���o�b�<� �J� ']�Tk\%'��pD��J�<9�_0Ve
}{u�S�Ml�ix1+\O�<Yvo�G�t����]�KoZ��
�K�<e%ș P�3DM�5S���R�JJ�<A�B�a��!�F���UK�A�<�� �^���plG# �lHP��C�<�P�мM�"!"� i�8�(�z�<yw�[�V�)��I4<�I*F�v�<���C�{N�%�婛=<����Bw�<���̜C�2�QJ�DR&�1C�Pn�<���1�Fp�V�<�ȹ��_`�<����`1��� K&	$Y��I�<�e�
H�(�CկN�R�ݠчX�<Y�̄�\��y�'ɢ0���H�T]�<�NМ(��ā����>�xRhY�<c/���(��m֬[�R�����W�<	�B�Mk��[1��/lO�)��O�<9w�'g!])�O)q�* ���M�<�6&5h.�!�ᯜ$$'hD�a�<��"U��I��,ҊX����cCp�<� v���=#"�)ա�y� ��"Oҵ`t�Af.�\���-�F�"O��`�aM�X�0�$M/��jF"O�d*R@�"z
e�nV)p<4i@"O���f�J(f�8�����ud�(I�"O<=x���<�Z4;W�L�hm8!��"Ob�p0EK!���C�ט`H64�"Oh�7-F�CR���K4J�M�"O�I���%F�T*AG�x�Yu"O� CǪH�A���C��/+	���@"OT�SCF+v���@�a�>8�6��'��ˀ��T�Д�o�L����Q>%��SG��!��!�ja:e�K"M����?6�O���Ї�5A���D�L�E��c>��Gf1h�� ZVF�*~�����M$D�(
��{lQ�m�r.��{P�_�F��&c�g�~88�b����!��Y�|��N�./84q֨P)��#2+'D��a%�[ 1�VYp�!
�<`x��OVм	�필�������Y���i��D�H4�����\v0TIC��^�azR�������H��T���� �֥���)ɘ)�k�0d��/Z��4�J�<AF�abW��/F����C(��H.E�����Ȣm�J�#dY�tр`�B�:�G	X�o=��6�KP��"�J�S�<�'+M� ��i��q}�h�$ Òx��(�q��e���!��J<4����K� ��ݟ�ʱ��)\@�S��B�I�s�����BT"�^m��`��� �oɭi(H9JP�Ԕ
�I1h�p��Њ��;���n�5 rH:0n�<=,
���ӺDԈ�i@	��u��`tn�-ԭ�P(fC����Ńq�����]z��rd8�O^��lQ81�P�Ȋݨ��>1�"6�Ms�N�U��Zg �-xqqÛ�����cGd�Hά�~\S�l�ZB!�_a=ĝh��Ȗ��"HY�}C��Xv3�@@)�`��e�w�O�!c��q�G4�t9÷	�&PȲA�h`��R
O���d+ـ3�U���7�(�B ϒ/�� 3�ЧdԦ��	C.���,f��;���H+6�@�1�kȩ bo��S�Q��j���G:)X���'���SUKI(0���0��RM &��	���c4�X	G9"��D � 1l�$9p�'9��@�õ��d���s �A�<PCah�^m|�� X�5
و� �6��D���G�q�Y�cю޼�2/َ~ة�0'@�q�ry���+$� AԧrJ�X��^�O��A�%�@w�@wU�"𝓤���aZ�-Y�'�pH�P�A^�M��U+��x���� �����M�����6�O
`��-���
顖)��8 �
ĝ�[F�Y�b̒�j�V�3��+'N�	��D&)�:�6� ;�Z�Dܱ\H�m�Ҍ�<�r���	��5z�H `GC�~�'�nx󇩙�����CH��h��� ǵ{��:�B�"c�(�1���d���w�$!�	
&J�q��apL�x��X* �I	mb���h�u�l��"��n+6-�����:�v@g,�>,dn�� az��S(�4�yb�fq!)��26�H:���8L�4�ڽ',��0�ʥQk�,��	��ȨZSAY�w̸ȴ&2K�ܙ��(2��a��L�Me$�4!����@�N8	hND�$wgf#$d@�sJ�Ro�E�@89�a{B� ��9@���CB�L�t$�P�iC� �7����k��KG���.ڶT	�q��ڿK�:l��XT�A5@5�����O.U���Ӳ+救%�%q�U���d�1C������ϝI���׆�A��1[�ɛO����#�Ͽ*�������@���9F�䃒�j1@����6����S/�c�䤋��U1�쩇hĭ�&�N�=B��#��H�Z��9g������7���׈į��C�Ώ�e��C����E�(!&F2?�J�f��8�*��$N>n�i@��/[|�R�+�e����&`A���"冬q�>�Q�n�����c��U�Ըu.֦5���X�J����_7(�I���ȟ_ޘPۓ	��s�ڑ�
���m^/V����s�O���:�DP&��b�	K�:L��A�j,N�I" _�U����$���
���~B�A$p
�<����OaJ���Ȁ��'�"4�@]+�� B�pNS�P�.0���(���G߯��LC��bIHb��K�
؋�o�JY����a6!<B��$/@=��OJ #�?x�aoU�p,�)���D18 Ġ @�F�8��Y��B��C=t�A�s+��a��26d�jM�7F����@��m�ăfN�7R���r�18�����5I&�	�E�N�`���lP��bޢY��,K �۱20���'h6I(�1n��d
�d��;�@s#��=���X�I7Ԙ	ߓ1#�����d�P4K#*]LpKV.Q�-�h0:q]b�n�Q�e�5`���BL�"7��)F��_Hx[fN�,�n<*QC�>Ѧ��a�T7$M�T%ҡęs�';�(S����J�� T�H�/��B�	3fؐɚ�O]<�ȼ�	�:�c�\���7mҙ�4k�c�b�*��d ?�wb�H�&�=#���Є�4�]x�N�j����ȝO[�H��ŞMZ�L�P�te�\ShՔ7�Bqzw&J��ژ#�Ԃ2�PEq�ش1�O�Z����N_:���A}��@F;t��T��ފ
hR�0��Y-e��	�g��� �Z�속P���Cd.c|H���'}L��A�!�\�T+A`��S'�Դ'\ �V�U�H�,vI@�t�HI�O?�z&K	��XiK���:tf�퐦��~�'��@P��v?!�G4����:N�8�� >R���`a�'��|���E�"LO�T�AÎ�+dzձ5�`���r�]`u�@��i	���!>��y[���0�XC��$�.|+�%ݗ�B�aG(V5�
Az��C5Q]qO?�	&nZ��t��#�dd�5(��
�PC�ɑ?�|p(�!<�r��R�^�\�6�	q<p��'1���DB�4�Pi�H2&�4�A}��!��T�`�@6`:Tz���p�C�.'D��0��N-͕b� "G��[�"���OTPh������(�`'F�#$�5�h�츹1V"O��aA��-&�ƵBf�E�pqr�X��,��?E��4I��a�E#�" [�̂�]�L�ȓ��ɱ��5c�\ɂ� ��8v��ȓ.���n�}�@�2�e<_��)���p�0PH��iD�x9e��L�tY�ȓP�Xh*��,4���tŊ�"p]���&Yҡ̹G"���۫,
��ȓ+�p����GL���Pu\� !���ȓ�l��ʩ*IޤP��:o���Z��$[��S�'O�Ae��JC�Y��h�]�^�)0��^q^L@�ȓmfi�ЯV��}�LT���-��w���ئF?���bh$����ȓ}	�����uRn��s��q�ht��:���W���@7<Xj�ΟEWB��ȓ"Ÿ�Zu㈍Ce��&b�=�`ȅ�k�D�:QD��eɈ`2e�1���	�m�UʵY{��i���w傱��I6v���Fؗr`��A�89���(����3��#
���1&��G���ȓ(�H���Sv<x���'-�<`��$�XzԮ^�*p��p�/m��q��6Wh!s6�J&�,����&Ha:���=�BXPʘ# }��:���4V܆ȓ��"�@QQL@��H'_rL�ȓ]z��"��C�'��%�[�[*��F�6q�`�ٴl$�<�b�ȓKlZ!D��|��y�P������5�F�Ŏ Z$b)�W���L��h�ȓdbȴ��A]��L�U����Ѕȓbt������=�>E�)��a�P��ȓd8�B�ͦDrC T�'�� ���V�c�,וDK����.����ȓi�^������@�Y#�f��u�9D��*1�"^D	��@HJ���7D�ta5�Y>F��U�ʍ!>�%*O �#"��Q��:`��V	�1�B"O��I���6<T]Q�c�z�P�K�"O~8��Z
F��{bC6)�^���"OHE�(P2r���6��T�"O�r2�$Ȫ ���)�V���"O��Z�阌p��Q���?���Rt"O����ŗP��
B�Qw���b"O���4�ըs:4r�aEth��iF"Od98" 3����@�]*1"O������q��@ןgL@(�"O,�JrD�.N65�W�W�q2h�;�"O�9�E.K�}97o&��D"O�ᔅI�W
�0�!�m�DiJ�"O�K� ��O�J}�A�Ҋa֌)�"O�$* �)�r��4J�&2R"O� �m� $ҷ4�^M���M���uJ�"O���JF��*$̎r��H�P"O�	���O�6�Mc��f�>2�"O|p*�F�=o���0aN͋1����"OR	ÔV?|rE�͎Y8ڵ{�"O����ß�P��M{R�J0*�|��&"O��"�͕�y����:j���"O��0'%GF��hg�_�Լ�W"O��S��:l:�Y�1g38D;�"OP���F+�l��JG$|���"O(DI����>�l�1M#YBR"O���@�$���`G��K[���"O$xA̛/IB�I�Eߎ\� ��"O �@�C�8qU�����Al�#"OVYR�Ȉ�-%*U;��/{9��u"O}����҄	k�[,`颠"OX�8�E> T��
�_Z�"O´�d�IڒE镳�0��Ў���y�j��1HM�G�4e�q�1ǘ��ybB��{}Ķ�-� !��q�A%^.�y�'��p���1'�G�
�F�b�e�8�y���VD��'}��� ��I�yrS�Z�d�pC~����3��yR@�?|�������uʵi��y��*�0�CC�eP��)�i��y���pF���b�
w .x'�@��y�	Αiqj\`%bI7tQ❺6h*�y2m��:~"�SA�M�L�̀�#]��y��E���z����f6� �,�yҀ��ZZ(�35��-�h�D��y�*�0�x��+X���6�y��ЭTq ����
}ܙA��y�L4���8"Ej"@��yҡ��'�j��!��F>&�[�J��y� �lN9Q ᖟ5��<k��߃�y�	/��*��O8U��}kC���y�C	m{�u�R��Kb�D��Ɗ��y"�U� l�c�ˁ5~�"Aj5��/�y"1_�S�������.���y��:� H�䇢��a�MF>�yB��T��u���l���X��y��3G+���4�ۧ�q�e!B��yb/�4KXa�K�Bq��h���y�Ú)!L��!惋'A���cJٌ�yr.[���4���ٯ.��)k��yF�Q%!e�;%���;#�	�y�$\�c�J%*婞%��g��yr�W�Y�4��nF[�٨Ō%�yN�������)D8��;E뙆�y�푷8v�AR(��t�V��gO$�yR�L�0�6m�@#�d��Z��/�y��E�T��l��}(���yҢ.e���g�S�8@�T
�y��է[��]i�T8Q�,(��3�y�E��:�\<���?�~p�q���y�܃lk�؇-��	ɱ@ġ�y��P�
e�0LX4*��W��?�y2���#F���H�亰J�h;�y2b�/Q��h)5��(}�̠F��y2��6*rR'��ME���6 ��yR&���pCÔ�6j���y�*fP(tx 
C�G#�s��	�yR�:�Z�M�:����b�^1�y��
��pi���Q0��"���y
� 0Ͱ'e���Uˠ đ3>���"O�p��4�>�����Nf��"O�m2��N�m(�y��E�R�,�8"O�T�CE �P_��l����U�`"O�1��nӇQ4�d��r��h�F"OZ��-��@���2��,5��:g"O����iې�&�S��ߎV��:�"O�����ې��Ū��#u{�H8�"O�@�v.ʲ8E"K�K�*W
-�$"O��gF`�!���qK6@'"O��脂!$`�KCݤ0����e"O�<�֛/��	��۬zta��"O�Ua�OЁ'R�0���ZD̚3"O���41dp�"e��k*ٚ�"OrDG��4����K3���@�"On=2ũ�[�nl�0N6��P+�"Oj���F�����gEF;T�@�u"OP�x4�oU0��d�*H`u�"O�ȸ�͂lD�U�5��he|-*�"O���A��C�8E9���ɐ��"O��DO�:>@(j/D.�<��"ON-�E �7 ��+WnGp�ꐃ!"O� �*��J����> ӚA�"O��c�-B��ض�X�#BA��"O������?Y��2�ZD`<�@"O*�ȷ̜�[GH����(5O�$j�"ON���χ5�|i�BU�%7��'"O��r���@�� ��-{& 3�"O\1�Cd�h��zSD�G���F"O��ʱ'F.823���}�"OС�tl��M�&n�KU�)0"O�h�#��-2��9�知w��i86"O@5�TjM0WJ�0F�~�0PS�"O�8g��"-g��jt�$T;2���y�)J�}3z����A!LP����y�ϓ,Z�t�,Z;(��a�C��yBkP�H�̝do-C ��!����y���_���˅�W�b�q)ɞ�y�b=V�x��37R����W�yR��$��� �.�$X�h���yB�
:wt5���O&	�}���,�y�"�����%�JDPr2���y�B�We
��̓�{[�A�Rm��y� :�v$"v�U�pA��� �y2���Gݠ�#�G�9E�q1b��y��p��X�7Φ [�E��]��y�-I�&�>�{��?}�R��PB�"�y�DX6&�U��;��Ȣ4,ͥ�y��Q�W����4i1e�m25�˟�y�K����mDF���5�F!�y"��Jj�p�L�;�FI�T��yB�Z�8�2��D�z���1�mI��yrO���<��ڛv@�`�ҧ�y�ɲ�>���+O�i+<�����y��N�K�(�C״i�`�$�y�ŏ}u��Hs)��st1��K�<١N�)��T��d��"���%�{�<��h��$��3c[�y�`�ц��u�<)���Pƹ92���U��e����x�<!�!��U��q{2+�g?~���X�<� M'2/Z�X���@�Np;�
�V�<�q���W����`@ގy	�\""[W�<�U�E;^ɣpnʜ <��g�[S�<���Ld(اe�T�!�.e�<� 4����ǰ���i�n&Y܈ɲA"O�){ 	�`!��h�� ?�FE	�"O���'08�#��LHH�"OV��ei�P�"so[<3>��7"O]�'CjT�i�oV�6�!�"O��e�B$>hQ!��L�)��"O���U��S�l�%¢0ar��"OƜSdL!�*5�2Ɲ"@��;"O���F��;�,�#�{��p�1"O��jt�T*�zAP��P9
)dي�"O��J'�9r��A�d��
�� �"O���B�z�l9��O,}2�-I�"Oty�
ԟ��-	7
 B��d"O ��A΀o.ԑ�
�mJ9�"Oji���{.��l��$�8A"O:TcF �S��5R!�����"O�B�		?�&Uk�kM+
nQ#b"OH|YU,�)K0�{I�=��1X "OJX���@�.����C�_�Lhp`�"On��Ɗ�����ZP�v��m�"O^�#%'����� R;=�mB4"OH ���
4
�ŋ��_���H$"O��SMǣ�H훳��E��A��"O��IM7`��HJ��s��̓F"O ��Df��a�&�8*�/>�
��"Oz�8E���|c\�)�P�#�Ip�"O0,z�%4�N�딁F-#�V-1"O�t�`��f`��&��3a�-�B"O��A�8Ъ���Q�6�.UY�"OduiF �2B�XB�C�2q:��"O�)!bY �#��#ik�d�u"O�Y���C�8�T��� �B�p8��"O��d��5*��� �!�2f�x��"Ot��p(ػ&H<l	�o��eVL��"O���B�G�:�L%!�n�s2|��"O>�"+��+j�%��A"O�8�BL�n퀱D�.:����"O�JS��>aȪ�sB@dj�R"O����V�8*"�2���c1�u8�"O~��E�8���
�*J<��"Op��e$��Ἡ�w��F��P�W"O��a��BєdRŧѸ0�:�!q"O	�CT,C��E3�*��A�"O������3A���m�b�z�"O�� ��1!��YqD�%Ry�z�"O�Ya�%a*aZ5 ��/QVY��"O$1K��!Ai�x/<&��p�"O�������٦lO�Ep�S�"OrpS��+��`�Q��;�:�x�"O6m�#��L�Lp�G�G�~��0��"O0���@	(_�4(���n�T���"O:mp�T9����J�X|2"O����5��p	@]9&'�e �"O�񺠤ޤuV� 0������1"O,������J!Kq��¤9�"O$���m�v�ha���Dq8��q"O�P�e��5Qr���J!'k��`6"OR؋&ϮEC:1ڳ�ޫJ�����"OC��V� ,[�])D� ��#"O��/�/�T��e�G�x�Aw"OxI�%��?\�r���9c���@"Ox�ch�Vq��;�b��tx��"O2�2��I�O�&t�B΁zs�r�"OF}P���E��M��,E-ag��0T"O� �I���U�wit�S`)*`!�Q�a"O<� J�;c�˅iۺr(Th�"On�2��U�.�؍��C6"��Ӕ"O��Z���^�l����!O�5{""O
H���Z�nܘ$�ޜ�*d�#"O�1�ʚx���"��R�,r�"O�IqQ����ƕ�Ǝ��l��	۳"O0|Z��dFx��Rm�#dL�`"O�<f��f�|����!Y
�+w"O� b�IQ��̜KRf¯k!��g"O��B 
�)��SD����!""O8��e�$��M�%�┸�"OnM�҈ Κ����!K�`�b"O&�Ңg�zchl2G`�S �0x�"O���NU�ް�S��`��i��"Od٘&a�
���چ%�f��"Oح %��Z A��8T���"O��kB�ͧ*1�JB')b��T"OH�Z�˱&H<��FF���"OB]�!oK��>E3]�H�[�W��y��I�zВ�#1"r�0� �F0�y�� g~���k���pd�y�H%f�~��+�r���4�ƈ�yB舚l�4�D�R�'I �h�����yRG�,�x�������Իv*�y�OF?�@�C��Ÿ������'�y�]�1�&P�-�A�PЂ�U��y�fX_��0�w�	#F�p\H�� �yr��	R#�[��$f�k�J�5�y2& ��20 ���n�`������y�G�:�6kdg��r�Nԫ��y� �?a-h�"�n=	����L��ybLޭx��$��,ܡe�
$S��D��y2�וX_a�c�O	f0���j)�y�E��~E	 L�Y�Ȩ�a�7�yBJ9Ub����R�Q�$*�Ӱ�y��-%�8�S!T�I� ����yRʊ�E�`���E�8�h$)�'���yB���*M���"؊5!`H�t�4�y�$1<k�u��Q&�A�MR�<�e��|)�YS�e<�l�`E�j�<Y!��E6(��#EJ1�ĝ[@�IN�<)��!Jܫ�cW-u
������\�<��㛘.zX�'#G(j�&��a�2T���s���T!�y{��Z�Yh�C-D��[B�Ю2^)�'��:W�Pa�g�.D��)ԫڼ�<�C������[0*D���US&9m��x�L*8�����/D��z�I�SV����鍢7���6n-D�$k�@�=�8|�fF�Cg�	��*D� S�"�3�P]1@c�,0ؾe!��,�O�����Y1VQq�L�W0a84�Y�w�x���I�AU8G�쁕<єM�d��p~�ծ����'���Ö>�S���)��+xBmc;�&��u#�+i�R}���֟4�sHB^6�����*�a�!��|x ��*�\�jV&G~��I��ǧ1 �=�B��*fdp���/G��� si�*�s`�;H���z��ψ2�T0�¼�?���(���jwiɣ�U�0 C�k�������.v��8�������&K�?Ya��I��	��� aꀵ��M�E�H2�����H���\�J��Y5� ۉ��tnz݁���(eN����Jղ  >Y)*D�,N*�Z�Ě�V)���@��	�7�豙����Z��7�
�"��Dp�^	��yY�)|"�T "�O� q�Ƨ�.k*RH�q��F&l��+P'h}麶ńfLEpD�&�0|J��;;D习�W�r���E�4 �尣cK(�x�	�\6M'?��|rU��c%�ة��>pp�]q	ԳWD\3F"j�E�.4+� �r�'Dd�qP�J�{8�� �%PN�JT�{�b]ac/�u%R�$�)�0|� �p�W"�!D��M���E�U2�Lˣ�J7|$@B�I�Kۛ�j�ix��|&�,�uA�-)FT�!7�:�>��D/D� P�-	�"��BN W!Ģ�)/D��R�ޚd��fI�x6��(/D�����ք��c���)6��XkM+D���ˇ�w�F���$Z	�Ĕ:ҧ*D�pq�����e ՎY��@6�3D����DR�A�U	�ȶ.�x��$$D�`��3uh�X
F-�D��B0D���w�&d���C�53��!�-D��Y�#��{z�L#k�Bd-z�,D����ʩ<��Ɂ2��"��ej A)D��Q�E(R�<A�����XH�yR��,D��7j�]�&���&/`��� =T������G���Θ�.xT$1r"O�mc�L��R!:ҳ�I,\�h�B"O��7B OWvhg# �-�<�R"O������xB�٥C|�v�5"Ov��F�H�4�؋�^�q�b)��"O"[D �%x�p�5��8�\�0�"O�r��+V�  �=��r�"O\I��+���d�Hݙ&����"O��c&��$�TX1��5hV�d"O��Qg�)B�(Ťƭ_<�k�"O��`���4mڶ�S�-	68��3`"Olb��; a�UPq�Vq0<���"O�#�A��/�	�@�%�0�3"O�e����2�)\8%trQA"OfA3����&m�%�@�}����w"O0I��G.H��"�m�#�Q
'"O�����h@���-H
3���3"O�z���K��V �&��"O�}�0��Y��Oa�t(�V�<�� ��r<�f�8.8��f!Q�<��N�ȼh���6V���3�C�<!�ݸx�\�'d�V��h���f�<�2���(ܱ��ݘy�����_�<��;��l1�dL D�4�Y�H[�<���ԢB6�@�%勼2(�!���Z�<�'#�>��E�xZY�rCDa�<���ϔH��d �M�7o� ��b�a�<�����W^��j���1�\$9w \[�<�ţ\X����6��*��98��
Y�<��R�&s��U�1�`��Pg�I�<�F�P�U0I!O��$@��0��E�<秒�Kj�B��̾	D��MA]�<���.Vm�=8���;j�@��C�[�<V��=4J�PeMI5&�`����W�<IfڛA�t)�3и0bi�^�<��΀'���H�l�2O���d`�T�<	p-7xn���嚬gd� J�KM�<)�m�Ơ��	�����L�<�wm����\X�)CC�$�P�VJ�<Y��ВM5��S�b�4p8��Wk�<y��A>]8���)�l
���B/�k�<yGg�Ny�0����5z�"� �O�<�@�-}�p@���Z9A5,�3�N�<Qӥ��<���ԃ�3L�+G�_�<��Vf{��&)�h 0H]�<�FD�o>Ta(r��2��*T+n�<I��H=�d �'Mv��aūV@�<�a26���	���Sԧ"D��3+L�e	J4z�e��	G!D�����`�:���A�ڐF?D�� �:Q��t�8�叚w��djw"O
!ؕ��Y���k�B}"�"O��)&�+*�a�TB�	?����"O���1J��8��d�W?%3윣 "Ov��� ՜_BTJ�o�tyE_��G{��I�L4pSʛ�^�2�`�Gĸ0�!�dםT�Z�"�W>n0R#��l|!���9\ T���+7>1AO\!R!�d�)��4��ɘ+0����ݖI!�$[-#���Ia���9��#^�[,!�$�i���ŧ�� tR�P"!�%[tQ�e�����E@�;o!����5�w�C��"���K�$I!�$�y�	��ύ��ɉ�HPq!�d̵z�΅ɧ�r��8$?P�!�dG%P����n[�N���p�`T!�U�O�p�q�����ъ����!�^�Pu:xX�� �@�ԡ��N�!�d��zT�X��p�R30O�	�!򄕨8Wda ��
�~sp4��� �!�dЪf��A��!��gb��8��3!�DӸ;c:��@*ԡP �|*���s�!�$<)�5Q��ÑK�lHz� �g�!�D�NZ��Ц�	�v4Ce��Ll!�dȗ6N�n�$���i��#%�,a�"OpD��"Gۆlu�]P��B"O�2㤍�U��}R���y�a`�"O�g�V�l�ݚ�eB +�H��"O|�ӔK����Ԃ�#oƘ�q�"OTDz��m��|�t`$t����"O0���-���ا$H 3�����"O�P�I�1b]d�*�,v�X�{�"OZ���`�JNX�PB�,dx`"O$�!�!�=%�,���`�kcf�F"O2 ;p�G�q�Beؔ	ʮxZ��0�"O��B�
8��AS	�A�e�"O䕓f�2h�c'�J=x���"O*���n �~g�d @��{�P�0�"O�iRP.ƻt�`j�L����j�"O��B�ŅI6`���B+c$�3 "O\	�X/)�f��l��;Q2 �G"O�qض�`��p���E��F"O�ظ��R0O��ܩ��ϞD��"O� ��.�>�D+H�61fjA"O�s�OS!]�D-�r �)�u �"O�)����$=N���Ǚ�J� ٻ4"Oȉ��+�JNpp��]�"���"O�U�dc��j��& ��>쑷"OT�@�(٥E옭+�%ު=h���"O"�j�"]�u���5�ç`&a"OqŐ�*�~��NU����"O@�s�i��
�Bz�T���"Ox��1N_�O�<���_�H�f9��"O�@�%
ҥ(:�<�&�G+Yd�+B"O��k0(ƎN������M%;0�`"Op��SȔ.��E0 �'905��"O�*u�ͤ-��H!�D�^�c�"OΙ0� �XҊ@8�EV;Lr "O�¥�S%P��##J�'��L��"O�$����#\���5HA��h<1�"O�����7p�Ή"h+n�a"O(��hT%x�.呀h2gDh50g"Of=��
�;O�Z�(\jL Pa"O�|��E;M�;�kɤQ*���W"O� ���F�9A-L���k�/J���"O:� b%I�0�N\qG
�h��1�0"O��ol���+S��Q��"O2�SF��H7~��$%Y3;=&x�"O� "���)dU����4��!�"O^�R� ֎?%�u���w�bW"O�0ROƣ��j"+"e]���"OJ�{�-߳+\��4I�"H�=�"O��bv*��P���(�I ���:�"OF���ҳQ��"�׫;rޝ�F"O��uE�=����	�#TcZŉ�"O�H�5��7����6c��[�"OxXb��PT���ED=N�n\��"O�m���d�V���r-�"O�CV�L
i��ģ�ִh0l[P"OX4���� �l�J�O��z��"O�񴧇�A���ҕ���-��S"O`��VgL�=( h֪hPyK�"O.I$�!]���z�f��0�%��"O�|QT�Ҩ!�n���%�Cl�Ƀ�"Ora� � \ԛd��7����"O�\�$�J6�����/R�D�5"O
�C�KWS���ck��9,�9F"O��@�Ղ@V�}���ҠV�2i��"O���o�7;�}�DȔ�&�,k�"OB�zŋ��S� �(�H`�!�"OR������ԡ��ϒ����"O��%�J$@K8t�e�F�Ξ��"O�����,z}x�c��Q����"O|�S�7.N�����1L}>���"O�t4�J�#��H����y[�Y"O�@��(K�^�X�
Ѳ=ȁ·"O�ALE��Tp� ��jVXT"O�Ā���8��D �� ����s"O�U��F�!1��A�o��D���b�"O|�qo	t�VL�S�:9hAR7"O�;5NG�He��RaOoQ�,�T"O  qD�eӆ� �Ӑ	A����"O��ɳ���+}���-��U�P"O<|�D �xƑ1�Â$(&�E"O�!����Q�VxiRCX�WAh�P$"O�٣LK�?�\ u���1�,QB"O�u�P�5~&Q#� V0Ms�"O�	�V�-P�)X����>�� "OD̋��+����N,bޡ�"O�M��ND&��qB�m�
V��1�"OV��)�/S\
��)^�9F�<9#"O���nR�2Q��ä���f�T�z�"O� �C���B��FÅ
�ɀ"O�H葈�E8�I���n3�EK'"Oj̚c*�.����`χ�)8���"OPl�QI��|Ap�x��?<~�� "O�|�1�;Ɛh�
̅Su�Ds�"O��A�Z�,���R1oP3`�Z�!�䚉m=
}��`\ ��<���B�!�DC0I[vQK��܋kO��Ŏ�w�!�LD\a*fk�	;�QX��F�!��](��0��T�=���*q��3l!�䞵j���0è��E|\i�k�<b!��NyU.љ��]�M�H����DO!򄃪{X��#%%'���Q?X4!���4wR4j��1=
�u�N��S!�d��]�mx�BQV�0yU-��!�d�O���t�$g�2%Rd�$	!�� ����)�!=Ԧ���S�Q|$A�"Oְ+d��m�|��hH�:��1j "O{�,J�Z�lt�۬9\��"O(!ݛ_0)j���0[Z���"O�hB�/!��I��)Q�?D��cr"ON!r�Ŝ�EZ�M��A!�5��"O22��Dm���ta��i����"O��;$-��b��\҃)�_I�ᛗ"O�R��B��JDb�2[:��s"O*��*�,~��å7FT*��"O�Q��V6�q�&�,42}��"O�}�#.���yBVe;DH��0"O��h�����jd:C�I��*�`�"O�(	^f�����m��x��"OR-*����ei�a��Q��� E"On8�sB�/+�p��	U�FQ1"O�1   �   +   Ĵ���	��Z,t�E�=(���dC}"�ײK*<ac�ʄ��iZ�Fm��x"�
��6�Y�?5"�X�h�k�:Z���0P%��ނ��m��M��^WI�� ���	�z掅��ӟ`3�b@�)�����)Q�������^' �@�Z�|��M@H�H�0���ݡ1 ��81���#S����C�[����Iը'��� k����S*Us�I+�t-+$��8b��	$n`�L�RdҀb��8z���DpU��)Ӕ$������,H�('>9����ВL���_�ț��t�&(ˑD	D��&�>�*�����G�d
��iI�nLU`�K���$3Խ��)�,�Zh�ɁO�8���i���$"�0%��M�J��HxW(�s���A��-;�X ��y]"O��B��&�-�L���d�!^��+w"�&	�B9�����:1�b�#��[`��q)=�$Ɯ`���C�r>-�i@�ln�qye�U<f��2@����?�o�'=�N��dYjyҡ�5�H�bU��q�Ԙ͓�r�bd��&�����!
B��BvnD!�l�$�`�%-C$X��&>�vGa�6��p�r�I]�t�@��lūWg���|Q4�0֊V�ʓT��B��\�D�Or�ij�	��:p�#�r�T�Bg��� ��O@J4$Y1*��'��ءf�B,ى҄���p��[��&�耳i��|�F�OVd06�C	v��@�:�r5��Gʒ �hq����6%�&XX��!����O26d���|"-��4ގ1�ֈ�YN��s!�z�X��	r��I�?�%�<Q��]�$��
�
��5��Jt���j9��8V�Ds3r�i�NH*?B�Y�3i1�M�R/�3?l�1q��i���"e\�ZNy��4ub�yK�������QO�4�m�=y��%
��'�&��QFз*,��qK\<�&�����u�5R5�x2i�l1J@��y=�}H`I�&�b|��FXǢyi�"O�����  ��'ƩJ��t�� ӱP����OB��W,�{/셺`a�/�������}�xй&�~R��]�J�x�S� � Z.�<B�H�	�v�����E, ��*TKY�@�bWMp��S&��i�C�m��l�o՟_wnOj���'��6�l�O_�|HȲ"SIJj�Q��]�!�$�.2�XmX�S�T
T}֨��7�xB�>�f6Te&��y�>����ުm���,   u  z  l   �&  -  F3  �9  @  ZF  aG   Ĵ���	����Zv)���P��@_zX�B�W4T��,9Q ʍ;A0X�d������66�L�w�Ԃ��C9�@ ���T��'�j��"��Ԋ�i�NU�d�"Ea
��C�_S8}@(I*B�q��$�$.`�%�D`�j��t��,YY�pȥ���y�:d!�f ?,��xX�� �bn�9�(N4}.�c2M��+J�w$ϚV���d58��3��~V�E �lӆI����r/��%����dՙv�ąYE/2l��X ��?���?A�����-a�
-�aȈ�#�x@:B+L�$G�Up�ɚ-�b�+�-�#�$K`T޺#��#�V��~(�O�i�R	�U��H�C
.q��b�� ц�L�b0�|�K��!��S��UI>�©T�l���c�Б9Q�@��զ��I�xc���`�".���u�'�
�Pԯ
oF��g��U4��H&vӠCቀ:Ԏ�Q��"��@����o��m���ߴ�?��'�/�ؑ���Q�J9��g�<i���Q�J��)#@4���O.�d�O����#���?�O�x\�7�=e���SU�-F�~L#�L�����k�aI�o�X���)	���J#,Fe�'���#3�D$X��h8e/<�b$ �O�?�n�`�i�HqR!h{�X	Q
G�'��q�E�­���}� �:d	^�%��0#d�i�2#=9�����?`\���'S�:8���ɍ[]!�$�73��%!���F���hs��EK�ɷ�Mc����ӥ ��1�OV�ܟ���G��<���K�5<��"@�iJ�����'���'�	P0B׳9н�u�?-X��z&&ހ>x����ǝ(�ά��aː &��@��(O�� r!J�8�,§�Ƌr�\(��Y�(
�����i���#t�
�u.be�E��(OPXy��'�7�U̧ ��T{��|!�0�`�;x��'��~"� �~U��;5��)!����e��6�>A0����Ȋ�$�5�qcI�o튄C%�>i��F����':B\>R�i��X�	8+
�`U�-lX�C�b�"�T}hߴ��-�RC @���&���{�l� 3y��ĊS-��c7�MZ~�#�#�E��)ӦB�ę���(V����09¤�O�'d��i�E';yL�K2��M,��xS���I��M�WS���f�{��q��i�U� ���"&�eS�'��(F��?
���2��	*Ȉ����c�O<�%@.�.^M�g����X)�)k��d�O����$�!�d�O��$�O�Y�;�?����3�\)BĢ� ~i��U�F�D4�1�э�?�Y
��>f�,��U>��t�����'�>�(�z4��1��{�P�a�W�	�8�V�RҒ��	I(��Ԗz��:M<�FQ���PD(I�5�\Uy2���?a�i��"=��'5<�L��pGN����-6���
�'���0�4�<��H�(	k
!�4����Sßt�'j�27̃�d:l`p��1!ێd��ʔ7z�k��'<��'���i�)�	˟|�'{���
A-�=��%s�
�%N:x�� ��h�r/!�p�GM�����N+��\H���4&`�����"v�������Bi� 7���4�b�0Ƃ�/�Z�<�B��՟Ԡg�\hT�:��R�ѻ���M��	|�']���gn�9 ?0��L<ȘQ�'��]�U��<:B`B�jܹtr|�O,nZ�Ԗ'Ū�a�~�������5(1���C�C�F}���OQ��M����?i��?���~XK��<�"���gӿ5�u��g�-���a-߷+{�<�r N+kr�dGy"bF�2�tXj+[&v� F6Pd�lP��b��T#vr>	;�(yW8�Ey哙�?���i��b>](�+��Ù�{\���'%�>�	�K���+焑T���$NP���	���$�P}�\چǗ�9R � �I�e�	6��Iџ��	x�tl�U��'��:$��vހ��ɸ9�������d�X���5w­V��G�RlJ'��E�T�X��1��OQ
�M� ߊ��%�U"�����L��pq�O�HT�q0& "z$��ˍ�7�q��A�F�8T&�|�$G��hY� �f�O��Cu�'*�6-@TyJ~Rʟ��yT������
#�����(D��Q���"0��]�bC�uטxR��9ғP0�?%���5j�Pk��E��"<#�G��M;��?)s#A�5eL[���?���?�F��t��ǚP��gKW�;�})v��$��LhVo[NØ��lSb���H3L�_��	�w0V]'��Z툧o#�8`k'�������%�D�SU%�	��$���xK�'Ri�|ca�-�5nVx:�E�~��{�瓄/��I�)����ߦQ���䠟�YZl�@�mD!%��@H��)J}!򤖪S��q���;��˴R��e?��|����.K�r� A	i�H�q�*H�+Q�l����b���O��D�O�����?�����ġ��?PbL~:q��#�^f�p�1%�:R�}B���~�\8|��j%A"鶜br����>Y2�����m[��&D�$�"θ�b�
^��y�k�5�R=�G�[)GK���P�Շ�y`ܶu0r�P��׋B�beA!o����[���$�̓�0�M#��?�O��r��P�j���A��Y�t7����4D2���?��\����Ø����<֚�P5g��~ژɱ��͗�hO@yP��3� ��8����	�>�`ҍ� w�D;A��1?�d�z�O��A��,4�@�z�A��b�����'B��$h,�*�D�;X��{�	O��( N������*��@N6*$8�U�!���i��'哥s:)��˟��N
}Ҿ,h��?:6<c�����M�ѫ׌�?��y*��O�k%�O��P�����ڝ��'%��Џ���l��$�̀q��#�D��D���ɬN"���x�)�'Zݤ0�3 ��4�D0��4RV\�	�'�����lI�.��Eb��T�FDh<A���]�O&$l�Ei	���/\5|#��8��r�F���O"l�+�2�8���O��$�OZ���Ok�ف�����j��K��U�"��:��I:N�����C:n(z'��iGL=d�tx�I�g�n��D�����SCb#mվ	�c(O�b�Ɉ_����^e��Pc �}R��t���:7�>D�l�W��d�H0C���2Q�}�tEz�O��':\5ʷ-�*MK:�a%cV��R�c$�U�0���'��'�"�}��I����'uN���	�N��	:6ڸ0����D�vҸ��'
(�(��8��G { 04����M)N)��		O)B�dQ|0&)i��H(Z����-m�&���!�z���%W/z����II�f�^I�ȓxS���%@D�+�.��v�5iC�$�'��6�"���:!%��mǟ���GJ"g�9|l	C�Ř(��27Fߦ]�$�B�0��ʟ(�a������<��d/ !��ɔ^�d�@��E���D{����
=�͈�xM8}��!BS�d�I�@ϰ�$�W�O�&ɪEk2�z�*�IP"}��	�'�*ѻ7�Y�Fm�K��S�(L��	�5���"�l�[�ɕ�*jFy�.F	o�N�]�P�#�i���'�哵k����矄����Nn����HQ""A�Q��;�M3�϶�?�y*��O�40�ꙙ=f��`�ZR����'�@)����Y��`�(C zep�qCaV�]�|��d�>��X�)� �.ȁ�I,Ic�km��:2=9�'�>p� '�nQ�Q)�$cvxR��$L]�O�� �ǐ!II۰%�&	xT�
ds����O2�i�Ð�p����OR�$�OD��;�?�1*�0�S+"7�X��%�B��LoZ�@��BK�|Kn�YA���0<9��� ���1JD/}y8��E�yWn�j�����0�ޞZj�ؔO)�P �OW≫�H�n[�z�����dN(�|6��O�ecTO�O*�m��Y���IR?q!בJ�!���1��@�b�'>�x�	۠�4âɝ�'".�X��M�ði��6 �D�R���<9� ^�NLdۗb^|��QY㉡zJ��2�O��?i���?)�:^�n�O��D�O�1HQ�;�&u���X�#�A⒯�-N3h�c�G�Z��P��'�2}
�ܹtLx#O ��Zy��J�����;&d���d'F�A��yY��gљ��I�
�O%��+�̚I!�k�&b9t
]צqsM<y��?1������(�	�����'Q�cQ�j`�x��'��س������R��Їw���O�PoZ�M�*O�,0'զ��	ȟt�'*Yؘ��I)U"���p��Ao4i�����|�ɹK;jВ��Ȋ7r"�{��Z�����#�]a�i�ի�0�	)r�_�hO��	�`3�Ca�����A����1�0\;"�qf��h��[D'�$}�
�0��>�f����"ʓ[h,������n�@e�!C����BA�<*�E0�"O��!����'@�!�H�f�F�;`�'2��2�0�P���$�n�.[LP��'�4��aӴ���O��'wr�����?I�l�	�F9�ᖔ$ZR�i�OH5fq�&���l�s�G������C*!c��'��O��$�!G!v�4Dh�Fȓ_����C�'K����N�el4d������ �h�0h�j=#��p�)�+LCl�2w��O��32�'R���������,SwM
 gԔY٢��u�x�qV,%D�̙�̿(U��S��L ���#�I�?�sL�X��E@���m�rIۤ䈋�M���? �K9�"���?����?����^��,2�4���('��˖��[%�= #�(#]|j�G��Z�$���^�4�	!5�1�WZ�6Rt������g��S��D�ޙ��Ú�o�|i��|��V_�d����)�k�9��U;,OX��E�'���'��O:�85��9`���R��a�bH�:n��B�!��	:����ə�,jwf6m�I�����'��!U�VH�֮�Eh|E�3��#p����t�?r����	ȟ����� �\wn��'���@$ ���
x��`���	j#�U�f��5!d�(��M�*��0	U��Y��b��d�5  ���d��:gR@�,�B����T��7�)C��X�(��,��~�
}	��DЖ �2�:� ���J�m��P[�8u�<��"O~��S��1��rK�M���"O�iC��t���a2LT̰�*�W�X�ڴ���`�� U?��	`�5�� 8䘪��C�}�����Ňئ�	���ߟH�	䟸�a-��&78@ VA_���6�������"g<�R���U�����O�hOj -���b���  �IQ Ca>-��"�18��,��FR11�$�2C)ړ'�d��	ן��}
 @�!�dK�E�_�@ �B��X}r�'M�|"��3� � ���	�`�����o>��.��L���)r�*��7k�($�GN�:B�i�R�'��S�u"���	ޟؓ��T�A���#��G�K @N��M-_��ب���U~�HiD�4@�4��С��O��1g%��yo���S ��4�'�1�4 !9��Hv��dl�,8�#ׇC�)�}��C�}�H�E� 2�÷��	�?i�G�˟���C~J~����~�g+�`1�K�=4P��aߺ�yr��)f;3��Q��	,�HO�D��l�J�]��M�?��@��松r�7�O\�$Ȇ�i��O���O�����c��(��!Iq�
^�:�  �m!�a���<8p�O5*��u��1��Se�'B(BF�4O^�-��b�$:1��b��S��ŪԛxAv�q!#٨��);�L�T����SD6"p;��G �̖'Bٸ��vaz�A��c�� r�r58A�+C��y"�w[`Eʬ+֥��+m��2�4f���SW�8dt�p��U��;�#s���/I��TPjUJ֟�I����	��u7�'O8���3�$[$G=&,��+�~}�� Ba�8kՂ4)��*&��X���}�1n
�Q��ir��blj�+.4�j�S�o\0��	�G��B�����Z�e��pشUN&�<a�dџ0K�F	+�ݨ1�ܴ:��7�;�y`̌R�sgNפ�<�Ai��y��N-"t�U��h�<�S�P��DӦ%$�$h3'��M��?��O���õ`CA�t<��C�/+��"ݴ"̢|P���?��X��
����<�m� F3��3,ߩ�"$�+G�m�E+Q,��=�PBA��y�'�",ʕ�JZ�D]�����<Xt����Tд��Ɗ�65�D�;�k�m:�)���r�'�b)��q�>`�I��4	5����ub�:D�X��I?T��AQ���	M�F�y�N,�Op�'.�H��hǈCP�R��֏�ʪO�V����I�L�O��E�'�"��,R괪R�@�"��Q��ƛ(�v6M�a9bHW��/z��r�%�Y��@F#Du+rc>ձ��+<���*tD�1��hkӋ�ȟ���l�tg����� ��V�2�S�B�*�ħW�E3E���)V)L�d'6q���U���	=��S�O&>0icm΄.x��+抂�il1��"O� ��M�?�r������"���>�ȟ$x�0ə��$F]2FB@Kgʒ����Iϟ�z�M�W�Dm���l�I럴�^w�Zc��؁@hX� >�i��l�&�d0y����?�n���eP-�Y�����I*)�̳��4�
 z�iÆs ����B'"��qX�O�a���9FgA��I|ȣ4-�5��i�'b����jZ��O��D#�IY��*�G�PГ��J&4|���c�A�<UML�D��<�e�ϛr�����u��4����<b��#w<6�ڲ��	Eq�\���Ɠ���Ѷ
X/�?����?y�C��N�Oj��n>){� ]�{�h���G��❁~WJ��s �*8��ss�W| �Id#	�s�؉�D�$WNyr� |��@D�V���;Ro�k���`G�TD�=!2�=���ˍ��\��KUR�؉�����s+L�Y��4�?a���s��<0�ipQ2����r,-�W�'�Q�����Z�m� ��C����2����>y�iE�^�Hs��Mk���?��Oɒ釨�(m��(�a�Q,�����41p��s���?���J��Pa+g�.�ݴV�����H��eВ�
$��``O�!�iА�۲wQ�0ʂ�R���Q�i��&���S�[).� W@�7D����ӏ��d>� 0׈�Db��2Ǭ�f�ɭEbZ���⦝�N|
��Y�[D�!i�e�fg��KS��B���'f�'�"n��L�0-a8�ҁ�֘.����ԑx��i>m��4"�"ٻ��Y�!ȹ|j��ڂ���$�"�*�	CR�i"��'D�:ྌ����������A��EX�ކi���R	�Me�Y*Z�b�{��_�7��Ѻ�8kt��"�+��O^�^�P�Q�a
�r��-���'�0%pr�ؕx��t�Қp����R./��e�}��ɉ+	�eP���h�����?����ǟ@zH>E�t�A;��=�6JD�pe��;�'��0�!�Č�]{�b2 Cx�9�f�+*ݑ����I��4r�iv��2�e�E>y��To�ӟ��
nܖ k�Jٟ��Iɟ��	��u���5��7*}�Sií[�>�E%�.m~0��\�/�,���Bs 8}�-�t�3햳�ē����t,��o�J$C4B� k��4y���@!���DIr�s� k��Ȁt�̝$����G�MU���Wu
���ʷ<q�j�͟���S�? �l@�`��V�1�	:?`�A�@O5 Dܼ[bU��o�iD��a�#�ʦ}`��4�`�O��!FԬ.�+ �\�T�\��g�R�z��ȓr$���	
'q�h@8����*�������c��͐[���a���&_����B�Hq�
�� l��n'91��ȓic�՘�"��<AȬH���Wئ���d�ڤ�v�ݵb��@BD@�TӰi��Ia~Ѱ��
�
XRT TK��#�r�ȓ}ݪ貥`ړp��e��7�Y�ȓd� ��mƖ��ͣ0
ˬ��ȓQ�8�@J��H=8E$uJu��;�Z��Fe[k#�8�0���h��}�`HǨ�yTB�!!$��$x�,��X2��*��o���mF!O����ȓi��b� P�; ���	�b��ȓc�&-1�g�7s����̊+{<	�ȓ@;���p��$�Y�`֍'��,��~�2�p%,ס3p�9��'U�_;\���>{��$l� <KTM��Jֹ]b�L�ȓ*Ƙ}�G�To���p��	�����l2�ࢍݲt����Áf,���ȓY��)J��ɱE�8�4�͹t�̄ȓip���+4p��y�@�%X��ȓV��IUb3@~8v�@� �ȓ?�H8�6iO�:�fq�sh[�;(�9�ȓq,B񴩉�f.��g�ܒC����ȓ�P�PI��z�D��ץ�`]6<�ȓx��VoZ��A�Rş�`��X��d��؉2mӅF�8���[�D�ȓm]�e��aD�����U/Nl�� �،q ��s
*�p���>�44t �.4�`�$~w���6/��1�B�-[����ڴy�橆ȓN=�Z���I� �x�(L�}rL�ȓ�!!�,ɬTq��`'g�8���y���G���F�`�j�N4��+���x&��4�d��S�H�W���
�r�aQ$�H�\�T�9+���U��y�jё3g�+�.Ƚ��t����Z!�_;�eG
^�)�@ �ȓD�Y�ɚp
�mv��{��~�<A��Q�v�RP��L�/L9c��Ls�<i���c�.\��G;v`cb��w�<1`Mɢ4�hD�ӆ�IΞ�8���Y�<���*�R9Y�[=��(*@U�<	��W�<�ܙ�͕E��Yq#�o�<�0�W�!S�)حd�Dk��s�<)p
��.rp��(B��0ᩙj�<Y1F�6��$X�C!��H��F�i�<$(k�6e���M!&�
��ǤRa�<9���aw5��� 2b�CA�Dv�<Y"a\>t)4CDjɢuL�i�A�|�<�V-��M��i�f��uϖ1Zf�{�<Y�%��N�S2Þ���c�O�s�<����O4}�$U 1)�d�F�NN�<�R��M�����!\�D��Rc�<!��V�`L�R�F<2e|졖�F�<aFDF0��re��4+�E� L�<�&_�Z��3H��B��!$I�<�7$/�:0+۴$�LC�) ��y⥜�^\�ʆ��9k��U-�
�y���v��u����`�1��	�y�n@�b�0U�����@�G�ւ�y
� ��3�m��tg�E5HӬ	�,���"O���G\̆�%�� r�4h�"O�D��k�5pyl}�kѴ�C"ODm#�2^����L?��3�"O2p�uG��P��HH�n�>��o.D�([�G�xj�Qb���q8-ZU�>D�,r���*�8�I!��;� ��d(D�4��}S�-�׬�,j- -*D���s�#���s�72M��r�B6D�|��l�*A<�9�a�
ab��j�b1D�$`��
U�)�&�ɣ�E	V�9D�x�FɄy�|���R�~|8�m=D�( ��#Z���*փ�vL��p�� D��vN�=A�4��A�L|���ƣ/D������w��!SPP4���-D���·{�D5A�k͓RF& �R�-D��R�H8�$邗*��F>Q���(D��I�χ�#8�%�E�Z�<��3-!D�@+%ʦNNBp�Ԣ�}��I#D�`Y���"TH��!h�4?���I��.D� �Mqwδ��oZi]�-@�,D�$,\\�re�#`�����zB�I�x��2��B�,� ���$�TB䉃5x(�bL�!P<E8�	��:B䉞	�K֡zA,�*s��,���"O�]X�i�vhp-�� ��/�ybe��x��e-��L�n�!�(�y�ˈ)O7��v��0J4��Gߘ�yB��>V2]�6��+^4@��B��yBL 89�uC�'�\<��W!�y��z����߁�P,� ��yR$�,+��2A��<�Pl�:�y�H_8 �6`�tk
c�<�rs/¼�y�L\<?�ވf��'��b��y"�+dzE���U�KQ�]���X��y��ȓKiP0X,��J? �J�l��y�e�/VɌ�À�-���$����y�)Wk��uKg��zd�k��V�y�@�?Ff1��'Ǻ**�k`a@9�y�&ר�xyPB����c�/�y�Ļq���J���Vd������!�yb�K�}��	��.NRD((�C��y�)S#��$/ I����K�=�yR*żK̬�s���E����݆�yRH�gʹ�$��A�	�猘�y��ٕH����ͯ|���Nĕ�y"M��I>�Z��ɘn;��Q���y����	;��*�
g(Q�'��y�	\�*Jв��E7b�j�[t�N��yr�ĕFӬ$��#q3^�*GKҹ�y���
e���&ENi.�E��\�yB���"@Z���������y����X )�B���V8A4�:�y��̇or�|Q5BW���XFH���y⪒(
(r� 򣔔#��d��bم�yrnL�^����'h�.T���:����yR"!u����@� ��9�!��#�yR	����2���'X��UB�����y�ն$^X�Z��2O��1Ӱ'N��y��[�%HP�K��B�5�����V;�y��хn�]!��W�e���s���y�g91GnD��m��!Ю���y���;�&a��m��Z`��hO��y�����р->#,$:����y
� ��d�҇k&�@F�&Dt��#"O���L��U���s\)e"OjU�M���!``�RrR� u"O�����M�]��$UbS�$��E)�"O�<���y�0L31L5��"O�:#(�-�0��eΌ=��*�"OREa��g�|�j�k5G�VY�v"Ovl�6�ԡ ��tb(��(8�0bT"O�3�a2;9��0�̙:>ӌ��R"O�h���0AY�B�C%j�1�"O������4�f [Ck 3Iܥi�"O|���gѹyx�+�N 6R�T"O� �f�%�Uף�IEt1�u"O��Pb�2��U��G
7�H`�w"O!+t%@>e��a��Zh�N�Ҵ"O6q�*�1���b������"O"aPCƴ-?�5�͖r�|Y@�"Of�h��Qx�,�ᅪX(0���"Ox!ؗƁP��c@�5"#z�9"O�Zd�7
T8�"P�͘78���"O4Y{���~,���G��y�Y��"O�MJƇ�f&�0�$�yuvir"O�pgMO:��Q�$M	GR*h1D"O2��$̟�&�X���!P�$���*�"O (�a	_�,����Eg�&����"O8C`i���q1�e�r�L��"O@�x�&�H�\����M,D��l{%"Ox8����1�N� �+ϟZ�@=��"O���Pΐ�N��tۥ�D�b��1CT"O&�cH�'��1�#+F�?O����"Oر��ͫl�̨ȇ���<�&���"O�� S6��i��Y�-;���"O�䓢K0$l,�[���+.��"O����Z�i=�ٙ�El#��X�"Oz�B�܌o�'��}���"O�YQ�l�r)`@��X�*PEq�"O�D�Y�k�'΍J��iTAD�C�!�D!Ԉ9�A�,:X��Q�Up�!��N�E�����W
&�fZ�HE!�d��O���N
�fh1%%K�m�!��A��зֻ[��@���!�!�$I G��]�a�Ӻ^$�r�
��!򄐼u�	�Gxm��9A���L�!�ėx�qrGjزST�a���@e!��S�(y�$JX�(A<Dz"�<A!����DtXp�(	��8`#GB!�d��;�
p(��ۙ����Դ�!�9h���@0N�"}8H�D0�!���O <����Mz ����ٌ�!�O�t$M2�b�(|0q��,� H�!���+ľ���䑯�����l��ZZ!�D[T��98�R�7���@�İn�!�Ė;=���ː�1�h@��?�!�D�8��P���m�8xB ^H�!���9s�i��˱"�v�Iw�Ρ�!�C:RT��RGސc��5X����!�=eZ�8��<�	v!I�]�!�$�d�J4�ŧ�E��v���P�!��G��|A�ƛ�Ts�u{���I�!�Ù�-�b��DR��f.�<w�!�D�3L\JYA��Ɋ9��9 6���#�!�ة(�����W�	��$h%m�!r!�
� r��Ti&t3z���@�)U!��@�h���_�|O������*MH!�� ��  �V�L�"�񲤅�X��PP"Oxq3�o��6q0�ءs;(y��"O]y��0M��%(�� �$؀�"O�r��v��lWiϹ��"O|!�eLؒW�8��2	�
r�L�"O� ���1ц�se����1Y��'K>)@������laa���~ے�X��e��B�	�C��1�b�2c��X �֧?�B�#�6H�m��QP�k� �B䉶 �N=	�KJ�56*�3�i�j��C��7?�h{��Y/�Q#T!i
�C䉊i_R]�kư\>�1�(�%^B�C�	�Z��0�J��3�.x� ��f1�C�	�x��x����x� d�T�ǢǊB��L�8g�?U�8�QH"b$B��xG�}%�H���8��I=4G�C��#+������U�,)��K�U�C䉘ò��3�G�h����q��0�C��4uþe�P/�	nh �S�V�|�C䉗a:��˅�o\>�!��%�$C�I�i�I2%*�3>���@���7��B�I^�|Ico��v��	d�[�B�e���XpB۾ZH�ɪ��	Q_�C�	�����˖/,��B�:tǶC�ɞi������<
���uj�'*e�C�	8|��Ʉ��*ΤMAPɌ�AڬB�I1e5<���IřB��m+�b��|8:C�I�v��{���#n^Ÿ��	��B�I i��ZV��=i#�yAo�g�fC�I�F����D����DD��(C䉄	�:0	�-�Ui�2S/5tm�B�	Y༩��$d��̡K��?��B�	�{S�-(׌�4[h��㠆�CF�B��4~ٶIp�E�}�$d�#x��B�I�3�4�g�Z�<L���ߏ`��B䉧RsRg��m�A����t��B�I;u����Yb����gc۱)��B䉴6�j�1�ͳ���2���,x2lB�INI4)��  )uP�Y�gY.c�RB䉳y���ps�Ƈ�d�oP�$B�I;'�7	B�@;��3��u�ti��" (@@�N��Lc�Z]�<̄���]Y�m�9O�n��gJVy�ȓ4�8�y� �H ���@O�V6vͅ�a��L�7'��t�x�
�.RE.�����I1擐t���zUE� b�����\!�Ü�"���vM֓q3����Cej��T�Φ3�^0K��bH��&˂d#�Z�j�N��D�'M����P�$5k��z�D� ��#1e Շ�=N
p��Ρz�*̠`�M�\����=F�M���; �~ۅO�{����ȓ<��`�H��!X���k}l=�ȓUhn��ԉ�>�^�� �=a�����:�h+� �	A�1�&Å:r&jy��M��y�.O�=���
�ř�=F���7Sw+׶A�ǟ\�r��	\�<Y� ֋ +�1��(ߝ�z��;T�P��R h9�}�v��6����l$D���̏Rtەl�R+�9A$D�H����>#vMqT�F�#"z5�E.D�Ĺc��3�r�+��2�p�i�-D��+��ϷWwNQvOֵ}�"yۦ`'D��2'K	���#Tc�m��[�G$D�� ���0-D6|f��Y�a�c�
Qp�"Oq0t�OJ���B�I�`#&"OP9@�H�::�� a�[̓g"O���2�-6�l�堎� t��"Od���@V�B��4pү�!����"O&�9�鏸3U��r�/�=S�9Xw"O��c@�*ސ8�QEW�q�$"O��cnA~�4x�%�&2�6"O~�#pG<5����A�"���g"O�$��l!��S��~&�Q"O�\(a�݀q&�@��G7���a"O(l�1d�~�E*#��!F��"O<�v�O�!���#WO:�t]�b"OJ��"�K�\����J���
��W"O|����Uut
���SL�}�"O���W/�cڲp���i,���"O��)"EH�%��B1��,2'�4D"O�ݲ�g�?Jޘ9Q#R2�%L�y�H�:x�yr�c8R��"�²�y�GȻS�,��iJ���&��yᓯa����I�<��a���yҪ#Zz
��vf;J��P�+���y��I*�ˠ#�+��(��i�=�y2+իB��t``m� 
�#��"�y�J�%w2��&��2~��ItD��y�K���*8�NU4 ��8� �'�y&1з�2<��Ҡ��y� O" Z�]��"�=����I��yR��G�r���E��C�T0�nK��y�M f�}�G$¸UΠ��BI��y��R�$q��a�X���E��ybbO�>��(x�Ǔ�yv�ej5i��y��0PF0PsA�	�H��@�T�_��yG�%/�b��J�?=>��6L�y���N���3&Z/`��&�J?�y"�'�r��G,��!(ph� �]�y�́l��)���8�`���y	� X�#�U6	8pؑ'A���yR���F��!��Q��m')ѿ�yRc�2*�A����F������y҂�?����$���b�b�Ѽ�y���8I�
�$��yWF8Cà���y⡆+k�:���b�D4��(Fص�y�
�� ���|�L���Q��6a���h�A	|��բL&(��ȓ$?v̓�c��R���G�n��!�ȓ=�29	���73��h�0D�p�D��ȓB��
B�"nü��͙3��p��L}˦K��p:�ğEK�-�ȓ�)pV�[f� �� ���27���ȓw莰*w&:<M0�K���?h2�}�ȓ��D1��)%��*EA˅H:�F{�'Xl�1��+����C�� ;΄��'O�Dp���&jBh�!P�ss��k�4?.���^�\YS�ǂ�HY�(��L*N�a{.�B�	lѐQ0!�ʽG&���@FS�j{PC�	,Y!�E���'2����	�$��J�
��ا�'jO$��M�<Ynћ��7G#�Q��& t�sl��:H7K��{- P2��N�/g(�|�'��T��@2y�4S4T\Z�y�'��=��(��y��tXf̘wAIy$�W����nZGX��Z� �G8�eR�G�s	`��E	/�O�p�۴��$И:!����M��ڶ��9eG!������g� '���PF�ɼsў�yaC-�g�? J�{UKS��%�B��j��"OP�#�͓	*���4F��d��XB�OP��<���O�³����e��ۥ'��"O�=��с��I����'�!�$K�df��u
D��=����,m�!�S��R aÂ�W)5���Q^�!�Dݍ.�4���N�I)l`�r!�!��=y������m��	Q�ת^!�$��@d��&³E��б&Т+)!�D�,Fa d��ܱ#�P��Ug�`	!��8hK��̵����O��!��S4ƀ�R��ܮ!���VD�?'�!�d��3q��Js��Z�Za�5e&	�!�d�h�>M(�m�r�l�9W��8Q�!��L(�2��A�S�X@C����@�!�Dچ{4�腄 �r�����"�V1!�*C:<h��ʵU��}���#�!�/b�B�2f��T��p�a�,+�!��8k}�Hj�+L�
����P�W�g�!�d�{�L2�-)@�Io���!�Q!u[�����N�?6d�.¶:9!�ïoLI�f׽<*�8;��VE+!�䆏*ĆD��b��M���p��Kx"!�DL7�bg���,b,qĬ��g!�7xr���Ҥ*Tqb^:Jf!�B-�X8Pn�E�Q�a�Q7W!���Yh��;�  z-iu+�"A�!�d�DE�2����2��� ���!�!�V>9�p�%���#7�Daʯ@�!�$�5T�7�(4���D�R'9�!�D��s���bN) , ��'��/N!�d�	y[l���C��!�u�ݜ(N!�$Q� ����iB7��P��Ro�!�HP���#f⎧B�@l%"��>�!�حTD��A�BW�v�j�!Ԍh!�d͸J�����n�5f�ؑFՉ!��\�H�=�API�*}q�7�!�D(^��p���H�n�s#�7-�!�$�sJ�|C�O�g>�ջ��-�!��W(%�䐰��d���p�䞅#�!�A�9Tr��	t����Aط/�!�d0�%�UF�@�-�E�:B�!�$��b���w��6FdH�y��;!�d-�d(�"�Mrx�v��R!�dGw+숳F�ğ#��i ��Gg!�$" �X8���@�I;�!��إa���8���;&��9[썊!�Rj�։(@�(�vkB�Y�Zb!�d�=�� S�K� ��E!K�_�!�0c��K��?��(9�OW)b�!�!Sj�X��)Hn8�X��J�Do!�M/Z%v���� vb�}�����!���^��x3��.D���Z�8�!�S6H��)�6�Ċ_�2)���[A�!��@T�ؑd�� �B�a�ˍ
�!�d�1�x�lK�o���b����!�DT�4�l����@�}E�5�(��!�$����i�B�,B�A�fə�;�!�$B9�ڲ��Yz%���7�!�$� ]`-1�LX�\]�2�~!�d������ҵ3Er���΋|!�d�	;8<�P�Z517�D����V�!��>'*Ly��זsy�S��5)!�Ē�kfj�A5H��)~�(�Bb���!�� ��w�G/;��ĺ"�F���Ȣ1"O��%�	�,��x��@�t˦"O�H���Hw��hĮԥ8j�D�%"O((�U�˻-o\��4�K�W��R"O�����ˍ�dq��nΓR�ڌ��"O6�+7���r4� ),�@��0"O�,: �C"K�D4���϶Yh�"O8�%��.0��%�pk��Y&*PZ�"O��RV��(aLH�
�9�p���"O���LE +)��[ĩ�hԈ���"O4ĠW�  �   =   Ĵ���	��Zx+tI�:.���dC}"�ײK*<ac�ʄ��iZ�Fm��x",�9
�h7�� 0�<٩&lV�c� Y�N�HhƼ*S돖h�n�:�ܦ�Q�)L��u�'˷e�n�]�O�pX���?��ԲBDn�1��L	dp �(�T!�g�<�-TCH��I��>9�)�1��E�j��/ZD�"�Qzz]2�
�8E�d�FM�lJ��p�,������!�v˓4&���k��-�`B�i�3#��]`aEH�
���J<Au�ޟ=\iO|�h�*��0B�LK�)�n���Hp-.8�7F٣��	�T^��H_2T/�I���؉C�_>e��.��q&�(VEڅQ_�e��G�%/����
k��*�Eþ3K�D;�D��/4��sh<R�&_�Q�ֵq"J�#I6���H�+��hM�ۓ&>mЌ�L�T��G_ZȬ��F���eoɏ �p
����n�J�<a�bTY��SҀc���'d?��D�
�7�vȄ�WI ��ɶ�`�+O4<���z�хK/���g�4͠dǌ	2,Ʊ�sΜ)������Ew��<>c�CC:(��(�'dм������'=��)�j� L9ީ����;��4xz�$ �T0�O��i��������>�O#ג�����PՐA��N�MfT0��}�'m�D�J�����|"�R�D��sQD�$0<e-E9}����S�_d�	;8��e5���3Y�r�SQ0O.� �N� ��5�WaT$1��	�q^���&��)-���OHdx`��'��'�(�ha�&,	u ]�2��3�(ȟ� 6�`����{��u P!YU?IA1OZ�Pщ\�����[9��퓥b>�1��+w�V����;G�E0r�BC��z���� "6��4�rހa�'�: ��*x��ِD
��Y.O|h�a)=M(�'�Ak1)�9�ēGq�����܌/f�I
&��p&�h0�Y�gAj�%��I@HM�OS�c��x�(H�e��T�3��F$��9u���nJ���KV�x  @�?�u����� 2�1�A"O8M�`@�OB�;���]���"O,�KwK�!�(��F�ӓb[�x�"ONDg�%
�dM��B����C"O�8��%�~����ajih�"OQj��V�X�Z1��b�zgp ��"OR��hً��Jb�� L
�"O��	*^�v����7�6	��"OH�s��0T��ۆ#IX   �  �  �!  ',  w6  sA  �L  �S  Z  b`  �f  �l  @s  �y  �  !�  d�  ��  �  �  ��   `� u�	����Zv)C�'ll\�0"Kz+�D��|���b�f ��yr�N��yB`�X+֜��$��y�"T"!��Fc"�(D��vk��I�iFQi�x�T&5D/뎇qC���bF<��	Nx��Qc�:�(����i� �sf�%��]�!Ў$"���>�୻��X;�'�?	Q F�h�*e����7=K��g���>���paX�	vB��V%���וr�7-� ��d�O��D�Od�Ğ�T�
�H$��)�V�[�cH�m.���O<�l�M3(O0�Đ�&�I�O�DǙr��	S"�Y.1��+I^�$a����O��nZCyR���H��u�dӿSI��Sn\�1����q�B�Y�z1���Y�����<��OZI�'f:ʓ
<�a�#I'_��p�U�hE�a��n�����r� &����6x��H�Z�}��(xz&�I'�U7e�
�Ó(���d�O2�$�O���I覥���T�O�>��PQ���Qȵ�"�U�/n���mZ��M`P�t��4g_���i�����,#�;'
�>�(�"v/P;g�pY ��;�$�Ι��jr��ݳ��t��0���9����*�G���r�S�l]PE�SJ@�ZC�lP��~�hnZ	�MK����T�LͲ�����l�8P�3,r�bP��J��MC��r~��FnQn�pT	BC�L�Jq��G]>P�F�vӲ�l��6����@�o#XE{PZ2L�@=H���-h� �BU�M���i�V6�Q�| �}��*��reb�
tN�J$ �U��ا�X�	�}`�HL(@��Ս y�`n��MS4�i�b��F� :�2%('�C�G�B�	�kJ� ���"�5A3�����k��6��!!~1Hq�Z�a$�Y �3Dp��;�	 �8�*�T&�ZB���c���In���?���?1��i���
[�E�'�`u�EPAD�Z�8�d�<����?���`G"��'��hB��1Ҩ�*Wn���E��q^ڼ���F��Hɰ��$wA���tC@`�'aΠ���V���s��,^$vp	��X�2���CPOB�np��K��;fVщ�)�b�'�&(�*Ob��'v"1#��H2
x��I�*!�����?i���䓦?�������O�����(�21�0�̠xƈ��O����<u���q�C(�d���4�>D�I0���z�Mص
���k[m�J��<93DĥjT���'N�R杩�X� �NYY���M�@���O�<�v�-���p����<	q�hn8x��?1�t��Q�,yj&�P�pQ�ѻ�HA~�;R�|x�V��1��M�`��<_�Z�;���Ӗy�� Q��� P�}J5K�P_��SB�$���M����|��I�8�Y~zX�]���O����O����OB"|RP��&3:����W��{AN[G�'2�o���mZ�<�ٴ�����/v1�m+QIB�FC�� X���'���OEt�����I��x�'�`��4ʔ� UN(X���x"LI{b\5|Ɣ�a@��Q�㙴C��?e���zL�J�')����*]r����K&��ā��Zʘp��ᜭM"�(�L��OOl�Yk�E?�0�G�r~x`卓^��r�`T�MK�Z�����O��	,&������!|���-	�׶i��`C��lF{����!{暑I���o�)Q��R�Tp��d�O��o�M�L>ͧ�(Oʵ�q��1'n>��uk�v�����[0e�r�'*��'��D��8� ��W�o��1��k�m��Q��	�Gm���I�$��-��i���b ڝ0 �Qka��)�؀�t+��46�a8 bP�,�D{""�� 
�����տ�0��F@^�6@Naj�gI��L)ғ��'Ҭ�	�e[ �H]�v͟�Wg��r���F{��	�F��3�P�^~8	1��R4_2�t�r����]i�4��i�c��8nZ՟P�	�����@7�n�����X|�	JyB�'I:��q��&k�����i��1���8β�1��ل/��pQ�O	�Q���𪅅tWQ�lAD�����x(�Hͱb��-�s,��W���y5,����1�A�K� 2��c�2�J��D�	�c�����Ŧu�4�?I4��-��8��M�&)l+DH�/��DiӶ��	y�韶�>Ѫ���p��%	<�D�>�	f�I��O�>7힡N�ֵI��H��v!�;g��n�ݟ�I۴9h�ِg�S�~�$0/OB��������9g..�v��WŌű�١����؟�Ч*0:��� gBn��eL�`�q��  1.��k���  �l��q@Pj5?��'(�*�ⱥ��6L�I�dI{D�RKR6�s��-�
2&	�Bʥ=��RV#8?i'L���|zݴ!�OA1���i剜L��{�M�6\i�IY��|��'[�'���'~�$�dԚ3 [�!Xİe�� ��� ���۟�nZ͟��ش�?I4-"
��H�Ϙ��1�f�қ��'.R�'����F��'I��'�.L�0,��/J�v/�əQ-��H���u,��\�|��dہ/��9�_>������0K�@[#�>E����Gю�qb)r�l����.²m�K�v̧�j�'�vaA��Ļo��p{�˓�	�t����i���'�8�#�����?!���?�Ï,,&ؘzs"�;��]�B�����0>� R�h�@_�Qm6I�� FWy2h`��nZw���?q�ey�
��I��⤫�(�l��f+M!Rx�=�fop�n���O��$�<�|�S�ժLb.���(Q�~+�d2�Pb��bp���y�R����G���e����3<�Fy��<N�ą�I�]`R�Hgc�a]�(�윹/Ct�%�@P�7mƙ-��9
t�z�
�O�5
dÛ>U��kF�#)vĤ�폩���'2� §S4h��B�'�J�y����s����	[̓{fb YBj�?I�8d�����~�nL$��Aش�?Q*Ot}�EeM¦9�O@���iP�3�>(�2+�(0.�B���$�O��$e>9S� �9*lT����|Ă��Q�&� �Q'�-�\�@�)�&B��{w"�
)𠡉���,��	F�0&q����Ԧ���K�9�>�v)&"'�e����U�p�����\���'����m�O.�oZ����It���g�(lL�Z5�=d��'u��`�����-5v��᎗�BO����
��'�ў��ϦI3����t��\�������c-��M.O�	ʓd�ߦ�	ڟP�O� 4*��'Z�P���S� (�FEO�v�2l���'��lH*P;,�j&��. Z蛒.�i������T���PGЂ�~qD���O�I44]:M�j�?m@D���k(��:�C�!�T��gG��n`r cN~�
�?���h�Z�ɠ`�̔�֪],AȬuS�8u-*B�ɔ^�V��D��U�0��v�g��#<�O�Dz�
P3t��G��95Tp)Ԋ^2v�7M�O��3l�����?q���?�+O��u��1��l���D0f���@�<����J��
mj8�F��% ��$ bjڷ$,X�3@��Z��C����;��5+��q̧�b��'h�� ���>�9���P1��ڲ�i��ʓ$[l����?e��� "&�"�N;8�|��H�J�NY���?�+O^��2�Sg~�g�,_r�Z���-1�Zl�$��.��DŦ	�ܴ�?�еi=���?-�O@���)�^�X�b�G��?u$8�Gx��6��O����O�ʓ��n>����2�\ ��K��8!�ׇl�B�I�<��� l�>?�,�D�Av��h����7��ebP&ŉ|u�I����zK�">�І�9N/f�3ɕXLN�H�K&jEf��I��M����C�'r��2b�<��z�X���x�0zM� zP"ΥX� �&��*��'���'i�b˓Fή@�,O$���q�BŸ�b(9��X�`����O�ݘ���O��D�O�}����(9�W�:@�d�c7C�؀���>HW�b�$�Ɨ/nQ�H��a� 5��șp�ڊP2�|���B.2�1�@�`<�Z�oeK���$���HO��A�'�B7�����I%����) �w.�=`b�[�b��e�' ޙ���'B�~2��(^1l�9�T�\�0�
�s¦ї��'�ўʧ2��+�Up2�i�	0%Jh��,g@7m�O�LmZ���JJꦩ��[y��OL���'o��@��ܤr�ŲA��7��-���'yr+6,S�'xb�	��E28��#�GF�sB�۵v����PtBȿQ�䍩�o�;�h�����J�d�C�&G�H�:�3В�܈�.�OxnZ��H�h擧aH�Г4N��;�T���V�O��d�O@�)�]��A14G�<~�beΉ�F�
xD�s�$HoZR�'l���U�_�W3�(pOթV����޴�?9��?�ē�j��2��?Q���?ɟw{j���L�>�HAǒG-�\���_o�&i�¡�/B��$b�%��O'�}A��~?��ǔ�]1����а(���.i5���R�Cr�S���"s���24������̭�=�i"��J'i�yƫN'F����/y�4�d�Op�����O����<9���?A��v� �_y|����Eay�t�'w�U�W�)	,č�#��,��e���?i7鉄�M�������$������+����͉� �<�0q�X}�'.�X���OO�i�i��k�&�W��9� B�v�8Y����L�R	��r�u�4*�8�"Dj��
? �0b�R�m[��H�	�t�� ������<,F�9�J'�����,ʓs�P�g��攠v����
�@�l���0ٴg���TGx�#W�,���u�Q�%l�ۀ����4����'"���g��!1}��P���$9�<��N>���ic�7�<��C�7I��'�bF�R�"}{�������U��	���'�Hh��'hR�'�����L2�j�w`lӈ�<(S�����S�*�ҩ"��J0x�|��d5T���8�陽t3D���@��1�\�V�TE��ߦnRX !"�H,���ѱad��ӤIlZ�D�0�����-����s���(�`yb�'��O��N~Bd ��h��)^<���J���'�ў�'S���� ���h�O�<+�zƥ�,m�6-�<Y�H[�,�4Y���D埊��'�: aa�9�&��֠�P֖�p��'�RKJ�QaࡥO,��6���F���x����U�t��-#�b��'tĈʃo�3l `���P�*�p�d䁭=��O���س�7}�`�K��V���O
�ZG�'G� $D��5��!�XZr,$�r�_t�p)��|��'���'6?�ȅڜ>6�P�c�Q�[$�-j�o"��h�fb�4c>�(���	���8��g�bD��`�i "U�(�1l��?���ԟ��vy�" �!"&�J:�~�Y!�J]�����8j�Hq����vBF� ����w�t�{% S/YI�dh��ݸMp�:G�Ġ`frc>I3d�*?��Zs�����̚~� ��$��M�[���O��	-&�ġ ���
�d�	 [�)0�Ԑ�g�r�'�a���^6Gª�+���z�q����^Ѧ1�ݴ���|"�'��$
"3z�P�N�3ZXD 
M�>0�`�g�#{�����Oz���Ob魻�?������h�l֒�����"ǚ8� ��xfh�I��^d��*��e�L�ҡ�> �N<Dy���� ڝ�"�;bi���tE�
q)T���e�9
�bW'�]n���I�{.%�� 3An%�R��ŘT��b!�Tp�Us�cJf�N��G�i(��$!����іK�$H��KT�ʈmn0	�ȓZ@�-Ȅ�T�>a����f�'��!ݴ�?�-OlY�iy��'>,�I��I.>
�P���_9}JQ���'�bi�8G��'��5�虊�S1^n�ᨢk>�\�Re%[*7�ia@ƚ3R����mٵe"`��\*:x0�`� �;q�n����U/_T(u┯0S��m2�L]HL�x�r+޼~�x�B��;��$��b��O�n����/���$�&�	"q��0��'�a|���28�*D暵omJ�ٳ����?qR�'Qh�0�ğxCl�[F��2� �`�����z]����OJ��|�6Ok!��	v��xĪ��:7X8��@�,=Ω����?)g�(m���嘈+(q	��ُ	R��R&���I[�vt:Qq劄�H�%a�K3f�ɘrwX�+�ʇ�v���JBH�>*۰!��&��ȭ����$
�
"Hu��!o8ƈ������O`�%�"|�V�� c�R�{VJHA$����j�<��3:X ��N�j�2�i��h�'�Ɍ�HO�����Ee��ϊ>.���D�٦����P��xx��(#���P��͟���ἓ�OZv�N�{w�Y���2�ij�(���P-E��8��I,P����|G�E�d�&�ɐ\���3ʚ.k���J��Z��Ȅ΂�}�5HG'4͖��D,�>�~9���Oq��-ȡ[S�q�&��hfh�� q��'Z�@;��bΟ�'���[�D��`k����ų�^��"Ou�� �0H���D��.�=�`&�>��i>���Qy�^�Sj=S�Ԓ���:0�Icp��$1�'R�'C��ȟ��	�|���
(��p3��e(�DQ���'MlLI�BM�, 0Re8EDʀgd��'������<yC�6E������1�
�6�g��B@d�h~|={ �_�P��Q�0+�<1��^�p�� �x�����2BŬ1����M�"�	S�'���*Ŋϡ_�BY�1��`b�@	ӓ��'�Z�h�l�9D�`xA�,۶f�&�3I>�Q�i�BW���BΟ�Iğ�(t@]�)иئ$܏��2��\ڟd���W���I�$�'
n��IM̓�`4��$�B�� �lp��	��D"<�קɉ3�D*7�%�V �Qi�Z���g��O8�$�Ts�I�K�0eI���x���#�B(D�D�e��V��!���i�]҆n$��]����,��s!:Y�x3��&�H�&�1�h���M3��?Q-�����O�|p��Z�PO)���W�m�p��"�Oj��S���+�|�O���6I��.p��z�+ߎ��1Iv��<�6`;�S�O�r��bo_#1�Q��O��`�Ol�K��'f�O>]s!�)6�����7� u�6O$D�L��Կul�h��)[e�t1r 8���D@�'��Z4d�b�ĺ�	�s�.q� iӄ�O ၄�����O��$�<B�g؀�QES�-Ψ��� r��X�ʕ}��u���F��X��ԙ|RLk�<0�ģ�0�P�c'�Ȃ=�āɕ�bS��hI�A^P�����|� ��FY 4&�<"��ik���?��O.����'���'��O:a�*�u�c'�[�p8�*�&!D���q��]T;�%VZ"�q�7M�<���i>���yyR��#�l��c��7�F8qQ�3l���{�aX<���'���'�n����	�|1i�1!�`�U�R�a��}�P)ӽq���Z��n��z�.Y�8��2�E3!��<)��ƄnU�p��́	P�N�2U���E����La)ʙy��݇n;��<��cJ�<�8��E�O�W`������S*�����?�&B��x "�E<a�t��S���?qƊ8b��@�fE�=�p��cʙN���M#K>6�ŀ����'2j�'��U��/S�mr(C�C�|MB�'@�}���'7�2�L��B�'1O��)d�e
l�2j��~����'��b����{7p�ҁ�Q�ze^ػ����ax��?iǓ|��&)��[��۾!�6]bs��&�y��I2/�ȱv�ۇmA0x�w�ߣ��'@ў�'T�� $V �*��1M�!9�n��������ǾieB�'��ӖL9l����U�M��C:Ş�r�I���֕����ˣj���<���I�@�XP��/�0w��e3��}O�DDx��)ӁWI^ �D@[���yS	["��I�b���r�)�'��-��j�o��Bch�!TbL�<��H~�\��h�Q"�=�¥v�'V���HO��#��D�:eHT'nA7=����������ğ$�	�x X]Y�#U˟���ڟ ����;���s� A�6�ͼ�`���_�\x.���I�'���pΗ�h�ę�@���>j�c���� )LO� R)j�F��$�`�(Tl��X�hsC7�������$݂)V��Q�j�'� �`��O7	�!򤁋m#`l���L���r�J�s��I�HO�I6��׶j,����D�) �LyF�n��b�I�H���Oh��O൭;�?����do�JBq�O߳>0�pe�	>'��X3���p��m�p�xY~0z���Q
�Q�h��:�0�Ad��"Q�Yi�E�H����s�m�Q��N�'k�e˩i��̃�i����#G��?�r�'�cbC����t�/>n<��'1��{ LEW��d��7,ȁkN>��in�'ΰ�)��w�����O��*��H�f�eȈ�l6�!h���O��2}����O���/��!�$j�|p�	���w�¹B�͓�
�xA��b`H@��2s��ғ�	�
�
�BKrB��)C�+F�8EP6�ݑm���! E2�d�֡Rb6����I
X|���K�	�V� ,]0� H�q�޳tB�	�#!��RiW>�N@��4���������!��\�x���v�B�cF*���.w�~m֟���E�ԁF1Y"�B�@��X��i@0v����U�ҙJ���'�����'t1O�3}	�nK�W>��ոc�}����5Fx���]�m�<�	$cH' ��A�U-0Y�	�L@ ���o�)�'2 ��j�9DW^�b⏊)f�ȓw�@�BlK�]����A�+�LG�4�'s��0�Y����sX+lh��4�?����?Q3 Y<@RX����?)��?!�w`�|�r�����d��#O�/���4��>k��{¬w��z��;ݘO~,D�!l�`?�C�	�sZ&���O�%B4Iye���VDZ�e�+K��4@3�cl��|j��Wy��	�_�j��b�~H䈨6c��A�,$���6��O<c>c��`��5���0� ё-p5B �0D�l����G��k�ˊ�nsfMquA�Ob���D���t�|r���E��Rgi��hT:�3�#�+�:��`�6���O����<�|*�EѪL���b���t��9���"���r���a�H�h�h�
 Ax̓���.f�v���a��� SD�
A�j4��8(�)��.�����FX�'AB��!�!e6X�q b�-zf-�Pl�?R�i�f"=1���F�r,I�G^������ڮ,�!�\4Y����gᑄ#u�UKw�E�<��'� ���D�j
%?�k�IӦ�X���΄i�YG��O˓�?=Ҩ���&ow�Q2���:Z<rw)1F��m�!�����rv%
�Qι�J(��O��C4�T�8#�����jX`)�͎�]H�L�w���*�?fPɟ CڴG��I�+��YI�AG,�Bd���
`˲�OZ��C�F&(�E�<j��Q�m+<��2��O��"(�l�j�$��G܆iB@�'��I9Q<M�O��`���'��pR�O	�l�lka�l�ҽp��'���-"B�����Uh �{�n% |�?-x�m�k�\蛥��OiRyb��"?��mL/��Ǫ]�9{ve�"����O{*��k��|��� �L4�X�O2�z��'N6��#}:�O6d��@*
E.n�P����:>pq��'���-Řn���jq�ɶ/�����d�H�Or4
�� S��臃C#}�|q�uU��']��0�O���'��T��R�4����O�Jy��Y�
hx@)���p�e�����)�|�N>���V�|�d�Ȗz�'��iP�	Y�͗~�zlq��J?N ���|J>IG��3=	(AX��Է}-x�����M;�V��s���O���8&�<���F�c)�+����4��`4�{�<���k7ڈ����T4*|�PIPQy��%�S��T�H��kÊi(���7�����Ke!D$��M���?A�����i�X�8Y�N��S�F�F�a�P�ǉ�:1:ʘ[�����
n�'b�*���g�rUz��[� ��)�Q�O�-Q��U)S4�RA�q�М)џXI�ШF�8e�"���hr8�;�	�:����ҦAk��;:�0x���0 �2DU`D&�Ą�<��"%�o?�	Rh��a$���O��h����ן�g��S��(b�Y�l( �6�+�?�-O|�$�O��� ]z<�#�x-�LO�k�L�a]Oq�d @� �Q�+
8pџЬ<݄�b�ՏW�J���6`$S��N�s%�Ĳ�g�0R�E����>:y���ڦ��.O�p:eiʴp�(!�w�گ/J}Ir�|��'�xa��tF �I I\�C����� )��{��@
�Z�N��1D���?-Oe)t"a}ʟ8˧�?����W��M!�=ڸ��p@���?q�J���0��"9a���$�^���d����*�Fu�1FP�tĈ���`��:����V�,�i�*�>�`�R�����O.��{�Y�)0�0)���XHC�On4a�'�6HO�O��� �L	4`�4v�"���0p����"ORY�v$�I�>��A���<�&��g�	.�h��@R��*
��Z��K�/."���ˠ>�.O���!����$�O��D�<a�J"装CSx�(�&�[�1V`x���'cQ��GB�8TX�`����|���H�����ͧ@~�s��]������&�4��f�#;3� ���T�|+�O���S�@½�2	I$$��f��<9"�]ߟ ��d�L>���ʟ)��\�7i�x >h�#Ύ�y(��a���u+�~�
�鳩���dR���	�<Q���i�&��� s���J�-!���ƽi/r�'�T�b>i!���tլ�B�o�Tz�4y%�f�t�27�^����c6�����ز�|87DĮK�����݄}p^Աp�
�a,�l��nN
(
�g(�(�!0��(��,01ʑ'����צ�ԟ`ڴG5��Fx�+�V<CV�ޱ0�����`�9�y�B�;W���8,qV����� ��Ey�a^,6�8�4��dA��H?�p�J��M�'6�䅱=>YkSB�������)Qtd�r�%O:`��I0+ 2Yj�ռE���	�,I$FI��$R�l��.��T�(����%�Jse��4�!�d�1!P�4`��2��b5!X7�����O�����^/{Lf	�G�h�bT�|��F�T��c��>Y�N=]�p�ꡄøOl�` ��9?)eE혔�C,�*WI���l>�' "H��f�����S�������'f���@� c���J�!(E�D�̨2:�x7�!1Pv�3+�����;BF�tӖ�F��4�b���*�'8��!BĄ�pb�"O`��2e ��{�̙"��Z��ɇ�h���K���9'_�)QDl �XX�b}�`�D�<1������I�)�0y���d&v�Pu���,`�b��)�G-LO�Bg�Y�C� pb3(������R��\�>�az��LP�1i�,S�i��%[�`�s/�'��%k����Ϙ'��b��3|,��ႊnO���	�'����UÊF��	Sc��c(2:,O��Fz�����
� ��	�p��s"Y�� \�~c`X�Q�W�A�j���˰�.��B���h��-�*"�ݬCX܀K���U�b�T�J���D[�Jh�$�O��$�8t,f9��B���u���nXK�Õ�H�t% GkA�q�D��¼���e�?�(O6D�7͌"Jd�[u��v������s��Z�@@�Y��YR��ѡxy=S���(O�|+��'��7m�c���M#���Z���,'��P_�t��� Hɹ�F��&������W���$oyb��u0����O�{O
��Wb���
$��9m���p��k�4�A6y�r�'����� U)H�h�(aoޜ<�����'�)#�k[�Z�4�$1�,�q��Lf����e�}̧�LMҧ��N�(����:y��M�UE�t����h��y�M]'����D�0z���>1���-h��PyՊ�+/U��h�a�Ěvi�Ox�nڢ����?�*�+����W&^�XN�y��j?D�������ti24�ȷ���r�=ړ	ʑ?��n^EbRc�Y=�%��ߟ��I� ���X	58���ǟ��	ԟd�Xw~B�Ζd��)�`��9(_���o��{6�H׬�6���+"���
��K���� "6,@	N�(p%KA*q�B�.-^�����C�a��0C�&�4����u�Ix��j8a�&-1}�Ɇ8
�V��P�Q4 �L%��-��剘F�������Y��䓢yb@���,����]�F �1�ѡ�y��+Zڰ��c �V�@��Wl@$�?YR�i>���y�'�\���Ʌ�ߣl��9*p�Şż��5��^��'�R�'��]d���|r D��q
2�q�ʔ�N}�vC��V�Z0K�(���@�P�[]iA�H�01��<�1��#�q��g]oC@��*	s2@	án�
\Zq�� ��I�%��(���<�b�Z��ysh�>[R�@Y'���H����G���M�E�h�'X�쩷G��J�4!e�"�R�'�RA��&\R'��A�f��5I/O�`oZ�'Ǝd���~��S����T�� �<H�N��������c��ȟ�����("K3(�51D�#~�A�R�/:��Ev��9X$���A�{n��S�$]*T�2�<�w�]3W���)	�M�z6�ӷf�����,W,W��A�
�UL�cU,ѿH���<�D��`P�4$��O��U���R��G��T=��;/O���Ŝ�4$�&mݬ �`ѲgF*
m�}B��<@g��7���(1c�=h�h���n�dy�E�!��7��O��$�|I,�?��=���7GҿN�y���]���X��p#�-���/Y	�=�r�|��d�d���t������D3/n���b�a-0��W]��y�#�T�i��
@9�:�^.8d*�j�L�'8�}zs�W*N �j��U;���4�~��I��M�P�����g�? �}���%�:�jVD�%�Ԙ�@"OX�򇁼����D�����w�	��ȟ�l�m��>L�4�A�*%�:���O�ʓd����i��'?�]��B���A�M4k��)b�K��AA�i�Q�4��6m!��y�u�3
�K֧2-��'���*�5�+6GK̍�����8�e���s�@X
��X	���K��=�O��Bq�@��&@�%�9.m�)��Rnyr�S�?���i��3�y�Q^&�4@!N�WU>�@�G�}�!�ѬO*��ğOr8��匾.�K-��|r������\<�0s�.F�D~�R�JE� �v�3�)�x���O��d�O�0�;�?I����T�)��<󂀒�]�^h`-K¦�x��P�1nhQr�j�_�&� w��mS�}Gy2��*��
�-$F�F���l. �p��M<$�*��dU�F�B5SS�DdI|B�+��|��O����'���	�VA"a9R �x�"��6�nӶ�Fz��7����6f��>6ҕ�Ao�n� C�$o�%Hq�_�:��ct��h�˓ ��6�'|�ɭ��1�I�L���|z��Ҧm�@1:e.B�x@@`Rc����xՏ�៬�	��X@FjߐW��fl��M5�tjA��p��ܔdX�)@�j��A}x�RT�[%+�8���ٔe<��A6���h�1�K=|�I����Y�O������QX ��B���<Y`�ܟ<���$��4[>���(�X~B � �yR�*m�8T� D�&�|��rDO����!�S�
�<	��"hlr`c cE<)���f�Vy��'2�';��a��?��&�>d�Yi3)_ld})1�>��'��[�أ�Oq��u��;�8��I&[���@��SA�'�a�If��'J� �z�h�aF��j����,c�&6��O(� rp�Лu��O8�$���e�\� O�C��0z�	�<e6ps`�6�Z%lП����埼Γ �<����}�͟k���_40Ċύ�^��sgű6����?�o	+�yR��H���ON���O��Ɏ<�n ق`]9Q���I&��M���	�O����f�n�����钀�?7��:��'@�`�lȍ?�5�!ǅS=�X�P�'Έ�����?Iգ�&
��ٟ��	�?a��e�\q���AL*�:�ÃyR�j��O�����h8�H�`�CE(=���-�u'�[/v$$�9A 3 ڼ)`��3�M˝'-� ��?	�
_�_�b����$�O��I;h�rL 5�[-Cq�	�G�b[b����g��j��OL���������y��#a��i=$d�Pc�6� 
4
�X$��1�R�:21O$����'�R�ɑ����O|��<ޔ��Ǫ.��cS���7�l�lZ�
�Jg��C������4����y���[j�T��@-�܊E�O	�N��0�ÂQa�F	EP�j6���Ho.�2۴\%��^?��S d&��.�n���a��1�nm8
�'LF���h�!հ����\)4ܛٴ�?���?����Ol���O��D̗7SDL���t��Ű���]�n�l�͟�������IO��'u}��at�]�n� 9�E�S�e�nZ���'���'��S����O�T�pi�\�¸1�KvO�nZٟ���R�	P��~j�����r��2��yČ��HO����$�6a�%��Vb��rN�؛�W� &��g�şdA�.��LF�B���:*�8Q�A-�;����OH��6�i>�O��CN�R�$|��BO�|���K�"Om�G�gBt�'���.`�"O@�f���f'V��p%Ѻf(TIF"Or�B"�Џ.�z-Q�NُL����0"O�qZS�k{�XBn]��ȵ��"O�e	&�P���th�+��4�x���X\���A� :#l�%`S�0���ՈZ��^� CHÄ]s��8$�P� ���k��4���uozYj��_�X/��i➈ոb� �BB�,yڝ��ɘ%y�|�`c�q44+R&�P@2�a�ኝL�j�ؓ��gݜy�æ|��)�(��7���K���Q 燇x��I��[�l��@��S��Up�?}p@���طg�n��L�R�+�;4��a%�ZѲ�ȕ�4NRY����i�v�J����^���L e�2HD�(x�4ѵ�R�
�.�$�O^͛�&Fk���	�=R�R���s�dY?A	K�]����0��	'�P5s6�>�އ*!:k��5�Q��N_�d}��>1����	&�4�iCBJ%��Y�2�dD�J;2�'y�>�nگ^$�1*Ę�+�H���I��R����'�\�ɀ��~�U`Ȧ���,���p<Q��I�:��p���,'�H�JVyRz���?q���?��N�yuR�����?	���?���Ko4�ӆL�!|X��a��J�c��˗@Ǯ_������iI6� �?P�1���
�I���W7��p�(°i�8|����m���Џ�a���nZ�']ތ�d�������N�� !�jҔM�$$sB'�^���t�'���9�X�4�P#=i�|0A&�6�B�D �1�p�h�"Oxe���D�>N*���"J�9�6q�ė>IP�i>1�	A}B�)]�RDɷ)Z 2XHFÐ�?����(�Q����O@�D�OJA�;�?����tJ��@J�ha�X�*���j�f(��pg���!�8���k�s�r�bE�I��� *d���I8W$����c[�D�vdy��-��8BF`�S�3w�	���O>�ZdF[�fLY�
�	c����X�Eg��'ub�,�S�*UQ�#E9S~]��/�dB��+~ 
G��V�vi�"�?Zb➬�ݴ�?9/O��nW��iXT�҄P;�f`qV X*jdyH���O(��PI��D�O��S� ������3,��)��'���DnB1:����@�6�&zg��~�ΰ���	?:�����[/�̡dIuaB�x�\�X�!Җ"���'jjUH��$HKBwQ�89t�O.�o��~�H�Y`XL����yWO
��'�a{2�
� �b����P��$Ͽ�Px��ff�сc׳��6��f7�����O��\�$i��io�'��S1���mړ,4(�r�ٳD1,�p�
,U.<���?�F}U����cϓ�MSsF\)]��mZ��z�'���h!��	��,@A�_Z$��8s�%�¬�E��)->s��1FF�#1M�6U�E�!�<��k���{�H�"�_�ē�X���M[������j ?$]���P�	�>�G_����P��l��a�^�$蓉ï��<(6(��\�^9�5�i>}ߴ&q���x�b�?&��٣$��(��zd�@gp��o�����Iҟ(�1NŤ@���	Ɵ����<��#`����$\�8ՄхG�4:3��3q�>��t�k,f��t��1����7�λ�?)��V[�H�i�/�&NV�$��b���nZ�f�le���&PX�Z����E��]�+d��Ɍ�a���4l�6u�|�k����m��O7B�Ę����c�"���r˙B�!���X3�fG��x��JȾ,>���Oz8Dz�O@^���p���;U6��`��.zU�hǞ#�t�[�!�?���?�������?1�O��8�(Ҙ�.�ȱL_'=�5�g�]� ����.�,ѣлi0�6Ǚ�CQ�؂��͑-�v�i��.�>�S��"8���2���fF�E��(��Rd�5�����\�UM�)a�o7�n</�&�1 ��O��D?ړ��'�h�:�)��F�.�7���;�t�
�'$h=c��ޡd2!X'��7 %#�{�z�
���<9��ЦPԛ��'����^�P�Dh�6c�?xA�5-S�H���D�O��YU��O(���OFpy�eǔ})�݁6/|�l7�Z�hl���*V"~��䉄�ԽA�ay��4x܂�P���M��J $�	3���*1
��B�s��ۂym�8Q�+��(ʾ�Ey����?Q\��9�v)*5��k�\xA�6T^	���?������O ~Mڑ�/ �\���'ӫdW^t� 1�O��1�Πq���S��\?pL���t��oOyb�TP��6��O��Ĵ|2��%�MrM6G��W#H����{��!�r�'%"(k��7��!! �&u�H4��2,�l]
�_?)@�X�h�r+�:Q/̕�U',��9Oˀ *BmB&v���CƛG6��[d�H����ז�.�P͟?�B��N6�'������6�&�'�ug�˪d]���	��*<Dx"У�y���� �1d��'L�9���8�p<����+���(3�Q�"�@p� R΢<��?)���?�-�+U�f٠���?A���?�S(w�#�ڝZ��EQCf�&jD��(p]9��	Q$�-34���|���C�$[B�D�_d�T;���+'��i�`��"���Fd�%G��[�*\���0�7�S71'�a�w��p)��FV����M/V��ᨄצy�*OLt����T�?O0�rn._/��bY6���"OddXѩ��ܰ���]*p�`�t�>���i>���B}�a�!+!�hk�%�v0�J�批P�[р��+_P�$�O ��O�h���?Y����<��mY�Û%��b�H �pR1K^bX��x�
��`@��'/�:�Ey�I��h� �"��/p��p�3��4}�h
ƩS����+T�@.J4�b !��Z��FyZ]��#���|��) #M~X�y�`�O���ɗ1�P5�e��$s�0X���(-�򄞚-���p��z�(���)�5�qOn�D�ɏn � ��T6-,b&<@�☞G��)P2ɐ�YɲY��ǟ������|���|ڗ�V�NҀ�a1Kb��ZU��:?� h;���K��5�a�����H�8�\\Ȏ��U �qs&��C�@����+jJ�+�P�e*�!jp����� ;R>��*���]�R+��'@�Ɍ|��G�<���Bmԁ6�v�0��ZX�`R��	E��4��oN�i�,1��+(�Ը�B4+2�u�vII*`D<3 ɜ�d' @��Ay"lW�e��O$�^>�1ԇB��D�C�a&�adl�	:��إ�!�?�N�xH�)��j,j0[W@�fA���� ��n�TK͚}0�p!q@
&/��Ӗ����8#��@D+���=Pp)��M�B��j�'Y�u��+J%? x��,�X\�'�����O��d&�'�M�� ګp�v��J�O�Np�bɟy�<�����@~�\����Q\�!f��t8�2��$��.��5!H�h?`��
��4�?9��?� &CG�M����?����?�'S�t����3�F@Z�l�j���BƩŶ ��i��,I�N��� V+��ӘO�Y���矌�*�l5��k�/�%Z����ِ̲�a�E ���v�,@�5�}��f�?��� �X맏�(Hb��
�	_}��DJ���\y��)�3�$D��t�J�[�8�H�,*4�!�ʡ ��Z�Ȑ�<�ѣ1kV�*��f����S}�I�q>Q�PlψP�fU8WN��U3�`O�!�@�`��?��?�@��@���O��S4��B��.��k%�|'�If�7bN���Ν�Qpb<[4%�J�'�N��«�X�̽hV,�,"��ZP��"���v��Q�>I�P	�45iџ\���+ ,�g)�Md �[���q]���O��0�IF�@��T��4�\U��BDZ`��#��ē' ނ9*� � )��Y���=i�i�Y���c ؟8�����ӊˋV`Ŋ� F[ P찷�_��?���v|�t���?)�OV�uKħ@�iF��m� �z<��C�2u/���a�<��:3�ߞS�6��(O�Q�C+]���' U�Zz��FI]���!�L�4��ģLR�N�l��Q������O��O0v��K��[��а�e�
�y�(S$"�H�[A��f�JhJ�B��Pxb�<XDIFK�!s0��aW(_l�u�s�4�G����4�E
A��|��N<e��(���'	ў��uN��nJ�� ��9�X@p�-D��[�K5y�z1f!�y�T0��.D��!�̻`��|ف*���¸ F�,D�H:�f�6?Ӫ�r��*פ�2PF,D�\���@�w���Qț�Vwr��"�?D����C���BVO�"c bУ��8D�qؑƂ���O���<LSF�8D��(��"�a3M�j#0 �M8D��ɕ)�rЀ�K�4ZI,��7D�|�V�ۅ,��L��P6-���6D��2e��hp�Ț:湻Ta:D��kU`C�$,�2� 9E!�х6D�0�q!J�jp؜�4���Y^%3��!D��xbȿ'��i),�;Re?D�D���J�i%�)*�e#"�0D���P�ϟ1iD�0B�w4m�r�-D��h n�?N���b=]=lU���!D�3�˲4�"�؃�� � ��&>D����Qڮ��Ɓ�56ұ q#7D��H����P���'tұ���5D�����2 b�����W��GB/D�@�cd�M�4�w��@X�20�+D��S0	�n'�U��ap��C��*D��GE͔#�41����PK�`�%D�,��l9$d��Ԍ�yW��p�8D���i�B V�)χ�5}P�U&8D�`SScŇJZz�:v�QD^.� S�5T���&��GŎ�r�� �PE�0"O��jP3zA2�jKxʎ	��"O&Tڢ��s�hA��`B�;_�A[""Ov�5�G1^(Q�R��}j�X�"OF�kv�?��iUg����5"OV�Qƪ���zui@�4n:�2�"O��9%�.ZBx 1h��U;0�W"O��Jΐ�m�4@;ufʎM)T<�7"OtT�'��d#Ѝ �;�E��"O���K�![<yS�#s*��w"OHu8�lխS����b�
�\z�"O����G<^��ez��F���5��"O:��u�ԥ&;�1s�3d����"OZ�:F�̭K@r�H6�[+o�H�!�"Op�
@"�W���H���;sp�8��"On��!��Wf�)�;+Hd�B"O,��l\�m�.��d��{��!W"O��������D�f�F4��"Ov�IG`J�	��ѱ����į�y�$�\�.p �kZ�
��"dCԜ�yr��G�xQ �˸PqL�rG�7�y
� ��5�Pj��]C�S`"OX�q�`� /�:�3@O�u/
x�"OV�8�S�-!� � �ED�9��"O`(fXlR����֘u��)@�"O���C�;[�|!cHJx��H�"O.��F� 8X�P����l�AD"OܛRi df�`D��8�^���"O�:E@�>1�s�AK�tI�C"O��@�j߈,�P)�%^�?����"O��B-Q�'�Lp�5�Ȭ�N���"O�u�$bӟOM <�A��z�x��"OV���%:���")qu���"OH��C回$�XP���Y�$��3"Orx�ҨDrbhX26D�9��	
"O�D��̸$�̄�D�,��xE"O�� BLʠ`;`�i��N�`���[c"O8	9��,L�f�[`lѳ䲜��"Od����lf0J�
צx���H�"Oi��Z7p���1GjZ� ����1"O�I
$S����d���F�Q"Oj����K���Z�b�E^��"O��@���Tm��:4�M�	6�0"O�P�U��/Z�G�տb�p�a7"O���aƝ���s������"O4@��a�D7RE�J��R��"O452E� 6����O7~9���"O
�"f�ĩS�����ȓ��`�w"O"ss$8D�ȩ�Ň��m{���"On�x[��B%"�ĩ=�|�2�"O��抖yLY�����Y��	�c"O�U���K3�B=�ED�w�����"O0��c!T�_��	Y����82"O.1hgL�Hh>Y���,<{ά�%"OVX�f��P�T�9�Ȯ
�|���"O~�#�aT84�08�P��_G0${�"On=薅�,@Fl�e�$<�!&"O,�+���;ND2�I�&�
Xt�"Ol��#��JʂP┠H�6e�s"O�0��;X����Ҡ� A[�b�"O��#D J�:'�t���]E~)�"O8,ɧ�E�*��5z�� �m�b\��"O�u�R��0u���2TnR�s&��"O�E��핅u�f�y�A�$0P�"O���Hֺ_0��q��.�Px�"O����Ç�y#�4�sa
���$��"OZHa�AZ�7ZP���n4J���"O.��Cn��G��`��͑�� 諁"O�M�� Hv�x���,٥��"�"Ox �K�)]W �(�)_�B�<i��"OLEKMNRo��Pԉ݈t��Ӡ"O�������!���STOd݊"O���� ܍a����rI��)Wv�:�"O<�8�KC/\�`|)��[Z?��W"O��+R��h@Mɶi߽44ޠ:�"O��RP��C���ԾjRjU��"O���P⃆Lq4�yq��R8��)�"OdJ#֐Z�1²�)���"O\A[�R#r0j�hcǁ�fp� �"O��A���r������-����"O�����@3\Js��*4�*��"Oz��D%e^؂U�� %��1"OD�)DX�l���4��P��"O
e��ۇ �x(sP��(��Ȳ�"O�1I���@݈S~rYk�"O� �İ4��_�-*��ܓ�9�"Of$����(�J�1��/#�.���"O��Q4(�1"��Z+��k���"O�<�t�^�����Jڢ.�x�*"O�Jc(U.V����`���*�"O �薁��~�	�d��	� � t"O�EQ7㜒ДpRD�̌��"O��1�e$���IW�ݟ!��"Ot�I�C�oP,���@/B:�Y"O2�V�C�O����EZ܁("O���v�è�PJ¯A<'H(�w"O&�0R&�,��8�paMg0���0"O�x�Ϝ�e����@	�Q�����"O����4,U>�9R*	'9�`0
C"O@pkd�J-�f`䈃u�"9�T"OfbѪۏ<�P��T�P�<�z�Z�"O ��ׯ9i�уE`#��X
�"Op��v�O�n�����7����"O�%���:
�S.�0}i2��"O�Ya3�A�������E�Sj�""O����L��6s:y�-έ$@¹�!"O�1B�鋠vq�!�L�L-J���"OvQj0.�,����`P���T
�"OtثB�@�i�D�P�l�$]#�"OL�b�XJf�Z�,I !ݪٚ�"O�-1g�̜V��肅��);B0JC"O.t��"�E��0�k"C.L@�G"O�x��G�j+�P�Ŋ%9�`9"O\) P!��3�-s��\�Q�.�"Oj4QwJ1O����hȦ���"O��ا��<;��RU&B�y��"�"O�D`GG
q�@�+Eǝ��e�&"Oܹ�'Ƥ-����9uqP���"O���&䕇b�ȸ�b��R :t��'Ը�"e��F�㔛
��h��'��4�ce�N��6 ����	�'۲���.͏A��YC	O��|��'!xتD�B�{]: ud��H��x�'����t�J�x5�Q��h��,�
�'Y�]P�↳1E�h`�$[���I��'^$��n�>0U��I8w�L$�'�bx�@�ڠd`�y���^�o�}	�'������;!�<���J��kG��J�'�>dg�&PG~���*�v}�M(�'�
��"�f'hd�gd��d�& j�'	ZTq�g��\fb�8���#��h+
�'�*|�R��9.��h�yX�X�	�'��`����M�ĵPw�� v˦u�'�����
Unn4�� ��ir�5��'b��0���0]��4f� r�j��'=�C��	N�U�5�F�i+�A+	�'�Vu ��8q�ˋ6��I��',���OQ+,�d0BE3'�)�'\�}j�;%�q�a�&�R�:�'��p�ȡ�Ƅ����ʼ�'uj���/�?R��}#�	 S�~���'9�4Хŉ?M����voʈ`~�"�'�ڠ�V��1*p�餪��
(��'B�DA�	:`�$�z��9��	�'w�i1 Ѩ���s��S�$e��'����M�q�4�"������'L�=�i��1�  +��L�F��'K`ěgC˳kE�:��P,8.l�A�'�dp�K�0;��U��閻*t$��� x��A�B�g� �Z&���:8+ "O�u �d[�qi�}��"b���t"ON���;8�:���,�z���"Or��t��.�&��.�jM̔;�"O>�ɰ�׿iA��8$��FV<�kG"OzdX���X���뗅 8�-J'"O �eI�WUJ�c��.U0�"O�<�uM�j9��l܊K%pI�c"OF����،P�,��C�Xx|�]��"O���Vm_!�"�a�.�h4-X�"O�a���[����P͕�2`���""O.S����B`eEL�Pؓ"Oh�ɐ�ޕ���/-���`"OZtW'R�*	t�ⳮ�7�d$j "O2ȹ� UJ�<T�V.G�� ��"O(AD+��r�Rl4N�_��M"O����g�΀�ӪMn�ܫq"OX|�� s��m8�G��P��"O�UJ�9bł˵؈)M�̺T"Or,ڗ"?�ҭ�%����e�C"O�bT恦?1��Ke-�݊eH2�䎖N��$��O����#W:K��'
Py�CA��x4�E����2M�.X�	�'��h����rs�%�ՂV=A�H���'��a���$M�eJ�)Ch��Q
�'������ݳE�X�����ec�\q�'&��t(J�Y��ߡ`�إs�'��	��M���i(d� ')0���'59+&,�$��i'���(岙A�'2z�vmƄ�JB�Y�o߬�#�'LH�C`�r���CǫT�k͎��'q�8*���*��IfbLp.���'+�L(I(��H��H1{�FX��'��`"CG��mY�����.?8���
�'�5q�NW=�ia�b�����'N��gF�C.�(�f���*����'F�4R�@��	,�1�LפTJ��!�'"PE#dA��2��TI���!_2ڽ9�'���`s1��"3�Re�Q�
�'q�I���9I�@��Bb�7�}�
�'*B�+w��6����-f˲Y	
�'
t��-�+L�܅ ��=/����'ޖ�ʥ��q�)"!P�9��:�'9�Q1�eS>J��5��2�z ��'ԜB�I�}'���i�:� �
�'�H�:��ZaDUZ��O�5Մ1��'b0��u�J;]E`Uz��:-���C�'�>� �F[�xr�Y#�-[�����'E�B���9	��H�NKA�g ?D��z�j�0C�"D;t�Ԑ0T���;D�X�W�4*���,��U�Y�Q)9D���مs��ƭ[�Mfу4�$D��"Ƥׄ^���#RW4E7*�` $!D����DA(��P2�d��0���.D�H�o�5*�t�V��9o�<d���'D�|����cV�Y+gJ�=[�\C�k%D�q#Ȁ(i����Ծ��@��>D���v+�x9��ۀ�61��@hu�<D��'(��b�0�Jp�Ƞ$��C�I�vT���!E���K��A��Ą�\]���d��A�,͉�)k��E�ȓ�e0p�N)
�F��0�R\ب��ȓ@�U�P�(.I��l��#�t4�ȓ`�v�� �� 
��%QGAl�̇�8��V	��V�Z%,F�(*�݅�S�? �(e�@e�����G�[��"O��K�*S�r���c�U�{����"O�Y`��.Kn�-���N�
��m �"O�v�Q73��i�6)
H0~�[4"O\e�gD����E���5��e��"O�L3�*Ԇq:2,K�۴&�v���"O8AK��~!�����,�
4�'"O	��Y8Ztv�Ht%���\T@"Oڌ�Ӽb|���X,rܬ �#"OB�:P��Y(�E�$Xg�x��"O0M!����p$`=��*R9}��Y�"O�BЈלR���)Cj�{`�d� "O:�H�b̧VBJ`��ρ?R���"O��'T�K�H��Ug� ��P"O6ĸq�A�|���⎈
t����c"O%0u�^� e�E�R��
H�q#�"Oޭ�i]�]Y��	!�|��:�"O��X�+�)K@�9A�1W"L�b�"O�xa�� Z4�!�g$�=r�(G"O���i����su���5). �"Ol}Ƞ+]'a��ݳ�eD_�.E��*O����GN
(έ�5�^$<up�' � WfS�BCD�X�6 z�%� �y�"tU �
N�G�l��,���y�@ǓPJ�br��s 풱c��y�瓍,�.a�U���\�p��yB�ʻ֙HaGS�d�L��s���y"�/S���TN����%L��y�hŦ�آ�T�~� ���y2��0>.�@����}� ���yM"<����QB�O�L�Sę��y�!A7Mw�@;sE��m����&��y2��.	���� S	��+�'�yr���@�!���L��ES`��yR��Q����,�C��yX@�	2�y"��9](]��RP���s-	?�y)L�Q"���i �@����J�y,�ޝp� �7{3u[@oE��yªڙ�P�pUe�q�����Q��y��^�t��և	�di�����y"��L���6
�'m��U�rL�y�a��[��8I�$	�8.�p2	�y���Jި�3��^5�����ɯ�y�摒+�LqY�C	)8%S�I��y�ۚA@��.��b�\��yrB��e(*�b�ΡC���Sᤋ��y�!�C�l� ��܍v��	� @B��y��ς5�����X� �� )�+�y�J�B�L�E]�I�d���)�y®�w�]X�Å5���"U��y�iʕ'���y�B� �P��E�'�y�ύ�(�vH�QB�ZR�0U� +�y��X/|}A� g�t�H�/��yR*ߦ$���ǋK'_@Z �
1�yG��Xl����\u����y"(�6g�~!c�A��s)�p�ͣ�y@XUb@Ys�I6f7�I
�!���y��̙l)|�1A�˜U��i�'�߻�y�蝽b<X1K�%I�EYZȺ�H)�y�nX`��L��GY�C�.��EZ��yh�!YO:��ƈ�f��1��"�y"�ϥQ*�H �(w�K���y��w�h���iO06p� df���yR�N��푶��3a=r��6�y
� jP���b�3ce݂R�	�a"O��D��� T|�`�f��\�X��"OƝI�`$ih�#¥�V�~���"O�!dQ���qS� K�JXSP"O�\ËՌk���)��B��`��"O��B1�+#8Hd���z�
�2"O�J�C2y?�� ��\��yB�"O����Ǜ�{��U�bOB���HB"OPȰ'��3q��,P��W9O��x�s"Oڠ����8	a��̴{r��X�"Oڰ����!�x�:�LU c�j�c�"O^��"*_aNYC�Wgf�yzV"OL�;%oX�q����D�2LZw"O���5���>��!`�d�H�"O�Y{a Ʊo=rX��ҵi�P���"O�@z�d#W�x��f�W���}:�"O�0�weا-�� ��Ţ��d"O�؂O��K���0��,n9�`q�"OK��,�h-��'(��`�HU!�y�	F�
��YQ��;YC:������y��^]�`�+�L�za)0I���yR��&�n3�]$4lY��Î��y�g�� �Dѐ��,�T	����+�yR�	��~t{S�ݏ:{5�E��y�	ٟY���SR��G��HIƠ�yҏ]i0�}�aӋ2�blk���y��݈D*N�:6 M�W��᱓��y��4a�68��OJ*Y�p�kS�ˍ�y�#ƕ�`����X+O�N�Q g��y�X�i�W��GӮU��J+�y2狡D��	2�e�0�թ7�^0�y�N
�c���㍝)�<�['�_��yr���r���C��/X#�̍�yb���fM2�2%��\�$�F헪�y�GL�n,�ɟ�S�:m��n�!�y⬌�Zƀ�'k4=�TQI��E��y�E[)���L�l�Qa�)�y���V�����<`�^؀p�}�<��!�R}����݃B#�L��Og�<���/0��Z�B�%g�2�z�@b�<�@̒�S� P[V.��:�f��� s�<Q�Ε�_��i2fG�[4��:T'Fv�<�g��4y4ف�O�s� �3ȋs�<sgG���
�k֞D�	���N�<��BB�}�x=*�.H ]�,D�(R�<���8D���s�[�����H�<QрF	B���I�]�P'A�<�0�'5d�E �_���д�[�<�Eb�:IZr]ʧK\�+*x�Kԍ�Y�<y�A6vVu{���^ʂ��@S�<A�K�I������}s����ARt�<Y�������D��5Bݬ�j��F[�<1�hR�E}�H��Ə_.z��¢�V�<��L6h�"���f�N��m:��R�<QP!�;Dx�	ƀ��Qj���m�w�<��$H �<�)���L�<���r�<)�h0K��!�!pW$���mJ�<������i�䝥��Ĳ�+G�<i��אb�6�s��%l�Ұ�#EE�<�!�Pq<�ArqΈ_�I�է�j�<PN5D aXq#ԊFc�j�"H�ȓT�ȰHY�'j��#�Ƀ!�lx�ȓd0���iJ�EfmCD���|�ȓU�f��M�4F.�[���p�M��S�? �����(�|}y�����-Y2"O�z #ّ֮[G���S�X�T"O���E���H��ׯ =DXmau"OL0 ,��Y�x�ө
�7��H33"O\IK��G�_�b���<2�l��"On��F�=,����
��Kq"O�0(CۇZ�Mxu��)!j��Y "O�,@'CN�b:b��0�8�&�c�"Oа���I&@�Z�I� ]�.� f"O��i��Y5eT�T��ܓ�)'"OV\�w&_�(>���"��kl@ё"O�U�C!�����AXi�"O�0	%��#)5V�9�F�cG�q�"OrA��:�
����
�v�K�"O���
�w,�M�Ҏ �Z��Q��"O���'�Ʊ5�m�ԇC�0��"O�%H.B�&� ��I$%���"O�����V�RV�Ee��\�� �"O主�	ӸI������{7�	2"O�e�F"P�S��(�A��e	d$R�"O�%P��Е�������>o�̹"7"O ���V�R�pX;��J1J�l!�F"O8���� �s�#�I�x�"O��� Ά	[�HR�%�Q��d��"OA lS'-p�i�A�f����$[�^�Tq 
@ۺ�i��F�H�' V��D�I���,��M��'�~���EG0��b4���s��i�'�F����ŀ6��(5H2B0���	�'g�]j��M�F�F���c>xvx��'u��0���ZΘ�ڴ$X�8�"���'��	ɮ �t��WiǮ5Z ��
�'r~�4�
\����&@x����'[,�s��K�	\8�8R���B��7�y"B�v �nȕ�ڢ�ӥ�y�)�(���{��D8�|����yEA?&��,���@.����i�4�yb��s14�(�ņ�e���K�/<�yN�`r�]z��m��%J%Ȝ�y�G�PMX-�2	!s�6Y�����y�eC).���
f��%�!`C�y��5�<����.e񀤂�� /�y��,K���WA�F��c��_#�y�O�2u6T��N;'Y�@�V��y"�Ʊ]K��p��hF� ���G�y����R��A�D�]�
Wj0%b<���嚸��H�$p���ȧp>q�ȓ[����S�K;;���4�P�}�`��|�P�X�^�Ew^P��%^$8�!�ȓ_ʅ���J�;_nU���J�4p��:7�X���*�Kٲ���2�,D�����BJ�,(�(�3@�~ ���+D�����ݴ0�b	h�DJ���'D���F��z�Ą�6!ȅ�58D����͐U��X�A�@��5(��8D�T��+��_��y!b�T	x����*D�43��!3iٕKS,4ze5�'D���@�*�~�G��:e(���7M)D�(���8&Tl�V��=F�Dx�E"D�|B�L_%�!5D�[$��+�$D�t�@�zB�\�����C7d�ru&"D��`c�-!"*��!v$�`w�4D���L;db� �	N�	� a12i1T�<�@MXJ��c��m����"Ox�y�CģF�<�Xu�qH�ʦ"O� �`r R�-M�I�����Crp�"O|Q�P� *�Y4B�Pb���"O��#ާ8#�rq��"&()�"O�Ѐ�)�X*�єI *e�x`e"O�d� %��z�<��!��;�P��"Ol,:��H<E�ɚ���O;Ĩ �"O��C�团>0��A�!@H��`e"O���q,��A�tA�xYhU"O��b�ɋ1/r��O_�=�@)"O��Ac�V8"�Z)�`��	dAl�a�"O��:A+ԀVvR���J�H4*�s2"O���_�I¢�W
�n!R@�"O��1��\&9��m%�,���t"Ot�@��#*r��"E�&+���B"O��ҕiO�8�v�s������I�&"O���af�"Ax�x2"�6D�����"O�,Tn�?4�� ����!S�؋T"O�����Lz���E�C�2�P�*V"O���5E��4��� �EӐ@���"O�x�S��-?�)85e�7���
D"O�=�6�[� ːq�#�*���D"OT���MȂ��P�UKR|�ٰ"Oj雓�A�b"&<a�*��k�,�0"Oaч��CH�9F�2<dRz�"O����љj��A@���xf�05"Of�p�ED�[t��K;bT�{�"O�0�b(��%J��A0t�B���"O��7&��r1<������b�"O�	&�G�T��42�i�q�"O<��`�<<����'ۆ�S�"O,��,�93|x@�̞�@���["Oĝ#� ��$�M֢"���2"ODz��43����˖t��aIp"O���d��,/�@�8!�Vm�
�:�"OP�Q��J�=G���$�)Cm�� "OlQlo�.���Kd�:�"O���V+\�pb�8g� �"O
Ԫe#I2���8��8:�h`Q�"O�����U� �\{ѬG�F.$���"O�D;�WD�:��D� ����6"O老U	߬04���T"�~lH5"O�@* ��"����@(K����'"O4@�&B�Z��)�/	�l���*�"O^�Hg����(DNI�L�d%��"O
]��aQ<�����L�r��eq�"O�i�)���Йb��6����"O��p���>�&< �ڎ8K
L`�"Opݫ.ޝq��(���\��7D������>svZp�'�>�v��p�5D�p{��L-B�(�2b�-9Y �*C2D�8�Q�2��"��U�C�m�$/D��1�_�Y%-*���iJ��B",D���C�½g�L�#��Xn�ػ�+D���4	��M���^��4�!b�)D�ˁ$�Y��(�O�Q�d�8�h4D��c4��d�f���*�� �&���,2D�xʤ��8�Sm!-;,%D�lT��Rv0��%A�, <�F!D�(�E!^��6��:���V�;D����0
`PtAeFِu��#U�+D� :'���kPh� nW5]�y�$)D��;�cD
/�B��%��/i��5F<D��{S˥"�p �`
,����;D�,��� ��cD(N�]Mpm��:D�� � ��E[�p��A2`����a@"O��IA�	n�޵�o؃v��AQ"O�)��-��e�p��%.B�)��`�0"O�y�	.�)۶
�K����"O2=)�A�[5��ȗ��|�>p "O�Ȩ%�.s����N�&m�ZQ�"O�(�N�(�|!�L]�NA�W�<!��/v�B�N-����COL`�<�*�4J8$�@�ė,vറ�ueW^�<�_#O�>i�J�*~�0�dZ�<1�
�t������Z#� A��|�<�`�{[�T1�膃Z9:��i@@�<�J3hsjUqq���İ6���xb�'D�t���\��a3�mMa�����'�0tP��hP�-˃�_�]� t��'F<d��� N�	�"���N�FE��'ݾ('��&v��hQ��$KȚ���' ԁӧ��@!���#?��T�'��mb���3���X�`���'���bE�4H��+�� +�'e�)�w�;9�� S�E�	}e���'r`����Ƞڤi�� hݚ���'h8��@�	:u(a���\�P�r �'���{F�!e�����X?5H hI�'�n��D�Hj���	�%�I�	�'��i� ��7T��,���X	�	�'��D[`�݂{�Т�b�v�H
�'GĐ��G�1uXj4�uI�%"�T�9
�'�����MŜd��y�D��1
�'W�Z��/��h�ŨQ�iݲ!A�'��s�a87 �qb��<_WB���'"���M�	��yJ��P����'���RbC�H5���-W �m�
�'�f�#ѢŹm+D��a��#L2��',�����2���S�۞d ��'�=2E+���줫�I�r�̻�'AhM�R�',�P��b�UȌ���'�Ε�W�B�M6)�b@�aP�'�AP�oil}�kQ*x�$� �'X2̋V��k�N��D�t����'�D��B�W�������	s����	�'j�)�a�	O�q�g�ٔ|��q��'X��["��4 �J���(�|چ�c�'}�(��A�^�|,I��9Bޞ���'��9�B'�	"	�}�V��l���

�'�0M+�+Bn��#�x|�	�'V�T���5+DYy#e�Z��,Y�'3�<��Ι�Pռ�x��K;
���'W��p�jJ�I��Ȋ�NYz����'6����KܜQ:Ь{�F;bl�'�6U�g^8�� �ɉ3����'ޖ��E
~���k��\^ah�'x��Xdg�g�����B���'/@upӢ�1d�p�i��O&l�b�B�'�ZŊ�a�t
rL�Q��-/��e�
�'������ʵ��k��v|h��'�B��W��F"[�f�,t!�}��'��ae��!j� 5q �ȷh0�i��''H�m��I����&��vV8h*	�'kn� !�O H��8f����py�'�t|р���N#�K�ʟ�[��'�,�Zc��o�Y�W �PB��J�'�6��I�#1���[BOM&y�����'�r��3� W@l��W4mz+�.D�� <���D[	3Wȅ���WA�|!Q"O�9�ʕ:@�
��p�ǧc�UB�"O�Y�&N-%��YZE��>|�"O�!{"-��TW�`�c��8���""O`0��*2{m@L�r�N�W�Z	�"O�d P�[8�x-Q"c�
��:a"O��iglĖafT`��!Gbp02"ON���<W�jt�1j���l!"O���h�<�"�	E�Z=�@1��"O �/Ib"�JQ�7@<H�b�j_��y�f��H��-�*�$8���GD	�y"c϶{���c
�.FY����y҈N�j	�tJU:z9�tY����ybd�%2��+�ʕn���!6oѹ�y���V��I����l�HHS�#���y���=g���p& �.���P@EΞ�y�-
n:vf�:)i� [�����y�)Щ'�vm+�#0ʈ B��y2�^�zUZ����ٛ(��͉AG��y���	��$�� H�#`"t���yҦK	l@Љ�6�fE��(:�yBeԒ�T���33�H �c���yrG�����1��3%vT�ʣڈ�y�$�R��|���i����,�yR�έ:���&��1�t�M\��y�Y�L�(���@N��T�ܬ�y�M��mF��ɗeD�"�2��4�:�y�	"Cڴ�rBoԏZ�Es�����yBe��^�ภGd�:Y<� �����yb�
�6T�J�eO"��u����yr!1=t���1}�p��N��y�m�%+ly�`C�<茘C"`�yr枚.��`���RGPdx���M.�yZ��C���w��Eq��
����
�'
ስ	� ?G�A�7"18���R	�'"�[q�+%<�W�>0�D���'���ځ�׆"�Pk��>4(����'�|<SD��.\�F�鉭3	��Y�'��@�>{w(��ҡœ&���#�'ќˠ��!�l���5#��Up�'}����"[b豒di�k��X�'j&�BUb��C*��č	���'�)��� o	Ze�P�GW�T�P�'���3G#����i�L�J��!�	�'�fxi��ɇ	EB��E�ƛ;�B���'A`+1�I(Ț-�؀/��[�'=*|�H�*mlZ�*�,ū26v���'W �СB�D�&��3j�%MD) �' ����:H��	f�(2>�8�'�v�bF<���A��K04�Ԉ�
�'�>��0�Zzcj�k�c�2�|�	�'LVhi�ò K@��t�L<�� ��'zB@�g�&T	��p�x0���'\<H��f\s�:e��L��w�X%Y�',���йע�K�tۦ$ځ�y���0oe���NڱD���$���y���>az-;�f�Kɜ�[���y�G�gM><p��
C�ޕ2��!�yRa�'�hXՀ�.��U
_��y"&�;�~L���=�ړ���yB)?�"�s' �-�xZs̕��y�����5���¢{���h��yR�֐+�b�c�j\�p($��G��yr�,F�^I� ��� F֭�y
� 
ͪP�v,(q�Ŏ�=��@3�"O`��!D].%2:��6�@�h ��"O�Y"��aM��y�mO�28`��'"O�� �i�8V����)��E"��A"O��k�+C�[m�d�Dg^;>p""OT�:BLӁ3�DA�@��F%�"O�Y
�|�a�R��C�x�"O��'���B��=�����Y"�"O��z�m�1Y+�1Q!i�K�R�$"O���B�^jǒ�!�NI�B�.�y���'_B��0g.F�sth�����ybꂰ	��҆��l���#N$�yr�I���d� ��0!���D���y�f�F�\���!���Bcʖ6�y�ŏ��Ҭ�C(֡f��L�҂��y�D�
`X(fhQ�e��ݚ�g��y"%�.W�H�x�а*x� a���y�KأV萀sփ9!�����'\��yb���Mfn(��	�L����$Ⱥ�yB��+~�:iڡ*�@u=K���y�'�"�@ S�m�9���[@̛��y���x�0�ӊJ�0|2,��a�;�y�cP),@bǚ=q�TM����yB�1pr����խ]:�dyfL^*�y��L�6�N�0��N��q����y���<0�ܙ�@@��`�Fh�yR�P�|ۤ2�ʐ/a\P�F����y"��5A�h1C��R�
�fF�?�yr�W�t�P#��΍A��`A&n�2�y�.��r���p�^�1�~��2���y��L�m�(q���I�/DРy5�yR�	&�8z���3&�ƹ�q,/�y�-	'	G�y��H24ѶaBQ� �y"(T���I�F�%N���eR�y��6z,��/��V��y*�ǃ0�y���=f7ҁb�kB�B��;���0�'��183#Q).�l�ʓb�(v�Ys�'b���f��>�N�����D����'�J,�0�VfG���Ő_V����'X�)1`�in.�je��P��1�'鮔� ��i8D,�ͳC(�*�'ޚM���n�X��MA�8\T��'�d<�r�R1e��%��$1�a��'�]���@�����?@�Pq�
�'K�I����:xh�UX!��;:`"���'X��K�U9���N�<1���:�'VF A�	"q\�Qv�D�[!����'�r�R��DdA��销~����'�VY8Ek�o��ip�śv{v���'�N�Csa�5{h��M[�s��T��''���a�K$ � ���	��j[���'Ț�"r�P��A�I�.Xh�	�'cD�J��Du���〫? Vxh	�'H��a�ڈ�a��#%��+�'o
������&���D�(x����'ª��"��{��`)^�&	�|{	�'����+ƫ+:BX
��O�d!	�'�1���{2lUc5)S*�1��'��b��8�|Y3��S�����'m��GM��H���۱���B�" �'�NՉ�"�&����R�9�(���'�`PF�ϬQ�`%�V�5m$���'xJr"�ԡmEXu�3��/8����'�f�+2	�mߢ�8�e�2d����� �LI6��:mY4���k�SrPq"O0<
5�_�����ĨZD�#"O��ʂ�Z#^r�AP��N�q��[p"Ofps'ηW��U��ET>m8���"O⹊VGM�Rzٹ�*¯l<�P�C"O��shE:gl��%��#*8"��g"O��SD
 �����Q6zW>���"O�iF�,s����$���=MR�;W"O�x� 	��q��T&�4��U"O�{%J�iO~�s�Y����!��'D�D�,cv����@�X�L�!�D2=��ؑm�;z Tl��	V�џ@F�� A�8i���Q+WB���,�y�
cż�!�h�S�a������?�S�O� ���4Z%���b�ب��'�,�ibaL j��a�HU�c1Լ�O�`��v؞�¨��up@e���H��b���/D��`
�gM��v�����p�F����x������aFk΁u&X������<aE+ �IxBy�L��+���G�xj:B�I�3F��$�K�,U�%���W= �^TP�����	-<J��h�臀x�Z�"�lȌ?�!��8	�F�"�	K�B� `k�0B���	�"҂�B��*2<��f�S;9�@C�I'(��Xto�53�����3��	�'W�4� G�	5�ȡ�׍U.P�"��
�'a�iBSN^3u׮���拓Y
�A
�'��aS��-.��p
Uo�V��c�'gp��F�BH �<�7!�9X5�
�'�- g�Ot�k��/
'���'L̘fl�O���z�'��}Qv{�'XJhD"߆i%�y�AJ@}����
�'���A(],i;����!#(���	�'���0�mC�C��t��0p:�
�'ظ@�!i��N(�B��\�[�'���b�V
$C�,�����	tj���'��|�B�(o�H��D�~ }�'��}3�� Q�Բ��>DfF�X
�'0p%�D��#U�`9����8�ex
�'Q
��"��q�����$�*�� a�'b�-��"d8�r�D�x}��r
�'�PD�4��u$&��r��7z�ը	�'�}x���+A��
!��w�,e;�'��\��ا8RX!�P���#ɺ��
�'��t�щͿ���z�a��5F� 	�'����i�*p� ,Q��|�� D�����*��|���(N$��D+D��!�2R�<A���HY�E(D�89wI��qH��:`ЯX<>�!�(&D�$�pA��*��E:�	Ҝ C8U�6e6D���%̿/ּ�(o�Tŀ�d3D�8�Vc9.c�0���8�0ű�d5D�h���^��p �ɧ]J��!2D�0 �c��$�DT��!G9|2E9��0D�X2��I���
�=V �� -2D�hI��ى<
��6�Cv�;��0D��x�ŉ�LC��æ�1%1@�R1d0D�D a��*bD$��e�,+:!j�/D�H�!��=���ǉߞ~��SC�"D��I���i:}x�i_�b�T��� D�h�D���m>B���O$gqP�ʅ�8D��8���v�V�I�Ü>�L9���!D�t����:ؾx2�\�!�M	�& D�h��(Q(>1<��p�ۈ^��3��!D�� �ceaR#N�"�cF��w���c"O��T̄a4��Q#�� �I�w"O���٦&"��Ԯ�,N�$�@%"ON=A#���������./�~���"O�Hr�lI��pqbҞ|&-�"O�|��, Z��L0�ֹ4~T0�"O�X5��)bZ5z�H����@"O�����N7`�A��A�~,��d"O�q*t�u  E9P�R��"O�1Ї��6�E�đ����d"O�ͳ4�ٻl�@`ڶ�8� ���"O>d�ׯѪ]l	B�gɮD��w"O����,ʹ0��\����[�j��"O6��q��I�Ip@�?](,+�"OBe���
�GǄ4�VU 6��d4"O<m�����E<�ဵ�ܡp�By{�"Oq�>�d�ԉ{�"O<LS"��m�$$U;4�I�"OJm�&�>+"�}�3I7�� 8�"Ox�;�I
 �`�&X�H��"O��r&�l�Uy� �" � -
�"OZ݈�)G�T��T-V!Q{(�X"O����U�Sdz� �Lހ@����"Oi��&�*y#�JO�'���"O��,�;f���(�H1~�0=�P"O�Q+Ì;c@��GA�=Ɛ}j7"Oz�h�/K�d+�YѲ��(l���@�"Or�A�k�k��	sc&Vs�� �"Oʌ��EԻc�vLa��b�zQQw"O6����;S-��р�� ,/d�R�"O�P��j�0���KQ�O���"ON�Y�JV.���9�
�7��	��"OJњw ן]&�AE�Z�p���	���G�0��f�i)�@8i&��� =�d�e�
�cTqO0�$����x�C�Upd��1�6 ��ұɎA� ��Im%�X ��H�z
���	�*�B�ڦ��}QF�!祅3
<InD�f�֔��C�6�����	dl�1R
#CJ1��0�M[Ŕ���i�&�%�ג����MޡP�v�	T��O�"~�I�"��]KA�!P�ɚ$`�-Ig��'�"?aӱ�U�4�M��c��k��r�*~�ܸr��[?)�T����'r�i>���n�7q��q�8"&���Ғ�y���/G� j!��~���0���;@x� �c���Ͽ۴O;�pL���;%��82[�k`� ��*�E&�Y	,�h���[0!y�H�$?ט&���+�"��H �1S�M� �6-Xs������z��i"�
TM߅ol9(%�G���Di�'���%�cAh����(�������rD-ʓid�a�^��Цm�	�?�;d�rܹ�! �4pZ�0vC\=x�CfZ��?�R�oZ\X��:��x�ʳi_�Ge�a3�R6�h�×�<�h�p�@�Q���2��T�k�oT�	�{Dö�@�VS̅���v<-K�aL�UkP�ecT�%�B�"�A�~Z�D6��$��*�,�3'u��s�m�;W� ��A�>�ï��X�ߴY�'���'��I�lYvE�rb�.HU�L�s���f�'�a}`� '[�µmȭy���e��'DhAn���M#J>����(O����"'ڕ(SD]>DT�ŘhY�5c���O���O~��(8����On���_7`��FS��� �J�l2��F�Q�P#�!�ʉ��4�;�����#�)ʓd�r<ҡ�����m�+H�z$[�k���)�"�ަI��m#wK�TѨx�&ի<C �O>i�&��X7�W
e���5�B#���"4�#8|Kܴ�?9,O��D�<Y��DÉ:u�����+E�lm�"��-�y®'#a��0R���M����Bj
�~b횞R��6-�<)�Zk����O��` #jZ��wNP�5U�P�q��O��y�m1��rA�ԷR�7G/+i`�I�^���p#S!��j�(�v��3t<�<)�F]�7�$�3�ǃ�P攬5$�*dE��*׌"R������X�4�*D*��Ex�#���?1V�i�7�O^�t�:����5FnUBE)Oq��K��'��iy���'�8���P4y_���h�y`h{��M���i]��d�������67KJ��F㖜�~B���_E�qY�'rP>���	ퟤ��ܦeSb.^�P�B�1��DHP�%���Y�-�<EHJ�:�� �Gcٞ	�|ѪA�r��|��'�5f�]�R5 	�f��:�=i�%�/�M��J>Q���ʕ��6�`���Ƞo�kK�)o��Qh䋧|�q�? �i�hIK��qJe�]��r�q�i�-��0���l�<��Z��M�&%NW��{���j��a%#�T?a�����hO�t��{���xGt��-c�N:�(O$]l��M�O>Q���u��G4$��0�֑�İr�_y�O����=L� 8  �   =   Ĵ���	��Zx+tI�:.���dC}"�ײK*<ac�ʄ��iZ�Fm��x",�9
�h7�� 0�<٩&lV�c� Y�N�HhƼ*S돖h�n�:�ܦ�Q�)L��u�'˷e�n�]�O�pX���?��ԲBDn�1��L	dp �(�T!�g�<�-TCH��I��>9�)�1��E�j��/ZD�"�Qzz]2�
�8E�d�FM�lJ��p�,������!�v˓4&���k��-�`B�i�3#��]`aEH�
���J<Au�ޟ=\iO|�h�*��0B�LK�)�n���Hp-.8�7F٣��	�T^��H_2T/�I���؉C�_>e��.��q&�(VEڅQ_�e��G�%/����
k��*�Eþ3K�D;�D��/4��sh<R�&_�Q�ֵq"J�#I6���H�+��hM�ۓ&>mЌ�L�T��G_ZȬ��F���eoɏ �p
����n�J�<a�bTY��SҀc���'d?��D�
�7�vȄ�WI ��ɶ�`�+O4<���z�хK/���g�4͠dǌ	2,Ʊ�sΜ)������Ew��<>c�CC:(��(�'dм������'=��)�j� L9ީ����;��4xz�$ �T0�O��i��������>�O#ג�����PՐA��N�MfT0��}�'m�D�J�����|"�R�D��sQD�$0<e-E9}����S�_d�	;8��e5���3Y�r�SQ0O.� �N� ��5�WaT$1��	�q^���&��)-���OHdx`��'��'�(�ha�&,	u ]�2��3�(ȟ� 6�`����{��u P!YU?IA1OZ�Pщ\�����[9��퓥b>�1��+w�V����;G�E0r�BC��z���� "6��4�rހa�'�: ��*x��ِD
��Y.O|h�a)=M(�'�Ak1)�9�ēGq�����܌/f�I
&��p&�h0�Y�gAj�%��I@HM�OS�c��x�(H�e��T�3��F$��9u���nJ���KV�x  @�?  @�?Fh�� gO��V���"OP"���~D)yp�G()V�!"O0�[f^-�� c&���2K&��"O��&�B+\I;G)@�z+ʹ�#"OH��c�	���������f"O�|���n!6	qsn���@U"O>�+�K���
U�B/�굹t"O�`�%e�"NưX�*�-t��d"O��SVE2$   �  1  u  �   '  H-  �3  �7   Ĵ���	����Zv)���Hc���KB&<��N�3T���1ѡ�;A~@p�d����)C�'ll\�02��o�c��%��ϤV��9�y��y�L�"�@��=�~i�F��^���/ uz`h�cȸ	IŻ&�5# 	@Z�f�$C?tv
A���Yθ����s�öH��   �x&U�"O�� �4f�l9���B�:��#��(���J�9p@���K=�A�h�$2�|����[�`X � T
���p�-3�}�%�'GB�'��~ݹ���P��!�T�.%�����_.D�R�
`+&zw�uc$�mg�Ysg��1���!�	F`��Q(�Y�$�DbI%M�D��c��'������B)yH��E�Ib���I�z�x���虾����P�L���d�N|��П��Iv����tD�����8`�H|`t�t�\��y�`�2n��`Edؾun�Is���M�1�i>��	xy��ܵTڸe��L�I�A�ԊڟfbP�!�Ҡ?qR�'�"�'���؟��I�|§��%Z��8 p��S�ހ��GK�a�D�iiR0�pL�S�F�i����	5H�P��G�M�0�$��Ζ$� M�I�7��	��:�4�lZ�i��r�I��F�����p:�e$eWtXQ7h[ H�(�mZS�'NQ������!��	Cj� ��`/?D��ȅ�O:  D6a�bE,�*�>���i�U��c!����I�O��S���k���sW��@�!Ĭ:r�7�IT	�D�O��D�#'}F�!�"M"�j�h�L��`�ΧK@�Y��τ(+\���]?e�5G{≞B�zmKB�p3�`�%	W�@��	�,Iz�p�ʜ~'�X�d%K�Pў\Y��O���&��v7`ҥ�B�NHl)g
;N�X꓏?I
�>� �6&�6x2H���L�X��	��I&��$Ҿ'j�i�G�a��5�W����^L;ݴ�?�����鎩Itb��O^l���P���JS	�I[*�bQ�C��Y
R�ۄj���5�e@
8É8:D�9�f`SŖR�� �m� 9�E��P��&��5�3 ʉ z�4�R��1K8x����<>�>qP��[���c�.�T���ПĨu��O>�m�������?�� F�)|�E8���/�*��J�<I@
�(9�v�(7Ɲ�S5.� 5�D�'��#�&J�[e�˵%�	e%9�GW5v ���'�ro�52�態��'���'���oݑ�	�2�Zջ�*�-mt�m� :r�;֩�))� {g�i�����á�MkE�O�ah���ēL����Ո7�8�*��x�N��W+@�P)P�*�����qvn�Df�17ߔ$���+#���V�UB3��Tu;F�����	UX���GŦ�I<��?��'�HA.%=����J٪xO�>��"��<�s*��ܸ0lK�x��A�it�6���y$�8���?Q�'��ѩ��T�R�
�;�� �K�N��/;���5�'K��'�"�w����џ��'7���P�1z�ۣ@_���Ԑ4ʯ+B�U#�$d�����b,��9ʓ6z){�%Y?5y2�CĨ� gu���7�!w�>�A�f����6%ԁ �0�
3�P��(O ����'E��pEC�w�b�:S$0}�<�GDo����1�	��M�lD>	v�(�@�&k4��ª`X��FybU���}��M�(ZƦQa�S������Sy���mp��'�?��O�Щ[�&�����R��N�`�Ŋ�4�n���?���P�qz�.K�H]j��lR�+��F���i�*�xCᓣ;�j���VJ�\�<!�OK�/�8�2@��:��X��44��-����Z�~@
vN��lB=R��Z�<��#=Q$E���IF�'W�8�5aʹ�R}Q�I)l���'P�~"k���+��"0�!�-�>����L�fA�_ƌ�'�F8U�D)r�>	��+~6�F�'rU>ӥ������}��,�%˒�<� !�a����4-���ベSn��p3J��?�*���g}�k��+���)w�8�Dy�e�?)-P�b7(��K��nb*���M��+� !`��"�ӕ��4�mM�X��c��P�`,���@�������#,O�T�S>�,Ta�EÁ`n���ga�k�P�'@B�|�i݁�p%� ��i�ƈ\��61�g�1�s���e��OX��J�J��A{�GV*U�X�`'��}�� n�����	��w�\ߟ����|��3�u��'���Y���M28��Ǝ-?i2tQ�獇U3�qG$��[s�܂a�OF�'&D�Ȁ�+�ؒz�b��G���:}@��[�z�Ӆj�)f�

F��=��l`�l�!��O$8;H<�#`Oȝb�h��I�%���]y��#�?���i��"=q�'���Qg�K�\% "�[qh�+
�'@9��hB�O1�u��m�R�AJڴx���П<�'7�X �4h�&���̗.-�XX"��(B&ua�i�O����O���Ǻ���?��O�֑q2Ǘ/~���f`�0�j�#@��+>���2�Y0Sj���3��%9qR8C Ȝ@�'����T�d��H� Ы>,�p�C=4��g/g�=����|K�`q��P�'v�	��2e���ӏ�'ovp��B�@�d�J�i3�#=��$�v̐�	��qn����{A!��zļ�B�;3k^�"u�":�	��M;�����QiN�nZ۟x��^r�OC�, �e�"(E�LVa���B@�ޟD��ß���9��XhC�y$@��S��.\�B��
Ը!�­��)Gؘ;C*ͦT�<q�Jԡ!΂���3�R�r �&c��]R	� ��7Nބ�&��V�~4����p�'�B3��G�>��u�κ��x@pB�dZ̒-2D�l����]I�,�
�t�R0�Ob�';l�:���
㺔z�mبc�]+�O�� �`����埔�O�b	:��'�2�L�a��c%`��l�C��e/�7-��J������d���Ѡ�ϡ5�����̎�G�c>EI׈H5N	x5��@s��820� ���gZ�V,Ќ0/G>4C�۔�D.Nh��q%���"����th_�"@jt(r�M�Q h�D�H���'��)�I�ON��37�1g���<x��⊍�l'
C��/8�x���2JkZ����0��"=9#�S!N5#����=`&|3𡞰%�JU0۴�?��i�Da�A�X��?1��?����k��Y�g_:��$�߀_VPr�ӟ-��偼���kb'�"$/l��	�� �H��7�<�zV��&�4qy�ˈ�U��8p.oӀ��4�֦./��01��F�Ď�b�d�O�30A��"e��H5m���_��p�M�O��D"ړ�~�o_27G����11�<\� eS#�y"GQ+@2QA�EՄ4�,��F7�M���i>U��By�@�X�N��'�X�cZx"k����X�l�~3r�'���'v��Οt���|�ˍ�g�Y	��P���B0
�5'r���"*ɗv;��ȢK[�6�z�Z�!��N�<�#jɎvU�m�AHˀtJ���:l�Ȉ�à˶z�8����|J2y����cf�<�pfF��$+����y��T���^TH���Œ#�y"��0y`h@@ǢFѬ8��J<�y�Kc�Խ��	�q^�]�AM.��ئ�$�p��a������O���;TA�q;�@0(��*f�Dh+�7�C�C�����O�d�F��t[7LP�84��:V�ڒ��Χ-��yՍ�;W�
�"�.�="��G{ʗ��ے�Q u�T!˗Ɉ�Q���B�Ĵ�uF*����w� �ў �!��O��8AZ�C��ɾ{j(q����K��꓆?i�)!�l#6�%P�!�	4?X��ɭ���āp}��&+�6[�B�`��.i�� ^�����џ��Ii��@�>GR�'��<�A�r����ʃ<��q���h��a��_��q�B	�r@rg���u�BטOev��FA�f�90� �tUH��'S��c���lp�h�#�%S�˒�=���+��OD�ӃF���I��d�6���ap�':`��JEɧ��z����)@��I �ܰM�r��.7D����%7nV ��%HtjԠC�)ғE��?}�e&��70�T�W�B�]�B����&�YzA^u���ğm��7+F�5
�$	b�Xr!�D�v3� k2�WP)� ���Щ!��*�x�0����`rV��3�!�d�*og`@8�HB5����F+�!��G�-�x�Q�{�44�%Fr�!������~�$��'���� -c
�'f��P�מ7�^���+���)
�'�~�k� X�f����v������'I�\9�� �4�R�\�70��'?<�KA�Ő;
�!�����-j��H�'0Iá��K[���͐/��Z�'��q�o�.@ܸ01��O��8��'1�Ѐ�	�<C85:�/ēH���8�'}����ֵ�*L�C�G�@a�@r�'�L���KF*F�2�S z��I��'���1f�=�~��B�CG��3�'����`+�R�d늏����'_���V��@� �`\�x�*���'��$ِM�_�Xa�g�@8c$2̹�'�x�c�55�'j�
*X��'�D��#�M��1�B@� 頸�	�'JH����Z�c� �ۃ䓐�y�ܲu��*Ԣ+Y��0�HI"�y"O,�ixb�#X�T������y+�M��jP�]�P'j-C&��yRF j���QA��:HI��h�y�L�=A`�(�5��:WP� Q6&]��y��*�˦.�]���F^CC�I�0�| ʂ���%��U��î�C�ɮ'_
�C��V�B�e�QI]�@�@B�	�n��G����P�f�EA[�B�)� ��"��Ů"Z���� aK�� "O�S0K�=�A��$.U�����"OH-IƀR=U -���-�q�"OD躧&�e<tڡnH'iE�,��"O8�06*�@P�y�b�/e��)W"OR���N�n�|9� ʟg�a�"O,���n��U��s��T�	�5�"O��ڃ!'3U�L���'^����7"O�]Q
űe�9:��P�!v\B"O[샓�H�b�C2:�;r"ON�U+M.B=�h��wĔ�"Oxc�,E'kH��;b	r���"O�ȹs���-��`�T��;u"O�]�1�$0���c-��s��;"O�4KB͔ Сh�΅ur4�9d"O��x�.��*�����W4di��"O�T�1$L4GH9a�c���$�JR"OH�� �/b��#؝O�*��"O��:�b�����VA�o���J2"O0`�F�_�[�B��K�Fq��["O�1�N�/ۂu
���%Rp�t"O�Y�Ӓ�ltS��Z�8AJ�5"O@�S��^#i�!"F��D8�"O̠h�K:��<��NX/0jؓ�"O���C��;` ��Zvndq�"O�\h�o\C.��G»'�`��"O!�R�Իv�~�@���"OR��%��Z�Ie$	/<�b�"O4�Cb)�v���͜�|��E�"O�P��ɩ楀fj�;Zg�#3"O�87(ȫ3���i[�;NF "O�2�"�.1�|��3�J�S�f��C"O�:g��
s��9��B7G���
�"O
x�䀔�E��H�JR����"OR��'�;%�VE�Sʜ�y�Z��7"O0��T�* �0ـ�7E� lSg"O�e�b�3!7L��4 �5*�̡w"O��A�@Z�ԽŁ��aX8�c"O����Ϲ(Nq"�!! �Z�"O<3�o�dB}ek��0�� �V"OT|�ւŜP���K֫(ר���"O��۶ѩP��i
&j@�kD���"O����EQ�y��i�w�RGO�l�d"O2)bco��6.(p*�`Ϸ?�����"O��を�jD��K3�J� ��Q:�"OR��Gg�m�t��
U<���u"OR3�ʛq���+��ܤpn���"O���9[!�P+���$2�"O�٪�ʘ��6�	��F/\V|a"O�\�C���
�9�A�/�9��"O� ��H�#T���5�ÍX`��"O𼫓	�4"!��T*AvJ�S�"O�͒A��C�r]!�@�"dY�k4"O�Q�c�11��!I������"O�y�m�3�T�f�+�H�"O�h�t(�}t���K�.��"O�\����{��*��}"i��"O(5�6
�D*���E��!��"O<=�V*-Q���&�p��, �"Oj�C�3Bv�����ϣAOv��"O�պ�%׮-,2P���`�X��"O�8iპ%l"=*@���$ճ"OP<xW�Y��!��� �G���ؑ"O�I@V�΋ɈUb�ˌ�?ORyB4"O� �򁥏7Rv����Y��@0B"O�)�GI˨f��=�q��)���&"O��y�@ښ>����M�qƈyR4"O�lƃ��C=�Xqơ��6'�h�"O�J����IPz-��A#����e"O�Xaņ@I~��%���3�b��"O>8{2$o�����c��}��"O�)�PM[=]K>-z��H��
��"O �K�^6f^���!έ
�x���"O.h@0��;���W8w>a�S"O| ��xLc��D�N9�bC"O���O�b���$L%X2� b�"O�I7���tua��ɫO-"< A"O|��`���S���Rh[�\��"O:t�vL0L�R���"[���"O�L�`E�g��mFP@�4�"Oܘ���θ=�<��$aں�ؖ"O6��ұK8ySd�@�<�@�Y`"OD���J
`P����$p�uh�"Of=a2�j��ivf��\]kr"O�|�!o��0�eS�3%h��p"OT��'�f�|��!`#�0�"O�|��ƅ�-D��ҋƄ%6@�"O�KU�E�O3�	��F��ȑ"O��lM(>!t,�*��3&<��"O�eB0�!�D%y���;;	��''N��sK<w��A�ՠ��N���Y	�'�9�a�B��l�w�Y�A���'o�pEV�6���>7��H�'{�yk!n��~��[6�	d2ͫ�'{��"�̏/,�fͻrJX�-��'�A��d�1AW�Hzs@��B<d���'PdB�ԭ:�C���;}	�A�'�~�r�Fd(訲LYu�v0+�'���,pb�M)�0$3���'��<E8"���q�*[����	�'ElX��Aݔ_0!��	2��'�|U�!��r��x����K���{�'��\� ��$�hu�w˦�(�'������k�`�ل-+A���'�m�� <q�����C:g=��Z�'����@Nf(y�ɁW:$�#�'��5��m��2D,�6�K�>�vѨ�'�"���aN�.����̗1!T�!�'ϔ�۵DJ�I�1���5"<�x�'G�% ���2~`MI 䉤VEt���'3t�5 �dHa#dÈK�F�
�'��9F�e���r�C;xftm��'�!#��Wxr���G�tZ���'?H��S?�(��-=��HY�'E�Q���~�+�Y0_[�$/D� ����\#0�t��$hD֜�ì(D���&cR)c�����?���Z�6D�t�*@�:�$-�@B�%R�C�4D��r�DX�Y��T�J�]4D���2D�l�%d�3I�j�Ac�.2��a�.D�t{��J�I��2��X"[bE,D�+S,
8VR U�%�Ԕl�TX	��>D� �
�-*!� �i�	qoN0� D��{�石6_��Q�/*�Z0�"D��Q��5"]dI�S����r�,D�	�Û ���q!�B*���{�N>D�\��	� ��s���8���h�;D�И@g�D!Fq筟�tu�At`'D�� ()*���y�v��a얟D)jy��"O IR�S�u�R¥b_O:�1"O2�#P%�i����#�O�p��"OPH�3b�9U�l�FlV:$�H"O$�eS�rr�:��.R.���p"O�e[A*P0B�Dad��%�Ȣv"Oz1���%y$��@�W�D��5�B"OP8�Rk�|��uh���= Ւ16"O���V"5㎈�/G�H�(TjD"O��f��SV�}ؐP��"Ov {��#s���ڵ�؝c��U��"O�T��Q	k?Vd�Dj~5X�"O~�A��.Yd9P L!nj��4"O��Q��	p�@�3 �,Q�5��"O�8ED�o�L�c��!8��ݘV"O�R2D�r�>�{E����"OQ)˔8oJ����\�za�V"O��Ҩ�gU����+T�>��"O�!S끴rM���eJ��]#j���"O��w�ɱ\�n�2 i�$���"O���D��2t��f�N[��
�"O��H�nQ�}��\"��
?h���"OB��F���7�h���ʇ[UV���"O����Xn���ЮG��`H�"O��׏��$\3Ԍ��.���Z�"Oi�FlÑ
�f�R��!?ʱ+'"O�x�6�6�X��$�JO �"Od��&_3/� 6��c� �$�%D�4C5�X!�X�X�VK*7B�I�<Qch�E��H�,:���jU�	{�<g��!:hp����DY�����t�<�,�"n�� j���}B���"*WN�<�я\;X\�j�,���OT�<��D�#���I��@sZ�2���P�<y�K�^�rbȖ�b��ի`-�p�<]+3=��A�+�%XI��ҋVG�<�S�.k����y�a*��E��SdI�&�a}�!��Z���jC�W?O)tHb�W�y���O/^� $ ˰CUV ��e��y�(4��ӣ-�4G>u �Q)�yr�W1�<��D�.�!��'J��yR�ʁ"܎�H�"ƿ(W~� eA��y"��"8֐����m��f��y�G'=� �K�� �h���I
�y����ma�)�|�8@Zҭо�y� W�JF@��b+�s�X5XU���yc\�|MB�D)x��������y��v�����#�i��s�O��y��W�:�#7풾g���#B��y2�8]���N�2sҜ����y���>�� � �8 *t���O��yO�(� �rN�wV�T�2���yr�#++*��(�$�.�rb�/�y��*vs�� W1��Ô���y��E�+GF=)�S:d����ߢ�yb.Z�Ǵa�҈�?��3o�-�y�,'&5�D�9(\����H��y���7U�X:�AN%-�n��7l��y��ͅ�ؔ����wbL��WG^��y�L� X.�ʃ�̞v���1���yI�CU,Lb�b�&E���ګ�yba�%AtAõ�H�\�y;�AX��y�d�k�
���Y�N  /��y2���'v�YkSk��R9LL�g�7�y
� �1:U��%�]��G�3ܰqk�"O���T���+�e��#Ь)�8A�"ORq���V9eV,��`�oǼ�"O�d�(�s.�3 Hi�te!U"O�C�)B�9Rp���3�*�"O�hR�������P�΢e��p1�"O�i 1�B�@a����4k�4թ�"O��@#���i�X�Oc��l#%"O�0o�v>�����)\�(�xp"Od��rd�Ut�'�Ԅ^S&1�"O|L�b�8�0đСS�gڄ%"O̔!Sh��JK��� �۵e��q�"O88j�gٴ�6�2cFǱ]�v�8c"O҄���d� ��D�
6Ԡ5"OVVCJ�.E���-Y2���f"ON���	�'${�����>����"O�t8�HV�~�zC��Le��"O��	`��u�*@���۔`T��S�"O>H���	H���UEK!
R`�D"O��珥Ú�@7�Ϭ#ZY��"O���ZU��I3�_av�� "Oθ"C��.rb�@\Pp�-�s"O~]`�BϞu ����,	 Ai�� "O6��ܯZZj+�7zS�E�a"OPly�cO\
�`�b��E<H�"Of�bt	�ˊ/kb�T�f"OZ	�/
�zh���A��YG"O>l��-t�c�/�+0#(|a6"O �p㘸6}��ꔉ�!��:A"O`-pV�[�W�.����"O?j���"O<�2�CKe���ڦ��28�hiY�"O~,+#� k(��+"��\�'"O�e�ц��h�^��V�N�x�D�"O��tcX=C���4*C8S�̝�!"O$AwJ^�&vpdY��6l��ʃ"O��`eԺ96�M��J�w��<��"OʝѢ���mV(+��$9��)j$"O�P�R@B�t��pÅ�0� �Q�"Oӑ���^��1�j�R�l	��"O`JWN�	n���	s���>A�"O�PZpB�'��Yv��ejx)6"O~L��M+9�C0�,1�����"OL��u	�����p��&gzNA��"O�5D�$�ʍa��ɤ1_�Q�T"OF�y@H�;�`�R O�k+v�Y�"O�5�#.�,���VMG6�AT"O����.I�) �ȆS�h+�"O,�ᕣJ�uj2�y�k�C� !��"OX=���y��4���q|��J�"O��z�e�$�,���[vʥ�T"OX}a��(E��"�I�m<�2#"Ol�GAE6W�ĩ�g�T>X��"Ob���d�;� %Z���1mD&���"O�	�G�N�A����C�		4�c"O`Q�W.�{��T�"`A�a[�]a�"Or���O��<q�����!A]�{$"Op�j��@�*$�����yR�Y"O��s��t��A�#FM���"O*�s�ͨ6	�\`vN�V�y�"ON�eE=y� k�MF*
�^�	3"O�̋��xq�Y Q#�Mь(�"OU!�9� �3b�Y4Z���8�"Oxlqq'�Wa��qcW	E�����"O� ���_|#���,يX�Fd�6"O� �U�s���)�ܹA�*͍VO �
�"O�Q��$֛E�|�j�l�WBh�Xt"O�\��4&j(YS��.<>��"O��� 	`X$���B�V呤"Oִ"�h �I��l�@a
*6�
���"O�l�BҺJT�{�oر3S�1�t"OZ�����0=��
��� .i0��"O��3��o�8�SVk�W�m"O� ��L 6����(�;�nT�d"OZ\�v#�2�biSi�0%ґ�"O��h�#Ӟx ���gF�7C��P�"O���g���J�P0k��	�3�$��"O��`�D۪SD����ͳ4!��*5"O�Hc���$���u!�R�a "O�M�FI�?s0�:F�^v��'"O���Q��9u��m�4�ɴQlE�"O԰;&��kѪ� �ʙEN��x�"O�@肿]���{���C8� ��+�S��Ռ&@��� �0yJՙfL =%�!��ֳ��4�tF͗�BYp�@�%p��=E��'r����  ��}��*҂I�I:�'����7�\�n�&Kw���'��B+�"�@B��X�_��F����=Y����g�qb��"r�)�$wo�B䉋j������9�j� �%K���#?��I#`UZܚR
R *@�����)!�!�V�d����A�
>*��a��A���(O?ٓs�[�^ �!#Â����d>D�8qTB��7?&�G_?Kz��Y��OD� D=�OP̡�k��R�� �IV�;!�'���<=ANm¦NMZh ��Ew�B�IX����
H&Ht�*�1���>�����}Zȴ�����h�Κ��\B�I� 6n�5�M)2�&�Zv*Z�3�NB�ɏp2j�KT)iʶ@&`�m��C�ɵ!��(�Ι�3n�I�k�#��C�ɋ+>6�H'l�'@��*� P'�C�IL���ޗb���tF��xn!��*=۩T�K�7ErV��_!�]�XZ.}��a�,p,XQ���n*!�$1/�"-	
͊=tp��V.=�!�	�$��t#w͋L�F	�a�J�!���BS�d��	̯k�|��I��f!��ā0���@�`���f�!e!�$@�;M�a��IN��#fM6G!�$�?��8@���@���#P-Y�!����@��܏8�����9 !��ш7,z���MM��\��G���Ռf
Ud� ]�ڀ+MQ8�yb�� :V| �ecC�W��-����1�yB�Y�}�>�3��#�}��5�yR!#?&����-9�rL%�ye�
Z[b�3b�'~��$�1N��y2�;(8K�ݸ*�x���S�y��#�I�q�(�rx� i���y���Rj\4!�#��T`�[ ��y2��Z�l1����H������yB��j���`dB����B���!���2b���6DZ��I��M!򄔼 6���mN�Xq�"UA�eL!��DAR"�ʮ*X��# X�v=!�D�GnDd�3$%� �F۫T!�dH�|��|s�@�oH2��^�B!�D����ss��8m��tk�+/
�!�� tI9V�N��j���m�>�v �"O�- 5���m��:UN�"h�ȅʡ"O(�#��ڭ7ʬ���06O�X�#"O�S��R�SP0T��ЛJ���"O~ܫ��Ov��,8�Y5ϸi;�"O���QKծp��jG�9g�pÀ"O�B�^�+ѠdR����k�"H�"O@<CS@^3h�NM q�=p�1Z�"O��j�œ>�.b�c]/5Yt�@E"O,!��B��CƲ%��A��CJԬr�"O 1�שE�(��
��O v0����"O�j�锢X#pu����e0Z�6"O&H�nX+f�L�Ѓ��'-��*�"Oy�SBA�p��CT��6>�H��"O����	�Xͼ c�_�!�~��f"O$xS*�X ��V�Vqd�m�c"Oʩ���H�<yҡ��-(A�"O ���LO�mAQ  q�8-��"O,��	�;f(���X,0NJA+�"O���:�2u�-ޡYF��v"Or�B��ރf<��P�Z�</�]"O4��!���$r�c>&�X�P"Op�I����nH��λXf�C "O�4Kel�xFH�*�y"E�"Ol�:��m�vS�␄U����"O����1.�M&��?���"OF��@@R�_������(��5G"O�<��+Z�IJl��#M�xSp�#�"O\�ȑʘ�|�)Y¥��CN��2"O���ҵ�~-��^�V`̌ڵ"O"lc��ƒy����EcB6�5�&"O�P��Gc�m�b$���δ�"Ov�rm�EE6H��/3m�UQw"OL��D�f�ҁ�aĕ-XL1"O�0'�X�_\]���	V����"O�ʤ��8�,mkUB�!��$�P"O� FX0J��[��$�R��"O��
�I�.WZ:5���8z~�h�"O����	�kcz�r��6;tf�@�"Op�!��9\��c֦��Rj���"O�r����@�[��p�r��S"O�AJ�  �   9   Ĵ���	�����t��?���dC}"�ײK*<ac�ʄ��iZ�Fm��x��8
�h7��H���rя�+�l�WOL(d��4V%��0�K���Q%����uG�	za�	��IX���?��IA!L�p1��3r�Pr�,��OȌ8�A�<���]�g`:�>�be�W�<y�DD�6����GB�M6�5��ON�� "���p��=��˓{|�9Yb�
6�B�S@9*p��R=�I���$Ő��C!�!<P�1M<����LNL�(K|��s0 �2"GW)��ԭ����%�Q'���ɧ'�P��0�� t�I�B+U�Z�l������0����Bj	9%��]�r�ߚw���2qFq�B������Z�X��+��;���|��(�`�J6i3�� �fv2�8!��ߚi�N��!�jV�4�N���g�Q�#�L� ޼YY�ᄎ�peQ�Kn���'C\YjG��By�O�0��y������Y1d	�,8G���%X��?�eb�h�剾-��!�

���OH�M<���q`F�#eB�ɳ�\)V
`y�*�>Q�D�O�]�����DH�?��o�1h���˟Qu�!��A�<l��U�RN�����9u�[���=X��*�$	^���'�،�7��g:UB�.�����e) 1u-�2��d�ӟ����\$o�R�O�D��ػBXACо�bx3 �"���K>A�o�� ��&��X�d��H��. �\i(�՚Yh� v���e���B�����Ge�	�O���*-�ۛ3������?}�^�SM�3Mֈ�2�~��:O�m���P��uqE(��@�'6����,1"�|�#C�����G
]17�l�sB��G�8�2э�� #3�̐Gь����������Ox=rٴ8)D9S6J�M�|�!��M)]�`��'�H��B��� #\�٤��g��h�0����&K��b.��>�*��BC�4�̓O���Ɂ=�1O*���K� DVqs�IJ%q�P��Nɂp��C�	h��  ��4�2\��n]�/T�s5Op�X���OD@����T���$�O~���OB�)�Ok̖�RV����Bߎ@�����&r�ɚJW����W��*�8VN���l(�o	 n剨B���d�`$��҅2��h���;:��H��D�r��x;éM4wHː͆77�\ES�"O�I[��M�}aҠ���F 7Y��y&�i�"=�'��(��T��+��8�!Bu+S�K�@$�L)+�6X����?����?Q'������O�����DO$�V<���'6˜`�b&K<Q�=����=4�I�V���"-~���lZ�:�����Z�:�Ri�b
��ì
�{C�l����so�C��T\��G�Nt�X0:E`�׎C�ɱ|�q�H�B�2̠2�݉T�J�8���|"�4m�7��O����?�u%[�g����G� �
�����~�ֵ����O<���O0�����Oxc���>dB��0Ä+X?��/�'�ģ=)E��I�O���K�+Q.�����i�:0]R����&e��"�'M�R�I�n��QJν[�%�Y��x�ȓM%~�z�o�!���!����5��=���������"�0w-h�k���ɼl����۴�?�����ۀmL��O<��2��t(~ȉ7$�]�9��B���b��֟`�<���'�\��/1����e�<s<����HaGx����`R�PRf�}M�yC�8s�(��%cR�8��63x����b���<� �Ӄ5 ��Rj�� V�ȆkX���f[�?o"=���iM��=�d�V
\�KM6U�Xil��0�	�[�$Q�o��8������	�u���5	ѨiJu��{5.�zf���M��M�0���Ɉ�j��:��'ﲙXsJ�*9���f?y4�,��	V��~a1^sf�0�d����Ɉ�IU%XI<�A߮~�؀
���S�fE�����Q@Bt�	��M[�^>˓�?1�'��Dj�0^�h��bF�f�<����3O$p�	�#S��P����YW��8&�i�7͖��%������?ɗ'Y �)�ҧD��P��aޜEd�6� ih�k��'*R�'��nݍ��ɟ�� u|���� �z�Cm��=A1�2:��U@d�S�d�����ĤAlP�ǬW7X��0P�g��p� � X�4��E��7Y��3������^o*��9c
]�G��#E��p(�g_/'�`6�P��П��	Q�S����"���z�d�;sJ�ʄ�
�ē�p>��m5M'ʉ(6�E�3Z�y5�J}r�{�Jl�ry�	�*a���?��O�`*�J��xɲ�I'lǉN;�`�4l{�R���?9�$s�	�u�#B��5 ��Ն�DH�4�ր�2��t��֖x~��2r�	�5Z$K�=<�2�ڶ'T�]�Nl�'XZ�QX��YZ��R��1u�uD{�a��?!����OH|hz�ɴr��zE�?��)�O��$5�OS7�mE�}Yp�L/F�:�2��'s �*(,\�l͌{�viW����'�a1��h�����O�ʧ38l�#���?�s��M:�x�疵.�ؓC��8���(�,l��	Q��0����'��O:~�V�ԭk���o]�n�4�'֎Å�]�����E�G�iߚ�ѕ�S!b�>\k��T5=X��h8Q�	4�����O��S�S�l��4#nL	�����c�L8dT��\R|X90,( ��+�͍�6 j�Dz��8�V:�1d�On 0��$cҰi2�'��Q�@�X�`AR�'g�'�v�]ӟ�2��X#p���Y3u����O�m͊��EN�{z�2�Z�S{X8a-��"<�⌄��0F�ӆF���#PB�n�����RF��	�iD%q���O|�ī���;����u-/	A$�˴��<�N���$��՟��?�OW���Afb(4hE�G�Ԓ�'[�]��f�N0x3���f��4Α��S��\�'��`x� KΔTa����H1�4$r(�&i�O��$�O���ͺ{���?I�O2V�Q����P,��s�";h�&�8�/�%�����Y�1�+�#�џ���������G]���RO�����갡�J��-	����XF����?��� FH�KS�m��ؠ1���B�*��i_��D)��]�3���52r;fگ+��m�"�;D��#���1{D�
FHf�1��>!Խi��W���0"�#����O��;r6����$P��0.��q
7�E27*�$�O�DõG~�$@pa�(c�|S0c�/N����'ڹ���q1�	���0\�^MD{��A�q8 dX[5`|c�JY'g��|�`��@�J6H��i�eў�9��O���+;VX ɝ5�Z��g�ܭQѤ��?��	��ݰA�ݴl�9u�2YZ�̄�	����C-{-D�ؖ�԰i��	���̓0��:P&"U�ܴ�?a����;Y�4�$�O,��%�2�~)���l` j�ʦ%�T�4s��р���!B�
S6�-��C�'e��y�!Fo�9��ڢa9�6�4�7 � ���B+t�x��.�r <�>�8�f�8qs(`�o^M�X�F��ܟ�7��OV�D2?%?=�	V?1�ǟ�Cw>�cB'Ɩ!�-�Á`�<ٷ!Z�<�6�[w��1�8� �G�';�#�V� r���a1�$�8�Q��f�'f�o�!2I��'��'�Ҫ}����?t�V=�@��!?�p!t�>Z��ᰔmѷ<"�B�B�]���֕�� [�	�J��c��ȱ��*�$ ʖk[+��@�k�=zP1���}���	�EPyQTJ #�����Ny˓H�P����0=�D�~<����3t���^�<���S��%ң��!?l8�@�֦����4��O,U�b��`v,��:u�����OI��4#BF�O��d�O���Y���?ٝOZԨA��/m���L��DC���C�"aLC��[L���cׂ1�6A�(O�� �(�&������'���(T���z<�1h�Q�����x���npPQ�L!��O
QGh��M�ҥ+�۫n��C�)	[�<1�P,~,e�b+����U�Yp�<�T��k
��`F��ND��b���S}�B{�:�O���%����]�Iٟ(�����ї-�nsL��jP�d��dl�����	럌�I/L� �]�jdK�Q,r�j�ӄ܄60�X �$C�W܂<��A55�NШ��"�)0��w"��d��š��㎘Dـ�X�j��:2"�&UX{`�5��\��ɤ��*9�`C�?	f$�Y#M޾w8�q"O @{b���S�5ȄΦ�L�"��'����!P��#fR0��lQ�h���'I \+P�i����OxʧJ�R<��?�gή)���9�&��-��yH�m�p�6D�����QP��4+�vS�H�g5�͢0��"Z1��aE9��xk4!BR�y:���O�(��Ϗ�V|�hvÒ<W��X��ɢ=�.�7��V�C%j��>���%<���H���OXH�s�'���O?����1��0���Ksl\#���y�<��kP�$z�9J5�ǧ,T��CC�i�'e�"ԇ��v�f�/��-#&�����&�''� 2�F��#�'��'2�{ݹ�i��z!Tt�|3A�@�9��{��_�7@�]SA/*�Ҕ�"�����'�O��u⍸#3�#w�1�@@¯�sH:X2��e=��g!Ε4DN,�O`�4#��!"\���ʆ�`=t����<I��V���Iȟ��?��O�����x��@k�( �x���'p��P'�1h��)�d���Bݴb����ޟ�'3�u�ekM",mT�2shL�,H�Î�bI��'���'��%ݱ�	ͧspl٨T� fmH���"��px�τ$N����N�5C≉��C�������%�S��P���7�a�J�j
���T,[X(�|
vAZ�"��Ѕ�E�~�p��v�!�oDx�I�"�t��a�;  ġׄ4=�M�ݴ�?A���s�\I�a�o�X!�M�}O8چ�'�Q����B�á��h�H�Y5E�>��i�Y�������M���?i�O�ȡ[���){�Yr��I�V���4f��ɂ���?���p��5.�?H:. RشWF�e�fI����S�ڱyv�Y:�ͩl�6ȁp�G�b�Q�H��+N.ٺ$��4^��Lȳ��
V�`#g�Y�m�`�[�F�mb�u)Ю�F�NE�5țc�ɐG�������9H|bEO�$+�]1�DڠG�0�z���6R��&�'��'�
#n�;v�=[� J,o:@E%#Fe�OҢ=�')���n�8)2��@�slB�vAW&	<T�� Y}FϤ+ƲI᳎�$�H�E$�)�HO%�������A*5b��i�"O&�Y%Ү*�(0)Ⱥfq�Ҥ"O=�����śfh|UR�"Op R'aQ�+?X��nCnd#�"O� �7/��Os����P�b0�y!"O����
�������B�pE�W"O ���J�?Fpp#IB��t4��"O*�YRDHU��0�R�A�{��tX�"O�a���>i�ĻTH؋�����"O� �MR��(���i�/�)�ŨW"OP�W+�k�j�Hd/�/Jа"O���.��;dUt��BXܙ�e"O����猹a�-0f�Ϸ:XX9{D"Ojtkq�,NV��e�T,X�"�"OV���H�bP�Q�Wv��d"Oh�gI!#�T��Z�E/�9�&"O���$[4m�b<�"�@t(��"O��Y���K_�逧mĩk|�02W"OB�aa �����M�)iah黃"O�܈uaB�Tx�,�dp(�F"Ot<1A��u:@�3a�%2^�`I&"O4aQ�&�=k6l|A�����1�d"O����cQ��h��\���q"O��h���3qr ���X�h �#"O�yˡʜ6B�(-��ʵ~�<Iw"OpS��T"Q�%�\�.��Q"O��ZLV�����K�OT��c"O�}�ij�x�F�7w>���"O �a�c��E�m�mS$rLP�z�"O���(���C�b����"O@0��iH�o��![�L�W�(��"O9C'�Ư.$���c��ƌ=y�"O4�2#��/��q�7�
c|=R�"O&	rtkܣV^:)2 B�� W�E"O�h -Ða�"�q�!�=\Ni�a"OfM
���dd<lx��A�rY0�P"O\�w揉Kf>�:�͇����aV"O�X��-�:��-���X�7"O���D�m���0o�E��آ�"O"�ioEݬUx!�Ӎp��$�3"O�d�&N�Vqp��FW��I�"OD�Z��ϱ�|�fΝ��\���"O��q�-���H:�g�[��4�e"O���E�� !��ť��W�R@q"O =IIU�M�>�Y�%�_[�!S"O<h#@�ɜ~���anB�!Z���"OHP�#\E��$�D�P�ȍ"1"O��h��[�Z���ѩ7����W"O�s "�A�2�1�f֠Xy0]�	�'��z/�C�ʨb��:��qs�'c���Bc_�V��j�/ȁI˴���'s���#	��%�0C�'��D���R�'����bҒe���%A^!3�'m<��wH�	/�0@+ �����'�z����V2K������ٮ�`DR
�'��T����6�0�Q�C.U܍��'�*V/�*"��M���ق�ډq�'Rڅ17k� 3�L�#I� 9�U
�';��I@A�>x-nXc�.?��X"�'����T��]-����d�C�ҁ�
�'�B�T㛵�z������,(
�'�����mв-�j�������',~��@�L^��h�
��Xk�'�J�RPi4O�|� �81��1�'��)��jըW�4p#��Z<�%i�O�<��Έ�p��y���0��p��H�<�t���n���2�H�<�|p8��E�<�6��&�xb1`I�"8�%�^�<)�E�M*z2�mɯy���+�NFY�<	�
M�M�:��T��-l_��3�I�R�<��,�d�P���~|�<�BFPH�<IR�Z�x��k7*�6v�����@�<�-ѬU��BЇ�	_<6i�Ճ�r�<� @�ra��e�p��ȯ6����"O��$�]��|E��@Q�?.r���"O���<0�RŇD@ =�"O�a�6NQ�)���2�f�(�"Oĵ��!W�H�@���>p��p�"Oxi��(�
D�><��i-\k�M�g"O�\x7��l���q��!4(�X�"Of��ENm�-a�D)r.֙��"O�he ��yt	�v�؏��0�"O����+}T ���2]
t �1"O�@�WGv&�S���Sm
�g"O~�����N��;��͋Ll@��@"OH�4�٬�zI�7�[�H�t)�q"Ox�H7��HB���З�}��"O9H�+��c	��L��< "Ob-�TD�6�j��e2r��"O�E� ")uQ���ʾQ�,�@"O\Њ���0,��I�1'�0Q�~�S�"O&�2@���`/�E�0�R��6	��"O�@�vk-mT�iv�X�
\ DJ"O���ʸ�X�k6��l�
Ԡ�"O�T�S.I36A�afj��X�6�u"O�W��'�>������&�h�:F"Ol��a H�\X�(�!�"O&�1��=&�X��o�p���r"O|��Q����y�.J�Wn<�F"OHx`f���9�I0���K�����"O�(��ֳ&J"�dbU*
�"O��H���X2��aH3'v^<z�"O����璌[���q�پa���"O��K6��$8��ɑ!�G�=R
��"O�|�c�ұ}K�( a��
o���c�"Oĸ�2kN�3^���%��96���80"O�ĺ��( ��0C�c��\*�"O��#��?C:^�;���o���:"OZ��ɟS�(�kd�ſw&:9"O�$��`I��1:ף
���1�E"O
�1'��:/f@�FcX-n��X"O�-�c�:'����F�]'S���s�"O0�C4:(1�"Ɔ��"O�]�b���l�y�!r+hЛ�"O�H:-�	D��sF!	�S��Y�"O��`#��p���jZ>B}d�"O���3��&:pɃ���;e��#"On5��1ka\l�b���YZĄ��"O\h�cd9'�4(���CC1�E"O ���!X�
�Фi�wE4�9C"O��a�9!����V�'�8�"OL(c��_Yx�y.��9o�ؑ�"O��qmBN�����E2~A#�"O�A����[%��|��,D�DX5$���C�*%�
,D��#我O�@�:�N
4}��X5H&D�$#����,{vY94+�n��)�3`"D�|rp��Jl��#�V�6���t�"D��I���`�S9;�Y�7�/D��pt'ß,���E�U"ܛ2�!D����c�):���.]kW�-D��2"�O����� (��a�*D�d�QCU/@����j wD��(D�(�ƣ�[� �
�CB'a2S��4D�lZ#.D(Y�Θ�g�Κ�$��2D� 20�M�&����V��sXX|"�),D��qA�%V$�iA�ꘚJw5D�� ���2�0�`a@r�iG~a�"O�D0���l��a���<$���@"O��!I��xG$Kpa�|���"O�1����a�,� 7A D��P	�"O��+�@E� �0 ��_���""O�	���3t�H���)�^���"O��`�@�9]v1YA��,*HY$"O����h�*�Jy��3)�!�"Oҹ�v$�9Q)���] �)��"O,�9� �+ ��8��'8� �"O޴kVoB�5{8�Рa
*e��s"O�iɃ!��GVn����֢#�!R"O��(��I���}�'ڊI�lA��"OhPXr1�V82c�!ug��"O���)6c�DF�"a�iC�"O�ȉb/G�n�\�0�f���[`"O^1 "^�e�m�p( w��I"O l+V��&(�t�����9��	��"O�e�e��9�6�c/Y.���	"O�3��4<r& x!eԩ`�2�"O �"��e��PU��%u���8P"O֬w陯U.
�B(�7/��u�"O�̛V�K�-|� q�x�6"O\���_�D)��1��"Ov�ԂΊz��dq i��,T�H*u"O��y�f�x���Uƕ5kkf@[q"O
��$�MF���@F	7N�~}�"Orp�1@��xŤϒIེ2"O\ �m��G��`�I�2o�!"Olѩ�dZ CU9?}D��`"O���r�_/K~@��lҗB�i�c"O(�ӣ�J,*���A���	dT8ۀ"O~���
�[�4��T�NM� �d"O\����UXI�bP{A���"O����k����5$U5�T��W"O��a�L�C��U��[><.���"O�����gDZ���L�%'����"ON`����1Ġ��+��&$ЀP"O|�3�o���(^��|��;�y��:F��d�J���U���(�yr�I�����k^!6���Z�m���y�b\2���P	
f���j�Œ��y��4��0R��Ĺ
��A�t���yR�CQ��K��^Lh����y��	)<%�ɹ�ង ��l��̏<�y2�N�X���2���5X `z�"���y�C�2
Nɰ0G��++XiP���1�yRHE�>��T٥�1(���kS���yREM�A	�ȣ���]*8(8c���yR��.1��d�4R�H�y����8Œa�=M
dӵ�s�!�dC;;�U�A�/�`Q���/a�!��1� ��ƪC*+�� 2��!�䇲���T�Եuݸ��s�2�!��L^0�l+��߆Y�"(�h�*�!��,*��e�2 �:^�x�# Ꚕ�!�D�Av�J��W�8� ��P��!�>d��Q' ��p�4l�@k�'56!�N�{;�y4�D>��9'+V�#�ɳidr���"�)y�:�#ƭ=5^"=�4+��mE����O `p���T�<�%MwQ�WO��ɋ���Q�<1�_�j'&[7�d��O�<���:t�PG��U7��#$b�N�<A� hA�xaЯM�S�J�z�&Rc�<� 8q�/�Sf�q���Ȩ;�½B"O����ٻc�(`�p��<z�5"O��h��.��՚�iz���2"O6E�P%T�v��S�g�z-�mғ"O:�K�I-I9�Q8q���j<��"O�xcBA���"�po�aB$"O��2��]� #�T�?c���T"OF�t�U�7�Ű�d)DCtI�%"O�H�� �Xt�3FBx>6��"O*�8WfY.m�� x�D��}:����"O��e�[�\��J�e�9
$pԋ�"Od�fθ\<�˦�(e&�g"Oz	Y��D�F���_Dh2�"O$H���c�L4rF����B��!"O��p��ғ|��|I�i��r�J��v"Ol �q�O-b��4��H^?Wl@H��"O� !�h�JZ�С�E`�`"O\�q�ׅy���1#�q	�d0�y�+�Z�Hr���!�z�sG�/�yRMѥ!7򥚓KD(NPQ:�`
�yr���:�%�A�U�.TR�S��y�L�<� �����E��(fb�yB�7T��[�Gr�����ɉ�y��B�;�����-��n3ɣ�k��y��B�K� ��Z�T��"!����y�ډtN������3H���%n�-�yB�K b�$`IV��$D
�P�vo�5�y�(	�1�r��HǼCØ�&��2�y��S;��l�T��q�:��U���yr�8<;vq2�ᐚkO�@��W��y�� P�H��7i�eh�p�M��y"�̐�y�hïs�f��5D��yR#+K<];u	��.�2PR�y򁍾�@H�TZ�Q����)�yҢU2�P	b����TXRT1�➅�y2nIR�b�@(�xJ���հ�y�N�t�B[�mF�ALB�b����y��GC�A!!�;4�I�v�^��y�Cʯn�.��p�2�>�Kv�O��y���lZ A�,я<�`�5���y�câS6�:�E�7q���G�0�y�kt5`��H3*�
������y�f�f��#�+6L[� @�Y��ybڂg�P��J�A�&DP���y�L	r��ш&����*a��y�O�I�Pt�`lO�6�b���y�A� �A!��I&��0*��y��B���:īX.I��L�'����y��I
te���B������@�y��1�lyȐN��:A�)ҷ�ú�y�/»5�RE�afO�3�`�����y�.C*J%�$��c�ĭ�Ќ���y���U��i[Ԃ�^���gi9�y�	�^8����$T��K�H�y�ÀCȖ��w �Na��Ab���yRd�!F�ܲvE�Tn*�
2W��y"��w,��� �B�K�B��AQ�<	�ᘷ	�(��,X�i��Z@�KN�<�����m�t喇 !��A�cP�<(  ���uf]�k�0$A7��I�<�R�7^4�I��C<d�3` ~�<Y�d0;���s�@�����Ԍz�< �G�]��pEׅ4�\R�#Zv�<I�@���*�?`|���J�y�<� :@a&���h5���'ckEB�"OD���0fvn{v�\cj��s"O�-WA�N	m`�^�W<ڱ�"O�Ebc�Qn& ���ZKx Z"O�a	!����R��V��ZUx��"O�t���O���`rC g�q�A"O���i��|�ܹآ%]�]z��ʤ"O�� ȁ1x����%I6��q�"Of��9��x�D�kP�L�"O޽BgA3p+i�C�=Q(#"O��U"m�T�C�S1@��e"O8x�!�1,���{� 	4I�J� �"O\���D K4UK���V�D��"O�4���V���L��<����"O\���]�Z���S�

J "O6i�� D�C�G�7�H��V"Oȵ�N��0L��+�+4���3�"O t*
�0��S�	Fnq�ͪ�"O�%�dc�+qXՉ&&Q�'R�!`�"OZ��jS�#%r�1�%@#Ռ��Q"Oܰ���o���`e�M�$jjE9�"O:�`���uD0��J	)W^���"O�x�&�Fi�`���
���"O$ܘ�&ܫ;���箎"����"O��xfg��!�i
� X#�̔��"O�p�Պ�&Kk�����+"��т0"Ol����!m�T� l �9)��@"O0m*`k��8*�ik���
�	��"OP�Q�Ƙ!��3C�� U.����"O4��ɑ���|֡��{��z�"O�u�gj\�bp^iCG7(PJP"O	s��!� 0� 
bћ"O��ܪ����o�X��M4"O~(����iz6�3��X�a�<@! "O,�Z�͍�a��,@�� H�\9�"On��2�["���*���ެ9��"O8�	5ɞ,#�b٫���[ܔ8hp"O�e[&#ˎO2�ph&��4vѾ�j"O�02��Ѳ[��B�����"O�Q��D0scPL0�H�K
���=Q�y� V�3�lM��i�- �(����y�	�E�`���ۙP?�`������'7ў�V�@'��8<� -�7hB	`�ˣ*O\��e�ݴ#�F�I��u@źd�I��H��ɽb�`�6`�)H��1�5�ŭ _�C�8:.�hA�X�KD�Q�O�u���0���~��7C>jd�'*��e}�a� ���p=�m�A�I\k<|��E��n�q�(�B�IF��7!�$t;Hqpj_T�������5oz&E�$�Z;u��R���'GR9ADN��y��$E���*\�l�X���%̖]I��$�)��<1��J��6#ؙ@+�y�. N�<��._^6�Z��wA�1+tjLy�mш�p>r�;p?��ѩ�?�\���HBG����ux�Ϻi�~Dp���C�i�񮙙3!��L)�ΐ*`�;lθ0Xf�Ȕ.�Of�=��"����Y��� A���� p2"O^��B+A�9�T���S�޹:�*O,x�D��=Rb�HR$وA�Fq�	�'0��,��TN�%�q"66|�0�' @8d@ݐ��[�$�-���'ff�KA�IH��h�/(a8Ī�'��\�kB��ѪCh�;!� | �'#����f�0G�!�#�,`JD#��� �D�+@�o�~-�@eY�I���#�"O^��5#T1=�	0u!ܜ[�n�x"On8�Ce�&�֠J�晳rT��S"O��Zb%�,���G��"��(�4"O��0�$_6#�z��.�\�Xt"O6� C ����P�2�,�e"O:`)���F?�ɺ��ߢ:�$u�"O`e!�PPx�<��,��u���"O��4�
o�� %fȶ#�0�X"O�UQև�v��a�۩-C��h�"O&��A�T�n��=9dcųS��	a"O�T׋�I��B��h�2�c�"O�(	E�I�cz�X�!*~�����"O����ŷH�Ա# J�k��@��"OڈB"K\	M�L�xR�_�F��t"O�४:�j���E��3�L�6"O����e�,p<�����~��A�"O��F��6	Qވ:�ĉh�q�"O&��h�|����G-}^���e"O,��T�9UY4�+�0w�DD�a"O���u͏� `Z�2�nI�m��$Q�"O�R0��)f�pWd��a��x�"O�׭f�F��DJ)=n��F"O��8%OV�G� ��b�Ljh]�Q"OP�Z$aa���*RO�%Sb�s�"O �b��Y7mΨ�A��4t��JU"O:[E��T↜��ߝ���"O ���mގ&4*a�w'C_n�I�F"OHH�ȕ8">U�Ӱ:|Ĳ"Ot���k- th��D�L�	��"Oz��e��D��28P�`�"O����j���(��uM�\+��Ʉ"O�  �5������X'@@0��"O: �6�"m�~!�' ��$<4�Jw"Ohd��O??)�xv���^�nM��"O(ԻS�$��0� �'q����"O�QA��H�2��p�F�9�&��3"O)2�kȩ L�8"�GN����"O�U��$�@s�J�_���	�"O$-��.8#��I	�+F˚u�w"O@�(�m� ��D��f�` Z%"O MP���+v�QE�ǏC��L�"O�uY1O��$�`����#��UJ�"OH4KGAD�	|JĚ�eH�,� �D"O^8��#�0@�5�aQ-~�Ęp"O���(#KD��B@�o��M�"ODQ�V@Ɏ@]�a���
`O���y��)$҈�r��c�-:1�F8�y�"�-ج�REĔ�0���"C��yro�����@axa�l��i]�y��*	�p�h]�p� �:�y�^�$��G�:\�QQՍ��y�%�3W����R04X5c���y���+�XtyAf�(^6hu�E��yB��"��p�A�'�t�1�+;�y�W)s���i��J&�d@����y���04���R��O�F�$�����y�N̎g��a��ŝD��y
�j*�yB@�/�xن,W�2�J�0��4�y��S.:�d�`��Lt�|�P�Å!�yB��7gs0���̆��Q�S�\��'d��6A�D���d�ɰ<�Nx`�'���3�+ZO⨔�7��3�\� �'^�Ԋ @ ��      Ĵ���	��ZL�v�:P���dC}"�ײK*<ac�ʄ��iZ�Fm��x�o�
�6�ٳ�PhS��͋O���B�K�AL��(�=8�0lZ��M��#��Y=2���+���I��L��FU�o��x�ɝ2L<�F@0`R1�Z�Xy��B����QM�آ��I/�8��*�A���gY���bFޢ+��LE����L�[5�	��mYd
L4��I�r���`"'t�(�R�L�*>���֌�P}&��6.ӜN�&>;t���n��_(�8� G'N"jE�}�ā�=,L�D��M��α;D���B�O�xHk�;� ��҆	0����Ozѐ�nC�0O
x"i^!$��<ȻBe8�*8� A	�b�k#��I>�6(�8}s��%��GH�#[aq�V����2(�� ϠhW4��',�d%zq�X��F.�OALx�qP��~
�`�]H ��U��#/a�I�QE�՟@w-[�r%�=�J����Ɏ����I��y��ߢ/'1�c�.m<8��V)
[>	��c�D�		d7�LH"1�$�� W�xҐ�i����G�I���7zr:�i�4�~�,~s�4����	�Q.ؐ�J��z�ə�Ob :m&T~�񕋘��t�x�g�����+"�d�j��}�s��x���H3ǟ�c�.!�����gz|�r��G�v���� ��� ��)֬�;CL��)��T;�W��'�EW��O^-�a�O�'v6�	dB�Y�* �$��{�����	�[ij6�u��8�%$H��+X?Q�5O4��èC\� ݂���O����v�r� u�-��Y��ύ�W�,Da ��R�ɺ�[?��,ݒp���;��:�l���m�6_��K� �-&�U�'����e.#�$Ū[����xR���1�T 'Iе�J��ū�`���d���0#~XB FU��h�"R�y��z��[7A|�Iu�8�y���m d  � d  � �O��xw�ɳA�0����]����"Ofu�V��@�8�N�1�V4�"O:a�+øH�:ݨ���R����"O�1DŒa���xH_�#J���"O�4���ߥڰi��\%d>���"O0�i4抱I��0봆�bҌ��F"O��I�j��hf\�Ē Ϙ�2�"O�|��bӈH!XW���A��\�E"O�2�)R�j��q2���#��`�E"O�uaP��5*�"RJ��d0�"O��Kƣܵ�}�޸;T,��Q"O�a �8��L��oW>�!�C"O��Y�f��A�(�:O�~�>��"O�9j��ΑA�<��1��h9�`"O�tx�D�j��AK'��9p�,�k"OXU1��đ]0"`0b��'���"�"O��ӢŞ`�����[�hxq�"O�m��&B�'R ]�6[Ĝ@�"O�"�c=��
��f��k"O>�2qM�!7/��a6@F�\
l�C"O��MN�ڨ!f�:S�Ȕ�"O��3�ʄ�^��yR�b�']�����"Ozh�Q�/W�|��!�+i�l��""OX��S��;ET��3%&�VL��"O������K#b��	ͨ]��"O��2��șD�@�J�'��5�8��"OLɈ��U8!�\X!�ES8����"O�4�Ao�mjx���� 3#|>8�"O̼`�׮5wD³�ͰO{E��"O�:����o�:��c��i�K�"O`k�G]viJ)H&��T�vMI�"O=S���(P�0�"��+�|�B"O`� eաm��;��
6>�]�"O蝙B�
�����T�k�:��"OH�)��O%����	[v����"O�dI�*W�u�� �BHGX\Q)G"O�:B�V8>:n����X态��"OTaIQ"�b�ty�X)&�%�G"O�рC���R�P� E�,l��!"O\D�%(�Y*	�cC�vV��p"O��H�,��}�Ǣ^�M2	�`"O8-�Q�V,���P�_�<���T"O�e�f�Ɏu��EZ#Cz)x<�"O����I�G˨E��M-��"O2ӓ�I"�2�JP�%����"O�)ɣ�<Ў@��Ӥx����"OĹ���[�N��1���^=��Hx "O�88#i��B���g�r���kg"O ���/1�\� F]����q"O8-�ma�.-#����^pz'"O<Eit��)9�*�R5�� v����"O-��B�E-���!�9=W�dx%"O��2��sB"�*�`:vL4���"O�1C��X?+�2$��NM�h�PH V"O� .��Ą��GGĹ��m� ���"Or\)7���K%h���*	"�޵�!"Od��lY�{�~�B��՟t�B�;r"Oܹ��G� V�0�UȂ�Px1c�"Of�����	L�֌K��M)M��і"O�!* �L7 ,*�8	ȺѫAM6D����J	ՠ�ʔ�׵8ܑ�qb)D����Ly� !���dhby���%D�(K@
Z!*G����8e��T�=D��v閖
�0%]!Mi�t�D�'D�X���8[3��K�ah|� %%D��r�˕9}�z��d�T?HT�׊%D�lqf��c���+��D�L��k1D�ĲE([X�N �OȜP�P1�J$D�aFꃊ]�Б*v�E%?��Re�"D�hE��	[�z�¢x�ňӋ"D�<
 �K�|��|kw���(J�i!D��y�h$�Q*�`J��&�$D�Th��I�
�mj�H�t5�6�#D��b�N�D�r�jgW=BGX�;g/D�P��U�qN�Yq����ZD<�!u�(D�l*���Z��Ab�hP ��2�&D�4Q2l��q��M0GEm8�1�R�$D�@��#�0ф�Y�¸Kj����"&D�p�˅3�Vt� ʞ9J�A��?D���@P�Fj��QE�+P�&$�� >D��#�R:+2��i�真!�.�[�i<D�@���:9�|�e�[4]kJ�[ti<D������0H�;�H�2I����B(D�x�1�=Z3�4eb�F6��Pp))D���!�y��p5B07c�T`3C'D��i�+	<e��	��
T�Bk�@��?D�8C�-�=Z�����W�G�8]t�>D���V�#����勾_���">D��� (1 ��lq&k�(yԜ8$O(D���Q�#�Π�$f�5r~�{�3D��+�(1��
2�	�
Z�[�+0D���S�[F.�J&+r�T@q�.D��KЎY�
�d�W�aO��K'�!D���w&vn�	G�W	:���iWE?D��a��uzj��O��z:�ܓ2L<D�lC��B�n��d�f�1V`�ʃ <D��re �+Mf�����S�髴�%D��[ ���P 2�S#H|��ɱ�6D�3��]7.��Cp��Rs��yb�ׇB��]+���W� x�B)�-�y�� �� �#��-��N��y�lɢX�<iCF 4����M"�y���K���ؓOӨj��p����ybH͙n��;�#h&H���ǁ�ybhA�P��4Iɂ1�"��PD+�y�J�0n� 1sԤұ�lDc�M@��y��&#�ޥ5��%��p'�C��y����6�~�em�������&��y��	V�b]xv)��AqU ��yb�Է?l:8�&�v6�4�	�y�EU�"�~�xb*�S�*,� ���y����m���Jc6�y��D��y�����"3"�;�B8�l�/�y�ƑYt�����O~A�xs�D��y�AޏExV��P����`���ػ�y�FM�T�VE�tI�P"���yR���������wP�=�v-خ�yR%�T(DQ�"N4Em 8&mч�y
� ����!��J�H���R,����"O�]�P	�E���s�G a?հ"O���H�7HA���(/<��Y��"O|�)M4H���q�
�W�6YR"O�3!o�)K"��Z�[�Z��<0�"Or���4*������"O�����P.� @�l��[s"OdH�GbL�\+��tn��&_��"OF�s3�� #\���.^'xQLh�"O��B̑*:�e����>I&m[%"O�ȑ�`�������q�D"OZ� �VTYF�H�T����2"OD��W��3�n ���	=t9>�"Of����A�c� ��S���D�W"O�uk���r�C�>� Z!"O
��fn �=9�M'�-�\A�"O���c�VA�L)>xY�"Oa�g��~ȡX�BK�V�칸q"Oҽr&�/nߞ\"2!JQ�e�"Or}�S�2N�x��/B�x{�"O`�:pHY>
8��
5�ڌo�H��%"O��+'Z�i)QK�
�0�Ӆ"O�l�pl����ِ�/
��䱓�"O tA��Z0�$���B�B`��j'"O���� Ţ&ШC���jP��"Of��o���н�C��(|�	�"O"ѣ��1<����ʇVl����"O�D����x�i�n��S8�1:�"O������N�M���J��|�e"O��BK
�U�g�x�԰@"O���C�Zʘ��Qi�+1[�L��"O���G,>8����獭g82�"O�ɸS-�4N��sf�ʲ�v�� "OT�*b��ywE������"O���ꋿ?C�8f*I |ԁ��"OH�����5[/&���N�In�3�"O����gh�3�aڸrU`�Qe"O�AB���wS��z�ω�[<l���"O|�т̟#(�,
'��"�<�6"OаZ��O!�H�h�픋hbֹy�"OL|�J�hnt��-|INa��"O���'=R��y�Mπ1=,�z�"O(ESG�-��/~#���"Op�p��5<���5�O�jtkQ"O\�ӣ/M�|bR���� �"Oz�3J8I!i%	�s��|Ð"O ʄ喋b���(i���T���"O$��,T�z������la�r�"O�q�s�&7fp��b��I`v�"O���O�S!���]3RHTAB"O�5s���m��s�`¯1��w"O�`;�^�Ux�@��7k�4x&"O6(b�+6.�� �&�99�@`��"OF<90:�~I�#�1t\02"Oޔ� ��p�*�ȥ�� Y���"O�[@ڿ;K����� d�+#"O� �B��I�Y�gwO�h�"OD�s.̵l�"�0q'A97D��:�"O��� ��"�P%i��)��E�"O�b���o�6�xP��b�ؙ�"O�H+1�Ƙ�����ǯX���+�"Ob�I�%�,d�饥�J�j � "O�����o��)ф�)]���"O�L��Nh�I��RT�I��5�y
� ��:�ً)>*���H��"O�yQH%/h�Y�!aә�
�)�"OZA�p�� �t) ���1P6����"O�=����}�V8�.�="�)�a"Oh��c	!�J�3��1: !��"O�):�L�&������
����"O��N#���y�'U��z�"O���ꗬ'D<�s��8���d"O��
�͕,Ae\�b򨁩4�ś�"O6�i��8"8ؘs�T�x�(D��"O�a�<M٢RE'Hrp$`�"O�Sf��7I�	��&F�%GtP!�"OX��Ǣ8Ci| ��P-3�|!"OB�a� ��RK@`:�Κ�K2N��7"O�%h0-��,hb�lR���0"OR�K����b�(ٹv,êi���3"O����LH�*A��Ҙ��"O*9�wOY$#�A�A�ݫj��8G"O$�ٳ�)1��eEM�4�0�b"O
��nG�gr.���91^�(�"OX���G����ID���"O�Z�K:+�-�ah�'N���v"O�Ig����$�IK&M���*a"O �b׻˒��b�g�B��b�<�a
ڤX�D�����	`�N`s�iK^�<	�J؛\mp�نȈ@��e�<&��%/,�A!֭�#8|c@k�<��h��)H �P��2�h�<�cg���u9��%`��Xw�a�<��MI� Z���!�ǡ3.���FZ\�<1R�Ҿǜ��Fm�P��Q!�l�<�% (p˶P*�i/�q�p�Pm�<�R�@�O>~)��̆+3��b��^�<1��l8��s,M-����'@�<ѕ'�m_H0��+6=2��Ł�q�<a���j�l2hQ&mo�eA hMp�<YBmY��Iy�b�"W<	1�Ru�<Y�)��E%����3&]r���+�j�<��LB�̌AI�=�\ �K[l�<�c*���#1��>�)��e�<�g�*�a[VKS�Bh<�����`�<ٲ�`���(Aɜ	�DL`�<����	?��(�T4����@)t!��ʜ,��O� ��x(ӀV.�!�Ė-� �S�LZ�|�>Yyq $<�!�D֙;�����A�F��7J�s�!�68��`ԉ�:'����4��*�!�P,Z�"0D�ob���Ԃ�+${!�$/U~�`�0N��YV�q�̗({!�Ѻ}�$�.݄[��LS��{e!��A�=��X��!��4)�	_�W�!��܀E�����M�I,���h�:0�!��\�2@*��j ��g�k�!�D	:Y��DU)������!�؃!���&��aWR}#�R)�!�I�fw�]��fI!0芥"DmA�D�!�dٺά�Y����Kg"˵V!��Z3Kv%�b��}�
p�2KM� 9!�$
(;xB`�����0��="!�@�4�h��%��"rhac��"z�!�d��}w�ma���0n�	{�F��!�$-a�t�
&'�lZ\ 2(�!��D��ԍ��R!w������<7�!�D�<��Y d(ۛ�D�@����!�� ��gG��V鞸1��<*����"O�8��GG=�ʑ0wA��Y\�Y"OR�2o��v��a;#��.I�R�`"OH99'1��-��V9P�Nhh"O(��C��ziZ|r�����R"OF��C���T�xT+a*'�>1�"O>���B͘%�Z��Q�E	��hu"Oj���D.PW����؇W�~��G"O�D၏�&�� #��{���'"O�i��p��y#����7aV""Ob1q��Q��������~I�"OR	���_oCu�@� �.9�"OD���4,���4�����Y�yRϜ:O��X�A�i� xe��e�<)�U�r�����G�3ν)�]v�<�Ѥ@�+(���a�~�0���W�<����u@`,j�^9�8͇ȓL�P@�B�L�p!hB��+L�	���.�����X���5B�D���ȓd�A�DDoN��1�R�/����ȓ#f�(" ����q�/H�7��ȓ��R%)DW�,D��*�4��Ն��"�(O�`],�P'R�8�t��ȓ$�FA8��&22L���m�{�����Lۢ�Ҧ,^ZNx����&/��F�Z Z���N�m`#��W�2d��s�(}�g��+zCLh8��k2XQ�����&F�:X����fEuN0�ȓ+�̹c_6Sn$�����5de�U�ȓ= J��D�~����O�/y��ȓcTX0GǞb̤��e�04	P��ȓ'���Q��W�`u�&�<yՆ����0AR�07����ߴ
����ȓb�,�����0V���4F�d��\T�Da��|��T��٬N�I��N����J |2��J�D��\��o0�-��Eз �<�񲦉Q ���ȓ@%`-9r��6e��ѠL+ l͇�y,ā��"?��� I�/-2y��F�~�Q�J͔��`�h��Նȓ�������7D���!AV$��ȓXCRĈ	Y���p�҉f� 9�ȓ(��I�1E�`�@�J��W)��o.fQq�'�qH$�r��E�֙����y"���/I:�2�h�<Gp�ȓ��,�$C�b{b5� hX�@E썅�#��=��$X� D��"-�&I=>��ȓ/�� !�Ů7|ꀓ@D��~����t4%@� )M��%S�|=��
�&��ѠA���VO�2nي0���6ljHC�-q�14 ��H�Ʌ�P𶬩��˲G%�xa�N�g�!����p�D�Em8 ��ӕ@���ȓm.�9a�X�}�@e
�;^"���UL��VKK�\�n�c��es-��,��|	���ߘM��		%R%�ȓ{Vz4[�+ƭ_�>ى����uv��ȓ�.�p �
4
ZTX)�gP�ao��ȓq�֨��|�x�o���e��(�I`�,
�*�Ř�M��.e�!�ȓxNLIQ�(�m$�`����}���aY��B-Glh1� *�_�Nԇȓ.�N�3B�ݠ*�:�q�˚_������Я,9Zl@��Zy8��[�"O� ��u��-`2!A��y4NE�g"Ob@���<�<0�J�zE�9Z�"O��{���W�`�V��P(P+�"O�I�@E�1�9B$�`#�A�Q"O��˵�fk���'\�0j�I�"O~�)��߬X*�(X2�C�n�Z��"O��жn].��jW�X��t�P�"O��:n�O���[�>tFE�B"OJ���\��V<S �F�{f�l7"On�*V���{�lsA
�X=Av"Oh����Vߦk2爻|��I(p"Oh�#�7G~���%�4wr s"O��� ��*:�8]�&jy�䂁"OV��f��9�0�-gfnu��"O� �nN'B���svk�rg���d"Ox<�5�E	4{HarlA'k
�)B"OV��`���&���JE0U�pa@"O���#s��UI"���S��"OʐCU#)B<@
B��G�QK"OHU�2b[����� �(9�Q�A"OTP)s�S:[@ʈ�� -xH�"O�Hj���$����*�G�l�1"O�T���$"�`s�FY5��,��"OjEeh]����Е�̬�6"O ����
�4�hl�E��trv�Q�"O�l���&O��j*�.`mey�"O��Q.��{;��H�~���a"Or4"��ю_FT�u��?~sl��"OXX;��I�0�n`�4�\�i>��F"O85�F1��%ۜI��P�"OB@J�zb�녃EE *Y�"O�q����P�ޘ� mף;�B!��"O(���9V'R��ʜEj��p"O��T�1V���Z7_�n��"O@��[� ���2HQ-'� ��"Op5�p��9g;&���Ч�0;�"O���bhG�Ό�.�J�� "O(C�K��N�����x"�jU"O.�!4fK> �b6!E:%m����"O�9��3y�:8
�=Cp��3"O��	��Nn����-b$�Y�"O��zu)!8��uxѦm���A%"Opcd�T/aM�	����,{ �1 �"O��QC�KY����j���a$"O��e�S��H�"!�8�h�"O1�F�%�F������� "O���c�ݩT�X�4�ղCn�h��"O���v�$j���5Gߎth@T)V"O��C hF�=ΔXZU��:Ȥ��"O� �+�cv
ԛDd��l�N1�W"O��C�k��S����Ec�L��\��"O�Ԓ��V�e��$ ��<4��\��"O||3��7fJ#%��7�H��"O���%�Wg�)��CM�- ��u"O�d��ǉ�`�&1A�!']-H�W"O��!��!e�(���`��@� "O���A#%~;��#"A�g�8��"O�@GlG�IH��(vnS{�^�"OY����2c�ְ���w��3�"O�壤�V��Fa���?M��<0"O�h��\4��c `�;AnXi�"O��9�j���8K��L�>�ܓ�"OX�"X0�j�Y�흭_.J��s"OlE���
'
�I5l�S/��4"O� ���̆9>��jY�)���31"O L�#H�&��Q1)ǭr�#"O�!�"�41,�U;�g�?xdRr%"O����'(C�1�&=��z""O�U�s匤ݠH�Cf_g�x�2"O��x͍%.dı����ݼ$3$"O��q� ��)m`XZ��Oښ�4"O"���*��0��5*�.ĳ�"O�u�&@���(B?%�Լ�@"OD�Qk��f���V�
��q"O^l��%�-D5"Sf҆��A�S"OR]��2uDfe	bWB�h�"O\���쀚J=�XkŦJ\s4�
�"O¹Q�B�	"����<���U"O���K�ten�R���LF�x��"O��y7A^(
�<�R$�"ٚ��`"Oȼ�d.4>.4�JDD���P��q"O�`�LU	o"XJ��~���a�"OH)�!^�G6�äd�!'n��@"O���� �:x;f�wsΡ(3"Oθp���F��� � �vUV��"O�![��?�(mz�b��O@
иv"O��GCݎ(�I�A�(�q�"O<�t*8V��q�� �`(D1�"O��*��Q�u���!U��y�Ř"O��
���U-R4 ���:�n�)�"O��w��� ����×,D�\�g"O�ͳf�I,eA���+�*2��{a"O�}H�*� "��Yf��x?�tv"O�����=4��Y��!1Y��"O�l8C�ׅG����ԩq��Eb"ONM�m�l���j
�s>��*r"OJx�#�^�� ��b��$hA"O2Q��	R z�2Ș�ȗ�~��1��"OƑ�3,^ta��5G�-wl���W"OX!���Ҏ~.��X��ײ8�A�1"O͑'��T{.䂗_*t���`U"OFYЁɅ�0��۶@"�&T��"O���43Z$��#�V�vY��"O���T�B�_Fq��r}�i�"O�m��ܦ�*WP
^B���"O����B,=M�8���^&��"On�`�G�U"����sJ$Yu"O�!�)��U�+�2V����#�\�<�e�'9}�թ �]8bM&����Dc�<a�N�]Ht�����/r��i��@H�<��D��<��\!Հ�"�F�貀@�<y`�R:q�}
��>$'ڤ�.�x�<Y3�şjR8{�iӹcb`2v�<��.��_� t�a�rtB�a��t�<�3	Q�9j�pS�$E�->����n�<�C�ƅb���Q�Y�{����"A�R�<Y�,D6c���8�)L9Q��xs(�C�<�r�+2���CӇ��Je.$K�̉d�<A�'�]�vi���4b�p�3�v�<��3Ln�#��܅%���K��o�<Q�K� gm$�u(�&bJ����k�<9�+V U���`TM�<'�xe��ʓs�<IfP�m����f�;d�"�{Um�<Q�
�.U)ƉY�!5"�9�L�e�<c�ߎm����u�J�RTÑAX\�<�6��G� �p�W?:�nt��e�r�<9�K?V�����G:co�H�*Sp�<�c� >���t�1��MQk�<� �U+%OȬ}���Cb���kH�"Ov-�կM�[A)g$̥(�AB�"OF�z�!�|��p�;1/jm"�"O��[s��2*�V!t�`5k �f�<ٕ!5�M
��Vi6��UKb�<!�нZu�ax���k��#�!Fr�<�w$H{��;ć�K:x���H�<ied��0���ćY�|��f$EG�<�E�BDӸ	i�'� b�Idg�F�<��%C�HKL����׋'|��9��E�<!p
�;��QJ�ȇ
!���p��\�<9v�շ�ha�eɔ/t �O[n�<�����~a	�/���kFEB�<QR.�=�(�Z!+1��I ��T�<	մ"(&%���}�scOE{�<1R�'b$�d
лR�;åu�<�q%	��&�sJ�Mwl,��dH\�<��ύ�$Xr�Q��nɲS�AY�<aP
�$A+����1.4}2s�y�<���Y�n�|�����J�n��@bM�<I��7.gT5A��J�6���tmBL�<�(�Ҁj�B :�Ȃ��R�<�"O�1"|֥8����Deֱ���W�<9f$��f�DK�g�+l������W�<ɇ���ɡ3�ʱ�����CP�<���9t�j�h �
�ּ�VODO�<�7ˉ��r��'D�<~4Y`�B�K�<y5��k! ��ZXY���\ �RԄ�B2����[���zUbE�6m�8�ȓ^T�LI�o��v���e� GH���	�!��.��퀲�
�^��:o�]����S��L�@_��D�ȓK�(z��M&&i4t�!�Fq��?$h�ae?M��a8�	9&���q�6���ᔆmR�T��
�&�Ҝ�ȓ&��<@A�٘`�֍�b��s0u�ȓP�)YRE?5R@1�W�ߔ4zp��g,N=��K�b�M�s�S6z���2��e��J�J���cI���ȓ?S�Q&߁I��xR��2N$��r�V�kVO ��"���Jg���'�Ji��>4~Z��a��7��B�Ƀq�T8�dX�Xt~��Ҙ~
RC�I�y��X��
?Apy)��܏>��C�I̰W���~�8��b#��TJB�%vɒ��QaY�j�����mN�C��ئ<�h�dܠ��kV�C�	�H,f��,��&�Af�\�<B䉆s#��c�	Yx���3�� <�C��#� U�bY�> ������*Z�C�	%`�Чi��Xހi���0u�C�	��<�H@ں'ސ���A �w��C�	�|�%T��%�4�	�˩nh�C�FV�\���*:q�#�ܻ6��C�	.q�ғ��)N5 #��'c�jC�	;/�P�&E[��0ݩd*�'B<B�	�M����WG� ���G�8B�ɩW��ٲ�K `���!���J�C�I+4z��f -;�(UQ6�ިv[�C䉍	�������P.aj��26JC��H������'EB�Zg��?�4C�	�,��qS�aԡ/���U��r��B�I�:3
5�uO	Hn<�s��L�`C�	!Q*�ȣ���[�d��G�Q�C�)� ���$�; :�X4A�U�`��'"O@�Q��%d�)"�+�5��"Oz�c��?o���1n܋S�j���"Or4����'N ��7��Y &"ODC0�+B"i9�`���Bܰ "Oؽ��Y����P��z@#"O��5$RN�P��˳Wĺus%"ON}�����#bܔ8�ȐU�:�A�"O��c�ٺG�\���_.�8 �"O��s%�Qꑳ�!��B��"O��r�0�g`H�$��I��"O�Ya�B:v���ߟ6���"Oz�u�1��3(�:K��Q�"O�*�+��A�ԃ�`�Ա2`"O�!�!Bw��M됇�Z�,�p�"OH�`ᖎ-�4����	O��"v"O����M�"(M��	a@I"O�@{u�N�����.����YR%9D��(Ʃ,���I�,�; +�M� 9D����`�7�,�0f炮%$�}��7D��!�Đ S1Jp#s� �Q���R��7D�첑��uBM����=�Td;�` D�d�j�c�e��k 6Z� `��*,D�t�Rg�?�)�(�%O���c�%D�(z��ϾnX֥��MA�+r��i��8D���$T(}����E�1g����7D�\a� G�7O4�ࢅ<5�0y�4D�[�됧���D��
����F�/D������3ob�I�W�	&s���bs�)D�(�p�Y�v��p!>rK����H=D�`���Hr����GR�^��#?D���o7w�P���
�k�>@���=D�x9�c�7�d�۶N��.��Hy�`0D��� ��)�a�G��:.Լ�`�/D�Ԋ''�
���:F���@Ȱx��*D�x{���2nT�I��gɋI�εCU�)D��y����Tz<�a�Ų1U��p�:D��uM�*<���(e��xZ�c:D���EF�f�$�S
ƫI\�ԋ`7D��ɁawN�	���Z��pyG D�t*@��Z�pxk���T;��=D��X�mDL�����C�O�T����9D�@��#�z����'��� ��-,D�p+��ʲ+���bA[�V��k�,D��0R�X��0�fNZ��li!AB(D����oG=D��M��pmN���*%D�xّF�=DH��2��49zn$D�X�sd� Rz|�Ǯ>��yi� D��Y��Z"U�T�91�P n�IA0I=D��°���6�T��p���
���!�.D��ɗ��~�]�ǵO�`͓� !D��[sOޥ2Ɍ����W�$	A?D�P�_�:V
x����)ڸ!#w*D�H�'�EϺ��B*�yh���A'D������=��=��#�T#r|���#D���ubL+	�\l�Տ[��nh���6D��RAN�.A�t0䎙!G#�4	�3D�(Bǭ�N���	�"�Tjh80D��(4H�%q�ډ� ϕ�Vf(��,D�l��AV�}�4�2+�����Jw�)D�d�����~` �Љ3��=�F)D��E��`L0�#H��z���
)D���B"��lXx�e�M��*�J�B%D��PLL�_��{�}9�l�Qg#D�� ���4mZ�K�A v]>s?T`k�"O�pqg�B�:lD0��5�꤈�"Ot��V	�[{Xh���<ƶ�p�"OR5{����1B�]�vn�-��C"O��k�j�$W�JSm�2[%�]�f"O}Q����0Ҩ�TKֆ=��"O���5$u( ��&,|R5"O8=�s��oǸq� P����"O���$���� �@,�"D�>�� "O�{v��Pt�A��G�d���*O���c��*`b �e�ESm$�c�'Y^��v��&E�W�J�J@p)��'DL �Wg<\a�"H�w��P��'zZQA��

+�e@Z�@<j�'_F�yծ3b6���C�F���'f5����z� V�55f��`qF>D����Mˈ�]r#eP�V�t��=D���Ɣ�y_x�ېE�wP&}��=D�ԐgoƸQ���3A@Jq'D�QwE0[���V�>��Jp�(D�xk�֭S�2�2�Cգ
�L- C%D�X� ʟ:9�d�ǏQ� ـ��@$D����A�2MT���9m|�#'	%D�����C�:� ��Y6�f8T*#D���ҭ�wި�Z3I�,J ��!D��%"�:fB� _�>��s��>D�XkQ)\/*����AǘiҬ�(� <D��[፿}��#`��0RdI��H5D�����5[1�1�A�6�J1JB7D�����3F.>�+�,�-�t%;�4D����.R�cl5�G��6&Y����M'D�8�v/
�sn��p�gݯ<z� �m%D�8ّ�6!7�	7����E>D���d#�I��`� ؀DQ�����;D�,+�hׂd������as�$�I;D�tk�mˮV0�� Õ�b}�5�S�#D��SNg��x��В~ל�(5	=D��*"�A�!JdfE,;h	�R�:D����&�<qz����=G8��fE:D�� 0����݁�ɗ�v^A�r�3D�,b����91���D��m���%1D�L ��|�!E����8y��.D�(�iT3a3,E�晚7Ǝ���.D�<���#A������
�e(	,D��	�h�$G��L���J7s- ����(D���a,M�z��3���a:�|�!�'D���@ͼ8�����'��c?��@��#D�L���,����G�\�J/D�����X�P� A�FiD�yz�9T,D� �@`��d8@�%)3s쨝�Q%*D���w�.H��F � G�,4	��#D��ɣK�8���Iݞ)�$�Aw�-D�c�Aڼm���x&OF���*D����,T_*��%�Z�+Ȱ	�ad;D�t@7N��53	W7˸`�f:D��Z�N]k����iV�	�L���+D�(��H���0k��u�0d3��5�ɧu��z��zy���6�14���Qe�7�yrC@�WQ�@bӇ%�T��"�ק�y�A�^�R������jy!����Mۈ��s�T�2A�շ#I�d��L��F�1�"O�Ց�(I�vϠ�����eQ���"O5H�@0Zˆ����ѭx�l���"O�88A%.��\�cE9}H��T"O� :�5�ˍ����CU�%�~��"OД��B�"%td{ҩL3-��1+VOJ�DFh?��d�>L����
# J!�D�M���2%oC�h8�ꆃ��(!��X�6��c���T
-�"ڵ)�!�DSW?�$"�Dɟ4�����"Ja|b�|�m�4V��!�"��r� ����yb��,��]���, _�0	R�L9��<Y��IU��Pf@uB�z�CGL!�D�!��1+���/	�j��fbշp8!��RQ�1[���v�ڝ2ע�!O!��koލW��-l�����!9!�����v-�h(���.+� f"O�MCCBV+�D1R� Pn�@�d+\OD�
�8<l����'|3 9��'���@� �4VZ�P���U�_�`�YS+D���N&*��p��JT�+1\ A&�(��e}��?ţ���u���b��th�5���,D�V�Z ���fj\�� �V�V!���p�|�ф�]�8.B�Sϊ�Jr�	P��(��y��b_��I�p��\��z�"O���7@�s>ag�#�XH��"O^�+���q���
�:$�&��"Of�1��v:��0�	8#Ǿ4P�OB�=E���y��d�H�,�c�� ��y��C����镄G��x�H�����hO����H!�ԐyP�,���a6��1HI!�䒐 :��[HS��9bMcG!�$إD8b��6��}�ܹՋ���Py2�D�1�e�����+ܩ�ҦS��y��;eLf!8���͆�Õ�Y�M�-O~�O?7M��;�]�� F5h@Wj�5!��F�1�x1(C�
�C�Ȑ�ђ3+!��̢Uꌸ"�ț6U�r1�"!�p�!��.U��#��K�X���£6՛�
O�!0eT)d$q�f��w�t�87"O(T#w*��4�ܔ�����F�7"O69rj	S�R0�!�/�0���"O�A�a�Ux�Q��Q�|����'4�d��Hxf�bpB���i\���"�O�K%��bf@X�%;����A�'+1O����
�,Z@���#��Q�P"O�I���K/�q�Ƀv�T���Ot����(���{�� �$8��n��<�t�p�"O��f��-8���͚>���v�'����O	8 f�W��|�'�P��*�c� �!nQ>[��	�'2�h!��^��M̭*Ș����$6<OT�Rg웭?^"�sgP�
8��S��B}B[���|R�<$���+s%��[�v]�41!�D�8&�����$��*ĔP`	�6n����HO�x�?9Rf �Zᢃ�T�`&�95&s�<-������z�ڠ��y0�Q�=�!E(�S�qT.�����
{�Ibi�Y��C�I�id�� ��v�����D>��B�	�k���c���3mА��)�B�	I��JT0iJd�8���Z�B䉹mR�[Ō�K�dD�>.C�=cmZ�)�*%�ΐ��m �B��/@�&�+�Ahlq!e��E����hO�>=�!��Q�� ��Ηq�I�a*D��8�ݫ�$T���ڵ���&D�Dɠ��:
�ŋ���v���<��哼W�@�ƚ!c. H�$&� (�*B�	�7R�	r�=����D	F��C�)� ��;�O�[
���A�;��D��OL���	���#�`]"8a4�[/kԑ�PE��'Y2v`�P�Va���.�KuC�yA�5Z��s(�%	DXH,��y2��:8\����<��e�T��y��D1������%������yמz��kV�\�"�F=��W�y�,z#��B���6!����U�y�@[�F��V�'�4�rM��hO\��),4AY�J<<�M*��8+�!�	)\y���	�dpu�V�L��!�D	Y��zs	G&uTN��G��5�!���#�L� �EC&P6ڴ8�+yH!�Z]���*e�T����b�D&}R�D~���ie�p)Ke�\��Z�7�� �1�'��<آ���\�Ȍ$iǗ@��4I����|G{���=�P�$,G�; $H2��=Y�!�D�"L!���ҥ�8C.!)�Ƌ"���G��H����[��<�	D##v� a�"O�4IѨ\�`4�a�X}(A"O@vkPjc��ȥᄎ&��Q�'P��<5��'jQ�Jah���=d�B�	FZ��)�(0W�Ή��

o�,B��/n\>�c�^�CP�Y�!�L7'����%�IOs���ٟ'�͛U�I7?��O|�=�}J�
��r��}���T6FA���O�������{�&��O`�`�����Tj�������'����ۻ��t���D4,����b�'.!��=fyD����tvp}�"�V@!��P�|�Bq��!��Q{�u���k,��(ON"|�g�߄'uXRL��j+�h�T��G�<�eǐ�C���a���,r��2+�A�<a�EۧR,�P����d�C�LY�' $�=�'g���1��8����֨�*&?����-�PYc��� ��:#��E���H<��O�r�'ܬp�B�0Yꨘ��``����'�85 U�:*3=5�C5 �$Θ'V�{��%m�� 덦-���!���ē�hO��^����I=�@C�&V�~y� #"O\���o�@�ࡩ�+�v( y�"O��pG�5��1�J<72A�24�|��+	�8s��Уn�Z�PK"D�p�g��39:�@� n
9q@�7�?D����nuX��&�� ��=��+�O�ʰ�
�I�
x���,.�@�"OD�����@��$jw,C+\#\���"Oy���Y�� ��G����"O���0o. ��� i�2�t3�"OI t��j2���f�L�Uv�e�'�ў�gm�
U��4�V����b�>D���.X�t��:b�_6j���;���<��}�����8*)��1�nP;w� ���hOq�|��'섓S�F��"mɴRz=���.�ŞL�h��d��~@�բ���6��x��hO?m��Ѫ��Y����3�n���/D��� oR�/1�$#����5h&�3D��H���5�"�TʲR�"��q�&D�XvGʳ$��У@�K+g0����8D�4�&�Q�8�ei�-F�&j�����)D��A^�MF��C`C L�\,ұE)D�\�Ճ(}�xh!�ᆄEH<ȱ�!D�L�����B�cP(6(K�ZrO*D����hɔu��	���`V�U�
<D�0r@΅'W� R@�15��=U;D�� >����]	��)���8�@IS "OR�R��k,��A&�T��$!m$D�|2��Xv������k�B��)D��kc�^/ �`Q���C�*}�2A(D�|��N�7(�:�1WN�/M��y[1l%D���q��(Ud��9�HCX�v���$D���B�(z�nit-�LF��$D�0������x�*Gr�O#D��i�ʁ�D�$��@Cd*� &�#D�| 6�Z�ZFh}�k*s�e��4D��0󂋪*���`�� #�ޤrp�/D�0�G�J�C<bLX���O	� a�.D� ��Yt�����D�FGPH�Ł,D�d����
L ^���A�Z�8�5�)D� ��h�0��(�+Ә|4$�{2�5D�D�jK�)e�)p�џpr�
�!D�ȈVGK��b��]�A2�A�׆+D����7$�h��O*B(��k=D����ĿSf���)J�1�� ��o0D�<Jbe,/�(e�R*�`����(D������ELr��7
Y2BsƨkS<D���b�U�G_&�J�j��2J���D�8D�\2� ��}�Z���D��H\�d2D�<Jd��q+�MrEG��a�30D�����}T�%y�!_7f��e�,D�P��g5n#�];f�4�B !ա*D� �$�	$&�N� �XT\
�M+D����$	�{����
)9��Pdg��SA'��Y���S���Jh��a�(�\T�#bOB�!y����^�V(Ԅȓ�}`%��6�MB�nʋ3�܄ȓj��(Cc�����8j��R��X�"OtM�F".0�i��m�*P��"O^�H�gH���!H��*i�)��"O�C�^t�)sQ'Q�C�`�I"O���qf�n݆�$�K�=�,cw"O�}��l�z�

``�Bꊌ8�"OV��1Љ��Y!F���{W"O�x8⏀#��Ԍ�
=h�p��"O�D!��i�r�r7L��<	�x���'D��#P�?ba�]�񯗛p�:�`��%D���@i֚��g�<������%D�,X4+҃h�J`jG����6D��q�M��7K�m� V3sĀ)G�7D�DP�'�x0A�X��'���ie0C�	�`��Pi�i�"�$��U���B�	�G� ��ҩE�o�m�L����C�	���$*4�R<���Oͷ0�B�� J���*7�T�4���sfN�)�B�I�5��(��"Ϧ���k�tB�<=���lS�b�$� �R4fRB��+O\��w�Mc�X�9�ˎ8`�C�	$M��J�7J[.��%�!*�B�	�9���j�I%6�uB�0F�B䉥K�� Y�B1 F.��1 ȦB��.	��� ��l �4�c	IޒB�)T���'J��%y!��	N��C�ɭ\hlU�c��;)ƀk�o��'C�C�Iv|<:q� ���C�Uq�C�$��=�`a����y�1��$8��C�	�p)�h
CA��il��C���!*�,B�I�<�~����9Sx�0�wH�8��B�I�(u�E�"N��J{�����%�xB��,(.=8�b�g_HlHq�`�B�I��̹pd�3��27��/8zB�)� >���0I}�J��׺Qd����"O�GdA5 (T�EG D�L�# "O�H�a[����i�0Pj��"O�hg� �Ψ���J8dW���"O�ۓ%z�邊 m�UJ�"O~|�p瑤Fc,�*釣^|�ѥ"O��5f<�� `�)��4���;"Ov۷�1"Ȅ�����B����e"O�MZAG�o����?o��K�"Od0a�խV8�H��ҤKr�QX�"O�����7�8��se�!t��`"O�M��ň�K_ �8E#Ⱥw��@�"Oz]�U$΅ZQ<����m���5"O�Q,/;�Yj�	�VQ��"O�]s��:�r����S�_��]��"O���q# �V:�Å��/�F�92"O� �PC�9Uܥ)��mTlx�"O��tk��1�f�&A"EI2"O͡2GЫ<�yq��9~��myt"O�Y�+CM%�)Qь^2d<-ñ"O��2�K�M/�xx��XͶl;"O� ����W-�U*F�b��,�7"O�P�AoI$o�����o��y��ֽq�H`�w  �2�\�� ��y­ҟ(+�l����,F4T"�.���y"�� uF���IMh[XȣR�O3�y�6eE�y� ��l!Na"��J��yBi�6w��aG�:vV����
��y�꘎k����ҧ�m��pe�'�y������3J!1M���U�P:�y��#Z�8�k�� т�r�*��ybD�p�d�����6���Ѯ��yR���q�(��ۦ3l-�6�:�y�!�=:�bŻ�%�!
��RU�6�y��(&R��/Y�B�ݔ�y��؅,�pa�#��<�,9�-Ќ�yR��>yL:��ŵK_��"B!W�y򌋰Q<�QE�?隱"S�Z��y����'����P㑟>��qk���y�
��6�&<)�[�0� q���(O��=�Of��1`"�j�5yrn
f<�h��'Ϩ��t�*TVP�R g'���̊;�(O?���=�@Er2$��5Y:����O5
!��X��u'/
\h!p#�&h�l�,�D�5�g~�B�=��襉ϐ	n~�NR�ʐx"�V�F����V�\v�աQ,�2 %XŋD	��?A���PlxiDki�xh� �Mb8�H��E�/�}&�Xp&-�;)�θ�!f@��2T��F D�4%�ǧJ#�%���_�z����r����t)ķ���s�Oހ}9��s�Rex5�E�(  @�M:�j��"O���y^l�H�jӖ`���"���ᦽ���Xa�b��<Yo��3�"�pH�,bd��b�C61�H��ɨ+�>hc�� � Xa��`^�}@�%1U��`SK�<f�)��'͈y�TNUA����Ȍ9�h�;�}"#��$�a�WR���oQ�#2�\��SbX�=xfbĂZtZ�����l��I�%Q�~��ą;2<!)0΀';��E"%�_EB��s��R�O38)���e�+7 ���HY�"����Y�g� ��q�M�_�4e!�إ{��A�O���X��+҄�U���$��=�nU2�o�1,��0�tI�Y��y�/R�-��$���Z�5�(E�2�9Ӣ$9Lpɋ����0�\8S���,HƔ��I���CeR��N�D⑟]���OL�	bў^�����oN=\6�Ap.�C �ѭ��B%�R YB�`b��+n~�:�"O��Xv��W��P�w� U� ��Ϛf:d0u�H'x^p`8ňZ���PN~r�X��.J�dS�'Q>J2���O3�!�DA�? ��s�n�v�X�i"� Mr�LC�/Y?g�<� '���#(.)���6`���[��ӊ�(OP��(�\�J���Q}���Q�'�R�����+����Q��(s���3
2X����6���k 舻Uت9�~=���
8n��|�
\(6�BM!T#}T���
F���'����L�kfS�/�~�+"o�� X���OQ:i��d��6�����ޓ.�#�'V����(4<��i���hq���>$�P�*C�@������-R��'?!��!�&�yG�S>B��E���Z�8��x�N���x��P$&,�H���4��l_�[%�Ir�� e�p�{��R��	��b[�$"HV�I��0�v�-�2]�PF\�vW.��N?X)�y���:�d��bÞ@�ht���W&)ĵA�	�L��Pt�G�{�rq��<�O �+�W������g�I�8]�q�xrAυ(��m����x�>���C��P�R�&
1�i���l|I�&�Y�T"-� R!����J��s鉑i�΍��ȟS�}���+8��,�6H�Lc��9�@��Ik��	�0��8���l��a��(*[n$P�Oʤ�'�W.� ���aM�`Θ����z��oӛ\΄(�FM~B���gא-�2�<�v�C8H��2T+�`��dyf�qX��U(��B�R���g��@`G��	L�d�rn��R��2_����4�	-���6hG@)6��*[|P���#C10O��@Q3D�r@����*`��q��E�	�1kD�?�"��F��3�&� `/z�2W�"D����J�<R1�.¨^,*�C Zn�D���Q�W�6���a�!�4����$�� #�2�](a�	�0"˷s��x���\=K�tC�	�'��.[����W�١u�Z1@2@љl�^����ެx��='I��&��v鉠��QAw%��O�J-� ��=/����N�B=�`A �(����i�ʀ��֖�<)9�f��s�ͨf�=�neA�#��u�^)\J� >%F@�<A#��>!LT�P"��R 䝡�A��6��)�V!�W�_8_?`��"G��$J
P�""O4M��3}Bh��G�%�zk5+ӥKeD%���yH����V�Q>{;O���P���(:�Z���'�xQ��"O���P�5wwr v�]%��,�4/��\k7��c2�A��	ȣK��"�w��@P��<m��h���+?��[g0�	���'�xj�� �r���1%�mnj�۳��&�4M��,zE��llh����$�Th��
�@ݢ�`���#�E� �E'H����E���!�O�\�i"�t�3��(I�,� �b�[C('�����]�B���Ox�+��	DB]z�%�;����i��t�ȨJm�@J`W�"~n��Cศ�c�9""B�3ϭYZ�㞈�5�.�a�TMǘ8�b�sj�8	Ֆe���Q��y��$��~��ՉNE :X�����Gܓ �X�|�'� �Q�l+[���r��0?%���'H�X�V��6#�j�)�zU �d̄m2�q�sle� �ZB"*�����7�n���;]�	�O�����Y5~����s�Ȱ�"Ov%�G�X�+� A����$;1"O\0�-"�"�`���HJ�2�"O�T��ɖ+O��$R��M�_:���e"O�iдB��-�%KOT�|,8���"OFl�th*�8X94A�e?np��"O�,�G�V8~8.!���T�|�к�"O���GB����sC^������"O���2jT�(u�,�CX�g�\�07"O���QN�dU�!P�'���"Oָp'M�A��4i���q�<1�v"O����J�E-t��e�.\�1x"O>�9��^Q8�rË6t��Y��"O
pA5��t2�
DIY^t�ɕ"Oi��@V���	Yđ�T"O M�%.X�(:h�;�ѢjQ�L��"OPt��e[2��R�EM�?�| �T"O�p��I��P��-c `�%��"O$رRn(y	�˧E�^�V"OFxŏ]�m����֨erT��D"Ox�"���"���c�L"-T��hp"O�(	�ė;?GxxA7#�D�3c"O���[�ƅmNTkb�e!�d��Hcv�`q��L�<)a��کNW!�� V�0�ct�(��ɿ3���D"O:p)���8r�Q�«Ãk����t"O`d1҄	F�����2�R�"O��"Ʈ�0i�%��NT���`�"OԑrQ��.i�@���J�ܼ���"Oluȡ�_�B���84냹S�ʄ�f"Ox\�e��4,~�1�,%��bg"O���C�Q�"�
�nwr��"O�Z!�Pa�	�� )`�l�'"O�S�gZ<N(H��L�M��x�"O���,M���4��:JKl=y�"O��8�FF�S����/N"��KW"O�A��¸Y�����Oˑ\�&�A�"O��a3���\Hp�.�%)�\��"O �&FJ�d���(����4"OHɘ��\Ƃ �⬖�-� �q�"O4�w�]�t�'+�<1�j-��"O 
��68(rT� (iL�<)"O��%hW�x�|�sDd�+l>�!q�"O��sk�VBA��Ԉ~+p�q�"OkgLT�}k�" 
B�-��"O��W�ڑ �����&��3�"OZ=`��թ9F��#B�8GTұ""O�I�d"Ԯ'��)�&�-`کCB"OtibX(r�f�� ʉdƅ�7 !��Yd�{�&/<g�e��%6)!�d̊T���uT\���k#!���fl4�Q��р+a`4���+X !���kh��R��Ũx6�9�$��!��UmU����Rz�T"�7Z�!�D��p�XlǮU�s5,*6�T�E�!��H�p_�I�$�/]�l�ҥ�L��!�dQ..� �J`�\�|��N��i�!�d�+Q������5�\L�D����!��d�P���;�V�@����!�!�$TfV�h�&�ŖI@�b�*T#!��Xm�ɉD�ȵq��F�2�!�$\/N��ZЉ<�y�o�}�!��]�,�)��t�,�J��y�!�$�Q�X��KD�C�X5�2v�!�d�*���O�3 ��1V�KcX!�$_1!��I��F^Q�0�Ä7*_!��I�*Q�D�	Ig
�)���<	8!�$�b�H03�Ψ[���T�%p!�d��nA�旖:9xA����>�!�H/*����2(�3�1c��6-�!�ā/,;F<��"S�?�����;�!��=e�����" ��³�U�!�$�)J�$! ����O8l�!�D¶On"�
U�]!'Ժ��V2KT!�D�F��<����%ɴ+�	ZE!�\�02rL� H�2q���"��A<*N!�$՝M�V���*=q�����$X�!�;uu4	:P�X�� :�ԟd�!����X�qcGd� x���!򄚲6;8p;��D:;�)Y��#|�!��5'��EcTo��N�`��KH6�!���7��q�P��<�QS�H+a<!�dS'�ndsC��5 �â��%!�Ge
D[�甙I�<�hE��=C!�Z+}����%*F����ZBJ�,k>!�d��=�Px��Φf�����ם}!�$�V� !���v�$m�e���Na!�D�af-GB�3�X��v���Yn!�� j�����2�LY���UV�:T*OPa*s��[o6�����/L`�y
�'�@kΟ�
x�lHF#L�N�{	�'��[G�=�,Y�(�,Z�83�']�5�A �'9+%����
�'���s�̒ l4 5z�g��LӒlc	�'��H:@�Q(eВ(z%cд�p���'�T�U�X�OQR\�W�
�h�̉�'��x�(\+�p��P�� Y��p�'�4{�G��@�b���c�Q��u�	�'�ޡ�ECį:Ct�1��ܰS��|)�'�d��K��L����!�{��Ш�'�ڰ��Kˑo�I� V�{n��Z�'�̉�TNˢ
FR�£I<9����'.$ QON�m�D4�wIOg4e#�'�@��%�#��Ҥ$�)B6��	�'�v�*���u� (Ӆp�.:�'y�i�C��1����f�? ��'�&e(1 �{;��P�َ4v� z�'_$�B�e�6�窓�,
ps�'���f�D�S���mF%�	s�'�V���M�,��Y�l�8 $�i�'��Pr2���^���G� � k	�'�DJ��k�廁`�qi����'͒�P�+���������y� �
�'���S�J��&��
�q ͘�'Ѐ�iH�~�N����D����'5ƹ�2���W׌�#a��)c(�d�'��)#�I�\,bA��EOZ�ht�'h��Ѓ�F+C�Ԕ��kď@�^a*�'i4}�U���Wx���ᒼ<�2Y�
�'��$��#R(u�4C��Q�1��5��'S|�;�����l��?3��)9�'Ҵ�-T���e�9�n�Ⴁ�<�y�+��Yk 0�E��&;�����;�y�eؙ5���;QTE
���/F��yZiH��35k�k]��0o��NddC��:c8��𭇔��1���I�"C�I�21"(2�Y/iaxDp�#���C�	r�`���T;o�`�2��5{�B�	h��(�©ݡ#�DX
snR�H2B��7'���JA�H�v5���z�B�ɸ(U����%Q����l�*�JC�IZdN�Ɖǜ`�����S�VC�I�>L��]�W-����/Zq@C䉪ZrDdxtN[��C���V�jB�I%n�A�Lq̰}�0,H�#��B�	$��Q:ЬԬM���IT�Miv�H�?9M[�����-s�@��N�O�|����6T!񄜡	%h-�P�?'��R.�X� b��arꞭ7+����Ö�z�0 �1����p<�_^��E�H<ـ؜��1���W,H�Z���	N�<�R�VT�r��q@׮SJ0�2F�|��@�X��\j6���Ƽ]i��b�+�_���I��k�!�H0V8��H��1s��L
S��;q҆'�\2�MJ�t�q��'������VZ$i��YB��	�'�Xq���Z�{�,���%�e���N'<��i���'���ˋ;b�*%��%��H~ܴ9	�-�%�$̇���v|Z%ˎ}F|��V!E��q���@-C���o��K��t��P�OX�c'��:��O��|�eݚM�F��v �XpT�["O(�$cQ�G��� b�R$:�l�bA�ɤ8x�D@R��|��ԐtIvQ��)�3L��tl7��xDݒ,6���CS�;�,�Ѵ�ҜD�9��Ͱ?� y�6䓊<�>lr��ęo$D}�&�'0�xe�|,[i �r抓�Ql$�Sn��y⌎�0L8��@gʋx�I��aZ��y"h���i��$��b�*07�ϡ�y�+J��Q�˖��� f���y��C ��p��
|�^e[����yr陒w58�Pqc	5w�H@v�V)�y�ɖ:���vF_�lj�mq�C�%�y���q��	]3\�	�����y⤃�g����"F��I��}�fK���y�&�-iI��bsǊ�}Dh�l��y���3�|Ua�f��pW��Z�I+�y�����	����`�#�E��y�C���d���#!�񴣙��yBc#\i($Ä�,{��1�7���y��b���,���B�������yB�ȧ9��p` ��M
�#��y���a�l�"%Я�:�*�@��yB��51�x����
�������(�y�G�V)@)Ң�USX���=�y"돰pc0ƪ�R4�y1+��y�HT�	�Z�(���xL\���̄�y�+�@8�9XCaJ s�UhT���y$��(�"PI�v�X n ��yb�6w�4���m�gN��7F^��ybd�_���a.���{����y�/:}y{�%����X�a!�y򤝂r+��P�)�$���k�1�y�@��!��|07��+�����P�yHj-L�s2��&$��0�/��yBkO?HX�EI��a�%�͓�y¢_Z�T	�oΉb^�Un	��y�γQ�T9KtA?y�Ő!E��ybN��	�@ ��:)XZK ���y��^��\r`an�	]Հ�ȓ!RJH�aA�_e�0ѧo�R���n��� N �Xu;F�޶z%8��!�+�^�p���3l����ȓ�X=Q� ��,
%Qn^�B�*I��M���\��x���y����.�n�<)ro��"f8���T�zdv)�/�^�<���_�s�|H�q�ޟ%i�mgVS�<��/-01<�����d��;�eMO�<���,g=���4�I�u�ܓֈF�<	GD\�aS����8L�r��~�<�$O=5�p:A�ި(���:w�@@�<A�h��th6����T&;����Qi�<R���{R�*V��d�l�XB�d�<	�hS�4x8��T�|/x�0f�O�<��j7R	�x��#�Qu�H�J\�<���A�gP�ڕ,ҊS��\�<��*���dA���)��hp�I�`�<q 
�X�iF�ܬ2��T�CX]�<q��E�,e4<��g����G�]�<�S���z]�u�?w)�(V��B�<����

lK9qp�i{�BD	#��C��+-�r�cY�`Ȥ�x��,5��C�I#q؆��KA�DȢ0�G�\q�B�	8)`-23lǷ�(�3F@���B䉯oG�����r��١�mު9�C�;,���f�Ƭ>���I"�];LVC�	�-r�` �"v���'�2;B�ɩW=<\5�Q,涉�g�F$A�C� &(z����% ���z&�;G
|B�)� ����x4�BdLY�+R(��"O��0"��2l�Pj�<�E�"O�Y�@e�;���H�;�-(�"Oʽ�BJaJ@�h�ڋ,��=!�"O0u�d*O!h�,q�Q�	0��:�"O�H��%C7�e���'c҆)��"O�����$ =������oӒ�"O�ij�Aez��㏁-=xD�R"Oj5�T�n�@eq0�͞jA�[�"O>ar���wE�<1P�i>��p"O�1[v̟�aJ�#���A���C�"O��S��,Qܒي�� 5kD��3"OR�9uL�z�ԣ.�3�&��'"O�i�2�ˍ)�0őb�DQ�2�ʲ"O@��G�Q/^^ұ	���:���"O)���8%����S��r�V)8�"O�5��CX�mI(�@�%�%��ЙE"O�c�MX�!��y�� �(Ѹ(r�"O���ح�	B�ϒ'���2�"O����9^2 ;����&!�9�R"Oʔ�"��� bF�%�	�F��v"O*x���8�@�Ye���YQ8�8A"O�SnB*=�8�c0*�}�����"O���� v���W�A�=�j���"O��a
\4(�k�FV�b�$0�"O)i��ӫ@C`�[UD:O`>��"O��	Vb��M�
����ھ[S�l��"ON�:�JTm��#��(?��$��"O~���@7/�X �W��I��kb"O
�x���
9��"��9?�i�A"O��;"ᙣ]�J�9��n�b�QP"O�*�-�{y2ԂDO	@���r"O��[	E����Q�D�C�ɡ "Op9��HŘx3�-� zIn�;�"O�����N|m�i�d�L�20��"OЕQ%��/Lf���LK^�2�u6O`Ĳ�����X���B;Vi̩)��O��V催M�1O�("���k�X��]�V��B�����ڦ&	�&z3��X�7���h$Q����S6@�52��8 D��01ǎ,���x�^M�'��c>ik�`M�vnМC�Aެod�)"ri�>y[��<�{�'k�U:��� #X�)�N��z<PK�4J&��"~�dbբoZ�Ul��U���a���eўD��>w�Ȩ�U4��Y�KƦp��#<ь��?�:��<l�<z@ɕq��}0�N?񤒫�(O���I�Q��<wR%�&ɒ�U��3_�䰃�)ҧ[j0p�C����B�q�20
j�oZ�.~Q�"ZB�^�<�~��P!W��-9�@ �(O ��ӌe{b�ۅ'qМ���̏=�M�K�����?��󧖸�M�C�Q�
0[ƃ�Q���1#l�I��Q�b?u���52z�rD��#(XXz҅�>���7�S�OAtA�ː�+,,�ӥ�ĊV��#ٴh z�<E��˨w�-(C��![L��� ,��:�Q�l�çf���0�G��r]����0�n��>	����DV�E'��y�A�v���g��+��=��y�IX.`����գ�9T�e&Gރ��7ړ^<�O(h2���/*j�[�'��]_��t�'	�#=E�t$KR~䑲�T\�{�L]eX*Ey��"�'�����6�,���"���-���'y�xGyJ|�b.V�*�bp���3�J��6��I�	o8�D��kJ^:4S�Řq9�-��N���'8�)��n&�iO
1��4�zI9�%�Y��4b�ٱ�tu��^�<���4Z�d��jP�.j������Z�<q�曨�|4s�\*`�l�@ ��Z�<��_��e	�H��=K<0�bW�<� J@I���-ˎ� #JT�4�d06"O$0KҎ��(W�ѺQ�Σ8��Q;"OF)A�'�*W����*�C��u۶"O`�C%P��.E�7j�`~8x�"O�IRA�Kl������ !.����"O"��"�G3lj	��@͟]�2�I�"O X
j�<&Lt�A�p��dз"OY���<��p;S�˟$��t��"O�lZـ9-�q�W�Htm]�"O��Q�i� G~l �ϛ���h�"OƱ�Wc	�z�r={����Iu�A�"Ox�i(SFڭIU�lt��"O�3��K�\�A�Ư4j�9�"O��ؗ�(n���Xc�H\�@� "O�iB��lh��0���`N�E��"O"��g��7�d����r��ea�"O��"@�i�|�䭈*���i�"O C`"�8u����тl�,�&"Ofy�q�C~�ӡ�lg����"O��5%��A�Ұ3a�Pcn(�6"O��;犇,w�����x�#��-�y���Y�tآPZ#w�,�Y�h���y�ѵX�Չ���4YW Xy�*هȓad8�S�{�HrÞ�k,؇��RsG�?/SL0�5�cCppR�'�2 *�;OXء{�k����;�'�V���Ҩr-z�FE�"�H���'B8�s���.��`r���E�@��'H\`b�ȒC��%1&@'1
�0�'��Њ'�׆;�^�H%��)(� �'���#у[�@9�3���N���'����vEGRع
t������'��(%H�6�0��JW����'�؀Z�M)P�>{C��o�Y��'����>���LP!Vi�M!�'Nb5�o�Y�s� ��Pbp"Obݪ�ʋ)F���� y�aR�"OR�$�Aef�R���Lv(�R"Oh]0���vՌ*���z6�a"Oҵ(��ܾ#��i�([>v�pȠC"O����<$�y��M�US�1�5"O�X6G���t��0M N�T�"O�!���4VG��LFn�;R"O<�eEً\��\�'�%�y!F"O2�`F&!��X���>9�v�#�"OT|�V��T�l9R���0� "Of-�L��8d��b-�NnP�"O���2]u4 ���Xw�r�y�"O٪������3#[��u"Op�����Y�H_z`�z""O��R"��
�6ui؅QJ4ͪv"O�L�6�CP�b�
�l�X���"O���C�Y
�<�Q(@a�X�!0"O0�p!a�9T�|�!�&o)��"O�9��i̻;�i��9D �W"O�� d F�u�z�@ce݁Q����"Op�1�
ދj
�Ȃ!eB`���Q�"O1��&�	*)d�#��^τ��"Of��2��E�Lۇ�K��܋f"On�0j�$Crq˲юQ�mR"O����J��<c����JJW6�E"O��a"嗇� <�׊�$lД	e"OJyz˅��M�pKB�x�"O~U᥍�D��"Qk��!f���"O� �@[ƅ�rn���k��^�af"O]�f$��&���KãV�>�1�"O �A$`���ᶫ\|����"O�P�$��.*�l$iI�L�@�"O� B��O���F��U4�H�"O�D�C��\Rr�r�0�!�"O^ �C��1{G���Ӊ��<�18�"O�e�Ye�����W:(5Е�/T�1��;�L�j��NX���i��)D��	�XQp�Yd�f��|��&D�I��}�ҥ@bL_P�jD�0�%D����`��O0@x
��P�,X�r�(D�,�C�M�:��,��zY�9p��)D�d�� ��=�\�2ڰ7)��5D�`y��ȹ�8��d�V�\�ERSD7D��3F�Jrl3�wtN�*��6D�Ё@'r�n]�7eC�-o�*Q�4D�	ӥ��5�,x�g�S"(M�)�i>D���n��B��D�'��>��R$�&D��I��4C�d�kPQ�T�~�R��2D�$YD$�:\C�-�F
�豫*D��h�
�Y���	X?�
���
�'�쫁O�1{~�5�J� v�Tc
�'�<)r7�0G�Xt�E�Y�E���"
�'Q`Qs�d���< ��JR�=�:H�	�'3|�h�JYش��@��a��9�'��tcv�P�V[[��ޤ`6N�H�'q.��NI�W�4$[�ْ'+���'C���3T�ne�e�H�M���	�'PV�3�DβS=���Fn�C	�'�(���' ��
I�ƃ3T���'L�����4	�X��'� ���j�'���s��F�#W�Lq�̉%�P��	�'i��;�DM3��ل�'�Z��	�'� �S�I	kDt��)J',�(�K	�'Rhu6�V	��Dj��G)8@�L��'�R�����Z�¬�3�X�(��`	�'G�t`�K�8�Z,1���s�0X�'�T��G�0*<\�����'ºE�]�9{�M��Gh �
�'&��ᄥ���e`��� <@p�'J`,���m����"���'KrXL�<Yp�#%D����a՘�y"J�1h5���W�R�?0��֎��y�雅v��5	��f}�Q�e���y2Me݆�b��V�y�Q�� �y��z΀�@�­@RX��u�U��y��U�g��Y�S���3�� �#ݽ�yr�qH~�c ۱*���v'��y��
!A�y�s�&��ڒ�,�y�
��v���2�Ť~�ت��߶�yBM	���i�H�!,�Z割�[�ybi�n������EvL��E��y�����XW��
]����yR�ۢ�d��,��T�-G%���y�葆)	�q��"5�!Rv+���y�,g���[�O�m|���ȇ��y�F++}�Ax@�V�`f|����ߟ�y"�E"�T���_)p�\��A#���y�,Q��X�5a���y�g7�y	6lvFe�$�[=	�BzP ��y��лZ�HK0$�36X���N �y¤�!> p1	�n���,�Гa]�yR+=P�i��Jv���3���y
� ���a*�.Fr��a��0ih�!	1"O����*]�"��C�͇�+QbAB�"O>�:P����a�,�RJč�F"O�����Ďɜ��2��/w��P�b"O�!1Ŭ޲���g�pτ` 6"O��S�B��l�t�0q,�L�RM�C"O���(Cd�
m�&��$w<((�"OF�PrN��e��1���`g���c"O0p��Y�-��X��ꃈ}L@�:�"O ��"�#D��R
��GZ�i "OR���;.K�S�S&C���s"O�81c[9$ڼj��R!?��t7"O
�(UFFL��t�&��B|(�"OL����(A	fg˱s���q�"O� B�*�I�K�/�c�I�"O��c�"̔������^�U�$�f"OH<b�n���2x���?`�
5"O\�Pe�$ (��"gn	^Kd�0"O��{@���$��!J�I,���"O�=5�5O�Ti�@�:8>EJ%"OH�&F��
��������e�����"O:�෈�w���i �ʢ��m`�'���"a��p:ڼc2b�#s)ve{�';��S��^"Ӵ:�t�'��x�,��}Ǝ�±L�5f� �'�>\1��ڼb��с��}� �'�4)вi�:w5�m�WK�6n��HJ�'�V�"BX)���$�X�D-��':ܱX�"Y�*�pBWG��K��]y�'I��UA�}F�s��<O���
�'�b��&�A�rɠө�F~��
�'���ዄ ��r�N�?��q
�'/��s1�ɵk
,�Qb��b!)
�'F����H�tT�L�&i���T\k
�'��J�څ,ݾ���>dn(h��',�ؑs�#Tlȃ b;�p�'���a�ѓI�`xa5�?^j�`��'��ygd�& 7��؁+S<(�|�
�'(<�xDM%�|8q)�h{�Z�'��d��.yk^���G��^ް���'M��3��M7E��b܊ -<�(�'���x�b^�E��]�P�y@
�'��hB�	!�ؙ1D]�nM��'��!X�`���TU?U5b��'��1�A�Q:v$�(��Iœ:����'��	�3!��bat׿'�Fl�
�'���׭B��8�� �"K�Vm�
�'�V0"2�W�l�f�	�a�G"lDr
�'$E�P�.��lC�A�<qn�ʓnAf��K�B�l���.��ܱ�ȓI2(��!K�F��=��Å5�.Ն�k>\	���I�rJ|��ۥ|�Ru��cX��p��.6=N�b�U��ȓb9bl8$�ɹ;[L%c�݃p��Ѕȓ,�Q���@��3S�4�^�ȓ^!�l��!$�bHY�������'4õ�n���f�Īk`N9��D
^��u`�I����aT����M���ks��8]�T�Q,4"ɤ1�ȓ�����mP�v�ء0�jEՎh��J�X�C��2�Qh0+=�h���y]��#���&O�B��J
%N����V��Wi�"����m��b2M��;YR�R�m8Hʴ��3�:Ml̆�S�? �H`$
!��E�]x��cq"O$�&   ��   �  �  �    �*  6  �A  M  �X  d  \o   {  6�  	�  ��  ��  �  @�  ��  Ʒ   �  ��  $�  x�  ��  3�  ��  ��  �  J�  ��   0 � M b" |) 	0 �9 �@ �G >N �T �Y  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0��	Q���鋚Iz�@pQ���bEd�)l!�D͢w�Zp!7Jی���Ќݳ �!�D��G����U��/�2��ߍw�!�RI(�:�#�E�|!b
�7��N؟�Y�,��R"�����M ���I1LO�⟴���IH��� L&K���B�-D��;A�C�Yj�������+�Q �m��P�=açɲ�'	X?>��LQ�/�}��M�ȓp�гv��?3F��u�Q�VN8�'xў�|2�i��-F�)cTNG�P�L`�3��G�<" l�}��G>㔀ȷ���u�c"�0�q��52Eс���|f�Ň�IG�=}��c�j��H���!��#Ȩ���BE��)�(�n٠�㔰/�`Ą�#��#O�"����4"�ȓ6Ѐ�����:�P�C�L[�X��B�ɏ`��A
V6�"ݶ)1�C��r��� �Nel~9:C�Tk���3���6��'f�>)A�k���,�`�9D�HU#�Lо�چ�ު6h�� ""D��`�\2/��RZ�xe�1��%��=��q�'��=a$a
5p�ZLk�g�>g�J�P
�'�R@7	ˌQ���U�̟uvLL��٠�(OR#?Wf27�^�1�1��8��RI�����~+]�u�K6tx$,B��9B䉹+E(�+c�]� �����O�K���$������Զi�d�Q�5c�$���- D�h(��#'��AP��i^ά��O��	��O?���g�2.>��!��ɲ3Ѿ]c�OY�<1C��=��eB[�BJ)D��R�	q�@aխ��6T�p��fV;p52�h��%D�<�@�tӀA�@#<0
8� ��>��<����1�+:΀������ȓ3����q*�*O/��Ap�W�6��Xߠ�:a�����,����1l�"Q��K(K��ݬ n��
�E�@OB�ȓY�pѨ��Tء�ckU�}�ȓM����9@À)Z�^'lM��X�P�sCHZ�xg� �DJ�����yt8��Şob�Y�kb�Єȓ<��0#�D�!��ud��F`5�ȓEt��V����IӋG��e�<��O��D��=�����E��T��	�	���!{�"O�hҔ�\����٩P���K"O�iذ%U�$�"q���"	��E"7�'��u#T$�0�ɭ��ЬՂT<�ȓvdH`ŧ�C�8 ����w����<G��k�E
�ԜX�a�E�ȓ2�,+r�N^�p�:k� ��?yٴ�p<�ࣄK�z=���6?<���%�z�<����h�\=�� 
:?R��G�P�<� ���`+E4vHB�a�D��y1��'�qO,�0sP14�)a5E֙v܀�]�����������E�h �H��i�0KZ�hO>MsG�S_[��0�#̧i��%H�d5D�00�J�(VR�[��H$s�n���6D�0�B��:l���s�.]����2D�@Q�ǃ>WV�L¯-=V���3D��CX<��aR���Y�%D�|1w�F?dLH(p�#_�`*@36�(D��@5o�w��)��@�:FQ�����;D���! +O�����ο	�p�WO:D���d�A�89����A�_xڤj��<D���J8=�{'��2Tq^�9&�,D�Ȑ�O��_V@jC陻"&����M&D�`�rڃTq�f�"o�>ID�#D��@�6\Z���
�L@���2%.D��z�ֶ#RޘQ�%�^��-?)���)eKP��#�ĂZ�,����թ`+�B�I�JA"�JSOҼ��$"�Œ9�B�	5��̠R/_ aȚ@c4f�'ʢB�	A�Ɣ3V2 �z�[�*l<FC䉽9t��L�fN��@a�(j���)�IT����ǇU6l$م��4V�RC�	4^����vGN�7ᇼM{C��D"$Q�F/J�=!�t���)-wLC�	!#����Ɵ$���5��6.<C�I�7�f�������л�I�,�C�I��:�X��;]b���!��	��B�ɭu�� d�T*Ř��EW#[jhC�I4F������ֆqv��g�Hq`6C�ɿF����Զ�H�����0K�B�I�i��@��팼7n ��'�,-�B䉋@�*)ʧbd- 1RW@�!�B��*
��Lؓ�E=^���Y�Zq��C�Ʌ	aЀsgU�]4v�1�W:�"B�I�K��H��� ?T.-�5i��?��C��.��'3��h c�7h���+��7D�4�換�[�D��e�5W�P30�)D��Yŭ�
�D� C ї6�.|�"�*D��(���(�,h(�PW�r5�)D��*���|V��ÍV����T�%D�X�a�,_ti
T���t�1&(D�Lqch��B��郑MJ�~s^���F9D�K�̋7c�2% Ă]�i�lu.#D����k��\Cfi�=Q��ĭ"D���ʛ+m�ᲇ�ّ��p�`3D�����Y�]j
as$�0�(l0D�P*���W��K풥`�\�Q��)D�����8���Oҫ�MQ�N2D�$0w���A�T�F�;6>��{�4D����ž�t��I��Depr�7D����.��y�F�b@��8C�r<S�)5D���G�} ��C�Fث��4D�`X!��~�:�aR$\�B8�� 4D��
7�܈�2E���3	5
��l2D��z�$\p# �P�m�I��]�e2D�,p�nP�#	�5�KU:N���a�0D�,xC�څ:t�$�
UcK����+D��w��=�Z��kѤu+^ɡ� )D�8�V���a�%�J����&D����H��7�*�z�@̙k��d�0D��(�P�>�X��ť�.{x�%[�,D����6J]�ȣ�

l��7a,D��7��+t������9w^1Be�/D�� ����[WLȂ	�?7@�:�"O�H�S��U9R�H�^��+�"Oj$K�͒�V��Aa��+Y�:]�d"ON-��IH=*=l}s��<���E"O*piAaTZ/��r��#�"`�$�'B�'���'%�W>5���\��C�	:�L�w��4zC�V=C�^)�I�X��ğ|�Iß`���x�������$�8!�P/9�X��)��x�	ɟ|�I۟�I��`��⟀��ӟP�ɟs@^���6zo��X'��g��I͟��͟8�I� �Iݟ��	����ɢ���)_�n_��j�(J	t�����П �������Iß<��˟��I�m��C
�Q�z([�'� 2��	��L�	ß��	���ɟp�I����	�?���N�]FR�gH�x�`���Οx�	ğ���������ҟ$���uo&p�2k� �F�5�F�YSb!�	�����쟸����I؟���ן��	��Т7Ν��!ZTF	+��I��t�I����<�Iğ0��՟���$G����Ah�8覊C�;)`��IƟ �Iş�����p����`������Ʌw��47�Q;#@P��b�@3Lx�5����@�I� �������� ����	�_���rB�@���SL������������ �i>y�����������I5k��lbGj4|n0�f��)2D�	����I��T�������۟��4�?���r��r��E��ы���0��G[���Wy���Ol-Nj��#���R��͑$DB�}�.*?�i��O�9O�tn/U�*���/͢;�E{���3��Yݴ�?���#�M;�O*u�bf�`����M?� c� �@}���Mτ�S�k(�	ş��'��>��k��N�@Lڳ#�=_�y�M%�MS�i�H���O�7=� C�e	"mw��Gͪbm�Ȓ�AY�-Jܴ�y�Z�b>i���ئE͓�r��>�2�[ƃG�|�N��eo��!�h�f:��4���#1R<`��e��)� ��Z5��<�O>��i6~(�yB�'4�|�t��:���r��#E�O�a�'Ŝ6�������dQ!xẵI�O�73��˲IT�]�	o��	�b�ۯ#N,b>�¤T��'�xc�ȅ�(l&����)}	xpQ���'��9O���ō�z�H���NQ){����=O�`o����k���4���4"��t��RDnT�Zi��S0<O�\mڌ�M��qvY��4���S�
fH����h#�z�o�"#�,�
$�P� Q����+!�$�<�|�<����xcG ȱcH�ࡥ]A~�Mg�R���#�O��d�O��?}S5Û�j�`M��l�:�S�O���d�֦Q��4��S�'-j���F�J�D��I�+��J����Έ�.O� K�ꐡ%O֝����'2��/3��@�Z�a|�b��0��O������9h���Ȳ*^�c ��O@�on��X��	��M{�iN� �,
ܑ��[�1ߚ�D �V|��A�iy�	Xx�!���-d$?1��#�Td��j=%ST��Ô�z�@�	��@��۟8�I����y��[e�Qӑ�4,Z�b$d[�A�X���?��]|��+H�I��I��M�M>Y(Q�
�ѩ��-ai>��D�O���h�&�p��ɐm�7�??�(E�.�*!҃ꂍD��QzTn�#&���h<>��� N>�.O��$�O����Oɢbj$w�x�A�[�*��%��E�O��$�<�w�i�d���'r2�'��"8lQq#n͍l�u��fP'��S��I��MC��iVɧ�iFk�~��2#����7B|�90nBo�F��f��^����|R�럃�u0�DI $�����	� ;���K��Ho����O �d�O���i�<��i͈�8��X��D�$�L���׭X
A}r�'�V7m#�������H5%	4��{E�@7�RY�C�4�?y3χ��M3�Or��aO)y_4:��<	�g�[xjd(r�
�n��2R��<�-O����O`��O����O��'4B8�F�]�Bk�e� J��'�xHA���?	����'�?���y��WӒ��M�Tl1i�m@�2�7m�R�S�'
�Z���4�y�+��O	&5"�ѳn��b�e?�ybaR=:5U+��:�'3��ş�ɎE^0q�D�$����޳e9����ܟ���şd�'B 7��4z$�d�OL��T�_,�3�/(�J�{��C�\�D��O��o���'B&|yQ��EN��`Ƅw5����O��� ܭ� +QI!�IL��,�]��?Y�AJ�|�pL �|6��Q�)b�'=��'���ӟ��S��&7���b�]AD-j�I����ڴR<������?��i��O���n�<�zŬ[�|��刕����[�u�ٴ�?!p�%�M;�O,Ń�i��t1��D�FIP
�3��!裈��#�b�O���|*���?���?���z� ֆn�*���/�5a�)O�nښ���	ϟ,��v�Sϟ���O�<S
�Ka"a����\���ʦ���}������lr���(���{��$'	�T���rV�I�#�t*���Ⱥ+��|�Y��h��e�i��(��R�ܫ�����,�I���	���WyB�aӀ�r#,�O�y�[8(&�L���*<"A��K�O��o�]�h���+�M�"��y�F80��	�UA�LRnXvK�6_S�l`��i��	*y{\��d��i�zu%?��=� DQ�gF&;�bܚEO��L���b4Ob����0oO�'�9~�t�pR*��m,0��O��������
%z��i��'[90ԫ��;�X��Ŗ�:|L�:��|�v�x�lz>u
S����'{��+� ]|`�u�W�x8:p��_3n0>�B��0X��'2��矐��쟸��:H�
$���>%<�a�I�gu��I���'�7�$e�˓�?�)�!���;e��RF�I�!B��࡭Om���MkH>�O�A�4��gh�ݙ�V1�|�,�E�YxԬ_|9�i>qD�����|��]�1����d��-t�6a`A��D(��'rb�'H���\�4�޴N��5�� ����B�>v�*`MS2�?y�4"���$�K}R�zӞ�D�mNB��04B���e�AЦ��I�w��QnZB~A�>��H���!��5�jM�S�C$7nvm��B� ,��IUy��'���'K��'��]>5��)N�1rd�K2g�&��Kj��M�7�Џ�?���?qN~��8e��wQ.�I5���X(�D� �0űar�0�>�|�D��M�'�����) �fQ!�bؽq@��ә'��0�`��*����|"Q� �I�t)�,�(j�: (Eh��=1 �ӟ�	����WyrK}Ә�g��O��D�O��PE�=HT� �G�_�a�LLcu$?�ɭ��D��1�4��K��Bǎ�.|��
R W+]i(�'}��B��M k��d	R��$��W��.��h�4$�g5p�2���/ |\y�S�I���	�x�I۟�F���'K�!�҇�)����ԫN�*y�q�'F�7��(jt����O��oS�Ӽ;dL�5C�̱C�4���a)�<1ҹi�X6��O�!{Tbu�8�&�0��i�@��]�7I��v�6�`��Û��畛�����OL���O��D�Ov�$R�tX�r�@�84Z*�ڣ`�^a ˓Iܛ�U�������&?	���>Ŷ�!D�5O|��pl[� �|}��O.pn��M�K>�|��(F�:����BG��pM�U�8��IJ~2���.(|��Rx'���'ej��2�jsbe�C�36ȑ��'c��'"����U�L��4)X�0��R�@�����'^�dlPAĆ�,�8�Fv�����^}�.bӆ�n���֩�>��q�b�Ef�h�ȴx$ �om~��*��=�%m�dܧ��K��� ��͘q�D�L�!��J�<��?����?1���?���kG�A1��s0�Yl�I�oV��b�'��EwӜ�*$2�h�D�Ȧu%�$A�ʟE��X��AןKk�a	E#�ɏ�M�PZ�T �LΦ��'VYs�I
�I6����h��_�����eӘ1��[�Y*��'�I����ڟ,���pɦ\zr��%`�PS����4�Iៜ�'�B6��K\���O���|*0�޳����f+B������J~�D�>ᦰi�d7-"��? #�V�T��N�iN��aRc��jB0+"�M����|J�jF:�u�.�Ę(*'|��AP/x����.s!���1�cbϖ���+T�[)�<��B	�:W�|�I��T��4��'D��>v�6�*ZÞ\Y%��=(b�� c����6-�O0�qӠ�pO��r � 7�צ<�KVRR� 	�DY�M��<9-O���O��O����O�˧��u�BcĆNΊH�f��8dD�����iJl����'�2�'�O��i���*A���u�Z�	V�Ѭ�z���q��i��6�;��IIJ+�7�f�x�{�;��N8��`ǥl����KB�&�Xل�_L�	Qyʟ�E��K���| q���PHYV�'o�7-χB��D�O��DD�m.��s��	�c�pfDǪxT⟬:�Ot�oZ��M{H>���7N �ÐL�U��a&@Yo~r � $����c��&{��O��Z �������~�<#���RF�$�����%SB�I��0F��J��A��L#Ao�P�	�MCcǼ�?a�D8�F�4�4�f��X�P\��M�eZ�qJ�3O�n�M��.� p��4���aK�HZ4�qa�X�(x�j�cԀGV�Y��m%�D�<Q���?a���?q���?��*�g�T��Wⅉ{6���S�ܳ���Ʀ���@ޟ$����'?!���C�&\2�䃫6p�adė���Y�Oܨl��M�J>�|��o� <R�ӡ��2$޹��چ}�⬙�c�n~�,ة}l��P��v�$��'�ph��nG�6W~	zP�ϾO��ģ�'�B�'�b���t\�|
�4zRAI���Jxi��A)3Ь��"vU!1�X���$�F}B�m�XYm�˟�ÒIW<����U&�j�aE+-UTog~ҫ՛b�<v��k�'��K@Q������<&�tt�V�B�<��?���?i��?	��T�� T'6P�f��{���^vb�'<Bb{Ӕ9���?��ܴ��GO�M*^��b��3h:�:L>aյi&�6=�v1�nq���HO�]�%c��m�脘���&�� 8AG�&8*��6�E�䓚�4����O���˽s�p	�W��%{��y�N�
�����O�ʓ #��Ş<��I��ؕO������@vA��Z�z .��O���'�,7m�Ҧ�$��'y`(��^,�*�nN����i��6W�z��ؼ��4�@L �/a��#K>QaH%]+�3�9_[BT�Q�QZ<���i�R� g�EP� -0�H�#��Q-r2��'-�6�!�	/����ʦ��RgB�K92�����<1�^ rucċ�M{��6�JE�4���ݥ�l�BR�n/��S�? �Q��%AB�E��՛P�z��2O�˓�?I���?���?������4MWl��*�dTF�I�.�%<�o�7�H���蟴��K�s������RN��n�3��

u��԰A���~��O1����#�m��ɃS@^2C��W���2C[�9�0�	'3�>*5*�	/c��%��'y�ɩ+
u[rd�<`��T��J�������]ݦ)
ԟ`���p�A�O�R/��j�)ܼRK�I�0�E���I�� B�q��OG���4蓠)d�j�i��L�'K^�P��i�O�![�����uvr+W bLkiL�o0NY���ְb���՟��I�0�	k�O�b���v�� 3�Ġ`��HuHɞ8��h�ޔ�W�O��N��?�;\��ĸ4H�L�p���
(Z��ϓk���muӬ���2�Z6M/?��K,�\�u�EP��� 'k��:��0)e/��b��]z�iy��'���'���'�"	
n��mP<#��a:��n��I��M���?A��?�N~R��6���#1�J\GH���?}ߪ�G[��)�4/+�&�|���`��c�ꥸB
7&�BT;���	�`\�l^��d�^�(0�x�q I>a)O�L�g�Ǿ>��T!ƠO��h��
�Ol�D�OH���O��<�лi׶�+��'��E�'/�t��Q�M�Z<���'h�C�$_H}��q�0�l�dB�-�;@�,��dY^� ����C�ckL1lK~�#ƹ%�DDܧͿ{&E�#]t�&�V*�ɔ%�<����?���?���?���Tf�+n#�˫�����}a2�'��v�Zt��?� �$Ԧ�&���`�C27pD��7�N�(C8L���x�I��M�����D�S��֓��ঁ�y� �V�2h|�q��@��܁����5UV�Xy��'t��'{r��R��(��ڢ�=���!Z2�'��I4�M{S"H��?y���?)/��<��c	4x)rBO\�dEP����T0�O�m�%�MKJ>�O]���S��CUv��ٹ��x}��y�ku3���c�<ͧ��}�_w�O�����޿	��b-ܢE#��S�&�O���O��D�O1��˓U�F��p�����nX�APe�,P~�y��'�	`Ӡ� `�O �n��F������ƬhU8���=L�Xrܴ�?�#� �M#�O�QZE�Ƕ'�RMZ�Ȭ<��G z0K��&7Q���L��<)*O����O��$�O��d�O^�'�����ޝl��3u���fL�yƾi� ����'��'��O��%`����)�=qD	4�ܩ3@�
o �lڅ�MCJ>�|r��M#�'A� �q,�j(`q���ۃv�h0�'�b�#fJ�2f�}i��|BZ�$��ß�叜:^d�� ΋�9?����ş��Iʟ`��_yRIp�ꔉ���O��$�Oࡸ��##��jU�P:O)^�q��>�����U��ݴ��<@F�CSh)O�.���&�~zH��'�d}���+������D�����ޟĪ�Hڵe����!Ș�RP,\+�I��������I�xF�t�'��C��M������a��\�S0�'[�6�>gR0���O^�mZV�Ӽ�Ǭ�)C�����J 	-�8�{#��<1�iR7�O�����w���<�(�ǩ!ʮ��SGP�f�]3VF؈T��*ξ�����O����O>�D�O�d�	pa���"�@$	��;��6�d�+�F/�>��'ob���'_�L�%uaXP��*ȑ�����>	�i�6�"���܏Մ��DA�\�u��==D FV S¾�z���ꎲ�u�e?�d�<��͜&�:u����a��D�9������?Q���?���|�)O�]m��|M�I��N�2�CB�Q��۴�Ɏ[�����M���˸>	��i�l7�OązR���)��qC�*L1�H\�7M5?��L�2���[�$!����P�̕S��{��ɲg4�
Q�u���I����I�8��ߟ8�� H'����@�w�tt��]&���O��nZ�5�:�S̟���4��/4�RuM�#X�m	lM'��J>	$�i�J6=�����~� �?$���ˁ}�i��Y;=t$<�A#�l�X��G������.���'�"�#W�z3�Ы��5C��"<)��i������'��'�哣\�H�0'�.-���2�g�^6�V����Ms��iGɧ������E�ˈ++��3��L.�jPhЉģ{<��h �<ͧV���^w`�O|���J$�����ڜ �����Oql��.|h� ���Q��h䈃�.p��&�ϟ��I��M�����>1��iѪ�1�_: @"͂w	� q�N���z�B��"b�*6-5?��/	f�J!��j����$̆.���R�W�7���g�	1�d�<A��?9��?����?)*��������h�ޗ-c����#����؟��	��H�Rº�y��P	F��p�ᔬ���W�&B7M�_�Şg�{ܴ�y�j�	z�APO9J0��DÙ�yB��q؉P��S�J-�'w�	˟����E��h��T$0M�֠�Wz�����Iޟܔ'�L��J}�'zb&��OMn�ht�ʢ:�\kG���Rd�O�a�'�h6�U�@�
���H�.#�H���;TD��'Y�q�S(^��ܫ���D�ߖ8��F��PƋ�DjIBC�W���{F������	��G��'�F	� ��]ڙh�T%62�� �'7�;<BT��O�n�D�ӼK���V��ω�m���e ��<!�iP�7m�OTqy7�t�J�f�j���`څw�x�� ���5M[�C�^�Ȅ�о3�2R��+��<ͧ�?y��?���?�K�/��U ��ΖED�)�n@���$�ͦ�"�+�џ���ԟ��r�כl=.�r�
��UR$�n	�?���M�F�iSɧ�O��EBQ�;�vTY +�&���Ӏ��Y��Oh{�f�=_��������c�TL" �[�21�)�RKTS6�D�O���O�4�ʓp�����+�2$ȟU���㍜�{C^�5e�� B��xӰ�dJ�O�lڤ�MS��g�j:j��t�#�%� 1�^������M��O�h��ɽQ�B������w�f\�6&M"��ԑP�4!8�'��"�K4LW�9bW1d��T��'Gb�'�bv�*�q��?���4��I���Ôl�)S.ޱ�0�ߟ3��L>��i' 6=��K��`���Y���w(�:ZW�찷��%]+�٥/C<�&I�����䓾���O\���O����&���c��BЂ��2��m��'�\���޴p]�����?�����.>D��)
*}n�����SK�	0���LƦ�ڴ��S�d̏�a���b�W2n��k,R� ��蚖���pejcR��ӑv�خ�6o�'�B�c��j�����HS'.��̪��',��'�����O�剦�M�',ӎsF	۲��uBLQ'�V�����?���i��OR��'�7m��LH����1n,���b֠mɟ���æU�'$�z7)����FW�,"W�S</�"�B�"X�׺�г�|�̗'h��'��'���'��=a�27��X��"g�ƥ�E+�4�d`@���?�����'�?10��y��Rm����&�
ތ!����3)*7mHЦ�'�b>y5'����̓:��I��X4�=������A͓4� �c�=�NiPJ>�)O�ʓ#�<頌�R�֩�* �.H��	�M��I���?	��?�'�E*׆]B��	3���X1d����'���a՛�u�t�OL��U��3MAXժ:g�8�Ü���0��l[�J��{�ky2��C�����Z�������Q�R��+
�	�b�'@��'������R�D�u��9� n,�=X.��p��4K�\"���?Aa�i[�O�.]�>����ڙHR$�2t�G�Q.�$HɦQ"�O�钤�w���F����u(��w_��pS�O��F�2�h	N+:$@e,Ѯ������O����O���O���2t(������h�����R�9�˓"��
��p��	���%?=���Z�5�'�L#e�`�8��%�`�ȭO� oڽ�ا�OPp�� ��R}�@�f��$�L袏�\��rWS��X���i�h�;w|�'x�3<��욣O@�G�ѻP)�jO`���Xʦ�惆�hń�M��!W#l�Y����H��4��'C6�&$�&*m�2����?�a�8�j)z`��uF�j�KĦ��';�9���R�2�H�{C��t�w��5R��װ=�|��Jׁ\	�ɛ'���'���'���'��F�ٰ�Q<yU��� @��������O���O<�o��u���D9ߴ�� �$�XDa�OLh)s�^8J�,H>)U�i�6=���� y�"��4��7�G޸��Lf(P@"8�h@�� ������O��O���O8cvR�#�i�Z#���D�-����O�ʓ;�v�<��'gR>1`1E�A|���1��(�^m��>?��S�l��4f.�v�|ʟ(�ñ�w86=���6�|4pbkQ90X���X�2��i>�ZbF��f�|�ܞEς�Pu ��ʨM(��'�2�'���U���޴X�B�#`�á;',� u��E�eJѬ�9�?��ۛ��d�u}��y��@���7oz���L(k���!��L}�KS�=�����f��>����S`lyB"ß*@Rё�9�����N��y2T����̟�	ן�����,�OG�ei� 0{čC�Ϟ\T�5�c�f�t���O2���O��?����3/�L�ÑD��c�<Q'��#𛖅`�`�O1����5vӈ��;k��ْ��߼Ũ�A�5E���I*i���yq���`\'�Е����'�f�Sɔ�uG �S��������'��'j�^���ܴ�,r���?�-,�c��OFX` �ED62��R�>aƼi�>b��ڕ��D�t�j�%u��K"� ?A�*өD�ޑ�������q�]wLR�d]�j����P�ԩQ�V�Jj��b�����O~���O$��:ڧ�?q��[�`�m4ON%#�&�AD�T1�?�W�i�$H�D�'���p����]�+�ʽ0�B.���R�� Y'��;�M��i�rD��暟l�R��#\=����6Z���� 8
Mʔ��)Y� m'���'�"�'���'�"�'�5�BU:)���BO���-��\�@��4j�*U���?����'�?��W�FB=��g�j����@���a=����M�T�iɧ�O��*g��!\S6���f�HE����!�"�u��Q���G�ťc x��yR�'��m�tģ�eك7,�"�⁋}!jh�������i>��'�4�D_5
2M˓ �h)�iB��^�AO3��g� ����O2�nZ,��$�>Qr�xG�8 �>��u�N�0���p�l��4U����L�;t�L~*��Kۚ$�g�Q 7��g���/�jϓ�?����?Y���?I���O粽�Vƕ(r�@h�EH'f��yQV^��	�M3q�G�|"��-,���|R.[K�\�B��7
��
�W0�'��6-����@�o�V~RӀ �%rW��7}��XI�/V�2٦h
7� z}d`��)���<i���?1���?�DG"��@���u�������?����d�٦�K��ߟ0����@�Ob�|p�X��8]�4+�8\r��x�O�@�'��7Mۦ�%��'3�`r�Q�	d!M�v@0ɓh7rY���Z���4��5x�.o�%L>��k�S��Hpa (��Yȁ�O<9�i�"|�ӭH*�9s��)X��y.��<���'k�6�*��>���Ħ��#H+q��%�Ј]0h� � �o��M{�JT���ڴ��䑸~�
IxE�5N ��v�>ղ�a��_Ȕ�g9������ON���O��d�O��D�|
d���i���J�9%��1�P��8X��v�B�RK�ǟ,&?-�ɠ�M�;0����l<L���¬8fI��i��7�3��Iҿ�&6-s���EȜ�N\(*)1�s�tP���4�4��RB��Zy��'�F'�hQ8�A۱@5��+ш�>@w2�'
r�'��,�Ms�-�#�?���?Y��I������יz
�Ca�ϒ��'�T�(��֋{���O�@�ϙ�8�4�SF*1��I���Lh����E���#(��@j��� I"��"���$�+���A%.ڏL4��'b�'��ܟ�abÒ\��Q��-�2ڨ�����9�4z����?���iz�O�B���'���X9�;���(8g������4�?��P�M;�O:���GO*3$,!�.Ûh>�e"c[�Q5�	��T�\0�O��|���?���?1��,#����+k�(%1�I���d�Y+O��n��Oc\͔'W�����'+�0���+M XXQ)&HG��2��>i �i�67�(��)W�	��T� �-��Є�ϭL�J���f�K`�.�"]S�狅�u�$?�$�<1�Z�c%��EOv�Z�	s	�?�?����?a���?�'������d^韘B >&�> {��'e6����韀�4��'��/˛&hl�^��D��Є �Ň�0ȄP'���Cj���a�$�9v��	���#7'��>��]�Ķ,A7G::�vͩV�x���ҟH��؟x�	���I~�'ud���+$�����`�Z�mB��?a�&1��o\%��)���%���r`�45����V�ϝ@U@���	�Z���MC����t!6ɛv��<�rn��zn�m�#�]8�pJ�A�Y�`��G�U�xj��%���'a��'��'��)!�j7�ŁS�w3���!�'��R���4�(,Y���?q���i�)>8����D�`i� A���S.�I����J֦�#�4��S��iOh�i3�S >m���a�1��)��;�0E��O�i7�����a��Drr.�_&�0[b��~����?q��?	�S�'��D����!�,Kn(�pc3��i�Q�@alJ���̟S۴��'U��,���jǭEiUPdB�9b��g���r6m�O�e�֤~�z�%�:lRũ�2���s.O���Ҩ�%F���GM��=�V7Ol˓�?y���?���?�����Ӌo"�RE㆚#H�(�a��2XElZ�X�v��I蟀�If�������"N�$9��&T>/<�V �?!(��`gӶ�O1��r7Kw�h��&-��b���t�}�֑߶�'V5���^�3�j%������'�X��w(#*4T9w!AK�zu��'���'�]��:ܴ��;(O��䄆A��ɸ%"��,nJ4�0(6DD� ��OB�lZ��M;I>��`�m��B��"*HQ�E�v~��?M5�) �M�I7�O��q�Խ�&��I�,м�)­�6%Ƣ�2׬�VB���2Y�r��E�����l� ���ɪ�M�h��?Y�0�v�4���B��,Y�t�s�X;hD�
�0O��n���M+��&FPĀ޴���\;y\�qJ�$������y�Tey��Q�y��M�t 6�ı<����72��ٰ#�P*b�H�c��w��ɭ�M�!���?����?Q����_����k'E� R�B�(ee�7���Iț�gdӨ�O1�*؀��&nb��(R�1���M"~H4��P"�<	gƖr����\w%`�O����E�4�X�.�J4��WB`B�P���?1���?���|-O\n�0UL��I2U��P�jK�)F�@�3�K�-�d)�I-�MۋBB�>���iA��j�b�xq��md^�i�C�j�L�!�/ț�M;�O���6�ʢIRĐ�h2����;҂Q>o� �So�>�"��"0O�$�O����O���O��?�H�@@\X[��=	���K�.�ȟ��	�c�4}�b�ϧ�?�r�i��'l�X �N�b9���"\�$�q�|�Bw�f-lz>A����Ǧ��' lA�@�Z U.�y��*M�R� eL�%��]���ۆ'�'��i>Wdӌ���O�Ȣ��Ɣ+K4�J4�8���V��O �d�<W�iG`�!5�'��'��#,t�rĆ�4~S�H��
��M��!�����Mc��i�ɧ�i�1D^xE�	ݬV�����"yh��$��V�<��7����<~�&a��!��'L�Z�S1K¢I�Q���+����'�2�'U��Ob�I�Ms���X� ��sGG?�����D7(v�-OƉn~�9�����Mk��_�f�PtE�A���#�J�����':X�3�i��	4�.�BE!M�걔'D|���(B�W�0�����=$�|���'��I��I֟��	����p�D�� $]ԅ �C!�TY�g,�7���'����?�N~��v��wH��&Sm�v9br$�"!22S�d�Pan�}�)�S�q�X mZ�<� @e��U+����T�I�d�)�2On��#+B��L���0�d�<�Oj`��'��$O$r�x�-n�bJÓ��F!G�5���'g�7e.&��t�.�+6c�yq�OD=�'�"6��Y'��X�'	�b>�����J�1ꂠ'?��ҕhQ>��E���'._z�XwvB�	)�`D[[�@ɺT��4$�
(1��'��'�"�'��>���*���C�� 0s��kŠ-}xM�� �M�fE��?�g6�f�4��¦�0,���j�$�	.b9`�;O<o�#�M������ߴ����1>l��P+A
�\kPB�4'�4��CB >:@Ȃh/�d�<ͧ�?A��?����?!�aE�b�ܹ!c@I�v��eQS�����
Φ5��Kڟ�I�%?�Ɇ}�~0�tC� bЈ�(Ƈ6^%&)��O�o��M�N>�|Z�H�,65���	z���'#�VыV!�A~�NF���bt���%���'3h�Д�LH~�/V"��}��'��'�����dP��{ܴ ؔ�����<�QO�7N~.т�PT�>Ժ�W��f��G}}����nZ͟Ԁ�3���҈�,��D Z�J��n�Q~b��`��Y����-�O1G!�$"�ޔ��;q%p���/�y�'L��'W"�'�r�i,6��+�M	q��}Iqbֲ���O���[ئ=Xq�b>����M�N>�ԧ�#,����Q�p��F1��'Z�6mE֦瓅{P!l�e~R�O=V��eгd�W��ض�>w���0�#� Mj��A�|�S�T��۟t��Ɵ�Ó�W"paP��U�@{�u)B�����Ay�fo��	��<�����P.l2�Ӆ��R�2������Y*�	�����ݴ��S�d��AAܑPfjP�L(��Cy�(��FLg+
���O��'�Z֝���zy��v��]�\���^/D�M ���?Q���?	�Ş���Ѧ���N��Tn�)��B��f�22�.����	ҟl��4��'J0�=0�v��D���ke�Z�#�PњWE F��6M�OB�b��z�p�J��
�mЏT���O�]��U/O���y�����'��	��P�	������4�Ih��m�>�f]Kc���� �R\�*�
7�,a�h�d�O��$:�9OȰoz�i�B��%N,Ȁ(�+@'��
��&�M��i"ɧ�O�����i|�Dǐ=���Wi��뜰�dÒC󤚘)�DJ0	��@��ON˓�?i��H�R���.nX6=��&Y�`���?q���?�+OL�o�!,�A��ߟ��ɋF�Ra�ơ��	�l
�GSiε�?)�Z�`��4y���|��� �0�S�B	؄F����$�X��[d��������kb�	����\i����E��$��L&^x�-����?1��?����h�&���,A�z1�@ZBk�q1�@�.���$����Q�M���	�Mc��w�ME��9����GÛ*Q��'dn6-�����Ix�j�lZz~b	�"�x��P"Q���x�ϱC���F�VYp8���|RY�$���0�I��I��0bw�;9�4a��� g�"0� �ey�Gr�<����O ��O���"���Qt��Ð[�"%)��O�#�^a�'F�6-�Ҧ�%�b>Q��dL�g��I���G�Z��!��$��I6�Ty�
R� w�5�C��M%�ȕ'��� �ܩW �ɆJ�!�8II�L4�Ǝ��r@շ5�}C�	>F�Բ��x�{�"�D��ODmZ��M�;)J���2�FA�N�Ã��ju�����Ms�Oȫ���@� SF9�	��z�ҷJZ&GW�3�@�Wj��<O���Q�Jei�埏G� 0rҍ��L����O�������.5r#�i1�'R��Bq�!gd��g�f	��,��s5�6Ay��
-L��6�7?���V�+o|H��L��)���|������b��Y�N>�.O���s&�t�:��6��J)V��` a���Mv��'g�_>}@A��3ވ����B;�0t� E??�eS�t�شo*�֜|ʟ��,H��p��O�+��!W��Kܖ؋�ɞ�a�n��|*��9�u��/��D�I���1�'�S�r�Pt�,U�!���զ3�)�%r���;Ƣ>D���7`W=3�H�����1�4��'��Ze��jND0�)S,ϐ@ M��J)~��6��O�� T$x��3��Ir'L#��-O��!�-ܫ2��@樂	w�V�8��V�����j�����P�E ��p�֡&��� g��k�&�$�S� ��8�Ŗ�@P+#cK���#g��F5Di������`��ޒ,^nX����6���Ȉ�y�U!"�#P����/[	���')�?epY���b���1P�B�u�z�󐄒X��=�W,^�@T��*�1] � �v�p�b4�X%:q�)k��J�Y�T�s �7pw����F	�v��a"�CGmI�^\��W䜛|��I�f?zȾ����߅:yReQ ᪼ �gV�R� ��c�'jR�'��Oe�	����	?��Z�h.ֶ�1��,�� *ݴ+�f�Fx��	�O2-�3��!'"�SV�V�,���O����Iş��	44��R�O ʓ�?��'�֍#���}_T<��m��/�����4��^]�Q�����'���'��x;!$]&Z�HP�"���>F��yӆ����9[�\�'{�I�$%���r���%�F-�h�mτgb����Y*�����O8�D�Op˓ �n�G·�$~Ll�@fOKb6�	�����Dy�'��ğ\�IП���ϖm�� 욲Yޘ`%�A�t%���	ݟ��IiyB��3��_�Thx(����;��\��n��`���'|b�'�'}r�'lh���O� ĵ�cvlm;G�K�> �U�t�	��X�	yO�:jn�'�?�c/F"�5{�,į9�D	�F�B�R��6�'��'�"�'֊����'����XV��$9�h��,�� z��n�����Imyb��F��?�����\�E��Ts�ջ� �5���H��'"�'mZ��'�'�'���C>p�<{1k�1��l�b��$���W�8����M���?q��BaW�֘�zz�1���KC*je:�P
8�7m�O4��V)H��㟤�}B#bG#v�H�W"Ҿk� Ast(��]�hϟ��	�����?}�'��'
q�"땊Yr���K1z^@Rv�a������)§�?q�*��^'��� $��:���n�)���'B�'d�KͿ>�(O��d�����ưDS�H�T^bԪ��=���q�%������ɺ�\���&F����J�~����4�?�' +����D�'ɧu�X�0���!r�I5B���P�L��ē�?�*O~��O��$�<��� '�p�Ǯ�
'zmԭ˸9
�4�F�x�'3ҝ|X���)Z)(��'����V勶1�6��O�ʓ�?)���?�*Or@��F �|����&(>.��	F>V�^�q�nOs}R�'p|BQ��S՟��D�M�ws�3&Vo��4�
-����O��d�Oj˓H�*��֝�4�]�e�ްAB0s��M�u&�1;�6��OD�Ot��|J����1�j��Qi[7�(�9W�5Zr6��Ol���<�0��ȰM|������Z��P�e�B�Ӹ���D۠/���'�t�'�R�'<��yZwB����Z��͢��[2�����4����٦q۫��$�����'��2!D�g�d��jX$AS�ۦ͖'"�'E�����F�̇U��e؆L�� ��Ը�M����!�?���?y����,O����qB��΍AR��ʃ��3yY&���O��i5�)�'d�T��ӀÒ1���ͦE��`�ƾiW��'er��K��)2K�DqqO/0d����$k�J	��!���O���~��~�[�L�n���gM#W��J5��MC��0�a,O�x�OL�OHeB�G�5	�3��<����WND[�	���b���	^y2�'�,𱗦ǆhzFT��zi��Bʆ|h�	ɟ��IZ��?A�'p��{��<[� �	�;x؅�ٴ����<�����D�O���0�?��g'ɩPfvE:0���U�*�0�`g�����O�����XyB����MS�Ѣlh@b)K�X �цiD��ٟ��'��M�
OX�S��DZD�
*��;��UV����/�MK���'��	�*�PO����C>R��"�� hW���i��T�D�	���O�B�'p�\c��+e 5:Sg�4� �H<a����$Z���]�8@�"B�N�0�1i�d��t��7-�<�#k�_����~2����������=t4Ö��=������d����?��c$�O���MK�BÆs�XHZ6�
�A�h��f��ѡhե�M����?����#�x�O6$�D	Mi��G�'V�`��z����O����Ot����|҅H�yu���M`�`Ի�*�i��V�'�b�'[D��3]��'��	�=a���m_�R��#1ǰH��,!��$Nh�������͟��� 1'OX����O�2t���
�M;��B�v�ia�x�O���'6�I1'�Vpѕɖ�^�X�& V�zAjڴ����O���?����?�+O�X1�,�2D8ى��U�X����� �'��I����'��'���N	.]�A!����0 ����Z�,�����'2�'*R�'c2S���S�
����(&��`#UaL�!V�����MS-O���<Y���?I�l���ΓVL�I�$�H<Fd�v$�%IC��%�i���'���'��	�HK,� ��x�Ē�	ȑ("���r�Г��<�VmZ�t�''��'����yB�>�	��M}�	)B��	\��@�a�ͦ��I�ܔ'`2��%�~���?��'T2(})4܉.�F��2"O�\��� \�p�Iן��	�	F�IU�$�'G�I�_���.C�p	>8���t��fS�� u'���M���?�����^��]�v�J=pO֚A���4�װ�<7��O��D�+y��$1�1�S�0X�ek�!�r;�� �эo�*7�әXbD)l�����I������D�<�쀈WE��1�gϘ.�~	C׀I����T��y|��)�O�ᅯP�9�&�)�g�;~ ƙ������	柀��!e��`�4�?i��?1��?�;kg���đ�*oRj�C�-��o՟0�'�������	�O����O��6lC�*� �3Åܬتd�ߦi�	�xX��O�˓�?).O����L<
�.+Y.p����� F ��P��A�u�$�I��`�	ğ0�	b�ԩ�E`��3�%4��[@��;�@!��oӄ���O:���O��O
�IߟtS��ٗDq� ��X�i�@��@�2�.��П ��ן|��ܟ�O�|��%�eӼ$Z�_)T�E�mV2	� ) �jSƦ-�	��H�	��h�	}y2�'���O�J= ��Ș}n�2W�j= ���At��d�O����O:��O�4K�mw�x���O �`K�$�ؐ�Qń�(h
������m�	ߟ���^y��'e~���OsB�'�$����2��,��վ[E�Xp�l�����O����O2 "�Ϧa�	џ<�I�?��ū^z�K!��V*L!xW��Ms����$�Od5r�2�,���O���� b1�`�E3;�d�2Iqv����ir�'�|h:��nӺ���O����B���O֙!T�27����Cnڧ l���`}r�'�a���'dBY��SC�)I�?P1��ۘ@'Z|��C\�e��&M��-��7��O|�D�O��� z}bS���K�6@	����A\���h����!)��,���O�˓��Oo��w/��r�T*xGH�J�Ɨ���7��OR���O�MD�q}Z�T��R?Y�Knk�̀���&g��V�0a��	uy�`Ԣ��4���d�O��d�D?|�;��8O"�!Wi[/X���n�ϟ苆H��$�<�����Ok�O(!���e������ ���I�$��?���?������H�#`���B.��;�F�<O*\�{�Yi}\�<��vy�'���'d^�B���rӀ�@Q��/Fs�E��y��'Wr�'O��'��8;���
�O+�M�v
F�4�C�L��k� �޴���O���?I���?9���<��C~� ��������"��2�� o֟�	�����TyBD�~��'�?��B��@���+/�1A����n🼕'	��'�"�J7�yP��r�&	*0 zjE9	�,|R5	��Mk��?!/O��C���U�S���*��@X��ڟT7�	�g͎S��̉K<���?��NՍ�?�K>�O�nIX�,W�B��B���P��83۴������nZ=��	�O���Qh~bSD0rm;�R%k�P5u�<�M��?����>�?�O>����K�(Zz��s�,�#w&0
b�[��M�p��m�F�'���'��4�-��OL����%un�D���D9{`�Gi��QC7*���O�b�Bj�b�����o�"7��OT���O^ ���c��ğ8�	{?��%2ٓ2b�,;�eJ���ڦ�$��@b�ʻ��'�?����?A�W5jڜ�e˗�Q� u���Mf�v�'g�eK�%3��O�d)���\AG��'!B�����z?�S�_�da&��ǟؗ'���'+r_�\P�����:6�b� p��M|R�A�I<��?	J>	���?�Q ��V���3�9VKD�R�b�"D�P�c�����O����O��[�C?��A�B��6jq,���Ɇ�&��+śx��'\�'���'�x-i�'\h�r@	Q�GM�|-R�L-K��F���	ҟ|��Ɵh�'�(�P`F1�",�BDAf��=��� K�O��YnП�'���IП�p~�`�O �Q�/	�V���H`HO;Dbr�H��i�R�'�	�U�̈�O|b��Ҥ���jx��xPA��y��,�`�De��'�b�'Q�8�@�d�?�A�lD6�R	�qL�r֬�ȗm{Ӟ˓B��S�i���?	�'F��I�u����P�Q�7�p�Gꗬ5W�7�OH��ֶ+�J��*��&��k>Pu2a!�h�p1۵擴8A@7�})d�l䟨�	П`�����'9Pq�4/��0�Й����%R<��m�*��s��O��O��?��I�1j����ڷqd�	
Af
�{��H�ڴ�?���?!��W�'�R�';�D,=<���vfȅ1!"�r� ����|�MR3( ^����O~�������	Q�Sa
�!$�U�'�67-�O~P�*�A���x�Ib�i�Mr�	P%w�\x�e����à��>A�� ��?a/O<���O����<)�cR�,������
8ld�9s-S">��
��xR�'�|B�'�M�7n'\�1�@ߥJ���+Y�D},(f�'
���	ş,�'��2T�b>�(�i�x*�ؖ	��+�v�Y���>1��?�M>9���?i��!�?����#2B��B�ב���ˎ0���ן��	����'D�lC�O=�i��(:�(Cf":DXvM�f�����oZΟ �'��'8�ɝ���>i��́Gu�T����8�R������	ܟ$�'�z��Ո ��O����*��TL��w6�g_� �������<1����u��S�J��\��i�ga��' ��mly����7-�[���'��D�=?1@f�*P"$�րT�w�քKt��c}Q����b�S�ӳ$s��葆��� 2�ـ8��6��#/2���O��O��i�Ob�D�|���w�96�E*/RhuKI!C��	~Ь"<�|���bd4��8Bda��Q��Pz��i8�''򩓁M�~O���O��$�8��I�-څF�5X��H n��l�>��b̓�?����?)���4�xJ�6�H���Mx�'-�Ḧ�'8B�~b���4�.�A !�=vp�1%�ϐ0NQ�x��� ���O����O��6�^Qb��sx��D��]F^2�&*��'�r�'D�'�b�'F]#`K� ��F*�N�<��CH���'�"�'"_� �%��������$�#W�^,i&�A�,���?H>���?��#�K}�⟶'$M�7�	'0Q<�y���9��d�Ol���O�˓;^H�3����Ɋ8�~<@�;��������|{7M�O"�O��d�O�����X
F�S�[�� �R�A"Q#���'gb[�2t�	��ħ�?�'P
�����y�V�%�'"ꙹ��x2�'ErK��O�S:�,]Rk�p��-X!�Ag,6m�<��	N�f¢~����"��� �eǶ �0 �&G�D��dv����OD�Rc�)�S�`�ҝR 
�`�b=��gE�.��6�`�Mm���I� ����'�҉��(�Z!b"�-H.�W%j� 1D�d���?�U� �<+�蛷r"�� i�4C�����idB�' "��� Dc����L?�ŉS�B� �qrj׵3X�ʄog��T��<����?Q��N��a���R1E����VQ�@qZ��i��HT*�Db���	l�i�����
u��,�#Õ�4^�%�>��[D��?���?�(Opi��]�@Wz%�`,/0�=Uǟ�O/(8�>������?���#Nvɹ���<8یm@��؜n���2@W̓�?Q���?�+Or�� F�|⣅�<>����G$8�0 E��v}b�'_ҕ|r�'^r�B���2��9�ÄQ����d�	d�������	�$�';����~
�2@غ�5h�4WM�<4�I�iv�W��	����I: ���	@�D��9S�)���&||���̤��F�'��Q��!)�&��I�O<����L��UqHR�q�) =t�Z- @�a}��' ��'��i��'�"�'�՟�P���Do��Pӱ́� �i��ɯ:Nʤ
ش�?����?��(�i��;���bn�l;KZ,Ƞ�{5�o����Ox��6O,�Of�>�0�!!e�"xr4���ؗ�m�Jt`WL�Ħ=�I�`�I�?I��Ol�� �� ��!"�E�歅P"�P��imɜ'��R�|���-Ҋ�8���R��`L �~B,�i���'UB�����O��	:/�\�X�)�9�bmx���D7�=��=('�?���\��:WB�)Z�f������0oܙcߴ�?��8���{y�'�����6M��`�@�	P����ڎ~���2Xx�̓�?���?a��?A,O(Q:Qc�4���لCĝ.ZJ�:����':FA�')�	ǟ��'(B�'���W�x��#��Z��D��B�tH	�'���Ɵ����'�z�C��t>��GƮNx=:��J<ˮ�ؕ
r�x˓�?�.Oz�$�O���E����/�%�/^�I�\���L�U\��m�,��ڟ\��[yR�־r��꧲?I��Ύ�j�bA���I�n�P��;V���'?��ڟ��I۟�8#mv����Ms�4��-Xa�K�&�3�WЦI�	����'�Z���c�~R��?��c�ĥ�$H�4zr�� $CE�d��M0�X���I�� ���V9��	��'e��ߍTX^X ���
b��C잪t��Z����*A��M����?)��jA\��ݺ=0���&�_�+[���E&T�b7-�O�������Ly���/'B�l�'�ñ��A�)@,����
Z"6M�OF���O(�I�D}�Z���	H�:L�)۽B�$I�D���I�6�NMV��5��?�SȟЪ#j�5��5
&�L7���s��)�MS���?��3�����]�4�'��O0P�� ŧr�R�{���|uɪ��i�B^�`8��~��'�?���?�� κ~��񠬘.3(�9��L�?ț��'�δ��i�>)O����<��+3�ÀB;F5�`�	���@p� �����	4�x��_y��'���'~��'y��>"lP����"�3T� ̮9-OL�d�OB�d6�D�O@��6`��E�#.E�2�4	Y� K��6-���I͟��	����'Vb�p�a>1"�e�*46�STC� :��tǎ�>a���?�����']������a�D�.����Bt�>Lr�_����˟4���4��e���O��@I�[8¼�1�$���)a��J�t6-�O&�O��<q�	�v�	�.�1W���e�� ��g�b�7M�O,�D�<i���r������I�?u�W었K�86'��^��@C�3����O��$�O(��8O���?a�O�ʅQQHŲ 턄��7=�Ҝ��4��D�g\�mٟ�������5����>��"�DQzd�t��&c$�1�iQ��'��(�'E2U�P�}g(J�� K'	�	I�LLɗn�צ�	ES��M����?�����\���'jؓD� \S�9I�&"c���/m��e�'b2�'ur�	�Oz ��H��)�6�3þz��J��ۦ����d���@ k�O6��?��'�b���.�+"V9D���p�צ��I�,�ɦ~Y��)���?9��V26�R���/w\��aN���0��i�2L�l�>���D�O*˓�?��c��a���t��L����l~�Xoן�!�y����՟��	ڟ��Iiy�~���j���<���[f+@љW�>a(O��Ħ<i���?Y�>�\{��L�c��آ�3k��x�D#��<y��?Y��?Y���
�����'F�VhXb�N`Z�j�úY�TlHyb�'�Iȟ�������j��� &C�H�y�'��N}�`�g�(�M����?q���?-Oڍ�`F�g���'ZF�q��J+���W����C�P��<���?I��,�2�̓��i�l���C2{u2���bb�:�0ߴ�?i����Dܒm��Q�O��'~�$��Q� K�iV3R����V&���?I���?�W��<�,��?](v�إT}��)��,֐��amӬ�*�|XI��iU��'|��Oѐ�Ӻ��k�!D��[d�M�d�5�����	��� ��g�$&���}��`�.��P�F?	a,�����9xF���M���?���"CQ�X�'���f��8b~a��j�z�x1��m�Z��6OB���On�D-���Y窕�q��S�AI���j����M����?��d�� �WT���'��O���ύ#@# y�愆5U��=I�i��'�*�3�����O����O������gdLʇ�[7ɒ�)�!ZǦ���+����O�˓�?�)O���Ƣ<��'��:�/�F<pA��Q���T�s�(�����vr��AL<�{�? � �1e� K�^�c�HǾt3B%��"O݋㇜�+|�tС���\7&���	>�lI���8|������ƑA#I��Pv61)w�D�>V�EH���6����$��d[btH#D_�:'P8��K��|.�Q���I�
>�	0��(,�LihWF���	㑪#Qi!i�>Y�	��;�R-�����>�K�M]�;��|#�['��X�n\�2$��"��9~�a�i�V.�#H����#�'�2�'��A��� �/�QQ��F!�5�@�6��$����5�()����U�,�"J�A�'ԐC/]@�����Z1x�D�v�:������(&
�)V Q�}���x��H|�'M�����?I��?I(��u���))�铌u9:�H�N�Od�"~�kQn�(�C��M0@R�aۈ0����I=�M+��?�IM�Ut<u�,M6L�F�;%��<1ԁؾiA���'��Q>Yp�Z�@�	՟H�ԦU&��Ѱ�Y����A#��e���2Ξ�
a��>-^H��7�Y�(�p��|�](�*� P)!&8���N�;N�%�C�1eBY���X�@�П'u�ic@�=���؈ e8WQ��A]ҸpVmA	R��O��S�Q�I(��y�%ؤ\_L����Gx>B�5`�(u��EƠy��r��4)�"<i��i>]�I�N����Aϗ��BV癬I	 �	؟`@�q*���	�h�	�Zw�B�'ҨC(0�1����Xr�dƁ:ꄪS \#o�fx�������8����<	�$M�,F�I�I�-Ecji���̚'(Ұy1��z���+W���9��'l ���2扮 %@�ّ%�F��dc�)ɸ/� �	-a��d�O��=�.O��&�1[L�Qv&V:6Dhxd"Oډ�@��"�`��+V+���ABW���D�'�	�%?��4c�2x�@�өw 8�CЇ9d��9���?���?yʓ�?�����4�ݜ���+<��@ʥ�bHکi��F�o���k� �u����bЂL��lDyR�Ɲ]�$y��=VbX��S���M�PAz�m��*��� �@>�h��X�-��ADy�?!�?PD�yĪ�'�ȪD_#�r��ȓ~51��6r�VL���Q�A��+��M��`Z�],����ɐD�r��򛦛|�'���?�-���Z�ׅQ�����&�0Y(Ĥ��ɜ#�h���O��D����PQO[�A�d}у�W+Y]0��OҌ�h�(�F�-��1�c%d�u�	`ն(I�o˳=��9���>w�(if�u����%erM��^5J�ބ�剩 ~���O��?1�S��"P ���*�@�����n�p��mx��Q�͑EE𬉧a�L����!�,�OR�%�DK��W�cL��Ï
�%z^����p�X�]9�M����?i/��M��O��$�Ot1ӕ�� #�|�&%�`�M{ Eգj���o	&p�f���2%����К�~b>�N�]5�H��X�E�m*�d�4:4ѩ�A�qh!�q@�bm�����jT��w��w2XI���B�	[!f¦i`�8!��$^�p�tDl�ڟ�D���i�Jk��٦� �
�NR=̓�?�	�݆��7jP�g^T�a��*:��Gx�(?ғ6����j��őV�Z�M"L$�ק:0��r��?���Ru�I����?����?�����$�O`����Z0P7:9c�ՁĨh���Y=@����	0��)�(ƞ���г-��<0�y" ��(z�a4�\�L�� H�.lL� �`]6G�I�f�DdB���O�n�;e�Gn�TZ�!Sl۲k�<��-�9!צI�aߖM�IW����i%{$�"�R�p��%�0�<D�H;W"�X��$²�N�l��A�&N�HO�)-�d�a��oZ�s�r `��_Ѯ��6G\�x����	���	ȟ�:"*��$���|z��ѳ�6�D�Ϭp5l�2�IU>и&��0ttk��R�q�=j�g_m��<iW�W,ET�җ�cF�@�`H���H���k�@3�Y�"� ;�^c⭈�8�:�<�#�ğ���A4�Pe�G�5À\�햜J\����ԗ'���?��PhT�&�J��,ZH��w0D���@�ڍZ��"Ң�g1btp
m� Sڴ�?1����z%F��"�ަ[+paI R�s!��ٿl��D��WN�&�{���z�!�䚎0s���C�#Rg��	�ӯy�!��Z82�n�j"�n-�9�w�0�!�D7o��Ҍ�hȆub#d��I�!�+(͊y��b��h�L�I�a,5�!��Z�x*������;�&��ÑI�!�Ȝ;�X��!"մ9���#嘵f�!��]+*d�X6�Q�kr�e��D�� �!�]̊�"��[g��S7���!_!��2"q�Q���?���
'�$KK!��4�԰� ��mP�H1�Ŷ|3!�ĕ%{,��A�{6$��'*<j&!��%_FtBF���7-�쉆ȕ�y!�� l��0��<(�~L��<S$<|�"O�t.�!4���2��.H �"O@�� b�ri�:�H5`%"O�X!�FNUz�bL�n	hŊ�"O�T�#�2j��Q2���#����"O|\��Z�c�$]:�&�!�P1²"OJit�Ƹ}t��Xv%����t"O��K@�L"u֜΍MJa`�"O����[�Ƞ#.1Rh�G"O���.��"��=9g�#uT�Sr"O��Y1Q�Y!����`�j���Y�"OD�9V��>�h�����!h�p"O��	�@�EMj�*�O#3XHRB"O&���.O�y�PҠ��$�|pR�"O��agʥ*��aÊU�@��yk4"O�P�ê�>�"�㑤϶]�8x�u"Ol�`f�N� �2��"�R�X "O Z��%fd:�P�bɤz|Z%"O����6����U ъ �u:�"O�Y�M�-Kaxi���'�M�%"O�h�V�USװ���@�O�B�8B"Oj`CŃ�4u��8+��\������"O�S(��-n0�� ���@"O�T�phU�!z�頄B�
i�P�4"OV�P� K)P3�1�a��b� њ�"OVY��Q�@V�hC+I3w���"O||Z��i��Sw�ҫl�"�a�"O�'LF�eQT��d�X�u�����"O�T��ŀ�M��P �-�f�� {"O$��'C��`2
�J2��Ss
��"O�E8��F~ F�� @T�c?,t��"O2�b��ۡq�ty� �q�((@"O0`S�,J�A��#!�5j؂�"O�-��MhS�uQBbMQ["Ђ�����)xa�>�O���qd�2���{��Ϗz���3�c�1���a�N����跮�<�p=�CÁ�H�r���l8B�����8<b���"�O*2ъ�ϰ}�mh���~Rk�	ECJՀ�Oƃde̐:u��0�y��R�Va�����]�РY���S� �jun$O 88���Ahh	{5]?yF���4f�A!B�O�),^<QD����p=�o�G�+҄<z�N	�.�T�'�]�%�(��Mɡc��@��Iԑ����CO��S�?:��ص!ϢR���-̐Vu��O�%�A[�%���%��?I9�Nٝ28~isHG�`]l�Y�#r��i�$5�dDIV�'LO�L �R�vb�\ˆ�A/M"�AB�H��ēZ�Tx�@0�3��D[�\!��=9D�GO׸K��$��Ze�D�N�^�d40p��>s�<�ЦNd���I��h��	t�
x�1hܾU���-L/��k`��b��!&ZT�s��< T��!l]!!�$�0)�����*���9� Ô\��P4~�)�@�-����O������qڀE*���8�};�'�0c2�W�oqZ�	�m�����5�s��<E� ��A��|rmZ�,��A��?M���^
��x�&J7e!����kJ��ƼC2�Κt��
.��~�:v�
CŌ�.����vi�:�p=q#�ʤyg��}�ɛqcQ#U	i�e�D�"����)��<)eA�	qZx�7ƌ(���Ϗk�a}���g�4�Z�S�$�3T���hv៥WtP�g�'��8���o����M��d��U���6(�F�v@+�	V+�$"�T���l,V9��H��!�r)Ї����ABӈ؟
x�'L(��k*�j 'ب{`Z������u���A�yr\+^��Bn_u��^P�'�l����TW�M��kR���=�ȓ<��b�ڧe�DL&GR���E�@�h֮|��HADDar ��4��J~�'�8�-D8�4h�PŖ//�<9�F�X�J>��癁h�t H��6��d��$O���2B�T!
�b']����$� &ԶS��ʒw��!)C��q�I3+�ް����4�!X?Y��d�H5�fT� �q����y��� %$�;*��
�)�|��I�<ގ|�u�D�i��ϵ <�$���؇!��Dd�|K@H`}b������K"Z��n�9ު��t��(�ʑѓ�դU��c�X^&�ɲC�V�bY�4Z�b����`�(3t�!PB��@�E����/1,D��p�����VH�{���-y(�P��B�¢?�c�ɃZ7���oP=D�
���*g&���Ϛv� �[�j@�_~��I� ���k3И%+U��퇞j�&�>ق�N%jG��&��9v����Dy�f��R����C�W���a�W�ʱ�(Ofl���Ǉtj$$�� �Ø�@nֆx�~}J��5��� 蚀Q�.��Lߊa�0[��M���2OVA��h�U�`HQ�A���Ǡ�]1� n&�OfU�d@(��Jw�#Ƥ�P%��K�=�ԑ9-�\B��רq�:U�$��r?��_�`�#��),`��®��'���Z�~�@�
F�jlj��� �$�0�#�Aj\�AVHENM��+��P�΅:$Te3��Ĥ@$�>	�䘩aA�(p&�όZ�4�A ���<̙"'��ͪ�@S>Dp��dGL">�#J�FK�@��H�9��u���~"��b��:�O�i@�BY�3�H&��*X�(rÍ&��$��*V���λI��RAn��RCh�80ߧ
ɶA���<_�%� iB,�]��L�>/�zLS+1PX��I�5�5���+u��B\'TV��	��J`!��@
Z(t#��TuX�<AQ��qn�a"��P*�t	!��8�X墔m����	��AZ8�Y�
J�@�$�DI
1 ���C�e+��
�G�!-0Q��bbJC�{�4�����V���Rg�@Ff�U��B�,P]i�`H5��`fBS�;j4���$�J	�)�(žK풽�"EE�u�B񨐈��p?1QǞ�W�^�S��ؾN��a��C�S��8{���,���Lf�' �p�wN�iS�LH�0a�Ր�B�,t��9�%�'��A�C�8~hP�@�G���`U6}(ՇE�vGў��	g;$��L�� �J�c����x(���0������o4���$�	�?l��LX~B�����Њ��^P�J��Ǆ�ap��M�s����Ѣ�*�?ʀ<�Ѕ;áK\���Ì�|�'�2L���ٯB��e�L��
&�4\��y'Hƈ=�� �0i�p 2M���ɏS���a �$�k���7��)��X ��(;�R����.�p?a�\�c<�HQǗ���z�L%@e;�g�1��\��N���Q��y�\F�@d��_!�f��dd�
�`��j�B�����$�Oav��G=!ž�"�ȥ8�t�Bdȹi~�P�<A�� �؅S��u�Flؙ)�~�I%q��J��KK�h*�J	$i�#<�"a��.*��"D!�4W���P �2R&�S�X�H�A��Z����k��$����X����ο>0�@h��X�!Q�@���N�M0A���2I� ��j|��r
!$al��1 ��H�HA����!a�_~��^�P��Кu���,R�N�]<D�
�`�9�~fQRV�X	!�	6��R�T�6�R!K�=�f.ɖqJ�I0
X#�3I6��T�3�y!?�nq�b˂�<�k�ɚ�p>�%��d��E��#	�9j��v��U�5j��C�Bc�T�1b��c��$De���)|��>QA*T���1�E�Z�q��`�+�R%hH<�vc�<��I�����#�[��P��C���S�A^��ų�����.��%��䂵�I[;9[��2O��DS�M���QSkQ�^5XwEF.E, ��4J�15T���E�5�d�P�
B�	#���}R��^{���0f�+�����f̭��	�5�x}�F�'0��	^�D�Cb��/$V��A-��Ra�1BD4�V)�Fj(�(O�D%��Q��]�� ڇ��{R��EL#G�OB��'EM!O�5�����33,���FD)hU�sQ,<Y�>A�%�̱G��:Q�1�Q�}�I�arD)h!�]k�y��$�C���Z�G����F�V�O�*ӱ��k�"1x�"H�!�D�@
�K*����C�9�%�aV N�����J����a�Abx���I�?�Bq�1�U�A��m�Q�&�d�������B�]��4��OC��OZ(�b���V����iɨZ�lՒ��54��0�NN��dI��,?�Ԡ'C��I3���ଞʎ�O��բ#Kaމꂪ�7i������;P:^��S�=$��hC�t���Jr�ͮw�2�C1�M���'2�A5�]�`�$�I� يdG��x�y��GB��HS�#7`w����-��<���W.@����"�V��	�>�jBj	��p�Rኗ(_�!��S+�f]������D��4r�'XD ��Z�<�`T�S9T} [�Z'��q��97p�B�I6��P1����aZ�C���^%�EbgbuܓRN�>�f.Шcb�L1{������uYN<�ȓ%xe���4��5 '��.WXl�4����'CD�y��̾]z�lɘTJh��ۓϐ,�B�<	F�B�X�PȦ�U�ҍ2B��V�<���njBE�F �K����G�<t�!��'��*��F$�T�Ճ�n�55�2��S�? 4�����[�&I��\�%h���DS�I��pj��Y�TS����S_$��Nŵ(\-�u@$D���uL�:O*�j�m� E�t̎�7�ը����>���
~o�5�!�Yq<z�'d�[����$�^=����O��(�_�ed���b��?BrXŪ'"O��� �'�ȁ׫�<V�V�:��;V�8��ި�$�Ïԃ����}�n��"ON�B�*�=�P��� K6�H$Kg��$)@�O��J�� �g~�M,j����C��iA�Ɉ�a͆�y�M� ٸ�Qa�5Rv0�F\�{��E��>U:P��zE،`i�~�~�6#ʷw����d�,?�\����~򥍭W���@*��PA ]B2���y��Ɍ��9���C���Ba �ʸ'�b�2��%ϑ?��dB��(}*�S�������`o;D�p���t�p�Z���r���ħ4D��Tl&Y ��C�+/&��0D�t���ˋ�|i1��e1b؊�;D��)%�Z^�5!�M\+t�����:D�&Y�##jA�A�9]� �)7�6D��C��)���ԃ� SV\���2D���c�ˈz�vL����% �l3��0D���(@(:��h6��><�(�	"D���	۶ub\�q�c\/���?D�|d�A2~rvy�-V&$$�B1D�Tt���@, ́@A��~���@=D�)FI�s� AAA�l��6,۵�!�dB�9��)Jƫ�rX��M��4�!�D�
0p�\��`�6W�@a���{b!򄓸 H�'
d]�{��ѳE!�$B?3=�`�`왡Q/%��h�L=!��U
I=��0���9��}a�A�AE!�d��yq����,�ڙ��H�'!�$Ŭ �<L
W��DP��C�n���!��_2u�
����B�s���+S-���!�dE�un��F C�X����b��T�!��?,Tk��@!?e|�E�p�!�Dr�zEBD�V�eOD�g�W�x�!�dފx��D�W`ās��i��L�!��
�a�x�{�&�	%�t!Tj
=0!!��#d���˦E���ɜ�X�!�DU	Edr�9W�P�=�� �ǂ��!�d�%���,�61�ĝ5!�ć�yk���C�d���Hi_S!�֎=�����㄂t@�h	A(��
�!�$S!1�@qe)t@:=AG����!��:ND����ގp�B�+c�8)!���� �d�Z�N�r���B�k!�䟽tD���"W���5A���\`!��PP�e����8v�h
�`x�!�A)N�Xd�s����pdi��c�!�$�
Zj�A��9����#�!�]<S����$���@8|0!�$��?���e�ME^z��TMߕ_3!��V���1�,�e�dF�V@Y��Q@�j�I^�C�8�j�+3�8�ȓ_���	Z75��\P�
�s��t�ȓlҘ(7�����ˣ��+�؍����|*�B6|(9qFKK�*64̈́�Vs��Cѷdզ}x��=2l���ȓZ��P�.��^{ިY�C�%L(�ȓ Ql����	�6H���1��d��B�(u���R�#҄����7��1��MW������#j��s�ȭ�͆�m�N4�U�	�|��8
v#Y�g9�T��S�? R�yt�űAw�}q%aյOkr�C�"O*TCt�����1�ic^Q"O ]B0b�5\ ;D��]~f���"O�\�̕(A%~Yk�ҁRO&ĺ4"O4���O�3K��p��5#Z1��"O>�c�ؑ0��=�ba6�~�h�"O@1�eN��U�*����Hy"O� ʐ�ɫwr�	D���V��I�d"On��"�(�4��S�Xo�]3"Oe�A�1!T��F��
D4Dđ�"O��� �=~��Q�L�9�tD �"O,쐒��0���Y�#�7{��"O��Z %�C���Q��2kk���G"Ob}�3����L5iVTdJ�"O��ׅ�� �'6E="O�S���6@"wL1�#�}g!�Dڎ����&@�TT�0
��[�!�D�2@�����X�I�x��	;�!�ZĲ�p��ۄu�EJ6�]*�!��+�zAQ�m�CϨ�Y��O�!�-[y>x�a↵��-�B�os!��(qy*P�n�X�1��k	!�$؋oYX9��ь���X�dD'+ !�Ĉ'���"׬�"�ԆW!�[	miu��^֒yB��T<�!�ݷTZp�oAl ���<�!��W�dOXa�B Îe8�fP��!�ГVkz�0�A�Rd�'D��bv!�D�U���1P�#gdY�7�	x�!�J3myܩk��=L.U�6+�0�!�d��$w8���i�K<V�����	[�!�Y06�be�&�^�F$&]�A�86!��
�#'�10��mT�� ��~~!�䚥�`��`��v�p6�]n~!�ڈ	"��f���4
��ۗv�!�ۿr#�dY���(s�Lh�cgͰ-�qOH�=%?}�a�φ��}�6�W6'!�l��D/D�0�7��5g�ҐK�dצg�L��	.D�ؚv!`��Dz+J�9,� т�?D��A 	�1�<��ԯ��@�6kO=�Op�5Mj!�DgU�K�)b��O�Z���6� |���˪q(4��' -%4�Ȇ�F���b���HX��J�wY�=�ȓfy�T�J�3EL�Zb��)�~T�ȓD(Y�� ��� ��&9��,�ȓ*2̃��@�hld���T�N��MM���p'"0�hL��.�E"�H�ȓ>�F4%�V�TQ�̐�|�@��&��q�J	�y�&��SO�2I��؆ȓb���㡉�b�
���B�RA�8�ȓq�NjM
�6�H  �ޒ{<�5�ȓ4���dE)r����ˌ$(�xa�ȓVzɆ(�N�
gP2�j}�ȓP�����O�ihX*3��#"ن�^���xC���N=*3�Rn�(�"O�� ��,I�B�LD6K�"O�l;@�M ,	���m�`1D��"OF�+�f=��C�cŰO��lY�"O��QL� x�F� �>�RF"O1:�A�^�"�r2m��j�X��"O��pE�� !���"��T�N�Z�Ж"O�cAL��^n�:%�W�_��b�"O��K�BE�IHzE+���?w\Sa"O�H�q �dx�;b ۞sjZ�"O� ��Ae�z�f%j�@	2<Tp���"O��]�H1P!g-�a�bA��"O��C�<zz8�R-E/}��Y�"Ot���,	�i��Ϟl�N��"O�	#�*��.�z���I��@H��"O�	�p(Ρ=�(I
�J�V4p��c"ON��Պ9��B&��k���r��5�S��Q��@��R�PbtՉ�gnC�	��:��4ƽT�h<��(G-�
C�	�Q�B�au��2 ��*�FИc�B�I�x��d6)�7)�fّcӾB��B�	"Y��J�	�"��L��C[X B�I�H�9B�nX�V�άR�ǚ� /�C�	�m���O�=3�dp�Z���C�	�[������sc��3����Iy
B�I"3�;�#ɑ�)ӥoͮk��C�I�fR3�ާn��13�
�D��C�I%0��L�2΋�k]�� ��h��C�jR�R�Wu�\��ߤG*�C��9+�|�0�2&�ɡ��[8tC�I�Al�s��[�e�^i�I�yB�ɪ� ��(/*  ؀bE�7��C䉴vt�Y�L-;�)&j��%�"C�	"V�P��O��!>���9_>
C�	#���s�Ee�4X��*�#v�����:}���}?�EB!���ũހ�yB�C��m������*"pKA�y��=�����xYVԚn��y2%,�h�i�m���
��6@T��y�a[�G@Z��z��1P&��y�%����@V���rpʈ"�I���yR	NW(\KP�\j�D@��Ɩ�x���1�^�{���"6A��x�m��B�hSZ��E�/�-p&��adC��$8c��G,D��!�u���oPjB�I>8 =I��%&�^9�ԉ��(jP�	M�����|�TI�_;����<U<
��"O�Њ���8u��1�0S;�TX�"O�����W-`�P�ɔ
/*�-pB"Or�h@3.����iR1z:��W"O�h�q�F-9�̬S����&=��	�"O e)BN�3P��*����P"OVhB�#�,�{�+�6�XcE"O���A�ĜD�x�Z�@P�f��L1G"OR$�`��aJ�S��.,ĐR�"O��S��S C>�<�2��+"�x0�O.���°b�y����;%N�*��2D��t��"��t��-ݘO�>��c�$D����)"戰W`��h�4l�F$D�ؓr.�>����WP+��Z�n<D�S��>�� ��`S3o����0;D�p�TF���4��A�$ b�Q���7D���U蒼[:2d�֎�G�*7gLh�<�GŌ$R^x��fܖa{$�R�p�<���f;�̓�g���n�V�<�`�G����U��'�*��g�z�<�S�߯9�`���B@W�`CUy� �O�hҷ�ܨkV�b�O7n8�"O���5�T�7�hճ��Z�,Vš�"O�	�̮q�]B�5-�2Xr`"O^�1�{�0����Lt���"O"Xa7��_�ܠ#��(&:���"O�$H5)Y�>����)qfU��"OF9��F�RfIr��>hu<4*a"O� �4��H�n+4Pr O�MS>�1&"O����/<��1qJ;wnE:�"O�1��ނ
1<��g	��sq����"O�l�@)(BF��8(�R���"O�=���N8v
�Y�E�O-0���"O���Ȁ<>HDaS��P����"Om��퀖vS�1`
؜-� �1"Ov�0�ώ>�bM��C� J�Rْ&"O�l�Q�.r���� ���"ODŋPhC'a5���Q �Ӿ@y�"Ot��"M+3dE�!B��VŬ��v"O�|S�/t�B��P�y����"Oș&�B2 0�Z�Z�7�ġ�"O�B���1mz�E��jX�"OҹB=�L	)��ϧXxH�"Ol���`B��0�aA�]`�p�"O��j�GA�Q�pIS��G�Б"O=��Y))��
"��a4ty�"O�h��*Ф�p����	�\��"O��j�� �A�u�H�'x���"O���ev�x8���.hh"�"O�c�ᘞ!B �!�^�A��QZ2"O̜Zf�	�py1�$���h�"O2�(S
C�uf!�2��9��"O�H)�e��pH8���	�x��b"O�x1BE%*�Y�(ǉT�H��2"O�d�Ioi����F]�8��`�"O�s���5`�FP �J�,��]��"O�4��k۲cj&���S�%|�M�&"O(�f$W�uqF`	�Hʓ]{t�"O�P���Gp~sd�'\8��"O�A�ы�v�H��B�J�V��Ԙ�"O\�P�Վv�B��Y#5��t��"Ob@ӕ�J'/�P��D�8��B�"O�x��F��@S2�(�(\���A&"O��*@�f��ȩ��R=<��"OFh���< _>�w��[P!�p"O��;��Lz:5C����"!���<�H%N�v�F8�$�Lh!�$�8�@�A :s:�tb�m!�d%TX���O=m\�m�!V�l�!�$ HL�Ff
Ui���bA2I�!��S(]� ]��S>f�tQ2��0Y�!��a�`��%�ؕ)ZИ�e ��f"!���?<�Ɯp���F�@�7 4)!��W�́��:���I7��?!�NH?�a�ƃ(
	�Ϛ6�!��j���Iϥ,��ik�d@��!��Ҩ|��a��o�d��A�"(!�DB Ey ���
�9ch~����D !��}�����!aX�����:�!�02OV�Y��B&OU��i��PyrEŲj$hR���o�p4k�$R$�y��ph@2d\�e�bdp��\��yr��|�@ӕoV$H�x�c����yr�[&b�:	�̅ <|B0K�e���yR��+>&&`X��)P��NP��y�"[�f� $�5zI����%��y�`�c���@ �D�r�T9(���y��T�8t,��c�φu��`�ֈV��y򄊩 �t���K�cNM�Eê�y��K�r����e�$`��������y !
�l(�vC�6]2ze�5�y�-�VT lq�^(ZV�uPT�V5�y
� n��lYg����6��xN�jg"O@PQ�5`8ڙi$��l��݃W"O$y����]p����G�5�"|؁"O�L���<xDl�E#Ζb��,3#"O��p�)�O��@d���;l�e"O��!��R>VQ+�#V�(�"O�  @ C	$a�d��EPб��"O�l�ЌU�9@�dk��C.��"OL��4/�4[QxY��k_�+�	�G"O�mCU��)G[�<�k��kF��"O��A4�C4bn¼AK��7����"OJ�3d̞)e��qJ�.��#�"OZݢC�	p�Z��1تK�%�6"Op��bئd��QL�j�1"O.p�����9��;�μ	"ON(c�a��;\B�{�![S�D�X�"Ot����;_���`J,dAF��"Ol�Fhص`��Y�����V?�a!"Of! ��Oͳ2�D�]��v"ODDò�V,5�ځ:���g��1c�"O��R��]*�ȕ��\8�\8�E"O���Pϐ>��e��$K)Q�L��w"O�����>{��D�MF���9�"O���&;;���Q#���`"OdБM=F�� �Q�Dp&"O�Ź�'�>��r�-@�XEp6"O"`��	xH̹@���.P�Z�"Oxl����j?:�Qe�؛j+� �R"O
�x�FûYAL �uf	�F���"OH�B�I�~�؉`%S�L���4"O"���-ͭ;�JUpPe�Pa� �"O�"g��9aU��FDF�X��Pt"Ojq��#LѾ,J�m�&	|<\�w"O�!ƃ��`x��k�LlD�`"ODl`�m͛dg*�kV���C�H "O��P'�E ���ȑ� =Ȭ�s"Oހ�@Æ�Tnn����Տ:�t�D"O 1c�fܭ&<�b�'$�"9�6"O:]��	r�݉�D��5eؼp""O0jR�YO�� ��8d 5y"O
��AY�Jy(��2H���"O�qC��
YH�<�S�')���"O }��b�".B���Y:4����"OE�F�RϢ���	%�yH�"O��`"@�lVf!�u ��O�,Р"O0MA�B@1e$�1�ϛ�,L"`��"O`l���žb�Ts��א��c~!��MSHbx�d-��Č!�/X!�$G�NUR�3P@A�b���K���9`N!�DG"P�mZ��-w��U�@,!��Rb�*�[�I	V<�`͐�F!�$��)��T��I2F^�k�bB-L%!�D
�	�ZlR�G�3ƶ�hb� #!�$�'X�a�Uǖz��Xz�f��!��Ā�%9��S?|��愳@�!�$M;h���bCԈ�J�8p�!�d�78H��S�+_�hi�䌑-$d!�$��b�V�Kg�#���1���!��Ŵm��D�$̯V��)�a��p4!�d����$��eO�Hy��)��m(!�D�"N��rB�ֽ��2U�P+!�d��y�,�9q��>9�F`�T/@!�DJhH����k�J-z�a،8!�Ĕ!S�b�+wAX�\�Q�n*.!�� �����1ll���(^溥�"O@�Ao�7(�H(2�3�h���"O��x�Kٽa��Bs�©+��!�"Ot���a�Fv<T˵�E�\L��"OeX3�؍�Tb�;B��4"O�@���F�d�6��
]`�9(�"O��`6#��>H�|qW�ʂ�L��u"Oh�#����L-�H`�b
`�0�g"O��l��E�@�R�C�0%�v���"O�P��bԦ<m�y@"F
b���Ȃ"O�јc(�w_�a:��F+Қ��"O��XA��x����V�I&MU�Ի�"O��C��P7찅��Bɘd/�D5"O&`�g�%<z�A!�'|�x�"O`J4 �:d&,ې/��fV�!�"O^p�6�߾��P�.�nB. �!"O�j� u|
!BW�м[&�ܠ�"O^�z�M�g8�y�U�� @�"O���W�Kok$� ��o�R@��"OY'�;
�@TH��q�Έ��"O �s��Ct�YH ��� r���"O�p!�-E�v���+%�^�`^�AB�"OĜ�3�}qfil�8�b��"Opq��ֽ#�d�CCʏ����b�"O�SLV6g�H��&�8^�ʹK`"OJm�f�UT4 \(�� w����'"O��sG��x"��!c��e���!"O��8�a&Xs|��+�@�X�"O�d*T��'���Js^v����"O�
�Q04����l��,y*�9�"O�Qj�
�z�����HYV�y�"O��S�1@k���Ҽj��I�<aA#A)R%;$Ƈ�����ĂE�<�q���j�%�S�V'X��|P0&[}�<ѳ 
*�xr&+T&d���Z@�<��W!o.&}p�¥�~	��%w�<y�K 1=���z2��<2�����b�p�<Ap�ҽuҮp{��;��(�W�[p�<���Խ7�z��3��n��YXwm�<���eN�9�.7+��P�dEk�<�娔�M�$��v+D>=f�8��A�<�CB�4X|�G��#H� @|�<�pÉVb��ƭ�6ލ�Q{�<���R,T�T$�@�:��Vl�s�<DDعT�0�ƈ�u��"�AIr�<��23��zf��R8�!���W�<��%�Qݞ�:�)S�+�\*U�}�<Fi�}pvIx�������K|�<�f��#46�s��M*��Q���_u�<i"�˄P.l�*d�\{�e�%�[G�<�*�� ��hӾH,�|s2%�Z�<iR�JV�fY��>R.,�aS�LZyB�'rd�+��1oh�$`�V�2#��p��$ O�c㓂E�BPjQ�<o �Q��|��'HB�')h5�Ǭǜ^(pX�����!�<+	�'Xe��A�82T�7V:e����'צ@� ���ᳶ�ɶ%���R�'�1�c�ŋ=UT��eoԳ%������y2Ɯ-l)v��7E�t��Q
޴�y2�0Ҭ��Eǎh�Ι�i_�y2�dI�5!#��-�p��s�3�?!L>����~�/�Bt��
�Өy��H�|�<��c]�g�JX��#�:P`]I1z�<1�E]~ѣQ�7=����s�<� �ٗ�
�c�2�+F�9?d~�y0�'��D�hSڨ02aN�N�2\1�ϫ[���)�)lP%z�~�<`�̛?(I.T��'�`��!�g�D�및�!;�Ԣ��hO?U�"d�l��%іG�v)��Bg�<DP�<#��tN� nH���w�c�<q�X�N��`�fMK$J�$��3�Z�<��ȗ!y��k��� [��$͛S�<	0��	��`D��,���q���G�<����1"��h3�h ���z7��W�<A�	��i��h �\�O�� ���m�<�q�
J�`p��&�0Y`C�Mf�<)�Æ*~X�qď1c~��Z�+`�<a�,�9R�E���J�I'h�;%�UZh<�7���t1�DA��x��.��y���7�(\���ίjc`�P�$ű�y���v��Đt*�.\�<������'^ў�_�f;p�j��YQ�5�dQa
�'�!���^")��IV��t�H�
�'��`��>j�&Bc��:C F��
�'}j)��>f�@�/Y:PG��	���d`� �K��%�����g=a����O7��hO��@P�F`W$p�lF$ ���3D��CS��VhuűS�Z ��d.��0|��mq�X��AĆ/�L��eIWx�TEx�L�&1Jt#U�Ӄ�Lh��PyƉE�D!������׊K�<12�O*#�f���S?+���[�@J��̓����ԡ
�t�D�Rc�ؼd����CG�1(��I
Q���:n��I�'wў�|"�+W24C��O�;��@��P�'Ma��.�T՚��Ĉ  	���t�_��hO��iRI��GH7!�&�v��7u!��O�~H�2&��6"�1����!F!��.%�25�b�F�nZŢa^,=!��A6
��!���� WO��C~�Ov�@fVYt�C7NWX�b�|�)^è���Y1M���JB%��C�I*C�8� �ψ2-��a�a�^�P��?	���у/��e!�-L�,����#�3P�!���TLO*wB�0� W�G%�eH�'�Q� �ה2�Up���/y<��'p�1@!$�?��0�U" �}^�)��'}�c��o�8��:}��\8�'(L)�EJO;��!��\0pl���'��l)��ŏ&���p�_�{'��{�'	JcP)г4�eH`B�"	^|���%���`��U2��<ɺ�3��p�<ɵ�˨rԆ�R�!�I���f��C�<i�+��f�=����	nF8}:wje�<����E���Q �~��ЖE`�<��O0��mq��	��K�ąȓ'@��"�-Ln��i��˓D��0�ȓh�4��בk�l�扜$�5��pH�Q��K�w���֏֖��"
�'�D�ЗɴG|naz% ��q	�'�|�4� J�t4Hݣ���8�'��Ɂ5螕_5�塣!^'~��%a�'�΁`�@�6?<���d��'�Lq����'�a�T�G-KN`�qa5�xɺ�
<�hO���i+1�М�か����8Q��2 �!�D�zn*�*��@";�*�T(��gV!�D�t�,��/�o���c��"D)��D\�.�.p��ٺ�0���e��kS �O"��� ��p���<H�-b�HX�>~9��|��)��,/���'#\�W�M0�ӚD���՞V�HL���А8��Y��e��L��'��O��<��΁P�Ψ� �Rk�yj�ˈ��:C�I!��RIR�Rй�d�	�	��B䉩}M64J`��6��a����9[�C�ɕ8���X&�=r�v� �@;V�C�Xw��:`�>G� @�R�B�n
t���{��$��W"�\�d�\2<�f�
�A�O�B�ɐU����֫褑[�Ѷ	R�!��HD@�g��!��3|��Ps�1D���V�:OA�8�㯕�H�H�� .D� 3r	P�, �@c*R=c�� ��/D�� k�k�����9/*Te�&e.D��We��s�j��4�*�!e�+��-�Sܧo�8=��+�:�����k!2\��or$S��
,_�T{���mN���ȓh.��G����:6�L�?��@��D��U�7+�t�WF�G�rx�ȓb�R���k�9��GݐS$����[;��!��L�,
 D�6�A$Jt��� x��-�R�,A�+ "^��'a���eO��8�!B#�����9�'�v����Z�l�X¨�|4��'h�����)f����3�(���'-��ڶ%<^5B#R�ȥu�����'�����HM>(A���dXJ):�'PN��g�KWx��˓�Z�TX�'�h����L$o)\�ȢB��UPJ����hO?ś��\�Mf����^��1cJ^�<1a��j�r8؁M�}����lOW�<9�a� (@�H�f��U��%�P�<a -
����򯂂$���a��'D��@�ؤ-�JE�q	�0e5� �:D�[$P[�@\�sCذ�DC7�9D���Ǥԕ`�l�'�T�1&�����8�O��fg��*1�PH��M�:~$�ȓ9�Di�A�^�g��HC�a�#2� 9�ȓv7�����̍<�tdN� 
)���ȓ2����o_3N���B��� 殕��p�84�U�ٸF|`�#�Z�w�1�ȓ*�,�[�ՊjI�J��Y#&�ї'aa~���=\�j9և��l͋4�Z9��'�ўx���<���\@��AbФ�<>��p�L|�<y�I�	�`X�g�$A��"4��t�<��΀jv�Y�)�h�ظb!JK�<���_,KgvP�nب/��qr�jBP�<��� <e^�y�ʼcS��A�a�v�<!e���!�����S9wِ1J3�l�<	��Y���T3Ď�m����@͉韬�'4ɧ����8�c6K���#�Y�GҾ�"�5D�p����&�m���3r�̱�5D��	�ĉF�)�6��=c �$00D3D���7�>E
h�P()l�tK4�<D�p�RLˈt�&�D�rT֤:��8D�������r�&Q��0�d�1D�t�2IW�D�zs��KffH�A�/D�����e��XK�IV'��0	�O�C���!�JV^*Q��|;�k�	%�p���'�r�$r'��dC��ᘸ��'F��`H�)M��*�m[����	
�'*|�#�ۣV�"3`P�S��	�'0����&��u� 9M�6x#�'��� ���-X���L�$���O� �8K%�uh00�F�Xܥ�"O�- �L�e�f����"gO�(A�"OL���jÈ5�0�c��K3RzP��"O��a��%V�V�0�N+� �B�"O��i�B� o]
#��|�*��?��'�)��/P+���
R�S�c�����'������t���0n�(r�b�'ۚ���'�P���'�$T,$��'��(s�ȍ�Z1*p�N�&m  ��'�p<�Dٕt�`8�
�r*֌��'@�%�!k��!d��
B+�`���	�'�*�:�����VqA1�Q��@�'�0`9�"�}�I��)�����$4�h��Û�%G�гE*3�x���s�lj�=e?�(��@O1E�tx�Ů=D�����œ&-*��Q�ג/�j�)D���sl�3��;��S-I��A��&=D�`�uMC�)|���)~:�Ҋ D�$��FE�x����*j�*5�8D�H�r�YQ#��i �@=Z5��a�c;D���cBsd��H��G_<�P�3D��c���������Iu����)0D�4r�ǌ% V�y���xa�%��,D�CH�?j�`0g�-�v��A8D��䏔\�LT�[�b+b%"�4D�@a�A�LL��@�'N�|���%D�Gf͒G��\��F�@�d�h�.D�L�I�>?����#�I�Q%/D�`ᢪX�L�\�  O "4�|�S�+D�p�
a�L���.]wG���B*D�T�Ч�~^έaAB��J��u(�O)D�L�ס۩k��e�f���p�F'D�H�TL<[�b��g�H�P�
�%D�L����g;la�q� pp��#D��h�L��7�����4Ӫ�	�d#D�,ȓ!L�	K̤1A&R��t��w�?D� ��V�*d��@P��$@&��rDl3D��a�P�,���r��S�C�����h?D�4��$΍)w�I!��C��PE:D��9�AC�L䘜giٔv*���#�O�所 ߂H0!)i��PŕJ=PC�	@����V�RV���jT"?�C�	 �N����72��Ж@P�"{�B�	�ֹz�	^�-�0/�+Z��B�	�x�F}ҷꁋSφ	G�0gp^C��th5�b��p���B�T��B�I4P9z��`L"U�\x�4��>q:�B�I�0��t�'7a��[`��8U�C�I�zj:�s�m �=��Qs�B�ZB�	! J�Y���3yp�@��M{��C�I�F@���	��aR�%��2C䉦�:SBɜR�8��Q�NC䉉dj�#�L՗)�Ҥqp䍹I��B�Z�V ��ˤ'��y3A���B��:�ZppW.�+1���"P�S>�B�:D�H�3#e����u9fB�	�o�=��d=Y6�"�
zB�	5`���u��u�����ċ�#��C�-��Uò��C�1�'Ɗ�l��C���P�� +O���:Y1(���	�'�dQ�݈qx����ĝ���k	���y2�U`i�m����7�08�Q0�yb�X�\ �Р2D�`�����y��b&�X�%�80@�0�ŕ��y
� P͙�� �|PeI��1m��M*U"O�� �%o�^!���e��iqW"OIsюN?^
6�Y ���~e��"ON�a�P+�Ԙ�FGS܄9�'�'Q�0ဤ̥��aP$
�$>���&"O���E�0Nj=�%�*.DY�v"O��i��ؖ�܍X0�GU�%j�"O��P�j����M�BY�{��i&"Op��\�~�i�áf���"ON��V�.��t�ѺHi��
&"O>tQO"prA8UB�U=��"O8h�@"�#H�LX��`C4�i��'YB�� ���6�|�ZiC6VU����5D��C� ��s�X�m�E��T�`'D�|��2Pu��b��3O�&ܑA"D��ҥ\���❊0��d�!D���n̂7ʈ|���\�2:��yV-D�h`�����]p2曑������ D�X�  �@�X�'G	S�iT�<q���"�D���p2��;����3&��0�ȓB9�q���ĪIܢ���	)�Z�ȓ//��JqE��zL�r�!�ȓP�p�p$�������[��X��oƘ�;C(*Y��䅛	]߰i��{@�-�Ӧ��#>�is�R����ȓbܘ��D	9���9�n[�s1�U�'��~	R�'�u*���,�h���Pl�<9qDժ3p�(eYN�b\SeD^�<Qo�F�R�� ��VM3A\�<�$�d��w���z"	\�<y!�ĒM�p�\xd���i�s�<��B@%nޠ�X�/P��	�S[��p�<�Ј]��$M�ԏ}E���YS�' a��� ���=fމh��y"�.|�X���O��H�^ �ybV%�^9jA��C_
5Q��%�y�˲&x���b	4g^Dy�Q#��yBF�4.�B�k��J�-�H��7�]��y������W�מ&3Ҕ�T��y"AY�@ &5�U"�!)��Y��h�8�y2��JdXh��@�q��щ$���y"B��4���0
�.�5�Z���'���,t�-����g�.�zg�.�y"	�(�1��<\�"�����5�y򥂔%q(�@�K� �F�C���y2��/fO�����@&�[U� �y�A��%��)Fڔ$�:�	u�]��hOf���ɯ)�`�z���<I6�U��H	�r�!�d&)�D�c�F�9'>UKc��^�!��>\�l��^:�����&R�!�]�_���$�9�X!���H)W�!�Աf��AهK؅m��yJp�@4$!����á�J>W�y2�!!�V+kH���C�]#X�����?;�'|2�d$执X���5N� a��� K%c�B䉢�(|玗+( � ��ˉ�@,pB�==�v��2 ϕ)���kc#�7zBB䉁��X�w�;&ĕۂQ�I�C��ǌx�v�,J�腐����V�C�IT�^���c�-��A[�*zB��k�
�>Föu��.&C��HLd���G�fՙ��K
\g����6�lU��� HQ���B��d��ȓ�lI��%��p��<�r��8,Z0h��S�? R|:s.O
[�|m*q )Aǲ��2"Ol5��(�)���4��ٸ�"O*`�E�6��4�́�oH�Ç�'��IU~Rj�70��E�p! �^k��"BM��y��M:�bAp�ݿiZ}�QȈ��y��._jd�	�$��(�QFU�yrC�����W��9a@b0��yRNXC��٩Qύ�d��l��U��y�A�y�z%+#,U#_��+dH�3�yr(�c0����P�^�>�
T��!�y�N�1m����c�V�>p � �y�#�!4n �0t� K��qX$���y"�ԡiK�5��	�/;V��ɑ��y���r*�xrc��O�TM�N��y�,X�'�n��BW82�:Q��.���y���94��W��/2�<�ylO*�y�nQ(Q/h3�E<_���	)��<���$Q �]�	�7Z�2I��l\"M-ў��)p���ڳ��,<nZu��Ŋ!5XB�	-X�� ���ud<�a�g���C�I 2J5�V%Ґ"�&U"���~0B�I6�˰�f��pt�?[�C�	�z+�����ԏ�|�qʊ�>ǺC䉨j�����hu���i^�B�ɲ2��t�k�;jvY�-C��C�I�$ (��eՀ8�r�r��B�	�t�T���A �!"�B��?aC��sD���i��lJJN|�B��"}�8�"y��й�f�3?LtB�B�TD0���Obp���X{dB�>
�&t ̌�r����['V�BB䉹)rL�򧋓�d/�90�
ܷb��G{J?�[ӌ��.T�I�We��]ᰱ�ŧ0D���U�!���qt�Ϊ��E�a�8D����枰@#Hm�d�M�fG����e8D�ԋ3��M_rH	�J�&/iz���A7D�����	 �)@�n4/���jE"0D��ȑHƹE&���I��6}��R�E.D�l:V$Ҭ��UJ`���;r�-��N����J
�1-z�H���q��=D� P'�9�fd�fE�&��}���=D�t)�͌$r���Â=u �0��1D���Qc�cT����ߊ?����wo=D�d(	�!�$AF�vi���7D������"��h(��rҀ!D��Q0n)o'z�;�`7E��`��<D���c��}�4M��
ɷa 81�� D�p2#�B�M��4����c `��o!D�bR��.O���s-Y�K���z��4D�l+gO�Oa�9�����Ȣ��4D��+��Ϫ\Ũ��������4D����B�}��}��NșZ����2D�\`�ŉ ��؀���t�ɸ��/D��)6M��!�b���S#V#�t��(D�<�BEP�L3؀���[�tP�*'D���g%�k�|���+kt�c$'D� SWb��� j����h��0F:D��B'h֡F�РK�$��B��-��B�	d�^I�5���;BT���W�C�I�e/��I�KM>���NɉWB䉀{��z�
�L���&[�}8�C�/J�z�B%;��:��Z!rC�I�oNl ���L��ZClZ�N|B�I<Kv2A&l�EZ�<3��Y"�:C�)� T��Ã%;�4���ƈ�8��e �"O�(�P�]�F�t��ʛ&�>Lr�"O�ӗ,s��Q.
�F���1"O Q#6oמ%�d`׋r�Q�"Ol�Q��#s8�q1����qh�"O�xB �&EPpAr ��Ij�"O����j�$'�����_���*�"O������|�@	J���!"O2���dѐm	\4� /��l� �"O��Z���]8�1�.�g�M(�"O0����<a��d0S�z�a"OT��%�S7Yz������@g"OTؚ�"<<���G�:,=,�"O\$���T�l�>e��KЩ2��Y`�"O��`5d�� �٫F���I�v]j&"O~4��h7J|t�8'���yў�4"Op�ض�\(	��zR��1@l|Tr�Q��D{��i�x��2U���|`Z-A��!�āD�E�Q�nNnI�3D�6 !��	;�T��bˋk�@�c�C3^x!�ɭ����AO?!ƚ�A���l\!�@Cג1A2%۬r�I2� H=@!���2<r�*L�I�<P�.��!�D	�qj4���b�0oH�D �Պ}��O����6K~x����_A���D�,�!���-5�L�	�
��*0`���.�!�D�Mh��A3�, M���Hځ*�!�/�������X��,>I�!�J,4��w�ÿ0��H�s� 5!��� ����U�9}�d�z�%�
�!�I$ �5�ӅУh�&���Cg��']a|��<�i�b�!����tL˃�y�������%�	"�(��/A:�y�a�$̱1��GQ�������y��(.��ٱ�ΫP,D0B/ۼ�y2���>t�'��K�TH:殟��y����pk�����FZqFiY��y�kY�Pm� 3��O7=�؄aC���y�B�;.��j���$�):�M�%�y�Z�C8��yp���pO������y"*���-���?]m� ��/��y�
�"�xd��oɖV�����y�Jђt����"�IȄ������yR�]�f}dy��B������y�$G2�2�ҳ������S��	�yb�J�E\4�yv(V%66X�(c���y�oQ�N��Z�h�7"�X�JA`��y�JI+��.U>A@�N��yb�
Vo&\��#�>��9`��ē�y�)&@��[� �19E�-�w�ܠ�yB���w6�����!B��;7Ɣ�yr�AI#��s���¶*��y��Ε[[X`�"�H@\�l�Fi���y��kȭ�bԚ+/u��-\'�Py�.�hMb�x�jS�[n����}�<!2�L�R�J$���AL�J ��r�<�%K)���b��@6;PIRG�n�<�c��&ym��� �?eZl�@ ��k�<!���&L;,s�G�}�E�R%�Q�<�@f�)-uʱ�����L���a�O�<�!@Ā|��5�ք�zp$�!%* a�<�%�6����j�č���VG�<1R��S#�JFo��~m��Qf�J�<�i�}��%�Mj�dmr�oXA�<� �}��oʇn�� 9#���A|d�"O�p7�Ҫ;�pP����P.�84"O@���@�&�Ftv�s�а�s�<���<y)����M�SÌ�"� J�<��N7N����6B	�丂&*�E�<1�9|�4
�gB�^DN�B� �C�<��4@LTq`�T/F�ɐO�Y�<�ggE���Z���$l5��ȓB�h$����	�5�U��8W8����$O�X��D/z���qI���d��ȓ84�La��=b��`٠�|���Z�&ܠ0#N�	p��҅��s��A�ȓD�0@i�ǞDCh�i���v`RX�ȓg�}�Ч�({�4,�@�M*$�ȓ7Ɉ�ұ��U ���[�S�����x9��*޺xG8���Z a��ȓ������u���BE�&�X���x0B@��.\]59J`nY�h���6Z1�WnՕR6*��h>^e��<.Q�%�;e�8�t�K$(�хȓ)��óo»=&��S��!(�Ԑ�ȓ]���0�'���A�t���ȓU�����?Ppz`%\\��Q��^�`��lO*1n^����{R���ȓHm�1���Ӵy1�X?VR��� ,�S��5iNL��@F�W��ɇȓNQƭ�3���9E�ؠ`��ȓX�8uh�wL�.S6-g�1�ȓ��d[��͌3͢���fZZ�a�ȓyd����=�.ԲsG.c�!�ȓt�R��4�ċ�*!�ϕ�C�,����9#�ָ~5H�`b�{�a�ȓ=�
��O,c��Q�Y*8L��
��w�9;#"أ�De�ة�ȓWK��+��U���Kf+Z�6���0���K����p.`��Ja��X��]���e�
�hX�� І#g����t�>�a�%���� :,I#>��ȓx�eHb��Bݙ�A )�����wo���dJS(Qd��0�!m���ȓ~�bճFP�S�"!��(�m�r���JAR����V0N"[Q����䤆ȓ�x�@HL.[~$�a�2O�0	����	���~|8E��D2_�Q��~alm�.J�d;ŀQ �l�LɅ�7�p��p @�%u��3@�V��`0�ȓ#B�p�S�e�dM��D��^䵄ȓ^G�z��V���As�@,?q��ȓ[� m���y�����A+i��m��h���3'��@QX��7�$��,��	M�@z�F='yXE�#3�py�ȓ1O�q��Ãa�:|p�,�]l:(��G�$Y��o�p�-x$Ϫ|�P����P� �átDăVfϽc����ȓ5�@�G�4 r$ɠ?�q�ȓFq5��*�v�ШՂ̷{e4�ȓ^�������'�h��u�_�Ea`�ȓ8�J4��Z*?�!kDȚ>S�q��%yVA���B E�0���
�1�pU�ȓV�|��`�[�Y��tƌ<9�T��Ī�Bj�,(�J� �j�1,�ȓץ!�J�8�p��pH�1Kр*D� �gj2:Lr�2b����)Ig�&D�TRw�L�}��8A!���})�)�4'#D�� �}�f��g�Z��G�>6����S"OP���L���zS���v�v !G"O$�w�i~���`GO�:��W"OMx�&�&.x�/�(Mrb`�b"O<y6�ϓ���s�ǖ'[`�( �"OB�֬��WƸ��� ��T$�A�g"O0(� !O��U0��(��"O�-�"��b� H�j=F�MA�"O��i��"#�$��iG�_Eĥ*�"ODu�4W4- ��D�r�I�"OZ,I��I�H�.4�
�	f�:���"O�KK
����Z�@����Б"ON��Kłu�J��GM�@��A�"O�`q$@ &
��]�!l�z$��""O�H�ЄO!zE�ꒊŏ$xda�"O�L�̀�7i�E��Hm����"O��ffɄd�E��.�=(�ʱI�"O�1T,��3���� �0���S"O0 h��~���r�e� ):Ό��"O�Ts"�	�"QZ�eA�(U�E��"O,䂁��vOp��摳S�Y�c"O�0�0�+B�:a��B�B)F�:b"O�aPP��F}��sa�:Q�*�"OH���B�<Ѧ�\C""O����<a`Lh5���W���d"O�Ue�y*4��	s� ���"Od�åG&_�\l���pP,�q"O�M��*��\ab�<?Z�ݓu"Oj��Aۊ6af�a�1@P؜r�"O����Η�/	���@$fB�2"O�xq`�d%D�I��&`�8"O���BΘ$�>�0ǥ�D]j0"O��yU)�+2��E��oX	!$"O����X�#���r�%��i�����'�0�ta��h	���j@W@tL��'��i�c��I�&�j�şM0p|��'z�ظg(^�*T�)���[�A�Z	�'y0M� ۈB$
<:��F�EH
�'`�t;��^|��A�Ǭ�	mGle;	�'i1f�Mc:�)�j+����'¶�+ȧ0��={n�Tt��'V̊��~���"���
H���'�b�a�+D�<a���{OfhZ�'��}�fôCm�Yy��@6 �,@��']�UංPy��E�-� �(	�'�����J��d�$jQD�*�ε�	�'���f#{j�ɉ!�7-e{�'����(h�8���B��c���[�'�LJ����;(*���P�a����'�&9!�,�YoX�Jt��V"n�(�'Y`�h��%X��U�p� �'?rY��dK1o�y;U˄Y�j���'T|��Q*�u�B֯N!l���'J��94�ԏa��B��ZB2a��'f.���שl0�SeI} y��'��h��"S:\��tS苷-���
�'�r��!�&D����d�*�hp	�'3\=3��0��,�>!�z���'��A���B
 ��m�B�\�
�'�"`�a�A�D�Iw�S?�>���'m�p �a��7�ݾ�x�j�'G~���f��wْ����
 �xչ�'�N��7hH�c1�a�!&B8��'� �兕�	�������|�k	��� jXR���.���p�':,N�1"O6�B�ǔ��d�UG�K�f�S"O�A��N�;��P&'T��t��S"O�y0-Q�mm�I��F�	���J�"O$%S2���:�[s�	 0���K�"OFQ#��E�P��erT�O�j��!�"O��S�G�_�L��@"}{@���"On��p��*����A."ͬ��0"O,����uHleS/A8g�V�a�"O��z�L�&��j��ڠg���"Oj���H_�B�0�+Sxms�"Oz1�!nխ�U��N��#��HA�"OL�$!I+,�����/�6ıt"O�8�� ��"���+]��L"O&h"�`�q� �q���r�h��"O�e�ЎJ;�v5�G��f~���"ODd�ń��S(��/�7B���"Olq���ւ^Z`�o�6AR���f"O
s��X�M����c�F8P���"O�%c�G�+�ܐT�M>CC<<ʕ"O݈1����z�+�G�,A7��"O%Ǥ��ckX��ś���A"O�P���΄`C~`�q$I3zܽ"O���[.v���L��@%|�"O.��Piם\��
�,&&VŊ�"O*L�ƈG�RT)p��`t�iY�"Ox!S� �6Hǘ�)��N6 V���"O=��mˡu$@g�=R@��"Ol�C�� 	Z����B28�L���"O�"�hA~l�挘3{���U"O�� h9#�KȣW h=�"O.�S*��~��XA��F���"O�����iJeeH�^�"h�T"OV�(&"��O�ޜ�fZ�H��@��"O�-�`f�,��i@u�M1G�~�s"OE
6�0m����4Ϟ�Ip"O� �3a�%@v"D��阓 ��jc"O\p2�=';>�P����<c�"O6}r�-���H-�%F��X �"OȜPS�R�\���ۄy�0� �"O֐�ԣ"K�:����R���"O��[d�Lg��q���R�"OҨJe���4���A�4D��6"Or,�R-�,oK�Ի3�F��� d"O*��`��&�;A�r�DUPT"Or)I�I�_���T����@a�"O(x���, �8���F�>��"O����J�J�J7GӺx���5"O�
6�2A�!sG�hR���"O��ѥ0<Q�|�2fJ'TH���E"O�M�Rn�c��3��	A�;�'_����)D}2� @�P�^�VHb
�'��5��d�(��(Ҁk�'cf 0)
�'�4A�E�@(���"�[J�Pp`�'�Ĺ�eN�D��	k�kE��
�'w �QGEA3E<F�q��� :�L��
�'t-���U/C���V.B!��
�'k�Ks-ѕ^db X���77���'��l�S'	;��@rՊ3_�B�Z�'��EAd��Aq�U�DF�J���	�'Ì�9` ��h�T���Ձ4W�i��'H���Wꒀ@_�ˆ�:|C ��'JL�����p5(4�JA�x�'�z�@a�ԩQ��,
��[)@f*����� \�����p'X}�K/8Nvc�"O�$y��YCଘ����,;�"O��:3O޵��Mҁl�����@e"Oh�G��^~fŘ���'��}S4"Ov��Q�� ^�D�k�陆$N�t�"O�p�-Ȭln�� 陨W�p�
b"Ox1à�!"���ٜ �8�z�"O�aAI�9.$I���J�E�l0"O�hS��ƫp��0��$l1�Փ�"Ox �0�ƭ:dI���{�\Q"O�rg�oED�'C3@W@ٻ"O��DnE�B�HcEa� AD&U+"O����n�1��X�j��
/�K "O��g��S.�q'�s2�%��"O�]��ɝ^�z�c�L�X �"Ox��R܈m�|A�I	kN��"OJ��s6�8k	��2���b"OL,٠�J4i�lcBgԝO1�p��"OV��P�ӊ TK�^�!�m�E�<��\�՘(�IF�����E�<!�c�=�d j�&���ܠ� U�<���I 4�a��V�+`�k��}�<�� ޻fr]��@5K����φu�<A����:CxT��Nѱ=*d&�V�<�5&ɷ\���-��0�"�$GY�<�&�vc���Ǉ��pY����PS�<1�ƨ?K ����GE��:�F�Q�<��C�a|��r$�P�cyJ���JF�<����(G�R� ޓ!`�\�7��w�<��ޅ2�޵�$"�p0��g�u�<��.N�{h�1�LR7̀��Q|�<� ��9Ԟ�ˢ��K�r����O�<)5jT2t����&�O֨HeOu�<i�G��pu�t�F� a�	��\k�<i��M�4 Q����R��4�R��g�<@�Zn譋���L�̈�"��a�<Q�d^�Q#�����\N!0E
Ԫ�g�<!�Jֵ�`��+��-[�Y�A@�e�<Y��E�BI��9���4x�I�i�<��+P| �=��CU�,���	Ib�<!��ݳr%�	Z���hB�ԸcI�b�<y�(�$�9CP��&-H��hg�<����S�>ᰘb�]
h���s,����#�39����Nh��C\p�A2h�X�x�Â�*
�ȓN,L�3��
=
����jS�̅ȓ,���0fD�+�d�����8���ȓ3�6RUS�G����fS�9k���ȓ	���e&��"�����O�	N���+U�a ��A!��p�ߧ<�bl��y����'[~� �ju]�e;vx�ȓt�0�A�V�cƈM�$L�bZ����=N$8J��,�jP�s� Vf-�ȓ	J�����V9p��A7]����gDt�rM'$����Q8j�z��ȓ0���C(�6yI��慽*��r\���eH�]=�fCԵ�,)��(w�1$)D�T�`�yĂ�6v�$��ȓi ���C$;��� �M�2+u�ȓk�J�@�'���I�2���k�Х�ȓo����k*�UK#��+/;�A�ȓ7x�Ԁ��±{��ܺ�@�'e����iH*X�CL�^���CݥE�t��ȓ(�Nز�HӎY옠�VK7WV,$��S�? f|�t�H�d���3���N%�!"O���ak��9<P�
����B�4K"O2��3H��Vv$��?K��y1u"OB1�7�V,2�85pD��>,(��"O��䦉�vpȐ�)�-��A�"O���j�?!f,Bs�.pA�"O�	V)�����9Ȋ�%���G"O�ű����b�@�0!uФD"O�)�P���A�(�[sM KF���"O��gB;E�B��#,ȵm��M��"O�,Suል
tH"�P�J��H��"O�Q'��S&�);7B�J�0���"O����C�eqX�p� ��!;B�j�"O�-��N=Д�ů�.P�jh*$"O0��T��Q�ɩ�1�TY�"O�X����|��Ǝ£��pg"OmA@��T��,��]�����"O�$y7.ט.��9��FVm<Z"O��QA"0#��
F�kV�}3�"OZ�[5����H�G%�`<����"O��pg�69�`Q�E��2���U"O��h ��
�ZP�$�(;��˕"O����ț8#�F��@�}@�#"O�W�B�4��eF	.N�\A��B�<)�,>׆I�v����	t"Ew�<!��#Pfy����.P��8x4H�<�7Ɂf� �걇X?��|{��_�<�������= �F^;�����	q�<��n�,6 ��feǳ13 �yE �S�<�D G�>�T`�J�.=�n����O�<Y�&�
Q���FΪ�,EI�e�<iD�� `�2XfD�2��d�W��`�<	p��
Ί��e���/�����a�<�V폎@����"s	S�"×Q��B��0�Łej�+@6\���b��yR"�T��DuJ�<��Q!� �y � ������x�d�I�IN��yr��Tɚ���Ox���[UJ���x��]1s��܈�$��[�`���A�c�!���K3pb�B�M��$��C�!�C�Z4�A�\e(�E�+!�D9zA.�q�杼c��x���'E�!��.t����	Idv�"�5�!�ǈUHV{�G=��婇��A0!�$L� Hp�Ȃ�!��R孂r�铈�>����%L����hUirz�f�Gk�<�v�Q7!h�pڴ/�֊[W`d�4%� ������H�@5?L��v�9ړ�0<�a�3D�,�G��& �|���T�<�m� [Ȁ��1,�R�.,�,e�<i��� XZ�W�X64��t"l�`��Ԕ'�DŘ`+Z�f4��9g	��i��'�803�CL�̹	&�zv�����OEɕNʰ��D��\�@��"O�5��
"�$�`���4@�����"O<�Ӕ�/A��x�i�Y��GQ��E{��IE3t��U&���<9� ��V1B�D��b?˓SrA@�\�b���#'Θ�x�'�0n��/���ԟ����(@ര7� �f���nm�$(���/�Ԅ��Cˊq�$ı��"��
�6�	%��O��$��i�$
	2���D'	^�P��'��t�C*C�0�x�!�΀W�U��4p{0����]�}!����!!ì���0*��\b�Pd"OtD:@�����������d;LO� �Q��Le~5��/�$t����dZ��(O�O��3Pe��&���j�����'s��6��td�#a�B=T��}C�Qx��Z��s�h��s� �e�|h�L5D�X�B�N*KD�x2o��M��q�����T0 ��1ϊ6p|(Ba��[�����m��O�����BV�1����h�J��"O��! (�X��	Z&&�c���v�i���`�=.ZD�Q �7pp��IU��(#�!�Ő	���B��̈��P˂<P�D{���"<���R+��ؤ��B� )Q�/�_x�d�'���8d�	������Y�W2���4���O>�=�O�\����O�m�2��EŐ���<[N>�)O>��-@���*S�޴�8�H�j0�!�$���R�N��"�2��K��OH��D�!���uI3��8(7�+!�Č0��D#7�Q����,S�s���,�0?��WqI8��MA(sU�� ��{�<�1��o˔�j���V������A쓏~��ӆmǼY�楋�2~�
Ň H_�C�		~X,] �
 �b������Y��h��(��-�"]�`����A�DM�"O-�%��>j�
��'(7T��hq��>��'��zR���m���[�<o��r1`�-��>����M�4\LdjE���~�J��0�O�$�R���Z���Q���$��pFf� D�"�'~
n��Έ�YȀ0�ɔ��)�ȓn^��rs�--Ę%���'#]�'5���m��;b�h��<ҤD>����D:}��L�'�Hԉ2h���顠�*�y/R�@�q3����
((W����y��O��5a�o�N���f/X($��	��y�*�X6��ҭ�(u �@x�.F�yr�I`,�S�j�^�̣�l˸�yW�L��q�����:d�"˚�~B�)�'0"�C��B�%d|xA+
$����R������Z֨�!���l,�T����`Pb��s�Ha��IY�~48I%���'�qO*��z����Đ5v6�2��S�H��"Om���J	Rq1s�G�s9,�I��D5\O���g C;젃��P�H�����'��ɠ[N}j4,��Bp乓E.�c�����xe���(#αXB(Z��&�<a���Oo�س]��y�8��4�@=�y"BC:�P��'��i��it�3"ʢ=E��V�4�#"m��b!�dᕸ?��ȓf� ���NÍ]���B��eQ��ȓ{h��C
*�քRW�� �x��ȓV�Z!��LIj�� ��!���y��CȖ�[�H4��`J (N,avŅ�	X~�jC&��A��b�B$Dؘ0N�8�y��[^~d3��)l}j�����yr�'����dG�|F ��o
dN\�R��2|OH�O(9#g��"�%�T��(j�tU�c�'��|0j��0�CD�N�R�X�l(�I��HO�Oe`�؄$Q��B��SjC�Z���U�)�d??E��T�M�!m�.u(u	��BVP�'�'H�)Z�O�m+��̎T�9V$.)�qH��Ot��*Od��d�?K8Ni1� +���C�JH.N ��d/�Ӻ�ݴ~��[3�|<�0G�%R%
��N]����9`�P��vi�Z�x5�ȓ��|B�68D��S�	�&m�-EyB�|:U�_�T��ԡ�L�5'�P�gy��)�'2�a�P��>�*��تT�f�m�g̓D�F���L�� RlIF�T�V��т��ū6:�k�"Ol�	d猛T�4��ϐ�7�9+��i����#p��(�>m�@�[����̆���<�g�VD~R�߹w94�4*?l,Θ�� ��y��Q%}F ��W��%bm�j���y"H�7`��P�� :.��X��Ȗ(�r�<,O�@t
=Qy�U�C�X�zE�ɹO���6t��F�[M��	P�,6�!�䍗a�p%S��ۦ1�$C�-̼,�!���0���"��D���s0��#�!�Q�f�f(��%�"N��d�=Z!��Y�x����UM�AF�-a���sK!�$�΂	)��9A�h��և�!�L��-[�j'Z/�aS��?/�!�Đ�A��Đ�*��(@�q
N12�!�$.c|.�cӅfH�#�[~!�$	 �>y3�K39{�8S�/И3!�d�&#6���h��;��es4���3!��|h����I�S�����S�N�!��
�/J���N'mX0t`�"�&�!�$��9����SRL���a"E�D�!�$�+# m�$�4j�r��`�~�!�D9��@�앖i�(�H��	`�!�Ƽ]*�1���N��ag�!�G�@�||*G�1.b$�@-g�!�D��K���λ4x��;L�!�$Y!�l�pB��
Es��ݷV�!�D�6g^q��E]�o��� �&ުj�!�7ކ��T$(i�!l;O!�d۹��|ö�9Xa�<P�-��+�!�$ �l~BL "�\�~J&���mј6�!�G�e �p��=z���a/�7rE!�D��G�e�RlE	�n: �[=7!�d�v���V��HX��Mԫ=�!��05M�@��O��d����LW,�!��WD\�"KY�?���2l�< 3!��B��pu�F��@�T�0u�!�$܉m����
�!�2���!�d�-�L.�v8��B,��q8t"O���f��<9)�!AB�z� $"ONYy�!�F9H�v@��B_@9�"O|�+s�R�z��2
��o&v	�"O)q�L�$a�8%*׹#��t�"O^8�h�	Z ��u��a�z|��"O��Y��SG���b��M���"O.Ez�#S�@)jض� ; "O���%e��Ge,9�Iş|�L�"O&!;�Q�]T�2#C�X��I��"O�H�/M�>�<pTA�Uw�t�d"O����F�q�^lz��-|�1"Ob�q�&of�LZs-]iC�9	"O¤���Z'!H�(�I��>?���"O.T�!�W�"�n����4\�ҧ"OF�Hoӂʪ	�4 a[� "O�9AN�0e�������cW�D��"O��I�H5*�ҡ�`
�.�z�r"O4�;�JC4<u ����8�'ٔ0�a�*�6D�ԁŚN"�!�
�') �sa���-I �����B:�ɱ�'��"�懔`Vj�0)�H��x�'�>���U}/(q�Gס8��=�
�'@r�A	�j8���IO<,��e�'̤�9v��#p({��� ��<��'�Y��@�a��mCb��dh����� B9ar��h@y�%%�F��l�3"OvP�V��!^($=j'#ПZ�a�"O��f�dƢL���"Ov��+O<(\9`��w�.p;"O���tc�:P3B��c�I8�:��"OdA�G�/7>:X2�a$U��	S�"O��P�h�?�ny2�E�Z�/�yEO�Dj��"s��)v�*a�!#B��y��O��`e�B�A��T3�y2� ��!*Ȉ/ذ�������!���M�9i%���Z�|A"HA0	!�D0'�.�sABB�3�<�Q��'-�!�DR,E�&�)�&��R��E�!�?p��<H�-7T�� S��;I��ܚ�� �ٸf�o�-׉t�4��i� l��U�%NI Y���q��2D���f $��Um1
����#�%D��� g@�8��h�$��[�ш��7D�`���WF���o�bWZ0�*O4��s�l`bo�-��}z�"OR�q����)�d�A� �[��ر�"OXa�ga�?2`<1P�❖4��`3"O	�pFǽp�d����t��c"Oԙ�3�
�qmC�c��,J'"O�����K��LK�g�r:!`�"O�}Rt�Ӊ" ,�t+� mTȨ�"O����/с
�.`S��<x��q "Oj�*S��77�e@�aW��`�"Oh���ØV;�՚����Q1�"O,dQB�L�J!E��� :"Oح��J�U��%�%�;��ˡ"O��b`�� >)��M_48�"Ot[g�0�����hS� `)y�"O�LR��@�0en�����dNH"�"Ob�H*m���P�!bfrXrS"O�Љ��8.p�a�܅#4��$"OԔ	�m%d�"�:���5bH�]��"O4MaQ�o)�ϊ�\*T����D��y�՜,�	�Aߔx�"����C��y��H�p;���+;�hSD�>�yB&FP���"�_ĲD	#�J��y�T�a�l9�co�E�$���F��y��F/ପ���af���Õ�y�H��B�Ce�F�Z��XS�A�yB�6UӦx!�lD�` �����"�y��܅@%�I�H]u{z�j׮���y����D�Dg�(j2(�G�$�y�
9�l����YJdh	����yr��KZ�� ��&��!�M��yBlZ�?����#��&(ʬI���yRi�"��P���o��jtㄅ�yBh
F�����ޤ�@�!����y��%ǜ`���	|��*�P�yRk��uଐ�ʳ1�$YË���<�0�J�3�,Q�O�(�2jP�Y�^T�w�*Ϟ	��"OD-j��ߞ~�h��C���>;xB���<�i6��h�O|�����pc�X� �!�'����&��	r*�넪V���PH�o *��Pm0�F#�3�$�54�yB��j�0��ٍ"����d.p�"�)@�AsWF^C���z���5+��2d`9�OF �T�k���3�l@;5���'��݂�O���8j4T������(M�:y���9O<@�B%D�h�vH�4f�U�f��K>J��"}��+�b����ȅo֑?)@5K�iI Lr���Y/�5�B�>D�DhRdT|�V)�A*�!N0h�pdB� OH��/O|,� ib?�3�� l]*�Lߙ%X��RSbXE�"�
O*�XV�I�/m�4+'ύ���z7L�%8͈l�r&L�!t���dK9n�`S��E�II�-���x"���`�V��MK�I4;���H�mÙym@��a����C䉌BQ:#/08W��K�`%
4 O�$�Ǆ��H`H�����/�����Y�g(��2ѩ�o!�DL<N\ؤ�P�j��`��T=6L��3�|���=7N��&-v��5���W��8����$F���]��Ҁǁ�S9PP�F�	cl����b	�}L�#%�O�%Z��T�mP�0I5g^�W������'d�U���z�R�:�[��Б$�<go��8#�M/���J��'D���@JN�4<I�3+�,Fgh����9}b��/]����G� �}�?����K%81��Y#y=���F4D�H��o��6>��� �V�6P�%b�d�_�x�y+O�T6�����9���JL�4դ�*�.�
d��-�B�|�	2Cǈ��]7,T�ki4��C��&<l�h�,���>9��>�0�MeH��&�j8��3�D	/�.�q��Z}b�]�E5��#���Y[lT�e"�)�yB��a)lq"�@��_��q����'��	�J���X�K� �D����F�Pya��f����f�N!�?a�MG�X��D�a��f&�@�Be��̋�@��(�py��[3,A'>:V�6d\���oy�}�5.�-[��e*��)Ck�u�ēf�:`��.m�R��)Qx\�Sv�[�N�Ա7jU�<�Waվf�}�t	�q�R��	1�S<4��`�7*H�d>����Ф0����Ȉ	f:����0?I"�.8��t�Z\��<�T�� �l����ޙB�q��M#H��D�,O���Ɇ살�D�sS��#��I=�����I��~�U`c�lT��%�4Y��>Z|a�JG6Uǆ�`2�S?���u�ə(Q ��t���
�Z��e�d. ��R��M�N(���
JQ��~��K	M_�qfBA�-Y4,{�.�1��)�7�?>�����K�r�nh�R�Z����� "Dh@ʚ`�,E�	;{|b�Sp��U��iW�N��g�;:LpU�
�c�(A�'|p����jO��<�	�Q�eD!�� =	FA�xz���"��#\�bpJ��BL��LQ�1-���ek$s8$��I�g�2	�B
c�'��՗L2ve�t�L�-�bH���>��'U�d���*�pܪ��YP̀Re�W�$��
��Xɂn_�s� R�Ln��Ԉ��O/���Z�A$Y��&�/�yԒԛ�D��t\� ǠP���7mH>>G��Q1��6	�z*uJ��{֐ʧ�8�a��c��y�^�⤊�-B�z@�h�.�]A���j؟ȫǌB0���&׿tuI��=y�"�q*�f|�+�G��mf����,�0��H f�=rya�Ff��,t���o���U�^����B%;|O腩�IX+Q�U�B��$z��50��3Q��[;|v�l�'���� X���'X�;GF���O�%Z4d�������Jm�u����·mu�-z������Ԗ�>t�7�N��tO�%���x��
 ���qC�>�"�9���æ2Ov̑p�.?�Y�kT����G�4Ų�J�4#�Ih�X��bйP�ip�=���k��� >�&�q#+D���Ɗ=� �ƪ��h��ى�,]v�؃@l�X����Yd.��>�"<U�h/�)����D�\-Z���b��h`���!3j0*u�i�R��!d�5/�LQbS�ѰAp�,ɢj�J�p��$�0>���[�RN4C��y���%GZN�=��`��J5U��l�/1Q������~gˈ�o$.詁((���âN"�yr&�.[|"�i�h��=�\	���4c���egӟ��P��4+C�m��f�����݈"��dkBM0�<]5�Q��B�ɑ���K�Y�F}֑���B4i�\9���f��9P��]�H:,@o����Fs�'0�m�bbܟW�"�� ��8�iaۓc���:)�n8��e��}e�T��e_�rŬ𺖏D�~�B��D��2��2k�l�{t���H���8� m�%zQrw�SS�]�~�F�� e�����k������J�M�<�C��Yd�0c搯a@�5��叏8,�dȅ�ۃ7n��'[��D�,O�e�ӡ%�A�5j_)Bd�t��"O:M�%ίN8��v%W��:�SY��ܺ4#��n��q�!�_iX�l��EP�R��
��W"o����u�/\OF���Ț $�h���CF��3�[y~@��I��d]�W;$��0rֽB��=�V� � ��$;�ɐB
�""-�m��5���t�
𮀑D &]�RFD�j쭄�G��hG�=��8CCM�0���@TA�s|�siϲ55�
HK����5V����8�4� ���%!�� ^@�P�A3e*ܨ�	� fơc���@(S��C�o�pH�!\:W�^D��	��J	�`oT#s1T-2��>Qk���dF�G��p��jL�)���g"���d��#'LQ�xkr(��$J��0Ζ��>i���]�|��N��m��ѫ`�{�F�bHY�L�|-��9r��u�Ko��j���$��cŝf��X�j��y¬�^||T	ʰR�$�.�@�����gr�;E�I U�։9��-ʧ�y�2G@�I��:ov�c� ���yR�$��	:����)��TC� \0_���x� �޴�"�5u	�-��O��#=���*RB�M��b�
���5�rX�,��+��d؛��&t�2���5qD��-W3^���!���,&��Ʌ��|����b/2��{�'ϴ~jp��$U�1��'Ǐ���d��>�����͚=~�|hRQfE��!�D
}����Ţ	�x��U�&��'�p�ѳ�ԇ"�ܨD�$��9h��jCnѶl�)�#�y�ٴ2��٧�d�&pA��53<�U�0}��ia��`��4��|�\*AѩJr���*`����#�d�" �&$���"��9L�d1
�s.�S�!JB,T�$�L�\Q��I=2Ö��`E%�<eM�9��N ����[��7D�ظ6J�`���Ia�B�}^n9f"5D�� ƥP5hfM;�îD퐬a%�.D�ę��iq��:4��yN�(��3D��	��#�& ��şc*��!'1D�P�@&L���P:�ӵ.�4crI.D��3��ձ:�ip�oQ!7;�r�2D��9Iʽ�b�p���Α�T�:D�$x�j��H���pw�6P�vg9D�\��(ڋ銉�禔	.GB0�]�!��[#k� |��A8w�|��T !��c5b�	�" !4��i0W�6h�!�d��
#�4��eC
U���x��C�I`Xr��Ϛ�`��d��B�U�dC�	
J ��`*�Q�AB䉨}I�A�eE�,�U{�m\�.C�5`�ة3��D3:T�=Kb�W1C�ɷĺ�pČ��K��,��%��c�B�	�*�^D��K	5�䥁'�J�B	HB䉆O:���Ҩ�%���C�F����W�k�p��jMl0jls�(R�'!�Ğ/����r�r�Ƒ��!�� 8�܌�"���v�n�U�ۮ�!�ĝ�Ct���	�:erq«�!�$ޘi�B@�	3�r\�/�)!�$���J���nԉ{zR���� @.!�$��7�N!(�&�(�J��k	�3!���;FA&�Y�"��v�`K��F�b!�DH��� 3�G$C�#�B�m/!�d�k
"MQ#+�=:}�-':!�$ƃZȬ��D��N?6��S���d?!�䆕Jڄh��G&m�0�ċ��?%!��b���'Fj��Q#	WA/!��?=x�Abv���j�V� $��,!�䐀e=���R,R�\c�4�`�Q�h!��%6p�$�IM�f���EF+uH!�$�J���E�y���RЇN(�!�F�G8Bl��M�}�H�C����Py�	�"Ȁ�#'X�G�>�R⮇�y��������W�M
%Rbݷ�y-��p���7e�7c���
��y�Xc�A+g�-SS���%/�yrƃ$�d�`?8W���wh�
�y�&۸��)�w'�7R��1Bn@��y�	�=��9�	9��bfK��y¡$-4��0��)f&��ց���y
� �Y�`��&�M��eP;%���Z�"Oy�Q���O���!��(Z7}�`"Ox\Rcb��+�Jq=(� �h�<YԮK)t�TۤM6�+' Zr�<1#!D�E�q��ȓ%<�E�L�n�<Y��ܑ%ʊ\�V�ܣA� d@�Jp�<I��ľ\�ڑ�E��b0�'Ep�<��n�`l �i� WM��sc�r�<)@X(���/��tQ��KD�<aP�A�W��;��]�f�Ca���<�3]�N�Ig�Ѐ>I+��Ny�<��8H��YqB�W�p���S�<�ч�%�����"
|�XЄWS�<�p.�����D,U�5���L�<�]?lNx�"�ǃ0]� (0���S�<���N$�f�E�M�^�RMf�<9Ҭ�j��Ј@aS�y(D{6��a�<�#hJ]��;��@���Yխ�e�<�4)�� �Leu��rX���[�<yCJL����+�@zT���x�<I�ީ*<��Sg�U��d;�ώz�<�/]>��ؚ@B��|���Eu�<� W� �җo�����*��]�<�n &�"@u�R'F�j�c�h�M�<�Q�-x0�Y��Nq� �k$��f�<`mR�"��i@T��.(��j�o�<�𧇫8bF��JI?A��x�aHd�<f�ӂr�F��� �<p� !.j�<����6�Х�BL.G�F��d�H�<)���Rjr���/�<��$�S	�g�<����]�h�����:�2e��^�<�#K�%v.�(�@��=*�P���A�<!AD\����Ń>{d�	�㊖[�<��@�늘1V�]�����Gj�<���V�KW�]�B�=rt�� `�<Y%a=�Y�Ԧ߄mqb�W�_�<�Rk�;3��Q��OI�p�&�G�<1�+Zl��}C$Ú.�x!C �<�G����*�o[6$�q�A)�z�<Q��+l���0�Y��PQX���{�<Q6�j��@�0*ӵ~T$��h~�<��Ȏi�����7QU�U���T~�<��
v�f��R��/��D�נN�<y��\/8h����}3�Ԑv�G�<)�ʊJФIB�<����{�<a��8<��{S%@�"� 4)!hq�<yE�F�!Z }FʬE4���Im�<y�.ұV�ʝ8�H�6}b��p�<1�S���qB���/�`A���e�<ҁWC��<Y�m�%',U2B�Md�<9�m�*)〥�d7j. :��g�<Qw��}a�����<hQ`%��%E\�<1��U�+�Du"࣒�Q�f�yŪ�X�<�g�����V�͗X��X�B�XZ�<�SI �[~�b�� ��@,�r�<AD���4t�|C�MՊԶX�[�<ї�^�<h)��:K�"̒�Rx�l9��:J�&��'ٌ�#3�a��%��)��!Lf�i	�'�� C�%4{�������{I<�ˆ:<r�+�B1��H�}"˚�A¤ye℧
-^Іȓ���ڂD��$�R����}���K��,I��>W{���w��|�I�F�*MX���$<2��R����Px�ď"t򨹳
�2Q�B����� P8r�g�>�`03��'��Qi��-^�<qʙ�QBq 
Ǔv�v�R0��*a<HP�O� �L����3YU8ġ�r)$��"O� �bH@� P\������I҈hu�>)E����(u"r%l�q��H���;Q0����W�<�����$���b�i6*^���n�Lda�[��P�ʸ;Lq��'���bC�Y4Mଐ[e`Ǆ ��%{
�'�h�	f��AT�	�d�vaqс�d�.XJDA��c�a}nG�/T�����P���aC�2�p<Y�
hX\!B*����X�B�a�f%4�q����r�!�DX�%� �#	S!ڬӅ�� P �'�q��6�G��oΈf�ɑc��.���@�� �yぬm��iN#�T0��S]3��N>9������� f !w��GG�,鲋ں\>2C�I�(�5ۧ�@<k{T@GV�d�)���2�ԣ��'n�JD���$42P�'`ݢ)�t4�
�~`���0e_v���کO�A�c^���iݍ3UV1��"O�@��.�Spr��v�I�]2dpw�>��-P�5-�L�`.F�ȟ̌�Rl��q��" �%-8`�@E"O*y!��$& +�EQ�_)�MR�"�w���'�t�,:&F�>�O0�!�ɯ1.<�+���+C�mru
O�ۡ�Zu �,�r�K��QP E�(�i0��O�/���ē���r��F��xY��ܝ0 �x���O�"#%��pu��-]Қ�q`�&�A�eLϔ2�|B�	2�X0@�a~*|� �/]n�'��L�$�IU���A��(���p���	��Ղ�ӗf��d��\A��'.��K˚�j�w
T�Hgv1B��*`��)Q,.�ᵘ�DK��Q�RL��O��b劶����,!���#$O�P��撍/�0iHƍ6g}���Smi$��b��y�0~�0	��R,�<iP��Pv�'3 ,B�޴p&�ls�.�:M���牴q$�dc�n�z~B��>����C�,�ؐ
f� �^L��c���O9���*�ag
�ۍ�Y���(̻<�F-��	�V���)7��v��'L�=�B%���*�Zj8��"�!?�1��V�ty�!� j$lP(���@�>	B�j7�0�	�ʝuxv@���}kzT
#�r��Qp��G F�N�)���� A�R �Ǧ�'5�=�v�P"�l�j4��4U����*G�h�"�'ܤH�剛�(Ev�5��D�����]���"�ǁ[tyK�i�?&֪`���=-N`4�A�6G����OT����C�7�ً���+��t ߓy�,(�/Ns\љA�Z/@�3�Z�rS�!7N�/��͂P��8%в�J�Eϓq����)Z.��O����X��a� -��y%˜�;v ⟐��;����BE]��3�
9^v�S=Rm��HǆO���?<B6�;��M��zt���<"�����C���O��
�	�:	d2��_� ���ia%�5�~��0fB3KM�)" �o�E
�|�4$"���)��I�4�t�Q��[~�t!sd˸L�=�1AͶ=���-nv؍��I�1R夈��ʚ
M���'�	�~,C��

������lp҅�)�W頨�J�H������<k'JپR�R4X�i�T�f��dE�6���5����Qq�n��S�a�~�hg�ɢ�!Qǹ9b9�Ny����D�����µMC�B��űZ�{��Y���'��)[�$Q�h��"���
a��9Z6�2O�)1���{4L�!���' y-�C
(	9���X��DɢvH��S�Ӹ"aʀ�pZ6�4*'��9j8�B&���U�� #tJ�
�]X����@�
X��0�a���c�B�.x�(��-���zp#�$,H���S O]��Aq�7CJ6���'8�����D�'v:���@�_>H��ɠ��?��{�ϙ	v�ء��=��E.CHT��d���I{��14'ٳ<�V�b$�L���DM�6wZl�FDK�O�̀�s$_#^��O��Sdk��Ng������9��?D���,!�� ��Й/Ox�
ۏwB.C�Ƀ_�h���͜������B�΂\�|$�7*͝�y�A���,�u�ݼ���N*i�D8B�k �"�p�w�X�<��Ț&8W4h^?<1w���w�F���Z&8S8t�U��r�����6ɑ��d��V�"�+#_'S'����[�&�a|��r��$�%�'sd��F�C5:���k��J�q��4R�'Si����T9r$C��Dg:yR��'dQa���I	spν�FJ�X�2��f�)z�!�$_��:�#MP�YI�`��e�_!��"h�Z�F(�s4���p�
�4n!�dNb�B���M�<E$��0�@B!���hhP���;$��q���b�!�MB�����a�Y�8Ru�M��!�� B$�B蝌x���U�Qq&HZ�"O�aӀD8M�<=r'���} !"O����Vg����d\# �r "O|8)� ȑ+�b�xr��=�V8Ӕ"Od���C�@$0���|�qG��
�qO<����Y� 2��
n�b2nS�fDx���#D��Ї��M %���$8B�D�|,�e��@Rx�<�t(H�>ˌ]��-G��\+S�1<O�U�͇9�P0��DBwY��qS�^H�1;[h �"O����E�\@���+8����y�%�*<�����o�Ol8S��!p��}P�(�z|�q@
�'w\�S�I�#;�1j��ŏi����GD����'��9-����	�,xryK��W�7a�,PEjڹ@|�B��.�T�k�#�����BU+p�Yy@�<a1�Ux�'Y�m�CW�y���� nٮO�ϓx��ģ��X,L�{c�T�e�ƴJ@9���%B���ȓG��s3o8M3��s�96u'����<&m[$�SZ��$��-E�-ٖp���)��B�	*Y$Y��c��A�� `Ճk���u����I��0��O���Ń�z#Hx�S@���p�#"O�p�`R�sGJ$��e7d��!�� u,QW�$�On�����^t�ZE��6��@!��'�Ry�g~�$A�2�P� ��H�G�E�mS�yB��-\h��O̚�t�C�$�y���Ag.ԡ�/@�
%̈�����y��ϑ<�tP9PB��5`°
c��yB ��K�HEȖd�0Y2�Ց'K�y��?[�����Ԥ8w�����9�y�LL"We*���j[�>���Ö���y�Ƶ��Pi�a�b����d��9�y2�O:���W�^�Yf���Q�R��y�;7^y��Z�.`ѕ�ռ�y"+���hfiƂnGv\��e��y��,G��T)��^ZV����yRÃR�����U�$�3�0�yb�V�I�ћ���'.l��H�y�/ˤzM��̍o�@��瓰�y��I�#����Л[ify{��U�y�$�0v9
�sC�ג z�UQ��ʊ�y2 _�@�(�2�N�?Ji�4���y�j5Sdˀg�
�����y�K1$\�F��a���'׌�y�f�+�)s�D�\�b1)�`]��y��4+8>Q0/@�#y������y�IY�uP.��'/�5�r��y�BL����w�O�֘ B*���yn�Z�G�.>��4"E�yb#J�UOH�c�2h!�d
�y�K��ctɒ�]Z��I��B�y�M���(YСS�'on��!���y� � `D�2R�F $�T�q��yR�W0����	;~BĪ�yr�-1f���fdBk�5�#-O��y�?��4X��
�e���д�ա�y2B���U��&?b����o���y!	!}f����NN�t�����y�̓0o�H��.�5G;Ĵ�S ��y2%S�X������;�8���̳�yb�_Im(��`��?���Ӆ�]��y@>Wolx#e�ѣX� Qx]^�����(F�A!A�:	�)��"kJu�ȓ6rh�*3f��\ �;��N N��ȓ)��� ��9������Q��J؆�3U��'��`~�Xb1NӍG���S�? ִB�늎����V�*,�a�s"OZ�Qc� �6�t�&R��"O
5��c�&n:9ȧH��4V���"O�bsj������G[DD2g"O� xD���m@4�TEK�7Pې"O(�����#4>p��,��T"O����ۚT���Q���A��dӠ"O�QuhU�+-�8��!�:���j�"O������8<#�H�I�����"O�8ZV�L�Lq�*�֓0H�80"O�d���P�R:���� ;+�;�"O8y�w��&��å�E�)�~���"O$`�)CH�(I
#�,��\��"O����`�1n�(ȱ�G��h@C"O�����_���X98��2�"O*	3�Y. ���a�F�7.a�V"O�|Р��ST�$���"�&"O��c�� ;����$%�4dL����"O4\����`�D�@V�B�B1����"O����*O)i2|b�f�3m?Ji� "O����m�;"�\��A�H
w&F�Sq"OpV�<:) :A�oP^<�U�w�'7�P��ģG(���� �����'�䀰���:8�[q��p/�@p�'���e���ȡcI.j`p�'�$� �..�� �ώi��ac�'h��;T�ֿ\�D��'�Y��8�'��R���5ƝK�$�.ɴ��'���A�X�t �u��35a����'���Z�X�=����0)����'�^)bs�8y�=�"H;
�P��ԫ��6����G�iU��I�<��!�:��SD91ʱ�m�s(L�I�?DV���\[є��!�"���eF�@�p%8B�Ј~_�@`���!^�b�$(#�����Oa�T����Y��EK�*l "F�"f�B�Slܵ:�Z@��'c�,j�'z��_� �w��f��A���*����?3\4�/�~ʏ��\�b��<H���Nf����b��k��˓G:�	��
5O���Ӿ'"��8�)_�^d�I���$E��3���U�4-�"�S�Ot���b*߅z�8		B+F���e�V'ۿ,��Y�7�� ��)�P�MԼz�|���Ԇw�h6�A�j�Fɣ��<�%�p>���螳��s�P5A@�dP��,��=����w?Q��E����)Ѳ'�b�o�'p&�`��0Q)a�^�F��|*G�	W�	+ ՟J#}��f_�A��E��}E%�ç�L�a��Y	X�m�G��@�:x&?�O�G�+�ʌ�`g�"�( Da_�G�z ���,�)�'��t`$�(	9 ŁMGl��D�+$�X*-�U>���-[*�jA�D��V�(����)��Q$V�*�ۏ{���cG�.��QBEk��p93����dI�l�i�{��)_)A^�yQ$i�d�q�FÊ�b�!�$�B�<�H��#�^Q���TP�!�F� 6��!�M�m�"�P�D�!�K�M���BAg�3o�n�K�&�&u+!�͐n$��*�%n���ƀT�7!򄞴(D��P���Ř�IF���#!�/n (P:��P��V ���&#!�H�w�2�a�ߖA���ʓ�='!���:'���bN�X��0�&F!�dV#S�T����(0B�|���#F6!� iW@�!�� y:� �3�$iI!�h�^�)q$��6��EBq`��!�d��i`
!�!&��m�6�xA�,�!�ğyK\)�P�>���h��]�3!�G��&19`h��6�H�	1�N+!�D�(��{@�>���1G�-K!�$�B�T��WC=wn��Aŉ=!���+�<��-�.}jf岳�� �!�muP=B�+d�1�@	$�!�� �D`E�N�x�^�����,{��!�"O�͉0J֜�3��'�� �"Ox� fչr����̤jxH��"O�pAӧ-��ŉ�A�1x S�"O�`PbީR�J�@R�֟i�lb"O�x���F�.3D�2PAB�x��Hh�"ODX�u ��d���`a����"Ov[2NP�G�	��o�)y�%�#"O
�����w�dA��號��|�a"O|u+v��K{b!9C��*[�,M0t"Oℊ1�D�	E|���gltzT2�"O�$x���Azf�!ćA�8 F�[�"O�a0wā�Sz�����V<
�he
�"OJ|�Ѫ�"U��Q�H�����3�"O^�a�L��@��+��/ټA{�"O�t���{8@�����q�"O~]�DᗔC��a:�d��W�P�"O�u!�bA�L�$X(����x8�"Od	�bN�\�f�Kr�Ǿa�jɠ�"O���$�Z?	�d���xভ�&"O�H���� ��1A��E�ja� "O�sr�!+�	��Z�q�p���"O:h1��A�e�����+f��4��"O`�v͗�AJ@�Y��IJ�"O��8g�2$5bb1�[/��PR"O��0�)͎�jV�)+�8��"O,\��҉n�ΡY$;D�9��"O��(�c[�+��5�C"�A
r%*'"O��)wN��Cn4s�aO=U��"O���ǫ$Mez]��a6
�Rh&"O`��Q�C3:�y�Qg�?�D��"Of1�HL,Iߊp���F(]�%�s"O�m3���"5�Fת?9l�#v"O��13N05_,yZ��İ5t<2�"Od% ��Y_��X{��³\/n���"Oڡ��{�(��vc��3B�0w"O�X�+0&���Ҵ�ޚl�>%yu"O�<�T�W޴�8�̀��޹32"O|��Ҫ��E�j�r��.�X��"Of�vNCLU��O3c��dxv"O�0A�ک-�X8����D�<"O��K�:3�A�F�"�	C�"O���HZ�o��X�Q��v��"O���oÜ6�L
!F��c��mg"Ovp#�A*Y��3�Kؑ]��0B"O<,;4��,s��1@H�$d�D�٥"O$s�ϒW�B%�$� �K��L(�"O���qC�M�Z!��'�s���b"O�H�B�ð<=�dcv�ʑ|��Ӣ"O�(p��ô.$���Yd��"O��>,�TX���I6m$�҇�\��y��Ѧ�	���3�2��î�1�yR�Q�^4�#U<{�Y��Q�yR� *&���B�{Qe8��̤�y�n�`�&�c�;���C�y�"O:�a��g������R��\ �"OR�{3o�=+r~��_H��A"On�!K�.BVl� �g���\C�"O8�xL���@�#&^�]�p��"Oڬq�f�>Mp�!�.��=B"O쥱@ W7x`���^(�(�"O(�h��K1�B�2�E�$�p�v"O�D��߻US�|[wR� �4E��"O荓��B�Yv�7�Љ BD�Z"O� `�K�G_�E���w��[-@<H�"Oq��D
�P0 u%ɻe"O8���ĸj�j�xV�B�(��(��"OT|  +�O��%�� ��"�4x:u"O�{ӄ��3Ɋ��C4W�Θـ"O
�rW0M9���E	�q�$5�"O���1��=(���Bŝ:3krm�"O�=�ǒU4Z0
̗wZ@d"O�h�a��*���z���9����"O�8e�	�mVD���ҒM�T��c"O����0i��q�)�7f�l�y�"ON�j���^.4i	 j�%:X��"O��@R��Z� 52�������`"O(:�\�<�f՛'O< �T��"OLA�E/7���c�G�S�|���"OX$�3?\�л���F�d��c"O\�U���Vw
c����jJ1��"OT�k�ʙ�]��u#v�8�Yt"Ol�9�FT�Kx�p.�5~t���"OZ�
W/Ѱ{U@�Y�*S�lad�k1"OH=�5��$�d�F�$BP1Ұ"OPeZD�=b`L�
`�ˮbIʹ��"OrI�6IB�Pgx�jf	���ls�"OȨ'��.9I����:�F,��"O��'�
���j�B�s(f��a"ON���=V�^��Ĥ w&��B�"Oz8`Eӻm'�9z0��[�&d�"O�%�Ɔ��0L�Um���1+�"O�5qf��3m
�ۦ�i�L��"Ot��IS'>�������;U"O���UF0Y�z�R�7'
j��"O6�`�K�0��K�DH�5K�A�"O"q;fǈ�p#0c��l�x�"O֐{VjK3-�P)�c/AT.|�4"O���pOĈ{ߌPS�͓�H�D�#�"O�!�i��v�ظ��AA#j��];�"O��$�:	[�$�t"�3d�A�s"O�H��5o�6h:��ʴ:3j4��"O:e�a�`�*��ԃ�G���'"O$���L/r?jt!�ԕe1�<��"O:AA�q�X�(ٗ"�0p�"O��d
�˼�2&�Nf��e"O)�gJ��k~��U����"Ol��Iϡe����EC k}����"O��c�a�(�|	�E^�lSz�i'"OT��w�/<��@�*M3Y��I=!�$�mE��"��RH�����*��\�!򤚽Ub1��*�b	�&���v!��ۺ�)ʧA�-6!� ��6u�!��H�
:�*����TIUe�iv!�$�{X`�Y�j�2V�,M:P��9u!����Ȝ�5嘐'��,�Ң�xx!�Z�Z���9�oU-���8&���!���F>z� �*�	Ę��iGU�!����d ��ʶ-�rFG�z�!��&Y������u�R��A�8A�!��2mX��1b�1��-aWm���!��@�bk����-z�au�"�!�D��~�P����v�`��5�)ar!�H�Ҽjf��'��9K�I _V!�$��!�����0d�<�[�*��W�!�d�m��| PL�	W���`�L�8�!�dV?ܝz� ͤ*t�����(N!���h�&f�;���	H�!�� ��k�@\�8"*��#L r"����"O��Aiݍ
7Z�9��q�(Q$"O��Ҁ�E/׆���'M1@��L��"OtlK�(��1�v8�5�ޡc�@� �"O�� h�:�֤�s�8��"O�E)���&Mfy�ϳ�(��@"O8�)�۲{I��3G(�0o��4�"O�)w�4�Np��ǎ�d��e��"OPA��Z�W�p�ʣ��1R���!��L�N�L�x����S,6$�Ɖ_�)�!���-.�㢪4����.�!��Ѥ^�:���L��e�#BG���!�d͔'�P���[LY>���6�!�AJ�:���)�E��Q�F �t�!��Nrp2�P�1[~��hU�<t�!�����T)��˕tmܭ��J�\K!��R=$�
�y�
��0Y�q �G�b-!��M.7i��0u�P���"�H�!��`=��h��B�`��@�B�Qk!�D
��t�F'�)��괬�>f!�D����j�-ߝ0GV�ZR��'!���z�H�+��N2.4eS���(e�!�D�!;5؂�2{0��`����!�$�=8;��P�Gk���`�$�!��S#j�t����S_
P������!��E7�Tf2Ti�č��!򤃎f���sj�|F���VK�<\�!��7[�}�W�¿4_¸�E)5k&!��T*��(��GN�f�-&!��G15=��%�!2NP��,*-�!��F�e���B!FÀ�-S�!�dê+Ϫ)`e�ʕB��
��_�!��M4lɢ��5>����&�L[�!򄋨b��}�BǙ2M��d[!$ˡ�!�X2=�r	@p���f|��[��/q�!�$֢0���Qq��/FH�ajU�G<&J!���)�x��"�rG�mK��Z�4!��U>J���z�I�m��9�����GL!򤄸JV&�9@mKi��� ʛ1W!��H�� ��GY�?Q:��eְU!� �a�&�Rh6�Y�D�OD!�I�-�)q�o� W,��(��6A�!�H Q�����
$��(b�Ūuw!�3nθC!d�,0�d��!B!�U���X�g�v(n��M� '!򄛂��DȎ�|z�2�L]�l!��B9b�����TD��T��1^!���Q���B\2%:b�г�ϼ`�!�D�2�٩� ź6��p���y+!��އt���W�:2��xdFE�!�Ę�9Rfy��/	�g02V��c���ȓ\'��� @�?�     G  �    �*  �6  aB  N  �Y  de  �p  �|  �  ��  Ӟ  �  {�  ��  R�  ��  ��  (�  l�  ��  M�  ��  H�  ��  @�  � = � � 4 �$ {+ <2 �9 �C 2L vS ~\ �d /k rq �w �{  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+��6#\��	�<4�d5h��'�B�'���'	�'/�'�B�'�♈� �X$ܑ�ƏMm���B�'��'�2�'Gr�'2��'���' M�`b���ЌO� �l���'R�'�R�'f��'>��'���'|Ёb)�/ܘ�s�R�j�h��'��'V�����'���'���'����a�)c�4I9$F�&ؑH��'9��'��'���'�B�'B�'7H���j�
^����@@3uw�h˰�'�B�'"�'��'�b�'}�'�LgJ�����eC�SG�6�?���?����?���?i���?��?�w�ܙ/=�I�p�,��P1s�3�?��?	���?I���?��?a�Ӧ�8��"U;E�q�"��:hZ�-������H�I؟@�����ş��Iǟ�	pX-٥M`ݪu%Zjy ��7S� ����	�8�I㟄�������B��R$@�.A#���������M�I����I����Ꟙ��ܟ���쟀:Rj�\W� ��C��z�%��aџ<�I矤�	ӟ���X�	���ӟk��=X�m�N�P">1{�(ߟ$��ٟ8�I���	㟔���Mc���?Y���;|���C��)wLzq�i�>R��I�4��������#&�����SP�^�nH�Ő���3b�.��?���S�<(޴C�̥�6)P37
�遢i�E��:R�i��e�%#I�F����B��Xᤙ~�T�%���d��9gɕ��
c����Gy��L��P׊/���0p��*��\Aݴ�Z�<	�����y�.�X�z����"g�u��ꌇ4. 6� Ϧa�����N<H`b7-u���v#�Ji���#"U��j�x1�D�(5P�� !'u���T�'�vh��+n&�a(��9����'y��a��M�2�UH�����ဴe�|H�u6���Y�\�ش�v=O2�5nH��w�P�'��487CՓ,�V��'e
%�EB##D��a��T�!B��ڟ�у��2V�b'-�*H%Hdҷɀ^yrX�`�)��<!&(��I�VɊE�<B�:��A�B�<)�i�H���Ob��4�i>��F��,]3�h�b-d<�������ݴ`̛�'��s7�i���"�"X�a�PoEx���̉S�\�Ո��"�4�@��k�iy�Or�'���'��fY C��|U(��|"���b��g:剬�MЏL�?����?!L~Γ�"�A����8]Җ�@�G���R*O�Yn���M�x�O����O*교����@,����E�v���ꎷ_k!��'��EZ�o�KҠ;V�$�X
(Of�� ��bV��1Eͮ�������O���Oz��O��<Q��i��e(v�'��yeL��6{��ӖA�)N�Xj2�'�����<ɒ�i���Za�D��]A���%� �kg���@/�M#�'�&<`�L�U6��I�
O'���O��NG�ߝ���6ND09��O*I��c�l������I����	���b���x��`DH�����'���?����?I�i�&�ȟO�2�'*�'�L���2ZѨ� 2��6x:�2W�$�d�Ѧ1���|�2!/�M#�'\h�2W�D�V�|��Ti�K�o0`�g&C�P��>�To�<���?���?ɇ�\�Z~��A�#�/b49�c���?����D���± �����IΟ��O��"��P;V�5�̈́+����OFʓC��&�p�R&��)d艻p��7Y��!i��T�@��aB��<�l�������Jٺ�Ŏ�5�u���<�;i�@,P�#.�:����-r������?���?�S�'��\ꦙ��e�k~f��@挨<�LA#q��.��8����p�	v����D�ͦaY��ѻ�,�XG*�
*c���B6�Mk�i�*A���iO��< ��*�+R)6��' xM��]���u�ƙ1Rmzm�g�w�|��?	��?���?1����iLY��ǧg����G�U�~A��
oӨ�'�OT�D�O&�?Q�iޡS�J��9`�x�VHؐ-)X�B���M�D�i�O1���4nq�0�	��L��!E�/��Iq��X�d5�扌Zph���m���'4d6�<	���?�tJ[<�tDڡ�Ț.������?���?�����D@��ғ�Ey�'�>-�� E<���{2$�h<R����<y�i�6-�Z�I��"f�LB� qXw.O
p���Ӻ�H�.(�)�<�S��
�8Ea�A�^��3�JE��xó�@������?1��?���h�~�$��?�Bj� q,M�G�(w��$Y���� D�$�	�4�?�;�l��(�W6�s�G�X��}͓J��v�aӾ�m� ��l��<q��9x�!���	�����J1E���2$J�D�V������Ц1�'�B�'�"�'|�'�IQ`"��8���;�I�E�$kBU��k��$����ԟ���p�ԟHs�k�:����#I꘹[Dn�iyBo�\n;���|������`�0rp�)�;h ���H�n��8fG�2��ѳ�,�b$x�).O9o�dy�C�(5{�]H�Ke㘄)F�ɢ�����O��$�O
�4�`�Q��F�1J=ܝ��1I��8@�|�qg�JSB�'��O��`}�v�zӢ�o�'A���0��7bΈ�������#ūæ��'D|<sӁ�/,�5zaY�t�Yw�� ��H� U7ux�<т
�i_�<i57OR��O&�D�O ���O&�?A��FE7���oC�#s�|B�`	���	,���4��Sߟ���S�d@P�� �t�@���ʠ���"I<�2�i>t6-��t�	�erӚ�����:�F}Q.tA�jޟ:n����>Q�l����W��ٔ'�>6�<����?i���?�e*8�b�(''L�
TP�V ��?1���]ͦ�1��ɟP�IƟh�O@B�ɩ(���@6j[|܈�O�˓a�F�o�l<%��S�?)P�"�3,(`���m�+X/�9�����m�ፊ55����ɖp���P �ϔ�X��m���  	E3 �J�c�5zʌ(�����?���?���?�|"-On�nڻV�B�14�^#RtR�H	+�l,br�0�	㟐��R����dAҦ5 �AF7c�t�&�ǗV�0 �kŰ�MW�i�Xisc�iX��O�+��Q4lD������<��Âv���XGh��Ib�i�y���^�H�	��t����I���O��Ih�K�~e�b�����ëz�
�j%��O����i��O�2��y��T3�0������T�h@7mEǦ�9O<�|�Մ(�M��'��AN�9Ě�+��q��q�'˖!�䘺��Xw^�S�4����On���%:?f���eU�X�t� m�->����O�d�On�iV��\4R�'�2��TFLZ��l��9I���:�O��j'���v�81'� ���2gk6�3�h�,v�(�b&?�f� @�yH0��<��$��C�$���u7��Oj���D�$�̥�"&N�k��Z�n�O��O����O6�}��=�R��7�#�Buyc�� ]��`Ûf�L0)m�'��4�|j���	W��PR�o�"�:O��oڲ�MS�i��iI�i���"��i�o�Lל�9$� H�֝ ��nf|W�_y�"tӤʓ�?���?)���?Q�����9S`��``��#���)O"Amp�2��͟��Ik��(:���3bL;%[B�xT/7r!��!)O�ym��M3'�x���G�bp$x�
�7xq�e�Y+a�0�±���g��I�fM��� H׺{�Z��c޴���#H�X��,t˾�uEB>01T�d�O��OF�4��ʓ_ɛv- r��B����圷
���;U#�= ��'X�OJ˓
țV�p��lڙU���8�kƹ j>壤Bޤ/����L����'��tx�.T�U(B��Q^�p�Zwc���3d9d���̝I��x���y��'1�'���'`����E��T@��\��4�Ác�6��d�O��D���X� z>��	䟴$���׫�-3>u��k9���v���'��
۴I��O�x�&�i��ɐx]�]3
�'at�A ���_��]�#��v��P@�C_y�!oӶʓ�?���?�YmF0��Ba ��{W�W�>�P��?�/O�po�FC���'�W>�ڂʈ6Rxp�y����E(��jP�6?�(Od(lZ�M�v�xʟ��95-k���&k�&��+�lL�#����L�Cr"�&h��vy�֝��4�L�t፿k�X �L1aB�����O��$�OV���O1�d�#����6,0�C�n������Y*�	!�'~��'B�O��g���n#������V:�䭂���7�C��q��b�٦i͓�?A�/:nLL,���&�� �  R '8Ϯq��C�U.�<���?��?a��?(�>P�2k�� � E�� "`6�9�ɦ-Y�A����	ߟt$?����ݾyLN8y���d�H����@�MJ���4G'��f9��]5:]�6�|�0���
2H$@�����@Y���a�b���D@���q:4��^�Ipy��'7�F+r�0�ʅLJ� ��5�EUO�2�'���'�	%�M�!����?����?�B��vzR�E$��AH%H���'��I��M{t�i6�'�``��iԈi���s��.(�ݘ�'�bNI5��;/Q�9���?eq�������'2��+�쏾�80�+�&�����'�b�'���'r�>���>M6hB���&q�|L�0A�b���	*�M30 S��?I��?i��w��)ʦ�*��B&I�+FO�)��'��6mЦM�I�K$!nZ�<��[�p�J#]��e3��< Vx�yËK0J�j Z��W������O�������'���'����Go?l�D�b�-[;��!��_��ܴa���)���?������<9�\)�^-q#$�ʮq㬍1���EѦ�i�43̉��O] �����.��D�vǕ�)��:2Ǝ�\���T_���׫
<2���;N��'��	�^�n!����
��H�*6r��	������i>U�'�$6��4�V���>T�����:�!bP�^�S���$�Ot�0�' 7�F���4u0:�[d�B�\b��aL�qV$-��١�MK�O�Y�i����z�f7�	�� ��q�Y�\�Z�R�m��C��$J�0O����O��$�O^���O�?QXF�Cqo�ab�e���2��şl���H�ߴ\D��'�?����tV��3�ֲ�,+�d�)�D�G�xR�hӴ|nz>��g�ʦ-�'ˬh���8<׶�tl[�O|Z\HU@�O0 Ѻ�D�|�_���؟t�I���Z�'R�ci���p	��o�ѐe^����IOy�Ee�r�8���O|���O�ʧ����I���Q��L%r?0��'r�		�M�f�i3�O���S$ PcB:<h�D���5,��j�%�n���vy�O������|�_6dѤ��woD0�j�d�" ���'�2�'f���U�<C�4�G�V)lxԽX�
��适����?����?Q�X�@X�43dL��l9k�m�qB��ZԈ��s�ib �!��=OL�d�)�� �7fG�[��S�? ��3�L�'k���ɕ!+�A��?O^ʓ�?I��?����?�����i�L+���ӛ;���jN�W�Hhm�xϺm�������E����iޥ 6 D5h�M��A͌}�@c@�Z�M�D��i[t��7�b�`#��H:@�Sv� 3b*���fu����cb��s�RX�IQy�'��O:<�e �. $�1Q�⊚M���'��'剗�M�e�J��?9��?�h�ZQ�m*�/�lH�T�!���?�M>*O�HmZ	��'�
%�F%Α
,|8ˏ1y,$�q�' ��{S:D��g���?Q����źs��'MX��p��O&��e�[P�XӒ�'���'{B�'g�>-���/�D�{�'@(~t�آ�U�_]���I��MK�O��?9���?!��wC�Xe�Y�3S�ȹR��#Jfx�'��7MHӦ���0I��m��<��%��"'��"n��ʕ�< �M!��H{3����H����$�Ox���On���Oj�dM�8��q�w%W�y��+�-Yu��Gm��ޢY������&?	�	e8Xm{�Ü�u�($BT�5ur��'�D6��a�S�'_�(�����d���i��)�D�k�D"GJ*+O���fOѻU�֝ �����XP��R]��Z�x��H�"P
�$�O����O��4��˓,�v/ͪ.BBg�@-e��W%]5A�GX�u2�'��OLʓ.���ø>���	S��9�U-X��ȷIX�F��]`ٴ����&])�Y�p�B�Bmޓ���nm���Yb��Tu!$��'��O"���O����O�� ��)���[�uV(}�ti��i H��͟��I8�M{F�P�|���?AO>��%��j�r)�C�w���p��B̓����>��d��M��O�pIdhY4�ؑ���F��abu�8����
�#�L�O�ʓ�?��?��1P� ����|f� �4�,�!���?�(ON�o7(T�'�b�OE�ĉA�L������H�a9�,ɵ_����<٣�i\b��S�?E�	�Y���l�u�;a�C�l����Ī]<\�Vɔ'&��N��J��n�^�ɄUh@�!B� S��#Cc��)����h���,�)��oyB�b��a��� ���;�C��:�ڴLIDn���O��$#��My��k���&��$6�"ic��H�P|�ಓ���}��4Q�<�;�4��ė$2�:Pss���Ӹo��<�3�Ѵ8%�!���!h��	cy��'�r�'�r�'2[>阇ɟ8EFi�v�1S���B]��M;ǉ��?1���?�I~:��?ͻ2�,�#S@HU���-�t�T+��i��6U�)��)~�nZ�<	&�U�f_ �;�(D:@�8-Q���<a��D�D2�oؒ����4��dؕp�x@�$3�e��� �?���d�O����Or�� �u���'�b�>|�m`t'�2Θy���EC�O��^��vlӌ9'�H.̆<[�:<\�5@�`F��h�dx�D�1�сL~��ß�uGg�O�Q�Fe�<�`arC?iҬ(A �O:�$�O����O��}���8��<�"��:� KTiS-jt��6b�I�7g�2�'R�4�0�!T[>\u�*�K�<��r0O0�o��Ma�i[��j��iu�I suL���&�'?�j٠bJ��9Ȅlrpf�-|�~1(�	YM�	myB�'�B�'�2�'uBK�\C� 9壈�X���� J�/s��I��M�$�Ԅ�?Y��?�I~�1p���E`�R�<=�bdVhF�P�(O�%nZ��M�F�x���l��i�F��R.��r��J$<;f���ć;s�	�+�Լ
1(����|�Z��Ú
@���%U68�����j��L������I��AyRh�R�:���OΜ��G&^��)siC�J�zxY��Ox�d*�Iry��h��t�'���gH� }�Y��ȕ\���� o���3O���_"���1+����:��U�� ҅G�\A4��G㒵W�(ϓ�?���?)���?�����Щ��0���VL�S�����'���'�d7��o��)�O�D>�$�{w��0��<j�4ics	��1O�eo6��$߫��6�!?qq��)�L�82�]�W��a�@�:M\������ 5re�J>�.O��$�OL�$�O�E Ba:[*p	��J��W��H#$�O4���<���i� ����'��'��ӄY���g�īa�0}�5/]�_�z���$�M��}�OR��+_W���,�3sx<(��ѤJ>Pse�`��h2S�T��-�r�;y�'4N�PsE�~�^i(2b+j��h���'w�'Z2���O}�ɀ�M�Hʠi���y��ĉ+�$�x�fĠa�0�.OR��,�	Wy2�pӲ�t�WoY%����*,H��ۦi3�4q��)�۴�y��'�̌�AJ"E2��wQ���3.��t�� �[�{��A�6�l�@�'4��'4��'���'��HT��Հ��~:��j�&��c��4A������?������<Y�Ӽ+։�'z�����N�x��H����b��`%���?-�ӯ3$XmZ�<�s���B�yX2"�	f�k���<1u�o1�8�� �>������O���]Yl~�e�S 	�Ѝ��n���$�Oh���O��ӛh
���'����t���@��3�=9, j�rP�D�۴`�OV��v�4"����fgT�,�K5O��d�Sf�96i�<����*��ۺ�uI�O��j�l@2u3�#�q4<�Q-�ON��O����O�}�����ku�]�q���H!" ذI��H�v��(-"�'A��4�x��B˯��T��a�Z`�1��<O4�n�"����~�(6�=?�#�2���I�K�? ���C�=�2�S�`�� i�TS%F1�ī<Y��?����?���?y�Hb�@�%�M�K3rp�Ɩ��Ȧ-�!�������&?���x�z���`���p(�.��|�'��7��@��|����?aB�KX`Qʑ�t\9���N87+B]������Е��f{�Q�I>a�O^: �ƖB��i�`~�Ω*�'^B�'>�����T�$�ܴ�����9�8 �rLH�i(V��5�ё��?Ɉ�U�2ܴ06�f�'��X�g��-�v�;������HC'�b؛�9O�$�ayH�a�R0[`˓�b�;qs%@D	-8%�Ի%�	2(� ��?I��?����?�����Ox�D��gW�*h�i�6�Uqh1§�'}B�'|7�v���O:��"�$��(1�
����?� �J{�z�O�l�5�Ms��hZ2ݘ�4�yB�'��
gZ^��8��,~Ν��iد'��� ��
5��'������	����Ƀ���b@���iC�y�V�?�6P�I��X�'[�6�Y�xN����O$��|���Ku ����z@��V/D~bS�h�ߴ:��&�"�?�(#�K���u�Z�v��5��$�2z�T���X�(��|�mR)�uG3�{����E U<M']˂�8H/^���O<���O ��<y�i&���mA*%�8`#��S�1�]zp�ΌS���'���'��'�剱�M�f�[P-0���a�z0��Pn��o`��T�FNr��I؟x J�
��[&�)?��i�`��,@�oJ<4�S�<�.O��d�OP�$�O����O��'|����P�[���0�59�@�{v�i�^=�B�'��'��Or�y�(�j<���t�MC�V�OP�p"�i��6�[�)�S)G��5oZ�<�e��P�h�ǪCQ��b����<D��6�~�t������4��䅾j;̠CҫB�9]��1������Oj���O&�4؛V,Db�'��T%�����*h���DBb��Oxʓ2כ��p���'��u
]�F\��s�	�N����#Fr����/:�t��J�8<=���������u'E�O>ͺĎK�S��H�W�Lڝ���O*�d�O��D�O��}���{"�M���l,;$P!��� @�V�b�2�'�"�4���)1�	5(V��A��S~(*C�>O`oZ��M���i���g�i�����t��@�:�l�EU���Yk���(MA�STdv��iy��'�R�'��'�R�[�'cl���l��
�^E�JۊYd剾�M����?9��?AN~2�$�Dђ*%/%@�#ߕ0̚=�)O<�l/�ا�O�hɫ�Oք�Hp���}�R n�h�\���w*� 
H�����'��ɦI�~�۵��|P���W�D�B�"Q���4��؟��i>��'U�7���>�Df 4�r���#8,�Sǈ�U�"���O �D�'V�7̀{}"�0 �\�RM���$�c�'�a�i���O��#��lx�)ĥ�<�����s���x�`-A�X��'e[�<���?���?���?y���lH	)r ÀG7Y.���%*���r�'¡�O ���O��'�'�p�'+��=�|�C�H��(q(���y�{�bY�'�V�01�ih�	�/��]��!Tz9����ԩ���������ǆ@{�IUy��'��'�I(BȪ"��,"�h�R'�+G���'"剐�M���Ɋ�?��?�+�F`��C1c�zu)��Y:����� �'<p7mw�S�Daڞ[��0e�ۂs�2i� �8U��#G��y9�[��@�칮���'����Ӂ��<H4=���B�M
TTZ��'HB�'�����O��I0�MK�AչVir	C��J P��b���`B�s���e��Z���$�ƦM����/�DD:��8ؼ���ȴ�M��i�H�!��i��I&/�ftH�P9A�'~��v!W%�2��#i��F�����D�O^�d�O��$�O��D�|�t	Gx��ģ�a�s8 ����R��FN��B�':���T�'D�w��Uf�ib>��T�C�"L�B�h�J�o����Ş)#P��4�y���Q�M��־{�:�k��y2
��De{�mC�f/�'��˟��
=%�ͺ��U��0���w1��I����ܟL�'�6�U*tq����O|�d��P�r�����oZ8&%1�2�0�'y�6͓⦕H<1��Z�E���+s�ܖ$K�]�q�]~b�F�$8���&�-Z��O��� ���h�	��T�����+qb~|)��F�In@��ɟL������Il�O�R�RW�����b�5b0D��)>�Flӊ�s���O���O���]q�-ɇ*J����S�%?*���"�MK�S� S�dAͦ�'8�� B�oX�����=���̋$?L�a�ɘ!��'<�	�\�	�����՟|��);K��D�Z%*�n�H�FX�X�'��6�J�1ʓ�?�L~��h�dD�'�na8�Xd�ɲQh)-O:�mڲ�M+ �x�O����O�0CEM�'(��+��T(ܨ�eFƂ9�(��O�Q�+���������6\:QC��=�x�K��c����O���O��4��˓�3|��⍡d��rV+�/Bh V�ŋ�y��'��O��A7�V�e�@�m�1�=�bn�/�`̉�H1T̮UCS�M�'�P3F��Xɠ��}��;}X�yB�4�Nd���@%f\��?����?����?�����O�0Ѱƍ1>B�Y �U0�ޱ�QQ�8����M���\M�t�'U�'q$ .ܨ�Xw�οx��K���3
y&OF<l��MϧR.� �ߴ���D�� ��@�>=֚��FoB$(�8�q!+�;���+a�)���<ͧ�?9��?)s(�%E@Q��*	�b�ޅ�#�N)�?Q����$�ĦY1��ß������Op��I�W8�X4�ʒi[T�S�O�ʓM(��)�)-�=Wɦ%Cg�4"�zH��Oт��!��!G`�M`(O�?��݄��r���&�7���e�2/5p����?����?�Ş��d�Ц%�B���ɻ�̛wo�P�,(L�:T�I����I埄&�4�'a47M-Z9q�#�>�3�eC ^`,�nZ�h�.�ߦu��?���
2u�$�@oR���d�RN�x�"ی�"i��aR%bN�<����?���?��?Q.�����AK��P{@H!d<N��1��¦���A�ڟ4��꟤%?����]0�*�aw�D�o&*Mht�1YB\�۴\�;���D�apH7�}��jb�YsW��@�26Y��a��0���.C#�9Sc Aq�Iny�O�
B�]�4�x1�� �Z`���S�1�R�'��'��8�M��g���O"�"5���w�4ʐo2"��	�$3��`yR�s� nڠ�ē>��}�R��n�.�/�>4�'����?U:�i����7i<�	ߟT��+Zu�uSd�+h��{� �ǟ��������0D�4�'
 J��Ϙ!Y��`�-��O��Ja�'&�6-[9�����O���%�i޽����`E�] �S� _A�B�u�H*޴kD��`�*A"�myӈ� �@����T]��Ѽ[�  �uB�"6H\!:TJ������4�����O^�$�O���	#�veQ���*m������˓9 ��NS� C�'���'+�t�f��sb������q�q��U���ڴ4d���:��	�K�u�
�#j�Ș���/9^�J���G`��.Ȧ��Ej�u&)�ķ<��n@2f�ʴ�L�M`��a��Ð�?���?���?�'��ԦY�'�	ş�s�lL3I|*�s1%��&s�1;ǀg����}���D�Ҧ1�4|���jވ4�$����^kpy-u�jm۳���M��O޹ʕ�G� vQ��k4�)��a���H�^�t�+p��k_��cE3O����O���O��D�OJ�?=��!���v�`���*��� ��Dӟ�����+۴sEr�̧�?�����TNyE� �
uX��Ѥ	C�4�hM>���iF�7=��@��Bn���D�Y�G� �~�1D�4'�H�RF�p��A��������O����O2�Yخٳ���}�DS�$����O.�������k��'Q>���#�>E���@��9�D�a;?�.O"�m?�M�O>�O����>Kd&U����	����� �᳤��3{L�i>ŋ'�ú���|�Ǵ=��#��-sv��ꜵf��'��'���T��i�4.+~e�%K)H ��q�E}�i��"���?���?	��䓢�˦u��h�3��5`�:@[.-��@ݤ�M�A�i
��iW��O@�1䎓!O�
p)�<��Ƈ=�P�`�N�طN��<�+Ov���O����O���O�˧9�&eЀ�N��E0�m�0r=x� �i���'���'w��y��y��ۓmr&}���^+1�X��%��=��7M�禙�O<�|�r��1�M��'\�5��ʇ��J���	��Dn>j�'�|�����3�<`JԖ|�P���Iٟ��FԼp.�	A��V��<��Vן(��֟��	ty�/z�~%���O����Op��c�9��ed�zd)!�I@yr�n�d-m;�ēRXd���?4�X1�2o�B���'KV����Ď��jw����F�$����J��_'f0�l+�I!̈́`g�������t��џ�F�T�'=�I��j� [G�|�bJܐl`<��e�'�F7mё8\D�$�O���3�i޽(�o
<�� .�w��!#U�v����4:���'DNIQ5�is���O.�3�M��w�Rp5�A)�D b�\>l�#��+ ���Ofʓ�?Q��?A��?�O�@q�v+\&(uDCr��*�*�`*O���%���d�O��D+�����R���=F��J�7�N�
ry"�d�<��>�'���~���N�KO��s����Is�JE���J��.O�ItɅ>3k|�]/�䓕�dF)K-�eBФ�|O�����A���O.���O<�4��� ��&�A�E7�Oʰ^J�q��&��zpB�ͅ�8�B�'f�O��]��֡�>q5䍻o�z��F�Q�$�R���Z2C��Ŋ�4����W�X4�c)�44n>��X���vZ%���Ug�>ɂ�F$1���O��D�O���O��d2�~������M ��!���1-6��ȟ���!�M f%��$�O�O�([����6���e�ܛ=\��I'Kr�ɩ�MS��i<��	��f=O@�$��c�Z�J�5��mr��iAL�T�¬t�Ȕ�k?���<����?���?�H�'8(���Fq������A�?�����D���	CD�͟�I��ܗOCzј�LHݳ��[��t��Oz�g�6hw�R$��'B���RU��E"���F1��;%�(xi�G�U���4�Re�$Fݵ�K>��K��*�9�E�9ij�c�*�?I���?A��?�|�*O�=n�5}��r�S�V�  �h\�+�L!P3�ڟ���ߟ �?Y(O��m��I�"�r1 ��[~t����	$�8	��4Q,��/B�_�V��b�`˝R\�����IybiZ0X����t��L��)p��\<�y�X���Iן��I����I�ؔOX�]�MɆ"j��1@�
�ܩ���ӌ(����O���O����D�O��L�����D����4���1<�Mm���ا�O	�	�Q�i��� ��A&D�����>�x�E3O��#n۝cB̠Bq�.�$�<����?ٳ=L'�rH�f�UA̐�?��?�����Ŧ�2ć�����ڟ|���t
@�,���xW�w���_���4 >�'؞�H�#��b��<I��6O$zA{�'��Ȑ�e����	�?-�t��պ{��'>��p�N��=�\e���1dUP�'���'cB�'�>��	�o�j�@v-]2q�,�j#@3W�A�� �M�3����$�O�杻3�Ty�@b�+58d�u-�:�扗�Ms��iQ|7MO)G&47M-?����3<N,@�*o��M�Z�6eNY�4 T->&���N>�,O�	�O����O����O�ݠ���5����!��&
�|XѲ�<��i<6)���'���'���y���&@�\�ׁ�|���.�Hl�I7�M�ִi�O���J��O��z@:�gX� hO1L��B͉�^���,�(5��c+�u�K8�ĳ<�,�x�`��-�488�#Я�?i��?����?ͧ���H��u���̟,��K<���zqn^9��Y`t�p����o���ަY3ܴ!�vȒ�;��B��Q�F T�)VK�'>al퓳�i���%M��X ���x�P�'?��*N����'XV����֗K0���۟���͟��Iɟ�Ib��I(d�4D�7�ű'�N)Fa������?���e��+����'M�|BbK���ЦQ��:��];�ġ��"+�����Q��|���)�M;�OliƄ55��`����@/�Y��ܵ
F�C���dNȓO�˓�?Q���?�9��ݚ��ȗ�������V��P��?�(O6�o��t�d�'�BZ>���]�@V�X�r��4{6&Ũ�j"?)O��l(�M��x�O6�$m��:h�����X�qb��p��}�F�!l��5"�	��O���I1*H��5���2,����Q����4Ô�xFe1��?����?1�S�'���@�Yͫ�N�#$G	>^x��BFL�%�Ұ�	����k��� Ҧ���Ŕ3pIѰ�n�t��H��.ȫ�M3�����ܴ���\� �p�r6Fл��ӭT����Η�<��m�0l�t��	ny��'��'��'FbR>}���X�P��B�1s����g��M�j#�?!��?�N~*���?�;u =A�F�(Wؒ���� �RU�ic�6-�U�)��<,�|�mZ�<��-L8py�7'�I>0���<�B �#9}�a�� ����4�`���%�YU�=*����#ў� ���O����O��d�힐���'���#q~��ԍT�a �\��� hJ�O�ʓX����u��%�Pr$�D�d7�ÃO�?:>��Q*?1���A �a��$��'d9PXw�*�$�ΪU9+T!�1K� [����$�O����O���4ڧ�?�!�Ct�J��1:��"���?�E�iuy�'V��'��O�nȢv��y��;	�h� ��+h���ڦa��4+��&NL�^?�=O���	���'�H�[�p���D�_�	c�*<"��8u`/�D�<����?���?���?a��8$�h���o��4hO�(���N���ӟx�	џ%?�iIBKH�
J��rgZf��@���<)ӷi�6MO�)��3��I&��h�7Čv��)R�ܧ8ä�)��#@L��u'�+�Ġ<��Ɗ%N�����IL�C�[�� �?���?q��?�'��$S˦	��H��/���^|)���	=���`� ��U�����LŦ[�4\��N�'tZ��!Rc��&��vΝ�~�G�i��	=8{�A�3:��$?��]&>��IP�G� D�4�('�	џ��������,��Y��	K2�9Ī��DX̫R�7?�%���?)�4�����<���'�"�|��sj�'/�d����P�>O��l��Mϧajܴ��D�'#B8	�h��*���K�Q���P����A�j S �,���<�'�?����?QR.� o�ԑ�E�`Z��r"L��?q����$Ħ�#'�����O��D�|���^7d�J��-�x*�LLX~�W�[޴<�V�&�?���o��qĄ�kw��=P4]�'*��y�4��#L��u�
��|�!��uW�>��@Rn؝y�*Û*��-��A/
L��D�O���OD��I�<�ѵi�����&_�F��=�fʿ.#j���}l�IƟ��?a+O@�oZ�R��@$��0"�!�5ݴ���U�q�����0H�";D� Қ~:J�`^$`࣒�T�=���<�)OP���On���O��d�O�˧u�,��靇�X"s�`����P�iX8Ŋ��'f��'/�OgR��y'JT<z��pA��WIȞ�2�n�� �V7��Ѧ��M<�|cf��M�'�#`���Q�N@�g��{�0H�'�i�e��E pٻ��|RR�l��̟t�� �Ȕ�y��ϰ ��!��������՟��	JyBia�~<���<���I$����د:x>U���A2Ia.���r^���ݴ|��5�4Q�B� �GLu�Q1���z��	����ida�6��b>�Dc�ݺ;R�'�~��B¿P_T��"OT*%��)��'b�'���'��>�ݴN,@��oW?k�t rnŭ
I$|��
�M�eC[�?���?9����#V>fO�px�N�~�4x ���<aдi��7��O����e�r���`���:(<���.ߓH��1�Nӊgq$���!]�!��1%�̔'Mb�'b�'���'��yp�/�>w��!Bt��<=�0GY��R޴A$����?�����< �5:Q���ѭ�~��P�&�3������޴ul���O�z\�� n�pԤ�z�D�(��4cX8��j�~ʓU#���D�2�u׈'�$�<)É��$w�Xdo4�����Bڰ�?I���?���?�'��dI��a���ٟ����l��ag)/p�\��Env����\��������ݴX�F	�R<�����CU�)�mO� �p�襻i���=�&��⥛a��y$?����D�CY�.4H=xÉ� ����d�	ϟX�	�����_�'\m���򤔾()�A�Z������?�����E����	ɟ$��В ��<��	JE�I�r(8���	�ē,��e���4�
6�1?a���$�"D�>uۊ���>�\x�?A���KO>	,O��D�O��$�O2�J�-U�Y��L�wdI�(H0k�Ob�ĥ<��i�Dݘ&[� ��z��cM�8O�e��Y�*���;��+��$�<��i��6�H}�)z�딁3��������+J�v�VQ�D�͜ 	(O�)��&&4���WBi�"��(L���0���]�X!y��?y���?��S�'����٦5@�/�U��� w�����BEZ5��=�'F�d�<�2�i��1
�oQ X��#SiD�g�L�I�N{��%nZ5 �Dpl�C~r-Q#Q��L�0�ħg��ɀg���7Q��K�
����^y��'�r�'S��'�"Y>��gg�$���R��߯�2�[��5�M���Ԟ�?����?9�����yW�"�l�`���w�1��;n�7-W�u'�b>�"4EN��q̓�!�S�Z4I�
uz��܇r;8-ϓ,�l� �S�T�x}0O>�(O����O��B@��Wq��{&-8l��J'+�O����O��<�c�i�����'2R�'W�`Rv�����,�P��0��&��'d�ɽ�Mc·i$Or��CP�*\7	*�X1㛟�դA<������/�&;�2��;?�.C��ċa�� ��yyPH�f�B�'�B�'�R���P�Ůx�f ����AH��PE
�4$4%�.O���1�i��1�ER3&N�8+k�Sn�S(u�4z�4GF��t��D�)~Ӥ�P��T���T�= H:uk�9k怡d�^c?�mF�%����4����O���O��L�;�����R�8���p�V�M�dʓP��Ƭ�y�B�']��'
�3�@X��D��=2�W�4)ٴ��F 3��I��?9T�ЕfK�5�d�b�M������P D�r���<C~	���ɺK��|\�� �]F��]��,�'�d���ܟ��Iܟp�	���SSy��o��a �k�O�t@`fF$~�\@D��"�`
$�O���*��OyR�w��n�Mk!�e�̝XP�M�hp�[���
x��m ڴ��D��&;B�#�Y�ܸO/G�>(��!tF�fR�PǮц�y"�'B��'���'7��	�p�śR���@36�;��d��j�O���OLTo�@��� �	K�ɉ}�m���:m�&,�#l�5k���O<Y �i�7=��ڧ�lӦ��}b��̀7�^�i1�#/����I͝\j��IӮ������O����O(��
a�%b�J��*S��0�K�&�P���O�˓7ś�,7���'��U>�k��#�� KE`H[�|K��+?�-O>,nZ��M�K>�O��Ј��R�*�8�U�+b�"h�`�pj�d\�i>q``��Ӻ;�|��Ѻs� 8��F�9:V�SCi
����'ub�'���R����43�*�JE��
k�\Q�k�^�j�S�����?����?�b^��Aڴp��L0�$[2�1�L�;
���
U�i�ҩ�1*͛撟�r��hhqEy�ǁ)`e�cEV��ر�/��yBV���	�,��͟�	��,�Or"UOԁ�U��8d2���쓈�M�6�!�?)���?�H~"��?ͻ?�����3�܁0bf
+v&��A�i�T7M,��I�5S�07�~�ȣA��(8y�)�`΃
+L)�ćc���I��t$��Tb�qy��'�r'ʽ`)�eӭ�,z+�P��D�G��'���'+��M�ABھ�?i���?�s���"3F/������o���'%剝�M3t�i<�'����%c��ݶ�{��϶%����O�m9�ML�au�$�3�Iݝl��]��?�6�ݛ	#:+`˃�ƀ�V�ޭ�?���?����?a��	�O@��#/kF�����9 &� �G�O�nڱo���������B�Ӽ���<_���KwGh�b�M�W����?����n���d	�^!R6m&?�b�Q���l�u�������'�!�j �Q�i�4�H>�)O*���O �d�O"��O
Q�c�Ƒ'`��W͈�E{\U:D�<��i�^T���'���'i��y�'R W�Zayg.��P8�z0�P+	�	�M�װi�
O1�$j��J#j@�*5͗��9z���[Ύ-r�<��hD�R
*�
^w��ON��hU13`�L�� ���&��x2���?���?a��|�*O^�m�_,"e��4��Qᄤ]�;^,��N?^w,�ʟ`�?�*OD�nZ/�M�ưi28�H��Y��P�W�M(�
�`�a��QO�����*d��("}S6D�v���ߵHq�ûᘵn�a����wN��<q��?-�M���?���O��}�+��ªeC�M����8V�'���'��6�m��)�On��4����l��Y&��7r&f�pA�bu��<���iW�p �@�4��d��P��0��C�Y��=�Ѡ�(J��PR0)� x2\1ǩ6���<����?���?���?cV�(Fl�;�� cQgR�?Q���dCѦ���)����	ߟ��O}�� SJůCˆ��A�\K���O|˓E��֋?�)� "�J`� ��$BW`J�3�u#��A�8vv����^�6��|��D\&�uWL*��G;;�ԅ�7�T�$�p����m����O����O���i�<Iнi ���g�Ɣ6xu;�aԂ	�@)@ C�z��'`"���<���i��xC�d�88�TL�Öy��z��>a3�M.�MS�O�L��
�d�n��� �<Q�+�2q���׮��v�2ݫ��R�<1/O��$�O`�D�O���O�'JǤY�٣4��i0�$N���u�i� ���'�'��O	���yw)�	2���U0.�T��pʃ�XWF7-��}&�b>���*NϦ��rX��J��d1���+:�` �h.jŀ%�i���K>�-O��$�O�!)�Ok���!�C��99s �O��$�O��Ļ<�Ҷi��8���'�2�'Km1�ʓ_b"<#�#ʕ!�J��4���<q�i�$b�(�c�7mθ;�&>�j���#?�w B"ahR��c�7��!ff �[w��DF$6\@��
G�`�jGnS6� �$�OJ�D�OR�-ڧ�?�&�O�z�X(� \2bq�M��?q��i��[����p�Ӽ��c�G(���8>����<y�i�6-�ϦQ;�����q�'X~��Q�O]qp���c[`��i��O'1�`�Qp���D=�'��i>���ܟ��	ן<�	!n{���+}�u1���zC.h�'�6�XRp���O���4�9On��t넅>�4�A��@��
O�<�r�i(6�l�)��1Y���[g>Q��c�L[�xũ!��v�@�j5>��-�u*?���<�bC�#>��R���!�|�A\!�?A���?���?ͧ��$ʦa��ן@�fC�E74�X��,� 6�y���J����D�֦�4L��&Ͷtp��3���=`�2��󁁲_v^���iF���\�;�/��m�q����3�Z���k\m��1㠇�
���O��D�O
�$�O*�D>�S!�F\����sm:�̎c�j��՟T����M[p� N���'��'�l�� )Y_�,k�-M�)�l�R�y�am�T��'z�	�iM�I&c�u�@P.�v�bn+F�H��I��^�mвl�O��Gy��'�B�'%§ˢl��ôk�N�r� �m�''剏�M+�����?��?Y(�*�2�c�J�}[��"a@8������'��6��n�S��L�+�L���ꋡ �dQe��6 дY��P:7�L�\��>G�, ��@��'����Qw���!@�]~*�u���'Cr�'O��O[�	�Ms�D6	�tDB�h^�Vpس!`CLXU����?i����'8�1�MS!B!���#w#�>ErP�4$�(����j=nE~!!rfr��bj��	�w�M�h8L����.Kf�Ey"�'cr�'W2�'#S>���HWM��{�o���tG�%�M��j���?����?)M~����?�; t���0h�j� ��˻\�dr�i4Xc�b>ek�b�Ʀe�X��%�A
��M^�la7�N4"XD���I� ��u@DkH>�(O�$�O��"N��q?H���E1mi�	��(�O���O.���<af�iX��0�'���'�
� DD�'0J��\�5�����$�<�i�Nb�D���Hjp'�iä��2�$?��N�9����Ř���O�y�\w� ��\�m�L�� V�1�H:�.ݰ�D�O��O�$>�'�?��ݛw�T��ұ����#MS4�?���i���Q�'vb�'��O�nE�Iu4pQt�����4�Z'��D�צAۯO��d�q�j�7��M�2I��/��Q3@�%�p�Q�>Wd�
������D�O����O(���O:�ĝ�d|�K�����D�!AA��˓9�2���?���?yJ~���I��ls���.V`=SGF���D0/O:Um���ا�O���RE䉣�H�:��RL��j�l��_�t ���j�Z���z��'G��k:
,� ��Q�f�](��3#Aϟ�����d��ݟ�my�nrӆ��F`�OȠ����w�B���m�}�U��OL��!��ty@u� m�'4����<rȾ�HpfE��B�����+�F��
��-<�J�Jv�`�S��p��G�"Z�H�D��?�\h�FF� �	۟X�	ɟ@����j`e�U`TkA�cHp��옵�?A��?q0�i\��؞O���'�'���R�H W����闝�)ɏy�mwӠ��'M>$V�i��I�g�t�Is�I�A�s��c���t�[�3�j\(t		c�	}y��'`�'�r�F��,�澌h���9T@����?�/O>��I�e$\�$�O�ĵ|���I*��q�K[<5Ɏ}�uk@~b_���ݴi�O�[� `�� �6�0��惜��ν��@{��R��]y�O��y�0���$�x�$�]��a�C�X/N$��G�ǟ,�	֟�����b>��'iL7�לQ���A�_�oa,�r�ʇ�[�J�i��O���Ol�t�'��6m�Yw�%L��,Z8���]�;Ѷ��'
FicQ�ii�I%yڤ!@0D�&t�R���e/����� �eNt4r�hQJ�<�/O����O�d�On��Ot�'D�2cˊ/T�1$�G�g(6�չin���'�B�'��O����y7�����|sdҗ�n��S,�{��7�E_�S�'u�"ix�4�y"F6P;X񻣪�?1Ƽ�3�C��yB��3-&�Ӏ���>J�'(��ҟd���R���7�Na�S�a5S|�$�I�����'��7M�0z	���O���+n�4ؠ����F�k:��'G6M�S�? 4=A	C8L�D�����
�N:e���c�YC�.)
$όt�S3D��1�;3�� 

7���10��ji�X�v�֎)-r�'w��'���ß��qh�"�,)�d��,M�D�˟��۴)"0�*O��$$�i�Zp#�X�D�)q���X�Os��[ش(���|�΅
��eӲ�'�ة��a��C�d�Tk��$Hn�#�ǆ�V?���q�M������O��D�O���O`�$@0tr�`�I��<���úV8�ʓ~�V� �2r�'�2���'an-ZJ�99 j�	���&�
i�@Q� ��4)�V�0��)n� �bT��R����G@�R-ehj,k%^˓R����Q��uW�5�D�<�P��)nf�y7gL�<ъ|����(�?���?����?�'��M���h��ǟH��+�y����/]>����h�	G����ğΦ�ٴM6�f�ѡ}.x��F�#�T1���W=V�ͻ�i�ɲ^�l\�Tj
]��&?��M��5��n�&vGĕ+ஐ�4R�	����蟤��ԟ��Iw�'}�@s�$ń?||�t������?��TכvᐯR6��&�H�Bg(0Z1�dAXW!�咆�ēZ��v�m��i?C��6M ?�QO�v�Xx�c�Ϝ�"�rBU�^0R��ȁ	<�H�AH>�+O�d�O����Ob�J �\�~|faæ��)al�0��O���<	��il\]�D�'�b�'4�S
�d�(�e�0J�Y���ɸ]m����d����4����I�%ݼ��� �i>B���� FRB�1�,ДuHl�J�o�<�'	A���]w�@�O��٣��ED�)��Y�(bM�@��O��D�OB�d�O1��˓~_�&��*4��s��5z�e�18N�Q�b�'�B�'��O��Gԛ�IN���hAo�_nb	iAE�.>\�6�ߦ�8�������'����Q&chnahaU� �&� j�j �`��7,����Eh� �'���'JR�'��'v�S*
u�8���P�&u��c$NbAxx"�4��$����?�����O	�w�����T�uo�}Qb/D�i���#1�{��nڙ��S�'Y�0t��4�y��L�R���I�h�N9낢=�y"X�p �A�(�.+�'�ʟ��I~ټ S�h�	l�z\ �nW=x*��I�����͟��'��7�Q�Z2j��O��D�p��)Q�N"=�1��I-f4��'��6M�঵sJ<aTiZ�,J,�{�덠oA�)+��J~���H�ha�/ϟu��OXL�Xd���5�ɚn�%0�F������Sc����ӟ@����,�	K�OhR�;X������6QR�q
dΎ��nӮ�#�*�<�����yW�C�L
M�CD�JV���R,�y��qӈ�l���M�U`W��M�O�$�e���aV�5�ε�"Ǳld�U��aE�=��=@K>�,O����O<���Ox���O�l!a
 cÚ�U��kx0�z�B�<ѣ�i�� ���'��'D�O � �"�WfZ^�TEB�-Ӓx�I��M�#�i�6O1��]��b�9%.H0�� 2H@ڂB�|a����<q銎$m�epZw�,�O�ʓC,f�)C��P�H�����?Y��?���|�)OV�l�8p���!zq.�[�DV=Bа���/ �	��?�/O�xm�?�Msd�i팜 ��[i�8ڡ�J�kΔ�Sfdۢ��f���S�*�XP���Z����e��ڈuF�Pr���M�]�$`w���Iݟ��I��D�	ݟ��*v�H�6�x���A6�JS�D���Od�mZ�
x|��˟��	N�	=R��p@�P6.��}kf�T�eTX�3M<���iј7=���B��m�r�k�d!�4e6��h0��T;�Z�ƥ?A"�Qs��������O��D�O��ǅ&p|�k���j<@�z���1���$�O�ʓ�V�?���'+�Q>a��ߚY��BK	��)�p�;?�/OPl&�M�xʟl��iX�R)h��fj�k肐��Ҫ8���F��Cf��|JGJ_�ugF0���g�2��؄���H$�ݺK#���O ���OL��ɠ<�@�i'H9��)˲6h1ie�����q�4Z�r�'���<9 �i��L�����m�W �"��rCo��Yn�7��nv~�����x4� 剄!;�Xpi�p�9�7� �1���	Ky��'���'{2�'�Y>�B�̓Tj��1V�?P���� �ˬ�M���Ɛ�?����?9L~����?ͻYz�x�ҍԳ��(Cg�
�B�^U��i��7-�n�)��?f"l�lZ�<�d�tk2����.w���i���<Y���g�XC�j�������O��DkpPQ�c�~�\��L�}����O�d�Oh�e$����(]�R�'���6T.,A7�Q�]OFr�L��4��Op�w��6�pӎ�&�� R�H�oz�D�@��E�H(2?�!��	�n]��f[���'@�*��]wQX�D�7$"��B6)�n��HiFgr����O��$�Ol��0�'�?1t@^,԰�2b�͜CA@� m���?�A�i:N��CX����O�Ӽ��H�e�����6�Fl΀�<��iw�6����if/]Ѧ�'G�H O	q��B��&с����8�wDZ)E�'��ş��I�`�	ğ��L��j���2����EW�(�' 6��6g�@�$�O~��'�9O�%�Lm5�e��Q�&�h�sǅ�<�P�iH:7��}�)擾w���ԻN��}[�,��$�Ȏx����'[�B�-�=��{�	vyB��t�� �R�MO��@bI�)���'L��'��O��I�M{!�C��?Y���2��U������ƒf�r����?�.O�Ao�"�M2�� ��
&È^_F�'&��,-��"V�&Z�7�3?�f��l��)B�ܗ�䧥�ۅdP�w�����Y��$� � �<q��?A���?	��?q����C��Y�%f	8���^�3�2�'i+~ӊ�[�6�d���Or�O��A�җg��bC\R8�H���I�	��M�&���4fJ� F���*Q�Z���4�Jx0\��)G<q->d��ò- �8%�p�'O��'���'(V�iX0��0�����g�Op��'��I��Mc�� �?����?�*��ѢC�%E���&�NG� ��Ő���'Pv7��P�S��c_Ғ����+l�s#,�0$���/FI�ꍊ`���4� T�t�]�'C2�"uk�(?��T"�q���@�Erz$��O�{��6�X ja�%Ev��pY��e�V��c@<*���I�OyV�1���4S��(W�Q�8�,�iu��h#�	���`AZ���/X��H�1e*+�*ϕx���$�����Hy�ܴ0%p!֭j�<@�£R!,��K �Uq=:m
&M�$ e���پ2^�E��$ݻ^����A�_;,T@]�ä��I��d�pg@;N� Yr�#�28pr�8�+M�[^Cd�� Y!z]#C��e��+���8~���S��+��ᆇ,�<tK�ֶa����`��N��Y�}"�'X�'��ɮEP� Ka�W��j"$�
X�&u���"�	ß�����'N��Tks>��Q��6s��cC&��M�PeP �>���?�N>�+Oʩ"�V���HܤOx�(E�m.n�c4��>���?����d�* NҨ$>1���L��dc�j��!����M����䓂�D��)�O��P����- �IS�"�n�
��i�R�'h�?>D�J|��R�[
1��z��=o
�=���Jf�'��ɤid"<�O�P �镥z�R�E�d�!�ڴ��-j�Z�l��i�O(��L~2�Fj��A����Nq� PA*�M+O����)��"$l�doӨ3���EH�.q�n6��">�T`nZ؟�	�������'9l�`D�$/����*@��h1�w���B�)§�?��CN7y���Bf�ͿL���B'��f�'���'�L�qbH2��ߟ��ɩ@���֣� �i2�D�94&X�}b@�'�2�'Kc�^>��a�g�����ց�<#0�6��O����B�^��ϟ��Z�i���(�*?�WO�;ᄐP	���D�E1OX���O0���<��#U�F��x
��Ѧ?�0�s��ϓ&��)��x��'�R�|�R��P��T�M�ꀹ���N�H0a_j�c���	՟��IXy�Ez���Ӑ�%��`OLe�V�1��O���"���<aC@D})��$u�c�9oE>%[@�^�����O��$�O�ʓ@J��{Н�$-E�^�Ve��"�"} ��)�Β L>�6��O�O~���U�d���r�C�Q�@���Z�q���'2Z�p �MB��'�?��t�FPi��0l�<���1���e�xb�'��*�N:s����BX�k�H��۴��DE�(��Qo���	����������5��f	/0ndـF�=f�h��i2�'�N�b��d:K���ٓ�!��x��fj��6�T�t��m��	����S�����<���7��BOפ)� -])=ě^M���!��ҟ��g� u5(�P��";<�Љ >�M{���?���)-�-�Y�Ȕ'�2�O����f��"��l�@��&�D	��O����O���_ \(�y��)J̈́8	�-��U8p�mZ����N������<�������Qh��+���Ъ�r�� ��#E^}�LD,i��'�b�'�rW�|JыǞI������\�ˑk�"�f̂�O���?�L>!���?c��p�����^	����S�4,!O>9��?�����d�s���'EU0y�@&Q� �~M���!\��<oZgy��'��'���'=@ف%�O�u��X? ��)��S�_2��5\�6�iW�'��	*��{��f�������ܤF��)[�뇑9��nZ��'�8�	������}�t��ѐ�?F�pd����B�nZ���INy�-S�=-�꧞?1���*���M��qCT�t&B1p��ӃcF�'���'w�	�����?-��ʇ1]8��gX�j.�Pr�eӰ�m��A(E�i>��'\b�Om.��[��{��|���Q3�:��pMBƦ��ݟ��B�G�ǸO#�a	R@��\Rd�1l[ O՚���4:~�4P��i-R�',��O�r���$M�c,� ��Q�1�4-���W"HYZ�m\��"<�����'�L�0�1�D���(�+p�ZImӶ���O�D�!gD���'���ğ��:�:\��V�_H���JP)��$m�8teH�=�Z�����'g��'.4 6T43����˔f�@ő1DsӤ��Ќl�&|�'F�	���$���*DiJ`�G�E�4h�q(wkܮX��+�f!yK>���?���򤎆�� W��b�� �[�Az����@�I}�T���Il�����ɞ��	Zt�S�q�تc�$E�Z��Ya����I���'���H�u>ɀ�����(�	�x\Z��J�>1��?�J>9-O�	�Oz9��J�"Wt��Qֺ/B��;EXe}b�'��'��ɔZ4`AO|Z�(�<$�5���O�УvI�����'�I��D���$�'��'V�\��jN�J�(���+G�oZ۟��Iey"	08�(�(���kl�u�l��&�_,/b\���F5E#�'Y��?Nή��}�Sb� ̨��씆Q&>���A�-N�\�PSZ���	 z�pM��џ���P��tyZw��b�@W�"(D�AB��nX����4�?�u�v|�%�TK�S�c�d���8_g�d�6�ʸ#(�mڤ8L^��	՟4�	ğ��HyʟdC�G2��RW�� BW���ܦ�����,�c�"~"S��J����CgW�a���	�� �+g���'c�'5���`U��'��	8�<�yǩ��&���*'��2}(�yR�Ň"��b?��Is?Y`��>n��4@�@���eǎ���	�r�|�'`���'��9�!��� �h^�dx�ˤ �>A$��:��'`��'C�W����!3_��G@̿ {
�$��)s��M<!��?9I>),Ot��N�
r���
�l��َ��GZ
U���$�<1��?Y���dB/gut��'m���h��S��;_Y:F��'*"�'��'+�ɵ2�<��2s$e ��|��Q�iɶ6	ЬO����O��d�<�PG<~b�O�`;�؃9���{ ��3��uZ�l���$7��<y����?�M?�yc#Т&����oR�Z���9�On�����<���7�(��)�����Ov���0����w��9�EG�Q_x��b�x"�'�� �t�.�(�y���Ӕ�[�~-"��-/0dS!]�t�	$I֬��ş ��Ɵ��ZyZwt�5!�C�G"\Ͱ��������4�?���;�$��E� H�S�'_k�r�+
;^��(ԧ��(�!o��h}�ش�?a��?a��;������^߮�p�9W[ ��Ġكv��6�q���O����<��DW�(H�I�f�:-r5`��	��akc�i���'�r��k��O���O�	�*�m�7�@&��%�4����6��O$ʓ~W^�ЦP?�������z-]*b�z5����|�j��� �M[���L���x�OY2�|��*i�
��� �|�ܹ@C#+>��M�<b����D�OB���OXʓw	�a)ߜO&耵���9VD]�l��'7r�'��'6�I�����h�8���P�9s�����?�)O��$�O��Ħ<����;g7�MK2�p*��^z��	[:��韈�IT�iy"�W���KF';�j�`�N��X:��= X��?���?	)Ot�p���W��Z<b�X�n�8�q��5�h�ش�?qH>�*O�	0��O
�OSZE���+�EJ/�3OJ1"ش�?����$[��r�'>y�I�?�X,w��A6�_h�.	��%��JiO��k��=Z���'�����&N.n����7{��Ӓ���M�,OF�@ME֦�������?IӪO��QP��āY2㢔`��?����'��L��yҗ|���\.�еx�N¾&�\(��������� ��7��On�$�O��I�{}�[�p��O�M� ��6ԕ�WeP��M��H�<aH>i���'84�1V�1��i�*�!K<p˥eh�X���O@��ͱ[�D�'��ß���# �( ΋H�6Y��-J�B$Aͦ�	WyB�  �yʟD�D�O��� U��!$��N���XbCJ?	��oZޟ4g����Į<a������Ok�CZ�ы��v��T��mO������+�'2�	�?u�I�̔'*���re��0���z�AU��I�7BS�-��꓈�D�Ox��?Q���?��9Y'<�#�K�)hIV%��([�Nm��?���<v�����?i/O�j����|�u�����)&*r9b��ݦ��'��Z���I�����%̠��(_�H<:��Zu�� �.8|��OV�$�O �ģ<���C�e���ş8:!m+�Tv�Еry����Q��Mk���$�OH���O��1�9O��'������ݛb����@G3q/��ٴ�?A���$ϸBp�m�O���']�d[�;/�L� ΟEV�q�\�$���?!���?��b�H~RT�4����榑>�\�So� "J,(ݴ���_)O���l˟L��̟h�.����T��CJ8b�9�Q�ZH���iUR�'��
�'3x��<��� Z|xh��DDK�q3��j��!�MCb®8��6�'�b�'��h�>�-O��ǆ�*"��ˇ΄�D�̕(��e�t�u���	yyr�)�O ��u�/줁C�N��_�R}��i��������l�I#�$��O���?��'12��"����P�8��K�Su]��4����P�S�$�'t��'�PB��5�(�c�bЇx�%���|Ӕ�dU3Kc��'���'Zc����d�מV��yR�kM&����Of4��>O4��?Q��?�,O���	܏{�����!`:�
�ض�0��'��I�,�'���'�"�X#ʘ�!�5^��tI%�N�8���'��'�'8�Q��ae������m�n5����K9'
�	�cn���M(O
�$�<���?!�PD�� ܰ�0�hٹe�4-vQ@�����
�M#��?����?Q)OAa#�S�$�'eMq�b��1����.4�@:ĨcӜ���<����?y�Z�q���I
0Y¡[YB�59&��S6m�O�d�<QĀȈr�ҟL���?u(`�
uS���E!@3*�hY�������O���O���4O��Ĺ<i�O��]��X�@�L � ��Z$Ș��4���90�>�nZ�x�	��D�ӹ������a�M
_[N��l�+]��%��iM��'+<d[�'cp��<��D.D'>�HEHa�ʩP,@�1�n���MWjݪj*���'j��'���"�>+OJ�q �YLD,�tN��zV��"�GΦ���c�<�	@y����O��� H����]"#)��`�&�h��i��'M"ɷcF���$�O��Ʉ4�l$�l�$[`0U�+o�j��򄎨��i>��I֟�	"��P�!ʟ�fQ��$Z2��Cܴ�?���/3��~y"�'?������)<�"a�%�	r"^�r�fO�T���Q]
!ϓ�?q���?y���?A+O�!q
,|��i�Rl�Y�)ɀ�0��'��	ʟ,�'�r�')�Z����Xr$6�"�AET�(�'A"�'�R�'�T�`0������˂9��0��W�\��5��4���O�˓�?��?�6/Vg���2T�0`��!��D}
��UeY2��D�O����O��z��s�X?��2T�X���D�蛓G0`a�P�4�?Y-O���O����s �O��ە&��X��ɹ��V�!��p��i���'�ɔ��MQ��<�D�O��iU�kh��v-C� t`�{�E\&XL!�'�'��d��yQ>q0��Ti�G��2V�˅H��:=Z���ŅݦY�'�^x��oe�h���OT�d��ԧu�C��D�ꆄJ ( ���O��M[���?�gS�<�����D$��_�02��9[��ٰ���$~6m״si��n���Iɟ|�S ���<��^�. ���q��c�T�C�֛41�� ��O��?A�����D�R��!�
^5��3ٴ�?����?�WoN�%��Ey�'�D@�P����L��
�����|�
Q��yʟ����O<��í>^�i3�*`���!��A��n�ß��㍪�ē�?Q�������K	�V�hr��x,T՛Te}�"˱�y�Z�l��̟��Ijy��.=DE
���[����D�3u+]�c/4��ҟ�'����ҟ�k@�*5����%d$p��C4%�l��IAy��'���'�	�]RJ�H�O�:��Ǫ�Qޘ��f�:24K�OV�$�OB�OT��O��[��O��Kc�7?���  ��N��I�#K}��'��'��I�u$hK|����,�zu��=3W�% '�W.u���'��'��'>,ebt�'��o��=�$Ū@��a表��Hu ym������wyj�,d�������=r3&ϋ^�vy��$�q ���H�I韌��G���In��e�C��+�Ѣ��(��d �"���Ք'<��P�Jcӊ�O���OS2����8�D��T������L�7;��oӟ��;Ӽ#<ю�t�S�;�2�`X	RG���Db :�M��%����'���''���7���;����L�%%�̓a-�O�\4��4f�������O�R&� (�QK��6+�>� �@���7m�O����O��y��u����d�	U?ytKY)�a�§ˆ_� ��l@�!'�\S�-~��?����?YVJ�R<�����ȉ����/9���'�"�@1� ��O��D�<���s�����i��ҺZY.<��Q}�썝�"Q�`�������Dy��H)w
բ�����3���*`Hw�0�Iٟ�'� �	ٟD#��M�7�RI�D�׸?�ta`��Вm���	Dy��'p"�'�	Y��b�O�`��tm F$�<z��[:�E�O����O�O����O�E.U�N���wɃ%%�����J��r��?9���?�-O6��W�Ja�S�?]��F"F�E�|�t���rR8��ش�?�N>���?aଌ�?�N��Ѣ���@_��k	�
�i���f�d�Ob�x�6T�����'����]΀1HU!�N�7d@
�q��?��O��dH�*1��$"�Ŀ?��@��/~�u�a��=t(F*|��ʓ?���&�i��맿?����f���a�� 9'LxC�� z���?9)��?9K>�~���j�xvg�%��"�ꦕ�@g�$�M���?q����S�x�O��Yh8i�h@�@�\)1�ǜ{j7MۊLɈ�D$��ȟ�Cc-5�y"+���8��t��	�Ms���?��9z��(O���'/A<8r4_"e����hæ\���	���ʯ2�&>U�IڟH���p,���[�Wb�@vJ��k�4nϟHrS��Wy�~��S��'9�xQ��]�VC�:B��
�,ђ�`�>Q�X�%����'���'_��	���Xbv�
�~�x�\9: ���'"��'Eʟ�D�<�MT�{ђ���ڸ���'�5K �C��F@~��'T�Q�����i#b�'�\j�j�p8�` ֵ *m�ԟ0����&�4�'�T\�����M�A��fjN�i�1Ĵɩ��ZK}��'��\�P��jG��'�~���,b�8(#GV�Z�X�S��M���䓉��^2B�,(0�x�L�W����P�@�To�p�����M�����O�՟?]�'����հr��]c(8\�x|:�
;L�O�˓8�6ي2�T�S��ǣ >�Њ����e5<� ��^,����OR����O����Ol������Ӻ+�g�^4�y��#S+|4V��ť��ɖ'2,-PB��ј��O��8p�L&���)p"7����4O���i��?���?�����?�9 ^�8���Ce�VE������M�b�/J�V��<E�T�'��bFĝ�3�.I�s��$mv�a�rio�<�D�O �DGY\N�S�������5y]�ep�T��5��d������<��Ht�O�b�'�2�Kk9t�yu`)�ȐI�@ţ=��7M�OFԀV@�<�_?	��d�	<`,c5b�.�^H���b���O��i����03�	��P���X�'��� ���wAѨ-��9fE�{F`V-W��'�2�'��J�g���� R�I�Fݹ@v[&�d�O��$�O"�d�O\e�7!�O�ᵬM� ��ZT��z`�H�e�榥�'U�|R�'T�3<\���4S V0Â̫	��� ��F!��'$2�'n_��#r��'��'B(	B��,M$�"���3��1�i �|��'!��!��'�$H�aF��R��,x���(�Ƚ��4�?����d-T��$>����?	ʱ��Z}��`�#[P~}�1n��ē�?����j}Fx���,@�.QP?����I<H��R�ii剕:^P[ڴu�S�������>��c�����	%�ӡLh���'M�G�O
�>ك$��<7ft
�R�H�i�jӜ�;f̦��	������?-�I<i��a �ZwbU 
|��u�L��-�E�i5���哎v�$y	uL��k��x��눴 �й���xb�|U��A:.d�HʡG��p?�!GBz��%���?v�8���<)CJC�S���E�r��s�Ư>LQ[����#N����6=kB���F��r0���@<Z��aR�ŏiѾ4�g4#�&��/-i��q�nL�f�(�S#�G2F嚁q��}�"
L"M��Ģ��_�H�\ٰ�G�,�(A&�M蟬��ğ���	4�����ޟ�ͧ��<90O�7YLnWA4&a<:v��5M 1S�\1�*���#Y0yQ�#ߘ�(OR1��.�*}�uj���*�t(
1^3G��=�w	X4<�.��A��")�*�R���j�'�PŻ���?�2�H�7iP}#Sm�4�����ɲ�hOĢ?ɀL$b�T�����, ���A�Km�<�惼3}:�����~U)Y�
��<�$�irB^�$��H�&����O�ʧ>N�!���i��H�GԅY�/��?��?��P!�N�B��&QlҌqEA�tk�bɔ(O�|1&�I�J����^�m�1Ey�d�{~v�IE�(}��i���Vx4�P�GG�&���,4�la��*��� iDy�l��?q���OSl(�T',d�t�+�k��*��p��'s�2Y6�����؈O.����DI��0>�F�x"IƘV-�����+F�h8�Z��y� ��Ӟ7��O����|��(X��?A��?R偢r��=T`�q�R���O�)��c�n�;vc��d�,\�+#̺H�d����;/ڴ��6,ҕE@��fg�x �ʋ��|�z�fن#Iv�`u�@�P���m�*'"q�(��y��$S��Z�w�Vݷ}$rUf���l~J~2L>!"�vw�� ���4!������k�<��׼8��iפw5c�B�N�'S�#=ͧ�?��F�|=p��P�Y$0E�TO�?��,},pQc���?!���?A�{����O���T\a��A�bAb�v�3�
�7�ꡑF��C<4p)��J&�Z��;���H��MU�1O��6)� (�j9PW%�
Y���AwO�T����cZ9�MU�@��	�L�\���y����, �����+����~RA���?��l��'�B�'���0��iu�]�Sq6l�� �!���hO>]؂N�3�<؁��4,�� (��M�1�itɧ���O@�O�dBE�D#��9����
����y��� Ah`�yf�Pc��aV��y��_�=Ijh��I.pv
�VKر�y� 5�Đ�ҫ�%>��������y"�8!5������D���FK��y�(Xqv��#�!<8���aE=�yb�A2��D�!0���z �3�y�,�"�&l��M-� 8�
���y��K�Rd�5ѷ� w^��e&��y�ƪ���2��jƖM ���+�yb�Ʒ`�(I�嗓tlԉ���	��yb �n�f��g@b�&��$�H/�y���8hJ�@�Z�:�sE���yR�̰~ě�D	|_�8���C��y�N�Q�&���a\(o28�a�N��y����UB!eP:3�R1�4"��y��ǗM2�=�QG߹7y�ItL��yB
�FZ�$�M�a��4J�y�)��bL:�JS��x��"�y��ω#�)+Q�A�;d�RaAX�y���� ��q6'�
�de�SA�
�yb��xE��"tBO(Nq�hՁ�y�F׫R��\+�ߤg8�O�yB���~hA�iVw\� h0�ʅ�yҪ� D<� M� vv ��
A0�y��=o�[$#Ԛo��ҡƫ�y
� Z`#`a��WE���I�U��:�"O�a�ǧ�"uArQ���Ґ>%�"O�aS�Y*�(A�0����Р�"Or���e��"�Е���[�(ov|�"OL��*�!Ix�W/z^�d3���?+M�9��Fz�O��Sf�޸(��Ibm�/޸M��'�p�1'ج��=:�.B�/����Gy���I�:��<Y��R*Y�F���-IŪq��R�<u�Ǚ;@� �f�;Q0��hS�Qh���d2[a���I�oaH����K0AA:�1Aƅf����DQ�
z\�1��#�yr,S4<:�j�F	�N��)p���yҡ?�P�c玥A�:�q`�N���'�p�'K�
=8�E�dD�
�N��w����><����yR��=;PPj��ޥE4yY��?M�A�3���6vQ>˓T�̤p�
� �0���Df�R}�ȓ�<������,����kw�����=�iAσ_��ن��&^�"��q��)�8��C�"\Of<�b0
����0����G�p2��U�Je�l�ȓS"M"�c�K�,e���K+[$5�ȓ]%xgD��zV�������Y��EZ|����"7zv���o	M�ҩ��?_6��4+��1r���������~��eG�R���e��B���_��Tc<�h�p�N�>N�|�ȓ!ۘ-���� v$>4;g���$����ȓ�<���*�s�f�u*��5D�ȓF/
���JE�,�
DyQ,àsD��ȓr�t��Ҋ��Q��F� �:=�ȓ����QLP�( ����G㖑�ȓ>`�\ɰ��5XCn!�p��(P��	�ȓU����D�3�@���͢[d���%�L�����7Hvp0��Ȇ~1 Ȇȓh�H�Eǜe�6H�oԖZ=����4��	�K�N��C�|h���E����W,�"Ay��[g�͒26�Ć���4r��@���;�cA�g�݆�2yYi�D�
f�m�$�x`\8�ȓg[�pc��
Qz���J�,��ȓ+����~�(���N�W��l��Q�$���_3�� ��ٓf%H��ȓ8�:$>Pd��⒒jL"$��O��yÕ�J�T]3IC�?`��ȓ;n��5���]t5��%D�c�Ja�ȓ9����+Ѩ�Y(e��
 �5�ȓz���P1
Pei�8�F�ޞCB�чȓEv%�!I�U�biZt��p]��WrQ���Ϣ]-�i7�ǀrJ�Ň�Z��Q�T垁6
֔�*��/X�<�ȓgT )nEϬ:h�AC��=e�A:�1��8�H���2!0
������ZDBc�X0BtPB�mc�MJ��_�/�" �f�%�6m��a�����S8e@'mP�F�z�{�O''Q� h7�K6R��*r��C�u�O]8����șKc�t�� +qr�R�'�����G���9��)K<w�4��'�� ���#y\2��W�z��G�$ꏇ��-;��0��n���y���� FT���84o��I&���"�(h	fL�����@�jB� �:�i,�Q�� b�M|R�ё��K<���u�-�O2��s�:D�vH��L��L_r	H��N:}�=j����N4)��)��d��|b�P�O�r���'*�
�(gBR��hOn�#��ܣ"p���R�"�J��ן~�q�Mڷ$"���"��x��mj�"O�Ѕ�	�[׎��C�7��̢��'���s��#��{��
��҉�	�.$�%Jbi˅��@�2%ҝcB䉳�*��mD��
��%$ֶ �9�קʊlPƅ[����:��Lhl�|Fy���QD���e.1���������>�ť
�0�L�� |ܺ@��k�d!Q��D�L#�h���ߝk��q��C2�p>ɶ��W�z��"�D}�sU�'Y�p���D�!^v�T(��O����'d� a���=��@�qɅwN4����V,�::�^��Gk�,����T�j�V:��e�͘��ȟ�4�ЈXC�q�ߥb�[!"O��8ƍ�{�
�VΒ�O<���voC�#\��I %�X��o��7�g�s�"��f	?[��p,�&[���� W&dD���p&�y2��1�,�C$�0 y	c���0?��'�is,�����i~�1D�
D�H�e�ޗm<�ML<���$>�y�bG?}8���NQB�<Aר�*5x<;eiƉ43n�i6+�@��¬S�f�����ɀ, �a��9J�*u(��f�!��O�	�D�Pf��0?�Xᳲ�I�o�!��? (��'�5o���Y��L�5�!�$ʢ4������s�����f\9&�!�'t�:��̎#l�\;q��!�D�*]o>�3rm��;P0���jΛ�!�[rD��@&N�2n>i����94!�d1&Rt���'"Tf�y�@�%]!�d�3ς�
��Ҧ6�l` �
�
-!��֐dB�؂��4#�{w�Ӳ2.!��DG������ �`Íu%!�$5M98����3	�*f��O�!�ė5Q�\I��HR�R�PC�a�(&@!�d�"<Q��A��&v/<])��L�!��Z�\eޙch�)�6`d��ik!�D�=4p�8w)](��3B!�qD!�D�C�����m�"[P�b剺d'!�$��y�8���A0z�`�� -x!��:fsF�!Y9"C���u(�yY!�$�I�
D!6�����z� ��cL!���$3�H!��oK�1��=��ڎ87�Fk��;��'���PɆY֗"9�zp���%�O�+��)�⽊���%;<��㜪lb��[�'.����T90-1��VzZ�)��I-{ለ�T�d�H'!X�Ա��ɇ	͆�'J������ϙH���ub XaT K0mH�QZ�$T�{��>E�4Ă$!h��@(1h�C�(ϫ��'�ԁ#�'N�b�m�`�"e�W�`�v��*OV@����'[�ayR�Ya�cG ٗ��!8b`��L��ѕ�'�"a����
�;"��S+�D�ţT���r&�N8��h�M��x�7+�02"��;�b��eM�YF{�	�4���ʉ�	ιZ�(��΀�bֶ[�SM'�wͼMy���dNV�6%f�[0�ѷh��T�����?)�b׼]�O��j�O����8)e��X1v&ܡ���U�?�� I��Ԇ�ɱp�p�PȞ�I�`���I����	Q���T~�'�69�aϖe���z���:p��X�
mc�=X��}��'�pYJ^c��h3�+_�Ύ���
2�<����(?��C6`&NYb��S�pi+W�4c@k��Y��i�v(�*�p�
�x"��/�y���0~`�k4��e�J�хg��L��)��'y8C1�حDN�P,��[�Z!��$c 5��Ƚb1�* �@{,̉�P[�r�Ԩ"O����U�K�.��V�p��\[b0O@E�D�S9[�p�Hw��"~���az��;��9Wl�D�G�<ac/�"t(����#�&0��B�H~B�3OZm �˄��0<	f@��=�@!�ɔ�f\ad]E���B2�C2���I6O�K���ŵ3i���s	��`�4��@�z���|�A�B�qyS��+����K�'2�B1C�2*g|8��T�\'�P���$3J���	gP���N���Iӓ\�&
0����7*W�WF�̓K AI���b5��O6b�۴�P5����]��A�Q�.!�פ[�hi(4��?m�h&��y$�I�{��hPL_�X��/	���[�e�(� J�,7@���SH�r���i�f؀(�����&͆}	��k�\ �H����?d���J�26�������|b��|
� 4��Ѓ #��Y��킘k��Ai��'�$��P*:�.�Z�� d���0'L�b�`Ov���N���<��¶���Po�-CL�K�"�x�'�~h��"�d]5T�mʰ�_/DY����O��%Ȥ��xB��2��%huEO\Y�����]$%���U.�O����PA,ʌZ2z 2�
 _sDA�"Ox�'C��e��Nؠ����X���M�O�J<�'p�O������ hn�ڧ-��f�~E�u�'����4e�J� T�I,H*n��#�3_j�OD�:�G��<� ��,�Ft��m�2�i��KN�'n��[Q?��C�xn�𡅞� �J�����5���v�_CH<Q%�8[�|p1\<Ö��FAByr��.t�<,�=E�to��V�H邊^?w����K�y�A��T�d!��!�\�Se�<��'�|��e;,O�H2���?�A�gB6\vْ�"Or��e(�M��	sƋ�OD�`p"O�)
2�L%̌L�4&�+1�@�@�"O�ڲ-Ъf4�0�*� Ȟe�&"O�xB&�+��y"��)9��́�"O�m[�;��=Pi��{�x��"O�Th�B��!��J�G�=� ���"O.��G�t��Fm�}q�0� "O0�"1.Qn�[4�GZ_�hA"O�1	P�pk��It,�9[�Ia"O������;3�H `�٥K=���"O!��!�7H�V�a��p:���7"O
 (���$��5S�O�!'J�hb"O$y:'ș�@��:C�}հ��s"O��m� ��2�L?*�J��g"O�)��� =�D���Mܫ|�d�r�"O�9ёI�a -�;%O��ҁ"OR$�p�G����pL*E����u"O"p�B��T~�2�ꏁG���"D�@�@�Y, `P�D����+6D�`JbH�.ڀbg�ӵ8�̔���&D�����(~I�@��Ѹ<�z�qu�"D����]/��DBT�ܡi`��0�?D�\!G �/f�u��ƌi�d(��m;D�ě���<��pq'G�C�B���+5D�ܰ�6SN�pP炧A��#B�2D��U#
V�����ܖX�C�4D��Z@�,$����E�°g1D�`���'$�v��'m�l$�2�$D�KQ�YRPd�A���{i@��g$D��@ ��3*f�	bi�'���p�"D�{��J)&H�\ Gh�;�Fp��?D�(!�ǡq�b�ղRzH\Z�A(D� k���.#F�tJ$��/R�]S�l9D�$��/"� ]�R�B�'��!M6D�0�Q�ʮN����%m&S�I�.4D��1�Z�JY�P�'���K��x �5D��Z���jE:��',��l�0�)T�'D��BT��h��=�R��uP*��`�'D����U�1��e��\12��"D�H�@/�{��5见�:6��IA�"D��V.��Qa:�H�(ؠ%ߦ���>D��(��z���(��5NKTu�G�1D� p"�c�|�X��(z�y`eI<D� Y�i8YI,!�ϐp@���eK'D�X�4��� u ��'�ώ>ԈFl2D���1�ޅ*�ȳ�̀��@��f2D�P��珵E3|1�Ȓ�[�(�/D�l#D&�=^�x 85!P�.T�%���*D��K�Nٜn�~��T(��ՠ����4D�� �9xR���e�d0�ed�w�D1Ʉ"O�1�F�N��f�H:Q�t0f"OjlT�	/��<[�j��X�A"O�Z�6\����w
ڿU�v�r"O"$�`<c��i�	R��`��"O�}�KX�3Hz|����60�F)c�"O���Rmȧ����`�]��	ӵ"O�I3 �@�H��'F�+��PI "O���aF �2�� g�"��-�p"O�5���³W�>`@�FB�W�8�"O��Wشbb�i1�šx6�`��"O8�FG�Ґ(�@��<B�"O�(z��ڷN�)��EC ��"O��r��<Z����e؋+䢤�q"O��肫�:nA�d�Su�E9�"O4���'�IE�'�$6��,�C"O*��j�-crB8�^aC�h	�"OJ����+E�Pk�ޖQ?d(Hb"O�@@��2K#Te!�	 $�%��"OQs�a��DB��*D�,5��d"O�l������La�-$�n��"O����)]2z��uC%Bі_y��q�"O�X��J��>;'@�}��Q��"O�C��=,�����Zs��9"O @���U�Y>�t
�I}��`�d�5�Ie���O~AHR`M�f���+d��n����'2VZ���:KF6����ɧm�:���'��q��E��{� ��1�
e���'Y\��V�T���!�K�4Gf�' <"��'.R�#�<'�t��'�(<�Ui��	�����4)���)	�'�N��b���R=�sa�=#-<�(	ӓ��'���s��!^�����޽DO\��'N�B��Z�f�tʏ<����'g���R�+���C��4�� ��'{B	��mP�3Y��RsA���~)��'X�yֈ�-"�4�*3B���'����MR�Bz28����\�'#���r��F48C�# ��#�'flKp�[�j<��۷��	�܍s�'݈�@T���T�N|Ѷ-	?x��T!	�'�Z��  � {er5֢��r�Z�'���JG��=>�*� ��ȼM�x!	�'�d���5|Ll"��D�7��':(�VL(<F���-�|`�'b�!p��C"]]�-C�J�\
�'ƀuj#Eϼ|Ɉң�Y�}3�@��'�nDbj�(����t(�rL���'ޚ���z�(��P�j�z���'A,��5�V"r��@��W�@�I�'�p�P"��\(9��P�����'֦Q٢o� dS4K���'f:��ׁ_$,�{+G�g��A�'Fp4��A1����)�!�f̩	�'����\�A���D��=\���'�����LT��d3��+��-��'�p�Bʗ��e���]3�\u��'��
p�F`�<�wm��*����'�J��VjReE���ǡ�!�xc�'�l�1��lO fLE*h���'C�\��N44���U�\�0�rp�'�荴B}"i���\� �x;�'EH�B�
T������C�����'�~�Is�$<_ꝓ'K'�4�;	��� �8S��\�W1��g�X�g�a�A"O�pj�H�Xe�3�67��A`"O(P&#�Q�8H3c�R7r�
@�"O��`ц9�RL#��� �LA:"Of�2��+�:l���6�d��"O ��
P�`���bႅ�����"O�a%/Q�l�ޜ8tbԮ8 � �6"OB��wK�8j�Y��_
�/�y��\wM����xָ��B�w�<���^H�R-���B�k���6. P�<��C��@���{WE�1^DR�@J�c�<!E�8vp������es�Z���j�<����7�YB2�Ͽ2�⃕g�<AF���~0��2E�� 7� ��^k�<��8fS���e̐�9D�
o�<���O�q
4bՁoCt���h�<9�b^�6І)@�G�8$5����L�e�<9�%��:��u�5����m��ENj�<q�.a���s �2u�=!���A�<I���C����o.oY����Q@�<q���"��$l��C�]k�I}�<a�J� ,H�j]�8jG�N�KD���>��|qa�-$$�s ђl`$���.���@7Y���*�/�s�͇���E���J�a��a����i��s��Y��כi#�)K�hO}��T��3� �Q����Ȋ�g��m ���ȓ[�x`�7)�TR�-��LL7>mt��ȓ"-L��&�Մ~(�귌��o�n,�ȓ�v���ƵR��,2���^�6�ȓxFY�살F�pj-Ir�ޝ��G�N)Ab�Ag�Z���)0��w�<Ae�nU4͛�i7�茡�'[X�<)pi22���u$��#!�u!�Fm�<�Նy�4t`�I*k5�&jSk�<�A��"�89�C[�"�e�IX���Oi� �׶3��'��
1*�)S�'7tm�����q�����Q�_�a��'r��S�3H- �M�(Z�4�Y�'���T[�4�
$j�!E��E�'�,�rX�s����E �>5���'� h�%M%s����A���Px��'�9@d \w̎YfJ�(�*P��'nxZ3$>Du��e)6���'�P)q��X.�&�
��װ�0Jϓ�O|<b��_0\)��0r,Ϟe��HU"Ori�� �n4���a���r"O$��g&
 :�uXPɓ<?3vL�&"O��Х��G>����G�`L��"O�r��h��pBӣ*b-�'"O�A�hJ6/�$]� ���
�
3"O���,׬	5���(ʢ�%�>�yB����<I�s�U?�ШG�T��yB	�BGv�H�ay�L�G��;�y�'��z� xp�V�q�v	B��y�%ʜv�䈷#T� �"�'F��ybFC2��Ѣ�iI�En�t �Ή��y�N��f@P��O׋?��� X=�y�tk�֖D��ɦ�ʏF��1�ȓ/j���N\�,z�	���J.����h J9�1i��XЊ�r�L�p�|ͅȓD��}X��ˬIf��?@6���X3�icAbϼ��X�,ށ+Դ�ȓB	�\ &��>B�H�B0͉=�B��S�? �0 �C�}���fC
�	O4�3�"Oة�C�Be��}�q�Z!g0nD0q"O85j�b��x���b���n)p��"O���/ķ%!�]BGi�>�٘�"O,u����%r �  �m�$7#d���"O�`�6�Z�:aB@����o0B�XS"O�0ˀ �"�8:�ʏ7A�ڴJ�"Oc�g��\`�3�T;f���"O���Y�D7pPȑ)�4'v��Y�"O�����סJ���qeK�El֥sU"O�9�A�_ |�Ekg3�Pj�D&D��xq]E����2ȉ<r	T�)w#D�d��\?#��CS��pN1�m-D�����-3)�Y1D��	�.���>D�����{0���FY�a�<6� D���cN
�R=�!�#i�AF@{eg2D��7��"q���$Q�	.f*��=D�\�a��RV����2�zْbN:D���R�����031�ˆ P���c$7D���gF�N�,8cM]�[�=X��4D��ɦ��$5i���'�Fp��1D���ch-!�8�+G��c\FP�@h.D���&��
�]zwI��7��B$A-D�,S��D"wn���#ؓt���R6-D��x�'g�Q$lp���+D�\CS�#)圬��Ҋ|�w*D�T��AX#`��J�j7&Ib�Jt-=D�,ڄFE�C���)�L�Y�~��5D�x�u�U�F�RE�SQ���4#� 5D��X$!�7�A�q�T��D�X��4D���Vm�^m8��������0D�H	�	�+]Y��!����A�+D��� �&_��y)�gU	ow�|Ѳg(D�D�"ƞ�;?F!� ,f���j� 9D�x(���%d����ή1���c3D�P0��
�&b6}	�!IB�P���/D�h	���6H����GL.9�F�z��.D��p����*]5+t�Bh0D��������˚�5�D�)�n/D�|�q�D���C2HՒ[rBh��(D�x7�L<�#"�ѯ5�$e�d�&D���Pȝ(D��1U푅k4�Y�Շ(D���u��m������<d��Wf%D�|:��D4eT���vh�8;>�]�w�5D�d+��P�xb�8ċ\$b���yҢ>D��*3B֟.)��k`.G8����H8D�8:'A<�]��OВ^l���e6D�D`�k� t���H�S8�`Iñf4D��c�Ɩd����C�+v2�m��$D��G�M�U�lPQQYo,eQ��-D��P�I�zP�դM�0����`*D������2A*n����I>jre��=D���w�X��	��O�(�ZI��=D�@��Ȕha��f��w�-���'D��!)+?��ٸ&"�2��r"D�HCg;�E�/ڸ4Xa�?D���v�U�(��t��䗲���q�>D�����3^^�K�@V�kC`MxC�;D�@#7LJe��4@#	
o�>)2��%D�$XS�?}��ys��ҳe�&q
��1D�8hKʙ�V�T$K�P3sSN1D�\����;l���!�	�E��\�#D�D���Ch��c�k�Q=�xk�H4D�"wN�*ߎEYac��X2F0D�� ��F@Z�(ŉюҼH+���"OFd�hA*�d0gg�7b*l�C"O�P�+
�k2FN�t�	3�"O��"��K���ԇ�IX��ɕ"Of�k�L
4E�<b��+�"u�F"O�)��o�?;d��4��@�$�""OԔ�4�ē5�
	�E�Ó!��\S"O�D!Y�-S�:).ʅY�"O*�)aùպ�;`O�)l�}c�"O�!�QkQ�5V����S���I�"O���"���بtFB)w� �"O��(�C�$�0��P�Q��Q��"O�ݘt	�)7 LJ��Wn�52E"O��r�(�*l�ЊAA
 sôM�v"O��4�;83F��%aP&$�t\�q"O
虅��}v�����X ���"O�%�7�1X;d�h�����Iy�"O���q��n��X�Q�����+w"O,�R��68-8Xiՠtt��"O|�0�U�Vui� ӄi<X}1"O�$!��G!F8���#n�>���(�"O����DK�g@�`k��^�g��P�"Om!�!�+2�����K¦,�2 [!"O���qgX�)j ��
͠}��@��"O�ĤX�q��:Bj
>�XP"O��jD6$���3���*1���"O�����/�\�A��V�oA2��"O��� #&`h3��BP9ڣ"O`yX�)_�}��u�ƭ�;$�t�t"OX!M
�n-�5M]	� %�"O��2ŏ�o�,Q��a3!�x��"OX��Ӫ��6�����F� ��"O���!�!l@"ԀG�m�:<��"O��1*��."���o��b��hT"O�Q��ڢc24��L�2[D�I�"Oެ:��Y�vj�A1�ˌe����"O��SÀ�0�p�5h��F����"O�����] �݀d^�z��PBf"O�u�b`8a)��JwE�-���S"O:��͖\}�Q� D;v�Y��"O$�)�D5u	������ # �"Ou�fƁS���o�>M쀅z�"OԵ�m��ixHlc��8p�}j"O�L������,耆ZY�jy;"O���$KE�BQ*Ȑ0��yi���"O�<�VŐ:"��x�#�؉F�d)�"O^���můe����[����+�"Ov���*��+"���F�_�/��"O�=rׯ��K�TzV-ٸ\t�8��"Oޑ���v���&��0�r��"O���V��?s�4IV��9�l�zg"O� ����M�>(P/\�M���z�"O��[E��6�*8��DG$-�W"O&UH ΙYŀ���,ǈ`8,q�F"O�lBTam��hIS΅�.���5"O�y�v�E����ʁ�&A��zW"O݃5+�wN�0y�i�b^0��7"O�|2�D��&��P�W˙�'�|���"O��A-�i� ���49Ղ���"O(���Zz
u C�ƴAØ�P"O$ɑHϦ(! �èNI�� "O��P"ǅ�T|�����#O�}k�"Od�xEnZ��x�0�-D�3.6-�5"O���RN�s=�is�б0�3�"O� r�yU��d����i��<	�8!"Oĸy��Q�%��E	�%n>��"O�%aƂd-��Ȕ�D�d��#"O�؃�+>U+�͒sm�W ـU"OԈKDH�DP��v�F3�iRE"O�A��Q=J!�P�"a���QY�"O ��KŨ�1�,F�L�C"O�%�H�g��ʱfO (��<��"OBDBm�2I�c%�(W�x���"O�	�C�R���	cdFW�v��my�"Ov����f�pU��3iZ��"OMauO?]�PŃ�H*b*<X�"O�X���&��YRtBS�9]X�z�"O�m��	:s����3��vJ��!�"OY�PM	d8b9G	վH��"�"O:���A���H �ݠ%1|�!r"O����)|����F�:�����"O�`ba�d!~�p�
��,�Q�"O(�� �A�RU��@�b�B�<�zp"O���B�V�<$}�2hՙx�H]��"OB��q+Ւp� �sf~�2� �"O�1��NL�I��<i��"4���XG"O�}QJ��̬��dFY�1y�"OU�J�vԚU��O,-h�r�"O$�riN�GbnlHdbCB|Lb"O`3V˘*SO�C2OC�1��,�@"O�):ӂ�om�)�΁�
�mBB"OLŲ%��m>����
�@8k�"O>�C�Bɲ[&�����y��l:�"ORT�͍w18�9�a��U�$��"O���׭�!�Ug��q�`0�R&^[�<1E��,,4V�)UO�TzzI��J�<	�L�h1� 3C���
�Cw��@�<���A�[�䫔 Է4�R=s3��|�<P$�n�&�Q6@E>4������`�<AV��
N�,)���i������T�<Y�⏌y�DJ��Ƕ�����ybə6'��p@��T!ez�3U��y���5/>5#!�b� ٨$!���y�K\!Qv�(Q2��-Y���9D�C��y�n�#0�6 aq� 6L��aj�`	�䓏?)���T��fԾٲD�H�.P�1b��C �y����[��av��'��Xa�D"�y��G2Sa��凃6�x�y1IX��y�mH�u B3C	ֿ�|�q
?�y���	���Í���%O��y�!U)N�Ւ0Lύn��r�	��y򌆂P�x�S�\6Ι�sm����hOq��@��!Ȋ!4F����վm�� C"Odi�4�F�li��.we<��B"O����ƾ$t8�N�:88$�"OJ�3����e��Q��ȓ�5`@�"O� �w�A1CJ���'A$b(�"O��2�kۦ�%��Da���'�B��y- 4d|��Gn�?J���`����x"NQe*�[!R?f-��`��'e!�Ϟ��7BݔKnd��m\5%u���8K�-�d�I�q��-&���y���u��8�% D�h�u�0I\��yR茾;��r�-Y<�5�'��y2��W���$`ƉDdybBf���ybo�%���kF%s�i�6	݅����'n�W~�埪`�bq���1�u�Cے�y���c�Z���J/7��0���y
� zhb`�	��|	P%��F9�H�"OZ��7
ؖn�R�pr�S+@b�"O8e�VL�+m�V����L9�����'���CJ�Q~j%* ���H�bu�(��0|�E�
�j�i&G��!2v(�g�R��hO�'�̌j6��gjX=*�kկ>+܄ȓv����S�Ϛ>� ���bI��L��.����CT�5��t�oĬh�>E�ȓs.M���YU��"�]��d�ȓBL=qwN�'��CA�G�W2��'�ў�|���fxV���e�)�%��9���lD{J?	 ��&cnP!B����j,��'|O����OZ�I�m�iVHD=4�z��׆ű`n�C�I����/�Q��q�a�D�c�C�ɔ �B=�J�m�m�f� �	7ZC�	�FC����86����m^;'��C䉈p�����(��I���cD�1!,�O���0|:5�̠Ic"����~��T�!DWg�ICy��O��qj�89)|�ruMI9�ܰ�M>�)O@��Q�i{'���s�<8`�LB2PE!��/�В���C�ݸՋZ!�d��j��ES5a�2.���*�5jK!�$�"pn��b��m� `)#��;!�D
W?�E�����Z�`A׺8!��glB0���D= �b#�7$!�ě�t�(Y��C�9��:��^q!�؞3Qޑ���ޏ��@A��~�!�� �A�ć4L����z.!��'�@��;�����"JB��d�ll�X�/>}��zԊ�y�*I���J`.E|�4l����y�É� fZ|���vgكWj>�y��a�z0I���q#&�Qֆ��?�,Ob��h���䒳~��:��Z�wR��/�p�C�ɋ`ﺠ���kY���IB<n^C䉧$R�����f�2A�@�fC�G�"���� |���2#
C�ɕ"�P�里QVyIdl�~�C�ɰeS�*��ҐU����F��C�ɯ2;��@���? !8A��4QԶ�=������e1D�\c�Zс5�Wu�"O@$�R��0R`7�nt�t�0"O�[���C�n�xT�G� fR���"O<��U�S˶��g�H7�"O4|�C&݂&ӺEI��J; 097"O��pD�D������B&��ق�"O@�$�)`��K�Q����"O	ٰB�#i><��̇�[�~�:�U�DE{��I�$G��2�3�����%:M!�$Z�^���@⋟(-"TkӉۃ�!�L�>q��i���gi*R�D4r�!��%D�9��2 'p��.M�^�!���wB��H�+��q���2��O��OD�� �I�&{d��@(C�G�N@��ǧXO�B䉅�V ���U� ��q��PThC�I;f����K��p����E�[^C�	:� p3@%�Z��aRp!�2f�C�I�i�4�@�� l"�5��JN4@>�C�ɽc4t�j���:�U�����C�I!96� 
��.=�x]HH��r�C�I�*�dD��j�>I�����]�C�ɑC��X"�&��n�ށ
6jX9�VB�Iu�����C	�н���&8&B�I�v�fM0��%FӀ�2g+@>jFB�)� �-����{, ݓ��֞I�x�Q "O� �t�M�Ϫ� 6n���P�"O0�Jt��F�>� ТҎ%�0�6�|R�)�ӝ_f�(�g�R.l\*HZB͑�Gh����*�	,�}�S픍u9��!���`���#?��L���EP(\�j�	�f�<	��S���w��-�� S��m�<����<T=ḇDb)���HQOj�<�g��|
��c�1LtI��Dh�<ɕiP;tVq(R �1O��0F�]ݟ���\���R�ҍ�ހ�
�1"�(�'ў�|zS���iwP�����(TBr�	O����<���8���O���b�o�OyBY��'��g��(����%�,q�����Py�\�kT�X�a!��s`��v#�#�yҦkTh
Bf�> ��w$ݮ�y�GɈdS܌�3H�"P���6�yb/����}�6B��blt�J�Q��?�(O��O?��T-8A�	�fWCh}H���Ix�|�'J&��!�M�>k0����5��) I>�����Ȏ����6tI�i���۸E!�䂿/���bN*<Z(
��\�!�$P���C�.���jU*	�^�!�D�^W:� @�x�)&J
+4�!�߅c�����a��d�p �.s�R�)�'O��{qK9[s�y���*?pf<�'��QG	<A�M�".��.�	�'V�]1��)�4Q{��(���{�'�l ���I�!�Vq)�%!��S	�'.�lc��G�v��&�N��١	�'�@�A��F�B�q�9Sn��:�')R� c#O�V��c�␺E�V@�'3��X	�(K�<-�v(B�J���r�'ܽ1g�3B$��o��kCH,9�'l$�I�N�? ���Yd��,0�Qa�'ߢ��3l&O��@�"�/m��	�'�8E�2l	�g��d�Œ*hC�5Sߓ�?)�O��RC��>�R(	�շX�h��#"OV)QEA�43dJ#fgp�� >!�dʙҞk��	)o�US�HM
H�!򤂡k�D;�F��N�e�ۧz�!�䝯]p�;�(ʗ�
a[�
S�&�!�D�Cu!�#�U08��h�
���!�DFza�Ec�h"a��(�x��}�����j}	r�ː`�4�,(3re1D��@�-������Ѱm��jg�*D�djՀ��&9�=���Ϳ7�U��g(D�,�v-ɋB`�����>��X;v�'D���$�@�}��AK��H�a�ɉ��(D��x( �Ba�=bF"�l|�#�&D�x��GAj���B�X-B�� 1�&D� �ĭ��Rb���Y�N��)D����W��lJ�-���R���1D���6���N���0i�x$��@�*D�L��� ��(�GBƅh|�9 �H*D�(�F-�#,��<r�oĈ/$���,D�$A��9,L5��;F�0��(D���wnҵ_��|��g�nzČj��$D�$�gC5���P�eh�Б��$D��+�g�&����8��:�'#��[��pB��P�b@L<�򃋵<�� ���,�O"�I .h���'�@:xc I�.}�B��5���mF��b8��f�v-�B�	-&�Hȱ0��#5&�����(��B�)� �XDNӆQ��0hQ/$8+�5�"O�����B�h.,���.���(A�e"O�TAà�(Q���z��ȅ.?�����	v���� .2Md�#����vX��:D���H�x���s���8Xۣ�2D�ԀJ��<Y�rD܁R���3D�((c!l�^Ei��ٳ[q�H�*>D�� �`�2�zi�*� 2�x�1��:D��@Ʉxɪ��íU�3@>�&�$D��QCʐW�f)����b� L�" 7D��;WǞ,F	 0�դ�S��U�P�7D��
f�$�}c�o�)_�I�@0��v���5���M߄�����a��;D�$S)X�#٘-��%Q/"d!�tN$D�ȡ��3-��xNI���4¥�-D�,��k5e/�4/�Y�p��Sj-D��h#�Xj���P���*Y"��/D���uNQrr`��)���2B:�$*�Oܹq��=@fJAᔲ�U3�a����'�az��]xl9'�[ �6��B�y���6n�����p�z� C��y��k��Yb�W�j���kH��y@�B��x�։g�J����4�y Ձt�V��`���c�"� �V"�y­R��\�[U�V�CFx�P������OF��$�/	��a͜{�$�2f?��O����C`�=S��� �F��fc�<P�!��2��4��荐S��0����1?�!��̣2�l�4J�8�j�p��.-d!�;_��K� �7t �H�D�,Ho!�RU��!��NcH<u	��!�E1w[��JV�XJ�0��E�W�!��ޯJS�Q���tA<9Q�E�(�!�D���#qdǁ)(J�j0��`!��2}�� �"��%4���	��g
!�OS�^1AB��
V��	�gF)Bўd��6zX`P�<� ���/��C�ə0˶��
͕s�4�(�L�d�B�I!'Y��J�,#}�'��ْB�=Y�$t�F�g\:�ۖ�Ŋk��C�6�0�S�T,J7bL��-�v؜C�I�kjj`9S
�;�d�{��7'i�C�I�S�tA:���bRdk�L�9E`C� D�0�9�� � @V�	k�(C�	�Hf����W,%� l��ۅ.-C�	
�����0Gi�I�U��MB�IDUXmy�d��/�����I�hh��D5�S�O�����!��W�^�Q7ό'w4 H�"OȽ�oZ(x
nу2�Z,�A�"O�(t
��@��E
�X��1�"O������	W!FF�9#�N��"O^D��V
I��|� $�]�N��"OLyXSb?] UZ�Z����5�'��	����zaQ�>9@Q@3mY�B� �	h���DE��'e��x�o	=(��q�!*Mؔ��'ޮm�3*��"��Y�����@��	
�'z0x�֏ ����@�l�
?4j	�':p�:w�L"�h0зM%3'�(9	�'$�M��G0{@P8G�P$�:�'|Y�۴~ڙ��� ����ybH*��::j(�
#l��J�H����?9��I��y��$=��t� 	�*� Pc�� D�8�"�����ō�5Z٪��?D�P��4K�`!�2y� t�8D�� ^��J,'���F��!��,�s"O\ĩ����j��%���$�,<[p"O��g��NY���dI���H�e�'�0O�-����Z$�"7"P%S6�$�_�x�	Vy�'��9�'D�*M ��AŒ���yz�'�8�*�C#(Ʊ��� �����'�p8�u��e��8�
���F$)�'�����	ߒ+��21�4�R�!�'.L8�g��g�`)��Dڀ��0k�'x����$ $sb3����o^٫�'�Αr0���i�:�@��U�-b`���'�B�'�RQ��gܓ����nکb�(�c7&J*�t-�ȓ#X(0� ��=x�­� �	��x�ȓ�l� O� F�F��/جA��؆ȓR��3��G�h#��	#��*7����?��\���)Ǥd���Ԣ,h�݅�߆�z�jڢ#&p�sw�XDԄ��	�<����N��LS��@�[X8,�G�\y��)ʧ?MV�됛bfA����A����U�er�EKR�4����hPFd��(��9tn�>&�IA�Q ��$���I3XK�`�Bʽ!�P�0LЂ{�RB��'c9((�-o��F�"c
B�ɑXxT$ ���y���g�:^��C�ɥU�0���H�&�*y��d�:=PL�O�=A�y�Ӗ���#�#y[d� �b�(�yb-� 1@ t�y��Y��թ�y�
N�m�� F���t:���䓻0>9���*Q����̐��1�BFEz�<)U)κ��a���ԌYR�(x��~�<)�j�3��������8�6��p�<�-Y'%��0W��290��CP��qy��)�'-��C�O7�l�9��d��S)�)���
���y��������ݱ�M�k�Xq�b�UІ��?iӓ"�NT�96�Ͱ��ҟ*
����m���⭟(\hHi�Ǔ;ɦI���T%��V�O�AydfA�
�����w�pa%m��V�ʅ��Q(gR��ȓ1�> h" ��G)�@*��L$j��H�ȓ�����7mz2�pfU�j��ȓ�����b���ެQ����:��ȓ>����@�|a�1�d�ݜRUv���uP~�9Ҡǃ1r�1F2Q��)�ȓ���kX�&�9�� �7V�ƍ�ȓ�L��Ŭ�/}��p9�%�0D��d�ȓu���� HO�4��"�D�4)������rP��do�t�p�W�r$晄�Ob��1��V��L⦍ё*n���ȓ)w����.�:]�Iʢ&�D���ȓQ�0��#���U���T�����|��p�L�Jmƽ�� �3����\�LݚJI�KZ��O�0b�L���u����n��S%8T��S�#�~��.D�dY��-j���ز�P)�F��w�B�	�J��i����i��e���_tB�I.f�(��nD҅Kd�A�|�0C�	,Z!�;�l�n��	��ۇh%,C䉼�}�Rƛ�*��+�	F�!1d�=�Ó/ݘH1��J� D�$X� ����@��L�����h�0˛�1��:�E� `�:���-0D���k�<����?(\��F/D��YC�cL ��iU�C8���,-D� K�cȦ\��-1���N�(p��,D�� <�����JZl$"Ǎ V�
0"OHIʢ	�P�J��ƹ���g"O��Ʌ��g�舢��c�$0�"O�Iv�P�
���4lՉ.��k""Ox�K�Yf���HD��	t"O<���a	��݊�!ٴߊ��u"O�]C��yv�EЃ@Û6 ��"O���p.[��ȃ���x����"O��3�I�K�n���X�����"O�zh �'a�\�0�@�E.ࡇ�|�'�Z�X���o�2�3ъы� 
�'3jE��� m��-b��N^�i��'���{%�|���Z�.�G�� �'^�	��͖W��(P��<r�Z�'�$e󖌛�귯��}!��'����ɫԤ%@�-7oml���'� ���I�sc����V�PeȢ�'��y�#P��Q����C��yQ�'� T����,��gT"9��U��'��iK�O살�pNW&1p�'D��U䈍{�\8	�8�P
�'�D����mD�XǪ^+�$Mb�'(f����UJB��a��^�+��,�K>��`AR��3gA�*qB��A��'[��ȓ=����v�G(�[!��}6���ȓQ��,ŔWު-#�/g���ȓA��-jѯT�,.(�dބA3���ȓ�9sY"���f
�
��Wm D���$��E���aI���Q)��+D��`��E�B)j��i�2r#��O^�d>LO��j�#�?�T �'L�ۦ�!�"O����C�Lt��s'��u���kg"O8����;c�d��4&�;� ��6"O�`#���6~�P$Q�/��i�`��{�O/l)f% #�Q*�C׼G�BYK�'raQ��H�14�11-�@���Y�'�2�۠(NX�=��A�g�z<��	L>�jF[�W_di
7� u !�#5��V���r�k8X+�z���)�Z���'D��SB�9������ބ'�Fh��C0D�X��f5h�$V�#l��QR�N��y���'��PI�gʝ��c���y�	Y���Eñ å`ʌm��N�
��x 	�w!�m�f�Eq�P�#n��џ��IF�Oش��b�/fm:���*x�"Xy�'�B�yQ�S�ɜc��F 9~�S�'B��y�d���$!��4iLP��'�kr̀�7���WLE�,��i�
�'���(U�_�
y�;@�V�h���'ژ�Z�Iں�� ���*�d䳍��>�'�(�W
_P�vP�lˉNuv���A�zI93�o�A˖��D�^5��
7U��K�6�ꦇW�{q�ȓ.���	�۾Vv���o�'m���P�h�*�Y�ˤqJD�˘vJ
���IU�'C��������0p��R-C�i��'�tA�7�B2�\	T(�[P���$0��ua`�:B�Al��2���}.|�yE+�"n&Z&吺X�5�ȓ1��cΝ�J�]	ǡڲ.��ȓ�ݡ�@3֐R$F�5�u�ȓ(��� �n�6H@�p:R�Z==Md��՟��?E�d�ɯT���H6�'P���Ѓ�߈�!�d��`�Ё�%`XM���P�D�ϓ�O� ��a7n��m���qY�g�@�"O���#�+(�!�T��5#7"O�� �V�FT��I!
�PM�e"O 
ĭ���B���+4z����"O���,V����
���8S�"O���*_�>��H�~��,)$"O֜�6a�x�u��z�r,c�"O�Q�@k��>�L�yVƈK�	+S"O.��gc�f	n&vt�8��"O� ��$T�5@�,��bI3Ch���"ON�Y�J٠RX*l�'f� �R"OxAr�3M}�0�E�Y˂m�"O�����,�21hvHǙ/�0y��"O��"�'я(�������q�w"O�)�`��2=����`�"`x�Bb"OB,P���`�$]��N�K�LQH�"O�`ѝE$ꅘfnD��D��"Ou�5�B?O��80�]�;0Z�S"O�
�m^:7�$��D�������"O��(`��B눭��J�Jl` ���|��'��!�gޫF���.W,1d t�
�'��u�� ],E�0��� 8yv��'�K��_Z���P�V�<Z�5Ɂ��m�<��B6~���$�	� 59�i�e�<a�O B��p��;T��9"�I<T��*g\65p��!q��h��PZ�B+D�ӓ�6�<���N�(���pi'�<�ON��G��oY&�@SmS7M��+"O.��2��8��|���6` 
�"O��[�	B>o�`�ֈ)�dy�"OV���-��N��U����;g�tLs4"O2�k����I��ѐ /H&!��A"O��r��4�{ulI.x��u嘷�yr�G�V�\���s���्J!�?I��0?!�fC�4��9�nյ���!��n�<a/ 5�ܴ���\�f@Z�A\l�'���t�h��N�56�+RCO�:6��:�ļ<�|�O�	&OQ�e?�Q��U
1Ϻ���"OH��24fv����;s,�9$"O��aQ�D�+�0Y��W�LP�"OБ����S �y�@E��<��"O��e�E�G�4tJ#��o�j"O�u���$"���3�M,i�,�S�I�����f�O��4���>�и�%W�-; ���R�'�axrHH*?��Y��P!&�\qF��y��R5�����E�$�t0SP���y�CM�X�6�z�,I�����ޤ��x�	{S��֎�2oR�:�/�Y��'|ў�>u��D\
x���FFb���0��O�㟔D�$���BEd�K���!T��-QƬ��/ў�'�"�ɑ\;r� g %�֠��d�����)��&)+������8G�K�����'��	�ƌ�N�\�+ge[�u�0�#�'�&�B%O��D�F�\>���'��P�/�'!{)ٲ.�)�Ҝ�N>� \��`�Ǵ$����@E�@����ȓt7� ɢ�>,p�"s�K�HO
TE��ӯ�$Sq撱]�(9��လX6�B��p2���À.\X���lhB��*N]!��]�Ph�����30B�I+"�Xe����2H�J�0��y="B�	2�R�[b�^:l&���ʖ.-mJ⟰��I�M��؁�ܹU��X	��ݸ*S B�I,�����ޓ0if���m�$Y!�� LZ���*B����d�Ψ`�'��O�}�$�!3��g�<E��ǖ&i�j1��8���y�E�Md�1��O +c L��|)���JP$�lX�DQ�.YJ���<B&ԉu�ϔ��a:��MN*���'�L%�`��­p`�A��ܸ�'P�p�L��R�d!`�Q={�X�R�'A��4�Q�/~�8g̊�LA�'��$��/ҸB~6�f�E'���'x�x�V�^�z�heaC�³e�X�
�'LJ����Ƕq��L�-�1g�9�	�'�t����K��h+n	,;B1��'�����剖c����␆���
�'��qe_<!@��s�)etz
�'0�\�������P�iH�+�p�	�'�tD����	�[E�ʠi�,9�'O��*��@C�I�d
�8�����'����@	�x�q�4� �+�6���'6@Q7�̕d�����5��Q�'�j�y�k��o��}�e�#1`}��?�K5j!r����E)4�X����y�d�o�������nI4�s�_
�yR̉�W��4'�^M�B,)@!�si��اF��VTBEi�`�3@!�d�&R�С5��c�.T� �[�8/!���&x�|R��2-�t������ O!�$	�sdZ�e�]����f�0o5!�d�3*�Z����q	.����z�!��_.q�pu�@�?��� `�M�D�!��F�n�x�S���jô�w�HR!�K��>A��_E¶5��X	M!��S\�P���H�,�z��_"!���t�X�S���M����6N�h�'��_>����Ԣ"D�����V��q@c�>�D3�O� ���#f<�"�1t�~$�"O�Hj�aQ�8h�ժ� �^�@�33"O���v�:r�$��X�/�tu3�"O�1Cq퓹ckpX����=O����"OZ�s!kR�xԮi լ^�z �A"O�eX��ͺ2��jց��f����"O2���^014uKP��ex@"O�DYU%��C��$���=8�
�j�"O�la��{=���mH !��G"O�Tô�
7|9B��?���t"O��Pe��B��m�GB"\,�CW"OtyȒ$
�F$�`�1S*�Q�"Oظ�,ٲ\���#��HE����O��	kd�	�&��Q�X���JӪ !�d�1��AHQ���8@Z���+/!�dT8JI.���nen��`��0y'!�$'OS"�#�H�u�
I���ٓe$!�$w"�m:��$� $���O<u!���������.VZizsj�s���dZ�J甭8��Y��-r���(�䓌hOq����T�)�Y��3;T8d@P"O¬!3���1w>�R5;�!#t"O*��FlA7VjL�F9i�,h�u��!LO�ԓB�����{s��0a1�"OT@���"Vx�Qkƪ�$5�`�ps"Ox��61e�̈[@'W�U�֬!v"ON��5瞂tRh����ɞ��|��i>��'M�u�@O��[���8!��:H�1��'�� ��n0bT�PG͉��@6��$�O�⟢|�bjB^��!�@�><�����S~���0=� �m���B��-8E�!\���9"O��U(Yi���1WD� r�
���"Oμ��LUH�h���V�9ܬc�"O�Yxե�9?ЍQ�C�'d�< )��	G�O���V�ۗ�r@�-<;���
�'5��v��:ʈS�FX)y���+O�=E��N(�.8K��N�5Y 0�Y�y!Y,�����O��<Z<��7j�;�y2��~�i�W�݉/'�u��I��y"�\�`ڦ�P�.�J 7��y퐓\�P)�%]�9������0>	�J�ܑ��-smDQӢ��r�<�7�(7�\0h%K�="�H�'��x�<��ʜ�kg��)��j���,J^�<%ߓqƈ�"h�m4 u˶	X�<��+I�~{|����d��US��I�<�DĔ rS2a"V	X,F2�;j^�<IcO�)��� jĐYո,�r�SQ�<�ѪA/���J��E'jAz�:�d�<�d��T��6��!<����`e�<y��3���]�J'h��rE[ڟ�E{����>r�F}X�H	(s���N��B�;H�T�1���(B(��Q
��r��B�	�W�\�{�S<�H�hi�/B�C��0��C#�;a��mHT�����B�I�b0�5Q��1|�%��25,�B�	�a7��0��E��,�"D�4^Q*���IO��~�"вm��j��%�8p��8�yZ�VI�Ŋ�a�L��CF�0��ȓ+DF�y��.;V�d��H�x��N�D���F6k������6���ȓj0{G��2~D���[~��l���hQ�#9Hlq{��XU�� ��C,0E�7����zgL\�orB�?9��0|q�h)`!��-a(��eݒ8.�4��	5)� x�s-ϤV��]�d�&2��B�	�/��D�W�@2��:rE]�B䉣o���qs���B��eZ����pB�	 W��l"�判:DZe��!�7iCTB�ɮd�8�K���U�����N�V;$�#�Ը��/@�\�Z���g���.D�d��a$jH��#t�YU1��ȶ�-�d-�Or���aI6:jD���e�8
��1
�'��т�#ǅ{:��2���H�%;
�'�`�`i7�j�Y�,C4F�R�q	�'���D1v�N��Y�9nr���'Kt��wD�:
��֖�r+O��(<OL�I�G{�-1�Ct+d����{>�B�	 {��X�L4S��K6�b�C�	�^ ��3J
�>�z�
��-f��C��w� S��#&_f�uÆ�9h�C�I,R�(p���b�,C�&H�U�
B��4�U˄�M�X�gG�2��C�ɱvX�)����ur�F�8����/?�Bm)��{�K6&�0��u�<�0jб9i���/n4����r�<���>��i��N�an���l�n�<I櫙	-�(E
#�$%��sqZe�<��2X��I�r��(lc:P��kW_�<UJ��6^�� �!.���C�D[�<Q����"�r��l�%f;N�d�<�?��I�U?�����>{X��M�[�!�䒽(֊��U%��	�%�wlD9]!�W�$�֨�&J[3��!+�;�!�� �;5���	��� �N�u�~Tc�"Ol��S�ѣS���@w�I'{بK�*O^�KVl�H�Ҡ[���/�����'���)�D�o1�a��1-Fe�
�'��8��$z!l�k6�
�%��e��'�8��Toֱ�\t���1Z����'�V$h��0v���; ��L��'��p$L�j�&0��O%���'� �@���%�JT(0�\!X*1��',Z�Q��]�:*.�ӧ(�-R�DY �'K�Q P��J 
_�fW1��B�I41 �2�IE-r�e�'K3z6dB�ɉu&\�R!�5?X�8�	�'�C��:s¦8y���
�T]�7@� ^�B�I�6n`�(�)�u�B���R�B�	�|7p<��$�>�j;F$W�B�	/V��k�m��*�V�Q�O�5{��C�I�dz0�����t<�u����a*�B�0I:&M�u�� � ���&%�.B�2�A�q��<u��)1儭VC�I� n`�%�Z����!�c
~�B�	�~8��4FB.��I��FL0B�I*�b���	�,1�X4�����D��B�Ɏ[�0��j*i�A����5ݮB䉅i��E:c��)��@p�@C Y�tB�<d��M �YxܸA�g��>@.�C�=v���pΈ8Cy����߂P�C�	3�(P;�#
��D3�87k:C䉼X[ZȻe� �F0 ��2K��C��Igx��CZCk����T�"�C�ɲ?�$mكg�#Y���<|����"O�y��IM�����\
C^�U�"OD���L�� d��&B;Y��Y�"O��Ʀ�##�H;�$%R�NY�"O^�$�06�F���)xH|�A4"O���(Y�2�EY�V�Z "O�M!��]>�T�rBd�+Y���j"O"a�Bׯ�`t��f�F8�w"OԹ*F(�5 4�q�A@�,�����"O0SEд; ��c��M���c"O�H�sh�la��ڐA�)��`�"O}�'*H/�t��\�?F�q2"O��"&��4<:��1��L�R
��� "O@q[��҈U��i�&�2�DԨG"O
�C��7%7^!K��	�T�R�Q"OFt��
m|�v�W&>�,�"O�
��(E�Z�C���$�Q��"O��Ч��a���Q)_�|D�Pd"O���)��z�֩S3�`�(�t"O�U����4|Xŏ� �V�"OԄ@B�R4z\PScZM�V���"O���Q	ҔPa��w��+�"O*lR�
ňƥ���4\�Zͺ"O|�$�Όh���J�+	rt2�"Ojċd�փ4db���+��'P3�"O����?A$�m�	��O�d7�#D�d��`�7Dh�R')�`�����;D�èƒ7��dbF,�'p��x{&�9D���!���Z�ȃ���j��%IvA=D�ld���g��$�Ɋ`�����-D��cDFT<e�:Q�ĂBvr)�p�+D��ˑi]�y��Ȳ��#J��H�)D�8Y3סM��%�=*��&D�
S�Z�T6٘g�<dVa�V�>D�� �������*A'��<tp"O�xr"!����$bĤY�{�l�""O�c �pH���J�C����"O8�8���l@z����!�a�4"O<Pq����yy���%t,�b�"O�A+l_7Mc�@���!da����"Oyz�I�.g
���Y4K����t"O�p�� d�L1�1GL�����"O�	ckͼeZt'_�rn�� �"O,��%ʀ+v4J��@�1��Lؖ"O���7�ˆw��A�NP�D��1	�"O�� �S�+�� ��<Bd�cr"O����N:SΈ�&,W$��)��"O���u��*H��ґ�̾)���(V"O��+�-O\8ظ+C09|)�0"O*7$XM�T���iL�z�
�;1"OdxWM������E� �����"O<�0�C0p��!�!�����"Oh"��Jo�aS'��x�H#A"Op�`%��<vƅ �a˂)#D�05"O��v�ġU\���,]�v��%"O�XD��l�y�I��g�D(�3"O&5qCaH�l/�闲�T�*O|a	��W$t�#ɘ|`��'�Hݙ"\'.m1��]�|����'sbm�Pḋv�BU�w<(@�'�h"7�D�!�ppKcǎ<�Ƞ��'�<�8��>H|�h���.p�XP�'ؼe���&i���gƹ%,�9�'/R�á�ú,QXU@�I��|��'bp;�f�1i�N�8�b&4�2���' �ARtK ����
&(0����'c>-��(�nH���(\01�'��a�ӆ�S�*��6����%�'����C�T�nF�Iv�\�,�Pb	�'Le�7��;��hu�6�4���'{�h�Ǭ�I�����O ʂY��'�
x0bC�\���v	ǌ#t�2�'4FDPBj(FRH�4�K�<[�l��'��Q��mB�-Fr͡�G�9��<�
�'���#���@ �C�͖.�ju��'��=i���4e��s���#"�)��'��XD41|2Ċ�B���8I�'i��Q��m��`3cS#9���s�'�(���NI�H۔�sd�+A&��'7#��CvR�S�@��Le;
�'ǘئL	2L����r�ѓT�3
�'*fe�"�W�(ȭr��4Vb�"�'{�AE��T_��X�m�"Ta���	�')�D�++Q��\��J�O����'l�-�p�ӡa���*�<0d�{�';D�YW�P������9�'(1�B_�j�����D̚��
�'-`��$,F'W�LJ�a[�-��D��'�pjrH�d�0�`�_1'`H�'�����1�Nx+r��a@�'9 H�D��)nz���%��J�'�b`Z5N>�N(I�B�5����'|�9c˨:���3W�
��xH��'<�@�ZJ���6Ot�H���'���S��kh:�S�!Y5\U��'I�Y���Gi�!2��&&�\Q@�'
Y�Ή�^�j��T��*����
�'�������T�|@P��X�6�f5�	��� �D��K��t|E�!'��"��EKr"ONP�FJ�Rph����: �:��p"O��ɷ�56zYХo�,��A�"O.����'N�]�%�_��L��"O@�'�˦Op�H���~m@�"O ��̀�A< ���"T�}$"O\<�3N���2��:V��t"O���RL)tv��JV,(�"�"Oh�9Q���T���0�&��:���"Ot<x$��1}��%S"g�5$h9"OB���]o�桩%�X�"O����]"J��Y��
Sdu8g"O���	ǳH�P�`'eȔD�*d!"Ot$:ďX�S"�ҦFxNAH�"O����� �q��
��Q9�"O2L⁌�U4jq;����!,����"O�a3`���J���1��3B:Y��"O���0��<�| ��K\=:\�I"O�XB����d�^82Te`����"Ol��f���y3W�ʺWV��g"OP �׭��$�C��A7����"O��!�J�t���瓀-�Xł"O��� �W;�Z��vgV�J����"OQȤ�^�����PE�^�R�8V"O��� !Qp����13uJT{�"Oi�b�ڟ���TAkQ��aS"O�`h���&����č
�.p0�7"Oj���Ɨ|# ���bO�*����"O"�qh��^��Qpe'VV_�x!�"O��Z�F��i�\`Y�� $JJ`�2�"Od-���a4 X��I"5x�B�3�S��y���y������;�"`�"�yb�"��m)n��8 ��9��D.�O�%�'F�>a�b�`a�Y9s���R�'*�5�m+4P ^gUb�e�7S�C�	�xSv!�)݌b��(�C٪g��"=Q��T?��lE.M��(�̞>[z�1� D���gJh�@ ��0bu�'g?��p<1�U"RL�@��S�E��O�<� �١m0A�Bʄ<<% ��Vr�<�k� J�p-�$�ޤ@��srdF��A���Ԙ� �m�N�l�sn�/M���/&D�<��M�c"�s�D�1vlVK���s�IҦ��_�g�Ym$)�RO�3/����元��E����?I�i"Prb]��؉5(J���
�П��6�	��hO`�C$]4d+Z���2.��qQ �'�2�'A�%�2怇\�Q(�Ûh`Lc�'8F��	�s]P5����Gk���uM���t���I6���ƌe(Ċ`�Ɗ�^iP��:c!�ܧ4�J�ٔ�����x(��5,-�$���$�<D���,(�ֹ� e�e�kbj΂�ybDSu���Z��Hc�p��R
W��yb�O8����e�,s>}Y���&����d<��^�:L� ��6H/L��C��*iXI��]�x� ��!������V�2����?��V� �@�Ĺ@�𐰭L�(z��� �d!00@H%79yPr���B2�,�ȓ����F�24s �P@�G|����I�x�׊F�a�&�#0	M�oIT؇ȓ���c�Wf�X��Ӂ2�~Շȓ=��-��E�:��U��"����<���	@;@�h-�C����1c㑟�F�t
�
'
8Abɏ-[�dZ��1�Ox��d�J%�M��W;�`-��� �!�� �<ⓠ?��{���:��f"OX�a%ƴ N�RfEQ��v(�ºik��$C�ۄa�f�D!f����v �W��z��x̓[�ؠ0�^yU!ّbɠ`��,��M&-)D �'ږ�`B@9�~��>a����'�n�:�p�j�X�R� R/�8L��ȓ-�,=�BZ�e)�@[���F�>���`�� dL�
9�	�s��!�\�ȓR/rɉ���9� ��W�,* ���F�'������*o� E�]O��q�'wtsW�Ъ"�>J�'�%FK��i�yr�)�2"v̸�����a�FO�!��B��+��C�K-$���݉�#�>.O|7-���0<�T��^��)�s��e�ĥ)ƭL�<y'G��E!PA֌��]��rh�Ħu�R���df�0�Ry���Νj0�$� ���O�8��"�p�C�'69�P1�	�'Vڕ*��B�2%a�댍+P�=r	�'e0PW���bv��m0Kށ�4"OxH"G�  �t|sB��� �"O��XPM�@`�╘6�\�r�$:�S�I�=�P��sJ��0I�h��K�!�|&�}SUi���{whݿ�!��֙L۪e����!{� ��g�;%�a~�R���&�G�h	<0���'�*�JK6D����$�RJ��4Á��!�E�O�'ñO��i�� �
�xM�3�B<�Ե��
2D��1�V�_R���E@�x�r�2'nn���>��ԟ��s���2�∺�	>^�̙�"O�ARN[�!��{�f� �uR'�'	��ĲdL� Xk��H�M�.t"<s��&O��=�!l��o��iZ��lF���H�}�ID8��� �L��H��������Wh8�O��əh-���;"g0tzV���Fy�C�I�G�H��a��������+p0B�ɝ>`T,?i�5�!�B��!�D�l����dB��H1ꇣa��y"52ړ���#ʧ/@e�54n@�`����3�ԙ��elJ�	�'�&z28A%I�79h,���h����ѐs�b�pp/�6Jlb`G|��S�f#�c��!&yv���H�+N{r˓�0?�@�>n}��%�|�ĵÇ"P�<y3�O�P�`tOչ:�0��Ai�H�<��MV[^`<ç�K���୉K쓙p=�5�2XJ�E����RtT5#2O_�<�᫛i�F���AXX��fY�<�!��1��ؔ-
�|h��GW�<IBK�+Wj,|�EL�R	�Z�!�n�<��
��o�6�h2����a���c�<Q.@�B��Xv�R6�LDs�l�J؞��=yA��(0�p�Ib����n���
]H�<劏8k�:�铒�䁇�ZB�<���7mH4�m�
Q1��yD�|�<a���4����$aH�)F�w�'��x�陚s!���u�ۑ] �٢ ���yr��	9��h��L�q��Dx7�9�y�T,L5�S�es��f���yN$zL��y�h� V���km��y"哞=C�ɒ�A��d!�"�n%�0<1��$�[
���'��k��؈�+��Eb!�� �&�	� �#���S�s!��� �ไ��:�Z���b��;X!���
��(2��fz"؈�L8@�!� !��ҧ�$h�zT��x�!�� �-��J��{��=R��	�i�� ����q�O:�y��Ұ�dI�AA�=d=���(O�ˁ��8�@�ʃb''m�-���ONyh��)�'|q���7#0 ~F��Ď�*���	g���9��]#=l�`��
G�C�I�J?T��AU!$�]`�H�7����D.ړl.���H3n�����K����I��0yXI�$��Y[�xY�	S*^��]s_� ϓp���
�S��<��Ope��Jߖf(J�� ��3z����p
O@6ͅ3^pж���e���`*�5m���-�O��F��6h
5ᱩU9u�iP�I�.ʑ>)�I�wJ�D�0��!L� !%�<��Q��i�Q�%�x9���[��)&�$X���)6Sv
`p`�Z��S^h i�"OpY��(ܫ9�4Q�S��&Hʌ
ґ|��$|OԱ�%�0i\F�7�ƢoQ��!
O6���X���j�)�t�Aj�
͏���Iz�'�\��W� ���� a��'QR\�����O�"|E�Î9	�X�[�ʐbi�a���=yQe[��z�xOb5"Z�<�"�	�(����sB��j x ��X�<��͎��F*�HM�����7��^�ey2�O�bd �S��`U`�%_:����'���0���gv���D��EdL%J��yR�'�����3�	�G|�y���^�g��hy%��/0�>C�
w;f���D�F��p�5�X�C�	�y6R-P;B�ހ+mۗz���'ֱO6�kh7���s���`ې#z�ԓu�K�#��B�I	�0Xc�i��-踸��ʖ"�|��H<q��$ڑ#��\��4y��Q�C_���xba��c=~8ae#zV�XKUɅ�;x ��~�,�c�u�'�.�It�X	V���Þ�"@̀˓�(O��r�:9��A�d�i��	�e"Ozq��(�,-�%#Q�Ǧ9����V"O�4	�nڄo;�PZ�"�Xa���"O0�q!�Z�:{A��d����"O��S�`Ƃ6j4� T�J��(�V"O�e1f-_^@k��M�V����u"O�y�,āՂ�R�V�z���"O�����]����"�K8\R7"O�	��׼�:��"�K+��Q"OH1����;�L���+@
0�:V"O�9
�F�S U�q �X���"O��9T@e���Pԩ�a����"O\����4-m4E0�]�I�a�"OiL��s]� ��Sl=�ykT"O�B����0�X)5��aR��v"OP�����}K�(-ܔ�p�\.�y�<`�0�P'�8h�G��y��W7P�D�4Ć�%�t��+��y���y]H�X���(�4"�#���y"
�!;(�E+��95����#��yb�Y�6UnmH���3
e`E�p��*�y.P?^,����B�ڸী8�yB/`������ �@�&�J�fʬ�ybϚ�.C� ˱&��؆����y���X�̨��H�*|:Pk�$�yR��$kg4��4��U:0��.ʍ�yr�6��	{F����s�_��y�$ 6%��aG
(n��Z�,]��y���Z�&I"ѩҠl1v0c���y*O
z���#�aĨSqԅ��$�2�yB�\+$���x��rApQ��y�l� P�f=��r\z$p��y
� ^ݐ�ۃ\%.3��ȅ5�$u��"O��HR��Sr���/޴_w�����'�^}���5�LAc��&�b�'��=�"!�'���b�(E.'�����+�(xt �	�'���P0ʙs#(��Ge��0���
�'���HZ�?�E�$��+��T8
�'0�̨����JP@��N�"º�	�'���S�5jD �@�u��|��'LM��bO����n Q�����'�5pO� ����_�"\(��'g�AӡJ�#�J��r*қ-~�j�'�Е�6ˊ��z�-r��i3�yb �_F>q�Uk�mO�t����y"G 2:��+ ���9�e�U��yb쑴s納AC�7Ox������y2&F�&,0�pF
�=��U5j�=�y�J�]"����W(��)`N���y�l����p)��(��P(����y�L�O�����\/zO\��V���y�d�i=�V�$�h��j8*<�C�	�.�0��S�XPUH(yD���B䉋zH�`R�
�t����I�sl$C��:y��GƋ؜	Xqh��0��C�`�c�O��o\i�A��&C�	��*(ss#m��2à՞vC��>^�\�b�����=r@G?���<��?R`a��ׅ`�U�TG��}�:�����yBМ��  ���Bfqc��sq
��P�(�$���>�T��<X�»k ��1���3���a��������C���H��U�6�ȸ3�i������0>)�cZ�#+M`D ���́	�lx�D@$ ����б@�^,�?E�SS!bDX��jqzGS�<I���{�r������ޜxY.V�Oh��Wfň$0B����X��H����Ag%QLV4[!�ѠN�� ��"O�(�%�6=�|8ăA�/�JQ�#���]>H��I�<�	Դ>ޱ��'� �Q�� )̶�[b�MrhH1�'�ļ	i�'V�|`BeP�\��+"-Ѩ3��L5� X	���'�N�`�)��8��*���+f��Ǔjf�P��Y(p��]˒��M��mUJ|<|�a�H�suD��!�d�<aWj�X��0CEZn��e��]�D^3����K�=�RŘ@K?ҧ��{�%ۙ+�m�HG�MFh��X���b��$L*���^�.Ӆ͌-�pP��'����s�g�I
P��UrnL9+9�$��=30C�(Y떹Y'�Z�1�Hu0e&��R� [�)��s�=Hs��PcL��	)JV`���-ŧT*� c�+X���[��F�X�l�/cR�ST�'������e����Q���r�����'e-�Չ�_���C�/�1[40�J����B�;`'�|Hf%��D�?�qA?O��@(āE�RR\!7I"D��#�7&x+V��" JD����8�pk�O���QN�g�I+ߔ}q���k*ĉ�rN	QzB�ɲk���ٴEϼ8����D��\���ϘLZa"�F,��	�P�M�ay@�{�l��y�o����
�¸cn��	GI��y2�B&J�h`�J�W�8u�c����y"Î�D�-
��[9D���q���y�ȅ�r�J 2�f���5ɋ��y�O_�Y����RM��ve�!"`��y"Ͱ�q+#�g���m���yR��ZT%۷m_ ^�Ľ��%���y�J\�r� |�e�۪V0��BB���y2�W�z֨P��M_EY�@�e	���y�/ב30|��00�e95�1�yBm�6О�+b�ǰ5�j4�����y���|�,X�F@�)���A�9�y
� 䔀%e��:��
�
KZ�Y�"O�L�2�@��V���ě�#��h�"O�$���N�c~�mb�S�:,f�"O���OA��JYeǃD�	)�"O�}��&Z�lS�	tc�>h٪5"O� 9$k:XH8s&ݒ!R��"O��$V��*�J�&ޖCL�"W"O��r����jRt��S�4"(RpƉ+&ʝ�6Ǽ=g44Psa�"f�>�ɻ`�.ejD�.M'��5͝�`b��#[�tm2�{��@�S��KcEZ_܌H�dN'N
�)ի;6R����m���bSȺ#���(�:������7�&��t��_��D:�ϧJ����O��6�S�R�h���A���\U��e��Bh�P~2E	�`�|3fa�)���0?)0�$f� ����g��ѕF�"�d�\H�z&J�[�|hP�%l��u�N�a���ŏ�ü�1#R���g-�$I��Z���x����s����D�A#�� &�؅ S�����/=r#��[ E�1OKk�Y��F�!�N�N[p��2$�?�y�HTL !����><2�!RgT ��O�#�j	&@=����ǆ��MUH�!|JDr�l�2}}�ܐ�iѐ�rЫC�
�7�<�'�I��%�p���<˴8B�#�?���E��3� \��
���`��]0*�{sIA�k� da�M�BY88�k�� �k�(HyQA�73���5fՁNu���,ĕQ�Ʃabg.[oN-�$�LJ����e��o�2@�Ӯ�z^���Â�]������C�9�r�XA���,<(��%k�j�&d��uB��b�c�IC�R,��I�%Ӻ d`�Q��'2�<zQ�8����*	)|�Ԅq�JגtQ���al�����'�M0�n�eX(ª�� �I�}�ԌY�
֑r]���1<O�)��3K.|3�E� m���+p��"lS S�lB���:H�*��ɐs���J��j|�!�&�{�vmZwi˩��Պ���Aa���gΗ�w���>�U)[�6B�X�.G5��@�J�ޟ�ssd�7?�h�9J\�b�Ei�5E�D�Sn4��H�JF�Y���CS�$0f	Y"l�H�lIɵƅ�7ք�Y�'�ָR�FF�� !��hI.a(����M��M�%a�%_��B�'WQ���MY$r�EP��D&)aD|�`n��K�l9B�'�@��$%�N@ڲEL��y(��9$�������&U`b\�tކP�ޔ[�ʜ?MdZM<�S9��|�F	H1�@!F=a�Iٺd�Z�D|�/�).�4��!�$H>!���݈���(6�h���I����"O���2f,}a�K�&1:��3O�){�bQ��Jt:��  =�>�P�CVA0d�s��_
=��(`�,ż(���O��[ 匩y�X"c<M�D�T[|yr�L=v�j �BŒ��S e�({�T:K>������$�>e���S��ϚOb$��ɦ?i:M����?t��{P��=(z�����o���+��ܾ�$��bךi�����>E�$�M�<�H�0O� V�J��F���O
��cㄚ>{���% ޴��O��)�gؔP:q�I�=�F�hI� ���/q|����'��"�HQ�(���K�9��I��K-%��8թ"}B�Ӹk2Py���q�­9&@��8,p���	]&.0�O.���dײY�P1��U/�n3��'N~5k1Ŏ�T-�':8$�L�>YV��O�DCX0'{�!!���N�B��N���=��Ĝ8��x�t�Q�g�N���흹���0"�O0,���U/h���O��}�`LX�@d;�E� ��,�l��@���A2i$�"}�� G���M��
�z,0i���Cr�d9C�LH���y)��	1��0��T'�<�Ԍ�ld{�IXu�B!AH��F�t�M-a/(%K�ҙK�]��e��d���Z�'�,��������-��\����_#b���	�xײ�1��Dj��ֺ����m'ɧugG>�*�c�ŵr���c	S#��=!7,Ν3�>-zF$g�2Ta�I\>Ȉ��O�u�x��[��0B�?XIqOQ>e�KÉy��t#��Pfī�5�x���2��h��=�0��/@y4}�᭐�=�ݩ"OvX��ԥ*�����f�3���Qh�5K[DU�����O��h oЅ��k��Y�7��R��'��,��A<zp8�ԉ#f���ЅȽBnu�ȓC@(�+��6E�<��ԲO�F�D|bHy@
aʶ�	�G&�]8E��,�4�)vJ�*E�!�ԇ)i����07�(1:CH'p��A�Hx�C��Rc��S�r �0��pn04A�^�X��?j�ف�fyi�,��J" ��}�'
�yHŴ.�܆�ID�*�s��ߪ,u
5�D%�!���dؑ"��!�O��P�e˂��X�X0Zg��	d�8=M>IWB	����rD6	PUM�S��$@VEQ�z��E{�ܐHJe�`�x�'`�^��?avj�k��V_.��;��5�	���#|槀 ��I�I��.�(n֚/:|�;��'��E�r��G�l��O?mҳA�![�xX��㝂U�V��f��<�5��'�O� ���'��ï�/_���U�(�_�lq`b�x���|�dɦOb�1�/��z5N�8�LNY�D�W�'�P�'�V �^$!��#g���'���{�C �r�I�N ���ܼ� <���5n��p��	�6u����W_e�p�B7b�~L��Y�t܄
@��w&�㞌(Т7�g~bΝ�-�dTٗkZO��Ⱥ���~2�J�]�>|�=E�T˃�:E�X�$�)"8��" �8T�cd)�O	��eԻ7�jU��C�#m�H��AQ��	��T�S�O��i�0*��Wg�a����'�pq� ��فA��*eFȫO��sc�<W�az���}���Bd�%�����S��p?��)��g(F���؊2�9����(E�g ����'mL�lqO�>wc�;ո�r�
޺�����-�s0��!;�'a�`8��	G���l�ǆ;/˂��'2r�� ��v_�y�Zr|�US�.Ep��(�%V��~�O�r#��=%>�P�%C�~��Sg�;Ā�XT��4'~��y��O�>t!��^�#�
9��) �A�q��	��DH!QN�(q͂��?�7��x��<2�ԏ�.��?U
W�U7c�Xm���Ův���ʁ�<�O��$�@�J�
�H�^	&���T�{48��f+���u���_�B��a�C��k����OdI"������Dύ ���Q��'���a�V�qZ�1�2I���H�� ��q�T�X�)��-�\܎q[���WX���w��	��äX�M�^�FI:�hh�}�����z�� 9��V�y�&_�?㬭(�K�N�\TХ�ՁIC���f�:$���g�V�m�Z�B"�W�{p}"��On��+����:��,�>^�\��RܧZ<>\��k���P���
�J���'2����b�Ny��)|鬁@�]=�Zƈ�P@��7.Z	���� P^T��>bَ,0u��_
2QH&-�Cx�X`Vm� &J���ԏ�}���!�2A�Z���H�"��ɚ f�A@�dЪ]���O�B�j�J��7�mrG^��ў�˳�A�ΘAeM��Ա�� �8qpa����P"a̻M+�9h��Q��zC�}���%�;K�� lA�2���H�|Vl��$�Y�r�������e�I1��"�� �%�션殘���	a�C"D�l�F'Z�L��z�Y#⎡R�db�L���]�P�=�Y:X!A2�?�j] !�q�>q�cL[����! %?C$SG��A����U�t�����B��!��!G��Z�G�$}��(� ��֠<V"���:s�|�AB��5uF)@��3#�a~��ِiXڅ�@ՋVk���K)(޹��D-`P���F�R�*5�F'�"�W�fDD}rj�.PV��qd�i�&]+ �� �& K�!�D5!򄝩3�yi�F7L4p�A��� ?�	7��q��铻4�&	[��M�XN\@��`��D�tB䉻ge�Q���<*�����
�,B�	�-u )Hu�ο ���	��ȕ$+�B�	�V��񋐤^%;Zl�z�H `I�B�	�@K����g�XH� ؽ|��C�ɇ5"�("���9[� T)�(��C�I6�\��m�6r:�a�+��C��"�!Y3�\]��B�6I�nC�	��i��nR�{lQq���
[ B�7��DR6��3yx��Q�/�4C�I)e�z�+�,D/�x�v�Ѧw��C�=��ٱp�,�R�+a��eA�B�I=_���㠎��M'�U8����zzB�I�P��Y�Z�hE����H�"*�C�	mݾD2��S�t<(�@���-QjC䉥^bA���Y����U�hB��/�ʰXa�/O��bB%��]�^C�	�3OPXw�3+��q��%qx���^�f�J�j�5`����1�.BS!�D�:g%�� �A/!YSde^�NI!�d�27ZXC�CR�}��iB�DK K)!�J�\�Gɋ�}�$|�BbO�/!�� ՘UnK�9�T$P(��&I�""O����m�'���G�H�1�"��"OJ-�s�P�X��ӱ=��%�s"O�� ��`ؽ�s%[�+^"O�%���#w���fU8$	����"O���r	\�cY�LQ���3�f$p�"O�Eqt�I�>@��̏�4�$�a3"O̕��&���p=��x��e!�"O�b�!�.�(�x	,�ନ�"OH���N�F��X�O
(?�4I�"O.!�����<�����Δ;(~���"O�HP������q�l@$)B,��"On��a��J�h�{EL�5xUԜ`�"Op1�d ��Z>ڹr��	��<:�"O�2��'�� F(!?��*�"O2�s�CF~�-	��ǜ�t���"O� �0oƓج J�dӐ�|5�"O�m��kY�.�e�����5"Of��tG�*(O��7I۠j��}*�"O�	q1*R�#�D@"�bK�-�L]a�"O�p��+O�R��42��>�8��7"O���#↓���a�%�+B�8�a"O��yG�k�$E��䓥7���j"O�I���Ÿ�B�����A��"O���B��A�I��udR-p"O \��Z	*N��e�$7p��p"O���'H����ViN:ws�)I�"O���M96 @Uq�bGiM���"O&�K�"DqIU`Y  Wd���g�w�<��`E�w��ݪ��	9� <X�OAV�@�ه +���8�B��p
����O�t�Ч"Opqr䊌�[vm�#�7���b��W&E��L&����5�g~��*<��)�aj�7�<������x�gK�'�v4�e�p$Z�1���jq�@HB��KUޙW�'��1(e�S-<Q�HQA�VY|�;�=U����U_v�+��'�0�5�l�@(��J ��'A>�#Gf�X�a��:.8�O>B��<" �[�Ӿpf�#}��G���*]�W���i��a�<��=C�F��E�Ҵh�X|)Ќ��>���c�h
^��E ʼx�~&��Q�A�\p.�fMM�B�""�*��8��Ҝ�ps�^�XN�#��R"vv ѹ1��0��ؕ$@}؞Dʂ�ȡ�V���fR2�@�-O6@jQ0>P� �%��7��6mG	9q\ j�Lߔ%��X�H;N!��9�vMq�i��)`�,�Ф�g�>�Å.|6�)�OQ�x�����IVm�O��.4Y�#���wt!�
8�rc��9�J]@��+W��@#�-3 ���I%�8�:���|Bk��N~Ԭك�¤`�LD!�ٻ�Px�j�&f� y��=(�$��kY�t1�a�2�����3Oa{ҋP>=)��do2X{JIsP�
�p<a���(�t�U-�P,����>d�:"l#qbEC`��c�FB�	2R��b�'��P�8��ǥ��kg �'�4e�%o�" ��`f�Vc�O�<�r��@Z��uH�13H�]��'�l����6���eoH�fpB�k��AXi*�`�����x���(v�B��#$�4#���/ :��x��!	b�9�,B%V,]�䦑�psz� FAX؟P@�c]�x⢨[%LՕ$��X� H)D�0��,Q%��d{DAV0K5ƴ��� D��S+�N$Ν�p��N��@��?D�ԙ1�ʧw�x6���׮��D)D���ւ8�"���b"5{�'D�Tc�-P��� `h�.<]	�#D�<�ԉ�`W���F�L�O��8��>D�<r1͕�3����J�O�p�� �?D�|�B��|<�/�Z���F�6D�� ��ӕc/tNeҲ�C�XhA�"O|tvNX� "�ٗ"�<J����"OґQ
�_zҸB��ќB1��B�"Opy�,|Rj`���'g5��Ô"O>����H;*,+!�={-,#�"O���/ɯe�Yr���.ra�'"O �I��3Io�5[��2O����"O^�8ㆉ�*�`C��܌H,J(�g"O`Y�'�,��`ID���E/6���"ObҌ�$(�l�*�+��-�I!f"O� ���̨5$������_[���"O���Z�X' :����G�6�p�c��
�!�eBR�R	tk4-�'<�>�ɋ�|��F�X�в (�vp�B�I o!��RD�AZ�%���'LD@�b��򕠊-��A"MS� %�$���vE��V]+���:;��D�OZtl4K%m���xrc�8o�:��W�ǧC��h(�߳/�&��c��y�ph*��'md��fC9=	�\��'S[�T�i�O��i�G�>�����ϡ24p�8�� p�m��
m�T�;7�����������@��y��%�v����7�#ʮ��P0ҏ�*|аI1���d<��I?Q��"O"[�lP�%2Oڌ����G���AGOC�T�ظ���',��(�F�);0�ȳ��:�ųC/Q�v ��=~S���A�=>�Uь?6��G|©ȶVF�8B@���@䁸w����O�xS�� R�1���}���`)ɵP��%��ea*}��P�s��i\�YV�% �g` ԋ^82P�Y���6OҰ���_�̹�r�L 3�Y�&���	<0��o-�X ;��Z�|g�*�gƑ����,
t�<�-��Q�  b�-���B��E2b��*EL@!%��] ��.2�R4�����`B�^b|�`�'O�}2	�;X���+�!Lt���u0�V�*Dl �����y���b�/,p>�b��*�ชW��!+����RG�(G Q�l���Y�"t��"�L�K�@X�T@<�:딍2�M�.��<��K�N�e����l�~u0��>*L�c���<n
�DѶ�ׇ��?!S�[��X��QK�������WX}�jX�����|��Ʌ4>ͮ��� �n�C�ʊ�Cf!��)~�=	�E c�ҭʳ	�o�'�֥ړIQ^X�4����sm��@`�!lu�	,D��a����ybH��A�4B�}�vg(D����6S��u
�n�-B�`��'�Oz���,=|Xu�������s�~X�
�'$Jm�M�;BD�F
ߠ*AQ��D�l���1� �S�u�M�G���?�~ea��&�$���U/�@욘'u��-֌C�Hъ��.jFda�'�b�6j��?ctU�O�>�(WF��*pd��)G64w���H.�=r�I.��h�|0v,M�~���uhvQU�>9M>;��̒`�,Oȡ�a�TT.At��4y��Za�\�B�qE�Rt��,ʧ[.��#�C�U�|���A=����J�piEL!����	���h�w�KW�"����O���
4y�Ta-O�1[bg(>���J�����y��|x�*bL~u��ܕQ��{�D����mIu
�����܏X�.hQ�d48�*t����z�,l<��>E�D�	[o�U)���>��s��!��'~��j�gE=��F��@E�@"�P&�G�	�>���^���	��U�� Ƽkax���)w|r��!�Z�xS"p�WK�-,_������'ZQ>����K2P��3ը��l��5�gAcA��^�#�O4�v#�M�\��A�8��� �'5*����*\��'��n�%r �T%��]<h��GQ�.��)�d R6�J����K .�X�
Լ�M��l��5[�|X��P�1��b�@�ky�!YCG��=E���*-R,�	K�
���J��
�O~�z��QVX��}j�dܒ6�����ma��(Es�<iq��^w��:b��*tI
�IqᛇVn9�U��h�S��?�E,~5�$���#"��GF�Z������	J�䘐4��p ���E�C��"O�y���tR)"���]nP�3�5�M���b�'KZD�� ��,�P�1#�;�2x�ȓ+�>x��뉼L AĬ��<�ɧ	�����R@��S�O�<���
�8a��Eڮk0ެ�"O <2��!�f�  ��Q.2Dy!S�,���SV��0��� bdI�*qgNThrC�0W�^@#3�'�T\s�G�!�v��ũZ)z� e��C=�2���WKH<i� �r2V����޳c/z�I�R^�'{P$�DI��P& ��~f���*��٭�u��X�<���ɤim��ś�,��ԟD��F3~S����>E�4�k�Z�Ce����m`ݎIj!�$Gl� %%ۈЀ��B�*5A�	�n%>hS�#�S�ayR�
d��U��)w���HШΎ��>A�N��a����ILԼ3l[�6���1$�H�C≌DS�l����.&颤��(�"9�\#>������؍��N�S�|�4n�� ���!�A ��yBX�^�37��<�p��~�b�xU���=E���j��l����)�������y�N�X(d��L�2�|�)'a@�y�"�"n/:�37��{N��j�2�y�,ܝE*���d���
O&�8eJ'�yBᓊ?)�!��o����J\�y��&v�neKT�
w('�(�~bkۢ$T�=E�$OB�&��a�r�;����슒�y�o��8.~]H��vU�وE�M ���*w蠤�1�0<O@�B�f�2w��IK�`��PS`�'��Dc�,wh�E����'Nh�
&*UM�J,���tH<q��D&\-b��S�S60~8��`�@?a1��Ƹ��'�i1I։d���~Z@x�ʉvp�Y�E�ob�%�ȓ%���e2Cp|)7HI�N��!��+|\����F�r���ʔ(B�!-�O���B	��=J5�cƃ#�Zas�'�^u1O�?,�`�G%ï�ǽ%�zK�2�t�W�'������R�N��	�oJ���!�5��Q�'��Ţ�=�'���zQ����1�?���ónx�a�Ė
~h�� ]=;t��2��0nOhC�	�C��X�s�U!5(<h F�H+	Cb�$�8�B%2CB�a���dV=@��h��K ��OC�-Z"ng��!� W2MZ��Y�"O #��\�5�`����#?��xi%�'����K�Y����JNT��ӬZ(r��(.}�?L�����&�,t��A��@��|"��9Z��Q�5O��ya��1� ������C@6Z��!�	�Q	&��`�Y8 `��*h��w.\��!�ga�agў�A�
��kN��K��@�Px#`YP��������H�^��rG�V�R��QX	�'b0��Pa����G��|�s��)�i<}B@���w`:��������|� ��<iHT���B<BC4���$�y'5��$"�oz���mա�y"O��H/���Ǟ��R�̟F�Y���<��	�O�
9q�~8k����X���'W�q�\��f$��#�tY��͆|�F�å�PlG�I2mi&̻�j�/G��x��նEL�!)�(")Eˇ��0?��cFO��5��M@�^(��з囖Y� Գ���
�B� ��4�q� H�����"'3�>���� ������rL�r/�)���Qc�޽�y�%P�r�ި��&��ޔ�2����dե4�p���{���3\���k�L	�L���_�9�!�ӳ=g�HH&��i�|]ab�T�!�qc.Ԩ'M�*k�`��"^�|�!��ԍ�|��6�ZOK�с��ǡG�!�d�$ȶ��&߽E	P�P�խ}z!�H�	]&�X'��^���lߣ?�!���}b��Ko�jeE�<�!�҇	���3�	��TUJ#�m�!�A'%^��1aW�?�x��M(X�!�$��x�(�!�h�b��,߱4S!���1M�ȼ��A���tQ!���]�!���ZF��+��X5��J�\�T�!��P7�iY0 �8����Ue��Q�!�W9����]�(&����o�!���-X	�Qg�2!�(�3"�0�!�ډd�x��5�+�~���Y�'^!�Dλ{�:���3u�^U����i!�D�=Xh-bD_:��e�MJ !�� ����_�	NLё#OD�7Z�3�"O���ϔ�T?~ѩ�/�#I��2�"O`D`�E�-%�\���O>W��re"Ohٛ%#��X�8�^:~�2��Q"O�9��&m�A�f�
���W"O�`;�iH�{��Xp*��Ti�Ia"O��H祚�?���yƩ�20��˱"O�����P_�u�Q�*:�nE�"OZisoת<5I8�F�%��B"O*� ��}V��`��6޺�0��'Rp$��·w>�#�	+&�h!S��A<a0(�J	�'{D]�%lK�V������n0�"�'_�8�F��(:4���ٜ���'M�-h��ظ)�lI��޸w�
�'�*�*4An,0gI��.P�'��8!�)S�B����S�)|���'+j��`ǫR�u���RϨ���'������13t��%+ɤ!�(DX	�
�Q��b��@6 ���W╂Fw�L�g�A�fh`'�H�w�!��e�j��DJ���c�7CXv�B�ff����o���X�-�q#V ��Y��� ��>gQ�KP�����C��A��>E��ƍ	�.`�m�$,��p��J�'�y"�B�n�DI��.��ӽ<~����	n������D����×-a�|��=�g�Ӻ���- �=X��M|�h1�$�fH<!��}!�E�D!0+�E��F�!�d�1-P�BG�7\�j�d�!�Dֈ,P�uA��сm��1P����-!�D�&I"@��mݏM��1�%=��K��䨫���[���sB*�y2��L.,�g�ɳT�4 ��	���y��i��lҵ���8Nf8�`�,�yRW�N�xI#���1�)�!ׁ�y�,(� ����_��=�'�yg�:.��A��?�H�Nϔ�y��O���0���W�l�bAg��yr
�S=>p�� ��@R��i��2�yR��)F9�-��I
5�������y�1B�X���	�U�h��7��+�y2L�hϊ��0�^�Q64e�g�C2�y�ȏ(��ዖ�R�X&+	��y�B�7�j}⇢�}���Vc�,�y"hI� :8�FA���ЋvE7�y"��}8��A����>�=�ՠ�$�yRգ3�t�6.��j!@Q���T�y�N��]v@M#��יYj��Ya�Y��y��(6�ba��&Iz\��7퓺�y2ė�n�H9��)O+7��1 �%	��y򉜼h/��ū�̪Mb��,�ybE�0:��㤪��n�.�����y�D�63�x5K'k2e�BI��D��ybA�( o+L��~4{PiЃYz��ȓ!�>�J��0�2A��I� [v:��ȓj��TGM�}:!�G#_bwFņ�,v�Y�眽301����;[͖h��-X,P5k
EWT]�K�.uX���\a4���.I�rR�i�kW?H�\8�ȓ�@�%.a�8�%mN:<NQ�ȓ0�
�M�����(�
6J�!��&��Z���*��<��)1l�$Մȓ�	3'G#�]1���$g�t��f��ݰnB�/��Ɇ��J�����TLF�H���(XL,AƮK?Kn%�ȓ�@%��J� ���p��X�}�Թ��hC*̰4�6�*����LҤ��S�? f�&'���n�a"S�+�x(��"O��j�F�U.�
P���QD"OL�&�`:ly�I 4�Xa+7"O�kjDA�9K����!��"O҄{%��,s�`lБ���V%B_�<�"o�����#W
P�:�	C�PZ�<ypL�5A�����BQRe���Y�<���Q�2H�g�Ǘjl�D�-��<���R���X��Pz�ҭhuƒ{�<q��ǿH��ijE���h%,R��H|�<�'+Y,H�5&�w�%��,Ix�<Q����g"(�L��-�SK�<A�)�Hn,�
d��r̊բ�p�<Y�b�<�@���^�����Ϟn�<	w�����c�hM�!P�k�<�T-Rs�5�U�-��XCDRe�<1�ˑ�p���+?������a�<���Y����4�ɣu�{`B�]�<1��z+�,@���<=x���ZN�<6$�J��*F�A�� ��F+OG�<a� �,#���4�x*X���k}�<�1!ϨJ���NP�G\��3ׂRB�<1g�\t���@ꈾl� ��wc@�<����+I�TE��$�>�F��HC�<!Q� �N��aM�O Ȁ�cJ�}�<�E�~x}�R�sg�u2�E�D�<ae�V0&h&a�G��\���4'�K�<��̲A�PS0�]�Kk� 2��YQ�<���C�Qp�@2E�e�G�W�<!�D:o3���͉:pY��m�<)��_8�����փ\�ČKt��P�<A�Ɓ���N��id\x{��_J�<��'Ty*Bd�����j&�%��o�@�<	�!�":���u �Q�~�Z��MF�<�CΊ7�a��͎c�-!�
_G�<�'����L|!u���N<���dH�<�"�1K|	q���L`HBƮXi�<7�̐r�d`��/���a�g�b�<Qd	�y�``�NC(I�.<r!�i�<��"3J�R�3@�٠�b��@�<aB��T󬑪�ʞBq���P�<�JX#pX��X���[ڂ�i6�[P�<Ʌޜ���fO�p�@	��̚I�<15�'U�J)2Ql�99��|ytoZ�<ٶcE�+":(`�#H8 �f�⤦PS�<�B�_�~X�X�~�Z��t�<����"9 eQ��5cm�<����p�<a� G*S8����Ny�s���y�y���QU��Jt#+��yB"˸�@ E	�0<���� �"�y��3I�B���c @p�!� �y"��"6w�}�����ڠ� ΀��y¥9�${P��)	Hʵҷ ���y"��>�. ��F	�( JB.V��yrI#��l�p/֌~�`����y���$:z%��!;�pAf�2�yB�?�Z4��.�>� ����yBL�JCn0 �`��
H���7"�y���,L�9t�<	��i�J���y"Ҏ{��0w&��0ݢ���P�y�Z�~Ҭ9��9\�r K��ϲ�y�L���^(���<OO�H����y�Y�M;,�CW��-8|�ťH�y�� v4B�����_�rIjrN�%�y
�  $8T�̎������I-
��"O��J �-��0�OV�\HH�"O�����P85����aD�6�&(�U"O��X��� =��A��ͪgyt�2�"O��������P�ȗBf����"O���Q��05�^��0�>k��Z�"O��jR�S1#.dE2G�D�9w���a"OV�(�� Eݺ)Õ�W.w�}Z�"Od��!l��y�-Qq��<nn���"O�����LE�}�fYA`"O��vf�X��|�����vʜ]�C"O�$��^'���'�]�Uʲ��e"O��G59��`M$t�\]�A"O�9�bM33��x��O�5'��|`�"O�m���ǎ}�1IN���$��"O��(��P��d1aC^7t��ȣ�"Or y� �/K���{ŢWe^��"O��
7H����@�"�l\$���"O��x�d^L���8�N�H�P�17"OF=���%����3��*p�NpJe"Oxc�E]�����jE�i�*9�"O�,3ĄO>Zz4<���$*��E"O�D�sG�)z_*�Q��
h[ "O�"�g�!^5l\�Fƥ��ѳ"O��[�f�P�j+7�+1h,u�*O0�g�nm�t�s(�Z�Pi��'o.%���;T�9ʕ�Nj0�	�'�x�I5 �rK��'��H"ੰ�'CT���A�6� ��?K�0���'���ˣW�0C���Ga�\H�'=��h@�64�x�aܥ<&x���'`� ����'ymVՑ��2-d9�
�'x�p���E���꙱+�l�P
�'|l�9��x�p����#.�2
�'ն��@:�<E���%�|i	�'��r�Jȕ<[zU�C���.Q��'2|!��aZ7U	��P�N�7,�U�
�'�6L�lPD��'��-?���	�'>J����Ʊ`d)��E$:<"E�	�'���TdH�*��	�! ;1���
�'VT�7B�'�2IҀ���'<d
�'�:�PЇ��(�}� AQ�"J���	�'���R�ٙp�PAB��G�lZl)�'T.�� @ _��h{1c�4����'-����&�!#C���,`~���'?����%;��kA��;u�*$��)��Š|��S'@�8r�f5�ȓ�ą3F�	7���[v�Ώ$C�݆ȓY���E�*LB����ď�b��ȓ?;�hԨ)8i��:�G����ȓ<��|���(�p� m@Dr���d4<�GmЇrPm:�o[E>�ԅ�*�4����N �[����)�^���cS��ˮKdީ��$�
q��a�"�� O�$a�虃�R�L�|t��z��bO�H���ɰF,FB"1�ȓ:��(햨D1��!��/`��9����o\�x-��S��5nTF!�ȓ~�^!�4�1@�NӴ�H):��ȓPB�D�n�H�Z���4
�nL��@d ���I�N
���%΁�g�^�ȓ;[��᢮��X�JG�{�N��_� uiрG�@)���3���az.��ȓ0(>l���ًW� �k&�$	 ���S�? �X�5%�_%R�1�l¦XV8��2"O�	��	7>�Pp�IBnAq2"OT�Ku��Ue1�Ɏ�c"R��"O�yS��2|K�-���ʀ8:�0�"O`��� �`XP�օɗ{'pѺ�"OʭYiۈ�����#�Y�s"O���E�ƃJ%Y�#ʊy�X��"OJ��LÁj�. �d@�Y8l�v"Oxx��dv| �&�M`��;g"O��q#M��EHs�^� 뢵Q�"O���6H�w����叙h�p���"O�����0C��\��Շl�L��"O��2B��l����c��|��"Oh��P<r0��e��-
7"O�8�Bb�4B���aB6d��y��"O�����U?.$k��/?�H�k�"O~M;#n=6��	 ��&~��哕"O(!�$�Q:�Z� G�x��i2"O<<{G�K�=o:�Bq�ޱY�A0�"O�����U>���� %`E$�@�"O����ˣU����]< ?�u*"O^!�$M�2��	V	

4.�"O��f`���	��
�9��4@�"O�=r��΀�H]궤ҧH�j�:�"O�e1`�+��r"�
/{�E��"O�i	�`�&q:�E�C!�H5��"O��;C,�9��ar]�#���"O�uVOS�X�DDK�*a5Ĥ��"O��
�P��[gO�
c)
YSv"O,������R�$h�/�B"@��"OH����F�PY2I��m�0��{!"O>���aA吁L� JP"B"O��J�ϛ�{Y m+� Vi��Q	�"O}����i�U�X�X�"O�E#*����9�fmX�-F"O�h��)�0k�r���4]ɬ4��"O�����y���,�'�E"4"O:4�ߔ&8�3A�ޟfW"O4�'�E�K��2b�����!�D[)c �  �d�a� G�Q��R5�fǦ��"OH,�b�O3�D�@e�D-�`�2�>	�tD}���˦}5�m3a�ѥX :]���?q%�̆#���X�O�3�9j�b}�<�ǨĲ�r(j�I�?��0QaGx�'i����i���S���-�̘�f��<]򄙳&Vg�����΀5� b���Bb�9YS���J>a|r�|rI�=>lʱ��/u��Y1l�=�xR�'`��4O�Q�潫�@��@0� �����ȟ�mS�^�.��ć�4���O�)��ʆ�$Ԕѻf�W�>Hj�QpE�ܟ���2���`�� -�R�*Fc��GČ%����ē�(��Y�M�='�|��J&NH�f"O�i��e_24 �"Q���`k�04��D=}�1O��?�cJ�;IҰt��L=�<h�ڟ4���+�|h��g� �r�r�JU<��l���1��'�*ub��B/(����d
��C-�,�˓�(Oh�C&bsD0����x�|!T�$d !,O���yʟ,�'��a�EoD)2�
��L�(�dߓ�'(�P��P�8�0OĆSH]���'"<O����O� ��
�HP��*0��'��w�i�V��'`��>O����g?٥�C�:!H )�.��"�m��U�<�"��й�񨞂p���r���P}��)ҧN��[�E�lde��̇+[�L)��#P,�U�6�b����c�@%�4����%�qG�<��,�����i�`B�I�N8�)8�\�G������;8B�IOa6=�B-֧D![��Lx���=Y�{��x�-�C��xp��T�J�������M3�'O����Ӷ{eT��cM�
�4��'�T3P� :�B�/Ɲz��'�zuH �E(f� �;�0`�'sʉE�$4��:7 �,4ڽ��'�^�C�(�"DbT��l̲L�^,��'΄)zäT-m"h4�%�!?P`��'6��VA�<b,~D���"m��a�'�1[�*��GN�a�X��H�'0(�����4h���H�' Q�
�'�h%�r�]�,cl����rɒ։�d�<i����q�P����9O!RLh��Fb�<�F*�';�^	8` +�N1�E.�c�<��f���(c�.'B�4�ӣ��\�<�`�A=��HS/��Yx���&V\�<�1 T!�����jǈ~�lx�7`MN�<���=t�d���|/�ɂ���c�<�qȋ�m`�5S��&w�v*d(x�<�Ch ��R-���$n����b��x�<��B�:�*��,נ*��q��w�<QO�9"g�<����>�(g'Hu�<9�'�[�D�	S��cd]��IOq�<ٰ��4�kU�Q.�ʤ�w�<����,z �&&�i"f���*�v�<A�EӦ>�Bv!�Y�6�S��v�<�d�G�i֬�Z�J,ql�qK�[�<��m��^�@q+.yܢE9��V�<�GcO�"�~���4d�Й[�QR�<I��ϵ(�d\0���2r[d\���y�<����Z�j�
P0L-��"wDq�<𦑒
ʁb�FG�K1�Q���c�<i�L����	�(|���9w�S�<���-~�2`��Jp�4��E�<���&1�<R��$5z��B!�D�<���2Tqy%�^H�����j~�<� ��'�ε$�b�Gs~���"Oz-���L�]�"�Z�;v�3b"O�8`����0�"L{�bخqpP��"O������TKI2f4XZ�"O�hC�M�3 ��b�ɀ�c��&�'��P���Iٟ��џ��	���=M,ʓ�8[,C� �I��I���I����ǟ�I��T�	۟\�	�ǾI�d�Y`�<��"�� ���������	ޟ����h��������.<xs*�&�A8�a�7u�����I��������I��������I�0D�t8�J��S����P��`�	����ٟ���џP�������ߟ0�ɋJ���4���9Z�ͪ3�:��	ȟ�	����џ��	����۟P�I�Q*@p�UnR'�Fi���N�;����ß �	�$��۟��؟��	ܟ�	���=�r��(T0�e+���J�j,��ß��I����	���	����Iݟ<��)�h�h��K\|�0��B�������͟��Iɟ,������П���"o�"4J��"������!^4u��������l��ȟ\��ӟ�I˟��	/�qA�õrD4:�ҳ]M�)�Iٟ$��ԟ�����X������̟���!{�m�hT�|$��0�K;n����Ɵ�	���	<�Iӟ��	͟����;�v�
�m#�s��(�d����������\�	������4�?��b�V!����VP��� 2Z��#^�\��Cy���O��m�Cv���&��X�\ P��L�n�1Dn<}�i���'���/�9r잴Q�g�4 R}���Pi��7-�O4�R� ̪O����'���xR-�V��^X.��j����5@�Z����<I���7ڧqn����g��J����N��9r$Y�&�i��#�y"�����* {U	��3����&�j��
��M��'3�)�I,r�l]C7O|}����+OH*�ؐK�;-�8��0O��r�X��l�KO*��|���a�� b���f��$�5N���ϓ��6�d����s�m)�		�&%!僕m"���`��-%��Dx�\�������̓����:���;u��^^1�+�/�	�5l4p7�-(�c>aAW��,	���I�/����ƚ���1gĖ�sW&�'s����"~�yL���C�o�4�#�.��Γ7p��N"��ᦹEx��E��Q���Ym�0��7d�<_�Lp���?9ܴ�?�"ċw����'��쩷n�$����fح�D����]�k_h|IY�zjў�`y����6|��x�BXfv��6J̎������C8�J��P4��JB�K�=��Բ�Hc�z�[���	�Mϓ�ħ���.��@*q.V�ML�9��]�6�"�[��:"��'�2����7W�z)�f�$Hy~�"�M ⼰4�O�h�ҒU)R�8�'(�'x�6�Y�l��B/.�*(;��H�K6>�� �<���iӎ"<Q.O��D~�
�D��
�0t��N�]2 �剽K�@��%��m��ǿRQ��;R蛻	�8dI�O?����)B_c ┣ǈ� t��P4�Qؔ�*�'��]�d�����8zq��(Z��c흁1砅a���Ҧ��c?}�i��'�)S0oH>mK`�z�+S�dv����?O���M�r�i���E,d̒�'v���to��ZT��$g<���M�U�1�����W5��rF�x���{y��'�$�R4�6.�L���l˝����'�'�
6���1O�'�|��Ȣy��F���S �i�Odʓ�?�4�y����O�X��O[V���f������k��Jn����������Ĳ��9$$�O��׮��D#(�qW@�n	�U���OR�d�O2�D�O�	��0E��]��zٴ<��Jp�C���#�"��!����(��<Y��?�����4�ʓ<���C�~E��Dy�`{G���7m�)p�dW��$�����!=FNqJ��gy�kVO���j�x��U`g,K���'�r\��G�ĨD
j��ֶ��vh��l[����+m�|��E��b>]mz޽r�ML�{�=S� Y �Ez�A«�?!�4�y"T��	����� M� 4��>O�Mj!I؂v 0Y I�1?n���1O�-�၊��\k�;���<ͧ�?��f�nS ��Elr�!Z�b���O��d�O�Y���IV9�y��'=��q2� G!?�<�P��¬sh�'��Y��ݴW���O*�1X��r/�&f"8���#� &����?Y%�W4P��� ��3������"��v����?b�����6.�(�R5���?�˓���O?�I�*o�d���� ��A�"��r��牫�M�`�u�z�^#<�ӗK6:@H#�;S�͋��BdF�	ڦ���4�?�%̘�n�l���?��4���2�@�,��� E�$-(@���ܤ��4�B˓��'V��	��\�G	S�%J���!?�ֺi�(:�y��)��L¤ʥѫ�H�S"
"<�'���iD�)�	����a�Dy*��o,��H�˰Er�8FE�\�ɑa[0��,��)��E{��O�{tx`��LQf�jL��KgRW�d�'�'��6͑�U��\�T\���R�,�R�L��
��Db�#<�,ON�Dp�����I�dy��-�,^��$��:UĹ�nI'��ON�)%e�J�li	������3�5� �="��Զ*��9[&
�ZfQ�2OL��O��d�Oh���OD�?�ڑN��O����N�Q��	F��y�'R�}����7O2���O��OT3QI\�v9x8wːo˔�@�f�l�'&x6��Ʀ��ӊW��` pNi��mڛC��:���>��%�W�V�?."�¶�+��LY2�hO>�į<Y��/��.�2!R���!Y���*3/��<IO>��io&u��yB�O^���t���A��/Ř�"˟����`y��'1��<O�d�)�,�*����+m�(p�A��' E����}��JW��\��66�2h��DE�2Qr��I�HRIf��7j,�'�2Q�b>�~���J����{s$�;J͞�a �g���H�(m���l�<y.O6��4�.�r0�,KlJi2(V�}��EnǟP�F+5A�����d`�P;[�r�� g0?&i"Q��:w��nD����Bi̓�?�*O^�}b�@S�`f2I������r�f�;mE�����'���I}��צ��q@i� {l�Dӱ�W�6�pi�	ڦ͓���O����'a�����S��y�N��\"*�w���YJ�ZŨ5�y��x�� �%ĦU�ў����v�ۻT�|���4N78�v���'��'��6�LU1O�Q6���czn��T�٘r}m��'/���d�OD7m{�p�'���R�@_�L`�Q-P��V0��'� ��F*Xq���/���⟜L��_
Fb���	d�ظ��N�JKu�{q��$�O2��O&�$�O��������4L��rs��a�n�K�\�Z����?���i�Œ�'fr�xӦ�O�9��If�.id�!i E^)8���
�:O�0n��Me�iOBLR�N��y��'�LASĈ�-|M��j�E��0`���( Ϯ,1d��W��'����Iџ�	˟ �ɭ�$`�pc�xo���q�C�:�N�'�z7M���O���?�9O8h����/b"����퀵(�Ձ���gy�)g�NM1��n�8q&>Q��?�C�Dս���1����j�6�,A���J�5����0a�*)�&�;J>9-Of	sB&�J�����W���1eŢ��D�O��dV+jtfo�jyr,{�fH��8�$qX���y�f���G�W�s��O1oM�i>�@�O��l���M[��i\�z%�83X�c~�1MV�C�j�@F���y"�'�d�JE�Q"}V�I3�W�l��5F�1�j�↨E<7�*���R�y��'���'���'�R�)٠N�� ���U�)M�9p�k�.|�I��O�����1��w�����M{L>i0�7$���jW&�5vfB]1đ
��]�0��4[v���O0�y�v�L�yb�' f�GF�9�.� С��Y�f��݊�p@�h vў���ay��'�l�!��T!L{ϖ0xQ���'��'g�7���r1O�ʧ``�{�	��yJ^Q �������O���?	�4�yҜ���O'Z�w�
�"]ˤ���D�"8�!�՜s��5���9��$���["`ѤkdV�O��f�D�Hۆ�AeE��v�BTI�O��$�O��d�O1�&�'"�F�	���ReU���H� Ӄ>,���'���'ɧ�\�0��4�2�E&��n����3~�u�i��6�/o0��:OD��ҙ� ��r���sW�$���hc ԝ,�6Pb󏁕b;H�Γ��$�O"���Ov���Or��|R� �.f��x����c^Њ��A��OV"M��'9��O��d�'"�i���1��4B@�Χou�\�f#@(�4n�M���'��i>���?���g�PZ��	Qj�2r�+\�\�Hb�PBh�%#��q�n��&!l|%��'^��'�<Dbq��I�a��H��ϤY�4�'hB�'�"X�x�4z�A��?y�MZ�c�cֲ(`j�c���d�>Y��ig�7�C�D�'N)�WBɁ���ʴ(�+z��O.�pk /k �횑�,��'pU��
���O�z�n
"�
�"rrEr̘�D�O6�$�OP���O��}
��\���1�-_�O욄��nõa�Hh�����v�݇�y��',�7"�4������q��B��brLE�m�����Rٴ(���M��E��p��'��C�t�"�[EËvlb�ڗ���
�͘gf��d�(e�w��� �'g�Oƨ�� �f�tis��>]��@�O��o��Ojpc����@�Q<΍`t��x.�-�P�F(��џ�l��<yL|���?�u/����4Y!���&%�榙#"t�hkl~B�M�DuH𐓈X*ў8 ul
>B`�Xp�Er�-�g'�ß�'<�C��M����<�C,
+7XqHW�G���a���I?��4�O,ʓ�?iٴ�?��\u[ذ��	�y�����E0m�p�蓅M�<��
j���@w_���'�$a�AR�Нdgdɹ��+/"�$�7$u����\y�T�"~JGb1Pf @fL�,\l��C�^k̓7�ք�����Ц�%�P�W��s���Z1 �����CdR�<)/O6�ߦ��	��1K1����Ƀ|��`+���#M����+
H\�@�?���(��Sn�A\2">If+Ըgu��y3f�AN��wgZ�<6�á ��h�`P	:�p��#f��`!>"  �"����6pp$�Vc�'���S�*�6�B�A�t	n�"cd�9'��%�%◷F2=�֣G*�I�aMTd^���g��YQ���c�#�|��䚡jZ�]0T�L���BT�|�:�B.�����(FܕA��Q=)_h��(��P����٦��I���	�?u+3�V8G���;b&��g���1�a��ē�?��0ц,����?�����#c�֑��Z9.a�4)�4�l������)-�����4?������S7��� ���G=~�%��)�+��� ��i9��'s&I �'�b�'��v|�F �>4�`����^P����_ɦE�����Mk���?������x��'��u��I�h'��H��=]B�$Bd����O����O ��~���?��DV=RH0��DF0}�P����R��F�'���'�����e<�d�O������Bl�z�*yXD��� `��@%�lӺ�d�O��$�72���O��iʜ=�Li �oB�� �a�͈�.�� �n��b�dl�&��@h<�b�,�RE��KN�6�lPbiHK�� ���:�xRr�^	E���#"8.M����^�Q
�z��]�$�q'K�EO��yd���M�e�� 2:e�d97�U�}RB�;w�P�~��@��8�,�a�v�H�����#��g*�6J0W��,	C�¹��dц��h�R��O@���dң�mR��P\(X�D f�:- ��'BrJ�M��'
2E��u�,I��΀B���iCF}����ǧ�8h�ʰ2#b߱*m	�̒Ʀ�R�1ʓ`��	XTA *U4��������C�#Ղ]��IC��G�����o�!�M�#�e�'�|Q���?��i��o۲�"���Ā���13h[�K��ҟ@�Iɟ�F�/�F�,@ڧ.N%�n��b T>�xR�zӮ@2U�E-_���R6ni�
5j2��o�]y���+N�7-�O��Į|"E��?���Ͽ!� �� ʓ�Mp�H�����?���1���
t�r�y�$·8��P�S޷wj�dA.����5�<p����a�De�Vd��>AS�,��-PvB+6��a�H�+:nH�RJ<�N @V5�COA�\ 6b�T���&$��NdӜ�oZ����J`�T�L8���7�	� �X���h��?Yϓ'�ؕb%P��8� N�<,(��ɯ�HO���Oξ .R1��"x�Ъc������Iȟ��I�PX9sD/^ޟ��͟������1�+\Rڠ� eN;Kf�;DJ �R��⃀��?������ы�L>чΒH���
��[��ވ1�� m�����Iз)���QΔ�}&�p����	�H|����Z0�E2iK���Y4�U�)�3�DS7�1�g�/:�}�0�Ǯ{Y!�]��p�W�8J":��pN@3&M�ɩ�HO�#�$12���@�B��G��0��H�]�n #���#V!��d�O~���O�����?q���?�Ѩ�"t��ܪ���n�DXւ��&W�I�w�M>]���J�RJx��!c�B�\Fy2��8i��)&"�&�.y���O�=K�Sx�+B�ҝ������ `DyB` J�4�p-�\��A�����r�Cԛ�D{ӊ���<����$�<Q@���n� `V� '�d��F�R�<�"=8�v����ToF�Q�R���t��lӮ˓}��,6�i���'K��j@�&h�.�9D�%30�sq�'d�M��'W���>Q'l��Bb�<��Q�H���mɟp�j����ɷhM�@Y�ьKd>�I�n;ʓb�RE襭�-\(r�X֫\xd��ó.8$V~p�A���$=r`A�L����Q
�#
�.��O@���'Y�@!�ԵL4)Y�@�"g��ʰ�`�H��ן��?E�$&L�QXR��0��?u��M��x��s��|A�2H���S�8�i��g�Oʓ �,\H��iq��'��Ӕ����ɒc(Xe�5d�9'yJѡ�A��v���I���A�p:�(�t���sj�9�S��^>u�@K2F�@�D��Jzr�+}��h�)��������I��a�q�g�[d�����	?�"�4����M#��i�����9d�,qL�4������l-1O��d8<OX����W}��2�hP�Sʨ�'��#=�Ӏ����	�v
�;M��p���8�X����?��S�����Kǖ�?����?���7�N�(�$`:�?R�g��Z��D#	���ⲹi���s�
{1�*!zV)�y�_�s@E�� ��D�����7 q�2��L��K��ܺU1h� %Sc�ӠBʊtY�4��$�#��E�|Hb�"^+]T� ����O`���O��EE�Oq��ܟ�q�����{��~����AG�gq��D���<1E��`����v͕�B��ɐ�HO\�)�OPʓM� ��qdCQ���
u�J�t�b!��7Bz��h��?1��?Aa��B���O�瓖,�PQ�Cl�½��S`�paU$t5�d�U�� 	q��hVaC>'���;��.s/2jRE0c~!�v�֪ b���� ����K�1��ݺb�ٚ/�Hp�N��(OХ��cZwd��p��پ9@Uj�S�Y^��h��,o�̟D�'����Z�#@P����/ʸ�*R��<	!�I�;`�z�ׄx�� k�� %�1O��l�$�'K$\��f�|�$�O�lJ�I$��B�* ��yrM�O���I5�4���O�擄�TTs��9�DDq��T �"�R ��-�wbI�2�H8�2�3ơ)s���x-�t�ľ"����1�V )F��[G�]N`4��oȎ]��`!t��B�2!X�Ƀ7 h�HN�Ƀc���qOȱ��m�!kΜd�&C�	2v��jf �4���#��̍Ny0C�ɍ�M;�l�^�QR� D5�.�AI#��F625iQ�i�"�'��ӱj���ɌV����BFYL̝7�����I��p���p-��q�	Ē`�������k"MA�TG��ȁ�Z�	.�>w�JA�d���:M���X�AĴ/Թ�ě�
 uC����}���:4��.UKm걋�I�z�'��,j���?AJ~�L~� ��q5F͸)�N�4��Q��!����O��D݄-�N�r��'cP���&ax�%7ғ;��0Z%d� 3�ȅ�VΙ�\�|Hs�i�B�'�	���Tt�']"�'��w$vX���d��+��X4NND�hP�ʍ'��@5l��ꕎ��--J��1O�e�r/��X<�pf�d�@(S�/�X)�G�U���(�)��"&q���b'T���tK�=�$;pڳ�Z���ϟ�X�4�?I& [��?�}�'&I[�T�#'햾\�L��fӋ��{"�|2C_�rڒ�saA@ZW�J�.��$�Ϧ��4���|�����Ĕ�~1`� I�f��D`%��v�d��@�,=�6�$�Ot�d�O\�;�?�����E�Acf��˄z�dɲ�b	6v(�0�'$��d@7-�h����F� 2'��x�7@��3g�J��= ����������?A��E�AYf�1�͇w�B1��Ar�<YP�١0k�thv�V�W}�M*�)Lt�(��O)1d���9�	ӟ҃(��~�^�"`�3Z�H��Ў��H�	�f�����']��aZ���*i��l���O��h�㑃��D�w�É]ux�4�'I��ҕ8A6���aܬ[\�tц�$G&�BR(�g/�@��4T�
���q�')�c�E.�'�f�B!ʓt�(�0g����Ţ�'U�)��
\��`e��MΣ�nP
�'�x6M)4]����N'2q���
�N1OXq�lIϦ����O�L�''�U�r�ԡ8>�ċ�LP�wj�u���'��"��>���T>�u�]�anY18��XE�:k���O��H��)�8\4�@qg��"X*8x��`=_1��'�\p����ɧ�Ox8T3V�N�jܬ�s�(p���[�'�<a���%,X�@ԆZ.,|��
c����=VHL�S�Œ&�p2�7D��(fC��d�.u���L*~� 1"D��J���q?�I##.D-^)� �#D�P����c����d�)X�@#"D�t���ޚy�^yK'�.��=�E)-D���Ǉ:R�=�F����)+D�h�����\��Yhh��0���h_<!��ψp��(�ę5W������e�!򄌚*d�S�"4D�T�!���5�!��/%;*MCE&�nxP��p�!��O�F� YK��D�)�p�k���Z�!��6�ʒk�=X��J�n�a!��P���HiB�(��u�'�?	�!��2~�PQ���P��������f�!���m����+�D���_<Y!�[��P�@ˇ�,:��- �!�5pbj5Yw��\	~����F�!���q:ŧ_�E�*cC��$8�!�_�u5��H�܉7�p	4��r�!��Ωs����jK1_����T!�{�!�䌋�>�Ãj

���h��E2�!򄃂 ��p�vk�@oN-��E�*]�!�sC�	�̙QZبq %A�m!�D@���9��:Bz�X�c��!�d�S�~���E'2�����f�!��QB���eU�'H-�Si���!��Y�?�Raӄm�6&�K��B�!��C�^���梗�����M(v�!���F�<� )�![W$yQ"+�3)�!�$ &����DQ� CP}`QC!�!��C�nճ��g����Ä�H!�ė�w�@Qr�U�ijz�Y�L-!�DS0[�ȳ��YH�x����^�@D!�DD$qFiއ:����1C!�:zצ�)o��2 =���)4!���4@�MrS�Ɋ�Yåm��Q��3��� j�LpW�٪UqX��e�<���K*x��ǆ�K�D]1!*Io�'��YP�cȔ��]H"�zJ�CK�i1�N��`�3�!aV�0� �6Snꕓ$&{3�|n*C������f0�5����v�0�G+ݬ7��>�|��l�43ޕ᳎	�6���<� B���Ӛ0�z5
��E� }�-1K�!�܇�kVGԚ\�ԑ�b�̅E��|�b��&�D�ˉ�D9hf�]Zp5��hctӄj I@�_�|Pt8y��'��iap�Q1�:�	��^'"��Q.�
��$:FiŃ"��t���Ĕ�1�,?)��͋E��͚Ԋ�	��E1�-VI�'���2cBr�&M�̈́���5x�
��G�>1���W	Q��h�Kٲ!���zp��z�|�q�[�V;�,V�'.�R �F<<P,��W����Erh��=q�@&��<��O�}&4Wo�T�(A�a��e��	>��F8RDҒ�3QT���%��]��a�+Umy�2M5�	ނ��ԭ����L�!V�1�'�Za� J�!e��hO��%4ڗKW
��Hp��2pw����#v�|j�'��T�r���B�%`�%�'#VH��G�l~�DY����{/T\S��D�O��ӥ��~�V��d��+UWT�Z%I���q�`�T<El@�bG�)�A��'L&H�aT��o����c ON��L�,:�	2DC�+˜�B&�'It7MWAijpm�H$��ó�dXFy�	��?4X�ӥؠ��0ՆQ�z��ϓҘ'��0C�� �E	J,�)$q�TFtkZ��A�'@�|��J��y�=*�m�n׎�r��c�9��'Z��jl�fǮ��	�dZc��}K�) �?B�LK�&1))�%ȰΔ+^{��V�?����'���a J�VP����i��8�'���Sr�'�:7�B�UԼ��ܴOcv�I�ϕ-w,��%L	sJD|@�,�z�H�p���P�2�L�'TO�=���o�xxr�N�{VI�'U�@�}�������
)|���M�/�7�ى;z�Gy�X*r�d�B�G�E�2����Ta�� ϓ�~�S���uI�Ks�@�� �����7��t�0/{PQ��;ea��;���Y+��HH�@�xT�e��$�<����W�$���#�䅲�N��jʨI�"�1�	�	�c!��	a#�
U<�S��U2K��QL�����M�"�|�.��2w��I^���O��D��<�K��d���D���`6M���0�{Q��H5T�����CQ��t ØWكPK�=m\.m3�*O�Ų���?]^�5�AK��~�n8��'97͛�F�hH��'�-c� �a����Dy�nI��h�3G�gH�YԊůjh�U���~�꧟�l��8Z��b�ܥAa�0��E��QM�h���U�o�Q�\��ߔ�nZ�6Xu;$�_�^`��˙ �2�p��j`�堟��O����5W�y+c�[.x�V (�,Q)�$H'5m��R΄�pf�T)?�u.��*`
i�� �Iz�Ey�n�C���?q�s��а�Q�c��(�&7K���<(���F2P�lQ�*Y�MxZ���œ2Y�l%��a+�ـ�E]�0(��~�dH�q�Af����wk�O\�D�$]��bR�Y?7�1*��1>UQ���.B.Up�ŋ�ժ`#h C�	A	m"��%�I>��Q��[�����M���1�g0�Jܲ���.H �Ґ����Q�G]�n�Zi��+� E�ؐ��*�	s��|��z*��y���$�
	�t-�=�`�Z�ÆI�'kp�2������J�;����O�\�#ǈ;n���)�Õ�W�9�G�E̓�B	m��s�%�tex���49N��ݥ|�b�%c.{rf �Ek�~�n��C%��6�#o�4���c��8{����'�H�.��s�PTG�S�6i���tk�	�=�tl0��<t	��(J���7j@*{�X] d�pȧOj�=%?qP��7Ɋ8b����}.4U	w�A�|ᕤ��Q����JC�0���M���h��L�Rl���Mԅ�ڢ<i����u�Lb�c̞J���DD���9��5�G<b����׸}�<X���K�V��'v�l�s!��s-�C��.~!2��e�=�~���9�J�np��*Ӝ�5����5����*]�g�����a'{���UI�.��z"�H�:��q�c�<�3�Ʉ�	��\�q7"0����gc �3a�܊���"Ğ��4i֙"B��GyB.�o�ʘ���c0)a ��|dB��rV�<�A)}����R��X��1o|`x �:W���#��� �X���ɫ.�aEA�g���eO�N<���H�1��`�Ox	F��O���f�K�\\�'�))U>�K�"O�ݫ�O5,�90p���G;H}�P�i��ৎUG�.����@��EȖ�-d���lُ!�����r�,�5Lӕ�yb`�Bj�kS�Gi6�Ͳ���s�<IQ�)��񇥏�z�&A��[�	ƥ��.U����}�V �� �z���P K��qr*A|�<�IƐ! PQ�둓ow�jD�d;
5��	�H��I Cp�@�e!P3�n��W�@�wĶC�	,P����ٴ���"S̙�o�t7MG"=�0<���O���=�Uj.�ab�c�R�E���l؞L8F�H�z@��'�l�x�Ć���{�%�N��$��'Z�� QLD"8ҘP����?і���}�_�%��ic�TQ�π �h C�m��K��/�V��"O^�[v��#��a�l
lk\�Yv�U�%'X�5�?}��"�g}��'s2@I����Z�\��R����(Oh8��3�@H����|\��VV�����k/2ɪ�㗤aM��+fMk���'�p�]y�AF5_?$i�N+��qnZ.�BU��4yw��	d�~�`'D%!\A�sOI� ��C��'O��ڄ��=�X��÷v����R�Pa�fL0O_ڨ�+%)6`�sG4ʓ]{��õA �!����獧1Z��۱�Y<�����c�.�`G#5М�82ږ[9r�@p#?��ױaP��&�e���~�P��#S����d
Bv �RGA�$�4�p"�@\ؤ%3��($�C6���N�Nh8�LN�l8�H�'��L�B�,$����P��`ٌ��1R0��0�&ߧ�@��mu�y�`�f<j���~  �q�I�'I� P�egփF�(�R:����
>)i�Ye'[>ZV��p�4k剽,��i[a�Ӆ'�Э��GZ�"VB�<����G�2;eAԺ)ƹx�^�+�^����Q��S�Dx�%9�E�tM> �M_u	@��C�!�3�\eH��м;�	�%L��쎯IB�xD�UK�OH�'#D)��Z�ۀ��4��CG�D�O����i�j��"<WE�;,�%���~|L���D~"[�@�ȹ�ta�Z2ѱ'�̘22�6-)7ۮ6�ƣ�~R�O�p���$�?�gG��� ņK�6nG�'!؀@�+��Rm���Q)cv�z�(D;qzD�|�8d{�q�'� &!A#N�!0�RA�J�� �5��"A*��	>Qq��SC�'V�t	`-�+&/��@�3tm�ir`�X���G�Z���Ē�N�?arq�����ɗC�SE���U�W�|��5A�<�Q�;Q��
����-1D����M7j��4LAi��G\�(�Xt�OR�F��B�m�Dl01���F<��B��9?��(�h&Y���dj�x}a���2�� �'��*p�ىL&޹R"!G�=�X�Cݴ~E.5:���+w
�O�]hp.��nI˕n�VzPH�ӧ؃3t)3OϬٶ�R��^��&<:�I��rs��X�e�ȟ���b2�$�1�X�Hw�ʹ�?	7,F_�,�b�-7�*\٧�wyr����h)�tm��*\����G�(OpM�����!,�h�DG??ڑ��)��'J��"�)�Y�|"��n4z��݄m ^h` ��Y��:7�V�h�L��&ƨO�����3��nJ�r�"Q`b���n�Q�&#'3�&�)!#���'&<M�QF.��	�g��,up�xp�r��T��/�Ov���D?j6���
7\dj����P�$"�'n~�藬�5J�>����O"Hp��ߚ^���O"Ir��Ϻ	�]�@�ӏa8P� *�!?{��� gl`M)A��Kk��OM�N�v��ƴRD<����-��I�x!ueU��?9��&w����AǞ4�LCqyR�'�@y�h@MExB���=�(O�ų$�V0m�6��Vc$>��m@��N��'<J�ڂ���V��G�D�Ɉ	�-A􋞅(w3��ҩ$4���TI�2?�XF}rO�3m,�H�weޱ���ϔjNr!�k�5� �CU�;+8~L��P���Az�T�YN�$M�7,,�pөL�N��+ fD�o漩W$,wu����C�*����SHܨ����':2��Ŕ�W�@�c���o��$/�2�����wPj@�e�������:���Z-�?Q����:T�`)VL��۲
�p���	/1�PL�jմ޺,��סi���גxR�c��9�#�ڟf�(r��8��L� �k`��O� ����c���@�'v� �O*Q�����#�JM�.H�W��qB5#��@K�OZ��nN(��D�$OG�i�FU��f �T"bi�s��'rt���`D�-��G}"*��{'��z�w�dB+Џ-��Ri���xT�A6��G��^�®D[D�^���(S�::����� 7Ҡ]����	N<�ēU�R4�t�(p{bk	��}�aV���'�- �$���.��,"�,�5"��kgyՈ6~X�ڃ�@3X� ������`��}(5�� (����`�m�z�l��'Y���ď�1q�
�)�P9"m�M�,OĬ(��: e���3�C�-�0�e�I5�����Y��|@�S��Sgi>���x�<�G��N٠�ܡV�� dGN�pAƗ�qn�����=*e�D~r��+r>�ͻv�.�9��ȴwZ��g�*r����'��l�?E����� |���-��q��,A�xȉp�	/y�n ���I�Z���I(p��#dଚR�]�H� a�-��w���'=2��|�bZ�6�2 ��E�(��q�9x+z�0bl9-<a�Lֳ��I����*cF&���-Ad<9� ��o�ax���T�s`cǧobܛ �5��đ�]F��ugPW8�&n�;DQ����*@>TF|�5d�� ���q�;-��ɐu�B})��Q�i�m��KL6'�X[�&ķ"��y�@Ȅ�5�D>p%*�sA
Вf0x���ܬKAK�
7p���ߊTP�0�ȓ��h(@�$p�\0IƊuz"I��p����Q�Y�Nq�5XՆ��G�P�ȓ#:p@��aM�U�����E	A�
̄�ev�{����c�\�8'C�#bR��ȓ$�
�k���Bi�Ё�=S� e��S�? ��k�#0�uC�A�1>�<�"O��d�Krz�-�s�}�t�3"O�٩���+$�*����B����"O��t�ë=�4y;��ԝ2A��"O��!�n(��!��$0 ��"O�����V���U��P`��y��Ʀ*L�L���W�P}s�$��y�͟"mwY�@�&}@8Aq�JS��yB������O�!'vE�e*N��yr\�B��K ����`�$8r�'��!`�.^!%ܱ12��3k�~@�
�'B��D+U ���☎6�\�C�'���@����j��ѣa��D�A�'�hy12���Pe�c��atS�'�@@�H�3v��R�-s���0�' ����΄���!�BT0li�j�'��%�/Bh���b�Sj�x�'1>ܒf�@�q��R�Y� ��'��Q"�<�,�1�ΐ~�2$��'j$���
"�)� +"��uq�'z" ���FzMc�A�*Di�I�':�$7D/9n��f^?;���J�'f�*f�*l)��#�gכH���'� %���'D��XUE�^,`�'�j$��'��H��M�4�U�r�Y�'�P��LI4z
���aˆU�0l�'� `��d��]�N}�ӥ�;�����'_�	kQCH�&&���7�� �����'H (�+]�E��U��B�0;r��	�'�,�bצ[S�BM	F�ڵ"'J�'4��00�{����V�="��R
�'/�̛C�G6ߢ�1��&H,��'��}�R�ؤ@lZ�A����']Z����C�ia`aH֫LV%��'�d���N����{w��:Lm��'�н��%Y�q�����:wǤ�'��2b�kGZ`��+i���0	�'�2��ăE	!��B6!Z9��I`	�'�x���� �&-�*T�7���:	�'-��Ӭ	8|8�0E 3O��q�'�9*��:�6 ���Ǎ.�(���'|�{c���H�d$�"D��
�'D<i�6A��+ap��G¶^��
�'f��ƃ�1�Ũ�O]$	$�b
�'���	�ߖ��]��U8�< 	
�'t�r�lA4hY��� ���I��'�B�@�B6���g
��'�H��5�&��"�"hV����'��!w�_�76�
�bŊ[��r�'��m�ԯFRB^�)�CT��:�J�'%pA���D�zu�I�%�([�'���B\�0A´ ��)|��
�'>��(&�ן#����H$�N(	�'dNh@dNѢ'T��Ґ#��q�'?��*� &c }�0�fR8�
�'���ᏉN����G�[�.���'1J�r ŗ�^��l	�O���',�u� W�}�� c��r����'�N��f�,\��q@"�Ey� R�'#���JD�ٲu+���nN
���'<��3��;�(u
�c޼i�Z4�'�	b��S#Q� ���c�����'�%ad�_�}ݼ��k�8a}�D��'b��C�/%<�"J�$'������ �����p���j��<�U��"O�M�1&��J���#ri�9$N���"O6����6�\xb��o"�Pw"O``�-Ԃl�i��F_�J�;0"O�ѺG@�]y��(�IP����"O�<����t�p�t�ѽ?��P�"Ol�B+Q�L	�A��Q��"O(}���3tސ�u!�=�p��"O�Bv�	,�Yh�O	%4�ěs"O�e³����Q[�.;��2�'��O$ԛă��%Ȭ1'@�r��Ek#"O��E�-am�	H�l@A\T��"O��E�D�M#pmZ;*���"ONcFl_�3,ġ;2
��z(H+�"O�T�W��Ii>��/�c	$��&�'��*>�)I�M�)h�)@��r��ȓb�
���j&�"wh�M���ȓH<����
+�6	Г�Io��m��X�=�!$-+;��K0^�Ld<���m��5I�!�34����y-�Ɇ�J}Qh7,51�r1*̍C ���1�P��wr���Y�OC"���C�<!��־b�9!��&W+~·�]~�<)&�F��)���V R,�E �LQa�<i�IΪ�"�7���#�ppÔIP^�<餈ֺ|��
נrp[�l���5��ϸ�����,ȷ�jȬ�@��� ���8����ġ>�5c�('rd�gD�H��`�g�y�<9���~0�Mb�煆N�>P
�nt�<!�bƖHk�h�揜~nT"R͖r�<	%�������=�����F�<���Y-	02y��\�e�tt!h�<�w���W�6u�3��#t�M!uM�b�<Q�#Noj���L�1�j�e�]W�<��N^�*Z5��U�R�ub�B��%�"��a`8cVR	:�
�+~��B�I�&Kv͹�	�7!$-�7M��*M�B�_�l@��GS����8��B�I�B�4�GD��r����IPs�B䉭`*��bǭ��V\�|31��MP����e��Ӱ�_�.h$�k�$��@Q3��&D��p-�m�4`� �%�8���%D�P�$� �̱a��\?KF���s�0D�lS��H�2Zm�@c>9-�l9��.D�X�Dc�0l���҇�&A �<��i/D���g��.6X0�eˍ]�Z�1�1D�,z�%�u/$�9ƃ
X� ])�B;D���/R(�f��@'a�!�S�9D��A�W�����C��kS�� $�OJ�'�5�PiT'"�8�)�
F��"�'�>YYv�M�v	>y��'^�9+�|��'�ĘJ��}�Ph��N�#�\�'Lh$,��HQ�%�JT�R�'���r%\=1v�Q���%@�pU �'�$��E)y(�,!�!��2���'�MR� �dV�9�T卌r��\C�'��� Κ=Z*���П4�� ��'���"`A�}���$ND:&Z]2�'ސ�Eo���p�gcY5vht0!�'@�⤇��3-���	n�����'��}�r�H�� \CDJ�Nt��'/���!@בk ��G�ȷE��T��'rL��g�H�75$"w�S�)q���O �=E�d���="�"q��k�pM��E_(�y
� ��s�o;9n9�����9����"O�9��z��h�F]I�.�(�"O�D���O�� 4�ѣ	
H#�tZ�"OZxxЊX����"�#�.~�`��"O�PAB��TbP�Ԉ�7!h��&"O�� G	�7�P����2��P�E"O 隤�
z��#��6ob���"O<} &k��t�#HfD�x"O �+��K>\2Ľْ�]���U�t�'�O��z�)�N�y�(	.$�p��"O ��'v�x�P�\g���*��-�S��yB�	7!�A��17��i f�B$�yҍ�X�4!�a��c$A@���=�y�	���C���6aR �I�'�y򢌌Bάxs��o���P��ybJѷ �&@;톡��ӆg\��y��b���!�Iª&��q�u�E!�y�Eͨc���틦(�]���ͅ�y���"[��G��@�P�g*�y2��Q7j��A�����p΅��hO|��	�t�Q�ɒ71�U�T/:�!�D��9`�)�[�1v�`E�B�d!��^���L�⇕�jf((�K��!�$L<�Z�b��R8�PWk���!�dJ >�����E�x�(�� �h�!�dW�2�l9(`e���@��k�!�ۊ/��Ś��ǂP�vɻB�ۉ�!�dD#r�~!��_�`�zp+�!�E\��,Ac�^�5�d*�*��nT!�G)����m�3?����?U�!�d�
�:�C���X�P�DQ�t�!��P�"Zd�B�4�L�J�a��Q�!��Ny�d{@�O�p�I� 
:��� ����c�  Ȁ�ӈ���'
az��#%#�@��"�抝�2�Ё�y��«h�
���(��F��G�"�yR����r 
T�ű �"�q)��y2GY�T����W�����a�!�?�'��}�O�~�
�!�!�9�"����*�yBf[.i��H���SiVd����+�yoO�����M*6��LZ�$��yM,$��|��ʄ|�D���EϮ�y���*4�� �r!I$sg���ꊮ�y�@�tp���//rV���dm �y�(�0Zw��E��m��A���y��-�Tm�E�L�_�ޭ�ԥ���yR2)B�ȘgN�"iĨ��֐�yR-  ,�%���l��J�y�_?5�@�tk�"t���b�!�yR�ĉLt�J��_ vV�Yg�8�y"��΄��C��i�hs%%��yR�P��	���ã`bĈv�yrH�Ly��Q)Ʊ\m
HJ�FL�y2)8/`����FL�U7�`%��yҢR;%�$Y�⌵EMڡHBM���yr'S+.�^9�c��:s��4���y�A�tkh�Q4b�9t�̙���y� �V`t�Cu`�����S�K��yBD�,_@���S����Flı�y���9�}q�胾(�L��bLÄ�y�D�
s<��]$��]iRO��y�E.sN S���"��0��#��y�^�p��j <v8{! B��y"�/s\X�W�X f��ER��y
� X� e��**�⋾r�� �'"Ov�Qg�	��(0����9���J�"OV0���l+����K=6����U"OA�
�^!z��9E��`8�"O|�#�X�2 �8`T�إa�0�6"O 	��&��]��� BI�
�(8F"O�`�ҋ��m}(�J�����z5�D"Or�s���'l��2e\�,�ڦ"O��G�{A�A
�,t%['"O&�!� ��$��i̥��3�"O�y���<��b��Ý+�$4�"O�yPu�F� q���C3z�<���"O��[DF�\x�"H}�8Dʂ"O��HeE��+���b��� &�Aآ"O��1���n1z`o�#@	~p�"O�A�bCP�*!X�A�M�A�N�z1"O���� 4$"52�&^*@8�ӂ"O�s�Ô�f��5ɗI�{�e�!"O0���o683A��16��y�"O�\��h0)#�͇bA^m��"OT��p@<2eг@�4*�8`"O�<�DI:�X�B� 9p��i�"O����Oπ%���T��<i��8�"OEyfJ�e��4����-mT�}{�"OdZp��,�V%�Bo
����"O�=�gdF�k�4(��OU%:�,p"OtLs�* �Ld�AJ��f�\��"OZԹ ĵ [�)��(�Isg"Op5�τ�͠	�$�K<V�X�k�"O$���k�?nXH��뉤)�މH�"O@���lHo��+'��?�te�e*Oj}��i��M�v��&I>Z(�'k�H��!	�S	���
̺6`�U
�'��0��@����ԏ,�n�Z�'��@��/��9�����.2+l��'�V�*�$�*<��HSt�V&����'�6-3O�-�Y��K1�P!Y�'Ξ9�M�#=:(��BǕr~�,��'�R h�´xf�ђ���e��|�
�'�U�G��4+U�)IR�A�\Iճ�'�$�pK[� Ҽ0�Ҧ�/Xl���'��Hj� 
�0�27�L�U^����'��|��D��M����L�\�B�'���U0i���V��$Ii���'k&����r��y+��� lH���'���g�X	Z�ްK0HS$e�Y��'�p����pi3�b�{¹��'=01���(tL��B����k�'o��8wi��BM!�!J=
]"t`�'R�`BqFѼ@��E�lR9�� �'.�#��F�~X4T+���21A� Q�'b`� #�q87oŁ,����'� e�C,ޕM�)��**����
�'�P�j��bW�U㴯�,x�A
�'4��Cv��!�,�t�bA#�'�`���HͧU�~����A�d# \��'!�����O�)�nQ�Dl��Za8�b�'IhQcǒ�\34�YM`H�''r�C�*b�T�2n��Tr:��
�']p%�ƿIJ�=��m��w:y8
�'��]���Q�+������ȇc�`���'�,Ȩ���&��a�W�]�6��':�0��X(�����MۻK4�}x�'2�h�LJ��z��F#X�8���  DCg�@�0��5�GX��E g"O"h�D��\� �� lضw���"Oư�p�[�:����K^4kb���"OޙY4\�qoz)p҉��Xj��"O��X��͝/2����%�� �t"O�Ђ陼D!ظI��4M<��"O����Ĕ:{����&��4��\K"O�i2&СWæ	�.B�m>�)��"O ,#î��jv��{�B͎'
r���"OH	%h�:1���Z!]4�<�j�"ON�Jf�
Z�6A��F�C��w"OJ��e�c�L9 s�_�D��Q�U"O\���3��rQ��1y1@"Ob�wjH�Z����N�\I���*OV\�2�I(��{��PL��	�'��	�DA%%=�(�F �;� l��'�p3�cW;(�J|��Y.@����'�PT� #�* ���A�$���`	�'� 1�㌊w�� ������	�'=B�0%E�<],b� �C�;����'38\��NR<�.L3$�fD^��'Ҟ9�D ��u�e��c�m��'_i���I�d�8��R�ʤ^ඍ��'���z�Γ��*	2���]%j$
�'Ϯ�K�KS�~�d����ҝT�.���'�^�$J�qp]�$��G����'0���)	�N��%�smW8
h�'zp��m<#F��S֧C��:�'ܪ���bϤ@S��"�I�8��`#
�'LBTxW%ɰa�@�rR C
@|:�p
�'�Bbem��Y��"�"�@U��I�'�0�2M <�bŀN�D���'��{�&\�G��)��b�1�P=�	�'sD���iJ�XsDkδ7t=�	�'S)r�@̂``t��8���'�͡�I�)T�q��(�)|����'�v��u��H}�CK�"mQPZ�'���فf�;A��@Jd�x��8�
�')J��ƌ,� 1:r�G�A��'�ZV ��1p�U�I��ի��ߐ�yRH@VN��A�P�6(Uy�+�y�ώ�RL���@�a��Ń����yR��<�~5�q��(8���e��y��
h��z��,p���oS��y�bX�Zd��O�y�t�qį�y"g2$/�B��#d�6�ȠH�2�yr�$q���1-Z�n�����9�yM&vc�ȅ� �c�!#u*��y"��c4��BR'�f?����y"(�rv��g��^�Lq�ϯ�y�^�o�@��d�D�J ,S����y��֍A_:`�bd�Wڸ�P�I�9�y��@�S����rg��x� \��G[��yr�B!^3J���ejC<�2����y�-@:p�4u�E̗OHj�����y��ΝH��8���ρD�����y2�A ���@O��@�
��y�j�n��"�&6�j�x&��y2i�'
`����#B-��*͌�y���RC�ǯ2b�`�ץ�v'�A��v�f0��Q&T��3j�.5n�ȓC��I�v�i����cF��ƅ�ȓk�J�i��Q�/� �ec	�"p*���|T��+��P&~�D��L.q�̆�S�? ���𡏥^�pI)�@��t�W"Or���J�P��q���%my�Y��"OSRoW�7���@�	`����"On����n�Kҍ9�.ċ�IY��y�"�$ ���h��#?"�1rဝ�y2S�qw0�U��*�r1`T3�y�Po �d��cĂ9�f�h��Z��yk� ~`Qӷj���(��7n�7�y��+I���(J� �`'-��y"B�����$�0y˰��6e��yR��}$
���ۭs��\Ж&�yR�K:<�BQ86��j��!�vm��y�I��}��a�WƓ':����y�G �|ds�H��
����k��y��:1���� T4�����yB�T)ʴd�%�wڠ�2l� �y#�/
" ����}��,q'c�/�y�Q`$�j �D s�$TZ��_-�y�OP:� ���Ԛ`�%��`ً�y�����E8�(]�8�s����y�"V�.>�cB�@�t�I����y��6VH��R!U�w@t];Q	ۋ�y"��r��L��k&w��-��j��y.}D�(i�\�ؖ�I!�y�ŌR{`��6�ИP>bqB���3�yR�C-PN�irsE*@���j��J��y�P�A�йZ3k9g(�f�V��y�C�yD�	����9z�� ۘ�y�̅� m���㒆m��Đ��U��yfV�Y�<��C]�|�7!�y��U���"E��U&��@�I&�yB	̪o$�r�ާ}���iֈ���yU���ܲ@�~�f��K�>�y�F@�:�<m�"N�JC�E?�yr	�a�|,H$�;Q�"k��y�'T�EX��(��D6T ����ԏ�yW�����5���q!C$�y�@�<��E�E2R��h��y��E�, �1�����@STDkVgD��yr*N�)��yG@�9�U�&aW=�y��#a�$iؔa��0t�4��[��y��=F0Q�D-H5P�0I&���y��Ӻ�X��t�+�\�"�� ��y"-Ў6QЙ� ��x�x�Μ��y�FnJ`��l
 v:����>�y��J	e� �AӅ�}�
pJ�!��y�,T��-[V�$�x	���yb,C ��iN4)kb���y��.]AM��KU%��mBWf;�y�D��W�������d�� �����y���;B
"3���0a;����'�yҬ�%� 0���@a������S
�y� ��	���y�� �pՖ����y��ƁGj���ϔ5�e�a��yb+C�Ƞ��d�?�x���J[��y��[-K*�T��Ύ	��Z��à�y"l��k`dJE�L���9�͊$�y2�͢oX4�u�Yofp�#a�#�y'�o�0e� �aN�x5����y"� ������D�T�����%ӈ�yr��I���'Gr^I�J���y��kƴ�r�ƅ5������y�k�5jI+u���4�4���HG�y�D .Y,����%���U	��y
� ����D8�C�E�d��0�G"ONP`���_e�\P�cS�#S@	zd"ON���]�H[Z�x��ܘqb�0ˇ"O����}12�4X�(�x��"O0�s��ϋ^J�ʵƛll�Y�w"O$b�{�E�SG��	X�@c"O��k �8p*��Y�f�	o�8��"O
��ɕ�k�Ÿ�R 5➑�"O�;�\�l�ZQw���uҰd��"O�L�х�'��]��G�6Z�b�+"O�ͱ"� =i86�"�U>z0`��"O��bv��<&8�h��Ӣ`-�a�f"O������U45k��3�I�T"O��&KۀH���!^�PWhL;�"O�tRW��) !@:%��-u\�]q�"Ofh; ɛ6]���q��� I&0�"Oʅ;dA�k2zl�É��Y)^��"O*��W�Y�N���0D�S���K�"O8�	fMS<˖��u� �L�<���"O4,c�,*]�b8H��(@L���"OF`4�P6_�v�{Î2/��Y�"OZ})"�U��( 
E�
T�� F"OP�2K�2Q�ܻG/P;�JD��"O���[�j�P�@1vH�ɰ��ô�yR�4A��xآ�R!g�@�3e��yb�)2n0]Ð�R:t�(�E�I��y����K���� Z�qO�pxeF���y�� ;+��Ȃ!N�aո��D
��y�h��'[��AV�$)���1芌�y�H��
r�D,�/+���@B��y�M�� ke�=��ؒQ&���y�ʓ�oz���	�p���eW��yR�GsCN��wG[ü��2�B'�y���?l�i	S���٤�����yN�
��a���Yު��7�y�-Q����G����Z���y�JY���̺�	��M[4採�y�E@�l�tiB��]%3�p2�(C��yRŇ�-��K�mD|9B�f��y�+�T�$���L�yϾ���aǎ�y�-���ba�u�ʄ#iİ�yf�� cA�u`B8$�r!�4�H��y�i\)Z@��ÀX��������y�
�~)�f����Y��X��y�ƠWITE{i�6�X$G2�y�ȓWDl�&��B���� ��y����#���`�D�O�p��Y��y�oܡ� �+�L��N"|��� ��yb�X@	���@G"?U��bJ�yB.-`I`�F�[�9�zHc�a�=�y"�Ɍhq�`�/-s���Go@�y���:L����'�Ш!������y"��I�}���V8Ghܿ�y�l�(j�0�l�� �P5o_��yBD��9��DB� Ӡ��!�̋�yR�ȄJkj�P0�
rI�j6C���y���;��t�ceX8\ר,�U�4�y�菽#G�EYA�� ��j�)M	�y2"T�$8('�CJ dx#B��yR�DRm6}���U�h��qiǈGH�<�d́3c����ϙ�\#�U6�LN�<��ǜ:����O"��C�J�N�<�р��E'~��i��W���k�J�<9&o�7\xs� '*4*HSK�<� XP�@N+1��	Dm��u,^�
"O6�ypƝ�+�z܂�nԋ(����"O�dX���	R���y/�F�"d�B"O�������$���^�f�
�E"O��94�ҷIҀ0��-�D�@ȳ"O���G�ë��%��-�k�L��"O�QŊQ�N�zij^��eOJ�a!��-r���Y/ *����6LP�E!�u~*D�D6m�%`�̛�R�!�D�5nΜ�s�L*LkZ���
$�!��4+�H`q�L�2^YR��!��u[!�D�9Gc~0f�1*�� �hA�t�!�D�>XNˏku.A����!�dΈ?��p$�C� ^�����Y�.!�dڟJ!K�"�-B[~}��%��!�UT6zF��adF�=XC���"O� �7���|_<,�Ţ�=>B�qZ�"Oґ�&�����Q��z�B�"O
����^U��<;e ),mz4�g"O�x���L�aH(��/L�\�-{r"O<8:�M�2�*�aů�]���j�"OIs�T�uk��k���I�a�C"O���'Q m~}0��O�!<9�c"O�00㯞&w�z�̏�s<@x�"OJ�kDN�$X��U#æؘj�A�a"Onl�iD�!�d��GI-F����"O�}K��A�I-*��6�Jik�]Q�"Ox�9��Ӏ���S".Ѥw�Lq�"O�yy�K#� B�>I��j�Ck!�����L�W��|��i�/�%W!��@P��9�
�>���b�g�G;!�D�}�Jy�a����A�y�!��7>�xI�%	�J�Ph��E:%�!�VmV�qR�רQ�pi�3e��~�!�D��o����l�!+���k�K7\�!�F8!�>� ��ΆT�a�("�!򄍵7����c��&1��#7�!�ă�
�`��ԻD⵺ԩ�;g�!�D�>�4�hT��=v���Aj���!�03ݚ4�s/�'�,@Sv�C� _!�$	#W����B��,�v �i�I�!��;0�P���
T��!���$n�!�O�=��D��j.��d@�3g�!�d��_H��� �y�q�� }�!�J9�]y��|w֘р�\Y�!��Z
L%p��//vT�I�B�9Y!�䇘]����自TB)�޵4�!�$��*\d8G$�&��� �p!���JF]�"1G� y��͝�!�$
k�詁���@Y��d���	�!��.��I�&�m�0�����!�d�#njd�Q�B9(�Ҁq쓒!�5ond᠈Ĺ/dй���j`!�$��z�^1H�MJ�3�z=�q�ՓT[!���C��ᕎ�
�Z��S��">!��F� ��ФP�*��4�&']W-!��z�6a��0W��B��ת%�!��Vl@h�_X ��ANF%�!�A+yǖ��`F� L@4*�L�'!�dИB���Ҍ�&�u��k��y�!�DU�)��5��Ĉ �P��Í�w�!�� =|�P)�C˙&��캧,Ζ\�!�dV��
a��K�,��{�k�-!�$��V��k�b�=�\�1!�� �`j��S*~���EL��#AL-à"O��YѤ�P��h)qd�F���T"O��� �;[��P
ѐ�� 8�"OTU�"F�Js���ɮ��"O��c���zVq�.ޭQl8H6"O4D���#M�0Aː;�L9r�"O�ճR�^&v�9!L��]�|�g"OX���!��/�⁺�ȑ0w~��"O�m(�� 0k�~x���N���"OF)�MR� ��1�f��Ӧ��*O�(���Àkʴ!�c�a�J)C�'V]pr�Ni����@�^%W�~\��'s��3@Ǜ�q�`���U[>��'��)�A�n�f�0���8/�h	�'�0�J�@ 
�ɻ�j�)��z�'�x�&��2�����R��8p��'6V5��aԊ�t%���S@�"�'6�ٰ��$�a!wi8=d���'n�Á���S���k���:	�E)�'wvl1���lc��P�.�:�@�'���iΟI��X)�ȅ�P���������g�
�
��E�ʌGN���ȓy`ɐ�Bٸz` D	�^�W#�L�ȓw֦��r�:
�0�0���	I�ȱ�ȓ?8�q� +��p�lŁq��t�ȓ�8}(3�����M� p�d`��=���M�,��s�nE8>n�d��(��q�C��g���E��`����ȓ4�j�� �ڸ�dnW�R��t=`�k5��7ư �'-��p��ND�ĉ���'g�����/����M��H�W
��a���͌+	�	��WȈ9����;)����'t~L��>���c�=V��+Q&�<=)�� ]�uS��(��Q��D^<�ȓ �qP(�#,�)��EN�;|l��6�[uB�h]�,p$�c/�u�ȓ��:�%P�M��"D8I �y��;�ኀ�g� ̡ �H�ܩ�ȓ)��e�נ)�(p���(Nr܄�g�P���@:2i���u~rՄȓP�C��ڤ$�P���V�vTɄȓ)�X�m��,��&C�=X:�ȓ-�����+Sr� i�%��R�L�ȓ^�ڭ�1�PnDxз)�:(	�(�ȓ�������_��ɳ�%��[�����G���9�c,�J�c�i����}�ȓ1��hP��Ky��Tb�WS��F'�)�&F��n���˱r���ȓ�y���Α7��(�V�M�4Jń�;�<Z���Εbы4L�ȓJ��@1�`�C�����ޅb-j��{��b��	E�
��%���l��ȓ2����@ǱL%� j��[=7�����6b08����}�ܱ��<B������d`��� oV!R'�ܸ�1�ȓ}0ST����@"�(7
�����#�Ȑ���U�U��m�-�3�����x���!"��>�6�G�vꄇȓ ����ᑧL�P�wNPfr⨇���Q�	Ւ_)&`kC�_�������D`��5�3b��ȓdY<kQc��85N���i����N���
M�"�I�3�G
&b@���S�? $i귦��V.��ԃ��:  �g"O��R�
\�9�U�J�I)��[�"O�2���R�ļ���ֹ8 D��"O(�i�?�q� -C�W1��S"Op<c�"�K��M�w���"����"O����m�"�A¤��2芁`"O@r%�#T��1��[D!Ru"O|�+RfL+o�e
�Ӭ%j��"O�S��
�qY�	B��.E6��G"OFh9CC��Q����s��,G��A�"O�b��^8Aa���C��w²HR"O�,����j��$�6���Ё"O~��ŉK'E-
���T
,`��"O�diDN���G�J �Ԃ�"O��Q��zpa�e&L�]�vX��"O����o�
)��Ӳ��/"��i"O�$3����[(��ZV$�"8pU3�"Ol�C��0F��]!�"C Nȴ�Q"O(x[�m8H�&c}�x�ča�<��Vq<�%��G
M�<�4a�<���^Z���TE�~j萁��S�<���̵-V5	7/�s�,a��M�<�a1�\)�2�u�9Vb�T�<a�o׌�,AZ�&�>�E㧈K�<�G'K4D�,AC���a��㖥�~�<Y���\;r����-8�z��{�<Y֤�#W�\����8���z�<�R`��Q'*<
�˚B��lZeL�t�<q�Ɍ�A�d����&8l"��Vq�<� ��2l̘ ��,It����j�<9R#^Q���%@��RX��eC[p�<i��"C�����U&
�Z�cv*Mi�<сe�$txܽ��m!t�¡���GM�<鑪�T�S��QUb����L�<a��N�"]��IW��E��I�d�<�c�I�E��Tٗr1~�Z�^�<��΀�[(�����WT�U�FG�a�<Qs䈧4k���Go�e.AR�N�]�<�5�NB�B�Z�@s�����Hs�<Av`�=`��h�>'R�C�D�<A�̕�[�dP���H
�z��E�<��`��hӤћ��aՐ���NEG�<1�"��
�<9�H�خ	[��YA�<1�ސW���[�I����v�^h�<��لjܜ��J�#���!t�b�<q��]�2�q Oڇ-�&a��`�<��$S�*B��yǡPO�ʱK��a�<����5��j�/\�˓�_�<��F�>(��8I4z���SDM�^�<����'��N�6Bd����A[�<1���l��1�D1"�R�k@o�W�<	���Ka$(�#��vB��PCQ]�<�V�l<�k0���I�HT�c`�^�<��o�-���&��*; \��i	A�<�`�U�|�6�X�
��w$p����T�<"�� �I6/]#{+����*DN�<��K�&��2�F��@�'p�<�!��?�X�Y�菗nym�-Kn�<��![.%�f��F��JFhD�q��r�<3�,V��
%�քZp����
H�<��b
#H�lzW&�M��C��C�<��"��uP�I���ړ7��4��aFg�<I 	�(o�X�3M��	�n��-D�IA�Y�3Ϥi�H�nJLuQI&D�� �Lb��gک�&9/t�!"O�X��wft	��h *z2!"O�4[qC�O�)y'-Y$A�$"O `�Lc>𳅆�2Y�}�D"O<�#�+_Dm�ǅ]��NI�F"O�D&�P8	<$��c�&_|�<8�"O�����?1T����@�<?m�B�"O��Q/�"��� �Q�y;�"Ov9��B(0<�֍S�S��`"Oh�AրK�N�2���0IB�I�"Ob�{B�U:���0��"M�2�u"O����QM.4���(����`"O~��,`�.�%�E>k(�b�"Ox���b
�90,��(Q_��c�"O�d	bI_+,�l���;_e
l�#"OT8��V�t�B�c�F�N�`���"O1i�h�54�$Բ��߉Yy��2"O�-��� *l�����. ^0l�&"O��a����x���W��3f"O8�� /D�5�1�R)hqnp0@"O��s�S%Ƒ8Ca�9ol8)"Of	��(��=�s7�CaH<�"O�����б.���/�+J4I�!"O����F�٘1S���Rc��{�"ONE�B��4�&��"�qK��! "O6E�`#@�tf$����Dv.���"O���1��F]��X�$�2K����"O,��s�ٳs���d@�#=��0"OR!a1��(��T�D�=���"O�!�
E�Z�0h;B�×(�&HiE"OB��h�� ��S�
�7�V9q"O􈔤��<~�=z���.0����d"OJ!���E4 ��$A�AF.>�^��&"Oڐ���fp<�E���&�B}��"O�H���>�Q;�e>�P4�"O�U����%0Xp 2/"��[�"O�ӂ6��i��Awg,�Z�"O^�!bΗ�4W���A�D�Uȵ"O�0#G�۫:�	;�	 튡�"OLHb�̚t�"��2N�#�*)z�"O, ѣ�t��H�vl��Z�"�q�"O���BO�=T��Q��]�<hQ"OSt@�T��0��'+�Zy!�"O�bS�h�JA�2�^�}����"O�d8&J�'B9<q�
ɇ4�:`"Ob��\�	ކz"�<E�|Q�S"O�ŉ3���\�x��һ��I1"O~�PC�8Ar�(&��+��eP"O�0xGf!H�(�O�%R��z�"O �'FQ����s��;��dK%"OXA��/9?߸Y:��<�P"O�2bӠ$1�Ѫٿ<�-�@"O��2�d��1���3�� "O*5	�V�IƔ ��%�2H�"O�h���]�x8���k��0r"O�#�l��^�|�zG�<a�f���"Odq�d#Eؼ��W�e)�t)�"Or8c���(����1���t8a�"O�rB�H�I��ȱG��J}44��"Op`�2���'<i+���:Y�Pᨶ"O��)w�x-����'��� "O���#d�<&h,-���E�b�AA"O�,�&$�-AL~�ɡ��2�
�q3"OH�� 2�(B�fՈL|j�`A"O� ��ÔE�.r�����%%L�x�q"O����7"��3feoEP�z��'k���R�D�9��/��0v�y�=D���j�(�<颁 (,�Z��h;D�2��[�5�&}��-B�}�:@K� :D�Lڷ�!%È4ȁ�\ t+x�@�<D��
�K��3��M��J\CE4C�;D����`��;���a�Xc2ȕAa$8D�0
r+�)50�,H�h�+h�൒�%7D�|����1���IES�*�ӱ�!�	l�'��	= �t P�Oϻu�4�@�*�O��B�Ɂwah�S�Mϥ���4$�*_�B�ɬ$�$M��k�3��a�2m�.5��B�	��D��.�1+�A��/
�_Y�B�ɤ�X���$�h]��7ȦB�I�EE.� �G�^c���E��h0�B�I"1�R�p!�m^r�����nB��,,�n�0u��4�P�H�#c6B�	��]I"M�R">�'�u��C�I�8*s.��w�p�����_e�C�Ƀ>zp)	��9k��QCŜ�\bhB䉤C��<���\��Ƨ� �B�I��D�@�lZ2L|e���=]�HB�ɑ%���v�˥! j�PGG:0CZB䉞Qu8�3�+@�R�:��4�#r�XB�I?uz�u�������ev�B䉘Vj]9� P a�9���_�D�B䉉��R�?\x��`�L?.C�ɦ��'
?Q�8��V&VB�I�$n���Rdˬ'���2�� 
����<I�'��p @ǂ�#�xI��@�B��X���x���3c�Q�`^�^(y�C_��y��ke�����*D�>1�tj�5�yB��N�eq`�Ȕ6��#̈�y�`��6�v����Z>H�L{��5�y�iӊReY�$��8�hB�����y"�V8c�ZPX�I��.E:h�$�yB&�PY,�H�@
	�H��c[�y��ҝM��hP���p�J�H�"��y2b��-H��+�-Ѱ~��ԑ��y��ʙ'j��b��طK�h\�@)��y���4k~ 	�A�4hz10��1�y�M��ua@�#��
0(�]���@4�y��&*0���ᩅ)!IƠ�9��=1(O��I�r���r���XK�N�?a�C�?� �y��^��U�*֋�����'�HՒ�N(5f��"�QC�1�':T|�fM)&Wt僴ĎY̌�A�'`�Hү͌uڀ1iC��eu8��'�V�A�I˚c�����D�S���	�'l|µCɅ.@qCf��4���	�'J&�rgÓx|(qgG*)��a[	�'H�պiR�y� ��Hҵ��@�'D�t��o�<�����̢���'>�-pg��}d�@�ˈ��m��'��9f,�tE��"�2$�z�'P�� ��S�Q*F��	��Y��'��m�2�N�g�H ¥��Tg���',���x��)�/!<��H���xR�ҁdpT�Ԡ?̠��[��y��������5�	b�.Ѻ�y�jR�wӌ��' �xoP`��� ��y�@�Oe���������y"ÛW��e���0��ò�'�y
� ��K"�L(���E<n��܊�'j�D�AX��LZ�`S�i�6!�$�!B�T,�ф�	1C>t��J2Y!�d�Rc���2Cʘ=�"DV�;!�$�(8|�$e��&�ޜ��ԛF�!�Č�w9��!��ڮ0�zH��ߟI|!�$@�D��ԑ���7�P�;���_w!�
�(���u��8*���Z��
@h!���shf�귈��)꼱����8!���
-0�Y,� \�bf��2�!�D߅ ;�dp�ctV\QSP��!���D���9$aD$rE�	ڳ�[��!� |�(�`6C�u���;�/ƙp�!�D�;f��x�K11�h@�-J�x�!�d����oG����z�lB(=!�ƜN��Xh`뙿Gx��r�
:�O����2?UZ9H	��Yې�$Zu!�DG�/�Xi�a�#چX��N�:Q!�dW�J<�5�E�].onB!��,l7!�؟-`�\cQ)J�mba�DGMB!�$yw�5��I��`�	����!򤟆N?�,� �.��U�P�N�!�R�?��U�A3�Ne9%`�4�!�A$B(�4��@ĭ��9�4h�!�$S���$+�͚�~�>i$�@�!�'�X+@�p-���ރ/�!�D�C �@
DLz�� ���*/k!��13�d��:>ܹ&o/}O!�D�H8%Z���2xg(�%�ʜ@!�D��/�h�&	�t`Fi��
I"s?!�Dǲ}�mh$��o�� 	;]&!��Y�Q����J�[WŠ���J !��F�24Z�p�`ڽ6vx��J^�q!�D޴�]��K7Ig��D@5!򄁡KP`���R�Z�P)�A��!�K���s�"H�g�P���
ԶM!�D"5�����Р">����¬v8!�D��!K� ����%s�հ�מt$!���vi�X����E�Zq!�dзo���� �Z@f<
��R�!�D�S�J���h�R�u�$>!��;�~�Є-S7��L�b[�\�!�䛩��C�̓fFkQ'�D�!�dīO��M��J���䆚�o�!�D��2����ٰ]x4�q%�%P�!��� ���)��']A���#$ӡN�!�D�9{~�3�D�qh\�'A�&s�!�ǇK�~$��@;o�8��D`���!򄋒8��$A�(Q�u(dU8�.з"�!�$��(lx<��M�.t��01\H�!�D���)(�	��=T�PK���$Hr!���&e��)��݃hOܹ�$��U!�d�/_qGY�sX���	�n�!��7U�*İ�n��A��Q:&�>�!�D�r>�@�!C��>��9�T&��p�!�$�!�l[� עT�Ig��B!�d[z�e��دP{���5蛫, !��Φ!�&�ӅAt�(�5B1;�!��ɾl�����$߱_���@���!��^Ŝ��Wa��{��]q�C�*�!��<H��}adO4Q2}�d��( �!�>)��I�'�S/+�>�0�Ƚs�!�$�:���P�ŏ�4C�$z��C�/�!�W6c�A	��J\&��C� ġcL!�� (b%G��� �.��j Ńe"Or]Af�@�i
h�`T�
�/��@B"O�9�bA�i�" iq�I�z��"On$A���->��H�֏�"����"O��e*�$p��0 NK�|�bd"O�y�c�&Qz���d��19�"O����O������)��G�
�:0"O��j�������L6G�25��"OX����'�셲E�E��lS$"O�	�T@/vn�W����4Bw"Op@p��k��C�aA�K2�1��"OP�e�;F�d���o:�R�!�DPu�N�B �:I���U���!�G�9�lD�s,�'k���V�Y*�!�ĕ/vH��eM B�"X2���:^!���8#���1�F�� $���jU!��oP@�F�[�kpd@���9d�!��*E��\�׀idh��q���;!�DE,u 0S�J�Ml���s*�(H3!��[
�
�[��N&=�5*]�!�$��j
�jN9a�by���4!�D�B�T��Bʰ)�FW��!�d���$��E�8����}!��84K$�q�*�	�&���Gc!��ݙ*�<�;ńʯCϤ�3-���!�́F9|�bB���'ɊqX�A�CF!�䜥�*�C��U��ukӀ�p�!��d?��E�Z�z��� @�"r!��S��P����5T���2 �"�!�$Y32gj0����MS@$��;�!�D��@��!��h���-پ$�!�B�����zs���;��C�	M��	����9\�
ŭ �4~C�	�e�X8�a�������� 4S�B��jh���'#ů����Ă�4tB�Ɍ'x(p��/p�x&���HB�I1�X��Q�Ωq9���g֗t,�C�I���Ă�����I�T�*�B�	;k��H��B*� C�6ϪC䉾���ق`�mæ��FHЭ.M4B�	��:ᑲH��JfڌrG���DC�	>f���^�bB�(��_GC�ɱ!�ư���W+;��A���r`�B䉺=V�XG��3���@�-Z�B�Ɋ~A��WB̿����A6d�nB�I�@��#e��P������t� C䉞 q:��V>)��3��@��B䉇,l��c#�&GlhU���J���B�I�a!��RG!H�-����$	� �*B�	)L�bSG
�r+�M��Ɛ�P��C䉢[��x�Ц�<,*�=Kׄ�_�B�ɠI�ʗ�ּ �zQk �߸n�|B�I�X���C�@�1�N������F�pB��_j�y��K��<�Yr��g�PB�I�b���k(����\�lB�	;9��ɕ�Y�H�ҡ
�T4JB�	�5�̡��]T��kV��T�B�	5~��<�'���{=d$���R7d��C�I���zh�-=\�� �5&�C�	�y�%`T�	Vo�%*��˝dn�C�	<f�ı�DH�lʉ;QDɿ#KB�9�tŊ��߬}��p���ZF�C�ɠ�V�A��H؝�B@�b�2B�I�8l�5��7p���b�nŐX@C�)� ̠8�c3+H�,�U��$Ҍ*c"O���bD�\�̝ĊO<��
�"O�����,D5�{e�?�*9��"OZ�b�I�k��(a��<tɦq�"OXи�F*\���l�{�v�y�"O 0�υ!ڈyà�!�$i�"O�	�t�[ W�(۷�0��mj"O�@s�L+]&�1kV�նm��i0�"OХ��-�	��lje�D)	���C"O�4	��p �'O�Z�D�v"O�A03�]'��L��v��E�w"O�}��l8�iE-t�98"O
�J�HF/��$�(k��t"O�U�(\�ܴA�-��$6xrE"OU"��O�w��A��mJ� 7��*b"O�h��N�m�P9��J�/3�H��"O�8�B�)a���It�RP 郡"Ol�I�#Af������$[�AU"O��� &D��D�q*/q:�+4"O�����X7�;�W���F"O�P�B@��u~��zǁO�cV|[�"OP8���ǓU2��f��'.�R�R1"O�h��
�jc!�?V��$�"O��B��M���bbT�u���#�"OThأV�e�DM��ҏ;��� "O������6�:ucZ9Q0��`"Ot`#�O-I�B0�d��?3j96"Or�p��kQFI1���W�*��"On���d	!�> ��1�"O��(�̌�t���G	�H]�E"O65i�Z�DE�K���6a�Ѵ"O��w�޴m&m`J��`E�"O��#��4�BHz$g��>�\4ч"O p���ѦJ����pf�&*��C"O>P�پ{�Ld�ԪG�f�2�"O.�R�ؠ/l���G�vI��"Od y2ˁ�rejV�ٷf�^���"O,���R%g�Q�t&�A��'��� g�O�fu�p���$�	�'��`j!
D� �Tii�LL	6 U��')�	��J�%;�x�'M��{t�!9�'�:���I)"��8���wM�X�'�`Q���0�H�ZR��u�,A��'4@��(��@���3v��2�'��H�bb�*kc|��W�=ET�8�'�`�>g+.�z6N�5[���
�'Yj%+EjͲu��D�0�Ս3��uJ�'Z�:G�C�}Kt����C��!�ȓ!�P�s��k��8@�%T��܇�X�̄�#ȓ	�h�g��� ���5K\]Re�<!,��ZҪ3.m��.�@���
���
����ȓ<�0}I�%h��X"p�Ӗ��(�ȓY>�p�nC3gBv�:FL�w����z���kQ���"�V��$F楄�.0vx* /ҏrZ�q���E ��ȓ}֠��3���x޶H�� LxP��sǤx�Ƭ�#:����Ш�.BA�<��):�� K�"`ެ��GB�<�A/	�P	p�S�=��Q�S~�<�4k�* (�t�B��]�!��|�<�2��9���caHN4)|LPf��N�<95��?!�.l�V/D����EI�<��jI.u�z��5g2sm�9+�HK^�<� J\�wo��~uaP�NԔD�2y"OV�hJ^4V�����
,��"Or9���ՈK�Tz��۴2o�	�"O��`fB#:��B�,L
!^z�S�"O�-���+5�`l9!J6B@��X"O^e��]3�%yb�Q�U��H�"O���0/�bl���֣�E"O�]YU劚Ò���<s$��w"O��3d%K7	��+�C��($"ђe"Ot5�3i9Y�4;��Ҍ8�i�#"OX��H�D�X)�5jC�}yХ�F"O%P��Bb�T AO��bm��3�"O�!�1E�y�ZI��'��Wc2"O�q�0��`�xР`H�1ax� �"O�� E	S��1��t����"OrP�t�ZVɊa����Tѣ%"O,j�CM* c�X������"S"O��"��=���q�A�~��MB"O5k� x>5�W��:�V존"O����f;�Z͈y3���"O���eo�:uhB΍3*'n� "O�T{�^>9�,4k�K�'"^e��"OVɺtLE>pCX�4)� �e"O�Ib_�R�n�a��#��E"O	�CdN�"��\��/n3��"Of8a�m� E�P�bh�!�\�"O$!8���$wT��'E�<i��W"Of���k��fJ
��E %ļy�"ON�q#GPn��i(�d����x"Ot	�w�ўM�
ِ�� �~p�jP"O�]�k�7G�rIQ#D�8W�Ų�"O&T[aB��I���;�i�%p8>�Bq"O��
�%��D�2JP��"O��+����~Od%3��M�> htA"O��ǆŚH=�-�� �5H�s�"O��b$Ym�:��Ca�+��!�"O�}�'�.^��0k4�$&��!"O��s5IX6s%�� �?ljH�3"OH��$V�M\�R2/D�
�&]�R"O(36	�?nKZ�qu+Z!:�ȓv�*��q Ya���@6D@��J���*���#� �*��� W����ȓ!0��#N��G�L5�$C��/D��p��](V�e�!'�A�pl#D���c��,j�SD�H��=��/4D�t[��"v/&������w��њ�4D��
&�H�Z��t������r��0D�dr�޽U���ivmsxac!g+D����.�&G�0�*WG�1/rT�i�i)D� p!"U:3c�h��a..��p�%D�4Qsn��d�(p��/ЙC霼���$D��Ga�Caޡ�J�Db�q�G/D���D� �"�p��˗ah}��M,D�h1BB�:sl�2�̖��@��)D��� f̄�"S�u+ڸƥ*D�X���'wx(���Ͽ �$a�3D��`/H5hB�l�7Ǆyɱ/D�������=�^�a�Lʋ�XɃ�7D���DyôX��`�=BBp�w�4D��hP#�5�zY!�0UX4⑆1D��K��H�_He:�@�>+BRb�/D��C�͝>\S!ED�B;�ip'2D�������E�Ӌ8X��u��%D��#$ͩo��jO�A*��Yd�%D�� J�;� �d�ƍC��A�
ي"O
1jB�ʶo��p� S9�R	�"O� � $��ɠ�ϑQ��,Pa"Oڸ넇�d����C��,�4���"O̽���)p��2�aS3S�p)�'"O�8��j¬v"2��OG�L��!r6"O�u�f�[���6�liy'"O8�g��>A�q0�kH�2��q�"O ��b��a/�|���3Vq8���"O� "�OD N�	'�A;gb��"O�(H���R��
��\	�Fё�"ODxP�	2X�ypF)`���R"O"��N�x� ��f�&�Z�X�"O��hӶ�4� �z�H��"O��`���M���� �A �`��"O�]�DN�G*cC-R�zț�"Ob�G��xv9��˙���R"OL��С�E��T�֩>~�2�"Oέ		@tjddI�Q��Xk�"O|x�%V@
T		����"OL���M!�j��ǘ;o�ճe"O:aaa��9!YDM�$�R�S���90"O"h8@EW:)�r-2�L�|HR�"O�Y��I%(�2�`�#�D�9�"Oh�ZV L4tb��\}���ju"O�<�fC�n����S�P��ꕑ"O�����D�"Ծ��C����!"Ot`�*S�~�J�c�#9����"O�i(���Q�gc������"Odx�d���ʩk��)���9V"O4���Y�T�y��Ưs�D��"O��࡞�190��#H^R��� "O�)2X0|����@��sB�=��"O�h	$�O���E��""[d��"O&hɒN��$�����[H2��"O��#�}�Vl�Q�֙34�`Z"O�U�
�/I%��D)��V򅂓"O��b+6S�^X���u���s"O2��cؘ��঩۽}��TAT"O��*��� n�pda@��y��A�e"O�a�oG�V��8�U<q�f ڤ"O���g�Kz�a⤎�aҺ5ۤ"O��8S▶1��Pk!m��S�T�g"O��C7lQ�ܸ�yցf�*-�V"OB�3",K�L�ņ�b�$�)�"O.|��߯E��DЅϲ�Y�
O�6��t`����2$�VAáa�=�!�� %�\�����f���+�'V`2Op0�e��@���E<\�X�"O,a�%��+h�8�,��uLBd�#"O��d��G��YSqM�<"O��:e�^�q)��3��������1Ӓ�A3DvCva��u����F�Z��%�[*U|d�2��+ ����*�4iσӒ�RR��>P�$)��}^lіƂ�a��]*��2m�:���u���E�+z֔�F2?Slņ�k� 1H��Q��)�C�Y��$����}��ԙ:0�i4%�)M��I��m}t��`Y� 	$TA��h�9�ȓWa�(��aئ�.�
��V?9Y�!�ȓ��������d�^�{�HFV�U�ȓ&iX}�L^�TƼ�+�K���ȓy���g�ۗW��t��|.T��S�? ������6*�����M�z���"Or	�,�0:�����׉^�Ԛ�"O��j�M%�iq���[��4��"O$P�6ćt"d�T�D#3*^%��"O@���3C´��E$�\�y�"Oİ �E��xxQ�/r��$"O,q'�W�ڨ���J
*a�"O��R��W��N��P H����"OB�c`�ζAXd{2B:�"��"O���P�gh8�*V4�̥P�"O`�z7�R6Rj���@�(k�X��"O���oñT�T��`�0 ����"O:�sE�5I\�3.ޔ'Ҫ�"*O��"�Z9%o�4A�L.cL$
�'�����),d��`�o�Z���#�')br�Ջ7��Q�]�F�����'o��b�� r@Y�-�E��
�'�:Is�� �JDr����A��0H�'�P���f�0���`�]�4ڶ��'�8��(=,� �IA`uVQj�'�P�#�C���=�AK�/�:�'�j-R�ʅ�X�|��`��x�j�2�'ʦDj��~)r�Pw�F�jNFݙ�'�,��L��+��kݢHt `�'�ĸxaa�j@�<*��UoL���'qL�Y�:`!�䊥��!uJ���'�u[g���*U>�J%آsbd�
�'r�	��U)�
ݚ4Ŝ.X錘�	�'�~��w��PG��bcM2x\r�z�'�,b`-0Lۦ�B �mX�X�'\�9��O�?B�e�N�1>�i
�'�~ԉ�hI<f��8�b*A�.��1k
�'u21a%cА>�����i�Q����
�'�K�yU��b��1z2��Q�<)7ϙ�R PBE�PWH���(�M�<�� ��_�<�5*�kF(�y�oDL�<Q�&U�z�J�³�N�4Sz\��*c�<�7bpw�JA���o��|�#�j�'�y��/������9Yh�$�� Ǧ�yB�A� Q$4��f$R����=�y�[h���R
Q���b�%���ybcJ�8��Hxc�ĜE�v�t���yb�F�¬D�a�$+����f���y«��lj*��^�V����q�.�y"BŮL����֯�0(������y"I�#.;��UO�%F#��r$��y�HS�Z
�j��X�EB �����y�!B*/��%ZƩM�EUT������yRKS��`��@>�:�ie�N�y"�ό ��h{@�ȗ$���ӭ�%�y��d��S� ��^�k �K�y"�	o���qᙝ�������y�d�;K��-Z���R���yb!�Ho���5�	H�I1�T��y��^��|�"/H>M�R �7Ɗ��y�D[@@Q��gO,e�	*'OE8�y�eG�WRơBQ
�|���)�I���y��/�H�f���g?�샶X��y�̑<�j* ��*�|صEY��OL��ȢJ��h���	A�b8PEb�!�DV9ef�$ȠD�H���P��_J�!�DL-�\iQHO*��8�%G�!�$\"�$qcUN��2�0�O��_
!�D.h2��I�4�L��eKO9s�!�� ���Q�;�H��f�-D��5��"O�Aې� 	A�dFo��^�H��"O�(�jF�g���-�>���8b"O�,+�M�)�^M�'�7>��L�G"O$�F���]��B�����"O �T�Z>MN`D��g]����A�"O�Y2%֥5�$�w�E�-K�k%"O���V�6SB Dh��FK4`��p"O,�0F��8��y0�(l(L "Of		��S�;:9���]<Gufc�"OJ�d]V!���jD��3F"O8D�%eQ�G��xr�E�CR.�"O���(ݨ��9��٢,��% �"O\	��"�&���C�G�)!��8�"Oܬ�wn�br�wmȽYZ�q3"O�mpC_P~l4� B�2�L��D"O D�eҋ+�L��A���,���5"O��|Z�C5�ʻ���pn�v�<YEւn`8�U��*P��}�<a��ۭ S��vBH&(r"£�C�<���Y--n0a�$'��i��-~�<����n��K'��) "b�h�t�<�D>
�R����G*��e1�#�m�<��̜�4Az$%ٴ0&5��A�b�<��(J?�Y!W�I�Y�^�	�N�W�<I��3B���֠Md瞱��!V�<�3����\�֣_$~~,�4f�Q�<ˉ158hXpMY�eQ��@&R�<�cvj*F��7������Y�<�7Œ2Bh۰ʯ)r��`�U�<&�F
/A��S"���(��a����M�<q���@@#��N%fV1@�h�N�<	�"%��P3�J�5�FmM�<1��[ ܼP5�L9�j�`�J�<��]�u
��cJ̑~����M^P�<�&nM��ܠ���)0="e�E�<�OSo��ǋV�;Z�A��A�<��iIE|��:A�]�1�wh�|�<��9�r��� �-
�%�`^O�<���Jt��Z�oR53JXy�G�<�%F _���S6$�es,�@�<�ʂ!>D�떃��"��H���V�<��˞(V�;w��5fIq���~�<���6.�9[ ����a�łIs�<q�σ�%�������e��݋2�Wq�<�I��4�D���a>�`��r��l�<�� \G(��E��1pXӦG�r�<�FU$3m&z�I˩	�-�`�o�<aC� &4i&o�%S���áb�<����i�� k���<��$	g�<)2�K�~�U�KΜo3�@I�+�b�<�3�� c�ȷ����$=!��TJ�<��� $��q��gA�+��iz"��H�<	c4`帍!�
β_����wD�7�}{�n�����+�X����*[�Cl����n��\t�����.D��0n�S�����ʃ> ��3�.D���Q�1�4*D�jS0ݡ�-/D�P��S� ��T �"@�"�}p��-D�p�Q̉P�Xᔨʗ�>@ˑ�9D�����³:(����#+A\�T�7D��@#kS�n	P�;�,�5��l�5�5D�t�Ԏ�$a����a�ƕ�h�yS�>D��(�AA�m"� �8Z��A��*D��@"��8�8��w@8�J1K�+D�� �Q�,Ԋ��e��%�T�����"O.��W��?=��=���;$��T9�"OеC�KTK&L+��V	`�8���"O�)8��S�L򁐌Q��9�6"O���*�ؙv�^�q8L�RV"O��eL�=()v�cl�_��$"O|��ƇtaÄQ-�� �aQ!N�!�dϖ9m���ڋd��� �o�>|�!�Ă���(�Ҭ��)�`MQ�.Nf!�Kgzt0����������-��cQ!�d\�-� �Z�I�ɚ�"��!��5�L����>Zȶ	��aW�i�!�Z�� 0EK3��ݪ
H6Q�!�$��_�ܠ���|�R�K6�]&�!�ȫU&�Da�H�N峇���,`!�Ą�H�v�Ht��5��0�2�Z�t!��QR'L�$���FI�K!�ąu�$��R�����K���!��\�H�$R�	�P%���äs�!�����
`Μ&x�����'�!�_JP�ub��x��xa��>Kp!�$�T�uBBO� %��['g��m!�5\�l9B nq�V�G�<o!�DLX]�@#5���1�I��43�!�
;B{ب��M� ��p4�� a!��>*�Q�E�ݰ�V�����Xc!���+|a�c&���|x�D(4!�dT�7!"{�Ȕ37ڄ�z�$ԅL!�$�`J��y���8I�p��!�U'R�!�$H"&��Ip'_�k4b +q»Rc!�D�3UN��*��5*D(@䎴�!��PO����j�=�:��!BG�(v!��C�ldN4�wƙ/���;�y��&]Bm�������.�N裢J	$6J�3�΂"�y�o�<���B�!b�a��Ϯژ'`�Y�On8��P��C�$$�%��F�5��Cc3��hb� ��1�īߝi\4d�R��|)�
O��t�^�mgL�� ��0�����'��@C���lܓ@Tq�T`�T��c��S5Z��ȓKo�#R ��c$ΠPb�&`&0�'�F���e�S�O�z�Y�ςMٸx	 ��&|�zٲ
�'�`%#7o]2[�Q�玔3v��K�y�.T�u����7^� �!�L�2E�A�B�8]{�Bቯn��tI��44��f�0z���B�WH<i�jҵYh�#�f�4S������ _�<�b�I8��$9� �'�Xxf�W�<)�@1|������6"��u8-�g�<!�*F-]�H�ҫ-��@6�b�<YAf͗(ZxY�,)sF����ʕA�<��L�6u
 ���epbh��͏f�<q���+h3�������J��s5l`�<�m�,h��������$'X�<���M$g�"��ǎN%z�R�P��[�<)&D�N� U	gJ�&_ST((��M�<1`�͉&��`� �L�z\��f�Q�<��N�'
���REnP�$�v́��L�<��1�R=�$�^F(���O�<�!bX 9�,}kS�T�a�h�H�<aP��?QRdIT�Տ���yE-J�<A¡N28��sl[dxl���y�<��G� ��U욍0)���(�v�<�g�[�bo����LI�+�考u h�<�㏗.���AG d����B��b�<ٖ-ɽMDd����G<H��P�<�  ]k�
�ui�`�2O��	�L��"O��f��v���5���$Ţ"O��23�P�p��%���K.%�L@"O��P���;�R�vbF(݈\�"O���ƫ�:R�h�PBH�5X\U:�"Oິ���3�΄��lƘZ�h�"O. �S����mXrL*y�&	X"O�LJ��+��;�L�43�~�� "O|@@�(J�d}�17JY7C�@X"OR���ϕj�~8X£
k�b	3�"ObhpC	@V��	DD>��b�"Oܴ�I��D��"�U��A�"O��S0�7�E
����@���ȓY ����M��/p@=�сE$:V�݅�u0!��h�L��7�ҢB6��ȓ=G� A� ���$��'_9��J� �1"� y$��C�+P'|�*�ȓX�eQ`�>pn���� �@��T�ȓ8��hpĒ7 }�y�D�F0@����/x�]0���<<��JƂÖT��d�ȓf�䬸b 	|��M�@�M�3$�͆ȓ:��`!�+R [�d�p�+�\.݆ȓ7\�a��+Z
mKډ��HN�sQ����;�&y�W�"�N��F�H,Zڶ����%�%�B�9[ �� �ϩgxTمȓ޼�[@���b����S��` �مȓlL�v�A�2���Ď�=���ȓpY�9����="��������Ԅ�|��� 8b�6����{�����P�a��J�[}����/)�b̈́�Z4V)9�̖k�e�qc�Ӥd�ȓ@=22�иK��e��/Fg��Y�ȓ�V�`I$(�:����<0�y�ȓM��,Cf�}rP`���I>v/����zI#��آ�i�e$s���<�u�r��b�״�h�\t��� �ȼ�����Ƙ��"O��p	W�LC��H�d�9a*�;eH� �v	�$K�?��R�BS���'��!��; G�!��.�����'�d0P�߭*8A��	 8]hU��&�͊��9�r�c�E�����H�����1$�<ul���*-O,8�VOǎ#�t�3��Wm�\y�/�C��B�OCB�����̟�]k B�I?]�\!�JU��a%� >�ʓU�ZR$UZ� ����׽"S��Bu� ���m�H��E��#�:���m �B�ɿ�tu�v��P��(���*F���3�׆i�P+�i�(�JI)�$���'.����ż42������M��X���*԰]��ҙ-��HD��`O��BÎT �څ�"N%B�Q9�$��6�@	2�=O�ě�͔�4����%�F�t
��	��D9bC�
�X�Z �I%��ܳ�ˇ� X���q���Ga�]�pȐO�}ۅ�U~�>t�0�ȑ(���6?O^}��k	��<�-n��Y�!�}�6x��(���5�v�#��ʷqd=�$aU� �!���.J����Iǟ g�ӣ�H*?����ʞI�f�!`���?������?��#`a|z5�'���a�IԿ�B�����P� %"	�n�����̪HH�_
@�����&A�n��3$��X� �<j�`p:��F���O�����^��\y'HM�r�3��I����R���.���`�[�u��9RaK�
z�0��H�l�<E2a�����ৌC����f�R�I����o�)T1��uKy�|��ؼr�6��CX�V����֎�M���3�Bi�S4U
$T�S���1�B���Oٛ`�tC�ɚ�p��W�#��xyf�Y�`���Q�ƻH1d)c���f���[�(F��,�B�/O�L""ҫ[y��a�K�+�έY�'�м"F�Ҩ��dꍤ-̎�Z0����$3�A��J��t�l�� �]#��M�rџ����֮%��d蕄D�����4�{��Ť���� �"N>]2��g,$�&���@��w�}���ٻS2�0p�����?�֠��
��Xs��R��j"$��<��A�6��hb)ϩ Oh��.��h#�J���a��ղ��Hw���to�"p�<���S�? H1�@�(0Fp���iz�f�
��R���J���k��S 
�2EM�CyB�Q̬�⥈�%�$D�B��0?)FAA�@�ޔ�$��>���!AFEڶС�+<L[<	0P#ɽp�ԍ��x�T�ˌ�$�#t���PE�zp��0f�7%���jTN����O�D�6�^(D0����T.QX��jO	}���� ��J�����=�����+��0���Ad�3:��rOI���!�d׃��!��!�?*��&?�`'J��N�@�nƷ-��K 	2D��`�IX�]�.X��m�p�b"DB��Ř�zwB���G�%E��O��@��O~R�.e���Kۇ�v�ڷh���p?Q���=*�vh��� "`d#%�A�]�E����60P↷QU\�a��,ܼ���X�2�8d��>e�}1�f¼m6�����A�RY�1��K�6�u�1�ElU��kVFKW��`C�"r���v�Hx(<9B�\&`p�#�X�6W<]s�qy�i�b��H�$�.m���U������~�`&V�
p3�gЦN4���bp�<�VcŨ������rup�z����Å)��#O�rwt�b�&r�'��r�B�(�-I|H��)I/h��U��d�۷���
|(%f�Z� e�d0|hr�H�@�Pa`d��-2LO,2h��_���;@E�)Y��X��'�PY�W�J�R�t�� � EA�3!f 5V��
oAx�H�+�!�d�;#%dR�!�+e㔉�c����1O���C��碵;Bb&ڧC��ä� =����c�]�>T��ڎ)����4:��D�C��8����B�3!8m'�9k�H&u�Ć�<@������ �`��7� ����ȓp�N��ҧCW��h�ЋT�=��d�������-l���vB�y)L	��9f����	.t���b[4$2E�ȓ>s����!�� �э.\��ȓ&�X�#�ۥN�>|�DK�����ȓi�=��(��+r���t��Җ��ȓG���/�0�U2 ���B��'a6����P:�L����X���!z�!�CM����$͢\�V�3�n�!�d�sz4��Rꌳf�0��&��	W�����'#��=��>I�B��;���⬌*_/�!�i=D��b��^�-��Da5�H�:�����9D�)V�0�v�qB�2:��� 9D�,D`��a��� 	�(C��r�. D�ز�\xW�J���:!� �!D��选� P(�'��al�d�?D��9��d�ڬ��ոr�h@�0D��z��tV6�l+L/x2�q�0D����] (vU�g#��K��z�;D�t*��=�څ�"�8L���/%D��s1�@&I�0�áEʰBh�\��?D�Lyfe�2x����I%+/p}���!D�j���=��Q�bA6(m
�-?D�����.8�R��׬S���צ>D��+A����P��2 �)D���r
����i"T�X�:���1w�'D���dI%)���$����5�cO%D�|;�A�>\�������e�A��!"D�P���L�2q��(]�x����V�"D� 8UhBY-X��F�d+T�#��%D�8�a8^ y�A�q><��@"T����hJ���2#��>���"OXy��\�1��
ŨQ������"O��1a�MJg��3�ǘ�c�x�4"O݀%�ۜ"M������c6���"O����E�1�"�I����A�@�1�"O�Ւ�d̻����w�WE�8="4"O�e��gߚAjr�`w��a�Ȥ"O�
�(T�
�I���+2J�0e"O�q0k�<my T��+-d�գ�"O� �۷&�	`1;��F�	��	e"O�%:q��T�|�5ዩ �X��"O��a�n��h4�ŏ�(S8t�j�"OX�#bT.�p��m��l-� @"O�1b���3�����mK�6B��`"OV8Z�I�04	���6\�X�Ԭ�1"O��A�jR�6�M@g�w� ��"O�̠��~UR��vl[�)�$z�"O��!a�A�/>1P+X��HI��"Ox�����(�к��V)�䡩v"Or���O�K�NaB0g�$<���j�"ODe�!��3l�,�ڃ��<\V��kt"Oz|��[#~A��P�X���"O̅�pj �z�0@T�L�*�"O�0�Ŕ��~�"
Z����٧"Oj<A�:8$m���M-.�t!�"OʴpD�
�o�.�� �4���"O|�%N���-",��%�❂"Of��C$[�c+>�pu��E��,�"O^� ��Ԭ\P���7
�9�Lц"O�Y۶G%�*yaG+�	pPP�h�"OT!ƁQ:)�I@dI'r0��h�"O�lx�g_�p��c��43:,3g"O4��
7L� ��f`�:�!!3"O�Dk��N*m��qrO�4`N�iڵ"O��U΂�r��U�#.%U*���"O8��d��)����C��a�"O�	Ht�׶|f����N�^VH��"O�g ��P�0Q
�NR�L3f���"O.8��O^>�ҴP4G�,7�q2"O�Hb��DP6�Ӷ�D6S�2��"O�� �-"��A[�&焅9e"O�8��A�6V,��0�5>�H]��"OZu��a?.�v�:�BO7�6�"O��RrI���x( �dьUc"O�%Pc��.
���"��F>;��	A"O� �R��� �m��VNmH�"OB��0G�"&�l	�*�2zGt$"O�B��S���+���i7"O^�p�D�HJy	�ʰI$���A"O����&�� ���J�dU.X/8U�2"O�h*��4m#=���-[�}��"OjŰ�
��	�#�	q�U�"O6�25�U?_�v��sV~����"O e���.��cB��7p0@ɐ"OHe
�� �5Ж��),Zm@"O|�s��a:��K�a8���"O�̰��E�K���p��.w�~ĩq"O�=�j�4��Yb�
����"O伂�B�7Rc�ĳu�U)Aj`|�u"O`qB��wM�:G�Z3�"O��#���Jx��Q:D8R�8�$�h�<��'��1b 0,��`�/WM�<q�_�EDr�Q�
�g�<a��D�<a�)W7}�Ա�F��0n��B*A�<Q���+iTu@f/S��Rl��D�x�<����*<��ۗ�ůDd�,��-w�<��%E>
�`o�%#�z�I���t�<Y���`k�\�l�qRz�WMY_�<���N��+��+Vi
�(P~�<�ҼB�*i�L�2"�	�q�<!2�H�jȑq�I\�S!��qNEP�<���8�QQX�J�93��P�<���ٛ92ZP�Ү�nm��AEh�H�<� �%;2Ń�+�ntb�
I�5T4�D"OЭ*0��}KXU��Q
)��"O&�FB�
�b�
Ʀ�T��`�"O.���R&�̐��@)Р��"O�|�pM�sI��q���4�؄��"Of�5�*�(��
��-�"Om���C�([��K#�^�>��F"O��$ۉ�\\�E ��\�R�"OP��F]4F��v�5/��E�"O踳ÀC��p�#��2 ���g"Oz ���l��:���P�jm9B"O��q�ɯ>����r@�ku8�8�"O�$�#��aj��#HA�p��"O�����~ʘ5���޷*�Μ��"O�e0�C���ã�
L� (��"O�5��'�=82Z�T�T"���"O�y��ɗ	��SD� +n���"O8A�$�0rFh�'�T���"O�"��ڑF@�i�@�(w�Z�ّ"O�(�d�<Z��L`!��t��;�"ORpAv�ö����M61��3�"O����&�Q7�\��ɀ �N�j�"O��(�1�R����qƶ�R!"OHr5�)G[b�0����n��r"O��[SAQ�}S����\>:[� "OH���L�Q�(0P� �o$:���"O^U ���3G1�ȡsn��b�.��S"O����T����$���*�"O>E	p$V�?�y��߶Tz\��d"Oh�Y1�ؘyP�IYC��8j��Q�"O�]{4�V�?@�l �ϕ�[��X�"O
�8f���+<��g��Kx�CD"O0"gnJ:(�tX�d�wߢq�A"O�,y��D$-�(b�F:r�%J"O�%B�*� �bls���Hj�"O�9R*W�!�^-+���e$Y�"O �ʀ�C>��4�5�ä<�Q˔"O5S���{�jR����R��"O��C썠i��( RC��a}�A��"O�Dz0T�s@���5"UB���"O�`���8'�H��!�Q�l��"O|�3���0���8vO�<f&�5��"O�:���'{�:�J�LR�a�95"O�ɩ@��:e�� �
�	'����"O
��qgˍs���i��ϨC2"OTx�%Й#�������q"O�r&FS3>�b���*W��`-�yr�f�:����S��]��lA �yrDʍ0Ϫ�3�c�x2|�UI�8�yR�Yt`a�ń0x�يm���y"d�$CdTm��cO+��A��CR��yb�E�`��%�:)�� 򔫍��yIِ�8�!ǸV��$⣀_�yr�5\anm��ė�bh�f���y���Q-��r����2X
�F�;�yR���p�]is	���܉j'��=�yٳ8'���K��(���+S��y��8/�L{DC�-=:.�6�yB��2� ���#�� �F�ڤbϋ�yB�K�b���3�jV��|����>�y��PT��!p# LO�^��#� �y��v���.LE�l9��A��yBɔ�RE�UoՔ*� �u�^��yR��4�E��/�@%q�S��y
� ��0͘�ls�$HW��$X��0��"O�D�����Kl�E9���;X~0� b"O�Se��a�r�`gI
=k�0q�"O�8���	ژ���gH�[m~@C�"O��z⌛,�PS�FR�rt�u��"O���	�d/�L�!BOֶ�"O<�V
�L��tk޾H����"O4��V Ë?��,����(W�B}s"O�M+ J}�(�Su!QU|e�"O���4���/�:1���H/X0��"O�Ȑ��7��t��	�o8~D� "O��z*�W[4Y�(6�p"O���¸er�,��>����"OlH:e]������\�*����"O�hS3 W�@# ��:�&"O�	��\�uNEP�C�2��5"O����FL&p��H��L�5�V1��"O���'�>�pt���F�Z��#"O�\r������*Ԧ8�v�7"Oz�ˑ�(���ϼ�MP"O�(G�ڜz�]*�O�R��12�"O�(*$��'s��5���+h�"O���*����A���x,�0"O���S��0�!��T�P��g"O�ڂD�P���5�1x����"O�����>������V��5+�"O�� ��/�*E	��͝X���
�"Ob�h#�קN�^usfo���}��"O�t����PО�ì��)�j��`"O(�X�d�6�iT���T�Cv"O�\���#�.�1�R�s����"O���B�2i�8K��!~v2��A"O���$KE�j�p�D�(+`�0"O4� «,a�b��qh0S"O�LX��ƐԶ)x�ػUwd9D"O��ya�S�vO&!ס�;Ħ��S"O��U#�:HӴ\���	j�"OJ��$�J�XI�����96�6[�"ON`��^�)0���GIA��0E�"O�ā��.��%sc�;q�8�4"O }�lL)O �`±cE �����"OƑ��K:_�zISl�5H�٠ "O�5"bt<y��	�)\{�A+�"O~�
�'5��Ъ���$.,9�"OJ-��X
�� *V��j�X{"OR��!ɰa�ujH�K����f"O��('Mܪu'�-���0�����"O�h j�*	��]��ΐI� ��"O�I���4�L�E���Q�j��E"O� �r���o��	���]!O
 �Y�"Oнh2bPKLJ���o��A��k�"O�A��mV�s%�@� btnd{p"O��� ('��}�.P�Zhhy�"On��6�^;5�8���CPF6��"O�Qk@G� A>���ĂRK~�#�"O����Q�*)�l;bl�t2��2&"O�
r���&r$!GMK572���W"O��PaU(Y�$5r���j��	�"O��S)9qm�DI�5'��L"O���aMЙ^�v�����
c�p�r"Oa#���#�p=rvBŔs��<�"O4�qqDڌI?|�� �Da��9�ҘH���#�P�h��I3�(��$�����ce$��Y[��2��-W�����Gx��TÜ
��S6�
�9"J��cJ���$�2�(O�>� ȱ��̃�e�a�p+��Q�jx���i�}Dy���W&n���
M�^h��r x�<)�O=<���Nļk�^l�u�Q���H��}B�e���'3��=����&}��S�Q�vVVy'�t�%�)��":r@�D��,�<���K<��J7d�<E��'�DhE��Ο�]�(���e�"�MS�(�S�OD�ms(��7E���@�a����S�	��0|����B�r����h�f�:�H	X�h�d�2��O��I	B[�q��
&���8�L�056�O���a�,akn�!QHK�.\%���	�_����-"�D�#@_�,Ȝ扏I��$jq��S��"�e�2St�y��+''�@��Iv
�.?NbYp��DP��}�'{���#Q��jlyj���a�T����	e>�Ѐ"Ȏ`��`�"Ň�)Ծ����0�I5o�Q�������7JRN8�e	�eǂ��6�xb �R���	����2���U�`ʇ�S�zr���U��>a�&3�S�OD���əd�HaydڈҎ��ٴq�<�<E�4g��	̲֔�� Ff�����rQ��b	�'��E�@-%̝��ဳ7��!�>1��-�S�S }z���d��)'�����7_f�OL�������d*x�h�@D�w��"fĴxd�	�#Q�"}�ダN[Z�Y#��m�:py���Ц��I+�S�O:	d�Mx:���B$�$���'G���3��_��Pб倊2�|�	�'i�q��ެkz� �f�ɟ*�5��'��Mr��1άx��
���fC䉩}'��#c��75p��ܔ6UB�I�9j��jB�TQ�Ʈ�%}�C�IJJ��" ,ޛj�����܎1M~C䉔M/��!��en�Q����7��B䉽.�f(�i�� f�1ϔ��\C��:%���,9U�l�0ā�1n? C�	�4�����OӒ&������4O�DC�I���]���FH|R�D;5�pB�I�5�J �P&^����F ;�C�
Y8�h����5���"��)V �B�I�!h�hy��]� ŀE��H�fݪB�ɦi�l�`"��hxE��ޠ�TB�z�5���0P�ȤG	��C�I�6������e2���ؤp�C�Ʌc 0��e�4z���Kw�՚ڠC�I5PJ@��mR�d����9JXC�	�o)�))�NN X�`@ �-�PC�	�8u��H�T?Z���Фn��C�ɞqT�<�V(͓r�^�xU*O2	R�C�I;F�<q�en�5 @h�#2��C䉗b���;I��VzPq��M�|C�əJZ�����|�T��d͆�fC�	=Z�!�q�_&.xj�hʀR0C�I#��Y�ecڰyXr�((2RB�I<�f!��X�.֍؁�V�BHB�	+S�nhQW�9�! ��'oFB�#L�-B�
5i��a�JS%cA���@�L�[3���H�ٺ���*j !�d��i��I��恪,��I�IA�!���I���B��S�!�%��<x!�_�
�Y�BnΈa�e;�eS�+m!��{���ArJʐ)R�f�a!�$�mn�k�%5���^9�!�dP�# ��tn��I���I�!�$��r��-�V��k]��"�֙�!��8.�楹��B�1Z�|�H�4-�!�DPzN��kA��%k���ǡ׽g!�$ձd��K@�Z6D:D��r`kZ!�Ą2�9��O\�3rȡ�fE!�� ��E�e$�a��^:��ҵ"O\U��F�Y~�PO�#�
U�"O�0j��A:���1O��}C%"O�����
 m�AME��"	�"O�iqSaũq�@U���)x,�3�"O��6�P�.ABQbդ��|P�+"O�(҆_�Ъ�c��I�V"OT��6�1oy��ȌL�(��P"O��J��\�2k�MySВY�J쒧"O���'{f���M�7��@1�"O��;�� 9��Y�>�8E"O�	�`%�
[o����Vr��h"O>���ΓA��P�b�Rp0"O`�d!E[��+�E� 	��"OtP���t	��JE�P!yޘ��`"O�Ҧ�ڀС`� �5��舑"O���D�A"pU�`*�_Z����"O��E�b.�܈O�7<��@P0"Ol}��&��I�2��у0��� "O��c^�E E��SRh{���y���P�رRǆH�
U0`���?�yX28-HlpA���*�#���yb��.0}&�^�J"d8�J>�y"�_�\ �% BU���
����y2!��L2��`�\�ZQ0ԅ�kW$T�QJWC/��8w��qҌa�ȓ5��+�*Ј]����b_�hԚ�ȓ6/R;dB�]�zH)�,384B�I�v���0�"�>jV����G�"B�I�a����/S~rħV�B~8B䉸(~�u����)c� �Oc6tC��.k���ф�+h�:�{�*C�ywJC�	�`D 4s�(V�	�L�b"O��J�f��Av��f�I*:��|��"O6}�!����ȱ����9!ft=@R"O���/�<g���Ui�+a�4�"O�(�5jǂ^w>�2��)5J&4C�"O��{w�B3.Ȣ7�Ša��	��"O���TIٸ���!�,��V��"O"*N��N�A�!N�m��C�"O�y ���_��y�`@�%xc�"O}��̌,� �鄀ۄ+�dE�V"O�X��0�L��.�9��1��"O��@ ��M.�1��n�S����"O@ �� 4�ƴ�� E�bP��"O�ah�@�$o��ԫ��1��ij"Oz�a1"δ���
�ʜ��U2�"O�;���(�αS$iФF�.H�e"O��i�]�h�!��*J�d��p�c"O\@9������HKZ P�Bp�"O�� ' �����S+o��`"O} ��	%��d V���0}n@�3"O��C�C;HA��N+w�VQ��"O"l"�.�a6���5�L���Ԁ�"Ol���o�L]Jx`
��E��ؚ�"OxS��<J�-���ձ�l�hv"O�Ą���[E�L�"OPir�%�_��e�Q�CaP	��"O^P#q�|�r(Z�ˇ#l	rX� "ODqc�x�6���Z��4[�"O���ϔz3r[EG�[�P"O�7iJ�no�fj���.��"Ot�D�Ja�1�ө��5_ A�"O,\�@'=�����׭PD��bC"O� |Y���	]j���F�)b���"O�<�W��T����"zQ��؇"O$<j�/��]x���A�I
s"O.���Z��4˵C�;�BE��"O��r(��|-�F�èe��$ �"O�P����8����O̹�B 0"O�}��BŠ}v��8d��tB���"Of�A咝0tr�P�ְQnD(v"O�5	�O�D'ݣ6A�La*(Y�"O�9��@ (%������&Z@��"O�d�1����gڤudʵ4"O�4{���<Kv99v�фaSV���"O��Cv��)mEJ;o"H�z\��"O��Xe:f8���;]^�IS��N�<A�=>,<�2��C^���UN�<�chѨ-⨡Jce\�N����fW~�<��K�\���n�?�����y�<�dh��5b��F�Z�[v��	�w�<��!J3M[ h*wcaD%>� ��d�@�	�3^w�L��˝;��H����|8�,;V��]� �� 0̕��X�����IA��(;�#R�z⨇�$F~�[U��!2�4y��ИMd�@��1sv��Q��0W�v�@6fļQY�Նȓf�R%P..�b�v$۸F\���ȓVx ���a9H�Y���\x�]�ȓd��P����~�P bТp.q��``�B-�]��r7(��s����ȓ8�0���ݵV�J,�2
>$�Y�'��~�
K<LY� ��W	�x���O��y�M� >M�%�w_0ղEe��y2�b\�f.F2N�E����m��C�	�b"�}��ឍp��$��ή.7B�ɴ/�Z,��Ȣ��0x���<HB�	�C�8�@=-.d����Z�qe6B�I7�@|��cW�nq`dc&�����B��/u�����$0�.N�lA���[�<i�☒w;�}@4 �z�>8�Qd�[�<��G� ��ܑ%�;&����eW�<٧�� h��CWEm�r��C�S�<ٓˉo�Ly�Vn� �5Ȇj�i�<1�>]% �PO
�u�2U��A�d�<)����&c
�2摀��k "�d�<!�c�?�� % =�:<�g�{�<�u�Vv��R�E�Zv�����Q�<I��K�c���J��٢Akz���*VL�<���үJ7�Q�c
�w$b�����F�<���Q��R3B��*g0`����l�<A�FI�~�")��f��I;��$�Hi�<	��)CbI��O��U��Y���d�<�b吧� @S��i9�};�Qi�<yW�dt����C�x��Ass
�g�<�c��M�L+�!_9�ys��c�<a-��IX�8���=&�qc�
�c�<�tj=k�ĕ�w�D�<��fC�b�<�&k L�0ԀS�ӽq60��vBMT�<i��N�h��hQ���K>Ś'M�v�<a���
4��z��\32[ Pd(FW�<�V�J��L`����s���U�O�<��D�`��	��pڲ` �Yc�<��
Wސ�Y%B�7[V�Г��y�<� FZ!	�goM�:�����\q�<р�^�'��h�)8��zЍd�<ٱ�D�R�X[F[,da庑��]�<� �SV#�"�*��փ4��b"O
�����|�dEj���H.�DpV"O�E+��D�FR��Qh��\/�xd"O�@���K�(��0IR%�+h|J�"O24#���(g��  �=�L�p"O�dh�(*�re�\>k��"O��&�)�(�B��I�"O�%zV ��4���B�*H����C"O��1s�G�x�<s��Š�$I�d"O&UivE�8����"��T檬�"O~�B�����jݺ�p'"OV��r�b��-�f*�=�p�"O�$ V�̩�r��cD�[�PMj�"O$������l�X�BQ�{��4�'"Ov}3��;i��x��{u���"Ob P��m0ܘ���C�8N�9�"O�V՟�^��5�1y�PͰ�"O􅠇A�������1��"1"O���1�9st���%��"O�	j֍S�Tr��,�2�Yy�"Od�ńG8_ȴ��	~�y+�"O�0��H�
P�V��V�]�P<�3"OH�K��U�K�����l� �H(�"O�P3d�51D������ I��Q"O~�sΐ�[�1��A�0=���"O��5�K"5&�:��5`���"Ot��Ĩ	4p�X����h�tU��"O����   ��   d  �  �#  0.  V8  C  �N  {W  �]  4d  �k  �t  �{  ׁ  �  ]�  ��  ��  <�  �  ��  �  F�  ��  ��  �  T�  ��  ��  �  [�  ��  �  ��  �  ^ � f! �' �- �6 �< D �J �P W �^  `� u�	����ZviC�'lj\�0�Iz+��D��g�2T@���O�6�M���lc"�¥�V���E�q\I����:&p�\C�
4��ӛgή�#�_
�@�Xw_����O�N�r�O)<4`�MƐHhXi"!j|����CmX�|�|К1�],dD^��Ǐ�.3�qs�nݽ�Ն]�?�r۴p�z���J�����7Xúy�I�\��б�'���xRB�.8e��2��iӚ2@<ON���O����OB����m3�-A�M8��D���O ��ح$L�oXyB�'����f�Oar�'��i��G
T��� C��0�y`�'��'���'u��'<�\wK��p���j�eh��HtԆؓ���/?�64�JL.�	\�D�(Q�P� ��\{l(bo��<G��5�T���'��5�d��<��٨/+��RD>���1���Z�K͹y����*�?a��?���?����?q���i��#G� �K��@k�F�#V�ZHKu��O~�oZ �M�u�i��7��O<�oھp��<)�4;�@X�3앝w0$|�VM߼v{ʥ�耓+�8Q��iU6M�O@��{"�?+�H~\@ @�@���z4��	˱;��p =jX[��O@o���MC����T�OP�kgV�:rP1=dqЇ�s��7��
zJ� �tG=j�v�I�5�.�t�F szTlZ7�M�½i��xX׀N}
�/\�u:���u�$s�Zy��QvT�7MTڦ��۴^�E
��;�`�S���kt�� �2vA��s�ʹQ ��YQ ��&���2;�ypR�i�6m�Ԧ)���[�"h�(��������_6��$�]2f ��lN̜��4l�R�F��R�j�!�i͚E��L�����'��!�\�`������N�Y1�'�ON���O���ۦ%�O�"�J���a����7�9"�(�Z����O��D�OTY@p��^L���6!
�r��͛�xl@���(N����D�.ͦ��Ԁ�F�Q�dH��(�ѳ�@H�.�(��GT<{&�y����:^Ed�C"i��BKJQ�t��=uQ���S'�<rY�Hq�`�*	�p�{ዖ�\�������OB���O&�O:���O^˓�?�TNB�6��IpJ�H��Y�iF�?��q.^���������|ڦ�'���x��Q�s/��/��
���D�d!�0oß��j�w^V9�b
Z�x����?$������?)��ʡ�&aB#L�6H2V� 3IGi�� � id�$�Ou�
�B I�]v��c��4{��	�-�"�a��:]��9Ȱ��=\}Ƚ�M�V�' �� TЩ?p�9��	�+N��'z�8��rT�)%�'��� ��Y^"h��m��ؤ
� ���?Q���?�����Z��]qA��n��c'K<h{ў����M�G�i��'�=�։��dJ��x���
4%.\�W�q� �D�<Q�J�������?�����S���L ��Yq��Q�CI  $kpi��P;:�@T��8�"�A2�|z��mF<�+�DC?A�[6A1f4S�P�X\ 4K�,.,Z�:'��>
}3��7@��`�|WÏ�t��	�q�h��#�;����Ԩ�&7d�n���\�F���O��3����p؊���M�Ţ�
H�ۢ��$�S�O8����+�:u���2�h[�j#���'�R�mӘ�oZJ�i>5�my��[��� ke�àP��� ,s��}�ah�>���?Q,O�˧���I�u���g��Z2&��T��2I 4�:;-^-��eb@����"M*{��Fy���<沽�0���@� �6�L0d퐐��NX8>��JG�
Z� �2�	I!a�Z=FyR�գ(���%ȝ�W'��!��Z6������V�0ғ��'����M�>cs8]9`o����@�'���'�ў��<��L��	sp���	b�
��j�ɶ�M�Ƶi&�	�x���4�?�'����@�/jRN,@fB]�_�:�������O|��v>�m�8jn@�,y���!V j�<]�N�~_l��A�3=t����ߨ,N<�<��J)� ���ػ
d4!æ�ҵO���q`�:4�̓Faט3F�`�G��(n�	� �]���o���I�M�ļi��j��O.�ƅÁ �@���J?g��٦������?�}��\w�>9{���p�d��Lr�����?A*��Io�*��eB3��
A2�p$�иd��jٴ�?Qӹit��)�tM��	AY������M���J|�q��/`>$b�h�*.��9���?�����4���a��a|4��ɓ�\P��>��Gn�4^ ��`d��7�y'�^~2��O��x�dD�	�=�7-(tF,�@d� OX���O{���Չ�Bx%R��2Ce����O�4J��'��6�Wq�S^̧QG�a�r� �A�Z�a���4�$�P��^�I����Wy�	w�����#�,�1 �
�N�#?�$�')�v�'�6��OJ�Kf���1p��@VяUo6��G\�����fyB������'���'�	��5�7"Y�<�. �#)׮-�"	
(�MJJQ��H�=-�h���m�x�D�O�~��vm��~�2(��M�f��B�^�0��ƃ]d�)�Q/�-I,�I�jV	<�E&�(��S+mK>, 3F��AR� �"5�4��&n�
Q�$�r�q���'�P�:��٘�?���?�bh҅k��� ~,cAr�z!J��|�)�S{<6ujd��|w��*ׅ#����O�@o��M�M>��'��/Otģ�%�8�H#�"��@�@]
�oџ�	��'I�S�|r1��C���2Nя	)� �0Q��Mzw�[1I�Tɑ�
��8�V�:�j�9C�d�<9V
(Ah�{e��`h�#ѧ��~�8�� ��Z�����% x�B�aL>a�I
�����<b�y:���w���K�I#D�,r�ڟxb�4葞�Dx��Ҭ~�TE3�O��jЌ�yd�B��?qO>���?�/O��O�a��9^�Fxi��R-U,�� �O2�oȟx�ܴH�F]>툵�	'�M����?Y�^Ĵ9��l��w��I��L��?a�>.Jm���?ٞO�r� $َF��m���YHH`�� �iWέ.�r������=_p��땶A�2`���Dɮ ��5�cj�;��7-٨A�(Ȫ��� @�ѫ�$#kW���
�,*���3�& ,�O��3�'D2���Y"��^Z�tj�2*��x3pe4���O���Dv��$���Q�`g-&��O�=ͧ6-r! �'!3�*ܚ3�L��1nc����$ۧ!�|�D�OL�d�|�2$�+�?��)9<բ'��1����` �?��r�X�
$8Р!Y�$�3
^<�t��by�ȟ����H��8�����%\+@(Ӳ��Њ@oR}��Q'�S�,����E@^ �=�gmR3*�����KK�8#�0gW5v70�rF�I⟨F��9OLu��F�>,~D���A�5R��af"OZ�2��,,f�E�qf<3.8y��۟�8��dق*�IS���VzU��++�(lZ��T�'����C�O�B�'�R^��#����7�D9��`�I j��Q8���L�-� ��C%bܢ4�O��
?���O?�E$�'y�4*b��
+�p���l*�9	�AI�#~`	SE��V0(����%-�2cB6�hdY�K�U�K��q|�H�B�fӾ<�'uȈ����Ο�'��j�V�~�d��SK�V���'�"]�(�IA�'��$RA���S!L����(g���R���'�B7�Oզ�����M�-�>��|
�d��u��P�3���l�* ��&vn�r��D��?q���?��5����O<�dg>��rm��3�\�R��`5g-�qF^K�)�55�HۓJfڡBa꛵kJ�)K�nMP	�l�U(U�#��劥ӪC�a{d�?Oq&t�s���3�f�Y���)	>D���?����*e�*�	�f|��YD�(��|��/A��X�/,7âe �	�&=�h�$���ڴ�?Q)O*��7K�W�g�R���˖�<a�!��1 ���<���?���*0�f�B[�:S0�$mHl�J��K�ò��A�aS���� ������F�'������V5T��Qa4�L���F�l(��Rf�hP躲��.|h��R`�-*��u�|" 0�?�������;:Bt]�f�+`�6�T8V��J>Y���0=�)'u��+�!lu"3ʄM���hO�)�A"�߾d�$Ls��:|$)@�	�ON�E8�l ��i��O�����p�ډp����qƇ�D�a��j���4��K$�T>s�F����B�@A����=p�H�#b5#�*�D�L�SB��]��H�O=C��@^~�RRL6Vj�an�0cJ��5$�-%�������2�mT�1p������	���)5c��$���){��iq>iyb��7��l{ө��e��@ׅ0�	p���S29FJAjCC}���v&L��=A�-���o`��OJ�̛ۗ�Τ��1l�
eaE���}�I�h�ɬ ��iȒ����	̟���ݼ�&FG�r�
��Kȇ=r\��->�"�xl�P�u#��9;���Y�c>���T�*��"q��u��eِ34q�P�w�R��R=6X!R�U�؆� u�I�<1�Tiq�'���:fn�o���:�e�WCb�2�������B�'�ў3���,@��iqpK�?u��!��R�<I��=мzPfC�w�Fc!b	Gy>��|����KChɫ����;'D�1%	h�@v&��[7<���O����Oj���O��v>a5�۽p��!@��G�$�#`a--�*�7/�tI5G��%c�D�A,�G�Q� ���T�,��w�Ӛs�d��B2H#�`B�*ߛX�(�Y�	�+�°�'�E�c��m��I�B�=b��ݛ4G߬c�.Iӷ�IA�T!� �O���4ړ�O��T�U�*�q@d�70�%�'�'B1Ob�*�CԖK��<2��R �x낚|$mӀ��<�p�'"h���'��ݕf�ܚ���9vQL��7�2�'�
��'�b9��`�#(K�`4�ZaJ���V���@Y�8
 �ִAw:��C흩SZ@�?q��1[�Faطd(@Ȅ�G�
pD\
R�ȮO��)Fmȸ13��e�'FB����'�*PsR�;�����{s��0
�'���Y��[�ve�8��O4��<k	�iIR�`��ѣ ��*"�bӷDM���y��ۣ�i,��']哥u���I�erQT�X�|�@�KI61��5�	ȟ� �NِC���"`3	�9iW	��j�y	�v�t���U�&�����H��i&��$^��E�Y����v��1�M�g�>3z(��O?	�֦	�@.��Hg�_5^���ôh3?��Θ����Ij�O��[?;.���"�V(�۷�ħ�!��$J4m����8���i7��j�џ�+��I4�lpY�O �\�x�gA
kV�6-�O��D�O�%�ڬ;e����O>���O�睑K�
��$��Da�iJ��@�6T��E�7��D��o��Q��d� z�d0a���Kn�K�Z�ڈȕ�K6��y�F��2�\�$��+Fnʓ7f�"��8����]�����l~R��;�?����hO�����8� �EO+^
l�+�=D�4�!�4	�$+Ύ;X�x�O�<ad�i>��IMybk"JJ�ܪlV�VH�Q;w��>�6ዧ�P6,���'j��'��������|B�iP(~>�y;��[]�r�3�,��|��0��CV� �Ih&,Ӯ4����HR��<Õw�? M{�؆8f<�"!o�)K�L@���� ~�Uar��0��QI	_��z�gԎ	ғO��z�焘@㢍��cB*�M�Ѣ̛F5��'�b�d>�'=�Д�B��Dܙ;�'0?��P��	x̓,mTU�!��<Ri�x��(�e���%��;ڴ�?�+O�E�p��Ѧ5�	ԟ)ҨΪ!rz}�� <%�L��b̟��ɴ8���ΟH��*�����$��}�1Ѝ����M�$'D�rB�X��(�H���7H5ބ ��9ʓ0%r[���/����E��q\8��tk�7.&�!��
��ĉ������iB]Q%�|�C̄�?�`�ip�ɢUf<yi�E�)?�,�	��Q?(�O�?�# `?	w#ݮ6?B�[pJm��u�}��hO�iA���+RN��XZ���%�~�:�vL�O�4sb>O̉����!�I����O�܄R��'ݰ�qGL�-N���s�a��S��H��'�b&Q}��:d��E�r`8����t�Tez�FF�d��SpC��G�OI��g��>D�n�'�J����N�lIa@�M�]�~4y�O�n�]z\GY���M�,�S'�U�NP"�Ȇ*F#����� N�)§HQty��$}�ő�ߵVF�ą�M�4��!�,+����� ��G{"�'C�#=�,�v��%���n�AЏ&ț��'�2�'u��h���2�']R�'��N�?�$@ShׄO���#�?}�(����Ol}")��+v"i���y,����58�
_�M氘��a��c�>���ZP��|�<a��+�>}¦f�`�RM`��ݟ(�'�x����?��+A�nP��OY#Tnv�2p&�Y�`B�	�):2�#�Ԕ[v���C���˓,������'k��3��}�J�Ue��U�d7�� l�7��O����O�˓��b>��b�.���P�R�2�x�YEI��y�@�sH�=?U��c���`���$���Q�H"s��Mh��u�Sm�d�ဌ�k�JM��&?TGd�s����*���K؄zR!2�d�{JQ�f�oKB���Ֆz,��e��O&$m�HO�"<	����u"|�(�mҦhapH���Ig���񑁞�E�h��N6��%����4vg��]�$�b����Mk���?�c%�+|���v
�{�ڕQF�4�?A��iG�����?�O�H(�B\�J�����.1�hs�oXMdh�Q'�չ{���Y�/ԡ�ZAp�`�B�'^p�)��1L���p����*�Z��t,B2Z6�0)\D����+��B��Ȁ0����0G�|B㞒�?����$�?$3��k3E|�����[;zn�'���'�� A�ԥ2B�z�`HKل�ً�i>����=���9'��H�1n��	VyBn�(��6��O$���|
7 ��?0 @�L�!��DJ�V���X�:�?��Rb|vI��R_`�� ��K����Ƃ�l�aQΟ�IS�ڠ��F
A%B��@�C��T�j�|��Y��#�" ��������ѧ�40��:InD`��/�8'�m���v���rM\%��џ�E���' �]{�f�X�X�@�30�FTs�"Ot�PQ�ٺr�����e�H`s�I̟h����D�7�؁�%͡%lD�����*l���D��ǟ`[aMTD����̟�	�D�;B[��� F�n��D)H�`s��A3c���GjZ�Z$C%G@̧m�Z�
ց��<RVh��Zt2��Hb%���S:u��`��	ɼ����&�L��#ŮNE�4�_�j��7=����1R�d��Bh�&����'���'�L�(sݬXcs��%J���'E�t	S�F9X��"���_m@<����?it�i>}%�d��I�z� � I
5ڒ�A�hd�|��Fʟ@�	��D���?��	П�Χ@h�2o	
e�5�����1lӠ3��k�DN�^�<�$�!*���3��G��(O�Ȼ!�k��1��E�`����	P+��˄h]�3CVTB�F�:{�4)	�咧{�>-qЂ)�R�{� ��u�_2\�+gF�'���"��'���[�'	�� �f{��#�۞kD�	���'���*�K�X���ҴeV�g?��YI>)C�i�2S�Dx�C��I̟�z)��%�2�hq��)< �M�c���(�I�aiƨ������ɦ��:�dƱT|y��E5�y�
	�0�X&�_�>�:��ƌ�m�ĩ��+a��u9gO�-P̊�F�_�O�H`2�x�ʡr���hW0��$��!s��wӎ��'�p��%�����W� �U����?������i%?�B)?K�|�vAD2��m@��Gk̓�hO哔�Mcᎌe��UI�!�"LS2
�Y��X����˔"�M���?�-����O�O��t*O;`RJ�0���z^�p9���O2��V�TȮ<��Ǉ�s���¯O�ST�ԉESen����̉�Q�^0��䛌-E  �e5F�5E�DW*T�DY���B�� �4���	6��'d�>A�/�:�b�,Y����`$�4��p��p���3�G�cД!������E��1ڧ=�Z�k�d�@c����æG�68�۴�?����?�!�$�������?���?a�w�����tF�9q3"��KW�I��Z�
���9fn���K�t�g̓3) qs�˴-���R&Ȥ-v���Y	 ����b�":x�8J1d�ȩ
j�*O� %І�8�36\t��'*�ɣm0���O<�=�@`�F�0�s�D�t�i�	@%�yb��6�0paN�68PcD�ؿ��$�{���$�'��	p�%1aOF7f��p+��K��l�
3s�~4�	ğ`��� ;Yw��'x�i�3v�x!���B�<�豠CEu�9�g��}O��Bf�T؞J���Y��&[l�<����(;;�̰�b�}#p���UX�ʃ�A/p�N=���/�\I�,Uן<��^�'}��yV+h�5� S���-��/D�@��F �u1�����P�3��	.�$�ަ��IZy��,k�6M<ʂ�E�{\�⨜X�Y�~���<����?Q�O�jP�Ď#S�Ć��5<dm12���D˖�j�\�'�V�ː(��H�'��s�'�R��ѝ7��p�冈�
H��*�3`�Йa���(�%3�NS�q��8;��Ą-��Q�|��Ą�?�f�i���DN㤏W�|`1�%oI�p'�D{��$J
T�r�A�&ݮ�&���ƒI��OҢ=�'D�&��*�؝�cKl_�C�5�掭�M(O�,A��IЦ�����D�Oq
!���'���׮��M3�l�E�$+e�TH��'�2�iЮ� C"�^�է�,�Bo���[���*r`�0I�G�f~�B��g�@��}ΖHj�P�@�\�֙�t`�%G�R�`���u�,��[��od,�����S�Oo��ò�X�QSQ�"&%��
�'6l)C�Dg���Jѣ/���Bl�O��
�`��N�
�I�`:37T�9$�ic��'"����j�9��'���'�b8�v�j4)�x�6���O^?u֩�P`C9q�r����'�t!��v�3�3�|�Ƨ�"4��w)K:%~@L��Q��qD\$k����2��X̧Y�\$+)O.��1.SA��"�K�.�ȱ���r�^�m�П�V���T�|�'^���:ږ�A�|��,�_0��)�'m)��
�52��А�
�/� ��/O6an� �M�J>�����.O
%�䌂)J�ŒG��@J�[�$��7�O��$�O������D�O�擒l��t�1�<�Fq:�޹�Fp����������L�<S"7�Q�}8�e4�?�I���ԚR�!�a�l`뛞m.�����N�mڟ6)��r +!�b$�|RK��� � �<��<����(~D���?i��d)�@ĉ��Y��x{�/ܢ H0��	v�x�h�X�`�=�"|yQ�W�<T
�&����4�?�-O���3%Dt�4�'r�y!�M�ml6��f&��1ⅪC�'��F�jw�'��	��Wj���� @>�'�.���@�2�Щ(�&�C��Ó.e�0�gH��i�Z���dC�Cy"��hۑx*�{�e4O<�c�'�r���-�ܤ��aР�[J܂W�ҒO�����H9�4C$�ʇL��܋%�g���<���T>��: �	�RI��rA���U�-Y�0��vyR�'�26M)���|��aʜ#!b�*|N��� 	NCh@���?Q�A�)=� �'
�+h@R!��4��L$:B�D�ؘ<�5�:%��0���`8%m@'B.�a@�ms0Ԕ(E哒6O��ڤ,@�%I$�0��\��$I�|�	�MK�����'z��5�<T��h��0�3%�2A[��HÔ|�'iaz����,����#`�;<��zHF��hO`��TA}r�IY�?�.�-�1yJ�B7E��Uu�����B�K���I�O����Oʓs\������Q@�`pI>¤<
���<l�������6������+��O��'�~��רֱ�m��$f�,@P�S�K���;RgЛN���J��O��'~ }aj@)5nű�OĐQ�"M���D_�!���'����]
v���WRd�d� 5��C�I�ZѪaӗ��g`l��!
4�����O�Gzʟʓ)����Ą9��8�i�&2�����8}M��'�b�'K�)�Ӗ&� UB!��-7ʩyg�6z=���J^">`��q!VL8�-���_���O.tbEL�b_d)�B�ֵL�V�{���
PT)��*k���Ս��}�H�?I`�\\�6��u�@��,�e�y��	��`�Iq������'Ņ�6�$ݛc+�f�I��'�1O�d+�^�M�l$xG�G�:,PԐ|��>�(O�5c��A�S,\��] &�Ɍ$~�����&��$�<a���?��xDFA񥄗q��B���9ޔɃD���t�p#)I�.�E�\
hџ|Z�Fϖ���1ۄE	���aH~Ӡ��e/+�S�1Q�dDBF�=�?)�����X�`�S��	vq~t2�ʍ��'d��'r����@$>D@S!��PK&X��i>�A��_&�a�"S�������cyP�Ixy�獊M��S��S>e�I�k�	;���gJ���䤒�#X���锢Tz"je_:P|��C�'���O�բ6̅$d���0k��:nFh��O��_3_i@0�/�J�Xq1�j=��1�ԼJ0�L(�$��!#�#,���;S�M�IF���'m� �����LE�5�%�	/>]�S�"O�x��%�N���
'/�|R>K0�̟����*?��L��(��Seo��s�>�n�<�';���Q>�<��B�U�vDh�h�_.y9�JEY�|s���ɚ9��hB���[H}c�mȴ�b�` �$LOX�A���=$�F�p��TFj�A�'�T@B����y����c���l�цC �,!�$Jv�q"�ʜ)a�ř1� +`��I#�HO>��
��R�~E{4��_�T�Ƌ ʐ�#�4�?)���?�(O1��)u�a�����Rx����+Mp�.)�r`��hX����'`���L�,]:2��A�
)�I�`�C��P�$�_�Xy(5��;;Ԙ�+��Z��٣�NɈH��,����O|�mZ��MC�ҡ>�;2Nh8��Y���P�d�d�$C�I�kP$|)V�@�, h�dL |�O���'�剕:b�(۴��iР�ড�!A ��%o!��'����$I\��*@?z�P9�7� c�ax�G��O���9;�mz��<�v�P�'Z�����ј'(�Y�%��L�KD&�8�D��'�\eha ۂOD�:�D	h\~����F4��F`��'�8kr�\�u$ܖ��a��\7L�'����?��H� *� yG.�.m
����	�_�Z���s�ʵ��*��?E��[>g��)h�Ǐ�t;2��U���E���;��<��Ђj>�'�h���ԳGzB�2V ��.&f(�'��J��?���)y������~Zjp�rjǄb�ȵ�5�1D��bGG��(���@�^��myAi=��^�>u�%��aSdT�cAL�L��D@Q`�Ob���J�<�e�ր�?����?����ę#kt�8Q�͟�9k����次��#�s� ���+IZ��b,7�3扙A^��Xӎ�|�`̡cIYx��eA���a�Ɉ�F���M6�3��&���Aa �� �t(V�h0�6?i�P䟨�I`�'����`*��DY���&4ct@�["O
�+�#�?����p��,�"��dX�����?Q�'5@%� I!�=�e;b��%P��i"՗'��5?O�M@���6���\0���;L\�����Y2]Q��8`�����b)0���?��#Hae�^fsri�A��>�'	�^x�'Y) S�`�`��<A̰D|"�іL,�Sfb��."�l����,w&QAL�?ٶA��h���bV.�-�ў�
���OF�d �$8F��
tÌ�l��*���#?���0?� ���5��q�'ghw�q:�QXx���(O�)k#��8jm�W��\U�pS�l3Q��͟D��ߟH�O1�<�'>"#�O;x��D��/)v`p5�(K���wmRAsp��q���d�i�d)�Ϋh@Pb>����B�m��X��_7.�peKg�v�d��OD�K!$��.�-DV�7MSV����g�M�T2�Y�-�Ƒ��dΊ}���cw�\I8�0O�؇�'5�������;Sҩ�r�H	|$xau	r/vh�ȓP�D��
�>
�9�g����?�� ^����q"M����`S���  �1N��ݟt��q�q�F���h�	��<�	�?��,.����d�6̮�0!)��-��|��ĉ�.%����LH������o�deԈ$I��O�S2�׊@�d�4��s"�M��#%%���G�P�C.�xAդ]'+6��'q��i�X�L�~`�;)�&�8PHťj\�9�Dሥy�0��'ҋHڟ���R�'L�䅚>z�!�H�d������oE���<-�0ae��XT.qk���v?��d�|�����'���"u�ޔ+���*\:b��3�Z�t��b��������џ��� #^w�b�'�󉋌q�V�:C�T��f��t�F(���)Th��"�[q؞�:GͫMb��ÊEк0"��N���#bfZ�*�zhXۓ~G���Ƀ_�F���>kh�Z���)D��I��d�'��̂��� �h�n��`�k�4Ov�=	\5��(Ҭ�N�ʐ��@ �l���M����2.Pf�O�9���Ү�8=A��s
B�4�ĩ:!�'�Z5���'�2�'bv�
a(X�+#�=��,N �
��B��+����q�Y5X�z�/<bv�(j�nD��(O�J�GT.H��h��	�V:(B��*c(p�A����ɴ���&Y$5�q�ό*T��R�.2�D�*U��'�1��ݪď�F\r̘1� *6�U��_�$�Ih�����&�[1%=t�	b��{�|�����<�ӏO�Q����掄9I�%C�c`y���9�6�O��$�|�0鄴�?���n' ��E/�pC�0�g� &Ԝ���V�Xs�� �K� I�ǀ]@ \b�)M�J*���/73�(���<>v	��y���z4:X6,!��]�r�:`���j�*��*jܗO�$���!��dC�k� 뮬!�'����?��O�OTb2O� n���ڂS�@Iz���H�F�@"O��hg�T�5ظ$i��*�TqF�D�O6�Dz�O�pl���2���ɢ������'���'W��x�.�6�R�'�r�'��֝��b��"9(��&��Y�f�ȣF����z�6$Y��W>^���O�B��!�t���;�е�J� ��!!�R}�����Q#�.ڡH�27�]�&*�|���Q� t��G󼋡���2(��L��vP�&)'}ba���?1��?ɍ<�����݆&��ؙ�11.�A�O�y�w �$|I �G"3)�y8P�O,�Ez�O��R��yC.�c(�����VDոl���%C���O6���OP���?�����4�޺`�����e9+[\-�T�W3C�u �CªK:����C��|rx�'�
S�Gy2@B,UZ1�R!�3x�89�vO�K�x+����sB���9_��� �O��F�Gyr	��?9Un ���HSl�c�:,�P̨�?Q��$%�`.��9������r'T�����<R�Q�"�%�F�:�m����}�'�h7�O<�8r�U�i�r�'7���.5���%5�������R� �(o��'r m�5�͌-�p)�'>hqTd��'�#M���
��R�s�HB���sװ������#Lݠ$&^�Wf"���A�|��,F�e<T2#d�	~x���Y~��xXSF;,H�O�hX�'�J�?��b�&w����
$%��|��e5D����C�Y`ո��U���:'�=�$0��|��T�h��^�����P/>zd��ǵ<)��?a����ĩ|�ɟF���
��f���ʭsvQ�W��̓�?��O��S�'<�N$���
x��؀	9�?1�4�ē8� $FB4�8���͹F ��SDbB�9��'���w�H��I���S۟@ϓV�����b��d/�i�+۱\y����U�Mk��!}p%)���y"Ʌ�������3�?�Xa2���3%�^�J�#�KW�5h"%��'
r���Z���s��Iϟ���͓$��X8��"�ڼ�Si�a:=K�hH������<�d8���<)�nknz�-�'J%
��%
F���Ph�4����'\���?�&��?��ȟ����?m�	�jD�F$M�a*΄:% �,��{��oL�����l���C��@�c#�x���]��u��P�UI(]k@��vp�'� �M�'	v	����?��w�d�'2��O_V=���=d��] �ƞ_���%�!O��D�2���'K��]��Γwx��m��Y�J��4�'NЩ���1�\3Z`�=��4�yr#4y�F�}ӚMB��Oh�]�?���Kd��(�� +g��ě�ǣ���ܴgN�k�'��h���?!���?��'8��I�Oe�ɱ-�]A"�=L���-DD3�40�,����$��?1o����,O��Û�1�	��6e$��ʂd ���"ORe(C��|p~ �b�V��4���i&r�|B�~�/O�'7��Qt��4�~���[�J��|��X�(%��F{��Ov�1�hB�s�]{n]�%�q��)��<ʓ.Ql,KT)�aK��ſF9Gz"�'�����+�>[�و��iBb���'��9P����5{�Ol$h�
�'���B�eu���q��!v�PIK	�'a�1�2�T�x�"�j�`�x�K�'}��c�`�@��)��kC�\�B�R�'D��:.w��PJ�FI��9
�'�p�T߯=4	�w	R�i�2%r	�'QP�B�`�h���q��q	�'QJU��j_'n���a �%=�M�����O>�D�O&���O�P�e��_^�*ch��)����]������џ8�������@�����A$ւ�&�'�/GL,��Ƅ��M���?����?���?9��?����?a���9�n\	�`O�L|X�J%͛��'D��'n�'6��'$R�'T��~��
�G�<F���а6-�OJ�D�Ob�d�O��D�ON�D�O\�dX3He�e"��ĵ��ũUIԏV#�mZ����	���؟��IϟT�	�ɾL�=xy�W)_=�hAY��٦��I����I�0�Iן����(�Iҟhi!��5se YfʷK4ƌ�ɛ�M���?���?����?����?���?1f�+q��h���u{�Yb�Z�
F���'6��'���'��'"�'�2A� isf}�V!@�Oqx|;��E�p�6�O ���O���O����O����O
�D�,0���䋱"��иpaM[v%lZٟh��ӟ��	��`�Iٟ��I՟��Zpڤ��73��@A�Z��a�ش�?���?����?Q��?9���?1��F�@��A�G��@U/M�6�!q�i���'���'_B�'A"�'���'Ӕ<r�ӥG�ƈ���\/F2�I (x����?�,O:#~� �,"5�&�G	U��I���M!�d̓��Os�7Mu���V���f>WO�&u�T���M̦�Xڴ�y�Y��&?��g"�����D&�6�]� �j���9e��I�o���������E{�O��Ą7 �H,�&%ڮX-����?lX��$����41т��<	� R<;≜�r��j���'z~�=Bt��{}�)�imZ�<a/���BR��^�p����H#͌��S�P�e�_f�9?�'��	Zw�x��/ap��K�� @e>\����!��˓���O��}�F�6U�4Kخ"�]2�Ӂt� ��	�M[��t~�p����S�3x��#��@�N.QHӄ�;4[�5�I��M�ǹi2C�i��F���H�n�%0Q<-	����
�Chn��G�D�eነ�&��̟�'U1�X���i�0��C��	5�I�Q�p��42O���<���4��|��(&
^)2N�k��[�
��1��a�0�IR�O|��&���Th�	 �i)LhP\�HS L$,;�O���GP:x���=�I>H��}�!!>$�G�$I�Z �ѻnN���A0h��3��0h�"�8.���<Y1��8,��P��G:>N�A�3���#�"�#��O-T�+���� |��
ܜg�tq)ݻ���Aàs��eM�+�:mj"���o��[dӂ[���Y�/С,��9���"g�L)� ��;Y(�G㎗�yR����I��@C��BE
��Z�ҩ���\�{˂�x���*�d�B3.F��X�ȓ�z���KƔ7��±&	@Q0�O����͓-��H@P�լy/T� ���$T �L9�9}��.>;'���1� GDP��=X�z�S3CM:����N� bF($_r��{t��`�'l���)@�6�ػ��C	,��@(�� �z�:����8.t�(����Y��DRT�&LbR���q%IM#O��02A(Ėm7�%P3�ڋ����4.C��?��?a�����2����"��'�^,�Q�])5��ڥ ʆn�@-#��'��'�'�B��7`pP��O�Q�V� 0W���f�ҭֈ	�w�<D�\q��S�I�OT��0�:,O�=nK�����NN�,a���	�' d�R�@���a'�?q������#/��@`�+b��W�-ԍ�! l�ZP�!�%E��m�3�5ܴ�b�ٕ3�)9��
3 '���@K�0b��I�a��YL�TӢCߤ:��|��@��-mN�(FF*x�ˤ�S�_�J� f�*_�Z]`1gߥL�eR�d��'��[o)�����"|���I2���w�8}0��@]��rf�A��͹T��n��p��D�G$,=�5�b�>y�W���(�I!����I�p���h�,�˧ń�Bh����D��3�~�O���'|7��Ŧm�	ٺ�v�S9�$ �
�k���Z?����h�� 9#K��B�c��O�I��,��'�ў�S��~r(�>:���QƂ(ƭze��%��˓LӞ�)��iC2�'C�;�1�	�qA��*cI��z��Ȑ3����T��?����4~����H)~{Lpyߴn�X��cL�f�O�Us� H���p�ŊFԤp��O��iD��W�4�4C	����:��e	��ŗq�x��'Ae�q ��]2lzj )P��N�x��'�a���X�F�f���<ҧ �V5�F�:k�D���k�/S��O���>lO�l�D���=�@����.��S������3��di��#�Y!� �t@i� �0n�.�?Q���?��Y������?���? nfޱ �F�	l���aR�_���ɇ��D�	�'l�"H<	"u.
K����͑���3;���ep�,t:�Ƅ�3�,9`�]`=������!!o�t�/G���I�52�V 0�-���`�Y�=�&��W� �^��-9BN�
L��Wz����M��'�������?i��P���V�`��Pb�C�<	fC�*/e�;Ff�u6����N�`0�	>ғ2�V�'T�I�_%�D9���8e�X�Z�D��d���5Tƽ�I���I�H1��p��k>Y��g�亙`Q��%}av�)���%}}�ջqKU/a^��ƛ"��䣌�DVi�z�	# �0ނH0��]�ǀ
u�� �f�8�!'P���O��1�i�ER�_�|�¬��
�;�� c1O���ڴ�?*O���$��b���Ŭ�n1���\~c����"O�	{��Ŵ#/~X3v���ZRf��G�>��i��\�8C�a�M���?��4Y;����훌0q�����~@�5���'S�qa��'r�';V)H�c�H�Ar�KEE�2&��_1��Q �l��l1�C�0AѢ=�U$V��(O�	��M�Dl���-z�~�P��ہ<��Y����ft�D��f���HR��(O,��E�'�������|Հu0�Ƀ,S��%&_X���O⟢}���@=7��8k4#M�)���X�'�F����'vn�'Hb!�]�``�\�eǠ<Cb �wH�V�'�Z>���ԟ�lZ�My�I�!HԵu	�)#0�L5���Κ�b��/��a��OY�T:��r���O`�*K|�D��j9�®@7a�@%d�e}bN�Ec�8 �I�_��J�U���`�F@�OO�5is�T� ~4���CO��"�2���ş�ش�?)K?uh�X?���7T`y�ք�g2D�p�/}2�'�a{���8�q�F�(��*������O�mگ�M���O�PFJ��H�-z�*�Cu� 8�6��Ox�������Ov�D�O|��A8�yW�K�Z��H��!X9wW6t�Hx<�6I��yZIkD��@	�(+I|�ը�U��ʓ\�;B��!�,���ġL�e�g�M�3w�31+G@*2b�hy�ʧbd��H�nňSy�Ε�N̪(�hF{B���׍X<\��,O��V�'�h7m����nݺ��l��� �8��C&�*!��6z
>���%Ϥ1�,�y�+G):u���HO�I�O,��M�d+��!'����O�>���V��E�<�   P�II4�|��ɜ�G9 �
O��D�7$�X� ��G�n%2q���y��̮'���37왴?�,�������yb��2y�J8�W�F*/ p��B�
<�y��U!���yU�U	@$��l��y�&ALjX)��x\�}!���yF���f��T��{�$�˦G�+�yB��)b�.��P�8{�$���H�'�yT�,�^Tis��K��[��y���>�\�Iw�ĺ�"�B�)���y�Ɣj�Z �X� ƀ��#���y2�����[�y#n��SL�y�R/7M8H뒅B�F�+Ƃ�@u�B��B�`*d�ԢV�4a$m�zF�B��
w��Y��g�,���.ޘ4��C�I.,R���ƭCE�=�3/��C�%��9p�.P欑�W�͜49�C�b�&�pr�m��ICNJ�"hC剝B>b�s /5w���򖂍�`�!�D�j:�j��d��(S&�5�!�D�$vp�����0R&|�j�E��4�!�C:8�j�	��М�T��ɤ�!�\5n\N����1����dC�UX!���Xd<�����p�0cc�$6�!�d]*8�y�Vd�v�l��%']�ԡ�#�'oD1O?�6i����� \�12N(���L)-�C�ɞB�i�IڢP�~�����{8�dY�>��=*E��o��#����tl�ţQ�;-y��,lO|8�'gE ���f�it�R��'=�z�8p,ƣw�8�{�'�`-�f��w�d9����d�dL��{" Y3T5(U�v�Q4q��|
���"y�0�0���m��ŮHa�<�C�Rn��c����vT�XP&�+3��iu�9e/L��fʤF��ODM)��P�|T@`o$,�%�2"Oْ-�AcjPP���$)��b��/��YB�����R��'���	��ڶ#����b�3��؉	�ղ)F�W��m�t��KQ���eOi�Yq�<'pĸ�ªO�<1e���.�0P�	�@Z � �IybM\&�
y�dcA�)R-�q@K&�>�T�،V�pQ��L�r=ĥ�<D�<rSV)��H����}�L�1�K��2h~�JO�[�X�g�����<i�b��n�s�J9�# �>�b���ϮZ�ZPXp�g����V�P��%Xq���n��eI怀6p�C5�Z��y�Gԙx@Ppu	�0S�����O�s�(�<eS6@�"�:q�)1�q��산x�����"  TӅ�04�D��N�3X:����#ğ7r�QjQ�f�8��c�
L3T�!���'�px�wn˱[<�������ֱY��鰣R�<�|2ѧ�y��F8 ��M��Qrِ�
N"55v�{�(ٷM� �07MX/&��:˟z!�1�p�I�Q� "k̀f�|Тf,�8����dŊ:�����e���#v���JL�W��h/ʼ��h��eX��s��E�y����Xu���U	q��� Ea��	��Fz2��9	X2"JE�NTl���/�o`��  �V[���&)W�8�I�-�]ʔ�{�'�h1����SFlP� >��Iڴf[��aҪI�L��{4��&F��6��!����|�1AC��1@g�*A�������\�*��ȓ:w�yX �G� έi*M�e�,�Ӄ�\}n� 1�Ȉ .C}��#A����aM<YG�7�` ����8��tX���˓m�������n���
�� �\�p)��17T�挝-F��aH�ω�����$,aI�P�'+C d��!"oĥ/h��ta���2!X���e�q9�7�>����P˘eZ<C�e����c�^8L3"�Z�'�j�J3j��H��|�3bT%��$ݴXmJњ���i}\��t�� �F���ԭ|���kL�,��PX�a/ٶ�ɲ���!��%*ٛ��
�B�������6V�L�!BR�J��z��ZƊA3eY?�`2eW#ܘ'p@+mܼvBY�$]�`�1	�%��:�B�lLX<��\������ɪ~��$��j�)�UJ�L�����I�u1
��G,�!1ܩ�GN@�}j�=I�����3��t��3�_Do��cM�f�rD(�t�v ���.�y
� R-�P�ԁi�ѩ�K�8h�6OL��표Y������GlV%�@��*m���W�<T��	Q�ʛ0��B�I�2�:YF*T�JQç��a���'�����&N�|���O��A�ڠ
���ir*O��f�Z��'j�y��j�1oz��
ɘ#@�l�T�p@D��'�0p�{�&r�O5A�N	YB7D�����4c�D�R6mΨ
�t�bqe5D���0R����f��Pؒ�ybB-D�tj��=b�L!�+	F�x��<D�R��ՠH��,C� E�m
�qR8D�$���I�n��*W��]}%C�8D�����Z�,�t59�j4,y�@
��6D�Pu�O3$Y�yb���P���:^�!��Â!�0`T��?B��i��OD1@�!�Ҋ'��iJ@���h��#�$�!򄕺�l�j$��|�
��W�=�!�X�ĸ0�LZ��53���!򤙁��|{ҥ�k�d�z�A�h!�d�r1,u���2.����1ɍg!򤖞�"�ˁ,?Az�uz�jמ!F!�R�]?^|�HW�A��p�ș"<^!�� <��᱀�%~����g�y=!�ƀW`�(�UN�u���<�!�D� slLq�tHΣS=P���K�o�!� 9���w��EJ�@u��3E�!�䉽u.�@�S͋	~��&֚r�!�б;X���f��2�<�a���yx!��<���T�tԑ��� |!�D�%�4+R�TXvz���A	Wg!�d&p���$��x���1$��3[S!�d��P�jEb�����ҥ�DΧ_@!�dA1p};��B5I����$\�-K!�$Ve�l�p&N*fL\��D� 8H!�
R�*�(���OB�)P#��!�54>�0"�n�'6��6��>xB�I9�̲2�YP� �C�:�B�� z�D����/6_����eN#n�xB�ɧG:���G�Ի4�`��O�F�BB�ɉ���p)�������1�
C�t���)�K���]놆�$ �C�ɓ!(F�	h�A�)�T��;-�B�I�}D�u�酹X~� *�h!s�C�I�Y�<P C�)M�\��eE)>tC�	�I[�oL4H�u;B���"C�	�ePL��2�D�i��u���D��$C�I.Ue�!At����+(O�i��B�ɺ�@�`c�¯kgn �@d�w��B��`��|��E۱h.�U��M.B��=h:��	S E24B�cR"#/BB�	/1�P�X��O>��	���%2.B�I�v_TՓeEX��;ᘋz�B�	�G,�l"��J����Z�'{�C�<h�Qk��Ѯ&~ZAA�f�4B��h�<�"�%'�VU��fA�pQC䉨>���Av��K����ܞ!�C�	�0E���L��N�gH�$hƨB�-�ȉ"�6<Y$���DzB�	���B��=�ܻ�I�Jg4B�	��4��Iâ�$�V%�B�I�Q�D���Όa�T�Q��C�I�l�	@�L5H�����58�C�II-�Qz3�ƶc��Xu ���B�	�	����f�Ӑ**zPtH�Z�C䉈u�HƑ�i�
Щ�qݦ]��S�? ZU����/y�v\ٷ�D�[0v�`"O:�`��)+��H�bC�3m-�\�2"OQ������t˥bʯ��p��"O�9��FǢ��q�tv���"Op$Q��ܐ{�"��N�71��q�"O�\�H}�	 �m�^��t�#"O��8�꘾}�hQ�썵6a��"@"OHE� ̀�_?�q��K!6kls�"O���E�&��8�IRSR t��"O�$H"��/j\���3&�^G�TX�"O� ��N̈:Q���Ee��n"�}3�"Oj�I��ۡx�b�c'S�B����"O,dKD��{�K5kJ	�<Q�"O��c׉�#u��Yd�ǀL�,�s�"OVā�	�'C���v��kbz��"O&y���G�ܞ�p�1����"O4Ԩa�)�$@���?��5rD"O�@f���y>⁪�b��P��"ON\30+��)Q�"�k�l�Q�"O�;Gb�)q����59��#"O�d{4!�G����� �0�H�ȇ"On%�MT�Yv��(@�P~Z9z "O��S���:V\|cA^�	}��q"O���ұf��L�(��Ae���"OnDٲ�өL[�(kP(Ԍ�$��"O%��@)���G�4xY�"Ox�)Ba�|�{%O ^�Ε�'"O\�j�!��T�8� �V��%�"O����,Uf���#
��U�0"OD�* F @�b����D�D�bv"O��k,	D_H-	RD��ZPp�"O�	hE蓍bcJ��TB�*�z$��"OBE�児��!"D!�R� ���"O~��G�@�|�|�/՘>���S@"OpyA�p�t�q)k(�"ON�	F��S�dD�[�.�p�� "O�Ipj�#�dIa0@I>v�Nm@�"O�4	b��
��Zѯ�Gi�M3r"O�\�S`> ��͒�	34��"O��A�(�
!�bm�6�@�.6*��$"O��h��#���P�L�5kvH�[�"O2LZ��ˆ<L�$���X�f:x�"O���ǡK����`Ԥ2?hi�"O�!RѤ��"jp�	�('�x���"O��Y�$[r㴉C7����t"O�b4˄o���8IG�	���s"O��B�%��^� �K`+/b����s"O�x*!��/�*��tj��ȍ �"O|4Ⲫ��	0�;��B<ݼm�U"O���B)G�O:PX� ���\p{�"O�|�����t$*v�	h�X鈂"OF	�(j� L��┘8.���"O����+�Đ ��$u Z�*g"O$QG�8O�D��E�ās����"O�#�h��-juBf[�u��0�t"O��
�CݑP��c�2y����Q"O�آG)�>mPY1�F7��0��"O>�ҥͼu74�P��@�b}	t"O�)���Q+�V�C��K�@�ȐP�"O`T���\>2���
dƕ�{����"On�Y�L��= �DY����}r�"Ot���n�͢��C#k� K�"O�%#¶U]�ʡ�.�~��"On�b7Q�PD� �e��O:�Z4"O� ���A ��O��a �O60N���"O|9Q���a�.��oF�K4�q��"O>�yD$��~�ҎJ`:� �2"O��0a��&X|!3�#ֱ�x�"O���pɄ�`�}ˡ"��_>>�A
O�}��Ⴙ/��� �� e"��2�yҪB%>����!�5y��E@�ޠ�y
Tj�R�R��F�tt"�/��y2�O�A� �8�
ؔFK��ԇ��y�� 
"�0b�G%?�~ѩ����y��]R�3�a�:�|L����y��;�l�+@)��ڞ�@w%�9�y���w�@u�憔�x�.�7o��yRJ�����jS#k�f��DO��y2$O�2nV��%_�ay�{uj��y�P1tǢ԰�j1�H8��b���y�_����ֈޟJ�b�����yR�
�g�5�ЄʺHU΄QE�;�yrO�J�HpRJԄ2.2�2呝�y(�~\�Y����PQ"�'�y�@U����2��h�|��ių�y�G
%�Z���IO,.q�-(��O�y��f���W��4۴ �t�H��y����PN
S�"+B�������y�e�?U�}�B��R7xH��+��y�	�D� Dct�N13)���$
I��y�@0J����*
�'��D�Z�yb@\0%���	���10x�cUV��yr��?BU6��A�(6�uҕLQ��yB��c��A��D*��ůX �y�K��]^"�iFB ���GD��y���$,�
W��iJB�B��y���{����d�C��~��PI��y���;d|;p�!�iu%[��y�CS�;V�x֭� �h��ⓒ�y� �&y?�Y��#���{��Ԏ�hO���F'B�`T��OV.TD��#�
�"!�d�v�t�#JB5T����3 FpjFGa؟����!`����!��A~q#�&=<O���%��7C��?}hP������Pqe��_=�9�ȓ{�}�qO�S�������^x�'���ש�;}p
p#�/�n"}�D@O?&	���&I2WҀ�6�l�<��Xj��R��1���a���9p����M�6-}�����L>�%���t���õ$��G�p۶Ji(<�荚N�Xx�ɒ+�\��F�.=���`���W�-���݀9����ě�>�9gE%#IJ����ʆ��x2�5]%*�'Jے�𠡗4>eV��BB�*!��P���G�f���'�^E0�٦?��mȶ�Y�Dָ|"�OVٔe��"I,p�B.śh�`9��k-�S"�v]��胺QJ�E��%�-w�4B�ɪY�d�ۤmN�d�1��'z|���B��-���­`a�2��b��'��H"�ӓ�>	8��B��jt�� "�I �a���;W�.M� ��D�(���+7��e����*��y�*ƞS>��P���HK>�-J�����ɣO.Ui�#ʢo���`����D�v����MَI(� �JP)P��C�ɑRw�؃�j�	N!
��#���SB �K�3��:T�(Q>��Q�A�8�ƨb�/�h�`�Gh<D���5K��y	~����z|���3��?sDi���ϸ��V��>�&4�}&�EN����8Y4ҏl$�� %�� ��]�pn�����D~Ar�ۢش	��ά,���KG��p=Y�F%�nd�R%�8l�%ES~8�0��EZ�ؚ�S��$-9�ŲW隓fꌸ�+��PnE�Հw!���1��qA+**Y uS�g�6��Բ� �<{��ؘ%���@�Q>9I��H��=�0�
���0��=D�\i�@�8��Ԃ�5{`�mkb˵6��`U�Ơ�?��˖6���>�O� �t*�te<���>~X2���O�u(��7�<���k����@�˲yS,q���<���E.f�v����ӛu�d�� �ªj�џ�a����4���l��BM��x ��ԐQ+�1z����y"��-$|��r��Cά�*��Y���d�!F\8�2��ӄo�  r��ĸ�)�-�X�C��b�j��b YǊ��둬,$ؓO���が�<I�K?,u�[��Kx7V��Ǆ�k���H�[�nL`cc@ۘhn��A�W�l�4���Q����4萠p���P�<��EB�À��?m��#C��3��	�A�@$D�Ի`.?}�T�i,A�N�!���<Qծ]�D�:➢|Zu��)[���+g �	t8�7��@�<�Ѯ�`���F,�%p,�Đ'O�0��Œ#G,O��e�O"OǬ���/�?A����'̼�a�R|p��	1�֢/���C'�߰_",d�OZU0���E�:ıO�8
�0�!�'�,��)��8��'$�e	P �B�bԛVeͥ�V���'d �A� �0d�Y��B.0}b$���)��>yd���$OP�#�P-`����.�r�<q  �S!6��g�5(�}��EG� Q8j#?�&���`џ�������CE�l�`��K6\O�Q�3
�_~�h�[�V��!]$.�T@i!Ʉ:B�Vl�Q`%�O6���g�#;�`�T�*	~��R���$�n��'a�a�P�"���E�����T��%�@��'H�!�E�\��)�.�-$��x�deI�P��)O��!�Ń�]�$�E�,O �Z`f̵x4�I��6�Iд"ODmIӄ1�8���gʮ*�TkdMĶt�(��OH����h�'W�Yp��=��c�K��7�j0
�?u��Pt��8i+�)}^�$qEU)\��B �Z�V0���Q�T���	�CF݉��}>DлV(��n��\)�C_�����=�Dѭ�<q�'y��[�슲#�M���
`���

�'Xt�AT��J@. /X��+�MGqyB �@<`D�'��a!��~�Ӧh޽�6�]�^�zAzA��<E"�	��$D��[׎�3SW ��E�v���sf�Z}�x���Y��H�s�ԭi�Ɖ����|��=%bB��KI3o��a�L	��0=ᡬ��w����E�x��(ې`^�vs���lA�%�Ÿ��M��k3O�+KeXfN���<a�i��}6����W7sS`ѐe �q�I3�`Вa(j�2Z��V�u�|��'G��$Q'R{���G$F�i�C�\�B�	�+�f���@�Ac|�a1��4K���ֲi�PJ4`�|�����T?1�n߼K�,�/����@�P�I���ц\bh<�A��l%���c��txd4QE ������y"��
B����d�R����X��Lo��2Rg�`����r��l�N��> *����'N���
K���B��t��1ࠁ#5S���4�|AA�^�z�5r��'�H<�[
�l�+x�.9!H>	�#%8U��H��b��~r�id�(۫)[� ��Nd�H��D?H	���%m�, ����',�D���^.}' �	0��y �'����s
 ?���	^gV���엉>@.T�uD�TpC�ɊR��=��
�'x���'��n��*Aaͳ��D
A��F�%��RQ\�J�RW(]��B��k4<OJ�PS M�H_B��c�UE��h���6�*Q8f�ޗH�Ĩ؁�<�I��T��J>=��ꤍ�F�p4��Vz*�'fp5��F.:����'�܀���?	En
��� ������,u��	�'R>1p��\���0�\�1"�#W���#����<����<������>�&"J�_NB=)�
��2f�l�3�ph<i�JN�w��xP�T$� �7�q�Z���^1X�� h���0�ORb�<�& �� ����c®I˸�!$1<O���gҎ	K��%,�/�|��kL�C���	�d����L�<)g�ݏps�BvŎ�V�2M��`�}̓8�ƍѪ;e���f�}�O�X��*ȿ	��!�%g�}�Q��'N��Bgm�2%؀I�S��<y�Ե��4V�,Q����S�O�L�q�㞳&�<(@4ǁ)l�ꙸ�"O��"�ݣ/HP�	����f�|�2����&M�8��	�Pl�H�\%&}�,Z3CM*]Ql��$��h����f� ���S�ItX����cԝj��(4��)7%�rPN	"��Rꪜ���;ړ/��L��B�B��qJ1@�<4I�
�8b0�"Oڜ�p%@�z����H�V�"݀A�'�r0�W���O?]��˸2i"�qr�\�7�*�K��<9�oJM9���pW�^�v�xg�St~���=����'��3&�Pd��R�B�Y7d��!�1r�tq %���M,��s��G,{�9�'�ԝ�rB
�3I:m���#�$-����)iT�%����%���@��Y�i���F�<6��?�:�XG�[>T� ,��Cy"k�.yPb��|R����(7����H^71p��rM~�<!�GBO�5(�E^&!)�(IV�I<L�& +	�=l%H�H3��Y�tH��W-&����}�$R��9qh��Hq�63<idI0e@!��@��0���?=�d����1�џ�ƀ�/{���>јCM��A��F 4f;� �QO3D����&N0YG���f_�	Q�h �o�<��׻=!&E�<E�d��&L���vH0^�¬�r��/�y�n�}:I���A�ĀX���=��-āZ��,,OBtp��&Qh�}2f��+��Is�'GBur���K����!�!uа�A��2O�zC�I�i7���eB�58B�1AnJ�I�4�?��b�)W�Jչ3 ���� !4NX�M6 �"O������ ������<���qqT�l�ׇ�
�ا(�ҌJ�b�	��2�JQ�V�時@"O(�j�iXr��Q�.W�mXg�|�&8����D^�y�Xixªϝk��J�N-iN��LN�9+Z8	��efA���"�vaq��54��3��2f@$��K�1a�({T�$O�06�IO�p��C�&�R����Gl�C䉉	~VMy����J���A C�ɖ @���'n�b�`��$CĴ]VB�I!{xL���]|@���n�B�	 A�j�M�+wކ*���2��C�	�&��4�5�w�
|�2E��-FC�	0Ɩ4Q�$S�/��ݐb��	(C�	|����0H�6=镠�7��B�	��~}��ܑbQX�2��4S?�B䉚t�␳��� .�$%#ȗ���C�	+sb hqʇ%��8�hX#��C�ɴq��} ��+"�L�	X5(�C�I�J~H��Q(iƒ��ѧQ�Q(�B�&`~��� E7#rl@�@�(:xpB�	�2�tJԃԂ.~P���"Pi�B�?kܝ�H�1qE8,bb0�B�ɾ6.l�k������D��m�C�	�3�����U�ک�e� 9KB��_:|3�/����Q�E>C��2{-4�;"�ʓB�RY�BN�-`C�I:W�b|٢FU�aĊ�3	�(C�I�p� C+��?���1��(6i(C�	+D��)�EU/,
lDa!�M!�B�	�r0��gˊ�b�-{3��C,�B��	Ii
����"q��e�Q�)I�B� }�V�i���'Pnt�zR	�(;XC�R�aP��)f���ر(�C�$C�I!]H㶬ݫ%�8�juA; )C䉫N	0�X�	�L�,�9��� C�$8*���'�P�t�!r��N�e�FC�ɵa�d��U&H�C|L�Z��;? C�ɛ9�M��\
ZPs���w!�	_6ʜ"�cé-T.d�G�ΌJd!�D���b$�dLO)E.,v��!F_!�� ֍��R�wZH���?��q�"O��,6Z���fW�t���C�"O���Q@
h�{CdE�S��x"&"O~|#�� 2�� �Cлj��9	�"O�2�$�v�1���]�`��0""O4P2��#/�zm(Dl9��g"O�%����`�A�4B6�Y�"O��e
ũ.P��Uc3�x	d"O@J&gL�;6|8$ė4,��+�"Oʔa�j�$&�2ą\��Xp"Ot��)�b��Xr�C��L�֑3�"Or!�FE�6��Q��'�!%�x��"O��2�!O�=`���쐢D��mЦ"O|DhQ��/�"�Z��Od�~�i�'�r�YR����vK��	lS�'�����2YW�!�.T�.�	�'d�U�ª��-��j�f�&��=��'�t���:�|A�SJ��:�|,2�'08�K��C<>�����?L6���'+������ Fř7I��Ѯl�'0��B1Q�sfH֡.�֐C�'(���2ظ�$n��ق�'JU�V�V,1��𣢘�A^ء�'��<[�J�E�4-���:�88h	�'�\4).��{*�,:�b��,K���'��j���a��U����
����'�*��wEPbYP�KCϑ,G&,��'���e�=pF"��r"��l}S�'��	��ӱ7�J�� ?zB�"�'���J%傛T��i�C�T�c��Ԙ�'� i�q$�$(�1 c��$]����'?�ţ���H&�J���\�4K�'��;�1�:*��Z�B�0���'�cpJ�R`rQ	�ϔCM�Q��'��a���!�=�`���C����'CPU�cc��K�"�q5�W;z�R�'7�� {m�L�ԃѨ#r(�
�'0<kGo�@�~)�t�	eC�y�	�'\> ��nY�Z�� !���c��}#�'��% '������ Xި �'b��#%�Y�(�t��_�'$�1��'&�Q���s}���o�9"�y��'&h��b��?JP6PW��R�lP�'�A �jP�
*2��6d��"#�! �'�6P��t( ����i�' �(�$6���{�F�6_Z$��'��ma�:����׹|.1��'#�q�Ŭ��ik�R"���	�'c�uPr��14�(�@��xdr	�'�8|�k�,|/P�b�B�7���P	�'�����DC����jK%R�h�'�Ls���	~���B��
��p�'6ك�5�XxR�n%u6��'��T�?�r}"�$�"} ��b�'�^Ĩ��Ԯ���戌z"Ap�'k֨�� ��mjLu��M�uG�BJ�d����F^|���[�w����aW� �����>��/GY+�(X�AP�U>�Mc�d�q�<��N}�l�ƈV�AG�D�Cf�<��T�e�Q��3�"%�)C`�<٦�����3A ���v�)bN�a�<�4�%��|H�J��E_P�1���Q�<�
�~Ę�	�=�B(�P��e�<��d�20���"E
9	���r0gc�<� ��9w��3`�"M�b�T+�8�3C"O�I Bʕ"s+�4�`�J��YI#"O��ҧʈK�� ��Qu����"O�� �@�T�u@�m�&]
~�ۆ"O�1�ф�TбK��qb�<2�"O�����hX�����b�dѡ3"O����Y����Ȓ?9ל��B"On��&*E�P���F
�t`��"O.=�k �:! (/}f@�"O$Q[��W G`f��$ɯ]B
��4"OH�2�'���X�eEA�仅"O�����I�|�i�I[�1��P"O�T�f�.gzPd��	�0���"O`A�t�"<�B����B� �S"O���s�Q�{P��P�a%.x5��"O����Â�rp4a·v�5;�"OH!�a�T�Za�Y3�EK�r�I��"O���tE9oʴA�S� 6���"O�Ix6��2 ~fP��c�6��s"Oh���h�#�60D��$w��I�D"O�u�f�
�������,��%(�"O�`g�E}�>�Х��=�*�ۣ"O�R4�ʅu�֭Y4a�p�����"OX5�4���(��oQ3�]�"O��q�� ^�st�̯7w~M8d"O DqSፗ'"�	��knl,�&"OH@sR�$R���
ИZQ
Q�"O~�(Rf��APj�;�*M�F��,X�"O:A0vA͐<xڐӒ) ׌�"�"O<�CD��;b�v5�T��/o*d�D"OTZ�C1N eH�eәU�-R"O�;�����R��S��a"@��"O���N��(dP�7�`�h�"O��ce:1��]r'쒕GG���"O��ȇp#)@c�� ��X�C"O$�Q���D��Ģ��с`gP%"Ovi{��L3x0�;�(
 g �(�"O�]�w�Ê�@k���Y=�L��"O�uS�Z�'Be2�F�`��"O�H 
Ӑ� ����?�q�"O���E,��\��҃\��(�"O �b�W�	x(� G���B"O�E�e�eȤA��%�,��)h "O�1j��Ǔv*����n�� ݸ��$"O��z�lT�ҥk�N�:rX���"O����_],��e�V�&��h�"O�p��e5 f
�E�: @���"O�F�ˈnipC��_�-�#�"O};�U�-u��8��~!|�!�$>P*��#ʚZ���:��J(]M!�$� |s0��S�~Ub��K1&D!����tt�}x�7n�&01eA�CX!�䁱`��Ӗ�~��Ȁ�"�-1�!򄚱+ "�J��E�d����I�!�	�'k6��.&�(L�#��!��<����J�0���Nұ�!򄜃�0Ċ��˔T���;m���!�ީwм�*���iMn�ˡ��k�!��"_@xm��ǂ
�����
/�!�dɳQ20(���֎m~�5[A�ʳ;�!�d��V�֘�%7jM���R�)�!�č#��!�Р�h��XB�7^!�d/F���x�D�5�*�
�!� a�!�D�>N�00᷏\1�q2���{!�� p5�
�2c�Z%h���@�X��"O��g�KeKD�U#s�=�P"O�)�AA�P��X�_�_X�(3�"OH؋R�X�m�T �D_�]A>�i�"O��f��l�$0�<t*ՠ�"O<������	�j��&�? ���#c"Ox��sD�$��
�R�FװiAt"O���fOG.1վEӠM�,'���"O̠U�O��i���	��Q"O��y��ûF�� ��L
E�"a�2"O��s�J؆�d�/Px�� �r"O���7Sq^�s��43�h�9�"O���@ �R�Ȍ��
�Xhv�0"O�%�5�2 ��Bbڱo �;�"O@�pkQ�� ٚ�&I[��v"O��Y�E㨥�tX���'"OD ��Q5�Δ�c��5�x�R"O @��Fȱ
,����B�-n��ۑ"Ofa�c޻*m�Izȃ1 pD��"O�7&��8 q�0�P
@햕3�"O�"ǩW%�h���$?��Ẓ"O>�+)]�}�VjG/u�F�Q""O�D��D�g<˒	�Ś�"O�l���Y+�F�`�AD�b^�8�"O�\�#@C�pvʘ�O�4����"O��B��c�d%Y�S�t��pw"OV��SN�)N���0�/έb���{�"OVI���,!��pe!O8U@�L��"O*|p�G�W�Heq`�&� "OB�"��A�r�25��$}����"O���QM�$<>�ѱ�b� %g�D�"O$�Yvi�l��܃�d��c�����"O|���B�j�,�rAFN�ba�"OLEµ&R�t;��SB�h�8#"O�Y�,U�V�Qx ��,ĺ��"O>�1�E0^�5�DAף9a�d35"O�[�~y�uбO��w�,P�D"O����+W;L�f.�OlRPb�"O^���L[?���aN��uI""O@\83 �-p�\C��49L�ku"OZ���O�<?�PW�!Sᆜ[ "Oƭ���:5�^4��Ɂ>(Иe�V"O�Y��$Ӳp����i�N9��"O@�U���WD���e*8*fѹG"O��⧧�r����RKQ+����"O���P��.�A��ڵh�i��"ONe����I<��S��F	�Ɣ�'"OZ�V�G0DrⰪ�#�
�D"O2�����;\W� �RI
O��	�"O� I����:� .���y""O���Q�Z�zR���mG�2J�M�"OZԂ����4hڈ��,T4�`rV"ObDbd?����ҧ�86�h"O�d�bm�@�q�]�R5�qJF"O���`������(Q�z0�u"Oq��̉i��Q�)��q�b��"O�i��* �Q�����T
R�~y�"O����6�Ҽ
pbY�Q(���y��L� pY��30M�2(��yB)B�eܺ�H@�����AQ��yҋEHpVA;B��i3�mQ᪏�yR)?A����M؜fCX�+���y�Ɔ/gCQ ���W� qd]��y�e�W"��yS���R��sp���y
� (�Ys���jW�A@M�H���U"OTʀ��)���ū^�(]��"O�ih4��(]�,1���U趽�G"O�QF	�q�zm����{�} �"OD|Zrk��g����)�>F��4�S"O� �b�K�eqBI�.!x��"Ofy	�G��\6��s�I�	o�	��"OpL���p����?�R(�0�љC�!�v���s� 0B��<�!��� ��9���_4N�G �!��DgK����C�Y.|�F�D�!��,$/��S��G�|�м��N�!�D�����@���-�t	�f��!�F��TP�k�U&�d��_@!�ŽZ�� Q�ϻ=7D4�`	U4!��Y�)Kȼze&J�NMX!)Q!���v��!Iw��-aqΈꥤ��-!��4�b�Ƨl��a��)Z�!�Dj����u��Z�"�S�!�d�2� <s�FI�G���R�!gG!�dP�y%xc6ņ�M#$�C1$͍lA!�H�F�A�0Î���+�!��U�*�DH؁Ξ|�����f!�d�J�D9�T#\�6�rp�E���/�!�DR��H���P� ��ϛ�!�R�L)�%S�^-�aB�K�8@� d��Ӫ��"J03
�LcpJJ�m�M�G"O,`AA??>����@�iSR�Y7"OR��d�5R�b�Ih\�h�8�"OP乃/"0�`�ږ^6�L}j�"O��y��գ���@�jP$ '"O��g��l������5^p�Ц"O�H',Y�E�Vy��GQ:F`�z�"O��R�F��O�j�9'�C!xAD�D"OH{�M�7��Dէ@�a��"O���@�o8��`9J�R�"O� �ǃN^�a��7�r�9�"O�����ܺ+�����u���6"O(��s�ޙq�e��@��U��9H�"O.̢�튮J��z�M�ĺb"O�I�2L8�(� ��@�Vq"O�i`�ڣW�x�r��5�M9�"O��F�$}�n�z$\��x}��"OP���ץO�h�P�&{B��"O�a�d�J9j������|��"O�$A��҉��<�i�0P
a�"O=Cuj?^�p(���TcR���g"OX�������F�7G�d@"OH�Ku��z2���wH�l>\�)�"OB8���ٖe�T���F!z�@"O�U���׹ib�  ����+�"OfP��!ڸ�bx�C
�-LS��X�"OH;��d0�����м@:Щ��'�!�H2^�Ds珉��1H��@z!�D��܁�e�I�uU����E�$t!�d� �H#��E�D����[!��Qc$�3!ޣr�J��aGj�!�$����u�4�*!zX�s�N,L�!�2_�ܻ���r����DG�!�$Z%0�9��ޓQ9N��E�J�R�!��h4�!�$�S�YHR��K�&!��A5��As�c�2,aʉ
�'xd��
�3k|�����Y�ـ�'���x&*�61I*!�V�Y�c�֨��� zD��(�. ��k_;f4$`��(�S��yRk�,
�tI��ܯIM\Œ����yr�ճ1^F�
��� �5�yBC��	@����?�`�Q�ݰ�y��U�n�(Ѻ�Y�
l� �O�y�B^S�Ƚ�����i N��y�L�lP�,12�Ӊx��hK#N��y��g�T��N��w�r��#E�yr��+�	r7a](l��D�L(�y��A!� ��6k�.�H� ��y2���6iF�¿��Pm�*�y��2��AK� F���=c��2�y� .�t���p��A���y2ֲ_����P�}�0���[?�ymI��A�����9��� �y��ٙu9��b�!��s�������y�԰FB���#F>n#VdA��O(�y��P!��c�K	X��(�A��y�!n36����I�8<f��yBŜ�kN�����M���udؠ�y���9y4r]�K����Z�jC��yRO�	GH��&��tj�$H�y"$X2_��ؕn�8�ʴѓ�ފ�yR��6�p1閥F� �y�4���y��I�F���Y�%�w�Eڃ���ybeG	F{7mH(s �}y�:�y��E�`�\���x����7���yR����XT�oU�i�J �g��y��
=��x�$��&3cN� �!�Đ�1�.x��Ѷ��xbm��T�!��V0�i#��	����>�!���҈`���_�9�Gܨ})!�]�q����@���bWl��H�
=�!�dǌ04�+���3?EYrs������)��<9�"�*OV>����D��*SE\v�<��LT�z��LS�Nr���n�<�TCW�E�Bek�A.Pd���P�Qa�<9�GP�&ĨD
���-`���kaU^�<Qwę)Ty� yS��[ܔ2��W�<��-H%`�8#��"I�X�2�Y�<��m�M߬��
�$#~���i�O�<�aj��f�P�2 ���?��K�M�<Y�C�v���!��'1��⃠�I�<!���2x�ͩ�.�9m:�R$UI�<�4/ċh l��V��O"����eG}yb�'O��Q̎�>��t�� <$|����O�=X#�P�x:!�2�$���g"O�X+W�I�@�Rc�	F�3A�� D{����ԂTs��-��%�(j�!�$c�Ё� ���^��&�^�!�!�$ܓ ��ʱc�	y��c�(Q�!�$ɂPָ�yf�C���E��G%�!�̝{ڐ9a���GY�aKw�ٲ4B!�D�ZOp��FڭfC2�[4�קh@!��=3�FD��I%nMZ�iT(!�$��t9P5 �'鬁����!d!�L�P��MJ�F�"!�E�N�QT!�d�4�T�s����,����E3?!��#����d�%Q��!3%��F�!�D�yCv���C1ly�݋ ��}!�ɊP�j�����&f (w͔#v!�d؈&<V�hY�~GEc6mG@j!��4�:9����p0���ըvQ!�X� �HS�`@80+��5�'a|
� Ă���`[wF3�v���"O����'"nmKF��������"O�e����av%��b
�}p��3"Oĵ���F�Q[��r���Ued��"O�P90�����5�KS�6R44S"O�10΁8Z�H,J$?H(���"Oܭ�um��aލb#M��]��[�"O�%��� Sb����_�j�&�)�"O֌R�`>4�3����@�"Ox�(�	۽J=����ш*w~]`�"O((�m�W-ri���ɐ�2���"O��""����~a�Uj�&V��"O� �B 2)�h��#��F��Lap"Onp+��D�"���aIF-��0�P"O<K���V��
��Հq�؀4"OĝhЎ��v"� �E���J%"O�A���T�24��%���Э��"OpqK��/M~|�d�x��pɱ"O�͂VA��8��u��(M�p �"O�1���ڒw�B���g.}q�"O��z5�3T:~����_�U��"O�3��J98�X<#����Sd�I �"O)��#�"���8����fR�v"O|���V6+τ@���1yC2p�U"O����JL�U� �g Z�����"O�3�B�IV8�t�K��|Is"O�-�5��5��]ᠯ˸�r��"O�qQ����h�-5T� E`�"O$��B�%�ޭ[���,;���(�"OD���*�`�h} ���p��@��"O�U�+ޤ�nE��c�%�F���"OHP��^�W=�0(�blaD�Q��!��X�q�V��C�8N((��BK1!�dN���T����h&����c�3�!�DA���5脮4"�����)�!�d�2瘴
��:w
4ݱ���#S�!��ƓPA�� n��j^�8 ��Q�i�!�D̈́u���7�B�gS�@ q�N !��1 I��B�KJ�I*!K��sf!��"����5�ٯpߌ�cP��*n!��J	aM�|���$og$��t�/=!򄁊[; ��N�fh:wi50$!��T:��j�BѱQ����畡�!�DC�l�YT�=l�&��'���!�ğ[X}ju�Y�W�T� r�R"	�!�D��;�p�C'����E��d�!�$;:MDqғD�0.�"%j֥��-�!�V,p�A�ϖ&.�}�"_�m�!�K
, �����ȗ=��T)��Z,DG!�.}q�"������ۆ3�!��
�n��2+в��i��+ʓ0�!�D�'m�<A�b4Ґ�2'�4#�!�LaP܈ٗl�PȜ��G��j�!�O3)-Kƨ���8��Ӗ�ly��'x��Xg�&P�)6\J�(p�
�'@|�$J��FH䆿>�A[
�'%����ө! ��b%#^�7���!	�'.lX׉B1p�V�5��Y��	�'Ԍ��!�R�U�Ĭ���"�~�R�'N��@Y�n�\Ap�mG<��$��'&��{�kļL����Ed�(��'nFx��@��B|�,)5\��'�	A�ƒ�R3���1�� &����'lj�i�T�h��]���I�<���� ~m2e���~�����4/��D"O(���V㐙"��:�W"O"�A���5Px8�b��o�P"O|C�G�;MR�:�@֮;�N,p�"O�%����nٞ��ѯ�={��B"O�e2�A�1?��]�LC�*�|X/�ybφ�Q<$�ӗ�B_�*܂F�[��y��վ%U�`Q1�,U���H1C�
�yBHȒc7�@�˜�L�� �@�^�y�͏�%7n�ц��;Iyx��`� �ybKّn��a��K!?	Ψ{����yrڎ;*�C0E�B�6u	�;�y⧖�^��Ȋ�`E�9D6E�1��y� *s�r����83�"��kU�y�F?b�v9ö/&3�����yB"�M�yҊǤ���c�-�y��]�M��|h�nJ��@��*�y�"O�z�Й+��� )� *2���y���U\���c�� �!ʕ�yR��[Eve!�D_+y�jUB����y�F�.�\9k�6x��5A����y�W�D6��e	�t��t���W �y�+��0��_:fz��@�� �y�@
`L���]�q�ǀW�y2%�� �(��qB�=[in}��bZ5�yr� p�����/��]{��[�	�)�yb
ǥ`|@l�n�',@���yb� �*Y|���/ �jE9V����yҭ��2���:���{�4��N���y"��84��"��Y<q���:��� �y�%�ĉ��[@6��p�H��y��_(--Qvi�?�T��I��y�@բ>֐�%0J���.�y�I�.[\Je���tk4NH)�ybOӶp�9tƁ��в�K��yrƙ8��ܫ�QFH]������y���d�^��BLԄf�<5�!���yR�(W���c�'�0^���%l�}�ȓ-8�@2�l�$ZQ��z�Α{"��c��-q����%���"�R�%Z�,�ȓ0����"c�?qm<���O�XP��x�.𳡊	0Y�>�"	B=l�(8���H�rnK`$��=2��!��"��4��ېH�<��+̴z6؅ȓu����KX	_�l�S��͹�4Յ�5����O_4z�]��')],��ȓ8� �X�y̌���ٌ`Φe�ȓ$ኤ(PAN|�ӑ��� ��x�b%Z�J� � ����_2�$�ȓG]�����7A%���	R����ȓ����bM�*2n���Á1��}�ȓ5�$�&#^V� t1d��Uf~��&c��b���*k���Q��0C���ȓ7Y�8���_5�ꄉ�#�z��ȓ9�Ձ�c��p��y�L%b�,1�ȓ6A|e�J�Ti�#B�)��5�ȓ.Q ��*��]�� �dT�,����?��|@�ϑQN� B뛿Y�$���]��0��E6W3.��5(K0ZN ���F���q�Ӓ��4P�m	��\��+���i����-l�-�p��&�E�ȓ7&֌˶��7_���{CD�c�*Є�#Kp�ң��N�̫��)�f��ȓZ�r`��d�?Z	H[��R%-/Ȇ�S�? *1iЭ�s0i 5�7Twb�"O�\��l�8�n(� ��
Ci���"O�i d:V��HB�G�%{�p�˓"Ol0����6P\܅���0Z����@"OH�sfF�n؀5�&�
!܂�"O5�!
�'� ��l�0G�|���"OnX��L7FZ��X��\�R�!"O@)�5�+~���ĉU��z""O���V�K���D
 ��Lȴ"O2%@�#B�YՌI�Fȋ�W��T(@"OZ �w�Tq����Λ �V���"Ox�zR���%���I���:�I��y�� �9��%%;V(�f��)�yr��]� �i�B�.grf�ڰ�yb�Jc`�B�+G�=��C��yr��r��@ǃ�)%����$���y��@ Wtn��(�j��BE� �yRb��b��0�$^��y�Ɔ�HA�,��n��V��y�ɅJIR�0����͊G�P��y��%_\�: �U6{~�"����y��R�����"�@�R�y�/ƦA�ニ�e��� �ܫ�y"@�Z9$h��a��`ۈd0�
��y��V"r�`Xc2��.� f���y���pF�9 �I�
(lД���y��KLqQ!'a�4%�%��h��y�43iޜwa�0hN�����y2HO�aI�aQs�ޘ#��{��y�È0�b�x.�&KF���T�yr͒+n�hq��E@����$�y�&��f�!�!��7t� �m��y�*)�%��m�>k��a3�Z�y�_�C^ �P�g$u휅�� ���y���) &�����m�}1�$Ծ�yr��-�4	3�P�fĖ�)�y����FQ�"̳C�>�3Sg��c!�D��3Ȗȓ�� �<ճ��1_�!��Îl�a"�k͕>��9@c�	�E�!���0�Q+�h�FFu�w��X!���?����b�O�����Ho
!�ĕ ?��T�E'�/-�F��f��0�!�dݺ*8�Њ��F�z�0�D��=�!�D��x!�PBf		8��m*�)�j4!�����=��̏S��M��O�d3!�O?�B�ᱠ��~x"��r���E@!����0ieR2/\P��/+'!�=�������)��I�:!�˥t�`Axvg����`mE4-"!��8!�P ��z�Ty#��3W
!�D��̀�uɑx��ݩЊ�{!�D��!V|���ٴQj0[�jF�g�!��X>2Ϭ8�pE_&]\񂇩F�!�d���,]8���$`�9�+޺�!�D�g6�Ӥ�:$;�2��.>�!�dٰRf� ���Io*���t�$H�!��M�� �q/ �"��O41�!�dC-oH��ע�$}vJUd흔�!�D .uJJ���<y���R�V�!�d	�Ry����S�2n�E
Ӂ�
�!�d޵,l��"�GZ�M�S��v�!��A�D:e��6	R^�Q�)�I�!�W$D�0�j�π/zU�  �4W�!�$���HHb�o�tr�/Pq��� ����F��T�V���..��I��"O��c���#\�BL���'Sj�b"O�p`g�
_�b��"r�p"ObDzq�@;z�P����3R�@�"O&��!�!o��0A�䈅Pƽ�P"O�mhuk��?��M�bë���k6"O"U�a�)f�ܴr�(���"O@���� `~$pta��64v"OƸA��� �Ń�
Z�'�� S"OΠ�ՙ3#T���/� ��"O�i�ק�.fL��G/TI��Eh�"O�xaǂ#R�jUNO2|tqG"O�-��Nc)"����E�dd�CS"O�ҕ� >*]�1�ƨ+gh��5"O|�R��#�8)]�yR0\a�"O��$O�OkH���$Y%�p�"O�8
a�U�uA0Őb��"(�1�"O�P��"z>�dx��2����"O�����F�+�!r5��;~�m�"O��j �����"�:u(&@��"Oԩ t��Q	�ա!A�.����r"Oа��$
�A���G�=����"Oм�*c ��5..]��G"O�b�=k��0l;rKf$��"OP�x�(Ɩg-���D��b�Q�"OX���L�k R�#��E���W"O� )C�̝��,㣪Ѻ@�٩�"O�l�2��;oi`�q��k��A�"O���I���@�k�¶
=\�r�"O�I�5��s�d�5��#@*d	�"O^A(t��0 �!H�#'����"O���A��b5��H��W�@���"O��􌟸�D���H��=��	�"Oz,`������L�#吚""܁��"Ox�cB��
(2$��ʉ��h�"O�jG��@�JabƌZ�E#A"O�}�1I��C���r�\�(�Us"O4�BfP�\`�A�L��	Eh"O�H�癄"��B�k^c5�;t"O,�y�Aw8 �h7$
�.zl�a"O|�ShB�x��С��U)ʐ��"OҕHuk	��2��V�CY��"ON�t�>aiCQ�B\��V"O�V'�.:����#둂:/�i9�"Of�3¡�;���j���2�"O$)�v┖&M\t[�Imz`yT"OH%aa�h\zy��b� 7�!�"O�u�EJKMv��b�3�}0e"O@�r!�ָR9�"��J	�}k�"O�HCQJW~�i[5@�D���"O�J�^�f�b�"/�I��-�p"ON�����'����g�����I�"O\��qa�''��&��4�`��"O��X�)A�RQ8�!cP���HC"O
��h�;O�As�	�d�����"O0`*1��.�69�1$�$a���p�"O�����!�,�hGm_h9���"O� Hs��Y�&�ҶKբH,498#"O��pqL��R�>mc��K>$��"O��{��6	iĥ��l� R���#"O@X�g
)�b�B"*X�T놽�"OF`0ʐ�܊�)�hR�[rZ�p"O�����$M0a��>a\�0�"O�ꆪ��Y)��;���A`�r�"O� �������l1t�#�� "O�Xj�$U`�+�Ĕ�B�ƹ�&"Ot�(Q�.^�ȕ����p�`%"O�<�#�خ{U��!��7���"OD�*�/G�p��pScR�a��Ӥ"O�r�o�Mw���D�@�|�z�"O���+D?8��@
#��N�\�!"O`eإM�b�Yyp�_*3h���"OZLB�-�9_�lٴ*�8/�9�"O��x�� �7p�h��̘5�N��"O|�o[7ǂݓnƹ�*ĺ�"O����逻A�
y�$,H jR촠�"O�\
`8�^����:P@��"O&�q�"�5�LY:����tL�%ʃ"Op�	F$�:s0S��:W6X|�"O����
l���2e����"ON�0�"E%zE���+�r�%"O�Q��F�04|��Ǘf�j�H�"On�s�#�����k�OQ�Z��z�"OL��#B�(��L�N>R P�"O`��FC>%a�X`�	fA�HJa"O"q� )H�>���ɼ�ī"O���&��B�(�{���bX�Xv"O�$!��ŷ2{�c�i_+i�@[�"O~�iG��5��w&\�
@�V���<��
O*���ͤZ���#�R�<�� Ǽm"�Yv̈\(�h�FNj�<�c��*~8pA0��"\e�t�#�b�<�ĉ� E�`<d�� ��YS�u�<���1:�
�a�,,x��Q��o�<��fY.�HؓAF��>h��Xw�<�`@	s^`�F�K�P(9 �]i�<�ĩ�� �yP��tF|���)Gf�<VR�,
���S��pHQe�<�BG�FX<ԉp�Xr0�a3��[`�<A�G0�����,� a�C�Y�<��U�L��,��FS�=�di���R�<A��Y�v��Uzv����@dm�Y�<� ` x�2�5&��P�LMV�<iw�ՠR(�4��̚+�p)�e�y�<���O��Q����"���%��w�<�� I**�� �ݦ[���/�J�<�����`����Z��<�)�hH�<QP)�h��AJ�@8��!A�<�)�JCf�� �L���:2�F�<��gZ&XN}���x8�s7E�X�<9D��F
�S7O�>�Rآ6#�_�<����J��T�Ѩ�Ϧ��6�B�<9�(�f� 	)�H�Ez�4��+@�<�M�!6���C���Z��q��}�<i`�W46��E��Q\ebd�O�<��
9LlH5*�I@��|o)�I�<�` ֙^j<�R��B�8��NG�<i���*q�01���uAq�/D�,�b!�O|8��mG@�����/D����OJX�J�
� �z��G�,D����g�g�Ha(��s�`�p�7D�� �*;@�s�Փ;P��a�7D�<
�c�6����kA�"�����c7D��RV�-!v�1�A�+��0T�!D�����F��l��K��2�DIk3e D��8#H�f���§䉟	��� �g<D�h�""��T��@A��P3�]br':D�[ -��'�`$�d��Q�\�Ѱ-8D�� T��X�� ��F�Y��;�"O��&i��m+�`JE�~@)1"O�(	�NO5L0d��Ź"w" �%"OV��/�Ω��5tn&�{p"O~Uc� ѯI��(����Ȋ�@�"Oh0hnCA�y���͞]tpC�"O��#��L�A^:U�3.޼d�d�t"OR��ݽJ��pGL�-�L�`�"O�ݑT��" d�����g�ک�"OVDj��։_��p1* :N�\A9'"O����ۇ%�n}s`�
-�X1�"O�p�%Tל�C5`�1N�
H��"O����$~!���EԳ]�Fh�V"O�@�q�	$��m�ADB�z��p"O���4G�5j�:��6<p`�T"O.�{$͚2[z=���N(Da"O��:aH,c!���B�;~H�p"O(��#��6�
���c�<�=(�"O��x���7��|�0��^V���"Oz]k񌈑7�2�Y��O�6��	j!"O���*��^��p�ao�'ɲA13"O��@�;s����c�E!NP��a�"O�����M��:E�J�dD*u�C"O���#� �Mȸ!�IQ$"O*̋U�],E0���e���4Ӈ"OP1�bK�F����ԂN=��)��"O��"� ިE�ECQ���}���"O�Eq"��NLN�����6�Ȩ�C"Oz�R��{6��+2�A$�	;"O���c�lH$�'O#���"O
�SD���� lHs��3΅��"O��[ׁ -2|4P���׌5IҘ`�"O�5�W���A�������
�l:�"O8����3�ԍ;V���Q�"O�2`Y�	�vƉ&Ȱ(*Q"O~���d��r6UYs"��S�"O�tI�iș|0��_���
�"O��*�e�N����N�J�f���"Oƈ֧��q��s��^m�%��"O �7��E��`.�JYtt{�"O��p�CU1e��X2vqXEL��y⏛H�$ rk�V�65V�ބ�y� B�m��l:�昦N�� U���y�H��Uˤ!��M�C�<�ce���ybA�u�Ta"�K�6C�Tɝ��yb-�>;���Qs%©~x��y��yR��wK�M#挅�$�"19��Q
�y�B�l��� TQe�Yu�߷�y�E��4]@�%�ƬWc�<����ybX�(0�Ճ!%� � ��yr���`٠%iw��B�:M��jA0�y)
�a^V�Ȕ��Af���*�y�҂v��p���͏%�dU0�A��yB$?E�ؕY���,���aܸ�y��9*�Y@��!O� iЃR��y�댦T�rd�c�$?X�X�]+�y��B�?�(P@�Z�:o�*3Nٷ�y�-@?*��ѳaC0��Ā*_��y�+a:�9� "�Fd�$�R>�y�NґqX�=��)ޮ`k�K��y��V9/�ږ�89�hѫS�y�X1V�	���!�\)A��yRmQ�U#�0)��:�~P�@C�yB%F$?��p��/��U�@��,�y
� �]��y�ҡ�,�)*�����"O�
��
G�0= "*�,�<��"O�e��*C;6z�����<�&��"OFQ���3���@��'4(F<g"O
�	����@9%�D
�	J�"O�D[e&� ��ȪQ��. �"O@��&n�\���s3�����a"Oqh k�gb��lq����"O�A�@�{����.��'�h�R�"O��p��S��T!���sWJ�Q"O&suKVc���,��c��;�"O����[���3,���6�1Q"O����@�)`�ZX[F��i���	R"O\"T/��vpެق)W�YIz�"O�X��.�'��r��ЕC�H��"O�Q��1;\��㇄�F(�8"4"O�b�N�/K�U�QfYOĤ��"O�%���~��]2��(�h���"O��Q�S����*�% >!J�"O�9X5�XTd�@u��/)���@"O<�2`� ��eq��_G�$�S"OP�T��s���֍�	;(@�zP"O��5䚗l�dY�dM�.$�-�"O�tʢ���f�0�@%���(Db��"Ol�;E��b�})V�R�]2Ԡ�S"O�H���T�,9��E��"�ѐ�"O�8����$l�v�e�%p� ��"O8�⁩3q����4KD�I�P{�"Obi�d�G/���G��`��l��"OtQ�s�#qѮI�2��qt�� t"O�$�1 ��xB��K��F&䥨�"O����@�_�huY�*�%\$qc"Oƨ a�U>�p�i�\*Hq�E"O�x�����gH�!�� �%"O�ѣ҄�|�P �D���y$d��"O�Ce��$kf4���\��Т�"Ov��󤘐"2N�3�OO Ӓ<
�"Op(��� �b ���"O���U'z�R���m��E�:)�q"O�(B��ͬ<��m�%��Գ�"O�X�텞@�X����3���"O����O� ���+��Ȣw�3�"O�9�T�I �R$+�.>�2��"OTE�G����q  *
�Y��1�P"O��#��E�F@ZP����~J�+W"O�``r`�z�u�BI7 �4tb!"Opp��ˉI�6��)�/#!.q�"O|��vK�#@�����A��1"O�\+��Y2�!P�ړ}[t؊�"OEcp�X&*C�� N�B��j&"OD|�G�B$��"���.��@��"Oz��a�_�	Or��̪*n~��"O��EA_�'�����@ԟl_��S"Ox�ڦDCPp��A�K[Ql��"Oب�t�����3�䙘.X�E�v"O����h�i�N=�G���BUt*�"O���?H����7<��V"O*���	�k���RR
^,}�r"Oj�1e�2_��8�g��~'��i�"OҐt�B.�bhɧ���}���ؐ"O��BF\`�AK��z���1"O$�fiQ� "�\�����"O��u��*9MÑ虊B�f"O��뷨T�6�젢$H-0�~a��"O� ��;1ئP��!�']�:�6h(w"O��sせ�'�����eBe�E"O�]�To�R����
=&^�J�"O:c�E
P�p��F><hH�"OL�F�ߖQ{X$k%�q����"O��	 ���(�����>q�͊�"O�}��P*R��W��U
2Pz�"O� �m&X]�MBӭ�){�|�pR"OP��V�z�HQ���.P߲��2"O>��*T�fU�M�5%̧)ct�""Ox 2'<\t@���YZ�̨e"O�3��'���ئ+����
"O$T�҄Ʀ"~��!��薌��"O��2dE�-x�3�_�>�dh�"O�]��͔Ϭ�U�U�
ф"O
q���`��^D��#@"O��r.VDu�Ą
V؂�"O�9!2bUHl�h&��?��"Oũs,�qk�X���7kZ���"OX��"c�+��Z#
�yc$]�"Ox${� �l�zظ��>	F�8ا"O�����[p�zƊ˯LtL��"OnQ�k�^MI���d<(��`"Ov�cD��;؂h�s�ϒ=�PG"O���� �"ϒ<��&�hR�"O`���j�<G���`�Cu
j�"O�Ā��H4wƜ�ۘx	�-�A"OМ ��dR�����Ge���t"O֭x�LW�kĬcJ�1{D�"O�(4�L5!�*�kp���_�]!�"O�U�0ƃ[�| �IC_�� "O��`#�͋Y	��!�����F"Ot�p�G�#�T]�I��M��5�"O�p�E�g��YE�G�l��U"O���ԬӟMj��z1���"T�A"O, �� ߅2_&( ���'����"O>��#�x}��3l��r4<���"O`�u�HI@�1��8B�p�4"O<vAU;%U��ժ��!
�"O��#��9�؈;銭I_*���"OĜ*GN� ,�z�m��pG�y��"Of�bS�Sn>�a4lҽ.�ZUR�"O��2T�W�g�����JQ�$�pLd"O� V�?%�J �@��&��*`"OXI�2�Q�=����V�O������"O�� �ǣ�@i�ʖ�;��p+�"Oj�xaiNl�F��RjM�aN|�G"O���D�P:}�.ɱiޭu�T�R"O8E�p� # �t�S��q�2MsE"O.8b�L�E��P���oZ�f�����=�z1�ԗX]�D1D����ȓ<�4F�A"u�ĺ����F����Xm���@�s%������I�ه�\ �aqӍZ)(�b��1h��J��ȓ1�(�xE@�"���e)Ѽ{�.T��F<��kr�9 � �yq����l-�ȓ��0����9�,t��K�_X��4��3�(f)��O�I�Vx��;��$a�`.��"�@)8�T]��6�Љ�b9n:�11`h�,zu�͆ȓN��5���H�?>H�`��T�:���s�&̓M�FŜu0��G�XcLp��,�hI�`�,]��`U%˺JFl��g�h��@Ԝ7*��A&��5٠���S�? ��p���r����>���&"OVE�bⓟJ����C��t��5r6"OD�5�1���S�$Ê]a�"O	���b��PcOȧ,�
Q�"O�:����:Q��rD!�>����R"O�80VQqH�ˡ���Mt��Q�"ON�A���g�HP2T�~��"OR��(��O�j���B�+|��"O ��=T��"*��9��!"O���3)X�r�m*S��~��B�"O
�Y�h�
v����䫜�_�N Z�"OI�	�=p ����MHi,���"O 0B�F�1dI�s�g^�B�R�"OT ��H	<x�YCMȨ7$�ay7"O�QI�&O"p���b�'��k�"O6�{����81"A�v�ژ�r"O�`QE��8`00C`�R}��w"O�� _�!
�����TR"Om(�"/f�E t�"`�i�"OL����
�p��r��Πn0��%"OT� VfQj��y#Y�7܆��A"O�t�s	�,�X�92�l�(-�&"Ov8z�gҕ$�R���O6����4"O��XւN�+�lH5�ףbLf�r�"O�S��	->+��9A6���"O0��UNE�P�p)����aK�"O����kĒ.:����>����!"O������C���������"O��/V�Lq"b&<��T��"OpPs"�]}��E��"�0�[W"O��%���"Q�D�W�V��"O��8�,$d����ql\�S"Oh�1���//�!�"�ԣ{-(�ڴ"O�I�� �,=&����K�]&�i�"OЕ�G���J��p�N5,��Ȳ�"O���㇜Z��A����0�VL��"O6q(4
��-���51\	�&"Ov$i1"�6���m�( �J""O�Yxe,�O��<�q�(܈��$"O\��cU7{�5�gL�e�l�I�"O�h#�h��^*���h�9%~p��S"OTa���֢d�֥Y�QgQ����"O^I���Q�U� ��%bx�`"O��+�䓪e4�J�N�%N�,��"O���V�D
(S� �*"�"O �Y���aX2�R��V�L�쁐�"O�Q�g&<E��):GN�1(���rc"O4Y	3ǲB�B�
�R!k�|t�Q"O�P ����0��J�<o�����"O�y%MC�<a`�H�m���"O�|Iug��|6�pF�Q�^�!$"O,� �
�v� P ���=���2q"OX���%1mzpѢ�؍a�n9��"O^�P�A�zrٛ���J��}"D"ON���f@1Oh"���+�/����"OD,z�h	�u6���5jڐ&~@�0"O^��%���oVp�A�ԻOg\Q�t"O���t-��ѐq���2H��"OL)������A��"V.&��"Oh�Ä�Q8�yP̖���3"O��zSf�f�:���HR	 ��I
�"O$)E+�C:d����R�F~�}��"OL�)Al�O��ui�H�.oB�"O|*7hT�q�Yz�+�KH)#�"O� NЀ 	����X�*H�b�q��"O����B��.}����o�+1�h��"ORti���-0���a�S�~�d%�P"O ۦ����Sc�C�|�΁�"O��� ��-['�����"x�d9��"O8mi%)�3<��l�bdݔ6m�(�"O�i�jW(<_��cT�T�I�q"O��:��.Sb����ΡS|aU"O>	�u���\��I��"�;k�ź�"O�(�S ��.�L�(���wj�W"O��*�R���〠0j|�u�q"O.�D/H0��9���k{�xb"O��b��C�[(�:�C�ot��P"Ov�$��Bd6���!`;�\ӓ"OpT�E͐*Q��e�]�d2��3�"O4ɸT`���d0���+)�e�"O����	uP;f��@M*�P�"O�(�F��J� ���F�<TԞ5"O�)���$}$v��$8�6�6"O޼c���8!$�r3C�lj��"O>͡$�{,>=��"_g	�-`4"O"����!�Z�*Q���6�  �p"O�xY�J,���o�,�:�(�"O��'E�����s&G\r�tU�"O��7��Q����P%0�|H�e"Op%8#��jA�hyգ/+�J�Q�"OB4���L�N��u�vlΰ%�Ρ��"O<�!�.��~`C"�U�Z��S"Oq��l�:7����K�uX4E�e"OD(A#Z�4
���ÖQJ~1��"O��pV���o��=B���M=���a"O����3&�,Y�!>|�H�n.D���d�ܑ_4 ���]���E #J5D�P+w�E%u����i����&D�`�a� -		Q�,U8;g����.D�H�s)�غ��"֐L�Ҹ{r D�X�d��[*� NӁ�x9C�<D�H��S�mt��k��>*l��d9D���0L�sH%�'Ȁ0cTbA�"�3D�l�1���B4-I�Ȟ{��aX��1D�x��`������^�6ut��$�/D��Q�,�c�\CA��,M� )�L9D� Hre�%y���)���8Fa�,z��"D��!FN�&�k��+l"tl�ak4D�`���)Sؐ��W:�v�h��>D�(AC���~�BI؂퀉C�f�X",=D��y� ������$E"�hC@�<》g��h�lŨCv� v�{�<�PM]6BHE걪[.H9�'�[v�<���U�	�(�*"��8ŚH^>�C�Ɋ[MB��Kaz�j�鑒�>B�	-#y�i
�)�?>t<|s��eHC�I�C?��ؔ��-_,�'Z>.S�C����*�7"t�d Cd�*|�NC�'~X�<i����/Y
�� W7C�	.}Q���n$���#�*h!C�	@��Y��L[o�53U�ޭ�$B�	8eiR�:�xr���� v�C�I%22��.D��5��8��C�	ǌ,��KKG�@ԤԜG��C��y7��B�)O�r%SG&ԟcR�C䉢 9�kv#'���ۡT)<#�C䉈��@pb$\ْ�c��;�rPh�"Oڨ�r�@���!�d�F)n�8C"O� �ː��"]��5C�b��U���c"O�չ �H^(0����\��"O�H�� G�|M�`�J9i��j!"OL���F�C�����\�nb��ѡ"OH�P!�Z|\" ���*s��SA"O0M��E�,?^��u�Х0i(Lsc"O2A��$�:A>�$ö���NT���"O�X`̃�q�0�GVP�EӴ"O�|�acқs6��Q������pr�"O�i�B�3V:�	ڷ儶82}$"O�uڲ��s��E�;9��Y��"O�JbaZ0zB,��(P�J��"O��
�J. �h�j�Na.���t"O��*�ݸ����2 
���"OS����\�VN��l��Z�"O��bd�B�)G��`W�߭�%K�"Oਲ਼	C(|Kl�*Uh�*�"�j�"OZ%���"�T�)t��6N��"O��c��Ԕ2-(tȕ�F�dV0��"O�uPlR)J�J4ÃoA*AH��@"O��� �'1y��qAͶ*G�%��"O�Y�c/��9�`�x&��.0<p�5"ON�҄�GePV�j�kQ.h7�$�"O�U���>	��ȡV�_CL�b"O��3t� A ��©�iBt�r�"O 쑂BI�atҴԧ�:)�}(S"O��i7��ĬE0@BE�0�p"O����X�>��{&�i؃e"O�\0'M�,��!�»,�Թ�"O~(�����Z�P���(����"ORE�m	�aP6��e�A���"OtظA$T(+ozF@߿VJ(1'"O��C�G�|c4�����y[�@�#"O2�FR$��ES�#n�P	�D�<�E�F?Z"LCDW��Xp�*Ru�<��ɖ"B ����_�)��Z���r�<I4eζ �
�9W��"�D���y�<�g �.EZ^-p�)�]�HxK�Z�<&E��Xa�����T��b1��D�<��"ר*�pAp⫊�Rj݄ȓ<��<�GΘ-
m��M݈$���ȓc`�=���&%�Ta�I�>6xQ��0�n=�h�3���&Fp �\��L��AE�_�Q-~��D�7�����u0��c��� �v�3'B x[���ȓ���a��8�P+�JĻU �Q��e���alJ�A �"p��1o���ȓ@�*ź�,g��@�ƈ@�Ly�@�ȓ"�-�A�3t.T�u/��6��ȓm[J}P �ܧPz QA��� ��c��2�Ƣ	k��!C0~V���ȓuP�ph��3_\6iZ���(u�����
e�x��,g*(Zŉ�<�5���쉫ӅO��13�O�B��ՆȓW�R�ɇ�^%���{���ȓ~��@��@�z�"� ė[%����7>V�3fE�Sj �¤OI�Zu�`��h���el(�k
�6l��y\���V�T�elP��@�m�ȓ9h\%�T�;JN=��I�G���1XP�-�p�	h`�	��)�ȓ�9�BE[z�v���I�4x�ȓ�f�R�	�V�P�����݇�#^.�Ï�>��d�S��
'9���S�? NԈ��L�Q�����T2D0�P�"Or��5�	�G��v�ۇe6HS�"O^�"�Ëb%:�i@�A!�8�"O��`��7��T������|�5"O\Ī��+�:��c�İB�X�yq"O<�Ƨ%N5�-��¿����"O�y� ��	k^�Q�[��l�D"O@3%�j��1, m����"O��&�T�a0�l�46�)wE�p�<��A5inC��D.�����T�<a&B7_�p� �'�le9��Y�<���6e��)��x��q�p�I[�<�El��O������qX��T��Z�<�cgؔ{_vL�"��7��I{�T�<�2�W�(��@b���- ����G�<�J��2P�({�dh��G�<���Z�5B(��!�ŉx�` 1�B�<Q�T������p����{�<y @4t�|q��__�Z�(Zq�<yF��8�v�����=y(dȡ��p�<�RlK	�����[9[��(1#�h�<wĐ �f1���Y2u�~|���b�<AD -*v��pB.cn�0�$�E�<	��K�1f�i��$(��GGZ�<�"�:q�����ɥ"�� ��@BY�<ٕ�u`d嗤D\�
5B/T���O� Ԥ�7��zI(e���(D���2N�	,��󄛐", %#�C:D���

�'����'�Z#$�I�8D�du�9I+@��%��a�q��)D�$����v�"���p��@o=D��F֚Ĉ�������5D����c��o@�*��eYUum>D�4�q���5aEM}<u��(D��P��.e�,�#͊26c8i�u�2D���D�������>��S!1D��(���d޺舒��;��\1�E$D�(�E�#.��O�$�ܛ�$D����̆}�^I[�bd*��w�=D� �g�;@`t�JB+b�����D0D�,��I�s���XP�][��%y5�/D�D8&ʎ$�cs�Y;%�	yR(-D�hѢB' �r@	Č#&z�S�0D�x�t��2�$��A,F�>�Д�/D�\��fa�1���9W��PAq�9D�,�4͍Y��ڐ�W	��H�5D�8'OR�U�������\�,5D�ĩVD�8�L��n��`�޹:ª4D�Qd�Q?f���b)V8�}��%7D�< 6�ȋ{�$�Qe4h��Ҁ'D�� �"�5+�0��
�t����k%D�Lˀ*Ɗ\ߐ�aծ�L����L8D�ܡ��ΧT� q�I�/b�� ���6D� *e�C�`8(�g$ج4LaJ�6D�,���ܒ}�,�4��r��7�>D�d�U�����r�f��3UH���`;D�ؙU/�2����C֭?T!��D�<Q��2:F<��$� 9��u��z�<#d^=(�����Y~Ԝ�pj�w�<�����ۤ'��!QDL�O<x��m�&-C�9*�}�5oL�q����X5��iB�3&��!)U��M����9⥃_�w���9�GQH�����A�Q;�cL;AV�+�EҶ��S�? D��$�$(6|0u��:(�(��"OD{�j�M)�8h'I%u�<�3"O��X�C�|`,T1��z�R�8�"O4�p�֧����� ��}jQ"O̔C��kY>]�%`RvFI�"O���JVks`��C̛n�a�a"O$�x�bG�P��"�$�X��"O�MB�E\�k�Tq`�'��}�8�)�"O@{g&�*	��,�7�5E���p"O4��&
��Y5z�yg�02] &"O<��
�'N��	���Z8�E"O.	�F��k��+�ř�"�f�rS"Oj���|��h��A�aƱ$"O��9��Y&�%��(��H�|�"OH�fPUKdYPGݏ栈�"OD�� iF�Z9	������"O8�����8�hH0��* ���1"O�L��
4��b�gI*P51�"O��
���� ����:\u��"O��k���0KC�U�?G`>��"O� �'ES�'%ƴ8��/_� �D"O�8�b�]o׊���@	�=��ѷ"OZ����L�pF���en�<��|y�"O\�@N�y��}�L6�F�b'"O��R�I�J
E�%�\�Yv�)P"Od(��j�nd��١1b���"O|=3��08����K!rY����"O��`V����@}�A,�q@*��ȓc��Q�� =j<���L�!!@jl�ȓT�&�K���_k�5��_�c��E�ȓrg�Q:�얗��0ao� {ĝ�ȓ7�l9 �!��a�H�9�-,�H��X���Ё"
�Pӱ��GH�d�ȓg�"U "�S/@���*�e�
p�!�D�!;�v@0���1�t�
Ei@�=�!�Ҥ@��`��ȝx�8d��H�!�&z�J�k�
�q�y�%B��!�Ě>`����Z9����͉j�!�D��o\DqI��4���V�K0nB!�D�&1IR���I����Ga˵W!�d�0&
6�3䘍+l ��M�g�!�䝯U4\��⠌�h����B�!�R�|�D)�G�[=,Yȝ3B�27�!�WF����I��t{U��*H�!�d,
}���(�?b�e��[z!��*�^ҷ��D^��С�W�9�!�$�(N!��e �*/�V��eg\#c�!�dI� �ސ� ��M���q��=!�#}�� ��+?ŪQ�CG}!��2��za KC���t�^�(�!��	}t��/͒ؠ���+�*\!�� =�F� �j�Qpv�Sf�W�,�!���\_�D(vN�+-È�S��F1�!��l�倂�W��8k����6�!�$�5f�S�� �D��G'c�!��K I]r��"�kt�6ɗES!�dɬAFT���͡3t���슇$!�䑦<�fA������X��FA
(q!���@���9c�Z�p������F1q
!��o��壴��/s�G`��~!�N�p���Z&��P���9!��$똱�!Q�I�>m��'ƠmL!�
99 �+�-�8��h��#!�D�04�H�A+��O_��SUd�%'!�� *����)r_l�8�$ъ6C�y`"O���#j���� �-bX��c�"OD�6�
�*��s��Re��
�"O (IUG��*B:\�u��4*0���"O��`�� /�>mڦ�њZ��(�"O��x� Q1X��)��'F��%��"O`3��D�d5j���eC�p�|y"OH9�hZ�	2�x�F���	��"O���Q&ޤae��pE��s���P1"Od���gE;{��aE�u�&�@�"O��K &��H)4��P%4s*qSP"On�"�@K�2�)I���W���"O x�l���Ȁ��Y�#�ݺb"O�����T�T\�����[&�bW"O؀Sa�J[�Ҕ#f-���R'"Ov$kP�ʼ'���!���
����5"Ov���CH1q^�1CD�%~<�x��"O�ĹY�̘3��Ǝ�.�)A/
�y�L#Y5�у�BX�e�|�Q�C�y�B�+�$ě�d͛�N�Cd���y��6KM��p �	{T *��,�yR���i{���(N`i���y�+�|4,��V$ڸ#t"���&�yrdݩ,a t���ǈƆ�k��y"���M��E#�^�H�`- ��yK��1��q4-�/#�p�Tצ�y2Ł�0���0O�2K��2����y�Ⱦ'��Qi�,� �����]4�y�`N0����q`I?U��Z��y���Pf��c�'l�X� ���yR똕%7� �s��T��L����>�y
�����(EiM����O��y� 5��{d���qp���!�y�ǜ�
�ڄ�<wNvYj�bZ�yRg�,;�*%A6B�/FN��8�y��_5MЍ�Bn;D�8 5�C��y���;3�PP�1��<b�Uϭ�y�%�$*����A�}bTpZ�b��y�cߝy��e�A���:�J�-£�y�`U�k��Q���'�D��"��y����H�+���E uዴ�y��na�$țR������J��R�'��L1�A��%2t���B�uެ���'+�HS��R��-A���l���'����R��$����@	k�ds�'�*�b5�[x6�:��.f�fe��'�hlh����z��3�F6CX0C�'Ԗ��C�En9����� ��'*Dʤ48x5�$�2^>��'�dX;R�v��1�Ѫ�tu��'�zC��R/�p�ǌ��l�:�' ��ɇb�|f�b�W8u�~�
�'ZB�f)��K�$@�Ć�`?$5�	�'����%���M�����-p�c	�'J��+��7C��3�e�(w4���'�d0��G�f�R�v���
�'�0�I`�B%a<�aΟbQ�
�'h�l�W�W�S�L\H�D8,�E*
�'��i` ��B<�ݙ��O�p�P	�'༥�dN� Bx�1�G��G�\��'ղp1Wϊ)�`��eP�Cqj=A�'�"d��O	�J&�����=�6<��'�@=1��=V4� $�յ_�|t��' {��#RD����c�7*"�) ��� �)(c��Mzѫ�!5-:֌��"O4�R���+xB �%��'+Jmxu"O���1e��V�z�N@58tX�"OLy���/��4Nʮx.,�8�"O����Y�9bmx��%zG>9	�"O>�Ģ��-����K#5h�j�"O�Q���W��Q�I͠}p���"O�q��	�(*��� �����}@d"OfuZ���w�Hi��	/�"���"O�pb���'5I���lF7�:qq4�'�'�T�R��})PT��D��6�  j	�'{�!!T +�욶ֶ1�xX	�'c���˖�N\����W5uز�i�'����be(�z�;5�s��b�O΢=E�$�E�k����M-Q��Q��5�yr���u��x�B��$z(*�3g���yb ��rh�q�V��p�`��
���y2/�#O���;�o^��&d��hԻ�yR��y��A���J$��''�yrnƀJ���sEC&���Z�y�L���h��ߩ1)�hr&BD����.���P����J�H���ض�13SN)kQ�K�:�!��<xZ9Ԉ��L?l�&(�!Ot!��;P{��A�ɰƚ%��M�$yW�zr�P�)�Ty��R� D�#�ܦ}p!��ج{p�M0@�̙_)^a�wB��!��D*Ϥ�3��,iB��S�U�J�!�da�=8�#�_&�1�9Uc!򄜙xN���S��ȁ3��in��dA�,�@�J�$���9��	]��p0�'La~��M,2l׻<�6 {楏+�y"�* ��`r�P�3Ҍ\#�N>�yr��#? թt�
�6�&�"� ��L���OdʡStͅH�Du�2kȫk}� Z�'u2�u�B#94���1J
9�]��'�r,��.K�4Rf)�P� 0.�VH�'5@����MQV=ۖe�s, q��'�d��e�M	��m_j<��	�_,|#<q3�SIF^�[VOP4{�ԕ�pU�<Y�̅#�
����ӭ3)��u-�J�<a�%�@v����({#������`�<!W�I8ڤ}�c�4��]D�<Y��W+nV(ۣ.!B�� tʊAh<Ad �C�ę��$��n�~�c&���y�
KS�.���#@�Yha����<�y�@6	��j�k��U%`}�$��!�yR� 8��9��R����Sǌ�y"(n�LYyQ+;8R`���y���rM�2�Y�8-BA�7*��y"�Т[���P��2iͲ�o)�yrbTz������<8�j qΈ�yr�,7�=��͇=2\�I1�ԛ�y���@����O��.���J�OF�y
׆Tg��:��ǭ;��������y"�D8�h�!�I^�.�'����y���:�V�;�J�F �q��+Y��MsOn=r�U>l��B�#C���"O����NJ�"���C��B�<@8�"O�L3�m�Z�$y�?4��``�"O4����9y�D��W#+�����"O����@N���k^�Jt)��3�S��y�%�-��Yҕ��5�2���y� Ӡ^O�AH��܊{�DL�D��y�*U�$�<QO~�'G�����
W��G.W)D���� ��'聹���K�^>qB|��q������@��=I�ٕ�̺��؞D���.� v�X9&�\�rh��B��N9��ȓ��ub1e[�X� ׌@�v���'��5�)ʧ:|V�	f��9_lQ���(KG|̅�����"�NzT�G��5�vD�<���ٰ�i��(���B�`�jԄ�	l�C��혇��q���ךH��uK����K�E���t�ʙ�>���?Q�g��nt<h��-Zk0*ф��yB�f]�hJ0��P9>�9�囱�y�g��tr5��A%E��M8�䂣�y�����H�,d���w�1�䓶0>��"B96�XҤJ�-V������E�<�qn��B݂��ϒX�V�˥��F�<I.P�t4{F	�Z�F�����D�<��Iن�̠��F�UV� 3��f�<�t�ǭ8@���)����Gd�<)%��-F� ���@��S� ��wcM`�<!W Q��q3�"��vJ�]�I���I��Iҧ��h�J����^9U~C�I?�0�ңG9�,Q D�+C6B��&j���3h�	��-�.�m&B�I<ž$Jc�ԑz��	�S��456B�	�p�@m:�OB�Xd�F��3G��� w]Q��}�Q7a���Ao��4u�X�3jI@�<�`�ךI�|L#�	�E��-�#��<1 J�{?Y�����R�p˕"�b����5�z�#`\��x��)"與�M�z�*Qi�/Mʌ���B�؜@��-ı�e㞠�Z)[d�m��L�ȓxv�=�1�� �6����9��L����pÅє�V� �c6Y܀��ȓcT���G7�h 8����
�dt��0>��ʰ�Ϯg\�P��b�݆�i3~=��"5|�E����zy�ȓ0� ��뗓%,)�SlK9"�\Ňȓ4d��Pn2
V8h17�̸@v"<�ȓk������L�`�ʹS���67�p��(�=� ��g�b�� �ͩ3�h���r�h�#��v�������$��\�=A�2LOj������ �R/Ê��ɑ
O6m�9hs�CWB�q�.����͔g�!�Ě/ :����#�+�TyITH�i8!��0b��x��ڷ��)3M��+?!��P� ]�YK jT: �PD�+C$w �'�ў�>����֭O�(��	�6j8=S�j6D�p�G�/(�髣%K�9�%�4D�|�ԃL�U	F��6e�ؠ�� D�L�Ra��B�|�c掸X�9�'�?D�4�V ���zuiK�D.}a��?D�(B���Eqp��C�
�8%(9D�4p.Ԭa}b��AD
�E�8�t(7D���+G�'B�M���ۻ\<�u{�g4D�����U�h�<��E���HF�<`F�$D��+��6E��R (e�����/D������6�t5�Tm�%>)�!,D�t�B�2[���ٴ�Sk<�6�)D���B���[��dBё;x����"D��Ҵ#��G��
D�z�\9�� D���7�V�M�-�d�C�T��$�?D�В�n�.z$�0FD�?8cN��"+3D��g떅]5����Vu$�J�
&D�$�D怗/&��1擿s����%D�� �8�ȓ�~���	�HD�e"O�h�R͕�6��z�_�>�Sq"O�M �5X|E�43&�z
�'����Ȥ�֨	�Οzv�y��'"�
�dޜ3Wtٙ�e��rS����'X�r�+�I�i���	m�zѨ�'��o_~4"M!3� �`�X�'ۺh�iR�1�h�(�@ʄ����'�x�vk�����S�_�	1�1p�'(��a�[�h�a�V&�n�9��'���+�0d�@����n3�m��'��Ԫ�d$\U�4JG�O�|�
�'X�K����H���YSG؞Ay���'��pA �$�0 rrj��fe�a��'D�=ڱa�3�N�CSgN�c�9��'UZ�Aר8���g�Ւ]MV�X�'Y"A3�!eN��g��Z/D���'⠡�)�I���� ��:��)@�'�� �JӞ%[�u�#P �ڜ�
�'q�) 4n�b2���)����
�''���LE�)�D�Q�-���	�'�8���R�H�y�
�ˬ�	�'&�h[���V"8 ��(t��-J�'Pj0�B[�D���)טh����'�Pp�PnAr�e VL'�h�'��i�킕;;|�%�ߵ\�z�#�'���C�CC���)r�MB�X`
h@
�'�԰a��2RT���f߲E����	�'V�\5 ̹����6o�`"��*D�$�犏6�>4�0� \Y `)D����/|��D����=6d"`+D�PT�[����Q�n�>���x�O6D�8
�]��b�[&J
|N�إ�3D�l3�ۡgg���v�;	$����1D�y�q���q�k�+�6��GF1D�p���.TU���s:�𽢡 +D�����U�<��ԛ���*�&ѐ�o4D�x��_	|���P�/�6��a`E?D���'P����G��B��e?D���D�	v[|\1	ZWXp谍>D��Ь;}"8ڇ"��n�F�"�,)D� �P���i�� SH'Rj�H$�"D��C&��)]ؐ��Z�#5VI��
 D�Db�J��``�u��d���ڵ�m!D�8��%į����!臰PB~X�.*D����*VV�P�3g��.�P"'D�X�Q.͝e�b#�כD~���(D���p��) � "S�3�lIx�i'D��P ��n�8xJ�mGg��4*D���G�&$Ќ���#G�~ǘ91��)D� ���U�X���1ժĖhg,lp�
,D�"M?]2��Q"̟�)�Dp��+?D�L���5*���S�[�4Z.�j��/D���g/NZ��)ٷ���p ���!D��J��E�(������4�&;D�@;���/l�q�ӌ�8)�,�m>D�����*93R!�6��+O�*Īi>D�� ' �%p�
ܨ��W�`0�%�(D�܂�C� ����aFJ�@9,s�$D�tr���R�*���������-D��&I��g�� ���x)��+D��jTJE74���0�K�=ixR)D�\�Q)o�d䳠DD�f���*!D�,��C��'f��OC<�z�8s�)D�� "��Wί1.���A�%z��xӑ"O��i)@�G��IC��?��t�7"O��#)��t����>uʬ�W"O(�S�͈.�%�1���g�vQ�"O��`�O!
D
��5��N��g"O�)��+p=�4�U�� :F�aCE"Oy�f�S�E����d/W7�b�"O�$m̈́T����d�4��W"O�%���ҥu��������u"O�YPwϗ#r���_�-l����"O�kG�:A�a�LY���P"Op�ۥ?���12@X.8A yA�"O4@�1%��@]O�:h�5HS"O������5tZ=�Rm	"D
N49q"O�d�0aF�*5(���+�FS����"O��0��Z�2Ơh�
K�l9�%S�"O0`�a��0�XR�+_�l+nȡe"O�� ��Yn�5�a�ƾ_uN@@�"Oʩ���It��p���j�ac"O`T�]�O�>�c���?8�nL0%"OĩRe7y�41S��C^t�!�"O�qKp΍7asz�bq���>��1#�"ODU��L	���Ь�6���{$"O	��ɍ+A�@�!�"v���"O�q8��\& &�$�'�0s�d@�"OL-����D�4L`į* ��)��"O�����&����LM�>�PL w"O(�r�<���R����г`"O�5�3���0�*,i�ꕥj}Q�"O$�c�A���ڤV��x�"O.H�D Q1@�>���g!g���P"Ov��@����3��'F[*���"O�Xi6!ʄR{r�2Fg������"O�p����O��@9 Ź�.���"O@��"H� _���1N 1�ҝ�S"O�d @�^��$*�2�P;�"O6����]l Bu�4���P"OTȩB��myv`�v-�(m�!�q"O��z����#��QB�G�u�
"O8�P�!�pٸ0���V���U��"O�ex&�sm���u�6��u"OR�"��4uC'��:a���"OpCt�����!�S�PH-��"O��Z���(��R2�тm�u�V"O���2-�0�Aط(Ц2���C"O5ó
:͚�r�'�>Q��� �"Of���'�*TDY��M90�f��"O�017,�R�A	P��7mfh�u"O� �e�b��P��7d�a�`"O�D"�*V.�b���C5AlU�"O�=Ze܋.���A�U":5Z�!R"OHٸ En���#R�T�*�Y�g"O��� ���A�,c��� r����"Or��� 6LD�R�rn��k�"O�=[�럧��<{7�8=Qr��"Oؽ�#�	K�x�*͸D~�Xd"O�@ 3$@�e�du���%_����"O0�Ҡ�2|ε�
W�l�&�3E"O���b,�f��UkEgR��jm�6"OДI&L�g>r��F�L�D�/�y���&Qg��xsIĨ!=P���g7�yB�;)x؄�U�>gr�Q&o�y�a�-Hz  �kZ�YL��1&��y��,{�Rؓ@c9N�@�еg���y
� V$��n�mz��f�U	$�8�"OR�+��ܳt7�H:�(H�D��*�"O�G��6`>��0H�:,�vH�"Oz�2�$�R��a��7#����"Ox��h_0�t����	eЎdB"O
D�u`�(%h��E. �c��H� "O�C�$�`8#���:�"�`�"Ot�K��[��KT�"O�l|�"O^��E��%V���c��BC�(��"O�1��M�)z���hҙ��q�"O~x��\5	�<�a�g�!.�\�"O����m�8a�EA�ux�!�"O�	����+�(����YUXpbp"O��si4t%. R�-݌K�@�"O8T�3���2&NH�d悓U4.�c�"O�jce�9:<.,)�")���F"O�!��Ȉ$�AÇEϨ�"O-j�b�)��!�Eh���"Oh0���j����CĹτ�C�"O4M�Tχ%K��iҥ�N2��+G"O6�)���
�j� �',�z�@"O��iZ��H9 !��u�^-���N�yR,W&:�r�%���r1��"�/���y�aьb��QC��f�q ���*�y�Đ?B��R�� ^ �\��P<�y��^B@�2�aZ�Of��� A��y���i�(}x�牨GG���KC�y���/��H!�T1E��J�-���y���.����4	!ha3dC��y���+�H7��J.ĕX�hǸ�y"ÇW*J�hVU�E%b����yBiE�@��D��<>H�9�#���y�DA�Y腓amJ�� ��æ��y�/�ν�b ��{� ���yr��"���v.��@8������y�c4D�v�*U/,&��a�H��y�7lͨ6�]63�`0�'Ë��y�CF�w砸(0�?-n�5�6/�y��:��#+U�(����H�"�y���?z4�Ib�ټs3p�-D�ա	�'~)�s��O��K���u�̅Q�'K�x�W Ɋ�,��g��]@�'y갱�&����c&�U&]�v��'��U�*W2&󪼩U�H)'��@�'Ġ����%�0�jpMǳn���p�'z,� �N�qJU.�:9����	�'��p�`D2_�`M�3眐-Rf�+	�'��l�%��Bb&�"o��)�'P�k)��9��(8$�º2�9��'j��ǝ>���da��b��E�'<�!���W�8�@���_Z�k�'C�IC̖&ǜ�ðj ���	�'�(�Ȁ��,]��X��JAu<lp��'�L��b'u��D�h.u���1�'�8iKԔ#��ز�ՔC��\#�'�&D�j@�J�{Ҋ�DMX�'- ��W�BL�:��E.�F�q�'�j��wʊ�):\)�.1 ����'O\�v�ٓ)pPMBD̞+q���
�'q�TpIb���_'6%��
�'���[��C8�E���)�줪�'�0��0���(�!F�SE|q�'�� �cM'����ր�Iƹ��'��u� �:p����5�6LnxA��� ���Bf�	+�b�+Ew��8U"O�e#D�2Jfx��gkY�YE�e1�"OT�C�A����
 J܍\X	T"O�9�:%��vҋ;�:��"O�,��΄' ��5y΅�ݼQ	D"O�:d�+lZ(���;<�F*�"O���e�(>���$,���8S"O^EpB�E�VtuY!Ι�`܊��"O>Xc6MDf�����^�VH�"O�%h��W�jϰuqd���uê��"O��:' �	f[uj��<�2ܳP"O�P���Η@�| PDH�9p��Q"O�QPG�V�e$���qc��8j���"O�L���F/{�~��C`Ix]�m0�"O�!�D uj� ��ZXv(s�"Oh��
�;�p{�I�^�j�iR"O�|�2h��d��1�C#��hr<� "O���#Oq����̣:� a!�'Fb��f����xa�ʌ3hx�R�'�8l�4ʏ�y8�ĢTY"�)�'�,a3.O� �R�2C�P�#����'n�}s��?Gа���>�M�'$X�
0�H,U��2�j��q�+�'���B��/O��B�?����
�'�@}�U)���VɈ�
ڋKzlX�
�'L`@�c'[��x�1H6�F��
�'�N���̩StJU	&���	�'�ds$-N"@"лF�4	oh�h	�'�K�Uad��p��Bo7Plp�'�� bR��6V��bc���dt��1�'MJX��� T�+s�K���!z�'yx�8Q��=j�!����@��'�`I�ਉ>HDɷ��+U�ݩ�'ObТ��U;J8x�wf�Q��t��'�(�ֆ��9h��;�UQk�(��'W��Z8I;T)ޓ^�h1�q�8�y��R�`�L9e�.L]~ �n���yBEّ*�,��G���0�ls�lC�y�H *���b��_>)Ln���y �.Vh��EGW�l�z���Ċ0�y�%�,+�&�Pi�����T��Pxb�7���):� ��F+��M��u���i��%BD�Bq�۔2�|���UP�%�v��"B쌐bm�ȓ @%��>(�Y��DP|��%��
T�F�8�"9A��X�H(\��ȓYF`PBl�%�X���Lt�l��=2��P�!W),R����NY뾀�ȓe�a�A�P#%�F|0���d�|�ȓM�v�����=�-��ǁ*kT -��ϨYX�@ѴH���b���E����ȓ~u�mkӊ�X�;�%L�x��q����l�7��,t��D��� =v8ͅȓ>f�V�>���U��'�^I�ȓR�P| $ �,)��aѢI G|`8�ȓ�hu�⨟�Zs ٕh��f����zy�1)�O�15j���a�DT���ȓ<�r���ޢTXd5����1~�"T�ȓg�4pAfX�Q����+Ү\�襄�Lv�{vfB�j���Z�x����ys,Hq���~Z@�B�n��%z��ȓ$u�e�C$R�}���O;�dD���R$���� �0����1.R��ȓ <��"�`�l�����␄�S�? ����l�q� �L^�dA�,o͒����s��K��M��$V/�7�R`P�%D���"%ւ�Nq�Ɗ�����H�Of!�pn&Kb� ��9k��5@D-j՚��%w��䚓@��ă�.¢r �v���k���P�i�`h`�̌��yƅ�,�,CtN�Z5��JT���'�\�ZUʀ�3)r�@A%9ʧj��a<t!4@Th�gf�!�ȓQ�"24��0|�l)�#m��"C�Gz�����<��Pa�����*��
k�a��ĸ�� c!��71;dQ�'�3c� ��q�]$H�u;�C��}z�cf�:�az�.b��!�n
S�~�´�M��0<1UNQ�q\��F�T%bԑpw	�1+8��E#�?2!�P��75��S�:�C���&�-����'L����-obS�(,鞼����Z��Cw!فx�N��g�&/�B��|T�"g�׫Pd�SKƥb�ΘI���tl��ae��'�hD�,�IJL̓v���C���|�qYc��5Έ���	�#��E"#���-�/=A��8BX��B@8�!����k�Y�q"����ՐV��y��]=M�.	:��҅)L�����5k�,��7霧D
�aҀ�H�"�B��B��|�h�A���b�(�#�^h<yǣӴ(��P��.��2E�%�OS�<���$�Ttq�D� D�.Y Ò�,��@���	�!Oq�S�P�G0��;�h	�:�!���%��h�%��h/,QWgQ�6��e3��PTdI�ւ�wx��?��vŧ�ēm���"�N�C}2X�	d�����`�����w�ȡ�B�!T�P�#r��{r@8
�oݩF'
 :U��8'_ҥ��'��\Js���T\�E�Qb2������y\ �qCIB�s%���6�O�6�T��'8������
�v$���, �
T�3O�u��̸}�� �M���!�i:��!7O��f�=�P�U7k���pc	�u��	 ��\cx�Ŋc(�!3�I����({H���''�U5��g�Zd2CJ�a!R):��Wldx ���4�̕b��T!����2l* �Au�xr��+�q���[�%��	0�%ھ��> 
�5y4���&�%KQ`QsC�'(U�Ue��D��d�ąA�3:nL��EߔS��5��ɷ{:K��P��Y S�1���B��*G���h�(��r�6��bPN@��M��R�pa��Pj3��@�c�&EHP��O =�"�ךl����'ؑ!.�c�i]L�b�T��0[��D�Ej�$2t�D�7��c?�X�t����eϴ$� P�d��Y�B��
B��p��Y1����j�y����Q$�$$��#�^��a�7(�~��A��1O\� ��[�ֱ�bn��*��`P�'T���@�ˉ-��*����Z�Q�h��`2�]Kŋ(V�V1����<��%�$��X��dF��U�A	��wp��E{rf	;:Qz$�!��;g�b@bcd�9f��	B5�DX+Q��x�$[	l!�$&*o0,�AEޅHA��S�CK�x�DQ�E�tX�w9����`��*n?h��	����~2��r9D�8�ϟalr 1P.�P�(!6�S~B��
��q[��䘦3��U"1.�[+4����ana"�M1LeX}I�AR#`�\���/�.( ��D�E&C����@"��!��Q5!�RB�	xؠ@����~��8��<N,B�I�Fx�I�Ga۝R�d��(H�(~�C��� O��=h*���+���C�4]�Ҩ��(�2����.GLC��sG�̊��:t����4C�ɷ0�X�1�M	��b'�ߢ|�C䉓[����bM 7=~��ȳ	{�B�#,�hJ $B�]йsG��8�B�	��4p�ЂE�*����/á)��C��8�>)*"�[�`�*0�H��B�	�9J��GO[�NIp�� #�"�rB��	�1�b� XPٰ��]�C��'3zl���
�2���h^8P[~C�Ɏ$��	$�˿h��$��Z�`ÔB�I�*%@�8qJUB=�pq��y]B�	S@ <��Z�#^���\,C�ɽw��: ��l�敋��˦02JB�I)N��RE�/e�Y��\_�NB�)� (�`�G'�t�@���4��*&"O�@r��Q "Ȧ	�%̀�$�\@�"O��2d��A"F��+�\�"O����!ֵ0#�Q1BC	�=��yr�"O*m�e��$yx�t� �#��Y@d"OF�r��V�8�asGYF̶�"O�h���}梴:�EE�Zo�3�"OZ�˵n������;=^����"O�L�7I!.���`�b�<�)�"O�4���}B
(r����$�9��"Ov���m����P���A �xp"OЄ��#EL?�����<���"O|[�,�-��0���0WȨQ�"O܄S����gy�!c�j�A�T��t"O��2Psy�!�����b�"O|)�F
�PKL�{��m��0�"O.��N��2��f�b��V"OhP�cF/r�)���p�Y"O��QOӓ�r�j��Y3`h�3�"O|�FN�<��`����k��"O��s��\��(s�B�=��3w"O�I�Q/��'~*@�
��� R"OIXףLy-:e�&D#?�yc@"O`��≋'p�|�ɐ�����Ӆ"O�A��e�(+w2U������E"O������+����GM��x�"O�|�t�#ͨ�{�H�? �a'"O*��O�cT"�2'�j�b  `"OB(0��_�|=b�d�M��P�"O�X =d�8D�cd�/U�%��"O���d:g���I�N��� 1"O��+E��/q����H���R@"O��f��;�6Pxp'_4)�2Ys�"OFـ�`�1 ��%̎M�´�'"O� Rꚹb�H�k���6��	P�"O* ڡ����d��-�=}��A�!"O�}�����,,)'ԃ^pl��"Of�+ ��Z�1p`(UT�T"ODH�@A� �	�ζVP�۠"OT- ѣ�*$)���1	�_/4y"OhX5k�\G@)
0CG�sRX1"O����S"0/}�Sdֈ^�u�W"O"#ŉ��X������O3D�h��3"O����EJ#s�R�Y5�?�b���"O�8Je��� �Tq!m�+G>����"Ou(�O�uZ�yꇬ��Xh�"O2A�p!�-O�
�k�mX5[��b$"O�\�����X�;�
p��ܚ�"O(�"�8)�Q����E�4�	�'bQB�#�\1�5��$\�b���'���!}���Z�bI��<1�'T�S�(�?"f�ݻK�m��0�'��س5�^�C�\�&��=Y�Y�'��h���/\�붣�Z�d �	�'Q@��嬎�q���V��$� ���'c(H��G�)���Ŝ�����'�j��6�E��K��s(�8BLGH�<9UF�5[��S�����'��E�<�6l4��!ՃS�2���Mu�<�?Y��HrM!�,4��ȓ*�j���l
�L����Aʉ �̅ȓ!�d��(�7u�	r�/J��`�ȓ(%�����'�^4���
�[���ȓ[�h1���qG<�@	6dbf��S�? ���H�<4�2���`����B"OP8���V�9 �ʵ�rd�c"O��A�Aޥ����A�T�q+"O��J���!|܂UAx	� Ϳ�yB [�(�2�0 �:��TDH�y�H�5G��
a�nY�|���&�yB��`E���pD�*Z
Th3̅=�y�
8� @��̝:\<11b�B��yR��mn�ĐF/Z W�X18����y�`�r�,Q��V(�	�K\#�y"�E.]$J��� �[Ƃqp�ƹ�y�.�.	B��D�G=D�<�8�F���yR�C�-�ԵxV�G��,���Y��y2@Ž6�4T��j_A����C$���y�&�rǦ<��D; `2܀��M%�yb�[*P���"�ϗ�y��Pl��y��S9�Z��R�t�tWN���y�A�<0^~9����o���r��Z��y���\��	h��[W9+V��y�$
��y����8�N `���yB�L�L`B�&H
4<�3�ό��yBlX��o�*O��EI䤘��y2��7p" �Ǡ8` P�#G�0�y2��*s9�����jWQY�\��y�d,+���bi]�gR� 2���yb�G�op���ҧ"M����R�E�y�L���P�5AR�|3���Py�GĎ/.:�0G(_�Z@���]�<ya K�	�`�¨f���b_p�<9���
B���A똠
y�-hc�l�<��i�%E%0�SA5Xz`:��S�<q�G](#��y��D�01^��7�P�<)�� �1b���#m\4F� s�d�<��@O<iJ�)��Θ�^�:��T)�a�<�E1Y���R��]���'��_�<y&#��.��J"�ײ5����n�Q�<aga��c�����gʱ}lV�9�.�S�<�fD�v7F��*�3`锌�!gLI�<A��S��z�±D�qT\a�ÞI�<���1zm��W�U�Xq���^G�<) g� %-<��@��f���1��G�<���~��:�Ɗ���u�  �<�BO�$<�K�`X*[��]�ZA>B�t��g�3~�@Q���%��C�I�a|*���(¶3�ʼ����iyVC�	�< �P��D��H�0z䊞�K]0C�ə3m�ň�E�;I��D1�\O�C�Ɋf��Y�s*��$SN ���L��B�	E��q`��D<D��D)�B�e�����e���1$��o�B�� _�<���^ ұ�g`Ğ*v`B�I)<P|1I���	~Ϧ%8�'���y ^�f+�`�	Fp�D #��y�F�*'`X�x4h�_� �8���yB�G�Y,�l��� ,d}cSO#�y��/�J IB�U�uXl(��Y%�y���3ͮ�+��׊�2�bcߊ�y⤔�/`ډAD��5u
Q�%O[�yb@g=������>5A��HՋ��y��)MR��aK[�>�<�;��$�y2��*�b��0
�cc��`Ņ�y�k�3yۦ�ˇ
R����
��y	����[u& ����>]�~��$$�5jvmͶv4((�%ǹIv����S�? ��P��<i٬�{T(_+�(�@�"O�hP&��5�H���H4d���!"O���B�"^X�h��ݖ{�8��"Ojl����0N��,¡E�7
���[�"O�1)q̊�h�B��)O��Ӈ#^�Ũ�Ba��s���I�.֖�`�
-	Yz ��1D��ʖ(Ok��@B�ߢJ<]�S"�Oh����&�%��Ɍ|	��p&C�*����.�:{���D�Q���aoP����L3����*P�K���@	6�yr�J��|c��JJ�r�y��K�ո';��z���`��"�[��(��4X7�@�Q�c׏��B��N�!�D>[��9�fI�$6j����V����e�߁h��Y
p3O�-K��3?Q-��j����U�X��Bfj�d�<��߭����l�Nz� q�#:c��
�/�$�����M`���W�>z�U���+ �`R�:O
��s��w�pa������jJ�^��{!%̓!1D���"O��`JA5D���i$$��\���/�&yx����^�!K4�jp��M�Ob>Eb�)�\��6�Z��VE��'���ѐ�W�V�}@�MR�k���s*��
F`�#%Y�t�.���Jۿ�ħ�1On �a�6x�͒�M;w�84W�'�E�� ��)Ѓ��(��:���&\~���9#���Q.@��ԅ��^a� �����}�|�J�C%�#>��L�G���{'o�-W"�\�T �#(��D���r���{S��,|(�Lq�<!E.�:��}K�Ƈ)7T�7.�:�y�/]9l���hU��������cG�;§@�q�&Nס_�v��c
=g�d�ȓ�LaoF�~�����2��Q@���p@��,έ$�2� ��Y��OY�ژ'��81q�^/0��� H.g�41
�f�<	2̐��z �
��&h�"]�m���J# ߰��qn�e�j9�ӓ}�ي�AʹK�4A9E��
H4Ez��ȇ=�|�p��L����`��"��p؃�������A&�R��GU.xB�It�r����
'mԑ��4z�V6M��3��
Q�=�H���	��(��Ik��sCn��g܈<��BB+ �f�j�<�!�E<t�������(CVp���#�B�;��J�{~Ʃr���$6�� �O_���s5�.v�ub֤�%QZ��0����$�!V�5m"�	�4?>�W'A8�r���bݳ&Q�H)3��?ss���	>m�N�zQ.B.7@�qS�C���HO~����] �y�5f	�k!l�y�F��Ꙙ� "qN�D��M&0�2a�]c�<��O ��B�O
�(Y�B٦�����^�}jQ� �!��p`�.4���\c��5��hZ[9�H��g(?|���'w�9a%<��\�F`�֊
 �^�U��ٻ,L'l��9�͙���)^bb>㞰!1dT��,`��&R��Q��+�O��+ ��2-���v�-~�(��D�
�A -F�i�0��� ǈ1�B���'�5����ZY�4��!�/�.�C��D�?Dft�e��)J�}�ˇ�	���1z
��Z*@m����#���&C�I4\q����h�Qj�	/�"牧��yZ�J��ΐ��o�5^#~2���2=�E��i8���fǛ�!��%_}���Q)׸I��AP�f��p�@[ê
�\�����'��X�`�<�619��	.�\@��h١$$&b��P��1 Ә��5�"5�h�0O��"@ÈV[�$����4p�"Of����?8�r(;�D	�P/�lҦ"Oz=9g�_�pJz(���B<YL	K�"O���/Ӧ8Ul�iu�M�k�!g"O69֨�:JR=���B�`UEA�"O.��A��Q���Ϊr:���"O�5+-�.��0���DJĊ�"O�@�ӄ�6�Mx��VM�^	�U"O��bq�ލ9h�t�[]q�s�"O�� F��#wz
��W�i���c"O���Ԅ�M{�M���}�;�"O�餀�y�P!�s��f�d�"O±0 DD;G1�%X���@��[!"O,(V�љ�`Id*��{���yF"O̡1��� qTE�ǃs��P�"O� �;q/��,D�$ce�}j$<A�"O.�a���TJ���ė�Xζ!��"O�H�KL/Ti��p�F�L����0"Ot���!�;I�Uk�H�L��5U"O����0`H:d���c&�s!��(IqRHBĦ!)Ҭ�'
���!�dG9�$Ub���r���ć	�!��7D�\�Hē��:q�A�3L�!�D�$G:���D���"W�.+�!�t>��!h3'��T��O !�!�J�i��m�G�"�����0�!��0�Z-� �S
{���A�N�~�!�$���< ���~�@�Q�
�-X!�d�'�b��l�Z��Da逡q]!�$�2o�&%��B֠��i8�cʗf�!��g@B�z� A�n/\���*_�!�>$��x$Ƹ<9&8�bU�X�!�$�&7����!�1��M������!�#!MD�����N����*%!�$ձXUP�:�#����l��o�x!�d��l}3Ck@=p�Bqq�'\�Hr!�΅?]H�(3�ҧUI�E��!t!��7��z�fӆ�0P(@��cc!�O2:l�Ƃ���LBů��^!�DZ�y�¼�k��nHd��.�G!��
P�a�F�ܽk��QQ�3G!���nDu�3A1>�0���.6@!�$~��ti0����01���y
�'Y��� J�@~�PQ�g�	-l!#
�'��u෠ͭRa�����"����
�'��0%� ��W��eP
�'���@�-R<f��92@�]���S	�'�|�(0^!9p%@�Ɏ�@��#�'�r5y��\�8�ቱnϾi�,� 
�'���r��O[
4Kf����WN�<�"+J.v8�	�"�d���ч�H�<�0,;mbPP�ᭁ8z��`c�<���7¡:�쌍>��9��`_�<�e"�qٞ0�1!Wm�<�e�V�<��C�*R,j��G��"&�9��řh�<�AO����� 3��*c]���Q|�<��,ȷA��!�
�Tq���Yb�<قGݩY��i�o��0L��dNd�<�E���%)�E ��[3�"=�"C䉭��a�"�
�m�m��Cb'jB�ɭZ_n��F�]`������FB�ɓm}&)�̉�^��f�K�D�XB�I)��)�qX#�^���	q�`C�I0�}��YO�젳�Ec�4C�I-2e�֥�@U p�$�U��B�
]�X)&E	X��9CӤ04B��qnz1"�M8n
u0��U �&B�I:Y�\�V�E nʈ|����&1�B�ɬ"C�l��&�?03�,��L�Z��C䉬s#J07ݞg:J%F��+��C�ɞ_"xqz1��9!.`CA��l�0B䉋�VpR�|y>(ӒM!�
B�ɿ`a��8�"	S�,+�JZ�1�C�Ʌ_�����NڧR����$WQtC�� $�pT���]CA ��`�]�?��B�ɫz4��Qυ�!࡙�[�B��#��DK'�W�R�^8�$A�aǄB�`N���5.��`�Q#}9!�$��^�*�D�Qb�4��a��"O� >�x��2J�X��F�r�X"O���GƔ\��=�U�ֹ�Ea"O �bb��� ��F»"	�]�w"O�AHviV�r������*"�d�U"Oh5�� .^O�[�&S�K�n�ٵ"OT�r"`^%���4�Q�
�L82�"O"1�P�a���UH�Qi� ��"O`�ZT#��fԈ��W�VKs���"OXȫ��	�d�� y¦�-<Q���"Oh�h%�C�}ب��$�$DY��"OvuA�?v� ���▒9G��G"O����D;T���W�iYJI9�"O���Q�a��q+��7�(�"O��(�nt�B���+[�T5�b"O�ݨr�߀4��|p2�G�gǬ���"O�m� ��cvj�����Wʚe��"O�d0�N�$y=8hu�)��\��"O�h1.�;g&�0a�Z"2�x��R"OЀ:���Q=�H�)H�2���"OP�(�(~�j���GY�(�]["Oh1�I�o�lR��]@�ި��"O$A��K�m��\ش0��"O�y�v`̅'�؁��G�[�6�"�"O�`R��$:AL�+�!�S�L���"O�]Wh�f��Y�f��
���d"OmH�jӧ^ɐ�
�Kǉ`�>ݘ�"O�!��j-l
~��C��m� �"O��x�c��3�^ ʷ�&@z�F"Op-pԨW��v�o˝IF椈!"O�1#�OI(��,���i��"O�xPR�� (�qE��gR`2"O޴���H5u^�)���F�ıB"O���kÏrW����T!@H��{�"O~�"*H\�Z�qA%�Q!�Z$"O�i��
]�&2�)dd�LB�(��"O8�p5k?+
D���	�l ���"O�,��=-h��J5��"ON�{�g4z݈�a�BK"7��Y�"O�����0!hmǏ�3�2�1r"O���V���eՂT{q��$2"O�����?���{�kހFOB�y�"OlhP1��l.���ʝ�+�8�"O|+'�0U\�-I`/,����"Oz�K%cM�&�jA򑍈����"O2P��l�*�@���"O��҂V�|���������6"OR@�W+U>X]pa���P�/�T�@"O�u�ޥ�ԥ�$'G�n�P0@"O8�	�f,i�@4 ��-U�ř�
Oʸ (��*����v-�"�x�`�&�=�~�.G6��'��	��"��'Q���&��+~��!�"cW#)� �� e�?ns���J<���|�A�G�Kd>4�aa�*424Y�&e|�T�#?a����0|z�k׳�:�!�V�=4�� �C8G�t�'zj����ȟ�F�M�Fe>#4ΙDS��±Ǌ
��Dܳ��9�C�U�)�'k\ҵ�W_|b}���G�p���]�z!���i!�S��yb)N.���X��Z�o���kDM�q�P���.��۶*��c�ۤKO�=�������U�Sta�Td��Y�@�#pKO��&,�������]�?�%A��������$˟A�
Pˣ+
��$�r���M�#��@igA<}��i�1[K̔г�Ď+*qcv���3Jt�	�=�J��Q��Y�Og���ħd��b�W'�ޤ��-gJPY2�`��/�|�x��m�vŰ�lI��0|�E�A]��8�dO�h��U�I _���5�m��m+M]��H9ç.Z��Ѳ#�!7ݚ%�cٞ��E�t��2�F![�� r������|֧���[�8���& �RN��s!�K1;��Q��-��m��a\�م�3� (9���_9��M�PjB�,+��;3��3o>���'���Č`�g?�O�NB�KOe[BQ!U�*	5���`�b�&��	�3�
ԣ�*G2����ÈMt�O��� B3�)�IA�w��U�g�v��y2� �>�'��}:����3ƚ����~��.I<O��I�X#6��?E��H31����/[�e%����+�?�C�9��������1"�P�z"L��.b8|���S�+��+��	]�Ot�i%��U�����5���^V!��%�̌p#��+e`��u'��L�!��+��������X�!�d	=B�`!ۉ1ɤu�$J�r�!��V�[3��1��]� v(��䀎D!�ā�q>�Bw �]dYÑEG�?!�$�?A��:p���\�T�ڃb!�$�#pbE���B���Kvcʴ+!�䖠\0N��l�Y����%iJ<V,!�\�m��YYp��<9����!򤘚c���˩J���%G�4G!�R�xF�X� I�C^��!��hS!�d\�a����kX.M>����i�x&!���|�Y �{= ��$��5�!�D:>ɸэ�H5($:C���5!��q��$	�o�'SqD���!�䁴H|.Y�c"�� 4�1���[�!�A�2���5&U=ED !��I&:�!��I+(����dOY�&V����a̚C�!��E'T)H�ɠ�ڞLV��ѡƅ0�!�d	�M�@��G�]�5:�aH�o�4�!��3iL�a��\#*$.4����/�!򤁤I�T����'gҌ��lVlq!���ARCC	�<�Z���GY!����9bT�Q&\�L
ӨJW!����������4֤`kt��6Q!�d4Wt�Z�:9߮����ҏ=<!��38Dv�sp��Q��5�f)T��!�d�gf��x M���	$h�!#�!��:dl�)��O�P�Nl�$%S=r�!�d�z���ࠜ9,��L:�"T?��򤂇"P��R�K�L �a��A��y�(v��%k񉔁{G��R�l�ybKO���y(�.�?&"��Bu��(�yR`�^�X��3e3,Ӿ�D���yR��%:�d �I�mb��È���y�-+%" 3J�h��P�C�y�
��_b�bq�\���|{�#��y�׮J�$�P��|����di��yB� /�p<Iï��l��T`D̏2�ybj�5��!y�̟�,n�d$���y�(е�a�#鐯3]�pl
�yr���gT\y�p�T�yu�0�d��yB����h�U�D�FY�s�܇�y�H#~�L��DbM�4��H�b`��y��ݴ!p�y�3L�9�gF��y�-�/l�r#f��<���0���?�yb���uU�d���߲*q�Eʡ�yhL����rA��h����-B-�y¯R�b �f�B�o�Ȕ�dC���yr�)a���D�~T�4Q��y�͘�p��!q"�)InV��T
�%�yҊ
��Hفq��-G�� 4��y2�DeF���镅A�ݩ����y� PE�$�ڐ�?N&!�cN̈́�yRGIc�����������)�yr��r���+U��jq�Ǫ�y
� ���%d��(�b!���9W"O`IQ���d�����:q���W"O
�ە�ˌk��-�P�@�P�Z"O�@P�m�%v�0�h��EX�"O����ʈ6���bҴj�^�a"O�����Ύ,��l�R�V��^|��"O��H�A�b��I*��6z)����"O*ܣ�,ېLO4%�!�I�JI ��G"O�Q!@u]©�b�/���%"O<��4@2��SA�?&� A�"O (9 �:r��`�@P.���b�"O���D�w�<[�.�o��10P"O<���.T?4�bU;��I�s��b1"OF�9di�=@��m��	 ��i�"O��K��,.��#������K�"OvpV��C���9�iC���"O.�g��C��|!B�
�'s��;�"Op�B$%#b�k&S4�S"O�$��E�;Yj�%�2���"O��`�ڞ��sD�9SF%i"O�D��i�i�JA�!D��q�0d�`"OR�a�,B'h�|̡��
+���E"O	�a�q�!AE�8c�쪓"O��F�܇YV���R#Vc��R�"OJ����~1*����^�fjZy{!"Oʹ���" ܨ7aA&����t"O��%e��7- 8�v/�Aj� "OHia���m�N���jLX�k�"O�R��܌V5V�
tN��\1X��"O"\���L%���Ԯ�!+��a�"O*@�p�C�q�����F)�l2D���e�{!b����
�C��%D���&��j����X
s\�I�8D�t�V��D��ey��I�p��+,D�T*@%Y�B���'�F m�^-a'+D��ˀ��"E��iD�q4.eZ�*D�<�"��=$���C�Bd6��ʷ$&D���'ʭr��Q{ǊA�Fu���4�$D����e��3�t��ç66cʅ �$%D�p�%R�
�8��&��#ӠA��(D���A�8��͊�;7�( /2D�8�5!S�Tׄ�k2��~^!���.D�T�v�F!l�u���,S�F9 O+D�p�Q� �y?�){D茅?h2�A�*D�$q��T&Te!�ʍ (����&D����I�#F�}(Q�J�i��(�M9D�<2�aMo2�����G'4��I*D� ���0ec<�3�	 �*!c��,D���[)�r�˅�`I>!�re>D��PTG 	2���Q#�<�k@`<D�d�g�� NQ�MT���X�!<D��y�@�&W�8�ǀO��1X�$;D�4��j��m��X[lϑ2{n����7D����$e�,�B��Ȗs�nY��#;D�����2_�(@n� u��E+D�hT'��l����&� 6����	+D�L��A�y����jǉX/^��d$D�h�'S9	��ۡhĠF���{4�#D��B�L�l�hU�\�@�	S�.D�̫�ɓ�^��t��\�!Ql]X�*O4��V�|@bŮ(sR��3"O���Q�p�4��W���5"Oth�#,X t� ǎvu�Q"Oz-jdKE;~ �&^�Q�H��w"O� �M`p�@b�l�`��0
�h%�u"Ox\#��J�S@�e��F�^Q�u��"O�����o�&�q'&�3��YW"O��kW-	4���p儥`O�M�Q"O6����ŚQ�hsF�67���"Ot��� �t8ѓ%�"BTv�h�"O��;"h���M�7��%/T�1j�"O��ペ�ss�����ЭGI�dB�"O`YAD��:n���Wc�W>N���"O\d��kɝ ĺ�*��6�EF2D��:D��oGDP�� �]���S�I/D� �ƏQ$�`���<S�Nt�$-D�؀���(	
��xW�V�FAN4�w!D�p�T�Kj�4�*Ӓ�0�c'I;D�4�3��S`�p�#.�(R��qp&�#D�N� =@k�$+s��S&D�:G�*B�'�	7$S� ���i��H��C�ɫ.*��ِ�G�U��l@�'�*v<�B�ɼT�p y�5z��H��P?YwjB�*�L����[mEx�H¦�u?6B�I�e�$�q�*E�)0L�����Ӎ��P,��j�"?�N\B�E�1�����Ĉ��eO���ؙQO7�@��L�\Y�f]pI�=�V/TE'� ���hbB��>/��}�*ܾ|~ A��q�,!b�ʞb�֜�r��:"e�ȓWtX�Eӕ+���aN�Eq����{]�ŹS,��=p+�'�9m�,Q�ȓ*]T5�ʺ�4 �5M�9�ȓu̍Z�AW�}gh�����gDzE�ȓf�����e�W�H��S0;@���t�B�HviO�,j��:��� ��Շ�'��:I�8���X�ĺBD�ȓv��$aׯM4.��� �+E��d�ȓ�)���4W��Up�N8��̄ȓ�Z�0��P 2XPeJ��5�ȓI�
���E�/��K��J�(ҞL�ȓZ������TZ�!����=y�@�ȓjb��k��G��F1Zl�� 0z$��b���BS�W;��J� �]s�<�ȓj�*���
D�\���D�V��]��/�E�Bߵe��y0�]�WG"�ȓd��s��º8,vu`%+\4A�&�ȓ/eL�8r�[��L�k�l�����'��Q�b� 2,��E�v�|���'&�<��J�	@L
v-G�:��|`
�'�L�Jeg�*�	jr�ֳ4�� ��'��T!�(ԡ,L�Hr&K��X�'��� �-)�ygaZ;��H�'`��v:�taejH�c�b �'F	*B��^����L
c-�X��'N�A�k�5Ċ�aY%UEnu9�'�&��PE�&K��h	�uV�)��'��l"���TM ��`�
q��$��'x�)V�*��hK��`�j��"O�xp��^��d� a҆b-R �"O����
��� � F�AyV�0=!���z� �pJH$	U���3��8!�䝣#�K� ҌD��tB�b!�d�q'Xp2���E�X�cv��\�!�$ɶ]P�R��$N�3ҧk�!�DD4!JԩRQ߷2)��'%��zl!��ЍN\򣊀JB���#ģ,�!�$�~ �P٢�Z%H��a\ �!�� ��bB�I,[���b��[d"OL�Al�:c�m8TH/K �"O���fBh�Y(�7.��#�"O�$�����&>���f�(~2��Y�"O8DP�AU�D�>��3Ő!N$�t"O6�`g�ѩo��j�Ŗ[I�a�"Oȼ#A��ڮ�	B�V2: `�`"O��ق�)�����N�Ƀ"OL,@�h��3vܼ9�C5#u*�(�"O�]*�F�NA�C`��*W�	v"O0�PpI]�`Pt��J	 B:&�`R"O��J�)U���гÉ�=P4��"O����:V���	aÈ-�0�q"Orl��
�Q"P��VAf����g"OFQ��ʀ�����/�h`I���O2R'�/�M+ϓ�M0J��f��@FJ�C��Y:X�;�(�U��7D&�R�.�%wN� j�*\�.}	�r��1��a�G^0_g��37�W���P�I�{,��D��B��!JXw��	� ���'��|x�^�$�4O	�:
.lJߴ�j�4!��`%�h&Eۂj���z#$���
%!0}��'w��O�9��Ãh��-���tG�Ӧu%���ݴ�.O�]S���am�52�^]-��M�T��;PZF(��/O:�䓙
��Ѹ�⑏
���z��D�-�DH��"۽�} ��%Ր��RlI�,Zy"c�ɷ	���hs�[�H��C��|!�h��fY����)LY�ͣ��[�C�����	��'7�@������eX��KC/ž m�-Q�!۞P^ұ�O��$�O>�O�˧��D˅*n�l����7=`���,ғa2!�dUl;����]� <HQP�l��0#V�i޴S6�F�'Ҷ7mA�;��o���'A�\�vءf@Пa&��BW"؎ֲD�s?}��'"6� ��D'�����
?c��{�$׍�\���ZU�)`o��NU���#Щ#��$�>a�l� ���q��1��Ḱ,I�@�L4�`"XϺ{�OW'hˈ���)$���
�GLE�'��	�ɟ�M�i�"���h4}�b���75����%F�|��˓���O>�iz�(r	N�<���s�L*0>pu��I즁�۴������^�	FL��F��4mW4%l8X���-+ɛv�'�i>!��\�^�Bu��Rt����ڒ^�����}��HV�i���Z���"�[f�?u�S�D+�.�rK��9s�-��d��eh�}Z�J9M����p<l�)h��ܠ)xr��U�^��Hcޙ�q."U��|x �K[�^d��L���?�7�i�ʓe��D���߹q%�۲�Vm�QfO5n�8���L��?��D�<�Н>��+��D����
�m{�9 CO~ܓ8қ�Ck�v����5���?������a'm�$wX4�6��_,�0*���d����M�	ϓ�MK�HCYh��䉑(�Ȩ;c�ҿ.p��8��\��Y��ς:(��K�B�s-�A��B���lt4q���4F�ѳK�P`��S� ;5H�	O	�""`ݱ�e'����c�((���s��f��)$��"r�pQ��',N7-{�	�����T��)Z�2$H�Q�6�r����&���'%�yS��5��`8�Ë�LenȰS"
�]$�4h޴��*O�đ1�E��oچ%�����?$ܠ!��E�Cwt���O��1p�J��Д��kφTpU��
�vPPp�çC%b�Ce��W�J��S�I�2�Q��P���p�a�Im�0M�C���$���e۾@麬�T�^�?q�aqG�'1Q�y��O�m�7U��a�BU�sf�%�UI��&~~�ޟ��'����?�m�5F}4�ѐß,$v�)r��!��B���՘עR�t��"S� ����G�P11���|��`ݍ�IN�I���#�O   ��   �  }  �  W  �'  �0  �7  *>  }D  �J  Q  IW  �]  �c  j  Vp  �v  �|  �  a�  ��  �  *�  m�  ��  �  ��  ��  Z�  �  K�  {�  !�  d�  ��  D�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ��N~��\	?Cv@ӎҿF��(8`����y�DG�|�mYDG1E�>-��'��y"	�*]�MYԤG,Czr��v���y�M��ۗU�~L�S�Q���(O�pD{��D�� o ���G̿%�v�K#�^��y2'�q�
�1N	�%uJ%Qq���y�ԆE��,F��H���[�y"�C�@�h&��5F��8wFU4�yb���B��|�g�Q{I� �&.Ҡ�y�a�3���C�'Ǩv���p�7�y2�" =��9��H�vVXt��kA�w�t˓��S��?i0A�x6n�ڡ��L���˶�t�<ѕ�צ2(=����j��{Ro{�<yF7BX"ɓ6*��P���Ã�Ju��'���%�B)ct��և
?��q��>D���%,]>d�h���K�S�z5���1D����`@����yge5R��P��,D�,�a��Q,�|KAI�
Ԏ��a�+D��c�����0
 e��0�|9�4B,D�Lx�U��� iL]LifQ�@}�
��'��|r��=z�t3�e�rC,�Д����y�#Ɔ_��,�!eO�ky��2�G��y��Ӓ0j����֘jЎ	h�/˘'�ўb>� mI���"��M�'� �o��'"O���U͉�P A�sFQ
0��!�"O@�B�¾?l~�ѷ�ΝpƂ�l4D�h�P�K�:B�`�e�$"*�
%D�\ɐ��y{�yc�F���M�H$LO��{�{��C�R��x�"�"D�|�y3
[��y/C-�n�Z��ȱ<M�9��+	%�yjE�R�e� ��Q���K~F�C�-,���7��>f�y����3H�C�I>�0��A�W!���'�A�A�LC�I(B��r
�.Ml�+d���P�X7M1���҉@�0�Lqɇj�0:��%��'(D����оPX���G�@���:&*%D�� "$�v*���#K6���e�.D�|�֧YM'Ĝ���J�x�,�(�H!D���F��p�@�h�u�2��W�?D��"�)/˶(S҂ܩL�52?D� ��DT�l��c��4�J	h�:D��X��W0\�l"��5��8�@6D��p�Y�\fp��7=ƺ��'D�,��,G.��� �_4;�h�Cv"8D���`қ1�D��1��m�Vr�M7D�HBwf�u�\ �[�^�dy�ƶ� �
�U��Q�5l��kf�j��t��W�`� 6��{s0T�6����⩄ȓ=�����"HغT�R�6�X��G;���c/H?52�*�%<;��L�ȓ!$l
g���p"���.@��	v����6% "��OŶ�$��`�f�!�+'D��5��2H��)��B�L�怣<�'�.}�U��&?�������!CG�W��D�R�C��C䉱]��Cď\�a��U)P%l��O����G�U�������;��Q�re��7��z�d�9I������8�	�dJ�K�!�\2y
�PB�O�U̤Q�����'��D)�)�S+��!�i�(X�܈��d֫w"C�ɺ:g:���	� ?��Q�ĆF���L��'U?j���
x��	
�ÝI�����(��T�2��8`�V��� ���{Y!�$�;R�d�/P�l�@�2SD��$3Q�,D{*���mCX��y4j�17x���HH<�$kԒW��6&�$.x0��|�<��G�:4Lm�T���PC�3�h��<Y�ϵ"L,�`Ҁ
F `cfH[x��p=	��yW�U��)U.q��I][�<A� ��yDA��D�I�`,�LLY�<�L�"
mN$Z�K��%��)jf��R�<a�ɚ��i;�d��X{H1J�g�V�<�C�V��h�ǩ�O��h�WP�<	c�2a�p35dU�8�4��H�<���X����0ݳW�Pܓ�M�ϓ0dx�Ч��1�V�I� V;ڤ�ȓ{ez���Ö�uVH�R�H�/��ćȓ#X�r�ʋ�W]zcܢ����M�ȸ�T!@�#����Q+���)�`B���f���.Z�6��a�'�YFy�𩃣E~�;p��S}h�f�Z!����)�wӳmV�Y�a�!�P�xk��"�P
��$�"-]�Y�!��q���I ���3b,�%|�:��ȓo�4�8��NP8�@@ c��t���f��6(��jP��X�Eܴ�ȓ��j�M5sn2i�II�$��a�he�`�W&}�R��e�O�܅�S�? b���H0��q�$�7I>9;�"O�Tb��ۨ,�D��;�N���"O�TC'��by� -<����q"O���)F�����,
�{v*�Z4"O��:㋦o�ja�d
<pf\T��"OZ��V��Frġ��K�O�\��"O ����W��8�é J��p�"O�<⶯B24UZ7O�i����'�I�R��x"D�2Y�(SN��x���&���yң�x���(^m��(�a�_��u�8�8�I�Þ��g
\XW!���*X�\����:���z7G&rn!�Ow��ĚF�=+���ӕ��(�O��=%>���Nɪx�����!D�!�:D�x[U�>s^A����.ZǤM�be&D�L[�.��B���� �D�8AdK�n&D��a%���j��X��+vu�y���#D��2p�@�Jۅ�;ռQ�A�!�y"a�� �J�B�3�X�ж��+�y��ܠ�B��O�$�ZUQV���y+A:/$�5@�H͹�qQPD���yr�ŏ;b�i�%���0Qh�8�y������W�T�s�j��IT��y�l�9�q���W�f���!�L;�yMX'(��\�G�$�:�&��yR��� D4cC����az����yr��;Zd"݌U���Հˁ�y���+�XH�E��I>晘Uŉ��y2��WM����

oӢ���n���yb�ЩX��(�0m�QH��bUJV��y�!ֆs�V;��*ۘU����yҍ=zE� !a�7K�����O>�y�9ܾ\����:pN��x���5�yB��'uS�@J�F;cFd �ea�4�yC]>�T)�k�(��)�q���y��ZY��A��a�����,��y�_�۸���̑4,���p����y2� �&�`���3� �7#��y� e;��$ȃ�
=$���!ڀ�yB�Z�u�l�p䒊�^r@J���y�L�:-��q��T�q���'*[��y"��7U�$���Au��Bn���y��2Pe��`��qȸ�v���y�撺)���K�pX��6*��y��VU��q�Ҧn4��q��y����-
!]�es���0j_;�yr�ɣG^E�`�O�p�52Ǎ�%�yE��'�D�C�셹W�ԑ��
��yE��'^��}�U�UkA��y"b�x�|�A���LX5Ċ��y�a���H���~j2� B�yR �$ln�дG6t����FD�yRBD�C��e�v,��ã�ʋ�yr"G�%���[�M�h�T���T �yR�ī>�������j���h �yR�7���h��g ԟ�y�D�P7A�(Y�
�+A`��X�'X�k�@��|����T*�>j�t[�'���K���6`vi�A�Cgm
���'/��H�bO� ���"Z�l�lѣ�'�Ȉ0#M�w���0�@�V0�0�'~��cFmFV�JɒSz&�3�'I:q���m���ؑ��G����'m���̙c���ʄo�>�<	��� r���^�k/i�c�ڶj�f�;�"OV���. ?��ɕ�۪:�jT"O2�!�g�� ��92���	$$��s"O�L8p�u�����l1���2"O�%C���\a��̴)�)��'�r�'.B�'F�'���'�B�'�fU�'�O{��P��[��1+F�'�r�''��'E��'���'��'��1����*��dCأD�⠢�'��'b�'�2�o�������X��!�l��r���2NT�3�ӟ ���0�I��,�IӟD�I��8��џ�`�� /�Qj��J?n= 1�mʟ��I���I��Iޟ������ȟȩ�ݦ���RbE�7����I͟�	�D�����I����	ן���ϟ(""�B���2Ŕ{�~����$��Ο��I�T�	ӟ��	۟��	�� �Z�@:��k�@�$���!��(�������������ߟ$�I��Ĩ����SE/#����afFҟ��Iǟ��	ȟ8��ΟX��ޟ���П� V�F�v��9Eh�z�tԘ����h��ğ$�	̟����`�	џ��I�PR'��k6F�kA�E�t����nY������������	�@��ӟ4����2e��1b���6�	!��E(5�ٟ��ڟ|�	ş��	����l�I۟,���(6I^Ve�Ǡ�z�Dߟ|��ߟ�����������I��M����?�"�6SF��g�����:�*[)����\�����ĆȦ���ӈkkJ��f�ZO
a饠�]u<�;����4����!SO�H���{o�JR��M���=���ݴ���K�=T�YrBG<���&o7��;��iM`�9�쟜b2Bb����\y��#CGQ�g˰o�)��]�c5@��4�d�<y���(y��&�H�(�`
(~��]�6���en�M3�'��)擏B	|�lZ�<�B�������媵�qn��<	�!�A�.(81�P��hO��O���@Lɍ8�T�3���0�x��6O����*d�������'}���E�B��⁅G�ph���m}�icӠoZ�<��O�����>bЅD�N%2�j�g��b��K��"T�5擪N�;V�e���@j��	��� K��Iiy�𧈟�R�_z���c
f`�"�J$&{�D�̦AaK,?���i#�O�)�-,��	��Hz��ҋpt�Ц��ڴ�?	���M��O�Hz�݉u�HS�B�s6>�ѵ�)d�t`��vY!��ޛ���e�+d�F���ޝQ�!�[�x����H2�6=�u�ɋU����g)�	.��h�p��&R̸ۤŪ�9w�Z(��ꊻ�f����́A��-��O�%�Z#͕*T� Mr���O���/K,(��#f��!������B���t�Ȟ<�u��D�6�F��Q쁱:�u�U"3=��D{�@�4>�v�0�Q�b_4�:�MF�hw��ϓ;����a+�d�8l�#�W����PE]�7�ہʌ-;���(M�d![��Qz��U`aJڷ9�b�24��_eD��v+_�܍{��"Y����V���˔9=,���s�ڋ�tу2g�#:Ք)���ؾ6�ͨ��8"_~��Ο/����߁ �1C�d�-r^<Lـ$�"?�\�Cd��k0| cdB̋,6>(���Q���?	���?YtV?M���v9T����n�*��1��"��҅���N3���-�2� 1��?u�RkN�Z�1O�I�C�;T� �1��K�<� �oX! �Ru�#�D��֌��v���1sx�}�&
�-Rr��R��q��;o���*�+F#���#�a�L����s��nz��Y���	qy"�z���e�_,kX�{�k���xB�'O �X�R����0f��a�h�=��������&�DlZ4W|��ӯ�D�|��� �z|x������P��a������|�&#Ls8�re�bd2$���0^��V/� ��YU ���i��m�+/�4}Dy���qxr�� 0w�I�5c�(x����W��y���M�������*׆2�O���'� 6�
 zF���@�!�U:����j��i��Y�|�	N�S����`V
x[ M�z���C�O���0<�����
1�HX'�	h ��w���W��^����`y�����'�?Q.�.��
V���#���ϼ3�l f����OL�������LF�mJ���')�VC��L�Q�	I�0=
T�܁�d�r�LL�f�Q��s�J��5o�)�$�{��@�Q�rE��uQi�F��u���^nȀs���J�Oƌs��'�N7�y�'Ӷq �]&y��|뷊׬"��?����]CF�^�,1��]�QJd�'�ў��1��j�Ti��1GA�!ۥ�۵	���X�FMj�U���Ie��@��b���'�q�Y7J��K���y��ިB���8�h��YՊ���͑�gH0	���M����v�e�� \�\�D�p!�Dڈ�C�+y��rF	�9	c�&D+r2�F���/N�Q@M�$������C�,���d�?��i�7��O�"~�	�c$Y�"�>�ʰb��E���I����	x�����$A|�@4BR5�#<�����?��	m�Nh F��,HZ��gۯ�����ʟ���&���U����?����?��r���O��I��B��@'n���B��P����#��]�S��8)@�H�5��I�6�� �yf�1~�r�sAC��q��dy7�πzj�B4��-,��s�A�^V,��O�m���h�S�? L�#F�:^�&�H�IT�EP�)ʠ�O����'���|��'��_��Q�n���Vt0%j�j����1�'D��:6ʈ#)�p�	3��4*��`�,F�HO���O�����e�i�Z��Յ]�eC��jC:����'w��'dң�"���'^R��!)Z�e�BhIX��ECV���aH��@�5<�
�s��W/t�Ԕ��Fz{�ᲈ��;����ӳF ��Ç��P��e��'8@�E��$K�8-Ո��vq����<;R�'5�u@���n*�ȹ��J�j���M������U��}�Z��J�AB�� ++J��L� �S/j�!�_�� �6�P}�Ġ���d���Φ]�ش���>\�N�l�՟��m��N�|#�1��ٚW�d@Y��T�����'�b�'�h��fȔ4jA���o��G��pAo�d�FE��T�T�˲ L�ΉicV4�(O�ɂ�D��!���E\�-@��Z�`*2�0�D]��,��e��R~Y��,�1Q���VN'��F1PR�g�Խ�~:`�����A _>.R��iŭ�<I���>#d�#"L�!��P;
�h�z~"�i>�O<yTn�?)�B�h@�:,[4ѹ�eJy̓�?��V.&�bg٨� usC�Q_ڈ�ȓs��D��)G�	����J�Lj�M��N���`E�%}`��� ؟
b�}�ȓ88��2B�Z�u�fdZ�G� {Tl�ȓ0�pd��?RډX�� s2�|�ȓ ��(����'D���IK�sO�ȓA����fD�XT�@����v����P`Ĥ�� Ύb��Aؔ��?��%��BD��3�,��,�C���|u	�ȓ_���k�.T�
[���E���PU���U!X�YYԔ��Q.�k����R"O�2���6������&겄�5"OJ�3�l�Kg�}kC�Eޮ<�"O� �
H��p�u���Ќe�g"O����-��J� ~��dp"O���U	N-qa�0{��@�`����"O�<�4��9;�P8AC��%A8�q�"O�x@��Y�W���ѣ��)&أ"O�Q*�G����Fթq���;&"O��X��|��9�dl��o���@"O�90���(S
�	p��.�����"O�L�bn�{"��#�gQ�T|���"OP���i���֘�� hV\h2"OJ�2��P�:��7o@13�Y��"O
]�d҇|%Z<�B�ȾW"H�yD"Ol���"W�w��u;�9�(1��"O�ir%�Ͱa�� ���[�� �A�"OH}*����1� q��Yj#"O�0��N0I�PSǢ�]պ��"O,�y��I�FIN�b	 7(dW�'Q�oӡq��t��OķvF4bSn&D��Y�
i\�i{a&�/J����a�<٣啹P?�OQ>���'L1o/����-C1m���5�)D�T��
0j9th�d@�-\����#�4�Đ�8(���'©��E�*|�{2�K(W�Bh�	��P�d
��_�{�ș2�Γe>\!��x�:��c��	3Y�=��I�7
��H3J@�C�����">��V�A�`B�!�H�pY?	�����8��[�)�0fX6�)D��"3
B�U҄kF��]���QD't��U-]�&$�-��<�B� 7���Il�}�b,Ý}a�Dss�*|��B�!5�:�Z�Z�_�He[iY���P7�S�U;����D�U�du$,Fx�A�,%L� H��H�O~h"�F����>!�N��l��P��8��h�CM6>��=�2oɪ)op��琭f��e��l�"a�Ęg��hCFE�&��\Gz��ʩN6n�2Vj�� �&d���M�'1��R�a�A^l��p��Is���2��)�NL�v*a�V}��_��-YW썸@mTB���f��.�d7�s��Z�g��/Zq	͎-�\�0
,D���ရ?���1�m�6A�J��v#�i���G��>#_�l��D)���g�'RFyk�#�$o�|�i�AO
X���
�GC�}�6�Ks�? ��0����
�L��n�M9t�6$L/3�
M�d�DMX�Xꕁ*O>�rs��(@@D�N(�=2qC��נ���c���S3�r���]�p"c��#�ZB�	�#�mzt��Q�%���ABb�ɆǾQ*�N";J�# ���ȟ��yq,�,r�Kd��6>�4	Z"O���e*	(E��R&�}��t�Ԭ�&��lځ��ų�GB�n��g�'%* �����Pκ�bF��((�d	
�T��+U	ؼhE�Q6
� 	�Μ��
�}����R,�8%# �t�'�8�W��9ȞAC5��5"�V�Q��$�3'u�0c�((Fq�B̨|�W�ҨȢMȢs��H�O�<i�ŤO�h��E�UH�����L�@	�Mܴ�[��hy��i5'����w�z>�L����pL�C䉑tA��!����"��D�P�z�|�w�y��
�1Ǔ?��Xs7�D?G������7�1���6��xa�i�����jax��C�[cޢh��"O�|��b�&B-;�r�����>�{C�S�.l�$�u͘�:7ⱺ X)>�C�	�nnZ��
wS����.B�F&�6�]�9�4�"~n�����!瑶[r�b�Q��B�I�)z�i�Iöjh�����I������TAg�'��!�*4,z��䌕$�M��	��8�6��O���&���	����	؊<����"O� ٦OF�B�R:�Îfڨ�鉞 �m�#�"ҧqx����1�� rk�(31����{��Eáɳ4B�p��u�xm��(�t {�N�v�)�����˧Pm�X"�^�[yH��`*O@���&���S�׋Z��)�_�� F��j��I�ua�L�WD9I����F�&���$OPe�I\��	G/�v~񛖫��4ܸ�+'� �v�!��\�l��-ڃ��5a�l$�n��}A�I�+B��J�O�p(�`r�O�"�b�ӆ�(�x�7�@��'����E��;�F@(aM�t�M{�Oܻ2
R)��A��g�M�r���.��x�0��m������lr�	�.�3tyP���	�WyKP� i�	>{.�5"
ӓu���rU�C�Q�.��jلd�ቋr�ڍ�(O�˴F���4��Y���Cԩ�%`H�'��L�4ӿ���bR�T9*"�ON0s���I~2�0V#|���(��(���%�>MzE�y�<�����6�0c��ct(�y}�)ǠY��=�$�'��c>�D����̮;��3�#�.�tH�䯇�7!��܎F�~���1���P��(>L��iT��u1��w�i���ɟ�O �!��-�ąK��]EL��K4�'��i!&�<�`�q�>ɢg�(��U���� `�<D�&A�:�>q�V�J���|r�%j�����.���b������D�P����'��Y�����#O���Χf� a�@�E�0q�*F���ȓdW�MH��u���E��� �HvˤT� 9R���<i�*�O�S*��Ͽ+fFI�e��Aap� 2ņ���LF؟h�TĜ�.\��`ƍ��� JV0h(��4��$H�]d@���-%��1�;s�ĹFx�
P/M�Ԙ0T��[�B�R�K���Ozhx�Δ�
��$�k��`�6�x3M��4$�aJ���?0Y)�bS�wS-HG��za|#ۛD�t	P2���7.$AA$��6��D��Y�L�s�q��Њ��]�*:�h�4���`gD�,-�a�$��/h�zs"O�LQ�#��.�`"�jVK�����4u���V���	E-~��'(f���4���	�Y���@�a�e�TQ�cΰ}_a���3h3l����]*�`3�A�R����Ц��l���I
Z}��',;T-Gx�KÈ,0F���hL�h��t�0"����OFe�5ʗ�<�äQ����U猿;�xPp6,��:��?������I������&.��s*��Q���o6pSa0O֍0��D��<ͧ`SH���P��ư��JZ�J�F���x���3(���#EJ�C�|���:y3��
�zҤ�;����g�i�aQEݥ$p�[�GK������m)�O�,æ&�o��]!#�5�)�ٟ������<QW����/����sD@�46T:㮆�&ޔ��t� �c�ҥ���97��5���D���^��][Æ[�R6P���\��	�p%a|
� ���!�:�J�2�A
�H,� rS���Q�M҈�Bfi�[��#|"�O�`!H���00*r�[Ղ9LN��	�'����vωt���$u���x�[(,w��I�m�@PӇ����g��EK�EϐH�9s����RɄ��,�M�2��fcP�9����n�+A�ݺ"S�`j2U��X��Dɠa�L��	@�y�ŋ!�P;/"a{2(_�8�$h��O`������#F-)<� @"O�`�HB)����ct��M����)�T$
�F!�'1
0��;K�IX f2���ȓ<�2�х�c*��TI�%�v��%�?��'�F��'�z ��bMv�$�)�H�w�8p�
�'"�T�V!�07�u�S�B�d)�ش
\*%�N�a|�k]%g��T	q@Y�B�l13F���=�R��&F(]�w5O|<X4�Ҍ/T�ʆ��A��p"O��"�B�w;�;@��#uB�2���^(�2<AA`5�BHd!�5B����b�B�$%*��ȓ#Y8��e��	�ҽz�o�>�p�l�2>,ء�}���i��m�1�/}t;`��ob�� �'p�Y*���p������/qWt�@�O~��ѧGD��ʧ�1+~�j�e��"�� !�O
lQ�<�6�C8K�~=b�엡n��|b��}�<��Ϙ�[�"�:¬G4T�@H�d�'j&|�a� �.�y�K�7��	�a
\�s[�L�ȓiӰ@Cd��&��zgOA;V��n�B�����s�|�16�ë��h2>��/D��b����<B���$�,�ԥ�>���	�_�$%���3$��F�Ϲf�ي��I�!3���dճB��]z��iI ���+)�,t+���H�z�k
�'3��ZE���Z*�� r⍨>!��ۉ�dξyԬ���)X�O����^9K-vE�e@z2!�D Pd���#ƥVy�ܫ�d�"����<��c�"~nZ2����ۥl�z���!�%yjrC��}R�i6�Ьh�IH��,T�YE�D�p�'��xp����8�cY%V���r	�
l�L��>O$a���[�	�y�
�d�@=Ag"O" :�i�Vo��&C�, ɠ�9��1ѐ��iCJpֈ��*�����Kb�'�!�#-K�|��E?p��ݛ��a���m٬/\c�"~n��v�\��-ܷ$W ��ǅ�5X�&C�IO� [t��.*ޱ���>k˓z䩇�I�sp܁Z�ʂFS��	ш�-��B�9E��Ds�M����
"��!��B�=\[��z�MʀE�8ѳ&�*:��B�I<ix̥2@���ExA���f�lC�ɸa�lJC	ʹe9�Q����/7ZC䉻aG�-�'�Ş��uz�I�ItB�.Җ=9'���v�����kd�C��0W$�!1d�Gn���04�@ 2r�C��;UP���
ޫ&'r���J��C�	|8 �]<���y@ �-e�B��>�M�s�T�~&��#�܉NC�	��D8��� ��$�Ċ�*N(B�	�Q�N�rdc��/����G��X�XB䉊"\�ҳ�J'MȰ� nʁ"�dB�C���@!�8<�� �"�9w�FB�ɐ2�ę��"A/����A牛w�ZB䉜*n\1���FH� 
�[HB�I.#�B���w���QGE�:B�	�5�iÄ�M(JV����T!�B��Qܰ͹sKVkrP�T�?^�HC䉦xF���͙�d�\pkwE�i
C䉙GV��we��)�|��q�;!�B䉖yH�a�VkR;2 쀲�ë �dB�ɝ��dz7`�0(Z��fA�a�\B�)� :����1y�-�WoI�p|��"O(�Y��>,I�Xp���|��`;�"O��C�Oܢ:����⯀�F����P"O��Q� #K�����-R�q��"O�%��N	�1�ⱑK�$5Aj���"O&B儏�Y�D�q�LP&DF÷"O�L���#��d`�,�Ƹ���"O��-E*@N�B�L@�F���"O�T�@���X�$ey�k�1�B�*R"O����J���K�:q��r"O��1��vB���-��u0D���ע�3�Z���,�d��0D�,���	���a��A(k|��� D��	�)�98��*#�ʘ h�L��3D����d�P<����-f���)bh0D�ܰpA�9!4$�d*Z�o|ʰ��`"D�D�2M��H����}�8��=D��P�o]�$#��Bª4u��A��6D�(��*��x�֩c%�2`�~S'�)D��p��ì*`���锗/(B����#D��f*FCb�����ӞA���I�"D� ) �ՏT�8R����
�S4� D��!Viϲȶ��%�̴~����S�<D��ʴG(	� �削�þD�CN/D������>�6���O ����f�.D�����M$���˓�@*pY�� ��-D�L��h�E�ᛔ��S?�)�d(D����NT�mZ��#'��
r�l�RP0D���6���8�F���2z�Vx��!D���qЕibĕ*R`��ewT�Í!D�Ȩ2�נ
vfI�����8�J��p�$D��Z�kJ�������SnX�c
$D�8�Pb\�C{0�A���T7>�� #D��z"F� B)�p&�[/=p�K!D�P
@L���P2�,�,d� x#h1D�|�E��?�>I�UȀ�/��SV.D�  �� ml$i��Z*,.$i)�*Oj@#W@�	pW�L�B�[Y|���"O�!�Rk݄d�qق(�&
{5a�"ORT��)�p�h]Ƞ�O�z�2A"Ob!��S�V� ���F�5c�!"Ops�)�U��X��O�vC���&"O A�@��!�$�(w�ߓo&�LB�"O�TB`���}��K�R!0��"Ol�8��r�V�1��эod��"O>��s!YE!.�1�c��g��"O��з��0�bȨCYSZ0�j�"O8p�hC�T���т�
I]<��"O�92�@J�)��d�-Ax���"OJ���^$^tx� c�_*	�"O�x3��B�A���y�7PhL�"O�`
vk�r��xd�P9r08��"O>D`�Q�D�G��#S
(K"OP�qՁ� ~ߘ����y�ĝS�"O�"�C�-Wl�*S��4P��"O�����4~�t$��O�<��\ �"OX���?;�-� l
�0�vmq�"OH�rM	�hf|%�d�G�a����R�xR�)�ӋZ��U�.n yɣ�߁+�C�?E2�|�s�L6f�	�r��)X9C�I�-��i@�P�:쪤���N�MU�B�	<X GoU�I|.�:��ʾWLB��O�v��C���ΕB�B�2x*B�	_�Z�r�
��h@S�eM�C�)� �]b�p!�P�R���u�ms�"O�����c0���c�@��֤3�"O��)�@�>��%0�����"O�бABD� J<�qu��$6�6�(�"O��c��=P�i�@N�S.�к"O�L�L�u��ҷ��rV*��'��� ㅘ�p4X�/W.X4� �dJ.D�Hj�Z,"쐤�p+.Y�����+D�Ph7��4F X�y$�O��P�+D�1b�ʋb �!囌%r��+�=D�@Ic� s�:CX�3Z`I"�L;D��CԈM0<�fX��e��)�x���9D�h
o A�8��G	?"Z���!D��h���']b�Qh��6�L�'�!��$'�T#p�Ŕ��`B���c!�$��<��Q�0�³4��Dä�<z!�d^�qE��{���
lŐASDƮr<!�d�?z$I"�����+��r3!�$IbX��M�`�H&
�%&!�ė!�� rksfy�
�6no!�$L�^��9ƨ�
������'B!���^�<#ǧ�/��% �iJ1�!��Z��4I�D�*���8�!��
�<- �(O�<p~T��čB�!�d.
b��K Y�m^@l!�g�"�!�DЂc�����n8B�J�Ɵ�q�!�dR�\�`c��u+�U[VǽE !�$F
7��9Y�e� <v�3��,!�$	`e�����E�U*j<�a,Ȓ`!�&̄�`��M&-FLS��^!�$��`0����F�\�ɹ���)x�!��(8�n��^ ���7�!�A�"��m� Р�-���D:@�!�$ F��P���4?���Z��J�D!�� )h�`c�x���R�ꝼ~�!�d�K��XC�E�V�F��Ê׭2!�$��'���kcS7I�fTX�i˽p�!�d�}�����x�ԑ0h�CT!��;: �15*�t��I��ᑛt?�y��I�.q�����V�c�N�>\�ZB�	�m��µ�;1�jQ*�[��HB䉈 ��B�9#�`��E�)M\C�	[;Jhj�f�� �v*T�_��B�I#j�.y��'�p����Q&os�C䉌��̀(�d�`�c��{�B�Ib�B����{%A�a�ܼ�*���'���*�y.(���K�(�����'������UA�u���64q���'J��l̏*��5�����A�>|�"O�@ץH�4����2g`��$6�S��4}���EFؗ{\x�3NK�ZNC�I�&����y���E
�k�O���Ĉ"f��ԛ��Ʀj�`-��㙃o��}r��� ��Cò�Z�`=wN�x�a$D���T�a�|a��f�����"'D��Bc�I��igc�kZ�:��"D�T�Q�(���-�/KJq��H D�+ Y��H��&�S�<A;�A?D�lt�b�$B3��3D�*ՉW%9D� ƺ�zWG�scV C
+D�,x#F�rUn���.�@�0�kU�,D���7�F�g,�i{ ���]E{q%*D�03Q�N�=8���a�<	b�x �L;D� w Յ~]@��g�<X~���'$<D�� �Mႎ�:.%H��V�R�Pf"OP�s���C���[��]�t����"O� (�k /9�T��C�j�bY��"OT�"A�T(6��MIgY�K��i�"Oh= ��=�� ��o�7��X�'�Ib����@�a*�Q�`��Np��k��$�!�\)d"���(�7o������j�!�d�[2Z���`��X�Z�	��A+r!��!j���v��P���Pǋ�e!��FH�Xs�L<�������Va!�Ϭ �ReJW�ӟ5|��.D�!���Q��p�@�7^S��e$��g�!�V�Y,��j7QR�K�l1~�!�dVPu@M�� ?o�&��bL�M�!��u�ޱ��������y�!��'�hA�IL->���D���y�!�$B�-#�ٺfC4X���oo�!�<M}���`ڗ'�ʩ{��6!�䀖O3�,����.	�6��Խ[N!��~-���O��E�G�� E=!�gi�QB>zv��7
f;!�DҦ܎`"�`އ	 ��7OW!�$��5^���o�V��h3��b8!��Y3 �qB u�q�V �J !�=}� �zt��!�>DY��ܲ!�DJ;L������8]���C��S>y!�d#]*8��������`���!�D�~촄"!Oׇ~�b,��}!�d��
�����D�t��7�Љ!�K�uX�jWe� /�����ˉR�!�d^���)��)��m��xB�;�!��׫W��=k�Ȫ�F@�R��:o�!򄐀t�|!�NT�dnd�ڔHF#;�!�d�)ŠC�FSF�������
�!�dH5n<����"����ʈ?�!��k_
钴�<�扐G�]�G3!��ɾjb�l�!R��ʐ�W�o(!�d[m}����L�D2/
'c!�$9>�PREmB�5}�E��9st!�D�&=���+f�׃J���#-�6q�!�٩vĀ�qT �64��O�8`g!��2B$��gD	����3�2�!�N���a�N�T�F�ǆC��:6J�xk���X��B��ѳ'�C䉩>�*4K���sa�T���н}�tC�	t�h��̖�q3�xQ`�J�\C�	�=!��9�N�3l�
7�9w� C�ɖl�pZ�E͈t �=`'=j�B�	�H����@4Si>Vpˠ-* "Ov\S�d�y0�$�� ګRH<�1"OƬR��84Z4��j�K�l��"O�-��'ǳ9Q4��pd�%A1��5"OL��s���!R*ïD@|C"O!�`K	ک����T��2 "O8�pG��
g���P�!)"O4�W��!JY�=Bdo��Q�t"O�ڶ��#�8��c�I
r�"TZ4"O@Ę���<2 4ɂD˺d��b"O��s��۞O���B��U�Ġ�"OL�JW�H:�M
�#pǔ�	"O6 {���xl�Hc���R�p�"O:� dD�o��%��� �-��4�"O�d3�i��0Pe=�d0�"O6
E��H��1�B�&��W"O� |ՑQM��;� ��\�?j0���"O�D��b\�0i3Q�VAD5��"O栋�5OAn��fM,K�kD"OJ쫒J{� ]��Ѷo1Nd�R"Opڀ�.��dq�gEJd�9�"O��� 	*�[�3'�a���"O$)7�R$�
�Ic,Ir�pkd"O(��Џ�&h�僇�*n���"O���CI��+�p�a�J_�|@�	�S"OX�zѪB1vB-�a���7?~HI�"O�U	�(���R �V�i&�Ua&"O0�k�	�i"ɚb�"o�R�� "O�H���Q
w8�R�&��IB��Ѡ"O|iwi[�aN���`��)2�(�d"O6Ԡ���1$��Cvc��!�{�"O���ګI��#��^3,��$�"O�L� .�(�(SЦ���~�k�"O��1@�B�]@4�c�βM��<j�"OX8����RD. �s��'�5�P"O$y9ਝ
a�����A�t"�"O83��/�D	���3	�4L`�"O�����NRl��p��hY"0�U"On�KWL8ofL�䋏�u�e�"O�:@*�x�����e{�"O��)%�I,F�ވB3��L����"O���N�/O�E�c&�3;ؾ���"O�q�eFK��,M�af�W7��"O�q�Č��q�%f��U�A�g"O��aj�߸����N�uC||��"O�i �X'�̥@�%5��(�6"O�I���]j0��Q����9��ȲC"O�h c@��^u:Sjŝj@�:�"O�`+-@,�2�a4ꛂ>"p�V"O����*���;V�=\|�b"O��
����P1u�2>3h��"O�y�v8���p��q-j���"ODG
�
'w��F苒1/Ry�"O�ej�HD�=לMA�G�XpB9��"O:M� 
�],������"��dP�"O�%J�-6���+�@�
�T�0T"O�aA"��j0ҏT�>�>  �"OL��jˤvЬ�aN�,Sv0;5"O:D����H��s,��y��E�"O,�ć�&��Q��<Y��,A�"OJ�q���0	`ā��LhQ��"O�uP�.��n����L�:Q��1�"O(��"!������
�Z��E@�"Ov���%F7������K�P�6�ڑ"O�����YL���.R�n�*L��"O��c�֘"j�S L��	� �1"O$l�Q�^�/)�I��^��"OhŋA�҈i�u��X�"O8��aL;L�����FM�)�,P�"O<�c�OW2`�f�cE@̀	~�(rf"OQ�e�� >>�J����X*�s�"O��ԆR�G��ԧʹ|�
+0"O���ዂ1馬�'�*�}	�"O(�A3�/j0Ї+r��s"O���tMʭ�0��N9M�H]�"O�"�2'H��8�/S$�:�pR"ON�r5E2Z " 9@���~|*"O�h*Š y_T��ǡR1|Xi�"O�͓c��/8��P0�S�2@�pbT"O��A�fP�;`, �kЭAׄ=R"O� �hq�'ʚk#���T�I#^�h�"O ��LɣKD�:�J,��"O��� ӎ8�v�S� E�(�!"B"Ob9ːL�!+����/�nyhb"OJ��EK�q�puI�.�[�=�s"O�e��Mܖ1:��8cmĝ=�~�R"O
�"ף�L��)S�Ų��z�*ONI�vo֒.H�q$�7Oz,2
�'��t;U�ڦ Fȼ�U�˾q�d�2	�'���0�I�'���!KU�����':���dΑ*qZ�q�[l�T��'�p�����G؀��i�	]��%��'ވ�"�A�qP��)��I�|��'wai�ʓ�y��0��������'�r�A�O7c�¨[V-�}j��2�'kNY`c
�;tF��5`Z�w���h�'�Нy��ۜC��i$Eݭ e��8�'����2��nj����-D��
�'���j�!�DJ&m 		.XQ
�'�z���V�<E����
7>��'����E�ME� �1K�n�0���'� �r1���V��`���l�&E��'zPi�� ���-3��@�a���'2��@�!jV�5�_�8h9�G�<�I
	�*�rsC[�P.=��C}�<	�![
�xI�.\�|H �Bȃw�<Q ,Y�1.�I���#4�2��Vt�<�$�ɫ"��: �	�֤��i�l�<Q�&��h�k�O�h1�XX���q�<уf��]!�b��P��ׄ�j�<Yp-[�}0.���@�tPLEb7�Mg�<EI#��J� T�.���d�i�<2 ��HXp4áh��W���� f�<�$�^�l1P�i� ����iJ}�<Q.Rs~`��a�hM���{�<�q*̎Ph�Ys�B��0�X�j�z�<�R��;el�j��Q�'�0Mآ��u�<�m�;#q:���xLt-p�`�o�<ٲ*� R`e��\<h(���OU�<�HE*C���n�0�X�#�JP�<	ek��żu�&HM)��� QM�w�<	���i��!���I$"l�t�c	Ew�<�2���(��9"�ϊ7'i�-���u�<a��F#X`�F�ƶDA����X�<)��^�I�(�z�MX���J�m	V�<ႭÄNQ�P����e92�Bq�MU�<	据NV�1!� �(�$
p�Az�<Q��	6"�⼻'/W8Z0-U/y�<CC�2-ReiQ��q�J�:�Ȟ�<Ʉ�vT�:��[�G��AR��[B�<�#����In��L@��K�{�<��ё+��-!# 5 V"ma�u�<��dP�tQ��B!��2@}n�@���r�<«��m� �
�ė6��{��	l�<�s虅i���@e�ʴh.5q'	l�<AЊD#l$�9��ícV�� �LPk�<)�n��T�V��;䱱�ÔB�<Y���I����PJ�[7dD�eH|�<F-C���uzG��
�2��功{�<�U�.���Pa�*N0��C
v�<�#�3gk��#c�l�*��.E]�<�s�I�,�"�R MōOfV���Y�<y��E�!4���E���v��XōHN�<��*������9o@�0�UF�<� ���F���pFb)A��
�0=llʓ"O���J-8���џW:����"O�@r�Ͳ[t� ��� d����"O��3�@/;�r���-��S`	ks"Oź� �j��>8:�R"OȌs/�r}�%�� 	P���"O�<�GO
d����A�|;չ"O��*���v@��� ����}��"O����:����	<t�H�9�"OP%c��N�Q$�L���߫.f�mc"O�}��DG�n�^���G�^RNt�"O�`	��N8�a�ǆ?a1���"O���#S�(l>��5�<���'3�}A	] ��p��΢p��0�''1!d	�ږ��J�
QB6��'�R��!�Z@��2�0s����'L�A��Q<cD"�Pd�0�'���,��KD����gЉX��i(�'�LlqҠ2_!�iö���V���K�'�v�eȐ,E �R��K]D,��'|A*Ra��)��)�V
H���	�'�`��ϬZ����d�"A�:�	�'��Yb�f���hD� 䏀UԵ	�'��5xB�E�nL;�!ǇвMb�'aty�c�^���Kx@����'̪̂�Π]� ���dZduj���'�\eq� ��R3�� ��G(nH"-��'C�3s���c�	�cX|��'0B4Q�V�B�0��LY#kI����'ݴD���_`��А�@Z�4*8�	�'2}p��C9l���e�<M^�	�'��zb�!g��<��L�����{�'��B�*���"ҧ5� }H�'Jd,�����<в�f�O14%�B�'B�ذ�n�K��KG�N�/gp[�'UF��@�ܦOB�)���OH!1�'�&	�$ԭ/i�|R�]>ܺت�'�/3�a`1�%=���c+��y��P3j1���&�	����HP�J��y���#D�t��%�
�lB��y��I�lQc��L�Ԟ�G�О�yR�ȘN���H3F	�TQ���y2�C�9�4QC�f\&?��1j&o^��y���0b�0pj��LF����p��y�!_)2X��K��j�D�#�?�yb��Xr���cZ�LعS�ɜ�y��>jX`���5���wN���yb��cA����.����"A���yr�>5x&�3ĭ�#ܹY2���yɓ{Ĳ�@�7s/ع	Ugԣ�yҍ\����tlG6sW�`�T#]��y�`��2(n�p6��>_sV ���ǭ�y��1i����*ٞSb��Ku����y¡ΪBF�y�4Ea8l�6�!�d���b�@���O���0 ��N�!���
�p"0�+��ѐ��J!��J�f��XI�%é	 �{.�N!�đ�~+�]S7)��#�^	�Ƌ��7!��C�vE|�j�M��0�:�)�P
p3!��ߋ?���У�
�e*��r�jL!�dү7qX\�)�%<w� �d��:=!��UO��r�)I�n4��k֥'}!�Ċ���� ����P��M[�hޣ{z!�W 3`jR7�+��34���Y!�� �}���<w�8!�����N��c"O>Q{ə��@a@̎!�^@1"ONģ�#�!T��bE
�d3	I�"O��K�.Z�ն�Z�k�z4�ؑ�"O�iA-�3��Aɏ&R.x �g"OZ��0O���P���Aְ�"O@$�уZ�C��� �Jf5�ɓ�"Or9�6��;�t8���2f2���"OnL�s�چ�����8�u�""O�ف��]5: y�ˈ_��9E"ON��P�]*�!�����9�У "OL�� 
�laR5Cs*I�T��J�"O��2�.��Ļ��V�)Az��"O�q�#`P�/�W�Ӌ0@�)X�"O���C�>z����&�8+rpQW"O��h���Um,�S��_�6��S"O�=k�)�?ED�8sE��3t��"O������+��A��c� Z�Â"O��7ȧK��h�߬V�u� �7D���B�T�Fv���d��8WZ���i5D�L�Ł�-Wi�$�$�]1g1q3�3D��)�'K�[��§�Z;Vv<��n2D��{�o�"�U�@�Wu���@0D��A�DN�9���D� �%�f-D��A�*)�\3BH�'h
��f*D�|��F "l@�١O�-�����2D���#i�t��Z֯�x[�����2D����R6qeʰ���\�N�~��E�6D��G-�5y��Չ���])TT�"#6D�0�!̈�$`�����?E<i�4D��%�P|�J�Q��-p5)7/'D�dp6�T�e
Lx)ʏ1]8����*D�D2�o�57� �P�N�t�����*D���p��B��i0Wm�`>�A�H*D�,*��S�T7n�R��Mk�,��,D�0����3w��-�jF�}���a6D����iY�,��\+oè^o�耄�4D�t��F��6��P8Ҡ̓O:�0I� 2D��iT'W�a�ܘb�IJ�f�bA� J.D���'�� s
���
�%HN12L/D�,�C.2�x%�8yz��++D����̕ 7?��q�4!
"T��a3D����o�*�"�o���<�t�#D��z�-A��'F�8&�p���"D��11���s:���_��J]��E"D�!�� .t�nP�c��C��5D�(�Ҍ�?�6h�$���ƌxg�4D���"T�rn��ſL��ȗ�7D�P0�ݙ$���Ƅ�hvp��0D���#�=&;��	c ��X��%�c.D��c���8�Q�"�_�etN( �-D��0�+�"
_H �bL�9$m`u�Ec*D��Xwn�?*w 㙹q\CGD;D��RT��^쐅薯��Dq(xum=D�(Pe���/8�@!�μv����B:D���e�D1�5�c�u�y��,-D�肧�C�P���� %�)'���a*D��+4ɇ`L�n�*�x]PS�,D���V��t�����A�8�v¶�*D�����ʚF�D���F�^JNj�k;D��B�ތ3E�<�0n/e�Xa��M7D�8��1k{� ����;?�`y��
+D�� �@�# ���UE5�$����6D���E͕pp�s��@��t 5D�� �9(�8�<L9c'��)�����"O<�ȕ���uVԵ(�E\;�8�{�"O�����4;! ��C^+T�:!5"O.|@�1��� #C6}�N�q"O�ԫ�o�Uo���ցH�R��9"O����oG7n1��a�FЏl�d-j�"OX�q��\t|�4�^ R�80K�"O�Qc��3���Q
^�" ��٢"O����iHT�R�r�B[wd���"Ol����8z�T	{�BُN^f�R�"O����(�����NM��Q%"O����ϯ4t�q����5@�"Ol����=Dn|L�NR1z�h�"O^d��GU����qlޗB:�]��"OR<K �Ċ �BT�W�F�#̱g"Or����ŖZ�D�4�6?��9s"O����T9;/pu�%M	-�X��q"Oڑ�r X=n�m�7l�JH"O(�i�G�5=���'wOօ�A"Oܱ�F��^��tP�$����T"O���D�U���h
$E2�`�Z�<Y�EG�8�9���[�~A:�mR�<��N�^��yE��_?�ЗML�<Q&/�+\�u+��I��@��O�<	��X¨P�&�J�}:v��W|�<����Y��m��(�0q2D8�%�v�<���O<!��]�U.�.";&ɋ��Mi�<)�#R�%���AJP-;`�k���J�<AA�����iP1B�>p�4D�H�<��d�&�4r�m@�ڱ�$�JH�<�-G"�z)�b�+g��f I�<1vi�e��ybDƛ��Lp'MF�<i�L���'JχJ�CfB��<�JVϘm���S;&����o_z�<	��+X�6@Zd�I�f�K'H�^�<��⟴��t�j��4� 595,PY�<���-2l x���I)�<E $ |�<ab��|8Ҕ�e��$E��@�RdV}�<	�M���̺T�H�c�P��`��x�<)���p��K�:����+�t�<� Y-{�DS�b\��>0��v�<�`�4e�`�c%+�C��˶�PK�<�Ǫ�<V�pY�G�w��A�TN�<�Q^`}$��⊄�0
�Y�j�I�<I��� �� �7	�	`U��-]�<�$FP�&Y�ԺR�H�d�V,a�`�X�<F��S�Z�"a�j���(P��U�<�p�W>���A��Q%{#0�(cb�R�<���d3ب� ʵi�(��aDT�<A�B�<N� z�%�U>Ҝ��@�S�<	F@�9bH�3A�qb�f�<a�_!���x�ƚ<�L4p���H�<��K�*��y���}ͦ(��eH�<	5��I�\���φI�����P@�<��E��9`���]�؀X�<Yש%�l��#֢��r�D�L�<Y�#Q�U����jG65�	��EZE�<��`�) Bhh��F��s��A0C�^C�<�E��b�qA���SmL
��d�<Q"�ı
bl̺�ɚ2ih|���U_�<)�B�T.L��d�8���f�<Qp�Px�
Ma�
9�䠸S��d�<�/�4 ���]|�\�&�G�<ՍL�y��#�.V�Y�.�`�h�[�<� �u��h�I��e[�J��l����"O��9�I$Gb��Q	α�|:"ORU�7d�^Z��A�
��Q����"O:�����A�~�YSCB(TL2e��"O@���L�%G�Q�4 ˰M.���"O��3����u���oT,�5"O8S�ȁ6!b��5�T~�P"Op$XfAO�'�R}�d��g���P"O��I��%3B޹�����q���C�"O"��fŻZp�T陱0+ Sp"OF�Hd�I�Hy+�ʒ10*�y�F"O���C8P����1�ۆe���2"O�5� �>��8F��Wg���"OT��a�]�W�E��(��C��A�"O:�ǅ�	-ll�PοfH,��E"OrMZ倉4\��sR`J({W$@�P"OTEC��K*{  �O��+8�9��"O�i�$�����r/�5%�H�"O���S
2�ջh����;S"Oh ��N�2g�JY�q��& ��a"O<T��(Y���`��z��<�"O\��ɒ����wH���"O��I6%�"i�t2�^%�ܝ��"O�E�ri�8@��t��W"�Xɳ$"OJ�sQK-t(Y�@�	�G��i5"O�y���|F@�32���o��k"OX�Yyp�y�v^7{����Vh�<!�� �r4�iƱ �.����c�<��z�Z�`dm�y��`WH�<	T�R?A�v!��L��d��y�<��`��j����[���&\r�<G��9G;�hS��k�&=H@�W�<��G�z�8��D��(�ҁ���H�<i�ŀ�/����b���;aX���C�B�<���W*"|c�-�=W|�]�'��g�<�HK:b%� (��I��y���|�<I2�-X�ๅ�ךd�#�ɏT�<)��N�S�BaZ�OŠo��ҧ�N�<�r���	�� [��XI�Å�DI�<��"x�D�`cIK}_qkG�B�<y֪Y�( �b�N�<��eõ��|�<�W��-A��y#`�'Jʁ�sH�x�<���O�Xࠂ�/`�|x�ār�<Y�.�(�lԈ��30�����k�<�!��_��`Q�[�B����g�<���K�r���oެfR@��p�a�<��@��3%JǧR^��U"WE�<��Oѐ_��:dH�%'�|��\�<��1�p���'�h�C�,@Y�<��N n.�`Wl?/�E{�"~�<���L=�4�Ӈ�N�t�x�r��z�<���̃?�l�j�7|�aR���r�<�T�N>+2,y �͍�_(�!� �n�<�#� ad�tz0e��8NP�f�a�<�#\.u�]�Ƌ�v^���FX�<�D���#Ϫ��!4=$}����V�<��@�bkl F�ʍE��-aƃ�H�<I�^)yAfDA���lX�؀j�C�<1"��i����,ūh� ���D�<	g@M���9��-���P�s�}�<�*O6{z��{��S�7Q�x9l�]�<�Gˎn�ũ��%_Ɗ����N�<!��%�=�&��4 �7$VH�<ᑈD��R�+���HJ�X�AC�<� �h��A�5���UM����m��"O����b �!:�������(""O�� /�p7��@�� Q��!"O��[�/�)b�P��F�9d��ȧ"O:���-^,8f:�8���&Th%�"On�Z�\�1p���%��r]�<$"O��q��{۲��Reʨ)S�Y �"Or�{�GQ.1���4%�9�}`!"O
H�f�=�ڀ�pƍ �m�E"O�ܰ3F�7!��9#E�<�����"O"�J��Evv�*棍�#gҵ��"O:�pM�1�X�cE��%��"OZl��/ ����倳M��*�"O��7n��C���I"��k�"O����W�n���v?
�h�"O����OF�n�$��-���e"O� ����R�zm��Gٴ:ۀ���"O!��I�]���s�9�&a�"O�Ա�I۞0�܌����%D?8Tk�"O�H��б&��U0�`�M2�-�"O�p`r�¢ �X�!���r:LBg"O���4JJ�kc�!��GZ�}X�T:�"Odus�Lʁ[�F�F��KKN�C"O����9a5+!o("��F"O<���+i�+˕3T"�r�"O�}Bϝ$I�Y'JA�6�؈Q"O��˖��5�@p"d��y:L���"O��E�Ѕ,����'�-�``1"O�L����@�ά�F��I�9v"O�%R�� 6b 0Ħ�38b��7"O���teF�2QƸ�%�yu:4��"O,H� 
�	D�(
�䎄fFj䉥"Oy�c�L�6LK��c_,��b"O�FH�"�:���3]�����"O|A8�쎩+�����(F� ̌Q""O��h�'J�F�$�1�$
:y�8� "O�p���.R`i�,,:_���t"O�H!ׇ� ^���vLؾ.Y�� 4"O��˳�B�T�<B��28&�a2"O9
W����E.1pu{U"O��C� �H4` 	wfTFx8�"O���%�N�h�fA�t�
 [�݉"O&����9{��y#$B)&q ��1"O؉y�M(`��9���X=���:�"O�����;3���,Y����"O�i�r`L�"H1��Y2!����"O8��P@ Do\)h��$f@�P"O� ɒ�
>@��$ �!ɌN�bp"O��$a��j�.�9 o	����1�yR��i#��D"	9o��H��%�yB�B	Z{vR�/�6`m��y�64.�0S$χ�<��<��'��y��˵r��HÜ�a�"t������y��U��Ep��W c	��;����yR-�.`�B��W�"hY����y�(M-1��E�sĈ�Bb�t�j�y"�-qV4{!�-8���Iq�	��y"&�P��ْE��,4�@�`��y���P��-k��F�Lj��y�3nY�Ѩ�E��vq�ӯ@��y��AS�rlk��'0��K$��	�y�,]�-U�@�D)P#)(a���&�y�A]�v;4�s.I%#2<ɂ+��y"�A]�l�1 'N5j����y
� Nd"S�����db�߂
�l��"O^ib5��;�ts�
�-;�L!�`"O�Th�F�+u,4U�%@�	!�"OlΛ )|:����0кP#"O =*��J�BN`d
5ėQ��Q��"O�Y�.??^T(jQ#�-n<���U"O%#ƭ�g�c��΢O��؀"O�yZe�)ў��n��L�B���"O4Q��K�'���(�E�����"Ol�	�
C�&H
�B��+W֞x��"O�<i�Ɏ�q���P�(Ɍ�r"O�u�-D�w�j��@��!O�ɨ"O�@9R���	�'zf�3�"OH09�jI=XCt��K̿=��D"O����+=W�̛PJdڢ �A"O��se�W
0Բm����ʝ)2"O�%9f-ǱqK���s�Kp]b��`"O�ā��'�J��q�]�QC`�HW"Or����..jp��%�,8>�K�'�EHg�0w~�ˢΙ�����'�╊ �C�Ca*ț�"O��Si�.y(�-�&�!g&LxВ"Od�p�O&j8��D[4n(��"Oz)K��Ci���k��D�R�4�v"OD`"���'z=��e��j X�"Oj�`���;BԸ�b��"H�rq�R"O\`1�+U�U݄����	p�켸�"O@�X�嘡7U���V��W���!"Oh5����>��@��ɶU�$�8"O��1��B�G�0�!��ߵ�H��F"O�4:V#Y v(i(�)��<���1D"OJ��W ϩc��BG�4��}�"O|@f��R��,��[-|���"O��Y�Ή)~�
y�(G�P�Y$"OV��E͙3VܹU�ȜC�^�K�"OZa��h��sÂ��G�����@0"O�b�)Or� )&�V�$�P�R"O�8ৌ�,#�����/]����"O��[%.�/�v�{T�7_(i"O��7�C~�J"�<��S"O ��� �I>^�Qv#vKA��"O4�����(S��E�
w0v���"O4,A�W�6J�X��A�.
���"OP�4@�%�l���ۧ�>�Sf"O i�6�ɻ'i����ڳO<�Z�"O��bPG�^A9A�8E��\�%"O�	��M�����#�Q��a�"OT��­Z6��){���m-��"O��� w��03��q$�@�"OpК!�В�$Z�ew8���E���y��`ش́���?t=:YB2LE-�y��i ���c���q�W>�y�'�ʪ0@h �f!�8"�VX�5I5D�tI4��o�P�jǯ͙/��1��4D�(�Ș.P ���̞�C?>�h��2D�<J��68�������#�"�$D�$K�g��� ��A��6r����"D�P`ގ�2�1m�"A��*��6D�{D�<��B�J1r��y��i"D�,S�	нi�d2�-S�r�ҁ��;D�ԋ�F�� �9I�-�(�#9D��A���R��C�Ϋj0���ӊ:D�L��ǵ�!���N�uF8�ѧ�<D� :�oO2[ �Q*T��k48�Pa9D�� �0�`�^��+V
����"O�t0V�ų�8y�ө���-A"O�{sI��W�̼����
/EF];v"O����HW^�,�I#�����P"O���'!A~ެ�$��&�����"OL����ɨ��f٬��"O���o�N��<��/�.$Q$"O�5�%�[&F��� _�j��x�"O��f�0K�> :�	]9����T"O�,�k)C��iq��r���Ȇ"O^�"&f�2]z��8 ˎ23�� �"O�����G:z���ק��/�4��"OJɉs�ۘ)p�� ���!�P�*�"OFE�� ٥B�B��'7�$T1�"OtA����R�P�a�2�H�2S"Ob�z4bQ%S��؛�ޟm�li��"O8��j *C >����@�(-f%��"O0%�櫓�\�]�#�X��$I"O���͊b���EL 1��Xi�"O���L$�K���H��z"Ot3�Z&5�c��@����"O�� ),�l�gG�B���a�"O��7 ]�y��}CE�N9G��ܳ'"OL���gS�x	�`�b��4s�I�"O|� �͜.�R��R�F�V����"O�rJ�w�����S�^O�\��"O�1�(ɟ*8Lb2G�:f<viӲ"OP�``�^�k�P���FG?7���"OfQ��ƚ9�:��û9*�yQ"O�e���!I�<x�f�7fhl�w"O(���kO
B�1�æ9;a���6"O�A���%�PL�g摆FF��c"O�}��Dr�n$	�$�=�*C"O��1�� �D��3�Y4�<�&"OD5�MX��b�-�A��"O�@f�02V� �H(V���"OL]葧Ws�@@
���I�"O�����W;@�p��^\x��4"O�Ӥ(��s��!a�ԲB���`"O@d���F�t�a��ꃀA��QV"O��3�)#>�B���i7��l��"Ob��q�\
FJ��g�05�nYi�"Oj��`a�+T�(� ��D� m�s"OH���C3���3�Q*���W"Od�x�@٨s��a B:aP @�#"O�Y�RhՏ\4by��oΐy�I��"O�HP�ǫ��-(�n� D�Lk�"O��̑�P���$g���"O����.
�CU��ZB��,/`naV"OČ vg '8���p퉉TP�r"OP���N�F��A�)�}a�"O����?~�� {A�"~���� "O�+�n�5(�Q��C �*�(B"O¤b��߁#4�q֯3r��s"O�m�
�R�@�� NUTр�C�"OX����R��HAcF�\*ʢQ��"OH:�a(3��܉�޵I"X��"O��p��g���[�lL.G��t�"O�����9LMs�n��X�,�"O�	 �fB���X�nd�6"O��5L�ۘA��-P70bj��c"Oe�P�[pQ����X�zM�4Zp"O`����<k��A�&B�P���ۓ"OtL�weR((�p��B&L1y��)(�"O� ���v��tWZ�X�$�$r�n���"O��@��,s~��`��̮�J�"O�,[&� �]�RO	6�v��a"O��ɴ�<Lޠ�G�W�N�zś�"O�k��P�x�ƕ�g��?���R0"O�D��%����%(����P"O�e�g �/[R��b�ǆ!�"`1"Oe�sjPHR�2SX,P�"O�t�7���8�����n�: ���"OR���H��8-��Н"�"O�s�	��`B,�c,��i��� �"O��Q���+xY�|q�k��:Ɋ"Oн�U��+YB0��֧K<.�|H "O�q2��23^�3���(H�"O:����7_��H�nœgzX�2""O^=ѱ~��%�d�"0aHx`�"O���� 
"j��rk�38S��k�"O��;#(��d��Y�� %PMF�e"O�9�jݓR�0qIG
f6����"ON��6씥7�Y�v'^-7"O������I�4fߑ�H��"O i���#����&FIs�"Os����w,H!��"0l�aB"Oh��A�!Dc<�걃�+l r��Q"O�@�NX2$�4hZS�ãu�P��'"Oh5�G�J4�v5��f���Q�"O �7l��@���$�BhkQ"OPA ��!��Y��hB�wd�� $"OH�#�rϪtY���zr@ۖ"O:\�7�HyV����Z�/gt�x�*O���`�]�hph�0�:�;�'8H[�b���{g$
.%+|�;�'e�e��t���і	U�.��X�'nDM�Rd� r ^�S�ƙ*�x�p�'26�"'�V��#Ц�+vg��K�'yR��f��{
�3䎚�s>��';nX����BC�p �E
g����'c"Њ����ue�(�� _�`1�'V�Ra�2D�q�"�P�[S�(�'���{�j�-4Z���^�U�.���'�����P�^��>e:M�'�2Q���L�.�^�3��Ȗ^��
�'�#�ǚ�Ԯ��у5Pl��	�'�N�I� N##��A	�-G��a	�'qp5�"�K#��E{G��J��{�'x��cg�����K�b�����'��-r�/
+��趆N�-���'P���G�e����um���D���'��,�R �$5���� �����Z�<��b:�Nh�eC��U��|�<���ƂA�d%Y����3����C�|�<��$IG��������`̀2��z�<�3�ҏm��,; g�`��!dc�R�<�E`�XD��k̕FE��Dy�<q���!"�UW� 6pͨe�K�<i��F4& ��0+�*V���p0�A`�<A�dA�sX�!�j�%ǚ,P'�X�<���*b��Q㧫E/�pRC`�^�<���DrQg�b��b%�]�<a�-�/�h���]qj$��MB�<��й��*�K=6��K�V�<���ʃl�
��/�]�Ha[�GJR�<���T3DZBa1���"����a�C�<Y���.^���2�'I+#��k$��A�<� N p�+��6P��h�E� t�"O���SN�^wh�%�e��y�"ON�:��ڨKvh�qGV4D� X��"O��sL�(<��h#D-�g�Z+w"O��9�`
�_�L���2h��ɓ"OH<xQ/�jnP���jH���2�"O�8�����vHl9��?��ź$"OZ9{��ٛV�6a�@�;(��M��"O��8 ��j`q�J�zM�%"O��@aX7� A����L��"O��d�F��D���F���F"O�r#LC����bA+Ռf2�)��"O0Y���${^�M�A%wȂ���"O��3f��h~xq�0�9JZ���6"O��s�Ń\T
�ӆ�;4��c"O�iZ��~%J��lM,38�`)�"O�,Hя��yn���7�.,�՛�"OD����|0h@�?��7"O���eU2nTks(�T��jf"O�,ɥ��<F눬(X�S���#V"O�$���ܠc�A�a��<�RM�A"OXHÔn�,h�DY�q�D#�����"ORl`&�S*gX E`b*�4	�����"O��C�?O�52�T)zt��"O�=��f�x� Q��خKqFaa�"O��#�lјj䜻W��[�1�"O��zs��JVp�`)��fN�IU"O�<K���^�5�iA6�z�"Op4�@�,O>�٢G	m��y5"O�� �3z̓� ��L�V���"O
 z�`��1���+�6d�3"O��(���7&hȂ� "��H""Ot�"��Ц-�40��4���Y�"O����l�*l�ؓĚkaJA�R"O��`v�G�@����<B��2�"O�����K3x����V�K]�Ԫ�"O@���%��O��9� ��DS�D9�"O ���dۺG��|���S����%"O�a�Re��	n���SD�N����c"O.�3�G^U���0��&Q���k�"Ov��KG�lJ,�@a�w�blCr"O�Ѹ����v��o�W����"O�:�I�#�L��N�*g����P"OűR�ۨ\�t�03������"O��;�&-Q�<�
��)n�
�E"O���D
A2~����[,I�h���"O(��V?3���ȡ*כ Ahuc�"O��As@��%+�Z�C�,=+� c "OP%���R�l����aL�d6e��"O��jUC�.��YB��M=Q
LA�0"Oj�B��Ip�lP�Q�B�\~u��"O�uI�R*8q�l��(F�i��t��"O���СW�c�$(��ڨ��%[�"O���P�A�o��Ȁ4
$
n� X�"O�퐠f��U��B���)�0�a�"O0�X��I�v�Na�OC L��X$"O�i��f��l'�a����gݤ�{�"O(��AT6t� �g�{�60��"O��1�m�S�ʕ@��ןQ����"Ol-�����R��fL�C�X��"O�H����v���%��d��"Oڥ�p��9t�渻�iޅ�\�P"Or}`pJ�qA��*I�~Z�(Z�"O��H���j��� /I?lo�,Q�"O� �5@���%WMT�@7�-��"O&#��j4�{�,�>\��"O�9 �Bқg�b�����T��)�"O��ktA�;(ɮHk�K5eo���1"O�tb���J\�5�1��_~����"O:��a��H�7�� 5����'l������a�`�a�`�IeV���'�깒�
�gE�ᨆ��E����'L��23NJ0iYL��e�V=)O`��'Ʈ�x�}
f!SeG2n�JH �'�*�8�\(x����Ɛ�a)td	�'�'�v������{��!�'�`��� �sAʌ�-�`���'���%׳�&)Y���6s�`|�'������|h.�%$�X�|�H�'��SEJ�%6q�U�X8J�\t��'R��q��"$�n� ΐ�kq�a�'�p�p��x�� ht�B�.6���	�'���S&��5h���/~��T�	�'o� ���pG�90OU�p�$�H
�'����j��8�I��N��1��'ܔ*2(�l�؈6����d�	�'�]:�&�"f�iA%�)}-���'���*	����Ⱦs���
�'24-�ƍ�	��� fr�����'���s+%K`���j/Y�P��' �F!Tv�v瓂x���'! �Xt��+[��qO�4id^��
�'L��۔� �\������[|�dC�'����!N�5�Lܪ��Ii� �X�'�&�dn�� i�B�*Oo�c�'��i��˹z����*^�F;�,�
�'"��PD��[����'�,kxb�'�H!�7CÉi�D��ʄq�+�'�(x�`�U8Ȳ�[E��o �ٲ�'��-�6eO4�|h��_�dݬ+�'�а�A�EH����b���	�'��ԙ����&-����
	�'Ű$�k]+o~HA���m�� �'�ƑS#��t�&$a�鐶G����'�u�@���?���2�C�	�0��'ìᑓ ݤ4�� b�χp�d3�'�-@$
YSc@Y�AmS4a��'\.A��F�T��p�LƺX(@!��'�ts�(½p
 ���5L┙��'�����ˀ1^��B�L�>�ι�
�'_H���`�P�Js�ĩ
��	�'P���-;+|I`��^#k���
�'��Ȑ�=/0�A鎷e�~љ�' ��T�[�Fa8$m�XUԘ�'�NԩT`�1JX�DH,M	4	��'B�{�)P�I9��a�H4�J�R
�'��b� �!-�>��"N�0%���
�'"~hڥ
��*�P|x�+H�!����	�'a�Eq�̘�U��4����-���',T`���a�@����y�U��'y�Y�WI#��������[�'��@���]s�j�CܟF���
�'�����&ձ,��yS���w7Ԭ�	�'4�C ��;b0h�d��[jN�+	�'�z�U��0ҳ#W4T���I�%i�\�AE$0�����Jm�ȓ%f@�D��h�ĩ+�Ϗ�gl����7�@�	���}��s��=a��؇�S�? �)U+tMjh)�l[� ܂y:q"O6pb1��%̘�pM�T!x�"O&��g�1�p!��J�6��"O<���r�PX�0ʔ�S튤��"O�!�b�`�� ���z�ji�"O��1"6_8
���LÏ>ٖ�J#"O.������p�bA�E�4kT"O�l��I� (���{0��e�Hqv"O�р�`S�OO^``3��;f� �P�"O��(TaY:#l!�cXw�4��"O���%�A��u ڙ=��(%"O�i�ЫG�-�P;j�
I�� 6"OR8�m@.,���Y�I�V�Np�"O��D#,< ��@�E����i0"O��B��>7T���=6��z5"O���t�٠E_�t�UO&@p���"OT�[5`���(rf̩B$�"OjŘ7���M�8�G�ܵ�r"O��#�[��[�bP�|��#�"O�X�q�ϊ�� O�W�jh1�"Oވ��ʞc���BD�N���F"O ��"�q�p�D̓8.��L�'"Oȁ��̝;D�xj����v�	@"O�A��J��XPL9���V�w��X��"O� � �:��MC�K�I��I5"O$��Nԍ`N@;&nɽB� �a�"O��� ��p#��$��x�$���"O�,�ϓ	>��p�#Y&�~���"OP��A�^~�1�ݕr�xx��"OV�X6��"{ږU)��U��\�i�"O�)�e�2�Zq�� �)N��F"Op�?�j��ݮd�ZJ"O��o�)�
D瀶K� 
"O���gk)#x�����O�0��"O�Z���}���ٰ�v�&�)�"O<q��)�cw���shT-3{���"O��K�,�wn�P�C��8���"O��i��9]�yT&Q'���"O�H
c��,\�V��HCE"OXq��:@�,MA�L��@�x�"O�!@Uǜ�"p� jȚ�ti�t"Oj�M�y��삇FT)��LaQ"O�0B3\�<�(�0�����Acb"O��1#��w�~$Aa��$pNT�2"O2y���<]�#%��D��Pu"O>LcVN�7OP���D�.+�l��"Ov�c��V}�鑂ջY"v$�7"O�E�e,P����� L�b8��"O�ق���\���F���7�̔�E"O8TJR�ܻ0���L p�f(��"O���L�.:�$���	ߐ���"O�21�	N�>�n��pl�%�"OP�ס0!�@�M��Y�"O=����{�p���)K�<�!"OtU�' W����ʁ
��db�ԣp"O�d���4=a���&jZ�RQڑ�s"O�X�SÑ�9R�b��Qhm��"O&��D疸B����$OئA�}��"O������I��=� !\<1���1"O��"Po��zRPd*�� ���x"O�jA�O>��٨/�pX��*O�Qz�ܓ��t0�A�$.��-@�'�
�A���^�6�˦��-j
)B�'� !�o�)LD� �)X�pX��� ��a��%�d����T"O�X��k "�}�3"`�hk�"OPS���B
���F(ƢE:�q�!"Ov��.��+�عZ��8)L,z�"O�Xe(�8$a���I���B"O��c�G,L3�ôC��D�^�+S"O�-igERT�|��a	�o�r��"O��W�4n^r�A�y0ܠ�"OD��Rj�CS2}�с��SZ��9�"O�̙���f�b�CF@ոK�C&"O
��aI�'!��A��1?.L,��"O ���\�1�tCE,�9�v"O�X��`<5J�*O%茥w"ON���o�kJ�e��R`�s�"OD� Ν�;]��k��&o�(��"O8j&��'RzU"����g���A"O�m#�M!J�M��O��B��"OT�	n<]1&�F[�
1Z�"O���h
�l���˫Um
�AD"O��U	�r��<�,C�:j5�6"O$E�Ƈ�b�K��*�P )�"O��#d��TL|�-�^�b�!2"O�H`���ku~���f#3����"O.�D�Z	v+h%r�e�e٤0��"O�Q��Ą;K��c�% 0�B�"O|�!$M3 ��܋�E��\�A`"O��Q��G�@�� d!K��Ų�"O���d��mT���H�Vn���"O��K�)M��]�G?k��tr"O���@͆/(	�CA�=�hD;!"O~�"��&*pͫ%�F�[��l�q"O ���ЕLk���f�ך=� �"Of�	Ȇ�Lܬp�ӄ��w���"O�����VETk�a	!��e2 "O�S��B�UR�a��T#�`��"O�M��KC���Q�Յs�5�"Op k!`ԥP�0��-��Y�����"O�����6vf��KQ�/�LV\}�<����	�d������1�J\� ��C�ɽo�\�@�_�x}8S��#w��C�ɑk�jݹ�N�&muh�Z�l��q0�C䉙m�� ��;|8	�D�E0&�B�?,]� cFԢ]�jU����=m�B�:6B�;��,eZ��jՃߍgr�B䉥HP���^9��Z�$�)��B䉸Rg��C úH����\�|�C�I�]���Ka�� �b��; C�	�_�p���b��!��2��6~|�C��>,N(-;�@�?`���+�jәN��C䉧B
�JGoL2L��tpg�vfB�I-�&�3�bN2g�� jUś�B��	2<<�`��
h�(�3lٜ3�C�ɮY�FA���ʒbӴ` "��d��C�I/qz4�0�B.s�P���"r�C�	ZI�0��/��y����C�	��`-9T�� %/��ɵɊ�3��C�	�+�,E�>Z�r����ʃP�2B�2fk`@��o�L���a�I�R��B�I�8Lt���H�,���b/�  $B�I4Q�R�I��o��&ʙ�iB�	�!/�q�bQz��6F?C;�C䉛?y
����R7:�V<��M�Z��C�I�i4+�o�(qDZ��T-�PC�	�|&q��i�a�4�y'(T�cu^C�)� H�1�g�D�6�y��=X����"O�آ���_�����O�O���"O�蓴��4̾s��F*��m�"O���0���-�U��&���h&"O�}j�,E'�V	��`Y%��9K�"O�QY�-�;Nީ+��b�P}�"O�aQ֫H����3(T��A�u"O�&Z)�Zu�S`�?YX" *"O.yJ���B �Xj0�!:�5�"O4���mZ�%��cD�<6|]��"O�]�F���_wLi"��
�"O*�@c�R"<4x�fn����1"O��k�Ο�_{�$�V)̭,�~y�"O� �� ?>�q3
�茌Kc"OP�&��qa�X��W��eh"Ot���	�=HU
A�# X�3�R�Js"O쭐��^]#��G�n��"O�)�&e��d�� tA�aϒ�H"OW� 2���0BLIt.��A�mi�<Y��ڀi�̣��&<7�lIa�Yp�<�B �0`j�JN� U�qH@r�<1�Xk� ]�cD՞ �Z�k�<)[聸6,Y��<FF���8�ȓb�l� 4OJ-TPB8�u��4:=���ȓ �4�圮'`��b�&/RY��9�V��f!�)Fu�tk��F q������i�2��b\fM��_�/�T�ȓB��]8��X	2Q~%�d��#Zk6�ȓ��=���_�-�㎡p��ȓ?��x�FO2;���)B�:�E�ȓ@7���3l}�j Y��¸^����ȓy��=*�C	�H#f��WF��v��ȓC�H�I�o�{]ش�,P-������H��Bl4�ٲ�ȧm�LA�ȓ��]zGC�_����/{���LA����In�ŀ��ܺz��X��R6��v@9~�B8c5�80��	�����1f,]�&TL�׆�>����ȓ)C�Q�� ��pP�����\��ŇȓtAJx0c�CI��3�G[s%��ȓ9����L�'&�\s�m1 �TЅȓ�Nqpa�L>�^azc�ɯF�vm�ȓ?b��B�X�Wn@�ã��Iʾ؇�&H����[�z��H+vM,quJ	�ȓQf�M��"�6�"]��%J�hфȓ3�J��g@��t��w�j��ȓnU�� �Q�]%��[!�)�ze�ȓV.��I�����iC�",��ȓ����g�۪$�İ�C�~���ȓ/*���(97����M4h�p��B���0F��rA���3X�`��q�A��k�u����bF�������<�`/s�A����0}쐆ȓR�����'��+V,0�U�B̈́�Wm.�q�,
�v�s#��SQ�A��I���@T��Q��aC�-,Vq�ȓoq�ɊZ0>w��lG�'�J�;p"�v\�I��;Qh���
�'8B ��=/��i F:P��tQ�'�tSsFWG&qykDW�<
�'��4 �H�g��T�(	�'�%3��1�@ �$�0~�H[�'d�l����(51+� |���a�'|\�%:4���AIFZ�Dc��� ��R0���m�v.��I�����"O�tB���y�v���?���ۤ"O��9 ��<IFdۆ��?{r.��"O���AĹ+%�0yE"̍S� ""O�]Ε!9#2(�ۇYA�ȱ�"O�Eq*�x!�u�ֆ)n!��[a"O\��N��7��U��B����@"O<sw��#��ћ�e��iY@"Oz��
��K�I�@e�&Q�$�@�"O����+ɼl�V�y�c\�D���"O(��B��Hav	X��zh"O����]�K$�8�j �.i��"O�ap��Ш�Pk'�D�M�8i��"OBT"���'.�*m�w������"O��`�^�!܈�������"O`��ϬV��A�4n�R��<��"O8�ѡBO#tZ,I��d�]�"O�� W�[�k��u��\@=�h34"O����
�y�p���"4�X�A"O�$@���m׶�Ɂ�،d'ʐp�"O�œQ�F�,`@��	�|눝
�"O6ABH@B*�h	&m���r"O4x���:e"�\
�%W�Q֢��p"OV��s�.B�B
�E���y"O�ԉc��9u�(�CR8ydx�j�"O��zG� y\���"�8,�L@8�"OI���<S�4}�����\�i""O �@��=w3�ݓ�O�d����"O�kF���C0����;t�*)�2"O���"��^���#�m���	��"OL(�Q&�|մ�8�b� }E��s"OFݳ���00�⑰p\��+�"O�-�⎘;;
e�tAY�g�\,�w"O����ҙ5Y�(s@�{���҇"O��"*B�FYY��`ݬ�CQ"O����E6 P�J0�P�Eڼ "OV0�vė=P&As��֨m"�p�"O�%����}Ќ����-cA��1W"OF *r���8)�ᚈm�`�$"O�8B����ՋG+�X4p��"Oq���ȟM+ƨ`�IM�$�Q&"O܅sb�ZF��S���vӶ=�"ODh	P�,Z1�+��ŝt��YC�;O������2cF�1�_��ZTq��IT���"�`R�L�#��`�VC�ɷ��H�ᫎ�~\�7W�=%(C��'�<ت��ʉ"�d@�ƀW�I>:C�I3aN�al��5��R��8DAJC�I<5^D�a�\���Iw��:ьC䉇`�lʴ�	�,Q��^l�B��=p��<2��G�8[��C��:Z2����g�UW,�m:t�C�I�&��9q�7_�0��"ؔ8uJC�IM1��P
�.~��X��?d.VC�ɞ4�$�0Ӄ	�>I�*U�zC�I�x����#�}\y)W�P�=�LC�ɵq���!��X�1l����:jC�  3�X��b_��+©tN�B�I?Qa�X����o�*X�w�� �`C��T������Q�^�����;�B��7(���T��U�B�K2�ͼ��B䉩^YRT���j �(r�ϭ�B�I�x�$9�M� �μ�UJ
)�B�I�9�Z�#�a��0� ;�g��&fB�	$@$`�򆉆N�$A�V'�/ņC�)� ����T�w��3�C��+[v���"O4�B��/L�L�S��K�TF8Uqc�'�N�C��#���Am
̉3� }^苁 
�w�B�	>��H`�D�4�}��3;�'k��r��f?r����	�ԎF�m���	�%�T,!�����4i��^�:�L$^�|9+ �ߎYZ�ɲa[r�B6��|�bTX	(4��ꕮC �X"�C���x�T[���������*^�0x}�B@�l��8���>�O�k���+fL4��7W� �v�����ApAl5kt�D�2�?	���G4*fޱ��-'��uf�=D��z�����ڄ���5%p4A6M�<a���R����aDضb�X�G�dl~��H�A"�hk�L@:[f.���'��Â��,�����b�Pl�p��
2*`A�RO�M+�pHu�����,��D�6C�k�$�"�~���d��"�$hq�%�4�)�3$��)��D9��44zrIK��X�:H`����/�OV��0n��u[%Cɀ�b����>�\3�`��m��A#���n���O(��*EgӘoe����È,X�x�I
�'�r��w���M��d�����D�LW;�Dt�t̎7�dd�@k
�B�z�G��we�t&�&���ˊ�3=H����U�m�M��鱵��=r����K�JT�d(��_B,�k���(q��IĤO�Q���Պ v�dn�"D�Z����Q��,Z$NŮX'�0���ԃ3|杈�.ӂ@~��)	��5" `�
n� 18��*�O �PqJ
�$e��J��I�x�җ�$_��l"qB՗D�L�eH�w�H���ߟ&�C2c�9Q���ăL#YlYb"O\�L�{Z�0�O1%s@��f�AB�"x�W�� K��,+§oL	��t�`�y��I�M��8b.Q�f��HF�!D��P�hȚ���z5��m&�]��B] ���QI/QL�D��B&'��X��H�Q��p&.�V��N�4P�F�	��=\Ox�;R�>Tz���"X;w*���,����	��nH9�X��@S�i��rYO��|�G���HX��
�йG��߸'�Ԑ�b�,9�� h�����l�6�L9a!���3W� ��v�Y�a�����A�=�FC���� 壉��1���'a�h1hࠌ�W1���_0yW�AZ�V ���ݓ�wG�b�����K�B^dִ�I`d1D���dM��
��P���c۴	�Ҩ�:K��q�`��r�ua-Z2+�<��$�\&�Q�dq�ORQ|���D�O+/�%��'"\O A�c�	x����P�H�M>d�W������BE0&��y��}\t	q	La8� ���5x5I�AF�4-T��� 3�	/@y0i'��H��5��Y�u�����|��4hf@6O�8T p��%�y�攓ru��"L��F�V=@�dT�:i@aǇ�)�$UZ�UKN)���(gq�.�)GKn�kr�J�F����[�!򄞠NTXJ��I���P��I`�V^ O\@r�O���L��� & Q�DS�'Z�\�*B&Y|� ��
�;09;
ߓR��S�� \�L���&Xv��H� �p=@��#�ם]'�~��8A�Ph��l��:9��-���O�)��E�r�:�Ƞ�S(MB �C���<���{f@l�B䉞.p�Is���n�-rS�O>zՄ���4Vxx��x���'<��1L�+�f�'�����	�'�D��)e�y�6-_�-t�y[	�'&ʜ�m�6��IV�ɏ Gj�I�'���j�&]ɴ�xfE�3��}S�'�N�k D�)t�� U�[�%p����'����0�:��	���@��B,`�'��i�q�ی\�n1���Q�E�	�'Ќ ��\�ZɘK?Kԕ��[�\�p�*V�KWri����?4�x��'�Zx�K*=��[�(�9_1<܇ȓ|��{��X�DɆ$��"]�i~F��ȓF
���r+�;���bO�4���;����	��X)F�����s����ȓص�ף�{ʆ8����3A�҉��7L��� Uh�0�E���=��ȓ � bD��D�����[Zz�ȓ�}oȲ6��aҁ�X�	N�Ѕ�,�~�c����=��uR�G�P|x��S�? ��)5�7+�L{5�\�z��9�"ONP����U;Z`��ۧPbց�"O�y�E/�=[������F}�U��9���pC@7��ik�i�pvH)��w1z݊�JF�~��{�H�9-(p�����M�p�n��`�E<M"��V�<�AO.a�\��a^B,T��`�n�<YN_	��42֡8A�(���A�<��B��&q�a��nFxe~�l�A�<�2RlW�b#US&��6*
t�<����:JN�X ��:^�vy�"O>H���$QgL���-�;N�"��'"O�=��-E�6�����d)�"O�mj%��Mx4
QKR�M�(�1"OZ�jf�!/2jh�
ըx���"Oz�)g�ͫMC��bl� ^� ��"OP2!RO:m�%��A(���r"O����B�7��XQ�2�p�bN{�<�����P/N��q9}"�q�Hr�<��D�g�f|J��O�#~��)W�n�<�#
D�#�}S[0��� Do�<�竒�B\3�Df��p���yrk��m��Q�S�ŻU��X�(�ȓL̵`$��0pQ�S�n��ް��ȓ1D��ж$U���i���F<P����ȓ-�����Ю�R ̞<w���ȓHax�K@�9��	�  ѽi�v���$9r�Ksn��7&�!"�ȾN���@w��00"D�o �-r1�ݎ0C`D�ȓ7(Ԅ[�nW* ����PnA
.�i�ȓ{����c��g�
9�f�څf˾؅ȓ|J��a�&O����*�$����x��ӧ�K�>���K��)d&H�ȓ����!C%b�PQsep4�ȓt��5 �^�;��Q���Mxj*��ȓ:@jV�	;^vxأ�j�	?�"x��O=&�S5��-;�$�Ce���6��ȓQ�L��4J����C�ʬ3�|B��2�d�� ���}S�E�t��C�ɹ�F��6���5�xY���6�FB�I
Z����d�`����K>�B�ɂf(�0ؤ@�3&ԝR�+F�O."B�I������P*S7���<sj4B�ɮ;�4d���L�DY����vB�	88Հ�#��YRd��e��v�C�I )�H�2��F�g�t��p��$0��B�I�+O�����-a�N��dX
`�$S	�g�Ksc�
[��9�@�R�V�뉖o}�5����U=f�)��1T	R�	  �!���9 ��@�F$F��鱊�-c�1O����*��a�f��!"�'vJ�.O��q�f��'(�|�ȓ�)А �=F0F4wA�v��E�����=G1�$лR��?�' 2���cZ�}	�e"q����	�'ݤP@��>\���A���.0���v"
Wx�̓��w���퉷X�V�d.L�R���V�Q�<�����օb��/N�$m�6��G�t�nM
(zD��%�7ݸ���B>	��ˊ��r�p�D�3U+��%��p��c�@����%"2p]E�D12����"'�%�\q���Q��yRC ^�
`a���(�~\BM�� >�5�U��%���I�u�j�Y��L<9����3͚��-�"ވ����vH<��kT6p�i���I�y��)s�B�B�LyCЅ��,ٷ�Λ�p=qBk�ۂ4������QpH�qX�q��O?YJ��Pj�6`Kn%C��P�~M�G
Կ.��Us�^�yBo�4��ہ聉5�x�W��'�ēh�����I��)٦���(�� ĕrG�Ϗqp�RwJ��D�d��V"O�u�VoIȲ���*νn���g�h����Ԭ���?�f
�rs���'n�`��2w���ԯWN�n �'x�D0p�K w[��qP�g�xU�`�I Ю$27�Nʉ��I_>�p9"�7fr ��Ԭ�5I �󄖷gv*�äL�K��4|�T��sm�h��̛p��u��T�"���F.���
���+t�>��<�ȗ�v�4�j�K��h�:X3&��M=~����Hm�����"O^�!Sk��-����i�Y���{�U�3� ��"�>��f>�gyBk���f���L��MjTiD��y��B�j�h�E�J�ܑ��?a�&	 \f����b�P�"��W�^t8���Bg!��ǁ���BC��{\���&A1[!�DG���!`XeXR9�q��=!�DG.ѠD��I� ���9!
�4�!�$�(��`ǰ�,�H	F.N|!�d�4P�Q!I�>�r��(�Ao!�D�/8ͼ٘����p�8၈Z�#�!򤗳6�D�v�a��9IV�MR�!�71K�M��
�**8���#gʲ3!�dB;O�.U�4�� �b��F�l�!���)O����$H�3���Pr�Ҭi�!�$ÁR)(���MT:�\Ģ��4�!��0��@�go��,"0��/�!�X�\��`V6!X%�g X�!��<75$p�/V�N��"n�I !�DA�͒�Ӑ�]�K|���'�t*!���Dbj�Ñ@=P��j�`P�A!�dJ�})��(�MN�Bc�͋s�!��Y��f�H����0��B	C�!�D��N����B��9	���@�!�$ ��aR� �&�Z}3@(�!��Š:*�IPeҺ�
=�f�!�d�R�D�����+B��A0m�::�!���R��t�sS7k,|��L]H�!�Dۤ	���A�.�=-B��+	_�e�!�2�T�(&N�tG���0	Z�>����F�`�0a��*&D�ɑ����y����h�% nL(��Lш�y�!���Yb	�U�����&�yBN�5<g���ҦX�C����$��y�ND4S���J -�\�7�܆�y��ݱ��"n44������+�'�b ZcO�-\CΠ���w`؀�'c�!*Ղ
g#^ͩ�f���'"ʄ��.�8+��lBÈؽN:�y�' w��J��Xa�Q<9�F!��'�L���<UДs$�ũ2/�p�
�'/؜[H�A���SZ�����'��e��n[86h>��qI�x��D��'��I�@�~�x�tEU��#�'���%Dr� ����|>P�;�'��p*Db	�O�f��ƄG�hC���'YN���f�b�5H�ܩv����'
4�f�. �>�m���
�'7.���� Kw
q�	�u����'�>�RT�Y	1���Sq�S�k��$H	�'���Ҁ�3O���(���:lZ�j	�'��H�#%O*���_�lH4��'$�D`��Ru0-B�lK�fD��q�'h�C��*S2�dICƯOrF��'�*АA�Ğnv���BG�;�v��'cb�@�V�������<w�Z�'��l��[�KY��&f��g�F����� \���C��ک��������"O����UW� [%���Y�dyB*O0ip�Y� m�i)��I��E�'��zB�T��0��$��s�(H�'���٦d�T�F����mQ^�c�'�|I�����\�y�V�P�f����
�\�q�v�M�D�-8��I+�+�&m�X#�ծQE!�Ą�{�ы0G�W���Ao�=YM�'��9j�	z����)N;嘙�4���&4��MT''(!��
�?�����1�j}���7q�����c*?�&�m��>�O�-���NY���{!��M�NQ�QO�!�҈��|��ӢR=vi�1���')R֕"�'�9),݇�	�."x��(]O�����&�_ �?�1��!wy.i�C���;�x�'H��D�2�> !#������_
�`��	PmbF��>/ $�' TI4�ا{i�@�`W����h���̓���(��#RQS�"O�5�ޫ>e���A�C<1�H�^��C��*0,<1����U��3�
-�٠��>y��i��/[�?��9���6A|lSa�2���I@!C�l��!BG���#��l�0
t�@f8�����o��f%I�O����#�Y�6��il�$��J���؟�y{"�5xn �"���U�"O���*��q�)Y�� �L��cf���@B�NΥ�uK΢k�����9�ʡ�#.�(
��[�cF4@�v�S"Ov�0ܓx�� H�E)-�PX��3u�=�'hI J��bAg�$gܒ�(OF<�%V� =��O�q�
h��'��!W�A$JP�2EJ�@r���N�6�u��	�qM�p��h�X�p����kQJۋ8�~��Cn]�r,��?9C:I��5|:���8Q�4P�'@�eJ�qU�J�� 	L����J|X��L
�X1*W6lg�<`�$�74C�h��n��lY�Ʀ�Nx�?�a�w���M�=$|�Ò��,7�N�J�'+|��w�ߓ)��HFۥ`�$Jf�֙xw��B�Lsn�arV��"c+~��'�Q�'iޑAgS�H�][\lP���F���"e֙�$����8N
	��Xd1�uKj�� ��(@ �	-�p>iԮ��+��-�#�®p@
Bd�<,±� p�`�t���~h�8�ҡ�	�m!*���·ϒeYr��Z�!��� E2,C�A�c��-[��M��,S���6�  S&J�1s��4Ɉ���O�>Q�;}�\a!�!G.�J�ӯ
J&	�ȓ+,LC�������P��� ���.4HS4�ڐ'	��a%��5Bz��2AB�G���<Q�D70��9��MĘ%��Xb��[��t3Q�	�D,�,�"��=�.���%ϕ��������o#�X���9mT�|APj،�p>م��#+��Ӕ�69t��2'C{��P|�3��!e1	qg\'�����+Ŗ��iɡa���U�<r����V0y�!��\T�Y��1<I���/��Y �������wC�wO@��b�<§X\���l��D�EQ�&Ȫ� �)�C�ɘ
L���6�B��.A�ndK�팅&i�m#1k� k�D��oF�����Z�'�z�! *hU#v�Ϥh}X�z�c��X��G��d�b��X�m�T�j�H��(
I�V�n�M�fn�l���;�G\�y��d3�$b�07�[O.�|��I�!y�%�w�)�'VV�l+���Sg��0u� � <�ȓ����B?B���2iO:8
���Q(@�3��8���O��AF�4vl�	�E �^�E�W"O�D�V.[��̲aA�kҖܒe"O>l���j��+G@I&N���ke"O���i��;�ڱ[����v�^���"O&�Jé�*H%: ASO� ��p*�"OR�"UG��5�a�ɕn��=Y�"O���Ҕ^熕�� YL��I�"O�5C��
0ON��i�!9��@�"Ol��/��k�p��k��r�c"Oj���.�,�уL�
���"Oj 0 ,P�$�ґ3	#?jEs1"Oy.�������CӰ3�A!R"OV$�&��	u�X�'ǲ@V@�"OfȰ�W��M2$A�^�5�"O� �@p�o�)Rsν�C���8L�"O�m�Q���,(*�W:SQ�y��"On��$m)cSj��A�9@|,�#"ON�F���l#����0�"�"Op��U��XC啻w�0]�"O���C�K�L:T��4����$X�"OH{��L�jHJ$�"-��Ţs"O��%�f.�\�  	"3z2�7"O��+���)��ʃ��D8���"OL1�0	\�4x`�鑜���5"O�JR�M�i,8���4v_�4�"On�h Ɉ0��%�v���AHZ�i�"O��Z筒���r���8I�j�"Oh��6�)]�5� �.7]<)�7"O@�s$@C�C-�H�F��_%���"Oj�BE,�=e �pSRA	Ap.W"OPYql+7�T�gI�.UhP���"O�Y9��� t�dQJԽNG�c�"O��`�d�')�hlKP��P ���f"Od�0�M7A�dU����6h�f"ORh�� ǁd�A��N��8Ӈ"O�xvÃ���7"��A8�"O�Y*��ї<�,�I�'��z�"O8�B��������	o���+c"O�p���Zo�L�4*B�5���a�"O5h�]�F6<�ѫ�,,�����"O�e%e�D9�J]�K�R�"O�]J��Y��t}hQu�Jq�"O  C���?�Iy�S�6��@��"OpA#�D��r%$dG��0�ܤ8�"O�\ Q�՟tV��d ՜<���4"OI���`���e(\;l���&"Oꔃ�i�-kh��%@(3�> Y�"O@���!IX��i�Վ~Od��E"O���E�
�4rf!b5)K�b<���"O����8`K����'�@�"O���"�HbL���Ӱ�u�"O��e 9r0~�Aa�l���"d"O�ys��#ig�ո�a��A�
���"O\E8��g~hq�DO�w���h�"O�M���͑;Bp}Y�w�~�P�"Odx9��EB���A.د}.�#�"O@ ۰*7�)+��KP�	��"O��k�(�2w{|x�A�Y�(H"O��A��_밉{�T7<e�	b"O扩T՘>|B0ĤAh��sD"O�؀��ڭmc�X��
1dUƝ�"O���! �lGH��&^�C��"O`z��ͧ\���B�DK�\K����"O\51��Q
<Z�հ��8h=��3"O�Q��@�Y h�c94*0�"O�,�&��"mӐ�S�L�;�"7"O",Kc��]2��)BJ?>�!I�"O���%�L)A���1���)8 Dр"O��c.�|d�y���0k9�"O����-~��t�C&I����"Oĕ#� @�<�J`"�D��y�"O�mB�b�)N�x�ċ�"5��s"O�8�+��1��탵��+}���
"O"���kȔS殁�M�m�hY��"O�X�P��J��B����eEJ���"O��X���
B(yy"��7@\ɵ"O�`�`ő��$x�,F�3:�(�"O��h�"���b�L�#C��"O� �+���F9��Z&��G��4�6"OF�[@F�$b$(�dL�0��0�b"O�e��֧0���p�	�.���ж"O�����Ϫ`�t�Y2ʎ�H�H4@7"OZ\����5���B�u��5��"O�\�@ ́)���:F����`E�%"O��p�ΊI��!u�������b"O�ɸ�)��M�� � >��H�"O�UqԨJ/�|,�&흆�T�"O�$(Fˇ�$��x0�] !�v"O�x�#HB)\uP���0��0�F"OtU8�S/S���� L^l 1"O���΋5B��𹦉X�:�['"O�h� ȱ|�� ·	�!Kxp�:�"O>d������, C("���Q"O���B�ő"��p6�J'E�Dɂ�"O>� ��Ҩb�E(Ul�IǶ8�"O���������.NUl��d"O�My`ď�z]R  �'�>#�a��"O�ċ�żg�<��dF��\~�TS"O��Q&�Jc±R5��Z�%��"O  n#q�`Rf��DPbr�!򤔓8!��� B����E%�;�!��)/�z�Z���@����J�}�!�D�F�P$p7NتMSh�k���{a!�Y}�<�6%ɺ��pa�j�L?!�ǫ*�ab C�2S2hDȡ��Q!�%�!��"�7��Z'a��!���-�q�k:���PP��!��uc�\XÌ;S�Ū�L�!�ę,6��%�U��+"u��h3hU)%!�d
(�JVl�1��xQ��8"!����ǧu�t�c�ۡc*!��1
�^ysF��Ϙu���@�<*!�Č�T�� ��$�8r'Z�8s!�D�6Fx<Y�Pa� �\-���!S�!��&$*��^%�Yp�O��
!�D�$<�8���ÉA�~tsՎӥ!��T�<�����-D�,:�͏6�!��?Pa6p1���d����54#!�$�-jD��(�i?��ЦM��
!���|��T�}L�Ǧ���!���u����B-ڽt\���%Ǆ?,!��b��=@���}In�B�ٰ!�d�g�(���$m�)�u�W�l!�DP
e����`�wM�Ă�N�M�!�dĹt���yǬʩwHܓ����6^!�DJZdp �6Cئ	��[�<3�!�Ц*P�r2
	���hS��
�.�!�_MiNa�Т!8	�P03���~�!���6&���C��)�.\"��/��S�1*T�(C&��
�9�	L+�q*0��.�>:H�ճ�$�~��'��lX0E�.�ɧ�RyR�<(����Q*�(����M��^8Av�=B�bUE~����3O��:@f�2G�5(BJ@y�8�tjP)e�,�O���	K! ���4<
�m�I�Ab�u�"0�$Ӗ%����iS&����I?��H�M9O4�'�Ӂ�ۤs���iM
t�lqJ�BS m� y0 -P$TH�	*� l;�#�?㞨q�#@�P�F���$Y�I�( �De�t @�)�'�D!��i�-���o.�5�pm4�P�?a������l�у�E@(�����	y��1��>	i��pkr�;��E�s� �4���E\���u8��OB��'�@�h�����0|7B�v�����Ks�N��1H0q"��b�4T_�y�q�	t52>�N)%>	�O�慚 ���,�r��`Úr����O(	3��"�7�7�"V�a�T�_+�",�"�}��ȖBKT�A��
�� P6M���Rl�q�� �~� ���헯�ܩ��d��2lv�B�'�|�nڻU����B��N}���ߛY+T��6Έ�.-B��Ï~���m�
6��9ąhy
ç,�V�S,�W��Lx��C3tH��I�=İ%r��O��O�ͣ!�T�Z9�,�2��t�@L�
��3NA�>E��O�hD��$��q�
Y�CϏ26��I��&�;�a�D	��L�]2G>i�!/�(��'[ṽ��4�F��7#[��3�^a� E�7�F:�&ON��O"�)�e�F��՞Qy¼j�	��r�<��Fx����*s������2D���g�נ>�"'HK�����@��G��"�-ʇ�h�z���;D�܁Q&��d��! ���V�qd�8D�8P+����GBٽf6�A�,,D��i�gJ, *��Z�dإe�>�W+D�H�Ai� �v�[�U4m�^8�EE#D�� ��Rh�u�K_ Y�h��p�!D�8b���(�~���Ú$�6��@a-D�h��oҏn��I	�j��*�	.D��Q �[�/��h�
�d��K,D�����i��HJ�$uQT )b*D��@ҡ�w���)�苜I;L��o4D�<�7�PO�dL�¤˳v� $��1D�ta�؝ER�1�Qk
�&Υ ��.D��P��
)R��d�3M$
����2D���A阊X�|8��[&�m��0D�X��B�}�P����*<�R=���,D�`b������@=L�L���6D�T�0�Ʒl�6�yA�t��2�W(H�!�$�Ebz��)�W/��gg=u�!��$���9��]�A	��ϳN����E��b�h^j����lI�~|�ȓj���bs�T; jL �`�@�"J��ȓA�XH�k��i��=�ӣ�
W�i���,X�$�[��0��NCR<��A�"���X���Zai�v��I�	�,[�%��J�A� X~���x[��:�-�Y�̉��M5m��|��E���CFZx�:"�V=2�ȓ=$@be��= m\2'�Z�䵆ȓM�pr�+
�LE9ڦ��R��ن�?��2%��5-�A�1�Wn���b�Aj ��jc<K�I@JN$��O;�P�&�ݩ`W~���`�s*|��}�-�TL,c�y��.Z�	���ȓ^V�H3��N�lۅNK�<� �ȓ^$
�pb�_%���@C��¾-��:RH刟5ICؕ����0/RE���2�2RgG&~�~0�b��${\�ȓ|i҉k%�8w(���`x0�(��?W ٛ�#��o��I1��A�i�t8��v� �-���4�TcX�XH]�ȓw��\Ӏi�+qR�1#I"3�0�ȓoY����ya���'C�JmP��ȓu@�����&C#�) ��G$?�r���H𡂄
7*>t4��@]�&�~9��"�	2�n�I,��c� �bjt���ؚՂ����{n���(��ȓXb��a��ؿ=r�sP�_ Twnԇȓ,��� g��v=(E�9". ��h"VͱE��$�ް��mZ1^B����P�E�\�C��`� ύ�.�x�ȓ�V��d��(o�vY�1.٭�`��j����㡄�qI(�`ai�$i�هȓE����a� @U��D-�y��q�ȓsߐ�c')�y{��R(�]�T��S�? �� �Nm���z��ϮaGH�RF"O��j��N+��(�	S�b�H���"O|�(�S��.4�0���''܄�d"Oc��,�*���a�<�6�rv"O0Z�-5ΐ��'�X2&i�}Ru"O�<[ 	$O7n���՗Z|*���"OX({��N�0�(�!�+�6H���P"O�8�m�"��������Rȹ�P"OD��#�C�_v����M7ֺd;f"O
���ٟ4��<�F(oW, Q"O�E)�/6�x�ZD$�
A8��2"Ox��'LΚg��A�O>��YV"O l�I�P,�1��7���b"O�Fc�U��L!��@:ꐕ#�"O AP��4�f �q����<��"Oܹ��䌃h8*���H,� }��"O���%eB�+ZL�P悋CӰ���"O����ϐ�N��$�#�����"O!X��N�Z:!4$�q�Ȑ�"O̪���	�>|�d�щl��A"O�`궩�1Y(�Kd��[g�X�"ON����H?���ƅ9<:Lܳ�"O��ppGt�f�1��_����"O�H&�K�a{�W9jl�3�"O��Q�gP+3#:��'��yH�q�#"OZ8�5���	kn�ՈS4\(c"Ot�9�ʛqb�)[��OF*�d"O@d�3��7�J`�����8"OX0�)��,���KR+�������"O��8e�"]�ƈR-�;�J쒱"OH�z�&#���K`���S\$�"O2�Y�jI�%��	�B�%AI.���"O�U���h�4���c .F�2��"O�x�#E!S�����,{~�m�T"OR���@�og��2 I+x4QpT"O��K��O�JD�8�W	ߥ`�\�p"O<|����0"�s$ț�BAt�J3"O����F	<85����ŋHp!�"OHx�-� B<�Hr]� ��q"O���w$�Q�eY�6m]ڴ"O�Y fE�K�X�p2�2v�q+�"O½��E���d)T�Wn�r"O}�Po�u>h��-]�+_�m��"O��sMɔ��tZS.�0+9���"O؜��D�x�CCc�+fʊ��"ONё�m	�C�����S1k�H�IV"O d�Rg_4V����b�Z�~���"OP�� Y�����'P��	"O�9a7Ǚ�.<�0�lH:#�Y�V"OB�A�bݵe�p4ѕ�8Q1p(2"O�̃�aɥ'��z d��B�K�Ye!��91 ���+ߦFBА�P@[�!�(f�D3��@>$���`% �!�$,T�Q� �D��FMz`OQ<
!��=_�b���$v�&�"t��1L!�C�N���Fą9v�(�@d�Ŧ�!��Γ3B�p�SI9�|!�iM�h!�V�G�*uA�(�=.y�Z�.�>
�!�d9T�5��eԶ|`���h�!�ͭ;nJT#T^S��0+��P0!��Z�S�5�U��%9�����l!�+%�vt�B��(�� 	T�W�U�!�D�MJ i"���=8r��qk!��+���%�X�=��9ڦ���
��� zMs�"\�g����3�^��~"O�LB�(�	h��U�V�F6<���"O�i3�d�P��"��Z�m��`�@"ON�Q˘�/�6���F"n��y"O���e�ҟT��k��S�^r�X�"O(�Q��*�*�c�J��S\��s�"O�ro،]Œ� ��R�sE���"Of4�b�%�h�4�~:���d"Od���Y�T�S���d)��"O&i3����+�~����  Y�nݛ�"O����ם�0��Ծ7��p"OdH�B��H���cd��=Nʀ4��"O\�K u8��h��+�`�5"O�KE�.0i,��G?h�^́`"OB!�㚥H�p`�V��S��X�p"O�DB�o��JKXAP�n[��K��7D����`�v�d�B��ŏ6��9+��3D�!dY C�J9�'�	]��� L/D�@� ��m%�:��T6�2���-D����C�̅��D��*�b��7D�ppeH�/]��
��F�cE!D�pH7 �!��a �,,���He�#D�tr%#��.����K"G]f��!D�Y�˗,a�Q��(�0�u >D��8�L���A��?�jH�#�<D��rB��K%�x�v�0G�>��"�/D����sвj��¥%0�p� .D���G@֜
M<���*�q����"#1D�\Yu��
d���Z�t@8��:D� �b�V:1����"o��q8D�$�vO ����UoV�cU���q
6D�l�r?G�PI�!�"��<�"o3D��!&J }�rā��9��� �f<D�D�C)�^O��r�T*�84N-D�,���T/&�0Y �呬 ]zp��,D�d�F*-LP� �FH���-D��2��R��b���Mv���S�?D�P��ˆmd�s�l
�|�PeY��?D�4S&��5d�>A�$[�6���1D�,I�)w�pd�q�W.�ָ9g4D��JS�[�[��E3� �K��H��h<D����G�9�)�dM|1�''D�TbҬ�xŨL��혥5�f��)D�L�Ah^pU���0	�=n\Ve�RO<D�8���Έ!���S!�@�";Z���9D�2�@�# F�(W�S���#��<D��s�m%xX|!M�P#�i<D�T��I�xez�AK�/t�	���:D��I�ձ�BH#�S�W�xE@6�8D���b�ڗ�<֩�N	V�r�;D���Wo�7;���Q���Qƅ&D�Գ�L���⭊�zV��%D��j�-� w@y�2���d48y�/%D� �2kкleJ��3�YM���#)D���7@�< )��� �� �;D�;aHN�|O��bBJV.0�"yK�K&D�̢'K��A*��S6 ���JS�7D�&�B�y��S�*��	�>C�ɲkVҝ��c�HuX��ϋ�jC�I���	�(�?6X ����B䉍�r� C*� {\��*���B��+7vt۱�W-�(в%��NF�B�	�\Q� �ɋ�n�b5��
��C�	i���jFi��!�P,u�C�)� �ݳ��T�{j�]�P��)"�u"O�5�r!Է]�&�1�g�>*vP�"O�����7�������$�tzu"Ot)�� ��g������'�� �"O,�����7q� pC�9i�	�C"OĔ�c�����ԏ�"ML�r"O�ɚ!"`f���Gt>DE�"O6Q�<;�RYPg�) 
�3�"O���D��I.,�RE����	D"O�a�0�OEr��Y����T"O�XP�MH�L��m�)�%�)�"OV9çg�4+t�����C"�b�I�"Of%	�U+J1��1gNI��rD2�"Oj�30�\Z|4�	�ظA��<�"O�T���O�l�p�K_�JA�A"O��a��b 
�h��=~�x��"O��   ��     �  I  �  �+  d7  �A  �K  �U  y`  �j  �r  >~  �  `�  �  ��  Ԡ  �  Z�  ��  �  1�  }�  ��  �  D�  ��  ��  �  ��  1�  ��  � e � � �( �0 '7 j= �C �C  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!��I\���B[��|/,�X.�V�H(��iKN�q1DN�l��u��Q�t�=)�O��~��%	@�D��ĉ�5	 ���C�<)@a�&t�wE�e_$�kf�_�<��{��'����Q��"w�t���جg��u�
�'\����1(
d��ר\�p~Ah�4�M3	���x�3�h�e�(��r����l�D�16�,�ʇM�J4������A�!�$���pň'7�f�"��
���XF{���D0ևQ+C@����,�I""O���E؊p����dI�tEY1�i��c�d�S�g~R+>\���·��@*ad�p<y��� Za�A*� ~"p�BP 0�`�"O�IJᝤ� ��C�^
 l���'i�4O8�x��\�z����H�$k����"O�yJ�/}i�����3��E�e��.�S�iѣiX��&�k�j�׎�<!�$��{s܄3ե]�K�l��M�!�D�-D6�b�.�4(]��P�Bf�ay�剳� ������`�ӎ[�\���V��x��˭Lo L	�E��ةҠ7�	{���	��������(c6�H�<
��W+1D�耖A�)Q�R8`��Ao�4�&H+�I{������Q<�&e����4'F%qd//4�0x�(�I�H���̱Pr���'_u�<yD����:��B�F�ʈ�SJ�v�<Aw	�!0�`�s��E+,N��+Ng���0=���7�V�{3��*���Ȣk`��@�=���Oґ�㧍�y�FxCQ��3�y�7.�2�1��+xnBxˀ떦�yb%ʺt���l-����:�yR�5.~H����9]��yߚ�~�|��'��0E��{-8�dV�_Z4�:�'�8}K�[�3p�s�[8ڥ���'�d�Ox��q�[���2|D� %L0n�!�K�\X$ݢ��ǘ" j(���z!�d��v����,Z��Sp㉾�!�Ė�N8AJs�0.��53�B��O�!��<E����0����u�0"�7F�!�DEA�H�	���?0�2|AFBO��!�˜M~� �
k���@�R0!��� ?HhC�(��7�"�k�P���B��H��|A��V0M�i�g+v�4	��"Od9t�Ѵ{Gi@���<}`ı��"O�ᩕ��]�=�c��&'O�5@��'��-�r9�,8!'N�9F�3������­ɒ�0q��"I�.��DzR�~Z�a�J#�؉�Ȟ\g.!�1�C�<Y��cZ d�3���1Q��R�A�<���Q�.�����C�	NPEK!�	{�<AAf�"ojN� �'K�\�(�"s}2�i\a}��N7?��4rwo՜jr��eH��p>a��>�����^@�)�g��b2�Ug�<���^i��+�@�	�����_�'$ў��;\��\�s�FVVv��$� y�<���I��&o�`�B�[;
�L�=J<�����;�mjS��>�%V��"h+!�d_x��킜*��hU����!��:/n��T���?���6�_$!���O\�x��*� �2�y��xQT"O>� A#�1W� ,�� �!#��i�g"O��5I �v��0�٘1�z( �.AzH<��F/;(\�6�ƶN��}��jSz��hO�O�p����0Ua�� &B�8-� q��'f�@
�n�n�p1*�.�/*�@y�O��ąQ�?QI����&� Lth��Hg�Lrv��A�ar�O0æF�V7*����N�5��S�'i!�$ͬ/\���Ɂ5s!2�P%��K�a{R@8�	6��Eڣ�H�|�ѲN�u�B��L�d��"���6m��@:��C�`0���#.!�y�a�I���B���@�k�bN�&�����[��<��T>�
���\���9�Ŋ��jL3T�9D�4r��e��,�G��*�����+�ް<� ℸp}%��%E�J�%IU�<i1hA'u�&���[6�6�B�P�<� 
uJ��ܚ�
�+���pI>��dP�XF{�igqO�u�& K#����A�2pM�C"O���"�:���F# G+��0�x"�2���O���$�S�Q�T� ��� �:0�'��|��L8{c�1��)��`J��'���ɡ����L�L�q*�+�y2�
4z����,�:qJaK(�yB�R�:;~u��4l��$�0eŞ��>Y�!�<)硟0���	����J�Af�<��D�,R�l9��E��!i���d�<��&�TIу@�6�S�V[�<a��r���3�Pn4bLkJW{�<)��3uDx�V�ŋ0E�����y8��Gz�!I�}ҕpM��
u5��yR��=~),��G���Z)񁮒)�?��{�O���8!D�t��0�(��R��!�C��C�dE8TÑ�g,�qh.��ڴ��?C� �'���YZ8+we�n8�l&�l�1!9�68"�
*L��<�q��O��=E��ێRn����ΈJT��7M�!�Y�.?�}��ؼ-
��FY)C�!�J�[` ���b=X��;5!L�z!�DR�{g�9������ђ�/A�<f!���^��Ykҳu�h�Z2a�!�$X�vy*�F$ز ��*�l��u�!���w���e�H7�ʉ�v.ߛ^�!�$AKj(���kA8=�> �N��9"!�D��w�:���E� ���L'��	A���)u�P@b]�FtZ�)rDۘlkBC�ɣ:I�Xh!
O�vdF}��MX�X�$C䉀��/��0(��Q�~힡;c�%D�k�o��)e)��Y�&v 9Vk0D��qw��8d(��hi�ܙ��I3D�HZ��� U��QS��Q3ri�bc0D�h8C�N��@��j�	UV�Q1�0D���F���pX���ɷM����$D�0�T��5N���.��.�����4D�,˖�U�:� 	)$�\�>o4��!�.D�4�	L#=�,����qz���b+D� `T�.s"D�(֤حNY<d��*D���)�,#�ԣ�☢j�+`L(D�0�dFF���9���Ӎ!��Y�L'D�@���9y�����[�0��ȳ$D�X�ũ�?z�<d�C�9)�48b+!D������5��x����ꂔ(v�)D��J�jD�i���F ,�1�FO&D��9vfҋNܒ��v/�r��	[R�%D�,�t"���\�f޽ �Ui�E8D� ����j��㢛`Pـ�a)D�����ւ��0���W�}���a��;D��a����b��h;9��!h��.D��y�
0�
(���w�,ȸF�*D���(�_��PuN�8��acfd'D���Y2UVT��
��jC���L D�t8bd��:#������^�!9)9D��@kٛڕ�!�Ĝۦ��,!D�h�$�ߚ!���X����S�+?D�gbîRv���틑\��ijw
3D�x�$��6D*�(�A�d���[��-D�l
nU�:��ёg�^�5���ঁ,D�P@�*Ϯ��`ZөݿD��*O�`Y$���2@����c�*쐅��"O��ġ�#��u��!�	�tT�"O*8aԯ�4fx
����)�651�"O� ��(@EЧ-ʒ���LR�����"O���eP�H]􌁷��d�Tջ�"Od�@�-�C�@��0b�@��:�"OB��S����XeN�N��8�$"Ol���*��#��B�eN�
�0�#��'���'_R�'!��'���'�r�'�D��1��+�@�Ȣ2�D��q�')�'�"�',r�'U�'�R�'
��81NS�W��A��Dv�tU���'���'���'��'���'���'�J�t+�9k0�IPaT�Μ9�'�r�'<r�'�"�'}��'�b�'�Fp��Å�U�GA��~�Z�c$�'r�'0��'���'���'�"�'9��Z%��hX=���+H.�*b�'1R�'2��'�r�'H��'Q��'R�d���"q������>j7�e�T�'9B�'�"�'���'���'=��'7����FGz���L�94�t$���'t�'��'��'�b�'�R�'z��y��ȍbJ�Y3o�#�e��'er�'
b�'H�'�r�')R�'kd��&E��4��a�T/�̩&�'M��'���'U��'�2�'��'C�n��p����<��%m��2�'p"�'�2�'���'���'�.�T��kE���<�[w��!r�'i��'�B�'"�'���'���2�b��p����W��*h�'��'0��'���'U6��OR�d��W�,	; �Y	[�J��G�R��`L�'$R�b>�@���'W�Z����cl��t��$���� Irq��O�Ym�_��|ΓD��V�J�8>���Y�@���|լ6m�OvI[F}�H� 5�w�|��O�̥S$�A9H���V�L17���yB�'���X�O�zŢ�-�e������A�'�f��}�ޅ	��d<�S(�M�;w��=�Ы��i~���C�Yt�r��i�x7�x��ԧ�O�xI1r�io�+\��BOZ(��C�ܻv��Ĕ�z�T�"�g�Tʣ=�'�?Ae�Q�wX�8E�HU�d�2J��<q(OV�O8�l�%z�b�( 3�Q�&�+^�}����B��j@�	��M� �i��D�>	c�W;�V�@�D�$Y�q3� �J~"!]Z�1�e6��O"���܁�	�<��9�m܊
�8����'sg�'*��"~Γ~��DP�+N�=����
�G喠͓l꛶�6���V�a�?�'*GԑX��V�X(�`r��&M7Ƞϓ5	��/kӲ���2φ6<?�s�W%q?�@�dw���t�&qq��]���:�M5��<�'�?����?����?�K�~X��fH{�|T9���5������`
k��I��X'?�	=�b����B�4�&(@f�>�X�)�O�m���M[��x�OG�$�Op�����Q��AE-��IԦͨ�LP8�P��8�Eղ=�$鯻3��'�剺/�`�@� R&�L��O�e����Iğ����d�i>ٔ'��7���3��$C,]A>�9�ǐ�.j��3b�O�g��[ۦ=�?�$W�XP޴i�� v�v�BWI[+9xLi	�ƞ� ��=�v	�;]�:7�w�0���G�hy�� �U�'����w�$qyq�ș�����S�H*�
�'"�'���'��'��jԃ�ꐸb���%�5y������O���OxnڿT��Ԕ'�47m'�d�2�,�P�!tJ�9ipH�E����@}�jm�`�oZ�?BD����9��?yvN�8PuP�"O�e"x-Ȃ���$�ae��-F(d�N>y-O����OH�d�O`��JT�y�E	���5I���O|���<���i�d�9�'Hr�'��S-�	Zp흡z�f��O�J,��f���4�M�$�i�O�i�
Q��	�;+���a��T��=�6e�o���b�\��"e����u��4��"25 �Z�k՜��+
����O��D�O���<�ӽi�*�#��
�7Q�lf ��QG�x�����$�Ŧ�?Y�P��ٴIy�1(�-o�b�j���$Jpʙ;�i� 7-N{��6�j�L뢌�7@9(�w�ƚ_&q��?��� �H@��G�9>����D��m�*O����O����O����O@˧�2Ţ��SKv�+�M�U���{��iĲD�C�'A2�';��y�y��NP�����67��8�c��G��=l�-�M���'M�i>���?ٸ�&�Ӧ�̓,�@�u��Mּ83	��`�6�ϓHw�����0�j��N>�)O���O�=#dmϻ4"JI�uj�-�	*fO�O��d�O��Ķ<���i���P�'���'4܉#"�i�H���� 6������D�}}"�pӮ�lZ���`����t*M.z`u@�d@��ϓ�?١��s�{s ]	����V��D%mݕ�8;�����¢!f��J�j��)@��?����?a���h��nPW-�x�u��h�TQSbD�2��$�Ҧ=��:?I&�iU�O�N$l*�!����
���%���6��DT릙�޴a�����>O���8Ma@�Y���%[*������ntP�[�t���5Q!��O���?���?����?!�Y�6��3Y���+��2i�,O@ynZ/96�	�<��o�s����+ܥ>A����x`:�;F ���M����4yƉ����O��D%�;z��I�D!�y�t�S�KI|���?+��	�2K�t�.ם�����d[�
��d��OF!uo�钶�+U���$�O8���O��4���z���yRn�39~V4r��Q1�xp[�/N��y��f���Y�O�ml.�M�'�i�>�H@]\��e�WiļR"T����ׄe!��7O����
O�:$Ѓ� ��ʓ��&Hu�? �[��1ky�����\HC�M�kS6@�f�n������Ȋ*8�w�?wA�AO"� ��&�$Y7�PR�� ���X'��WڰM���'�H��"69�d�
�g�`��1�DW�a�@*�p�� �68�5��F�a���{�0���P����ƀ4w�P	��/_�U���`/E48�7���q֪:t�η�J ��>c� �{&,X�I��[�-�^@�P����%���p��\�5�dЈ0o��Q����'��'�����E2�D�Oh�d�� ��ˏ+U0r��X=7���p�A0�ɶ@��|$�������I/�؃Fӓ �Z�Ѕ��42�iI۴�?��J��b��O$��:��ƶ� ��R��e c���*U�X�T�,��� �ڟt��ޟP�'��1���0�&aP�O�1%=>ЙTG�t��Ox���O�Oz��谁�n��h��!�L�j	�L��B[D��?a��?�.OҜA�e�|:#&וd<���j�xt���1�
G}��'�r�'U��ޟ�	"YO��P��-��7�jq¦,�l�'�"�'WrP���`�U��ħi�(U B$��+��j�dQ5<�2E°iB�|"T�xc�>�ӭX=��6fƍm�FPf���6��O���<q�懯j��O�"��5� ]"F�H���HP�E�j��C�#�MC,O��$�O�-��i�O��i�ūF���fxtY��I�@H��4��DV9 �bEn��I�O��)�d~�T*��t��A�lU�c�Ǭ�MC��?%�
-��?��3�$h_�Ÿ_�d�� �o��v"�G0&6��Oj���O��	D�i>m��݂q~N�p��m�v�d �.�M۴-q~�_� $?�	�����~S0��eRf��(z�BH��MS���?y�;�@5I �x�O6��Oy��k�}|�����0"���dV��'P�ˌy��'7"�'�~9���ġM���sR����*-��"k�x��.;A��%��͟|��cy�ĆE�8�Pv�H.j�{��Ś;(x6��O���a���O����O6� rFy"D��!Z BB�J�a �5�abE$6�'�b�'n"T���ݟ,����ZK�}`J-���Z �#��b�8�����Gy2%�!sf�0a4��瓑T����ۺ|6��<������O��$�O�Q��T�t{G�~G�A�ߚ��mv(`�j���O`���O˓B���_?5�i���3{�(�A�	���R`�7��O�ʓ�?	���?�s���<�,Od�8�����XFnE�v��5�I4<r���O��H���TR?)���P���Sq#�<�(  �e��Hc��0�O��$�O���E�}\�|���4䝜rqN���� 3���yA@�'�M�+O"��a˦Y��ޟ��I�?ay�O��S�M�����:�0�@��-Λf�'��`��y��'4�]�'0g�U�rᑊA���Z�����мi>p�0$eӦ���O*��v��'��I�j�j��LZnM����0ʊ  ޴Wb���?	.O�?��ɨpu����=*��@��A[�C_��ش�?����?I�$[�-��}y��'H�$�?qz�!�%ٗg\����G·
�O�a(���O����O�M�J˿�H�0t�z0 b����m�	({ ��y�O�˓�?i+O����<�@���~�J��!�
/Y�p�P���u�d�Ė'q"�'~[���JK0B�IC 5&�Qk P�t/��h�O���?Q)O����O��FOd��b�2�μ� ɽ[�8�q�2O����O����O��<i�#�:z~�)\8;�,p
#k���1�e.и1y��W�h�Iiy��'`��'7����'w����% 6��{0L�:
'�5��F�>�7�a�	��'�B��"�~�,�<���:@�Q�D�N��k�i��Q�p�	۟����(���g�ܴu�ja���3��x5LA�4O�o��8��\yRENB]��'�?Y���*u�ۇ���!�"6A��!1$�)Z���?���?��HA�'Y���^4X���H��F�B4�ʔv���[�؛S��M��?���24R��])��uj�����p*f�Q�ߦi�����H��c�$�'%� ��	Nk��u!���;B,��DG�&j�� )�6-�O,���O�)^}�Y��[7�� U���g��H�R���M��o�<K>	��D�'ATiȳk^�!�h48���m��9�E�~�H�d�O��D�b�X�oZ�8�	����	ϟ��Xl.`�$�B��See�+� 7m-�$��6B�?�������I����s1�Ѫr�Y�k�5%��ߴ�?y
�:7ڛv�'��'��G�~
�'}�]�g�(�6�+�NӼY�V͂�O��ұ7O��D�O\�D�O���<�3�3��{��6;ִ�{�J3pl ӆ[���'G�\������ɍ^/�9�A���VE�@Ɏ�N�O�<���?9��?a����DǕ�\�̧�x��'�*sF��vc_���\lMy"�'��I͟����`���~Z#BN�ϲib�n
�"���yti����	����	ԟ��'=�(��~��8���C�c�N�H󇓩w^v��e�i=B]���	����S���I�����k�>$kf��  $�.P	2�m����I@yBT���맄?1��z�M40j�`�3�C�q�� 3ǈ�3`��ߟ�����D衯t��%����&7*tSB%Y�~}�v�UD|amEy�K4Y�6��O>��O��)T[}Zw��,q!̜0����	�x�b!
�4�?��}M�͓@A��~���}:�"�(v���-Q�Ak�Q�"������3�M��?����W��'Y�`�LJ���M���51��q�t�@E�2O~�O��?���7�� d��c�,9mb���h
z\y�i4��'v���.,7F���d�OH�ɨxCV�`0Ȗ�#P�́��B� x07��O˓wl|L�S���'��'BV4M̴8�8�+�*U�J�-Q�NrӤ�D�9
���'���Ɵ�'�Zc>,(8!ɉ�cA�U�>��O�#�3O>��Of�d�O���<q�n�1�����)ޛ_+d	Jh#�:a��_�ܖ''�X���	��	���[��Q�pɷ'�*=Q�a��4�	���I��$�'��m�s�i>��S)�wz���)�:M���a�<˓�?�*O>�d�O��$�F�S�K��@��ԃcB0j&�ˢC�"�oZݟp��͟��	Dy"�Q�맍?��W9]hP`am)�2�G�=��6�'?�	��|��ğ���q��IG?qRM_3`A� �B� .�f0�#M�즩�	ڟT�'�`�&��~���?��'u�����L��;⎔�QF��}��x2Z���	ϟ��	*p���ܟ��'%��|'�!���9R�`S�Z�b���_���T�5�M����?���bQ\��ݜ$!J	; �R�X�4-�3��'yR6�O��d]�U��ODʓϸO�}�0oqanY�խ?3���4��PA�i���'xb�Op�����\J��@
b�BB�EMH .�lZ2s�f�	ɟ �'K���$
$U�>�Pg,� K@�2@�6aN�l��@���
r�ͷ�ē�?y��~r��蔝����u��<�Sf���M�J>�[�<�O��'k��9D{"(��j�&(�X4�&D-�7��OT�%�y�ޟ,�	p�i�� �b?��]� 9n���>ѓ���<I+OT�$�O���<YfJP>%�D�f�$��0!��6��`3�x��'|��'®��v�с�(����ddM9�'����������'�4�;&/v>q�'L>V��Q�av
-�e� ��OΒOv���O��>O���d$$`���?	��Qsd�h}R�'��'��	Pھ��J|��]����G�ќ|��U�	,K����'��'���'J�s�'@�|µ��&	�۰B�,	�<m�ɟ��	Cy�@���"�d�\���B�tr,�+�7�� ����G�	ԟ��	�0�^Y�?�OT�W��>��&M�m�����4��&-]�eoھ��i�O��i�v~��Ǥ�v���]�dU�uiF���M����?Y�^���'�q�������)�ʉ&t��x!�i�B|Z�/t��$�OR�$��&���	5��qkT��+$���ƀ���ŒشZ��p���S�O���a�4X�mJ��d��ׯ���H7m�O����O2�)&��i�������_?9�cϖ~H�Ԃ�m�+W��4�e�L���'J͗]g�����Of�D�A�x���ςQTP�R �8?�@lڟ`��b����?�����c�Dާ��u(��&s)��FHB}�F���y�U����П���WybE+�� ��ő*:����řV▩�BA-��O�� �$�O�H6�6((���8_v�����̋.��l�����O��D�OJ�A嶭��5�ʰ�W( `��%�߹@D:,84�i��	��H�'��'�b�R#�yR)�;@Iw�_�{M��N������?���?��?�g�����'i�)35H��і�k���"E���'��	ğ���T�!�l�\�O��#�ꋫ����$�
(�LK��ѧ_�LXO�t ���c��/.0]�L�2+�l�8Ǡ��'r@,� ��H��$8�ƢE��r�׳P F��ׄAd�v�G�q�-דf�,�Tʕ�P�V|��@�O�xp��A�L�N�R��DI6ph\�)�F,B�B�f��ELA_(^�ȵ��s�J��gIʚr!6��TnՁ|V�tfJG�H�L|����%q���i��A�U�\��OǀFI���kޗPp��H0_���SVX��ea�ʫ8��`��*����v�׋A�\T��*�)^	X)���Ӌ�?Y��?a����{��D�<)�LU���	P�!�`c�I(Q�?�h��2�S�* 7O��p�� O{�YT��
�H��$!�g�ܱ���܄E�ʥ� ��J2q���!��|?a2�#~�
6��@��]+�R�?��O=�&����ɋYJm�!MO�x?���ə�6�C�	0s��!y%l - ���W�\����������'5!h� ��aw���Ek�'_�\�w�D<H8v�'���'g2 `��������';��Q'�ʐ]��i�(��+s�)��S�s�2��F/F&�@A�1�<��r��.�o��J2�, ��'c�>F!B��ҫ'R��a�I^4UZW���&�m3�<ʓ>����!|PFUQ$^�N���o[����	Y�'g�O�����&s���i,՜:��\�V"O�x��D�0he �*�쉄�ly�"�V����ITyR�Z/l���'�?)*Rd�Ԑ�/�t�	
ǆ��?���,�j�r���?��O�
@�!o& �=�$���"�ի�)v��5��(P��K6ǀ`��u)��t�'v���)ՠg��8B�"ˀW�����"d�֭�b��[&�, O�����W+B�Q��:TH�O
�ĺ<V�G�5ʜ��*� '/����v���=�V��%1>�sq"X�-�㠯�v<A��i�������w��aǪ�8kN��Q�'x�	�D��q!�O@���|���3�?�2Α�.����p�=L)N8��IZ��?�����d���@'�@��'�S]��m� 	�̐2��H�*���\���Iq~�x0q㒱a[j}r�g�c�����'�GⓂS��0(!���.��Щ �G�YX��'\t�I��u���v��d2�3� 0��`IV�0	
ңP n/Ę��d�O��=�*O��qȋ�w��p�х "����'�^6��æ!&��)AԠl!��M�T3z�l�9����O&�$HJ��S5��Od���O�����=���N$�|8f�E?�.�*S�V�`"@!�J�a����O�(2��c>e���ϲ���"&6���c�S�vap4�p��U鶵c�g����hG�	��� Su��۟IRK�'�jp�fM�-0Z��RD���'S�ɣ���4�Ģ=QRF`h�ׄ�[�\̙A�q�<��*P��5{��׌}�����q~�,��|�����$��h�x��e�2#BY�'K�#Ӡ�
4��:v\����OP��O0|���?)���t��+I�t0Re$�<|ND����)0�`��ˊ�b łt��/mP� C��F{ެ�Fy�)�n�tm��jWxO&q��h�7B�~��&�Z�	�6����@ ��z�
�gm/�y���#���(2���L����%������	$
$��S�B[�1�3'Jˎ5*B�/E��a6N$\6n��P,�/�b�hbߴ��p@AԶii��'\x�y&�;x��	s @E��,<	��'��&	��'o�	Q N/,�;S�ɐ���#�]�(�t�çG��<�b�(s�b�w)ފ�����dƧF�����L�4s��LV�RE7^��&�ӖS�8Ir"N�?;����Dـ_F��H��d�d��|��2 �ћ`j&$C������y�AC�0���p���"~*ia�S+�x2�|� ��� }PnDq�	,mb0P#w#2���JqTm�����@�D
���BFX�3C��w5T� F�� *��' �EE�S�2�!�$\q]H���GA�LqU^>5�(Q�mv�;�+^�C��I�A8}�Z�R=X��G�+4�ҝC�� 2q�A�E��n�4N߶1ol�C���#䣞�A�X�'��U;������O;>�JgmKF%Hs�-b��% �'�dq1#�A��zȺ����X�f%�Ó&󑞴�#ΎW��ASwD{�:M�dm��MK��?���-C �� ��?���?Y�Ӽ��M��3 �`��Ó�:Jx]��%��9� @�~_<����s6:�����`�I_�̓h��5%B78�%�e�*Ŧ��3BȇiSb�ʀ�/+y��(��'��(6/r�09W��U?�9cV�190��#.[j̓:4���)�3���!jꤙ�p� ����T%�!rg!�?=� �gR.���R��'7��	�HO�I-�N�m�Aø��,a��1/��-3���36���O����O8i�;�?������(Z��Qb���J�]���4����.=�����]�����#"j��q�O�4=X ����F�9���G���
��'�d(�bH@�;��z7��)@���x��M��?y�Q�r��'��A�H<r`*�n��i��e	gh^*(��WgQ�H�:t�<)��i��'x&��raa�4��OL�Ӵh��1�H�@ �ҘM0r��Q!�O��)f>�d�O"�S,��q	�@��]r�a�q����c���!JFe�$�	>L"��&L?O��y֯R��	�ᦕ0D��6��o NY�a��^3�AF�	{��x͇�?�I>�� B��ግ�,�l��CoR}�<Y�mB;:,�a ���@�J�}�!���Ȧ��� ���X�7h�48#BNn��/|A�p+۴�?9���I$=vd����/�hԻB�ݿ0?ܡ�r ˯^.���O��r0E�'0SK<�OY�ӷ$�����ӟ��9�Eòl�~�'h�� p��E��O��J���Q�e+�$��w�up�>��I��T�<�b�a 
�����4 �6����H�<�pi�2;��e�E�:"��d��̈D�$��R ��� %#P�C�l�7�<?^
n�֟��I���W���:nfm���X�	���ݼ[S�1s#Jź5`5��kM����<�`�Vx�<�f	k�^�ׂ"8/���%�� ����
�a@`���4��[�7�c��{��Oq��'p� �EEſh��AV	�c�ܣ
�'��������h�F�T+�y)�O��Dz�O��'vѓ0W�(�
�p@N�X�8XY1&�]�����'���'s$g�	������aW��;���%��s�/RKP�(ƕ�u��h��&Q�!7�'](��j� _C�Q� E�Xz��Q���	�A�A�ҭr�#,O��c��(��b���"e����'�O����O&�O��D�z<~̡C�ٗ��� �@�}$!��I�ě3E	wf�!��Eۓqn�O��lZ#�M�+O�<��E��-��ğ�R0�A;�H5��E�+��b�����I����	�H�	�$���8r�@� �&�bkX=�Fl9(���aL��J���ɠ Q�D ��X[��O��rC� �
A~	����>�� "4�'�.��?�X�p)��+��Y�Q@(y�1w�f������$&��G�� UJ����l���0'0�҂O
�m�yiI�νR�f%�!���\�[ش��Đ�E>r0n�����Is�t)�0�b���hZ8����$܀���S=���'�Tl ��&H���ѓ	��xh�H!����RU��]>�x�&�Cߠ�IA舧?D�	yF.}�f�
}Jpz��%��#3�V�
LԙPga�g����|ᮉ)�'�E�άѦ�pI�O\�Q$�'�1O�Lpr5�o`@��Y�ލ�"O��{Cf&�Z���Űsk�m�q�'�F#=��͊�P�z���%xP�n�b��6�'�"�'��Q�����2R�'I���y��o��#ӫ�[]��0�mje ����7�( �|�
�)Kݢ4��2U`݃���7�Jy��+�'B�����X�g�	(B�z�bN�+�TyY�!ˤS�(�<a�!���>�O6����t�(b�_�hP�"OT��f��AJ�d^OA;ҟ�Px���S�NY�e�� G�~�>�2w��Zʺ;e�ԝ6Tx@�I��P����,�Xw��'��	\
dNj	�#���A�c�X�����!�&|O�m���M�ZpC��
�%�dAP��n��ũ�+'khP��M�6�B(��͕��(ORi�e��*d	2H�P��X�*iyr��hR�#�O�-��F5�(Z��rі,Q�"OxH���-zdH���gź=� �!��Ŧ&���T�����O��9��% R��҆ǆ=��ui�k�OJ�d�i`���O��S�<H����К��iW�J%� sK2]�r���ϐ�1�ƨ� �[�'�������7i��a�8f,�J���"cst5�"_�z���q1R,Dџ����'�	U}>0�&�K�'���"!CTC䉵)�:�h�+<�cB���H}"C�I
�M� P�9��+��5pUQ�����?+O�	Y&� ަ]��П��O��1d�'PՉ��S�K�&���3)̨��'z��ڄh؍Bp��%e�m����r���'��I�q���[�3g�T�2�H�o��	H��c��X�:�ț9X�f=ʉ�d�&�\\S�	��z��۶-K����!?�.��V�)��ew��ۢ�Q�j��٦���-y�C�ɯd
�`ǅ��o�n��a��/3����$�D�'��M
D%��*ecE�C�Y�dQ�}Ӽ���O��D׼RenlJV��O ���OT�4��4`2�W�8E* 
	������d/��9:�t���
�m0HKc��s��G�H-4qO�0� �'��I�&�=D�f�X��� =<8ð=�D� 9��L>Y���kP����~P������~�<����R�L0�w-U]�&(R�A{~ %�S�O�~pS��N|�J�z��ĚPD����R ���' b�'�r�n���Iß�̧p��`c� ;t=��8���{>te[&�&��xB���W� ����T8��3�7+�� ��/���]���ͧ������>�J|Z0��dg��h"�[�k���a�'3>7���M�	fy2�'��Oh5i�cP���m1���u�	�4"O�]�Δ�j�pma���6 F�1O~���'p剐uzt]w���'�FP0&$���2M���0Њ�R��'R�&EC��'���ը:N ��B�l��'8���GG��8�D@�6�A#��x§�� �{R�5}��Y,(*KT'܌4���u��?�p<�D,ß�ߴ����'�BAJ惛+�p%aU�Y����t�S�O�r`�s��	1�0�0(D�4���'X�7�R�#�f�B��ׂ;���'bFs��Ķ<���
��'r�Y>�k�+某[߈D�
<R��,C��h�sZ���ɧ�|3t.îcj1:[v��{!+ñw�"l�O���zV@�,ݢd�D$_"@T~M�M�p�'E>s��;5��Q﮼��b�{�`@2�?�+D���@ڗ�� $�9@��5}��'�?Q��ir�6m�O�?���-�myv��FB$$~B R�3�I���	�.�V�`B�%	�΅�CA�19X�E{�O��#=!e�+nɡ�ÎT�n�K��@%Nכf�'���'V�c�B� U���'���'���$!�T��䎍6"�Z�Tނ`�1O�qi�'��t#�/ؒk(���S�V?TX�V�A� �d��e��O���EE�޸��Q<E�e�6v��Xe/!;r�Ae�|�!�?�}&�p�7�E�O�y��D��"���%�"D�(���J|��(����*-����4�!?���i>�&��R3�!5��a�M�h�p��<"�b��0��ݟ�������u��'��=��ꆃ�\S��sdӢ(������Y�n(zq�5� �e$�-�ϐ�-RM�Ņڌ�(O&q���
��j����͒��`�1`��jP���]1��$@���	;<Fx����wQQ�LY��u�����i�!W��� ���p�$"�Oj�c��F	t^Ԍ{���[	�x0�'	ɧ� ���Ǎ��9X����r�fL��d^զ�$����(I?�M����?A��J6G����̌�X(�U��`��?��A�x8���?Q�O�,0���M{z��wf�L|��"�?x*���Ǘ_3�<C@N�w�}"�F�E�'-*�����hU��j'�	 ����ל6&(hХ�-G츨y�ƃ�<ʤq�b�Y�'1�I��.�'L��&k�S�`����4)tYJ�'�xm�vK�-hN��H�B,.�^�3��D3��|�1�i�jQ�5�T�A;���v�֩C<4õ�|���$4M>6-�O��d�|���/�?Y��'Y�f�"��1v����(��?���ƩB�jAA�6ܳ�4_�0e�&���S���P_>���řs��	k�Ȗ�w��;W�1}�"�6K�z��VJ���V9X�H� [�a��NT;O��{ӿ��W�!@�U�HB*Lk|��G���I�V�����j�)�S�|���r�QO����!�դC��B䉄E�u��Z�z����/tU�PD{�ObD#=����{����Ņ0j�Z���_���'92�'z��� %B�r�'���yw�
�r�ȹ�NV�_s���� ��?7x )׸i�~]{����62���*擧}�$x#3O�����4?u��b@Z�+��aT��W"��P'ð2ؠ1��BEG,l�!�m�$�ʑVtƁ�;b��Ŗm5.� �K�$ς���|RMK��?�}&�trfN��8�a�UM�X|CB�1D�p���6���s����x�H���n��I��HO��$��S.&G�P�K1r	%�\"(gD4�f(���d�O@�D�O��;�?�����$`�@0��͗� �Fm�w	�q��!%L�8F�<�sëٮS����I��bT�@�ڭ� `�(N�t>ՙ@�J*�B�j%�Q�Bh��_F�'R�,_R2Y{�BA�Y&F1����3�����$��?��$��W{n!J3E��Qx�8�"c�O�<�p��>:�)�L�mD2$�G̓�O$t��A���5��ҟ�0�D�<_��mx1`GAո��Q+ ٟ��ɩ-Y~�	ٟ̧|�&ے��v�p� �� y�N�9K �5�fcA��>���	�:�����T�<E��+]X8����67=�q�������D�K�B�|B�B�
�� �Ď�kd�p3@@���yr���NzڱF�T>B��A�x�@~Ӗ���H�N��	���p� �k#��%N�<��'��[>���֟Q�-I��v1���S�I<���G+�ԟ$�	�h����DN�~��ū�>ћ.�^�'o ��H��liH1���D�2�`�OX +�N�Nl�|qp��)�MG���(���Ä:7���2����ɼunv�d����������\ເ��1�٨�g˕>O���"O��pT
�$�F����@�b��%�q�'^"=�"J�a���"�M=tQT�і�N5(����'I�'�Q:&��2�'��yh�1:��`�"[�(�c#
4D�*@s�g�Mnx,&藦0�rD3�iz[��B�'Y� �����d�4
ņW�T)`e�:V`ԈkA�At��Eh��Oo�����<� X�l�X�ˁ�;(�\L�P�	�'�TL��S�g�I$�fpJdH�&aP�i�f�[�u�tB�I!c�6��֣�:�Nm�!UΠ�]����v�ɑ,S��3U�4��ѧ�@�qq"�C�U�4����	ӟ4�^w�B�'g�)A9�~�G��2n �͹��˼u�\�`EO�z��.FW�h�� �&9�.��(O�]�!�d/F�"Ѹ%��p��`��O�;�ݰ5�'���$+o><��\�<N��A��v�!�� F�}��j�%%T��o�Sy1O���>��/��-?��'"�	5i�����۹x	�+�iB���'�V��'�'�":� �q�'�'2��R���'W���+�,��* �Ǔ}���?��aڭn�:]�F@A�K}X��ɓg8���tE�OV�%��+q!ԪRU��8��Ů+�L�Z�I.D��#�5ttı�Bٝ�͢��?��ܴf�L1c�)2�����#P�]���<�%��Z���ן��O�i��'X0��'�W��@"�f�9p��U�'���<k����!�9}9�T�$b�"m�S\���^��P2�I)CV���a ����c���aNl�*YBQ%ݍz0T�?�VH\0e�(hq0���BD��H/}� H��?�бi	�#}��'	@�r'�	}��p�Ѯ)!���'[
�6�N4U��l�r�?#}���
�.���$PF	Z�C����G#���N9�I��M����?��'�p�5���?���?������0N����ΝoS�9Fa51���!ǰ?@20ݴD��\��!Bl�g�	+KhX��a^�s����be�6x_���DO&G8����ir���y�g�ɒ��m��m2hϠE{2��%f��5�I>Ar����>�Op9CFG�z�r�"��B,q| "O��1�ڮQ:�	A�LY�Y¸YE��8���3� �]!g��0s�`���kR>;���/�
'�����)�OD�d�O�d�����?Y�OmBh��o@dɈ̓���#Q&���
#q��@�	��
Eڹ�C#�p�t�����R�'��@���l׾���
�"}bҐ�p�
.,�x��GhU��@�Bu`@0�pdc�l�P�'ͮ	!mʀp2°숎J�Ȗ�/�z�I���?QӧL�q��,��`A�8Pq��f�`��%�|z�(U�Q�]�7M�)Z��
rn/�I��M+L>�@/��+J���'�Ҏշ L��/PO��� ЪC���'L��)E�' r:��A��'E�'+��4��~w(uCU��rQ�Ǔq, M�$�Y�mr��SB^�M;Mߛ$� �s+ۍN��90�da8��#�N�OȒO�XhE�D�0�� SB�U�.�V�Z�"O40{�(�9WK��:���91�� p�O��lZ�3�l��E�O�u���҅+lL�`%��c� ���M���?�+�P��pe�ON �%�Un$ ê�0�0)�0��O<�䄓��Ap�,W5&���%�Y
`l��q�,]�2�'3�(�C����*W�Qs0���O����ܸƀ�`@�=@��a�`��m����?)K�#?�Rv�@i�"LB�d(}�l΁�?I��|��U���)�,.>�����yr��)���ī�/����b\�ў�s"=�
�	��Joi�l��G]2��f�'ab�'����2�'�b�yg̑�Oj�1���).���P$�./纩���Pc��4Kq�݊C�X��q�IQsƊ0�'�N1��l�%7���c$�2C����+;2�R�[�I�(�(+I_��OvJ���O��<!�aC��h��F�y�ˠ���'긩��S�g�ɕ6���*ԁ� fg�d��FQFp�C�ɠVv�aR�D�5�8���M�w�@�	ڟxя�4�b��#&X�~� bVN�M��qq1���"w��:% �Oz���Ol������?9�O�Tl ���>��`yd��Qz~�k`O�(���y`*��M3�CF{&X@���(O�U#�«t� �`��Q�By:�g)ca.�Zϖ ���Y�7
4Ce�B6F��Q��$<�B7FEHa��T�sL�x9Gc�#�r��'J��D�X�mp��Б��U��hF6o�a|ҟ|R/�y���צ��FL��#錩�'��7m2��ƛ=�p�oZ� �	0]�pɇ�$o">Q� ���Q����	ӟ�؅g���	�tQL��gX��#��8a����4Jav|���oH�<b!��{FZ��	�A	PŨ�lH�je ��&K��'�mJ���.�Xsgў����^�䝰�� �yy��h2��O������	[��m���"<���_�/'X��'*��'hɧ���j'�K���$��N�M�A�'�2Ep�����:@$C?!a�M�ǈ�����I4�M���RdR�f�'�B�'���D(DGB�AS]X�y�k����0��n�7���'���[�'�1O�3?Aq$úC��u��l/yp�m����P��-h���?�2��H.nv�1��ʁ J<��'}j���? �|��4I n@���#+X�+��yr'A$�y��z��x��ȟ+J�q�jƻ�0<���+0�&�1���i̶�Ӏ� �^�
۴�?i���?A�fY�]����?A��?�;�P��񁚕_���A� �.u�&�j��ٕ,v��%��_9�������d\8h3�l�<y�A*L��>F�L��v+U<�@�Q���pj�l��j�j�j5��ʄcej���ןp��Ƭ	��y7c�(k=p�����ed>��N�ei�j�<�.���>�$�Oh��^��p@B�^�#��y��Dà�-�S�ONp��#	ݑr���j`gJ�ZvB��?�Ѿi^�6M.�$����ɧ<����N�~�������a���[�j�p����?Y��?9�I��N�O��s>���BUz��	�-n�4T����~8B�I3u9����h�5QWf̘0��H`,93a6����蛱7�΁��F(t%�t{�#Y" ����X؟ ��b�	5��`�Ukߥ5�F �� =D��i���#�]�����-扭��'���+��z�����O����+�&XǭE�T���O��䕨]�L��On�S�������,͊Q��ܓ$yZ��*ٗ$�p�떁M��p��e[.�z�0��I�$�������=�2���'����!+��P�E�rf�1X�Ѷ�Ƕ,��=pf�	ev��d�y�	�
�Q�B��0.������S�R�BB�ɢ=�Z:�^1
��6����#<���4��nک��p8pk�l>X(F�Q���&�4��&�0�Mc���?�)�����Ovu���,��Z��F��-�O ��y}`�D$�|�'�9H���9%U���dŔ�_��:O�,j�O��{���&�>=��1G�����i�(p�C��.,"��Bg��_XL��B|�)��$5:$���A*R��ZUg�1t@,C�5/��:�%[�?<2TIĭ^ >�����	n�'~��CGn��'��8�@.Z=zL�I�m���D�OJ��Es���j��Ov���Oz�4�� �=z0��R	��"�B11��Ia��95��6-�G*.�a�f�9/c���|J4@ޤD��/"P��sI�4q��pc��Ӊ(Ű�q��?�\�jD�
�6�����,� }��(�0O���w愩M���%!b��-���O��BƼ��)��O���O�ʠHB8I�����mU�(<6�S�44�t���4:������D�#�`��ɠ�HO����Oʓyo|�h2��{��P��T��f�b�f�x���?��?"������O���Lpm�d.��h����������&��D��&0�)#gP��"L�s�	��(Z3"�	��@X���-,�l W��"8m����쁘(x{3�ĆE��(�0�I�T�h��Ǐ!O(�б�
>=4�8+A��O���$�0n��cw.;
���+��W�fxa|��|�K4O���v�ëi2��%#ӧ��'�h7m&��A����nZΟD��698M�@�G�n�Bc�����П��n���I�|:6��!}��CB�]ͦ���`J�'}�-�6%C,C/̽�r'�5�~yɁ!�
W:�|Gy�'�,q/ )�S� (ò��ǝ�������_02HX��2ǔ@yS��m|�F�Ξ",�'t����*-�'�6�u���p���(�ȩ�	�'Wd��eK�m�UQ�$3$�fҋ�$3��|BմiY�E��E�5Ԧ7dϓC<:��+�$�%_$�o�ן��I{����\T���.����,?A�`�I�R�b�'q��P/�J�*%�i}H!T�t�`�ݏ>��<T����䦔�x�ʴ���@�Pg�'�")�a��n����6�$��I�E���Q-�9N��֬l9� ć�5�����Y�a�uipM�I���%?%?5� �F��Ӥ��w��@���?��ڟ���g���(�B1r����K��D{�O�t#=i�O�]J��4-�$*�Lq�Ē7Q ���'���'�n���p�r�'^���y��k�E�Q�:�c#;E'�٥�i�<�pmՊB|\u�)擓u��c�=OQ��H�3Qr}�i��+m4y�Gi\�8�(P�<�F��2��Z�q��``O���y�Cлi� %9�A�*�D��M� Xf"��H�R�Oq�R�';�B�$R�DXc�0"��ѱ� 4��Аs�@$�q%��+V��� &N"���Ol�Ez�O�]��z���-�4�!����q���ݫjj&P{΃۟\�	ş��	��uW�'�B7�$��`ظ\������'��vT�ã�
�a�,L%Gd�8`�fإ�(O�s�Fh��aHN�L�Ar��;}��FZ&� ��7M
�)�T�0��(O�j5(�'Q:�"@k�s-��%�W���'�����F��T��l���#M�HEh㓴�G�R�*�mH).�ά��i�*
�8�<I�i�'>�`(l�>�$�O�!I	Qw6���eW -��iɑ��O���T�3Z`���OX�ӆf�u��cX�d7-��șЦ�ş�0i�H]� L�)H��_�,� ʓؠh��Q�!#N�0��kcHl�u�QL��CV ������;o��U��u^��8K>)�ҟ�3K<qЇ�ئ���,H��D ��s�<����B*��!@�2`Q�P�Tf�g�'�ў�ӈ�MVn�	J&��AXy�V�4QXNu�!�|r�A2EJL7�Oz�d�|"7�X��?AQ��'1D0(q&�o�����?�/&��(�[�;�PШڴ_PB������U\RgQ>c�d�8\����J,��`x��#}���j"�	X�R�^��a%��P���&B8{��Y���`�a�D�r�D��d>G��Y�>���埌�K>�zR�Wd,�q1*�Y�"dG XA�<A`Fۼ!I>�*Dd�;VR:�bfHG�hO�m�'�dݙ`�ЀO����g�%\��ov����O�y��aJ!E���d�O<��O�n�:e� t�P��y3����q���H<��	+fx(�|&�H��`����S��[ �$���K��'��� c#H�g�� M��qcAW�k�lI��B�����4Ej�I������'}B�'$�<�U�D>!b��b���ac�ʘ��xr��[��J�-B�hr�
�/v}p�Oz�Fz�U>͔'�.���%�/�|*S:.ih#����X��!�'���'�"{�%�	��̧H�t��ę�2fP�C�
���D9��CN<�!B�>C-���b���ZQ�pڵ*��Lx���@)�mX0L\cE^]��O�� ��{6��ǟl!��q�����ȹH�*�.1�Y�ȓ���@�d�I���v_�\/$��<��$>l�Zdn������M����������Y+���I���c�o̟�I�|�A���$��e�Ȝ_�����>r:�x� ?O�����'*NP{C-�2{P< ���H��x2m��?	�xbl�.8��AC�M�XR�E�	�y���4�t�����$+�$���͐��xk�0Xc���&U���KÂ<]��mcv"Of-�Dꊮ>��<�S+֤��i6"O� R|p%F6�q�RJM�|�$"O65�D�K*>��	̂B�\ ��"O�K��d��&[0��d�"O�X0l�*~AJB��3��XQ�"O�å�7�
� ���D���A"OVDZ&�R/�& X�O�4Z�!h�"O���W	�]0�%�p�n���"Or8Z�V8r���'�J�e���9d"O�7�	��Ā���\�{�b} E@8D���v�C���C�I�3SD^u���1D��s*ݒo�(Qɖ� �{ ���1D�d+�B %c���kFNC�#x�x�0�-D��PU�,m>@�4a��]�ē�K-D�(���K
}��թ�_�RF�o0D�x)�� �G��i�␴)c��)D��q!٣���۲-P���M�6�+D���	܍~��H��JK�(��)D�H�e�R�)�b�Q���1fH��A�&D��bS�R�\�tY*3m��M	����%D����kӑa�f���Ș� ��e{�/D�ܻg�6b_�ȳn�,9������,D�(�4��7�@� �Q�d�#4�/D�([��[�vY�\[�@>yM|����"D�D@Z9wQ����"W F]Z D�L�#�} 4����Գk�,qy�>D����E���5�� �t�Ε��=D�
p�K�Hx�e�ǂ�;%=�M���;D��l��",�t�Y��h0V�Rq�<��Eݶ Y��i� ;8`K�+�n�<�F�Kj��i*qi�%#H�0`��S�<)��A�v�౅��	U��*g$�P�<�Q�',𐥃"͙�nfn�B�K�<yuEF85  0����s�r��E�D�<A�EV|`kHh��x����|�<�B%J��h�d��,}^8��d�<A6T�9�|#���Dꞔ')@b�<YT��-+�z̰�Ӓ� !�L�Z$�)�;Oh��J�nU���y�!�輌HJ����TVf�
�G
�}h��c��<Q�"�~8����	D�f��@1!��#�.Qa�B3�$��cs.Pc�J#�3�$�(X���7n\�&�܈��O �!��	$zu�2�G�-2�)��X$���B�{B��<ч���i��'���!����lX�M
��
	�!�9P�ڱ���5_=��"�J�a�iu 5���с����Oڰ�~�q��|`�D
�eۄAH7Q�v���I*U��dـIHv7클OSԌ�f�R��k��3����5�i��-�JڳA#t�0v�{X��Y���+Gt�5�S��*��"�$n&��+Q����X�yသ�Fa�OAy��['uŎ�g��$@[z�s3"O���2�8zL
����E�"c����۩o�
��ì��yZ��?��b�����>�RDZ@�a��x"�.وY6$��Oh�'_��	36�K,��Kk4��<iR�J@�<�di@#�Ȑo1dO.u�cZ*���6�W��"E�	�OU����k��L�m�?vH��m��iP �έt�59�ºx ��ӕ��&E���H#�@�#N*���'�� z� �tPd��a=(�J����# 0�
ߴl>>-��C)9^���$i�	�>13*>.\��WJ��-9��J7s#!���#�����1��M���ӵye<�B����%n*�Iğ��!f���)�i��>mƸh�E�M�d�ۦ�+XZz	�Ys��!���RN��54+U��vDM�f��>S4�'l����A��i ����&%�9�����5-֌b����cb┢U�� �l��=)�V�)6�+5nL�t�M}�G]�u#ԥ�p @&F� B��1$2��7OM:KeP�hT+�p>aeÔE�@��)�:0ܔ8�����0M[���h���E�#��O�N�W����re��Sx��F`]�4!�D��~=Q�I�mK a���y�� �uq�����ږe 0pZ��ǜ�5�	��Eڌ�{(O κ��$�?�����1L�r9�we��Z�� �9���IY,,�J�%�$�h�>Y4"��\ˮH��"@�a�V�{&!��|&� ��5�$��ʇ�g����F?�=��a�k����%�2�Ĥ÷Z�H`re��Yn��b#P�+�:}��$f׶�Z���n���dZ#p�P�eB9Lbv��&�)�
*]!�`jAݮz_�!�H�~n�2��1S�]�v�d[��ܘ�h�uh��C\E+�',I��ʩ,�Z࣐�1nrpT)�����b�l4��V�$@E=�v,��@�:w���;Z�Y ��;���L��C����I�$|@�FFl<YY��͋_4���҃�0)�U���<a�.Z/>C�M�R%�?(�Vma��m�L<G�ڂ~�rq�$�W7>��c��e�'�px� ��EuĠ6AΏ.����Ӣ��9��I9�M2J�����Nm���է��#\԰"��y�����$��G�K�}����0�T�S�lC�		0��9$���4�'��sӸu��2OH�8�O��s�ɭB� xc��хu�0
�(I��x�!-r$�B�HH�$������
�y"O�4�7m�8\�����Ӧ18��ڟ�aB��D5��8�ሉ�MPZ����'�i� ��jˌ@ c��hN:�Kq��q�S�D�����ԀS=0��Oݞ�?I@�(��}�	J�6 "`��`�4`&%Lb�Z�A!S�($�d�����?I��m��r�0z����uH���Q@�'��9B��y9(;��7�gUrA��� �eY�D��}p�1sR-�q[���<��ԟ�I�<�_?�6e�V�1 -Ԍ-�&�1/	*Ӷ�k	�pr+D�kP�X �Մ=~D=��IA#c?B5�O��xD	��F~�'����^}"���HnJ���Q'4L���ds-�qk��:f����@U� r��Ʌ�+����Ӏ]	I�T%	$/ڻ����OJI ������}���%�����ĥUC``X��t��<���O��Pv���>�L]XI|�z�x�ei߳[Q�=� ���'}�����ɍhU ��$�)����$��4d�t;�Mˣ��I;4��1�GM:r纜���>��d��?˓`��a�n²9�∭;nt��P�A�t��eBY#
z(�BZ,A�a��Д;�8�j@(_�O� ����l�w�RHy�d�7$�y���1�H��2��J�J�D�8Q�Ӈ=�XI4�'*Z�jq�R�^Ĭ%��'�E`��� 6O �u��h� �1�!@$Fb��A}	�y�ӎ��D)*O�U���l����c��!J6>�	����.��M�xPlb>��'�`d�2F�4��9 v!�U�
���V&h�$M�4 l�.�R��@aX�X�%].l���4H@O\ܨ�D�7����"'P���D\d����'e��͝؟X�	(<|p4�7�&^z�u�#O�Z9ހ�Ɠ"���d%Խ
%���@dּ;*i��Y�L^�Ɍy�vT
�'���S�T�U��͚sa�~��⋡	(�����k�XU�JJ����Ԋ�0,�Y! ������iN,@�	������h��Up�'�a�$	<?��]>���Ө/#�4a�5�ԔHOh��2�ɶ�x,��¯~��0�F����f��\YuɯY[
�Xu�ʨfv: J��ѵא����'	PE#@MH���X{`nF9�B�sDBT������Gff7�P*q��'��^w�"�;�B��ˀ*��t$�hA��#`���o]Y�<!�F�<�A��|%bDD$�J��( �EZE$��V��80��lyJŦO��b��+� �QT�4�"�S��'��)(�:��Kq��7{B��J�-����8�g&��!�ގt_�E\�#��`�Ą��0<A��D�Bt�JU�'R�(�ҊJ���)�ւ*$�H�+PIW�ep�<y��9y��,�zԆ�*$!לG�ΐ����>����V�zh�U�
	�
�i�I��H�iᡗu��B��@}����6�y'�ŀ}N�=�� `�ȗD �ybG��!U�B*�?D�!��F���y�e�9$����6�0�>�#�?t��E�'B�0%��c�-H�	z�\K;G�����$}⮤����A(C�@̽u��9�4����P�P���T��Dۥ��6!< ��F�c��QFx��c����G
��9�/�O�dA��?:Gdp#��#�=p�Op&��oZ�A
 j(B2XM��b���Z�� "%#�!�O�`P���HR��|^�4���� I}0)i�m,d)�Ao�Y��j��z���6�4�F��GO���d��.\�E3�ɱ#�'F�l_d��&���,W	��tr"{�>�>gED�(�j	�Τ`���,:v�3��C���6��8BT�D~2��f���%U����(=�M!#ݫ-R���)a�<AfD�jy�'S8 '��A��1+B�J�b[��(O�`0'3��H�`�1B�L`qT���'��1XF�0�I�1v���4��O(�&*�p�� �ԥ�3N�\mZ�b�)"�9���p>��^�WiY��,�3B��\���9���{�N��M��8!P�;��S�s�y#���M������%x:�r%K?�O\�����U���N3�VAK����Aܠ�1�{RL� .���ɪ{M�Y%�B�dN��*�F䓢e�I>��a��\�Eh>U`f�ɨ<Ҵm!7�״t�T��� ݇JLl6��P��2'�&i�A�	]��y{t��(O%�d��Y���a㋗w���gW�� x5CŦ�M�	q����r��W�Z����0'��Zգ�
7�x��~�<�s�ж,�>�z�L�"h�h��
�y'lɶ哈H�)��I/R��09b�%���ց9�� !%�>��(E�NT�i����w�5`2�t��:CĜ�(��1h	�bf|D�0�Q+8
1c�n�Fۄh`&HC�t;h�0% 	Bb�h�E�<�q˄ p��D�'��Д$�nb�H� F�u�7�ּ7�,��kN�?�|�y��ė�wƲt�3�Ɯw,��c^�<���l1�"O�5�hY��N�]_�0Ф�oz�x1��i�˱�8F��I�>o�#<A���V���a��v] ]���(~�hqgJ<�� j���(LB�O�i��T��Xk��9vG�|Asˉ'���	��z��as��7t����$z�:�%�[eB��� ���1[B���|����5S�O�9�������y�<�V@<j���f�'2�P0h�+~n	XsKج�#T&�.C>��Ya&���lWH��������0�MX��MzqCȌT�PjɌw����O�f�����ǬR�ɣ��9yn\�+2�.�V��OZ�a$'���ܱ��Mg:Xh��xyr�¦J�6��d�Q*^`�K�!��O�	A	]�PY��MY��D����ơ`q��� 
ku�()����t���9(b�>ag�ґD�p��W"_�IA���6�,K��??��t��I�!u.h��e] � зb���^eZ�狴OV��H �O�O����� 
(%���F�a!. z$�C;�0=1�#؂tא<����4��S��Ǚq��i)b�P=E�����$u�1O���Y���sE[1+r�+�O�&�X�s~�y���̰t+����N�k����y�O�&����K�'^�����&�:��$�R�p~R(�@�W��n��Q� 9��	=�
E��+W�_ �I��*��T
,#<���4�GJ��%f.͐Ū�r!�qr�ӉA$�I�s���'!Ζ��0K�<���� M=�0��h`�(GO� T8�Լi�氳\��0>P��)�`�8p'� ~8UPG�7�(�p��g(*��uŋ⦽#�
�#7�'
ZPz)�"/��P�U�1Һ��c�Y+ܰ=�0NB�w��0h�3O�)#���)�����#�VY���f�BL����Aڽ/�R h���O�7����y�f�#x���`���qd��+R4��'����I�9�"~��x9%�,P�;eδ(֤�1�>`��kA�@ĻW�\��y��3�<[~aۦkV<�$�"���`U������:f�O��G��O���{*�bt�Y�8}���"On�M�-VD	I���Oo�����'�%�dI�pX�T�N�Z&���r�W=G��U�9D�xK�i��!���b�l�Q h+8D�$�ѤW�&�A��C�0���7g7D�0*R�X��i���FRڠ8ZЈ2D�TZeL�<�h|�UJؒ;X����i=D��#��l}HY����tӕ/&D�p��� �8��IM�Z�Jcj'D��!`L6e���0a��>%��d �-'D�X �;�����m^R���pN#D� �
#i��ـ��*U�r0#��?D���A���i��X6/�3~L�PA>D� Y4Ɵ�d<pLy����9~���$8D���L	�P���]1i�Թ�E1D�hq $��B�,�!s�ٸ+2�)� G1D�X�rLZ�R@ �󣗎=Xz(J�g)D�����]=@�����/�5���'D�(DET#%L�%�D�*@��/D�@����.Ζ�i'���p� D���רP"��X���`s�4�A D�tٔ��7B�M�FB/n�,b��=D��+�A]᮰J�ۇT�f��&D�@�VN�!1�B�	v�ڽ7���p�>D����e؂3�YZ̘	g�]8&�=D����cO�8fNܪ���xNX�U�:D�0i� ;� ��$*��Ga$D�LCa��+�^�c��fw&�2G� D�����q�eX���U�p�ǁ=D�8k��1+l��⣬����aF�6D�|Q�gS�y1x�;�"`T��])�y��L*G�b���A~ݙ����y2�
�H7�%8��p�^�����y��X�>%�8�b�R�jƘ�Z�&���y�%L>^ xHv�[/,��P��U�y
� D�jG�Y	p�ܩ)U@�-`�P�Q"O,4�vK�)U:,�E X�mO�m��"ON�R�m�>1�-�%N%;� h{"O�����T�R-�0��Q����"O��[��J=}Z����M$j����"O�
�DZb���;�"�?8��"O������w�8�[�⏪4F{�"O�,��eՠQy"m)����{(	�!"O*����F���$ 2�S��U@"OTdR����m ���y����"O����ٚaK��qnL�*�3"O�E� MS!F��!���h�&"O��Y3�C�q?��h���$�CR"O�ubd	حH͆ɛ��T��v=��"O��������@I��e)f�@��#"O������?����D�m���#�"On�s�6����Kf"O�j���*u�����$/�vT9�"O����%&���mEx��ɑ�"O�������cЍ��O��4�"O�	kqnV[�mC���:]�H��"O� �G�
�|2�
!0q�U"O ��Y�/,l��0J!-I���"O�9�k���5J+�؋�"O\9�o^@���#C���W"Oh�C�E�9L(�@c��H;⼔#"O�yа\��3�n�z�t$ T"OX��u�	�<���*æ"u���"OV-X��#X�qK�L�	�q8e"O��a�AN�t���C�+�
|�PW"O������~��u���>Y*��b"OF�If��q��D
��hA"@%"Op��Ť���<�ŨW�i�Ɉ"O��sĕ V���F�"~H8�P"O*̫�ڈ����ś�FX�A�"O��Qꖄ���04�ľl�nA��"O�a�6c!N%j�B�F��h�"Olk�\�Je�M�!�s��D�"O(���Ǳ����}���o-D�|��-ˁ2�(��]���t0q%*D���3-߇��i���(�\rh5D�L�vD܀>��`�������=D��0��O�.�,Hà5o@h��;D��B��$K�,���֌���#��:D�����f(}�ѧ�&~	B��2D�4��� l���m�:7�R�چ�3D�`��2N���K.J�*��fg2D�@�B�O�e*��^�{���Ej/D�8����p��S5l��y#���-D�p���N�-�6�k$�����!Ro*D��@(�� زl2���9<�NH3��(D��� .I�L�����L:c����@&D��Qa�]@���⁊7�|��*#D�t"��)�l3�a��O����?D�詠�T�&���#����[p2�5�3D�PjEh8�I��'S�8���+D��� ��S����'.���ص2�m?�d;�OZ8#2����$ض� 1��c "OPu�j ^�\H	G�@3�bmЇ"O�����G���q l�^��p���$�O��}��^b0�x�C;o��bAK���h��ȓC�$��6������G��"8J�'-,����������'8�D��'�aS�@�Oz��2 4���h�O���� f�ȣ��~�L�k! �(u�I*e"Ory	�DB:È��7��|i��`�"O|H��� �V����P�h>dIw�?�S�+3���X����,��&���U�`B�¦�#$
�;�XC���8~�B��Gm$D��Qw��-3r�P&N�!�8e��D'D����"
*��z4n�Wv�!1?��(4���AJ��蔢��X8&���0���� HE�5�����-
��7�d��,���ɴ@?C��Ex2�'#���go�F�^ [�DK!s.� 	�'�H���-�2DZ��n!��'��t �.�'^�\!��_�c`���
�'C� h�@�n�L���f�0^�*L�
�'&¼��C����e��Q;�
�'9iCe@����à�[��J1�	�'�^�!1"�LHTi���`�]��'W�q�Vd��T��1
iۏ(���'3��2+�a�L3A�{u�1Z	�'qP��(~�f���@�@�~�8�'��XJ��6kL��`e��$疀�'#$l��I�si���䁃�!f~u	�'�:|kQ�X)��%8�Ʌ�c��i�'���U���G�ΠH�o�_�I�y��IA�'OD�9#MG�^�l]zC�.@�~Ą�	k�'�*�(	E�����-�"��e��'�n��C )�Z�R5��$1-�����*�S�tp�di��ȕM������%�yBd�	q1�e��`�;��)`�Y%>ў"~�4Ѭ���ȅ��� +B��~�hl�ȓ&�J�i4��?x6$B�H�__����=�S�i|T  BB��I�%P�K��,�����2�	=T\�`K�?N�����@\ajB��5(u�(A'F/uz�e���c�HG{J|�1��)~���N'�J�*�`�<�Ɍ�J��%@1��R:>̩�
�����Y�����ͯ]���D��m����g+D����b� =�a�G�ͻ~`�`FkӺ����,p\XP*Ӱj�p8r>�hl��J��T��,!�̌�mĄ����I��B7�?�S��M�c��?]����/T�1pҩ��Lb�'�"=�O���@޻Z��H&�B�ċ
�'T�P3��>������4	�%QڴM����Љ�Y�H���m,���LS|��< T,%D�T �ޮ.�V��B��1ưԲ�ơ�0��I'wH,q��٬`H�R#
�w%HC�ɴR�!��#&��.\�E|�O����c����W�I>9�ͱ�B,�!�d�OrMZc�_�yr��v�ݸ7J@�"O�hk���8�=`_���]pǐx"�)�Ӭ��0�b�	j�:@��kZ2WDB�Ʉs��s�a�)!cX��FN�*���O�=�}��S�u���I��T;&
�G��q<Y�:f��{�	]$l�W�ҁ"�����]X�	1�D�6Y񂵂%GT	\v�1����?A$�!<x��R5bC혗��}�<AćW2r�v�3�@�m��h�u@�x��e�O��0���qL�yq���P��S�'!��`���Gݺ}R a�(ELXh�'*qI2)�;e=��P�/��9r���'���aAT����k�/�4;Zx��'E��k��.9���Ł7#�W���y��	'�<�J�l�7f�J�`B��y"
�?i}���@P&�YJR��y
� �X�GҰ`{�U'a�e;-�"OԘ�>s�i�0�;���:��x"�'tE
�"Y?Gt�$q'�� OLp���'�8r)V'"��
��X�{r�i��y����Q�R���,ҡm@�x�� ��y�#�=tmX��\%y44Q�I��/g��čY��(�5/��%ӑ�/ML�D,�S�O�^ܣP��"�$!�H4���	�'��0��=H�����t�P�y�)擱0�>!�/�9rF�]3��^x�pC�� B�>]��C�4{��]�dZ�f�*�9�S�O�lI9��SU_N1�a��D�nxz�"O�|���K/tf��� U�Y-�H�"OB��#�T%֢�y�ǋd$��8�"OM�q��E��px�.��2"X�C"OTH��q��a�@M\�$�N���Pj�'�O0b�$�r�
�6�b-�0a B�E���>D���)ϙ$8�<�iUKL�� �8D�h�G�A�&����Y�,�TKD*D��pql^�~����W
b�TѤ�"D��9E��0g"V:B��͛���(OL�}��&br�[��� �6�
"��p@�ͅȓA���1,�/_S4��3'S,H�D-F|���`�����K�2Gt�rAН �C�I�RҰ��j�$�2m��ިB�I>?rRU��0)g�!��l.�"=���T?���@�� ���<Y���`)D����DW�K^x4����U��jc�%D�����!��E�VJǻB� <9db!D��H�)~�y��ƽL�0*�>D��+���?X1!�h��1��k�e=D��J�k.��`ǯA$�$�J)D�h[���j��� �V�����kg��E{���X_*�e�	V����
�:9!�d����5����\����9C"!�]6�3�c�1:L����ޙ'!�dJ%}�+!��SYx�x�_�y0!��ܔ*��ˆL�9P�n@k�+�]!�dZ+F,6%�P�9(� �J���!�$Y�+�Z�ӁM Z�\��q���s�!�D�1:{���N�y��1�F�$g�!�@���d��AD�F��c�T?�!�DZ7��i5��u!@a�d��0�!�$��}�^�'(A�{���`b�@%�!���1G8����טy���e��S�!�ږ\���q�G��8"��J��I�!�D��s�9	 #�b��X���_�!��X�~h�0�k;
�=���Hxi!��b(�`A1��2¯[2@�!��C�k�f��t�T'����퇡%!�D+b����Y�83���LI��!���4if�R4YO v�Q�W��!�D>O�b䩷뗤& \i:1�֔&�!��������
�<�|ʤ�W�%!����e��Ӱ7������}!��1:S���C�X�U��1!FÂ4!� �a�<�)e٤8�J�"�^
(!��"XDƤX���AҔ%��,ɰax!���9���B��^ 2�L\3r+�p!�d��~��@[��X,1���cJ%U�!�$U#�@���F�(7ָ�tk��_�!��W�PSJ9C��o�p9��A�k�!��wX\A@	1�>0���_:Y�!�[*�2�Z@&I
7�ja'���Z�!�� ځ��K
6%R@�	��C%���At"O���U䗐O�n�@�ߵ^f���"O�l3G��TǺ�����H�q�a"O2��T�nؐ���$)V�+�"O��Hr�@�D,C+�>/<�A��"O.� 1H��o��)�2J�V,5��"Oʥ�4.	�9���*���&&ˠt�"O�4�܋J1�B��Иi� ��"O\M�tיL��PI��P��i "O
l�Co�P.zP���]�-u�dh2"Oj�q���ꔠ³^���g)��yg"?�pl��ӑ~vhpj�N���yꀮI����*ظr2�$ڧc0�y�EȞ<�Q���ΐi?ę��芾�yB�_<Z�a8�h�\�5�����yb�G,/�P���+؄&vN��M��y���$�V^
F4^<k��F>iH�B��4SIZ���ɓ)AR<1�$��@q�B䉂1.�#�Ҍde���h^1B�	�A l���ߊO��Q�h�.>�C䉙}DK��KOu�t��zC䉇[ۨA���1��$�`o+Y��B�	,,�mx���
�|�Ӣ�3Q�B�ɏ���S$��p5z��λX~C䉇y��0�sQ�9rR	�e��l����ڑ4��H�F��B�X�Ē-�!���ɀ!�R �t&����(b�!�dAbi2�S�Οw#�!ڲ`׉^�!�� ��y��!z��p [�!��  *�aD���q���� �i�!�dΏS�~HI�ŏ�#�t��w	�?Q^!�$� <p^��F�%
x01j�H�#a�!��=�P :�G���EE�S8\�!�� -
�hu�"]f�2�M�:�!򄔴U�fl#�b;(����f\��!��V�����E1*������	.!�$S�G	���!2WtE��0i�!��п`ڀ��f��)3/rT�"K��!��4)��lBs��*Z$����	V�g�!��*EP�x$�G"8� `	�1[!�d�;�x*�������[G�D�RN!�䑉%xt�8f���l����T�\�p/!� �,%"@P�!FbI�����s�!򤋇M~h�c�E�(掑S&�$S�!�όW�
IZ�����p��1�!�����Z�
.Wz�����Y�!����2 Ac��o<��g$ݒT!!���]�^��ϊ�:qv\��}�!�d�$Cs\�f��8�@ٙ�"\�b�!�dزKix���R���� M�Vt!�D��M�b�&զWk�q�ӯŋ}!�d��^����`��,�`��Λ�t�!��@3 n���AH(�nUr&(DV�!�A$X��� "Yj�Xi��)�1Sm!��0��I!�倜�Je��߳\E!�dG\/LL9Ԭ�2}��P���
Z!�dZ�b�(��՛O��a6$įc@!�$�(��)��\T��R#`�!�d�� ��䀃�� ,����O�!�!�Ė0u�806��w^"�s��ֿBh!�D�v��r��@�!%MN�!�D�0fi�1SM�+��hɐ�$l�!�D��m�4-
���M*���ƛ*�!�dT����W ��a�%^�tx!�� �����?�dy��*V!xNbp	q"O� �u���~���	�	K�ݱ�"O��
uǓ-� J2藅iG�S�"O�@��?W]85�ІŪX@���"OZ�ٗ�a`��A �ьA߈��d"O�В�'�$-�� ��䆤\�D�`�"O�r*M?K*TgDF�0�P!*c"O�5�6DƄ#0���?�nm{"O��z�e�#�ZE���Ωo�Ztҷ"O��J�Ă9s^"��Ў�6~h��"Oaq���7jf9��홿k4|��"Or4�a�%�X���+�KK��#"Oa�f�Q�҇H
6�M�P"O�a��F�$�$��	�m�"O��z0+X�A���Z�*^ �b�;�"Of�*'��V];C�
`�rI0"O���ጜiT��c�G<+_jA��"O`q(�kK�QEJ�xI�9ri�= "O&��E�/G�0��HS�= `t!�"O$3FaTO��}1�D� ����r"O��ʣ��|�����N��٦���"O&�����5Qq�E҆$� P2 ��C"OBE8��F�`�W�C �!G"O����G�1h&ר�z�a"Ozu�J]LB��3OFxI4"O ���M�+7&�`�cF	.J`2q"O��Y���#c�ء��d
a+r"O���Q�-E�N��2��-��Ԃ!"ORa��"ɝuq"$(�$nl�A� "O�APg&J�
�r��0�U�wP��z�"O~�k2CP�0�6�I�#Ϻ-��s3"OȰAq�V ���'N
It�"O8��"��@��ar"�\Q칪�"O��S��k���1p��N�[�"O�i�5LMT��4�;a�5��"O�Hf
�$�V�X1폻Rd!8"O@�`� �*8���bY�2CRu��"O8��-	�t��i1 ˡ2���"O �#ꔓ
h�0�@��AH����"O\�gA� {f  ��F-����"Oj��e#!tr���'M�XJH�"O�!ӇM�Ix��V�(Q����A"OX0�Y�J�f� !�J<4 ("O$�!�'�b<B��D'\�Q"O�!�`�7G%��pttm˳"ȎI�ݷGr���V_r@�"Of�3	��5�SF";&D��"OJ�Z��¶z�( ���-:�"O><�W��m1n���Ȟ��Hs�"Or�ju�*��a��V��Z��v"O�U��ox�3�F�r�^U��B�t�<���9*�J�QVOɏb��Ж�Ct�<����^��!a���5��s $�l�<A���VQNh�V�E0	�����Ve�<IBV�4JTT����$}4R �H�<c#G�v��GN�r��L��'�C�<�êg�>��`l�s؀��v�z�<!����[�����G[����n�<��,TK�eqT�_�&��E96�j�<�f�.����O|@YI��`�<�!�VXyȂ4Ο	���� �t�<yK:Et� 4��T�J� ���H�<��1\�H0*Q�}Z9xKH�<��U03Q�a�@�y��ѧ#�H�<� z��%-�+3	�ܘ��vgjAU"O� �C�9-��h!s	�=dm��ش"O*PU	�v����U$����$"O��:a@ʌ�Zh��/FFo&�iD"O�uBP��^IH���/��hV���"O���<Jz^�0��ĔPeF�{W"O����[�@{VQ�Ư�$1�W"O6�9�o$,N�pB�<zQj�"O~���V}X��fg߶B���Je"O�P2���,t��8p���9����"OA�6l�V%$$� �]眉U"O^,��̈́�%(!RA)�/�t�"O,|;��=Y���n�I�!p5"O�<�6��4��|뢮Ƭ)��G"O^)��^1�Z�Y3��J��as�"Oxˢ��-r�l�͒�-��R�"O椙!�3�L��s�ٰ$�T�"O�����&�Ҕ!W���A��ۓ"O���FТZJ!����b�:�"OЁ��	��u&��!����>}J5"OF9��JC-� ,�6�>(.aK�"O�S��[�,s�`�� ��h���qC"OR�2V�޺(��[��1�r�2�"O�e��e	����R7Ef��"O �yt�M(&<�!�l��CW��$"ON���2;dj�F��#-�F��T"O����I!B<�gc�FPH��"O��Ġ-i֌�*G��1==�( "OH�Ip��}��ԪEZ�$=Rr"O�ر�\�̙fmU�8�hX��"O Ix�D�\�9��nU�#l��Xe"O��hG�/4����>z81p"O�� bb��wq�-���a��/�yB�L$�� �_�D��l��jO�<�E [�I?V����9q����*�{�<�4l_0O��z0@!L3�$�7�t�<��B��u*n=v!V/����Jo�<섞�@hx�oI|�.|�m�<I��,�����h/,rdE!�p�<Y2,[rj}��D�?����c�m�<�u!�7b4��U�[�;�t�KWfi�<!1��f�<PK�둗d�4km�z�<�2�L	X�\b2��:R�0=#$"�y�<�&�4X�
��A
�ֆ�:F�Lv�<ц��v��Іe�9~�|�VIv�<1�(� ��(s!#��;<>̂�+�u�<��7k��! CFbʮ�AN�q�<�Gj�!��,�u ؘI��`@��c�<y�ꍑ>x��e� &>��M\�<�T,R�'�ʕr� ;.ΪA ���a�<����^$B�;�߰+��3��QZ�<��N�$�dȨ�C������g�V�<	R쏈���ѫY�<P��9�$Q{�<Ѣ�&��(��T	w�JKKt�<	%���[qƴP5k	1)�l��C��"r_DH�SEF�^I�ԅ�#��B䉃s-���'A�w�!�l�(bB�I|�vTd�
�P'@�w�D�y
:B�	(U�.���揻F��+A-NxB�I
j��yDH���꽐B����C� ��]�`*Q|����� 4;�C�	�-&�#���~H�[w���C�ə�����撖`�B��T�o�B��H� �*���	�m �;@�B�)� �|���C�l�H�y��A��в�"O4r�LB2?��i��Sd����"O��6��4�z)'ϛ�r@�0q�"O
�2K��@� %�nՈT<�*�*O�a�6�mu����� �
IQ
�'"5[�-��=�ȴ���U/	Հ���'��1���S�q��8�Pi��z٘!X�'.1��hFA���@/U�f(:��'4���S��1�ڈs#�7\�`My�'6n;#$�#)[}bg.��S���p�'��u��
�/)x �VeܵH� �`�'U
<QC�Z�pF�`��ӎ>��3�'�D� 3�����8�ph��4�
�'Ȏ<*�c�4-l���P.�5U���y�'�FtXR��;_����!\�V:��'F�P�K��[[D(h0`ЙI���'�2��G"-��kJ%G�rc
�'e�Z$e] V��`Kǣ�;�(lc	�'׬�8sQVO�9�!�P?e9
��'�D�ۓN.]rؓ�ɉ_� ��'��K��yP���	.���
�'*8�r @�~��I2A�r���	�'�:yPb�((Z5����:.`�s�'ERA;�eW�B��P̆�,��m
�'|���[N� H���K�/X\�!�'�KO,�E8 ��%<sb�p��U�<a���+̂��w�*M�P�'��z��0=p��=5Y���S�	�.P�׃Is�<鶌
�vDUj��^�d��J�k�<9ta�D�<�#A�r'�����j�<�*܆T�����ص3M��k���h�<�ĩaD�B�`�(q�)JT��f�<��@GI���vB�c\ �K�H�<9�F� f�"���/�4�DhkE�@�<�W�
�s����C�!�29�7��{�<IE !�Hht��1��`�c�Wp�<	�OWI�b�sq�A.<]��U��m�<AN��w$}sVZ�_ю���j�<���Γ7�d"���"v��K�fPj�<�1��H�б�E]��  #�gx���'4�R���(�Z`3��ۀqLl4��'P,��C˪Ȫ���i�cH\	�'�H�۠ R�+9����U_�E�
�'`�p�cn�1X��H�=Wt��
�'2�0���4�cǀ��	�l��	�'����Q쀍Y�!Cf�� �])	�'�����¯'dd��"%R� 	�'J~5�V�y�Ƙ�v��QJ%�	�'��Ёah�=�A�e�]�����'=vA���;Ry��E� @B���'oF�e�"���0��,ihl��'�|��Tb�3
p0a��#�P���'H�D8�AT�K���Pg��%�eZ�'l��f�I֤] 7�Z�?����'<��pC,W�G`Wc�>���'a�x�"�Uf>����>2�:�'YT� 3�� ��陗�L/X}i
�'�l�D�{),�ӑ�5,��[
�'|(�ʀ���yp�-1&Uh
�'�� "Fgy���n�+-�֡�'}jir�k���%h
U�*R����,6z�9`���E��oD)y�ȓ� ��r��${8PY�˨~���
P0bA"[�rڀ�0U�L 5L8���S�? H4p@���k	*D�qA<Oے|��"O"������I1�Ͱl�-8�"O��ڔ̌JV�5�a�R��pX�v"ODi�$�Ԃ3x��B�珃Y�
�P�"O2X��ׁ3��Ap��;$���qa"O@�gT�?'^��Uf��Y�n1�"O�\`&P�T��X���\T�U��"O�I�K�K5|8[7�UeJ��`�"O� b�	5Ǽ���N�|L�E"O�)�	V1=�z��I�&
}2"O ��툰$�%�F�y&���\0!�d�{�"��� 9CoT`p�X�_&!�$�1��%�1������an�74!��^��w�ɹY֊�G�ՆF!�L
U�0�n��	Ұ��P�=!�$�-��0ZbN��
��(� u�!�+z����'� m�1�ѠO�!�Ē1�h����������#��;�!�$G�Dx�IH��Ia$|��H�F�!�C$.��\����YpL��g�x�!�dYG"H8��6p�7�ǰ'�!�dP�:�b"��9-jt�ܕ�!�d��?�ؤ����Y)��˒�ؽ�!�d�V�|��bC�<mL���ݕ �!��!��a�%�^*`�� ��S!�Ā�R���s�?��y+����al!�䗝;�����'q�]��N��'�!�DG�x�5����i�� fh�O�!��Q�����1 G薃p�!��92?��g��@0���"�!�d�&	mڝk�#�'�� I6���!�5<j�8���]����O��!��6��ȕz����h&v!�$K�����D��i�1ʢ�B�Qj!�ĻbH	�$^l�
�+��	1P!��Pc1�8BM��;�ĭ8F�7Z<!�Df�ţJ��B!��T!���'(D�a��ҋ(�@9s���&!�V���q�S.|��Y��.�v؇�k��k�bCB��c���紩q�')����o��Q�ơ�
D,��
�'?~u�TI3K܀��X�{1a�'�d%a���P��H �.>���'�b��o��-B��#�M�|�.�x
�'��9RP�̑'��li�O-"��ՠ
�'�d����M��:��ֶgX�'m�Myf��5v�\�bg�k����'t��%U�q���f�՜_�X\�'� )��,9�%�fJX�OE:,��'��g
�;�$�[V͙�F�N{�'+̽PRf��p|SH�@�(���'���w��<9@�](��U@V ��	�'����0˔��0.F�>z���	�'�*,2b�Z:p��*�H�Aqf���'�v�h��3zᮍz'h]�-�0�	�''�PI7�[�l4)�E"�&+�ر��'���X��+Q[� 㔩K�R�.�I�'X,�q�@� d֦x����4I宰J
�'U\��!�	�R(�u�� �p�j �	�'���Тw���
5d #e�9Z	�':҈b#��z]�,a��,�����'�҉�t� �{+��q�DE�\��R�'��4cr�L>Z�4��w/>d�9K��x���OnN(��L{��ŉ��y
� @�@c5GP��R����b1"O�QA��M�l����B���d� "Oh""HG�#���fa'�Z<��"O��cN &���OĨ�Љ;6"O"i��O0%+"��`�*d4K�"O�e��F�?����.J�
���'�!��ͳn
����S<��
�-�(�!�ű"tq�%玚Y!0 ��GX�<�!�dE*�>@��\��\�	BƗ�1�!��h�|YB�䁶��S�� ?�!�$�)wdP�C�%�4e�������!�dW�o�����_�(�� �)���'`,J�&��2�{ ��6NX�J�"O�H�Ҍʇ��٤��9j4fq�0"O���n�4���R��V}��q"O<�r �cq(I��=pc�q�"Oz�jPF�8�d�!_� �"O��+�Z,q�����G�["�ˤ"OdAHԡR�v�N���LN0*�"OX�P��72^�q3�m�Hy��"O�C��Qu�m��AJ"e��`�2"O�q�b��+H���#ġO��4�S"O�� Fg�G�lQ�7�Y�w�@I��"O �@BF
�'o(Q˧&���!��"O��y#j�u�T��&��!�B-2�"O|L�#�� �4#���a~��Y"O4��[  1�LI �60q��r"O�@%FU�Hߢ�K���X��s"O,}R1�O31�aY���/N�X�"Oܸ���՛�xI�0n�LjJ�*"OHu�C ��As�((TL�gD���"O�-Z���iĆ���U1}L�!�U"OPQ�MX#i�"i�1��Z6>\��*O��3
). �s��N2|��`�	�'
�j�-�_���C�-_~��
�'�jx��$�����fT>"J<�	�'�JC��"о=Z�@�Lk�̓�'��ȩ������d@g �n�H<��'��$㇩ڨ#1��lIX=
�'�,y۳G�=�Re�'��<�Q�'�wa�h>�x� �X$D��'2��p��I�ܽp��� PO���
�'R��sHЫ"���U�b���k�<�P�Ht�|�1�.Q�yh�E�l�<i c
� �%c�臫Y�x=��Ao�<�S!N	� �V爦
�	�D�k�<�!�΄��]X� �uȽD�h�<i��� C"���~p�T��l�<9s�]����Ǔ"�P�%�n�<1�@T=6��$�B�{�Ti`@�q�<	A���9rf�T�"Y���m�<��<Y��ce	�iE0�(C@�d�<�v���$5�!ab�_4$y�e��A�k�<�7��;t| �QaOJ�1������d�<�t�L^��qK��KM1,Di��d�<QP�5Od�h�u!ٙF�`lB�#�`�<���F�.�����M-rꭢr�[q�<Q�jI&C�Z�%�-aM*��@��m�<����2�f�� '�-+ ����oCh�<�MQ�(���R���&�<x�Eg��<�2r7�l)��P�@	zd�Jy�<1�W�M�n]�3�V;̐����J�<��J��0T��c�)E�(��Pk�<�S�M�|�r��ůՏN(�J'g�O�<� ��+�)+7J�"��)r��F"O�q���
�rdq%�C�td�8і"O��:4S��A��D�y�����"O���4�W*^U��˴ᛧf�L�F"Or���C�hѢ�lS���"O���C x�����V�B(�`"O��S�@��6�:�i�r`}I�"Oz����g��u)���3��L�"O 8p��m�4��ՈB�"�D	��"O
�r4JL �(\��hߧv��:�"O�9�gC�J��}��оi��"O��遊�H�:!J��҈lf�a�"O��iU�J�y¤��D��m*���"O^`�se�;���(�͚4) D�"O 1�խ�X�`p�&B�N�n"'"O����J��]�׵0�X;"O����U�/�h��@�Q��ZW"O� C�F��	ֶ�+�hV� �Ƙp�"O0X�d׹S�r�S�$&g�4PYv"OhXڣ	Щ ����`�Z$�z�Q�"O Հ$�=���#!J�����"O���K�T��ya�>_.1c�"O�e�#��L`TI�G.x�ִ#"Oy[�H 	s���F�>l����A"O�]W��M��Ylǭk�.��"O^1�DXkҪ]��#�d�2�"OD����F�"A��a
��YsW"OʡQ�J�-�h�(E"�^ʸ�"O�8��O���XQ)p��1oЁ�"O�J�&ȯ���l�+T�t=��"O�m� �3W�X2 Kֻ1�0��v"OV=�t���`u�X�0�� �T"O�]�B%@�Z	d�K;vX���!"O@2�.O�e� $���<V@�M�"O�����Wnp���>&`MJ�"OnRB&V>q�$���H����2"OH�c���06�`���'GV�Q"Oa+��F���g/�5J;��"OVmI"śPB�)����sӮ)�E"O���2��F��H�B�ޏ2*�x��"O$�e�q�P͂㧜�v�(��"OP��GުR���jdg A��\�u"O�EK��g\[s��%S�e@v"O�T{����:�ϞT3H��"Ont:B)�>3�< ��cϫv��"O4�:�h�8�X9S4bfp�0��"O�I�%�(��*��SS�=�"O ��4l���D�7b�>M���"O�L �n�H�q8q��:n�S!"O�J�k�?^��;�/�5� $k�"O|�7D�	(x����-�kX�Ѻ�"OV`�d��Z���O�SX ;�"O�(��ٶQ�\�j'�H1rS���"OX	��V�1���E!��6F\9)"O�\���ȕ_̲e	!N%E,�� F"OJ��Gș�oS���4��<5 �K�"O�C�)�?x���B2dq"On|
 �M�B�SaLG� �`"O
�)a��Z��h"�Β%0��f�'"��f��!p���6��ؖ'E�m<=��$N�`�$��D��R�� Y��`�آr S��	E~m8A��I���n�9
����W�MI�H��v~�Q�M��c1��Eۼ�H؆�S�? �� %Q�-l�ɡE"=�b쫶"Om2ub�?�ZyS0�Y�8y�#6��d������A�V�zŋАO�� b%�5D��YW�,#�
�i鏨I�&�E� D��#�G�
ŉ��5i���&<D�d��a�eL�d�Fc�J��a1T�;D�tq�+φz�*#�wZ�\:E	7D�`��
Ӷ	/vd;#H*�s��^�<!��j��5�m��h�Y��E_�<��»M��;���
NЪ ��^�<y��ߗ��14�>a��Jc�So�<�4
�am��"���>L+=�#��g�<�B^�>�vu��b�w��� wO�H�<ђ�Nl��E�5�����H�πD�<��9T�X� g<Q}��h�.�}�<��m�(�TGŻ(�T�0�b�q�<���U�8�M	1�4/����m�<	TL�< 7��RB�0Pmƕ�g��h�<A1'�v�P%��+��8{����h�<I�OC7�v ���7��Ҷ��b�<!A�?#�i�ሌ���ӂA�e�<�cd��>Q��œ�jX~�q��g�<)���|*L��U���Ia�O�c�<�CG
x1
%"�_�wJ�aDǅY�<qeg�k�t!��-���"�CX�<�r�M�f��Q+�aQ�v�r"(k�<��#Y>F����e��a���
b�Tf�<YP��[�Ĥ�Ј��x�����F�<mO���LK@ゟU LBR(E�<����'�Y�,�+�0�HH�~�<I�K$Uk0�X���I9X-�w�V�<��ݍE&�@I�$�@2q��P�<y��O��\��H�A���3��I�<��$�=)bM���z^,{�K�F�<�We^�2��,R��[-5����'�z�<Y�*�\�|��L$R����Gt�<�gc��Y�(��G.�d�aE,\t�<ad��.@��"!� �t�c��y�<�@c��7X�`�ŝ{��R���\�<�ْ:^txZ�I<Z��-C$�!D�����\f$*�`0c۵h���Q�@?D�xD�;Z�@���ܒT� 8D�x豪A�fV�D)PI_�{�&��Ɔ1D���솛h���lB���q��.D���'o������9K&�� -D�8I4��qj�� ��>Y�8�*S -D�,�d	����e�sJ�R�]�A%&D���!X?9:��N�>4ڔ�P�0D��B@�
%T�E��N�*��,���0D����1&�iRI�m����b0T�Ђ�e�Aw�1�bƄ,y��L��"O�`y�E^�'����Eī5H���"OL@��h_�z+>1*�$)ry�"O|@�4�Do;�xFm�_qV��F"OR쬌)�Z�x�'�-k�l����e�<����Kd�Ȣ煛%[zI�f
�F�<��L 4W����P�Ne����%HZ�<�혓{���yR��,x�a�d�<'(�(���G��0Q��@���z�<)p�
<>0ש;.�HW�]�<�a2��u�V��?������`�<a�ʎ4vvm"���|��}���]�<���!>G��c@��*g���B�\�<��*���XȣCLͯ+�\�cɆ]�<� � �f�>H2D���#<xy��"OjI���G%3�<ŰS�P/��!D"ONx��!U�.�`c���L�;�"Oz����)c���a��ӻe��j�"O(pb�g3]<$���G
��S"Or�U�ŻE���#��^�9��"O�=�q��1-i��iuÈ� C�x�"Oh"��}��7&ր0\��RQNt�<����]&�1&��k��E��/Ur�<I&IJ�^�Vl6X�Q�~��n�g�<I����
��`c�iΏ$N(�-�c�<��#W�<*FqjЧ��f�5
���\�<)���D1��.��Ip�Z�<�3�_;Qz.���[!pN�0�v�U{�<	���rv�< e�Aw94��T�Ww�<Y5Я"�b���)���@�aZL�<��f�"U["�Y��i�H�Ą�#����d�����;����)ü؄�+#l% Kym���J1+¸��D��8�	^8[`"��EȐu$}�ȓ6n�\B��\ f�b�g	�~dD����b� .¼����4�M+�ȅȓ�
�x`B B|� ��o�=��ct9�	Gv;���?1�Z�ȓ"Z(��6.Y��%�p�0m�؜�ȓO���U'ڲSH�3R+P�n@��OY�(�E��8m��!P��.O��`��r@2�U�`�<���-�����TG�3�N$*���zGj�&�М��opX)hgE[2��h�E��d���|"�m)���V\4x����1#��ȓX�@�`��`Lt,���.&dB�I�I��嫶E�f���y5��)&OxB䉗:�������oF�P$�ӶXDB�Ƀ^F��B�
&h�tꦨ��v}*B�	!�h��D�}l��c�	�b�DB�1]DdQ��Y��4��kT�G�&B�	'U�LUH��C<pK�x����6��"O��BB�{�v-�SD��2���"O���qnT76�A�`h�%��9��"O�A#�<H<��s��K.�>� "O����╓(�*3���8r���a�"OȠQ'��p΄#0@+)Б�"O��)woK_BR�&�b�"�"Op�0&��
S�j�3ǂGa
���u"O�����yA�b��7���a"O��3��U
w����/�L@(B"OD�[1b,�#�cͻ�ڝbU"O �P	R͘MÔ)��/�,�"O�����$lɺ(ƍ4�b��"Oȼ0#���Yt&x�ѧ� &��2�"O��#!Þ69��8y�@��6��"O<d��L��n��<+�*_>蘰�"O,��b���6�hH3�H�>�.��"Oz�j1e�#u ��P�F�dZXZ5"Ou�A��j�/IĄXbφ'�y"��6��P�`�p�@���@K��y���='��dٕ'�n���S@�R�y�h�a��D�E
�k���և��y2���@Pl`a�b�j������y�
Y�\�(2M�9�X<Ô"���y�K�k��p�#-�R�`L@)�y�OS�w�� ��ѐ,������y�Ɲ��X ��[! �8�"'J�9�y
� |}iSg�}�F���X�&���
 "O��x��\�hlp��@\ V6�,H�"O��s�hY�|�R�9�/�
��C"O���Q�.'�`ѩ`oO�d
�,4"O<x�+N�P���N�EKj�P�"Ob0�l�rp�R��D2�D�"O������L�@-{#h�-D�q�"O<���:50��d�/V�\���"O���BB��5W����ڭ�1"O�K"�֨9������*t��""O|TS1�tbP�S�ar���"OuȖ��W��`K�d��SM2 ��"Ot��hBQQ��{��G4�5 �"O��6��+gXf�00��/J-�\�"OP葰K�<w��-9���D��"O�u�D`�a~�bQ�%Zh0�"OV�`.��(q���KF���x"O�-� ���%V���� R�C�p�"O�bC��+f��0�I�$%�x�B"O��Y�+߯:^$] U��7<���`"O���u�w*��nݔ�N�
�"OJ��Ӆ�P� �ڗ�b�i[�"ODe�C�'It��2fm�L�w"O��r�OV�@IC���)Q,K!"OZ]+���7yD��0'�-���"O�k��=$n�x�f B����r"O�����,G���3��IU��qa"Or�N��B�r��o��4Q�ѩ�"O�1�!��3A�84P�XM���H"O|�P�܆+RX�`_�B�X��"O��䇙���3T�-&��#�"O��jqE���Gj�+j	��ʵ"O�P9�LC�6&rx�T.=%�B�p@"O��*��B����ыo�X��"OTc�R�Ε6��:l��Ԋ"Ot��g��~�[u�P���Y	"OzuA�ؒd�JxY� �4:�j<�"OZ�9�/��G�:M�� �K�s�"O$5� _9Ѐ��O��d��a	�"O�) ��$Q�����o�c�2��"O|��ƍ��{��5�IH<$����!"ON�ǌ*�UR�i� T�H�{�"Of��b��2�L�#4С7xLT�D"O�@eV�>#��A�	�)jh�"e"O0Eb�؄Pj$ݱ�I^�FQ��C�"O�d�0Jě�����u�d�@����y�ԭY!8	2i#���4��	�'�:��a��C��Q���<hb%��'���1nY?s�]@��O<7����'����*	Lҡkq���6A�mR�'���9�A�I�<hD��+`n~���'^\�8B/�x�i`��Q���X�'X��YRǏ�%p�1�p��!C�<���'�|��ǍۜK��I0 �0I��ؐ�'�^Xu��2����cT��U��'�;#M�3�A��ɱ�>�2
�'̐aC�-��o�!Egyd�*�'�xcf�a���N��\�����'��e�6"�$�"�A5Pv���'��q�J�uw��ie�ȐI���z�'D�,Q��7���it-ՕX�$���'!P3�o�v؊�qt�يF�a��'z��"�H������?Нs�'�b�R"%%���sGX�3`hM�	��� ���Z��h�%S�g��q"O���咿5<�a��ꐟq[r��"O�\(2��v��5icj�YwFH��"OlQ�u�IX�\��׮ʎ0f��"O�y�֎�����CLǌTN��1�"O��$h����[�*�5ј���"O�� �ϫ\;X���l�v�x�G"OD�hP�,z��D*>4<`�"O�y�����@X�)۲<�v�:�"O�p�N�	g�� ���	?�\ �"O�E���B�LQF�ʗ	O������"O\hdC��d�2 Qg�KMd)A@"OF��G`_.�Xh�e�5}J"E "O�٫�'I�:�@t\�xEf�ZT"O�{W)XhG��XPL��i�����"O�X��۶(u��2�����x��"OT(`��.La8�S&�G�3'>uZf"O��d��X�L<�sN��f"O"���/��y�7[�{>�F"O���'��{���	ebʡO����"O>�2��qO���#�kBr��"O����E1�*�/|�.��f"ORlH�7�Z�k�F�r}X��"O��#����	bv�����>hBS"O�	���;l������o'���"O������TO�I�de���"O��t" ݬ8b��]9n��ٳ�"O�]q5��
#~&���#��K۔��"O���%�0*/��C��s�����"O�]�p.�KF�YT����1�"O�x�Vɂ�b tT�����Ār"O~�`�ʆs�sv@[;�rE�"O���С4 �R@P$5�8�W"O���#�/y�J����,q4��j�"O\���͕ d�(cE��.g0x8)�"O6��aI�(�u@7���9��z�"OD�3��ݸ�b�kT��<q	�'���"��:���U�#e:��Y	�'̆��U.�#�:�ЖJX�Vw洹�'���5�3ɨ�36.?|�*��'3^h;d���3 ����2?�"Ek�'�d��i��`��I��E�3���'���v�,X1PE"A+�ȬC�'�葸ҩ
I��y��TND���'w.��Sh�=}^�h��
]#�iY�'=0�/�����Fѱ7�f��5-�4�y���#.����*:/w��uD��y����aF&�*3njr����yrF��&�$劳fH(A�TPRL��y��N/N4�ê�$(1r�;�y)�-i: M��K�]��piу���y�&8�yEZ�4mP�BO��y�M�x|ltbi�P�P�wD)�y�$�.0�<F�ډZ4dP�@���y�M+MmؠK���<H��`N���y���&h��q��K�-}p-�K���yb�N�EFL���.��"�:�P��@��y�#׺S�C�i�,FV��g+��y�]Km�}��CFA}��ٖ�ۭ�y� ��<����c�3�2�Sc��y����4�x���$��yB�A��yb[�xP��3�/.�M��J� �yb���B��H*qbS�4��#��� �y��Fֆ4��+��v�6��Y�y
� �����ɰ;�� $2.�D�a"O^���O�\���Ba��1���Yw"OV8C ���&zP!�e3{��P"O2�3����)] ��OS��"On�5�O6��r��Y��5��"O6M�7NX�	-�I:�X�b�a�B"O ��cJ��/�}���ѧkt�dj�"O���eIC�@fNi���f^6�9�"O0	�6@�%n4�-��G�BU�)	#"O��iɛl$��W��8hB���"O�T���8_jqX�ċdSn|�4"Or��vb:�&�*�	��<?2���"OR)��k�2%�:���l�64��"OT��W#*x��Q�C���X�"O*� ��!<����V�|�Y�"O��CC��t�2����U�0e#"Oƈ["G��ZN� �s��" #�"O�����	W�Q�Fe� n�. +'"O��a���o�8����˵clȀID"O<a���5 ����b�؀�"O�Q��������gH�>\d�2"O����`�o�Tq���Euι��"O�Q���äU���^(ux,S�"O�`�\a+AjY�\��I�"OvC��}t}���ˇlRڄБ"O(�A�h��4�x�� kB�_�s�"OJyeo��.���
ɾ4����"OTh��ۀ��y� J�)v>|��"O"5Y��-�N����+@�D	"O�Q�ɋ����^�@�� w"O,��eU/ᖬ'`�H�"O�X0�DS�M��J�]�[N�MZ�"OhC�ȃqմq#�ڳlC D��"O���� ݹ)8�xs��Q;����"O���@���9���!u��@'F�r�"O�HJ��A �8����Z���"Ob4(�ŝ�F��9!���u�DE "O�yг�ys
T��Ā�I�|}p"O��X�J�+	VX�E��$�s"O�詤 ��M��xG'��d۸%�F"O�<�S	��#?�c�CX�\`�"On�h$JBJ+$��+[�C�X�%"O�\�U��uq.�:T�Vst�l p"O�4�S�XZ�DArP�4�TU#�"O�ѫQ�ɪ����b�"O|M���I89����gQ����a�"O��х�] 0+���f0q��s�"O���D.i���̔| �"O@<A�gƼp��Pp�A]�ز�C�"O��Y֬�!Wq�`� �R�*���"Or����Q!�L)�c� Ą�1u"O�lpfևP�Ј�oͭ:�,�p�"O�\`�ȇe�)2Q22���e"OTL�E��,]JH�Dς�fs��"0"O���Dм��i���A�6j����"O�P���H�:O�C����:^؜�U"O�,;�$�->@,���^5Iv(ʅ"OT�2�12;�����0-���7"O�Ԉ&�=i�p��A�~���"O�`ɣ+P
}jZ����N&b�Ų "O��%��^ �)��у+ 4�K�"O���B�+Y�N��E *�<Y@�"OXQ�⏈%#�x�2��:�H�"O!6�	j�t5 �)�Ԙ�"O� R����B	s�n�X��}�!�"Or<kd"�m�$��[�Js �J�"O �A�f�t�6�Q�5q��0"O\�� �-��/S�5id"O�]D�;Hi1� ��a0��"O0p1@����y����	�5#G"O ��smC�B:��ֈ��3դq"O0Ѣ'C� Cx��)K�_��"O|U��쀵o����e'&�CA"Od "@ '\�i� Z2aXjH2�"O��)0S�7����g��	*jP��"O
��3�$o��
���	Q�L`h�"O�HH�B��in�I$R2���r�"O��	��T+d>�����9X��	*�"O&��M��D��)�D��'��$� "O����"713�yxu`�!C4��"O�Qz�E�.;�`�A�.q`�"O�P*%��"Fp�-�w��Q�j$�"O���'�/4 b2�Bz�q�p"OLZr�R�J��H��jH���d"OD�Jŉ)q���L�T�8�"O���
-2�Xc�n��� �""OHH�� EKX��Lɻ`���2"O�0zעX>���˲�Цok����"O��	���4l*C(��%�t��"O �0״*��i�ĽpQ ᡡ"O �{�NI�QE�ŋ>S8��"O���t�܉�z *���<~�3"O�EXgK��RpɁ�'MJ=@��� �y�Q����w�ܻ:^��rL�y�nW��Mi��ъ>�T�c����yR�Q�)���ۣ��5!&@���y��%F���2�?d�Mࡪ���yBjL0yu��P�홲]x:�$�"�yRD��l�ZկFӾ�[�/��ybM�B0��fe^:' |H�ա�y�'G"��LٶF�*4��	�����Py"��<^`�Rb��]5�$8��Vn�<�`/"3��'J�d���l�<1%GM�HS�Xytn��t��aӬ�k�<��4!�&y�%��v�,�:S��e�<��A�k�8�pTe
d�E84Ta�<Au+S:{�Q��ώY��%�g��`�<��o��A�z�r�#�AGD�cbMM^�<Y�_�)�8�ؓ�ظ,��NVu�<`d�=Z��{uO1l�x%�m�L�<ٷO�-��%�Ah��3B�&��\�<�AL�%si�>%���f�N�<q��ƢCq������0V��c��E�<I���|D����I;6_b4��R}�<ѐDԾpdN<����L]R�BP�<��iM�\��%Q�f�"� H���K�<�@Ö;��E�t+4��m�5MR�<i ���� B����TʂQ�<����t����t�Ub���!��M�<v/s%X�@n�GbF}�U��39#!�$�&_mvi�(K�g���*�$y�!�ć�O5���RF�Y��Ir���B�!��S�Ao����n��C�
R
^�!�dLH Ѱ�g�6�%c�.ǡ�Pyb���	��0s��I�@�����yf&�,9� ��-�P�XQ.8�y���l����gتu���I#�yR��]�^@#G�)tw@�r$Ǩ�y
� �!�E��t� ���3(H�	�"O�lj󦒫4٠�Fߥ���k�"O2,)�h�97���Bf�I��=;�"O�a
8��R0�Jp���"OTM����4B��\����FFq�"O6,��)�'=������Q�N�p�"O���f�Q�7����f	�m��0D"O~i�#���AX��`�:D"D"OX�����ؓ���J>\�b"OR�(�G
����H�(\�}vu��"OHa�
ߗ0�ƨW(וv�(��"OؠJ�HG��Z,�C�'d�����"O�+��I�=�L!�R$�.�<�c�!4��C�G4)�|�b�Q�� ����>���.����d�zC��ӧ
Hx�܅ȓ�,��$��	�Dh�#�h�8\%�9���i�|�H+X�P�vE7�$�!�䓏f����pf�9Er�m2��� l�qO����сS�b\ PF��Ya����a�ўHF�$��`�;$��2����h�{�^C�	�^� x!H�q�µ�U�BX?<��d)�k�T	�*,��K%�8"�,���s?���1XM�mW�Kx]��'�y�<�2m�"�p���A�*��!+��l�'�a�� %t�R��ũ)'Б�@썂�y�fߣ<xb�R�?!טuP����?!a�)�<&�%Q���/4�n�)ҧūT��b�'-p���-�dI�!����IO�P[�'�Xh(7'�x�"�8Ɖ4U;6@k�'6H,"��U�G�B�&ƏL]\)��'�4)Ar-���zUXO	1л���yR`ڊoH��ALH�yN��$��6r�	P��H�8IY0'�T��m�Qb>;� +��'!�O t���5n���nKK����"O�	�� �7� ��%��vy4|Y�"O��_]�]��B�uΎtS�"OؽҒ�MX\�m�����Y{ӿi1O*�S�g�Dӓ^62Y��S�/(5s%@L#@�x�/ʓd	hE�vMH��d$�Z>u�)��O&J�Yn�(w=��JG)�z�'���O���%FP�$aХ�0n��0,�m�<y��݋{��Y F8th��aG`��0=��ƖvvLr�-����cd��Q�<1��^d� �Į�3R�m �P�<yȁ�J�6X�u�ǯdY��R$I�<Q��B��>m �٨���0���N!�J'Oz��K�V<���*AcؙPDazB�1}�3O�@�3vr�r�fS�?�D��W"O�$ �7Y>� �K  �4��"O���n���	�v�I(Xl*y��"O�ؐ�DZ�l?�X���XH|��/�B��)@�`����%�P2�ԧO����@�̼��;L[��;�͖'(��M�<����?�Ⰰ@ Q� lAS�F�ўH��S: h���B�.c-�!�gB[#�n#<a
ϓ6��`%�!](x{�4q:^����@�a�Ư'���Є�Kc�Rه�5=�b&��4�*����-���ȓY��)�k��k�
�`ǎr�$�ȓi�(H@�A���`K��_��ȓ+e|I�Q�g⨘�QhL�b_v͆ȓk�$qPP�e�XX�%�O�d�ȓPwx�Ea�5��(Ȃ���s�%��r�'��S�N�&I���W�r������� D`�%+���Xv���>+�"O���䬛��VH���9�$�`�"O��A@Ϋ{yj���t�rd�"O�Ɖ�F#|���"_�z�:|۰"O��(� �v�ݙ��� �i�`"O4��d�IVܾ[�΀�Mp iz%f-ғ�h��d�� $���&��l� 	�!�$C4n,yPF�P.Bnj�ǍW!S�2�8 �<��O�m��(XH���{��=U����"O�К��ɪ=��㗄��]E&�;D"O1Z6��W��Z�#�����Oj��tJ�|<���*��mqy��<D���m�*;߰)D�L����3C9D��1���s��-ʓLɊE �Ј%	8D��QQ��3F:�������$,kw:D�Xu��E�pl�ׁQ�x�a�:D��׮7��`�+�w�(��'$7D�ԡ�ա?ޑ�oZ�d�
@�t.4D� hÇE�|y�T����uw�u�F4D��90w,�*d�W�Ӣ�Ⴄ���=�r��"AL���ͻ$JZ%ڑ�i�B��Ʀ����F�@�5��"*�Yr�k�z٨���s�68*��Z�~ |�6��$��R��'Ց�����[�V$���%�ʢ"&.!IWm4D��R��Nf�5�U�C���  G�1?y��)§Sr<`��^�pd�dM�f$��fT�����5q��ȷ@�l��'_�D3�C�'���95�@�����0h�BJx�����yo4|�Giۇ��`��O�;�y���F�*��O P�2�Ar�M��yl�� V�v�ҿOۀ5AQ�W��yr
_G>�y#�]��+�J�y�LД<֜ ��H%� ��e��yb�]4��S��St�XP8P*�-�y�᙮*c^�A��Ԓw�2�2�C�y�IP��J ��Y�zm@ş��$<�S�Op��ʗ��
��1*��qOfH�	�'5<�b��8U��Wl�oJ�<��{��'"XMs��+g,���3jU9oڰ��	�'�p��D��B�kF	 T&4D�	�'��\�#hB�7
r���ȟ�[zr�'Ӡx�&"���VU�b��T$	��'���K#@�paP�H��7�Lx���hO?�y2n~"Ҵ�@�E�p��DAUf�<!eD$hl��$lB�2���� )�J�<�e�(�T�
�J�70�����_E�<1���|(^��Ӧ����(y2�{�<y��8j��CJ&
J ����u�<A���&D��L���KLqp���E�<٤�B�8�K�+,�*�cg�B)C\,B�	&?8�T�Ʌ=(0���\WLB�	�BSjj�Iuo�����_K�C�I�X���QC�)F��y� �'db�C��D�� ���#NM�ݰ@�<lܚC�	 3�:��ԃJV��°
��AOpC�ɋh��k��֩������qVC�I!%��6n�<j�z��
��-�LC䉽rj���6	�ep�"�M*uhC�ɪ~�P!��n��X�ə&^�B��<n ^����U��h��B�
zC�Bp���5�H�1��1����Jx�C�	�Va��9ԫY�`W0�4%X��B��9+���+�Y�E��cM58�C�I>��I�&�dC�4"�ȧs$�C�)� �pK�����%Ŀ�,��"OLK����)�c�P%��U"O���c&D6Ě0S�b\��4�A"O�x��
X�&>ZlK�D�N�T9��"Ov��Qn��n�T,�EF{pM�c"O���Z$Rr�����[�OͶ| �"OD�Th/j{HBb�@�HЂ�"O���#��k�|��-@"F� �"O�$j&/Ƹ9���R�l�S�ph�"O��:�W��܀a	_|2�Q�"O��0�쏷	��5��g�2C�5;�'Nؘ��҃<���� O��! �'$���A�G	WB��@��Α �#�'mt=rV��$t��M`I[��� ��'x@�P�1S12|hw�L$e��H�'�j�P��8��P˪Z��0�
�'��"���<In�����|�2m��'��J�)ď],�u-2m��2
�'��,����I/(�2o[g1��z	�'li��,�8[v�(�-hp*ų�'��!���^�`n|ᅒ�4e� �'v���)b� �[�틘D3�d8
�'q��Cr�=D-#e�=C�X��
�'�fp��p%�A(�'�4��(�'-��٦lP�I�*�1�ꃃ ����'�j�Q�>^�d�JD��|�<A��'�:��$@��ƴ�T�#<�2�c�X�;�,�����<�� Ӌ��I�1O��ՠA=!/�d�'����"O.!��X��Z� Db8<��Ш�"O������&����β	�HyQ"OI�ˉ�)>�j� ڔ�biڂ"Ob`36�ޘr�<4����И퐆"O�Y�e(�¹*�ac���w"O���EjV��@L=?�`���"O���S=��QŃ7|RЌb"O��N=E�����8?4��@"O�`R*ޙd,@eDPL�m!�"Oڽk� �!1������Թi���"O�%В�Z>)]��rBÂ�	���xU"O������)8�j(QI3���"Op�d�B�`��z]Qό�p��z�<!!�X��b�J��D�r˺�(u XR�<9&BK9%N�E� O�H�\X���t�<�e��#6N�$BϹ02�	0R�AH�<�Vù,E�t E�eP���VJ�<YwHӤg�L��c����",�F�<)�٦�,��4�4*K�X�c�@�<���������ǀ3oJ��Qf�LV�<��ޜV��E��'ܖ)���C�o�<磍��\i�b�&}
���Xj�<Q��̹r�X)��fB"��D���B�<a���5H:4����d`vb�<��b��C-��r r������Y�<I��ÃC"�`4�XF6R�9�(+T�8 ���c7��#��+G5�P��5D� �!�G��a��-O4`� ��4D�4�� �% ���cU�J���(bԮ$D���F@� uqb��"�x�K��#D�b�R0}�4H� g��L`�*OP�A��B� ���,<ҡ�d"O�p����Y��lʕ�I�m�|��$"O��:�Ȉ7K-�!�ѧ#���"Ot���i�*�	�"�S,�f�3Q"O��yc�je�a,W��<X��"O� �)��D�S�����I5��F"OF�:ׁϩ`�yJ���Pβ%�B"O"�;$Ŋ�"�b�p��\���"Ojm��J�h4�0�g��j���"O8�����+I�4і��'��|��"O^����-�4Ijp�.�0���"O�2C�K�$V�I2�C�;���y5"O�Հ1�_)S�ԅ"�#+q2`�"Of�I1�-wD��#�b����m4"Of�x4�G�!u@�j�b �R|�V"O0lc��׸ _@u�&A�'.ĕ�0"O�;� I$e����1��R�"O"��F@�+Q���d��(	�9�"O���P�R"Bf�9�n�"~(�"Oz�0��C2����mŽnȢ �"O���A���	 �
��F�<պ�"O���H�?7�,Z�(�$t��A!a"O:�Ӫ�:�~A�E)��4�&q+�"Of��&�ՙmH��z��c��تt"Oz(� �%xw^a������C"O��Kw�Ԟ)�r�X�b�*Ӌ��y2K��X_ |ɂ�Q��0�G���y�	a:��"Z��$C�n�;Ht�ȓ&�֤����oϸxĮ�[R���ȓp�лLϘQS�.S"bڮE�ȓf�Y��I�%��	�f��P*<���wY�hTn��-�UPB��I��T�ȓ%r�ȷ�F$LP�pa �
U0�ȓ���Ҁ�nh�l�!�� v����$ђ��/A�q�dx㏊4��m��zɴ}� ς�:����$��#LN<�ȓRt��z¡ǂ WF�I3&�Sa@ ��P�d+����A�&\���G¸�#�T)V�Z���@�)�6��ȓ&�H %@1�z���R����ȓOi0��-X��|���<����7��`SB�j0q�R3\�N0��<�a�B 2�P^�-�:|�ȓe����3�J�z�AӾi`���Iфp�q��(Kv�c	�?k�l�ȓ=F�9�3�
�P�
%����ZZ̈́�3�й�ECɦL  ѩ���:mƠ���@d���"'Ι?S�<ZFٮ0��ȓP�=[���9Z=�AŅ�^���ȓf���QD�7O��=Z����P&��ȓI�\8C��i��!7�ۋsby���za^b��١eA�v����b붩B�~LY4���@�RU�ȓ9l��xql��B��y���O%jx�`����Ȳ?�
��钻a�Ԝ��!�J�<�AmJQ����;$��ᢓ�RC�<9Uc����BU�H�����Ht�<��#�$2��;�ީru�i2�i s�<�  �#o��= �Π0%v�����j�<�rhӥxמPp��	'i�9k��e�<)2́�yTZ�bkF�6��0�6`�\�<A�	ϊr8�� /ڼz��%QSǐ_�<��@��uִX$.]�p[�TP���B�<i$ŷq=v�K�)��|W�X(��r�<�$�
]
�H8��7K*��r�L�i�<iE�κ ��=A�L�.B�FL*Q�a�<IQ푊o$�%إ�P
⏎p�<9a���$(�}׉ƧQu��	�Kf�'�L�Db�
b�q�����S���IQ��à.���N�&�y
� nI� K<U�D" �~S�|��ibE��'��J�
К�/�>E��4H��[FWW� �*?ZN\�ȓ-l�'N�7�d��������ɚ'�X��ɇ�V�O����O��IA�q40���Nė(�P����' �T����,�̸��'e��䂃�ۏue�x��eW�w~�Xq�-.�O´I'�7C.L�2J�=.��P"��E�L��![ �����+TDJ���~: IW�b|��OT�63x�0"q�<�P$	
�{�Fӷ1%(P��9��`" �>rc"QC#�� ��G��'�T�qÝ�E�f�z���K*)�'�b��d�! ����"�B��<QM� J��ɃN!�H�A���F}R��Y*P��-�Gh5� Ū��=aDA��
�J�B�)�^�t�(12.̉�cEu��@00�5N�z3��@���> ��h�7ge���?�l̘z���z��Όjd����!n��S*9N�!S�N�>y�aX7�R�:rC�ɦk�l�cq� *2@�	��G�g�>}�v�<
�4���%nCFʓf�O���R��*Г@!ƹ�To�Kt!��zry	g�S�;*���񧙐1��4@��s>,��B�>p�=y��O{t�=1c�74d8��#�nH��4�P����A�N��,iՃ�!'��B�b��B�d�i� �g$8a��Ϭ -ʙ34�'�Ј�ܷ]ܥ� �&�H�+�r�'p5c��M�d��A��!�7hQ�� r��bDT�f$�kC��p�Ȇ!]e�<9��T"L: ��W/�<Xq$��s{L�	�DC MTjQ�"j M�t��4���Q�A�H+M
�]b7�_�wE�y�!�:D���R]K(���/�Z�j�\b�I���$J�س�hD�A8�H�VQ?�Dy��ȗaLҕ�%LD�`:0IQ�L���>YJ�
-��@aV��	`�QJ�n�4:��0[q���!�>����Y'g�E��	;�"u;�.U����BY��X��(p�a��,�)5*P�!5��2R��2fv�����5��,�d�r�*B�	�Y�E����D��i����-*l��Z�Yɂ� ��\�����R���[ ?Qö���	apj�8mP~��G��<��@Gj"9ka�8N*܁�.6�@�f���t��0D��Bݪ� �Fk 1KnWz?q�v�=���6i���S-:Hо1�%� �O�!�U��O"�����p������T
�zQi�E�2z�xr��O*;HBU��˗՟ ��&u�����d4批4�Z,*c�$�.���I9�t�O,���C	�9�p�{�� 4�B�8�6�X�È�7�R���a3c�K�8]"2I��*\�=fi��wh���eBdx�Hh�ϊt1کh]���1V��-ly"<�GŇ;�B��4��djt��G�"|Qz���΅+Jm��&�,n}*(�'E=4pc�W�LZ�᷄�bVRل�	*y&�+'$�;I)�z$�G%&�v,@ N�vKN��4BA�A�bdrM���K��8O-
�JD�Ƨ#�l`��9pGX�Q�M�#U�hEa���)E&(�FL?��m�R!�ue����h��~f�I��I��^8Z�a�0�4�`�����Gm⦉�Æ�	�������8k�18H�ఖ�M="�԰���N�m�(�qE�<A�n�8٦��4�D;�5S#�	�3㰌��Z�L6Xh�PC��2/�� ���E�TIHt�JLVT��O!(��8���B˼�����u8�Ca�X�(�AF�Ψ�������3�E�qH��`.�:JKh��!;�.���:�qB���Dوw�m�r-�2��}�[�](���.'�}�
�'�e��MM�R�ک��aX�Y��u��MS�б�"K�eT�)E/�N}��]3��� N(y�ft;FC*V�
���@�$;j�RB���٨��$�,6�	cFё?�f$�ŨF�KV��D:�t C��&C|��@�\#�MC� E`䍊4c�-td�[��rL�(�&�*K5�ԦOj��g��.,0Ǟ,0���V�|�0X�<�~��FF�30X�+F��-��/�kcfuQ�D=g�n�9�OJ��C-Q!`r(YHsK�e2s`�U��d��H�xB�XD���Hѯg� �j`�U�|?���!
��R6�i訪ЯG41�8��#��\ʄ9��@�	�rLsK\�޸����>�@P�r�P�/�ȥ	�/�½Q1�� }Px��@̖��/�)OS��S�zq$ѡ�+{�4���E;y^p�瀒̒��G��LT��/F���b�UgG�{s�B�O�T���d�ts�dYw)X��j��7홆U��q���w+�X�4�1\�](��ڥ|���	�bL��U��W��i��*�t-�@�L��A�����@�N�E["�<y��^�-B������F��x�B	�joH4�WjB�g��p��J��uV�"�O��a���h��I��0� � ��W���2F�8O<��I�>�1�i�'R��l����2
����M�:�R��K4&�IЄ'FN�����h�@R�h;���O xq�ڈG1�,��L180䋡`�W��,��EUq����b�ީAP`��O��~�8���*��Yb����O��H�TI�'�ꜚ��[��1���%k���ɞfj�d���j��T#�WNQ���0��#��`eB�}�M�@@K}��H��� �%w�[��`$��D-����d ��{��t��?|��RS���`��)��!�y��Y(7��(&���0=a  �X�t�u�H���<Nh���	&x��` ��� Z�酬VZ��k��є�c"O����P��lI�ĕ�\d��"O�����VR�je#6��>P�f��"O���-�G�D��C6%M���"O��J�Cͦn(�Б!�_P(j�{�"Ot`���T�y�OH-f��Y�#"O*hk������겭Ƈ��a� "O���b��Ⱦ�{�팄g��PPG"OP�gC-a\:q���ڦa>���"O =�P!��2?�D!�G&;��"O����L_��:7�ӹ(�P"O9�!a
�^T�$�2L���"O�1/ژ�ˑ�0��e�vE���yr�J�o�Qð���x�`$�F�ȡ�yBCK8����*� �@Xa� �y�@��I�¥B��I�(Du���R��y��(3��i�W��d��ڣ��y�ƄH�\`���E6$��<s�*��yң�!2`訐����ju{��	��yR��=qGF	��A��i�r͒<�y��K�C�q��P%
�`� #hY��yK0b��ze�u�h�2���yRMҦ'�z�����v�Ԁ�"e��yrf�<�t4�we6��qBKL?�y�)ƽ<���r��ʗm�*���$�y"`�3!2�pr��{�� ���y��5N�4Sf���|�����y�����+EIM�������y�+AM�l1���O�\�	v���y�솊D�̜��K51Cx[��9�y�^l@�r�EAbl���D��y�S�����I"0oD%�PG��y��\;kJ�9���,+�EQw-֗�yb��F-x3%�>�˦f�y�A�;/D�x���?@�k�b�1�y�g7�`FAɞ]P�ݑ�E��y�/2t�N���˕PB^�zo��y2%��"z�x��������K��yBˉ5�t�	#lR�Q_r��"K�:�yr�?6;`��N��iJG*P�yBcʅ	1�����D[�!p�,�y")��P��0A��-D�4`��I��y�⓿v	�����/��x����y3�����˩#7`��u"�y҇V�Y.b]C�mZ�������y�(ώr،��*�]M�)�yb&�f�V\#��˼_�"u� J�y�E>�(���.�;8����b���y����}���P�؄LV�%(�]��y2k@._�Dm�E雷s�a(F)�y���?����@�nl`=��nP�y�l�83~&y��胊\Lx��p�Õ�y��SM�����O� ���wB��y�D�T6�)��N�	�v@���1�y"�)ʪ}�bZ�~3����9�yb��-�M	!�.�I���G`!�D�.\7�Ɋ��F	6;E��D�T
!�$Oi$�)�#e��pB*R@S�;,!�ă��N	�#�\�R"����I�"!�$̒d���a/��$��D��c!�d[�oX���ĵ:T� q�d�9!�D�6
\L�"(^��RAR3�_>c!��V"�(��bK9aݦ99��ɭ!�d�:J4�)��+��h�漡�,�n!�� Љˑ�I�ۖ������b��BP"O�`Q P�Z�l�1H�%JP��"O�|Z�O�;�
�sh�6;�.� #"O�Ő�ы`�Xc���vE�""O�4�a�Y'���d���N�xA"Oj�vnМ3��� p�X�;H9�"O��Ů�0O��q1�;%��ɧ"O�mj�Η+���rW�اeΥ�"O�xȄ&e����e7;�x�2�"O�di�������ŃȢu�h��"Om���W�hϺ z�eY���q"O���P�;���c�D�`=j�*D"O�����ь�L��eM� ��"OTx�r��_i��K�v[��B"O`���D
�7�R�⊞� 3|y��"O<�;�.V/]e
ch�1V
�"O�,���R�F�q�׉6���"O�)�4��>������"��dq�"O�@Y���(L�%�$ߜ}��l�C"Oy4l&��GDE9�xY`�"Ob]2�8<}�!a0�b�"O(��a�P��T���
+s�\���"O�U[��&���T�$.�|D�"O��1!o�X�~�����I�t�	U"OB�`��ο^�P�ԩ�5nk�Թ"O$Ca��M2
����0P�x%"O"x!��	����� ��O ��2"O��Q��S�ѫ��E�-.LX�"O��Yw�,3W��bc�M�\�"Or��G�߯cѲH�ԯ 򅂐>�!�$֩-(�[ ��}u�	p 	D�!�$ύMF.��s+]e.i�舊�!�$F-�l�(����F��H@H<W!�I/ �(I��KC i1��'}!��`R� kDmK�w�j�Bs�`!��W�,S~�@d��@�Na���B�!�dR�I�"ݳ)��sS\X#�dՄx0!�DU90rl�2�F4Q,U��dF�3!��3<&�X�r G�"[&D"�d�>	5!�V�J�,�2�az��o�!򤓬sP|��k\�	�d�1b�D2!�y�8C"�#x�����'��S<!�GFCl=��� E�4��� Xg?!�$6k]�%���pV���H�f%!�W�<v��d�RBҽy�x!�Z�n��!�ؠ=I+%��P)6m��'_�,j2�R ?�|����&q�J}�� ���'"A*v������R�VM�d��p� �L���0���t3fU��!�©��T����0�i�r�%��&��d�*�eH#_�e&�1��Iv^0�1Ɨ+;�.��$�Tfw2��ȓaO�(�� ��,�eY�l�9EM D��ÓdY=�� �ȟ;c�h�dc D������T�֨�f��h]<ruG2D���@����1$�۬m�
��N0D�L3�L��VL"��l{
L�e8D�`�6,��6��n\�p�$�0%D��xף��.Q�}Rud�!|sYA�F#D���d"`��`�X~y&�{"H!D�����́H��F��7$��Թ��:D�,����v�2AB�A�9#���@e�-D���4�$�)�
O eH��g<D�0
 $GtWN��Ԋ
5�ڀ���9D�� \�JP�]�(������:=��iA�"OtD`ee�-�ޑx���\O����"OH��)W;&U(4�@-@�e�TY:�퉦��u����,�>5a��,+��qIN�$`鰊,D�`�í!hz���??�HcT�jӰm�u�M.w�8M�ק�i}���i'p�2&I��NA��Q�˕�|O�dj�'\����J�\�މh5j�h|�M�u0O�h�E-�U�J	���[џ\��b�	nb�A�_�J��a8�@6�OX�������Z�%Ǻ)�Z�RU#@<,�BL�_|��r��i؟T���2��y��JB4]�%2�)��1EB�,��Pa-4Ż��j��O�|z�G̟"#�5����O3��)	�'̠���,�b��3����)'����)]�Lq�`߿v�\i�"BP��h��$�KU0��A�+5��c'N��!��g;�|Z%���V�*a�Q�Z�B�a�CI&Vڑ�D+� ���ϨO��#�X�x-�D����0�'�$�I��L�DΦ(��#H����e��|-��y&
7v٘��1��(X�a~2�A(@J����,ۦ%��ذ���'�,�S� W���M�4ID S�A�|�w�D$�)@F�*fO)�'�]j�<II�;
N9Ȇb��Z<������V���{a@� j%�t�uC��+��B���p�y�ּt�&eX2b;X�B�)��0D��JK�5E�x%)BD
@��`����)w�.Y{��'O2�hdJN�!��iu�'K�%�F�ɩv���Q��Y�$�f�ߓE���s�Kם4@��\���q�f�2����$e_ޑB�h%i"��d��|n���甒���H����j��P�m�d��P��"8Pu+���L��iW�iʠu�.��Ѡ��$�!�٪7�40cc��{�2�� ]�3��R0�ɂ0?P�ӧ�B�/ƍz�'*�H�wj�=S@�C2��N\��;wo���y�#�9U�j��" �G�*\ E��*5t�k�+�=$<0�.��]*L���\�<�Wǐ/0�������H���#4JWx��T�Xyx����b�H�b�)eO��� ��	rNy��I5(b����D�L|L#$����評�%�ўH
1 A��59�̇%(qx�P I�?����Ǧ4�]��ua^�Q�d4D��9shE�Z�Vy��4:b�A���OR���JT%o�}Q��A'��S�ӊm¦(sg��N͚Aŕ�?�z�ȓpٸM�+Z>#����G�t�*vҪQ!�kZ> ���e� �s�8���[���bkn?��e�EJ�2L������ײj&:���-�O>��v��&2$¸c��	qR�$假\�&�y� �8<ιhgA��BUh���ޟ��c��t\�0de!扣>�'��!͈0��ȆX�b�=��h�Mܵчh��%Ar���ֱ��8`
Al�T��oݥKF6�iH2���΅�O��E�ă��y�b�>>�T���ȲK���B��?�c�U�Z�����H�b\F,� �V�=�Z��U�H2J���zv��1-h��3K�f������K`NHCTeT�3��B�I+xeV x�nA:n]aE��e����D #���&іQ���Fk	�|lD8�9hu9�	�+b���z�0�񇌷y�m�C	�ZG���$شXA�i�'��
�� 鐬&TА	��x]��.����
5I��Z��Q.(8�)�3��\F��y�d=}�	�"4ל��R�[Jx�kŢډшO2�r�ڱZT����,}�B`S���@a$���T���2�	�T�@ّ��(.W���m�u��	�ɔ�p<F ��j��	��r.�Z0�X?A���	C֤a�n��<[�$��z�c"Q�0�N@��f�d�vX�}�X �� 9,씸b�o��C�	&M]`�`�"Ť�~�Q���X1\�$�ǌ$LpJAkV�{b���Ob��^�D��s+�.���7J=�H�Y?HOL�$�S'��~�)�$�8�`gh�>���k�	wi�i�Qc�;�M�Gav�n�rQ.L�I1f�@W��{h�����ܧO�miv�� �͊�A��>���*���3*���l׾q�ى���Y���/�L�¹qC���H<����\����]�1{�H�腡��9�㉶!�س�l@{��A�-�:�ʓ j�e[ �4�J�{0M�9!��#�F�q�M#An�א�cҦ��,��<�fQ!.�D��l�3hkr��o*�!��ɪ3O�g�+Z����A�A����d��3q��R�h4�I$��0K�#�)\���;+���zbMKZ�DCF���8|�V�j��pF�����D�_�e��K�	i� ���/wB���ea�6_ɼ�� �O���*����\���ԯ�)�*1�d	B����	O���y� bߊ0�P%3	�t���ӡGs@%��H
o��9�pA��n�.1"�g��[Ȁ��f�'�0��	�
1�ԋ4`�r��a0�{���9�ł�7�zLe�B(�*`Ǝݯx^T��/��'�֕[q��=�н�ON
H� `�
Oܐʴj�]}���A:p��0��Ü7B�J3�+F�z������-gZ�]C�Eׄ[c�%W�!�� ��؆��8cI���SɃ�TV=(E�	o�Đ��-<�8��h��D��e�T��j�N��ٺ� .G�!�X�Q�&8� ����p���#p��$B�	xhK���7H�az""W*H����G���i|�8Iȋ��p>�d� .|����
R8I\��j��Ofi�	��&��C�ɓ$�Vݐ����-�`|yp �Q9�C�ɠ,���!G�ZDx��c�jZvC䉔&(v�p��\�3&�K�jO�T�zC�		@��� �P.f�D�#��$#�C�7.�z4i���;F�t�oǾL:�C�IgL 1�̜^�L�S�Q8}m�C�P��1Hs�" ,�����f��C�	�qFT�y�π1��tQ$�oO�B��K8Mi&�_4��l�g�O�B�	�|�i��M4e�l���M��C䉞F����فt��BË0N�C�	n�Dq�\7^w�zW!�9m�C�	�_���dրQ� ���ؼ��B�	9#z-���D�>9{	T�xdB�	#g�����ʜAKy�g�[NB�	����g��>P|H�@��8B�ɢ)ڨ�U@ī�$���C۫_�zC��5A�E˄aW���i��"kq*C�I���� ��}O�s�k�D�HC�I-�p�z`e��wo�ͨ����B�I���x���tNd��Ɛ53�B�*:q���̕8�6qTDZ іC�I��nI�r#5�ؤ�!�-MB�	�Hm�=��g�<%b�<����0B�	:�|�`A
��W���+�����C�I;T^�w`��"BE�=[��C��)��M����(psX��-8U�hC�0pC�g��x\���瘰)�@C䉡o��X0S`�'�����>@C�I�q^(uj��{G�DJa��
s0c�x2�f�+|.�`e�$!c��ɇ�+�u��h�L�S����ΐ!o(C�	-0k$q0�AE=un�š�*�CsU٣fRGy��k?���OG�'L�Z}H��%&��3mG�bj]�ŧ(]��%iB�@>�t"f��E�'��)T4���F��A����S�M�t=�`Ic�:iUj�D
�9t�`@�#.�4q��Lߩy�pxp&�c_,eSwg(����w+ǇgC�u9���uv��Ӎn
*rV��@�2xYƦ�%��඀�g4ع�	�em����M�'��Q�\���q�L$
�Г�D�i��U���`H�`�OB���'�䧐��E}����b�.P���5Ȇ�V����|/�(A7ΰ����'��P�2nŦ��WO�:%~� �C�A%!B)�z��-͓z�O�q�8a�pB�J��Re��2F�>�Or�qS��Xy"do�$>���B�a`�@��%M�`�d�����O�E̓_а6i�<E��� � ���㇯�+[��H��B_8FH�D^�|�\ݪM>Y��?M�	����I�Z}X%���F�@��*�v��E��U��B�H��$��iU�|µc�I@X��mI�B�nɘ2Λ�\:d���? ٔ�#$��)��ͧ�h��II]G�V�)��Ԩ
FT����D�ֱxDL�L���A�)^Q?���|�����>��pФ���\����I.[�U��a�L8�c��J�g?�O���'�8�){t���|Xĩen��~�>Ք'��=h��蟴�`�o��VN�5`C�Ԫ >��2�o;}Ҧ)U �6� ҧ��I��f��x6�	�aJ�\p�dߍ|��0qN:[�Ƃ;$��S�O�P����@+V:��D
 (@�4p�`�jǜc=��ȟ�-�9 @l��I&D͊�d·$��	- �=(P<OF�	ݘ�y"Q?�`0�+t� ܛ�i�L8���ުb��'z�d�A�g��O���"QY���(v�`+A�YWf�8sZ��;�.�>��)���~REɖE@03q�M�K�iJccC9e(��ȓ4�
1���7z�4�b�E]5Y�T�ȓyF��ٲB��'%1aC�-9n����V?X�:"B��dY$y��V�k�����z��u���0	�B��N�\�h���2iTX2�D@g�Ԛ'!LY��x��S�?  �C`�-�̘R%J�,�}ڠ"O�H�7 V�$����6�ι2�``��"O�z%"� ������	�X�Q�"O>�1jѤ?WZ��/Ct�ej"O�����\'`�i�G-]�%S�Ix"O�L3��۬jdf5�,�:Q��zT*O�$bT��A�M(�B["�J=b�'�8�RDf�,Gm��H��D�v"xy�'�<$y��C�d)�$굊
#{�Ȅi�'��U�/J�2��"�^�!]�E�
�'�>};�@Έ�A��2g�t5;�'����-��~((�[sčQ�'z�DAv��Ot����,Ml�@I�'�F���>h�59��(6x�'�����+�@<�'b��
h��B�'d�;�J>�^4�r,	9H݂�'_���V,\�,��P{��O�f����'�l9@�-*����H?0�A��'� ¦ϹE��5d��"#t�Z�'���IV��Rμ;s'��#$��'�:��r��U�6jMU�g��	�'r�t*�`�5�D�b�� :`0�	�'��	�kGw�ر�qK��x�@	�'�ș�jC�#�E#$
̏?����'x$e eUy��RDc�1�<�Q�'��-�ad��I.�pcB�ʍ'�$l��'����R`���ys�+��@��'`�
P!�X<�a�,6򐨛	�'fT��@��JZF�h����z�TB	�'��a���4���Б�y�r��	�'�����A2v6EX��ܱnt���
�'�p	@���
-���J���	bm�	�'F\h@!ʕ����`UL�=6n���'�"�x�+��`�
uo� >��2�'�d�yA���y>d�R��R�~��-
�'c�J�!Ѐ+������ۘ%YI�'�P��4hH�o�,�B�N�!c�$��'�ҭ�F�g��Ep��?l�D��'7,Cv�AO..lRwp@(�'�z���]��1�+S�(s���'{���ۥ3�n����p�� ��'I�1"6�̏YwF|��	��h�l��'JD����&���@ "ÓY�F�X�'�9�╁=�s��9F��%��'�X%P��ƎAp�#D�B�Ip��

�'V���Ө�]EH{�J�<,��	�'O�5"Q�˘Ґ{#(�2�%��'p.D��E���]�{�� A	�'�d��%DF�v��+�BڋF�(k	�'�,�;GF�+/E�"f�9;��� �'T�C�)ɨ|��Ԛ���b����'3��#�Ɛ� �� ��)Ub��
�'Њ�dJ�`�\�k4!_U���1
�'T�m�d�	�0������-E�H�	�'�Ȗ�ٕ����$9�l @�'���z��O/%p����,����'Z��bF�M�"�eRa@("&��+�'�Dт��"R-B��Ed��L*�'T������1A!E�5�]�(5rܠ�''*�CR��� U���%*��'�E�F�̯j�ڀ;aE�*$R4��'�^�+��;+*<S�Ʒp��L�
�'�̍)�d@H ň�!�2jg`��	�'��\Q�Q�����
�o���	��� zɡ�O1WH~�2$B��s�@�Qp"O��YЦ"
��``aEwC���"O��?a�D��[7'0䌲2"O����,�26�T[4��%	��۴"O��k�B*���G�L6��"O
|�2	�	n��������"OX���O!��X�tÈ�u�<ЂB"ORH��NF�Xrq����	�*4K"O�A�aDD%aL��u&^fO~m�p"O������,*^��D�)Eמ��e"O*E�á�x(��"f�V<�|���"O�	�ƫ�5.����e�ѣo�`P��"O��	�^LWP1��c�L��AS�"O�TKя-h�f��Ì�Cxzx��"O��!KE$�Z��㕊,��P"O�p�p�83��9�u�ҳT�����"O�Q#���"�
�)�F� O�0�"O�����_�T�Ă�]�6i"P"O��1�]�GV�`�p"OhDH��q`6�`�NS�[ ���"O@,��I&`Df���R�~HD�W"ON`	4�Y�"�8�҆�"�� �"O��I���4g�1��DH�a*�P�"O����]�@�h�&(WX��"O���@慷v������=X���"O!��� 6~�yb5d�4jc��p�"O&a+�Þ,o���Y5�w%
)��"O�sj��~��,�Z�{����p"OR1#��jf%�A�9�°�"O����W�X�$9q Ŀ�4x��"O��9�T�@���;�NT!IV ��"O�Xb�S�;���Qύ+����"O4$�v�G��"P�����٦"O�"#�	Ml�X6�K���I$"O�\бA��P���'=� �A"O�Uaq��5	�Ex�*�� &"O]"#���{I�(B6�M�2!ҷ"O��3�K�z�2��p`��i{"�q�"OnMr�b^��R��/�	��Y��"O|�)s�Ȃ1�
4����Z�`%@�'.>Tq��d!��'�ֱJ�'#]�f��Z�3�O�N(ܒ�'8�X�IL?~ڴ5Ȓ�X"�$���'l�y���et���YC~u��'�tY� �$����N�xT%{�'y^��F�?gA�y{�[=l���'_�%�w��M���p��:
ش-��'��1� �6ɀ�����U��#�'���@��Up����jS?ܤ��'oh��%iY�h-d�����@h�'��	'�0hTz1�Ѯރ}K^1��'Y*[P�Σ]�b�����v�:i��'�dP@�g��\�{4@�#k����'��Y{RN�r(� �3�P-�R!I�'�h���$ƓI��
�U*���	�'
&��'���'�&��rc�$SK,8q	�'�� �C���x�pC�A�9pTI��'/ =�	!ᾌ��DN�7 �l��'�)kD��O2\���Z�3b|)+�'E���5�¤~���u�U[�XԚ�'<��ÆN���TՏӌX�J�*�'(
݀���3� ���OY(%�](�'�8������rqj#�϶�Vu+�'Ͳ�I��aYJ�y���+e��T	��� 偁i]5#��{���!^5ڃ"OfI����N�l �  �#<� �� "O�$�Df�(q��]�wO�lĹ��"O؈���0�Z�Gf�6�p�"O�SB��L���(�'}�~���"O4`�4(�*U�N�"��S(Mv@5��"O֜C� ʬt�D�%`|`xC"O��
�LV�!c2��4�	u|F<��"O��3�A� �9��*���m��"O���g�Z�=�
�k�J�(�\hC"O|p'�i}51Fş�B|�t{�"O,�IG,9c�q����N^�ؒ�"O�ų$�Q�x�,9�B3r�� ; "Or�s*��2|�D���j��-�"O��WÑ�3�0+a���@iS�"O ݣ�Þ#kGН��)~F\+p"Oʈ�r��,�XBs���5t�Թf"O"�1%/�6ʍڦ�āLg��0"Oޜ'�Ye5Z��'P\m(zv"O�X�JC��3u�N�bj�a�"O��be��(�rik�
��xj4"O�P���^ x��yU�M�q��H�0"OaC�"� EV��	Ti��}8��#"O�X��#�
.#�(:��23��d"O6�a h 6b(��T�L�b'"Of��5n�30�s�DT�Լ��"OR��"��2&��&E�41dq�R"OH��v��n'>Iq�?��7"O~�a�wl6������"O�I"�D!7<�K	�9H��IS"O�[��^�$���*ܙ%3�eR�"O(]Kw�	8$��0lxً�"O:���DN�=��
��,�"I§"O�,�'�R*,XA刄:]����"O�������nֶ`0�.�ջ5"O���WͲ¨�ɢ�M-	��1b"OɇAз/B>���ڰ%��ͺ�"O0(�V�ܒ)9��r��Tk�"O�a�I�W` �D�V&b�l��"O�`���@��1(�
J�b��@
s"OvI��M82���H��@�c�^�`�"O(�QthM�ha�%��0~`���"O�dñ�� V�ĸ���2Ŝ�!�"O��#��R�$���`�)�$|��"O���K�;1C����2�-r�'�"�H�)��M�m3"�����	�'L�#w揄A�&�qFb� /L�@
�'�t�1#�>EW�%��Gͅ�� �'l��F�32�4슁gF�|�(�'�*h�ƈEQ�j���M��v�:C�'S68s$#:�v�h�
��t&Ɖ�'���Z��--�T",G�h�2�R�'V�L�1�L?#�9�̈R{!C�'b$Yp����%�۵ �B�l[x�<q腇
�4%#�h�*.�8��fEr�<q�.T')�&�qa��P�*�)��j�<�!�N�>Ob��4C՚T���"[c�<��N���3�꛲|z���I�j�<�v
"�� ��.i�n��f V@�<�'i�''�R���,��]�n��+a�<���&��d�L$s���VCRF�<���<:h(1ХN��WP��x���D�<�½Hb�ڢGM�1��x"��C�<10�I�p��Ũ�"�)#��� �o�e�<�E �P    �   `    �"  '-  q7  �A  �M  3Z  �d  :p   {  �  ��  y�  ��  a�  ��  z�  ��  ��  3�  v�  ��  "�  ��  �  X�  ��  � $ f � � <% �+ �1 ;8 }> �D �K 7R xX _ �e =l �r $z v� �� �� !� �� 8� |� �  `� u�	����Zv�B�'ld\�0�Fz+<�	�K*�ac�'b����F�|�W'Q�H ��M��uA�-�������ú&��P�h��%N��bH��J���[bo��u�E�"g�t�x�tB�J1��f�q��)���=�j�"6�._>�R���VD�!�F#\��]�r���ʟ�R&e�#�~��ر4�}���Ik[�4�GF��?Y�0`�A*��y�V����'~2�'�bl�F�,�*/hB�P��]�F��'�R�|��˓�?�# 5���쟘�P�Z|����>\5��D���������IΟ�	Ο�iG k�� C��f>ԃ��
-��Z�̊,�@��@B�]����'c�	X���Dy���	�4%`����3��UK j	�er\������~�-��R4
6`%H�ӷ.��m��ƀ5g�1ӆ)�!��d�O���O�����U�	ԟ�OJ��G%J���"D�<��Q��!ں}���j�D�l���M�S�i���h�P)�����Cd�_��(����PC��iґ�5/����Z�HO��T��!s�6��u��W�"b�$hh���?\�q���$� �uM�~��y�'@E���O�i��4��O�Ը�>]f*٥{~��amZ6v��h
s�s�$�6�Y�F8<L��N�Ya�}��Z2_�|Ak�Ì��)�۴c��& �cxta��*5$�\)��٩B���/�%KB�b��iӦ8o��MC����1�r����H�]�lm^00_��0��	/��Tb��ʢ ��1#�%I�u��0A�N%2����u��pm�<	�BX(�f�\MV �A����&�2(P�F��m'z @����HdXٴH�.��rH���AJ�*hp����'����A�[�9]���� �:��'��O����O~�Ě�A�Oǈ8�F&>Aw����o�3j�d������O��d�O��`�ݕ�𭺰
V0Y �r��8��1paV�RŚq��gY�@�R�D�4yQ�|a �[<e��=	��U�&��@��
?�`a�%V�vk�ek�dբ\ ���%B�0Q����<�$W��hAI�U0�XqiY+#��!�%�O��D�OؓO����O���?��ͷ%&���֍��գ����?���"�0��c������|�A�'���Kek˛;�����.��[�����O3|jr�oZ������w�H���	�Y����ΈL؈%B���?�͖h�R@����H`A��D�j�beF(F��Ot֒��7i��Y�~p�)Gte�	(pڴ1��!�6�(;��^K�f9��-�Ϧ�O�PS1��(y����#��� �Oxɕ�'�f7��m�O��QQ�nt��mQ�W��T��A���'���'�"�'�>)s�S�"�Q��F�>��p:a"<ړ�?�$�i+<7p�nZ�|Z	�q��@�U
�w��K�'^6�MK����Ė���	�O��ON˓�=��j-tҌJ���1WZ0L�잊��Qڅg�5p �5Æ��)���챒*��;u�$K	z֤u��BO�:Mr$`#�P&4�R 1떏0C*L�����6�Ne��i�N�s�'�r8�CK��n6��nõW�FpC�i���r���	�?����<.��CP�)C��+q�G R�� ��hO?!8�MN Lf��pdֆ �8B#�ܟ����M�6�i�ɧ���O剞	|�=���w��0������5!Z�����O����<�)�N�8?�z,*u%׾*��)��^�|�|��!_92�
Q��r�H��� ��. ���v��+^"�ex"cT�A�D]�!LOT�h�$	*|����X	3{4����Q#N��!�����iX ��	�?��d��O�l���HO�"<�4#Ǩk��H)���}�X|�dC�vy���k̓m;&�[ՏԗxlnC�ja}'����47��T�C� ��Mc���y�,��Q�")p2㒈JȬ��7ķ�?�-O0���O\�!dRL 6D:J 7�_U&Pk$�R�h)l(i�_�$�KT/"t<��e+ʓz'V� �S�t�37)�@[8ջ��;���`�D�:�F�A�$�؂l�#�L#��J>�3̟P�ڴK#���'谺�g_�,���vE�M�X��oگ�?!I>��oܧ*x��p�.=U���$W�N^���?yI>������ߦ-b��ӯ})tS���7`� �%���M�C���!W�5;jI�f��0����?���4��Ŏ�
-��kW*���Sh*�?����و-�L���9wP<s�;L<�h@�L�I
h�0��G>���'���"�N������O��b�����$i�x[�*�N�����&0���s�U���#�*K����ثt�b%u�f�%>��|� +H�MA�i���F0ƹ"aRK���p&�������'���u�݃F�6�ht�!#�2M��B �n�¹iC"eq�Z�d�:<�����P�|�	@��>'�l�şԕ'��@���OB�'^�[�|@@B:<9a�@�
f�;2o��0H}n������aӖ�B�_>e�S"c�m1ͬ���2��)���qBK*���LP��o�$U��D� |��-S��e�OR��9����y�IHe�(U�2+ �:pe�T���e�<� H�ҟD�|�	؟`�I X���ҨN�	b=x�Ⴘ}Y�%���	�i��$sZ�`l� $6خ���O�mZ��MCJ>a���(O(xy"�N�A����m�\�7� m���l���$�	ȟЖ��O����A��(�����Īo2@
�8.�N���͓�lH�[��O�PV�0��ʙ��(O:�@k\"3�|�xU���,��� D�� �1
񋅜G�,�k�Ѧљ��ԣrF�a�`.R\�	"sF��aaUhީS6��1_VJ���
�O����O�,F���ތ$\�Z!�	0��%kp`��=1�y�͉BaJy&L�R�܃wB(��-��'}剢g��Xi�4��	Ɛ+�x#��7:���p.�<krX������(�'7�T=sKX�bG��+:��� F��d�Yk)��)��E�sڴ�B�H#z�L9���$\jM��`	IW�~(���2� ��Q�ɒ�AT*��1��º'e�cb��1v�%��{b#�OHm���dܭhA�Hf\#���pW�>�'���G���t�G����Rp�fn4���c#��'�ў�s"=�F�=�X�x�I�2K�{@�Æ�MK+O"E;�o�æi��y�\>]��?w�J��Uӈ:S�0"ҡ@,P20���ş�0��8qJx3&�	�L�
�v�����Oz�B$��.(�v]�S	���XA�Oa+�!	6\�Yp���F�z]s�6�Ӆ�����K��$��ɗ�
=��޵�i�6�'�'�?���D]3�FU8L,1 0��68���ȓy�� ���J"g�!ТBۗ���D�%ڧ#S~�%F��q��+��#X�
)2�4�?�+O��cM���O0���<��� N~�[ş1wX1ђ�߻��D�O�u)&�'LO*�C��^$4�.Q;q͈�_���"���7�0�C��_����{%nܵ:�1�
D���p�C&M-H���	�dS���F���)O�����'���?�O�h�eaǢV��M�df�}��k�.�Of�d�<	����OS��	U��9�EA�c��=��K�8��ʓE��F tӸ�d��9�O��d\>��FN�{K���d���:x�bc�(**\��4�?��?y*OVʧ��$`��֬y) ��	f�ڈw8�
�'�@dP8CH!ց
4i`���F�;��́�Z�Wq�%1��J	u��#��d�9\z�)�̌?X�T����7��P#��''�6MTL�'��DCB��	j~@1����m:%"f�OC�I�Qʶ�2tM��u����OX mZ��M�+O8�a&IFҦ��I�<�0]��#�K �i�\(�ş`�'1b�'v���M��'w�`�!�5:�M�:N+�Aʦ��#`ax⋜X�[P(߭>���p g�41��0@��3"Fx ���3�ʴQ�đ��O"�z��'�>7�zy�`X�=�_1� Q"��䓂0>)SO�fl�4��It y���
gy��'�47�T,~�<,4��J$GټP�p�����y�'��bg+e���O��'N���#�i��� `&��v���F5������?� ��%Y�4y7eMI6����<��{�n4��i��u���K^~�&�����*3L��(�X�T�N�E4R�����C!�u:�/�>H[4L���@5(�^vu\�֪�\�X�@����'�O���+�'�y�B	Y%�ǡ�Vm�Bo	*�y�d
~6(`s#�%M[���$�D���O$G���Q�k}�q��7�����W,Q؛��'���CB$�ʮOZ���O��k1D�����5g��Q�g���, *O��$�=Dk�$��p�6��a��O�
�S�	�}�l,��ΆtN�W����i0'-N�'7�bѩ,O`�
��ƑM�0���l��0�&X�C�v�)�'�����ʟ�'K�-۳�O�Q��1Sj���(���2?������V*�16�B&v�e��G65/剤�Ms��iu��z�@ʧ�"/���X�f�H��tJ�rm:����prnx�'Q��'��I`��1��0:��S~a�If�ܐ��'�*ZҨ���)�Or�HԠ�kԄ�J��\C�tY�l�#=����� cB�
g� A2�?��Y�dYIk`	kԌ�>Ք�3d؟Գ�4D/��H�?�7���(C,��B'��p��4b����?����?y�WE���P��<}ʘ|p"��p�h$���ڴo��FY�T�5`��x��̟0��>z8�萪\�>�hs��Xڟ��	�u��5����$�'5�$#�)ب0t�zs�ՙ�Mk��80��R�ZD6('阔w�"���w�'-0��ɟ�m"v44oՎ@����i��%�V�5#�n}�l':��	��O��[�x�B�)^�I��J���O��B����
���J�)H.|���'���94�@��!�Z��F(#�n�+ ���]Ɵz�
,s��paaB3}vp�����O��0�4顺i�"�'���o V����9� �YFE��G�2��/�|gԍ�	hC���Z��d�tD�!	�ҙaE�+u����&�M��eL5�(]J��	N2���1��8��d�!%�d�V�F�U�~<�B�%q�:�nˈ���X�dxj��N�l8���vnQ�W���	�p��	:��S�Og����S�n�˂�׎M����'R�u+� ��dr�,����t�����D|�O���e�U-\��Y�q"NBO��3�i��'�e�"�O���'YbQ��26���u�LT�)=Y�RV)�'P��X;4��1j���x��O&f����|Ra�C�R�2�	 ��"Ӎ:I�0x$��X��s�/7��4�G�FG7*1���<�pV��OZ�Z'���/�t5�Ă��S������uӔܔ'�*�j��
ȟ�'L1K҇�5H�P5;PK�c���U"OB��g$Z)~��C�nv��D_����4�����<ɴ��}�h-�w��r(�1��@�v��[���?	���?���{���O�dz>mkc��U�4��3��|� ȃ�)@�F�Xu�^-e6=��H�%}t�s�b�Q� XՌ3� �L���ȡ	�d�9���#�88�ʉ4�L�q	��L�4�-�N��Ccĩ*��$���c��c&�`���=Cj�Q��ܷWА�dIʦ�����/�.D����ǣYzI�2��_�&9�ȓFs�]��C5X��p����'�T�ݴ�?�-O�x��$[|�4�'�Z�6���J��t�G.)���"W�'�&R�#���'��F�p��:��K&
�J#v�Teu��)�'GF� *�"#U�;���x��=	���*.����*  �9:�nQ�B�`�cQyz�2�׬$Dz�6@��K4�a���2d��Q'�tB��O�Qo���d��!)����%YyX
�s�#�+��'Ka|R-\-���daȇpF����O(��?���'�`�cD�#���a�u�X�����DD>dR����O���|r�
^;�?�C5_��b��U{�t`��C�?Q�^���F�GQ�~@H`e28�(S�l_�oz�iΟ��c*�+��`��K�$7�^�����E�Z�~N%3�'�Hp�ِ1\[���~�t�W"y�`��j�.3z�q���L~"a�:�?q���h�j�ɑ9Xj)�v�A$L�8���E58�$B�ɝ>���q' �
�1 8sV�?���Ӻ����d����� �Hؗ�ܨoZן��'�`L�O\��'��Y�D��ƶ8�`�cU�̮�
89u��Wyb�'��[��'�\��$�)2�E���(G����͍<h;J#�'vx0�q�D6��Ϙ'Jpy�V�I�Ga|�����XrD�y��i��������?���o263�G�;��0jt&ߓY�������?�+Op�d+�3}B�#J����k�x<��M̌�����ݴ���|��'���[�w��x�l��N�����4i���5/ܚ3�t�D�O��d�O�|���?�����ڧ�x�(�?Z�]�C_�a)C�^�M����F�'�6�ׁ�x�N���
��$aإt�
�Z�=L�3/	ytL���A z�'�+tj��@���(7��0|��&�C��?��'}�ԛѯ���ʈٖ�HeL�1�
�'�����\=���a �HH|<�L>!��i��':����,�~b�y��Ii����fY`��V#l�8����?IG�M �?A����b�-@[����$8��k݉m*!�ō�]7�mZPh[�X<���]�b�f�FyR��0iXR�"3nhf�ݪ��YKL��3L�JRRy��kC�Mep�����LDyҎ��?������$�hT���I�7��,�&�+�P�	|���l��/P*�H��^9P�Hiʲ�8�OrX�ɟ��B��$I؅z�a�47��Ĳ<��*KS���'�Z>���e���|rP/��is�TkЈ�_@��C��П(�I1%�0�@��
� �̋^F�3���p��?]���� %�abQ� [��ex0�'?�6$�����"Ȗ>Ȱhh%J�{B�nM6��$\ � �t� ;�@$�-%��v�	��S�O-F`�T�$����$�ʏR�X��'��c�b�N��$�O��
�Ls��dt�Oڄ`�C�K��s�шo��x��ir�'�2��t�*a0 �'+��'��4�Nx��8'�D���(�=�}��%H�~)�U�Q����p��}31�,lZ����0<r�za��Q^�8�#�˼Nbᐑe��,��T�v��3
Vn��iD�y���OJ���Y�j%pH���_*>A(;�6�d_+>G����È�V���O&�B��.=�!���X�*-3@C��7C�����#��ɲ�HO�I(���OBT��WJ^�
�:���ʠ�#�F_Q�����O��$�OL����?Y���T�ĆdO���/
nm���S͋�\d��c3���<�Ⱉ��G�X����	�,X��@�Mٖ͸H�7/��e!��n)�y�Ո���b��S�'��� &K��ʸ��gآpkl� �&ܺ�?���?1���>\�l�+�`�2��i��I�O��B�IT������g�.�ZƋ�$��O�!m�ןH�'#��+E&�~���{��	�qE��#4BC���('�1��?٠D�0�?����D L+:&,�S���P08�!L��,���AA$Z#����V�U�׉� 4r��Gy�@�mOab��R +"Ԝp%�ޝ�Ѝ���/"�vP��W�u�Uj�� ks�DGyBgO��?�������h�b����N2$�*�0�L�h��'���'�4���-�[��Ӎ
{�L|���i>!�bͲm�V�h*,HUO��O�v��	py��)�>6-�O��D�|�M��?Y6�W%�t�;�)4k���C:�?���;�\��&M�]�z�ڗNٸ��(�P�u�	@3�:�ˑ" Ft��D��f�c~b�A&"�$	�F�I*u���{��Z��ݥI��'mҴ�G��dKXX(`�M`�u�'Ξ���������)�U�T�{�^��팀bҠ|��"O�%���%;���r��:a�$C@���h��H  /�O���y#�],���A�m�����O(���Fs�u@ �O��D�O��Do�!�p�J�<A�y#��=B��櫀��fP���7w�U+d�´a��b>�Zwi�.V����J*|��(N�L��k�`ɹW a����-�,�cgF>pD��逥@j�,z지 �`���DpD1�oU�U=��
W�2��U�U;���Z(�$c���!
J�Ɍ~�!�E	
�R�2@��%q�:��S(O	A����HO�	?�Ē0�R�qP@7	@�hI� N�\�bq��٦5��ޟ@�	dy��HޓbKޝJ�/W+n�&\�"B o>���mв4��5B4�L�<r��Q��5�h�6�K4��R�>�q��O�0Ј� 5��r�<�j�\a�$q 
���Oı� �L/��yeJ֣=��{`���I���'{���-�'u��p2�-��QuT��.߃C�BU�ȓ��� �%D��/!����S�.�ͦ��I[yRdB/P�j����rGI�?���6`�8�fa٢�'��ßL���T�W��vZ�)G�/b6����L=m���;�ʶFt<a��H��;�P=������a�uF+� �C�-۴���Q��O�kF2�˥F�"�*�`È1�<�����X�'����� �2�KQI�2ڕ�H>����p=��2�N5�g�l-�qIA�"�Oֹ���YP��D��4\;ph�74�<�d�<)�U�,ߛ����Q>I�I
W#�	Sd��7�����������8{#���w�8�J�c �lM��+G.�+��O{�h��-��ˌ|Ȱ���`�:��O0�hc�Jg�:�j���
�f��4�Ӥ<���6j�9&��H��<�*�pO���ڟtE��'�$�҅@G�SF���B�<���"OFE� E��t+��E���8	t��<�h��YA1��s��$Ӱ�X4��t!`K~ӄ�d�<�F���z��?����D�$I��Y�! ^(���yU�ѳG��ѓ�jW�
ʙ}!�0�n�8g�1�H�O���6h̘!�eS#��d酬�4
�~ق�$h<H��F�N�1���O�4{�c=B��}+ƃCs\4�#�'�����D�OX��4�I�A�*�aA�Tq�"i��#b���ȓWLB�	��s����$�BY�'�0"=�'�?A,OJ��T �"y��8���R�J���ŤyL|(o���0�I�䔧�O)�}*a�C�Eܢ5f*��D�l0X) ���X5�V�C�R�c��y�ڢ?�qE�29�z5q��.;x\�J��PF�z4�@��.�us�`	5p�� ���ùN�Ȼ���5%�b���Ξy	�h �'7��H�'q��BȳK���!�Z�ȃ�l.D��iQ�I02,9�K�l���X%/,��Ef}BS�Ժ�A����2I y�A!�%����WtM��cy��'i2�'�����F:����p����)������"°�0S��?12`�w~>49��`�����H�0ܔ�aG:xE�4 � Vcpp����P�5�Iq���'p01�A�(v#ك/>�ѰN>��K*ai�'N�n)rUa_�
�,��	��?9�m��@	��'ԓY�d�3�oB����'(�ثϤ>�ON����A�\%)����@�@^�r��t�����,��$��.�'{W�M�mС������n��0�h,��`�p�	G�^
���P�%�p)��H��6�.���h; mZ�?mPf�9B��Z��I�Tka1?�$ڟ�3�4 �>�'W�F��7�±P���0Ӧ��aH�ȓ	ݞ8��j�{!���f	F�\]4GK!ڧO�l���F^d%�#�P�r���O��r�f�j���?����?�/OX��vm�	�-�
N"8}FyZ%�3�t9��G����@a۽l�c>1'�hx�fN0%H^��ʢyLP����$$���
v���T����b>9'���Ӫ��<�L�"U��5M���ۦ5�+O��hR�'8��?�O
`Q�֦j��eJ2ㄴ%d�)c�$D�dєjQ`@�� �[�������<y��)�,ODi��@ "`X�H�g�se`A@0�F7mZȟ��	��d���O	��rGۈCa��c���9����Ek�_�fE9�@74�J]��,��b�^�?��Ù��,�1J�Lĵ�� ��i>�ؑF	�.c(P	��ЧM{�������%�L�c�̀+�d���Y��m��'��6�Z�'���z�h�]pp�AWf�/]<��0D�HhR�,���5&�&mXV�:��J}2X�L�+����m<J]��bÖBH*�0�@6N��l��qy��'���'֨�3���e�Lҋ�<�d!�fMU�~mQQB�=I��\���I+���?�wcH�]�dAp�ef{U%ʵ]3z�j���$GTE!�#�:軎�D��kK�af�|�'���pGā�:�T�sa�<A����L>��2DX�WHW�eo�M;����#7:a����?�ӎH�;Pbآ6�#�N)hf�N���',�W��>�O3��@�vV�GO�{��S-	��\��i�ܟ$�I>V�5�Cm���X`5��>s;����D	�0F�����GRM԰�
!-F���?6�z���V�2Sر;�/�,�?aY�K��аI�!*A��2�#?�Q)�럐��4KK�>I�g�? H�
����W����G2OO��B"O�����P~��2r��u�j�aB�ɰ�h���� ����>Q�Q$���Ȭ8 ��>!.O�8)���~���OJ���<�1ʝ0A�zY���C2q=jq��PŜ:w+������E��*ޜ�x��D�|B@�e���y��ϛ�dZ�Kob�y%L�!Xh`�˻)�pQ�����|�G��f�������2*<� jM4m�Vĳ<�a�Aϟ��Sp�L>iv��jҐba�׷����IU�y�QXEB4��&&�F�� �פ���o�����<Q��V�d�"����5.����1A���2�i���'�2Y�b>�WB��n�)�����IZ��H�! uZ�Lb�![�j�}X�Epl�2��$X���@h)i�B%_,���@�@���d�5$T���aC̑=bџ�J��^ZBX��`�U�Ǌ2UB��$�Ħe:���2V�]q4+�;x}�x�_+�6��D"O0�k��8�� S'�[�q5,��|��>�)O���7M�Ȧ��O��-�F�����j� A��hOV��$A�"|�2�܎7 !#��G*ԭ����m���Î5�gV�]3c�V�d,�E@�� ��(��	���DTh��p}^����7D����cΉ `LB�I <�dH* @@�"Ү�Cvl�$���������Gn�7Q.qa�=HGrd�(>�$��a>ld�>�}j�;ptp䲁"�+�b0tK�w~2�.>�Ea]5P��@P�O᮸�`�.�A��[+d���O(�� 
�F_ ӑ��-��^N�O+�lc2i�7"����gJ�r)P�O�p��'�6MN�O��I�1m~���6��gHjňtA�3Ty!�$ף׬HB�a&�*!
bKJ�^џ�H��	�!W� IC0�3Ir�]Su	
"WVr6��Ol˓Q1,��*�Q�8cuj^�I��Ҍ�8P�҉Zb�2�	�g���Dĺ/唨��Mɝ}zҽ{P��>H�1O\�'�,�Dj]Z����R���A�|�-��?���y"(�*Ck��0r''M��P�B���yi��d|>��oڋ�^8*ء���S@������uk�G
`]�d��T��ؘ#H��[����^��cN��z�:B���T֛��+_ ��2�2�@���0@&���$ރX[4W�'`��*�'[��'5���`E�"?���ӘHiܜ�4��;���F&8pȢ5hD�Q�%�A!C���(OĔx���#`�n�XC\�	wf�r�
	mB���:k�����!E�������(O�����'�6��J�OV=H�D(@b4:�
W��˓�0?��b#`�M�sd��/r�qu�DQx���*O�EbFEȠ3P`�!b�'c����U���fj
�M��?�+�dl�D�O<��1r��%˒*�d4RC�Ow���;^-`��я�:%B�X`��B��L����fb>Upe��s6΄����d9X��2c}�@A$ā�(X�J�&�E�y&�ԛD6��c��ħD =�U�-r0X��4�u�Y�_6�E�������'��$�v�~x�	P�� T,�!�dW���,g���o�vMC��>�ў8!����_����t��OP�C֣���D�O���Д#p� 3��O<���O,������đ<BF,`*�m@
�	��^0]5\MB�Ͽ��Ph�  b0���g9�3��/�'f��y���-��� �%fHԉq`ҁ0�$XA�]ت�@��)��0ܘ%����/2a�>lr��ݜ/���
"?��"��,�IH�'"�D��t@��lϰoU�a�҂R�b:!�D��S�ԭ�`j"�Ҫ�l���3����ş`�'�z�ZU��D�:��\�R�c`W��k$�'��'��O���'?�i� ��	Kի��:^@��8�:�� HDS��L��ř� . ��s�0<��XA��dC^�����;�$vM�ts��a�Y� <c�nM)U��b�؁DN���T ��m82D�xf��z�D�Pc�N�2�	@�'t��V�	+OB��F"�*	�r�
�'Wh3��. s(y�U�>~zx 9,O�1n쟐�'D��5��~
���L��#S<���Z�^zإ0Ӌ��?�VJH+�?���?���Y�X4��ާj2}3�
��8x�lƒ
�&�#��3>Tp���;���DyRoF>��p@�V�w��;��� �d�åX6{�x`u!"Y
�˄�H5Tݲ���b��Od��5�'���i	e�dM��HQ5iP���'�3��g���� ��S��ƫ]�#�S�?�O��'v"��cg�,�p�t-�9<���.Oҝ)���������OBtG�'�2aJ�\�C�"�j�\Ir��u���T#GL��F>��Ԯ�>%21B�]�d�?Q��eK�VwW��w���A�*�yRG؀qZ��S��-�*q��N
J����%�F���~�`f��H��I�<:4�������<��̑��,��a~J~j�O� 2�q�ڪ{;���@мz�q��"O�	��EÇ*�L!33�<��%�t�	��ȟ�L�`G#_і�ൠV'm����u��O����O�e`��'tf���OV�d�O੭��?�W.M:]p�bŊ�_�<3��,�8|��A�b����!K�Dw���̟�m�s�����	S����$��Je	�タD�&�$|�"$���`s���������ɔ6�l��S�(��n
/Pl�=��&yC�d���wc��L�����O�=٘'��L6)7c�dY�O)$K(�	�'n����#��Tub��F�"��:�ő��̟t�'�5i�����F��e͂����$	�;��y���'ir�'���d�E�Iٟ��' ��HQ�.�?&A@[����DN̡*�Ӧ
�Z!RFI�S$�@aGb�7@���o8��n�+�@���d�B�ϣ�X�u'y���J+uU�tc2�nI^��t��5��#$�xL��?�tZ٬�r�.�?��E��܋4՛6f;���O4Y�Ć�L]@�gc�����T"O@[�h�h6�ۓ��戩%^��#�4�?�.O��B�Y��'��)٩,N����C�R��������I�@��O�r�'z" �=aJ@�%O7t� |�@a�stX%s�'V?|�(����=Ѧ���88��I���Q?q�Ė!39�؀���2���׋�=K+�	0�!һ��Q�%���f�r��"�[�'E�	���?!��4㐊:�ex`�I�F/>�J���&��$!�O0���H=^�B�g�;HL��b�'�˓g�9�%Eƪz�|YrF��Z0J��'��'��U� �O��3O��b0��eV�zJ� �P�RP�x��?,O�է�O~:-(�g�H6�����<�D�C��S�ēx=0�/r �&^����c܁x���,w~R�F�<yVk�g�T>�	6f|i$�"6\�c�����B��q~�:}�D��I���'`�֑��ߥy�hLpf�߭Xcvm"֍"}�쨟TF��'�p�
vNԁ֞�(2��@��1���+��	���I9R��'�f�'!V^�pt�X<pI�;u�U%<������D�p�'fU���I�'AB�zA�U:I?�ŁN�)`���D���W-�U�&�O,�m�Z�������>sUx���S8E���v�ʩ�OD���'�>a���%F��wbT�TY��i��٤�~",�=���|�P�Pa��?1�O�7<��h��H�4G����DX�3���'k� i�O� P����<8�����4j�b���ŧ<%��r?�Cȿ�?�K~�s!<��<vV�yn�U�r��H6:q���	�qO��D�O���7擞�fM�D�@�fE��C��RB�$"|>�R��M�\�!��E�S9�7�O��d�O����<���?����?��P�����hN'6�Dq��D5�V�'U"�'�b�|��Iِ-t0��AO�;G���!�Z<8���'��	͟��ID�d�'Rԟr�+GJ�8f�P{2fJ0$�M҃�i���'d�'��Od�	�8a��1�#Y�{�`xy҅@�FF#=��y��P�F�V�<N>P��-�n�o�Hy��|�O��P����<t�SA�G X�фK�y�<�௏I��-"��
P�6cZ�<��PRR-��8�X�F�Z�<IgW(#"<�X�J��94��gjJJ�<��KY&\$�֋�!PMja��C�<	���'�	��O GO� '��|�<���hX�SӞ}|�x�
Oy�'=��'�B�'}��BE�:ȭ���y��#t���4�?I��?i��?���?9��?��J4�sW30�.@��U��,x6�i}R�'(��'���'r�'i"�'hn�@Rܛ{jl�qX"(-�dfy�b���ON�d�O����Ob���O���Oȁ��R�E�,`��H�zO�[���%��ğ���۟d�����柤��ޟ��ڈ*�����ֲ"TRD[3	���M���?����?���?����?Q��?�S� /5�	��(K,�����| ��'��'"�'I��'���'���0F�~  ��L���!���w��7��O��d�O����O��$�O����Od�Dԏ\N�9�%D�E["}0�
��z��oZ̟�����I��0�I�������p��2:t�i��� u�P�ٵ��_h��4�?9���?����?���?!��?��9��AK�C�K���(�JM�Fe�##�i�"�'���'_��'���'���'��E��� %�V���(���`e�b�F�$�O��Oz���O�$�O��Or�Y��)���tF����'tmZ���	�d�Iޟ@��ϟd�����ɥ:U�43���3X��E	�"@$8;�4���ONʓ����ͣ �ܔ(��pI����[��<��BvӠ�P�/�S2�M�'�}�0IL�6|(j�h�7*K(]2�i�$7o�$�'f�O��,#%F	��~biC/��q2����:��W@<[Gb��� ��rnè|4ў��<�����N)^-@bD�+T:D��Cӟ�'��'��7m�1O�� �؃��x ���M-,~�Ay���Nq}��c��l�<9.�l�����}B�0��ٚ?Xl�X�S��Y0(Q7g�,��Af#?ͧR�`�ys�Ɔ�yҪװ���r��ӈC��u�+���<����h����Fc�C�*'t��w-ͫ;�R�k��<˧�����4����DτFB����ͥў]yŭ��[~"�{ӂ�m�d+���<z�w��"U �3<~��]�w��(d�H�$�ģB�B�`S�	ៀ�'\1�8Ma�E�i�l��䊉N:.���]� 3۴=W�d�<��TN�I:��4Ƒ8L;��:SCR<���Q����j�@�S�ORl�g[.(H���"�6 ��[�GT����OTd�B� �1`vi�.)���<AR�ێ������J~���@^�?I���?!���?�����d�˦�R��`��0q��0��0lA ,p@P�㟐��4��'/�� �ƭi�:���!@����m�nXq���A ��{fbS�a�$�O����S
�XP��<����yW��~��0��(Ovު- t�W��?����?9���?a���?���׆ɀ������fY��Ձ~p��'$bk|Ӓ�j��� ݴؘ'��|�L߱^�
�A��I21�T���x��c�An�?�: Ț�B�牨H ��ʧOܩ4t4����"Pt������I	!FӲN�'�H�*O��d�O���O�[΃�jת�&Q�Hyy�d�O��$�<��iޅ`�'R�'���n�l8ƍ�x����� ChʓS@��-�M���i^0O���$��IQ�xU�|�N>7a܈�DKE�2��ЈN�sQ�˓���\b(E�K>�
�2|ې�Qvd˴'	04�1�C)�?����?i���?�H~J(O��o�~`%PtZ�7H��q����X@�7?	űis�OT��'�n6-�WS�P�B�7��/2ҨI PmӨ\nZ)g�D�K�"�t�ɔK�:l���H"wY�(�'d�)#�e�?A �[创/�t����'[���X����|��,�	v��@�>��U��.�t�~�u���i�VV0(���'����'��7�p�hA��@�>ͺ��
�	��s�N[¦1ٴ�y"U�h��?���[}�]�@k��F#��a1��Ya���~m�p@2���(���2<z��goS�cy��'��A�-��L�q��7�r���E2�B�'Er�'��ɨ�M��V�<���?�7�����Q����&�
#a�~�x��O�<oZ��M�'�xr�6\n�q��!�����m�0���'�nXh�fCW��р&U��S�gВv��<���$v�l�v	o���� ���	ğ����HF�$<O2�
A��
O�j�E4�HM*��'�6mռf �I��M�b�O���a)=Pj&3���8SX��J��'ֲ6m��Ep�4_фHBE��<Q��6�l
�_�S�pRg�;%��qw��!��A��(�䓡�$�O��d�O����O�dF��J�򉓜Ir��e��[Iʓe"��_�*R�'����D�'��� ��CĨ���2O�|���>��imX7�t��%>U������Zu��M�"���eނ�
W���C��k�ƉPy"(\Z����n<'�'���"�|�3ʄ^H8��Gn�u�I՟��I������p�'� 7�=θ������h�!�"x�y�&��*���$�¦Y�?�GS�k�4;w�<O�Y����fr�ա�KS24�5�۠P�A�'�2A�uS.�"�Hߒf#���?����v&�h�U)�J�x�S�Q-l�����������	��D��I�O��\�"B�o/~������UXx����?���i�&#�����ZĦ���L~r
�5`^Q:��@�x����!�����'�H7�����|^���F i���I�S8�LK�%t'�z�aUTmR�.O�3�IrG��H�	~y"�'��'�RM��t(q����QL�9S7�J�]2�'��		�M��
���?a��?��'��d��V�>���+�0%�v�k��[7���a}�"�`Tn��<1L|��'@���"�7�욤!�2�(4A������������� ��;$�O��"�ؤJ/�y�u.)AG����O"�D�O����O\��Z˓|�V·�	O����(L��;�f��~����'���b���>Aƶi�-`�kG+�FPP7�A�B��#�cq���DA$\��8h�9O�DЎV@��#�^K+&�]5�-���ܵ���fFQ����"����$�O�$�OX���O���.�D%��*�>�f�;s�5s�a֝�M�R%��<���?AI~�c��2O쨐Jژ?�z��r	F�y��i�0�h���o#�ē���'��wշg䴨�P�\��f��&{�}�S/T�.��I��sFx�r�h�/?��#N>y*O����O\�{�`�$g������A8�>T����O.���O���<"�iu~j�T����A����AR:e�d�xD��l�K:�I�������ܴ�yr^>�Dϗ'~pQ��R�cr qm�O���	q� 4D�_g�������H���'��z�t�C�hݓ_xֈ�p���?����?1���?���	i�t���w����@�ҬxA"P;��O��mZ_B]�	ğݴ�?AJ>A��c���Xg�'r�h�9taݹr���1��U%���|Ӗ�DЃ[3L���8OH��ׅ!�>,���3>�Yk�!F�᫓�&i�I�''�ĭ<���?a���?���?y�CZ�4&2�e�<z��qg����d�ɦq��!i���	ٟ�&?�~,�9�׫iw�u�tIŸ#�ְ�OހoZ�M�G�x�O��4�OԢ!�� �	Q��et��+U��=�&Jup|U�PV������?K���eB�uyү���H���U=Ur�	�/�_��'1��'�b�'!�Ɋ�M[�K�<!	� �=3�H�C3��)��)F~]"�'�7��O֒O��'��6͐�IP��(Ѱ(D���h�~m�1g� SҨ5���%B���՟�3%$ݖ?��t��nyR�O��n�: ����u��?	E�����J$h���'ZB�'�r�'�b�=�n=x�HS�4@s�Rg��d�O.�����L-?�4�i^1O�m�B�ҽpR�X#�H�*�pE�=�DHæ���4�B#�&;�Vl��?�nI�V��A&�9w_�U[0���G�`�	�IA8g����K>)O����O����O���I��lʊ@�c��xB����O,�$�<�ֿi�tU��'��'��S�T] ҇�wH�&�.˓a�	�M���i�(O����4�e��kn�@a0m�D ��l�V��-V�ʓ��V�P�PX1O>���>6-�)!���[,���ϗ�?	��?A��?�K~"(O@�o�gD5�%�,uZ��e��38��y�5?��id�|���>	ѸiMvV�<��Y�!nJ|_�E�&Ӻ<oZ�c*ּ�i���I�g`.PA��*2��'�|�#!�$sU��ҍ�g�v�Sv�'�	��t��֟��IƟ��	m�E҄*a�Mj&�K$di~h�Rě�3���"�y��'X"���'^�6f��	� ~2���n�#|�12�
Ѧջ�4m��'���O����׀!p���'�^�!a�`�j|p�J	,i��i�!�'� A�WeC'����|rU����ɟ0�4&�cn���O�L��ty��ß�	̟��	Ey�r� ��t1O �$�O`A��sv8�R !���c!�9�������צqߴA��'�⭘�A��:%2& �4|L��P�':�� �S�}˂�9Q$�V-���Ju
��;����ъv��P��"�Y��N=f�3VI�O��$�O��$�O>�}��'>Ҥ{���6F�vd�gZ����i���F�[��d����?�':����aן^�tː�L�B�	Z�vDh��nZ�y��a��s���I)Z�t�'��Z(���%���j�(��hp ���C�	|y��'�B�'��'.b,ƙ3k�)ɤ�MT�D)ɷ���t�I'�M�&
}~b�'���H+Ѥã0o�2D
�Q��i���{}�v���o����|:������&�^YC�G�#:L�:��7��l�E�����#3������W�ԒO�˓5M�mQQ`䆵�3(P�;q����?��?���?i+O�LoZ�2���78�8A����A�{E�M�a!F�4�ٴ��'F�`��6al�f�	��T�!f�:*�����=`j��E
���D�O س�"�'��L%F�<A�'I!���X�^�31`�!D2<�#���?����?A���?A���?i��	�,<�8�����y.ͨ&�&t���8�45 ����?	6�i.1O�Hk�GS�np}�gfM?$~l�6O6�8��m�N�d@�,�����4O��DJ�֮�� ֌�"T���c�K�h���kr
��-�ؒO�ʓ�?���?A��X�:�!A��#[P��6��#ap3���?A*O �l���|��ӟp�	P��%�-�&4�P��./��"���D�v}B�u�8lZ�<�N|���5�i
��U�7d]ؑB,"�EmihB5��F�Sj���?��햎'٤]�fيR�L�h3H�$F7n5b��αOo�=��*��}�ȓ�v�A����h%���6���F|B)Q�6�H��������gV5[�:��o�ij���a��nn�T�C��P��E24����dr�$1@C�
����MUw�8�e`G	l�����7)�j���R���(�-Y� �R`ֻs�n�@�/�	6ž�Q,�"LUz�M��G��lX�Ƥ���AW�y; А��:!!R�A�Z��!Y��
uf�QP �E�T�w�H�싐 �bibLB�Z΁{uJ��/����J�d����'�*����J�'�9Za!�_������οqE�Ex�h��
j!%���'Y�����|J�Y+�W.�8���#rp)�E��XrP��儞1F!�a��H2L��f�kFv�Y@k�7/`�.1W���k�DƂ��ȓ3@�|��a�ꚸ_'����� wΔq􈒨d�Tq�JK���::~�ó`�e�Q1�G\'^�"S����[y2�'
��'xR$"�'6�QA��Z5@x��G��Jn��Z�V������x�I۟��	7��1��4�?)�4���Mw``���P}K���?Q���?�/O���O6�)�O�ɻb��:�g�'�6��͛?*����O:�D�<�UH���S�|�I�?�k���@ֲ���"Fa��IB�]Cy��'�26O,	��O����73�
AZ_����M+G����Yy��[7��O��D�O����c}r]f�2AY��:df� ���Tb�'��ƚ�y��'��IY�'����T���F�����W*���4�pq�4�?���?���_��	lybAIv0,��!I"K�l}���G9�r*$�y��'���L���?�s�OU �D�hZm`�{�� 1>����'v��'�`JF�>�+O���r���/bE��f���S�H,��b�<I+O�Y�Б���ş,���؂U�!�8�0�:o���b���4�I#U�D@�O���?(O��݄g��L�P��#Ni6�2�<8�˓IZ&e̓���O��D�O�˓P�*��Gc�378�j�φ1Z��� B)7�IIy"�'�	ɟ�����2`R�Oz��cѠ�-��M���P��z�	|y��'1��'��Ʌy�������0��+�-2��=GnM�Ily��'��	쟌����(��n{�Ȃ�Jو��y�$�W7H�I��hFߟ��	�,�	��'j��Uc2�Iā2�h���\�Ex��2o�|�����O��O��vO\I�=�4%�;����G�)�:yPQ��� ��˟0�'�Y�g�%�I�O���YN�4�U#�	�Ԉ�w�A�Mh�O�ʓD*��Gx�π  �P�+ϩj]HQCEg��~c ��'�剩`����4����O���`y�C�=�ΐ���P	#��Yɡ�J��?�+O�1"�)��$�ȑ�� �rFh�!� X������qlş���ܟ �ӏ��'��L�����Y֘��`%��&�~�"Q�'%��#����ܟ���䚰Y�ԼZgj�$�ʼ�4��5�M��?���-�,L���x��'��3O�� 'V�	�H��a��0�$�C�d٨?W1O��O��$ΖA�V0@wɜ�aS&t���-&�D�O$a3�e�p��?�K>Yg�7I<���#B�<}n�ʡ�����71O����O���<��_�:3��r��5�\�P��J��p��x��'ҙ|�R�H��J�<`�x����-H�!zV�� Vb����͟���Wy§�H��	��,��(["O"2�R�+��H�	C��qy"/��~�JT4���i��=�TK�����d�OV�d�O�˓,4&٘D��T�¸=逋�W�:I
$"��N�"�'��'��	�"ݰ���S�r��yB��e$v�����O��$�O2˓Fk�	�#����'���뗯w��@���bG*��'�剾�#<���|��H,���c��[ )�N��my��؋iݢ6m�|J���� U��ا$���8-Iԡ[�.�v����O�ʓ"w�)Fx��t���Z�x=��C�ul��Dؗ�?1�(�08�F�' �'��n'��O$q�h�%$��!RI�*?B���
�O�)1��)§�?��Jܜ
��}�T� ?� �H4����'�B�'j�C �5�$�O��p�x�.<W�t�0��zA��c���(�5�2�	�����ß *�ى��)X��	M�E��HП����`�ڼ�L<1��?yN>9ѥH$o��Sx�e���Z	C��*O6�2���Or���O�f�DxdH����  J�Hk�@�� �#��'���'g�'��	�|Z����+ʏSD컃(ɈZA^]h�h%���������'׾����g�o
� 4�&�!�Y�������$���'�� ��'h�C!��&�$f��p#,O���O����<��R(5a�Oyp�ȥ�_l 4�9և:�P�!��'��|�W�tC�`>�	�F����f��f������*�����OR���<����4�O��O��| �*U���V��!t�PX���|BV���� �S*�AR�ׅ�
=��
c-�T�ε�	vy� �2qT7m�|R���ʕZ�����2��0��G;(M3��Oh�q~*5Dx���ڧ�~U�C�E�Hu�j#���?�N&aW���'l��'����*���LT�q#���@��d۲��m,|�ɁP&H#<E�$�'�hI���K;G�����Fϭ:�d\X��v�V�d�O��d�I�@��>���y�'V0��1�!i�W<v�r�'��'�6��y"�'�"�'a�ܻp�[�!��pg��D��Kr�'�"�
�pc����g��17d���p���aehQ����F�*u�'q%ُy��'3��'��� 2��e�V���g~$2�j�P.����]����?����?q.O�ʓ�Ɛ�4(˸[�t�c��!-
,�룭a��?)��?�-O�͘�R�?i"7�
�w�ј�o]X܀x�e�<Q���?q���d�<��Y_���`��P����t���T��Wy��'O��'^�	�B
1RO|��M�F( D���:�x1I�M���?i�������O_rqOJP���Qz��G#	�myf�H��'7��'5�0�,�L|���z�/�i6p݀�n1_� ��B������:#��S?"�.�i�+ξ|Ͱ@ۥjGB���Ĳ<��ǩCJ��T>����?=I*O��īӽED�st$�KP���'��	�q;�#<�}*��Ѝ5���ӥ�S��}�D��0�rD�M���?��"��x�'(>|�r�� R)�ǂR�I���P�'�4TH�����PP�ʋ.'�E�	Љ`��Pdȁ��M���?!��
����xb�'�";O~0�D�0�P5)���-T�D��c�d��^1OV�D�O$�����(����af(��@Խvr���O�i9��z�ޟ`�	�ɞ},��ADE+R�$�C�� ��'�0��y��'���'��	"_��9�f /,0P��FN��:���9ԃ�1�ē�?������DԀ1	��bA�߈$x��r��y��}���O����O�˓��Lz��OԞX!� �6��U�(!�64�+O���OĒO��8��'�Pr���bVܼe��#O���'O��'oV���4ḿ�ħJ�<�hA
+.Z�l��E��&rb�2���?�K>9+Oq����Tg4By���P6C\� �CS?���'+"T�耇k7�ħ�?��'
�BA���j2��C�2���HJ>�)O$�cf�?ݹ�i��~G�hJ�L�+�Yr�(�O�ʓC1���R�i��S۟��%��$C��:Pr�N!\��aJ�?�X���`$�Sܧt?:���IE�^ ��d[�e�4����6N8�ݴ�?!��?Q�'��'���Ԩ8�,��C�X8\t�&�'��	���O>e�	b�? �-9u	��~S���Fˣ.\3�xӲ�D�OL�d�)+.'��������J/��x�� f9L�Cu蛘v/ހ�?)7)�B��?���?�Ѭ+_9��NE�@�iWg�6�?��2�^�7�x��'�2�|�K����]q�GԽ���d[�^��	�Wtb�\�	�p�	Pyǃ�I
����,�;s���bݿxP���$�+�d�O��D<�D�<Ydʌ���	�%I�\�,���$f#$��<	��?����� �`�H���z�$�F�CY>Ԛ6J��a���?���䓚�D�!U�����QQ �!O����b�x��ɟ(�	ڟ��'�(�G!�ɕr\KP�E21�胨G4(���O�O*�F�j��=yP\	&���*  [Ov1 �F؟��I��'�iW,"��O�����Z����wEɩ
�0�{P��-cn���<����?)�o�f��O�)��3�L��`��f�R��w��c�p��<qv"�*כ�_>����?A�.O��U�Ɓ ��5���i[� b�'�r�'jದ�D����D`ޱ����0ixxJ�R5s�FL P��O�BD]����ȟ�	�?A�L<)��*�0�rqD�3O.�B�m�7��)��A2��Ϙ'��'��l��rA�N�/:h�Q�b�J�nZ��Iϟ`��A��ē�?����?���Jh�11FlB:�2�y�։��'_D�
�y��'C��'�>�/B���a�~�hR���?��7Y�� ����O����<�wfD��v��ajR� �Vȹ �L�����:�1O��d�OX�Ģ<) ��:�!��l��?biX��4�d�����OƓO�ʓQ���+@�z�B!��Q��$p2�5�Rb�0�I����I@yR�ѝY���i�%�F���Fčz�t��3�^����ڟ���T�ڟ��I�N�l�ɳ|bF�y)�1r� �P��iȊQ�'�"�'R]��#!����'<m�$zP�Y7)�й`	ط���I��?�I>A���?����?��O��׌�4hE����OξL��9*Yᛶ�'�_���P�_��ħ�?	��n<Uy4�lB�Z��ͅH��#I>Q��?�EV�?�N>�'`�И[R�W�lDW��we����yy�ND�d��7��|"����^���%�Y�q�Z�Ï�3��k�n�O����O�j�6O2�O�c>MY�l�"\���u�H[���O4-�������	ß����?q)�}r*_Rb �0�%��oF�:2OHir���y2�|2�	�Oj��r)ͣ�&����� ��Y��ݦ���ğ �	�]��K<y���?��'<�"g#�<h��5(��ԙi0�=q����s��(qK~���?i��r#�jb�9mp�+� ��<��8��?qъG�.�O���)��]�!��=v��&p�� �e_"w��&@�80K>����?q����_j�a�,#t���p#jpY�P�q��V쓓?�H>���?�S��mGAL��(�Q ��>L	�����'�I��|���H�'������|x���Hx��k٭ ���q!Q�(�����'�,����0!���ğx��H�e��eX�i26�� �J�vy��'�"�'��I�|�xK|��(P�0|�Y�D.O!P"@��aZ�?�����?	��<\:�
���Tht��w�7T�xĩ���	m��'�X��ӭ���'�?Q�'2����t/6 $x|#�8���@N>���?)���?J>�����x�	���X9�O��I��Hy�i��S�:6�|���
�Q��c%L
?x{0��=#������O���O�ɓ*�O��Oq��@��l�� 0rt&�9"u����'�\�b�Ng�^���O��$��$�$�d�	2{�P$P���S,|��8�	�X
�	�@���?Y�߮c1Z �qo
x��������F�'=2�' �"M1�$�O��Dx��R��G:=��s�� �2u��Ot�OL��Q�:���O|���O|�*��7�.��f�S�D��v�O��dŭ`F1�>Q���:l��D',Ff�u�#��L���*O��Q1*�O��?q��?i(O�Yh�@K<)-h���u���tD�'�,�I���&�(�	���p�+�5Y���#jňw�)��� �.hrX��H�	<\���F��hP�x!�B8-'�U`�ďg���#۔{3�˒l��k����Tm�5ߌ1���?A��?K>����?IB��"d�ld����PR�)6#�?���?���~�ѳN���)��H���?S��"B䱛��"{�j�"�Ā�$�	y�I�D�0�ѥT�>��
6{=�:&i
�2���yD/�UŬ�ic#�!]p�[�H�\��KF�V�k*��@ ���,`H��DN&��8���).)�e�����p�&�پ>[FQ1 (�)~Fq����#p5�dK��H�� PHצb���20�R�Z�<�+ ��\=����55O�U	�N��|}Zia�Nس^�v�� $��� b�BR:%Y6
�]����S-ϖ�d$P�k��Z����BgN�sx�hUG�j� div���Z<̝R�(^C @���ǒf{RP�u�'��'���!�0hD��+�i�dqW�Ֆ� �g@I�8�� ��!��A�'Q%hQ�H�B�E���aS�:5�2�x�޾-Z�� ���X���ʎ(���ȇ'\_e�-AB�L\�]e��D�\�Ot�y�Sl ?�
l�a���|L��'6ԺS�^�=�hDZ�����h;N��D{�O�6�'S��@���Oظ�� b�����'����eļ>�����	Ќ$&���O,7� �i�A, ��NѐS�΄a��U�(�29�� 1�*X��$�yU�ۡ,�8�
%����|�1�H� ��T��#��M92�ln��*A|	+���C
�4Q$`��uc�%���)5Xq�k̊�(βq!5�2}K��[R���9_��Y6�?���i�6��O�#~nZ�j0B���kYפ�
Ч�h���I͟���	2��8�GE9^�L��
�$�h����7�HOr�RA�l�
y�A�H��	�0�[��]� ��ϟ��f:TM"��՟��	������u��'h��H�eFJ䑷FKH��Sc��)	��5cʖyf���T�+s�,���|t:�#ʿ��lȊ� q�U/~�0j#�i�(�aJ�g����ie��9 jX��I�4Hqތ[H>9�
�
E����+W�s5��Ы	y}���?�P�'����d.�1�ۍl��p��'�6"N}�$�0��#O&��5_#)Fz�O��'``T�����wPX�)�/�}鬤���*r��Yw�'�r�'<����wYB�'��6D#&�yV�� 
�0��g�
i-�4YӭV�i�q�ӈN�n�fH8�%����*��䑵 r���.=&��!0��+{8����>*%�ݱ`b����� ߆|��P҉��%�B��$2F&�!\�:����ݤjQ2�*,���O��<��|:���X����&�0^�p�r.�R�<�P��3�МAS�N�]��<�d�y?�r�iD�[�;k��Ms��?������n�"�����Ƀ'�٨�C��u����I韼��	YP�[�-�3{\ ˦�Md
A�e�?A� p�̈́+,��ݨ���9� �Ҡ�-ʓ.���R���RI����?���C�����@��C�B���6��4H؀N6ʓ�d��ɟ�(�X�  N
.�8��͎G(�#"O~T
��I/L^�A�r�
��>a��4�Z��O���-bF}�"���	q��g�O�D�� Ԧ��I���O�J` S�'��iBj\@ d��� 1G�a#��3��9�|�?	�N2#AR��f�>�+��S����唊�O?7O�;�|���A�#EL�W�Ɗce�G���?�b�|���i���s*��^�ZX{af_	 pشQ
�'��9
�!]�2Ũm�5�Խ{'��*��R���IB� <���E�|��dX���d3$T�	ş�7��/��i����l�	˟PZw��A���g��;��ip�燢IK(Ye�R�EPȸ�h�C]�����E� ��z��'�@p@�ǖ}8bd�vDF�e8	��0���&!���?�p�+��?^��:�e$��R�H�jX*��R-RI,I�pO�(<����&�b���E��Pk䙫IN��#4�F�-�֙�I.�,m��	*,�q�k�-4^�� )
�X`W�i>=$�����O��"�# �_��+U�M�/?^��7������	��	�FY"��	̟��'P��hd��kt�\�2 ��@�T� ��B��rsą����"�8?����b4�B�s��� fz��*F+7*dSv�^�����'Xϊ���B�S2��A''ʓpr���)Yτ����gX�E�' �[�<pK"O�ȃ��I�!#j��6�^x$�%�'_���a�ɤBǦ��� \�ણ������4��'�:M��i("�'G��(�@���@*5��i�A����I�:�?���?�$�3z���#M�w�}���ٖr�"#��B��"PrWV�$¼e���c�̭Eyb(с7���
4R5�p��^T�(��Z ��Z'�P��يр�2WfIEy��?15�4*�trs�Ƣ~8���d��i�nB�%9�)Kg�^$Pf����^�'�ў�S��k\�A�P(��7I� ��~�<���C��թش�?�����ik0���On7�[�$�I R#]�N%c��/C���'�Oß0�<���'��%
t �<�0�"7*ď=^81��4g��TFx���i�
�!�ԈP���Z3<���ڴ|&Ā����S��M�2i�
E�<K�-��v��%;��L�<9g�3b&p�
b(U�[���ڤ� K�'��#=�On��v.��8�`�j2/P?�v�����OL����P�n S��O��$�O�d������!	5���{��aBQ�^=0�h�f��yf��	Ԩ'.���2f��^>�'t���]���2Sx�1���)+*�i�/�l+0I�ax��BDqӸ`�	����̷*�bN>���M %��:tIp�I�eܽ=O�5�	&��� �M���~�'�RQ��)�8od���_%V���x�",�m�����)���;i�Y�E�HE������I�?�	`y��҂od1a��@����
½��pA��T���'���'��a�'��8��d�,�e�,aQc	Ɩp#R8;���Qd �a��ڏ�l	�	))�0�!�(O\�q���4����b��UM����i�#?:�ٳ�H8O��X�aC�s�<������(O����'���XR��h�N�p�͕�<�|�E�f�<I�D�T�}jԢ��r�8ɉ�m�L8�XGz�!G2I:��!�K2�:1�B
M��~"hӼ�OhdHOЦQ����O��0(��x \�4g��BT���B�� �"�'"�ͤ:I$�8a��3�\��L1!$�HeON�? 8YGC�;n�ʕ٠b��/�$}HD>�w.<�X���3V�.����$� �ʦQ�4+��>�^)�a#�n�>��n�n�'�.��g�Q>Yh��\�V�>�KI�*py{��+D��Z� پv����%�D�k% �ס$}��i>��N�Pc�JC%0̝bA�wP��F���Z�E���M+���?Y/���A�OR��u�|�Xd�]�#*AA���_�hQ�·fi;��=�R����G�� q��Q4E� �|��-J�Z`�S'�$#�͝
��o�8`gD|�a��tTzqBgN�D~��F�'hq�kL>qJ���M�(l����-�Λ��N��?��|���i�i���P���4�Ɇi�.� �'b�̰�
:���iҔc�U;�{R�'T"=�'�M㒅��6��q
�:5*t����..M��'74�Y3	�!8Y2�'�r�'/(֝ԟ��H3�ȓ����/�t�E=\A�|��!XN|���Ϋ ]�n�~�"͚/P0�Op	��1Z�x,'l�<��[�!`���V'G:A�&F�o u8���{�'H�Y�D1�O���C慙>/��5�@�.6����T��>���ğ� �+��{����NTx$�Љd`V!���MS��-��I���\/�A�G2u_�#=ͧ���t����K*��r��;5�\"�+�I>����?1��?qԣ��?�����φu=ʅ�7�3Dj\l�ę{� ɴg�*��=�ߴ}�X�z茏�$����"i1x���H��� �`D�H����$�K����j�F��%����$[)܈��%�ȓO̈��'J�)Y�&�7s"���"#�ƁH��n�<	q��7�ꁊ��J�h ]��*�q8�XFz �
 ��M80�Dg@|U
���~ҁ}�J�O�a1E�@������,�OKVdA��4nX��CD>� 8��RY�����O����d'�'��?���F�O�ӠG#��F�K<�F�e ޾i"=���ݺ����#��^�>QZIүd��Sb
C6j��aq��߶6k���J�<�T�N��(c���[1y���q��Ma0��4�V�|!�3C��Y��@9�EUj	�I�|�+}K	PP���mTX��u�T��"�~�@ey��'��V>]������$��ʦ��C)A+b\JA�S��jMkeX	0��|#G��"q��@�iۼ.>bE�_?�$?���rw�dc	�l9�}˖@��Ѫ�n0N���0K�K�Ȝ�7%.l��G�\c��9��핦��q��,�H���1شg\�Y�I)�M��iVb�sӶ�J%݊e�<p�4KE"*أ�O�ĵ<��"0+��%Ʉ��dɺe.��Fz�i�J6�.����"�]4�$m(��:W*�l�t�_tE���?��M��2$�����?)��?	d��h�dt�̙�Rۤ�fH� ���!w,��A̘�gX�Q�	�e(qE�3"��S�'-�p�埖<�P#t�X8A�\hb֠�N)<�ae 5tP%)H;���#ʓB�Ҽѧn�i�j�_X�a�'|�M�����z�8s�\�0� �*�����Y�yύw�X���41���[Č�6�!Gz�OL�'~`}S&��;0*v2��6	,jt�uh�8���!��'��'�bb�0 ��'�N#8Bv�))������6�,]�g�\1t	12��!i�ɠJ?�P��q�ġ`���E��#��ЄR�]��ܡA�
e���Hq��3��Ox�j2�'Q��QB���C�-��?�T�x�XD�<9Ƙ.�tX�7�ۀZ�U᪛z�<y�(��C�4lY��:P�6]K�{?�P�i��'Wp [4�|�.���O6�'2�B����%W%�A{#F]/0� `#��Z7;���'R��-.�Ų��-}@J�z"��3
���S�]�rLX��EK� \Je��[x�#=�q*ڷlUf�p� B�T~n��w��5��TdJڤ�  @&3%�P9����HO2�*r�'�D�|��M�)���(�j��1fz�K�Mi�<�C3,F�E#4�H?��!I�JA}8��I��R��	Pk��̊"d�श��!@���M{���?�*�����O�dd��i
��\�lV6i"C�N#ezd��D�"#�u�VB޻ tj��*O��f��u�tE7U�, ��;j���z�!m� ��T-~�H�Yo���3.Ɠ_�B�1��\c�1!de�#&d��H��tP��ݴ%����I���S��M�%!�8�����a�&$c6Mw�<y�/߀�V��J�I)�\��t�'Ep#=�'�M�s��i@�P�%D:h���a��Q�9���'T��Ǡ�K��' B�'���П�.?��8w�B�ufr\q��p�Q��fh6dT�_�1��X?�B���:�'�`�I�9
���=׮P�eCʚ2b��g`�91����2ǘ��i
�3�5�O>I��
�X^�'��{�-Qhs}�g�<�?�T�' �5��ؠ�l�*T0r���'M���fo�[�����у��&3�"=�'��9Ub̨v��tXA��� F��\Ä刭0|�`��?���?���?����?ɴaE6zV � �C?.fB�'�[6��A"�'��9�����I)R�X��3�	�M$��v�t��  ��#�V

r�`C�X�@aM�&*1�!1@L.��O�yd�'���D�8PtYRE��Wz&���U�uO$<'�P��� �?!��M$ �3�Pm���T>�h��Z5A��'�L�����|A� z����T��'�f6-�要�'b�1 �Of���D�O��'zK�y�Fˇ
X�E�ńO<�j��w�1o�r�',bN�0L�,�n��$�5�τe�'"�X����4�U��q�Fzb��J���!��Ǚ-�vp��å?���i��d�%H��䡓G�mA��p+��O�`G��'_�`��%! @�4�Hq�L��yBDP$j]zBf��&�NSPn,�p>���>�Ъ�LC�a�A�Ɇ!=R@�b_~?	���>L�v�'�B[>a��͟0�I�Ҵ�� W�Z ;���s�Y�)��2kA�%��"W��%C޺���4�s�Փ�KغΊLz���8"Ӿ�`�x���:4�Y�Y�2Ѳ��T�|~�
4�:��s⇰W�Z�Z�a�5W� �@��[��0�*�O�c�"~nڥE$�kT�" ]��ɧBĸ$�ZC�	<wT��3+ؿH>���f�p&"�<���i>�l��`��@S�[�o].ݣ	^G�4	h��?��O
�8�Tuy���?Q���?i^CY��w~��@�F��H�R�E�ypa����!H�>,���0� ���Iʔq6$ݨN>Y��1��qjOX�lJ&ǚ
ap�K�\'����׵@n�O����
$m�F�_P�	o��Gv���s
�$e�Lx�'�<��H��z�Ɩ3(x!��f�.{�Z�Qd��7�y��ۧ2���H5n��P��B��B�Ez�O��'�4�E�S�!�Z����ߒ�#��e���WBƑ�?���?��� Q�����?Q�O"T+��k�4����I����A�:c�0�;�(S�0� �o��2~�,����`�'�0�H�d�p�pR�D(N�jY�v��
?���1�I��r&�ۘW��)Q��BV�'�$d1�9�d;1�K���i�$l��g�,���A4D��CuhW�d�9��W +�2��3D��hq��l�8��&�bn48Jb�����4��
�A�_?%��T���->ð%�
��ΐ؂o�6xv8q��O����O�Ep�	$��9�Ç+��6�Q'2<q�DS�|��}#�K
�".h���BϠ E�<�bsABmҿq�f�q���=�GbE�^���xBΛr�´R���/ �v��cǑ'Lb���q�O�ln���O�^�H�;S��d�ټtt��'DR�'���ss��J�����ꂂ����t��|��E�2��z���*B����Yo��e�iQ��'�哄Q��A�	Οln�5�VQ2���9L3*�`�jC,�Y�ю>A��W���� ���(!ϊՓtP�̘�56�N>F���P/��@K��Ƚ�M��D;~2"��棚�XE�����V NNN�㛡hj��5�%�);pt���W2]0ݐ�.�M�peϟAN>E��4c��p��f����s�/ށ0v"݆���dp1"��+�*��7��(6�LDy"�6��|��4fX���F
��,�֪A>"!��c��'v2�O���'l��'�B�aݭ����qI�JB��uĴ���]�)�d��� \]iD�ћ��So�����|"��%��Pc�)3|��7��$e�0��!-ĿQ� 9+#�@�a��#��&�jG���qc�q���g��dj�,��!�'�l<��;z�z⣌"��I�$��B�g�م�M��ZV��]i�[� �"a)��ހ3R"=�'��.R��v-�~��!1u$7<���˸F�jA���?����?�2�?��	�|ZЂ�3�-�g(��>��Sg��|	ƅ�9��O�$S�ڭXen�
T34�<Q�N&'���H�d�$(�J�L����/�<M �M&ˎX���H�o�T�<��O�̟�3��# ���Mغe���3�ω���ش�?9/O�D*��|�Pl�;~ID!S�d�I�s�<���+3���2�E<9;8���Ho?� �i_"T���L�����O�&1��W�D��w�J]��Xh�%ߵ���'�,F�7*�:�K[	$9n(��E�d���a�.z���8�m��*�X��E�v<��ӌ��'t�b(9t��>
�`�c8OY�I�_I������Cd��օ�1<h���6ʓ+�n��	2�M���i� )h�E��2�>��r@�|���OT����5]��y����;�m����铠hO�s�ę���Eƒ�`��lJV�Zb{��̝I���nZ䟸�	X��X�>�2�'"���F� �t���ƝP�Ak�D��~�Hhp��k
�\���� [s��o9��@M���ʗ�m� ���+�=+�T���Kp��;{���"�T�4����-H�'C&}>Α��5�y�&	6T���FI�=�b��üi�d%���bɧ���Ƈ	>�>�2�%�9N��bϛ��yZH0���s�:yH�_A<�Z�{��'�"=ͧ�M��7L^aiת���({iъ��nZ۟dC'ʁ��VY������I�Xw���~�yā�eM��q�ު\�����<�"���=��U�牸'B�S�ûQ@.�����	u�a����d���D���"�{����a�S�? `�i�.Мg��9;f�U���q�!T�0k���On�l����?A������}�P͖�8F �F��?\!�D{�A��S�J2��4*D�y���4D����|BU>��'vHW��ub���^�`B4hc4�'L�s7�'%��'��^/uh��'j�)�<1��ESf@� >#Nq�E��|tq�@�$"�:L��={��,!ǓF�P���B	S�~��s
[X�-P�f\>D��4�WoεO��f5O:��'(����K�z1#��J�<������3�y"�C
O��	��$��"�8B2hɿ�y2O߂m��p����u��ȲK���~�':���8���4�?y�����X�,�D%��.%����ńEGC�5��T��t��ğ�H�bV)z�]��A����qCL�W��y �m�riS
d���+�#.l%�<���Mc�!���_V���R��U6Z%����Q<��p�&ϙJg�p�"Rģ<)�@\ٟ���4S��O㛶�
"V����D�;6?@#1�E�w���(�)��@��߇$I��pG�I�<�&�4A<}��i>RJ��P#?ɴuq�fE9����.���k����M����?�)��h��#�O��$o�t���t�4�S\�R���\j:rd:A�j��eӲ��0�d�����.���F�?�s�E�`X+t�i3����)?���"�jӚ�
f�,Z���G�$i{�����+aL��\ㅂ+;֞�)dd$96������MK%��ҟRH>E�ܴl�4H �b�N����KI58@���)����L>kh�U�C�@/�$Y�=��m���S���rG̃>+Ĉ\���ŨuH9�	���?���p���
��?!��?���t��O'aй��ay�D%CȰ��¡� 82�	�2/�gC��3�yp����>��R:��F���X�bխ_�*�z�A�&N90��7Ζ���5�i|����K�����i�*lK�y�gC#�%�V�ڝw��3��P[}үɶ�?)W�'p�[qZ��:�BCNo���
�'>�f��)VB�aCs���u��L@''�)%FddEz�O��'��us�+M�@��"��m�U���P�����'���'�R��M���'��IJ�f!\-Ѥi�>��� W�F�d7���R�,i� �A`W����̰o%�iЊ�dW�,���M�}�p	tgy��aD�).���[���"zJF���k��+Fj!�qo�a�'�Nz��KF$�2̌7?'�y�mBtX��L,D�X��F�8�5�6*�R����)O#=a�D�=0��&J��_l�d�L?y��i��'�� 0RMw�R���O��'''�A����!��U�G�w�0�q�I��922�'�"���D��!��!䛶�$%������ݲRe|Q���E�+�x;���8F�:��	=g�Q�֎K�k6��M��iFtsP&%o����b��1�~mpQ*L�� �ґ|"��?��S�T�d�s�(���+���*%�B䉆vgz���%�B̀	c�.��x��'�ў��<��	�n	����N�f��X����Z��v�XT�ܴ�?����	�N�D�Oz7��N~�Q9�*aD���l: �<�sfA��	���E���2t"�M� ���Q�՘�5��J�Gw�D�W��옓Յ��MrC��n$��BބC�h� c!E	:�&��������S!LDd�E��%;����i�u����?����?i���i�K�$V�7�t��ŧ_����'�B�'�YС�/-~I�#,Z��Ӌ�D�A���D�i3��
R�B)y�lYtK�	�p|�2c�OH�D�4/��Hr)�O����O�d^Ѻ����Mk�&�%P�B1�G肻p:P}��S}bn&�>��+ː_��*���j{�\��dX}B�Y��>��l���z��󣇻C�QrGV}�K���?i��'L`�cH�Z�}�,EO�\M�	�'Q x�4FE⍺5NנP���A�$ʻ�HO>i���E�o��s&ܮ�Z�+�ݐ/����P�����L�	�s4�����,�'�q���QQsg�A�V�(�����7�O��B3_�D����
Jtas!�}"`���.*�OJ�`s�'X�QS�I�V^�<B�U�/�B���ZN�<���% ���)g�9���HQ͉o�<�`��s�f�ԅJPK$�P�k?���$�!L�^4m�ן�IZ���VEH$�D��%|�i���[�Ph44��O���O�Q��@C�'hI��%\����b�g	ܐ���r<ؒ�#_�59�,�"�#Q�Q�<�6?R�x��!Oz�!��:fǸh�cm�7(��R���(c��K��ά�Q�Ē�k�O��n��M�����Ǣ~g��P��E�g��t)��B�z`��E��?���?�+Ow�مtk<�"5L�ݜ�+5	;��	q����|�P\o��=���0Lٶ�2�\����$��@�	{�d���%�P��-ȱ'N��3b!^9�0)��h;D����O�\p�H� 9��U�����C�A��1�G�+�D�Wk*�!�p3��)��J�L�8"ȇ�S�? ��`�N8}n�P{�i�+� ��`"O�CG%"TP)XA��}80T�"Oޅ"Ə]8|z�H��',g..� t"OV!�`G\901yp���5h>���a"O��@�l����g��B��!"O0e�[�H���BAG7����"O������XF�k��ӆP0"O\$fߨmfh�"�n�!CQ��y�"OU9�iЫ/���Df[*S�z�{e"O��Bp��f���Y�ˎ���ؖ"ON��e@0��h�rH�63����W"Ot��)�f��Q(X�8݈U�"O]fOT1c�N�j�a�g�,Y��"O��
�D�6.�$�1tOG��
�"O
��T	S�(�h��; !p"O�c�k�i?XXs�ğ,X=�\c""O\%�cA:��k��M��J�"O<�/�TK`A�jt�!jT��yB�	=U�$IbϏ��~�����9�y2�=>���! ��2�Wk���yR��R��H(����z_65��jB��y��Bn���!�/i@<�"�C+�y�%J�Ma`)���\�ain5���ڹ�y���\p�M:�*:�����ybCk:L�9E���pA��!i���y��˺?�E��>jvh	p�'�y��Y!ɸ����I�`�������y"����K�FR���桒��yBHH���\�ѬE�vD4��#ܰ�y�]$AH%� �>k�ԍ��)%�yr��+H���h��݋g�:`�G��yB� �NMI��Rm�� ��
%�yB/�3�:0����A�.E�C��y%N���I���T'Vzh���X��yB�܋Z(Ș8R�LY�ii�Z�y*ޕ$Xz�� +O�G�X�Y���:�yb�%(�4Q�2'�~�g��y�A�z�ۣ�֫zt����'�yR+�l��M{���+5�D5�y!&T8�(���.����W�L��y2°Lt`�h�jޓpܰ ���q�<i���9Al�# �t��3��o�<a���V��@�� �@tӣ,Zs�<�#�P
rΎ��tG�?��,G�b�<�T�O�	���B��"i��y�"O(���%͒�n���G5��9�r"O��fK�7��1��><�F��"O�����׬)"Y�TA��Pb"O�tQ'l�;%-V����~XH��"Omre��i���sC�:6�V�p�"O�x�#h�_�H`�����.�P8jU"O�"榋��0*P���{���y�"O��Zfm�,u�6���!�8�.XH�"Op�!C9i@���eO�,Vz��x�R�L��7�Ol�A�
(�ν)���y{��3��'��������q�#0>���/` ��!<D��H�=y'�L���U�V�Yj��=K�>�S�`o�O;"=8��S>;� R��%m(�j�'����I�2
rj�@/�5�K���f0��y��9O*��� �5���nU�!)j-�G"O�Y1G!�mC�<B�V}^i�B4O6���$�!'�a|
��t��,0��5^��E���N��0>a��R�qj�̓b}�QZ���G�j���MЕ�~E��.�ty��52|}
�H˚-p�UDy"��-�p�~� ��0�@T�P�Z�)��4;XP�$"O�����_�U�N� ���>�����i�x�c���s�6�Pa	Ǽ#GNz���5eK���Q"O^����L�`����w�Vͩ�"O��S �v�x�(Y�v	0"O$Q��g��kRh$�(���ٳ"Oȁ˕#Ω9����6AZPy@"O�����H�Z!,�k�g�ZUZ�ِ"O䊖�l��l��'/N�`"O�9Ke��3 ���KȐ<Ff�h�"Ohvj��{��A)֡088�"Oj�%C2>�<h��H;v�����"O1r�SU��af+_�&��(�"O|��&#�Y�ڍZ��Ҫ�%�S��y�J�/��l8��]6�ܕ��/���y���=�)A��� N���]�y�M�EW����ڋ}�^ +@GK��y�)� k���1`� m�ji2��ت�y�%����3u��mІ��@���y�%�<�^�a͒g�����y���n2��#e�U�\��f�Ԗ�yB��q����`�g�n�
�e�
�yr�9
~�E��\z���⁬�yR�	�L���w�T��P"c���y� �
v�B�� )P�u���+��	�y�Ȁg�9��*�p�Qe��y�f�f꾵�P�RV�2#
p���_��xD��9G��2J��g�t�ȓ��-8�M��z����R=kR�M�ȓkڥS`lQ!Pr�Ү͹o�����0b�r 8F����4g�2L/�]��!|��������5%�RB䉿O���ꑇ���0x5��.��C�ɕW�r�Kf,�v{$����(�B�oI�UⰥ�X�4��M~K�B�I����E�&2P�$�R��B��5.*�Hh��T$h��ĤD�B�ɷ8�n��q�E�7��IYpaTL�B�I7�!CۻCg�͸�)�1��B��4h��Ա4�D*����Ĝ51*\B�I�,�d���l���X�bB䉆J��e��֢<)��Y`��V�2C�I!�r�[�Ǌ/V��x���(D{�B�	6?����@�,�p�� IJ�O�C䉀u܉Z�ER�R�.�`���4��B�=�JY���O7u�p@��b�P��C�ɫ9U�xA�$P2Z|LS��ܓhRbC�o��uxץ�$:u�F`�b C�8*B��##܇6���0t�	OmJC�I;|E��)f���4���1��:$mB�	��u��%��>�Apb���$*B��
N�*Dy�2wc�eH0�O�B�51� ���4��}�d���B�I�J����8	�N"�T�M��B�	�� bj؁jZ�YB�S�"�B�I.*���i�''ܬz'"�	�C�	ؒE��8��irc�q-J\��"OH��VeC6<�=�f+�8Olz$"O.h��ûP�p���G.< b��B"O�a��<�Ȃ���1�΍��"OB�Ñ�
��Hu�U�x哂"O�K���5lʥ�ƅ�!�D��'�Ը9��ZW̓64,UP���:��}�g�D_���ȓ.@��CB�6i���ȣM^>T��'ڠ��SBO�x/�T�OQ>� x���ᔥR�	�5�vN0���"O�|r�Ŕ[�n� �=\+F��f�I��򄂘^�z�01Û\�3��1�HR���>s��aD���EȠ��D��)3δ3���s���"T�`�\��ׄÌ+�B�1qN?�0?a�Aº?'t�y�$/Yꦄ���y�'"��Bƞ3E����x��J�:rk�!���� &ZPZ'c�0�yb�:x�ݙu��0c��kWj.�y���[ X,���K�r����r�S�v�V�J�_5�)Q!X/QLNB�	�}�Hd���+p��-�Kt�7��\�R��3~�TL�d6Fx�+܅M>T����4\R�(����0?�q�X�8Xʶ#o���Y5!�lբd�#\+j6�I��˚��>qeJZ�u��<)��Bi�QYǅe�'�J]s2�!�Ne�`��+��9�4�(W�
p�l3��
 -�B䉽 �+��R�	犅�c�݉���?#�"e���>]Ƚ �
}�OX<q�b��+B@~�aF�X��yRV�T,j���8`ѨC�-ޏ3Ml�Q��'�f�3���Q���p˟�,Hv`"6:�9 $�On�襣6�OT���A0!�����������>X�V���m�*ȄD�``*�O��%&V(@	g�ěO�����!9\>�!��t�@�ᴛ?�8����,�X)e"�4�'�-D��I$��O5�i�g�V E��[�+��x���>(�4*Ф2]@a�tO�)�T,[7fݽH��
��
,�y�#P�59�`hS�1z�T�SL &8�'��]X��2����O��F_�P-,$BN an(�:�'�
��FO��6�Y4�J��ڑ���G5��x�@/�^؟���d��*����A�O� J�$�#O���G��'�"��S�V4.�@���c�{iDl��'Fh�b�<zv�Ab��)9�L1�',�t�F�_5Ѭy�a��;�d���'��At�D�TDQ��6j�e �'�. @b  Y(����l��R> ���'��j�OK�r��w�ÉKJ���'�a`��hz�{ �ɫEz4��'c@���	w��H2k�
=�T�j�'���b��4���B��V(�|�<�`��O����"�iЮ�Q{�<���܀Sg4�cf�:@�� Fep�<��%*NX �BM/=>��a�
�m�<I���l��@��ȃPB4;���l�<)t��3<fq��n�m������Q�<��Z>9#��cA���x.�L��j�z�<�uD� B��@�#��6|a�O�n�<	�cO�BV64�ĬC2��`�S��e�<�t�<��<5�˩z��͑b
c�<��@
J�^�(�A�b;<�U��K�<�G��1z��r��]�i�d�Q�E�<�.Yb��Q���%]�4ek��e�<�6L'WG48�s��tt(�P��c�<��=�`p2AN�4P�!��R�<�k[O��}% 18\��y4��I�<a�cÌR"b@C��-2��Q�f�H�<Q�+B�_����Xzz��AFL�<Q-`�l@Z�O56:���sHE�<�OTx��5�pm��2h& ��I�<!���x�D�d�2���+�n�<Q0�S-�2l1�g}����P&�P�<�&$ȝ 4��pv�������O�<1r�^�����!�R����a�b�<a�`�.sv0��)	=��sR�d�<A2��ofXy�EU���BqN�I�<)��C�u�z	�P�M(�X�R
n�<!���G�$1@
+ijV@Ҁj�<����(q�qa���n��} ��d�<yfB%N�S)ɨ%���r���~�<� Vyye3����ꍙM�D�ؠ"O�A
c�J�@lR�S@	�V����"ODh*�/�2B2zU���*[($x��O�-�!KSG2H�:�!�p-*��g��g�����ېRȤ���VA2�C�	�]:B�G��/�p��ţ��	�dC�	<Rq0�r)��U�T�)���;\�VC��
I�:t�Ǉ�����+�/b^LC�	-)�Rd+�FS�}�H� "��<k�vC䉨J���1��(aJ�;���}:lC�I"���y�%^�d���{@���C䉐=�a3fi�	0J���7���(��B�I] �Uc.Z��5�'��kq�B�ɁR�ޘ�Q�ؤo!�<�S���,��B䉏#o.!Bf��?zɀ	�C�@N|B�ɐ^	^a;�	)�P�s��� F>�B䉷d��0���"� ��J�~hB�əzf��*܅c�� �R阀4]TB�I���HV�Q����$��qFC�	�vR\9�BמY!@�|[BB�I�tv<�`O�Ljv�K���	��C�	 |wb��ӅI�i�"�A"��F�C��3|� ,���]��Q���v&�B䉪�|��7�1fZ��2q��1��B䉜��A�B�#�z�PGcXU5�B�ɵs��y��V�
e�֧7p�B�	D^T��Ԝn\.��b�y��B䉇sy廦fW%xm���蟈lL�B�I	:�ԓ���2J��@2W�S1`�NB��(��3֥=v6jH�O��_�C�I8�*p��B�N��, ���<D����
7J2��dN�{8:BCk'D����$C*6�JŘ���}��̣!@:D��v��=bA�P�gD-J���!G8D�l �ʝS6��f��6a�8y�5D�d@v��T���s�	�e�X�4�]&$���B�e�pg� X�㐥��b>c��z�nȦ7S0��c�9D���{�@�o�mx7S�f�A�c��i �FzZw�k��f�x;�M�c�0Iք��h��kr��_4�:��$�qO�'����>m��rf_%4/��/�6E�������(O�tnOt�	��'�$��� J�Y�ɋ�4`�t��`L=���la4.��$� S�Z�ޤ�g��VⓊ>h��@�\o�LY%�]���3��d�6m�7}Z	��:<o21��)�<\��4��(�&D���V &Zs���уY�+��hF숻+�pa�1�F}"���D��`	�^�L�W�(+B��3�F�N6�a��I�%6���c�Mz|MC�蘉D�6͖�A:~�r�A��)�1����&�Q���Ǝ�!�S�Z䖜��i�;]�����"O�D80_� U��� x3�A`�K^�C��Gy��@����-8��@b�3�8bG�]�0pPM��/U�l��ɵ�'Y@R�clH��B���iFd͂��b�h�<�'�	�u�b��3�݂E)�i�E�'&D�R�#V61�*��'�6�"��� S�z(�#�8-���o�4�	�5X&LXb�ay�AS%���[O��X�mҤe6���'b60��ݎv̎AJ��ˢz3�H"�4fٜ��Ն��u[Pg�9	��mFy��3&�A�2��x1d�P{ܤ�k� {�<�6�^�8�(ҩ�9^Z�Q���.-��D����8�*֡���S���μۣ��3"����V�	��@�BEX���C�J�4}{�� c��y�V� lIJ��
���DJ	��$+5�6jp6�$�H3��"|���F��]���_2D�Q�q̀�m!��i��ɥK:�$A f5_�yD�tU�@8�'��T���b�ӣm�������RyH1�,aV:=ؒ�.}��:�Ͽ�1�N*�4� G�Dk��[3������S�	p)_�v���l����a�໦��4���J(o�P%���gɅP^��'倥���$�v��8)"
]	P�m`��[;��]b�B�s��*&M)��lb��K9{a�n(�r���#_=6.*�ʔ���~I�O2$z �/��?%ۀZ�7�i�]�.!��Em�<c�,��'�B!ృ�9F�X���c�B�)�}ZwL���@�k&���IK [��T��,�p��j����]VL���I�� 6\�'4Mئ�)j��ݪ�Zo��� Hä-�ꐠ�#�M�S�O���A��X���<!$Si/n�jݴzh�I���g��e�$�խ-0Ey��� ll�7C��v-��!1T�v���xS<"(�O����ʲĘ�m�t�`��9e2��B%
�lˌ�Gy��-Ju�d��%���@!:�
��c�Շz��`�VgF%f�R@�D٧;������bhǋrQ�mZ4�58�@�s�
Wy�a�(_T� ���	k����L4���uM�"z�N85��$�V��`�OQ�,�?y��OtB�tbTɊ��F�R}"�\r�*��!��\�F/��2B�pR�-�G*�)Fx�g�F��� �E-�6�(0i�)3�`m�=�@���+Φ]�&�3�k<l��<�s��+*�a4�l�1 �A�&a1�+�dP�LN>��۟�r;��k�ߨ\+�<
����µ!��H�VQ��	ψ��=���[R´ϻ4�0��L�) � T:�J�#%Gx��
U�`�
�d�nL8��$"#�0����d���KvU�88Ĉ��^��dPs'�5�����8�mþ�YU,L�w��pybg��q��`ӊ�DmC��[Q$\�7�q{fo��1q���o�Up����|��2�������L%g|\p��	g��G�T,�5��,�.���:y���l��e:q ��Ʌc�pP#ǎ�V�<�s�U:W��!�\@�E����Ar�� �	W���O�M��&��z׺�f�>`���'�<���:W��n�]����w\@d#Kۿ$F�)�L�T֐Ux���*�G(�!���,�
J'%K�N��x߻V"��3�W��i4�4<oZ�����B�H�V�#ʓ|� B�z3&<C�U�� ʋ�d�|x  
F�#:�&=A�E�M����4���� �%.��zPL��*�ʸI�Q:/�"�S���X�Q���k�I+�Mv�� ��@mZ5�0Ȃfh՟)A��R�E>h"@�<�s��s1FӸ`�*}��!��~���90C(�T���OX�P1o)
��Ԫt+�mbt����(Us��<�	J-�ըp#�--�t�	�w,�\�P��e��=)�Mik�-H�"eZ�'���(	+u,����]�g���Vk%e�H�cgF�<aFJ��L!A��9U�4�r���Ɵb?}$#όF�%���7m�.�R��� ���*e�M�N�\p���'�J�?]��Z�h2nW�C�*�b�BH
��x�t��`vt8��&��&K;O��%?	KM>e+J�Xxxc��E!�i�Ek�
//L��q�
�h$<�� �&��?טw^q��E��lJ�$�A�%׽��m��#�2D�k9�|���ͼk��=5�&uǭ�U�H��7��f���Qg�i�M�"�K7f+l�sg&�yǉƿRV:d��(�#�h�v����'��9DH�1�����)��bI~���:1�,�S̏/#G �"�`�J�'{Ρ���B�OS�)�Q!�m�b���Rب��5�ܸ'TL�D�,OJ �W�>1с��P�R�`��Ov�5����h�� ���&�Ј�1f^�VȌ�10�0 �L�jV�'� Ș���(���W*VD�@��N�I��D�dqO�ذ����;
v�q횹z�����'.���f�R*bf�����[�L���t��]�=��\����Z�PoT��d��1���N�Q��	�NQ%�>�!���;J(���cd��@�EA��=ي� q��<aC� �^�JE��aJS��� �-�v
豣D�/���25��([r��}&���U�I�����i7|�4`��A9u�y��+_�p�cB)��E{R�wv|)j��
!t�rt�������`χ�&��@�$W�~aH�{*�6@3g9�8-I�J#Du����ȗp](�!`�òD)t1Dy�'�����ط0�(�#d3�� SO��W�r\En�!LO�f=�d���	bEq8y�%�%d�N|ZS���č�vAG�4��U���iy2��%])�a�RM�'�(�
��?�~2rƂ�
����-�(DR�XhaZc�,I��i�/l^b�@ ��O�T���ʬ>��B�t͊}jD�ˆ3sP��D��^@(eKӤȇ���՞9�$�%?m:7�>�&L�2�`xQgc��	�2�{,�M[,ojl�24�@�>o� �aN�T����f}鐄�\%�|���޻c��H��hƷN���Q
�j��9��>%?���wZ*�����1���%�T`m������(���O�laf���]�T��Q`ܚQU��X��%Kb5xL�P����%��A���*4f݈�?%>��`��)������vs��ؒ)�<�g��2b����rj[� �<��rB�͟b?y2T�]('�dXc�(��T+ŋ�܄pf�X�uN�@��'Ѽ�?5�R\���	�5{F5��n�|�zl�SJ�Z`Y��iDij��4|���� �K���p*���T�7d�U��Pp����e�Ⱥjw���Ʃ�Y��5c�$��?��� �K�P6Z���)3�E�2G���3��D� d��޹r#X*O<%>c���,D���ɖ�]�n��сM�I=J�2"aϽ,آ<�S/?K~��U�]�	�J�0�w���Y�	��^�z�`��#oGR�ɡb?}b��^��b����-р@X4=������Y�>;��u�X7B�kQ���d�)#]u
��U!6�`-sҠ�.<���D�׺f�¢䝦 
z�`Ã&�x��d.�l��h����<j��$�f}�k�&&;h�zt#K�9�F	8C*3*>m`��֋��5n�A�HDaB��4o#�d�`��#cn�)XIh���F�ā =��,9�ImT���@��(O�\c�:!3G�Z�H�l�?")�ċ#&ˁS2�1q��5O���'~�� R,�ň��r���hV�	\��8�%�"8�Fy��2r�� `F�I܄��O5F}r0�#y( ��k�(�9���T����D:h*<��H|��*���d��ʚ.q��X#/oy�)
+:ĸQ�j��P<����ѫ'\���U&K[P$	$��ş�xv��
Z�D�2	]� ����+9�Ε�ő�:��QU�T�9���W�,?�$�ԉ�yIM~�=a�rPJq¬ǜz���#V��V��	�^�jAłA'��g��v�,x"�)׋l>r� D"],i�8x���*2r��
�d|Ԑ���	�2����A�0Ur���$q 2�� �<�(O�����"z0Tp�����	��d'�ܠ�|��"���� ����<P�������'p�th���.�%:�F$P���'��9���:@�h�,��
�Xp�ˋbQ�<#LQ D4:��	,p<�#�)�	�AB�O?qCpF?1k�@�T�ܤ1���#�D�����O&����L�_����qO�DKp�U�:d�܊RÚ�N�t���SD?!'�N�z�uI�gǦ���$N�(�.m�׋�*|���Iu��@,���2��;=��c�	���<9�iP�M��1Q2��)1�&^5P���(D5ES�����	�:[(3�.N�����i
��], ��t��#hѓ�'�8=1زO��ܫ`�8:4��ND��M�>'�ę ,N{b�7[���o�x��@���ΌS6p���?�'<Ұ�S�%F�y�$g����	�Ye�Pa���.�6�r��O?3Ս��NSz��?]i�e���<U��0�1p���ӑ.K�m��%?��<��c�/?YڼS��ΫPo�C�HZ�/����d�ބy���&�g�I��&�x�$��Rq#�	Y�)0R�gcӉGʒ�i�� 6���+�'���{� ��^��E[3��Z�>噂��/bV�a�#�F�UQ�DZ1��1(>����&��`�'�V$�R�Y�Q�3���14�R�#u,�F}�'�5 �d8G(#c�O�6��A�\"�*2!��-0F�p,O��P��2���Z�� �M�b�#��8�'v"^�`�� �b-��G�-m���'ǰhg�]�h��O�>%���R3،��3��欤��S�>�8�2�ň�y�j]�e�Z�N�0��jb�DjA*	�2	(F�Oha������	�RB�l�E�3?�4  �E(����LD Pb-(�U/�� i�j��jOD-f�¸�˓E�*XKT͒yg��/d�����Y� XHR	5��r5��4�����%�h2����#�5Sk"	9Q'S��4��'fVEt��$&l�8X�A�DW�Ĺ4���"��'E�\;�� Z����&�S
�䭲Ѥ�2-|�T"�I_�d��C��;̤-��׉]�,e�vGK#.���a�D��~b!Ӗ{�p����{b�N1i VPH�j�2:�e��X?��?1e�^)��!K���x�ǚM�,y[ׂ�t`�\�ti9�O`r��-c��q)݀j�(U���'�ni1���iU�AQ��q��Q�AV8c�ܭZ&p����.D�`����_�ݩ�[/rW� D�4i���t�C�f�
'6E��=D�����8-��+whM2x��R�:D�ls奔4|�¸��� wƲ��d�%D�p�w�J&m��Ai>jD�sn!D�h�A��n��Qre�;_d(M�w?D��b�P=+���6$Y=I�����>D�HP2�)UN�+&"��4=D�����G�da��c,q�Nh�Sf9D�<qp�λj�k�ǹ�t���<D�h��K�p�x�#&�J'�K�f D���D-�ps ��C��3�XYb%a>D�L����"x�`�#�K�I����;D�0Ll~@#��ʕՌ(rF�7D���ޤ-dt��A�Lf�,ّA�h�<��]s��V���w$�J�<�F-��Z��LU~�d؀`[E�<���ĝ1~�IB`�,�MW%��<�����Kp.|��n�q�n��y�<�7��4Qb!��x�`���]�<I ��_͘�v�U�pR+�Y�<�� |�`���O¡8��U�<y�#�b�I%D� C��M�<��S�kEP�q���<B�:lz�_�<Q���(a�,$Q�oN�h��)�k�\�<�����<j8$��	����	��]m�<���2;�x3�m݆|r�� 	j�<� �1�)��P@ƊSe����"O�1*���. �\ǩD <h	g"Od����^�,��c7똽E��@��"OȁĬw�tK,��t�ja"O�(㈚�nBH;�+��o�0�"OP,J� Y�i�#��T�n�ZЦ"Oʐ�1癣y]R钣�W:#۪ա�"OD���w���H��F�� ��"O,\�!晾�Xv ���)R�i~!�d D���@��N|�݊��=BR!�$1i�DQ��"
��!%���!�P�P�0�xA#Р7��p�%
��bo!�ğ.6�\,��n�#/�qZaj��!��P�{���� �g��bW��h�!��H���s��=
<r���y4!�D̚c9���wB�= 
bE$�d!�$�C��@nˡ-�6� ��m�!򤔣>YT1)U,�>+��Ⱥ��˓R�!�DO���ԒSa�*C��h��ΏO�!�7[��1Y��PԈ����u�!�ϖ�F13�
̏D�Xi)�m7�!�d�1:%̀��R��ƨxW��+b�!�ĖCX�"��ۨ)�����Y��!��.r�깸��4e��@�s�ҕ3I!���1w�����8��P��1E!�DúBK�e)�a�Xo`0��;-!�ɇf��I�(�*6d�����V!���4r��Jǎ�CW�p�L��bQ!�DX�"�q�R)�#T\�*5�Hj.!�ĉ�q&�H�%Cָm;.����g0!��+�\� T�>6���غu"!��G�poG	V�u����oq!��S>A�LH)�.۴I��J�'�!�䜖Kvm��*K4�b���FU� X!�D�%$����sȗ�Grl�����:5!�DS�R�P��HȰ-�0��NmJ!�D[�7�)�����QƤ[6K>!��q�6�h�H��\�@H��ᚎ&!��\=l���a�<���R!��h!�$	�o���)�A",[j�����^!�d�?s"�� ,qR� �uM�:I�!�D�6V���$��UD��A��t�!���d�fIQ%-�ɋ�JQ�'�!�3�0����W2��t�5u�!���<H�ڠ�VA=t�I�ꌀLx!�\L0��"無��G2w!�d!�PЕ.����bG�x�!�DI�g�����K�p�ڡ(X<W!�d܎0�mC �Y�T�A'L�Py���"2�~�	'�x�(����y��_t�t<+LG�JA����)�y�VrE>�P�`K
��M�QJ��yȆ�5Z2u�g�W%b���I���:�yB�-voPC+�=WO&�*���3�yBe��)��t�UN��OL,� $���y��\��PH�I�����yrA�%$b��6�?F@�pP6��yr�3Ī�)��O�J\�u�ˎ�y�*
>o��	u'/{��c%���yr΋"�����Ȇ��<����y��ۣ6z��8w�M
8M��A����y�j֘V��0SJ�4�fm%F��yrOM1��p`F�>C���
��yg�9
|�C�+]�+�TC$�ʂ�y
� �U�#Sz�b�� �2!Ȅ�"O���tf>@��i�%�Wa��h�"OP�̝�f$0���f4 �U"Of-����	f&�)r��&CS\eK�"O�lp�f �e:d�B����L4"OR�(�N	�T6����J&�
��"O,���F.j~�\����(`���*�"O�	��ߍg�<�U�Ѝaw`0��"OJ�2#�3º��M�&�H��"O,,���/nt��eKبa����"OD,�e��5uTN1k�8�*�q�"O�,��̇�R�q��A�x�"O�`QB�^025P�;�+�g��)�"O�A��H!v������F1pY��J�"O2�a��S�R��a��S�{2DH�"O���D�J�.\�ÞK4LKs"O��3��-V|��25�O�%z�P#7"O�|�tN;b�l�b��,0�"O� !���j\�YZ���HN
�(F"O�5b$�����8P-�te޽i!�$!"ٻ`'����sE#�n~!�䂕/)Lh�"�Y*ih'Y%p!�P�L���� 0��t����!��E�L(p�Q'�1��8A�!���;�2I�4&�ި��I�)!�Ǥ,*^=�Kޒj^ёU���f!�đ)x��593L�da�Y��Š&j!��oYnq���
��L)��$S�7O!���F��$ O	��T��#�L!�E,p��Ty��3�6]v��E!�d�)���c��c��r�>'!�	<kWN�Ô�>-Jm���!��X��,���OE�ՑmB$�!�D	vy�#���2Y#,]�d�߁x�!�$�h�����ۺT�1�d�&hf!�Ď&/
�뗅%���c�̙GR!��M5&-���F�� ����$KD!�dP�uG^0�mA��*2mV�A,!�[��"��㇀{��=�P<*!���2^W���+!�
�3�%�=!�6sr2��.̙�8h�D��+
!�dִ/���:Ţ�'� �X�F���!���\��]h��Ҭ`x�)ҵ��^�!�d�t�0DA��N(v�`1�O��!򄞸|k��qbEAD�쑚�O�x�!��:}&�vfX�b�H���J.w!�yC�2�R��� �P+_!�D79U�5���#=�Nx��#�{�!�Č�j�L�q��.y�R��� �!�[�`�L$��Z92�T��Ф�#m!���WL��c`٩x�����"��:!�7D���9���jz"���#��Py")Y(KT�d�f�M�km��OD��y皽`� ��%C p����S��y�G �~h�Q��W9:e�G���y2��8/���d�[�PS�TB��C�yB�D;y2�b�#9�̤x��y�@�/ܑ����`*�b`�N+�yrk&-:pY�4�'���y�C����m�. T(���y�H۪C�	4&���� ��k%�y��� IA�	5C�lu�u���y���j~:�C#l�(�V��2MG#�y�FF.tۘ��U�;8�p(9�)1�y
� V�5��?��es�^9x��Jp"O����75����V(8���"O�8���11���W�B�x���*�"O&T
2.��=��(�K���YV"O�mB�gL�B����+ƦH��%`�"O���fG�9wc���#j��&�aV"OL�q��S��tࣦI<Gw�}�"O��1��ܹ:{pM�L�=`� "O�����3��pA�l�.�ʵ:2"O��³! "��`��E���H��"O�V�ީ'����T��I��"OT�Q'�\�>y���S%���"O��&n\�z�W��X����"O�����z�j����?�\�H�"O�����kXVt�1 ՋV��ݫ�"O�uӢ/о8*lS��R�0T"O�	b�IƸb��H9A��]�@5��"O�A�A�5N�,E���["~�F	��"OBظaE�U�b�q���"gPH�"O
 Do	
#��;d,�%YG  �	���'��1���.1vH���-�>���'°=�Ui�UWr%a@��'�δb�'0|�S3C�u.�AH�%�
)�����'㜬�SB�H���r$V���'�����8O��$�̅����'��H�E��/L�҄œ%"c�1��'sj]���F���B�M��T���'V��&��[� �B��ҷ]� �'ϴ�P4/N2 �`+[�3�bQ��'pr�*�OÍBȒ	�G�3�J,�	�'JB�g!*k��1�g^�&�&��	�'�@�{�L)<<���
�1L�NU�	�'�Aw �A0½��-�+K�^ɰ�'�h5B�1!b�<��ݛ?��!�
�'jL�jZ�d�T��(����
�'*i�vnǔS@ʌ3��#2T�8
�'�l���Y=hji�a�:OD��	�'���#Κ���L�A@�J��2	�'�.��.�`Wر���C�Bj�-Q�'�6���$���%�4o*��'4�v�Ɛ@o�����K�)�p�;�'� АP�Ҙ%B���
W�R��9
�'�N
u'ޜ+s������P� #�'H��AA�0�0���T8����'<�a��(ڪO�m�$��X�@�Y�'lt0�t��L�� ���1M��[�'Qb�§a��}bF�h��#&`���'jUpf�F=�|x�E�X�_V^|��'��K��ʖw�����U�^}0�'�|p�e��sv��h�`�R)L��'�ڡ��䝐.w �xA�}$,��'�.� �5Q�,1P�K�x!H���'�5��-_���! ΋vF���'�h��].N��2�آi��t��'�nI+Ui��X]Q�"��_~����'#x��C$M�`�L�g�R� ��'mX�/�ڔ<X�G"?N���'�Z��Q͟�z�&�*��@����'A�T�c�0:���3�G�?� P�
�'�ֹ��W�6�����JwP�q�'=����`ΙMʘ����u��[
�'�(� P �b�0�8�ᙩ3H,��
�'y�p룭ǁG�68�u�ѨԸ+	�'�n��A��s�.����؂���	��� 6dys�S�]��e�)r��b�"O���3/�$8u��@�DD+!�����"O�hr!D�-Jv�Ku�5J�U"OV�j�Iܛ"����!�5�Pu�a"O�h�Øs��Ⱥ��	�~4���"O�m:vmӯP�Z|@g�	ު9�"O ���'�I2T��B��tjZ<�#"O��/�v���)�DO2VM��"O0z�\L������%N���h�"O]���ѻW���X�&�A��}#�"O�t�`G�,<8��F&��vx��"Ov���o�0pn�,y"�6��`�t"OD�R������i�f�0��4"O,0�5F�7;6h!΄/9��\�C"O��BP(�+K�D��6�ط�	�"O~�����:]��
vȝ�r�pH�#"OĉQ&C��|�y��H+%�@���"O���b�8�Н��O�*��@��"O:��`�1I�(�c.��H� �(�"O���$�6�x��C|�A �"O�l����I/�聲�S�Zvޙj�"O�ɲ@�&eT�fA��
_���"O$�6�K�Td)�j;��8c�"O �7�_�	`�!�r�I�Q����"O�њ�]C�Y%G�#Y���b"Ozx#C/�7��:We�IZ��"Od���5{\���#�+kʀх"O�D(��b~Ι�M�a�xB"O2ؐ�
�+����	Z$�YI�"O��
fO[�>� \s��'q��퉀"O�i��Z(@�ǔ&bt4C�"OvԉI_�̄`%�����I"O(ɂ��7k��%Ʉ�̷e{ɀ"OT��t.2 �����M�etm��"O�t���B��m�N��|W 8b�"O�]Qj�ײPSa"�3Xk�U�0"O�@#��R�Qh�qǁ�5C[pU�u"O֨���^�$�y�AV�Q��	q"OH��JD�=�f��E���P�"O�2��(��SU��*���R0"O��z	�<I�۰X2R�z���"O�zq�IMƦH�QEʍ���"OܡA�����r1s��O�^��x�"OL��dBѾu�x�GM�B���"O41��F�6@����ȉ稽QV"OA0�\�s1�m��C �/����'"O�ȳ�ȫO��h�УL8:Ƚ��'�Eh�'!y�U�$ʗqe(���'�~�lJ-3��o��e����v�.D��2��C�(L��狶��93��[ʑ�"~�	�::��;v��O>��pc�+"�*B�-6���%�E9�|a��_�Fc��F{��|�%Q;R�I��$ْaR��?9�'�Ve�o�#^�֘Y�MB�9i�8��a�Σ�+�
.�=p�DqY��ʒm�K�tE{Ҭ>a�@�7eǩ?B��"A'�Mی��'�ƩAa�_�"
�h)��(f:y
ߓ�M[M�4pNVQv(C�익i��ˇ��>�	�&�H(��9k�l]�h
�AI
��ȓx��y��̇p��ԩ��O����ȓ$�T�b��	^�������ńȓc���;uN�󆄃8z��ȓlkeh5J.D��a��X�Kh�u�ȓo���$���:�
$��"�����S�? NK�fV�Z}cp�S3m2��X��b�'��V�"�B���L٤eY�4:�
ʸ�y���e��2G�Z/��xR��N4�y�d���Q!ѵ!��k�k�'�y�'�b�(Cbܙ,ChH k�EӾ$��'.��ZcD7b��mp�.7]J�i�OR�'=�S�>yP�P���(�7Ѡ|a���ny��)�'+�~�+��7L��	�\�$�XFxb�'�,8$��"]�I�� V< ��=+OT�>)�}���<$e*��^2����f���y��X+G��Z��'{�V�Jm@���'�ў��̙6��!YB��$�v�q/�yb�La@����"�� ⦐.��'�ўb>�a�)KT� DG��Jlhu,���<�t���I��-t#�v��8cQ(<��4m.��UEY�:����E'\?lT�ɄȓE�p��w��$%�N@9�?- 9�ȓ���h�O&d�3@;�p4��u?YI>y��
�Mhj�d�qS���s�]j�<�rC�Qy�(ye%���`ū� ��!A_�xD{��������IX%���b������6�S�O�����R�!y6�'C��~3.h�'wX�f��:h��89��W	y�l̫�'�ʑJ��B!	��� Ԗs����'?�e
s�դ0O��Zv��\B�S���/�t���@:.��a��:o�x��r��`�O�꩛т��oo�9K�E�	j^���
�'u���9X>�͈刊+Li^��'�ў"~:�i�$<�b��R����E�M�<Ac)O4}`��3��D�P���A��<q�gӤ��$^q6@��&ɝ�0s����� 30!�䏦:4H���a�l�p@�'&(!�DL�}�Q ��J�h��j�`G�H!�J�,���G��u������-� &������" ��R�2��'\�V�lCK���D1�S�O(>�F'�39�:p��$֥�Y��'���
ӫҧ	��`F���O�q�
�'��a���_�F<�ԘUl����
�'�D�ka;��Q0�P�O28
�'{�r�ς#������g
����'a�IR��ԬD&���N�e���J�'��,�'�0�D=iϒEx$
�'�2%�F�1t v!d"�#(ox	�'�䩐��A���93��~$�`�'��	x ._67�}�/x Z�'�̈�g�H�v�p��nJ�NU<��	�'axp1��T5����1	O�0��]�	�'V@4[d�5����4�4��9Z	�'84���M+|%��4JJ�/׶0��'~�<���O�(����N'{,�`��'$<�J��_�_���Y$q����'^��AO1wf���Q�q���{�'�R�7��Tw��Z��,g�>���'���w� �D���hC�&�|1B�'J�q�_q:�8��6o��|��(:}B�)�S�Nm�;��L+ud��s�L�H��7"�S��M��ȝ�7D�9Ä�,��(9"�v�<1R�2gu�m'L��m�����F�<	�����$�u O+v� �i�A؟��DtLA��/��� G�ro���ȓ#���C�Cq��2�c�t�"9��Yi�D��/:��Q(��� ��<�����!�v�	���*{�V��u�x*!��ǄN�.�SӉ�O�� P�ɓ7!�� @�Z�OɎ(t�Q�� #$�A�F"O$(�ce3M�|0uB��@�B6"O
�IC�O@�Rc��=zH��2�"O �0�B��� ���9���s"O� :#BA�a�d�[ǁ U.�<�f"O�5z#,UE�Q�'��1j�yE"O2��� ҢU��\���<D��"O �� .�M�l�tle�.�0�"O����&t6jY���L��"O�-2s)W��Ԥ#W�ƿ=�.�z"O�(Z��M����Ws�}c"O2 ���� Kw��77�P�
"Ob�[�ǔTA�`��ӑLe&}Ò"O�]���[����ԇb�H��"O`ٕV\CE��~��0"O� ?]w̤���
 ��`�"O��s�ͧ�!Z%L��� �bC"O:=�w�����"6@C
Ď�AA"O�%�2�(���� �zĺ@B�"O�I�
X� W��G!_�^�	�W"O$z����o�HD*���r�� "a"O����劣lj�#��X\�pXp"O���,R@�V\ЍNT�"O��,�P��	1L��v����"OZ�``��0`�M���	7�Е�"O<mR��EW`Y1��s�w>'!���)5@������nG�(��!��![ j��2R���҉-�!���3^q��A���(�Ъ�'&9!�52�j����6Q�c��J�"!�D[�k�	S�$z���(��:�!�dQ5m�X����&#R��c�ײ5�!�d�$H@]{�
�m]�8��H�!��^s�Ir�A�Hz���P]�!򄋊x��c1�	��S�ֳ{�!�DQ�n�~�ï��k�hI�Ǧ�1�!��A�,��e��Y�R+P�؍K�!��3�L�j���iX4����
<�!�C�f��EX&1cZ!�� 4�!�D�;2YJA����g�J��&���|�!��	^������~ 4$1'�pz!��	%-�\I��7e�
���C�h]!�$F�B�ء�2���}9�#H!���|�x3�͝��12���AB!�:(%��%'Z�t���ۖ�F�A4!�͹B�*�����?��`�r� #<!�D	�t��u!��a�9q��G!�D
�޲)ѥ@� \(��ʡ�ޝD�!򤌗P���`پpp8�bD��!��B�D�cBh�Y��P�9�!�䆯s�(��g֮X��e2�AX�Hq!�$��+K�]�C��6sw�A8#!X>Sj!��-Mc���jI�9b��0�A=�!�$�3=���"��F,N���B5�!�$^�|��5��Uҹ��A��c�!򤕗J_p����[-0�B@�F`��9�!򄛿(�B-S�#A�_�:1t޽\P!�$A�W��U��jL�����Dh�!��Z;s$�ATC��9&*����^�/�!�E����ɠq�	�d�U��!򤀓K# � V�[�^�l� �i��K!�$�=$��L* �b�~�C�Â`!�D<ZM�Y�窖	 ɞ��DH4!���k_`I�c��3l� ):5�QZ!�� �X�u$V)p��l�#QA��0�"O�-0(3�~�:g�&Y"B���"O �#��3:0 q$kַJbY��"Ob\�נ
(0��$�0�)Ѧ"O� ���ؽe���� �,��DҀ"O��#�Gԛ> ��]�3� l3�"O��ũ��2j�H Jī9�jي`"O����kF�>��%���x�RQ�"O����/��(y)���K�H "O�� ��J����3�#z�"�)�"OF�a��D���AS�PL&x�ȓs�JLЦ�C�tܙI��C$[zm�ȓ{��9�ꔼ#!b(���ɋy��)�ȓ="��aiФV�$�g!s������Ta��H�4�DÄ������'��pU!p(`����~�P�'�����k�1|n>�ڄ�T�E����'<�� � �/@BL�4�8�&Ձ�'���@  �OX���K�;0|V���'��+�bq��Г@X�E���'�tJ��[ Tl����aʁ{�'�����[/� ȒR7i��'W�h��ț$%�A�!"�	��Ճ�'q0Ia%S�HHr*�!�pM�'!R�aO>:q�=�tkm�z���"O�X���'8�\���G�/��&"Of�H`�&uZى�C+Ұ��"O��U�˦\�n�9S+��'�a�"O�8+�C�m�6������c~��U"O4�Ս̇>L�#�,��l�@�"O�x�"��t���ۂ�7-��+�"O�;�o�o���)R�j�p�"O��q���\ᆕ	V��!����"O�, ��+`�Jq�#�L(*�Z�aa"O�s&$��N6]���]=ih�1�"O| #c�"Q�:��� �?���{"O������	G�p$�Uϓ?\�蜢!"O@�Ee�U��	�>��雒"OnĈ�/O�Δ sG�Z�8t�#"O���dW�3�Z�e��F��#"ON=�Í�g�d\���vU��"O�ab莕T���GC�"F��l�"OV�W��&����З.��x�"O�:�狂m,t���C%V���c"Ox�Z�p��Jp'�Ab��� !��?��H�T�kk��3Q�ʢ7N!�Q�Pl8�@��0Y�٫E�̓zJ!��X�4��0��@S	%*����G[7r�!��8������Q��&���G
�!�C$�*YrP��2aFH5Q!�d�5<[τ�	��U�����!�d�d[�E��nР9㬩��.��	!�$�	e��ra�P��P�'I�Fx!�d�C��I0�睑���Gƴ�!򤇬u���c6�A���p�GZ�!�Q�<-��ѯ>��@v#�:�!�$�!٬���O,3/�-�C�8�!�$�[0+p(��UI��Q��!��Z�3ʄU����*ZG���k�!��&k><��J���"�"��;q!�$�yW��x!CZ)
y~�i���3Fy!��%EM��6�(Hf���@��No!�пm��xs�&��%���Ql!�$��Z+x5Y�-ܢ;�pp�˥#O!�� ~؈ĄԩM8����â-�~9�"O*d��
��}0�h�#oʆ��"O�X�p�7���x�dR!��m��"Oh� HC�P���N�y�j�J""O||)A�]Vj��#ťU�.�:�"Ohu!�{�j�"�m����"Ob����C}���!Z�L�0��"O\�� �F|�CU*�k� E"O���ӈh���8@LR��P��"OJ�:PIB�,��dPF�9[�<��1"O`�I�-	�n�����b�0�b��v"O�T�-_��P�"���
"O|(p�T0&�@���)|�N��P"O�(��܂.S���/R�'�
�J�"OH,���P��vMB�"$D��!��XT�F���ͥSU�$�� 
j�!�	�[�����ݤ7hTH��t8!�S;x|�4"���v3�ij0�J2#!�DL-~�l�7�,W"L���e]4!�UW�`xe-�88pX����0�!�$�0=�Ԥ��	-+`N���Ǆ1�!�$9EGZ�B���\>4�"5-·�!�$�i*.@�hBl=V�� ��"L!�$��~5��H�cW�& ����V+2!�Dߐ-q>�2�Bs{�-�$k<!�$�PN2�@V�'�Z�)���-}�!�$��꺩Jt��s̊D�\�Q�!�dX8z���*2Z%�֯��!�d�7v��
Sj6(Mn9ĀM�+�!�1�@��G	">����U5b�!�W�%�.,�t�ڽ�,��D�I*S=!�dp��,�G�y
���@���O9!���U<LS#%Q%.�r�zPAP|!���7��}qp%�!�2����K�!�Ğ>,�*L�'̜4 ڞ�z��e�!��]�X�[��d�]��O��c�!�&c�@M�f����ڤ�⮟�!�DA+�i+�fE��%G��x�!�D�sp-�"��7ג�[7��$�!�daG���4,���s &K�z�!���i8@ ��N8o�l��N� !�$C�f��"ĩ3]L���
��5�!�D֣�x����cNy���D	w�!�dY�0���9P1�H�J��
�!��(i�4qQꗠ'<1��ވ` !�$���Dj0.�����*�_�!���	��QǛ�v�� ����Fo!�BW��#҂���m[`�O�@`!�5Df� oL
ѨU����-W!�Y��V� �k�x�����{H!��6kӴ�s�	 ��apZ4!�X�~ >E�&@�Xk�D2�/��=M!򤞑\b��)��V/DK�4iϖJ3!��ɱN�D�����L��k�I�f)!�$�0��]r���c]��@��ܕ
!�ʧ�|���	�|A<	�͇8"!�dV�.�9gȢ�v��g�)!������j��)���l��*!�d��x\��+7�8kv�ѳ��B�!�Æ\8�ܰG�7_\�Pq��:�!�Y7v�M��Γ�]Y�)���;C!�D��(���XV��?�~)�J� !�$��R�`� ��Hz�qʀJ�!�D�[N�ӑ��9Se���n!��  c6�|���s�[�X�!�f"OZ�(q/B�o��}
����r���K�"O�$��M�I�,�eT3�&�*p"Oz������}x��sCW+ ���R�"O*�sO��;�Z�`џE��<�"OL1 �G�`p�4BS�n�^Q�G"Oиq�l�*yt�tJ�'�1W�3F"OV��!�(T�!`�VkRi�"OJY��Ût��{e6��Y��"O��۴���W]�6�ʉ$2\<��"OL) ́�|�4���90 4"�"O��3J� J���E�48A�1�$"O�|Z��[9;��+��R 1�.� a"Oڤ�̀��>����ܪ�"O��XլV�gA�E�����DC"O:I�w�P#a�$-y��MQ��Z�"OV� �jnhP1��d3^7���"O<�1DL�
 �4}�Sn�@	����"O�pk��І,Y��,T0d��f"Ot8�	]F�d����XL$(*�"O����ф�n�2g]�<
#�"O@=�N̏~���� +,��d"O(����X�O����BְXL̲�"O�#�+M���%�D"O4�L�|$�{��*�l� p"O�ك���b��P�T;5�1y�"O���C�L2.�j��Ll�Ȑ""Ol�g��.(�I�&	�sm�`!"Of���C�$����n�/vT"�3"Oؐœ�p$�v��)@����"O��KP��D*>���͚�8:���"O���@K�EdLTx�bܮY�u�e"O4��gB��&2�XH#�݄5<@�S"O��)q�ʊ/�xy��Y?:"�"O�E�v�M$�du��͐I���"O
X��@:i3�D�b, �B1�eq�"OzYK���1,��Y�+σt�x3"OpH�w�_pj���*ɏ&�4v"O@�䋟5 ���lN�\]p�	�"On���I@�p�+$i rYZx��"O��%��^�vh��HL�HH�e�!"O�A�Dđ�X9q��'RlD"Oޔ	w�]�8�jp�§W�"g���"O�F��5~�R�`�-�'RJ��8�"ObY�Kռq�$��A�B: �ؑ"O�X�Hߗ;z��R�A�	O!����"ON��@"<<��)���w�td�t"O���W �� � �l��Ձ�"O�]���9JL
 	�����3'"O`1�2� Yj���2HU�mܒ�"�"O����~���1FY/k��Qp"OPk�`֟HD�!�� �k�"O��C��À��à&.�%�F"O&�h�˒yD�S��צ��Q(b"O�bE��g?,�%���Z��*�"O�L�UKƿIr6hYRN;<���"OV��U{ee�!JHB5���p�^�<Y4၇d����ԤJ����R�MW�<aL�� ���+q������U�<I1����rF/R�+l��U�<��-�7
��j��!3��ca�M�<����ة;Q�
��V�Sf��q�<�gGN?.��+���MG�ECP�Q�<�7��F$�'a�-K2���_T�<� �4a$��'E�Q��x��t"O�e�2��X���I8#&d��"O��f㐽q���f��&*#pa��"OXDi�@3l�JGӚ��-(�"O6A�uGF;9@���h����U��"OlU�A��K�X:P����H"Ojq@��Q{��%c�Dݳ��D1"O\��������$)RygH`"O2�q"�qĆDT���g,ɣ"O���O�6��F�qS@��"OfE�P̎�,�� Б���><X���"O8�Q(Jd���%T8/2��"Ofh��_�t.��R�ح]�"O������.<���Z�	��s"O���(�c7!,´�`IG"O6�je.�H$�J4�o�[�"O�ٛrmV%ahh���.��T"O^00��5xE�x��#���!"O��B�L�����wB"i�"O@Dq��
%�.%{��c@n��"O�)%o�7C�����;{4l�{T"O�`䧖�wn,�oׯ"���ٔ"OTi�BB��_A��  ߥ�U: "O�y!`'��
�` #W��I����"O��as�M��@�k���@ר���"O����H�f;p�Q�M��~��U��"O{�i��[2Dh�<�N� "O�DВlt��l��L�&"����"Ò�qφ�Z`)����>4|��"O�p����X��̳A�ڰ'���"O�X�V�&!�.uTmy�����"O�9�(�9��J� �0C"OM�� Ql0I3V�X�5_��z"O��h�9�2�z���
tWpeA"Ob]BE �%7+�����&C�sw"O�0a����.&�����΍J9��S"O<MQ���K5��2�h�x"��c�"Onĩ�X%a���ۀ�Z�w��b�"O�}�"��'�h�)���*�"O��Ӣ.�k8lJ�^e�L���"O̜25I�$�
L�#�Ƨ-<~up�"O���@�
�%ψX�'�X*|��"O~Pr���P<�X�Ē&�N҇"O��˃)��T�j��D�Q4�X8�"O���s�ͱBHm;g��@ڨh�"OF��&��)7��c�-ȒĠ��"Oډ0���� \�A�L*_r��"O �˵OHa��AI2�˷+9H<� "Oz@	��ՈqNf�
�7X1"O|�� sr�2bܵ ����G"O��s!F�.�B!_3����E"O�y��aL�$���˴�K�c��	Hc"O�YK �J����e�-d��@"O�ț�ϵ3|@�b�Ժ�Q�u"O:H1RM �n�`��7"YX��A��"O8lC��V@�A!��ݭ|�*<��"O4�b��;�yP��V=�$���"O�HX6E�C�t��W�ZH|��"O�y�1F�F��t��7N'��p"Oँ�DI�3�u�b�,���{�"Oҍ�'��	��P+"H\{��$"O�j���hG�K�hއ �<�9D"O:�SJUF� [��J�W�J��"O�y`�	�M ��RVЇE���#"O� ܃�eF�Bx�A�1YZ�TR�"O�|�g�7^��[C`�F|�PS"O����^�yѪDun[+F(Lr�"O�����V�2�Ba�SCI5�����"O~��C��.bk�W�h���"O��a�Ea��� �铰M��b"O��6����q�T<O����"O"Q:���S_4�Qp��CYT�RA"O�Ļ��	�0��o�/@ʸ� "O:�B�fRgd�(�� 
�P<�"O|��@�Я琼�vi�h�z6"O���%��6���#��ջи�sT"O�ѻeOP�h@�����A"O�[��yW���o��YL*��"O����ӿ���db�9�"O��D��&CƽA#�O�D`<�2�"O��C�Jس^\�el��=y�j"OtS����3��(�
��gN�I"OBD�	ёIa|�j�I��bE�Tbs"O��Z�d
�:���I��p�(!�"O
�*6Ua��x�.�l0�I��"OR%�a��>�ٳ�$S�v|�%�"O��F/�3cn<�#'
ע=mm!�"O�ȢG�4��a��$Dk(!K�"O�h%hÜL�ޡ���[�x,���1"O�	
֩ -o�XY�V46��%A`"Oֵ����!\V�QLR�
�^`S"O�U��*��­��jWx6�x�"O���U&�'J�F<Hv(NnΜ�W"O
�s� � bD\	��R%X���"O�	���	Y�hթa��v�\�8�"OP��Q�΃�TD��>r��"OP�CՅ9gv6��uDU�:�9$"OJU�扂�����B��=�n)�"On�Ah�?�
��n�;$��Y3�"O��i��8��v�G^��DB"O�Ƞv�A=QD��8��ͨz��q�W"O�T��O� A��Y��%�./5୩A"O�D`g.WT�b��F��51�M�0"O8aɦ�?�:��~���X�ȓLAN�x@!������q���s�!�$s��k��A�B�:J�+ �!��0�j���!��Y�T	����)!��2.�!���.��"D��!�$��H�4O$Z
�2g��9�!�E�W����G�,x��i�V)��d{!��5s&��� NZ=$�F�b��E�n�!�d�S:	{�̛�Kb}�aרE!�d['��!�qƞ/y�>5

Dgs!�L�,ZH1��E�t�rυ�!���"%� ��|ڡ.]�R�!�D�
Ԝ@�gѺHM�`�q�Ůi�!�dM(/����#�1j4��@l��!�X�Ռ����F�K������&!�� Bj�\���PN�ZT8�H_,!��-4�<	�*��9��UЃt�!�X'e5VIBb��3J�xP&�Q	�!�C�=�XUS�DN�"��Bq�Y�!�Җn&�|������P{����)�!�C��V�)�b�|���=U�!�ėe�m�B�Y;W<�a�͙�~�!��=T��G�Q�S?�Z��6=!��l�H%o՝0
�\�a�9K�!�D�*=��x1"KC�JN��'@�Ta!�� �(��Lڜ|���]OM��h�"O����(��|�Z�#3���Nc�H	�"O�%4�؟!ъq)F/�.3F�]
�"O. ;�U=�Hy�g�ȅPy�`"O�ip��c� �WcԧR�L���"ON�#�_"�2��Ӣ��+o�EX�"O��hdL
:P�'E�Bf\pcV"Oر�����LI�@���7_Rp�"O�T�煘�V���{�!��~@��)�"O �𗂈�H�<�C &L��T"O�1Ba���$�ZXz1����*���"O�Ԩǎ��N��qk��%� H�"O�"3�S�H�z�X�g�K�05�V"O P`��Yu�$�d�!a񈹊�"Ob\�DD�Zz�#�j�*�
&"Ox�:��S�]Xt�Shl�|,V"Op y6l�2tI���fﮉÁ"O�b�B8M�q a��E���S"O85{��O"!*D���W/E�$�"Oi���%=R�@s��9[��|��"O� 7�A&e*�H���^���"O�t
0�8�*Gɑ�Rf��"O�K�.vy�qE�1)�j�:�"O&� a�&{�4�ė�q����"O�a���'U���q��7Ƅl��"Ox���Ǭ%��@��ų3��J2"O�9�*���nL;ᩒ�F%�Q��"O(���P"&ZNܘ�g�)e�&�Q�"O�`�����؁[D�h��Y"O��p�+!:�0�d�4Q�T�Zd"Obe	5�O6q �M Tm��`��P�c"O��З�C%�H;��*p��A!f"OniI�/19t�C4��V�p�"O��2��1�� e憕I��|�"O�y�I�,���ӵ�
����s"O����E ��Y0u?�ZԂW"O�����[�eK����<��"O�3A�A�w a�������"O�]�C�!�
�)5�/���p�"O�\���̅h��q���CO`ЀB"O�	��̦ ��$,��k7.͙�"O�x���UFH����1W�${b"Obػц&s�4���9Nk�-2�"O�Uc԰A!d|���=ebb�"O��R�#\�>}�0��}�r}9�"O(Pa+��[�@�x�t9�""OP�S�˄�Cô��e�C�6т�I�"O�)�WD��y�H��_��p�"O��PFW1j Q��K�C�^4�@"OX�S�ۧ	���" \�P�aj�"O!3%��C5�@�
΄%�XHRG"O������N�����Lv���u"Ov��$Å� �b�+҆Y�jmL��5"Ozs"hۗL��uPFh�JUQ��"O���gj�2>�Q�)�3Q�5"Ol:`f�Z�@(��ȉ�&k&1��"O&#S�X;�f�H$U�$�t"O�Z����EVV)ʳĕ5�1j�"O�,��XMRbw�����@s�"OtxC��={�^D���M�x�`�"O��ՈO�xD`�Q$O�("A6���"O�	�fA,=�^�����>Υ��"O2����ˈp���,��Hm�5"O q�d#�M��aSg�#/��D"O� �@E��=��sRm:͢i�Q"O�ĻA��G��xB��*C����4"O����I�Ґ1ǋ��1�����"O ���
\��,y0	p@ҽ��"O�FEEq���zeQg/ԥq"O����<�B}h��z���WU�<���H��1����,��hK2��Q�<!c�jE\��OF�-�Rc�GUd�<y�	 `�Pj'�F/2n%0R��_�<��7oJ $��,p�LY)fʎ_�<���=�R��!'�J������W�<)Ӌ��~@C`���q���賦�U�<�s��u2�Q�3�����R��0T��Z5��|ܕR"�%=4���O0D���wdN�]�b��X\إ���0D� 	!m+(w�q�׃�X��I��;D�H9-�eApK� VD���Cf-D��3�A1?/�@XQʟ��t�6`/D�8
D&E�δ�i���$9^��N-D�4H�K�`z,�B�A�>%0�
*D�����N�^�>9��CKC���R�)D�`�e�i@�P;2eɉZƶ��T�<D�����\/����VDF'HV���Ve%D�����*jS�A���t�x�b#D����E�!�$p�q#�
3Y|g`!D�T�ĺ`�`�2dS2��2�l�<Qf�ѕ$��{S'�L=N�Ս�J�<a����7�ޝ|��/Q\�<y�)��TIanYv��ㄓN�<�l(fڜy�Ō��YR�XH�<1�n�}�nE�DOd�l��p�F�<��ԐX>TT�V�ѕ,��XC�6T�xڃ�@;�TA��֒q�F�!��:D�t�2���Qt�$(tH�:p[ !�r�8D�,XPB�|
X��"R�PX�ճGi7D� s�/� ��<cvT��*(D�T�L30���Ov]bH3��1D��#b'F�Y*Ԍ	T�_-�>��n:D�xs0&��,���I%�Z���8D�d�3�՗CK�8���
Z�8�e*D�а�+ �%k���s��&-DP(D�p�g�Ha!����ZU���;D�L�'+C$J	���tk�1� �c��=D�(B!��y�d���T�c%�1kd�:D��;��k�^���h�;z��ʂ�6D��iG�%.�Դ׉�������1D��AF)C�	�T�Ђ�H�qT�-D���D��A�x�� �M7TD=� �*D�ts2,��Q^��Kh��&6��G'D���bٹ�1��3��}"�
'D�X��m��(�	@�)�q\�1��@8D���D�[�\s�MBV�C'^�()p��8D��C�jM<����� ��b����7D���.����<�� ��5$�3D�p��%��A��!-���K��/D�<�" ��2�X�%N�4YƏ)D� ��	މ{@~�X�Ϛ=@��}ȓ�*D�,˂�W ft��N�!:����+D�`q$mF�C�f��v�Y.P�Z@�uK(D�H[b�I��-裃\5�P���'D��Z�˥iz>)d�j��*D��a0eVC!�Ƨ�';���#��&D�0۠C��h}�dߑ_�����7D��Xs�'?��%˦ɞ�Q����`+D�� ��c���ZvD �G�Š�u"O6�
��:o3��WGɿ���t"O
*,�9R����#�l� �"O��Zb'H�>P,���=1�ĸ��"OV A#gפD���:�!��,�ҹQ�"O։F&�&~:��G��@�YW"O�L���'�pdL�!moT��u"O��$�Q��b`z�j�`����F"OXѠ�/��m��-�F	G�Pj��"O� ���� iJ��Jt�"O���F��>��bq�O�nm"J�"O���!M�2A(��F1o=d0!�"O��x��Q,�r���	��UǍo�<������r|���R3[hp�E@�<eeűkp��E)�9>�Pl�U�I{�<i� �i<%��+�1]�pHP��Q�<�C�|�ѓ���/h� t9��K�<��
�*�)��k؁`E����UF�<Qq K�W�PQ��?5��ڥ	�y�<�m�5��d"��˒��@�e��B�Ƀ���#�q
�@���QTB��"��}����v����ZJB�	�EބAQv�ͻ8Δ���E*�XB�ɵ`E�t�!|H$��`N�=d!���=Q�vy���4N%�e̋�$!���eh %����i,&�Hv!.��C�I� ���u��8.�f�yŁ؀��B䉐Y:���w * W|� Do�;z��B䉔5*�p��"��"�"8���Zo���\�\Y��!R6FcȢ-� 8!򤀳c��X�q��#eDŢ�,ŠQ$!�$�$-��Ae�~W�i��.Mv!�$V�m�H�VC�5wc����?[!�d<�<��cE8Fr	��@%,/!�$���M��ƅq0��i�O�!�d
.kv�ءw���`�X� �͵5N!�$�+E1���e�ЮA{��f�!��ɯ+�2�� c>o��9Z�ʒ�!�DNT9�A��-�)m�����H�;z�!򄈍4�d� �)��O���J�-��#�!�$�)Y�4�x��X��5{W�ٿD!��T�*F�x��O�fv���AΉ��!�DH/j��r��</YxU���K�@�!�D�3U:ͨD"̞(�`�a�/�!�䂒�����Z�)�$)�`aKh!�d��#g<|���b�t��bx!�$X3~��8�RLLb�6x���_$�!���ld�%��Ձ@�b�
�My!�$��X���Ò��!}<��:�)�'\!��N�]�%�qLM�,:�⧉S�AH!��+*�B�c�-�A�/�!�dZFc��L#b�Fam_�2�!�d�?z�=� ��5��i����i���=E��'����Dσ97Қd�T�]�Z6�*UO��CT18!��Ш��C���C"O���-E��dӁ(�)�zL�"Ohz3�L�KU���G,���HG"O��@׊�mli+�A�!.�\+�"O�W�Qm���z%B�W0r�Q�"OD9X�G/=��0X"�8H0V��d"O�B�X1�8��1 �./~P�#C+���<�'�?QI~�/̴��� �[�jơ_3B�$�ȓ6:(�	��¬*���K��u��$�ν)��n����@NQ�HF6Ʌ�S�? ��Yg*ޘ'T~,�&�Y6Q�\�:q"O|��b�K ��Sw ��k�5h�"O���)���l�F�IOep�"O xs��7Z�Dӄ ?����ISyb�i��Dq�q�Nu�D����bh!�ğL�>=r�=ݤ�wjX/�!�d^����q�b�e��@XG)CN!�D�Z8�Z��2�>m�#	ƽA�!��:^��yJD�F(8��1D�Ӕ
v!��@�`��p	Q��S\c�I�K>!�dN*'%�=�I��H�^�W�U5'��M����E +��9�a��s��Y��"Oܑv12�8*g��<F���"O8=@�+� 7��I��O!7��$�w"OĴ��R���K"NޠP��Q�e"O���O�0|�Bh�'"Yr0P"O:%�$��k`�2�0uO�A�?4�8������kՁN+�Z���6��?y���PH��I��(��Go<��gaҝp�!򤁿��EiD,teb��̀Y�!�d�
�l1 f��Lb& ��$�i�!���D�R�1"�Hm�L�⣈_��!�-pr�+�����1��ʺ�!�� G�5iUG�0g�"c���_�!��V��r��/�d�ۥ�\�&@ax2�ɛlX��w�˳��#B��(zB�ɗ}���0fφ�olu�rY jB�$o�t�мk{��Y'��x�C䉡O�ލ�b�F�2�f%�T�z�B�	6)��ShE�%5
�@2#P�)(�B�I+,[T-x�E��V|��h�� �����>��+:~��hC���7R�r�9�K�<я���*FZ�;�*ߒT����@�*d��C��.h ��Wǎb���XE"��F�(C�I�@��-���1Xv�R�ˈ#}�BB�I Y����6n1 ~����A:q��B�/Yh��D��\;"<(4��g9����(���xk�aR�$>n�8�6B
s'�B�ɹn��U(�ϗ?\I�sƐ8F��B䉦ze<|�paQ�o NXH��Q0��C�I�)H(ܡu��L�L(�E�B�zC�I1�4������w�E�PLC�	!	\F���I[����r� O�>C�I�zP���UA���&k��Z��D�OĒO����,�y
4Ҵ�׶1�����"OD�`րl0|��ݢ㪥)P"O�}��#.G�A�6��{�5��"O��vF
tZ([�E����"O��e%G!j��8��wK&œ�"Oz�[QD�=O���pt�0��t�!�䂒I�6�Je�݇
=p�A�"�,l�!�DD�Z���{#��쌅�!��D�hp�%�B�j�i�ذK�!�[^`���͌'-��$��ޫ.!�Ok;� �1g�H�PQi1ōd�!�$�R<�"%߰��p#�d z�!���n5z882���'��X���d}!�$����	�Ĕ�V��iQ3b�@F{ʟ�awC���xׇX*n���r"O(�EBO=
�!(��6j.8i�"O�#��.��4�6b\��H�"O� ke��k�� �㋌�>r\�!5"O`��͐��̘�red��M:�"O��3q-��jCX��Sg�/O� �a"O� �ુ_�b���ό6f"�� �D/�S�'fub�H�%� P}��*@'a����p~���s"*xE�DOڈyV���(��Ԓ�˕�3��<���Ft6��ȓ+� ��%?��*�e�!�t؅��1�GP�n9֕�$� #?�%��.,T�T!��Z��H
����TT��ȓ ��|sT[�A�|C�,�4����ȓ;l�[���1}>�y��p݇ȓ16��&��
�Xݙ2˒))��-�ȓo����6�\c��ӯ#��%Dx�'�F!)֨�ZK y$�L�]�u��'��@E�W�vn�aԃ��Qld1��'�L�*��tPC��FN|�1�'O�� RbF�2E8e���[$D�����'�P�*��wj�<
�Ai�]��'�D}���3{
]#"�N�Plz�'ml@3�F,,=61���NAxA�yR�'�:�*��H�Y+�4���g��
�'�`�20��^Hthhsd��� ��'��}�0�`o6(���Ӳ}r:)�'��%����2���C9Rzh��hr
L�ah��6�̜��-R�&�^	�ȓ	H
�H�����P�	4'*��f�u9g&�.M��]��#ǰVmA�'��}«)�Xp�4�6(�	\+�y�Φ?�T����7��ɂ�	�yb�X?*t�[��	�6���������y⌘3Rj�)����5iR�rE(	%�y��8;+�yP�B?uU>�1ejӢ�y�١w��\���Nr1h#�cD*�y��'S�|` ���y�Ejޓ@+N��'���a�B��`V#�5Mv��� "���y2C�,i��
ǋ��n�t����y��^�e̒�r4`�9ȔP��F8�yR-�F�"g&��ʛf4�|��'���Sb���	�0+�%bu�'V>�ypÂ�E=� @C�
�'~@��pJ��4H 0+.(�8e��'Iz�0�.R�`0�Qr ��#�9i�';H�{�K��u3tt�Ƭ j�,��'[�|���,�xM�ѩ>gødb�'�0��t�̑QV��#�J�LZ�'�D�UI^Wۘ���̰@#@�8
�'�:4���Ȯ@�H���<NH]y�'�x݊2��nq �0N��L˖���'DΈ����t�hy4Ɲ;?0m��'�:����zr��R�� }�ȓk�Pa N�:* �4O�-a`T�ȓc|�b�m�2r$�A�W�X��4�ȓ;�L�h���
}��(h�L�,�A��V~,�N�Ϟ�SӣÃ8Y�Ȅ���:�j7��#�Q=3*F����d3��+�h�;Q��5, Ňȓ~�|ȴЉ'&�%3��úy?I�<��Ί�X��l��&/�YCBf�<QL� `׬t�@.VR���^d�<yT�w �pS�Œ3��MB��z�<��R�o��Xۑ� -�4���s�<���X�p�r��h���w���ȓ4M�� �� '�����K�iW������!Xp�:�z�J�B-f�x�ȓC4���n��2�V<R��שX��i��s��@gK�/wc����V{*<��S�? V5�D�!���@iK�%g���"O���dLͺ+K�xK�
C���`p�"O8Q���P&y�x�R���E��64�����G0��yڇ-ߗql�Y�,D�@P�H `��9cb�l݈0�7D�`�I��d�8����ZR�tĸ0D�,�fȆ�D:�[��Z�:%ˠ0D��6A���ơ�׈لmu�u��3D�Xa��7Hyȱz�痧���z�%3D��{�]'9�d���=wG�����>D�p���ss���R�L^�\� A@=D��{qΆ0Y+���;!��YuN9D��`�l L���#��X�.(:9D���G,f�B�a-аo,Fa�Ī:D�`A�$��fD���N�E�Yr��9D����딠L�d��m�J��e�@7D��Sd���N Fe��l^�C���C+4D�H�s�`���[�M�����S5^B䉜U;���a�ב/��M�g���0�6B�	�p� �:�s�qz��U7�b���'����͛���2�쟃L���'�d)D!p���ʁEP1�(�'gl؊s�̫3�&��QF+:l��'hhUl��&V2H�g�(nb����'�l�lR�n�F,)r�Ӳ;�By
�'���"/lt�=��ϒF���'(i��V���Qe��	����'J�TC�'G�{���H1Ē�y#~���'b��W�����#F�j�T�
�'a.�P�EH2߾�	P�b$��1�'�&+�,�:BA�!G"������'���ѥH�E8\u��?����'^ \!`�\�=��#��?
���'ڮT!�d��9)F�h��)	n0e��'�z\�R�\�`\�r�A�|��`�'f�����j!�g��0}ߪt �'H��J�!ɬoRY��;g:Լ��'Vq�����*�//�h��'�@�1��=swL�XB�|ܤ�'cR:G�֍��Q �� �M+�'�b����_�^.p�₋9���
�'���Ht�ʰ/O(�Q����z�j�'�����e��(¤���#ɛC0�r�'ʂ�{4c��A��x!!H�9VX4�'K� �0�72��倃kޞF;v���'���� �,f��7*�1x�ؐ"Oz] ������6\����"O�ԋ竘�I} ��q��'6����"O����PI�����2k��e�V"O��X+�`���) IIsݡr"O6��ըB�gKֈ��!�>ox�u"O8�K��� 7V�D�叓<bvP!"Ol����Č����0NŕN�@*�"O�=�G��4L��,RD-汲 "O�uy��D����4B�!@�P"O�$8���E�� @�.f��G"O�5���7Hw�3�.71�%Z@"O0xB c�y�������~L��p"O���`�7ᠰ"֊�8m`ڭ�D"O�}�-ٍ��̻	�TV.��"OH�S�cܞu0��Ϲ�����"O^�j� �Sp�ٚ�@E����4"O�ɁC�^'5�ïO��ŋ�"O6$��)i)>p���Y�@�t�:"O� ��*P�݅Q�	n�`��"O���1�-I��)������R���"OR;�A�[ڐmB�s���"O��X"ISY��\�!����S"O����4:�t�֌^5�<�"O|�R#��,_D�����,����"O�ũ���$2��j�,X�<5��"O� ��E�3�*���,m��a�"Op�r�ϾU�� ��H�y�r�p�"O���a��~��!���B����"O\@���Y0L3ܕ�7쟮|�@���"O�1k���
��0��<��ũ#"O�lk%��"q�&4�e(�N˦�a�"O���ToY�9d.1������$3�"O��"��7M!���`�W�^��D�&"O4\��;u��;���j�bTI�"OZT���ߜ�t��ҫ�>T��@"Op��Q3L�d#�%��G9�9��"OJU�bB�{�Ӣ�P~:$	�Q"O�Q����9K�>����&0S�t["O`�"�H�-s��DDlNR�E"O��bD���P��-��H�!a���"O|�*�	e���SeJA��a+"O(�PR�~��8�r�@ .��E�C"O�%�+ց{x@X��kаS��F"O�ݣ�^�Q-����I�3tO�!"O�8p���{��X��W�<>��"O�t"�f1�~�ӷhH6CBt
$"O�@p�Ar��t�J�>�;@"Oh]B!�H��(���q���p�"ORi��싇�D�2�̗2|>ӧ"O�1`BĮHO����ŎP?�i4"O�뇁B�cL�!g�^E؂�2�"Ot� �/N]�zy�e�CּHg"O:�k��~6& a��Ǿ[����"O���K#G�|@bd	?6l0}"r"O�e�K=u�<h{���?oT<���"O(Y��	�=Xݸ hP�}#���2"OR�SAN�8����@�	TxH�"O���5�ĿYxY���'�|�)�"O��+��'l]^��c��U�)�S"O�	�M�`���oXJ�L��"O������8E��|�_�b�T��"O��SC��dd�g^7:h��"O�Tؗ_� >p]�ƥ��� *�"OXX�&.J7E�K�}�e:�kX�y��A�i�ָ���ڄ{�DL+�hA�y§Q�'H��d��z,��`Ƨ��y�(�Ta���Ec�(k�`Q��h�yҩ�
{��Tj\�[��{�-J�y¯Ƒ_��x��Xtd�D�Ĕ�y򄞚<2<�̐�F�T�Y���%�yR��
|�H!�g*�?�Z5Xs���y2/ւ7��d��7J�B�jA�yJKTqv�vƌ&4��lB��$�Py�I˺WM$�Qj�g��a��H�^�<��Mhi�A"��1�ԝ��"�T�<qr�����K�h"@I:�ST�<1qlʕ����jM� �nq1q��R�<as�ݯV�x��  ̘k�Zq�p�OR�<�'X�M���Ō
�l)!��r�<��K2%_& �$F�͞� �n�p�<q�m�Bq����KW$w[f�K��C�<Aƍ�4����DK�
�yR�'Tw�<� b9A2 e怸A�[�F��t�"OH�4�0A�zQ�s"O�����s���E�+t؀��"O��P�G��5_�B�C�.�ָ�"O$����XY��$\�O�fX��"O�����^7���T�P {��d��"O�<p'C��ݪdo�o��m��"OQ���V�p� 1#B}{��	a"O2ݙ�H��4A����nӢS\0�+�"OJW�NU�$ ���!p>�""O@�7��bF���c7�P�0"O x�u�Xg�����U*a"�"O�u �.�"��-ꉴD�2f"O��i����xaވ�'kC�UL9s�"Oz���ӆiq�ݙ�@�,�x��Q"O��p��<T"���@ ����< �"O��a�N�3lp��� Mʠ|�F"Oȭ�GN]{�l*4��@�<�v"O�@����%�V9�̀7d�r!"O��I�o�
����,���g*O��p�#�&D���Pd���<4p	�'��)�g���4,�I�h>�t8��'�<r�	�+��k�"��!��'� ��#�jT����;y��(�'�2��'��:�:�2c�,����'�̭����Q�\}I���(#�(l��'ܴl�Rm^%a��ŁF�\ �'�h�2�KUy���4�� ���'&T��N7Y�v�Z�*͢%y�'�����բ6]p�cס~��:�'��P
��gr���ď!_�t2�'�Ĕ2�d��ˢ����
� ��'�r�H�Q�_qtܰ č|��Ų�'L`Y��#�\L0���z@u
�'_�܂�+J�&�&�!�Koc>���'���a��%�vE"1�S="�A�'�v �e�Se�@ʼ����'L��Q��ۮ	t)�p��F&A��'o"D"�O7��0�Q0|%���
�'(�d����.�@�1H�Dq���'��}3����P�1	�d�?����'���� �J�fTe�E�
 ֒���'��b��',�eõ�4~Q�y:�'�؉������h$�N
EZ=x�'ud�{A�C>C�4 zg�=r�j�B�'��0R������#C�#8�4���'���X�f� �����E��H�'[Ē�&�1�i�(ͼw���s�'E2�h�#Px���0/1W����'|&�)�� @���++� =��'Dᣓ���L�	�c���e1�'y�8���& ����X����S�'�TyX�gµ*I<��aѸY�h���'gV��sȎ0K�2����B�?���'��=;�+���Z"0��]8�'}lQ�S+�$~����]� ����'gzMq����b�T�� ���$!�'H-`6 ھ@  ��@	�[,��'�yPgkK�*v��a@��>v����'��e��!W*n�\��'.�P�� �'2S�O�ڤ "�5h=r
�'�>����3C�h�b�����)&D���%�64�1���7\x��0D��i-�����X9]r��/D�� (`jPf��B�b�,5�!��"O�b��v��9�����'
 ��"O�l�4�F$��)*R��$C�4x!"O&�[��(y����mCp���`&"O*`6��S�5Ҁ�X,p��"ON����_�85�H�pN��i�%"$"O� �0b�22��	��}�l,Җ"Ope�0�.:F� B[�qL"D#���v�'��?g���dH�)q�D0�����B�IǦ�"b@�$�V� ��O7tȂÉ12�98���H�@� ��VoI]�v$KB�Y/w����'w�����o�|����I�N,X���kzqO�6�ϨO�+��ȕc�*i�f���­��\����ا���i��I��
I:��\F����2z/x��I|���3CI����ҠI	)��b7��hO��t-���+��<��a@j�(���� �$�/<�YS��3<��g��`�!��69�r���( ϒ���H�!�䍆	�H��ؚ�tI3T#B�N�qO��=%?���␰�t�R��6F$8+>D� )T�G��µ�ע-�`�=D��BJ'L���؆�ՠU�L�j�/:D���U��y��h)�(|uB��#D���C��3
���2��8���-&O#=1@��E��L�@!	�VH��a��'��b���3��{C^�J�E.L$��i�<A�	�<Y�S���DJ18֥i#�_�~���@����$�>�ܴ=l�)�'F�Bhì�v�4��/|Rȝ�ȓ'������_�4��sk�o��'9������j0��!"��ʩ��d�KhD��[04����5O0��#�	
B��J���:�I`�'q ���^�+��Tj&%M�?G���:6H��BD�r��2��5F�l�ȓ?pđ�"��y���A`*T'\U"m�>�I��<	�{��O�NO-SZ����)A�2��M��Q�uw!�$ϰ/U�U3n�`�6��)�{s��Ez��s��UipB	<,&�-B҆)*����
B֟ȅ��1�l- @���R����BY#kT�����O� �S$��7��-SD�h�.'�鈟�$J�3	p���`�ΫM�&U�`��+�S�IL8^�v��G���L�;���?w'����(O��A�7��q�g�ى�` ��F��ȓu��s�`��>�m:�B���'1��F~B�Ov�	,3%��b*O �Z@I�/9b{�B�Ɇ9L�@Q�O5P2|*��k�"=A��T?�C�)W'TQX%��@^:=�
���+D��p�d�A��z�W�v$����M'}��)��s���	�N�J4��`�5?�Jl;��i�O87�<��A�:p��č�j�"L:��Yz�<��a�=ފ�PB�w�TAZȄ{}r�'�B�q�a�z��9��*� ?֠m��'��1�#E�h�xa��,9�ˎ�(}2��O�'H�:���T+9r0� u�VbT��L֍�n_�#�E�"�� z�imR̓���sӴ��4BIT��/�;p�Ш�U�(�O\ӧ�g~�-z���cX�@��5c7c ��$3�O�)kSD�E{��SGD5.J ��x��'�h�ҁm^ �p���g܅#u.�q�'�0�r�	Z ���%��#k�D��'�`$x� B+�� �p�M��"������R�Ob�Г�҅Si*�����$ ��1�'�h��ce�=)�&D
F�AR��'�>�ʱJ�Tj��3�Ѓ;IXX�
�'�9����vh0U2`
�(3�H��K<��S�? ��"��8�|̹qoP/7]����"O�C�O_�3�F�J���ư��"O�1��Y -�V�Zւ�4����T�O�d;t���VS��U�ÅG	�i��'e`��L�R�0�B�+ʺ�,O��=E�d�L\!8T "��!O\�JEO�5�y�DI)�X��㓠
���N���y�,'�h���GK վE0����?A�'�ff�5��Iɐ Y�,�
�'ɘ���+�3C�p![`A�6�<Ջ
�'��$b��W��t�D
 C)>�)�'��{��	G���H݈E�TX�*OZ�=E�t@�"{�T��TA�>�a��&Ĉ�yR�����7F�?A�
ě��R��y��-T�2D������:1�B���p?�O��KԧT!R��H��B�o66��"O�aR�L��j9<I$-ͨH|��Z�"O��F��9ls��aEצ2̉�"Oj|`��+OF|M���жӮ@��"O�e�,�:����bV�U��YqE"Oz���ϕkd�IGaۗ9�M�"O-�5�V2�)�т�8H�Z%�b"Ox���[�l�s�C�L?XX�"Op���ړ%�T��ZFf� "O�X�fQ�D6��2��Q	e b=�r"O��`Eӧ}�j�y���2V��a"O�����ސ4"���?"���#"O��$LːK�8S�E�phY"O(-�́|�$%#�O��EbZ�Y6"O��f�%����N�,l.0M��"ON�ѳ��2���BD�O�1CZ���*Oj��[j����RO�5!�r�r�'[��d�?�l���C �HDB	�'�(��KG-f����6��`�'�\���ތ h����ľ	�l9��'W� E�ޖ�0�� *K�9s����'n��"���=���P�þgn~X�'��]��f��l�p#�Y�8 R
�'sb�aM>\����ލ+|���'�x��	�S��Iԣ��w��Tb�'���PcÞ�;���)��D}+�L)�'c��
Q�$dx����y�⬀�'֖t����A����;�~m��'���N��1�v�(M�7L�Ɂ�'�h�Z�V�rvr�ä$`QB���'"��窝�W<���g�"���{�'�>X f� PXe@2�م�:H��'��� +Чr�|���`�Ä��'�갨QLE%9i4T�5�	!	����'�nLё�ʡ3���h҇�%olj�2�'�5(�l�N�1K۩f�D��'�f����^�2�2DO+c��	��'"��P�GĈ}����LM$#6�s�'��=;#�@']S�0r��0[�x�
�'�6U�PC��O��`J��X��	�'�&X�W��&%�`
C,�xO�;�'��Q1��ƾ8���#��j�����'������ݧ�VC@#��h���'��S�	`��@HJ�Z1���	�'d��1��V)Al$���ѬL�d�b	�'J0d����Hlzq���C�x��	�'�\��1���h�0 S�FS�� �'�ؐ��,[�:L���ؘC͹�'>& y��޶�1���5��	��� Q$�уQv���L�:F�n��F"O>A
�~�~��r�N�#\�Q"ON��D��86�ıQ$ٿ}�.��"O�LHB�G}�n��Z�a�"O�`B������V!R��h�b"O�ِ�	�k: �;��]95��QH""O���w�F�j�X���"��#D"OV��w N�&:m8��p��8�C"OZ�G�?(��f�\RH1�A"Ox�Cb%6 F��cb��ik�"O��z��"��u����V�h��"O��R%&R�)0f�/@��|  "Oxq���N����+��`��J�"O�ԙ��Γ_|d��Z{D�!"On�8 �N� [P�Q���6?l�1˰"O ���C�U���a�N�,�q��"Op1�vN#%,��(�!�9=��9sr"O����E�71���OKk���F"O��jaE:�4ja/�*D�z]�"O10����'�(�ò��� ���v"O�՘������Fɔ*�ʘ0�"O�6��)V:=��DZ���"U"Oѓ��E�~`�Q�	<�:��"O(a
L��y�*e��nҎ8y"�I�"O�HCc�D /� y�5u��5��"O()qTB��H�		�O^.%cq"OPa��O�x�	c�O�=sμ�s"O.�r���Jl�����Η` �@�"O�9�d��Z�ƌ:�EO�9V`q�"O��`f#��+�l\h��ߦ)8���T"O:�
d`�4����7�-��"O�@�ufx�$���H%,��"O��͙�g;T9�"��Ff� �"O�}��\
�py��aߪ��yw"O�a�cʶ>�
s�J�,6Jx ��"O�E����1iR�@��)�x���"O��؂�ת/�X�2I�2Yx�]@�"O��ק �P�h�kШ�(\rDAr"O^(�n�^�*xaш	"�`���"O�ld(ÎQV]2$.��2�@���"O�����ݛz&���C,��1j,"Oh A���b��a-P�"��P�"Ode�U"�TNB0
�P����f"O�������\خ)��)�5W����"OF���Kx�Պ�iY�jH�'�j01s��`�x<($�8J  U��'�	r��N�)�ؕr��O��l�' ����MԷ[:���� Q�[}Y�'$�58��ȵU����qF�P���A�'��e�S�R� �R�
�J:F�|�'i��W�_�4P�	����'���D�I*��·��	ԩ�
�'��m#���ˌ��j ��
�'�ʌ�0G٤���Ҩ 2|�2
�'��=�%˓X]�(2�ڌg��z	�'���QTf6-BY���ǅ\ʸ���'��|�!&r��i�U�D!Nޢ���'�섑E�61�pSR�Hm����'<P���*P@��(bK9�*|��'C ���o���'���#��(�ybc��%c�\��-!�!��x��,�ȓ@ε�a'�"g�|�P��ǻ���ȓF<�Z ����`�t�,z�"O	S�A3t��2./a�f��"O� ��u����<�������"�"O��YgY�D�H(J���0�~�x`"O���::��5�̷cƬ�"O�R�L�E�b�;���(�2����$1LODT�._��"�ړH�24��͈"O�b2M�e���{T�:z�q�"O�����q��7�8���h�"O���2L��(�왑=��=@��I}���Iצ?�v��jQ&R\Ӆ�ͥi��'fў�>)w�U�;���5gH�3#���l�'�qO$�V@���)hH��s��A2O�*4(f"O�)���%4�1��(Q���yV"O]pto�Zbl�"m�H������'c�O%С �
��8��,�J��h1�I]X�0��̒�wN2��i�n�H	v�*�O֒OD��%I:Sߎ�P%d�#/^�:"O�8�-�
bɥB��]R�hæ��7�S��$���!D�ph4�k� G}XB�	�'�0H�áF�IB�+p���x'�<I��T>�hG�^�H�2�$�5k��0�<lO㞴P�$�v��{�#C�k7\��<D���$ÚD��q!�/@,7:=�;D�X���i��p�I_�p�
����$D�����5W�&$����7;�H��`"�IA��P��j�,K�a\�#������%?��p�p��4���O!��� ) %튩�ȓ^ߘɃc$B,vVᰐ�X6TE�ه��M���C�|�~l��E�gޥ�u�X9�hO?�I���Ъ�Q&`�b�^��E"OR���� (y�S6�+�� "O�|Y�N�6�5 և?fX�C"OxH8K"�\�8�&R0�A"O�<����*Xĝ���(�t��H��-�=gYL �#H

!ҝ�'ܽ*<DB�ɐ�dM�1KZ:�%ف_$B䉏�0ՙQ	͚qg6�R�ɖ -��C��"Y乡bÜ<�*���`�����'Mў�?1q��T�H]6�Asm@�B��! �!D�4�@�Q�d�7ݕ}j��!�+D�X�l�m�Iy'K�7A��4�5D��[�̩_v:Xb��/݂���3D�8��̊D���B �";�&TAR,���ēd�)�)9��2�B�y�̀�i��10g���C�I�Q�"ʆ�� o���	��a�0�F{J~jf^�m<X�� �9�PRS�L^؞��=Qtǆ��4y�
8�fٹ�Ic�<i$Ƌ6Z�����_5?r�QǠ D�<A'ɉ���� &^��e��%��<��aŽ7����yK��薏Nx�<����+j0�RRi	8b*�!��&�u�<�B@�)v�C���>&)�2�즍G{���iMt��%%��(\m�ԁ�'�����HO�a��)��"��'H@:jv�"O��{C.�g��<:� N\]r�˶R���I&)N��XC�81XP�a)#k&����/�!z=�e�e��;8(�Ҡb��O��=%>	�C��3���私�c��j��.D��@&�~6�{ՋE6C�ܥ�w�2D���Ǌ��E�Z��Q(�!.���	N2D�4x�`N--�L�2��ޤ��tA� 0D��K0�+C����������8D�$�p�Ѧ{��5!�N$=�ֵ U5D���A�i��A��4��l��2D��*��_�2�8��ܜM0�¢1D�� ��ǫQ-���)�+C�6$}�F'ғ�h��dY<8��jV	�J��8�e�?!��a��
d'�.�.�k�N�T*BOR��gD�gA|ț#��I7��`��'qO�u�ǘ1�J���36�8d"ODa�G* x�n�R₍�p���B"OX�A�b�	A�hulP�!~��D��^�Ovܘ����U�oޫ��,��' �qbJשy�T�����
DҕA�'�~0@�n��k��z�j�L;.�ȟ'��6}r�'����Fj/ q��"��6X���'΀{�K�Y0p���
"��`p�'���PbK'�����aJ�z,`�'!���b�Ӄ-%��&X�^0 �x�'�rTs�o[�<�|��a��`�b�'6�(���ѝM�~)ƀ�Wv���Ǔ�~��>i�4k��a���;��( s�A�#d�\�'��	w؞��O��D�})���=�^����<������ O��b	���ޅ��L����1��`�3�"�� ޙ`n|ꓠhO�>�S�D�v1e��h���D�&�O�&�ZȹROޥ2Ō8P���wj��ȓ==������o�b���1��&��F{���H1Kk.���U�{N��OA���'�az�D�>*��W/Mt��m�cJN�~�)�'s��I2�	۽s\�p�+/2-�T�ȓ��`�cD�}H��-,Լ0lZ@(<��U;�t8��fr�����}�<iČ���͠�'�+h���YGdy~��)§6_�� I.*|��e"؜?��Q�ȓ&�ZiI�
�1^2��Kb!�jH�`��#�d���N]�a>�p�&K�l�Y�ȓz�����K�W�n�`Dg2f ���'��D��u��)P@�[�ml�m@D%�5�'Pў��<�g]�HG��J	�v"�P�MB�<a ��N�֝c��y�E���WF�<aL@�/�M��$�'�(�p�OB�<�� 3N�(��.\�˖��Q�Y��̇�,�(�ǔ{�����%�9B��O��8E{�"Ԡ)���[�We4���Q�7�!�$F�F����ۯ�r`2QaR�V�!�d�I�$��$��(x�6��ǥл|!�d�ZƈU���Sr��𡍆c�!�DȈ-�,!��M�u��m�E�Jў�H>,O�i��c
��o���B��.E;:!�M����@,�B�@���$Q�~!�O�jf���O.��\Ч��
Z`!��
��p�fj�>v����%�<l��'�>!�#�j~� ��z:�䃔�,D��Do��\��h���G��H��O*D���so�|�p!J!�T�gɴ�Xt�4��(Ox�J����2��0u1�i
�&X�N��ȓe4,[��H�j�dDhE�-������(D� T<zF6� �׆i�i�ȓ
�B����,o���q#��C�|�'fў"}�)޸��n±k�j�%��t�<�Ae ��l)9]b(��+�[�<� �˹�l�H�ɨj|6; ��Z�<��{ �}'I"jo��Q�C�j}R�'E��r⚫n�^PX�\<4XX{���Ɩv���v��Ap�,�"Y�o�!�$G�I�Z��p�_u��XP���-2Q��G�d�	Q�����9{���h���yb�-�Ŋu	�@��
���~"�)�g�? ��x�蚡4��<iV̓�VQ���W�	~�ax�,v���r�nK6b�ȸzg��y��DI��@d	�]&@�;����y��	rxQq��% i�a!�<�yBNώr5��DѤ Y�������y��ؙ9v�8 ��$H�p0+0 ��y���9.��w�n�0��S��yR�åp�Ь�5�A����N	gt!�D��0�(�[�� �2~�!�,H3.U!�dӕLS��+��J%phŒ���1tR!��(fd	�dU�sb��ـ���nF!��]>}9�-�@�G2S&J��aI#f!��$?�6L��S�I&⍫�.K`!��~��0r��T����!e!�(N���A�aU霓#l!��$�D�K���9]&0bӐN!�d�XƵ(!GC�DE�`P"G�SC!�-i�U�0���B3�9H�F�2.%!� �_��$�B�a �)�E�)M�!����jMd��ENֱ.`t�S�!�*�)C�W�����lD9z�!�=+�	@�a� �N��鉻zU!�7o�J0���&DSxӔ��?-;!�d�t�nLA����L��q�[�q�!�� ��!��� \=�� �٣�!�,	���1NήL;~!�0F@1.r!�d� Z~���[Ѝa���W!��&L�� ��5(
�*�\�*!��M�6N�(xq�҈{�� ��M% �!�#�H��G5����C�\F!�U+e�QC���~ⰂA��!��-d:��AF
��L@ ,�=8�!�$^M% p�O�s��9�e�	/!���9|�4���&D�y!���f����5�� ~!�$�c���B�C�M�&�3C�Y~!�&�i�֥�>x�\ӵE�%!��ѦjM>��ǣC(Li��I5��!򄃒?K,�b���Nzݳւ�s�$טJ�&Y"_6��C0�"�ў`��+�[�Xl�W�ԝjP�g!D����(^������A�qB�` Y�B�	�TLF	0F�ޡ[ ڥ�WcF!l�^B�I�4 ,�� �ӕ[��=IV(�$G+B��)q�<,��D��Q�� �:�B�	|���b��M��HVZ�k�C�ɢ\جX�BȔkx�<9��کK��C�	�:�JQb"��GO�(�6ǚR�B䉣D
�A�k/h��� M�?��B�	&K��}�ɒb�f���/�<F��B�I�b
`�8!���XbxB���+3�C䉵F�����C�mb(q�D�̣�C�I�Z�$q�$�8��Q,Ʒx�C�ɿf-��_��|���.o?�y�"O|�c���;q��4�݅k�Z��w"O�d"�ンA�>�D���d��7"O4-t�#)Ȑ���d�5�L�"OzU����a����#�;j�|�"O۪�V3"V��R�5mገ��"O��%��0^պY3A-L�h�J��r"O�����T!��p�Oلj�4[b"O�%��O��#��(yMS�zIF���"O�a�V�+O(�lS@ƈ`z��ȓ�\����).�)c�I�LV��ȓ,՞�Sc�Q�V����"�LiVM��S�? ��b�D�9��(�_�����"O��)B�+rD�q(��ZVM��;T"O���LG�w���j�$@�t�ur�"OJe�a
J�dԫ��u�r�c�"O� �2LՐ5��H�炔�~�V�c�"O�=�FĠv]���v�32"O"X�U����N0����(P��າ"O�H:Vc�,N҅��G'��0"O��5g�7ID]*'GȐ���0"Ỏ�DR81W�٭Kƌ�Y�"O� �nI0 �Y3eO%C�ɓg"O ����I����� �	G��� "O2I�N��H� ��!�I��"O\��1�J�D��{nʾ	��E"OYr�.��9���؛P�e�"O�Xf�tn�R�	Q�D�̘
v"O�P���@6̡�϶.�Bl��"Ony�e��@*��Qeh��)�*�"Ohi�S��=�r�7��0��$Q"O�9*���6B@\��ŝmwN�j"O��Q��Ja�)#�#VU���"O�1c)=��,�b��F�|@j0"Ov4��F���ؙ #��zyR"O��8`���k=��!� C
w�b	��"ON5�u��9	�8�so	y�2��G"O��[BG�)�L,!�ڋ�Q�s"OdL��A�o'�q����f.|�j�"OJL�1�?D�(����(F��G"O�=�P�J�c�NjX6
�J�"Ox! �G�Y�,<!��n�܀k�Q�̢F�)�O���3�ٶiق�*��:A�N`���'�M�I��@"��^"S>�Z���Z���6D�\��Ā<p���e^>H@�Is��6iJv��rc�A�O�l$Y���.��4�Jˣ4�1;�'cvղ�b�[���2�Ǌ��LA��L&x��y��9O>P1T��63��� � [�st"O\C��-j�%ʗ��"9�	�76O.���{a|b�S�ܼQ�H�<8��+�%�0>q  ��[V&��z��-�EC�9B��d��5%0^1�� ���Af��=Ō��b�-�PDy�Έ#���~ĩ߿-F
X�d�T�+N���Qdk�<iPI
9�IQ�d�?�t|
����M1��<�S��M3����U���vꎻI��"�b�<�D��8~A�3� �2R�i�7&�Z�<�WmY�=�����ċrv}#��QQ�<��e��f]�lX�G��J,㢀�d�<�(�5K:\}���V,B�BP��a�<a��vU2�JE�F#���t�^A�<���	�
�yb/ʦ�D-�Q�`�<��	��4�ܙ��:rr�����v�<9V����3ЊS�<t��P�_2�yB*�~���U_#;�8t�����y���"�	
�#D�D��(X��y�	>�.D	�٭/.���`���y������P"rM�|�%!��yr.�~��峓��9>n�phͰ�y��ht�Ŋ7hJ�]������y�&ߐ��}#Fd�Q$��9g��9�yn�$QEh	r��ؔMcL@wGP��y��5�j6&�#.|H��G(d�!�4GT���"ƣC�6l�Ά)|�!�DP�{���؀؉cv��֤�,�!�d��t-�bNMc,]Qސ3�!�$\�0��hv�Q�	���V�ҶJ�!�� �!��H�T$A8�/Ȅ&u*�ss"O��;�#^�nXzQ*��Q|q~��2"O�в$ ʹV�J<��MO�Fn<��"OE��g�=h2У�ȅ8fZu+�"O�]�mܦuq��0��kw�1��"Of�"�
q��t3��W�%U��w"O�x�/���$@R`�A �)D"O
�I�$W�n�y���ʑ)�$�b"OVeS��P -g�qj���=	��"O��f��;e�<�g�,Ql}a�"O �r5�M N�.�+A��'\JL�"Op��S��c����$��$E ��"O�M1ղ@6�,��Ă�YI���"O�yA��ڏP�tI7c	0�H�b�"O��K�{���#�cҫ>��\ȡ"OP)	�$Y\X`�(�3Q
G"O�L�$�ʬ1�N*�֙Q7� *e�!��5Qd���4������Ğ��!��̹3/08Ae�;y	�):��G�Xz!�$�i<>00!�T%2����)�m!�� m/u�%O��<q	�A<7�!�$�%����e�׋�
1�F��!�@�?��
 ��eL8ԛ�fK�`r!�d؆2�@<�D�Ͼ{Y~�*PW�!�$֫y	V�
QU��p��e	�!�[�<�ڤ)Gf��f��k�C�2*!�d��FMP�0�E�8RX��s�bU�rz!��J05TjB�02��
gőT!�$F+1�Кe�Y	�4#Ч�5^!�DYhp��%"L�##ȗ>F!�d� m��] �l��(����� F!�DȠ�D�� �8E8
��ǜ�l6!��U����Ft���#���;�!�d\�h-he��8��D���D-!�$�W�U+f@�5$�:���*�)E(!�d"ұ���K�UV��is�D�u!��\�s�QVB[�KJf{eȓ�mU!�9%����e��R#�0A$f�<`H�x��hH��<	��ڻ_�h#��/Dv<@���M�<)�E�(��aq!�W��;�|y���mZ�k�O��6er1"c_G=�tc#gY�B��B�I��~a)�&�>`��c��i��9�_��iT#� M���#K|�>�DOW9��	����/J�0��O�U����V�S<^��q��.��y�.����Q�TU�)���ܖ~��ŉ��'gz<�@#�-�b�ӡBԝ5���Ҋ���2L�Ba-�,L�I˟��&-ÄC�HMʕA	)'H�� �"O�����eЊ�q0
A�+l���t<O��qV��H%��2L�M*��ӳk������ �1���ͷ7�LC�	:h�PI7���2�� 9�ꈺY�6��ѦH՟�1��G�����H2Fx��lg�l��*�^jl$��$L��0?y"��sݞT��-�9<������w���x��'���3A��>ae��B"�K�gQ�[���P�\�'�@ЈC'wF���ұ(�S�~���A�����"�o��B�	o��� �,�z���1.�d���	�Q�l��I��q��O�O��]@��X�B����c�� �U�<9��2�N|!d�ٴ=wX��⾵G�%k��Bu�U���*�ZX��O��:0�И��a�&K�*R����'(�eZ���T.8-��!�� ��(@B��3����A��i��'����vFD57�
�+ǻ�$����OoaJt3��)#�z�kȟ�X��ʤ.��,`�d�92�,�U"O�x�$�P0�\�gI��"�ؙ��O����D¼H�I�N��0|�4��
9/��������0D���_Q�<i7��1Bp��חQ-���$CwA�˓^]@�0�O�9���'�.]H��޴clp���,�n���1	���*QP� �TKw럊 �<P`!�6u�y�@�5u������d��r"�Q�R7���3nV�j������G�N��yr*�IHl�Q���ki9$߰�y���c������R�f���#CP�yB�T87�X�t��R�	��ބ�y��� ZZ��5HI"��7���y�f�l�gW��S�΃1�y��PL�^e�pL�L�<Qу��y�%�nࠪ�뛅M���ba!E��yr� %�j(�t+�G6��p��yR����!Z�_�0�d�`b���y�h�)J���a�1;f���'픁�yb�]�	C^�R$���4"�S����y�m�<��u�D�+�>L��
S��y�� �6��l� %�����Q��y �$I��P�(J��!�-�4�y�
7�^���GKF� #���y�A�U�|#���1ܸH"�g�3�y����/\��;#bC
-��0�,��yR$ĸ~�~�d(P]{vb#�yr��%qo�� ��ےF�6�A�Q��y���:{$h���7bR�$ڑN �yr�Ք�L]�C2F��cN�'�y2 GB�´̛�)�Z%���yRl�"^�8�pTR\�Τ11��y�Z z��1)n��(�(݊�y�ަ/<��f>9(I"�
��yB��"�:V �!|Ǧ<˃Fׯ�y��X��s� t��|�A���y2��	����wnŉuW,�D���y�M�-��)D��9�Fh�p�V �yOچR~bȀ��ݤ�TrqJG��y'�>9
M�sLҮq��-(ɖ9�ybh�'���g�lގ��P�yB�г4g2��sIW'f�T�����y2�� �xH	��UV�P%-R��y��2N0H���O�O�^��q�E�y�hB2t5jY�d���8;&�#�;�y�ŏ�i��Y�)֥4_Z��Mα�y2��G��tB�F�$V@�z7��y2�ܽJV�ș�`-*h�چ헏�y��n��� 4���y� �����yR`U>/$���d��*R���y��7e�6�0'�RI�)H���y�#U�K��L,0�̱JL-�yb(�6��4�skM�0	4��0OW,�y��=ͮ�K��C#+n��'�4�y��H��ZEsV��4V�K'�H�<��+K�Q9��SoH����2��L�<�A�߿R�Z��lHtX��RJ�<9E���7~���۝|��)(s+�@�<9�jK�f��|�bi����V�<��D�x~l(Hf�<���K�e�L�<�1NѦk,�ҧ#ǘ5v���0_q�<y�ߠt.Q0��0��K�7_p}��o���@L#C�v	�pl]�B�*̄ȓ�@|�͖�Ki��ce�"T�l��}\@��o��+r�P�aF�$ ਆ�O��b��=kih�1�a� t���ȓJ�t�m@2T��& e^��x��	�nR�>�h����	ir���c�|s'9�fEPb�W�Vԇȓ ���\H�� 0D	��=�ȓ2:ܑ�l�>� ��M���S�? h���'8�:�@eĵy4D�$"O�\���4͜Mk�ذ{�B�"O�(�+��,�dد$4�-��"O<���h
S}�tKR1$�-��"Olp�w� (��Y:��&���q"O0H&E$/�Ĕ��
x�=�"O��1�.
?�1�� Ǵ��+�"O0 ��ۀ,�`��C��1��`x�"O��Z֩�z��G������j�"O�<ScG�a��C���� "O�!VCĹ&ͦ�Jc�"�laF"O�|�d��'�xi��a��V����"O��g��`�d것*>��+�"O*�`��ѱ7�� �5 )S ��"O<�xVU&}��p��O��[-6�W"Olh@�捱0��*�HG�"X)�"O�A�`�Gt�%����"U�F���"O��c��Z5Ck�ly���(:�쵺P"Obpم��A�$��i�	���"O0�ZU%�/�&�1��r�4L�"O�]����5W�XP1gÝ�u�l���"O�0��
�`�``_�f��a�"OR���J=f��%��*.^�{"OФR4�J&���6��%F��"O쑴�G�^a;2�V�TR؀ڇ"ORT���"m(�� ĉ$"N��"OH�J���y<�����A�(ԝP"O.	Ȟ�uyn�[��:)� 0c�"Op��ǑuОaC$'�3B���!"O�Y��+Ʊx����晇1���@"OR<��RO&�d:U�ϥ=���4"O �#��	�|�QB4!,�"O��	�Q)
<8B!�*"�`{!"O)k�	�?d��w��+�(��4"O9��c�K��مhJs֨9�"OJ����PZ4,�$fD�i:�8�"O&m��H��cF�e8AA� (�)�"O6��vb�R��h�E�`Js�"O�P`"��F�\Q��m��JP�{�"ODE �?f�TD��,Z1$��$"OhzC$Do�j�!���0z�j�"Od���O� �
-�U-@
6���"O2��T6��JO�%���s"O��;0I
a7Lh��CV�@d�\�E"O���%G^�(����F�ۜfx� S7"O�q�Dk
'g�v��a�g����"Ol1Y�*C�y��9�vң�܂t"O8!��Y<�H����\`F ��"O:	�B�@"t�*A`aRi_=��"Oh����WH��ƅP4 /�`�"O,�Q�� �R�J60nl!������y�)1^�u�v�1\b(᱑�y"��2E�1�A�?K��S����y`�F���x�"� 9xɑ����y�ע6>$��P��<��l��D��y��0<���c�(e� �T��y��K �P�z�(�)m@���O�ybHG�v��V%��\�f����;�y���s�R����U���Q�l��yB��>NT����Hr>��B�֨�y�O��X��D�>4$����>�y��*����Y�y�.��%>�y2�%	ᾜ)Ug۴|���bu���y��y`谰g�ʾaV��qB�ݤ�y
� �Q�ХN�{��2v+T�.�(@"O4���G
+q��	ط��6<��Q"O�$� I�H���YD*�3�,,i2"OP��%�
��n8�����B�pW"Od�2�I%<�Hb��?J���1�"O�P�V�M��=asƃzD(��"Of��k�5{����J� ���{�"O�]�CG_7�Εkw���C� 1�2"O��c���~��倄�����"O0i���5�D�C�N�+��d"�"ORUbҍ;
�}W-�(`n t"OP	s-P�Z�9{#�$-�t42"O~M���:�A��W.}��4�D"O^-��F��%��P���B���a"OF�z�Hz�6	S�޹/����"O�a�!��Z�\ᰨ�7u�A�"O�4�T�Uح�!��x� 8�"Ob�&�%,���Ơ2݌,R0"O��u�
�R��1������A��"O&��V���dL�iqMF�m�~$)�"O��J�:`���kE�3l�) "Oxh���vj�4��F�If�F"Oʄ�S
,D����7,�t�i"O.X�%�2oݰ k�k�8M�`�)�"O�d��NV�^;L��qȖ	~� !�"Oz�P��! 4��$K�Z�d��"O�	��a	�o�$�a�NЌ��Z�"OT��6��W���8��P�M��,��"O5а���n?�tQ��Lg�����"O.��ѨH="1(����:�L�b"O���Ů�&^��eբHi~)� "O�Xɇ-�6����I>)lF��"O�L��w[�mxӈQ�0�8A�f"OH1�'BV=#���ņF'��#�"O4y�A�JjP������Ѓ�"O:�c��Al�l �����y�X�3"O H@`A-�Y��f�1|� Q��"OJBD�$|��r�E���$��"Oj��d�8QnRqY���b�vD��"O�1�%cP�Z%�}�W�v�H�X�"O�#ӎ �2���k�@X��"O��;�)S�?�l�e�Q�$L��"O�q�'%ӂp�AТ��8�x��B"O�|aGE�\��%p��ݡ3�x0��"O����ME�8;� #A!͗( �f"O�$2��WD�݀W���f�N��"Ox��AhX��<���xr"O�+��+R��҂�Hc�]�`"O�ܒ�aV�'�V���<kҘ�t"O"�A� !Z���R���(�"OP�����6C�ԘY7a�R�|l��"O�T��kap�ֿ
źQJZ�LA!�Ĉ�b�,�y�M�5^���W���
A!�D�9]Vf��#��f�x�0Q�!�d�p����w�0up.���)E�!�DU�:��@��2�4L�fĜ�Nk!���b8���A� ���%�q]!�ŕ0�ā�6�$L���ELNH!�E�$ �œ5D�J�C����
O!�$Ձ8��%fX�o�,)��	^�<D!�$Ȝ�*�ӵ盵G�P����!_ !��9RA���lQ�����р�!��%g�dM?q�Ġ�1�R��!��XA�6�;G�
�J S�C�:|�!�� �=:u�±;��@�J�,�jٹ�"OX���F�Ŧqk�ڭ-�Ip"O�<�3�%�A��C5�,P�"O
�1s�_!0�B��rc�7���"O	:f���=�����*^B�	%"OH���<9z��Ů�� Kbg"O6�ԔAN�j�2C�j�"O���@�t�>UQc�Ӗ8Sf��D"OUD�̝H��t�	MR����"O�+��Ϊrݖ�zr�ޞ\Z�:�"O�-�C��~��͈6�OD��"O��R�M_Ek�Ө6O���G"O��;C&�A�ԃ��**�p�`"ON���]5�1#�%���ɲ�"O�!"�e���hH%�1�J
�"O,�z�G�&�z�h������0"O���D'+�|af�#yn���"O��h(� r�J��\���X�"O��2w�� K��\� M�u�*�[r"O��R��#j�
�� ���C��%z�"O��A �Y*c���՝R�x��"O<��	(_J0�`��yJ�u"OhYj&�A$8��er g�9b�@�"O��'��F�Јq��^����"O�5{�NL�`i�ၑ�ܧr���5"O�Q%쎺A���G�)H(|�s"Od�Ѕdv��A+�ꎷ7*�p"O���wK�8m�� u�ҽu��g"O�<����r�fԺH�@�B�"O��{c�Y�8J���m���"O�T:���<�z-�5)\ 2���"O��l �- }{����i�`e6"Of=�&��BTauO�+ɴi��"O�<AJT�w����GD�X���"O`�)3*Y0"KtTb�h&_�v �S"O�Y��V�%����G�����#"Ot�+B���l^�I`����(,j�"O�����30@�$����}��7"ODh:aͰD.��u晌~bv}��"O�ͱ�dYk �q�F'k�a"OH�B�,	�L�⥏�2���q"O�e �	ߒ�r����%���"On���^x�T1w,�m��,"�"O`�h9}��%���iY�1
"OH}�(CH�@g Ȁ6 ��KV"Op��T�ޑH�F3�FS;I&pq�T"Or�xR�L--�U�g"In�IS�OvQ!�h?$�8�K�m�d ѥFW�r���K�'����vkF]nP	[�cՍ~u�mҡY�.���&�0E9T���'��p'Pu�gy��'� � ��ވ��陒�ݝyn̫��$"�S��2�.�cWg��n+
1����՘'*ўb>%؃lڢN>�1�BΫZ�"���J3?ً��Ӭs5�}�o_1� ��(�.G�*C�� 5���bC1q9u�ϣ]�C����H����}����q�N�<���q5�+�hO���<:>(��	k}���Ǝ�?>*Dc��G{���▢H��] �f:0o<��A�J����-�S�OB@��焔�lJ�T�U&J� �2ts�'Oў"~�a�C#b� 2c��0v:M�1 
�7:0*�/`}�I�Pz7��t���N	(S�B��qG��,	�e�1����ɖSX�����'��-	u�
����ٰK�"�z�@��d��^ɄYn�)/��p�<ڤ� Q�d�օ;���aV${��Q0J�l@�Ų`�<E�4LϽ ��LF;S%TM� %��Z���3@�@0�f�;�OvцᓪFkSdx���1%�%!JP��@T06D��) .Y��O�X���-�܅��ҳ$bt˄���~�\ ��y �f>� $4�`ËgY�D(s,��q,�"o�ep��d�e�$��_���)�W�:<{B�R�~�~T
EbY<Y��{5��3'�.Q�G�%P%����i��?�@&+C?�n�"�Eϑ2.ƕ��m��d�0D���F�"^�!�B\l�����S)G��b�n�2q��Sk�J�<�z���&��D 'J�%�T����O)�|GȊPE���fŭTa> Z�"��@p�� EČ1oT�B�C"���Y�'H︔�B����Ta�B%xOE��������' �T��D�?�G�T��g�4!��n�����+�ē`� ��G5<O6	Q��	�(�8��l#kr9�A"O��� �ԟwܵ��+݌sM��"O�8��Ş��=FJ�19a��"O��XoK�/��PtnE9c%�l!b"Op�H�nR'R�� �+��7%�A��"O<P�䢅�BV &KG�($��"Ox��CĞ�v.���
8��"O�)�p.�O{�L7 �\���"Otx�Q�ҡ"`(�3t	BH��y�1"Oȕ� �Ǩx*Й�I&� P"O>) V���y_��b4�"�T�q"O��(B:jhљt��H ��"O��2Ä��Jl1�@F8�n���"OLۂ���q:�$JD�M&N�h�;�"O$CU�ӭ<�<��i�lpZ$��"O�����r�*Ġw+39�l
�"O��Y��+h�ءEm�5��ؠp"O�9[3���O��u��аw�nPQ�"O |�6�,)G���H�=�l�Z�'
��)Ƨ�D�b�OY-;����'Lb3,�;j<mS��=�� �'��q@.��ĝ�}�ă�'4�9ys�Ⱦo����'y�Xq��'�.�B�L߆i8�#R+s}���'RFI�R�ՂR�T���ƙk*����'��<�3�̧;�0�S%�m�(U�
�'����EӐ1�y;SER�8��%*�'T�Ei`H�+>F�ABFV,0C��'�FСVƙ�}g��V�#�=��'�!j��Q�D�.Yi�H���Q�',�a�6J�{��-(�-��|�,#�'O ��C��D8��撵q� ���'tP���
)A Z�`X�f�$�c�'��3P=f��� �iH a�pp��'�D��φ�Bh��GFʞY�`��'>hL��j�'e� ���͜K�l �'�e��U� �L�F�4���X�'r IR�!T�aD��6j�|(=(�'�N��D��>{ł5�����w_��3�'&�1�'B�`�p�%Q�A�Z��
�'� �U�f�b��T�W�3����	�'�Z� �K�^�`0Wk��1`���'��L���ʇF�l!��E�+�p��'�n��cC�I��y�T$"�P8��'e�����7�PY�n��Ja �'Ҙ �r�߼�T0�R앨�T=��'�P�����#7�u�q��K�y�'\��D-W�P�!S�l	�tW�!��'K�}��c��q��-@�n�<0��'�@���T�L����\bV���'����n�2oԮ�� ��4pT��'�� �B�\x�Ja�/St���k�'��u0h�:|hyC��x���C�'��Ƞ�HQ�/V ��Gl��:�'2��G([�4�q�l�d׬9��'UDq���=?Ą�Y�F��Z�P��'o(,j��Q�+��]j�T�' (����� ���� �*4{�	24X"O�\XJZ�|܈����>YH�m"b"O>� �Z�h���▀ 5� *�"O�H�*��|��XC5�	�qh1"O��i�n�o�:�A�o�,X��:"O�!��o�$y�:���J� !d"O���K�mL�r �on8e8�"O��VA�B9����I<1��qV"O�)��Ό�a'�`Q�D&{҉��"O*�(e�ѱ?���9V,�V��Rp"O�D��4E����,[�Y���"Ob�����B>�;Ŭ\�b�n ��"O��㍓�����7O��"O�x�0�E�d�A���e����"O0�9�$.<Rd(:�f_�}6r�� "OFyJO�� �����B� 2��0D"O@��K�<֢i���|�ށ�"O@�r�H�F<��4�N�y�*�)�"Odњ��ȵ|7����6�d�#�"O�<(��F�;qؽP�%W�UhBPSF"O����J�2h� t�ӭ��X"O>�{t�S)3&��q��3L��pE"O2q���eD)QGJ�"0!�]p�"O~��G��<�S$
�IV�hs"OZ��aLT*R?0�QH��vZ�c�"O��8��̊V����'"SL�t�"Oa��F_BD��I��>;�2�"O������Y�uISF�r�R�r�"O���VFqydB�-�`�
 "O�D��#G�sx�Ce�H�N�.li�"O��� �OrtE�)@Jb1�q"O��[���d��CHӳ@ߤ(a�"Ov���b��0崈�L�Q�~�1�"O^� E�����#�����	�g"O�ũ甪s�D-���&�H8Yb"O�hA҂"W0��%
�&[����s"O4����2�PD�%n�7 h�8�"O|L��зc&�,
`V9a�Ph�"O�m�4��\8��:�/�$^�p@�"O�����9\��@��/ۯW�V�"O&u�V��+�r�p5�,��8�"O��X�ʖg^NA��L�Ms��YS"O��"ӈ�$L��=Sm��o\\ZW"O���$�R�dp�!�7��
ܐ�1�"OBl���lT��dd�85�~�AW"O\�Z��ߴ+�,�r��t���"O��te�'d� ����]6W�D,�"O ���O�G�\��U.���"O.���"�5u�93�%B(x�rx�"O��6K�k�� r�2��4�"ONE����;i՞���"�5�$��W"O.<�q�
;y����Y�J� -j2"Or�GWy��S�
O RԊ(
"O����-��0��HZ,I�,�T"O�0ؔ�V1m9�1Z��*ʪ��"O��"l��w���M8B�v)�"O�	P�i��Ĥ2��8.��x"O�yt�>)!����߽	�t��"O2�3>HDmRp�
A> �"O��D�¥sV�]����1y�m��"Ox�R%
&x"b�H�%̇�Ґѡ"O�,2�G]Ǩ�:��k�.ɘ�"Oҍq�,C�xCj\�q�E	f��"O�� 6E�R	>�@1H��$��T�"O� |� �()7���bU16EQr"O�����Y�@�`
 !4ެ�9�"O��2 �7�m��f��Tk$��"O�١��7	��IP�@%hTl���"O:���B>������4aAL�P�"Oҵ�5��9���B��RP$�F"O`t9��՗T�h�7�n@��Ҷ"O̵sB�W}��)f�T�9�-��"O���̀��<�#��L:o,t�&"O��KCϗ5K������
��)��"O�XQ3�7U�P1ـ�� 
� �t"O"���z�dɠ�[=cq&�#�"O����,Õ\)���EĘY�`x�e"OL�i�H*8bĳ��M`����"Oj��E�
M
%���^���(6"OP�⒚=6���g+��iz6I("O��@Vn0l���Lύ=v
Zd"OH4�c�\��:���$��Dn
��"O �g���=B���VZ�+�"O$����ҧc�np�a�=\�2�+v"OR� �PO���"�`B<J��q�"O�aaC�M��t����,:��"Ofl��D-	�j (ڬ38(��"O �C'Ě����:� 	)0:(�V"O��@w�S���!�T@����x�"O|u���8o2��[���D�ȓ"ON�+&!̋4d�hC��9?Qf���"Oj���ؗpl~��.�46iZŐ�"OBq�Eb�r?b�H�헹WR"D�v"O`�	3!
�,_�!qjV>H��"O�qct"%-r�0�`JՓ9-����"O���%�H�0���c��B5�ܰ�"O��&�.5�8!8��83��u"O���l�z0�u�b#ڔY2��"O:���:a�Hc��"b��"O
�ˤ��J;�|BBʶv�6�F"O��Zg]ov�Xf@O5V��Ĳ�"OH]:���IB�s��8ɸT��"O���h�!h��Xs �r��p "OZ=A7&D��F�0o��p(�L�5"O|��0*0=�ekӃ�	�v9x�"Or����YV��S"�I"��Ң"O\h� I�/^LcjRG!� ��"O����O����iA��4����"ONq��·�-i��S��F
M� �"O�#��VB0y��Ɍ�
����"O������ ���.�j��"O t�%N�9gY��R�*��ɩ�"O衚6��IДd�bGI,X�n�� "O��Q&���ˤ#<�"�C"O�3��f�,�Y��"p�:�cs"O�,�����/�V0z�AD�Dj&Er�"O.�����=^�w@8�έ��"O���7��+e^=�E�Ë~��ai�"O�����!��y�
-.hp�"O�PR%�C$�>d����[��r�"O,�b��
h��f�
�Y�T<8a"O�pU�����´���*T�4��"O�����ܡf_�"�-�H�.��"O�� �V���1������H0U"O��C&K���m�u��#6|���V"O���$"�'?�����]/Rm���"O������J�Sɖ7X�10"O�YAD_�h� ȍ�F&���`"O� �q���p�TS� 8'(���"O�qTo�;��ybCoF$IX��"O4�8!�#��<�,�d6� b"O$І���bX���̦`�0�"O�`��'�:T,��3�u��8�g"Or�"V+_4��$��\=��A�F"OtX�ҧ�(?h�}`2Lτq�) �"O�5b���7z���)<D�� �"O��B��.+f�P�"�1Tb�ӕ"O|��X�C��pڥ/k@"�"O�5�4���0���ς�!;R��G"O���K��*^x��[�17Bi2����I?�\	#��i��?���臏��8h�	_�>�.h	�d����	�d�h �G�;���Y7�j-��C���2	�)��eK���dE�բ%�B�� 3�xR��Tp� C�%_Iʨx�#j�iyA���)
+w��4�0#�1ۨ�-�~��'f�QC�$��D-ҧ�u���RBHb��.iT�P&���(Oh�=�'^Ji��JL1j%DX@ҍ3o�vI��I;O��lZ��M���J����i��<�ӧ�U�[P�L�M�|�"������	ey�Ku���G7ju*��)D��J9i/Y�5��Њ�!N8��xa�.���z��**���'f2���Dx�9R2��]����S	Z}6\ɺdo�:5�8��~�RP,x"��`k�L����|����L��ΒY���P�+��\������u�,�ݴ6�	�\�����'W�i�Xݙ�OZQ(���'R�X{� ��0�$ lO����*�'m��u��g�N��jg�>�Դi�`6�5������)�>i�ş�30z�ۤ �ʸ g@�v�d{��`�H����O:��%�B-{��[g����9�p$ǯz���W��&A�P�{��\
3�@�d��J+Q�<�g�N2U�r�:tʚ�ob0TCG�y�� 㕬��S�|�����qGt�:�b�YGxB�
�v����L�Lr���>g6���p���-��O���"��>jq���Ш<�T��A�#�&��������T���Ç9�����D�;q"�O��n=�M�*O�e�������Dm�6h�"}�4m� �V��@�����,��ʝ�~X�H�K�4���5�^���U��!Ң<�� RMX/`�b2Z�*w��<�`�8!((I�U6p�ȁ±h/R^ j�b
=�,��N� �\q*�FɾNhtH�	�?�4�i�:�ɁDp2���lQ�a�Yٗ��W������	A�S�'��<@w�����%��� \v"����>94��,Ω� �	3be􇆳.�*��i�$f�.x�������WyR�O�D�i>�ɸ�$SBbU�^�%s��!�'���0Z���qi:��l+��)��	�6�����)I�L�X�����h���/��'w��pu�$~�0�O]� Ћvb�
Y�0
����X�J�>�FH�K����|�$�xbO���?9��i���\�h�"��d�( �G�����X���D�O�㟄%�xPE*�@��4��YX�4��=O�in��M�M<Q�+\���ؑ !-�V����_G��7��O�ʓM㎩2�'�HO֕�3
2���1���J5��(!G�5!�����ӗj9>���O��4�Xr��;_!�!�7�W�x�@�ɡF��O#����Ec�u���Z�*n ��C�fR1�.Y����@M�2t1��
u�ƹ83�Z�6m��I�	�p/���)�<��4:d�8�v�+x�\ 
�V��ء�T�(��I$�����:d��'�[��O67OԦ�&�P cc�?��'�����%f]�񳦏�#@P�=��'�arg��\   ��   Y  $  h  �  },  d7  ZB  lM  1X  c  �m  �v  ��  ΋  7�  ՘  �  `�  ��  �  '�  h�  ��  ��  8�  ��  �  P�  ��  ��  v�  9�  � 	 q � � :% 0, 3 X9 �? �@  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��nS�R�p�<��4�O|�OR�Nȇ|2N����!�YBB�	n���	� j�I j-S�T '��R��'Ē�	%�'�����V=M$NQE)K;:��	�'�1Or��@�'�M��|�c�<��8��jӹv������>D��B.ك�I`A�2"��8�f�|���ۦ����'>�X �s�t�JWA�+:~�㠃6D�$3��O��yA���_Bb}�'H2�	w؞�j'b,�H?�Zaά<����S�?�l��!��
���s�B�I�!��unáZ.E;�_2ob�C�ɨ%2��h5/�9��A���37���>�r��+KЂ;g�`Z��g�<�b�^�h0ک���Оz��@��$OZ�<)����}��!Jf��f�آ�XS�<A1�Ǿ'o�k���&�0u��Sk�<i��۟N�p ��'�0)<̽*��.�hO?牂~�lmx��&s�R�A��U�p	�)���V1O^�?9�I�f�Y3Q�ԉA"&T��e���C���$8�O�)!���(?z&̺Qd��ba���>�ش*'�|R���T!P �7f�8\���H?��<��d�!W��r�ʔ�Q�dM��,_W� G�4�#=K�1���2�x����(O�=�π P1��Z#D�d� GO�  2��b5O��	y��hO��
$ J���M (���"O�@��žs�j�;Uɔ!�f���'Q�[���3�Y������`�{=ب[aI<�$����剰b��Qp�ղ���p��$F{l�=����؟�!�ȩ������Z#(@���&&��y���R��p�#��a�<��FЫCx�?I���ܺ'���a��`1����GQ�HR�)�.�1�F&Ƥv`�`R-��DS]`���>O�t�v;�`##$�v�P"��xb�'t��^�=� ⢍ό �nL
�C����D{����:�, ���xPT(�.ZW�ay"-M�Q�2�6r�H� ƎE�	ZY�';��%�)�'c�̉y��=9�J��0��
Z��-�ȓ=��p릈\�(�И�&�YE�=A�np`9�F�R����(ςY*�$��� ��E.@�� ��� MP&����=�۴#*7�ٟu�&}�3��J�᪐l�&r��u�ēz
����Pp�씈F�����\�'��ac*χ�͓��+���	�'�r�@�ϋP��1�6bN}�U��'�v �Q(�vϾ��1
)�y��4:ʓ��)��`��(�d��7=ʙ(Šz��y�jL��&7��L�BG� ��ٔ�x�'��� O`ӐY�",�X�gU�_���Ǔ�OA�r랖.ibu�����e�a�'��O�pr �ܛL0l���p��Q"Ou�Y�Y�>���ǾO��
�"O,)��H"f}-��L� Y3*Qy�"O6�\59�̑��j�!�(=���I$�0<!!%�.C�"���|���i��Ub�<�$G�N��A�eŐ	jj���#D^�<I$�=t��c�ʛ�H��hAe �[�� �>��/��N����wT�G �Z��Q�<g!	�B*�RǦV�Mw�b�"O�<�0C��0�rܘ��P2$�x@7�K�<��h�!Of�eѢ�6�FA���	E�'�ay��U�^��u�֡L��H�"���y�.�x�\I�DG�(�����M��'!,�i	������*V2���'��U�0H����(���//m����'���3��{>d⠏T�$՚t��{b�)�	�2۠�1QC˼�@���d�!�$�(��j�"��7�<�$�.�!�Dċ�8��UhO�����H	,�!�V�7�]���ZXK`�Ae�.G7��
O�T����+�0h�d"
�K!���"Od��$f,m�l��g
4,�)��"O�k�:�Ψ�1,@J��@F�D$�S�'c�a�ƪ 1�lp*0IH�&�؄�Y�
A�Ʉ�d��h���	":"���J�h����6ƚ5�֧�=TN@x��2t��`�����qZQ��r�<����D<� HQ$:�YB� ��(�FŇȓJ�0	�UE\�A�B�7t����3�pt;�Γ�wiĔei��~�z��ȓE�H�Ij!��!1׮(8���Q���$��:-&�5��;��ц�}���bêȚꬱ�!�Z/t�І�f�.z�*��W��R��.�,ņȓR�|\���H�&�(�X�'A?T���0.���šG� |L)1��J����so:�X�h M��x��ͯ{ș�ȓ	�~��f�0 ~`��@�ˡ&�]��S�? α{p�RY^�H3BG�0j`Cc"Ot�"�G�>sW��C�G
#U0Z�;""Oz�{�A�	�١B�G*Z�H�"O"=Z��!<�`�P�W�XJ�	B"O2\�G�*仄E��7Z��[�"Oh�W�B(|$b�e[4Z2�}[5"O�ذq��]Z��B���+4 H��"O��Pg��=�l��).�`�"O�t+�'��t�g"�=�AC`"O��څ��?k�����]�$���'"O��P�K� ��ԓ㎌H*T�1�"O�ɀ"G�+Jܘ�RGn���"OB�wM���^�4���p<l�#"Ovu�'ĺ-�� $�O4L4����"O��âJ20%F���+MC�mX�"O��vaהh���q�$/f5�"O�m�dÅ�-����e`h��"Oԭ1s.	�8J>`�EF:�-`T"O�E)2cџ*f<�;P�
9v�bJ�"O�%��>c���L)R"O�D�r�]!�"3�w�$�D"O&�SD�N]Vtx���Ҁ:��q"�"Ob�+�v����,��2��4�"ONH��HJ+��]��2_�м��"Oyb�N����p��0$��ܫE"O��ѡ��:��x��]KL�D�6"O�(X�B w�
5qBa-V8ڜ��"O�鲳@T2fLn\s7�׼?����F"Oȵ��ڇ4B��ϓL��Th�"O����ɏU��xY��@c���"O�TY7 \%*�T���B�\3�"�"Oʈ�G�5.����P���'�Vbu"ObՂ�,..�Yskπ1���"O�����P�?0ҍ����6EP�"O�MP �=G��aAPBE18�0�"O�$
��Ê�ʔy �͓Z��(a"O�$*to%E'L�[b`�\h8qXG"O��q,E�4�\*0 #=4��S�"O8��1�@�7#��:���(H�����"O�ŋ�!�^�4��N?q��u"Oh�@0Jʊa���`�o�� Ǿ��V"O�!��LZ��i��2-I "O�U�g7��� �[�B���"O0� �&�$ꀔ���/Xr���"O �+��Sm��-��&Lz66)@�"Ony2ק����K�ۘ9�Dv"Ox@`���Cn�ęa��]����'"OȰ**@�
�`�ԧփ*}��j"Op%��EG7v �e��nv��b"ON(�C��t \�#�D'>`P�"O�(Z�G�*T ����c��d�$�"O4�FYs��4A�)Z�\�r"O��C�lH�f%K��Һ0�Uqf"Ofĳ����$�h�=4�H<�"O�IcQ m��ي�홸��%cP"O ���a�+@u:��A͓����e"O��R�cD-N�����T�I���&"O�4�E�|A�b<B.��"O����7�F�j�U7zOP�Z�"OB*�!��3�^	��؈ljA04"O��X&����Ѫ�F�*'J!9"O��1�'�()���8� Y�E�H�`"O<T˰�ƍE��KdE�$|��ܒ�"O�H"�وP�)�Ĥ����k�"O� 
��.C!�e�w$�?~Y�P"O�D��H� @r�I$��br 8"�"O(�)�N.xa��r�=rm
 Ʉ"O��g(�����F�0OV��"O ��#V�n���@�qWFЁ��'-�'�"�'��'��'o��'r�P{6n4-��V�}i(P�'���'�B�'I��'Q��'X�'���)w[8�	��~i@9S��'���'"�'J��'��'2�'�Z9 ��K�P<x��
3?r��'H�'���'m��'���'T��'$-�'�N��eYq��@��u�'f2�'�2�'�b�'���' 2�'G�y�2$�0���t���'$��'���'���'4��']��'�Eҁj	)0�[��TѦiq��'�2�'�'���' ��'���'���ҍm�rEK�G��f��$�'�b�'V��'�2�'��'���'ՎM���B�_��`�WC̪�4�f�'���'�r�'�'&2�'���'ڬM��/I�P�T�#K��/������'���'�B�'B�'�r�'�2�'��yB`�����8₋���u�'I"�'B�'���')r�'��'G��a�&�4�\
D�α4`(��'w��'b�'�"�'�"�'b�'y�|@'����HT�LҌ[E�'��'n��'���'(�*`����O��h�KO�X�8�K��7-�9�EOy��'3�)�3?Yc�is�H+��Ǵ=�X���<.��;5$Ƞ�������?��<�i>��a�bI=�����<	��J�~�z�DIm��41Ù�\XҪ�F� eQr�~j' ܬf.��ѯ�8+���AϘW̓�?�)O��}��G�!^�X��8/Of�G�e5�ƈT��'���=mz�i1���2^�F�D��XK% ���M�W�i"�D�>�|B'���p��̓&n� �KD�6���@�!Hni�g���P���L��4�L��N8n�4��W�V�N��c��&Z.�d�<YL>i¿i��1�y�o",l��k���,n(���dK���O���'��6˦�����ޚ;��l!�)��֠�xR�%9G��q���
wɟ�H#Fc>U[���KrF��	.�XPp�&ԛ.�S��Nz���'n�	ٟ"~�x{0A����W��E;�FI�,n�ϓb���i֯���YѦ�?ͧpǖQ3ūH(D�Z����\�~���3����t�\��!_�[��hs�B;q����Z5a��
�2b,�$&��%�$���d�'r�'���'ҕ����4
��!S��{��$�T�p�ش~F���?1����<9���}|DI d��0DC��,��	9�Mմi{�O��韊��������1؂ ��#ݕ�L�*I��(3+O�]��C
�(��?��<�G%��}�	9�o�2t"�ݫfI�3�?y��?���?�'��$Pڦ���ix��.\|� �ۀ50d)���$wx��I��M#�"i�>Q�iR�7�צE�'�S7m[�A����9������[���۶g�x���	�i/¡�F��6n(�!��?��;o���BZ̑@�&�5J��aA��y��'*r�'Vb�'"��D�t.qô l]� ԋG�d�|���?a��h��������ڦI'��8���.'�`A"��"�4hq�G��x�6Hj��)ZH�4	>O4���dq�ZE�o�fq�f�I�R��E��~���iUO%��<Y��?q��?A��Y<,�8�.��b8��2b����?����BӦ-Jf���	�(�O�Z���A�ay�-�R�E��1OB~bD�>��i"7C�i>���E���R� G!*G!��ZD�͵Vg<�i@#DyB�Oo��f��4��'���� �N7C��\���*�W�'J��'5����Ox�ɽ�M[�M�0�ґ02C
-t	�=���J�q�����?�v�i:�O�%�'�7-��G�꤫�Kϐm�څ3��5��5m�џ`:EKXp�v�I��<I׫ �z�;��[ty�
ۮhʄ����Y�"�)ƀ���y�\��	П��	����x�O/X�5�N�F����'�H%b��h�n��e2O���OH�������"�`@,?���7ϐ#{5�@Jb�Φ��4a�����O@�,O�"%��'*X��%k��`��(�B�'m�P[�'�f��M3Q�|�W��I؟��*�"�L�wت7��e+T�Aş �	����Ibyb�a���k�<O��OCqAVu�#A�>�q��/�I���Kæ�+ߴ\��'ڮ�B���=h��]�A�
~�<T�'b)�tNT\: /�)<B�I�?�#����l�I� ��p*ǂ��jv�Q��S"6��<�I�� �Iԟ��	I�Of��C��l��j�*#~@ ���0%Ҫo��I�5��O|�DBȦ��?�;Z�t����5
R��熀�$�A�1��6!kӖ����ҡ0OV�d�V2f���BV�P�բ�n�+���+ҡ��Unx���e;���<���?����?����?�0�Q/���
��l'ސ��@�,����ʦ�;�'�şt��̟��.A�� �ƌ�v Lb�g�=bڈDѩO<�nڴ�M��';�O����'�x\S��[@�X�d)N~�5j�lO=$uTܘQ�iV�X��`�a�jJP��My���w���4�B����,A!F�'G��'��O�剧�M��]�<��B�=����JG\��Pǘ�<�A�i���|R@�>��iUh6�ʦ�割a��@$d:\(u�ע%Ȋ��PJ؃�y��'�xm��g�ẘ�	gY�p���� @���a^/#O��`$A*��p�44O����O��d�O��$�Ot�? �]#��8�m��%Y�&���|�Iȟ	�44����'�?���iD�V�d�Ơ7jL ��bYZ}�d@�d��<��O�oڝ�M��0H�a��<���P�H�U`V2�B�b�g�(;��
Ɖ�"K��J)�����O����O���D�"U�@�M�Qá6fH�d�O@˓]��F@'y�r�'R�^>� �CJ5G�Z�⇀��5R(�7?�$\�(��46��v=O��<��W�]m~Ly6ׇ�T]�qO
0%͆e�P���
j`�Ug�<���v��ș��E��������
I�^��'%������?Y��?��Ş����9:��	��d�	�Q
@甉S��3-���$�D}b�r��qudK�\( Z"bM�iu��%�ӦP�4;��9P�gZ�<I��?jR�h媃�6{@Ց,O<��4o�O[6��� ��\i<���:O���?����?q��?a�����ս�( c�h�W�x��H)���n`X�'N���4�'yf6=�=��A
f�@f���92�\�a�צIa۴�y�U���?��I;h��\��C��!ڷ�|�c��Sڞ��ס
�s���ۼar�j&*+1
�O���?���F���ѣ(K ��B'�(D�u����?y���?�.O�o�? �J��	��p�I�GL��ICMDuv`a��T�qk"���X���d�Φ��4�y�]���̊�6��(��)b1JGGx���	y����:w�L��'��#[�s���1��'���i�!��@ ڼl�^�P��'�R�'��'��>��ɗVq�C&�?vm˒K��~��H�	��M����C~fr�~�������v��j͢�2ä�s
�	:�M�f�i��6�Ҋ��8@d;O��QnЮY(Q�D�}R��S��͞��5��H1VI%�<���<9���?1���?��?�Ʌ	OQ"mI��ȏQ��+�������2f~�T��䟴��H��'|�&cƞ7�iq�
yx��5�>��i��7m�s�i>����?�����"t�k߹w @�Вf�Ba���^ayr�O�^��=�Iǣz�'�剺h�,}�`��|�������,O$�������	韈�i>Y�'�n7M؂��>h�Œ�ၟyg��g��|���1�?�[�(c�4ZC��&kӊqe�^8 �Rh�e�`� 1'&.�2�B5O����XN�ȫge޹�b��:��;Ȭ��"Ȇ!#4�eѥ��S8@���?��?���?����O���K�f�TaZ2n�C�*ћ'�r�'��7-N�w�I1�M�M>q��̮E�:��+�A$�ƅ��~��'�6Ŧy�S�(��|��{�d�I�D�q�Ǯժ=O~���H7�8�*�)k�����N�Iiy��'���'��o~f����z������Y���'��I:�M�v���<����?����RE 
�3}؀�2�� 7`B�K���N~�>IԱi�6��_�i>��S�An6�	��]��(R%�*x6T��D7 0�Q�̜Dy"�O��X�Ň�.s��'�r�rF�]80B8M9�@,o
�9K��'�r�'�b���O��	'�M�aR�I��a��i�����sv��UG��';`7�9�	��dܦ��vK�v�x�K�2KH����\,�Mk�i��W���y��'�|�;s�9� �(�R�H��Ѐ�f=3�ҽh�x�B�l|��'�2�'_B�'�2�'�����%(W��B���_�l�(�4R���Γ�?	����<���y��9hA�I��)�� h(9E��};�7-@�!RK<�'���'ta[FJ��<1��� u�4T���}bPQ�o��U�m��P�HE Տ�6J"�E��˓�?!��`ȰUi!h� [������^���s���?����?�/O�$oZj�������ZiH��&Q �	S�#��_D,8�?iX���ܴ ��-9��0p����fL� F�޸*B�(?z��O,	��jY�P4��j��<	�'8��Q:6ʏ'�?��c5#�	h5L"�rE��a���?���?���?1��9���`B MD"-�$�ԍ,���2��O$,oZ�e��n��F�4�*-���3b�X��#�)��]ۄ3O�o��MW�i'�lCLY�y��'�J��'_3L��I�3戩Jb�@�P�7
]���"X���'\���������t�	����$}�1�흧v yg#��:��ݕ'�L7�;�P��O��d3�)�Oz��eh��6_�2С�-�n�*�@t}�izӪ-oZ�<�N|���?!��E�S�vm:�	�
 -��#bU[+�)�����W�u��!$��]��O��G��RgE�M�Xa{cb��|�JP+��?���?���|.O$�m��X1�1���G��j7�Q�"�\L:U#����i�oZx��R���4�Mc��i�⌆DP���B�6���Ҡ�(�|�7 H��y��'xJ,`BcxV�h��W� �ӳ�5�ķ!� 8� �ǃ�)�`$��'
��'>��'�2�'a��9�ơ�_�bq��/J5O6Dy;+�OV�$�Oxn��oh��8ٴ��q��#�o,� bbȑK56<ۙ'8�	��Msg�i	�D�>V�X��'� N_�6�5�D�h/��kP���ʂ13�dU_���J��Ţ<6�L	R�U(!~Q%�ȭZv|j�A̟6�6U��aPK|(4K�Ǟ�:����&B�4C��AO�b�p+@JeH]fKU/�p�7ױ�Ov��b�Ȭ ���ق�ʫ7و<��N�,�2�-�(԰���J7t�\�k�K*-��!��N#&�¤�&O�8��=�.�A�DX��R1����HӸ���cC����"c����Q(�$)�@�Y'$�hqXqJֲ��R�@5(�:xrMN�M�(k��L�25�*���G-HP�:f�i#��'�B�O?j���?2�8�񷤒 o��ͽ>Y��?���c%Ԙ����bP%�6E{xu;�CB�S}�(���	���'��%޻�6m�O���O�����d���^�? 8��-�6�����J����@^�l��;ajT��ǟ ���T�~26%1M� JN-{p| �v����=p��B�V@�I͟|���?u#�O|�a��9W��6-�����ʝ0g���A�'>H�'��	y�'�?iU�M�|�����&4��冘�x�V�'>��'�Y�`�>�)O��D����ca!.r%��D9G��R���&���<���D�<�OXb�'yra��*=��B�%�F��$��qT�7M�O�p�gDH}�U���IFy���5v���\�zm��?
@��� �����ш'��d�O��d�O��$�O��35�[��?ȸӴ���N �l߳9b��dy�'`��䟀�I��p��!ʡy�rQ!�]=<�I���Y~���?Y��?������bp��'(�R�*�N�7|��
� )�lZHy��'C�	ȟ��Iڟ\��$k��x�Z��Z�
�Z�*��n���D�O��d�O�ʓ7�(df[?�IZ��%�@��0��dM38\2$��4�?�(O���OR����V���9}��A18�	���)6�LM0�cnZݟd��iy�������?�����"&LP��zR��%V��)u��M���ӟ��	��S�)b�0�IIy�ٟ@����ޤ� ��ԉ:�����iv剴("T\�ٴq��̟�����ܲm4��KO�EW��ya��1ٛ�]��j�d+�S�YWBX�㎟1C5�aH5K-RQo�<���(�4�?����?1�'yƉ'�b�J$W��!i��Xs*g@Ag�7�P�F-�"|
��ڼ�������2��ū�"l�5�i�r�'e�F%r�O����O��	?	O�WD�7�my��N�b����.��ğ��	��8D�N3J�zBa݇]l8Z ���M���{%"������O�Ok�� q��"[$+������W��Ɏ=c����ǟ��	Oy"n"Nּ�/�*JLJ$i�$x@5��+��O���'�$�<Q��F�u�A�$\%��d0�FY-&��9�<���?Y����D�'�H��'|��U1��2\��u���9Y(BO���;�$�<yfc}�IU9�fE�ǂ܆!�l�C��QByb�'SR�'�I	I���J|
ǢC�%v�4�N�uA��B'꛶�'��'5�	m��b�|�&���d�����G�KS��˱�`�v���O^˓Ko�XSǓ�d�'��$�G9c�:��d�89P���q�BOʓ7(`�Gx���e��D�A, �I�� Х��i��ɦH�f�ٴu�������D��q���%]�z�P�zg�	�w��&^���wb:�S���+��Р;R�Q#D�
s��nC�J� �4�?����?!��~��'YB��p4��2��[�N}�3Nħ4g�6�
w2�"|���D������tl\ �Vj�+xw(�;��i���'�B�C�{��O����O�Il2.�à�]�n�N ��)NAxb��0A#4�	��h��ߟ̸�CG"�v�a��1}�j���#��M����Ha��xB�'�|Zc3~���gìi(t�ӟ5К�˨OD<0����O��D�O�ʓjۆ����*}�>���$�
�.Eʳ�/[��'5��'��'4�	�f��c@�XΌ��$"K2T�h�c��(�	����؟ė'=���A�}>ys�
#\����~�4���>���?1M>�/O4 �rY�DR�W�[`�PKS�:44I��>����?�����䕛�d&>u�e��Mnl+#V�LU��9�ƌ�MS������Bq��O�]��9���� Hƕh�xp� �i��'�	0Tf�}L|����(�<y�b��
dv��皕��'=��3e��#<�O�R���L�`�xx�R�S-02�`�4��D@�$�m����O��IX~�/�:�såY0{�2���MK(O8�s �)���(E�!m�+]�n8��JǛ,��7�Z:*<�m�埰��Ꞔ�����?	1hRj����)�h��,��yޛ�M�)�O>��I&CwN����%s�`�P! z-���޴�?����?!��pܱOH���豕�=Wj>]"�ΔM�@����=�	�Y��c����Ο��	"S��P�gI)0"��P#	]!i>�d�۴�?	��Ԕti�O�$9���T ����y��t��Z�B��TJ�W���Ƌ/�I��\�	���'` �!�o�2T�ؤ͒6LZ-�X�D3 b���D�ISy��Y<-��Qq���`�b��
Sj{RQ �yr�'SB�'F剃P��MR�O&����@=_"��ՠ��Q1��[O<���������vh��OtAR%��,V�37���?���?�)O��T.�jⓆr���#�ȍ�`�(���B*:0pٴ�?�����<�% t��O�e�Ӆ����!u���Ei<���i%"�'���0G�U�J|J�����%ݳW]��Sց�Tshh��DU�y��Z���'�J�hϟ�i>7�OE]r0r/�cq8��m�g��X��A2h���M�&Q?5�I�?���O$d� �#֐8a�f (N�L52�i�ɫc�#<�~:D��8!B����9;|њBæ��ֈE$�M����?	���ҟx2�'��L�`�D���U�+J�y�~�B̨C�)§�?�$�\�^f��d�0K`mT9�=0���O*���;�X�'�\�	�0�S�? $�0��G�c�	f�Q;����h�1O��d�O
��/;� �I�+�/��З�0F��qo����34����ē�?�����s��ι,�!#%)�;�P�"tap}�����'i2�'��Z�H�Ƈ�y�L�)5-T�����	�♋O<��?1N>	(O�x�˖�jl�Y��?X�B<Y��J��1O���O���<)d�Y^��)�}4�s��7�r� d�͇9���⟼�	h�byBL�3���H�-��黲���_��Ia4�I9���ݟ������'�ā�p�3��K�`���i@�~VTa�RN��<�n����$�|�'t���}��G�nq��Z(o�� 2�,H�Mk��?-O�[R�c�៴��G5�՛����_�X�K�m��4�L<�,O�����~R��(Z�c��& �\a�G	�ͦ9�'���Ef{�R��O���O���=����d��J��aaGH�Tn^�lpy�j\��O����1�
�"��9�q�/f�DYs��i��T�@.v����O���X��>9���;Vǌ� S$ ��Ȩ�I؛vO�*�O>��	�c1�rE�	�T���%�?^Z ���4�?1���?ٗ�[���O��䡟�;&S8�����b^*BX(�7�'�ɪ>�c�<�	��$�I�L�ȃ����(IGզ5�ux�4�?����A
�'���'�ɧ5�"���qx"�B*p6��ëՅ���D�Qd1O���O��D�<�ק��Lr��RՈm�1�f;�顶�x��'MB�|�S�̩�
թoZF�Q��0^��R���=��c���	�����xyB��H^�����I��Qk�<�:u�W�[�2��?9���䓥����������"9<y��-װP����?����?�.O�訂$Zg⓼jΆ���ߧ2R��W�� FAD��޴�?�M>Y-O��3��dQ�%y��;g2x�6!I��N2ћ�'�_�#� �(��'�?9��5y� x���`�D��э׏j��IS�x�S�$�ǫ(�S�D��_I�!�aB�r�r�xB�	�M�(O�ź@�Ӧ����$���<�'�F`�:Kt֔(w`��$�6|rش���^C�b?�!���3)s��hC)[/@E��a��XK�P����IП���?��O<A��-����U�:s��*�,S��pj��i\x:v�4�1O\�dS	;���j�I!a%Kw6B�~1lɟ8�I�P�$ ڑ��'5b�'%d��P�ƎAސD� C�$k3�lhSc?�ɢl����I��|�Iܟ��IǟбA�Q�Bxq"@�/_+�F��M��lE��#қx��'�B�'��i����, R(�A��5�`�J�>�.CP��?q��?�-O���F�;�N�:C
�4� p2�mƵ:b$�'�X��ԟ��Iyr�'S"Ǚ�bOf�0�M,���(ӫ"��T�y��'���'�+l)�(a�O-�H����F!$���F�TK<A��?1*O�$�O|��T?�AWc�o}�uK��0�$X�� �>i���?�����$N�-d�$>�XGޤX&��m4�<���M-�M������	�O�}���D#�01�/�4GU��y��i���'��5\$�L|R��ičNbX�X��܅!��ݪ�Ć�[�'BB�'�d����'/�'*�	�?�Usƫ��?"��J�0Z��Q��U�F$�MۡU?)���?�y�O�X�^����E-I�+�����i r�'�.��b�' �'�q���h�͏�}גi10�ӯp�T�B�it0�Q�zӈ��O���z]'�t�Il�T9򵯑�b�ʥ�Ǩ�~�ȑ�4ꮵ�����S�Ow���3q��a��KP��#t�XrbJ6M�O~�$�O�(�N�I��?Y�'$����̦n�"�ʧiчx�8��ش���6�S���'��'t���D�%�N��$\
m�
bӖ���Vp��>������c�FH�=c�<82�[1L �:��e}�L��yRQ����8�	Ey�M�o����oC�rwϕG����q�(��Oj��0�$�Oh�d�;C�~�a`�#��] ��/t��!9O,˓�?	��?�,O@�a�(��|�%����>�~�뗏ש��O*�=���O(�$�Rs^���_<��a�L�r4ɦкd�����䟔�'�L���) �ɋ'M8l��i�*["t�%k�u�mڟ�$���Iڟt��)ğ0�O�4wf�W�|����{��ѻi���'1�I�>� ! K|�����w��� /��1�K�r��/0���xR�'��E�
U@r�|���%�󂔇1���@�)U.sG���i剐$-h!ڴn��؟�������t6��&���T.�$��f����'����|��IS$$:~�"�*ܮ �d$��כ&�ݎV�^7��O���O\�)k��ǟ<�a��3�|l��RX��0�߅�M���?YH>E��'�0̚�B��U�`^�y�|��ux���$�O��D�>�'���̟|��*1ęXk�V�X�;1��q�lZy�I2A�$�1H|Z���?Q��q&�4�p�$ c۶��.~H��q�i�Íf#�O,���Od�Ok�D�Y� ��q�K�61�� �3��F�I`yB�'r�'���;f6V�ӓ*�+z����F*�hݻ7�Ă���?������?���>�� ִa��_̎<xg�Q���`@��?�-O\���Oh�d�<���	r���R�OY.e�wm��3�PA0�NM<4͉'r�|��'�B��Gk�)�7�X���r3�1aV�Zt`t��?i��?	+On)i�n��Ӱ^q�wƖ�ZY�M�d��c\`��ݴ�?QH>y��?�d
�?�?)L�@��Ŧ��]s�L�u-����Z�u*���SlШ�@5�$$�}����g��7�.�rQ�Q�[v�I�P�a�X��CW47���0����Ov��VJ)D�����W~��W��-4=3���3�­;u�_�y"���!7FP���߽Yc���F�%&)Z������'���84���o���'�h��|��o��ywTxu	߾W
����K�E�9y�Ɔ�[�ؽd"�D�,�U한l_��c�ͦn(8T	d�Q�~'LLbV��:�C�E͚|�}
�0gnݱ�(��������@��2�u�)*"�F�ܭsU^U`1�˨a�b�Q�i��	�&iD#
!&��Č3�:=@�}�':O�m{G.U5	��ٴ�U�Q�D"6-^&@��2��A~S�q�1�H�m�r�
��l�$�K�d��;fJj���)�r9d��DfÑ�>���|2�Ñ�?�}&� ���'e��b��s.~T0%,D�{ �
+�@���� =`j��g����HO�I ��#�B���F�x�S�ΘL��x�̪ k���OR��Ov��O�4�����_��B��C�mYh1"�����ɈqOރC[�Qٷ ��8)��)S��(O���Q�����h��8]G�p#�:H�2d!`�P�al|<�v��H�+��(O0�P���c"$� �ePʸ���A�#�� bӔ�n�ԟ\�'B��bd�U�be�$ȑ��c�+a|"�|���&�@�U%�Dl8bǄ���'p�8r�'i�	/i���^w}��'x�tc�ˆ+o���J؟
�J���'�b$ǿ&�"�'9�)N0Y"r@Za��8����&��<�<XBwj�8�x��{!z �k�D�D-����9q��I�
�BG��`����Dn���3�ҧn����Ɵ~��)����*����D�Y�B�?�dPQ�����K�#� pDo[9�!�䐙@9��^��I����haFxb�i>���4v�2�ؠnp��R��C�g]`jO>�w��j\�F�'�]>������H2�#e�|�"� ��D-ε{t�[˟��	�{{�9��X(w�b�(�ᔯWĖV&�pB��O�Z��b�Lt�vM�qCӉu'��J��C��)���R'�_E|��i��>Y��CR�?5Q���\]�wOm-����.}¯��?�ҳi�L�0�����2ă�Rh	���D<�d����OP����*G=<`2�@�;K\ ��=.ax�,�M���S`��"�}k��Ї=���[Ÿi b�'��OO�^�z�'��'�"�w���B�1r���I�X0f��sB�#|L#��V9�AhA�991��aPfF"�yb�A=_&$�Yw���d!�}��Ζ�4���6��ee���u�>���
���	ND��=̓�nH��F.8#2�x��
�f���c�|�i
��?�}&��"2�VPz�= �B�3w>�YĢ:D�$�7�փrT���C@t�
Ecy�$�� �HO�*���<�>ȑ�ŝ$�|�#5��d�/�d�R���OT���O
̭;�?a����$t�H&�K�YP��g�ۓ{�6Pb�'^z�B#떸6���T�خU�nM�Á�9�xRk�8,��L8�����6`Xe�(ן����x�(� W�t�z���p�r��)���$LE�EC0)���I$k���<YF�d=���lZϟ��	!(i�]�$��c���hPƋ�2D-��џL���͟`���|��"�=Y�b\�aG��1@��?j��a!�f<��'��5�� s�Z�.y��<�`a ���;W�@�%��ӑ#V�8��t���wێ���_�6(���g]�L�f�<��i�П��L<�����jޏ3nع��^�A�B�ɃI����d�^@D����$��#<A��4��m��*|t��0�X4Q%L����`%�P��̐!�MK��?�/�@��� �O�e��ϊC=��#�8�Խ��!�O<���
��3h�yX�����vH�U�0mR�0��˧G�&l$�W�D�,�R��~1�O6�k�� ���N���D+�*V>g$���?5���M�SĚ-r�2�8�'?}���;�?�P�|���&R� �v��˲ktNQYW�M�y2��_ U+�M�6e���3,�*Uў���HO�0H@�=u;�c����U�Q*��Mæ������Γ0�)�3˟��I����iޙ�pOP� �@��A����u�D�&��1h�@8w~Q��(Z5WȜ�|�bV�8打X���{��$���(d�_�W)����Ɂ�>X��c�av�z%C3�ڽ�B?O�I���)�ظC`N�t����t��|���|�$�{&D��V�	^��[�@� �y2��G�n���!�z�L5A����y��'�<#=�'��k`�PC���G� �΢N[J,@�fq�Hs���?����?�S��
�d�On瓑J#�5�V`�'y�tUj��1�܁�K6�(��)s{��C@^�^�����/=ŨB�I(q{ҵ:bL�5SD����[�n1YT��Oj]��)� ���d	Y�E�<�#���q<$�['"O4�¢�7[o�R�Ҙj)l{�Dg�U=tq�ӹi4r0O�	�1̈M����a�����'��@
���'��逑�M;�e�;6M��x'jZ'tD.���� vv��q7��6q�V�&܇ϲ���Ɋ}}�4Ԥ�EŘ\ja ؚ-��d"tAޙf�`0���=]�*P8�k�ux8���I�Q�@�����]�ش�?ѲL$M&�P���٧ Y��JFh�4���OB�"|���'\f <���
F�� �@�\�'�ў�S��MC(�2����կ'e4)ZeLE��?�(O�16�����ޟĕOd��"�'�0X��i���8b�m�)Y�=P��'���C8`���'֞��X����*�z�k�JݑX�S	1��M�!n��d���@�iG4j�'�����$^�E�@� X��	���`"^U�� !a�Du�fİh{d�kA���	�c���$�J�)��<mF�9!,6Y%D]cB	�k`*B��<+XN�p��`)@�A�`�
Ƣ=�',ؑ����/^�n�ܽ���C�u�0ݰ�j��M���?��f�c��T=�?)���?Q�ӼS��R,[vʸc0iN
r���·��Q����3/�2p��o��y(�\X��ĩҚCA2�͓X��Aǭ�Gr���/O�M�fG�Ly��
z��:�4��O�,K�d��<Y��i���)R��Z��5��)M��'��5��S�g�ɒ-�z��[%�"`���>A��B�I�	R�YR# �(tҁ��=�^�	�|s��4�B�O�p����5�攋%gY�pmh$ӣ�9�@�I�O��d�OZ���Ӻ����?��O��<:G�β]��+��,46�U�{}ޔ�D%�' �`Q%޼f@<eD�r�'Sޜ��WXĺU@�o�eN�B�a�+�F}�&�_�f�
�C�c�;#���YL�'ؐ�p�W�@��Y�)@�,�BPk�I�?	��'x�RQM>�9�M�&Wބ�s��� ��e���,2���HH�1�<��i�'�:`�`.n����O!`�ŝ>=W^�i�匃�dX��O��d��KZ���O �S�
;�Y �ニ%��6��6�V4��?>"j$�Id1�Qi��Ʈ9a���?�(>&�kDMEE^J�Х�58��� WUg��y�fJw��͙fNJ�l`�	P� Ă]t�HL>i� �ß�AL<	Q���*��h�עM�A�h��Z\�<i�ƜB�taZ7��'V�H���Y�'�ў擔�M+̈�348���i�(�
M�� M>�aASL���'{2^>��aA�러�� ��+`�@��ϳa:��� )Cȟ(�ɅW�&���Ӧ:�2XmZ*2�
Ө��]����/��3�E�!�"@3��P�b]���>��b��.	�U��J��a�"[_/"����P�q;¼3\w3Z0p�OХq
�iۼ0����R�>q����kI>�JF+X���� A�U^�J@�_�<��*
D�([bm�"v؁��Ņ�hO�i�n�'vVHy�.N� �b@:U�>H��� �Fe�����O���N��}A���O ���O��4�8Q�l�2"Pk��܉B��1��G�\����O���3�ԜOQ1��'��;���#��,؉Qpf2t��#��}���u��`F�/¸O��<�0+��<)�Ē�*����� r��`(�a߲+M�'��`�S�g�z��x�����d��PA�62ǖC�	�]� 1$��w+�`�^n+n�h��"|��
�^H���q�	�sF�!%KI&�������?����?!�������?9����<:3C�8]��,:�a�
���`�#{V=�/�"tn�Q+�ђMџ�p��ޫW3�Y:��Z�?�(�3�ß�Tk$릅�X�.>�Q�4h�?��O�q�R�
8lzL�qdH�Z���	���a\B�g�2l��'�Z���'�$��靓w$�(����c,�=X�'�~�(��,��M�f��bEh�՟|�nx��]l�]yRF�U܄7�O����]<����kϝX<�D�J(�?��p��m�i��1�D�EH��)ԴāTn��@Nr C�X&�lxS�D�,�X��Ō�
A�X�?��T)��SR!��2%
۰u|���3f@�b-y�d�=|��R�!C�'"Bl��&��'��Ujֶ/r!����N=8�)�'���o�(T BK]1L\�(��'87-��Jޘ*�c�p~���V�V�oWp�O&�s�����	џ�O�2�'| �2D�* o,c�$�5��(`e�'d��) ."iQr��
|�}3E#�6:��'���&gP�ID�2s
��k�G>q�F�����KOJ��0���@y3��4)6~t��2�&xa�������O6p�W�'i��O�(xU	Ӿy�L�����Ch2j"O��Ak rY�X��F��r��F�'\�#=Ap�W-G� �EM��v9y����F�'���'2$x�EkعX���'g"�yg�#���5+�11!n��҂�t�l��$ųJ��Ѳ �ÂI�Kv�	.�$� �,�A`�DgK��X�dG�� �.�3�����c�R!~����.�)7��h F�B�M5.�J�‵n�
�&��j�b�Oq��'��!भ̥
S�m��E_%�� �	��� ��YB�C
� Y��� 59������I��4�
�O�}��&^�|�"��PC�,P�!X�łs��	�O���Op������?��OLّ���	`h����n�T��D
{(�8��`D�;��{�f�ՎXJ⃅Z��I`�+�<��3��	�[���&	ў1��tZ�l�!9�B�Fy"��-&��݊`N*Ĭ�f�˥W]~UC�}�a��%�L{1�݌<^ĭyD���yreI0qን �Q�]F��KTN�Ș'�6�<��ڱI�@l������"��l���L�!M4�P�O��T�����q���|���|�"GA�{|E+S,,�	��
6)���\�����U� -2A�I�,�<�O��\q�M��lF�n�`mh�����-F�5��c�2Z�u���h���<�f�K����K<�E�͏ ڼi�̄<!% ��@��_�<"�X?wƶ8�W
tmHP�K^<�հi��jG�rD 0�:]X��2�|�%U,DZ7��O����|Jծ՗�?q�듹N�:�ctGO~F��9��@��?���N4,���b��/H�c�,��V��H�Q?�Ol�e���I���ъf��2���H������"G
ؑQ�&�05V�pw�Tb���Ѫ��
'*��źeҘ̧O��%�'r�=�	*�i�9<du�1��0 (����1O<���Ob��<�����_I����$T:x:!CØ�ax��cӊ�n�D�6z��P���d�p��B��
T�-i۴�?����?yC�A7w@xs��?i���?�;4�th�u�(N�T�5�֛4( L0�J�oPR	b��CnH�h��ό��O$�'� AA��
�`��;b�^(P�$tҡ��F�À���9c�HB|��ē9�V]��ʚ�'��q�!�F0L
&�;��|RF0�?�}&�"����C���5���67��B'�<D�ܻ�.ǽ�2C��\�V�:t�9?�q�i>e%��pSl�D����5�T��f'
/(�Vm��!^П\����ɉ�u��'�:�.�;V�Y�YI<4C��6��5�`&M��%�dO;^�n�q�ѿ5
�?Ad��M�\�@��M�k?�#R�E�C:
 ��ˑG>v� Eũ��Y����.G�@f̂Nc\l�'���𨻄�'���jY�M��-��a�uτ	��b��ybB�a�B݉'h�"�>�r�G����'=�7m/���b"H�oZܟ��	�h�,�c�DS�K.FX#FCL�g�.!�I���G�D����	�|Z�^�q�EA�W���h��K�J}�0虃wH��ɷH�ZP���ؚ>�B�<�1���Z����.ẍ誔(�^v���T�V��2E x Ɇ���u2rI������\BL8���u�� ħL�h���z�g�(9!�d[5:�8�{S+�?|�Ā f
�j3!���ʦ5�cC*�b�`ӣO����$#s�I#a�����4�?q���)�;4���ĕ#)^��$i�s�Rb����H���OV,A$�I q��P,�	:m�w�K�DϺ�W�|
Ѥ���N܋�mѩQ�,����\���e�n�Y��_�TB䱐$SA�|�3v����	ڲe� ��T�N�:�a����'[�Wq@5�I���S�'j�b@��ܥ(�^<`ە}����Z}��1en�@S:��nB; � ф�I��HO����RE)�a9ƮL�^���ۦE���<�����B矘�Iݟ��i�Ś�I�8d=��0��7p(�e!֫d�a�+*�6M��c)�iԫl�'QGR� 'mh�(�ӛS��h�Y�?���@%H1��u�iԦ����?vI�$	��8񩇲O�@�8�w���Gf������I����~Ӗї'�bL���|����'|2I���׍x��d!���U��4I�'�tXG�� �,P����W̆u1�O<�Gzne�����<q��+r�^�/�B� �TBZ��r8
�^,�?���?I��~��.�Oz��q>	�".S0~?�x�䉙$|w%��aɓ���g �]�Rͣ�!��[iz���_0HQ��7��=R�Y�
_�Oz֝�2A��
�~���a͜�:љ7��,f؍�#l�r�|X�}2d��&J8��C|q��3��)'�MK���a�)�%\@�JU�"rb�4L�(��|�� T$D$a�$ͺǢ�&���<A0�iL�'ު4�Azӌ���O�M1!@ZGP��1 j�,��ao�O����.�p���O�瓀p<M�aȊ��I�bm*v�=@%�*�Y��Eq#.1���T��%XC�(Y�J�aw��j��m�i�o�s�Bq`��M
2Y)ee��\�^U�S�'Y+�_(�'��X���"�h�Ҁ�2O`h��	�'�"��γG4M��m�<O�Ęj��$9��|�iV�IT��o�BL�' �>D%z�p�|2#�b?x��?I,����a�ON��/�|;���N�v�X�TA�Or��ܡe�6Ph�DC�rqT���m�IN"����AAu�ʧ	>�1�rf�	G�����?n��|�O��@D)ӿV�.��3AJ,VD����C�(��̟4��T�,�����O�G�v�j��>� �ПT	�4zz�F�'b�~ rB*�pK�@�alZ�h�*�)����ON��D�	�x��p��	^�8̘��]�H�ax2$ �S�? $����u�i۽{a�Pʆ�ʦ9�	����I�����������������ߍy���$�B�Q�V�x�s��O�Tɞ�	�
M�������žef��|���#Qu��	9<�D0�`_.�:lQ�"�>+7L���@�$m4(�ˍ�L!���A#(�S&';(���2O|hsU��=-;`�c��%[JTa��]����/O ժ@����O(�Ol�k�gF�n�Lu	E�	�
��R�"O^,)v��W��d8�n =Ov�Ta�'_6M�O��`�p	Zgπ/=n����$N���:'�������?���?�w������Ot��
��� ���;$����b�Д�A��I^�<S`ie�֦� ��1�1ʓ;����RdĮA�v�1%���Tܙx#�ܛ-ZB̫���	W�
�3Ð� !�2�Ȧ`Ƙ IN>�ZȐ�&Rt˘�$M5S��8V@
؟�H��FT�(��D�5��0��M���S��$�$I�
�#�hܺui�/fi�x���;�I��M�L>&�,2�f�'�O)7l hqUM�"��+ԤY�Y.��'y�|	�'B��'m�����0��LJ�O&08� �=�@�; ���vfƨI6�'�4Lb�7�
���10D�(�&ϛ6m��
a��Gcvh1�G�R8pD}��ت�?��iz��Q��H����JP�L2���?����������MĂ>��Y2�L�v�z�O qnڮ�t���K�m�������K�4����u���l��4��R��,	�=���=<�p`W����	)g/	�<���'�q@����b�^0��+'ᢼYTZ>ݗO��P;nM�0�*�I_�X�h�I�|��`��f�VI'�V ^�I����#P�	�c��BI

Tx1(��#}b��?��y��$C^�MX�# K�!KL���o�&�y'��j�c��@<e���b%���0<����]gEzr�U]�0īO�
� ���4�?Y��?9D�C�c~z$���?����?�;`����uO��T=�I�w��
 <��-��k�tH�'e��L����A���O��xQ#f��<�I�`��R"��]tJ��H���H�k��'����E����!�}���Ir���ɚ=&Z!䤈�%� ౕlF0��]��4��ɭe3����'U�'��$�fJ6
� h�g\�`!��	�Oע�8T���c@�l���R�9Of��d�'��4�'���S��u�`\�J#���g�B�fl���[���ȟ����Zw���'��%u����"�(I��\<�l��
T+{�l�
��k, �i@iMؒ	Ì��Q+zd�Y�0N�K�P !�Ƨ'�x���'��ˇ�a���S�(� �囋��Y�9T`f��ح�c`Y.(�����O���+K7�Сg��� ac�j����� ���נIpvF��qj�����J.1O�`l�C��7c#�@�ش�?a�R@����,�zH���B�|`(i ���?)�쌕�?�������@��а#0K(�sCɤ_荺�߮>W@���+!�l�C��!�"UGy��_�W�� �cX7�R��Q���v	�  ��9��1����jF&�7� Fyr�"�?ရxr.�/6|�JT�3c�H C���yb�W}$#���,;P|��f�OТ=ͧ����G%��@ii=0JD��,H �%�@�7oL��M���?�-�x�@H�OZ0�u�IO��	ɕ�+{3
<�%��OX��]k�Ƹ4��d���u�z�4���nαL]ʧ>�I�o4gfDia��2;� }�O@p��L&u��z���;
	�%�C�"͟�P�bǜ9:qY��i��j�>�����\*L>��( :TWKٷT����q��w9JB� ����U;9w��ڔ�K&2� E{�O�x"=)!�3[��)�E挓/�V���	����'�b�'����d���'?r��y'�1m`�pğ'J�zc��81r��҆�in$l��&ʁVb�9bd"擘a��2O��c���:dX䐚S�<
�f�rw��5n�Hyj��G1i�d���(tu*'hUc�tkϥk�I̻'لL`��@KT�Č�{Q�����|�D���?�}&��U�C�x�ʡ9���Rp"	+D��M�%�$�m9m��5Q��k����=�HO�<����+"2uCCJM�z�^���L�@��D.���d�O��$�O q�;�?��������5c�t1&��.-Dް�#.��1.�k��C�T�~��Qb@!����C%��|DyB$��*�N��>u�ȅ,Ώ��mp�ɖ9%�$9�@!�k��0�Ӊ�7��#=�7�ܑ9�]I㢉�)Ă(��L�5^���̟���H�'"����6*�zcwF��iK��!���D !���,OdYiu��!g5�-QG�F,1Od�n���p�'�l���v�����O|)K©^&�Xym
�\�*}�#��O�����Jհ���O瓏#J�$+�D�|&�y�G9|E"��&d�xr����'�t�)&#�k�@$KCo:۰�R���	���sl-��5t2Da��R2k�����`�!��ƞP)~M)c�±\� ����{���صj �諃%�(��ƌ���'v5jU�o� ���O��'8����S�? P}�pgV5u��� i�-D�d*�C�O����;9���d6�|�'2:bC�P�\b"0�d��D,8x�I�XAO0�S��1ˮ8hU��.����	��e�OR��'5.�O��cT+���(bE�2s�����"O
H�ԇ��@L�U�ޣ5����W�'#=a�'��S�Ru��r���#��zz�V�'���'X�uX��>!���'����ywO�0� ��@(, ݹ!��Y֢�*b���Ay�,˲�V�����e���"�)�j��'Xv�t/� ��`A����/����bʧP��d�3��
|�ڢ%K���O���pCA�<�M7�xM*��Rg �(��7,�Dz��DD�H/���Y�$�	����umX$�"$aEѸ�E�Iɟ��'�������4��%���rVi']J���y���	��M��i��'����O���/>
��b�e^�(� d(�睷��B�ɞj|!�O�,(�u��QZB�ɷQv�@��6�A����M.6B�I�$�iĨ])]��] ։�'Z/nC䉾wj�0��r�jM*�YNC��9-���AP�.KGf���nZ?L� C�I�BQ�L�����Xo��H�HDG(C��5q�Լ�ͼ3������A3WfC�ɔG*�Y��Y�����^��FC䉣X(l����n���\�3"�B䉛Hd��!�$�Mj�IԛR#Vp��O�x��Q�ܒ0�И���O&I����{�fݼ��4*�Ɩ�MDh���x�Tqs���E�݁&`��;,Մ�%�N,�G
L(��b�JHٺ̈́�1���ɑQ,��l	a��
h��@�ȓd�2H8@�5`�Q!��CO�h�ȓ2r��{�/�Kx���2��,"���}d�d�Ph@�:�`!2�˸%�Ь�ȓ|�ȵ�W�¾d�llp�d�W��a��h�!v	�qs�����0� ܆ȓgA���q"�Tz(�THAd��j���UܣkĬ����W�%�Jt�ȓp�q�+Fp�Qb� [*���ȓ4�6���&��k&��ɢ(�.QŅȓ��pR���_���a��$��]��f4�t����6#�Tق�i����[�D03�&��/s��+�ŞC��@�ȓ ѣ���]�2�k��$�Hq��@�(����I'��cF@1z0 ԇȓQH ��7	��&#�m�˖:�(���gV�qd�$ ��˥��#��݆�ɜ�0�;V�'�V�w��%no�ͪ�L¢b��i�Î�� e��{�S�4��I�`1 ��.{2�Ɂ46@�,13��8o� ��O�>F��O��Ѡ�AGR����ܔJc�X��>��n\!�p�*��&I]2 ����'�y�W�B.~h��-�*n}��fLR9�>ɛ2j$km;_�(�B��̳n tș6b +�<d(�@��ܓ. t#}�'	Z}y"��:L�����d7�d$j�홀Gk@1��640���͟�㟘A0ば%�v�IG��:�fݣ��9D3	YvbW�4����`�l`��l�S���ܩ4i����:S�)C��3G�ʜH�.�/qoX��7�(��?)A��-�Q�]qb�V�&{ID�2u��� #��$Ԏx����Wȃ$b��P�u�Iٍ}BI�.�vp�WGOO�<���bS)�ēb0��ۚw!��"Ɠ'�v���/�ބҦ�D0XϞ�ؑ*ҥXJ����S�JR�a�Ĕ�%�dT�B�T(+�8�� m&/�L�Z�CVUX��S��� 3`-�sJN�4|�7}��
H�h��#�=�8p`����'3n����
{������_����5�&$� �7��R����%�J}��/�;��I$��1Z�XDy�'MJ|��'r�	d(C)���IIގh�Dx�c,� 0��F<Q�T! k�q�N	��b�(��O���!��Z��E�V��)���9!�x�g�3�X
E�\�4���b�����p<�f!	3��M�ƃA26Z����w�HZ�L�=����3�ޙ�|�s�%��EJdAٷ��Sꜛ˓`q��C�Ts3(�Ҵ��B��D�OfQ�a'mt,�$1T㈑�e��EH�\���? �h��t�_�V�^%����*o�:��
��h�D�S��iS�*���{�E�R�.) ��X-6���N��4�+Q�"��?)"��6��� hL�W�U C�hYAU���v�^*�ִ9%Z2 ��5�~�j@1��>�'��fj\�~�B�SR��#V"e�Lb���!�����1����FY�vp�Y��g}R�G�b8�g�"8H�y�E~�*b���>�&�O�'���Ez����Z,ݡ��<L�⥃�ۍe�����=:ٌ��%N����?%?���iE'���rC	7�n5�T�+}�(�R���h��@�SY>�j�,I���'�M
Wo	�v�*:��Z��A��i�D�4Pl�=��|�Rύ�5����_<E:@IQ5�\�hu�	JT+ Ll��Q���O�@HS1�L��s�Ax�}iIL�P��=s� _������AL�)g�����At��� b��`��OHx<2u��CkNAz�!�˶�>�j�D�]���:����ez�$E�gr�����`��A�}ݶ��M�C�,I�%/T�W���2!!f]ĉ2���rBD�u�_=o�"㟒�Tt(��X5M�>!I��[��|��q�>A�їb�t�"�댪NŔ��A�G��w��=Ή�(�(�K6b)��z��ē�0|*�EђҊ��v#V� �,��F��r�,�%��*,�b�	���OI,��B�ܼ+e���汻f@�fWX�J��ۦ���)�'�u'�`hg�ʁN�h �-<�f���}b_�>�����5k�:0���Dŗ[I�0�N�.j�u�'���y�,�����=�{?��II;�\s�Nշ�Z�
C*��J�dpŧ$�bW��p$��C� ����dHBJ�'�	�zhn!J6�8�5���L����Li�a�9*MCT�I�!Ex��Y,@��o�e%�Ѻ�lA�J���<���ԟh�"�G�fypTjD<X�(��ƅ�j�~�h�'%F�<�SU(���=����s!��Y9���%�B�0�܄Q �'�ў"}��Q# ��ң�I�胄�@$1@�b��!A�~�F��$J[�Z�$�Q�"�y�ڰ{��XqF��@�� ��IN�'l���F�Q�<�{q<��X	�A�+R��M�5/��r�L� �T��*�n[$\���^LQ���'�L�3O�%z�v�� ��0��I�젣I"?�a��ˌ�b��ȳ@� ��4�8�gޗ`fJ�O ɨH���:�Sba��	C�%)���]��*���4V6�8�4LI���!؉��O���(���ԼK�`Fo��p�M�fd�xB	 ��F{��IѬB��d@0ş!Z>�p�+��Q�L)�}"j�Fӊ�H�	�4?i���͏��,��x���t��I�Dم7��U�'�Q���g�=x�R-Sr靌!�Q��e�"B��Y
Y����ܔ/�&�$*�=����1��q��LGx�gycO=>|N)"�$T6��-�@����I�z�ڔY$��iO`�Ï�	���dز�[� A��"� ��ӡT��?	��!K���t�x�J�ݢ.i�S��)�����ݜE״  EEܮU�ּ��` ����[pEb��AM̎��ݧ>��R�/� H���@�Û�hy�|��Þ~�O��'A8q���cQ�7�Ok�2�c�u��Dr��:{�@��}2��>yP��C�H�QH��x��j��'9�V!���Y�,궭�!ˀ�:!�kޜȦf�
p��zd�"yV ����((8�%zt���q�ޔ�7h��1}<���kM��ʘ��]�>8��yf����P� ��T��Aٔ�߱'����d��OB�Ba��)��g�'����N�6T��D>h,qq$IN�t�����)k�QPB��M�6�ɱ��%�B䉍G����v�P~�0y�+�[fn�z��_-qOa�D��2� 1Hׂ�?2�dlAn���0=i������' �A��J<L�y	��BiJ�
�'ˮ�q�l�w�S�O���J�/
q0�2���œ�y2��W����=�|����±�$.܆*.��SI~"AL�M�T]��	?�-0�(�,{
��O�6����$I�Ia��� ,�FiY�,9=]:����.�0>��I��4�tJ�A6,����%�c,�FC_!<H�M��C
�ݲ��'^GX�'��������O�d���mT'�A#��(�l�
�b茭����A�ˈj��� N������f��Q��pՌX0�a��TT.�	>]�ؠ	SŘ%s��xJA��B/f�G����kݚ�K�ߍc'H}T�I�y�^0�ҥٝ4���:r�ė��7�S��yBcųm~:���*k`d�'�#y�V=����Y@�k�,u��r W>Ń�.�&Gh$�IS��xe#F���k`b�DR�t��@KU�G"��ɻZw��O�O�,�wf�D����K��ܐ�A�Ђ<�f��E�ZK�Q���[�V=ܑ�w�>H�R@��Rrȡ�fל	�\���4m���h$�>�~�%�B��&p��?�	W�1.v���DP<V�\`��!/��W��t�w.L�;D���\3qX�T>�"W�l�m���wJ@|��Am���!��m�bu �F�O�>��A��(�kLL���W�F�]�"� �17�����A�4-h5��� 
2�2�)�'w󮉤.n�B�O�|��M�5�I���T����)Y!Z�X?#��Đ��=aee� U_>�zb��R����3�&(q�ÊW�V(q���J��:�Ȓ
J�H�����X%+i`	C𨃫l)���`\����<�Sk�p(t0��bӇ(�~9seMGuI�`�e�K0Z�6|���'}��4��ą]��$c���� {e�53B�ġ��<^�[C���wֱ
���]W�	��B*t*����SH���?L�M�e�'P�83!���{`���ǌĔ8�b��t�O�6@�Z'^�yp��;e���qkS0@̸T`d��A�<�AT��ɟ�|�u3Hs�4~H�E	P#y�a��-�T7P�� 4��c -��%Z��Ov�!��Ϊ�J�:Ei�	�����f����xT���v���!�9L�뎜���)�iӀ4�D[e�� Җ��D�6KU�Q��FP;f "ʓ#� В��V6IQE�=n����F�#G�b֠�l����Q+>��'D���'N6�$�Y4(��>Y�N {�<o
��dI�e�Xc�X��K	zd$8�<p�R��1,N�c�"i���L%#� ��xb%�*� Q
L:��F��o1y�E
A$�,=c�p����	|��c�@�P����7�O�MF��O�bf)о1at���� Z���D�V��J�� Ҥ͵���� {(�9d�Ƥ)@R)�MA�P�m�q�ؚ0X
^��!�j#-s��1���1���
j��&��g;N8 v��,3Jx�<1���=J���"���i�bN�E��q�ێ:��4�#6,O
����[�y���*�^�?�b���#&�P���xA|��ŠJa�_pd0�V��)r�?	�iH�m��) F�H�-��J0�D�
v�`f�pS)ʠ�h���ɕJ�����֩4�x�k�]�)t��D�N�/��I�H��I�>jlYw�	5s���1@�&EQ*e�%�٤�И��a¶(�T��xr�A3��y䇕�%��\�蔃�M&`������Kay@X9MZ��C�"� ZP�įOVL�Т)H�Z��)$$P�' [T�ԏ�L�Ҧ!XeŴ��U-V�y�8Kƪ����I�8���b� �~���QR�'����F�O9�lx�����"!�a�a��I�t �wX��K'�'��5<e��yd(��S��'㆏8��O��C�=�N�����"�h�* �G�)�P���ǭ3��w��Ĝ�V�}]|7m�4p�"}�'�$�����2��ƛ!M�<�JDBھQ����F�OhX�mOR�g�I]u29�f�U{�T�#��Q6v��Q/��)XĳCAERd�0ig�#>��f笍R2�ݡfD����f���phr��E�Xi@��(O~���n�&RS�Q*��Ӻm[d��U�IK7���@�X�l|f�ٲM��U�#>id�V�Yܨh��׬s��b�A`I5@��.���q"�:��'�Iò���%áe� ںݑ��~�D�2(_V�[�����Ar���n̓H�@p��۞(Tj!����ͫD^1Ц�I3��x�i�	(ڽ�E�3A�Ӱ+۪&����d?)���N����X"�-���rQ�yT�1���*o�>�i��u�k؟T���r0n\=&�Q�Ra[}0��K��Ck��a6��ۊ���*aPbmi�.�:�x��kO,��-ƶvi�0�ׂ'��?��c_ZW��R��H/8ƾl*��B9F�v����mَ��g�ۆ��O�uHƊ��d9�;Ƥ����]>s�������r&��>�Ơ��I����o�6y�6�ߌ�ħ(�v����E
��=��. fUEx�Ԍj���F���S�Z֤ ��J�S`B�YkH�iX>t�aE� ��E8�'0����Y��a,Wi����Ɯdۈ�L� [Fr������'Z�и��U�Υ ��D���4ZW^����əT$�tYg�8<O�-x'�2P�́��AYN�@ٵ�'z<)Iǁ�`;V%Y�FN�A�Yʗ"S�Z��1�ˑ)<6T��2�vl*P��<fzA�b��`�>q���D��qٵ�P5Zs�?I8�P"���
gk��T2B<D�DBFc6)��z�)M,z8�S�J$�F`�&�wAX˓�h��D�/��i��
�t�`:�/(�!�D��O�	R���9u4H0��~�!��D7}�
q�쀾[���hl!�9m����`	 T̢��(F��!����`�b]�)1��E/�!��J�\����A`���
��H!�C/Br�1B�نE����	�\3!򄝏yS�܉e��J:��F�T-!�����5nM�>9
pS�d�k0!�ެJb�b&`^�KP@12�B�lv!��ԣ#z�]c IT;>TD���@!�ɘ_���pu�S�Z�6q��V�!�0.6��`�Ȑ!{0‡�)~&!���3����#C�8SlVl"�%�r�!�G�Z�<���\l�&C�5�!��܍^1�,�Q�V�EX@�5��g�!�H�b�b` bNe�&�� s!�(/N�t�  ��^*D\8��\]!�D��d/��ZU���4�$z�j�2@!�� �x�¡�J�����L��JRb"O6�c�=��ŐI<�*$� "O�ā���Q�IjE�ɱ.�n)�c"O�P)��rXF}s���qz��
�"Obؒ�
O'2�IS@�3yLX�"O�<*�b^���ӣ$J[v�"O��@hW�N�|%P��4^"v���"O 9�煙kIn|�����8�q�"Ox�s`��Yo*�9�eL
q��2"O���Eƣ".؄�#OQ!���"O���%��^`$e�aL߁}��a4"OV� ��,A�J���DHd~`$"O�I[�
�$H�ؔP��E�j��$"O�A�W��0P&�<3䇔[	6�۵"Oz���d��/�8�{Ң�'j�r�"O���+�x��J߽&9;�"O8�q��Ը��įZ�#��;�"O6y6h��y�R��5N\��)T"O��)b�%`]�x����+R�a�$"O��I��_��I��-�P�X8 "O�D
p�3���R�	
F�=B "O�(#q�HAS� a��#"��dx2"O�\��䌀E:6i��K3w�ftRu"O~����mP�$��'4S�ܽ��"O���E>0���� uОAr�"OX���$5Y�t`��X�L���Y"O�Թ׃�`-lȹ�,\�����"O�(SE��C3��K�d�t�X&"O��`���	P���򨎈	�����"OT��&��~teZ�hO�EA�6"OJ�)'m�
 �p�J6'�>AH1��"O�����#��x�s��E>���S"O�9���}��jc	T��.�˂"O$QC��.���0q������"Ory�%]>� �iT
]Lh\�U"OpP��� �)-��Mur���"O��F�^�T@�b��#����"O�� u�X�VdZ3㐯m�
�"O�	�A�=���P�`����"O虪V��i�na�t��*W̾$�d"O��)����Cn(a`+̓T��U�"O6����댱`&Tzf���d��؆���t[� Z�\�񲈙�|-�$�ȓ]d�9�]��Di9�Kƀ@�X���g R�6hL�e��1�A�;�"T�ȓ>�p5+�� k ���Y�2%����h�Xȡ����Y�f� ��ȓ�(0�F%"y9e�E(�ȅ�A�i�! X�iA3�Z76��ȓ
�ڝ!��W�|K���D��?0��ȓ$����R琦Z�:�6��/eFꀅ�v���f��s�T��AK�#D��u��Uz
p7 X]�A�3���o���ȓQ�@2p⊍m0�lQb�іjpf\��if��@J�v�j���d�
 ���y�BM�Rr��ѥ�Œ�@�1��(��=1�y�	Y�����Yw�@�R��7�S�O8��Q׌���M�Ȑ�t�l�{��)���)�lh �<��b7��=X1O 7-<LO�A�C�A�"��T3�
&U���h��Ʌw��O���O���r�ͬxP	��@6|d����'g���T��	 ]Ce���`|���O�6=�I^�O���
 #4��rT��T�,Q��'A ��0g�m1��J�D�Na���� �y��)L	#��T�THqN�:�"O���ؔq(�R�'�4��#"O��S�@ħW��#'Cb��h�"O�(��+,-�Z���� 3N(��1"O����i��߸	y���;>q�A�'����5p�Q�K0qjx׭�*z#<1���?a�u�ʒ<�� �6퇫�^�ɖ�)D�����W�M=�eƆ"1'RLj�3��舟2���/�%�9��B��Cdd"O�u�#ʊE��Ȳ�7dD�-2e�'��	�x{�����X�����g�(o���0��9��V�$"H��&��*�.0�B/eӢ��)? ,�j(x �B�m|Bq ��nX�HEy�.^����QǮ^%��0����y2�)��ܰ�ҋk)ʄ#a) *I5����|Zp�a��k(���A�]I�O����ױd��]0r�Y� !�Ef��:�!��̒)��|�-ձ1H�R�[���Iox��'R�!��T��B��wHL�YQ�hP�'7��!c�-<�jR��Rl������#�S�t��h�]z��
	Q�ʓk��y8.�L��g
�D���FZ�yR˓#R:�{��M@��(6�J����	e�S��?ya��?X*4r4b��9�JE�.FN�'�̡F��B�0#H��!h��b�2᧜ ���%�O���CnF$�x��D����i�pH<9E�<;BZ\2$������V�K�<A�Ij��.�@��Ѻ���ȓi��8!Dk�A�~Ń��>@�x���Ntb�I7�pn`�D@=����>qד
���쀍>Ċ!c�Z6:8�TGx��'(�h�[�@t� ���M��lb	�'�j(��7s�J���n�<0�"On4
�NO8�B)!P��?g4�����'=@���闈PST��V#������L�/p!�DϠ@Pu��̏ \�1�O�FW!�$�;����m, ��sLJ.j;!�	VR,b���v�e��@��"!��OڅP�L�N�-�I��>$���$�����Ip����b��\�n@��bEX-�6�;��9� �m�`q�� Q�p���"D�8��IBӡ�!E�8����$D��X���@��I1A(J��6�:��!D�l9��/_�08���FO�ٚRH?D�t�3����\v��O��@Zt�'D����M��bl�Qc����ۂ�$D�YȚ2Q:LX[�$�4*� �C�#5D��R�vl8<y�*��ث�4D������5��$颩�Z��8K5d1D���␑��I#,�A����Q�2D�(�l�xoT4����u�<�/D�t��mĳB{���wF@0A^��Pj-D� 9�Å\,T1����(�i�)D�8Hd/K?H?�!&H�2o�h�O(D�h `N�=8����u/�E�'D�����4$��M��ď1v~�AT�&D�B�Fc���A����_����$D���Ԧ[5l�,ܢ'�����R� D��� *>�y� i
-/���A D��@e��q��" I�=�D�r�̄�I����㭐!M��i�V!�L�!l/D���������g� ���+D�8s�I�l5� �B�S(/Y�?"!�D7{���A�2%��S��qO��=%?� �=	�\`�`	���"O��S��E�ǦQ�Ҫ
��YC""O0�	�EI&qx�\	�,K�d�*��[����I�	��]���/O09���,8�B�	nW�(g�$=M!��& bB�	�[��Z��U�V��@��4�<B�I�bP�����MB̓͏%E|�C�I:P%KsE\�&�8`�����C䉚وiГS"2�8��k��dC�I�^�Z��c�f��	с�D�|C�I�DSd) ���c��\ҢHY�s,�C䉋"���+T���M�R�ukyfC�	vV({��D6)_f@"�/A6,LC�	?>y̱���3N�Hu�R�<<�C�Ɏ� ��T=�,�+E�{��C�	"3'�#�E;4J�FC7$�xB�ɜG�ؙ�bgͤrN��"��!�4B�I�r�)"@�:X��p�OX;4B�I�R�DA��'�T2�-x��ԁ?r�B�I;$���˖M�Q"��X_<C�I�)�l!rW蒴q�>hbBR{I
C�K�lT8�L5�4 )�K4j�B�� w�z���
5(��Z�˟2S�B�	�t\Qi�@��:���� g�
ڄB�� �4+%�--t�����`~C��5=>t�͖:d�r|颯P�)�C�ɿ :�-;��NI�X�'�E��B�ɳ�䛲�@�oG�kы̢*�hC��&^�|yp�F0L�� ��Y��B�	��U	���1"��!㢤�5	��C�I�p�+�׭kW��B�*FW��C�	�<���C�*��_�mX�/��R�|C�	<rj���V�+Ū%S�o^:	4�C�	*%���f@�_��t�� [
;ńC�I�d]��#�N
]��J�"�S0B䉘^��x�@�01`����*�j�$B�I�i�X�˄� �>��T����R
B�Im]~�sq Y�Ps�J�xZ�C䉰��XR)]���Qha�V'{,"B�;4,x`Ӑ�[�%���At���K��C�I3�����o�@eY$aE�r�C�IL��(3ХɄ- lQ�A7�C�I1-C��I�GM!2(�=��*Èd�B�	>/�����ò~���7k��$V�B�ɫ�СHU�R)umZ ���^X�C�I)cl�XA�.�0C*H�fH�I@B�/5Х��$�1X����4�2B䉶p��r����C��1�VH�-2�B�I P=p�Aģ�7o�ັ$^�2��C��6Z��Px"�[�	F����\�yQ�C�I*x��US�i��&:�#pc["X��C�Iz�Xc7偹H;��$�DGpC�ɗSD�	���CL0<��-J7�XC�	���u�
M�*ԛp 	&a-�C�	�	0�u��C�;;����n�2;X�C�I97�F�:��ŉ+�4�
	:oE�C�I�c����6���pɧ�ӽT�B��)W"8��tgݶu�%Z��HtB䉗;)`(r�!��.(�Eg@�(?`B�	8@YjxFN�#4����ď�(VqNC�I�-�p,B.^1rA{�)>�C䉌G��X���g�8�҂Ďv%PC�	,�Z�۴GL�zi�wb�(L�C�I�2�>@_l<�;���>;��C�)� ��B&�J�)n0����R�E
7"OlA��? ;�Lp�_ ���C"O4�Ч)G�%�P���ޏiNt��"O�qɢ��XrНC2h�"��1"O����E� ۸��'K9�n���"O a`�M�~��˴�͗<���*�"O�I���|�\�a�܎��U��"O�Q�!Ď{*\���#v�"��D"O���7���i�&�Q� ɪG�8�k�"O ��T�5ޅ�@��P��pr#"O�d{B@KT��Yz#o�c}r��"O���G�]��b()ѣ�q��ّG"O`�2Ue�:��lȑ�+m�b�"OȤ�sō�
���
'GEtu�"O�	��	0U��|�wJZ�q���I�"O^d���S:"�����P��&��p"OfA� @�o�0�P��n�:��a"Od(!2%�d�t���匉rn�C�"O�u���ӽu�J���΋6Ha�
"O`)@�˃e��XمmG.~F�h0"OJ�8�c�d���̑J#J�`�"O�U��e�9N��[B+O�#�p�Zq"O�DU�_�O�D����7�|u��"O�qI�JO��\�sÎ�=|�����"O�麱l�$Й�->�^�à"O(���>m#�d
T.
�S���W"OdT�a�U�q������_ղ�Qs"O���@&Δm�"
_��|�A"O�@�cĬ�0q���L�}�4���"O�����
~P�ƇQ9	�jE��"O =���Y�l����~�d�&"OX�@ׁP�t�.�PU�5�Q�E"O��̜ ��i��k�N����"OD�vMV�:=:d��B�D�Q"OP�QE�h��L�(�>����0"O��&	΋>"6 )�P-1���E"OyS$�ơj�Xt��IǮs���p"OXi��$�0����QHL/M8zP�U"O��S���5M�,Ɂ��3)�x�4"O��7fn�P�7IX�)���"O�{c�ݐ�T��b�:�b�"O��
Ə�(�ʱ�Dg�+rL��!"O ��L�O	����%	�&\��"O �R��W"��*��/1�z�#�"O��D2&�����F(?��Zw"O���a�%hIɱjK)o ��("O0}2Cn��������Yn��E"O�!���K&Uj�ȓ�f+S�R�1�"O��XÂ�f�&��!�O;~�m��"O���"oX;+V�#f��F^\@�F"Od{r��6C���[�}ZzT��"O�];'S�c��t&2ĬB"O<ݨcj
�D�i��!29"O����a���1	tGI�t Д"ON	�D�:~�3X�&)��J�"O
�Z6���?�d�ĉ-U%0-)�"O�e R�C��:h�I�:0��R"O�dh��#uC����W�~@�r"O��YN�4Ȅ��G\�p x�"O0Ip6 �3���B���$W&�+�"O�R���(<��.A�y=Vu��"OD���'������A̋1����"O*�Pd�7�мc��#NQ ���"O�2�'ܒ-�l4sq�;&E��c1"O� �(����Xu&$�SJ�!c*�
F"O�)���(A�CƂ�4e�j��f"O��h���c0j���aI
���T"O~l�V�ެ`�"��nK7x��A�"OX��6��<�Q�$-��{�
E�s"O�Y�Q,����F���HЪ�ZD"O�uB���[��3 �ּW��=Y�"O��a�ʜ(�PŃ��-/ܤX*a"OlA*��]�45���䆷c�����"O0�ACH+=)���#Y0n��蹗"Ob9{�nŸK?mx䞥^�BMh�"O��!�$L�~I������Z ��"O@���#YE*1��N,R)�	��"OVM��O���J�'iN�x"O-���N�n:V�ۇb�In�U@S"O����MI
/R����G�R��&"O���k�*C���S�
=�H9"O�l����6E�6i�7j�3V(=�C"O��"c��d�͹�)�'�0�c�"O�@�a͍B-jXf(^$����"O �P�NE�c�R���G��D�}җ"O������>u&*�A�擁/�F8��"O|�QDA��Y���r���$j��}+�"O�<Ht��J(�Pj�		�X��"OL�[T
��yi���\ �,j�"O��#����@��T��hɬIWlM�"O����_�pQ.͛@蟊��A	v"Oހ�%/�5x? ���v�����"O�!��Pk��J.����"O��F�
�Ni W�/S�p]��"O��Rs�ΗX*�������"�"O�� &螁h��ts@ܬn�D�x"O>ݨ�+��s�ق�)�bqYS"O�i0J��{�Iؐi�yHn�q�"Op���[�u����58��p�"O����E�	U�*��U��So��c3"O���g��؍Bȓ�=aƤ9�"O�(�m��}ޤX�$v�8��"OZ(�3$�X�C�!3,x3w"O�ujRK<H��ƁY"i&"O��h�a	"`W^LAW��1��@"O���\�#[*Ma#.
�M�6��"O��*��\�N@F�ip�əf��"p"O�e���X=c��U��N�~����"O�!�G�΅/��$N6s@4�a"O"	���ì�t*���`Y�8á"O����D����0�ѐJ��3"O\��"G�\���Vg;��k�"O�h��O�qP���ȆV0���!"OୀW!M�<�&�p5��-�es�"O�c��N�k�lQiwGU"d�YYT"O��;1KI�\^P�����q�"OT$&�;ETb):/Ļ���w"OL�Qg��khj(P��:���G"O��J�� r���ե\�����"O~q�V�F@!�� �V-��"O ���R��� c��V�j@"O�L*�JƮ{ ��J���c���`"O������I؃&\�N��I�"O���P���K�x܂�EE����w"O�qJU�
%K*P�[�zS���"O����$L.س��	M����"Oĉ��a*[���b�
*/�%��"O��W��K6�z�J��`�%�1"O� ��S���P�H�#�T�Q� "O�̲��^'/�,�2���W��ճ2"O.��bj����)�vgU3��U��"O0p�PA-��Jd�O�x�l�(0"O���`&����)&�D+[�^!CU"O�mH��@HOR��F$��:�ܵa�"Oސi��8:��i%Â:2���Q�"O.�B�e�*7��(���*Vp�S�"O�!�#�
�|���� �5{P蔠6"O�*S�V���� m�T��RZ!���,�$���ς�
�F���-ȃg!���0_������a��i�Bm�,P!�$��w41�`�@#�������
@!��Q ,>�A�Pb�1�f�h�(��s7!���0�8�Cad�6B�Ȅ���s!��ψz����FL���!2�O,!������1��%P�� ���W!-!򤞤7L>��P�E���u��H�m!�$ȇ�\!P�A�
y�ٸ(P F!�D�U�,�9���V�g���8B!�H:{������VGR���O�E!�@�V�� �S��~�+3�/:6!�d�!@��ra�H7z^�d�V��b/!��Z$`�,��S �)�Tj��L:((!���5y͂H��l�g0�]ѡ]9p!�$U�K�
���&D�MG~�ST@� �!�d�3t��%�� َu7�-3!@��7�!���1��h�B%.��1̆�Y:!�;:e��'��k@�`��!_ !��eoJEa4��Y��ēs��:�!�$��;�p���1Z霡#C@Ƞp�!�d��d��p�D@JC:�\i$a޷O�!�D�x���E&��t4������?�!�� �ؽ�#��-\1X	9T�ގ`�!��+FI�㝃^�y�C�7c!�d�%��H�b# :;���yP!���uHB��F�LB8A���x>!��҂R|䡕CT$��m*3�/!�Ď$?�@�b��X���Q4.E�!�8W���4L�%��h�d��M�!��
(/ШđaE�h���u���+!�d�G�<�S`l�JkH��H�\!�DB��x���gLx�y��CO!�$�X:(h��R!E��"�O	,�!�Y�l\\���[NpH�Ęl0!��ͅT�|)�&�,B����m�-!��L��B0*LL_ ���p!�D�	&L(�r�<%�A!��-&
!�$�E�j���Mb��Yn�!�䚑v88��q���z|�Ж#I!�$�7C�1��#�
m�D\�� ڷ#K!�D[! n�iK$aS�=|^ %ON<e!�d��������9q\�B����!�d��/(١ACAQp�G�h!�D޹4�����c��<K��k�+��z��&���A �19��ZRc�#|%�݅�Alj�{���c@��B&X4`�ȓN�����-��+�����ዯ2P�%��� ��&]�b6nJ�B��u-��k��g8M���
�XZ.B�Ɇl4�����M+"��tR�OL� 9�C�	p�"��u/̯+(�x�L��kJ�C��J�JUp�&��c�|����4�@C�I,�X�I�D�XT��ŤEG��C�)� 0���)gdRp	ƪR�s"(�s"Oڈs��Q�a6m��I. �Te�f"OP���b�N�փ�%w�&Ѡ"O��)���\IZ%!P!v�n :3"O��sEbC3.�n�����ɨ�k"O��P�"XL�i��ѹ`�F4�5"OhX�I7�>1��R�~��"O��%�ʪ��@�t	U����"O�h@!F����u怹E�m�"O�p���$,VfHq#�K���Ճ"O��!�  �?nQ�q��h¬eI�"O�T:ID�@C�%ۦ�C�?C,� '"O<hS�l��l��8�"O �;��H�"O���^�~7��MƓ5Ą:�"Ov���fH�f>D���K��5��pxd"O:�*�ЩUʴ�	��=-��T"�"ObؓS�����rǗ:m�x��"O��@kͲeM:�
EF�'�q"O�8X$G�����&-�M�c"ODc��_)�uh��с1�0mC�"O��i
 4m��2���:&,�S"O\�qA�TvN�`i��ZA�� �b"O��B��ЀT(��M�c�ZUj�"O�,���ŝ|Ң<�
R�9Kc"O�Hq��)(afI�r*�9}�0uI3"O�<Y4+ɫ"#>-0���	����"Ol�c�.�����@���Y���h�"O^�X��	~D��2$؜+>~�B6"O<]� ř4;,�:��ے=��P��"O���R��G�R1��3�T��W"O� 򥊠]/ڔP���$!@���"O,8�` ^�l�8L��Z3�m�F*O�XG�F�b*e���:{'�-0	�'O$�� �Q-��XA$U�zP�Ԇ�|f��)���W�B� ���:\����ȓ!���{�"B�V�~=�u&�7U.D��~@hȈS뀯T-�M2b�]7a<蘄ȓAL�iӠH�N����4Kdy�ȓl��Rk�htd��O;T:�$���4�R2��4F�<�4@R7q�<��lz�% īO�qr��tg1]��y�ȓ_�4�!Y&�0`s����v�Մȓ�T@a��%{�� �E�����:��}����H6��V��]�h��"���sed��q-����oÁg;���2R� �(1l��Q���*�LU��`�JȈ���"7�H[s��7�R����H�J#&��#:��� V�ȓ`Od�;�O�6gځ2'��;N���"T,���@�U,�Z�!�,�$�ȓ H��P4`WC6�pr/ɒT0�p�ȓt�� ��+\�R�*���	�{��a��0���:�T��䚧Z	�|��_�&X� �"_s̥Zڤ4[�lI�'���*q(�<=_>P�NJ�4u���';�8Z �jd9�V��~{�R
�'+ތ�S	��?��1!"n)�a�'v�(������B��T=j�-��'K�� Е0���a���	�'jr0KeN�AG$���
�.e�R=��'X�Z�eL�)�s��W�0���''�%�a�R1Fo�$�AX����'�@��N�T~�'&]�?%���'s��11	�C�|)��Sc�aK��� �,�lQ�~�J�F]�NF��v"O������!:�.̼N~�iA"Od$��IN�ѣ0��XN�$�E"O��"�.3�j��k=b_Hpӧ"O�9��У�x �c��bU��p"O>- ���(RJ
u��ٮTeP�[B"O���nҦ^0�O�u{��Ȕ"O�d���9v��h�P�)-,i@�"O�#�%V�./$eRӪM�3
Ġ�q"O�E8�( |�p��R� s�ڑ� "O��ʳ�ˢd��t��	/ת|C1"O�A��ė�NV��[�L,5�X6�2D��2�H�#�0E%sKT��)0D���M�<莽� �5"y@����#D�����ާ8PV�A�舁R�f|�c?D�T0��Tυ��0R��q����2B�I�Y�����'0ڭ��Y�XC�I^�@�POK�:M�SDK�<;hC�	�n�̡C �D�X�����#ƚ3��B�I`�0�����  Z��%"�:M��B�	.q��$� I�'�e��B6"V�C�	�>��8�C�)v���3K��2�nB�>��M�cg���}����t�XB�ɦn�m�B��9ho�Uh��vu�C�I%v��(6��#mb-�J����C�ɘ'b��
�e�5G�4��)@f8D�(���W?fhS�͓hVŹ��6D��!���#e+�{q ^6�M���0D� ��B�,��T;�m%q9��#ע9D��Z�ˠL�m�2��
i;�̑�m;D���$@�Ӵ��5,?x@�}@Wm9D������!�P��a�*	�P�*2D�<�U!�=iTY��C�jkXa�v,D���2�	�s5� ��%��/�6(��+D�x��h֔Ur!�A�==z�p��%D�@�!�P5w�=��h� Rn�����#D�P�`��7;���0�����6D�hU(
,7+�,��oV�|	Πq�8D����Æ�P6R�!S�^��[�$<D� ���
������-lh�2C=D��q �A�F���k�]�n���l>D��A��;)�>TY-��,�N�a�.D�@�a�n�Q%��	T0p�K8D��0�AH�((��P�d$��18D��d���m�@12׌<_k�)�4D���ģBBÎ� �4c�M	�N2D��"��PF|�� �(QB��	�$0D�4��M�V�D�	�%ͭT�P`�-D�<�G�[;V��:�H�6_2��t )D�ЃR��m-��Y׆�6ƠX��:D������l�����j��y�*O6�#�(�q)0���n:�YK�"O�a0�O~��9G�_1j{�l�P"O"x��a�:c�v�6	տR�"�C"O���r�9,���K`��7x���@"OFa3t��d<&�4�^)h�]� "O.8�`N� 3��dܱANb�1"O�q�2�I�T�&(Q�L�+4:���"O~�k�g̈́c�q���*+#�q�"O�L[ ��O0�8��jܑf��@C�"O̙�ck��6�����C��E����"Ot����99m�����ɨ[R��"O���
�zA�t#ŴOd=kb"O&�B�$�a�w�.����"O� P���J�4v��� 
])'��mbS"ON���Ѓ=�8��
�,K���3"O�� W��NZ��T�0�����"OBm16��8�<D06&[�W�tL��"O�!D�K���e�_~vI�"O��z/�c�����D�U��"O �#�	e���Cn�� �9w!��Y�Ai@}rň��@����2/�!�d�3<tX3�n�l��T��!�D��i�lY$@N�)uu`��W��!�N�2�Z���8[�1�KU�!�Ė+l�6K�i�h0�P7z�!�	t`h8G��0�X��H1�!򄘍i��j�b��*��{���#�!�!�qqǫ�tj���[�Y�!�Qi���y��3EX�*["I!�dT:8��H�W�`as�U�*� �5"Oj�A0A��f��`�F�ތ~�:4"Ob�a�q�8���ݾGh��"O�@&G\��J!C��4R���"OL��c�"�f����E�2^��F"O֜1 jO&A��[��#x֔��"O��Y��M;V�K�s �:f"Of؛�OM;h��rʐ�G��!xQ"Of���Y�?U���T }y���"OnLc%h��	���*Å��1y��9"O�pk���F��E�G��n6H"O�X!)TFMS3jؤ��"OV��W@GFJ�ك�&Ra�)B�"O����O�4ĸ蘣GF*�3W"O�=�b�O#�P�z�f�>:]js"O�1ː�D�Rށc�G�)%��`V"O0L� ×��`f�_i�w"O$��D�)s�4���g��	J*u:�"O�hy`l	�oF`��B,�1�*(��"O@A���/���*ڸ2���B"O�8�i�D(���
F�#���"O,PS�(���h��IR @2v"OqC�"�"'����& �Fh�"O�$�� �R!�q�sE�Z�]2F"Ot�ñ 60�������f'� �""O��H�dB�fz �悽#(�,��"O�u����f�b�d�M'
�!"OX|2��OyPL���F�_W�i�"O4M32�N�αR% B�D�ucf"O���SD�@�ꔩ�lK?�~L��"OH���l�d�8���錔u��ȉW"O����P>&gR�h��G谄"�"O
� ���`9v|'�)1�\h�"OhxI����H�)���0�´"O>e:��U�<��y�֔7����a"O ��"��Z�J�yiB�l!�E"O̐��m�W'��3#(V~pPy��"O
�R�+�Y��,�4���XF8%�&"O�1����вve�$S�6q��"O�����F LE�5KϏU���d"O]�5D]KP� ː�q�J#C"Oи��tQ�g���<\�v"O���ې(Z�@�S�C$~�2�+�"O���g՝.-"���%�/Or�僷"O��Va;N�D<��e p���@"Oʵ:�Y=�D߉�H|�G"Oν��������vD$e���1S"Ob��"�׷Q�1Z����-�FE
F"O� �@jS�D�)Ŏ-��ש<��)�"O��Z�[,kD�p#�i e��H�"O���`�
�@��5��(��l�S"O��jD��+�b`��˘n�ZU²"O���D*(!~P�S��7��Z�"O ƧY�h�T页�èm�|�+�"O4(B��S�iT���@C�!����"O���e�>.* �qFS�p\-;"O0-�ֈ�4F��EvD[�
Fj`�p"O�u2�EL#�y�`����ӵ"O8q���i͸e �:#�KF"O�5J��� t�@�	ȵ\���kB"O�1YGg@�T��`1��;,h�""O4YT���2�U� I��Eyv"On���;���ђ���[��"O8i��Ǐ~�´��Ǔ(Jz|�r"O�!��f�u������2E^΍ "O���ą�7�apvg�$&I��Q""O�m�����S���f��p#��p"OT��v�W1Q�؀�k�7yb�2"O�1	�+�4��y#KX"`��"O�i��C��>������N�Q"O�MyeH�T���hє���"OR1��Oڸ4 j��P�$�����"Oȅ�t�F2p11G(Gi\ux�"Op�	ۼ0WN����3^)��x�"O,��seI8��H@��ތ�"O��
Q�+��Z�Q�H��m2�"O�@F���;߾ق�H1H<u��"O�8��E�a銘;��g�8��"OXQ����=N5��K�*G9>,4�"O DfBƕ�x�q'j��ww����"O������� x����R��
=1�"O���a�!I���ۇ
63�Ʊ�"O��IM�;}E )���ӻ�8���"O&�p���p� 3�U#
r `��"O��YB��7�ځ8lP4$�0��E"O���
�9Xdx27Y?X�H@9�"O& +E(�*,}�$P�'I�}p�"O��a2N�I�$�׮�Y)��k "Oa�ꀕ0 L�����H)���"O,i3Q�^m9*��w���c�jd�W"O�J�L��\�0G�؎��-�P"O��h߸-�*���ą �T�s"O���GFX�Z_�c�@# �"O~L`�تP����Զ2�J(��"O�R"��(�NZ�	�.����D"O��X�O�/�슕��w��õ"O�:�/T� �9�%�K�@0"O����ǅ+d��aR�[�R�؉��"O���f��ά��ү�3.,z�X�"Oک��Àf@�e8�Ob�h"O8a9։�A�a�6OU�y���"O��`e�E.᱒�J�(�� "O�ɲ�ȇ[��@��L
m�~���"Ox����7>X4�TF�,{C<��"OF9j��Z�,0N�!ģ��Z0
Y�V"O�#p)`�v<��H��/L��R"O�yF�0<\�`P��&(L<�E"O  ��6�Np!b˜�	�ċW"O\Ax��S�9�	��C�5��m��"O�Ā֦F�M-0Hb!/Ӭ2��@�"O[xGL͏^ǆ��Í�I�l"O�A#���o�B�	���$��I�"O� �d�D�� 0��FU�Ie���b"O����]֬L �W;|TIU"O�̋Q��<z�t`@�>s�.1�G"O^�g֟H��{ROC�6��}�"O�� 'X9>&��ђ��9�j�ٴ"O�E
ƪ�3�4U�MR�(�DtY�"OHh:�e� `�0��K�K��ղ�"Oҥ�S�+�\�w�/?ӎ��"OzDzŅ�?��"ю׃dd�� "O��sa�ۂ�l�`��:`�u1�"O��x� <j?|e���$3`��"Op���[�
��,y6��*骁"O�آ����@���zĂS��Ȉ�t"OHhRe�T1h���I�B����*O�#�&�B)���"�g�VM�'BD-za�H0[0��qË�WI4 Z
�'K�B�)=��R��N9:���	�'1�=�caC^���UJ���4x��'�����	7d����QkA+�.%��'Æ�C�.C!*�+�e���I�'� �:��9x���+�}3:\�'��]r`�:�B�0%/	�E�Z��'��`J�,V(Q�'%?�ze��'�����!J�X���"�Bb]2���'�J2��!p�Jѫ�&�
��	��'
d�$�ѩJ�<��rO�$�	
�'�5�wc	7�2i�+̾41	�'S�U�t@@�}H��C�I�&<r5S�'�:�B�@�N��-�2�L2_��P�'��D��H��$�b�I�~�RyȎ�2��4R�$m�� �#����f4�"OЄ�w�ٴ4�NLx5l]b|�"�"Ot��T��=K�̩�P�K�Q�t��"O�	�@� > ]j�r"7'�|��q"O���a�6H����&��0�pz�"O��YQ-�(`�P���X*�	�'"X}+Q���pB�2��7����'jqe˱�2���L3���
�'Ur�S�7j�{q@1���
�'S�L�BJ΋Q����p��)}��Ѣ
�' �1vKְDIF�� G�	o~��p�'�黕b�e�I���˱n��1�'��!��mC)g��(�T�3��\�'eԱQ�DF�e����vI�%�x{
�'0��B-�+�2qr���")�,
�'�\����I����u�����
�'�����t8��Ĵ�$@�R�<Q'M�5n@��R��=�(ak7Gh�<qpM��v��&����cO�<���D綅�C��MN>����WE�<�%"O#}̢M��DїR־�r��L�<�u��P�	(�������6�F�<)Rg�>)���%,�x� D�<�͊��R�8��Z#<8��u#�@�<)���%ꐕ�-'=�D �I�a�<I�♜A�^�� !�3��q�Ce�Y�<!���;�:���� �~��x���W��\�ְ=�K�,���&X�v� @E{��O2�Lq4fX�-������/?[h�_�<�G��N�����# ���}�<��P{hZ��&hNu��%��u�<9�J��M�|��P,�޸����s�<ɤ��k�l��wMF�]�*�CcSX�<�#�Y%@�|�Bk���#%��X�<� 2&��	F=F��L)b����'���ޠKQ��9�Ε�_a������r�'��'��3ʓ{�6��4��%IkZ�C �̵�$Q��E�鲗J�;X8~d��쓶~�8��)��e�D��26J��q�װ2k���ȓRTh�F�	��Qn*^��Ն����vC��6������ '������d!�0]h�F�\gZ���a��5�CM���kCO^�r�*��	~�	dy��L�����GD�x��Z"5>�J�#:D�Ш�(I,ry�I��\���$i�9D�C�`_Az��7�ԍ2c�p";D��(�S}kf9ҢJސf^!�T�.D�x#!�٥:"�����"Q�&=f�>D�L �X�\8���ϑC16�0D�|`7��UȰ`E��<l�X)�OC��5e2�(�#��m�!�#��Y��C�	�sk^A�'#K�<:\�g�ٿnTPC�	n\�$�5���!P*�jQ)���0C��:'�4;W�P�1Z���E[\
C䉸.U�5��E��XN���U�2!��=�ç�����3 @"e�À c�}�ȓ/�Q'�۳W(��BTd��	�H�?���0<�'���h���zU╳w�`IHP�[l�<Y���-)'��Da�_����blUc�<��cU�a��8��(#%�,QR�B�	!~r,�u�^�7 ^�ɱ�Y�b�B�	(p�Vi�V얶	Z�qJ5L[�o�B�ɱb89���X4� �)���B�I�%)�8���f�9H��3�	O�h��>( ��뀃�4XG��tA2D�0����0�2�NS���|��"D���Ơ�2�t�ǎ�(~�	a'?D�l��`F�1�)���)g�dH�"0D����o�g�����ΥgL�V�8<O�#<��nŚ$�����а[
-p��SRh<iS��R1&���Ć1_�X�q�
��y҉�,L��ɐ�^c��pp��y¦�,!��\:�$�U#j�:� ��ybj�&p�,0���P����%Ǩ�y�� e7��)�˙[�.�KƪS��y�h#x� !��W�|,��CD�?����(�bE����.l���ڷp�x�ȓ`5Px��K/�����$��GTM��rhT��M̸.SD�#k��n�ć�m���1�
�(��Q���M�\���-��0C�ِRb
�0�Û�UI"L��<�L�ѕ�o������GV�p���	��9�5��ӡ����*U�	؟`�?E����'��=B��8��mh$��J!�	,]F��p�AA+%�Ԙ���˶3!�6"|(��#�v��q`rT
4�!��6�d����:V�҄ؖA�!�$X�GX����Q>,�̚�,B�5�!򤘅!�8��$P�UH���z�!�$�S�Ę �H�S���Ԫʱ<R!�G�a���cG���=A)H�@!�dٿ\�*M���	�*0��H��(�!�D�3k`�j�$<������%6!��M�tQ�̃�Hŵ`�dA�oB�3!��B@���L�
��R���!���)+\8�gn��O-~�%kʊ;k!�ă�k��c1���������m\�'a|�,_�m�I�.�%�#`��y
� R��U	�=Vi�]��.�%9:m��"O��Z��6��D�,��|0���"O±�@��%o�`q"�%@�ؑ�"OV<QЪE?
j�����6V�|Ps%"O �� <S�QaI5�x��"O.Ց���7���Q�힩#�v��"_�p��	*Gbj%����N]�9!��5D'B�Ʌ/��q�MύD`��`7F��#G�B�	�[i��D b$�l��/�B�	l����Z�I➱�NZ�`MJB�I�	6��&S�e�%BWǗ|VB�	;oH�I�i�H�@( gN(72B�Izi�S ϕ�Z��=�D�	bZ�C�3,x\D�2O�zh�qS4jǻ_��C������Ve��d���Ӯ�%J\���D ?���"2��Q�&��9�؁h��O|�<��e��S:^  �g��8#�u�<�󊕀C�y��IO�fz�H�\W�<a���,\�n���'B�Niʔk�h�<)D��.p&f�2ь�,s��P��k�<�/ �ljF�dB�,��+�,\�<�cKݝW����0k
"6�ܸڡc�Y����<c��6@����Hw�r�ϘW�<q���|�\q�D �A��1 �Z�<���&��h3/Y�yI1G�]�<!�o*|[��@�!��+�Jm)`��\�<I&�o�>8h��>��,I�DVZ�<a��[%a�옢nK���و7�U_�<)�a
>cg��Q�	XU�@3E�[x�tExRM�N�(�J�t��\R ���y��ۚb�d�����>e$Y�T�ë�y�"&֬T9@�ҶkA�u���Ü�y��X���؂F���\���R%Q��yrÊ�D��3$�Ϊ(�XXQ���y�b[�|���B	׼���2����O^#~��o�  \����gAzu;��]P�'�?a:v����@���ܗ'��
P%D���<:>x�Cɝ(`�0�r !D�(P�\*��[� ��
j��� D�h����VX� ���F�b�����+D�0�g�vp�SG)ď+�}�ª+D�$��皝ER�)�0�����'h(D�p	��Z��5OͿG�԰u�%D�4 ���� �L�#⊎m��4�Fn'D����	Ƭ	@
��F��"W:tыu�#D�|�w�^~�d��`��e	b��b D��`qȁ`���0@���9�V����=D��:��M�d�V��K�|���!D�����uB�\k�N�8�X8{��2D��m��;0"hy�`���^�*�)1D�<#�`Vf2A��k�6إ�.D��f��-se�)�͊�)���J:D�h`C�r�8,�#/�c��4�cO9D�h�B�Iv݌,�&� ��r 9D�q��F�p>�3G�:��x��:D�xhL"�~$#cY�/ZLsD�8D���g�ֲOI>3��00�@��6D���Aڤ�T�:�X�Ģ�Pt�3D�\KD�ʟ,}ةI ��#<�d�#w�<D�<�0�˭QVpi�&%ӞA�uJ%D��{��B�El���/�
esL�D6D�����5/l@i2ClJ�#u!��0D�8
�O�7<��P��#�&x�}�R�0D�̓ō"pzt�V���~�̥��%-D�� �eg�����2�ð�B��g"O�`A$�,.:t�1��_l�r=а"Or���2{YbQ���0}�DZb"O��G�ޛv�R���.u��*�"O.��'ׇ3��ȆK����F"O��q�!�(���U�I�~pw"O���k��vH����q������u>���f�	����ih�J�F?D�����5��pȲ'J�&8�hSs�;D���i��
�0I�` L�>�:��9D����Y#>�N<�����@��إ/$D�3���e�����a��5�ީ��@"D�ܒ�
�u�0����%�����$D��I[_��y��$�&r��aS�(D�� rj�@2&ѫ��6$F�%k�(D���E��#cvH�pZ6��I���%D���k��o)����[����"D�����2
8p7�9�rA� �-D�tQ�ӝ@=�F#Q�Y>1H��=D� ��B��m,�k�lN>�$9"�+<D�x��ϒ>�z����,:��s1,;D�ȺG�Z&C��+�dܓ����g4D��Q��ѧoo���$��L㞩� c4D����nџkQX5Y��R�X��5>D��S
_�j� "��D�|BA�bD;D���qmC�Nn��1S$�f�(�R�:D���2N[j��h���W I&�p�$%D��(��	� ��J�4'��%Yd�$D�`��C֍�Q$cҥ/�ةЧ.D�8;$-~�.,#�˳/�=�'D����Οa:Mؑ
V>a�ys�&D�X�뒐}D��2u�4P���RM%D��abńQv����!=-݈5�F�!D���dȗ�b������*K	��1�� D�,�"n� ���!6�D�Lݣ� 2D�`�'T	/���e�ڸu��B '<D�h�a��1g����u�,)�\ݡc�5D��
D��n���PUB�<D$i��K5D�p��k("l�*ƪ��@�L/D��y3	$w7
�b/ќ]��8���(D�h��K		m6̺���"�P�(D��;CO�:MO�\*ƃ�H���3�'D����b��5U,�@�&� ���s�&D��q��D �+ƍ�h3���#D�� e۟[���Iwȇ1��mZ5/#D�Lpn�gc^%�3*@1j��v�?D���nұJ�R���ˊ�/�!�D?D�k��5D���#��2���g>D��E%��_+Js1+T1P��܉@�&D��*���79L�"w�R#|��� *D�\j$�D�jhڔ�Tn�}�ث��&D�,�&m�!P�(�Ub��0�����6D��´l.$R����3IV9�P�3D�����FV����/E;	!��0D��r�̞.U���!�E�0HC-.D��BT'$Y�4CuD�6r+dA��)7D����l�/~����U-?�4�$;D��A�NϤ$�����O����@8D�X�Ǭ3�;"��
<Ҫ��4D��kԂR�X�\���KD�6ջ��%D���wk�c��4a�#R�(��(D�xz��A�"3���'EZ�\��sb�*D�`���N3~%�A(u�� x}Xq'D��y#�C�<�Z4�@镻"��e��b:D�� `�Hr�4��h�a��tY�"O|���� a|����˿��e��"Oxe�b���\=2B��|�
c�"O�q��
�r1P�1U凹uGHp��"O���*C�T4b-�>	.���E"O��pG�J�=�D��	Y+�y�"Or��dN��gJ��̙>N"p��"Ob�;B�ǁ.�F@��Jɡ].L��$"O�S����"D��1J�'nP�	�"O�����Y<m�8��#@qp�\`"O�a�%M5A�*y��	�����c"Ob%�c�ӊ���!q��-.�<�%"OH}C�$�
C/*\���Ϥjt���"O�iX4#ߙp�xU��&��N���У"O|y0w M
n8zD�:�,�s�"O�ڃ)^4Be|-�r#�)Z���{5"OJ�8���- �����?�̀Q"OaI�è_����	]f#
�`�"O���F���t�@�paP�+bd[�"O���AH�Rs�$Jā�"���"O�C�i�<�@ ۱"	4�Q "O̝�`iǠy������$��Ա'"OM��"�b���{�G�L{����"Ox�����$(�'�j���"O����1c��hD��Ir�,�"O�Eb���:4w�����xf�)��"O�Z����6ic���/=zV9*Q"O�A�-�69
4C�'�3g���"O�����Z�� ���лPs*��"Ob�x7J1h���q@E�?[Z��{�"O���E3@�Ī�
\�Q.qP�"O:��p�6@�̔�'/НnD��3�"O�C�D�s�5�t@�,~VB���"O"�;�G��QF�!n�.���"O8�#�$��[�R���ʨ;
h��%"Of��G�,��0ul�fj�hW"Ol�cZi� �kdm�4mP�YBH�`�<I+�&Nd����Ԯ$�b@��`]�<�w�J��TIRK^��b4��@�\�<I4S��$��`�B��-i%.VZ�<��#�3v��rD*��c����֍��<��!Ѣ��p����1hhM����w�<����,gHrK���N6���b
�q�<Y�G��DM`�A �M71|mhQG�F�<� *+3N����z��X�J�<Y��E�*Ø�0��P+_I�%8D��F�<��AҢU�h1��<�Ƀ1�k�<A�`W%7�L��D��y���CGg�<���O2$aV��Hdk�؃g�Kk�<� ��E����!��h	�R�e�<)p��.���*�kb���*YM�<�g#�
�*��4g<lz0m�B�<cI�6�� a�J�aE��@~�<��F^k���'�-J+X���bV�<��bCJ�5BB�,p��K� Z�<9�Hυ	�\�`��"l�V�##�Y�<Y��}��y�E�B'�>QK ȌA�<�")��JF���P�]Fe�R�q�<Y3-�U�z���J,	��S��m�<�`�[��R��l+JO���2���<Q��I3�� a��^��܃� {�<�p��I;�!�2��HyKL|E�C�Ir=ڡ�3o	~J$�k4��bAPB�	�`�0�qD2,�`0 
�G�nC�)� �<Rdn ��f��6�V�WO�D��"O��{���5BKj�"��?M����"O���*ݳ���ks�Яg����&"O�x�
x��Xӗ�G�a��u"OPEH7ϒ�;����+�IQ�� �"O�A���Q/P$�$
�P	"O\�Dd�y�y�)��!5x)t"O���,qG�`�H�ML3u"OR�d�C�=Q,|x��ȀLs���"O�Lb��P�c;��X2�VJB��"OZ��S��W@T��f�<90U"ON�p��`o���d	Q�L�"O���gJ0\�r4$Z�iCKʽ�y"�����U�b�~��Ѡ���yr���[��4��.�*C���!̀�yb\�p�h���76��a��6�yB��$�P�:�Ç86� �,��yR�^41�Z� �l� (�����Ѫ�y�%ҳn^j��ķ����E�
)2��C� o�u2��$��������<B�	�4ʚ(�6���6m�L�2��t�B�ɿ".�`���׳ �XKH]E4C� )��J���%^tz(� t9C�	/��E~L �E���@.B�I
G� �+��>���g����C�S� ��$ȏM�T�5�;G�C�	���pq�=�2�)G�H�Z��C��$@)�Ey#��1n� ��Am��[k�B�	�_���������� �0`o�B�I �*�1���=���V�S�Z�rB�I�
�J�8@��"TZ�Z��R��LB�� Q���㗗,.ܚ�b�%"P:B�	������A�Ig@�'��EbC��5q�~�h���*�D!,�z��B�ɶqw����䁅q4�@�O?^��B�I�M�l"��G
$i�5��&7|B�I�?y&�Q����8Ys���'�8C�	�\zҔ�0�%p�>9СK� \3*C�#-�S��ȰM��(P�^ *C�	�\�8�Bb�OJ�=/��l�W�0D���K�$	̺�>n#����"D�PC�)�)s#����%ѳU�p���!D�pk����	�ǪO�nݐ]��*D��J�8;@ ���j�~	a<D��zR;BP����J�?�h�qQ :D�,���L?R��Sr��-!�*� +D�c�g�?���Peֺ:�Cu�*D��@@88�,L⒉�#"��� ;D��0��X�z�CÆ,�>X�1+$D��ڕ��T��U	ţ�VnU�d D��xU��MF�e�Aυ1���"�a>D���7嚴����b��< �8�=D�ԩw˚A/¼j�dI(GyZ Z�0D�,�6�S�C�q�"�0�]	5�.D�(ⅫE6M�PD�U�%��d��.D�"�Xef�C�L��ȫ�a8D���!KTo4H�;��N�JO��u"6D���'o�=!Z	x� 2|6�A)`h4D�������~��p��ݽUبY2�2D����`ߋ"LX@`F�<	�x� 1D���Bg�<Ҙi�Sɔ�6%B�[��-D��r�o�6���"�Ѓ%��P@5f6D��3�f��t,`��M�N�Q��l3D�L2�N�8b�\�	�&I�J��Pǀ,D�� 2T����
��9G㎉� ���"O��۳N� ����b(�6���@"ON�ٓڿk]��"1G��~L����"O>� 5J5lO��#씰}>2qzT�'���z�K�,@�*������@0l���az�g@�9�0	K�\;�f��ȓ�p9��З|K�!��A�[��͆ȓsՐ"����u!ŐS.�:��ņȓJ�X�IA��@�!	�^/Q�H��=ۓ..=��m�\�А�%��=���'3�~�떸6I�Kd���Ao��8UV���d�� �=��c��fb�Z!��4�� �tɅ"�y�\(Re�@{��K�B6�9�۩�y�	Y��jI����@.ds��Ҥ�?����I�<1O�{g�Y����&qi�h��dVZ�<a����3�$���L&)�2�1v��Ty��)�'ah����J$^�1�r�R�:u*��ȓw�E:��Nh*�ND ��<�'��}2��(O�d�2!�	�FnYP/�y��1n1��+]<@���a���'g�{�eW����� ��8]�+���~��)ڧK&��H@�v(�U0�o��"}N��ȓ?�iu�&;$��eY�_�8Ѕ�c���R҇,cZx�0�ݳ5�x��I[�:I�xQ�6Ίe�Ur5�׃r�&�� l�J�*n��OrZ� �V!o���!�P(�E,�&.y�{�F�BH���H"�#RM1l��+A�9-�1Ex��|扏��h`� V0Gx�	��8KڲB�I
V9��#��e�����A�1Y�B��/O`P�4l�E[nI��bC�C��B�ɰl��8"�D�}N�����>=��B�6B+ !�b�5;�i����#L�B�	)qV���(G'���b3&JP�Iq�D:}J|�O��p"K��MuP�����m�c"OT��㚦^eK���+RV $"O2����<?�5�B�׆C4���"O�i�/�?b��jG�J#b�$��=Oh����Y,��q�I�Cw؃�/��!�D�%u�^�����	mb "E`±|!�Dև"7���EF.`����O�,p!��Z;V�)�
�����k�-11��{��h��8TӜ4���V�^V�E�O;8����>��DY1U��-�f�е`nN��j�U�<a���@t��6YZZɪ��P~��'1�es�eO�>���n^>����'ў�}�	n�.)7̅;�V�+�F�I�<�˅�2lD͊�f!�H C��B�ɪ���Pt�0�U�C��}��C�ɯ��D�"93ٺlY�b�h%C��#,{��E�CX���re�<|�C�IĦ����.-���cA��7`�9D�XA�^�{�,�q�к&� ����D�����$�g�:�	����wȱ!d���ay��I�9 ��UFO�|��ȫa�[�
C�	�O�8�Z�+Ő� ��R�ӆCf��hO>9�sJ��s!r�u��$8�!`�.}R�'���b&�P- >�(�4Ň�{�ƅ!�'�
�JÀTI<ThԎQ�u�X��'c`1s�E[�A�����Q8u�,l�
�'�̀UfZ��j��c��Zv �
�'����#
[%|6��(dN�:T�����'��c��;V����!7�>=R�'˴Q�W-G�%�88J��Ҕ5�D���� �0-Ğm��i2��
Z(d���'� � s�CI�6�#(<W�C�I�B�Pu��'Q?<<��A
�	�"?I���V03��	� ցp�hKP�ג2j!�d��`�����1vS"�3�D M��(�S�OI��*��B L¥�CN���lB
�'m���w�ņI�|Pr��4&���
�'�$����/����򢖻|-ى�#O�0�#�ϋ\9:�s�ɨb�ESP"O�u� �1b L@��L5<����<�K���'U���s���m��t�XL�P��$����a���8P�ށvY�����`�E�E�X�:��@��/��l�ȓ �ҕ�'�S)r�>i�wh�&O���<���+#��9���CV�L�H�H=��sm��0�� �f���W#
8�H�ȓO~��{��BW6�	�CBЧ)U����'{��?����i�|Γ\%�1�#�3x�ܹ��x��=��	T�'����w��R��Dac�מ/�:=���.�'Au�}�E��$_]֘Yq�ڋI��?����~�ǡZ���CZ�<XȺ�_�yT!�'u�X�A�d�^�#�D���'�ў�>��slE��92�O�����)9D�h�֢O�q^f�Z��ˠU�j��C�>���ɟeְ�x��H�OS�� D�į`�tB䉗Rpx��BÍ��Q� �T[jp�Ɠ+ �i�`Ć!:4H�&���|�D}�����4�W��b�f���:�4B�� �@]���mp���E�R�q�*B��]ٌ��m1 -� ^�}���$1��s���
0)(v*>~Y���&A;D������C�|�ҟ>�1J#�6D�p�7ʓ%R�������D��A%�2���|`�ŉ(���A��Gb2�����<�	Bܧ ��)ӕ͔1I���������'�ў"}���M�#D`LJ�4Q�Й�Y@�<a���3%�━��E�8_���'�@�<�T�ۮ�ti����<Ubn�z�'�Q?A��S���0&�}Ij�V�7LO�㟸�m�#p�p�qe�ef@L#v�5��p<I� N�y��ذV�.�ԉID�d�<I��յjY$!���I(P�����I]�<�#�S���h1�(8h� ��Y�<��'`�T��L��u@��0�LV؟�<]�1���S���B)[!��'c�I�)�O�$��L�:�i2��N5_�8Q'"O��  �7u~����ڛSgj�Qe"O٫��M�q6�h��ȕ�h�p�(3"OT�r���)�0A�ŀ��X�%�v�i1O��S�g�D�{�Xr%�(_���� dR$5!�t�.�j�f�RTh����8a~S��J�mG�7�R�v响s�`��
"�$&�S�'l���TG��,Қ�`�N�`=^-��IT�pdB�O�R�*��?�腄ȓ([�D	1�O����$m@"���}�l���
����c�t�Zm�O
E1D�kC8�p�*[�e��c�"O�	Xg��+[(��ٗ��mR�U�2"O���@C��LS���C,;q��;��'����ha W&pk��P�T 'r�8S�,D�xx��/)����L�nx�@���*��#�Sܧa<�, Q䕊u��J�ʆ#ӂ��ȓ)���kSNJ�)��i��>�d�Exr�'* ���/�9�́�2	DE�
yX��� L�R'�WU�,bt���cyR����;�O&���'��u��F��>K�;���7I����'!4-�2��UP��@��A��I�'��9G�\~M����'
�f���'
��!bL/}rL��R��`�'�����)��M��F���.�C�'
T� �8y�8;���9<Ӏ!��'�p��@ҏ*�Fj��D//�pb�'�Ĳ��/4G`��J^4V4b)0�'�J��6�	YX! � _�4 �'ݐ �r�ɝF��ಮƟT�V�a�'���p�q�T�"�˫V�0(�'�LQB�UZ�¼���M�lq�'ju�A�[<fM0#��E��$�
�'���ҊK#}d�W O�O3����'�詠w���l���@��@��$k	�'�̑�R#P3�l��ln� �'Tf}c��U�vi��
`���R�'a�A&8bu�EM�T:�P��'tƉ� �S9qS�
,U�J���Z
�'�8ź�ؾ8�TI{�+�H-��'�R�f��zV�C��
I�$�
�'H� �q�$V0��� �J~s�`�'4�-+��&b��ԁ B�|��}	�'���"�ޟP� �'C�/n���j�'N�-6�߱x���J�k�|P�|��'����G2Ive�5�ϠupZ�y2���ElԼQD�[En���&P,�yIM��m�$|���h����b(��'��P�/X<������S趠`�'��S�D�7��%:����F<ȸ��'�D�R'��4�b�XrM' ݇ʓ(�����G�O�}ʔi��XB��ȓ~?L\YD���jE�-�G#`P�ȓ�L��`��J fA�VFW�.D�@��-����'�S��9�Ո��� ą�َ���"i�D�.
*d�ȓ50(�Hc�9S�8�Fa\�qZ���Y-���pjNXO`Գ�
Bn#��ȓZΙ[�lB�96T�d�"	D��ȓi��#1��K�����mӣ3��цȓF)��2���m�B�cFB�\��,�ȓ;ܬZ��Пfp���LK����ȓO�Ҥ��p7}���W�J��ȓ!B�8D� m����.�i����ȓlא<�+� N|F��b�S���<��d��"2
��XE��9(��Q��=fp����_i�(��o��~T�e�ȓW�ĕu�'s@��d H4yj���bʼ�Wދx���3"e�6+[N��ȓX
�x!�"1b�@����GH}��}�0��dM
�x��w��5����$l���f�Q��f��Ng6ć�&-�0�Z�~G�p���S�O2x�ȓ4�����q���0���.p�^��ȓ^���C�C-'oh�P��&T���ȓ���!T�Лi~F����C�~�,��T܆ �ʃ[^mX�d��&a C��&s� ��6m�.�4���1( �B�ɬ3�F����4g~�j L��[�B�	;@��`r�%�������-y&�B��_�Tm�g�E�@���*�'�S�DB�	�zxF�Rcj�Ol�k���.B�ɪ=�f פ�/��\Z�f؜|��C�)� �I�t�W�uq��.͆�y�"OA����b�VHq���rm�"Ot��iZ�L.�JwBO�)a*iȐ"O��C�ڧv� M�@�M\P�<Ʉ"O��!aLuJ�1�0�?
�,M)%"O�lc�N�-u�~��s� 3�P1�w"O@��D�c�� L�pHq"Ob(��m�j��l�4a�&JL�u!"O�����%�r�N�&9�|{@"O��y��F^�$9W�	:N<��"O�Q%��|$�P@�)EN<�U"O�|`�oI�{���@�D�,;u��"O���:���g-��T��"O��z�
H��dXp��j�*�a&"OX�㇣�+t�mP5Ŕ���&+�L�<Q�*y�JĒ2�X���AA�y2nȹ[���"�><�&�y��Ӷ�yRk�
����14�����y2��#W3Ri�@�D�,�<���P��y��T�wX̙�E�a��#��U,�y�$^Om�<�f�ґ&K��J�U �yB��.Ӻ0)�KR������yB@ S�.-bf[p�0ؠ`�G��y��"���Sb��%,0���y��<iY�`Ua˄��ڂ�\��y��.��P�ƒ9d�e೧�y2 A�
'�C5A"����L���y2�֛l���c��N�@�@�yBLKc��p�B��nq����
�yr�L;p;|u	2d�,p���jQ+H-�p<��e�P�s{��Y��Vb@v��y����@�꼳�*X��	Q�X�N<���', +S�&�)�'j1B Y�E�8��YQ�-Y�F�A�ȓg����1��h���⣂�V�P%��#���/U���ף8/����	{�va��oT�u7�RC�!?"�9���I�՘�@ߺ?�4��e�Px2+�C���xW��"b<J��'<��O
�C/X�q��Dь�X4�§��+`�(H��"O  ����3��Z��´��heR�d�GK̈�Pb��|��?V�r�p"C�7Y�B"G�<�I�1i�����'m����J�&i���2�'�jr�U@jV�!��F/���'�^=�1EA�WB�(�#��D�P��+ ��x�@�:�B@��+�A<�c ����y2��Q�� Ӓ#��N���m�y���*I��Y�S<8�&����¬�yb��9���`��f����'@�y"�,:nbyҁ�!/k�����$�yҺ9Ю�XDĥ��0Z�a@�^!��DTؼ���L���7�C�Mb!�d%
x
�؆�@�]��|��J¡O{!�D�{s&M��#x*@,��׶H�!���(7�ʶe�?�����B�!��0!Z�g8b�"%�%��5!�D�?zh �`t��	\�!���!�D��|�����J�Q�8 �ā2t�!��!v�F9X#�F;z��*�@��!�d��"`��Y�6�I���!�$�'�؆&���z�䑡s!�$N/� E�K�9%{(0��e�S�!�$R�O�QGT�2Ǻ�D��&B��а��n�=!����d�88�C�	:X������	"��C�s.tB�	�Z����d�C3h�
�Hu�e�BB�)� `*pA�d��}���j>i"O�]�!�Ĥ@R��!�FHIR�"O�`��]:��IՁثn(]�"O� v6S����I�IG"O�5����� ��Kgހݼ�H�"O�两�پaj�4�ğ���8e"O�IH�E�b�St�T��qRv*O������b\���p 	�Yb�Q�'���YׄZ�	o��
�+��S�x�j�'���d!�=m�ia��E�+fk�'�V5��	UeK����J��Ʊ��'2&�p�)�$T�3&�G.	�L�@�'b!�Bٛ/�h5�u�.}�( �'�(r`T�rB
�uċ�s!�L�'L��22� ��$zE�F<|4rH�	�'nrXBAdO�^V�ES�v�2Ey	�'�uJ�A�=�Ṇ��Ѵ'�P:�'��0�� D�u�r!ɐ��'4�Mr�G��i��]9w]D�4���'��9h�յ'�hy˦�@G���
�'=jL�tY�dx�3 �$5�q��'N��A�F�H��M �ʟ30�I�'z��B Y�q>ȸ��\|��@�'�
4�æά?�`8�*�<��'*��g���3��ɀ��>{�N���'�p!�(�6>q�����f��m1�'����ԭݣ|�(i��2S���K�'̌���@;v���i�_�T��
�'�D|Hscؕo������C�L�L��'�J�[�j�2K���A/�,N�pɍ��/���F��$�,� ��A���N��ybF d�"��çV��2m�-Č%fXfl�:��	�Q>˓S�pd�,)
FD�ӄ�J�̇�#@���EeF6������W�X�;"�ZQlp[�o_8��=�'Q�r0ڹ� ��
�ԕ���Vix��	Ǡ¶	�ډ��j�)yc�&NFq�<���Y�dF�Y�%�ۛ�y2���ء��o� 7�J�Q֭��6�B�iV�	
e�� `�=�'q7�y�$O��(�d���8hr��ȓ򉛦�K�]J�Q��ӌ,��=rA`:m�������O>��R��a�g�I�6���zr	U<�|�	V�F;�B�8<F|c@@Ţs�����'�+
�$%�2G�BbGKZyT���	�Ti= ����7�(�HA) '���D��ah�-Х�W
^|��j͠[Q��C⏤>�U�5�׿J�:\�ȓM*�L���Tݹ�H��U&d%���#�`�p�r	�J��}D�$F�/*�[��r[����e��y���"�vIŰj���)�5%�֤p�o�c�R�IS�>|��L<)獙	H�-�"!Z�;X��P6��TH<i� O D�f�A ����!#*E��dA�6j��@"K�(�p=���W�jC>Eb��&pN�T8$i�`X�x���e�����4q8T��H^�U��"�����sgͱ*�Z�'�:�!��>�!�m\����H>1��܏��쑰H�pz�"}:u+4c�k���}_�KV.]A�<9DnR�/,���'�8J��r�@
�@�(�ȲA8���V"�?�'�4P���Xe�H8��� �U�� �'<0)s�jS}C��K`�R4q\��CS2�<a�gd�7�{r+L|�@��#��!|��s ���p=)��`�Lj#Gx�L�u
T�+0�;���l�����!9D���JƓa��V�@R� �`2�I�dDj���G'���&F"����נ K$C�� y���j#h��J���6�-u�
C䉈ZLps�4��mCBf��n�"C��x?�a��I\�H����h�cC�	&���7N��fĸ}��	�(��B�	�a��J�!۟UTy{���%k$�B�)� �Ŋ��̑Z��cB�$G��A�"O	��陙QR-���W)M0<�C"O@]�1K+$@�d�Z-�h�w"O���d�16a��cD�	Z`@�"OVI�D�I���"4a��,���"O�����?>E����+1�^��""O*�k��M�GrU��.?ˠh��"O�e�hE&�Hԏ��kA�u{q"O�q�Ѱj�IH���L��yw"OX�r��Qm<��x���Po�V"O�ĩ�f�w'.��T(Q�S5��D"Ox�@f�޻O�sg�D�mZ"O򴸐��(�"I�r��d�h2"O�3�h�(3S&8�ĦBh~� ��"O0%�W�@3�p{���*"2l�&"O�%��	R�\�Qb4䆢~M�0��'����Ƙ�'���2��
�L�'�n�Ac*=dP쨐C]�*zjXh�'�̼�&ˢJbԑՋ��$��|	�'���ʒ�T���q H�)
�'e�X	�ʏ�sUR�`b
F/Ё��'�x��S�n(V��р��x����'��=��
!Y��i�/2䵫�'Պ��E�I�Kk�e��&#�2)2�'�
�p.8�l��&�����'��X����~^��r V�E|M�'F���"W��tHb�B!�0�	�'��V�m�1�A��\����'L�}
C�.}��	fM8]dA��'�����X�:ժ��ѩA�Y#�'�l��I̭x8*��@��qe����'�T�0�N?Q)��{d��^�Z-C	�'���+ W������\U�a	�'���{��:c�2�k���
%A6$�	�'bJ���`C����� ��6Sb5��'�� ҫ@�n ��Zª�,*L��'p48늓B��C�%^�� ��'�p�㠅��vV�)��G3��[�'6�:#J/Xv�B1,.���Q�'���d�;>M�) Gү8�T��'�Ԫ�l�z����){�ĵ@	�'�D������H ��0Yi�0 �'���;��*�@� �:H3�i��'�α�WAF�.Ap��5PA�Z�x
�'� ����@=4
�1��@:D�����'�u��4p����ڱ�4�Y�'b�y�,ʃ#wX����B4�'Zh��%Zk�,2/�	$�q��'J^D����-7*D]ɔB�=�
�a�'�(�0._N�<|������9�'U���7[�P��V+R&� �'J�hJ��˱mT�E��_�"����'z��a��	-��3�ɀ�xl�	�']��"�ߙ0;ZqCBL�H<A
�'et��E�_�4�. 0VSy�H��	�'��ݨ�m;�vtdK)-|Ձ	�'^��4���s� Ȫ��Dvc��Z	�'A��+r�A�7��EP��m��%)�'�z��f�]�Dmt� ���ؙ�'$�TI�//T+G��P�&̉��:D��2�"_�<*�Tjsပ*��X�@	2D�����[6�İ�N�!|�@�,3D�p�@%դd��`v"܀[��8pd�5D� �D.?y��V3yVd|���2D�� ����cW	򨨣0kY{̪��d"Ot���V;C5� E �7?�nx�`"O��@U��:+��@��]#Y�Nsd"O�Q��^�Tb,	DY�߮���"O�hz�CV�B+%��A���<"O���ŎN�J�NX#��9S��,r"OU ��?�&H0��9��|A"O<��$L�]x� �X'
�,�a"O꜋�H�Qu`���N����xv"O�U���>v�lY1���
*�4�"O^[�iܘi��W��L �lB�"O�]c�Ä1u�&���	Q|�}Ze"Op��
�Jȸ���G4�!�g"O�q��3Q�X�SB�/T�(�"O�� ����Y���X1N�I�"O�����Ӟ'P�|a��͚\p)@"O�P���8"��4�
� !�b�rc"O@�ˠG�)	?�M��@�3�
���"O�4�����EAe�T6Ȅ�"O�q ĭ� {�,<)EoQ�<�h��c"O�e�Qo��#yZU�ul_��y��"OL) ˟�i�j�WI08I��Y"O��X���M���b�5)���a"Of��t!��C~��`ȇr��@3G"O��A�.�c�DAɆ��R�(j"O��S!V6F$u�T�E�<�
�"O�����I*n�@4j�f�2���S"Ol��+��O2�=�� ]&���V"O��$�J�M�ms��v&�K�"O����YRp�� ·$혖"O|@0E��Sǀ|�7N��R�
e"O@a �o53�Jͻ�`�[Hö"O�=�����&�jqDLZ����"O�u`2�P�A�BY�aB�&&	R=!t"Or\)Љ�0f
�u��y�����"O�ģ$�̀J��JG�I�4�V"O���4���<bX�IY&/<��"O�)@1G͙X�x|#�F~#�!8P"O���֛o����k��;�P+v"O@�K��� @���� &���Q%"Ob�J���*l�i�Ǐ\�;�^ �"O��Uǁ�^���dNF.}�rTZ�"O٩���k�Z�'C�R�Z�ۆ"O����g/c����P�ؙrf"O����8|�TXĨH�D1�Y��"O9�e��˸�;%G��6��U�"O��1�Zhl�rs�_�G�~��"ON�Q` �V�h�F�.�(��"O�܀��ڍtJ�cM�p���	s"O�9��8r.��z �ǧu���"Oh�ɰg�:0��4<I�"O���#�P�Z<U�� �|��!�"Ofȳ����� Ԋ۶<Е�"OVAyK�pR+�c^'u�8�x�"O���b�_�����L_
���R%"O���&�V�o\mj�ŐZw$���"OL�RK͟3�4�����0S>��"O<i �@ɲqP�`!̙)Iv�e`v"ORP`�e��}l�'��7ci�Ɂ�"O��K�#G�/��Qc�Df�[�"O� �Q(^�%t���"�2�c"Ǫ����;J������A�]�ȝ�0"O<$ � ��[�8�Kf�&��U�"OHl
�CO�F�BH `� �K�du��"O� ~���/��*&v�R��y*�@U"O� �S+&���SU�,oj��"O�mb�� ML�9��D�l�$�W"O�|����t)J����w�X��7"O
�	b�#Z<^4�P
N��!Q�"O4I� ��D长bĘ*2"O�H!B�0]��y��ˀ-:ċc"O
L�e�	=��f`��R����"O:��Q�J�X�H���e�P@�0"O25J�j�E��	�4D�d�X�r"O�@B!�S��T�t�+=�^�H�"O�Գ�*�(�RV�:P�2
4"O�@0�ӀLc�"O��f��Y�"O,�a�!X�{,�����%yg����"O�͛���W�6��Ҥ��{k@���"O��{P�<s����6���@UX�#"O�Q"㘢 %�E���C,J���"O���5C��_N���'=4(yv"O���w	ݟ]�,Z��]�t%��8�"O�djؤsBrl�U������C�2D����-Q�l}�T�^�P&��a/D�X*b��=:VlQ��6O��CU�*D�L;Ɓ �Oz�%`�t�^9(��*D��QR�ݲ�N ���ox����:D��1�)�}��x��K	+ld)`��8D��Ztf)sr"d�f�ñm^�Q�F9D���B�V�I�-1�d˴}�X���T�<q�b�=<J��V Gw�m�Wbe�<���ۅu�D�Z
�,�2@��e�c�<�c�ݤ#�t�#��Gm�)�#�\�<q�k�^i��3�E̤@�|my���a�<�/ܸ93��	�|T�Ю�X�<��߆J�`U8q�������m�<��k:v�D���M�aW� �wMC�<�g_=|4je�ۮT�1x��}�<Ytm�	K�i���/	�ݣ�O�z�<�ǏH	(f�]0�.A*)o�̸TOGw�<�F����3g�I"09)Un�<�+��mk�鳆v��0���a�<9"��[�b�p#&��C��1�f�<�`�Z�H��"�#�Ru�@�`��<�W��Vv
�K1��=��|x�MM{�<���^�A� 벦_� H�;�n�Y�<iP��<	���R���pG����XZ�<QǮ�<���ƣd�4�to�<�t�ӏ$�� YR��2?�1;@�d�<Y���+R��
A�P�*b�
�(�a�<����6�@G�}2�4��d�<e$�[�*�P&��zLI�)b�<�΁���ISj��T�����g�<��fȰ#i��h�*�)Q"1C#Fz�<����gx���-
�Z-���~�<��$ыUq�]���)a6IH���~�<�@f-*��)M�����t�<	��ߡZ?а�mT$!ґ�Wˍ_�<٧Ι*E�Jy{����~:(��Up�<)�c)�L"��ę^��p�f�<���Qo*�.�0S@�ޟ�t8�ȓ0�A����y�btJ��P��ȓE!����H)uf�rI�=L��ȓ4�)��$zJ�XQ&�"w�؆�-�H�ʴ�U�w�R B�.�ڵ�ȓ}�X�'Ez*���T�܄C[�Ԅȓ=�x(�k��rvغ��i��S�? (�(��bc�@�K��`}F	�"OhX��%ىEBx@�6k�7T���"O��"��R�LcT���+J���"O4ȳ�#J�wQX)��Y/+�$��"OF���A��=$�a���Ƚk�"O~���y�t���@�,.:�8F"O���m e 1�%4d�@�"O~a9u�K!P��i�E� ?�R=�"O \���;_r����Js�"O�qi�+B-����<?,sV"OnQ8��ş�$x ���%�<"�"OΤ;�,h��)V$�ua#"ON*��v��eS��K��qP�"O���g�ƙG��I� ��G�֨
"OD�jѭ��Dd<��!:�^���"Oi1&��9\0���ؑb��!k�"OZ@��.G�\+�!�W�պ��M�"O�5X�&�.��X�N�v��xx2"Oz�H����,8W�4�|�5"O��C(?e�hC���s	�܁�"O�4"��L2D0$��u
Ш2^��S"Oj�hA�КC� �ըӹ��!
 "Op��!�7o�dq'Ґg�j���"O�mXkGHa������H�Y&"O��%�W�sV���$]���l0D����Ɍ�3�����#N"��C5D�@��
��y�=�6��7J<�0�5D��8s���-UH�(4�5%�ԭ�f0D����*y�a�*�"��Sf�0D�pr檌�B��Z�F�qp�.D���� =&\Q��kU�S6%�b9D��
�ǃ,pHth
B�ĝ|u�h3D�<�r�S�c�Щ�q� �G>�dC-;D�0�d@��8�Xg��'�4$��:D������;M�� ��B�XxY�R�&D���G.��栐Uo��*��%D��a�΅�F�T�2/��Y�h��,D��k �F����"0 �"��!D�,�V �)D��f n:���;D���E���Y�\��@��*|M��K;D�˅팋%R���dOˠ)`���7D�\S�+�/Bj�iE�F�l�n]1��5D��(��ݿP�a�$IWe��F2D���DZ#9�D�k F�9H��2D��)��2�f9�`�.x����3D�@�E�H���g��M0Z�ZG�/D��	􂉽)�AQ���d�R`aҀ*D�d"��+HdzeKDg��-�$�H2�	�BR��T6Ot�Вi��M'?��|J�Y�<��[��S�|,���@�T�c��F{J?!XT`�,<LJ�o�7�򼃕�$�D#�Sܧ�64:Dd�	{� y�FDf�~Y�''ў�|j�`�(n^*N����e�������NL򄁍9-t�Y�(�_���ȓ%*C�CC�r�	ۂl�N���?����~�$��z�ج3�	*f�и��FY�Ij���O��8�$ޗL��m�
R��Ȉ�*O0�=E��5` ��Q#&0�D�iQÙ�?	����xr

�*�[������G�h�=��{���H�ZՈo��Ȭ`���-@��; �Z�%�H`P����h	�L�� ԛf�DF���ĝ�-��cKS�.���JR0f91O,���j�渧�O����	�S�$8�	�U)��Ћ��p��6M���%է��;��?��G�]��Ja����=d
<	�#�)z����T���D
�ħ��O|$��#D̴98�Tq�Ū�gB�y1@��'b���VM>�+Q��%�$��` f$��P�<D�I��ڜ8#IJ-a�� �9t��-`J�P�ߛK�ecr1O8�
��D�5���t���M{2�>����M��I��N��H(�'�"�\-c$��O����4�̈́"|`�(���<���h�|�2MС/B��a!�ʌ/A�/�&)��2D���pٴh���çJ)��8r�_ˤ�@�cձ�E����#�,���l�T?T�W�Qd>����, �=��Ɂ�>�2MC��ϡi��
P,��\���C(�����'�����8'ȠBW��D��)�Ł�H��c�L�t��DAt��RZ����C!�!��\1��I2姎>h&t6D��?!2���I���ُy*��	�\�^��HB>Gg�P��N*k)0C�ɶB����M��z5D��w��W�&C�	�n���(��q��D�Umm�C�ɘ:� ���i�)J��S%NT�|>C��:<b�e�E�9v��r��	�C�	<]�ʨ���O:	��8Q�o�B��C�^��52�&�KpvahS�E�_�rC�	�kJX8j����DZ�`2�ޕl"C�I�`)= ��G�(�c�#)lTB�I.t%�h��N�+V�TkG�G9q�:B�ɟzR�P[�
S�CV�PɅ��<E�C�=��}@��	5f(v h 唯e��C��3_t�A���!
�`��,;}��C�I�3�t���	dQ���K�m\DB�I��\��XM�tx��7�>B�	�/#�0�4�' <�k�>��B�I�zZ��P��կ|��$JQ�)z�DC�	f�8 �Q��85����
X26)4C�I�3������4Y���A��B䉁��
���R�����U.�B�I�R&�4�TOJn
&9�2���+O~B�I
V�h;q��$�.��A 1��C䉧J��I"&�C1'��bWK
�R,B�I�*a��D�
����GlC� *�ژ��lW�@�x��Ƣ�R�:C�+o��x���!� �s#�i�NC�ɴ:a�uÁ�^^���� &U�~C�	�hƎ��G��A��9�2�@(��C�	�V�$j`�Ol�Qꧩ_�+��C�ɥMf!�҄���I�C�"�C�	N.^���
�*�x0��Z
>C�I-[���iBa��?����G�`R0C�ɞl�h�XB���i*�� q����B�ɥe��h"g`\�pX|4�%N"|��B��9����̏ �z§��	`�C�	(	Ş����^��%x�`:,C�	 �p9r��c��\) HK"+|C�I�D��諑�D�E��[�j\�2�B�Ɂ@b#��61��T,��aW�C�IC��)���y����e�6t�C�jC����+�~i����v��C�I;yl�ڱH��v�j%B���G��C�I�1��I`è۠"J���g���|C�5'I�a�����A'?G^�C�	:x$��đ& �ţ��զv�C�I�"7���t���?-�|j�#J�0C�f呖�W�:�&�HצƘ[j
C�Ɂb�����!l�\���X�o��B�I�`uά��b�Z��i�-D?b�B�ɖHu� jJ2�uXEdB�`�nB��&}��P��C�*�|)0π�U�B�I�bLٳV��1^�Mҵ�^<L��C�I2A>��t�W�ᖉ��5oZC�I,B6�s��l\�8����C��4��	z!�+�)���Ĝb�C�ɘ4�V�<eP�P�iX%<T��'����p��&�5�D�
nL���� $�P'�;j�y@�ٖ	��	��"OV��A�[�H�٢[�7�xp"O�[�E˟bqj��1o���i�"OfE�Dƀ%"��Y�/u�ة�c"O�m�Ҏ��?x�s��زN�T�s"O4� ��]�"	09a.��)"O2�:PEN�^����q+x�f�a�"O�CP��18 ���6K�5P���S"O��EN���"�J�;4�y��"Op-j���hd�-�`�ݟR� �p"Oī҅��<����5_�6��Y��"O1	�B�?YY�#!��1Ӑyb"O��qF�ϒgF�h5�?���u"O��@��܀%̶ѡa�O5V��@;�"O��@��"$�A3�怢}Z ��"O�A���9}j����Ȳhln���"Ot�嚧H:6�8���0T�1�"O� g%
�x����nL�|5r0C'"O�G>Y@h`�b#T� �P��"O�|򔎆�Xh��B7B�'2J)1d"O4y��F���d��!�]�Z�"O�cWF��?*���4Yj%�'"O�y6n��5Ȍ�CV�L�$U"Ol�S��G2�0 �E�gʘ�s"O���^7Bh�#Y�+ pu�"O̤{�Hԥ;�Ա���V5��́�"O�$���	����6P�\4��"Ob�R�[>XΘ����}�Ɲ;"O�ɱ���F	��S���%"��"`"OL�Ƀ���y/2P�O��/�hx��"OH,�K
�]�8B�y �c"OP<�%Ɯ~�p�಍�1�8R"O��"ϔ�.�V��Fv���"Oz-z1"Z$r��!�$ #j�Z(sW"O�Ģ�iQ>l��5�V#мK�r�"O%�1͐�{������W�͋�	�!��#S�`!k~#�Ux��<O�!�� �G�0=9�&pne���;')!�_�R�)՟#�:�Xw�Є<�����'h��RU�[T��5Zc#��Dj�)�'�0p��m� ӓ��o�m[�'�P��W�{�Fk� Orf�I�'0�atk�B(����\�4�0�q�'�
]��h�R��G�3'�앃�'wz ��B̎YP� �6O�N�}��'$��[b�W	��IH�!���zL!�'���p��ע������Ga�'-b�A�.Ȝ�
P�=���o�!���<������?� U�r�@`�!���M���Hh�~X���4�!�J�]��V��0�|�J�l-T\!�Dt�6��}j�Px���	0�!�d�D�n�XK� U(����h�!��Q��T�R6��>f�l0qMV�g�!�ė:>�r�`��Zq?�<��ք2�!��̤R�ʒD�j:��QE䏫'!�=h�©�gC��2�q��a�>c!򤌀2`�Ti��?
 �!�X�!�T71��|k��Ȁ��ъaC�!���J+�M:j�r�&�ïL�Ko!��C,Pf�a�eU1a���4��6�!�t.L%h��N/���a�܂�!�
�C�r<� +�<�BDӢ�~!�DT6*��0�JR4D�")�bd�D�!�� �$���G�m�0���Hz�N�I�"Ov9�5��=s��#�a�3x���"O�PKE	.@��Y �LIi�8Y�"O�@��Ԅ�u�a>sg�y�b"O
��a��h2D�ᒯ++����"Oz}�qA�,x�f�4��EpJ��"O��:�R�e�3��H�	L��E"O����m��>�	B� V9zͶ͉�"O8� S�{��5WQ~���"Op�s�LXA�gBJ�"Q	J�"O�@Y��+;���I�j��NJ~JT"OzU��N�Fe3�ɖ&�\��"O� ��-�-M_b�3Ũ��]� :�"O�Ƨ��[��Y�E�f�,�b"O�=���a~F}1ց�wj$3"Oj� ��/;���"T���aD�"O���u.�`㔘"p/(^���"O�i�b��2��CW�ҋ_��e�"ORPHB�Nt�	�����T��iT"Ov, GiX�e�v�8�U$����0"O�THw���EP1�w�2gu�Q�"O��ࠀ�!0$��N�*(���"O!1��<A��hh-�/cJ i"OD�#�HC�h�ɀ���1M�@��"O�eu!W��,��K��iD�]J�"O�3DY"%�qq��	(��A"O��Z��%3���h��ԷL��8"O ���Ï$��SK�� �t� "Op�1�NM�_C1�&*@�?�� �"O:�QtI�	xS� ��ˎn�ڴ��"O0 �%�Ҩ;�����G��и"O������FE+$`�	D𔀋 "OXy���T�9$ϟ5I���2"O:�����[4�8��'Ep�:�"O����܇cL,����� JB��Ц"O����I^4�M��˺W^���"O�U�6n4UJ�S@n�:MEd�R"OD4�f'¾o_��p�K2.4"O�8r��E��d92F�p�b"Ou�%MZ�X�$iӤ�>���0�"O:�;7OO�Be����M�~,"ON�[���Mk�m��, ��]�3"O�Š�FN*�*4��k��(}�m��"O��B9}� �k��ԉ>{��Y�"O	:���|V�l�3�>PZ�Rq"O��GC�(�,�it�i��2�"OƵ��"4�,�q!.c��H��"O~�����
/`P)�\�0�lx8�"O\q��K�~�@P���]�%{|���"O$("!��q�x���#o�� ��"O�}
ca��T	`�c�frP
U"O����,R0p�$��Y ��"O��K���#w��c��ƽR�p�"O̕8fIЌY!tU@6�Q$ 5�!�"OʑQ�X�~tޱ+�b �=&�0"OER�Ɛ�����B&2�8���"O�x��* u�X1�`� t��0�"O�4Q��H[=�h1$ ͱf��1C"O�I %!ע�
���8Όas�"O�\�$MWToBx�nծA#dQ�F"Oj�;!���D1���,'a�*O�Ɋaۃv�x`¥(�$<�����'?jӱM�\7¹ȱ"8H[�8R�'SB<��Æ�}�Q�/� A��8��� B��)zM�D�C܌1pt� �"OJ	"�b+�(�+��1l	��"O"�pҠWF ���PC3tZh)��"O���ѧQ:xp����뛛v@�$sq"Ov̺���H�����4+�I��"O�%j�[|K��R��Ů&��p�"O�����mG�4jC̀�&��p"O꬀�;'�l�ð�V�a˴H�E"O����/C���%儬gQ�"On$8�,�g(��E�(�����"O,i��k��8b��� ��H�"O0���V�N���I��1S���0"O\��$   ��~���K*�y4iM�)���͑����I���0Ҁ���"~Γm#�tj��+�0����ò%�|�2�]�v���	��,3��3�3�	V�`��IT*j����C`X�&�	�
D��b�Y~��d{$�	%a��X� 
M�$�v*ݗhZ��6!��"�ҠDR(!'Q�|�b�U/*�杭3G�Q��m
'!Hĝ�7�K���8w�	�X_�q�L̉?s���0�Od��A��6w�r����I�Y��@���	�9^d��E��7r��~��kC�G��+#�S߸T�P-s�D4'�p���J<&�t"����]���Jt�V4{�!BEu�<�kB	���cf�Z�?V�e�V���ȓ}*<�S��dj�)'�ۻFͬ%��?���� �¿F(���R�_;R�(���"<l䨃Ñ3:��Ì��^P��y��D�CW������D�GX���ȓVDxa��
�_x
Y(����4��ȓc�v%rA�&{�(&-�S�n-�ȓ�����#B��l����y譄�S�? ���hQ�y7M�+AWL�IA1"O �r0�Àn��tK%
�8��k�"O��C3Y�X�R\�s�!V>\l8"O\rW��4�t�c�ѓ8XL h�"O�Rgȑ�w����ʞ�=�^�*�"OX��.� ����S+ĳ����c"O�J����QYc�Æk��$�v"O�"��	1�(�eߞo��"O���4NX�h�e���O��QQP"O�5R'�T4%"���*t�m��"OD�D��Z�6t��)��i�"OA�@�d�������
^��`"O^d�sLH�&Ą�Y�K�9k��P�"O�x[���_<$��9T[|��1"O�B MZ�.��I��I��ER�U"O~8!c�O
i�B\[3/�#pCd�3�"O��*�)�ٷnK"z$Ω6"O
D�c�C��-�0�s�2��q"O��Q(� y����+7��h:�"OL�����"��$�Ȍ�Ml" r�"O,Q ���!Z��a�"O��7K?o��`R�:>��"O��f;]�x���TO7j9�E"O$X�%I09	#�[�"U�q�@"O��ikʗ2�y�'���]n��#"O��ᣥ�έI ,F�,eL(��"O���R��LI;g�@�`^� �v"O
Y$�Us6��,^�[T�V"O�-�w����=���S�JV�@ "O|qk���`�^eH��\;<�4�q"O�Xv��'KD	ɷB�9�N���"OPA�F�~�2���A�.3Z��bG"O���$B/H)�!��*Ё~G�=87"OQ��hմ2#hػp�ʡb"Qk"O�عe�	�B����e�|C��"O"���R>a��QBD@;�I"O�i(��M�S�5{� C"*/���"O�!C)$��@@�>'*�y�"O$��lQD���&a�&��"Oz@;��>���t�\/h�LkB"OJ,�rK NB�Q)#��15{��"O�X���G���@�K��l �c"Op|��G 5&�ibj��.d�[D"OT�K0��x���R�C�*�e��"O$� R⋩D(6�
C�y_���"O��i�jO��<;ˏ�sOT�P�"O �sAԱ&�P,Չ�%S!Fxi3"OPty��ɪ)�
���܊� Y�"Oꅫ��n7|��A'G
��2R"O�=��0A�Q�B!����"Ov�) �Qr�d�Yp�	��z#"O�)�sG�b>hp@��J	���"O��@�Ӽm��	�oY=�t��"O�1ۀ�	
�2�s�.W�l&y)W"O
4m�^�K΀m	"f���s"O4���Ŏ0;N��x�i_
!���Q"Oz��`a,(��X11��s��<0#"O��/��z���kY�[�+s�<Q�FG�|8 ���1v�}
%��n�<����h�>����B:V�th���g�<	���&!�E2�C�T��;��N�<a�$;#\��	�A��FMn��q	�f�<���>a�bŘp���/N<�R.^�<!�LG�r��4�����t�S��W�<� l��h�' ����ܤ`�H�z�"OԥxA.D35�j�$a%/����5"O��!�fQ��z� �2e�<�"OάAVMU4"%Έ��ZSn�"O\��ڎ?k� �TMF�7�T3B"O�x��ϧAX��s喴~����"Ob�ybǭ��Uy�m��o��۱"Oxh�&���3�hA��9	��"OHd��n�זa�¡�X	��"OtjFV�3�>���!@i�6T��"ORY�7G7Q�nE� c���V��"O�E0&MZd���u��� �\���"O �X�oǅ��D�4��~�^��"O\�
�^j�k`�ŝ`���!"O4���ӂ&gXA��H�G����p"O,�uC��5��|��욲�N4
������B&� A��~%�I#�AJ�IfP�>)��)��]�ty���*aNG�-K�!���"�La����lo�%��"�yC!�$^�O y�� �7
ɾ�Fa�&q[!�DO� |� ��a�J�G�U3t31O�����t8��u��~��I���[�t!�בLP�<���	!1�N���,�C��3(H0B�V�sx� r��=aT�C�	4c����gШm����Ƈl�C��".}�r.���|��)�'�C�I	��`9�Ǘ*l��0�u��4��C�	N!Nxg���-Ґ����
��C�	�+LX��W��*:o� ��,
�V �C��%+�4����H��
�bȶ5t�B�� ^��"5�KByp��lF�U\�C䉅q�j�3�Π>�D�	b�C D��C�I�CN���'�QZ�*��mE&C�	K�,�j�2�хKЪYg�O����Y��գ��a����#�B.d��x��I�2P�Hg� �<�Ay���<<PC�3A�0����I�}�$�M�"�C��vLt@�b 5*�|y"	[;0?.��D���B�Z�&a�x��\�f!̜�70D����W�91�\�$��L;����.D��C�%Gx`���s-F*eG��s2�'D��;&J��H5(&�3'�Dhe;D�t���	/nK��GC�	 ���E9D� ��H�tz��� ,QGAd����9ғ�hO���a!�	��
)3�O1�PB�:L-Ľ��_�,-�[���NB�	(b��3��t����bC6B�B䉍pZ�U�
+�ʜ� k_�m�C䉈A��-���v<}���^�T��C�I>����h��E��������C�8a�%c���>��p�dH�1�B�I���!�B	8y{�����83<C�Ʉ���@���-9s(�B�@��B�I�Bh�p�6�ҽ{��e4�^�d2�B䉈E�D�X�cC�hy����._�s(�C��*L=1� �9t��\��AB
>�jC�?[��࣌�#W�\���-2	BC��h�V�;��Ʉ;͞��լݱ�C�9-��[b [
M��Q�Ϝ�!��B䉕OP�\	�e���=)d��0ԸB䉯t�µ�����R��Ȫ�L�:Gx�C�ɺQ�qB4,�9�4��fL�)A�C�	6:�h����I�^��a�SdC��
vM�2�)A�1RFQ�C�D�E�8C�)� b!x��"p�~ �@�_�K�p�B"Oz�`�/p����K�'�~� "O�hzQ�D�yn�\��'J1�Xv"O.Q��QRJ:օ�s'$� D"O^�`��^���t �D
xk"O��!�h��mCX�1f�V���4�*O��XÆ�.O2}�hΆ`����'c<|�&E�V<� C�c��);	�'VF��&.��)���6!�&]۰�b�'V&�#��b><]����ZBT�p�'��� ��Xm�1f��CA��q�'�@�� $��z\�1 �ޑ3e&y1�'�6�p@ҙK`ũ��Dv x��'a��cME���	z�ˀ�{�(�'+z@�$�/U2�c� �x��i��'�ĵ����+�8\�cE�m��:�'^B�%�4X�d�jr�8X��C�'W�(`̣@�hR�!ާTu �
�'�0�E����fN�G��)�'T�=��K�B�zh�#bY>9gR�I�'�^��W�E74������7?�X�{�'׈��	�|�c��j�岏�� �zĀ�E���Kl���gnC�O��ԇȓ�Y�AA�@Ú|����*;��-��AOvY���$k�u�3$M�|9��K�a#�Ӗk8��1JH�����lJt*"�¡X����*�	��p���i7�<D~r� �d� ���4�����h�4�y�	��<�|	��o*W꽸�(\��y2dZ�2����'NU'�BU�2���yB�C�pӪ�q��/���
��5�yR.^1v��ԋ����L�����y�Y.i0�0`F�]��pS H��y�	�q >�6�D�]`�0c��ŧ�O��=�O��q*s�< �,�b�m�h��'f}�3��D0�,PtO˕l]|H3�'�2�YG�ބ;>�h
$��i�����'|,A�R
J�q.$�"��/�>p��'�@�ԩ޶%����dW 90��'��aS��[��9=:*��
�'�*!"�
	>@N����oޚ/�N�[�'wv���fǮV���qK>$z>��'b�ڐ�
�T�9q����J�'�̒an���ȡ�gɚf� ��'��E3�+�3P���p�@�^m�!��'��%Z��#��t�׌W&�)�'��%��O:
����g�V���
�'Y�Aq��Y6�ca�UݖT	�''�}�y��L�:�Hh�j�"(�C�I�T8�r��^�#U��� խ#��C�	'VX`�%�=$�e@����B��>+�ٗ��;qbza��
WVfB�I�4h��#�Ǡh <���C'GB�(8y��ŬST���� ��o��C�	Bk����h��cc|�{e�,Q��C�	�!�paˆm3
$��Y�e
�G��C�Ɏ��5[�C��V=v� תD_�~C�I�R�b�3�܊�NYj7.D�X�dC�I;X�( �CH�;�MJ�f�
?�C��l�>�c��^��`�*�^�8O�B�ɤ���D�;{&����ܤ%��B��?4�2m��c�+�LA���E�8�RC䉖���{��3E��B&0 �B䉻O"<D������ U�j>�C�)� ���g-+>�T�Za�X�6���"OH�%-V�r��7�R�,���Ya"O�;���/x��H �MQ��e�"OlupW��a6�tg��%a*J���"O�8aV�#s������z��6"O�����I��RnY�Ì�Q�"O±�6�\F=��G�&��"O��qP͞�`�a��e��
����W"O�IWj�O�a��A��d�6U�v"O�q1 _�l%(\�rK����"O��r�
�;-�� ���G��[�"O���` ��F��m*����=0�';�ؒ�(8|�u�,�) �H�'�\�Qp�Z;m������n�MA�'�t%��M�U���d�͚|�RAI�'��R�(ݗ&�=�ԋ��p��I�'N�豤��/�Z��d��$\��P��'A�Ѩ�&"y�y1��՛A��@��'4(���
6��%b���f?d��
�'���cN�/y�<e��
]k���'��a���Rǀx2O��[�d|�'��-	T�5]���1��^-O�nL�'f���G[!wqz�{���8��h��'�X�$.ǝ�#ѯ�
�h���'�KF� i�3�Ɵ�x`���t�<��fįG4�H0�
ݱ "�ً�Mw�<)G�ځ2��34DRr�l�'u�<!�!Ɓk`�`�����U�]n�<1�G���`��@C�Gm�<i��H/i�XJӌ�.!u$)���o�<9&+�&u�����[+�j��j�<I�i��*�IPdLU
?��B�L�n�<�`NبtK�I�MD�����j�<9�a�b�����ٻ_�1[3��ȓ7�����:Xd]�ω'B"X�ȓ=8J�y&I(T���%Ӽi�@ �ȓyl�`[)9X�Ѱ����	�ȓ�hd; �P.xZ�M�u�nɇ�N(Ҩ�t@ZU�z�¨Z_쑇�-���̇+2��1s"�,d��ȓ?P�\rF
�nŮ �� %�t���N�d�7���V݀B
C;!e���y�*�R��Q�4��0#׋�m,:A��S=��"��9�<�d���"-�ȓ	��i���"+�,��@�ؙ�h��ȓvx|���%�� �E���ȓr�d<�����v���J_=f���ȓ"� �b �O�N% �)u�ZZ����v<��O���PzG��?MM�ą�r`�y�-@=:�b�SN�I�|ąȓ�֤!�IT�C�2�r��=:DE�ȓ^Y�hP��޿*�b�:�J :ʘ!��^�́��ʥ{�J���Ԟ4v�	��!iڕ9�Q+�(�����@��4��Rԭ��V�ڸ)30��[E�х�VΔ=��Bߩ?��"v�1�u"O8 �UM#;,5��JQ�<j�y�d"O�uc���e�.�*)�aeX	`"O,��Ƥ�;s4*�J�C�E_*x@�"O<��uFz�~���dW0k�"O )J"C��v�̏~S�YÇ"Oh�@�H��6�^'`��5�T"O!cmoÚ-��c�/f|��b"OtQyUjԔR�
���!��9Ѯȓ�"O� �8��RpN�9"��P�+^ʅ� "OVmkBGM�-�d�(�$Q'-M8*�"O�P0��4������*�0"O���6�\��q��{ `� �"OUCc�R��5�aUGT�|J!"O�.X�Lqm�!�T�Lਤ�n�<��JMD��B����O�ְp@�Si�<9&K�oF�	a��
����"��K�<�`.=��(XJ���cmƹ�C�0��y�������x#d�Ŧ@�C�	�xݦ<!%'$��x����I��B�=%��Ӕ%ԒAؤ`s�eϑk��B�IP��vc�,���A��M(��B��<u����2��r�����(��B�I0�bEP���y�D�Y�&��
�B�	)'HN=��T m�����ZC��;Q�x�Rec	Q��3��>�C�63G��3��O�J�� ���M d�B䉯 �87M�h�ޤ�Dm��>G�B�I�D5��c�H�7A��)F$L�zzpB�I�hbl Ȱ�Z�U 6ݰ2LݡW	jB��=!�^��3��3?t`!SD��9gՐB��5-gZpFbP�E�#���>!�$إj�X���S
$�����SX/!�D�1(�l��i#~&@�#��pv!�$F�>4E[q`	�r$��Ǉ@�zC!��mj�Q��	xf��I�'�6�!�d��l �A���W,���fR,�!�$��B�$��QfC�`H���@�=�!�$��6�JHe�P������ �!�R�I���YcBۀ-��5R`�8j!�dZ�lWT,2��V�[u4����;s_!�$�l�h��ɇ^����̲B!������hZ� ����� �4!�$�4zD�;6]�c��V"�<G!�$��S` �Ċ3x.He&�@!�dռ�%3�͆Yg^�	+Y�L!�$�4+�X�)�l�3t�"a��ρoh!�G�>����S ���Z�HPh!�DDPiP�y��V�L�
Lå瀵}F!�DÒ8j�fW�h.n�rs!�	!�
J龜�L_�c�h���*G/!�D�;8�a�B&',6�p$�wE!��"�tp�H"S{���F5�Py"'��}��bS� m,�X���"�y"�V@`8����.]���S���yR	�&l1AvkQ�%� C��+�y�W@� ��k��D`�핬�yb��:?�ІjJ� �N��y�C��a���(���DP`��U
��yRU.ppx�[$�#6+�!8u
�%�y�.�)� ��1hշ,���"��A��yr�FMtN陧'R'�vEB��'�y�H@]sL	X��{����ʣ�y�BBZ��̂�� Pi�b؝�y�HԾ?qxD�QN���U�P���y��ơ��@�E��}48��&V'�y�@
dQ�8b�ͨuT�1`sW�yr�.�ؘ��(L1"�D��[��y��q�šA9�.!`��S6�y��\>X�؛���=6n�P�[��yb�,S�8	+�ΕX�����y2�ܵe`�%@�E�"bs�)��Ʉ��y�ۢ_� �W���ڵ8���y
� �y"�Y!��1
�.�G�hܺ"OXTA�/�+ݰM���O�@�x��"O�4�R�B9FM���m�$$�"O����ԃ1$�)�r��	@"ONq��h�5�=@ÊQ�*��b�"O��;gO�) �@]�	�D"h퓥"O���4ʎ#	F^�rhZ.'>U8"O$M��dɍ'��D�*яuʪ���"Ol zm���"y����2�h�c�"O$�S�
_�Bz|\�g�؉fx��H"Ov x�bB�@7�THrCY����`4"O� P��.[A&S��6��4Z�"OT�
sɈ7^;�<y�Ɵ�(}~�7"O��K��p��f�=?�~��"Oxm[���*�*����(��9�%"O�$Zco���t�Cǖ)Wh�1�"OnAQ�h-p�^eXakʸ4V`q�"O�p�`�$�<���Q=2;r"OV���dG���m��"Q�	:V�zA"O�Б
AHq�a�ǚ�5$�s�"O�1�f��:��Q�&L uAH�0"O��@F�}y65��&K�[7R���"O�����d�`�e�.0��]��"O���`N$Q�~�r�DmPtS"Oh��-[vl��$��)�A"O$4Ф�N�3JB�0TB�'��9��"O����+vF��Y6c��QG�U�W"O�1�aX�~�D��^�襈AN �y��ݸW��y���$������*�y͖҄L�X#���J8�ei JD��y�o�"�)*腄E~8������y�`��:`�!�@	[�
I&ɂ�y�$Թ ��}i¬P�st�pu�y��P:�
�jF���^�	����yo&R@0��7c�-O a�����yªĘ?c�0c� �1��p;���y�J�;Z p�A��).�ad�އ�y�.��
p���6���3EJ?�y¡ܛj�@y�݌��aa�LѶ�y�b
o(�d�Y��M���y"Cʱ&V,�a�"á�V�k$(U��y���W ��i#�{���"g����y��A�"D��&)I4
�N�8���yR�<�|���ҝ~.�ppC���yR�d�v�xq+�pܤ���,̰�y/�n&j,R@�T���Y0kZ��y"-n��`B���E�7j���yR�ޜ
�8�*��JɁ�� �yR�G�B>��; dK�=�Hͩ�ͻ�yₚ�2�*���~�$E
�@C:�y��!8ZRprWd��D�:h����y���'��J�aBɜdK�MX��ybDX.J�TTKrH�'<���0a�Z��y�o,�dTɡ"H�0>�
�Ý	�y��Y�"UAKю0�X�q���yb̙�ug���O&*09z&�� �y҉�.o�j��U�%;���0�L�y�́8��c��6uf졉� U,�y�%�W8�po\�YkH����!�y�A�f��� !��A�=�Q��;�yRdN��[5'�|�6-9�Ȑ�yB�ޭw�|��AZ9\[<��e(�y�ƀ4�^t������ �A�'�yR�^���Ar �_�>�ԉ�,��y
� �0z&��DY���.g�T �"O@�(Y5�D�h��!]�Ţ�"O2!qEH�=70�\����<M2H� "O��a��M;�xi�)<$Q$"OTX���"�$���
�i$L��"O*�h�JT'(�����O��%�b"O������&YQtL{�&P���0D"Ot�ْ!\Ԡ���=p����"O:x�şxޜ��qd-'�͙u"OP��Ɖ�/�x����g���D"O�����I�8�H1��$��"O�XC�� ���(4�F�ܴ��"O*)�2�� ��4r�Fl�t�"O4c#��[���1�d�����"O�x��FZ=hZ���S�rz��P�"O�h1���2�����5o�+"O��R�jX6(	jiie��~fZ���"O�Q���3=����1����"O��)aES�dp�����6x�G"O>���6W7�@�S�M;@|]�c"O��H#,X,M���P�E7htC�"O)2��M�+�&���P./gX�E"Ozp��č�
����׫�,2Yl�1�"O���w�ŧLM�ܫW�Jv��F"O�<r�-�+Z�Ѻ�1=��"O2��?�5b�ľPt��"O�H�EM�4��铴N��l� kS"O*\�G��<z����n�t�b,"O\��tm֯&�4��&�A1Z�0�33"Ob�c0@8b�(X;���$}��� c"OJCGD-�1Iw,�6�@��"O�YГK7g��``,$�|q"O��ԧ+�P{m��0�pHG"O�(�固b:�х�ҐfV鑒"O����yTMh5���-b�,;�"O�� �Ʈ�`E#��Q^GDxYU"O�S+� ~��"��#+*�)�"O�8���� F.��,����2E"O^8����1_��+�2"��p"OB��a�"8�հ�J�(�T��d"O�	J�8�F�pь�9gO����"O���3��*4f�4�6jg��P�"O�4`0� �E���K Wlp��"O�l�QbʎZx.%�G�.*c8Yg"O�-��jM�cL�,8�n�OR�;�"O�x`s�C�nɢR�B�8=e1�"Oҩ�7N�:�6�^�X��,�E"O�����`Њ��kU�?����f"O�q��[�?�T
�+��{��!"O�d	� �X����ꉙ	?v�ȧ"O�̃��[�@�7IH�1�u��"O�@x2�άUw�1YT��-H�����"O*0��e�w�dI�/�l�a�"O��hġI�]��8[�@��d�hd�'"O~�`Aa�?P*��p� ҏ]��$�"O����@}vr}C /éN���PG"O��rH6,HD��p�1"Oڼ"4�E,E�n\�V́�^�=�"Oν��A�����qa�/hl��Y@"O�M���M5H8�!�h���Js"O`�bE�J=]���`����eb�"O\@iĄǰR��Y�SB����"O�-A��8Ty�@`�nSH�4�K�"O �Rh�p�^̂�l �~�T}��"O� �@�@
�-<8�� � �Zn>y�`"O�ț���N���m
,lOu+Q"ONj���N%rPj��K��@�Q�"O���b�o
d���L�$����E"O�蓀�G+�z�+�1ͪ��0"On]��#�t��k�-�+R���"O<��sJ�N#��A��\ �"O��n*Z]R��!�0I�nH "OBt�2h�2͊�I����B�~�D"O�(�2�C;h0��'��0P~�z2"O��jG�P�MSL������Z�"O�����l�@�BQ��)�z��G"O$���!�$Rz�0%(�X%�D"O�A
g�¿fۜy#M��%��1!�"Oxp�Ү�I=Z��L��z���"O���)9<���EڢP���X"O(�*�F�x�:�j��	8M�����"O��h��U=�=�R#G"'�0�k$"O��`�L"
Kr�b��܌��G"Oĭ0�B�<�h��ć� 6��	�"O�- -�����9�� ��r�<�b�Y��4@�&�Hv���t��k�<A���)cm�Q�L�&�܈����k�<�f�E \��tf\�U�NA��Țh�<I�n��p3�8e��y��Kg�<�a"�6��`C�=��Lav�]_�<��E�\p|�G�9��D��nZ�<ْ�?�ձu��2T�6�)lY�<�cbX� -V[')M9Z9��oq�<�To׺7�pe
����t6�x� m�<I���(J.��wK_�T�j5���}�<a�j���<`V.D�p�\�5�F@�<��),#.�H����.v��� Bz�<)���LC�l(>K$8���v�<9�×�Q��@��$�Gؘ YIu�<�C�4l��b�>0^t�G�s�<I�!	�2x�T9��������s�<��E�1o����.�R����6��q�<!@nX�
r|Iq��qÒ58p�Rp�<Q��1l�dPGڭӤ���Oi�<�pț�h�7hM<Y��%�f�W�yBZ"+�D�	�� �șq�d���y�'I66`T��C��t��⢏K��y�!B�AJ�1;r��mA��y�� �y�Қd�P�R�O+�����yR`�),}L )��	4������yRM�+���xW+���2���y�-�?2A|��I�;�-��n��y�F٨x�¤��	��d"G4�y�Ü- ȩ��	$�p"!�*�yReE9���)5�[�=0 l��yr-5{������h 1gÝ�ybo�j��i��*Q�v���ѢK.�y�@�6B"8���K�l�� ��μ�y¢@�F�x|z��!aZe�U�M��y��{���	�B6V�HBu�_��y��WT�PeYFD��=�j��Ej�5�y���[7 A���B�$L�	H	��y���-��!��$�����yrL@#�F쓰b]̔s�L���yR������*R10���Y ^�y��ˋ;|T1�H�?a�1D��ybߐP�@�#��M�����1�y�����`C�B�m�������y
� � ��B4�޵��,�9n�X�z�"OىB��4lA�I �:d���p�"O�E�֠�%k*hR��Q-G��Ph�"O�H�&�',��v��#���"Ox��錂4F��g��B$�5�&"O�yS�!t�$�t�R�m4Bt"O贂0��=pd�@�L�Y�|�4"OZ�& &0#�$8D��UH��"O.%x�m^1�T�����	A
�
2"O��q��i"�D����l>\�"OT�Z7p��M0N��G�I �"O��X�+d�p�����2a3�"O|���vr�yj2��6-ܴ� �"O�@��*_�n����*1<��"OF���f�{����iX �DB"Oj����PG�t�M����p�"O�y�s.��"�X���扷k�*��"O�����ܞb� z�K��UwQ��"OJ���ǐ�& D��#J�	Gb����"O�9a웿=p�јc)��j�N��R"OP��nڍ*���pC��w��x�"Oʭ����	$$���pG�Mν��"OZM�$Y3;j�Y+օ����3G"O@�{�`J�a�����ɕT
VК"Om +B?Bpع{TCF����"Oh������2�Z�:��J(=�&I#�"O�YP�N��t$J�!Ǉ�-  T�"O�d���=��y��FY�X|j�"O|e��aT�\�ؼ�!OE�2��"O(i�c��N�B���:�Ie"ONl���ÿ!j�0b��R�_��P"�"O�Ū��8~��8��"ǂE� � "O��Qu�_"\�����z�pu��"O``RhC�I
>���n�BE"O*ɺ o��(�D�^�2"O�tä�Is��qun{̲U�%"OM�E�U�u���7�R�c��4`G"O��r�]�n��r��T�h� �"Oԭ0֣̱_��cr��|$:��W"O@u0�k������䔀z��"O���Շ�9.�=AgN�=����P"OTHbF�Q�	Un(��*Q��"OL�Q�	�F� �y��P�9'
��"O�4��E�~ �uW�V��x�t"Ot]���'�@�a���0�"Ou�a�_2]���ː|��"O���׀�5] ���Fɋ���xI'"O���Tl��t��Q���:�L��r"ONQ21D�L���Q�喔���"O�a�sh�*>�و��u�B1�3"ONa�bJ�/� �3��^�Ĝ��"O�X�$�_A�6`��]6>�p�z4"O�(�"�'A��� ձ$jp��"O~`CWC&"d;Q
�"���u"O�p�����p�bܠz2�A�"ON%S1L
$,�t���J�&v��W"O���f�1�� gc�(4ψt2F"O��X4Oπ���`�"�W�l�[�"O��:���(��t9#�~�l���"O�hX���--�Aʇ�1PJ%��"O��ّ�:HMJ��o��9�DcQ"O�p��ĉ���Dwg�>32T�A6"O.娗�W=xD쥡2���%O̱"O�s/=&�<���+gK�Eڒ"O� �Ei��@(5'N�S��=m/&$�b"O�)����
,v�AbV̄�Xx܈@"O|�`�E�)�@�Q���Dhd�ۤ"OnH�5D�m��ip3��nW^�*d"O����	�%�������l`!�	�'��xbwa�Q
�T�bi�5<s��#	�'�D%����d��5AR�P4$�M@�'*���@���pb���'�~ �'M�+�,E2�H	iI
31�0��'�z�)�+�7���bw��-B`@P�'$r��t`���	�FU3�B�'�`�����=<J�*V.,���'����|�Τ�� 34 "�'>�pPTYE�"=C6��\Ӷ���'޴ 'c
Z�(ǃ�+NM���'�4E�l�;?��
�:���@�'o<˶K�mb����F� �����'K��� cB�0��в[&�
�'��]��D�<��%���+C�]��'���R���D����� xPq�'� �a�.��8M�s�f~1��'��-qR�յ5K �i`�Z%7���
�'�쌊m΂!װ�HP��u����' (`���"txwAya�dX�'��Ųa��� ���E�z^��b
�'b���(	����8׏Юz� A�'K�u�g�K��3/�=n���j�'�ld�6���gP��xR��d�؄{
�'�D@���)*>�y��U�c_P���'VMz�bYը��K�Q�rl+�'����U�G�q���M�Dqz	�'锰K��2�1�I]�ڐ3	�'��@�,��B��#��
C8�	�'����3�P�A<�J��Q_f���'�z�bV"M6Y�mIeK�3w
5��'�@H����?�H�Ӥ�c(��r�'���f�ߌra���"h�+S݀ ��'>�Y
�+���Ҽ��`�W�xQ��':����:0Y�F���P� �'�F@��mF|Ic.|)6�@�'N �j��P�L�\��(����e�
�'46(jCK3)ԑ���$d(�)�	�'������w,0���S�U�=x�'��u����^��5�$d�N���0�'�1Zu��9Y��]�t�u*.$�'��pB���	}#h(�E!�w����'j��d+TbŰ�I�4"i�݋�'$�!�U�T
�hV��p0^ ��'�6u���Ѯp�T���؈k�s�'Ғi��"�bW��/!��vC�n�<��DL�O�5�C/�[@q����n�<	d��u{ �f��@T�W�H�!��M0cs���Q�Q"D|Q��Ž�!�D�$l�r�@����|_�ݘa#�X�!�ĉ_^�8R���TJ.�rq�I�K2!�d_�g�&� �G5Ld�s a��!�D��Ld��0��fT��5�G�"@!�$M��V�(=��`��fƲFl���l���瘆��mK�o�<G�	��|�H#c�$�t\�pF_�nø��ȓp>	�e��l�Es�B�h���ȓm(h��R�8��c�S�\m�ȓ9�p��A��%E�X��,�.x��_����q>F��!���Y� ���S�? �M����Xw0��r*��5��s�"O��*�ȅ�!��U�3ߞ$�w"OzR�.�-<�^�#HȈi�!�s"O����
�;#ځ0��7h��!"O.}��C�}8l8�����C�ؘ�"O�y��R�k�4
�@�-�Z1��"O��!e�ā7"`#������%��"O�yC瑷4B4	���z��W"O^�Q3�B�!�R�A�f��Z��)��"O�Ġ�N�:�z��* Np�c"O��zĀ�0�0S��|�F�s�"O@�U�B�j��i��������"O^��t��?^�A�Ac�2\60Z�"O� ��CX� $ ��g��#��$h�"O�} ��=���"��ǧ9��B"O�4P�*ܜ�Dy� �Y���I�"O 5��ڔ0��es�$��x����"O��� ��������71���"O,{6�ґ|ѐM����%�5�*O��d��E�h��U*��
�'���E��x2C`'a�X��'�fPX&��7����
�v�D��'2�%���U_A�UZr��<^����'�h(�B�D�a@���	6S�tH�'ּ��fHޜ$�!oR�R\.�`�'ن$�3�&ax�JQNȅ��c
�'_t��t/� ��)�@��P�4t��'mn�84O�kO��h��@�VT:��
�'<`l�"���W�PH(�̓G(� H�'D>� ��˖i��y˱��B��M��'�Ds뒊r��[�"��>v���'$��p&-҃OS�E���G��I��'�aB��
H�`g�&Jm҈��'�,���%*V���]�$���'^$�â&@�?�D@R�ٶ+��'�P��T#�@ ǎ�,}���'��ܘj6n�X0ʶd�(w~���'ܲ=�Â�2���
Do)f���'��HVeȇ52p3*��1L���'gjI�T`Ó8�6�1�%�G��r	�'.l-i ���_��!�G�Ǡ�&��'w����\�d�ȼb�M��6\2�'0|�'� ���(���,��A��'��=(���	'�v��[��@9
�'����A��5`P�bN��y�ꇣOYXt(b�9-&�Ue�v�<���ۖ!�Vl����c	�͊�&�f�<���X�A���a@�
oT�:2��c�<����2=�AI7.�B��ݓ�_E�<i��61��@�0�t�g�h�<!`�-�N���/�2����g�<9 ��&q���g��)i�p��Qm�<ᒉ�(PT���\��)#��Fi�<��ጦBy�`)��hZ���d�<��%�h��A�W#���"���^�<�)-$9���'�R� 㰅�bEAP�<1 �
X��#Cl�iw� ��f�K�<��J�:嚔J炈 F��q��R\�<Y�%ƺ	-�e[���@�����%�}�<���>��ʳBE�^�hy�T�Gw�<�c'=@�!pi�ADĵ9V�K�<����'J�\,qBΗ?� Y	�fU�<FڤB󶰺uD�(OƶUI�Fw�<ɄkS�-�h�!��; �����~�<� �҈���p�C-�3p�pP"OAa���" �]3gA�o^8��"OF�rk\�-$ްCvB��v�H,�G"O��%a��q@������y@`�# "O�л1NI!@����"`#Z","O�,�!��E�všF�3r�Ч"O��C�i���ġ[�#F's��e"O�XQ�B,vn)e��o���e"O�@2�ՀL�|=���ϡZ�c0"Oq�$��;�J�{	ׇ���"O�h)��Dg�fȖ#Y��X� "O")��T)�uG	뺵ڃ"O^2�\���G�R�v����6"OP��S�܄c��&�&o���AC"O�	�vk^�R����U��g`e0�"Oة��0g��9y���WϦ�#$"O��ʆn��\SD@\166�BSH�<Yr���հ .
�H�A��nRy�<р��E�d}@� ]�b>duIt��q�<Ŏ��a�^�ҋ��OOr�C6�k�<`���
$$W�E��ɐd�B�<YS�D�9V�d���ÝO�2<j��=D���W*�KHA��Lc�@��<D�����v������H~ԅl>D��rN�1�3-��&����K�3�yb�<l@��!��r�	��ߝ�y�W����Zu�P��+�;�yR뉅Dpd���ʿd_~8����9�y�+ �ynm	��?d"=w���y���7|��]1C U�Y�x�`fCB�yR��o�|u�DjU�Iji{��Ψ�yR��F�"�(q�I@j�Q6��+�y"�Ծ�P쁲��/=�t� ���y�Āts���7јFT���>�y2-݌V]�����B�M��3�j
��yR�O0�麐�H��X�X��y���s:�Թ�D\���آ���y"�Y=ib�5��[{���{�A���yb�A&���dE�n1��bGo+�y�CW�Pl*���*b�f��cЩ�y�Q67BH�FbT[gh4Ӡ��y��u��"�.R���0D'�y�gO�PB���d��H`�����Y��y2�U*�ذ�QnV���M��y�e�`U������b#A��y�+F��AJ�d0���)�e��yrO�>T��
�.K�i*H���A��y�c��&8�ۇ)�gTZ�֊���ybn�#7q�=P�0�ʨ�	G!�y�`C44�0�&�O�"i��Y����y��M����W�1��,���J��y"$M�r��/uqX� `�*����0��e��J�%a��w�� ��	^�� ��P�P���"ԒM�z܇�KD|Yj7oR$1������Z¼!��=� ����KcP�#e%܊l�T��ȓ-�0���h=;���c6�
��ȓZ�Z�Y��1O��yT�K��e�ȓvE�U��KE�k>�Yi5�-qp��*a��	p��/v:ِ��(o��	��Vʚ��a�J��x,��	B�1�لȓ1����#��-;�
P�0͛�TD�نȓ� r!�0O�J�Ûr-����.��9� �ވ=���j��*͆�S�? h�9uf�� ������F�Q��"O^Es��i��ѻbU�d.�ˢ"O��5�ޑV�l�h�'T-R�\Q�"O�Qt��!q%,dI��w�4I"OVD	�f"i��6�º(��i�"O���FX6���C�5H���"O�P�f��3M��X��ׅI2�r"O���1nkR�����)u.����"O�;`(4&����qOU�&��\��"O��������y�  �ixVl��"OX��B�fZ�I��-Jv�!I@"O��!'	�,w`,�Ӎ]/'j�lq2"OxX 	�.; ��ծ	�wa���"O(�`��(<U\I�-��S,�"O4�	4OV�<���陆5Į�Y�"O$PSeBÛT����9l���F��P�<9�ď({�hcT����@��v�<ɓ�Ƣ,|a���#|�ĨP���s�<�gF�<��u���$8����r�<I�!�|_�e
6�
� �lrҧ�p�<I!��AL(-ۓ#��G��c�n�<QՅ"*���7�IS�&�f�<!���*��A��K\���PĘb�<���
0n���vH��L�Kv�^�<I��G��d�9�F�F�j�+��[�<iW�5��2��'�x ����X�<1 ��Y����B�S6C�4��7�W�<��űz�D�K��@-j�"��d�RV�<�1�B�9�|�aDC�>G��r���I�<���e池�@\	3,6풵�]H�<��V�R������- �:���e}�<��'�=;��*��L �؉�H_d�<��HH�+�vu�,[~Y�Zc�<�� R�%Qs,�~�:yâ��H�<b���$j(ҳp8�h��_G�<�A�@�V��V�ЧZ��8�e�Y�<�Ù4h�L�����3�v%�3�T�<��
0v� �fýAmF ����y�<q��5
��Y��O�W&�:@Hq�<y5ᜲ{���%Í�4��)3�Ru�<q�g�E�<�!K
�t �@�o�<ٰ�h���5I�>�&'�l�<q���68	t�"�����5�q�<��mU\�r���B&
�8�9���d�<���P�~�J�y�J$y��SL�a�<yM�0�괫�3�Y4C�D�<Q �=Y���j���[^!��{�<�pD�xO�)A�V�#���T��x�<��%H�{qX���@n�F$Ғ��l�<�R�S1K�4񃵀Y�h:����f�n�<qVL���8eP��^B��IW�s�<���*6�@��3CЕ|KX}2��u�<Y��C�h��i+P�K8x^Q�欖I�<��d�7eu��@A��1B�M���\�<Y���;(X-J���H�nLQ�Kn�<y �׸�~}2����&�V�c��h�<����m�(1��)=����d�b�<�F�ޚ���AG��$Ɔ�x#@@G�<�O�2hؔ`Ѣ 8����YK�<�CI�R�� c��2Qy8Ո�^\�<1���'_��)��NÆ	�\ �JU�<1Ǧ�=F��R�T!`@� �x�<�&N��lxq �>N�F(���w�<q���czy���](�أSi�s�<� AT�F
�*��2�� ,���S"O��bcA,�i�5&�A�"�j�"O��`DiW%Y�����'�<�`�"O6�˥P�On8���Ў2� ��""Oҕ����^�`!�2"L4B�p੕"O(%��ӿY���J�%���"O`�S����/����1�
��y��75F��pƄM��jɯ�y��M�+r��/J��L(#��y���)I���A�!
�  xg�F��yRa�.~3޸�I� �6�����y'H�@�X̨P���J�@l��#��y*ܩr�<ؑ #?��L�PNʄ�y��jlT�	+�:�5sS+���yb��>�n�QRm%�X�!�>�yR
W�t,�i�hg^��&[��y��V�*0���oپb��i0 �*�yb��%i�8�%.��xh����y�'�
$�(�
#���",�����T�y����ԑBa%"��A�W�
��ybd�	��e��J5.�Vq�V��y���* �0�*�'���b��=�y�N/8\\�`ȁ�l��&�ʹ�yr�5#�(Pk%�"D�@���y��w�H��G,F�"�2Ż�M:�y�K�݅I'�p�I�Hӡp�y	�'ƪ�8�ɓlk�-�Dȃg]!;�'� ���ڵ&� I!#�L*H�0�	�'1�A��*B���KV&<��	�'����Um�}�&��!/��u
�'�re�E=��tS���t�`
�'�D�3w$��:���R@����'Bb��JJ,c^�mh�N/�h3�'�|� ��֞T��SFΒ'?��!��'��gMѠ\Sz�����5���#�'��;�� u	�HT�&�����'�\��4(kz� ���"^�j�'s�%;��ɪu{�	�@k�&�%��'�-(�E�������!_5^<��'C��jT9DB�c�
�w���	�'�ڕ�ԅ	Fv���+ޟt~*h1	�'Ԇa�"N������&<Y����'���3���0څ0� j�$h�'�@MCVe��p�@�� ^�4iR
�'�|Q ��q���]�e�	�'
���c��%ZYQ�b�U�v$�'�xy[�	90������ޅ_��$;�'p,q)4l�2w�6TpPK�g۾1�'{��sC�z���35#V�]ʼ�	�'��ҮH�8�j����S _��0	�'����,6���w)�\X-��'�J�[ǈC=2t�i;!���H�Qh�'HI�L gz�K1������'��'�IND���3JAR�'����3�آu�>MX�CX�����'Ū(2���tņ r2`�3jƒ0��'K��ڐh�$��K�.�"%x
�'��ݺ�
*D�ax�.�<#, $�	�'2D=�#�S�����2�D��'�Ћ�UKr]X�%8�Y�	�'8~8�u.Z�L�:s+�)�b���'�����U�U玥afȌ"� )�'�v<�ƅ��0�TlT�d,�D�
�'D�ԧ��a��ʤ�	%�f�3
��� �< �b W���s�E$��"OެpAi�c��1��<w7Ę �"O��Di��&D4����.~(lDq�"O�#�ċ� &�qBam!Z���"OЅ�@��"���`��
���C"O��3&E�,3��%�WG22�{"OJ���8A�~���_j)��"O���JݠZY��q���V(HuH�"Op0�I]���t8�i J$�`"O����ju4p���#���"O�U3V�5C��)���,
ș�W"O�!Җ�Ϙ<>>a�� ң(x4`2"O<)ؗ�����Ć]	��*F"O�Ӂ�!{��	@��:��@�	�'*p���ȿ�v)���G~Q�
�'1+�[paZ���z�\x�m#D�`��)K�`�1�G�Q0}G�\a'7D��2D$Hr��9���
���eC��y�07_�,�*�6����%�'�y��՟+��3r��.@$iq��D�y§֖j䄅�  �x����y$ٚ- ��15KL��Y�6̜�y"ő+C�H§F�,�F��=�yR�2��|bR�_0?f��Pm���yb �0|���?���Q`R%�yҁ�$;�
 �Y:�!
�I׃�y����Ƶ�r�_$5Oz��@��y ��(=8ǘR(ڇ����yR$�,��20j���F�M,�yRlߗw��(�I|	�Q�U��'�y�k�)������{�����η�y�c�����eD�y��--	�����U0�1��R;��3��?Npp��ȓ�����k;	lI�C��L9��U�P���nN�|��$�����b^���ȓ-�,���
u�V�>Oļ�ȓU}̭є+�j����+5eV���|����@>�P`���3c,H��U� e�0 Ǎ15��o�Gf���ȓQ�U�"���x��Q�ߊWS�d�ȓ$�,��!)�J�����m^�5���4q�R�.:rm�d�		oD�ȓ��5�����!�����[�#tЅ�,
�L�'mN(e��X4�TPa�݅ȓ_��Ā�ۍ4�D�	s�[� ͅȓq����ئZެm��܀k�0�ȓl����ï��) C��Y.,�ȓ8tl����	P�=�t皌>��Y���$I�F=n�����bM)��;0�(�A̖��>,�A�15n,��Wژ�/�v�x��&�-eέ�ȓr,��"3�y$ A���O&=�X�����́����1)�M���	p�`�ȓ7�(�V8���>�"\�ȓ/^�����/-�6�h��ȼ�,P��]�p���R�-7hh(��<?�n�<Q�FN���m:��I)pІx�S�x�<���4�s"�4�|��&E^�Hh�C�	�%�F����1|r��&�ܜ��C�I�{����.B.Ifo�;9�C�I1VV�����Ҙt����wɬC�	�V��d	<������B�?��C�I�,�nl��.ۛ3��5�4b�;x��B�I����A(�?#�!`�b�r?�B�)� �	��I�.#7�%��^��uXu"O�YPA],;!���؈4�~�s�"OL��AӀ7`��
 '��J�P��G"O�0���Y+d���m�(Hр���"O�)A� [��r�,^Uݾ�!"O�uR�U�a�
������a"O����+�v�d�V�\����%"O� � O1��ʃL�bBU�1"O`����=Z8Z�۴�Q�u񼱙&"OB cK�n�`�(D�2K�25�"O.�Crb�����Ba�-o��tS�"O���K���rP��\�bAf�Z�"O�M83I�&`y��ܞ$,����"O�	X K�<L1jBn�]&��"Ol=�Aᚊ,�F���mB�ZX��"O.e�H3 .�q�"�,u
�"O&��tt�̠uN��\Lr�����y�m	u���`O��j��%�AbE��y�g��OQ�����P�Zf@�Z� ��yR�/� )S׍�!IQ�%yU��?�y�e�/-J.���&�F��X���ޖ�yFY4��1!ϊD�#��y�g�j��	�$ ΁e�j�xF�)�y��W;1ld2d�Z�^h�u&Ŧ�y"�[�LTp�!�*VԪ�R��&�yB�T��
3Q���KUh�03�xJ�'F�Θ�i,���1"�#D�l��'���j�흕e>@�h&��#�N���'Ҏm�l�`�����(�Z�a�'�H 0��?���㒇T��u��'|���%�V4E��8���R�pX�'ؔ�+p-^9g�)��Μ�]��,R�'	J�I �R����S�YY����'��|[��%���˒�R�LF���'�@�(P#!`h��g�K""9*�'�����&	e��#����p���Y�'�4�l�Hn�����YyҸ��i,4iU*�?�� YF�ϰ�ޭ��!�8|�S��| �XJ̳{�j���b����3QjZ
*׆);z�p�ȓ"4��4!��|��}z���$;�n��ȓU8Hx�6
�+H:�9ʲˉ��^d�ȓe��сU���
����*B�`�ȓ@�&Yx��(I_�1�#ϣx.�(���`�R�U;�*|�ת��o�z���~:��dC�aɴ�4��d�2`��q�(r����JP���ԌD��tn�%�!��&!  �Oϯz�~�ȓ\�~q���u@2l���(3Dɇ�v	��V�ӌ2mR2�(ݚ�� ��I�Q��6Z�z�1㓖ss衅ȓS�HaCB.T,�N�١g[j�����'9��s�['%�!!�՝(U���ȓ�8�C2�	�m�(��0����ȓ.4|��ޗk�� Z��0�a��Db��a�M	������C�;���ȓ|R̠S�5 ����_�T���%xL��	�.ά�[��;Y��E��m�|�r]�*�����4]�؄ȓL�S� ǏK4 P��ظv��Ąȓ��<4�W�Y�n��3K�$6�l��5��`�Q'>r�k�ڍ@c���ȓ�@sR��Y��}���
����ȓf���Ȓ`�j���4.��i��y��S�? �8�V�P�(��EX��E"O��w�Q-z�d�4��7��@"O�Ls� ��JW*�מ�@�"O����1Ҭ�Y�	�1�HiYP"O�=(R_�Z)B�9�  8�"O4d�@\HL�#&64��� "O�I�"F )���"&��!T,B��"O���CAʟX쎵��Z��~�[�"Oܝ�3 �kYnP"S��g�����"O�����jDM�,K� �R	x�"O�e�ܰ� ��N�x��"Op8�5L�=\����w ď0�H��"O�(R`��^�M�=d��0K�����I�(h����'C�|�v^6*`�B�I�v���,6:P��ɥL�2
�B�ɻ��\��B71�J%��c[3u��B�32l ���>b���b�M���'�ў�?a��N��x{�0�E�P�!�Έ�;D�0qsN�yd��BC��3�Z�p�bc��=E���&��,@ Z(։�a��!��C�	ɦ�PӨ8h�\LҬ?��Q��;D���
�G�m�g���z�j��8lOh��qd@ǜ6��h� ��LH��5D� �U�[%�^�(0nW�Q.����4?�
�{�N����I&��t	�8`
�t��@}B)[tI H������hڴ%�ȓW�28@�*m�-��B�p�r���Ϯ$b��Sd"<�X��]2d�왆�D)H��_# ��8@l��^�z\FzB�~��B؍o��3�!Ło"�-�j�m�<����h��'k�kdZ�F&Q�<��"�������; ��P�<�`�^��B�b�phS��ZP�<��!�S�����t�@P�GEҟnZn���O�x��'St�WIS�� e3�M�[	Vq�O6����(_Ŵ���VK3� �RK9P���4�O�S7�ܻG�9�b���Q�"Or{�c�#e�&��o��x��}"C��!lO�ʲφ�TJ���д]ɴ�Ya�>�����(v鮕س!I�dBSk�9�	Q��H�,�����S6��ƙ�O�A�"OLM�!	 Z۲���EeG�%��"O�h׏�>yrL�����K2`P���Ij���IO�J�f��I�0
�тHj��xr�	�p�1��eU%���,�&C䉗3���� ˧I8(��c��<�H#<q���?)����!*��т��N�r� �wM4D���̗�v�~��a@{V��Ƈ�O�7-8�S�d�$��T�^i��5`'�1v!򤒅V���G��<6���O���v����՛����h)��C�ˤB(�3"O�DF�٢�`y������4��'�'p�)��xBiW�7���(���T��4���x��'����b͆�����2]�	�(:D��X����5ĺi� �.=��[D�9�	w��r�'>i:��	]=��A�b�03:�m��'
��2�%�!��A�.>\)��ēI<k���WW���L9,��Ey��!��+�<��-^��"���%G�B�
&h��Ε����f��^U����Y=��DeӦ	j#F�~颔Yb���PxI�A"O�X�!�E���{��%
pj��'��'u�̛3	�i���H3�B�����O������Qr\�2���y� a�b�R.!�� 6�qAĕn�p#1
ۂnMnc"O����-?<lP�ToX�4xb%"O.��6d�1M�2�H��0�b"O���4��b�� F���"O�L�@��yP�#C��,_��u3%"OR�!/�%O}T�����p�P"Op�� �ܕpȬ���V����"O`�+V H�f1LҲIXG�n1�B"OX�C�I��9hnП+�>H0P��F{��	ѿH�0-
SE�Nx:�2�K��J�!�$�R�h��� M�e��4X�H*k�!��#
����.�΁��j��!���m�T�2�"�"g{�$�����M�!�Ĉ�(,Ѕ��M�h���ƌQN!�V	<�PЕ�O�I}l�����g��y��I��ѻ�DS m� *�3:C��
[��qA�P�@�.f�fC�I�fs���Ï�c�Dy�N�A4C��!gB� ��6/~��2C�� (�&���	/`��h��ȟ#���$ �e�bC�%-� @��?M����s#��VHB��,|�,�� �܅<XTC�ᇛOp@B�	�)#���ȉ,��uSCe۟dv8B�#5:&�he�
?ҹI��רq0B�ɸ)�aJw�A�'���kpHVu.B��!P���%	�P�	0�l%-B��!jKj�cqǃ99Ŋ�wi�	����e��0��%qb�M��������fF1D��ӣg��d+n-��/	��`R(1D���2a�ߢ�
&��7-��dRgD-�D<�O���-�6}��ż@,���"O�}cs.�9�Ȝ �MF�MTL��"O���dбMM<��D����+��>�I>!�%(��?�)c�A�?���x��L���x5"D�lp&�ǚvE��ze���z���b-=��ȟJ���L�iP��3C��u 8a�""O؛Ąs�Lq9�a� 2�t�w"Oz�����TH�hj K��0.:�z��>�נ;�S�==�6�ʬyв���N>C��a!��.D��s+��M�� �
�0�Q*6��O���S���.Ay�AC�'V�{(>0����Q!���O�� �lй*琁;��Dm�d4b�xU��E{��� p�♯6�(��@�[�D}���'2�'�:�����#��A���>b.����O��Ez��iF-�t�b/��xbD��
�*�'�ўb?i�� sa�)V�ܗ>o�a���<!�B�6���c�63 HD�K�0��B8� �>q�o�`yF�Ȁ�ê%έ	���w��$�LZ�[���m� �+���el%D���0C��Z,	��# ���e�"�		����6��DoD�{NXIQ�-R.����Oz�=E��GE�  �x ��.�v�� C<��=�b�|bCG7-.9��@Be������~��)�'QΊh�
��7CTI���[==�8a%������� ���&,_6������P/d͆�>�,�3F6Nib��5b?:aF|2��-d��L�e���FlBT-W�+C�	5K��H���^�,d����]�6�	����,MAOQpp�P�R +�Nŀ�"OJ��JI<2(�H�3!�yn�Q�v"O̹��F�b�:*B/�q]�B�'���+9��y`�̞	V���"o1�!��:O�fġ���7;�~��	4�!�$Ӱ;�c3.�y�2��UG�z�Q���'4�>�  �QD����a�Ɋ6 t�� �d)lO�+�,͔r!l�q���i�Б� O(�d�g�ʸ�ub�/���b`kԶ\"!�D	�JN��R�)%��ԉG	T4I	1O���$�*^����r�Q�5	J@C�N�6U
!�$߁R-��P"
�*�)C��!���Vc�kB�O�w�l8j��6�!�dӊ|z���k�2�6����!�D]/?o�������<q{@C�q�!��Lje�=z��Fu`�*��ȸF�!�D�*$r"Yg�]�i��$�T��o�!�
�a����X�iB��!�Dɝ?�8�bDm�	�@:c�6W�!��>c+8�s�ʎ�G����� &j�!�β%��� L��i&* �!�$�Є�q(��5̢%Ѐ�Ջ�!�DP/o�I�+��z��FΖ�f�!�dD�F�Sm�,2��� %LQKm!�DF�K^���/�;4����!l�N8!�Q+�  ��'��2z�E�3�6),!�(yVM{��[� �\m��i�H;!�d��'�� :#$�3=hJ@��
	� �!���jL����U�J��l��z�!��?F��3�σu�B�'�8&�!�T(U� ��qB�3�V��4�P�a�!�ۂ���SѷX�h�@��v�!�$��M�)�k�9��x���G�/w!�$	�@L��`,���t�J�H!�DA�ր@Z�X0]ܢ�rt��'hj!���`",p�Qe��BM�&a!��_)Nd��Rr��1a�8��,b!��A�z���J�]`�#��� hR!�$P
�E(b$C�N]z�Y�M�\&!�D�6�v9R�	
�8@�9�T)ϓ"!�D�i."�8�^�#I��'��'?�!�D��3G��� nï$X��u �x�!��6�L]���+�	[�+�!�dK ��hRk�7U��,4��(3!�dC<nc
I�rh�(n!n�$ T,Ʉ�+�Tiʱ��52l�xH�S� ���G���V�
�B;I��
��h,�ȓ-�c��Q��0ˀ'�чȓ7:	`���v$���R�dN�	��#=*0w���K�<��.L:"�jD��~�$.D�a�Ѷm5:���&�8��c�}א�҃�Z(@�p�ȓ;��
t�9ؽ�2$O:3"���'
�����_�{���WB�h�ȓi	�\I�%�.�r<*AM�]��f ST���� ��D��I<`=���^�P���Æi-ZB�8gZ��S)۳$,�X�+ Q�B�ɥ4�`��U%ZA�X0��AiZnC�r���"�Yc�Ȼ�&�r�B�	(!8D!�B�J���*R( N�C���Zڂd�H(d-P�bU�C�	3���H�Ϟ*� /c��C��:���뀊	'�q7��#�jC�1L�N�X��GH
qh��]��C�I �(AQN4/�^0q�� GM2C�I*P(��y�lN:o=&�A����B䉂N�U�'�"0*�'*C�{�B䉸O��([!dY�b�DC��j��C�ɻNS�%Ï�z��Oڇh��B�I�0FH��(�p�(�"��:3�B�)� , jVoX�E������W<$[!"O~Pr kL�"� \;`n�6w@�B�"O���v�8D�T9�eC��n<Y: "O�)At�9=�%������ܪU"O(\�R#�-�4`��ɳG���r"O���D���⭊�%��@�"OR�[<Cht1��Մ*��D"Or��O���$4���
E�����"O@�5�S�c'L�J�(� Ӽ�"O��æ@9G�F�Yri˭���P"Of�2d��7m���C�A�Z�"O���Q�Ҍ1R�Ar�ZmC��0�"O�Q -]��t*��CR��"Ob��E"_���R$κ!!�e��"O.IB5EZ7>������U"�Ԃ��IZ�ZT��*
�o}"]��5E�\�0P�cI�e�.0�4��A�<iT�B� >�mY�N�l��[S�G�.���8�L���O2dF��O�}Y��&"����-ߝdː�r�"O��� Q'Goj,��b6D��1�%�I�Byj�&Ɠ}-nq[ʛZ�axC cs���oR�;�����0=�iz�V�b�#�4
	�T��l
:tB4l��U2�jG�G.Ov����]u\X`5LE�<���D]���&���$]�z���5U�^`�3��, J�O���1�уXو$J�m�Dڂ�h�'t���-Ʃ��=�Dj�uWX鉊y�tU\��=�|�&剷T��8MA
V���@�So�<!
��"�t!�A�6~���
JNU��h��dȵ6M�a�V+�=A��Éw!�T?`��U@��@n l)@�07L�[��֨_�I�a j��ɡ���G5y�x�R��F�:����-(��W�N)ۅ�s�����C���iC��T2\{��!g�.�O�]C�S8 k�L�����h�W�d��nm�p���t� 	<
1٨��йQ��<,2�k��^[Ԛ$q"OB�#��Œ5������ؖv��eX�Լ�^(Qs�O.N��uQ�K�w�D�+X�?���k�t9�L����Eb���T���S���{p�'�� #�)N<�KyӘ��'k�� �)*���_�65 ���~�t; ��OH�х�St��Dˁ��(O�}� �J�2�օ�š�B�R�k����0U�偧�%+7�扆	v []w}�m�P�I�=-J4AʑN�8y�jR 1̊P�s���@��D�'ۨE0v#,B�V<97��/[��1�-څ`0,�
œrW����*�"`���
�1av�|7����T��#������Y�>*$+e J������]>�M�T	
a�8y�0g��d���C�b5N��6-֧-�ܨqQ�~�F��i2��CY�?�(S$M p��̀;\�P�SD��o�]D}bဵ:�� ��EHD~�	o}ur�ɞ$�*,��ԡJ��ѥ0y��Ab�i~���)C��]?M�(Exb��(>:�����.o�1�m���~����c=eq�`~"�_�;��nKd
qoZ�*PH��3���w6��wN*m���".S9bM�!<~⢩��I#tݲBA�,��"
цPa\�\4���T#���8ڴ]����u�jЇSgP�P|4�Bv�Ք4P�s��!*���$�~	N��P
N>L�xaW��G~�tID4f����t�i��Z���)@(��ּi�<�';f�(�Xw�N����T��N@��ߑ|���R�	9����@7�/�����O^���.�+u2�����.o��3��4Z�֜j`C:�Z��H:1�.l�ol��᠎#�O���j��T�����AmR�6����<�q��l~R��(w,��ƵH����S�0��Y��L�c��8�D꘶j��%�^�����p>qV�ѥ��4R��jk�ɑ2]g�M21�i�(A`R�iv�Hs�П@q�R�%�� �;�y���
�^�D#hї�y���%,oHx��́�� �&�D��Y�f�%~��@AX� m��q��%���N �l���?���E:a�S�
4�YX��B���2������>=��:�酑3H��I�-ϩ\�i$�X,C�Z1K��
���Q�3�������[zj��;P4��1� 8zլ��08`t��nO��Ӷ�H:� H���Ta�!��"OHԨbǚ�ڤ��ŹTW�9�鄌/}�%ÀJ�<YU�p�6�}��yC�1PFy*���/�����b�<���B�o��)�����شط��<�foQ���'z���Q-6��l�FF�ti�1sg�],y4�|⬝�v��ɇ8a�L�##�,^�|	dZ:e-H6,�H�@�-b ���N�:n�^���9D�� ½SS,�?7�$x��oŪz�|<p�"O�R��\�9�����/��"O <1�d�9� =Bf���DtSS"O�E��֘b��0�ȁ$F�4q#"O��A�d%I�\4Kg��8�2��B"O���W�ӫM)��'��2F�N��w"OtQEd�:m������Y�P�5"O� ��Rq�dF�&%����C"O\m!G-˫� @�e���);T"O~y����u��B҄�.Ū�$"O�DDB~��r@�ǁ|�|8�"O�|a#��z���� =>���y�<��ǧ6��t@Å����*w��z�<1P�����Q�b�`�`�-y�<�H�n�A���
cjh���Fu�<�%)�<M�YRj�=��yq�dDh�<��^?b��ǚ��f��Nb�<)D�F9䲭�� �<5�(���d�<���8�8�Ă�
�2��"c�M�<Y4A	�3���He��?~X(���@�<�NO�cqN�����[�|M�"IUe�<Q��f+.i녩� \�B��W@J�<��	[�!;�����6z ��w,C�<�Sn#o@�D��kK3j��D�ҁ�C�<��(��b��`
� �N�E�z�<���;-��a���x���{�<�Q���ҧ�DU����&Au�<��Fp��u��*���Q�Nd�<i���2�~|z$�T�X-<|��Oi�<!��=�� ��e���\���gJ~�<eQ
{T.8����{ �q�Jw�<��Ш4�N4bA!F6	��-�Ԣm�<!��A�b@���-u:H����m�<�E�*$aV�K�����4@o�c�<ɡNk>V�Vi��F�[W��G�<����";�&=)�'Е[bT��i�[�<A�<h�����������S�<�Wt�B�p�Ѻ`��Q�QFO�<��$Ȏ�8�&�6B�d��'�g�<�����/c>�yrNQ0"|Ń��c�<)u�Zz��P�����^�<�V��g������O9W��y��.�L�<�T� #��-��@0|�P�Y��@�<�uhU���% �Q�M����J�D�<��땕A��� ��A�uAb���	�D�<�A�1xB����l�#M�¹��E�<�!�TCFҕ���oӪ�2�A�<�D旿h��p�dA� �(6B�<16"أZ¶scP-�,t���{�<���0t���2E�*y� #cmZ�<�u�%p>�뒧[�Y�B��NW�<�W� BB�e���T�(��E#'$�t�<���C2Obn}蓋�< GLmced�t�<aF�D-~]��J��&l��:��Lj�<��,H�B[�������jX��2�
I�<�Qd�26�(��SK��@�<Y'a��7G�5@��Ռq�seJ�|�<)�h6����N�:�RI�,z�<qbɃ3m��hР��5$h^ ;��Ku�<�L�H� c�ǆ3b��ʀn_d�<���H(z�)7��g|0�����d�<�秘1w���'-�'{�-���Ko�<YF�2_F���L�"�%K5.�B�I�0Y����b��-�����,�B�)� ̘	���t�D0X��Y��Ͳ"OҤP�
=jj�db���=^���d"O��g�2�<}ɗK���v�j!"O�41�傫|�a� D8����4"O0]�ׯV;W֦B`n`Zj��"O�	�Wb�p�����E_ⵘ�"O�=3����R}��铗9v`"G"O�B­����P��D�>(�4�g"O(��f�	|Wh`��(2�C�'�L�y���19�
���.x�<��'��M�uB�?^�X�s0��+�X�J�'��"��B�J�F�RǪ�7kS�u��'l����9$d��v%ǜm�h}B�'+��l� �I��A�^�j�X�'��h��t_8�qA�� R͜�k�'��P9gU�Rf��c�J�TBLyq�'�V�!��ԧfǔ��fn,A��1b�'�@��Kѻ^Y*�0g�b�x	�'�����O�'V��fڟ3�DA��'blH�m�5�b��؊Z��mS�'���装˒Up�x�Y!��h�'Y��a�
)<2�y����4|i�'F(�2��{.��Uu��]�	�'��Q�6�P�A�6�Q���h�,���'����ӈh�hpH�c�0E��'���!E�Q��y�!��f�����'
�A뷈�$���A-̖R�� ��'�ԽirM�09D=�֎@!����'�D��1�@L�$4���>BN���'dDA�ǆ�=��0'+:	$��'�8� ��=���t��)��QR�'�4	�� ��U���OR��p�'NZ�	Ğ�B	2�{��M7���8�'���9�&T#8(=���F�M�t�	�'9�I)&��,s;@U	��۵8��pr	�'ö����fWƴ��_�>7�< �'���9*ۨ\r@�(26��'�.Y�N��l"�� �ǃ^Ȉ���'O$@�a�0O�(��Gb�NB��ʓu��a���#x���ݥZ����ȓoI��e`�}��=��edф�_rBL�0D�g�T,qqÐfʶ�ȓQ��P)���mY��|�
i�ȓNy܅`�hg��������$z�t��A���ǃ��v���&���ȓ<fx�J�k��Q3�h�v.݌J-t��}��$R��P1�8ѡ"]�B��4S$�ᢁ���b��S��t�\`��#�2=ȡN�6j �p�NY>����6q��) �weʈ藇��-pЩ��G�ԡpׯN�EȰ�����Ҥ�ȓ*:��y�D��ɥ	�=��ȓ-�Vx▍�� ������H���:�nЅ�ַȸ�EE�;Ӻ��|螰XfkP
+B���
X�~9��s_�t�SE=����(޸n�>�ȓ ~���b#6&G�IZc�Z7#X����=B��CA�	�z$hߟ݆Ԅȓ5V����ˠdgV�2��ŖW�%�ȓg
��:$������aN�B� ��{�
D���CZ$�V� 9��ȓc�\��ĩ2a��0��ɞ�?�����$[���␢N)�e`��"ޭ��&�Bd�⇗�����!A|,d��S�? �4J��\�I�&@�vU��]c�"O��2�(̙[��ۇ�L=�ZD��"O�(t�P4�8ňD=KT�Ĺ�"O��B�Q�D�B`!�ꀱ^f��bT"Ox���Ι�1 �ػ�ʃ53Q�9 �"O�9����	d8�
�7J�A�f"Ox��P�8�yu���$Q�M�"O�h���˘�-{���TJ:�"O!�q��9Kx:�i�7��@��"OB��o�L�6�H��5H�*�a�"Oj!J#�W�Y&0�S�����@9�*O��ys�t|�� U�\�yb�̫X�L�_(�R����9�ʓk�^lFNI
m�FUDjӝ�4��K��t�M��(H�]9���'��]��<F�\;��]�nW�D����H��	.j  �cʵ
�����>�B���� �za�&b:<#AI�?���uxp�ō�]�l��dEX�i^q���$xō��o�Ƭ�� �Q��M��6��q���{��}R���e�n9�ȓG!��jgaU4%�i�Մ�|��)��@i����Y�<#�"D��Y�ȓn�Xѕ�\�P�����vP�ȓ�Fԁv	�v��%�S���{�x��ȓ-�vɻB@]�X��q�$����ȓ^�ڕB��T�[]�<r4�Uת�ȓ4/*�JTlm�V�A0�Z�Cr���fhTiҢM_�)X���%��xd1��C!&�a��>���'��2�=��@b�l ��I��e��@�f�������glȍM�X(�s��<ZT �ȓ�A'.��=�X���Ǒ~����]�`����D ��
Tڱ7&�Ȅȓ	��ɖ��H>��6i�2]�<Ԅ�3#���0���{�����k�>!��k+���lK**-��sC҆A�܄�q�`�h���H(D�ط�������ȓR8T��
�3����FR�fŅȓ@]]�SCBKF0�Q���Z�х�H%�2W��8p�L���%�|ȇȓfs�t�F�[6F�p$,�'_����(T�]ꃧܔ6���/�>���/D��Q�K��x2!c=R�ސ(T#&D�)`����u�u�� G*����$D�����#v$�i��rk��#D�����7T�����ǉ{-�X[Te?D��� �f(\����
W���"(D�y ��/����o�OG�(Y5�=D�Ȋ��ިNu܌ p�l�fـ�N8D��E�b�b%^#/vٹ�m*D��Y�-S���ڱ��YXy�6�<D��@ �ل5{�ض�ے�"r��:D�xP�2@`.��	����2�6D��0]u]0M�g [�>g �"'�Ң�yB
�H�i!"L]�-v%y���y��:�$ a���~a�qA��?�yȇs���"`%�*\Q�&	��y��F#ι0@k��Ⱥ�L��y��V&a˪�9F�K�Z�������y2���l6�d��`�?!�ej�,��y���*xWx�y#��2A�(+���y���B@��)��xZ��@f*��yҌ�4'PY��/=uH�Y�Lء�y
� B!借Ha��7m]�X�"O�di��;j96	�lV�P��D��"O�a�C��Xz|���@ �����"O�P��m!w��MB�)Q;P!�A�s"O�a���?L3$aj��I�z/Z���"O����H�۬Q$�1;-�s"O�(����)]A��	7=�q"O2���d��l�wIEA�s�"O�H0$"H������@-vf�d١"O�82W��9v��A�ʖ!_���W"Oh��A�[(-�P@3�5$FĔ "O���dO�B�����g����"O�!� ҙ%
���Ș�~���#"OL5�6�>g�2a��n�h1�"O��y�ѻpE:�C �N	����"O:�[A*X�a>6���9��y'"O`�KE��<��vF�:	z=��"O�� @<�Q�
&d��V"O���"�G�-�=�4d��z� 1��"Oh4Z6 ��;~eyg�S�{d����"O|�#4��o�
U�R���d�	P"O^qC�۝F�\mh򡓌z@�q��"Ox%2�f�0=Px(��Qb]�"O�����ޗa��q`�L&LLe"O̹C�={�נL b�J��g"O��'M� UPW�o�ȥs�"O�$���X!G�����h�:�0}�*O�Y�Cけh9R���/�1gج
�',LD�dO^)~�r���a��O�,4�'�4�CK	�!�^�sa�=����'P<�����k9��EȖ�t �	�'�@���n�6U�*���cG�f8�	�'��c��.'i�%����|�'��Ր"I����#,V��	K�'�8MSJ��	Y�Q*E"�pV�d��'E�L�"���H��(��n��o�@{�'m^%:3AՏ{0�;s�I�_10���' &���A�N� �����<$�0I�'�0�əH%v���҃1İ0�'�>�jv��:5�fy�R��5�8�!	�'�t0	�&��
�q ��8�EK�'%cP����I���E%Z��'��#�N�4�Ba�$�f�B�'�~�P3��y��a9�*ε.⹢
�'��r`�02�01%����p��
�'���$B�d���
5���	�'�v�����q���7�S103��*	�'Dh�S��H"�!ۡ:QR`*	�'�����3�"�:��ټB2���'fP�ԢW;G�����$׽,��	�'m ���C
j$�d�W�>娑y�'1�aʲ)9rPp��W��n��Eh�'c�9p��n�
���(ZB��'~�CVM��e( A��8=Hhi{�'�0�t��Z�2�U"G�$}��'�D���Y�r�j���-
V�-h�'���a����XP�݀B4Z�
�'��y�7���C$G�:)�.�	�'Er�� �LV�$��'�ּ�'v��a��Um��3e�ΛK����'�d��eҰJ�����K%9hN���'%�� �(�t��xAt�R�:^���'��U ��Iq �:��_0m0�I�'�+5a�2n�B��$�L���� ��s#�
`X��iŃI�>�0�"OȨP@�r��$آ�_8���Q"O��Z@ݝ{ް��K�gv��Õ"O`y���R
�@�*
�g�(�"c"O��{�%
�d���7%|\m��"O �P�&�pL�5�Q!pZ�9��"OL0"�ŋ&k�(1I� C8i��"O�mڕK�iN�r��W�~�I�"ON̪���/�	���ׂ-�L��"OP��ĉ��49��U,�)d"O,�E�N�xVFu���.i�x�R�"O���K1i9(� l�.�<��"O6h���<	�K�3/@U"OfYY���B��MҢG@ b�ȶ"O2=����*v \PHdf�k"R'"OVm0�F�'(Y6�I�.)4�[7"O���r�*!L�ñ{��j"*OF��a�\+�	+��=V��a
�'�*I�j�1�XX��ȎA��E�	�'Xf���ϗ
}���G�t��z�'H�|p$ϟr'�RWC
N���'��\ v���)�bѺxF�	�'���a��	qr��qw���'m���2
�|>25A����^�n	�'�����AXA��qS&��7Sj�$ �'����4�-4અ�$��[dz���'����-ޭ�e�d�PJ��3
�'-�@PSf�&�����Ŵ4�dJ	�'�ʳ�E��ą�=H��'Rƨ��bH�p0T��,��H��'Zhh�i�PNv�2�D�	SF�mJ�'&��#@��P��b�D�TL��0�'B����J�$7�e*7oK4Wɐi	�'�:����;L��f��g��Ek�'��Hcv�E�
dr��G8 <c�'_)@rH��.���$h
44�*��'v�(G(HeK>LbD��#O\�z�'������!�i!C��Q�
�'���!ႌ2����B��?B!X�'%��X�/X�þ�hR+_� �,��
�'r �kea�/D�t�iܚ4*T�
�'d�e�檍;|������!;2r��'u��H"AS*B
䐣�
�?ʒa�'j� KPޅl�@���K:3�q�
�'���Q��+ �5�EOQ� �vŀ	�'A���W�Pq eϹ`�b}a	�'U:t
����JO�3�B�d�\���'+�UVKɦf��D�Y_�,�{�':���tȜ)v[ܠ"TJ�F=�p{�'��Q�`� C�!��p�'���#��u,^y�uңsD]��'N�V�L�
��)됪HR�'z�yzFg���T`���}g����'id�إ�Z#k�8�(5-�2l�p���'���1�3�zh�с/p�jP��'uv,B��Yg"�2���d�T@��'ٰ�x0���O8zSҪ�_p�-�u�ڌ ���tC��"��t���"\֮� �h�H6f=#2:O��C�:��%ʟ��t�7�ԗw��9T��[���y��|NyqaG(����J�#1V�ؐ���T���iZ����)�'"ݬ@�@d�i�01�� �%7���oڕhQ�"2�` ��b����#��ēR�`�'��\}ʊ��4�'R4��
�5L�Oԣ=����(3�G�*�d�XA�Ř>Ô�yp�|R�)�ө�NMr1�S���9n��"��hO�T�?� �y�&�"~�-��bX������'j�#=E�$F�;��� ��O%�Z$�¡��Em��Fy��)��"�6�Jqٶ"A*�x�$���%_��ӧ�7F�xK��x2�ǡ_�`ʐȤ��8�0|�
�E>"�;ԍ���R�B��Z���'(\� �|h6.�r���ز��'��p(t�x�E�OXe�=�~���I�b��a-�3ú�R4�C/�O�|��' �x���"<P�
�Jwb�&(�|h�>�)*�S�,C������	��*��Q�SȄO&-Fz��4���r}tiA��46���S��3��dKZ��(�b�X%��R�P��$ŝ�Tl|����'�ў�~�q�V7J`�a��;x��M�Tn�'�a����!7���圴k�<T´k�3��'�t#=�����I٤��x�mA�2��c$�x" �B���Oy��86������aѮD9��ʬO�@����i&<�`K��>����0N$@�6�A�#�T�«���E
H��T;@����+=|9F�ƭZ��x
/��6��"�jذEk���E����i�	��H[�i�Xx��)F�-(!�D��,3D=�w!�/kA�M D��}�!��X�]Xv����T�c���!�ę����g[+6�9���
�
�!�$�=e�a@��+P��0*�`��!����e�-��� Q��+�!�E����qN�5 �Z�CY�=u!��{�Xk�kQ�w*M�Ee�H!���*`a|A:�F��q�E�\:A�!���%+g% s������}�!�[� ���]/4�ŲT/S1Kn!�䒯M��0`�b���zeq��yW!�$�,*�$(
�ݜ]��Q��j��%9!��N�g;:��w�B;y��%�W�=%!�D�f�r z�hT=G��I�(
�m!!�Ė=�����#
R'���f�W!�C�D�n �!e�7;�� ����<l�!��mX|a v�F��D��*��	�!�X�A�0�I��l����g
�8�!�|���s%Ȥ}�X��gj�=�!��\y����-ħ/�N���鈭SE!��)i���#/Q�L�4����S!��80@h Ƙ4L� �����?/!�$��#�`�S��&q��+FÏ"d�!��|����NX�}e�ɂ'��0�!򤊸q|�P��U52\�)21�ѥ@�!�$W4M��a@��4YxD�I�,��+v!�Dn>���v���ek�	aA��u:!�$_�d�rѩC%_Z�<�A���Py�L	f@e��.���`C˃��y�Ƨr��ےKI�q�t����y"Cؘv� )-�l�
�['���y"
T�bv���#Q��pG"���y�N�$+����G��  [�HѦ�0�y�'S,-��p�n^=�P=�0�;�y�Ê.\��5��睶*�B�WN��y��e��l�� �.Oy8�C��y"���|��Kuc��XP��cIY0�y �f��l��5e�m	v�H�yBÑ�W���x�k��� /�p�A"OV���Ȅ۲���*֪X\��`�"OH$hS��:g��͊�O?�D��C"O���f�,2��*NT���$Q"O�����l;v� Sg�#p�t�7"O2��#�,H��9�p��+_��$8�"O�Maej�&�qѤ���.���"O� ��%���#�h~^��T"O� Ly��H�O*�!�Ť^$��C"O����$yŃ�1$J�4��"O$�P,X=��C�ɮA"b�q"Op8Q��t�t�j�c{k�i�t"O����)W �Nh"�`¿B�Ve	�"O�)�Jʠ�R�Ư�);��hIq"OX�¶���L�sq�I(j{��;�"O�$cvCس;�R�Bn�\h�5rq"O���e��bP�bΟ��fqBr"O�aơNY���8v
�x�銐"O  1��\i0�[�gS�4��C�"Oj��dHҠ"�\�-91y"��"O����^���{���c�`�%"O*���Ϧ-�`{D�T�9���w"O��
�넝e��ta�*'�Э)"O��E�%`8�غQ -z��OL�<	� �F6�5�pIʺcf���*�M�<��'Oކ<뱨�+<x읓�cPI�<7J�"3�}�������㧉�H�<Q0���B���-ю(+q����_�<)S�/bC����GB�b��&�\�<���+.P�y!��U'*�Yw�Xl�<�V��_T����j"u�$�j�<A��Q(O��0	Ε�-#4ȳ��m�<�����"�l�§O�1�J�����t��Pg@@-~ڙ� ��6? r��,�d�
���z�\��`��f��E������#5�b�2p�"C���ȓv�8�"hܧZ�0Ղf�U
�)��:��23�X�U0)@d��w����f�@����3;�\s'��
EHe�ȓ*8J�#nA�0�����L:z9��kk���Ԃ##Qd��/_<G�Y��P��T�7�J��,�� G1S�,�ȓ>1�b�H�mE@�`�L�0uX��J]�e`�`Q"J�@��ë���앇�#�<�j���7Ě��� �L:�@��;}l�p�f��O�^�HR�
�y:dP�ȓ+o�y�v��u��x4%z�n�A�<ـ&(6of������V:�Р��F�<a�c��3�Dڰj@�	Ĕ��'�{�<qTfΎr��0�j$Y�J �'�p�<9�	�=/�,ዓ͞ �*�����V�<�� ��z����Qbt����A�-�y���p����^�c�ҭ���y"�	2�쁣����U:6@��� ��y�� /Vs$P8uL�H�*,"���6�y��Ȓ"L�(���6ᬘ* ���y�ق(��9iV��-̠�p��6�y2��Y�ze�&ݱzRjGGF�y�K���3 c�r(���ϝ�y¢߹r� ���ꊸ}ΤM�A�D��y�戽j:�0��U<?�T	�A��3�y� Z�0�,M9�#N4�Ĵ�����y�C�!L���cA'���rdX5�y���?#�����,Gu�L��$�yR�F�h�-@F�F�D�= ���y�N����6��W���>D�X;���@l|�s%�4Z��=D�:���B��|`Pn�"���D>D�<���غ>�KV�>�n1�ea��R�!�'I5���(U�� 
E�H=5�!�$@43w~D:!��=	��	9V��t�!�D(�R���ꏈE�ȕ¶��%�!�� �XQ��Ja$}�S�]�W�@pұ"O�TQU�ДA����#�t��$�"O>v��ksVX)2(ɰzXr��C"O��	W��$k�:��'M� G9D��""O|H����t,�y� 	�D"�E�"O���bi	2(�P�F�N�Dg��""O����j��A!��!���'Wbp��"O-��i�	�B��T�Z3D��[P"O�ဇ�=P_A�c.G.N"�96"O�0a�f��K��~�6<ɇ"O�+�H�D��2%�`��"O�����C:��s�웱l[���"Ol<� C�4X�� �E�ذ/���f"Of��hHRLЇjڌ:�L�hc"O
 *[08z0�Ԯ\瘥�d"O�`s�㞖D\���I�Vn���"O���2kȉ^p���m��|e:��E"O@�1������eŉ;~��m�T"O�Q��F"�^�"���~�i�"OfԀ#(�Ms4���
��6��t��"O��j���A�l;5�֩\�y"O�Lёb!��	���
b����$"O�(�Վ-����Ј�Zؑ�"O:�uLC9P�H�b3#�4]��7"Or�b�AN� �������-����V"O|�RM�[���,�l�؀"Oj$#Q�m.�4iP�H3)K��"O������=���C����,Dj�"O��ȃ��]v���5P-�|ʵ"OȕX�&=O�L0J�l��*&�$�p"Ob�k
���q����-�E"O.�QB��� 1CٓD�h�"O��6�ܨa���)�Ed~8��"O��ȓ�Bo���@Ls�1
�"O�d+ �3r:�r@N�)g����"O ��c��]`�S����A��"Oy�Ő�_�F�ĩ���d�0"O \���Ƅ]S||�"�6h7����"O���
8h�M�&�\�OW�y�6"OP�@@�ȟ
b�4�F��<j-���t"Od�फ��c��)�#�T$ 5""O[�J�=N0`H�rIF�����"O�c����1��yb�i��>����"O��j���Br�| �j�5��y q"Ox�!�б0!���� 5R-:y2"ON�1�L)uԶ%j��_2Jܸ�"OpW�?8Ҙ�kvhNK�@X�)�E�<i��� ��@����m��`���U�<��2y����m(,d���� P�<�&�=�Y*��)���*u�K�<9W!��u��uK0)�&@�����AO�<���W$b��)x��PN�<����>`��p�づ�rZ2n^K�<a`k֋z���!t�Û ��i�kD�<1i�i{X�1��6v�`�H�{�<���A#6،A�X�Ro���@�u�<��*�	Zt�rF�����Ѡ'�s�<��n�eD8�0��.r�� �Yz�<�$�q�~A��쑨��\���t�<���	��}�f
վf�	Vd�m�<yֈX�$��g��<rnj1a�̈^�<!h@�=޴�!��7-m VF�T�<Y��a̪\���ɲc�.$��ah�<	` ݎR���7�\�D.L)���d�<� �xy���RWB�6�LVIXDqr"O�y[��Ll,�E/��;9��x�"O���#�ʙ$� H�VȔ''d���"O܄�G��0�F0i��K�$�2b"O`H���֠NOH1q4��._%�Lc!"O��iS9��8bG��0bp�d��"O|����.|9�āG�֒i���s"O��dWH��j'E�+N1�i"O,��t�&8�����c�] U[d"O@�k�Fj`���@:;��("O0=�U��:O�0d�p��e�ZY��"O��R�F�<X Q���٣p�8��"O<���FV� k�: ���g����"O�*"c��a,��+�6&��"O���i�8�HD�
˲.V|�0�"O�4+!
�	[�ty'�T�P1�R"O�1;�g�!|�	#(^�J3�� D"OT��"ʝ=QrځP�L'����$"O�q��-���F�G-�_dT��"O�0��艒Hx^H��.޷i&�xaU"O�t�4m��Jխ�= ��0q"O���5+ĩ~ ��7m�=W�Ȁ"OD|-T @  ��   i  �  �"  -  H7  �A  �M  Y  tc  jn  �x  ��  �  ��  �  ٩  Ѵ  �  W�  ��  ��  d�  ��  %�  h�  ��  ��  2�  �  � 
 N � � & Z, �2 �9 �? .F �L S Z g jq 0x *� � � %� g� �� ��  `� u�	����ZvIB�'lj\�0Ez+��ɰK*�ac�'b�T3���|�W'Q�H ��M�7H�`��?4x�3����n81����W��T�a���v]P5�Ѫؐ�u��[�(�t�>8�����]Q^u�#�T�z��U��lE t����Mq�6MB1윻�˞�<��]�p��M�S��M�E/)�D�G�M�u��:�_�`�Qf]#<F ����n�6-�$>�D�O,���O��d���nl�����@�e.�	ED[+m[�q����v��ܢ�O|�������韆���O�P�����"`&�aY:�����Od���O\�$�OZ�$�O Iٗ��M�pړP���A-J�fQc��"y�Q��^ո���dP�Zը�<Ѳ�K:f0�ś��˻o�8]�fA5)&���O��{�\?�t���=�v��(b>�# �--���O����b�B�O����O��D�O�l�֟t��V��0���@�TX���[T�`�9�'|$6^ɦM(�4A��v�'}6����oZ�t��G�x�<h�0	� O���gJ��o2�a�'�
�DB�j��!��[<HJ����Ԙ?%ޢtZ�6&��5��&T�T�,����Yg�hic��O�mZ.�M+�'��D�O	�ڄ)��(�ӧ��6]��*Ǝ'�7́�Aq�Y��ҾN�HUh��]5S�YW��5m��o�M�G�i
��!�d�&B�	"��"I��`ܸ`jD�&a�P~��۴|��`x��M�DO�7G���$�*�� �#
ʎO�<��#B\�w�P��oS6~���N�>"4��q']���ش8����ֹ�Ӈ��}�*$�GǜA���1��~,�a������В�`{��X��Q�3t���@Y�%Jh�D��O��lh�X�j*�QÓ�B57��YB"e�ğ��?����?��ml��?=0�ꚲRmxѰ�`Ͷ�i�3��O���?��?��	h��1�(�C6�L맆�7P� 4���øQ�h)!�L/m  %�!�;13�4FyR��gǶ� ��V�_L �s�B&
^��A�Μ.}���zR 5uh�D�� .�QGyrh���DZdy���� b��gl��C���?����?IO>1���?�.O��_��t9�F]�<��=�׶5H� �$�OL3�e̽��O��9O����0����;����*�&6���i�O�ʓQ�*�C�i����t�q�ĉɈ'dMz�O�8O�D0��OZ��R0������i����ˏ�����ɢx��� _��p���7#L����/�'4�p]�'|�J�5_:�Y��:�H��b�*%2�N?]�A�F5 �8
D��=>Vm+�<?Y$�^ğ�޴��>��'Zc�Q1#�M�^��&�n�hq'��IΟh��П,E�ĭ� ��Pq���P��� Q����hO�����"�4�y�iq�I�t\�;$ɿ>��ts�/Bh�6-�O��X�����'�?����?	-O�Z����m��L-=��k�P��A��!��m�r�P�>� t�+�|Z��A��D�C�Yt?ɖ��r��)�vEX�vs���%ޤT���*�(_9�u�VgJ�Or���|���ǑO,��j|�`1�ޓz����.ē ��0l�;��D��u-r�O'�3��ǆ]D@4�!ƞ; �yµC��gP���'�S�O 8�� B7��H��Lov���'&��{��mZY�i>��~y�-֢Q�����H�k�L�wh	rZ��u��>i���?Y*OJ�'��$$��e�	i1�#��=�VF8=n�١.�0��qn�A  Ub�![�'�l	Ey"lۍ0x�ErG�}�R�rc���3Q&8a�!߷@2�h�T�ɳB:dI�Oȶ,�Fy��R,V ��ub>c�L4pD�.�d�y� #�Ƃ>��O�)��#�XN�Y�$X�C��j3R�@EB�DU�MO,�ãB�)A1�P �'C<7MDԦE�'�h|��s�@�Da����H�*Qު��t�F,y�& ���Ovʓ�?����t�,H��H	֠�M���|]���C�"Q@���MI����C�YHv�P���^�,"�;񠅘r&f�4eΒm<�A��- �Ef帥�@��l�cV<��aG��o���O�-�?�p�i�7�On)��������@|�.��¢<�ߴL;b�|��̸Ot}��]�&�4�b���*}�bˏ|��'���>�M���F+!h+P�׮fe��v�t����'E�7M��{���{Ă�dR��rw�i��� �*4���h𨛜c��2'�5J�"�'�u�e��4	���7�1$�Xi	coVEܧy�j�A�읇]��<��F�(,�Ե�O�������a6`�*��W�hH%���ێW��"�V'�z�	�6Ov�бB�kj�9�6�Χu�I����$ݦ��N|ʋ�T���I�ɏ!-��,�$����?)J>a���?+Of�r��W)}4s#	i�~�!�ʘk�'�t�DyӚ�d�٦�� W����a�e��%yw�G�s z�4�?�*O�E��
���$�OR��<��gӎLw���� ���٘$Eʚp��pߴo��HK���y��|��'�t]9wC�I?I�$
�(ԄY��a�<�Zq�M�zD)�GEx��P�*!����C���P�ẍ́`ˠ0�`���[�ޜ�`#�[�� �"tӤ�'��ؚ���?���?Q��ѳ{Ϟ��U��	%�
d¤�
��䓃0>��O�eP�� #Y�D�:�e��꟬����MӁ�iq�'8��O;�I8�������	�^AK�m_�=]j�"b`��M;���?i�����)ׅ2i��w�ƿbXJ�z��
0���$ɹy��d*!�Kl9�`.C(8(z8�t�I��h��Eܪ(� ��B[gu�ȳ�B�*k����K�Tf���4N���X�O�fq��IJ>a��u(R�xp�	F*lr��&�X��IҟX�I`����ֱ3f`�Mc�+Qg �8��e��'s1Ov�"Q��(�����PEt�qǛ|Rzӈ���<i�4ћ��?mp�@���bő�
	��{`"�O�˓�?!����Ò!kq<0�!� - ��H����ڀ ͙��:b�|ɧ��T]:9q��\98<Ҋ�$:�4�D,ڝp9���D,٦%��ǜ-9���B�e_�	��A������3C2*I&����L�O�Dn����B6����ˆ�Tf��Q���%��'�	o���hiՁ��,^��(0�O�,@�F�pE{�O����:m��Z��)Y&����� y,6m�<���Ƃ(����'d��I��'e�ՐWEQ�":�is���+0Rx22�'5"�Ʉ�����/	|m�V�ܒ2S��?���ʖ-d��t
��ou\�B#�!?�t��19��9�Ď�	7�˦k����Ob� T��'2fM���\a4�2�Oj��4�'q���ܟ*���>�n k��=m��X�@��~�<!���9#(Nٺ'��4]�-J�B�'r�}�YB|[�g��z�@�2�U]g��lß`�'g�A��O��'@bW� �šB6)Ō�Eỏ^��Y�7,�Ny��'&���'��iC�&�0�<�k�%B�3�HU0P*R/$ސ�@l�7Oo>��CZ��O�\2�O��� ��
���`	�� ��x�$�'�rL���Z̟�'��Q��0��t��X&�:4v�'��X�d��S����dV�J�x��k� f&�{� Ɲ��-�M�׳i	�'r��˧��,�.�h�b�<�Œs�=L��[� �;dH�lZ���I۟d�'���|�ʄ�0��xs�
�e(vYNܼ7�\�����"��D�Ae��U���G&]�oI"��d
wa �iL��`�f9�rHE|d�J:��	Ǹ\�r8yrl��je�1��[���O4ғ�O@�y�.U�".��wB.1344��'�!����,ab	Ic̪h�D��s�4i��'n6���M�'��(y'�f�F�Dq�t��)��x;�]r���,S��kS��O ��?Q����S���?�`�^�(�*Ɛ1j������0<��o2�DыR_-r|�P�3f��ׂՅ3�qb��E)�Q�s`�C�'�\���:��V �<Q��Ny	�q���P�������O��a��r�I�3T ��m��rL:7%�<�	ߓL����U\��Ѩ�T�⒧66�<��
���?����?I)�x�Va�O�h��ĹFw� ٗ�K*7�2D���O���K�J/js��O[(��m�
@��(Q	
`�a�S�|zd��c��fH],�:�J�F~�A��v�ݷ4��F�˘�*8�R��)׎�0" Cl�����6���؄Gx���FlbAd�W�2c^��}8!�$�.2�n!�bǞN\�4ȕ�=�џ(@��遢q:��� �7"�l��LO";6��O�˓wV��9�P���I���';�?2��i3���9��PЁZ��I+WZ � �'�`�y��ǽxx��9�ɒ)^M���6GK�p��p�3�]�ИO�\�� X�����H�F$��c�>S�,CKR���+,O����'"�$�?�OP����;R�Xe����^cb�y�#�Ik~퉡Rh�M�$C�Q��A�%չ@����Ge�D��香�O��4S>����J�R�&�c0È�M����f��Yw�� �O~���O����f>���#I>0�t����l9��Xe�I��q���ny�YsjͿE.pp (��U�
��\<Ֆ@j_�ҬF�24g��cs��B�'�-�.�PΥ)S�2p�x��nR��?iE�i/n"=��2j_�����ڋ\�#F���3�R�'SB�'�0hٴ�ڪHM�vg�}审�O>)��ijB7��<G���?Y���?qJݎl��s���X��Q�İ�?I�yf҈J��?��OE>Mڔ���3>��SBC��XǛ��N�Ɩ	�v��J������|1"|"#KT�(O�	`�&��Z�~P�G�H_�6�X��� ���?f�xB��;�V@�A�%�]��F[�ē#(JX�	����'��}i�N̉G�����J
hyR��M>��J�VT�e+�0`��Q�A�J́��ɗ�?i�*j��Mb$�"��|���Vڟ��'�&�(Q,n���$�O�˧q�@���0��Q�<�~&�"ci^`2���?A�J��?9�y*����k0��	%��"'�99'f��'�����S:$�����)�&](�%�u%>��N�P ��c�S�O�4P�`+Ȱh	6���j�fM��'�@�VJ�9s<n<huƆ aS`,���D�>I��55�,����"�ĸّ��2���R�4��$�\A���?���?�*OȭZ�$�+34� ���1d0X4��H�UX	S@�D;}�R�KV"�8�Rb>Y:E������O�kS��[���qh,%2��2yx44�dbѥ5<t���a�	6p%�u�ɘ99B����'p���Δ|>({5�̴0�9��i���d���I�?���I` 4k�#�V�F]1h��'�� �D�1t�=�4/V6r�t�,O.�Gz�O�b[�����W�d)�C@��d;��(q"�������	�����u��'��>�d5`Gݗa(��)�j(0�r���KK#lF�yit$��Qٞ0r�[&�~��%�P��(O�y��� \��5̀&	u�-��Q����!U<|�8ӑ&����&mQ�,F�y��
�.* .�$��d�� ;�H	NQ(z�"\�i�UZ��DԦ��D:�w��y�,�'~)j-P��<jT�x��mn��+�*΂E�,0�MH7A{i$����4�?A*O.�Qu�_G�t�'�"�j σ�4���S�,كw�R�J�'�r�G)w���'��I�~�,s��ՋT��8K4��3<���w��_�>0�#� �K���ʅ�EN�̈���R�����J�h�j@ˤ`Ɂt��ЅB7@��T�.�ZґiКm\�̒DӀv�t'�p�%'�O��mZ���gW����F8gVI_�H�L>��D�T��Tn�;Q�Ź��ҰKܜl��		�?�J�8��9���R0�
d��̔'٥�'�b�'L�%v�R��IBs~$(dЦHwT�)g�ǐ��Iڟ,
���E(�@�r�@1u~�^?z�I`���_��d�CLb%��P"/�������dû~7^i`�*őVX@ �nE,^�\�C�"���S6D:���d^O~r䰗B�m�f���x�	�D�T3O�� �P����5ޒ8�p7"O&���!��Ցb@�5@>uA��I8�h����T.2�`�"�Y�d�L ��i���d�<)�,Ҹ����?����$� X��ZF-����)���ۺT�
��?��͋��0=�Ƣ�;Z؍J�� 9 h�#�2QD0 "�Q4�?��M�,|��|�<IE'ַ.ⲉ���]-D@�<s��M;ES�42e�O���8&�|�tą�Ep��g!x��h��ɖ��d��Jy�'��� �fk���2,a�DL�Pn(͖''�6O�A$��S�?�'���#%��g'�в@P<9��8B�Dٿi�tP��':"�']��fݙ��͟�ΧL�B� �!Z�1��ڷ�}�lx�$^�b>�(0I�0F���4돞QJ �`5'>ʓes�� �z�:5k��2*dPSk�T �;+]5hݖQ�Ř�ep��/ʓ8����2xu"L�1GS�t�p�P�" �� ����?َ���;6���sKڥ5�m[A�AZ��{�ăh�Ȕ#1�߷A� ��q�!i��'�7��O&˓!l����i$r�'�8����
;l�Z%�R�X�kL���'�2ٴ+��'a�M� [4�E��XY$b�3#�0Q�D��%��m�`-��F&tJ��'.�e���V-j���1���qQ4�{��ּ*K�0��[��t��G�	XAs�����������'?
7��OV��d�D
T8��5�E����<����=���͓B�|����4Q��b��V��O8�=���M� �P�t ph��-�M訝�0��	m���'!�7�=P�2H��*�O��D�O<�i�4�>���:�������Q"v�sƅ�E� ���On�`Ƅ5F=R�8WF��zAb��D�ԝ?]�4�����GƏ%���&;?)5��(-f��2�+R�H�*�!G](aJ~rU�7ФM�	% ��&Kr~��?y��i7-�O�"|:@���m�Ҕ�K�	$�k���l�I̟T�?	�yrX.X-qr#S�u<��x'*���O��l�;�McO>q�&ς:��t��.U�r ��Q���Fk�,����?��P8�S���?q���?��Lj�N֨E�k�6q��Hrc��EȞ,��)�XѪ�A��$"Qd$��C�(��O\���7
x[�.��BP(���	�E5<���E�7��\��DR+81�䈗c�0�~�Ƈ�;%�����[|xؒP �?)�O���%�'�B�ɝ{��أ�k����$�
;(�ȓO�&��1�?U��tB���@�h���۟ ���4�8�Ħ<��yv\��q%�?Q���q�5��8@N��?����?���}��n�O<�d{>}���8<^EK�Ɍ�	7�i��K�X�,�!ح�&X�s�пD�V���f�8/Q����TS�R�'��%X���M�d��`8�Ɉ�[*�yP�00:EJ@d�F���;��	����s�&��!��a�cN���2�LvR��ԧ�'���+c>����H���fb�l;�$�	Z�p�8�'���4���?�'�i�"�'�� 1pJA,_�D�C� `�&`���'�B���9�"�'R�	7g���p���P���S���#7m8N�@����X���KV �q!��W�Tx,O�I�'�O�D!�+S�Np�Ģ��'�vx��}��#�<�Eʑ5a�MS/гk�ވ����t��Z$��'�b�'`=O���A�2{m�p@
��g�!	g\���'�ɧ�O9��G:)Y<�C%"ωN���XFl��XU����D�6�M�����|ʚ'r�ug͐b��i�U��^$���OR-���)�'m��US"n�d���B���j4p��'�������� I�B�+�R�kG�ܒw��I)V^��}�)§�n�AW��, ��t2�b�L6D��R��TR3o��;Y��2���l�F��2ڧ\	�XX��k9����f����ݴ��)��]��'�?����?*O.�I��+&wp�{&���y�U3����4�PeqM�^V:�"��T.�Tc>%'�X�6גw E��5V�����M,x���?H-�{6/Q��c>&�� jQ`�b�L�3�NAq���7�'��I+.��d�O~��>���U؞H�DB�]��T����=[	�ȓ~�>�	pD�,#��1���Ю��t�'Mr#=ͧ�?-OD��ŝc�j�X�X*8�	��̈�_F��lΟ�	��\���OGrq�� P0!� pq�c �*��m�r,�!@ڵC�]W踩#lW��ʢ?��¶=���\�Q$e��hX:*�D����n1hy�fGV8�n!�2SY�\#�᜖GT��i�AH��HC�'���'�O8#|:��"r��n�Z�e�6��Mk�<��Ȃ�6Y�UN��Q�0��2�K^�I5�M+���D�'.�t%?ձ��5��Xw��w�9`�-�O�ʓ�?y���?a��*3M�s�Y;py������tCq�V��Ae��8����c�	�}y�I[s�([�<l�E.$��0���3<1sD�1Jк����h�'L�@��?��O��𥂃_$�d�@��0J���3�|�'Maz"��oA����$"�I�&��?I��'dTPZpǓ�V�X!��$�u�ƍ����$�=/m�,o�o��}�4�'
pu�n�gl�X0�Ж0��1@�'�r�L�<���B�ߞ�����/��?��#� ��4�D�7T�̉j�&8?��ψ,X�%"��+-$��#g߂��O�(�f��$�Tu���W�Xd�OH���'g���X�&K��6 ,�l�&��%�*�b�<�dO�W�8�@t��T �Hr7�`�'7��}��l�;�^�P���y�8
_��M{���dP�h�2�I�Ob�D�O$˓w�J�2�_(p9p`� ����I��лt �eE��F5����(��ɘOY�'��� ���f���A��,�/̘ P�t-�-H/0X3�����OC�'6�%{C��,� I �&cL-q����Ā2HLb�'z���Ø�j��D%\�����[��C�I�9j��1���O�hZ`E:+�B�y�����П̔'���(Bc�"p��8�d"�??��j��;&7�ON���O\�S�'_�l��&ǌ>�ě�,R �([T Z�L� M-K�ʡ��	ܯEiџ9�G_�p���Cėy常
wT!YDEa��
�~�� �*9����g��q�*J9C࢑0���de����O��oZ��HO�"<��dS�)�4ҶN��P^nl"��IX�<�.U-ݒ�2cMÀ*�D���S�	?��d�<Ѡ�ٍy��OLu��^-u��,yF̟�J<9���D�O(�D�O8l��M�>kZ���.�~�`ܑF�ÎFp��t"�i\I�7�Q�+�\ER��LG@�F�ۙt)F��#_�gڐq�ѮY�?�4���E͛R���a��:g�����Ӧ�(O�XPe�X3SHvm�C* �i�p�5�|��'�Z8:�j� ^��-�$���B�<D	��n?���1Ю�[ �ќl;�)P�U8�?�)O|��Ԡ�{}ʟ�˧�?��O� gf`�D��W��4��B��?	�C����VnD��h�rJ�	��2��)һ2*B��e�'-�6�7%��n,���y3��0��?1���� �a&��B����5�dӧ�ֵc�t9�A��p~�/��?1��iJ�#}r�Ou^�+���%h^��%��� �'����5�Bt�F9b��
��$i�O۰5s���~!`�4�@�x�	��Y���'V�$J��Oc��'�rT���'�EAXT,*���]
]ӓ �,K�� (#�"v����d�ݫ	{�p�|�O>9�!LtD$U�̇*��M��`9Xx�"^$�2|0`��>j�t��|RK>A3��AҭR$S(q�8��%[��M#�P��SƁ�O��8&�0��`�|KVͻ�
S�%�h�pQ�f�<� 	�.i|d��`��0x��My�/�S��U���� 7��"���
e���B%
'�^Lp�4�?Q���?�)O1�R,hdd�:�м��&\"`��yda�9J�,\1p�@�i+e�Q���}o�-F"A��?ɐM�Rn.@�$�3 �6)�Q�J��&�{�#;j�Q�ɩ\s(�@BF1 ��mJ�����H��)�OtYo��HO�"<��K�$5�)�5¿׬��'X�<YSᕦJN*y��NV�$	��[�I���D�<�e�"#�O�Ii�搾>�䙖G�G$�E+�����O���O�X7)�Yb}P�CO�.�÷�Q8*/>=�Q�9hw��h5F���F�D]���h��3F��O�ك��.��S���5=&��E�����D�Φ�s)O��	����/dҥ0��r��'a|2B�^�4`PE��	Y��1����?���'rdY���P)�$�R&!�T@`����$�e���֧�ɳ|
��P	2@ڴ䒰lY0� �'V�5*���?IƁ�I>�*�^2 q��K$bܮd5��p���]�	��@�3� ?&�8%����aa5^��)0�Tu����\D�'0�0 C����P$I�Hǅa+$!�'��h��OЛl.�'��� ����m�%�i����`"O����57,D�)[�)˘y[F���h��)g�ybSh�\���#�>�)O0p�柆�d�O,�$�<q�G��_��[&	)/�@9clR.��Qs�|	zt�҈�)z��E����|��ėY|@aP�T�'t��;ň Hl�F�Z�y���o�L�����|"%@�RH�Q���!)���V2A��b�<qA�O����Sj�L>)�FQB���]��@�Ul	��y���Wؼ�� 58�qY�C����}���ɫ<9eǐ['����es��H5Ⓔ.���u�ir��'�BQ�b>XS�C��찐WB˄H�8,��h�'h>`b���J<�I�)O>o�Dx��$Ũ;x�����3��b���8)�ಧZ�Je48Aȗ�DH��B� �i^*�rO_�))�`0&�X�_(F4( �ݟD�4NՑ�@Fx"e�9q�D�C�Ƞ>� uX�����y2���� �U�8E2�����$��G���Ly"�
$ �p7m:��&�*?���dǃkiB k3Dl�'��$�2V�>mQ�)D��b9�k�U=���v.4O�xQT�I)	g�-���B�4�  ���l����b"��W(xR���W�X_(�x`��)!���dT���[5pNBe��� ��m�O�,�Ņ��i��j��k}ұ���|«@?WrRc��>���>3x�r��T<>��@��;?�'JZ���
��6]��$�R�O�����׫U�.!sT�\�s�\�O��e�W�V��4�b*#NJp-���	/v(����O�6}�&����	��F�D���1��	a>��3)��H3�1��ύ�D���!D��:ؘF�$R.LA���;!��y�'n��}��� �����?��3�ط�MC����ʺ�g�'nLD�`�íU���ْS?ưH�y�Eԉ�0=�5�&ȳW (Bd$��h�M̓ab����I�EV���FUd�e� �O%NN�%�x� l�O�c>c�D�P� �gG�c��3������9D�t�Ĩ��|�S�+>*����L�<	f�)�';�$y��1�Z3���]� �	�h'*x�#�im����O�B'Er��@�r�� Vƌe���D6�8�@���c�!@�$�(!4�%�w�'�ʩ�!�'YB�'�4�7K�	�(��0!:(%;d��t�.Ѫ1�Z<~��W�U%�e�]���mEy��E��`i��,J����Q�]&����.
,�4K��ۥt30	��#�|xGy2����?����O�(�ʎ�
��!��e��4(Or��$�"]ׄ8"B�1Dg�T��H7��}e�<a�(O�8M���^=q�j��Suy2@�x��6m�O����|
q�Ő�?���2P`<y6(Ăzd���@D�A�(Yp��oӜ���K�LnP����c$�6]>��|
���;RB&�u��6��x�r���<����6fy:�b��&�ɫ��[�L��-�!����GK&P �	5�����O@�S�E~Z*2SŃ�n{V䊱D]��
$��[#�!s7�K�i^ x�Ɨ8
�F{�')�d^�IP$T~w�`a�L��jޘy���?��~�T�Ӄg���?��?a�/���O����!N��)Y���+���ҡF\F��2-�ENR�*T0'�'�^t��5}�ǻ3h� � jN�WQ��H��K���#���	<��@���s.൲ϟ�qHc�G���ɠA��AC��� ��g*��w �����hG{�=O0My4"�s�h�P�ʘ�; �a��'%񰦯Ćvj��蝊M�����'�#=�'�?�,O���2+�\l�Q�ޚAҐ8�Q��1"!=P���OJ�$�O����n���O2�ӥU�5��'��Q��3��W�g� ��8K��Ah�A@�c�i{ƮN�>�%��I6K�V�£�jOȕ`W暢p�6�#�%�.t��)�'�ВFe �kT��?e<�I;$�I5B����V�l_ �3$��7p�M��(%DŊ��&���O>\0Ѩ��e��(�u��#V^��0"O\!0b��$W������y'�l
4R���ݴ�?�)O�����~���'��P���I�l){�6	�$B,.:�,�O��D�O(ЛUM@�!�^�"D*R�;�������2Y�>�[��َ{�:HWjX����\&RQ�$[b��L���v�Ԁ5�ڠ����=%Rv!�uI�sjf��aX�]�1d`O�j��ܑD@ˑ��s��}��ȟ��|2�mÅ��i�h�	�JhBgD^y��'����oֺR���S��9E����p��Im�F��%��t���`��"#b�'�*��i���'�ӳd���I��Yf�_	@��@I	]�:A@����R�M�J,єkMe��
��ԕE\�Ezo�j���?E)�l�-H%��Af�C �*����u���� Sv�l ��&SZ�� �K6%Z8��C:��y����dc�8}&~D���V.W�X�!?O���7�'q򒟒���S�? ��ZC���A���D^>K>�0��"On�����U�`iȅ��9x���{���ȟ^p��lU:��g��D��� B�O����O���m�#$���O��d�O����?��e�y��8D�V���8��-�� 7\Y��N��uKn�#��
�^�2 "ɟHd�����5ܵ��D6H� c�ϒ9��0�3dѰ���I$$��2"91�����9!M�(0�Ŕv󎂔9�bYPR��o�� `��Y���,����OΣ=��'�0���12�ޱ+b�1 �� A�'2z PBK�9b���E-|�hp���:ޑ��ܟ��'�h�Xa�u�ـn]��H�;�� 6��q��'�"�'��`�]�I��H�'�0�C�DY>����o�j�]A�I�)&�b1C��#x�83@T�6�vH+!�;ʓ:�V�:q�ܸ�D�B��D�I��E��-��Z��*!O�/2
���.ՙ� )�ê&��Y#S�x��?q$+
'�Ȍ��ȣ*��d mW�\����9���O��k�C��H�r�:���Y�Q�"O�À�˾T1 ��2r^��P�ȫڴ�?)O���&_U�4�'Q�����S���<B@1x� K�D���*�2�'k��ͅ<�sqN��dr��yT�G1~�X`�o�"���"֟��m7fŧ*h��P��D�Kv5����.�z�G��<�hYa�Z�n"� j�G��z� ��F��/Pxɛ��dW�Y��'�1��Гh�H;��6k�0I&S�4��I���1��d!jE�� >f ��D_y"��;"��g����1m�9��D�O<�d�O������OJ�َ��4���D0����6�Tꓠy2�'?�	����C14����n̊F�>��DC�)�Ob�Қx�����O��YG�b�f�Qp�Ί ���O�ͺ�'(B�+N���<� !O�uW��ZB�@8i%D��w�ɓ5A��ONȤO�P���>�����J �E�$|����wI"�yb)��/���O� ���h��+iH8�f��OpPECD��Z�a�>���>1��[f��B�C��.�jth�f�?�\񩗩P��?ɲφx��S"G%�?u�3�2~
�@��c@I{���e���<���4}�k#}RMS��ɞ�M�V��0W4p��TC����L�rybϤ��ɷv���+�'0F�t�f��,zy����/���Z��O��`!�>��y�i�:��'ܤpAd�ϩ9��A@�ֻ?/-Pa�KW��P�w|���9��>�z�(�7���hSꋪPOP��J�O�Ek�'YH�j��'��y2��~��l~��� $��I��?�g<�	ǟ�������|zb�3&2�A��?,KFD�{�<Qև^&Y��X���ԼY�}Q-\����џ�������'AB�'�r�'�2Y�s!�b�4 b���3��`G/w����O����O��O��>�����'h�^�+���v�-i�ds�(�D�<���?A(�����O���ss���C쐦q�I��ÅB�X6M�O��\�?Y�'��#UCv�b�!s����P���$O$D@\"2Qވ��E�'\�YE�i��IM�)��a�t�D�����7F̅�ê>D���#X�v ���V!6,^�y �:D���'Gϯ5`��ď�2A�|��R*+D���i�>4��B��q^n`3G�;D�H���
" f)��"�9�~)���?D�p���^@��1b�ݝ'���'�>D��B�g�;#�J�@ę�	L©�A�=��?����?A���?�1@U�"Pٶ ׬9�8A�7�ט��V�'�"�'���'
��'qb�'-��Xd� �mF1V�i�WlY�#�6��O�d�O:�d�O��$�OD���O��B#m�P:�IJ.D0*�I1�5}��l�ݟ�����\��h�	ǟ����8�		J_,qC6�ʱW��q˓vG�I�޴�?Y��?���?)���?���?���^Ȥ�����hk��T�t��i��'3��']R�'j��'a��'btB�)Gb�����O���֡c�"�$�O4�D�OL���O���O��d�OV��m��B2#���0(�Ĥ(��]����	矌��ٟ��I��������I������ ��(��%׈*���p�2�M����?!���?���?����?A��?i���R:�3mEn"�����K�F�'c��'���'��'���'��A
`�F:�e��%]�J�z�|Ӱ���O����Ot���O ���O����O�-za�ɓ?v$��']���p� ʦ��ϟ���۟,��֟���������py߂f��t��~�X	(ס^��M��?����?����?���?����?�S��J^"`k�m��T��8b��E#3�6����wy��S�C�xP�M�7�p����wp��lZ�^c��b�i �DY�>1rk`���&�ª��7��禉���+�i�w�R6��b��B�M��Qԯ��W+�x���O~��q@@@�Ɛ�"!��|:�'8bu۱
�!I���rH�}��I0���+�dN禉b�=��N�? ح�T��.7\��Dˮ�Ĥ ����T}R�g��n��<�*���� b��i�*iYOZ}z6�*�U������$)*���/9?ͧBF�3_wɲ扒W�
 8e$��7@ C�b��n�����D�O��}��D N�03)��o�� ��'Diȩ���Ms��|~" w�����?A�@ e�$K��6<]���	��M���i�X��暟��6�"Y�.����|9GG������ҙ~��[���ԕ'q1�h��r"�j�H��'ѳS
�TzdS� ��4%�<��<���`*h��4�ٓEn���@$��͛�*h���IZ�O��Т4��,LY�A5`����\���� �O����D^�WV������D��e�<bPJ!E��$z���y3����Od���O����O8�2��F�y��D�l��%[�#�J�>\�jʐ5���x�p�P��Of�lZ��M�W�'�b�	EY���m�T��j�����
�M˛'��	w��9wJȮZ��	�?i�;/ovX.��� �㗪Ѭ0.D�(��埴����8����T��A�O�&���^�6�]eg@
k�fmj���?!�s@�����$�����<���N�����p��?X8���#�� M�f�q�b�I(~~6-t���	O<�9��L��TkA/�1ll���V�� �)��V�Xy��'���'!�ƙ%)n�5.G��z�#  L��'���>�M��l�Q~�'���4�~��.9'�}�@i˯@N��0Q�<�O�l��M�x�O;�D*�b�xiOU��HÂ�
����PW@�2��1�Q���*�~Ů;3��'�&��S��Q
B��3JH|�"��':��'r�'�Rl�1x���#S�4+ٴpn B��׭E�I .]4_|Lr�GR�<1��s�V�|�O��GN��G�V�x��TM�h���匍S�V6��劣��^ʦ�̓�Mc�ȗ_z��P��q��I�^��	�1m/��@g=H잹���_]h�be�J�|9
�iW�0<���9A��jM"{�f���K@�<)�H�'*]L�Q��+*� ��ɓ�N��)BD������* �T�UJ�->u�Э�%6�P��2˖�Z����F��Ҹ�:��<w.�<�ã�c�q:�H�)~�&�θ!2������tz��ʰfȸ���дw�D�� ��L��IPBk�
�Y����N@!d��/��8!�M�=0*$�	p�,��q�ċ�r�T�!��%xB<�Х(�:�!���s�\�� L�i �pT"��P����SOV= ��;F�� Q	�y���Y�$���N�uf\��!��D��%��M]+,�x��U&�	T�^� ��\'V�|��VT�Uy���i�f���Jдv�(%��$�H�.�F�Y-ͱ|�𑊧��~0t�Ѓ��1�A+��L�Yq<7��Ox�d�OV=8�+Sg�i>����4P���f�����6�0"'�
by��'��l���'�"�'�"���.�r k��U�h<΍���$Mg2�'����F�<�4����:��G�}�D*�d|�%��d�{c��G�:��<���?	�����2�Y 4C]�&�\-`S��@3�DW�AE�I����ß��'���'ߴ̓$���v�d�w��({��C�O���'12�'��Z�88�?�
��jq4HG&�5���5�Y}y��'�B�'��	X�Ɋ4���4�8dA�#�'V"b8���K#ܴ��?I��?�.O8�S�"[C�ӇY�,%���I�'Uz ��bҒq�H��	��IbyR�'��.���O��ॢݒK�
4`fb� vNH���?	����Ě..��$>����Ã��	���ZgM-	��T��@`�	my�Ge�D�48��(en�U�L�a��>, \1a��'��I#}�4kݴ��I�O���ky�N�M�m���H�PB��S$D�?����?���֘��?��3}�׊X)0�hA���e�jU�?�"�'��x���`�>���O �D��,$��>m��X�$鉒~l\,������I@�����*�9O��Ă!}PĴC��2��saͽ 
n�Ο����\ @�B���<���yҳ��7��
�x����#�a���?a)Ov��®?���O��D�O�U�����(>HX*��w)��5��O����<��'��I̟4�'���B)9h,��ŧ'qF��
�K��n���*�'Fr�'.�t�')rT��Ճ?�z��q�@�IW2qX�#V>��h�O���?�(O����O2��@�9+�o-�*�"�L�-@�*%`R:O���|7��?@��$�O�ʓ��5��O�� �e�'(v lhӌ�w�&a������O���?����?�b�o�Q�Y��P@&�'	�nyۂoџ�I˟h����' ���B'�~j� .�*VkHA�@P1�J�gN:u���?�,O���OJ��� p���� H�%��I��! $c�!�sH�O�D�O ʓ��H%^?!�����SX����H��"L˥)�����'"�'���ư�ybP>���|B��4	?������9��i��c	��L�'��iئ*w� ��OT�������'Ӵ�PQ�L�8Uʀl�1���Ђ�'t2�'zΈ�'-�s�,�|j�g��@�IK'c��T(@Բ�\ɟT]�Mc���?!���
�^�Ԗ'�JP�UdJ*6j��X%�-T���1��'�X�K�'�rX���� �0"gj�{�mB���(�1�s�i���'�b��� �������O*牸����7-�S��(��ה:� ��<1TK@(Q	p�L~���?���`�Ɖ�ԏܾ�Z��d�4e�x���?�S�4���wy"�'z�����P�;� 2�\�\|�]��$�sy��ܤ�y"�'�r�'S��'S�ID�? he�Э�2El�s���bn������%|����Ol��?y���?q�c\�K���$G�f.0�'6q�0�ϓ�?y�@�ܜ���?�,OB[�B�?13P!'7�r1H��[~4j@{2`7���OH�Op���O@tk�2O�"��k[x�jP�W�|��g��<���?�������X%>��E�W5~���p�@�o������_����D�	�����er��	Nyr�U m2��;"_'l�҇� ;�b�'RP�T2G�6��'�?��'��Y�f�,!G^l`'%�i )�O>i���?�d�Ⱥ����t�3���:�H�!�jh9�L	��?1+O�ĂuE��m�O�b�OҚ�ܰ���
�C��h0�.U�zZ���I�t�I�2N1��}�)��f@�	{�Åof��#�P���^"<xQl���	������ē�?���I�l`����B�,:�сth��?C��<�K>E�t�'�n�Q�ș.t|qkS�[�Ŷ����fӄ���Of�$]d�$���	����yC��ʷ��)Y�x !a ��>��	o�I;$H�%?�I���I.+O�
Q$�+�zus��8N�p����PV��ē�?)����Rv��# �#[���R��K|nL *O�|��o%���O��$�Ojʓfw��Q A�j��=҃�>y��Bڍe�'2�'��'"�''����)Z\k�=+%g�<u�Fh�C� ��V���Iܟ�&?m�P����:5�䄰�O�h-����+�Jy2�'~r�|"�'ؾz)Ү]�! �A�H�#��O�.u���$���Е'��K��4�@�m�t�R�"8�Tʱ�ӯS��d�O�O��D�O��2��O2�V2�q���v�$���J�i�^���ן8�I|y�d!
�Z�"���0^,�Q�"�Y]l�P���^����?��+�x������ʕ-B�T3�JPm҈��+��?�*O$�`��黎�O�b�O�x˓DlY�G�A�r�ɒ)�����ş(�	�����]�j�'e�ƅ�F)���agG$NV���U��ش�?���?1��D�'�rn�%��A:N؂A<��`A֠	�bѿF��O>��I-RDP!cJT�E4*9���1R�@;ݴ�?��?��Z��'��'8��*3L1AfMF1ȂX"&L^bҔ|mI�j���EK!�C�����
�b�faKkƮI�
,	���)'ߜ��oT9L�@�2�K�r��,
�L�I������xAed�zP��?t�V�aR
	�+�h��	ǟ�oZ�$Q��|����?A�O���^ł��ѝ�2�{3�D$#����O�&&���)@�"b�R�#�r�� ��<��� �w`�Pǁ�7#G�y�B�μt~��"O���0�§�@��f�ş�n��BO^>�
0Jb�Vb�f�0mĘ8ؼU�a*�:�������<)�LY0���*�s�hd��O�%3�eb�
Pƺܑ�
D3G�.���i,`�X�@ /�g�8��5M�//�~��fɖ	���G��E� ��X��a,�:F�����̉)��x�Iҟ��	ޟ,�Xw��'՛��^�D�1X����d�x<�qO�_]!AD!�wDJ�/�-�x��]w-���4�LF���օ�gBt�����3 T
}����*vO0�ٱA��\�,�J�C����ѓ>�t�N �'ExĢ�$�F6Ma�D�����'���o�=}�>D���/�q1�ۜmI B�	�Q֐c����6��T�
�RӮ�<�²iBS��k@����MC�4b8�[`%ˏL�ԁaȝ'R��r��'g��'�h�X��'!r0�Ph�⋆�xX[C��[��]����?i������Ӊ
G$���T�EkA�E֠�(O���=g�DʗȐyy�3ĕ5z�8�����.G�2L���ޥq`���t����(O6i���'�0�I5$�.$���كG̬�pT�߻/�JC�I�Pb�������)�J�>��	Ԟ{�^�pgNޒlNd�QG��Y�@Bش��z��{�X?)��V���ȤAA�h�F��"A��|(GdȲs�A9�'�2�'T&�����S> �����u�|�$�D)Cm6�H��S��7A`��'���I��y ��d��Ew�DY���LTp�"�N"𤰷ϓ�$PJ���7NZ�,�5`rr�� �F.�O0���'���S	���чF3
@�PsB��57f�T��'wڙ��+K��8ȳ��-F�דF�qO��;Q¢l�q�hY.���4r���"'�i���'�~�'W�2U����?a���M#Ƨ�Z�^���`�ٳ*
["���*�)Xy��b&�l�'���$r캐�ǘ�GK d�d�</m@�ϒB\�B7��==/�����>a�S�a���)�#�
?������'��	����˟ $��Q�MϹN 25��%�:��'�'D�,�5��"�D���Cٷ�&Ĺ2�1�3�HO����92�-�':1��٪<��pS��#�?y��M^�$����?1���?�����D�O����!h���:J?����!���'!e����O�#ZrD`��K��u����A�?�0eD�_ ��w"M�}pL\!�ǖ'2%P��$��]H����y�;2��� P�:��?s���CF��[>(( (5�V7휵={RM+�O��)Uؑf�49�"ĉ`�0�"O�T!1mR�~��'�U�H�Bm"��	��M�J>�A�ܬ8:��i�$���f�Hث��ر$%�z��O"���O�̚��ON�$~>��`��O��S�? ��q��F,������;[�YY��'� �XL<	w���"!����M0]j�:�n�i؞�)F �O���2�DX�GĜ[�v�Zck�8��ȓU>0=���&g��Kԟbe�a�ȓ ]H�a�c�3[�쁲Aj� ?�l j+�I�9$���ڴ�?y����Ë��p����bIb����+j�����O.�$�O���a �hɬ]��J��bi��*V��l��~���v(�3q� �bwnτ-��tCbe4��:�XXa֍��aɗ�fZ${���f��D��7�����(��(�����P��'�r��.Q?�8V�S�R��L`��ߖ�N�t .D��"Cƿ3�Z��T�@�]����ʭ��E{�Og��X�.g�)[T��g��l���l���a�i�2�'|�O�&�r�'���'r��
��14�dEU(d*�� �X�c ˝q3�����k��xь�$Z�b>	�wA�͐���G:y�Ъ�%!'څ���׌>Nz"Rc�8���cq��.j7�(�y'G�1X��k#�Y���;p���&r<�D�x�I��H���t�M2f��lb(�ȃ��:e�C�I/h�z}"U��
$x����]�t���'N��6��|B�O��KW,��,��EٚsG�1�@����A8S���	ʟ�I��t�^wa"���3vD�鲢�!8W��x�Ȟ�v$4G�	?J����i�Mb^wwF	D�
<HKQ���Ԡ S5�TS����pK����2��Qsi���ҫH6���Q��%��ɴ[AD��b�7\ά�!*�)|,7͈�|_��#�Oj�;vJ-Ĩ�qkyA�l�u�'�I)I2ثfg�:�\�PS��&~<�<��i��'�(D�F
p�27-�/u�F���D3}�\$�p��';Bu��֟t�I7������̧^��DpK�����M�+��h3�Ϻ{M�|b�S:	;i	��ӗ 38|�$�#ʓlM��c���!:�հp��t�	b`�4 _ �W�ՋG=:�9T.�(���=ʓ#4ܝ���~�,��\G}Aa������b�y�RXQgB?C�̀a^�èO&#*g���!����g�ѿ`�-�e�ϝr9�6�<�$R��^mZ��p�IN�T��2��1��3_�L9jPh�H��I	s�'���'�@��� �0�r4L+_ކ��3�E�x��x`���(�����)+�D��W�u#f��R���R*��v9���*��Tb�85�X���wD_�_!�Y��U9W�Ba�@y�S\�%������(�"�,Q�[�h�x��יR(��:"O E��`� �=`@
���)q�O:�=�'x�qO��ҥgϒO�qʵ��Y��9��m��,R�t�ܴ�?1���?ͧ_ހ$���?q���M#�	�S��v��F&����&A:���!I�EhDS�D_H+�.ҿd�1����;i<�3��C�[p*H/�8p����%�^:#G��a��D��Bd,�=^t<
 �o�ʧ��nF�C���T��{"�1���_8f ������'�t̀��������H��9ӌ��r��`��ps��'0%ە��?-;:%��L��S#ȃM�l�I��HO�)�O@7M�	^�E�c@ZOb�H�I�E�T<���!D�=[�Ñʟ���џ��ɜ�u�'j�;`����9\�
�Ci�2פ�o�np���dӢp{�5ӕ�ڧG��rs7��k�)
�R���@�� �����^4�I
�B��� �?���'��uHAEZ�fgtx�l���Yb	�'����Ԭ)n|}�6 �~1��ʍ���Q�/:�@`�i��V�>P0H�6��q�x��fW+% �d�O�� 'qd`�D�Of��F���$�>yWg0C�v�h�D��'v(����U؞4�5B"�� "1p4�ɽh���� Ǜ9@a{b�U5�?��O���jJ�,8�aǨ�$O缜�T"O�-�쓙���2�l���l�`#"O~M�0�۹"v���°z&
�����'
�}�����O��'h�R������=i6�N�O<Ċ��*�?���?y�$N�:�.0� L�"����g��|k�@+���uυ�H�t�g�b�dap��2��'_ڬ��l^�1��i�KĖh�^�"և�9��}�S,���l[�*��)�)��b�tjr��O��F���!n��������1�X#�y���%c2���C�T�Q��fdצ�~��i>iq�{R��$�&���P��f�M��L%S�� ��=�	ğ��i>��c��������o�:[��ͱ0i̕~�>�3dKד%�������'��3�E�>H��J-k}8���)*@�0�C�QDt��坡oX���LR�����Pm��d�z�z\����>0y�	���:�>�L�b���FK�W�� �q
=8�JE���pD��H�n�^�����;D?\D�=���i>��'����p�����öt�,���h�OlQ!�� A_��d�Ob���O�ٯ;�?I���Q�Bi%���ᣪ�/9&թK��T����	̊���\�Z�d��4b\$B �� ����9BY��9�a����N��xh��]�.��0���&N��^� pT	���P�q��sn[S�.�(��݄�M�q"����C�-��� ��b���@/�� �����E}2�A�-�.9��̡19b��D�	��(Obm�C�I��2�4�M��k^����kͺq2�ɛm���'�'�%���',�i]R�Q���_�>�0�A_�hqe�!&\.g��Y�ɏ.cL>m"u@ݝ)Y���Y.f���&[)��+���^��:���+p�4�!'� ����mQ54�*s��DB1G������E`�$��ҁ�S��-Q1j9D�t��P,C��[d�RyzdcN"��ȟ�8��ɘZ��h��LH<(���>�MK>�߬w����'`�Z>a7�ׇ0~�K* �Ap���Q\\�rQ�I��P���<���ۙ F�nZ#�4H��eQ��f]�XwS~�EfrzZ-x@NV"<��}��B�7tV�� ڄi'i	&#c�"�aC��+7���GZ�*��w�t�F6�'�0�#Q?�i�o��zB��{�d�Q�"@��.$D��y6$m���	0n�}���%��pG{�O�8���#[ �:�x�MÆzw��c��>,�Τ
��i�R�'I�O�|�A�'���'.����%7�R��E�}NZ�*�A�J��]r�)Ik��6��b/:��@��<|��|��?���rW��� ,�����C&"ӆ	�2wz�U� E�P�`�3��߰y�$ s�g����U`�|�t?�����3(�T�9���B�T��Gޟ��J>���>���&"�TIq!��T*�i��'�^�<���;��Р���5��(���JY���O��Fz�O���9C��x���G�%��[�x����d���3�GT(�?!��?��M�.�O\�4��˶��a�R4*�MV> ��3�B�7[7�z��Ⱥr��9r�M
"�u7�I{�Z�� *�	(���Ì������J�?�J,9�VoL���
v�G}�L�}f��l��M�Fŀ7���MK��ퟨ���$��u�C[����!26I�ȓ I>�"ԫ��aoޙi&����lEy'uӐ�ON-���	mڃ:�D���OK������X���=���?)��x:� ��?!�O�6����dϭT�<X۵��-�H!�˒i�a{Rd2��qVv\�p���q����'Hf���I�|��$Fl?i4��7y�)����:3��x8��a�<a�)F|%�8J��	�lŸ�c i�_�<���B�D�B��,}Ba�3̆�Jߒc�t��2�M���?q*���r�'Պ��`	�)�+:(D���/\~D�$�OB����g�R���a�E�h��k^�O��s�)��kF��ud�����5m�� s�윧(SRc�$B$��c��ݨ3��V��s�۪D�J�0&�O�2\���I�R�a�-ޅ��m�h�t�|�ɉ�����0��t�ԼZ���r�ՀP�!�S�4o�����T�J�u���Q��d4��|2��$Ɗn�`�dFX<5�`d��]�pSb��偈��M���?A��|"��1�?����?�ٴ\�$���϶JF$�y1�%��(��HR@��d��i�e��]�E�:�k�h;���y���< �A,A&C���
ğ���qPF��,�R�2ĨX 
ʛg�������Cmޑʶ�B�,�
�2@��,_��\�" ��?���|R� �g}�+-�~�ET�;�nH0�@���yR���3�J���!�";b��a�,����ǟ츌�4���X;��ħ�]���E-�.`X�)���'er,+dNϏ]���'[R�'��]�����A�@�,0R�鉀-�0���p��_��b��Q�>��-a�J�9=�n��Y�
� �bH.d�erY6^���`gbv�<Z�� I��V2iw�<���Hպ���*>'��$�RB��~�B'�� f�"DoN($f�(���?i���?�*O
�$'�G�:����'9�P�c�`$g�~bY��hD��"�b�/�Ʊ�e%H�UQ� A�4�?.O~�#��H�n�>vh��L
��K��J�8�Dϟ���ϟ�G�͟��I�|
槟�p0\����1;z4Y�̝�H��82KC�4��ǣ��6��7'V��<I3C�ct%�ġ�.ô�R�p��r���@#�$pt���� wk�;G�V�<IDo�ן�{�'��d�W��r7�:����y��ғ�N�8��bʓ4W2�D}2�����cщ��eՒ�jj��RȈײi-�'�Z|�q�e�N���O:˧&YX�Em��LbL�sGۤ)�L=c0C)�?���?b.�(43T�C��$�M��-�,s5�!s�GKe��.د~��rQ"�.M�&tp��$�O҈�A�Z̺�CwL�|�����9\T41u-�7�J1h���ٞ�x[�J4i�hV�H��'�B4I��e�Q?Y9�ϩB���B�902��5D�`�b� 59(iI������J����E{�Ov�➴S�k8T�&���~A�4q8r�#��^ϛ�'�����DAW2t��'���i�r ��V!a����v �>H�� �a��h>���
m'y���
������6���yg���XA����dP�w�!�S��9
��FC�� �U1Aҋ�j�~�1�� 2(�h]�*s�q�#�J��T&�󟰺J>!�>Q3�,'�1�s�X3d�.Q�` o�<)��y ���sK*V��m[�CB�$�O��Dz�OO���u�(���9C�P9d'�.7����{Av�b1L��?i���?1�H���O���wg�- �b.t�U��)v�@vU�&�E;�V�=��	c-ț�u��ɑO��A�?��H�0��k�E�|�-9����MQ0F±Vl�)����5��E�ߴc�9FL�k �IL�<���݀LE���a�>J���(��2���'q0���AE�l0�$*�hOl�bq��*J�~�U�ls(΁w~x���d�G�@�'ʓ~����|­X�0�t7�l���@ChO#`����I�)�5 �ʟ�����p91M�����	�|�a����Y��O��h�D<gXj��TJ\�5�� 	�'ؔ9j���	AF��W���|X�lה��� �l�2u�zA�ʁ�u�����' =����r?�Ԏ�7>5�����Ր8�Y`�jOV�<�B�X#6�jƂNצ1 ��Uv�<ye씬$�y�����<�w��W9�b��RC���M{��?I/�
�@׀M�i��9 �� o�Q@V?	��D�OP�d�2X����%��Pb�S�d��.��'O�-=Z��	V0;�n`��$Ơ-|r� � �h��eã�������HB��juɞi�d�ZM�I������b�Ś)6�L���D��4��"O�l��hV�po�H���
�ʝ1a�'���(Z����~���2OR�h]� ��y��L9٤?R��':�O���3�'��'��6"؝av�P��;O��Q#�lN&!OJ݉e��%��`�G,��M��ҟ�b>�Kܦ���NB:[]B7B���xهk�{��$wf�=BJ,�o�>�H�����*�S��݊Ma�l)"��6U2���X�'	:"}�'�<�yCJ�y���I�
Ŭ��P�	�'�X|�"g<$������c����{"�>�S��Y�:	� K��:����] v'| "��Y�PA��ˋ��?����?��1���O���w��c�a�37n\)*%Zr1j���Au��!aeȈdĂX�V&׸�uG���q���ʁQ��43��Y6��X��=Y`� f��(yl���Q�f�٨��XX�'tX��}�� �X�O`I�شH���ɒ�p>i���:n��u��㏳8�K"W@ B�	8 �MQ�n�- $���'�i
�<i���ªYp�o�ަMK�oFoV$!���:�H�����4�?	��?1$�ߺ�?�����C�!�?ѫObax%�ӾQt��1�!C�F��ݩ��'!��)N<1��2&�R�x�*�$��D��"�q؞��$�O*����9���6���V�B�	Y�Ć��`���]�l�F`��Ϙk?j��A�����D�jC�a��3d��&%���h_,�A�4�?y����)V�6=��S�퍀7B�W ���� ����O��$�O�@�soLj"y³K��T>��;a�2���J̦o����@��>>%
i�>i�h�p�"���aW+�>Ɂw�
w���Q�1w��5 �"3�	�}r��C�`�4�?O|z!	(��ظ�썴���W-����O���<!2�M)m��x��/ 25#BВ0gDG����{�h��z�iM�^�u��N1��i�sh�ᦁ���d�i>�W%S؟(��ޟ�nZ�������� �B% ��U]����T��,�CXg�n�Xf'� �L]��!dމk6`��Yy�a�b'ȟ
� U�e���T�Y��Z@�ٳ
P�h�$ʥ�vܧX�����D����^	TA�U�*j��h�����i��>������e�'[IB���,Ϗ2T���@��( 3l��S��W �PT���!�I>�HO�>A���@�@�Q�M� B�|P!!P?��lZ9|"��p��П���ß��	�u��'+��1!���F�sV$��G�W�A�NnZ�E�1u,&�*Ec3HҴ�0<��B�iZūej��TBIS�M��A�O��5%2A����0b��aI\� v*�NP�o�^@>���kX���C��!o*�j$�Ń9K�,��"O�\��ծ��=㠬F<DB�1�	��'X>���fx�86-�����kM�`t�w�ɔ���I�� �I�D͒`��ޟ�ͧn��H�) �J��� e[RT��e�d��4��h�a{�(��E� �AK���^|�dH]JJ�5KR�1ϰ<�cj��t��yB�R��?�u�O�%��ԹUj� ���#;n�"OhĒQ�S�W,���%�L���f"O:���*G#G�p�# ���*|^�7���McL>�JK����O\"ԫ�-�*^y���3��E(#Z��B�'S���(D]p��B*�"z4(��Cj�D��/���&"Q@��G�K ^��իM�}��O�)0��wU؜)g�ے%��yň[/U$�r��O����.� ˒8p�/�7`l�>���ߟ��I��MC����g�? r� �BF&/�(Z�e�	)h��9$GX��?E�,O��iG-�,8?|�2�cG�8��Oh�=�'%E���q���\��yl2�X�������t�Dpp�'-b�����Z�'�´i�0��/�_�x�1����i!5��O�b�tX��hO�	J�	�:��sS�Q/pt�� �y�'R�"}�'���S��5���a�(����8���O8Y'����Y�0�S/�[,ژ��$,܋Gb9D�,0��A(�0��Ś�Z��P*�g6��HO�Ox*��ģ5�l� E���[`�)���O�ٛ��C����O��D�OF����?����I���Y�p��!�0<�@���(ҙ�h�p#�Iʜ�`�!����1-V�dq��d�+�D���0B���)Q�(,8��ťt{ڀ�a��I�R���09��@��7^,u�@�M4 |`r�� �toZ�C����OD8�hK��
��0T�V�e�`���;�Oh���)1��]:S��;�GyB�uӞ�O�ųpA��o����c�9�F�P��+<&a#��?�tx����?��O��m�BgZ3o��Zp	S�M1���A�.<!V��G?FabC�	xF��7OH�'�.4Ud��WO��P1%[�qg�!���8���hR�^Gl�Q�@�_m���0�s�'�"0��	F�$
��Tz����[ތh�E0=�!�DI|���@��H�&��1
U�L�Q��E�떌t����1K�%���cQ!1��4o�T���.ya�4�?y���^�Y���g�)�D�X�n�(I��:S��O�D�O֐�'�R���D�=�X%Y���1~��C��p�U��#'*�qӤ���庤c6�+��(�P��Q�B��^�ĭ[=4+Ȕ���2;���C�KZa��	�1&,�	�����'d�4����ȟ�D���Z �p�Y���*R�!�"O�Y�s@�zP�K��[�
,
����'�➈��T�zņ�e�'O$|p���OL�IoܓӈO�[�
T�e��h0���(#l��"O�|��k_?Cx�i����H|�v��N���KtG!�r1	�h4jx��?9��	'�,�`&���S]�=bQ�G^�<Q����~)ʌ����#��-�aIX�<1V�ɧU�P4c��?�B\0�D�q�<�@F�32�|�
m��}�`$ ��s�<�������� MD*2ԐVKJj�<	&쇲|]f��*.3�>Qk!if�<y��Ҙ[��K4��g�3a�$���Θ�w���t� �&�?�E�ȓ؀�@w�žrM��PiV�1�ȓkD���ǐ7YI�\J'�2�J��ȓ�0�P�Ț�:��|���%�Ry��x�����!k��(ZT�T���H��r�<��,*	[�����^�d��hXx��B�ѧ:�"	�c̒�'����ȓ$f$�B��Zuz8Q���.5J���.�HJ��Ư5�&� ��_�A�b���Y�MK��r�zQ(���+;*u�ȓo�*���-G❡עL�E8v$�ȓt�vQ�4��-���;1�۴�}�ȓ
m��U�8:�];B�ºk��m�ȓ	�(����Z�+���&d��`0<��ȓ* ldj�]:Ce�i�R�N#F��a��:���v�د����F�!G���ȓ�:��5E�n���Ɣ�y�<$�ȓm��c�L"?�D,�fjV�@�j�ȓf�.%x�-Y�LdeS��50�F�ȓ~��	��Ǣ!�jy�T���X��u��8d�*�d�{�Ѝw��/~�t,��Eǎ I��⭪�eP"!^���ȓa^���b!�$�T:�	>M�ȓy�PZSF	,���`LԆ~GpH�ȓ8��=8�O�_�PY�3O��s"��ȓr�:8�6aX�b��M���ϼZ�6��	V�����E6{�q�a�?$���,��)Q���-�|􈆂p����*�d#v�M	a��8�]�B����S�? �u�S�^�C��<ڰ��"O�Đ�g��n�ӧ��O��2F"O�ٱ�C�F^*0����.%Jh���"Op�����4=��z�&2n }1�"O���"	�u�� ��P�di�|@�"OV�!Ԥ��/�(��o�G�KW"O*�{�-v�t�!�s�:�Q�"O�U9Aݿv�	Y����n��ɩ!"O�Ĩ�c�0o��my�ɠBFZ�a"O��(�@ө)Ʀ��we�C6N3�"OnT9�a���	9��Z�x(X�0'�'�R�8A^�+�6��ы�6eB�!Vh�)$w8x([(��B�I2c�&����ʹWz^h`�ǟ?ZGr�<�EDG3a�.�Ƞ͵UyX`$?�w�O�"�C)�ls>� v.D��3��ִDkzP�"�W�Va�䌿�`U{�f� v/�8KU�E�MG��'|x�R&,I���b�^�<Ɗ���'`X��&�n�6h��&N�T@jB&�;jJ��V�C 5Vtڤ�ť�F}⡗�{5�mÑ��%�����H���=Ƀ���]��$!���{�4�I$i��p+�*#�߱�r`��`@�����'>�řG�U ?*�T ת�:7�x���}���]���P��S
��*h���RZJܱ���	8����ؑ�0ą�TL��"�}�Tux��݁Jt�0� &| %���QD�9p�D�V�O��	�Z#�"�+ڏy���8���	jA�B�	�xu��W. fȂ�Z��!Z��7g_�z�t4v��*R�� ʥ	m��ɏ���H���芃T̉��&�0/Xa{
�^�0i�ʿ\4�(��	�96���Ֆx$mU��D$Ȕ:	2���:6(m3�d�"/�x8Is��-7�O�HSe
�y��V��UBX��Դ!�V>튶!��M��m˷��1-C΄Ce D���B�6'���3bW7�f�� �8*zM+��:.hI[J�M�����)���+��
�"Èx32b͗8�h�2Gl�l�<I��مn�dQ�Zy:Z��	 ����X&�[�[��PB0�D����P��Q�f�6�	�.%:�@�5[��h%a_9
$���I
W���Ӡ���4�H���00�b �c�"XI�C�6�r���	�+6%��ITe�1�B�*N~�m�󍉎y�z"<�o���P+�%G�S���V���(����Ѿ��6ep`��^[s�e���Pl��O� �`�$��+�,=0�o��A@����N�p�Z���� �Z|����w<"��jߒnAN�$�*9��Y�'R�QKu�I{<�`$�/(���e�7P����׃AC�����3��	L�F�`�X.M&xzŢت[��,2�	9�O|5i��0JЈ<C�''�"x�e �y��S��ѷSt�Lj�MÕ]@���Ɍq�� %O
�9�|�0�'_�p1;��4����ڗ%r1B$roҬ{��1��ɩxS��"�JΪLH�j GF�����"Oxu�����[���u(�h�vux�i��	���9;��-�:Ċ�A� !�b?�Xf���D�O�r"(eҫ�(xC䉌z���Z�{RH��C��C���Q��#)t�����<5�C���~�3m�-/�I�/�$��C�U�ʀуi]�$:u듪�#H>a|�)�W�
u�QeC����$ɐ+2� b��%5���I���K��J3l�!"���|UpT�HԚ`��u��Y&� ��C�Ҽͤ5���6�HO�I`�҈ZD�ɰɟ`��%"ڇv�:���j��h������$���'�?�&�ɀb��=`��1����,��幁�ߠw���hB�t6-V8>0��CD�S�F��j��[�9Tv����>@�1�k,Ũd锁c�U�x)����=FV��'�l�c1�?F�%�ȟ���4��516�D�o�<,u����L�PlsãΧ>�jؑ���x�8�~*ձ7CN��.���̧M-y�#Ƃ 6�
4b�i���3��P&>g* jӓD_��$��0���a��x�� ��G�"�a$�Ͳ;p�Q �� �hAԯ��G��4�!CF#r4�A@��<i�O�p��flY*J-���T8�0���d�.Ѐ5{��(a�����܁!���b�M[�#� ���/�I����[���*R��3<"��r��6xI����"��|n��U�ܨؔ'��x�g�^�'"������-ɧG�P�$	i�^R���X9H��є�4�i�Dt��F䜻y���b�(�r�Y�lGġ��(ݯ0��Icg\?#=A%���]��I�C��;���C��R?"��)X�<�\P����:e��a$>��P��4w�>U�0��6�<Rp'Έ`�` ��ǁ�o�Za�Q��rꄄ�I#ݲ�)�
�}@Hi��a�N�R�M���ՈG�E�V<Y&��,Gݰ�1��~JP)`�Eӟ�j��[��4�%��H���N)fn���
�9�	�-ݸV�Ā�1�C����G�4CF�!k*;��|�� 6�|��V�I�&�v!	�ǕNҏǙj����}nڣ
{ΰ3�	�0�@��P	�r�OD��p퐈�f�`͸u�z=Ӏ/����Yw�(�)� ���4�\��ȓ%�$G�(q�d�Ks�T˕+�=ZJ�h"t���DO���I.�d�i�e>$��j)�9/st���WcP��;B*Q) � ��"��.�`�q��?&��r2Is���a��#]i�1��
/r�2��h�31���!f�"���:w�'�f�y���`n
PW��)�\�0�j�P��RV�7uN��Ђ�Ԍ7�:�Q5n!`nD3�K�-�J�PS�C�T�|����;�TA����CpDC�+,Od��&��2���v�[� k'�߃v��H0�hS�dQ���r���,�E�&y0A�'@��.� s��P�S�jM �$�
q���_7��� �e�vb�H�&٭��}��,�!1]���S�^1k�0�.M!o�(�K�=g�-�rM������lLa�e�e$ޒ.�<yqa�[���X�YITh)�'D�7M\���cWo�:�R E�TJ�	���q���#��W�TY�p�	�Wvb�C��?�DP���O�	����s��r��<k�E�1�.���'��`ކ���
Q��=9��10߾�+�lݲN�,ܸv)%���k-Z8g���d�B�jŴ�r��޼7��X���TcZ0h������6k��}�E�%x����l]�B8�I*������y�OZ1sF��Iͼz�d�K�z�th�եO�6�>D�'��Y����ʆ�^U��Z#�Ä}w����눓�zt��E�.2�$x����9\��8ّ!]*8L��e�$&�>a��Đ�<�R��+[zQR��Ҥ>A%�a���-&p��֧#�,E�s�Q0�Y����N���S��9;�R��R�ɖ}�q�d��9���3�T�-ڀX��M�6Hr��Dx2a������h�Xѡ��ݪ�$�a":\�І�_ ĥځ��)�'�H�k��c���a��o���R�6U����g��](M�v�O/pHeG~�׿�r���I�D9��Y���!jx�rd�A"E8��`�t-th;��������u��{����H��@�f�F��z�Bg#ȷj�b	N;Æ�Ey���t��C	5o�t(-��$�ÌY�d�J��R�>�Ƒ��œ�h���#�ĘE�(M��)��h_0���OF�	D�9�ح�&��l���[�
�C�2y�W�F�}=���C�0^��#��C�{vd,�Wc�;Ϙ9��!N�t  �ڧ'�z2�ဳ��6�Y�N \����n�=q���*�kǬ2 :������?'L�/6�`�r���aF̱T�T�t���r��dV���i�r�G7l�zb"h�x��э.�t`�'���MS$�i�xd�'�'ڰ�yPjщ��1҅�ǶSg�����+$��ì�H��Y��X<Q���!ba�'s�MiaH�8��,R4F�<���.pĄ�v ո-�&Moڒe��	���Z7�X�l4�Af�+?	�Ί0O�f���+Xgx�Hgn\�[9n!�"&�E^hݰ1E��Q���2An�;"�h��WW�)dM%Q[q��A������ґE��xJQ�;l\�H����ꊣ	q$���a����}r�hYLr�Wa�"�`jA��N��]	q�G{�MYrn�%kR�$�f ч�XԦ%�d�ͫ>�����c��o���	E�28��ڂBC�#�<��x�ˋ	bh�`֢ǫvzJ�Dxb��l�B�S��w��!�bH�TO�E�F�U<3Hl�QP�]Q,�y�d�j�T�����Iu�	�E�7-�l�c��S�f8xS��M L����kgI�B���
�#=���ͣ5�F����-�� ��T��ۢ�ݼ_���#�ˀ���UȀ;.���k�^�:�� ��J�T� ��{���3�qQ��5S�[�h���}���Y�2� �ͿmnB(X�P��& Y�6�0��@�t���	�"�H��N0#�y$�j�@�� ;J<9�A�/�}h�DC�"����2)^Җ��PǈqM�|H��ϙ,��q��	z�$i��wI���r鞘՘�� 'HuG�PG�*�����M��j$��`��q���\�l���Z�<F��&
�6�e��?N��Fx�C�8A&��� �X�2	�G&<ܕ#$��I�!���PuJpa"#�G)���`$��;=i���"9؝�.õw1L��F�$!�ˑ'*�$h�# �zh1���$�!0�) �lV�H[�}�����`��80�n�6Q��J/y�c&��E&T�V�5̪���A�e��P�Ci� u�0�ʯ��5P7����ʌ%���:���8<�1O����Z�9��d{��_����k�*��.�,-�Dը��1i�.�ѕ,����4q�K+zɬ�&+�_�,�l�c�����LZ�<������,A���{���P1Aȹ��͗ ���%��.�9�$]8]��PY"	.[$4�¡�����Z&4���jP0Et,�0P������2%��1*�E͸#�9OT<�!��"�	Dl�|�<9�/9F���QD�T��9��Z	C�΍+��X�BK �5�]���8��\�C���9�$��<1� Zȼ�@�8�%���-}��Hb��t>���0C��FxB�ۃY�hM�����`"⇻Iv�b���'K�Rp�e&v����I�� ')�1�j�3��d��`c�@*GX 5��N�8!�`�2�6�ɰ:'�D��
��0��:��P"HY�b>a�7��=M2uxRmN0h�tH��4?��dd�x5�@�B�O�.�G�����w�$�qT��7%�:� iN;�d#G*��B��a{c� �A��3?Id�ƶr��U�(Qܩ����B�|HSA���<�R]�<S ��|�<��
����˽{��`���	(ҢxI�O�3{Į��J7^o����,ȸ�(�@�xl���Z#X�.�� ̚'�ƨAT,��(Ovl��`��[� ��p��&
�=����\�%
f���U��(���	r7|�+ُ�XA���~�0*���^pq"��U"͒c`0��I�� (�h�dXDk���ߛ &h1J"gG�0#8����9w�AbNh@q�ŵmt��c3�� >�6�t��:�&�"��E<L'��K��M���� D��'���(���9'P�y3H޶X\:�X1(܏0���l��`����xR�$[��}� �߰.y̤s5�ʍ�y«\'@����,\Oh�c�	�M���c��b���2��̘@�T��Zx��1��I�~�Y �D���E���0LO.  D��J���滛����V����D��{�0���'���(U���_
8��2I�B�F��'u�P��S�t�V�a���+?d ��'���;��J�r���C�:.�@����� h���=��H�R�� r�|��B"Ov�y�P2}t��(��|�<r"OT���
�0v=�d��;g�z42E"OH���숧f�U��Dj4� e"O��y�柣jZ�����Z�9|�]p$"O�MQ�U;0�=
�A��UȎ�p"OZ���Ka3Z���@a��a��"O$�H����I�ȁ{����"O��Q��WXtyW���"�f�s�"Oxʄ+W�&d�TƏ_n��"ONd�BH�/Y|)I�@?6H�d�%"O�=�a�9�<�`�H�W*����"O�`p���*z��{�,W����"O��YԦ*��bV��mr�Q"O%X�C^5+$f� �J�3].��%"Ot��L9t���V~��"OL�:�f(r�ـN��)0�"O �Р��3+SN��ҩ7E�rq��"O`�`���E��y*��D�}�d�9Q"OP���N�_�r���������"O*�)�E��qt��@��g�R�w"On��f �09>��Ĝ�2��ـ "O����
C�Z:)���W`�}J�"O-�l�h���LE�b�t��"O؄P�L�
�L�����pP��"OΈ[b��]��U�4#�[;ސ��"O6�䀅<��@3�U�J�v@34"O�l㦆�8��1�e��-j�3"O<��,��M#Ġ���Y\��J"O�]S� ;=�x�٧2\��HW"O,�@k�ka�@J��#5:8Z@"O|�L�-M���ЪZZ;v��������@���Y�E�V:.b�?!��J����1@�*FnΌ�b���yr-/�����B�Qr��؆ޜ�yB�ƅF*� ��)Hv�8iV���y¤D�	���U w���p� ���y���)�B7䕭Y���W�G�!���pc�����ȵ<���xV*�>�!��Żv-Xݓ��TJ�,����1�!�$�_�����NC*f$��C'x_!�$�Қ���� ��Ņ�4m{!��ΌV��t ��Ѝ^��GdڒP\!�Г��US@EE"c}�Xc��K�J�!�D�� �q%DG[s�\tX&:�!�$ձh���c&#_Bj�5q��;ij!򄖺K.�i��C�`S�X�dAG3V!�d�*�N���B�E�r �a��f!�D֜}�&����k���%Ɠ�!�D�"������BHP�G1W�!�d�?n��댚��Ed2~y!�$�2G�*D`2�!:���2 bݫ>�!�dY$W���Xr�T.M�ލ����_V!�dL�)*&%`A�A�'�fT㦀	�O�!�<P���v���v�����@-G�!򄔬d���F���Lb�䊑D��>�!�d� I�E�dCR �Ĕ9x!�Z����J���"wCY���A�%a!�$�h+̴I�ď���8�+׳U|!�ʡwuD��@gJ�e�܀1k�0y!�DՁE��Ԩc�ГO'�<���Ԭ6?!�$��^F��JRLX#?&�|4M�-9!�!�z�)u��!q������0-!��59�iq��X�I�q&�7!�	�p�
�񴊌�4Ab��F�$E�!�� ���1 	�?�u
 ċ�BDH	Z#"O<��#�:qQ�8�B��-��+�"OH���œ���x��U�P_�#�'$�:���+͘'H��I(�'b�,y�o�/-����'��Ea���	�օ�W��\��  ,O&MY�O�Gpr�$��|ڧ��$
�<�T�*��Q���[�<����2f�e�T����g���ēg�04�6��gܓڪ���W�p#V�
�Æ�k2�9����FZ��K�(C���kg�D S�ƍ��l��dϰ�0�6����4+�!B.����iS�2��}D�8��"������;�u���w��+��/-�*)&W
�yRG�G���2<>�N��,Or�j��/pHA8�CC\�����^�nT�Vf��m�p"%c "gA C�	�R��x��0#O��� R�k��(!
�w.�1��O
]ᤗ���^'1�I�(y�
Rl�*��8te��B�I�h��h�vO	X�@Iа*
�����`'��.w��!�$�MC3�������N����y2��q^�u�"h�_.��Y����0<�4K��p��ߪ\'�ɛDn���a���0mPKbj
�E�N�1D�P9f���d&��[ϓX7�U��f۲m��UPh�9n���'K� hSIP�Yfp��&ƭ%�`���O�^�컶�K�r3�U�S�K�Ć�B �ߞ��x�A(j�t�����cД1�&矢	~��Fױi�DzR��(JT��G��kAM�7)^}�fIɸb���æ�V��lkEE�s�D|���T�C{L�%������?�� �xf���B+ω��,Zz�d��>�@J�gϓT�NXi4N��H��B
|���0r�Z�1,Dp3�p��U�ƅ3���
��0\I*�N�~�\�2`�@��č��B�ax��z�,j5K,T�؁�b�?�~�lA��`�0��P[� 	Ĉ�"�hO&l�����{^�`��/��l���h�6�!��"N1rd
e�0�v�E$�(�p-�+W�֞�?ٕo�\#<9ͻJ���g��	Z ��F�� o.���ɻK�*�@7�l?p��DM�Vщ�G�~�����'�PX~�8Ӂ��s���A7?y⚰?9����²���0G�J�'�����a�*-kD�N/3D��z�>Bf��d ��tH�e^�] RU�'lF=���_�D��T�*%O���C&�.3��0HQ�.!��_���t ��
�q�s��=�Z�#�I�P�*<�ae���xẃ�`���A�2�4W�ݑ��i���X��r!K1��[U ̱�����.lQZ��=��5j"�	+�&U0�˗�A� p��'��Ӡ��~��� 	O�dA�ƅ�>.���<��O���N[����pE�?���U��p6%�,tİ9WNްa!�(�e5�'�R��FO�3e�ʞ��V�}ӜՁTn�(X�|�������p�iʌ#��C����	�\�"9���$אU�xqDkQ�(n��3����ě�Es���a]�d�c؊��'C���q{�	(��I�Dd�t蒅B�;�py�/��R��~r��=��0b��hP�����+��`�w�A.cf�x�K����4^�i�N;C���cđx���!��	z1j�{~xW(8J�Ր�%!`��=��'�F��g��bOٔZ�b\� \b?�"B�/X����DR'I	�=�/�k�'�����Iȏ�$t��h�#xp¸�^w>��C�d\���ȁՁT�Kڕ[t�i薍��(�=y0:�hu!S�2�q��I�W����5��i������ ���i�TM�$F4>���s�ȋ����k�N�P0�	�@ �I�F���a���r����<��)hQ��,�&pS��Y�G��9�w ���?�c2?��Oj�����d;���O�$+tȬ@F��2��Y��u�'�by����5/$��Q�Suօr��9h�R!�\�<�IN؝���1�4��ݴ^j&��OJR [�Jw�B����'������+o�$�F}�&T0/�}P���hΞ��"G�?�Q7I�@���Ư��S�(D�#	���A$�ع,�
�:ٴ�?�f�� t��O~P�O�<�&���K�`�&"$vO�	a%�@?Y��Q� �yF _(kaY�P>�?牸}�h���b>���h�7B.=�u�'~��bb�E�ZA�6M؅'{��"!�I�lJѳR�F�@2��O	P�DyĮkulk,S(������?�@��D�g�J�vJ�+s��C$�Tr��]: e�4/�_X����K�4�A`��I3Y�\WT��8��L�L X�x�D��Z��sEҮs̥� �ݻ��r�m��;�t����>Hf@ږ�ZB��st�A��hO��b���Y���R��GjbT��u'��/6J��yFI�9k�6��g�MJRL�`����TT���g]�X���t��Pz���G1�Ќ��%�O֑W-��X�60��'��-�h�1U�1`�.�Ѝ�����y�==B��`A�!sd$94��K���b��H��,Z�d���0��,ʓ#f$�s�M�n��3B��06y�4jV2���Q�t�k��{>ӧ��4/���KDL۹4w|�⠭�1<5lԀ���54�Hu��nZ���:lJ��t*%� b���Jڧ?\e�� ]ׂ���$�I���7}�����t��w�, �B����7%���W�)j�"���޳wj��>yW��	9%��ɾq�<y�۟��N�B
	�'灻^��c��<i����c.�Y�A���7q��%>��D�#U�����*x��'
\4s��;�n�P���`���$�ikF����
8"�)�s�h��H�9t
��D�H\69t%�&*�D��~L
��БK��PJ(�qO ��d�[���@�V��%h�)����dht���M;��`�V����'�0��⯂I�<5���ҽt�|usT� �d}�i��K3X*����i�z��V#'��i��Z	m~R�a�=Qh4p���X�����_�d�Q�@�R����T��t�ڹ_V��1oW"F��ͱ���0=��#�7n�Y`Y�+T��Z#��(���Vs�QY�@̦���u� �6�ͬ�V�)���*aǘ�Q0��⋑=.��x�0�#���n��y�4�ӎR��8��S%}J��F.B e �W\*T��U̓-d"P��
1�@�ANe�'��P��E&��p�&ȫ;2k�%^�$@ca���{��H[ܧ`/�S**��-��)�/I�)�JߕE����Ɔ�2Yr��d����h� a�B��0$܂^���b�Lb�	�&TK��,�A�:�zʅ!��w�|ui��5�0���''|tk��u&0����ObU�;j�Hj"�ܒ^�F��%�<1'�� 3�z41NJ�X��C���z�4Z�3'�h�R�ǌ;�*(��+�&{6*)���q���J���u����|¤��03�l};���]Re�G�L9L�Z1W�ƗCڑ��-E>�ȕ����Kwg�DÂ�U%SN�P'*��׼Ers�Zl�\T0��50"�i>#<9�B6(m����<
8i Tg6U>(e���.�O���Bk�|#S��*��]�#%�<��\A����ͥ}�B��Fc'v"Dq�)�-�2�Sn_�)��">�@�^�}Ȇa��Lm���o�y�,��k�u�p"� >"�-
�,��hO�4	#�& �,��!���>1I��O�9�R`�~0�Z�`���'�6�Z�� q*���O�-��8ӎ�������Q�d�Cm��ǯ�����>%���:�8|:�:Ť��ΨO��ಿ5vrT����F�P�)�+�,n{��-O��'IP%3���s&nN���qJԏ!� T0���M؞��5<��dCǆL�y�Ĩ�6J������dGv�'8~�;D��a@�|'f=9�m΍~N�D|� �}�i��Ԍg�̻��Y��ybʊ�pj�Qz�-�eyhE��f��hOv���'��6m	�`I>�0� �O� ���O7���`!DB_�����'��ua��,V�$U�Qb0��CR'��b��3 C+�<Xj��"��$�C�0��$Ó��J}"VH��"CQ��! �r��0��J@�2�$�#�H;��7'�qd��Lk��X 8�>�2ׯM8�0���ה�����#LO�I`�3���e@��8�l`׭�ji�5�F�'����*��`y,���
#�*yzp��a)��E|$�%1=4!SeA�.`2$��yҀX�iٮ�i1��xF�ݱ�ꁶ|��EzB�ϔ,Wڵ���cg��b�HK��u7E�?x�A9���R���ըDl������%�Э!�\�H�N�?�HO�6mȉk�*e
`��	��]8�.�.��$C [O�I�q��7��q�2�ԕ-����P0U>Qhh��Rz�A �ÿJ�U�e��MI<�� g�d�Y�%�Ƒ�h4\0n@u��&)�$[d)q	VAE~r��c%4H�;vcpș��ߜ��`1D�z���ln~"�x��IY+6�pɋ�D�u> \�CoO�0�Ш��^�'� ��L�&5� ]�Gg_�pvЩ+O�]�4.\#^��4+�3��b2�'cQ�\�0.L%L�^��0#�G���`6G�O<T�7�.�z�o�'W��E���ix�A���!��������Hx�y����L��Je���[y��c#	�2��$��4]��#�;	���c.Ƣ3%ўt(TU�J�v4؁�\�	U���V�P����'����@�p�T[��0n��d{aA� x9 ���'\����:����&R�v�z���h�yC2�1��I�|f\#=��y7�����fb� P��\����
v�G�'�,}BD��8r�$3jWp)���'4E���	�.w��R��\!�ĥy@�ixў���T�{�F��D� �;b���=|��i�j��1̒Y�&q.���!]C,(�Qȑ<@��Ӻ'�88ЉO�|�D0c�$�?`XU�T-r�:���(&,�����j�Drt�I�$Y�m�N�1�T`A��t%B�K�̶�\%VĈ�FxJ~���V92���ɫx	��#&'J<h��D�>��+!@�Q�2NL�x.�Ai��x8�'q\7�:X��O�����)
�	���a	З8�6HbD�]�7RB<�ȓ�H��A�G�i,����
%(�,D��:[~���O(@�c):���@�`��*3�U��؃�CE�[��� C�xҩN�>��p"��$_����g��iq�41O���ɧT_L{��,6���N��\ >B�ɬ ���@��P���}1�K2��C�I��bYÖG��d�����K���C�)� L`�����W	*P��I�Zf��qE"O`(F��H��@�GO��,��"Oj��+���8�
���Ny�X@S"OQ��.�6�H%�2�õge����"O\�A��^D>M�A�M}aF��"O<�	w�?��PR��.-y���a"O���v� �\���4X��"Op�ȶ�E+-FF��5!��r씅��"O �;s��1X�m�ve�8b���[�"O<IB�&�=HTy����l� K�"O��i��_An�;"��t��[5"O,��A���N+��r�Ӧ���r"O�`2%�h��Ҥ��~v��0�"O�E�i��(�\��ã�8D<6$rq"O�X��S�S��p���dJ�=�"Ot��"ڂ�"aaN�q5z��"Oz8�Be���4��O�X�"OF0:r��!3/*u#���G﨤��"O.���DD=L��"L����CW"O����[#S�f�w@�2U"\$��"O�a���-��jӄ]�Ɲ�T"O�5it�Z)qۦ)
EG�}�\s"O� ����I,�Q�7N�\���x�"O��[�����"HͲ.�dh�"Odh������,ۯK�^I��"O�����(^XҌ�ѭ�s����"O������hRY3��թb�2��"O�+��O	x�13��ޗE��0�"O��)��ʹ1�4�ӛ��X�"O� ���t�r����� 2� J�"O�|��H�nRlqK��ҷ��ЛV"O��j�̖%�,u�&DV�}J-9�"O�,��%ډcuܵ��C�+P\�9"O(�	�?U:�]#� ߐQW���!"O�yY�K�`y0�[��*M�b"OE��"W�򵩁cZ��R3"O,Yr�ҧM�I�s�0{�`г"O�U��	O%����DS�>Q�Y��"Ov�z�0o�2R��u9X�1�"OB$�ǆ��0�B����P'|��Q"O ŀ�E�hOV���β}�8�"O��@Хݣ)�`�� �.��9"O��[e�%v�"�_# 	����"O@�5$R#n�i�+Y���B�"O�5��L�'(;LI���YV���"O(P�q�!{jѺ�� �h����T"O�iQ��Ig���f�+̸��"O����A;|�ld&�pP "O��q�^-"�a�EC��<��"O4��璆l��g*��_l��"O�m��M/!t�j�ʊ>a(�ȇ"O ��b�]E�:��وnS��"O�1�udU�UT�s�gQZb4""O2�P�j� ��}��`�7@��I�"O�e����<U�HR0 A�C"�#2"O�\¡�N�+U�v�@�^@4!��"O�d	EO`.�pS�:V�(��"O�<uDã��COJ��.��"OD	��K"tZFE�sk�]�8�hP"O:X�Lɔ([�PAȅ�\���;Q"O�(`Cc��6i��i�fU� ��� "O^4Ks��t�$�) �	�|��	�"Oxy�D�\�WZ�����7Y�z�J�"O�4��$�6Z6<��2<I��Mx%"O� V�a���7�n]�üm�+"O��p�N��x�8�� P�t��"OF��Cm'R}(��r�Qqm�hXs"O`����#F��&��?I�"Ol�cb��l�<�8��w�*��"Op|�aÛ=��Eb0h�0PР��"O�0��N04��x6Ɖ�v]��4"OT��j�U;�I�ELHt��A"O�]
ǧ�F��\�%W�}Q��'"ODDI�Y���1u�Ǩx>D8��"O�Ti%ɐ��h�(�L�%v�0!�"O>�����7n��!�kؓ�ܭYE"O8BŢAI������C$s���"Oh�qqc�8頝:PT�I�� ��"O<��q��:y���-U!.����"O��ʦ�,C�X������/q�,ʓ"O\��3�Z5��q�� _��U"OH}��ʅ;aB��v"=xG����"O��6G�)H��,�FK��ʡ�u"OLAf �m�z9��dQ`},�"O�E���Y)f�f�!��t{�!2�"O}겅>9b����ѶK����S"O��3���#.�4C��խA�.]�5"Oĩ�p%��oZp᳷I/��(0"O� ���T�Skb�S�ϻ]�s�"O.H��\�P�ĩG�lQz�"OZ�3#�	_��)0�>wGz%`"O�Y�䩘�Z'��A�بF��3�"OZD@4b�� �ۇ@ʏ97>��s"O�iz`	�͆!R�l#=-�&"O�� �F��yA� �h@#l�xh��"O�y��W�6G�|I��ɺ]~��'"O`��A��"��h��I7p�+�*O�t� �T�' <�� �V�
�'�>ĉ�,U�v�z���/Iv���'@e#g�ͧ�}�M�pN�2�'1�h3�)@	t����چh�y�'/����#�-H���Qtn7Y.4��' T��LV;P��d�PM�:z���'>��� �$��}�H�12dh��'`��2T'�M��M�U��� �'�L�s�%k<$@F�K.��Y�'�VuIt�O�W*��JGFQ$I5"I�'S<(��@�C�"����&l����'�`ģ��Y��^����;k�j:�'��ܓ�(�	w~�l��EP�[Gޭ��'\��/�-,k���S�Z�L���c�' ��苁:�.y��?l����'3�z��ʻtK:u ��A*��K�"O�ڤ@�":��d�ׁL�$`��"Ol��Ub3K���À�3a�0�"O���d'�K���˂�P!5�J�@$"O��j��H�X��
�0��X+P"O��Cd+�O�@S�m�El~U�"O�L�AkY�^Q4��U㉡U��TP�"O�<����>tR��Tm�
@�l���"O
�)��2�6(�flP)F3���P"Oj�)ƦS��!�*�GI�Ē@"O�` �:�r9�aiQ�C?hi#�"O=��J�4�� c$O�4DPQ�""Od��3�@�)&��O�<l����"O��s��ľ|���dn�7�@�{$"OxtA�K��H����MO:����"O��P���F��h�ì�[_��!"O� 4ܛQ�>��(P�"��\Y�"ON�[��Ҿ�촃�`�/jw�e��"OF���J"�d9�`W�f<9�'O �k�!^<i��,Q�@9<��U�Cc_s�<�D��V��pV�4s �]x %�m�<1���=ê��򅕌M{섂rBh�<9�$�Y�q�o�l��*V��l�<Cΐ
;	.���`��_mB8��Ar�<�dOӸ["��R��(�8����T�<y��I�"iQ ׁ�b i�C�j�<�a��-o��T�W�BH� ��k�\�<I� �������������dW�<���C%>L�:umߌJ��Y↋XO�<	�
�L`E�F�����!6��I�<9��Uxq2��6d����G#Zn�<6O9-#������[:䤡��^p�<�V�:�̔��W:;@*�S�*�h�<I'aR�4�/�9M� Dg�Ek�<�%'B����$��w�ݪ��Wc�<	�[�k�=
D��r���BXS�<��A�D�Z!���Źf�� ���P�<���ҩ[��!���4g�]���L�<���Pb�cO�,*p��x�oI`�<Q�'�3W'6�" $�CWd	"q,G�<�85�R���(Y^��iȳ��<A��+c��#�u�bR�fY2�y�kL%d�<T�P���	s+\1�yb��$��@�u�޾7[�1`'����y��
E	�TG�?0g(5�.X+�y��8ma�8"��]7�$�eG��yr!�u�UK�EJ%YjEҷH��y���6m�S�虡"��w���y`,pZ�)���= �ԝ�'�N)�yb�j>�y�Ë������b
�yRL�9 �&��р۫t�]��\��yR�ɤ<`��b
��	|0������y��͓<�03 �z_��g���y�OA�I�����曫m���yD Y��y2%� �2��&�h�>�Tl�'�y��Yb��8$(^�W͌LAdC"�yr�иT����P�Iʖ��_�y�ǟb~��G��U"��;�yR��Y�0	����B�*���yRW�|��}�U�6�( ���O��y"&^�Ri�%� �qK�,���yb-��Q�0(���/�d�����yb'�?�]`���~}�-�ӓ�yb����P��0r$L��.���yr��?(��ɷO�9y%`���$�y�D,��=ȃ��� 
^���Љ�yr+F�1�0z6L��Cm�D��]�y��L2FH���[�1�~5	���1�y���15��2�U(���9A��y���e��8��'d�]#�(L��y�[B��S��G?@(pr)��y2�)7\0����g��C��yr��M!�5i$9L�U�oR��y�]D˰\	�L�4`��0E^?�y����th�
�7) �5�]��y�*�v�5� ���JR���1i�C�	�g�V�.�&X����F�^G�B�ɔ`w<c�JI
^-�ф
�
S"O�e25��:pLA�*E�rJ�� "O��3L�?H��
ҹ7�V%
�"O� ��J���4�t�Id*$���:�"O��!��G&>DN�K7� O�@HIW"O^$a��V,M�����9r��v"O6��q��VͶ	�V;6�ra��"O���@��Rt})�iމ��}�"O�=A3��I�.����&��3"O4���L�g62����Z�|�X��"O�p����h2����K.Pd 4�0"O(��
�3R�fi�����kX���&"O,�
��l�д�c\,+I��"�"O؀�u�0y�"���|A(1"O�|��-�}Z��:���z2"O� ��V%Z4Ը@ӎ l̹&"OneJ3I��c����@�����"O�1K�e����p1�Ɏ~�m��"O�@�DQ�$��2h�	��x��"O�LX`�B�g����gH�<(ڣ"Ov+���W/�eʓES��%��y��� !�T��%*
���m҉�y�d]�j>=��+�"%@����%�y��D�o�
�Z#g�,�,�����y�&�*������%F��1��"�y� ٮ��US�M	��l�".��y�C�lX�}+�� j4B��K��y��K'Qڱ;u�_ !�~��Q��yR�P����"��(�� �;�y"h�0W٠KK��Q�p�^'�y"+��T��B�+,`x{��Y"�y�D 14�]�Q���}���p���y���p9#�; x�%i ���y򢃈0!�	aF��g�j����yr'��L�r��t��J�N��S)ܫ�yO�>�z���\AA�#�C���ybb@u,�pd�7G���8�h���y�nܔz<�h��O�FI�P�W�Z��y�i�VCH�!HN�I��KW'��yr�8Ȅ�@��?<Q�U�F��3�y��#]�.�J� F���;��%�yrk��/`:بq�9)�T)��f�=�y�l�2x���M�5s^��U�4�y�a��B����6B��_A�l�5h��y"�90�$0�b�ۧR�z��u%�(�y"�Fg��`���v���4���yr�I)��%���t�������yR�N�I�ɳ��Xr��E�3-���yB���9���颈l�BI���Ҕ�y��-1uT=�S�Řx�v���k�=�y@�6� P+2�C	Gy(m�Ei �y�M�n�D��C*��3�&hG��yүȇ"��=��߅%rܼ�&���y"��/|>XӠ��N�j؃���:�y�	�!���0	�J~6���ʗ�y�O��B=Ń��nu�eK����ycYy98�"$��3SqN�Õ'_��y�"@v�����Z	N��R����y�Iۜhˎ��u��$MJ����ٹ�y"�	4D��!��@= :����y"揯/�A�3D;�@-Z�陈�y�`L�$D�A�	Ҁ5ϲ�q혳�y҆�"K�2���	�'|v2��g:�y2�A>K����G`J'ȜXq� �y�@R�A�~<��DZ�L�PO��yR�ؕ`��0C� nrUbw�J/�y�"��[��[�����H�y
� ��i��<=򂅙���i�`@`"O�(��Z�(�T�͚?�x�"O�jcJ	+Qʩ+���^Zfe�g"O��3�Z]�0�d��Kyn'"O�tK�k�?@%T��@�|N�W"O~�7�Һ{F�`�eY0MxP$��"O�p��$�#*���A��%b�u*�"O`D�W&Zv�T���B `�p"Oz�B�fȁu-��J1�Hd�`E��"O<P��/�(M0u�ȏT����v"O�嚲mғ)b�(j��e�=�"O���4�Yg�i3�.�%���p"OH�{%K܂p�0����:1�8iS$"O^)�I�(.��FIS��Ж"Od;�Jޙf���h��R�}p�G"Ol����N�Ap���?B�#$"O�hҔ*��lU�4�\Y-���"O E�p��:b�T�k��Z+�� �"O�AAv��"g�T�W�+[RP �"O�[��+g���h�f�+a�;�"OB`K'�����c�Ok��8�"O�h��N2{1�5YU�P"�����h���'�ĝ𠂊�p �HC���&Z��'�dtA�^�J|�R�gO!!;��'fH){�,H(T�4(*���ӓ��'�Pኲ�ϡvAp�p�(�,-���[�'�(�� �O��V@�A�G�Mά=Z�}�IŞ,��E�~�z�G`�D����ȓX}�#��u��٩FϜ�s�n�Ey��'A�����Y�*��̫����~�F5{
�'K�E)��֓SgF1��É�}����d$\OTA��I'_OvDb�d�*�^d��"O,ݰ���	�������]��"Oй�d�ºϼ��A� }���W�If?ɂ�Ӹ�:�iwk�0 Y��Em�6jZFC�=3���8�D�/w����!e�C�F�������$R8U<�18S"�^g�%�D&7!�d�';�%bA7yP��F��n!�� %z��&eˣ|a����R!�D_ Al�p�A� U�=:B��p��
O(YR�R��$8K���9rV���"OL��-��1qE����[a7�y�$�$�E�P-�9`I��bO��>�M��A�,©\\ )��:�\*!N$D�<0�R�80Q�#J�8�����J.D��z�`�(�h0�'L�]m��c1D����M�al!8�#	�IT�hcď-D���u�@�
(�Đ�m�"Y���-+LO��'���D0%j�1�D��z&���HjB!�$��Ik*�����(i$���_�]�џDD�T���Z �'�D#t�H����yB�)k�I���/D~����(O^��ēk|��C�<iP��1��S�!���W���{<J�Q�!�G#[� +e�B�+@@�$q�!�DV8禙#���v"�{�C+�!��;�@��p�6�L���X8�!��Ãw,`�bd@�<�� )��.+�!�ΣPz�
&���xn�}��/�1W!�$��{�3えw��Y�S埆?�ay��O�O�
�V8���d�P�FJ��2#�Aq�����)�2q���V�V..�4�:"�:��'��>��v�z�)0���5���@Z�w�(L�ȓ*܉��-�R9z@K˴+�<��S�? 4ۤ�=u>詑`�\��J�j�"O���5엑Tw��FD< ���I��OX6�<�O��iŐ�#r*-*�JJ2i�PI�r�'��I
`e戱��-^��0H!�*qXC�I�Z`	B��ڲh�b�I�KU;1�
B�I�T!`�P�dS4*Pd��
T�.�C�ɸm>�M34A�(Hi�QN�,��-O���f?���'�b���G�]G�-q1�̀D"Ш��kX�q;4F-P>"�xV�#��"O��sCl0���(�!�3w����R"O�1���\83f%{D 1)ײxY��� �S�S�'ڈ� I�
<�1��꛼:��C�ɨW��	HP-^
L��K�5tjd"=�Ǔ���y@hΟ6D���E:E�h���L>dqJ��)����$�
F�݄�c�r����8P���؁1� ��ȓ/�(�QDZ�qj\h9�"Y�r�N%��S����$놰w��|:�ɓYRH��ȓh{v�aG�f�V�2�J��݄�P�>t"�k3WA������
g���ȓy�4��G�i�*�*�b�h����TQ��(c �,�+PLk����!>�9�G�|�4 ��?
� Ex��iAax�OS�U�H��#�#O>��iW&��y��ɉ���AEi��E�Z�C�ˀ��y	��������� 嗂%h!��R�GK�1���c`Bh��#��T!�DQ��DD��
S�$V���A#O?�!���6N�x23g�%f��"�!�D�+�Q0�&�-��pj�/�7sQ�0q��'���Q��$yϐ���Cv��l{�'�Z�XK> <��c���=���1�'Ob�x&�'�I05E� A'pMA�'!T��a�� ���W��aouP	�'4��#�R�8��"�0M�A	�'����w��M�Z�CsƓ�[�x��'v|��`�܂bst��Q��_� 5���Q>�1�Ƃ�l0� G.A���"D���d�M�+���J�Mǅf�T��!O�<�����a)��.X�-iRt���R3L2B�4**�B���V����SF�B�3%<Er%�޳`�p����
'�C�I�d
YisM�_�JAD���C��L �I`b�?S �h�D=��C䉱c��MsL�[ ��GȇJ�C�	�<\�1�`+ X[�l�<md�C䉮8kP	ѲĘ'?���X�Î3FC�	1���G �n0��k1*L�q��B�	;]O��1��<0�r�c	�;
B䉿Į`���^>\��O�4�
C�I��Ѡ���]6�Y��#h� C�	�!ʶ���KL��"��p�D�o���(�V�
�+D�O:	�&Ia� �N�!�$��|�d�"Ȓ� ��|����/!�Ć+>�8\4䃻}7�ٓ�Z�l-�	Rx�p�3jU=x��{���Jح�AC>D�Ps��U#8'���e�:CZ�۱�<D��Іa��T��}�㣛�y.,�!' ;�D,�S�Y��'�bG�s�6-,��ȓ!��@vĆ5*M�=2`���B:���OL�A��4&pքIu#Q3
I����� ���4���d��-c��Q�'1�}b��=��b��W�sZ������y2�L S�L���]"h��Q��M-�y
� �]�b
�w7��Z��<pA�"Ov��qKǏ\!�E�ɇ�-�9�"O��S����
|�f��j4҇"O���h��^�F]��kըs��l�V"O|��Y ��Պ�)�*�1�"O�+�}��v	�!Y��X%"O6�Ӆ�� @��$��N�b붸�#"Oj����
=`΁�G[{t(�6"OHة�'Y�4Đ兏`p<��"OѲA��,E`q0��Vj� �"O��k��P�"����U d��f"O��X��ȗ(��Hx�G]��*� "O�� R�ЏU"<Y5眝S�,k�"O��J�͇Bm�y[�܃3����"O�Sƥ�l�Dٛ��M�g���P4"O��ki�<5�q�@B��a�6%��"O�82!�>:�(��D�D�ب��"O��B�5��p:��P�'�,���"O,�Au�F%�V�����C�챂v"Oj�B��Jw!��qFЄ
>�A��"O�i Q��<Ad�@E�[�,��*!"O����
�T����P6�%�"O�$���O�j��Q����c�&8� "O�ш��f��0�B�U�t��yb�� 0r`�!3����҅��m�$�y⧝D��q�u��t�P��F��y"G\�	���RD�Z%� ��a��y�J#m��u��@�-u�T��&��y�^�m�H�f�L�n��{�+U�yRhݝ_*�]�Ɖ�O��80��;�yR���.��i� نpy D�@a��y«A9-0��a��:Xi�G-P�y⣙*$�TЇ ,.7T�	7=�y�㋪.6�Ck��#[�p�vB��y��7mr�r�Λ&K�*\*��\�yr����D����R��,
�l
��y�*K�~�e3[al��ab�$T�,��&�Y�G����x�b=��_��9lJ�0궵�l�=�δ��'�0���(ZVތ�j��-����'��ˇE=KhN�q@
�#�h] �'t(@���ah0 �!�Ae��'����W=�){�cL�Z����'68y����i�`C�MA'`�a�'���	�J�*q(�a)!�.Y	�'�`�� 삄�4�`!lt<�X�'�"p)b�^x��1D�>z��)k	�'�*Т���9@�\���Mtk����'�xWhEV-6Mj O�f,N 
�'���beL�q�(�D�PCfi��'�6-N&�ت���S��XQ�'F��3�ޒ1��,;�GB�\�L<�
�'�>�0�N;���P�ݛ$���'�����&m�.8QGAp ���'���0M���u��(>9|�9	�'�F�`��*��$��FƹK��'[�9sBL�`����s
�<s_�q�'��e�3�����l򨌉e��IC�'�邥)��]j؈C�bU._����'tHէR7Bp� ��F�-X�a��'W�\�q���xE�1�m�V�<y�'�MS����`qѪ��U�����''��*���$�M� XQ�K�'O&M���D4C���;Kₐ�	��� zؒ��J<�D�BQ��:��P�"O�@��bS��h� I�t����"O ):do���tb��ȫd6N;$"O8A��%ܭ(D�\i�ă%%(�H  "O$���/<��d� �2"O.��6K�]Ű�"b� Ӽp��"OƤ��&�� ΓD�L�z�	�e�<9��ϵÞH:@ǚ�!`ġZt��{�<Ac� va`i�tf�n�|� %��t�<D	كWB��������n�<��� �9rU�P�^, )��e@n�<A�G�'L��u�MV�>�Bt�C�<�f�=oC��)}��H$�W�<�u��a2f�"jȞV�@�����R�<�CD�(SX��#Ǎ3[ä�(�%Tg�<I�`[6���;�β����@'c�<��jӚ)5o�n}M����_�<!��F�q�V�
V�%�A��e�<�&
�c&�����+#Э��)�|�<��/�3����g�B�W�Jl6D�<A���,N���NQ�(�� �}�<�-9 z��歑<Z�Y�%[R�<��O�ayN���Ƌ�-�Lȁ�Q�<��EJuR�xC��D��aX��Ce�<ġ	�(@{���R�q,Pd�<I�$*\Nth�&
F�kb �Sj�`�<���;Q� 	9�x�����`�<�Z7.�Y��OƓL�h���$NB�<�Ī�$�hK�q�|ڄc@�<�s�3}@l	�`[d!A�^}�<ї�S��n�1�K�.�pH��K�d�<Q�bZ��t���)��\����`�<�IVN	�5�␷m���e͍]�<���0�� C�zD~\�Q[^�<�c�K �%;Ƥ��"$��)�[�<��*�;'�<�ǆ[�Wֹ�E�A�<�ŀ>B~����F?(��=Q�ie�<�T��*=,Ma��f�!��-�|�<Iůˤ2"d���+�vI��s�<!�
�
m��iR��`��0�Ld�<ui0H5��%^?6�;�K�g�<3l���"���圻�Z��A^�<�ũP8���P��C�x�s$OR�<�r)�=|�<��R�N-����Z(���M xc���yU2@pv�_��t�ȓ�Vk� F��LA�̡!,ą�.@%�6�q��ك�� }1���ȓ(x�M��ȣi#�vo]%<������\� �-�"�2����(��y��o��(ҳ V�ƥ�@oD��2a�ȓ{�" R&D³��"dcC2�� �ȓlY����)mz�x�'��zJ��ȓuX2<���S�	�0��!~@���ȓir��*f%�-Q� ��,�S����~�|�%���s�\���捏	ˎ]��A��`�A�'������H�yF�t�ȓ}�dJ�M�3|oMR�o���m��\�:р�AӍP�\Zb{B���Z8����)
P_.�����3q��)�ȓ77É�:�2ɦj����-�v̲��.:��d�F(S$^��X�ȓ ����D�~<��D�^�F���-t�"��A5F.u�S���x�Bɇȓ��y�R��y�h I'i�,Q+P��S�? ���Ɏ��rYʴ�
�,�Hljw"O~%j���a�����'�LH��"Ofx��e��x��B��[�|@�Z"Ot�tN�0R�3� DH��p"O�����K�d�
 k&�x+4!`�"O�+����4܀��Q�"�TZ%"O>�ֆE	�����߮x"���"O
y���J4^��TwC^4<���Q"O��w霰o�m0�� �Z��"O�\:`�;z�<x@P�D9� �ٖ"OZ��QmJ5d��@X&j��=R3"O��yw&�3��%��S�v�t"OVԛ� /�2������>yXR"O*����&]<�;r��Tj�P3"O��H�A;B�̃�;D��q"O�͒R��in1��E$�����"O�����_���
��qϲ�;�"Oz�)Aj=z��};D�0�&d��"O`�#���/g4��v�̘U�h�D"O]�f��*Y *�c�.$�j��"O��C��A�t�Q6�K�'{����"O�qxa_��N��xA֬;J��yr.C�H��`b��B�m&��ѐ��y�FVo��B���1{�`�c`�^��yR'���@�6G�:v	 �٢���yRM��z��#�lȬe�q���yR%���9p։4X��X��,�/�y�M\�5]p�A�\c(:U���/�y'�x��%��T`W>�ʵ!�*�y��@`1І���V<ju9m���y�*�#��1���R�੺ `��y��G *v8�$�\D��P�H�4�y��ՊDJ�0�n]�'/h��� ��y�NH+�6t{2�E
ސ1�H��yrg*aI�T�FI�\���K��H��y�)�E�t�å�J�򘀠�R��yr��b$���TKQ>H��-�w.ٍ�y�N��N40v`�.8�
tH6iփ�y�o�%Uk: 	�6L���`���y��N�&�(�(���"ht��Ql "�y�KG:��͒���h)��c�Վ�y���n����$�_�%)����yb��y��t"��+e8`�1@_��yBO��C��eeM�;��&M�*�yB�	y:YۡJ� 5X5)�[�yR�2h�t�Ơ	be�(���і�y�i��5�,T[G��!`
6�b���"�y�C�s����:PI^L�b�ރ�y¨G�n9�z"e�E�VܐB����y�d�*�d�TMY�`!H�.�%�y���<A��u"Q'�v��pL�%�y�E�>y^�����xrP�q����yR����yz�C�k_��:S�՜�yB���K@�<��F�\q��{2���ybD�C^�	��B�v�H@��yRR޶UKC�� 8���e,�4�y"�a�h�jgF�).กؔ̋��y�"��
.Ta��.�v`�֬�/�yB��5pn.<��m��*Jj�i�X��y�Vs��\��iH�4�^ir�
�$�y"g=G��R��;�jT���
��y�H5,<u[e�.2~|A�-ȇ�yBhKl�D(�H1���t��y�L�
�X��T#_�+�`D�E��y
� pЋ!�A�&d���.��q�Q"O$Ձ��5B-Ј�ã[ �F��v"O�q���'!�^��#�I!&�
�"OD� �&
�L֜
V/]�q@blR"Oօ��f��j���;a-�#�R��"O�Dc���f�}��C��j�Kd"O�"��]�m��2GJ�X�H�ɐ"O>)��aM$!��e�ҧ��6�j5��"O�����\�_`m��G���"h��"O���%�ǃeRT9QF��oUb��G"O���c���y�����/G<B%"O�gˆ'K�q8��S�w�����"O�qB��({��t��*'b@�*�"O.�iW�Țf�f1��������"O΄�C��C���鰄e�� �t"O��0��[y@�Z�c�+\s$`�"O�%!I��4!�5��"[n�x۱"O*
�H�N!D��D�4���hu"O���h��I�Z�" Q�I�$豗"O��ȇ��X�<��� KdH�`"O�]��G�*D�Da+�m	Lx0�"O^�ҕ���� ���/�XӢ"O�jD̓#KK���c�<�(�R"Ol����2DPjl���!ff��"O��@"� ��HA��9_���"O�|Zs�P0+df��Q��#D���"O�!w���>�]�@�A�d|8��"O$hP�k[�j� �c�)�t�(�	�"O�8��4;��娰F˱�ZiD"O��(���8f��9a�Y>=�M)A"O���_5�dxjU�J� 2ҥ�"��e�<1�ѢD@�L���U�~>�ܘd&�_�<�A̙�s�����m�<���`�VD�<�2CX#Sg֥�喋g�ԙ ����<I���'^�N�* ��
Ɔ��u�<I2��pl����ӑo#�i����{�<��OU�{�X���Ǝ/�����{�<�3AȘ8b��PbG1��iv�Oy�<q�+�
p��<3�hȩmcj��rh�u�<ycL��胵'�j�9 �Ro�<	�/N�3\�l���|˜E;"I�T�<��bޓv�Hkt�[~q&�"K�w�<��̱+������E��ՌL{�<�fM�n�����@ĥh�$���s�<ysǂ�s�<�$��L> E�n�<��ޣ\�Tc�N�	��")�~�<�G�.���(`�WW����.ZA�<��8}6B�����a�Q�A�<	�j��:\e+���4l:u���y�<�Q�OA�x�W�|�nE�r_�<1%���'��C�+J,�g w�<1�.N�F��Y���'/��I�5M�x�<�P�7s��S��##3|)Y�"�u�<����Z)�0Y懖l��5��m�<⠟v���A��t2 P��O�<���1?�)! C�=826�L�<�EB�'g�(a2.$�T���]�<!�bT>ss\ta��'��0��[�<�uI�
j�u�AǦbV�Qj�*_V�<�f`<(���:Ţ��iӄ�� �|�<���Aՠ�)U�lLl1U&�\�<��C��mB�Ua�@04=�H��]W�<y����Թ �ժA\���tg�V�<�F�fz�>6��".�X�<� ��clʮq�Hq�Fn�uR�=�""O�y���b��Ы�B�KX�Yi7"OY��>|�
�Sg��c�q�"O��ق�߳V�0A����O���"O�A�t�T�-�(%��n5F>u�"O�9��Ʌh��2M�3,�`�"O�3'�^���J
�<�~���"O}�⁖�t=�(��M�Z�b�P"OPt;Ú�2��Z5��]����u"O\C5�T)�V|
D�
����"Oh*A�8i��M@�J��B�*�@ "OdͲ�+G�.2XY�c #E���0�"O��"�,>p���+��D(@"O.ݺ��Q����/���a"O*�2���vA[����^(xG"O+OV:l��	�B�ԩb�9eJJ�<�q�ɇD{fTzTÃ�b'�ڵ�]�<������"4ʥ"����B��\�<Ad�Z@#�M"�)Z(c�-j��s�<�5�S�syJ{v�"{F5#�]n�<1��Ō$8��kш r�x�sOf�<��`�:_��s4w�i@F�e�<��
dF�q�e�'4-���b�<a����EK��@$>W�HA�<C�	oS��E�8I�8�I�C�I�ۈ��c#$\�����L7��B�I/܉���6���K��K�q�VC�ɆsH6��4ϛ�Kn� 䨈<r�C��|���!sV�Qʪ<�DlC4�xC�I"�}�&��o�ZD���P^C�	 �Pq��ףo����ܾb>C��q3��K���
H�`Ix��[
�ZB�I�\F,}�`1-�*- AϬ!E�C�I5 '��Òΐ-��=�V�_�x�ZC�I�K����Dֱ/�x�n_�=l<C�I�V��	��Z4� �Hr�۪YG&C�	�bj��J`�֖}z��[5[6�
C�I3}�>T��	�{�~4k�h�e
B��8>`�b�*�X�9Fi ]�C�*v�ڴ���N�WR� �o�;��C䉨.e�@��	'����U�G�`B��+q8аBA��'<	�F�zr�C�	1P)�a�a���o�xm��"Ob�`%-"�P��gM!��̃�"ONQ٥��i(Z ��(�湊7"O$u��,OD���	���=v��`"O����!pR�����9auF��"O�#��0I����P-��<cf�٣"O��B���c/0{5�5I�$K�"O���O6n�1I�(}?�)$"O�q�Q.��F�5*�<ώ�`"O�R���u�q�e'Y��!�"O��H6�4J�j��T&�S��K�"O�$�ૉY�,|�H
�2�@=��"OF�`�+�,m�Y8q�;n���"O2�;�*�]Y�\��ۡ�XPj "Orxd�G '��%SU�/S`HjU"O��ф�>�&�c%�3�a�"O�e(3jC�U���ɀ5(j�"O[�!��7��|����'w��D�q"O�|
wb�VV�Q��C$��M8�"Od�3��-C�jT#f˴-�d;�"O����G��6C(u���#���
�"O��� C	3T`@pA�ײ;��q�"O� �u8�o�Z�l��L�l�ܐ�@���	̉	u"T�p�=7Vb�����*�!�X�T1D�t�V2h 顦܅9g!�|{@ �%K3�D�Ğ?��B��}���B�
"nf<ⶆ
"ChB�I�J�|�k2,��fMBT+�ȉ??6RB䉓H��H�`�9<�݀��˸h�~C��	PA0������&cK�RJ#<���?b��0bk�D�0+��MH����F7D���c E��	FO��4x��*D��5Ӧ@�B�rR���?D�� -4D���`I�#�f�$�σar��r�2D��a޲L�0<�6bO�d��ZTe=D��J�m��)#���AÚ\#��4�7D� �a�%������^�ng��� N2�I]���O$�j��0uaQ�\�<���Z��y�Wvs���d* �>�th��D�y�刲�.�,ޅ=�pR�4�y2+ˬh
���@p<��B�R�y"E�����ϵ0�$c�&X�yR �,2�d�Q�*]�7�L�B�ǎ�y���
<Ѣ�SelB<1j`�2�	���y�o�@x#��}\U+G�!�y�/XQ$�#���Q�M�vEه�yBD�#ǼeZ��S��9��߹�yA�8Ĝ%3�-)S��a ���yr�O0DnD����4l@Xi���7�yb�)dՒv�L�-���Q_Z�<��р�x�;B ��	��}���KZ�<���V�-��dJ"Y�:�Pu.�K�<�ҢˋId�c�"J�0�B��fI�<�Ŏؿ��� Ӭd�4|Q�F C�<�D�(���a�M�0�� �Zg�<�aÝ��Vq� @	<�`���Jb�<��j�`��\(��0�x�� �Y�<1��DB�2�oT�0�L��Y�<�5ý+tT)� "�!`���SNZ~�<�Ԁh!��±�T#>3}�S��z�<�I�ZcR*rX#dt�%ou�<���lܐ�Iq��O���r f�q�<����u3��ƌ��P�W�<y��ۖx�<��N�R��ŇGh�<����KM!&�<��@vC�I��i����{��Q���B�	"���:�FTP�:�ɷa�O��B䉹?��͛�!|���F\/0��B���.q�PRo��	�s� !+�B�	2Z�|%��P�i�4OݤQ�C�ɥ|E�pi�P#hp|=s�j�?)W�B�I�3������Q�f���U���B����Q1�[�a\t<�p	��%��B�I+1�Z���8M(푄,�$�B�I�q�
���j�V(��G�oI(C�ɲ>��2R�l�"(��jѫ f8B�I�:�����ē$�����	Z��`B��*=� rC,�"�X�q!�Y�bB�Ɇ&BL�`'n�+����֋>9B�	�$��[wC��Y@��kw��.�(B�	�0���ȃ��C�)0/8NI*C��!Q�|4K��?��Sf�Nz��B�	�Pe*X�4�8. �s�р-i�B�Ɂfo^1Z����Z�1�F�� \۰B�ɑH\��q�]t~�r�g�6:��B�	�9��	s��aƨt��F̢MulB�)� 2�S�oĎGdH&U�qxDAx�"O
���c�'>`fp@�TY@���E"Ojq"dlKB�����n�4�ӵ"O�}�-�N��xs(�i�Bѷ"O��a�+�����G��,.p�5"OF��1�0N� X�`��;E�T�d"Ox��7�,E����7�̡qN��"O¥��oEN���a�M�O?��K�"O�="�W+Ek��q,�J+.��P"OԄ�"�ѦwR��[+W�K�q�g"Or��c߄v�[���sk��"O^�#�o�#QP܁С�t��"O��k�)A,���b�W��nIA�"O�	��b܍\�,Źp��	~�P�r"O�1�VN�PPV�PKSvFmS�"Oh�@	S�^�v��1)��Ѕ"O9	�听NS�B��?(;���"O@!BhΖF+��L�� ���"O�쀤��w�&�*b�e���� "O�L%���MaptԮɴV{��""O΀*�86��	b�2��)K�"OBY1�)�`�QBc�0Nz���"O�M�4f�h0ZH�B��;>�|�"O�1*U�.Q�"�z�"]�;-�z�"OPة���y2�j���!#�#d"O�Л#��,>d��o� �t�b"OX�`pKX�{H�ZC/_FLbu�$"O�*�..M��x�3.ϖLAb@f"O.� ��˝^�J,�C��_���2"Of��pk\�n�:����F-@B��C�"O����U/7�ݨ���)8(�;�"O�Y�6m��>�R9��%׾M2N��v"O.9`�[�Gd�P�7��*e ��A6"O����\����
�-P'r \���'�l)s�K�2��0��kh��[
�'v+M%op���UaWt��v)D���$ʮ$,^E3�G%�p%-&D�2�U�P����i�-R ACw�$D�,��䆀=��p���ũ-����&D�$�S�Xh��\�"��7f�v`�'D��+�LC�wΕ�QOκ�ʴ�&D���N��X���J����0D� ID`�0�:y��b�!Wz0�-*D����� 5~h���T-a�ZX���"D�� ��\�4�ּ�b�17������>D��	C�<H����g��1f�|�E�7D�l�@��=ex�A'��!�L�Æ�0D�(�)^%6B�Q�#U�Aq$0D�Hz���*^z�`��O4M�U��#.D���!��(s%Zx�B�c�ȣ�*D���.�v�����Y�>�r�&D��b5�_�"Hhs�g'-'v=#Ǥ8D�X�k��AG���QlA�$�T�p"�!D���7 ��ryhT$� �2�A>D���LUG���b&
T&M�qat�:D���J[]c���ş=(_��R��8D�hXī�e�ŚG��/g�h*��4D��%k��`h�H�!�1u��Q�2D��� ���T�yq�Mm�t�X��2D��Y6����l��6g��x��Ss�,D��JFi��25�iq�� ���B�G7D�p�Snɶ)� �ipc� @(�ey�@5D���3�ЙM��5�6h��'x��b�>D�L��Gԉ/N�%����%X�&̒&�;D�� ��8EB�*��<�w��8d�v"OV�c��Mv�4���X0����"O���E8,�&��OVW/	��"O�[QP��1I`].Xl�R"O6 2�! �N��W/��<�ͪ�"OH�*��2W(�0�M�/4�B���"O�A���1],��U�ם=��<�"O���fo�"��2ҾPܘ�в"O���4��1uL+�"�bҝy%"O�U���v�3��"
{NA�"O(�2�f�m���YD&]�V��y1"O�M��^�tPP�@F_�|��l�7"O��E��3[0��S"
��]��"O<�"W	 `�r�J�ċ�o���y�"O"Q���+x��0���X�5�p'"Oh��sG�6�����9Ǯ0xp"O��a�KH9�Z�x'@K����0"O:�"p��5kʀ�P�H�d��J"OHP��/�>r��<z���]pd��"O6x��iEh�zB�3aa��9r"OP��W�5-��6�MWM�`*"O^���@�ᮼ�A2"VB9�T"OH�Ӈ�Дk���Q�Ýw��:�"O���s�^)-  �뎬C����"O�DKc�K&���$�,
�QC"O�A�H��(�s�BX�x��"Of�[�f�e�W�P�JB"O�F\c*+[!�m�hʀ�y�E'{l>ȉ�!Y�r��5��y�H���� cMCJU(��U���y�D�'!.eZ����A��<�����yBlD[EX)A�E�u�ibu��.�yB�7]&���k��o7��9ŀ�y��ƞ6�~�r�� �nV�/,Մȓ ��r�X�>��}���!iUHq��Q8�8�u-�@���惖:�� ��A �l�G��8)�P�{�n��gT!���N�I��� 75��t�]:FA����ii���6 �:j]NƊ&�*|�ȓ��QsuMO ]��i�S�K�#zp�ϓ��?�G##3h�(Q�T�j״���(�w�<� �B�����Ůg�����Y�<�7@�%�ZmؑJH�0����'
�S�<9�L;m��@Q��y]� Ձ�v�<��OJ�H|�Q�)�ĳ�+�u�<QQŎ�@��p��A�%hbDeSg��|�<14L@;l��IK�`���4;o�{�<�2L0E��%�Q˂8x� (�}�<�I,zx�ш�8	/��B"�Cd�<IR肺V*����=\�RD�%��b�<��ۀEJE�0!Z<E`"���u�<��F�,�.[`&[�S��MJV�Dq�<���<���@#T��i��Kj�<��aR�|�i�km�b�@�M�<���P3v�
��}�j}���F�<��1��`�V�/��tH�LZ�<�b�23�\ �i�8h�-�Y�<��>q�pDh��9!K&��rd�S�<A��/<��a@h]4q�v���J�<����D��]R��A3�Fl#�Lo�<�cH��)��tc��Q�p���e�<Y5ÒPGv,:6 �*����d�<Aw�`CJ�w*\����u�<ِ@<<l�g������1�A]�<� ��t�%w�*scO�wht�S�"O�ȉ�������.�"\]L��p"O"x �iW�2�i�FɯZX,`"O���v�}t�q���{X�t�A"O��� M�V�*���V4^V�˔"OB<���6!J� �B�"4�iÀ"O�K`I� O� ��4�;*$6٫"O�\��E݇z頜��� 5edy"O��r�Q8���jZ�*&��bU"OD��D�7Y����)�;[:H�r"O=gF2:60(V
��q�T���"Oz�sl��N*�e� ��) �m�"O�}�1�4��+�P3V��0"Ot#c��-0.Ȥ.)�D}�"O�$	��'(�p4�'[O��$�7"OP�Q1O��l�x��.��5�"O���p��vH��x� ��U�7"O6J�'�S�D�U �X��ې"O���''��0&�Q��!�����"O����ŴY3ve�"Z(o���hB"O�����8���WMRl��+R"O���2��/���kөpJ�b�"O!��a8y�K�-aڹ��"OrL�Я�*i��r4�.�L��"O~ �@�]�J���FI�w�1��"O����	�n�x�D+Ҟq����u"O`!�rD�\�^���$/p4L�2"O���$J;l
!�v#�'+3�S"OB���6h �|p3�
�(%����"O2�ꝍ;�) �Q�:,}�"O��	5�6*�* ��K�9Ԫ%9w"OS�b�6���҅�"w�PEQD"O@$�e	�(�����N���J�"O`1�%țF��H)�פs�uJp"O�i03�R�\�ƌ����[�0��"OHy*��5I�V��,�Y�|���"O�U�b'Q!/�L`�CX��M*�"OD��"�*F<H�P��D5+$��xB"O<Łcd�#V$n��PO-l1����"O@U����
-WΆM�D<Ȣ"O�C#��#$��8�����8k"Oa�D���i�m^X����"O謱��>s�"� ,� V�5�!�ށZt^D��O��~�^���-<`�!�őy���-�������&�-g�!�d�-$di�L�@Ѧ��j�!����������>tޤ �Ff[�OM!�Q�X'$���o���)#f�aL!�Ğ�dR�����>E�:5�F��!�� TN���+�q��9d�K�Z�!���<U8�!��$ʌ�����$;!���W�����ɬn�& a�%͍M!�DM�bY��0��'��]��dR�e!�6]h00�)R)�h���!�d�'�9�q�Β8���yD�� 	!��.&�@�&�~��铢%P�C!�D�A���c������p$�9!�ĕ�f4P�啭7X�g��,l�!�d��DJ%b�4lT���2M��Y!��
�.�8���℟Xhը��V5m�!�d��n0H2�
fjP��Ev�!�d�O �5�W�>Sd�Ԉ�BƪL�!�d�Qְ��$/]J��*YA�!򄄬�>�*��]S#vH������!�� J5�Ĩԑ:���C��D�OӰ4��*OfeS�k w�h���R�H%��'�,p �2��u!��R��%��'zt�'��z�<���)z֜e��'����q��D�	Pd�W%vJ=3�'B0���%�1�yfd���'������FJd��,�=p�vP��'!ڀ���I�W���vN)f��M�ʓt�(ŘQ��3V��t����%?�͆�k��t8�i�ª��5�A�X@|��X��RI���d! "k��Cg.��ȓX�bY�vj�<u����qnQ�~[N��ȓ{OT��v #dOfɪd%��~����ȓ3�`aw��-m��ҁ�Us�ɇ�R���W�Ąc�l�g�W]LH9��Wꎬq�j���d;P��c���ȓc~��2B`��vG6q�iKY�X���/����"�t�t%�)�kQ,���FmX�Ϛ+/���A/��1|�H�ȓv�.�J�1y|�V,D�N�.��ȓ5��u��n�:n��`�j�`�����-�̀��ɟf�0�KcI��IZ ��V��"w��S��҇p��X��*yz|)��^�[:F�ѓ/�<�z=��OI�$SBL�R�����O�n�Y�ȓv�<i`�&	�M\��FΧJՈͅȓLUR�1�+�� U��S���2������t��٭\U���w��3%�J��ȓP���jɌ~�,=����U�\�ȓ.Wt�$H<H!��t� �ȓv;�̡0�^,W��6m�Me~���F4��j��D� g�X{c���7Z%��Osn��DI]�4����7dэ|M|��ȓg�v��!l��b?�U���+p� ��w���Οen��K&�B�����O�����#�d����T���ȓ I�80�I�\:�yr��0�fU���.�`��9S+��YW�?~sF��ȓ��8��-B�,�	k��iO&(��Q�l��զR�t^��Ǝ�&xĆȓM��X�@h�!t�I�riI,����)~��ej֚L�h�W��J�<5��J΢��'�*d��\@�,��7��ąȓK����c�[��Th�A�H�����h1���ɔR��#e�Z*J����G! G���_ƴ�K%l�"I��!�ȓrL���!�6����\�B�����pf(	��#��4� �4�r��ȓqRP�h!N�
���k��y,ب�ȓ4D9��aѣe��yc�e%r�9�ȓg����ƾ�>�1�E>�Α�ȓO=f�,�T*  )8�`�����M�<Q&)E�*Td��B�f�]-�A�<��J�Ve�5zWOG�c�h�0g%T�|�!�݈`�v�8�d��`��`�Ɗ5D��H Ș����ң.šg8 !�5D��8TG�:H/��;tℲ)�̬�E�&D��x�Oףh�4���T�V�yс"D���̏8,��e2c�7*[0�j�!!D�0��ѺWEd\bӥ��x�P�h#D� ˕fږk%��kԊ��B��͑��6D������Bf�a���3t~���3D�����_
n�m���ըg����$3D�������s�h_)b^`<�D;D�� v�A΁�t���G�FV�:'"ON�B4�N*�={gf�Bn���S"O6�b2��WK�p�Bg4G� "OT`�$�	bbJ���惙j�}�a"O�a����PL�Y���6[j�	8�"O�bѠ̜RYX-��&M����U"O �Q��Q* H�i�#�9hy�"OjXc��������4^�ɚp"O@E W.ӨhoT	(�a׬YY2��D"O�����	%��d�Aa�3��#�"O�!���X�d慑�\'L�"OTM�DCWzF% UfE1��\R"O�9ee�Vǅ��X�i�"O��y�G�t<P%�&��8�"O̔�7�[�F] �`�2t.P�X�"O�0v�ڥ#jّ��)#�5s"O�-��l�b����c�u� 
4"O��Q��,��=D��^]����"O[W��@7ZAYc	�Z��`�t"O�ES� 0�c�ؗq�`��"O��Zu�_������b�8Tƅ��"O�����3f���d��4NH�d�"O���R)�N�BВ'��
L8��"O�t@���+�H� 2���E�i�A"O@��E$�4=��(k����-:�Ț�"O��*�_�T��0BM����3"Op}�a� $hizaÈ�Hr�!�"O+w�=���C��A��"O� `�i�&��t��8�Z�y�"O��x��G� ^
�h�.زF"O\p��LP�.ٶ��G.�+�JI�S"O6�8�W?H�6m� ��>s� ��%"O�si�B�L�3�뗇��}@�"O<����0�"�KckF!.#��3�"O�X���	⩨��K w�Z�H�"O�u��_���9v%#j�4�2"O�XxRd�x�� ��`��e��U �"O 
�\
�S�/���(kp"O�H���\�`@����T�s�"O(�K`���4��m@�c#:U��"O��*���b8�P8X� �D"O�T{r�PxJ��kw�)_i8�"O�u@��6s�t�����"L�A "Oı{�/��'VF�P7Ã2P&�	"O�3猃1�:��=(
�r"O�a�4ͮ ���mɺR��)�1"O�p��ЫQ�nL�fտg�h�B"Of���c�`�J1CR����=��"OL��F�<�x�PH��'׾H�#"O�=�G��FBHE���3��E
'"Of���@�kPX�� !�� ��"O�BSB�&+3B�h��F�l��aK�"O��C7��{E"9h�f�`���"O����A�e3v�Pc��
=��"O�g�F�>�RɸF-�E��hs�"O�x���\��`uK˜	��Ce"O�T�Lѹ>m`�q�']F"�!p"O4R�NY�g��UiP��TJ�B&"O�,:V.�d����ef�8P�)�"O�<p��i"�h��9���"O��i�  Jj�Eݹ0�F�jp"O8���� o��rG�M�.q�"O谶�"E��!��y�&�T"On��V�ҫl;֤��đ�}�CF"O� �i#�(Ƚ;W!�E��5��(��"O�1�B�	`=�L�T�4�#A"OH�ٳ�ǆu���p Җ�j���"O\d���ץB��5HG�Z�*0�"O�i�g�!X�:EK#�N?\�)�t"O���RF�VJ��q)W%A_����"O�)ۡc[-�T4����2cl$h
�"O�M���|I�� ��	=}S����"O~�A�#�a1X��Z�8�"O8y��%�]�d��̞�b$�"O\�9�O�'��J�M�X�DG"O�,X�F_
%�4'[Q��QG"O8��F��o#t���/'��mb�"O"�Xf�.L�h��V7z{`R�"O0�q�L�����r(�=��`��"O��K���r��r,�j|��"O��#��$rz%�0,�q��"O THP�\H�0��"ZX�R�"O�Ĉ⡞�&X��8�^�"O.}���b~D4����,^2���"O2�a���,Q�мO���1"O��r!$�4B���0�fYe"O�p�Nb ��B̵F���T"O�@*A����k��^�(a�e��"O���-W U���Ʋ5dS�q��"OD��@��+-dt2��I.�9g"O��GhJ�0= �)��ƌ_�Ҡ�P"O��:�h�$m^���K�Q�⥐�"O��H�je"��6K�"Q� �+w"O�}�sgƧvд�;f�X:F`|�Ap"O���A+�,@X�'\�/,��h�"O�����+7L�p�=q�b"O�����C?wEv�䥊
o�2% $"O��˴�[�e[�� bd�l��%��"O���v+ټ�ʔb�'6��93"O�Q`$D0ɾHQ�A����r@"OضU.p�����/4�9�7"O��(��H�z�ܻ5O�)::��s"ONHSW쑜lӀ���N�(u�1r7"O�����N�4�SO(&�E��"O��qT[o-�P��� DLKa"O�AeeK�Dh��##C[���P"Ohyr�����|(�g�ȷA���"Oʼ�F�>�^< T�N��ɇ"O�-A��ڑq8b�z�hD�Iـ̋�"O�I봅[�+Pн����E�n0�@"O���-��(t���	X�n$�"OVI���	@�:�"6c3?�y{�"O,Њg�/q�b�@xm�'"OHZ�P
'(��FOȪ"��c�"Oؔ�se�J]~����B�z.� D"OB��VE̳0m�}YC��E��w"O�]"H_�Jd���aՋ�*�(U"O�L� Iʲ���H'ᏗJT�w"O�pD�[Jh`�D�šGp�k�"O:	Z0���:��]����6&x)�"Oz-��A��H�T�3pj�@�p"OZ	���X7J�p�)��S{��5"OZ��t�ȑ��!��g����"Of��s	�nZ ĩ�.[��Ț�"O^�JA�/����S�$�\�IR"O
��g��L���	���g(��%"OL�K�3ؠ�ed�H4tyI'"O�1��*l�R���Mw�-cd"O� �y�eKS"���"d�T���Jw"O�$A��q� "Ă��
l+�"OdM{��C(}İ�Xd�ِ5��	�"O,ؑ��ٞR�[���%5�-�'"O�]�� W�"~�`�@�Z�/.,x�"O���!oI���x�:h+Н0�"O�L�%��B<��+b$*�I�"O���n�|�"ŗ`c���"O�MJFΑ-�,��� Ud|��"ON�Z �ߌ'ⵓ�JR�9^H9�"OX�J�KX-�Ag�+$8���P"O��;��Ƙ����46Ȣ�4"O&�J�J�V�u��%5�vԈ�"O,�S2dX8b/� ��m  A�Bp�"O$���h��P,���r+8p&���`"O~$Pfa�,NG��A�=^��"O���Û0+r޽)0�ۃq���s�"O\L�0�V�d��Xi��)E��l C"O��b����rh��p�d��"�H�`3"O�9T�H,�����FY�E�.yF"OJ��.��=�\��F��?w��Ic"O��@W�:��&f76��aR"OfE AM�c{�I���25��A�"O�Q�%
�(���M$�`	�"O��2S�A<e8=c��Wz,���"O "�դ0PT�X%&�KHL� �"O�,����'�<|�5l;^��"O�� κ �Z�ڼp
 1ؔ"O��Z��@>E�ecwC^�r��Ɋ�"O&U�A�cV��B��6+q�"Ox�� C�,F,���M�4��"O<��RK���a�ï.X)�"O�P�j�j�1�F$��\����4"O���!
�1���)���4��M%"O iK�	�]��ŧ�s��hhp"O�;�GMe��1t��!���q"O����̟'5��ʆ��AȺЃ�"O��0�L�RӐ�i�+E�0��z�"O�����5	(�U�	�Z|H�"O�PYd �0j��J>v�\��F"O��a^�`t 9p�B�m����"O��6e��T�$�k4���{4�w"Of��F�L	������rT*U��"O�ӣҗX 챺�Esd�S�"O�I��ʐ�!ѮG,&S�X�"O�t��k�<v�8�� 	%O9��8V"O [���-�ƍ�c��9#Y����"O8aX���(f�r%O�`Yx3�"O<����2x�N	c��(=����"O$H�E��h�}ɱ�_�b"����"O��@�U��r��wj	�W앫�"Or��`��w����CW�.N1@4"O�	9�\7��y���$�P8"O6@H��.l�x�����r͂�"OxX���Xz��u�E�^ABLaP�"O��
"$��k<�-P��ް#D�L�u"Ov�cU�ۄ��Y���:2���%"O���BGJ�(������y�.q:�"O�P7��Hֶ��U+��T����R"O��k��LFbtqU�$Y��p�E"O�S�(Z>�ف!�P�dz�@��"OMh%'�(*���Ƞϑ�<r~Ժ"O�$�T	�E��-&���
�"O��C�D�\B�K�,!�uz�"O� �Ր�n�$Oo(�(�[�- <��"O�AS�i͚j����Q�D1nX�U"O�pj���/tĆ��"��U	�"O���I��0^H�����l���"OXi��o^>TڌY�P� �.��"O���5a��Dr5�E[� ��"OΈ��"��,r�;CӚ���"O�Y@C���� �5���"ON���b�Ag�Y����	��i�"O(�x2 ɞX~�0
Dp�rR"O
��fE)gѾq��-�$8404"O��t�ږE�8(�����2�p���"O\`��ƌS�<qBwEǛO���ʀ"O����
\�y��d��,�D���"O�1:7�߶&^tQ�#�b�`tR�"O���A ��W�"uD�ӽ_kb�0�"O�86�߈9���!3 �:Bdt$��"OR}����|� �`�^�E�"On|��W|�C�԰2BF�Q"O�9eM��iH�'��@2��ru"Ov��2)��J�"����h��GK�<�F!� .@���Ǌ�=���$ �E�<�S��?�`�� Ȁ�{���Qc�E�<��o՝$��	$��r�D(r��Z�<)s+@)5��Ɉ��&>�r�D��p�<aT�!�@D��@�$cTƄ��gAp�<���eNha�-��+�
A����h�<QF�C�@Mh�Lٞ\h&1�e��i�<��I޸^���gĂ�`��� �k�<�2fŻ(X�;R!�<A�6L��f@d�<�U"��B�U����z/���^{�<�ԥ�?m�H���%S_�6X����Q�<Y`�_p�LM���_�Wz�y�b-�M�<��d��Cx~�5� Ae��C�K�<`����쉺��߷���C�<����A�b@�4��92c�{�<��-��q�,��؊9��	Ӌc�<��I
���@�
u�B���Ü[x�LP��%�=�l�C�&����$��yrA;0��e)E㍧EX�Z��΂�'��'��>e���*M���B�C�.�иk��3D��Ȥ)N*%��0jr��gH�p��0��k��8c��̤q���BS�Œ6���ia�"D�Ā2'":EC��ĽY���ħ,D��4m�D�(�t@��:�Ip��+lOH�<r��� �p��B���ر�qF)D�`CQJЮQ[4����){T�U�� )�Iu���5
z`c$폞����J�\���uBd���Ŗ�qC�*N�Y� mDx��h8���C@	;��`Z���]'���5D��6�\L��P���ټ"0*�B %1D�ؘ�!�������%��4Ł+,O�b�������RDâ���$�6@��xb4t��ʧ�zqHD'ŋ+`�D{r�O8rI#��[�U�J��E�zo��i�'�HD�� 7eF�hb�쉠dYT�!w��$�H���)
����/F�z��ّ����RB�I =�堣�7 �-{d�U4e�B��r�{P��l��1�'iF!_�xC�	<eQ %,V`I>�Y���b�d-�����F
D���A,T��VĶ�y�M�9>؝4!J�B�zuy�lO%�y���8\xQt R�?���֮@�ʸ'na{��Bk^�=��2j�Y��Y��y
� 6�f�эu�C,��hK,P�"O*!�P��s X��T$O�_#ɔ�'{�'� `�c߱樫У`tpy8�{r@,\O\�����C̥��@�!^FP����<a�����Yr����W�Z���cW���!�d� dYr8��sH�1����џhE�$;q�,p����G\|lr����yR!�j�,� 2��1>�q���)��d4�S�O��[�*�H`��2��p��G0\O���=yTG9s�2��!΃�UM����S[�'��y"	ŉ�
e�І��x*����j@!�y�i�"Wz]ŃR(u���X�$�6�y	-x�T���HDfb�%) ����hO:���BP���@ {H�q�O�)j!���M1Ԅ�U��qi�d���#(�XMDx"E;�S�T*^�+�QP��v��8��D����=y�'.�I87��������W�`IS�H�\�>7-$��b���~&��A�-X�mQ��։]6�� �2�I&�HO�'yLd�Y2�	��i�B�� $ZX��a�ظ���\,�����+H�	
ڴ��' �>�iaw`� �Č�u	5kRz �g&D���2�C>;ưu����6�P����1ғ�hO�
0�n�K��e^���!dC�	�p8T
�Tfr���ܮC��4�t�Y���m�NM�4f[[;V�<���|�"
�^�����Y"=�b��a
@�<Q�n��^������C6�y�d-\UO���y"S��g�'��Th�CW��zx����P,���'��ݹ�1�&�H��MH���'����BЫ�����<>�c
�'��-�� )�R` 0��88��L��',���$�AY&=�T&Ƒ1�v�	��HO��(q�R�@u�%P�\�WD�Q��"O�{��"��D ����84D��"Ox�'ʹq��跪�
# ���"O`A�;W�b��&Zmp�c$"O~�ذ���A"��Se:��A"O \C��E�~�q��F��}+:�2�"OPZ�ϦD���b%��C�(�PS"O��3�۟4T�u�RA�
_�:1s�"O4-��L�������E�;~r<*!"O��XYx�d졵B��]b���"Ol�"4\hH��T�Y\�8��IjX�Ѐ�,-.�~��#AL�:�VJ:D�� $k�7߼At*�0B[:�)�+D��P�E�<��ȋ�MC�W/0)�C.D�,[���/jY| ���@�@ě��8D���Ț� ��1�;�T�W�!D�Ș�5,����o�7u��QA$D���.������˙4R��z�& ��<I長>���2�1+H�6�Q�<����5[nd�G��07"A	t�K	8��A��D'�O+Hhr�L�[<�u���]�<��ȓ^�� iv�H*[kV؂C��,�����bd���˴:��}���M� bb��I�����pkb�Q� �����
��{�!���n��`B��36�>��g�M=}�!�<C,6�2�M�tL�Z�)ߌH�!�dV0j��2c,��:��<8�L�J#�f�)��9�t'14!R��g�Q�q�/#D��!ӡ��)��@)�v���@n�>!�u6��Xb�ѥ���k����9G���ȓ'5R1�o[�%��}C���#i.̇ȓ7��I��.� +z1C�ΝW�f]��S�? �d"�ɲt���pԅ�����R"Ot���@��d��	�|`9 �"Oʀ�nV
{���Kw(.uq4qqv"O2Q�C�[~�HQ�d(@.#g�L�5"O�w���}(.Q�!D>4X����"OX�AЄ�j���X|* ٩�"O�-�Dƴ=D1�Wo߄���"O���F��'�,('-ݥW_Bp��"O�s�c� .�@ �"SIh�,1�"OvX
�>�:��eE$RQP����b���'k <"�wҦ��3!�4���S	�'w���)f*�(h�Ø�0n���˓�ē3�D�=b��`e�ۙg]z��'�@�z�!�䍉nxt1J@��#�mB��އ~���E�4)A 0�T����S@Zc�LP��y.�!zI�-0r��F�Ƽ���Z�Ը'�a{ҁۮI�.X��#�>� �C�h��y℀�e^������4I��ڧ�7���0>Y���D)��$­���B�s��\�'����i�j��T��m�y�'!n����J�RA�H��m�1�l�j�'�P9b�K��O�Ҭ���H�~�R�'Ǩ���G�"P���3
��a����'v0maPN�8K,�C,���q�ʓQ�����������iΘsrH�ȓds�����Ak��s+A/�����qF\J f�Z��D�/�v%�ȓi1
��&(B�%�8@wL�`FNՅ�5��ɣA��b۞�I;z���	Π��1��y+�d��M�c��ȓ!6u��!�rs���"�L�.m�ȓz�����}�`�Ƀ�	m����ȓb�P�$�ԵW?$��)T� ���vkzp�XP��Ze��r�+8D�Z /RR)���Q�Ac `�p�+D����ǜ�)�Flb0)��+��rc5D��� ��.�@���`��<]Q4D����L���؀�GT�}<�2tI&D������*>��}(!CT�J�����.D����ďe3�̓�?��Mi��-D�Аୁ�C,� ��
�T	�N,D�\�5�:b��,�`
��%E�EO(D���1-�y�Z��ꕍ:���1� D�����ĸ-�8��Ԝ#X�D��o#D�d�IL//=$�U̐�wF@('� D��R�Cn��7gN \�d�5�!D��TEܠD� ��b��b�h�C�;D��������Ԩ�l�&H.DX��9D�����#�Q��/x� �VO=D���kW���H�ISsi���`�;D�T��C�$n:�8��+UC��3g >D��1ӆ@�~��q�� h�1�/:D�H�ېjY�����"7r^x�V#3D�0y�ǘ�!~�	)fk֗BJ6 ��1D��AN��I���^	.$P�4D���kO+O��I�U@OE�N��v�1D��H�	]=	��=;r��"?�H]yt�4D��yȘ#A$Y�HȘ2�%+2D�x �F&��81t۽AO���V�/D�|�e�C2Am(�˶�Z�E�b�J*D��j0EF�@�b�����XG�fj���B�������y�b����+_�:B�ɘ)vԀ��Π5�~��5�S�8B�	w�䣶�W�?�Vy�b�3=)`C�)� T�"��{O��o����m"O���!(��R��dQ�K��ي�"O��(%�3���t�q^P�v"O���CH˾@��e᎕�Nhzmɐ"O��j�.�ш�B�m�
Z�����"O4=x���5}t��t�q���"O�$�ge��;%�z B�
����"O�qiנ¹ X0�a�s,����"O$9����0���bp�>G��p��"Ot$�D@laaK ͚#� |�"OBD���,h�x�����\�^��""OLm@��)$	Q'Sq��#"O���w�]�^�1�қuN�0"Ox+P(�6O�
A��'`�Q@"OJ!�e���B�z}QGhR3Ohݺ�"O���`�X%V+V�pU�N/��A�"O���Ԉ�馽a@$Øy�Э�$"O���͝e�!���x@-��"Oz<*�-G�2�Ɓ���-o��� "O8�p4 �3lt&]�g�۰�Ġb"O&�Q/��Z}��Y�KL��yb�Y#IW��7#�>��`���yr�R�"�YH�f��)�x#4���y"MY�]�FH0���#�blBd����yoQ�����J�{�hm�d�!�dS�+`(�K���y�40�A�H�!�ď�������� \R�{!�f"(2�l7c�xE��Ú�c!���uM1�B�7'pE�1��"kU!�U���A��:a	��Y#��PyB�C�o������1w�b�]��y"��=>&�BV�+p%�0�!/���y�E�"{l�@�.b:����0�y�X'V��"�"�]j��!��4�yR�X�srx124-�b[4� �A��yB̝H��ֈ�5��h�� �y�D�s.ĸ-���9����yBĚ�2�-�'!�J�VYR����yB���"��A�foNy^A�(��y�C1Nu�� G�z ^iq��y� �,V��T��ak���#�)8�C�I�?�
9`���Jl&�1��D;ZXC�I�d�2Ģ�4*��� ���Y�.C䉱~F�rbU271���c�9w�B�ɠj�Q����Y�4����n��B�	<��b�P&$� ���+��hC�I�#NL�Ǖ*9�5��eЅ�nC�I4�L��k�)T؜�
;�`C��/$��|HqL��O�԰X�!cłC䉲N�����M<_ijm���lZ7�:�h�@O9�أ��Ҁ���x��'D��RO�PI�3�[�@Yr�e�!D�DK1�4X�.�:�/h�B�2�:D��C��O�P�0D#�mLm)�=��l�A���Y��^aK -ۦ�ͷ��C�$6��WA�o�� �i_�f��C�I���)�3
׏ay�%�`��5�~Y����s�:�B�A�\�Ѷ�ܸ3� 򓤨��0@1�Y�"�ȼ���.W�Y�r"O$|�2Ô�F5�@��H�#ZF@dQ���M�ON�P��Hқ1�$k�6h�2��'�n��4�'�iå/ϼJ��T+�'v�ꦣ�V��ł9��Ii�'R����h[������N)D*`h���� f� q�U��։ۅ/�72s��8�"Oh� g䇘�����]q��;�"O(��d�1l��D(��$4If`d"O@m�Gg�T6��I��5t/�a��"O�i���E��e��JnH "�mX���p���g���OU4F�� 4�>D�XCE�Ӹw	�����fq腮8D�d�O�0a^Q�v �K�^I���5D�0 i�6$�S��+%�ٓU�-D�dP��CvjM�Ҥ�d����Q*8�k�T�OW:o��yJ=�v�V�z�J�I�"O�R��k��ܫ�A^
� a�"O��J ��ph�`�
�.��r"Ovm�#J��8R�)8�K.&���"O��2֩��t�i٤`��!�B��"O��v�2F�T}����:���""O ��`Ô�_7Lt�2���"OL���c��G�������B��C5"Oh-�`����%)	P�=�&"O��a�L�>�D}pHڈq8X8��"O�h;ucʹe�ެ�%�@�*���"O�,q�B�j�D`!5�	z���0���$�S�Ӆ1Nj8��Џ��E� =fC��*�:�T�y����J �	�:C��<��H�k�$�Hɥ@�p�8C�	�[�pa��j4CF�)᫞�MN�B�ɬJ)�@ 4G�>i�PS�NЛ/vNC�Ɋw������MC�����9:/NC��>���@��Wd�p�q�0�I�LG{���IǷn���JB _��zM�P���M��' `A�&�ۀ��T��Z�'P8`Б�!��c�JאL�(�OX��oӐ��Sȑ{�8�̀]$X1�&"O���p��$2���W+ݵ����Z����'���0�'΍e���'ʙ�f"P��'7��C�Ň�3�|`�&�\_9>���'���C4�F�5�p�f��S�`���*,O��� W���H7�7]� y�"O��'�5[�>�����9�谶"O^����(�Vtr���>	��1w"O��f��Lo������cN`��"O
	�1��4)->�iW��:<y"O5b���/?شz7�!+J�!""O=���	n�h��0� �t"Oޝ�hV�w�1���5]	��æ"O�!�
O�Jӎ���GR�R��S#"O�*�j�B�d�a�̖(Uz��:�"O��bH�w\J]��׵b`���7"O�pQ]
�%�6�>$M�*�B�I�ޡ�r�L*t��` �*
��B�	�R\������9܀\so�5Pg�B�	%jL���`f�NR��B�M[�C��)���N"
��YT��jX�B�	:$.Гtc�+t 	M#��R���	Ǽ^
��'EDv!�D�3g�JPx�J#\v�`�e�a�!�L\�:�(� ݟsR�}�6$	�7�!�D�>��Ed�E!B����:GV!���N�D�eCצ/l���]aP!�d��=t��hS��!A�1�lJ�e�!�dD.D�,��! V�K��c�$$�!򤔯v�H�#ɚ%V4�ʅ�2�!�D�k�ĹhR�"Y������7���I��H�����쀅g�b��"`���L|��"O� 9qC�>b���8�H�=o��\jW�Jx�(S��'�|Ź�͈x��GM)�e���)���Ui�9l��(���!<�L�ȓxg�L�3�4�T�'��s��9��z�,���ܚI��4K��2B����Ib�'ev�8W��o�
��+Z�0̺ش�Px"�ۥ6w�9�b�N��IvmO��y�7<��@�Bm�l*ǥ���y"f��t墐A!!*bbL��g�ޔ�y����ez�TbdGЮ&^�3��W8�y�JC�j\���f+��ps�L$�yR�O0k_t��ffŽ�Ҙ�5��1�?��'�$��7�I(`Y�i�a� }�)Oġ����,�� �!οA9�\���T�^�LB��ej"hy&��)0�^�v�dc�P���S"���
*T&\t��)EH��į<Q�'J
 �H4IR�b���J��g�<��)�Z�Q���? �Bq�]f�<�� h �5i^�7>t8��ba�<	3`W�{kL���X-�t�8�I�]yҘ��$����͉^�|��A�S}~$�Ӂ�?q!�2����S�{�����_�b]!�$P�+��3TA� �5����b<O�$�$Gߢ@>-� �ӄCYf%!%"O�|I���dz�J�,�A"��
�ȟ��KdC�
]]��J��aD��C"O���M�ql�ь�3b�p�g6O�)�����s��i��-��.
� ݒB�I�EW��[�4F`{`�F�[vB䉠)�l��ԁ�U��{�@?=z�B�%=`|hÁ�oΔ�z`�.yhB䉓����.��<z���@4C�I=k��0jU��6#��1����B�	��@2u�V�o~>e��(�wZB�I(F�e��Ɠ%OXP��H��B�I,P�I�%(	�Bv\�uk߃�C�I&2�p�3s�	�y��Y��|
�C�	���SQ�ĆH0����&�V�rC�I�pj8�`UBO(#X��xeEZpKB�	�*��`aN
o�Z�A�*�?*�&C䉇9����⋼<R���VnC䉔h����L�)$]ʥ�:f�B�	�QE�-:���p�\\i�� s�C�ɮNmf]��"b�.,����y�"B�	�?����f���0@  K 
��C�	/�B�y�Á#P�� �Gs��C�+<ц�7ȨY���I$g�9�C䉼o���y�bǛ-��u:2���dC�Iaݠ�r���#�,XZ��$^kB�ɮp9�(�0�ά_�HC���/�PB䉄%��y�!N�T�"��B��0a�찛5A��x̠l޾w�6C䉟��xvFDF��u���N6 1C�ɞw��P¢닚�va�	T'C䉮G
���E��I��耔"�9��C��+
�`�d���hn��e�}a�B��:,EF�(U�'_�$x��^� �B�	4�(EI�� ���PFFۛ#��B�	�<h0Ej�H�AS��Y�N��B�ɢ_L[A�Пn�DT/E�nrB�ɧt��uiX��t��*���pB�ɪ(-t�Re�	>��A�>e�PB䉩P����U�lNE趁��TC�I�`FzA�I���%22�F��zC�)� ���k�16Ĩ�1��,+�R�x�"O4��p�٢	F�!
��կ��2d"O�hi*��No��س���D�	�"OT\�5���>JHt`N]1H�p�ZE�^��Sd�4��)�4�*^J�?�� ��xV����A8$:J�Q�<i��W�e1�M;����p�Hh�+�O�<�tH�B��Ȃ 萾Hnq�!�H�<�d��*�:ٹb+�"`|�!�v`�F�<a�	��娧F̶�t�[FJ�X�<�`A�&~R����@���「PX�<���ÖZ�h����+y&ʷ/EU�<)p#�%���A�M�9`p���+ZX�<��/�g���9ǏP+e(�-y��	T�<�@`W(I���u��0@u��	PT�<��$ۨ$�t���9["��hp(GP�<�@d�!��E��#H3�Bdp�@L�<�O�>���R �&��#��N�<Y���3@�B�HS��4WUf����@A�<�_�'X2���:n=C5�P�<��I��Jh��[)j�X�����H�<�d@�<)S(N_��█]K�<y%
ѺC�h�I$�-�䡪R�Fl�<���l"��$b�+~���7�j�<�REʌW.�m�! N&����b�g�<�����0�����e�l�PU�E�<i��ln����kp�xT�TF�<IE�!��,��6
E���F�<�P�E>@�z���
��mPrX�<q$�ν ���R��2 xgˁZ�<��K��i��L*�g�x�$�#��NW�<�B�T�z��x�a�X"/L~$��TL�<٤I�T����!�֢4��A�KNc�<	� ʍ�f��`�-�4P��r�<i���#6v�(�,^,R(�ţƖa�<cEّ0�T�QF��!b:�UC�]�<��4w����kJ��t��
�@�<I¥�W\����,I&��h
Y�<��eX�6h<���u%,����B�<q�o�9T�\�3�
9M������z�<Q!��D�L�ٷ�1 (r���Gx�<����r�%�$f��[�A�_�<��!|���%G^=2֌\�$*ST�<ɱ&�$k�D�8�eH=t�@�(c,�o�<��ɬ5h�rgE_4$�8�ǎ~�<y��g2��#1GY4
k<��vǚw�<QQ˘�d�D+	J�B9*� �e�<�s��
_��Y3Dj��O�y��E�<�Q�K��r�"�oI� _hx�no�<�tc��n	D��%�C�l�\A�R�<�v�0~�T�b'_��ƌ��i�V�<9��(,�|y�3CW�b�J��b!BPX��2ǅ!��P��9X(zirQ��2Kl��S��Z��j���'>Ե/,2�����::(C0!J@�'���.]�q(:�Ѡ�͸��'es��l}��놊X�����x��J$z':I{kC�ˀ�Q���]��Y�b�$�<Tё�鈟�˽h@�f��N�x JF�.R2!�d�u�)#!b�L� �Q��PPޕ�q��3%���D���6J 9��ϨO"-��P�����H�$�� 	E�'��k�ӓ$��`�/لq���@�%�q���%A��Z�iP'�Hf^�����+q�Y)���M�Th��7r�O�0���7������E�KM�N�'YY���ԭ·cݦ0�3B�M�ȓSr�e'J�ef6-��`R-�e�[{��0�ƒ�=�Dp�铺�y�)��l�0ԣvF�#�}�>�yҍ]Y[�d�QG�(l��ĸ� ��4��ݠՅ�xʴ�&ˋ\ � [w3l#>� �h��i̋WS��#��$$����'slM��������#�1Ϣ8򡈞-o����up΀���DE6����pMN0  H�`Ma0Lѿo�c�s�[�x�Q�`A�'Zf0�EE��D��Ӕs 48�%7m�|��F��{%�C�I����B�	T�m��|��G>hL���ܯq�V����46`n��&����Ҕ̻b+(��̈k�T����.ݸ�ȓ��LcC��O3~�Bc�۪D��y�!��56Q�q��Ö�0��2��ź���(O�P�U۰���+����x �'�� �I��z�A��1x�y�&B����._� �Tr3��sg,����>�O�X���1x���S�\�]C��I6j�� j��+f��\K�K�%m��q��	�?%�v��G"`:�-?�I;e�%D�X� R�P��t@�'�%i��,	0 ��
$�:u
�1u|d����`D�@�����Ͽ�@�Ctxl�G�B�����p�<�c�BR\��R[%�T�B�]�8�>���+Q��b���*[ƹ�Oc�M��Bo�bTQ�K�e�a�C*�a}2�W/zq�2�P�/���a��"R<Dڄ@�!Z�x���ΟM8�b�%åO+��
4��D(Ꜿ0ٔ����Q\Ǒ��&�Ec{<(s���k���	eH��gCZ�a���ikt]�g	�#`��0�d���y"�Ρt���@�W�\�֬�[8�M+Ԯ����`��Ac��AF�ؕ���ư���^�,�͙��raL�z�"O�uIᐒwHiXP![�'n��h���C�����y��	��Ӈ9�:�(O-��HB-�2h�U��?�L��g`���6ъ	�_��)�{�Dz:�ń$��Gۨ6&�'p���P��M��51PT��kƈ{��d�O<��*_��h��M�K~b�H�j\5}Q��Fzb��,�x�%��9�r��N[=._vI��2O��南$
X`@�kV�A@)�I>;R�ha� E6�b!������В��N���:L���3�i[���U	�~k
M����\s�{L�]�����\c����O��`����[� 0	��K���DӼ<�4�2t@�1<[�3|��{D�=þ=١�?��]�w��8QMp����[�܋��W�4�ݟb؎��Ş�o�����~'�E!0J�$v�;�A�H�D<��az�@V�K%��3-B�T�nE,���P蒧r����UÂ.P�tyT剃�8]j����\6$�2uo�E_���%�yB3��,`I�?�|�A�O�^Т�����*�r�'.1�N��&�7�,(`
Ӵ!?fE�"�5je�X�U��Q3�Cօ(��Px�×�D���C��'<`MD�ܴ,Kf�Rp)��?�8����i����J���)t@,^g~y�`�"<\ؤ��C��M|"�Rd
�h�7Mg�-��,@�`�����T�U��F��+�H��HO��HV#����1ME���r�b(����bQ\��	�t$�-܉O���+�I�xQ�!�al�R���*@�J�Z�D	�ȅ:���y�꟮ �}���i��d�CC��(ؐC��|W���aښD�(pI�KL2��� i��)+�A�� � �'_���!�'N�z�!č]��,x��O�
�򤃈�@9`��
��)�!+Q�Z<!�HC�9�~�֌�	5��I5�D�c�2ۃliĘ�x�j�ON�ȃ����MSP��'��A�C: 	uph��ɺiHqhN� Π��B�<�,�C��P���n�/�*%C�b���A2Sm��p0)4Mҳ$)�M�� _%0�a@a*A�.-S��	�"�<���<}������f]p����������eR��q)�"�0����=����fd�U�u!�
.���ADNܒdrR�(��?�;P쏝G��=Q��'wq/8��W�Z�&c�0��G� �4H�Ȏ���#��K�	v&xx�̀���4( oZ�%d�� �B��
(x�|�ȹYFmǗht���@�<y�,�++��:�/@��@\�p��
�X�H`i�'�p�m1:�h�i���0:b��
!���6#��N�p �!&��H��ܞn64�l�,k�\��C���m��x�HOl��T�/�n�p�L?<Hp�c>H�d�2ϗP�	G�CJ�x�3%֠0�BL2���q,L�t� S��"4�ZxZQ)
t(����:N�,8Z�DT-ÄL��I7����(C 2BZ9�¬	�-�E����;L�"
c$��(Ȓd��)Q7� ���(�d�DI0�L+K;��{q��/
��2f�U�7�¤��_��"tN�	�F$�X.̼��LߘD��ɠH�B�-����]���Y���&
�OKd�pc�V�zn��§X-iƈ`c�AX�Q/���z6�	�#ېe��#t�^�I�e��%�n��w�����EB�'E�d��R#�qzGJI:V4HD�G<iHB��%r���ȓ��#N�X��$�&�]� '�t��5; �U<.�G���<AGϝ��V��2@��w�V����s��	C�L�+��Z׎U
{{
Y+�R� �bh��d��|�"!4!8y`�ǵ_��E0�)$+eS�@��X��瘀E��2�_�|��{7M�=p�5 ��"��ቧ�]�q��u�S��@��i�8W�_ƺS,�{�0+��ZۑJ�-|�L,�G珱f���S����V�`�S�B�<Qjny�Ԉ4�"��"��)Z�]3�f�!H�x�l2?�F�M,-A�.�ں�g%��Z��öj��*Qv@�aG�q�bx�U�G[��p��DuW�~��HGK�rMD�d��p^h|�Q��V�:p�� P3fJ6��`N q�.tqEꃷ>-K���П2׎�P�$L����bC 1���w�4@�f� Xp�`�	@g:x��
�fn��uǐ�2��v#�F���	&�Z�_�c遈`5f�zt��bf�=��^�5���0�fՑX���s�풗�?I#Hʊgb@1����2�0E!5��=0���h��An0�j���K�Ƽ��DD(�4i4�R�r��5���̊�M;"�iA����'.�
�"C���TdQ�6�>�S���Z�8��gR�E�hQ
�IB�B��,�u�C�'��T�!��Ll� tm3B��[̰�2S��a�A�EW6�MS1��<qs�1�Ț�!��a�'b�M�E-ɞ�ڨ��̚�AH ����8�ȤEx2�70؁)�X�.��tj��Pz�!C��ޠҐAE$�D��W��#sبIbm�@h�Q.E)y��E(���c�Q������O�0@�ust����H��Bw6-�#�ݣOd�i+nH�I�>�	G���>9���5�t��40� @��8A��,��]8x���'ᕎ>$�1���f?�ʓT>�t�PG� ƌɐ㮟�o#�YX��dX@���̙.����׻Cw�ը0eE��Ƅ�rJ
�s�|��ٌ	UX�ːL�-���CW�8G|����圢{W��h%�s��!H��C��҇Ŝ3Xl����8u�8�.Ȣx�ջ�¤czz$0G���qF鏶�&T
&�F {���!f��P�&g| ���_ܓ4\8A�L�C��'�rl�>9�bI�4�� �7b8�GB�@)��1C�GXp�Gg<+�6h��י�;�JĤ|q$����t��1O[y≅+9��R��_5tN���o�Z5p��5
1~%�5&`�Z���c�X�^�i���^h�1f�UX3~��E�ԝ2y҅Fڒe�D���c;ƒ qd�ǕJb�@���?�t`�s	�Fz�4*;N�KA�ƅ>̂<YT�'�=\Q��oZ����$(L{��J�#�$o��]�P�@Db���Gή6He�oږ��a��Jw��b�c�%Nu� ���� ؙ�KȦA�b,����:�0R i�'G��e�H��� �i��h��ÿM\�]Z@CE�u&D�`V��H4��٤7R(Ig��d�~5��$��NU�e:�c�s%@�P�'2����L	��9ǧ�jHH� �yr��i@\�x�����Ը�qAIp��ġ^w=J� 6�Fo�j��G�mD��",�5� ����|y���F�Q*ɰY	ïm�h�InB��B�Z6�(��^wJuᕃX9xS<��'Ӭk��Et�U�X4��뇥+?v<ъ�L_5��':r4ݚ���4A
Be��$�/]�8i��o���B�D�@D���匒�y�I�@B�x���._�3�	�"hN�+�j�G4�{d��;�,$�:W�����B=cH���!lD�cu�QI,�	�8�$�]�"j��ZBd_�5���ҭR7Z&J�prƊ,#O�ii��!�,i)0��&i�R��qTڼX�IZ%���k�I�y$�b����hOi�&��7y��QJ�^����_���]O�L�KA��[�1OH�{1�]�V	y1�2~֍���i0H�p}�׎G}�"�"TN��7���� �ja��H]�dF�1F�;� L{q�'LC�I��FĴ9���	@`6\Z]��dܵXh�&P���	S���QO�p��U8��ة��%Q��&�@�Ʌ���R��>�3�C{�y�.ݚ7�p�Z�nʼb��})�g\j���1�/�,6��#������S�ıF<pE�co�4����8AD\03tCV�9�9Dyo�7� 9��BBT<��� Q��q�n[*��Y"#T���OF��C$Y9i�(�I�z�d)�Z�f߯9��S��� f4d�>�Yߜ�p��|�>�Bw�B6KjR�##�	O��9í:}bHF92�H�f�4Z�ʢ~"fʍ)o����@
�:�@E��ٍc�Ԉ�&��g��h��	�bVT25`�:��=[I�抅h���q�,���L<�Q�ݔb�`ת�&%<�]��@�<q0&��p��`Z��'Q���'g��@"�/�kΉ�@�9}�ljf)�Ox��M�(	�>�y� Ѳ_S��z�'�q�(�/��D�#C��A��i��"��A$Ak!�$��"�f�r�֏{��Q;�.Ӣ/F!���,ӄő%o�h,���֭\�!�A$<z��eeҏn�0eY��P�'!�d�#z���E РW�@Y�ʗo�!��Q;W˸x�d�4I�/͐E���m�x�� �53��h'��JB�ɟOW>�#���Z���	AY[�.B��f�}qE�R�42v�K���(*Q�C�ɖ���:�d��8D0k2��q�C�I�eM�]8wDH�*�:�z���=��C�	�Y����n
bf��C���C�/v3@D��A5V���u�c��B�I�eP����=v����Qd�XB�(U�PX`��/-�i���CN�FC�Ʌ~x֍�d�v�F�xo�)%zC�}<V!AŠZ�moX1�L�<КB�=Uh����0}f�|���&XB�I�PX:�8R%�cF3&�R�؞C�d*(i�w�Ϗ}�p]�b�W/nlC䉮b/�U�/ߠ/} =�vH�)^�BC�IQ�J��#�W�p�����1\�C�I�t��yI��5 ���ɒ�W-�C�=v�r��E��y�J�d�бK�B�I<��K�A
D�T�`�Cؠ!X�B䉣n���H�g��w�����Y|��C�I�I��dN��i�dA�GH6o�\C��D�8ȹ���v�l=�ƫn,C�)� ��y�D�Nyh��U*MV�I"O� /��� 0�W�	в���"O6q���	K��j�����""Ob�R���#U�ʝ��S�m���AA"O�(�Ą��x�X���:@�J�"O
� �H��^Z��b���U-�|�#"O��Q��ŢT�R�����4rFl�u"O�z��"�4�˱Ù2k�h@q"OlA��5c2PT��Lf���A"O�QA�k��)זl���քwB:�C�"O�RWo^���V%F;��"O��˜2´��k"��� �"O�Dc�H5h|l��K�3j�z=�"OΕ�h;h�0P)Ωm`�0�W"O��3�OƸK���� ⍽b�8`�'"O���4au�P�1bp��)Z�"On�9�C�4�d�RUhE���q"ODu�Q�زgQsG�p�y�"O���e�/$��P�;e8�r�"O�8rT! 1
��/�z���j "O�mB&���x��]`������S"O�(�c��.4��(Ӊ��4a�"O�]���P��S�7&�-I��[��y2B� v������&}�h9z碑)�yR�C._6b�GC�wV|��ʓ��y�!��(`�E*u�����C���y"��Dڊ�{�� joR�P���yBh�"Z`$1q�<`��pˀ�E0�y���fg���'���Oô����Z<�y"���t1���,O�>�1 &C��ybo|�!�G�
D%���n��y��̥s�,�e@�t��E@M��y�+7��8�4%��>�R�*u�Յ�y�AJ�u�"��b��*�Q��@� �Py�G�X��ڣ׽M�����\m�<�5�ưf�4lR��@:��SgFc�<ဏ� 8�!� _���Hs�<�g�o7.+��I4V(�@�B)h�<�5jݢ%x0r�I3:�ެ�1e�j�<a���#�z�y�*ʆL4
�����n�<)df
����X�n�c�N��e��}�<����5�~�[�a�=ͦ���~�<�3��*s��g�	�Id�e� �f�<��ٸ[T>�� +ݲ{�DM�2b�T�<��b:~1'Y�[cV
D��R�<m��;�*U��
0zB:�m���ybO��μ����M�:q)\�yr!
G��+SK�~�0]3��'�yb S�-�t�a�ܛh�f|��!Z-�y�%|墜B�E��as�ؙ�M���y��D�l=dP�˄a�}q6�J�yR�&r��X����LEX�g� �y�"M��PHH�O�M�d��5� �y�&C9w�� �R�@=N*��#hQ��y�bB�P�Bu�ܸG�~)*2��>YD$�+�\�ah �]q�I)GP@�bd�h�8��Oj���ۜ
��� "�TMN�s��ɼF�b�2�۝���b'��X5b(��(6K|���J-�!�Ď
\���6υp�����hɺ.��$��E؏m�D8wmN.
���o:��<�!�/>$���h�3!�@�K�+�k�<A��-,�D����%v�(#�ȏ"6���b�(�A�gH�A��0�3�wy��c��\�<�D��̅�F��l!rC=��Cd/�4޴a��hE9HBtx[փ�72��r���&�0?Y0E�7���2G��jZ��" ƃP�c���� �U�x`'��})֛?� ���+*kѾ�9��/w�J�y�"O
�@P(�y��P�ɒ@8\*Ri@� ��4��M�(e�QA�!��>��'t���"��:��B'g�	E��H�')�U�"�ͨ$l�ɆjזRU{�ݔ+�Ш�k�hQqန7�uw�*�3��.юJ1�[��D>N|�E��	�`�ܹ�i75x�C�U�Ai�����X��A���#@ByRD���0?�%�pG0;e��8�1��D[�l��ba�׻[�)��x�����|�6�DD$��R��(��,SW�<ɔ��� 5dՁ�HFjİ�ȋN>z!S�#��}�~Xٖl�;��tд�ӗ�yG
586h�z��� ��R�k\��yb�H�rB U%`�,}��Q�����w��� '�U��m^6@U2_w8�1$剪2��h������aG�������.3x�� -�(7τ�1k�);2�B�'~xKL�����2�?R"v���Z��9�Vo	)/� �%�C��0�#�Ѵu,+VM�TUPY@KA�8�]��s��zB ��R���[sҒ>��B� -
x��7n̙D��(U���b�t	��ָ$�T��LKkV!.p�Џ���)3&��d
"]�$�҇f�%a�q�ȓK�HX���ˑm�.��Ъ0�Q�T�ŗ{^����ӫ$�rC��F��7V�qO�����ֻ�~ͫ%h���D���'+0����5|RH��'#�0䱣��ڱyxa�1dx=�< �c_�N����g0LO�|�ǎ0#ϼ=��+�/,����ɆEh0����Y`� ��,�	��L8�F�8<���Q��'�ByAp-N�jm��'�&UHq�r^|Ԩ�̚
Q6��H۴-B<��nJ��e+�*�d�}� ��?江k�_�X`� �+�:9�Q��	ȆvH!�D�w�<p� A[�"A	R�A�oz�	�+B������'� 胖Q?A��M�Ƙ'|�� 
);�=��0>�P��7dp�� @�\}��;{rZ�G�=U1�/$*�V��Gǖ"Pt�s5�'��d ��6��HP3��`X4ڌ��ѧlk ,S�BR_>�qf�7!I¦�àR�ѦX�\�r� ���3}�T8�'	�Y�b-S�"��e�R�U����شT�yJ�Z�?��}�j�<Y���ś�A��|�1�iW�^���7�:` }�ȓ(����
��(���C+ �>��"n^�,�4��bKmq�F�a��i��j##O/��I����B�s�VXS$X�V���d��	P��y 蚬a�(i2��#X`�F�*�"��ӥT�
P���bʰr,)O���@loBpf�m}��"���.��O����/°1�Y�(�����ؐ
��ސ9ĝ�4U#��R�cM(����D��=�$���$�:���@�y���%]u�q�Om
|�CЯ�~R�
�����|��UBC����&"��\��1�"Obx�
��	+��P�Aͽ;����Q�Ǵ���@ �ȓ���(n�O8��W�2P4�ā�V��\�3�F;�F�k��E$L^!񄕦���� �$iCR���nɺ-���0�OH.�a����:; �"�����b ��nNH��3�xr�.V����K&��Q��CY���<Y3�/D=�PC�1��#r�5F�0��ᒪ}Nhi�F&��q3d��<,����*lhb�O2T�b��	4}Sz��q'�9"��A�P��'0��`��T����d�Q�CO�a�Q��F��H��*�q�5!�D�P��`�+1(����0O`� �M e�n	��j\[�'k2!2/�	#>pK�"D�~9(Px���$�����43%X��C�fh0!	O�'6`k�Bċ:$D`���"�X�;��5U���� 9o���[mE9 h�MKE�'��2y�3¦H?"@,�P �X
�k �3'g��k�䃉!Vٕ`��y��f�>&I:�0 �\�uI�-%+n�c&
(U뢨�4�3,O� �L��U��i9W�I$)栙�E���A��Pe��d.�I�!Y]Hb䬀�]�d1�f�B����E�%D���p��c �qd��Z[�fi�+|�X҅
+���5��#R��k��[2m�6�J�eΒD�lY���qŨ�-Ҭ_���1}���r$<[��;��A�pT)��̭-O`�ӵ��2��Y���U�'����sn	\�%�T�
#x  �%�/;蘭��	�HZ����Zbg�ϻd/fm"$��.�慀P��q��!��D�Nt:��}����$�W�t� �/D�Ұ=a�╏;y�1�(��C���[4�h�3�Ѵ����M�0%3�e�%#�'<�F���4��~�x�@r)��E�`���+|6�Yf�S��p�{V�	3���FX�H�0��������\��`��fO�~���'ә��-����:b�ڡ�K�#|"�AQO �
|�ӆ�*u��bRǒ��*w�5��`{�o�>�&���<)��̶e���s�L�26��1Q��Q���\�ٽ�4!C��vle�Ԟ.�褒���K�|m����
wNű�HO�_���D(�!�����(��Fx�l�,�M{�눾{,N�u � Ǩܰ 7A����W�Ղ_�8��(�y�'�DQP�x�Q�6��5\�³-Q&@�!i�l	h<�Y���?�aF~boI�f�D\��� h�ḇ�l�_Olpf��<�R�F�ƜZ���Ք�� d�^��u�`��(�LF"p�X�-�@,��q+�2Z/^u��/ۚ~�ֵDy�}����ǜ.y�~� e�=kf��#'��*q,}����9�x�q�`*6)�̱��R'����ϗt
�r�h<Y�aI�>�f�)g@Ϩ0&���F ��� ��u�`.�807dN�V���C/��]��`Hv�LuN�� �KП<�
���iʇg!�HǄ�Q� ���/�.Y�|  g�!�v�P�N�KB�4c�'pn�c2V��Ra�ċ�6�b8x��9$���P�A�n:���b�["��<J��a��!��a�iI@7��n|� �vzl֞�&�$���ě11�\|h�M�
W��(��ƔR��({�) ��m�0%8�a�����[�㿳EO�}��TC��O�\����C[�@7�R�hj�d�2d�c㋟*6�:y�����H�&׾Vkʴ�tC�	c$���U�֙}��Z��^ͬ�1G	G�VxsG[.5�8�u�q�p�: #�,~��I᳁&?9�����,9���ܖ;^h�Ov�Ϙ�.q ��T�=y�Ũ��M]:%9�m��E��J7�?c��e��L ���+s^��k6h^#HW,	Q�d�p)Z%K9x�
�[t	
$#�`q�%!<3�JLy)�qi\L�(O��
qeA�"tʁ)�I�^xU8DO,X�<x����V'<Q�a��2=�����B�~3tC�Š1�s��?_�"L�G��U!0I���۱;��͛�	æt!�tz� ��Ec֡I��9B�Q ��$ ��bT�Z�'�ҴP��]#	�6�+q�S>(��\�Ť�@s����f\�z��2ȷ_D� KD'H;n�UbA��.��H�դ��FvqOj��K�4��	���&L�&(˗�$�1�����ү.�.�[�K"�<	���_<�$�F���'\l����#@R�KV!f��1rE�Zb�@�$d��'ƭT���N�b�b���<v�a�����L;T�MvM� gX4�Ec��7DJ�)��W�u�y#�L�6��PԄ��`i����4�|��W�S�J#�Ђ��̡^�>�C��*~u<y��'���u�B�S�j��'�&�O�q� ��!(�Z6CP�N�6�P�j�4*����C*a:�D)���-!S��# �b�c�I�,�pʘ�5�@�]�bI�2R*C���V�Ȗyv�a"��,��<���إP� B�M+��\ ��O���IC痓(s�t��Q�J���6pv5��L�:>rqx`�!���gV,|�x��cw�8:0D��(x>�Z�.3fc�|xb"6�I�gf�\(�B� Ln��2�R(Q�,)C&mݝ�Ũ@\B`x���#�\a���A(#�:5�ʪ%¡�&H�XȢB�"UGh`��'�Py���+%� Dfݡ`cM��w0|3A�_=PlX��S�3�.������q�F2����+AEƁE
:�@#͓�U���� c�č�f�sy��Z2tL�I�jPntcGǑ�Wº��Ϙ'O��C\$A�n" ���Z���K�X=0�qjT���x��k_�7O��#c��G�t�<٥�\ۼk�K� �|l�'O�0�R�� N�2��rஆ�z��Gxr2c%<�
e�]�1ozIdi!F"��[N%c��iC���9��z퉈'�X�K�)ٮn��-n�����M�B��8�'eh�h�'-�gn�0`�L�r�HaT�"py�c>�J4�!]����B��("�(�1�F7?�ET<UO�m���,V��iE�Iʖ50����LDy��L!aO�U��@����Tع��m� ����3?cͅ.
	�L��>/0�ɱ����7�J̚��L�<�B_�bҝ�|�<�EN�:�(�D�7sd�i3sM��!^�l���̀N�|Us7��2֑���n_���5Ƌ+(9����*�)���t�N\h����c��(O������.���N�]6Ԡ�W+C>o�d]��"�}��KD�	-��}�則H���dq���I,~
1�s`A�==�=��!,��pK�e8�C'z�l�9��I�+�>`�%��~P��fM�bJ�`�G��Yg؈q��+����U��FQ�� ���+ q�2̛>l�`�����$8�g?�E��T�U�`�fa��%�)��8V�I�K ,8��L<��T�u9t�����{#�*@D�<Q��`M��'�';-��oӠY���d�O�^cx��h"�>�J/�O&�C�/TlT��J?hWƵ���'+��"�_4���Y�n�eeކv�(���Eˑ^r!�D�Yq�͢S�]�M@$��c�I+F�!�	s�@��!_?���U�!���7�B=8�Oك_��c�f�!�D3W(D1u �.�����b�!�$�hޢ������h�Lq�!��F�&-�Vتx�*tT�P<)�!��U����B(� U�İ�$�ݣ,�!�d)�.�[#"�b)��.!��[�#��0,\(n^L�Ń��|!�$H��έ0"�3!Sz�Z#�"0
!�$�	I���a�O1{n�pA���!�$���:}�Kw	�a�S_"t��'MV�2q!]�=��iCq�����H��'�(�jbƐb�}�P��x�:� �'O�����-T�d h�)�t���2�'���fK�>O���@�4��a��'�L5��GJ�9pȉP�O
�x��a*�'^d�! $�t[�ͳ�LN�Agƅ0�'9�\`ALūI�v��4iØI봰��'(�Z�e��%
	��K�T܃�'�H�w��k� X�����'U�[��#mz���wh�/C���'cR(�C�4U�|��!Ƙ׈����� ��wJ>u"� �?8V�q "Or��a� D��ٙ"��T�"O�UYb�>V�2���ݺ��h�2"Oj�ڗ�.Ix��
��W���*�*O:�RB�շr#��"�h�Oc�`I�'ih�`�IS�GT��CUN@,=eZ�c�'��yx�C̬�8�M� 2;,���'� �H��S]��=
�N�&-� ���'��GH�j*f`��aža��'ixHcl�P�w���!"��'��`�  +��hD�1���	�'J��2�Y��PB��ռe��	�T�N͈`��"���q�-��+E����3%P�u0�|Z'F��.�tN��:R 1�?�O��>up��!�y��	�6�b����&�h(��e>A	��S�� ������i�dD@.>�I�=�蠁O vHD���֝wܧ]�n�� '�E���S��\���5�ƈs0�S�h;Α� P���v�:EHU��>?���2�% �&�i�4����g�X�`Ź ��|����^����fO��B�FL���T��m镪��m�f| DL��p�8�)�'Bp��q5�H�X�a��<P�*g�WR������'�$o>q�a�īL�,}*���9�����AX��H�¤�'�y�^�������ޑ����I6��"���*�5b��]�<�t#��~��ʡ�u�kR�4�eÆŞ�=�8�[�h��'��ֻir�9�W�~�	�NE�'W��H��*��njl=:�GU�2�O��Γ2�Σ<�����@+�.-(	��ҭ=^�<�g[��K���6��^��V:I� h�S���,�=��ddD��O�`�0̑���;�n�=h�-J�ue<�Y�c	/]Fy��|J NY���lK�C�0������0��Ob05��,G��i0PƮH18���2�@t{��aL<q�E
�6�~�+O|�ѕd��� �B�B�,�*X��(���)qO�>��d�CNеsQ�Ð\{�Ua�s��u���A:������u�t0=Jj@�#�F�+:��3n�	Of�ۋ
�'(�z��!L�"Z�4��*�j�����R����O�(d!ȱn,'��{�o՛z䀓O��s�O�[�Sܧ?oZlʃ䓸C�aE�([`a�'��ʠH��Mk�U��Iʟ΄��X���a�IV�]�f zm��5.nD�R�]3���1j^؈�V(�d���M�Pz}��,�(�ŀ
�H�!�Ă)�����-v��F`M�z�!�Z7 m䐘(����Qcn��!���T�!�Ģ�u׎��♃}�!��#`g�$Hw�Ås�
���!O�!��#9�xd2s�#�<J7�A:
�!��H� ۚ=�U�'�nl�sBǦK�!�$b��<��E �s�:�˵�_�;y!���4�D�J� �+
z�)�[ !�d�w�P� +�71��1���[��!�DOn�d�G�	*�Z�z�)��%�!��μ6�Tq���ȕ�X�)�N�!�Ҵp�$]ԋ�*�4ݳd���!�dۑ.G��A��23����Cɑ�`�!�� �6J�r��L3o�F���&*�!�$I)Y��ɱ�O]%���x�O	+{�!�ߖ#���s#�7�����̝<)!��^���9u�#�6-����(!�DM!v&j���ט��8�!�>!�$��5�^(;C�Ԛ
�T�c�l	�,!�dǊw�JH�IX(b����JJc!��ӬEh����N�wt�a��O�a^!��>�����Dq��2˖2jU!��6i*Ȉ���5>OLD�"��tF!�,n2�8j�ɲ;N��vH��2�!�-d���3i�7a��q����L�!�d�#6�TT[G"ԛ{���f'�<V�!�$ȸ)&�spO��1v�!ug�>�!�$ʣ)�����i
0
�D�C��	B�!�� ]�SFG�H��i��i�2�Z|��"O�p�� 3v�!_�r�U"O�a`gƃ,z�����2#��B"O"��1*���9�ud���Q��"OD{�`V�Z°�J4�ŧ4��Q�"OT6/�(lX@aIq�K�U1(]��"O�9�,�,'%�
x<D��"O^hsv��w���q�Z	_e&=�"O�����/-Lv%�1j/W��R�"On��wƋ�H��̓�qAB)�"Ov��� ��R���Z��Z�4,4Y"O$�`vhU�w��8���n�~���"O<dJwm3p���s�Ƨ'��v"Od+�d@�d�210�9g��@"OfB�H55��(����.B��;!"O�e�a5Gr �a��M����"O>$jA�� ��� �.v��"O�p�C�T���!��!Ǟ?
`�"�"ORt�&I�C�z@Q4��=
� q4"OZ��bh\�F�4۲M����A�<��j�	������P�����w�<�##��U $�1'�O�v��h�<� �־�h�Z����[:Ras&Bg�<YP�֋\��Y!l�%S�L;D{�<9��:9z��	 d�#YM!P�P@�<�s��zEb!��*�7m�0A��ʛ|�<�!莒e�ּ�ek4i�$	�O�o�<���
$g���Ǆ��@����j�<�DG�:��9�oR#���p��m�<'P�x*@�1���(W��p'Mg�<qDJS 2�L����6���$`JK�<���A66?��T�?>����K�<�Bj�!R���pB��h�c��A�<1�NH�:� "%��*i�m�WO�D�<)2�94XEcS�� J4��p��C�<y�B�!r���铫��#��J5AC�<)P�E)R�%S�3� �BR�y�<�p�	�ad��q!�ҏo�l���-�M�<�ToA+�F�A��_�Pt���ƪ�A�<y��
u+~���W�9��rWJ�}�<���10Y��B�L[�����|�<)D�M%��UZv �YUxܩ�O�w�<� $��Q������h�JM gA^�<1�J�'�����Ѽ�vP#���R�<Y6+��t���)A(H�,�M�<��Ă����vƂX�j�:���I�<A����i
��I��\&Zc�%[�"E�<I3G��Sw�L*��"a�j)BFLA�<�dS;F�R�$�
�j�"0�d�<iG�Z�9��L8�CH<68r]�D\J�<���
���h��-���C�<QƃA�n8
��AJe�KS#�C�<Y�/��I�ԃ0#��g�P��Z�<i6�$�t���Dl4�bs S�<���8w !� ��C6b��&PN�<Q@f�+H�|��%<|���&�L�<9�hԽwCH5(�O4��	�TI�<�M`;�p��ɛd�$!	0� B�<	G+����᪅`#� 0�F�<�b��WW�5"���L�`�
Wv�<q�n�E���V$��]<'S�4[�'�n���@
�1:X`��΃�J�d��'��+�M�#i6�P٠��z��\)	�'��Y	`D��8~1���\"#nD���� 9ѱ#��Y�t��t/ޞZ&
�3"O�@�vCH�(�1�p��3v8�"O� k�����F��ԛj�A�"O�@k����g.z���L�c���Rd"O(h
���p<�� �3k��@��"OD}��#M7���u߬X	����"OP�
Ь�����4GɆ)��� PE"D��*��6Z�hA��mA��xw�?D���5�*W�HmReHH��cС<D�����Nެ�p�ř�0�~���9D��B��w&
|�TH�U�naA֭<D��s����SYJ1�蝙iK�H�B�8D�@%�	��4���Y=ph;�#6D�P����-�����L,QBm6D��	T�Y#z���4F�2wz���2D��Adϗg�Y(�Wg�x�3�1D���M��i�C���18dj4D��S�Ll�8F����eqwh?D���!N��:��U�uA��uo��K�M D�؉���K�F}z��y`��X�!���jC`�W�Xj����D��!��G�
8nAb��,���k�;)<!�Ē�r�4�#��Y�Xs�	C�55!�P�Z�Dt��� #X����I��K�!�$+d�YR��v�S��V�M�!�D�J��,9�M�	l��XK���c�!�ĉ�i2���GF�����$81|!�
) YL�1��R]3�#\�~�!�D�-A�r �#��Da���,�!�d¸S/JG%_�;0< ��\1A!�7�B���L�.E�|1�e� D!�dL=q�t����E;m�Z�Y񪊄D�!�d	�s�l�;�G�nЖ�*���!��S+�^��6`U�g�q�I^�i�!��	C6݃��5 N.eB�'_��!��e�-a����GA�񹆍]-Zk!򄜜1c�s�`��p;�� @M�0vR!�|k��br�$AB���D�!��B鶙Z!/�990�yi@�ھo�!򤎰��Q#�X�F;�\���S�8!�䃍&���bْF-�a3Qj��O�!�DPO}���V�Қ1D��)[{�!�dהy���гt.@u�jM�$�!�UI�"����>x��I���N4!�d1X��(�㘀8h�����":�!��ϚY����p"�*Z��l
��B�-?!�D�mM<�ڕ	�uO�\�M��5%!�d�(g�d�TlS	P@,,�W�Pa!�	kvdĈ���5-��Ʌ�<!�D�%(m�0z���\oX��Un�P�!��љiҸ%P�J1[`�d�6�u�!� qz��` ��Lz���eJ��!���p.�\�s$Ǎ'6<�{%l�!�}�B�,�)b�8�ɷ7E!�D@����� \+B'.��ˈM.!�dܮY��'HE�<t����Y!�D��*�ꐈ*ɠ�M/	!�DE6�$M@s*[�)`T�F�WeT!��nي�xM" x�!��`كv@!�D�!+����W5h���%Q1T!�D��$���E%�X���8#�B�%>�~d�7GT���hpP/�"�xB�	,�H9X���)˂ ⓪�pB�	4[�`m�5\�t���D�?<�XB�)� &5z��:����+�#p�Hx2"O����T�:�R�P�ٱ'�2L��"O6=�3�8l
HjW�W�X�Vp %"OJ�2�#H�M����Wh'C�>X�"O�pq%=�p*��-'kL"�"O��q��8$����3xU��Ц"O0\���N�~��U�K�I<,`z"O�ՠnu�����l�gY�U�"OZ�)�{!�cf((PT���"O���,��H��i�Z0���u"O�xP�gݤG���V`�;/s��e"O���3K��+qD�[uo.8@���"O"�r�j�-F��u��n�!+��z�"O2z�KA2_u�t��畁g���"Ol�`���HVFH�	O1���y�"O�����'��hsϏ�bza�"O�%��N�v_@8���=�N���"O̥�*�
Of����C�n�
��e"O��3�ү'������J�6+�"O�m�ģ�pk`����[�8���(�"O���3́*9�"vg�`��0�"O��0s�(i���eS�t��Y "O��5GR��l��N�r> X1�"O8�HT_#��	9�CK u�.p�"O���81�z�:�̈$�RU�"O�=�V���G��@Qa�;.F��"O��@4剹9iC�� NAxt"O���aN"?��g�2v�JY��"O����BN-*�L�5��PC"O��X�g�^p�pѤ�5c<ɻ�"O���T��/��)�� J��i��"OX0�*ܣ_�|�0�n��8.ةy`"O��C��g��� �H
1eȐh�"O
-��C+p�tL��g�n<q)a"O��[�O�wcl��p��o�0�$"OX�%k��FV2��3W�Fq�c"O.�j��C*l%Ф񤊊�La�"O|l���ҷhg��*0i��6Dp"OF@�g��_�}Re�CC�<��"O�YjCD4U\j�S��5p��tc�"O��h["5h8��U)�TS�2O��$�"��bش���+�p4�f�(JgR��[�b�����1=0�w�XF��UU��1;�p�Q ��(p�-�Ͽ��(�He�:W��.�ޥ��_Z}�Ę!Gq8m���{��@��:y�U�D����'T��	�)�}r�����J�L�'n����C��v��T�OS���0�R��AHz6J�hŵv�0��F{�OmZ�	*:���g �{�,a��RP�>��i�L6��O(m�k���X��{�؊Ka��y5i��) �$�<���E�:�V�I3�j�ےo�*N�(�����r"���0*K �fx��iw��ht�?i�S�z}�hj�f�<�
��o��8�Ɖ�9v\�1�CO�E����(]����w�67V'>u����0��l��3�)Ҷ ��'/?a�V	�օ�<	�����P%�����?����MCP����aS��D�|���e�A��-�O��"D/l��r22��8j��Ot�l%�M;N>q���,O��DV0C��FJкm삜'��@iX%oZtx� �	�s�:U΃(ch$�saP#,u�8��+�4��#� J�ԍ�Q��ׂ��'ʓ)�PB�&�*t�ȍ��΂7G Հm]+LLB�rҢO���JGG\�eKY?!�#<��#Ԧ!��l�.�J$�rBH�l2Tś��<�D�O(�$:��>�YWM�!(�\�sq K�57�l� �>�E�)��wZ��g���R��CH�u{�'
:6M�䦽�'�kC�b�\�d�>Ir�B�PP8a�v'�0k"d��`f�'b��j5x-��	�k�ԑ ��N�LJ@�+��e#��?�p�;��ũ��N�'�4 �)ߥ:�
M8��R�[���猃�|���b��b*�](��5��<P���O�� ��'TV6��d��N*QPBG�����k��Rs,�����d�?E�$#4rҕn��0c�Y�O�912B��d��:�F�=R(U�h��diR��F-M4��I��M��'=[���'��I�?��D}
� ���ゝ���0����~�Bę��ܟ��
8�h�$*iCj|���
1����SI$�]]��c o|
u;.E�%D>�Q�B0z�JV(`N(�P��<,��G�$�\�&>I�4E��B5�a�A�3,���c�>�A���4�&�O���*=A@HE�@$�L��î7qs��>Y���'��O8El\�ʾU��?�0����?�M;#�iR�'=�.H$���L_2A���ȀS=����}y2��>^�6� �冹�#�7
�I���ј~�H��h����;j��Db�4��4�O��ߐ��D�DBHÑ�{��A#FKʭ-��<qCf�E�]�Ď�3[���������$\�����O���"���2�`��=dQ�&kڸb�D�m��0�g@ş�W��,O �c�lM('"9[��d��f�3�,(�W�O�����;�n�	�Cah0�e��\����U[ش��1AȪ�'�������r��Y��T�l30X�eH<q���   ��     �  &  �  h+  �5  j@  �J  �S  N]  �h  qo  �u  o|  ��  ��  <�  ��  ě  �  O�  ��  ٴ  �  ]�  ��  ��  <�  ��  �  �  ��  2�  � � � �$ �* 1 85  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����'�#=E�tF�@0ڳ�ޭ\��kD��yrMQ{�<�q����5�����?��O�U�O�g̓*u`���k�heSc�~���IG?Q�K�H+2T��N�|g@(�c�G�<&�?8�@A�3��w_A h_}�<��eu�t����Vゐ��a�<�� P�VV��k��R�&��up��u�'�S��Xe�!�uo��#�'Ʌ�v���A�.Y�vKD�kT~�s`���<i	�@���$�ǟe���;���JE����;@��fD8d�QK$߃i� ���J
�ybR�wـ�SvO!��Bb��y�j��r������(��ڊ�y�Ã�0y�@�K� ꨐ��@[:�~"�d�M>��Th�>@�|�1���!j@�# %D�\1BE۰!z�����.J�>�z�"��p<	�EߦJ��(��@�\�TaH���~(<ɥ/�Y˲���į'�~�����`��B��.PT1�eȽV�N�t
ŽlB�	�I��ɀNOP�T�P�d�hB��&��䃣�F�oT�j,�	��7�S�? `��e��')�Ģa��%@�"O`1�P����G�6�I��"O�Y�
�L�p�J����rIñ�'��ɲ'&<�7�_�@��x[Eoc��B�	�c��E���=ںpt�J6X�B�ɿL�"��Nj
���T��;��C�	�(i�r���fCؽG
�lM��Oܣ=�'A���-i�.!��
%��
�M��UbC�	'FM`�# �G�5`��	r	�Z����'�1O8�?�ӫ�#/ �Q'��/"};�{�<!��F�1�r�ʰ&�/+d������D{���i��+d��o���U�<q�xyk�'S�X���	
sN��j��p*�}[�O���D4s��Xð*��8ع�M�����HO�O��$O6��ȦhD$�$�8�%e�!��R�WĄQ�u"L�"��h��ئ3�!�$�2���eF�X�beH���'s�!�� �WB�K�Na�"�I��`_+8D��#�ˁ&~F��� 	�+$jP���#ꓣȟr�C%Ťԅ�pI�>%��@��vx���Ԥ��9�}�ˬepԛV�*�dd�l�>�O���U;v����h�) ��%A�@��*ZdcWOZmIrk�1��}2 .��#�B��r���I��|y�
��4�|�	��� .�ll�";$�<�T��'?�5��ƨQ�x����Ֆ�M�	�'�5��h�@��5(��4+FH	
�'j\}*���U��@�� �' �1��!,O$qɧ� y�(��Q�V�U:���"O�d0 ��`�`���#C�q(t�ò"O�MJ��̂k�y���uh��߰<1 K��4޾ �l؝w�F���Cx������䙶��:S���.c�!�c$R+��h��'zP��Ì�#�+�UۈdhP�Eo�<�fh^@:vj%�֍C>Apw�E�<Y�@�}���bF�*� � nCY�<�!�Ŋ�fya�EW�N& Aзo�{�<����lP�V���� e@@�<Y����[��M�T�G?6�-�b�D�R�C��`�9��V�8\3�	D�-��C�	 G�8i2w��#eJ��HXC�I�'ţ���,G� !1��l�dC�	�A��}��JZeD̘:�aX�tHC䉑^��صE %S��94���JNC�"6�-����!q���2F��09��C䉺nG���V�Þ%�Td�&��C�ɉw�ƹ٢��
\�0) ��9C�I����v,Z�u_�1"�Z�h�C����h��a&y}6�	9e�h)��.D�0��9;|��C�ױND����2D����g�.y��Ñ�SG�|�WN5D���J�6@C��1𡐔A�: {��-D�J׎�B�,ek# qо 3�m*D�DJsᎪ@`�s��Vݎ�ZT�3D�HsM�'l��!�kw�|�4�%�OX��3h&�Sk	��&:��W�A�B�."�Ԉ9��\W$�<�iX�tw����Kq�'�����[��f5�ChV��nL*cO�	1���K�m[��'�Ȁ'"O�}qt�X	@�2�*pe�<&�t w"Oŉ���%z<�:�ƈi`������T���>�Ƭ�Dg[!�5�Q���K��ن�ǖP��)�8�	�#�;n{Hd�ȓ��AB͞:LW,��')��Q\8t�ȓ�칈ݤl�(H!Aj�?�t����)$�� d	��ӫ6�´Bg�ڦ@���'�'�O�ܹ%��<de�iRD�[�x�~���"OPt�1	$���2�&����C"O�	Rc�C�!Ñ(H�@��aP"O8A+�*��� "�C�n�b"O���!_�S���C�_ �A��"Oœg�tf�i��	-0���xB"OHp���ϪU;@�� N�k�81�"Oޤc���]�$Ԑ#"Xk��1�"OH�ç�U�լQ��u�pT�R"O�q�CL������	3��S"OX�h �2d��s�ݭ#��ɔ"O`�;�%��T)X%��0�h��V"Ot �o��DXHC���%�p"O�@2 �|s� p��s�, ���a�&�=�O0�X�������#�4m	��'ҡ"�77�lhC���\���'#�'a�S�O��p��퍿\ɲ	q@+���'Op�B'��1t�HpW*���		�d#�S��?!����(y�C��{�`@��^����'�D� #a�����V��B�'3�Ab�K-�t�y��B�PD� ���k��r�ɒYJ��i$��2	�C�I��ڴ�$G=�ȡ��=7�D#<����?EQ�R�1��R�gH V�fU�#e0D��ɴ�@�ؒRTiH�8�ZEr&�;D����ڟ)���G�ɓ<�R�bP�9D��Z�!B6Z��굉�8s�4ɂ1�#D�XbB�Z��ۃC
Zf��Hg�"D�h��n� 8X��AW@�����e D��ciO!	�Q�v��:EX���`,D�P��f��萙���,���/D��������z�G=�Z�F/D��X�ݦ{ ����㞱|	|}��3D��a��V1i^�M��%t"�a@�.D�`��V$,\ƽ ���Jy�j��8D�D�`�((e��#�ǌ,t��@��f1D�����%bY¼5H�ܨ�7�0D�<���@�S�S�,ʕRȼ� !D���Q	~/�yWI0��,(q#$D�pAC��9ن�!$ ��+�$=D� ��"@�cD9ӱ��!`���0D��B���>Cf��d�D��@PJi*D����;3d��QBj��;��!Å�:D��)���;������_���n-D������	m�(�0Ѝյd�М%�)D��Qv�*e���'�R�:*�:U�+D��I7$5CG�1�'��n
�xd'D�И�ª@f�E��B	�U��� �9D��
�IR'~'T��cΈ
M:�m*��5D�|�`�-(�N���G�]��1��,?D�ȉЅD�W�Y !�D7=q�Q���/D���Օ1@�IK��\(I[�ur� :D�HAu\ܠ�V/٨g\���/3D�`K���9>|��Ц�:?v���2D�\� W����bU�;sB��B0D�t �DO}�ə����X�>�+Ʃ"D�<I��^��̙�#JqhL(&�#D���kM9�:8��2o1r��o"D�ฦ�خ]�V���Q2������,D�@��IuEp��o��F�V��,5D�4 ����i)t��"ޣ" 3�3D���Y�mdh���\ n�[�b5D�찧�eg��9�[�2��D��>D�� �0�CD�E6�4�`M�8( �܀�"O|dB)� O8�J�
��Bܢ�"O�)���@. �"���S�B_����"O��aM�L� H �8�5a�"O2ܲgd�X�("�Ά	g��g�'Lb�'��'�b�';�'"r�'l�	�KN�n����ь܂a�&h
��'���'���'���'�B�'���'�*��s�Ƞ-?���ʅc�����'U��'���'&b�'m��'�r�'Ny�e@�)�ȓ���<k%�F#�?����?���?!��?����?Y���?�X\�C!%Z�dR!+���B.������	�����ٟx�I���	ӟ,�	1r�"�e*��z:�y��ra�	���ן��ן4��ʟH���H��~�~��A���`0�pY�,����	��L��͟0��ݟD�	���������6c�,m�K�*h!��`�ɀ�7�� �	�����˟�����	�	��� �Tj`��=�̵P��ב<�|L��ڟ������	ş����l�Iӟd�	%*`P�&ڀd�A�P�������x��T�	���Iş��֟��I zt�s	�+cY��;�j܇�����؟L�	�h�	ɟ��	��Iş��	F
Y���L�J����g��~��I���ݟ(�I�0��Ο��I������¦^�&���Ag@�*hq ��Ɍ矈�	D�Iߟd����,�I��M����?Q �����HA�
!�� ��`� (Oj���<�|�'MP6M�*a��J���b�^��G�B"10���d��̋ش�����':T7�G0t�̰�F�� rn>t(�G�v:�o�ܟ���b�`�IvuvYZ��B������IBĉ*M �%��m�FX�<����=��j ��K�/�B1���(�����E�Φ�)� 0��~�'E��w���'���T���W¤h%�qӄn��<a�O1������<��_;_���@Bн'����<��e\2.=J����hO�	�O\)xOݔ
ݪ��6hI4"��x��>O����Qj�V��Ø'k�ᑃi�	J.HPӣN2y*T
���HI}�Ew�ܕl�<9�OnL�K��.�<��T��Ny�������C�"[�d��>�'nO����'�?����-|tCnN����`��Z���D�<i�S��y��\ Re:�X���`%@�惦�yd�~4㓟P�޴�������T)X�Ê�;f��*��ymu��]m�˟�8s��w�	�YO�`�ܑ�:�i��@T�"hp�V�G��!�\��My�OJ"�'t2�'1�b�M��Y���R6=_~����L�; ��4�M�����<��?�L~�Ql!;Ҥ��=Z%�E�Ժa��U�V�,�ش}(�M?�4�$�i�PR�I�-kX]���K�S��`)b�#Ex�*��<��R:E��x�������X�e�a���5&�F,���~����O��$�O��4�P˓�&��y"F�$�lI����Hz�L� �S��y��pӪ���Ot\m���M���i�d��&I�P��4LU� ���d�\"S��I��D�R�J4p�yqA�[y"�O���ӺA��9R�o�G8F�� !I�y��'���'S��'����Z�5��X����}��D�ƠH�����@�4:�(�'�P7m�O�ʓ�"�� �(e>홄�>8���a��x2�n�0Lo��?ͳ�Hly�'��MH�Vx�@�r��!�*0����3$u�l���(.��'w��⟠���p�IJt�8��(�a���hs�x[�R� � �'s�7M�hb��i�O����<���/Qʹ����@���I� b)���O�Y����4]��F, �4���)ߣM�x�iA��k����捙 j�=ZB+�
h��!��>Y�O��{�G��[�2=������ٻg�I>U;��bG�[�^�����>]H@��D2$�Y���'�V�H�P�è��Ɓ؍!�,A����;A��6�[g<����EX�:�	�Â� 'T
�l�E���$���'�a�3�P����ԫ�B^0��B���e�3i�q�2!�����hp]v)ҸQ�JY T���-�-��A�:�J]��/�V�Й{�iӅ��S�(��|��-�V�Ӥ�ƹ��G� J�@��С0��p$��a�A���U�<O����O��d�<��?��$�+tV��Ҩ_.kSB4���	G��m�J>����?�����d4+�hnz���5�C&P�@��*U�r��:�o�>���?O>�,O1�_� @`��
ݨ���StFh�I�>����?������X�ν$>Uh��W1�,UB�A��tEy�,���M#���?�*O����O���S��ҩPƈ�� j�|��	g�f�'�R]��pAU���'�?)����8XPt@F$2�1l�ئ5�'3���EIf�O��ܴ�Bh� ��1��@=E�0�ohy��C��7��~�4�'����>?F��@ź��ږ2s�i+1�O����I�p���uyʟ���x�LɸӖ�-;���;�M�S�I�<ٛ��'���'G�I;�4��p�H_(EPx2��Ǖx����͓��	���&?1/O���O��s�\P��c��t0JӖh�̦��	����IU\M�I<�'�?���p�lē�DK�*I<0��	9H�Z���R�P�I̟([�K-��ޟ�����LxR �?9V�Y\7Q�B ��B��M���$"δ��x�O	b�|��O�T@��:�E�E= !�V(�n� ��<���?)����UR�*�k�t�fM3�"\�WW=��%�o}�[����Py��'���'[�� �)Ff̴EN� l�<%������<����?���?�����ċ}�<�ϧ �n䊐�џ>Έ��S)Qx8�o�Oyb�'��ϟ<������wHj�֘+�θ��үmc1wQ66E�7m�OڽB��O^���<��X�E��ӟ�:3cNS�-��Jz�L�����M���D�O��$�O U��4O����O��s�+-�ܹ�`AǻD�p�E�V�xF^��Ov�I��,	�P?��IΟ��S>��](��Z�R(J!b��F�8�4�O��$�O��D����by�ܟ��:�ԘP�l�a����Y_`(��i��I7�u�ڴ�?q��?���r_�i�Q0�/
0X�����Xk�cD�z���$�O��<O�O<�>����L���w����r`�#mӘ�hE�
֦��I����	�?�ڪO�˓,���Id�T-K#��N�>�,A�2�i�N���'��W�(�"�I�h��$�/B�|y��F81 l��i���'�bEX!Kɘ�����O��I�0Q��eA��yR�A�Ke�7�O�z�:��S���'�r�'0Ys��C"4p�:��
2�L�3Ev�z�H�j�Y�'[�IȟD�'ZZc��02A�.5��1顬G,L��OJT*g;O����O8�d�O8��<�1/����"�KT+[�6�i�X�7{����]���'B^���	�<�	�C�<�S�$I.,a��aӁ@h��")j�Ė'��\jA�'�[��[&���d�7g+���a��F&�⦬٧�M�.Oz�$�<����?���y��ϓiΪUˀǅ=[)F�8��Hl\U�`�i��'O�'�*m�|�k�� �D�����KU�e�d�0�r	q�fc�L�$�<A��?9��w����?A�l��	�
s��#���*��G�D/�?����d�/P���%>����?�hsa�2I-xh�4�k\��	�=��'�'�Ջ�'��'z�i��]i �Xd�ם}����'��x؛�[�lz��_��Mk�]?!���?�O��)��9t�ix"(�fv��Büi$��'ʠ�q��'n��z�O�H�[F���6x�0ᒮ��8}�!޴k����it��'w2�O��O��D޲U�0���O=�ԥ�P��M��nڊy����?E�4�'�z`L&T��0�V�'	>���g���OR��	��$���	˟X��~z��Jr����4l2-��n`�	�%�	�M|B���?Y�A$��0䛷3����F�
�7� �3�i2B�~ �O0�D�O`�Ok���{�Rq��=?_��+��r��	"h6���yy"�'�"�'���4s/�"��v4�Y�"���e�-9�J��ē�?Q����?Y��2 ڈ�Vlq��`1��"�(�q�iR�<1/O��D�O6��<�.3��	�JT)L�=�z��V�����(����,�	(~Jq��V��\��M+�P|�w�Q_
E�'jB�'�BX�`S2m0�ħ0��(��������I�4s)���w�s����=���O��dB�FV�%}�^+|�ma�"�+OD��O��M��?�+Ot��֯�~�ȟ��S/|;B
�Oi��pZ��@�_1p1�6�x��'�&ϟ�2�|��ع���NOr1����0���A�i6�I��ℛٴ4�����S���SJ�@��v������!@�)1�V�'���0_>B�|��t	�v,�֏�;_o��@߷�Ms ��Oޛ��'{��'��d�;���Ov���m"H��[���6N�Τ��ɦI���x�|'�h�����r�y� A-x5p%cU'�j܊��i.�'���,]��c�t�	~?�"�hچ5�WořuX"��o�ߦ�%�� W�0��'�?q��?�CF��8tus��V[]F�Y�ѱ\a�&�',����+��O���+���p������gш>���уJ�T}2��9��'���'�2]�ع�5��%� Ŷ>�8��*0z"��I<���?�I>����?y�����]IP�\"%N����@^|t2���D�0>�HQ'g� {\�W�8 )�Y+b��ze�i!������}@�B�M�X붊Ɏ-YА�3�S|�!��	m���y왔=��}���	�-��n�rL�i����,X�5��1�˿!۬\0��+Һ1�1
��k��%�HO.3u�b,&����_7O�,T�@��j�Ӳ��W�(�R$M@0���V��� @"I�MzDA3qLLe*�Yb7��>��:d�1Ӝ�1Bƕ�NA,D	c�@6��z�*A�SD��:V��O �Se��`�o�8	+�� �O����|�0�`�6�����e�0��邢>E�'m[�M"�C�.i04������|��O�ԃ��֌W�y0�K�,}�(B&��?@�|够�U��KC)d�,tx��:]�P�>��
���s�O�b��g�xD���^���``Jݾ�yb���X��e�b���L?T9g*C��0<A�I�pR"�X��E�)�	�T`�M����?��;6�ȕEE��?!���?1�Ӽ#"aZ�M�<4���\�	�4�с�2AN!���C�S�!+�n�t*��Ĩ�
-ƹϓ_�x�	wFM-"M�ҁ�~G�����CG
L#�cS0�8M��Sܧ��`:B�{�xЀ$�l�2QJ�! 6*<u������)8e�)�3���3� 5B���]�\��@��;`d!�;>�@]3�¥�꘢�dW�X���O֡Ez�Ot�'�R��cK�_���������1{=�0���O��D�O����Һ���?��O�2%)����&c�DAF.�77�\�'�l�Q@N�V�������E���`%�G�'2����	�\���-��L�a�{�r)k�č�xwt�z�)G�/V���T�/  �<1 � ��8PJ��k��P:0�ݷ6H.ͳ���O���*���'���i�b��ę�`��$:baJ�'n�)���� x����vN:�j�y&oӞ�Į<���ˉ;x��ӟ��&��Iv()R,��T����ǟ<��5J��i�Iܟ�ͧ`���g��g�a�!���]�ԍBd��m#�В)�n`��w(4O��F�(}t��,һj�¡�d�z̠�\-h�qk�j_��p<�fl������Ny�cR�L��|Ҷ�M�*� 4��<F�1O ��'<O�|�5K��M�zy"0��xzYj�O�lZ3Vۨ�B�
���`��⋦hu��	{yҦ3?��7��O����|2Qꅝ�?I�H�	2 ��DjP�$��[B����?!��A��%hѮ���J8Un�	5g�8�����R*�hs�G�w�>�S0�?�^�`ǒ>AU��(5��,LZ�~Y1�_EdD��6jDFEt+HeX�d�<=����D��9}r2��)�9o�j�QTc��H�+�t	!�J0Jt���hģa:F��$� OaxR�"ғjY	5���1��@c���jjuB��i���'Ar둫G�<@���'��'��wh�����O-+$	{p`_ˢ�*���i��yҏь"��+��~tD���bֲ��'�>�Z
�pd�qcLI�,$T����'�HT�|�l�'�?�}&���'��!�� �Wʍ�VB|��6`>D���R	@(YXj1a�M˂x��->?�5�)§}���(���� �����5L��XK���V+�H0��?����?���Z���Od��*hn��	R�"y�{w��zh��B4넁�`ي���wg�u����5sҦ��s�	��L�X����d���B@dN>f�A��ϖ��
��	�4dBp2Ս^�<��� ��		 ��-9#�߈R��@�Ceײl�,Y{���O����ɪ �Hm@�j�2�|��*������d(�dL)b(�$�J�q.����΅>r1Ohmm]�	�R�L���4�?q���$J�ǒ;H��HR!0E�h�a���?���
�?����#� j<�8c�L�r�hH�?E��\�\�6W�qX'c(mrԘ�M�-j�]Fyb	ܾW4�Y&Ě4^H�t���4��`�A�M�^�(0$�ҫK�5I�í/tEy2����?��x­��t ��M���R�BU'�$�y2GS>=�B��ϣc����'����O��=�'Fe��iV�w_�9�%�Y/$K���?��'_�x���t�$�$�O��'S�J����1G8HVe[$���bĭa	^�J���?q%ܱZ,�f�+�M3�F,rT�SV��l��Ө2�*�H!KQ�C�HE!�lW4v(�'�^!�A�3Q̼�!P�;H��+�.�2dBq˅	L�f�N�7b�~=�Ui� �\E2!����	��S�'X�& ���d�b|���ǹ+���ȓ*��4h$��d��͹ŏ�-a�r���4��4Ezr䘲'�T��1E�>Cbvi���uQ�7��O����Oe��l�,HKL�$�O�d�O�NY�IB��h4ۂo]�$F�=Q�H��e�B�q�i�L�wo4|
�j9�S�w��sV<O����A=�썹���7Om�b��Q5,ƨ�P���JЋ��w�q�0��� �y�.ũv��8 '�1TH⠨̓\�P�OZX�������	,���\.Y�4�6�Â_
e���p�����91�tɡ�a�\"�Γ�?�T�i>U%��zb�';8�`�Rd��W�@�C6�
��R� �N������@�	��u'�'�b<���*�k�`�$8�E�Q���6G�	[�TD{�C
a��1�Q5U� ��m���(ODk4C>Il�<�q�@H����a9���6 �+<V�P0��.F�$huE�%�(O�H�K�<A>���'�
��\���ȑP�B�3�O@����#�It ��@��s�'o�'0�P��H(���7Hھg�8Q��y§e��OеCtL˦�IƟ�����G|.���LɦG��������L�	+��\�IʟLϧf���1�M�t� !���G�Nu�m�#�m�84��tЀz��X)^`홵O.�x�:����1TJ��X�9�a"�}����CC��i)�`0G�7H��G/�ZV��M>�g/�� �	Ly�E�-�f1y�%��a6D-p��E��y��'QB��S�Tzj5���A\ 0�ꉁ8S#<��4��YmZ�l���BBů4dpԁ�:y����`y".�}�6M�O �Ĳ|�`D��?Yd��1�Z�k�%&gL� O��?���@��������	.J&)�G�S|���E=}k�O񟦁���@v�έC�J ~ON�#V�>a��՟��O>�2�WB��uY0�Յ|U2��E��p�<�r扭�����L'PD	 c�l�Pc��$O4o; ��T&��U��#`dH�^��@o�4�Iޟ$���_�R�~(�����I��]�Q2�yᡮK�HGXx85�	�z�q�<�Bbx�ihV!s�$U��xf�t#f6�ɭ���$�V�BX{gB�|nl�� U= �$�p�Ԡ�Oq�ɧ� ,Р��w�`0B4N�A�^ �p"O@|�@jޥ���P���6dr��Ӟ�����ᓩE%L�P/�VXD!2�# V��U-��:��5��ߟ8�	ܟ�	XwFB�'��)��[ �6�V�%r�26�ہ�I@�$̀o��p���+s�r��I�t? �����Ȁn���R�AƃR�4ݚ��%�Vib@�*"Q����ޭy�(�a��6��S��$�0ԾQ�^x�BƢ����H1�^���,�O��i�c��(	ry7/A�7-a�'�'n��"P�ҥh�&��sH�y�ƥ�y��sӮ�O��Ч�u�Iӟ<���{�^�3�'Z/拉�S$�� �	9'����؟��'X҆���]�	�i D��kV�lq�v�0r>��T�g|X���#իR�.���t�\�j���[�vXpJ��*� ���'�fQ���2�'�<��g �+c�M�7ʒ6[T�Ȃ�'��R�hQ,v˖�+��ҧK�(� �'`7-�VI@�㙇y�@�2�%C	LrP�O��e�ɦ���柴�O���3�'J9k��!��!�k%6NPP"��'�R�� ���c�	-e��*�H���*	(�L�>O�S�36D,�5�8Q�4mƔ9Hb��Oʱy�"Ђ9\D��@%����#!�ɟ��q�ߣp�p�X'ߤ0�x����>��N��@�K>�J�K�S�QrFW�U��uc�G�Z�<��k
*%��P�ʿ`.@����hO�v�'��=�iH�X�2 �v�F�D�y��M~�&���O��DA�&��DF�O����O4�4�nH�MOR�Q��Dwt(���B ;���fߨ(��xC�Gňp�lb>�2���G��$�s�\�K�+�'^���prƐ2!���9n٦W�d��Vϗ'd)���O����'!,���f�w�P(C���
4��m���2�D�4���L>q6�� �Dp1�@B�����g�<�� 
d���20GيF���d�R�<q��|����c�I5=��HEl�a7����a�J�����&n����	� �	Ƛ@]w1��'`���A�1y�CR�1�E����B�f �pJd͢b�i��L��;�t���&:� �B� Z(�C�
9�zU1Wg��[ Y�AD9g�4�c-َG�����,-h&��Җ�:2T
���8RRJɊ���r�(�d�e؟șb*R�
W\��T瓉Rj4P�2�=�O@�O�E��F�0Z����/
�I���D�Ц5&�������M;��?�%"���1Q�'P�Y����,A4�?��;�����?!�O�F���`l��Jݴx֎�XP�ɦpŊu�7����:�(K=d3T�����(O�u�w��-,�V�[��$d~�pb�M�Ub��	ǯF�<ݼM��O�Mݘ*V� C����0+7�$C�2i7�d^.PҘ�H��Q<]��mC3k�,�!�D�8h��3�c��|�,��沎�D&��|*��i�VE:�F˞o����N�[;~P�s�|B�J�f.|6��O����|:�ę�?�W	��y�ج��NP�S�F]����?��s���&�٭
�-�$Ώ�a�<|9DX?	�O�~l
�L�4�♻��x�FyO��J���FѲ���za0���AXg�GQ&(iu�/�� �"R9L_اO$9��'���O�V<�b�|� ���˔@�! �"O  �
�&/B�Q��O�|����'��#=����F9�P⤐$!.��0@M�p��v�'i2�'��;��L��'"b��yw���V���E"^
jP���H61O����'m��!G|��� H�.��{R�Y��<qR�LGv9�1*�Q��!R��W�'���S�g�ɷn�&���B�n
���h�(��C��0\��$���о",#���vH�����"|��ە5��Pk��P@ͳ!�
�G�T0$���?Y���?��4��O��`>�*��@�&T̩Rd��p�Lt�
_�J�(�i��X>3�i	g����'L 2Q�i�]�	�Y��H�����������P]�W�@Tz�6N-�ـ�Q>�Q�H���A Ѹ"㗴z���:`"@�I>�ėM؟� � �5 ��N`.�=)��$�O��O��� ��1[$�H�H�@���p��ަ�'�\�
���M����?�'�	fX�����,c8�6��=�?���o��j��?��O!�(Z��5_��ݴk >��B��Ob��!,J:R�eB!���vb���wۀ�(O>��a*ʧ`���"J�f$D��썸S�ݱC��	s�P�"�,J�ƞ�D%yT+-�$���-�$�hFݩDB�T}VU���ްC�!�䝲<x����D�Te�) ¨����E{�Oj6��9nЃt��W\݁��C<k���O"Mk/��e�I˟��O�0��'M����Bն.��X;�&RT>�qY�'I¬�)�5@ćU�T@x����Y,�6�2��c?��-h��D%W=HjȀ�Qn��r*��'�44XT%Ж&��,�c�*�t�֯�G0U�O�L���,�6�1���/t ��N�<j4�O*�D�O���;�ӌ5��S�� Ѭ��?�b�<�	zx�� �y�a�
��P�0�HU����h<��|B�鉐%�i�p��wH�8#"�L����4�?���?ir-	8vc�����?q���?���C �i�b,�'	��)�"�=mDD\35�?����&Ɔ9��S�"G.ØOni�E���<	c�/Jo8��<�|i����3��p���(��Ɛ�lڱ	��d(�-<���l&bD{Ԉ�/4�b��a�v�jtkq�|r���?�}&� �C��82Ҳh��c��)�c�9D�p��Z�v�<���ru,�\0�������4���O���dE(��"bR�2\�� q/�2�E���O�$�O��DFٺ���?��O�0B� ��
�@�G*ݎ6��(!�R8\c��sm��M��ß����LA��(O�ZŘH��$�0M���2t�"��:R�a����ܒ�+����2S�X�r��d�#�%�$X�r������Q7j�CP�R�CJ@��'����D�#{2%"@����1��'Fa|"�|­��H]�A�bDI�e����ɕ��'m`7-3��$���n�����5��0j���
���Q�7p�0��	矈	j�ٟT���|Ru���0��A����Å���4��¤��kUL��A
�J{�0���_�8�ˍ�dŪj1L9�TG�#}֌���#Ħ\��͔�#���v�
�4�ri:*�x���EzB�L��?qg�xRI�#���Jt���h�`sEIM��y���b
�6!��b�-�����O�=ͧA��֠nH�-Id�� ��@�N1�'V��v�`�v�d�O8˧&s>d��dB����e%�@]��H�� ��?����+��ME8X'��s�	ܜ�1b�ŏ���θ-�
x��˓�V�����^�P��:�&��gȤV�0�y9�ƅX$P�>!��2��NU�JX:�(�n�p͹��"��2ؾ��I���S��L�
�C��E0pΨ�
�b��I>���ȓD�Ih%�˾h��E�#%޾J��y��4��tEz,V�!�Z<����Gq:ؘR"Y�0�`7m�O����O�xS�O�!G���O"���O�+��-�� E��)�b�N$eE�#"�>iFC�H�,��|&�02�]7��YrD��(w�.���b�:3�8�r��=pg�֩�+^h�>�ⷧYv}�،-wv�������H ӢQ�X ��O�X ����=rl8�eP���k��8����ȓW�l�Q�B4)[ڙS��2F��'�H#=E�T���l�ٔ��q�93G��;�F��`�OX��'��'�n��ԟ��I�|"S�A_"�9�{-�5� �*_���GX$X��$
WdJP����K1�U�� W�@]*h�=pٚ����s�T5/�ִ	P#�
���s�x���W؟T�d�/�vH-IՊ��f�-#�!�,Z� XE*��_����1���'�1Oe�>���,J�v�'�"F�h�!���� �X}���_�1��'��(P�'��7����u�������h����*^�^LbG�,Ƙ0b�Ȑ�p<A� m�R�J�"�A��,-�4�B��:�p�7�R����$	c�m<��E�8�ACa �B���5'RD&!�Dƿ@�2�U7-z��Y��m!���9�a�Y�L�����QV��8#�?�	0r��`+ܴ�?!���I�%���D���1�d�1�����X%T�`���Oƭc��);�f�#F5?k\�{�Cp�t\>�t�Gzh|��V���c���
#;}�IW6}����$ʭ"�N$��ɁO�hmSG��d�P'~���ӀN�(f&��&AG��ɜQ����N�)��5X�L�%�#���w�!QC�	>�����@)A�z4�m7Y���WA�'|�
��ҍY�l�bH�%��(h�Fz�D���O"��J,){���Vl�O(���O��4�Fl����d8Ps2o�( �eQrE$�	������R�UˈD�4��,H�tȸ&��=WqO���4�'ـ	)b@��o�,x�d*ܽ9Ob�臝|�ܽ�?�}&���ϔ;�`̡Ҭ����sq�&D�0�gJ�{���s�&�?͆�C3�&?��)�'z��E���R�gR��0��wM��(��Xl̜���?a���?!�Q?��	�|�VKœ|d6�q�/�q�� (׭��G<��D	�P�J�aD�'�l���gHf1���;_�}�0�^H�hH'(�����/�1���!\L��)@���&�'v\6Mɦi�	cy��'��O�Y�`\�r2�H���Mk$���@"OJ�5HW��YY$�U	b"���V�$�v}�U�<2���M���?��F�xY� ��K[	_��@8��?�� �����?��Or�1��]�m��ta�NdlY5D�� �
``�֋_,(����	e/T��H�Z�'�
@c�hJh����	RHTܰQ���MbEn��+xh4#'ރ+y����V�'x`�C� z�'�4�BE �������B�3�������4W��͋0��$�BO��o:� �x�@��Vw���nA�B��ID�)�$M	Q��mџ��	G��4xE���$vblx�h���¥�m�b�'0N��nO2L��l�4mE�$��m�|�/��d�W���A�)ծZ_��r��>��,P�8�`��H��{���0a�SG�Ј3�Gԁ��q�c��]��'B}���^ɧ�OG�	g���3�D����.W=�I�
�'Jj4�����Y���x��߫I���1
Ób둞�@��ԜP��A)��5ͪ���΁��M����?	��-�aįԨ�?���?Y�Ӽk��>7��aV�Y�~�~�0��"��y�OrA"�� ,1��'2m�3�	H��hz�eK��Դ�߭�~��'�O8�;�J�/����nnl��g�=�\��%��%]w�x��|Rj�%�?�}&�������4Q��Iͼ-��ePFg#D�ԈK�r7��Uo(*�tQs�4?�1�i>�&��k�9`���Ǌ�4�4�5�P�sҸ��� ͟$�	ӟ��������OX�-9 �L�$kA73�����"�3#�~ �Q�Ȅ@��t3b+F#
D�2(I9*tb�q7�I�̥$�Vzt����ʅ/�j�0Z#3�X�h�A�%`jF�Y���C#j5:p�ȓ�(O�8mZ�G�L ��C�tmR��	J�����OB�o�ʟ\�'��D�?����N*=��ܱP�J
K�a|��|2f�������	'$pI�d[#9�O�� d��]�'Llf���Iɟh�EZ4%A#0&C�fX��e�쟴�	89:�	ןHϧJ�!��A�	�`J����r�,x1�/YNJ��D (P�O��!���I��1�5��	�!��'y,��jE�'G�%Â��a2k�_�*D�
�'<.i���<m�d	�1�Y�@����'��6�?b�05bU0�ȁ���u�1O�i	��ĦM��ӟ��O��"'�'m0�`��s���I�$�54��w�'6��Ƈ2-R�r��B�AfJ�I�*x@�.�� �c�(]t<
����4"[t�'������ˌy^|����]��q��H
�"ռ��OJpuV$P98 ��hB�Z�0I�\:���O$0%��?Ak���!���r���^{��3�7D�H����'�~�c�(s]F�q��U���T6�o��s���(Q�L����̋��1��iD��'�"S�T�6�ZW�'���'b�w�&�d��A\�]a�<!�~��4X~�P���S�lȬ�{B�ڨI�1�f}r���y0u���HB*�*Q�H��	߮m����D/����%��8��6��B?��Q�'@��p ���*ݐY���x]���N9�d�xY��L>�	�%̢A��ʛ�VӤ����JB�<3o�3(�h ��"�6f�rr
��<���Dԑ��[�)��X#� �&lt�RAg� S
X@���XRhl����h���� +^w���':�� O���ӁʆE���i���{(�	���;rd�06m�� ���e;z+� Ҋ�D�;RH���@B� 0 �]8XQ��'�Y�lP�d�2�A5��c
A6H���d��[װиD���P�@�Z�x�	23�'���T�D��A����Id�ã�yR�/q!�T�����}�p��I���'+�6�1�S��H�=c��k��W>x�X{�̋��y�@ _y��X&�Z�n�`�b�L��y���N}�e�5Z%�E�W$�yrE�ԩ �	L����D^2�yB�I5�6�;`.�����#�yb�ۻw��(��	&�0��c��y�kIt���D��@�sQ��y�GJ�4KB��4�ѣz*��r�	��y�*X U[b��e%�=�%p�� �yR˕ 4���9�͙j���&�f�0�ޭiÒ�K������;��	$�M�	�L�;uh.V�1�ȓ j����'G���8��ȓzh���daR 1ِYѱT�bJ��ȓ	��9�n��E4�蘠�5+|��ȓI��C'+S�~h�9�K��,�d��f7��1M�<Aބp�nǶr�D<��u%�+�2+ƅjQ�E0./�����z��˧~K�	�kF�(Q�!�ȓv�X�s�13t�q�3K��	��p��j�Dz@"�
���K�-
n�u��:]�@�a��e#�x�+C�;�����G����%�ƭs�pp���2�
<��S�? ji7�^""/��(�ƛ�2�й��"O�]b@�Xd$Ń`�K�1�	k"O�[��
�7}�ix4�ɔݎ!��"O��b�LZqE�P`al!_j	aa"O̐C7)ȇܼ���q80{�"OR]�ঞ�7dB��a	�/U���r"Oh�i2(R�J�\��Q*�$�Nq�g"Oj���'��h��C!D�{|�d"O��Zp2)�&�J�Ŏ4�j<�'"O�l�ӣшs�Z|�4�N�#@��"O���B�:�>x�0!@�1���{�"O�}a���Rg<q���UoRd�v"O ̃uh�;�T<s��D�D�X�T��P���/����\��ń&����Iժ���PB�'�z�����pU����E�6eO��z�	s�Mp�L/D��� S�{ް����!@^��t/2ғ;�L����/�>�0�gZ�e�Je�e��46|RR�:D�jS�%+��M��ӹ���ेk�jТ`m�Iq�t$�"~n	�r��CYJ�$��uC�M�B�I:_ ��됈P�ex$B��� T�j��蟘	dZ��Q4�:@!��~Fz�!B�K$N�*�� Vn�DӁ�>	p� �CK2E�ua��0�J�h�>
V��qOJ�F9
��D�vψ���h�b1Qa䝒d��Q��5�d#=!"��1��2�FY̄��Յ�z?�e��J�A�b��GѸȲ��R1�y��ub� ��<�$�G���?T/�@��Q�'�Q�!�Y��e?����O^�p�	�Q��C��2$М��"Ole �����#�&����@,�6�����On1S�_��	�?�t�̓���f��{���d��P�Y������z2x���R�y*L%���?�Xg$ݛ6>��O<}��X�w�|7m�*	��z��?�I�c��;���6pu�$��Z�G�d"=i ��"�Ɯ`gk�z�� q��C}��� n��W�	m�pѸ��;G�H�Μ�>���Ҳ�'� ��vj�7Ih�c�I˟4f!��4RVN���.�0�6h�7����@F|ZcB8�	:"���*�&�C���A�'+��(�%A<u��q�����z�@�J��rܑ� �Gg���<��k����՚?�H�`Vs��Q2��z���7g������b]"o,�9i�e�r�"�*���Or� �%jo�$��
��vض|�T�䂲�$H�M �~-(�A����������%%��H��+� }ZQp�'?���L1A��I{��M�"�@͚2�"J��B��y�e(�$\O|�2"+�J��1f��*[��0�v�Wc2"ɢ�ɚ;#�����b�/gџȺj�(T��	�c`׼�����]r�<��M��y��� �zX��G+X��$��&�z!�;q�(��ү��y�Dքw2<���x}���2�M(�p>qb�۴w!�=�1)���D$X�.�8����M#pL�(��]�ː�?�$��eܓ}�"V�U�"�n��S�vaREy.U�?�� R�E�b
n��C��'���;����&r吀�N����P Οj��e*G.I. �� Μ\��i�L���a��h��� 'ήH�0�[<~�1xZ�JtsW��Q��̧H3��a�Y��}5�Р�͋�'�ȡY�K��s� I�K�;}�������e?��,�' R���FO�s|"�ݪd�������� х�Y�B����tM
�r`E!����7Jy��:�m��?�<�k����?2�4C���)Њʗ��!-�O@����a�@��S���&RR% ��I�D�Ё���K9hB �����5ͤ��W�ƠR},���C17} %�剘 1�j(��B >/:q��'�0�G/I#5��\�S`� R���qә0t�5P�C�}�F@
&�ݞ\�ў�S9v��5�o�	}��li&�I�-���a�'�r�!G�9�P�ǎ+d�H�R�!� X�d#=��c�����	R=��ݹ-�t�E�	%��T�e�-_BX����a7|cqfےE���pc��r��Th&gҁ[ü5�)O��W���	�n��@V#;98ݚb:�����H�$y�ia�MK%h�剖!)n��@�9B��ke�]b��'��$���(qN�%)�Ń6��Z�d\ �?��O��<)c'���QB�%����
TcDi���M�U��Ԣ�̑L3�QB1N��_��5[��]*K�oz>��?�	���4��'h�]��׏L$L��e���>�l|�2����0?)ףݎ�ơ��
/��	��fI�2����������_���n�D3z
~�[���O����,��5"E@3#lH�/��
�IL��#Af����!���82s�H�_�={H��W��R�䎡P���ߴ:�:��]w���=�H����M� $|�wM�.hv")��-^d�r�qQ�Ks�*H��� P�EPKK�hH�X�$l릮S�5W�4	c	ƒp��hȑCӔ.j�'aȓ��:$Xw�Z�p`-�'���A�1%Ӧ�̟aB-�W(�-^4 �W��-J��",`��
�$w>�bǤ��u��������@����^6�j�ZD�<xɸW�M|����eJ�yaA�-MrȲ/	`�(@���W�4ܰ�,�l{���O���Q��H 	G	���.�"�0���@�5��r���L8���k#a�֩h�wP�|���˰CX��1MP���]��gy����jmHrM|�}����`yJ?��1�H9\��G�1;$Ȁ��V�@�2ᩴm�$ � �rQBFD�M֧��ܨP��"t�[)2ѫ�l���M�	9�Nuj!Q���(����Nڧt�)��Od�"C$�<ȋ`eӲ �p|�C� �2E���sӬmX�	�O���L�`p��$<�X%�LkJ�dB	y�����`�hCeAѩ,(  ���	J��鑢�>Z����AUg� � Gk��A��O�`Sq�;�I=PĽ� �
]�lz�Ú�Aƴ!�Q��=4�H�iކG������tcI��KU�H�i{l���7;����ϭU�嘪O��:��ub�o�;Ct��=�)]���9ۧf�7!ܲx��DC#$��� +�&^�:P��Q7ȋ0.ټez��a��Ʉ��m��I@�g�t �%�V�=�V!ߗi������> 5$�S��M#���`�w�Y-%W�!� �ҟ�2��9���Pv�J�� #�<�����fi��A	�	�G�+BF8@�O�-
t@�z��Y4�1O([1D�<�ZG�5=0��:�ˑ�U�$M��郕fǁ��ӊ����c��)X7�Ldw�)eSC(Z�@	0(a��
H�	�lηf�:���w/�0���@�}ir	Ɂ�M���՜V�A�;@3>5��<O1��|��z��i'dDD┰��ɠ,���t^a[�! _>u����Xծ�B�"C�JX܂�fM���Q�t�2��H��#|�'7N�{Bȉ���pSU�T�V�\h�O�����r&
����Rk�O�N�y�H۩Z���aT��0��0�a�����A��;�\�
�%�0=�� �ur*��!��[���&
��[���h6�	�y���S�)�w���xF�El<����c�2.�7S�����-V�8\�%m~C�(����z�J�`�{ʟ8]�!e
1>ô)��4�Z5�h�)����.���i"�I�-��� #�S�x��Iv���M6x2��r����ЬI���4��T�i�I�N�@բ�٠~�Kg>qA��|��Fhna2aʮsp��(d�H6��ӰI�v���EU{Ĳ�j�At7�i>�y&J�{7eĳJ�ʥJ�9O���c�D�7�F=���L�D�J�q��'x��1�7dt��#�#^x|�ȄO��<AB�'5bMr�Ƌoo,%��^'9�ĩP+&LO�pS���\��U��	��Pb!8� <���#N���"��'B2Yr��F���B��Ҁf�xܓ�m�qt � ���-
9�b���v�R�g��\�uGV���Ѓ�8��R!`�a��΋�*��t!7E�����4��'R���@�4���7I�L��N<�c�	:t�4�A�^�i��$q�)�|暡A�BPD�d�R X22=G~Zc��s�M�
ca�5���?J�>Њ���]T�2�L�o8`��P�3,O���ݩ"�6]c�$@��X+ߘ�Px��L�0�`��'��<Ϝ�㗍\�)���M�'����B���K�c��A`�K��a�K�,@�Dd��z��3_��e����d~b��V�F�&�K�-^JąX�}b��21�����J�Z�}�öi�'0Fr'M���	&�/��1�bkE&#`� �F�0e�`,0D-��ɯ @,�z��Y?O30��S�H����wk���0z�PL���'Q���*�=3�X
7�߆���hM�1,-"�1�瑅0C�l��Aٯ�0<	���!Uc}��)z�J�c`fB�@,���^G��l��Ӊ�C�tu���
X-%���ƿ�p<����/k�`�J�<��!�DH�,C��J�@�?O�n�@�1O�Q<�<�;Vn�B������<���kU(^�-D�s7�$�6bO��gg�����M�q�'2����ڗi�ZiXb)��)3(� �4�M�J<��YBt�xB��-4-���Ǵ���&�CU�͵!A��� ۭZdNm�gBU�]L	|����'����";u�`�,Y0@?�1���=W>,�Wo�,N��k�,`|�q�1��-��Ũ���mƸ�!�5܌�$��G{��d�L��q�)��Gw6��r&�'J&�%kǓ��۰�ڹx(�]�=fp8Y�0}b�@ޥ,���a��'r.d�+tE��{���G$!�wB��8�N5�����'�4�C��F�����))���9I<��KM_$�����7;��4����b�'y��Q@���n>Hu{@��/�Ɣk�O��q��{�H���D�1F�|8��ެP'ZM�#��9��a ��cyZ�ON�@ŃL�m��S�w�����X���69N8��u���z�x�P%i�E��KH�!�"~�@ݲ�D��t�,z��+!"�<��C�#!��!ʦ�'}P��@@�/k�w��(���2F�\��AVy��M%�\��AF}��ݦ���Ӻ����478��89��$	���ļ�ጞs�q�l9�Xc��,�>�H�:N�A�{�? �Tr�-�J� I�6~��0@3�xB�$-|�6�,iy	j��f��Oę�oF�:w�0*��	:f�i3j�>�w�A�mN�3�D��P���3;��'!7�_�E���E0��׋��nA 7��=�b���M�1}a{�G׮2����-�4�����"�HOp�cG9;@�+NQקu���
va9�`������%�y�E:2w~��ե��xAR%�8�?!w�����j���S�Od�e8R�,Z��zt!Q�-_�h�"O(="@%�)�%�$L�2F����"O��P�y�¬"��W5&��b"OP��0�*"U
�:���S!�Yy"O�HK'�{~A��ϻV��c"O�	ь
9�� x�;_���X�"O<�`���'�-	D��L��2"O��$�2�2�V�\$���"O� �ŝ�=�Px� �Ǯ
��H�<ѧGuJE�⥛$(
�`���E�<Cf@�3pb�(�n��@���y�<i��\�x�z�EN��[�(���o�<�d��`.��E�NH����j�<��冏Q��l�3dĀu�&���G�{�<-�~D���9gD(��,�.N�C䉪
 ^i+ġ��=j�l�go;HC��Rz��R�ے:,��"jդge
C�I�H�\`G�Z9J4vP���<O��B�	��bQ�sLS�9�P�����O:C�I31O8c��ʎ"&��)͙wp�B�	Z%�|r%
�h= ��kS��ȓG��`�f�R.0�MӳLE�6���ȓV��@"��A;�PI�$"�:"��X��#8Zg��%�T9K�,8h\�ȓPI�ʩq���2� @�xM�ȓq�t,b��O�rm�
�x�,��ȓF,�̪CE�-2��!E��,ri ��,��0y$L")A�!�A
����8ph֧ݵ&��0)�$x
X0��9�r1�E�OA��êO�`��]��Q���%��$/�np�u�^�}��\��P,�!�f�m�x�IĀ&�j�ȓs�Xm��œ#HЭS��U=[�ڽ�ȓkq���/W����3��4?@�\�ȓN�4A2�@�X��q�I�x�i��{&��[�j�Z΀;B�I-u#���ȓ=�,�q��'d,�!Z�1����%!J��r鑏D.^��t���n�0Ȅ�|� h��ַ`�"<�&mǹ&���ȓg
|<�D��,���!��_009$���(�r��V2W�x�ujI8C��,bI*,1��
Q��8���L�C䉋.�м���ڼ8�
��UFS*7�C�I�&Y"��V\>��ӆ�%�C�I;0��-ͪ3R�M�B͖?�tC�	4 Բ��DHs���"H�
�dC�I�:=bul7EH�Q�4�qxXC�	�<預d%r
���B2@O0C�	Zl:%y�ܩ(���؂�J6pC�ɬ
_0����S<����."�dC�	�t8�Q��;,6ls�G�gNC�If�(,�N�@L���;t#�B�ɞ#Q`�Ů?0ԩ��5��C�	�V��V�w\  �$'L�bC�1X
X�S�TP�
�1��ZC䉔OН��īQ���&BL�2C�	I#6�Q�G�.̬A!�9,^�C�I�\p���ڑK;�1*aA�^�C�)� �PI!�J�r���fۣzkb�a�"OL\i�J�|�)�7��(&o8 CC"Ohy:���F�&M��m�$}Q`�t"O�h+�V�W��p��,J�"Ol�0%Z:��$�5&�(hF"OPb@G��� I���%+�"�H�"O��Bb/R��(���S�C��P�C"O|���F|�@��r�½9c"O�|PF��
0P�5�d�P,WrP���"OФQBӂ ��q�f֬;���9S"O<�KՁ�t)b$%Ly�):U"O���P�I�NPSqC��Fx��x�"OpZ��G�|����CBEv�s6"O�̛!�܊~����� W.ڇ"O�����ɘOuy��G!HT"I� "O�9(�c��͹�̉�sܐ
�"O���C^hOT@��[�}4`p��"O�u��[�ՠ��L�����"O�%hP�"pL��Q6R���q�"O:� Z9pHJu��4Sդ��"Or��U��4z���ǌ�RΒ؈�"O"Q���$B���X"GV$[�H�I�"Oά����?A/�I�u+4cEJ���"OREI�Ŝ\Pd)Z�U�$���R�"O�ݓ��W� Sj�13:r�"O.Y+B��<�bM�!	 w-�P�"Ov�#cbh}i���o�� ����a@�>a!�dQ���()���
L��=D�X[A�
�6�h�c�W�.����9D��:�́-�� 鰢
�ZO�����6D��B��#8� ��Ŷ ���0`N1�$(�O��`�NX�lH�a��_4���
O�6P�<��!
����H? �O����Z�
�8�ᓈQb�r�kAC��ax����e@l� w6)��E�C�B�H��,�E�[A��E�C6�n�>I���+
:R2�bn16��t�d0!��W�)斬t�Ǥ�j��E�0i!�$3}�B������K�`�р�ްj!�$�/l��K��d�\�9=6��O����KY�4��׽3ڹ�Q�˘8���󤹟$%�8p���t4�	�2uҹ)��<D�Lb����& �1����.:����#;D�$#��5"�	S��U�Q֬m8�@+D�T�6o�&z7�]� �!x�~u�-}��)�S*�xY
��r�Q�J�S�B�F"ب`Bk�$xP� �e�VݖB䉃%VR]��޴�<�P ��(C�(B�	�W�����~fr�'�����<
�LF�I�� ֛,�68�Ê�J�����t�\���h�$`	g�Q�޽�ȓ��:DJP�r6ՠץ1;���ȓX�1pd�^1B���X�vf��ȓ�
�����U��ʵJ��\�v�=}b�>%>㞴���G�j,p�ʐB��f����f�5D��a��K�i����d�ѾH�VG��>!�<M�]q�]
��q����"�Ї�IG�'_,���5NZ<�+`#(.eBu��'��!B�ЍmY
�sd�G�&+�=��'���h�c�1�j��c�,5��p��'"� �.��������2SA2�'�]��?$C�@��/��"��ɣ�'E�}ٗKT�� ����&�쭹
�'Ŭ��&l��3B@I�"�v����� T�t���B�Q��%��gD���@"O����.�t�"�Ǔ~O�P���>��'*1O��<����6)�Ĭ(�LF-)��kv�#�Ln��!��1�M�}�dql��%����k<�c!U8�����E K���sd	�<) (S�f� �Ti���a�Ձ�y�M7N�����
�J"���Îy�i��b>ͫ앐X|d҅�H�X����#`-D��@��	O9V�؃-�g�i*��/ғ�p<Y�JS�^�����åg�0!
5��`�<1�O6��̲��Fo�B�Б��F�<ᄉçO��Ez4��o����$QX�'_������2.W*!��ʶ�4s6��W-�O�<1��!!J0�����$u�@a�'LG?I���S��(�c%�A3����ťt�dC�I5s� zJ;&�$"��D�w^�C�	�Qq F��l��q�2��6��s�7D�d���nɰ�d�I�cN r�G!OF#=��@�3��yF�xܩ2F!�}�<	F8	���sLǌ+!�B�
}�<�4��m^8h�n��
�<?�C�I�%�A��,���>����S,̊C�	.Mذ�!��Y56��P�D�v�^C�ɶ ���%"�����s_LC�	m�K�f�Q?:,�d�ΫdWC䉸2S�-��Z"�;0�2��B�	;j�z�!S�E꾅����s��B�]QwkSNpp�гQn�?��4�(�x͋��_�!:C�NPb�m��"O�D`f͍���q�#RWB�Qf"O (�N5� !RG��R�"O���tJ�M�쩳���94��"O�hy���d(0F"ES��HR�"O���p�P�$�J�H��}���"O��:vi��=�̪��������'TDy�N�5.��<�`
�;c�&��s���y��\!�4nT6-%�u�eGM��yR�U"d��iQC�ӣpGJ���Ɏ4�y�(7 ���%j���q��y2���=n楲�Nȝ/�`�E$�y�dښg�",J))~�XP��y��A>��s1���r�T0��Q��yBf�^���H�<�n�⤛-ld���%��;���c�@3�X8�B���	g�dΝ<T����ְVcd�$��1!�$Va��r1��#�(Qq�#	:'!�䒬@pd�qg��{�,���:|e!�dE�~�6�a3��#��8:���y!�D-�R����ޭW� �DO+@�!�ĉ-^�I�o��O�j�� �� �!��e�LCᯆ�h���A�DE��!�H�]�����5�~XB4�äA�!�+L�.8�q!C&04y։�1o�!�Ā*|G��g�D92�M���J;N�!��1c~5�5���Cv����1:c!���0�x�Xǆ�,i<�!��Y^!��!L8��#���,�0Q��(|!�Οt�FQ˕��]�D��H�����	?e�"����|�~�Y�IǪ?��B�� ~?f��O�F2��r��hL���E{J?��!�86���`#��:�`�)D���C��4�Zq&��/� }�%,D�p� �؅=MNx���iX��A�k6�O��]�nD�yf� i�C�z��e��S�? �DYf��2B�9��8L!��ё"O���o 9A,��3ڸ{X�R�+-D�C'���x\6ѡ��
v�@�"E(�	^���S?b���G�I�2pB)�d�7�.C�	�C��T�CCFsX��6F-d.C�;*��P"#��!R�����o�&^C�	2WXjaY�IxA��D�&k�C䉼@!T{��	1�Rՠs����B�I�S�%�NC��~08���*�B�I5Ue�e+F�'	h�3k�.�.C䉍f���wJ8��C$E)G]C�	�i��֋P�V�\PX,G�i��B�	�p�>�`S���lo��P��JPJ�B�	8*����f����a�L�-�B�ɋUP�!�#��I�h�$�$
�C�	 =��y��	kJdɁGU"b(�C�	����3�6U�����\D�C�	z#�ڴ.֠)m�i��C���C�	��]���po�$���a]��
�'k�b��%�����f�|t��0	�'^�|aD���Q��@��&t�q#	�'���[􈖒{:�"C�=j��@�	�'�֤�� Y�f}��"  _�`� �'Ũ!�Ǡ�˪Њ��F"d��Ġ�'�5�b.j\R=���% ����'��Q/X+%[-�+Y�;�'�$)
T%��{66	� �Z�]���'�`���̊D4p��f8H)�'�mꕤƑ ^����n�+z����'�:���Յ�0e�2M7��"� D�l��ɖ<L�0&[ a<P��R=D�<�&kJ�}`!�cex�	� ��yB��e�~E���`���Ц��yR�F�IdV�s�ꂀY��R̖$�y�n� t���H�W�` JQ��y����1HޱU;
= �V��y�nܯW.�=�Wɑ4S~���C��y��9d���Ã_#BkldI�Ǐ�y��Ν#�@)c��4@Z�l�T��yB�Ŷ Ңa�G�̅=�\�p���yr�����eQ5&G4b�� �7d���yr�8�X�)Q��m:*��V��yjG<#��������a����b��Y�ȓm�8=��A,_DD���V��L���l3�����E�2`B�ȘSL���fQ� �G$j�r-
�i
@� фȓa%�D����*#n`8t�ix݇ȓI1���T�Wj�<��f+_��M������5h����c�C)	�ԅȓV[�a��H�$[��M��D�v`��s,�(�N@[!�8 7](r���c��=����h����N=4@�؆�n�*��n�TG^8H���{W���ȓBS���U� aIriɸ-$��ȓxz���T�X��Q��8"N�݅ȓkt�8G�*ok�qY�]�A[�Q��#�Н@c�����)�K�j�9��R�r��u��	�J�81(�+�U�ȓ�����&oz`i����}��-�� ,X���ʜ�S��;R�[
d\D$����y	`�Bwu�uA��+d<Ї�K��p���8{g�4q��(b~�͇ȓ	�"Qkæ[�c��8�ۺ8rnA�ȓ
��4��BP��n�p�ͶU���S�? ��ٕ�*ND:%!"bQ�[�T���"O��!�2�iy�@G�B����"O�l[����a?f4�FMC�@�� �b"O����H�Kl<=Av썿a��)
�"On�Yǘ�~a ��J�&��a�"O� �f	�F��@(���UJ�v"O�<� dD�ẁ��rj�
I���Pv"O^��QS�H�5B3j��l�n�ib"O2���O� �Y�򨖝]�b}!�"O*��Bk�,,��drW��9��"O�Eq�fE�"D%"7'͐MX<��""O�x��nRsf&M����'J4qp"Ox:W���Ƹa�=h"O��ы��f:�5-X6�X��"O8!Х�ʶeu"T�&��3>i@!"O��j�"4��D�ҁ;0@�s"O>�a-�M�j�� ��l.��"Ob��� ��T�TjI]^i��"O>� ��ع<���Vi[�0&d�"O��$#Yʸ	���Ӆ? ���"O�=(@[�%0؁y��@0�À"O���b_�2�����'�zh�"O�H���H�����"3�8h��"O,u��+V%9��@�0����չ�"Or��'�!T� ��:Iw8� r"O
鱣A�w� �@��cv`-�c"O��Q����HT�8ak6ك"OhQAA�,+xI���^U��"Od� �թ1�6� �K�XE\�C!"Oh8r��O�`�m�`�M�C����"O���r�,6^�]z�IO{٩"O҈ҥ¾<!je"�N�2>�ر6"O����U�af�5����-$�ɱ5"OPMʱ�^73xT`ɛA��"O��`�hߪ#(���W Q�����"O\��  �}����T��H�8A3�"O@1+u.�7bzY0�G-|f��f"O� $���F�J諁�u<t�u"O�X�G�$J��������:Ԋ$"O@ IR�~l�D��C܋�$�R"O�<��J�gTf8c�K4ڤ��"Ox�C��U�5%�\bwjN|�|��"O��	���~�PB2�D�6qj��"O�� P���i�E��$T��R�"Oh���)� sEhC՛c^P�"O�IaX��m���ޅ,��:�����y��1�%񄨈='Z����&S�y����ބ�VE��$3�@�v`��y�Ήf���� ��i#V�C���y�E�(�5�gZ�a�!�K��yҪљ3����b.�7ch�@����yR�3:8s�f�-dņ̃`C^��y���>02H�QF�/a����O<�yB��&2pv�J�Æ9��T(�D?�yN�@n2��,�*~��6`�yRa�<~�@T�G-~9���%F#�y��@\6|�J�$}E:�ReI��yB�8��p2�G�nc��{$��y�ˍZ~��Hg��3��(��E��yRl�&D������.1fe�f�y�/
� ��`��=���[��H��yR.�N����D< �y������y�+�$Ц���Ə�A.�ہ'�	�y⣉&�T$p����l�L	� �%�y
� `�JP�@X�x���P6ؤrg"O ص�J�'&B8�͚(+���"O�=1w+�2x�jXqt����p(r"O��pg�S�4r6	��wy��"O�%��ņs�<Ad(�.vdP��"Oи�g+G�rt�3HU�~����"O��z��G �I�e�/ ��1�b"OLؠ�4y|�x��cB��m��"O�Iʱ+��K>��#ë��Rj��2�"O���F-˄ժ����( T��"O ���������N�sQ��Rs"O�H���8֨VI�$��]Q"O�MӶ�2\WJ�"m�*���"Ov�R�U t
]Z�H�ׂMc6"O��®E�x��pfAO&� ɗ"O�BD�M�T%8�@�O#&9҄"Oh@���#4���!�"(V��"O ��@��,/81�V�]�K�B�ag"O�T��@�s������<L��ٻ�"O����LG�� �R#�1��]+�"OL�
��\1͖Is�FJ���g"O�eɗ,+)�$ �F
�,t �´"O4EA�V��U�uƀ'7Z�U "O��s�G�t�3`%�/X��r�"O������gw�9�
L�g�L!۳"O$�+�"ڜM\�p�#�Џ8��aA"O�Q:�(�v�m
a�U�WԚ��q"O���Bךa�h%0%T[�����"O��q�%����т	K�U�F�#g"O:幅�S$g������eUnp�"O�	A�� Ɏ��0 �0S U"O��f�3��ꔀ�~�ؤ"O�Y	f*�7��w�ӘJ��A�"O�Dq�����)(�i�"OH��Ӭ��~�p}��<C� �U"O���5�غ-^D�0��\�ιɒ"O��زlL�*����B�v� <H`"O��§ 9]�LT���O�Z�Va"OQS@#�2�ѧa��)s"O=�R�^&9%�L��oVn�8�	�"Oes�s!�����o�H9c"O(����ZH(�����{"O~0�6�B�*��5�%�Q���(P"O��8��Y�rH���,�#{n�"O�ܳw�R!yoR�!���m���F"O�)qC$	�j��v(ܜ1�p("O�I	P#B�x�|{��:|.lɚ!"O(uQ� G,R�H�����~%d�C�"O��k��[� %th�FG�f�R��@"O
�BSi�G�K1��=}�\�Z"O�`��'م�N��	�'�ؔ�"O�)*R#�8jh�8.\���"Of�7,ѱj�����O�{%��"OP�z֍c* �1��_g] 6"O��k�	�Q$qs���tD2e"O��*��ׄ|d�RcF�YH����"O.�����Rw,d����$<M�"Oj���0L�p)b�WmC�� �"Ox���о��A�ӯ�\AHѐ�"On�p��ƚ�Z�aGH�5P,n��'"O�M��!r��%����~���9u"O �B�<a^�8�U`
����"O��F/˜@|�p9�H�=g���b"Ol�Yc�t:Ҥ+���}.��d"O� d����N3G�8��S�-J]��:�"O�[R��!�hH2�Ŋ��x�"Of4�E�+G�f�����Z�����"O���E�2(�@TSu��<0xB�@�"Oh�/ߞ^x�𲯐���u"O�y����h=d[��	�����"O��Rւ�@}L ���A�D�S�"O��cÔ����fX�Byι�A"O����燾Q2a9�Gc�ԥ��"Od=�b�K�*O<��(ϱ;Ոӳ"OJ����y��� �G^��<=b�"OB1)k�|3��b���E�� V"O4�P����J?*�@s��~�\Q�"O\=0��E�}) �9X��4;�"ONLC�.O�'O����#� Q8���"O"p���ܙ�l�T#H?���SW"O`M7�_�ޔ9��ٚ��@"O�`�ի�i[ڑ�%C�'M�	I�"O��bS�ʶ6�$Caမ`�8�"OL0I��B�FH�����]84["Od�Q͊�`B�	f��
v#l���"O-sf��#c>ʑ�R �+J�4�0"O�|I$!#U�e;b�\67�=B�"O����{��7��]��,b�"O̼ag=}�@���T#��l!�"O\#���X����EcH������"O�-���N��1;�kD�f���W"O�(QJ_�}�-�#�W�Ei��"OL��ď׃]�l̐q''\Zl�)@"O�ss
͈hb���͢S>��Je"O�����T#%Z��C`Ɇ�6 ��"O��0�L�
��'ח\�v�"Oࡋ�٠'؈���a��OH*ܚ�"O�<0��v�~X[�/�4,]te�G"O�9���L7���n]�i>�"O���3�$��D��?$&�P�"O�yJ�L͋,��]�B�	^�2�b"Ox��#݅2�h8ۀ�G�6�x1y�"OfL�'��9��̪�ѽY�p�0�"O�t�R�ǊWjJtz�@��?�18�"O`��dnǻ���"ϓ;��q�"O������\Y@]8�*,R�"OD�"-8w�� �Ã\����Q"O�����W~ƀ
�%�F���"Oz�c1Cөk |@����I`"OȐÖo� ��9e�F�v�ƽ3�"O�esr�'b�����+M@8q�"OT�3E�Pu�F�JqI0�I�"O��j�����P�X/`E8cf"O��� >^�0rGoD67d���"Ot�c�n�9$��I0.�rڐ�D"O��tjL3x,L���/D�
t8d��"O��Pc$!B�r��N�t���2"O��`a��H����ȧsj`9�"O�=��D֤(d�3&��\g�8��"O��z$�ߊE�>��Ћ^�$"OX!�C�[�(ӺYuK�<q4���"Onv瞄��|K� �8"p��X�"O
Ճ�ė�9V:��4J�oBP�"O0� �O��3a� 2�
Q 	pb�($"O���I�C?j<��H�U1�	�"O %���@6>k���f�.c��S�"O^�2�K?>���O�6�A)`"Ol�Y�G�&r^��k��J�q&���"O� ���#k�w��z�
\�up�(r�"O���kc�L�u�KIbx�A"O��;rg�5zǲ�x�C�Zʦt�'"O.�A͂�N(����M/�� �"O �s���R�¬95�ݓ"w�m��"O�0@�	I�eC����,!t���"O���sP��^�A�bD8-b0�s"O������ܜ� ����E]H逆"O�I1*��]��Q��oV�7�T�C�"O�`��;V�Ti��C<�(���"O�E"�A�;$� ����@����"O.Xs���3�$�ˑ������E"O����h�L��{"�߭Q����f"ORe�A�� b�B
4sn8; "O,([��ȿ@���J�0q@�"O�ty��	bc��Z�N�Bb�1"O��f�mB`�7&?�x�`d"Ouٷ�T>��`%"~����"Oν+CdJ���T���аo�b�W"OJ́��T�z��"
\`���0�"O*A��רt���I�+���F"OԱ�r��	?�r�a窓�kǬE�R"O����w:��0��G���k#"O`�r2-�{gP=�����7�*���"O�����^�3lʵ�¥ܠ=���"O���a�TH�z� �m�&5�6�C7"O q��&C;S�D(��	+*}y�"O��Z��Q�K�0�I�j�%`�:p"O<�)v�&cģ�H��R0��"O$�� �Y�m��(k�K5����"OF�y"�>��)E�O ��2"O�h*�)
�W��xc�\+B}B��"O����6+�hqU�[�Ppډ��"O��� �����"̟qmpa��"O|ڤ�Eg&��V�V=u�ڜ�u"O*u�����H ����&GT̈P"O���"Hݎ� Y��� ��m�"Oh����P�+�$�*!����"Ozй�i�B+���H�&e���d"O�S @�E�X���j��0�"O�D��	�
:ei7��ph��9$"O�<j�OA.3²$�P ;	o. �"O*%2�Ę�R�I�� k� �"O�Xh��?�j	�0�D,<16�w"OF���B:�`���BW"#u`�`@"O��Q)[�=��i�$��g_r�'"O�"�ǖ8+���1d�>C�����"O��K4b(�.���@M�U�H��"O� �l Mݢ���^71�<4!'"Oz1j'��;vQ��.�	;���H"O��;�-A'�e	��&6��`�"O�ـ��� ����c��}{�"OZ��^&a�V��=�V��"O�E*Vo[���eZDϒ�<�ɠ�"O�- Dc
�J�XC���F�H��'"O�y�bV5Q�\�Cѣ�Z}���yb�	&F�*��Q�;XE)VB��yB�
C��� 
�2к���y��:C�\�%lO�{J�-3�`V1�y� .Sg�����=)Dv b�J%�ybC�!���QI�$�TH ޺�y��ޢ[�H����R��^��Ś�ym�%D'F��9%\��"�Ӌ�y�E��+�i��~�X@:��?�y
� �ř�c������E�*˸��D"O��`�F����e�Q��e5"O�=�fń"xz6Ă���HȖ"O����Á\5� r'"ܦ8�h�"Ol����_�tEz�R,C���:�"O����!?w�S��يz� ��O�Q#􃑿s�:��U���EO ��%.D����0X�V��c��1_X���H'D�4%������UbM:Dob���"D���ċ�j<�da��J6 N|�(=D����Ç�z��M�WlG�W\��6D�$x���E��)
�8D�죶�L�n�B��COF�5�X�q@64��XĊB��0�$�9�1��_k�<I%Yv��q��ƌ��L�`�_�<AƆJ"jp����V����^�<Ae��x�hAi�&J�����X�<��I'$:] ��� \��7.�j�<a�D��n�\-�&�� -&B5[!�e�<vMF�K�����b)��gE�L���͓���dɆ�Q�� yWT��t�ȓ����rKF�bm��nǊu����/)�4�5F�B���p�C�\�൅�bXx�R�UdW�m�b O5f��ȓZqh=k��@ %J�X���^�<C�	��N%c�삖I�����@��C䉓3����ac�z ���-Ñc��C�ɴ��)�RC�i����J�C䉚Z.P躱�:"�L��)�1��C�I v�d]҄�- ��\)4Ƅ���C�	�W�P����*%y���O�9I�FC�	����x�.�:�:)c�L"C�I2 �慙�$ �ec���&��c2B��3e�X���ݏkq��d�ɦ�\C�	�$ 6�R홻 E����M��mr.C�ɞo��ґ/!Udpй�fؕ0�C��>u���־e����E�q?�B�ɕ^];�,�B	��%�	�B�I�,���Q�bU"3rb����,$�C�0=�8=3���=`2������`�C䉱;�"���]��nmj��P�Y�C�	,2��iЋ%�4 �%��B��P��֤�-�n�xc�AےB�ɠA���2nWw���cA�m^B�ɻX!��⎺��f��il�C��yB��KC�%O|��aNT#.B䉌5�}�$�XV@Llځv�� �ȓ.�����62Қ�y5EZ�FP����k�	�7�à_P�P�M��u�\��W��xc叴Q���(U���m�ȓ=�b�cD"�>%Z���??:,��2���l��m�����`
�-*����wX���#f�hP�=h��D�ȓwj�eIÊ�F48�;R�Q�]�^�ȓ	m,=Ss��/�6x�B��5MHX��g���3����D;�i�9W��хȓ,� ���
&:G�r���2_ V���a����� ,f����]% {na���q���+��ʆ�>���ȓ}|
$�$c�72� r�+yZ��ȓI��U��9!�<�wa��o�ʔ�ȓ/{@��gG��b�d��'ω2ncƤ�ȓ�f�P4OԿ_~�}r5�M�5�ZP�ȓ����1#O(s�p���-
�=��S�? D��\�"�y�� R�2xC�"O�e�7Jz�� a1�LC�����"O�9e	�*�r1�ą��b�^�"O�;���zh�E�a� Ųd"O�x
� O�b�@�isO�������"O>���&�/`Tn���л�*$i"O��4$ǀg�ޙ��Ú}�@ܑ�"OP�#�P�ie������'tVh���"O�x���	�l�>I�$Ï-M��x"Oh"c�.Tt�TB�k1z��!"O��xfC�`>2����I�c��PzA"O��p�!R>�B}��H͌:��<s�"O�t�']$�Ei�hU(,`�Z�"O��#��
1:�~�2�	A(o�y��"O0�ۑ:�.�wϑ���Z@"O�f�>&V����G�$��P�"O4=��_){Z�,�E.SPPTq�S"O@�E.C <��U���W�s<��A�"O�9�!oQ�Ը{&���3"Ov!��@�f:H[�
Ю}ӆ�"O��V��j�Ҩ��� <lVЫR"O�5RI�8,C.�Z�P%���B�"O��H`�\6;mj��
 e��͡G"O��2� :ԼT�"!�3F�U�"O�\�C�36:�A��A�#��a�"ONxڠ�D�t����e��Ԃ 1"O�鲥��U�H��O��|5�B"O<8�"L�n��L$��#@�j�"OLq1&R�	��Q���H��,Ƞ"On�C�D�5Nҽ� _�x���� "O*q��ꊣ��U`�N n>}��"O@�C�iS�{��4�5���S�~���"O�eJs������-6f��I""O`pPd /5A���A�6X0�ѓ"O$��WF��}�Mw�[��h��"O(dȓ�O/BH����͸$�z���"Ot���=�شȜN �ڲ"OTA�CA�Fp.���P�8�"O���q��ad��!�pH���B"O�q�'NS�of��8�mY+Z)qD"O,y�$3�D��fo�PQ�"O�m���{����v�W���e
q"O.!�  �)�nɰsL� ^�b� "O ���� j��Br��L+�Cb"O��(%�*j����f·C�����"Od(y��T�����΍V�4s�"O��q�ʛ�S��bgl��D�($�v"Ov�̆�I�𱢡)�0�"O��S����e�8�Z�@@?� ���"O��02ʍ����aO�
 ɫ�"O0ǏS����YO�)�"O�0U�#e��Phd�ɋ3��0�"O��ڤ$H�aN83p�L� ���@�"O���&P�MN����ҵ]��� "O~�{��������t���"O4K7�Pjfޙ��Рp��t�"O�9��Z���p�m��j)S'"O�y�r���d0Z�">3�>���"Ou�r-E�t�J3�= 0�]ٔ"O��ے���&m��%�:n�Z:"O4�w���r\�����V��5"O�k"n��aEN5�&�0�˷"O����� |K�K5�B���3�"Ox���bN'd��(��M�;v��є"O� �4��
��a,��ˢ�	�t�`i�V"O��@��Jp���Y�皨7ø5K&"O>I�P� �`��#�-��D��"Ol�Ɔ@�3RE�WGw�����"O~���g�zh`8�#>DĪs"O���Ӄ �qS���)X:G`z�xw"O�����\���Ii�_L5�U"O�,����5r� �\���yD"O�=Y���0b~�A���z���l"O6�s����G�(0l�>W����"Ox�2�+����z5��O�b��B"O�l���lYS��$�ȕ P"O8�ٕ�T�<S�̇C����"O��!�_%e(�8*����w�4��`"O<lB��~��!iK�_��i�"Odl�` 	�<�$7�ݾ](���"ObL�� =>��Y"��]
�`pW"Ob��o�I���-���"O ��W,��A��v�G���(#�"O��b&�r�O@5w`ȅ2�"Ovlx�+�j�f�C.R0 Y�[t"OЈ���f���[sn�74$|
v"O�$��t��AcD��C2"OJI#�B9��YR"Eԉjm�� &"O,�D�@8�wB�H�P�"O��@g��xR��#����"O�02KVɲ��*���p"On$�� �#������"_F�Ta�"O��j��8� �cm��p(��"O��I��/XԴ(���N@X�"O (����ꪜ;���\|��2�"O���Vj$ERE�!
�aw⤡�"O���B6*�F�c2��`@Yw"O��P� 6 ޜ���ʛIFi�1"O܉r�gD�(n���lG�f��Iw"O�A��T���s̟
i@4("O9e�I�qd�m�Sk�0���#�"O�y�Ǒ1B��X0�_�0z��CR"O���C�>f�h�akW�,��|��"Od��D�Łz�ԱSӊW*1oN�c"OV,z����5A�"7�7wmi["OΔsB�%h���Ё/�90iR��"Oޥ�eL˦lET��$�]�!�2"O��P����fO�R�!^�'���9&"O�`�G'C9S��K�J�Z�0`��|r�)6�>����P pz���-�!s�B�$<(:�j�� E��}�%H�ttnB�9�T�"��)U����d�B䉪\ම���߷F�α}FC�ɦ/:�j�n��a��q�Y�rB�	�=	�h�#%�bp�D�>�B�	3lH,�pcLV�G�x�� �^� B��UVZ�$ܠMe�4���"�$C�	���A=�0}��E��3�(��WN1D���&�6 ����ᛛ@*@ě#�-D��� �ӷwZ�,��FVlzY ��'D�4X`�K�gҰ���Y�!��b�'D��
"��v��0"A�{̶���$D�0 �/�(ݶ|�a�A�8�Q�.!D�T�S����d�q-^�C
��z�.*D�x��t�~|*0�%��	��(D�ܡso;{��(��-]���{ˀK�<i�DP�S�Fyi6mM !8�zr�Jp�<��o��P��Xg@�T�� ��%o�<� �,���S%�P��퇭ct" �"O�Eg�I����94j�Th���R"O��� �&_HQ&*��`�8�"O��&��,���Y�K&(�"O��)A"�3��t׈�)C6����"O�8�% �z@����.y8���"O�l�%�ۼ �|���<~e�(��"O�p
��Fdm�a; E�`B��5"O(c.�8w�D�C�E�2Z�҄"OF��q��\�T1�	LB=	$"O�B4�R.�`H�qg)G���"Ode�pUaS
ѕ�{	׀�yR��5,k� �5 �yv��-��y2�Љ(�j�a��Y� w&��`'��y'���4TK�#֗�b�����y� �	"^�`�`;Al}���y�ƛYoȝ��CM�x"f���`���yrl��1a<@& �V�(�Q�y��~L�IWe��C��l޿�y��լh��}ہGޝ76��Ɨ�y�"�BsB]a%�'�X�qш��yb� � �6�p���REB�(A�I3�y���<�� $k�8;V;�	��y�V�9>�!s�'^6#��������yb'���^��7��)4��-���'�y�&��z��Ԙ�Q�6�yR%�<,d�Q&�N�h$n=����yBA�m��Ϗ��A�cL��y�/���!�w\,�i����y�����4R��S?u@}ǣD��y2�E�V7�8B �ǩ�hQ�C���y�,(��X#�"�@�4d�'�y"I
Q��3�g9{�![�yb$��i3'�*;� �w��*�y2̚�C�����`�!lֈ��b��y��%t^Z��ܖr�1���9�y�	�JPxs�#h�b9b���y��VAN��o�XF�\���4�y"�q7@t��Z&>�rCW���y���iv��Z�H�0����HҾ�yB A�6��A5�q���� ���y�*
m�)�BM΂5��6�y�F^�h����;\�x{�k���y�m�=i@��CB�\���j0���y��x��S4!�����i���yb�ǣ3��pӢhV3d|�jRl.�yˊ	 �5����`���F2�y�MO��}����'L��5��N��y��Y�o�})�A�2Hk��؅�y�X21�M�Ug��1*R�S����y����QB�	0T�B]������y�R/""NYꢧ}��AQ�<�yrOL=V�=R�cR~�*�!�#P,�yBI�@�0��A���l\��y����w������)7�,dʆ�R�y�G8d�z��'%]L���e�Z%�y�.L�2�VH���>C,AJ4��y���)Of�Q�Mg���IT�׮�y��@������� ��$"��+�yB�G���{f�ʶ0d��7�^9�y`L3Kс�i��(���v
�4�y˞�Ig�ɹ������e�,(�y�ឃevN��%�,���w�O�y���?()�!+�?7<YZ�딞�y
� �	�Ц�*��U �@�j,ʃ"O@�����|Q��8-��\bC"O<��`�33�2u@���3��*P"O�aH��1d���!	���ɨA"O~�(Ea".K�����?w7��7"O�$S�n 2I2X�֯A:76he"Oڙja�Q25��pö.�E)�t��"O �j��0�x83��N�����"Op��p��R���MvAxI��"O6���I���Y�G�&`2YU"O���J�+g��8�U��;j(Vm"G"Ot@p�MZ�h���"�!O 
2��"O
I2�ȕq�R�(bÉ�M6I��"O`XRs��'Z�:q��⋄az%��"Oz-hB�E%Ju�ݾl���B�"O�L� m[
Of8�&�@�6����P"O���@T�Cy�Pq6�+Op�� �"O�l�p�
�e[��'Ul�*W"O�\������EJY-.8#"ONtjq�;j�Tv��-H�` �"O*�A������@�'A�J�D"O}�U@G���D��G�U����f"Od�V Xg|D��`� 3�D�y�"Op,Q󩗿S���w�؞6��,q�"OM�.��f�̔���>�dܳU"O
(��[b@��BjQ��aJS"O��9��4C�I8!�S8z 9ˤ"Ox|�7��<mi0��TāI���2"O�Y�ǚ�\�y2̀e�8�Jt"O�0h$�Ҵ�A��>��m�'��N�<�#ؙ+#���G�#FLX
��M�<�e� 6�4u2�Ě&_�����^�<q%�R)S��L��"F 3��4�@nJ]�<A3J� V�K!�FP��K /�\�<����xA�1��$r��B��\�<�#-N8e�tp�B��&r�("&�l�<�S$2@26$3���Cp@�����e�<d��?��͐2厗;ߊ�j�NS\�<Q0��!ŀ��m��b��2�IC�<Y�.̿c����,��~TbP���D�<��A�u����Ϸ��{��}�<�sċ�-M�9sP(,\����5�r�<Y6�?_D��!f'Y"���a�k�<A5� cZZ`���)��'��e�<�c���4<���8L�N\A(�F�<�FsT-�ÂE7��u:R��V�<��g�5e|��+P�Z4a�4�hW��l�<��˳&� e;�*�����T��d�<�5�,a9VH+�.ٲ]�%�W�<Y@��4:EK�&F'* ��dIH�<9!����0x��ɥ>dt����A�<�3�U?��"C/�L�Z��Si�<��IȤ:�Q�f��XtX�c���{�<9� ͙!R>�U3�ư�KDu�<��FB�uî�C!Ǉ1RֶP���*T���LH�;|tJS���\z��p��+D��C(���Z�N��Xpѣ"�'D�L��
ǕoU4@��
�]M6!�q�&D�\hf��yD���1��<K����%T�\iቚ0(��9�fE� }`+�"O���U�*_Nf��0参IH�ۃ"O�!%O^=p�R��α{����"O޼���L㈈ӗc��.��8@"O���qh�7|���a۹0�@�1"O� \)%*/xٚ����q��� �"O�9	��ʾ�ΌX��F���}��"O �%̐eP-D$G*e��P��"O��	t�,4fT5�Ԩ�Pn"$3�"O����׊{�&C�޸D8��b"O�)Z�Ř
�zq��L�&"X%"�"O$H�����!{x<�f�25L�"�"O�UH�+����xۧ�B�4,,K"OlX�A�H.�)���a��D"O��TH�O(���%{���I"O
y'cU�K�*Q�q� ��2D�l��ْc?�]��QT� ��=D��0AL?�Tx��8B�V��;D��0(��Tsxc��>5�ͩ��8D����"����3��S$ZQ�*D���3-f����ׂ/}4�rd*D��z��s�1B�b+#����2D�T�PK�V�6|��T�^����R�:D�����Ū1�P!�8�Z0�E�<D�|;f�˴[\�Y���L;<!��.D�� BG�IQ�h�Ӊ��F�.�ِ�'D�bf��(X����k�P��E6�:D���T�X/z&\d�X7 �~͑�e9D��a������S@?i��(8D��%�I�TF����\�w���(d�9D�lcq�B�O�LU���*���H�h;D���$JyiJ���R�=�@�P�G9D�|�C��'vU^����+Jh|ъ�%D���0�$�6�:bHY:)�t���h&D�L0��ʏ^M0-�sI
)o�)8��(D���C�2������D�	�	�&D�hAqo��e��sDY٘(Z��$D�����ʆj��k_@M���F"D�xu	ދD���à�\ ��hH%D��1�D���8!���R.��*�7D��H�+��&^��0������r��8D�@�Ȃ%x�p�؇���4����+D�@P�DZ%K_���m�6)�� ���%D�haĜ���H�U
�=Q�@.#D��	5K_Kjh��S*X!8��\Jw�-D��jP B�hٞ��蘎D��0B*D�$*C�,|}����ؼ/��D"�f&D�,kR%�0/�E5IX�'}�,�S+ D��c�A�IN(��b�}�U�=D�(r�m�ZyR��T��q.P"H/D��z�@�?L�d��d���.L����
-D�XXE��`8F,�ֵ-�����!+D�Tv'�	�\0z���sj�"��'D���%�K�A��1y"�8c�X���	$D� ÇdH��0Ç��� |F��#D�XRB�
�9��L�刀<A"�RH D�S��T)aL��7�H1xZ�(�F"D�hc��8g�܌��ī0�2���o?D���0%�n|����~��ؑ��*D��`����*>�y��:�,��#D�dS"��bRl"�ߑO�~�`)!D��p戟�f��������bۢ b� D����e,-�%��l��Is0T҇J*D�P�o_�4��I�~EX��]�y�ʟ		9�Y#Ң�B�Y�׭ !�yr�%\d�����g�ԭ��JD��y��w����/�9X�VL!�X��y��ܧDB�ъ�� N�d!�L��yB-ӚVyPujO��<qD�Z��y
� �5�/Q6��Q�P]y�A�v"O�dr���X�B�A��@^��"O0x�F"�pXق�k���qc�"O�r'�H!+m��r�L��R"O��1��-$t��A�J8/V	q�"O���"�h��җ��* �a"O��Y��'��: ��;@�F"O��BQ�do ����	�b �B"O4]s�5:yr�d����Q"OFy��rC��P-���"OJ����7X�
���m�1p7`1B"O&8x�g��,��0b�L
�+=$��"OLؓ�&\�ZR!�J�r)���R"OA��6!�Z��CO�2#�d8�"O�xuV'%/D咴"��E��ۆ"Oh5��ǅ3c<�� ��		X���"Oh��EO�H�%I���6?z�x�"O��P���)�U!�(,4{'"O�%Qa�ަ5n ���ɉ	��6"OL�pf&�g�\��c�;��� "O��ٲʃ��w���B$��`�"O.͘�ㆪ, lbs,=;���"O�<����Q (F�\
7 � ó"O��[�I����tb'L�ZS"O��r��ί��HQ"@�9<�Q�"O"\	��)�V�i@.J�Lڒ��W"O�@Sa1![x	`�oչQ�T���"O��F�,�r��,
�~��b�"OҌ�Ы�mL] � W�[�4�ɳ"O2���Z�U���mvpZ��'"O^Ⱥ�D�)!�@l��:�""O%a5�O1�zȪI+�Mʔ"O\|��'%LrA�gH�yؐ���"O��#d���NB�lY�aW�E�6y�"OF�ࢦ��=�(�vA�r�(�[�"OdY��n57Ȑ�$���"O��X��'ED!�
�|�0"O�(K4` �!4�q�B��@L����"O��䅙�?,���!IPL���"O!;2���=*}Av�@�7��{"O����H�7P������Y��"O��h�ߝ3���1�ɝT��I:�"O�,�Q�_9j{�i#�I�'�~}��"O(��B�R"�~�`�#{�(5c�y"Oڴ(��y�݌�l����W��y��M�~]��teջ`p�U�À��y�N^%�P��W�V����E��y�HK�Y�M1"��9���ssbB��y¯R�Lwd%�7�@2]�T����yb�T*a]�x�3mE=y�t9J���y�ˌ%Uܺ��q��R]�P�V��y�-p�5�s��!Z�� @�N�yc��:m�U#�Ǚf��b�S&�y2H�[�^�4���WA~ɲ�� ��yB�ʷ�0�E�/g����D���y"-�
g<d��BI2[�ʽ(�ĝ�y��)��A2�A�V&,B!���yR�͙D|��3CL�4M"v`�1�ּ�yb��9��HQtD�%K�V0���ļ�y�e5�i�BmKG�z�6㝴�y"�ܺ>�� FBB �9��]%�yR���m{��r@)H�B��u��@��y�+]6��D�$m[�?���
H#�yR"��E���(a��)�y
� ��#`�-"�"�?3D�
"O��B%��"]k奅?0  �v"O��[2jߘ2E@�k$䗳@�Z�#"O����P�܉�$�e�d�A�"O��(�B؜t �@(��0,�R�s�"O
���`� �RxY�a�w�d=;�"OB��רߌh⸈wΒ�bg��D"O����%P�M��|W��xXX�H"O���B�*�beJc�8T�h)1�"O\i`���{{xp*��� �t�"O�Ѱ�n�!B�i�������K�"OV��J���,���,+�j�b�"OJ�C�M�l����F��u�T U"OBԁk�&�.<b	��"O�\%��
z<܁Z��B,A�����"Ov�Ǧ�B����_2L�tAq1"O´!D� z'�$��@٪P�"O`5�0��[O��33d��>��"OZ̊��D�ih(Z��p��<�"O`���L4K�"U�ǎ�n�U�"O����b�		=�$���+0(Г"O��QK�$��<���=N�� ��"O�L!�EGG��(��Ǘz� ���"O~);&E�02�D�
Ӡ1��`"OZ�b�OF�LƴA@䎕t5�1�u"OT�*�
�<��	�~$r��p"Oj���B�JI��l�q�P��B"O�a{mVo�r��FKB'��a"OX�ҁ	�2��$RFJJ�jC�#"O��{Am��J:�à+�9: �Xa"Ob ڴ���/�F��H͉sS��1�"O�h�fHU�
<e�+�X��"O�!B�DP�J�谨Q��-4n���"O�C��0����3��,$c|ճ�"O�T�%ڢc�J	x�hфd�L;a"O�x��A4)s�����
���	�"ODt�A�wV� ��m��S�|ҳ"O�y3E#ާ)R0��^5�s�"O�I!wjM�>+�eArL�		K��Ȅ"OP��@���N���e�ȲzBN��"OD�� ��G�x`Y�ˑ1&��DB"O�9�E��x�Ĩv\/ta��ۤ"O|붢�c�ҩA�[C�D"�"O>��%Ǽ��P�p��On��4"O��R��0pe��qV�Mu��pp�"Ov�Y��-|��8�F���&I�B"OD�ۢ�N�%�XP�F ) ��["O�(��I�{:LZ�fبO���9"O����5��xqń�/:�����"O���'��I:d ��Ko���S"O�dC�E�A6*�#��΂��"Oj���#�t���o��j��谗"O@�է�/�m����
(��lH�"O�Q�
_!`���	sa�
��,�C"O�(Hw/�D#@<pfb_/H0��b"O
����=RKHH��/+�5��"O(	�b�@"� �Ɇ@B�!��c"O^���Ȃ�?���o�	h2�r"O�A*F��-M��Dk�4'�l��"O�q���e�V��0�ݚ�H$K�"O$�����}0�]q�*����"O\�`��Ril�Si\8�$��A"Ot	���[1OJ���6H s�>(�q"O�ј��C�V�(MSŦ9[�����"O� V!)e`��ap�! fJ�f�V���"Oډ�� J�#�r�z󤑚:����"O@Љ��B����@�-#x�c�"O@��b��2ZѲ�ȣ�	6m�%#�"O�0���)i����KWE���R�"O�1��W�ɂ��*��l��"O���W_���!�i�����"OD��gd��K�����)��� �"O����'��GF��Z�����y�"O�Ě�ϐ@p⑻&�<A��1#�"O U�OT7������]<���"O��I��T�8"���e�A�)QX# "OQ!E�ԨD�3�N�Eh��"O�0�����:��p5,�6ⅲr"O�,[&Ǒ!�P�ժ@?^>J�p"O�����G8�2I�e��0,�D�v"O\4�d��lJ �C	�Dxa�"O�4�p�í�	�g��-���"OBT�2��Y3��HU��E�*h�"O�JƠ�H�hP�t���^ �e��"O�m��c�|O��IB֛��pp�"O�䈢��>�( �BW�C��PӤ"OB��c�սe����|2�5�E"O�I���r�R`��'[�]2.,[�"Ope��gZ�u6�3��z0U��"O�c�a�@�:2e�^&N�S�"OP�)�*��E{�%�E͔s��� "O�r&Kdǌ��B����"O�hh��,{=���t��P�$�U"O���E# �>������}����v"O2���n�&? ,p�`��P� 4��"O��;d�X�o���D��Q"OT��@F>G�2����]�ll�5"Ox��l/��@���<�x-R�"O,Q��ZLڡZfD�H���0@"OT`��>Z����E) "~���;p"O^�2!�؃�@MR�%Щ�$��	�'`B�*r��]��C([����'*ƅq�&A�/6(�I�j��rU!�'�T)�P��K�n�r����.X�'D̝��h"70(۴cԶS"=��'��|�e��f~��)����R�>	)�'���eK�0#PY�׋�)~�ڄ��'���K��M(�I��G
H{`ě�'
.���*iHq�@j�;D!��'�̳E��gʂt��	�!�&��
�'�>��eB�a��y�!�d��Y
�'f2dB#O�q���9D�G4%�4�
�'J�@  �i>�k�Z-K�H�	�'������=?�n�󆀘K�D�K
�'ӆL'�e�r ��l�ID<�	I�TE{�����lY�3��<�r �p�A��y"�Yf�X�ZR �'����K��y���G����R��4�<���F^��y"D��sX�Y���-�+gWV�6B�I��Y��-!E�0aF'"b��Q����0��e^�t�ڰ�@-L�#*�"O@�H�A�#]��(�5GX�gq|415]�hG{�K:�0�trEÞ"�p�9gkS�J�Pцȓhܙ�w��_]��Q�g	0?K�0��ڰ?)����|&4��Ć�/G�y($�G�<Q�eA�IzA�%�'�Ĺ�4�A@?���c5dH�e���O(��*Ϊ@�ε��5e�����V]
�hu⁑5��S�? �qB7g
(�T|6"��>!bl��"O�RU�%�Ra��A6H't��"O� w,�&�i�`����"O�q�)�#o=4Y�����=���3w"O�(���߹^�,��Y,a<�{E"OH+"*v�Z`�B�βq�*�@��'&ў� #b]<:����J16�	��3D����GF/"	�J�}m,�p�-'D�8�!��e�¨��G ��;�E/D�t1���9��ͩ�KEl�|L��#,D�k��ڗZS���/�r8�g�+���ɷ~2���!ߦ` �1��a��˓�0?�*Y�c�z!��5[$2Vd�t�<�E��]HL� aL'8T"��g*BL�<Qń� `��ʁ#��4Ĳ���L�<A6��c���,�2	�kT.:�ԅȓ���a�DFe�D��.�*lY&x�ȓ^�����_E�n�� +/"�ȓz����̓.�F�3&,5�zԄȓ]U
}q��_�x� �è���� L�)kA�1�$"��
/����ȓh+����6Q߈����R`o~��ȓ�.��r,F�S�-�Y,4T�����?�&�x��]x��H(9�P��'Ox�<i�`ǀ#�N9�w�O�,��ps�GP�<yd�B:C�0�K᧓<� �@�%�v�<i6�S� �K�(�T��f�i�<��Z<7�`�2jP4CQ �R ��a�<ɷ	ނZF�8GHE�4DP:��R�<y��Ù�#���/6�
Ub�v��t�'pVq�ADǩ�<��u�=8<R�K��G{�����$QZ�[s���*�I�2�� �y�eC�R��dPT�W�",��nH���'�ў��<%c n"P��`j��R�V� pF2O�=E��B s�0�g扺o��uصM޺�y���$�=kvD�
e&|A8�O��#ў"~Γ+�lhS%��`�<�b ⌠?Iޑ����QQ���w%Dr��%N��܆��S�'�l��я�IQh,�S�T&=k��a�'����5Q
�t�֍��8�Z�'6Q�#��	��5�5��+u�\��'�iò�5"؍�Gϕ�p	�؀�'��Mp�*ʲ3�)IV�K�u��Q(�'� ��cGȓi���:ƥ�:r���	�'�h���N�Dנ}{�L@�yeJ��	�'��p//���$�rh�Q��'1��!�i�7q�C�`Ψp����'AD��ԉ0/�>X $�P�c�5��'|�<����4.�4��˯b�TS�'�dA�Ё�ޱ3��̯S�L��'�f|	�ĝ�G��� �ݟM����'ږ���g]
j�,A���H����'T�[���+4�֜
����;b�|r�'͔��C�T�zH&y��j�/9H��ȓc6̑�T �:x�Tᨀ+�5� ��bV��q˜�D���Am��a�Ն�Y��!��@�������D���E���QD	;g��:r�	Qd p�ȓQ�6 �K-eͼ��X�-�Ѕ��x$��	a� �@�����K�n�݄���A2)?D���K��-��������H�,�XlC�C�/Q�}��a|L�3l�+N^�1`%�M��Yj��޷|���;��H-�u��IU�)� ����͍�
��7�WBv�(�"O��3���XZU��TI��E@*����ތ�c$���S��&R��GO�D_!d}ʠ�V#�~�����Lݜ%!�dS����֣����Q8�!�,����%��ot��rI��T�!�D �N(�
�JF�x�h��e�	���	��hO�4��u��	�jt21a�h�*01"O� pƈX�0�M�������"O|Ur"L��'��٧��s�����"O���F �A�l�.^�)Z��Q"O�$�ҠD�Ix�ǚ�j�*xQ2"Orl��٦V�8��7��v��0�v"O���`/�,<�<,��	+J-����MOe���O�Z��'�&E����|R2�ɐ����'��ْf�b�����J�L�f01��$=���!�/��h\	9u��M�܈;�"O���F
�>�Z� �ֽt�,�a$��l��2d��qs<����X:�ZeD*D�� ���l����H�%^Q;��)D�{��٪|$�\#��{��<p�*������/I�@)!��-f��Y��э�ȓ9�]�p �=\J�T2#�J^����2iF��%[88�����o�$���p�*%�L�j���t/V8e��oZS��������F��a#� �l�Іo�
�y����+��9�Ed�}���Ba		�?!1�'��y�0K�>�t	@�*ޭ2��b�X�O>0�!���ukh���j��oW�4�"O�8B�KTl�kG
Y=D9�Thb"O0��BБd}H���c�H8T"O}A4
Д)شZ�h��B��xC"Ot$qɛ�u�jL�*�k�j���"OZ����S�bT����a��R�"O���l<�4�Ǌ�30U�pã"O��Ñ��F�^dK��	f<��y�"O�j ��=��)q��	O%N�cQ"OLQ��1"���S��(5`�b"O �&�\�զ�� ��#-J�)""O&���$W$&rd����4K&���w"O����Fl�0�����M#ZL��"O4��5��� pE�G&��U"O�B��C!��p� �,F��"O�- ��1Z8��y�.���Rv"Oz�)���?�`,���씩)�"O꜠񫑩͆	(�o��t���"O���B�qCRIi�)S�;�0�(�"O�����)l�ڄ�犌l��U�q"O2��b��4Ș��dW��;�"Ojq9���:im*9"#��:zJX5�B"O@AP���W���X�V	W�Z �"O.�Af��(���KN�l�T��"O^sCd^�Pt �++y ����"O���0fCG-�L��*�9v�:䙁"O(is�b�tn��oSdӺ[�"Ot`�M �&�(M��mI$�i�"O�5�t�D^,z�	����@9ݓF"OB�S�鏃'� �p��R<X.J��D"O�`3!M�w�U�C��sK�T��"O<�(U��7b� ,C"�?kEfm�t"OV�xrH�	.�P�+�#V�6��"O���pAԗo���X��	O5X!��_E}�0�ă !��Xc��A(N!򤈰`�R@J 85԰XbG��$e!�� ��Cs!P/�.�N�Mc�=("O���hÚ+�n�:�cD'k]�۳"O���BƁ�h"�� M�����"OҌ8p��`�A"�l�4��0i7"O(e�S��71(v�zƫ�[�ɻ�'4j��d.H��a��Ɋe�����
-�"f)��N�Έ{�'�bԀd�U1"�$PFKA JnP���'kz���燰m��M ���~tʽ�'��0��Ėy�jb�˿n: \�
�'u�C�,�&@,#o,n\P�j
�'c& `�]<[ǘ�����a���Q�'O�ѓCb
	�2�*��\2� 
�'^\-�'d�;v胦C�&��H
�'E�Q�OB#,�h�"7F�m�	�'��Ԩ��8�PbMBkL{	�'.8�rr%��o�f!��G%%��0B�'���d
�{~D+3(ѹ+3 41�'%(��@NZ�*Y�qx�-~:~�k�'��A��@b��Ӓ)ޓq7@��'��)�(� W��y�.����'����&���1�����B�0z|���'��xn��@��z&�	�i���
�'�D�h'K�^�DM�%d�o��� 
�'l(���,d��Sg��$��'&�� �: ^�S�(X���L�
�'FH�Ƥ΄(n.���
�<�6#
�'�*yr�_���!9�L7c�a	�'ʤ52Q`�E9����1y�:	�'�9k$E�#U� q LT�6�����'�d���+̅����4��-t����'�.�at@V ^�t@ZQ헱^�i{�'HA���\
Ug:� �ړ@t���'�4@2`���S}�|�Ľk�"x��'"��GHՏ9x�{��� ^� �
�'�ڜ��N��#=^��F�̲^>D��'��T�.K�p����6� g����'t���6�~�R��D�A&auv�p
�'���� ���d�Zq�F��_;�X�	�'B����k�����EA.PN���	�'���J	�f�s���MFu"O@Ujԩ�26��r�,�$V�^��"O�h��>H��#͓�e{��yp"O |���F�q�@r��՘Z�P�PR"Or���
P'b^)C6�G��0�"O���f�n�w˄�\���j#"Oj]�b&��k�fi�b`�� ��	2�"O��j��\�k�5v�%J��Ӱ"Ot�ѡ�� y*����3gf�9�s"O������9t�|�B�H�4VQv�S"O8�qQn�#,���FN[X��(�"O�[�@ARb�a��eʰ"P�,(C"O��Ҕ�@�$̞�k&i�E0�� �"O�a7,�2k2� (N�(<j��q�I9�f���Dc��򄝏"L������9z�HA!d!�����	�OOpF��@%��|�(,�@j��4p@�ԘVazB!U��"a��C�� >�U�F�B���<���Н8�M�&ASXEA@$� �
t1b� ��\Sv��F��dO�J���K0��*z}����3��'�R�ʀj`��1'�֐v�������ʝh�U�d�xXXԃ�i��yҡ�_���	�ؔg���x�K����[���A���d���XadK��O�f�'P���P��g���(Bd�V,��'�ftW�.�PDؗD�-�΀it �s-�l��k�xB򝃂��D��$C;lPRsM;�Pt�UD�H�xb�M�jQ�P+���D�u��f� �"��%�J�h� C�=�[fO �� 0��FP4`q��!uv�Ջr�>!�邿6�����ׅP�<Җ�N>!�q�6��a��B�a2Q���:@��"O��w�Y������`�~�pɉ4 �v��p-�z��g��Mq�\�Of���Q�Z���� Yd(ܙ�t
O��1Q9�ޘaU�UJ�z!ᯅ%g$i��O̚PXDY�D���RTb� k, ��ɶ[��Y���-��ɯ&�`�296�4����¨kTi����3A�S	D�k��̻D�R���U�5�� ڑJ�$#G6��AΜ ��IE�t�C�ݻE��G&��A2\U�d��ħY-( WjH�b�@ ��7�:1�ȓ0؁��c�3V���Q�.z�h�pc]�\6� �nޜ ���MY���m��'�D�� ��ROF�YNF�b)(��'RJ�D!L�Z;�u¦�H蕡WMh	����3d~�	����Tb��I;���F��8W,�h[���iX���$\�^��	�횷+M�y��׍w~����O7E��q ���/�d�0��N=H���ğ�Cq�o@�K���	��0�qO�I�tI�W�>!�'�z�y�@�M���'j~ʬ��K�?=Bi���P�[�̄�{�\�B��>�zh��i�Z��笔�,�u�HF�.�4����y�^c?e�3�rj��7[�*� T�8�	��Ω�yb ��F�J=��R�E�]�%S��bD�U�'e0i ��Z��Dce@��E�XFy"�� pR;Hԙ0�B�s��p=5�"T�� ���uY�<�����D�@hwG�	��\���0�T���tu�|"!��"�� �[ � �c�
��'R���!ĝV�h�!��&�����8P���4���A�/!Hy�AG�Ff�B�	,x ���q`�9i�,)���_��ʷ MH�`f��H8!��-z��XlY�wC���fC� q��@�ND�6�V#�']b��U�ݠS�Q�
3��0�>\D�-*���3�Z4Y�H�]f��%���O�� �ʅ�Q�,��7P�)u�'+�Y�F��{�T��3�ͨa�~���b7{9��o�	 �a�	�,m'DP�ѧQ��y¯Qg�b��=�OA@ �	�i��E*�D����{2q�hC�"�L�`|�7��"�0`'M�5!"�U�_ڈ$`g���X��Z?r`\���툂wt�O¢}�!?"�t�#��ɉ�e5)�x0��B�B���	b��oU�d��OV�%7,�3D,+�ɗ��˅�ޚ]@���t`ӟ%ᦴ�1f�O��E�O�L<�A2N*\O(�	T
[�̼ 5%��}��mAD�P��Ŭ��PW����v���iT�Y��� eE�)w�%Q7@�C�����V8ga�� !��qq�����'�Z���%߄?�BE�d@����[�o�:�( 2&a�5(	�tR�h�2c���qi¡`�x��L���!#�'�(��L��Xr!jk��F-DV܁Cb�I�$��D����w-p,&b��CYƭJ
�y��1r�O�^�j�xX9JGcڜ'�*鸄	ū3���D�v1���~�'@t5R��O�>��U��$��!��'��hu	-/=��'��&���hN�Q���>U*�*G�t4e�FԑZ��4)�"%#�~� 7!R�i�R=��+	Sx����N>���x�iV�6��H���Wu�p�#n�R�`�qC��p�'�:�:��"� Q�ϝsz�f�X�R bGҝ<jf)@�'�0��k�<f|d1�
K�C��ԇ�=��#f�7���AD�Lq��P��dzf=XcJ
�D���D�K	9�կ�\|b�#��$���iO?�E;���sN8����:Jv$ă��8���9�*�r���Z��Ȝ4�ؑ�@A���HK�l�) ���Y�i]98z���7r���B�oȝ6�Н�'ִ�pcQ�d�P�׫{�*��'ZޘZT�ǘ3�H�3�	M�l�h��aL*B�b�a��<G���ƭǊ#3�T�/�8�
�3aG6����ɔ[�V�ü�I�AF�������s�T���Z�y�|1%�R�>B-I���{��-�pgU�<��DАp�Z��wj �*5�r�q����[Uдs�A�p=����+g���%����0>�ŀ�-f�5�l�*T��5�R2v3R1#��ǐ4ǒ�rE���Su&+���0`b,	[w�T�r�"��O���Ul @�s����4��bK1pR�$	� ��O<Xz����~/�({'�ĲH��0�@g�'1N^嘳晤8�ѱv�[�9��10 T>d�i���k�Q��*ނ GP���FY�<� ������<��I!=��j2A�	bc��IUo�p�
��ѫ'؅h��S�Ȍq�I��:� ��!܋ae��y%O̙v� �s��hU ٛ"$΁d�E ���0O'Z��%�?-I�( � ����(�"�@�'��1X���M���Iw@��f�#�� b_T��Ϙ�d	�'���<	0��06���O���G�A���'�t��ej�-#z,x�:	�nYԭr�i���������/���wd���B�G�ݎ�ʢ-l��Q��+g|L�1��rЋ�lY�'jX�UjVP{��$#��k��U	�d�1�&�>�Jc��Q���Q��h@��@Pf:X�'McA�$S�)	bJ����:�����'�+�!Z��шS~��:��J2E\��E���4iUgY( � �[kT�h2��)abi����SV,x�ՆՊ"
��؂Fץ~�e@�EC�\dJ�� ڋ/lx]�w.�VY�ɗF��Ě�
�%��H2�Dg®X1��/._��"B�L�D�Z$)�
A�Q�<��,�r:N�s�ʄc���i�Jt���R�N(s�4A�0���0�^���!qC9D��T�N�g��I���H�#�jIp�bc�;��,A�ˊ�O`(�2�	�Te~� ��#%`@fOڲ�8<��ǵS�.^ f�=kٴ?��6�c���;��?7o�li�ʝ?��}s�'9��M�aA�IF�DA�Hz�ɈHC�d����"v|�;1�'�����sN��B�� �|R���59<� y�M$[ɸ�m�&V)�U��c�>�"�kb$��۞~���0F�)�v���2�rԭʺBt�@�O%� s�J��Aд�S�gK�st�0)���15� 
$�i��6��8N��+��{U�DV��ufӦ{ ȝ)2��1UB.|�1���\l Y��"&��C����#ڼ� 6�TDB���J�#�kZzo�E@���
� ���D���BhI8e�B�����<yuNS�c�P ��=0���c��"Q�&		�M5�HP�3pw�,+\c��8�AfL.2�D��C�gF3�db��c���<,.�f���w@���n�
e�P)P�M�4e�P��,���vY�u�� ~{Z�&���+�<��0eFM�M���`��,���{�Re�L��I�2�q̝FJ�c��N2J0���
3���'�d4�ɕ�e;��+�a�+yk��Y�'72�jEe�%q��0Eo�9� DaŃ�,Q[�ej�]�P��\����W<$�2�%��u��-H��nAe�U:$�R���`qU@�Qq\]���dT RTV���O?vg�Z�鉂��%8��Zu"�U@ Νxi���5f��۪%`G��`���7���Z��o��S1�C�}��c#�T�7��薀��)b� ��|<@��E�4l�⠖N�'�|�P�N���pB�ټ��G	A�(:
�����?1� ���
O&(���S`�,;��K�.�=>��tP�*<�Ŋ�<O��cj�49��:v&�'.�ek`�޽.'��N_�5�F�[>|RP����� U�ܸ]"m	�ɋ�%<jw>%��l�*h�cɟ�xx���2JY��Fl�&>����J�O�牎h�8L��/�
�v`!���� �W�U�NI�57��8j�^���$ֱy�@�$D�tk���
��xDp1�mUOM�)(Gf��k�^��d׳}�V1WÇ�hI�t窋3Z((@ �@S2r7��H6r���ubC�:=W�	'f�d�(�,F�X�فQَ�$���Ϟ7�v��P�٨j�)`���I��\����.��*���2�j,�+N�]�Re(H]qJiR����6����o5�X���9(=���$��0jl��U[�~��g�tZPU:d�4�E�.(|p�YߴK�����F7i��A����<��'l,h��4�|��#S��9��Z�f�'fD�{wlO+l�@p�]ܼ����F�3���p��g�-0���唊,@�����Q{v�"SlX3.\T����m9�$-1�2�
,A�S�T!Q�^���$E��^[  2�a� ������NT���e��c�Sk̓�@%Bt	T�I��m
ń�#��It�ܹD��$UA��YR�O[��y�&ǤS���{u(��EK��i�&R��$� c?Q�8�8d��j&!��Ґgr��ת��F��+�f�3.u@`�ǁ�=ξ,0�� l�<�Gd�
bW���$�qQ��z>���ֲ"=*���F�v���F{��LmfM�e,�����O?RFMH8a؉u敻��È�<i�TT��C҆N!��A��?g�T��u�-M�- �䉹@�>�dUY����� 7B����3�'U0�iK0��c��3�/�H^XštCY7Ep=+�'�t\��e��ɘϘ'<�UB��ZHb���T(�Q�#�<a!�E�= Ձ�����%6��Z `	'.�b�̰Fd�@P�oA��X��]8���C��?�,Y"�O��*ggG�37씊W�&��hЉ�$X�S����2fFS���&8_�Q���29 1S�@S!��>��@VJ@��c�s�t�|�Ke�Z!c6����+uꌒO4���K+t�lD���0��<i%�5��|P�΄�����`���z�)ҧ5�2��œ�S�03,޾hЦL�ȓUs�up� Ǔ6A"�@�gȒ�X,'��H�'H��Z��;$�.P����)^�qHS#w�!�B�tV�P��&�M��P�nUX�!��Y�+���b���a�R��c�L�!��"xs��t���$P@��LY!�D�>@�L��G;Z�����V(eD!�ԧXblP ��g���u�+Xd!򄑲z^�x����(���MsW!�D�Bz�� Ѫ�h�qk�@�JD!���d)h��i��U�d��J!�QBO�p��':�����A$�!�9t1�i�.����Oq!��:656٠����:Jx��CI�J�!�N�x=�y�� t9Z�eA;�!򄇤N]q�A�[� 6�y� J�E�!��ì�� �J�L(La!Vş1!�ďD�R���I}�8U`��H:Z�!��6G������f[8p�1���!�$Ѭy�����a��A6��J��T�!��.69�z�U�����U��!��v}��r�� e&|�P�F6!�$�+^�.Ty��A�!X�Ed C�m<!�ċ�I�&�k��� ��J.ߞE!��F1����`�|Ҙ�s6 �!�Ğ�(�zi#F�SȪY�䋁�!�DG-D�BT�b��T�d`)GF�3!��A~ᔜڤ��5U�r%���z!�� Ġr%H[�b�DAQ���8w�dB"O$Q �A�.h�q��^���"O�@�QO��[��4`�A	�u�"O\�qCJ�8	���U��6bm�E"OZ���ʷ�TD�R`�a|0�"O>��&N_�,�q�T	܅G�(���"O�1aB�u�(�KB�TT(���"O,����K�x.山	B�@k�!"a"O��@��'Z���#�� ���XQ"O`����_���ꧤ]#F��}��"O(��93������,v�`�j`"O>؋��T4��	d��Bp"Oθ��(�gWV�[�Z`�,�B"Oi��g <����6*���A'"O�)���˞m��տnp���"O����xm��gX�o����"O��R��
)S9k�D�9O�4��"OL���;&\��D"�.j!�0�6"O�Xh��y�VZ4^���AȂ"O���'#��wrD��^��:U�s"OR�9!)Rr�Y���w�\��"O�!P�^B�ᢃ��@��	B"O�C��ؖe��G���� �G"O,��g�n�pÂ�h����F"O��X:>�(�P����m�"O�}I�R18Ê�dK�w��LY6"O�,J�طF`�!v�Ɔ"rP�q"O��2�cނ3�=����'p���"O���� u�p�Vs^�h&"O��'��^t�S���<�e0�"O�H����3�^]�u��h`$1�"Oq�J�$��Jƅ� W`XYe"O21��ɞ(�f݉P�
)N���"O����JO�>Wʐ"�H۪ �N��B"O��,V
�8]:�GL�<	J�jo5D����lH�4zp��Vg��RhXȑH=D������3{�!V�Z�d�2�	;D��#��J�,��YF��J�>��p$5D�hja��H.��r���0��)D��cשLI�Ȩ$�<�FxX�+D�����@�u�f��t��>z�.�YA/+D�� +V�$HJ�:ՏӾe�V��u�&D�d��A���O�lez	r��&D��i�iJ�$����'̐B�P]j�$D���%��4Z�9�.�?���"D�H�ow
�3��^�1y0H&D���1�&�<��#�V�v%Z�B$D���sb��cSV͐¥�<);S�'T��Q��跫�!��ܒ����yr�C���5���!'v��`����y2eīQ�ZA�� U6�`\"Āҵ�y��0 ��Q!G��|q�1�ybɉ=*�NQi0/^s�l"�Ǻ�y� R�9�]��d�Z-�x˰䋙�y2+�;]���e/˜Z_��8 �A��y�c�3v�" @`�؏K��\�G�ϼ�y��� ^�)�L���0`���j�� ���Fe�'���D�,O-��ې ���0�����P�"O�H N�sk�y³�2��C N��1�F�&>��9��')l�0�F^	.��Q��.O���/��E8�//L���b��R��#�'�/5��ɫsB�>�Q�O��F�7�&q`��FM���x�f ��t��C����#$��O��p��55���Æ�3A����'�@ձ���3�ȭ�/��W��L�-�O��r�;#�f�Y�J�6ʸO0�ҧ� R��X���@U	�W5��
'
O����qFl��@��)I��9(f�C
Q�8UIפ׎_���o�a�8���e+,h`0�T$&���crL�d&������P����V/��[刭P�'����z �ۮ����c �]�C��l(<�6L@- Ba�p��IWT�9�\m��#�������;]ј5re�oƙ�}�ue�bJt�;�)^4���Ho�<٣([���(k�DH�O�ʀ�o!:��9���M1`C�X�$n��9� $�}2�>)W�ܬ)n\T��A�Q"d�� �`(<9��'#F�ŋ@�#�D���~D�`z�?�"eXb����0��w�+O>��ĥW�DٜQpe��I�l]0�'�qKƁT2o0�륡+	h(m�p�Ɍ"���3���1=��ВЮ
���8
�X`���5��(o��9�B�G.p	�OIS�e�X� X����U��]!���5e\����:��5 ������ҧ����"OHq��HQ@�SOH��lP�hD�4�ʵ�䥅4��@�4
�6���$��ҡ��L8 K�{��P�w�N1v�
��f�54�h	ul@�{�I�bfڽ鰯֤S�
���6~-�l����zQ5��`�'������=|%ço@:%� ��?����G � f�IJǏ�L0��b*ZT@%��N��H���c�-%��-��7Ԣ�:b�s���ц�1Nr��=asc�#3x�����h���׈52��`���5��@��D�:�bErmZh��"O �V-��Dd�J��
E$8PF!@mو�0�Ǝ*s���d�d,������ļ��)K(F@�b���#45��k�<I��[�Q�,�*�`9[,j��0��!Ǥ�Պ�-ex��5BG	���I�L�;R�:�<Q�4.����ţ;t(�0�GQP�����O<R�)�\�K�i7 ��f�Y���&�E3�C�p��"����p>AD�N�l�H�!�-�6m������OܓT�r�CFơex�XӴj�i>�]�׎>m�)O)SI����Cś9�p��ʝ;f�!�d<.,-��휵5�L�Q2�֣��4�3"���e#�)��"|rBa���O�Bϻm*��
����=*��V��ȓg��@���0+
r�i��y�~6
��$Dl4�r��P���7
F�g��x��s�'���kCK����g�(vH�?�����\9k"�͋�L?ah�����?Mh��L��gvj�kvv�C��>Nn�N���sM��g~di���,�x�0r���h��08�DUn_b P#��!c�y������#g��A�n(I aIB�8P�FON�<��&Z�!%��'�V���G�'Yk�=�uOۣS;�] ��^rhY�UƝX󸓟pu�;<{������0Q�m�C��'?FA�ȓ����tC 2f�x"��8�1��iۏI9$�1�^ $[�T�ӯ��?��4�3`��<����T>�ݳЪńtV���n�y���R�ּw���
D�myn�ٖ�H�Q8&�#͚2n���fWjT��@���?֪!��I"}�0�s����Ŏ�<$�\�{��I=G�����߉ ����`�#�F�3��Q�_������'0�� �b���[���}H<y�L�f�}��
���A��g�{?9�M�;\���䯓?;�	��7޲��C��I�v�Uk�9���#)�/ ��	-��3pB�$��<�RM&p9YC��jD1ja���7�4	��bV@;B�� �!_�ɦ�b�6m*C'���ef]$����l�:��ŲE#��!�+;�O���m��;���C#m�Q��e�'���{�� ��>1ݜ�ieL]}yy���ϑ:���+�MI�U��Q؟'���[w���)�@�?@[p�҄�R�\m��ɑf���K�㲩�JI�81p$;Ht�����!H�Q���M4���K��@	R����46퉃$u���iј+F&�*���h�뎍~%2mh2��;(�9��⥟�3ѩ��E<���oH� ����g��$()C^���XP��)\rИ:gM�0�X��!��,�����M�r�lp�������آ?���_�z�ʹ+���@ԃQ��?��i��I]8%ETI�0���-D��*�$y�ĥ�dTZ؋Yw����I�D��(
��A���D&2-8'���a|��A�BfUp��ǉ~��ш�k\�'��)�fK4 h�Ї雌K��98�͐j�pC���q��,u�l�A�.�H����'g�h[Rn�4f]��:FL�^�Q�([��4 ��t&�Y,d��M�5N�1!lԁ4-�%ht
p
 n�V��L��ܫGܬy�6 ���(e�5k�Ɲ*t�ۤk|\R�N�S���~����41֘�a�c� ���!i3(Q+��ș6�5��Ѳy��$��S�5є�Q��آ�%���H#aT���E�e��$�e@Y�xYbyJ���:^-:�0�i��_	����喦��Of�!�P*`��ĳ`b�60]�8��G�:Pd��/7�>�(W��'ƾ$�q7O��R�/Ês��ӋPvXA�J�>~nM�B̹6� �8��F����
0���p#��[q���Զv?��"�P�ta����&X3@}{�'�[�K�K��H���^�6S�p0h.���%A�:	��Yw��fU�����@�>��b�������PO�ia���(.��l	1� !"�yC�%�:4D�v�͏g �6^6�cS�AkK��P����'�]�B�3x�������eƵ rl���X�H����S	D�NXh|C��dƔ)�4
<�V���6v�`LYM���ѫO�p���ݦQ�)����B��2oϥN��Qb��_x����D��%��L���� �0�����h��HѯZ���ˆ. �*���`���튕�˽n�
�l�^7D��\�u��ݟʡ���J�g��A �ၐ*�P�BC�8Y��k���Z>
�<X���Ser�s���?>�qB�&!]��x��#Ֆ:,j���&�M3䋓mrx��E,}x$�s�<��֧�)*zF�7'�d��U�b�d��p�l�$z�&�t�Q��&l���	.(�9f����tZ @�)c����1"�����UW*��eWL4"��<2���+)�D��g��!��)-��"���`��١oz`Щ�S=#<'$�4v�)�V��=o �K 3tJ]{w "�M˃�i����'��@fH�O���V�B1��ݨ +a�Ru��![�n�>|H�K��%)��G�'�\!�@�� &A@�CW�n�^�h�)���mZ$	�p�J��+ʛ6�u
�Д!܌X"�Q"%#Y�<��B�3�%�%fAl��N� l�u12F��(����(��cp�C4LL3.eD�E�Y��5���0kl�,�"��Y��P��/���d,�v�0(fF�'f�x�mLcW���U
��wo�,Z�B\�2oXQ�$'�dE�,cД�ɉ�T=0G�LA�@��Z~@e�Ąƌ_�X�d�7t  ب� �|	*ѩ�÷I��]������n�2!�v����ت"�$9q���*(����R�U�J1��`.Ԁp�)�4��J�2/0�)��#�)���S�T� R)ؘ*�\�C�ڀS�AX�n�zE�GQ�/FJ�`նu�����B��<�mPi�'�L��So�H�XWB��iB���)�8���d��v"T�V��E�$���H�K���UoI���	ӈ>��YN
>,�Z!��<l' ����C���S�2ғ�l��A�_5E��nޙ���T�w$J�Z��� ��)ɪb^��"E+3P��` �O����ᦕr,Z�:�
�D(iH�˓�(���H���1�@9'?i�,E8/t�����vtH�`Ձ���^�C ��:���0$�)�!�.�:ekn�!�
��#D����S��~���@*�yr[/*�(A#�N֣����'J6̹%����)A�',/p[R�\�`�Θ|�m�RBF2!N>ܙe����5q�g^', l4҄C�Y�����lW)"�x,�eE�$�&���Z�<1�N�{[L83B	�b���GxR��5r��ca�\�3J��&����&��-|�L�HGM{��}JU�Z8h�6���.D�v���W�&VS���vO��y�PШ1�Ҽ$j%I��Y�F�#Ĭ�H:�{�6�{K,�"F�:�����X&?�l��ľ4P��jĤmBz���do�D�kӁE;�@@��4_ؚ�-~`$�0�
M܈��'�z���5��X�aS�$2��RC�X ��M�'w�Ј�+L>d6��M3|�h�dg)��N�ee��4�R��\Ft��QR�Px���2H�U!d�l E�A6�B�5�p�ɯG�`� �i�nq�@@�"���"T�F
 �p=�VG΅$x�xI~��yrLH��U2d8O�R-*k�3�?O"�Ä�̣'�������|�<90��?t�摨�
��j�4�-֦m�~�d�_
,�j��F�S�3�`iF|�mT.6���3q�U'z� ��c�2#Rx�쎂gBY�� =�OB��ǉ:`M���Nٟ:Ȁ��;,�i�t�L�ttL�瘴b���=���KhQ,�@S�F�U�쥟��ӑ ��P{�9�t�΄}��T��	��?�]�Jאf�|(����̃`�0�H�Ǉ�<ʀ���]8Rl�'uh��lْ��]8�?37�ܢ�Li!$�O�:�Fq(t!Ƌp4�1 ��<�C�Al��|�<�ǮB�Ae�i&d�.��i�퉙{�(�ɶaF
�0)�bҐ����'�,�Qb��5����H�xb�4�!���'�vD��H��L����G�pd���a��A�xIk�b�<y���A�RYV�)t�t�'/^��g�Ёz;]��OdE����$��}�e厃[y.�t�ɤ+�`�{*��\U꒟t��'+���;�88�d��|�8:�l�k'�'T����C�I'�DP+����-۪��'N<��gZ0n&O�>2f	S�3U�I��s�P�%H2D�0�� άO�d�	�FC�o��0{5�?�d�n��8s%�'�p���'T�3ڎL����rE��'���`��i��h����c�
�'� �֎��l��#�5YRP�	�'A��iaeK"7�~;f��I�,��'�`&�^�M�܍���}@�S�' �aR�̈́NG��E!Z��	�'"���Wp�U:T��{,�)��'<�	��!Η&�̐듃/p�d�H�'2�"0�V�>�.�Ң�Bn�Z "�'o\aB��1ZF�C�@�3*;P���'ݔ�Q��x�:���7%���
�'.j�8L��1Z�,�Wϙ�
� ��'R�㤑�h�H�1W��2N�{�'k��J�Σ8��m����O֌
�'�<��hБ0|��˧-�@� �'6LD�pe�I�8yؓ/��=aj�a�'� �d�)-J�SO�,D��#�'����ɟ�\Bj AcF ���v�<�ӄEtT���vn^8 ���KDm�<�r�$����b�PN��IZi�<A�NHjP���UDr�A���^�<!��	�D����?u��P(�l�<� :up�-�M�h����
�l�  "OH��ՋQ�^2�H�SB,�и"O��vk�4G��|YƢ���9v"Op)D����� �\�z���D"O,���Pi��	 ɞẑ5 "OT|Hb�ɘOc��`�H�?	�"O�!��jP�NJ�8A֢�	Z��)�"O��c�J#+O<�@�
5�~QxE"O� ����TU��"�L�f��"O@���a�0[�2�ڤy�� �V"O�y��?\� ���
� Y��DY�"O<��i>E29�*B"+� D��"O�ph!���rĲb�ڰW��@���'6|eɑ�(Lo>�!d��f,�93�n�H�N��1mE'J/:	R�O6D�f<�)�'z�p� H/ ��a�S�*�m�o �}���@����$dw�Q�wk��st��En�*U�nHJf�^�y�Ľ0�'�$�Ze�O/�ٰ��Y 	C�ء��e���0�ٍ��0dɝ*:�}X�o̍��I�?}������-7e���#�o�@x0�K{��zCo�x 8�U��@��	�9F7\��0Ƙ�i��S���q
b�kd��O�ݑF�ڻu.X$��O��UHTgVΈqy��
���z��'td%h��X�~ũ��/�0|Z"aK�_{֍q��>�L=��E\�%�@�G��'Ay���y��	�"�n���&K�p ΐ���O �b�)��*m�p�l� h�:�l�}4D�;��1Z��?J"d #Z*@B�m�-_#��$`�P�g~�OC�NN�S�,�����!s��+.�1�����<E��ȡ$�0y����p�pA� �=/qO"��^F�O��)B�wƎ���+�0����5D݉'��W��A ��)�����ŎC �iAgjDkE�H��Gx����IH�'pV�I�o��Aej��0J	c|*e��>Y����~RUI!0����jK�v&�h�Lq�x
�4��������O�ӏ[,:�(Ch�8�ui$j�	jx�0��D�5�a���T�g��1SA�^5kC��1��Ј��	=jׄ|�s��)ϊBm�-T[�`�	Z,<3�ɇl�`�j�}��)����Aj��`��sE�.Ϡ%�OQ?��s�L�&�!��H�x(&��:vb�Lz	�'N�*C�.c��IRЎ�%M��`�=a���&GW2�o�!��'��i��{��x�@x�}�C��*��ݲ'*���N�JT���SB�Oa�4��.Fo��ш�Eш0r���'�2�v��e���2VLמ�*�;�'W�L�9;vva{�n��?���'��Qb"b�-S�8±I�"Kz��'Bd�`r&�5@-�����B�vY{�'�Z�2��-�t�q$h�.
�ฒ�'���*�)ۢ��L���}Sq�'�p� ��.~"��L:p=���'�.�"�ĝ,U���X�I�j�b��'�z(X�*�~z3�asj]��'�$�ІU�2V�(� �;<�p�'TTa��Fm����0��P����'�f,1w�'@��pH�Mw0ܰ�'�:��Q%E�h���٠@�bH#�'S$��fO#Hzz���cP�Be��y������E���+�^dH�.D�y�j6��a��.m�=+�����y�MS _�p)q��
UA6u���U��y"ǔIa�i��X�� ��L��yb��Nh�����	|��Ȋ#�y��W@�xK�Z�!�$��T��yҨ�Z�`��S�h<a`눶�yrKR��y�SH"�LEL��y�� >��aB���q����y2`E
>�����"[��Bą���y%4���^)^�+�Z�yr팗,�ib�܋}��m9֩���y�KcYh�lH� 2D赆��y
� �A�G�h�$\� V��R�"O�Y�!���
#��mٕ/w:t��"O�4�S��5얱��K�L]���"O���g��]:@���P?
P��"O��E�sV�0�'!�iC�"O�A���KER$ct�t��B�"O
�K �>E�uA/Y�w<|�"OR��g ��c]�-f�C �<�1"O�q�A�h�\�ꦁ��D@�Cw"O��7)PN�~�u��Vy�D�p"O�h2 C䮥�2��9t����"OBPA�m�@x:p�2Ņ�l�X�"O�@�@�D�_Ď��E�.�r(I�"O���'�G���rl�h���"O���B���S��U�!~p��"O�,��Nѭ�tS''�
Eq�u
$"O�)�o��G��iF�ӳMjj�i�"O�� cN�zA�e
�#��Q"O�"��%	�p 
� �-'�6��"Or}0��HZ���Ӎ�8�V"O�H�1OփXvj8Kţ�%9idРr"O&њ1����(��%DԬh$�8�"O���V��),%�UB��'��\2�"O��)�.L(�� ��ϔ��Dm��"O(Y�C���z��`��p�pIS4"O���$�U5F	d8���6y�b,��"O�h�FC��@ ��
�r��"O �(��P�=dT �d��7(�,`A"Of|S6h�Cf�q(�N�Ѭ��"O�q�c�/�>���)C%�8"OJ-)u�ȸ^���i�-���"O@a�栐#8:�G�G����"O��k�@׀jw.aP�c�8*U��"O�҆OՈ,]���gD��L���"O�!��EL�d#
-��C��u��T��"OlAh��D 5Q�h�sN��a�"O������,��k�X<b�
P��"OM�d臊B_��6ʀ
=㲤�"Ox�*�T�N�J$�Ph.#Ƙ�آ"O�����Ӣ=*���FĮ�,�C�"O̐d��N�.Y1����Z�Aa"O�"תQz�n�`�c=�H�a'"O�-��eA�px�bb�/w�e��"Of#AJ+�L�ȵFn�t#�"Ova pG��a���y1h.�\A��"OH����=nn����$[�����"O��@q�%7a�}Q��I|��{�"O�Mrd"ׅ� P��̳,z2i��"O����a�#[g�ȣ�R)H=��B"O��K����/se���;6���5"O)k��*��{�-T�9���"O�bU$�}	����*�s��IX"O6(B���+�P-y��S��6���"OR��q�ڊ!P�|��G 5p�L���"O����Hd�Q�G� Z�,���"O"T�kͭ����6�F70XT`�"O\�eҪ�*�*#(�a'x	h�"O��`�X�&�"�Q��L�1�u"O:pJP�]v����dH.f'&uXT"O��yԊ���貦���%8xI�%"O��t�MBY
�1��Ж>t)��"O� P�+��^ X9��B�N@��"O�@3����96�9qg�L̤�`4"O�u(�^�h��( pǲD�G"O� � ��� ��P���K�I�H4BV"O
�����" Q7'�� ���@�"O.u�U͟+]Ӭ���+|��lxQ"Of���J�B������'y����"O6����W+i�&P����]�b-f"On�bGh���z�@��)� a"B"OL�򁄕b�:���VTv $+�"O2��#EӚg�l���>C�]��"O�Q�$8_�9p�_�	Z9��"O���&\$մ9�����Y�Tl�`"O�@�G)˘�R5R��a2��z�"Or��S��"	-$�J�,֣eHlq�F"O� @�b�2 ��;A�ڙ!C<��"O��Ф��>��1�#l�D4�<)a"O��s�ǃ^��I�c��"�]�"O��P����(Є�ԯd���y"OT��u���7�A+	8Zm�P�"O�Y6��C���J	�^X�]�U"O���#�p_�tJV*��'�����"OY3d		���[�(�&p1bT"O)+�F�i2��3�g�mX�9�"O8A�e��dC' 	$��m8f��U�<��N\Uz5�ďY�P=�Q��l�<yV-�-!��|iq�B�^��,x�`�o�<!!'ڂL����7D&D�8`���j�<I��A>ldRr�H�tQtm��_�<�fQ��XV�'�ztKT��\�<Q�@����0
��*.e���q�<��
�,���,@�6�<�r�C�<QVD]]G���Ei�!C�L@��$^|�<!�g۔o$�B�X�)Z�d ! �N�<)�Y~��B&�M���+�*H�<q-��4�*�Gʐn+��Rz�<)QM��:�hJe��%�e�J�<Y��@���� &O�pxW��z�<����3.�B寔�����2ʃu�<9�̚�C^���V��'�jl����t�<đ�_�$�Jw����vC�w�<�'��/4 1w�\42uxêCq�<iA�IoFh��TK�p2���c�j�<A��Υ-H"�  �[�M���SoSh�<i�mZ�]E^���Y�] ��0��`�<�+�A��&�^�>6�a�#Yw�<1���H%��kA��$!xtxiuO�W�<B�Tf̅��Dף0J����Q�<��(��,��D�<tX�q�iL�<��f�2�N}��g��2������D�<�W((�����d�M^D�B�N�W�<	`]<��t*VJ��tM�}�%fO�<Q�D�5��aqM�x5�QŐG�<Y��J��b5���x=*�a��<�P*X�(F1)�)�>W4��F{�<��>�,�X"�JS�n=�m�x�<��˗�%@� "!RO�[҄�~�<�7�E-
�m�t&�q������t�<���@�5�(���%�"�ys��q�<� K�?䊙0�6RD�a�g�XG�<�g�0# ����&���r��n�<A��w�9Xm�y]���%�Vh�<��H\�.�
0�E�5
h:cP�<�Z0����`�=k����DAJK�<Y�� �7T�Dr����0�[��G�<������烞}�
5�3��{�<1���=\�"PP�X-��AZw
s�<� ��*f�J�p�0��D��!Km���0"O�r��z�J@��-�S�9��"O�ER �ϑ6]�����:[L4��"Oz�S�%A�
�2��T>�j�"Ol�:��I3�v!ЂI9t1�X�"O^-�0I�(8�h��Җ[�j�8�"OR�{ ��%oZ8��	�>�2|i�"Oh���\^f����*T��DR"OP9���t�����M	>��d"OL	�ĳ:�ai&H�<�*�)�"O�:�؄!�A!�KE��0"Otq�Q�N^�Kr��U}��"O�:c�ƒ3	���f����#"O�� ��0L�����T*"P���"Ov����ƿB��5{���!I���`"O��cAI8`�:��&ټ�IE"O�$��
>N�x��`U�%�u3!"OR`��!��B�hU#�d��3�"O�E�F��L��]��@� ��b�"Ol}"b)�A��Qz���#\��`��"Oġ�j qA�&;LMq�"O�q�����N�ν�ad�2J����"OA�4$�	V��R��Ŷ���r"Or��BH�#�,��e�A��N��C"O�X�!l �x���'c��Z�ĕy�"O�`+l�;R�@��1r��h��"O���Ѯ(�%�J��%�|�s"OT��׆�!83*��*ϛ)����'E֭��-ծ.^���DS�۪��'NX���OH�t4`�n�
�t�'̸�U���c����l��'
C�ęQ��$h&��
�����'�Ԍ�s��9l�X]cfǞ&q5.t
�'ԌH�CX�<N�Hv�߇i])�'@Ȭ��$޾Uf���[&`�"�'x6�;0��(��$�Z�;P���'7�I�4� B� �C��#5{F���'h$��F���MK�[��eQ�'b����ӧ4�x���HҪTvHb�'uXaR�FC?�4�ږ
��}w��'��C�ꂢ@|��06�1v�"�i�'�n���iV�����u�l�>���'>pɻ  ��O��X]t��� �N�� t"OvDh4
��/�:Q��o^(}�D"O|1P%��+3έ��c� 8	�z"OΉ��E��G�tx[�A&	��e��"O� 
�Jclź��\;L�$%
w"O�p9,��x��-�����J�0�q�"O���щ�)v�� �b�=mal=�s"O���lַ{tV}8���YXej�"O� ���NE�y:� ]��c�"O�	J'�J30���Ɉ$HP���"O)#ԅA�E�z��5�[8� 4"�"O���AD�8S��)fZ�r�0a��'g�p�BF�nfԉ�t�E�81j, I�aH�HY6��Pt� �D`�<gɴ7��5�vk�<\�q��Y�<�@�D�M� �
a��&*\|J�IZU�<A� %D�� F�#Q&ġ�LBH�<�#BD�V0�Hgt�P5���[�<aE����#�㗌e��E�g��U�<A��j(�љ��H�K>.؂ ]X�<��K�(���т�c�����[k�<�4ႫD"6IG�U-e_�8�1��~�<i�$(�|�j�K�)J��1��,Pzy�;O*c��|R�֮,7`XY�hH,���с�Kݟ��b#�U��b��~rt9G�b$�j�R>B\��ǌ�Gf��{dr�S��M�e�',d���>֦`R��p_�B�5CNĠ�� ����aG�ϝx.�B�I� ��p���ݬX����*�bB�	 V��Hi1a	v\K���SC�ɒ_�NB�ǔ*Mnf�2���Cj���4�S�O��#���b|�D!Y&s+q�"O`=��N+s@)����I��p�"OX]um�.b�����ܱ4is1"Od!hV�Ǚls��P�J�}��a��"O���*D�Q���K��S
R�8œ$"O��`�)�6�$�bK�A�DIp�"O�`��R�j��2*�"h�Y�"O�q&W& �r����Lh,��"O���v��)|��R��0j�X4"O$)a�ҷx%6X���Q�p�|kV"O|�"+�?�	���x
�$zT"O0xX�ٖ��}�dF���h
�"O���2��,@V�����7���	�"O��"�A�_/ѩ��Gv�RC"O�i����*5F4��SF�7j$@D"O�ݒ���J����"���c""O���RbR�v���U�V�;�J�W"O4!�M��H��P��h�<`ڰP��"O��R���}��(��'ݞ4���d"O�!���:���A@Ǟ<�XB"O� �\AS��P�n�+������P"O:!���,ST�@�C ��h��"Oj�S�6�*Hx���uM�S%"OrI�E�'�q�s�#����"O�$Q���$бG�#[�^Q��"O������3��q�}�*}�"O���P.�~�� KJ��5�Q"O}�T*��h&�%����4Qܬ��3"OĜb7eGU�b�+�*��8���s"O@y2��U�5lp⒪֒(M���"OV���W�!(��ەi�*(Cv���"ORH��ݺ~���z��M�S �D@�"O��K�o�@��Э�(	B�:�"O.� ���a.DU��{���h�"O|f����k�s���z�"O�xip���X�h�a� ��Zc�"O����Z��!����0b�F<�"O��!c�*�4�uE	��] "O�h��Ɔ�kt�%UO)tD��"Oe�dX�X<�9�B@��vjn��"OH\�G�I�R���Qo�0
j�p%"O�M�V�:q'_�8_�|i�"O�R��٫ .�0Ǎ>V�MR%"O6py���,a)6d+�G�R�)ˇ"O���E�M�Q��j#H�h���"O�� �D�aT�h�#��6t�e:�"O�+�����6�^�q�"Ozxѡ�l���˜-
|�%��"O*Ir���f0i葋J���3�"O8�s '�@�b�j��x��Ӳ"OJ yw��MTZ,��#��\l��H�"O&��]��])f���X���z�"ODt
`E��q��¡��
z����"Op��j���Zx  �Z�#[X�Y�"O�XaoV�A�"+!�^>�-�u"Oذ�C�2\�ˈ R�J��"O� *Tģ{n|ɒ���6d�U"Op]�q��O�yȀ%�8"$��"�"O�0���m�F�t�^�:�{P*Ol5���S�~w�,P��i��d��'`RQ�P�V/-��L��c۷_���c�'[H�P�_�xr���gG��XvJu��'�vD֠ W/��Y�Ř�;�ݢ�'o�  �m9|�zРm-^���!�'�|��#�
Q j3�I�e���;
�'��{戒�J�D}Q$�T�ZY��	�'����&�-ö���_
H�8
�'?�=0�MKb����=T�� �	�'�jM@VBĽQ�:	��"��N���3
�'����  0g����@C���'o��h�`�zs�!��l��M��e�	�'�PR#�={r�%quF��Z��t��'���d���)l^�Y��Z�3n���ȓ~�`�a���J>(���aHj�6d�ȓj�j��֬�2M����
Ϲ!n����(� ��b\ P�*������i��ՇȓFF����ߞJ@2�Yg�ֹ2h4��NU���G�uAR@�m��y9�@�ȓ\3���G_K�9��R:]�
��ȓ'�@��
5��d�Y�[o ��3R@�K��-d��X� /��QD�̄ȓ;N� /]!2�T��� ��=����tcE�
-G%��8��L�Ρ�ȓ�,=��Ύ !z �b��p�\��S�? �#�R8H�qW�ɵ*����"O�i���3'��m�%��Q���R#"OpQI��H{���s·9y�܌ `"ONx!"k #����lǓ;��$HP"OJ�PA-V�\��� O����"O����OK�y�q�w'T*
��1"O��k`����}�Ś:}�&�cF"O�\��Ǚ#7U<����F$FD�0q"O�0
��*���*vCJ�#��"O���St\飗b�X�&���"OxȪ���fx���@�\����"O�����Np���� @�;��P"O&D��S�o�:U ө�P/�8�"O\��/@^�Qfo�E*j(�"O�P����XO�� �F�T:�c�"O��`�NB��ɐуæv%�Xx�"OtaB�I��v�ڍ�����	�|��"O��B�R3Z;L�0� �3����"O �b1�-j�F�E��4��l�"O�i��R%�T���1��C"O2}��`T�LL�x�"m�vO�ݸs"O$-cÌyV$��+?N�1�q"O\���B؞Y�4i��#��%"OH��$뜡w��E�i�'L.�)A�"O&t���к4��9���$".ѱu"O4��f  g�d��� �Q���A"O��r��8O/j�Q���t�ZHy�"O`D���]	"8����?0�d"Or�PSF���I
p�Ͼ5�T!"O���홓* $�	���c�zMc�"OЅҦH�G<(���:�2�ٷ"O��
el7E��-��L��Y�e"O��")άu��i�-�"�4�2�"O���ԭ�.U� ����b�Hi�F"O|}�@)�%?�< �%�4R)p$"O@���D-v|Α㗯���Iy`"OzH��ɘ)ch0�E���O�^4�0"O�@;Å�w2I�7�U�i�����"O��H#�2NA��h����~�Zȁ "Oڐ1B�9���H�Wn����"O�����d(���h��Z��C"O����EY�%j���n̰ZIn�6"O�)k���m\8��ԧZ�h���"O�I!�����d3tj�3:�^��U"O\�
"�Ƀ9lı��'@�Ș�"OQ��S8d��!bJ;T$<��F"OVup��V�E��w ��X�;@"O�0c�Ǳ�����,XQ��u"O���4	Q7\ #LɎH����W"OVi���4�@����4!���yb"O�]xF-�2E��{����x��u8�"OȰ����"�nTSՎ
6ٔ|��"O��v(�!�晊fM]�=�t	�"O:x�1�v��,:�mT�!�B�!"OZ�
��P5b�@hɓ .6��JV"O*1BIűn>2�)�C�z�}�"O�q��ȏ�(7.�J�A��`kZ�YG"OnUQ��P�	2�Q���.aL
a�'"O���sM�F���⑩H2���!"O��`f�ǈ D�7�[�ØX�3"OH�2U�;k�Y��H��.Z�@s"O�ղ� �}���!(A�ؠ�"O�0xƏ�4|\�� �>0gpx1W"O�U`���}�8)�Q
�1\�c�"O� ��J�����h
U��GP�a�"O,�c�T�L��j�#tLby�A"O<�1��LV�U��i^8&C��C5"Oz��H�*FbB�S1��9BqP�"O�I�p"h}�Lֶ7ꐵ��"Olup� Ns����5��/� -�S"O��2e�k��pHd��}��BS"O�p���_t��cH;��a��"On�aGI�.m��$Ó�utN� "O@�� � E��rǄ�igx50�"O�ek7c��Wܮ�H3D `��"O�4���kl4x��#��a�^��v"O������B������ޢh\6l3�"O�p;���1R����M�e|�"O6�� "�7]�� l�PC"O�Q��EI�:���
6b�gZ���"O.1� �k����"�A)dL�Ī"O��)�C�P"����NƦh�D3"O�z%"��<a�J�	tL�lJ�"O�ݓ�� !W�
0g�o:��K�"O�u��&K�Ddt���GI 3�|�J�"O��6B�WKJ(÷��<m��͹�"O����ŜKN@�����vxѲ"O`��Di�52N�P��~��P�"O*���&H� ���*f���b���"O��A`JW8a��腫6�9�"O��be�6w=��H«�"��� 6"Ola���/���(f��!i
EB*O8�
�l��v�L]3��LyMQ�'u$0!N�V'fܭK0����(8D���GA�U�.̨4Ν9yS|��6D��a��@�R��M�P��6�`]�!D�p��8.���c�F%�`m2D�8�w�մ���TC�!�6}�F&D��qq��b����$�V� 	hg1D�L�b�6WB�;6�ZbHV�ą.D��sB���]Ss-�:`�(P�*D�ܡӯv�\qѧ��DVo'D����ЕUW����f�����%D��I���?A�<��!B
�)0�.D�t����r�����'M���u24o.D�@sP�\���3�
K���&8D��`M�+=�@1��v��=I�L6D�8�� �~�z)+UeE��a;ŋ4D�����J���q��S��#3*3D�X��Wk�h�*��M^Љ{�M/D��[�M�:R+O�k��������y��@�9C�@$:���Qe��yrg*M(,q�C�N
[[t�`�)�y"� r����\6W:�0@(���yBm�,Kn�y����Z�*S�݄�y��94�6EA�`U0�^�b�.(�yR�YE�@�#$ ��>Xc����yR�)2�!'L�w���[�)]��y��D>vM6MсȌ�025z�n���yR� ��5�`��F
�T���@�0=��ƾ�٣!c�6-�l�v�x"�V	P����ۥ@z�x��'$�1[���i��W�_�Ĝ�e"߬=���֭�K���f��aO,u۳����(ORѓf�?r�=���+��P$U�Y�@�ۯ*���+ޫ3$��f���Ms�,Ȳ��O�Yn�:��9KuC !fHepƔ$6�d���	`�'��	�JZ�PB��uQ���6��8@%��<��'���P�G�:
�"D�P	ҾǼ%!�k˦9R�4�?��iΐ;V�d���<���h�����%;FJ0�J�0B|���>�a��(`K (ͻtA�6AX�R����\h��n�N���&ԛ8*�5�s���Nb��T̏?%6�{f(bo0<����:D��D�u�� y�G)�u�2F�E?�>�0E���OP��~�t�'>��O����#�</(N`�w�A�_�:���<���Oj��<�g�N�.��p��:X�8�bbkb����۴ ��[���h҂n� 8�B-��`=r(S�+��W�iWrV����?I�>AAh�W`р槅�����i!.�qp�[�Z�SC�]��vBO��I�<QY�w�Լ3��a�6m V�8R��-���0��8Wm�p1
�.�(�0�,�&�y��TJ���N��)���M��v�D^�y�+O�� ���OǥW9?�2{%�P� ��+J�\��$<O���O���7%��9�\�Ti҇D;:�J&�����޴�䓧B�'�M�
��`$��GS9%�� �Տ�i?	�h��1����'z�֣�dX��E"*F�����TI��s���D"�4'k�+)�`@Ճ�'Pa�}1��d��7��ݨ��6@��!�BG\�n��9�]c^$T��<�K5��F�C��؏:����1�,�FW�9h7�UQ���2)|Ӗ�!g�'}6MId�	���Im�ɯ Q�EEV�z=�RN�$ s~�If��h�l����{�d�޲t��ڢ���M��� ~���'��6����ʧ,�f e�i�����:DU�SaH�X��u��׻�p<�!	�m��,n��+c"�>&��=z0��R�̸A�Y�[��HaL�>3��(��@W�'k�����h�`���T&$���CI�%7qv2�J�jr��PdG&���3�۽�O�p�'�'��6��T�,)�W0Y�l�xfK]"u���O��I�X�?�O|r�B�a�4R��H��L�An�r�<a��L`�,�0)1;�$�:�JY7��6m���]�'��=AѮo�2��2�i~ݝH��@�r�0:��1�Ԑ!N4}b�' ��Ē�2�XɩhY�qЛ�� 5�,j��O%p`�ͻC�-Ҕ��>2]�;�}b�A
s��%����4�N�{��]!�L��O���u����"9��#��7G��#���'��H�q�6%x�\�$8�ɂ���ݹf�*5~	�Ϡn�,��'���"|�'"�<�g�
��� )s��(f��2	ۓ�M#Դi��ɲX��?+X�����]t���'����"�'�'Ñ����   �J��%��	�<y�Nт$��X�D�*.�I�/�s�<���5n��xb�ň�R�+�H�<��-\�4��t��F�
5�<!�JMH�<�3a��M��H ��?�8�I�o�l�<�ƂQ��2�T�J 4��" �@�<A���.!��I��d�ăs�<�� XX��dt�Q�H��c�l�<�3�˥B��uX'.Q/5!��KFNDk�<a���v�	�&Q�i6D˧`d�<�u�C6)ʅJ d0�ɐ��a�<IFOU�e	XY����� OHW�<�mM0ˬ�"�j� �P���W�<�f���|u��A��B>����}�<Q���l90���%i&���z�<��J�}�%�� � UA�S��|�<1O���@wl�5��
�d�<	e)��BJ@J�I�
���C��Y�<ѱ�yVp�sI8d����\�<Y�B?�}p%O
�M���*d ZQ�<1u�4:��+�S@��r�/�O�<�@D;�VЫAmQ*|��R�<�jX�'���a7�TR"�%z��r�<�c�D2��qKŏ22�q��C�<A��@ ^��	�u��Kz�@!�lt�<ᢄӸ]���	u˕5��@���H�<�*ʱbjl�k��S <�p��3`�C�<9����B��7'��3�̌�t��A��HN|��κ[���#����1��Q�ȓx��,����6n�U���L����ȓ��dJ�
�YN��3��Ć�dh8�i���k%�4*�Y�ȓT��  T	�*�8u"q���bL2��ȓ8��l�`���iӸ��v��h��}�ȓ2S���o�\m�.��X��ȓo\��P��x�ۆO���xɇ�|ae�d���ѓ�	�a���ȓP?�Y� �|`ኃ���P�ȓ?j��c /ݰ��:q*�u�:Y���������oŰ<�ì�1A"&t�ȓi���J�L����+�N!�ȓ}W I��Fa4Ą��.ۣh�\�ȓx�J|z��K�B�0��W�LT�A����C�D%5z��V��I|`ń��	rp`U�av��$	��w�a�ȓ� ���K��O�D�c@��'贅��z����q�j�����@�*��'<��g�*b��p����;"v<�ȓddȔ!�&7���j�L�a~V��?�8$�w`_(e>��i��>����ȓ!H��g���h���Av`�m���ȓ��)k։ћ@D�A@�<#jP��S�? e!�I,#�Z}@��}�i�"O�(�WgQ�J�^q�n����aG"Oh��u�XY^�(�,�+WD0���"O"����9Ҙ<�+�(KE�!t"O�cĮP�n�j�jA5 	Ȁ��"O�-9���j<�y�Ald���0"O��4cN�%�qS5. �[B�� "O\�D#|�}z�,߁,��X��"OꅘwԚo\��91Ɇ�zy�rb"O��9�S!y���X#��6aH�д"ONQ��cY"/hRRJ�6""���"OƩ�&%	�@�L ��19L�x�"O�t����W2�ݡ�̊�,�* ˃"O,5"�.~�� Am/>���!"O�X�d�<c�0(�K]+%5pi2"OTI���['=�NH��ґ+�M�6"O���*�	���sS�R�XX� "O�5r#��*�@�C���ZJq9�"OЉ:sE��w����Ck�6#�(��"O�5��kǺm�|��/IH)i��"O.�ѕeF�[Zq�qJ�Y�t;%"O����JԘkd�9��)o.�)�4"O�e�;?�P��V��HhIS"O¤ �Z�굣fm�0�y� ��Dq�,{go -`\�E��	�y�ȗ�G�Aӈג[Uf�����y��A�����VWe�-�w5�yRŇ�Ul�X�$i�#x�(� �7�y�ET�WwH��)�'~��IsN"�yb�ݛV��r���s}�e�m���yb� 
d�s��Zh������.�yRl�7$1�9K!]�v�I�V&�y�-7�Z$�\*WdƝz��1�yRL��C�6{�)N �(�Dɚ,�y¡�/5�m��?@�;��:�yb�\�<=�M�mT�woH蕂+�y��MnD,1�6��!s��̓u�_*�y�LB�VK�RB+d�*q҄���y�&�=<��eXF�
,+�:���u�
�'���EdX$N��\�qV�$/���'H�a�e>}f1q�Պq����'�@���1]�<9���2^���A�'^����l�$T ��FC]`q�'wR� h�JV[�I�Ĝ`@�V����'S��]�ʘϘ'�R��$k�DC�|�"�߼�`F�_�, �">_]"���	�g����?�s�'V���NS�N(ɣ�j[��!�r �3��{vF_%:�zŢî_�7Fq˒.�ȩu����8���DF�3q�-Y"�؟��4��I���M�3^��@�&�O�0&�`��d�Sǘt�!i�����6�hO��s�'T��x�&��]VA
��;9ິrI�(*�4YΛF�'�H6m�|2����iĴ+Α��H���%Q�6"F$S�����M
ϓ�?A,X�}�؁�$ޞB>E�#� �;��R���l*:}(���`�Ц@.O� xDy"��!#�av�L�|�1�$�YO@��¤�Ot�B�3$���%�I&L�-`�𤉸l��p�!�J�E��ͺ�-I�A�:��6�'2�6��y���h�Ik�ަ�����*�2����q�PyZqm%D� !$jȩ<��mxF��8���f���"��� lӜ�D�"PIÿi�;0�r��&E�
�`��!"��)�̹G}�'S*� s(�q⌳�K�������oU�jW�1K@��R�BHR��8A��ݪ6�Ѩ�(O�-sCƂ�B��ȱ�l��%�^�]�f|�e��Wޔ�&�?C,%شL>o�XlFx����?ɔ�iN��ɜ`���)#�����!n��7�O��d�Ot��?9�c]O6���gm��n)ְCU�,�t���J��~���G*���&��T@�R�4��яy����'&�O��D�i��H7�G�k0zm"����!iB��'?�Z�W�$A��#t����5"���n���%�0Y���(�Dg�V�!ɉ'~���ĹB*XeC�f��2�"�S#���LCӟ�9aA�"e.R4�Q,�F�T�HњxB�X��?���if~�<�� H��Ր2pu1r���`�x�����O��%�$U��SL-��i�5?��d�� 1Ox�mڴ�M��Q�f�i�"(��NQK)j�ۢ%Ͼ}����Ѩ���	��y��J�e#��鉚CEB<�Əi~ �L��0Ǣ�R	$,�5�-j���0��A�4�O�09�!%Pּk�H�(Np��X���@>>X�7� Q��A�,��Ԡ��I�p_´��鉞J7� ͻn(�ҵ�i�i�jH�5�5[GGQ7h��V+�<��Y��>���O�6͂�a��)K�Ol Ҳ�6s,d�?9
˓g����aE�qTRl�3B�.F=`d�OV�lZ��M�I>A�'��O�`:"	�#[��������k� ��2- �D��4��<)��d	�h�qH�a�ҭ�G��U�T�¬[�JA%��1O�ތS۴0>Fͪd�2�(O|�2P� �vD��
YD�2U�GO�����wAa�	�+��I��x�����vv�"���5c�Ts� S�W�$)�"��j�VQSC�'�67m���	iy��'�e}rF�z�|�a%�$��Ճ� ���y��O	�x�R�	r� ��)
�F:�O��(�)�Ϧ�'���Yw��;oZpQ ` @�?s�a*����1'�O@)o8�M������O�˓���³m�}[7�^)@�Rm)'�!6!�D�	FIL�ˀ
[8J���!�e�'{t�$����f؇�MCM>����<��w�|�� ���]�JV� JJə6�Epͼ��#沟D�r�J��M���4���)<��R=erYr�$���8���I#.���9mjV����;��l�8N�w��A���Ͽ[t�Ǜ>�͈�����ڤ�A
ߦ�1� O -褆V�$B��@pNB��̳"@;�s�����iS��S�alaȴ��bp��E�'d86�	֦��I]��MC���21��7G^�u�beY���[?����d3,O~T�+�'�� 3�W<H���A0����Q�4��0���\w��C3e��y���ЦO
�4 �A,��6lO$��S�  �M�ƽ�# S^
\�cbJ�;�x5���l05�V(�D�S��4y�G�]\�)�l��d���
qRQ@ F��� aeY?	��n�2B�O:�k$�;g��"�$�X�p�1'�����c���Ɵ��ݴ|��gy�'����OX(`�@���%K�N�[�v��f�5$�$(�H*z��``Q��LC�bқ�i�6M#�d�;�N�)3��j�)+ù	>  ���
�+�r���1c���t�fͣT���>9b�iY�6�+�}��P�B���t�e�Ǖ*��!��iNRU��������M[��$�j���E�v���	Ie���2(D3E�Dp�	����yݟF�IM0_O�qaR�TѤ��,O��+&�:J��5mG0U����r_P���CU�Vɼ�|<�4&�2U�t�ɪ@�h���E);�	('��4%`�J�_��8&��O�I|�	���ߦ��c��)c�2:#.��A;h�1f/��j���'M�t�O�e@��@iQ�4����x��h�,���ئ���?��w�4)�2jQ2���8Y�Ɯ1�ᄳv<��$b�R���O>�1o���(�$���h8��I���D��j`�	�AZ�xuBÖZ�h���PwAs �
���tjPlH=X�����/	W�|��C:?�Dl"f����iC�I;la�6���A��mseoو�b|a�m�+,����ܴ*!�'��'�O�7�24;`���OU�j��i�&̓�T�!�$��bʨP�7�UvĈB,�#��B��fhӆ���p8�i�P�D���+M�,�1fG�Ff]��3��?��	0t��$�r�It2��ٴR,-A��FB��Kt�}�^�QO:D[��P��d�O�*wOG�FնlC�'r>��1�BPoM�;v�OJ%�uoҾ4Yqh��	��2�$Q��a��4�?�Zw��=a�E�-3��KR҇YB���؟,�'��)ڧq���D�U?] ���a�ԅ�	�QHSl�z���'o�U��p�KL$ [�&�|p�H䟸$��$����   �ޤBS���%P H����S�pӴ7� Ц�$��+ql�?�&���}��U� @�?>�p�I�?>驢�A�N��lRAˡ'�~%�SG�ھ�����/!tl�q�W/Q��	1i�H���Ͽ��&�20f���$��`��G.���[��Dϴx��*Y�e����Ư	�V*pI��
a�s���a ߪx;�]+h�6}�R����u��[�'7MBiy������l��
���p�L
�, �� ��~�'�O0#=q�+�	{ϼx���`�����L�g�'�~6-��5���M;���]w��TP�	`LY1��	��(��Ȥ<�q�*k_�f�'|������$8=�3��4\�U�P���)�>�⑅а~�+�e=;|����0)Y���|bGM��p ܸ%�&���	�p0�'G�*
�r � �R�>�1��V�1S�Кpu��MF���Ix��S�@�E�� �U�@�s��O
in����?q����$	�ܡ�k��#;|- �H�=��>A��š+� (���M�Pά:���~6mF��q&���?a�'OT�bA��!xь=�4PM�m�3�
�m�d8�'�'L"� Z����5K�.Sh�BlĮ9ਨ��"W�����b�R���v �b��@�r�I�#��2dÂ5A�,}@�'�H����E�+d䁓��D;�(W�Ղ^2z�j�F/�V��t�	�4�l���T��(�#q@͕<��P��̖��M�����$�O6ʓ��O64� ��Jm��'ަGLl��'"�����3^���3��j�!��'�`8b�~�(�O�����?�L<�%�# .  �F'Sa��=b!����H�fz�Gy�[�3v����5�R�O1P� ��GO�}��{pcA9e���D+~6��t��O.9�����7Ι��H��~��l�"�'aZ7��~�	ҟx�	H�������KW2J�F�{�`-x`�)��HSN��`� ��V���%q�����?ɴ�i�R,y�^�m�H����'
�7��Ok��)����E�S� �GbρͨO���/6?��0�,��M$<����M�)�:@��':�La1�Ԗcwf� ���?i|�J��I����0�m�P�H����'^G�L����{��M���TE�� 7��4/�
͘4�4����I�MK#�O^0#�T.�d�g��<�N`Q�OX�d�O"�L�~B�i�!$��iCC ?�⌓�kG(<	���!���8#�R�CR���C��v�"���i#�	�<4 <#޴�?K~��'�M۔	R+6.}�$)Cj$(RT��A?���IJ���cF2c����]��M;���jx��#/���S@��
U��$�xQz-2f�x�'E�#�pD[E(�~(�R�M�!X���3��	ԭ,q�=Rƃ
6Q�ɛ�^"[�'�����3��l���;��qOF�Ȉ����c�ʇ�l��ty�'�)&����"��1��Ȉ�	���YA',O�6���y$�� �� kR#("X�cåН=;���d"��&1��]�I^�'3&�� ��$'�3%9� �o҆'�H�,�$�|�B�n��a'>e&>e�$χ�O�.�beN�.
 �!���|�?YL<!�ܷn����!H�'G�&�H��Gx8�<z�4͛��'�x6�`�� "�u#��h�|��h=J����V芡�M����䍭i0��"��  e��TZ4ũ�!*�
��*�Q�^�	V�_� ����,���i럂Y@W�8�y��A�425�u �=D�+���A'�Dq��(dt X2�FT%S� U3��/�S�d��U�wI��`�e�p*�ݫ��ά_�~]�dG̦5x(O`������?���M��&�b�l��)UZځf�? �O����G*e�*]5jW���"��$��Ǜ��iӠ�O����(�u]�}Y�@I�jg���Xa)S��]�g�6�,<O����R�HLcgo]5:������ RLŉ�H��Q���\j�d7M�3�Y9Ō6�u��a�bK_'i��[�J������ܱ��9���ѱo�W�S5iY�j��Ro�'/��;�k�!^$���<�<�A�?�?A6�i��7M�O�ʓ�?!/O��\Ӱl�"j
"��+��Ȥ"Ed��|�2d;6	I�!�݉u�Q-�Hi��|��-n7�'��ܺ���߉#\ l  ����#��' 6  �` ��Gm�����fU+����'J�u�΄+� !iB��M��4�?��i�Xlz6'v���ĭ<�݊�"��nV/V^b�QЀ�m�.�,��6i~���$�<B߲���e 5dXȲ�gEh�k4Å�d��8CbkI��+� <���e�3MpfmY dZ�Y%K�3�\5����.\0����)9oD�˶H�~nH"<���M՟ ݴ0��O-��,�
��MY�KV�b�μ3g�?�R�d:��O?��p��ūgy*�r�-ϳb�x骓�'�t6��ܦ�o�({�	�%�נ*�����%)���ɼ
#V�!ߴ�?�(O��쟠O�e97�S�4	^��+�*�P�r�CPl�E��*5Ҩ��*H�9L�@ԆS3 f�����?yE~�*P$�W�v0��gG*7�D6�f`Rt��|4l�v ՑF��,i&�<�1�kl�s=^���A�5 $\x����m}�v�ǋ�?Y��in���?�E�ܴ`<�:�ȝ~�!Pd�߭>�d���?
�f��$�Kc�m��K��y𴉸vi��Q�\��4B��&�|��OQ�N�=���hTDW�xvZ�sF(@�H��'"���1�xӸ��$^�(༓�Ŭ�����/��F0����!+F�����ڰz���!�"�?�ˁ���t�O�Pq�G	�'���;2���@%}^3�828�+ѦA;�� j�&ј��U��-qR��j�AE�D�ȵh�e>�	#*4���y�N<����?	�O!x�G/8�jY�$ɣ������>���I�'X�ʶ��F4���f��t���4֛��'��7��O<������' T�����.v6�B4o2Sx��8�)��J���jϓ�?1Ӭ÷p���c��^�#/���2�Է0BF� �X����ĒdH�BТY�;8�HDy����b�y!�&:P����L�nG�I!�mY
����#����xuė	f�\�8��d+ R�E��H�D놡^����"�������ē�?�����'���N3���m�%)�� c$Re�TC�ɰcqR!" ��%{�@u`b�Fv�ɱ�M���i(��%6;X�Kܴ�?YK|�7+Y�}���!l��!��Q��Ob��?y�"\�`��$`Z�S[���4'.��w�1JKB�P`�L�f2(Zr((s8�ҏ�dH0G#�x1c�+]2�J`�5E]\���#�.�|�Z� �|s� �8{6!z��I�D/��ĕ����ٴ�?᫟�+Roִ2��� MS��q��ƈ����'w�)��pXw��\�Ո��D8���pg,�O6٦�o�4B��l�n��\�B�b[�r�d�'~q���'k�'9�O�|(��  ����G�^x���{yP][�� T t�SA$no�<�ȓP
,H+dM!�ŀê[�:�F��ȓ���bAD�|���&�f�P}�ȓ<vh�g@�o�,;�o����ȓ|0����9u6����/G�[���ȓ�,p��P,y��A�FY�2�ȓ!{�-JTK�0@5`w
^�x�ȓV`�AXVN��\���#��]"�ȓa�&<�5�N�HK(u"䭉�}L���#��!z- �Q�
�sfn���o�څ0���-�P(�d��97+b��h�`�KFO� �����(J���mBT#Y-j
T<�ӧ�4y�L�ȓ2<4@`"큪8
����AOo-*���P6�tX�
��Ia\]Z�CQ�>C�`���Pzt�L�����N@�E�Vm�ȓN�&d���У8��XBG�bfʵ��䂰�ѫ�-耰2b��L(�ȓu�8�(f0v�P�NZ��0�ȓj`9p<�"LZw�p��\�ȓ)v� �����'I9u��x�ȓAq0oҼj��1s��Tg�Ԇȓ����<_��¶$�WȲ1��"|�M�Յ�r�b���+Ie��ԅ�S�? �YBS�>/�)���N�e+�EB�"O6EJ�`Z�4����H*�ј�"O� Xc���W�B�ć1&|�`* "O>y���J"K���矑vܙ"�"O���)]A�2QH@-�^ܫb"O�uB�%��ф��+.�d�#�"O"ۅg֨g^ �� ��m��<C"OF����6N�S����ap"O�t��Ԟ�`Z�4}��3�"O����Y\B��8nӢ9 2"Ob����Hq@�����˸�>�C"OШ3���D
��΢���"O�%�J�n��K��N�֝��"O��+�Ǥpƒ�1�C�a�Ԅ:W"O�I:0��
c ������$���ے"O�0k����>�>��sN��#�2Ր�"O�uJT�J��]b�m��5���{�"O�i
C؅8Z����N`��"OPh��^�r`���!��=@f4� "O��d�=EJ>`(B��GҔ�!r"O��8��]XM���gj%m����0"Ox����A�,�d���=�jD��"OL�� �[�E�V �G�&4����"O�d�(��L-j�&�"Ƶ2�"O:р6���`�VE	 E�9�.�qR"O6�)����V�j ��?2��"O��kT�A�=&0�wMX�z ��U"O�50ƨ�����J�LUt
�A�"O>I�v��!�Z0F�D.,3�"O��*b���ŘFO�d�\��"O��Ȇ(T������a1"OV����1Q0e�f�"��qu"O�x�$�B,+\�DE��3b�`"OXTrr*�pU�	��V.{��"O�a����\V�`�Fzf��;�"Or����H% �%�[:I\`c"O
aP%+vu�l	��R19�e��"O~����m����w�{�"O� ���L%,8m##�[�Ի"O.�b m��Gh܌�C'U0I<P�#D"O��h���`����S��t"O����n��8/Hy���!a�j}�V"O@�9��a�D���F�	��P""O��� ��<�|p���ƥx���"Ov�{�
U1\�8�s�Z� w�-�"Ot}�`IPX)@�Ǜ8�%ZQ"OL$�ѭՉ�>%�!��I ����"O��cT�f���o �L>Lă�"O�`�t.�"Qq�m;T�	L*ր��"O�� �.��d�x���/�<��"O�d�ˈ�!�h!��LJ��H9�"O��0GD��]��hQ%��!'��F"OD{CD]� �l{�˂��z�"O��R#��i	�) ��3)( y	1"O��k��6-C�z�>U��S�"O�e�aϱ	F	���R>Y?`t�0"O����ˍI�;�LǉG(��"O>��$*Մ6%r@Д��DD`	�"O��Qa�T/]ބ<1Ν.aΞp�u"O �h���#춝KTmơ�9	F"O�����Ŋ!0�<Ƌ�	}�(3"O�|Sᮏ2(k0X+���5耬#�"O�,Т��_K��	�g@�4z`�"O�%R*˷,y
e
�%�|�P�"O� r	)A��@�)��..�\��F"O�DY�gXjO�zy�ÅȶbD����)c�搵;�N�A��)�@)��&��z��T}�8��*�n�^=�ȓ8N9K� H�r��(�q��_�`�� E9�x=���ZHӒԅ�!�	y�T7~���T`ȉ=TQ��z��1DC�@+4X�vaQwf�Ņ�*��a�� 68�q���O�2��؅�zB�����I":��,���4&��i�ȓ��YHWl�#;�Y���t=Մȓ=ؙ���g�6e��dE-p�"��ȓ
�Α��hY4qB	�1��,q�P��\'�h+��,q+rP7�èF�HL��3����	ڭ$�f�ZtJ�go����"%(��S�J�R��)^1��L��0�򑑣�͖En&X���&�@!�ȓC�v�{�mɎT����D^�)h+"O�q'�F�$n @��+�
r���!�"O��2�m�:Z�Ȩ�u���!���"O���uA��A2��Q�{��4"O�(7��i��$s�,���#d"OT�vJ�5��iB�NZ9zli�"O�Xh%��$��[��^u��P�"O��s�Ȉf��b�N��� �"O�����L�G��)B	T��X��"O*]+tIH��|("��'dt|,[�"O��
�B�([����� KlL��"O�5�k¾8� ���FN  ����"OJ����,=�J�1SE��+��""ON�0��p���{�D��YФR"OH�#s�?g'D�%Ɉ.�Dԡ�"OԱ[�CX�1��ypdS�a�jR�"O��3�0 ̦T�-F3LTF�j�"OZ�ӏ]a��t�Z.:�p�"O �E�A
:$�8b�]/}�(��"O�yrD$T�S����!�?<��"Ot���� &|��D��/�=Z�(��"O� {UR/y�T\�S��} H�q"O��qB��5�p�g�)o�(�"O,� b�BEl�g���"�L,2"O*=�5`2c�<�g�\�U�~)�"O~=ST/�J!C� ��/s:��5"O$i��+%V�����5�`��"O���4�U8M�$����k���e"O��\${�:Y��&����u"O�i��Vb�-�sbWxKd�Kf"O��
�ش>4D�@b�q=�5B�"OVt�E.R�m�8����4.��0X�"O�Q����
.�Qs�FX"ek���F"Oހ��I�Y^�4c��V[\�� �"Ov܋V�R+TF$��L3� ��"O�e#w�ЩQE��۵+U3=�� �"O<���G]kl\��
�+M����"O���F'�kq���t�Ή0�\��A"O)�P��5%��!ш��I=�y�"O�A�7Q�� �!]b�8�9""Ojp@�Ϡ&p������"X��X4"OVu���yn���a��W���"O�XRFE�e��@xp����ekQ"O�m	�cѨV�����U+��u;p"O�B5d�<j�����)� =�@X�D"O���G3D�Z �㇀Yj��$"O����� �����ȍgM
�� "O� �x�Ì^% ��}H�ԽH�!��"O�� ��J�<� x��ɼ?ʈ�!`"ON�`�ȕ$Vw>���-q���"O�e+2nV���"�I06���R�"ON���A��Q2t@B @:N��d2�"O8xr�̷m�&Ph@J���A{�"Oh5Cdl���H{���+�� h'"O64�����0i����
Z|J8!&"O -!��}��R"�́w���v"O����Ʉ$\�� �"
Q\1�"OƥǢ�
tK�(aO-;u��1@"O�ݒ�a���HI
�@V(�@�"O�ex��f�2,�H�v* aK"O>�sI�Gax=�,�D�"�b�"O�\z��Ѫ^�b�`���'K�,�"O���r.��&RVd���Ի�fh��"ODe*�-�) G"��P�(t��"�"O���	X�y\X�R���0U,4��"ON-)�JͿR�"�&�޲�4m��"O���
KPB��H��B���"OLI��2}A����L׹
�N<�`"O X�,�]��Y��lƅʂ��e"Oz��g��mc|i �&/[�}�"OrH���\��Ӏ�'J���t"O�M���V�Bo�Y�ꊢ2�l �&"O�$`Aaܦ4wRٙ�茉E�TAK�"O�飀��?j�������*t�'"OF��I�L9t̠�)
$�"O�1�&!y�� I�h���V"Oy��c�o���{1"
<
�D��"O��K2�>.���!�6_ &�x�"OhA�V��'Ar�h@�/#��mHF"O��beM@�2�
�I�ڡ�b���"O	iA�Ӻ~)>L���J%��a�"Oe���5�d� ��Z����"On��SJϽC�4q)ƾs՜+�"Oh���� p���#�A"t%��r4"O����1DQt�z��
93v�ʐ"O��2�
8"jh����ں*��"O��(YԘ[���$�Ĝ��"O�m�;E�1���"�R"Oxq��5(2@�T�èl[�"O�ѱ4����>���.��5��u�R"O�}	���� >A�do�7�H��"O<X8 �ń}7h`�$���1T"O
 HuM�/9���7�}��M�A"O����)u�x�K��[;����"O�ʢ���|�x)YVH�?�Rp"c"O�$g�ל+��8��e�;W���"Ox$��@��W�2(��N��L�,�yүR+ssh뇁=��� g��y��d�lLA�GF���u[5,ٕ�y��H;3�VqJ��\�a��#��yRG�
޸41���3IL|p����y���	eZ�b���@���Jܭ�y2�ԙe�ΡCPKL(�	�"J�y"d�>>���SE
M*��4����y"i��K��Y��!I�|�F ��ހ�y�(�8��(p`"�{X����^�y��C�c�ʽ��a��ql.�"��$�y)�<�,�ɘ�o�T]30ȕ��yr��0���Y�n��i 0L�
�y��R�r���*�l�/mB�`g/��yFФ>�ؐ�!ʐ t�$H�ƃ��y
� d�����|n*�+V2M�(�r"O��c��t�X��º%"�ٹ�"ONPp��<S ����
�L!2��"O~ْ a�vjX��*˹I��s�"O�}!��^�a�:y��"_�KLX�y"O��zǣ_����g='g���"O�DZ�C�:z>�s��-EPr�� "Op�e�xkr��S�G)�Ҙ�s"O|!+ %��5�l���D jC�"O\Kf�w9��;�A��%����"O�yJ4D� ����SA]�lᐉ�0"O��r���x�S��O9@���4"O�
�l�X&�aՍՔ{�!�"OT4��PE��4bR��|.L�cV"O�D��k�
.�@����1+��1�"OAY�OL4-�P<�U�Y*��"�"O"d�n5 �F'>z-�,�"O��$�ؼwx�mJ����k>P�*�"O2EI��\]6��UF�8?4��C"O�D�+�	�Ґ��Z4�Y��"OA�㢟*���:B�4/ &���"Oj�2�ǳ;{�iS�d�)[�^�w"O9�h�3<�����3QxF)��"O�������4��	�<�"Jt"O5�pKjGȱ�tH^�dкU"O�q�G)L�=q�FDz5!�"O�����0j���s�l��
š���yR'�E�ХPV��&[�F�q'��yb��0yy�I�cX0N�bq�vBΰ�yrM��~�!�׎A�X\�F$K��y�Y
wx�H�`֟p��Z&n�#�y"[d3<M[��T�44�6���y".�8AL&4*#�X2x��[vI�yr�7{�<*Ǆ�u���R��]��y�e�H��画eH��VQ�y�,V�'2.�Aw��S�Y�v��3�y�+ڙ)b����ɶ|�@�	��yrEO5����dD+o�ĈUŜ
�yB�{
iC�`H�b�N\���_%�y���_��\� �`x��	DE©�y�$u��I��?�R�S��C#�y2ID��`)`)G�	Mvp[�F��yrC��?-�<h���{S�i;RF���y�@S���K��Ůu�q����y�O�%'�H�UŔqK�B
L��yrK�� �4!�"�V��iغ�yB(.'�(����'F�1qD��yB�Jzf�0��)�&D� �x#i�'�y��N�B������7�܈���%�y�ʃ ���`գ,2� E"l2�y����W�>49���U� �� ��y��N�v�T���ǛZ���G+��y�JJ�T��� �|
�P�f�y��(\�:�i�v�:]�DJ�y��=zl�h�eĖ e������	��y2��Amp����U�h�`�P��yB.Ҙ\�ҀC��a���^��y⧌�F�u��똍ifR�A�,O �yb��?mB�!��v�R�����y��'�1��Bk�f
�dW��y"�L;f�8X�	O�6�@t@�"�y��"0�4�x�垻d5�)	Pŗ��y�ܷ�H�I��Y�op��1�H��y���-}�5��)\�m��q�QB��y
� x-���;�h]�n�
/���"OΜ���K���۷��\@�"O��@'B���i@�K�IV�"�"O�3��s}�xV���,��ɕ"O�l2D$�j6\��$cG�^���"O4\; �4�ltC����� �"O���IH� ����@�~���8�"O�%̊��*	�
����%+�"O�ġ4.B�2~�X *�9u���#"O@��DiE�	���2q�$��"Os/��k�=�gB�wW��;"O�]�wE���d`ተL��"O�|c#oƕ3$���aOX�3�����"O,x;�ϐ�:��;i�$Jh��Hc"Od��1�	*�XE��	�d$æ"O ��5�Ȫ6�"����Ղ6�"O�,i�r�Pxz`&ٗo^���"OR�Q��8jƖ�SC�S
zG��+�"O^��r�Y:c��,0��S�v��E"O˒.�l��˘��h��`"O��E�%5��ك-ԿK��9�1"Oܑg�U�]���$�ɈT{8���"O�,�w� A"��#p�Z��"OfI"֢�A��xcm^�5a|��c"O���u�ִ&�Lh� �wrQ�'"O��+�EF�R�N<�R�Ғ)�\��"O���g�> �A��3]����"Op��u�\�O52Q�u��nڄ""O��R��җAJ��4K��o��`�"O�0s$�
V�T����u�Es�"O����,�v�Z�@�!<�� �V"Oj��r+D�O$�E��O;��$)w"O}��'BM����ύ"k���$"O��� ���A���8��D�Q�R��"O���G�6GX�!�MN�5t�B�"Ox0�(յ붸��b2[ �"O �K0'ɍJ�p��bѪ:%�5y�"O���&*��=(��"A�&��x�"O�%@c䓵v��ѐ@&&:�u"O� ��[�Q
^�� ���X{�"O������U&��0�I�*I[�H#V"O�����#U&т�g<R1"0�p"O\ ґ��|^��jf���}̺	+�"O��)�������,��@}��"O�M��_�0s���L�V��@"OMXIR�T,(-���ɵ >�KQ"OF�����~�]�u)���dP#W"O89�d\(5��(���?^G�)[A"O}�p������O�`� P"O���Q�V	��V��"t�T	�"O�5zw��#m�Rmj��(|��3�"O:4��B��o�|��G��Q&�3"O�e[%��%&J�\� �	�$��i#�"Od���у2Q2x"��O��&��"O�a��4{s��aL�-QȲ8�"OHq��K�3TCf�ڣ�
{�x���"O�y��^�fv�pQ�J��0�f"OBL①]�(�w']0�jу"O���a��.�6d��ݐH�����"Of�$O3#�BC�
�Pzl-{t"OZ1I�GM$^}j!Чl�4j@�а"O�cd��/�I8�)�T�u��"Ov��.�*'�^ �6��l�5��"Op�����(��E��4^,Z "O� |t���N��J0��cT�t
���"O�y�a� @0p�p�B�0���"O\����
h�ca�)+���{7"Of�p�
�'�D`��K�H�h���"O�}JD �/o�8�vL�?p�1)�"Oppze�۴{�*��`�A�fxf"O�R�$JGh��qb�e��L��"O�m��� -�ʁc�b�v]��$"O���3*E+L[vua���"PL2I��"OV5zP��%��@�����d<>���"O�!� %k7�p��M=<,��kR"OV�9�a�Ix���$��K�q"OhdY��ioH0�(M�!�a@"O
���%ՊD������(��}��"O~�С�М	��I�s�:A��
�'G���v�;��L�"c��z�*�h
�'!$K�|��11˟DԆ-�	�'B���f�Y$k�����<h&���Ug)S&�pM��	�!ú��q�+D� `�&P!f+N�[b�Zy�l顫)D����!3#��� ����?U���G)D�T���Hպ�y6��vdv��k:D��8�kM�9�U1f��������8D�xӥd�<X�Ai��?B�T[�(8D�T���*)
Z�2W�F&0N�lB�;D�l(�#F�Nz��C�Ȓ~��3PA9D���λ"D1xU���$-�0���5D�����_<'�b�� Ę%���q�2D�1�n�'����}猰���+D�9�T�*O�P�o	�2�~,a��*D�(C�3�x�Kg���@� 
-D�$[3�(;�P������x�P!� 5D� �� �EÜ�0S����aB2"3D��(Sg��R\�Ф�e|\}*"1D���7��e���1�XM�v�i��"D��&��#���C��q�d�2UO"D��Z�Kڷb����'���\P�֠>D��+c�\�]�^lIGl,e<��PK=D��أ��Nq,����� �i2`=D��S�i�XT�C6E������'D�$�Qo�aLxs�F�i@ժ%#&D�,�G ��O��Bも4K��@d�(D��k�����T�C��e��H���$D�t���-L1���P��;mb�1�L0D�袅%@�d���gC���X!8U�-D��5Β+C���0�����*D�\�2 ̚�Z���I�eF'T���#	0A���Su�G��29c�"Oz���cgP�*�I�!�ƐzA"O��S]F��P:�%V�&�d��"O�5R��������?�b�z�"OАr#��)}��	��%{���r"O�0�� ��:Ɋp�Ưf�0�"O�����X"-L���\ d"O�<+��#��B��$X6�A'"O`P�A"E�r��lh��U
��C"O��`�M�).��Pq	�;H$���"OrHj�c΄C� �#
"���"O��ʦ��EC'*���R3��[�<��+A<Zz�
 ߬_���q�YQ�<1�#��[�P�˴��$&�� ���K�<��AO�xS2���^�@X17	J�<�4ퟑ�t�B�D5Ճ�b�^�<���?�t(2AF�Mv�5�6�_W�<� ��4�d��m��'M&�"O�W��� �#MМ8��)f"O������9q1"\�1���h���r"O�T��*¼N��RIV�&�V\��"OD�Y�R�~�T�k��^j.1�"O�ᩄ�QwY��I_�����"O�1@�3<T��j)I�v��1"ON�����p3�j2�"�z�"O@�q�,&�9���7f�5�&"O��Au��4��<-!�:Ȣ��K3�y�¿#MB�a�n������y2�Z�R*LЁDh��JF�� ��R:�yB/чnA����Ғ�R1����&�y2��_��X��EU�^`f�����yR��b����U ��b���!���yr⋺id���X�l���\9�y�E�&�R�1��a#�i	���y�d���C$�*���Wf��y�dO���uѲ+Y�u����Á�y�(�3(k2����R<,�M�pB�5�yR�C�b$�I���3|a�x CJ�y��A�R�\蛕���)�Iȇ���y"'��~��8�фX  ���*����y��13ǂA �# �zEz2��y�m\��P��]2I�f�hu��9�y2�	��li�afT;�8ŀ���y��͎[2R`r�\�a���.F+�y�Fִ�*}a��o|V,�e���y��F;C���䘆c% !����?�y� Q�H���(��(l:���yR.lZ� ��"]�MO��&� �y�V(d�AtO*F������y���Y�@S�Ĭ? �K���y�	8m�����6a���xQ����y�Fnw�[W
0�h���y���%G��ು:wv�o�y���;���K͓D�|�෮���yr��5)��Z���1���(�8�yҪ �c���P�$I���l����y���KnL�a��9x��ެ�y��&E���0RlS�{u�a�� ���y�X�:��%��#ml�#�%^�y�	�|��t�e�b����ޘ�y��,��-0���0V�\ s��y�IϨk'�$��.��Ld<�7吳�y�(F�	��U�4�h�舠�y�.Nn���Aټ��B�#�y����> ���(�S#�:�y�(W�\���fIп#�V�{���y� 6lb��I��ޙK&���yrC��`��BCQ��։��*�y2�oA�� �� rb��y����K�R���'G���a����y�#�2����D�AE�=�2�yR�E�-8��&K�� �i/�y��/3��ЀG,_'���A��ybl��'{�IK�{�z����y��X��4c4A^�sb�C/���y�X6�D����c��ɋR%�y&�'��qpr���L2nz����y�`���S%dFn���T@�,�y�hĲz��h�-j �Q��(��y��	�y�('��T)�dj����y����n�)�$
��H�\�灈�y
� `��� JOnݓ��րN���1A"O)Ȗ�t��$�'
Եb� �"O�u�/��|Hq+�!(���"O̵�D�HV������E�w�RL�f"O�Tiad�D8����*?pǀ�yT"O�m�p%�..@RSd���ȅB�"O�Qz1�ܥ"��q�ύ�5���+�"O|�r$�M-C�X���-:�sP"O�{t��R�9{��K #a~u�"O�A���YT�~���Gi[����"O�7ǃ{��#%l�/HJ��&"O��vG*t{q�vj!df�a�"O`�	���tЁ�.x`����"OȈ�d��	g��Rv�E�/P�Y9�"OR)���Վ'ϴ��%��8Hv��"O�(�Â=��UY��<02�Ii�"OʱH�mE(d���K�>;�n�cc"O����o�$����ˇ]�ډ@`"O��9AL7G7�h*���!�1P2"O�H4fB�	�����N��l��S"On�q��#J��鍒<�\�9q"O$\��ˑ�0�Q(��F��}�"O<����uA�p��G�(/���Pv"O�Y�� ӭ��d֐3��р�"O��s�*Zj$��Ę�}�U+4"OTA���_�(���>~G�$sW"O`P�F-��lSHĘ��Z7��"3"Ofa�����h�z��)V(�"Oi�V�T�Q.DT�1��7��Ч"OHx�1�˵tΌ���]��(HH%"O�䃆/G Τ�Rr�د=���"O�lks���d�)O������w"O����Cʢ<Z>(CCQ�
�F��B"O*U+S� �b��}�V�\j�(�p�"O�E��h��
Ep@1��p�:-�Q"O�8��],����'�1;j���U"O�ي3%�.x�0I�		MJ�� Q"O��́�$�`X҉I,u��"O p
�@Ҭ]L���(3�xhb"O�Q� ���D@IxfJ:M���s�"O��10	�N܁�4j��A�E�"O�(	0��4oC��A2Iz?hY�"O|�I�B(�.�sH�!�\ɨ�"O|h�q/Ͻaf |q
�b7��"O��Q��P�p�A�iX,N��T
"O�	a�F�L��B�H�--�0IP`"O���O�9�ִR�&D=X�)x�"Or����*)���
�+P�I�٣v"OP�����l��)Bʄ<?42��C"O�Y[�I��
��X�i@-D:d� �"O���g%�"UX��QhB	/*> �"Oޘ)/Ċ����1A�*>H� �"O�a��0T���g�0��"O�<�w�p6lʑ�Ϳ~�l�R"On�*�X$ `����p�^��"O��� �y@��G�W��b`�"OZ�x���wl���^1J�n�G"O�u�R/(���(�/�%"p5�"O��7�J�-�LY$iG� q
�"O8X"�YjK6�x!��� y��"O>���$	�~���mA�)��"O�0NFmҘ������`��e�e"O��8�Ƙ�_��R%�]u�H��"OΔ��%ʛS���Y����iED���"O� V��c�R� �eN�+0V\E*O��:`�QZ6�� ��[bD�`	�'�0T�-��!y�:!k�!E�lDy�'nQ�4�L!Ba0��K�/7tS
�'��l�Ъ<#�L�w�M04o��	�'V�X����0|�@�,�̥��'o&\p�FM
-�֘�6 �4z	�H �'��a�,�}����H����'�!H�Y%CתYhE%M�q!���'�5� E>��*B.��@*�'�lu�CȘR<`������'��7]�!����R���'�pPړe�mX����[�(m*�Y�'��D���R�g��(�� !RnD��'6�(0��-~�$��"ל2���'�rXh��;@�\`2�5~c0�X
�'�TY�a��:K������y]�0
�'el�����m�b����G�t��9�	�'�`�	v/�Z{�l@VJR/B��`�'G~H�pL��a���A� 1����'�.�@�Z{���ʡ���)�l�H�'�� �\"Ř����Ų�e[h�<������B#D�� ���b�<�����) Z���ʓ=k�Y���i�<iԹT�Ux3�G�:����b�<扭\"� �D�8Pa�c��S�<a������'�7"t�E)J�<�2��>o�MB��6��t+��F�<Q4�G��A��CW+W�N���A�<��GZ�n�����"s�.�x_h�<�$f(c��Ȃ������ F�|�<ɢ)�-#�`Pcf,??��(��̛~�<�"$I�v�<���8q�QGF�q�<�$+'!�tx 	�fW<%�E[G�<��+̨nź����X)F�N�<!�J M'��a�F�|M�iF�J�<��`�s��p�T���U�eZD�<qEU+3aR]��� �~zT����J�<����6x�*y�جk�R �W�E�<���<e�0y)�K$W��ۧg@{�<I�D�D54�ԦI
�ћ��N�<�揕�k�X�ʆ+Ы%D:9���H�<��	� yx)�@+3}R�FUE�<q�#�(9� �ܮn<��'�EB�<�ɞ�mRZ0����d����N�u�<�7�@�r'��c�F+�v��&k�j�<�g�a��R�� � �#j�h�<Y��\�'�U�uO�;B�e%h�<) �H�T�T�j$�b|`0�҆�c�<A4jݔ0SXQ�gE1�*xuȀf�<Yu�Um�H�[r ׄ`2�3�!j�<����
E�Q Ꮑ�s#��[B��c�<!Á�&��l0G-܈Q\�"L^�<�w
���)��JP��3b�Y�<�A��=�&h��*�T�2�EM�<YWe�dh5��/�<B�ᛁ�Pa�<��^+6Y|ڦJG�M�l��S��x�<�Qa�9ƾŪ���+ �q��Us�<��DE0	��A@'H�Iy]�!��q�<I�.[�c��E�:+N�8�rk�m�<�6!^�|	"�E^!?��ӳf
T�<���	�bĄ�"�3lb�ZHG�<�Q�*:��Z��Tx�B�*�E�<�/_5 �8U���WvDRF��{�<� m�,�:\W�D��͈�G�f0�G"O,]RfI��oTR
K�V~ �C"OЖ��6M�r\	c� �]�����"O�0����:�~�Ł�:;�a!�"O����a�D���	��Q�BZyP�"O:ŢD�1+�a
e�ٹrLfQs�"O>6X8[QBD���A:NtB�˖�)D��I��1L����	�j8y��%D�����*�|�����(Q�U��$'D���A$
$?ʉؔ��h�	���7D��@Oq�p�$MR�N��3��2D�|(����qD�3�No����O+D��JǨH<NX���� tdH�R�)D�\c��J($�&��ӆSP'@�� 	$D�L��� `�.i0��
D8��D�=D�0�$*�Ơ�G�,HlmZJ;D��ҕ�&w�|�{n�&�8D��Zt�ϫR�R��+�)X�����y"���=����('�PiŇ	�y�@��d֥	�N_!�@�@��y�+�8q�Py!��K8�4���Ы�y�.�	he$��0�z�8�Qk�
�y�)#��xr$	�q��̃�Γ)�yb.�&M��Swd�)4�
�+9�yr`\/ΗO���	�'R�R����ȓr���zҦϪ(�� a��=-j�ȓ/4�r�+S�c���@Ɇ
ްɇȓ��А@H%l����G��x��8�U�V�
A{�!ڶ`N�-�j�ȓ\rV��f.���y֌֮S����� ����c�XW���"O��S��@33�e��㊁I���h�"O�-�A��8BFř�S��P"O�����5����c�<���@�"OT�x�/��B牰A�̈�#��fO!�D̓R��;��+nq�:Si��N@!�d�k�ZM8���3q����艉p�!�D^�OTp��A�֐_���h؁F�!��..�@R�����Ĉ���y!�d@�@W���VJ�Zמ���r!���L׸	���.z�$�YB��1k!��o5�Ġ�#�:-�x��%�߃F!���7 q�8p�)M�&1�G�F�>:!�$[>`4�4s�V�%k��#Z�/-!�N%C�RM;A���ue�����Ў;&!�F6��{p�֑'��4񏕨B!򤚲[��D %g}�Y'�N�a�!�$�R��	� C�a `c�ȇ�!��V���y�� �9Ib%Zp�,�!��2t)�=T×3 �����߇�!�DM�zt���1~���"'�P�v�!�$k��@B!h�|xp�L R�!�LGI S��3���#��J2�!��V�e%2�#DbP�4�ФQ3�Ԟ	�!�S����FGC/4ؐD�RI�.q�!�;�H�DE�,/ϘՒTg�1�!�Đ�ARt%hV	��6�d4	#���!�$ &�t����!M8��\q�!��ӂ�@G�ڠt&bI �h���!�$�Y8]��C�{@1ړ��mn!�dD%:��}�4�۝G��Kq&
7D>!�U�,�H�E~�<`��e�R(!�$I"[Ŵ@���s�f���y!�]9C���a�Pz�V
3��K!�� �X�kQ�/N�[s��-YN\��"O�
� Ov�����(@�"O����	�=���ġE�/�Ԣ'"O���T@֓3IL�{�`�{�*�"Ox�Q!yd⥂�"n8��"O���W�		��Xk� Y6�`�"O@ �U�=��R7`*@��rb"O��ض�V<:��`NT{5(�"O����
�{�鑖���x��b"O^uzbS��t��5GP�/�L�P�"O�TAS�L��I�ec�B��Ѓ "Ovr2��Hp�\A��V�'|رZ�"O����B�)Hb��[7nW�\�"O쁃Z8����9Ū��$�<rh!���9�&������x�ѦInd!�F�w��u�M[�x;�Z�]b!��0�A��I�� �Ƙ�B]�'_!���:H�S䞂gq&�����4�!�D��\�J��R�R�o��V�3O�!��7</ƌ5)�4{���Vi�L�!�D����H6❚*?6ly@�]
�!�������+
48Z����B�nZ!���+o(b�a�m֌BаX���*|�!���ꀤ@�U��$��UKָe�!�DF
k��J��M�e�V�RT�?y!�ͺ�pt�&��0Z����%\9!򄝇w�\��	+��@qѪ� 4!��Z��%3�d��k�4Y���R�Y�!�$·�DD�%̔�8�` ��_Y�!�Ċ9�-��a).mЀ�D�@!�MxJ�+6���ɰ����g&!��Y9 a�P�4G�7' s��!�d��.~]��+m�%Q'�5�!�ΐ|k�q�u��3��)��2L�!���?�v�suD�6Ge`J� �K!�䈸DS4�@``��bFB	�c�(M�!�DW*n�HS6��BA����^�!�d�+F�"r����@�ؐV��	�!򤞅RPP���U&e,��#G@'6�!�d��)r`!#��d'*1J,I;u!!��	L�>�BB�34�H[BL�!�M�ck��x�f��?�0a4�ɨ'!�$ZO�!;B搞K�นĪ�Q�!�ۊeX�ŸK�;����J�!��֠d�9!��/}�r��k�!�D�;6.��BHں#$
(# -�w�!�F�$�+q��V�Źvl5�!�$� �("��[�L����"*K�!�DI�(���ԉ��=��c�)�:l!�D)@Yf�����9�T8`�BU�P�!�^ '2���௄�@�^�!�Q z�!�՜a�ޱ�s��Ovq��.ޤg!���U���E�-��K.�?k!�DQ&��0jƧ6�<=ڡ��)\!�ȫPҎ�	r��#�ʤAvl�B\!�s:j�w�J/�d*ъӱS!�$į<�8tR��o�T�@�o��d!��B6x����iT�����>�!��1!�ͻ�鎽+��8fM�6�!��GK<�	 �B�KI|i�U��X�!�d�-��y��M
>+f�	�)��{!�d�v?��+�M��m#he��-1Jq!�ď�5�i�ϟ�\(:���v�ȓua�\��B¾pt$40f�	@��,��S�? �{�6S�
M3�?���&"O�I���:JF�Mk���#����"O���)ַ��h`5P�>���"O���b��n�Ph�bч�R�J�"O �� �طn
9;fB'��h�P"O*�r�9#`�`B�e��"OpLA�^�F@\tZq�W��@�9"O��Cs`�������e�xh��"O
�����q� �`g�_�vDX��"O�I@I�00��9��B�?jh9r"O���%7�b�1Ĥ=��U(�"OV� p�EL�Q���֒l�<��4"O�8��Sl:$���A�||t��$"O�ArAB��a�"'Œ_�ް�"OV����L�.˸�����"]��"O0PQ���NW�[&&�)v�� ��'BLy�OFa4+X'FB�)W%XZ���"O��j	� 暝����O��Yic"O��K��+�@��������T�'%��<��`�iP�T�D�
XZ�*��{�<�$d���`q�+K640�_x�<q�nV7;��J�i��t����cF�Y�<١�1}:)ᒀ��=�2tCr �U�<�b�Q49���ׁez,cR��N}��'���@��"��Ũ��-_��c�'NP-Dy��ɋ�M�d��#)���y��L�AB!�䛫���Q,�m�n��w�/������7�"�U+��t�Rq1���=iw�C�	ʟ�*Q ȇ7W��jw�4<)4�Z�Ow�6B�IDUrA�U�R����_�t����ͥ��';r��݌I�tC���W
h9��&D� �m�x�"p���S8-�fMh����P�~�|© §<ǎA�����I�<�d����E�ȓ3�(�@��L�}Bư���^�Q�{�֟b?���<ygC@�n.�k3��H����Y؟�!��'���:2B�,� ��d���^ h:���4ON��H*�&�� ��	,\�=��'�O�h2(�'_1�u�uY�0�0�a�� �!�$�=H�ԑBg�طcA�qUQ�H��z"�Ѐ��'_�|B���.8�	ZT��&W��ȓ:pؚ��}��<2$��k�0��>	+OܒO�pu���*��h�㏘8G�D
�'��P@��E�s(���T�)_�b����'Zh�q��;YE�W��;JT ���,�S�� ��wE���QC�Y���J�7%Q�$��Ig\83�I�z5�!ar��0� B��0[{�Q��郙I DX���`��D�U�8�+鑐^8q��")%�����DPd�Id���O����+�s
��)W�,�I��'1x�jGȘd����
v]�[�'P�����̯/��M ��Υjz�s���n�#>��	t!��X58�Q%�L7@����TϸP��,�7���w.6R��ȓ#j�P�ĤQ�zP17԰Z����ȓ@�Z��� C�#�Y�e�f��%��F{���,X2L�����1�Jd+�	 �hO� F�ԫB�KhZq�Tf�|7���G!�y��H1C�G��<�*��-��M�`b!�S�O=��fm�8T�z�: �X���gQj�<�S���J��Êٴ� I�sK�h�'��x����
}���c���k��y2�	N`D���ş�W��lgK٘��$#�OBԛfb�<e%����W1��ӗ"O������D�����>�,=�"O� $ukU�}��鰐�
�B1��'u�d�<I�L�0s�H��΋^�  �F�MM�<1�E�90�K�,ĉ0�T(R$�M�9�v����)���1
l�f�3�"}A�=�ynP�s�P���,
$���ʰ ���FyZ��O�2�3pW�D��$��"��17��Ӧ��>�����b�Пl �M9�I�&̸��0O~��d%P�"�1DN����ً�lZa{��DQ�oV(J��k����t+�s4!�ۑ.E1.R��D����ժ5<az����|�ɁcG�gi �x`�^�;(!��ԹG���� �=;w
�� �7���'�ў,Gy�� ����X�Zp��ƨD��yB�Ea�n]��Ȥ}���(�CB,�y����dM��LүLE�h�e�9�y2��<�*�M�I�(��Ξ)���y��'

P�c��[H0�1��B�'in�@�腹[��4��A�j|��k��?��h�-~��A��ɒ;0 X�F*��q�V
�i�����Q��
�<���KY�/� �X"OvXj�Ȍ����"�d�nA�v"O�\2v�ѐ'&�Q&�I8^��r��IU�D2�S<n��M�2C,��`km�(��B��,0�d�`�ޅJ�lA��7	U����l���p��J�|�F�]���((D��0�&�9\����\X8�5�!D����õF��×C_G+,p��)D���h�|.�DSh�:�� �&?)	�/��lXQ/*u�(�vd
�g:��Ez"�~*�I���:�8�"��B����^�<�!�G�P������&P�(xb�C[�<� #ٲ��X�
�v.�S5�~�<1��W�b�&��.��L�^�kg�Nu��p=1��D,Y���B�G	�wn ��f�G�<)�Eͼ0��`ْj���2OF�<)��K1xu&H��㇓6�>\����G�<Ѷo��;U�u�G�y��	`�F�B�<��b��%��@Z�ع�D	���E�<9�f̣6g�i���2�8RE�X�<	*e��B��/o���	��l�'��+ҧ*Xx��E��JC�oPY�ȓk��9�j�>e���%P1J�ȓG+z9����R!�dK�Jj�u��`ܓ2̬`چ�Y��l�'+@�D@���'��}�F+-���Ȥ�@�rR�8���_,�y�
͔#��x #�qgd�`��Σ�y�9RV��B)f���\��y�<'��y���V�g�~	�`���y�"*$��;�/^1	���KP���y"��/ $H��NM�u-FY�\��y�:<��� �����XD*��yB��$%���i��J?���^'�y��$_��(���0�J,��#��f�^�!"��SNjC�.�z�w/Z�h�40�'�1����Q��䉨�?�tW?�����B]0$����o�����@��?E"Y��Pn���̄�4L��)Q�*��ȓeֵ: G�"�|�0�P6R���7oܥ��@��
�b��]{���ȓm8"@J�F��[��i��̓8(ԁ%�<Ӕ�)�ӅF�UȀ��+a=��W��[ϠB�	
�Z������x���h�Ԑ���OL�"~jA�]�S�ҡ$_?Wz�S�`�y2�T�@����W,еl#����O�<�'&���f�A
|}��9?M�ܴ�(O�~n:� �-�V P;v�p��J�%��e�'K�'haz��؞_��%�%lν{��9���yR�׆�bi#�C�
#dT�r ݟ�y�a���5��h��_z�Q�n����hO���e���i|D�C��p=���Q"O�D�u�ř)¼���SO��"Ot�f��Ѩ�:fX���Ȇ�i�ўb>�O��9P��:.ll���0"����A������4��أ$�J��p`�-N"<�	�I%���)U�p��d���S~ �ȓ"�)�f�B#y&v�ؤ�؜nN�͆ȓa�@]q�l˱n�X��@�3&`%��*Z e�6�0�Q3�F�4UӐL��B�|"���pt��.J41o$�ȓo�"�0�(��D[`�tQ'q:����3`����R�J��hSںBF�x��@�
��ǃ�s��{��.i_<��E���8֏Dc������+m���ȓR���:�	�T�Z�*�c��`����4M�y�.����d��k�#T��z��<q���4��X��d��I������l؆d��8|b�Ew&����q��l�f�� 2��6 �0�ȓ.����Ǡ�0�6����qk�=����#W6P�'"I�z(�a�f�c�<���;�:�L�	Z(�tae�F�<AR�N-l�	s�_ s:��!b}�<�f�&'��� D�0��T���M�<IB&�G^0���C�(R��)�F�<�R�X2��� ���^4�K�~�<��� ���Q�����D�<���<���sA�ڊZ�]��m�B�<��#�"i+r��,ֻr�}�S��}�<A��A�J��{Qb4CuZ�{2kSq�<�"�\��ꆃ�,T�[d��b�<�T��<b�0��0A�(q��C�<	H�?eƀ `�	�M���q�J�<ـ� �=(]�G�E���d�q�<��n�
LN.t���m�t��A KY�<ɲ�ϸ$��a�m��4�,����~�<ɒE��}��0�`�[�id�u�\y�<q����:l��KR�i[�aA�w�<Q��[��.��J�v�z ٧	�q�<�'U�q��VhT5;� �rG�i�<agF�~[�ͳ�G��e&��P�'"T�����n#�dA�+Υ;�\�U�$D�P���8c״�@�o�B?>t��%D��3�ľ)v�x ��V�p���!�O&ؑ@�V(B`�Ι%u:lj�Ï	u㸼�R"Oa�V�ǻ)2R�Ð"�x�U�"O �3�]����@��d�p�"O"X{���+G�,ɱ�V8Kh��"O��a���/Cmt��¦J��L�zU"O�E�b��4���e�(Ŭ���"O��j���X�2!c��F���r�"OpŒ���/�T�ps�ĶS��A�S"O��E�>�f�
���<oOhS�"OSj��Y���W�U!�"O��:�Hƛ")僅�0e|:A�'"O��@�#rx09ӎ_��2s"O�ĹeI~>u-t�4×K	�re!򤟾��d݌��Ix��45l!��	Z)�A�f/�'P�¹'	 K!�����	��|Q$I��4J!�� �"DZ3y�(��,R3/j�5�%"Ov��P�ٜ�:���m:tR�ջp"OR�7D���<���!Hm�L��"ObE�Q�ݡBm�����y�����"O��Ƀ�V�5���Q)�:�2d��"O�YpgN(d|��yp�7{��L�@�'xj��^�>�	H?$�(�0�hQ�Q�QȦC�I)3⸙�e���@SVH�	E���O�HCf(�D���"�;�'21�ܳv�^>&���Crɖ����	�&���Kb���Γ��
���	%�4ySN��>���qH� "	x�X�'���)�0�3��F 'fn��fg�9�(DsN^�@��s��]�4�\�O��ЄL-��O ���W��E�xMp@OU�g�>e��-C ��`�k�\�j��'�D=�D_�����,s��%�7˔�LN�������^8��'
�����Վ<��Ղ�%�:Uה���ie��q����Ԙ�����%��֜p�g�/\O��I���]*�h#$G]`q:5� D��b�E�	4D|�E �'V*)b�X/].�PSć ^nm:%�� F�瓩.��a� O�Tu48
�N� �N�?I�M?mB��`�\�?E��D�t��`��EU�Ĺ��OY�����[U��a/�������2�̭��˫|za" �(�f�ϻ֨�YǊٟrưiJ�Ҝ{���'����M�p���+� ]n���K��y�S�j��	@E�#�,�"4��i�u���Xp��	ӭGB��FAۗ���Y�嗠�6�r�}�ɽE��8��H�"
I�P(���'���
�-�(9���	fF}2"�I�D��,�2�!C�L�$��!�6mE;C7��I�#��=L�;��,DP�#�p3���{�(���"� �,L�|�%�G!�����iȑ>�8��	I_�n�xKY���(����p��\���F ����Ai	<�>�0gHQ91d�xR�ڤ8Byj��2��O΅	�GA�d�8���J�
���p�\8t��C`J� f�t [����yV���'غ�>r���t[�%�GN	<}��cp��e�zc��}_����;v4HH�OV�lq��s���'�v����
Uњ�k�lW8
0���n��?��Y��x�����	�8��
4i�'��.1I��1�˃L��aX��x5��*d��D�_qO���Ǘ�9�,�+�0<T��" (N{d%ʃ�ӻ �H�Ӆ�+����G":� �c��3<UŸ�@X(OxV!ig(�f�lYB�H�t����soԓr�y�NA�!c��Z���O�SJ�B���"|�ԩ��f����v@�a/�� ���i_�y���l �;�4E���c�K�8�LU�C��R�A1��Gy����2N����͜���O�@���(- ���5w�RD�9*����c"	]XxH�@��o���!B�*5�8��e�X��˚�"����#!Q@H��l����6� ���;q	^����8a���b��5P���"5䎝BvFͿh� �O�H(*�٪bj�6�>B��:ddW(q� w䙄(��;M��DKp�B7���tJ�a�a�F��r䄗)u1O�"2���C�&	it��8�p5H��Ϩ �P�F�ِ���d��BLA�6-9�a]<�j= F���%΢�����V�`�&A�L�4�P%n�P0�(��5�Y:$NI$L!Q��D�
�|\����Cތ��ЈLiD�jԎ�|0�� M	H���D��C�tp�!��D̤�DL	OoJ�R��>���w�B5L�xt��L�h�j��~eԕG|B�)�,ph�I�-\�~�q�ֆr��5����Y�,X|]H�
�^hhEq�@"~l�B!%��v�6�̮���A&v|�rQ%���®�&>�jF��;U��Y	�@\V�'X����F	N��Y��?�:f��C��U�&�e��a_�]�| �rF�8P�kr�P>��5��.o��+C��#�y�!�[�f���'f��e*	{�ѢS��}v<#�4�J5�0o��Xq����OgE�锒��)��'��*;��@&����!b�Aǈ'*��5� �Z_�A���� 2d�����/Y��u�&�C&��9i��\x��,�����)B�_gx�Ȓ�U9wnvI��X>�&L��F�*&D�[��W�)���CIÖYjf��Ժsefm8DL��9 �E%M�j�YI�씩F��s�[P�1O �3 �R�ɸ&���G�^�*d����@U�C��%��*/#�0�=\^-z��^-։������`�!F��ȅB��-%�5p �<;��jQn��$ԛ�A!uK�Q�ry�4PFA���C2/WV�x�	�c�]Ѱ]?��"��&���Y �G�JJH���6%TQ2��� Xf��d��m���89 DDL�*8�Mj2��5E�I�sӠ�a�Β�'���"�Ɵ:��Z�D�<M(҉\�e1xĩ��#E���J�d	/U}ph��hP%l}��5ET�Jȶ�Q��d�Շ�XPR-�4l���lP!	�Wrڅŕ�O��'��*��)"&� �5��CpH
�jɕb����΂]D���DF�6��dYƫ�q+� ��$h��c�TN� ����{�:f`­LT�0)Ĭv���2eAE;e<�*A�ŊB��'�l�բ�	�0��UΟ�T�8� W�@�X]��`A�țw֬Z��W2@	+6%ۋ�����L(a���9��T1`Y����	�|΀
�U1@;E���P0��jE��L[E�N#K�����'�P`�q 6S9����i�D���lc��c�I|����%|y
��bj�#{}^D�c���:"Iҗgњ)�x!��ivj��[w�*��ӈ͖U���s��y7���9lf���슝E�,��cdG�h����CF��z¾�9��>LjP�.��=��Q�j���+,6��
`�0��K���(,ܠ��[. �V�!3kQ;f����2��~)��2 U_�(,��b���B���!ΜJ��$����с`�}���.�L���qNL��'�O�J���4�mӂ�1A+_��IB��39���"�,=���!&�*5�H>�偟"�>� ��;,X|�#ޚX���f@�8.�����۞s��07�M?i��{Q"���a猀s��6�Y�/����.�q��g �k���6JS�1�P������
\���<s���[G�1Q���S*V��f��92�^����Y�����5P��) �i�% �`�T�G,O��K�a_@��D*�֩D�j�d��1��OL-�eC�!���'H���Z�w���xA��`�⩃� �n����:AWb��e��(�*���O~�{������ςT�����!s�ʄxԭ������I�U��*gZ���'��&��܉����P~������ �&DS�/[)9�.��0���?j�=ூ�����cOS:X���&�0�4d3�/ۨ:�&�� 5�� �0�2`)+U�I�Cp�D�U�	� �@M� �y̴�C�-yn�x!����p/�4��,CԶ���K�'q@2Y'BLO;J�r���-(��MJ�p.�<��E�BѺ��+�d?�N�7Bz��p������AK�qy��B!7gH��F-����3��['8Jc�'�j�BQ��8���6
8钲+J�i�}��Bd�41 r)��Z�T�,�Xq��2ȨO���g�`�( yV#�Zfʄ���'��QV�a9�(�F�	.	����i��a(G�`�ҠqQŀ�8����!�؝vVBaG8�άB5)�T��qG'st����L�T��xboŔD�t�p�g�8u۱k�i�XPq����M��,\�o:x�Ѣm�	,����@�I��Q�VC�*�ꡀ�螇8���F���D��ѺqM��
��u��,!lO�=)�!����,�"b�� ^,`���S~ʤq1�J�'L��"V�w*��'l[$o��"�՜]$r��1'�yǼ٢�$<ٖ9`�G�w�Z5sӆ1�6�dI	"C��i��#�9]���Q�h�Ԧ�����aX�i�N�FCJMSw@�)֮�H&%�5W�\�D�qlī2MJ	gU�ACN	$BI\}��O��J�m�2mN<���]b/��!�悙�#��4��BV>O���B�T�n.�I#")��+n��T_*B�L	����&\=��. �c�Ly��
��5fH��!U�px͕�O��dj# d�'����s���Q�-?�Ur��ɾ���O<��x;$���nP�7��M��ӜdP��F�5���
剕��P'g��1�~\�
�R�Z���YdF���&T�x�T��.��}��A���&�A��G�DN��b0�^mr��a��p� $Ȯ��A��!���>� �F���{EN��+`���˝'���Ez"Nxv��J��5̜Ѐ5nL�I������ه����)��kon1B.T7bx�P`�*=�tp�v�"�DYC�A�������Ƶijb$y�NU�p�ɢ�tD�P)	Ac"���.x�7mT*:�s��0���q�ΰ@"T�Ba�=��d��Y�_�4c4b^�D�2$
R5*n�s3o�J�V�����@�0}�2�<1����4-[�V�F|�K!�ҍ� KS��6јpc��\��<�.�	�0yi��
5,щ�ˋ!�ܥ�ЫR�"Š�OW��UT9kzI�`�={�@)��f��X�T����TX��J`��$���W���$��vp�t:pHD(��m`0�� ]�Py''ˤ�^��2�݇ ��V�)[���b�A�u��+7A�cR]Q�� ��9#�.ѧ!k�#=I�- �5����`��⊹"�(���~RcS
<���sR�ׅ`0bA�p`W
m:&���i��!�h}H��W�t�����:���K�W�a3jU� ��y�#c"��(��*f�6`��(�%�MkT����3ulJZ ��D����MKw�ݰz��U� ��#5��a�4%�J�qp�B�<�=Z��C��(�kR�Ԛ�$��A�ܡa,4�k��$�L�>���u\,!�(�!w|�,Z�Y�%"�Tz祂�b�lb�'	�$Δ;��m�u�;a�~<*W!"Ê#�bͥAՀD�w`J'U�T���T�4� #4�H���d��j��1�֤11G��(���;�riZ��D��[�@{���_�>����Œ�Q�1$mЭЕ�ۦ}R� 35O�k�	fe^�!�E� K�djc�hO �$"�wi�V(���ܐ33f�C!��ٱ�Bi����`�ӑO�n�{']�2<�����:᤮F���{#F �\5[���g��''�ɺf��7�:�gM�,ZiN�ڞ'��tQ#S�r��؊�f�l&�V�T,iU���]�܈��'׮�9a�M�p�h�	�H�VIH��i&���F.]�7Dj��	a�\��$M�:�AӷcC�dw��IA;,��\�#�':2�r6�	)��b)�8 ��';@��(� ]�Ln��)���%v�A�b�ؠF�,d2fJ�*N�&�@r�'�REp��]�/�ԍ8�吅zu�h$�ÂK}�y�bn\	Z
���E� ���܆*�Ʃx�xv�@T�B Np�M�®�']�LY��@K��2�V�Z�#!��F�_�|���٠`Z\��%`��qxp	�/�*,ז"��;Z�E1�gW�C�l���-��fPL�� ��r�'m�,�wa�t���&#+
��Ó
�Z����ɷ��p��P��?�r��Q�V��P
I9<�(	e�6-e%P,�9����C	T�t�B���E�N�(�	]6g���7�I�ID�l�|S�.͑8�0�P�(��?��4c*С	�S�o�c5��T�H�O�>5�hd�J�9@\�05�Oj�"���%�
A��f�3(�42��׮f��,h�O�E���Ѹ�x!;& �P���P#�B
���u
�X���.*4�#S	/�
|�ד��X�󫄻��%��%l،�ȉ���TWV�2�g��oҘ�'HH%�܌3��|�H
@�̊x��`Zp�L�5TP�*�ONy�e��Z�K�&٢�HG�x��ͲD0
t!�.�(�F���b�v��8cT� 묐��
T�xyB��� w��R�,@;C��`5h�%1��5���)��CQ�ˋ��O��PA�@�#k��0�%
,@�����I�� �fH�`_��"�/�>��@qN�� ��eW"y�t�1��vlp @B&T�J�kBB�b�<�W!F`&�����F$�@�~%JUXã�s���s1��1i	�̸�b�>��p(�A;�O�(����;\y�XG6�b9i�o';a�r�A�y���9�|�4I��Hڕf�ˤ'O�z���!���F�1CF 
�(��#C�K�����#%H����˕(-"p��"b�P	ě}n�IA�,D4!;ɨ�(P$�&+�� t���M�1Ǚ�	�Ա�%���~u��<�}���	IP 8)��kW5{�F�y�Р7@�|�d��%�h�ڇ�y���'q�dӅĂM�����R���@`�V5[G2��P�3] ��Re��dE��dBJ?1�שu�| �׫�$���N09:�k�E�,]@��"�8��?�TΉ�GR�`)Q�9?�`� �,��BW�I	9-�P1�	�q�I�r	K"�~�g�	oDPt�S��JX��Rdşs2���>�0�s���%��T3�! S��J��#���R��r�	þu��TpR��7-ZE���$�w
�5�((��/���*��±J}��1#�1}�"%��ϯD�:$�t�ޝ0�2˧��,���z)�2Lv��F�D��YP�O\�G��d2��_��~��)_6���R��'7!�	+Q��A��u0s�B��Hb��3�~��W*G�n�!t�Y�+\�P`&�Bq�h�2TA!�y��%bz:)��(�hO
���gS����Ab!�,�N�iv�U-q,�; ���%xĨ�Ea�F�������ʻp��{��ܺ#s��j<<�Cą��2�*7������c�'e��C=��`Qv�՚K�� �	
�ʍ*�jaFk��xK�TŪ��G�����h�O䀓�
�P��
D��+�lU	F��;}B�HCE���C���/��!�Y� ��i�����xaT�a�>��a�6��e$ �)J	FMR��!Б��$'04e���fJN7(�B��`£�O`6$Uv�µ[��N�%6:y��l��dNH8G(�:G��扥'�\	AAK�:��x8��ۍq��hri��Z���KI`[��g�̤%�Vi�;�M���5㪑���sq1�ɺw��� n�.(�
���'�����4�v�R"��6Cp$Q�o(ғ@z�@U�W,��$b���=P(�qV��Qj��g���G(��0C�)�r�k�Q�u��b��3e2v���8t�~��P�� p��qj���w`h��I��HO�I�!oQ:S� 	t�N�3�©Kd�C04��q���pL��b��DW6+�(�%����(7~$�@{t�03��$!��X�rD��bζA\.$/A7J�.�ѥ_ F�$k5Dr��?E�4f�ɹbJ��^�:6��=H� Q�ڟx����i΀�	��E\�JB�./�����̈�� Ta�/"��͢��*lÚ�QP��GV�
Ҭ��<��f��dS"=�#��*D��)vIE,(c�<+�%?��*��d�NV�?Mb2���P�TY�L�
^Y$b4��ct	+_�@��잷)��s�<B���* ��M��Yۂ� 83��G{"��
%� �p�'9���0&��N��P�.��]���;g����O�#��i��$?��D&�N��Q0.����c�0")긑Ѯ��P�ӢH�9:ў� `LH>dr��� � (Πz�X��h�'�gS2й�f����}��Kȥz�ycv�Ia�
hX�Y��h�W�6fQ0ԡ���#��M���;v��0��,L|�Y�f]���Y�$�3(L�+A(��'������.9����:7&��3A����l���� e;n�9A�S8=d�j��L>R���3,������p��� d9剛v[��zG�D�Hԉ��dH�)7��.t�DH���şM��I� �[�T�Z#�d*� ϲ'ڼo6Qx �vj�r_
�W�_�.`>d��B�c���hwE |�����',�R��(�"�	pmR�HL���MҫV���Ҝ�.U�D��Ms�� �?�s Z�)���S�G$T�(��M��b��q�&�X�=�l �í"LO�|6��X3
��f��o8��D�%4v�����1<�"�Ig�CKT<LJSg���i4Iϻ�?���Қ��	�u6�b�6��� S8]�:�r��Q�iV8�=a���(HR��L4����AV�g��X���M�|��c�H(P��[��
����qy�/E*��h�W`��'�Q��BV/AYS��r���sRΙ�9-d�@P�Tn!1��{�ӵUl!)/O�m���*�<1�M�[�5а�O��@���!�0>!�a&[�L�k��2r��D(Х�oܓHk&�B�7Ob�Xe$�5a��t�C�_m�	y�"O���T�W�T���ݑyZ�IA�"O��q�̕�3��t��U(!��"O���Iͽ#EXɺ�)�P%L�I"O,���9 �&L0g$b����"O�̪ ��59M�P ���kl��	P"O$h��a��	����ަ:D��Jv"O�aJ��@�gL��x���h9^���"OF��֦IX��A���3I�J�"O�;�GL)
�B-�G�3Cd�ș�"O ��i#6��Q�;i�Xd#@"O�Չ�eB5R�V�Ѐ�":���!�"Om�7�"Fd�h��C��P1 ͈�"O�E��+Zk�h�s��S�1�"O�`!�.] �����K�H�(���"O���nM-N�^�� $�w��}1�"O:I!�^�ִɔ��+6�Qp�"OҸY��N2�p)b���joa��"Ov�{ E�W�L�k�0`�=�t"O�M�3�N@ ŧDW��IA"O�; L(yk�!Y��K6{����"OPDy�nP�@����b�՗>�:���"O�`�7jQ NQdk�e�<db"ON����_�_��PR�R*]ϔ�8�"O�	�L�WJ=�6'�(1��m�W"O8Ae�~^iS��E�R��=��"O�q&+�!��\� �Ey��A�"Oд ��$i�\-*T��8a��"O�D����']�&�H�x����"O��B��:�x�,C4��Ȣ%"O�(t#�lB�Z���.-���;"O�|IVɟG����#B�Ad�k�"O^���A���`\�#��8���E"O�8��5ӄx��@�?E7L	#"O��c#�1iɤM�p/U5& ���"O�;񄋦}k^ ���I�W�͢�"OJ�	���ms��i���o���3"O� J���<�� �@|�X(:�"O�ǣ*�L�;c������"O*5z��E�J����D�l��)ZF"Od��E�*��`�擻܆X1�"OTxq�$�9���7��-�ؚ"O���36���[Co�;����"O6m��i�$f�2hH���n6RiA"O.ԣbI�6� 8SG
#$<�y�"O^mAF�_��^pq�	L(�"O�ȳ##ݝC������%-QP�`6�'�|!T	˔T?�	/z� *��܌�9<�C���@{FbR_B9P�k��$h�O@1@�G#'n��q(4�'z|� �$H�e�1��4E�\��	e�9 ���5G�X�o8H c��M��Bp���c�J���#D����'�(��?�3��T0�Spmώ�%+��f��1$lSfl^	1�lyz�Ê���Ov\��I.��膅�:O����2({�����Ћm]�����'��6k��'�:�[��]?!: ����b�l\XB�Ӹu>��3�C��#H�ԍ�qΞ@{d�i�d�U��	\9ZI�B2H���PĜ�Ѕ�%\O�Ȋ!��Hu�=sD$
(�4 �!k��(��h�$�\�EB��J�Jà���ٲ��Ou�5K4��)�:�1+H�)��擌4("=!�%�1Ͷ��0!�%UB��?������Æ�D)�B�͊I"![!d��I���Qǚ��&����@"CP%K�v7���>u�ѲC��j�v�0�t�E!Tƌ�M=�9�BGh(���>�A ��S���	�BB�8b㦕�����F$@j�)('A&X����'o�'�Xub&� vFM�5�Έ}�Rt�XxiZt��tBI�>qu.��b0p&.¹t�8���OV9R����`Gc�*�k��ҹJ�~�cUn�h,0��C�q�6�ˤ�V�U�f Y�v��m�%H�4:��p�� �-S��ޔY�jU���,O� �l�X��X���1r�Z�a1Ã�"[:������e�=c�o> `QbX��4(0�^�v�B�i�#�'S4����e�L-����3w��Ѻg�"�F~B
I?7�����&I��[�I��`����U�V�V��U��#	�sS�œ�O;_	x)0�,ߕ9�H;��<(����� VV��I���ɵpV��ۢ�N���"�!�6:�%G�>l�yyA#�>��!�,3��	s�J�tf%�0bC�������Q#�J	sh1��B$(�bC$�Wv4���b��a����b��9�J���4]�1H�'(���=) �(5�9���90ݨ���;�2c��!WB�!���~G�dI�C+3�-�`�E�70ٸW��:���%��Jp�l�5i�)�XRa�p�V�w�6�m�q�'6����
$�Т F4/r1���`_p|8�aJ�	�j\c�֣�80��g�y�B�� �\��h��5�]��!Ȇ,t�z�^�\3`���L����E',v�2�́h�����D�Z��P	 ��:,ҕ�7��mb��ڟ� �W�C�^�ph�
�%`�������|�.�U��2��uZ�{�y�ъǶ���p/&v�Jtm�<�6 z�2��%�Q4*�p�����%���K�Y�u�B�fӆD!G],��� Ɂ�[���s��ɔcq�}�B����
���K>3�di�܅(�����$S�8h^��F��3���Bm�88���F�9"m� 0h ,�.=�#��9;oP�#�Fς6����͓>*��SƖ7ft�14L�5vhE�- ��vQ#�GGk��k3'V5<��j I7�j���q2�P-d�H���aɬl����/�&� �z�N��.�䒆�˝�f�Q��Q�c�T��R!��o������$�����*-��#v��o=� �q�Կ]�V���q�
1��!1��ꗫW�[�p5�T-c�d4�s-X �a�U��1MBR�rƉ�;ߜm b��$_�`oډY�$�P�皱	H��dw���g s�����K6���f/ړ<*�h�ܺ7}j|�ʟT��nQ;@t�e#��0�iE���H��cǟ�R��l A\�Poj�$LйEy�Q{5�̄3�91�f�6�''�8灗�`�`��ɴ*�`}��4�:��AQ�	,�Vŝ,O���ï��q  l^��녻같�`B�2\��P���N�҂Z�.��P�Hc��9�n
#)p����+�I�j�,�P[0�J�c�;d*r�"�4�Y��M�5;´kv� &.y��A7�ԘC�`<)@�
��*Qd�=�&���@l ;5E�0rl��A��1iurY��$�hqxM1�a1RQ"��Pf�9�&���,Q�7#خc� �2U�ϛl�2a��m�$:��Z��+VH���Γ��>y��CY,g�*�5�Ιh�"}i�**+J�#mL&��h@ l?Qq��je<�0��D��j)�I�����F��A��ӪI�����#,r�1���מ_-�D���F����g�0sh�����eњ� ���\2xrͱu�7fԜ�l��*���` ��8F���"hՋ4V���R+
���+�j�2,�J��~�� �"Rm�Qyt*�+�Lu���:m(�b�V-P4�����QD���{1�.26|�b�#[�E �)Č�8f<�&��(ٔu!ؤ���:�T�Ü(P����ϔ^z*���LC�I>"�-?�@T�G�̭8r�0&�@���-�Tp��J�-9D�����S����'�X�a֐`!���jye-�j≫9�,���[P�6<�e,)H.�꣭��<�Dk)=�.|irÛ4H��0	� M�С���Õ"?�i�D�����+�+;�:X)c[4H��8@!M!vI��q��A�A[�	�4MW�nx�	�v��J��H�`Ua�fW#sB��WJ��DS���~��.K8#z�CR�4)�ҋ��y���<"%P0�QҦhu/}�Ƀ����  �q�]R�]�`�,ݩ�Xv�� �O�-J��3v�+nH��ދ!�r���̰|��%V�|'���kR�E���Ħ��I��P��H�B�HH���:c����N���D�@� t<m�CF K��'v:y����M��=KFF�Ih]���VSÉ[�al�Y�'T�(M���04��=s�Ghez嫒��M+�f��`�N�瓭x��I�� ':��eĮ(~4ɒ�)�$.*x$�§`H�a��h)0b�._^P��b^GEF��E�G%OBA!�G��s\��ht��@�'DTmy�G�qX��P4D[qv@ʠ�T�"y�,��DA��SU���3���s l��<!cA�{1:U`s�J��n��G�@1BI��2����<Q�� ���@I?�:��mJ�V�x��w�9�h�!jÞ*Ҷe�F?z�����'�\�� �j7���u�li%o-u�MSu�J@D�a��IW�<�
!'��TD��H�A�?���,�}#��Ԙ �
���H�CC'��<���K��Uq�e>�I�~(�G�I�@����/0��@хh�d iRk]�)�l�aHΔ\�����Q&��m�R�G���x�EH	�f q!�ݤ(��ŕmV�,x�)I��	�=ڑ�h���:O��\/�L2���
�(���+���xu��@�.c����船'u,����	 *ѓ���,]���#��Szq �?*i��������K�Z Bӏ޻6�� "tN�<a!H��{�ܬ
"��9X= �éӳ���� ����#p��*�.�?B'2��� "�x=�5���d�{���D��(p2�ցY��B��D�(mC�����(�Z}��^m���*5���R�T63������{@��FP�^������>=��Z%m	�"a�!Ce�[ |L6Y�v�r��U���T0aє�!�'ht��Geļ8�PM�!�W$l1����+xRL܃۴H1������!>���Տ�}{����c��N�p$��kM�U�6�Gሌ6t��bAK��2���(p���D'v�Pb�N� |x�ԩG	Q�m�AY嫖�G���7GL{��6�ЗS�h
�o
#}{������l�]ae� B��$���/.Lm�4h��5�<4�DK��#=���"�"yJ���Ml�� �y�rmmڜb�$�&q��}�LE�Ua��qFO��%VpPrw	$j�JX�&d�>�`�$t��]��,D%Pk���GO�5�%�݆E��U��B� B��I�e�6��p�Y=n�N�� 	�"���S�8����&��0	��3BH��8�h�`�\T<�y9U�61����c�ǈ5v�� E#��W�XAS��>>�Q�XA�G�et���A�_⩠LZ�v�Q�G0�DX4//��L�2^0��T�=�M��%Dd잝W�Ǖ������u����f�ػr@vT�	�1�>��M�2p�^�˗A#J�^A�Ó�j��:�!Ÿ|2�Dn�P0,52�FZ�aR�뇁�"H�PAU�S!b��Za��x���ΐ�"<�p/_�PRh���ɇ�T�#�h���h�'�/�U�?s���sǕ?pA����#�"e_;uV�+��|��<a�4$��5���T>xU�W�N��4MS�'�lC��ɃL�@PrC̖
;ʌ��4m�� 9 �BAz���!��w8|��ꋒ�*�� �G�.~�9g��i��a�N)�,�6���P����Cp��́iNb(0�T|�)$��`;4��B��X�aq樘�dSN�Q��(=�ᙖd��!c���a8<�q"�0_�U!�H�?-�q�,�x}���Jʦ�p�_�	":���o�&�ay�R>{PD��Ş�u�0x:��L|viA�U�&Lv�ywk�%W��d`���FI�$�v�<`:�L��sne	���%#@`�1���?=�����HZ�\�a�O*{�d"=�C_z��`�MI�K�n�p���<�~�
4�<c ʘ�E!�@�D���<�h��O� ���bL�AI����mS�2�[P��D"�T#��Ͽ�yr�޼,��e9&"�=�"ɻ�Gޕ�M��Eӳ(�P����&|����FL<�Ms��5�ۤN�xUܔ�ߴH0~�cN�IYA��"$϶�×���pfĝ��	r�[I3x�>�1�P7:��
�2�Lᩗ囃�a��a�Q�^�0S*ԟ{Y���p�m�;R�L�x�
�}T��QL�6A��K�F�?q4��� ��+��0%i���D�	��5
G��D�Ή�&L�PH"C2�a@�*݋;f���d�A�W��z�#�B�Խ�#��O�Lp�4A�|t�(Իt@V�
f
ަ��roE�LF{"iݐW����ǩ�#��Ȼ7�.��a�JڻO��i��#dsX����#����a�ޚ��8R�E�1�6Ӷr;��C���F�����[��,	IvU!Ӭ�>gO��b-s�̂���0���[�dؘ#�6�o��X���¦X�yɒ+T?C�Ʋ+� ��h+dz� ��q���@��ő":yI��[�%��Hv��b�ɜ5�P��%4��%�D��O��I���\��q�K���S
%�t!Æױ&��$*'��qѰ��6���
��B�1pv���b��X�� J�t�E�ƿx�N��q��/UJDn�n}B�'z�:uĕ"O�f�R5g�>y�J��!@ǮWOL	��h8%xhAG	��c�/L��Px"�Ŝu�!��M�:X�X@�ՄL�z��[0G�4�#���CV]��Y t�-���Q���>���X!"VȊ��S<y�����GTx�̂��Ӽy��'��i����<�iWH��z��h��އX��Y�Ҙs�,���mA$��#?��A�E�L�:���_�^4�pf���clƭx$ hP4g/'�� I!j���Um�A+������
�e�� �ƂR��hC��5Au��C���m.,����'m�!������Z�M���R�5"��q��w�E��o�?4P`2U��W�H`*��'�H`��վ���A$	W?BօҠ�V�ܱ ��FX���d�+
Te�h�	�fl�Ŋ��@Љʐ��W�ܵ����Y��I5<���'��2\�2���GO� E �	2�(�Ƈ�"�N�)&�Q�Q�P�H#�?��*�=4�ڶ�W?Ef�y���8��A���,j&`��f�:�l����;j�Ґ��n���B蓋>�����a@���`�櫟1)�8����k���_��uid�D^��y���\a��4�JH�Lժu;�cK�܉96�CX��#�'O��m��o܉1�u*b�v 2M��^�L�ޥ�'�0���$a��	���.5q��:�6eB6�����b�汰��ѣ)}ax2OI��<;��x�i�sǊT��#�Kޤ*�� ȱn~61ʢ���Y�#�;�z *��0u�j��ԥ�<�ͩc��<y�$ �;#���7�Pܰ5�SgMذ#�i��:��`�BPZR�Ȃ{P��O]##*�I#��E'#�ҍдK��&�G5�����B,�e�d�	eht��ш
(��
Ób� �Wˁ-��<@b$΁<�(II���#yܠ$�"�ɀ I� �shҕf���'I!G��F��+� ж)���3��?S��i��]T�`��k��'�H���;tth\q��J�8��1��Va,d���c�R��aj.~=A��O�D��V�HI�뉲=1����L���He��]�V�A@B",X��Ŏ�n��E$����K�m��Y��> (r`�T+[���v[�L�;���>z��iF�V.QʨE�"D�\�Cg`�l��e�(V^�P`2d�48w�R�i�|A����+.A�� yե�\s�S0�i|� �F��TU��u�ܱ5��v�_
We][e%Zx�1�c�lw��8�F�O���N��W�@a�CM.Vm�i��Y.
�D�@U��t9��"UƟ���鲈���8	"��B"m^ 4D��p�M��<X���]-$��ZcDʈa�B�Y`��"��2*O�QA� :�<��;LN(���S?�i�#!�4՚`�t�� s\�)Dz�.���&��P�nE�\"�!��Z�N��0_�Y�0)S��_�"Ղt�u��
��M��2d���@B-�Z�P�� ��7_�0;6�^!ݒT��	
��a[��y�����u��OL��aɖ��"��a��n��q/ԙ�rmq�NӒ+�����1htp)әz�(a�Đ)@�-�ɔt�"�1Ag�� u\0�ڰozlG���1���<���U�E��	����	5&ʲ?ED�:��_L_�y��J�Pa���-G����i 
l�j̗bp����gVr^�)��&�N�i��%Srt�I7E dE�M2�nE�6xrU���HO����DZ�s�Nũ�e�
���;�*$MN�1x�)՟nW@L��Y?S��t�$��t�Zѡ��E����+�
�'KA�	 0�Wp��H��+]�hs��]�hl�9�j
T�'R�Ա�C+`��*wn�0��P	�A�uL,�;��@,ώQ��J ��9DR�^��b��-��H�a�rC0�c�A�/ΊE�j��%�<��A���0;2_�+1DЀ.,�$�>XPr�Bp�b�.Z��X=`Lr���F(���!)B?���C�9~��pb��J��X=7j����ڏ!�0�� @O�A7����W;v��P2�(���X�K$ϳ���� O+�����-ԼI�����:���2�M�G����Y`��GjfL���C�0'Z�r�o?.�b�DFZ�}/:�X�*q�8Ń�-<Ml�%�"C��hOְ��h� e��ç��,<���5.���(Jпy�.ݪ�jMY� ]�!h�#b��gN���5���8ꤠrX��tØ.)���`1$M����%�u4�p6��2?L(I�@��e)r�9D&��'Ni��댜}&H����G@e��� TX����7"��[p�1t&ڨ'	@}����}%B��E��Fn�D�B�Ҥk��<K0�Ԇ��S�x� (&`�b��,]Dy���b4���t�b�"��M�f�D,����k�2'��$Q�
݄itT�b���P%SIO�!��e�ƧE�/����+�<���@�P�@Qp�O�<s����(<�K��T�$��c���3�ޔ���,4�Ǡ��}��ɯ6��0oZ&�a�aǍ�aM�y`� 0V"6a" ���~�8ZV�T$k5�'���3�A+v�B�i4'TƩ���ɿ9*�N�Id�&Rڕ��4t*$X��2�hi�d* �2^5�'��A)l�h1G�	S����_�t���@(�jX���ʎ;��z�(�t)�C�R�����T��9��>��	���r��@��ɟ�P��ؒ-H�u`ɱ����C�9|1���^�y�vj�H�����_�!�ɥ�ֈ�C�&��E�7K�WQz`X�)Mq>�|��ɦ5c���1��<}S�O��c��2mw�BG
ʮ$]\����;'^�(�f'[�u���R�ծ��O���Z��<!AK��:v(1r._�<�6*�U?�S�q����Y�64�U���:s�{!��.BqO�� �.׀�0<�7H�7	���P ���
�
52��C��BT��p�i=]�f}���P��C�ɋe��s�jN+w��S�A)i6�C䉔o��!�	��K���p ��0e�B�I�N�6d�'�٪��������zC��x�ȰI�,Ǚd��e 1+�%x�8C�I�G&���E�G� )P��%��B�ɵP�T$z ���%	�8� �9n�B�ɛ.�V�D��P`�p��OSF�B䉦U/�`��`5^��X<,Y�"OЁQ
Ѧb�6�bFF�+Gi��"O.t9rm - Q�$V�ORв�"Oq��@�5��L�΁1��c�"OF��#��A�Չ�\Al��"O���bD/~��H�*>HFP�C"O�0��č<Č���(�:�� p"O��i3w��,��͝�w[�ti�"Op#�$K(���iW,I�B.���1"O���,��jR�aJ��ݫV�~\�w"O���m� �D(�+I�&� �#"O�D�BN/�t�)�I�)X�5��"O�p�b)�s�=����A��@�"O�\aM�0b���OXl8��"O��Pi���Ǻs5��!w��I�<I@)�1/\���I�d���'s��H�ca��M&��B�+FgRD	4�Ɩ1�HpÀ�6O�1@��Z�l+�]�� )$\�sv��t� T��J�>�p�IQⅼg��nWjX-�ᓁ^X�uS� �1H~��nE' C���E�5�6�x
çf������b��E1���!k��`fHp�O�����O�f��1�#�(R�S�aW�A{�I6�\'`¬���O���t��'$Y��٘hҝ(M<��#�3�MC�y���M�R��"���#U:�x�HS����V)Ud6�#�)�'{\�y�c�=uϺaz؁z��mZ�oz.]�=���i>� ���	k��5����x��$������'	mzӥ�7-P��RJɟjM��K��]\qO�%��MK>�����\�>�	3X�7�H��0�'�D
00n,�h�{�����'7��Ec��GL=�ë\��#�.<��{��)ї*�ڥcg��:�Z#$��F�;t��=%>q��X�x�;⸘��I�%���Q��ɤ>���y� ��?Q��>%ŭ?���iݪ>&��u��eb��!r΄$AYԩ�c"����Ls'&��>t�He��N�FJ݊��
�6�K��Or1b@�>�.T@��O�>���ưI��<��9x	��Q�sӺ�&i4��*�'2���� �p?aOҐ{��ͣ��߱p�	�B���&�&	��O��*+��s?%>�3��d�	5�\�!!
\�OQ���.]��T�p�Ŝ����it��S�.���)�bȨy�0ՊƦ��#}|��J<���F���|�M~zb'�QT�老j��s��Y���FR�$��-�>���3���A*$F:���g�p��չn�}�4BD103�����S�O�8=��R$/��ɍ�q��,�b���J`*A�" ,��s�"}R�@�%<[J��T!�1\.�E;�L�Ѧ���G+��y��)P�(�;��1hF�	*�~	�A��'P5r�V/^^B�43�!�b�ه0x.I���
�$B�I �J���"^���'�_�B�ɛ"r܉#JN�N48�nɽ$l�B�I K@����ɮA��p���0K>!�D�<p��za�	�P����4t3!��3i�A�$��z���a�
��y�!���.z��ʣ��z��	�h�0I�!�d�6]Ǽ5Ѳ��$�(|�'��
�!��Z

1L��̦wa6����!����f%�bL	�M��6�@�6�!�D!Aꂜ�A��5(.D�UFn}!��%c�`fȓ?G��$�&�	w!�dXNQZ(�?nwN�3�dН,e!򤛂��\�`�gN��qdь9@���K�}WV����4u��Mz�T��yBi���aP�іfA�8Y�%��y"�W�7��Ah%�֭^s��Q���y�Oӝ,k�Q�A-�:W�l��Яˣ�yBj�<@1(�0�8��Œ��E��y�)L�FC�@	��٘�2����yb%_34�H���#v���B��҂�y"Ǔ�l�d)sA��-vH���y"��;-@|��w$]��=�� ���y"l��ɑ�E�1N�*�����y"�
�r��GD)8�H��4���yrBͮo�!C�BC�2���P��F�yb*��a�ZX�a������q���y�*.2�9�%��#p���eg���yҮ;P����č�
��Z��5�ye�wN�P�A&n��,p� ��y"G�=4��YR��:��"�L+�y�H�3mt�U)� �b}��ȕ�yr�� 8 �Ya��H6���/�y���-��E��NW�J1BM#P�C��13�(��Ա)`��ӅIu�C�ɥZy[�^�����Ο4Z�C�I�,i�Xs3�#_��)��#I��C�I*��d"�Γ�[ǌ�!�^&��C�ɴ?���B�
*E�.�c�-�vC�I�#�n�I6/ף&���F��lC�I�qB�I͝����*b�C�	�B��U�c,G�B�|a1�D]��C�I3���å)a���re�M�a��C䉇I|�+1�ڭ4�ft�T�W���C�	�d��Q҈f\��2�B7I�PC�i�h*�3� IS��	�v@�'qn��]�)�����b��y���@��� n�tN�Qgh�s�&C�?٬I��"O�<�GjtLj6�Jp�2��"Of��'k�Q%ڵ+��9	t��G"O��������Xm����c"O\����F#�:`�v�˧f� ��"O�Dyg��%S�HP	�-A�z�`�õ"O�I��7KG<m���9]ʘ��"OQ	G@��O�tU�̻6Kȼ��"O���5�Շs��k,��{;:,�F"OƬ��!�E���{�ҏZ�b�{�"O8�{a�[;JD��d�D�r֕:"O��ʓ�zl�����)^H s�"On1JTl��d�����>�����"O�BF��
�j��#�=s8��2"Op|�g��+e�$BC�0��%�P!�$��iJ޸b��#b4�!�ߘa��D �g��Bp0�B�N!򄕦 �|��U���D��['ٍ/ !��||0-x1�2�����G�)�!���TM(�@#��@,(�;�D	+z�!���sVt��M*KB��!�֏]�!�d��Y���)�\��@��Ʒ�!�ʨ ~PSg�&2��`��Gh!�D�P��W�W9��3"�I�y�!�$ߠWyؼS ��Ь��ǂ��!���Nt���Soؔ`<�Q�E�i !�$ )[��XR�P�nA���Aܗj"!�d�!�%)`�V<�	��A�z!�\�c���P��,(K@��6��K!��'hɜx�@�=9�\�t��k!��K�kj��3LI w ���ǽu�!�d�*ИjD�^�o��p1���9�!�d�e� ����"�-!u��U�!�q�x�C�-Y��b�2�!�Ĉ�A^ ���]!
g,�LY�!�$��A�$q� �S�QBJ� r���-�!�đ�'[�!�瀗�<���e
�!�$Z�Hw����E�c�dI��=Zp!�Ę�d�(�	-� ��33�
�b@!��&:܁G�V��.�*��K�}6!�v�V̰A�>��a&-�x�!�D� FO�E�%�nd�Z�M��!�9L�F%Y���1fr���O�!��O�<�4ȱe�H��l�"b��(�!�D��@Tz�91
M'k⑪r���b�!���d����G��O8�`�q��� �!�$�5�ॲ�-B=�`�>!�dGr�ځ�(�qq� �@�B�!��J�x�4ؠ3�6TZi;�HO�!�DK�A�|���I�#?B��D�N2h�!�G}�2�s	."ȡ��D�]�!򤕙w��2���n�@�`��<Z�!�D�6k����QT�<%���7�!�d��t؆ s���8r˜�H�Ǟ,�!����TA�A�P�ԁ���\w!���LƂwIۉt��eV��
^!��=Ot-���0��3s0Y!�ƎV����]4c�TU��

(Y!�"uލ� =�>ظB���E�!��!v�U��[�t��Ύ.z!�ަ���n�]���e�
�'q!�(L�\���t�ؐ�7dK�`!���d����Z(\τ���BXkM!��+9�z���"�	K���AB�4�!�� ��E�Ǘ;$.���˚C��Ж"O�ЊL�w�\��(ג�aS"O�� �:�����ϻD�0�g"O�k��X�>���s�����%�f"O�`�A_r��b��*�D(�3"O�a�#T1��m���^)n:��"O�� ��цo@�U��U�e4E�7"O��J�!�&6R��q&]�(8�e�"OlYI�őʬ�(ԥ�t6hZ�"O[�J��Pd;)��0"O��0�`��Hm�tks�����s`"O H^�� � �P6Ԁ�"O���&�U��H��A�`��1"Or��+	�7�\����ˉ5f��P�"O����S�D Ƚ٠Ĵ�LA"O�Ā�E��C!�	��dÒ\"O�U[b�F�h����Wm�D@XB"O�X T��k2X���9{���t"O��`7��b��x�b+��0�|�a7"Oh$��$�vx��s��d�& �D"Oz�)��Oc�H�C�Z0<��t�E"O\����M�P���l��p�B]Z�"O�q�"H,I8���t%��*j�-P"O��R�(0L4J��� �'Xb�g"O�`Hb��,�*�ңT�6��X�"O�\�Vֽ.7D\�@Ӥ7ҼQ��"O�tQf��-@i@�p[@"O� ��L�����I�?r�q"O�rd��*ԓ �ȆO|���"O��;G�N6ABv���H8A�)�7"OP�b�J�'�P���3ܠ��w"O�l+��-u�f|"���,���"O���cλA}�xhDS W�f�"O��
�C�܀ �W��/��m��"OR�P���1��tC�P�^�d Ѥ"ON�9��N�<�ck� ���{a"OZ�Sg(�N_�(:v жT�F��"Ot `�&�:_#�`�0�֕^�@��3"OD�� 臽h�:4su֦ƺ���"O�l�ע^��/Ѝe�4���"Oh=�b�A B���`�Ι\���Bg"O=�eF��`���1~�8�!"O���n�%F/f�+��>�Q�@"O�=KCC=��	���S����"O���G.�f�;��@"�:�"O�%��P�Y��<���M1=��Y�"O���� ?+��Mх��e��}��"O�L��Տ �]�SI��gtp���"O^uڠō�N��Y5���8��g"O��W��H�H��*R4MX"O�|iv腲 C�`sQ�6=5 �zF"OD)B�KC h�fp;�D��y�"O��+ȼ�0�)#�P�s�<�Q2"O���Wn�>-����a��
����"O�J��U�m�*p��ޚ�I"O�Y�(�{d�B=ldj3"OF\�B��W׎0U* %����"OF��eO#TE���qCQ�k�(c`"OȘ`B�V:HFJ�I�a_5Bh���"O����3'l�� Ɣ�c �:1"O:���삾�$���ɾd�h�"OB-k4�P�t���X�� ���Y7G!��		��ړ�ŬKߜ}����+!��$Ku���(<Rs�1��\��S�? �	��54�X����/�0���"O�U�0�0%���r�B�:d���P"O����:,94!�v���B	�4Ғ"O�!���y*$"#	�=N���"OV���e����Ȥ��(<&�9�"O���%� -ra�5�Q&L� ;.`[u"O��(F�ĉr(� ҇$-�xJq"O>������b�Ղ��x����"Op��1kA��$%rQ��܅8S"O:�gmP�W~�J���
���r�"O�̐�IM,iF�X����"O���؈p��"2��6	����"OyRA9w2��ƈ�KX��P"O�e�SF�
��`'�8I���"O6}x��݉\�e8�^�6HⰡ1"O�Ivo�:1��r#��"[�l �"O�)��d��T�����gdT��"O�s���UB��)��>tN���"O��Q�A%e:��J��V3D3d	��"O�|Re�D�pq�C�M�k#��R�"O�)z�ƛ9(.�eN0��c�"ODH@P   ��     �  �  S   �+  �7  �B  N  ;Y  �a  Cm  �x    g�  ֋  �  [�  ��  ڤ  �  ^�  ��  �  $�  e�  ��  ��  .�  ��  ��  [�  ��  = � :" �1 (< CC �I �O �Q  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��e��G\���,0DB�1U7x�ȓfN����ģ���"'	(|�<�ȓ5z8uBFF�9!0\�4�C)?<�ȓJ&���GF�Mܔ��D-��ȓr���e V���)�I�_�zy��IJ�'\��ؓ�
CYP}��mɸ�x�'%��`�/5Z�}37�͂u���I<ى����VBYQg�����ر�̅�s�!�D�_b�	PT�Ժ�Bh��O��v��O�����O�S5i2p�$> ����H�Gn.C��u�P*5�Y/������(�7-.�S��M[�hQt�Lia�Ā!%���%%�V�<aWn�E�z��uK�(J����(WQ}����ɰ>��IoǨAe�e�v�Y������ RrG�G�0q� BC2b>X\�"O��#N��Of�� �@P�n4�
F�'�ў"~�A[�W�~��14dҥX�f���ybL�2|<����]c����m����dw?y����$�	z��(�;~،�R�����<��m�l1-OH�R��L�=����]m�yK��)D��  =�d̊���\?j�2vBi����S��M�Ҍ�pۂ�AwI���h�:���G�<q����;�T|� �%,G�ҕ@S���o�M�d�>i�y*���b��\h\0�D�/y�x��KO��y�l@�p���+��{䫏���'A��'�d=��"�9q�LA1A�FknT���d2�S��ȟ�;�`$)����.�<1T�����'Aў��
�c�����;\�y�$�i%ў�}*%�G�,��Y��t��-L1�pC�ɕ(�Q�Wf�,2q �kS�O1:C.���(ʓY���8V+��~Dv�W�F�` �ȓLe����!<��Q�'W���|�O��=����Ӽj�,�q��d�z�P�C�Q�<��(ɚ�Tx�"�H<0��b�Kܓtʣ=�����'!��H�T NZ�D�����|B�)�S1%� �8��	W����/��4�"=��E`>� �A�=^�����	MOt�Fy��;OhE��i�N�`�d�w8����V}H<3bA0Y
@��1h�!�*��l�s�<�O� 8v�IP�ߌI8��MY{�<�!�K�����쉅P�@�u-�v�<9dځQ��A���ز��}�<i�K��
� ������c���� v�<�Q��<3�9EH��N�*�F\�<1��S�|�"I0���⢔{��Z�<���7�V�rV���w�|}�զ�S����<iw���Y��
s%��Y�r�����S�<	1�F�T�rq�N��
e�.2��B�4B�ظ;�e���Du�� ߝ*\ZB�?A���"��2a�x�ݷ/�>B�(�^Ig^��:H
� ,-�B�I�Yf�̘�����a���ߐw.�B䉍2��9Ç悸+T6٩�&
�1��B�ɂa4A�S�U�[F��q'�R��C�I����S��%eȄX2B�	 {�	��Ɣ�'>�B%'(�0B�	�5��q���+HL����"B䉚k?��S�#Z��$�F� O��C��۲����}�C�k]�C䉘9�r�Z��N5e� �7�
�:�C�	�vRvd������ �c�+M���d��lnZ�i�B�*U;p��a��,G����&D��E�8�j�٠�T�j��,i�&��*,h�'�>�p'+B91XN��#��8X�:D�ё��A�dȉ���I�  ��6��������u)Ģ!v.t	� �..3����"Ol�3�AW�(̮�� �ظwV��a�O�7m>��?A�?qw�ח:����Bi�"+vx�g�{�<Q ���EIt[�ߠo������O�o�<�|���?#�<���
��%�6f�Kx�,�<��^���1�]$(N���� �<�ϓT�����XX7�]�4�<!�|GR�2"L�*�ɞ�<�Dm� ��c��B�I	A�p�K�EI\�l�'�Z�U����z؟Tڶ��.�N1PK4.��S�)�O��7,V�3�a�eʔ<��K	_V><$����	 n(��3�E�`��r��<��#<��韮�	�F˸=�?ݎ��e�G�C�)� �yB�(ֈ}�Ɂ
�l�r����X�E*Q��D��;~�p)�G��l�ڀ{��	����ȓzb�1`��=�%Sw)�!M=��p���Ĉey�}���@�?N<x��gٖ�!�-��T�}�(����E�-��Dr�����R�K�H���R��T����?�y�kµ&T�|��ω�r 8u�+0�ybv�R1dl��88��DI���?��'ᾜS��E���R*^�D�S�'!t���M#N�ܼ���ߧg��n���
�HĖ��I8G�
�8�@+:D�����pD��,?p����RI7D���7'��%x�4�E�^�D�7<O����$��ҩ*�)ۊ`-�BC+�4�!�D�d0y�a(�"�p�C�B�ў܅ᓰn�f���X�ƕ1��W%-W�B�	�1t�H�tʐ^\X �W����	^�'��<��JM�d���`�M�<p��TPHS�<Iǉ��s��H�e�9	FP0`$숏t��#rQ���=ц#�"� �W�����;�	�m�ў"~�!oN>w0��*`�߂�$8���y�*B�IfI��C�BՌv�"H($���'ԣ<Y�OZ$FxBF�N���Q���/o.E8aT	�y'�x�碑/Ԅ��'��sq:B�;'h,�8��_���B��4}����Dۥ%t�O<qj�)J�FZ ���i
#��@j�����hi�c�����	?K��t0��J �0��F)�+bh��dk�R�ߴ�M30n8m�>թ4!�\��G Og�<!�͐�IXh���5s��!Cc�<�W��nE��f+O2[�l�Ck]�<i�Ӿ(8�XQ�P-gɚpQiRS�<I�j�huP�"�(	���p�M�<��,^`�|��g#S�1]�%y%n[K�<ɕ �~�
�G�Zܘd	KC�<���F�T�=��#݊ �Ʃ �iEA�<Ѧ��!'`�a���^}�)"�U�<ѤE� -"&�nK�vU��6i_G�<���H.v�z�oj�t��GO�<aS`S�-��I��nF����K�<���. A4�s��7y�̬Ȑ(_K�<ٕd��"���{��\�=ːy�@��[�<1C�G^���:d���{�li�C!�\�<A`��L��� ])㍻�Ȯ�y��X3*f��aH�W| 5���y�KF�	*PA5jJNu�C!�y�-�הA�dhǠ����R���yB�S䠌�i%L�����yri��P]����cY ����M#�y�4V���xWC�tV�&�P�y�T���(x�X�K�eaiW�yBO��^� ��G�N0��pÍ_'�y"�nh(�CVFL�Bl��:�٤�y�+W �bĉ� A��p�B�J}�<9�J)s�DZ��ٚ^�"�5`u�<��k�e~�X��W,X��ٛ��E�<�s�M�}a�Y�ć^%a�����L�<! ��B^9J����Z �M;�Or�<IpNԓ7҆�5�7"X����o_W�<ق��-W�u ��5Z 
t��R�<�6�6�~tp@ �16T�a"�y�<�t@ܰ���	3-�.$�	�Sr�<��C�- 8x�펪���!�S�<�gn�"g����F)!�h�*� JO�<�A�T-tN�m��n;-�^q
!�F�<� �u8'���,u!�ƺG�Rт�"O�H��F-L�vԺ�m<Dk�(s"O�=��r��C�,�@<��{�"O �����]cTL�W7��b�"O��R��8Y����2+P� V躢�'��'��'��'���'}��'a��{t��$����rn_hȺU���'~��'��'hr�'���'���'V���n���4H��K�LaЁ�0�'���'���'nr�'���',��'���y�#צ����[=Fr�'?�'!"�'���'���'3�*A)��P���P�>h�#c�Р2���'�2�'Wb�'���'{R�'���l I����U]�D�B*F�C��'���'���'�b�'�"�'N���"a�h�����(A��MO�n*��'�B�'���'���'$��'�2M��.��А��4ItL�Al��'$B�'���'6�'/��'1҇\] K��4��0jr���y��'�r�'�b�'J��'�b�'^2�ۚv=sKH�dE��؁��'���'ob���l�֟x���ɦ;�I��BX��� ��2��I����	ΟL�	ߟ���Ο��	�����82/|�����-?s�UG�64s�'���'tB�'�r�'e��'y�R�t-� ���nx����
.��'mR�'�'���'�z7�O��d�>'��8a� �0k����$�� ��'��[�b>�'��6-M'I~6��F�N�
ִ�
��
�ppBǗ��[ݴ�?�I>QfZ����4udBq⌧S�|�Z7m�'t���R��i=2&D(�m�O.�8�<Z��USJ?�#����	�bU>*��(9�	ҟ��'7�>ͫt��[.�m��	4K!�\�0�W,�M#t�Jr���O��6=�����!��$(cG� "0HA��PȦ=��4�yX�b>]�R�#(��I��=*�
k	}x�=9t ��y�_	gɂx�g��Cў�՟�"�n�Pƺd�D��.l"�9�s�4�'��'$7-�'?�1OL����&J���bEFز+���	!�ɸ����Hݴ�y�_����OO�\_�b�K[�hq���"?i%��gG҄��Z̧[M�d�fσ��?���@�!�\�Ҧ��/�����_���d�<��S��y�-�_<��)aA�#.�Nl��C��y�'l�L�畟,	�4�����-Q<��<) e��t�n��DZ)�y"%k� �m���$Hs�D�`�Jܣ��n���eܠGg:�B@ǿy�D`2b(E�p&,��W�j�L¤�#-�j4�'C�8h9�a�e�)R��r�*@�l\=��>Yg΄"���!�`�{�'߆.�@26aB5$r�R���Ye�H�$u?~��#��5�0;%ڌ2�0�ڐ�@�o��(�6IM� �*|PEd��ID��
�7`��0� +� [X.�i�eB�|�訣w�	��z��f��q~���E�Mp��GN����[bʆ�G �ɐ����K�l���o��+�T��\`x�R��Q�9�틵1�<(1���
�B�r/�,�x0�)-]V����<�S�N�h��nZ��X�Iҟ��S����{���j�K�4Uy[V��G*�f�'��̱Q�"�'���'���~JG-p\0�I�0�V�
��ɦ��ݟ��˟����?��'*�5��p�>s�Ȗ�!Db"�������E��Q6c�"|R�� �� �tQc��~~�a�i��'wҨN*;$�	z���'4��@<9K�t���J�gQ��Yc&t�9�<�6)Z��O�R�'Z2g���f���H��X��␽;[�6��O �+�)�O\���_��'��'�f��ҳuv��r�V(��* I�>a1ItIĽ�'&��'�"�'���S66�Z�Sg��N���գL�(�<��'7R�'8��'��'9��'��Z% 4vМ7�U0��8��n�����O����O����OD��,4Z��|����]7QV5XU��N�mZ{y�'��'��'��-����M�ǋ�,Z�yf [�*�t����V}2�'�R�'n��'(�UI��';��O������y<��GK�{��c#�i�2�|��'�BnF���O<ɑ��%,f	�ܜ�ڝŦ��I˟��'��2�2�)�OV���b�i@V|��QdT��R�9��iA��̟p���<�V"|*��a�$�]�CT
<p�!�a�`���G�&�[T0�2�i_�맫?���Y0��,r�H�3�tE:�X��ĉb��7M�O��ɯ���S�t��ēj�Йꁭ�17����L�&���l��Y��Ϧ���������?2N<ͧa��l���̇kwȹG��hv�m��i��ݓ`]�@�	ğ|�3��Ο��q�)6>�{a�ؐ�U�S���M#���?��e�� �x�OPb�'e��3&��!I#$E��#F�r�����>���?�P�Pj̓�?	��?�@N hf�X�C(lZ�3PeG�&:�F�'�\�xc!�4�\�D�Oʓhn9`���0H��Q����x�Z��P�i�2����'���'U_� y%�]C�n�q����8��!ާ��%*L<i��?Y�����O�����`��Ád��ӷ��V�6 ����O����O*��vp��0��1�c�Ltp슃��K��A2rR�l�	̟T��Qy��'1��Y!����O�ʀj�EI0l32a;���t$���(�I��'�ps&�I�$e|�=��`�$	��5��*� ^�\l���sy��'�b��$��Od�T�\Bf�� R(���Jٴ�?i���H=� &>��	�?�XX����5'�$SE���H�7� 6�<!���?���t�O���t�? J(�6��oݦ	@B�>�����i��ɫ|0��޴)_�������䗥�Hb�`Μ�7-�Ff���'H�@ߍ1��)�g�	�x[���J�	����D��R�6���5�2�mZ����՟��S<���|��R�O������R��T���f��x�I��I�?c���I�BK�i��6`�p6h�#m���9׵i��'|�8:�O���O���55u
��d/�%S@����7�!�'x��'Ȏ�s�yB�'���'z��� i8����%��$)(�hy�����?�l�&��S����ry�8[
�(�w �LyT��&�?�|7�O�����O����<��[>��i��+�H9�i�
TɮMJ�����O\�d�O����)f:v����b��-��"Zn֩��Q'����?�����D�O���Gn�?��A뒪1v�p	/��bQ��{�Bw�z���O �$(�I�ȫbFL�"�7��+#,T���E��}:`�����Iԟ���Byr�'�vP	GP>	�I7t}�d�6- p%��3~@6!�4�?A���'8@d���N~�&#^�$�Q�2ԑ8��n���L�'�� ��8��ay��O�
łU	=�t�w���;oPT��4��۟�������
c��s)Bi)��:)8�Ek�	�&��)�'QbI�.H��'�B�'��P����L:�eV�2���P� z�,��?!u. �-�<�~�tITx��aB��,i�̩b�����sf������H�	�?����D�'��X:2�Z���P�e�Ϫk} (�8Tbw�ȠD1O>��Ij�&%���V�`��xXF�� @��A�ݴ�?A��?�Vn˽��4�>���O"�	't<��D�+�n!���Fa����y���.V�D�����O����Wt b�Zg]f�CB݋7Y 7m�O�Q9��<���?����'Yf�9u���y��l���ҟ]�JQK�O���U��:j��П���SyR�'H�	���� Gn���4nf<)�H�<7������	��4�?i�'-@%8�*�>А{��:HȚ��4{����'���'��I��p��E�x�7E*v�8L�i�9�ʑ�ve�ɦ��IƟ��I}����O����"�66���rƚ,�x�P�@U����O����<��o���P+�0��J�<L��80���#0�9@ѐG&�n�͟�?�)OH�·�x��G�N���̇p_`��1�Mk����D�O��X��|���?A��z��0Q�޵R�pRE�\=2`���$�O>X��B4(1O������ ͱl�B�ǃ�:C���?�$b¼�?	��?���+O�����<;&��5]�4 �5/[�}����!�'�&c�b?�Ұ�V�d�����,���e+3�{ӂ��b�O��$�<�����4�$��V�/�A�f��1�xGF��/)�l�U�Zd@��9�)�'�?9E���	�2�#{p֠	7B%=���'T�'�@"�U�����P��R?�ţ�;�6yz��I�y�]`��"�1O��2 �R`��؟L��i?�Q���,��&�W�x�QƐЦ9�������'���'�����hɎ�#��<ɥ�M�%;�	�G�X�f7?���?�/O����mm��[թB8!������E��`"F�<���?����'���BY�A�CHiD��X�R��f*ċ����F�'�����4P�j4cV7`�\��C	EP<Q8b�Ħ��	ٟ��c��?YsgH���0oړ"�ܵ)3 �5�:Ԋ`lA�Wiꓖ?Y����O��TF�|��o�Q��8iu`����M���-D�V�'��O���ƠSi���$�xmʹH�v��O��sN��cG���M������OP�;�ż|����?���{�,����e�Rܻ3H�_��p.��'�R���i >��y����2G�ؤ�a����/JA˴_�x�I�+Q�X�I럼��şd��AyZw���ѩ�6Rm�0ʫw��O������@���4�Z�I�O~�(Cf�&/%(��D�`���� ��a�L���I�4�	�?y�����'%6ui��K$7Z<L��oʃd�K��f�*鵠T8v�1O>��	/V<�vFϭ,�%��N�b"�^ʦ����4�I:ƚ������'|B�O$e,	󸼒QC�$,@\���ģ[m�c�T��E��'�?���~B
Μ��a��Pmv��)��M��;�$"(O��D�O.��"��*+����VL֤��-�'̋6���H�Ar��C~�'UW�����s�����E�O�,aj �9���� ]y"�';��'d�O�$�4$�<Ҳ���s긹C#�Z4ZJ��g�R�	�����hy��'�\��Bڟ���GF�� r�(
�g��J*���e�i���'�R�$�OBp:�H�Rћ����B��=�@�ss�5���O����O���?�ië���O�X�oߔL	&�j"�ٯ��%(ď��i��@���?i̗֯@��%��I��E2^V�����9QJ�F`s�P�D�<Y�j���+� �D�O����� �����Y�$)���1�ʻDL��>���g�p�3e|�S���
��yP�S����jG�P8����OB)PP��OB�$�O2�����Ӻk�/WPb�ܹp�&�!�!�c}R�'M�q��������D�O���/��ԁ5��nY�{��@��27M��q�����O����O���<�'�?yWFLZ* k���,CȾ�qn��?��v�0IR��k�y�O��OR�I%� hPA,׹_�n=�v�Q� ���iob�'��'��r��i>i��ǟ��p�T�+�H "��K���?H�8����-_kV�%>Y��ş���P�����^�RԬ�0�
�T�&�mZݟ�s5��^y��'}2�'kqO��pWE� a.u��l�!4�&0K�S���4V����?A�����O$�⇉HC|`� �JH/��d 5��ʓ�?!���?)���'���a/ɿP0�T��dC���!�a/��	l��O�D�O�ʓ�?��ۍ��D +��x�ğ9Զ��G�A��MK���?9����'��B��/��sش4cp��� �
΄p ��89O&u�'=R�'r�Is"(�P���'�X�'�@�G/���N�j�����z�F��'���LS�DFTO�A� ' ��zv�Oq�fhp�iJ"U���	$iM>m�O��'L�� N���)&F͚S6�b���a$lc�`�	�K���K'�~�q ׁx:���´pHZ��
l}��'�l}���'�'���Oz�i���hA'ʀa�aB�+@��BB �>Y�Y)��2��m�S�'P4��9ǉ��HM�	�H�cZ,m�#zq&����L��ʟl�Hy�O,��|6"0k",w��;1�	16�@6M�z�9��S���p#�II!r�U�*Vd�	qÃ:�Ms���?Y�?�BE�/O��O>�d��\���os~ܐ�뇹[+�|`+*Ę'�'�O���'��'XT$�v����ݸ�&��M��f�'B-��P�H��ӟ���G�T��ӥ�\����K\@C�h}�58���OR���O�ʓ�?��B�dL�F!$���[��b�y�(O"�D�OJ�d �	� x��b�	M9����b��S�����X�Sd�I؟���gy2�'�l��4ܟ>���P)*{��A �'J�^h���i2�'iB��ORm�4*�<0���I�����]�<Du�&E�����O6���<	�b4��#-�p�dԤ0"�d2�|Ҷy��7���o����?)�"Ǥ`#�D�I�"�X5H`J�L%.-sA�ڛv�',��'/��R_�d7�O&���O���J�p�l%*	ҢsC`L�sL/x)�m�퟼�'a�(����'2�i>7�+�N}ʆH�v���@�tZ�v�'�A��{�6��O���Oh���$�3�ڇ.̻j�]��k�{@���'`�&["�|�O�'ev��)�(�|8R�3�M�x�%oZ!;Ra��4�?1���?	�'�j��?�� x�A%G�V��9��+�G`��r�i��P��'�ɧ�Ě���'��0:r�%��ub A�'y�d v�z�>���O4�D�G�To�ǟ���ğL��ǟ��<7��U��?���!o�b�|r�E�E��O&��'��i��e�4�UJ��X�� j��F:��'ҕʓ�|Ә�$�O��d�O���O~�d�5"��l�4@rQ��Q$��ɥ&���I�����ȟ��IP�ӷ�ԉ����,�1��m�;6SY����M���?1���?Q U?�' RK��e=ֽ�����b��WA��#����'6��'Ӫ4�e�'drS>�آ�V��M��
a��83��5X�̈��Ñ�p=�&�'n�'d�'�	��|ڄ�c>U���G�MvȥWæK��5�MC��
>0�
��?����?A��?��F�'��Q�# 81�%Ta0$}	�͚P�6-�O��$�OD��?����<��'�Ľz&a��t-�Ѓ �/��@��4�?���?I��6W����	ß��I�?�zf��U�|��+�Dڤ���Ò�M�����OT9�;�`���O.+>���/S���#�K6K��y�я�1�M��?!�iA�>�V�'���'����O����<n�����w�j�R��$�\�l��y�b�?�g�	8
�Y�1(Խ bU�Q� �w3�6�^�@=�n�ן���ΟL���?y�����i�<M��&K6%�(�����u�$pش	�p����?!.O�	;���O�݉��=�M�4�]�>�0���N�M���?���>2��w�i�b�'���'�Zw�b�[䄗�P�0��'�_ȅ��4��Sˮ�S�d�'��'�EP#��?��%$��2��w�v��ףs�P�m�Ɵ��I̟p�	.������CgF_xe����>g��
��t�2���T���O��������O��d�OD�sAl�Yj�����ĖM(��v���\��l�ݟD�Iǟt�ɦ��ɥ<���n��p�F�]$TV�`��-K���T �(��<i-O`��O���O����%m�,n�52��i%@��VH�����Z��k�4���O����O����<������۫O�� <*^諆�5QR�8sش�?	���?9��g�7;�@H�޴�?9�S�9��(N�-�u��+
��t�q��i���'s�]���	�AF~���0�^ޭ�#Is�(�J���^�~�m��t�I埼�I��@�4�?���?)��+>�k�N��h!Ej � �T��iL\� �Ia��S񟘖���4/�F=�c��2%�|*ʈq�L�n���I�H����4�?Q���?)�'��.��}RF��>bpD81�(�!^5�Y���"g��I�,���Ē~��K>tKD%�d�U�.�.����ߦ�����M[��?�����'�?I���?�o���x1�N� 8���A7ۛ��,'��'V����t��t�OX%9��0'o j&�]������l���'g��'RD�K�m�Z�$�Of�d�O����4��&��抙T�:T/���b�ЦE���ܩp�2�$�)����?q��'O�H�R=	犘�O������Φ	�I� vB��4�?����?a����Y?�rE��xX����cX5h@����G}r�����'K2�'���'b� � ���}.��2�
.�y�'�5����'PR�'����~z-O(��ޱ~h6)m�f =�G� +?G2��16O>˓�?����?�,O4�X�$��|rEe߆1M�s�ՃKIĐ�0�K@}2�'�"�|"�'���͉>^�o�p��H&�:��	��D���듲?���?�,O�豵G�@�*:���9 �N8U�[q�8Jڴ�?�J>y��?�'G�.�?YJ��	Q���1H /�2%4�r�DfӾ���O�˓+��hĜ�4�'+�T��H��jY~M���R�T7��O����O>�A�3��~�ǃ�n�JTY�*αs��t��Ֆ'h��QG����O#B�O��s�@��TeF<-�P���3ajLnZ�����۴���M�)�S�1	`]�4,S�{�� ��%��u�
7�
A��hn��p�	㟰�Ӥ�ē�?i +���М�ۼ�ʽ����>Zț���Q��|��)�O�j�I�xl�y��K2W��1�c�զ�������$m�b,�J<���?��'ט�� ��&u�4���%�J�bٴ��C�\���$�O<���Ok�E(�q�f"I7n�՚@�ñB�f�'q�F�3�$�O���&��ƞ]#�C��9@H}�8�@�P��-b���'B��';�_���De�`�E���7ym����2�ج�I<!���?�M>)��?B.��?In��J�b:�����d\ġ�K>���?	���dS5@|ͧ��1kA��H�u��
^���'�R�'@�'�B�'��E�'�)�4o�&gK��hU+��
��H�sı>a���?	�����-R��$>�[��(1>�,�7��.����$���M�����?�\<I����I	�|9c���!N?P�� �pӊ��O��uЛ���'$�\clre!�������kY%~���i�}B�'����f�'Pɧ�i��o�����ѹ7Rx�B��ec��]���+��M7V?��	�?�!�O�8�R��@H����M�
�P
4U��I�2~|����\E��V�K����U���۵K���M�Ao3��f�'���'�$o7�4��\B�]�!Sl��Co
C������ٟ��'��#}j��`E�P�!(J�9��
�mʆ�i��'��� J�2�'��S��l��n���Ĉ���v"�<�6���$�F��Q$>�����IVPN���'0Y�̔�2���<���4�?� !B�nY���D�'��>�tP)fr8�c])RD��qF�~}J�-��'���'�2�'k��U�8�p��I(I0vaS�˛����SQ�Д'�R�|��'��b���M2Al� ������W'wn��
b������O����O��	r�3d?�nud*ڮ�����ŀb�ژ�s]����ݟT'����ݟ@{�c�>9�� =�$w��8"���2u�SF}2�' 2�'��ɳ"wp�O|2%@0$�J���L\�#+��Ǐ\8[���'��'3��'{���}��֨���@���1� YR'�΀�Mc���?9.O��k�F�S埌�Ӭib]�2�ٔ��0�v!r4j!��O���[����'B�Y���֯K��y���.`�`opyBG��i�r7M
v�D�'��dC7?YC��3�pq4�,.^2	@�J���������S�,�S��x��4�U!%%���j	 p�m�6x�1�4�?Q���?��'F��'��/�-�x���A!�ؤ)c�PPj6͉%��"|���E�$��O��<�Tͪ�&��/+�՘дig��'p2�b�'x��D��2�Ri��"�P۬!1��Ώ����t���{�&)%>��I��	*�n%��,ҫt���C�	>MlYqٴ�?ٓ�J"`>�����'�r�>1v��b�rmg�@w��� �DG}Bυ���'mr�'8b�'%�<>�гG/��	F��R��d.����'�"�'�R�'�'�B�'�$m`�.���y�+];P�V�q��+5��O����O���<1r.R�󩋲�䱨��̅J�4���R#	�������H�����	���=\bE ���O/f�ţ	X�H�'W�'�2T�l�� Ė��'Y( �vj��h�r��)жE"=)ƶi��|B�'�B����'TV�(�C�&GX�	��I�?s��4�?�����d��`$��$>����?�(a�ټE*v��c���3%�A@�� ��ē�?���u��Fx���%2���{����&e�k́	a�i'�	O�&p �42&��������D��C� �*�!*�"bO4 �f�'DR�>�O���]���^��9��Fţ&$�@�'�i���1bLuӼ���O��$�|�&���	�j�!����� ��
���4Z��]Gx��I�O.�" cǬ+X>M��l�"�h}Ф��������d�	 }j��N<���?��'��59ŗ*\dh��k�Yre�}"nI0�'G�'����+-��m�-���0 ��v�46��O�y� �|�	˟4�	B�i���Q 3m|0���N���'a;�?���?Y,Ox�)����O�����׼u��A#�ę�Y���$�4���0%�0�O\�
��� 	��!4��J�h�$��O�D�O�ʓ`"D��5�~$�2/<�R�J�q�"�k�T���Iʟ�'��Eyb@=|&�q0��8sF�\zu�G�����O���OH���O���
�O,�$��� a0��޷i`�Y#놾rE�A�i��|�'��	�&�
O`��s D0>��2RdZ*Ka"lp�iN2�'G�I&�I"H|����Rs �(���b��պ^�Q�dkX7G����]9.S?7��#-:�,sv�Iy��XZ���6(���'���L��'^��'���P��um>�5/�:pQ�W�+�6��O��MW(eGxJ|�Aƕ�"W�3����
0v�ڦ��M{��?���b՞x��'�܍��2zE�7�:+e�Gj�P�4�)�'�?)U"�.?{��K���F�d�����T���'���'�� y��*��Od�d���ed��G*6���G�>��T��&�ɡ1}�c�����4�ɑAv�(��ͩj�R�ЁfT0Y0�xٴ�?Y�A�	i9�'5��'�ɧ5�`E�����΀�9$UI! �����/~1OB�d�ON���<i���7b�d��0�Ҷ/��єk�mr�A㡜x��'�|��'���O�/4�*�G�%)"px�D3jĸ��y��'Rr�'~� #��
�O�J0�q���2��3zDI:�U� �	̟�%��I̟xZ�+�>�� ��W����pf�:�^5i���V}�'/��'��I�x���KO|��f��{�������u�r�2�ځ &�f�'��' r�'-�젉}�J�N*�0��q$)1�M�I�nh�dɚr�n�T�8�f�9t��7bO�L!�- ^�M��m�K�bDsM�	���)S?c�9���F��y�J^YH�BL�)'�Ds�bL�u��Q���ݓ$�L�0>;JT��KTS�m�MA�8��C� C�a����Wt��	���N��)��͓|����tl���I�f ��Afj\^�Ap�C͓h\t�!o˙h��5�Š 7M��A�Mv��d�윿Rk�BgnR)ti*@�T-pHP� �HǊr���'���'c��]6D�R��%2_�&:G�S�KX�rg(\�40����\�m����	v̧[��a�g�d�lB�b�p�R�	�E
-5<٨D"='6}�XC� 1�eъI%��>)Т�>%��A�"��2���\|��,[�B_��d4?�t�Y���d�'5��`���ˆ 3ƎJ[�p{�'�p���)M���k��P-���Od)Fz�O�RS�hBtɊ�>D H� Z�M�!J\��h���Ɵ��	Ɵ$����u��'l�7���9�Bi�~�3�kŜu���#�F�Z3���t/˴U܊HXǫ��v�<�v���(O��0����6�� �凿g��t��Lo�v�!��0Vl|z�)@�l��0�eJ�&�d�H�#*��ڥ&��t���]�Z��Z�g�9p��{��'���w��m��va�0j���_? A��n�:���q�&�,�ȣ$�,�c�(3ܴ�?9(O:II�I��m��ʟ�j�'U�M�`�R��0Q��4��䟄�ɃD<�	����	�k���y@�In�	^`x!�I�;x�|�tbD,�(��ݿq�Yc�݉nH�I��1��eX�b컰K��n����aA����O��n�䟸B��{a�(��W,衢hjy��'=��|���Ə2�ᡓl��4���U� �]D!���확�2 	��2�[#,l�JgF
3�M*O
С�@:<R����O��',Y�}��/�`�K��b^S �Дt"�����?�P�Y,���(f�����S��^>��c�W�B�4�K+Wnl� f`%}RMދF�l�R��
 ��~��)��D`����)[��X��O�{��ٱS����hnΟ��2�/�&4��0��:/U8�CT_��?�ϓ.���0E�9r H­ ;G����Ó,ˑ����@�A��͒#$ǹ2�J�
�o��M����?��=�4%	'���?����?Q����K#�|����
�e� 
Q�	*$
ui�lD)��O�"�R0CK~R��x��]�:g晒��Cs�ՖRY�e���<F��S�+5>�=�噇+w��3F�xۣ<�H��Ŋ6q| [
?MV*\�7KBy���?�}��ߟ��I1��D��㘃D$�{Wo�
#<��ğ4�')������W�s�&9�p��<
Z���N??�5�iS66�7�D�����<Yqō�|6����B�	ʖ��WHK�h�����?A��?1��t7�.�OJ��u>��QV��b�
�z��p�6�@o1���4v���0��.h���gvQ�4hE�L`�P4�kޫ;�>��qg6tF� f��*p�69#�,��`3t"AV�Q��y�KZli���cg��.�� �=��d�O���#��v��Knn��6�۰U�AJ�@U�6B�=�ȓ4�l-�g����t�8!�� r��<�F�i��P�43�5�M��?yd���m�X�i�ȃ�FE�W���?Y��P�	����?Q�O��d����]Q��A������/�%JE���b6��#a�DZu�#?�rH�0<!���W%K���j�,[�@����	�h�ŀ�d�Zl#��I�o����O��`<��B�"$���1%*�4�ϓ�?��������Wȗ�I�,���׍g���h�OX	m?c����0&m��Ò`�7����Hy�I�%�6��O��d�|Z�����?��ͮp ��@�#̐!�Q$M@��?	�|���dՋ�D,�P�ʧ���*3f2���/�^F�ѱ�Ϊ2R��V�PBgE `���銝r7��b$���<n����M�DB�(2x��ɍ�M{@�i���� ��ٰ�"��M����<Q��1���O���D�.Q]���@J�	G6����Žj�ax�� ғoT<P�AL�.����)!�@V���?a���?	v��be����?����?1F��ty��pP��#�(L���@L�#�Na%�\41b�G�ӻ=�����Wk�!
e���u�Љ�Rh�.��ux��X�Q������"�|sk��>ǖ�Q�-�G��O\��R�`�ＣŅ����5&�6 �:�P��-;]���<��G��>���OH�D��7�j�b#���.p�[`��I������O�9��*�(Ѩ��gKb��H+�7O��d��"�4���|������\���pCj[=uv �J KӪsƚm�kܖt�����Ot���O�鬻�?I����D4-nl`�A��G��@Xt-/+�Zm�f�	2w�X��F�r�B$�m�.X Ey%H
~������<�u���Z!1��#7�U-@:d�s	nX����f'H����Bc���'����&�.!��zfI�	����$e_ �?������?�����'�x	p��_�'=v��K��3L�M�
���p���C}A��
��V��<9c�i��Z�$����MK���?�FCU5j�nL!v��� �"Q�1�@��?!�4Ò�i��?I�O���h0NӅ2����'�����%@!���-6�li Ǔ_|�p�)-��fJ�z�K�}�D(�a��/#Ї�.X��D��9�O������L�8�Q0�11�,�x�>O��O��"|
T�ݬG�-�q�3,�)���Vs<�i����J��)� �g���[��'*�>j�	��4�?�����	�:>� ���7X(��0O�t��u�Ȕ���OD��D��<o��� �E�14!�`��C�*ыU��|Ω��<�sbZ�W�ZШU#Hk��L(	�Ƶ��mJ�r�Īs�U��򰍜-��� &�a�= 7���R����\� f�8}BN���?i���䧮�lt�tkr'�j?����ɇ�V����<	����<�Q 1��!S��0 ��� ��&�hO�_@�'��0A�9Y����fM�`�$|#��a�*���O�����cX���Op���O��4��at!I������Fvxv b���prH��lL0N��Dt
�QY�c>�%��X!E�IfΡ�f��H��HS��7>^��`R2&i\�	��7%�lhY"TD�4-^�\j`yͻ0��P�p�K�j�v��ÃCb�
p)��i�˓ZL�i>!�r�7m���b�	65��������"��ȓF�
UJ���m��� Q��)��?-���$��O��3�l"�&F� ��$�&]�u���CF�)/�nQC��?���?Qն��$�O���5ϒ*7�Zs�8P�7�TQ�(t��@�@3*5����Ȱ=�O��g:�y&�ҩDJ�3��@�T|.E���\�V�:���/c��$c��_9�hOV}9'nL�e� ��! \4@�t��n̸.���'���'��ܟ��?I¢�xB�P��`�l(����j�<	2M�4����τm��P	Ze�	��&�'���B�8�ܴ�?����p!�"�.\*<��4ܻy&Z��?a�	S��?������3��)	O>	��ϛW!�q�âë%�Aav8��9����H2@FM��~r�	�y� ���d��Vqt�S$��p<t�͟���4S���'��(���+}��1!T:'���Z�]�x�IH�S�O*���ҀюO�͂����x�
�'�t7��N����'I1-}L�A�nN��$�<)RA��
ٛ�ϻ?R�SSZ���ɵ8*3�ަRʔR�^�fDi��ɟ,���2G���b�ޯO�%�p������|*sLR/E*��1g�.<j%����`��3�dKEEÑk V�kV.QࡃC�p^�P@��O&h�Ǎ
�P��j�����m�K�8(�.�O2po�'�H�f��K&ZR�)2u�u�H9!���y^�B�I$K��sc�*��!x��*�hE{�O"#=Y�&�:i.�*���;P�0h �_8���'N��''2Q�r*ǝ-z�'�r�'+r֝�ä��h<)0���WTx �J��u�A� d��B2�XF'�_̧��7��=�1$��FH8s��8���y`�֓+c�����Ψ����#(T��T�Xʟڑ�AT��y�IۈL'L%ɲ��-e���;���3e�7m�ky��1�?�}����If��I��D\$v7r���p���Ɠ/�`1�@�ΖUE8���b�)|���'Tt#=A���?�-O��8�N܍V6ε�0�F4	i̡�)��`!Q�C�OJ���O����ͺ3��?y�O���jr�LH�����n��=����EaM5e�3	LD�*�x�U�'��p���F�U�L1t�Q�-�:*VXB�:Y��
���>���0� ��v�|B�J)挳W�K6_�}���X�d(��měF�~�$�H����O� ;��ˣ��1}��H��0>!O>���
b�{àѤM�(�2E&�S�2M�v�'剂G����ڴ�?���E3T$���E;dE.XI���"wU�As��?a"Җ�?���Ƞ �ј��9AuJ�:f�HH�q�1Z�Da�%%��^QRh��I�s���w�`���#/�0Tș����L��d�䜴z|ؗ�'@0E����?����?�k�`|�ժ!&���.�Z��'%���3� 0yRa] ��a�1$�v0�;�O΄og�f�Z�q���nK$#���	Hy��W�;��r�'��Q>��I֟�!�� �:��Ĩ��G�ah���؟p�I�,��8I0b�hI�P��@��
 �ڟ��'�pu南*���1�
+)JѤOzE Rd҅+!Rʓ�ϛ�v��a"�-"����#�~���1L�ڵ���]� mҤ0p��J�$��
g��'��'2�BM@�眹+G.�"�߃DDY$�$�O��dN�|�Uy��;!�v��`V�&�ax�C5�[9 �ńH�Y6Τ�+Gx3dA
�C0�?a���?q�NN�-�85���?��?y���l �Bϧ t��h�HYQ2�9<l6�CG�[�`�%ӏ%�n��T�aӣ���d�5/��I9Ԋ��efQd�.X���"�s���X�@��L�ȓh�(�FՔO J�x�����S�	�;���4&�
Z$��P�6s6��op�
��	2=���Y����#hz�1i��I�E}�RUM�t^l�'M�}�F����x#"�3��x����yr8O7-E���$�T�S�?ٖ'¶XĈ�2$����r�� F,����sh
0)��'Vr�'|©v���֟��I�1%
���ߛ;l� �!لq�ر��	O|��=!�@
�-}�4ı��H�s�Q�s$��p�L�$���+���P@��o�lA�'�}'j���L2��h�UJX�I�Q�����şD� ���cX��QF���(�$�O��m�֟H�'�_��'�����}4��A��)1������]|yh$
9Q�9�����I�M>)q�iG�7-'��O��4�,�:�ߵ)ۜ�sL˛x?�Ax"Oր*zJţ�J�;R��˥"Oȼ!�
�*P�I3
֨B|�<X�"O�DP6� �g���K.r�4�"OΑ��L�V/^��
��3�"O*=(7鈸N�!��,@����(�"O��1�Q<x�@x��M&�z &"Oz�bF�j���AD��tf8�$"O���ĉ/��"� �7l`��"O��9�oC��hx�.�1w? �X"Ov�K��(�H��uHK�t�� �"O¼�DŞ�v%�(h�@T�q�����"O,X�Ӫܟf>�92���6h�i{�"O:�8&#D�h�Tp��41^��s"ODy�,Qh �"�$�;o�"OLI9�d�t7젒fC�?M���!"O� �$ꎙF�kG��J���Bs"O�ęg�J,`\>9��AU�>��Y"O`ၓ����=RF A$ko�d85"O�X����9AT)8��.*D���"O��1��p��)����4[��!�1"O�0삖�h�
��S���w"Or-�'���J��y�BX$�`�V"O@x"�n ���QeKǹ�Ƥ�A"O����"Z9�N�p��b����a"O�)@�Ztrd��W��#V��U�q"O*�h��(ψ}"�ڇn���f"Od�&[l%��]�umz4��"OFœ�ШF�zZ"υ1wl"��"OEjmq�n�s�/7O��8"O�RDG�-�p��N�0BV���"O��K�HF�����&���:�"O橂�K�5��zu!Y�\`9"Op-�e��|��@J!/^�'���$"OF��W�SV2�{�M���	:�"O�, �ݤe���Z �D�xB�`a�O&,���"P�����+�����P���5�a@X�T��%qcә�!�Od*|p��JRȍ[��<�@a�@��'G��4#щ̘ް��t�?Q�?QlW.qm�*��$#�D;�"I��p��� ;rP�@��B��\Rub�1�0Ÿ��5Jt�Y)@������	���,̫y<�b�*RK�V#>!���#A���{1��lRDHd��
�J��Sh6��&.Hk�|�w�c�<�wH	(�٠r�7E�E{T@[�<��-n�)3��J�����s@)�h��=�A���f$zB�V"W�H���*O�$��ϔS6�QࣅqE�I�R�_��M;a��@�J�S�l�6���6�)� ��VA�-3�8E�ZBZ@(�' ���D�Nú���8S�Z��A�&'f@������=�.�qѦ�\T�{I%4A6�rA��G�(�!˙��O"H��.����s�@"�d8q%�X�&��cX� �#ƅo+��Ȁ"Ot��s�]�ew.EF�6uh�ñ1O��Xr�C���"׏WX�t��w�-�'{6F)��
�G�H��"(I�^8}�gk�b<�&(�,c��̊�LZ�0�4�#R*
B�0҇ߌ(I��K��[5�2��|JK>i� �/X�x}rᏃ�l��*�.r�'j� i�(�yx|p凓�<)-ON����E%Q�PIX�R9>8*�&��
-?XU���U�(�ᇫ2�	E��Q�J���4<޶�j�h����Q�D�*H��eK�f�G|%�1ؿS��l|�p!f�1�0�"IY��'�$(��A��'됭��� � �]YQC�p�'Hb�q�l��?H��k�j��;��B,��uw5����/�T�!����<��	��oLT̻���	�h	E.�؃M
m����@I(vI���/[�<<��?a�B��<�E�[ �E{�j�<{bڱ8�Ά{�''��rÃ^?E����9v��'4� �5C�3I>N�Â*��3^RX
��>23�9���l(BY:�%��@��!7�|��O,��2X���Z�GMHѠ�X�[�c'�-��!�Q�ĕÐK�����i>�X�O];Q��ɑSF��dM"%u��u��D�<�r3�ױY?�$PVO9��Ǒ�֣?�B��Op ������;�$ ��͔�o4����xW����Or~�>ф���mV�n��7d��עFs��YS�n%<Od��ӪW%7s�xQF- ��zB5x�\ �����pXў`GC >:�@� �5p�O����3T��l�` RM��9��7wG00��V?# |xۀ�: $��	! ~���nޏ7B�L��b�k�L|bS
�O��z'�߄{���	��XTiK�8����Gy�eT�x:;���b=&�X��
+V�F䉳��'T<h�k�˨�`�'�:9�����'o�IY���(!˚�z�g	*���X񦌴u̌�O����=��Z�l�'P�m��Kw(�:� �1��<�Va]�p�2�Gz�A!0� �� ��x�GF̜��q�GVaA�G�Wx��s�OF>%��@�ON�a�0�k0g�
J(���B�$N��=��k�`��'�"Q
�̹�p�#����Ma�I��cN���F,�]����hVU��8����G�a��v ���2��I��O��u)D)���"''H�d�`�
����e�>�P'O���$Ӆ	8pE��R+�$ ®ԋ'+2\Z�H�!�Hb1�_"blJ�z�:O9rA��&�1O2@�S�"2�  &�C�N���('*�ze(! O���UFDf�'_,9���my��Ņs<�=C�͂��yᐥ9WL8q���	�����
,�Dh���V�K�}��a��\@���Z�9�@���IE�<�'
��\ ��dPI?)��>q@d��-`e�M6��; J���,�5w�(�l�C�he q��6YZ�"<�"C[�w��=�U���Ȝ��Ē><w(��	��0:p�H�O�;_B,�'Y�_�t���C�=��Q0�Y��K�C�[}�dK{�t�kc��<Z��u����W϶峓Aכv�^̡�AL�?I��Om�e�?&�T8����;A���aM�$2��7m�:gxTty#�O�L W���On�س�ؒ��ke�M$<PQT��O�,K��	�I�h�	�hp�`��xpi��.= ET�>ꀴ���S�Gơ.�p<i�O�vP}�;S\��"�ӱV1Xd�7㉮Q�f0�'m��k�y�X�͓~��"���1��,F&&��w�ᢡC��GW�vR�*���(O��xw�2Ea��A��W:���OF����q�����(�m�<�@�j?�yR7O2��$��peF��ŭ��~��	�Ɓ�!�V0��FR�B�'Õ*`����a�1`��	�'i0��7��8� ���/B�
 ;�
:�j�I�uX|P��	N��4+Wj'
��	 )߼T1���A�2C�`V
V0(y椈�'.���2�H?)
	���V�_��̢�J
�ns�u��I;5D�mZ7E8n�CW��J�8��\�@ ��Upj�����q��4��iRe����z8��ф��=��e��
	�}"'�Z5�X�A$ђ`�ᡖl�2r�扸�-�.n�Q��,
�&����BE��x���4&���4�O����:D@hfˀ$t�����$
���b5OI@#%��P*�F;h�Q��E,M�ns�1����n�TT�o�D��2
.��2AU%a}�I�Y�As�SZ�w:Rpa���<MؠҖ�ψY� ۢ+7��̅�ɨ^ٞw̴�U�]=�`aS��؛R�x��D�<��I��-��l�rO����!�^>�a&��Gt4��2K�Y�Ұ�5M6�HO��3��z�|l�-Ҍ�Xј��?��˔e���Pao�2tˮ����`�p�0�dP7S��l��V��4���4K.����OX��ũ�7(�){5(���T��i>84��%/d�䨄�J��8��L�pp� T�u�ܻ�'�[V@9�5��~��Ν���4�)�������
�ի%V:�ⴢ�",�h�{$ J�@�X�Xf�����R�x?�s��]�APj��#~L}���B�~��'�ՖUV�<�s����y"�Ŷ����9Mt\$���[06c"0c��H������D �?a7^��A�NS�����HL�O�Lu9��Q�{H�8�1�]�V�h����=ғGo��`��dߌ��e&X	�f�է� ��@�-�10��  ���9>�rI��覅nj��y�'��"K�#����~r��(֥M�.���u�:\��)��cӺ��ҭ�r<~���|mZ}T4O
0jG�V=48́WV���2/C�.�H�*2j�7��݊��>�B�G��~r#ڒ.��E}��B�Yj���?B��� �eӮ9Y��(�i��c� R&���*}� v?���Z��V�4 �\A @�>]�~x��-�.�`L���p~Y� %�#nh 8I�	ϾU��\�s&A�=
d��� ���'�z��@�c�d���@hR�HS?X�WBʴS������=K4�2 ��M�Ԩi�m�	FE�*_\��7hإ&�>H�c�.ՠ��A�O.4�y����e�i��銵��*P�Ć4�����cW���r��U��+�5U0d-�db�0�>����-�y�C�0H.��I��-���F�[�>�z5�T.y�le�恜Gz�ɋy$r����t��=�G��M�'�Zm���C9C�8=�7���y#3�Ħ<N>O�y��fAK���0�~�n�O�5�֨�Z��e��-̝E���;v�L�(�l���'XT;s�p�Y*��˹=�N�[�O���B1&��vD���K�(a��'m�c���q�<������1UΉ�\F@4;�)�'o��x��b.B��(c�Fg��ː�>���W*�Y�ʚ�a$�-���kʛFmSP�FV���O�BXq6�ԙE�0�s�f���\di�k�D�,��i�ua�˓�l�t�[ �0 �$��O?�vЈ[�1YAG����B���?�a��U�$`ʠ��	T��	�p��?#=�Q�`���P~�1��D�?x�p�U˙����O
�]�D���~y��?�g?ySN-'�p�ber�8���O�we�pF�
�p<�nB!���"Ǹ��O���D��x0�)vT���o�O��3�	���X/R-���$Ոi���SRJK��PXF��VK�X
�b�;��+��|je�ux����
I�]�����J�� ��D�+3h�����:��G7�,��i�����BB�^��a��yN���42�\Ij�C!p���$��	v�&�#�g�'����0X���GB��9S��(�'� 	�aBO�?$��7ۮR���g�'�@A������!��ME�%�^-�3�8k~m�$��K�D��Ԁ��4��\�"�xB���a�����cO�}�r�A��E/!T����]�;�џ�e�W5�q#"fY
XP�)�
Р�����^RE� ��<� �]�^5FyZw�����	("�F��n�A����Ϲ_ܤxDx�4O�Ȭh��� &:, �Eտ3?�iD���@�lZ�	�m����>5�(-�De�t����Р�4^��dQ*�0�	�%ݦF]����c�::�ܴ�R��u��?:p<Р ��^�z ؕ#�WZ���/N��뱡���T�=���ƄZ�fŬ;���u�,Q�B�s1
n����;�.��%D!�@���=_p����	f���[�&̷Z+��`��
�ڜb"`�%��}�1B���s�ϧ�h���^e�Z�I7����DP5Ǡ��qm�%".��pK.m��?�v�֕���lӏPV�%S* �:b�9n��T�TX"���	��c� ���^�Y�F��'�~Z��D�~��q��Η7w��X!&�"�d�E���et �b�+fd�F$\f��̸Sbr�H��D�#�Y�@�Еb�ʍy�.F�0�^�zb��W?K��xfɌ�LD\+�O�� 	PAJ�3����W�G�����@��.l
�Ju�F�WǨ���֟���X�<�n���u�M�<��b%I$O�\��W���'Ϝ]��G�gY�@F}��֊t�<u+R�+R���Ё�	Zh�J�C�b���J]}"�Ǩ0�,�):���8����X!F�2e� /zF�qj[-G��ui�O8��&�E�-=Xz�H�(L7 `�����p����ȑ=��	$L�D�|�ۧ��
��Sf�=��4H�=F��� 㒮b�0FxR�C"��4X`�<N����	�E��i��(Yg���hI�!��O�,a$@A���5v:����x�:���	{�� Na�0�<��Pi΁F$���CG�Nc���g��.u��eLR�t%������'!�Nu�3���b��2eE០�ЈA7��ɪu$���'ߊ$qu�;b�i��*��:Ʋ���X2�ܰ!�*��~��"��zF��۟w_B)A/���C�cvP�E��4e���Cv�L 5hv�=�1iShO"U�����mK�	zt���5 ЊoZLM�4�>Ec�Uߴ���a��դ�z�D��~�ɏE�%g��1��-�Q�
�<ѢЯU�D�!暹'	�0�%�|b ƛv|B�E)P�DmE4z��b�/A 4�P���q�D����	5TV�'_��#r��7[�����ûF-Hɇ�ڸM	�FI^�<����-{&1��˴@�U�I�L��Y��dD�tCL�x�ؒ`A���#�5D��D@����&�� �t�cM�O$q�@�>.�\��$����y34F� N�hq*�%P�!�YSZ��a�J@ ː�U-�!�d�*MN�dX"�U� ޜL��H s�!�䑋l44 z�A�"����&�Ȓv�!�DF)�lEEi��x����Z�!�ĝ{ǒ`��يF�ؽS���?!�ؗl� |�׫X�z���dc�!�D1(�R$��W��[v�K��!������'��=P�mH����z!���B�
S��d�N��Кe!�� �mj�`C�P�6���l��kЩ��"Ob����*^i&�SaA�0b�`�"O4��pd�=R���F��XKL���"O�Ț�%#6�H�b�����r"Of�	vK�I��X��ڍz\����"O��$�#��R �I�?Wѓv"OzI��+Z�U[�G�(\���"O(ɓӥ	:��Ŀ"<<��"OJDS�	C�`J��aI�Z3�"O
�J��*n�EI�`	��>��"O�ċ���&��U�0h��"O���ET�t ���K�5{6��r"OND�G-
\x����h[��y$"O^X�t(F*;؀<!��ٿ]�0�pw"OL�6�3X X|�c��f�Z�G"O}��Z�PDrA����*G"O"���gՒ^̰�H�A����6"O����$�WL��g�t�����"O,5Q 	�j(J��r珹,�@5S�"O
e�y+���!^?X�f��R�!��ֈ�,pSTク4�q���9!��׋Xp��#ѥEF��6��0!�$Y�m^���T�Y�,11⊞
!�䄰sڨ�a�	��#u��� �{U!��4��a�!+�roV$vHߍ7!�M� �&Mr򮬑QEǿ !���
&;D�XE�N���y���'.!�D�7$���b�)Os�*�Ӂ㌅"!��ϒR�D���,T�a��Y���"!�$ �H�6�j�N��f	hE	M�!!�DU(���#HƸ&8�L���< !�$3-��AR����7!�dޛ]����_7f$(��	}�!�d�4B=��av�ڤ}"p��4&��;�!��<mC��	Q�Ū=4�`�s�]�!�Ę M�.LI��S?3XXH6�=�!�Dƾ��e�O�b*G�8�!�M�i)Fؚ���#B���ĳC!�$98E��g�E*՘0�Ϳ	!��%�v��CO��!�ǌY�!�4<f�hFf���|��	�!��O6U�D5��5 LG� !�d�3�H0Ɗ
��j՘�ꕑjp!�dG�ij1c�D)t	�S��Z!�䚹\�,���GO*yB ����$
W!�4v�f1jv�*̘���T	A!�T�w=�
��9�$����"�!��� t�K�.R�M[�%*R�[8c!�$�� NN��eI�v*کٷ ���!��C0������=x�JG�ʭa�!�$� r�hD�w��`�`f�
!�!�ΡV�8<���QJ��� G�!�DH*7�4� ��"[腱�I�Eu!���+7��!��Rv�AT���z�!򄀡p���p�`J��:���`��!�DB��������#�P-�do �!���g/(����rl�$�E.��C�!�d@�T�r�����w"�LV!򤌡\p��1��Q"? �!�9C�����Öc�t�̏� �!�R����3D��V��!��� �x{!�d�(@,:�P`&�� #�#ǆRr!�$�~�`�I6ƈ"\����-b!�D�$)`	9U�[)�������'K!�� �e���/��XR�e�rih�"OZ�05��G����NL 8���` "O.����8F<����7�*�"Orc�[(q������c�"Oj�R櫃7hiNy1��#9���{!"O0��@�Ѧ2�҅k0��/.� k�"O�0jǯ�X���v��4>!Xy*��'��'��8��iG$h\��fL�z$�� 
�'Al�QRl�3]^���DC:l�����'�*%���>��L�vE�c�.!�'��49���5R�=���Dhh�9X�'2*��)���\AvA��]L�u
�'��;'A�T@����$�&�
�'za�W�������T.�
�'>��w�[!
ö��'�Y,Ȃ\J�'�09��`��4
~���MS�\�E����)����9O3��gÀ k�m���S��y��;ĸ<z2����Ig��yR�M�1���Pg�O��V���$؍�yriA/3�<���gL6�F`J�aƱ�y�A�8#�y��N\m[R�k7��y�S]���%�d���Y�$ɒ�yB�H�,xʥ2oR�Z۪�K�	[���'�ў� i�a�d� ������Ɓ��"OBdӐᐖS�t���/Ȉ$j(�!Z�h���+ZM�$I���'_�s���k�0C�ɻ>�����Y-Ѭm��*G�x8*C䉩��"�+��h	b�Q�eBC�	�4Yr��Ԫ7�.5���΄!rH��[؟p���.#��x%�����e&�	Y���O&~1�
? 9���*��=��'̝��f��a��h	!\�m���&D�Lt�-�-���fJ��5#D��#�F:����3/��bu`�eD?D���Hܻr�Z�[�&�� ^:��ǭ7?��OO>yzgN�i}�<��nY;Z��s�G:D�X��
_��<�s�| �I��7D���b�7d1I�t��:��5D�hq�"�L6����  �F�qh D�����?zjaa�A�S&.��;D�XSN�8&d<��'J�!!KFa�wE9D������)���*M3l�(����3D���oúpvŁ&�
(p���Y0�,D�<�)�"�V�!A�۟`���j�%0D��2�V
V�NM���>��` T�*D��iTe]�٠1��?8lt����;D�< 㭋�mK|�*q]8#�r��6�$D�$+cHہ+)�]"���~�\q$"T���a�D�/�`�s-S/$��2�"O�����M� ��L�1��%8C"O�%��MG�nR"�Z��?z�
���"O�)bUII,�i��H����	c"O�4�u+�<���4�Fbt�ȳ""O\eȁ�F�얈�w`V�;��py'"O�P�mE�C���QƂ�R�,�"�"O.��.�=E�M��䊔-��Xk�"OT<hF� �Z���dL+��m�Q"O>��T<aۀ �6- �@�� "OF�:��2�h��E�%!$�C�"O,�
rU�s4>�s����%2JD�w"O�܈�m�F�d�`F
��2"Od�0�@�aDɱPKV5&��P��"O��2�O�F�Rɇ����Q"Op� Cʇ*h��-��H �;���"O� ���g�)@�4��M�S����"O��	���ͦH� &�b���H�"O�����i,U��B��X�̑(�"OZ��!�'�>�{E��"A��yv"O$hbˀ�YM��t�M.P;�"O�����	Q��!�!ؙI�:h� "OlPPN��`�P���+S��s"OxP�n��w���Q䎓 ��O��=E�$�Έ;�VTi�%�< �4P���_��yrӡpΌa3D�B ��(��yS<k@(ȱ@˘3f�H���`��y���6~�0I�B��-�� ������y�BŲTO�|����r;��Sb��yBk�, Mj|Q�M@�b������̶�hO��䙰n� � ����j�43@E^�lv!��Z>ɔd�D��n����O:cc!�d	��U%υ l<ȵZ�9+�y��	�{�k�A�c%�a�\�%��B�	"Y�~����J��:��Y�vC�I��t��@Ҧ4#x��4ş�r!C��$�n�����K}X��!�!�LC�I*c�b����֯MI.��!��#AVC�I�X�Q�j��|����J��}5RC�Izg.�CF�`%ʅ)�
8�xB�	�	����%C"�h���Ş9�<���<Q"G�Gb�$cP�[���f�@��(�Ob�����(w��!AcA$P���"O���N��r��݋ (��f"O6���U��tAĭS0f!�a @"O�4@��*T+(��v"Ռ5�,u1"O�<óG�~W����G�.u�"O ���HI:��Pc@^��Q9��'�O8�(���+C1`�3A)�i�z6"O�Qz�.S�w\*�H��gf4J7�'��'�P�U��<qv(R�-�8�P	�'��p��KV�Aa�I�"yR����i���O�:��A%��R>�ڰ��}8�'��I��J
�$�&y� ��*�Rߴ�hO?7m�h�x�@��^�0�h�����5�!�dǿ
�� ���*)����䆠�!�d�%V	���#
�:]�����ѥ(�!�WI���RS�'y��`�C@�g�qO���Z�P�����8POl�ے�S�O�axB퉮�&�j�*�#+�Ιs'B:"7�B�4Lզd*���m�b�"a�)R�C�	�,O��k�τ
L���`���}$�B�ɀn��iP �ޯt�IXC�[?i��B��W������L�j)��J#AR���D5?�uL�(|M0����n8�R%_T�<	G��@��<al(r>.���"�G�<��CE?'���q�鍠^��`F�KA�<-♈���MJ"��Dn%i��Ňȓy���K$�A�2e��실<��i��F+z5K*�:ff`QG� ����ȓ؝!a�ơ-Z�IIS &lцȓ�����k� ���[PK[�`,���@�MKF�C�%��G�@�@�X��~E>`3�g#5��Ԉǳy0����
X��a-N;	������1ez����!�tl�J�O�]���m3pD��T̹+�^%kc����̇)%����%#M� %�S���1	?���ȓ*�HZ���r�z0j��T�赆ȓ6h�\�M"Tt���F�G?9� t��S�? ~d�֌Q�b�B\�R�Ìa�X0�"O*i�r+XK�8W�@65!́B"O��*��� �.i�d�[�J���%"O0���߁J�\P��f
;l��Y��"O�,�d(	���j&��at��x6"O�!8D
چa.����� L��dҷ"O��C�^C?��VI
 �<mRf"O���;�0"��J(�0A6"O0A��]�!"�ɏD�%r"O�I!���	>v�򨍞~(�i�"Ot��e/k�R](&�u� �"O��Z��J%S��4��3�n�4"O���$Ж3���9���C�J|�"O� �3��*���Cdk�Ê9@�"O
��"놸���;w�1G�xP�"O�i��gʿ��(q���� "O��H�	?�X��F�7�4H�"O��ٳ��P18郢O��;��yV"OZ��
5-�:%������ja"O��A �[p�u0�@�[��Ic"O�p�d�%q�E��I
,a8�A"O���VC��j�٠��g\!x�"O��&lV;"� &���V�U��"Oq2+�<��G	A���t �"O� � ����=�a���+�%
"O��,�
ؑrQ.�:���"O<3�,��*\IQqNE�N�v�Q�"Or�!"��Tj:e9'�S�0� �Y"O6e��eߖ0L4H�RA͹�~�"O�(Հߪ-�q���3R�v�q"O�⇢_�!>��ѯ<K��T
�"OT)�M�=(`��o���ʸ*�"Ovd`"�M5+�j�QՏM}�6t	�"O�(Ic鈬w����,Y���hp�"O9��HF�N����KZ �e"O�]z	F7J,l���:��"OdA;#�t�H�`��7�M!r"O�X��e�%�N9�#j]�.l��p"O6�!��4��}���Ue��6"O��p�2R�܁�ïc8�8�g"O�P+��_5�kҦ\ F2ZD��"O�\�6��	��)iP�c��x�"O�i�fW�\�ee&��97"O���q��ML0)�%��E��"O�-RU��R����ўp�xKu"O���� ,N��C$�4t8D��"O�� a�Ze����$Ôjl��"ODa�	2�Td��Ò�3��"OJ�s����]*�LȀ���ܚ�"Ob�n�Ӿ�s��g���"O�a3�ь[$�h3!�8X�Z�B"O�d��H�&i�)�w�[#{5^A`�"OF���+�"mDԑ$�Q�i�`"O�()�D˥]C�T���&䄙C�"ON����KzB���c�u 7"O�Ta�EV��Ē���=�^���"O���	�c��p`4�Wؠ-�a"O�)ȴ�اg�8q���	�I]b�"O�@*��E� �1/G�y� "O�(����2DY?����d�<�$ㅐ�:8d/ 7�x`Q�f�a�<)g[
`� %!�*K�*�xhy�J�X�<��öv���(��Ȅw� ����{�<���8I:�٫��+Y�(��Wl�<�  �ɲ���h�6U��)�5g�	c�"O�tb�!^�t9��1�F���Ti�"O&�v�A�S!vđ��\�K	�dy"O�A����F���_"$�1�"O�}B� E�mź��Ú�s��0!�"O$=���ؿK�^������}��"ORU���&(�R��̺yA�- w"Ox$s�@�0GD��T.)�Q�"OAq\yܪ��B&75DT��/�D�<I�//H-V!�d�=*,j��SB�<	cC��z4���牀�w��ct�\|�<y@�s^iie��/#^���ǫ�A�<���G9EK�{�V�bDiU�E��C�I�]a�a�lP���$bv#J�
�!�I�8��-��a���T�[�B�8�!���V�L����	�e �Ȱ�!�����`�%��9�&P=�!�$	�2|�h�
Y�X�r%�&&ͣn�!�$��SE� �'��:�Y��x$!��2J2��! a#2�c��b0!�F�o��y�B�Њ@���O�`!�dWu,$0cA)Ξ�\�o�:\!�D70C�ЊV�H�����b�@!�P�E���7HH�(7�@e�+d#!��լ]�acb���\��+�(*!�� �@f���4��_j���p!�S	$ʌ�����:�^�K����s]!��Z#,���C�ᅴy ��4fC�ZB!�I�p����b��z��\�`�PI5!�$���ɗj�M�(,X�@]V5!�*�>@�C�7L��%��o�o2!�$H NB�pr��8#��-Y�@��Zy!�D۟;G��y�Dȯ|!�soX^Y!��:RQ�3 �td�ڳ��,!�$���z���OZ`���	'6 !��&1.=����Dix�ٲ�(\!�đe�0�S�.KBd�93�m�-^*!�dΥi���ʀɓ�>�2`�Ы�;!�$^5]ɲ���[�JU�M�� ɫ!�^~P��C��eP0Ě1N�/P!!��%
��@��3V�����o�H!�4�,�!�
0a"�(776!���I�|(Pg�VHzQ(�#�w�!�d*�̼Z ��j)��"M0N�!�d��V�F�Q!JH�tj�ڔ��o!�K4p�uJr�O�?b�|
�	��w!���Flu��,�3`�Z {��B,XK!�Ći�H�Q'�;t&�)pC�!�!�3.�*�(b'2}d荀�Ҕ\�!���-X]�Lr�DF�V_�P�E�&�!�X�V�� �߬1{z9KФ�@u!�M�K�&�A;uz&�a�	�R!���_~�d�DAڷJe*Xӳf�oK!�ȇ9�hA�#��Ot�%Y���9=�!򄑠^�D�R�ۂn��Y# �m�!���$[���1���0s�&�9d�k��'\8�a�ӛ<rp��'սm���3�'J�����0jf�kJ[5f� �i	�'�"@{���s�x#'�̀c��E��'��A�%�2��g��]:�x�'�q)�Ŀ4�F�[pFB.VuPQ�'J��Z�i��]�⊏�^��P8�'�Y֬�|�Y򯐭Y4:t@�'w���,~Lz�Ö%ܻTn ���� 4�0Ɣ�@��+�eX`LjyA"O��8� T,i���a#�3F58"O� 9��ݙ,���U�P��	 �"O�鉠��>E� �R57" d�%"OV�b1��XP �`a�?J�lؒ"OL���	l|T�p!�M����"OLuy���1����@��I�&�"�"O�a��X�j<	p���?/��R"O�� ���%F(L���ǄO3��a�*O~�C�ꌫSX������B	�'0*�*�,�I�8mc0`Y 4��'�\�"w�A=�l8q4<'P����'#�ɐɝ�I�XH#ψ�����'���iAv�h�K=�LQ�'a Tx��Z('h��;�Ĝ5�01p	�'.�(/Tx	zd�0.4�Y e�9�yD� ~>�U��I+s�be�@N�y¦?Bl]�ł��{4\�:�N��y"-J�!��1۔�Y�)9�4´���yR�ߛKh0}Ї���)<ƌ�cg_��y�N? ��!m9'�]�e  ?�yM�L�"daeV;�~�IRQ.�y2˒+<��%a#bD9�P� ���y�A��_��TK�	̉[��� �y�I���&E��ǋW����ON��y¸԰ ��U"oՠ�EL��I[��ȓfPn�[�h��EU��1�Yb~Z��`�X=�DJ��U��H�WQ�e�ȓz�xL����y��9Z�/y���t��T�F��V�B�U,P�!�䒠	�p@Ƒ�S,08��$�!��_�:��yVB�_b�+��I8s�!�$9^�9(@�rkV�-`�`�*<�!�Y:
񂃠�<6j��G�W0�!�Y�q3��GM��iT�<:�!�ʄ=�r��g�ˈIԘ��q��C� %���J2�4y7Px 0�Al�C�
:�H{�H�>.,\�7(	�YL�C�I4m���P%�6E$|r�� �`C�'k���bQ/S#`��F��J�:C��.�����ˑ�Xg(�x��)	C�	�3\���ϖw��̒%k<��B�%� �� �#ar��|C��ȓV�$s��_�7�<�S�K�vpl���s���nŻR���G�<k�,��r�%8�E��1��D���4��m��AZL��$BC�J?�Xb6�
S�f̆�e�@�%l�-\ �bQ�Lkv��ȓ_��$A�l�"҇��J����ȓ5�2��6�Զ_)���2���a,�݆�/�����4|}�`�H�����PP�󃕉w��$:% ,&"���m3*$x�kǂQ�b=JF�2c�.��ȓ�H��ホ)<�`�)wg\*^��,�ȓ�|��u�P�F��5C��_ j� �ȓB�̳gžZ���j�f����i�ȓEd*�����)D�M��ꜛb@,D��4�yrg�-Wà��F�>�J؇ȓYV����U�y&%�U�\�jt(!��8f� ��%�P�N(��8fi���j�cD�CX���bEЬ\w�ȇȓA����!�^㸱�&ޥ5U��ȓ%��t��M
$!���傕d����ȓc�,��Wᚫj�@r'��X��S�? �iy!%�kh�E���cd����"O���Q�6}�2�(�Hr�"OXȰ�k�@c�ѣv� }B��A�<�.E/I,�xu��Č}�W�RW�<��_,z��9�� 99���J��l�<Y@ δhux�ʕa���5�d @n�<��FKu;.Diր\�`����.�U�<Q��ǭ�
���ȫ,����@�X�<�q��]Ą��%Â&*Y�1f�W�<q�#H� �
Q�B�:�K���S�<I�+�5l�����(ĿqY.T���O�<m��p���#�D�zvl��e���y�J��,��(�6�2kq������yZ2~H)W��W>�z�Ͼ ����M�@9
�KG�&G�UR���5�̴��ZU��c���u9>�j��X�:��5h���g#���@��K�[�P@�ȓ>t*�+�3S��Huh��r��Ąȓh\�S��!1���JFE�=�ȓ|3�p����U��=�g��*z�y�ȓW�RdFO��[d ��&�����%�X\9���JY�$v�U>q�Hх�K��E�2�Ǭ���bP���6	��y~��M!~R
�֎ȕ Sp��	O*��a�3Y��sT��d�l݆�h��Es�&L�JX �ѥO�#?ڜ�ȓG������\ dN^U�#��aU�P�ȓ~��	����t��{V�N9���ȓ":4xE
�_�\ɹ#K׏N�^\��i�  ٢`1H8�۴x����ȓ*3t��1dÿ J��S�E�hx~�ȓ#� + �/��@��g.|,��ȓW����#�E/'��q�&�'.�Ji�ȓF�d{f.Y{�����9;��=��p��j'�D��Ȩ�R(D�m�݄ȓ3����юB �`��P�<��ȓj� u�Ղ
~��Q�	$�l�ȓ �`���2r�x�E�-j�<����&`�GI��,�p5&��!^��ȓ��Y�C��	������&���u����&�<M[��0WB�;z����z0	��S`�٘ �<mKf��ȓmo�D:"���+��D�aG��RL@��ȓ3ƪ�HS���ez<0���D�Q-<(�ȓ#��e	ШԾ����;�J����J
�BL�1젰x��]ara�#"O��+�-7�"�	�$ŔS�Б��"O�����$6�
U㞬'�V�a"OIR�*8w�М��B�
$�X�9�"O��:QC$r�h��A�Ԙ��X8�"O���@",4Ey ��a����"O�9z ��;P�R5�8�>;�"OfU
�b�'Cn��J�{����"O*���IL kHn�أ�J?Ҡm��"O,ݣ�c�K�\0���*֎8K�"O�<��B�h��0�`�ڸpZA��"O0 �樈��\ҥ�ؤ?�43�"O��QP�'�V���Ÿo&B���"ON�Y&�s��H�΄&��3�"O��1&��k���$rł�"O|��D�U�N��v&	�j^��t"O^�j�O�}�|��c	Yw�W�y")������@�O2.�v ��iQ��y�OJ��X�����p�I�Ɇ��y
� �5{Ah_99NA��_�E힐i7"O|$�26:>x�r��q�@1#"O���Ț�7^,= 1d�(-�r��V"O `h0䇢?R�T��J�.�) *O��J4�ǥE���0��j�8�B�'��0����%(�S &F,d�2Y�'(�H�b/�+9�Lq
 ��7VJ(��	�'!�@(���0�>�[� T~��)�'J@�9�
�l6�p����J
�'E
�k!`ۃaJ��� ���	�'u:�
1�RVSb�X��S�b	�'Jc�-��t7r�
�����\��'����͚!2Db����X�t"�'� �y-Ӏ8\I_Uu���yb*æG�Mj�p��8�y"�Y�eyj�7VU�K�y(C.�j4��P*C8�Z�h���y""^-@�4Q���>�����y�ȑ�<�ݱ6U <Pr��r�5�yB�
-KJA	��.�H�s�ď��yr�_tf	�����&�r�y��#�yB��A����p��*t'�	�����y�Â==V	q5��5j�r�C����yRG���P�B� R���Th��X��y����V��̣t�ŏB�4���-�yr��7 B�� �Ǘc,�17C���y�`p �`��$��JV�I���>�y�#Q�p�m���op�z��I0�y��sD ct��d�<u�G/���y2Ƒ	_"�pa'@\%�Th'B�9�y	T�\ "��DEfgJL �	��y�F̔j���@�ŲLH���yRgς.N��	�*>�,0��T��y�)M�W���j_�C���&CP:�y�cO�@0�(���1� �X�E^��yr��1�\�`a0S'��s�dÍ�yr�L�8���C�&�p��À�y��M9Up�D��T�9,�y 7���yRj�+nM3�M<5@�)�jǠ�y�@'0Rn�Iu�_az�Bp���yR@A6u��y���Y�J�Z���"�y�
�h��Q�TY��+�,�4�y���y���ï�D��v(���y�̓v4�2���4��]	�$��y�l|Z|�)B�/�>�*a��yRb	>nz��١K5%{ĕ�5�H�Py��-^��wMS�.<�"snA�<yw�gG�y{"�-<|�#h�}�<9�B�Lt��C�2[
�!"�S�<9�U�ƈ�uD�]i�K��Ue�<��'�5AP�9B�Ƀ�b�ꐂ�j�V�<�$�9j�4�!o�,f�HD@n]O�<q��&��q��<����'�V�<��Ö#�V����-
�x9ԉ�\�<a�j��%���{ O� 3��z�CZ�<ِ倠O��YZ(�f��𚖣�^�<�#[%ff����m�P�:���n�<��c��C�#�`يZ$dr��m�<���3T0zh���/o�` dI
c�<3���9�x��DN.""�D�A��x�<Y�'�b�`(qm��VW Sb�j�<�&�:V�,�[��ٯCn��wJ\_�<��h�c�� ,/�^<UB�X�<!��������Q*dL<�D$DQ�<� �5ɱEW�3����J��i1�"O�����VpU�K0v91�"O@��"�ӱ�ԑ�&~�,p!"O� �t�G2Jy"=2�CS 3"OB)k��(|ن3e�ѹZ52�"O���Q��P���҆��*��Xd"Ot�2�c��A*X��LZSԡar"Ol؂֯È
�z��$�T#g��D�4"O���#,A/��"�V�#�0�"O*UkԬb~���4nU�<�ڢ"O̍�$��:?8��Oh��4�"O�����n�Ј��j�-+��l#D������l�x��DI�hY�?D���g�ߊY6�d0��(�"�T�;D��:��PN^���.U�DQ��"?D��0�M?U$��
�
;aoZ8��!;D�L�̉<��Y�#i�4 �H+�N%D�P�Ԣ[9na��7Jr,�'>D��!��(E����Ў�u$fTҐ=D�,�6C��^��Š׉��/��p�>D�|�G (f�
Ӎ_CⲔ�1"=D��J�I�"_�(�S�O�~N��G�'D����+]3�Y@�EA�.&TUieF&D�`@��؊!vJ�A��_*��xI� #D��C J�`��EP�eK$WN9�6� D��Q���K�)	�ꉚ)aP���?D�8�"��KS������>U(A�3�)D��c�OJ3$D"��%d%%���a(D�$��W�Q���!se �y���8�2D�x�B�7�! QC޲�֍���*D��X� �t(CC(�6(�u��L)D�d�b�Q!e	b�@�	U�&���g'D�X��d>k�$��d��ȣ��0D���筀#<(%P$�P	63����.D�HP� �t�Z0�2��<��$�1�(D���3��13�.d:��)_���a�)D�@�#�7��EB�$�V�� �'=D��:#	u�>�ĂS�6F����	7D��ڐ���Q9����!�=i[̕[��"D������NPr|���ͭ|���B��&D�4Hu�{<踣�*��p�F�(�%"D��Y�$L���à�Z18:�B�,"D����Ƀ*S=�y��ł(�)�G>D�8��j0\ռi�5��HϮ�3f%;D�������
xM -1.�t�:D�<H�ƛ,Q��$ J0|
�Aǫ6D�\���-rh� �t��=OD�U��2D�����o$=�Q��a<F� �m6D����.G*[X2=�����Y�,be�9D���U���<PC���#��h���5D�<�q���lؾ��Ԣ�-ʬ��3D����(�+@�8�h�Z%h��zt 3D���3lQ�vo��%��m v��k+D�d[��ޔ;����T��
}>���tC*D���׏�'�z@Ѳ�PPn<�Rc&D��� ��D}�-�4h�FAX(q��"D�d����u���z�ͳW�L �g,D�P)5�
[�����m���Q�	.D������8��w�Ȩ��=��,D��4��*6N��T�۵K���e*D��KRm#X,^��3e�"<�<��'D�҆#[�r'��4��(���da8D�t�d�G�B��M��MҵF�ԤIU,7D��3���>"�X.P>"]�P�G*O� �����H����!�'[���@e"Oh<�"��=d<�ӧ��w��	R�"Ođ���0Q`r����W�yppq�"OJ䁖�Nu)��� chUW"O�I��S�vc�hiR	}:65+F"O�H��H�s�`[��z[�QY�"O)�1`�jTܙ�0
�>��mx�"O <�!��|�,ᗈ�[ָIJ�"O�9�gGӺ1'�-���
t�Ҡ"O�0��!A )�=㠬�-@��bf"Ob�렢����NV  <�� "OXu+ �J�i�����P�' ��Y'"O�� S˩w��y���2B@̀E"OrT/��L܋��?"��{�"O>����O?�uȗ˒q���#w"OyQf ����z0��?���	�"O�`��)Z�~}�g��?�|8"O�(HF�D���07`�aX��f"OVIP���8j
��2B���Iv"Od��ቜ���#�N]�1��EH""O�d��Z8����-@m�B	�P"O�W䅢/�$X"g�DcL�Q"O`Y��E I��Eۗ7�a��"O8��+S�WRؚ�X�O)d8ce"O�Xp���Q����C[h"a�0"OLԋW(�<KP���#����T�"O ��σ$c�n���K1;�fx�d"OdH{����<�����/E�&���u"O�� ".Y�2���P�eE>�n]k�"Ol��iRs(�؁e��CȪ�2�"O�p��(P���Hq�
[�m�^�S�"O���jB�<�=@��<|��E�v"OZ�җa�.J���jn�'k��U��"O��WE��QJg�Yo"��*"OtQ���>I��.}��E��M�<�K��H�Μ�DI�ܕH���E�<QS�:����c݄p7(�X7gLZ�<��*� ���C� �h<hB��z�<i�i$������94�p@pB�<a�ͅ,���(�M�[$�	R�G�f�<�j %d@:ũqhQ�t"<j��y�<Y�G92M&��@�?-~�y�KAZ�<Ѥ��S��4�����G���c�R@�<!�W�p}�Th�P����i�B~�<1�MQ�_O�	����>�D˲�O{�<QE��h~H,ѥ�/^f��S��z�<ip��'yS���hS.��tY�.Lz�<!w��"kx��p�1�}˖#_x�<9�F\�d�9�BȡZ��u�`�<C��	���B�C{	����x�<��IN@�ph�%� '�l��e�}�<Q��_l���PiZ�`�)�w�Ky�<1�mZ� �"1�n>q�b{�B
x�<ɳ���%j��2�=.�h��K�<��T�sq�0��aW�s���0�9T����٫~V���E7�̑ab$D�x���Ѿ�S�fH�}��qS
#D�`�g��a�PI���1�n��ua<D�d��Т�T��b��<�j��,D�I��M�ḧq�V��F�#�m+D�H���S�G>�}q�$5X�\t���*D� j�.ŰeE I����L�ӆ)D�p�f��;����
]eq�`(D��C_5�@��B�-u�� ���9D�� ~�R�JC8k��{�l Ob�H�"OF]0�*֢k��1(���l�4Ak�"Ot�z�x�I�j[
'�`�J"O(��pg��и��G�/�̓�"O�R�L	����#�0`�"O�P�bo�d�p�'�Ec��q2"O����Hn�z`f7`>��V"O��ӪW9<	�a�DU�*p���2"OB�馨@�P��M�4Ɍ�vi�f"O�Q!ƕ����G�$8 p"O�Hy )0#2Q��oV2-�T"O���H�nq�L*7��*4�D"OhPKY4O`�p�i�V N�9"O0��)zҪX@eT�m�B���"O,e�C�F�fz���@�2�VA{"On\��ē�b�+�aS�|(��"Ojd�R8E�d��W
E�
dRl�"O@
S�<D�h���)Xc��3�"OP�P"D �`���GQ��@"O��[�&�dc�sw�8R{�a1�"O�q�cn[/P>����5hIa0"O숢�]%ye����Д?���B"O���R��{b����S 2�� "O@��«�ˮ���±oJ.`D"ON���f�7F��*AM�*bEp��"ObTiC�	�=��(�m�5:��(�"O��A� �TSb����[�C*�D��"O���#���-@�廔n��5"=K�"OV,�"a�/4D��ٓmɰ$���$"OIH׏������,-���0"On��Z�x�
�-R�`��c"O��7��_=<�p������;�"OND �$Ֆ|$ڀkM*��"O\d�w��Q����"I[&%zjИ"OI�J���(0�ӈ
�p���g"O,���s,8��V,:�\�A"OL9@��0�By�1����.l�"O��qU	�p���
q�L�c�"O���nE�,%���Ӿg���X�"O�K�m�N`�!�ՆH;ƪ�ڕ"O0��q
� {-���'K�	�,��"O�찃�	Wmf �g*ڑl��!�"OJqϖb�r�j*�G���0"OPĉ�
0P��Däz��ؙ""O$��7�]E�q���:�luk2"O�0j��	�� ��\k0UP�"O�����њ5/ 0�@dۍs�X�f"O���d��.L�"CQ�}è0Q"O�2Ro�3)��h4�Ť�b�"O����J��a_B⵫PR�M+g"O\���I��UF��D3��˕"O\Y�碘�Gs�亡���:#:�X�"O���GB�!p�P��#��vs"O^i`�-�:�\�D@���Y"O��Հ�dZ�	�^-p�JG�s����6��̉"�L��x�q��tY�ȓS��9��V����1�gҋ`v��ȓf�l�K�.-�����c:0��&M�1	ҁ�1�G+�:ΆЄ�=���Рִ`�`\a�߳_����4ܨ�M�KiĐDGK]w\@��mr8�2�˸B����Á��ԅȓK	l�04�1*�T�y�Ļx�d�ȓ����6��_69B�%P5C	���S�? � x��2����O�ftX�R�"O�ɻȜ��*�f��"O*i;�����"e���4�(��"O\t��m�?��q�-�'�Q{"O�1P�,�:lŬ��TeܠoS<���"O�U�6,E�x���PFF<LZ�h@"O4��UJ�&A��U�fL32D4�a"O��ҒDP-�D�Aŋl����"O��	��ƨ8�jm��K\1x�윹�"Oh�8E	ϰG��#�ô��qrF"O�KE���A��I��T�
�ы�"ODP�r��.�y#��=�|�b"O�dQ�H�^����Śa���$"O֝$��p�0P�	?� Y��"O���2�ߞ$XT���
�eٔ\��"O,ݒ�AٸK��M�1�˺m�DqB"O~���Ա��{�
��h���"O�ȠWM;KVrmx��ċ���K�"O�zD,�9D�H�c��,B�!�� }"��Q�en��Di�70�!򄐡� I�@]�!��
?%o!��>�^P�P��%�����O�?aB!�Ĝ�Z�	��K6w~��-V(!�d˭aѮ|@D�ݬ	b�Q��^�il!�DL�WiV�i'g?�T�X#��'�!��ī/� ���jz�H8��P�+l!�D� �l9�H]��q1�<XT!�$�ȴe����.X���(y!�G�+��\�P������"d�!�V�*��\sb֞	�d�kPLt!��K]��Ԩ�`�'A�\3���7?!���)O��ǃ[�_�HiJ4k��N!�D
�2�"�����:�dA%^)!���$�6�;p��S+*��1$!�ă�oF��J�+�7;:ֹ��#Z�yR!��)�8���F;P��01�@#!�!�dX�=�h}�C�
�jH;�����!�$�U�j�+��L�0z���� �Q�!��˿:� <X!,�=��ݘt����!�V�E��|�W�	�Qvd�Ϟ*�!��c�~]I��_,hA�x�/�7�!���d��P�-��Y��m��y�!�$  w��c2��*"��}jVM9L�!�$��E? �!՞ ���5�� !��45��l�'dH���� �?
!�DL��>iHV��5��36�3'�!��V,¬{c�.xcΌBG'^�.�!�d-�fT�%K��z1
�x�ƀ�^�!�ċ�
A�C]3�@��Eƹ�!�d^,<���2&lh!a�U*-B8�� "ON=�G��`1Ĭ��ϐ!�Ny�4"O�-zÌ�'"�	!���a��Hр"O^�P7�̬My�L�g�)��"O�u���ޒe!f�($�аM�(���"O����x���N��mrr";D�lx���+�H�Q�N�V��#4�.D��sN՗v;�`Hr�R�dP��� �*D�x�u��\��q��*%2GF'D�xcG��R�;f��7q:jT�v�7D���u�:W$��R�M`��5�"6D�8 �[/����p�/�z��+3D���%g�W^�<�bM�T�z�J��.D����
�>WaF$S$��
�*�۱-0D�hsQ=!�4h�C ������.D�� �T�S!#'��JE�	�G~� ;�"O� s�i_ U≯B��Njy���"OJU0���l��8���,bl� "O� 0�m�	��;F.���z`��"O�E��dY�F2� �&NZ�*���c"OD��c�1��rr�%X"���"Ol�cB�0�����l��!�"O�) 0��,�2pk��_62�0���"O�(%V�3ZZ���B�!�����"O�p0n� qPP�1�R5J��q�"O�9S����)�LA�b+(=��"O��xF�ƀE�,8��K՞� jC"O����7:�T�'lY4��`p"O~���߅^7�,j���&�9�"O�œ"E
D�I�P0|k���"O�V�VP���D"t���:�B�e�<aa�G�w���뇍�!��XB�Ky�<i�aY�#;b���j�41�f�W�w�<��7IдAJ�N�3\�� �D!Jz�<��(�'/�d�B�v�^A�4#RM�<A��t�L�����n��5C�u�<!U��}:��F�:a�d��@k�<��J�����p"^�]�%���g�<�e ��/��4Z��']�IYpKFJ�<���2:�2�{���IK���!��H�<a���O��a�+��>OLtC�p�<��-ԵP@�Y�V._3�bA�p�o�<A�ꋐ�Z�����Eg(�cь�C�<��G�q,l�c�� �I;���f�<i��g�������5 ��_�<	���!<�ROވ=��b�L�u�<���E�����4!O^���zfGj�<qq�C���I�i�k�f��j�h�<�R��j8ȡ��H��`[qQo�<a7dڹ0_�Mi�,Y4r����u�<���@�8 ���	be���(�]�<�5cW L� ��+�:^^2`���b�<�q#U�|;�v�tW��ҹH�"O^ҕO�7w�	��ʭt�^���"O1�B�R��6�Ts�*y6"O�!�1D��\$cU�6i��d��"OB ����?ɸ\�e	�g�d��"O���b/*E�(P���HR0"O��q�"�L�DC"a���P!{�"O��
-�%b�<����ڸ��"O�`��Niv�uළ�2_t��S"O��3)R<Z%$���#d�go��|!��9Lyp��'�Ń)Y�p7,��;�!�diF�aCB"H�9��öd�!��U�j�\���GQT����B, �!��oǦ(2�M\��`�Ұj�T�!���r��с懙�\1��
Gi�$�!��ҍ�����KX�Er��_!�o�����k9�̑���!�dM)B�	YA	���͸S��7!��:uW(!��cV9XK�i�!�Ȇ�!�ѩI�ݡD!]�<K�k%ʏ>&4!���s�!�"� c�ɨEB�.{.!�$��+覠+�ŃpY"��b��!򤀫`5�䢣 �9g���bD����!��_#��$�rcD/dˠ��b��-�!�d�t�� K�&�8UcE$U5!��9<�����׏9�8���Q0!�$�>H�y���.ܒ�p�C�<� ���ϊ�t�f�ؕA�~�8%{2"O��ۓ&H�L־ͣ��=&�blp�"O���g�TD|<���שO��q�"O�ԫ��:J���J7	S�$�T"O������k����ˌ=�V4
"O*�#rC��'a����Ӟ��2"O�1����(}���Y
� �e"O����0 �T���k�,�9bg"OV|xC"FA2<4�U�J7����"O�D1w╏l¸ݢС�'{֪��v"O��*Ei\�#�$񲠎5N��l�T"O�q�'��,� l��IX���K"Oȥ�E� H\P)���9t�Z�8�"O�����/]����f��w^�2�"O `KJ���G%5au�$�y�kh���It�ʸD��+Q ��y2H�=�0Wf��93$���L%�yb�L�?�@و!o�.[R8Z�,�yrn 5I�h�Ƃ�G
���bb^��y�*��r<����0g.��bٚ�y"m�=��1��!~���s��>�y�I�U0Yz���|U��D̵�yR�S(g�JU��n�,y\ �y�._)uݬ ��]�&h�q�y����&����E�5���s�[��y���1>6��Hv�� -���6k:�y�gJ�7,`A2��6�f��
/�y���^�mY2Ĉ*{��DI�a�e�<q�/K�N4�YZ�-Zo�\p�ҎZ�<�u38��d��ޥ@Y� �c�|�<�T.�*_8"a�,�"�BLFp�<����-U3���V&�o  ���Vk�<A��ѫvfFL�c�V�l� �mV|�<9��G!°��%C�YJ�jR
w�<�E�3�蕒�iŷ
PZMRsK�<Imc�!�5&629��I�<��E�:/\�@P�4sޜ�Yi�C�<�&앧8�B83q��0C�x9ֆ�Y�<�gM�4An��5l��C��{rn�P�<�"FA�	�dݗI�8����Pq�<q� 5z�ʅ��ۛ"�*m��
D�<�� ����@T��?+6�l#� �X�<�An|�X���?k�@'�U�<���c��&�9N��A��Q�<fO��T� �J�7�6L�BfK�<�цE0C��Q�⃀�`���P�Hn�<1�F����`�e�9�rA��g�<qGo]�Z�z&FT$��3���<	"���2�0�Ё�тm����B�<�D�G>M���EFP�E*���m�~�<s�P0w�����Ӿ��ݻ�EP�<��/��>p� h�)��օ��&G�<�3H�<d�����Ғk�q��|�<�@LЛ1����	^�|P�,�B�<���  (\�y�oS�Y<����T�<sS�1
�@�D�	x�n-�&HFi�<� �$*P�s*�[^V��ʔc�<�7�µŨ�;�I�<?z�[u"�`�<��$�B�q�㗻P�<��V �P�<���+Q��Y�S��UՔ����AI�<��,��'w���
��)���_l�<��+;��<Ѣi�+M����CB�<OR �)��V&N�B�#�@�<�"!R;�b��E+Pk�x8��~�<� �q�f�ʠ2�`�Z����rC��Ӗ"O��Rf�^�X�~I����)�x"�"O�gp(� �J�P�4Y�"O��y��"�V,2 (Q�+���"�"O���@׀tY���ڔv��D�"O��مN@�d��b礙�{� ar�"O��8��C+Y���b��O�_(>�I�"Oܸ@7��4	�4ɋT"��"Vy:P"O&�#HH�[j�q{Ҧ�7p��w"Opx��M	J���2�c�3FԈ�"O:\n�M��!V�X���G"O��B㖻 �n=	Ta�8V~L�#�"OZ�j'���p�� �9S�ပ"O,�BW�p,
��eT��@6"OTāP�0�,�Q����,��"Ox]�RN�Co�1�&�\1Er��+�"O���lĪ\g�ЄL�EC�Ur�"O�aJ�nO*37LѠ#k�!nJB��"O~�.
*e*�a��lĞ3�ZE"O���W�łn�8@�$�ף]���"O����2�Ezd�UM��p"O�i�H�2�C�@<`ac"ORqQ�F�,/ä���Ǐf��"Ol� ��|�PQҦ
,!�N��s"O��{���r�l��7�"���f"O�\�DiY�jz����b÷g�Bk'"O� ����mF��"\��LH��"O�����OR�b�|�L\�"OZ�)�/��22��Νs��]�"O��#Ӭ��1��w�]*�T�ɵ"O���F�ԹK���֤S�3����"O�ٸwGPD]���%Lw�=P�"O���fK�;5(�3v��&kW�-�"OR�	�D�Ɩ=���\ H!�"O(U�ծ�.Nb�Гh�K��kU"O�h� �B֔��H�#X����"O`H� �צt+z�A�d��5� ��"OzBUN�Y�2	x�Wh�"�U"OP��a�J����dB��Ģ5"O�	1���)C�`��.<�z���"O��K�臓m�2�)���=Ҕ�`�"O�,�7.�7v_������`�P7"O^��ܸN���дj�4@��@go D��R�B�#-ql��3d/GR�V�)D���b�tr� �e�Z/��0g(D���R��v�3��!|R��gO:D���7�I�W)Ҭ8���*�n���D7D����Y L{�����JF1ɡ�4D�@16��{hb]Pb#Ǣ^!:i�
1D�����m3�-pb��ؕ�3�+D��Qejؾ)JB��$�Ĕ1�pd��6D��s��{ �t��'B�xj@�`c3D��q/ւ����AI�'�Pk5�#D�ċ�g_	�\=�#�@�>�F�Ѕ!D��y�_�p.��&#(x�:�4�>D�8���=F*��ӂOr~����)D�<�ѧ�"	xB~�B�(r�>C䉗�N(�mY�oBA�C�G9�2C�ɣ �\��%S�H`,9r��$�B�I`"����ʐ>v:�3���h��B�3i�T���Ԁ+�t4��LN,#k�B�ɛ�Դ�f�N =�J�"��L=xB��W9�Q��GO��pa�V;�lB�	�"���Yb+ �J���J	X�cVB�)� �RŪ� �@t�4I80��I2!"O��h�B�f� ������"O6���ĳ,�h�X���x���"O�Ai� \�2?6�����+�b8"O@�G�1�Y���S)��Ss"O�lѐ!ZV�\!�#�̟y	��"O����9"2:dHS���d���"O�h�+�#�-� L�#[�aW"On����#8�F��Q��:R�̹Q�"O����&��H��R�([?g8=:e"O�MI+�1�9c��WVN2��"OJ��������h�&?I��"O�@�n �\.D�0�@,DH�1s"O�]�#�چhJ\�@� L!OCF�cQ"O�5j�B�#�VaHf!G��ƙxR"O�ps�d�t�r��t���v�Ҽ�"OR`�ᨁ�H䒉��,}}��b�"O�Q�Q��$?
�����\E��#U"O������ }pG(ٕ}����"O�-{���&=B`RfᏰ8�F��b"O���-<C<10�L��R�R"O����iY=@�aB%�7ư�ӗ"O�1j�j��!1����b�҈{�"O�T��뜝0�;1��$��P�"O����a���1�D7+(lM��"O�93� 8^^�x��ס(j�{d"O��A1�(�
S��?����T"Oze�!͐-,�,�y�L��8R!R�"O��%֐CGn�4e��J�u�V"O@��!�^�D��P�_��X�a"ON�B"��
2�5�R��ݐ��"O���쎥ya�5aQ(�
�r� "O�x�f��4}
,�s��=g����`"OFaI��DD �2g�"�eQR"OZ-EH�.UU����R��c"O���!Lɸ( ��ff]��v��E"ON=�b�\�Y�jC|4 ��a"O �+��/�V��R
�9'z�!�"O2yg�'3i���§V�\�0e"O�@*7$B%1���,2uPJ"O����Su�t����lݘ�"OZ@�ܧ'4�Eᱤ��x|
���"O&L���"eB�\�d�i��PR"O�Q�Dh��B ��@OW*S���f"Od1#�K��
,y���L�03d�"Opq
���w�DJ�nN�Rv�Y�"Ox4�� ��EQ�A���R�g�6�"O��KFVp.`լ�/�̭J�"O,p�2f�&I��؀�M8���R"OT��(u^��	�3nz�3"O��BqB��sT~,"��	5�
t"Oj4�P-̋3�r�2�L#�� "O(E���Wy�>�P��ÖY�2�"O��D�V?]	(���.���+�"O0�hE�Cbn,��*VV)6]��"OI�ߏF����Y�H�&)	�"O��,�u��؁Μ�!����"O������b�1�5b
���
`"O�I3cL�G*�����CJ����"O	aҁS��%���X3f_�] �"Oe�#��-�l�"umE�xb @�"Ox�a$N�0���- �m���0"O$�ivJ��}�x��v���B�PQ"O$e{��E�������q��H�"O� P���J�0eA���%ײ|�&��p"O�р�,�34���'�	��-��"Oz������<K�Q�&W�S����"Oa�rj�?C��Fު,|�X��"O�tؠ-;F����e�$��|�V"O����(F�]gΈ�E��(a��]�%"O%03�^#�~%���R���"O�`�u�ՆMU�3��8*-���"OH�i���|�y���Ծ@�	"OHU�^1mN�-:�B����G"Om��D�%: @�Vb��XL�Yb"O��+�9x�Z�YO;:�	�"O�8��]�\�Dr���1 I��"O�=�un��R.I�a��	x 8Cc"O�a��.�zz���j�-�לx2�)��2Co\��@յ;S�Xؔ	�X"�B䉳Z6
����� \��L0&V5`�`B�,6�%xL͓g�Dy�Ψx JB�	:?"t-�c�����+KA�C��RB���?L#�P"a$��^�C�	�~����&G@��.�B�J��:D�H�.��
�
P`���@�)�<D����D�m������X2#%�tK(D�,A�N:��@ug�j�����;�ɲa�az�IF������ʘD��HS��]��yr��9?tp�2�R);�:�RF�ǽ_'�7�-�O�1Â�.jf<;��ղTOX*�'�Il��߅Y�	�0���f[P�!�d��i/�ܰBC�l�H�;�ɷ|�qO����R��_K@�r���%i����iա�e}�!��^f���A�ͦd�!��� 7����9}�lQ����!%�azr��§S5L �R�Un5�$N!OK�7�)�����!9���zݶ��S�5D�*B�g�����ޞY����5D��AS�_�<m�Q�te��_4���01D���d��le�"�i����ke�0D�8zw, �Y�@�(�&�Hڈ��B�+D��Jҋ��;�Lp�'J}�P�k�O)D�(����Kd9��ǧW
4�q i&�}���O<��c-ZF�����"xy�!	��Mc�{�̇Y�4𔨆�3 9J���=�yb���,s�i�0Ɣ?
�xTJ6GS�yD��2}�d��b+Tv��I@�.(
C≂O���c�OX Fo�J�,�$$��b������%�ӓH����`S�v>\!(�kì!˂��d�<��g��ԩ��%Q�J�;���@̓�M#ݴU/�O��_	�Qs�F�>fn�т)ٮahf�����Y©W(^���m���hɇȓu�H{�m����1�'�Y�:DxR�'����O|ӧ���ޓH�V��E枚17�0�"�
fn��Ɛ¶H�"�'�x��ݫ5Z!�κ&70q�ӏ��!x8���ŲiNa~�T��� ��BF�e�,ͬ����)?�����=95���V��2!-{��P؇k�t�<ɕ��$`dd��ceW�S�ޤK2l�t�<Q���ڬ ��R`�]3W��K��%��'�`��y�A�H�	�d��Z�C�Iچq�B s��=����\��B�Ɋ]���4j��u#t\:w�u��B��,1~�S�C9_�@�Q�o�.��6�/�D�<E��4PƲ�X4�Fv���E��MԬd�ȓ{�6�a���w�P�Ь�0/j]��#[���疲rCj��n�
I�Π��Iz��1}
� ,�A�咵l������W(ѷ"O��i"��f}�ɒ� *r�+cl&�S��yR����p��p�F�!+���,R�y򥇩,ƭ��en"�B�lҵ�M��4���&}���i)BH!d��Y��*'H��g58���'v�48U� C@��3"�2����'��hRV]/���a��3$,�����'�I��v��6�Q6���2�Ɔ�%�C�	$d)�d	ϣ:�h���t�4B�I29R�I��
[����I�}H�C�ɌO.$���"��|�� �5�Y�o��B�	q���g��|�thQ�-�>~�B�	s����"V�X߂EQC�
N5�B�I	c��ku+�>�he��D�.��ͥO�ӧ��<�H��4�ߍ'���Ӈ
U�~�����_h<4NF4~.�dq���{F���SV�<)��6 p��mU�]6�m���H�<���A}Y��A��M&H}s�&Ʀq�O�ӧ������o��5i�M��� �D9�yR��[^d cI"I	�U�cА�y"�cL����q��<3�Iѡ�y��)�'s�p���L�e;�KE��(����?A�J *C����"ѩ�2���#0�.���
�|��%L�jz�iQ��DUJy�ȓR�F��w��s� y�L��&�<u��y Ur@lD���D����p��?ɞ'�Q>E�'u��Ǫ�%T.R���)h����$�@Ph	��X��qĨ(���G|�����~�vg�.Q(6��c����Y��~�<ia�Z�Z�B=kĨH���i�#���&��5�5���n�gh@�b��݅�I{�	�Z��i"-�>NY��JL�Z�	A����S�ΞfE�e������ZB"0D��襢�5���l$4Q��1�	/D�8c�6�@q��:aI�`X&m�ܢ=�O��O��A��Vf0�@�:c�ܠ!%$4���Љ��)~��5ꃕ2�lU1AL�O�ON���E�-�蝆V��BAV6!��>lqz�cq�;]��8�-�d�!��2_P��FEFn��e�4m��D{ʟ�2�(=
� T��o�%g�vx`F"Or�q��ZD�Xc�πd�Zu!3O֣=E��k=�R{� G2ad�@�mO�y��O�=;`�h�b� "�	��yB���A��d �K�fHQ�tHS��HO@�=�O�����1S2�(p	ƴ8�(1*��;,O�˂f��
��NZ�����"O��a�%M�6�\��MH�Y�� ��"O:��3iO������+��=KR"OV ��ds�|js̚��51�"Ov`)��H����f�4
��QH'�'�)�>��)�:�Њ7@_Z!�IX�J�'��{M�7+JpJ�K;�A-���1 _��:����M����O�>��f%ζ(�I��Cӗ��<���5��2�HVfO�-+�R�|���v�Cpi��#���O2���[�V�F�㇃E/u,ɐ��8�ў0oڪ]��>e�PB��y�(pC���W�@�A�D�O^��$ū���c��ADD�4�$dE�c}8ȉ������4Ϡa��Lܛ9���hW�5Q��X�c-��B����Ќ6lJPQGk�%����'�4 �2��z�S�%-�d�Ѥ�c��p�c˜V~��l���y������|rO�,7��Шr���2����<a�@#=E��'F��b�`K�F�2a1�o��zm��'H�}�'��9&+2lxL��*m`r銚'��
� ���M+$�<�q%K<Q�p�q�"O0��4�G {R���V�-��$"O��A�aеq�����O�v|�̡��MX�P��Z�8E`9h��j�(�
�H7D��#K�52й@7e�quJ�e*D��٥,�>4���ā3`����H5⓫���$7h�`t �����2�'I�|�0�y	ǣ.4��K���I؜��I�i���F�S�Of�4�#`R�R����Hn��!�"O^:$�ٯ�&��m� {f`XQ�	@���I��@l�<�fi��3�ܒ��	<!��rQ"XrB�F!�V��u@�'e(�Ҧ��*v;����C��F��y��'�T�	��NG�<%�29��Y��'9Z�*�j�]���4#�%|f]�
�'@�"�4
�� �]�hk�'�Qۥ����x�# /X�
�')�����UG�["$�%���'�
�8@F> @i���	[6���'�q�Sܠ$�����R�����']~yj&��'���I���"# DH��'�
q���^�k��C�c��22:�@�'�"�`
U��
6M�Vg�E��'�Rd��M�eK�JL$R���'�����F3{��1Ҁo]�G�Vm@�'9*)�cHǈ;���p#Z�9�H�'B���dCJ�w?.���&ַ%�^�B�'HJ��#e��)��� $W��'�B���@�/ .b\��l,+��y	�'�@q�� �%!���W�W�
��TJ�'q�H# �͕K#*���c�#:[jŻ�'��p�M[7y
����,d�$P�':��i�
@d%"���[Pԥ��',jM[���~��U�Lh{Фb�'�Q���Ao�\�rŕ�1��ի�'�Ab�B�z�͒����*��X�'ht������,Ć�����5����'C�p*Ѯ�2���8!m��8rBU�
�')�`2@oM�d��s/��0��H��'��%`w(Mo�=q�!Z�z�R0�
�'�,��f���L4;�@?l�Ȭ�	�'���k�I��m�TxU�j�����'i�tH�)Կy(|H�G�m*���s8�q`�^Bb��
���>���n���87�Ԙ�� {$���6�Ňȓ6ۜ��u&K�/V✢TM:s�6���c�@����(&づY�`����͸"mA/Z?B$���9"�<�:E��Z�x}A�fؑ[�HB��/U�hj�EY�I�⤁�L�� B�I�N*xR��'6_����U0S�B�ɠgxNIJ�\�z��Q�vHІ��B�;�9z�`� ZY�U��Α�M߸B������j�2B�����	X<
�B�I���)��'Rv�pM�VC�	<`��H��+,Z��m�T�)k�C�)YUz}jpk%\�f��ь�j5�B�	��f��vD��t]|A�(���B䉡`܄3BC�P}��N~ɨB�\ǂL�R���B6�Xca�6,r�B��?�����߽[���C䆚$��C�I+XQ�5;��?@<Q��e��5�@C�I�c��{ugݖ	Y��C�V�
�PC�I:K���a�$H��(���@B䉉�BXsȕ�Ir ���׍!DB�)� �(�F�~uh����՘Q����"Oн��@�r$�<B@��5G�b�`%"O� �V�! t@Xr�U�C��k�"O�4�ǥR�C���H[nB�h�"O���`iQ*e�4��g�]d��w_��$�9�qOQ>]�DL�Y���)�\R��(D����iNw�l���óxZ!�0�'}BK�f��Z!LO��c��^R���ߔ)�8�ʶ�"�ONm��^J��1Sb��G�j|)VG
3q���e�̐2'������!|^Y�EO9d'�#>ў�x��H�T�z��΄ �O��ݨS��*7�4=xM�+����''r`L��-;�5�N��yB9�M�<��2�\!z��0�g`��"~�F�,��@�g�k�Z���l���y�H@��H��'M`�Ν"�E6� %��$	�X@��]+WV�]I�����SR%f��C��#@Q4���+�O�d���rA��Iq�A����M.l���iF�>P90T�:�OE��_ �
 �D��Q�Ĉ'�ɼ���;P��\�(Xr�ON��R� .P0*P/�=4���NU(&!��]�u��x�hV�
$
�PT��)����ՙ,��"�!E���Iz��M�\#}�1;=dl�aj��$|�ˇgG,]ɌE�ȓ~���M�D������.vn���M�0+�P�!�9l�T�:G��m��Ƃ���'�~�j�i�`�<$���P����-Q���`xӌ�JE�/x4r��>�:�Q-�V�T:��3xYP�K���g��x%�!\O�\c" ����!QE�D���:�[��S愅"�z��/1Җ(��� <!kF@`A�+u���C�� n���S�>l��8@#۞Pц��b�BCN�T�ơ��#�A��l�F� 1��+5ȝ	7֌	�+��r�##�����C6f���1�,Рӭ�&�����َ����'bl(�C�6"μphV��5��@�P�L7P��#,ʄa�y{&
J�H3���!ɰdHf�5��h�H>�n��m.59ᮉ#sfuK�H{�'�pI���S��$�vi(䜄r��┪Q�[d�Q��̪H��I�aF�"K������ք���D��Ҍ��8?Ab&��E}V �@(��zD�TFC�<Q��E1� Y��F&O`<�R"攝@wB(���Ӗ{�lp��&�, aH�YC��U���˗vH�T%�J�5�/� �*�Si�ϸ'mVDҲ�ɳ�dhG�ʓ@h�hT��,��(;(�p��iT�ƈDbLt�2i�2�pX��KE~�0���/̌X�T��-_&���E	2#\L��l�M�L̈́뉗R��K��0}>A�#lK�#w��z��ȿW���'S8̤�	gX(U,��+e�3{,q��� s��J�⩟��P�Ӊ��Yy&�
,!��9u���}[�|""=.�~�8Ae�>?�(]ѥ/˧�M����=�:���P8 4�ˁ�Ȯ.v0�c���M0����:\���z��u�����O ���S�B
&�x����vP����'G.@���N"�:�%�;x���4�@�@�9-t��;��V�"��*��M�5IUa^�D��R�)�?QS��R�����:��������Ǉ�#��hf�H �䨁
��l#��co�,a�i������6#��(��	�����
N�[.�\;�D�,��Y:�91���EBȷP�H���I90������c��+�% +.���,ЭVr�0@V/_�[�
�B�;��r%G�g��Sa��%���CLP-Vp� h6��L;�X31�P7e��e�P�N�£>ф#	�[UV@��]E
]�D|>���G?obx�V&X+��fiƽ���lb|%��Y�,��ᩕ���t��v&W l`�����Yl��x�B��E��1,�|��n��C �O�ia�F	6H�h�\x-&J�/cw���4K�h�\����+�!:Ǩݳ��86����W�~d!�Sڼy�6�{s �x�jq���9���G{���.�\z&���.r�*U�_�]��u�bn��e����g� RF�!�E�4-�DB��ڼ+y�"5d_1\��Q�b��VY��#A�4�"�cbND�~	��0EA\2a{�o���08�3X���d���v��@Ɂv�k���:o@,-I�m�/
�0G��L��&��p����r����@u�4h�E��'Ӛ��'+�]�;���.����`	�����"A�T�dN5;�$"�[3�2�IB��T�#�H�%��-��� G�@�A7>�S��E�MJ�f5z����4�	���l�<�#I:|��D�a�&Wh.X�7iO9����,M�A�e��H+¨y0��Sc̩��Q�8������[�PXv|q�ƀlc
��C�	��hO&p��H_�k�́�'�R�CUfy 5dC����fʝzA.�$EׅTH8D�!H^�o�Ե��$ӍG]tUh%d���,��U�Mz%�6C�L*)�e-�-ZU���7�O����B��1|�� �AH���
��'�e[Z�`���	&B�L�&ď��O��(CBg�
~��lAAN�g�¬�©l~v1��I3hdXX�!͵9��уE3�{êX�K(	 F�#?Tq�C:7��y���O��!�J"�ȕ�̂&	 �(@3�Ў����17r�A�,��&�ru�u#�$h�1Ovy�#T�m�z)+����F�<A-�5\:Hy�'�R��%-�Z���E�
�jL�����:_�&��U Z[��<�d�=�F���	�b��8s$B3m��d@��͊J�`��6M0�6(K�V҈��g��P�dC1i��DUgL�M���x޴�L����`���Ȓn�	#rTRaNխ~�<�-�ҥ�Q�H�[�6Z@�KQn��b�������.!���h��++�̙�I�t�a*¯P[�cf@C1D����!04��Sc��1�`	,�9a!� zx����a�H
�X�57��F'h M֐>	�H�K�V¦�@�M�J!��G�S���I<�й��N�}.��֦F��t{c� 
�d���N�:q2��Iߵ3<=ȠG}�Q�U�a ��b��� ːQ�^-4�x�bZ(�\�A�2aq��b3ړus���G�-&���a��O��@w��3|~�r�i_�r�f��oK�qy��hC�V/"���	'�� I��&N�0�*���� �r1�RD�+tg�d`a��+L�0R�'�Z�#�FËZ�Ze��dW(=�&���	N�J�bI1�=Dh��cl=��T�$	�7�ZQ�C�V���䓧X�Rd��N\�z5rF
��O�*�����Zc�е�I��>�B�,T%!��Y !�J�o�Ό�K�/G�Fu# �Z��i!�gE=y���D�F����1,�����@¡����� �6F-��,�|<4�0+���?����<�E��MGw�)���=�`<Q�Û��]P$��q�@���ƒ?�]�p�A|�i7�վ
�~ � ʆ"
��a��F>c�����۞
�x`Qr�K�0v�c��m����*��hOl��0K�}��}p���c(�؂��������^q��1If��MC����9� �Ӱ.Q�'�@���ta�%(�w��K�.ӛw<���]�`�HA�}�'�6�Q�c��e�Dt���V���y��2�,��^�q�F��2E��;�d�A��u��qbw�B���z5��*m�YSF��{�����U6�P�+o�p�W  ��3�5@��ʁDe�cX,yh�Q`C �$�񭋙\)ȉ�"l�q ��B-1Ѧ��U�ݫ,��I��|�"旋q��(�!��"�t���6,`|�3wE�-@eN���<�F�R���p_ �j�F��Ed�s!��3"�'%A-@dJ�(�V��L���:v^8���uf^��?r��5-��)f���#z�<�s�P�Z�����	skD9�?��	��%�X�[��
s*�I{���~��)l��b�ܸh7�6cVh���L� �V�[f��S1��-0R�	2�F$|�b��d��Dq1��X&O|d��)�,L�uEy�d��P]Y`&�#Gr���KQ��kT䔡V�H��T$��z���a�H�FFBR���II|���/�;�ĕ�S�Z���-{��j����v�lj�,|��`��3uʱO0T��L�0V��ؠG��I���k�l�'^��%;�'/��	5�ɨn����uG��}�}A �ۘV)����i9[�4*`'ۗ'��%�I(o����%��!z�U�;A�	�&T�LZ����-���y14��<kV}�$勜
�F�	0��B��K|�`S�/�$�#�JS+HtZб���!� @���Ml� ��T�?��!BH�6y��X���S)M@��3�1��5��p5��8������c�i3�W�&��s�M�\׎X[6`����`%(��ܑ��	7a�y+�+�Cm�d���K�������Q\hit��H��d(�(O����&�RRpAF�&ذ1��	� #������^�B�d>�$)��	�j�.�2 �D>%Ӥ	V�$+������-�T�Zw	����� )֎�RN�O� 	��$�� eH�a�BX�-k�$(�z
0F5�T��a&M�R��Uf%��m�|��C�o�x�ޤe[~�';Ĩ��'Jæ�&P�wx�����4(a�!�e"��V.�@�f�:I�2�ۂ[%�eJ�b_qf�aA�*e�5�5�ߧT-��'0Uò�ڴ9Nur��ët[����D�q]�P��ԧp
>�j�%�.I�p(W%�7?X]2�`C*��'��=!�g��p�v���^�:�"�,�&r�+7��N�����#��a��1	�g@:v�l)���8�
V��� Ŏ�*�����\0:W���B,X����@�+̈́2RazlVq;B���[>�bѰ��%-qz�"��ĚLתِ���� T��W撚P��i0�ܚQ�1�����˜Ϻ���9�����޺H%>��v#�q��t�j)vEu�|٧#�?q�\Lw�G�g_B�R��|����G�"l_h<B&��MS����M��H�����e�N�=2��>��e�aHX�Y_�q�Ġ��-�$�"('����I�a&d�R l9��i��� 6	g 8D��`͐-D�:�)O`���'�M�q�Sy{j��AL,f��]R$�.(M��'�u�\�@h&M���}|`�<���
xu@h�6��1O�6E�$Ǉh1V�ȧ�E�iZD �4/R�zEfT���ċxvD\���D3L�:E�g$f�p�8��I8)��eӯt
�����@� ����bAJ� _�� �i;�l��6 � ZD�U��.s�c���e���s�'qٔ�j� A>b@fl 8��d2�y�8�_w �F�M�^|6��	4���W��;E�ʌ�����O>9�H7)*��ZG�7~��Qq���!6i�\�"O�tg�\�GC�;� �P/�6*~ȳ�
=8L�l�Ц�[�&�x\Pq��q��I8n\�畟�y����$��T
]����n���=���H���I���I�b�90.�2����J�]��¤��M�D���R2��8j��a�M��0�(err���,v���'܂�C��-�(�Ґ�&`��ʂ��=6Xl:K��@�Q�*d��[�@'�o��
S<���O�Y��s�$�0e�m��aS-N���@�Ο��<!���8:J5qQ�=��`b���a�` �Q�^�n�$��B��(�F!'�]�A�;/]X��O���6O�!!���~6-¶'X^qI����o}#W�_�H����F��x��!ڑ/���{���5����X�,��i����4�ާ_^U
'�>7K�8bg�^O��uJ�i��t���A�X�ӳ)�����D�Nxb���'9�qS�Ǌ;Ω�����z�f�&˓1.n�����;hl�t���Wm3�(I�9ƽ��N4y�l1���2�ȍ�񈟱_�!�$�M�t4��	fn;��S��H��Hq7#�b�ҹۉ��0�𕱃��)� ���� iR1K�i�;y���L#ܴLsp�T00��ѳG����!mK4aDcI�!,�����T�$�!���6�Br�8M�NMA���T&�i��+�8�bB�9!���#&a0%���[(���`�H7�%!�F ���Q*_($�����%e2-�;l�t��WJ��|gbIJU�E$$����(}`z�@��x�kʖS����f@�J�ⱐ�`[��\qu��bغ�
��R���XTb�N1�ϟ;�(�HUk��!h^EQ�핐���� 	��V���8�F��`�H!�aϞ9�8�xݴf���%+�0���ȟ�vYF(Rv.Y��P�1�ءx��!# `�ݚuK��:�=�7�3wYN<rFA\.j�>	�%#=�!�#��-Z'�q�&�`\�<B�C�#;9����ۅi�0!�E+�	�G����C&3o���R�3��F��{.8l:��(.v�x��k��7��$5m���" 0�ܙv@�{)x `+�'�����7v�h5K�ƒ��91��J�'Ҙq %I�(���;7Y3n1�,���ܽK���B. ��n�&�5X��ѫ�@θ.�������o6h����IW�LX9y���.U��utEG(? ��cŬ�r�;A'AW~"Ƈ�Z#��p��� *������ qet��5[�v/�8�B�
�/���� ��^�5��:Aְ�H� �<�p��	V莈;�!+	�����N�[�uNI;EƐ����!�� �lI`��x��%a#*�t�Q� ��|�G)7��)AG_# �ta ��0x��5Isʛ�w�)!" 
� ���iF��1���A�G�6hV�R��Y�g�& "�ʈ�a�b1S���9���"��'��S�e��_ʈ�ВK
x�XaP��ٌ)�(8���I0�����2̇]
p�c$J��@��HA.i:��ʔl�(�s��;#@\�Ë�I��ɹ1�"�I�a�����a�{+� abZ�^f ��)9����#T^������`EF��`�j�ѴG��}c�
�\bi�	F��u
zݙԮ�{Mz�R�	�j�����$j�I�+\��'L"��I�T��� U�V�A�BRJ�D` �}�{�k�%2�R!(�㐠H�`'2��U2CoP0)�d��4�Y7E,u���E �E���&��cPI1G����c��l�Iñ9�Lzs�Q�pm4�&�Nt�'7�%[�G��?�cG�M!�H�y�4�D/^�b�֑kv&�L!>��G	��D���]�dd�(�?��U+&�����Hp.@Y�����ia5"��i첵ۄBd=��#�l�S((�ΧKs4p�C�= ��I!�g�r�EF\�s�U����Z��Y���[g�aGxr�̸n�>�˶��26���L�-�� �Țr�T�PC�$[�T�B��1d��mXǨ3�4i�%A�/��;��p�R�HcN��|�;fE$�C�k�h� �;Eq�&��9���r���u�&~-&TG����1qB��k�$�4�p�y��-H(7DK�WD�AS��`���O@��SdZ�2�j���>�GG\ r�<Yr�[�O'Q ���{�)r��B'����Ѕ@�E�|�DBP�Dv�i��',k��Qs"J@�Г�O�`@K��haތ���R�Q2�(���{�@��(��dK�E۱c3�HRQ \[�ƭ��δ!V�v#�$�5��h�)����H+
�C@+Q8YDErV�ѕg&��C��c7�hA��'$��sr��g?�tq�+��U1BE��B�)���	B�kT iѤ[-`�"(�W�^ U�F�~�	=h�����4k,���I�1^2��O�	Ö�@�]5����fX�H��P�^h\����,A)�M�m��T���A\�hpp*�!�@��۟ўt���A�W�.���a8�R���)^�Z���xyb
�
��O�b��s>�j�+7�Nи֍�^����V���fŅ�ɬBۢ�2��ʘ{E�U c��|�^�"�mʩˮ��wD�<qː6����,�w��q�Ta�n�U�|��'�t�AE,�w}���u7x��E#4�`��I?�~����-����|���H+"h��d�	4s_�s�P �!��XK�9�<,�|,��C`�!�d�V+и��[*{,�hFi	8@�!�D�,4A��n��� �B�O�L�!�Вy�m�*��L����^�N�!�Q2
���.�H�������2�!򤒾T�����r)y���M�!�� U��	@�&B:�Ĺ�RN�T�!�ov������~�еj�E�d�!���=�22�J'vj��Ӎ�>�!���NQ� �2�Ǐ[o�6l 7Kq!�Ȟw=��b�2|ob<����0d�!�D�-/�P���D��PGn�9z!�d�rP�=��ś=X���R�$b!�$�=&�n�a�4@r��<.��
�'r�rǯ��&�F�HѪ�?���	�'�p��E�a@�ŨeM�1�.Ɂ�'����P!ݔ2K�$j%���)��[	�'�@:W���� ���	[��9��'�8�Q�K�+��Ƞ�"��c�l��'�\�i�&\�I��t1���e��T�'�"���fK�[�2��a��f��"O�|2ϖ�}�=�gi@-����"O�0;�)��n��\۠葮m:`��R"O,�*��V� H�s�&��//�9��"O1r",>\� �[�FA�3B��2"O��⋱2��R�L7�Xi�"O~�k�R�-���1�"«y��9�"O���v��6��$�#�[%@�<q�A"O������؃����E��"O��aQ�Wj���#�[�~��t[�"O�����&U���%n��r`^0*p"OJ8h6�� �ण��Ҕg(XJ6"O�s kV	��Y��g��QG: �u"O����a��\b�� �8�t��6*O�����c��Œ�	ǀE��()�'ȴ�C�ێ.�t�8q��aY�;�' ��쁒2y����.A3[� ���� �Q��&�=N�Bh���R�.B�"Oj��5jO3>�T�aՏ�0.�v|��"OB�2j�JL6y�U�KVw���"OL�)fH �U9��b,�?zi> �B"O�G=^���u�>��y�"O�r�	#t�J  G?D�8�W"O���'�2��ZfO^&6L�w"O�53�X2{��\�RȎ.pֽ9t"O8	s��<�I�!��D�:)��]����G�qOQ>�)�%� Sٌ�W��
���GB7D��`R��]\n��$N�D�ڀ#� }�	����@A�Ԉ ���g�0�b�>Oi����e"�O���r�j�^pm_L(j�� n��4
,)B���	b&�0&�K /)B��%^�[��=Q �~'��r`Kb��"���I��	���3�9Jx
t"O�{�h%+K��VH#q���'��A�¤I�h��,"� _N?E��h�rhX|d�P� ����L!�DE	0��cP��q��E�R�Ƅi�\�����D!��܆*�~l��]?#=��b+7�\�`�S�l[5A�NX�t�檂�H�8�Qe����Ĝ�gH��A6��)%K�` F�j���C��ð7��Pa`D�#9�<2��'ғ?νd��PD�pRLQ��� QM�D˕�	<;�L9#b8G6B�	6���Sqؒ ��`��	�#j�6m�6w-�(;��jX$Rt-n0aG�\c��6-�5(���ϬP�z@@�"O�q� /	��Xك�޾\������7	��Qj<l��٣e�M-��S�S��c� I-(1!D��T�H%64
���<Oƀ o��M�a��%4��׿(!T
���x:Z�H�/�*�h��r� "�i���	�p=��e�0Q����D�b���2C,�tybꆓH<��J"�L1l�da���-�~��~1�f�7k����! ���7�N���͙��<�y�j>@m��-����[��;N��e���|�
\�j޺%o:��dj�=Ha�_w[X����IM�0�];��p��Ɛ� �(0��
�A���DP�G��Z����Εb��֪
J�����;;F(Ν��j��pdY<'2��<XG�T\�X}0J>1%��d�a�-��w*�Y��)@Y�'p,�Q0��Ӓ�J��k��Q�'ßD q�-K.n®�R�ӭ@�Z�+���SզȂ��*Pt0��y���*Qv2��'���KR����m��	H�J��	��'4n	H 蜴y��@�$��1k�������u�WI�4L��%�6��<%,~�!!i�&�Ĭ3.��z�
����7}rlܠX�N���%��d��X������X�^�`1�\���ѡꏺy��y��L�_���G�۟^�켛竘X�<0��?z��١uj;SIA�_�V�hY����=�5�s���p=yp�O+G�h��`G� ׍��?[��Q��#=��Y���w�֔��e[�Gx$�C@YA���(?]����������#d�FQۇ�R~��q� �>[�\1$���m�H�3jϕ5N �E��ֺIH˄�.�{ �AZ.%�P� �^��bMQ��z� ��B?�ŢU�h���W�`�T��3���wE����=�gH
*�yN^�}_0��)!~���*w\>Y0D�%z��1�ʝ���6�1w��"w�\���t�1ͅ�c'���*sS�Y��O˅�L��O���2�=
@�O��J�)s%�X�+�|����~��T Q��1V#���B/�	?
D�Wo��A�	բ�9,�h\@%��qW�I��!�=I�l0 QK92Ge=<O�d8`��UAm*F(���\Eǹi7�H8% %e����WO�!Rr��F�H�S IJ���>x��hP�E8k4�L(�Q$f�jsƘEZ��$14�����I�ve�u$��2tf\
cc�8O[��. M��bF��6M���W� &����$�)fv�U�4Z�}h���ڮ OƑJ'ڷO���@@��k�iט�A7b_�@��eA���U
F5��'�~	�u�˛gXܹr �I4jOި��O㶬a�����\��M;3�u;�� )XΤ	A'Y�;Ov��0c\�1��b�E��~�q�#;4�i����b��ظ��PYSfAyբ�'9z�QV��y[͑��T,,q�c��f��Ȉ��Q�]YpMa�b&9y�iJֈH��̦�ZL��o �60�f	6k��p�a�%lO�$�Vm�`��0�r��,jȡ����# M�HYʋ,��̢�&]9s�R�DI`�� ���O.g֑���Z#I�T��
�p���ɗ��>!���K�=����+<��X�b-e��Ц�ܧ3s�acU��E�|�p*ŨQ=4D��X5Vh�04�?	�H����ds�uS�Ɛ@�j�����*U7"tS&�'�
��G-ǎZڞq8��J�4���y�H�$�ɵ鑭z�x����Y y����R�\�ݺ�#�4j�^�[�H�}$^<*��E=mӦ�T=V��(�Ǣ!DQDH�P���l�ў��6M�=�U�G�T�� ��[8jْو3�^':u��P�箙���9�e����Q���X0�[�kߞ%��)V�x6*]�3 t.��[EϏ��vų7�REx����LzZd���p`�D{��N��`��G��sL�Y��	6SW��D�-�+/s�X�u�H�Rxz�z�L�.4��$!A�:_�az+W�Af��H����bNT��#�Fw��y2�h
8|�,'���]�|�7i&1��X� ��
vF�O�$�1��8[���``,�?�� �{f*���B��o����
Q̓n���ujN�V��B�+~�6)]3_���(j��@Ѐ����B׉"2���V�ζ�����.q������*o��dG{
� r�!������@�_�.��X')"٠�x��Ow��K��Kr�j)��mڏ	�����޿#���)��ň����Q��ݢ/�=N��Ja��bL�#�/_mx�d@�%�~�T���i��s��a;D$1R\��Ŭ���)�K�5EGU8�@E��W8n�� f5b耇�,g��2$l 0a'tI��Ɇ~� [�L�YU�<�% N�Y��q�p��0��AZ���(��oZ�F�'&��	��7K�X+�FֻM!���3�ݟ�8Q-�k�q��K��2ȫ�:��s���s-�i�nTp��J>XQ�pA�:�V��jk,��Đ�*@� J3���7���F��,C���$"0	(�2�o�o:�=A�Ά�'�FP0�nI&<��S6��E�f\Q�D"�p�ӎ��c���TN� �^|x�.H�:��3�i����b�Z�eD�ө� G����V��Bڸ� цD�0�ax"m6{v��D�
���T�/���բ	,P�pt�p�,K��ɲ�/3\)��U,G7�ŢL�4��
h �eɘ�g�bx�%ЫR�B [5���O��ylҰU����6+!U���h�
ؙ�([��}}��S%
�@��4+�'P�H�4\KWllӮ\�4�ߘef�2ڴ��!c#-��{c,��EL21�Э�O�a( ��*H�����N�z'���؆ �"����i��@�Q,<̂m8��J��0�+��.�CYʢ�r%U?(��[�		�`
��iX���1�2t�*Ip�c@�J�jeХ�h�'t�QDՠL�ۿs��!��Gru@p(�Mˇ;��Kǩ_⦁���O�	-�}��G�z�6�kT��8���2n���3l���uZà �*� ��+�1�nt��lݥ0���Q����9䎚7�.��+v��11N�B�)	s�ӏ9S�r�N����9�.[�1�"���%A�r��qA�+c�̬ѷ�C�2|�I�R�5�O��tg�����b#F^�
���	�f�Lw� p���/v�$����؁v�RQˤ�x-u#0I�-n�[��=}���_��q,@9N��U�֌B�m4��E�L�0ލ#�"�V��	����%�񁀣� X}8u)�?�0h�q�Q5؅#�bԅT����
$���� \�"|Bᗑu,He�T
�� 5���C�p`1	g�U�L�ʬ��AS�_�6P*�AVS�x��y�'Nqs�!:��M�I�I�ߕ6{�@a�'�D#�4���&{��UiC'ty�=:�b͠I�]�w1�V�ð�\�V_����X7�f j��:�܅S����(O����ٜ2�|423�E�8�\1�aɖ�Ը!WL��v���C�v�(0/�q�tA���N9�Z��V��Ȝa�ׄ{p���s�TPB� e��P��RcI��m�<1�>�R�[)K�T}h1B�+7�d���L'(����(��xH�� }$���O#N
�B0�`Ͻi8�ɀ*�<x�*��h����6#���j���(�<� d�;2^q�&N�t���隺�� 0p�h����lλ;�������7Vy�N|Z�a�� l����v;�D���U4_�P��(:n�c�#ɖ_7Je�q�ͧw�-�rC�s0�p�E�4�	'.V$�(��IU^���}��@���B��D���優R?X�׬	�.T&�8
��\�r5㔜ŖP��e��<��]�Ϗ��q&�&=�3*����� q�9�(O�1��'%:�Cj^�� 25�_�nR�@�q"ՠh�5C!�ӣV6�ˆE�6�%i�1�����	��Qӂ�[�Qxcϙʺk`k�"/�Y�7�SCEI�e@�z�'��r�`��GT��D�Ϥ(��(��K@(tjAH��=?z}9���:�x�
J?�$$�sCW�Q:����>9��?}Cw�R+TٺÑ� {B}�e��Sf�)�C�2 ll$��?[P�o�5�`@p�F�i��Җ����� PcL��|�&���kw��
�\!+�^���D	AD HYt����w(�+>� ␐U�A��ٙu���BQ�#�I�j�R4Ȃ�
H�^��K�IZ0���.D/��̨dM�>#��=���S�k�X(�"k�N�B�[�+�H^:��6��s�\ɓ�<VNtA��	&
����@�ϗ8���Sŀ�W��D����&w�(��T�EO��`e���bVTuJG�S<5V\24䛏T5��!v�i�j}nU�9�Fct}�AA����ܚ#�һv���S�%�ԛ��d��{Q����'� �a�ѓ;F"T�J�^y0��	�K~�h�7SЄY��k� ��R��Od��V�˙7�DI��?-��kFm&��Qs��6;,� O���|㵃�i�`��_��xQ����9:a-� g`��B*���fK!�*(̧U'6��H�d��D�x4��!K̳[u���>H���'c�ղ�NȦ}:�EFy��R;	�ux�kY�4�h��)n�4�� �@�ty�e��������
�}$��\�8�h�
�럸��lK�u��) 0b	Tzx�x@��'�M#�Δ7D"=! �V|v�@ +��`ʴJ���T2d��q�Y�D��� N�#d�$	��ש��q(DN���j�+����X�A������g��hF�!f  Q�m��H%T�GC���I&\��C�m�h,9RF@�$ޚ)��"�|>ֽ�F�'|�(�TH�oAb�˃�́&g,q�G��H��9�I<=L� (���Xw���I�2��r5FP�w|��2�RZّE�1�L�9T�]B��T��D�X��k��ԛD������4DR��Ilӆ �6dC�g`Ja�& �qy�*��kJ&HSF�Q�XK��2b�*�()�=!��IPC���B�t(+�-
C���sbH�6cToF0d�,� �X��ThC@����ٓ0�������k9F�yd"ђ�ay�A�t�f��#h�� )c�bF4$�δYw���g�`�ׇ�u��X{��w�iJ��I7|x�U(Gﭟ��'�S�0F�իC�C�yj�5m`]���լH_P=+7��#P`�O��R&n��A�ވ���
�:��e1s�
�c��:��L-Ǵ�k��dc�����$*�|�û ��qI6����M����H��U��ݺ,�����KS���ɻ>7OI6Y/t�0�hR(fS0a.N묡�w�Z��bXt�Բ-�"	��Z:}B��R�k� F�H%����D಑�D��i�y�%"�_c���]&g���`f�Y%8=�]"�P��S2~�q ��I�l�6����J���)�$u�G�¡[�ʄ���A�=�xEZ7)�|�><�5�L8J��I�t�����I�!X��y�̕�q�Hic �dP�@7�5i�T��	�q�B)�`PaY��hw�]�j�Xa!阔7p��l��\y�E9�H����[?x�3��Zw�yI$H���Q	�A�uW�W�h[�%D2f"����Η6��a[��ґ.�OD)��FW�'U�A	��ăy�Ĺr�U�kfbeR�g�B8���s�r�2�i�cPP�&�B�q�~L@�
/c�|Kvĥi2�8n�u�j�
�)Ƴa^pڦ�Cr�F	�!��Y�r�MD�L�t����<!2J��(���yĭE�G�:��a��%��U��L�C�P�@D��?�4)�c��tĺ-��ؿ3���D0��SWl{	x",� f(���I�d��9��}��@ʳY��H4���vXZ�[3�K>�4����D��!'%�6��[�O�_��xD��uZF�K`>�� �t8C���G��d9FKI�2ca� ��5�]9�͏�'���G�3_@�YC��`q(�QAG#z���bl�_��c��kp8�a狻+�L)��!�8go�0ɮ��a	�J-
L�={3G	�2�xe��>9\�mbWmGވJF�x~��V='Ҝ�IU��t� ��7��O�d�"��U�8�3���-|�$E�Eo|?`U)�Y�<��U3�O�$[�:Ĩg#��4�U�cI_�t�.Q�5��:dY1�Ù�8��us���%X|� ��S7�!��AG:����G���)U���yx(���Zm{� �銜S5�5�ׁG�;����G[�F�(E0Ŭ	� ���ꔩ18�p�ŋ�T���� AA+n�T�rS�J4[�<mxELIIܓZ�<�#�;{���9��ɰd'�ъ��X�z7���7���Fl� SF�-H�-�wc9���!&�2a.���T�Y�?��� �	:�`���M�� �"ҍ]�м��؆�����i��$X��m�:TH���-��ݩ��Q*S0�!�WG�6z�څl�79Q��
�?"��d�ƿ6RH�t-�1�@����<9����^wX8i���s|��3�K�&FqrpeLp~���E ��$�K�e��D�4.�ﺓ�eƓ�<1�"֟�צA�\�� �ʛ#�lM"𩐙rk��!E� 1��)�h֦���;kvdqG.e���)��K����	�X��*bJ�qXE 0�!C���u�+!��<�}"G��[S��ӯ���BN��S�6pYTIы.��Z p���ze.��@��@���,������8^�pP����!�����oV"�&D���M�&u@��Z>�b%R!ςY�vL��O�����#�6d�UG�"��CV��}@6���f�)Q�8�o��f��ҏ�ֱB��L�'O;^�\Ib�_a�d5��ȀZ�|��ٙbE.�Q+	%�<�P�����a�ҋ�n-���H^�p	��Y���wPzA��	�s�0��/3�L<YQ`,Tp�[�h�-q4 ���r:��T�L��:��$.�$f�
�CްM�Јh�oR,H�`��6���$��	� ͒�NAf}R�T�-�paɩuv|���ˊ8)o^��R������	<���ۊ�t�W?������OP��͏L>N�Ro�>�X�P%!S��4�ģ��T�p ��5Oꐂ�`�=��<���W�qjՙ�� 
h�+P/N�n�r�;��Q9�H�@����i�#:s��d�A�-H�XE��.î��V��m�b��ϓ/�������i�l����d���J�-�1c�����̘�l�@��V�,eݾsvO�Ü��FlT�jUQ?��E&m� 8�d�<(�����X���'����̘|�Rp�N�S�O�*`�e��'̬���;[<�A趎�O|��0bLJ'Р��#��������t���D�E��h��3�JM�A.L��N�sr��~bĠ�0���2<�б���ؽrj|�R'�T���1۳/=�O=�v���~���3D�!F��Q����l����']?8B�ɲG���F�T��!�` ���+"d�i�`���=)R&��g��h�f- ��Zۘ��`���7��a��Un����̈́��S�OM�
��	9~� E���w%���'��%3 NL�1������k��MR�'%Z��&��к���K�`�jP��'d�4(�(T�j �b�؀[���3�'�
���l����	��«{�hb�'D4`X�꙱}4M��p�Н��'�>��%���SN��P@
;r�t�K�'?>�Y��N�_�������s�� �'~P��M	�rZ��P�r�@k
�'▭8�ǔ�=��P�����-B	�'	�WF�:���դK>B`�*u�%D���G�H�NT �`ږ1��Y�u�!D�X� ,�M��=��C��-�yj�A=D�(31iƛ]�R�1�� ��ӆH$D��yC��W��]AD�����J#"D�и6��S��J�M$x�����&D�`��"Β��4Q�fU[�H�de)D�D�A��6AP���Ϫ[q���F'D�(�dˇ*�A  �5F�$ta�l"D�|���/;!N� Ԍ�����E:D��a�f�0;�%�r�Kk|�0x7<D���mJ�`TxI�KI�x�U�'D�xbd'1GWʜ�`�ҩ}�r #��"D�d��Ú6@6 ���׌1X��x��!D� i�o
v����u���ufB�# �>LOr�B���4.�-x��zl3��1�^Ĩ�l� �r��$��V�2="vNE %cQ>%RiAZ�}x@���:��sE���	�7�p����Z>�
D��+�r-��Cө��堣-�<���V�M�4��v~��i��G�xtpbK�z�0��B��ɭM_�ū�4A��R'�c�OҒW�0��P���ۿ��0���O�+�OME}r�	ma��͜?N�5�#W�5'n ���������T��1ac`��$?��|ڒ��4eP 8��"�
Q� N�$�����yReC�=�a��JQ��m��/е!����eL��y���<r`�^�)�AVA*Qh�<5(r�H`M�d5ln��<��&��S�π z�0�eTr��L�y�8O��PV7}"�1�'F��O	�O�*�!gL (��YJ�k�����>� *�Oa�4i� A
�iE��NY��Tֿ�� �V���%��yZ����O�ɟ�|���
r:�P@"¤$��Ex}��'$7��!��)�'G0�ش��\�~4����!0<%o�ß�s�4�`<��ܴ\籟�a�4�S�Ǣ��\#�P11O>3aJa�S�O�F-�q+�9�U��
�%
ɰ�Z�L��`b�"~b�'P(`�DW7c�����L*���dŰ�0|Q�F����^�z 
��k�Ve��x���Jk��|�'�V��Q�N��
D8Tn
�{j�,�M��`�<�S����La��NL(�u-ТRBP;�'IB���y��霺ZJ,�z���q�DI�ơ88�έ���2�I���O␍&?5
�	�.��1 ��}�}�p�c?a֯i�����0|2@�hÄ���;Q��;�0�M;��<��'��韆 ���)Ҁ[X�9p��_�ry����l��?f 	����C?���<g��c����<��#W�^�+T"��r���#S�
'ʤ8z��U<B$�~�M_�%n~,c��]Z0
Q��$�ybl�7|h��PHVDh�؋0
���y��YfT���c�=��5B�	F��yB&3dV@0�"���ȗo���y�@� ꨕ;�n[�x�^�a�
�ygnII�,ӷB�PUK�<'^.�ȓ6��� �d�"6Nܚ�*�O[Ɇ�^ d�9�ȥK�>��_�Rvj4�ȓ���G�8B��q0�	���28��FTi��Ň�VH��bG�Ǯ�*͆�)�����.�;���Ңo�<��h�ȓK�)�e��*��6��Ą�R���KF�\w�峵O�,u��h�ȓC�(���鏝A��i3�i(R<�ȓ'�"�E\��!��J��H��6�"��c@V/^���R&J�:�2`�ȓ
�R�h��_y�؍�5^��FT�ȓT}�p�Sk��@K�����NG����w,�8���V2H�|M���6)4�ȓ}$�,+���;��]�3M�6Ui�D��40�+�iӡq��<�e��)6{lɄȓ
"`��bL��t��ѝ$�.�ȓv7> ���j�5��	�51jՅȓ�t�3턓o��ce��7]�����x��-�1 a8Ec�/�(F*�ȓU�HMj�	X�=�	w`W"U����ȓg�<[�N֚(�X09���Y�4����K4��/O��Z�M͉E���ȓLȀ�����Bq��8fG�8w�<�ȓD��XAM
�_!:`��Ǆ$Qn���fDy26�R
��d�g��L.݇ȓB�z &�>ڂx����w��,��l?��0�-�wC\U�%h�2
 D�ȓglMsf��>y�4�a��[���x��a��̐Rtq�(I� h��&������V�]��5��d>0���b�ZHY惛8]������ ��|�ȓV���1���*jnܒ�dO�q�E�ȓ�^��Q-rt*D��K�t��+0��X��=
$6��h^%��ȓz�H��@l�	jϚ�R �Ф,\Ʉȓi�ɑe��UҠ�a�ըZo�t��}y�,���K�w�z�p�@ƥ<� Q��x낰��J@�bSx��땻?���l)�d�5�ή	O�aB�0nj}��3�p�Za�0F�ش�7k�e�攆ȓ-q�a-�1�������y���ȓq&z� ���}!:�{�H��u�t��S�? D��&��:#�I�.�9Ϣ��"O����ū2�6�;1��<�.�q�"O��ѡX��&YY �ƶ$�R�Z�"O��"�@�|ST	H�M�9&�޼h�"O8���G��y&�`mN�l��E�p"O��JWE�/��ʖ�C�
�@�b"O���e��:=���4,�M��%C "O��	A�N�sz�h� �?I��i3"O�̩���6P2��l[	h(��c"ONX(�T%!o��A�IJ�7��T"OhDҵ,�!S���3�L(z���"Ov�e�V����uŞ\ilxx!"Oh�R�UqE"�wV�Kgh�"O���CkU�g4\Ucݴ<�Y�`"O|����
o-98䁅)}��
�"Oư��j�D�v�Rp \�+~�q��"O��*��Q�Qv��]T��"O�5�B��:4�֌ARW[~��r"O|$�� #b���s�Yx���"O<ٶaЩn/ �	�kƃ]�z8�T"O(��CؠŰ,G ���xP6"O�<���������E�v�0"O@������F�ɓnƣM��)�"OԈ�T�F�pn����D�J��8�s"OJ��ԖKXȹ�U�&�B"O��#S,�/$>�b���/C��=�E"Oބ!0dġ[�ڤ1�i�{t�{W"OPD`���~�%�B9C���G"O�C�P�`^̲���W���d"O	jB ��j�U����N�iS�"O�6-OW7RݹBk�#Um��RR�+D�0sɔ5�^t�G�o�t��+D�t����#`Jq�d�jОH��G*D�8H�)҄R^lٖ�ʚ@�X3w�&D��V"څLchD���Hp�1�w�7D��JAJZ�Ix䣐�Ć�N��:D��󂉃U[��˄�"A
W�7D�<�C놁}�i	��J�&��"��7D��{R�*;�h�V�G�B�ï9D�B!��1})V܊d�+¸��4�6D�Ԭ]$%���q��C�h��3D��*	>NJX����d�*�e1D����;*��"�k�:�(�s�1D���$��YAf!��+-	�Uʠ�<D�`:��)[��س�ʙ1T�m$H&D�ȩrN�,Q���Ȍ`�X�q�#D��XmN�D`���/Y� `�d D�x#��|8X�a���>�ȥy��8D����y��5k�%� cv�u�gd2D�����w��T����3��"7<D�4k#�)�����Y-k���"�8D��[���8tB4Ыr�W�c|X��$4D��p.�!L��bB/���yz��6D�l����)��2H�r��eX��?D�`!4�¦��yrDʓ�YuT]s�C=D�H4��9#
|��"������k<D�\����l��³EC�Ŋ�� �8D�( �፠D!��W�(	ghH�E�4D�d�!�ҐL���@�J�u���K�j1D�����=4JV����		K��Ic�-D�x�UΗ=_*\��p�I�[Sz���,D���d�]!*�>|Yg��vI��*D���fI��JE��8o`E�aH+T��di��g9
�QF%��i��z�"O� ������;o��3���3�fH��"OH�r�I.bԉ���@�~�Xd��"O24ۢD�����9���>Z��%�v"O4�SM�hH��9a�5,}ҕQs"OlwĊ�\zX�AE& ���&"O00�%;E�	��� 2�V��C"O�M�z�Má���v�`7"O�U*6@�_�d���N��6|"�"OZp�S%Ǣ2�P�ϊ�A�vpP�"O�D����'��i�P�J(uf ��"O.e� =;2���E�Q����"Ot�2���Q��uŉ. >��!"O�!�2� �8%��s g�* >`�&"O�L0c����q�� ���QF"O�1��n��a4h��/�![
D0P�"Ov��6_󘥈�M�6$q@e"OH����lM0!p���T�Bg"Oz�4[3}�X�X�(��]a���"O�x��-<�C�❸HxtՉ"O�%9�a��>���k�a%0�ڭ�t"O\d����5O��!�� ۊi��("O*��īW
�%h��á[�&P��"OPt�3���QK<�pe�_u�P�S�"O�,�t�ηFT��X���m�hĺ�"O~)��iBxuR���I��k���"E"O� p��֎Av,}�H��O��l�"O.m+��Ĩ.Z
��h�V��x�2"O�UGᄰD2J�bdhX���i�"Oִr&�h��	 G�%Ш%"O�THפ��K~�r$�Z2g�"5"O葙�EF�O�&��E�3�� "O ��Q%�0bH�A���B�"�t6"O8�0f̎
Uh�<Zc��#D����"O���f�5c~H�҅��$x�\935"O��C6�TT� "��i�H�$R�yF�4z6}�[xBn@B��^�yRCS=vP^!ތh(2����yb��4Cֺ�
T��)Y>1
1���y"���X1x��H׽3�x�P��y�JY�bb� � U9X0h #Af��yB�Ǵ&r\a�J�&]Qfq{�$ɓ�y�o�,~�t��P���Glؼ�yB��D��h����8|8Գ����y���6V�`�''�@���P��y"�݇i���Y�c��l�A0�����y¢�;`0��a
�w̄���HG$�yR���\l��2��l5~e:`ǌ9�y�e�3,�l��� P*_�� �t$Ѻ�yZa	� ��D�QPi�L�y����$��t�׫H9HCD4)>�yBO4J���3%��v8V}�Rj�0�y���� OҜr}�4�Ō�0�y�L�
B򂄨�Ïm�E�d��y2FDS\����rLI�OG��yb'�1xT^���E��8��!�� V�y��0c~��	<C�n�K��C��y���%3ǜQ+ R9qT�P�1�,�yR��35��H��E�$By������y���,���)磏�Y�e��y��Ӝl
�H�(�����A!Q�y���Sd9bFҳn�å����y2 J�Y2~�!�W;v@[�����yR(��`���p���>��1	L��yb��;��F/�3iƕ�pG�y
� ���&��.��h��E�J�BC"O�a�-#F��ףʃB�&��"O�ܒ������0dJ<=�F�;@"O�	qCL@NR ��>�40�"O.�Sa.�*�ڬ�e���Z���Y'"O�QO
hz���0  �/���b�"O٫s۱j6n��C.�/�Ƶ �"O�T��ъU�
��73p�"O���@4v�H!;�퓾j"��5"OԠ`��*H�0p�M�.
g2u��"O��p�,�gC\�^a��+��U�y-�Y�P�i���\�ҼBf���y�ޤN38H�7鐫`K����Ҽ�y�I*� � ?]�f���j��yR睨�:`,I�[��	���yՓ;������1[�*�Ջ
%�y2��R� 8iaFY�<�T���a�!�yBi�$�Z�	R�H�`�`#�Ĳ�y�B �PU�8�0 ގM���q�G�3�yrA�y�zH��J4F����ʞ�y�F�8) `  ��   �  {  �  W  #+  �6  �B  N  NZ  .f  �q  
}  m�  Ս  �  5�  ��  ѫ  �  V�  ��  ��  ��  �  ]�  ��  C�  ��  ��  (�  j�  � � P � !! �) C0 o8 �@ �G �M .T �Y  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t����	V�Oa@�H���*\�L� �'��O�x`	�'�6%� �6.h��B70xġ��'�؝!� �>"VB�$�*6�����'���vB
*%���׫�+:VP���'z��gn\tF�`�#
����'��U�bM���2g��Z�i�'(f���A�*4�� �6gV;�P�[瓨ēG��TN��!���0S�B���ԅ�Rj.�Z�����{�!X"��>9+Oj�=�;#o�h4oS�/>~�a�NTG~��s1�4X�H�iX��AAR}Z5��{��h�����%~"cw� ,Gv\�&D�a#!�dǐ*`P5��+MJ
�� F�,�C�ɧ� @#*Qg���җ��N-l��D�O��O"T����<����kY�@W�Q��"O�	P�Ȃ)>����>60�g���>A��� Jp�eS�.ͽ6�@QB�S!��ˌ��PnL���/,!�$��u��}@cm]&'<I� ��D�!�$!!�>��iگ� }�ш�m� ����#r	OJ(�@�ӫN!6z�@�ȓ\�� k���o#��"�c�f�Z��ȓ	��mR���Rr<917��B^�X��.'a�'}8-�� ���T��1g��:�j4S
�'���g\ x�h����*"x6�a�}��i������U�E<"\h� '�
 dh�"O�P!��"�g�X-ga���5�F8��Ѡ�LS`�2ԯ�:W���.)D��� ��,jH�T�G� <r�sW���M�����>�7у���Q摥d;x@�E��E؟���ݠ�l�0���&K��8=���iЬpk�Ō7�z]�qfP0T��x��|��$�E@\�/�����/z�ع��l���I����cn�# ,++�(�'�ў"}��J��]1�U
��t�H�����[�<�R&�5[�p�e��h�r��pE�W�<�ȉ�O�P�Q�];2z���N�<�adM�V�"�Hc��ْ(	*�B�<I�'�,_K�M��ЕB~>]y�`�}�<q��Ω
&��
�阕B�m��C|�<q�k�v����M��p>|sp��z�<ٷGPH@I�j�1�Q���Q�<qd�җf%F�B� 
��H��TH�<�ǭP��\X �@��-����Lm�<�󋉩Z�8�ID͚jx0��q�<Ѱ�^[;f� Wh�Z2��k��Bq�<��jڰzp�x2�N2Crf��&
�Q�<�G�U!\F���T�� ɣ��[K�<� ��$)H0[r$��$�5O���p"O6����jDY��&#܂LYg"O�L��N�e���E�r#���A"O�2�Ԙg�&P�b#�Q�Yq�"O~�W�D�8�cqKŐJ�t��"O��`do�
�|�b(��i�6"O���$�B��) �g7��azt"O2�	F�;-���1��	�+z5�3"Od�j�捼`�fMBQ"��m\�)��"O�p��F������G/�9O��"OF��Áĭ?�u����+:>��"OĤ�̤V��M�T��:�"OȰ��Ĉh�� a�I	T>��@"Ou�jԯ0& ���*ο�~8s�"OD�#/�!�8q���ֹP��q�"Ot(��N
0-�`Á�T	I�bP�"Oĺ'h0&��0�D
� �Z��"O5���Ie��m#���(\�J]є"O5��C�"whR�a��˨&��ّ"O���Y�w��䃡�?=�T�v"O.83�پ�I3&Aƀ*̆1�"O���sC�&uj�;u A2L��:D"O����W�1�y)PO��,��a��"O����A :G�Z�˙4Wd�"t"O�8Y���`W�@S��ی��U�c"O  �S@Gt�8�(�&����"O8|�
5���ݧd�0�S"O�y����=�f-	�NH�]��I�g"O9*�NR�SF6����kV(���"O�IX�j^3iJ5��lK�e`�m�u"O� �vk��rukR�$'F�a�"O��#�L�#S�ٻ4
��$��P�"O�Y��:V�^d��O� E�hȠ"Oly8 
�P.Xi���OݬlKC"OB͹Wiڡo-�@`T�Ǝ|fPL��"O� �����8��C��6c���"O��"�O�9�����]���cE"O�����8���GG�@� �Ȃ"O`d��ˏjѸt˶�!h��:}!�d�	��\����]�L���#]!�F�o~�(ހb��H�����ax!�]�	L`]�ƅE�Jjl1�lWX<!�Ɓ ����'N~}3AJ�*(!�D=s����S�.�r�G��!!�DՓ��M���?I,)"�Q�Q!�D�P(�<B萆~G�W�N)aX!�D�:D����GH+1Nl� �
�/4A!��O�[A$`с�S8RE��b�!!�S0����i�2M���T�]�!�D�n<��膊�WQL	���<�!򤊙�`���ρG򜱇�O.�!�$IVU����i��p*�	ڒ\!��H?n=��m����%�Q	)F
!�D�H�� �iw"=!C$�� B�ɐ+K@U�	� � ՀcdR�fv�C��& ��ā�΀Z�ݜr��C�ɘ ���.F0RWH�2Ei�B䉷z̤P�L�V�4ik7\��C�I'�,�wC����9+gI�3��C��1`��"�ټo��sO]�v�C�uʂ�jq�'�$0�V'g�HB�Ɂ`LT@�M�`4̱���;a&B�	O�lI����*#�8��M���B��8)°���oA�D�J�XsnL�~ZC�)� �0��� /p}1`B��;I��X�"O2��d(B�n�PI!7a��'�l��E"OT+�
��Lz���d�|ip�"O21��!��G☨CCô��MC3"OH�I�C8iA�R���9�zA���'J��'4��'�T>�����	G����.��v%�do*v�I�|��䟴�	���	՟|���4���2�ٸ����J��@�
+H�$�I����ӟ��	�����T�I��H�	�D�J���r�X,A��A.�������	ԟ��	��(�	̟t�����I�����;K.;"��!hD�	ПT�	ޟ��՟�I���I��l�I�N�X���$~�M���/~	D%�	���������0�	ʟ�����3�, C� �3���s��
H(������I��Iӟ��ڟ ��� �	�x�DȘ�I������_6S?@��I˟��I�D��ޟ��Iɟ�������I�e�����Դq<PZ����X"@��I៼����P��ϟ$���I���Ʌ3o-��M�PC��xAY�d�� �	՟ �	Ο ��ӟD�������ß��:�6�A��L�8��)�3�أ<�4T�Iןp�I̟(��ğ`��՟��I�|���<���[!0���Ꝧs����؟`��ʟ|�IΟ���䟘�	���	7��\����s�UKp�ͯG���	ڟ$�����	���Aش�?��U;��#���7j��\�A�17
�Q�S���Iay���O n��E�$9!E��J\��!	3.�Y�2?�r�i%�O�9O)nZ׊}ٷ�
Q�����4�%{�4�?ac���M��O����m��	
B�H?Y1b�7)��儆�H�r�ZCI.��韤�'��>%�q�LI�]�g�O�{V�'����M��)�w���O��7=�D5hM��7�6��F�.a�����Dæ)x�4�y�[�b>�CFڦ)�(?�5�aB4/��؀�I�y�5͓:fy3q.�k�&8���4���d#,,��S>M��#�ߢwY��<9J>Ѹi��i��y�#F�S���0�iеWu`�dB58�OfY�'�6͋ঁ���DR�qD:4B��ّpp��qwc\>:Q�I�#A��#H±%�b>�ۃHM�2�'D���.����m�a�N5����TT�T�'���9O8��P���GH�`[��b; �h�9Or�l�lK|�,8���4��aq�N z�Bl�D
��*���8OlnZ8�M�����9:�4���1.ڬ�`OИ>7���u@�?~�1�&�T2�y��:��<�'�?����?1���?&�:F9h}����qւ{Bf\��d���M slӟ����D&?�I(�.�r�N� �� FҊ��q��O�al	�Ma�x�O����OJ�T��(�A��2JR� f/]'S�ۙ'��)�&E�2a����v �OZ�9+O�0�#��rwh\hŗ��Ug��/�?9���?)��?ͧ��DΦ���۟����Y�
���
�"V��,$¡du����4��'�*�%���f�J�o7<�X�HPpÌQ4a��S���̦Γ�2l#C�&j:�@E���y��#3����d�F � �M�	��l�Ѧ8ۂ�ϓ�?y���?a���?����O��{�E�
\�F���J'=j.]*��'\2�' 6MI�H��˓n%��|BM$i7n�X��	�,&]���-3����us��|�ƋӾ�M;�'�����	�}Ab�ha	�<�\`�M�z��Tj3eB�5"��+O�rbi�<����?q��?9��ǀ ��4�F��'�N	�$�,�?�����$�æ!��c�ן�Iџ|�O
$yZ�̌<��iX hK�)�=��O�a�'7M��+K<�O$�})׭H+)4�AC��$Rr`ܔ{��R��"3��	�u�(���L}y�wET4㦆�!H�t�S��>�R��'u��'��O
��M㤣\!8;rTP&�S<�j1�w��3^��U����?�i��OJ��'<*7͍X��9W�@��K����m�M��K �M��O^y��=F�L����<ɔ��(�X,Y0��
�(���N��fU�(��Ɵ�IӟT�Iğ|�OX4)��	&�����H��{�v��`�O^���O����$�צ�?t�(�3�|�y%�_5l+*@R�4e��e?��)����7b�Tp�KL�\����X�s�Ȗ�`�8S@�׸xM	G$^Iy�la����?q��2¤�uڛ+�ʸ��ȿ= ����?A���?	+O"n�&c|��	ٟ��	�L"�|z�@�;E��d� ���*����ET}��c��hnZ��K���S	�. �����䂓����'c8�)�Y�$=X��EY��\w�������|]����)I�W.Hv��W@��z�4�I՟��	ퟠ�	S��yg�+.���j��i����DIS� {��a�\X 7l�O*��F�e�?ͻL��`�O�[�z����(�V����Ft��mڵ}J�l��<���H��
T(A�Jv�#��s���A��~ ���dC;��G��'a��'#b�'J��'TFl�e.Z:D,�zM��x���T�l�ٴx�҅���?i�����<��N
!���4��=KT&��5��2��ɇ�M� �i��O������[�r���A۝L�\-+��Q=Z��%�P�M�C��U�p#�MF��uGa�<qU�ie�2yJdR�gP,t�Ƌэ�l��	�����ϟ��i>�',7�B�S����Z4>�p��! �88�ɐ�+�,���̦u�?�TS�p)�4c���!g����p�H'^�	�ĭ�,y��r)8Mr�6�??Q�gF!u&h|�	���䧿�� xȁƠ�i)�9�C��]�^�;�7Oh�d�OJ���O(���O��?���αPFzkc�׿	H^���� ���(��4���ͧ�?��i��'��	��,xt}X�O�j@��(:�$E���4���ɀ;�Ms�'��j�2�����	�n��8ؤcӵ;C*YI���E���鶞|�Q���	۟p��ӟ�@��H���a�#x�Yt�Jɟd��Xy"�y�Zy�wI�O����O�ʧ&����9m�\Т-�:��'7��M���hpӬ�$���?)��e��l�\�:ɀ�3B(�Xš��XV[f�� ���TJ�%�ޝl�������$�I\X���=`/��!��ۉ�?��?���?�|�.O�4l��bu�E�@K�(Mܽ��7*�
Y��=?U�i��O̍�'�6MލwJ�%i�� ��T0�wŃ$kz��l���qh�ƦI��?A��ƲO�:�b�(�U~R#��wLr�Tj��;������y�T���ߟh�I֟(��ş �Of5"�J�#&�͡�,�8snakw�~���$�O����O2�����F��]���	�����z	��WO��5�4!3���!��)9�6�|����&W %-��ҥ�\����s�v��RR��T8M(AZ�Ny��'vRH؀ C���5�ŋK��9�v��$���'�2�'��	��M�����?1��?�g��4P	��<��Q�cT<��'ox�TR�Be�T$�虲�W�0!KE���<�[��/?A���1i�jh��D���'#�^��_w{��$�_��b!߈��!E�>y����O����O&�#ڧ�?w	@,�B��6d�5B��ѥ�ܣ�?)Ӿiq����'�b*r���杄l�+'V�te���*,ˀ���'u$6MZ���ٴF ��	ٴ��d��H�Hsq��7Q�挻��	��4��dΆ+X�I�F'�Į<����?���?����?�4�[�Ty$�z�ED�!�-A�`���OǦ�����I�8%?���0|��-���9T��5���ڒC,��OL�nZ#�MKb�x����(b�V�{d%����"JڋW,!��/E� i�~A"$a��St�|RY�4# لE� 3-Űb�Nų������I�� �	���Vy�kp��ز �O�Ⱥ��N�6U��C�A�>zZ�[�n�O|�m���=}����Mk�iaf7M�;M��� sfI�L�`@���`̳h���3��[�Т9:h�H~��;|6\÷��fla��Ժ5/�ϓ�?����?��?����O���)�X�B�
��Y�r�9���'���'�7�ǹ�����M�N>9�ዻ��ĀQ��9[>�Q�[�R�'�,6M�ݦ�S1A�>l�x~rh�;g�aj6-V�+B�2�n^_�0/��Z�nE�r�|b_�X�	�T����@��߉!w�3��A�Om�eB���8��cy���O��s�'���'��S)�.�
��M�	��Q�3�[�Ph�d�I6�M+W�i�ɧ�Isঅ)��^ ��Qj2n��f`�Ϗ�#?�������8Y� ��]��'���(��^<gr��D�¾l�´�D�'c��'T����O�I��M�u�ԇ}��`1.D ���j���a�^=�'V.7m!�Ʉ��dP�qp��,`�"����̉\"@y�ϐ��M{�9� ��ش�y��'��1 ���!~��O���R΀�u38a�j��Zab�t7O��?����?Q���?	���
�Am���dA@�h���#JFj�Hn������`�	U�s�Px���sժ��EV # �l���WBQ7����h��O1�Ri�a�y���	�QZ\R!���Y|�ݠ��	=7��-zzY�%�PY9��|Y����P
kٻ^�B�x'��5j+��&�2�'qB�'a�	��MK�g��<1���?i�Ğ Y�z�cEJOo��q�����'{��yϛ��tӪ�O8�bC��:l�آ����Hj2O��$�-FYL�`�m�.$�	�?�!�Tߺ#��'�V���CFĈ���� �a�s�'���'���'��>q�IV_�ȧ�N�7�r1���=9rA�I��Mk�\j~�Au�n���M#�=�Ǖyђ8z��6x.�ɣ�M��i���tt�6<O.���#\1
�1�.	�9��՛����B,S�@��
�i��=��<�|�<�%ʊ�k��Qr�O��m15�v~��d�\ɲaE�Ov�d�O��?��sA��@r��0�`�Y�Z��i�������]��4X���O��X��J�	;�49��ǂ�s�P��F	�ݙ�^�L9pHg��@O`��1M>����?���N�g`���W�?�����?����?����?ͧ��Dަ�@0�I�,�V*ّRX�U��c��$�AsŇ`yr�|��'K�0�Mc��i��7���8�Z&�k�����a�4��auӎ���4��[9v�8�IHay��Op�,N5�9Hҁ؜�f��7�
�y��'=��'�2�')B��ʤ4Z`̐Ԫ��_"z���h؁i�����O��Q��1�-v>��	�MSL>I&�{r����=X$�r1㓩e��'��6ͦ͝瓓ځoZE~�N
;�=P�N
�~��!���9��4"�R)�4�g�|BW�\��柼�Iٟ����	 O��Y�t��u�ڰy���D��jy�%q���Z�E�OZ�d�O�ʧ{��s$P9j���+�뛔q���'��Q��vkx��%��'Ƅ�p$țs��5p��W�^BP;��ͼ.�U�&I��4��Y��{�!xI>�6A�j(�8�b'\>�Lp�����?����?I��?�|B+O�UmZ�p��kM�$ z4)ϡu�����"~y�,q��$z�O��lZOO ��aW2��5�1�)y����4n��� V
|͛&6O"�d�6��� wiQ�KgH�S�? F}���3Y	����N?I�9�5?O˓�?9���?Y���?����	�{�|a��V� �l�HF��!S���m�9!Ԛ��I͟���t�s��
������)Q2-�fT�:�u@���9�&`Ӳ'�b>=�EJOꦉϓc����Q��<��
�k�?jIܩϓu�K�l��3�~��N>A/O��$�O��(Q�A�(�6L���]�rԸ�/�O���O@�D�<��i�&8�2���ݴ�?��7l��q��f�M�H�u�_�?�N>�{}�)t�>�m�$�ēRd�9봂��R��t��+Δp�̓�?Q�l��N��4��[���$��R#n�� ��20���R&��H�y���E~��P���?��?!��h���$�-�:��E�Ų"��g��J���ݦ�Q���wy�&v�T��݉S0� �ǃ��A����1��G_��	��M���i�|6��e?�6mj�8�	$�N5��C�PT���r�GsX��ᚊ5D$��6��\��Jy2�'Nb�'{b�'#��:`3!ڕ�I?_>V�g`V���M�K��?���?)H~�: ���/��~�t��b>J*$;�S����4/%��)���$M6%�!Nʪ��2Aj�>,�\��V+�#.��H�P��!�_��uwn*��<)q%� h�\r��]'���	�/�n�,�ܴH�\�
����|���X������C	a2�B�|؛����w}�#yӤ�m���MÄ �<溱���)fm����H�`ߴ��d��rGhX��F,j��8��Q)B�T���/G���;��O<�d5�O��	R�E)CI"y�b�2:��<ؠ��O\���O�9n���'j��|�X	l�� �γncȥ�#�>kr�OF�o�<�M�'k�ֵ`�4��D��6 ��h3%Ɯ�u1v�]�,����U�ψ'+nԁ�1�D�<i��� �#K��j���pe37�R��O�@oZ���<�	蟰�IQ��TwV�p��G�J,����ϸ��N}��o�~�n���S�$��5�\���G&Dh�U������S�<|� X�V��8� )��E'�'߄�+ �� �h�ԤY�}�$9��'�7�W�g�D��`.auA�F�D�S���O��妽�?)Y�<	ڴ�|40�'��9��H��Z[��,��iD�6-֢/yn7�,?1�'�r�Ty�BP���L�'GpA�ӌ�s$�$���7a��<	
�yr>L1�Gze�����H��+F�i�r]��'��'��alz�a���Ͽ�}����4,�#���M���i� O1���x�Go���0h����
(y6D��2]M��I0<��� ���%ZN&�Ĕ'���'F>��6M�
"���a
52���'���'X�R��"�4E�����?��T�����+W &\>�BJ�*M��`q��ͳ>���i��6-Hi≇l�r�9�/� ����%EبP���$$L��:��ɱJ~��N�$�u'��O�t��K�n�)���>'��5	��O�d�OV���O��}j��3���! ��rTF�`�4[��D��	S�"�'"�7-!�iޙ�Bg�܆��Q!��r6	x�P*ش#��dt�Դ�E��|�5�"m��-.0]H��2i�[-Hi��	U�6��Z�����D�O����O��D�O���J�;y�$b���$��	�,8)'��\��au"�'J��'̈q�&�Uǰ��gA���MS�H�>9ĵiV�7�Ty�)擜/;pq�EP#�����#Z���P3Z
��'L�aE���[��Ty��ƁY�}�K�6z� k�z>�'���'��OU��'�M��a��?!DO3*P�h��n�mPDi�$*G��?�`�ir�O�@�'��6M[��4F��ո e�Do`�s�IWȸ��H���M�Od]��únM"XYp8�I��R �����N����\.A�A��1O��d�OH�D�O���O��?�ʔG�#\qJ&�_����/����8�ڴ*��e8-O�=o�b�	J3��۷Ş�#ҾQ�� L�
��L<�D�i�&7=���ɦi�'[(�8�d^�t��B,�1m��Sac�s��ݨ#�˶-��'�����ܟ��	-���$%��st�T��4Ŋ���ğ��'�^6�Ò �"�d�O��$�|"G�5��i�B�
��8`�Sq~�A�>a7�i$7M�v�i>���&�V���
�pTt�FK��L�� ,�%/�VD8w��Wy��O ��r��^p%�tk�$c��E�B�pL���`*Tܟ�����@�I��b>U�'j7�_�rk�$�A�F^b�� � �<�2�i��O2��';7Btﮝ�E�:1���䎧
=�HlZ��MkB����MC�'P¯T-k5���Ȋ&u剘W��р��շ ��ᄍSN�Lyr�'Mr�'��'l2R>q�$�%pq�	!���(]Ф�����*�MSa厸�?)��?�L~�9y��w��P�i�	- ���Ɨ
'7�T��{Ӳ-mZ	���|��'��to��MÜ'(�����\�*���%���TX�',ʵ9� VN$q��|rR����������l�#'o��,IC��៰����Idy�)nӾH�7"�O,���O���eZE/X4`�"�
ww�ђm>��!��d�ߦ�1ش)�'OD���&[�^���� 랻&���J�''b)^.�T����;fM�I�?U��L�c��'� 0Q]0^@�ܦ,� r�'�2�'���'��>!�I�-BL:F+|�F�j�-G�/4$Q�	��M#��k~��k�l�����k�J�(S�$��m4�I�M�i�6m٘��6�+?9!$Ԏl�B��  V�? �@���*�\pi�FLs�G)�$�<�'�?���?y��?q�H���傀V�bՓcn�����ڦ!;�M���	��&?�I���t�#E|�,��g�2rZ��O`n�"�M�P�x�O���OD����w�`���R�5�V��e���;�S�O&��*�/"�z֝:�䓡�Z 	�|��̆�aa\y�*�L���$�O>��OP�4� ˓[؛FB���yBl�?t���c��G?08�����y"�~�(���O�am�#�M{&�i���@��2��uE�hךQ�6̕�!��3O��[3R��0�6FNJ:���?i�]�%q��JS"
�#Z@rB
U�F:��	���I�H�	�l�IO�'>�]��7�l[�MJ�lE����?9��,��V�����d��q%��P$a�	M�����<"��t9u����YC��t�(�)[�y6�7Mw�t��E�a"Ȑ�H^P�)�dU5[:��y͓w��!� EZ�IOy�O���'�L�s�,�t!�S�T�E�AC�R�'5��(�M7���<����?�,���`�I��-޼��B�ןguR�����lz�O҅m��M�M>�O?�4vU�$H:`�3E�3�:У�L�hM ��a��4��)8��c���J>Ѣ"	7M�Z�ˤ�˜*X"iƃ 	�?����?a��?�|R*OڰmZ��l�j��?cH¬�E.�?v����T�$?9�i��O���'1>7��Oq�c�m_��9aF�/8\�m���\��ӦM�'&�P����ܥ��YAJ��Z,�%��g@J�y63OR��?����?���?����i.,ޔ��j�3G�ś��l(H�oڀ2T��	�� ��g��� Q���;Sd^	B���aF84��9Z$F��%hӬ�O1�L��Izӎ���]; �5άd;�	E��ɽHl���ŷ :��%�`�'p2�'}B9A4�z2�0c��^�&qx}bQ�'���'��T�4��4II~!��?A��!���B�ԌSU"a��"F�O��y��	��M��i��'A~�H�'��F$���c�5X�� p�'2�AR*Q�!���	��?I8t���[ �'�`!��,��*y�!�tT�QH�w�'��'.2�'��>��	%+<�Za�G W��reH�X��e�ɡ�M+���?���h�f�4��<F�H�P����ҚY4�A�#=O�l#�M��@]��rٴ��D֚]%�x�jN2M����B��)f�Y�֠!f,�dA0���<���?���?Y��?��`��J�]QU�ݓU�������E(@/�ǟ�	ş�&?�	�z�Ʃ�¡�/5�pT@v��"���O��mZ5�M�H>�|��#�1Pjv-�0�����	S6��b�0��d�O52u��j�	N>�,O�YY`ŉ�;�vxZW"M<6��Q���O��D�O��$�O�<Ar�i���rG�'.�L�䑲T<٘W�M�p�X��'7+�	�����ۦ���������r#��*V�E�'U�!�%�K2�BP�ݴ�y��'��\���=�J���X����߱p�J�$Tt2Pʈ7e��9��,w���	�$�I۟�����P���\�-��x'Ǆ��Cg��<���?Qa�i�U��OT�m�K�_h�yxf���7��ɣ��L:KoPE$�Ȱߴ���Ol� ��i��Ɏ_P���DC7�,����6H������Q�~R�l�aȂQ�gy�O��'��FW=;�Qh��)N҈�蒃�9<��'���Mc��<i���?�)��m����k�F�s�P�4T�,kT�����OV%oڍ�M+I>�O��iP�g��]JT�܊KȒ�{��	�L�`��1��4���A�~�1�J>��ڽex�a�J!b��o�7�?����?���?�|/O�n&<��!�`_�.�0d���3_V��hg�(?���i��O�h�'��7m@�^�������A�b:͆�nZ؟`�`����'@p���D'?�<��  A�%Ġ�ֈb����! �A#;OL��?I���?��?����I�%Y� )j��
�vx��0�zEo+n�b�Iϟ��	c�s������t皏��06�7H"��,$ju��|Ӛ�O1�v�an�*�;�h1�QJ�E�X�t#�/��I���(
���/Jg��&�<����Sٟ��'�&	nXx�!C����&�ϟ�g�ԟ�K���My"�i�}p�!��?���͟�e@�5QD<�R`�����B��Q�Id}��ڴ�?�d�i�6mN�Z3��O�y[�#��!���犌����x�8O��DQ�%�vDQI΋���r5J:�u�h�O�!�#G]a�	fj
�B�t�X6��OF���O����O"�}b��J�"`�'Ǉ8��)�$B�g�����A7�����>��'�$7�0�i�	q# C�WƦ�DI1��@��g��K�4��$l�֜�M��OƄAwwG����aر:��\+'�@��D�a���,E%4�OL���O6��O��d�O����O��F�!A�
���Y����s��Ot��Ycfdc��A�f�D�O�]m��?�Gx�e��Ş���5�؈ �FT����?Y��i>X6m`�z`F�|J��#��v��A���~GdA3���4��q�DX�=���,&�D���Һ�Ӝ|"�'J2&A�Y�ȀJ��|��6O�Y^��'���'z���ПH�'��7͇	��Z�)v~���eлb|�PMьR����<�)O���O�����)��4�?�v�� VN��3t�=ZC&H���ڊ+Y���ߴ�y2�']�}ӱ%�=]���\������Ճplҭ_��T �[�$����ь���	ӟ���̟\������: h�#�D4��23t9cV�ͳ�?���?Ѣ�itH�Q�OAB�kӢb�زpA�#�}��ꉭ\n�0�dm���M����ȼ)�������� � �iX�='ư���;��I�dD	�����`,0���<���?����?�'̎f�����#ß
N����	�?�������8�fe���ʟԔO�!W�B)<N�aA��_��<x�O��'f�6m���'��Gt�cԁ  5�����:�ruA�<�R	3�X~�O����q��Ĉ%����a}��P�F�,�p�r�Q�`�IȟH��Οb>ɔ'��7�S�9��A5n��W���(G|PQdl����$�Ħ��q�	����u ��4v�ܚ7�\e�*���\��M{��VM��
�4�y��'6�8��"_�Oo���O����OP�|�:�݁���S�7O�ʓ�?)���?��?�����)	Kڬ��LK�1�Te�Q�F�m�Xm�B(��I���	R�s��y��������fR\)E���Ix�!
�׾	3�v�m�\�'�b>��@Ҧ�ϓIX�2'�bH�gd�$�ϓaRpq�F�1s@ؐCJ>y,O���O
�x���<��`��.ְ<�2��Oh���O�$�<��i=01*v�'p�'�H��e&��[�R)��R7���Q3���^}bBg�0�nژ�ē��pD�ɉJ�`I��J�oHRh�'��p)R+��4������ +����fn�'�*�	B�+���B�e��`�I�4�	韀F�4�'���Z�
��K�Z|� �5 ������'�,6mϦl���O�o�g�Ӽ��وx�q�d&̶�ܽP]����9�M��i)�7ME9Qyx6�$?Q�L\����b�҈d��$�%WQB�hcI�%h���I>Y+Of���Ov���O����O�9��!B�kC���� ׯh���
�<���iI4pp�'���'���y!��i�� "�O�fe����KT��k�w�İ%�b>�Ѱd����T���U�ExG��x���7��Uy"��~���8���P%�(�'��!�� m,�㦓{iRtP��'���'r�����^��޴�6���G��QCD^!*�#SE�7L�D�B���$Q}Bjj��)mڡ�M�ph�4]�t��@�C�n)cc���ti�T�޴���	|<U��� p�<��>�nJ�z�V�B����G��Q��냩p�D�Or���O��Ol��&�S�2�|��	;&,�+#�@�'��mdӰа�9�<�$�Ҧe'������x���ՉGB�8��n���ē��v�l��)ΛN�7-'?��G
z%��E�5#�U"Fɇ��X�"���8�P�1"?���<���?����?��gX$mz�)���%<C��ag�H�?����d���j��s��Iܟ��O�b�RqFH#K�
���ç�|m��O��'/`7��Ϧ�J<�O[R��Ǫ�QZ��H�x�fqK�'��rl �@�c����4��i� �g��L>�_�D��8bP�º4t8�����?����?����?�|z(OYnSyV���IP/4̨5PqO�/)�����gly2�e�n��,�ĀJ}Bjc�L����T�a����u
^4#��uz`EɦA:�4���ܴ�yb�'��=�$�E�o��q@D_�訦	�<0�\ �QD��y��|#��e���'�2�''��'���'���E�r$��?����II�oT�`޴ZD ��?�����<a���y��@ ۘ@��+��e�uq�mL�J6m�ЦтI<�|���MӘ'sjyjU*E�8H��r�[�z�K�'�R�)�˕a�)k��|�[���̟܊���A܈e���,�T�ruG����	ܟ��IyyR�xӀ�*�`�O����O踓d�_�],l �E�*�R�[�/�$�O>��'��6�JƦ�'�xxu��E�-��h*wVE˃�+?Y'���j�G���.�T�[wZ>�$��S����ʅ?SB
̚�lA��2�D�O����O��$"��+���+�f��Ѫ24�lAK$Ή��?)�iZIj��'�2�q�B�O�9�s�G�L�>9a1��Wݚ8�a>O��o��M���iH(5�f�iD��=U��m���`;�4���P�=�<���V�J�9�'he�I|yR�'R�'�r�'��Hq���1��Bc�@Q�kJ�,�	%�M�S��+�?I��?AM~B��|��o��37B���(dH1 SQ���ٴ.ߛ6�,�� �|��ؓ�!�?:H{�d�'`8e8��3"ʓ�P�Y����u�)�D�<��	� #`\�y�J�2��HeC�>�?��?���?�'��	��	�!����ŌǄ?�����	�~B:��
b�h��4��'��@��fm��nZ6���bs��*a`$��#p\���V��	�'9� ��IO�P�Ԍ:�����w���B�ϓ PA���b��mB� �'���'��'��'{�|��N�|@ T[fG������O����O��l��`f��ܟT�޴����@�'M�yd��iB�e���9��xҠcӀInZ�?A
� ����?a�� �i{�m)���JM�w�"lu��4�ΑjH>	-O���O����O�������
���]�$��AV��$�O �h�V�T6"�	�\�O�.��ŮB�{u�A�DD�S����O`��'o�6M禑�H<�OR�@�/
<=���dC0A$:Y�Gq�J�(Ä�%N4�i>m����Һ�t�|���7g���SfEDU�έ�ƃw���'H��'���^�`Jڴpn��s��*�	�<R]�H���?����f��Md}R�n�<X1��0kށ��֋yԲ�����Ԧi �4l�L�x޴��0o��
P"V
S�˓� ��g����k�)Y�5N:�Γ���O���O��$�O$�D�|r�&zV������",�y��̛�lo�FWu��'ur����'<�7=�\����޻s���&�;ߊ$JC̦͝�P�4u����O��ųi��� �쐧���w�$D��ˑ�kv��W6O��;��=��d%���<I���?�!c�E	����oD/PЮ������?����?����$�Ӧ����\��ǟx�B ;J� �X�� 5��&*�v�� ��	��M��i `O|��| �4H k�aR�� �y�'�d!"��I�Ta^�����Z�U������Ac��҂"��:��9
��1�2�'5��'��s�5Y1�	 q(ԛm#G����g�@П��۴b3�9s��?Aвi7�O��,^y0�h�f�N%���l����ƦMKشR���]T�����Z��-��ţ��8~Y�Љ�K;I��yʡ"?�t�&�h�'���'�R�'7r�'�x��Z�7��`�o	�y
U�Z��+�4,K��C��?�����y��6�~1pa�,jTl�7b\M��1�M��i�BO�I��P��ߊYG(TB�$26hmR�[/`ʨ���ͤnIb���a#փ��u�-�D�<�U�K&t2,�2�R��ॉ����?����?Y���?�'���R�ퟔ�֯��6f@5�E�s���� ��P)�4��'�Z��&�`��ioZ6E�٨��܃�T����;��Q˵�覍�'c��j�S�_0�2א���w�z]�P��898~	JҪՖ$@����'�r�'���'���'�����٭5�RA��bG�%8 i�� �O����O|om,(�'�,6�!���	b�����Ck�z�^�c�x�%��R�4*��O�*�5�in��%;b���K{֝JAK��v!�Bi�%T7�!��ai��eyR�'�"�'��h6.���RƐ�!eJ�T+�R��'O剠�M�%��?Y���?�-����Ӧ
�h��@T"T4Fw�0�����Omځ�M뢚x�O�D-͖8��&j@�|����
�s�ҬؐK�"G�ʑ(�_���S
��u��B��'��}8�! �)���V@�2���sV�'4��'b����OO�ɣ�M�ǮF?-��ig3D��M�Ҭӕ%������?	��i_�Oy�'�7��8�H���}V�x�e�_��	lZ�M����M��O�@{%ƅ�j.�`Ҵ%�<�⯜�)�:����9=�r-�6"��<�*O����O����O����O��'u'��j�D:2���:��B�7fr��i�aw�'D2�'���y�l��.�	r�:�(6C�,}449�mX<;?�lZ7�M� �x����W4^B��3O��9�ɚ�)d����
�-s(9ʡ2O��C��Yv�ߏ9��'#��X�	���a�M�7=�̱�N��T��֟�IڟL�'l�6�ƛ2g�ʓ�?�b���i	�Lc��'�Y?f[��,گO&}lZ�M{W�x�F$r�hzV-V(:��X(��Q	���^�hf�� c���6D���sݍ���0]���Mሧ�ғ3��p	��?����?���h�h��ӡ~͈�Z����L�La��	',��������I�Py�-p����"k��Iːッ������[�&扤�M0�i0t7MAM6m|�8��
]n"Uo#h����wl\
zs"S���@�2�$ O�	ay��'	��'���' O�*I�t��V�\���n�>���MK�*��?����?�H~��bI����?��Ÿ���$NZ%�T���ܴ?���)��A�L3 �H��!8�n}���	B�x���A 
>-p�$�r#��u�"<�D�<���o	��(W�c�����?���?���?ͧ�����aA�dGܟ�A��5S���Q���&f<1���ڟxݴ��'�L�bK��~��(n��	��؋�i�&PBA�Td^�yh"�ص��ܦY�'��.���n!������w̌��t�U���Ԩ3(D6�e��'F"�'��'���'���4�Ĭčb��9�g�*%P@0r�ON��O�%l<I$�ɟ�Bܴ��L�>�!�_�1?�,�S�
_n�؄�x�kd���mz>�3�V��9�'��]PC'��^(]+H51��P��$� +@����'��	����	ǟ��I�oF���	�RA�q�`�	���ɟ��'@�6m�7v�F��O����|"&�O["��0�e_@���^~2�>!�i 6��H�)�e�5n����AȖ�^����!_ >Y��	� W���/O�I�"	{P��!��\ܽP!��!IR��%a_8G������?���?)�Ş��Ʀ�J �L
��!C

}H`�)�����ޟ��ߴ��'$��8�����}@)Op��x�%�i�6͘�u�*ZЦ)�'���P`�L��HyPQ�D�'��1!g,Ёc�X�O��Ʉbr��'<2�'6"�'S��'g�~@�໵��a`	�@J�4�u�Gw��C3O �D�O����Ē���2�b�%ǁ$g�bBk�&2dJ9Q�4w��Ɛ|��d�M�:Od)�  ��r�:�3Ө� �&%�T3OR��V,:<�&P�J2�İ<�'�?!GoG2{�����9�|�bwg��?����?�����Q�Z�~������ؑ��4����ţ��sw�e����]�.��	�M;q�i��'�L�q0��,� �F0VW�%q�O��'��q��1˰�	^
~��݂�?Y�c�;`r!;�P"U��P"�΀�?q���?���?���I�O�Q��G�Y��(�!���854ȓ���O�oڇ2��Q���4�|Ms�͈�0X3�L�!�ȓ�8O�mZ��M��#��u��4�y��'0���	{��R[dAW�ӋzW0�@�� Z�Rʦ�|2V���8��˟��şx��"N514�#�!��BAb�F@yMt����;O���OƓ��$�&,؜ �,�+Pd�����u�'AZ7W���%�b>����"� �	���(@�m(��ҁr���1 ,!�	��4!+�A�ݺ�@�|�\�P��[�k	�))5�
W���B���ҟ���ԟ�	��SZy"�O��:�'��e��)m����r'W!,&�@A�'��7�5�I&���!�4�?y�aB�S��,RB�[�j�rÖ26iQ�4���UGO(Qh�!,��OM����Њ�.���	��(�yr�'��'s��'�R��\=g5�t��غ��G)��/���O\��ڦE�`�??g�i��'�t���NE@x0-Z��=C��c��|�i}�n0nz>qv������'�tqR!o@�gt�JE���}�cmZ3;n�����T��'i�i>�I����I���K���.>>�{C�W�(��	����'��6�ͧB��d�O��d�|�;lHX��E�9n��*��S]~��>)��iX�7m:��?��3ײ��I�u&�$ ,����=Ry��%�&\7���|VGH��uGm2�$J]�� ��̟<z�2��D��+����O����O���i�<1s�i���c��)2��$m:Q��!���L:���SŦ��?�6Q��*�4Q�t�����m5f`�2˅&O\w�iB�I�Yʛ����Hn�-�q��~J�\)l�6t�3IE�6���y֭�<�.O����Ob���O����O�˧(g���/�4N����B�Lx�1�iw���'��'X��y��o���Ԡ	u��(��ĔL|#��\_�nZ��MkI>�|��I��MӚ'Y2E��Ŋ1^��]�F���M6�'}��k��]�Q24�[��|�W��П4ڶ�^+ �0����M�O���m��������	Ny�`���0×����h"z��D5J���!�+��D�4��?�X� cߴJ��v�|2A߯m��Jr,X�%��Yy�D����\�jZ<�PAi�11� ����{�}��~�����8
���g��M@<9 ��?A��?9��h���dZ����ja�	:evT@�Фd������HWb�˟�����M��wG&��dO�,R����%٬tg��ӟ'�b7M���iA�4&�l���4��D���['(Hz��P���]6i��0pM�jP�wJ�� y:����5�đ +q��ت�&֡G������G�:��H��A� ��&H�"����A@�����uj��)R�7t,��L܆�t(�F�� �|����
����'�&����F�%���7 �"h�x��%(�	�r�ْ@	8fjxb�	�S���񩂗7=�P��"�(|�(aX�+�*�����S>Zy��lF�E�&�zd%���[&%��Q�N4�t適MBjp* ��f��4nC�Q�vH��&���H�� �,�cꆝ]j0�e�$ �M�f�N(�ݴ�?����?��'!��I�$����R~�t�a7���R��\�ܴ�?����N!)�"��G�r�l9{`A	k�T��h'v����.o�*6��Ov���O����E}�S�P���*,��Q'�7Hk�P�0�X��M#�<�?)M>Y����'�4�����4��Q=U��#lӚ�$�O��$�}T(��'��	���n�DD�4jI��H�����-���>q󤞦�䓽?���?iT�;K2 �D
'z���h��F��f�'�
�bģ�>A,O���#������̅^~hy�'I�+�V��k�dNr�	џ ����L�'�6��d�Q9id܉)'d�� o�A�E ��E�듣��O��O����O��@E�~` ��f@Y�?FVq�1�7���<����?������N�>��/o_d2g �.��$���o�h7M�O���O�O���OR1R��ONh/2}��U ���[RĜ�RgN^}��'w"�'r����J����22�qs���&V�ŪRKʄf�m؟�$��I؟��
����O�pJ�F�%� Mxw*ϐ-�H�'�i�'�剄!Y�R����D�O��)M��q뱈�,;����4�9Kh^�%���I�r2�R��'���'8`|j��E��$jm@;7˶lZLy�ՠ`��7��Oj���O��	F{}Zc�1P���7 ��Zsi�x�vI@ߴ�?���%��Y�������Y��#���<��q1#�&��9K�f��������	�	�����?���Ob�Uݎ����T�?�"�+�$y��il��X�d>��ϟ�â�R�Dvp�
���md*�pR���M��?��?o��5Q���'��O���c攴k�*Ii��Y ��t�D�~� �O��D�O��
2� H#��>q����Γ;p�oҟ��.�����<�����scF� �ƍ3o��mP�� �v}"�ـC��'���'��V�x��aC�G�4���Ȣ7�ɨ��4b�O˓�?q-O�d�O|�DG$("�̠k �~|A�`��r�0�B�d�Oz���Oʓ/����2��:���e��A�E�����E�ib��ߟ�$�(��ߟ̱f�Qm?i@�P�{A���D�O�ԤDi�R}"�'l��'��ɹ`0�h�J|"���u�jBU+QU�y֌�!*����'.�'U剹Q7>9�	y�Ʉ�)�����1?�� aiX(�?����?+O�lYag}�ɟ�;'�nus� �]?��&dU�	E~`%�$�'�����'��O<���C�p3�Px��%�\�fX�$U����M��U?��I�?���Od 	b�-O	b����$� ɷ�i@剷?��	��ħ���q:�F�6��)��'��g-0|���hӜ���g����	˟4���?ͺN<�'5����)�o-D 1��ܣ�x:��iHl}��'+bQ�T&?�Iџ�������cf�8t�Tչ�AI�M����?��Y,h�t�x�OQ��O�e�ՏLb?2�ّ��:(�娧�i�R\�LJ��6��9Or�D�O���W�? 9�������J����i�4(�RO��O�˓�?	�GSL��MP����U�X����Z�q�I>f{���^��󟬖'���5qH #�ӭvh&��(N�[����W���I��?A���?٧)�Zr�dTӌH�fϣQ��}YrΈo̓�?)+OR��Y�;�D��,;��V)H�3��g�F�	\�6-�O8�d+�I�h�ɍU�����t�F�z$�7K��7�^�9��$�xR�'C�ӟPE�x���'M��9�D� r<����r8"4�7Fqӂ㟈�	�,���{4Ox@F�nK8�;��ǰWٌ���i��^���ɔ@0 �O���'��\c����KH�VX#"+D3^s>�SO<1��?�$e�a����<�O�~����/�� X1JːN(
܁�O|����WJ<���O`�D�O���<��Ve�в���m��Y(�&��gRN�n�П����$�X�5�)�ӊ8v�H@�T?"4� �ur7��4��D�Ot���+O�S�DT�˔���8���Z�@�
ㄔQ}��O>��DC)�&y
E���*$\�t��M+��?Q�0q� h*O�SH��0�@�r ��w>|�b��54G@�Dxr	7��O����O>����J�?^$x�"�
: *�U+�U��XZ�\KI<�'�?�N>�R�q��}9cf �>�F�QR�C*��I�lV�L��Y��ןT�'Ur�K'I��h�'҂Oۮ�#GJܫ\��ET]����L�?���?qw�ı4�0��%ڜ(� I��B�hrh�$.�|~��'���'�� �L��OV: ����b>��`^DU�aP�O����O�O��	�V���U�0���P�i��Y����6j�	��_�H����	Myr/�<<��l��u�S�'w���#���kV��9����}��p�Ibyr��;�B�~���O�HrC'��n��4y`��u����`�'��y�(�)�O���N�#�c�",캭�5f��[�<2��xB[��`6�ʟ�%?�'�=R7�		$������ܕ9	>�'O�e�����'�"�'���]��]נ\�p�	�rE�\zp�̴7��O��D�SYPEW�����
1�9���{b��Zg�ҸUћ�@]5O56��O��D�O����B}�^������H��`.�"+d�(H0k��M�$�[�<IL>�����'$ �۰k؎J�ȈȔA.q�<��7��O���O�ă�q}"\����S?���ڪ%p�m�5'�!S�R��$IɦY�	uy�h��yʟ��$�O��ڪ+20��'�O�dl3GH���mZ��K��2����<������Ok�X;l[�p-��3���c$1G�I�N3��^y�'�b�'{�	1c�� �H�%{�(@��GΔ(�����<!�����O����Ov�x+�#?c��R���ҡ�m8���<���?�����N�y�&�̧Bl�"�E�P����#K��)��lZ\y��'Q�	ܟ��	Ο�A�oj��Qc%�	AJD���z�\J'��M3��?1��?�/ON��V��}����5�w�tj�tT�ܳ��at�Y�4�?Y,OJ���O�d��Ĥ|n�='�j(y�l_n,
Q{�b��*��7��O:���<)�'��6�Sɟ��I�?=�Qk�[=�A�'���8�F��B����$�On�d�Ol��4O&��<I�OV�-I��[*G��#�N�%~5"�4��.Fe�!l����	�������� �K�$Cs���I�z�a�i!��'\Ƞ)�'$2R���}"s�T+�xH)&���C�,���#��c��M����?����B#U�X�'�Zك1L�n�(L���	/��L:#,a���aD8O&���<����'���	�N�7ꌅJ52de�Ge��'�B�'��ȣcǬ>�/Oz���� ���J���i2h�%~�L#top�^�D�<���^�<�O�R�'���Ϻz��!�0�sQ$�CN�6�O�,#!A�F}RT���I~yB��5v�Q�"���x$(z�vAa��̓Z���\�	��	�����$�'-�x�/�8i��păV���+7犃_ꓧ�D�O(��?����?I4� (�]����sb�Z���?>։��?q��?����?�)O����R�|"��Ax�BZ뇓%���E����'^V��	ȟ|��"3
��Jh�֣�0" a7�Qr�|tlZ͟���ן���Oy����꧛?�1pQ>���d�x�x
Ya�ym�����'���'��D$��'0"��@��� D8;�T�
)�1�ڴ�?	����$�1�h�O���'�4*���d�@c���f��d�S$/m���?����?Y��P~2Y����I1��Q�<L��%޽�d,l�Vy ��&�7��O����O��i�}}Zw��!0&�*>��a+�䝟m��޴�?I���,q�$�l�}����;D�����! 
�r)�@����ch��M����?���B[��'���Z���'{�b��δ7��&-uӚ��?O����<�����'�(�����3��I�C�Aǘ�a�rӘ�$�O|�dW�8<�L�'������'��ؗFȽ6�TxQ�"ov��l����'Sx-қ��i�O��D�O��XFCN���c���fh*1жG����	�7��I�O˓�?�+O����	���T�	R�E���5_�(�d� �����IȟL�Iby҅ *���W��� \��
/�#"X���$�O�ʓ�?���?���0Cu��*��A�j�ڸ��� �b��p�'���'�r�'D�I�"
��8�π � $L�Q�:�Xr�X N��p�s�i��ʟ<�'�2�'+�!�y�H�@��Ĩ`���r� L��`ߪGWN듗?����?�*O�"So�@���'��\3�M0��Ã*�0�zt곎s���$�<��?��P�n����I�Ʋ���#{�d�р�)r�7-�O�D�<IF��Z�Sܟ0�I�?Y����~˶yZGÓ�U�Lqp �����O.���O��`V7O4��<��OK��*4"R5�Xb�A�=Ga�Ŋ�4��dVJr4n�����	ş<�S0�����R�/�!Z�n���(�<]x��h�iKR�'�x���'(@��<���$��/������<6ݨs*X�M+!^1U��V�'?��'Y�$�>�)Op|��dm&m���Y<<����S�"b��%������K����������!a;I�xIe�i6R�':⅚'Q
꓆���O���%
�@ t\���ME�6��<q��P��q�S�T�'��'$
�@UW%�ذQ���$F $��rn�����-1� p�',�I��L�'-Zc�1i�MY�q�tU��O�E\ȣ�OJ9��9O�ʓ�?����?�+O�@��̒�Aad���؁{<�3S�N�,�܄�'��Iş��'���'B�ϖc9z��v��!���	��z�'��'�2�'2Q�T��&�:��ī��
���;��Y�g�U���Mk.Op�İ<a��?���:`D�d��Y4�W�Z��@�Eb�(E��f�i���'�R�'��I*q�L9�����4p�f���EЖ/�� A"Y�$�~�n���D�'���'����y��'<�����!2d��<}���X����'|�Q�T2�DP7��	�O��$��J�)�bt��K���~h��0�_}B�'�R�'���'��s��'^�R�;$Ƀ�7���0��Ӡs#�HojyB��I 7M�O@���OP�)�`}Zw�*x�" 4�v�R�h��1��;ٴ�?	��&R|�Γ�?�.OD�>�A��G0�}Hѡ�|���b�,�! �W����������?qO<��=?Θ�7�S�N
�0����1�a[��i*�q��' �'���؄qJ�%�ELD���!��	ђ��l�쟌���ʠ�X=���?)���~R��#$Ă�zVFA�E�&UH�
>��'�@�y�'�r�'���q"'̒0 ��q�N�|�2�
�z�����w*�%���I۟x&��X�
M��83�*t|��E�1���iBP͓���O�D�O�ʓ��4� d��M��+���1~���.M�rC�'��'��'��' pH�@�L�:^\�EB,A-*��#H��y�U��������	Wy�X8iф�S5Fu���eZ�b�8l� ��HZ�OX�d�<����?i�������;�La8���'��qX+!^ښt3fT�,��럴��qy"7cd���`�H��4P�aG�%FqJ����@ͦm��ByB�'��'�m��'#�[�j��5��X��$r�~��ulZ�$��^yb`�.p]J�L�D�J���`�!\o������!�� %f�E�I�����m���Q�Vri��88@����@��f��¦��'�P�3�gd��,�ON2�O�@�H�^5���|��0#î��R�i�Z�M�DKԨ�?qO>�(����;-^JAẄ��옂K�2�$6��%�mZ���	����=�ē�?�R"ڨ.p��d.Z( s��G'̭6�Fj�!�r�|��i�O� C��Oe�u�a�n>���������	���ɠIص�}"�'|��{���ka8N\�Ճ�ʱO�L�r��O��D�O�%�G`��aKZi�G�f����#	�]�I�8��I<���?�.O�������So ?V/\1�C�3e�쳐\��(�Y`��ݟ�	�Ĕ'�<���온��o�EQ�,�0/�I6O��D�O�O��d�O�8)�C�=�a-�/�8y&��U6�Į<!��?�����[)a"���'@���E�jI.)�@��T��'�b�'�'�r�'���Ѷ�'RM��n���
�"�	���ZD�'�>1���?�������'U���$>���iԖ~���1�	�QCQ	�.�Mӈ�d�O@����O��D���#l���>�Cp�K�T�,���@o����O��s���Q����'z�\cY�-	'�~ ���b�T#Y�����}��'�0	�$�'�ɧ�	�-]�T �@ҷMV[� Q�@i��U�T�V"4�Mk�V?�I�?�X�O�وǯF�g+�����--
�ѻdV�8��9�~%�������O;�8)7ݨD±mI�1ӌ��4��`Ӷi���'s��O��O�)_�s"��hԺ)I��aǟ7��io�n)�1��ǟ�������U,�^؂c &��I�p��6}ЉoZ؟������ b�����|K�@p7���^�keF��xf�Ш�"d�&�O~��udBH�ԟh�Iן����0#*e��˻.�$��Y��M����=9��x�ODQ�$�CmA=J�ȉb��<���P��>�sIт�?9,O��$�O��İ<A)�'D�Pd����-�,�2!�����<C�xB�'lў��ɂT�b��	�%�X�cuD,s:M#ƦFş��'���'R�I����#�Q��P�q�.�T3.6<g��C"�M;���?������?����f��;/P�oZ�nP@4 a
S; #�0�֡W� r���?����?�+Otq aYV���	��OP?�下㮕�U�,�J۴�?iJ>1��?	�ŌW�q�&�𴬑_P:A��o G��xm���,�	gy�Eۻq{l��D��� ZpR7�8:��G	=	���0ƕx�'��O���B���6aA$E���'Ж:��6m�<�T�T�*���,�~����j��4�Ԥ�B��$_�qX�t���jӘ�$�O�0��I`�'R��}�P��.~��q[$�R����l�=C����4�?����?���a��'Z"�K<q�,p�m˔Ub�:�F�sx6M�)&���E�$���6�%hsGG�{S�$��Ǟ*s���3cQ!�_��`���R�/=m"c�ܚ"%�~ҁȉ}iD� P	�e*�i�y�*��G@�*E1 B_�$�>�:�-�c0����#W4܅�2k �m�z��E�?L�%��ݫY'Nx��bF4~<:�8Iʓ'���:�`��C �-����s�ڥE>�A`C>jj��i��7H�sO�4BU�L� KÙ"{T$��/�=�?���?��	_,�{��?9�O+���߶ �Tl�	͇c�$ ���(|��l�S�˼l��I�IB�T��c�@}�'��ڠm�4[�H��Q��=1�"$���2? ��ƨ�*��xb�*�. ����S�<�1�����ٟ�+�wB��Q�֎J? ˾�=����'�|!���9���i�׊h�!���]|��b�vl�qvMR�s��$�ߦ}��kyB.V6*���?�-�pё3�߆U�z|p嬍�$�j9IхW-n����O���#)�i��$P�E���y��˧���8��9 h�x�ÿ_�;f+P�	ݤ��S�:
1�4	N�OI�2ek�<�H|�@����[N~L2`����}���	&J/���OV�?q�$�<q��`�4�˱)q��e�ԇ�I�u�x5�7	�������8�|���P�I�<�p��;]�Bu1Q+Ì�`�'�����4�?	���iݞ{���D�O��d
i7���c� ���
�/��<���5d�1�LR6p�^W¬zMxY�!!�̘Ͽ{�
Z�7�2���$՞h�fL��ê7�~�1�O+ـMʤy)0xː�����}�ݿmZ�ز��7ƨ���P�r������ğH�	V~J~bK>�gK�z�h��͓"�$�@�@�<q�
�bǜ0*�*IP�m��l�C�'h"=ͧ�?A���2X4���ߝg5*����?���OJ��'"�?����?y��d����Ob�d�u�&��`="b��)��� D'E9a`����[:2p$��۟ ��@ă�'�F��Q�;U�<,���EN,��	ʵ�δ;e�Ωh(�0��C�:��$`�1Y���<��
^�k�z�s��"Tz�6'x?����ٟ��9F���R�5v�̝1!��KR��ȓ >�s���͐�>]1�}���i>�%����ہ�M����:��X�c�؉p= �ĥ�?����?y�l��h���?)�O7ڍ�E6X���5̕;.�Y���8U��M��ɀa��)��Ӹfh��F�R�'��E����V��h2�U�L�(��w��Ԝ���-A	���Z��O1Gb����+TP�'�J����?��j�'R�y��@�K�Hj7	D�<y�
N��-I�$۽��	���C�<�F`OI1P���Ɏ/fu��	B�<i�i��'!��i�v���O��'���dG^� `�ÔV�\���K�?Y���?�-�>���A��-����e�ya3�O4���`	�2�6����D��Dy�Lx����M�W�Y���`���!*Ru�W�50�l���M'\<�Dy��N�?Q@�� J��\�pE��@"�Pi�(R�!(�C��" �t�w�F0+f����
ݱ�����K�I��H�rMn>-�ǆMW+��ɩEL��ڴ�?q���J�0� ���O��tz�3��-C�n�BF��)[0}h�!���2D35LH�D`M���]&�����.���Ț�e��Dʑ#!e�0X_nB�eH=>5�	;gB� �����a�ZԸ�ǻU���>�܎uZ����&08ey����.��x���Oe&�"~�� R�`h0�+�D�l$8$)ܦNe.B䉭D8
����P�3Ћ� ��88��I��HO���Of$�@��oi��f���HWnTh���O��D�!|���E�O|���Ot�D�����Ӽ#7(O�&���QQ�xha�X�@� HkB�Pu�d/�$-Zm��(�P��0n �	9x���ɗG��C�l��F��&���ox�Tr��W�Ga�T(��?�� ܩq�1OD�pɒ>2T��2RX,��OJd���'+�7�����?A'P?�+��x�b��D��(@��ä"D��q�LT�Bl�$Cv.#y����ѫ���HO���'�1Oǣ�!.��:�H�l��i��۷�y�D9~��� ��	�3h�-�Q�&�y�* .\qf��rΔ�y�j�C �H��y�)YA���x���w���w���y�ʝD�N)Io�j����١�y��¦[��@�(��a�i��H��y��j����.��?Ơ`nM��yhF+8� `�Izҙx�$]��yRnZ<�Z�aS8�>��b%T��y
� Le�,ǯ4�q �(��L��"O5㒩�|SZ�*U� ��,�"O��(t�!$�� @� >{Nv��*OL��&��V؝�g ��%A:D�	�'��B�T$3��0g�ؔ�HH�'rB��"d�J\�
B��"[f�H��'X4%��էJG�Uv��?D�hՈ�'ﰌ���ǖe�Bq��M̌@L�i�	�'#�2�CA���ܡ���9O�e 	�'K���/J&�QA��̕`F��`�'�܂�G<Vsv����	.����'LĩiTᜭ#^�؛g'��#bd���'�� ���s��:W�Đ�MC�<1ՌS�#�m���!(��!�fTA�<I�̀d~��A-�k눉9d"SX�<���\it� ��	�nq���Q�<�Sď�=��� G�L�Iqh�g��H�<y�	��ʌ�C@	�q��F�<�M]�\��'�Ã�����~�<�C�Y<�d�Gۗbi`!�|�<��g��:��Pd�[�xAxX�t�Nb�<9b+5q8be��A�$�ȤC��_�<I�\=RQ~XRc�`�85cvB�F�<��O�1�2ظs�8[%0�c��}�<ѶbZ#��H�a��4M�!Sw�<�d���Ae���rU2�41+�t�<yA�!_L�8ꥢQs�ڕ�3�U�<�W	�Tp#C@�?����aIS�<�b�ѕ$?]g��1B�P�<�'��!�<𨞅o�H1�N�<��m�ZF�Q�d�G6��2�$�I�<)�Z�B���D�D����拝@�<1'�4�p �g�Q�d�ж	LA�<9��_^�:IP��	�A�x�@�w�<�fg���F�	!V�Ȩg��s�<#�52|M��g�'�f!�@�py�%����$�T��y"�Y�(|����j��}Rj�b��m���с�S�Q�la��gLa�!���(��M+ݰ�CW�dў܁�kF�h�TBw)�Ğ��� �p=�"Oxd�"!_��iS��C�ܕ�e�'����N�R�S�O�� �ۜd_ ��b��7H�� w"O�lj��a����'�	.�*ܳ�?�	U؞��q�8P���C�%G�V�"�KD<D���u�]�*Ӡ��7U���;D���a	���Y@秄�Wz&�	��9D�����s�y���6G�4�  �4D���s�F�w?����ɝ�����'D����Ǎ.K�Ԍ�6bQ:\���%D�����1|(�D�A�
�4Y�?D�ؒQ�ևO�@[�g��j~��u` D���`�U�mJD���j�D�S�0D� ��D)�XLj���6Y�.0D�y� E+0���zTeѣ�,�6d,D�P;4h*o����e/
Jb�+D��ЦO�:y�D�BZ�2J<	�"b+D���D�%��x)�> v< W�.D�4��(L�l��H���+� �b�d,D��!EDg��*	�/g�,��BQ��Py����(��
�,˂&V����,�y�/.��C@C��qETպ�BK;�y�JJD����$��lR2�JD����y"� /K;ri��+P�`��S�Aʃ�yB北S^ܹ��].A�z���"�y
� t5�r�w�m �
i3~�zB"Or]+ï�rH��J4�Z�+)
@�|2�J�k�(D^����W`ܓI���%
�"ʨA�Mʝʚ���I�_���g@�J�riA�H �%�d�1�R�����`�O���c,�)�ӄ6Š�[~~|��.��l�x�<ɒ�פM�6Ģ�
K$^�~}��&����I6}�R��F���E���D�PH�4aӓ'�/���[`���
����@V�'>\X��G�9�de���T����˕�m�z��'AF�XaK���?�g�/�<�0��$�|ئdS&z�,x�B�E3�qI��"	���Q�ɪ�ጂ3���� ���tÅāL�CU` 3�O��af>�P)1 �=i��ÀY�.�j��'L���p�G;/(��F�0{�u��*B�v��2�kĭ��6r��0��$h �sIJ7L/"����n��(�����I�?2���w��!5U*O�$z#�^�UZ!
z�((��nK�3z��Up�$�gF�4���[���95D��2a��OfUH�e�5���QGl\Sf�$���xa�����M�X�Ĥ�"�"Ql8��
<K�Υ��D]8h���O�yb�.\�"��a'>5�����5�Ő5'�`m���%FU�O9zyY�ާ5�"��(�F/�"�PH��Њ%�~Y�0aBˎi�F����d��B�J4��?_�(�F�/@,�Z��O�AV&��)  Y±dϿ
�m�t�J�	Ӳ :��J(D�h=����!H��۴%�WqO�l�ЋB�B �@���@���OL0���ֆ0"��i��f��
��>��,�^MI�*�+B���FE�>E2���OL1��$V>�z����뀔X��U�H�W*�z�X��p![�)FܨO�`0���&|4	`���v�y�@&�x�#FG�W���Ϝu}Bk3~1�f���a�#WM��@�5��Ct�	F��9p�l0�OGC�-Hʣjʰ6w�\��۱O<��Q[�����Ӽ|U�\����Ü<՞]��Ŷ<��(�E
�W:���a"8(��6i�^�Co�)S
0=�$(�45B)B��,'`��N�F��h·ŀ `���=�fH�HXt8Gh@�7*�1H�N^?�" F�>)*a+�)�.��$��`Pg�$C�i�\�K��р��JW'D'h-"��Fͤ>�&(V���H��ɃU�!3҄��4�b���]1�=ZA�	c��J� ��U��>�҂�b���nQ��q��gξm�HAs&G�K㖐P�/�ow���41j}X3�����')@1��.B�nU8��lk|�
��n����pѨ��(��*�Ș�+�%�v	�>q$@V�N�}3�$�U�,O�h��\�D�ؗ�
67v�ĀC�}�v��j7<Ov����S�=zv�@QbV�y!�p@S��K��2�N�
hGZr�n%p]�A��{2��nn�UZFŅ!7jTA9�ꀣ�~�JYr���HJߊ$�ѩ����'_�%�ա��t#�4c�(+	��u��>Y��J7D��6��l �V̺#<;��'���a-��ed�1L���xB�H�'jIA5��/�%@e�=���B�4�0i��$A �V8��CII?�I�7 ��6���	W8f-��� i�Ȍ9lq��r�k��p?y���B�!�=|��p�2#ϼ�M�Ī������O���7�ݏ�"��Ǎ��i������"6�'�<�B���AQ\����/,F��q�Q�[L���w����䆃 7�SG�'�Bq��͘c��ӱv�����1IzT���!3��¶��W6�XZ��V%g�������Nȁe+J`O��q;|�����7.��c���韈�ˇ^΀iz�_V�̘HdG1�[�� �`�Qg,�2ĮKs�(���I���s�l�2Ӥ�b�$�<�4��9��a�!g���r��謘�m��:�p
�0eꍨ�"ȩDw$My%FL��DI W�ΨZ���HpO¤7"Dd��L��<���&�!*÷'b��]�@�	C�/�"9A$�E�����ׂA����&�4m�(iP���5/����'h�H�Ԅ�$!���h�;	�d �=�FGд4cꅩ�a|?$���x�'B&�Z�#Ui{0��7(��3���A4"X�D�ΒZޜ��ЏZo��	�e5�8�s�'m� C�h�.4�X7.�"�� ��O�q�&-߈9���Y�2@��|j������Ǎ�?�Da#-ǭ1&$U"O
БR�ů-"���a�48���!e�/MmNܚ�Oݦm�%Å.2����'T"��A�S6RklCV[�R���ɡ>�8e)�P�>���P���N���T�L�#q��鵄>1�A��	07�#X
N�B�ja�Cs�"?��d�x	�Q��O9g՚���O��L�d�-)	u��E�ڈ�q
�'▜���?���sA���I5�a@�O|�� �;2\�L�'uCޢ~�@��4.Q`�wM^��x��Sk�I�<��c�*��qS���K �BvN42&� "�O���J'DA$>c�Ԋv���c��5+��ܠ͂��BO;�Ohh��5y�NB�����C�7[�����1���4�b��I7fz���� K�~�(C/A�`,L#?1կg��e��"�7-@�d$�iٹQ#�t�F�ߒ��4�RI��Q�!�dF�F��d$�ɓ�rp����*�I !�5���K�m<��5�'#�>-��jюf���l�oA���S�? p�c0��5_�^h[E$�w��x�b�|B,�57~y��B�P��9u�nA[��
�Lȇȓ3̰`����d��<Cr���9�	�ȓ[i^� d�M�'��x���2o#�x��5�A0���-n��˴�R�	:h��C����/��=ʈʀ�ުG��5�ȓ� mfdH.��Z����RԄ����RDZ�(�esU.�[xH��f��ң�!R���3����ȓ8p`y���Ɋ\�$)�HA;M��ȇ�~�|�;i�*�Mrb�*:Ȕ��r�����o֝n;��I���5;R݇ȓ̺虡 ˁ"��`�W�7>?v݇ȓ3��p2��$�.��D�^�����)$:8dn}��!��_���ȓ&)�]���y���U!�b��ȓ�����VP��p�0�5:��%�ȓ53nŒ@�E�<�8�p0�B-pP��ȓKrL�z���4�P�i�$(zE�h�ȓ-�^�����*q�AG�'1��ń�>�pS$I!f���"\�k.�ȓI�*(����wL�p)��� �ȓ>�T�� �;��qk��Wm��ȓ:�9��L�V9��SB�x��h��s����'铛%/���e�+s��ȓ3*,��V��_}�8�!��H�hA�ȓT���ↂ�zW���t A�Q:���t#�<iP�HQ�T!�s��h��ȓ|�la"sFٕt�\}*�@=	���ȓQ���`&Q1,��E��& ��R��SV�
�V���Q�I("�E��@�E�vGٍ?��0I�$Z�<l�-�ȓX]��k�e�1vF����&R�JI��o���S�S<fP@B<�2P��Ji��z7��2\�L�e,�/S�������i�P��_a���d�Q#�͆ȓa��U�ȿ8*vu��mdh�8�ȓ?�<!!��̪c��<+����Q�`�ȓv
�	@��;�2����ƶi��l�ȓ>%��!�`͚N�����&�9"jɆȓ�A���83�Ƽ�Q�V�*��U�ȓⰰDD	�Z�+���X��Ȇ�u���R�o^,=�H�ZP$@!MH���Nwr�u�$<�v@ץ�}e����.�D(7�__2H��E�E%$��ȓR����#�'���WB������/y��ZDb�G���*'t���=)���箅~�6��ԭ�U1���ȓUl`A���f)�p�S�L(���ȓ`pɃ���؁��¯�8D��;j����S�l�dh�6�-F^<I��6���B�H�lŦ5)R����&��ȓE��9s���9Ğ���O+-��E���Ҹ��Ȓ�� ��E�q��|�ȓA��(�%Ñ�[10	�3�_�*�!��09Ĭ�AlL�'k��;��աip�ȓ C�E�bd���8q��j��|�ȓm��E��	�W�D��ĳQ(Ąȓ%�0�A*�C���ѣ�ǩ��e��R��A0K�?-d�&�S
@�P��5���oQ�8:�iaNȼR�L�ȓێAz̔� ����Lضr�zq�ȓ^�!#�ĕeh
a���Ҿ,0نȓy�,	B��=Jq��S9l&��S�? >����%o��#g�'�h�h�"OD�fEPU���p0��O�j[�"O��y�j{L3j�;M����"O�U�C-FIe�##Q�y>Hh#�"O��F�8	*!�Ğ}O+�6�y�mA F����P�"�#ULM��y�Ɩ�
6�C�޵r��x%�Ӫ�y��ӆ:nyr0CG �8�
��Z2�y�l�:d��:�Ε�����i��y����	�^106F̠or��ׅ���yb��:f�J��摅	E(Aw���y�&�H*:��o�M`�]
���7�y���8%|�k��ܻ5�0!S��yR��C="�Lڣ#49��'&�yB�o_z���g���R0+w)��y����ްq�'X<{7Ԭ�q`	(�yB
�W]J�PDu	��@����<�ȓ:FkR�
��%׆s�V=�ȓ<=b	a��X�&b*p��̇��؅���"�W���P�Wl՞!֖)�ȓ=�|����$��8h��ݝ&(9��7NuB�f��7��̳�i�0#$�ȓ �ޝ�݃^؉c�l¬���ȓ����t������\�:�I�ȓb�&@i�A��&f|t��9���ȓC�B�'k��2t�ՙ� ѐ	!2D�ȓ]���-B�[Θ�0�FЂL�M����=�k��@���J�>U��Ew�Ͳ���1l�ȩ#!�X C�Ʌ!(�}�E�Є2��L��� wR�C��&���{��ȫM�� ;A㝣``B��!2�P����>cc�x`��?D�DB�I�E��b%��s��k��"s��B�ɣ&�b�h�ԘY�B-Y7�ӟC��C�I-"��l�S!��K<.I+�L�5t�C�3~��Rc��F"�ڤ,O��hC�I�^�<qcb�9fH��1vaA�P�zB��ik��8��Q6vB�QcE�1%�`B䉔A�7�y���k�
T�ES�C�	�]pգ��y�L�J5c�6e��'�a|" '�PQ��
�#�L6=�\��D��8`a =�ꭓ��4D���b��"D�ԋ���[x�$V�>�����O;�fy�#~JWm���1�r˚tkDHA�/�h�<���Q2OFbT�]��<�/�~�<�`��O���Ў����#�B�<q�$W�3P0���&QR}��`�c}�<ia̖9�^\�`�H8�̔X#��z�<Y��w�,l� ��`q��be�n�<�P�Ӊ&����� &�K��^n�<Q��^�"�y��^�p6XH�.Hg�<�Ѭ�"1��c�`�Bjb�
@^�<�W	�WH��x%
�*{�M�#��\�<�c�k	��k�k
^��A����Z�<	�ǐ=q΍��kÌ���z�^�<Q��ϰu�lh�����5Rs��t�<w��#]`�@@ŉ8w�p8��)VY�<����(���`�#��~���W�<��N��c�`4AC5{���ش'�G�<)����J⪤��a�:t:��B
�E�<1��ե-�α2��8(�U`�F�<���/B�5��\	xm����Z�<�̗�!�����h�R,��	�R�<ѳe\�"� �sa�(�"=�U#JQ�<� ���+]�u��mC��D��9���	L����L�p�PUh�Wu ��m"D�����6d�䍘�˯ Q� ��!D�Lk��� D��3�
%"�p*O~�#�.�%�h�!�)es8�"O���T@�=jn����JS7?iZ��"O&]
A,^��P�b� W���"O�d��E7m-��Y���kO����' ў"~����FX>e�W�6c�\	8��B��y��Q4��g�ҢJ_��rA)X=�y�o�8Ϟ��AWE�F���X��y2�̷Y�$8��Q�6<���K3�yb擘0������6��� N�y��If�����U\y.j����y� ���L���T4S��Ѧm���yR�Τ�@d�A^h�(-t�x:�'�� A�T=�U��b�>+V����'�<K�Q����%�����'��+�:���)3a "���'�0I�m�r�4L2r�n3����'�2a�B�Y>e�!�1*Ίh�<���'����N�l�� �1�A�]��%a�'�b䋰O�6]�Y�Ĥ��b�f%��'�]����z������ߢYM�|��'���J+7d%�a�K_P��u�
�'��x3��t��x�����i�
�'0 ��M67��#�^�Ҁ`h	�'.A�GeS5,��ʃ�řa��{�'���"kR�^�v�*��	�Q͸!�'����%M�P���B�G�L���'|��̋3/�╺��)qQ`���'�lu��F\�\9�]At�Ēq'�TH�'�ȴ�[�-������ه{n8xp�'\HH���Ĩ�sP�m��Ȍ�<���2��X�SL���ؑ7� YS"O�P�ӂ�#��9�h�� �h"O���`��s�(@����hM�D"OTJ0m�w���i��Ͷa��!�#"Oʥy*�3�����V<=�dHC"O@�8�+Ϊ\�Y����H�YQ�"OXɈFh��0�m�!i��`�H{g"OPy
�B"�ށz�է`t�Y��"O����.D�t���ڥUkPYB�"Ob�����O[6m0�CL�$4��p"O�\� �9ԁ���Z�((,� "O^x�H`;x�٣�ҥq	")��"O��cJMZ�vA����ٔ]Xw"ON�bʌY)���gɀr��=�"O�|j���$c@֤Aw Z=�B-aA"Od�3�إWr���BF��1�%y4"OPq(6c��>C�"�-rl��7"O��{v�,mz���a� #�D��`"Od��D�6~1��h��Y������"O��a7⏶72B`��׽w����"O��V>h��Ūew���1"O,���/�[�v��TK1h��`�"O�x�AoK9I~^#u'�(g&a��*OT�Y�ҕi)4=) AN�'/B�	�'o"�x3!ޫJ\�9�!M�!RZ� 	�'����Ȳ}���HC�b�~LQ�'�&�!�̟���%Z��ѹ�'�2}�"���<b�����y�#M�d��5��	ָ _�1��T�y����z�i��Y�{�e�f��y
� �hX���3,�̐�N	'LȾ��D"O<P�I\@q�ѐR��h�*@X1"O�A	�b�8cF}�#씋t���6"O�dP��� ����S�E��x�"O�<RR*�F�]Ys�3��A'"O�!��I[������9�2@q7"O4�[��%<~F1qS�>|�DJg"O���1Ɛ�UM$[�J޿<��)��"O�}hEb�34d���# MP�I0"O� y��F� ��|p�n�>d5���V"OH<�ЌQ?WP3�@�;Q��"O
�W%�0Ԉ$��!�� �}��"O�a���콩����r�Z�@�"Or8&�3x�8����L�v���"O�����>U���IeD_HMR�B�"O�`��kӭ|u
�d��L͑T"O�<E�G�h�8AӢώ5	Ių�"OX����S�w��,��NW8H���)�"O���r���K��!��b61�7"O� �g쀰x'�<�wH�dM��""O����m�P��s���*=&���"ODm"��ղ]��!�4ɕ+P�@ܱ"O�У�%�i�Ja������;@"O6�Ȁ�; �L!��
� B¡3p"O��� T�R�T$���F&�B"O�A��%�ܙ�a�:!��"O�yY�	B>р�`���N�ң"O���ׯp|% #͙�\p&"OR���'%:Af/�'N֤�0"O����ݐR�ڬ���&Q)��Z"OFj7jȽgIv9`amՌJ�h��"O���x��II�AƎ�n�"O�Q{�����\�DjVf��ň�"OJaۧ�)[S@U�f� 1r�"O�d� n�&^e4�����()>��"Od3D�*P,��g�{��c�"Or�QBƑ$؜��f�/2zF�0"O(�3׃�NR4���Le>��U"O��S��
& �&d�&�8%cz)�"O����"���XtF�-b���"O<�I� �Ѱw�[�!7̘�"O����A�Z��g��-E����"O:ؚ�f/wi��c��K� A����"O6@��Ah���OG991x�Y�"O��8v�&�Ni�0OהV�T�	�"Of�z%�0XoRM��L����"OB�ˡH�~&�x0a	�k��}��"O4Xm���1��W�:I�,X�"O:�;�H�3�gRУ'(p� B��9@�ʶf�.r��}�2O0R_�C�I:+�2ܪ�g��.G�A�,N�L"�C�	6%by36�3_b乳���bC�	�{��C� �:�"�̘=<�0C�	8(�D U�|��ؒl�
+����'�"л$K>�VxZ�(�Th��'C��(��9|{f���{�����'On�ˢ,��;�Eo�+t����'��T P�үv��ɒR�Βz4��3�'�J��5J�6;R����$u��:�'w�`J@��'L�g�Gd$&��	�'7ʅA(�!^�IA�N3Y���	�'�Z�{�l�$FE����O�Ba��
�'"�ʔ-Q�Bnz(��M��f�:��	�'�$q�G�XnZ�8`�X9X a	��� X�SfN�R؈�"I�#N�P K "Oh(�AI.>�Z��v	V�s���D"O���I���ȋ�n��dY�"O�u9�`��%��E�tH銄� "O P���	�Vf�X�����dha"O��{�/��D,X�:dB"y�J<��"O����7hi2����F=	�'��0�K�L��G��!S� \��'�`$ʑ�+\m�@"��J� H�'8a����V�"dPΗ�B��P��'*4X �̃|����B:�ұy�'���)���+?Vp�'e�G	�'46�j���!q-����[*t�hj	�'�f���ǎ�Q��� +eRI��'2z��� ��W�}��V�jh���'WF�0��;=;�d�����4[�q�	�'4��H���c@����}��y�'�0YQFf]�ٮGi�3}����'��ѩ��3�� ���oq1��'4���tn�	>%8}C `�1u6Pk�'W��"��,
1<;E'�=A� ��':j<��P�^����D#-N����'\����D��e	d��o�J�j�'��E�b�Z��U�c�d�����'*����傞�8��Q`I�`��'�B}�n�\��)�q�H�BL�	�'c��Qdܯ�(�j"n����'��A"��Ƕ!�%�P@E8]�4�X�'�Iz�%t(T*q��X�jt��'�0�j�-<2������~
�q��'�����e�^(����
�p��	
�'����풜l/���M�:h���'��i�)��腡6�M��.PP�'�QS�%M�$@<D��[�n���'/�ݺ�����UIT�϶yh�'�"I�@�<����0���J�H
�'��5 �kIx��	c����u�	�'!x���'�0)q�u*���'��}��%�9����kD��8�'Z)��aG)uX�d ŁM0r	c�'2 }pA�Hݮ�@���&n��Z	�']�J� �4��]�R�r��-D�`�πG �H$�H�#$"Y��h&D������;E~٨q�
e��b� &D�d9V#��Ra�M g��ŘSH"D�\CÂ�00C��{e��� �!D��$(Y,64���$A�=��>D�(8&#����9�7T!�U���:D���a. �L��Ir�mY����s�8D�\i�$R� �=v�r�Æ�(D�4ʤ/U�'����s	��6z4�UO'D����ś[�Ÿӆ�
 �A":D�*��	?|[`d�ƛ("�I��-*D�@���";y2�c'ə�:nM��l&D�T����4II����/��$�br�9D���!��)���	��S��hSR�5D�����.MW4=zt'!fn���2�6D�8yG�D�x�t|j���H)�4�J?D�����{la��ˈ��R�A-)D�d+4M�+�:ݹ1-��NFӥ4D�`��dD9F�d�cjn����e5D�,@f��$=^ ��A ΐ;���:%A3D�(���Ue����`�.!��jJ1D�T��؀QT)��яS�,!��-D�� |B�K�l�H��H�	?Ba��"O��2Ŧĉb����ԸN*�]��"O�T[��L�\߼�B���='2`��P"OV4�Iͺ(�μɔ"8A ��Z"O���+���q
s���C"O�(T�E+a�|�РŏKod�"OƝ����p����o[&ij�"O�p�.�7��Q��m�$���@�"OL�0�!M���#��T�L�s"O������Q ���߬n?�	�"O�R�&d[rAj���_*��
�"O\823�7K�\řQ˟k���F"O����2GQ=����J�N]�3"OH���Zrh�9E �5`�Z�R�"O.TI���i8uR�֐p��0�B"O��g���tY�Ed�UѸ|aw"O�Yx��]�C�Db�(d��\��"O�J�A\"&�>d �AR�<� C"O�Q�Q�F.� ���O4�n$�e"O�pG�̔s��T�.	�d�d��"O�m+`��j (Ie.�?~S�sr"O.�"�l��R<$��'EI̀e"OD�	Qm�>�&��4搓a8�`A"O:E�T����6�Q$3h! H�"O��I5j܈_�pIE���NV��"O�,`§�	x4{�O�0IH��t"O�)�G�&^"��	����{��!R"O�8T��h�����n�	�M�#"Od��"�P�!*2t�c�	9� x "O,���;-	ԑ{ W2q��U"O���Q�#HNA�b�F�bDt-"O���G��8sd}��
Ϋ0�p(�"O��2$�!KG&.d�8�c��2P_!򤛃a�"�����L�l	aG[�K@!�F�5�԰3�ÆMv�<���L�.!�S{8�)��H$L�2\j �ˇsw!�䍢���&E>i�X��F��:m!� L&�ɕ5)^�G�J�/`!�]�T�G��7[�<��	?8L!�$M�hܹ��Ǉ��J2"WsJ!�ā�-�u�Al�'J~��C��R.0B!���ye�ai�@�����UOF�P!򄎮2�]�S/�B`"@��n�h!��Q�3�xc%ۡ_T�)�C�CZ!�d��	�@9Ӵ"��/�<�Ё�M�!��Q�D�HtE�c��1�Td] I�!��RB�CV�ݏK��uV�S�!�DF&�	�`�4@�B�[�ѝU�!�$R>!�03�p{�3�B�=�!�$?���'��?Bl�AC�9~!��b�fU�NHi�j������{!�D�dA��%�(T�l}��hA�`!�d� ?�NT�NI�.��$SHؕK4!�	�l �BE�\� ��4!��$ɒ@谅F�b�0}��
j$!�D�<)"�q
��W6|��AP��:Y'!��V]q���5pd� k%F� �!�$�v��t�`�%sP3B�G�W�!�D�Ø��B�V�)�~��A�#8�!���丂QdC4(~��-Q�T!�d��d�h���Ϗ@�����ɶIl!�D��cj�1P�C�:�4�	�"żB\!��K�,���������KR�$�!��"�L����ʸ&܎ �s�I�+�!�� ���#gP�mq���R����"OF�P%�t���v-G�<���c�"Ofh�T+��^��,��ː�[��Ts�"O$0��)��9bԼKW+Q���,��"O���a�˶60��	� ��#"On-��G<�P�A�(ʝ��Yzq��e�O��y��+�>E-�ܠ�Κ�4YF��'� �{���J(D����X0܈j�'��\����:$ޠ�G\a�D��'3x���`J�>�)R�%bI��'C LZ�5o��-���E�aB���'��A�bT64}�d��L[�o��`�'���I�U#5s"L�j	��ъ���OX#~j��ݱ'�:�x��,jA"i�B"�h�<1 f�:L��M�WH��z0����y�<9&��w&��DfM�xHɲa�`�<�c�\�-�"Ԑb+6���)or�<�` -r�ݑӦ@�>kHUe.Ik�<�e�< 0��8���>g�d1�'JP�<�9/��<[E���$Y��L�'�?�z!�	�H��1AX�"^���7D��ңh��Q���$��.">B��"0D�pC�v����s���g�(���8D��1���s�
�0�&�D���3�9D�H�GElz�x�3K54���Ҡ$#D�H�6��g����ɱU��\s� D���qmЙs��q(&+����H D��Br@�
ϘH����>m�b0#��>D�4"ЏĂ[J�h�$ sJ�4h=D���g�2'�~[�b�>�x�G�>D��jQ��)*v-چ��*D�x"�%(D��HWdL�����'�1�Ƽ��$D���2
&i�	Ya��$f_�P�""D�X�g\�G��岰�_�:���X@�*D��X3��>@���+�
[AJ M)D����!J�T�����^�*0�@j1D�$�"�$�|-#QJ�-u����Fa/����NE+�KW�C�x��ɜX�v�"O���2̝�d^J�±�&v@�'"O�HiaDý͚,�''K��}�A"O8�*3E�%p��=��뀙�(�D"O����ό� �	�UbdaD�	y�T��HU@zyȑ V/gլ\��%D�8z\M�Lb���K�|��])��Or�D4§/�θQ S*���e��.p�I�ȓ7[�=Sq��<V�AI���d�U����R�"WA���y���R�����_�p�Lw Q�u����@���E�N��W���XC��RD�$2��`�'�a~B��-�Պ�ƠJ�4�ymA!*~i��˿f=P�����<��$̧%jV�ET�`�4�!��(`���#�ۯ2��6�P�
�!���{�F�!B�N�����ێE�!��H��`PV픴I�A8׎��}R��T�G�>��6�^�>��Uy���Y�<�����LR�D��R���T�<��S�:�yA^�{�Dua�of�<W���\�����t���$��e�<��&#��$���@!����a�<1��ۋ}���%"C�u������Q_�<��˕^˲͉3�}�4�`-�V�<y1��g1P��[��]��M�R�<��-;Qp�W��>�	�dHK�<� �Y�ʕ
R��%n\��ʵiF"O`]���{�����
�Z�<��"O�Y�L��xH@��޶h��Z�"Ops2
�@ɖTyQHX�F�4P$"O��ӳ����"�h��N�z!��"O��8!�:*n\��fT�q� �"O�tK$Ȗ�î�rժײR�0L� "O�M�Ҥ��8��1�j܎lZ�	��"O����F9t��Z���U���$"O��)sn�1�&���d�"O e���/o�z��K� �"O��l�W�BH�iP,M�2�Qd��f�O�ܽ���5��Ȥ�
�G V�P
���DG�CTb�sE�� `_� ��*�!�$�_�, �͐�\"r�FJܳX�!�dC�(�L(�b���aD	�p�B�w�!�G�@n�yEW"G��#*z!��H*{N���HLg�� �ׄ]�\!�$Ǆs̥Х��bsl�c�C�`Lў��_�O�@�Q��-��Q��mV/��a
�'�J�q
U#-���*�g�/CE2�
�'](4�4�1V!������3�e	�'(��'��^�\� C�"/����'�]B�K�"	0�B拕�R����
�'�����o��ț�D�zx,
�'F����j�(�<e�v�@�A�a����i�B�'�1���i¨�V�����A�ph�x�"O�(SU���7���2�'�?T8,�"O4�"��N	8cF5���z�N�"OHA;����S�栘��' ��A�	m��X͏�R�%"��L	����.3D���4�W*qb�e��ȉ�����l.D�8�V�b����v��I�T��R�<!���'���}��*������4
I<(�(UN��y2o�:9 3&�I�jb!�F��y�FD�f�g	�����H��x��EЊ���9h��#��_�Bў܄�~I��7�ҕD>詈���=f�LB��<)���a��ſE�~����+�TB��:�($��G	~�T��RDJ�w~H�=���?)���O��؀wh� -�v���${	�'����'��V���q�Ă5���'����7���l���,Az�(��d;�'1����ӴZopȳ �׌,�y�ȓb��ڗ �2!Z$�+Ɗ� !�q�ȓ.#ށQ��²��q�0�J+���un z�&!s*�} ��_�M��I��Q̓b&:��ˁ�e!�i(CL�)N[Xȇȓ/4`!��.����JΤy�x�ȓk"��acΘk����AќH����IP�	�<!���F��!��NI��)��\�F���O/~�SեIc�R �r � �q��'�)�#o�^^��� �KcHH(�'TD�1D��|)'����Ɍ"�)��^gF�)0���w��Y��$�y"՘�& �5�j��p6�
<�yRivp�	ƿ[֐���R��=�����Z)e�@��0�A0`�H�@4�V�N�!�d�	ڬ�"�_�E��! �愤T�!�W�	�5q�M�)@x�}@�%�#3�!��F{��*�o�gr��T�+?!���(v�U5�_ �hceA
x!��S�9���r�.̊VD� ��nF(.M!�$�F,HPЄL,�bp�sm�1+/!�� ��C���GA�a�B
�5�|S�"OZ,�dhי(�h���5L(
�"Op�p2�B�5�n(#��)^��u�p"OpՀ�&��.�Υ�a�T�R����/�S�I�d$E�j�1=D�x˕�ղ[R!�DB �"�C�(p*^�xqo )��}�X��W  B@dȥ郫,r%���1D�D�4@'uzɂ�(XYZib�"D���S��-��Ҥ9.�aE�+D�X��![I�S�풩m	�9���*D�$ ��H�m�t�rG�ۇ/�x���*D��1��H�$��
*��m�|d��K)D�P��+78=�Th��$��H��.�<����S>xZ=A��Q*}�T-���R5i�㟀��d�ࣗ\O���S?n���0�$D����.k�����O�;D`��)!D�̢�R��8\�4gB:(0�,A�!�$�;(�R����/I>ȁʇ#џ�G����G[�	A��ɔ��ϗ��yb�^�Ls
��,�}�b�H	��y"jZ�|���(�	�'l`BG*˘�?,Oj�O?������(��/�D����syb�'R�5A�Λ�b�h2�� ^�
�'e�<�`��OP>h�A`� �4		�'�
��ѩÜ%(\!��³,N��'Hr<y�ɷa  :���&,39�ϓ�O��CV)��Y\�-D}-p�"%"O����э:a���`m�-A6��Q�l�I�P�IC�Sg�T1O*$8�!�DL��)ˋ=��� "O�D
m�+%��ex��o_B�K7"Ojp��bҧx�8��"�M!biz�k�"OF�{�@��:]&}��HI6Ȗ�("O��k��nAjԺ���Q�-���'t��'��ɿZ�\��CaXT��C	V�C䉄4���!H��;�.�Z�hQ)sb�O˓��O���S1 y���&@�:���� �tC�	�B&
mhp.���2��C*�rC�IW�$pЂ�I�R��ZVh��K!�C�ɣ|&R,[TN�������!s��C�><<=��'�U�l�&h�|�\C��Z�]���<Jql!��jU�^�B�	1K H�!g���6$0��@:9���O�c�2BQ����c���F���?D�H+o �!qr]ڄ�Ωo��ʡ�?D��qš��3"��ӦQ�ub��KK#D��RB�rP�x��Nf�\	2G"D�x"���8)�� %%�2a���+;D�\��̠^���(R,rD�pF�#D�d�Æ�5Z��t#Gg��5�� �$<O0"<���v���&"/�$��(�D�<y��S�y�BYBc#�~�f���w�<�a&z(������3���p'z�<y���O���2�T`�I�D�ZP�<�GV*��x��ƀL��A7N\J�<Ah�f�L�#kA��H�<���*�ЭA�����e"�y�<Y5J2{!���Ѥ�:Rr�{�<�&�@9L�l�������\��/�v�<����]�� ���F6�调 Vw�<!'J"�DIz"
�����@�q�<����;��R3�_=;�$\0�e�<�r���AFz-D�9G��+�D�l�<I �V6^[V�zPg�3����	�i�<�uLYZwpD9F�]=j��c��b�<� 0�����h�0gO�^Ԛ8h�"O�$�g�}�ո����&�Nb�"O�u��73\�S�l߀wz��$"O����&ߩ�p u� 1g ���"O���DnK�J�ҕ�2GN��|0	�"O�ɰ�A�W��@��F6s�z�p�"O�1� f�a�����͚�yK�"ORm�%��)��!1 �\�7>R��"O�x!W.U^���AX�M9��ҀO�I�`��T~����aA�����0D�����JƢ1X��E�#֠�b-D����MK�1b���;^����0D��3f�ԛa�t��o0*�i%-0D��0R]��(�E�߁6l�Q��� D���@��k�	����0*��� D���EA�_�J�RtdZ�m(\5��=D�� ��0�Ua��mJ&��U�:D����!Su:5HS
!>��I 0�9D�H�t�L.z��������|��Ed,D� �b���
���E)D���dQO��u�S�sDx�8d�+D����׋�*X�V�~�n���<D��"�m��6f�h��8x�$��'D��q���a��Y�a�)�XZq�*D�8��G)�U�M/b'��*��%D�� �|�����ˉA�~�c�b%D���so���C�M�u�r��d�&D�h�ǫU��m���Ɣ�fi!��%D�l;�(� r��)�OG0��A0�&D�(;���o�T4RNٕz(�u��#D�L[� H�R#b��(X�M0�!D��91"��jl�헓`v� �O#D��S�fH�M�����Q*;]0�8R'D�ģW+}	�p���:��b!.:D��f	̀#��`���)���s�).D��A��8>� X���+#^*$�@�6D��[��دa�<���NI<EH8�2�3D�x1Э��a'� ���m�Jq61D�d�Gc<&@
�j��Q�_x4���-D�� ބRYj<HC��x*Ũb���<��N�7����@� �x(2TWz�<�U,^^`��.�p'�8r�x�<T�4�	�F� �~�)�TOQY�<�%�ĺa'�{�^)�+B�VS�<9�W�3m�MBԏD�a;���)SS�<���ԃ|'t#A(��>�
{�/�O�<QwDݛJ��	ʄ%�|��K��O�<A'��9QE�<!���h���yB�	{+`��Ɣ'v���V��y2�_���Y�s���)�y�jM��yr��* y���X3�������:�yB��7���q�,��=~�8vL��y�$��g�u���M�0k��녍L��yBCNjy6���fX�"XT(����y2���t$�� �P�`s!х�y�AX��y�
ܪi����ģ�yBl��V�H�8���������D�y�+�>J��31BĀ�V������ybFO!%GЍ-�������`D��y���&V��x�n���k3U��yr��XA���ڍE1`�3C�T<�y2!B7�Y��1+W8��a��y�
�.*����� �(���y2���.����#�egTd� k�9�y
� ,��"�w��z7NW�0���"O>,`�o��wDv�򢣁x���Ԕ|��'��O��6?Q�ŝ���	f��?_<8�G-Q�<�d��Z��ٰ��M
I� X�� g�<�����i2�f��.���	��Ww�<��*��
�ŋE���<��M1d�j�<9$78�\��_�*Z���(Mi�<�!��iW��������"�G^�<9�k���Q�cŇMLT�T�
ݟT��Ο��Igy�����@j�
?�<б���*����+D� ��(_|5C J�Qϐ� #�'D�����٘�h]�� 

#���$D�h��q����DT�*V��Rn D��So�9 ����!%�(����*D�dQၣ2�x2�W1�O$D�����F�g���s� ıq:HC��O��$>�$-�	�O���o��z��MQ�4aWD�W�yx�g>D�8c�G�ILj`sY��`��ȑ-�!�Dݹ�H���#g��J�D�?�!��(^}`�!�B-|�X`���V2r�!��^�(j�����]�J�æ��!�d�/;.%+�E۬N{dI8���!��F�L��Q�voX�.�q���2�}�0�	D�qv����JO�%Q�L�!�1D� �"� <Y�0XAP�P�6q�đp�9D���k^�sf���� ��u"�t�"D�0I�I�9�`���'(���@�>D��ۃ·8<1Q�燝"xF�r%(D����m �/V�Z�`ڣ^mܬ*�.14����R�h�����نb�����z�'�axB�Z&R�Z0ا L�;HJM ���y ޒ(���-���;qׄ�yb*� A���n
+��0���ybСE���2⋲x��-���=�y�A۰"��@�I��k�6(
3��y2g��[I@
�gӻ2D�I�ҏ���y2����,|ۦ�̩v������3�y£�+y����mb��hҹ�yb��)��Q��Q�E4�0�[1�y��Y�~� �a��^!E�9*��'�y��`���A)ޮn9"�څ�?�y�U�\%�ٔ%��8"WD�d�dB�I2^P���6tZ4:���0zTB�I4�2�⳦%!�,�{���4as B�	|6�к�%"�(Eg��b�VC䉇���h�OnR|�����dxVC�I7j�,�iU��7ItH�
2)L�y4C�bx�x�w�X�G���dAύbF�B䉊�D��2�Q�H�"("f���C�N��]I��=C��I���˫{ �C�	.`�}YO��F�����G��JC��44�$��r��]l��cwi�_nC䉻9�8)X�H�dxi��f<�B䉹}�Jtė�V��cW�X�b��B��Vz��cP�\�z3P��w��"�C�8�reh��֙^iH��u�T>{$�C䉣h^�\ʗc�8X�@�Y��Ӭ|j�C䉊)T���H *h R��r�Q��fB�I�&���b�VU(�	�fTtz�C�	�;���8��O�,u[�Lӟ|C�	�6�"�+�!�d��%A��O',VC��'�&��b�:0�~���_9.�NC�;HV��VB<�N�c���|FC�	8jV)%� )N��W+=e�(C�)� l��܈[OXl�6�W)�$�	��IO�O����G��LH!b��ir|��'��l�� Y(|����>Y�$eK�'ْ"mSd���ȏ0z��L��'���Ʉ��'v�֭ǒ,�s
�'��zсD�2�L�"���"~:��)
�'�RDK�(�;q㶵��*s_
�(�'e0!��S�L�ёP���i�L�k�'�lђ��;����2�Nh`�'�VQ�G� `uX��T/��P���'��Qj�KT+>�2��n�2v~�9��'Z4I٣�׶s����ӆZe]�R�'ez��KO0J��Y�T�>M���{�'i kV�_�:p�s,� T��\��'p����(���p��G�*<F��'BR�p�BP�T�����M��aݲ�z
�'���&��b��n"`z�h�'S�h`��3:&�+�����藶�y"D�Wr���i޾���!E�B�yD݄*� �$�\���;4�&�yR DD��m�I֝���[Ь �yrO�S��FFɵk�TyX �	9��Oj#~��V�:9��P���l�"�Kr�h�'�?�!�95"Xx1�O�8��E�s�5D��)D��.�0��1���Yv�5D��J�b�a�,j���J9Fؠբ%D��{'[�f����!
�t�1g>D�Ѓ�e!9
Q�!A�f�"@�;D���2U>G��x��0l�\]*7D��d��0a%��:�@\7fU�!�K)�	qyB�6w{���jP$h���W��y#�(D�x��Ì'���0e�g?�0��o2D���P�Jy2P�'k�P�px�p>D��dB�&;ܶ�C�E�s�)c�a;D��P�L�04�r�]D�@�W�=D���h,M>�����"��� �;D�HC0*�;.ˀEH�y�~��V�%ړ�?A��	ǹJF&�R�Λ-2���w"L'4�az"�&��'1�	�C	2�u� �;zi��'ʜy��]5�"�b����Be��'�b��v�ڕc��hА5 ��'�>43׉J>�ܔ��j�c��Tc	�'rD�J *�G4U��Ĕ�W�,i�'�v@��D$~Y��bJ���'��*�nvK(0�E��eQq�L񴄴<��O��	'�C�*�drIU(�>�F"O��T�@\��mh�&�6����"O�����F.T=J�̝��jU�"O���蓱i�^�s�YZ���2�"O��Z(�'�Tq�	I�t��ڦ"O��Y�S!'�:H6�WH/�D1"OS�&٦\��8Ce�;%b��'Z�'����/V�,�� �.D����X!��ǽi2칫�/>	)օye@ޏZ�!�$
5jZH�U���VB��!�$��hl[0b�;R�8�%O� �!�G�.�ڠ�B/K%�ΰҵ+n!�$�	aH`��Ú[������;X!�DB�P@�S'Ý����
:]Qaxr�#��D�O��(LT)�׀�*P�w��2l��B��7-;BJS� 2��#��;:X�B�	�4��@����#	�� �_:|n�B�	p{�9�E#O��z��`\x@C�Im9��&!�<WC��$n�3B�,C�)� ���I�"s�^�3D�P���m�"O"u��'e�DZ�j�$&\<�U�'��,�a�J?O���(�=]id��b-D�P�$f��hYRu2�,@�{U"+D�4��%�'Ax���S����3� $D��Bt%�,�(��v���	�  D��@e�L>i����%��5K�:�{#�(D�P{Gl��&���5�,>�D��(���Ov������1�#ţ"��hsC�
M�tX�"O��0E��d�I�`��	ie(&"O(8�Pޫu���y�@�
Z���""O.���.OjT���2�"OLIq�(�ry&�Y��%���ʵ"O�9�c'J
����/]	!J�� ��IH>�B�Ҡo��	e�+>w8�S���O6�Ԕ'n>m!cj�1��!h6G�]�%�w+"D�LR�DW�]x"�!"
YiD�tB�g?D������#2t4�ӆ 0����'9D���s�F:d_L�($�T��Ҍ�f�5D���6��/ϖl2��S�A���5D��m�i����-K 2$�Q��r�<9��&m�DH�tnۙF�Nt���p�<Y�$�4����6Gū��HJ���n�<iDC.�����,Z`-�g�<�����U-�]`!\M��XjS�Lf�<�a��g�<J�$��]��p#�+Hy�<1����n2�$;e��(`�0h[%h�v�<�s�Z*]�ٛe"*'�t%�]脇�f�:�+��;�8���-r̥�ȓ=��dZ���a�hU-p�����)Ru�A@��nȬ�S3��=&����a��Ļ�	��&���C�<��Є���`��މO�:|I@mU5=�X��g� �24�
�}�B�+g���(��x��F@l� \l�'
��axa��f۔�qb�քu�"<8���.
9�]��I]�H�⚀h �ʱNo���ȓv#��r2�QK�4`�C��7+���ȓAƆ-�4<:`�-0��Q�qYzI�ȓ9���Ӥ/	jA@�V�Y\���ȓ)R�h�6"*.-t!WF=[�~̆�/S�����|Kh��C ]�Bˀ��ȓy(B�sJz"@�)0��ȓG��ŊG�F6pG�HB��@!b���ȓKm�*&�
��EM�My(pI	�'\��SJ��la@��G�P��'�\L+�E��&9q!� _T �'�ԑ���Hj�N����òm��'T���kL8���M�>VK2�
�'
vHR�囐U� �'&Oc�@��'��H(���N �ƀqqp�'�����c��f ���Fl�m��M�
�'�b��S�NhH�Q'Jz+���
�'��}ru�[}4,,sq�(w<2�)�'BtՑDo�l*V�c���$h瀠��'����#��� qV [@���'lV|�K�4�>I���#�
���'�4q ����u�zx����2P����'od\���E�#w\��À��"��0��'�V@�� M��z�p���)R=r�'��(rU�0��%�(#����' :���_�g�]����	E��'kQ��3P�t@��'�P`�'n�d8ƆPqr��J6J�#D�� �0��T�� ֻ*'��C�"O*�@U�ރJE �	q�Q$��@�"Oh<xfP�"�J ��J\�"O4�����?6*M��iq �P3"O�9"w��}�Z��fP�q� 0J�"O~T��!�����xA��n�$͠`"O��ɑ!Vf"B�	R̓�.
�"O�}�oP�	;.W�</�,Mc4�k�<q0l�!���οp�|�I4m�e�<�G�>�8���<]�]��w�<���?Q���*@�D1G�f(1d'�o�<I.Ŵ^�HEiq�u~h��(i�<S�Ȅ&\�����PsĬX�.�f�<Q��V7T$�����<8m��b���f�<A2ąV�̽頊�Ӭ���a�<yp�T�a¹����~�,Pz��]�<q�M̆OF�L���!$Z��GFW�<9���U>$لcH�1��P�1�}�<�e��:�x3�9��D�x�<aCeN�4���\>�@`�Ot�<�o1hs���WFZ1{�$P҂o�<��
~�x�( �+F�"(�!�O�@V�ī��H:Q��m6n�zq!�d\�-�0st�ĦSgν0�"�h!�E�$�|(�A�*IƜ��?�!�R��q[��v����0 A1:P!�@+Y�2i�$]�aZI�W���k?!�$�y�xl�E�FG�����$!��ߋX��Ik�4�@հm
�g!��ɮe̪	�@\�Z��1��;eJ���e����@
��!BV��yB4#@�8֫��XF���	6�yr$��*�V�K��D"	��)9uH	"�yr�N1~�0x�t�\ y���L�>�yR��	+��q�(\�lo�ZF�Έ�?�����D�O����U�@�������'�B��O�&�!�$ˢ/Q^H12K��ʔy��q�!�%
Q�Xs��B6,����2,V!��4E� ��`��O,�-`sN��D!�$�BLT|Qg��y�ܜ��M���!�$ B1�%$ݸ�� m�
3�!�� 6q3PO[�1d�$Lڧ;�!�^+�F�A�͉�/-�y�⬕�$�!�DG�)\L!�A/-%\�H��ۗ�!�d"�V�:�`��8�2�(T��Y�!��Ё!,@!����U�B鑜�!��°l�J��r"C�e`a��`�!���fm�l��%@�hm萚�A�$@�!��N$-]N"��=E�,Cp��_�!�d�/c�	�s�D�x��ټ�!�D.y�yɰ$EJ�x$怓�-�!�$��M���6��`�(��Մ�!�d
< �J���Q�
�����],�!�$Y94B�P�j�@�.�q�W6�!�$�+8�<�q���!��-�1�7�!�:��ɠ�\�.����hZ60�!�Dƭ亘aƀ���TH�G�W�!���X�}3�H]h~�z��O�z���P&� ����+<�}Xl�#�yҏA���r�M����qb��yN�{(h}�v�wd<5 ���y��u1�Q��K%
� �V�6�y�)J������V�
$x�6I���yB� �
�{��\�Wp��aD��y
� x*L9/T�-)�� ' ��"O�⇧B�73h�i�2W�xp"O��K���P\R��&��6��l×"O �s'��/��y!��[e��Qc"OA;뉫'��]��#������"O���W�N!``ܕ ��L/{�B	I�"Oli�'/�#�+���[r��"OF�����@ O��&TjL "O���*P?�9�$R�V��9U"O�\�O�1X�j�z�KB<6���"Of ����7,�"�_���`D�O�<	���"�"�#TB�$In0��Gl�K�<���"�ܔ�uIIB��쐇&�F�<�0�?[�IOd��0'.�k�<Ҧ��j�(�!b�vEb���a�<�C�F��J%D�;\=G\�<���?rz|yR4�8�Fl���M�<�sl�	'=��jU��^�Q2��d�<�s��.Os��\�Ti`!�c�<	�A���A��P<�����$z�<����0���肆�/"k4�X0'y�<���с��d;A-դY.��	�`�s�<�6�B=
�@y���K���)w�x�<I3f��It�2�ٲJrj��B�Wn�<���%f,ĂǦ��rz������<�ec�q���p�־
n� tc�<�5�Z$��&���.��ώ`�<�F�^3pY����^<F\�S�GY�<A!B�?C��saX� ����&�T�<�4`�L@C��WF�XA*v�<�U�N�7�hs�ّ���&�LK�<I���zxh�$+�3�D��mG�<��iϫ5y�}i�j\�Wb>"f��g�<9��K$��ᰩ�j�4��X�<i'C�$C`��@��d����EJ�<�����Iwq¡���\lV����p�<�7��Vx}�e�U�r���ơFm�<��ȊI�T���U�{��+��g�<��,X���ǎT4I̬)��O^l�<��Fv^^aȉN��k'*^t�<��+��U�H���لfL�ʣ`�W�<YwN�20�\�)��V,Y`<�[T�<т"�_`p�7(*L]ش�XS�<a$�0WA�d�U�U�H�zqZ�*�K�<�r�J���Rg��p�
,�c�E�<�w{�c��lE�9(�H�p�����'���2�#D�n��{!�1l����	�'�NI�g
T�}0���dSD !s�'}Ƥ�DǗ������R�Z��'�J�BWC�pu��IS��!0�Y�'{V��`�10���q�=Q�@�z
�'k���D�����# �B��U
�'���J_�����f×<�n]�	�'���3��,;}4���NEzT"
�'=D����I�:���F7V���	�'���Wm׷n��E�-x�b�K	�'I��%�ȵi<�
�eׂB}�P�'�D�9�@
>	�=c�a�Q�M��'f�a�]�m�D�9S��v��%K�'"��eOU$��Ʌ�48�'�����.T�>YJ�)B�ѫ_��]��'�t|��,�~�Y�1��Y�"�)�'U)	�-�^ypdA`�C����'��#���:M�,59� -N%��s��� |�`&�)o��3b�W>=8p"O��%- �]�D��b��sN��p"Oza���Rj����DU�C"O�Q�W&l2Z��lލ2�� u"O(Mp�EcD� �H߷>��D�c"O`x�2�R�z�N�*��"�zȡc"O ���݈3���p^�J���u"O�PSFgZR(�3�ƥX/�h�@"OH�y�"�1��,k2�H�S"x���"Ob���h�86�D�qcM�A�|��e"O�C�@��EW((�1�фQ�����"O����S�!�%����x�X���"O��`Pؒ'^�t�HӤ�� �r"O�����76��ؠ�P<[e"OB�W�T����pdN�G�v%�G"O�8s��nn�4���y��e"O��k�]�VD����9�^�7"O4j� �3rp�	ZWgűS���"O48�����x���q'N�"O�}����t��B�a~�S�"O�0p��0Ȉ�:���Q/��"ON)BeΘ�1�.m�� S�4A�P�R"O��%o[�DȘg陠[^�E�6"O`�p�-Y���գ���nҀ��"O^T3�
��g��H�F˂qU�Db�"O�,Cf�$d�<e&J.z��<�E"OxD����
�Ha�e�le!"OxAB5�9Z��(��7T{n�XP"Or(R��3v^$��^�A�*�0�"O����'J�L0D�I�c��(�#"O�E�7Ǆ'>�,���N3eo�a�C"O !%FZ�0���c�9h.�h1"OXm��gS�1T���l{W�ic�"O�@�D�"C>J�qZ�:!�p�%"O\�;�o�s6�m�VgB:0$��"O�,��K�uS��(!��#$�9�"Ol���,~���B�C �$��"O��i)¹'zb\��%Q�U�T�Y�"O"��s( �G�0����^�Z!B"O�a�okj�t�h\�a�D,Bc"O$�S��!!C>u	����
z�Ԓ�"O��X��"}{0-�V�R����J�"O"��J@�-}T ��k��1�"OZ�i2ԥu��P���>��%�""O�(��^�J�\�T���R�_��y�#^�B`)�(�T/����V��yr�M?a��{D�=z�y�B���y��ƤVF9B������"�y�N��4-��U˙R�ʀbB�ѫ�ybP�z�U�C˄���L�y"H�Od���a�"@,��s1Ӕ�yb�7�X�9D [><z}�� ��yª$,G�q�HT�8��"��\�y"�	��xi8����g�q�F��y��\G'����`��g�݋�`�9�y�(y2�Mc!��-\���$�_��y�����L9E&H;_��Q�#�ɺ�y���N�k2g͔^���flE�yrA�"N�4}�͕/W�6u�E����yBi^ G�U����$>9T)@�-�y�Kǅe�FXH֌�1����ʅ�y�B��#�}�f�:+^,Q�����yb�F�w��YA(͗��H��O��y���A5���5zUP��ğ�y
� ��pluc�ip�֋('���"O��8�o�'2i���I�B)9"Od����<��%�V���M���H�"O�sàB;} �Z$@�f��LP'"O>U�0��c�ؘK󎄇~B�;G"O��R�!�+�؝��Tw��Jv"O��8���E�(��rF��U_��U"OpY��KӱfA`d�%E߸	:4ܪ�"O����$�PM�1b�O@�5"O~�+�̠d�Dpr��1�:1��"O�D)�J�;�q�e����\=[�"O�$��Ғ,��C��6�l�;�"O�$k&�W��PdP+�~'�4�4"O*Ш��N_���Z���67$)��"O�iA���4J�8�Z�J�^U�"O�����T��c I@,n�K�"O@��G�	���� �U0
�<�AC"O���"�BY�`[I�&�J'"ON�bbV,\M�9���k��̹B"Oĝ���ڞ�B1����Q�<��G"O �ѧdO�<W^`:�Z�Dr0�k�"O��S�j͸~1�Q���W��͋�"O���#z�b��%��G�$As"O�	�BN9�L<	T��C��ِ�"O��S�`�@jyR���!*�&1�C"Of����
4�܋�	ܤ5űs"Obh�B�Ӑ@�9�1)E�4,|%cA"O,h
�K�6o��H�a'R�&²y"O�] �h�P� �*D��&�ԋ�"OR��YI,f|�@o�!�
=��-�j�<�@J΋w���	׈6AR0�P�f�<q��7�<i��k��[Q���Wf�<����f{�h[���P0%�!`d�<93��9&|I�Ɓ
f�����\�<!��W.7�<��d�����v�Y[�<yt�Y=9��C�^�G��`�&�r�<�ЈN>7��EؑB��-RX)���r�<1v������Μ2~~��H�N�c�<���k��<��410j-���d�<I���G\�p�Ӆٶ7RV�Y��y�<� hڧT쨩Y"\�]�	�cCKM�<YD�·u���K؇T�LȲ���I�<VM�Y�p��?#[6@xQERF�<�&LO���c�Z�a�̍�U
�x�<�A,�<%�9��L_4UqHeCQK�Z�<	#l�
�
�h�@��I"T���V�<ipkگ���a%
��D���L�<�X�v�u"pi�-X�yI�HE�<���ʒ�۠�d	�_�P��6&*T�`��Ӕ?pT]�ĝ]*f���1D�hA�܍��!ǜ!uz</D�@�@+��P9xE����f�Z ��!�Od˓A=��6�V��	�sf	>���0O����=a�J�9�^��qiʧ{�"��c�cX���>�޴!>�xpk���*���E�m��=�ȓ:�6XV��%}�89p���Y�؍&��D{��t�޲u|p
B`@�&�8�`�J���yB������ځȉ<�xA���D)?�L<E�Di�;w����# |�*0�,*��d��Hu�����"�z@>nax2�'"�OR�P#KT,���i��A�N��"O*0�ڔyB����R��U���G{��;b򤫦�+!L4�r�G�C�!�D�)��ܻ3��s7T��i�(�!�� �#�f�$�*xz�BE5N�\�R[��G{��� �dj��! #ɖ�R�#].����,=��i�U �_8���e$	`C��^�b�:�	 �h�����GY 3�C䉎��Qbh���8�&Nا%NZC�I8��	�&��zid�-`��C��=1]�H��|Xl���f�[��C�	�-��  r��d���L�e��� ��~�e"PJW 1?1�c�VB�I�	��%�!��+B�Č��+T"d+C�I�q�4�k�)�M�<���ߜ$]�B��4^f� Z�#^�
�4	�ʁ$A�
B�	�ִ���N��@̣��	�����>���t���Q�J�]j|#�h�m�<��Aɽ��݀�ˁ�op�jA�WU�<1t
�"�4x٠�-C�~Ec5CO�<A�nVd܌(!m��]�a
��p?9�,�S�O~a�C#X"1��)�Ү̾Q$�'���[���7�\X��!��E�v��/O�6MJ}�d���J0r^���^jF
5��>D�t"@	P�)��r���*k��|J�/7D� ���,�J1""��g�L�`o3D�Pô/ٶ&��$S��� �p��F3D��V� =�$Q�C+D��1[T�>��PB�bc���L��d]6e�L��Ig��^�v���9�!�w��	ٱ"�#ZwQ����*4w��ATfW���0�	I�U��C��̡X�o� hrZѠ��E$��C�I��J����(���t��O���hO��æ,��8f�ǶA\�L�v�gKa��O ���#M�^�,U�6�t�\}�ȓTxB�#��W�����Ɂ@����ȓh�����.LI�Yu��>���p<�Pg��
F❠G�R�_R��k[|�<�Ǧ{tj
�
�
�j��D�~y�'F��ÊTQ��u�H�b86�k�y��O�"<��O&��#
�82�&���JA�1�f�q5\���'	�x"�'CҜ�b�ؽ}ze�T�?P�x��4��=I��B�Řj��8��p
ҼB��;�OVʓ1Ae�TJ�B��ޔ\l<�Fz��}���'��O���Gk
�0}���p	H%F��q��$3�'U�t�r̆�[l�hhWl�%�܉�ȓY�������W	Y�^����K�e��3�j��"�Y��Fzb���L�3+ft��/�a0x d�0D����iWh!�$�zX��O-D���+�*/&�)�fk�!��
��IPh<�SϿ>�R�H�D9G��xa��P����?��� �z�ȑ"�
�� �
�H�Iv���g��'�t��&%ME*pa6d5�O�	�<Q��I�x�JH�)�0~���KtVL�<����?��h5i�,w���a�H�'[ў�'.qf+p�LC��aʴ)�Ї�Q�����ʩ]� ���CP�6E��A�*�8���L��dc��3�$C�	:Z�4p��7�|d�a�Ԓ_�˓�hOQ>��%ݴ	R�IVa�/���� �-�d)�O�x��D�"�Х�@$�Fcb���'�Ĝ"W��Ų�]ԕ!х[�;Z!�ć�u����L�&Pᩲ�Q�:9!�$L�wR���ˁ�%rJ�S��V#)6!��%Z��+d��W�\�Xd���}����Q�e��aeb�PנЯ�t�V�b��⟠���Y��s� ��L������1Q�3�a3ړ�~r�xZ>� R%��,]�Ax���6̅����Ɂ"Oh���{����w�ʩ!P�'v!��ۓB�
`�%LG�2�b�b��t�|xچ�Dp*|J��=x����nW�yR \�!���)!��~��H@�"ܲ�(O|�=�OZ�8y����ae���W�Ƿ,��XA�'����	Q�\t��o\:&9�k�, �S��y�K
9��8���I{����R'�y�	�#0��TJRFS"�R��╘�hOz��i��V2����_�"����l��a!�ƔtH6E�Mmu�����]9;��6�l�	��?7��_��)� Ó
6HD��Ԇե}�!�ܸ�(H���g4��Ie��#bt��X��4� `�?��ʡ$��x¼!�9D���u�I�<Zд���H"�zDh1�6D�8���1|n����P\�N��D4��M+�4���l���'4j�h*V��8?x�90$"Of��6`�L[�F�O�\�	W"O��:���%Sf��e�уBWb y�"O���6Q�x�P5fO<�g"O��ЕfG6`{�%�agB\>�iS"Oԩ�$��oG�hr�f�<9� ��"OĬX«�`�#�T ��Z���eX�H��l�Z�̸��?����@�1��l7��A��D"6A�H�b�M&��D<�S�O�z����"x	�������-R1"O����o��}L�q���!jV�S"O���s�=X���"ˍe��a�F�'��;O68��#�_�r�1���3����"O��"�A̯ �h5�����Q����o�V}��hO�N��Z_b-��LR$����1��
�����i���bA�%[�����Q'e�����hӞ���OFO�g�$�1�L��c�ߴ+�����_�T�џ,�ɿ��Oy
шD	A]���G醌5��8��y2�ƙ5��y�Gǜ�>թ��NKnD!
͈��<i�O��'���AYb�ISd�P!3s���'ܰ;��N�4���r3L�0�b���}b�'�fd�įV`���ȍ9z� �	�'�\"5.!" 㶮�+B-�	�'��9��"(|Y~� u��� �d�	�'���q���*�a��lMD�ġ�'��e����. αKp� >�
�k�'&>����`��	�Ä� �jA��'QXm�O��, ����3}6�x��'L�i��˒ybd��Wm��s�ȴ�'"fLci�/MY���)�_0�H�'�F�6)�P�P�2m
�TY����'��-���ߠp��/8#�b��'���3��y$JL��C�/n���
�'���3P� �I�t�9w��!��Y*�'��,�v��y�<���["I�H��'�N�h�똾L���5샛 �XE@�';��)��>7�ؔ��Eid0��'�N�����X
.�(d]6b�� b�'aj��%n�	��QW"S�$����'�q��Ώ  Ad���Y�q��%��'����c ��o#|�JŲz��p�����ު��a�P�B�p�2dcW�b�<15�C�}(�	�B�%îX�4�b�<y 뒷d��v�M�j��
X�<A�逌1����eD+w*E1�T�<)$+	��,Uy�"�(W��`�aM�<�퍉ĐJ��=�T����L�<�C%������sH�k�.:�I�<� n�Bb 9��i��B�{t@I��"OV�)Ъ�/2;��GƝ_�z$;�"O�<�sJ(�4ի�/c����"O��B�(_�6��I������"Ol�Rf�
�p������O����"OV����I�^I���,TY0`"ORɑ��t��mڤ��Li�3"OZHv�Z��p�[���G�!�"O��ч�>f�T���d�$;��
�"O��Yd$^#SpVHBB�j
Xa�"O�Y���e%ab��Q�L[E"Odl��VQ�r��𠊓�(��"O�,�f�>]���"FŶF��3"O�}��Q:t��u`�ڨV��@S�"O�<bvKO�"P���WH]zb��"OD�r.9K�ɒ��q`��6"Oh�+6f�T���"��:U����"O��bոU�B��@wd��@�"O�A��D�7�hBfˉ6�HXK1�'+��`P�;Ci��PA��|,Z1%ƨRn�A`�'g�U90d��IV� %�FT����')~�ƃ�Lw&���}&v�
�'�D`��<�|�"�
�%�����'�P�T�M,d�=y0)[�'O=H ���)�2l�z��	�'����5H�$Z姈h�J���'�`"�\a�� 1��W;d���'�f$�F�P�(�����@Z��'$Re��@K��Py��;�>	��'�2-8bjI�gf���ª��(-�'L.�`�"� :�"5g��3}r�AJ�'���b�Z�#���B}� �z�'�>X
ʢ@>~�A�S�@�|��'R������`޼Ass�՟F���'�t�"�郦1��d)��g��'(�Y�w	�vv��3a�'Lɾ(q�'I��r�ƪ*aX�"O֋F�f ��'d�)ӊ��i��.ةHfڬ��'�� 8�N�;�Y@Q�Q�=��k�'�,�cE[%NV�` 	M�d�J̑�'>�;1��za�X�@�KHmD��'�X�v�M�O@U�X��5"p͘Y�<�T�"/��	gMÆS`~�y�.HI�<q&.�#�0�'�W�)��p/�}�<٥N" ��i�#􀀥z�<Y�b �^�Dԣ�*ݓ�:	E��y�<quǐ3z^��"j!=�^�7�B�<����4a��(r`ƕY0P	�T�Wq�<I'�2\���g��e3TeT�<�l��_@�������F�DkV�@z�<�Vgx-츶��&y�\v��m�<�5�S�)�4`i�*��c���9�Cw�<)'��=��J��3��S��f�<y�r����B��D�Gb�<����"q�G�B>D#�`R��k�<��
E5}?R�9��P�qq�!Bq-�l�<�p�7;�����[7�`#�O�S�<1$�<<��6�K�8��%#Wl�L�<�g��/?X���b� ]˂��v�<�rcef.�˱�^.�|��^D�<�qb����`���{H��
[a
B� C����])9��Z"FҧY��B�I=P�x�![r���i�@]]�B�	�*:��C� ,:�\�٢,�nB�)� ԼʦeZ#.k*��`ٟ]S���"OVy�	� :̢�k֠�<^Rޱ��"O��څF�z��=�S��0)e"OF��� �E�:E:�/ܭ4 5S�"O�uÀ!	�3��$K��J�0� `a"O0Ф��S^|T�FĎ�+,^�Y�"O�]���f��ՁD�$0 d"O������gB$	Y'o�w��ᰇ�'���*��>9�(ʢ/�8dK1MD�R�E���i�<I�T1<��T�+u�S@�Dn� ��5�b7����Ħ~��HXg�h��"OH2��(&�81 ��P��N�0CqO�A1��Y�țd�<W��k��=No�}�b�$D��"�Y�W��������mP.`���  �;�OH�8p�U~�r�0�U,>��R��',$9�kO|~r��v�����I%����&B��y�[/PiN���@���gM ͸'sX��Æf>�r��Ŀyp��g�B^�I�@l3D�H����+0bL�b6?r��j&��{��O�F�,O�̓`���LE��
�&$68u@�'C���a�?[WV
�L%\��1
�'#L@�@ܚ�a"	�� ���']�aqS��;w9����� �\h��'��)c.Z<E���u�B n��h�
�'�޼���K@��K^�W���b
�'���A�ĉ�@�q� @*2��	�'�l�2��&6��w��(M�z�
�'��QI`�x�]@�\<}�hb*O�ZT�	rW���K��|p�2S��s#�˘rJ p��b�F�<	bJ[9��2�gX�\�֨j�GU�"���a[z�r�*ٞW`���' c�֏ �ع��H�|ÌQ���c��lP�l�.\;V������_n�+Bd�m���ŃY�zQꥡ:��'�>��jީ`
v�@CJG0Ԅ���*�.��Z V1�`$�8�� N�h ��`e�
���p��K�
")yu��s8��y��<�N�Ô�њj�"�2ࣟ���b��d��	� �@�$>e���vI��O�5\Sb���%	>QZvk֋x�a~"B?%�u��A&� r#
�{h.�#�'
�,)g��T�B�3S�Ȯ}1� �p�I����r�W��P�H���&x�d͞l��P�Wk�
5l�]X6�W(����+�]AJtAbK��b�b��P�_�-����eD�'��i8��q�66m��c
�\��R�"
<+�ݔ$�Q��@H��8z��A� ���<Bձ��]� ���(��A�����T;��EY��;�J�#�˹?�Ezbɚ4+|����mF%�T4��	�~�%��m44�B�=;:H|�}B�䞞*$p��MKjR9��j�3V�����ҳ��� �� *��-s�n��:��7{ȺE@	�#A���ƫ�<�6�@�B��!f皬��i@͟0k�tz�Ȉ�`q��j�}�TD^�tnp�:A�HM���	h��Y�b��sny�#H���H� -v[ס>���0
�y��I�"�r�'�MK������
 �X*AS�<QsJr�t���*	fbPhUϐ0]�\ 7͗�[��h F�E'T�)���HO�%����4
F�B�#U(c�eɑ�'��}��Ňu�.p0w��s������$t��"+Cv�T�j��ـ:a}���Hy*D��S�Eq�cA��HO��h����4�D$+_��0�)�6)�b�GqmѪ��!="�LHG"O�Tif�s��2s(W�p������'���!g!�*2�~�3�k_�-l�?R��D�%J�A0���S�Z cY��C䉸7�4��B�<t���{@�-Tƙk�| ��/Q�c?O����\` A�􀎵
�����O ��v%�%-	�m�wN��0��JY�lU�T�
��*�>����%�0e#��U�OEj���.�Px�1AƏ;ev��N�u:R��ȓa; 
��6g�P��E�JB�����1s�J=�O�E�5`��������+ �1	��'y�H)1.In��H��ţ@�*�� �E���yR�$EAV-���ˮ v<�����'�fU!FK@(K���F���,eT���`��&l:�j��y
� �L�R��Ec6���O#	;E !NK�.�J�T�C��a!G"%�c>c�8:���2#�QK!t&���D)�O� aD(�#c鎠KWN���2K�MN��(���:v� ���߈/�a{�@��?)l(��Έ�[�JHв-����O����bƳ�8��K+�Z0C� mݩ��E�����e�5r�0��#D�����O1E�Q��+Ί4���a�!s�C��P�Z��xSJ��u*��30��'�QD��O�h�D��e�t�6�O�@����'R�Y;"k��P4R5��PD$Q�cE��&�BxJ� E"V�LiP��?V�]��+�d*&�&�ͻ\'��q��έ{DjȻ0H��̇�II��Ћ傈��t�K����8�9�^�H@���݂R���z�ԖD���+��5%K+%�""<a�e�9{�J0��h]�B��ȪS��{�'�ti��1�<m<"�����韺b�oL�VtI�	�jdB1��!��\� aĖ�a|����!��E�$mۢ|j3����?	"�%��u�fMK�2�(���#��I_�nѺL
�lӲ�yǩ�]~T!��U�
�8E����4�y��F�h�e솛�<a����()Լ��J�[�d�y0_���A���U<O$U�u/ *�y�C�(3���L�3wN� �thY5��>�Dș47����Jߑ@�B!�Ы�����G��&��)�U��U �1O��PR*^�D�V���$�>$�����O�`��r���'@ ў����I�?�~��&Y(����W�P��Ҕ�\�+o�����T�
5
�.�	M���RF��()�ه�I&A!Pm�R�ۯ{��H�����	�&�$U�(в��g�hȠ0܆t&):�*{>����M�Nb�i`@��XH�p㩘�X���Q@�"D���,� WT[�7E�<hx����<@� 04EFmT��1J�	�ܟ��i�I8�D~ޝ�%�J�f�ICV!�g,�bf&<�OF9+SN�BQ����F�j �]���E��ThK�:9h��V`�4@��	�,���Q�I� �<�J��<�- ��Ăs��>0�C+e0��QZAkL$(ߟ���'�fAJL �g�<?Ma��"OE�Սn�"|�1PHVd��W�p7�S0���P��>E���C��AB���*,M�l�yBK'F�Ar�L�"`
C�,���'aS��M8���fϝ1J2p�p�H�C����&�&D�eAF2��i�@�@>%�`ra�Of0ì6��>q��FƵA��Z�0�zY�%�m؞X�W��)���5V�	��6c�Da����:C�$-��3��!�ŝYB4�ɦ+D�*��=�5�Dx���-)�C���!�X�69s��Fق-��nb��=V:� B�\��9��FY.O�٧O<�C��Y�8�ៃ0��IX�▜!9��w!$D��yRON��$�"O�,n
��Lќ&��l9`˓�*� ���Q;8�r ����)�>�맯P�'q�zb���J���{�E��<Y�@�g��e;��V9_�l\�M�\�<ad�_5l8�;�I�-��(kAT^ܓgg��઎� ��#~!��+�0a�����B�>S'$�Z�<�2�ڐ`hN|ڳE
`}L9��/I�%I�fDg�D�(��	3z� )+%/Ǿ?��@Z��vzC䉇u���ã�:v(�@RiR;6xPgO[�?;�K�B)�Ov��Y�9��2�<�����'�pp*�'зZ�d��f�����&+�AD(!�ē�>��@�.92�8�G�/`��O���%,��ȟV�1E)K�]�)��P��Q�"O�PZeA�>$z+n�A^*���"O���%�X��)��Ҩ2D��Sg"O8!?_�hT���>(O��R"OR����:$K��GJ�5P�"O�z�/�� /p+���V	�8#U"O����}��豠l �<��"Ozm���/ ��R��í�d��"O�a�&��sT p�[��$��c"O@T1f�:K���q��|j��!"O���sk;��r`sH5f"OHE�q�),~�;¬t6���"ODyS@	ֿu-��#��"Z�`S"O^l���*!��ճ�g�bY	�"O���^�)���Y5�"����"O�%"�Q�J \U"��n��)�c"O� �9[��L�$!z��+�0��p�"O�|Q�ćlcƩKD(�VtV��"O:����A�BK�o^@!``"OL�;7(�(v���&K 1lv���"O2��e#5�ꖕ1����"O�A��揟\ٶը�HG�5���A"Oz@cˀ�F��%kw9�=��"O�ua���"QZH=�#��8g<�̀�"O�p�D�*h�J'�;w ��"O.��G�Z���J�CĻLN��"Oz�����cn��b҄�ܼ�"O��#؞"nr��'�:Z���T"Oґ〧�!s���,ı�qi�"Oz!�F���}_�@Yg�B8 j��"O���H�A�\ s��Y�7�N(�#"O���%&?l��]`Ga�;��AQ"Ovh*Vn�������.̘�{D"ORq���v�1���
I����r"O�l�_K�DC�n��5�Ry(v"O�\��DH.T�҅M̈́&�d��w"O�I�f/
W�@�àl^��1�0"OfT��Ŗq|�����`�p�`t"Ol�S��
�Pz`"�R�d��9X�"O��s�D�&������y���K@"O��+Ы�$l�V,��o\%��X�"O�[�.ߛ&P�ɳ�͜0ߜ���"O^�R��	�1��Ǎ�O��1 �"O�SW(�<�RsE^C�P� "O^p�%�;N	ɷ�R8je*��"O�$#�kԟ/�\���L�_|65s"Of͓2.�Z#��I��R4q1�"OI�``V�Ϙ� 7�$�u�"On(�dZ�0�j���.7T�q��"O(�i&FI�O��r�ƛX6�8w"O��AK�n���4��|:�"O�I7aGY�M���,V�H ["OT(�Q�Nw�M!A�ay��"O�Q�0�
�,��L��2��c"ODX�.|��u�PMP�C.e��"O��y ���N"��[�'U��<��G"O��8���&M��;Fe��|��Y�"O�y��ɏ�4g��DV-\y�"Op��CG��J��){W�8?���"O ���S���aC�j��؃"O��I�*���ӄxǬ��"O�IdA٬*����F��K�@�j�"O���C��/_P��%N�'|����"Ox,Ǩ !���$FXm�i;�"OP�z���;j�D,õ�P�_�h�s"O����Eа&#�	�s��K0�"O�A�a�y����7̌�k&�|C�"O\�A%Ž.�����[1?`I��"O�`�R*S*TkLy`�
кn��|�#"O�ƛ�R{����8�u��"OH��Eй�qh��؀YS"Oب�d`�b=Aƨ�!o���"O�"���0|�,hC$���l�3"O*�)���#`M�4���#��U��"O��U_j@Li�oۙ`�Qr"O� [�J�l�@۱��	8N��HA"O�� R��w�ԍ�d[}O��T"O�}3"�WeH��T���n'�U"%"OPX����0+,��i��JN���{r"O����`��T6�(T�3v�x���"O� ��`�C� ��P(�Oɀg�޵�"O��a$���%Jd�Ѓ&�@��"O(��BŒ�Vu�%���^�v�(y�E"O�ɳ�MC��J����2��ې"O��	cA��y�ȕ{i@y�1"OL b�Gә �FL`�͉Cq�pA@"Od��I�h.X8qˇ'{�哗"Or�IaI��P�����ذ[�1S"OF��R��`��Q6�..9b4"OR�)EJǯG\ʁ�� �%BISS"O�zT�R?0�QAi2V	q5"O.�� N�hE��{�!\,�8��"O =YЁ�8!���I�'�^�p��V"O�D� ��,{[�8��e	&t�	zd"O�A�#&� �!a����#"O|$�@��;^W��(�
X�6�C�"O��[V��M�>x�O
'�Z�˦"O���b�)�E�Dhv��"Ox#5�C� �*=&�J�n`dD�"OJ���j �#�L0LP��KU"OP9#��	xXx8GƓ'`��+�"O�p��P�K�V5���]<��`"O<�a�@T�k�p1Qe^�d�"O��(�%@���8dQ,~�����"O
�yD P�9�~��B-�1��9�"O��)�Z�=�J<���هk��ā"Ol�Jdan�"(�S�ك(f�D��"Or�I���)%T�U0稌D���S"O���K޴D��yS�`M(HU"O.���.�"
�~@�@�@���P�"O�8���L��b��L'h ��"O\8��IT���+�(C�@-����R����Ԣ�R�>E���P�q���2�D�Þ����>�yҌ�2�B�H�	I����s��B)K�,)�' (Rbn;�&��O�M��+�U���ΘES��B0�'�XF͌�1zI�ƾ�������/Ft8*@G�w�n� *��^�qO�#|�T���`����̫<0�)��#�\�'���qH�ޔ�ccR�4��Y�x-�7�D����Q��ē�n�c%#
��p<A�i�n��HǅQv�t����a?a3-�8(����fDm�?���A W���᲎ў�ajr�X���¥@\0-���[f���sW�E�5�M{��B�e �Eτ�tp\�I�&��P���+}(����"L@��-IRA7��ڧ2�r���K9"�6Ac�����bP�'�H��J��m�(ҦK�9&����iS2H�R$�6�� k���3B���?�:9����i����
y�'�MK��=!"� �4n�h)���}�'����bS"�Xi��r���7]I̠(�EF8u��j����P����AUp�'�^��H�Od���5*��6TA"g��(Xf�b �����"ȓ:�PX�BCWaQq��t�a 3.�^��CM�f�����l,�x:�!3�ɰT�G�8����*~���iB�U�cʔ$����l1P��/O�!s¤�"I7��0Ej��cx��2u�� @�5�t�ͼ;�o�	|V~���$ͬ$��a��K���(�/U�V���ϴUn�q��<u�h�KaJ��|����3��=V�����j��I�uGB���*Ea�"eK���y���,O;�a��犠t( +�&��j����hq� J�GB3fj=��Oꑞ�3ѩ�� +�m�<�^ث��*�O�pSO�(�F`�!]�5�޴0��\�J]�I[�:�͊1Y,���O�x��a���Z�,��aL6���dД�
�����@�T(iA� V>�k#G�l��ߏ\�(���/'D���FL��#&�%�C��R�M#7�Ov@(B�ۢ;v�a��]�p�"�ґ�� [ɲu��	wY�5bD(��y�O�7\�l9:e�/c| �Jn�3U��}'��ZF΁����ē74�� �	Cؐ�G(K['����Y�$�p�KP�a�ԹdeB�97��C��&���DM�#v(=z`�%k��]���Y�!���\�z&A�)i���{�.[!��D@�̩1���l��9a@�`_�D΍x l��S�? 0�A�_�F�(�r܃8��4�!�'�ԉAp�gې�J��B�G3:QA���yb˼o�21@��j:H��$�'��'���t&֗z�&aF��Gͫt5�	�U냤l�lkp&߂�y"�6��u��M�c#8-yQb�w��1s�Y5	� �'��>�I���Ѐ��I�zBE�L7{��C�	/P�,HԨ2T9L0�BQ8_����� G��#5���=E�ħ(��6ȇ?�f�I�&q���� -Sa&+e�iB�H"��x�N�RP b����'�n���:�>���HI[Nu�B+�K�\�b�E�a?���ZL�')^H{�e�*����� ��V�� ��]  � c�,w)iX"GZ��.0�e�	7���R�2O����N�2_""|r�wu�`��Wl0M��`�J[e�
�'���J��ix�b��3$����ݯ�.��`G�t��d�>�B�HB�O
�G�P����S���.�9P���B5.Z$l	"���C�-��!.2����	!�n<���?UߎJBb-5�����*8VIB䦁�l�n��c�U&�O��( ~���H�'8�I롨ތm^�̧E�P+�-_.�T� P �7�,�ȓq��9Z��� �P����2[�N� g-���R��'��=�eNŉt��1�~*�2��P�楞�Q�*lU��S1�O�y�.; 8��[�x�`N���{Ѐ�1Vw4퓅1O�`�_w�X �5[*�jfnP�LS�}�Dτ<l��)��	:-����G���g��h�3o��aQ�W$�iҷ�U�^��(�*��t�@	�2�� �ȍ#\�f��6��@��0�>ѥ��3�$@h� �ժ�_�U{�0�.l�A�K�	��Q��8<�DJ�"O6%��Ù\��0X
�c��%���3h>�����%���Y�
�3�!�#�ȨD�)	Ъ�5���b�"O@U����<Zt�xo�,Cw�d��KԅXLX���凈&����?9qE�I*n�`�$>W��H�Έ�/�\���ǒuD0u��'Z�03E�5�6L)�C�"&�P��	�'�X`�P��/�̔jF�8�i�	�'��)scC���Pٵ�M��@��'��hoҊd�R�kM�yaL�`�'��K�@�G���{U�ʌ)�)��'Utq�2H6 Wc�>����|	ʇ� �a}��� j�"09"i�AW ��	R��=1h��f::I"�'[0�ەü���c�WYcnu@�'����V��6n��s@Z3'���{2�ـ��]���v�O��1���G� ���وp�~�	�'����c��wO��� ��vy��i	y5j(iO�$�g�<Y�����!���u��Y+&��<�Ū�/��玀�_4���ݱ^��q���x� ��	�o�9�l��m�����S<t��$[4x3����#E�y"DG-N��-�tCB	%~jAG���yB!�Z��C�^���x��˂��'�v �5�@ Fb�F�T��<
]����~���'���ybA���H �O��i+�Mӷm�lQ����	�m�Q>�y0թ�B�,Қ4��W�cݢ\��n���đ�M��e���\G5�F� J���X�8b����h?�˖�F1:r�Ss�:lOP�G�zh�	#���)R�8in�C&e�2٬C�I���\0��~�l`7X@fh�#���5*�?a�%�iXʝ��Ƣ#�`��O4D��U��s���ʵoAr�f���5D��� ��6��'nR,!E�jф1D�,˃d�Y�:��f�κ
��8i�,D� ��	����� �$�|�+/D��#�$
`�XHQ�ÁNv�i�(D��9�/@��M�J� (�.z��4D�D@�F�2<�����OX#u2���/D��H�f����E�3τ�1��i�td-D���� �	K��}����<y���3�1D��@!@�A�6<U�	�X���4�;D����؆;_:̻��ž5.d�Pc�9D�� ���t�М[5�D	�!�<�f9�F"O`�'M�rX�q�  !<]��kU"OM{ �ɹB
�� �o�O�dj�"O0����1D���EN�y#"�I�"O ͂�(T8D�:�)�H�q-H���"O*���ƅ�jٖCt���`1"O�<z�� �Sr�i��æ&dXe�0"Od$���	)�`�d-�106�	��"Of��e\T��#G�U�^����E"O����h�?p�>���O{�y1"O����ܬY�J�s���?WZ��s"O�u��Lؘw�L�Ӿ!G̅r'"O\��r�	 p���Rj�p(��3�"O5��aи3�K&o8W-rŀ1"OFP;�AէQ���톐">6YX�"O�HH�O�.8��M{Ŭ�&��*�"O*��2�޻a���@e��&-p4�R"ON� 'E35�ڱ遈-a�Pm�"OVi��dߢ)۠a˃/W�lK�"Oҝ2���,���{�`� >7�%2�"O&� �%#z�uu� �v�}�"O�P7'
)q���ǎԩVM�"OفW�-20�OA%Ug�!�"O���m���G�^S�w"O���0�W�䵱C�JyBȵ0"O�A�82�|ŨR�I(;b�S"O6����K�)t�	f�s&��Ѣ�'��T�G��I �
b,P�q��U �b�-Ţ�i�'D�|�V
ډs���:��ב�d y�'�����;Cʌ�:g���$����'ߔ�3gOԟ=�6)���˝qw`|q�'�6���ޤXRpHY��I!yqJ�'&���@dJ?�t9"�E�HL�}1�'NH�C�K ,��u��@�W��,h�'����'_�qN~�s �¾Odj,���X�R!�5 d�6��H�'$YD2ڱ���է0|�T2A�dZE&E� ��=z�����J!� ,}�hA��uG�� _@T��!����H�t'�(\��>�r��^P����?�Z�p�ƐB�8����qVd�h5�Jp�A60�Ɖ�H��� �΃<3H`m:A%
#e�"8���i��y�w&I,M&�@i�O�?�
CǓ��v�K� EH��1`,0u>�O�8t��S��Q�'-}�9���z;@�F �-|�¹��'�!\,�'���{�t�O��0�a�M� ��$�C�5*�T0R�L�G�I�5ת��?��}:�O_� �4�ݽ��(P�I�"�(�!�K��y�,���4�$��g�S�NС��EK�9H�ei�D T�|��T!];\�b����ވ�$�]� ��T����@�{����0|� �_�`��MjfIէot`��p��q�oub��`��IٍZ�T%ӕ���F$�w�ܶ �!�d�b��I��(9fL�Ze�ܕe�!���%1`��Ҷ}	�aĐ>l�J�i�'�BFȨ2�U ��B��.��BI�6�y"*���x9�kU�������Ϭ�y�I��~ �v���!t�U��X��y��
��00��I:q�f蹠4�y���x��A���V�f�z*��V��y��T;{N�u��䙈_�t�EN2�yF�
g�c�	�k���c5ŝ:�y'�%�{�d�zXe���y2&�
J}��"��"fv��oV��ybH�v�����h�T�<��O��yҬ�?�D�Y�#	�6�+E�^��yb��~����vϒK�\�wL��yr�̶h[��B�`�;����t��y��S�Ag>mp�n�~g��K��L�y
� ���Pc�P�J���V��љ3"OdA�c�
��������F~@ҡ"O�x�a�ˊk~���%!ԗs���"O�E���O�)Ӧ�uWP��*O��c@��A���y�k�8X�8��'�DA�穖�H�p�ؠi:O��I��'�le�F���j96��`	-Z��k	�'DlP�sL�$X���1@ �	�|]�	�'=�Ձ1�ƍ]hH�ǃ��"���'1fi�O�#{p�a��� (�"��'0��@t��;pHVzWF�-*В�'�b�QqE�m����. '8�9�'<�����0Q��]!&�0j=��;�'�0`�5��u��4����%�	�'�D�$	]&�:�G�W�� �	�'6��b��E�nJ�jf��3t���	�'��y ���&��)���܎}\��'����fIƭw�y��խ_P����'O������P�`fH��T>���'�:���AuPi��G5I� ���'i�#�L*�����-E�E��'�J�N������09�P�'��DLل-�f�y�&\�4�Xi��'������p�� ʷ��%&T��'Ђ�8��{a�T��#)�� �'��D ՍЂY	(H��إ~�Y�'hȐ࣏	"l��!@T5Fc�ȃ�'"���#E&a��@�`S�;}���
�'I�,je�*1H�N8C m�	�'|0���?<� գ$�P/V^�	�'�X0��;�Ľ0��U�R���'_��c(^�'ܔ�J�HD�;[���'7@���NXJ��!:�D�R�'V,�r��,h����ȍ{����
�'K$]���n�; �#�J�
�'I��;�eY#9F~�Ūƶ'�*��
�'<,excϒv�NܳUw[|�"�'S��K�؎up�8#��Y9[�$M��'�<���#ŋ���Ѥ�GZ���s�'$<��FdW��̱ ���W�P��'k�!�#��3�� ѠiMMWe��'ČB�K؜J���TǥTk"h�'��, ��X?"ZZ��
��Ky ��	�'d��PΑsN �q���k�F0�'s��)���D+�P��B r�"Ob%zb��U�����C M��A"O����F�I��t�s$Q�J����"O��j��10d���� �a���"O���F&�:1���W영	s�}ذ"O� R׉Y	&���Jw��i��"O ��T��<�mӇ��
K&1�"O�5�&C�;����#@ӱn�b�s"OL�'�J�^�-#�HUŮ� "O,�j��3-�*�ֈź�&q�0"O�)�1mI \�,a�r��*�$]�"O60�\%�ֈb�o͑6�Z}���a�<���U�"H"�� ��j��Y�D��u�<�B����;&����<�`IFs�<��,؉9L�"�#.�V0�Ԉs�<�$�دG�V��[�g��<��(Gl�<Yu���=�����8;5@h�#j�<1� N(N��E yB��3pm�i�<a��W6v��r����J����d�<��E�?
� !p7�@�X�L����`�<� TIBޓr�����z]P(�"O*|Y���%18Ȍ��M�,C�#B"O��
s�F��@ɇ�E<z��"O����'ֳ*����� � �l�Q�"O �q��[�M�@��W��`��"O�i+��=q���è�.[V�"O���R�&Vll��a(5:xh"�"O�y�t
�5t,�r�"D |�2A"Od��#2	(ȅ�tN��B�|��"OVI�e �R������&�Yq�"O�Y�CM־M������;l�F@�P"O0�r$k��0q��sG�y"��ђ"Ob���B�^�^e�ƌ_�xJ�"O���a�����)��T-:<u�P"O ԠSSpk�]y�.�u�L��"OVZ���$�rQ�6�]�h�%U"ORu���.Q�<�2d��/\ݪp1b"O��SX�	����&�T�xS"O6d�䊕�q[ʐ��Q3�Խi�"O
-�S��"� !B&�XǴ�A�"O��V-^mF�ǥW�*��4�$"O���I��B��⧊�Ip�e��"O���' :bjQ�T�ֲgV$� �"O��(Q,͎�x%�$�Rn���"O���@BG,��e �#����r"Ox�"���z(浈'@k�<["O�Y��L�'��A�!�"Oء�� í�=;#��C4Z�z�"Ol0��GF�>p���+=��0R"O�9�f&�> ��:r�׀4
�"OL���!H�������8(Ҍf"Op��'�^!F5cQ��6��b0"O�ı�fI
Z�8��Fk�
��S�"Ov9�FF�D�0�x"�K�w�pa�"O�� �F ��mR'�W>/� ��"O:T�e�@$����(��X1r�"O�<b31�<���
��,�q�"O���w��_(�-�n+#�D��"O�p�6�I>�EG#�UB(�S"O�)+���e��(b��C7*�BA��"O��D�֔!��̚W�H�n���"O6A��81|���lH�%@���"O��㓬V/�x� P�l�8UҖ"O��{dF(c��k��^��<*F"O~]C��R@V-�B�j��"O"���h�4ʈ�.�/$ɰ��"Op-b��͖\:0ԣ޶v�t��"O0��ց~m� �#�C��)rB"Ox蛀�{'N�p���x`��"O�y�,�+.��BP�&Hp��"O�yad*�/�%�7�&(El�S"OxUIs��N�
L����eA8�"Oza�G�p,�2R���YJ��%"Obq	��J	e��e� t���R"O�(ۧ-�	��
u�ɩM��t"OB K�U�JI �U8t�D�K0"O@,ȃ�Ep��M{W��3}+�m�"Ol�
��Ә_Y�T�Rʻn��"OL���Hif�M��Su%�
�"O�@q����i�e�� o��S"Ohe�V�@�DzpI�(C8t5��"O�	��[�[�8I�cbXWZ�4r"O�H����31�(��#��DO8���"O��M�E��p���C=f�mZC"O� �t����l�8��r��=C��ș1"O�`!'�E�\�P	cUJ��:�R�q"O��[�� �u�ico�Q�"O0͓��C4wy�qS��\9z�Uڇ"O��M&9aʥ@qI�ZaTa��"O�Q�Eƛ b"	[!��S/���"O�!�gL��wha�#$?=&��"OF��2��W�lX�7/�2F0 �8C"O
��uK�X4����ښm(|�2�"O��zE�ۺ=T �#��.�ˢ"OF�i�)^*u�%�2,Q0t�x��A"Oi*pLT��{k��\�֐� "O�H���@�[����C
6 ���"O`t�͌3e��������ݐc"O��x��C�k32f'F�����<W!�$��Z���p�쏬n,z����6zB!򄚃��ٳ�hR�On��Sǭ,'!��T�F�@GlV)SX(�@WNլW�!�y�f�A���w^Tۂ��>Xh!�DPw�ʵ���z�!j�Jh!�#��h�g�8��&�08!�	%��Mڕa��qr�E@*�!�dY�t�,�ZQ���M��9��ZL�!�D�.��\ñƨ@��&��ue!���\�D儶y����&ŽLU!�Y#		�̓'�Ŋd���/ܒvQ!򤀀s���<�R I�{>!�$� v���ǰU��� 6!�D�*l�0��ㅖ�b�����Gġ9�!�$��.`Pq��⑳BƜ'�!�E	tt�1�Ɨ|�� ��==�!�
�r���rpʜv���geg�!򤊻*!��K6 R��p\!��<@�!��,b�dDiqD�c��ȫ�o�%Q�!�d�";����z���*�n��[�!�Đ2=b���חZn�Ȓ�	>)�!��YU�R�jO�q��	����f�!��G;������l0�CdԿS�!�D�&{��لm�.��@`AE��Y!�䇋:�h��j�=U��D� ^n!�$ݖC�j��&�P�,���e�&1!��C�]��I�a�Y�]��h�D� f!�D:b6����|͜9T���'�!�$�>ܺ宇5�T �ׯ܎Y�!�$�����B�h�{���`���.6!�Dʀ�,�暵�&}Ag�9Z7!��]�
I�H� �X�4��y�F�#\�!�Ր���1*	
?���eC�IO!��@5/J�0#q#A0X�R �6"N!�d�	(��ڤq���2lI!�$� X�j��5AY�p��܁��58!�$��AW��pq^�.�R����C�,!�䌱I��q��KW=S��TQ�K�K!�$Z�Y-R����YԦ�����K!�d�0!�JAq�#-����I��!�
v'D��jH)E܌�4�ߚ$!��x� �  ��   (  �  �  �  �+  �7  :D  O  wZ  ;e  �n  �x  Q�  -�  ��  ��  A�  ��  Ũ  �  J�  ��  ��  D�  ��  ��  ��  ��  
�  p�  ��  ��  � A	 �  B �" H* �0 �6 �;  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�kL���>�b�fX�H�ҢS,	aʄzՊZ� {���$$����=-jܨ�U��d�&m"�-�Px��$�#L�V�"��UOJm��&5A�zB���=�r첃��d34P��Ɲ64!�� -^�����;��)7#�	.!�d����i�#DΌ!y�ш��Z+!�$�!W���Xd��1w$���Ȩ|�!��b)『'L� D���%����'qe�u�Ѕ;�i�ʈ:$rH��'м�*@0Nx��6&���� B
�'ƥ�&@��{[��KC��.�p�	�'����b�<P`�2��%����)O��=E�d,@"W����&�&|l�
��9�yb��-rτi��ۧ�nHb�ّ��'=�{�+^}WP��L�	[
|q���ybG�q�HԀ'��:��ҰO�$�y��U�=/�l�5*�t�p����0>�L>�Ĩ]O��m�7��<b��C	�I�<��&�)�f��H'.�A�f�p�đ$�M�ד.�h�8R�L�G����r�U�B�	џt딬��E�����LA�6ʖ��w�+�?I������ɼlV�Ǣ�4�bL��NN.�x���3?�*O΄
�],W��A �O�*RP��r��`H<i4#��U+\�{��8r��U/ZL�'O�?�����6s#�(An�\(zE�v�"D�,�Ì���X*�A/7|�v@ò�'^ў�� b��E?�*����Xx�<�U"O� �I��?J�L5�&��#8�Q��"O��B�SzTf}ÕMě*%�t�f�Oԣ=E�d�O���:��C>hm`�
�M��'��I
`hF0=sؘ��<ht���$�H�O~x"bˎ�V��81�=4c�s�'TZ\A����xX�ɰa	.�ICH>و��	�I�dlK�A�
�$i���iW!�$��S��xᒧ�k�2Cw,�w%�'�R�'I$�,��G%<�0V ��ty�,(�'��CvaZ4j�ʀ8�N�r�|k�'����ݏ��i�%�L e�x��'Rv�ٔ�O��n��/NI_ �H�'��c4iծ^���ԏ��p3h`��}R�)�)��EP�a+RE�e!�xc��Z�*�!��.��LK7�Ke�zg��:c�O6�	m���{B
Q�T��m�C�G ���g�+lO��𹰏�;,-
.�D]��� )D����f�3>���!4�湛�k2��Q���O���xR�С6�����j����'t����Y�p�nhBQO��Lg�Q(���I�'��I�	�t���Pw�6�[�a�;t��C�	�n����nQ+FlZl�b�B�-{
B䉑0Tdl��kG�R�"���e�C�	�o9(p�w� �HR@�q&��X�B䉱�lDJ�玟\] ))`l�Y&B�2!�NQ�������@��~�ZC䉢+K�y2���-�h`��`�	�B䉍U����i�!�l�	��ɒt��C�ɀ\�2r �\�\�f�1	��C�I�
�!9b%�;L��B�N5n�pC䉸<��@�j�*'>Iz�/��8 <C��8Fr|1��K�(�&9�W ϚI��B䉼%�6�	��I$2P:��C�ЛZ��C�I�4sNQS�$j��ʋ)H�B�I�m�<�ŏ��'��|�dl�"N�B䉤5P����!��xD��p��B�	 2'��gJn��qh<f�B�ɅE���� !ٚN��a�LÅA��B��u�DLY���[�Ysg�1Z����6���52��X�lfL�0�i�!�DG0�D�����
X�V���4yQ��F{*��@�DgE�+�  ���qɛ����y�鄓7LT,�֤��QR�͑���y≄�.Sv��"n�=B�1����?�y�#T�0���K7	��!u�
�yr�)����4*@̰kt$���y���>	z��A�H��K�@}�F�ҁ�y��P�Ċy�piQ:X$��C��yBfU�, �`�� �=]*P)ir���ybK�4�,� �b�^�˖���y���G��3�΁ rI��᫞�y�/�3���D�5O���*ο�y&�"DF�)�S�V�"5�"�-��O�"�Wς�O뮑�2*PZ���R,B�<	GJ�甙5͈h}�\pf!�B�<Q/�B��R��`��g�@�<i���kL���ᑗ���RdLy�<��gH�/��V�Ch�}�V�t<���,�X�	D�ױ,��M�v���Yu`�ȓH�Ƽ�ʟ5DA\�P�L�t�̜��l��%�G噙G���'Kó4�L����~!`DK<+�Y��҄nK �������A>yN���+р�X���J �����U�0E�H����B�����S�? Q ����k�Tu��Lч'G
��s"O<���# �Eʌip���?(O�H;�"O��r��SWT��c�ЂRN%�#�'��O��a�@�#7�F��r��4f��"Ol�a$�C�-���)@R)]��PF"O`�t��_จQ$�N�`H�-R�"O�@�O�;Zd���JB�u"OV�H�␎K'0�bf���ی��"O��x��)����*�Ux^1G"O�y�!k�	�:�Y�����"OB��դ�2-���"�Q�f���3 "O�V/+�-��d� y�V�K)�H�<�CڇP��|��e��!�¼�Pf[H�<�D�ۋaC�ʆ�v�L�ssFQl�<��LU�V7r�tO��0�)��Wk�<��J�Anv	�0��\)�80��d�<I҉�?̆y���X����;�"{�<I���2�ҙH0hX5LhB���Ns�<�P�ֆ$]Z0;�
N����Öh�f�<�j�>�nMib�K�!t>�c�c�<� k���%���
�:���C�X�<�T�)}fHED\$9,1q�g�U�<�&���J�X�FMofa��Zf�<��\�VF���AX!,U��jk�<)qA͉����D�M�JR���g-�e�<�a�5�F�i2�¯`w��Z`�`�<)�>���1B֖hޒ�I)Y`�<q5퇸_��E��*�?���f�_a�<�.׼+Mh݀cI�"��TQ! �B�<����� �P4�=0q�$CA�<���>?�~�*T/]��)	�-�}�<�rdJ}����f�?T	�X�#*]d�<�GLxS>肴�V=c�D���g�_�<��+I������^�{3t�P�J\�<!�2%L� TI�v��e�t�~�<Q`���0s�%�e�K4>�ꐁs.I`�<a�뜂2|
�1.V��(Y#M�_�<�6����&����X�$:�v�u�<����;T}l�%�j՘x΄H�<�P00x؝����m�p! �'�F�<!��֭5�
�V���
���I�<�r�����S�I_'O@���s��C�<��]$|C�tsh�8L��au��|�<��!��j�@ r�g�J(V�I�$Or�<�L�w�P ����(Ig�y�w�o�<��� ��A�m�!x�n�@#	e�<�ъ�0s��('d�(,��+�Bh�<Y�bʰ.��U��  }���SE�z�<��,f��eKŉ	4X�0�v��l�<��ύ�x�|�`i]�|���1&�d�<�U�Ք]�x�K���̼aԪu�<q6)��\�f%C7/��!@�K��G|�<y I�k�h��)
U(���$�u�<��e_-SF�S��I/���㧄p�<tI�Q�������<�xeQ֏q�<���J%#3x+r�ج<z9��LH�<���_0+�H�ү�2�c)G�<qCmW�l$�*�KU7@�@�s��]M�<�Ri^	>N�CʵG�N��A�<���oRz� B�ݼ�z�0	�F�<���XL�1�w*��9Ǻ%IC�Zm�<q�Ĉ�vo.�\,Y�u�g�M�<ё�Q	���:C΃ :r�@ɴ�E�<Q -�k�VpSC`�$Y;�����<� ���6f�Ni�=;A��.;O9��"O��B잏Z�8�pϓ5��ؘ"O���FE� lЙ��͎�u��ɱ%"OZ���^̕�7/�>�\��"OD	�W��<�^p��˘��$�+�'��'��'2��'���'���'��8����=
Z�+�jm2Ε;��'wR�'���'s��'^��'c��'y���T�;5;��ރ`L�����'�"�'���'nB�'��'��'� �k`��l��Y�j�Pj [a�'92�'���'�R�'�r�'2"�'o4q���Tu�ā����6#��'Wb�'���'���'��'p��'_�,����Y^�����sd��q#�'lR�'���'H"�'V�'2�'��kA �@�������+��%�'<r�'lR�'���'��'kr�'sp����Ԣ�޸���ѲB�&�?����?���?)��?Q���?y��?���Ԕ:�R�r���'P��XvA��?Q���?���?����?���?	���?!�g�%��1b�M�S�ĔJ����?����?���?���?���?���?��Ʀ�T�H��7D��{$�V�?!��?���?����?���?)��?Q���-*\41�İS�<qe�S,�?Y���?���?Y��?����?I��?)Be�{��@�G�kAr�r�!�3�?A���?a���?i���?a�4@���'�d(~Pt����]g���C`�:�d˓�?�.O1��I��MSB
%+I����֘)�����
=��@�'$�7>�i>牮�M���q��UAf�#k=3ŋ�.<�v�'�N�a�A͡���+<Z`y(aH����{�d�9�iL$5�@��M1Lj�c�D�	qy"�ӗK:r�AŎ-���$(<_�q�4����<��t-k��NC�BašâG$�=XF��EߴmZ��MC�'�)��d�䚱�n��p��G_z���k�m;x���)u�| �OV�N�f!আ�k�����'��D@���j"(�фd��6ޔ�'��IR�I(�M�@��g��>I���Ut�e�cH��h�+�bJ�>��ik�6Mm���'fh!��/G_6�T�@#��x�O�l�)U�#<�E�R�)ک&D�])P��O�<XG��/@b�)�G�'n��|⧪<�-O���s�`�2EF���H�e	;` B(ɵ�k�H��418<�'��6m2�i>AC�H��,ƍ*&��o�p�ܴݛ&�' ����(��A�U6�	D���8`ܹ�����+n�	#Q*�X=��<ͧ�?����?����?�$$� *�N黗eR��^$s�����$Ц�㶃؟t�	ן��D���'���N : f@�p�Z:9<��2'�>1�i�X6MD�%>)���?Ba��^I�����BqY��Z�mʹcL���n~���垢5�p�ą0^I��IZ?�ᥣ<���L]:�*�n7*�@�c�-��?I���?Q��?�'������V ��� V�A��X��%���s��K��h1�4��'-N�!/��C}� o�;]��Z���T�9C�替���`w��*��������A�hqj�gyB�O�v�X�~I�10�$p'��&���ԟL�	ԟ��	���Ig�' �|}�T'��M������)w�-�'���l�>�Id���{ܴ�?�(O�$� E��L�M���D�tX�A���'d6�Z�����0 ��I}���	�di>�#���Ԩ�,'R���%�ԂL{flJCᔴHz�'�h�'���'FB�'ϰH�F��45�8�p딁|�E{!�'��W���4mX]�/O~�$�|�g�rĲaY'aZ|тXa K~�i�>aB�i?�6�\��$>��S�0�yƇN�#Ak� 
�p ��Q��n����gȄny��O(n�������'ܶ�yk%׆0�@k�!L�aô�'��'�B�O��0�M3�� j��LX��V�e]`(��kK�=�'��6�:�I��������Z'-�!��4Cէ��� � �+���M;3�i��t�� �yb�'D��3�ԆF�6L �V�X�v���T��eJR�\�i��'t��'X��''��'�S�>h�ib�A�c$���aǝ\:0�"۴NM� X���?�����'�?���yG���A#�2o�=-�4Mð`����6m|a%$�ڟl֧���O��$�<9�D���'89�cFʯj<,ͩA.��ih�'Z��QD�_�&⾨�Ǟ|b\����П��r
�2I_�d(�ˉ�����L̟t��ӟ��_y2hq�|�64O����O,� AkPN"]�&��X}�롩#�I���dצE��4Fr^�<Z��Rh��Dz�.��T�|�B��a���	�'���q �Í7L�'���531�(2��':~ �5�#%�͉��VB����'2�'R�'�>���I��@2�D�"L	�*C�86��I��MӇi�@~Rdv���]8^EF�a�L4cc�Q�@�JN5���M%�i�26-�]��*�8O"�DT*FQ�"��.j#<��H��]�����k�x����䓟�D�OT�$�O>��O��� �(Z�|{��CI��"����?(t�|��含����O.�I-�I�dP &�׭I�.@*AIMS!
��'�7������ħ�:��
4���ǩ�h)x��`2%�2p@@�'�8(�,O�`J3��2�tj� :��<!��6)PX��3 �/|��s,R�?���?!��?ͧ��D���*� �ɭ12�A����J\M���ڱ\)�I��M���>�"�i�7-�ئ�B���9'͊�+���$r�DHs�A�'!%LLy��m����1Gj�L��M8$\�͖'��t�`�� �	җ��4���7�rg��p�0Oj��Oz��OX���O2�?Q��fm�l�s��cj��s���I՟���4Z��A�',�6�.���#D�̌�E)v�T��'6�6<�IH}�d��Po��?y�eS�I/�	ן�p�O8H�����ӷY�H�{�Nq\�����)HJ>I&��'���''��'Ҽ �
���9`%��7 ����'��T�HܴFivH��?������/]}nY�b �$$�e/W���	���$OƦ�޴ZW��T�OZ]b�Ǝ<B@���G=y1��	��՗97��n�0m��?=CQeܹBf��%����C]�Z�yq�ã����6�ϟ@�	؟ ���b>Y�'?\7M$��*C	�r:�c�+O�E�����C�4��'���aڛvfثpM��;�Gŏx١�fE&7Mצ٪��έ^v���ɟ���U'Y�P�u�JHy�A?�����m��.��`�-ў�y�Y�����0�	�0�I��O�ƌ @G�q��Qҡ	�$�!$Io�X�@c�<���'�?�3��y���4P�ȁ�m��z}��`I�B47�ۦq����4����������/��L/�K�\I��.ăL��[�P;*r�D��x���YE�K:g�֓O���?	��b_^qi�'�����u@��'�����?���?�(O܌mڸ|%z�	Ɵp���A�}��ܶ%�Nlsg���%�ڰ�?�V�|#ڴM�V��O��v�0����]r�qg��q�PA͓�?���	xz!Kd.������(p��8T������3�)�3;*��D�ۗy@����O����O��2ڧ�?9-3����N�t��#;���	�M{��M~~���6�:��P�	r�T�I ��0(�P��M�!�iA6͝�zn}t3O��i�J`��	��;co^6g�0h�����ju�6���<���?q��?��?����6]j��F�ڰ�Є�<��d���� v t� ��؟&?��nr���7��#*Hڅ���e[�P�O�DlZ��M˱�'��O��d�O��T���Zr"p��kO�q��Ν�C�'���N3�ӥ��(N6�O�Ӳ7�Y��9ڰ������T�p�������ɟ��Py�OfӬyڧ:Oڙ�J�M�v12�
@WrTڤ3O�Mmn�Rr�	�MS��i��6-�73�,���H������u1��@�)߾����O������5 � �s�<���	�kй'�P��8�t�C�U;=��O��d�Od��O"��#���	E�yɈ�M�ȝ �����џ��Ɏ�MCg�X`~�Ew�r�O\7��:|�aDۓ
'��[����?a�OhmZ;�M{��, ��Ј��<��K�&E�r�޸=�U��m�5A�*�����_]$m�B5����$�O:�D�OD�D�{E��R(��֝�A�9|d����O��v���a'�yR�'�_>��u�GXT��� 8�]�'�d�XK���~��I�	L�S�?���k�:l���P�N���
B
H����wnåF0�	�'���^�1��*��|�gϢ;x쪶חl�ꅑ���me�'v�'����[���4i����b�'՚�b1N�,K��D�����?i��)F���x}"�o��Mj�I�p�dq�`���CG�����ܴ�h5�#��<���9�R8Cr��68�J+Op����_�]r���P!��i35O�˓�?I��?���?������P-^0)���n0�eK5-�J0�l�5&��(�	���a�S�x�����3Ņ Y�t��f@/�F�rE�_7�Ʈg���	c}�O�$�OD�׭��yb�H�Y���a��<�
��$�&�M4�� l�q��� �T�'I��'+��'i �#AH�v8�Щ'/�0�jm�1�'�"�'��Z��4Me��[��?���tsx��S�@�&�Ҝk���96�-C�R�>��i��7��ßX�'����P��P�h)IL�S~dTڙ'��� H�Ġ�H��I�?�s2靂�"	�	�|�:# ��u�r� �݈�<�������ݟ���Q�Or#ʉc�R�����v4q��$ںw?Bf��9���O��ܦ��?�;7�,a�Q%�ș{�i#�}�F���mp�� nY�.m�g�}���I@h��@��t;3�Ћ�!�(HY�C�L�\EB�0���g�	Oy��'X��''R�'��HF:^l��J���.����A�`��ɱ�MCwD]'�?���?�N~���+Z�Td�;b\%���O 7�^��R��2�4��f�OV�����v���i�z�H!��ᇈd,`���a;������<ad��r��问�����䋡L�@�X ��@�E�<҈���O��d�O��4�p˓�քJ�k]M!S��1Gз*���!.>f�bjz�
�D��O�l���M���i�@�6%�)�8�K�M�������Ǒe$���'�B�;dL���U� ��	�?�
]c�xrO�"3F�# ��+⾉�'���'=��'���'�~���Τi6�4#������ ���<���?͛���T�'!�7M/�dH�L�X����H�V�.@�����	I}rElӀm��?����
��ן��eW�'����ba�y�DY Ua�j�X�+!b.�v�&�̗'���'c��'�L��.2*E�� ���/Tb��'��W��Q۴D�Q�/Od�D�|�
	�L�+����^���@��y;���M¼i�*�D'�	��4��e��F���c���A�"5c��9^`�э�-c�.ʓ��&'U)����K>��"ߢP���a��;Uv�ۄ���?	���?���?�|2,O��lZ
,�\)��+�=��� ���D�lҟ��I��Mk�b��>���i`�2���	v�`q.��_鮘#�j�l}o�O�t�`�b�4�ɤo�f�P�@K��~��� ����%�"��lɴ��
��� Q0O���?Q��?���?�����i>7F��P��,,c�i�M�J$l�#���	ğl��L�Sğ�����a�:
�P���T�<|<�h�$t�FMu�����G}�OP���O�T�VLў�y"��8Y(U�"oq��{��?�y�7}�ta0u�I�7��'���@�ɠE��Uj ��#��1�%�1�� ���D��ԟ4�'�(6-�Ġ��?ٕȅ'}v��dE�go��������')���f�dӚ��Ix}Z!`�u 
*| �0+ T�g����y����Ф6�d��\��~Zw��Y%a ��$$ ӟ0�â�I���(M�d��ş<������I��E���'5��c�!v@�.�$�T���'�"6-��7E���MÏ�w�ܴ9���g�n�8����8�'��7���	:�4(s���M�<i��EG��ɴ%�Nh��7�F�7]4�$�
^�^���/�������O��$�OF�d�OR�����)Z!Dٜ9$����"�?i���jj�V/M���'���O\�S���k�/�7y1R}����*�H7MX&���Ʀ}��4�Қ���O	��Ԭ&�&LK�!O4Kl�%�;l�6��W���!s�I�$!��o� 	ӆ`$�(�'�J�(wMsڈ�3�O?Cð�(��'���'������\��2۴_ؤ��r6tK�
�0R�
 cO�����X������k}�t��o�:�MC%.T2)�J�2"#�'j���[��*3�q�Ĭ�<i�஑s��X,*�h�R(O �I�×�@�r�*qΊ���S�(��<!���?���?Q��?�����X�:|�<���D+"2LG�)�y��'��`�(d`v���2�4��%���k�ʘ`��ŲQ�2~���#��'<����M밺iq�d�,A�5ۘ'<"��R����t��T�B�;Ť��a"~� ���q��$I�|�S� ��۟D��ǟ4��S�'�6	3I�s�J��������Ly��`Ӝ@Q9Ob���Oʧ|�&��08W��)��E�jy<��'��J(���sӚ��	]��?� gA 0�]i��ω'oZLx j�rf��y�G4%���'�d�]֘p�f�|�)D0I�� �5 �j2aɡA��Y�r�'�2�'(��TQ��ٴ1���G�!Q8���H3>욂aVl~�u�T��s�O&)mZ�,il��d���"7H &�۽U�DAYش ��v��u��I��'m%��5$�D�f��n��ep<	��Ɗ2f��b�����'@�	����Iȟ���q�h�O^˧�4��*�P6�atB���N!:�i�@mS�'�2�'��y��u���=aZB�n�@��a�	p���n�3�M��'l�i>����?�&�ѽ�^�	�S����E׉i�4����2��I~-��vL̉[��&��'���'��D�$f�9ei�eؗ�</"��r��'}r�'��V��ڴ������?	�tHG�8<)��c~�r��ʟ�'�{�OP@mڣ�MS`�'N�ɓ�X�9�gV:4N�)�!΋����ן�Cc( ��`!��XIy��O{�4�X,�s��m����Qj&��zPl?) ,[���?!��?���h���J��BtY%�җ7��ŀ��	8r���Ѧ��g��8��	�M���w�f|j0 �(�BE²m�8o�lx��'ú7�O���4h��HJ ���<1��r�T2х��P5t4�UF�lCJ��H�jO`h�`������O����O���O����x�~��U$E�8ݪչG���Tʓ�։θx���'�����'C�m�V/!��8���H�D�!Dc�>��iH�7��'>���?	�&��*��*��W�L��(�r�W�i����Uryb��qrݹS�
?W��'�!t��xW&τ�d�Ж��!T,��	˟���ş��i>�'	�7S�d�\f���r T�, �SDM�� ��Ц��I`�ɰ��$��	ݴB�����d�btjq���}"�;��Kg,��F��y���Ŭ@�\m�Ŋv�A����񟼜�1`.����ׇ��$x��[�VtY͓�?y��?y���?Y���O:<y�L�%R,S�X�Fj@5�'�B�'��7m[����O� l�i�: ^�[�׹
���	�gΠT������W��i�4�*������7O��� K>�'�YC"�yAâ݀;r �PF�\�8ږ!5���<I���?	���?ir���3 ��F�>��x!4�P:�?����D�ʦ�8��^yB�'��ӱR�> kf) i�v�a$�1���%��	3�M;�iʘ�D>����z����,R�h�!��B"*o�X���#���B�&��t��PL>�ۏ00��zC��B��H���[$�?)���?����?�|�,O�En��kR�e����vjH	�"�]���隑s���'}�6�0���������uDT( �4%��qd�aE�ޙ�M�i�l%1�B�y�'��<�p$'�ʅ��Q����l������f�ћw}�<��i�\�'n��'��'���'J�S�q��dPQ#T0��Zp�G�J�Z��ߴp*B����?I����'�?�@��y�!V���p�\3�����S��|�j�lZ��?1�O������i�	2��{6O�a��'I�`�<�c��>ld�a;O�TI��$_l�Ɇ�+���<���?��΋�������6E�kwb��?���?������[!��ݟ����lV�"/8ze��.ѐ)=։b�GBV��j��	�M��iA����>9���uK�e�Q�&(�Y �cQ�<��n;5�NU:\,h)OH��K"s}X�X���O���a�h�A��h��HÜ����Of���O����O�}��,ljlYs"��?�B�p�AW�>|����>>��*Zl��'.�6�.�i޽��(7<���F3^]ӓ�s��R�4 '���d��aB�L�E��$�O杸�E�]��Mp� ��+u��c߀x2#Z�L��� �2��<����?����?����?b����V�Q��/E�T��˟�����9*"�̟d�Iğ�&?a�� ��d��֩(�$J��:��	�O��mZ��MC�'`�O���O������ m;
�zC씔+��uSќ?�n��U�ԛW��&q�\�5 �N�fy�/M�]@4]0��1[4��	�M�t���'���'��O[�I�M�%AG��?��!U\��h�1��&��᫵��6�?9ֽi?�O`��'Ȗ7��ۦa��4/_4h�6��%x� 
sD�9KܲE{COL:�<���?��-�#R4��Vl�%����x�14]��"e׸/����)�z�]̓�?)��?y��?��-��j
�<(�xy��L� ��ecX ����O\|l�:��ޟ`Rٴ��XK�[�!�U$ yTIǶp/ҹ���'�ɓ�M[��i��$�	J$P�'!�h	#N
%���>^�4�S�*g�L���&G�2u��|_��������	��x���!���{o�Q��N�S_����O^ʓ4��ƉÎ,���'�bW>���@;a��-�pbа�p<�'&?�S�<�شr���n�Ov����C��0�ɠ���j�\��cBƥFt$�Fio&D�s��<1��uf���p�ڝ��P��B�bR;.v��F�ņ(+ m����?!���?�Ş������A%�8�e�1�ѝ~�����Q�>(�ܛ��$O}��n���M�.@|T{g(J2d��ۑi���y�ݴg�L�R���<q�"���P�-��+���,O4M�4N�`%��:����K9REڳ>O���?A��?	��?)����)Ŧ��b��H���7� >nnS*����K�s�\���K�ß�Q	$o�
V�v0��Ĥt�V�v���Iu}�OM���Oi�x���y2��φm��b�,qfJ�o�;�yro؊-��� q����'��I�4��4hJ���fC̅l�B�)�y�	ȟl�	Ɵ��'>�7m6�4�d�O,�d���AI���~,�	�LU�S;��t�O4�l�M �'A�I�g��5K�MB2�t����D�O�lRdĄ�L�\��<Q�'o8C!��?i���S-�9	7��R�z-�`�K��?Y���?I��?	��i�O��eа5��Ӵ��A� ���A�O2io�t���y����4�(���K:� U"�n�E@�cU;O0�nZ��M��i� }��bM�y�'m��{Pi��f�� �r�)Z�;u�Z?���q�F�"�'���Ɵ(�	��ɟ �	t̐p�aF�y���H*��%N��'�7-e4���O���!�9O@�S`�ݿ;;��HA��W{����r}BjlӮ�mZ��?QN|R����e!��1�����$�r^����Ί&ל����&��ɶdRuC�ˈ������_�w�N�}�8�:�J�H,����O����O��4��Q����־�yo@�y�Wp1�R CJC�
� �����Np}�Dmӌo�?�M+A��r� �F��+�8�ɔ� �RV2t�b��<q��H��*�q�"�{,OR�����cU��V� S�R�Oa.%ˢ	��<��?����?���?y���h�*=3�MR2MW 1JA��m���yr�'�2�w�މB�����ܴ��*t�(�Gߪv�L�5�(^�8(�R�'��I��M���iw��	ܼd]J)ș'�҆΋֊T1$�[.>�Xz�k��DT��%������2�|S���I�l��ƟxoU3�T]`���C��AQ��G����	Vy�dv���d������?A��}���
��Y�:�&�:B���d�p�OT��>�M��v� ��*�	���N�1K��U��
���4�#J	7��1�宍�R (˓��a��5�h �N>���G_T����G4a���a�a��?���?���?�|R/OB�nڊ_�����f��yD�]r��2O�m��<?q��i+�O2��'[�7-F_0��@ׄV�n��M�ֈ�&ߺ0m��Mk��C�<R��̓�?��� )�v�sV�H#��$� J�dy���:���v��� ��ɧgC�m��qJ��؝`ih3H�fNN�9��.:�m-�>9�s���5V �g�<2���6�9�v�<�d��H��}�dĠ�B�a2 6A��a)���00]~\���V0/ʱ�(�\��ݣ�f���2E��#<U���A�#�R����E�,�.!c�d�$VjA�`d�g#d�j�l9 g��� &�zN0�w�@�0�^��0g�.~:�B�M�vH\E��C�5�X����:�.�yS��Ԧ��	֟����?�O��9b���+�5��̩7k�Sjp	��i��K�'�RZ���[�֟���"~Yh]؆�C>a�@Q`�B��M#���?��HyT�{�X�\�'���O�@�	ݨj`5���Z,_�"H#&�io�'�� ����i�Ob��O�`�G��/��[ �(PI�����q�	6i�z��O�ʓ�?�-O���Ɔ8�MnHX��[�V�ի!X�8�A�o��'���'�rP��U���'��k3ڒQz̛ã��9&�h`�O�ʓ�?I(O��D�O��$���LB�l\�)��t�1H �oG���P8O��$�Ov�D�O����<1W��Xh�iǒ@���@@5_��r��0!d��X���IOy��'	��'�좞�5�o�(���)n��)�X���M+�M�Y>�����?a-O�<���T�D�'�`,�re�,l���5�E�Zֈ9ȠM{�l�d�<����?���+0�(Γ�?��'�< %oG!@<J5y����p�4�?Y���$�΍�OD�'E���`&0�����<[����M� �@��?���?�RAu��<�OCv ��:Q�.5�6J�
*��hش���3O]m���I��P������HYE)�(`4l�%Մ4kN,���i��'�A0�'7�'�q��<H��L��b�(�-̑9V��0S�iTz��ňyӚ�d�O�����<�'s�I,Ԁ �	��)ط"��PҔ��?PԵ�5�iDm��'���'Jx������$pЀ�'	 �:0��l������H��	����[N�rݴ�?���?��?��nh�"f{kt�+`��2P02�n���x�I1�r��#k������?��*��%+�$�1Bf���聶����'�T��)�>�)O��$�<�����6& �KiD��
A/Bo}�Ҍ���O����O���|�ጞ���!��f˝0)\	�Qj՜]��i�r�'3��'�|�'��d�O�X�$�"p�$8#�A�=B�b��e��D�O��O��D�O�ʧb�F�S�iqD ��*Q Q��1l�$V�a�xӴ��OD���O`���<�s�@=�'R�$}Qt�ۭ9�~4��h�?$W¸�Q�i�B�'��'=�ə� �SL|ztM�,v>�-����=h�8҄��,-���'6�'X� 4�c�8�aJ�@EZ�J! �c�@t*�lh�����O�}���p����'n�dH�a�|	2���ʶa�5˜ �<O��6R��Gx��H�����Pb�Z����t1���i��I�l\�0��4"��ϟ�����$��Xwx�A��ܗJ��kL
()��[�hy��=�S�-N¸PqOB8h\���fԭBJ��lZm��M�4�?���?I���'_��zc �Y��	��|c� ԣ ��6�S���"|��:��-jR3�ڰh5n�$a�����iZ2�'�ҭR�qW�b�t��]?!��N�!�L��(�&d����W���<����?Y��;��܀AL�H��Y�#R7~��	7�i5ҋ�;�pOb���O��Ok,�|�튵�̔'4�Q���G �ɖd.tb�t�	���Jy�n^ 3�e��dW�xpR�nX�{ĞZ�m;�	џ�'���'b!�LN	iS���A�_�V
|rE����'#��'�"U�D��a���
���	��뀂k�l�{GD����O��;�$�<y2CU@}��9B��Mȕ<dcg�L����O.���O��{��<���T���_�U����OB��Q�ߥd�7M�O�O��s��>駭�'_B��8��.���'��I�I�Е' 8��ւ3��Oh��ܧe�ns� X�́PCo�^�'���'�@���T?1ӡ�ݲtT���CB� @0���oӶ˓�>0��iv��'�?���,���0X���"��<���Ŧ�v�&�<iRMW|���O�4\�댕zn ���߮}�M�4'�v��g�i���'��O:�c�(�2AH _���ha�w;�A�v�P&�M�B�Us�������WL�Bb�֔��a"��0V�Yn����۟ �5nK���' ��O��P5�G5�:��Q�O�YFD�����+�1OL���O �d�8��s5GOX�0-�0�R&���mҟ��&��'��'��i�q�dGC�qnN�9�k\0:�F�"TϬ>��j]g��?���v��[��ā�>�~}��E�h�b`���]�8�K<!��?q���<�a"۽7����C(ɔ �R��-ʀT��H�<����?9�����i�|Χt��K���+1�hu��aV���M�'�B�'�R^���'`p8x��8 Q�X%�V�� �Y��C�X��I̟��Iby�H*<�f����@/,���U퇊:j�l*�)��	�	u�	fy�G����'��x�ː��<,P!���A��ܴ�?����Đ/��&>u�I�?x]�隤�y�/W���$@ƌ�ē��
,U���Zq"p���Q����%V�L���mkyb��0+�6�_���'����+?�0��Y0ę�F��."�bq�cJئՔ'�f)�����ɩMG���J�<.F�ڇ�,CD����2vIR7��O��D�Ov�)�j����:2#\3(J�R'L	Q2��U��M�ej�a�������B�pY����J�rdR1I�96RplZΟ�IϟxoG����?����~rO��3�z���D;6��D� ��/��'2v-S�y��'c2�'�� c���y�3c̮$����b���$8k\��>	�������+N�>Q �J/w��L�r�WB}��Θ'��'H�W�����@��h ���Y:L� ��-��}B�'�'<�	�Zkr����9���P%9x1�;�	ퟀ�	�D�'1�튑�l>�q�bR2w%1aP�҂nBh�! ?��O��OH�z-�]�'���F၅*h|�#�!��v����On�$�O����<��H݌�O&�mі��$;Z^<�W\�C��� ��s�2�D/���<���[u�[�t��!F$���Z�&=�n�ş��dy§N��������tyd��B\P��� ��%)�Pd�	sy�ų�O���xr�O�!d��"�K� �6�<9`k@�%[�g�~����������!���)�������i�4ʓ:�.5Dx���#�f��`A�O�75XZ�r��\�a!�$ ��oi���D�O�����l %�`�If�D��pg
f�bA���I	n֠li޴8�&�Gx��)�O�d�!��-!�\ږ!�nN������ןL�� Z�ڐ�M<����?!�'Ά��ۘ5!����P=J7F��}"@��'���'��GH���qc�)s�8aчE�q�:6�O�h0�N�G����D�i�� $��1���E�̧R�Q���uf>��Ɵ���'�:�S�F =��v�QD[�i��x��M/�ē�?�������F�Wr}�o��j�];�H3��1:w��O����O����8�D@�L�5Ną�ꊒ� Պ�U������`�	ly��'�Bč���I�Jf��6'�  �ˋT�{�O ��OH�D�<��K�T��O��+�`Tv��*Ǉ]&v���g����O@��?A��R����ć�l�X�I�
\�V ��cM�O>�6�'|�Z����k]�ħ�?y��d�F��EH5����! 05�t�$�xS��:�F<����&:� T�ىa�ܢq�ה�MS*Oܝj��ͦ�i��`�D�(��'S�Ea��
(U8������4�?I�mr�D���S�'��}�2��r"�bul� ��nZ�=�|�!۴�?��?��'Cg�'���/)���V%G	l��z�G��E#6MH�N���d�<	1�ɟH��)�!?��A�m��N��p*EƟ)�M���?������Ҕxr�'Q��O U"�H��`{��3�	�hp���i��'_��S���i�O����OJ9b�Y�>��E��.,юH8�ϕ��1��) 0���M<I��?aM>�1i���U�DT��2���)�'?�(��y��'jB�'��I�!}:qQ ��c+ȸ�s�K�AE��k����'�R�|B�'�� �^��i��Զ:��DQq,�=CA�uP��'>R�'��'��\>m�@gQ*�M��~���� ):QPe�vʔph��'���'��'���'t6�3�O��BH�5Ĕ��j��?��`	AZ���	ԟ|�	Hyr��s�D���G	'<=��*D�H�5��%#������	Zy"�'O��'5��Zd�'��iݩQa��<<X!R \}<�ep�,�D�O��Нpe��t�'6�d�T��r�pR�ؚ�s���rk�O��d�OH%�F�Z��ȗ�'!l�&6��d�g��M�-O��SӇ����Q�� �����Q�'��5��ƅL�୓rD)�4�?��k�Uy����S�'>�j$ �Cڪ�0|�I�m+̙m��OfdP@ݴ�?q��?��'v��'�2#A;w��	2@�8�. K!�O�b6��u0��"|r�c�\����;,6�� �)�m����iN��'@b�N�zCFO����O��	&9#��@F��^�"A�q�~`7-�<��5A&�����D�OR�d�Ok�ԧ0���ۃ+�4EP��q���9��V�'g\�&g*��O�d,�����ҍ�Q�G�X�0h��ַ����:`!���!?9��R9I��pj���?����3);�=�"c���ƕb�L�9K�޼�&ETZ(<� ϑ02�� �#���avN	{�'����I	b�h"��a���k@�MM�ސk����G �`��0�m�<]`��@�qh8@�6��Y�n𪐂�5x&@���T��m�Fj�K�F�-TEmI���<w��,Y��*�5@��iG0��h��:�Z1�рߟ-%���C%d�� FI�d6vQ�J�_[�9�a��!h��L��?q��?�B4���Lg5
9��� 5�¥�$��@a$�v`��J�����ŗs��Gy2�&t�\hf�:z��Ҡ�Kvz!
D��:��� �.V�/�r)Aք��i���Gy��ؼ�?�����O�T1����i�!�@��&���3�':�r�Ԇv��T0d�S�l8��L��0>ё�x�d����ԙ��[fe��yR�ԡEn@6M�O��D�|b����?����?���	�?z�P��0w�B�)`n�0g�Bг�g
B�n(Z����5�&�D�y�Y����3�
�z"�Z�Zh���U�E���9SI�1r5�Ãʆ+g����L۱�P��߱�/ɾ00��t�޶E�ࠣ�)
��l�	ş���'��I	��Zu�>g2�U����vԄ�	��h����I��M�ӫR1è�Dx2�'��|���lQ�㠎�t��f�#�"�j���?��	L���`���?���?�f���D�OF�2�)�w^��$�#Y�`��1c��y�@�	H��8��ܭ>��iC��{�O2�I�Z�t�9梐�#e\!��`렼����y/ m	B	�x�u(�?]
��&1OԜc�L	/�8m
Į��'��}Xa�OFtY��'���zy"#G�&kr��mP�Aѱ ��yB��K
*m���F7S��u2���g��"=ͧ�?+Oʡ�VIȦ����Y|��4�W,ئ)�&�!4��͟h��ߟ,�I�t�`���ҟx̧���0
R�_�	�d��z�Q#�f�?ye�������� iN#Q�H[�IA}�'��RCi�!&����TUCZ�H�%��M��5�H�(}+��F我o=N-{���x�'�|����?��F��Jn �.���x�ʈ�hOD�?q5$ͻP�$���� �-F�Ih�b�<gI�25��P�ٛ:�H�1�S�<�d�i�V��1q�֣�MC��?y/�lE·B�aN�{�JF��k�IA9Q/�=N��O��f�M�fI ������`A3���a��0j���.��ؙG!Z�C��հEQ x�Q���.�)���8�V�C�VA�T�O��=����*e�@`bl�G�b0�פ_9iQ�(��&�O�ID�$	'�z���Q8�Xuib���yRKko&��器b�a"��[����*��|z0�x�Q5xt��t_�S�!kQN�4�y�L)F)�7��Oj�d�|Z���(�?y��?� ���ƹ+6���hX8|�6�)�!��;���ÁF��Q�L5��-ـh��/�#`4c>��]	yt�Yg�I�WoB2�J-
ډ����B(��1��i��Ӧ�Nl����w�Ƥ��C,x}v�j6�Iy֒=�ǈL�P��B7���O����]����p�G�S����"OQ{�	�rI���W�ޏQ�bi��$�O��Dz�O���
��qa�-&1`x��bؗv���'\$q��H/r�'�2�'+b�ɟ��n�r��H֬/���`Ҋ��I�rޮ��ǫ<U�3(
�:��-�qH�3y��DJ�w5�}2LȐ1���!�f���9s�$�~�dħ�?y��'�P��/Q.\������
�'S�L��@$0��h�V&_.&40�!�j4�S�O��}jӤk�x꓆�!�V��wƃ8�U�'$�O��$�O�D9PF
���O�� W{�Ķ�����KK��HfC�.6FpD!�C��� �䣃�SW�L��I$6G��Y��=�Q�F	'
}1PO:z��Xr�\<[�" l�)itXh��"�(�	8�M��+@�_�� �A��4S�x�c�q��&�d�d��y� ������*.[ڔ����=�0<Y���L2����v�Np�1kI&D?�$�I}�T��8,D��M����?+���F#�J@L�0�鏎5
صzWI
E0����O>���:@�l�)ge\�|%�4A�Ώ�5!D�D�r^ZD3Ѫ�K`�]����
~���Iv�DK���}2����ʦ}����Ц �=T��Q��jN���hw��Y�'�b�1�G��>y1&�P�K=�e�G�"�Fl��+D�8F"�!:`]�c̙
s6�m�+?���4��e$�x+�G�/rth2�/�к	k� j����n���M���?�/�L�U��O����On$���O�ܹ�!ɐ��vH ℳ�@��=�|Fx�@/>&��I��M�>"ypf
�M� �)���8Q��V�R�I�mzCv�"D�Q*p����S��?1���*D��s%����`�rU��v�<ن��9���'�.n���QG�G�'�#=�O�.�2��?%d����=xĲ� �'��n��'�6��W�'���'���}�9�i޹ �]�Q�X�5'uy8�ڂ��b+0�H 厁ksB��� O�X��������Nk���䆏i�`�� ��g�줹�N�<CN\��ołcn(�x�ݟH\1��ɘ'��xI�N�d蒱�C�8/4-��'w�$c�e�a{�+	C��m��o�C�Pm²���x��';��;��T!;H�b����#s��HE�&��|�M>�A��ʛ6�$1>���U/|�HL���?Cbr�'��'�ę��'m�7����UK\2rHh�;�e�&)�L%�%�&D����k͕==�i��hب'X�K�h���(O���m�
J��iΚ[��S�"XjH<[3�-�����O�����F���(OF�*p�'��6�6���˄������v��|T!��ܜ=���c�ύ�֕����3Gaxr�����b�næS��D�ƌ�9JP扑�M�L>�R,�.���П̗O��Y#Dղt�u*s��&�z�����7N��'�Rʝ��&y�ٺ\d8�c�/#ӰM��� �Xm��� ��"EN�&��9���D�
�݊Vg (7�L����b�``�@+Z��UA��N�'�И� )D�I��I�<Q����Ol�?ѫꀁb��E������A0�i�L��vx�0$�$Sɺ9��s�c��%?A��4��'��耆�9y�P��'ޮU��ɑ��d�h��m���M���?�)��ASQ�O0�d�O�9;��]<T�<�%��v��0�t�_"T�ţB%e�zXh7�G�~��J��':�b>���;�L��d��e�B!��O�zJ��H�u66�X����?�>D�Taɐ��т���wQ 4â��'���r*2{D@(	�B2,�;���O���Er;h!J�C���p��"O@s���n�5���/9��DY��D�O*�Fz�O"A��_S��[U�[�;#v:��1_BR�'h�Rș�a1��'3b�'9tםΟ�]#&�@���v�h(1��?ZZi��-ųj��a�����вi����!�4!�y��1W&N��q�ʨ!�EYd��l8�2&�A���
rE�JH	�O`�Ld����|�o]�D��2s�"dR�.�6�ʹi+������O����:2�~���!\'�= �g�� �B�	���hp�D��8ño۵^5�I�G�^5�HO�	"����U�`0l;-�(���^�IRE0S���/V����՟�I�����@���h��؟@��I&',0j�4|)D�C��4j<����<z^LL{ܴd��X)%*�,GŮ(��D�u�X<��jM_C��)Roۗ���r�̓�t�n���ٗ�X}�2�60�<�s�lX�YC^�O8�s��''2jW�z�f����*�`t%�8' B7��O���?�)O��?��%`��j�����n��I�n)O@�=���^x����ڎb."�"��I?	ݴ�&T����
�M���?�*����"�ȩ#
�]���6>�.��G`[�F��$�O���(Jh~%����4*h��Q�O�3� ���G.ߖ@���1�d�2�%��3)&l�c��r�N ��bҡ$�D%�ԢI���i�DSZ[`���œV��5� 割0����S�O����(Z�1I&���Bj��
�'���цF!x��HjЂ�s�ʬ��iS�'d&YR��qk��V�h-v���'�8�yӼ���O�ʧk��i����?!�7�2����K5-�Q�,,��S�N��f�T")��|����X�
�gT�n�E)��LD��%M�)p����� �c��H�A a��}���z��߁�f�d4�s�R#����E	�k��������S��?B�E"A�:��S&�6?�>9���U�<���J�!�9J�N0>5*��`�E�'^�#=ͧ�?��D��ntd����7�-��?���Aڬb�J�3�?����?����.�O�n�0ܔHY� ��(�N[Ή�p�m��jEre�Ɂ�J��B��՟*"=Y0L���жC�<9���b�����qa�_;�h��,��@�*��'�HO���L������98�V�Ca�O�4�W�'-���$ƟR7��0ŧ��P��1;1�٦�!��@;(�b����A�S�ܡi�a�2 �IDz�O��'E�p`��}ӶM�iҞ?��x� �v`rG�OL��O2��;Zt����O@��1zƱ�F�W�>�T`��gw��2U��>` �EC'��;[V��t��s�'�^�A��8�4<UH�T�hH�7��P�(f�H��gi�t�џ\@s��O��o�;T��V�E�bV�`矶o�B���X	�Ǖ?e�*9�杸%�B�0r��	��)C�w<� �@��l��I��ML>��Ȑ���&�'�V>��a�JXT��H�#��p����,Bn]����ɄN#��j!�^�qX�PSgL4� ������R%ӑLq��ypL��XT��z��	�sN9�s��L%D1sNN�a `l�O���!��X,�n��&��"�*����B���'���'��:`(<2��0Q����+r����Id�S��yl̆�p<{���Pmଡ!S�0>���xbNL�h��`�8P� L��˦�y2�˅/�6��OD�ĸ|�� )�?a��?Aj٣<�\D����H"�փ�6|�H����O?nK�oR����\?��|���U8�*Ǡ߹C�Ԉ�EF؛)��`w��ra0��k��id\9����eQȣ|�]0U�P�kB�"Z����C�*��9�ğ$!J>E���5�"����/n��qХ�� ^�v(��m��Tx�B�13J�Rg��>��HFxR�+��|���V`t�EHL+l�%Q�� K'H�Q���?��� U����?���?���8�4�ࡲ�
9��5c��5{>:H�����n���J�'��Ȳ�FN9��iH�f���p�y�2 ��UZ�i@�b� ��b0��#��>�ԈY�IM+��i)�O���7�Ay̓��h�<e����^��6��9�	���=A/�9�t	#	�{*9XE�IE�<���>`�^I ���OB��ā�W����Sp��s�~(Q�4GD� zU
 �>��Q(= �x���?����?A�DK
�?������n\3�MK�NDn����!�	Z9�8���Xv��\����F��%%��@j ��sJ���8T���z�A�F�Xy8QƑS&�e颬8��Oqc��'"L7��:�0QQ�[6,t���j,!�d�x�t3�K�v%x� ��"!�D����pG��/MDڀ)"jGl7���}%�t�pkY�����O>ʧb����/�NDh1O�"ZHX�T���?����?���	{�v=��<;���i�;,>�Ә}a̬��)͖)@2)���M�*�ԣ<1p�K������!re�A�����9U��`n�8�( ��)�Q�����O��lڤ��O%��aR�F����g�!)�,�ў'pB�'�.��!�Q
u��P���X��%3�'�p�q���{��1�T&�ꭺ�y�'��yB���_5�5$�7OzL��Q�C �y���70��1���8B	�2����yb�ޗJ��e��5��ٺ��J��yB)T2^�!�N�?)�.�㗋ӗ�y�O�E�,Pw㛖��hr�È�y�K�~��QC�,�;sJP�  ]��yb̪�N��q�ܑ;�b���ybDX�>�6�@�NA/^Xq��b;�yC@���	���	&iR�R'�н�y¯���ٙ% � ��u*��C��y� �z���Y�"�+0C�U�F/��y�
� �|x����*���Bǌ���ybo��p�*�8"�H%����>�y
� ʡh�4,�y�0mݚ(��@�4"O���ѥU�E>r�ۄk�!2�>`""Obx;���4�H�M����4"O���Ec_�Ey��̉1�ȵ�"OB�A��JHVT����i��4آ"O���A$N�"�´j�KD�p��e"Olŀ^�F�q���Jے�Q"O���h%aND�����1\""x�3"O�h+�#؟�(��E�+E/N��"O���W׹bo�e �ER80���"Ob�1��`o�+_.�����"Oz��Em�W�0���cڜ8�(�"O\l����/�fb���+�lʡ"O�h���Q��,��_,s��Hqa"O��� ��;�� �� ��u}���"OLy��茋{�>�p&�Q�uZ���"O�abU�@?e��u �J�-/epyRQ"ORU{�Ըb���9��*I��"Of�C*��:ڴ�0���G:�zj�@&�Sy"�.x}6��5�(�K���i�E"�c�q�08�FB�2ݛ���O�#S�c�$�c�%#LO�u�40�@ix��&zƄ��;'�jh���'.�a�cD�a�g��a�<	��3(�<���Zq@���@����<	��B6�`��F���?����r��t�$�N�)�� cD\n�I�i� �=W�'���&&Ǐ]u��פ��,T���p�ǁvp���;�ɱp��� �(�*��IO�|
e�9zM���Ӭ�G��8��K�'�h���
��zQ���S��h��9@��Q&2p<CA�,�d��usX�
V`^�&%��Jօ�_3��[1��� �f�L�$XX�7g��5�X�R`N�f��'sT�s�i��~�\�W�̳ �5���i�<��G�+y*�{�T_8�8��DL�J�$}"�n��jx}"E���UDD��L�56�6x������v&6y��|�d{mṕ'&��l9����x2��T ���c,^4@�=�	2}��a��"�*|� ���"%F��O ���)�	��?���2cސ�����%��hт�:��+�fՉ'��;�%N k:tC��������'1�xbR��L%�ٹ�� H�昺��`��D����V�޽f((
aPtG�'Ԟ���'K^�V���,�9(Q�c��@k�2��S�'N���G T����/[8V��J>�雍AeV�Z���,"$�s�E6�M�5�ܪK0�3�M��:�����ΰ*�t� ��=p��q���l�+�ݼ�k���f7$�B�|��G���I��B֭N��jq�ےL����w��x�݉�� qC�OV���M�I��Q@�=b�2]0d%}2��0��'q�H�W [u"Rn�ā��LP�fN�xKe��&4t�&����w�������p��I
kx\5���b@��؂!2��5��+WN(��'�\��L�d�0Y��٘��%��X_G��� ��(r"�Xu�A�_n��s�R�mj�	�=i���~>�U�	J=f��E�Ok���$��E!Q��4$�n�8���N�h�JՐ�͍a����i����ȶ.{�	��yu3�͡l���P����S�!�����'.���'�O4=��5zr�пK�#��'Q�q���9#?�h#���|p�@���B�ܵʀ��9�"T�#<\O2ᠱO��HU��
鋾��8P��E�8 ���n��52M<qJ:i]� hbf�6G*�؃�@a}�H����)><X1�B��y��:����q�qOtSAAgA��?^,��q%Eê|`�'�4e��F�e��4�g�ȧG1�`�FC6
�`�Y�Y3:���,Gx��#~��%	f�'f����+�>�x=��O�P�}`���|=�xZcڈ[�cT �T����M�6��`�H>�����#n���تn.�Qb-I !����DG$"+r��pO��d��	�
�(D�(�1���hjԄ�vk^C��!�?i�{�N]�(7�10�C(D�+�$-��LV�%�Hy�f_v≌�X�����,�`3d���e5����NL�a�V�S��Q1g��A��Jܓ6��"�f4����J�2t�8%�|c�jtM�K�]%2����Va@\�rIǤ(1�Ӊ{��	����X�B�+�-ݪ|o\�4=P�dcu �B]Ҭ���_p^�I�I(	
�0�H�h<�Oܣ=�}��G�h@�p;��U>���$���0=i�"*%PA�`P��|{FͭP0�D�5G��΀�@�-��`�1O`��h���s��8ue6 �R.Έi�~��(� �\�ӎ􄏖r�qG���@\�4�2����(��B�� 

��!Gc���R��O�G��OZa����*����� hP�:OJѫ��<�)�	� 
�Z���m�,���"H�AE�y���30`�ʶϐoLPl��7��<��I�E�8�B� �蚑SI�g8�'��4!�O8�Z��C$k A�'U=sr�O�qqi�K�1ƃ@4��X`�14�� �h
��h��U��(� ��u�i� X��� <*y[��?Nu�(Oq�k֬?�`XS�K�4��0�K� !�]�'���GC�
C�ȫ�K�#7��d{�i_y"��q���OzhIBSi�s�	�i����$G��&1�1��K�>�����[�~;����̣d�tz�F^;�tR1	ְ{n�<HE.X����XU`��Ɉ�\�!�l��le�0n¬Ғ#>�*�qD�lz�	����L��HJ�<A�ńwj�q{f��|T���B$���x�&��3J��%�9gQX\��N�牲0G�e�p�I4VWިK�L�$���)�S>+�*8�R�����цܲf�C��	��v
�O���*�c�n���2���/'`)��ǊK?���>)eIZ#�d��dZ�B �[��S�<�(?l���â��'OMr�c �Ŧ���	�8ؔ���Y�p��y��[�[/�(hK��p_D���D����=�曨xZ�	P�蟗7��s���5Z���u�� ���b)4�dY��:.�)��D�Y���rk.�	��n�˶�]�\5����O�)�Ec1�I&U\�h�aO!�y��^�	Z��C!U�v@ r�J���D��L�
� �{����W�������k!%�[�!�$
.sn\�B���~��ٗΆ�#��'}�$з'�mx��F`p ���� �Z�°S��?�O��Y%��<P�]��Ő�Z簁���$v��	�'�X#b>�la�O]3f�z���
1�0������+^8��bI,�"��\/�y�,M��\���)+z@I2Ζ���GHXˌ{��Ϳ+��,�$��
Dz8�fɊ{�!��Q�5'�l@�GW�([��J�rj�6!� yp흒ea���䓀���A�/Df %2C�XYa{����Hi$��A��쓥@8H���Ggs� �l�xh<a�(�B$v�#�߱�\�NQj�aW�Q��E�\T
��%?�ӎO2@� RF�~1Є��)��B�I)`�B��!�f6u�dV{��� R$/��c�iCG?���>q4���u�QA��E%?�68�PPOx�8�T@/�ihY_���P����|�&MФj�XZmrp�_)%���f�$*���d�0��9�
N�XNK̕�t�������98
��b�D
x�b8/T�%B�[����%i��+��	
��C,�{h<�f��f�x�LȬ+���i�́�aq�)�,\��qmF0xm�8��Ů<�}�1T`�xE�0PI�7T>I��c�rDȂ#Q�N�rXK�=VZ0�$W�l��I8\wPYkUX?%��AA.+I�'7�A���%���7Ā(hv������j��(�p��
������H^u.yXV��x͠��UBȿo�e�Q�"<OV�S�$�e�쁑dO�g���b��	�t+�(hÕ�4v�����8�|�I�hԠ�cQ�!9s���R�]��ȓV"��Q%ʋ:d��T*&�jy�ɫ\բ��G�@ }N�`ơ������*�f@�C�1_�
�+)w"�ȓZ���E����0(�$��������d:(%��;��Y����s��� @�[uH�$+\O6	�F=�H�f�2��" H�m�>��/G [+�
B�����0>��B_!m�(z�ǚ%b1����T̓e�b0�ġ�4h���B�gjp����!%. � ���3�>dys�֢�y�N�/_#�P{��T�#j<��w��ai���1��G|Hd9��/����L'|C���O���C�C �{��P+4!�DD�Ir�h)B��0l�PŲҍE��	�!XV��a'�[2��3A�6mň"<1��>�
X�֊R�M��� #_]��LiA��>X� �����w��F����!`�j蔥�N	�t�)Q ]�����Cf��"Wn_�p �Uh� � �1O�Tj��@|(�3`�Y2e�t	���S�6�8�m��/?�]H�j��8ؼC�I��)��O�Fl���%�^I�u�4���.���k�Ή���SܧV>��;^h���u�L�C��A�U�C:E���ȓ2�4�� �-R��q��V�05�'l�vG����胡I��u���F+Y��BX�Q�:iHR�V�<�џ�ӎ+!�F,� )X'U�9��B� ]Ғ�A���%�d�`�̀4���!%�;tn0�[&�'44���� �ȑ䗿
[$\J*Oe:0+W�~*m��!/Iq��!���T>���! 5J� +��4X`�=�'D�d2d
�;}����B�:-�p���LW.������1.d�ѮO��?����&:�� ��B*�SW���0"�+��\{@�'���F�U~P�u���$��̠����mM�9C�����b�"_�'��=б��9G.��L�rat����D�.{g�0�R�ؤ��.��?Is�%%jj��@vH@=8��]q�h$D��#r�	G2.�a1�å8��}q�+"?��jB��(���G�=�N�!��tl��S� I�*
F1����!�d��-���*�O��`����ʚ�?�&h�F�Y�b{4��	�?+�(����|��:S>X���nC7L��I���K?�y���L�q�B�U좵YVM�yiz����T='q,eZ�&J{���`�A�>�c#4h����$-<LOt̳�
�<@�`�Ɣ��r� �o38��w�Q9�~I��E.D��!�b��$�֐G���@0'n9��/_��A2#f	:��"~t��iX��jf	%(LtІa�l�<'���l�y�V�A�S���12�I��.*��[�(�� �d�f�I�vs��{$�Y3�xC�	�*h�ZV�^>7P0�a��&U]ZC��	U��IP��_�84�w���RC�I<�-4b��Z�2|���M�!��C�	2Nt��{S�΃�@�#�f9�C�I'~��F��0Q��W3;��C�I;t	\��7A�p�6P���;F�C�I�v��,P��U?cn�����V�LC��*2T��i��;�NhٳFى�.C�IC:a�c%ێ9�(A�;}�C�I�i� }���4�Ʊ�ǭU�]XC䉲d��{Iͩs�Δg*��B䉤R���H��ې)�r��fM>*�C�I,u(���D˲j�Fls�J�T�jC䉠t�>(H" ܟcGX��e�۶q�*B�	�G�A�ŭ�)pP�2 lY�^B�	�uF��'o� G[(4�ְl"�C�Kɂ�J1�Ǆ�ɐ���ffC�I-y���1M�3�J�HSP�2C�U �i� f�.O���w, �^C�5�i	�k��a���s��%0�B�I���B&��@��cRB�B䉃 �2�9�˒�+;�5#SG�K��B�	�pn ���� �l�p��z��C�ɸ%0�m�����ȁ>��C䉲I�|�	ɭq�|�� �ޜH*�C�I�� ���q�B\��ɝ]�.B�ɣ(����"!^�P��E�5��"zB�	�)��e�1��ǀ�H�Hڼ�$C���ij�ͩh���6� �C�I� �#��-;<Fl��tڴC�ɮK�h��r�9XBp� ��E��B�0w`���f�y�:hj0$֐Y��C�	C{D��ZC+
T���k��C��}(�	�'N>AI�AD�ҧ:Y�C�I�$����cHV�5��|�P�G�lB�ɨk��xbbQ�pL:��B?�vC�	J-�M#DC?-�Vx�@lB�Q@~B�	�HGbm:ԏ��$�X�c�i�tB�	�#�|x�D�4:�1���DmpB�	�+���s�R�����֟92rC䉦*�>���� �L�@��֗TbC䉠Q�\���A�y��j�c�p[�C�I�H�tّ�S2�������P��C�I�Rfey�*U-s�eA��޻hޤC�I�~�9%���k��aQ�$�Z�C䉳D|�*�ۿi���9%��<_9�C��Y؈9�����@�AC1D8FC�ɞI��P�E(b�p�� K<C�I�G�X�� �� �����DݧC�TC�)� s&�ء�H�1%@�8�L\Q3"O]j���8] Ψb�)�3	��PY�"OzѰP�U���<��gέ_���J�"OL�pH�6oѢ8
V�	}�X�a�"OP)(�-�&`��q�Ɗ�N��l�a"O�lɣb�?Uڽ���P�$�|(jS"Oz�k&��O0tŋeE���$R"OBX��@��Cq���.����`"Od���K��H�΅��OK#0�d�C"O:x�"�:Ş�iW�ŸO��[�"O
���_�>����&J� �"O��a�=Ta|��vH�-$>����"O0sN[�y���B t$|�"O�p@uひL��X�0f�"u2,� "O��H�C���B�9�\�Td�HP"O�+,�4j��rĤOc��q�"Ot���΁��(}p��<5�(�a�"O��Bt!�	���2�G�0��8J�"O�*���\���\�C��ݣ�"OX5X�J&i2ݢ�D4S��YQ"O�,� o��L�*l��G�p�LS�"O����'Y�i��Xb��D�!w��7"OH��c��p�<�q�� *[\D=�G"OBI�E��f*���6iW4R���B"Od�W��LR�̩caڸV�*���P����I7y��ɵ�PH@VF�6:v@�B�B�	� B�ILqBC�Z�K,�Z����%� "?ً����9(�4h���-Ij� �7�!�$)�h�ڇC�a�����<bG!�Uy�̍�"�4b�<!�Ѯ��,9!�d�+$ ���L�)����v��=w��	�n�}��1e�`���N��VBP��yR�"wCp|�"��A6���)ߴ�y�E
�O������4ϼ�p��y�E�2J*�����+�R��W���y�]$f�H-��C��e��䉰�Y�y2KQ�T��glݧ]3����F��yr�B��m�慍�N�T�+��
�y"�ޥ1��\�`�˗A��1�FJG+�y2cƻg��|k�?�(�0Sa�1�y2���B�w�\3����C�/�yb%č|P0L^"?p�����y2�¦R��m�烉+Y���pě���0�S�O~n�S����O ܠ�!]�i����'8�P�Ȳ<�~��A@ڷJ�pH�'#��	�M�<��֣W�m>���}�)�i�8W��]�0�M;r��t���!�$_!`�Q�C �������K�5��Iu�ۨ�RL�7E�'+3n��t[J�"�"O�@(b.Z#}wJ`�V�ګҤ�8��7LO@l���,T��A�NT�1��
O`6Mײ 6l�!��q�tP���+S�!���&�����i��B�4,IG�[�l�!�ď�j���Ë�-�z��'b�3#���dŁR� �3U	�t�Y���M�'	����7*��A�ۋK?����';&Ӧh�*��a�FG�Zi����'���S�j
&Wx@��2�=N2ts�'zNȰ�'��}�jh��_5!&,�)$�\�G�� \�t���H�hf ;D�|SWkí �:��1��8n�8 �!>D�\jtc�?���3�3�n�h��!D�t�����z��e0[ozX�4e=D���ƽzx��f͓p�y���.�$4�S�g�? H�:T!#2��;Q/@�hmN���"OH����Xp	�˴c��ofԐ򵖟���Ʉ1%�L{'e�%5�H�����!q	�"?Y�'��I�����	�ٱ�A��:���u��B�	(s������Frd֧��X�B�I���3A�9:���i�eK�B�	��R ��螒K���Z�E(?���0?��ꝯ��X��X1g@h�W�<Ih�,�I��M�4������P�<���gne�$���F�>$��%K�<!���=�֡�Fo�܄� �y��7o��S�
پ�X��@��$�y��"z` %$\V-�&���yB��]�@Hq��ìOo��"�ʌ��ybK�O�"����ZuE��Ju��+�y�Ʉ�|���A�fܢl�s�#���y�jƠ�4�V�W;k�� ���)�yb�.n�mQd�_B.t¡����yR΀( ���̍�lP49a1��(�y�k{��A�#ךU��ܪ(��ybhD.OM����H�.�6��Jʬ�y�\E���Ӧ,�1c�����]��y�ǈ�-n� Pq��	 Ğ�x�AH��yb�<ea2#"�ٳ�f䣶�A�y�� �q�%���@V��kخ�y��\�Eƒ�-7T��t����yb��P����DhF'pZ}�$)ۖ�y�@�A�^=�V�^�,�p���^��yR�v�|;tE�)yI�
��y��/`���FA�4`�����y���E0��V���]�g&�:�y����c��1ą�t08M���I�y2_�o�zA)�M
l،",���yR��|��0a���hU�8#���y�>��(�6J�l�r�	�OK�y��~"��yÆπsEpq���y�n�7t�Zdpu�ƀo7��eX�y�&7q��1AGh��k5��Qqh��y2��4DR���2���5<n�`C�D��y2���i�$l�s�V9�R|@�e��y�-Y���YmY�f���F��Oޢ=�O ���6�D�8����V�[îi�'�f�I��D���b��^����'�l5�Ť�#N|�	C�(Tt����'t<��fRC��9����Md�}�E�(�S��?9f�y��g��>5�媖��g�<A1�6&H���3�K/y���IKb�<�e�݁7Hn0p��,}�^���`�<I�H�?-�%��"P�xL�S�H�<I� #4��4��c�o��r��n�<��o�CԀx:2H�&��M����j�<A�I����T����i�<��A�:��ys1'�?K�v�Tn�<qе4<��xB�8\���D��n�<1&�¿B���9�o�h1J(3��T�<1����_(|�d���G�W/UN?���S.)`���BļXtN�;�(C�	,>o䑈��%�t�y�,,l��B�%	�̝:nZ�~���.Q4��B�	�n(��CMO�t����<��C�	�o�tK ����L�봂�(��C�I�4�%��%R�]�^�c�	h�C䉿]���b/㐜�t,͖U%�C�NH�����
>X��S� "ʈC�)� VL���S�y�Pb_f��d��"OR|�5/Z�*��;� F�z���"O}���u̤�"�T.o�Z�A&"O�\xc�Cg���ef�#A䨘�!"O&�(s�Ӹt�(�a�Ϡg��}��"O,��Њ�=SK.H!"��t�i��"O�e���۹U,�o4�|y�"O8a!Չ�ro2���[�i �ex�"O�U�Š�B�P��
4n�J`*4"OLp�t�Ăe�X�QȚ�����"O� @�� �~��F\)���y�"O�i		\+dQ���O�$ ��)�"Om�a��J��p�to1$6��{B"O��&Y��L��,D.8�P�!"O2��M��TM�% ($	�m)�"O�-�g��n]�C C��_��QB"O�P@�U�d���H3B�2;�hB0"OA�rC�J��"���I����S�Є�	�zt��A-Ǧ:��u��X�;�jB�tG�5C��ǢU���'��<&�B�0NBp��F���p��`!Ӓ|š��@�e��+T�`f���$�!���t�J�gԴ��)S!�ҭ=2!�$��}.M2�f̑�z�����O!��
}1��N���t����7�!�d�.���Q���?�t12��<Z!��5gV�yf�X��%�5EF>f�!�$���H��n�3�`�;0!�$�
k{H��	/bFl���l޿4�!���18m���O#^�K�l�%�!�1:W|�@�k�2uP𱊳i�(s�!���fМ�� mm��֨��oj!�䖞v����f~0~h*��%6!��%U��+�`O��pX�f�V!�$�q�r�����03���s&�
�	7!��0��R�#L�r��!��ݧR!�D�L>�(���'d��I�Ϫ<�!�$޺K��D�V.�4$���Yj2?�!�$�>t#�`f*�l��E�/��+�!�I�6�Aæ�I:b��!sv�T�c�!��<4t2X8�˅�0�����A��!��V%|�($߂ ,����e���!�d�gbl��cB2$X�	Ş	P�!�d��(��-I�'�?9?<0 sC	 5�!�$J7C�L;GdR>W[���b�k�!��țP���#c�,Z�lB�M�_�!�D�>�`I�iI�T��s��GC�!�6��*����s:)�"�X�t�!�dy�@ �EŇ0��1���2�!�"j���d�O��<���)͸:�!��R
j���# ��8�0I!c�!��Ʃ"#�LAe�4<P�9 JL�ip!�$C4F��  S�EĬ%�W�F��!�_����&�X'Q&<"#�D?k��
<Ä��C�o��0����y��7搄@bǄ�1���+'� �yb�܀8'2|	Â8&��x���C��y����O���K��N� �ҵ dֆ�y�D�C�� 3ˇ+�HŠ5D���y��U9z�|EA��E�r���)�y2�V���PT�C,̀P9ÁT��ybh�z&)�%	���l�[��Շ�y�,�=ȡ���ܔ	���yBK=)�p��ԏ-j���2�W�y
� �����>���;��[��p"O"� c���G�n�@ D�"(0�4*"OXx��a�2�­3��W~"�c�"O�L�6��ģa�+j�fl�b"O�S�O� X��0P��.U��"O�t��ñY?8����.��5;"OΝ�V僉1��+�c��w��h%"OЅѠX�C��XzW�6-W��"O�t#�`�N�@���Mv��"O�uzь�N��  �AŁ^d��"O��� ��
|ں�a'��3�D��5"O�E��cݨE�Ng^%�"O��(b\���J���P^��""O��E�,v�a��&K^�p	W"O6�s�$o<��rs�
�fy�� "O���E�\f����(2u�5qr"Ol����� �\�hD��p²1��"OB���.V���)� �O�T��u�@"O YH�UIe��Fc
�\sn���"OZ�f��X�XD��@̱B�]z"O�}92lװu`2p����*քӖ"O*9��	-tB8K��)l�� ��"O���	 H��E��!T.zF�	��"O~�H �U�L��z1�E+(B)��"O�(�gL|3.M{3 ��~Ϝ�J�"O��r��¿mC�y���?��]�"OL��V�:9ThqҠmރO�(`xA"O^�-T8P�MN�(H���;|�!�d�s-�m1�BӺ+a~ H�jI�G�!��J��@��B	�A%���iƄd�!�Ĉ6.�։�fƒ�,�
��	k!�D���ܬ���~ڢ��ț8!�$��!��=	WŇ$1|�bWf׿�!�\����$/4��GD�=�!򄃎Y���S���-	��ZEܾL�!�$��tU:��7�*d*UO��y!�Ζ$"�Ȓ��R8 1�"OJ��q�ρ&<��El�`A �zB"Oz�)�fǩМ��w?S@��""O�i��'�����X���j���Zd"O@��R4� �V�;.����"O8��C
]^I�ӂV�9,���"OB�p��S=GL"Q��L��[��Q�"ON�����6H�(�+�
�l�3"O�lP�G��9��QZ�	�#,���aw"O�8���5E�q����'P��<��"O�A�5������j"��I��C�I�Z�� r�!�p�)գݵp�B�ɧ=8rܻ�O�=��)i�H�)bTC�	� V��p IUUb�u��,.�C��4#��7O$�̃7 @$B�I���M��ёB*~;�@À@��C�I���bVJG,U�&0*�c��\�C�I�2���(��0>�2��#8�C�	,k�`hc���.|0"�<2��C�������ʖ�F��m��4ԌC�I*v�rA����V�|+f��jqNC�	�8�"�qH2}r�������GwlB䉥j.~t�`Tj�����ٚ@p.B��M��i �hЬCm�\ZB�I�K��Lj1�$0����ӪT�\�B䉶;
P|�fư�d����y�$���4�z��\]�� ACT�s����ȓL?���d��8z�33�P�\����S�? �<3'�g��@#}lT�"O   �V/c��DL>0��Q�"O\��j���@ J5���j�j�"O�`EL� +p�&E	�!̺�h�"OZ�"EO
�B��C�
�����"On�'�JS��! �Y8J��"OJ�� l�#8�l2���>����"O���RLӲR�20`\j��&"O�����g�jAC�H��/�f	�"O�x���0/��x�M�-ô��a"O����$8\�C�&�n�� "O���-��N�8�ZԈ؀�T,�"O\�2��E�/�f�(3Ka��B�"O<=��Cن)|���g���^�1"O @�q��2@������"|����G"OjI�Y�2�D�S�H�/��%a�"O0
�`�+C�Ҵp�+�6�Pmz"OdMp.�&Nd�H�Uv��H�"Ol�p�(\�C�EB�l؁gY �+�"O,�D��Ym�d��D�	s2�H *O�,�Mҫ6�d�i��3�fY��'9r�W!T7D����tJA�u���	�'�0��$���C$5q��|�'6���%�WC �MһeX���'3�P��,>Hr�=JեK��$�';V=�BG�}��=��kB>Vc�I	�'�D�	�4���j��Q���		�'��=1�[&T�>!Y��@�Jb����'Q8�k�G6r=�q�7a��=�j,P�'���B�[p���P6FU�A^ԉ��'�Z���?����!��:�$D��'ɒɢ�h&!���(����h���'�A���,"�� '����(��'x�r��Ǯ#F�(Q��_)C���'^�a�SJ��S5I��8�,���'��d�үZ�
k5bA�Z��,K�'�^�Y&f�# ]�%+�.Y��5��'��*�L�B<�QpUJ�*A��-+�'�Hlʰ��VvP� ����E���'G=J�o�C� bwE�i�y�'�4C�D��
�	'��^��'�L���C�V��0�u@�'���a�&�7��H�DX�A��Y��'�V�!�(Қa
aA�:�.���'������"/z��C��ܴ}9��' "�;�c���H���nn�P�'Ŏx���A;o5��06��2�xK�'0H�� ښBv�5a@�����'�x��� ^^�R��6k�;Rvl��'~�t�b�K~^L`Е !�*�
�'�)�`N5�j-#0H+4A`
�'��}�#hC�p�.}�W,�)��<z	�'��D
��TLh��1�cҜ%�,M#	�'��лNB��p:�#�g$Hd
�'"���W��q$f��.�f��	�'�hx1�iL㊑�b�D>	�%!D���n�Z� �	3����ܵI`�<D��:�#S���A�l�R\B��$D�h�!��0)"r3n��4b�����=D��F@͆�r����ʛ#\����.D��gE	���KV�ܬ|�D�'�*D�!�i3
g�\��)� p�FX1�M=D�h��(ʵ:W ��㘨BRf�i4�9D��i�?8��I��'=�(\�Ci9D�� έ�S*ŬGP���DTm3@�b"O
�ᦅL0���"�b���2#"Or��6�;��\��`N�7պ5+V"Ol�P ��0��Dڮo�.!��"O�o/ղ[ev!�	
O���%"Ox���ʀ�k�̥�sF��X��*�"O�q�e%2[E�] ���'6��)#g"O�=E��{�q0�D	\	��Z�"O�����-�&�����T�^q�t"O�����G��x��,M�5<r���#D�T�QB�\�D�H6	�6"b]�!�<D����I��E4��j�ŎB���y�)%D�p�p^=z�^��r��9uW�,���!D�l��@��z�s�m�N�m�bO2D�h2q#�5UV��ee��rU��(�E1D�|s�H
,�m���S�Pƌ@��-D���!D�1��P#��%a*�+D��X� &&�8�Xub
�-����;D���J�@
��pD"���΍�%�?D�8�n[ K���xfe�.bHrL�@;D����ڋm���e�ʕ,T�9�l:D��j�C�*��)W�q�(�0%7D������숀L�#_���J1D��!t�C�d��̉�)� o_�t!�;D�l�bG�ZF�uYF*O�>c��E`.D�𰢇�z��|C���*YK��i�*D����
�-�|S�N��
�C��'D�l��A�&e|=(SD�*W��C�#D�r4"��E���J"WJ�u��@#D��th��6CJ����>&H��`�<D�0�QV��=�C��KE`l� -D���0��&"�$��kςx��-D�py�(H�3����ME�!�T��%&+D�h�VK x�.1�!H�<�<\(a`'D�\�Q�
  ��T�-��]~
\ʡ�%D���Ҭ`�:M�v̇��Y�8D�@�j �l�|,"� � \W��ӧ 1D��[�l߸U\J<+��P+J���P@f.D��
��%0Ȉ�� ��+Al��()D�d�rlS�.���F�\�BB��2B�	�li2}	����|qDC$S�C�ɴ?V4�Y�ȝ�]���y�@�B�C䉳sW�3�i��m��㵎ȔLDC�	�����L�]�2�AC��>z�|,I���>���kT��C�:%"�x f<oM�E���P1͘C��<*��
®]x��k1H�nCtC�ɈR�Y�5�
s��)^w�L��'��a� 8��I牂�p�:1I�'&�8���3Æ4��%2u��A��'`�� �l[�E�A�Uv8)�' v ;!EY
�<8Bv��7V״���' x�!Fė�F��p�&_:!��,J�'BT���댋��p�ꝛ��-q�'u� � L?� �@B��as�-s�'�bH_�N��Y+b�6KS��
�']���Ǧ|�����@�A��u
�'Ј�
R�B^��PG�$5��P�'���9Ah�]��u,�*1?�d!�'��+��ȟ7�v�A0n-J�X��'-�Є�P�K�0���܎,���y�'n�)U��6B\%J���.�й��'@n���<�`�Ip�	.Z�|��
�'����4	�*E���7+4e�~	��� �	IM� �F�Z7�M���"OBPh�k��&�Su�����"O(�	��O՜�9EM'���E"O\�rqL���7F�>N���ç"O�Ï�Hw$�c�Ń�7b��6"Oظ$�h��`�G9q6�"OxLy3+]�g7>�b"�I��
F"Oe�㄀>x�`�����R�jB"O��S I}�%��CX����"Od�(ԡկ7�h�Wg�8[���"OR4c��!>�D����M?��R�"O�(�HG��8�E��X;��u"O� �E�3&RI�U$B�{��|��"O��@�D�~�5y�CBG�D��'"O858�C��K8�p駫ӆ}��a�"O~`�F%�}�L��C�y��s�"O�	�b��q:��C�߽r�(�7"O���+�
D��<�&K�#�%Ȁ"Oȸjg�0	T� Ũ�({�8p�"O��A�"�А��JW�|y�"O5R�`Y;���iEL�F�ɉ�"O���&6Ŏ4QBKd�}(�"Ob�%�
Xd~$25AB*X�8s�"Oh�b�f�W��4P�N�B�!I�"O a@e���9R �ֽ	��iba"O$l�A���A�1rA�4}�@:%"O4�K]t61��@G5U�$,� "O�@ �JM���1$-�-��"Ov�A�<V�b=q�A�-XD-�R"O����;_.mے`��+fȃ�"O�qBv)̾aDV4P�Z)��ˇ"Ov� ��gm(�J���	 "O� �@��q�ꑁ�]�I���O�<i�J��`��WC]�I�8)*�D�<IQ������S�+�2n����HB�<�5" ~�ĴCĪژ}9�U���j�<!JT�-����Q�K�*y�*�c�<1g�.~��K b <<�\�0�!�S�<	5ͅ�3tzX���:y�����N�<�R��>t�I����_b�\Q��H�<����Msм�b`�&>a�̱�)	B�<��CY/���k1�H�a6��°��A�<�`(J�	xB4a��ʡ&6
hZ�Yv�<�#�]�x��/�=�z�Fp�<�ED��L+�9��I�V�y�j�n�<�7�Ԕh���&"[f@1��#O�<2�ǯ%�D�@%��n�V� f�p�<��.�t!�񱠎A'���!�l�<5+A�M���!���P�����i�<Q1��R��q ��!��(�, k�<��Z����M��u�]�� ]h�<yFŃ!*�`S#V�#X��`��m�<�f��:�4H�0sH �i�/�o�<��n�8�<��+����!�K�n�<��dBA%RĠ���(`X��!1 �l�<��τ��:�IÆ�c,<�v�[e�<��t2�@f�Ͼ�b�@�{�<C쇔}��]	e�O�F1�Bra�v�<�e�r_�#׃��x��t�<Y�.N&#�-0�l� ;�:CGl�<y���?6��5�	�{����
C�<9%M	*���S�e#RM1���|�<�s�X�4$`�ZDV��J����^�<��F�F�n9��� xv\�T� W�<� r�HwC��(�ȣ`�R(@7��Q"O�c��:b�2��	�0A�"O�=�`*�<}�T	�}�8d¤"O�	�a?��xY�G̝��0R5"O�`�%�
0���� ���Hm�A�"O�@���2%�PmHS\:��"Op!A�kZ�����6~N@�ps"Oĩ��#p[P�CiǱIHd��"O���Ͻ;�2�Ƈ��88�"O��s���R����۸1"ONdK�-�+1b TC̲;�^�	�'T�+�oN�k�:܈PI�! Bݹ
�'�@xi����Vi�G� �pfz
�'�v!z�"2�V�BN62Tn��'�Ne�҃.H@�h)f��53�]��'� $������5iF�TwB�D��'V��p�ɿw��HXui�5@���'��0 ��"lOrG$�mw�i9�'%f��2�%����E��`��X�'�!��p�!�Ȍ�X}����'����ME��0+fn���Y��'y���F�S���BU.�h�Uj�'��"�Y�!���4s$)��'m��A�Ć0PH���Ƈ�x�`�'YJ��A��]0�@�V7��s�'���[�gK�n�I�n6A �0�'�"��e�H?��0�̲m&��C�'.�q���� y��Ͱ�Cm��݁�y�BՁZ �I"K|�.�k%�E��y2� �S����ׁ�o��4ɤ���yr��E�B`3r�ڈt�d	��4�y��?cXa��1f��U��Q��y�h�\.�%�G��a\P���O؝�yB P�KRܩ+#F�g�n��� ��Py�oZ�"��`��@�m������JN�<y���,\���e�E+[E�� !�L�<I�*ڜ;�,<BU斩a ��CDG�<�r��5f |�+�"�&9��Ih2��@�<�t�P��`A �G������f�<q�ѳ1gV��D�0i��pمN�w�<i��О7쉈P���-�ՙe��p�<q��Ⱦj-�l�Dj_.��ԣ�m�<�P��t�T�2��|��B4d�i�<	��B0u�093�)N5Bb� ڡL�<�L����5&�/St��RDQ]�<��^o%�`Ғ�Өvd��p�RZ�<1����<�`Pq@ɿS|�xAD��[�<���*kD鈵��:�ʱP!�\X�<�u��D2��G3b�^���P�<I�ƙ�k��FkDa�
�j��GP�<9cJ#Q��9c�@�/��DIh�e�<�5�R�~hͫ�b
�H�H�*TM�<)p���<�R�+r��'�Ι�G�s�<i�%!mc��BA�X����P��l�<��$�$����o2J���3��h�<a�(��|y �ё�A�]��Ҕ/�c�<y&d0A�Pzc�R1�8��T/\b�<��-�!Xhx8��*#�µ���R�<�g���B���䁎1+3�T�RON�<��
u��`*��~!�H���G�<�So
*u"��.Ⱥ,
��b�~�<	 ��D�X�f�^9w��)D�x�<� ���D�x�k�Ǝ�>��	u�<�I�E���ggؚ
a���'�E�<� ���ƈ��zG�Ś��,Dn@L�v"O�|�Ѥ�>Hi!��.#�2�"O������d�T�i�E�&���"O��86�Nn�^e(b��08��5"Ol�:���_F����!a����=2!�ă�;�(�a.H/1�i�lR�{!��32���1GE�?�PCƍ܏!��	+k�1` �K �Ha��f��$��)�'�z�F�{�恳&�\�\P	�'�6LIQ���l��TMR�U�� s	�'�����2����+��O����'�H�iW���bH 9'�R�e`�'�H�IF^Yh�,��[�@���' �0��(�?]{�(�AҰ�hy�'�u4��'$\iiw��	)b�X�'�!@�H�}!�c�oO�~�Y�'��-i3)�Y�|�#���
�'u����Ե{��(�5;�l�	�'ޔ��	�{H�S�A@�)�Ҹ:
?)�'�<+ j�6P��T`��Y��=����2O�偰�Ө�4,�k֔i lͨ�"O*��;%����O�:��"O2X��֗P���5fR�$��䢆"O6Y"�	_�[�QB��ǧ/�L �"O��0�c�לYY#�(�Da��"O"]S0����92�/|��x��"O64��#�S��ik�@��\�0��d�O(��)J)|¥��.�	���(�!�dK�gYv<{E��'���S�!�su!�dQ#h�F���w��YA@�P!�]0>r@4��탫�µ
�Q�BS!��&
<����ޯ Ȫk���
ME!�$�<E E�}�[%�2?�6$��'`輰��Es�P(���	nvDI�B�'#a��n_����c�J�:[�	E�̘�yrA�I���d-FC��i�diJ��y�≪LR DU	B�` ��	�y��y���{���%>vd!����y
_+u�8�PT��5NȆ�2!�y"nB& l$��B�֔����y�Xf�� :�ٍj)z05FU��yBŝx��	"�jP�f��	�\�y�)Q�v�`�ǜ*f1*��Q�^��y��V9o��y�$D�>5t*R�yrBO�/f��tFI�a� ��!Z-�y����rh�f��W~h��ș��y�c
#��k���lU�x�qBۊ�y� �"
&F$i�+�i��l����ybm�8���A)�/P!�-����'�$,��fĐKD�-ߏE1��'[�[��O1=� ����{�P���'��4���4,�(��EA#BhT:�'�p8���#*�����.W�Jh�X�'uzT D�ʕ����L�x��у�'|]"���Oeh�S��y�����'�L%��bÇfA�!"�GV3tFp��'��
�痔2��� ъ�
q=�̓�'>dy��=6ዃ�X<�#�'� ��+
��>�RVI.fҜd��'X���$-ْ}�v!�玱W�4(��'�Q��i�� �v�Q���;VǠx��'�fI#E�/q�z(�6�H�bm"�'�0�1�d�"�&Y1�*�!<l(S
�'9������7���P��M; ���
��� �����pR��cnJ�R'T�Q#"O�@���y>\�6�F�K�j(Hd"O}k�M	9?�pR5m��P2i�5"OJ�jBG�+T����j�k�q�C"O��;Q�
�z;����h�e���p"O�U+MN"%���z����.q�0"O�E9G�.4ȩ���D#�aF"O�Yh# d�H�s�!�E&�4��"ON�	��	j��QG��@23"Ox<3� �?u���[S&Z�h
L8��"Oe�P�� (4�xx�%�E���"O� �$Z#\����F�_�;ې	ء"O^�0�U�&��Y	�JL"���3"O�)���#���1�"�.c��؈"O����mI�Ca�H�C��=����@"O|�a��S��LA�A�"K�� �"ON�!�M� ���qà�~��"O>=�D&& a�m�\�"O�3�!L�D�2�V�U]��س"O������0U���Za��@�"O���厉�� �B/�	A�$H��"O:Ѱ���_��y�M� X���	6"O�ei�Z/���x�3D�Ph2w"O�Ub�	�9A� ]���A�Pr&"O�Es�BD��s��\ZU�8QG"O�y���7`�rDI�FY腳c\�xE{���� :"�[q�����<�U��8�!�DN��R�:�����$���� r�!��^��$�ݪۺܚUږf !�z�ҭ�]���Rr�G�S�!�D-I��H�0
����J��>�!��T(���������ÇkF�!�J��H�rϘ��ʼ#�i\	>��'�"�|����7}�D��%�ގbL��m��<)�C�	�ٮX
�� �fIh"A+�	K��C䉸P�d �D#E�e��8a�$E�C�I�:�4�S���u�s��� �JC䉪T!���jA�^f4� @P�(��B�I9Q�l�{�`K4co�,����-D�d0G��QN� ��/	�t��p�օ�<I��?�ӓ*!��ハZ~踄��bT���])H䋶� ,�V�!T������ȓ8�LL���]r��ivm�����Es:��u�m IARDH�Oe�<ѧ�վ3z�T��
2*]JԤ�D�<�7m�%vÂy�T���>����TB[B�<���w`PUQ�O��/g�<�!�x�IG���C�7[l���V- �"�aB	=D��GL�a���0���ڱ7D��p���2@�I\WM�݀�j9D����iRC����%�TQ1�n1D�����O>֜�
��2n�詈'�/D��Pd�5���g�Q<��EN)D�H��VV�&�S�	�P �⥫%D���7F
=:�H���ɖ���H#�$D��@ԦB�yI���T������ D�@��P<��Q2��4�N���"D�`�W��ɶ"	+�%A�l��� D�J�I�0#�:�  IL�m���Q3D��1��O��xvMK�x�
���.D�<��&�"���aRH�ޡR��-4� 2U#,h�h��U�2o�B��n�~�<� 8/�J����Mxi{�_r�<��/�5>��y�A���<s���R�<� 쉰`@1�.�:0�#U����"O��ŉ��A�����B׿j�  "OPL���yn�J%�3X�,=��"OdP2�H[zS�}0��V�����"O �k���(�)���¸ߺ�p"O,dS��ʍ^K���q�W�ֶ囗"O`5���A�#�*���nɫ&���p"OD<{�M"#��%p�,B�VŪI	$"OP��A,\5ΪY�k��y��`A"OUq�Ó>ZF	a�	:S(J\��"Ot}J!fD2tN6����r��ӆ"O���OC�E�(��hϖ<���	W"O� A�/�1v֜r�� 5d1"O,�CUE�X?b��pg�*n4՘�"O�̐��א?
 ���e�"��قr"O���n>��d*����o���5"O���f=U�f1��k��t��"O��S�E��VT��A h�d��"O.��p�U0��,إ!U���P�"O��Bo�}�T�"�y��	�"OJ-P�.8x|D�5`�(���"O(=raS�P�������i�:A)w"OT�`U-�^�s�͛X�I�"O*�Tv��E��R(h;�'��@�"��(��_���a���йH!����5��_�2��a�+C�5!�$��~��l�Uaޜ;����� ��~ !��V*S3(�t���j�a�h!��-mn��B �B�Wͤ�qc�H�D�!�y��Q��i��aGiI&!�Ă�o۲9Z^�r� )�ņ*��}��'���
"n<} CH,�f6gU�NhC�	�a�2�S��:dV12pCR�o(�C�I�L�h!B7�ֈo�!��N6"��B�I�i�ļ��B&_m&YD���:��B�	:"jN�3�HN�܈�b
'1�C��C]�X!�c
�����K�{`C�	 J����m�|�VQ�m@�w�HC�	�+L�A�O�U12-[GH
�8B�ɮ`�^�r���B��*�H�._�C䉕�(�S`hڛm��(��,�&�B䉱lr2	 ��M�H���r�݉mHFB�	"�p�G�O��]���Z zB䉑P
J�*T�	��V�0�b�($"O�A�J'A�Zy��IEP��0�%"O@ +T�ް`��D�g���g���"Oܔ���9�\���а/X%�"OT]˅�_gdj�)�#ݶtKt��6"O`�g�P
ʥ�VbW�"O􅑧��i�ް��&NfޱQ"Oxeb`N�#t~qS!G	@]Ta�T"OhY;�,V�N��p�OG��"O��֩�$�P�b�	-h7����"O�dD`�5",�h@Ů��N;��%"O� 2���ܥㆧWsYv���"OP-�#�L܎���JQ���b"O�$ p�6l���e��4�6��C"O�EbP*�J��X��� ׊�b�MQ�<YA��>G�nhphJ�}�4!R�J�<�͑�Ox�y�!¼A��Q�F�<��� gZ���C�Y� � 2ƚV�<�� �"��}A����Xp��V�<!�#f��EY��،%v���)�]�<1v䖀#�J,�G���B	�i;w"�B�<� ���Ph��E;j�y�A�%V��\k�"O�i�%ءL����R8fb�q�A"O�T���s�l���S\yE�'Y�ɦe�fi�A��YM,]�0FH��C�	��ƤW�٢R�F�[�X�z~�C䉼b�|X����&4�f�1ŗ�8=�C䉘b�Y�̐�I(��Q%&�`C�I.�d���,k0(�jϸs���&�n�s4g	�	����2 �3�!��@@tLhdd�t��IeȈ5��HyR�)�T 3{CrM!����L���"�y�+is��
b����L\�r�S��y� �>r�p�+6�U".t���'��yЬE ZDj�J�|�ر���
�y��#/�$5��O3E��`����y!ܓm�p���Y,+�BeJ���xӕd}	�D�*I8jx�G�J>Nr��$O�	sHču��8S�ˁ*���"Odd�R��!�Rp�Q��/Iv����"O��qb�U�H����)S_��"O��S�_0J��I@��L7���"OZ��P!�(W���#&?|18La�"O�=��ԇ����D׏O�H���'��K%Ԉz���/?X�sF���ўd��	?6�>	�5fÍdz<	4	�&'��B�I1tU�ǂ	$u�Rv�9�B�p�֐hg SqGN,���V�/�B�I?���努#� [�U�[��C�	;5`���Dj��;� ���O.]�C䉱�$X�E*N���]����:f�C�	*�b����\�l�vu#�P�**��D;�	m��~�.
�+�P�p&I!UD��c3�׏�?i�'�,�� I��O�n<�
J�3�����'Hti(V��K!:�i��F�a�'{$���l=a�T	a	WMP��'[:���i!���S�
E�=�����'	:tb!�W�%*�h�S��+K��b�'��%�v%V&4�,�B��Y����2O"EW��7@���؋Qǒ�q�W����N��X��V@ni#�b Vv�72D���
�k��4�N��'�ݛ��1D��pe$f�p�f�B����r�.D��&K+2BDm$A�y����-D�����M&*O<](��*ppy�u�)D�����Ј�E �ޅT�<���(D�4p�٫�|H��Y�� 1:ԡ$��2�O���pA
1H�����΅l_���"O�P��3Mؘ�Wj�0@_B�+�"O&A���@Xʔm����YsZ9�b"ObȀ�FM�G�$�GȶgH�]0�"OtaredѦH�T"d	U�IEf0��"O����)	n|1��^9*E�`{"OjI��l���13��ؙ2D� �r"O�l�h��GFj�b�-X*/����"Obk⇈���d�U��8Ғ"O���p�Ǚ�l�`[%;yްY7"O�q��%`$��I � �"r"O\QB�kT�*kn4��U���t���'��d�E��"vh
$Є�r��/�!�ιHJ�UH��hS�x3pk�^!��<}�U[%A�5Z���I`
�M!�d�O�&e�bP>c�d�9F�j�!�ċ�\d�η[��(�X����ȓdeV5;�O�8�.��a�_F`��S�? F�pN�bs�JU�fh
���'#�I._�8[ő�L�*H
0^���5��|z��C5�Ek��W�Y�,!\��ȓ�6� �$�@���{F�`¶�ȓIc� P�D9e�i��avb��ȓz��	��/_)��@[� ӰA	���B˞��a��*�j�2��)wo�B�	/��A"�| ~\�q.�fdC��LZ����mԓTD\�H#�S��@���O�������ub��i�%r��du!�Ԋ6��P��<�qP��Hi!��¨���#c�E�����dH O!�$Oj<]
męEx�8ٖeǱQ,!�ę;���S���(]�(���J52!�$ˍ&&�H��m^���\� !�d�/�W�
D�\MiAZ�U0����B�<	�Ԉ	<,ipuy"/V�X��� j)@(^%X4�dCo�ȇ�R�֘��+M.[:�����P����ȓ0���V�ֈ7����G��z�f|��7�X@b��W�Jhx�+3G��������ޛ7���ѯ�8�6a�ȓ�*�P7o��k@���9@����?��=����eY?�ܥ�7�"nV�9�'�a~�Z�G��HѲEΥ
V�
��ʘ�y�Z�*y"�g�|����sl� �yB��wC�����3mUT�1#+��y҈�1h2�`��M&X��BK˪�yrIցL+>���#έW�Dy�&���y�M�vB@�Uk��Y�������'�az�Ä8Zpl*�� �J(�)�?��.�S�O�m��NK�6|A���6�4� �'-�eÁ�L�j:�j��� ��)�	���d�|��A�'�
!������D�!�O?8���{�B\�X�R!��'��:�!򄃂���z$�6<��\ٓU3C�!��%c1 Au�ކb )�eٴF��W����ҟ�&?����Q�\�Y�ˇ���aA�6�D-�Sܧf,����R�#v�xA��w:|��cMr$�r��w�Rԁ ��#\F���r~"B�N���TAY�4R"�c+@��y�lDCC\8�fl�*�����I �y&C�B>��k ���"��q�/I#�y򧋋}�5̍�L�(|إ�_�yb⊠QT5��I]�@�!���'�ў�O�dr+]�[��)аc�@�	�'l�Qvl�5ze9%bǭ1��e	������@�A�'�ɞ�(���ÿP4!�dL�M�Dl�N�=8�؝S��R0%-!�đ$D}3�-D�y�(�2�f�]~!�C�H���{�p�Х0��'B^� E{�O�Z4��Q�SZ@��������jO>i���)M�6��ԉE�W39�liu�=)�!�S�d�`p0e��8H�>���&ص>�!�Y�6�~���F.&�4��%б8y!�K�]j" ���D�p�P�Ś$S�!�$WL������!<�p�ۆeƸ7|!�d	�J�p,��0Y$��{��s�Ayb�'_t� g�W�ap@Ш> /���
�'lD9�a�~�8�
�!�nl
�'߈�ˋZ�i0�c؎E����'_Q��	(�p����=�Y��'�J�b[2x �����T�:Ȉ �'�h-���5��9t�*B�d����� �Q闂��.X)t��~�R�"O~ɠ�е ^L�HB� -J�pF"O>Рs�Q	J����+ш:��HE"O$$�Ԡ�w��mB"�D�62`�"O`�ض,����QUF�)� #�*ON��I�u'����	��J�'��A�gF�z,���32j����'��IZ�m��
C\I:�&T�ea�'Q�!p%o�)L
��V�������'Z�=��͌�@��9���X2-
�B�'�j�v�ٌ{vX����ɺ�'��)�e�Ftļ4�v�����'���:��
F�]d�"jer�x�'�� ���;�h BB�MMڡB�'��1� �X���g��=C<`�'�V�*B Q�&o�A��C./�8A�'�L�ۡ�-,ފq��F�.����'ό�C���+Z�a���"�\��'tŢgd�4�@�Ffl�ik�'��!2V&Ӆ >�����Ι�'���A�C�,�� �>��Q��'P�D@��A�jl����5/k�K�'x��(5���
�@�&EK�%�� �'r��e�Q�"�n(��Iί"���'*j�0�jODMn,�F����{�'CI��HϘ$<��8�!ҤA�m�'M`���G��;�PȹՃ�]#2i�'��H�&�Nk,�aȔDؑN�	8�'K��rR���e��cnu\���'�,顆ϘR�̘(�EM`vN���'�P9�o��hT��Aw,O�Sp�b�'���0b�%f��k6 �H\<��'P쉓�,F.�M3р͏9UT=��'�J�p4��h�`}���>2Pޝ[�'Z��#�X�f�h���,5���'�Δ`n�"6�. �N*&F����'t��b�Z�|�`4)"�J�!��q�'�t	��;P�֐��� 2f���'��������,�^���hF�����
�'�x�P�&��- �._�����
�'۾���O�
L3ؑ8�!�9(�q�'����6e\�t��Ϊ7~p"
�'���sT��F��v��@3¹�	�'���SrL�4Qr�7��*.en�
�'��5V�"���K�� ��*���'�0 H�N�Y�z=�q���"���'�R�QcW0��	��Od��5H�'R��� c�2ΤI��D�W��hA�'#$���@�{�T�o�Oή a�'-��0�͋�`%�`���a�U+�p�<IօU�l�2�%
A�qEi�<�k"?J������+X�Q�Ώa�<y������t!u�&8LTr�]�<!�MY�'�n=;%GO�V��lq���Y�<a�FT-m�f�8w�+�Иm~�<��ͨT�E�P$ȏk��)H�"�|�<�4��� H�q+Ia�L�02BD�<��'��'��ѱ�\P���)Qn�@�<1��(y���`".L�>Ӯ��S���<�l�5>cJ��S&K�[G�|{D�Ox�<���2-Ƙ�"��q�q�"�Lx�<�eiM-h��B��cŒmk�fMt�<y�Hˇ
���u#�W������l�<Y��'Q�0��pj����݊2�]j�<�  zp��9=���]z��,�r"O�%y4�s7đ��Z)7t.�A"Of�z�J3f��1C�@P���B�"Od@�OXV2� ���	2wgq�"O������}�Z�o�z<$�:�"OR�`Fe��@�E�UMˊU,xк4"O@��NK=ʡ��E�|$:}q�"OnEYBKѱ�H�1w��=c�ʴ�""OM�@�&&Ff)ha��%�h]��"O��#�g�zt������}�	�'xj�)��	�q��u釫^�eo��'�x9����z� P�U|j�'m,@��ٷ?��Py�P JD9	�'Xxq)��t�����G�Bk �*�'�x��E�P�Qkȳ��Ք�^1i
�'Z�x�%W		�"�`�/��M����'��)�@�	��xs���'R`���,DK$ 9cGn�����'�z}1�.�uj���dI�s��%��'G�%S����T�3�6gq<j�'�.�2ց�U�hr�@>^6޵R�'*� ��=�U���O��H�
�'�n��a♷>(2��S7�{HC�I�]j���Q@A�Jш�gj��$�C�I�'Q4IB3'6GI5#��:"(/D��2�A���If@���j+D����N�c����K�}�\L�B���0�S�S.Shh�FX�`W�C䉕m{�i1�@�N�h�-g�B��u@#���-���	�B�	�n�t]3�N�5	�գ�L|x�B�M�]3DRQ����&C�`�nB�I.)\(�@儴#�n� ��
'u�4B�	=2��m��,k(,%h�>(s�B�I�A%�0�X�*�
9XS� �nUC�ɫ���V@r����$�q�C�I�A���r4΃O�������bC�ɶn�(b EǮt���f�
��B�I�ڶ��cH�>X���U��:��B�	>{��a�'F�6�����C�I-"}��pF��U6��v�=D
B��*��ku.G;O�L�+���!TC�B�ɚ�����#=�0��"G��TC�I�h�tH�%a�+0���.DbL�B�	#G�J9����?q��Q�v�0>��B�	-�M*�!�7&l��!�ХI�B�	!)�B�	B�]�@�ji�!M�(HB�'�X=R�n�j�J�#�7?B��'$_�d��� & L=��D�:w�B䉍Ls�M@g��!rP���E#W��C�	"�^m��W�x5|t*�@�_8C�	�J5�9 R'��5X�s� ���C�I��,�UM�)�����P��C�({���"��iX�r��C�!����/֍H0�#Uˁ"��C�ɤ$�ĹqɊ?p�-[�˅�b��C�I��R�ˆON�1*WA�z�nC�	�f�
��7���=5�0r��_��$C�	3@A�R��m����"�ZK�bC�I��4a2��55�x u�٠m��C�I�}�H=�"c���T����8lC䉓0���?�Dz�ƕǘC䉮;&���$
�1rR�4!��6�4C䉝0��й����A��Z��B�)� "���㕲$���J8Y|�@"O�k[�_�Te9B'Ĥ[d���"O"|���~��q�`JH����"Or���HԖP5h��RJ�@��"OxP4�ī5�⁘��,'� �"Op��c��K<X��7O�&P���"O0�R6Q�!�������I"�"Oj�GC��b ��I� P��
6"O����Γ�P�
y#ti��1�naP�"O��z�΃m��L��8�Xq�"O�)�e!�H�P䨒��4��yY�"O0�Za�v~D��Ӑ\��D4"O\-D��?AL�fK�!W���"O��;��%@�z�I�I�vDr�H�"O��80�s���ƨ�-9P��6"O\������R�,�g�))p1a3"OV��E
PT���a��F b�ځ"Ox�ٳh�p~�1�$"4"�(�""O�3GA�ND�`cs䔏b8�P��"O<�j3�LF����Lá��1�"O��P1�܅<�,-R,O?"��I��"O���r`׵��aaH�E�58�"O��2�E�O~|�;$m��"���v"OhZdHJ�J��Q��,�{(���"OJ����a�u�
h΀h"OD4c5��:�%�<`��@�"O�Y����Z~��W.G#�D`�"O��Ь���plj#�X�\��b"Om
�f#Sg~%�ejn!Be�%"O���H}fX��葷p Z��0"O�	��֧Ĩ#d��sH}��"Ox��5'kH���ԁڠU/ �H$"O��㱤Aͨ�1 �!�*-�@"O�PaF�U���Q O��r��ұ"O~utO�-*�3�����̺�"O�!j0�ƚf���5���t�"���"O^,�#G#7���aAK�zΚ�"O��5I[�-�`�s ˋ��] �"Ol���ߚP�*1�Ǎ�=�z%	�"O��If�S�3P��5R��j�<AVa�#}*�H���[�!���v'�j�<q�K~����
9KX�)��h�<��#ё`9�����N^p4ǥQ{�'�ў��Iӟ�@Q�ݴ}��钲���,����.D�л��R�M�F��A8�ƔK�1D����%��w���U�Գx]j�Z�-D�tI�l،ae��ra-Qym�[�)ړ�0<��jMs��q'�w�r}JSNA�<�/ݞl�E�Ǝ'7r���T�<�ME�o�v�8W�5hv�a`��F�<a�GB)'!@���*{���郮�<镊�oz(ؔÍ�{��]Yqj�f�<��MԔY����	�:p����0�Of�<Q��,.�*���3%��ě��J#5��,D{�� �a�� x���b��mJ	(P"OL��5���E���C�I9$Ұ(�A"O�]���ׄ`"�(��̧J�0QQ�'��O��J<���W� [V�Hu΍@�	h���R��4uSy0�Hձ,��ģ7�z��=E�ܴ����)[Ɗ���cŋ |����|�!t(��?l��	~r|F}R��"��u�S痍F���r�kC�B�I(�Ћ2b�[�ҍ�t��]��B䉂h���g�7o�l��F��
C�B�)� �!b@��+Tfu)C�7y��! "O���UR���$E���hr�-"O�B�V%�ȸppbT�V����'����~�5a�L�M�m�D�曆
O��(!C]2g�����/��i�9��"O�%���-ynPY��sv�e��"OpAPVMƯP���l�sl��d LO��"�ECL-@,�`ˎ����5"O��ȳ$^��|��I�N��*R"O��KwGTJBy[HB�l���"O6���=���lq���r"O���$��Ll}��o�cw�QH��'����<1`H�(�Ju�>B~�24CYO�<��
d5<��<N����J�<���1��x�r��"m�]:��H�<Y���2An�K�Z8��$��A�<A����9QC�Unְ� �d�<A^�G���B���@�����M^�<�V.W3RX��&��{0��U�p��hO�Oǜ��% RF��e$
1Ǟ8c�'�d�f�10��a�V
���L��'7~���ɔ�w�X4�ED��}p�ȋ{2�'s������*�ȱ�)_fz"���'Fa��'Ќ�O��i%��@7c����<���$�$�<@)��ƔJT�<�#�%9ґ����]�hR`��-0Ejt�L�Iݑ�G{�����>��=��#��dǈ<+�\�Ѝ���e�l��dA�9�)�o���f��$��(��ꄻi�uk ��<$\�
�3��.�O��s����%e�ٲ�l��|@�kW�I\�O>�mE
�d:>��5��
CX(��'6�J'��6U.Dp4����k�'�ў�'�r�Qe{�f��7nX98��,�ȓ~m�9 �ʹA���0�'Q`�N���-�� ���_�"�(<*v�>bYv-��@=򸫅��4E/F�`�� �܄ȓx�8���9<T��J,̄ȓEPMBv-�0i�����VRx\�ȓ�(!ħê9���@�+P	7L���Nt`!��&�3\I�a�"��(�L���VjL�D��1H��
���ȓfAd�SP�Oܖ���/H
���ȓ1V��`-��J/�T郑L\|��p�"��U`O�
����#�s{R0��j��=r��΀'m.Q⦇�`��ȓ20.q�#+��C݌H�1�?;*UDCO{�O3̹p���S�dp��Ⴍ|�y�'�r�ء�D�%h��#ع `�P�'hT�®��kZ������n��'Y��2���1$��+t�	�0�8�{r�'p���g`͓~!�E0����N4��'o�9� ���v����B�І	]���'�:�Q��$q���Js��{,�|`	�'唕҃&�*ؙ8/��xo6��'|ź��ޞ@�n�É��le��
�'K
�:�&H?g�0T!��V0/~|��'l��4���*�(�Pf 9��B�'�Kٝ�����ͼT�J�8��c�<Qq�G"+���X���Bq��G�<	1�X�2�x�+���rم�A�<@D�!CD��0�I�!�P��@��<Qt��5A@H�{Ҿ��G���ED{���i&>�9���Vjr�X���;YERD���y�C����a!P`ҎF��@�#�� l`��� $5���M S��sGG
&`N�Z"O.]�ʉ�#�5�W$�<t֡�"O�
�D�mԎd۷�,TmT��"OX�£kN><O�WL^&�"O�aON�l�e!���0����"O���'cx	�����5�V�'B.��'���4!�!Y���JL8D����'���K��tHD��#P"7r�d	�'���a�˫}9�D�Ǆ|-pX�'^��e�./�T�w"��B.ܘ�O�e:����ɍ|��ih�EͪY��̔�"2�B�	���5�cI�%^����螺R�����D6�g?�WOJhž�A�HϚ^�R$�)h�<Yd(̒m�V1T����H(���ޟ����=�雒����!	5��f�>��Ie�=o�h��,�) ��x����)��ybቇ�f� �(MRT�!I�UT�C䉸`A�H�l.V�~h*�@�<=hC�	2t�UkdOX�$~X��Q;Ih�'ў�?e�%aNyH�ժu"F�OK�Hr�8D���HK 6��,��0��\��I5?a�A"h\��`k|�Ϋ-�>8��j�I&!^��� ��dV(�N��(f�B�	%xy"lj�HW �2��0M��'2b�̅�	�)5�l�`O !ah��蕌Pf���t����O����%���N���b�M��O��C��,P�gJ�zjt�[�)���C�	$���b�M�(�@�UC�+Ue\B�I0u�2�2թ�1�J�Q �Z�~r4B�cHP���
N>vPk�)��iB�	C�P��L�>s�4�b�E
�>Q��ITX�P�!q���T�V�ap�6H�!�N�+�b�q��̟�0u�@��3��V
O�e�e��:5qՇ�ℜ��"O��u�O�H���Q�gD�u���3"O*�!b�P/<�P�X%�+��|�ýi'ў"~nڮ<�rq��5�p�p�h�?TЎC�I�u/\����[� `�a6O7]��<�˓ \�5�4��9��J�������&����r�ɕ^�Ќ��V�F���	��tA�֩*�fCEĔ�H#��Fx"�i�ў��>E�j��k�*S3�1 ω�-�\C��+��xB���.j1�F�Z�pB�	�F�n�u#-*RH	�F�Cc�6B�I�E[��bAE ,ӄ�R��N;��C�	L�`2F�I=t�(��A�!lC��~b���t�� 4C@���O-[q�C��)d�d9�3�6_"m�g��~KpC��5=��QKF�{�D$f�G�7�`C�	��v��4�Y�cZ 2� �8.��B�I�	:��"�1�,$�*{TB䉓(Lu�q	Z%h�
 ɡ�^�+�XB�	R��9�I� ��P�)��X�C�	�2��� �ϪHͺqb��]��C�I�\�007g�=iR�qq��ĂD�JB�ɇ�n$q䢇�.�P�$���B�	�k i���݈w�*I���ή<_�C�IRi�\�6�18�&0#��9=�C�	�l� ��,�eɀS`�>>}rC��a�l�c�X�h�}�U��WC�	�Q&�5��Ƿ@��0���֛G�FC䉛:g�qB�?d�P*��V!�2C�oDY�ßl
�`��H�C�	&4s��r�mT�5D,!؆�� S~�B�)� ̕���H[~ 2��і\�PPc"O��P���
o����
��8��"O I��d��nTAR L�l���"O�Y�BA�;��� LK4�Yr�"O
$A7lD;>�ԭG-�o8|X�"O,��
�8����K�4F��"Op��(����a��tr�h"O�X ���'����"*Q�b��1YD"O����	t�>5����M	�T�"OX����Rw��F��U���y�k����yxS��@0� au���y"O�, :�p�(�C�Q���	��y���!	�P�kI�	���9�H��y�ƈ�ww>���C s�<e� �@�y�t�c��'��\���c�ZlϓAP�Dj0�67�]C�O5x���G|�ɛF�D��-�o�P�PN�#�y"� ����ΰZ��4�A���y���T ���I�\�H�"0�X��y2�ۿr�p��IK %��$����y�n+L��Ȧ��VFyH�(_!�y2�F"uOL�i�
"��qj���y���')PVDB!�Bxm�)k�ӥ�yң�)s�fU���B����L�5�yePp($�i׀Tcn��1�<D��)��((%�恜�NA��� D��C�+_wz, bϟ�Z�勖�"D��BF+�� ���o�M.��g//D��D@R�p�ޥ[�mF3S8�T��-D�T�s�>&��I0���0���K�'7D�x�(:]Pt@fͮ%���/3D�H�s ��6�dHѱ��%v4���$D��`��P�� ��E@�R���k'�%D��� ���H�`!��P�r-��<D���MK�ih��4i#N�8�
Vk;D��5�X)1O�T��TQDۡG$D�$J�`�!"�X�#�99`�T��i%D���soG�/���9�J^�[]fhѭ)D�h��ǟ!�13b�_�J�4�h D�@��Ҝ=��ī�(v+��q��+D�Ph7.
&���E��i!����(D���*�/feΘ�8�ds0�+D��c����vb4��kE&@��ċE.#D��pR'ӡx�T�3��/�����!D� �`� k�ǆ"�����'*D�(��dĽPE����JH�D¡I+�	H:0aY��I��dP�"A���j��<:ֈB��?"2y�D�S�hק�p�P�;AS�K&R�'ឩF�,O^I:b�K"x�la�旹=���e"O�) �π\*��C$+�a ���s�l����9F����$$>����R�^�BP�� E�i��y����\�NL����k�hIn�GB�Iq���t�I�|}y3"O"��aP���7kb��f�8��hj����	:?a� �9ҧd
R s��8�ތ)��:.����ȓ��h	D�5Q�0���얊=�X��Q�D��E3�(�Ol���l�X�g�I/W�0�b��vy0��D+w��B≡M0� d�͛V�]�'�2θ+T�؃DLȌ1e��z�Ve��I9'њ!C���e�`��;C2������5�,�f��r�t��dZ�,հ]����:��tH��Xs�:��ȓ �	Z��Թz9�Q���׍+Ol %�P�k��[��(2BŲB��F���֖4��-�2e>FF�ذ`��yO�85Xك%�3&
�Us�X�<�N���Ô�[�89�ɵ6�����L<i�쌗4��Q퀍W�,\4(HcH<1�4/�=��LӘ*�M����T]JY�R��k� ���$�p=�`@�m�*xs��Ņ�
"�Ʉ�	nj��%(E�+T�сH�� \icF�z����QDQ�Z�r!`a"O��2eOt��8 2pò�|�e�95 P�2aB/j(G���4H��f@��-���P�+�}�<���^���B��&'0W�+7.U�.N� �� 9[3b�?�'���n��=Z�J�(�?y5�ݢ�'�����L4ȰK�!���Fo �X�bT�̋ ��{/\�
jT��phP�츱�f�;�p=t��:m������2}Гl��|�S�q�*��`"Ob=� o�RQL�
îG7�\��%��ӫV���r��i�����{R�I7g�� &�U�!�� �d����9W�i��6y�!�	\~`"�ևXQ�\�!C�6R�!� ��t	"E�Q>
�p�86�Xx�!��7*� Q΋�V�7f\9Q@!��-ҐZdiFN����4݁S!�$C0@�|X���!uy�y'&�*.W!�G�'DL�
�闱xX�UXG�J%O!�ę7"���)T��	4䍒G`��h8!��ª1�>`��b�N=�t�%e�--�!�$?pjMc��N~��� /TV!�1j�e�3��5f�ܛRNS�!�D���Ή�S	�0�mkUɑ�!�$V_h�	��搘=��I+_�Gl!�䃀2�&%3`�y|,��J�/+S!�DȯB�~�ZD�G-���p�i�}n!���Z�D-�����4M�H�7`}!���Il�H�T.O���u�qF܌r�!�ҭh�P8"S�x~0�ˀ�)}�!�d �N���2D�~�
���i�!��3^�@�GL(w���X��"p!�DC��a��b-5&i�NVs!�(�$Hs���UR(@O�0�!�.���E��F�Z9��0(�!�D� ua`mM0P�XP�H�x�!������4F�M��!�H�?u�!���l�|k�jV;��(*��L�B1!�D��.�N<qu��X|B���fϽOV!�$	��04��%
c���d�g,!�$E* �M�-0�<�a�m�{!����0�Vk�a�B�ɐκ�!�D�4�����˒�H�ؽ[�� C�!��ܣ"���� �&�Q��	,�!򤀳J����O�>k-\��!�1m�!�d�FR�pRj�9o2�D�f�L+i�!���	�l���3��]�Tn�>�!�$�8&:9�4O�G\��Arm%*�!�� ф�p�K���4��-Z?x�!���C��0� ��/�F��e[��!�Л�zac�yʄ�S�7%�!�D�/���œt�:�"����!�$��*KK��K����ĩZ�^L�x�'�Zx;V	0@��Ȣ� U�,T��'�T;��Qx:�S�"F'p'��`�'��q���"I������
$"rڰ�'�hy0�����I�
�nz�1��'B^$���Ψ+`^����e�d$ �'��� Z� \��i��YL=��'�jԈ��eUp@1�@n�F$S�'En�A�ME�.ph���eR$�8�'�l�C�F���@V�R:�EJ�'Ҳ�4�
�tg0DX�+�8H8��J
�'��er�J�.��6� �~�Z��	�'�]����9��5�Bc�#b��r	�'�����ڈL�Z� R���PS4���� �8R�熃F谺@���+��"O���+ �̨p��D�	���{1"O��r�A !0�1:���m�2��D"O8��L�JvH��!U`�iC�"O$9Q�J,p�[�V%I%qq~�"OJ��ӂOt"v�S�	P�D	�"O����Ӌ<��	s�jΎF$ }��"O���B�ؠwM������ &�	�"O��q���l9�͗�:���8�"O��{V	 ���v%[4E��Ly�"Oء�� �jH]aP��'̼]�"O,� J����`+�B�;Z��������-CI����-%wڤ�Ʃ�7@��R�-ؐX�!��R�&pH��qEl�Te������5hĨ�Pxr��8{�K��
3TzX��ˁ�WY� :�)�)qOd��a��"WF�3����j^���"OH�rb[�RQ��*:�I%�� "B͏PqO>�rw�R�]\Z`�Eɉ�8"�@�*O�	ˆL��TJd	��Ò2bn�h���R3ge�t�ǓU���P�63����c��!^����T����I	[Źqm�3%�~��6BD+"��C�	(z|��X!��t�:R�J�2A�'��������N�DaU�\KSd]8�cҬ�yBDA74�����8�tP{áF�y���	v��ɛ���3���R�Ŗ�y�N�	p%p�E �_�0�[�i��y��\�B���NH�W����O��y�"L&-F���W:&�y�%�+�y����a�� �G>(����y#]�5������=M ���o��y҂�3=�6�#�	�zOJ�{��Ֆ�yB�]�&l~��Ӈ$r�4�R>�y����%��q�m��X<�a�)F�y�O��b�DH�h[��%�"�W��y�@��:�b ���T-½�#�M��y�!Z���#�E�s��`b��X��yR�V�q�X1����n9())����y�)�[�0�P��׶VϬd����y��3db�3�F�_���D-��y��Uw��7Q侱8����y2�'#,.���$_��<����y"OQþ�H���>�0 �7����yr�_�N�������+x(Yk��͚�yrNʾf`�+&JJ(mqV���yR�Z�j�X�Ph�?w� � %� �yb�
,x,8x���{A�=��"�?�y����2� �9�O�`	D��y2���U_
T v�~?��V�
8�yˍ��0����Xqq����y��ȿ*�TX�B"�;p� ֠�y2��T�HQ��-t^�(�&�?�yBl�2\�8��a'_j �B����y�Nԯui,�3F��ȩ���y�ǘ�Q�9����l@�@�y"b���Re��j�ypt �[�L��'�$TEa�
4�� �J�2��h�	�'�
���!J��;S15Q|�	�'� XюB�We؂�ჷ9�ɛ�'Q�I��F�;���R�`A0hT��'^�0���]'؅k�������'6nx	_Z��q�($�l��{�<Q1	�G��(�5��z�4���q�<��j�5[��źe���o
�8!4�_v�<g�W�
P���Z3(�:�`� _�<� �!@��B�c̶Q�2Jָj/f�2"O\�Ȅ��<A��(YeIQ4x��XF"O2)'�P��ұ��K�5PW�p�D"O~y!�eR�'o��-lV��"O��q�&�4�ض	 `Xt�P"Or�8`/E�{�Μq$R�h�"O�( ���["����GO6<�d�Q"O��s�E'��!�+]D����"O�ܨU`� [���+��`�*"O���g�ǀ5��u��N:%��Ų"O4R��HjP��cL�2�x "O�q�ȃ��:�@����j�
S�"O��4k B�̍r'@GDj\c�"O�������œ� �\İ"O�`	s��'!K���[������"O�t���K�"���^�H�����"O�� Dm�}.Ґ�#�^�y�I��"OH)��IP�,�Q�H�W��!�W"OV�*cK�0w.����y��D�b"O@P{�	�m�4%��$��#��MГ"O�Q@BH���C6L�*z�@jA"O.L4���^� ra��Q�$x�"Ox	0�LCp6(��LŞ}Wtl�"O� �M߂���:�&�#.h�g"O`�jUj�,)�H�C�fŘ��! x�<A���Mߦy�$+�^	PP�Ao�<i��č,�4��+�qpd<���Za�<q�WL����fH�6������w�<!LS1�xEA�(E�s��	kBs�<�`(�1֪e�゛t������T�<�%�N(O���%�I�7����`�G{�<�&�¿+Z�)���L�)e�L�<yǕ�F�(y��U&lXt ���M�<����#z�D|�v���z���%�V�<���� � �d(Z-q�p�CE�<�DǤ(��p�����p���ZK�<ɒ��-IVkB��)�T�1���J�<	T� �L�a�Yz]��&�@�<T+W�_�򁈷�"B�д�Kx�<I��R��\%�t�4Ow�͓��t�<�4�H��2%�Ѷ��+��
u�<9���p��(��M2D �=G,�T�<�`$�,rDPXЖ'��K�@���d�S�<���6N���X���̒a �I�<��.�
; �K�CB9��rm�C�<���ۖ\eX|�a,ף h�S7��U�<qv�)&
Q�W��GU�ؘ!�TP�<)&/�?�����A����i�%O�<)!d��	(
i"��yqH���^@�<�3��el�E{�nݗgF��4��u�<����On��sa� �2}{�Sl�<��
(�,�!���
0���l�g�<a�*A2 �R�r@���4>�I�r+�D�<ɰiڶ�d ���j8-YQ�JG�<a��(�^�z���n�� ��!@�<��>m�,�qQ(�|D�3BB�<y�G�m�BY^ip��CVz�<ѷ�_n����1�G�
B2y�`Qq�<�Nݛt��`�/�oܴ�T��r�<�W���%x�}��:~�!B�$�U�<y0�ܱwl�<+��ô'�N�4u�<Y�Y�B@��v"ؙ�l�Y��N�<����#+�����J+X@1T��E�<��Lӈh���y�	��/��0�fLA�<� �!����xg ���#6�8ؠ"OH���)���VbϹ:��� �"ODxSƏG#MG�`��ϳ0�4%"O쌁A ԓ4=nL) ����8"O"Ez�BŃbr81� Y;^�� r"O�<2�ZZ���w.ʮg�ưcA"ObԻ�W$.�8��X46P��"OXH�ɾo�Z���˛1����*OF�X�AX�R���R�M�z�4i0�'U�MK��۲P�X{�͕�s�+	�'�&�s��/������'d���'��! ���#0X��r�[3k�a �'x�83�@=��ƯŽgl���'M��pv��3}���5���\�'��l��i�/I���kU�!+(`�'Il<�g�ў:(�ܪ�6Vh)C�'�����O�44�����A��'Q�-@�:������K�����'����T�Zt�nѤ;�tI�'���(��5{��-k����l�1��'���; b��C �TBG���cZ�QR�'�ț�	'pXpY��㛬[�P��'��yjš%|�*���b��U�Ѡ�'��a�b^8�t�Y�J:Sp����'�Q�Պ)� ,C�K��K]�U�
�'/r��eT)2ݘx�t� 9����'�����+^Ԙ���cr�b�'���d��e_t)3�N��dv` ��'�`���
�H��!ba��l�i+�'��2�M�^�����;_�ܺ�'N�p����,� ���ėQ���'4�jg,ݐY4xL��
 �Q�]�ȓK��(ر���F������D�g���ȓn���2"Bmh�T ����?�=��QT��kV��4N7�4Xҭ���Շȓ'H��`�/Ir�[�
G*k���iO0=��J
'x|3�-H�
@$��ȓZWb4Aգ��0�h5sw�b<z����ذIN<x�`p�7��=�������@�w�]�(f�d!�6�����o����3���I�v�z���G_����Z[L$	Ҡ�0ay�z�N�ve��ȓȠya�Nѷ�N	�у�<h%�%��1*°�&�ʛAIJ|���_�j5>P�ȓY8�,x`�$vr��3Ӎ>+V
��ȓ�F�IFjT9�t0)uj�9�,��ȓT��l�Q�W0\RY��\�`K�`��|o�5r��;G{`T�C���	�L�ȓ��!`��(�f�ySN��R��Y&  �L��h�{�Lbd�$�ȓxܼ���̒�GA|�&��J��q��'�
M�� D��3�{"r��ȓf���!eM��" �[0�ٿ��\�ȓ/%��:gB��&	��7�4:�0���dD.��c��\U�8��ʹ(�F!�ȓg_~�F㝒T��	�����%D�,�ȓwʆ8���\��y�r(�l�؅�(��QP "E���9X�8��b*�Q�Џ/�d���J@2w�����*��;4���	Oʑ���
�I�ȓ't ��6c��rï�:q !�ȓMƜeX�D* x����y�^̄�j�U¶�V=~o�����ՐT���ȓ9d�p�m��C�f qCg+z�m��S�? ��ᷣЅdb�I�3A��$�ry�"Oj�ReV'�<t�"�Ϡm|�a"Ol�ff>c/���%�S�$���r"O-) ��I�.-=�X���X��y2�އmhV�Y��:���"К�y	��J��񯀕*�M�Wl
�y⍀�r���G�O�z ����yr��9�AB�9��BB�M*�y"������7.
��L�aƗ��y��<>Up��dL�h=�|�wc���y��T��9b��jA���@_��y"�ޛs�A F�!~0`���j&�y" �u�B�:7-�q\رţ��y؍A��$��@�jhvdr�HZ��y��&��b���1W
���G4�y��D�J����,����a�W�y���06$��Ѓ�,#������y�[8g�l`r�W

ΰ������yBG�M���;���{�0i�0�A!�y2jj���8��ؿr�V�� ��yҦ��>�v�׫c��\��)���y�/Ͻ%�8Z�ǐl��TX!� �y��7�t`�a#��Q ލHe#T?�y� �/�ݩc���d��y�$�0�yB^�4ޮ�Q�X9T�,9�ι�y�� �,@���rb9��O�)�y���>�>�S��>�����y"�2t������>$�p��l��y�b�inPXp��H)��ȵ�yr��jI�uJ�ˁ�G�-ORA�ȓF5b7%�
`X��F��D7n �'�z i�5
��f�i�Z�	�'L��� ��_h���	�iÞ���'(�a��̪O�3,�:>)�58�'���C�V�	�+U�,�����'� �[�~�2�$G(S�'��IV�^�5�]�"dT"�4�9�'S���	�*j�<LH"��
�a�'����c��"�z��Ș��e8�'�k� �7
��K�2�(H��'�x�;���=a�E�'e �?�E��'�R�G��0��@�g�ԛ:�N��'J��n/�h��� �l��lh�'|����@��c�tr�M3�''|E�@H�;t(��
�jԐ��'��PA/�3��,J�II���'16L�7H����EL�1 T�S�'��i��#l�Q;�GP�Y��;�'�M���ٙwph��T`%R`����'*����#�h] ��UeҎ�I�'�0��U_:`�^i��˜�gz�Pi�'�Z���a�/T^]"��� Q�2���'&z��u<0�R�H܌IZ�'�r�[c�V�#�*�@u�ŭv��
�'���{B�#A�l���%H�	`i�	�'�\i� ʌ-{��{��|�D��'��H�.�'��q�E_�W�py�'�Ȕ!�AG�f[��{�����H�
�'Ĵ	{R�2Ff$-P���|��ى�'q���R �7]��;���h�f�X�'YbE�灁8=�(ZE���oè���'Gl���Ne�"\���P�[%�Xh
�'�v���g��P��݊#��X�8H		�'��@�*�zX��OҦ/<����� Ph�l[� ,v��%���4��f"O��b�#X0���BLnshmX�"O~��@)�*~��S6�\�v�Թ�"O̵��4fP:@���d��1"O������e�`xR)�_�P0"O�q�feWW����'�I�f��<��"O0:O��|s�XS��D�� G"O�=�ƣ��8�|��d��nqxt"O|p��(C�8��4i!��7y�|�z`"O�� ]�
xȡ�JC�;����"O*���	�L ���)F�G�p	s"O$����h����j_{�8��"O��8� CԘ�ۅ�k��H�5"O\�7a���AKu��6�C"OXԻH]�JrngE��N��"O��K�a����ڵkћ/�̢&"O��p��P�✤�KR�4FDRp"O�0�!+��.���8��D�z4"Ox)�`�U�|��,�G �9��Ib"On�x�Q[ ����K�d"%"O,�1&n�v�$Y�Ɗ}'r���"O  �.�<E#Pp� h��{+b��"O���t�L�d�Z�P �Q�HZ��4O�(3fll=�a�
YD�န%Ͳc�Ҷi���_�HX�=:@�)��DP2�ы�����#u��R}L��R�':���a��0΀dA��˻E�
d�=q�ŝ"����'8Є(*I�6��D�ꟽ	��8�O>��24�)�S�4x< ұF�s3fLQ�'_�A�J��5�R��?E�$E}Ip��\=� ��	���IN�S�O#XIJG�Mg]��Q3��n�Ԭ�"�5��uTa���W,�m	F��0���ʖ��;��'AJa���ԟ���H:�@e��N�BP����O������/!��c�h���O�O��Vo^�P�|5�qEG��u��.�a���Q+;(�W�SD>����ũ�QqF�F�J!��[�i��dY�*�J� F�D�w�@I��MG���ԷB�u��% dmQ#��dYKB�� �&�������l�4�b,�r� �{�����`
���C9�)�'պ��垄o�, �e�<N��T�A��9 ]�M�N>��� Y��UR��3mSH�'�ڱk>	���e?�RJW�֌9P��O����D�7vg��B��\=_����T�O��3�U�$�����O�f>�(�+��C���0��z�X���p�z�:e���G��	F�P��~���u���P�X��K 腘��U�:YX� �/������9�\��K|����NS�&tԩ�$R�aY>}�2-�\�6�bRg������i����S9Cu��;��·{8��2���[��;�'��ˑm�	,W�����O:�-H���6bB1�k�7��Qh��tj�l+� ��S�5rs8O�˧f[�`�������s��lo
@a�ŀ���O����ɭ~:Ǐ��R���NW)z�� Z���s�*�$�R����?c��O��%�D�U�,d��M�0<�0 H>��m��<�2����h�j5��ӡw��hԠ߱0�!򄎄oX Q�L�ڬ��Or�!�$� U�{�&KE��#�!��1T�l�Pw���h�:lA�d͟7!�D9L��L�بp�ıC�k��Z(�C�	mcS ¨{`d�G��>u�B䉹E�b�@�$&^|X5m�3ּB���`��Y�F&�����IւB�'\n�A�����C �j��\�ݎB�ɤ���*��	�_�HWi�	~xjB�Ɋ��e(w�X)�Ҙ��#�?A	lB䉸}A�9ڠ�J���3wd=T+.B�	�7�LX��/�}Ԫ��c�B�B䉌=89��/��TΊ�Ԣ�&�C�������0#�&�I�Vr�B�	�ΘHe�8!�-�N�wC�	.nE"9a FP�H[�=�cH�תC�I��4@فa�z�v)R���s��B�)� B�y����(�c��1"O�Tpv��h]S��P��<�Ӑ"O���#Ā�g�JD��
<~��\�6"O�<�h�3"��0��W
�ˠ"O`q��/*�(�΂��9I"O�����:f��b�ݮ㘰�f"O��
B'�*�XD*��]
"� �"Oz�k�g�"h�0m�).��-*d"O�A2���P�2�J����.�
U�S"O�$�c��C�n�qVHO��$�=D���_������c��=�%h��.D�@·I��C��I� �%3��[ӥ"D��)����3��@�ђ]v�ે�;D��a���.@��C��""�d����7D�L�Ճ�z�r�0�%��-��]���/D����"�B�إO�"ن��r�,D���ތ C���Ť�#()����>D���'�mè�A3 L s��m)D�,*��R�m�4�zGlE$�"�!D��0i�s�z\"��_#CJ��Ĩ?D��������Ȭ��>E�(|��@;D�Xag#��MQpy�R�̍,�X��7D��ӱI
6�@�i%lK�=��8Y%�5D�0�!#�tT�hK����"Y����i2D�l�F
V��xjt�R:s:D�EO4D�`c5`~�v�v�9Lp�x�D�2D��s��Cb���G�6$;�l#t`1D��B��U+9���I�o �&����F+D�<A�N�D�:&dʕ=��b'D����f�����͚-�� �o9D����R�Q)�-'��@MX��8D�<��cډ|U�];FH>|@@��5D�X�0�^Z�8x�/��k��PXag'D�� ��W-����%��Yy��I��#D�<����COL�`ĉ�d�V�%f D��{�
��7K>��C �� �%2 D�X�D��d��ȗ(S��yr��=D��#�'V0����:GVTu��=D��RTK�/p�Eh�0{4� *�O1D��[�m�J~����E�N(8�M*D�h�-�
G�����×#��Ds��"D��{b�ՙh9�݀&"K�����*O�d��$+��jq�Z-b�@�v"OjE{PI�tT U�A�@�PQ��3�"OhA���|lK�M,&c~|�"O�8�$D�4Iĉy%mW�K0B0*�"O���aU�,x�q�L�:)<�"O����..nq�@_u8��"O��S��(w�ܺ�	�	�-��"O$�C�W�#zReSC#�h��"O�`"@�70�N�#�⇬X��"O(���,	~H���Q������"O�U�BÍ�N��6AR7�(��"O0dp�ʖ�4)rP��B"k��ܱb"O֕X�(� T��fS�&kr�	�"O�\��b�6NL�ˆk�`J�{s"O84��AJi~��3�4w����"O
U"�`E4M�(��N� {�"O"���O�~��􃌩 ��5�&"O6�Z��[�����C����(�&"Ot��֦Z�\��"�G�$p�"O�`��ƚb��dPf+�*2=D��"O
����&CPl܈�
��-,�+$"O-�PJI{�:,	k �H��"O� ƼK�BϚ% �Qa�FL�J�"O���O�8GC��:�lT;y-���R"O�0����M4as�"[�|&�Xg"O��طeL�w��Yvl۶y.*mq"Oz��*I8�eAP+��lH��*O��b�d �A�p8�OF ����'�̥i���}�H$�Q�ɒyT�x�'�B�%
��#��L� � ,jQ��a�'�����R�Fz��WE�1h}� ��'ZaY5韍=���昩`tr���'�$�a�dӜ(3�D��S��"OHH8��ϧ"��]�� �|�"O0��g���᲋^�~t�R"O�T'��w�z�ʳ��m��ö"O~lrt�� ��K_���"Ou�7D?5$�6&�G�fh��"OԹpF�S� ���W��Z�Jh�"OT����P�  ��� �(���Y�"O�|���߫z2r��VDG���g"O(��D�%_=��1��D�C̒��0"OB��� ��5(��bΆM̉�s"O���1L��"q��B ;�xa"O�C7�\K��]�4!S4��s"O�	���2~���@B<qu�͐5"O���G�;?���a/Ѱ?i�)��"O�l1Ӏ��f�R��u���^b�T�"OX]"��(q�Œa�صmx��xS"O���Fȣj��X�߷;]&�[�"O<��q���qK�Qd��G=Z9x�"O���S� s�Ѡ�\%�DMh&"O�8Q�
�<Y(1+b��*2`S�"Oz�`! �%f!��n� 1�H���"O�Ehw锉g�R�zg�K?H�ԣ�"O �3
��;�r\��ȕ�@=1"O�0�-Yu�TAW�Ա'�V`j�"O�%2Ah�aE��k��=z�f���"OZ�H���	
"|���%\�tZ�"O���Bj�"uw���So����P"Of)���@��p��o�R�0q�6"OF��b�>k�$E�V�+�=RB"O����@?;'*��oŨws0"Oؒ1��vܠ�N��w_NKv"O�؂�jU,*wڰ��U)V�+"O� �֌W�I�B5 S- �[?�K�"O���І׆d�@�]^8���"O�aD�f�0���!U'�4�"OP�x�L�/zlT�$`&�x�"O��J�]�Q�Z��K�+	�!��"Otȋc.? T�أ�V
h���p3"O�e+T
T�^$�<����BNL�k�"O��k^{T��x�ND5M;���"Ol�"���9\f�x���ĸM .]@E"O����Ç<��yWFR� ��'"O��r�H߇~�M�å�#M��݁f"OjD��b�u�Ё�2i����"Op(@4nZ"I�P�"����Y�v"OTq��+�	+���3B��fr��K�"O�L[n�#yp�  �TN�Q	�"O�M�B�W���G��2&4yt"O���F��9N�6U��m�%Y5��!1"OƑy 	D%R�X��m%h�P@"O ��ta�(<�:�,
�
�U:P"O�e3���!c�"��w.^�8�X(Ic"O��id'�V�vp�S��&�.}�"O� ~��)S;>QA�A�3��(5"OB�!b�>rj�;%f�'I�z���"O�y���	��H�"̔:��|�"O�H���僣��c����"O����
� cYYdA��ys %�A"OR)����X�\��vOR`Z��`"O�8� ��:��1�`,G@L�I�"O�cV���(������M$hH"O6����^��IX���-����"O�H����e�M)\'��ȓ��]�X�U(؍6��o�I��G𔌒$cG=!�93���2(P�Ąȓx�.�9�-�w�,�͔2")���ȓ*��|�G��:�N.R��ȓ#�����H<W|p���B�5D���&U�.�L���1���tg5D�@p7/Q�)�ܹh3��+S�����6D�P�C���t�ā�^h7�=��4D�,��%��U$�͛� �'w�]I%3D�(��AO�\�X�� ҾI`��1D����eēZ�$4���3B���*��;D�T���ʎL�.Q�@)��u��)kte8D�V�k]��0)��L��l��f>�y2LI�Q�
�t���MI��h�JE3�y"�)̥���}$VhʇC�*�yr�F�aZ��c�d
y!Н�'-�y����@�NL��Jt��*�yfG�OM���N[�eΈ!���!�y"�9���*T�w`��@J?�y�AF<
����,ƀX���3�y�/_�c�	3y�");R�T��yB@9tNpPV����|4b��� �y"�'{�lM'�E?f���5���y2 K�\���򅣚9 h��@+�9�y�`
upn��E�0}Z�)��˚��y�Hڥ���jb)Jy�ƄzA��7�y2��J䱇��C-�@q	P��Pyb��v�୓�m�&{��y�O�k�<�׃X���;�KġDD�-i���d�<)��ɥ���ܟAV4����F�<�s�S�x?d*'��)�XT��m�<a��G��Cpa��({f �R�k�<���Y�Y}�ђ��P�%˶}[��Rg�<In̠.CL��w��#�RS2�N]�<�	 ht �w'@"�2Y��)OO�<a�U�E�����͜�/;�5�5���<�RI+y>���nY�+��@�7�LR�<y��ij\Xiuc�<,���q��X�<)Š�_��D��߱@s ��c�l�<��\K�H}��lH�ce��a�C]�<�c�K1s��C�$c7Z�qd�_]�<�D՝"\$��_�0���Q�<���   ��   7  :  �  *   <,  �6  ~A  >L  W  �^  *j  �t  �z  I�  �  )�  j�  ��  �  5�  x�  ��   �  T�  ��  ��  �  _�  ��  ��  2�  v�  ��  v � � s S �" �( +  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}��za�@AIp '�`iF�'�ay��D�3������ ��4�%�x��'�za�(Nx�0�A��Y*�Jד��'08!��~��Y�O��Q��,�ۓ8�>�O�q�Axh0:Q)0W� P"O�H��/r8���H�<+�E����<������KO&�0�WK�qs���1b!�D��/�*lx��K_���R*Щ*?�i����>E�$Μ/2����@ΐjG^��w	�M0!�j��؈u��C�pT˔�M<���~�C�SQ���'�@��2j�?����Q	I�"�|(#���'�r�BB�]35Δĳ�$Q1OR�d$��>�Γ>�"䋥K�&\�B�� �c�(���	Y̓<���`G��5A������dV�C�=�S��?�e�}�6=��%W"R����r/DߟG{��I�6�R�T4e�㳊P�9��C䉺e�Z OK4g.���θY�JB�I�'�)�!�`�:�ѡ�BA�C�[��y���F24�$�d��'�B�I�[ǆ�IB����٘b�ȼz/�C�)� ~��NP�� QN�B "�x"O, ����)��U 6n�~��م�O8➨D��O԰��OP�:�����b�	�'�B��M���!@fGo����	�'$jE�*�6*���mO�g�f����HO�|�5�H�QD����mV�l�����"Op���1d@�@��y	>=X�"O�}ѣE�d#�0v@$S� l��"O2�:!��M@�q� M�2�x)�"O��E�[�+�� ��7/����"OTP��&
����n�|��+��'c���å�+|�Y�F��K��q���)|O��	m}�a�2P�-Y��L�Bg��	��HO����!���|�q0�ף��Div*O|r�'J).�P��Ob�X�	�'sV=���Z�\X�d��@�H�tt��7ړm�<@H�4[�,u�gN �d�D9��l�"X'ԅ��J����"*Ͼq�@iG�~M����l|֑ÅoH�1u�1�Ā�����g�]a�=��.�M<ҙ"�ҟ"�2�D{�'}�:��ơ^���箕/�J���'�T́�S���07.Gy�����'W�����0bN��!���iQV�Q�y":O���9`�A�B�X-��xB��5mf�~b�O��h�&�j�]B�"�X���jp�K���xb���@|��@JrHy��k��0=y��[�2�|��ҁW�ZxiR�V�y��')�x"P�ڳ��H!ܬ�iۓи'\���S�G�(<ĸa��5m��'o�t�wG�b�A0v�z�xR�|B0OluE{*�
k@�=.�P8`/X�|G�h�*O,e� ,�e��eHg��hg`��'H�ʂ��.24b@���2[�t� �'D�|f*C��̰�$�Y�ܡ��'w��"!�QxJ��E�$[\�
�'�Չ�E}����P��y�'�h�;1COs�<�ا�*y�^�8�'��ɵ%�)�'b���vEE�>��C#*��s�l��ȓ#���5@�C�")�`T�H�������$�q@���!��i�4����%Ɍ~\�7�F�?��CL��y�i	-Ԋı7`Jd6�P��ϼ�M��O�등M�J?�xb�O�/C�>��p	�h���Ō*�OL�	/NXYza��5Y��5�RRr~���'�$<?�
�s|�Z�]yW��Z�X*&���D|��F�8���΍+R�bYc䧑Q6TB��/YF\`GH
�2F�./m�S��'�����tў�Q#��!,���ڵ�O�d�ܑ���3D�x�,R*jr8�%)$��Q�G'�	`��@�+��oՀ���/ܼ*�����&��e���F�n
'G&3�^h��	%��9��cM2�rf��.,:�����y���mڦ�HO?7�ǨVR �����%F�|���'7�� Bb֧J�B1I'�/t����
�'����aY1w��@��Y�rq��C
ӓ��'��x��O�M_��I��%� 8��}�"9LO8�2s\� �v��2��[Ux����Gx��
�e��mZ�_1 �$E��h��듾?�(O(��Z��L)������9;�铍��0��?˓;��8h��ph��6lǍ1�ȓ��I	��d���R��C�}�ȓ=�H�ӀU�h3XJ��%�T���#��'}�*�&y~���N�2p���#��hO�W�zI�r��+�PـS17���$?�Kj
 Yem�>s�$�p�
ۘ��l�����O� $�Z��E��1�EL��2)��י���s(��J��'s*�'PL&hAreɟ�|�9ҭ �6;���zX�x�ɤ+��c�_��eh��OM|�y�d�>��SzJ|bu�͊/ƈE���" �<�s���DX��'���O�U2 ߝ_���ԍP�3���>�	�bs��� �Ș;��}X�j�1miڽ���:�~�Q�8�-�dkX�5B��R5%�?�HO���(J��3�dT�UFX����,:��Ic��슓�	����6ː�VVP�8c�̮i;��շYf6Y[���.BĻf�M)�z��? O\# �@�л��9IB���2���:.��Ǫ�9p
��3	��~ ղ�'��O?�d����Z$zQ��B���Dz��D]d��!���S��M[6 %e�<�`�I�"�0�V, �y�d�l
(I)�c� ��$�. 6-m���'�.��D8��9Ȕ�`7JC�J"$�0f�I*!��^,[�ڙ��"��1�δ�
Y�?���O�˓�hO�*x�(`(bI>Oa���4̒�Q����i���W�a��&�L��sU��Oz�j���s�8�t}]`E �-Ԩ�ؑ�0D�����Б�+]qNn�$ )D�|;p+I��,p��W�t.>)Ӱ�9D���q�ȅ(�B�X�����'�,D�0�tIE�|L���SܨK"L+D��꣏L1p|���N�
�v��0%)D�t	��M2��q
g��j�@�	&D��ȱ���ydj�;3 �'�,�;�"D� ��f���у��S�Q����!D�yw�_&;�ȃfM ��;pE5D�����X�9'�颤**��|��l6D����g��p
hPD L"p��!�!D��3c{�	���G!r�V�+D�йSLL�4��<�a�B�(�<BwB5D���b�<�V:Ξ(���G.4D����'םA *%J���4K�>��=D����A/5��U+3Λ#��ʲ�/D��ӥ/_h�(HaD(�{��ɠr�-D��zÃ�Bx\�#s���a��*D�8����/uN��rK�"*�E���(D��@��	�y�Ʊ�ௗ�0�Y+"�%D�<���O�Q|�#W��+Ѫ���m9D��jE֗E���`��W���yqN8D�<����Y�����C,�\,gH8D�,36��;�P r�S��h!���4D�@J7Pf5�iF�<��0K2D�|#�ԈE�"����x�h1j;D��p M 64U���ؾ��鳱A.D����@��pZH��,4հ�{6�6D��A!��)L�|	�R6�~!ˇ6D���v��%����ˑ;&j��'�/D�Жb�1��T�� �,U$4JB�-D�<��%S��@� �͚C���S�,&D�\� �K�U��3R��9�"D#�@#D�pLǟ/�uH�雋G�N��BA!D�����"#8�,�d�X�T(���;D���P�l��m�o�lJ<� �:D�`f������r@�>��t$:D�d���2:��Q���5S���Q�7D�� ��9�F\�Ū�#��� fd7D�������\��X[ �ʤC�d%A�J7D��z��%"rRg	�:���X�$7D�������Ҥ���ڛM�%�j4D�̲G�\�j�(M�!k^�yܒ��0D�4�׉�x\�b�
�<77���O!D�� �<��M�/��R ��P
,y�5"O��Ӫ�k��"�o �xJ�"O�8�A�~M�N�<��S�"O� ��
)	�n�1�'��\{�P�"Ojh�WN[�'2pPk�%�Nv��hc�'�P���Iܟ��I���ӟ\��7^5Ҭ�s+7R�b�����XX�	៼�Iٟ`�	՟T�I����Iٟ ��5p����댾Wp�XtÎ 1NZ]��͟ �Iϟ�I���	�4�	��ɉH��	��dR����.�zưq�I����ʟ������ʟ��	ݟ���"�#��=Kд�uDj+���I��X�I����ܟ�������ןh�I�Q9�!�S��rv�uA&,A�_y�������䟠���	Ɵ`��ޟ���E��{��F(1Z�d�UAH2�\��Iɟ0�	����<�	����<�I�?I�pd$]T&UZ��w����Iԟ��I������T����������I��LA͎<k�	���G�ԝ�����Iß��Iȟ8�Iݟ ������I �h���_�0H�CD4r�f��IҟX�I���ٟd�	�8�I�T��	Nm�T�fb)A�Q{1�\�H>1�	�,������	ş4�I���I՟��	�{6�4�cF���l�Q��O�a�,`����|�	�X��ӟ �Iڟ��	���ɰ}�^US�%�n�`]� ;�D��꟨�	۟�����6�i��jh�X��O�7�[���� ��f"�5 �'E�Z�b>�\��6�N84���JVC�@�Xa�5F�$n��u~Dd����s�L��4B���!_8.FTz��I�!Ռ} ҽi�biۄn��=A�O:}��D��R��H?i
��Aq$� S�*���x�6�͟Д'S�>́ .�0Q�4��F��gw�L�g��M�'j�G���Oר7=�hAP�
f��q��_:J8r@s��NԦQJ�4�y�^�b>��GG�'i����6�i�@S��"��tg�0D���	)�*U��.M8L&�G{�O��+U��6��@,�q�d���yrZ�4$�h��4.�p�<I�D�a�,��lG^�>�8�E"��'#��֩y�R�	c}�%�	(�L#���%�lؕ%
*��dJ!^DaY�_�|�1��I	U��T�����7 [�HW�$?1���6�ۖu�����O?�I�[ڰC���H����Z$�	4�M{	JC~R+gӢ���&<xt�Zծ��z��i�uJ�� ��	�M�G�iO���M3����O��:��P�X�:�I�#��`��A�T.���0e��٭-P��=ͧ��$3�	���n�A�bʻI�&��#�.?����MAb�u���O�d��gA8 ,.P�qo�/d��K���>ag�i7D7�`��&>Q�Sȟ@;�`ڃ.Ԏl��MU�y�N��vK�����Rȸ>�t���|�����jƴ�'�G��p�`-�?�=(��@0s�@�{����<qL>�%�iֲś�'��I�N�my���&�� W;����',H6/�i>牔�M��i�2�J+�P��㓄e��f�J�
L�/#*�	�~l�#f���}]N�Q�B�?������0�j�͛�˂�[lX�C�3�P�#��b����Uy�_�"~uDW>���1��2i�h�jT�,'���$��D���e�	dyRl�A9���vd��i����R�K��ī>�i0*7��O��(��]gR��å"�ޭ��hX?u�<�AV��(�-��U�O�v��	S�L�|�'�*��|R,Ot�Dצ?a��C 	��e���2�&�!'(�D8��E�)��,�	D�T�A|���0��!��3`Mɒ��d�J}bai�j5lZ�<AI|��'(���A��'Dm�����W㦝���M ��[4b�F~��O�T`Ԩ�(��'���������۷�ҭ ;:ܓ��'g��'���OD�I"�M�U�<����+Y�L+��J��'��7�=�����
צ��5�@�|о%��_�/*�e�"��
�M㡿i�"U�克
���>H��p�M=���bE�=X�-�<~�P����B�x���<����D%�']^�QGٓ]���#���).��}:�is�lZ�y��	զ�>4@4;p�Z>b��q3��+  ��ٴ�6O���|����?�3cٴU@D�|�8�B�G�%�@��h	 bl�!}ё�OU2s�4 (��4�����33Y���(=C�"�{�-�r!��<�L>Q��i��]S�y"�:TZS�0DobQhF
��OH��'�86���������H6�VMҢ.��J{�ɡA�j[��O�ɩA'�N��� �����S"3��U�QM�џ2֬ӕSZ�yiS��n�����ay�U���)��<1���XE�����@�F�v�<a��iG�� �O�lZ�%��S?H
�xhѩB5l����7�B�h���7�M��i�	�8$)��'2 ި�e*��Җ<��!h����=��Y��893�i>�'�O2�TP�ϔ�g.#�n���n~�%k��p3��,�S)<�X��ϛ &r�s��:H6���O�lZ��M�'�O����'�|�1�oZ?)��3��B�RqHĲq'�:9����O������C~D�W%��<	t��/�^��d��'ВpP�	 �?q���?���?9�A���d��i�ĦE�?�ò��4/���RW�ޛZD��T����ڴ�?q+O�i�W}��hӢ�n���M���EW�@�PCׯw?�����\`���<���E�][5�WT�
�+On�)J�� j�����(d@����*��R2O��D�<I*O?��P�X ����ц!�J�C�!�ɉ�M��C~r"c�L�O+G%z>`8U��k��\��\ �y�W�\��48q���'�d|���^��yb�'QX�yRퟞ ���:�J�@�0!�$Y�y�����菸Sў�qy��''إ[T�XB�F��ì���쀟'��'�j6�;\�1O����"�y·;M����(&_,�hR ���X�OlmnZ��M[�'ɉO��g	�}��P�W
(����ۭ0G��RPĐ�!v��'�v�i��A��`��+E���i���*��&CJ�r#jPy�'��)�3?�3�i�VdZ�B�iA҅��Ђ&��"�i�����¦q�	g�i>�	�M�uO��Q)C� h|th �L/����'�d�)VƏ��yB�'���3Ӂ�/|�����O���h-[v��k�(T[�r�1��Op��h��]�3d���<l�Ѩ�R��u8Pa[֦��:���?)%?����c!�^� �6x��ɗg�ة��xE�mZ��M#�'	�i>���ӟt���˘��	�(��"n�fy�K����
���&2Ax�96g�7��G{�O�b� �q(��*�B�i�%���y�R�$$�P@ڴL9�,�<х��hq���U�2�������?�N>�&\�D��4<ě�0O��(X���b��^V@��A[2
:�XΓ�?QdЛ3^��+�#�E~�O�؉4
�Pb���F�r­^|r0����]�<��'�B�'��Sܟ������iJܸz�D��<��v%Bȟ��4��ϓ�?!��iɧ��w�sv�F�L7�y��-�1��'��6�Ϧ���43������<��4w߶P2�"�	@�Yr�).{<���	��D.���+�ў���^y������4.��Q�ђP�(`B������U���5�	y�'X�����N�L)JE�E�2]�CU�t�ܴ4��f1O��8���OA!���H�l[��F���U�#Ir~�߸c�P�&+�dX�'`�ɆS���*&
Kf��rƌ2ZL�I퟼������i>ݗ'� 7MN6"���W��㲉��Y�q剐S��
ئ��?��^�X���ʣ��X�4m'�uC�	<
�8˴�S�d��	W�@�0"����?���] Z"�rdB		��������1�aq�J��(��L�7���<p����?���?����?��?�O~Za���)��!R5�ԛW��P)f!mӨ7M�OL�S�Чk�l���H&��2ȰLX�����J�da�}����M�Y����M��'he�9�����<�޴|9���@%�g_,�2�ء#Zܴ���:@�FI���>3��'��I�L�IƟ��I�3$���_B�閫��4��@(�4Q֛W��:�4 f6\�'�?9�����)I0QX��K	\5���^-d�<���?�qS� �ݴ	 ��e�O�O�� ��4�L|�p�Q x �Fd�5r���+�3�E�P���S�M,<<k�R^�_�ּ[��:V�(��C�e�p=�'�R^�b>�9�6 O��>�2ćÁFBd�)��M�T2�@8�O�n�ҟ�$��s����4;�B{�-�94e���6Z8 |H*��i	�+@(
�A�'��[2t��ЭX�����,v��R�"�	RV2ܪJ�%��<���?i���?I����4�*TQ�D�;���p*[
T���Ʀ=�IG���`�	p̧�~�I䟠�iޡr��^b�����el�A`���M�D�i�p7�r}�O����OZ�;GH��y��dt̐��e23�yj��ä�?I���E�b�RR#��fў�IƟ��Bʉc`����5_��9DO���'��'�6-֯,21O�DS��H�6܂�+�b�!m���"��/�I����ۦ(�4�yR���gtY�P!�4:>��S&j�0�	r�� :�\=94����7K�yt���4D��@����p�~���P���C�6�e�eo*y`۶aP�d�<���l�{&��4��H�䈮i9đ� ��K1�h�"H��`�8:����qU ��>�\�@獤}�1����gixK�M��66��'W<=E>A���ԯ2[V����G<Wsg;d� -����1oR�a3$R6)mn�����%��bu�5�Y9�j��)��1q�Y-�v5�B��Z�$�1t+�4'���	ҟ<%�֘�.'L�svh�3D���O��@��7��O�Y���O���Ov�d�O����O2�dѻ,�D��B�B7R�|����8@�6�҆I�y�	۟���r�I۟���!j��Hچ�ۏg���E$!7`�a���埤�I�����ҟ��	ʟ��I���z�O	�E��R�6��#
�,)�C�Ol���O>�On���O�q����H����j��-j4.��G�<gHun��L�I͟`�I��ɘ~Wr�CK|�j9Gn���b�1�������!]����'p�'���'#���Ok�i���)H=�au���R/�M�2��-Bh�DW�m`�@��E��H�F3|ZL�8F��~ql9H��-�#�F��"5�Qс/@&㠝�T���Q�^(<�[@����']:%Z~�H�1J�M8D�=xnʝ+��U�@��Իc�؃M���#'$ٲ4~4u�eM�%b���ç_%�H,��I�6y́�S��.�cB�Q�̸2�G�1�"0�?(��|�uL� UM|�*���$>BY[vY,}G�!��U*{ʁ����Sr4���x)�Mcq`�7h�� +0gܱ�?I��?��\�Ώ�f̮h�w���T���k
'p�$�]e��bWc�/.���R���O�p@����<�G���e�]�Eى_M��0aaT�hW��su��sqDII���F��}R�I��.�	='���.ռy�x�S�%I�PM���H>i�%I���>�O$�Pr���A��0�F⍟C6u�"O� ��r�KŞwNɰV���
S����9OX�Ks����|""E������� �)�R�ڵ:�k���r�'���'��]��4�	�|R%l�e�@=S�g��b!`�/&|;����(v\6#�G��e����T��e� �<i��4TU�҃��JQ���6'i�!R�����r��>moP�Zq��Z�<Q�E�}_4a���(w��티��?����	�?a�� ;2��9� A-aA�!E"�T�<y�i]�wS�)(�$�"�|y��z̓hs��|ҨIq��6��O(��%�@D�F	�	?��`�IO���OhI!�(�O���m>Y��%��ua�y��3q�ӥz��qR��^s�Y�M� ����T�P+Q��r�iS� X!�X��U�.TZx�U��)��)��m�&mY�5�cέm{Q����'�O� '�D�����}H���l
jm�Bh(D�$�#
��iѰ�95'��.)�"%��ܴC��@B?l5��� g�%���3L>AĪ�-����'!B\>��$B_�8�@'
 ��P`* _������� �	�uΚQ �燶=rΕ�S!��3�h�I��02��O�PE��p�D�8Ҭ��N��WR8n�8�푌Z~T�q�Q�|�� K?I(��		f$��a3j՚O���ps�$}��Ԫ�?��|��ThG�8��-��`A� �r
���y�͜�I%�8��ɞ�i��X�' �0<�6�Ɉ�� �@�%��#'jJ* ���ٴ�?Y���?9���S���a���?a���?�;p�����A� U��*���m�h�	F�F����z�'� ���mK����^�^qW�/C�܅�IŮ`����L[/I1NuC�'ҊPS)�v�g�	/=�Lm���7�`�	�R��1`ڴu��	�Lp��4���i:���o�  �Y��)F	ϊa�٢"O�x{�H,k���8 ��KAP �撟����D�o}RT�(C�'A�K�8)T��/Mvp�7F�)%�|�
�џ\�������(�u��'�r8�p#��O���򕈑�pR��0����`���B�o��M��'2�P����Y	(B�I��!�N:J�a��$�:�6�p
ӓ&�0��7��G�թ�kE�Z[<�"a����r�82��@�j��8�]&����l�F�ȇ�B&�-�@��[��<9��ě�fC��n����5#�|3��R� 06�i�/ 2B e���)��ߟ�I�|n%\ v	~�(�L*p@�y����z{ @�@B��6+d���9��p�T!�;K(�<�A�;H$�If�4�"ׇ ,vP�Dr��	�F����י<��@
��?g'�<yV�\�޴Mq�� BĎ��d@W�f�Ph�	��������	J�S�O�Ԡ��&�!c�)Y���$V��3���>��|bP�i<-�%�<����d�^^)�Q�'^�ɶFVtA8�4�?����I��B"�OJ�H��շo�Irbq@��O��D\���ҧ[N�09Шլog(�yah�	,~`�'_QZ����F{a�a�3�pе�OlR�eA�2R*hj5�ư$��7��G�.9e�?}��c�
1����MĜF���:`�8}⩛�?W�iǶ6��O@�?�	fOE�z�,�v��gy�C$�7�	ş���I,
d�S��p�~��ԍK�&�V�F{�O�"=�TE*G��a0�YiY(��%�	�RT�F�'���' ��s (V�2�'��'�g�AL��@x�ιs"=�4 Z�V�4�g���mY8��D��Ip�)u�)�yg�IX�'r�CPC^�5��]��,�B��&e٧6X.]�lt��:p�aӸ�>�C�n�v���ޗ|�l	cO�-��P"�,�e��x%�L���Oq��'LD�Z�U�F�i�6�A�7,�I��'��z��>Ϙ��8jt�\����O`�Fz�� djJ���J�6�d��G�X��q���)G�����O����Ov��;�?���t��{)��i6K'+h���Ӈ�Eؾ��d
�R�zē	� 2�0Q�N#r?�uYa��4a�� ���!�N�k��RN�9t�D<F,�
�K�2��`ɗ�O�k�x���O�Ol���OD�Xc�C��aͫ�@(N���Ys�-�y�¢���B�A B���[A-��'rD꓌�:����'q�!۞g�`�&�$X�q�s�	 Kb�'.-aB�'J�2���3��	6:����W�gr��^��ShѾ�Jb B�y�p�F��'�Q�0kR+R-�`K��@����EG�����B/lJ��[�\hN ���M.H���B4[K�m|Ӽ��'@�s��l�-�U鎿|L��+�y2�'A�y�X�f�� 1d��D/�A2��'�O,�=�'c?�V�G	��@ˣ�
>������utR\�Iw!ڋ�M���?Y/�9b���OԼ�� ؞fTPB�G�1+©���OB��´#L��X.G�
��b��S!��3��ƫ;E��'d����ɫ9������^���O�K�OruZ��S�O
L��dB[VaĔ�'0��i��p�8��O޾�|\cw �c�Ğ�}� ���A?���j��ZQ�&��>tV!�R`�H�p�U�K�2�YZV&�=�'S푞� �yv�@�y`����S	��d�ۦ�	�x�Ii�j\�@i�H���4�i�9	����.Qz� [�A'$4f���z�:��ֱgz�E��Wڈ<�|�N<y�Bۏa5��2A�VqvUr�\I����D�{��
f۹ ��}I<GL\�e��]Bw`��R*N��EQ�)���ǰ<iA*@���?��?���+X	� �� �~���fBR�<��N�a^A�E&EZ
(�T~d3�S��Y��ee�b��c��^l�3�$ǻ[��x��������(�u�'.�<���1��	r9�xS�A%/t ��̋!�XH��ɚ�D�� �������#Z"48�(#V)�<`S)�^H�s�a^�8 ��G{�U
CvʄB/[��XE	 'j�
]��x)a��CS�J� Ͳ��h��!�y���nr�t��ҁv6H|������'ɶ7-?��G���ioZ��0�I�2�ZQ�u�� 4���h�1{=Q�	��h�f���(�	�|�W,��z���릅2 6'3P��w��,J�l���NҘ1(�0�a�H�E�qGy�-^�z�� qh�(�� �)nl-q�#ƕ`�����+�L�����&	 :��Dy��K�?)p�ih6�^��99�	хDc���5#�Eo�m̓�?������h2V�C
Kt�p����}.�Xi��T���įl�V���i'8��q3��?	L��O�O4˓2Fm� �i ��'�哬c���I+�4��0o
K������B�Pܝ�	��0���G�h�� �Cb�0-�t(�Ʉ�y�dt�e(X�$.H�;+z��-�)�b��Ҳ��?�V�ǰ_���u%�	�\� 6`m�� V�0��A)�)�<�"�#|�'Uzy*��[Eɧ�>ag꟣>_j�h�Lּy�X�;�'�����0�sd��n@L���i>�H��D�@nq����QQ2���'B�Q��n���I�x����uw��������ß�>yD��z���#eʞ��0 �RՂX�D惱=�D��5�i[�����T�����?����F�K6�D���h�
&��P���_�xT(�j{Ӕ]�O�����+gX�B&�D��C��C�(��F�i�~ʓ1ta�i>���j4� ґ�L,̈́5:@�C*q?05���F��F�h)
���(;��'��"=�O�	�h�q�b��#��,�uNP�/��ၘ��f9�I��@�����Zw���'p�)OT��Z1e֧��Z�m����o��s��c��5��pQé�a�Tk�򤈮(���8q��ɖℜ�J(U�'�^%"c^�_	�h�	Ifk(���d 	(�H�j��^��_�{������' 4����T�� Õ{o��S&$��$�a|��|bcH4�*5�rd��E�v����̘'�7"�ĕ"�o�Ɵ,�	K���aG���g ����c��@��۟XJӃ�ڟH�	�|Z�.��4R�(	��U�������+)���	�6ʴ�di�:?�d�q��]�l�<�I�/~4 7/�2\r���C�L`�鐏�zu�$�S�ؖ�<4�2�[��4�<� Iȟ`�K<�!؅���yp�L�gSz5[qZO�<a���2X�HS6%J�2 ���p�'�ў�Ӽ�MsW,�7R8�
S�8�=��ܯ��{� �i�b�'��(=�v���)�\��fN2o���� Ո^�`q��ݟd�d-�$sE���Z~*�Dʧ�9��E�,���#��٤h��إO��@.W*y�,�ɠ��"������+9�p�������'u����@ɧ�O��=;���'>�lxh���$������4N�s�����&�3%DzL��Ak����+#�!�@��ې-�FLr7AXb�1 �i�B�'��Q��`���'Q��'��w�,X��H6
��2�! �X�!�DS:��yB���p���'
#$�4��`6��']��K�^>b}����h�����\�`�所Ó|�L\��?�}&���SL�<O��!fl�'0�Q
dB$D��2D���&�
�E�>5g��Xt%.?�1�)§Pm�Y!�M
?S�H��j�1w�걙�L�c��;��?����?у��X�D�O���N^ ��eGy�b�D�H������V6(0T��+O����'.�lZ��a�剎TB,��ʚ��x���_J�Ht#�8"����\al����sV�,���	�*L����N:K�v<���=��®�O������TZ���#|U|R�]=j�����=+Xu�w�%#���%
1JZV��<�P�i��'�.�z �t�>�d�Ox���р-�p��U"1GN<����O8��@0r!����O����[td�%}+���ā$���!`� ���c�	$�:	�d� ]����M�'.R`yfj�4�豨�TMi��惚1<E���
� ��o��|Sv��P�j�'BV���S�'-�(�I�O��B�@��<Pi�'|���%���5K&��
/�,#��!��|��i���-�&y���cP��"0� �|���6�O�D�|r�ǂ��?� �dy!aŭ>_�[wi��.�A���O����.B�^���F�0J�6�x!#��*�e*d��c��'BZ�|��V��L"7��;�u�O�hR�D��z'U2���(�~���?�3��0��)q��
^��X�b0}�
��?���|�����tM��k�e����M�0A��y2(���}:�(��e5�܅1�ў��HO�(�t ɇoVNR�6��9��&�Ҧ	��ݟ8�	2gv���!l�П��	HnzމrӀ�6sY�tZ��6@������h̓cj iô�'c����
��?����G���­�aM	y�=[�W�m�0�HR��O�f�y^���d�X_@�8R�����-3������)�3����
?�  �Ǹ	p�k�/6Z!�Dܧy��H�͛�8U�����`F�I��HO�8���7��kA+�;R�E�t���aN0=	u�ݧ;� �d�O��O�����?�������قfa���E�ؙ��<R��gхPx����4#��	��FIu(�ˋ�dʢ
�*)�$N�oO`�� ��$��U��Rm��	��/b 41���*��f�ToO$��%��/G��4�厢&�l() )X6~�Bn.�OhyY�dٖt;�|��ŌJ�@�+��'`�'9t)���
=bQ�&�7"�*��y�s�h�O���k@�����9�׮I�zqqjטf�����ԟ��	?-�~���۟��'jˢa��j�\��u��t��-�R�T9� 2$˕.G��H�c����O�Y�@�зe��qru��� ���	�r���Q��R���n�BG^4J���Q9�G.�ĕ	S�,�r�gX�f�8Pʔ�wL!�$͂
$���=���S⨐>(!!����陔���VV����?��,���^�	�.�T�޴�?�����F*U ��D�jrzU��C4`�8#�EȗO� ���OXz��3BX�����\R����-W���Zc�|�I�����ʇK-#:�y��h��_l"
��%sU��7D�f���&�������
x m���jI^-�5LZ�+��qђ��I<��S�'��h����/�(vD��1A����2N)9��?A�*G�[6D?���	�HO�Y�խ;�pe� C�i͘4
�"Ѧ����@�� 5,�O����	ޟL�i����;T���{���9R�C�=`Y�eBum@�ŰeJ�k��1��D��Qs&5̓4��rqD@�k�`"�d7����0/X�,G� �ݴx��(���[�{i~�'>) E�-]��Ѿm���V(C}`I�Ť5(�R�'�T��$�Oq��'G��(0e���L#&oȌFX0�[�'l�Xw-�F���׏���O��Ez�O�'��;�l^,s��"b�poh:���o�G�'R�' 2M~�=��ßT�'m����v��Ww���� ےf~�Bg��]�rQAv�"[x^��g�&-�u�'��B�m�e���W�	�>F�T9bm���%)���J�r�bG�Z7�[��(O��:�`
�w�8�{'�W�P�0�ĊQj��#�OrHaaZ&	0R����E6v0e"O@��A��zy�Q ��8]�����dR�m'��3�@#�M���?qV�C�!&�-["$�wJp���(@��?���{6�](��?	�Oal��dcӞB>�=��M�@��dC3(�"���P�M�y�Ё��џP!ŕ� `��2S�T9x��l��)�Jju�#ʀ%W�����d�x%�g���?����q�-YR(e�f�_�:�Z##ʘ(DC�ɴ.+�@��X�!��q�T-+$�B�	�M;!�_�P�F�1��A8��iB��
��\дU�R����'��St^����|�0��&L�>;3��vbp��Iӟ Z���88[$��")�x ,b�Z>Y;�_�-�Ƹ�B�@�\7�z�K*}�9ն��n��_@1Z&�A�OҞu�t�E�I����',٤:,���L���o�Ot��(�'�?AP 	�%���)��� �!����xr�V�:�z)�5C��iΒ�&���0<�#�(>�*�J��ߦ���P':gq6��O����O���ğ�{@���O��D�O���R����ߜW����%�>#!"� T� �<}��_�jI��+��?��](L]R0O&(�B.�r�`��Y@����9��(�"	p����fo�q�BDk�,C,�y�mX�rIڱh�&�I��k���`��7�{y2�X��?ͧ�*�bH�U��mz��_!?ed�µ���y�FKb�1���<D��qu�ߙ��p�'@6��OH˓ZN�4Xt'�(:�p����A�6ețv����?!��?�d������O��ƽP�&��[Zt�	"�I
��d� f��5!���ቄB<0a��;� ��	�5#�����O��	&NJ�V�h'*���BT�� ��V���ˑA�Z퐢�	+��!�Hۛ`��Q�Bʆ9��$��K�O�����< ����&dhl��b-:C䉲b4�k2B�@�c��9�c�$�ܴ��"�*�� �i;"�'�L�(��<�8�{pfCB����'�b��l��'_��W�
r�i"�`G�rfZ(�� z4��_�Dt
��1!��&���2f�'��a���KJ3t��'�:�#A���,�ѵ�Q
\,���+O�%6"?q'	���zH<� �Z�4���Ë�w�ʐx(LG�<�2�ޘxJT��bb >�T�p��A<źi��)��`Kb����h�3.���	�y�F�-��듕?�)��	
Q��Of�KJ�sX�XіiY�,����Od��L�\� ����B�_H�����O�S^�TIM*�tyxQ��"pW D{G@B��It�p���l�
e�`��S ���3��M\���S�\�ur��'�
83����D!ҧ�rw/��P��a*�P��!�@S���xb��=|I~	��'[�z0 cԦ�0<��I�d?J��GO�R�.a�UHކ@� ���4�?A��?y4a��.ʄP���?����?)���BZ ���D����M�Bdڇi��{��+�p�� >��Yy� $��M	�h� $6Ot�!RA� NP�y���'�� �B����
��H�U��H�R`�e.q���PS�J)�y'E$J���s��N�@�x���D.P6Ӧa�ɸP5޴�)�<��eH�Z6K_C�\8�uD��|��d:��:����/�M�"���nL6v���Γ�?�Աi�7�=����v����<��8̼��wh� u�J���a�^��ƨ��?����?�����O��d|>�S҈�#�#񃚷	21�n�S�8!̅ +Rv�� cf���AFŹ&�Q��B�,W�n��K��q�-��8#�Ʌ��5�v ��Ɗ@*�1`��f1p�Ey"CW�6T���|o�IPR�ǖ&7.D��9/�V�-�d�O���>�I�E?��I%j��p�B�z)]�/����4�$�#[� l8��hR�PIz1OBo��(�'O����x��D�ON*`�x���aE!L"R�Bp ��O��H {��d�O��S�O�F�dg�6��(%�=�s=O hMb�]y@�����*Q�a�G��(O4M"��	J`B5*�%�:<�S��\:F�AN�>d��pk1��;YZ���D��(O�ha�'��O*%���^�+�FɑW�đU�:9�"OZ�
�@� ^Ă�$ۅ3��6%4�hO�I
Ҧ�V��x�*�9��G�5tx���!�Q�I�	�f��ݴ�?!����ӱ �����1.�Q;4Bݿy$���)�Us~���O��ℤѼ��e+VA��A���
#M��t��`|�aG�m�Ԅ)T�����QG����ɮe�!���ԉ<<�$YA�i�U�T�=d�Ӑg��u'�_�s��9�MO�`7.����&0�����@�)���W
9�� ۶}<���̣fe6C�,o������2\���;&i�!�"�F{�O	�#=It�ܺQW�{P��>-Q�٤O	�K���'4b�'=��Sc�w�R�':��ygPI&t���	��{�
�p1D�5�@E�w�Z�б��D�SEXs�I�!'��)�'�ֱ���B�&�n�*��$_-|��j�[����놳Dn�T���N�>	�n�|��OZ_K���>��i��#�S�ɳ�kͦi����K>��k���>�O>ؚ��>J�:�B�"u1а�"O:=z"mM"�Z�ct��6��8�?O��D
@���D�|⥜=�h�إKY����i��؟+� %B� Ț_�"�'4R�'�j����	�|�f�Ⱥǎ�3snOj���I2��s�F�Cr�Y��< ��k���Jȣ�B�<1s��+عY�GS:0*���F�8]�n9'�0�{T 	!G���S�Aƥe.�(Fy����k��噠�\�EH,õ�Y$1�4��$ha
���ǃ-L
U�s]��0>QJ>1�	ϜK�$	Q�ǉZ��"Dbh�%��V�|B�U'T�7��O�����0x���3Pw��Fa._��$�OR��7��OR��m>-V��.Gs��O�y�1݀0tx�G�r|�v�'D�p���ʕlnJ�Y2�Ԁw��L��?>"�HP�ǗB��l�$� ZX���퉒J ��h�ɤ<>�}��A� kx����M�C�	�asD	� � �l�	���AA*B��.�M��U*�`	bc%��|pni�6lت��v���B&�i��''�S�^��	g.t�� �+W���s�̙�o����ǟ��&'�^�Z5�SFA�x��O�e�6-: 
�q�Df�?@��TZ�需uz��Ѓ���ɪ6�:<�'	�����t/y��%Z۴7h�TA���u�j�.+�ְs�
R���q�d� ��$^���ȦA޴�?��$���^08\�5!ߢx�,�@�ј'�b�'�20�`�(L�
)���*�Z���i>%Ҋ��Ա3-!��{�^H�- '8�J����O���O:p��ꁡ),���O����Ov��E[޹ya���_&�̱SfH6v*��%�PІDǁZ������)ŘO5X�'=�x��K8L} �@�
�?G��K%��/Y�jPr�����ӗJF�ĸOh"�'�p���8~��젓�E�L�h�s�'��
	�\�4���=��jQ�n7>�ՇD��!3�^�<����!]�pY;vH�7�:a��ʁV~�/��|r���$��f�Z<��ʳ'H:��K,bMx#aꑞ&,����O����Of8�;�?9�����i��-ގ���	H�6�����k��L�	�'�Pd� rA���}�p�2/�lL��Ӕ�+�;A�=7�̌Q�K��t��H�G�Hۦ��X؟4���=؂��ʂ*"����ŏ3D�$��������$ӾO�@���%�	��'k���!l�6���OR��jс&[��16�ЍM3��cT��O6��H N7��O��7@���wVZhbT��*՚�WC�S{�i�HA~^�n�"G4��BV�ɽSy`i��N�.����,�;rA:��s��C�h�-�ZE ��Cn�6fj�AW��v�`�d�a�	�sm��#��=%�tűHTR�hB�{�Lܰ�c�9�T�a�2X,"<���4��%lډ��\!V�K6~�m�u�uz�$�|!a��Mc���?A)��}��OHpd$��Z&�����[������O���ٚKpv��c��+k��qdf��oSv%��g<~�˧M'�<�0�ؑ^z�I�lκO\U�O�H����B7:�����4N��I���ʟ�ЂEBR^�XprG�ZW�f���>٤���PxO>��Z(x�c����L=*DΆA�<����DL	Pt�_�lN��4��hO���l�'ŲX��c�N��Hׂ���l��k�l��O��$�.S.����?����?��Ӽ��da<�@[�o0V�~������9%
�l�����G��\���T	
�+���ϓ7�,��S�܅I����ԅt���zbi 
��b"�YJQߴظOo��i���<����?ʰah1	�L�.��D����'�&���S�g�/ 
N�ʓ�N�	�j�4��6�ZB�I0U,h 'Y$9�vȂVN�WWV�	矸i��4�f�O�hb�����\�iV?A� i��"O�*��\�xa��>%��s�"O���M�-͖q
ci��'|\�"O"�8�F�!�@
E.�6rxZM�V"O�4)���)=Jr�`7xn��6"OT��J](N� h�G��J�bS"O\��UdJ7KQ�M��M
5��ճd"O ��#�[x6���u#%p�	.�y�+�TBx0Y�k���e�1�y���j2N3a*Ɇ!þ�B�L��y�K�hm22�̘���㧘)�yR�ă>t� 1���9~�{�Eƺ�y�-z<*I{��D��|�1C�܆�ybH;z�����~�:	*c���y�N\7���H%oc,�ae����y�f��=�l@ ��9�^=�����y�#�_(���fg����ZU���y2HȆ[d�M���YNxq�U�O�<���&,��bmIL0f1�Ǣ�r�<�'*��Cvt�K�o�XK2�����q�<)�K>TG��s���x�R�s�<��#U�U�D�s��a��h FoLl�<����RSL��fkM�iAT���"�d�<�
	V_�Y���j���wH	_�<	���O'�s��6m>��0/�\�<�$)ͻ*u�}����M�8�`��D^�<Ѧ�O�A���x�.l���Z�\Z�<iU�M�R�H�C�^!s���0*�B�Ɇ f -�#*R:Z*5��H�^2�B�	�X�1A@�?l���`�5�B�	
=<�A�$ײVw�l3�Pi�C�I�7�X�I%B�	.�wnϜl٢C�	4&lP�"h\�	���;�G��%lNB䉃��Q�-L����4FI��C�?~��8c��a�r��F�\uC�I<&Y����:_f�2d��Q�B�	�,��@����o�*����8��C�ɮ|�T�rBJZ��BUɳ��C�I6KT�0���*F~>a�%�/I�C�ɩ ,D��J?c�6�I�I>^!�C䉣OtڥB�4=$&ݓ����C�ɜo��xg� �:��7.O��B�ɇb���곊^�wl���(�	���ߍ~+�{�.�j�y�d�ܧ"�S�지 �)��WRc
�2b��=�VQP�=OzD"1��
c���c%e\�(���I�9h�͘��	:�&y��cA��5��Nˬ��^���=��|�>[zqص�]�V��'c��1j ᱱ���p<�W���}��.�?*XL���]�Yr���n��A�b�����y�S�Of|��'ag&��

3>���#F��qDz���snpJ��9_�xp�������1�.��$��&F��%��H~���	WX�OF�ksџ��ˇ�G� ����������T0j�L�9?���oڷCx0��(�*-��8�O86��O�Y�Q�BA�Rx0I�ǑTz�H ʪ���g�Y�|!��#W"֎�K�(8ړ�\L[�"��KtFzp����M�4�Ք%��'sL�{yBo�G7��X�5���sҨȫ�e^  /z����H��M�rF
59����=5�blbe�Ɯ�RR�I�'8��f�w�.�,��'�"=ͧ����
��#l�"�B��f�Ӈ! �L�R��˕(vLX�GQ�G����'u��r.��"� �(Sɛ�3���z���O��v&��b' �*W���s��xT�'�d�S�,�U| 	W��ڲ�;ݴ>Ꞅ ���/`aJ��rKK�0'(�D~hV�����B�$.�l}i%kM�<�f��X�I�tM���Ʒ2���`V,Fў�Pg�#�l��ǂ�(#[2I��K>K�f<����k��dB�x�`���Y>5�P����1����'y�@�3��Ǌ��%����-ӂdsz@���d1��|���a~X��BҔ#JE�ȧ�����-�6���C%aڱN%"��R��(
k�i�'Vdɓ�}����C��-�4Z�	iP��C��j��D�Od�%���fE��%�;3�>�Ѥ'	$K���,q���nso>�Ӡ/&����a2���`�0��<����Ǟ��e����Ľ��_�r�i���	���M���3�p�=������`�_H�HC��� wgXP[,�Q�=y�A�~��O��xAPp���#Q "�
��.��ى�4.��y �'�pp���^�`��m�S �&Z�J���F5=΄����O�M�5�������M�D��M�
Ay��
� wB%hcΚ%/(�*�nZ^�'S�=�P�N�{!�3c��WdS�O��D��X�)xo�0[��e��'$%��#�F�I֟��@��"D��:�g�P�d�%�O^��1����4Yt��@Z`��i�FTK�f��@�X+Lڢ���{��$i����@��5Yq�ɍc���Ăg���I�U���:�I�y�,��t�� 5��=!1+�&�� b3��s$R�8�@FR3�(cf�ɨ�y2��P3�"B�gn���6�
p���IS�"�z�nZ8���l��L�X7K��٩䩊b.ڽ�ЯZ
Y��x�h]�	Q��'{�,LزnS�]�eHC���x�.�-�HOn�Z��_�n��0����IJ�q�S�Xa�#xv@����SI4B�8O�1��h����	⟈2�'оp��D�@((a�'��YvdU�K֍��S"3,L�	�%�V��lͨ]�8$0ǊѴ6��#?��'\$k�Ā�E��L�e�э�M��E���h��K�\�,��'L�hO(��U��%�p�s�P�L؂y*b����FR�d�*~̝�S�\�2�IB�"'�f��3�̹~���E4�e����L��M<8+L�2�Ζ1_��{���(��M�t���1��X�opf���n�"m.�� !��Y�'n�Bf��x�Z\P�B�W�l��O@�:ወ�zj�P��AK�U@������ʦ��	�S>�9����:��7X<!���ɪ1O`)Is��Lp��Ɣ�^��6�e���ޞ"�����H�㑟��=�L���jx�$��%�] ��ώ�V�\��	_��u�c��*F{�垫gw� D$�,E�T���E��xro.��8@�#W��r��n�h�SQ�KoY�a���C(	�F7�4�
|�Ǔo�BH�0���e�(,r�2��e��H�D��� )��J�t ��P�ErD9Q���Q;��ɡN� e
g��y"�*�/w��\Z��C%i��=��K��-�F}���9��P�R`�#):d٦��?	���$aKN	���".��P�+
�� d�	a�vA�Mġ]
~Dj!�!~�Ї$[�Q���� ��#�:P�dY*���OD�N�щ��P?L�E{�'#^H�P�f�X�w!�!d���*H����?�c�L�!��a�DgL���Ŝ}�̅���)Ѱ<�FA��y�D����k�=($��^XI����J
_������z*�� aʞ$�څ0�\�<!qM�6�~=�!��m2�UȦ�y���C;-?���g�V��ĚF�ob9ؕN��o�a����O$@*�.��i������z|Ę�	�͠=��@�����7+����Y� U�E�_.�p���	�GM�">1�kJ�-����	N
$]@e��,S>��6�'�.�J�H֪{Nl�[elC.X,QF炊4d����'9`�"dLi�1��1{Rv�i�nB�>6��B�)�O�QxƠL���;dn�h�4H	�\�.���䟏��03K�6���x���I/-�	�a �6#���(׉I�1�J�>і��Y�@l1@�2�ug�Tϟ��A����Ȍ�8h-�U�n��A�$ 9y ���4�ܛ��,D�(�[%���T@
���
C����
I|$� V�������d3�¢=� ���1�7(Ь���d�]_4�0��YC>y��	?i�8u�V�����D[�J���a�N١Wj���3-m*$I�w���Qu�ƖnՐ�c�$T�,/Hi�GҚ�HOF��â�ث1"*���N1K�x"=�ɂ`SG��8QH�R#��E}#K�4�����Y�{�N��.I���	�w��n��Ȗ,��*$�9�	� x��S쟠��͔?W��Г k�6m�t<(�ofӶ���b<:�d�Ӣ僮GE��Bu�	V}��:"OO05FM���>5uT�a�oK�cr��Uk�ԟ�QWO�?�D{ҊͰh����4zŠiJE,�`-����?��+R�ҧ��oo�(�q���Be�l����|����?�p<��)��
���7�Hd��`Ԩo˰�6�C�~K�k^T�ȺQ�j 	���
8$DSD"X^�'A���Pl͈���Rqf<R"�( �O��V&*�n��$BJ+��P �I�(�R�@��;.�"e��*(Er���&Eb88!,Q2�`��
�/|\��@'��$�DN"�Z���-��O2Ic�(h��-h�Z	X0:-��V��E"��D#+��� ����hOxM�r��"{��x�#��z�,E�r�i�N�Z�{r��T��(���#@ R�/�0�M���9UѠ�3Pe}����zdTD�;I �@q�|bxđ ��^�D�	.Tǀ@�%�OL~�Y�����)������%z@J�!��3"�ڨ��D�7�B��u�`%���	1���+O2��Ԧ��=Kd� `-��?��O��C�R0�y�S�Yڕ�o���,���D�?	B&]:d�#� S�z}��˦�I���=$e���S�O� �r�<��(h��"�"E�4}�e15�K�pmz����)g<,5K��5
ӮW.op��p��B�T��dG{�jʤm� ���I;+�8�A+*�M��"�5��l�eȧ��O��iӆ��*RԆ�{%���E宸Z6��-xz� A�'B���biޅ���@U��+Æ�#0����O�	V�Ю,x8'�b?�v+�n8
�sHϤ]d��b�$J���v鉖���;�o�r}\0`��.e���4�~!"�B�
eҼ��F�w, �'W
U)���fv���g		?�s�@���kb/��?��I(z�8c�-�rH�wn�#B�6M_4'L@!P�mM.i}�ly@ L���'=NlxBD�0�tEڄ����\�P�­thH;4��m���ۑ��AE(�H��S`h����hO<-8���@�&�#���b:R�S`�âS��@&��Rb�˲s�N@�m
,q���Y��͌�<������W:`=�6�5=_̉���Y8��� �(�y�
��Aϐ�k�.��/?͹ #W�H�Щ���F���H�"|�Q$B*��D�N�B`H8W"�-[����҉>ғt`}�f/Fp���)Ά��y�'�⸋0�*j�}b�d�BF��?OX�C���7v6�*f��1�⹉4�d�X|a�h�"�L��'J2u�lKd[�9Q��]h��@ߴN�l��d�g괸�%Ph�e$���!p(e��
�_ �]b6(Q�.݌�D��Zu(��d�&�������Q��?�F�=��&��@�F-�(�EF`@'M�Z��	��|"E���K"#��q��$��n9�����u)�g�>�P8H��('������L�r����$A> ��ͻS��,¦�G�N��	�7H�h8���,���1��� ��|�S�O��i:�'^���#�h|���ff�j �XFzR΂*o���	_~�~H1�a��N�kE~��'���@|v�qgM�"=��i���o�+KJ����ϕb?�)�=�\XP�D�7�?Q%��?E@)!5�,t(��(�=a�e$&��J�.E]��B&�ԟb P#��hS�`U�=�Ihq(�RY�q�4Af� �ȶϓI��"S"&�"6�	5^���`���x�ň\��Q�a�I*��A�֝��$�`��)<VY�p݄m�!a`��^N���i��K����$�&u���]'G/t��A��1�i�jK�up�JG�]��<1�2?E�ċ�2��t떯-ˊ`t�Ӭ+�MB4�[�y�*֏Q�:����$8�x3���y�*D�<BF�E��"}�Y���4�y� =o{�xJ�gX�cb��g��yr��/(��6Q]%d�cbA��y�C�O�hU�ef�XՎ���Jρ�y��(`�
!��Ǐe�0�w�H��ynR�Wl�W�F=5��E���@
�y�Ȼc�v%h�ƅ�1���w���yR�ν�@�g!ǐ�
�'H��y�Q4%�J�!2?NvUd�
��y��L�A��*�U4nB��03`��y�� &>a�O\<^�FP�Ǿ�y\��;��ݼ\D�#3�E0�y�D� ,�Ȕ[ώ&H��C��y"���h�q$W4R����	 �y�ꗅ�|�!�7I7TðH��y2P�n�R1hѽ�ֈ�k���y��$D� �,ߦq�.\���K$�y
� x���.�>1ġQ�S�u��b�"O��������wjB��V�	�"O��P4�U0Q��(�B�rt��"O��
!�Ͼsb-AR��_�i7"O�Hڤ��;E��U eF�%�V"O$�8��ƇC��q`A-��_-
��"Ovu���A	x���Ǝg60�#�"O!�bjر:���J$/��E�bj�"On	ĂK�F5��Ed�xn|a��"O�kw�G!b�=&��<Yj�P�"O�%Σ�]���ѶI��KS>�ȓB�`�#�@����D<S���'�r�
��͇>%yZqX�{��ȓ(À,����(a:�c��O=s6�T�����%!�4)�q��,ͫ����"O�xh$��:H�>ͺ����d��"OHq���M��!F�u��@"O�9{�E2���`O����r"O���p&C��8�S��4&�����"O�4��ڂh� Q���Ҽ/��ź'"O�AIe-�1f�:!�i��<�b"O�)��2~�$�2�N'+��MIg"O����ļ*.T�`�FnKp8�s"O,rP@J�k��Ѓ��S�dA����"O�x���:ka�����a?l��"O��Yd@$i]�0�eY5<)"Ob�ʄ�=7�堥b� |3�"O��Z�aޣ>���IV�S����"OQ����{w�mh��'Wa~=�a"O~�:��.r|4x�j4x/��e"Od 3s��}"L訡J�;2��7"O��& L8���F� X9�"Oz����2-"�=��U�9� ܉�"O�ѢWo^�<�����P�{�"O<��J�|���
Nٕ_�De3"O��K���9�V-p�⃆]�p� �"O�U�Ҧ�O��Ȩ� `Ȅ���"OPR�ތP�����ݴ���C"O(5�Q6Jm*�ZE��q	"�a"O� r��ϴ466m�3���fy�"O ���t��0i##�%w�Z%:�"Op�v@S�L$�t�Իu�h���"O�IQI��~SŸfB9a�`�X'"O��xw�K"HZ�y"/}���"O�x��G�B�H�a�Y�3uJ��"Of�)�@+[2%�	�R��i1�"O��j5a�"m5t|� ��<8�`Yz�"O8��B�Ƙp�{��
���"O��X�%>#!��nP
pk``��"O�pq���2n�Z�!�U.aY:a�v"O.��b��� t9s�	C�T�s"OT�q�e�@�D(����U6pA�"Ot`ڃ�I���|��J6E��!!"O@PAt�- Yj��@A2B��EJ�"O`�0b���g�����O���*0Ё"O|Q����m)�����-�^�ٳ"O��e�B�,�������1X���"O�RqN�~ӜD���$^���D"O�Ș��i�^��bIP K�}K�"O�1%�O�#9���&�ڭ{�ʥ�7"O���l�Ol��(��j��"Ompg%��y��I��G�1�d�� "OH����~ƺ��"mױ'�$���"O4�B5�XJ .�V��%���"O� �]�a��q�~��5@�az#�"O�=�7h�� /z�!�����"O@���)�y�F��$��L��@�"O�,�C��֬)d�J�Jt}��"Oܐۖc�L��swo]u�L�:�"O
�
0��O*�Ю��H��S'"O\��Ι6h d�ЍU*��!cA�'~�$[*y� ��+<�ִ��h�1�!�/ݢA�g�3Q��-����hy�����B �D�Z2��m�s~!�dܾ @�����PO+���J(YKQ��G��&i" pis��\и`m���y��j�AP�S�A�2�b�$�~��)ڧ <Ht�� ��fS:]�@�6���ȓ~6B��A�L�I��= �d�.~-
]Dz��'`N�jf��쩣��TZ(��X��y��'�f<�a
1g4t3I�R[��	�'���a�(_/+��I`ci߃H6�C
�'X�]�e1"��#�LS.?ʢ�S���hO?e@5�3I�R3�� �x�R�G�K�<y�(QLo�����Q�+ዕO!�$L���%�ԇ	/nm�(Y�G5!�d!��LȄˋ+@~r�z6h��B+!�Ԉe�T��M�5�9�f��!�$:$�6�����i��南W�!�dԁ�8����J�(��`��+�!��-��"�թ#z8if��!򤊒tr�U�U�Ѩq@��&�D�[!��B.1#䅱����H0"M��a}!��Ok�t;�*L0/��Mz��Oe!�ڮK��ق��ۯ9��au��:5!�[0ik:���c���P�ʁ/-!�Ȭ�<#�F����2�N7
!�d֋/�4{SI���U���Q�U!�D�O�eS���1gg���L�kb��"O�}q��Ll��`&Y$� K�"OHMR�9�@@��Xdh0��'��' A�&�\L9����GE)� ��'u4�{R'�����Bd82M��'fa�f�^Xai�,�)T��c�'v��*���8~0���		RIL�i�',�u�3,��I��*''4JRx�
�'�\�9����b�Ѓ#�� DԹ���$#�]��KW��|sh���BH&s�Z؄�L�T�2�OV!
Y��: ��I�l��zޔ��O�2J�ܹ#*Ӝ	R��ȓR��ai�ӘU�.ı�&V�@<"Ćȓ<:!:�a�)\y`w�4\��&����	=Q��Lr$P���X�/�5U�C�;O���A ;@�e"fJT���B�	�3�x�(��)������^��B��'zqJ�1w�>`�Kdۗ�X7� ��{r�T�JဥP%�_�l��I���4�Ik�'��'
��B���g� �˄L-�m@�'����c�73l�0�`�;��b�'SF�I3R5C��Ke�H<�d}��'��aUM���$�Ԡ�"F���
�'�l��H[�LSt\ԮO1N�<���'nd�kt.����z3$�4J����'>T�RK^$`��	�d3m�ԑ�'~jRFo�ԙ�,� ,����'(Y[ _�l~P�V�p���yR�IQܧ�x�Iᡗ�&^aI.�k�Q�ȓ,K�K��W� 9�\���1~��D�=A�S�? ld ��ۯ|�
��e��0"ʵ�V"Oz�d�� ��f�Z�1��q�V�)�	��?��O��aI4c�Q��K>�
��&"O�Y�j׆s$V��5��*��\�e"O���&+Vb��@��1�� "O��a���8 ��Y�S���Ts�"O��z��*qd�{��	,��(��"OL�Z0��	���"�Ոt�P����'��'�X�
�'f�r��i4%2/O���D�%:�@aE�}\
�!\-#+!�C�'�L=�&۾EgR4j�"��A�!���m7�q�i��*N���@a��!��U�A�6��J2DG<�h�@�r�!�$�G9�lQ���Ͳl���^d3!��LBuh���@O%}�����ߙd(!�R�U�ݳ�)�,%��Պ�B\ED�d4�S�O[U`�'ҵY=:�S�׈bx.���'-P�*|��![(]��hxf���~�'Xe�uɊ��I�Ba��`	�'6�	��@�#G�0)�`����'Q.�bq�C>ii�i�犟GrH�����0/ʼ�w�]�*��F6k����ȓL'<�"U/��b�h`���']�H��3X)�f-�c")Cr�V==U��	�D�'�D}!���1v2i��h	.n�P��'Ŏ@��#L�0�\%C�C��h58��ߓ��'�j��T�U�/I�tJ ��.i�L̲��y��T/U	�Ց��� Q�@H�aO4��#=������z��&��)k�U1�˚��!�D�����
U���7q�A��S�T��':��_��O:��?)s-��l�zT�f˔c̐���m��Xl��<9�@��Ш��̏81*l��Mh�<��f>v<��K�'��G�?��8��y�h�2Q�]^�b%�����<�� �ȓk8ܡ�bOʡ(�r�r�)�]��a��D!��4��em�� �(��?)"H�S�X���">i���׮k�e�#M�?��p*��<F5!��τg��i���N#S��q�C
�O��=��RLFe�{F��V�0yb��"O�p���H� ����1\���e5OFb�,D��'S~�@"�9���;,���'(�q���*0a�ǀ63�TD����?�
�w5�	����8wt\�t�
Lمȓe�d���L ��و!�*�XD{�'�8m��>[��I���1A=\��
�'��<[SL�N��ց@�@�	�'Q��HT|u����F��?��!��'&���ɚx7�p�*ϸ����
�'��Q�j�R�Vy�����3��	�'0�!��,X�#&:b-͖c`� �'�n�J"��:-p�N�
��x
�'�2�R���$v�VU�t�޿qp�I
�'�0-ˤ��]�F�C��2�l,	�'^Z�4j�������(�(	�'�(Q�O��Sj:�ŗ=L>Ҕ��'�\+t"�g���jsa$D�����',��	��ù ��͡J�
e�~��
�'�Ĝ�B��@����Q�ܵ�q�
�'1����F�=���a�	�\HQ
�'l �ahG-�T��@��?�PC
�'I~�@��A�E\h@s`�F= bh�
�'��Ya�Ls��Ms�h��t�Rk	�'BdyV�_%PC�%ҥ�O�l��8!	�'X<����
�}t^�0��\ò�i��� �<)A�E�-�8�O�O�x �"OvX#��J,n݌ X �A�nYZ�1�"O؄Q#�T�+�b��d�IR>�i�"O��ra��Dr
��Ed�ty�"O��@��[ꞁ(&����ZL�E"O��É�#rVI���Ph�"Oj�!��=*T،��O 2�@�R"O"�*���2Ul�a�f/W�0~��"O��ˀ(�=�L ڐ��$��:%"O�� � I�j�X�S�͑z�n�"O���I�9O�����W�
��H�'"O�a��F�l����h".N��t"O�Y0@MNHRy�c��F���3"O���"M0�\���6h���"O`���nY'<���HH�@uZ\��"O���ƃf��Ѱs�э>��a� "Ox�Q��HHʬB��'-"�B""Oz��#ʕC������Q�F���Ȑ"O����_@R�&�T�}�z�Hs"O��g�<&Ė�8�j�8.{��� "O�ţ0��<n46��0	�0o|�hD"O��EŒ�I�Q�5��KO�0u"Oȑ!�d�6#beP�ڙ\�:	�P"O,��#��7C��5L�A��p'"O�9v��L�VE`� <Chz�qF"O�d��A�w	$u� @k����e"O����$X#.<xh���|
�"O@5siZ����{#��q͖�S�"O��s�'�7 ��)z�h��l�b��"O&���ߙH�,l@��'t~��"O*�e!�!9?��P"�FDТ�S�"O����V#hT�QKT o<��F"OTQz0� �-��HɆ�EIx�"O�-�s���F䅢�i�	~���"O�5I@	�2n�pH���ڐN"���"O�蘡g�,@�l�0AҎ��	�"O�a�e͊|<t��զE��X�q�"O$|i�H��TQ�dt#��9��p"O���ס>+y�)��]�s� �+�"O������G�xKu�5gFI""O�Eٲ���^�SSN˻����"Oz��h�9*����MMW�-*�"O�܋s�^ 
S<#���/vO�0C3"O��i���%_�MZH�+E�-�Q"O\���ˆ�$��ڥ�E)0.�
�"O�%���?��i�V�B!P�.�E"O�ܢ�h^�&�&� ���&|�s"O@=;�R5xYP)�vΔ/�Ag"O�x��{�J(����
:�����"OI�eo[��v����=W���"O��yrBS�z5�52�+N6%���s�"O��#�7������2�4�Cd"OʄaBÓ?ev%�a��~�8��"O�9�(ܫ;���Qc	!��ĸ�"O qb���I�H8Y`h[,#"�D�v"ON��W�d���!��:�"O��X�H�(�pآ7�h�4cF"O����b�L ���A?�jY�F"Of�a�%�R��vO	#�l���"O �I�h�j�ЫC2�d�ʐ"O����L�\��!�_��p�"Oj)0eԫg����b��yA�"O���!@l��Z��"�j�H�"OAp��
 V�ic"�=oL�4"O� �t����\��}��P�ex�"OB��&�=�p�j*N6���"ON�z����z�ʇ� �U�Ă1*O���[
;��0X��0}N�'[~��ӑ.��9�C8gK�m�
�'Cʈ���%v5Jd3�=eO�	�'��(� �Λ4v�s6���z�'l�u�4��;4�9g E�&�;�'��d���$f+����� �F���'ݖ�hg�#W���A�zNft��'I쀓�'-x���=[��A�'oV,(W!��Ӡ�J���PHL�a
�'f\a�	�n�,b��&M��]�'!4UCC�3n試��S:��'m.Pp���%l�iJ�	��C��1��'e��Y2�K�"�0@h�'��v���'_�+� �#��iҲ��
�ب�'C����l�)���A� gJ1��'��HITgN�^�����L]�tx�;�'^.�X��xGX�c�%�<�$S�'h�-
w'�9T��Z�$U���}�
�'A� (�ǯ_��ɶ#�!�\9��'����0NC��e�։V4f�(8�'@y����=�zW#bR����'8�<��dG#��A�̕g@�'�����ؚ њ��rJ����'v�1�ON4Z-�GԪo�t�(�'���qv�C�QIx]Ҵ�>���'�Q�pǉ�`l�	�JS�=����'��3�mI�A	��wM��2�'�J@D�*:m�g�I�#�����' Rnd�Z��E��"V����U"O������
#�ȉ��Y�p�"O�=h��V!
$٢#N�_d�\c3"O1�� �9��pk�GF�4s�`�$"OR�W!1Lj�ز�.f���ڔ"O��j��Kg�:,	`�ڛ�LD00"OR�$��)׮%��T���T"O��+���_.�@qehG��VH�"O����:*|8(�GO�]G*�h"OX���N�:v� ����n!��q"Or���`�2���1+� g+�t�"O,%"�ȷ4��0!���9z�.�j�"O�u���dPJc�_�@JE�"O�i���ځn���8����@�)�"O�j�R�?"�pу�9@I""O���� Ġ>��,SB惮 ,2azF"O�h#FcKKd�$@V�".���"O^ �ڻM�hmS6�
�y���R"O�zK 
�21S�N��^}@���"O@����6�P��mà����c"OB8�d�N�%R��1V��l�|�3"O�9��c�a�p�sp'�5Yʶ��C"O"tn�{.�mцK�#c��,��"O�8��Ǵ8��ڑ��k�B��"O��J� ©t��94cE
��D�"O�%��h�hg��oq�t��5D�Pp�n̵%&l�Q�'X ����3D�@s+e��B�I
���!�D@)yh�����|���Ʉ�!�$X��{0��#�\�r��!�$G�K-�9�!��t��2��V��!�$���dj@��ZD-�G��!�D4�"��&eI�Iz���!�� H�Z��	�V���	W�� ��"O��B0�#(<P��B*,�8b"OV��&(�#�Fm2�jV�1�d��"O��B����� ���L̤٣"O���H�k3��p�%T4X�^8H�"O"ث��#�d�HeWk���;�"O��V�ÖPΆ�bw��X�$���"O�1	��5F&�E+���VQ�lI6"O��3n�}�>���	ۧ4>�T�S"O���ʿH�����.,8xW"O�(!�n	0RL\��"3k���"O:��FΦH� I��>�z��2"O�Y�^) G��������`"O�����_DL)1s΀�6�4ő�"O�ɑ�ƌZ�=rA�՞O���"O(��U�A&��D+���2v��p�q"O.��tN�pe�$���/^�(�"O 4X&��M�e;�n3S�X�@"Ot�8��^���#��Jܺ%��"O�=Z��4�$���MRĄ��#"Od���_�(��`��9H�$@�"O�1����t}.���U(&00�U"O>!(C��y���Yō�=/ �"O�1y���Rm2�6q�и"Oxx����&e�����J�0Iҙ�W"O��pC0r�ą��l0,\;f"O�U�4/�&I/�����#.��a�"O~� ���c4P���Z�	��1%"O��8T�F?f��k4+'ۺ&"O.$H�[�^�.��Q��_�ʠ�a"O~�e��*�,���֩I�B,q"O�D[���K<*��]��E��"O�i�D� e��9׉E-kB�*�"O|����<�"���*�$<"�h�"O��*"�ݭV^��B�+H_��ZV"OL!j@�F+��1� ]�cl���V"O����T�
��A��nV�5W����"O��$G7H]�	��FF>�e�"OL%1���=�v�*�F
{}�9!"O(M�%�\/�ݐ1%!C�l�s"O�P�Pt�� �
m���3�"O�����x�9�$(�"��HK "OX�0���/��Dcsf�9(��ɂ"O�%�ƏF]�DآR�Ǒ'�L%�g"O����Aǡw��񱎏(2�ځӄ"O��˧�]�#�L��j��"�Sq"O���6)��u]��㡊ؒZZJ�d"OjI���6}ⰲ��ޱdN@�"O�Pu/�1smt��1〾.���"O<Uh���^��b�H'b�	��"O�˰��/�����t��!I"O�li���B�*l*�A��mE��*�"OI�т�7X\Li$�ջ@���"O���r.Z y��I�-��!A�("O�ѩ���$1`�9���K6��"O�H��B��Y��Q�ra"OQk�O�G~-h�B!b8�$"O��-�z	��!�N�	Ѳ"O>�	��W�NT"Ba��2ᆨ0�"O�1��I��rl�e�b�K�u�X���"O �&)R�`[j%�m�d�0x9b"O�`xK>�����˂�_ҒQ�!"O��G�	6�H����V� ��"O�]	Ԧ�<S",� �2l�hDa"O� @U�=o[n��G`ޯ6��{f"OҀD��u,$��w�V� ��"O@��*G�:�����3�&0S�"O�Q�u��I�h�:�����t�S"O�H҇�\X��I��l1/�P��"O>�HC�}sh��s�P;��u"O�9rD)�*@�T���%ީ����"O���G�+d��h���'�t`f"O`�@��6�����(^��D��"O�X�4ኊn@ᑗ�ҭ�@�5"O|�u�K�2 l ����Fv����"O�����ϧt͜JP��f��9�"O�X�毙+2�>�)҄�?!�-Q"O�! d߫d!�Đd�;N��B"O������T��-�B��'�2Q3'"O ���o�\q ����"O�U�ŊPZ�`/�/%�$�p"On��*��fK�-?�8rD��u�<�'��3�2�C�"�����@�o�<�O����&�V�qd��%�]k�<!A.�<!�$m!�M�?�����c�<A����t�
�R�e��!�Py��mY�<A2&���t ������V�<I�e
���y�ˋ+x���CI�O�<�$�Hp30hP��ܜ>py�CR�<�0�e߄i�fN��z�z�Kf�<a����I4
�`��^�vp4� �Ml�<�͍�2@T�� �-X ��V�Sk�<Qn��}XT���͗2s͒�!��~�<�6���jY���
Ј_�ڽ�w�}�<�ď�O>>�ucLA���i��Q�<������#� Ʉr�fu� �J�<Y3���:-��2�S�Fͩ��D�<YGl
�E$�,2H�:{dMy�&�B�<	��
�@��,�q����0��x�<y1A
e��胧�+����w�<�3��9Y�I��	!`�˅Iv�<�F��?�dm+E�B�e#��Gv�<�֔+�T�W/��7z�җ�p�<�S��%]��lPCπ1d���'��m�<�$��"ao�(`��-��Qv�o�<i�l�;[�,<�� �$ k���G>T�d�g��yE� 呸 /b`@��"D�h�� YGv�KpP)�H�3�� D�|"���X��3�����`K?D���/�w	�@���w3�	z*D� �-�=}b�a���"O%��3��(D�D�'
'&��y��-F�~Z}��)D�����|P�0�L��'f`I�N;D��x�̦!\Vh�6�r�Z�`֬%D�l	L��$A�dI,1��۶�$D��Z�N�]� t�t�F�VΎ9(f#D���@� W�t[��� �t�R�B D���*��c���$}$�m
"D���R�)FE@��s`��D�Z�2V�$D�t�1�_R�(G��C��X�F� D�H�C���}�vM�� �W�dԩv D��1ğ"H�]�A�V$&�lm�R?D���,��o	��x��Hl����" D�8���b�N�۰NF"����Cc>D�t;%��E¤�HG�W'��=I�<D�p�G��7���[���Dl��e=D��D�<���$���ؘx�B=D�0������i���(�Դ�u�:D�� \�DŰL%z�	$*�#LL�P�"O�u��I�%C�Z42։D�'��S�"OZ�yG��bUZ(U�U? �Y�"O dx��յv�3��m�}� "Oa��hϝm���Ʌ�A�O04P�q"ON���'=���ps�X=x��a�"O.uKD��1C>|�r��U�j��͢$"OфN˩y.�"��YBl�
7"O��[b�C5V�n�3Ԅ )���2�"O����Ń`'�TqvD���b��R�<��@O�fyR���ǘ� ��M�N�<��<d�x�cj�w|L���H�<�HO-;�Pr�K�}d(�1b$�[�<	��n7��4b��P��K�U�<i���+K ��u�T�h�� (�J�<	�@ȝ/�8���-D�G^���FJHF�<��/Ǡ*̀59���)H��!/KV�<�3�i�rd�'g�%q�&)*A�IU�<qƃ�8=YX-�/_�R��Ic7ɇO�<�1�ń2��Kj�8^���JP�<y�j�	����;�*��2#[J�<AGֲpl�E��H�,�"�	όD�<9�,7+i���H�	t.��W��{�<��F�T�
��V-Z� ��F�u�<�5l�6�P���/�	HZ�a+C��h�<��J�|��CUo����	K�L�l�<)�#��ґ����op8�t�E`�<Y���b�4c�C�*N%��Z���F�<B��/Z�
Qa�[��\�zD��B�<Y�)C�W�$="�fV`���/A�<�4K	���I)�Β22��� �T�<�ף�����_�������e�<��fWz Y�kC���PC��a�<�FߒsP�����f��5���_�<1E�рP���F�S�>$<��OR�<�!�Q�C�����L,D�ZM�f��M�<9���'X�#n��F\��@�/F�<�uni?D�QÑMXĩ�S�MM�<1�"�Lɘ�/W�����p�<1s�[�I���Ae	�%�|�X�k�<���.��А$!�6mcD��s��g�<�cբ+�Q�EN7.�D����c�<i��b=,)�P�wJ�`�-�{�<�P���s���ٓ*�/3N6%Ra��u�<��A�mU�P�F`��O�(<� Lu�<	� �\��q8��Տq�\	��[p�<�uW� ��h��͉6'yv�v�D�<)4��$AD\��θ9ѰM�2,I�<�b	Ce�z4�T�Ǟb��Y�N��<)�.D�\{��C�Bm���P��{�<�!�>j�8�kD��n?&�:2��N�<���#���hQ)� ��D�<�#��-a����G[�&�Y@�c�H�<�u/��c�la	�D�Wtě�B�K�<�B+�
��)��]�o�l�CK�<1�A��fRa��V�RQ�AFH�<a����X�V�S2ה+��d��hLI�<ae͒'�<��_i�� �O�<�����@��C�G�9�\ ��H�<Y���1S�� ��L�,y�1��DP�<	P�K1��q�/�M�\���(�c�<)��&]��L�ac�rt٢�RJ�<iE�,�J�
5�K1r���L	J�<��BR��p��T��d�@��J�<� ����GٿyVf�q�@�A�]��"OԽbsf��Sǎ�
Oɍ�0!��"O"u{o!)�8�C=�p�1W"OZq/އS �����ђD� A�"O�`i��M$KʎD;�����h�T"Ot8W��aI�����N�$4br"O^������!K� B�&��p��"O
�IGo�	?Z���U�T��� �"O.�d�"?J�!�ʈ�{Bj�;V"O֌:���4�&@#T��/f;���"O
`YH���V5)�BܙD�ȸ'"O*�r��M����*�;��"O�\9 
ӵ6�!@j��j�rAQ�"O69
�ԫ@�L��I��|uJ�z"O"��W�:3�9����N�X���"O� zP�N8L���kŌ(Ɯ)�"O��P�B�7?j��)-Yi�Y�"Ol��K �hYځbd�:1Us�"O )R6�O"FM�Y�_r��̊��y����<���p�G1(������W�y�E��d�,�Oݥ98�� ��yR��-@le���z��*�)�y"ìh "�xDcA�k)8ыr�M��y"���֑��G�5�!����yFW
Z4�h� D�\@�XAFY;�y�Q�xJ!���WR�r�A��yB��D���d�����	^��yrj� �����a�b�Ĳ�I��y2Ϟ16�������v���ܑ�yR�O72�!���:g0�@e�V��y�'łn�XX�� 0	h����yr��`�B$C��,WJ�5���y�m� �v��A�.�X�nC��y�`�%m^��%Nًc�nQ��/R�yr &Dt�$�n�%a��7c�:%!��)P����"�� �
)R��92-!�D_�j;��
W��}ke`�?o!򤛁0�Hc�a�	�4�p�N�1K!�F|����E`��y�Ј��ȍVC!��;^�
pF�C��^�����a!�DYA�`	eޤAf��
�%P�qP!�R�((
��o�%TJ��E��)B!�$�;y�J�a����W��<�u�9t\!�ِA�$�ir�UVq�Pq`Ü�$5!�ą�j�|� �n�qS߉(!�D�?^QΤ�6$��a]k!�c!�$�7�T��쓉 ͎�@�>`!�$�9v��؀�W)	�xb'�O:j�!�d�
\�"h�L�U9�C���!�dHx��9�P���Id� +�!��6��
��F�d��l֨R"U!�1K�I�G�,�D���(\aj!�D�/(6vc�I]W�X�1V `!��@������a�`y�g�3E!�DU(sqF��rN<��H�rE5>!�K�g�^��3�-}�"7���{!������s��=ji�d	n!򄛄� �H����E�x�!�Ǖ]N.�拌�5t�݃�b��Q�!�Q(��t���Q\&0���N�!���`��耪�5>ނ��ХZ�:�!�$�{��M`U+@_�v p���X�!���~ �BA�Q�"A��A��.~!�D� gbsTOP�5�`m���ݻpa!�� �����1�N\���Z M|0��V"O���W5�숙���8b��`�@"O>I�1��b��ZԢ�9mu�P��"O8��DG19vA!�!�*u�S�"O�e:f��!<֐7A�&  QI�"O�,c�OG��Hi3�_3C�B��2"OY�N�[]v�*�f�N�RY��"O��2�O�"e��ȡ%�J�b�U"O$�bM,�r A�.��IϠ��"Op��/Y�%��.��ɐR"O�+�
��	�މ	���o����"O�	8�Dδ�L�x�^�f,c�"O�-�`��o�`�4�>@p��R"O<E'��:r�x��uǚ<UE�p�"O�{�噍��e���e���C"Ol�g/K�>�0��D[�&��)�g"O|PF�DwDĀ���XվU"O֤� #�6%���Մ;B�(�3"O�bf]y�v�R%ĕ={�Lۂ"O2��7+#�x�@"Q6CM�${u"O�1r2Lʤ9y��E�82/���"O�d�A�	�),��@gI[�h�����"O\��&5ST&Iڂ�(N�K��y���?�Peғ)ܨ-�|�D�β�yB��|V�2&`A?NT���` ��y"%ΜA븩�ܮK�PA��yA��|��%�g�ʦ@�Z\�0���y�k�?u����pg	?ld=y�(�6�y�G�Wy+�m��2{Be����y2�\�U�}���N�v����r�Y��y�5z�1d���la�,��k��y�/�&�u�t	&h�| C5�V��y`W..7�1��+_Ö��Ca-�y���taf1��dQ*H�|(�S���yRÉo(�!�Va��E}�{���5�y�΂�H�6�U @��؂���y�dݍD�0sK�8�FaHrn���y�i3r�h���h�98.0dR����yb#�(UͶ�$#�6��y���U��y�$��H�P��%nH8.���x����yB��#h���A!��"����3�D.�y��G6R|�-�g�ͺ H|P%�y�G�Sb���i��B�5���6�y�*E�(�1G�Đr�,Ɖ���yR �OZ��֦��R�ph�	�y���)�Qr �MLe�@��y��'6`X8�C�S��,���H/�y�$�%��`@EKMe����V�A��yro�=%}8p�b]XQ��궬�]�<!��T�qn��X���7�؅Z��LT�<���{.�{�%�W�z$*���J�<9��ʔdp�1��A�B0:��B�<�怭��06ń=d5VTr f E�<�r�ҜH\�В��,����e��I�<!�@�~�hh+􎛰FqJY�ʚ@�<�K�75v�A�wX/%'0(0Q��{�<aUn�'R[��J�/©N&��3'�z�<)�l��P��eJ4�A�}��=���NZ�<1���;1|!x�(#v��x���W�<I�.լ;Z����2�n�0�j�R�<Ӌ��ؠx2	��*����N�<Q6#�"Ęh�bG03�|ȱq
BN�<��P�^�8W��(q�����GSc�<!��2#�`e"Eٞ�f����QF�<� `��3����1��I���3"O44)�H�F�s�t��U��"O��b� 5���WG�(:stq��"OB�k�	��q����V�A�=z5As"O`��
�q�ʩ��@�-��	YT"O�t�@��Om����B�7 �Ԡ�"O�<Y��.EJ���C"���)��"Od�b$L��T�;���Q��&"O���pd�G��i"Q�Gǎ�{�"O@0Qd!�T6� k�M�Lb�H�e"O�L�0�#�$ܙ�
C�wv0�R�"O�qժ�4%�Տ����3u"O�(@S�84��Aeׂ i0<��"O��	��S��t�u�Q2]tiY""O�`�͜c�0�j EJ�kRp屇"O�2w�0$hH�ء��Nz!{2"O~�X��Q$�r)�L�s�v�Ȱ"O���$ەF�m�a�F�mی��%"O*(��ͿEF��Ғ%�.�\@�"O������ZB�����;�"O��a"M�&z$��C�2�4P�"O~��Ve1 ��<`E��!��-C�"O�G	�-�8�ڰ�& ���+�"O����M,mQ"Q�c7i��m�"ONZ`gL�x0�b�fH; "O�M;6LU)0I'g�$� ���"O 1�AD��	th��#[�x��AS!"O8�f���Z#
�(0LY>;��eHu"O>��!�?K�(�듳9�X@��"O�i����l�0IA�)��8�"O���ւ��.h,�(`�G�#�Xt��"O4I	����zך���?VZıC"O�i!L�\��L�W�m���p3"O�C2�ރ'����-ń�(�[p"OhP�#�H B�q����Ll�Y����I�P��2v�֠UN��q�y�B�I�"d�ԧ��b�c�Q/��B�	�k�.d���@�c�򴰆�3G��B�	�:��捤z��l��N,c�C�I�75��AT-�i��	&��C�#c���KFe�|���w��<]�B䉳��A��O�	VD���'\�7��B�	7i�����]�XB��т*D��js��;�8u�%)s!��6LInB��jXriص�.2�ԑZ�(�B�I�$;���$��%o�A	"�ۭx<B�I�Dբ2mY,z'�`&��d��C�	�J�J��TO$2���@�"��C�	%*��%D=����7�/OTB�	�-h�"�� -J\�`<MtrB䉪bNj��G�[<=�n�:�`Ά`R�C䉅<�i ��c:���̣'+�C�IQҊ�CǄ�gK��bN�!�C�	�x� �@�w���!��99�C�	�{NT@�w�K�I�<���b��~C�	� VpAt�ą{�$��#��<Q�B� L[1Y���-�е�4aR"/�.C�IӸ�"�+<X
�Ґ�ϳA��B�ɖ*��!i�+1�0<���K0NжB�I�}rx;�P�����<��B�	����ڼ�h� 阕S�bB�	+)��|0�m��8�|�J`E�
	�B�Ik8ĉ�g�>$�@���$y%�B䉘A�
�K�̕(2���g@ʹ�B�)� fdI0K�%]�zu��� K�T��"O0�8V���^N���-	��	�"O���	��xp�$�&8[�<a"O��d�݋J�	�V��Z� M��"O�l`�H#iX2,B��e���y��f>��c�J�W�0MX�%��(���&6D�x3�-8{��$��9��5yF)D�` To�+0�:�9���L�u�A'D�db��X�#X�+����N΀1ZT&D����^�p�a׊�c%ja!��%D�H�#�Ĥ?�ՋRE?o}:7#q�<Id�Q�"�(� ��K��M�u��v����"�'tZl�Ǝ/cW��IS"��ʘQ�ȓ,D)���@�#~ॱ��
dv`D�ȓ'&�(y&oUv��A�lC�P�����T�SNW2|�QqÝ�m6ڵ��eM������XGT�Oҍ}���ت�����~����l�~#�ՄȓUq��0`��"R+ĉ`��*`��6��#�S�7� ��#�x���G���p�)�C{�%�ׁ�M��m�ȓO�RT���X`^0R�ͪu��@�ȓb`��{kƎbj&��Oӯ~�h��Ht�j�w�x �Ɂ`�B��ȓ�j��@��	7s@���7���ȓv'���t��t�<���4Z��L�?Ɍ��~:�#W )��#����k��8St
�P�<QP�Oa\���O��
�:��E�<	�C��X�X�J�$�BU���<�#�Z��"9�B
�o��L�d	Lz�<�f����-1pG�)�L@��K�<yEO�+[�z��Ç�y�`Q��j�Q�<I�@sV\��&�[�4���j҆J�'�?��s�O�q�qR�O�C�,]��#D�t��mC�R� )��ͮlp��D�"D���C�H/e�,c�N� o��Dxt
"D�L�$F۔I�`����O��\"�H?D�����O���B��l���'D��`s̞�j�=K��R
p��0��o#D�(´,�!�(��l��%�l��,D���pih�$(�ALS!�Fб�n?D��
FݫXi��K�M0r�:�i?D��1b�0g.�L �j��YT���!D�D��� 6��s�C) 7l��1i>D���BeԞM��s�k��e�N��C� D��Bc�=�X�Cn_�C��s]pC�ɢl�z)1!�@�1=�ʠ)V�s���D$?!�H.;�іmC��`�M[]�<�c��5�0p�Q�_Y���q�W�<G��/[�0���$Z���w�\�<	֢ȕ%��(3��Y�7��@���Z�<�ЈX�Y���B��8p<q� ��V�<��([�u����.H$�fa��`Pm�<� i�+�l�P$��]K`�"��d�<�Dm��z'�l�rfˊ@F�DɚL�<�.�|���EI�}�I��g�_�<�L�m��YXP�x�L��Fi�c�<	1���OD���*���d���g�<a2a�	��Pd�'�(q�FfVd�<A�oq=�2�rx�9�U{�<�0H֡"��;"�Z�8��u��w�<9��0ts0�Ye��*D��J��I�<�vCW�H]n�!����"��hR�^�<V"�Z�(�ّ�K$>���V)�Y�<� �$�w Ր,�JU�UG�X��5��"O�9�qF��
x$����8R
���"O$����9.l�Pp�mG9�&рr"O��i�/j����&�,����"OP�*%dݝ�-��F�D"&m�d"O��3���@�C��
%}����"O����B���F)w,�	_NM!�"O"쉳 �q� m�@+��f@
���"O�U��YS�mB�j�H���3"O�A��ד��U��RfT��"O6�y�m�xQ$���.G�o���{"O���'=\!n��O�1y*��"O��@,�p����F5u\��"OEc���enl��͝��BG"O�� *D�.����*7D��胕"O�jí_7R~�0IR�M�F\�T"O�y�C�	��ʦ(��9k�L�"OH�p��C=Va@1�HR34b�-�"ONm��^
�,����	4����"O�$C�y��]J�� #���"O�X�A%=Y(Ѥ��8R� D#�"O>��.�:V�ށY� ߕ|���1"O��)�
�+AJ��s ���#"O��{��%�X��w��=��"O~�["٣]I"�����a����"O @ ��E/��1/^���)�"O,(1��կ,��A@�A#I��X�"O@8s�]XĀ0�Z?�%@wi�[�<�T'�]�B���k��+�x�s!�]|�<AA�P�&YNH��d��y��@P�S�<q���$�)��c	�m���D�Cd�<1��ӢJs�)���5cY�E��͇^�<y�'JSPȚ�aP4f�@y ��X�<�G�Ibe����wc�����M�<���L�X��Տ5�Lu8a��^�<��'ϱ_�h���l�D���u�<�s���d�lx+vΟ�Cd�a̅t�<Y1g��<����C�	��	aנq�<ɀ��T=80y�_�0T��BU�<	 I^�Z<
��c@�3�_{�<y�,�*_Nb�Q�-���ј���s�<�U��dM�l9f
�-}�F�0��m�<����A8H��U-�(P���+�k�<����![��\ڐ�ƥH �fdi�<%cF�T�r���bH�v)�h1�\h�<QAnBA��9X��?J;�� �^�<�G� G�dh��E�<h6�#Qb\�<aDB��w����	��܌�d��U�<�@��0��q�g��$'*iad�O�<a@&U�7hr�j Eϛ2^86�Yv�<���[``(�������Q��M�<i��PI�����ZI贸h�u�<AgF�e�v��_x���!Wq�<iv��7U�T����(?��DK�g�<���ƅtF8��a¡c�Mq�b�<����5p��s�/��%&�C�<!T%9�f5B�τ����b�B�<1��{��E�Λ=��xBNH~�<��yD0����l���WIE�<�s%�qC�eS⧀�#����G�u�<��'	s�򳌞�#�D�P�l!T��b�28�bf�Y��[��:D��`�A�$N�`��@��j��"7D�h��؍D�A��I��CQ|К��5D�� NL��dǴ���E� �3%�Ѱ�"O�-Kt�@�h�S`�u��k�"O,�i�c�Mr�I�R��J��P#"OZ �/BX*8 ��0[Zbx�"O4|y�׍Z�؛��ױiK�aw"O�-"���$tp�6�<,"�Hp"O�\�`�Q�\>�a��۸����"O@P�M�w�$k�,�8Z<0 "O��`�"�t���|�)v"O�H�`
C#ad�8e)Tmr�a"O*�ؕB\�VZ�1c�Fă)�t���"O����Ҝ{ff )5��U}���"OHݠCM߀t�l0B�ϭK�<��"O�ܠD	��0�k�W�/̶t� "Op,c`
�-�j)bc��R�X��"OX4IJ��3'BYd��Q�r̢�"O0�R.9V����-��I��0��"O.��#�:S��2��/e~�D	"O�ي����^<0�f�Ђ&�d��"OP���R[C|� ��Oh�)�"O����7���p��T�h�c"O�8#1�D�"�$q��)v.�:�"O��X�cH<ߨ���T/4���"O"U ��Q�\ސX�!�e��q"O�Y�f���'��h	D�@.L�l�v"O�XX6*��F+n��e_�<|dPG"O �:����.)# P4[BD�v"O�q�ǁ��cN�"�ʏT)����"O6��T.�>8��V G�T���"OZ��7/ ?sݒĉe�O
F,��!"O�QB�a&�������
�+�"O�i�
.`+ ���Gڜ&p�eВ"O�qJc�W�$���ă�F0Z�D"O��G� �d`�4q�c�>�ԁ�"O��� �ŉ*Y���WI� XV�"�"OԻ	M�dT]cu&�7T[zL�"O�(����f����r&�
A��q�"O�$��@�������(�)R"O�� g�F�B�&1ʱ��"���j�"OU��	I7q����5͕9� ��"O�q�"a�?`{�8z�+˴����%"O8Ě��F*.QH�+��
"��3"O�a+�A�<gD���J,E%"�"O�}�$�E�y�pm���>���"Ox��� *Z�.-+3@�2�V���"O,9 �(�;.�^�H�(�1���"O���]�(��@f�Q7$��$"OĐE�E�8�,�Z�OSl��"O � ����y*�=�� ��6�|�"OT��ď�%w|�!���V��P)W"O��tf,Z��X��1s�IXu"O\m�4�	j!��:�i�,]4u�"Ol��֧��[���	���*QVL��"Ol����� Q�\8	$e�5���#"O�ɛb��7n�\��#�$7|�a"O�0��#B ˑ�O2:�R��A"O�Y�P�X/J#�P A�%��)y!"O�x	��>��ĺ�OZd�ޜi�"O``g�A8P��؋�IS�4��aPA"O6�ZBh�:n�TH��*� t�d�"Oh��⭔2w��K�D��=k�L:C"Otl{�ٖEp�X�g�N hα��"OZ���I6fDsV��Na��3"OL��Ti�=�����AS0[S�]�2"O� :�1LNC�R���K�;�	c�"Op��G����f@�!n�N�'"O�6"��I�!������"O�ԪE��_�ɀ!~�<�F"O�dRTI�<����Ɔ.'\�J�"O4����v |�4�ĐG��B"O@����ΛU�	0�@\�H���"O|3!,B
h����@\>B�AB�"O���+�;}/Y)0��!`��-	�"O�y��;�j!��bF��:7!M�<aH� :l5x�GU� ��
dR�<���^f��B
��ҙ���F�<Q �7::�[q*EI���X5ėA�<�1g��V4���
�N}��P&\w�<q�
Ԫ����oO*�B=���Tu�<QWF��Hp��^H`8$.�W�<���؀!�M�:7l��k�
Q~�<�3͌�}f���ȫ���cV	~�<�v+�VպĹ�A�{����6�@}�<�2	�?���G�%t�t�����A�<Ʌ�L�����
̝aPi� �U�<�@�V�:��i�� ͂�!	NQ�<�$�.�t��sj�~�t`+�v�<��߹��Yq�JƖq6Y�e��{�<Q��L��X+��ґ	x�j� @�<9v)��o(��b��W�#�\��BYr�<�g&�36z�q���m=�M($�Zy�<��Jɟa0�A;���?p�, x�e�N�<�,ś^m Y����	�`�3#`�S�<-e�Q�2�
 �X��/�3�LB䉿)D<Āc
���x�P,���B�	d�d4D��8��`�#QB�I��t���*�b4����0D�C�I/R3�5ʦ�X�}H�����C��20v�6L@��>���9X6�C��G��� �j) t�#�΁h�C�I�q��h���$�2˱Ws�B�I�z�$�K��]����B�NR��B�`���3Z?u�Ĝ��>5b�C䉲$�{𬍚!Q���(�#�C�I�
�"���d2aĢ��-��(yB�'��h1m�:VΨ)��Z�V@8C�I?,�hk4��<ϰ8���h0�C�	H패���S�7	�:��-�fC䉠��ԫFa�=BAҍ#��0q:C�	� ��e���֑��s�b]�q��B�I-:��5�`i����C«Y�%�C�	�j7�xu$�.g4xH
M
u;�B����Ta��S2Hl�B޻ytC��(yZRqb�eٳ/
��6��y<JC�IO&ֈ��b��c��]b7 �h�DC�	�$r�\�AD�M���rCL�:LJB�	19ĉkbH��5�a�b�ʐO�0B�I�t��T(�A��m�	x�!�N�jC�}e&Yc��S�d	��ܟAKVC�	�V^��x6CP�?U:U{JMt�`B�ɠ���Y�;s��2ʌ�l�B�	(�p��ગ()I�U*fޢc�vB�	�`�P�S�aW% -d����$k��B�������԰M�����[�C�:j���1�eM2-��Ȋ�	��\B�	�~?�����5y�eAM){x"B��5)���(���a�HA(ʂ
yB�ɐ%�v�y��D[LպS$
1/�C�)� ��s�jT�>b�!�"ʱr5�hT"O&q�.�,0�$���!����"O��/H&��BA �?C� ��"O� :#cW	2���{c�ӧ�2Dh�"O���I�"�T0�FF 5�8��@"Olը� ��	��	s��-u��J�"O�tрϗ�W&���(߆T`�"O�c`��c�$z�g]�0_�|�"OA��$������ B�@)�"Oޝ�@B�"U9����B�+#�ّ"O2����	!F�.Y���U&z� T"Oll�ä�Z@�!���!��9�"OH4�IA)�T�`Â�>�)b"O�-Ic雑~�DYTi��BAE�'_!�� :C8�C4�������6v�!�Ԅ�`�ĭ�,|����ׂ��hG!�Ю=U#e"D�=��L�7➴D�!�R./|ɘJ�	����vf��-q!�� �B81�B�7MZ�ХA�&G!��!\F���$(:��#���FB�I�Q�J �KEU0�Z��ɼ#X�C䉃���Jp6U�	􇌥FrDB�	�+�Ԩ�6 K7��C$�(l�C��'Vd1CV$�ON��7�Z�~o�C䉫E�R4b�+;�+0(�Oz�C�ɎO�$�F�ӕ_R��cI;��C䉏��]�!!�N`��6��{KfC�	�d�
�^9�"tY�dV020�s�'�|�)��P�V���@ڹ3����o-�h��	/6�@g�Bv����3��J�V�	$@
��̶&����ȓy���:ua�$b$�37aPɆ�>8��A����M�B,Z,~�dY�����VJJ�	��yx'��&z��Y�ȓ�D�#�N��tXS��i�rE�ȓX��
�/T#� ���n�N�����.e��LX�!)��#�H	���L��9����S���C �s1=.���ȓJ~^��%mHj���[�e��YD~���J�����R��h�h�<~W^���V���񴮍�[�(��'�;vx ���+튤��=DZ`��!ϗ�}�"��ȓ}����*��#W�������W1��ȓQ���)rɎ�s���g �pܺ��ȓ1<���Θ�8�(�Y��{�F̅ȓtǈ�R,�^�(đ�i!xX�ȓe!>%�s-S1N������\�:���T��ѡ���d�)C�hY��A�J�
u��0t1� ��(vx��:�j0SH�, ��9��ŏ�@@\U�ȓ��¶"�y̼;���K6D%�ȓ'��k��7qM#A���mH���c3��*� �:t��E�D0�ن�1	r���C�pB���� |����ȓr��{0b�b���t���ȓ]��4(�̞
sN�c�I�2|iֈ��SF~� #�/I���j+uCX��ȓ9�z��a͈��"��G�*@�j���|�~=�,̎C��R�B�Nw���ii�)���16��cI"���ȓf46�c)$g\��%liZ��蜌!�%�h�����P,P}�ȓ[cJ�!'-��f�ҝS4��V�2��ȓg�"�@��E<BV���Js@ށ��S�? l�R�#~5V0�#n�9D�R�[u"O����_���ݘ��@<���A3"OD� �M�P"�a$��T�xp"O�1�N�v�0	EjҰ�6Art"O����۫�5�׃La���"O4P
Uc�(�f8��ٜ�fI�c"O�k�*!:}rx!C	�~[��C"O\�h`��"��K����Y`����"Op����@��@y�%OUa���"O���� ����ϮD0����"O�Q�EA/QlD�Zϙ����"On$���W	.�pYQ��i���Z "O�A��EǖlҞ�!DFY���DZ�"Oȱ�W���G�qZb�Ğtx���"O�����!(�R��G���^�$�"O��YA&s\�8�ME�tP�d��"OL!���DЮ�c2�I�nA8�QV"Ob�	"(�>�HQ���<FΠ��"O`!0�o@)u���F�	�Y%��"O���E���e��Hx2�"O`���
�$�@%F�gp���"OzP���Jx����R���W�xXW"O�U�%��v�h2�;g����b"O�AQ���)D�H1y2�b�|-YQ"O��6��>
8pf�7����"Ol�"�ۖ �Z�����P�"OI� h�n��=�/[:�"��W"O�(�s�;�~���ݐX~F��D"O|��N��%���XxވB"Oj$�6$�(bD� ��4��"O��U���2�O�,�jW"Ox�8�ɴS��)ʒV=W�@%��"O�Ѓ�)�[AN@�vkש<|� S�"O��8�OK8h�\8�ЩŜ	�v�AF"O&£�/l�f��i��twR��"OPl�"OL��p��'��7gd��5"O��1� �i�\�ܨ;�2ɳ"Ol����7D	�<!G�{�T�"OD8�b��
�"�%A'$xYZP"O��h�5��
��qL\ԉ�"OlP�E��%�3!�� �h]�"O�)�P�R?����  �X�&0
�"O<�a�ݡG��@�i��'��g"OR Zr��"_Xx0g�,a$Ƶ�U"On�+ElҼ,���#l�w��d"O���`LWP�T�E*Aa�Z�#�"O�UG=��Q�qǖ+�4i87"O��2�f�]� X���Z�'�����"On�8�/�Y��\��ӧ|s^0���	a�O=(!�(Ր*0�ȉqE<_�91��ē3o��"�#
PJ���G��Y����z-��v�(d�P)�PEͮo��ȓ;HB1�0㒝Qt�! ��2J� ��ȓI������\�C!�;YhQ��2�䠓u��L������X�Cކy��7̠��EJ�1r�*� �n�3��ȓB����7�u|�r�C?0(���H,XE�k�t8�\���b�R���^x> y��N�BZ���*Mj��9�ȓh��cqo!�"�aCD]�)�.y�ȓ7Z(A���Rr�ܸG,�`/f��ȓOY��Б	��W��檀3�j���zH4`-ECQC�]Ty��z���ƹ(Մp���"eH�ą�S�? r�P7n��f�r��v〉8NpÓ"ON0�p)�/P"	��F�|�=C�"O�ݻ�E��az��e��T�4b�"O84a@<ep=ɒ$�:K()�B"Ozu�K�~�����D�8y�Dl��"O�,!r��u�<��bF����ң"O��1�#�^�z�Bb��%z�t�d"O(U`��
� ��b�����ӷ"OP�`BjL�R���� 8�z�"O�]��iŘ2I����X$���"O�8�ƍˌ@�H���E�N��"O�h��o@<3|� �D�*���a"O�4�׎U	��!q@���h��&"O��Ӱ��^|>���+���!�"O�m�1�hf8�e"gy 0�c"O4�"������w�GM���"OL 2��[���M�;���"O�(B��=u6,U�VBG#�M#V"OZU�t�ʒ���h�B�#��tR"O� S�+D�7��r`oE�a�Π��"ODx9����tӕH�$;����"O�5���#^�t��W�6�3"O`�z��N�eZ�THSn_�H�"OĪ��K�i��, ��<9��#�"O*W�	.�Tr�"H�nbT���CH�<1�j��m�&� d��=�2�"��|�<��C�?6N����Y⧣���'.�ᛅ&�+�Z�b`��֦��` �� �荺t~�R 'J�X8|��,��q����i~�t*2��D�ȓ2Z�\rPmȱf�J�c���2M�z���n��
�7W8�U�1GE,x�ȓ�)8�X�x�J�
7�ج+���. �u�� �x �C� O�U�ȓ!����2@�Q����f�
'\n�9��RƤ��wl�85Jj��2m�%j;h���:�r��h�#T�z�p@(��!���o�T�EW�&w�Q��`K�0e:��?���{��V�(� ��% ��ȓ&��y�C�5��B��3mM���&`�Y�釹5�ܐҷbE�-j�d��L5��Ȑ��@�ó(��d�ȓ<l��1O��K��ա�	<�*i�ȓ�d$���U`�L$��JP�c�F)�ȓy2$	���N.�@(�0�H�1.j����D�D�7j��tr⍐�_�आ�|u�=�q�r�Iё#�;c:�iP�'����A-Z��ѠϏ�)T��Qش�Px�6~8 R�ܗ�~�1ӆ��y�/C�Y�Z��� �(D,V��yr�K&�<��ǫ �|g� 1��y���L��H�
a���EN���y��4;%@ӴcF1])h��d.���y���\.R�����5$�2�b����y�Ei���3��'e���$�yrj�
ވ9`��v�]�*B��c���#I�3�(0��oA�a�XB�	�w��qѳD��P�,�Kd% ,ϖC�	B)�e9�O�NfpI��\8�&B�Iu��x��"ĚQ���{pM��j��C�	�,� p	2�� ����X�C�ɿ`A�����(s�=`�[2c�nC�IJ��T�C�;A6fiS�oE�_>�C�I�VZh�)[4}p��� Ī*�C�)� ��"�iOX5��>��["O�0��!��_� �!®F*T��V"O�<�'��{�PaQg��XIL�p�"O�!��G<�։�¨I=?6"(S "O��JթU�BDTm��I &���s�"O
�0��0@�i@�KUP���"O,�sw�L�+��	x��Z/��9�u"Oܐ壅@��9��92fD"�"O�F
]<Xa&es'��X+�� $"O�$)�G�jc\��&�߀1�UkQ"Oİ�Pj0j�}(�@J�"�pI(�"O>(���I��՚s*He��`1"OEi��T%���L�B�d*g"O���cV�5�i� )~L9��"O,M���A�B1��ڵ_3�4(�@"O�A�!eܕ!��`���6V�d�3"O�8Yӟg��h�Fމ/F��"O��*�G��-4V=bc�שv�E��"O(D!��I'4�m�2��y�2���"O@Aۧm�$�F��gHªJ�13"O�U�0@ԗt�Y�喥&��X0"O����M'+��3�����pB"OL��2Ó�T+�@��AH`��!"O�Ö펽%�4�2��,�&� �"O��2N�Noֵp2&����v"O ���(ư���)��@�"O�M؅̗�#9Rу�BI&�|�k�"O��$@�"�dPS6G;
�X�P"O����� `�� ��5.X�0�"Oe�Ce@�-(��:�苖"¶��"O�A13�I�2�X�Iߩ8�"��"O2����	v����!�=1J��d"O�ph҈�*^�t ��݌&�B�"O��[ �Fr	.���*@6o�vu!�"O�C6�T�^� ��Q��AG(}�q"O�u9�8x(^��G��R*�y�"O>x�1��V4$$��$ �O;�	s�"O����?%�@��%!��N�^��#"O�����l%�ʳ��rx���`]�<��焲Q��غ�JN�_��	�׏�[�<a��
J�����-�Y��٦��W�<�A�;�4��%�0b�>]�A��Q�<�4FP% �<da�$�'8��mS�C�M�<�iܦk��u��"F��#Ea�P�<��ŋB<�K�S�!q��B���M�<	7��d/ ]�#���w
��QO�q�<A%��U� �q�ȽF7��(b�T�<�&*T<j�XD,�+������N�<�U�,`!�t!��_,���Q�H�b�<��MY&?AYC���t= KՇ�D�<�@�,���`��aI�x��K]�<� �=,��Q#�
6�%(w��W�<���W�BMYX�ꆌ 	pEB�g�<тg�1c5���f��=x�b�]�<y�D�?H�8)��	�SN&�a���a�<�%1}b��S�"�A�Ēi�<	�/�"��!�G�<��bsm�i�<�֌3nzQ�SÈ�kP|�!��`�<���@�I�L��M�6d:`}2�U�<���C��T��d��$ct����Y�<a0)�l[�Ѹ����e�: `W�y�<��%Y8K�̸:��P?h$��0�v�<!��J�X�ViP#��)*��� ,AZ�<���D�r���O�S����V�<� B�tB�Q֩�Ќۄl�	g"O�|�Ggʳ?�Lr���_��4"Ot���+Џ<��̂'kH�AY �"O�  ,��y��J�ZOx��"Ov�A�"ޒ	�^�9���<f?<�h�"O�e�!'�=hچ����w%�%3C"O���؟N� =�r� @���"OfO(N�eH�l�P�l�"O��Ӡ�1He��a�
�.ɀ��"O��XG�@6m"4��q���Ķ�2"O�<RV��n���[$�)3�d�b"Opq�4`MY�;'�N=D$.U��"O*�
���dM��ӕfG�{���"O�iȲ���ظ�-AT!9'h0�y��,�$�CR�W�q��] f�ڎ�y��'V��t��g_5o=@�u��y"j)yL��@�Y�of��t���y���c���#�具m��e��1�y2'Ԃp쐑0EF�KT������y"NȈH����E�PAd��d�D�y���<u*r7�
�C�t(�#� �y"+ZR�{�lׄ0��Q\%�y�0Tv�*�&��0I�����7�y�g4)�nl�+Ǖ?��ۄ�Ǎ�y�g[���4�b��-�����/���y�d]\x�UHO�_f�qrCc\?�y��_?W>�(�V�<�*4#�W�y���O����.%;���Ҧ ɶ�y��1Hm��*�*�mh�ߝ�y˜�'���bA&}c�!`+��y���2Aܪ0����/\��gm��y�f�����"ll
w�J��yL(/hQx4�6�B�0� �y�AIᬘ�7U�(xi	@�y"$�,R�Feа�\�1�$裣[:�yr���m�,q����> ��般�y��F��B� �*"h�@0�@&�yR�[���@�����wM*mӲ�]�y���,Z�Pp�T�.nL�Q3�@�y��?
��Y�@䄂a��Ɋ�y��N>c��L�.�I� �is����yrG�.��
7B��J���b��O�y�I��6C" �!\"x�*�X<�y�� 1W�<Y�F�Q�>	���J �yr`�;(X�uB��]2W�U����5�y�c���b(�t��TÂ��b�y2j�7^�ck�8�Iҍ\>�y2n�I$J8�DJ��82�����^�yR�ěC�.�
t�7\D�䤘��y�O4���W��5�0T�ް�ymY�(E
��-�P�1�S5�y��=8C4�r�C 6U��K!�X�y�ǚ/1�舠P�ͷs$ָ��J��y¢�/$�<��!x`&	+P'	�y����|��ԫb��?p���ʒ��9�y҄�91�杪�f�2y��J�\�y%M%9r0s�@H�}\< Z��F7�y��L�%8@s��ͳs\�ы�����yR��y��)U�ߝj�Ɛy/T��yR"A�&��@��,�3�T�rb>�y�ʼa��4Є�V�*��ro_��yR#F>RR] c��
������y�J2��	`&����H(Uc���yҁ�9%�t�b�$H;��'���y
� Pt�fMN�mԜ� J��h_�(�d"O:��4gM
=�x��T	�8nhł�"OT9Z�+�(�ԩ�	�oG0Y�Q"O&P[���'�X'�E�a8͙W"O��2�/��v��D rɶ�\Uh�"O�m��BN�%�j���^sЩY"O�3#�π��1\��|�"O� �J�aX@eh�/.�P���"O�]�"�Ð.�`�#���Z~xT �"O���g$ g��y�O�>�"Od�P4D�Y
�v!\�Af�#�"O���g�H&T,"u�M�J�j"O�B#� !)�^,V�m0��x3"Oα��l�$�6�Q/@�L!Ѕe"O���t�@�*��1Rn�i,thg"ON��FА'ij`cA�z��g"O�d�f釰?��x�K�� �bR"O $B�ȕ6qHvLȥ@�>.�90�"Ob��!�	�AW��ۂ�ŗ) 
��b"O�Ա�CH	�P��'7��)2�"OD��Ħ �;m$Hx�j�r'��r�"Ox� $�^�O���	[<�>L��'7�L�AK��ku�U�T�P���'i�X����O_�����,}9�i�'� ���/�?E�`l�~^��'�$X�1�4�y*�+T��T��'B����'=�̛G�ʿo�:��TO� S����{�
�Z�轟ԸA 5�` (�+X�n�#�-5D�8y��z����� 3�~1i�?'jn�#�*%�'a�M@a�A8��Su#�%Z�d��ȓ@��`S�S�v�8(r���`�4LKpَ3�4�"~Γ|Ѥ�2áW$G�R|��
"0@a�ȓok�홎hu@�i�}���؊��&g4�O���F�	M��ݫp�Q��@��'���xР�"-�UpS�E�;Ķ���hA�;."�kL6^@��'��b�+�
{Y��'���	�򄉞��z�K�#xQ�&8��խd~�|�a�|x�N�2"�!��ɞQ�⍨�)A>���W�E�+T�B�@��� 	Xx�A��"Ո��dX?n����h�1u�xh�֭I|!�$��]7�I�0�|R�j4A$Vo�`�uC�
`�ؑ��E)D�QB��O6��)Ckޚ�⑲�L��8ч�*lO~���b� �zD�3FV=9��c6 �u��J5D7P$�S� ~2�i
�S��" �<$�E��R)`FfM�=e��0!�����՘&h���
�R�N	;��8��D��EC�W����e"O^ #�M�]N�U�E+�KP*��f�@٨u蕄��[�<m�d%B<kZ(+��D��yi�m*��7��V�Z�%FS�yB�Q-1Ub���-K(y���lG}C�#��+ݼ��G*�:/�x8�W�qQ�B�%��p2Sm��a�����@��ɏ`��w���d[�/J� �~|��޾-���	�� m
��A���h���r��X�<Sb���53���3�����n*�Ĉ2�����n˱!l*��W*߱ƞ�	3�..��s)�q@Ԯ7��0�׹ ʴ�"O��6Ì0p���C�|���2f�йh;�PP�g۽u5$���k�(bV��&��4�O)aS��-\��E��	, 3���G� z��d����R�(C�f�P����� ���@�ߡ4�$�9��;����"L���j#"�d�$�BtB�9�֩X�炿j��x��	��ܱh��ýo��H)��M�n�S�K�#/����G�8&�L5�ĬG?!����bOH����@�Y,�0ۧ�Q����#%�䑲����D�Nt�%�
0x0�aZ�h3V擘5�����>�����R�l
�'G
$Q�x@�-����?T�("D@�q;���[!\�<�u�!BB(AO~R�B �y��^�X�R�;�yT��-���x2+H=S=(����R� � �pՠ~��#���:ij�Γ�ZH!��@H�Q;&�q��vVe2@�=ᮅ�� �X�����?䢝�E �]��x	�E�Z��i���7�IJ��07���
EhL�Y#�8�O��;�&؇����	_��x3w�|"i]��ds���9Vg�M8��I)��m����rE�� (���)G�z���`���9u�V�Z"O�x��k�&���G(�OIڽP2bO���A�눼�Vu��
$#�t�ћ���'&�n�85��4�t!��0����	�0#��^.><���Did󆉄!$�.�ʓ��#X�ZD�f �2j�\0
��î?(�ŋ%�:�@�"	&훣�S*<Hkϓ	}"��ӫ,l#�g��A�����H�����f��P�Yqf�<o��}Z1�и�0>���!2�\ؐGV�:�+���h̓V�<��A)}�\=b��ɇ	^~Q�+C:*�S?#3:hI���J�B�@�['fzB�ɭn�����CR'R��6cثD��ʖ�˩K?*iZP�ȯb5��z�,A�o�q�\-r�0�*91�E��sB�TB6�ףh��EJ�"OfݺAD��I������2hC`]!C�,Dfܹt�ڐ�P0�V�V�0�f٪a$�]�'�%��)�L�b
�lh��`RH��ZX���a��g�|IpTmU�}����g͘(ٴgׅE�^�k�g+�O�a�Qi�0���eQʐq����3��,���7e�)�eL�+ .�'a��@�C �-�r�8��<lTŅȓ)�x�#1nۨ�3ҁ�'Ks��"�G���p�?!�q�ǍA��y2��-%SȘ2�鈗,�Q�c�:�y��X
!�hG��|�ң�Kd(����s�r(rA�ǯ<Y�Q��hO���ш-�=�����t��#�e	��ō�0i���N�%�Nq���K&�໠�A�xR�ϛ0_\�׈��$�Vysd�J��<���Q<N�4�k���32�f�ڶD��^!��k������:�h1PQH�+��t��j���D�S��s&�@ĥ͂X����V�O�I^Tx��]ư��&��7���
��@�`@���u�%*��,W|�( C��I�@E�ȓn�Ԉ�f�Ε*�����$ŔJ�.���%�j�3 �rP8�	-]���ȓ��+��Zp�D�C�F��v�B��=RءxV�R�9Z<��]�T�<��HS�ԋ�fߚĦ�Y6͞2U� d�ȓkV\�Rt��E�v�"��G���ȓY�0�@d�X�Q��)�ȓw�2q+#N��z�
ʄH*^���W�`0!�=7�x����\�ȓ)S(��r̎�F�2{�胷k�p�ȓ`5��)�
j��[��l���0S��&e�(o_�r
�.a�r���}�v�هƜ����P�h�&�ȅȓ=�XQ�7уl<Z�"�e�]�ȓ��-��k�h`x�ƟX�Fń�!3̅
���~�U�ix���)
�ӊ��'����m�|�
�ȓrU��:r�_�dr�@�q�ʰ�ȓ:6~��P'���{����m�ȓF�\��b�T8�:��x�\ȆȓR��	P�'~��L2�'i3�Նȓ-���SsaL-B�8y�1�˒-��Ѕ�vZy#��@�Pd�QBb
mc�=�ȓ0��d��nD,{9����"WR�����]N�(4������DN {�&5�ȓSɮvg�$Qpzy��a�?,$�͇ȓrjf��&�QE�f	k�#Q�2n}�ȓ$��Q�N���`�r��H�nL|�ȓI��h2J�& .~�3Rd��f�ⴲ�-%	C�A�}�h�ȓ(
��[oҤ/��A��ʊ�_u�T�ȓ`��(�&&n [�,�L��ȓ_�r�ۥE�O��Ñ��<9��Y�ȓ=��m"a�!	���ѡ��s�vi�� r��ҫ$eA�����̈Fq���R�q2�� �t ���
3/����(����� %jG�}���N����+�ȭ�3�G�FN"u-i3p�Iץ%D�� �����k��<k5D�z�*t;Q"O��P )P2�f<�D�[�
�@��c"Ot�pƥ*?��4r�C��4��-�Q"O���C(K9R���׭K#N ��"O�=�o�)xP�}s`�$n�I"O�±Ǟ'�}fN�7	�� �"O�4��Fא$#Fڢ#�M;W"Ot8� �Z���i���Wr�D��"O���)*kvإkY�W{��"OX����ԖQ������U)i�0b"O"����Â}*�;��[p�`1�t"O�M�����l& ��ɗ>xFQkD"O�i���L���z��˴PVp��"O~�6�������#� �r͈"O��Seg�J��A�- 3��9�E"O\��g[f^11eN�'(��x��"O�MyN�^"�uA�@�y��Ѵ"O�q0)3L�|�s�"g6.<�c"O|�# �A� ]r�/� ��b"O��p���p���
��9;	��d"O���p-Y�m������s���"Od����Wl*Ј��P/Ma"O�q(�'��#�H�5��|��٨"O�"�N;p.�S���}�b"O�(y��ƴ*�dd�A�O�v��j�"O����8gH�$&��7����"OBxY�GA�p)"��\�;�
�h�"O�ź��BAX=Ka	"n�.�b"O�u��ψ*1�jPA�i� Ƅ��s"O���$��;��GG�b��pc�"O8��"a� 
8f��lY�:�� hV"O(y8Q\�Y�,�dk�Mw0�@�"ON}�	C<j���q�6 � �+�"O2��J/G��J��U�~<{q"Oz�{d���*��$��h��O�X�G"O�)�Ơ3y��E�V��>�-�v"O�(�X�!��l24����"O���O�1�����ϘV���[�"O�h��,X*7�BEAf���(�0�4"Om�Ь��u�R�Tm�Rc!Y�"O��HUB�/y��u������4���"O��U��2k0F��F��q"O�'bKH�}85ُu'jTas"O�Aa�˹8؂y�f�׮j�PI�&"OT� c�D��it�Z6׊�"OT=���Q:"��sn?���	�"O�i��@�-�0S�N�N��p��"OȂ�N�7?��
�.�5B�\�0�"O��e�ܹ"�����Ԏ�49(�"OB5�P#u؉�L;����"OF$�QH��@d����f�$�B"O���`ۊu�R,2w��m��K�"O|C���6�Z�P!�:���G"O YՠF=�Ts�Z�e�u��"Or�яP�Հ���;��5z�"O�=+�ј]ހ��#4#���"OB�(E�U�n�ۥ��Hd�V"O��K�E�`�zs��O~�4�D"O= Rc�A�����KI�.P*1w"O���@�
v����Lɣ7K�#t"Ofm�h��uU��2Gk�>���`"ObW큕�6��`�'E�S�"O��$�+�.J���^ӌ�ѕ"OX�3��̈́f����3�J=˺k�"O� 0hc��T�w#��:��O'��i�"Ol��F`T�>u��4�>�2i�t"O A�*�(l:��{�U:S؉c"O�+��#)���*C���w��l �"O�[ �@�O,>HQ#l�(D<�aX�"O����K�r��@�II /sи��"Obd�q.1_�8��H�;Ud�X"O:�ǅJ)'+���ƈ�hԥ�"O�pCB[�c5�I�t&I�>��'"O@����Yy͑r��
���e"ORг�a���b�
����Fu�4"O
H��C]6b)��ϯ�-Y�"O6D�r��;��A�X?x�:��s"Or���i��mN��A#mI2A� ���"O9 hR�nV�ݑL�%7�Ḁ"OR�֖� �`��έ?t~,c�"O�t�� ϲeul��k
�CSLa�1"O��01k�.K�n��@#z����"OJăG��:���g�#6~r�÷"O��p�dE?[���%�21\�I�"O����
Tr,�0 �|Ȱ�5"OĀ�w[�]K���Ӥ~�҄P"O|�4bߛQ���fO��^����"O�����\;���4�@L	"O��v�H�]��`PVa��}�앓�"O�H�1��"�9���Q�����R"OF�
�&F���a .���T���"O�`�y&�UHs���&�7"OV ����f/VM1���48{J�3r"O��F�L|$< #kS|f��s"Oh�"�̈́����ȥ�N�Sj��"O��@eˏ34
l��4Ꙓ'[&�"O���Dj�/p\0�'K��~\=i�"Oz�"��̝:�0��f,��|8�pp"O$HR�!��-A�����!
:,Q�"O,���iX�+D��#��O-y��w"Ob�E#J'~-� �8DB(�u"OΙBS�׻<+�MJDH�_K�]R�"ORŒ�ǠE� ku"(0Erp�"O��(�i
 T�<���ς
G���'ޘJF�
Q�$N�3)��:�'����ߦ 0�Hէu�|�P�'���æjBdٓ&^(kҰ�8�'\Vz�Sc�b�賢ۄa���'<hYi�kձl�^����VG*��	�'b���ũ�R3��@��$SEXX�	�'2\��7.`�	8�i��z��x
�'d�l�FI�&tDx�D��@��B�'��R�}�`���㘕T���h�'а�����+���G<Rb�2�'�r�a7	Y:N�P=y5��*�L�	�')!��U=��m"��3&3@��	�'~�#u�<C�J՛������)	�'�6I���0�`Ѕ�{L`���'q2eQtK6� �Wn�?}����'�:)���'<��Í�rv�(p	�'�2��S��h�89H��ٯv-!)�'n<0��gܐN�R�ɂ�ZH��	�':��w�vM�PQ��$ L0
�'�ܙ� U4�21 AO�y8�!	�'>¹I ��*+�h!	4�p��'�B(z��4�r���-y�V!��'��Hڨ@�ԙ�G!�4��'g�kT�l|��K���-r����� �P��%� !W���ѧj�zp9R"Oz���C�.V$4����c,���"OƬP"�RoN�s"�^(2���V"O|!��C�J�D�J`Ȇ�8�B��""O|)RDID"r{��J�B�xd�"O�W:0�p	�/Ťr�űC�^�<	���P-��;Ҍ�R�x�d�Y�<�Q��%ur��b��Mx�eAM�<�Ʉ<=� t�2�4X��ҧw�<ٴO��g����֥��/����Uj�<��J�X0�x��ؓq�.�3�nGk�<0�<w�d�c �ISN���}�<����EY���$	M'{r:������<�G\$j�h$�Dgբ�Y㮋B�<��iZ�Jl�H��/�eo��*��<)����@	t,^i
�lA�M�z�<�AH�<l[$p�Ɔ����Rf`�C�<!�$��cx4i���W�J�Q s�<������+Ү?�
�����w�<I���6/����J�9��5е��X�<!`ሠm�ⴘ���A@��W�<	���9$��q��/ލ*���X�{�<�DoZ5���`��l�\�@f	�p�<��&�.D@��8�o�퐑A��r�<A���?9��oH�v�ĩі*Dk�<�D�^=;�E�0J#m��-r��z�<� 쁠G��y�nT2@��D'S�<�2֨�z8�V��P��@��L�<9�B�6N:]�E�"�%�cgǉu6!�ăa2lI���CGd$�Y?!�d�+e����,F�( p�ԋ�1+!��2�n�b! 1O�]��k�� 	!�Z�G���愨��'Oէm�!�d��Y0��)t�ƙ)��U�n��!�$ڒ5��J��I�d*�*mʞ�!�dB�ء�Wh	U�SEż�!��^�Y-4�z���K�ܙ�&��$!��H@��e�N
OV�ເ�U�~1!�jt3P,��Wx=j�F�-�!�D,I�T�� F�Y�|ɠ�&>�!�Dà*����暮���4��1S�!�Գ%���'�G�f��	޳(�!�dȎ���C�L�g���V�
�!�A�ap䔊��|d�5:�ȃ�! !��L*uJP-@/�}��cF��7)!��?&���j��?KLT�K3ți�!�$?r>�̚�W"vUC�h�!�$֙�j(u��T����E6!����z)p6�v�NE�b�ϱN'!�$� B�h��L�N�&�Cc��G�!��߿X��!%�Q�4�[����#�!�$Z�z���C��9`�I��	/D+!��ԅnHv���J��h�8Q��(�#!��Ȱ)�"�ӆ �P��G��\�!���=x�b��D�ʻ"��Ձw��!��([TP���"Z�'��A�ү_5�!���*�� �T8�01mB�H�!��N���D+poX���!a�2�!�$L�cS4��nE���e���=#a�G$Ƥ�#ޑ<rv�iWN��I?lx�m"?þi�$c��yܧ�v�#�!̘o��Mb���v����`�x[����¹H����"�Ғf�`xU�P(��d��N�S�Oth�1�`�V$(WG^$=��io�&�ɰm�a��!$W��]��º\r����S"�'�T������ ��2Si�~u[hǛi͐=Rr�>�$�����O�aQ��1w�6;&�נq%���'���ä��Ӝs�4��d.ѰW��*3�G�O��1wn�
����&�8����f-���B�F2��ERO��u���	�w9�#�R,Z�^q�q��GOqO��0Q�-�)�)NB1����lَo�,��CW� @��]���Ta	;��Y�%ʷ<�j���@���~2�®iQ�O�>��HT�l"[��ºR���1��.)�F�����I��q��P�R�̰	V�)-ްT�&��Iu�0T�a��/�"b��s�Ar�Tmم���'���Jc���ԧͯ8��q�t$N�i7p9�0�9��	:�l��?���)Q�]�U��B��c�>��$�G?���R����h�2�Q���G��ʀ7~e� �!��EK*��?E�\X��Ǘ!]�-[A�Q~Dh_`��0���|§Ƒ����C%ܚT[QxܓnL�� ��O	�-Krܒ/�=%ph��,�9��{K��MO3,�j�KQ������⩟�+T�ٳtHS:j%�`I���y�,P�g�ұGL3c�"\�-"�y�S�SD�|;Q�0J��1��e��y�߉��	C��mT8�J�gP�yRgڄc�b���h�c���%K��y�Ü� Gl_"Vqb��#T��yҮ�H>���끍U��HU���y�3M8��"Sa�=V\��:Tc�y2$�i���&��=BLѣ�	 �yңN	[����B���a�9�y���9���R�%�;A(�S��Ç�y�Y�g(z[�7.��Є���y�nR>��]��h�25�4�Bs.�:�y"��*b��%-�&!C�퀉�yr(@0FZ�|�r�Y*B\�qj���y�.i:LjRχ�$h�g�)�y2j�&mR�uq��Q�B,��x�\B�'Z���U,��1�CB2`��Qq�'� �h�`�##:�$1 �O�0	�'@n�2�%yj8��P�E�Z�(��'�pQTLA�UZ�q!B� v�� �'^2t#g��35��%Ca�a��#�'b�xb$&
�!Ps�J�i� �I�'dX��n?C��x�Fʑa9|���'~�|y(A�7JJ��L�_|�J�'���ʠ��P���TZ@e��'��@u#¾D���X5�e��'�	(�\�IΈ���h8H�]��'�
��D��'�Fi���³=m�y{�'+�Y�M]M�έ��fӼ9x���'D��S����H�*M�B%�$7N�M��'�B|�_�ZD�l��+�3��0��' �xqk@I��1��4*r, ��'�j���J��0�]8��J9w��h�'�~3�	
H�8 �W��'#�ҙ��'�~�a ��@�{��o@Hq�	�'��ّ�C�����`�RP8	�'ze)cǙ\� d@L�z�����'!�q��L8R#.{���(l��'#@�3%+:Q L�� 5z>��i�''
 igj� q�h���ɑZ�d��'��+���s���Q��[�_/2ܙ	�';�����_3fI�L�YRL��'߾��P�\"'p�Y�lJPPXA�'Y�)��l�O��<�ҭ�D�P �'TIƧ�7
l!krI�bF�'"����OF_J��t�1ڂm��'�^��0�H"�`�t��6��l��� ��q��$x���s#��]>9H"Ol�CQ��?W�j��(�r|��P�"O������u/6|+�@Lq�q+u"O�yZ�" BlԐ��B�4����$"OR�8�NO��Cd��\W"O��b4kL8 �Yyp�?��eQb"O���@*��\$���"O��@��"O4@ٖ��r���2b�D=���y�"O�0K!)��U�p� ���#�~x2�"O<s�j�<��2a`�9::A"P"O�s�c���@qXE ˝&!�ɘ�"O(�!�ͣP���r�BF0�"O�ٺt
_�D��@�,�)H�6"OD��UHҦ%�ܙ�b�Ș�"O�L	��y{=�蟥z�t�"O�	J�c�,>!2��d���(���v"O��R���
`�qKT�(�"O���5n�H/�1b�*�rV<Y�"O83.3j��l�gP�|��"O�PH��>m�M�sO�#�ҴrG"O�(1��!��J��.����"O�����d0��G�ݭNVb��"Ohd"0CԌT�z�C�j33���q"O�;��)(f�M	��U3XJ�5"OR������h~b0b)����R�"O��`O�R�KΚu���Y%��"�y� ��c�ʠA�%%Y�z���Q��y���;g���#��O��d���;�y�K*"�D�"�A'�d�q�$[�y�hF�D(��K?���X�DƓ�y2ί5�&m���eŌ3G�C�DB�	1=���1Uc#���`Dǂ'6�tB�ɡK24��6�^Y:��끤�>B�2��B0�ܸ`3&�59zDB�	-W����V"n��X��52&B�I�`�h��� �'`�( ��U��B��S � Q�%�.� |ٗ	�1w�XC�I�/'��Bs���G��s�\3 f�C�I E׸��C��%n�1�c�Y,�C�mGr%5LN.*�	!X�r�C�"�0���̀'1 q1�F�R�DC�$���(�"�=+���7C�B��B�#p~�q��N�p'�|�7���.,�C�ɪ	�f�wS?v�܈�Q�!�^C��0	���q�=o��sC��%Z�B�IW�ns��Ǜ:nD�'�ƹnvC䉜,��Y`I���F��"c�0B��6.���A@9%ܬc�h��E�\B�I�8F♲��G�T|qR��`�"B�	�w�>M�N�5�2��s.�2��C�I�)orѐ� 
�r�ܨAX,{�B��3pF��R�K���B��BB����IS�Ņ�>�i�go��^��C�I@6���B���1]����ʃ*$�nB䉩A����p	Y�~�&a��o�	^76B�I-��<*׀r���"�g��}� B䉚@x���c��9����p-�C��3����l*&`J�)J'B��C�ɂ|�t<�@⏁b��3�mʥ8�C䉫K�ju
�B�8�X0���&OC�C�����8��;rNܺ�䝧L��C�I�G�`�a�,��$�P�r���U�B�"-:�W��/òDQ��/-��C�	�iƄA�l�lܑ�C�)� �)��IH!�\��H�̀@��"O����A�P�bl¦\MN�{Q"O �A�W���zԫ�_D���"O�I٣�#f�$�����-�R"OPճw��{��!PIF�T��&"OpL�Ӎ*B�D#�'�_����"ON��Ӎ�GD��GF�)�y��"O&��N�)�ҽ��ʧz��"O����ƛ 	LjA$[�,�Z�t"O�h�g�=E��l0t#�|�R�s"Oz9�/�"g���)�KT�d�8�"O*%����v������D�f+��j�"O98#�ъ9S���!`��r"O�]��Ϙ+�ͣ�`I�x�}��=D���0�ܖ�0�Q#�/GՀ���g<D�T���e��Tw��/+�b9D��D���U��AC�Cڲ�<���5D� ��1_�1�1���nXÄ!&D�� AfX?B J7-��D5�1���H�<��V�x�f�iF��'�<!�_[�<qCgH-�:�P���4+<�����V�<�vMӂnf <�rÖ�=N��G�G�<�G'Y�]Y��ì
Q�ůIE�<tj�q�>y�CJ&$0� 36�Ly�<!��7�:uX�/�x)F�Z�-Ev�<	�`V8ck�U����i+D�$��L�<q�	W�R��[�z��q/Go�<yt+H8^%(f~A��K��Ih��?�S�����'����3�ܶ^�D�ȓiո̠Ǭ��*���{@��	�L�ȓ<@L�ƍ� ,BAN�!��%��ZI�yc�k'~�`� ��8�ȓC9�R�.
�z4 aǄJ�.xn��U�bi�a�_��J8�ƬM5��@��tT����G�PQۤ�Y�+�6A�ȓ]ޢ����J3�e�Ů���t���l�h��8���3mP��E��v�1��܃OeLDQ��L1������;������o�Ȃنȓ>��<h���vϨ��#�P fBՆȓ�r8���̦!���jR���=☆ȓaK����&2�$�j$�E!	��Ԇ�}i�X�7�T�O�������(/vf%��K�%�"/I�|I�Ŋ��D&x-���ȓ8�ԭ��"o�⍂3E�x�����\����$B��5��b�k\,&�d�ȓ�4ݠ�;�БZp,êG�T�ȓ}��2(���9B�@B�dOV��ȓ;^u��& �Ze�t���ȓ��IQQ��?{��u�b�<�@<�ȓM�^I�c��[�{gc�~�:��ȓFx]pB�Z�3��Z`���⁆�7?��C�Fv
6$��-RG��u�ȓ�P�I7����b&S?F�1�ȓ$I��AB͜3���A�_�XˆQ��L�$��6��40���9��I+;�F=�ȓ��H�哊(2�4!jb�p�=D���\bH% 0�8�䭐l9D��R�ī�����U�Q��H$+D�Dw'Q
D��B�8�0,�7J(D�T��l�:U���[�%�/�PJ'�%D�\�R��MQ��bGZ?SO[�9D��j�W�x謈@iV�,�ȩ�6�5D��; �_%,�D(��	��zҨ�g�1D�� ��y��:d_ �`�NH����b�"On�0���!S��+�'��`)�07"O�0�n_�h��J���4L�� "OD���$�6o;>a�d�1e��"OD ��c�%��i�)��1!�"O8M@%�A�KԹ���.�̠q�"O���C���8��f�#;u���V"O�i����0L�1�F��d���"Ox�1�FA
D4����׶m�v1s�"O�h�&!"b��c��Y�f��2"O,=�!$!=���;���Nv�qc"O�x���Nz�I�a�J��9C"O�z#(W)qM�i��χ�N0�f"O*����9 t���6��djW"O�����,A��!�� ���2�"OhT�O>~tZ�8�/;<g,L��"O������9:a�[�Z}Ib"O8� ��\+_T�����^h��"On��I[=�H�	�d�-膸�"O�zD� #�"�#y��Pf��*M�!�$ݙ5�ҕ�d�L��@��3!��ƼgY�u4 ��c'f���L�3B�!�$�x�   �