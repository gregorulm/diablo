MPQ    l�3    h�  h                                                                                 S�Z=��(Y�����mB z0�Q�`�;��lR,~�ḌZn��\�J�����I�m����̅ ;��u�15������.gut�Ȭ�Ź(���Sd���?N7��~�?"�1�`EE^���0y�ƅf۸�O%�d��eAMHk�����sU��)�"��0}Yr��V�Oڝ}�|��Z*�j�0MP�AO���}ɨ��rs�
����=��Z� ��.���]�a8�_��v�N
��0sYԭ{Q�ųm�#C/	�?���>��VF�����E���"o(�`8H���,�QF�w4�7*ץa��V�QR�X+�8h�aH���t,(�.�$t�����
�����s\ղ4�U�T�޻�fѶ��x�S3{�Jf�~2����"\*
fj�hb��v��X�CpEO������!D�8�a̪�o-�mCR]d�kV� �iVQ-��u@2�<���Ev>����E��+�<�V��7"P�Q�Z��@fM��4�24?�����J�d�y�a:��@
f�Z'25܉T�q��Ơ�%�4����𪡵����g���E&�R
�
�w�!�bD&��=fM�1U���0�ͧ{p~�'�!�5�Ik��gI�mm)��U �hA�Am.��R���(�� ����	�eP�2t9F���&+.��I��[n�U�V����5���P�����\��� ��B�|��z�j�m��ٰ����j�����4�ďP��ᜊ�Ͳ=���g+
�)�4f rR�����-�3�P���e^'��������v=������e��T�ְR)_Uj��;��)��){M���ÒP�֖�`L˹b��l��ݱ����"�>�(�@�����`�gΙ�6b�tBB�5��N�h���ٝ'�,�*�6vB�hw��%�wE�wS�k���`�8���:�^$�7���P#�#wr0K��F�p��(�\�?���a�L�AM���/&u�Y�!u�y��Wa��&E\��`O��I+�^tzIC�8X��<z�Lţ׽a9�op,�R�Sp8�vԀH���f���*$��|��$��P71�l�M�#�����"��)�4��'�����R�#[<BI�b��y����s�9�
|H=e����^"
 �ȓ�J����B�]�3|�TX\����	��v%�N������=�sP8�
��ohی�V*���m�r��J'u����:� V����w�6�Ǆ�m�k�Z�-�������c,�/���4�r��~�)�%CL�pS^�&c�+@�8��p5gN�2��!�D����d(M��	�RA�v+Iv�E��];О� C`����n �䬧*Bف�<�6��]��h7dJ-pb0��z�!*��	�	L��\�~ڴB��Fp�}�r��8%�*��:eП��N3���A{��8�I5Pw��WFk�-�mim���T^شl��XحZ��<wI:�#�R��Ô�<����9cPbm�#��p3_HFzJ�Y4�ٛ��6:�Љ�&o���څ?�JOm��ޥ@\;ߴK�6|��i��{�T���/+��*oC�l]_�;L#J���sH��o �ި"�d>���q��؀	�����Ζ׮�X�5x���S'����X�4�،��((��A�]V����w�� �B��D<~7�RP�tb>� ߬��g��� �­'�I:0CXJ@��.��n��066�����t�D�ۜ���#du����ի@��5`f�-����u�r���[R�[�:�F�@ƪ��=�X�t�Z(�!�VX0�8H����F�"2��{�&��%�f�n��F�<{U���~�v�$r���z�,�g	H������;o畺+�o0�/G�Ъ����G-���O]�"�]�Y�v����t�.ొ�S�騯�G�~�CK��n=��%�[dSɵ���2+tόvrW�ъ�vF������D������$�|I�VY���/�5�4s�����<[�^rn��b�Q�{�+�攇<�(V��*����o�n'����˦��nwL,MJJO�b���C����ڇs�Qz�d����HeX�HZ0�#QΩ������g6���Y%�MC@�_��.7[#l�m�(~`F���yK�����$�gP"O�:�|�ϼo��+K�d��	X�X0��2����u�y�OC���|r"��X�{h'�n���7���,�D�t���eL��RQ���m	*���sy�V�1��T�
G�r�#�1r��T0��y���
�ڽЭY��hw����.0~_hp@	 ��*�L��ޔ�#ʠ!t����5)�gEC�]�r
��fI���,]��g��J��Jq��4�e�YtR�O��3E1��@�ƾ��Vn~e����=�B�
��OT��߉TL� Φ��h9*��h���^�~������ %�C�ӎ�]"0������.�z���Qm��Y	�Q�q���-��.�����3cj�����ڠ���E$\!9�����������t5d���t��@�@+��C�p��G{��Kɸov|��E�7sE{��V ����n�>��rC��r+;��n���@f��C�#�F�<�_~��ϱM �� M0\�Z��r6������|�.���lS��Jh�-�j������,�,Ȋ:�F}7�ʀY��E�
Ao{�Y>��o|Q���%g`V�����z��4���2�ffJa�m�D7��(�[�c����h�<*@�/�B?׫����
�k�#��1'+��f�x��� 8�G[_�S3T�p'��O.���aS'7}�43�^
.��"�jsd�hZW�|3�/�{6�@�� �;q�a͙�3i�Z�x��o���0�`P���m�C�m�,�������X9�RLUF����#m�mJ����><hז/W�FZ�Zb�G�{���*�f��,�Aލ PmRΰK�fo/(5������2��X�#�"\]��ժ�y-� ��� C���0�͆������=:2Q g������!���}��a��(ᙦ|�_>�� 8�s���*3��K���Xv4���������2XI�9gY���\�I����J��I�
H���u����梮�1Uj2=�Ѣ� �~PlP&�a�iK��~�*�GvF�)����*�Ԏ%�����sݳp�l��pj]:�����Y��y�H�͇V�F���~'x��Qz^Z-��״.ؗX�V,��[Vܰ���#��2ʷNI�����B	{fY�U�m��=�D�2�B�5AZ
G���d��^�kY_W�MS(x�h�PփRDx��U����`q�.I�ƺ�����e
�WBzE&T��dr᜼cis>�AZq$}w��D^��%�2mb�t�[�gc�C��v�\�5P��q(7��*�݂,(y��$�1����!3�`Cz�⭗/Z���fA�<�플���L�I��ei0��\Fy�+
���L��?����kljs��(z?E d�'�@��E]�Q)�`
U����v�98Y��gXz�PցIV/�l�s��$��!���==-�9��z��J�$aj�m�(�,�7B�� t\|ؘDB�m���i)?_�8�O����DNp�f����ߡ<ͮ��Y�ӹD�M0�x���x����b���QL����6!���P?�ؓ ��u����bv�Ei�e�m��p��6�&�n
���[�T��f��+�YQ7ֿ��H4�Ol��f�|O�z��H���m9ǖ<��N���(e��{L�%�U=���٢�M��O�f����}�f�3&p��	��^��������v8�>�.��� �T FmR���j�?Ь��Q�7�c{H����Ȉ��g`g%�b~��H��������>�'֛#[��B9˥6gI�6=�7t}���PwN�ہ���h,��`*<jBf��#Iw�BS	��]3U`�J�8��h:��틅�&ZZ����+Ki�2
�pB���w��?�_E�Z�LV+�)s�&�XY>u�3���ܝ��0\޾�O���+�8Yz�\e8͜��(�>��~&at-p�P��N��FH�ނ�,����"���`$�|������N1���M~~n�W#ڃ���N4�N�'J3����R��'��}�|��;��y�"9�UrH���z�n^x� >������8Sn���n�_T�y��d�	��%X��#f[�3�Q�N���k�
��ۇ5*J���(����bU��k{u|��(�s �͞��	6'���~�k�`@ǘ�C�x՛�$0�,d�ணl� ���9���@w���
���?�ﭱ��t��k2B��m�bI��_��g�M�Q�鍥��`�v��$��Yl�C{ /� 3nۛ����n�x��7@*�PG�#u(de"b�*z�ɧ����VE�WN��"���p�]�r$�E%�r����8�:;N.�&��=���oPJAwp�aFF�}��"��]ћ^Ө��&�Y�t�<���:s�R�5�#d�}.�cK!ֲ~Sp�n�Ha��JD���q	��k@�&z�/�c�i��z�,�WO�I��f\v�Ĵ�/�6w؛iE��aǦiC+(*J�glIB�_^��;GC&����H@�� �@�"l
���`�q�i�������\�2�3X?�,�<�'h���34L��w,7#g�AlT8]:��_�\�9Dw&7G �KL7bt� �XK������!��^�IuA?X�x�)A%n	�0�ly��|���ζ��* Od_i������5���H�(������ ��8j,�V԰:�g���G��c���V�5!�r0.�����HF�n����{������A����<�_w�����<R-����H���Ȳ�<����0
J�js����e�����Ϫ1G]p\��E�ˆ���ϝ��lS�y@��F~�F���yZ��V= ����F6�t��rҰ��$Y�0i��1������� �@��
�q�e�[Y�5��W�6g@��V2^m�����6(3+�7m��YVo�[��rX�
+�n"8@�WE�h�LG�J�]�b�p�~3�:�gs�VT¿4ĀQx�X&ܝZ����	��-6�8��6��δ�ߐ�T��__��.`l�2��%�F���y��R��)�$�d"ʥd:��3|�z$oKވK�ʛ�f.�XӦ�0��82���PL_���?��3$mS4���h����.7(��2�D�58��Ny��Q�-�m���2��� ?��]T2׉Gdƙ#
��r��0].�S?
ct���	�Y@b�h�����0~�9�@�d�3��ǧK�o����tM=����)\��E�`�ԍ�~��f����@,�����^�E�5J����r�t���X��{w1��]@�����V�����t�XT��^�*\���L�DΡyOö@���
������h�/����ӉQ"��N�����I�:(�my8/	�j̟�(�".�w���c�>�N�������8�}$��u����1�������6����{Z��޲���1��Qu9�*��&�e��z�E��t�:��n�����șR�;��ڗ�'f���^8��ם�~�5�����۷�\��ZA�Rr������c΃)�� ��Ԧ�h�j2�g���g��%�RFxM<�%V ��Ƅ���o�$>>���|�	k���V��R�'�5��4�+�2qM�J<UČ��X��[���)h���@���B���(��Ei(���,���T�%x�W�;�G���f_�T��M��IG.�+�a���}��PNR
�r"o!Hd��W�eZ3�<����J@@�0�j�Jt�t�i+�*x_o��}َ��CP��/È��e��H&�, ����T���*9=URU ���(����+����<���/��9U	nZ�<�%������(�AL.P��Ϋ�f�sl(јt�ݻ���Zk�3��F��\�M��ЮԑV-s�����0f���PA��K����2�����/G��gʁ��}�%���(��8�wJ�>�� � �s:(ϥR�&�sܓ`s4������r�C�織T�ے�d�7N����M߫�ڻD�.
���ȝ�s����)i�UE���� r�~Kg
`����@K��)���^v!� �鲾�iώ N6���n�ol�Hj؅킊��Ĕ�e������:_�w:�x�z���-������2�tV's��1�N�#�2��~N$*9�G��ݼ%fTW�ȗ����D�;RB8b#Z�ʜJ���}�kTQ!���0xY��P-�]R����6}� .���e.��!ʈ�����ZW�<�&/�{d�.���]�>�Ɇq5������H���2H5t�Rg�=~C� =��F�PC�(RKl*Qao�]�0y6C:�̲g���|`�˴��M#/�0��AT�<�c�'��5eI>��e$D��w�����
��8L�)�?l���j��(5޷ ��z'� ��QT�[`�`��� v��8A���lT���\'����lX����!�=��C�T3�ʇI�%�:$����'�OB�1 /��س{���č�c-)z�8��ֶ��3NbO�f猃����Ѯ���j�D�Z�sc���upX(�9o�������qܷ�s���	�M4�0�G��Zu��d�e����3o����w�&����V;[�7{�LOن�A�Ĕ"z�����T�Ѫ���!b|&�z�m6�#y>�OI��1|E��%��B�U�:s��54D��fD=�C����e�_f��S�g� �!'�3Aj����^ݸ �"����v3M�����۰�TձR$vj�u�5㎟�R@{C�A�y�`�L�`��b�;�|�B����X��>
�����v�����
�gĊ,6�t���k�N��z�p�����3,/�*���BA��#B(w{�S�����g`f�8�4:x{��f�/�a�%�Y��&�����Sp�JK㒳�?I�[s�LV����.�&�HY_4ug��uWҷ�v�\��O,�i+�2�z���8�4�|p���Y�Ta�c�pb��I��,}Hw���G�c\����$�f|%����P1Vk!M9�E�))������~�4��'嚉��RNx�-5�=�o�6�T3�9��Hs�9�u� ^��W �˓{��H���M��H�T��6�U�	U G%.�>�Ȳ��q�)�������ۂ��*�*W��*�����w��uWeFc3
 ��5��et6�t;���#k��n�&?�S��_ǰ,���X��[u���C��[�2�f��܈�*P�n^ֳfO�E���:�zǚ��"Mb�H��RX���Gv���9�?�C�*��{�n����{x89�2�ٹjb���Ґd�7�b&� z��u�@p��?���R�+�j_��_�_p�]�r��>%u���6���զ|N)-���+;��Vk5:w�xF!�]��������^μΑ�_{��r�<�Ց:�6VRZnW�^徇�pcF {���p��KH|gJ�,��c������)&u�վ�kĀP���G�Oc�Y��|\�឴�q�6rM�i�\�ʻ��=0���*%�0l�G�_�@�;B���P�SH�)\ 	�"��ղ՜q*�.�?����𦖍c�X��%�,��'����7�4�Ċ��=MA���]�E���ꕷ���D�.B7�]F��bϞ� U$6��5��O���I�r�X�Ѣ�$��nd��0���Bs�j��Α�e<.d�"0��#���G5֨3�c̍�u����+�2#Ә^�Q�(:V�(����:���N����*!>ۀ0�K���p4FC��f�{�$�������J�<Ld1�����,ԟ�|���"��]$���	��%���y �e�&��� �E�߱:���
]K�2�Ӏ�����ҷ*���'��S*�����~�i3�8K*���Q6��k	��Z}t�rM�K�����k���HG���'�{>����.��E@�֢�5���q�c�rr�^hl`�S���a,+���2�9VJ�\�.~쥱zn�J���q�#ؤLb�$JE=Kb�?���՝�s�{���ހ�GXA#{Z&7Y�$U����N�6����˺��؍�_�`�.�El,��^�F�D�y��M��$ǁ�"Ef�:���|F�o��K�Pw��sFX���0��2~��+Ǵ���D�<��h�Ǧ��h��A�1�I7�~w�XLD2a�W���QX�4m��3M�L�x�e�TmñG�9�#��rpF60����
�`�����Y{Y�h�����r�~+v@9��Nr1B�V�J�@��t�F���)��E��Ԩ(��\���n�,�� ���@�tJ'	��٣��hY�E& ����19@&(���؆V$C�iS��s�=�����U��L�AΜW�T]����%cêts�®;"A]��H$ӄ��"�S!�C|ոd^����$mT��	��"�,\�#mk.;k�Z~�c�R��� ����s0j$��ꦐV�ٌ1w�D�T��Wʂ�����d�ܶ�>�y���;�������?K�A��-
E�X0�̔2�/7jn��:Z;��TR;եΗ���f��Ϥ��Y�r��~��6�?�͖B�\7��Z��r�F�4k����r�$T��{�T���zh&�j�XBw[��������Fs�<ހK�Vgj[�oq�>f��|ǏX�[�V�ٺ�����D4���2�S�J+���9��y�[��l�RT�hA�!@,�B5Z��ĩ����Y��'5 ��3Ax`U��V
�GQx�A�T��H�Lؖ.���a	J2}R�ri��
$Z�"J�dH�%W<_�3�i��1�@�@E�'Ŧ��O��if��x�j��u]��FPr��ãK�9�=�#S�,;cS�E$��X�9�w�U����NU�c������<�]�/�"P��Z���x3����\���CAT*�P�}�Φ�sf%�)(������(�����t�\F^s���X/5H-.�E���꺫���^�|��[a����2}���Ɂ�	T����}}�J��(T�/�r�>l�E �%}sU��� �ʞ���j�4O��L�����.�o����B�(��!ֹ�F�ɻ?/�
���X�����>�U *�G�d 5�~F���$=��g[K�k�� Bv��g�$��`���4[�t���)�el,@	jS�euS���;����������
2�2�x+6�zT��-˚��MO��	V"��-��	{�#'�(�qN�Z���f��x�fOK��#�򵳥AD�d[B��QZ�����bw� �8kOcG��xB�PHޟRS~���[�#���z.�X�p���C����W8�&
.d�y��r�>�qOqګ�EJ_��-�j2#��tC,g���C㓿��P��(m �*�٘�8�yqƣ�g�������`�tS��/P�o��S<VN��:K�>,I�!�e�w���|򊺱
�e#L	�	?-��j)lW(�� �������N�Q�Q�`@���心vF68ϊr���pĭ�7[K�m@l��K!`�0=��>�o���9� ��$׾�����"�BHgL ��b�����c���� )��8!	���ؾN�N�!�׃*�ߗ'��Z#��I:�D,�;�n.1�.,+Σ�T����ߺ{|����3���Ο�o����N�s\�;�de������
�0����&<O�z�([�:�ǵX��wT��mm�I�ʀ �����&�|A�z
���Y�ԊE�������^���g�P��c=t�@��Q��sf�W^�¯c��SS3\ؒ���^��j�]�R��7�v.�?��(ŖhT6�~R���j��)�p ��m�{>(O��8���`�9DbEWB��V�\����>�Y�QҘF����g?�"6�#^t�M��fpN�����.��X+c,3��*21�B���^�{w��S[ʢ��`!��8�:�9��A�݉�̄��h!3����zp��R��~?�RU6��L���_
�&uY�L�u"+8�p�&�Zx\T]�O�~+�L7zZ�8C�MO�8�]��4$�a�̓p����D�����H2�j�b���|� �$7�*|����� R1�gM��A�DY�y/�Yx4R/O'�"
��ER�R�mS�v����/��9@L[Hݩ�p*o^.Ҏ ���C�.�������:T)��fm	�0�%�i̴Y�>�)����X���@b��}��* �k��e� ^���u2�~��T '�՞�6����=k�R�ǎ҆�.-FԚ~�,�������&��� 9�v?B�����o��eq�	hh�a�l_!����И�m*���M=U � �G)+v������1�C�tk��-�n��۬XS���-�E�Ŕ�ՙP=d�l�b���zry��{S|���ۋMjL�ż�� p~Zr�#%Pxv�q�<�p\�N$��R���i�H�@;wft�F�	΄�ܓ�q^��)��=����<�ˍ:i��R5W)���͇�%`cA�[�4��pd�hH�H�J:�j�/��&���&pm׾u���g�bN5O�=�o�\��l��F6m�i�8̅�{J��~9@�* �	l�l�_�z;=㲊�S�H�t $eQ"b��Սj�qe�'���������X�Vb�G6�'^"���v�4��a��Q�3�A"��]��&�9���3z���D�t�7}�A��b*� ���k����(��iI���XJQ�9n���0g:��4������l�7���dF/��z�Qݍ5��@�~;��`%ڭ�#� n���L��:�
��q,�U����*`��:!yM�0dҮ�]�F�gb!){)��u����3m�^�<爃��Qn�����_��a̲����`tk�f	��`Y�@�W��Ө��m�	"�]&l������� }��[��THS&�'�b~��ϼs�N�qf�LO���AM弝�t ^er�͚�{�.̦���g�|i��֡Y�M����B�Q5i�0Ѭ�;���^c��s�󸬻�++:�����V%.�i�w�@X�n�����޼�L}a�J�<bn.Ƥ���p��s��|�u����7�X\��Z��k����R���n˛6���jڵ�~��8L_U�Z.�ɞlg����qF�&y\&���$��"�F�:ix�|J1�o�c�K��.���XI��02�b�bz� ƽ�׎[cW�ithX4q�L�l7��s��Dm���"Q��~m:>F�N��ǃ�lV�T�ύG��# ��r�,G0�q���
Ym�a!Y�p�hH�j��DF~p<I@:v�iF�6��%z{�Ft��U����)KEt�����׋��v`�,p��H�;`PJ�pAe,��Y����Ĕl1tP�@�g����V՗$1��^g�|SJ���y���<LT�ΗUGy�c�@�Ѫ���.�|�p��#[�ö"A<t��o���m�0��m/T�	:��B�0��.�~
���c��(�D�4��T�̮�
$-�������o�����Ř�]���X�����@���e��(���Ԉ�\�ݒ��E����R���xn½!�ϓ�r�;�J�~�fnI���"��_~�dԱ^�5�Q��\R�oZ7V�r�vҴo���Mrσߴ���5�J�xhA��j(�}��
�[�2Fn���`n�(�-3o��>AB(|6���O;V����Tӥ�54瑼2gz�J� "�����R�[{�󪭿Qh�`@.ڹB��n��J������["�D�
�x�/�q��G�4g�2T8f��>.��ad�}�x�q
�a"%��d�yW�x~3߶D����@��]#)O@���**Bi��~x��5�ݍ}�A�iP-�þ����O���$,vKB����;9�Uw��(�u�ޣ��_y <Q�/(}�KE�Zs�|x������	O��MA�(�P>CPΡV�f��g(G�ћ����7���4��}�\�v������-�,�����&��ҢW��������
�2bk��A���$E��w��}XM5��(�~�m��>�q ijsp�Mϛ����-��	�4�<��8H�(_$cg���\y�v�.��!<�\:��P�:�W
Y�0�&̠1B��4mU����� �|�~A��(ؒM�K�٧�F�v�"��_)m��L�:\�υ���b�lGȱj�|t�@p>�
$��J�����W�����xF��z�}y-�@~Ɉx=�h��V���lHy��#BCq�ΐNګ������#fJ��~��n��D��B.�Z�ډ���>���kJ�ɺ^G�x�ޓPcJR�
Yd��� �1n.�~��9������OW�!'&�`�d#)��4��>�9�q5s� �٥���2���t~�g4]�C�&��m�P�$3(��*Gr���1y�ia��s�Sr�2+�`@=V�3��/��G���'<�Ĭ�]��g�I�i�e�����Gt��
ic�LD|�?�Iz�aj�߃(�{� �J�Mֵ��tQ�`��R��~7v��a8�����%�����=�l�7f�զ!��V=<�̊+��}H��۱�$��>�d�o�B�[g �{���I���2鍡��)�n8��)����Nn���F�E����ޮ5x��*�D����i
��O"�cc�o鴢��ۺV|���������U���ئ���&�+���et;G�%�yĎ�Y�&����5��[�]��B<�`�P�
%� ���̐�`n�]d|\�z����Zz��a?�g� �}3���w�����k��=O{��S�8f�9��Ѧ����3w�#�zn�^�FŜ����P�*v)���?u �Q@&TQS�Ri�jd�=E���{9���/���a�`��b~�2�g���\���> 1�֬�m���5g���6�{it.�"̡ �N��N�&�����,N/�*��?B��r���Bw��sS�3�n�`��N8h:n��/��5x���c�l�CBpsH���_�?|�L�R���&	q�Y�`u� kSE�M���^�\���Obw�+Ɇ0z�h&8�*}j�\fs�ӫa%Xp�e��?��⥖H��}�[R���[zc$rq\|[�$���=1��M�Na�_-p����4}*4���'�B�0�RM�(�1����e���
sH9{�MH����k��^��% o�^�:+冀¾�s���VTĒc��O	�%����t�����ߧ��O���J��x�*[ �Yة�;=�m��u�g٫S �/�����68����s�k����	��	�S��UN,5jS��\:��Z�j���ӹ�\�}��vv���פ�r�\�����k����}.MM��>��⽦v�%�:GЊD�C�ޅ�q�8nlR9��K��ц(�m� ���T�-d���b�rzM���V��u6�H(I� :S��)Dp-�r�/�%++p���l�2�Nx�\��$���kDw��F�g΄Y%�.3^�D��7枭F�r<��:��wR`�����Nчc<y���plIH�I�J�+T�E���"7{�<$�&kW5�t�����}:�OY��Jay\'6/��TP6h��iV�<�@[��U���*۪�l���_/��;8cc�ӴHq�� ?'/"ݺ��hq�/U�u,���fo�C��XpL��b�!'�rU����4�Z��HsIOA}t]B'��T���)���D(��7I�<�gb�> �������u���I&5�X����n�0"Ѫ�O���`��G`�	d�	f����3�5L�ę^0�k��ڈ�^!�	V��G:-:���,�t�p8F�D��C:!��y0�ޚ�~j�F���>D{D#��𮼦ҕ7����<��m��)���b�^����6��S�P�k���}����[����ЖO���h����]$��I��P�݆���*��-�SA�w��Ul~eܼ���+��G�o�!�5�w�t;9�rC��V����d��
��wm�1%V�w��±m�̕�5DX%����	�^^���Ώ��g5k+F릇(w{V eϔ��E��6n�s�hq����bL���J;\)bI=��/����s�%�������:Xw�Z�	�x�����	h�6���	ѐ9�kS��_Ы�.�.(l���Ĕ��F�]y��Օú|$��";G�:D��|�<ToְKǼw^�X�t04SJ2te����;ܪ�rl�^����qh�$�g��7���NED�9o�UȐ�~#Q`hm��k�i,��BepGg�T��G5��#���r&30�C���
ԙƽ<�nY�Ah�[��6[~�m�@����:S8��� ~����tz���i)m��E/�����0�RN��Qrw,Ih�Vz��6��J��� �r��� �;!���Q/1��@\�
�}^�Vڇ��.���Y���r��3���V�L��Βs���q�%�[�Ȫj�b�dA��r�~Y��z��"�DGใ���T$���(m
	uv	�M��P.��ЛQc�Z����~���_$ȏ|��4��B�c���Ԅ��P�����lp�,��ϯ���Ư��b�ʸ[���w6�#�qE}�w�B�e�e��n�҄�Y�ʱ;�N���$fI���ȼ��#�~�D��ݫ��\m��Z���r������٧�)��`�1�V�H�h\�^j������٦��gFiO��6�5��bH+xog�t>��|=��ԑ��V�;�8�;�f�4u�2��J�6)�0��)K�[vӖ�KVh�W�@I�B+]]�zޑ�����eO�Ŷe��x�8B�\^GG!�B(TsM���U>.���a��}ȧb���
��" gd�q�Wr��3�#R��{@qPz>���kO��i܏Fx0�����9��ڬP������/>���,�Se�{#J�>9N�U2��C�]�Y���:��<Td/��#F�Z΄�3�{�:j/�R]���7A�FP�(�Μ�Lf�<%(�F�.���d�Ģ���\|ߑ��zG��-�{~���2����}p��+���9�2�yj��\C�?V���ɍ}3�Z�(��%�h�f>"?| $�}s���q������D�K4�!�����ÔW$��C���c���;��`��||o�5/V
��Π��L���I�Uօ��c� C�~<7qyT�MS]K��ܧ�lv��洚�B��ώ`9�*k:ݟ�~lbpBjI(����E�D��묓��A�X��-�xa<�zJtd-�������;�VG��ǃ���"#]�L�N�C��^0䮗vfE9Ù�j��)��D'FB���Zv�!��pڏV��kE秺�؉x��NP~f\R�b4+��Ѵ��W.�� �&�z��fS��F�W.D5&���d^֦����>�!�q�Z.�������zs2�t�|9g�>C������Pt��(�*�*�*P��*y�,s��ҽ����hv`�%��N�6/F���Ll<̒��E�Ű�IO�YeU?���2��7h
D��LUS?P�u��j�rP(fz� � 2��ﵱ��Q��`vC���]'v�rM8E~u��O�fm;��"�B,�l)���!j\=���̥����wd��-$M�a�i��B�o� `Z����Y�M�|a�)+��8WB7��8�Ns�
�ڃ`�ߍ����:&Db�'�d$���X�g��V/�xӣ�1�X�"���i�t��+�%���a���A�1�eO5Y��@gP����&� ��Y�[��p���{�;C��EV�x4��8=ѻY��R��|wG7z ⩒�{ � ���g��xj��S¨�k�J��܊��=*G�َO��0JUf�;��x��R�3������^n������J�v$T1���0�8DTlB�R�;Bj?Ĭ暾�� g{48>ʊG�}�`�͓b�3��B��`��)��>��|�mI����7��g5ds6���ti��<��N����鹝�<�,iߚ*(x�B��Ʉ�\~wL S�,���Ԡ`�E8(�":���������*������W�p.�M����?}��}�L笤�!�& �Yp	�u�Zon�?�/�m� \�{�O���+���z'8���@�����꡿a`�p3W��:鄆=j\H�]c���ͱ�6��$�&�|�U!���1g�RMj)��z_/�o����~4ȏ�'��3��R_g�����4���}��B�9�HD"�f�^�< *�>�U3��$�a���~�Zk�T_0���-	f�%DA���rB�pʺ͢�0v�vS�s�2*��t�ߑ�V��1�u�w � ]�����6�g���5kŪǄ����1�M�,�H����l���%:������(T�m���� �?���Wf�:Y�N(
�ˋ����4M�؟�y��}r�v�m�J��Ew�C�hH��LnG�Ƭ�c*I7��#�Q�{Y`��bd�6�b���z(����y.��ҋC"�{�G��r�pH�r��%�����Ц'N���%4��q2��Uw\�F��^��G��ɓ�^��4��٠�/�<��:_�JR�ݔR���c7]Ҳ�p�U�H�j�J0p�� ��]����Z&fa������L�F�O�<%�_\b��R��6cl�i����ZD3ô/��*���l5�_��;3��ar�H,j� Z	�"X���C��q۟���o���햞b�X+b��}��'T���Vx48������A�i�]�ǣ�o�����$�DcaO7��7�b��Q �G��2��{��n��Ia��XQ����Snu-0݇�j�I��<r�"��d|-����Z5�Ĵ�m��y��c<��7���B��:g-��煡Ћ�ҿ���*!�d0��ۮy��FT�-��c{_r��k�������<2�~!p�=ZI�k�qɚ�<��F0�����眈��V�|����Q���0�+���]������;����;Z�X&S\���i�~@�X���Ɯ��B�,�|��2�WtV4-r�j]�1E�Nb����r�����ÅՀݗ��G?M51��"x�C��^Y���)^˸"ϰ+a����k�V��@�߯��vn`���j��T�L���J���b$lH�j�ϗ�2�s����+0�=w�X��CZ�v4jR�����$�6�d%� Y��(nP_K�l.~��l�Ρ�/F�5Py�+�~��$��"�gT:�|�go�hnK¢2��lX�)v0O�u2�Ц��U�v�jsYWj���h��\ۂN�7�A,)��D�zT��0��]Qi[�m��4��j���f."�5THbG�T�#��r�Y�0I5^8_
O濽��Y,��h~���H�~&��@�O��N �E���Kyt�#���F�)�#9E�T������0��,�T,��b��1��J8�2�1���P�N�z."1� _@�F(�xѺV5ZO�L�����r$g���0���L�tG΍��/�z,�ϬvC���]�?t������u��"�l��t�q����&��m��%	��x"���.L���Zsc񴳿:v!�YF5�$�g$c�����JٝLz�u���z ����Z��gW�JM2��s��Z��^���z���x?EX��}cm� ��n�dkXȅ�;&Kۗ
�;f$=��J���C�X~}D��A�Ǣt\��Z-A8r}�z��{L����U�Ҍ ����Ahwϳjj�Ӷi�S��ȑGsFd�eޑ�\��	tcC�o��	>�7)|x���,�PV��ۉ�5$�!�4x�2]'aJ�l��k�G�c[q�U�c��hrn�@d��B�x�U�N�1�#�*�{����Vx���5	G�'���T�T1�D�.�s�a�}��0�m0
���"�<�d���W�3հۂB�6@,�Yg66�|����i�"x�X]�����1P�����h�w?,�{��S��a�9���U�V�^}���g�ɜ<���/^�wAaZ)2f�"��Uڴ���ɥs��A��Pt.�Η��f6c(�g?�Ih���%Ɵ0�2��\P�޼��@��-_ꐼ?��̄�X�X-�����㴈52���V��Z�O�m�}����((%%�c�N>}�g �S�s��3ϑ���+M�I|4 �?�����G�f���J7�lN���u.���v��&�0��
��ȉ;��g���U�j���� �k�~7��S��yDK����'�v�"��l1t*�����p�Z��l}8�j����dĀ0w��I2���r�<��ci�x|�czŊ[-\�����؞�V#��"�W�:o�#x_P�qSN����3�I�f@ങ4�%��:�DB�'B$T�ZQ2��6(J��7dk@Y��xEx�P���R}�+|�w��ga�.�9?Ɓ�`�t����cW���&�d�d��ۼjp�>|)Rq�al�v�����2�Rut�T�gj��CԬ��#P�P/ ^(�_X*=���ssy"و8��om���U`�.��ic/������ <�Ɣ����jI�Z�e����=D���U
�DL�NV?�.�p/�j:&�(!�� ���5����Q@��`����\SvWQ�8 (���0�q��ȶg};�l�*�I�!qsB=�����m�sǫ�_$���tg��y�BY�� �������G>�WK�)f�\8�ݶҘN�VRR��{���x�����j�D�#2�_O��?D�\ﮤ��q��8��r�]	H�>˿!��bf�^��\{����Ke*��9��tԎֻ�&M���E
[(�8����Ā��>�͞���e��+�|���z{�}���v�;��ǝJ��s�����&�b��X��=3��ɶ�˘�f�]���s����3��}�p�1^ITJ���*vA��mA��OfT�QR.IjI��!L�>%�{/�����8��`�Ƿbtq*�M�����>�(�bOe�w�R�zg���6��pt������N�\����ӝ��I,��m*�K�B����-w�e�S�E�$�`R]�8Ca�:d5���F�Mh��zm�����p��A���O?�.8�#LB��0]=&��bY˗�uS�7�GC�H��\;O���+�Z7zk�8tԈ���\��Ő�a��,p�h��5.���N"Hc�廳�tH����`$���|�ҵ�z��1���M%$ܕ��������4p�'Qy���bR�����>�rI�[^��2�9�/H�t
�a��^?�t 啂�p[����d�o��a�T��p��X	���%��ﴪ�в��jʕ	2��|Y�n!�*Xi���q�c�u�hIO�m �6���w6�M��n�mk5�����&�����Kd<,kG�������v��vM��[�R���H��7��D�R�pv��	��J��sS�M�ʇ�Gx�Gfv�ո��� �DC��g�n"l��	���vI������ʉ�d��1b��z�ͼ,���k��>��֔��K۸pc�r�\%���"0)�A=4N�E�c2��e��!ow�JF���Ϡ��dh^�L���B����<nr:��IR�ѿ�J�3���c2�g�EKDp�_WH�}J�Ԭ��r�����r��&a��*Q�<"��rOO�� 6\�
����6^a�i���z�Nڛ�Ϡ*��lp�_e3;;.Ø��1�H�� u�"�%���Wq0L��;���\(��LnX旱˘��'�s��z�W4sq��~�(
��A3�]���슨��eMdo4D�<7N�2��b;�� A�
�	U�����I�DI�w�X�s���%nИ0�^ ��:��V������Qm�dq|�?�b@�5�o ��p��a6��>\�ԏ�?���=�:�����r�Ц ;�:��|
!*dC05�t�F�̓R�{z�=��3񦈹��6�<��
�y9��q�����z�I�]�!}S��<�7x��Q�Q�*�K�K��z{]�������N"��������?�Sw*Я~��~5E�$�uab`�=Z��ת���(StqO�r9�Њj(�WW��8Ko�m�O��/�~�����;��)5�)�]���� R^T���LW�݈�+|�����V�����]�Rn	:����+�LΕ�J1��b���Ƣ�A��s�O�JK��F>X�AZ!�EL$����?)6����{�g����� _�v�.YX�l���K�F�p�ym�9f$36~"1��:��|��oRK��~�-�8Xz��0jC�2j\+��k��hᐨ��T(�z��h��۝�7v�0~D�͜������Q�vmkr������8���cTY�ZGkH�#�xFrܟ�0G�/�
�R��YgvhLF��z�~�0@k�⳺�.��޶�A,� tT�T��Cl)#��E�������H3���A,�b����,X�J�f�������H�1�ܕU+E1%��@����sdDV�LU���ݔ��'�qc�A}L%�Έ��	E�]ݬ�#n�`A���~-V���$��p��"R�m�/���ʩ���\m���	��@�>�}�.�x��F99ck5���َ4���_�$$��|�I���P�0me����J��5�hܢ&������R�$���R�����yE3��=i��un�\��L��@�;A�-�f�橤�rp���~xdV�o��͂��\�f�Z��_rX�� l��5�@���JY�{Sh��j�Zn�������,�WF_����`�B*�~{o]�>���|����X�V|4��Ռ�ܶ48��2ح�J��猦�Y_�f[lK1���?h-��@�0B!��0�o�l�d�Ō��{�M0xL����.�G=*y�z�T�{|��RF.�U�au�}>!��Q,
8@"���d4�-W���3�]ႝ �@�߿t6���6ͻ��iR�xf=U�Ε��R��P^��t�%��F,'�G���z��H9A2U��q�y"��O��� �<��/�L�<Z��j��T�pj"�Hd�N��A@�@PTBΒ�f�!(xk��d��s��z�%mYk\��޷���P-yG�&�����3�h�lR�����2s���rp�u����2}��Y69�(�h|�^,�>�3 ��s�����mڛܺӠ4������#�9�u��*��qb��X:�~Ͽ�k3߲�u�+�'
j��D�ߠ���ԵU�oE�3�� y ~2.�'Nl�þoK&�<���vhҥ���̆]�����^�u(l� j?�)�� �Ļ��ǯ��͟�h�~���x��Lz@�^-7��9\��9�VY�}Z���U#�|��Nk^��n׏���f;�♏�����D]IQB� Z,�q�����"k;�x�o[{x upP�n�R��`�T�GYΰ�~.�����F�/V��%�W$��&v�dԐ$��>wQ�qF�ʍ1�*�R�,2���t/M-g��Cϟ"�~�[P�Y(ٴ�*��7ݤ{y]��Ӈ��-��CC�`qW�ӄNw/<BX���E<B���.����!I+eˆ���h��v4O
�pL�g�?�ook�Tj���(�ג -(�y��g�kQ{"�`�z���{�v�Oe8��	2|\��֣j�j�l_�3�!̜=mY�ۏc��6_�ln�$�����.B��� ֺa�:o��O��2U�)��8����N)���l��g�߃}���6��5�bD�{��Z������:���|�nT���;���d�� �˺7��7c���S�w
�'.�e�`ϟwv�P�ќ�&����fQ[+�緳�φ�Ļى��p��q�����|�tz�$~�j}�vv��8N��n8�	OK���>���T��d=�>��>K�f�fݟ"�.����FI3�(G��d#^$u�I��!��vN�PRł��T��R�@�j����\���iy{*ȝ�@�;��I@`	�b��yõ��B���_�M>�ֽQ��25em��g+��6_Clt�Z~�r�N���7$N�D�	,��(*?�B�|ȄJ�Qw��]S�~�eG`��8^<�:�s1��4��1˘`k�m�T>Xp����R�?s����BL}o&�˸.&�}Y&FDu.���.���#*�\@hO3k@+��DzƔ�8/�d�X:��Š��aֶ�pi���0�;��R�H]l��	��fe��G�$#�i|,o��u �1�M�>�ܰ#��eE���K�4>p'�=���R�aY*+�����^���B?9,�Hz���\��^�', ��*���X�8d�?D���wbT�������	2�%����Ÿf�}��py�DS���Ĺ�i}�*l3��LN��7R���u�yB�Ј �ꇞ��6IT&�)�jkP���zĞ��\\Ԇ�q,f߮��E�",����q��O����D�#K�Q[a�u�a�M��������S�*	���M����r��;�v�]{ q!л<�C�ş�xn�(r�D�@֙�RN�1��Յ��d��b�M�z�X,�g 1�F6*�9"h�1rQ�d	p~>pr��%���]����rNNz����Uy,�wRn�FhA0�
����?^� ��H ��wL <4�:UuR�:R��:��Oc-;9���EpP��HPJ&Y��ֆ�ӄs�(�&\�w��ڬ�����ξ�Oʻ �=�\ؤ.���=6YvjigJ��q�Ni%��*l�l�AY_ �V;)���H��" �-�"N�X���>qQ��F����TW:X���˳��'J$��U��4�,�HK�A��C]si�쥠���`�?�'D�͜7�-�tb�@� ����$8�}��$wI�HNX�l���n+$�0SU������?���B��Id��[�P��'5}���)���p�Ȭw��a��8��:У�]�����ҵ��W(�!eV0�+ƮoQF
����{�pX�a�]�c{��q�p<S[��tq����걜7EԚė�����L���҇�L�b�W������fk
����]������!Ɉ�ۘ+����wtS�zد���~����_�j�G��8��2c����t��r��P��כ̒���ӛu�h9 �Bo�9$��ނ=�05�B$ј���y� ^O���Z���b�+��i����V�P��U��2�n4�y�?�ʏ.L��J�z!b�)���j��5�s����f��6�X�f�Z��- f��>Mĸ��26�d��W�j���Ԝ_A�..4�lSo�e��F��jy�O���k�$N��"�:�w�|6yo��qK�Φ���eX5+�0��2���r���*�C�kOn�՜khD�X۸TJ7�����DY]ۜ&b��R'Q��m&���F���.�YBT�@G\�#��Fr70�xJ�
Eߖ���GY�9h��?����~��V@&����֒���ޑrdgp|t��D��`Y)~|ZE`/��/$���U���g?,��'=�'@�J�M�Q������	��0H�1`q�@-���n�V�^�l�����hu��L+(�|@�L���΃���Fo�FO��#��DK��9�h$/�O���k'�"����~n��x�	m�	&�:��s�
�{.(�8�c'A߿0����t̚e�$�r|�wq��S�����ӄ1�7��.��h����π���M��s=��gh�Ȳ����E����7Y�6?en�і!a���0�;\Y�� �fڰȤ�wh�yɱ~s�d��;��=،\��Z#�3r3��[|Χ�s�K��B�:�6	h���jk�����u��,FZq#�G�ˠ�j���&o�i�>���|���bFFVw���I�u���4S��2STJ^8��������[g�(��$h��C@���B��1�A���Y�`P}��vcx~��G7G�f�F�T$Û�S�N.�W�a�Px}��y�U�
��$"�
�doRWCh3�*c����@����%>,�|͖��i�GxB���-��@7P��*N��6O�j,b,�L'��9_�Uc������ʅN�˘Y<^/�'�7=�Z���d4W��x����)mA{aP���΍zuf�%_(3���~D��q��U���}\M�t޲f��Eb-�'��A+̺?��{}����L㪆�2�d��-�$ȐI��c'�}��q��([�+�Y�3>3�� U�-s�p�χ���H����}�4V�#��锰�O泔���b�V�YIa�H �M2]�&��
Ō3���.��JC�J&Ug���nDN ��~-� �hX�~$�KA������vC�}�K��g�h����;� ��el�(ej�꓂��K���8��d%������Ѡ�@�x��=z�n-�t=�����V	;�������\#������NF/~�������f6�L��]��Z>Dx�B�Z
˜����'�9k6�k��L�x���P�"Rs(�?��[�����.���7�,���C�"ĘW�k�&Q�d������>r�`q��H��ZE���2j,�tje�g�wCʲQ��mP�[�(�)�*3^���y�6��n��ٞ��4`,�Jӟ�s/����ce�<}������K�I`�Se�Z���4���T
՚+L0�?!�f�2j��v(�6� !c��rE�B��Q�f�`GF-�̺_vn�8v�8�$S)��J�~>��|l�QN�=�!'�=(΂�����i�~�G�$�AI��F�	Bm� ����Uf����Í)܃�8(�ȸ�N�+M�Gl��I����
��D�p+OD3�n�U����|��
��]O���ĺ»�����:��˵m-6-�ؒO���y���,e�&�
&{�Ď̝�&���!}�[F*��.����d�����tBI��<����'�x|ȑNzqv��E�3Ա!��q�i��dż��߈�*���1=�jw�?�[���f�����t���3�x�fL�^�Ꮬ�����	v{����b�=߶T��wRs�j�,���r��t��{%��ʛ͔��,�`$�bjLu���}Yg���7>�|��t]���	g�]�6:�t.E�K%N�XH��q(���-,���*�R�Bc�o����w��S�����Z`�D@8y7�:Z�c�&�����{��P���p_��48�?�a}�L�c�f4X&�l�Y��u���ɒ9�u��e\{�O�Q+���z!�i8��$��R[[�{Λa�p��+Q�Nw�H���鰭>�Z��!�$^�|�+��pP1xg�M�yI�˵]����Л4y��'��V��"Rpvc�[�:L�Q�vr�9g�aHz��Wh|^��C [7���Ǿ���NT0�^����	w�%ut����30�K�p�
�G-2�d�n*�.3�E�"��u��Y֛uy���X .�@��/�6�zb��z+kk�o��c�u8����z,������}}�VPz��c��H�_��ы䌽�xL�H��&O����)�i�3M���*��NP�v��[U�v�qC8ǀ�]ѐn���lV���f��p�@��d"V�bƧz��ڼ����� ��4`�ڌof���p���r�}s%�6���,��w�`N��>����X�w�|�FCq�E�ܚu/^�ԗ��sg�2M<Oz�:�o�R|Ô��ަ���Wc(�F��'p�uH�jJ��5���ʙ4���$&W?F���H������*�OE����\_��#�'6T��i���,��h�$�*G8l��_��	;$�>�r�H]ʃ �o7"����2Vq�����n���і��FX\c����q'����0�4����^? �A�	].j������w|!e�D�q7�?}(Sb��� ����?;y��N��69I:WX"�#��n��0l棻���L�γ#b�E0dMXs�X�.58�����WA��S�J~�uP��3��:x�\����܈��0P[�2_�!�h�0k�o�j��Fe`�]�{����8V�>]䬰�<��oɅ�N J-��R�՚?u��v�����m�A�G�o�MЂƒ���%�p�]]mC��5���cǆֆ=L�(��йS��ȯtc�~��n�����M��3�Mɍ;��c��t��r/F܊�e�����n��c��r���qA�.
����d5�{��� ���^Jfh�:���S\+��:�	�Vl4v��m��Gy�n�M��ֽ��L�wJ'�b���{%�w�s����<3��nFRX�m�Z����l�y���u�6��1�%�����_��./l��� ;�F�F�y#*�����$i�#"'�':�S|q�-o��K�����X���0��h2`���MH�'u��"�J*�0�ih����7l%N���D��|��*W�.�QzQm��i����.+q���T��gG��:#禃r���0z�esl
��t���Y��3hOi���>H~7s�@�R��Jx$�x�lYw�2�t������)�X�E�M�J���>���L,5�e��"H�JIU����1E1�'�ӕ�1�I�@ȅѾi�VF�C�e/�(���M�'���#�L[���~+?@��]O%��C��Vh��������o��f��"������O����mvI�	a��I���l.]�?�V�cB7���Bώꠜ��i�$4�A�rp�ٮ�>����L���v3A�����%[�є��&��θG���~��2E��G�.R=�Ѡ�n�f�|�qȶ�;w��{B�f������t��B~n�%����"O\يZ���r`���ݧTHh�vhҝ?\���mh�dj��`dI�c�bϨFUgLޢ�����K1oS�Q>��s|)Up��S�Vrى�vޥRn�4nA2��J9��A:�mW[bC<�t��h�rj@� �B����N�N��3R	_"�љ�x�5����G3�c2T_*���Ϯ.~ya+�&}��z\
gu"l�\d�zjW�؎3�a�Si@]��4�uN�q3�i��/x�f���C���PԤ��EHt��E Q,����硋��y9��U�s����Et��00<@�//"�2��Z:������>��\_A��APE�fΈ��fG^(��B��9r�
���0���$\�a�ޭJvQ�-����\Ѥ�������<�����52)�o���ȫ�2���}�`����(��3�T 0>�dj �0s����N�#�	�0H�4�ɶ�Qx��W
VA� Q�����4������ܻ!�i
 ��Ⱥˡ������BUB�s�$� �~(�ݢ��9��K\���iSv������L��7G��@݋vbl�P�j5ꂇ6g�1�ǷQ"������������x��6z6��-�]�ɯ>��o�Vwm�3�V�k��#��K
V�N! ��Ͽ�&�f1��ED��YD��|B��Z⥣�����Өk1o��%^�xv�"P���R���ԡ�}\�8>�.谂ƒ'�����=��W�&,ڭdJ��;��>m�q�7獧Z�`�U�o�2Eɞt���g;[�C��<�4��P`9(��*�LP�Z�.y�y�	�W�	ٞ��4`�BӺ.X/2)U�>X�<�T�d���I���eAN��4��l�f
�8wLk��?�P�a�-jK �(R�� <��v��$�Q�ʑ`�1���@vh�}81嬫?�R?��Y2�.)l�����f�!�O5=�b��ȇ��u
�"��$9�~EL+���Bj� L�y�p}��E�X���H)	Y8�4_��x�N������Kc�y�î| &쫻oDΊ��P�L�P���0��J�dU���[��{g���+˰ß�B}�M@����Ѳ�e�qME���]1�Ǿ�&^����Ȑ[a�~���S��Z��1[E+��(�'G��>O"|�?Qz��� ?����[�n���d���[�WC������=����z�@�D;fӃ-��W�> �3���SK^�ؚ����W�v���s��V�T�>uR|Ŧj�ι��Om�S�{ �m����i/T`?vb��y/���Al����>�_��s�9��0��Ng!F�6TtU!`̨��N|���b��ߵ,��V*��B>������w�V}S�P�5v�`��F8�R^:�P��ct���#瘖���O�
��p���O>�?i+�X��L�wp�й&�{mY��u��)ں>����Q�\�8�OiX2+��tz|��8�B���+ͺ#�VpaL�jp�]��&�↩�tH�܅�x����U$�;�|b�k��1�֫MV���g��[��{u�4��8'"�'�R������U�%�̿\�Q��9�/�H�,�Rn^P�� �����m�/����F�T�����k�	��b%0p���~��
��&��������_�*"J� :����<���PuT�D �� ɱ1����6��^����k�)��p}s�P4���iX,<��{���1��f��)��F��x���?�׫A��C����F�:��7H����KM_`��e�����v����ߨ�1�>CS���Un�ެ�(��b�X;��b{����d=K�b�^3z��ټ�F��|+�/���ۘ|��p���r�`�%r�����*�>kN�\�t�,�� 7(#�wH�gFB��l�5V7^�ț������<j0�:K�ORWl�����U�c#���Vƈp�<+H9/�J����Z�I��Cu�&R�p�;MĀm�����O����[\N9H����6O ;ip��i�߁G*"�ql!�"_6yU;����/YH� ��]"D��կ��qǠE�|�����@�
̒X�e��$�'@�5���4$T�O���`ADH]�O���%��m�_DO��7�#ԿbLa� r6�Z^��s�;�ڌ�IMK�X��b�!Dn�0ɢϣ����°Ύ$�b�d����$�s��5�T�� �4��+^���]���_a�.d�:������=��l7ҫ����J!ۚ�0���e�:F�Q��5
{��%�W�ڦ_���R<��jA��wB���m���r���#���E��!�B9b|?�=�����	����]H�I�p'tWކє+����DIcS�z�����~�ݫ��>�2s�.����3A��^t�`r�$t��3�3�	�ʛ^a������ �Ip��3%�5��>��௳^E�f���{�vp+�@T��}�VG8(������n����/�L�@��L�qJ��8b�g��V՗�Js���ם�)v�X��kZ��W��(��W?�W6��Ό�:��S���_7�.��lɏSě��F��uy~$�j��$��""�):��|�T6o#��K�z��>��X��d0��42۾A�(�N�b+�y�DE[b���h�ze����7�[��DϿ��\E�*aQՈ[m�����!������T
�|G<��#�m�r�2o05<��
;X���h>Y�h�';���)~�D�@�������x�G`z�Pt%
�����)4U|E���e�ҹ�ꘫj,p�9]!H�pCJ�|�Ǽ��L�!�Dѕ���1�A�@c�Ͼd�IV���6�0}��^F2�`��&�L�^��y���!�x_��3�ѫ-«� G��E �a "cN��`�{�!�.��mQ�	����P&� z.����w�cc]M��&�ũt���$ϩ?�m���	�U�aj��g����W�Ưv�ST�϶�e���)@?���j	��v�E�P��i��l"�n����7�qЮ;��]���f��6�6����k~i�U���ͳ�5\�L�Z��r����� �������齐��h���j
�?v޹?a����FP}Q�����sL���#o΀�>c�l|d��Ԙ�Vm`&��vǥz�4��A2IJ���W�0�[]�k����h^	5@ЎB�������`��7_�϶,�x}��څG�?8>>%T��V��>g.y��a�3�}o�R&��
�.2"GX�d�wWy�-3�$ۂ��$@'G�cf"���L�ib\x7������c��P�g2�`bT���� �,�\"��Q��-,9�U�[��ѡ���e���V<{��/�<7-�Z�'��ň������Х߾�A��P���΃�'f��[(�6L�����Ρ���U_\�R�ިN��,g-K�C�w���2����b6#=��l2����}��Ƌ��Y�d}z���v�(�\��O��>�=� ˦s���}�	���(�k2�4���̶\�J����Ҕ,��X83������߃K���t
{���u�8�����U>S��$� J��~#��8����O�KwW��}i�v�����[�~���p���e�F�l阯j�a,�b���l�ʷ����� �y=��O��x��7z�$�-�ê��_��
f+V��!��&��#���7�N�0��e��_f,�ԙ�JA���aD�BF�Z�aL�"ER�]�ok,ae����x1+RP��Ri��{�|������..�m�����`���Xb�W�б&��d�x�ւ�>h��qW���b�T{��x}�2 ��t��!gֺ5C�8䒏YPP7�(*t�*)��5S�yݹ�����'��T{�`������$/�̵�kT<�yk����0I�%e�a��O�E�矄
��RL�s+?W�n\?Dj�3�(Ta W/�������Q,O�`}=k�\v�
*8��Z�[����4F�i�al0�����!�؛=��,��_E��J�$tV��-����Bŵ ؋�����y��2�)R�*8^�e��X�N:��>�׃�m���M)�W8��k�DiB��K;����*H�w�XM����x��I6�p6˫9��w��!s�ț����e��k���G땎���&�Q��4[|�V�$(��p�l,E�%��4Aт�<��E�|�|zgy������'�J�	u�_]��l�}&�x�o=q">ٵ���7f�%��?9����3��\{�^������*�v5��a߄ų�T���R�7�j��߬MK����{��Q��$R`Z��b`�pT�Z��I��0�3>�b/��V�cޒ���g�N16�*@t�4��C �Nw�m�Hl��u�,�/�*�ٙBe���uwS<S����.`>��8��A:P���>�_�9MS�1���Nk�e�p�@z�jd�?�{3��L.�����S&�>Y7�u?[��2/��\�wkO�+���z��K8`�Q��H:X�1�4a�5�p:�H�!��� ;HO��_4f��}5$Ԑ,|���fP�1.f�MO�:���%��V:�4�0'�W�r�R&�&�ۉ�p���G n�,29ݚ�HK�\�M��^�w� �|��;���R��4���z�Tf$-��\K	-�%��Z�� &�k �v��}^k�ZQ�*}�}����Q��O92u/lN; d�Z��=6Z'�Z��k����	Ж+P��7
,ׁ��vh��3�0�̩7�3��>٢�?7���F+��>��ܧ���Na�R�Ś_�M:���<����v��k���T/Cn��S��n�\���iP�ۆ
̹Bu"ն@hdX`Ub��zoP(�
��V�*<D�Bʰ�7�Sp��rwd;%M�|��Э�mN�����*��tC&w���F�:���E���VW^�ܻ�Yz���<��:Ƃ�R25*�6���vcx����p�ƤHT�wJ����g�������K�&Ms���6 �(���c�O;�l:�\�3ôY�c6Ju]ix'ᅢ9��v���A*���l\�_�%9;U�(o�H��� �S,"�{0Պ�q�������k�e6XҮ��J'������4_x��C��l�A��]��4��H��m��ڢD��w7��Hu_b�!3 -!�u�{��{i��nI�|%XX�����n<��0��\��2��B���iE�=�|d��J�[��|5�6�;��Mh�ڪ����A��T�)f�:.4o��e��q�&?N��,�!�G0��*�`XF�,>->{����ҽ��H�"K�<$	f�e٠������sњ5���������-�v��=n��>q���"��Z��f]�]#����T��̆���v����pS�*b�j��~� Y��͸��)~��CL*���jt���r%#�x�V�C����M�Y%:�S�c�j�h�d����nQ5fMT�I��J�]^@d���E�ɯ�+豵�
cV"\����}f�n�ᑡ�)���}�L:F�J��30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���șs	R�KF�Ǌ�pxC?�ކ�m�$�������D�29쩑�G]��f����qm�O�2ڡ�?|�>jGG�ZB�x���;�_�K��@T�V(uz�;G�7�L.���S���,\b!��IeT�������懎'��3��~�K7$�!2"�fyŻ���r���������������C
�P߯&��"k��������;i�M�'Wl��s��(��-�XD�2�����b�3VCU%�'��f��k����D��z�0�1
b��{�Ug�tjx�Zg�<�(ݶ�I��6��$i���-z�w��'�?!~�*0��+��N�Yݔ*	�k�'�m�9ŝ�~o�F�G㊂����H8�o�l�k� �<Y��=U8 8#��EB.���e$*�$C,�6̊.��� �%�E�Ak����^lCz[�[�Fs�q���^�d[�b���N�H���z�S��E+��]��+uڙ�UO����j�����q��rX�iC��̆b"�hԇ��y��8f��Eʞ.�0N�o��zg��ѳasjT^��H·��n'�:A9�&F9Nq6���*�OM��a���!f3pk�ܭs;���<X��x�!ә�N 0����5H���� ��;Wȥ�A0W��^L����\V��H��mg[�ڰ��92�!���*�+������Z�����1�p�����l�´H��Sž4�������D���6�A�:v��c��^ ��i�����'я�wPm��V����I�fd�jM>����,羘�6�_g()�~MQ�Q�֦NV���>�cv��ʭd�,���p�~H�ϒ~4Pϭ̂�ލ�%B�>K3w� ܘ�����ϏLUԌ;�!�Ӥ`M��4H.j����R� ���+n=rMQx+6��p�_��k}��i{����8�myy� �6*��t��HS��g"������1��΃� ��yL�N֡��tR]�,w�K!e���4��Y�" �6�jR�����˕�]h�m"wU/�*�.VC7�<��.��f�O��j�ù���ƑD eb�7�<��4�vďȭ'��C����D�$8�5�`��_8���j���s��V��2�^Tb�U�6����F���A��y��Ka�� ������jNp�=�q]������`�ڜ���c��Ί��f�0~�R�j}3�3�u���1N:~��f��%l� �M�RY|���d�d��Lg��w �ߴ7���Y�I#��ٲ�0~��yX�:QŇ���Q�!>p�	�w�ݙcg`2�y���XK̔�K������a�4b��M�e ��߻܌?�Ul���dA�%w��ٸ�k���	����+����aW���	;��sn�Z8�L,o��M)���hM?ޱ5O|rΒ�c�u7�v�L~U7��>]�I��&���z��6J��.Wز�:�n�l>Y�,#���PdJ�oTk>���9��)�3�����i>�'^�eVI������h��I��*���y�4�ӵ�e��*��7:�:6�[ ?	���=*�V�WF�@m��sy�L#��mo�+?vT�DA@x��nF���ӽ���#LM����5 ޓͽub�h׈`!�z�[^����'�(j����3�'��C,�L-���3޸��j�n�; �Y�����?�x�~~E�{p�ͫ�)�a #��%��=��C��ތ�Z�N;抍��^j�����qOG����y_(�WZPCd�^
�l�|LF�Q�Brd�{��~�����Xd�8�Í��eB�~��T�Y�7�F\L%$�M�=�oHW*�o���b�Suv�g�[���\+���lT�_� �|�?���h\�	�Ԫ[f�0�4�E�,��l(V5qA@vz�Ph�ҕ�2�H��8 YE)��+x���/5t�V��M#4S��/�%��@>��k}�'��'�6s��қ�=�r0Ij>ɫa\�N���]���/�̦+�Rݘ��z�BCFv���נh����.u˖�v`6:�Cx�v�V�1L;v�I�[��ш��ҧ�/�УT q F�'}�H#��E�P�l��+��\��� O�N+b��a�U	*�
�UV��Lb���o0�4n�hDwm����m�*��]�ߠ
<-�$�:7�����w�U|�d���'�/��QK�{�� ��=)'��h���в��*3?i��Q�����#FQ�pN+�B?,��/��cZå9��L^ U8[2�٤�9+Y����έ}�-<�;\L߹F�%�8�R�]��ʢ�)b�
���6s�����׷���IP�n�/`-=*��Y��G�@���%C]-T�@��AD��{C���m1�5�p����z�(�
��k�~9�]ϡ�F������������C����
���yfF���Fz[�+�'�X�FHw8�Ơ�%|A�2	�� [P}��M��׈ma�y�q����
*�׿c2,ᡑ�S�ed��NZm��2���?���>��}G����K��]<�_ %�����{T y�u��Gղ
L�jY��L�?�^!v���T�*R���zLR�=��1�J�!��MfL3��4�r9�T������0���s�VA����t߂�|��؅�l$n����#���N#GT�$:���i�L���� u.0<;�Ѥ�B#XkΨ_3�u���4%Po�{/>�8'0
�9USGk�X�!�/[��L�k�H��Q��`�ψ����l�]��X�γ�%Y�s2v�M�;ge��8P��_����@�v)�Zh#�ӱ�pr$�p��B��K��vI�U�@>>sxܟ��s����『���$��."��}w2��`�� k�-9�KI3.����Ou+�J��쪼p9dxN?����'���@p֘ҷ�d�K���嬈�ò�o��0��*�
��O%0�Ey�9�:�ή����#�������0�L��Du�+��T�!��}�ۗ<�&	�FO8�8Q��]{@�Bv )����s�&��t)ʢiP�W�#ָ#��,`�?͒�������BCYC���ॽ�z��䚲�1S,�p���H�zB���1��i~�te]o�F����A8���d����%�n
=g��ua�.u�F��+f2X���w�*4�"��AY�����j����N$�����m�����`1*�w�h2�/F�����ۗۧ��m�$:2Mw?Oi >�g�G����k���R�_�O(.����RT�߁u�4�GuA�L!͸������`!!�#�b�Tr1������{t�ݲy��4��+U!E &f����i�r�x��B���_A�=ǘ����$���"�]��������.n�MZZ 
z�Ն�Do���$-����*^��W�b�y�C��)N`�gpb���v�����a�0z�[b����{�t}��&�����]��>��7Dj@�@"/�S��J�1#��ݴa��HN�--�@E}~�w�;�j��ξ,e[�����dc� �dKy�������(2��Gݐ�p��҇�c-���{���t�=|q~���p�1���/�au��\���>7=�J�����Y������u�$�^/�+�B`Q{=�$�1E��Yx��~��i��E��nt� kز(�$Q���x檶��͕
.�~��ߊ%&��M6k�Ã�Bb�����t́b~�)�cg�ϐ�����8�ly6��h�P�ȫ���J�¥�J����.�m��%je��{�20P���T�gj�Qw�XJv�GtkJ �6�2��җ�CDx�j��=��-ɭ�J�!�Ty��@�<��KY��僌h,1}@�vU��z�#��G�;Y#"���^+��X6t1)���2�/�w���j-a�Pʳ�9��y=���H�e��m��J��oG��{�/��y�Y�r{�}D$�c�EM5�V�t4i�9���L&�Ʋ�o�$(���/���4�����~����J��6����Z B�y�|���T~+kgc�-M������O�� y�Y<˵�PrBM��܁n���d���`!��x���j��X����2�_VP�*�kΫj��w�;�v���`g ^�[27�� ��D�O���Ό��f�iON��C�ˇ�ї���ntY5t��W�?�14��^�?���z��G�
�Y٨��Y�+Z��5:3��V4��>�BE�~�����j��1@�M:��i�3E� ���s߹DJ�k��Nr��@�-�e�E����1imǚ�@�{ ��)��M0X�c`$�EA&�<��h��^�bi��́�4��K0�(�tq�������ʏ9�2Oxx\����������������xenfNvZg�"[��A���Ǔ��b�����՜�i�N�U3�d�`%�����N6'I]��t �n��>u���uH�d�2��ͬ�:�Fl�O�j~��� L�uVG�:(�G���FZ��O��lЊ��R�g��J.۳�˶\�pf}��<O[T��~�.{ �h��)��2���\�)7��r�\?����))w�n_�����ez.ە9g'<��Չݛ�!���y1����}���D*�
�md[Uz�+���ȧ|���-�5IC#���Q� j�;K�(��U�r��"�ͮޢ���$_8�Lj	���9�e|���%*�����^���TU��\�	"!H���-y�R����%�i��Vjo�51o�z+C/��̎4�ažc��]�jk�k�)l2<r�9��Ʉ0(�O �xM'��mBk۠��K(�%i�|Cb�E�����K�x�5.�UO�
e`]ilA�4�=����E&7
-C*�bӈ2q�Y�wT�҄Z17"U��2���_�,�~�M;���xu$��q�Ā��)�
�ʺLA#,��ѥ~���y����f�_������� >Ԃ/˷�JO�;X|Ԙ����2k`�����ɷb�y��o��s�����^X�--%A����/��c���0��r�dҎ�rn�mѢQ�:8�"�ӭ~qrW؊�	�~7��b���S:pR��z��L*� ����RΨ���ʇ�U��-��X�ڄ�aXF:"Gn��D�$9�Ӳ&}u������P�O$�?a�d����3�5�3&b;�}<o�'�o�L�p\� ��-)Hn�w�;����XA=�̒�L������V�M*Hrv�m������ 9IѶ�� g��Slj����ٿ��0���"p$����Cn���\�S\���!#�D�������!A����˅�c��"����9�~Lp��@m�,�V��Q��J��l�	�h��KC��"���J���V��y;�ht���g�/����Q�P ���5(����ǫ�,�z}�D���A�����(�B�Q֡_`
����RA�}��fB��;O��tNP��W��.�"�

�J�o{�Ep��NMda?�p&+W�k�\�;!�O�誝`1CyJ���d#G	����O�Eմ�s������1���v�G6�gł�.��,�lR�������q�>����
{�и�J��%�]3�k`���7&C�:�̻=��-�*%�	枦r�PS;m�@�v;���a����I�@��nrҊv�#B@���#� Z�]tA ���k�iRt�#�'炦�A��V��0��st��F�ЛF*�{��5�ܹ�ǁ+6搏X�]ݐ�^��&�åk��=���T��	P�*r�J\S������ت���Q���e0� J@��r|=M�J�$�\#�h̺TX��Hk����Ĩ�u=P%�a�
�uZ@5�dUq_f^�e�=]�z&@}��'���1>��ga�k����!�s�i�t��P&��,�8	P-W�%M����!/�s����*Ÿ�M�7�McyO��G���R�$��qF$�O�9�-�|M�V;˓��37y�'��ب�T��'gO?&�4�I��Q4ڵdU�'��,o�y��ʸ%r�����]4l�D��������Î� ���'�F
�Ӯ��R����&�ܒE�os��X��r4� �8�sN#��y��]+p`�m-����2��(��!�7�y�b���zW�#٬]B�9#�Ƃ��z%j�0����O&��j�("�BC�K���Tߟ��/pМi����P��͌���᳗� �bIi��K*%�Ϝ��AZ��.���*l����Wh�)i�g���*;�G�;v�C�c�D�>��ڈ�<�4O�'
�P�s��H<C���
!��h�TU�^o^G[P���u���� A�&�&o��[�q���1�G,��d��x��?��Bi�����T�[���i��%l��	�I�K}I'��v^тS��� M˯�.��_��u��^��0���a
B��{��M�"��7�7�	��J^��C�@�p�ɏ��o�rEY�9�P�0i7���޼��0�O!�V�S�H���b��Jg��z:��^B �VTJ*�W��4V �E_f���[w�4�w+M$Z����Dl�y����_��>db]�
0���]9������Xl"�s/��0D�ݶ���͛N'ir*9�6�~�h#�V�$���������ҫ��t�_� ��x����=�7Y"e��3$�K��.i� XE_˔��]����z�܈[OѬ�Srr�����z���g���2H��z5Ta��7��?[�+��rԷ����$�L.���T�^�X��1��/GbD�5��Ay'�1fr�3E%J.	�9S�ϥ��
	���b꜓�δ���():v�S�*Q��3���em��w��[���͞��S}�{Df��Z����:�k�׫*E�*澚���ȴ�[�f�F@K�yAx��6��$��G�Aa"����8�U,~�ꀹ�~Ŀ�2����N�`�DRٲ��i�f�U� nL�Y�R�1�_���^��Fg�O��<���`AY�e,����OtE#	���5g�zl0湻Xr��D3A��q�E�/ŷ�g��Ԡ~2J�]�C�F�敧�[����~����
rʴ��>$��y�F/%o+(LX�Q�w�a�����A�U��o~pe�x�c�S�F]ImV,K����Ŭ��2�đ-L�����\X!m�w2B�k?��>���GUZ��E��_u�}iܫ�m�TUD�u�+GJ�L�ea��>Tؔ�Q!kce�-T[������]��R��� .���!�eyf�u��iX3r:��q��A��R����_��y{����OȞ�/���������Mo����o��0<9��uGK-�����S�b5�C�3t�~"&�\��K��&�ԯ6�F0�,b���ǽ}t�[0�����!���i��˴��5��@�	X��h/J��$�>��a�XN�4-1\,��w�wW���qγ��[�wL�=Qc�Od�98��j��b�(�ޒG҃dpV$�8ce�Q����1�t�C�=��Z~��pdH͕��na����qo3����=\��K�#�����m���9>d/vb�ܗ�6{���$d�QEˍ�M�����i��>�e���Ug����k$�ɭ�����+�'!~�=�?P��T�a6����B�s�˺��� ~��c�ې��O��u�yk�L��	Pp4��{���i�6�u���8�î��A��jݒ�����2EGkΌܥ���j��wj�Av��I� \��2��f��8D�|����C��l���[��Od]��:��f��\ �����U!�POT['��&�j�/襰!Hk�p��G�����ȓ�9O<g�]1�/v��4?��� 7��	K·ʎ�<����
l΃���c+�������u	�]N&��K*�Z-H��t:�rS���8�{��ƨ)9c��2@���A����Nh��$5m���y�l�����M�I�&0����f���:Jttp+�_���Ҟ�ُq�e�i�}��j(����J�]�Hr�\���k�פ&����B,�����(��c(��Hq��42�Ҥ(�N�N�/�q�h ����j/p��뢖 �np´���SG
!�ly�0���[�ls�Ag���~ɠ.����Fa�)穎��mQ�V����B%����R���dk�u�	� � 8VN��;z�h���R8��hbQ�ᷣ���(�[��� ��W�}�����f�,����3B����o
Z�%�}*�}T��B�x�O+�N��W���؍��
b�-o�����»9�d��(�W��B\ST��@��|�1�=\�vT�dnZ�	>��Z�l�}�U���1�v�XA�2�g&��6ר��:b����Y���m��S��{+����]���0��n�
&.4h1�=��ت5ȴ	Q��r�3S>��!E��aFʷ�8ٶ�+v���@� Sr����N2��89#���[�o�?w�έ�ĩ��>��Pf\�k�Z�Y��	�q�^l��=^W&a�h�ٙ�f9��^k`y���y\s���t��&��mu8jI�WK��=Ա!и�s�I�����ٞ{�xNeM�C�0��[�������UqG���p"P�n�\M_�!L�X*+2�d�'�%p��4}�HGO?g�0�`�nJ�4{��U���'h�R,pd�y���f�ye�{�4Uٶ�������"��P�W��~F��N�O"�R�@���|ܓxZ�(�s=�m�GR迡oh��L��)��>��`��-%¢�0�p��gb�������{az8��٭r-B��# ���'z���2<�ha8���)�yBd$ڧ�T@���
K�@ɴ�qhy��Ӟ��n? ��i���*�:���XA4Q.��=+no��Y3W��i�[���6�;�0���CϠD�������}���'�{�P\��]C N,�k����ATY#����^���PJQ�u�������A���G8���	*�h�p[|�����l��Ex�����)�E��[c
�
}�%-{"��W��L�@IH"��?7��\���W�Ȓ��!Rå�/"�ꡫ�i����j^jI�C�Ӗp=q7�Qm���=�YxRϫ��05���6�W�|qȅOǬ�"N��I;�.ٜJf%����8��#�*ퟅ�	�J���W �V���_������B w�� $�C��Ќ�l$Mɍ�N�_?��d.���V���Ȑ9,�����lnm�?xJ�|�_݂J����'5A*9�ޝ~]Ri�[���B=�v�vY�Ƴ���$�j��+�� �5*��Oy>�Θ�e��'$�2��d��.�2� �FE+8���c�L��z	�[[��퟾��﬿
�� ��#a�H��z���߳6���3�+cy����`�|ǘL=̴<����XS�����bp��5�ly�lf�1E�=R.U"p���|��|A�nism]��{f�s|��.A�j%|@��_v��}�o)�t{O)6 B�����/����Uꔩ���#顭�j���yr5]��	��{�#U����9'z�=&%�d/X̰��_�\ށG����=�e}T<SP�]��/b"�4�˫�mg���)�	7�i���<m�	��=�oN���� 1���	��N���73jZ�n&��g�������C{j/��Cc�0zA���F�,���h��5YgV��&���)����!���t0�RE���vJ`k%+L4۽�4m�E/�Q>X���՗V�gdJ�����\�o���8!�z�I�����Jt頲�($ۯq�e�2U���I�`�6��x��_~�2qc���ԝ�C�~8D-V��eVuQ����@`3X-�$�-2��	N�����
7��zvH�٫+NBb��#�+�J��z�ć�:��`K��'JB"�ŧm�yT~Ps�4S������f��������]�� UJ�i4�2*�~��B�A�o�.�s)�Z��̀W'��i+v%����;m�%�z�UC��D�HH���|���ӌ�'��P���F�C>��	����!�T�)����^�G�P��u�Z��~A�N˪E��B|h0�n*�+3��t��8�x�"��٢fl����[a�CȖ�%��q�(���J[�I뻈5 ��!Mi�>N�*�0�m�:�~�Ru��^������� 3��b�<�"76�V#���i^���C��#p��]�C����MY�`�o�&0h ���3��o�����f���I��8�ݡ��J9%�Ƞ���@���	J�v9W.r.V_�r_�>��l��ecw�w�$���Ãk�l7j���_�2da�����,���<9���He�l�����O�Oݵ�Ƭ�O'(]M9Fy$~��|�c˨^��|�ư�g��ERؽ%a�ޱ� �H���Rg�&4���_~|��ĵ�r;��� r�����~��ׇ����
:�#����Lz8��)+���d������d�٨&�*Яa��"�͇����9*GD&�R�؀s�¹Ota�ar�G�37Nڲ��;5@�<��]=��G� 7f�}H\W0�ǟC;����h=���L�:٤pVޜ�H¯lm��7�!9�HѢ��ЃR��_8�A�<��b��[�;��pt�����If�O��S���q�����0Q��Q�`A�A�����e���bd�K�Ο����Qm6��V?Aȷ��ɼ�Y3����!4УNܬ��PVӚ�;AR h������~��*Q<D���B8(��8���|h}N�@� qb�1��jkUB!�ȡ��^
��뢬�}��BLO0H(N�"�W�a�r��
��{o˵�������d��.��	W�~\83N��������1����dsP�	㻫��^������&1�_�v�@����K������V`E�1�������aa}۳�� ��Q���u�d]���U��39
&��YƼ=7�M�z��	6�\r2��Sc����Ɋ��cܷ�/�T6��&'@�hOr"�g�s�_�J�!#���`�]�\%���Ď!}�y�P��L�0~�Z&�+�
=�qg;+^��X=Cy�&��͇�!��Wʞ�Mrpke�D�xWsјt��&J��I�8/��W|�؀Br�!u�s2}k�����^�	��w�M��[��ր`�ťsoD�q,D~�����K�M$5X�6W/3ym '�B䨿�t���??�`1�o�#��z4��qUiȹ'�L,U?�yVP���/�>G�����4x�[���2�^�񊪎a��uXM��F�'�T��RU���:�k�x}󎭣�sbv[�i��_�fU�9�
ۃĆ`�W-��U�Ns��:���l �z}<ْ�5B)��#4�ǵљ�z1���x��h���F� B��i�ߞT�@��Ӝ�!��Z���ڔ�,*�Y�5�Ai&Q
�S�  �j�Vpa���cr���/��=A*l)�uNO�C��*�]�������z��מ�)����y:(��_�NgcA���g-mm� �,�n���"6f}(͞UMu��z�8�͂v�]c)��n���P�.�Þ�ƢK��6��P�	y�v���Iv���3��&�<e���i��3D԰{�!'u`q��E"j�]s���
���Tn�K�Mu��6ZQ���ٯ���� �{a'E���_�3�$�6�j�^�H�W�gF+��N��1aу��(�e@��F����]aV�o��|�u��*"�K��"$Ꙛ~˹JZ]�"���/[��.'��7H�{�1�ꁟ�O���g�ۛ���D��ze'��7-=<�?�a���X(F�	��ED^s�)<����ȵ��[�5k���.�e�V
ɗ�Wb3���ڇd�����Z��	��4ip�0d���6�'~ �3�;p�]�=�:���b�ņ�B����`��=���T��R-��3�ٸ����U��b̖şɃ> �YR�.��	�d]e�p����$�Lğ�Cy�m��}��0�kmy#�:u'�5��Q��>�,L=��g��cy*�|I\Kp����a�S�T��ŊX�h@b�sp7���`-|c�^�SU�r�����{�dT��-��n�85`+���"��F��Q����0Q�*�-�й�@���v:�&��������a��hGk�U�,�5P
9p˅t�7YQ����w�p,G�o5}|�"ik�ճ����n<�!Ϭ�Z�_��&_!ϳ�sy2����a��W�nh8JSy������U�|�D��i����q�@�SE�z�L�E�!���6x�*�����<F�$Z �l7�sg-u	�:;˷G�XwF-M�O�����bgΜ����k	\��}ō�O��PT[�`�!~@��)s_��I\1n�`�[��͟/���I"N�s)*�nr$����z�l��a��������<�cg���:��;)���b����~)8h��T�K=�r�C3�K/ǉ�u�v�UU��>��=���
	�c]%�>0�u�P�*�DH�>��#�"Pz��o*昳3}9	,�I_�~��ݛ{7�}ÜelY���~�iֆ�� Z*�:`��m���Ka�"�e��"*��v7�#6=rH?�,��@��:�$W�ٷ�3y�IxL���m���?��"D�x�[#V�3c���r��I�L��-�O8�ީhs�KRV�����^����^����4j�R�I�|�j�!��M��:gĸ�t�D�{ �Ρ]ձ�*�x�ZEw����P���E�� �|M%�p����i��Z�ۧ;<����hL�y�џ7Ԟa�ЧО�(��`Z�����l�<J��؏����,�%Y���ژ��\z84�;��ۋB����#2YD�nF+�%�f(zlo�X������8��S��(ҽ��[��i\�Fѽ�
Wp �^A?��h�	"�x[|��
�I�Al~C�5��vPg,hx�䍈4v���Y?���Ht�ܽ5�����^��_��)S򎎐�h���'=aV�=��s^kth��=N�/hˑa�S����1�s�<��,�b>*��gj��}���veD���-"��c�.K>��.�:
�Ìk�:&v�[K�/���^�9X�qV���=�mH��~h�ԦL#��c�2\�ЧY�����b�����.Q*e3M������b���o�=|n��yw�P��Խ�*��^�5>5<C+��h~�g�!�:�[w��|�*��e�a��Qa�snI��I�,)}�~���������?�~�Q�ͯ���#�b��ƒ�+�O,~�9�\P��������94��8�y���3+o+��W��}��<?�vb�"F�H�8G�]16ʸ")8Ny�x;ysm�5l���O��Mq��no�߄�s`Q쒈���Vפ�P�C3<�����`�ߑ�B�Й�1I�qp�'��8�zx�������#~Oc^]���F��������{��>�=:
����yĔd\F�+kX��%wiZ��}A1<���&i��D�R�Gmw`׮G�ˠV�pQ��Nh��w�--���;�9W��ewt�$_��� �P4�#��@ZG3V��Mܓ\��<*3.]T��/��4"S���ݲ��j�	N����N�<D���Ή��ƭF��W0�,6:	�r�N�,3��^ZP:�㖪��UZ��+C{����,�D�'�Y�[~n���F�g�Fhg�5���=������BC���+j���դ�g�J�}8+��P�9��<�M�(�ʎ������
�2nJ��_��W\����ƙ��ƨ� ʗ2�5��������([�q���2L}��KIc�6(".�;h�r�E_��qz-L��9�C����̡@K�+L����.[1�U��/R�X��� X�KY��Ѕ�o��2)\uZ�%\�Ff�)XI�w}w�`�¢@I��ʲ�����`%O$��6K�o�r��z;�����qΨ�������c����- 7��zB_3�Q�Ŗ�kM��!e��;q�g����+v}Sw�f���ǭ���~~���tD*��H��:�2:�f���K�H�x��o�����؏a�L���b(8-���=�ύ1���E=�	�3�!R�$���,Ό��s��i�R��_'�^yhg�A��)��ڰ���,�P�8=t�^����g�^l�����j��"A��LQ��t�����:��]�R����h/E�A�^�����ܒ��<I��΅�гB���-��� (�9%��C(�)m�z,v���v�a68��(X&M`N?��@��-M���c�}��9���{�[�N��ƍρ��P������<唭�R3�(�Ǣ���X��~�q�[Ѧ!2#G`�]���?�j��܁'���t�n,3cM m?6e7��r����2.�{����L��\N��W6��NA H�gqT5���1�����,���⁔4],!����9�������"�Q��9d_�"�$�l]�~,"ƶ�/�.G�7�O]�ܞ��.O-��2�{��gDGe��7x�<�w?�%���<'�5W�4FD�-8�H6�qŵ.g�@s��68�0�V5���;&&b�`�%,O��=��=
�3NJ��:Z�[o��ۙ T�~y�p_�=����6���QO�m���&��	�y��ds���UR80�3%����1���[��?����yu ��,R�����d(���ܬ6;O���>��SJ�-����0��y�C:���i7Q��>_ ���X�Kg�
�y��þ�;8K���ʊ6S_
�T,��Џ�������67���`���B`S��ح?��[�d���-��(n� N`��=�����*Q6��;���B-bz��#T�d���j���R������=nY�̍��k�3,�ψ5;��}:��Y\���M\p�;R���{E�9� �Z��y nG�����*3&���*�j2�F:�JY��ns_S�w��-3�����Q�i��N�1uW@lx>P��̷
���v�a�Oȵ�w�q�dZ¹ܣy"�E�vX�O��ZE`gL�&f?2wog�3�7
�"O�܇6/n4c<��/��|ei����o��t�F���?� �I�-6
J|��!���R����ђ�r7�7��2I�O��ܦpʨK�s�6#"��$IL�ֆL.�d:��W���,�0W�����#3M��P
uK�4 ���a��>�{�0%c�U�$����!�WL��|�k�ke��[>�O.ϣ΃�G�8�X6�����n W��T;"��䤨�$�׽�{�{��)S`�h?T�&I�r���杨�Ʒ�v��Uȉ�>�韸g/���G���:��	_p���mO��E>
� #U58PUoe��Nxf9�=��6%9h�ݶ��� �eGfZ�����̽��U*N=Љy�M��P�ӆ�Mez�2*�>}7k>�68��?z���%�U��W�d^�ģ�6�LT-Jm�4�?�C�D��v�4Ю�J��t�)L~���J<A��.�A����1�ke"^�og�X�j�o�G�%#B������;������h ��W� ai�&�
��#���ֆۻ�]�\kB�M���i_T���c3������ߏD4���g{� ʼ5iI|�*Yb;��$�A�0.���^7��ZIeW��i@|�Pa�;±��o�BC��pD�c���T��pC��ט'O�)Po�4�;��Cӂ��>:��s��TL���^8�P]��u
?�H�A�3���`�I�}��#����dv��E~a�Z`B@�pگ��Nq��Y� �t��	1�3 Z������G��Y�J��˅+l�j�(3�w4D�����c���8�c�[I@��J�&��3�/��j!���D/q'S��N��k@��e����1~��{���n��r���(��ު�
�A�2hap�������� ����KUkI�9�L[����b��A9�*x]j��G�6�"��}���f�4�e�:N�4b�)����@2���@�Ǜ�~�Zd\N�f3���`�Y��`t���Ik����c> �>�91�g>�u�1l������i~�D:�j����M�8����u��:M�[GP�F��UO�J��/�C�g���ρ*���\I��}W?�O`�+Tm*��s�c�MAM)E����F\�g4��y�ͱ��&�A�}})��Xn�-g�mz�f�>_�ᣀ����t���c��BM � ��/﵈2lU����A�M�P�s�J5��"��4HK��j�2/K���x���"ޯ�h�C����8n��jN����|Tm^J��ț���qq�Y!˼��'	g�H�#�����R�4����iF!Vop�5�Re��(N��Q��ֆ1�c��3��tk5?l�2.� ��0���O-�OxD�k���䮽j�Q|(��Es6h��awx�����i
j `i���yJh���yE�@�
R�d��8QJv�j����Ʉ�7{4�I���@,�CM�kÂ�$*8"q�c/�~������qVg,}�
q)����>�J�Msu��9,���>���|�J|֤�@��=�׆P�kE��N�W��\��G���1�Z�X?��%�c䰊9�A� Ej�7\�7@�rsm��G�3:}�l��dMr|A�f� ~�X��g��;<�:�:��_�L��{���m�Q���Я��eՌ0vzٝb����a��"l�"�	&�9?D[&��->�#�O	��aLyk�ZR'P
�@����+`i\n�Z@]D�a����v�=���>�F���"�xZ��]��Џ"�`��j����Z�B�gݿ#f��o8��(�X"`��g�q4��wӠ��|�U���qho��t�5���k /wBIJ�g
vI`|P�!c6+#)X��!�փ�7��I!fĎM�I[�@�$W�#�a�$:�֗*���e訄�,�0��c��s�#e��b&u\ڸ4Q�I��j_>�U0�S$U'���=R!����M�k�^����(���7�4��4���	x?X'�6�+=ל�n�;�"��5�r�^�׎���lt)d3�hOt��w$rP�w���w�v��-U�b>=|��=�6r����j�.!���|���v�>�
#��\P�c�o֬:��mf9��<�u��*����I�)9�e��z��tӘ�|m�Kl*��jt"��'Gӷ�4e�q�*;�7�5�6���?K-
��3X�f�WH'��6Q����L�%�mq?�?��`DØm�����ߜ7_ښ�5L���g��Ս����*�^b�C���^B���銪j��q�ut�`v��m��x!����d G���	�W�V�~x8�UE���r�������� �@%�dN����`mzZ�?�;�n��l�%���3�x����s�(tPZ�$�`��l��|Ȗ�����}�o�Q����A���+8���"�|BU���=Y��FW��%�����oJ'��F3��y�S����iL�[���\�XCr���� �-�?{��h�<	��[�g�ඹ׭��l*ɭ5�=v��h�~�4���!��Y�U���4���/5������ہ���`�H���n�-�s'���i¥s
����&=�Z [17��a��P�k� �����8��T�ɮH�čĕ�v�t�עc1�O�.����8��:���ø ĳ *vE��[��?�>Y��uU��e*~q�K�i��H��#�p\�RZ`���A�ބ��ӗ�P�
b��.��̈́*��������@�bJ�|o���n���w�5���HI*�ϝ��#P<o�ۼh鄓���Չw�	�|f��ɑ��1[�Q��6��up))�7����RQ��졀?k<�Q�@p�y�p#QN�rF�+;-,*��ވt�çb���� �q�8��٦��+���1�}�w�<�F]�J�F1�m8s�X]��c��#�)�t\��7�s��a#-ʄ���y�����߰��`�c1��P��Iī��s�C�Į��]C�߽��|�k1uΤp�q����z$":��ݩ�m��~{�b]Q�-F�<���0e�1�6�k��G��
��,��*����F<8�+Ȝ�X)\w��p�D�]A�X�<�N�+$�p�o��.�m�3���
��v���12n�0�����'��	�m^�L2/(�?qT�>���G"�9�M�y���_"@u�j�q��T��ou�qG��L?���E�A�!�aK���T� ��!�&漺�ſ����^L�C!�`�f��O��Zr;����{��fU2�_y��X���sv�����?`�M߉�&�M|Il���(&�&Hz��-F���g�y���-b0�Cj����J�I��ؚ�S���;�0\�4b�z��j7�tK�t���1��K{%��[ ��4��P@r ��T�J�P����(aFO<Nn^�-� ��:$wd볉�\Π�[��G��c~��d-����d�X3�(���G�3�p��4kc�H�辿���JtTq=~�b�p�2��"����aW���~�;�:E�=�c��58��U
��ڱ5�Fd/#J���K{�%8$�E��|z8`@i��	����A����v$s�|���	��3
��y�~��k�����6��Få��B�#]ˇ���cp�~���:�20B�v(��'�j�Xm���1���e�T������r���k���.����"��P��͙O{_Z%BW���jq&�^PC�=�&E���E5�vv	�L�0kD�7/�sp<ta'&���<	8N��W{{L�!�!4��s�O����Ž�W��9�M�� ��m�?�ե2܀�bq�y)�T�.���MC�x���78��'ws�>?A�,��?�� � ����T4_��U(0�'L��,Ԓly�Ÿ�^�]^_�߆S4����u���>�p핎��)�Vjl��F���3�eR΍�ٶ���܎E�s�Cg�+��xG�����ڨ�"��`�2�-	�j씞5�m�������B�6�z9�1�B�y�#sl��lz
h������ZY���Z���BHS��ST$j���
��1���Z�U2�
�A�AC ;M!i�!*
�L�h�Au`.�K5��T��нWC�i����/;�y��`��C���D�e��ߜ����yx�' \�P@��,��C�k�o�ÕıT��1��?^�?P.�`u��u��J�A�w�+�0��]L��ԃl��$��В��)&xK����6L�)ݕ[�V��U�%�p����4�	'y��n��_�&���b��2}Wx��W^�%(�LSZm��?��zD��Α�t��mE�����L?F!�+kB��U�'���ZW������^r��j�����F��>��ħ�Cmf� � wT��9@p󆾣xh�EӟW�n��i���z �%��n��Z�Dt;?�8�ؒU�c�-�=�a�,�i(���ZB����l	����4�խ�0���p�����J�E8�{�RD�B�+v�FgY �AF�#C%�h֩�ozA�����A�S	��ҙ��[�&\�7�����[ !��?��hNӚ	���[�P����^��lZd55��v,/�hԋT�dc��Q�pY���Z����a5�����B^���t�N5��;�]1'�ԙ#�s:k����=*n"����X	aN������ϱ��H��Ր��꣮xa��dIv�)L�Ҿ��F=.'v׻ha�:�b����0���UvusA['?h�nJ6��luЕ'�q2w&Ù� H��3څrԂ9��1��w�Ŝ���-b�8���,�*����J���bz/o"E�nֽ'wߞ���ױ*�D�?<�G��f��3��	�w��|�`����Xa��Q���J���-�)Y?S�P���@!�w?��Q"���5#8>���ٱ+24�,Z2޸y�����+�o��8M�.��w+���3��}�[<"G��Fa`;8���]�'�}�)��Ԝ�sI����Xʴ�cש ��J
T��y�`�#����y�ŤLC�D�24�s;��|��w�1���p��.���zT�������w�~��]��wF�1A���o�a�����$�w��
ϣq��C|�@Fl]�+�g`XY�3w��t�RA�;��l0����! �#*�mӔ��#�p�����	�V2�b��ʊz�W
��9��m�p�2_�3?��u>/��GRf��}���O�q_R���+z��5T��u?97GG�IL3>}��*��q^�!�Rh�	���6詛=��m����&0u7C	�:�8_��P�j:�3����ŧ��֨uz&�:�R�G��F��,Oâ�.�"��ge�vn����0\��%}�~�O��Tl5L�R	��0)�/�K��\�)�1��O�Ͱ�v����)�~�n�$�̵�z�C]������U�3<
����݊:���^�\N#��U�R|�z|����k�)�ً5�s����J�j�Y KU�3�Qݢ��F@��7��N�8mm�j-����4�|��8ɩ��'	Y����xb����	F,Hm�"�QxQRf߈�IC�i�	�V�`�5�F:�DY�=���q���c���,�k&�7lֵ:��d<R0@�_O���xqG��k�YN����I�|�8lE|Ɇ=[x:X���W
��i���XU�U��E%�
Ѷ�N��wu]�J��3Ҩ��7Ʀ���(�k7�,K�M�
��n$)�Bq�h�=,��.�y��|�,!���I3����ϝ=�=�,���+���>x"��ۗ�J�g`�_�C�<�����ykȫ��������h�H�� X>c�%e��o�9��fN��#���vo�r����F�X:\zL�"䭢�r��
�I%~�VD��X�:�X:����5LN���}<��v��+�(���g�/�[�|��~�|a|��"�֔h��9~��&��,������OȄ;a�צZ��3�ڲז�;	�<���/�q �g�]�H0>p�a�;�����ί���o�R�U�8E��
*ޱñ�J2���A}RU�f�%��l>�����C���(*����8��1�Vf�WK��/x6N��k���=Ga4=7��ZJ8�֛���_��p3����wW�r�UR+8б�M�w��2�|���AR �j_�D�^���g����C�4�k*�,7��˂9't����~gd�l�C���������AE@tХt���X�Z 倊��� �/�x�A�
,���l$#�T��"w�H��d8���}����u�n(q#�x��U5�h�m���,5y����6���(�bM�眺� �v�`�cS�����H��7]ǭ]����Ϡ�P�XȂ`���s�ӔLa3E_q�&ns���ϝG�Z�!��`�g�B� jz�C�����z�nK�M��6D	E����y��_{K�� "�{���x]6�	81Ha|+g���8�1-%_��Ao��O�ܒ��¹]�DȞ;ِf,�;�"-Q�8���0W��E]v�$"E]�/E,i.Q�7��k��l��kO����-�w�kD�q�eQ�7��<�Ԑ��q�����Ҕ��DH���S(_�,Y
�-S˞����ϕ�V����i�b]q	�D��ĈΞ{˃�&��I���Q��o�<�Q~�띿vp^G=�B���gM���������fH�>��Y���b�R��3�h�Ń�C��黗LP��E._�3 � �R稖��"ddǣ�����:��-ꜟ �e���g�50�]y��:=�X�Q��>~S�&)k"$g�̰y����&i�KZ���	�S~��T+���>���L�75�`����S�n�ج�Х�?�d~�-�>�n.l�`iɅ����'�Q5�L�_��T��-��)~m��i���v�%rk�����O-WH�,ck,���h5z���B��Y;-s��N�����i@gy�L͑�?����;n&stK|���
���|��$�q����~����F���;�x6���ÿ�bB�4�!��='~U5c#Tؐ����ð>�t��y�:Q�Z�P�x����J����1~�j�o��)djD���7�2ls��=t��o'j��w��v��x�i �ޒ2*���WD�E��u�:�n��]4����|��}iYZ���t��o 19�&�������_1JG?��YAy۞o�B+��h�
�3�&w4�Vd惪�Xh��~9^.�@\ ��ƈ3�$�E���X\WDϻ��[�N77z@:��e��wҍ�07끠�_��o�����=�޴9�yS�q*���N>�1�j��{
TAV����_��Ov��+�����y�xM���"�m`T3V�tC�'KHL%�f]$"$�uOL=m�=�?1nWD\�=�@�и�=�ڳ;LH)��T�"�N�>�������;���N7^[��"�j�L������jn��7g���F�l��	�! �)0�b�=���xѐE\��K�?�� �� f�%�@�a����~Zs�%;�:��
��>�x�l�S�f7@�uJ(��Z�.ٿ9e�l�2��`f�=���g%�����"p��Ӛ�8��΁'~BngK�O��YI�UF�B�%?q�_�to#������U
S<��[X�\F�+9��� �S�?��GhW~	'�j[!���O�?���l].5�#�v��h�/���������Y`�
¦�5�a��5��V��� \����8Q�[����*�'����b��s#�+͎~=S�X��Y2a�<�)�3�ꅪ��K�d���Z/�����]�qvJx�{��.�J�q�d:�w�1�K�Lw�v���[�4Ԉ7� ��p�О�9q[w�⻅H>�5cc��+���O����M�?.��}�bDY��6V�*JCr	ם̮�bc�Qo+�Tn��aw(�i�Z�*r���<h)�՞̟�?��wM5�|�;2�J�?
 �Q�'�3uՄ���)�E�#���tBޥ8g?D�VQ�iW��=#A������+{8,äQ�A��À�������m8VH�����+'o��fL}�`�<�F�E FJS8�3g]6F�]��)}3�]��s�Q�Z�ʝONײi��st!�))&`H��m���"V��@�C�0�;v�����6e��i�1.�7pẒ��}�z=�k��	��A~��)]���Fq�h�|T��*[ �����M
�X��4�����F�mC+���X"�w�<3�}�pA
�����k���)�/���m��ͮ������2�2�.��3�������-mW9�2H�?��>X�NG�k��;���/_���í⫊:�T�KuhR�G�@L�E;��j��#!��vⷠPT�.��ze��5;!�Xv���gc%��!�uf玂�/��r��b�]e���mc����1����q��~�hn���C��1耩��M5�E��!�?�;M�-�Q�����Y��bԭ|CC���䞚b�s�M����ԯ|_C0���b����C5�tR�[�j��ݤ�0�Y�s��q�E��@K����J�1��ݘa�ڬN�T-7�NX��w={��Zwι�Z[O�ڠ��c�-�d�I��#�1��(�8�G�&�p(����cH5�W�ϵ���t-�=\~�^�p*��{TJ
�a�'��7L��0�=��T�:���qp]Τ�s����/������K{�3>$*��EQ|>�}9��aixRY��u��Y�����$��:�3���/��u�~sL���7p񚧢6������B��� �z����~��c�޹�Jٻ�׬ؓ�y����9KPv�����܅�'�|z���&R؉|���j
j#���Q2�GT�@��'�j炦w0=v��S�۝ b�a2�m$�D����c2�YU�m.�<s��7��Xc�/DY�U��i���L18������C$q���kG���Y��랮/d+�K��	�/3zC�4�*�"{�˂<�7�,�.A@{(=�Ŕ�3��h��u��[�DN�/R��Nv|@YL(e�4*�l�61m-��N�{�n��j�QR������I������h�xӚ�n��a'����K4����O�s:�Uj��:9/{Bx|��F�ԂQn�J�c��Nن�J�errhN��L�&#���a�>��M?�f�%�cл��9>N�03�EF`�&����Ҩ�I
 ��l�� �ެ��%u����h������ͰQ�:&���SGXs�$��u���:,I�G�*F^�Ob�*Ў����g�<]��ʳ�I�\�}��}O�gT̻?��[��l�)D���?\B�������~� Ҷe(����)�HӑHq��kx�Ȯ;�1�Gƃ3���4	�������)]��7��N@��u���!"U��_2sꊤ��ʒ�]=cj"�'�/�KZ.��7��"�3��r
�Oӵu����>�D-(�e��&7�X#<�ц�-'�⢂w%��;1ZD����&>�s$ɵT�c�&��������V[���!N�b��������O���y��U��e7`ρ����.R��j���8�p���=�)���/�ŷQ���^�g�MA��)1�%<�R�)3�'o�J����j������&�zD� �0nR�_���Od�����{���Y��8��
�y��䰫Q�H]� ��7�7��rs.�G� :} �=��r|�gf"~��ڇgS;#:�;��_�L�!���+�����q��&��0W	ٝc����a�I("l�9�	��9?��&��q-��$�O	 aL�K��`�3����;��<��� �U� l~WR �H�P7���);�:����M�P�L�&q"lV���H7N<m#r����R9�N$��R����A$�ݤ�M��pDQ���Op�nW��p(�����fS�������ޒ��*���WA��op�ɚ�H�֔e���C��۰��~�m�)XV4�3�����X.kR�K�e%����ǤZݿV���;�U�h�6p����Xb`QQ
u���A(,�s�'����}����ղְ����v�B�l֡�
Ԃ+�7:�}N�VB!_.O�i�N�rCW����?�
ܯ�o`��:w�sh�d&�7�՞3W���\�a)�����1����n�d��	����T{��Y���+��1�Lv��[ц�!�����r�K����ih���;�6�*PiX�5�mnW�ʋ=]x+��n��hr�&hK� �=L��/~�	��r'PMS����h!���F�l�i$���v@60Zr����9��9#�9��՚��qR�����m��P�P <��e��Z�'��4q|��^fI:=�J�&����"����x�"�k�����s���t7fl&?�$���I8�d\���!J7��jx�.}TYXǽ�a�] ʽ:�Y�1=�Q����o���b�ߨ�97�ʅ��/B����1�{�B�$���E�T��^����i��Ҩ1��M���^�$2�9�y�g�'(�Kݢ~�����r�A�6��S�dQ�BcR������~5�yc�5��P����7�y7w�?ՌP<�"H��� ���`Z�ͮ�����+j)cmɼ��2�ZY�	����Yj���w��`v�����@ (�h2Af��j��Df�֟���p��j�B8,����ѡv�B
Y�-$d�9��t;�򒒻5�L�}�
;	�A�8V���;}�h����ϰ��Qx7㣛�u(�!�Ӗ��EF}
#�<ᑰ��զ�!B�U#���
��V��Y8}�oB�IO�/N��W��خ@�
��No� Q��ڄ�dmF\��p�W��\tY��[�q�6N1O;��Md/�	�(�[��@�;��XQG�1���vWB�(K�H&�`��ϒ�F�me�}9�=	��\g��j��h�]?��!z��y�&�,�%�=s<�6��	r��r��S�i���8���^���	��a�@��r��Vׯ�)��-#= a�N[�nͿϸ���/vOP���Zbm9�Ɛ�q��^mD=:&��P��*l��މ��k!2�J�s��mt/&Q=���8�ΟW������!�ڕs�|��
����x�ME�;��_���R��Q� �qhBAڱ�?���>M�YC���vK�(0'�e��t�ډ��?�Y�+�U���4<;�U���'ik�,�5�y��Ǥ��c?�@44κ�ٗq���ʋ�-�z�ɰ�I�	�FF,5��R�����vܴk@�iYys�㜠�}��Be�ՙ܉u1x�?ש`>�-f�F�땵
�)�Cbb��!�\�z9,��·�B�v#pT����zG�쇒�M�Ix���OJNKB���P��T���Qݜ�˭�!��r����
���� 8�/iw��*G@�E�nA�B.�XL6��& W
D-in<�>'!;p5�ݷC���D�p��<���Ck�'=}LPK��C���,Uȕ!!�T�3@wl^&�P��uxv���A�\V�����e����漢{�MQb�F��x'ߪ0�I�׼�1�[?��E�%\��TX�mO[I�c���m�d����-�>����A2�u�N�^dP�ҹ��Ck��0 �?o�"�+��ˬ1�L^��C��%pӧ���vȸ�q�YN	d�2�0�M�L%��R���3��xB��3���J����`(��
� �g�8��JL�3W1�kVY_Hc�6��,��w���$<�&xl:���jg�_���d���l:��h\�9����dUl�y-��<���3�/膱���o�L��ӏ���U�T�~),�3�f�\*�dy�����Z�M�#�F�)��nKTh�9z[���(ֵ�A��{��Jͳ�	K���ⱦE�� �Y�6U�L����4�!��^0�g55W�7� ���j�K���_��^�����ʦǷ[��8���ju�%�|;3�o�owx�J������7	�YiH�_
��|,R�l�đy}i�%V�H�58�)_�/�ܑ8>��Mbcd�n�V�kn�slo�ʥ�gW0��
O���x���!�kG�9�7xl����|/,lEZ�ǆ�@�xO�^�A/0
�=�iX��Ҡ}	���AEmٞ
dr������R�c�����7*{�0������,_i�M'��*�$q�Gq���w~�v�#�8��,ix�ё⇾'[J����tKT�����j�>�'Z�#FeJ߃ӧ��Ԅ���8_%kL�ɘ53ķNn��`^��_�8�h�tX��
%�K#䷕��r+��-���]�vwr�t,ю�0:��#����ƼrCNP�~#&ԇ�/��:��u�f',L�:w��aԔ��6�s5�[)�wM��M����a�Y�"3�z��L9�?�&�^t�/E�OHa3����D3S�R��(;Q�<[���q��\
� S|���Hxdf�cP;;����D��8�L�����VzRH��m��w�S�/95l������-Q��Eo��'���X�/�Np�&�7�./���k̘SH.(��0,��L)����A�z�v)KɁ~����^�g�_�j�J��hm�K�V[�|���"����X���.�0x�jlT��V�V�`;�<mh��ڇS������Q�=��.(sk��3 ����}jd%��NڰM�O� ;B=Ge�K�
����>O5}5�
B��XOL59N<��WAb���
�5og4���Y�:�d�y�\v�W�\�6o��7�1���w�d���	�����ՠ�Ӿ��&�\1�i�v��®������mXm0�r�i��ړ��Z����������hm���fQ]�ND��C�O��&/��-=�����"�	�I�rN�DS�P���W�bEM����B�(@}�Or>?r����f,�#��d�|g����a�/���*M1�!P'	��LT�Z�:�&
�q��^�Rl=߀l&�҇)�3�s�����k�J�Ps�xt~�8&fڂ.��8K0mW��^��!@�sN���@K�zjy�9�M�{��1M�|jѥ�`�q����+�/>�M@{gM@OKp�N!'�6!�[rP��4�?(/��:��o`�4���U��'ɜ�,�yrи'�HZE:�|M�4.t ��V'�N\إ��Y�}2g��Ui8=F����p7R�<��Vn��6��"3s�؏�(Q�����5��֦۟(�`��J-��c��@X�j�6����;�,���z��"�.e�BE1W#жE��(z�b!�����p������Bx䧰�kT!���ʸ�+G�������0�'���u�/ ��i�y*�g����;A\��.@wI�3��hϊWj�iν����+;Ўl�==tC0�D�����>y�v��'��^P}�	��Ca��Ȍ╁��T�����^�)}Pk�Mu�[ �B��Az����L��Z�.H�qLF�	������`xh���������&3�[dl:+^%na*�K���,�I���x^Z��S|�A)���07��C�u:�<^�9��2�3ѣ,�!����"��7�y6��b�^�+3C��p3�w���4k�Y�.K��{�0�Jd��γ��x��E���غ�
�*�d�tJ\̩K����S�`�х��6J�� W�y�V"��_��e��\#�f�w��$�]�Æ�9l��L�ʬ�_5��d��]�����Q�9"���K2Ql��u���ra��8dƏ�'k�$9�$�~a�'K�&�%3#�x�'Ɠ,P�N�`����$F \����/4������eH`&o��et��.cS���8
G9i�6�Җ.K�S^�E�
O��I�uOASdA��Kv��5k7�O��nڃ��,U;7M�'��2$��q���;���Ϻn��,_���GIG�������?�j�����ss�>�>u�D�J����9�Ժ�:�.h�k�b��Q���[B�V�c�����SiX�,�%����mK�e����� �ԇJtߓrP����R
:��*�a��`ery���~��P�D�C���:ҹ�Q�L�%���N����)J�y_��28ٺ�|Za:��"i44��8�9|��&_ !� ��%<�O�!a�Mp��_r3I����~�;��<�������6� ��O̍Hn|�g�;p���zL^�.�Lf$k�}V�@H��nm`�?���9k�9��K��p�N������k�歽E陵�pF+O�-`��Y��YS~������D���X��#�A����,����xG���>�]I� /b��9nm@�VQg�^��N�+x�裫b�����*�� �V�;;�l�hV%�������[�Q�7W�q�i(���)���`H}�*����C˕ռ�GB�����yo
��4��*�}� �Bs�OB��N�y�Ww���D
�
�ɠof�'PŻp)�d�}`��xW|l�\
Y|�����L��1%��ܪd��1	5wg�1����"���Tg:�1d�Kv�'��K�^�nj��;7�h$J����S/�3���0�r����G
�]�y��2�ŻX&e�x#5�=�6u�.�	ĝrDk,S�0��x�3��ꣷ	d綦�I��W@�Br4���Źy��w#���rI��Ԙ�����`s���Pݔ^��VZ�����wq�"`^C�*=}�&�EZ��a���C��kw&��_sc�t��<&\� �8�^�WN��T��!�b�s�2�U�@�p$��M���g w�r���ŏS֮�q�]w�D9��!jM�����A@p��'j܇��Ƌ��0?�h*��=���h4��ZU���'?XC,'��yh�D��������_����|�P�ĸy�c7��_RS-#����ְ��Q�*�q[����H�Iӂ�m�՞�N}�q�fD��ǳ���E&L���t*�#�������Zf�(�K��x](�r�� =ea�9����8�]�=7p�C����a����^N	�9w+R҄`�������y)����R''�_m2c^T?g�
 �U�	,�l���,^_ˉ��t�t���q�g�Sl+S����_���Al��� !tвp�i��2�1�?x/��A��܆&LtS�Ò��ɟ���a��&̳H]I�,;�|�(Xο�?��R5,��<�m��,|�m�<!�6���(��Mf�4����i~|��q�c�9��q��,ǔtƓ�l�GU�P$[���6 �l��s*�3LM��.����Di��m�!xP�`�3֩i�rj� ��Ǉ�����n�M�/6�J6�   �  {  �  a  �%  u.  �4  ;  UA  �G  �M  T  ]Z  �`  �f  "m  fs  �y  �  /�  o�  ��  ��  9�  }�  ��  ��  ��  j�  ��  ��  V�  ��  ��  L�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl��@��- G��D����H��I�H���9��ɥhp|$xun&2�v���>�VE�1zMl�2U!V*����-	H�<)#($�I!��E��%�b��G�<)���
5DU@�O�>5�U�A�<�BĀ4A��E�E�<^f�р�jҹ(!ў"~���f5d�w��׌Dc����Q�C�	 w�Ը��*�g�TXq@b�L\Z�
OZ�9�!
%Ių�@O��3"O�����l����IA��:�"O,��tWS��T�"
��e��=i��|b�x���π �u%l�8=,$�g&E�!K^Б"O�]2�]0!l�%�/I9���	Kx�����$u�:�[�o�j���"D�4Q/OLp@�8��X�a��q��#+D�D�l�8d�EH��J�]�
�P��%<O�#<��)�$-Nu��C�ȫ��c�<!#ߨP��H��)��t)�ɳ�*M\�<�K�4F�Y��o�W2:4�`Mc�<1%�{V�Y�v�>�*�ja�'��x�6OΊ���A�%�xQ$�
�y��<�t����!�^tj�����M3
�'����熓E����bj�d�~���'D8�K�a�BH끣.X�j� �'�ub�"�<9i�9��bE=U`Z�	�'3:1)r���S���р�d8���'2��9�gS���أɘ2]�+�'�H
��<��r�(?��3�'�^��'	A :=�MK�S� �^���'�N��$-��w&�����{��y���;��,�tk䗱B�Q�vD�7h ���ȓ|<��%聺S#r��!����T�ȓ#�T<�s�ױ���4W<���T��@�������C�S��4�ȓm��yɷ������N*<�d ��Ic~rI 8s�L�p&��;|�q�М�y`ڨ5x�	��]*j�ؓ� ݦ�y�iŹg��h��)@��
y�3B��y�E5U�	#5�� @J$\)S$ګ�0<9B�	!w*~`{2f�5��xr��T�"�LB�/#u�E���h�fU3��<a�0�`��"}���,���A� ��-�N�g��EX��O��"J�	�j��7���B��,��"O�8��7r����Ѣ\(�*B�y�D$�',,\"��[

@���`�Uh�ȓ��'�=[��Mj7�Y \� k �4D��b�N����\�#!X�g
�(�F&D�8*7�E�	L�}P#U+A�&���F&��<��}Қ|�"ܭ#;|�1埠O��DCP��ܐx2I �y�p�)Sd�VuR�@�e~ B���l
�Kܿ."�Q9A�57��"<����?ᓵ,E���D���I
M���5@&D��1!a�Xʴ�8#	'<�tq+2f1��=�S�'V�`C��/���p�,Xݾ��ȓ�y�N2AM�ȑ��/\$Y��$bz8*3ˋ&=��a�B*�F�H��A���uN�kW��v�(E��'=B�z�S�9���ӡ��q0�ȓ1��2�Q>�����H�! |e�ȓqh�Pp�!��&�s7� ~gm�}�����&��j�v��u�<}ln� *S:�y"!�3;�u��A�7m�L�p��Y������Z��m�U�ҜQ��c��Ҧ0|JB�+��dX�o�=���2�J� B���|u�u�8h��I0GmJ��2��a���}�*X�&�u�ȓO�a˖K�>IbȀp�6a1:)��8|��Si�{\���A�D�]&��ȓl�fLk 鏍�NxpGBŉ9Y���>y	ד_��D�"�J�X��1H�k�*d�������2َx�X ����L����ȓ[���N���h��a�q#�@��8����(�H�N�pD�	M	fh��ZD����D�E�F�
ύ5t���Of�=���C9�2\�RN��GI�����{�<� �,@`�D�I�`��Q,��43�"Ot*����?{$�CB���8�Y�"O(��à�1WeHF#A!$���"O�4�a.�,e±Qv���� K`"O s�ƞao,�h�z�zZ�"O����/���o�:XF�����5�S�ӷg�L���U�03Y��-*T�B�#��{�*	�J�@�s��C���C�ɀppT���ϞmFe��V�K/�B�	�9<	{��Pp�v��s(B��B�ɣ��B�I�	&0p�Pe������D ��`��]��eϏS)V�㳆�gX�B��T��tx7J
�T�~AۓdN\n~c��o�E���O���g�^�b�y�ġ�&i�1�
�'.�E
�?~P*�� �E�$��
�'`�0�ѦIh48�0J�Oj.��
�'�L=�cIQ,K%d ���[�^ώ��'iVqɆ�|B�xjS�\�Xlj�)�'X�5C"M\~>%S� �?r�ā�'p�ؓ!�"C���r3��DtX=��'A����̐Z:��n����
�'\n�I�B28؝QsOs�E��'e��X�J�����(�3e�⩻�'J�i*�/�r�B(i���Q�'�"\�a��
t l�W蛻28���'Ʀ��E�Wy jtɁ�R�$��'�ԥ�'�</[��K�U�D����'���e�4+�K����R��	�'��1�6B �	���ˇtb���	�'��s�̈́�H�hyr�����293	�'K&�⣌N9<�n��<b��i�'b!�KìHVxA�*H.^�X
�'�`D*���qSр�EH#̴[
�'[$�qD�K��&X���-���'�F�JU�I+k7,�"S,f�]��'�\��k2&d@RD�B����Q�&���-�,i�,xg�"B���ȓV����#�
�#�B X���>�Ni�ȓTV���:�|�C3��VU&���( �F7�S�j�O� Շȓh���
���0� C�M�N��L�ȓO|�1S^�z��{�E��BTR�ȓ\$٩���i��	[�ϨA�r9�ȓ\�֭�4Þ�Sot���[�1v9�ȓX�p��c��e��Rv�yy�Ʌ�+����"�"~�
�B���I��R0h!��F�<+�~u�+�;	H��_v�h�EÞ,�-;�	�&����,��(��	Lݞ�:/s����1���H@��C����Ԏ�'I��}�ȓE@ ����_L��b #1�t��0e~��e׻kL��P�H�)$bԇ��< S���90�ƩE�(!�e�ȓl-h�i�n;@ Dh�B拏"J��O�P p��E�haC*X	v��M��{\�����!vIΌ�m��'�0�ȓKl����_# e:��d��M��ȓ8��!��C�`��e���}z��k� �6 Ě3n��!&�2�|����N)�t+��m�����2�E�ȓ_�F�S27�&X ˄�j�4ч�l�����Ή|` �c��Z�R�b��ȓ*ɖ��e(��U}��E����8�ȓ�h��H�Jf��e�����e��S�? `p� �6/4�9Fo��x�䌳�"O�0�١2Ҹ�!Sl���v��V"OнJRf��nk��y �8z�L�!�"O@x�U�C�I\�t�C!_����"O�\#�o��Cǰ�pa��!���1��'�R�'S�'�r�'���'�B�'��\����<^�$K���S�R<��'�"�'C"�'���'I��'���'�,��@�Wg@��C�G��j����'�r�'m��'�R�'5b�'�r�'�bl���a�ά7���=���4�'���'���'���'�R�'7��'��@��I�t��y�M�:<D����'��'��'�B�'���'N�'�vq��6�����o�3��{�'�B�'���'�"�'���'��'�\T��7tJ�HS8#�zIR��'���'^R�'B�'B2�'�"�'�=ٷ�J(y,I�@�L�H�8��'�B�'_��'*�'o"�'ur�'��h�e�����R�G�u>���'��'��'|��'J2�'�'�0�z��2%$y ���
Nr~qc��'���'r�'zB�'3��'xr�'��D��"! �Lݶx�����'2�'���'{�'���'rb�'lX�B�[~J��i�!v}�ݹd�'72�'���'A"�'h��'w��'9�����%�U�],�M�'P�?1���?��?����?a�-��'�B��WDX������߾c�˓�?i,O1��ɰ�M��J�+~�\1e�E�G|�'�A�%����'�6?�i>��X"���0��U���W�c����sk�����I�Yg.�mH~7��8�w�i�)gDh��й����ա21O���<��i=��lPa�D(�r๠�؝-*�nZ�zb�(� ��y�υ��=f�:TT@�2!�|�"�'u��>�|��AN�M�'l�a�Z�TE���#\4Lb��'���@���i>��	(q-Du�(1}� ��D���	gy�|"n���D�D�ff�Lg��<XҪ!�F���Xuf��[�O.���O��IR}���<C4h�
�hʉf���`%�����O��I��1�����t�c!3--%l�K�+� ڬd��*�<�-O���s�@ L&MH�}K0ϖ�-/���eOe�J޴w	F��'ע7�0�i>���=�����2qY����w����ߟt�I��}mc~=�~x�S�+X��DƔ���i`/F�Wm�<��'�H��BM����'��� �X���'m�Z_& 3���gz�G� �S��Lp5!�4y��F!�&tp"�ZM�M'j�s&Ës *�"ƥ�O]�$ �P17�Ќ��h��3�"�q�@�;��0��E�>��#��5 �ۢ�['�`�Ej��'�ri���G�'s �/\�*��q�u��?۔��d�^#d�69K��P(c	�ӓL��S�$+��x��VLOi�<�Eg��"�=c$��Cn� *H	^x�AR�^�O�r�$'�le��@EE/3*��[5��WF��j�OB@���bl��֨�����2Rz�ha���Ȼ��i�6|�� D��p��i��=��;7��8F?*(����(;U��:�hd�??�([`�� e�:\*@$N�ـ�ɂH���?����?y��>>�.�O��dހ a>�R@�;.H8���. :��	?N���fI�c"zP{Пў s�F�%%֢���N4B\l��"`���?���G��l���eO�c�3ړV�ç�*�
(V�ې#��4���3~��2���?�S�'��S�l���m�����l8��)D���ao��tO���$�Z��K����HO���O���;����xM�g�\�|4���#D�0��ÅF���E��>gm0'�>D��b H� ^F��3]s�����<D���d��^��="��Z�({f s�;D�d��!Ä}Kl�e�����Q�):D�֩F?�>�vE�!7X�T��j6D�${��L?�H�X���
B��t��*D��B��OăѠK�B/� ��(D����fդZ���B����7'Ȥ�FL(D���� L:}�� ��\�����%�)D�T�"K��vP�`aCZ bVV̂�(D���RA�LdF���+Z�c�I���8D�(õe�r!2�B!ǒ�Rz�@)D���뛐L��L��j�M*C4D�����i�����]r��S3=D�xJ5K��@�t�F�fM����/D���4Hԣ��qF��U��>��B���1Ѥf�422�L��L�>,nB�I���h� �%9�S��^�B�ɧp�5kgG*
���DY-z�C�)� 
���`�<yS�10U풋}�h9c"O�%1����x�3�IO7�8�1r"OP4hc�28��F�&����"O@q삕R��Ŋ�k ��ޠ�"O���$���N=��'L���xz�"OD��D� �@�+'f[�jx�C"O��)cb�%-��S�0�%A "O��c0.�#�R�ض��M	2A�4"O$Ȱ�D.6Jt��rAZ�L�Uң"O|1�&�� ��ո�ɕb�P9�E"O���@Pn:\*`�0̮�Qq�<\O�hBt�-�X,�V�i��H���'o�i@p͔9Q�@ s���:��ܱ�'[��LB�I�>��9s�S��)1 �o�h"?Y#�	�k��~Z����d���V ���y�W�K�<q�� @3.��%��W�&tq0B�C?�u)DQV�� 3���Q�9E�d-M�di���!AGr�q�*,�y���6�=[�`S�r�T%SI�DY�|bgIo�m(Qƍ�$J"����?#<9�;$�r�;֥Y��zd%�S��<���ٹx���8p+^�`�A�ÔT��aɬC7�� ;D��|���-l � �J�w�,cf����Oz���Y�^��憌�%LL��9�T,x�/��,Q��qܼ|)�"O&�A �Q�m�	�ѫO�0_�)4�'t�� [=��	����&�C$� P�r�sw퍊{O&����
Lc��aJ���"N;G)��%B��p̀P�ʾm��� U�#D�R�	0��)^[�'Pj�٧� 2`���Q�"�4V���k�),����Z�q{J������<�w��6?����s�D--�\L�%œ>9wa|��2R�|��V��AԺ�K$����hO΀q��
_묔jo �.d�h�ߟ �C��(+��)��I��:���"O��hdG�=!H��f.	�8���1#7O$����(f���C�>s���F�t�ѽN3D2���m��\y��ڼ�y�j��\��Y��GJ1 �k��f--�q�o��I+�Q 8�"�sƔ?#<��ɛ]�f}X�'�*���QrA�z��(�$n����k�C�QJ��h ���k�����_�V�:��LY�ư>aP��kvf	;�� 
�)8E$R�'��q��!��`@)E'��'3�h�CGg7ڐɃ�Z=|sl��@�0���ț��:� ���y)Hy̓_
�X[��+ 	�钓��' 9�?��p"ώ"������3��9��"D��ɴ`���� g��={�8p@����x�	!26�݁�ϝ#G�,�g�'���٤<Q"�o����[� a�@�qQ�d��fŜS��;�����]�xb��^�ᰇG&R^t��_+�HOZ`���R�H��q��+#�//.
I��#�i�E��C�l��B䉂<�L��! J3{!���V���&�B6m�)s�Akb��sӪ@�ǆ�n7�y��#]�P)R�"O}afD���XƊ�:���:�R��2�'���{rf�|Kr�҆#~�
�gH!��>��V�O�`�N��MȬ�����"[T��Q"O�mHC��<|JЩ�CF�&@@Q$�	 1y6�#��)D#3��<�6�͵jR$�P���n'!�ě�T�z���b�.rK�=Qጎ/*��BBs�Tm�=E�ܴ`�fћp��K L I֮��� ��D^`(�V�����D;{t���'u���fG���=ɀ͓�PP�b-@��z�K��kX���
���x�t#�}���b�C�ۓc��y��2Z]<Y�wC�Nf���g���hO��k��F�r���Hc��9��E,ٺ�e!�&<�0C�	*G_�|�`M�/P�q���Ygip�+�|�P#���_N�ӧ�|BeTYoJ��-×5mt��QÓ��xBmD9����gfδ#�<V\>*�L��DG� �������$LO@m��cU��bM�}�&P�5�'�8��d'?�1 �61$��"��c?�\���Vz�hi "O����,��� �j��ws�$Xc������4���K$ ��E�D��0}E�2U*Ӏ<��u��'�y
� ��`s�!@�\�P���V549���Oh��
�}Ե����<�Ϙ' ��H�D�&^���ϤM�Z��'���JR,��g3.��v,�*���y�AбjE��d���'�j�P��҈H� $J��5E��(�ÓFE���(��,5�At@W�4�8�r� R+E6D!��t���I�F�9P7�՛4d�Ұ*��d�w��U�����H�8�u�'+�'%���'�W#avH�KU��;�()�ȓF,�CT��~���SJ��b�D��T&�y��>�)�1����ⴤ���Pk����Am�����DV�7O�Qi�!�1mh�:WH�09Bru��J�lЛ�ݿg
"OX�.�Ph!�J2��ቿ��y�!	C�e�6�A'C�F�N�?��I�LI���,D�8�'V�+���"�T�}��t�hI�U���D�"	@�أ�X��0>1 iͫ�qs��� 1�ѸSk�x}⇋#w��+ܴ{5��1$a݋F����y�Ok�aJ:
4��G����4��'\��sc �?�Դ��C�	g���ŭ�w��1�@=?9�3O�S+}��r��p��];���i[���(�eD�B`��$�6����a��BX�(IjsB�s�$^���ϓ �ţ2/�'�P����YGxHP
E!b�u���rM�}�2�R#��OR)���<i��˴a��a��8��+�&wR��)Cf�cG�1�c��]<2mp#-M|���ἰk' D+d�vؘ ��1�*�A�Z Q�;OP��Q��,���'���8O�	���Sm�X�ȵh��W�z�!��<���CѠ�	��]9�f�j�`����<��̵s���~&��&O��X$.� Pl6�ɔ6���dP3�7挋X��|�5A���	@cu~2c2�I�Ҿ#<�g�X?A �	�3H6J��ܠ�	]n�'F� �D �q��Qh�����)�/.����@_)D��i�W���������$Ѓ�V\���L�5O�`Q�ᅸY��I=京{�"N�����1�s��S H���y䪒5H@�L��g�CrlC�	0s�����V*���)C%�` 1��L1�y A�2�S���g����@H%m̠I�̘���-ܝ ��'dX���BJ�3�B���טS����c��`.�97'D�]�x����'ʓT����e�)*Z�jVLӤMC4F~���(m[�IS��E�"&l��l���)�L��I��v氬��"OBl��߰gl`�,B�\mR����̦��b�>�=	��6
gR������y�c�9 'LC�	9^��ѻ6fL/$�:�b�Ȩ:�8��!#�+��'Q8#}�'�6�u@P�< �m�DH�!�	��'q��3t$Ͼ;6�8e*�H�9����iC��0>Y /��#(��O	�1�Xݑ�Ts�����=9K@4͓~``E�sͫ�T���?&@��r?�Y��K�h���`�n�R�U�>ك�Ħ)U���b��bs $B�D9xf4(d�;#MvC�	�`�J�AAdC �\`҃ �F0
�;T�6O��F��O�o�~22�&b�eg���"O��2�O�{:�@p5i�L[�T1d�'��帣k$a|"�z��8�
I���)W��>!��C�F��dZ�8�J�h���9[�)fس)O!�D]�)f��S�-&�.�;CdȐ@I��H��ߤ鈟��G�$c%faIf(�
2p-I�"O|�a�M�8�j�9�gǳ{9�l!Ƕil ���!�)�禅A�Xq�%9 CX�n��zU�-D��`QiU/x�̝�s ����)T��>q`�D�c�a|b�4~�,��v(�[O�]���,��>��9�L�dԈj)�4P��Ӈs� l3��I�!�d\9B#$�p�e��S���Kݵ[ӑ�ܘ2��q��#}��/��\��F�FJe��Nt�<!�_�n��C�T�����E��	�r�hb�"~n�22�乑 
߄Ve��Qr��?V|�C�	��P�e���P9����Z�ll����9|Ozh��d�K���K�G>z�P��'tN�+j�ԋsi��;����P�ƧT���2D���r�.B�p���F(L��MS��4ғfVM�r��y��r��0qD0�Ƙ'�jC�I�[=�t�4Kܖ~����W�q�7�שN[��>E��t�? 8ȸ��Оz��a�`.��T��< �"O,Yc��<>t]a�!�?C�6�R�����0>!un�7z�`�M���r�+V�hX���S��	�yR+C6=�t2��8\$nͱF.��yJ�b}>��ŸML��&B�3�hO��� ��3.�Ѫ�ɗ�iQ*�iM�Y#�B�	�l����\-T� Y����|I�C���f(p�$J$$����b�I�K��C�I�g�d �BD��t�$�ƫ��C�I�
!
,�AjA�g�,1&�E��B�Ɂ#�Td�����l�a �5fzC䉿O)X���ƚ77����	I.�RC�	M���$�M.U\���/ƸhDC�	�����F��R	���΅xC�I�}��%{�c�.w�<Xq��D�	�ZC�	<!^�L3��ը9�Z�������B��y�"%�0��0h+"����}ߤB䉯X�|yأ���H!ʤZs&29W|B�	�W�L��S� >L�ly3�@mC�	rd��_�c�X�A��(z%�C�	��)��K�E�h$����4=0�C䉂=�M��G�3_Tq���q��C�ɡ�x�'ρP�H�&�S�NC䉔7��<r�Mk2-R����D��B�	�vk��q�O��I�Ȍ T֖��ȓR��L�`_�=*������Jd����%
PA8��Qz�ֆo�D���"K�] ��D^����-cr��ȓ'�t���
�Ej�(��ɋ�d�|��ȓ�j��nZSO�$H# �#�ry�ȓd��؀��Q�T�� (
�s�V��ȓ7}��+���/p���
H�z ���4�ʷ�\$��ͪӃ��s���j�)���iȜ�� `U>���M.DM�6��E��=��P��6��! ��^��<�����l���X!�h&LP�#��\A&�[�Y�X�ȓ ��Y���|��Hё�<f-�ȓnH|x��
�8���-� lH��ȓ&�SQ��"G�� GnYU���lqdY��W6;�j�Y�oA�fp��ȓ2[8��D�q:��j�&����k�T����S�I b	���Ցv钥�ȓ�\h�C�T:F� '܄X�ȓ.H�Q"���B)�	��ؖm�01����Y��E/@�d	{7ȅVM�!�ȓ:�<| ���Qb�L�6����ȓ=����O�A��9���.ai�ȓ)��b�Ȫ-�NECW�[� ���ȓ�0�Ԫ�-R���m�]�$��":q)pHɪ	y4p��*�j3���G����&���ulF1#��-8Μ�ȓ�H Z��
|FdS�LM�z;\0��=���Чĉ�EL�3�ƙ<����i�l�'jIs�L����|��w��c�,�*6���W�GG5�@�ȓ};&9ѕk�)&<�5.Ց��Q�ȓi�I3��\�:�T�(Q�#��]��v$ tY�E7��H�O��x�ȓE�`]	��U;*:̲seWv���ȓr�Tq��7<s��J1O��ن�dj��`�U�:˴��5�9������l�\P
p��w/���)p.��V)D&3�NJ���6P�q��S�? ��
 ���]�0�$k*���"O<�{�L҃u� ���摉Lbfh"O�]#�i+I�P-"�E�
b���W"O�t����i*���4j�SyZ� U"O*�!��4Y��T�*L�0�ia"ORP��nR� ��Ź�H��%B �"O�Т4e^3Ąl`�S�l��Q�"Op#��� w���T.��RӾȱ3"OX�wA�,;���h��+lV���"O�Dˣ.�_��e�:k�t;C"ONe�Q��ty ��D7�i	�"O�Ř�`��)��e��;N��1�"Oܜ�V*@"8���P�	� fD"OR4��,W���P�`[8[��0�"Ox� Se� t��Jā]P�а�"O�����"�ȩCB�n�Z��A"O�<"�Q�Y`и�^;P�N� �"O���$#H��ruEI�	��f"O���l	�ARٙ�F*_��i"OD�Z�J� 9�̨�h�r�֘b"O�:��r@�`J%�A�~�h "O���⧏�)TX,��t�be�"O�X���!H��"Qc�A�`�	�"O��h� V�D�� ���H�B��C"O�y�G��D� 
�!eQ~d��"O�z�o��y?<�9�f��!G��;�"O�i� ԏ"TyaH�P(:��"O&ˑ!˥*R��;�蘱��"O��)��eRN �(��6��d�"O�rp�^U䀌ru�_3U�`��1"O��Sd� ]����'5��t�"O4��
�<f�����5�H�W"O���7��I��XaaE*�$�:V"OKK�"���C�A<NL�t�<�y�+N=P�	IV�%7,����y�JR,r���ì�'��a��yBW�H\�=�CᖘP�@���`X �y���i�����NuQ�I���U �y�
�����*f�]�A�Tۂ&ȩ�y"/
$6	RQ���c��G/X�C�Ɇy��D+��R0T���s�VC�I�lG�e�R%��%>��)�
�JC�	�8y��&h\����։�%vRC�ɷt�����N�_	z�j���b�B�I>:AX%:��7^ �6N�p!�DC�l�䴣a��8`>���L�>j!�3NTFmgZ�
R�\x�Lɑ18!��K^<B;��R�z_H��s,!�D��������yR�|XŬ��S�!��I�n�@��������G��>B�!�d���4�JP�����e���g�!�_�A2b!�7� �`�揞s�!�$G"Pd+T��0�B��Ňh!�D6߼=ɶ
Z������I�Cf!�dR��ɺ�dܨ;��!c�J.8�!�D� ���Zg�,���!�B#_�!�D�$��t�YP!�5��z!�dH,���2ŠI-C��=hW�ة�!�E�.u8ɳ"�/]��1����h!�Jq�@IR��®7G�T2bCZ�xr!�$O�%� ��+X�nq���V!�$B�����@�Z�Rh�P�J�u<!��7KQڄ�� @5A�D������.1!�DIC�� !E
�=Y
��Z0�'^.!�� �E�&	 ck��{���b��@[g"O���m��9>�Ix�d�y�X��"O�kaM]��8	G�^_")��"O�l�d��-,�:�#�^\L �#�"O>Ш��63zZL�"��('j�)"Oh��w!�:$Z�Y𧞺`-P	R�"O�`zjvU���=Ouaf"O���Ê�K5L��Q� {���X�"O��X�"��7�ĥZ�ަd�ڌ�t"O�x��	3d�s�R)5�r� r"O�H��LH�Gm����$>��u�5"O̸�G�0T	�M
�WŤy0�"OU� ��/w��I�D�����D"Op���7fN6�p���-�@�;�"O��"�G��?&|��^C'b�%"O�Q�C�%n�RQuFD�ԂS"O\�J�RaBዧE�S��"O2���\=5A@8��g�kq>�x�"O���ۣv�)!��G�dW��"�"O��aǊ7M
zqx�H�#(���E"O�<#� ��1���FQ� ��*O(A$c�#`������M�q�<b���Ψ��R�ǏY���aND�<�#Dҝ	xԴ{W
��n)Ň�e�<A���"h�`!�֌	�B����V�f�<����>:%�=���
t��"��v�<�bAK����b����~e�Um�L�<����?K88Q�bJ7b�$� ��q�<y&�h�hѓȓ�(�Ldbe��G�<APf��l���˰�� ���{�<���Z�Q�}��)�R�	�ny�<I�	R�2BaxQ#]�x"~����Gk�<�Lʽ#��yH�@�Hb��O�<�"dR��6�v��rW�T�E��O�<a"C�)
. ��ѤܛlZ��T�\W�<1��] 8	|�8�m�n)�)�V؞T�=i@ףnzQkcE��=
ϙg�<�����l��ֈ�%Πx��� a�<I�i�:��3���.J�̰f�TZ�<!W	�:��ش#�Cf��i�R�<���:y8�ᇢ	t�����O�<����B�|1Y��F��Qm�R�<�3)�NQ� r7"��u��dA�_E�<9��B[�`�����#���UL�U�<A`艠0�T�;�%A�\��-*�mX�<���%�I��έ2��@&�z�<ǌ�X�ԩ2n@&Oy<���q�<I0C�n}n�{օ��C��5R���A�<i�gX�t'�Ps0bԛ9�y�Bd�<�U��3H3���U"�"
�J#��h�<��ָ=Q�Hӫ�Y*�(�EMYY�<Ɔ�0B�`�`$MO�@�:��F�QT�<i��A��T��U�o������O�<A"�H�.���7"�ql��E-�I�<�EǛ}�8�ѫF:��[���G�<y��|ǜ0i�J��_�Z�,�j�<��C��{¹���	4w�YC�gLc�<�ï�:Q�^,aW�u|pX��VY�<)Po�04i�CV<�&IX��A�<QA&#,)�څ�^�B�\�I��2D�̊�����}�3!�\ 
��re/D�d�h�v����$�8r
8{`�,D�dFa�H2�0K�+#���")D��r���lw���-����&)D�� �!�U囥y���� �Zl0��"O,�B���[�fI�O��B���"OX���`��im4�`5�4.�L#c"O��[��Әob6�Z�V�n���'���#��˛,Q�@��ϖ8�hT�
�'V>���øs�j�����4d���'~�	ElA���%�F�D (��'v̄�cn��}A�0�����F���'�"ra(^!LD���4
D�i%���'�JY0n��^.��/tHi�%h�y�a
�ěh��P��h��D<�y2._4CM� V-ܽIF�y���_�y�nC�>���%"H�CP��R��Ԓ�y���S�m�F��@X^��b�<�y2��0<���P�\�&��� �H��y� ��e_j��!�:��e�0�yrI..^	�Ăʎ����ׂ�y�/E�N��`Y3��p BMJ�y�CϩOD8�� >�vt�����y�H;	��ت��"�`��r����y��ң4���Ui^�[����M��y�ԝg�����hmbcĊ�yi̓0	y%Ȃ�`,���nӉ�y��o��j���	���
G��y�	>y2����&ЇE%+r)0�y�
2��cf�W��f�X�'���y�¼C��HC5�L' ��b`'[��yr�jظ�yd��D�E �Ɲ��yr샢l�T<���*R֐HR�L��y���%C$Xk��4�T�������yb�هj���#⪚�v9����Γ��y��� lƂ�	e$۷o<T�a#���yҨ�%	�$��0L�4V�Ph��+���yb��P�`���HA�{��@Ra$��y2Cϒx�'#ԊKȑ��HB��ybl]l�7鐞H��˲�=�y���	R�!;�(îQ��}(B1�yb ̼J�$�Z��ܱF@晚��ʖ�y��T�<R�w$�=:�Z `e��ymT.?�q���2]��ѧD��y�M�����ᖴ��@wNߛ�y�ĐNf��D�y��x���ȅ�ybJ��a�> �M:v��8�0k��y�`�taxp��CP)F`�X�뇜�y�c��ǲA1���u��Ũ���y��5W��I��J�$\.l�R!Y=�y,�<<΀ �lQ�.�c�M%�y��Z�P�!�c�=k�B�zď��y2ēI�D�C���):':���!�y򦛇jըy��I7�*})�K�7�y" +$��{ oV+zA��P�y|Z��	6���q�ag"�yR�M��!�/�����JU(��'9P��F�}>"��ύTˎI
�'��i���˩�ܰӰe��Ja����'�����H�v��s�MݺX�����' T9;�j�=)�m["�ŢU����'�f����q�8�2#�
Uw k�'6�A�P�p}zmN�I�
�'K���r��&i�he����M����	�'/\!)�ђ��hU,B�L\�	�'<��	�
S��2�R�eh��	�'����$)H�̓5��*d�Ƥ
�'��y���}#zٻ�I Ih}���� ����"|"g���k}�4"O*��pmЉpW�E9@��`��"O~,�W��K@Ƹs��C�e�2�cS"O�y�1�T3C�����	J�-�6"O���̒�r h��3���gu��i"OhU� ��=�F�1'&ޖq��l�"O&�i���g@��AdP=d���G"Oz��FG�+㴥�6�{��{�"O�Q"酏6�~�rDݸ�*%� "Oh��T��6�慨�%�rǢЩD"O�i� f��f ��*�;M�=G"O�5��.
�K�<i�i��L\�e"O��S��U�v"P�����]��ؐ�"O(���ϐW}�vN��-¬��"OX4R�OQ�Z~�M��E�|��a"O��ɓg�(*ִa*���#m�!�F"O�x3����LkQ�7]�.}�E"Ov0Q�L!!y��3�F�H��	k"O�(��Y�A.H�	�o�5<�b`�`"Oj�R��^�"~9����L����"Ob����� �֌b�GI��(�"O&�zFB��]�F`�!ƙ�m��H�"O�T��SuT�iՏ�&X�"Ov��w�M]Q��!�ۼM���ل"O4 ����u�cE	�x���� "OT�JQ�9ʂ��3i��q�FIhW"OvEA잞:U��#I�9UՂ�j�"OX�Ju�K0yn�}0��ϥ\�J�)�"O���M�V��e�&�e�u��"O�|��GΛ��A"4K�jYx4"O�Xj\1}�1:��T#e�6��T"OI�Sd޶]���Z�9�d|s�"O^�cp,+E9 �Z��X!O�\��"ON�[��M�~��u��fH
Ae�a "O�����]6�t�FhH�{}���"O@��B��֊+I�)+(�שs�<��@:�
l��h�?m���\u�<9�
��IĄYU�
t��t�2B�u�<�7KKir����FZ丗,�q�<Y�U�9|8q�Ԅ J�r��u Uo�<��J�')z&�sh�2��m�<1�i�1*�9��1lz�{���h�<����|M���w��8k$D�[-.!���+�-#��N�N��bk��X�!��5Z���Ic�^�H���rgi��!�$@X��SG�kߴ���)՘R!!�R/?R<��bhH�dҬ<Bj�2!򤜋@88���p�20��/? !�ĺ5w���D�m�z)ÀH��Z�!��Vt���S^P�+� ��|W!�$��zol���O� �ba��O�!�DN�����6� T���p�
7�!�D� R4��D�5K8Yaw*���!��D;�r�����HG�E���L�9o!�N0jZ\����>P(F�APi�6jy!�N����.
��!�ӈAh�!�$�x��	���%M� �B�g#,�!���qђHc���u]�Ѐ���!�D��S32���H\??L����DΤ+�!�DG�K8��$��cF<l�͚LV!�Җ�~ 5�ݵZ��8VLJ7S�!�D^�>b((�G�RmJ�R�+K03�!��Q���W��NQ�$�p,��s
!�D  {1�-K��=`OΤ��aӏ�!�� d�vEO�F�B*�
X�z��B�"O`Ͱ*@f|3��Z;!R�`"O@��%�	��Y���Ζf)2�"O*�*TF�2�8����ڈ3b�b"O�0��wk^]cå[�r� ptgFp�<y�d�!:3�I;f�Mr�
��g�@p�<����9(��)�!	��t�UP�<9��G����	{c��WN�W�<Y��Y�S&F��!�4/�°C�)Vo�<QĆY	N�p�%�� )��A�k�<�MB�M����fJ�]�(p���m�<�T��L��QJ@�9��p[���P�<y� Z����!+P0X!:���NM�<�mIb@Dpx`�#[����t�<1� w��c��6�nER�%Mn�<�v�W�z(x%����J~N��s��S�<y��TU4m*Akڝ4_����$D�Hc`GX9E	�Je��3 �VtiI"D�l����7 (U�alK�cy�A�B� D�葦���do�Q@�቟?Qp`B�.?D����f�&rq�렯T)x[N�P��(D�(�B ID��7`͙'.<j�'D�t!R��%������~�$TP��*D�d���&в!�gtV`�  �)D��3p�(R��A�]�5(��Am$D���	�� �1[F�N(3����� D���q�K����e�&l8��Rg>D�XYF
/U��Ka#�>����=D�@��$J�&+~0����bqC�6D�<"F�0p�\ "��.)�H�D3D�4��' *n�PJRUt4<�1D�h��3`�)X�o�6L#����,D���o��R8�wkˊs����"�6D��(��V4�P�Ah��OC�aHP�6D�$�uC�XW��D�-URu�n4D�Å�^"m���s�N�7z���/ D��)%��',R)���#��=D�4Qf��'��"7�R�S_�� %1D�;�	�!|���0��M_�ȹu�0D����wF> #X!t�b&� D���I��c��9	��+6Ny)�"D�1"��D��˦��CFA��M,D�pz#!ݿ3�5�T�2i;8���*D���gd�3o���䬄#Mp��)D��`DŶ0ڤxF��T��I��:D����%	Uh���W!��H�ȉ�'�$D�4؂CM�_�<T�&W@�t��sg"D����@>N��|�d�dG�]s#�%D�����U�-�f��C�w��{��%D���2�M`����>�� 4@$D����H�%�����*�,�H+E$D�lP���$�(�F��2��0s�'/D��P��ī_�h{��ϽP�H*um0D�H!Q��w�=�!��#�Z�sGB0D�V�ա2�j@se�
' �<��K!D��)D�m�4��'�|���=T����,��Ԥh'͠<��q�"O�azR��6���+愖h�X@�"OU�c+Z�<����
7n�4�{E"O��R��%s`��)�,{��5��"O��+�'q�(�`��^�֑�v"O0��cH��d�Zp9�� �̬��"OPd"G��7FD��.��N�PS$"O8��7m�Y3�H��J]��u�"O� ��C����RA@��*~4��"O���X����s�Ð _����"O`� .�B��-�S�Ү-^��"O�Q���	��EM ��"OKߓ{F��O8]z ��.�y҄�o��L��SF�@C�yrȋ>bL�咣�){���J�̊/�y2o��f�� �#p�-A�&�2�y"i�hf,�6U�hy�0K2g[��y�aμ���3��·[���e� �yb/��Uڐ!]�&n����

�y�(_���l�愳%AD��R�P#�y�Aƌ'�D1���қɶ�KU	�yr��4���"��<j�x�qc�]>�y��={S��/��s.�xK�F���y�Oߪ���؁�q��<9`$�y�,�(O�(K���_ߊB�DJ��PyF(X̰4�E�b����aEH�<YF$��P������dh����A�<I��9:g��7�C}��q��B�<1��_7!�D}�� 
;$�0�G�Ss�<IS�]�,=��1�F�sCl����r�<yF铃X le��!�.�����n�<�ʚ:%���2�A�&0�YR�^C�<y�`�4��@PFN#!��h���Y�<!T	ܾ���҆�!;l����h�S�<	�%�9�$h"w�Ѵ6۠�GN�<Q�/L��V�Ë&欂���G�<�Ï�	�*<`���
&��SRB�ɇ%T����U�*�j)۳j���C��:ފԳ���6dq��z��C�!,���1��1t���K,1��C�ɄKN��r���i鸡�#�KB�C�	�E�������
���"FH�A�fC�I�SϬɂbKֿR��y�f�>�VC�	14`�E�;1�]��m�<n[BC��?[���7f��-�j��S-�a��B�#vԬ��ݦd���r�ɡ=��B䉒r3�� ǂ�,���g�c�B�I
���d	^��Q"�ǅ9��B䉞+ :%���;�d�J$�C8�B�ɷwoxIpCfA�{�V���`,6OvB䉁5l
���fB��P��G2\�RB�� w��}9!�H�4�$ E�c�6B�I�x�~��f��Nٶ�z��`��C�I4�4� ��*%z}i�*7��C�	�B�na�R�Q�D��� "Q"��C�?q��s��؀��cu
5��C��_fDM���>��\�RJ<�jB�I�\�P�
��G�@At�ɐL�;�B�2Lƈ����/�-�ď�WK�B�ɕ:$��7⓯*�x(0/q�B�I&T�����l�����	�ct\B䉔�pQ���O����h�?#�0B�I�u��%��0Y���Q [0�B�	zB�c�J�(M�E2�A�
تB�	#`��PO�+>ژK!j�7%�dB�Ɍ$i���Ħ
5�(D�s/�J 2B䉪�����J�8)�4�am��<m�C���L���O\�U\�1Al[�-��C�	�`��#
��T̪)ؖM�� C�ɥgb���b��~�D�#�7q6(C�I�bh�`A��.]�P-�6hNc�^B�II��(��?)4Sh�b<B�)� �p��ѹ0�<xFHڬX�	p"O>���}, `A:�,�U"O�8��3td�1H��4+�\�c"O��ɱgF�>o0P�ϙ���@e"O�`�lH�O���A�l��h�v9u"OR}z��['5Ʋ00Fօ�֕"U"O I��/�sɾi�����J��`"O�����,/�愀�p��-y�"OZ�e`
$5&�c j�U���k"O��w�@�'A����c�e'B<ȳ"O�l+�(�=j�H�H��c	б#�"OlLӳK�Gj��� hI�Ya��!"OV��4�ج}zEˆ��SJd�"ON�!D�͵7��銳��,0�"O�\� �>*�b��ٵ*��܈3"O(H�GV'L�KG(���&�z�"O�`�%�?<�L�#ΎU�0��"Ob`c�A�)0�	��T�.�p���"O�=�R41��0NU�02""O��y!��PmQ��ƻ���C3"O&T֨�i=��j&BՒj�h�Q"On�:���\D�,�)&�z���"OND@p,�C��Qp����z��"O����˺_�Q�b���z�Hv"O2᫒)��i��0�d���(��uۦ"O|�3f��%F�ܤb$������3"O��Q����ؙQ��"�
�{"O$1�3(	!�0=H φ�7����p"O��7�yS��X�#�J�v��'%D���n>[#��@�Z6��Th�n!D�t�th&	>�%)����q�.����;D��1�iڠe����惥x���+��7D��o��v
�匃]��j��:D���t���Lw��X	�=θU�T�4D������#%z�U��tXp�k3D��1��7a����eV�L=��>D�h�e��8�JXckƃ~\6�&�9D�,���ٿ6dM	f��S�"�I"M,D�,@1i�L�D��ͼA%��7�-D�|:�@A8W8���OI�-�(�#�
(D�<`6�Q���A�5A"A��k9D��1Ń�d� ���B�{�$9�M4D�P�F0�U�pn�2+k����'1D����N�a�x�gV�j�x�x��4D�(�&+P�!�Y��T�9U�2D������<`,cF��,e�9;j6D�t(P��O�rq�J��b���2�H5D�t���ΛO&�X��삲ֲ�($�>D��p&"�nT$���FÜx�����;D�@��ս�l����V�E�n�!�?D�,��G>�xk���6 a�T�h=D��s҈B�U��P�+2B�9I���'��
7K՟s��I	2�G'?��!�'�����,����U�����L�
�'Al�
p�V*( �X�w�8��'&<�u���N�0�2%��5��'����4hU�t�:��'��i2����'�Ih�.@�:�f���O�\�ԭ[�'4�r�@U!R�Uk�h�OѼ�[
�';ޘ���_ QmH1�
�'<�,��	�'f�k7#�6O���b#`׋f��P��'>��س��c��C@)O"�;�'}�X�H�tĤY`ˏX��LS�'�̀91�A���o�� NJU���9D�� ��iS�Խ8�(�`�T���u"O��&%ơ:됰c��_�4����3"O|�3�Q�*Ф����R�J����"OFp��e�<�%�#	�<��"O�d����Y���j�k�?/�F��"O�e���Z$J���B�����"Oޤ�%��� t<��
�_�`���"O�0�v�˔d��١��X�L�y��"OV�����9��9۔'(5����"O��'����A�韕o0L�5"O���a��/S���"�؋t`�e"Ojy����4t5�ȓq�)	�@�"OJ�琮�v�7D����Q"Otј%��� �R�+O�d4�1"OF{�eȽgצ��g�̟q�n�E"Oʬ@a'A�r�(�@jY:g-b�"O2�P�)gj��zGC�,	Z͙�"O�Q��d&w���i�_?r��E"O:$�"��qnpI�%��7���"O�2�i��=xN�0R`�9#��	�"O��&��"<�i�eL98`t"O�Yw@�.F��{���,(���"O�S��L����l$�D���!�� \��KBlIF:�(!�F"��
���h���!�dT0z��鉠��=���5ȅ�X�!�d��$�f�E�6���BA'�7&�!��L�V����"(F��p��G/\E!�Ĕ?�Հ��3LRFl�B̆�l-!��9�@�AS�1<��C�D�'!�dѱ
��� Q�9����ʒTn!�Ę�V�5��.G+`�m�$g�E!�0y�= �ƞ	k�
��%��H�!�]xrDi��h��q���Þ$.8!�f�@��%�@0 Ap4&ա8!��]�#Hd:4n�R-|���DO�o�!�,67ܨ�JVj��骴dZ -�!��]�>a�C��-����"�[(!�� Dh�k���8$9�I�v�E�H'!�$��,oV��6��7<6�C��Β;�!�D�>zސE�7N^�o"���͈�at!��Ƕ!��$p�iW�A�VĊUcQ�'!��C�`���P2�X��GDy&!�  #�,i����(��E��lG�F�!�֓^*\Mk�D')�b��AL�^�!�G
�F���Ã�p,�%���!�Đq�,�Y
K>F��lQ��!�d��"��x��-z
�ڇN�!��.�d�"�*\R��-ͼ#4!��s��(� nI�x��E�d!A�r"OJ�0��G�jB�����6����"OL(xsEE�q�l�g#S8D'N�u"O�����	�-|�hQ3b��j>��j�"O��R��)dv4$�"��2���"O���N����gM4 �΅�倣�y�O�#��T�&����`���tW!�dU'6&Y�4!�*s��ٺ���yB!��-Z���mlЌ��'��'@!�$ț�֜���_Z�\[���h�!�dҬ[�\�ʂ
�2U�x�a��T�!��o� �s��$@h\����[�"�!��.�2��g�A�cLU�o��!�ė�?m�z���5e�苁n��H!��)���8�".X����� {�!�� r9P�L�U��*�mU "���#"O��!J�:~��!�G˔���XjT"Oڌ��F �1"������J�Q��"O�-qTEE�q�"䅍Gz@�"O�aQF�C��w`�;	��R4"O�H�P�I	������;���"O��� -�6=x�uH���*�>x�6"O��@�'� $x�q3v�ǀK�\!rR"Oh+�,�2���diT�J���AY�<��,�������!M,g^�8�`��O�<�JT�s��Z&M/�L!$�c�<��oB�h�G�0^NY��J�<��<:R$5K4�&V�赡�f�B�<��昴��[B�T$�%�/?D�L���?�<���VF��� �>D���wG��2��̘�T��|��<D��i��ƃ �X���E -wT���%D�IP�W/R� E��&w%�b�O"D��9��(Fb�уunN�|�Q#�g!D���&L�S205@�A�Y���	�/*D� ��;~�A�O_� �����$-D��C�eI�|��@vN۷
�jA� D�`:f&ׅb�<�iG噌uw���g
*D�0�%�ARjcW&��_�:�Y�&D�Tq1��\�P2�g�*�qŅ*D�H�U,T�~/����_5T$.)��,D����Ǣ58�H�򪜤�bu�W�+D�(�tAJ�M
��XAM�m�M*D�x˒��M��afȞ;St��;D�(a7M��ps�P���,kz6]��:D���	�"Ԣ�b�

<S��0)��9D��B@@:S�19�ݥN{����e5D��`v"�'��%P�ʜ�Nzvh�5D�d
6G�yF���x�2$�'�1D�XzBB�*`�e�1���G�$���*-D���1��;��q��9^�H)��.?D�H��-��Z ܽ�G�X\�t2ul?D�d1��$:�Lt�5��?:��I��/D�0�d*��Si��F*�Z���+D�PgGF�7t$E���?K�j���(D� a�+�6G��Y"ߓs�"��M#D��䏺K����x
�t�EI!D����^yC.���ƚ���� D�t��JH3q�L�ᆨ(j����D$D�l��%��<�	�� n����#$D���v�+�rͳ�BP���H$f#D���&Q4s7����΍92� 4�"D�И��^��>=ꦥ�]��� -$D�@Tn�.#Rd[�נG�����G#D����@Õ�ԛC.3'3��H�!D���6�
��� �p+I�=@�=D����/��H�qA���n,VuH�i>D����eR�.:�p`�^�P#Ǐ)D����
q�<�a��U�X���O5D�d��k��xt��z���%N2��%f.D� ѷ���0�Xq���B�Q��A7D�T�ai��b�zq��W�1�b'5D������H�Ta*[��M�dh3D��*P�L4-���'0���K��$D�C�fA�J�P����� K�PM��8D�	�
�T\B��`X�P��8D�����L���4����m1�5D����.i��U��uY~0Ŧ(D�(�D #;��ȑ/�^5���!D�� ָ����'F ����m˵6��"�"OPɂ����J�C��q��H7"O6X���^�1C��x�@�EX���$"O�1�k�#D�͸��Q���!"Orݙ�*Աh��Q:3�X��T�0�"O8{�h�Q�6����5쪘Hd"O���L���H��Bϲ���"OR��f�/V�i F�G�
�@%"O�eQ	T�u�P4rEg����@q"O�IaD�!�f8�I�%p�	�f"O����/��_@@=+TBK?���Z�!��8��T�� 	��-#���>/�!�߮E�X�k����(''�
o!��|���e��7
|�,97fL�ZR!�$��g7D8`�eq��K3��*3!�R�6��9p���,Vܰ��Cʚ�!�D����:0i�qM(��֡�h�!�D�v��q%	s�$����!`e!��7Vp��Ј��R����T�)P!�d�d^�%3M��: JBL�M@!��I߾8�sK�Tfܐ�@�&!�Z%h���:���?U���d�R<E�!�	�_��  F��
Q[*� `P�b�!�ۨ`����Vd�hKHā=T�!�ύm1�隠�]�P?�� �3�!����������F1�5��a��u!�䐮G<�P���*,��Zu!P�[�!��H�<�j�zCFۖ3(x��b�7E�!�@vW�,xe-I�oz�!� ~!�U�M���*S�˰`f\�Q��.]!򄓝[N�iu���{R�	�Y!��=�04�M�EIąs�b.(!�dDQ1�I�"���,�qT��U�!���WvH�a�*X܊ՊݸJ�!��! ��SÅ�����Ri��0!�P`��Ңn�i�TDI�N�)"2!�$�%\}�]z����zҴ롇\?/!�$M�E>&AD�$�R��%��o!�$�2	��U�̿z�B�k�_(k�!��!3���� �LQ��CȺ�!����0���QP���c�!�d׌QO\:`�ˮ*��y���F�`�!�$�`ϊhX�d\�1�
lXu�6!�đ�v6���b�&��Sg��3�!�$Z�q��y��2\������=I�!�̯4�u��K@XHpIc#@6WS!�D�2FK�hR�.�x/��y Ƙ%,!�dה�Ҡ��K�jL�i��. �u*!򄂇������_�YDh��oƀp�!��Z����i�0!���N��'x!������ '�ѕ �Q��	�VO!�
	?�`��A���9�g�J	d;!�d�K��Q���@ 90��l�!�DI�LZ�) �d5�a�ŋS�f�!��4�rZ�f?g���Q�ʞ0	P!�49�`@ g��.<NPrǦ��m.!��Wn�ܐ�J�&D/��#�e۳"!�d������cJ9F�,�����js!�dA*[>|�C�$���P�,�!�D��<s�I��hDi���$_d!�'���H�-�f�]x��QU!�P�6u�`s��G-��j�Oe�!�䄯Y�m�7)(���.�3�!�D�$BHb�k��&9��q,Q�~�!�� �L��L����;��p"O�P�"��zDv�r��Ϻ%JX;�"O`%���Jt��̣�f�Z�~�"O�aȲ���x�&A�SC�< �>|�E"O*�)�i�u("�nzV��"Oz���D��jH��A͢E�#�"O�-�E��  Z�"�p͢��&"O�y�6�Đ\dT�,�	!a0*�"Od���Ĩ���7�@�X<`K�"OR��AuJ�T�Q��1Q #�"O����S�Ȧ�����)�"Oji�	Q5K{& *�) ���[�"OЁ���T�J� �[��w�
�7"O��Ѧ�YiV=�d 8��dCP"O��y��l-p�1煖�z���e"O���mO'-p�Y��-/�Ep "O��G*��%���0�$^�Ռ��"O@��'@�04Fxy���V�\�"Od���&]	*�:�k`hA�Rل�4"O�����7XNΉ)(R�l1�)#b"O����"�3^�h�iG�D�Q@�3w"OrU+P�Դ�@�$�K�h���R"Ox���B��ZӦ���艢J�t�(U"OV�SG��G�B��&U�v��q�"O�%�DF�.W`�Pd�5cqA`e"OD ���:(5qY��n���c"O���Ȼe�¬⃊�+�B� 0"O��qT/�'`7���	҅$/$a��"O%��`S~�*�0��_��U 2"Ol��eF��g�@9�����!�!�"O0���MCd��@ ��A�n���"O���AO�+� �	(��0��"O��0��C�lE�q]�h�N�+@"OD��ǌU��jUB̴(�{�"O(� �cR�eU�!8��
, جh@C"O�t`R�̰�\d����Y���1�"O�l�6�T
c�􀒸>���3t"O��B��C��H���M�bW~�B�"O61	���?&�֪��3D� 2�"O��ůö'��`��R15.��"OZ�yd������+ɂ]~��"O��b�)׹0,~MەM�U���0"O�t�f�K\���0��%Q����"O��j�e�o"�H(��B�6�X �2"O�̪5�ց-���J� ��p�f	�3"O���@H�&�$YR��H� ��C"OāV@!~���� @��h�"O|���a�& ��8��:;����"O�	�`�PUd|�Х��lJ"O���h�4S��ܹ��C�q�и�F"OXQ����.:�.���H�l�H!�"O�eCC��7oB���.[����"�"O�H@���>�x��	�O���"O�UTF)�<�:��u!�,ٹ4S!��T(���bfu�PA2I�]<!�D;`�2=A��N� �*�"+�2!!�d�����9�DI��M+�
{!��&�j��!��Q��i�	�8�!���1@���6��2�`�i�!�$�-$�{ub�
�aIס�!��7f��#�UT�A�a�`�!�$�F�D��H�2�<���/&x�!��	_|����h�����/;�!�2IFְ{�)�T��0+&n�%�!�� B�C��4�h�rf��:ʬ��v"O䩉q��4�NY#3����l��"O���F�^���
Dm��u;3"O��6���\���� �F����2"O(�#����^�%	�*�,q�D"OHȩ��)&���)�	�:UN�P"O���P!A&!�|%(Q� %+8 +�"OL�bI�X�n���hA�rʨ�+�"O��SF@�.4=BPh��@�u�����"Otd ��91<�+`fYx�bli�"O�ijNN+r�0UQ��\?���4"OF%��i'�Hh���;J��I��"O=[veQ$]���1Th�\����"O�@���c���`��	+~�ѕ"O"����ߺW�C�Z�k��|��"O��T��"y�.m���Ҳw��� "O��XFǛ�0��T*u��&|)<��G"O
� �,���4�QH�qi�"O�p������`G\�e�¹�U"Or�0f��;%�����H�?���P�"Oj�CEA�4,,���!���0�"O���Aۑ 3�Hɐ�"Lx�#�"OL�pங84�����"�'n��qx�"O�{��ʫ{P��y ǜa�Y��"O�$#"�-TRh��e�_�r���"O��f�܅)�������܂"O�jaE� C � 5u֎�I�"O���S,�3�H��g��>c0'"O�ɳ)��7��	b��֗���b�"OȰ+��Z!T��( ���a��A��"OĹZ"�Dcd�@7ʅS�V��g"O.ɰ�ؼo'}���@ j�|}��"Ov�c���[ôdj�kP�G�p�a"Ov��e��_މr����K����$"O@uQbLK1K��h�@�$z����"O��!&�w�����i�=\[��"OR}��I�&7f��a@�S�*��aa"O���ee�u�H�d�)qî�a!"O0�s�$���-�lM�h��-��"Oh���	5������k��0z�"O����T(ʀ<b��ӑ�2[g"ON�SI˽|L@b��8ϐ���"O���ǥ�L�z�4
hF%�R"O�UI�g]�j�*���"d���"O��"����YS*���"Ot�i�M�M��	��^M!�"O�Q��Ƚ��kFi�Qަ�Y�"O6��ҫQ0 ��M��ٟB��	Zu"O@eY�طRTP�2H��N���q"ON"�F�gmD��G�9��1S�"OiK���*+��I�HF	*�dE1@"O�8;�����!i�k�.¦"OH�� ٣
`Mzb�R�6A"On;V�9U'�ԛ#`L0P��Ѱ"Ob�����c��Ё��U3�D�"OjԈ�|�̔Q��0#�H�"O�YS�̍{��p��ت9:���"O蜘��C0b��(7�Tx
B��"O4��5�M�G ų�X�3�ԝ��"OX�*w)ջ��m�%�Y�P8�]�f"OaXՅ�[Ν�0nީ���"O��r�%_�0'h8pBJ�P�)�"O�(�͆p ��
��f8DU*�"O��!���j��2I��y⬫�"O� �t*^�ZWX��ХE�E<m	�"OHst�<=�HC����"O`)W� ��m��Ò�V��)�"O�1����a
�1H�cV"� �"O���M�a��B_�(�f"O�-�'&�f�TqQ�n$t��(03"O�������,�1D��7��Pk�"Ot��A,!�h] c`˟9��U�""O|D;q�+�B�(eE5L?���"O����A��]�P��6F��?r�B1"OF��AA((���cƟmJxJ'"O�IY�O�R�B�{����(���"O���t���$���L;>z�( "Otّ�	"bJ�}����)����U"O����S�qDh=)j�'�$��"O��:@RT4Ф�P:08=��"O�i㒀SI�F�����%oZ59"O�4��ZX*ȃ�	T8Z0��"O�4Xt�(iU<�[ �R�fhJ(6"O���m��M��u�TŞp&�R"Od��2JWI*��Vj�P��3APz�<9W�X/Xڼ��K�d�9��M_�<1�Q��A������@I�e�C��+]�;�N wX�۱cȣ62B�	�G�0�P"!�	l����GI�"��C�I,͒,��`ų`��d�!�[#q�C��4S�>Uk�J>�Tؗ`�5DC�I=p����r¤�HT�8{C�ɺ�Hh����pJ8�2b�ݰC�ɎM��U���)#��RSO��K��C�I�,�rIѦK���MR����i]�C䉡Z�Ic"�U�ũ2�|s�C�	*P@�JF�7���a�mtC�I�*l�8EH�$�̋�ˌ9Z��C䉘�n��E�����i��bPC�I�$'��jb�p�D�EJI�d1 C���aJ�k�3��ۥʜe���d�L����$��(�vC�?J�!��Y�X�x��NW58�f��Tb�2�!�d_�KJCA{���@��I�!�$U�r��t�#�%4vFuh�"�.6�!�
8����mƌ>YN�����0�!�5$�$"��9FB2y�&@��!��K=y(���X�=N�����!�D�(x�@q��ʢx8y1�ģ#0!�N�U���-7|qB�m�sO!�W"�TMq'*�'{
(A;�&�"J�!��� �FU�ªO�m��'lN�w�!���&c*|�ذ%��&d��k�::(!�$P�E��m�pT�]�ȡ� �!��Q� lpD��� �(rS�?�!�D�N�]�Ҏ5=ڶ��0�Z�H!�D�4����2�[�`������)�!�D78�yC�K��{h�a7�P$d�!��i{H���K��각IC�A=�!�d[�#�Au�֝k�}h"�D	%�!�5'-�(��3/֠8Y�G�'?�!��t���\)-���k��
k���ȓ]��ٕ�̒F(�juF�ڑ�ȓ���zA��F�����υLp8t��"�p�8�눉AN&�h���p�ȇȓ爅"V��sd�[E�K: ���ȓbLd�ᡄM;��a���:R3r�ȓl��+bd |�>0Z!)U�
�\Ї�S�? �Cӌ��d�����ތ8��"O�S�N{Ϩ�a�q��a��"O�i�򁘢n]D�k�с ���۰"O�[�BN�'p@4��GY�úăF"O�	�ȓ�7HP2!)ZM�b"O>�7&�6�X�b�h  'J��P�"OD�zcI��Ae��=,J軂"OH5Qtm�v��� �ݾ:����"O�` �f�T����-$�2T"O(8Wnɐ�=sQ"�*+�����"O ˃d�� i3U!ɹR�h�9c"O"��ă2�Nt�5 �p�N|c�"O��0�O�LH�e�/��bм�xa"O4�RңZ9J�ȓ��x!qv"O��ò��]�f��h(dU�%��"O.}��K4�8�(Y
O�t�3"O�Qk?-�x���9�r�"O�aJvaY�a%�@��Ǉ�'7z��"OfiJ��]�1@ԑ����#4!z�ط"O0
d�<'L#�������yb��qX䬁Ң��Q=��Gቛ�y�l�fЀ��b��J��C�N��y"�/�bd�'��H߼��B��yB�\�1V!҉צn��J���yr�cXJ���l�-c�$	aAH��yB*H�
 Zl��!ׁd6��w�H'�y�Ɓ�`0�Z�a�+
�0�Sw�ȸ�yR��xOx}IՄ
���	G�G�yB�Lf,�" �"K�rEJ�e�4�y�)K70��(�b�=w�"��y��F:8��A�U�ߧ0	�4)�)�1�y��M*&6�qC"q*F���+�/�yE�;|�yf`ZminL�@F��y�.~B)ʔÏk���� ���y�?,yP��oC�__�9i ���yr�3^sxpa"	H*'�����jD�y�l�:X!�Q�c � r$��]��y����V-aDD�_�9��V#�y��<��q�B��Z�K��ں�y��?vcrq Oy�����R$�yR��y��YӅ��>���؄o���y��#]��E�G��?��4�# H��y��%p>����kM �	C��&�yr�@�A�|��/�;^$r8q@��ybfI��X�i��}�p� )�	�B�I;_�i�e�]�VP��PD� `�B�	?;h��3�N�M�j��勃�A��C�pQ��3p���v��\Rǧ_2l�B䉙$��T;�C({�\���:٪B�I&{r���B�c�maǮ\�����]�H�"̠0�����j+�#e!��Vk��<+����DR���e�!�:V�v�H���_��'�F-�Py����2%z���7-��XAd�޲�y�0	�M�"ҍ"�H�:4�B�yB��*N\1q"��������y��G�oF��K��cU��;�m��y���`���r�EL�V Y�RIT��y��/9�E1���=�`�y�� ]��W$E�9��$I��'�yBD$�ޙBT�*޶���G��y��
��9�V�B3�%�A�G�u�ȓG��ڶ%\�m2��c[�L"�h�ȓTMf02���f.V  �1t:�ȇ�S�? v�H�v�R�F�L���1��"OD�(��@�U�9�D�2��=aE"O@���Y��6I�^��Qx�"O�p�G�q�YHە`�%�"O��葯�!	�D�� ��I��"O���Iº"b��qgL��}5v���"O�]�4fвbZ�*sJR�Z��b�"O�;��ˀG@ʐ:���cT�I[r"OT��� aj)K�dK6O��aB"O��h�ˇ�|�,m�f䆪��Xb�"OlJъ̿n-  �&#����<D�(Q�Hy6J��1ZV�b��9D�hu'�*�(�ٴ�ѕh��5���8D�� 䊏8o�F��&9|j��!D�gÖ�%�6��C�;�0��&?D����+��R64  �BY �&G>D����ɵ-r�=�R�@1��ti@�!D����ۘ��I�
!�"fo?D�,��+�1t0@�Y���T��P6�;D��9d�a�����/zl���L,D�x���͒��l���N�JX���A+D���C���l}�HC���J�h���'D��@'׎K��4h׍�?d����A�)D����F%$9�	aqj�t}�ģ�(D� B�K$,9lAGf\+.a#E;D��`��جt�cdg��,�ܔ�ga+D�!%e�1J��`��*/���;i)D��s�ˏ�Hl@��
Y_��٧�"D� ����
{��|b5�R��d�R��$D�X�3DĹ7��aJ]�A@:@�S D�(s��#�z	qB��H�^<�C�<D������3I�N` ����d�Hf�/D��`U-�z��*�%�&�0��A/D��qȑ�P�d��D��u7,`'�0D��A0ꗐ(H��DFD+u$lz!�*D�D`5�2A��I��@*U�����)D��qJ�,�HX��݉v4�y�m$D��X3i�\|��ȓ\�R���S��#D���M�E��%��hL�6ɴ���>D����� �pcT���8)^l� �:D��������F-�3l"O�<��8D��Z��E!xw��jE�'�*�vE8D�4���ӱOx����a� l� n6D�P3�J�-+�R�J&���C���A�3D����)�"�,�Rc���S��:�a,D�`0�I#F��G۷¾�z��5D��x ᐃav*��>�D��gm D�H��P!L1g�,��� Ӯ<D�,x$`Ďeঈ��lZ�&P�ز��8D�T����4��M��X ���Vk9D���1F�W.���0��6.�&h6D� kc���*����KC�iXԌ�8D�h�Β�3�D�.����)D���g� /����^�I��۲(%D�����7�B|Ib�t	��J��#D��oY�-	�����E4jBN"D� ������t!C�y�9Р�,D�Xk��?y���4+�:!ʥ��B,D���dH#8��,H��\r�TmR��4D�X�'��g�5:��j��0%-?D�d���"���Hs�,]����9D� �V������B͉3A�X�k5D���4���W�"=���2.hp��L��y�(ޣ/x�|�C�"���o�y
� <�x�"� {lhQq����|ڐ*T"O� ⤉�s�JԨ�
�adA�"OJ1�EJ�:a��	���swvrD"O�i��#V�X!��?iy��"O�a�7ɞ�����K*>Z�!4"O��8$�"@$di$膥XF�=H�"O"�bҫԡKT��Ri�4,1��d"Ovpx��	D�d��U�5�"O&͹Uԏxl�7��%c���D�4D�T��̖*8tsEkU�vn�׭3D�D#�%�15T89���9VO8I��3D���&�WD�	w��9�
��/D��:\�pYi(f.wސ傒$:D���P��\�V�(�"r���E#D�����
�-��傐�E:N�|A:g�.D���r��9��Y tǗQx� ��?D�l*2�J�C5���+�r�� a=D��h�$с-�*�j�+�Ҩ���:D��c���1g6I �A0�X���8D����@D�-�ܵR3���:QLq��4D�ИS-�B��᠒��(F@AB�-1D����	��,���r��ƕ}�&�i/D����P%`�a��'U�d��k.D���!#D�f4��Dj�X�*̫pO-D�<`���yh���Р� ˼��$N-D�<��$b>��3f��Sb`0�gl,D�x�%H�,1:��l_Mx�R*,D��#���w)!G�@�e7 �g/)D�� ���~��}�!(��O�쭛H'D�����!V
���"�)j�j�� D�x�U�8�!s���u��њ��#D���!��d�@M�Yi�� D�`%c���
x�uR�>|t�Pd#D�(�O��|ܰ�,D���"D�I�/U�PZ:х:Ci,��qi D��ZDO�j��h@ S�vt�RW�<D��Pn$=�xDA�!П�*`K&�-D��#�ֈǪE���
K���s� *D��z6J��N��Ts�G
-��)y��&D��q@���#��YX́�e� D�dx�H�B��٣��k�X����<D�  ģ�`��u��*��j ��8�e0D�h��N�A��ku�(]3�;U�9D��Eƍ_Ĉ�j�"Ɇ`�P 	p�<D�����E�'.�b!n�q�x���9D�`�pYn��'AC�RH��7D��S�bD�"��p��1+y���!)D�h��Ƃ9����A�ht�BAB(D��Ȳ��/i���3�^;/�ĉytA(D��I!��/���2���;x��8�o9D��ҳF�� �Xvj)r�Ȕp��8D���Vo&à�'�Èy���4H<D��*sdԢw�]Z"ȟ-q/��0$ D��R��"� 43$@��a�^��H<D�	V���!�̘y��8Bt4����9D��:�4dx���Fd�c(��5�9D���*�*H�P����հm ����!9D��ФiΒ�@xt�Ɋ2����#�4D��`kO�U�̐Y�f��%Vi�6�2D�bR��G���ㄆ�}C���2D��QCj{Sx�	DmڱqT�����0D�8)�ι|c��3�$�2���Aa9D�4"�R��ƥ9��R.St�c+D�D���&7�\�A��K0P(h`(D�� ��hU�޶n��5*�.>u0""On�@�ٰjن#� Hp\И�r"O� �p��*���Q�$W�~>����"O�U��B�Bܑ+�#��c7���0"O�q*�Ą�Rb��b�
B�2��"O��9�#�"37DY��$I�D�}��"O*\i��k���s� �rZ�);�"O4<�vj�k���R��Ha�p��"O �cǃO����ª@�62h=��"OTa��[�<�Vhj��J>N���6"O\��R~|��[b��9�H�!"O @hv�X4t�HlZ���K�$�"O<�Y�A@7>2y���҇ed�јb"O�����!Y��
��
Z̭�"O&�i4�N�.@Vl�6̛�M���"O��1	��)�^��u��qG"K�"O�4('(��lW
��
�?.D�"O6�G	\Vh��Y��� E�FE �"OvE��D�>�6�bR(�,xv�k�"O�b����.��ݸ6�?ld��S"OD��`�^�i��)iY�T*�"O�H1A�rpe�r�Vx�X@�p"O4|��D{�ʭ�D��%e�:��s"O��Sfe{5N���B:_�n<�"O��� +����TGp�ƨ�f"OL]ZS&ޞu,�h���8�\L'"O>�T�ћ�*��'�_�k_4��t"O`��R	��.)��J�oO�	4"O�5��
�v�jl� #ýe����"O�XA��W0�+�F)G:8h�"O�ȫgE]&� `$Eڠ*1���"O�%�QE]/S���h�Ա~���"OԤ) ��ej�����[8{�TQJ"O&<�5�[h����,�<BD
 �"O�Lf�%;=���iZ|� =)�"Oz���ÄU���,Z���S�"O��yd���,%�^�V�h�"Oᒷ��Yf@yI���Dݠ�"O�y2�/(F�qP��R�r�v"O�E��L�%!��92b��D�ҵ�F"O>}y�@������L��J�"O���C�j>���!��6��"O�!p0��9������W�p�"O�y��Ξ�pI��lL�2�����"O��ʡ� ��T����;���"O�a�'$�,Pld���a�n�ЄYe"O�) WݒbRę¡�.�DApt"OR�z�WN[��\��h:�'���:p�¥fI��� �/2����'��h�.��1�Emļ#l���'�`��j@x��cܴ)L=K�'��@cV��$|�Ҹ�b)Ԓv�0:�',.�q #$sTX���Y�eu1�
�'�ND�����T#Ag��[�z0�'��A�7�]UD�Ы��)Z55(
�'�l]Z*��2'�>K6]!
�'�`�MG�9��]�r�ޔ2��(�	�'K*��S,ޔ҄���&[��!	�'�����X
mqΕ)��ֻL��%��'�f˔o)h2�A�d�T2Whyp�'����GF� �DI����u�'NPd�#���)�
!3���m�!j�'dV)�0�U�D��Di�p!r���'R�!X�d�O�D@�d��1�DdP��� ",�alHSv���CGS��P�;�"OT�i�kÙ`vܐ��2���0#"O�Tp��+h�<�:���8a �"O��`���:��D[Dm٭$,�a�"O��)Q�\/)HFh2��Jv&��R"O	�` �>�nx��:m
���"O
T��X�{P����˓BOf���"O��{��)`���`���?+6����"O����N�{�P��eߐc���"O$h�l��H�JT���R�.ͼ��u"O� Q����p��wC(=cT4�v"Ov���iK���RC��$I���"O���e�A�f9`ʤ,Υ3��	�"OB��G�]�)�k����P"O�Dӂ��:~\�แ�Z� ��h��"O|u�7�Z�b��� �m�	^����"O��q�(B=P���Yw�L��2d:g"O�I*#���3�Z�D)�"O΅#�Iֻ����G@�9vx���Q"O(y �B�U�\Y��N��w���""O�m�7M�ƞp�v�̲zrH��"O���B(��w!�Ld�^6Y��pj�"O�ıuA�3�:T��K�@��Ʉ"O�(�p�˛L�\�eR-H�}��"Ol9�3�F9o�x�f��1l�Z�07"O*�����}�腛QD� پ��R"O�"d�H���#�C�5<#��ar"O*�#��L&p"�V�`�:"O����� ?�jA�aK��R1�j�"O���F�je �ӯ8x��؄"O�D5�I:�^�ѕ� @�b�H"O���2�ȎQs.Iq
L�q�8�""O2`I�À�e|Z��B�X2b��$"O����U�&t�ܘ�Cɡx,�"OU�t-A�x���K��v)��@�"O�=(��pɜ�1w�UC���B"O�1i��K�r�@���4(�"O($i�C^�<�:�q�*�."�Y��"OLi���}�%�vCI��@�A"O������'w�Hg��@�*��W"O���$*�p�2�M�n��"�"O�pUbM��D���?38E��"O��ғbݪ$J�*bm���"O�m���\?
����m�d��Q�"O̔@'f� ��3���	.oh���"O���"�,E�2�x�kX�9��h��"OX��$eT'��48��	'O���"O�	"E@Cw?ܹD�?���"O"iɢ 
GH� `DHB�e�"O� �$ݹ@8���e�}�^x��"OX5*w��z�z�!B#c�ʅѱ"O��hR��|����E@ 8r�a��"O^}Áa\5J���R�[�GN�4�"O8����,w���C�8@�Z�"O�s�\�svz �v.ɏG��9�c"Oܜ��cR�g�ب�-َH�Ft�"O���$���Q�®˖Lֈ� "O^b��A~�<\��-T2\���"O@U���&�`����= >d�R�"O���g� 2��DK4��'��ز"O���h�AizEÇ+YP�9f"Ob$[D�E;6��!�3�ҢNC�"O�hB�\I0�@���q�黷"O���HO��a�d���~�~�V"O� ����C$@�� Fm�-!B��V"O�$�F� /��l��I5Hs��`"O�����"5�a#vȒ�!p8�D"O���O7i�rpIg�R$i��"O��;�k@0?�$2Tg��"�)��"O
���.\>q�����6w˰X)�"O��q��./��A��Qƶ���"O�@���GZ\Q �qQF$#��',�-�"�S�`�%�Dę�:����֎.��`
�'����ڟ<W �*t'�� �ޙ#	�'g����LS�i:�����&}��'iFyK  U3k���`��P��y�'�� �3խ�4-�腳#1�
�'w�4أ��d����J�'���	�'/ڔ�F��0m�NQyEǏ�/�-	�'ݲ�ϔ��"��ծCv��r	�'u �+t�������s�Q6+8 u�'c �֧��c���y d�$-��3�'�6����M�
p��
ԃ���F]0�'�����S7pB��s�B(L>F��
�'*�PZ��Y�.��p[Co�GXP��
�'q�Myb.J�kٮ�����
=b ��
�'��Ѻf��[
�0��92�zmH�'Ԡ)e%��V�n1�Ɂ�b�
#�'k<u�&��Pt)�Oc��xI�'���"Re�[zM��,��k@ \��'��P��T#b��]Q�@O2l(��2�'�L`�/�o���H�&o���'	&q�4���@��jĪo��hS�'����!0Eـ$	����c���c�'��"�ҷJty�j�Y,�0
�'Ѭu	rCW�L�V��ԨןWX��0�W�W\�ڈ�L�Ы"o��)�QC���/yG��W3$���@�J\������-)��[TK�"@L���%ڝ�0?����q'ԥt�d�.�#2�0���Q�D�!���
���4`0�Ӏ[*V���R��V��q�ȓX�8���N��y��%C@Xu�'���'�����C+�$�d�v��j$�q��R )�x���q�yN�G��X14c�vA�Z��Κ5�6�rD�
�B7j�+�Qj��𤟊5�D�Y�j�'Cn ʦM̦�a}�m�L=8�{���@
�褩
9"\+���+�XQT�A�K����3�'��n��1�b�@�M�#WY��*������@�+�DͲ+
T�v(�g��i��~��uÁ%]�IHIY[iƾ�ȓ	z��"L�_\��cE����J�l�/CU\�	�K�y��$`�@+�F�\c��Kf���Ixȝ`�构 j���'G�cA�S�8�s��ʇK�Mx���u���M�<d��`������<ʓ=�,(D���V�*�zf��*H��'�V5��C�o���I�V�H�Ӧ��7gOH�p���D[��%jE�h�dS��'�ġ0�F��b�"��C;^x�<ۍ{�]�=h��ҷ.���
�u�ujB��.?h���'(]bs��4�"���� �D���6�$9�Ȇ<1���q�"�<��x���!;�z�KS�_�B%l���O5� =�2�w�X��"< ��%*D�ʇM|�͢	�'��Wt*4�#OշB�����AM*n38�)�'�<�NIC�l���VӞS�O�%Nݘ���(�4y�]jW�'\���N8M�T�3���g�X�ɗ.E4R���#��A�gTvj�y�\\��~�� 1��ѱrR�a�ɴ"}΁�r>�	?��@y�oɢ
����`�G�tC�9��̔���ԄV�Hq/�f��d��HوA�"O"��U�@.dJ�"	?ATxP`��ҭ[��:!�#C'��k�%�S�.��e� �S�W��n�<_��4��_�1��.S:i�!�DAMT��*���H5��x֍Fa�@�T%�-F�Px��C�`�vhh&K�OR��rDM%�Iv� #�~�PdJC�>Lf��ğ<���xf�^�Mp��Za�T�W
������5&���y6�@�H#r͹��'%`��T����H��t��+�	�Z���QE��|�s.� %2��ի� _N���i00�����2�B���:M!�� ��A�@ �=s���-���d#�a��i�)�Seb���L@,L6��I� 9�S�O0�N�|�´賣pWJ���ꙩ$!���@/ҽ$�h����i�sҵ)�])uH0�жkL"�XM W���A*ܝR�D#�IV|�8q�(Ʋ4%z͂C�E�nT����\��)��ZH홃j\?�`r��]R:�����Y}������v
'|O�iRGOȴ0��5�tI�/'hɉ��	Xt,�;֩ݼ"��H�� �$/Ӹ��Ӹ�R�Ȁ�tH�;���!*�)�Eǌw�<i��2�&��BI�/ך��C��6�"�S�B�+���R�	�<��e�S���y�F��"�d�鐤1�b���Ş#{!���;Q80
�!]�>�*@i�8a�DA3 ��	�k�)��'��� 	�����49!�U�܄��
*�Ob`c3��+)J�h�e�1d�YK��;P���#�Ӥ���0>q�L�Z�̠��f&�����|���ϓ/*8%�wH����X�K)����f/�y�7�̲>9�Ԫ�4���#�}���ť+]L؈6oF6/<��ȓ8��l�C�Ѵ�rX��M�Z�J��ȓ/���oV&>B�Ls��D�1Z�9���.lPoR�H��h��P�h\̇ȓ{�����X�Ⱦ�!�4|�(�ȓNL����h���X���+[`n8��'=>ٳ��+
f�S�M8C�x��ȓ}̦����͓m�k��;8�H���^1�A@_M6]r�F�4K��5��p7\�o��*�x�Y�=���
���ǃt\@-衋ٗN��1��PY��QkV6�u��F
7��X�� <Z=h���/OV$��
:	ir���˄@S1��X�>��q�5-�$x�ȓ'���G��j���W��4���� �� sF'R�`� m0ub�F-��(U����*H4!�ҙhB�C���Q�ȓC�d�u�;i�d���n��]��RJL�Х�H�F�d(F�.*LI����Y@�l�plP �àD�� ��{���(�\�C 
�"j^<��=�l%�smǢ����6�ТSAD��Eb�8���`> �sG1G��,��t 	p&��z
��r��P g�D���3�,��M݄b���a�p���ȓ%���bQ)�6`��R��71�N��rfHju�KC����*p�ȓ�q����,T\z	��h��`��O�4 6&�zubJ���ĆT�ȓ��	�i�s[�YxvE_8��,���RD	�	�*�+����Ej��4D�l���<&q�ܯ	g^�Ht)5D��AmӀPNJ=�c����܈Չ1D�@*��^��hv@X�/*�=��8D�H�!�;?_���k�!�Ti��4D���e)�Ե���D'}�d@� 0D�T�dψ�7N�C!I��j�d8d�.D���_7R�r2��"sdԢ�6D�|)�C[�i4�!S�h9����2D���s(ʚ	r����H݉[xD09# .D���b�NbLJ1iPF�6z�A��9D�$Wg��H���:Nn���6�:D��D�'#j�*��<�|)�s
2D���M,S:� �!!�s?��R�d3D�`[!�)q�T�w�5b�j����/D��P��ӿ�aY�ň�&�Z�(+D�P ��[�ʀ�4mF���x�c4D��!�`.3�t\q��)[��E2 �2D��)���#Y��L�棂N����Ћ7D��  ���^5;�u��@�#]�(��"OZѱ���JA��!�Q�=W@��q"O,1� G]=L�h 3S�߸.�Nآw"O�ဩ.8�x}����HR�"O2$�d+߸}���R,N��"O�\Р�-b�>h0�P.jc܉X�"OP92�³~:��1pAĖwn�52$"O��Ç�$_`���S�\Gvi��"O����:{2�s�( K4� '�'r��X� �C	�
~�R�#i�'>�j��a%\O�@����3�xlP�'4�%Ͽ4� P�L�j���'0�R���\��٣I@@��XH>ѳF��AD��x�a�+dj"}ҕƍ-fۘ���k��v�^�	�a�p�<�4g�u�䭱תO��<0{��3Iv)x'��z����36[�$�~&�x�q욮G�(�c�O=G�8��`a7$���a�60� F�)��Ā�o��!�C� 	lP�2�`���
g,ԧ2�^��4,Ϩ4���qEe#O�\c�R1?��hZ''���ECA�g<�P�)@�>�"@*�y����D����-_M��'G���E_��&�Ό-���򀓉P�>���^�I���w�R�/�F�;�'#D����DǺQ��� B��=�r5	� �+Cb�Su!�)#��s��C�b>&�����F��S��<��t;f&:����O�!���Ug#z�V�;�F
TP�yZ�aZ�]y��Wh;qh�d����AHc��B|�� ���$�i����b��*=8,�Ў̊g���@�ڮ��C�aL�xV�L��-=4�8#O^�8��4�D·�^��;�@*?a�	܎b���C�& �l��B���OD><B!��&�a��H,j���x�'=F�q���'"�DaqFJ*kx�+��1f.Pbb�7g�D�=��Of�'@:P����Kh��P��R"�4���'A<@�5�J8� ��,�����r�h� ��ӈ9�&��(�-��y�aRcv���L ��d���?�0<��)��F�\I$��T�޳�|KqMF ������P���"`�]$��x�wU�d@��np(� ��������0,9r���Jj>U �CC�H6&xq�`A"�P&D��E68r��v۹k����+ŢX@D���iŲ��Ɗ��o�\�>�O�a  �hk��%	��K�j��i�O
��AN�\�z�IW��uA�K�b�L�EIG*o�~����8\Oa����G�Ę`�ǒ>:<���<yt(L	{&���cS�&�i����ʘ" O��(t��È8}�!��"Wf6vHG@�QR늄Y��'�Ybk��[��$jEF�p�OXL(���\�I�C�H}~��'�z �Ü�j�֤+��[�M��9���\2��N�tc"�<��E�4��1�
]��LⰦ�Z�<� A�A�R�K���j<D�)�C���h�:D?a}RC����eC�>e\�K"�G�y"�[�J�P� Ei1^84K�Ọ�y����$��G��B���!��I��y�$�%7�N�Q�ˎ`�:����y��W48f��à��[�AQ��T��y�� �;h��K�I3I\��3���y��&#�v���.I�@l��ʖ�y�Q�4TD��V�~nj͈�k��y��8s`<��b��,l��aXq�y2&X�wY`	1���}��p�ܟ�y���,�0��@u�!���y"O��,r,PȒ
hs*����׀�y���7l�����Y������Ծ�y��	]� �2�OX�Ws�C�ƛ�yB��Q�D	�2+��(�F��y2��$s�hI��	/��l��@$�y�� � �]��֋h�p0P�F��y��W�c6ʀx����RE��'D��𢍄��`�ԉ�8j� �i%D���w���X:Q#��U�,�t��9D�� �#�]E�H(1�Z51	$�[T"O�釧�n' =�@���%Ў�R"OB1+W@�#O�P�f8=ц�"O�EWƎ�eV�p�ǔh��0d"O�];V�$f���k���R�VT+6"O� �lѷz��Q�ŋUr�"O��{0͞Bc�m+�I�6��8�a"O��I�\/U� u��g�uXx��t"O=Y�ՍfbTE�c(
>M��"a"O��x	Q9��Gۏ1(���"ODx��o��4h�@G[)h*���"O�� 2GT,�)U���/f��d"O68�Bl�������E��y��"O�i��ګJ��Qxu�,H�Z��2"O��p/;%'�лmT<q�f\@"O��	1!ݳ!�@�k'm@9#�̀�v"O�h�q��'�<8�j�)��0JA"OL�ȧ�Z!^��(�A(ռI����0"O�ѓ֦�];x��3��7f�
�K`"O|Qᥥ�C�$�;@�@�9`%5"O8H�Wn����t!�*�QC�"O�9B�L�"���x��|���"O>QPC�ҽu����;-��p	4"O�h*��Q�:�4��I^3R���3"O���&�/,����e�;e��h`"Oj�*4���c(�����9�C�"O0`k��7�*�8r.Q��J=��"O�$YECW<R��C8=�fI2�"O������5���`́�%,�9�"O�!���>-��3�F�7]\m[�"OV�0A��+:����2R�"O
���E) ��y�����.�K�"O�qa`�ΐ~v�(�A�"@�tUؐ"O�9�P��5x�����/�'E����"O�ɥ���:�,i sKZ;xt<��"O�E��*R	��+W(ezD�9�����'{F�)���>�c&��E�	+ X7u۠��-PxH<��Ȏr\A�G�"l��<r�J����aG�x�a~�,�f�ܜ�!�$7��H����?�p<aC����ؒc��gy����u��n�"z2��p���y�J�*�LMs/��k0`���#P�����2W�n��C?i]E�t��	{�>�8�dD�=���('���yB�-� Xª��4�aH2�ܾ0�>̂юK�<A�`�'���CK~�=���1����cBG/�B�����AC�?5,Dkt炚b�X�k����P��̩㣃6C}>�֪5�O��դ�&;���pL�f�v�� �ɠ1�~=��)�=r9�1�V���0��72��)��>ؑ�lX* �B�![�P�zE�P֢U�R
��Q�+ʖ�U�V�
ԆF4l޼�:u�2�d	G�\c��a�,,��	��$��C���
�'
����8'��a�'�?jhȡ��);���S���x$�L�&G���$<ʓq���*��D�:�[�����1��I�7����o�@IT�=h
h����2��UY3�\37Ж���A ���|"�ÔL'�MӅi��.����Z���'�DL�GK-�\��6k��HR:Zc�Ĵ���MR/Y�p���(tҸKT(^��y�eX"wG>�PCH����%�4ȑu_�92ׄB�0�2t@	��M�
�a���b�O��.3r�H�������[fNӇ6�!�䘱E��iӇ�(*�%B�G�>tє5$�4t��m�Bu��;��O��Q��Ǆ!���{U�Ye�������S�a{��<Ǭ8��*�L$���-�*Kې0��\��=��y���$퉲n.�|��Z��Hy��Mi���ං��'|`k1�xټ�@�*�j��tSV�ƶ����^@8�j�;d�}�I��PQB�I.oR��(�$�vE�2�R&Vn�I�RFD8�L2����*�6Q2Ef�,m��Z��w�xx#�%C�zPq§�	6s=
Ɂ	�'F�Y:���+5K�y��c��f<�@ذ$�&�2c�[�j2��6��
F�I
��Qi��� 2���!ǆqRБbmKb���r�'v�@���5 �`�T��e�t(#�ܧʈ�JG��R�;m �4��a���8�Oh�UJ�v��S��A��l�&�d߂z�T��+�/Uo�Cg%_� ��� �wBd�/'WHM)à�;�	�a�_l�<�Ӧ�
;�F��)]N���0��M�?dܜ�����A�d���gc���,�Ӛ4���Z�kQ�(�'DD�<�����x�0�'|>�` �Z)(�v��t�!6��̀�'�ּ��R֙K܊9Zө	�K|<�HP�;�H�0�[A��*%����*�h����	�|����P-�2�.*=�C�ŀzx��z���Tl�6cR2<BR��>�O6x�'�B�%,�䓅F��l�[����C�����_�	���H��/	L��O_�[���?X����YZ�'��=	�jB�n~}r�c��Y%h��uꝒs�*LؖAצf>���u���h��$N�T�.�k"���C���K�4u�!�����t�'�U�0<�T��&��D�)t�z���M�az�O$YX	0B�g��9�����p>����/���Q�1��+��̾^MF�B�M1SY�B�IFY4�FU�fu� �)Y�C��UҸ[e���,����@ϨC䉦��m w"�.r �E�µE��C�	3BPyZ���fWu"a.�$AR�C�	.]����A�{^q�c�ȪL.vB�ɟ��|	R���U��x��AXW�B�I�;��z�F�l�ժזY�C��1G|��ᙊE�ޘ�q��@�pC䉷z�h��B�o/��k׆�0� C�	B\����}�P��J֛f_vC�ɑKvIb��t�D0!��Q�.C䉗Y�� �7�58P�(T 2;�4C�	h�f�`�Ώ�N��@l[=Z�B�I�D �fJ/q�،�f!�xjfC�	�Y�̥b3N:o��	7S�g��C�	�(�T���Z,ox�  EP �FC�	T�4�ai��^	� ��C��K�>C�	^�
���k�?@hx08P揺r�C�	�n�4�`cҼf�Z�j��:3��C�$7�D�*�/٭x�40�6�Wo�B�ISFVaڥ:�L���l���hC�� H@�� 
D�X��M� I�B䉜`zm�L̮vx$�t蕹
��C�I��Ȭ���/V��Z&
Q�C�	�Z��)�M
/�?k8pp!�8D� �a/�����H2P�H@r�H9D������2���+��	0&�jTA��7D��h�
�`�b�BD=
�:�c2D�a�C�*]���S �O�(�t�;%D���r�P�L���X1"P��	R�'D�X�F��#�:��$E�(	��1�#D�@r5�Y9Al��qCA�'%���C�O*D�Ⱥ2��&�����8��u�A=D�d���_@j�3d��FxHm˳D;D��b n	���jVAY�-��y!k-D�@IpEڦ��׌"Yn@��e&D� (Ǌ	^;�LxD�4H�>��d'D��A�DYh���f��6�(�A�$D�dc��"�H(�@��S\����,D�����=N��ɂ��g?pǁ,D�4AAM�D���C��9{��*�f<D����!\�9��s���-7��q�qf?D�$x��Y�uD���(ƪ�-*A�:D��; �*'��w),5v���8D�h´�x��SD��;����@k7D��I�Nܧ&�J]����=Fa��L!D�h��"V�+�.\�,OD���+�L D�؊�`#,����K�7.��E�:D�� z�� JZ�����1(y2�f"O�)P�Z1�b�1ޑgĲTa�"O*%!�
�� t#�(��4a "O�}7��:E�tq���>Ua�"O:|Kև�3��u��1耤�t"O��P3�ʤyb+Y*7�D}��"O�L��"]'l`�R��P.Ė��V"O��p��3��8��R�{��ٰ"OnQy�lJ]O����ټz�:(�"O 0a6�U�aC�lÍ�F9�"O�5k�l�2u<�
�R��\-�d"Oy)�F�c�R(Y�i�%PV,�q�"Ot�j�6#x@ف���*m��a��"Onh���8��&�8H����"O�M��*Ե����]����4"O@�Պ�#;ڢQ�%eX�N�j�X�"O�y�r��.yq�����1r�ę�"O>��f䀳Y�\4I �ԇy�
Dj�"O�({A��o��̩�>g�����"OV�*��!tf�Їb�w���V"O^��e�=8�%���BfT��t"Ot!k��!��-�`"&�v: "Or�J���%��X�2��/ڌU{t"O�pyf�^	%�J�3��'u-��`�"O�Q2�F�$M#<踗��?p��h""Oj�3�.�(Q�l���DO�]����"O,���]&C��Hh�l8QF�pc�"ONHC�
/o��+t��y-H�y`"O�e�(Q���a��`��+R"O,�!0�V�pFf�*D��y�20��"OJ噀���Ha�VȖ�e�4 H2"O���A*M�'��G�!]ܘR�"O� �,��I	Ra�x��}�e"O6<��+������'��H�"Od����a�yh��)�.�Q�"On�x&j�2/�M����!��9��"ONȈ�ꖨLm&Yq1*0?��8I�"Ov�3�#�(j�Ȱv�4��E��"O�(Xǃ�M�~�)4	�*-zt��"O�h�w?���rr��>Zx �"O�*'�	n�J����Ӡs�KT"O�R��f
��
	-���[t"O�)�e�3L��I�$Ƀ,����f"O:�ѵa���p�Q��\���)�"O����
� �`���#&�<�"O���b�I���B5H� ig�z%"O�Q�Ջ����P���^�H1"OE����;k�tёƕ�6NB��C"O��X����#��h�`�#���*"O@�x�_7�\�RQ���,��xp"O�ʃgH�x<x��$*˥e��5Ra"O�D���J�yo��:���@��"O���Wt�YY��X�7��((%"O���E�	�uL���W���HVL!�Dgh��Ic匲.~9��d.!�B��U����f�(��T�.!�V�}�$�$�U��ԍ:��V�J-!�%
��U�4��X�*Th��6	/!��T2V�bH���2]�0��r!��M.t�r9P����N��u@
�$�!�dh�g��&���3KJx� Q1#"O8P9�f�RL��!0*0���\�y�$��h	�4�c녁,& 7����yB�H,���@f#��h�j�u��y
� ��@4��.?��5�0�VI��8("O4�U"�/وI���i�@�r"O��S���3?��ѫ,�����"O~�K�'�v��94 � X�b���"O��E`1�Z1�F≒(���0"O�,cP��y�&J�[ �*��I��y��KE<�;�9ydXɐ"D=�y��@9
�bp��'\��E/
��y�Å�n�B��ਇ:�\i����ybꋖF���GH/����Z0�y2���x{���3�-%�ne�çX
�yb��{-�5Qs��$Q�ē�y�i��9�`=�5�<X�*]x���yRlO�9a��qp��Y֎ɣ	��yR�Ӄ|֞e�Ӎ
�]�R��d��y�!��E���%��U4#pi�����H0Պаf0���M>t�Dـ�+V�Pc�!#�I�|�#�[�Ot���Lš({2� g͒g90�kP'ܺl��'�pd ���"��D�6!�d� �2�GS{I����E�ul�&
�a���A��x �ł\	�D`���$P�
pup4�S��)�Y� k`�K؆]q�Y)��mA���O�0ِM��w`��&��}:� �E����Ԩ� 4����"P����*^H�'
F�g�S��F6p� ��Q!�M���=��'R.�
p�4��ɜ��` @ܴ(�:i4��.۬OBq�"H6�)�S�>E$-�7���^����e�G�P��Cd�O(�N1}�'�?E�ԉ����c�!�5AA�I��&�[������	�Z�a�T&�.�d���Ǖ5�>4{SNߐVd`�Z�h�X}⁙�Mc-�x}�j��N�����!t�l�BP�& ���ix8�nՍ\	��	ç.�uӰ	Š^wt�y�*��su0��B�i4����.5�P�b�N��0|ʥ��:�X�C�.�@��k��-
f�W��!IH$i��|J����~ڤ*5Hlĩd	��-J| ��M�@�Y�O��cٴPO-���C���K�T�B|0�j~�V��'@��*�yRɟ���dAxn=a�E��"]�`�G��'� Y�p�'�)擹llvaY"_�G�։yS���B��'������)
����$��#'�H��s�#��I�Y�#<E��
�� �$ �c�d��1RS�#�M�ل���ȟtx���rQR|H��S�!xv�`���'c�=�S��I�g�(�ɔ��
 �H���&���'a�����~
�q׀���M�<���m}�<�Aة-s��4A�"'k�Q�QIFu�<�0�6�
a/�X����i�Y�<it
�{���q���[O�|X�Zm�<) ��
Q�(�CCO��0�@�s�N�<)L��6���Q-��^��{�LM�<ICh�3[*����.�*|�6��F�<	���5F��yp#K�}����rJ�n�<��&�p���0<�Ή@R�l�<q��O�=C���&`8Se�h�<A3,Y���y# ���1��q���?D�ԪJ�M�ԸVl�U4���=D���qEK�0u:K#!Iu`�E�'�=D����.v�x<+G̒�%%LI�� D���D�V�vlr����[h�rg%1D��je���38�BA�	T���a�.D�8J���9ܢ���ؗq��1B,D��1�QQ/�.�"*=���1K(D�P�C���Z!�0u�\s�&D���0�'������2<܄���0D�T�%f1R�j@t䖡?���;��,D� ��& |z0kp�P-S-!��+D���RjD.l!�C=fz�$�6�)D�ds#���%�BP�3e�F���cI)D��p&k�t
B��0S����1D�0�6C�4���nV�r�[�o+D�� �@z� G%Q��X�JɖE�HAB$"O�L�����p�8�2d�S�/v��v*O��X��C�jvt6��K
*y�'6X8���$�[��b��j�'B�$	s@ 1�H��TI��X�1�'�T��m��E�ء��iH�p�JT��'�n��p�O\�XY稄9�޼(	�'#n@�P���Kovmb�͛�C��'wPe'퉵�@���啻YHhH�';�;`ǅ�3L�1�bN�i�� i�'6蛧�¾Om�P7�B�iK����'�:����ƕGf�X�`%�XC�'W|-Ic��+���+�a�Vt��'@�`�g¹lK��%�ȴ]g$�(�':d�*��? �nu)���QJM	�'��09�Ә�J�id�ɓDO�<Y	�'~�`"�n� ����ͩ49���'f�x�#i�"��1��0�8I
�'����F��	&��)��9*["!��'�҅��H[f~x|[���W����'���㗳e����HB:���'�����ؔH�zi!ri� :ܒl(�'��tˢD�=TUz�Ж׽f�R1�'���P��b�PiҫCHI��"sp-��\A�	 J��5i�L�<)3�U�4M<Ha3�ŝu
फ�F�<�s�K'���!�Θk����<	Í��B/2U�`S �us�ax�<�a��2-J�@��ߥO:�p�gmq�<�uc. ��
+B�w� �R&��s�<������9c�KX�w4��V��n�<����{�}qӬ
�mV5�cPm�<�"��O��A0���PU�N�n�<IV�~�&D�aG`j�jq�U�<!��@�6�X���R5%z<���GM�<�T$�r �Y�dǊ&�Z��
WH�<����'p��g�8zӞ�@2/��<�b�&rI�#�]<d��T85g�z�<��(԰6x�-B����]C>��b�t�<I���U������H�5�Z5���
i�<ɇg��>�|��$G7h�� �Jg�<Q �X�]���
���AJ@�J�<)Q흎u<|���+[��A�b��D�<�O�b�t���&3_�ר
~�<���f���3e�x���D-Bz�<�������M��!<ϔp�я�r�<��� �Mm���ŀL�]^�ᒁŕF�<I��َZ�>��f��yl�\F��A�<�����Q�
�3M�lh�P��}�<���R1)�����ʲ2�DecG��z�<�J����L:7M��j[4D]m�<AVf�Y�  S2�٫!Rpu3�M�Q�<��_�	��i@���*-�ڕ���N�<Y!�-a�4	X�-%�ezCh^�<�ծ�@��,�V�C�\���"��z�<�7�և1D���DR52�B|��́y�<�J�0X ��	B�
�I���&O�<�5%Ã�
������jc"��I�<�P�� !xX�R1�E2Ew�H���F�<�拓.�KW�_�N��=�6E�~�<������pls' (Z�{�<9���0(�Zhy��}�d`q��Qy�<�0�$��X 댅̂���^�<�rDU�J-��b�B6w1�����Z�<� ���U��2DM�P�O��Tӄ"O�\���&��5b ��$�|���"O�ȈҮ��r�ڵ�s�/S��Z�"O����ׁ@� i��\�U��k�"O���D�k�����
u� ��1"O��Y3�?՘xz�FOO�i3"O	��͖�����⏦eMc"O:PSaȇ~Avx�#g�����$"O^%봎�eN�XJ��#X����"OƤ6蛜єT2��֔opab"OF�X^e�|Qb%m�Y����J�<y�Ņ�o����A��0g~U���XR�<���:u�ȁڃ#�n,$�U�PC�<�!)Ɇ<���Ƈ?oN��cAMd�<�!�yu�E��NLn-����GJY�<,^�S:���oQ�`�
زJV�<�&�<O,���?hbXh0d�\�<96`��'3$�d�9_��I� t�<!�Һ.B��v��N��)S�f�<1�'?
�0#ScϷ\*d� ��Zi�<qad�$yG��3PH�7i�I�Òg�<i��OE������-x����`�<YBL/4j�k��Ŧ�"1Eh�<�� �!̡�h
#p��ٹ0�H�<�v��,d����ƆW�#|d�i+Z�<�t*�6]f�j�lJ��J�A�bq�<�D�2w��q��MĶ] Y��n�<i ��;(6��(�
�0>O�1�nU�<�� s������V���h�P�<��+@�2;��c$���5��T��`�J�<��$зEJ� ��~�ڳH[�<�T<(�X��� �%�X`��V�<a#�R	U���-.��Y��*j�<2_7>�u�D��������g�<)ԍ�3u���*�0ْ/Na�<�WA�o���z�ȯ0��jT��`�<�S+�&+�.�`�kR��`�gjU`�<	vÔ�@lЦ�D�BӪ���D�<� �����,�����e�G�<ycˌ�w�:\I�gGy�
��&��C�<���ȵ~�EyU��f#m˔+�y�<��&��f��Y@G,]�}��mr�|�<ǎF�y�������#j�!Kv�<1�Uf������Z��@Hn�<�m��=����b�ý3�*�:3ɖk�<��5k~
�P�+��2f���G� M�<�`j��v���zR�	�Z�*��Q_�<�%'Laͤ}e���=�x8�w�W�<	Wo��i��)ZG�/rGfeQ�W�<'I1q�+��G�������B��*k�-b�eO�br-��#��B�	�2MH�q�]'D�{D+�)y�C�I�8�QK'�37�Υ"7���g�lC��
6�5��ņ$�	��g�$2}.C�?W0x��d1TczE��L&$�JB䉟~&H8�@�*<0׆�3�(B�I�4[^���ٌ4�H˶c[ZC�	>:�:m@�/ /5�@��ђI�NC�I�Yf�VN��aT�� ��	2C�2��ԢP�
�̒�a˖-��C�	+1|0�w�G�ِ,�F��D~^B�I�|!�e9E*I*H9�y��F�Q�B�ɗs?D�y%B
4Z���qqo�/r&B�I�r2���	��,gb�!�Ȗ�^��C�)� TA)��pw���Y	q��TCp"OF5B�P�G���pH �	�����"O��cri�E�YbEH
����"O��3��*1���j�gR�O\H��G"O��1�E�t��#b&�2?�:"O�X:�gK�	2,�d��B���	T"O� �iR)q�b����?s�1i"Oz,QF�T�8�q���U�Ҭy"OTqSƄN����AVi�X�p"S"O���b�N>4P�fZj����"O<�I��I0�����c��[U"O�D; �]KZ��#ׂ=��z$"OF�i&�H�B������3Ӣ��w*Ol�D�E�^�Ҵ@&�K,i�2���'}�`8��^>Mhr�$d�ںx�'�VU�p�F�'ﬤK��
@�'�9'%� ���s���P�xr�'��#��T<�X�7Eڂ<�����'�~�����a#�q$�F;h��9	�'�Qq�X�kl����kZ6n4ɲ�'�rā�gp�\�
Ef�2PA�'`�}T�"��0���c�\}��'�eL�>*2�y­Жp��99�'91T�YР�������P�'�����U����zEA+NxU1�'q�A��HT8R� Ԇ�>�>���'����6�l��E<2x��q�'��x#�lX��(,!�=1�☃�' YA�a���4k$�!P��
�'��{w�ڝq\(I�����޴[	�'����$G?8<�*�� h�(�'�v� �%R��q�G������'
�U��Ɋ�T���"C<4�
�')�p�o�
Wc�J!$�fB�"	�'~`q1i��E�,m����W#��H�'��tx��AH�0%p��&H����'����`
�<RMp�l�A��ؓ�'!P��M�/FZEZ5iô$�����'��Z�
�������nD�S�'��uXQ]R�ĝ�$�ϵg�D��'\A�s��*�H�cbIV�F]��'%��IVg^ ����u$O�Ĕ��'�xT��� 2ȥ:�@H!;�'�ژ�%Ɵ�$����+Bn��	�'���u�˶-��(���V!<炤��'JZ�  ���   3  Z  �  :   �+  �7  �B  ]M  �W  �a  �k  �x  n�  Ƈ  -�  ��  ʚ  �  N�  ��  γ  �  R�  ��  ��  �  X�  ��  �  �  ��  F�  � � � V  �( 70 z6 �< CB  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)d�C��0S4���T:
b�lڍ�xb�۾b�24��d�\1F^���=���DR
X��£��c�N ���;h�!�D�\OXe��GW �t��V+ۖi�'�ўb?5IP`,P^6��uf �>�b6D�䩆�'cC�|xv�=3��YY��4D�P�uk0P3�M�4(�[�Mv2D�P%�	���;S�"u�pR�L.D�бU��\R\��-�.OЈ�a�*��3�S�b'�i+���({u�\r�c$���?�sΉl��k� Nr���/VQ�<!C��29�,aˇat�@��̑P�<"$�?(�$�pU�C���{̖C�<�4z� y �O�!	����LE�'va�4`�>#�����))w2x���I�y2�Oa��ك���A,]�/V��y�� =-|bu$۰&V-8S-�*�y�n֠0�J�+���7��q�gD���ON"~
�΄���T�D7^Ĥ���M�x��'o�s�bŃ=���w�˴/��;�O��=E���;'���&�l|6y�����?��'9NL�u�T�6*������~���'S�	S"L{a��T₋|o$�s��M;�ҭ/6�x��bہG	��{(��yRʒ u�͡#Ǝ�3��C����'zў��P��#ЯE�z@r���@�>�Ba"O��:��g~m[DE-k�\�RRaȦ����~�8O���y��eR�4�|��c��6M����Ox���IN�b�ʄ��H�@A��I��<�'Ta}bLR2�:2�W>!4��00�D��O�"=ɛπ Z]X��
֙��"� C��0*��iM��Q"+yȤÔ�%,���B�G��?�s��W�Oz�E�t�F�"(ŪRa�1
�V��
�'KHq�ؓ0�
T��`�z7��'"���)�'wN����	�7� ���Hi����*�� ��!�3U��XXҫ��2c �lZ@}Ҷi�2���O���,�C� ��%`�,UN "U�'D �1������8�CU�%lZB(<�g���b%oE;6�b�xW�r�`� /8�|��h1���3��)�@I0H��ȓB�� ���j=$�ES�<�*�S�D�<E���N�X��T�
y����&!�0ȇȓK]��q��U_P
t�F�@+�܅��>L�#�S<7Jr�q �_ Y�����Q�#�8Hh@!���?EB���#\,H	C��V��p��o��m��T#D�ᦆ��
*34��!O:�p��TFj�g �}���'"�m�\(<AqI��h[�d�)}{�:� $!Td���H��2��Č,+n�c� �e���K4���nX!򤇰"hZ λ,����d�J�	Yay���)q��a�FV�y�
�!�[��B�I�BQ��Dg�8}���D�(`B�I�e
�h
S�K�Gd��?�]p�'�n��@YO�p#c�m`q9���hO?yM]+8h(�d��vq\(��q�<Y�U�B�!���Ve�rK�<a���')ўl��i�]&��zh�P�P�P��2�O�扞NL��@�c\�p#bt��h�!��B�	0C�l0� ��`s�D��g�N��	P�'5�i�-mM)v��-;n���,_�~�!��T.i�2!�&mē�Ys+��m�1O�A��-O�b>��qk�?O�J-c���(#V�{uO9LOʓ�?��CʼT��e+T�=:�k�L�U���?��)��J�@���� �
�q�D+�CS	�hO��	N�Oi�������X�陳�lT�$�"}"�>�Óy����$���¼k4�@:� \�?yI�\$��'�ĝ�G�q��r���Z:���'�b)��N�4*��F	�j9����'��5s��_+]N�rւ�$W�~�(��d)�'m��Ր�BU5G���S@0_Jqʉ�D��(O��$tT��r�H!���v�U�:��˓�y���/P
�Pץ���+�jQb2~6�>��k}��L�<��hP� ܉��ʌe($#!����)����<�O��-'��Rp؛8�:B���{ �"��-D�X·Bm^b}��/� 3Y�Չ��.D�ġ��_�F�Z�!�u@h��d$(D�@0��ܬV��bu���.-�	*&O)}�d$�S�'�l0y��[u�:��i�F6��	Ʀ}�'�}�pc�<YO��E*_P:�I�}Ҩ3LO>r"�B�WFZe��%��It����IP�����'�4h�jڝ���y�� �/�&i�
�'����{͘Yr��Q�x2��@Ǔat�5C�}�)�7M���.̲^Ϻ�!��Q��y�(DfL�G!�FT��mۈ��$'�OJ�!��	b����HP'�J�X6�i�ў"~n��c2���7���9�4ِ�10��B�I%UԵ� �V�3��P#d�cAzB�ɨ%T^P�f�ؠe�vXJr"M-Ox��D�Ry�MYsrAYg��T�D�W��yBʚ*M��;�ΐ}Z�l���Y��hO���![o�8�S�5����DJ���!�\�Rp��#�wr����(-��Ɏ�HO�>11�!��<��e��g˞���/D�� ���5NWM.<B c �IL8Y�a�|b�)�S�t��2�/¢������T�F�X�IU8����p��cIB}�&E�$�Q�Qy���?�ӓ?����7I�#ǂ�z�*�
X�A��	y�V�!!ӣØo�Fy��X�6�@��>)�%�0;Y��0A"ަ	H��>��yR���4O�1y��\�-������ �� W�	Xx���j��@�h"H]��P��g2D���ҋݦ'�p ��Ȟ�(L��/D��95��+0Ď�P7H�Qx&ex�a'D�VB!6澡Ф&ėl:������<ɋ�ćDe�E���ֈ:����bqOF�X���0}"�A�^J2�`j����2'��O��=��Kb�(��$.� � �ղ9
!�$�$x�!p��]"��I�$�
�iJ��"~�@�#zV-��C����	�̡��'�~e��(�0h3��{evh0�/?I��i�ў��OX�"f�����d(<N�y���'�'�R�0�b0w&4���F�{�����'��:cC�~"�Rd++�0�����'�&��4S�A��}?�����@�
�!�䐕>B�H0��Z02�)c�ϩ'�铲�'1�|� ��gOLͻ�J��H���Vd�|�<	�'ϿG($iF�m�ɠT�Lv�I~���O|D�p!�A�4�R�C�e��#�'n�+P��2ݚ�+L�	����'b4R��7}(���D�n�7"O�"#�X�-f2;�$E2�@H�R"O5cWRS�|�F�Z��ɂt"OޠDA��	�Pj�kF&6��9`"O�yi���=�vQء�Z� 58U"Or<#B�R�/la�BL�Q���"O2�z l��6P�%�m�!V�y�����L��X˖�ȧB�ؤ�D�
4s�"@�B�3D�H��σ�O�>ea��/*��D'D��[Eꚗ;����c+K�s�鉴a&\O<b��!.ܲB�0��a$ďj��
$1D���BL�]%�4j��"D!�ة�.D������L��I%�ҝQ"+D�����G("
��Ҧ Ԃ2*��ic�-D�SR��0�\�KV�F�>8��).D��8���rN��+6�E�.j`�9d/1D�pq�@A�*�)�g}7��j
#D�3� �$����q�I�z,@�.?D��`t��^۶���C�y�4���%2D��� ���Gg�I��N��d1���/D�t��jM�vb"%����?]�Q:a-D�(r�� 9`ev+���/�ԉz�6D�d��fD&c�X]�w�]6���y6�8D�h��Ɩ{(\8�G�*B�.���k7D�tyF�Ŧ��0-?0��6D�H��'�8Cr]�jP�OVe��h9D�DX4��~\j�C�?o��@�5D���&�J��Q� P�0�X�X��'D���@L�DȞ W��_�p�6�'D�x�"�<�8�ŭ�0p�U��+D��j��ӐXX[�N��ѓ'I*D�@	Q�W\LZ��r�[1E�L(D�Ԓ�D�<#x�zϛ����a�-!D��s��/.��$1�BL;��#�"D�<���Էk�����!ZK�tR��!D��Q&.�v��ܨf�.`���A>D��*��9<]qe��=ƍ�P�<D��a���/�X�c!�$/�tA��8D�� �;t��	E�bx2�$��X��Y�"O<q`��qX���s�ҘTxѕ"O�q���[M���S��()���c�"O^��ӝ\´XQcGQ�T�s"O2e)���U�R���E�V2 �:��'.2�'Rb�'���'���'��'�=���)<��{�� 	Kl0���'���'|��'���'R�'"��'�b���\��B�;�F����'b�'2�'�'5"�'���'=baH K��^.X�4G]�1}�h��'���'��'��'`�'ib�'��`��A�n^��C���B��l4��'l��'"b�'�b�'4��'��ǟ�rH�8��K>n�x�KVa�r�'��'���'.��'��'���^�i~�T��+BG���q �9��'���'���'D�'9R�'�ҁS��Qh�#��p���I���'c�'���'t��'Z��'Y��� ȆQ�p/M��]bU���'?R�'r�'2�'iR�'��A�M���
�ǚL��%Hu�ٛz{R�'{2�'�"�'��'E2�'���h���U�ܐsOJ����T&a���'[�'WB�'��'���'��[-}$L�&KȻw��fC6&�"�'�B�'i��'gB�'�b�'��f޳`��`���=�t�ICCV��yR�'Sb�'1��'�ZΛ&dg�����O��;.J�I,�4eC1g&�M²"�yb�'��)�3?A��i�}j�b޷U�D�Pb�l�@�9�Mب����Ԧ	�?�g?޴w�`�7)�
�^0 V�mjlDx�i�Bhɑ"�������cf���1�~�&�N1͎`���L694��j$!j̓�?a,OR�}�L�E|.���0&� �����f훦�Ϫߘ'��6�mz�7k��[.�*��B��<8��w��i���<%?E�3���%̓	�ĀqG
�X���y�Tp���̓w� 7+��%�,�	��4�$�d�8>p�1�N#Z0�rP�*��$�<�H>q��iE!҈y��Č/�\;��� (�Iհ��O���'�ºi��$�>92�IkԼ����؍.��D�3�Yp~���*4c��?��O�&,�����I��tp$� X����g���'e�Iß"~Γ_6���O3 ���;��(څΓ7S���0���Ŧ��?�'2&,PjA)�s0493�mQvR0����?�ٴ�?q�-I%�M+�O�x�"'����(A	��nz$8�Lɜ>������-��O��S�g�d�I��K	FN ���D�f�	�'ۛUj�nʓ�?I����@�L�֥h2O�D_��&m����O&yn��M���x�����Y`�B���9����h�g�� rI[���ɦmk�y#qF:R���3	O9�"ѫe`U-s���5��  5F8�����a�J(i��N���`��5L���*��l��tx�I�,m��� ���UޚȨ5�A�-��!��Q]zl�d�DD	� ��\�sg�y'£D`�T��EZ⽺W盒C{*4J��N�ڔ��f��Mg�i6�U�D�n,�P��MJ���a�pt%�mŵ�Ұz�e�Os����X�p����ӯ �q2Ytf�Dw��qP�M�0v�`��F&.��0uo9��A�hGF4B��\d��倢��&R�$Q��<Fʝ2{Ӕ0�vn������?�bg����?)N>A(O\�:�W����3Վ��5��!�R=��į>���?����$K�`��'>����r�h7��]_hh���M����䓴�ē$C�OD�W"�3K�)
���+[�� �i�B�'��INDx-0I|����V���8���(��+n��y�f��2��'�副Z"<�O�htJ�͓} ��Ӥ��%�*���4��d	&�f m���i�O��i�R~�'�8 ��K�<LC��2O���M/OD�(��)���z�,\QkG4,��1������7�XD��lZ�l�I�P�Ө�ē�?�dA�I���1#�`��<���Q4/��C�H������T�l�L�)�Ƃ�>r&�st!S�� oݟ\���TAs�����'�2�OT(ذ�B!N4)�$n�9j޵���j�1O���O�D�2���@1̱cC�-|n�S�u�����2b���>���?y+Ok�^AF����jB�>����߳v����!#^c�t�������wy�l�,GZ��{�.�9�A-Q�,�$))���OX�D6��<��������C�|9�g�qV�<���?����D����'4��̡�J�8]|x�#D�Pl�''��'�'&�	)s��jbt�2�� �M�`,K�@t�'�"�'
R�`�D����'�NI�W`��e���_5h$�A��ix��|S���N0��q�j4bňE<0	*L)�˃��7��O���<їf�6�O�b�O�jxiŀE�jE8��±���c-��<�ψv������Dxʑ�� <���B�
ǖX���Q��P ��Mw[?����?�{�O�\ñ�� y�L3�'�h4+��i9��\�&"<�~�eH* �ؗB�L��,Pn����[�B�'���'��T]�0�	��I5��xO����2p�ĝ�����MKtȷ������Y<Z�F�F�9>L�S�|��%`���$�OF���K����?9��?��'��%�A�&����8
?2|��}�g��;Z�'Lr�'� '� �I�����E��l��������ir��R!�	ԟP���$�֘;fX�mUf�$��l� �t�mʼXN>A��?i����*L`�Ti��?�� �f��O�����<Q���?������?��{	^<���;vv�\3ЮW=SP��y���(�?�,O,���O����<���Q���k3��x2��,pZ���P	:�M���?�����?���xp�r�'�^�+R��/����VZ�~� �8�Ot���OP���<� ����)�O�	��=(�Ȫ��7rS�p� ��e�I^���`�	��&��=�p �;Bn�R0�[0A��i1���e��ܟt�'h��K Z>e������S ;[>��t���gK�1ѶC�(=�J�'�4���4���͟|$��J�<��w��3c���9���1�b-o�Gy���22���'�'��_���33��%�ƽk���k�N�mQ�7M�O&��Q1���b?�����Da�D)ȇ.���j��g���`�A�O�D�O�����˓�?���0m����/4^R�XRB�R���im�Ȑ�������/����p�`�){���M[���?��+0l��(Op���O����H�ԃ�F��m�S�J	_zZ]p0� �I��|X%��	蟬�	j{�+�.K���bR����4�?9��>����O����O��Ok�>�уuE6_䲣�Q�\X�ɴ)��&��������]y�B_ $T6+4R�朄8'� ���J '�Iڟ���$�����()��*O���c�Q�i�.����'|�%� ��џ��hy�
��m{�ɀ�$c��p�D<9�Fucd԰'!���'J2�'��'K"�'Q�p���O��C ө���0�������S���ß��	Wy�Bu�`���(òr�,V�0y2�W�,o֟P�Ify��'Y��L��.��ɋ�XLNy�Y/r"��i���'��I&~�t�L|������\��,�Jڢjz��!7�ݽW^��nZPy"�'���'l�����5fg� f/�%�r���"QB��MF��M(Op���"A��������	�'�Fl��w�\�%I"B��9�۴�?����?9��v�Sny�X>7��G���pKX?��UQ�V�H<����h7��OV���O����m�i>5�V���L��&$� ]���BӬ�*�M����?y���?A-Oz�g~��D)��k��ܻZZ��J�sB6��Oz���O*���NB�i>Q�	�t����=+T.���AE
4"��g
�M���?A)O�x��y��'Y�'��D0a�Y\^l7-J?��ŀ��d�*�L0�vH%��Sȟ��	yae�,+�A�23������"9.$6��<�������Or�d�O�˓�n`�I 	��4+��f��c���4��'�b�'k2Q�$��Mz���[�8�X�)�-wn�r� �O|�$&���O2��<���� <��ʦN���߹WS�(P�A�j�Iȟ��	���' ��'��q���'6�$3"퀿z�f�w��7�����K�>q���?����dR�v�^�$>E;p�0�0�J�.]�`���j����Ms��?�,Oj���O�p���O˧`�}0Z<j���R���8Y��Ȉ�iT�_���I�|��Op��'��\c��4�Ҋ��)c���� �&dL�)J<Y��?���H y����<�O���3��&��ؒ)Kr��4��DI-8W$�l��	�O��I�L~�١`<�I�d����b���]��M3���?���*�?�֗�D�O��s�Ҹ��͓�@�°)��[�bK�����iͰ�A�'���'|��O��)��6�jtP5iJ)��$��P�֌�>Uذ�y���O�����U���4�^}����,�����џ����{�eIM<ͧ�?���~�i�P��{�4����P@}4hc�i8r�'��µ4C��g~��'tB�!`����G�x�*ɐUE,�&7m�O�0��O�e�i>	�	؟P�'a�kՋ��J}�XR6$�r �[u���'`�|��'{�'"��'z�I0Ub�M�/�nq{C(�Dj^����W��ē�?����?�-O����O�U
c��*h�B���\~�NT�׈{��D1���O��d�<Ѳ� 
?��t�� ��*Y��Q�j��n8��ǟ��	ҟp�'"�'�X%b�'Ð! �-E�8<(۳aO)	`UPB�"�$�O`���<)oD�yx�O�R�ڥ@]> <��:	�9 �,y�lbӖ���O ˓�?Q��PG��������; �ᛰM��.�b��B
��f>27M�O���<rǀ�}��O����5�-n�蛖$E�#�~4CC��6�M�.O����O������O������ƌ���`V�9��"'&��Y���g�i��&F� ���4b���̟������$��T�R�أ�/y_�y(�dN;����'z�-J2"1�	����禡&MՃx�,��a�y9����s�^1�oL妑�	Ο����?-�L<���B� �|!Q�A���pW��ٚ�@�d��������?�O���BJ���\�~�*��S��;8���۴�?9��?��H���?i�O�����YA�"�G��W�"is���v�3e<<�6���O.���"G"i!I�' ���a�X2yS�7-�OL"〲<I�_?��?1)�j�f|s&h͕k�t�� n�="��I�J��`Sl9�I՟��'E� �E���svפ��!���Y?*��(4_����ޟ��?���?�D
��#��0��ۯG��v�P�_������\̓�?�/O�d(?�|�3� �i3���i8��Z��Ư?7�xڇ�i��B��?Y�79��#p%Fɦ��(�z�t���h��.`< KT �>����?i������@'>1�e膚U�*ݒ�7\���ɰ��=�M[���?�.O��D�OD(#VM�O��O���S��3����ϫ}\,���4�?a���dK�-�$'>����?��!
x���@̽0�DaR	�*]��7-�<����?a#'��?�N~J����lM�y��a�S�TЈ4�V릩��֟�h�U��M;���?�����'�?��^<l����a��C�֬��"��I͟x3+L��4�����O��x�0�IY?e��@�&��c�t�oZ�I�(=��4�?���?)������?��"���!��1h�\aSL�O<�c��iF���]�x����O��O��B�G�}�ɳ%2�ݚ@f�̦��	�$�I*�Ԍ��4�?���?A���?�;w¡��%\�%C^A9�+�(���>��f�\��?����?�̳�A�q��0J�P��ş3ǛV�'s�p�)iӨ��O�D�O%�O��dB-��x�p��a��iA�����'�%��'@�	؟��	���	ɟP3��7n�v|`z�3�"P)[�B��Eى�MC��?y���?��]?��'����h���H�f�����AA�?��a�O��d�O��D�O����O|Tb����� Q+w,�:��K�)�L#p����M����?����?y����O��9�3������tI�d�
�P�b�H���d�O����O��d�Ol4��XǦ��I���QiL�d�c@dW�2G�1�G���M����?!�����O����9�v�'uD)ZtgP7h�A+��Z`Ԉ�۴�?9��?9��_� ���iD��'��O�)�3�`K(�dI�4e����r�����<��b@�'�?�,O�i�bI�v��	!�B���E�Լjܴ�?9�+^iH��i���'/��Oq���'����".��%,HdI��ŏ\ ���?�hL-�?���4���O�޼+#�X��dr@��	����4y��$se�i��'wb�OV���'f��'��TK�f�5�Xur�O)]@-�@mӊ@ʷC�O���<�'�䧖?�2�&x��8��f]�X��̃5��(�6�'���'�xi��oeӄ���O`���O����\�ǅ״� gg�A� �є�i��P��" bb��'�?���?�ǅ٭5�`5OV�zH8Р����'��T��`i���O��$�O:,�O�5.���m̈́d]�!jo��`��		'�t����IٟT���������i��؃_N��zC����A���n�����4�?���?���s��SYyb�'-�U�$MS1G�Va�	Ǹl�,ec����y��'�r�'�b�'�哦,�a޴i�|�C4�/8�L���O˔A��%R�i~��';2�'AX�����a6�sӮ$(�?-��b5oH�A�6J#W��I��X�	ڟ���]�r��4�?��'h�I�6�Y=R2`!X��ڤ+�:)s��i�B�'J�Z����oX<�S�<�4��Ԑ���_��&��!B@]n�ɟ���ß��I/�m�ٴ�?9���?���15��(�~���t�Q�'f�e�i"P�8��%@w��A�i>7��3_�D%+��/]PS�N�=6���'��@X�dW�7��On���O�����Z�$�:2&�x)�%.�0��W���&,=�'�/�3r�'��i>��Lj"��)g�W�T��M�R�i�|q�A�wӞ�$�O��������O��$�Oꅐ��ݼ2�\آ���M2WF�ߦ�iF$�˟d��ay�O/�O�j^�rR�j�.P�\`B�\�Os�7m�O����O��!iQ��	�IşP�I͟l�i�q��Ѱ7{�Ax3MB/��e�&wӞ�D�<��`�<�O�2�'F����� 1�X�2�"<�S�a�6��O�@Q��D}bQ�x��\yr�5�k3�ۡ$ }�bp{�� 8����� ��d�O����O����O��'I4���(ś/F����$�(�8��p�M*����'���'~�ñ~�+O��d�&A5������;u�A�BD�%��<@0O˓�?��?q,O<�r���|*0-G������o�xsP�1e�<���?�H>����?i�d_�<��IO�BT����?S�yB&'�[���������'��4�t	*�	S#:J� P�UF����?F�
m����'�������#m�ȟ �O��8� +H4�ŪVm�d���U�i�2�'�� \<`H|Z������x��9��.=ʞ-9��,��'%b�'����'�ɧ��F%>��X8��^�e�܈q�}ޛ�W�ȳ�.�8�M��]?���?i��O�,���^�VjRA	��349���гi���'�!���)�}��ɜ�� Y����vA��HQx7-�O���O��)�o�Iß�����X�z�Ԫm�N��P P��M�#����?IM>E���'1|x�C-h��� د\P�42A�l�d��O��4(8�%�<�I�4�Lɘ��%Ϋt�`z���6Ԓ�n�s�= �>-�M|��?���f���Ba�]�B~�2���L�"�i+rj�6]^�OR���O��Ok4u��]��gZ-jߐuJ0�M>A����KC�c���I֟�	Byb���,�b"n^�;t�i8F��j�h�"���O��$*���O��� �� b'f(>�`ݓ��ǁ7������O��?	��?I,O��P�.�|�#�Q�8<�!�"/�E�Q��LNZ}"�'Pb�|2�'Q��W��y�(�F�nPZ�OQ�i�M�$`��4I���?I��?A*OjtZԍ
`��Y.1���m�0x�gSHܱ�ڴ�?!I>i��?i(���?QK�l�dŚ>���T��
����(s�����Oh�!�ZP�U��D�'��d�:� ���4t����,
�6,5���x��'l���O��<Z� Y��@�A�LȘr(D?.8
6��<��X�&"���~Z������fȆ*U����	�&S
�E���}���O���>OޒO�� Hfl^>��96�ǙQĘ��i�Tx#t���D�O$����Ԍ&��S?c��]�f��c�XT�'�FQ�y3�O���<�f�����ƋIz�E�����1p�G�M+��?���Ũ�x�Oq�a�*X��%�$l~�2���s�8�l�Qy�[��0I|R��?!�
����׵/�8��o (��۴�i�2��>58�O�I(�Yk����(��|(2�p@Ձ	\�lUy��'��	ş��	ן���˟DSQ�Yp*-Aѥͯm\5D���m��ҟ�������B�����V��aə5M��9�O	/F�$n�B����?����?y.Ol��đ�|�uH�E�����fǕ` ��BA�]}��'[��'��O,YٲW?m�d� �.�BAf�_���"bk�>����?����?��P��0+�d��
�0������RG[�-��OR� *Xm��&���IAy����� �n%��L�=`�LK��0U�N�l������ɟx���}�.ՖO"��'��t*�y '��@��� �կJ�
O$�d�<� +�G��u�h֖-��`�K�"L��0	��R�M�*O$1������Iӟ����?��Ok���@���ȲS�(�xՇʰ#��'���k�$%'��a�@&M}��WL$�`ܴaAFX����?���?9����Į|2b�O�*s0=J�޳8�ԽC�eNR��-
`"<�|���s,���dA���h�HϠJ|�I�b�ib�'�gnG�H��'W��K;L��X��ٟҞ��2)���BIDx��#�I�O.���O2E'�M-mz��16&6u��L�u#�Ŧ���5{%���N<�'�?I����	�
d��Pc�Ox�A)�\�!��� ���<)���?���?��p6D�C@fɝ	6.��w��>�
����<��$�O����O�O��侟���l��n,�[4��[�T5��j�n�$��t�	۟P�IKy�(XƮ擠,RzՉD�]�|ؘ�f��;m���?�����?���NP�'p*�;�$]>'� $0B�8�@4گOr���O����<�&��pE�O����06��3��!z��	�|Ӱ��$��O��$��NK�O��Hw� 4e��q�Ϭb`��9��i���'���**3@�I|2����wÐ�d0�UjGeۈ.v9��eC#މ'\�'����T?E�r��oi���V�}�V�{�{�˓<jB�c��iE��'�?��'Z+�	3U�����l�mq��B�N�?��7��O��F)i�b?���m�8'�4Y�B�/6B�g�j�n�y �N榙��͟T���?=�L<��M�@H{ ��7b�.e���=TH@��i��dGy��	�O����@ز��l:%�=^)���tL�榕�IӟP�I�}���L<���?�'m �����U@ts�D��7��i�}Ҫ���'���'^�Ǝ���u��2a֤e�R�߅A�n7��O��0��Et���(��O�i� &E�N���eO�Y��+�*�>���e��?���?�*O�xj�a����I�.�Ȩs*[ ?��$���	��'���I�S6G�%Y�]�gA�Oe�4�,šShpc��I������p�I2{%N��~򐉱c�$;�$���NS�@n�@��ܟ�$�D��\y�덀�McF�V�����3)E89Q�I���_}R�'B�'��I�|�:�����V�&+"k� c�:0�R*��<dN�m��@�	G���?i�{��A�~L�92��߀Y��̪��Mk���?��?	U���?y���?����*�/�08�"0�TI°!��zv�Ǘ��'B�\�<��n6�Ӻ���ߪ#�(
a���j���2EH�ئ��'gN�0�wӈ��O���O	x�� ��S�U�@�����$f��nZ@yB��$`5�O�x�)P(kV��H����~�xQ�VI��Ms�AT��?a���?��������QּL �C�x�e;b!��X����EV��;T�$�S�'�?�C��)}�U��n�X|p G:U���'Zb�'�pu2��*�$�O�������6�O�t6�%��(����'�	P��c�t��՟l���?M<Dd-Ɠ&t��
ш%5�T��ٴ�?-�>$"�'�"�'Xɧ5�(M�:`2q�d�(��Ѓ�l���ĕP1O���O ���O4����bJ��brn Vٞ2��L'�X AD�<Y*O��D.���O��I��<�n� N�s���>��7͌-x��	�(�I՟��'���Sc>iV K�~�B<" Z�v�8�2'�{��d�O�$�O㟈��b?1S�Q�l������j��P�v}��'r�'���'�:��'U��'������4=HP��әd�H�p�w�r��%�$�Op�i`0�$��)��%(yL��EЃj�jx���x�N���O
���O��"�O���O:������F�PQx�K�DA� ��1�O�F��З'%yq����rgS����`�HIN��pZ��i��ɵ�����4/(�SǟL�S�����w�����-r���d$�'��E#�4��'�h��F �g�H]�3gK�aϘpXش�]`��?!���?��'���|�� 2��N&P�p8t,�$/�հ�_�|�p,>�S�'�?	�(�1*����L),ƪ���#I\�V�'��'�H�:$>�$�O����h���#w�m�Ռ.
����";���Jrc�4����`�	4c�ɑ��9&� �����+*��s�4�?YM��Np�'t��'�ɧ5 ��r@�h9�/Z8�U[I�Py���'�R�'^B]���sAV�[c��H.��A�d�����xe�M<����?IL>���?ْ�Ŧ7�"X�1b��iQ8��1�
�D��<���?������,��ϧ+#"�V�^�,�H�X6a���'Zr�'��'[b�'l4�O�̀b(״��bJ�li�Y��T����џ��'Q"�+<]��'x�V/1V$x@Q��T>�k��P.'A�6�'8�'O"P�[�"��\�<����:�8��n�����'�BS�Hc��W���'�?���T�~4j�'��QNQ'��&g֘XXp�x"�'��z���$�*)�ו3��|�e�-�M;.On����E�)b����d矪��'��k�\�έ���Z.P���[�4�?��tF1��JP=|Q2f�"v���l�,HqNm�ش�?���?���Q�'��A�U�H��ߨ]2�)�g�OaQT6�#"��"|b�n$ ;E�I!`�� �l�%?�q�ǰi��'�"�	O��d�O.���/WJ�2�nE�A�p�b���%]�c���s�7��-c�PX� �؛B�Z���(՟,t	I��>��m˰�,X�t=��Z
 �6J�T�?��@sG�;�8h���D��_y���&�� �����	a(���B�'&���9&&��[�<�e�3"��b��O�Y���<Az��#Z%@��t1q.��O�F���%]z��7�D-�j�XGW�,��+gN^# =�sn�	'��S��=o.��At!�1��) �	P�8�ޤk��D�ry�]� �S��e+�tD��c��E��ӁT�"�r$c�'!�����	�@��|f��woa�Ļ��O�Lk���8��u(D�AlD:��'^2<��?x�̈ ��X�Se�ߒco��$��-�� b�O�g�џ��æ�O�o��M[��@�
 ��-��S	Y�f%*p�,O��-���tg�(��T�4+D=��m��se�̄�����ǥy00�gS3D��1�Q�_~BP��������M�'�?������B��?�V
X�?�B��g�'d	ę�rgݾ�?���T!h�e����2�,T�8�*���'w� �� ��i�@�$��~�R��OrP g��.f��%��T8P��Җ� H��O�L�I�	V�X��X��Ŝ?ZP��M���^�?A���h���$���d˔�65��p0��F�G�!�Đ#J�,�0扞����Y�DG5S�ax��:�?���A�"]�)r�AJ3xð���?����?����%=ؐS��?q���?ͻP�.@�%&�	�Ƈ���j�� ��3{�H ņ7/�
u���#*}��A�B����=+T��qI�#%SЄ2B�8b\`�AO��8"��d���|%©�oV0-�l�'<�3��I�|�t�a���䃓l��Ofў����J��$��\&9�	�&o+D������4D&ə`d\�Y��(�-4?i��i>���Ly«�6V�q�Վ��-G�����`���i2�' 2�'2T�]ٟ��	�|�βe�|Lr ٥F�}2���0�@���.�<^ ���v�gF�=f���@�\�#@xQB�)�<JFz�A`����=�t��?;�쬁���Փ�	��&$"h�ɭ�Mói��]����U��7Ql�HB2$�VH[W�D�c��ȓoo�T���E�P6d[ѥZ}�-�<�'j��<�'��=)mt��������*�>u���K�۵C��7L�ܟ���0Ҫm�I̟Ļ\�L�B"��(q��@�$J�}����>|d�sBaX�J���Tc��8�����0͓����
�>*�@@B��\�Rl�5@�*C5ZH/sFT��֪��kmQ����F�O*���OP�K�;�R,X�c� 1.	3��L>^�ʓ�?y���	�%s���SqA5>5�Y&'!��ڦ!�a'�h3����o@dv�ő�-_�,�'~l�&gz��D�O�˧*dd�+��4h����Xo����m:� K��?Ń�0����3 -6������i�|*P�d�.�{�EȷG� ʃ�Us�$�
X���Pf�ͫ_`n%B��sS�M ��S5�T[��Xl℧O����'�2�'���I��+��9��تJ��MB  �?�1O���/<O���hY;z��[կY�@�,�0�'4$"=����t���`�D޲]�Vt;�'�6y9���'���'lHh�fS;���'����y7o�%O�����	j_T%�u�T�p�1Oҡc&�'�J�B�e�� K2 �4m�Z�N�#�{��F���<�U� �I����u���b����?��O��ɕ��?����?��
$h�����N��z���R�����xb���B�������b<B�K���Čp����<P�A�,��`H�\"�2=T�A�Z��e�BD�?����?)��.$��O8�du>%#����&��	�#!�,s`<�.B�X��,�	,T�{3�+W��x�Iz�? Α �,ܔ"���!�f��pȐ3��(s��O8�h�'O��V�<m��Ί�=��dQSo;�?�ŶiF�7�/�	��O�p)�G�;�=�D��m�\���'7fUy�g��e_BhУ@ؓX��u(�yR��>a+OZ`�G&�q�	؟�y�/��d�zX+�B
Xd}K�	�ȟ���YC�p�������E��ذ6�\�I�cQ0��p`�%�l<��A?i���d�*s\��Ј�4$�T�؃�kp��@��#i���$Ү��c��	mZџĳW�\����0�&�@b��)�B~y��'^�|����-\:3�V�pib@�(S5h�!���Ӧ�a�BĬ�
i#$ �x��d�޵�M3.O
Mza%�&4�����O&˧`�����0"؁R���gO�}#@׃W6�a��?��`�*3t����C %#c�i��k�T"��n4:I��- �� ������
K��y��E* [�2C��~�O�0sWl�=m�"�#:���YI�@pGB�O���O���>��m@��K	N�$���(��y�O�b1�On�����;y�Y��o�'R�k�� O"��'�b���O��#�����RR+�9t��tL�}B�'2)*}��-���'q�'��w�l3c�	6O�Q��o�<.Fb)#d"-/j�0"���q��"R)q1�bO�A��l�U�t[W�ЮRe�L�D*�<�T�A7�B�u�UR� Ü�q��ORdcg�N�d��LR-Z�s.A�7+���}2,OD�s�����Oc�Oh�F#�c�A���ڿC�Ш�"O�LR��U�z����那v��Y!$��؍�T}bZ�\�.�T������ޢ=踉��@�SA��I���$�	Ο�����u7�'��5�����s�a� �;ƖP8s(�g�v�0F��,6 	�E[X��CBˋ��^0�c� �Hn�AK�ҀZ�b��2�
)?�4����-��<I�e�}&$z�G_�S��D�f�J���I�I��p�	U����O�f|@$�I>�@ɢr��0��]S	�'}�91��8 ���k��3-۴eЏy�,�>!)O���"@J}"�'��8�W�Ѥ4@p�h1��WtQ��'�B���'���+h� n9>���7�|Q�����22jl#`��%J�a�o�,��r'H�J2�6�X��}�DU�JnT��*:(8��ı�p<!���x��Ry�aT�&�Ѣ+���I��!�4��'���'V�ࡳ�'w/8=a��� ��3�'�H7M٤i�rD#��H%TB���T�2b��<�W"�RP��'�W>�9���� �s�J�YHXh4��M<�X�4��mR����m��,T��d�A��\>aI�鞥[�vM�d�D�zC+)}h�1�6���\����~r�$����X��ѩ.2�8HS�
N�D��S!R`ӌim�̟�$?��S.8�5AD�P9zQ�Am�<r5>��<�����'n�'1��G�
������2;�Ó<ś�~��O,�B�A�h�0�� �I�l�:ō��1��ȟ���1o�1ic
���IܟX�	��ɠ��3f{ ��3�ۃ(B�%rS���?ʎ�ju!M�`�p��8���|&��+� )pT I{�(�>bf�k�.�A*��#/t��9�sʧ ���>�O�a#%FЋ$�P*d�57����,�O8�=hn��)��O|���O\i �k�`��8�e��M��%�74�ز0$�3,���Ta@$1.2�4�1?���)*(O�����P8-8�y�z("uʎ(?i0ezV��O\�d�O���S޺���?�O�:l����/�(��gʙ2�h��B@МY�V1�����U
l���+hџ�B�/�/D�:Ԁ�,�?�!�����2|L#I�� �Ӱ�V�m$��FB��9v[��Ȏ?�m0r��|_�����-ꛖ�{Ӏ⟼���ԀI~- �0VǄ?Y! �p���B�	��h(��g˓5���2�q�b�x��OV˓$��)� Z����
U��*V�7פ�:�GZ8%ئ��IԟDx���	�|R6l��q��@�e��N�a�'�>�lY�D�2�=ggY������+�xQ��AA��9'�*� �Z��l�����h��s	�M3�=���0�'��������xv��[�b�C�y"�'��y�����l��֤d*� V��xr@rӆ��l�(�j�IƤ\ b�by� 0O�˓k� ����i��'��S�iy8�ɓ|s��+H�U]����-�&fH�	���`c���'"���K��H:��|�,��<�SC5�X9��űk�0|"2�>I!͓Y����GD3�"~*�K�L#p���M��x��ax���}~��qӂ�nZ�(�ZB�Ev�R�fM#	�t��Z̓�?��{��P�L1	A�YP��?��8�HO�U�7�È/��  )�t���ѳLu}�'���)h%�Er'�'P�'��w�x���#�����'@�N],���2LNzʓ!�ܥ�3�Vk�g�$[��Y��-�`&
��*NP]��*��)��$�3�� ��L>� F�0N�(��qk`���J�BD"Ak���i
ݴ�?����&�?�}�'H���� �w��XL�S���d�}4��r���Z���◾j��ɀ�HO�˧��$�!Jl���3Υ�s�EivR��&S�%Ѧ�$�O��$�Oj᭻�?����$�K�L,~p���S"z�洉� G�4t�tiD�o����D�d�D��ͳN����g��@�`��-�(���ɇ:[�}Ad���AD�X�1�b�t���
�O��m���M�����O$��[ת==~���_�-�A�2D���Bۀh ���D�ʺC�j�.3�I���<aq�ҝ�F�'RB�&\�Hz�>,�D�YC�:R\2�'�PM���'9�3�(�f�۬�L8���eK��4�t�H�!��q�q��=�p<�R�a8{���(Z�ε�	�*�r�{6Ș�HD�U�Ǝ��� ��CvӪml�۟�zìW7� +��CRT\؅b�hyr�'��O>� U@�Su|��� �9�Nls�>��ڴ+e��KCɂ�iy� Ѱ�11bd�͓��$��Y����g�O��d�|�]�?Q����F����͂�6��<�WH���?i�#��{��������4`�S�l�wF����S�� }�k�+�O�j�b�N޺�:th1m�Qr<@5�>��bZ�(�Iȟ���F�'*\���K�6l�X�W |N=�<����<��K����0�-� a`�a�^����dF$g� ���Xv@�qnI�-�`@n�䟼�Iݟ<0�߅�Tu��ӟ ��ǟ��;6��2F�Ñ_-���M��1A�d`�E�V��`F��W��A���]̧`��[��9�I<j�����#00b|��iQ!�N|��*��ow,��@$BG�'��U<hia�T6�U1u,6 ?�s���?Y�Q�0`��S�gy��'E��Ҏ� LN�q���0\���j�O�d��<|�&]A�a\�2D��b#���A���?�'����E-LL���0�X�m����!14 �l���'��'B�e��I �	]�
�!���$YT�u�s�X�Z?t!��怈qw���qW���D��&�uR`n��b�vm`	�}4�Aa&V�,�D ϓ|5��;�朷|�(���#sH	٥B�� �I��Mc���D�O�������<9�NX0��0nd���եr��G{���T&}V�!G��-$�Xw`3�J�O��oڛ�M�)On�����������L
�FO�Z�8m ��6f��b����C� ���ȟ�'�Щ0�1
.����#@6�X7�@ ��i0t�N=i �	��݋B��li7�)j8�b�H�:�ĐSsfd���U�WF��*Mp�Hy�� lQ�Ҷ!�Ofoڻ��$�:3` �ZoB_M5��ۊol�$�O�D4�)§�ư¡��3T*6Q���48!����b;��%Ł^��	SlI�#�vDW� �zY�[���Dڴ�M���?�,��X����O�Y�BD�T(���ɞ��P���O�����\�&9z���).�Tp�����ʧ��� E��	�����3��!���	2�'ЍB����$0�Nܯ�H�n�Q2�&k`�	��G�v�4�>�HU��8����p�	n�'-��Ȱ''ެ:�L�c�eD�n��0�<1����<�4��dJBh���]�^�KU~�ܨ���Ѐw�r�@w��0���*$	l�ϟ��	�|�0��P���I��P��ßX��z�.-Z���+Mf�r �Æ>�8�J���DH�>o*r��|��B����]n�@8bdl� oLM�WeQ���"Cb���|�+�Q���f�����M��(cd]�ܴa��ɶZ����'sr�'�8m(PH�a�T�$��2�D��O��&%O�%z��*L`��Z�������?y�'J��#"eŉx�@�3��@��l�v�!�%���'[R�'�bEe���՟�ϧV����:)�a���.
vnԩs�0��P����O��ի��*O���p�(+���	R�V+$�w�D�YTI��ۋ;���j��̙O!ax��xL�hS��}�.��
$fp����?�O>���?ɏR@ ��r�e S�T�r-�)��yD�XHL����b�"�V���'6�7��O���Lq6�f��b�ٺ���gHl��a�D�a�ˁ�	�&�����V� $��Fi�E�2��)nk�h�sG�����ȓB�r(�6k��I�>��եŔY����?�틂�Ӹ1��Yi�H�dḱ��'�t.��{S�ȿSm��(�a<D���ǀVd�Hڤ�/(��|)g�:D���b��	��� 叟+��$c5�9D� aD`T1/s���N��ap�Spb;D�� �<���J<.� �Sg��8?F��b�"O�-G��Mxz$��KY�pFT�v"Ol1�$dÿ>�P�V�3B:���"O6����fp,�q���{R��e"O�QPWi�1{�xs��&���@�"O>�с�Z�iP�4��)$�@!"O|��F�u�
��S���e��"O�d��M�\?���*�G��	�"O
�h#c��q2��ʿj�B!@�"OP�(CeĎ�,��3�P	D���"O �q��ҝE)��#f�]4|���"O.1�p뎞j����%�U�((]��"O:�뤠W$j{ư#�$�a�u�&"O:�7J1zUz�8�L���q�"Oz��tJ�2o��Y��ҭ4@4���"OX�a�������$<t5@D"O��كMB,X莬�t�'pFx�"O�)(�L@�n���
#��>��5�c"O@t{dl� S����JE��L�f"O�] a.4���Ā�<�l4!B��|A剤q8�Ց7.c�T��0
V�<L2��פS7`עM��I�Ur�u��J�i)B��j� ��W�̿z�)�S��-t��]�b����wE���l����@&�@���F�& ����1��^αOx�駌�CLq���ǘ&���to��G/��(��1`�z�k� � wFYz�n؞48SEKsN��2.U9&)�=���R�sմe3��KA�'�Ƥ(�,U�g�D�1lD�p6��
�(!��\��B�I�k^���IS����#eA�#~e�"<q��\�W1O,��O޸���&�~?D��c�>%�ȭ9�d&lOl�ң��uG����\�!�`���n�c�\�Z֣��B�8X"/>i�հ�4�f��rZ���W ��j$�@�~B��($�ԐE�Ó;er)�� +��'��,
�B�~"�i��K���L����i�l�h);��������m������@Kdi^�U����a.�	�p�;Ì>��q���E�6 �t �#���a�c	��d�|�C����J���fݵ!,N��3읤$��(�-��
1��2R�v�[�R&�a�U
KdؗL�~�N�o�,>����'�Tݠ����^�!"̯�_t"�'��K4e�!r�5�AG�y���ɝ: �r)_ �t���)J4<�����")R0��R$؈��@˃�m?>-Ц�-M���8�I&4ӊ��;O�UP0Ǒ�~J��3b�"�rU�������RI�<��Tj�����|rQ;B�����7�A�	@(Ļ@'�cTذ���1��ۄ�S�O�rPE|��T��x�R+@6 @���U�KsLY���-a5DC��~��2K|��6=jp�OyJ�c�KI�e�1�6�
U�� ��?"����cp��&�V'7�5�!ER%j馀l�\�4	����|�$hI3��'Bc��@�M�}(=�P(���3ۓG�
�˂�"����!����WjR(z�����6 ��q�[oy�+X y�O}JLAG�Z�P�.-h�Á�O��e���>- � �ү$!F\$�ĦOF�CJ��y��ss'װ~+�4)Fo�$ ���oKw�r鳊=<O����$ԿN;�iV�;�D���Z��B��H>��U��2�I>��Y0U�D�։��~�����.q�ĈY�GDh<����+zӦt�f�*%FC�N��89� Ey2*�72����F������(q�) �K�%*�p��$�E zȺ@-�EP\1��_�Wj��ZB@%\�� ��ANT�ymi��'��>~�P'��2B�(��S�4O��d����&�M�������&�O`�)Ch��U�\��3� w}n��x"�ڮ)�<�0BS�4�� #vc�<Ij���V��O�4�Jg"�V�� �ʎ�OT����]���RN��%��DiP�?����-ڟme��{U*�]X�T`VR+o�`V��/\j`ð�@%"�0��v�8�O��#F:1�0 L.[�j}��~x�ٰ M,�?�����Ybʎ�u��a��Ė�Q�ʑ���^s؞�P0�K?��i�̄=o���`���({�����^*�D�7�r���.X���_(�T�X��il�xa�>u"�I�ʈ(T���Ŧ��B�(���B�
u^X�u�Yi�O7#]9�PHW�� Uj��p�>��/D!M�T�����1��<���:h�R5�ܴu7��`��Y�,< ��o�i�#j�z�ج{J<��k��Ja(iӁ���( ��BŁ5�h됎�]�
�˅8m��H~�
:i�9���I�<�zT&�"�\�ᐁY�x����P�ҏ�"Ph��TN��D���>O40��.ǠGr�<���7Ha�Ԣ�J�lr,8��ݱ(N�p��O/N�$�A&�~2���4w�&2��Ū��ܣ 	�r蟨{ך��!N�j�L<	���MG��Q��K1_T6��A�u��1���܌RPJ��T`�(?@
�'����h��9�v����Q��խ;�uWR9V^���P�\k��� ��9��<j�`ͪB\�:�V��G�:=l��{��* `̨JL�zNV�'h#���s�P�Y�hة��ϔW��0òJ�9��۵���>�ll8�#����A�kx��e�޶H�ͻQP���l��K6}a��2q�Υl�"Ո�0�iن/���R"�əT#�O�����țP+�-@���V��`�I�pv��Y$N�=�`k�Q<rQd�c/�%"��pg��R�� ���_�	#u��x��ae�.	��	l���'z� ��F$4JXܻ�+N���i��l�܋�G�:S�	�S�A<Z����'؍X�D�����_5�x��� �b��3�l��"�p�Z=	�f%}�)U̟�x�
�fVr6�D9;!����.��rҡXC�[�c���#��ޚ �D
R>��!��$�'hDi��I�`b��ݛ�蒇
XDAJ�ł�� r7�ϞW�>Y� E�Y�ՄJ`�ؘqF�7/U0�����%;�(5�f��}�\�T�O1v�.�+MW�V�2�����I�(:R�ؒ���,���'��a��@g$�P!��V�K�����qD1���jem��D�@�rփP/'$���!��y<��U,,ch|�ac�/�vY��+@���0���H���C�V|��_���Z�捿<mm襯��P�,J��؜�^��ժɶ�p<i� �##��B��(.�4�U�wO�h�s�>)Ba�O�ɑP煐^ ��mӨ`W��Zz�QP>IV�m��$�#��ju�E�d\��G��²hq���ōW5�D�� [
�{��O��X��a�\:�̑$���20���V��i0C��"������zV�u��	��f�$�+4�.x������I:�z�'Ď��
D'��@G�=��I�u�у)O ���6_��T#t@Ɇ�t@b��B������N7l��B�,5�t���^n�U!tH�d�'ܜ��V'���,qP@�	re�}A���;-�[�!�2G���{�����~e?�TdJ�
�*,����"
48�V��CT�0 ���
�Ӽ�6(�����ӎ�;6�
��Rt��_��t�mQ$Hu�q��6fL�I�,X�2�脘o�<�&LJ�Oq9�P/�!�0<y�!�|�����:!�jpJ�%D���¤K�E�t��Ä"G@X\��.H�4=�J֌8Dh 2��d����C�! t��ǌ�X}@p�̌=��QAda�	5���jb��
�|��'ꀐ����#
������j,M3��dɦ7_�<�NαL/�`ψ�I��L:�'l�=�pj��E~���gنw��P@�ɐ�&0kC�6o,5Pb�/X ��b�v���c��"�E�w
>�~���ۏ7k�q;�Y7B�P���"��:9��:7.�� R�1LOrY�q&F�����H\���pg����O�,5 Y � =�!C�"���qT1O��C� ��x���"��+�tx�ŞH�=!%.�(#H1@��ϣs��}��Hf?qV&L9[�p]����J���`�Y*cmҴ�	�'���4�
�.��Ip\��+
����d�I'��!��C쒝��m@�������Ur�L�7�����M4#p��DK\%c�$9���˞��1Y�́�X~BU�c �5	K�� ��QB���/D�z�X���۾E��0[��	F�&��a$X�
7�MJ�ğ	h8qb�b�ZF�����f�'E1O�x"�,�
5V)�6�m�v,����b����k��*��hy0k�I^k,I�^��R��w���Ru!�Z���?�Kԇ:H�d��%i��ӭ�
P��!)D,���@�p��ѫ�@V�V�J��?9<l�Kc��%ᨐ���ʺp���?Y��5\zh�p��ʓ��P#qoS����C/f��5�6���1���lX��Z�i5V��bKG�yf4QچۑK\1Qc�	,�d��?)����>�ԲL�*=���P�b��ث'@Q[A4���gA	�����~
�Dx��-$(	C�ːP��C5��.+>�@戂0��q��k�W/�!Ӵ���["r�����[�@�q�J2IC��_�P�1qJ�mS��q×%���h�cΠ8�V��X>�)�o�O��(FkϢ|HV��2-J�(�� �a���+n`��>�F}�?��(Ȉ/ц��o���L?�$Ea�2(3Q/&�<�&璊k�R�|�MȟdRb*��&z�E��*&�L�Z�ne��\Y��*tGZ�9���1�F}�ʴ�OFD�O�d�hԣ�=)����-r|�A�E�Φt������S<l`C����mH �>3!��f����m+�3���'��}j��N�M���eU�3�z\��O�-|؋�� ���']�Y�)��3z��̲��]=6w̚ �ðb
��B�;��Ey�'v�͘$��П��"-1��qP�ν?�u��Ð�iRra$&O:G�����_�Y�л��S��*F"=§���i��D�Gi�&~"����0EQb�Q3�5T�M�a.�_�S�{��$�4X	x�s��؜	�µ��60�I�y����'�M�#6��;+�e��N�sh���+�tLL=�O6OlTl3��N�;b]C���O��g�i>��C�Z��|�r�d��[%��{Ĭ���K� b��
	��S!�>\�?�'f�.;v@�u΃,jfZh��hן�gD�ا�ɓLy��O�0��$��&�v�Zb!�jР�do3�2j�b�e��O�)�&*�С��w|���Ŝ)��
f�֜u�y�)O�	�#�O����S��K@x�,����5�<�20�]?K���<14�M+����/�"8���Z����<��<a���5v��9��[�kR���a�Q8��cW�@.��HSVk��c�X��u��J��D��Tx|��V*�:
��0��N�K��	/%���(O��I8@p���Mܡt�(0���+��i$aSd��8h�
.u���P�Sn�cCr�  M_7S� ��	e�I5W�0$�B�=��"~�'ㅑ*�<���B>z0͕�<�^K��أp��A(�J�n�
�^)�V��a�����nϡPC�q�� mm�ɜG��"|�
��`�G�W���_�C��q!L7�u�
��D�ΈMxzX�+!:��m:� Ne�4NM�Z��Y��μa�@�U$N��d�l_�qO2���� I�1r�C&R/"pXs�M�,Z�XYI�,갴�AHQ���ڪ�dS��U,
BA8ĮL6m���A�(b����HP*�y��n*a�	�5^�>��ԭ(��	
+<|�ӡK+�`]Y�eR,�6�YP��gD�[f��-���P��̰E�� zBLЛ�M���X����[2��Y~��4�]<z
��quL�?F"�9"kټk��ġ��H8GTA�g�'s��;G�\e+&3Rq���L�Z�3��T�iB�SL +���OPp!NX[L��Ee	|�汁T�г��O���fbOjH�A2���l#�i�4�{��T�DZ�8�RV�W}���IB�s�I )pq�'���E� ���V	F�����AR�3���ǫj��*Q�X��y�O^T�/@�R\@���ޣ#�d����i3�%hՊ
*���;�'z�5�@L� M�Ls� ΝF#
�9��~n�G��5U@�}C�H "i���'��r��F Zm�\�G6�m��)	w�h��.�?B08�c۔���0/O�)'?�:��4?!�y��h��>���ʳ%��cp:L�ʊ'Y؇�i�������2P�A�3C��
u�Ǚ-Ch�1�+�<�#ŏ[�c?�J��ƛi�x�*�t(ȢML�|���%�3,O.Q �M���u�C���p1�
 m�EXS�ݷ��rP�U>S���CT�K�1��]�'yL��a�2�kc�J�8�t8*�ҟV
� 2�����s���fPw�IVgؠ�CO݀.�K	�\�2��r�
�7d���'nA�<9�*N�68�82�E�َ؃'j�П4+d�î���a�^���'��j�)��X�p<Y��L	��Q� �߀F�H��׳�Σ<�S+I~�P��w��e�wm$pg�<I��)���87 AӢ�Q��=�o��`��|�$9s�L��*�!��O^d�&�,KAL$�&dY<2f8��ĕ>1UG]4 \s_!#��,ܠ����7A�0����
(up�$�%gEJ�IPF�Qh�A�2]pR���^t�e��;%f�����Y!nL�o�>�@`�%ax��90��|����&B�&)�U�)�1a�� 宄 �I�|6 ��'(�y(<�7ɓ��"UbC�� ��Xd`x~^�A�����"0z&x�hA��?�}ÍT�.�Y���D?|�dL��I�v�<�BNQ�5ƌ4���0@�	L
md�[g�X3L�A�	����|
�	$}��&h��y1�:ei:�j2,��Pxb �I ���@'%���HhD�P��̛ ��NN
uPV�N�dF���'ʆ�z"�A�n��&R�"S�b�'���`���8x�7� , Ѿ�`�'̀X��@^�0�Υ��K.ݨ���'�֕K2l̓Kn`X��j(a� I�'$-(��P�sPlz�/�81=�9A�'B�(�'@˫�>iI����'�fQ����5( ů��z")[�'�8�a�?�sd�Z.<��'�4q[�l*0MD�0�A� 8XX�:�'J���V�ycqL�(.3�� �'W��J�;-�����*���x�'��@�(S �b�u�W��l�{�'��p�����XC0P�♭">@s�'{�hb�)Ԟa���'��'�}Z�j�	S�*��rb�yJ�#�'m���]`N����I!uw���
�',0pQ��U�A��$��n�>�=S	�'�8��dmʌ|6� Tg�%h����'\�p��Z;`L ]�C	
s-⹈�'	2�;q�ܠ3�̠H��[h���R�'�Tt� C�y��0�'@į�~���'3���`��.{#[g wp>Ƞ�'�6��^"-�@5��N�p}f �'��1e��
��L*bO��K�'̦����<LC(d���WPM!�'��2-&.ڎP8���w���C�'�*���gN'|�\�1$�z���B�'��h�`�	�()tX��F�j5�\��'�&�+Ä�z>�Aјa�n���'p�h���2M�lHA@Ĵpި)��'�����_+VL S�ik��*�'3�eA��N�/_�=Z#�_�^�]�'��Փu�Ή���
���������'>,�ҕ�ʍm��m���O$%���'E�$�sE�1�x��Ǯ@
��� Ƶ�P�ݖyHd ��C�:�M�f"O����|��A�a��|@�"O�Ÿg!�8|w�Z!iT���4"O�պ��3'c$����	3`OR��"O&�B��,�v�R�Ӯ<Q��Q"OZ\�1�N /-!��U�(O��Ӕ"OF4RŎ�Y�j�c&�0^T�m�X�<)��4g~ء�j���P��N�<�i�7)�Fd1���CV@<����I�<�CH3d�����8K6Ƭ9�Oo�<q��*���v���+���y�Ɏm�<��㏮��4�'f��y$��K�,n�<��GA0�����m��0�Y*F�v�<	2��Y  V�6@�ly��Kq�<`��>(�"�`��3P���LCg�<�VƎO:�����*6��a�L�<A��O�/O�-�UL�mxJF�H�<�O�'�T!$d֪o����$�A�<��#1��
�(#|cb���z�<��HN�9��Q�S!w���ٕLQK�<��E#(�E�
���B��f�{�<�S$;��i�*R/v���8$�u�<IT@� )��E
f�,3I0� ��Im�<�lG�Q��$�T��&iX���.�M�<Wf?"�� �����!�s�<Q���.7z�Y�ݻ!db�S4c�m�<%>��)p!��)�13�E�<q�a�)*}H��Pj\�d-�@���D}�<�+��,�*��A4߂Py��UB�<ᠤ�q�h4�Р�3�)���<A�^	g��C�i�@�v��A.�y�D?�S�� 5�Z��L?;�[W(͟y�̅��؅�m�?#���CFJѡDc踅ȓ#��6.��c���$
� Y����&���u�M�y.~t{4hەPq�(��Ӫ�s�6H6�4z3���e:�\��"O����B0T$1+���d�x���"OҰ8�ψ%�Kف=BjQ������yH�dKf`��o##qX�Y����y��_��x8d��G���J�㍣�yb�y5��x��
z2�cG`ʞ�y��E�=�n�z6f����]�1�Gh�<рb��4�р�@�j������Pq�<���� R$�T��a�|��AaD��d�<�T��9�(hc6-�won� �"�T�<��-�8?Ѻ���LӶ&�0���O�<1�M��E��1>���#7N^f~��)§nEbI�B��EY��p%ĮO����ȓD�Xi�D��>P�G\�e�%����	e�Z �JSfX���E��}X�B�I�N���PD�M�,���@��-v�hB䉷g�&��V.�)��Ȁ��
>c�DB�'	۸lJ6�B4��Ӷ�	0/R2��3��$N|J�+���7v�2qcN�E!�ĉ�Xb6ؒ�I��Uή�`3#�=nw!�$S�4����d�\�����&-L!�DB�+0�N�37�����
�3!�֎���Nj��,�7�#z	!�,4;l�w��+t��2��
�k�!���|�	����=F��b@`�&�!��]5K�4�z��$L���Ζ S�1O���$��'�)z��%�}@��%H�!�����S7��A�����\<Mf��Wx��R�W��޹��M�
�li�m*���)� ��st��3e[&���-I���w�$4��8rɎ�X?���e��J�R�h�%�����̳s�FE6^�b`�oW�
U�d���G�d�fF��J䣏�oj�0�5ć�a!�D ���H
6^�7��0���d^!򤇌?���`#ԥ^Hh�R��fj!���2�q��_0+�͓�e�!�����p{�	ϷC
-�-�O!�ę7~���{-W:��U�љC!�D�C*�!*b���m����'��b!�d�.�����#T/�H}�(��=�!�d�9lc�10��}p��f�����rӘ�D��(SA<��H�l8�8p"O��)�l�7T�����q"�X�R-�	N���� q�s�<[��Xb&	G(/��C�	-���ڻ@[��c��Z+V�C�I5�(�	+,J��̀p/�%��C��43�x;'!�I��<�E�b�vC�I�Q�hi��E���x�&�>"\C�I�dif%j�G]ZG�|�SD���B�I�1=�8P��J�8<�,�"��BۈB�	�B��Q#aT�DnژZ7ş �B�ɓo����%!ґ�`�"���z6`B䉯*'����h��A[C�[�a�fC䉮P�Pz�Q���W+Ԫs�H���?	o���pfT�|A�,rSl٣n6���ȓ	?�8���3�6䩓ʖ�}%�%�(D{����ݓC6��hVo?2m�A����y��J�^���녅�?i,\
�D�y��G Te>��ţ�+/KLuY�`"�0?�+O�\�č�)��q�F�(m6n&$���V�P{lr�٤E��H��"�R��y�'R�,�&������l���y" �h�����ұu����µ�y���|��-��Xsh-{��4��<q��J
�l1�U�ܬFw�y+�-�5�!�$�T�bQk�L�KWf��,�%�!�d��o�(�����4Z.��s��u��h��JW	B�b�o[8�<�#fG$D� �b��v���6
�D2pY�0�-�{�?��� U�(��L�����fq�AO*D�d�zh����e�+VxX�;�e#D�3�`�+~*�rTՏ?� �	TD=D��9����okT�@����!����CG;D�P G��SR6�u㐿]�Ll�V;D�`����t�82���# �+��8D�DC�ά@��p9A�c��Ak%�7D�dB�Aږ'ƌ�p��Ao:ȝIs�4D�d���6;&���ʓ)pV]�&B4D��B�kz��Qc�?���9��3D���6��9+� c�ɍ�����2D� ��� �&����|҂)��l0D���z���#�� =��c��0�y@�;�zX���P8��4hu'�(�y���0'�"��b�_=[$���	��y��L�,n��9P����A�˅��y����<b��#$&Չ�Bp�gA�y�#ъZ=`L��h����j -��yr��ht))\d�fD���Λ�y¥�G���&�N$e�	@� ���>��O\���T�Q�	��iG�.°L��"OXI	G�ܕ'q"}c����'��]�"Ox�cDb9}��#F��!��R"O���N-�|��C�D5�a¢"O� ��U��71�#����Hda��'Q�`���NWO��1��ưI�X����#D���o��NQ�⪑):xX=1��!D�����۶"�p�y�I,l�b�a��>D�<p�n��d���)��?�F�*�"(D���EE{�\�����;�\H�7 %D�h��l�/�t)+��I48 ��=D��f�6W0��Pg
���4�)���<9q�Cu�}�d�p��M�� V�<��/%@~B�3��3��=Y�Z}�<�U��G�����/\��	ů|�<	��R�r�]X��çЪ���k�y�<1��@h����Խ~�@��k�{�'Q?�̏�(i4���ۼK!�D;D�PC�A�,I`dD0iؖ?2�ơ4,O�X��057|�f+@�C<����yҬ�,D���L�s���cA���df���>���d�5E`��ň.⾽��� K�!�d�}d��`� gl$b���y�!��Є4b�l �.�/)��Xh�$t�!�D��I�����2A�AA�R*r�!�$��^���a���H�`�!���$Da�H��X��8��'�!�$�UE<hG L?�����Y�!�X�~`s���%x�������_!��� ��;4#ߊ!����G�	�G�!���-��a��A�\"���++H�!�$�W�\+�ʃXtU���E�!��n�&�k��U��@2�F9%Z!�䜞2�d�"�D�J<�8�A���uG!�J3W?���t@8ށ���p0!�Ќ$�pX�K�T*�m���NR"!�d#sqLI�eϥ]D	�c��C!!򤐚#FRt�'f�+������:!�D�/a�\h�D-L�l82AR�F�!��=�JT��_�k>�EQ�	ƈ'�!��8N���8bC�	y�j����f�!�U-
�B�@��p�LAx��ޓl�!��|%�-�� O�q������!�DM"��br�އ�hm����G�!�d̞���ܵ)��cC ���!�$�!}�E���,ndD9���|f!�d�i螙�S�W�k%.1Q��(tN!�d�n��u�݈q�@akVG�*#c!�;W���Єɉ(8dR5�(�9nX!���\����'��3t0Lڄ��I!��/THFl��T="fD���@;?0!���m�l�r��)0�tز�Ē�L.!��
�%o\�r�*Ѯ8�2�˄��	�!�

v*�go��E��X�FNF7[b!��
_8�eRHp�gCK!��"���[��K�xa���&�!򄏴|��yzuM(Gz�õ��N�!��G� ��1��F((_Z�Q��st!�d�z�z#LGjy<��!�/t!�Ȇ`'kL0�D��b ��H^!��7954��%��T�|I8'��A�!�dA3g%�9�c*D$W�P���	w�!�d1���i�,��=l����#;!��c[����*7440`��$#Z!��/D�{ (�'C������n7!�$ӱz���X�%�0`��O�<!�d��<%�Xȓe�� �><�\|ܨ�'?�T��2z|�R2��#t	���
��� :��7�D�bT���#�]�$ՃA"O>,�qG�&��""C��e��"O���`lM�*��U!_�z<�u"Oh�B0.P]�Y#��#>���ʒ"O�x���Ky�T�t �5 � `sc"O��!���AR�/ٷ2�*m�t"O����>+ԉ%���F�8�y�"O�$0�/��Nl �����\��I��"O8���ϭ&L��[GY/;��y"Oh("����rF��"\���R"O�MJ�!��M��-�ь�:H���qF"OT��W�pp�в��H�$�պ#"Ol���*�G4�0�!Gh�#P"O���f�ϏFIR�y�� ����"O�I�V!���p"�
�2"O���}�����k��e7"O!i�
�>3H�s���y�T�'"O����L85T��*U�~ ���"O�pK'�Y�%��,�t�D��- �"O���M�GkX�I�ܸE
R"OT��%�л��
&�8�T5"&"O�5�B��R��Ը7(9qz;0"O>EaQ�,F�C�I 8��"OT<ɔ��%�TC3��<"�6Y��*O^%a��@A���i3�ߥP���S�'Z�P��N׾In�tC���H	�m��''��*"��6%����i��M�|���'!r�;vk����ʋ]��mR
�'�R�:�*H�X�yZ�ƠY�4��'��tJ��I�B�f��X�O�xA�'������8B�j��UL�6`-��'��l��'���hu꓈@2���'�*���_�~��D�C������'��	�*B�JsX�#������C�'w@���'W�܊��!ڞ���a�'V|�7�\�k���kW��#N��J�'4޸2�I�6"��E�L7Cʘ���'�He�,O�   e��b�ț�'�*t1C�Q8�XD�7����'�@�jbaD)+�ʍZ�X6+^"�B
�'��sd�	\PLԸ4i�	l�>9@
�';�k)��}yX`BÍ��h����'�p�B�jL� ֒Kwȏ'3M>�y�'�V���Y���Vcׯ@P���'78��J�9B��d�lH�3ؤY��'b�qH"��� P8ꥆ�(5���3�'[���C��|7���爕�2��k�'/�M�GK�M~5���x!`
�'��h��g���^��r��-+�X�	�'�	kR"���r��ҧN�E�	�'::i���H�$���kE�|T-��')�#t"J�9�̈��B��%����'E��*qcZ ���r'D���|�<�e+J�����Ѯ��)vB����_�<y����(�)�=n$��M^�<��$F,�0k�g74���@�<�"�yd}KW#Ҝ;\u��A�<I��[9L���,N.P�j�zG�@�<�sB8bA�M�6��9�b,�FD�<��B��2�$+WDE��a�g��G�<�0�2;)�Q�lŉH41��N[h�<q���TN��qU�U��~e���Cd�<����|�4���\ ������{�<a�M��&��KD�	!�����{�<� dtk�Ə�Y�~�V��2yp@"O|
r��kA��(&A@y��'��p�婚�)�r]I���,z����'!��е�]�.�LhG���j_�p �'���g�E0B�*�:ʛ)l2]��'�0t��
MT�eIg~��'��X�@���l�KE�i�Nx�'�1D/R�\hD��f|֩[�'�Z8jE�\�T7�@
���Y��x"�'ߪ90R�:a4�{p)6蒤��'ZJ)!va^a$Q��Z໦B�I&Μ�2MT�|sJة��΃M��B�r4��@�Ù�/�j�8P��+q>B�Iv��y"��2��q8�O߈O�bC�I ?_�A���4xH�!��E�TC��o�\�a$���a���3B�JC�Is��!�V. ��Y#6 bC�ɬW�����Mu����!^o@C�	����c�X�n�H5�gX,��C䉍Nb�(i�Xb�m�)h�B�8�2-���<=��ز`R�v
C�	;f�T�[$^�|�P��ϵ_�B��-_��X�p�Le\���I�x��C�ɰl�a��&�4Ac*����["~ȖC�IK����7��"�F �]*|�tC䉺�xY%M�p�N���	1bVC��9o�XИ��@�j�(V��tB�	I����Q���ݮ4C���	�'���2���	�P�gn��B���	�'����r�Y�K�`P;W�8@�@	�'�0s��Q_�HaV�B���:�'L���H�`�4�3UK�����'͖�!tdQ�1�00��"A0l���'7��#-�|M�(�Sn�
��Mk�'�d��6M��<@8հ oƹmx���'r�(dDԕ'���  �W,=(��b�'��1Cp�1nr��@��S�bO�)�'�Tm�Qf��eT����H��$���	�'����S��O?L�"���ܚ�
�'t�L�@�%�\$���'k��(
�'b�0���7"URl�A�6b�x�Y
�'u��@�>x��Q��`�dp�	�'�"L�q�ƶ3xNiطd��Z�����'�����`F�g���ZdL�K��A�'e�(ׄ<q��h�v�?$���'���7N�9�ΘHF*�>i�b���'��H0��v�~dx����o|h�S�'���m��P@!���[���3�'�.x�.��h��R4)N�	zn ;�'�Pq�wb�J����ʴJ�����'b����U+*'��6�	�A_��'ΒѐT� H�m�uK��6�F1x�'xa�d�	b�,+��B�)�|���'�H�`����3P�Ɵm*�\9�G-D�x����4q���emG!~�j萢)'D��1��yj`�vcG�=�f���d?D��p牀9�u�Џv�&<0.)D�p:�D1`��{�D,U,D���m*D���푹�:���jN"%!l� w�'D�l�#�>4#���$M�=E.��P�&D��(��&�rt�&��-/L��2D��w
O�P�ai��K���4D��ApN]�U���B�ʷ[�!��2D����ˠ^|ڰ���I�{�-�2H.D�� �Q���]8NO��[��М "����"OJ	9��� *F=�$g�����"O��`7*�4`9v�ƥ��y �icT"O2]�wd��?� �3��X���"OL��WI��>�IK�aț-�����"O0@��G[ B�±�&*�8��20"O�U3�+Ĥ3��t�<#��Dk�"O�e�w��\�8�a\�v��J�"O�1ۼ���(�"n���"O<�S2B 0�h"�Ǖ�|�6i1�"O�"�]�V�H8z�*q�|���"O�eZ`K�7Qrд�5Ă�J����"O�E�g��}�d��I].\�
�"O�;&�*�a��o�j��b"O����N�0:�8cOJ��v9
�"Oj���!C�sްf-�A��}��*ORsAnR�9��Y�V�������'h����ȑz�T�5�3v�1J�'�Μ�Dk�	zx]�j� s�\]:�'/�80o�3����҇��_��1R�'���g�D���A�ٙ0�݂�'�F<3�>p(�2��G�'4у�'�~��`M'<�x�`��Gc�M��'�9����X�2a�҆:�Ł�'�fM��o̊A4\Y0M�f�j��'�����/�t~�lҧ,��P���[�'d�<�6��nJ؊�iـv4�-�'�S��ϑXo��1D	5Y���H
�'4�X��G�8��$��_g��z�'�2�8 ad��V��i�p���1D�0�B��p����sT~(
��3D�p��й:���O�B�z�:R!.D�\��䝂h�@\��Q�m�,�O6D���m�'
�;Ȑ<V�)	�"3D�8��+��}�t�sg�J�{5�M�G5D� C'dH0���;1�ɓH]lq�b2D�����*�`Ȣ�,��W�U�/D�����ݫ=xƴE�Q��5��-D��hUK��%2hk2O{U�{W!7D�� �$�"g^-A�a��$��T�A8D�Bfh�/���s#46p�ܲ��3D���b�P8]
`���ȸ`�!M>D��@q'D2 pv�z7"D,4i���;D�Б-ϐL�
@ۑ�����i�8D��Ӂ �2z��v�k88 +�A8D��QV�͘?+6hc���N��pـ+7D�����I�ox�8����Dj��KSh3D���F �"@<�ZB�j/�`҇,3D�4; ��9`�N�9���$�A1�/D���dL�@�E�Z(I���.D�x���2Ue�|� F�+�ٸ�+,D�܁o�
gv8��X�_��m�r�>D���cÍ-Aw�k�l[�M=��9H D���ℚ�0� ��+^��w�<D��vn]�=a��#��Z 0uRA�Ʀ<D��h��?Z�P�FAU�X�D�i�;D�H ��^�}���"4lλlǄ�Y��:D���"��<D�_�z��Td9D�@Z	�9��E�O�"ɚ��M8D�t�6N
����#a`�5c�C3D��P U?:!B�ɑ��rIj@ �;D��C��ub�(�%��;[w^��.4D�`��
01wt4���*CJ�(B�3D��h"�4gF�A��B5e�@S��-D�� j}K"�йdА@+2��/El���"O�lHB����r净5N���!�"O�<���+!\Dq5�[�O�l�I�"O��#�D.z&��N^.q�!�"O�Ⱥ@�1�5�#�E:1ȉ��"O�M�$�C$�p�-?+#PI�2"O���D�s����!c��e�"O��`@H���Q�Ӂ�%�R���"O�6矖ڸSF����� ��"O"�����"@w:tiC	<%��Ց�"OJsbE#,>�֡_�Ht|��"O|� W*w�fP���/[���"O``z���2l����儎l�e(�"O�qb��2�@5Bw#E�c��Q�"O����e����8���w>�˖"O�x���!gV��'��)<p�yD"OJ�&���`L���T�%��8�"O�Ѳ�)�/NfMb��Ƌ���"OB��f�zTV�b�Oa�x��4"O�,�4 �u���rc�����u3�"OvȪ!�ݙ`xz�3�Hgzf�X "O9��v��;�LY�lt���"O��cr�G]bE�sk\Q��B"O��Ǩ�<�2|;�ǝ�*2JYj0"O�es�(��t�>`x��ȫ �z �$"ON!���Ǘvu�9J%&VA|^X��"O@�	�h�97����åos���"O��"�,�o⥚�D��'qM��"O�����J���J�����q�"Ot��&�Z���l���S+clzD0T"OJ})&�M-mB&�K7Dو�"O�}q�˗FR�1�O�</>BL�b"O0,	�&�"l����/�4���"Oj5��h�Pe*��0��hBb�<�D�����t� 5*բ�ʱG�w�<Y��o�]�&Ī�m
W��o�<��&�(�,�5K�2Y$�K
Qh�<Y&ԨP^Ll�i^L$���\�<�tk��|�@m�a��g���+���Y�<I���l�΅�5J�z%$+�l�R�<�V�F+5���Ӹ^���J¯�Q�<Q�Ӱj��yS׮�@�dx Fs�<r	�/7�����[���R#lZq�<��
A�l�&ܫu�<rd*Ss�<2a��a��1У �+i���&o�p�<��?g��Yt��K���'O�p�<�S��uQ���wa�q�hY��0D���T�r�
�c��a�<D�@{�F)/�ذ�%Q���H��yB�L�eE�`Ѣ���~��	�"�y"��2-��$�ءD��c��B"�y2��VфO=xupy�S�ռ�y2NU�V��) �:��"���y���p�)��e[�c���{̂��yƇ 1����QNP�\k: ��M���y".F&],a{ddF?&����N�y�̆5?s��S���%h������y2H a�T�ˤ���}��̉*�yRm@�J�ȉ۠�0��8X7�^��y���,e�|�H�����`
wi�y���[`�SbHÑ
�$9 棂�y҈ozE#@@�[X0A�i��yR�F�w����&"{�93��׺�yR�ǧlf�S#��.
��ԙ�
"�y
� 4tI�؞C�^�@�#�z	0�"O0 nZ�p��]@u��PB@���!D���W���칳"��2�D� &;D��p�OGR7!�! K���]2�I:D�x�͘�/� Ա��>�YA��$T� �靊z*�R����Ԓ�"O��ʔ��X1�4�h� bƊ�J�"O�}C � <���(N	w_��"O�5�̐�W���8B��[�H#Q"O��P��Ö2&:����Y4q�L�s�"O&yP��܃\�d�����!�"O(�xҁv�Qr#E|����0"O�EQbO;\ݱ6dŖFZ��g"Ol��B/��2���͕�' ̈K�"O���'A-�D��Oަt���"O�ka�M�nD��G��=��g"O<T13@U,�fQم�D$Zt�C"OF��BH�*3���@��<L#V��"O���C�Ps��HO�!U@�b!�D��
a"]ґꔽ==6蠓��U[!�Dܦ����d*߭	���:���(�!� q��m�q�P4?�i�%�[m�!�DR7D@���0ىR�)珧4�!򤗦zZ\�qpH�MEZ`�Fߚl�!�C:6��8�D�2�ܡ�0���6�!�$��.����5�0.��t22� �!���2r4Y !�9;w�r�$� �!�d>ie&�9&�ļ+ r�JD͊��!�D��WRD4;�̋��^ (P��0_ !�� b�HpCf��(5�+E �ȓ>C\9hP����Iq��I��Y�ȓ,�V�)M�V��$)6O�=6� ��-{FPH���Oچ���E����g^��U�t�\�(��n�d��ȓ)�t�U��f�i��$ʯ<5F��ȓddx�a�3aH`E��~E^��G� X�� �, �ԨC3-AUW���ȓM>.��7c�)ᔁS��P�sl�U��@�"m�sK'2�8�s�����ȓС��	#yt#߲|`i�ȓ
����d\ b��`i���1V�p1��rg�EI` G7vr��v ��1�vB�	8z8����e�Xlʐ+�+	�B�	�=0eCd�O.�{7��
*�B�I�F����3�<�"T��n�eg�B���lq�
C�E������s��B�	W�(�겣�FT0��J�@<xB�	[��B.T	z���d�`B�	^�}����_ ��ʄ�Y�TB�	6F�~Y`��� ~���2�?1�B�I9w�>1WnDyʙb�B����B�)_9���V`�5R6���RL�-�C�ɱWۢ	��H:St��af��|��C�I�r'��p��A/ �,���,�83�C�I�]��t21���7z�p�A�Q|C�	0z-p�QMB���)P `�+Q�vC�	ZdF���p����iЦp �C�Ɉ&����TJ�3(c�����/Z�C�I3p��d���_h�U��@<p\C䉾D6pc�D��T��U,��T4�B�'m�����R�B�&�j�a�2!�B�ɶ.\�Pc���,*�bj�m�50:�C��(�*�w$ݥ�  gb 6X�!�D��B������xzW�Ƞr	��� �-���R4F��8Q� %5�i�E"O��+�n�?O� �W�˭sҾ�q�"O�dh3�78����B�`�E�"O��G��&(Q~UJ"�3Y�����"O�c$L�l�}�.F�l�z�"O��	���;'^d���Og4��"O�ܫ���`�n ��.�_�d1�g"O� ѵj�S-�Eر/Q��b%q"O �QU�ٽY�28"d匛W�P1Qs"O���W���6��r䎷I{�=+�"O��qS���hy�#�3t�В�"O�E�c �$Z�v�h�bDD�"OM�  L�"-p�Sf��uzp�X4"OjT���]�x���;6T{`�=��"O�d�ۿd/J��R��3�d=Y�"OD��c���\,�PKZ� �f`q�"O��I�N^��|c* �,����S"O��	�	�)��m)���B��,�"O�t�ƊI{P�=R���C�@�{�"O�qBB�S�R�LX������F"O���o3;�\�r��7(���Af"OJ܀#E��%
�"�ak�R�٣"O��yV+�����Oҿd�(�r�"O��z���KŤYE.O&Q�d��"Ory���Ea�I8t�[�q����F"OX����"Bl��+�P��]: "O������ K��w���C"O�	`��;f��A*"nR�p���"OH��q�A�wJe�����6r�]"OZ�`Gl��?��Y��J�8k�u�""O\�9v���!Ɗ�[#�_t��F"OƸcC�	F�2�� �T9Vy���R"O��$ǋ�y�Ʊ{�_^��r"O~�ig�ՂH�}����9j�L`q"O6�R��T�p�X	���^:e����%"O�-�g�2F����DC^�`ԣ�"O�T�(�*4��ȁ±|�0�E"OȰ`eP�!vr��eN5l��\[ "O^��FP�=fX�жgi\`��b"OƔ�1-e���5��(C���"Ot-��5!d�VO.a,ڤ��"O������V<���,E�--�H��"O����H�7�)Q&�	�U�^��A"O�\�u��6@P~�3�!�!k��)"Oh�;�oջ\�,�{� ,k���@R"OD%J��Q�a�Q%;C|x9��"O�e�"�]G���W��9ol�M�$"OLH"���c.*�w�T�$ G"O�����^����O/@A�Yؖ"O�t��F�G�h��Dt��y"O6�Tjɜ(Sh����0YT8�"O�!���J,>q�Q�A۶(|c"OL��g�7m��R��5��<�g"O�ła/Y!X�"�ڏ)���3"O�uc�e��.8����%Y8����"O��R1(P�Gl�UΎ33� <i�"Ot��%��8qGFuh�K�q��h�S"O�9��
�V�,p�˸&��0�"O�ݳv.�QoRd�2"H�A���"O�h�(v$|���cR�I�z�!�d.в��BZ�C}&tf�M4m!�d�\�*�ʆ��o�<*�e�9ZW!�$c�$@HKe#� ��̍Hj��ȓ@�,��c�%���!# �?<H ��S�? �)����n<���t�\�BG���"O�xY�Z=8�V�V�N��"Ox�i��N�M��B&�3���"O� �$舝"<P��D�,"N�Q�"O|<�w#I�P��+5��7��C"O��8�kυׅO@��Q��B�!�$�_Y�$��߮H>,lp`N$6�!�N�2|b�o�1�N��#���"�!�Ē��*!�!K��e�D��4|�!�nHA%O=C��#��E�r�!�$1&�PЃ���"�ܓ��TJ!�d�����KdBE c�\d��aW�!�$��h�
����l�D�'�!����p$��*�����l�4^Y!��PIf���q>��
@f�/��Ԇȓ!�q2��At�0+����|�ȓv�z���t���]�\�&4��+�v���E�5)�HB��P�9"B�	�� ���ܝm�,���1B5�B�p�СйD��a�NְWPB��,Iɬi{�&	.B�Js�R�I�>B�ɥs���Bf۵GS�izf�$<�4B�I�H�И팙
^�-��n�^�B�I�{�iѥ@�?Ĭy�!��B�I6a������ߢ���_V�C�	9�6%�3LN�t�nU���?6�C�IC0zL�b�!#�Z�:w(��F��C�I�Y��K�%�^�	%+��b}.C�ɠr���v&��E�� �-1�C�I8i]^�ipljf�9� g\,HTB��.M;�M��BS-v��=��+��0�>B�I:q���3�b�fb�y�e@�� �
B�I +��8`A���Q,Tl��C��u���ҫ±A�[�1X�C� � $��'�~Ԃ5h3�Mk��C�	�7��A	��Q3&.]��(C��B�I<p!^4�F׀|(i��Dڢs��B䉒%��b'o��E�����XIf�B��+W��t���p�*���`�� A�B�	���5����
t�P0E���B�ɾ	5���􋈚^D�ZK��Q�"B��7'_��j#�C)eĆ��A	A:�XB䉘iצ�s-	T'6�+#N	�1�"B�	�ra�rO�Q�ș���D�	2B�I�p��i�@OͲi*Pౖ�ĩ]kPC�I�~Xv	г!IP-��V��/F�C�I����K�LƤp�"�=}/Ps�'�X��t�^!%�
���Ꮛy�@���'�[��W�N@b�m��`�����'��@��g��S���Ʀ�3^��%��'��˂�u��Uj�BՐR �%�
�'H�<�!gP,g4B����M�B8	i
�'�����*��b�5Q��N�8K<lc�'������H��E�* 8� �'���BGQ)��Kð�����'V��v#�4!����Ŕ�k��P�'g� B"ٖ$|P�K�MX�hu���
�'�T�ѕM�3@2�+�oH	`3�
�'��"�a��Vu�s�@'VZ&��	�'���"aό�"��A���	�`�ڬ�
�'�q�"��|�n����	�Q��xB	�'p A:るH���I��_�;<��'�^E#�Js�PC���B� ��'ٮ�[�j�K���)d���,�;
��� ʩ
b�دP ������'�T��"O�)��ƈ��� �Y9@��ԸV"O��3�Ŗe��s2�_�4���d"O6�z�eY�-�a�v(Z�j���"OX��p#ݍx�LuB�F�"jS�= c"O��P� U<�X�vE�i�6`R�"O�I�`�R�~̑�M�E�\)Q�"O�Q���kڔA1Mݸn�V�*R"Oҩ2G$�1/,H���Q�#�Zhy�"O�Y�;n3Rp�F+At���6"O�p0I�#e�p���d|U��Q�"O���U��*?�P,�Dd��l��"O*������qN���AK!$�h�"O.,;��/o ��*�u"O��B���lFQ�p�p�Hy�2"O�qZg�l�V���T{����$"O�TJ��@,f D��ą�Gh��"O^Y�oZX����ÙGfV�hw"O�$yF�Ju(��N�HZ2M� "O^p	��͢e�hA@���5G�՘"O�MGZ�jnu���7(�-p#"O~�9��W�3T"Pa�&���ʣ"O�=0�e+n׎�P%X!	~:(��*OR&�	$<ȝqS���9�+�'��C�mÊl޸2�T	,��Q�'����䐉~P(�r��
$A��A�'�6�����^����E�,C���'��0�TGX$XA�i#6M-&H��'m�ǥ�"��A2��=u��c�'	�:U�j,��qPʕ{XD��
�')rMk�&Ȓ)�ػr�3p�P�Q�'y�$�1C,~_0�;�%JoIl�C�'i{��կ80�y�`�����
�'w^8� ��h<x�n�,?ڔ 
�'�d�3�O�y� }�`���0�+	�'!BM8�W�	������US:B�I�,B$a��l����?n��B�I�GF��C�9I"��
�o�	��B���*�A�،g���:��֡:�B�	�xW �{E�G����`�)��!��C�I�g�����fB�_%����h�?��B䉠L��0�AD3d�n9�a����B�I�m�X}Ç��pܹ䡎4k�B�ɝh�z��eQ�<�`d�r��������h��N+Ղ
�gҶx�,��ȓR�n�xfb
a�H�j�>8��ȓ~���c^,p�FP����2oĵ��rb$���L�cKla
����=HFņȓo`��P0��=,�v� 1��*-"̆ȓ:F��",O�w,8X@�	�e-浆ȓ �İ��KG\�����e	�q��*\,�ti�n��y&o �:D�ȓB8���G"�Ei�,��J��+f���nH&|��$� ږ�����u�(}j�%ӫ6��0K"BX�K	 ��ȓV�0-3v�VH��"uA1Q�ȓI��#b��*�����Z	3�r��ȓCҕP 1<�@q���v�p�ȓZs`z��+X��1)��V�`U�=�ȓ%a&�;�ڭ���q���C剓iC�1��`@�?�a�-�C䉧}0��rF��d��(cт)`�C�	�xZ,JA�Γ2�DIW!Z�g֒B�I�f?|�hgJF|PY�	C �B�)� �d���E�m@�L�e
��ܻT"O@���G�n\ڔ��0R*�Ѳ1"O��B�C�j�f�8S쀭)�e`�"O��*�I�?ZDŒ�J
1T�D| �"O�0B��	^i��K�ʃO���"O���nQ�v3^�sы$47���d"Oz�S#✼G\R���#o;��
�"OJ��#��;�N%c��*A:�"O���"� �����ǠtT"O��AbE�<k��w��(U��"OL0[5��z��|�5��7��"�"Onxxt#P Jب���6�$���"O���� 4ٮ�J4ꎕ7��j�"O6�r�k� H��#�Q6T�"O�����d������3�a�TG>D�d�c�&%
���EE;j/p��rc=D��:dI�C�|U2�#4B��I:D��p7��v��M�bh׃}�2�(��6D����'�!(�3@葯%�̹�u�(D�� �!U+
ʡ�1��w����V�%D��D�H&q�( �'�����k�� D���q.��b��d:��G*6�)D��hJ줰���B= 7n9D�\���7rL�
f"O<��e�6	6D���WI�c�p�v��vm��#
2D� ����.H��Ps�U��g=D��� n*82��	=] �QtM9D�0X��]%K[�5���9HA��S�,D��ɓk-�98��D;>�v�2��)D�����O �1[ҭ�?��� )D�Xv�&��c5 �#&���%D��b�ʔQ����Ξz"��C?D�t�7��L��4�-�%�!D�h8����V���#f��bzI�� D�TJ���\�8��HXXPƢ0D�l҆�1qWH�[ L��D���s�+D���v�ԗ�d%S�� &.\�1"'�)D���5�I<���� S�cd0B�J%D�X3A2��Ȩ��*A*�i>D�(r2�:��mQ6M�#3�E��9D��媄��Ȑt�6NHƉ��O=D���AR�p�JQ�6K_^,�5�� D��@�L��y���d%I�\J��	�-4D��Bǩ�/6����(B�-���2D�dja���K5Ruq�"��À�K/&D���%K^񊉃t߆5F���m%D��x���f�~P"wl�2�XKb%D�k���A��LH�o�$jht��!D�`�׈��a�(��I��\�XH���=D�@��hէ`4v�Ƭ�4�^�:G�6D�!E+SX����n_	w���J8D�x*��ʨ3��Xز�:PsD���2D��2�J�f�-kS�ݷ���+D����x:�CO�+
l��"�+D�ԫ�!��2�Di�G���$H� +D�1�.Q�l��:׍W�2Y��X4<D���Bmф_W�(&����i�8D���@*�0��@�ȕ�'.�TX�#D��-��UR��-70�C�7D�h�bƂ�tQ��B�:_c&(�+6D�d�S�0>>i+e�DQ*�xc�!D�K��T�x�J2��-��x
�#D�4I�e�6 �Jt�x: ���#D�P���/!��D0D��P���;$G D�� ���̙h�V��tU8���D"ODl%��g����b#(I�"O�ȣ��/]��)����Omn�Z"O�M�w�"7����ԬC0	��d#�"O )��F�$-��32N>dپ��@"OT��#"�,P��=QE";I�0A��"OF����%�DtR� _10ĸ��D"O0z`GY�v0"t�E���Nq�A"O8M���&C�`�d(�]��P"O����L�!~�i�G'�ƴ�C"OF��f�=!���0��V.f���"O�`�U2f�(��c�A;k��5R�"O:��!��d�b�2g��!T�ҭ�C"O�� ǊI�F"�`��R4`�̠#�"O2�wm�> ��ѣC��1☥��"Oڤ{3��kX�"�S:�t��"O�����X�*����k܏"d�x�"O<uX�Èq��M��
Ii�ak�"Od�
�DN"��1(��T0��0"O��G�1C: y)v@�4 ���"Oh1sCH�v�ΰ��T����"OJy"���< `7�B8�|;�"O4�[ `�;����O+#[2�
�"O�����9V�������>R~��1"O���AY��b��
�jl���"O����C��=��f& ��q �"OH�v&�6x~L�W(�&\DF=Pq"O��"�@�R����Z� )����"O2�S����r[��W�{���"O��i (��/�����'= ��X�"O�١D
 )<�XCu'D� VJ���"Ox�!@D�j\l�	�B�v��"O��pC�	�-�d	 �Ô�=2<���'��uA"��;fh��'�4���'9sg� �49:��r����'#^QZ��G���HUK����
�'��tA���7e^��+L����'�p���㞰�%C$F��X0�`�X�<��h�'?�%x�ᛡ�Jܻ3�X�<Aq`rڄ�ۂE[7�3�)\�<yB��� xP���S��M��T�<��EC*��JfG֙o9�su��S�<�q���R
2�Z�>"���Jd	�E�<�U$��:'��SAC��1�r��E�<��O=DE@3H�jN���J]f�<iV��"MܜK��{@6��w*�_�<ya`�'p�p�� ��u��h��[�<��H��# ƀ��-�8u�T��f��W�<1d�ĀJ׾H��*�20�h��V�<�!�ʹ3�$$��Y��X�JS�<a�O�	~O�9r�H���,ҵ��P�<Qf�� |����W��2U�pc�#MP�<�������F��� �2�hRD�<���)&�0e��DĶ-r��B�<�ajU�af�[:ְ5��Lz�<!L��5O���f> ��Q�-�w�<����V���LB~m���' E\�<�QF��u�<L�Љѵ@��5��
V�<�BM	<9*�Ȁ�4?�4acS�Q�<a���pr�`�٠N�f�%B���yb.�,���"KG��*d�
�y��>c5`2�`��H��!�cï�y�����y��;����e��,�y��> ��!"��)rJ�YХަ�y
� 6���H�(B¥�æ�>����F"O��{�j�_EU�Z?��5[T"O�����	|Ȯ�J��@�g��Y8�"O|=�@T�n�e�
��u$"O]4���j��Q0*��n��=�5"O$��f�>qq��`�ILW���"O4�!�� hM9Q\=# �m��"ORd�
ߧI��.�	����"O�ZCb��62)�3� "*�4` "O��R5k,HL�4z��X�.3hX:s"O���&̇�1����IA�&�&a�"OdD��	Q~n��H�"`� Sv"OĤ�`MA�(|@�D��<��D 4"OV�j`#B6C��eۗ����д2G"O:�0P*<�&0Z�J�0h�,��"O��9�E7 ~&�s$,^� YL��"O������ڙڂLP�j[,4za"O�M@ �Ɨ��b%�ٴ9��X""Or�j���(A�-�s�ڛ	�0F"O�u2��Π���\�*��8�"OL �c���d2�CJ�=^�5"O��㑌*�(���U��p�V"O����IV��`l�5�2�@ �'"O�]�sj�>$��	�!�ƤF�����"O J%k�6�jl1�k�3��Z"O@���A�4�"1z�T�]��`s"O�0��!]���5c8r����"O�-i7
C/9�Π0���(R��q"O���E�a��UB� Cٲ�"O^}j� ĒO'��rE�G%`�컰"O�}(���|8�r�_9I�"O�Z�����p�bF	
p��&"O0x�dBL^�����$+���YF"O�Q)��(�lR�� !D^��"OP��C���R@��q!$^/L��8�'x�C��^/.^z0A�o59����'��e8��K����)I�eDX���'������/e�^=��m�Z=�Lh�'��	w�߁jh�E��&SE�5C�'T�rӦ�XH��*�(����1�z\�1K�Q`�yFj�H��p�ȓy��Jc��n,�4�A��@�tm��6V,���iVȐԢ�(�tU�ȓz���B�gTQK��A��:`R>؆ȓj;"���F�U{� F� K&h��;����$	�����C�SX�-�ȓ]4����,(� ������D|r8��k���bjy���)��ͧt�z���N�j����+�M��Фw����^i�]���'#q<-Ps
�""�N���{^���1�����d��(�`��&���2�X�67�{�/�9yS�m�ȓDn�z�@7TyZ)��FC�_8��P~r1���.Ȏ����P�qCzU��2gL��"�1|@����W0:"4��&Ҁq��'�W�r�q�n�!`���ȓ?���c���Z���z��أB8 ��ȓ+�D̹!
@�#YX͒��@�0}؆���qa���9
��	Ǉ�^[fq�ȓd�`��r��a�x��)>༇��N!��gE�?�n<9@Iʉ_� C�Ɂ&6�@[�� �TZ�M�}�:B�Ii+��P ̂��	� H<8�'�K3��@�t����Gd�YX��� ����B�cv�H�@�$?zl){2"O�������ԅ��� m�U�E"O�`�Ӥ��8��"&T�6tr<yv"O\��A�_�b��+�%H�M�%�7"O`{d�Z��Ī����h�:U�F"O�b�	��+�ܹ��-��)�ΈZ'"O���A���/
�R��H��%��"O�y���3Mt<�4Ȗ(y]Z��"OTQ����$E*<�#ȏ$!0\hu"O ��B䂵
-f��q�K�g>��A"O@�	�f Kt,!�D�09p�"O�!�D8D��UI 'vd��"O�(2�G!nh�'ɾ_�x�"O�����[���Fi �Bjp�%"O���7Yf� 5�D�&]��:1"O��Kbbj��+��κ`Z��"ON �Ϗ?��A�d۔h=,aX�"OҌ�u�F&~��pҍJ%ji�$"O2�9Уа2X,d���u��%�"O��eGP�w`�ѦN�2�*�d"O��z�ǂ"�BP$d)S"O��"�Y�,��MYbj�^6�E�4"O��I����1^���ϖ�Z�m��*O��֢\*#k,h'�ڈy�X	�'��P����6<a�H7�	��2��	�'����uJ�5:�97jG%z���'GM�Ӣ28(p��7�E�U����'�:(㵫i�u�D/U,��
�'�����
>�ay���S�l�y	�'�88��E@k6�d�U��B	�'e������� iߍ�aj�'��E���	0�9Ch�f׆���'TA��?b�����܄Yk@ �'���Y���K����9P�]�'E�y[�&%q�D�g �5lR�b
�'��mp�ŉ��x�P�֫5)z�
�'�1 d�Z�aY�$�쟖@$$�	�'2������/@��f�$�"���'_�%�R�"\� `u��$딄[	�'�f1A�*ǭ/��i��-ĭ>dM2	�'���� ��6��s��"Q���	�')8a�����v3�3C˝�o`9��':��"T�Ο
�F��b�j����'ijx��C!5!z�d+���q�'�p��Μ�9� m8L> BP�	�' P��D�p�"2�	�Ą+
�'�P<,W;g��� "�'gU�E�	�'�Ơ�bHK�RZ����6j�"!D�P�"ȝa�XpdD<a\��r��)D��� U�\�r�-ɱ���`�4D�0�o�3R�(�� B$�=Q��'D�d!���)n��X���O<zx��P�%D������5$,�]:�
�;B.�p�7�#D� J �J�y�wI�4t�Ptavd/D�{����~�n��e�#�tUr��,D�,;�LԸ9۲�cR�8=B���O+D�$S�䗽p������(^�k��4D�(IW��w1z�
C���sz��q��1D��Q	7�`lq��;(c� �E�.D�DI ��f���	r�_�=ӎp2
+D�P2e�#!�� ��(�{�,D���G� ,J��f�eHʴB�),D�4�䫓���w�5\�p��'D�t�&G�N�^��B�(R��p��*D�� �TJ�+S�ì]�r��z:l��g"O��8w�$$@P�C�ޏ)<�51W"O
��
� )%�8:0-�%mI`8��"O�x��A"8e�zDL�*���"O6��,��<r�L�7�QU"O�MJ7��G�ʵ���ӿDSj��"OЉ['J�T`R����4�(�"O�Y�$�0-c�@b��^�C1ލ@"O±p��	�]��t��b'u|Р8�"O��b���~�à���	m��P�"O�ՙ���% �!	�x3"OA!B�.D������t��hv"O�%� �
�BZ83�uwjR�"O�A�%�E�ߌ@����D�@�"O���@�A�Nu��Al�X����"OL�Vh��b��PK+pE:�P"O�uBԉ�|�nd����m4�`�"O�=��s5���V�'n<�"O���Vo߁6J`	� �2C��"O�@���N�Gztx�f�y�W"O�p��e(��<��C68qv�"OB���a�v�Bt9�lY��4L�Q"O2�`���T��AT�ȓL�4	�"O�1!�==.��z�L��&���"O�8B�hYJ1�C��C�Y�a"O�k��i}��ߘ'�beQQ,<D�tr�E��uю`�$k�3�DcR%D��j2�_��l�hH��8�kso#D�4�]''�|�#5�T�M)�����6D���`g��r�S�$�_l8�5�6D�0��Q]Z�z�&����+��/D��q+��Ń�	��K�����0D�pz�	X!n���c�∏=E�1�Qa0D�8{��0t�[��B+��-AQ�9D�xi7G5��T��J�D�K��3D���5�,F[�t��
3	q �I��2D�t�̋�c�H�d{����ui/D���LS��F���W4L�v��R�7D��H%�QP �:�h�7F�Zm+U�4D�(H�E�4j#l1{`�S2�.�p�$2D���� �?%$��t�*̴d�u&;D�@S�T����+�d�$D��#�Fۦ-q�	#G�	��AC�,D�8��VX��"�/Q.ɤံ�)D�4��T�1�Px3�e���I�g,D��#UM���ir�F' �Ɖ��*D��K���+V��CJ�#�LEۂ�&4��zB� "U��͹�Y�M�`��ш�F�<i�υ`J�ss�؊.����F�<��AzY�v��#����(A�<y���>]�b�	��{�:�g�D2�O��s��ݒg�*���ꏚ)lsP�'����VE8e�O�k|n<j�~�c��BP �p��|�'���Y穝%��c�*O�a�1q��HO���4���.�5ɑ�٨JD�`V�'4���$����OU���2�l;}R�)��֎U)�K�dC���3(HB�	�^$P y�@�W�9Ue�� �@� �퉝3V̉�GH�h<+@��)�O"�DF�XFF�qDh�d�@T��0,�'�ўb?�BeG@�O!���q�Ҙi����6D���!��@O��ο7���062D������ZN"�0Ad�z��(��O1�O2�GD]ѕޓ*�b��Z#\���S�? ��3�@V:]��Q�f� �q�I�O|^HX	���cc��k͖8q
�'ň8z��.#�L@�CGU�s����	�'�0� RjM(_�\p0�LP�j��p��d)�'^@�`���Lo<x�s͐>k�׃G�<)ʋ�pN<�m0=g&ma�-QAX�,Ey�� FM�,lT��'J;n��[�'�LCuj� �n��4O
n�Jak�'m���ߑ
��x$&�ŦJ�'(~-#���~,�U�1 +#L��L>�شG�<%>%�6aZl6i2B��b�HD���=ʓ�hO�ӄ"B�h.�P5d���;v�C�	?*
�*�ЛaG���j���B��$����*϶��L�禝<L�j7�@���?�G��#^��ű�(��3�L%��^�'�?9�m��z�����Ǌ%$���u�-D�h(��ۿV�D�-=8��YzB�m�� KO��*��O?7�3%%�A�R�@H�J����Oў��'���<�i׺����`�Ԏ���*� ���:���<�|�'sx�H���#'o�P��`��F����'^�Ese�� ��xx�B@�a�4e��9B�%k�=��JF�}L�A�p)՟V�tt��x�r6tE�f��%�<y�,�pw�:D�Ȓ �	�5|J�Rc�_�s�f�1�G8�$'�S�'y�BD�%%�06�̃�	�	W/N1�ȓ<[�1�gU7���K��H�)�����6k���ǟ${��9`KA�Wb��
�')�PJ��ڢMY$��D	'���j�'�|�Pk�n�^��ǌD�����'}�q��Y�#(9�F%��}���X�'�x�C�a�wka{���i� ��ĭ<���i�2xz}���� ���!���9(����=�P�M��@b�E��S�Q���O����O(�b>)!'�4�6L1bd��q�B)-,O�<YfB�%6-�I+l�l��QH�Wy���	À}�v+�#X�9��7���O��=�|ڇ�!u��1���O7Dń�;��"�yrd�>[%��n��Gv� �D���h�ў�F{B:Odq� d�"ad8U�c��O@�!���'g1O×�������:ڜ �PJ1]*Q�|F{�'q'tkƥ��w��y�n�9=��]��M��(t�T�ҸG��SUf��Lb��mZ�&�Q�"~nڳƢ���3|E*�Z ƞ���B�I�q&��C���l��X0�ʫd�B�I*oN�i��F��!��aJ4f�OH➄s�S�7�Bf�M��.UbЈ�Uo'D����*�|��-߅�`aK$�	��Q�\$���/��4�T1��n��(F�1L!�hO���w��;�h�6G��M(�&S�W��7ͨ<Ɇ,C��p=bdƫ=Y�`�	h�tئVd��hO1�N�C�!�8Z�e{2BL6t�6�S��54������(]_<�Eǂ�~��n����d$^���`��rq찰�ȓ��rB��?/fP�&��J���"��]�H��`���ȟ@���1>�l�bG
�BN�RB�O��=E�d���t�30n�5e*����L:�y"������@�'�pDkjJ���$!�O^6�B�h�0$xv�]3E]��� (�a}½i�0�J��� �;0!;��\�)"�@��	X�'��1��A �m�T���ġ�*�'�\#%A�65�iz��H�v��'A��"ֻ���0��C	^������ɷ�~��)ڧDR\!��ޚ4|��ƴg"�ȓx삷��P��"�A�.H���D��3� �e0A�m�z�� (�<f�"OTQ*��hb��j��*�b���'Z�PFy��3W��x�jE+�6�C�F�yҭ��	�f��p�v$ڱ�A���Ŋ�(OQ>A B��/o��I@ ���p�|�&�*�O�ʓ[�I)�='�b	�G�����<��O��	AB�_�xĸ�#)!ΙD|�I����I'0��u�6cS�9O2B䉏d�:�V�_��p�`��=5B�	�0�!x��3
w&y9��ڰH8C�� ���9w�
�q�ajY*#�c�8E{����Z�B�*#�46� �۵��+�yB��"8$:uc�+v5@h����'��z��צ?�f<��H�'d���A�\���>�.O����Ӫ-�8�R���~� @��T}���~x�h��g�\�励��ExΨ	T(�O.�'.���Em�&]���Yf�!(|8u;	��hO�c$�
�*��-���
F��� 1O�=E�T,y���ӥ,�T'��!� �#��7�S�O�0xa`��ia
)��-(2�q9�'�(�a�aO.Z��i��1�M�)O�=E����o�, r�^	=��u��/A��x���+4]n���΀�2�Դ�"�j"?����Ej����Ï��y6%��J	!�D��1�(�3��+�9�R�\�󄄾=~qO�����xʁl��9|"lqG)��\D9��'.�'��xp��? N����Q��*�'cў�}���
�m��8!ᇁ66碔�t�Kg�2���<����"�'�17�u��V�z^B<`�"O|��G��AA�P�F�YT��!�i��#=E��4x��7�͙}���)�|؄ȓ[�xM�e�M�dɐyǨ z�"�I���?�	\��x`e�Ŕ_�^C�IBh�',��y�՟�)2�Jh��%�%�.j�n�0�x������I�/T��1pH�H"�i�O:d�� �IE>5Z�===�(�*��M�~08A+�>��F��BB�)N�����ţ'K�u��[�`ԢC[8eh7j�9���U�6D���Ҩ�'����"� �C�l�e�*�<����'o^��+�@��G��y�bی��ȓZ����чɻM��b��Q��Y�ȓO���Q��� 1�T�HF�_�i��B��Hg����̥0`oF�� �ȓ/ʈ9te����f�ƺF )��Q#>�ٷ��<!w��2���3��݇ȓ5?���V$�<���r��1
����\n�B�/64c�)qB�� (���M;w��� ������˂� 27I�a�<���Ѿ-P�@􂈿4��ٳ �R8��Ez��Z�������$t:�(3�Д�yr�\ �l<�R,�v6����߽�y�6.-ε�Q�T�kq\���M��y�ȅ�`i"���k�:AY��K�y�	K<�=yl�$>�\*��<�y� �FY���q���	Y�8�@LЕ�y��U��B��(L |�Zd����-�y�#�t
��MD�Hj����y�l<+pPŢq*_��D����y��b���\$0��Xr�b�4�yr��?v�e��%0pq�=��D&�y���`a}���<s�� ���y�
_!fc�}Q��I,m�
���eJ<�y"���'Ӿ<�1��o�I��H��y'��! ��T�>�X�	��y
� ��
�a��!�ԉ3q���"OH��e�5w�v��&b�:/���"O����֚$hKנ4G�\��q"O:(Ӓ�Q�,��,@0`HEgb0�!"OB0�$D�44��@�E�L
�"Oڅ:3�<M�����T��3�"O��j6�ϔNbR�y`N�<pGm��"O$!��cEv�1��n�.H>��q"O���T:=�)��l���*$"O���a�ˇ|�\AH#��-�y��"O����O�B�i	��G8Q��"O��b�R9�-e�� �j3��Rp"O�hӤ�_!Z�� {#!=(!����"O��0�/�S���/Ji^$z�"Ob�s�	εQ?�"Eϋ�7[:�u"OX�k���'?�h�w�A*<?a�R"ON��3��-.��Mpď�U3b|�"O�̳5`��[ ��2�5 Z���"O����c��jfd6M{�\:W�'{	K��Z%:L0�Sօ&_�t�pVC%vKH��X�)���3�'r�U����2Y���%��~�~� �'u�=Bc�O���1k"}V)�'f�=1v�ͧ�Q2AEU�z��'�B���
2}<0�B�GS= ��8�' >�@�ԚYO<@!W6A�F�S
�'/���"_#6�Z���;3P4�'��b�@\J�P8�0
.X^�q�'SDhq!�C#Zc2I�P�Je_�=��',^\Xs�G
*T�q9`��
X�(� �'��|"ʇ�OD�5���Q+Z�!��'�>���4
ˡJ���''��y��S��0)c�F$L{xU��L��y�ȍ�*���i�lF�B�^H��y[��D�%��	=p��˲�×�y��Φ�*H���%>�~9���1�y�D�aR����A�Ny�i�qĒ�y�*D�"�`#�͖?��y��ڊ�y�ȓ�VGX�چ��c_HHk�L�:�y"ʓ�z�`�ئ�шR}�p�D���y��K2m�ƙpƈ^U碼���=�yR�DJD9R@��7@N����A<�y2Ü/���A�,U7To&ђ��|�<���I)1r颓D&w��ݘe\c�<�S��:1��@��E�Pi���'+�{�<Ɇ��	�jE*��	] 	0#��v�<s荬|�����0ҔY�F��p�<�unUOd��~���AT�<!����~��iD Sz9�,kR��V8��J��Ms��$�l2W�^�$�HԨ�"%^J��e)�O�$�D�=1^�k��
�⠹
עЩ$"�+OX����
@���L�"|2T�Y�a�بքB�*r1�K�'���3�o��kL��V�"������sr��#�L�á�)C
�C�R��Ba�F�3�ɈT�,���:J,���B�� �	0nX����8?��S�'	'^1�\8 3����Dz�i��G8�����"�0v���[�k���
��]�b��(�e�9�B��'��a�`J$uT��^$6�k�L��P�(O|�0��O�uY��+�Hi�R��<�O
�IŎ�v2hӊL�Z��baڬ{Y�A̓��y� E�(���W�_*��)�'b�N�g��kqQ*��Z��E|bl(<���Na�'P��M�v%�.c�4:���4�@P��XDy�H��ʔS��{�	 B!3�f�;��b��ٽ�y��3Vb���S�O`��)�&W|D����C ~��e�*e%ߦ
��H D�'�Oƙ�CL%IKh\Q@.N�M>�4j���ؐ��]�h�A�6Oj��D�I�*
��9Q��<����5[�S7��QS�xSqcZ��0?�a�@�rӶ�r���;7A�ԫD��)}�2��GG��4�H�	%S�D��ũ�=;��S�π vy�1��* cb�{����I.m0�XsPC�fq�Bp�b����Tg���S�ʐ� dDw�ɹR�Θ� ��|�ݩ39���_��c����y���Y��Y�A�z���%R>H�E�6�(�3UWY4����I���:{�V|���U��'�����<?����Uk�m����d������P�$���[5� ����k��@~�8Ha� =
f�u�'a���I{��æ�«��i*�'Q�>ѱ"ʠi�G�8_1�ȅȓH��܂0ω2=	�=��-߻Spfp�d�,	����m�ԅ�Cc;�3��W5�\u4�Ҕc2�XBN_8����a�8|h�'�,'߈YFR�r6�|��B�s�B�ͨ����I�m��AboH4��I�z5��Dsb�F�?�f����8pHS�ε$����*q�2����Ɵ+ښ��`L�;o5�B�1o�����,KHUdG�%���F��(c|D<��dԇGy�1���0��$%�;<찢r��|��Irw
|�� ���E�J�z
`;bE�����cB���\��Ȑ��F�"T��q0�� ���5�x�@V�x@Pjq�
D�c�fϊ^fP��Ѕ�5�p=��b�Q� \q�ٸC,%@@�]T*8��$�1c>�b&$�� mŘ�%²��dȂ �8�����']�} ���72,�j��$s�b�"�{��R�s�R��r��]���Q���7(�{[?��F�7M�
h9l��#���Ϟ�yo2t�-��! ��!�'�܁qs/��b�1q��&^��"�K�1����kCvyz��� ���]�̈�'���j'������"�1QLNL��O!Z.B�	7N*@b��*o,x��d�&S0x���" �6�� 9L��@b��6L)D0"RH�O"l��DJ'Q4p��B� �hԯ0�l��Ђ\.��@��t(�p���.3X�I۴KB����Y��L����N�򵁤�JU�Vu���L�]or���Z�g�Skj�	�.��-+��>3��➐B��_�KW��j�h�Oil����w�rl�u �(Qv(�@���(��02�kFX�!�Rrx�ܙ:u�d���)Ki�>����[u*��4X����i�X��e��)
��ܫ�V�	l�7fI>N�8\y�
4rF����,$�(��g�$~.I�a��(2p�M���͢Yzp6�O%H?n�0%ϻ,?$�1�KΌL4�D���M��;+�!c�ϊ�L�4m�gR"l%L1c
�'�fy��E\
4e<|$��cԴ̉���OUԝ8��6Cq���˞�����6`4t$',�Ć�wQ��w�[�9\�|��هGa{"ǋ�l�L)�`�ȍk�xS��H��q.�+GNmQ�kئ3����d��)솘J�`�հ<�g��{��T�";��$;0�zܓft�H�'\=Oy�ճ�&�j�����V~�݋��]� �úbXR� /��S����	��?���V�6���X��ۃYUj(Yș0�x���L�t��-�%�b��MYO�82���@��?1�rf�uVN�����0a]�Xr��3�23����;!ŊiQ0�I��ħ@�J�fe��B
���p�V(J�F�X�qf�E�Nf�%m��m	[w���r��&0����M<Y��+rh.���kN�|e,�sTg�Zy"fF�=3���O�]��Oqx�{����?<�$�V�խ*q���P/�'G�>l"�&	�:�̚�I��U:DC�Pi����	�@�vE(ǎ 1^���W�١v�^�L��#����F�*��ȟ/
�� ��\;�j!�6���҆�$A_�ܙ���|���2E���?�pD��O��8���
) H(�.CV�x� ��z��r`�Q�8`Y���)ʐ��'��!2��.^�[t�L�A3��`gY�Aџp�w.�.4����D���Ƥ[��Og��p.��C!i��tO�L(� �\D��'�ΰs�$O�'�E�7��� �RԣUf=-4R��)O${��כ���XI������p!bGq���˧�.�4)��I�1m��lQ�'�?ot��p͒�n�z	Ö�'��!�>�Ơ9	�m���j>}b�UC8�0S�U=-�q@�6@La$��5�Z��;bi(��E
OϘ���(��q�A���bkK6�9؆�X9`�X��ϐ"uo��n���0��o��P��6���|���4�����F�����p<�&ܖ
@b��p
�X���ɑ¿��q("��
�:d��ݜ�4Ի��!��'ur�ON-���T ��Cb6�9�\��������LW&L2PLf��p��_�D�h��ZLZHc��ر��5�	T�]�mD}�䅵$��0�i�\��p �	��,��6@� ԏE���'M�����X4 >}�w�<��3i�JA�-S��N:���I��DQ�3��e��R��(�̭xP� �ݒ��$I-,S����\��pH�M�@Hd�I�ߐ�?1��E�`:�������T�F9�G�MH,Z#[�S�-�9B�
e��~}BhH�XΑ�6��
K����(�yBdS�T�h0�p!�!B�8��R/�y�(�	*(��s:��$3}"��ħ#Җ�P��0A����N 0 D����Wt�=@"��h˂� A1%�J ��nF
2͹u��>E�Op��k'�3}b'>q%���śa��HA����O��Y2GO9z�D���	<� |`�5R���J��"�ܱa�lǇU=�hsukOhX�l�e��_8���	��EӨ�d�Y�^P�a�%#�	
��S�4�ąJ��6Pg}r�H�h0�"X�{y^
�����y��8x�^��s%ɇs�T��ӽ�y"���:P�`���4$$�;�&}��ħ&��-��3a�����A������,`�qZ�i��bJ^y�I6�� Y�6uᇤ��C$��O�e¢�?�玑e�1Oh C)�>Q��f�.4립Q2�ɒ 6�)�����}C��D#�LKF�\�M*� n��F��QtB�5f��Q%����(Y2\��D� GB )ҕL�F���R�A����]�.�A"F�M�	h���G`�խ�%`��D D���H�A!��D\PJ����b_�_�~Ĩ��B  m����T@ Q�/�k�=�Wń�c�@%���Q�ʈ�F��WN����L>,ЁEаdLF��K���Q�L�ЩPN40�A�ѳaKL�2��M��
)�;Os��(g'V�cİ"Gn�b ��ȓg����ЪvW-��M�Q�4r���y��B�С��1E.��b���7�9�4�!5IM%1�����	Ѿ"�D�c�"O�U�!�Y�?���ԍ�i�f���D����s��(N���闪H�4��<���>1�)��<�|����R���i �v��tuh��hx�)�u���GW�5 @ +�`EX�$�	'JO 3y`� �B�3Pa{b��xX�����͟ZsR$�⢃���'ZVh�CY.��[%+Aڪ��b��v��1��ʇ2Up�x��	&x��1"O��b�Mr�Mc�fLF�j�k	*c����Q�\4Dm���T��"���"�͎L�'�y7G�3(Э3�ӊ+�Н��KQ�y2(S0�+����J��N(z�~�4��'Fd�Q�@L�0"쌲����dZ$&����'�jܘ4�ҳK�F���k�1̄ +
ߓN�J�Hc	�!�n6��1Af��@+�'���.{?,��'2VD�Ŧ�C��{��"C�Vx����$G&�Y5ၤ��'�"(���"G���'�� �|��/X� ��eU>�$ّ��]o�<ɥ���/R��[AD�]��]+\x�|�r%�>��S��y)T����s	��<X&� סė�y�S�6���	��E*0vPMA�����~b��(D.V���I!D+�%`s��n�8�5bN&D�B䉎����1��b,����'�,B䉝#��\�}	bbѼL�������>�h����H�$�ru�?=:ء�発[@ᘵ"O��� S�; �����(1rX+��>�SÀ�Rg ����xP��	�|E�7��O�~��C��X�/C�9�J��H?K��m�.KU�<i�l��{��yh;9�Fd���O�'�h�g�OZ�OZd���e!�ļzw��i�TU[	�'�䜳r�~�0�qv��>H�E��'�~��&�Os�S�O������
ex"d�u�RYJ�	�'C�1��Z<��rS�C)}�\���!}��Q�t��I:Y>���%} � �̦!<��dD�v!�|���ö"��` �f�&��c�<�n��gX����@ l��H��X�<YB�T�D|�
R��h
�(�m�<���T�d�
`��Y�����,FA�<����c��)BӆBw��3P��~�<�f��6�u(@Κ �,�م��x�<7�	����"PIg�A�݄�y"KH�z`�����XR����>�yb$��I�� �ݓZ��q��~�<�a�)Ci� ɑ[%k�����"�y�<�%(Չ?,%���.:��#�͗z�<9"���B�]x!���_�֙����C�<��L�
;Ph���G	d�0��}�<QPT�1&d��F��1y���Do�x�<�֮\:5���4� d����ƐB�<1�)J0 A�y+s'�L��e*���T�<��	���E�SO.QFIK4��S�<�oU�0�9�P�{�@g Q�<���Լk<��e鍓�P\2�g�g�<)`��/d��e�|�xġ�Z[�<� ��& �,v�$dKGeփxc��9W"Op%ـ���F@3T�	<S$� �"OR�����:�tE��ą�h]*T��"O�a���IX�t��,5��J"O �*5�RH��1yrߴ=E!0"O�����?�<աҤ�7* �ba"O@c,:0�ᘖ,U,~�ܵ��"OQ�T�ql�X� �8�V���"ObM��*��n��ɷ`�M�b��"Ott���o@��q$ډceN-х"O����i<H9<	X�M�M���b�"O�D@'O�	Y@� �o]�x�@XP�"O@�Q���'F����65��4� "O2�z!�� �g�0�TmZ5"O�D@�J[Z��	2V�Y�RD�A"O�	Bu�9%�฀�M+A~��"O`e������bB���}x���'"O$�3�ؾd~����X�!{"iR�"O���Q��$"���e@,P���"O��S֫�&(2R`I�".i!5"O���L$&.�s�/�*l�DA�"O��h��O��5;f��.V�4"OjY@R�"�~eZ�!I�e@�"O����׸3�|;a&F�+�"O"���$V&:K���g$� �M��"Op�S� �:��p���	�����"ON @�*V�)"�䱇�®BHf���"OzU�WL�{>�����C'j "���"O�I@�#�$M"M	"F]'G9(�"Ox�*�AJ!w�!��,��6��"O����L�%�D8!��+��m0�"OF`Br�R/���H�{��+$"O8H���#9�x�PQ�13�5xD"OzQQvyr�Y e��J����"O60��Ƈ��ೄԝ9�dI�"O6���`�_5��� bI�\��0�"OP`R��.*��C���3���C"O��C�EU���J����(�9U"OR��)ޑd���"[ƴ�"O�i�t@Ǵ�����R�]x��"OF�f���Z�Z@��H��x`IIS"O��P�a�>24��FM+ �KΧ�y��;z�~����c��嘊�yB��I�E[��XPRM���y�e�	�p�j�mO�%_�̡3�֐�y�W6C���	£�N��#²�y�$>��I�M�&��EX�		��y��&?�TY%#E5c�I ���yRH�?FK&i�.	'N�a�ʊ�y�aJ�D�&�T�H�M�p�˽�y���g�6Ec�n�z ������y�p޶bM	3O�0+0Ǚ�p<�&��4$�44yJ<��&zt�qWĞ/������Lt؟��&+M�X@�')Z;0|X}
e��s$rq �X��q��Ԍm�ā�Ց>E��/�J�0,��Dd��1�c�'��O�X�D��#\Hb?q۵�6g�n]�D��R����a��6_92˓J�@u�6&F��g��Z�`H�@%f8JQ6$�l$ϓf�\3$�"'ҧ�O�x�*�B%�׫{z��2�-Yް� ���s�a~��M6J*,�V�?��zf�A�����v2�YuĂ�ybɀ� �6ܐ�gW��	%�,P���44���Q槃-Dľ�����`Xhp��C<O>RaS��і��u/��j{L���3O(���]�z �懤<E�����b�!ʞ���;1-�XE��G|�e�*t�ccSܧz�Uy6ei��+S� Y�d��'��Uy�|����{�ï-��$��6^���"fnM��yr��3d��X�5�Nn����.��� �M��LЈ/�� �J���<��Z�i���r�'F^��tD�
O��k5F��J���O�ثw�My��y�'��\0!AI<y��`��Y�P��l���qv/Ưtu\h��{��<i�\�`�,�"t���$bV90�.$���#(���%���1$�I��)§w������D�D�j���\k�8G|�nؘ[>h(B�Hh�':D4e���N{S�@��"�Xm~��S�|�b^Yoz��}&�$�ED+~3��"-��F�~���n���g�@+�.�x$�>E��e�<z��Pr���p��q�ݨ�yBV;g����H6ɞ�Z�f	��ɑm:�)s�"�J��ִ"�p8C��%?�%o�5����4��&j] �_؟���^.��d!�)�j�(M�s�����>q�J
⺕;�OHZ��F �>E�Yt#��f>�h��|���@ܟA��0Ŝ����'@��rW~��S��|���G�,��|��[ⴼ��s1ҳA8F�0�aE��}=���i!8`�3�S��>����-i��+�g��e� �X���i���4(�E��[�$�&΃ǔ)��(�~�.�3G8�dh��M�cD��7K�b�<-�P,���=j>��OF	7G2Uh���c��ի�c��z��DF?>a��w�,ѵ�@N�đ�c_'E�.P0�'��Q���,b�d���j_;�\�" (7{Yj���-/���ND)��Y���6ғ6�ы�햝<N��Gh�vG҉��	�j��9
 �\�p���2$�,�:�� L���馯űI����*�L��	4ܢ0�/.�R��C�0�OP��0��a@Tl� �B ef:���ž;t�G�y�B�!N}���C�ʀj���P����С��9�0i�B��P5I^f�°
#��]IP�����w���U�0�����!q{PB�I�-��@qŀ�kB���gE�#Q'����&[�چD�}V�0U"Q�,��">񇩓��>X�������B%�{��`@�e�)B:�x��N���9���	M�I��ǟ2�H,�6D���ҏT�1�tZC��NX6�7�	'-�X]#�뇖}���E��O�8,�j,�cD9d� L�cH���y2"��P��̸\���F¯Id�5[qbK��_��3�v9��'6?�����6�"=��i�[���"f\c�<��ÐVA��JRmE:!F��j�ț|�8 m��^K��@7��2Y��i����O��{ת��1��ǯ]�*�k@�,D���cˢk
�x�ފ)¨A"�ޮ;��,���Q�5����&��)K��HOHq3��6���1�E1=��H9��'5b���*���nڠ0;�4Zu��0� ����eNJ)ӃˡP��I*#�'C\@aMG�+O��2�揻{E�	ʉ{��]� ��Hb�	�M��d	(f䘓'� ��d�^)[H�-�!M���|It0�xr�^�Y��t[���M�<:��1n��`�M�B\�i�hȳ��.W��ن*����dK�#��`�4����{?8�²�Օ��O��� �Ҋ����H|� ��5]d����<Fqʱ��	��8�J#E.*z��s�47��Xwr���KWU��`���m<GȠ+�,-e.��'�`#�]�(��)�O�d���bUp I�0u�3��$���(W��;!\� S����G&���7	O���=��e�z��8���3E�2|�jR�-_�f�rE�R��$HT��O?2iYvhV�,�NE��O���3�g��W�줢�.F?h@!h��G���S�e'/���鐆��6�րP�'	$5TRE�2	�n�R��M�p�t"��S$4Q^Y�R�H�vĀ�W��S��� �	���O�U(��^�ae,�>�ȅ� P����'@T'.p���!-]�H*�Bu��-{Tm�r�O�̕�Ԣ�a�V��:��O?(k��9FD�/b���'����7綀�O�ɘ5㴔��&T�z�����)7=��Րu&�:H�}���x��@�s�]\`x��I�PE�cC��!~��[�I�;�, M��;��Zap�``�ɂ`�$i�B�w$�A�'Z���n��1=��0�m� 1��F;sU!�D�38���I�T�Y���#W������c�l�Q��3�l%"��I�� �)VQ�O�jԐ����4u:Q@QfRYd��'���dAY̓���h\s�U�3*��,�ԁ�*O�#���7��;�֑�BϝH��C<�I�M�V�����]����L�B�7Ϙ����5�0_ ipd�>�H�VƅE].hX��E0)B�Y��(DjwdTH��ըOX�r$�j�@6�YJ,hI X����	��ȀR�4x���D�)b<�z2��kĆx�O��.��uY��	f�؀FO&1_���t&�=^�����<��Bc�\�d���-�/'�&�s�� 66f|�e
����64bt���-�xq4E*���*���I�kK#n��9ѷR�aNӧ�	ұ'�X�����
���ʛ ��Ey�a�$D�dD��g��N!�� �Dhu�O|r���'@�+l��
1O� ����:v��b&���L�O�`Q�~2����#줝��	�:������h�	�h#�z��Y.O\du�',�;ܠ���eW��Ւd����I.. <L��O���ƀ���z݃/��l�0"B�&AC�]�1���U+>9hrɏ#c��ɢbP7���*��1$��J��_�(�a}�m��=�7-Y]����!h��9�XW��P�T>���l�-Xu��8S�l���K-`��a�@n�7.�p��4D�$A�A�+1N �
��Ҍ��ಱs�����*�"���,S<5QI�L�Q0���ܨW&��2��K�lD�"À6�p>�1�ˍ�Լ3ߴA�@�&��W� ��G蓤T�|!�!K�_i�I��5��Oiv�i�H�I�O�:�3�b_�]2��cb�fkd�Fz2'w��F����t�� 
k�?n�H��3�x�hg
�Q�����.�<��'�񟐠�r��^�hْ"Q�pd��#��'[��X�n\Y~b�V,C�>AqG �XG�q�E!�n�"�����?�U��49T�9J~�=�����F� ���@\`��.�v��`���!v@4�6�D`d���{Y�e���"m��d`T����=Q� Su��yF�4����N�'���@1���Qr���E�6��3rM�����+`�\ŀ�E
�_��g,��qO!�. `d1q�,� 5�t����[���"R�VE�h 3��/t�@��%�,$fl9�~λh����cO�QES�B)3"�ȓE�TQ�&��SOL�D+�T4hr$
T�l���!��C�1(��W�?U�v�PH�O�u��iL#] l�&e��`���'u�O��~)�m�7)ʇG�$��R�V
�9aO���T84�ҍ+)p����Z؞�b ���#ai���o��1�T$.���D���� ��}B�,�CW�ي��鉝Y��c��H���A�{�p�@FZ9g!�<F���7ɏF��p�F�1P��3T�޻~���@4)�%m<�Q��>B���}��w��� �ud T"�k˂3���c�'sD|�aO�0&���iզ��;q:���D&��9+r/Uh���3����1�2 ��c�����/�j�P�.����`2|O6�	�,���4C����n^:KȞ�)�`2��0Γ+��l	��=a�Sq�ɵ �[*��W��T���ٲ萾(��ʓ�T�맧k>ţ��G;J�)���M�(U�ơ&D��sd���r.�`Y#��m�I�;FVM�bHV�)��<�g�˖"8�p�'��&j�qGf�<Ѷ�J�^M�= ��F��nH��Řb?a"��,4����QaP��2��۰��VCԱ.�!��X���	�K�	f�Y(�c�.c!�d�Y���p����2d�±�:'!�D�-J�t)��[(.������?!�D�9�%�7L��y1�#��Py�).th`�g��}Cũ ��yrm�$h��{���a�		�y��E!U�\4��@@/_�XsG`]�y��^/VlY�7�DP�D������y֤[7�<y�&N)Q���Ch��y��E�O(�i)�D��9��u������y�;�A@��!�*��+���yb�
�4B
؃w��ܰ]���ֹ�y�#��_���g+��&i�5.֮�yr$U*A�Fi�V���s���Z��Ѥ�yr�W�鰰G�,h���cEƐ�yb�\�}0�1�!�T�r1	����y"BL�m&}Z���,L߰!�+R�yr��0U�H3�'I�B@�$�p���y���bU�t&��C~ �PgƵ�y���>Uj�+�m�*���`�y���
��uM�5�N9�GK�.�y2�2cp�zUiQ����ѤB���y�DN@-��J�e���D�(�y"�M6Z�00M3f� ���k]��y��I�ojZI"Rm�]�z�/�y���Io֝A�焏][��� ��yr��4@\:���R���$�(�y�mX-Yޮez���	T�Xa�Ê:�y
� ~\5��}��X�阈W��i��"OZU�A�}6҅A�A�2H��%s�"Ob�K6�B|z�H7��(�"O޹�Kh�> bTg�uE(E�A"Of��'��b�s�&U�]0� "O����ZwP���(�T���2�"Od)��d̃Q&��0EN@��݁�"O��Ҕ��?w?X�+�e2��X��"O�<��+!�`����+1�R�E"Oz��A��W��������;�"O<MJ�C_�\w��3c�^�d�X�� "O��pŅY	���cw�ō2�i�"O��0B��:o��S'B?p�V@91"O���	�|��c�f��*x��5"O� h2c^���8�&<VP��"O����B���7b��
�xA�"O�(�fװ�6���bç-�v�(�"O���s�:{�jz�A�$i�&�а"O��0��r��`s�J�a�d@�"OvX��]=6�=öb7o*�$�"Op���gF�BN EzE`�-�r�"OLYF씧7|�y!�%�%!�"O��S�?�8]a��5`�1	A"OJ���Ԍk�6lZ�"��%j�� �"OQ񐁉3ʔ�V@�DO(��"O�"�&�׸5���޻�L��"O�`�,ʆ������Y� ���Aw�'�f�lуD_Θ���aZ�(V⋝l�Z�S���:JRԸ3E��
�y�������4eͻ��9O1�L�a���/�m{f`_�5�"-Ҥ��0���>JjAR�i1�Tm���V> �z�6L��6=#�9Ol�ɩ`������"~*q�@9����F���P���� ��`�SJH/o��'.H"|j���uW@�8<�0R�ŭS�xi�f�ˣ(�����a�d���bv���GG�M�2���l���� �O�a���!1��N|��j�
%�qP�*P� ��"L�F�.�����O������#[p�e3��%=����H�x�v�e����<�2)�5H� 2�>U����,F�I�U���?�}���a�$� ���Kf���Iy�@�w��OQ>W0 @a�v��X䊵bc�&d# T&k��OQ?���a�7 �[�X�.�dr�LC��d�=a��O���Q��پJ�͓��7�`�?I�@��ħ�8$����_2Q���]�Ά�%�`�4�;�S�2h�R�aV,_W>��R�^��4a�'�`�������SU�]��r@b�6���P���O~�O��ԧ�� x�F]V$��B&B��5Obʓm!��	W�g}�O� �04��'#� �F�J$��r�)�T�S..�Є����?5�z�����䓵hOq���*P@ .�i��%[%$��:�R���A_W�S�O�p�1Am��^���c])]HH�
��Դ��b�:ڧ<�~�JP$H�H�@�p��y���C��l�����(ҧ?�D���[�?�y$F§E
����oT^�'E�̧L��G���ğH^�(�4�y]Z� W�<*N����ȢIRM�ǅ��r4j�S�OV� k���	�:�!F�
m�Q[cEL2FZ]���S�b�|�S��?��f@"z#���G*K�����p�<�Q�	���UC��&(D�bE�D�<a��O}�^<Yw�ןfθi��E
B�<ɢ 3���@�(�c��|���{�<�m�h���P�M��sl�C^Q�<�ψ<UnT��C.<f^���t�<�%���+&6���*&�4��4��d�<��-�8Ӟ��4�#7��͒')d�<AËկZMF��3���%�>8���v�<A*�8yR����Q�:�Nuz���u�<IuLPBȰ��F��<+$���Gr�<�"��.}�Ԭ�׫�1�h苄�Wb�<� �8�1g�1����A��&�&I�R"O��YaAC�Vb�]��&Y��IH�"O&A�W��0�$萭�@�:ճu"O�M�@a.��UZ�k���<թs"ONA���Ĺ�T����t�؀��"O��#���qj�'"��pq7"O��Q��/'k�U��#gz�"O����߃Jzh��'��dY��
"O� ���բ��L�G�6-S��"O�ę�j�#}���K��C�"s"O"<���C����ň���2�"O��ҡ�F:,�����։+��	�"O����qFƉ����,t�8=r�"OF5@R	��~CL4"7��/�<-0"O�i
�O�c���,�/�PB"O��. P���a5��*��=A!*O"��ꕗ_��`�E�� g� ��'�&л��Ea
X*����f�hxi�'Y�!�*d�>�x��J�(��	�'���&�D��Y+5��� �h�Q�'��]�wI  ��YA1�_� V.y
�'�8T"��W���3�˱Dغ܁�'��
�\?H�0*�n_�ml��	�'��c��n��hځŇ	b�q��'oj	����Z ����[��	��'� �-�8�Y�@@9
�l�
�'X ��#�)�hأa�~��u�
�'s�剑�_�gt�;P�q_�B
�'�"��1��N��7O ^�J��
�'[N���l�(Ȏ � ��V���
�'�mI��Ud�RgE�"�΄#�'�(Q���5X��AH�i6jM��'�p�3@�K�R�Pp��ۦ!��	�'I<1��DJ�e>�8�gn��x	��b	�'�(!s��
���c�E��Z�С	�'FP�J��U�&l��/��Zɐy�';�����8x�� ��T"�'���Y�ԓ.� �1��b8��'�Me�َD�x��J�~Rz�
�'�4�Y��ot�! 
R�H�p�	�'R���t�^�T����� s��h��'"���-Hh��{�B�o\�-b�'�]�LU��,�𨗇�BdJ�'[��ƣ��I��aKP̉�{b���'��5x�n_/���o�� ��k�'���Z�L�	c��'m�&f/X�'�d���c�&.z!J�#�#cP.i�'�~�I$ᛓc�4�X��]�d���'Ǆ��"` �_�Uz�k��XP��'�- � ��F�>�{c�ǛI�@��'�:���|����;}xHs	�'�d�A�O^�|��L�f?xZ��'0��w�?+���'�ɶn*����'�ɹw��.�,t�@M/c��j�'$(w-�
Dkj�7��9q�`��'̵1S��|-b�(v%�%fb��s�'  5�f�˵Gj4dv�C�Sv��'^ژ0J�	���g�u�����'k��R�\%8��0i�K�g\0�k�'�rx���]K N�SF��b�Pt3�'l����K>d̲���'��*� �':���eR�Kq�]
F�޵1̜�"�'/�@�F&�i}pBe)�%�P8�
�'�d4��W	?BɄ���/n��	��� ����5(��"Jə-A���0"O����6�E�W#�6NP5!"Or�r�J���2��B�p ���"OV�B���b�%X�ы7"O���BFT�.��"��$MW,Eb"Ov��DݾS��B�C�*>"��"OƱ��I,��c���
H�`k�"O��8��O;{v �c[
p�V�"O�S"�U�d�jw лC����C"O�ݳA�R�E�@J�Oىq�́��"OE*s��3�b� ��&U�L�Q�"Oha��d�@/�|K@�u��T��"O�e
��,Y�Pȳ�T�T��p��"O�)�2K�de��œ+�",a�"O ��Òt3�̸pD��z�ҁ�r"O�ђ�o�0.���a4C&N�,�"O�"	�i��sa�KhG�"�"O���^E��T����6A�U�"O�	��+ /�4q �Xϖ���"O֠i�E9\���ÐY�\a�r"On!2��7}b�*�"A#)�Ⱥ�"OtY��'�7�8�砕�Dܐ�c"O�ejb+]<���)q�ޙ|�4dp"O�T��bސ}JTM��L37�l�6"O�8���ޕu�^�B
K1%y�Q"O�� w!�,�\P��	�A�c!"O��3c��EB��Jfh6L@��"O��B��ӋB�:ePN�-��i�"OZ	���C�1r�o�� � Pѡ"O��BSiY8��؉���k�݂�"O(4[e�Tb���"q�(o;:�Z"OdTba�W
m�xɆ.��k�
"Oa�@��u~(y�L��Iin�@�"O���,˂'�P�K�+�
 h� "O���4�ؓ
�V-ȣE�20I[�"O���g�/0g�!*�F�%z,0�"OdQ9�(�%iO�4A�%�\,$���"Oi���x���%N�y�>��"Of�2EEf/v�3/�*vѼ��!"O@E��n8v�0i��U){��B�"Ot�&�ȸ\7�	�GDդa� �[�"O�U �`A2/�ШX�IY(�ٷ"OJy�/.1�wƔ 3>���p"OJ]k�A��Gݜ	�RŃ�=���"O��PװP�����(^�\a!��HU�
02���A�"q!�D�$�j9P���/q�TZ�MZc!�[6d6��[�o��Vh8�"��i�!��08H@W`�gx�XPi�xB!�W�$�x �C�\W&���h��'!�^bB6tr�F}L�)1��6N#!�d�H�yB�Y-~� �%N�T�!�dҨD,JT"'L�!d"��\;l�!��U�f�r6=�����S�!�ă�c'�����Q�P�@qƒG�!�D�U�F�J�mF!�x!Jg��7b�!�$�I��I�����=����Ǡuf!���3�^�0��Y_"��
U�>X!���3Ě8SĖ�U�� �g�yF!�d�:l�P�GB��\�q�EMH�,7!��K�k���	'%�
�2�Pt�BU+!�$�5<*�]���Fp� ����+&�!�dZ�7��٢�D�� 8�Q��u�!�d�<2�X�3���9�]�PL��!�� 6�sd��8L�ѓ����f�nd�U"OZ "��/zFT��l�[�d��"O ���.<����wK�b�����"O��fO�NV�)Jd���o�P� P"O*$��&\�J�y�ea�-u��)"OL���G�ZS��@�`� }�>Ԓ�"OP�b�ѓM`p�"o$�,iye"OZ|"a:#,L�b ��P|9�"Ol��f���N�%
`O\ iV����"ORY�C�3�����-�_*"eHQ"O^�Ү�xi�ϓ@Z�ӂ"O6i�4�̿���Zl�B�&�`&"OTLX"d�^U����v��A "O�=d��(�MX�Ҏ��p"O��1�.$J�Җa�2T�Թb�"Oz�XP��zȑ@�(&��MI"Ol��tC��g)F�����x�R�x�"OYP�/'��9�Ҍ|}T z�"O �y�L�C��(�Ȕn\X��"O�aI$D�N�LZg@	M6d1#�"O�<x�n�*�!��VL58�"Or�bA��%}�r)2�3h�C"O��q��n��R�IƐ;ԑ�!"O,,�-�#m��E���.,��[�"O�����G�D�l�:S��%Լ��w"O�Ypa��g�T9�q.Φ>]$E��"O�A�D(�2�&�z�앳U��ɛ�"O��K֌L[^`r�e����b"O�����̓ C<x�E�lJ�Y�"O�89��Q+�B���E4>�h+&"O.e�7gè8����]�)0.��e"O�2W��	J}�m2D��I.�,��"O��ƨZ�?�d�{�*J�9($!H'"O����J+������)ƽPT"O��a�!�8j�\���E����6"O"�@��Wft��ʞCՃd"Ol��v��2s<��{V���;@�y�"ON `s��/V���7�n��dQQ"O� 	���:J���'�օZÞx
5"O<���#Z��
'��^�ma%"O�`)G+ 丽 aJ�)+Qxqa"O���$_�SĠ��u�9���z"O ����E�p�9� I��jʀ<z!"O�|S�U�K���s
�����&"O6P2a��Z���JC�̖Q�hu��"OnX�c&�(�|��-H�H��X�"O���+�Rұ��0?�ZY�e"O�$xQ���sNe
�ǃki����"O"@0c�ךb\���K�'	h�\�"OdD@7N@0nk���HB�T 1�Q"O0];�%�0������3\6����"Od��ҫ�
/)��`%~�hyQ"O�D�s�<���ĉW�w����"O>�JӞ8�x����V68�B��"OxUkPeɍZ��0�gG��zKX��3"O2�(��k
y��F�=[���V"O�}ʦ   ��   �  P  �!  �,  �6  EA  M  4X  �^  Uh  �n  �u  [�  ��  ߌ  &�  h�  ��  �  Z�  ��  ܸ  �  b�  ��  ��  *�  m�  ��  ��  4�  w�  ��  ~ �
 7 � � V$ �+ �3 2: t@ �F �M ?T Z �` i  `� u�	����ZvIC�'ln\�0BHz+��D��g�2T���OĴ	g���?YV̒'�?��]O+�)Hu�t�ԤR�
�cw:17�D�MլY!�l������ք�C�N�",���)U�_���)\�<K�U�$�J�Y"�1%@�"<�DL�@ES�e��ۦ���y�>�:�BѦ^:(��;)�X�B��F�����+�N]j�
��,%�YCP
ݣY��0��/�T�4�dM�{Zp�a�ӌ6|%l��N����	ɟ��I��Ɋs��KS�C2o��z����<�b���K�����4Cm�F�'E�t�O��Id�O���'��5w�;R��"e�L,����'��FeӪ�$�O�|��a�O Y�v���|HR�Ŧ�u7�)gg��W��Q�-A��!�șZ�O��'�z����c��Fɶ0^�T��=-���m�>��'Z�'K����T�����4��%X|�A!@K �zf�U��?a���?���?����?�����|�%3fٯ.�eä��f�8�3��O��n+�MC��i<�7M�O��nZ�h��pߴC�N�і�[\X��D7Dj��3L._��4��Q���l�������=-N�韔�)7E@����UW%�B��C-P���q�߲~J�sJ۟4�4| ���O^�������;
z���;j�Q��N�+p&�oZ*0�x�aG�J��Ih�
Ξw����"�v��ȩ�4}l�6�}�Z���s��!�,&,Bs��S� ɹ�Ӝ*<jum�"�M��i��� PK���`1Fћ[�z� ��W
� �$H�++��15�A�`n�	z%./N�2�2(hӶ0l�!�MӇ�K$e�h� �ЪEj���+I�D=����8
�B����e�i[�xU���E�X�;#A�X�n���'��O� HO�'��E �$#?����O������xID�7�M�ϟ��q�y��8��]�lT�ї�'p�	��T�	�|R��0N�r�.�b3�Φ�Q΃[�xj5&^�,V������7�ް!�~�I3�� K` �	�9��e�ro�!��)W�r(���[�+���')�	���Bݢ2�j�z�a]0CI��	쟌�Ie���?����?�'HA��l��h�֙��J� .B:Xj�)�&��l�Q(�@��lY��	��Y�\6M�<�̀@Q�V�'f�t�D�'g�,2�D�(I�Z<K�,5)�J�QR�'*�菩S��&'�# �8��H��9�ZQ,�ug�)[^
a�Ó��:��dD�#�L9��SG�lը��"ڧ.�^��E��%�t�Z���S����'Nf���W���&ҧ����B5=�<5��M��Q��Ȩ�����?���?���i�3
(�#���I��mY�<x�џ�{�4-ț��I��D��J��ҙ"�ɀe�L��7��O�˓Vn|-����?���?�-O`�"�Q43� P� @4q��ٛWB0"���R���ئ��R�U�+�"�?Y���>@zY�
2:�죆Q��m{w���n�`АB�N:\8�|2Q�f~B�B	��QJq(Ϲ0?(�����W�&H�<�q��ޟ���B�L>���Eyw�|QA�& Y5��k;�?������O��?��'�0���֞��&M±4��+O @l�Ms����U>�e�tI�D��1��b�sA�H��K� W�u�t�>���?1*OF�'���θE���cD�=�A�B��y���+3�ֿq.���Q���y"K��GP��KP�01X�j��@�Z�R�03�XТC�0l}q'�E���Of� ��ŗ
~l������ m�7D�LvӶ�Ez��:L�9{'�ƈdL��d�f���Or�5�Oh���n���!��"wa>��^��ljӜ˓(��(8��i�B5O��6�O��5���x�Vy��O֟Ȗ'W��'8�7?�^h�6�ҵt�j��B��_�d�(�$�D����ג�l�� �'�.�]
60ɖ���j��t���g�6����]�6Qx��fN	���@��� �<�@
�����4|���'Vu��(�>^����1z�PH!BQ����p�S�4��,j L6A�q�ҧ֦S~Z�Yi?�Opn�hAbe�Ѣ� X�Iy��-0�L4��4��$ /f�QgbF_N&ʓ�j�i��$Ґj?t�[�EO;&O*a�F�Ąq(��'N\ڡ�>G��y�ҋz�:f��bܧ/����i�*� |�!g��4c0	A�OX�a�ł�5�,S.����bQ�_A:`�fȻ��	/5��8�r*:%���>��'�\����%rH|ʉ���A�X�ۃb�*z:�sciĺ���?�J>����?�+O�j�F�kݘ�ZP���~�bı$Ko�';���e�p���ئ5�	:JֱC�Xž %!B�&�(٨�4�?�(O��8������O���<i�LԊv( 	���.�n���P
��- �$�;ZJ��e��d@kQW>�j��c_�+R���`['UV�b��6wH<uy��ۡoEtq �0#��z��t�˰���L?hH���DC&$��hѣx��6��ey�`�?�����?Y�	(dig�#����g[��T��J>���IC�8��3�&
��e�@NIC��>�M��i��'��4�O��	�-X&��p@�
3�� �G8�!�f#H�M3���?a����d�|j�O���@�	b��ha�V�F�bq�i0.d^�ca�0��j$�'%�`� Z���=q���8rɂa¢O?R�]��՛P��E*�
U>9:�ۊ��ʼkxj�7N���7�Y�_!�?9��i�V#=���d�&Y8���6e��z���r U3V��|B�'E��im(�pF 5y�đ�Rs*Y`�'�6��Ot%m��M#.��QҦ����<�#dU8zn���,��5�>�+�������'���'��IĄl��t������E�q�b��� V ��ީ^�<�:��<I/.:��'��MK�X0v����1 H�x�T�"7�Ԓfo��h��@�]�|������DƖZ���bӈ��'#R�[S��d6J�c�k�%t8t(L>���D+��xm�,x���P�*1��&@�����Ǧ��JZ
k���ʧ�}S��22$J&�M�-O����n�Ѧa�IKyRS>U�	�cr��K�|a�M���;T����	�R%��)�:r��V$Qa�������f�;��Y+I���&M^-:ׄ@�b��xjP���lTp��!A��F�L��&鍫�Bc>�*��΀=p�c3�Y�_ߒ�:��8?��f���h�O�gĄv�����[�f0�K_)2�!���X�n%@�Z;T���L�.%�џ�@���E�Tlj� *��S
����1<��'��,�~��Iߟ��I؟��'m���!��iCL�8FO�'fHIBǄ�9�m��"Y��$ҲG�1����`ɋ�~�nPx�x��MI�Fk��q���-�FũT�"G�����N?A����c')(H����C_�4�kBiř6���'r�	2mb�d�O��=��HIƅi���F�fH+�G҄�yҤ� b�a��L3pF�4/ݵ����P����'��	�2O>x��ˣS��ԫ�Ǽ/���Y���{�������	ޟh�Xw�2�'��	߄5���ӰF�1��O�'&YT)�1�I��YPm�<�,�SBՊ��O��a��Q(Y*2a�/RR��h6Ą�SL�5�T��K����Ř`"��?!�L=0���4�V>${H�O��$�	�4�	s���rU��.(Z����4 ,P��"O$dZ���2��@�>X��*T�|kd�,���<QT�"�O��0)4�OC�����/�MK�����O�$�O��pd�0���ff_�ڀ��2���%M��ش|�ܙU6�l�?)�x�<	0�Y�G]���!��"�,lb��'M>����ȆZ6X1W"��T�ܳߴ%�n�DyF
�?�����޿kM��x��@.C����aDZ>%��'��'Bl��7c�� �.��'fa5��I���oβ~�9���ɠt�����D��?1/O ��v��Ҧ��I���Oo9��'�
�A�Kǲ	 DA�Ɖ%n�rE�'���"�j$Y�$J�q��!@G��O�I�d��i�r�$��x��1����Ā9	�е�Ԥʡ�еA�KV�P�\��#�)BK��T�K+8����� |��	�Tp����s�)�'*��X(�3�� �T��b}���a���5$C�!�L�jQFZ�RDbd(ڧv��h)�E�u��x4��cJ�Hiݴ��)�.|���?����?*O�L��F�< 8����Ó7.x)(G�K�/C�|b`%ߤX���q�%r�`b>} ��Z�E�����nA� �^g��9j��r|�=a3�[�4w0��e�ߣ��<Q5�iR��`� �'�Lj�*۷F�T�g�Y��"�p����$��\ b�'�ў�3�@�@}ji93O�>"�`��OQW�<�3�4\ʒ�j�K6H�r!E\y�E&��|����_�?`��q�63I�����z����$����	�����ty��$, .�l2���c-��*#�[0W�����=$�s�$���r���JT�����+�(�`iU#TG�)���#�$� F�+;ℭ�vdQ:[�>#>Y�a�$�4ͫ�눚~�R�
��#��O.�d�O�8D�d�AuJqB1�F>hd@S�CG��y��*q����ϛm�a�������'+剡J��@����$��������iD�� ��V
�4�$�O��Õ��OJ�Do>A��@%kiL!<�(��I"h�����*K�
����ф��?����$�m0��9D�C��6M(&�4S(�Av�U�z�(x�TĄrL`�+Td����To�O��D%?�5/`.j����؋C�^���,�n�	K�(a�����3%� I� ��3�O���	�4��`����.J��(��ŝl 
�d�<�Tb�Vv�F�'0�X>�&��������jgN8qjdK��џ���^� jD@R�gqȌ�$���?�O���/L1`�	��G
|�A�B�K��<�bǄҞu���F���h��!`� ��5̂ԋ�5!�`y!U����O���,�'�y�N�K��E�ĳ,'�""!^�yr��J�.�J#n�-�)��כ��O��D��n�N�Z�!��[	[���O�y���'2�'v���a���'rb�'��Nڬfk|�*�	D������hM� �r}�eY�9`����y���6��8�M_a�9���;l�]�$)�>��J�/wb�=�|�<���ۭJIZ���,C�Ȃ��ß�'^�8���?����V75�T��ЀI�a񢐋��3MZB�3_�}�����"|��0����<�q�i>��My�J^��r�3�0.mjݳ�'˯��u��U���'	�'����')�6�4��΁#n��Ԋ#�X	$�<���C=���G%CR�A'E2N�?���a�? �q�����Y��
r���x*�'_7����/�� gV��)a�@�%�ɥXR๘��.AȬ��C�[�
]�G�OJ�*��O2�9�FJ�f�j\em]8,_�Y�0"O�1�0��.fR�@ұC�tRbh2ŝ|B�|Ӧ���<q#�^I��'�2m�O �Fr�V���cߟ��'[)HG�'4��'N��q��g���0d��;Ը0�D�/�}P5�W�$�3ca��@ax�Hϲ#,B<�o��<�l!	A�Ǐ�XY���E82�Dէ݅ka*�q�L��>���Ey��?�Ƿi��6��O�ذeꌫf}� �f��[�BA���<���?IL>E��g	/��k0f�is�uc�/Z7Ԙ'rў�'U_�Fb�y��IB��Ƥq��5e���k�6��O"�l�8�+����Iџx���2
�Y�I9p��I��Q�\��u���W+�i��̟��gI�"j�@K��ԏ@�bq)�	U�f�\]��N�o�T�%6Yi�5��/g����e����d�e����"� *���'�ǡ��%��˚��S
I'�a1�I1iǚ=ZDʂ�jh�aю��	ɟD�t3O^�����8�^��,�2� � T"O�TAa(ôvRfE3�i[<<�x��I�h�R���� 	����� |���Uu����O��d>z���a�G�O6���O��$|ޭWDK�P�쁺d��5aW��j%eӿB)~Cvk�4E��k�C,a4vc>A&������xݤ��g��eր�z�
��;��$�4�2Ih ��( �pc>�%�`[��9
u�2R��H5&���r�ɁJ5*��"�3�X�fX{� 8��z�K2�ZB�	<%\���&-��h�IU�',�\g���B�	���͠�C�	W����'��]�(ER.0n"$�	��H�	ğ��_w���'2��rD4�)"�W�$^R��C0\,J��G�Ü]��ٰc؅z��bVDY3zP�p(��Ĝ4�Yq��֋RA���A�DI�c�`Ť=XBfo$L���!K�p���W�X��� �\�" ���r���`s�'w"�	|�'�Z=�ץE�+�ݠF/��1�&p��'��!qB�O�mp��)�'S���	K>�p�i�S���������Oج��&!eX�g�	��m�Ƌ�O:���I�v�$�O��Ӳ�h������UMӟ@;�K߼P�|IKS(�Qs��	��*O@	��W�R>�ڡ�@;c;n��	��&ܓ��X�lQ:����C�mFaxB����?����
2�����d]�� �mͫ	+�'H��'�$×D	%1���{A��k�6e2	��l�Bo�82���`�D�&���QGŕ3�?�)O�p1�B�O���ʧ�?)���3�p Ct?#Z�S��ԍ�?9�L7~!zqgذB��q�@F�4�����B�N��&�"^/p	�/���I�rȌ����'qG��Np�O��qq�/��IzbD��AK r:zX#�O�Ȉ�'�b���<) �&A��@i� �`\�"�@�<�5���� Y�/G�@E��:r`]q�'���}���c"�QY��N1_��(H����M����?��O*½P��ؾ�?����?y��y7��6f��� �%͉m� z�aS��z$J��A�B2L�e
=Cp�U�����'���*������ߤM+����9+]�1; ��$a�$�{'䎭�n$�#�	v��1c����H\C@l��Oh���1?��ޟ��	y�'�����-]�.���jA�<m�Ů�yb�����dD�=��!bdQ����Ln�����'�ɓ��K�'Ňo����uL\�=j@Q��@#Hl��ٟH�	៴C]w��'2R)1�*i
�IW?d��I�F(��;/H4:��`ˬq��W�Ό��-A�~�C�ֹ(��tjfi�5���o�&$��q�Q��q�W�c��">��$�4�� )���(�BaRD)�)|����	��MC��x��'����>oE�Pڡ%�0B�Љe�Ԏ&'p��D8�ɖ)����g 7_�v4h�,�V6^�O�yl�Mc+O ����Ǧ��	ݟ��VN���b(�@��}����Å�����zj���I���Χ?ӊ<�D�^�N�(a� �I�Z�)�/Ԣz1 +�`�!']�!pb\^����'�20�ҡ�ӫ�&�.����;@cɒf�� 1���I��߃7R��V4{���'��	$.������ C���'�[�}`�O���$?�5��Z>	h�ةS,�]p����O�ժ�"G�X�J���n�7�]a��'0�ɢ:�Z|��4�?A����)Ca���)WԪ��	}�����៧=:��$�O�Шl��)>"��r'���T>��ORL����[��2��Jm�xZ�O����,8�����R�O�U��Z�NIj���"V:���h�O���w�'(����<��m��`����
�7acH�S�<��X�E��|��)
�Mz�d�"fS�'��}���2�e`2�5Y��bWđ��M����?I�Z�*Œ�eW��?���?!��y�/��J��AZ+]Z�(H���2�W�
X|RD�� ��I ���yr���b$2�(W`*`Rj['��;� U��EbRA[�pZ��y
� �8X'�Ռ7��4x.ۅ\����bE(��ۄ\�r����5��Y�V���{���0�M�#8�!�d��6� � [1+���ڇ�K�P�剽�HO�)7���6�HtJ�W	F�νI�֕��}	�,�Z���O����OJ���OJ��r>=p��ɗv�)���;1ΐ�C&�� �����JE�	:CE��a���/�B��D�:i�6�H>-�t���)�v�S�A;`�!�<{�9���I2(�8�+��!`���@��xp
$�O:��;ړ�O�t9��	�L_6�P�쁨8ɸ5(�"O\��Լi�� oά56�)��/�DӦi�IYy�L�
��6�O`�-RN1�#gʈ ���m�y��퟼1gg�⟐���|Z��s����&[����w^��p����TC�� w���u�����OH!����ì9&H5�'�J$�Tl<GM�	�0k5��a��!����-$�G�D�J�X���!�~�ȓp���˒��69�%z�-�?	E�����?q�K'e���5)N�uа���A�{�	>
h���4�?����C8���5U��X -�#6V���1�.bg��D�O�y D�.�\t#�.c��()3+Z8Vz,��.(�7�Ӭ?��R ����T�@+A\~R@�=p$��C���>��g&�:��0cgRH��ځ5� (p�a�Eq����E8zk�	)�~��'��>�͓i#*8��>qe�Ak?�\T��C�ܱ�v��)+q��!�0�޼D2I%�'oP�%	��P�e0i�扔@�ti��4�?��?Q�̇=�~�����?���?��w0p�cSL�q.�9��B�R��H�gC���a�B���<���j�̘O���bV��\?�!�-��{��\f��Rլ6i1�s��M"U�pe1��+V����|B��Ŷb�
�I�g�΀ГL��y�@S%G���$>?�(A��IY�'gl}�C���d��i����L��"O*a5��9C#��Ѩ�?J���R�p��4��Ŀ<� ʗ�}K�#��Ҍ/`X\1��X��Xѧ����?����?��J��O��$~>�{#�.,9 HcS���Q�VT@P���;QFX���-&��z��\x�����pjE�7F�J�t#�"6j Yi�Bۭh+��3�.6�ؠf>�(�\lPG��bٜ���Ɋ%k�5`P���0���P�?ю�iCZE:�a�,A�ps���'&Ү!�!��B�+9��c�9I��Q.M^��'s67��O��Uh e���i���'	�b�lK�X7���&��+=8p���'�2�ޫoa�'��l�og u�7!(G8����7 �$��I�JE�8(�̨1��	�'�*���N6�aGf	p`��ӵ��W`���@��0	�Ӄ2�ta@�@�'V	0�)��֬c����اBV�s��:�U	�������?)���S�O<*��f�H�UN�Ug.}�T��yr�|��i�v4C��
��l���� � ��!g�����æ��ɽAM�}�	�@�Iڟ8�0"Zş�C��&	�ܹ�vʄ�'4YQ��ğ��	Aφ��Pǟ�!�@�E�i��[?]�O��@���.y��\Q�@_�����O�����Ț.��e
��N�#&��lR���G�U��Ԝ��×�
b��I���¹��	�f��̦�3O|����B�O.Q�j�3����N�"�<�O>���0=9#�e�����
9MelE���Cs�'���>)�����S�܉p�GQ�!5|u(�	�?TX�f�'�B�'��TK�*��v�B�'#�'��N�Qd�0�Ǽm@�u)��<R�㣈sO�zb��{Od-����6�D��+Y�K6��/T$x���}�`C�t�4�VF�Q�� �+�d�.>��A�M�%���L#��� (�)�O����ON��"��ĀI!��H���&`l���n�A�<����QYdE2�x���̙gy��.��|J����$�&r��c	�#Kג�p��4q(�I`�!�J�D�O8�d�O����?�����C�pl�$�f�əM�UqS�4`8H@G
Z��̠WGR�N!���ɔ,[��I�m��NJ��ha#�33��U+��b�h!��P�!b����k�'���5N7�eQ׌���"�M�?q���?�"�S!8G�h�&�R�)���i���C�	�k���3O�R�q�Vf�� ��O4�m�Ɵ<�'=��J�A�~���=0����48v�-�F���y��Y��?�c)���?�����Ī���ʙ�%���Hnzi��E��4D������<�<Q�W�B߂�D�B�&���'KZ�=N����e�N��b��[ ~Tx�E+���0��U�I�o����O��A8Vq�����@X�cA����L>��0=y!�!}�f8)�-^H����Bb��؁�w �i1��ĥK]��zC�4&�ҭ��Ay�R�`Ԛ6M�O*��|�Ɗ��?�b�C�N�8p1��T��0�ƠR1�?��Li0n�\jjE�FN�!~���R?Y�O��X��Dޯ9NN�"���dȐБ�O:��!q�\��A�{"H Z&A$�ӂI���z�̥;q"e"���H��Ht�@��џ`F�T�'|� V��p���6)������8"O�`3��D�@ͩ��R�r}^�'�	��h�i��U�N�P�����}����cpӈ���O��M�<�����O�$�O��dgޭ�pcE�7l����0�`��>[�ر��X�0��#�O�!w8b>=$�Lx D��")LMp��3��p'�5,�Vݑa`�|�� �1��D��t�|"�R.f@.	�c�{�r� _+Z2�'�z����Ϙ'@�B#��#r���7���N��y�',��S���7�`��@�2����/O�9Dz�O{�'��}`��M�z�lQ჌IR��x�� TB����W�'���'��mݥ�	����'q�Ut�^�`^і`R
"���Ƣ��P�&eK�M�Yg���d�%~�>s1��;R��="A��=�8i��+$��)*�*Q��p=��
I1 ���fbQ��4���Љ^Eְ����M�C�in�O���b��@1?Q.���+K�p	q��dg����?��#ɺ6{t�3��źN�d��7�c�	�MK���.e��m�h�$*6&���[�mț���6I��0<���c�'���'�]�z	��rq'�_�0��
Ó*�"EFxr�>T#� �Ո��
a�l�0�0<!1����<YVM��u����c�>�.P`u�t�<I�lV.BHZ�E��@���G������O8(�K���ir�}x �;"�Z$$��v����sl=?�(�2�i^�l��3�@�Djq�`_�dP���O �0Ǉی
!(MI��	�Z�5�)§*��)�Fnz��zS�����(�'�*p�`E�DY��xCcN���>U1 ��*�z�[b���Lq��x��>?������	q�O���3Q��E�'�Djr�� �ˍ�j�!���=cRZYI�%�#^,iSm<�џ�����͛ju��`P.E�H�0� ެ'���ղy���5C.���I�?��	ʟ�'u�y��f�*��X�B�@���eZ��[�j�O��hн%�1�1Ob(#χ����#��R�x�����2�qRi�O-VSA;���y���g������-^&���A��?��O�@"�'}��ɳ'ɘ��S+�h*|l�1+ �G#�Y�ȓ�vI�ua�-�j ��J
5��'I�#=�O�ɣW�*�SW��|�q�gļ?z���Ҹ|��$1@p{d48�aR�&�(�m�	 )��GG�F	���;//��W�I�@+8�A&��F3�=�� (����	ٟ(��@��I��s�H�+9�?�'[�u*a���$�V�V�/�fDE|b.�<zj�츐F��|��S>� ���@;���A$�ȸpDa=��Q�	��l�|�BI�)P4�����5����)�xy��'�r�V_HF�`�U�����y^�ɛTFdE��R���Z�^7$RP�I�P!���?q����i�@m����O��H�oڳn6�m*s���G�����O�}�%D�'`z5�̡b0I�i�Y6.�S��+��6#����H�%S)Z�JG�^�^�	�v�C�@ȵd�4�F(/#�m���ԿdGq�\�'��,A��	E�^�h��0:O���'b������>��{1�@�e�T�'�ݷ�r���.��xR f��j߾�� �CupZXF{�f4�O������/N���5�@'�������?I��?7r��Խ�?���?y�����e��ڱE^��8��L�1�:��F ŷ*<4��v�><n�b��׬��i;�I�[�V�c���f
����,gF�!�V�X$��"êz� Ys�`5��46�4��O~��e�0M���R��*\pq������OZ�$?��y�Ie���g&�&;���yЍW%�yB�\�Dtp����,3tp��=�?��i>��	Py� � ;�f���-�)J�fm����y�	���'�B�'��V�b>�զP5.��b!��!&��4A�΄��P���j�*���⚍O�M᥅P����Gy��U a%8Ub�A��J�p�x�"7g���q4I~�؃G���`MҤ�E,}� �Fy�h��?��S<)P�ӣDM3K��1�TJ��?��,�+IBlr7�S�AI�)"3�P �Fh�ȓ7@�l�FHϭH��b��#"��'H�6M�O(˓,�����IK
{������>�U@ 	Z�8˓�?���?aTdσWԢ��EC��}'��a0�V#}p�h���[l�r�؆ZxDe�+O��1Dy���og�m���h��cqc�6t�
�����m���ӴPx���A�
2JF�9Dy$��?i��ɘO��i�IƼ�j���$��4�-O2���	�X�i)Dkt������}�!�<	g&�(����S�18�Q#�őfy���z�R�'��Ij�T�'�2$�/q_�@7 �9%��4��@�<��dNj,$R�jG�H��Ԃ@ψ/G&z�Aw"��O�&����:��spJ�"/����'`�����Ʒ0�dۑ,�v�&��垶 {nD�}��� &��5�D�sf�EA5K��<Y�M\�x��X~J~��O� ,��bAz��u�&%�$?��6"O��z�	�..ʐ��T�7V`d$P!�I7�ȟ:�;���M�q�Z(
�8����OL˓x�4I���?9��?�(O�	�� �d�[���6���:V$B�0w�iC3��O����s*�tJ!�?#<Q���L�JS�eDj��b
���
���}3��%�1u�M��O&�1���+ɰ|���u��]{џ�|ᐯ�O8��9ړ�yB��=��i`6�B�.x`��)
��yB(_�lp�@0�G'wȭ���O �?1��i>���}y2��Eɔ��A�ӓ�X0��><I\tZu�'D��'��U�b>!�#R�<�Pa�ڧ_����6>�^�w�,&�8�2c]���<q�����xU2u/ږ�R	ʃ�}���0S#�&`�2���;��<	c#��0`Ǫ �΁q��9j� �����D{"�I��r(�E�Y^b=��nXV�C��yގK&��P/@�'����ʓɛ�'��	�x�L@����f>����K-5pȀkS�(�Bd!���OfTЧ�O`�$�O����B��7]6jҢ�0)�^��i>��#�]\���F���t_P��'�>�5C��l�d�RȆ����Z7�!)�f�xg��c�X/�D�!�O���*擟a����_j���4�țp�0ʓ�0?�s�tu1�=W��VH�Cx�)O �i���}�2��ƣ\�7�Y�rR�l��Ο���Z�'��DۼQ;��b�A���'ȹax���-5��$QRd����/M'⟰mZz��d
�O�Ҽ{姉4���3#�1&��9�}�Z���9"�d�ɽ�l��ON�)�O��	�v��5��J��?"��E�<H+����ܦ����6��E���<�U}nz�M�͟k����:5M��t���͝�H�K��?QG����y"��,�$�Or���Oz�I������
P��ZAO޶S�h� С�OT��/����v���
�?7��B������Y�@4@Q�J$fw��[��gL�	ԟHbǸ����O��$�����͊Ft����`�u�o�.`?ry���	�B�$�O��.�t�Dd�8H�k�?7�� ��;>W��Cc✤KZq�㟣%`�nZ�<�ԉ�۟���Zv�'�?������_�dҨ�2� Ρ��Уs�2=	�@�'�����?I�����h��r���?im�i,�A�G��%����33�&ii��ԟD�@���ID��/&���?��AbE�����2)t����%�BZ�v�H0k��DN44��'����'S�d�?)��}8���_T�� ��͚B�|6m͗]���Ĵ<���O~��D�����?��B����jY�bO]�::T|��)�*�y�M�|�ܐ�D��6s�1�c
�$�M+���?Y���?����?�+O��$�Ok씰�Ȱ V;HVL�8��K?�	H�	��'&�h�	� K�ɹ�A4(�b�X�!��W���'Ā}"`� AĔ��OB��%O�����!�pRׂ@�8@ "O6���催)��<�5a�1+$���"O����j�b}���R�|'���"O���E-�lJ��$ ʵB+L��t"O��l�"0d3�Z<�|yQ"O�}�w�,i�0����
k���	g"O������l8�)�m��G]��a"O��6�"v��U��K�j��њ�"O \"����s0K��L����I�T�Iß��I��Ԃ�l� �x|�F�@^h��0+��M��?����?	���?���?����?���mL���HV(Ci|��S ���&�'��'~��'���'�R�'V�	-u�r=�fV�L�T�'����6��O����O����O��$�O��$�O���].��x#�WY?��[5 J+0�jEo�Ο�����X�I��X�I����̟H�	*�IKF揠a ��Y��A�[�V��ݴ�?���?���?���?a��?i��X�0i����>po!:���01��Q�p�i9R�'�r�'!B�'���'\B�'����M 3�=ⵆɲZ4��bj�6�D�O����On���Oz�$�O��D�O�b��v&���h�@���JNҦ��	՟��I�$�I����	��x�	��N"Y4^�Z֍�%$�R�[��M���?���?���?����?����?�$+X$.R��ӺM���X:f��V�'��'1r�'��'%��'����,a�6F_-'h��S)�9��7��O���O ���O�$�Oz�d�OT����RN��v��PJAGG�)ioZ�� ��������P��ϟ|�	���ɤA�Jx�4���0�/=$���	޴����O��Ɉ�m��鉎~UiN F��0!'�v�Z=1P�D ���M�'R�(9����x� N^����7�'ۛ�0O�S�SMIjDl}?��b� 
dE"Ⱥl������OƟ��O �R"(�놌�o����1Ol0�o.�i:U�Q�c�l��'0�	m�I��M���h̓�� |� �?|
�V�j���Q���syb�'�8O�˓q�Ra���.	|��q%��Q_JY�'�$�jg��I�L�!�O�i�&�H���y��6g?�S'#T%$�<�1Î��d�<9���h����0[�t:�g�9� �t�����oӘ�cu�����4�������*��$mZT���bf�H�z���O�7�O��(
b���I]�,� d�]02�ݠjJ�Hy�ԇ\#*��FLZMF��=����"�
y�l��������C1�ةNzʓ͛�L���'��1ps�@8S��h���P�q�%ːEy��'k�V<O("}J"\�Z�P6(G��H�����'�&q��Zp~��7@b|���fNd��*%�X�M��ᓵ�+���%j8����E�<	�eD�f02\`���%W����aCJ�V���ӡ��$URX	��N����"�/5����|o�L���~������
�+,�`�gϱVRd @�+�>Y"v`��E�H��f�B�jY2e��2C�9!4a�+f%Jx1�bgm)�� �7�p`���?3���F �3�ΙH<<`�Q�����({s.�1��}0�d+"Gzࣵ�$a�@%+Ec+^��5�B/6D��H�m�P�VݣLG��XPw� ?�TcX���म��q���q!��H!@�D�R`0�����Y�D��L
B�F`V�+���r��_�I�g�ISp�5[ϖ6-�`A�4C��pr����f[��D9����Nq���CI�/$��	�&Ǜ��j��ƚ6�@#��#TX}�i�|XU��O2�PYݴ�?)��)��J�ሂ/��%f	BvXy1��?yJ>9���?��i��?�O��I3O��r+�K��F��?����?�-O��8�bNt��ßx�Ӣ#f�Żf,��~�l$�4l�&��%� ��؟�����$%���>���_�NP�=�dM�����ĳ<y��X�]śW>����?1.OT�� �6]���5��-,g�u"��'1��'m.��P�'�ɧ�O>�)w�� 3�1���N$-^|h��7��I�i�����S���$�O�ܚ]��M�Qoш(����qȠ\��d�.y�>���O���1�SПD�	�2�(#��1yͰpT)ˁVj֌1�4�?I���?�W���J����I�O牦f��eU2~}����	X�k����OH��O.T���|B���?a�����C$N�<�w ˑ�����O$�č#H�l�ş��O2Y�<�I�zC�|��L���ޟ)��+��ݟ��	����	����I����	V���'��i���ݯ8Nd�����Utu �j�O���O�O��$�O �p�eY�4�j�@`�G?I-����%��U��Ķ<���?�����$ʎQb���`ɒE/!��àB�=����?Q����?Y����b�%0(���N0=��PP��P�lk/O��$�On���<1C�[	q&�O����d�G,�,�E�� E��r�'G|b�'F��>P2���X#ϝ!Y�L#'�H0W�P4���O��$�O��$�O`d���@�u�	ҟ��	�?�&��	��k0��},�mx�GScy��'9��'��'	b�'�Ӳ2v�EXIT!
����%6�d���O@�D�S^�Un��L�������?��z�\�3mD�A� $��FR�vw����՟����P"5��ڟd��k��*.�)��T$l?Z�iQW�{<�t��UI�y�ói�Iԟ������O���9����d�+D��k���%kvl��S�cP��$�O���$�����Ɏ�Hq�� 1�}�����a� ���4�?i���?�'J�5�����'
�G�B��8���D
�a�֪D����'���'�,��f_>a�O��=O8��ō"m�0h4��	<�.iU�'I��A�����$�=P�f(��ݣH^���,�D,����OܲSc<��ϟ<�'�_���(ȱhڮG���"�-(�ԡA]��	����?���?Y��?5�4Rs A	W�:d�vH��4�LqFx��'F���t�� �|�Q�� |����O�n@����N֟��	ʟ��?I��?��+�F?I�E�X�D�@��� �@hAW��̟ȗ'eg���џ��4��t�{�,
� s,`ע�ҟ�?Q���?iV�J̓�@�Q,Q93,���C��z��	����?�*O��d�x5h�'�?���y���>a�h9�/^�l�$�FLI>���?���R���<�Οެ��a�F줸1�[e۶���'��e�֦��O"�OŶʓ.q ��ZШ�G��K����%������Ѓ�F�P&?u�o��'_s�t G$�?XL���2[r�W�uc��'�"�'��$V��'���U�<)j@!�ƍU����?�F�>���h�0�d�+��S��� �0FÖQ��n�ܟ���՟X�!O�9���|���?���$`;�Q�7N�S�0��ʑ�?i��?���>�4��+���'}Xq*sgQ�I�hM���Ù#$P��������&ԱC�&�A�c�1 "�s�iMm>ze�4�'��'��3Oz�:tDF�n�����[�R��Iۅ�|��'�2�'tB�'B�К'2�W=Xx����:_�.$��J"�'џ���ןx̓���֮S*wâ)f�0��G~R�'��$�O��d|>	9�E��k��� "ˑ��nl��c;��O�la��8*��)���O"������S�&-��D�s<��J�͜�C�I�:A�MaW囂�j9�F��V�Rc�pX�:V��$i��\iD#�A�odtу��M�lP"��4���;mz�R���(8F��ħǭG�ryX'�*O�f=�B�3s�,�������'��6>\H�G�|�� v*e�?��X�7�t���͂�]�f�#�k��O�d�wi�3��`+v��)<�*��HV-:���u���e�Չ��F&r����/J�I��T��?i���.؁��	H�L���PG��q(�?��O���:�F� ;r1"p�A7O�\Q'�+ .}�ޱJ �S�3ĝ�BFZ=\���\>��≟?2㤕� 
0&�!kT�.�D@`�2�nӼ�n�؟��~z�	��hLњB@Px)�q[��ߕ'��'42�'�P���	ԟ��� �t�g )i�0\�G�x�!|��LmZ�� ܴ�Mk���/,@HŸ���7����W�E?'A�7-�Oj���O�̉�b��hU��d�O0�$�O��X�n�P%�S������ nd���f"6f��Vȑ2F8�9�!��O~�6����?�G�V#��dy�	�DC h�_.h{�5x�	�
g�L� �Bǘ/D����D�i0(UϻH(��Q+��(ܐA�ꈓ4���Gz���'@��	��|����'�8�
�o���I�+�&Š�`
�'� �"�\ i�� �H� I�D�����զ���~}B�;g� �p�%j!4��0��]DBp��. <�Z���O6�$�O*�;�?)������K\��]�%c$�V��!*�>N����^�iE���K�-��!┆'�c��#.Ѳ{�(4��L�g��� .�88�t:[�����E0>����1&���Z��¢g2Ew���GH#T���-�O�Z	b�T����
�o�&E�� �y�!��<ṱB�*5���	��[�¸'c��PdV�M����Mk�C^.7�>�fb�: ���$��F{��'��*��'D��'��<hU��5)Bt����΂u:�[��Vap�l)9_��RҦ�TX��S�Ԑ{`8��F�9�R�*a��&!߮xi�
�z<f�7+�$�����v�Q��h���O�	nZ?�M��4LX��pp̄>!��!�3HR�K��$U�Drߴ��D+r��4֧tch���.h�Ѐ���x�*�l�F�+U��3!O�A�#�)�V����i�ªi����@I�Zg��$�O
����T�F~�ƼySO:mh�Mx��Ё*�@���iLٟ �� �ԍ�R�� O���蠩����3P?��O���Ѕ��) ҭc�m�h�t��K<a5��1l�X}[ aT(nD���Z,_��S�|I����?�P�9�O!�t�'2��O���t�fm�C�����U/�h��"O<ea��P�d�Z�ٳH�9R��=X��V���d�&ʓ|3$� mۙL�q5�W�)x�g#rӬ���O��OPЀ�O �d�O ��wc8�����i���R�"'$�H1�p �6����U�aӲh"��,t�t$?�CN������^����1�	89N���t��fa��MW�M�4��)-�6�`����i�k3�f8�"C=2�pd^6)��:�j���M�WW�X!`��O���=�����mڼs,������h܋a���u%�̫�'(�����)=�L��G�R�ԭ�~��'�X���?���h}bE�8��@)�%V�S�=b5��:6��6�%7T`�$�O&���O�D���?Y��������%Cw�T7�4x���� �@��n��`��`	�(�]���P%2��bw�S�b^��>\���k@N,LO��(���K�0���R��^������R���'L-2�l�;���Ƨ��B�Y��'y�E���S&R鐠��!��_
(�{b�,�	0 gr@"۴�?qߴt��Q6 �-���j�d��(�qJ��'�Z5 Ab�'��)U3B�"Fi q$�MY�S%A�P3��cw��0=�I��	:Ⱦ�:���-����� "i�ј�U ��h��19��Q�A"@Y��ß<�'�:,(Ї
��!޺�� ����~��'�2��I�,���R�I6���A?2����)F�<m3��T���K�2p����'���V�����4�?9�����&}�&7M�]��T�G,]�sw�� U�Bnz$��Iݟ�X%af��@��Od󄈀��P���	�~r�	��ZT�!i%F����  @�	���aHf��" �xeA�m�%$�ĸ�}P�
�NZ���"
%p�ȡ(Oy�!J���ަ�J|�K|*�*x�=�ѫ��MҼ�Ct�%�qO���6�d$���LTvE�ԏ��d��"��c(�����!��4��ah����R�bݢIq�!0�T��h�N�D�O&�$T�j�����O����Ob��w�H;���`2�qg�(���	��Ťz�D� ĉA
�(�o�b����']����D9��X�F��#7Yr�c!�T0:���؄Q�̐yg�J�ym^�>=�@Ê!�y'C��N`�&��8b��Q0L*N2��$Ty����?�}�I��n�B�@�KT��!a2�[D�8z���^eqO�X���P�	�T�D�1ෝ>��i�7�!��?��'��Ipr	�&�b�±kI�fb2�*�)ݺ�đ�O��d�O��ďݺ����?Y�t����%�/��C��DT&E�ÀȷB^jH��(6-���"C=,O&P9 oJ��p}����S�����2����-;����nPsX��Y��ҁ�j�k, ܅���^�X���O��n��� �'-���t��j��"t-A4�ʸH����	�$��R؞�K �̓i�N-"�[��&m��	>��s��&�w�˓"�u�%�iVұ� 8��wX�{��Qu�Ũ�՟����.!���	ϟ��I�Qm� ��ÖxL9�k��
����5K��	H��6G�#Y�����'^R�k���W�αh��#A��y#�ߢTB�W);9B�q��."�4�K���
�4��eh�P�oZѦ!Z��X�e#�%�rh�q��Xql
�����-�?���)�~���¡A�)tYd��7��$TC��d�J�=ZPk˙d�aȥ�uf&��'E�u�'�>6-�OP�$+�Y���t�^�Ix�����}�zA�SI$D�d�B��7ӒpH�,ԉK�rUҡO4�	�u�4ը���3�ʀ�fd�c�P�Ol� w��(y��]*rHH�7���8�"OFX����&ܺ�WFƽw�h�8"OHVeթ1�rR��B4}�&��"O��
����>M�.4e�8���'ے@B��?~�����P�Թ�	�'<��a0�O;1�tڰ�IP�
�'d��Yt�@%�R����Q�L�6xq
�'�H�p��<�8�)��޷E㚀0	�'���� �נ`7N�rW✔�j`	�'��|1���)ST�y��K����'`B�AAm����F�XF����'��lZN���,���N�~��	�'�HI�1�	�a��<�Iʼi;����'e.�#3B[�7�<B�E�k�����'��(E)(4���#��[c֎�;�'�Ν
�뇳GX����? f�Q#�'ְ=��K�*��V�%ނ���'r��*��w�x�e�3�6m#
�' R���l
2t1`&�y1��:�'�I1'g��O���Ce-<b��9�'�Rl��*��>��ܲBEb����'�x�EM�@���$�� �$�h�'��D��M)i\�Bg�����'{P��S���:��B�
���'�
�����0*��1�$J���v���'�1���*<��4i40�
�'��qj'B�}ޠ���F�yB�	�'�>50�C�!dm�m�S͕&Mo^�*	�'�BD��	^x�l ����o�-��':,Y�0�<D."���@��s�����'��h;��[yP��c�0L�	�'@�Ș֯���6H6R	�'������P�"�"в]ߨ�0�'��}J�HN;̎ PMJIW��
�'2�����_����7ǗY^h�
�'�&���
���H�;��Gn�.M*�'m�5�%D�q��X��'a�m��'ܡ�g+/	��\C#�"h�v�9�'��$X��Xj ���HX%k~��*�'����.��^�D����fh�a"�'(yZ�JP�#�8�"q.�S0X��'>��ҋ�6���)�C�7UH�
�'�HBd���Xֳ0�DdÜ�y���,�|e�R,]*��B%mڷ�yr��5|�`K��I$^ ��2���.�yB��X�&�CULӓM-*��#G&�y�IӖBG>�i&L��C�J	�d+�y$�9~j�V�(=��ȳE/˂M!�C�I��d��㋊]��@ZY��!�'SyY��_&�D4Pr���5��'Jܑ�Dճ?�Vā��8x��{�'kr���*��'}l4J�$�
LZ�x�'���R)�-&�:%
��k88��'�>H�e*�^j��įO2Kd��
�'9�%���ډ]��h��Ȯ)���
�'<DBcO�4)_� @�� >;�pq��� ���!oD�Y��)QM��k�=OD����2�p>����2f���p/M�*��}Y�X؞�q��<.�����'��L��O�.~��d@O8�� �'I�<�օ!6�;��S?:/T1:�y��ӿ;,\!�D�k_�F��!)�y!"C��$غBG �yZ(��a�]@7FT�*L�,ُ�!aa`D�?Y!�4����I�����H�i{t��S��C�It]P`h��*S�<$sSN�:EyX��E�o�
35Ⴌ��ɭ��l3���#��y��@Z�?�R��S+F~}��〶wT���➞c�H�4	ɺ)��q+�HƹB1�0�'����L��!D�&؝��aPI<�C�B�84��� ���=s@`$�ӈ
D��Vn?�a�$N(`:B�.���c@Y1'�α��mgV*�b !Y�=�	C���;.�0�@�#�SW�	�n���%c�-������H�
��$��{�B�r1҉q,�E�uf
�/�(�'�D�y6�x"ٶ^o�D�o*,O�ajt�R�8�@��sL�*Q7���'��h*�FN��^�0�㖺}��0V�E��lY�T,{Ԛ ����b�!��|���p��D P#n.��I;?�T��Rl-2�\���T�� t�ͩ焃4V�ޜ��$�
�y"dϣxeP����W��,�5�X�HI�����
dR��R�j
Z����L~r�J*�DIor�[�	쮙�d*�5�a��Z���TA���+%�	�di�/.�*%��~�
�M�#H�����/r��򄛉n��|�F�.+�Ͳ^�\]�����7lx�drCɖ�ru�#��'}�@`����I���N��9��	�J�B≓� 9�-k(�:��J8l���fbA�0��A]��Ã�
a�Q��6�S�Y[��Z-O�*�n��EJ��C�2�bX�5��
�0�g�s���`�+�7^��H��a��Pv�aw�*��C���Q���;��k�R""��>y���	�=r��z��)2�x�{ؑ�(E	]V�B@R�Q�'a��\�T��牐,W`��j7�n��0·�Y��">�e��OwH;#��{��h�˚�"_�0���D"���!���L���g�]O!�D@�i��뇪޹+q����X����޹|���g�MӘ	m�������=��OtBe��Ku8���,�m�P�+�'���y�ڧ~���Ũ-(	�	��PѸQ�G��=)@��"gS���>(BO�Y!���Ft�Z�EF'HIP�F�'��x O��h|q�惐$���""���C�<�rDpf#���b� /|R�8�2�P�<+�	�+����&!��P�D�-��	�� �!Tq�mä�$����'��4@�Q0E�b��N�R-&�2c W�� s�dP�z��!��d�D�6���dI!p��1�朶M��D��
K�J'܁{k�E���էA�&���	a�'T�:蒧lM�BlZ��Ư..~i�G�B�|�.��d�)��8���:C;8ı�1.y���@��'fP��c�OI�8�W>�A1�Qu�'eV�8d	)��(���ͨN��r��y�Ԁi�йhZ��pFP�li�1�K�&����&�H-m H�nV&��{�{�ӌ\�˧!�8L��h�jZ��*�+�lCRE}r�[��9���+Q�r!����#�>DQ�oJ�0�bAЃ��q�(��2N�%�?�`Fim�?���"1Rn\	�@ɠp��HB�JM}b�� N�k�'�)RdP����+4�"|
c����I��
�$jw�XطZD�<Q�&\KVX<�%啧\���j�l�7h�a�4%�"^QZy��˨tˎ $?}�<i���?.5��e�O>�J��p<a���$Y{H�*���R�d[6hܡE�����/snB
�/ְd����dȵ8zz}˄�:%�E/ay�)W"u$R2kJ� Z�II^��/��$|"Ү�:U�0B� JR�;'ײ{�2��Ճ"<q�CC���~�UCV�pcp��%"ʿ4�*�:D�|�<�bC�S�b|{��;6X�+S �G�<�=rYZ���Q�n�bpJ	K�<��ͦ#n$$@S�8B79s���N�<ɀO�3<J92G��2�4M0ČO�<a��<�~d;T�5\�]C5)�I�<a�kx�f=(a�ܲ%�vTSbE�F�<�D"�]�Ta���סq&pKA	JB�<qR'��BH0�)��6[�Z���d�B�<�v�Q,P�]�q�_�"@�kA'�~�<!�`�;?����G',0Ti�a�]A�<� �2d�LQva��HB2PA��"O�y��Es�@��D�&YJ�bR"Op�3$�C��U��%��Z�.Uh�"O@��$��C�Fщ�.M�$���""O`ِ��B�-$0�b-��P0L�u"Oxг��V4Sn��1��Ǩ-<fx��"O�� E������p�閍+ uQ2"O�� cg�j��Q(�(�>7�d��"O8���"�-̚�ز��[�*u{a"ON�֢�T��[�A֌����d"O�P'�]�����*��H)"O�e����9?�kV�� Q�j���"O���g�9KQL��7`�>H�Αi�"O@�a��F'H�tT���>˖ *�"O �b2 �6���M��i
\��u"O�DsD�S�	9���w�Kk����"O���#�F�c^
}RE�ӷc���"O����.���s�Ƣ}���5"O�-[S�b���z�lˠn�&��C"O�E�W�r?����KK$0���2"Ot��kU�@ư�he���`^ڲ"O0Ls&O��H�n�+x$���"ObT�jr���Y���& �I�"O@�w V����V,Ҥ7��kQ"O��9p�ø:�\y[ua�J(P���"O&`Z��_P�Qp�N���=)@"Oe13��*M�R��'/'x�0U"O�e8��m�<CR��9ep-k0"OB���摦m+@}P͗�lz�c�"O���#�\fؕ���I�q��(��"OD��!S�H�r�c ��Z��)�"O� 镅l6���;�pI�"Ob�uF �����ÇC�N\��"Oj�y��+*?�ѡ�!̬Ժ	 @"O��9ˊ0&Mk��_�U�2��w"O(ݫ��E('��GOP�`�ڼBQ"O�5j��D�=u�� �Oޕou��5"O�ܛG�ޢ)/�|��c�-8S�P�"O��i�i\�`\�P�3�Q8	B��P�"Oe�Ռ Fs iѫ�;���a"O@�Q�GׅpDf�Jb� &S_
A��"O0� ��F�.���$k3��"O����j�*D������o?���"O��`F@S�j�# k�m�ʰ"O�͢��[!**@ϊ5�#�"O"RцY�L�UZ���G:��2"O�ɔdZ  P�7&%L��1"O� x��ޯg�x1t�J=�Y�a"OĔ���G1jѬ� E����A"O�����g�TTQPᙩVT�ah�"O�]���b��,eQ�S����yB!�	�^�0�C��m��qDL�(�y�b�,p��v_/XfqR�
�y҈�&Yq���#�I���U E$Q�yn�,+2�%bļac�Tbn��yȑ0�8��GeL��Q�A�A?�yb# �:o�i�a!]O�Z�
���y�)�1+�i�	O��-z�j���y�dO$|Ҡ��9?�x�����y򬐊���0�ͼ$�5A)�:�y�GҳRv.�k�� UF��1!�M�<�F�9X ���֤"Z���Nd�<��J�xfn	�
O&S��e���Hk�<A��1����#vL�xC���<� h(��Kޗ����'N�M(,B"O��r-�MC��C�������"Ot}��F2S��ŉ$u0���"O`���eٗR2�s�OV�`�<��"O��2��0H�A�C��$Z6\K�"Ob�s�� h��sa�ǹW�ָ�"O��6�T�,bLC4@&����"O�|C�ơ?�B<ye`U�E��y��"O�PA1���0��PB���Bd��"Oz@x��x�
YSӊ&K���+C"O �)��ǅ|�>j���G��|p�"O�Xӂ2y��)q#A�V��ڇ�d�(@�bѻ�����#U�H��'��4�'jD�dr���E�Y-��9{	�'�ٙ��O�`´H��0{���c
�'(����(	Z�8�)���"~ ����'5�+d$����4�
}U���']�#�i
aJ����a��}�'�,܊!,�C��$@p+��`����'J"L-){
L1w�Ѻx3�Lsv#�y�<�v`_�U{Τ �'W�;�l�:���z�<	�#�gp�:���-�RV�Gb�<���3C�>�1��O<u3�q�Z�<���6خHQ
¡kL2pQsa�X�<� �6>4��nC�Jo
ݠ@��U�<a�D1s���#�{U�x`ӊ�k�<�1��1�6I��A1E�^��]�<��EB.m��k#��):4S6U�<�PbQg�&���(x��0���E�<9��N�Vx�,�lPv�.�:��}�<a���![Cqqp*��/h��"��E�<!RF 8���P`W�"�.�AG{�<�@�-Y&�kw�XUX<�F
O�<���*eH��(q�	����t�<!E	1I����5C�<O�v���DGm�<1t��)08͓� C�]�vQ�B[D�<�R�OfH�u����	b�L2С�K�<��J&jB`"և��t�q;��1T����(\�[��`�A錤&�A[c D��ʄ�˺x ��1�� �L<,X��=D��Х�%�ށ0��-��D���'D�$��剕)��Xj7��:~��
�1D�гB��0���Ţ�2��s�./D�U�&q'�٩��ȥb��)�8D�a�Ą�Pv���C��,D0�,��
K07�3S�RAG�4� '&(1��E����ݤb!�D�6q���͐
w�~,i�i��W�hQo�9`^�r��OT����Y��XG�]Pl�#'�R3[1T�˗�8D�D���G�8��d�wm��Q��%�W$\|5�FY�=W���/LO�C�nS�H��q�I�}�Hذ&�'��}��IR��1��wV���&������	�3�t�ȓ9dBb�� �oL� ��-@���=A�� ��#� L��#|rq���|�ɈN/��8�gIY�<Q��\*q�d���'8L:tY��/J7�̤�F�X���?Ѻ�|�'�J��D��sZ�2�`��@���!DpЉ�}��h�DzA�&�1�Drԁ�8F���j�L
z��\
��ɕU�P)2u�=}� j��5\OL�qK_?w��bq!�2f`.�����=���i��,�bi 
�'\�hE�J�Kɼ�	'�]TX�=Z�{�&
lt����P֊\D��"�t�$�&b�9}�\��%Lݪ�yB@@1a8<�� @�(i���A*X�h��˃�O�4���'A�EE�,O��"h�?q���H�+!">�s�"O6�ZŅJk��8�Ө:5�]0�i+�Q�g�1'��@��'U�ي$��p^�
�����#�x��P�V�p���FJ�*Qt�{�L!�i�QO>D�� t��Q��V�Z���@N�A1u�	4Wt��U��O*�3`O; �`�:`���]��HC��Cv�����x'$=�B�ֲ^҆�����Q*��sJ�3h�n">Y�C�0p���＼���Y!5A��Zހ[5K�:�y"���fՠ�n�_K2����1��'�2����<�Q�Κ9�~b>�(c?u��2��
P
�l<�O*D!̒�yR��*�}����H0�P�e@5$�>�S� ���J�AU����')��[�	:
�-����~u����OuY�e���M�&Z�-h6e?�gy���xU��c� �b�̠�wN��I+ZЊSM*�O��H%/�5,~P�#ң/\��c/�r\�������]~��O�q3����k�;��x:�H�����^o�����cr��֏�^ L�RrI�6lڂ!����~¨��y�NP�x(� �M;��$� C>��үG8=��`�'P�s�џ�6LZ�^a�U�c��� �� H ���.A�={d/�1Pt9���:k��lڒ'��'h�h�G�[p�'���	��'���W*��Bu0+O`�B�O� �h��ɜ"�BlcZ��O!����@ 9_vD�'Oڃƕ`Ĥ�){���I�0�0��`��}���`��h�h%w�*L��ۓW�(�)��>0<��G���oU%J������ēX�I���!�3��7@��C!^�,��\��J¦�����'��<Jq
d���Z/"��I&����1��(�4�wKW7T�?�2�׌{� �rH���Q3��T.�ΨZ��9p��8aP���laO>aT�������9����O~1�'��0 c�ƥ:��D)�h֩]�:�A�O&��VBɜ3{t��N�>F��ԺP?O�g?Y�$t�d��G'/��Q�a�?�#�����D�1Z|V��-�[�Ҵ:��L#IND�j��Ynt��%U�3��5��LT!F����^�?�$���1ϩ>�G�:*����&Y5<f0��);d����a����|�.��E{��@́:ސ$�'@�<q�2�[�#D�a{"�O&=Kv��W�]9i�D��.~��L3P,<O���PM0V��>�px>Z����藼B��Es��;�A��㧭	�h~�)�GIg�p�I�(dI�k�6ָ@�,PTH�e�R�49�$_0 �C�L��~��;+ܠ��j$�IT�KnP�r�G��բ�ꋄqd�ɷ;��j�%�$�!'�ׅJ�(#=A4��,l��	)%n�H�<�sd$3���4o��@8�)�3 s� �Ӓ~�<�h="�+V��5b�0TN�2Y���(R�"5Q��Y'�K e-� 5T��6��7s�>�"�ϣ|(�1QAMӸ}2��;<O�0SE	�9��:��\5�l��W�݁o�|�?9���9�qK�j�2ػ�Ћc�1+w�8�����#h�@5sd��"}�Y�c��>@���#����Ƃ<�|6-�,[�*�K�L��$�j��Ğ32Ͱq�Z�
��K$���&���6'�;W*�I�DЩd��h��Ծ��t!B� k����ݢ��H+S���0-�I� l���NJ�z��k�D�u��"=�e9�ʃ䟱4bٓ�

 M����+�~JQ$�n �O��I<[���jYV��&eW�0o��K���
&��E��mՊ(�v�����|�c��Jj֬S���*���ચ�AJx�����|��4cI+*�*�O:�IK��ߓY��tL�=r��Klf}�+�Ƶa�
���2�F�#����W�D" ������]P�x��K�C9$������Q^N�KW3���6�N�IS��d�A���ʔG����O��IҞm��`]/*��M{0A�� z�(�"�"�)[ч�K���E�<�H|��*#F�x��.qXT[�K̽X)B0@�i���>yT戦U\��Jb���`�"�"O�'�iY�iE�dV�y��^<bor���N"��ɣ(S��ٲ��f��U�K�#���dÓH�TiᠫN�K�����F����.zjź` ^��	�_���'h��2�$�V}�"ľ.�^���㙛VLV�!��� ��O:y�B����'��t{@H]"��y֯�([�zTb�$�ɦ��Gl-}R�ų�D~��	�[�� �nOԞ��'���ċm��Px��/}b��7��y��~�u(�_�D��sgB9{þ��c��pR��A4�O�- Q��H�hl`s�A1>�T5*A�>���@�B<^�kV��<i@�Ox�P�T�L�`�Y�_��lЩjL��+�L�f��M��|D�91�X����#<�L�Д�ೆ7Ox��L<��z��a@�lcP�.e>���g��}H8<�ȓ<V|@�C��. ��2T��8E �g�D��@���?�':�@�&�F6_�<8�.%H5i�'Q���n̥h������N�c8*�ہ'�|l�]����9��@D�QE:%��`I����DT��:$�H<��'D!Rt� �v�آR�hE���Y�<fŁ:h;0l�-������	z̓Co�豍��Ă�W�|�Q����j�*D��y�"�0�n$A�-?�P1��I�y�ě?���Ơ$y�(5q� �y
� �X��g�ε�b'�
?�����"O&$�U2T��U�`fS�Ĕ�+�"O�-� EϘ$��9��<B��̪�"O���t�"{n�y�RM�&�py1"O��C�BF�]TR�:E�K���"O��@��'E���@r�S�4��eX7"OZ7��͙��I���w"O��k�7`��`�w��'Ϻ��"O<�L�<��A�F&qm� �"O"�ϓ� E���ĦOi��Q�"Oz����'j�S�4M�فu"Oj@{����N]#f�0(� � "O=�����@�&M&�ɷ/n.!�
*��)3�fFT�Z�M^�]'!�䛪su�@E�F�q0�cW�$,!�� .��0TmM#z�ޠ��_�}�!����� �5�Ġ��K1�!򄒷 uH�9TjK*��l��D�T�!�$�k!2ujt�R>G�"h��C	�y�!��D��A2���s�,y&�Py�!���yX�ka�t�V������:�!�D�<�A��#۾��ѥ0�!�d
�mR�銊~�Yq���$�!��ҿ B�ծ[���%c�?+!�T5 �����ٱv؄�)��({*!�d0 4���ڃϐ�BՊݪ!�DI������m�.��\���_"!�\d�T�9$cB�7D�5�t�'�!�ċ�a�^H�S'���7��)d�!�$Ŧm~m�P�;��o�/h�!��W�$��q
��|	�H27�&^e!�dQ��	�!��{�ج�㉮l>!�$��k6U2��P>�L�Q�� i�!�SH���N_+sǞ�JZ�����'����}w�g���>r���'`L(�UI,�yq���@9Fl��'�l�9u����U�1lL1�p�
�'Ⱦx�aM[���Q�d*#h�h�'\�z���(�ǀ��%�\��"OB�B����<Fj�J�G�r���x"O���B���_l-�1��X�J "O�s�G��0Na�D��B�����"Oɒ�Z>s���+K/q��Y�2"O> 3�0��z�i��q� ��4"O��Q>���wB�3h��1b�"O
��5�3�e�eAQ�,�"�i�"Oр�ҜJOԳ$���($�3"O���f^8;��q�6��(f��z�"O��.��1RV�5S�A��"O�X�s����\2L	f#X���"O20ؖ�˗�)����"#02V"O0��������%i��8u�Έ�yr��1685HPM��2z��/U��y��E���ɨe��
f.�6B��yb���dyޜ	`��{]����y��z�NDBkAd�  ���M�y¬�VL��T�\!�P �y��N$Q�4(�&��Y���u�%�y��PM`	PeA k�)����y�`CWm�ٺ4��+�h��M�8�y��Ԥ$z6؃$�!2��P�;�y-L�1C�=��̂	���+���y�d ����%�L���6gX�y���#^|�e��.1:�T����y
�  
�W�or��Ĉ$>��"O�$�2_/�d%�z���g"O��+�`�0�C�Y��zc"OU�E*�L[4�(�Yl�F�xb"Oj���%��Y(�'K<j�~��"O.��`ʹ,�`K�EW� ��4�"O�,`Ǌ���7�O6��"OԩY@�B:YK<���ϰz��}A6"OrŹ���׊Brn�x����3"O��yp���?*4�1���Q���"O��	a�Z-���a��'�P<�"O�QD [��HAB {�� �P"O�A�kE9hQ���Wj�n\4(ȑ"Oj��
R�:j
����k���"O����,�F��8r'����ģ�"O~ [��s8%���Ԍj@p�(�"O>�8D�g��p;�A7[*.��w"O�8�s���g|�Gc�,>.��"O��0���	��D�S���%Ѥ"O&����E�4�J�``��*F%�ģ�"O��{"�-r��u��X4~B�ؠ"O4]�2��L�q�Ñ5�n3�"O& %9E���Bc�0�J�+�"Of����  ���ѩ{*�1��"OL�p ��U��؆�̩g7�X�"O��9& ��iHd�`�E� �����"OЉ��0l�n��ĎR5��9��"O���PV��e�#g�N,cU"OȁI�i�2�x���jvnp��"O���� ��1g�Q޸j&����)D����MX�3w��ߌ$����`;D�Y-�e�$|���"d��aV�%D�@�FE��]Z� zAf �;���z�"D��y�n�:a�e(h��e# D������a�Ш�"��?���	>D���Q�C":�@��'�tQ�E&D��)fh΄]��u
�Ď7x�����b#D��s�m�c���tD��d��%���?D�L�W�.<랑3�#4ٜ�i#c<D��A����Kva
mк9}��3�h6D�l���2K�$����oM�A�6D�0��
�qIf��H��~o�M��i3D��æ	��oڸ��v��c����1D�PS�IR�ը��`l�0�t=�Ҋ1D��$M2|�B��d�=XV�����/D�P	�c� 2G�¢Iɠ���5+D���C�(
h��#jG�9j��T�%D�lZ���J4t����}B1�+$D�$+���Q�<�SC�S�^i|y�>D�tRT�G��-���Y�1D�8U鉋	I@I�%P�e�Y��/D�p@���N!�:R�� (�̰Z2-D�@���< ](4��$��B�ɓ	�
9��&���K�掲H�B�	�vL��1&�B�HD�ArE�E5 B�	<D�D9�'���T�� $�B�	����]�R	T�⢌�:N`NB�ɑP� Xb�1B @�`�\Z2JB䉘yT�����I0d��-� n\0:H�C�I�^K��p��̱S��APMA��C�ɛI#6틷��<��'F�Zy�B��o�|*�BK�m�nX@�E�v��B�	�[ �m2��
�ud
����%ZjB䉽g�.ݙԪՁ�}���;g�LB�)� ��U�pˊ)X� �64!va*6"O uX#�C��E05N��G
�J�"O��2��א�(�*��FO*5"O��x�����ū�0NJ���b"O�=#S)N�f��cpØ.VBQ"OT=jc(λ.�ZL�q(
gCyCS"Oء�#.P%*�>m�SI�	^��p�"Ob,�'�ݔ%�v!�Ce�Db�0z"OB	#�CB�V������I�bx�P""O�(@b��j�2)�HU3Cv��B"O��1"��|Y�a[H�(WF�Q�"OZ��F(Y;����f�5۔�q�"O�\�Ή6B�	��&χa��p"Oz�j�����j���*:�RG"O�4ڳa��a,�*����n 
v"OB`I���T�H�"7+у<����B"O�:��Ȃ6�Z�r)�/G���0"O�GN��yx��kN ?X+�)+Q"O��Ãē�s�	&�+*��KR"O��F4l{t�jo569�"OL�Y��,��gor����ÿ�y�˓�9l�8'M �n�z�Æn˰�y�J)_Į�ƍ�a;y6-Һ�y@  ��Yj�G�D�N�s�����y��)��̛��Ŧ;�đʗH9�y�KY�S�N�I�IBt�0� ��y2">'`$�� ��f��E�gP��y��=R�����Q�ZA�Y� ���y�M��Jՠ�lO�	<�i#SE���yR+��)���� �{f�
3�D �y�c@4 ��pM͋x7*�S��(�y��*aX�I�hz����B� �yr�O�H�p��@�Ŧ�>�
sEA�<�rDl�t� (H:��8��Ef�<��*V_�	P���m��1�Śc�<��P�Rv���b�	^��r.�c�<���k[��ɡEE�w���qB�v�<�`J��z�=�$��@%���J�<a�`O+*p����1|$����NG�<���: ��G�zs���e�E�<�7OK�l��GF6pPx��#�V�<�$i��%�6��B��z�>}��^P�'�����*nz��a�k��Yf�`�Jպ![!��K2�كf��?Oj�ys(N;qX!�$�6k3��J�@On�fļU6!��M�{@d#���6l r�*aē�W�!�DA�{����^�4��1��8N�!�P�zD��:b�;LH1a��}�!��3���ZDnϭkSRa�E 	U�!򄈿�B�bʉ~��`��b�7i!��7��X)v� �V ��!Ϩ<�!�DLh���G��N�9�Fށ_!��\�8�ر�O�0:�j������b�!�38��a[��ռ !|с�9
!�dU����h�X�$Nuj�B^�!��Q���kb���i�P�a �ͨS!�$�@��(��P'о��G�N}.!��9z��c�E;z�8��e�.O!�$	�M^�@�蒩�2	��$�c1!�Ě8<�L��e�A�s��$�3�!�DV�U��՘D�!q�@�A�w�!�d�R����OU�DWtih�A��x�!�dZ�S�����Gv5�a�$<j!�.t��Hh!�ȉTֱЀ�\� K!�� �\3go�5V�4q�� ,a�nX5"O�1`���D�� ;,	��"Ot$ڥ�W_:��"�!k.84�s"O��cw�2P�6y�G�N�zL�P"O:�ش��6y�8�� ��p����U"O(鳥cĂ8�f��d/Ν��@�"O.Xe�_�K ec'͢Ag2{F"O ����8��Ѡ%ԉb�^, t"O�h�@dU����ADǑ7�Q
�"O���ntlE/dXM���G.&!�d).]�i�H��/��5rr'��z��VH�
VNאy_��U���y�i��b`\�#�\��T�;b/ݗr�*U�ȓZ�q�C	���Cf�s�p����dA��>����2<p�ȓ��"�� ]#p#F
����ȓ#��I����/yj��I.U�NɄ�E�	Ӆ`��fd�eC� -��8rEX� 
rږD��l
�?2���Z��Ԋ��zA��8��9(X<)��}���Z��]�{�4h0CP,L�NՇ�Li���5��/vXD�C!_��RԇȓV%�brmҩ%n�ͱ�H,xOJ��l0h�%ؙ3W�!P��$���ȓe�������r��%��B�=��(�N��U�\x|�k��$V��5��@��!��І���' ӻU�ʑ��A&q	�&̘ ;��3`(�r���ȓCI�)�s&Ŏ��LR��'uY��ȓ+~�k���?m�*I� @M)x�d���i�9rb��J1н�-�,c���j�c#�&\Mʼ�o�~4I��]1@xa5�@q��!g!8b�x��/劈�B�J�d�F 	8[[��ȓ|�D� ��'0]L�:u��6tC�Y��w�X�Af��.���P.�X}ʝ��q�x �lG��<����1t4������YI�
;`^$P&bU�Lv��ȓ]g.���5�n��0Z��0��ȓS+��ЕKνp��%Q�L�OC���6<�)2u\>fc��� �Ŋ����X��u��Qt%�ā1FJ���2�9s�
�*|��0KϬO�}�ȓ"�Ș��d�c���KDEc�� �'����`ʴ=�8AԌC� X��'wP%���B!B!@�cSl�)7͚��'U��A�{9�RB�,��8��'�2��LPRg�hY�g���Ɉ�'��i�m�6�n� r'� ��u��'5�z�Z�����S�
�NШ�'�D%C�.��k-�`h2��NH��
�'̪��n �ij��^����H
�'Z�)H�&�: ��\{�� ��-��'ax�a�4: �fn�*b�<P��'����C�9&Gt��@A��.6RՋ�'�N���h�N<�@���'OZș
�'8��і'ѫOb�����30ChI
�'z�$l�9ED�W],�d	:�'���Zb��:I��m���	W``���'6��6I�P2#��]D���'Հx��+"�DҒ�S
gd|��'|H-c%H%u�x!@Rb�&Z� ܚ�'w���v���Ҡ��(��a�'�<3@`�Y� ��V#n�
��� �6��^�`�jT����"O�yc���K�X���&�9���z�"O,H��#�	�e�<Gu���E"OȰ�G�	\�I�F��l
e�W"O���� �Hj�Ѳ%	�|��"O$Dr*jT�3�J�"�~�P"O����Ć �%�t
˾}Fq��"O���=l�:x�J�k��$�"O4�:��OӾ��Gd�ex�
�"O��s��S"�RyG$�D&�`�"O��*V֝M'���7d&K�"O��9P��h&�`B3��'%�h���"O��x��	l�����~��<�"O�	;���x.�Z ��6��	��"O��$޿-� �2��e��@A"OXͻ&
?.�Z��ªr��l��"Od�1�Y%�:�R��N7�T9 B"O&�w�����*�^�<hG"O�%S�Kҋ���q��X1�\H9�"OI�A�E!+�񡴋͋q�Z	3�"O����ӽ\�ѻqjI#3�܌�"O��ٰ.W�xr�x���\�4}1�"O���iB�9��U�L�D��9j�"O5�v"ѽ5���� ,�2D�()�"O���/N�]��$)'�Ġ���Q"O"d�¡ߜZHx8A�.�F�R9AW"O��"�O� ���s�ګ!�Ԕ�"OTQ0�$�Y��JF�u�8Is"O�����Ϫ+^hQ�C�I���"O@I�Q�Z>N��V%[�e��EbQ"O1��ǌ�Ak���Ɔ?>���"O� �a��%hn,�B�I"���"OƄ�`�$y8�ԙ���S9���A"O��)� P,D�x ��F;�Ƞ`�"O�z�(V�b��#�(S|�P0�"O�*@�P(n� ��%Z6!���2�"O��Y�G���BEʇw\�|�p"O�cङ�$p���	�m
�K�"O��`Ë[z�Y�����.���"O�iB`�	V�@�pBa�3�̀�3"O&�P�Ǉ1���
T7e
6%�2"O�K3
D���y��ɳ�FD"O�9�cW�h�բ��U C���E"Ob ���9=±�c�ل|"O`��G�I>`i���R���{#"O���@�;_�V
�l�1�T}H�"Ox0�0�2}����&!Ŵ���F"On��2�B##+|8(�H�E���2"OTH�gE
D��m�7�ԻR���R"O�LJ����J1lZ�ud�"OPEbRK�"tU��]�EEr Z�"O�(ǈ��l����j]<0���"O����)H�ęF
�>�Ԁ!c"Or�KC���"5�Qj���ҍa�"O80P�M381F�3�8�Π�s"O�̱S�A���JY$h�b��"O:��aHɽ:�xLb1�W6o�)�V"OliA�;��A���!n�Ό�A"O�Q�W%�GP�,�7Ş]���c"O�Dy3m��2�xM9���詁�"O��KǡC9{�|!3bE1h2��"O�as��U�()zƀ�H��$JU"O�yj�$C�`׮��&-��"O:�q���&��"ޠ#���( �'�1O� ����6�T�˙'k���Qg"OR8��jk����c���Gt �0�"OL�2��L�lQ����5xe����"O���v��4(�@qx�η0Z��z�"O�9��&K���#�=#=�lЂ"O�pq�����+ k,���q!�$��`bX|#Ć�<_�)!CŞ�_m�}2���Zccߚ1����c�w�R�E(/D�L���A�����,O�6�pU�g�+D���w���h"H��F���o+2YY��6D�8"�-�:F�źb&��@���c�5LO��d	�'�'%��W�V�9��c�!�]'E4nԙ�$�-Lٰ��дj���M��(��8S'"_�Q耕�6���M@�9D��:�O@(�Vd�w�\����v�5D������+�l���Kݽyj�\�7$5�O��I��|\QAAD�Q�I��L���`C�I�^�Z�#��[�Xj�FC�	5 z�˥�̪=`�az�S09NB��Q�ƼPG=�v�(�
E=4B�	0k�df�Տ.�AS����zNC�	�a���A-	 L�M(�B�	 J! �kT�=Onu�ը�@�B䉜i��YYg�кp�La���$~(C�		!�����@�8wB0�r ��`C��Eˮ���N�0�
��5@
;xR�C�I4��jUd֑=���;���P��C�Ɉ����f�UhA�� ƅW����'�	�>�vD
$%�1���Q�.�G,~B�I"*7����F��P��2��
�C��7P!@I�a�8)6Ԥ��.�4A�C�I*�<�p΋�M
b��M�%ɢC�I�!'����ܮ|:��Xp��6�8B��7D�6���۩Ma��*���JYJC��(3�H�HcO�o������YB��gsh��'�थ���+y�B�	#0o�� �A7WI�E�"���D��C�I(K�D�B��Q%g�ɀ�J�	g0��h��p(��եL�L��؀B��'0D����k��T�l#�%W�|��P�C;D��a�t>&T��e3�a��.5D�X"uc��?Q~��S�qw&��^p�<��T>u�f��X��m�K�	V*l0��1D��ӆ�R�
��B�!,B��1��hO?��&����F ��A.�!��Bi!�Əo����A�C;g�$4H�Ywh!��_P۶\�W��E��21?HS�|"�x(�EO.��%�
v+T�3�L�	ϸ'�<#=%?�H�ڶ#�,�spd�0 Ԏ̣ե.D������/g"�D˥n�e�v<�#�1D�hh�*@�M:�,����P�(#�g0D�8ڴ�%���ٶ�K:z�F�أ�1D��BA��P(����F�T)/D�X�F'��\{B��p���Bܙf3D�(�i��$�{g#M�l�
3D�,q�fC�>���Վth�]�6b-D�4:p�^�iY��7W{����)D�\ԭK�X�u+�i�\pt`0��3D�,�-
�K(ā����h=N�W�-D��m�<��T8T@q��VD)D�P8b*
~��B�-y�JJ�*"D���uI�ު�{g�I�3� �`�&"D��0��U�/�Ex"�ǈ{���Ж�>D��ʷ�1mY*؂wFح=n%��� D�� h-��`�=d����0#�PS6"O6����I2�M�+��A��"O��z�FN�@ �"�m�<tﮑ�F"O�`�n�4��H���ֹ� �RG"O*��c"^8�Qq,I�� �$"O\	JP���%!��j+W'��L�P"O2$��;Z���Ћ֓ ��P�"O�1&�M&*����@� 1!"O�U#"���j�	G.k�ș!�"O�d{%�R�w��8�sct�"O������4b��v�ŤnRn�""O�ɪ�.�_����m� GX] "O��k5+O�i_�P�e��4,��"O��q�eE%�����e�,ol�YC�"O
�g�LZ�𺆆<o�d��"Oб�Q��' u94��)O�9�A"O�p)CDU�q`������0;�"O�1��>Z� �����a6&Y
�"O~m�3C^%���dUtyF��V"O�[B"N��L��$��r�93�"O �Ӕc��+���c�
��5�"O�2@eN�#���`Ç7��L��"O��[�C��Es���Vl�g� i��"O�Kb��$y>1PT�+_����"O�,1�HV"*�ʸ���҈@��A�E"O^0�.��j�ˇk�lg�I��"O���DN�\(�I�JR�+Pe��"O��-(D��X�Q&{�-8�"O�]9u�B�0�����]<:����q"O�X��
	'�h�wH̴?L���"O*���hN�N.��Ð�`/��qT"O\y�8({��;�$X�"O"u�t�M�9#�űx�  p"O��9&+¼}�ԑX��Nވir"O�eiVlN�)��<��d������"Ob�p���h��r����M�g"O,�a��<B�<`�������B"O8Q Ԥ�(���bC6X�B)�7"O|�6l�--��p�D�ܶ)�}f"O
��t�تSI�R#�� ��!���>������C��	�.��%�!�$��/��賃m���v0�%K_�L�!�d�k���Cf'�^�h��S(H��!��'ot��@ ޘg�
��5'�a{!��	9*j �JP)�-_�Ε�@f%_!���<|�Ha�fȡ?¾D3$���MM!���!t|A��(�0�T,"ę+$,!�$B!�4�I��ѺU��@C���N!��8$�z�zq��,O渨���3!�$�)Q�x��&��k/J��p��=xj!�$K�G�I23C�����IV� �KV!�䖻z�ָ��L:N�x�k�%r�!�D�M��ⴍQg���-�Q�!��V�ƥ�n[=ae�u"��@�C�!�$��$�-��F��bF&���D�x�!��,B�^-a�: H�9p�+|H!�d�[�zA�^TcRQ���C4!��>vm�!�ա[Gx���/!���3uM\)���#м͸���;^!�$6.���5D2G��С��_!򄌍5��1L��^���@�+L!򄃺V����2
�1RH\���Q
�!��A���j�圶f�*�붭f�!�d�Y��h�2���n�Ҁ[w��# �!�� ��`���QӼ5���_B���*O�Q#�ėh�N�v),�3�'l
l���x���yU����PyJ�'�F�AUDV=�Ș��V�nʹ��'ނx:�J�'R��u9�-�$}����'�����rz��%�P���a�'�N�h��E8u2� �R/��C�]��'a��*�O�,M��X��B�Cc^���'D¨{�#U�AB��Q�-A�x0�	�'ռ��Т�A�jL�Qi�
JO����'���:GI^,7�np��6H�J�3�'W��XON�n,�������>�&ٹ�'l��C!e
�"v�`肯�.�v6"O�IZ �\&�Ne��C�9d q�r*O ���U�{;�Y�&L� ,Ո�S�'�����̄Hq��0�@�	W���p
�'�M�#�[���qb�8&|��'�l�w,� J,RD�q`(<��'`��A��~ڌ �C���L�b�'�Ȅ`�|֮�A���@��'}8����I/��U����^z��
�'����]>Z���c��U�&Y>��
�'��`#-Q����&�=��'� �X
��m°��)u*� �'�2$�S�O���j����4�'ڤ�a%�1!|h8�iVo��dr	�'ݒ-pl��
�d�Yr�N�c�FY �'趈�0�֑W5�JcZA��'�,<��-�r�1v	�U�:���']��2���a�T�U�`��4��'�h� CJ�U��!�@S���h
�'� �bO�Ѵ�`�K�L  
�'!9�����8(jK��ٓ�X��'�����]���ɢH���Xh�'�t�����Q�j(3�l��}���
�'vi�tBO*��M�bW���PQ�'�����	�x�Re�T�Z7j� �
�'�N�����,�X������p����
�'�fXKaZ�@4DEᓇn�~0��"OH�a�#Ģyhp<���P�B����"O�XsFS+.�� :���jOD��P"O�8Z�7�(���C�f1�"O������n�BP����%(�Q�"O: Fh_8" �{cb��3�,ʡ"O����g�P;���!B-lU�]x�"O4����92��c'�8<�P�Yr"O �
et������P1���S"O���!!P�J�А�#Ȇ H�{4"O&��$>挃s  ��)�"O`8PЋ_17�d�!t�׾�>eF"O��c%��]������_��q��"ODdӅb��9������N$�� "Ox�J��W�ОH�! PZ�a�"O�Q�A+��K���1dY�V"O��Ɓ�9tn����ƾO��m��"OI�v��!���FMzH��"Oj`X�D�	hY��FXNJ��s"O>|�d�P>�h�W%^�B=h�"O��%#�����1%�V�#y2�"O���M˾r2���C-8r�"O��S��*Y����B_�#' ��"O�K߀}V�QFL9,?>��"O�X:+��_pAf�'+6XF"O�D�T��B�SPE��@
��s�"O� �%�RČ�jW�4�!D�p�$�2�"O*0��Y%v���C�P/G�e�T"OZ��%B	P�B ص!Q��G*O�	!E�O^z\��E��C"� ��'�B�t�n!EZ�H����'�*A	��� 0�����#�1����'��q�NB�$��@	ՃY�0�|��'�j�
b�ʳMiX ���.�ը
�'����@�O���"o2!���'���Y	D�7��leD/&Â��'��8�p�\�!ʴQ4�R�
�P���'L�����X0De6��T�~����'^&��sF9Oe�3�% A&��'�V��_� ?p��'�5�X�'��RC��E'�eP�g�*�.��
�'w��k�[�F�LE �^�nzpI
�'Y�ɲR���x���8o�9P	�'L�(�LS�KĒ͊Ua��7
h0	�'IR�Bb�S)��C$��Y�p*	�'J�$a#��^?J`I��z2�	�',�`
Z&G���i�c�m�
��	�'��e���G�NVܙڕ�R�bxdP	�'�t%ѣ����V�`��/]��mJ�'�$��e��VFDx`Uʇ�B���'���w�P��@;V�� KN�ti�'֤��%�MuJL��5ݔ@��k
�'��-Z��Į?��Ju�^�14��	�'�\�ѩ܅%-���o�9%\ u��'�:q���
	" a�#�43Hmq�'2x�d�?-m2C�
9�`)�'���Y⫓��ܠb��2͈H+�'�:+ �1�����GŨ�$qK�'���7�҃.8���_�q�Ȋ�'��1�sP�����&b�+g (���'��9��ׅK䈁���Rd�Ѐ
�'�c"�!Gz�L�UlI�O����	�'�ڡ�k5�NY4k
I憤��'隘RB⏡o��,�D�Ƨ:���'�0�!���
�4I��5:D����'%F�3��"�J�!��4UtY��'�dE��ET�+D�T!�>jk	�'���5�;bF��0�M(3��	�'D� Y����C�Tp"-ז2�8�'��!�CJ�:!z�x��U)�fp�
�'��� Mt�t��֢Ũ �P�'N����)�3 �Jɣ��D��'-^iǧ�Q$�RF(� ���x�'��	G���y�������
��'���!��Z�~QS��v���'�xL��ҽQS����Q�jN���'�N1�a�V�t(qe��f4�x�	�'p����.�""����X������'hDA�6!��0��6�ԧ��p0�'-L�@���W����  ����'^�T*���j��b��d�'J�m(UD�.e����WX.Z�x	�'3�bu ��y�V�~�����'I�܉6��9� ���A9.�N���'��@(�׃M&�T ߗ(�6��' 
���LN����&O
x\�"�'�"��Ϟ�InVȩP� �����'�z	���c8������B��P�'�񠑧�u��C-��?Z�`
�'DԘ��U,
@LB�2fn�
��� R� '�g�>`��
�� ��"Ot�z�ϑ�G�V�Ѱ��S�^�"O��X�X,���	7�� �p�"Op9�)��a`�!ч	("����"O�̓с�\W�`���"jj$)
P"O���El�9��Ţql	4fF�z�"O���E*[?�����F39X�1"O�����2h¶Al:� bD"O�\��٦A�2 r�3�T��"Odc#&�"�(����	�I����"O��H�!�N��8%�!d't���"Ova��΃?w���8|2�"O�f�1j�NPc4J jt�q"O�\�m�7z�p�Qo�]��"O^X)r+L�p�Rq�&��8S��1�1"O��RDC��G�ԡz��̶�ł�"O�lyG/��7�Z�Mݹ"꜀K�"OR��r�J3B\yy��J?�M�@"O��*�k�%���i��<��"O209D��1����j3����"O�+��]��܈R6�ɬ* ��d"O>���Yj��,��$M�-���S"OP�V�ðZHn$�Q���Հ�"O� �f�ڃF�(p��ܝ_�x���"OF�S�~�>A���H����"O24K
�R��,��6�Ax6"O��Be(��pȩ�SMPId�$y�"O��EgD�5�����v?� AT"O��:�k�>f��@D�>pa�"Ot�B�(X*���yI�BR��Y"O9фb�B�~�9��h�xٛ4"OҵC�;F"�7n�{�*A'"O���\*#^�m�C�G/jt��1"Oy��x�Y�v�5Gh�h"O������EG�̀�jÜB`8�ڤ"O�drd� z�.\Y6�q5"O
ЙJn4<iR���>���"O؅��n�^A�Q0X�l�0a"O؂R��$��  �n\��ݠ"O��`@���8At4��l��(
�"O�`X0�8sf<Ys��~K<��6"O��b6�	�bW�p�0�^�"1�)�D"O"�r�B��DNإ�5���8(��"OP0B,Bj#��Y@��D"O�a)�>H���2��~��+"OI�үϊW�8�!$�4Y��)��"Ol�p���5H�D!Se�Zk~�9�"O��4L6&O~�񗊊�=�TG"O8�x�C�:�eℯL�gQb��@"O$��qE�)I��b�C�"OPA8wl(Z.�#�� 2f��\#u"OI�P�ų4%�%��<�8���"O�A�"�ō7o��u�E�0�ę��"O	�d���(Q�6���ݶD�S"O�@�&�@�f����%���?�*�k�"O��ӱ� (dm��,��E��"O¹��Dv���򦕦%�z��A"O\%�vF�(/��Ѐ7#E�u�z��!"O���N�m��1ip"�7)V�k�"Oʀ.��q1SM�>L!��$���U`��d��xv-�(!�-G��y�)Ϧs��u�C9|����cM���y2Z18��,	�b��t�$]�ӊM�yr�]焥��%ߒ{,@*�"�1�y
� �x��:�]Y1.�2�h�S"O�y���\��AZu♚_�2i�"Ob=�A��`��6!�z�|YkV"O(u ��@�<G$�X5��10�rՑ7"O�m������-ʶ/F�^؆�bS"O���t=�Y��nհt�>AZ�"OB� -�rX�b�G��
�E"O�=I ��R�P��gM4��i"O�TuE�!mo�\
�L	�wT|`"O���D�V
/1*�i0�
@�=�"OV౔Ș�AqZ��⅒K�0�""Ov�B��*Fy>L�u���E�\��"O<�U8It�i#�ۻ("�\�T"O�2؎�_��2`�-���"O:�wFA�PEb�H���.��u�%"O`$���
����R�t� ]H�"OT�����5L���H�� �0U"O�<���E�]SJP��h��T�$m� "O�B�8��QI!�i�θR"OTQ��/=�R���U	7�¬W"O6�kP�Ai��RQ�ʢj��u��"O~y�sm�
%�z��������J�"O�l:Q�G�<
ȼ�S�Y��(��"O8Q�Wf[�5��`�p��u����"O���9_�*)ࠫ'S�uy�"Or�!�Aϴkm��K�q���c"O�9�M�V��	B�k�	wn�u�"O��X�f�yv��U*Q*AP�[s"O�0p̄{�Ż葷tiF�5"O"m�Q�ɭ.�N��e��GW��b�"O@����x��̫@B$�u"O�S���Q�&1�%K�&P5��G"O~����&
ހ}q��΍�\H��"O����.Q�c�!�ǒ����W"O6�������c(�?r���A"OR��P�	 x�2zC�ʤ05����"O6�#�I%Z���;% �>  �l��"Ol 2Fn��L1� A�ao`%i�"O0�CA���^�N��o��m=�Q!"O���GF^V�6Hs��
LI�Dc7"O��@�+�RH=	�`�/72�l9�"O8dX���O�|�놡��uL�""O扛�!�]�rT1��7�l�I�"O��b�F�m�JZW �0~H��%"OPQ⣮Ȃz�P����Ԟ@���f"O>��ψxa>��4��4��` a"O��{���#'։���%l�� 2"O�̙��*:��*���&h}�"OHD)�Qe�� ���[�4�<jt"O�V�)mR�ᐥ�Q~4I!"O��CC�N�M
*E1P(U�|�8a��"O���mڇoN2$h�'*f�x��D"OR��1�E9R��'È;�yD"OF	�f��I�|�YS��
�J��G"O����h�:TT�:���t��A3b"O�Z�ߌ6��uX�KӁM��1"O�Xy��:��@7�޽=��a�"O.y���٫c�>��7o�%�����"O����g�0!idl��֣4��|�"O,��Eԭ����$ݧH�6uh"OƄ8��Ոa98�)�MͻgT��T"O�eP�n�	#�xC3��4O�-�"O�JR�U1K\�5aت�Ҕ"O q�&�[�
��2-ҳ\��\(�"O� j-8��Ԙf��$QE�	D�ޔ@p"O(1 ���)X5�G�\����"O�I Wj	8L@d�bΡmOpK"O�e���ٜi�|a��D��r��Q"OT�)��"�"���M�4���8�"O����ҭg��� l�^e!��"OT����>C�݂p \pcl5z "OH��2	� ��9��"jƨ*�"O � G��O����#C�z9�"O��0$� {QD�)bH�-�&�Q!"O6t��M]�E��3�`1�2"O���M�*�݈�ܩw� i�F8D�8��!=1�$M
 ̕�-�+&�5D�|�Ɛ�K�f���	XXĨ�g/D��9AKĮ3�z3(��-�ā�g+D��p���p>5c�C��=�!�Dȧ:<L�W+�$z��(V�
/!��H�9	��֖!z�!Æ�.)!�D�����&JEC�|��Κ-]!��P�Urc�Z�iDt�Sr'�7�!�$�BTT�Z���o=��Q���s�!�	
��4#���\�����-�!���c1�X7ď�XڬZ����)!� )�,;��F,HUkTAV�
�!�$)vVx8��f�_L:��d/L�Kg!�d�%n�ʡ9''Z���+�)g!�dB8�p�E�{�����/Z3!���eaD�[�J�@a$�(	̽-%!��#�p��D#�"%0䋴�֕F!!�$��P�ꑘ��8#�؈���9U�!�$N�o���S�HV����A�;!��
&���:��I�5�ڹK�嘈'!��ҹ0�� ��	�2XSCKL�!�d��Z�Ty�j�d�X�0 ���V�!�$�x�|�yA-��D���E�_{!�E� H4{g#��n�f�+Q�!�D��n�H���L�;}k�m�E����!�d�?UN�Pg��\M(����Y#!��ڗ"�����.�����s!��&ud����Ǝ�E����v�O�5�!���s*�`���R1Q8��b.�.�!�d�	U�E��JW���s-۔K�!�A6V4T}�dܦiBNԒ��Ysi!�D��/>8K� ٬r��y#A���fM!�d�*at2P� @�7?i|�ئHؽc�!�D��cC:����
Q8�d`D���!�̦]���S�B#2��P� Q�!�$��d-���5��<�5E�nX!�d��H[���c2�9*�N.W�!��N��@�����r4r�#߸�!��%2�.���I6z��l�vCb�!�r�,m�q�_=>��T��U�V�!�D�+{FPe!	Q+�t=�g�εu!�D�1O����J>���:�*�Lm!�$�$��H�6lZ' �>�a�H�r`!�D6ْ����>8���֘I!��N�fW��T���>�2<�VL��o5!�䚐l�^��nX<e�,���Jψ5!�D��v�R�3�b\�2a�@׋Fw!��;.ιJ�)Ǽ4�6H�Cf�c�!�ĝGk�����co��9��R�a�!�IY0�%�`KwӜ���� %DC䉉c'���M�,�x!�3G�<O��B�	)} �\{DG���L�z�m
�^TB�)� �%�M��*<�)�9DN�: "Oڜ`��]�{��ؓ�� 9<.��"O�cK˻ry�<�6�bE�);u"O�(F�5}��rQ�K�H&2��"O�)S	5�*=Z�d�F1��4"OTH��D�:8bL8����YD��0�"Or �V��U`ؙ	R/�xU���"O���$�J��d���ŮBXU2�"O�q��L�&Y=��ӄ@�*8ld�"O��pׄ������ԋM+��Y""O,���,�&��%:�.�5W�<5"O��(�f�/\L�W�ńW$�"OZ8)�ՠ|�`�a��h��\ �"O���R�8Ω� �@�s�Bŋ�"Oh�Q��P�x�`D�}�� �"O����ț�	��Z �	~�$�k�"O0�0pӜ6pЙ��<Rą�0"O�Le��"]��h4�	�_�0�"O
���j1��
�gE-2P�"O��â�5Qt�y���T��W"O
�@�o�$���h$�.��j�"OPɪ@��1G͂��4�ʄ��"O~�(g��!BѴ��
��p�ۀ"OE�%��61��Ɏ��@59�"O@9�	<C6��1G�\3S��蓔"O" 	�OU3q�TI�;����P"Oʉ7$Ry�,��U�D��"O~}z1lZ�"~����)43*�5"O��R0�߫oN9�0%߳*d���"OFt�שհ=����cѸb �#3"OYA��0/}����Z8I�R"O� ��T?0<*��Gˎ�8��0�"O�,�$Ī(Eje��ʂ�6@0r"O4R����?�^Ahr �����"O^������A�.މn�\��a"ODR�8:���-V��f%� "Oڵi��E�4z
r�	D�
4��"O0��c��mvʴB����jʌq`"O�q��N�>�0OH��jt�"O<�d�±+���)��(�����"O
|���$۾1��%�d�lE��"OY`q&��%k>��#�/N��8�T"O�K�(�8Ѿ�[7�Sd���"O��HG��*$eDk5J��*>X�"O�	��+�3s��[¨[�-60���"Oy#���g��p鶧���8��"O1��Z"��@B�aC�/"L��"OP%#�ځ1V��Y��=���K#"O$�S����Q�q�_�CV�p�"O���7�B����@F�C��X�"Ot�@F�B%�XU��T�oݒ�"O�  ��JW�x\1�qXĀP"Ot�Ro�$W�*da�ㄤB��%�w"Oڈp'�J�j��) %t�X`1�"OtY2թV*Wt�ș1BƖslli�"O0#*_�Osf�� ��O��J'"OjE�"a^�e����W�s�!��"O�٤/[36���%�`��2�"Oƨ�#ʂ�+Z��ٱ
�i/n�"O��w	3����ɺn!�"O��P
A!,�v�Р��6!�dp"O� � 	x0H���	$D�e"O�]�2kӶ:?*y9�O���Qc�"OT�X"��>��
G"wЄ��"O� ��;W�ڿ:T��s�HB;MЀAd"O���-q���J�Όfì���'�0H��Jr�3��!Y�l�C�'>v�q@�W�Jh���\���0�'Xٹ����r���A�B�)�r��'�n���+�R��q��L�N�P�'_�D��Q�WOx��#�Dd��y�'�Рk��N*�E�2�ȳ;���	�'�8\ط��	h ��P��/G�ꀢ�'�6<�����~đ񧛆F���'b@��H�@�Q����G�l|��'��0З`�6�����A�H@��'���@(�*b�)�B�ê,�Z���'ZM�� 5��}��C n���
�'�F��-�m: #A�ތk��4[
�'����D��ڲ%� ���d�r�{�'�A�!�ٺZd�uh��+A�p��'�Z�]dN��6B�"�)�'.�!���L�
L��&NS�l��l��'C$�`d�\a��؀��N��U3�'3���hL2�5@0�� |���
�'�z��� �
���,�)���ʓ������
U ��$��-9�ȓ8ZE[����T�*   �>.�̈́�z����I>��c$I6 #���e0�U�q(�R�z��w��$��(�j��R'[�_���1ӡK�$�ȓD�t�iv�
g�i���Ϳ�B��ȓ'��2�W�$��� �ȿ{<\q��&��0�S�ء5>�%�g��:"�HՇȓ`�H�����H����GS4_@LՅȓ(XQ����d`�۲�h]�ȓ~Z�&�"fx[RϜ-����ȓ�����H,��F'�t�����td&����<,B�dK�1��&5�b�K�}�0�H#���^h��ȓ��h��Ѡ�21�oG�N�p ��qdJL[�� �t�S�&��犸�ȓl(�#LOݼ,(l�.3Aj���=�����8 x����)IpЅ�[�l�7H���V�p��+4~5��*T�n�~����["o_,�ȓXx��_7�j ڕGW��=��#%|���#E�8���斎uఄȓ6��P1H��[���ɶ�U�2&�-�����ӧ�-R��ˠ�t	�%�ȓV}����ݛY��|s���f��X�ȓo�$��L�9l5c%��!1��ćȓK.�A0'�(5���0� �9`���ȓ"��l��9;��p8V
 0.�*%�ȓ�إ��Nٚ*UT顷░/��ȓ{N%�� �4/�ly� �9�r��$ޜ�7jnA(I��1O���D¤}���'��EP��.*��y�ȓl���@��_t0 �bN�"m�ȓD#l�� �qF���ŏ6h���ȓ\��l�ª�4IvP��Ā�]���LZ�s�/ķh�&挌I��܄�%�T(Ӄ�*RN*deB]rxԄ�+�ʐ5(�;k��!%N��f������э?C�D8CeG|_����&|��r��R5?s�a
�@	�I&|�ȓ[$�%F���p�Ɲ�4�
a�ȓS�8`�藞'X� ��Z5(l�P��S�? �i �«'㌕x&!ߙ!��Pj""Ov!V���Й�Ҁ 4q�\�B"OZًUdP/�b{����wh8kc"O�	J�ƙ&B"2l����)W⩊P"O���Pl�3���;�H*6$�F"O\AJ"��f�@���#�*���"ON 3A�X0B��+�bQlߠH��"O*H�Ib�f@B���$?�b�I�"O$�#�%ڱE�z��qK-��}r�"O��)g��&�v3ri�!�41�"O0-�Q��# � ��1�M�K���"O�X���-�dibGf����-=D���BLJ<��(a�i���1-=D�xᒟ/o��)P%&!���U�.D�d�3�K��*�J���|�l1�E.D�dQ�
��!MB��H@�k>f	�eE8D�@����.���61�i3+D����M�Y��]�0��K��%D�j�A,cX�S��ژT���u%D�����=��Qڒ��_��`a�&D���Bb��9Ϫ-�$ ��!Ph��h7D���P@������R��7<rx���8D�̣bFV.wF�h���	q �)��6D�ؘU"��I����(�[��,Cpc1D�d��� :��l�ċG.%$�fK-D��#G� (xHه��o4��,,D��P�{Q�d2f傝s�Tq��f+D�PX!�/q�q�U9_)H�:tg4D�9�����`L�w��O�N��g%D����B��ԙ�`-�dmdõ
$D�d6䕍SK��@ @3���A�"D��P�[�g���xL��_�0Q�<D�8z�� +�|�v�]
r"
1��G'D�0� )�#**����n/���h��&D��jGk{����R�1+@�5 ��(D�Lԇ�(�����&��PJ1G<D���o�4pW�(�u�X�
��8�#;D�42��Q�J��f֜U:��O7D�Ȓ��������A��,��1�8D�D�Q ~U��A��|k0@T`7D�8ѱ�l< hq�@��A�SE5D�!�G�-_�" ��&1'<�=��F'D�����V tԂ���>Ԥq��.0D�c$nM��,Ds���3fyx���0D���f�1���Tj߾O�f�+.D�D{���5f���'�A�Tm���+D��8�"Z�4p�HǸQP��`B7D��3e��<+��kN�SĈ��d5D��(�� �Tx,E"̎A�$H��G2D�Tc�
G�d�¥	���Sb�O;D��c�.�j�(�lؽ^b\�D%;D��㚵N��$�ӊ�Hkf��P$D�p:'��&�R8⑫��Z@z<�F� D�Hi�͉� ��	�1��\��y%�)D�8�F[�9��E�&e��0F(D�;"OX:^�����-�)>,����K&D�hI�n�9���kˎI����%D��k��G;����
 u��iBP�-D�`Jg�i�
�J��j�΄y�E-D���ǃC� }���	DO���E�+D��y��gF`q�w�@V~�)��6D�������%M��M�t4	��]z!��;�^� ��u���!ʼ^_!�DL�s�f4*���+tcP9�rmӨS!�� Ni�!�A. ��sT
w�z� �"OPY���ª�0
�bԚc�<�` "O���C�(%Uܸc�]�|��1j�"O��k���~���`�Ab?0�
�"O�pc��@�{G0�/]>3\(��"O����Ә
��EQ"E9F\�5"O �0���6M������O��҂"O�� 6 
2���t��\��ba"Ob[`��'p�RI�B��*S�8=��"O
ݺ�*�j��E��X�$��0ӕ"OP��p��^�Ū3��5r� �[0"O~P���O�?|���GU��J�ǒE�<A���z�x)l�z���f��<f�C�g	�	AfkĽ|ڜ`I�
�{�<1��@:t��AQ�94�T)�L�w�<�^.��d���f�꼳���q�<AT�:uY+�LFb����j�<Q��$��\��L%d�2�s�"Z�<��D��ej��٠Q>�hS��l�<�w�2�
 Nm��V�j�<�����-y�\ږd\_1�Y�lL[�<��솕<^,��m��%TaF�]K�<���	H�ȲaK��iKh�҂Ga�<���_�qìbt�F�j��񐥱�!��V'�&;�L�	4�Er#`J�o8!�D�8"�
I�E����0-_ ]"!�!n�:9���-l�`d�nK� !��7qD��'�+�*��0�K�Y�!�y��9DB ����7�A��!�dϝ?�v$+́�6����Al�&Y�!�)7�4hF �*�֌�ҪǬt!�$�[}b�Ĝ�G�&MaR�8�!�D�k	�T��
"�B��ɽtS!�D+o^�Q3#jK S�h�!�N.I!�Ĕ ���#7A����}�ƏE/O�!�I z~5`�"������\��!�$M5Qε���.�G	֞�!�D׺vI�@ �#R�>�ۡ�ϡ*�!�D��j�8���NJ�m�z��F��`�!�dR7Q��$q/D"p�k� ]{�!��^fLi���ܲF����2��p!�$��GWPyq��1[� 8�ƠS!�S�Iȕr�A��~�@5sQ-�>O!�d͋0t�M����I�\Ȣ�ʪ<!�ˊjD�easj��HpaC/�A?!�8������Ύ{e*'_3?!�$�(B(���c��l,!g�}�!���/�6���)]�H¦L�!���ky:��!�('�=�CѦ=
!�'P����́�bs���!:eN!�d� 7Z��;CB�L�f�����>!�0g� ���Ǔ�:\u�F��&!� uk��@�ՖR���3��_� �!�$�,�L@k&��D^H�͋�f�!�D��o���m�^aZи"A�S�!���.�U �!߲4(ȼ:b�ɇy!򤅆Q�0r�bY�8��`�&��+b!�7�ŨAaZ7S�РZ����N!��B�v ���F�%4�i�/�?(=!�D{�<y��I<"Ѻ��g�n!�䖉@/du  �mb�(J4��N!�Dٓ3��PV�ӵw]\I�е|���'�f�Ja�?\�N�[V#6TL��'���p���:RY��o3��0	��� p�K��ɒA�z�ENL��`(��"OE����*�h���SU���b"O�8�Ƃ	Ԡ=J�B�
o>,�"Oh �0K4?֍ِbσ-;� �b"O�c@a�Qߴh u�Q.G��11"OPU�'f�=;|r��T�j�`2"O|��N�Q��j�$�'9��e�"O���悟�<���B�@�_�<�{�"O`��SNU4KLJF�öo��$��"Oƕ
'�;^�8c�єx���&"O
��1HCk/�DX�-X�G���@�"O؝P��Z��у#��><`)�"O�x��%Ȧ1�d"t$H	hش �a"O ���!�|U�f�Y�y�\�w"O��"� #)=V��p�V(jhv�S"O��F-�7l\��H�=��ݘ�"O ��5.�%��B�%_�|}��A"O�i
3�߰q�ڤ�!d�9j��?�y�mXd	I"M����
S+��yR��<^�)�@�(=����y�9�L��Տ�?kr!⑆�(�y� H7B��HV�+CT
����  �y��Dh���{e��>b�i�sb$�y��"����Y�6T�+�%���y�H$\\��ui��y,�Y�g�-�yb%��w�^|��j�xY�=S`ႁ�y҂E�_l�ZB�D\�v0*p��*�y��ӍaV�#C�'�:쁔g���yb(�9B㚱 ��2&���rBW��y�ܹXr�P�A?��0Bh�7�y�"C'��Ȕ�~���s�?�yRֻT�n�d�@�z�F�k�n]��y�/�Q�\��R��G04��bZ�y"�	I�Y�2g%D�չ�nF1�yBo��c���+6��/ 4�b����ybOT�s��\�@��n$�y��Ug�����3��8����y�dYӶ����5�xY�e�*�y� �*ӂ��ǌ]&1���qF(��y"�Խq3-� �ځz�Y�Ę-�yR��1��<���SkΤ9 ছ+�y��'DJ��q#؏k�yzg̜��y"��9��	���2!V!tDV��y"��g�0�s��7�Zı�̃��y�.�|�(� �"�>Z�H� �T(�y����8k�TP@�g�n�K����yR��HxL��A;g�D3���yR�<	F֭��JƣK�@��"C��y&Գ?�h��kT#p.^�RB����y�<i��0`�gֽ|�R 9�䐺�y�ݖ޶�q"J>���(#F�8�y�\fw"UCA�'�������yB�aKf(�L,9vL��m�yb �;dl�R`� �|{�bM��yRJA�	Q�|��[�EJ��j��
��y�@�zڐA��ɚ$2��قѡ���y2ꐫW�9ASI�(�y1`&�yrk�'5b<Ѐ����%GX�PdԾ�yB�חM�ҵ�áy\HH3Ɋ��yR�O����.ԼC#r]����y���|[��!���-�N����<�yb-��� � �t�����h��y≟�'H��1�S�l\�p�Rg���y$
"|(�@om���/��y
� ^M���)G�x)0w͘����"Or`�@⺌��O�V����"O ����F)�`��G�g°��b"O
đF�	�Ng�����^)5Lj��6"O�´,��Zw��L=j�o|�<yQ�7P�ՐS+W$����`JN�<���
&1,ԫ�( V��G�G�<�L��m��%F�4Kg��<� T�V��|qV�6.l�+�b�z�<)��G�;�
�[ӥک °�9�c(D�Ļ�Io�H���:���` 'D�$�Vd�����To��X�~%i�j?D��jQ$̔����hΠ;�͐��9D��K�l�<D<�ʇe��D�6D�LZ�G��2�|��e�Z�W��� 3D��C4n:~h$}���˗|�Ƥp�O>D�� ��X�܀�S��7(�����<D��Ye��1����rh�Hx��&;D� �'N�K�ܐĊ��@�v��u4D�(æ�\;E=�	P�
�'FX=y3�7D�x�`�W2����cʉ>��*��'D��0��w�X��)>�ɲd%D�x��� \yz�"	6I��|��5D��dM� �UP�ҭ�L����
�y�%H, �"u��¾8����Ď�	�yR�\=~�ш��FZ ��	��y���I"��3��ݺB+x����5�y�Ʉ8u�ĵ��ʲ6YT�!Ņ�-�y��$p�� 6�G�+
��H�Q��yb��"}�5-��s�:����#�y��Z�vi>2�ʔ�p��ir�\'�y҃R�R�eM�#\fv��&�
5�y2G]1�tB��@3K��\���ƌ�y�MC#V��h�ʦ=?Ј������yB�U�z�8�KV�i�r�҉�y��͟t9�}��^�="��h�oV4�yb�Sxa��Q�� =1GD��T�Z��yBo�� 7�P��J�$f�ZUhҩ�yR��1!~�3�W��6,$���yr�ݺ,�6, � �&8{����y"h��]���Zt�ƣ�֬��Ë.�yr M�fg�I3P��2�3Ѓ���y�i[�r�0�oϻ<�^ 17�8�y�oho8�D���.a0R����y2�J�4��p�%�T(ʗN�1�y2lM4R��u��^'",v؁f��y�@�cM �`IΓL�	K$�y��@-X�s�g��+;H2u�D��y"m���T)�"B�Y�jdXt-[��yr��4�~5��PYj��c���y�iF'm!(�آ͚�@
���͚�y��Ҟw� ��cKS83����@���y�K�K>ֵ�G �99X�hv�]��yr�,L�2a��i�5/Fĸ����5�y�cL�W�AH��,,���ŮJ��y��P�p1jQ{`�[,*	f���NB��y�#<%���# ]�nR@�2�K�y�l7 V�)WÑ/(�|�/]��y"�ؼ�*�;Ca�\��+�����yr&�d��������Z����y��:��!X��(Bj�$r�M
3�y��C�;|.��%�l������y�f�6TGr��,G�yԬx�N�y��@��@���Ei��
d� �y
� >-bፒ��09�L��~v>�SG"O��HTO�;)H���d��Yy�Q��"O�A��CD�(К�8���Lr� "O|D�b��%z�����8� �+P"O�8sr�B<f(��x�g�{�L���"Oj�� MP�<��'��>6�8\� "O�<�c���xD��S"C��|y�@��"O�I�ϒ+Q�*\`'aN':_p-K"Ov9`��R�1]�,hQ���l��U "O�CB��kU$ٵ��.R��'"Oh�闊E�y�Ɂ�g�T���"Oư*5�0ᄼh��܂Y��+"OB���HF�2j�.Ak�|���"O�����:I�\�t�To��� "O$�'N/&�$8����BI�g"O�*2G�7W���r�j�=�0my�"O�M�p�[T����×%?����"O:�b֠�+}N�l
`HA�@�M�"On�J��C�B��5۴A�|�NP W"OH�a5�}D�`�K]�`����v"Ou��'��z�F@3R*ΛO�*��"O�8�%F@�l��t.
�/��uW"O��Q�ćF캗��>��q3"O�{��Z�1�@�E�C�αB�"O$Iy)�#%B�Hwˊ�b1kg"O�p�AƼ8:n0Jw*[�'��q�"O���&Ϣsΐsc�:�K#"O|��AW��bQlx5��"Od��N/3րz�A�c����"O�q��BN��k0O�5j`4Z�"O�Y��A�l�^�򤎖9dT�R�"OtQ���@��:� �[�1�E"O4\q�)p  ��!��,=V@	�"O�Ia��ЋdE�tdߎm�h�8�"O�a�BB˴ 1N qg�G�@��Q�"O��)釂6������gG�Y�"OH�a����ه%�3�F�m�,B䉴�P����ޓN�E��o�& B�'E{�����K�	�B,ܻA��C�ɈHm�$�9w�#Q��a��C�7��2e䁕ư�P�
V5g�C䉧�XA�tl ����a�q�C�	m�>��W0�����ԉu~<B�	�L��	��_� 8�1@T���B��C��0i�H����%�dX��D�
�C�I�
U�ˢD�/^�^X{�`�SR�C�I�RL0��O<V��eU.��p�\B�Ɏ+��k���j�6E@@bőg�B�I=g�"d��h��i"�QFOF0��B䉆t8�
E`�bw��He� �\�jC�I"
8`��υ7���ڠH��+�C�;hG,uy$	O�l���o�e�\C䉦4�EH�h^�A�AF:�B�ɐ������Vx��v��9?�C�I7����Q'>5�$1�#c@'u�B�	Dv� ��<-N��� �jY�C��(dS��o�K��y�/�t�C�	�q@��R��<0s����-g�C�ɧF��@��˓R���)UM�=��C䉱P�\��ѷ7�fM�-̑s��C��31��[*m���(�rC�I�[�1��c����Ce�,C�	>�F��S/U�i��!���&��C�	�$ox$�d�"lάHF�D�!��C�)� �10�`R�x��Q۶g���S"O�{�Ȉ8�J�Z�A��T��	�g"O��H�ӏcr��p���m޺���"OPHAq�WG�� w��Fي8��"O��#�)V.Aرo�B�x��"O(j.v�0-P����k��#7"OxU3�/�){dyc����)�b"O\�gBF1ݐ��� K���Ti"OPp�� ��<�@�[*�csz�:�"Oz�R�G�
m;|M���[2J��Ƀ"O@ȱ�J^�}��qq��/X�ȃ"O��:��[g����F�7)�ʠXS"O����*@"y�$'�'�m*�"O�ԡgG<IE��d%ԁY||�ٰ"OFm�C�#$m2<2ծ
:q&ȡ"O$��FKT.T-�J��ǰUp�p;R"O*��b��Y��վ<^� +b"O�1*���% `6��2-�""ON4�0ECq
u@B�W�!�>}B�"O����Lޠn��А"�����}Y�"O\(�GML�j�:���IтW�8���"OR���d1U���[�!FEZ"O����X=C��;A��S�y�"O��lE#fz��IR]��	zF"O�4!t���r������Q} �� "O�<`�%M���BD\D<y�"O���N�0NK��� ��/LUI�"O
$��BK���u��"�ͨ"O���f��lW���,O@����"O<�!7gV�B��!A�C?.�Z!��"O�9���Q/yz6�ص�V�4��	��"O&9sO�y3�x�qΌw��0D"O (��M/u�`R#��0q�AF"O�Q�SmI��q�L��?�^I�Q"OF��LEL�\�KT����	!"O�-R�J$���&�{EĹ��"O�q�`%כO�>�sR���>(&���"O��I�	ɳt� �Q��K�'zi	�"Oj��EbZ����v��	T�*!�"O������a��p4���h��T"O24C�σe����d��L\RA"O�a
6l�*�����Gn�H�2"O$��q�9  P������]}����"O����-|�hy� sjD���"O�7�I�m!L���hA�9��H�"O����ӨQ8EAF/|�4�;R"O6�8-�EE001�&҅ =��!$"O�� ��,R�x�zq�'h��0"O�]	�
�D�l!R'��x
Y��"O�, ��'�4	� !�*p�"O���3�Ѫ4 ��A��2X��z@"O<�Q��q��Yّ�ʝpnhD+�"ODU�C$O-$�b�U�օ4g���"O.u�Ǫ�:�fXďhZ���"O����T�%5Xt�q�� N��"OޘөF�.����!�;��J�"O���oQ�9�цkǠg���"O���J��V������	{U�M�"O�h��nжj�(��
Q�K:f�J6"O�"�I�p���C�ʗ�?��{�"O4�s�,�3����vv�"�"O�d1�W�,�z��/$u�"O�P[u-
T��*�`0 �"O@���@.
�� ����R"O�  �³�Fk��F��`���;6"O�8��'y����եT<k��P��"O�Ȗo�� ���k�䁅n�p��"Ob@��EJ�n���4�U�C�8�
�"Ox�b7��D�|8����"d����#"O|��B�$fr5��E	+z����"O���������N	�	��+�"O*]���������R:��څ"O�EdN"�D-9@�Ya�N̓�"Ojp�fN�D$�D��8W7� 1f"O���CW�z;�tr��C/��ZC"O4��S�ܱ]zZ�f��;"I<L%"O��s�H�Nq�K�M8�Y�O���7m�I�D�J��& �@^C�<Q��s��!�E��#{:1S@��e�<en�%6��i�'������J)|�<Ye���vn�I	ņ[�Z(��ץK��hO?�{;�0i�EJ�dgBQqf��rF�C�	�,�r���X	)x��S�T��RC�IG�~uj��=*9~�
`'��b�b���/��$��E�d� }	f5���0!򄆭�YQ7!�	<��|7:kYax��I'[�4<9E��g�ҙ煌R�\C�I�1�tdq�ʗT"��8`!O�"�^����Y�L�"�b52�ʃ9q.L@�"O��vNU$a��k�i��>XFᐧ"OޥTi��2���R�H_$oF�d�G"O `��@����7�Y�a�NIR"O�@ê[��d�1���S��u���	�0|Jb�	h�輐ш�D������s�<I&N˂A�q�T]�raD��V����>�G��2��9�n�IT�ARA��O�<�E� -_������Q8��2�r�d/�S��)�JUy��w�Yx橑�\�0��V��0���<:p�˰�e�ra�ȓ+t0�"���� �3g!�D��4�ȓF=���1��0W�vM��#�2v��-q�'/Э�jҠ;��4��N(_�t\����)�t���2S�A���	?N6H̹E���Px�iK��Xա�4kxcT
^�jD~�"�'_J�K6��6i
����G a~|��.���3U^F�J���>����U�C�I�Z�]��c$��REeQ(=�#>a���[J@��WeH+$��-���
K�!��O��	RU��:��9�ǆ��i��z��%�/�.ypvl�>2~��#�UN;tB�ɮ4f��2EG�K;L=�-��O�>x�ƓfU�䛒/�d�nY
��X�T���� �M��y��ӊ ' %��+�s�b�3�b̉�yR�*bQs7M�;6�\x��b�
�0<���$��H�TlK�a\fxT$��y~!�J�$���b���)$���5� �HaxB�ɵr(e��J�Y�x��ݖt�"C�I�aIQ!o��v�B�X���1;F C�8AV�b1���Mml���hs��B䉫{����@M/��H�Ն�+C-*�D�>y�Z��%>���~��˴A�z	����+ �|��n ߰?��'�*<0�Mnľ�ᇪ�4H��q����M�'�%,O5i��4i(�a�{��!q�ə&�Q?y�@,\�f���GLX��� �#�O��eX^xkQf�&HT�#�c$Lh�m���y?q��d�~څMV�%kv�' T�g��i�Vd�@�'�"�i�Q>���c�FXj�C��<}2ŠcM ��-�O8xPP��/*� 0h�M3^d�b�'W�������j� x��oخt�l*��D0t��F"O�u�IMJ/ք8q.��z5TQ��xB�{��hO"��1���zJ��y���M�M B"O�]�i̖E+`i�Ul,);�|�>Ƀ˄Xwp��)g��'Πl�Gi&;@���J6�v�ד!̶�O0��@bQ�p��dbU�S��+��. ���DǕ�C2A
L�fg��60F���O����#K�S;�ybf%�#^n4mK(<iu��a�6욵Q�}�@�s�
�M��8k�{��\�d�0��g�>�`��C�yBʚ�T���۷�`�C��=��'ў�Oܼ���,?fx�3c
]�:�r�#��HO8��dg�1`�����a˔���i��$���L�p��aF�+�넠*�!�Ě-G�z���7)�YIlms�C䉮lv-���!�8@H���v1�C�<�d���G=�$٥�Z$*�B�	�nL�s���4��$2p�2o��C�ɏH��U �p
��"��$xpC�Iv��h �7/&�<r6F`C��N��PR�׋ko|�Z���+l�8C䉇`Vީ0D��#2�Vt��$�OF:B�ɥ}O�[s��W��\��A!n�C�漴�K7_ζ��@K����C�I�N���'�Y�0���*�C��M=��� L*6-NAٕDF�x�C�I�p��ݙ��F, 	baä0I�B��4����� B ��"����dB�	���Uj� �U <1: _P~C�	���p��W,&� =`���) �xC�I?���$��\ �f��`;:C䉵s��4A͝x4���ŏknC�	IԪ����O��"l���C! �B��$@��mѮ5ȍ�����B�I�� ;%#L��Y�g ,]"B�	C�b��� ��(@]:  )(�BC䉗;��`�V
�H^y��@�%vB�I$ks@`��R�y`�(�ڋoC�C��,w3�u	��r�x�HvMV�(܊C�IJߎ��h�$f�\Hd��YVC�ə=j�4�f�
����$�ҭB�@C��5Qi�d�pC7u:�f���E�C�	�|�P��ҙe�9h��	"��C�IE�<���"V�,��0��A�>B�I�YC��p���"����p\x�B䉞O��nP0�F��S�D�B�ɻ8ĉ�e��h1Vp�B-i�C�
��yQ�F�/�j�*��x��C�	-}�<��j��P>$D�s�:"��C��6�dDUm�<M�d�6��2W^C䉯iT�l{1�׾RH o;yRC�ɛ;�B�0E��~�^e[SLÈw�C�ɛˠ)���$�PA�p*���B�	�mx�����s�6티� \�C�ɟC�B��𾐊wh�UW�!HW	0T���6��h�V��ĆAZ�t��"OFt��G�9:l�1�q�۰W�jA�G"O� �f��*���y��Y���bA"O�T���\!����#Js��"O�P�%��8�`�P�-k��)f"O�	QBG^���Q!�Y�Rr���1"O�!8�\�?��Q��\�)]b̢"O:�8�Ȏ:#[F
3��<JW��*�"O��3��2���K�,�� ��P"O� �-�#\-��(�F߀P�t<��"O��x��\+�8UJ�&��+�"�"O��I^'p�d�[�E\�Sp��ht"O�m��$��	����D�IV���"O�A�ԡ���<śdٞ7���Z�"OX��ѪڻTհ9�@+@�R�,I�`"Of�a�ĝ�)cR��q���!�h�%"O@����*N��)���3H�6 ڔ"O��
�KL�b�\\:@���~��X�"O�X����iC�в4�G�!��D�p"O]cNi��9[��ٴ{�1qc"O�4�Gk,�|H�eM"�B8��"O*� U�ð`��)�����#k����"O�(�gViȮ|����Ji�ԑ"O�	�� ��g�}�P�B9Kr�$"OV1��U�Y�	��`�k���@"O=�`�6B�,�F�-��=��"O� ��a)��1+�m��\�a"OVU8u˜\?܁�u��}�h��"O|!�1嗆ʦ���B��\p��"Oj}��CJ62@~�{�a@�T�p�"O�Tj�Ė���ړ���PDR"O�Q+6��?�|�2�#
�X�H��"O��9�*ݑ2I���!��B��9�S"OUf�{$�L���9��;�"O����*η'���aUKݾc�$U"O�ѳ�/k�=[��@�"�:ݠw"OX�RE�җB�t5��˙"2�]��"Ǒb#�ۢK�A��K:X~�Q�G"OR�낄Ƈ$2���ұn~T`��"O@0C�	�|b���i��hvU�"O�Q(T���}��X��Z�[��a�"O@ڵOG.~g,�yҰt�\x*a"Or�s�욁nz`�Q k��`��a%"O8HYb�۝KF՘��ظ;�,��"O4���lã�E�#��f���"O�:�ǋ�8���5u��r�"O0s��=,\h$��+��7�2#"O�ի%�!��ajS��=)lLp"O�x0�޺pAr��BO%o=��@�"O�a���E����'.�U��@�`"O88iA �$��\˳mS�F-$`�"O�!s���&T�u����t�C��+�x�u�C7n7<�(֎�C�I�y�"���Ņ:�.	�c��>X~C�8�|E��R�j�:��͏-C$C��q��8���ō&�{q��J�C䉊,�ĩ"$��[/�؉�-֓L
�B�I�z1�`��)�p�r���CE�C�ɵ]e���{���6�׾C�	�oo������T�P�4�Z(T8�C�	�"���+e/��1%�԰Gi�%D��C�ɝ�vP���C��-`df�uͬC��h �<!��M6�d��eŉBB�ɂE���C��Qиx(�%ЌYB�I���j�"=Xz��� ��C䉵m��Ѕʃ�Lj���0W�B��1�ʥ����g��$��>nRB�I��Z(�7�]�K��T�`��i��C��W�
%�b,�9��"f!�!V.B�ɦAh��@�(3_*�BQm� B�I�WZ-z���4�PP�WP�b��C䉬)��k2dP�6c�ka/�&I}nC�	:��e�ᅛ�L��a(�"͑d0�B�)� 2�!VB��,��ճ��إw�V�+�"O`iP�BV��(<��+���e"O:JCKK�?�8�b*U�}� t�"O�`1��'����c(]FH����"O�ɘ�-û:<����'I���Q8"O��@&��x$X�q-�=,q�KP"O4]�"*Xݠ��V�@�SY<�C"O���
K����I��nMx���"O.-Su�G*B+j=�P!D� I6��'"OT]B��40��U�G�P�k=�`aW"O} S�̪O>p�B+�Q.��"F"Or��2�D6E̺y��C����A�"O�|C�.�2#f<�`�E��rlw"OH�@gڛ<��d �
��zǮ�r"O�4cI���� �*]�F���"O����u�bA�j�g4��W"O6c�N_0�\�R�Ϯ:��M��"Or�E�,dH�ƈ/�� iP"O�Ѡd@��4�F�U Q"�#@"O��;p $eWJ@��+�H�Q8�"Oиc4�ÙcN�	r*�5R%�Y��"O��#H�6i�Z<���֩;C�$ؕ"OlT&��!�V�BiĹD,�Z7"O�D�C�//�l�*p��/��9�"O2}(��(TY�5j�ŉ��R�"OX��D�SA��B*lx۱�$;�$;�'/r��"��L�O����Xo��a�ȓ V��#��p.�����]wH��Rb���4�ɫ2i�H*��̈́ȓW���XR�`��Y���s��Ʉȓ��U�V��=x����Z�g�($�����.ҬH�����
m�Іȓp�Pd�C����D�Q���ȓ;��Tص�?�(�S ��ec ��ȓޔ3������G!�d��ȓ!��@�E�Y$?�Zm�K	 !o)�ȓq��q�S��$`<)"K�SkU��)��9X��@�&%��c���4C��Є�d� �X���;b���rۯ��@$����I����o���\��e�i� (�ȓ)��tK��2%�r��W�*	�����O���O���󒅑q9�Ԡd�|R�)�SJ�^QI�H�����
�%U�C�	�4E��A$��P'|T�"ON���
2���x�k��o
́��'sў�Z��: P ��OT�#�Qs�L5D����K9X��U�-����)7D��ǯU�SF܌0�Ǖ8��5�9D�p�E��l����#Hv��9D���d	�
����/ĕ������"D��Ӥǈ�^��{��]!�p�ٗ�>�	m��ħxy�`	�-c*��%��.x�.	��X���rD��D?���F�r�v���M9�#�_�h��uP����KRPF{r�O��� t�,bXQ� �^����'4t@R�R�?��xI��F E]� ��'�,p��R�)�l�qP�E�~l��'�و \ |H�	�GgY���0!K>1�'4qOq�n�[0��9uv�m����4ܜ�
p"O�)�Acb��ȍ�cl�2� D������cVi8"C��%�b4Ȥ!D�V�^���X�� �<�8�2�*,D�|c�A!U?����^�y9ق�k�����+��1�cD�J�����	��C�)� (���՗l�Q{wF�t�t�V"O�T�5#΅��@c�ꟹ�v�0�"O����y��D����u����R"Od��F��� �vhX����b)�S��?��iQ>[zL��ό/9�8��t�R�~"�'5`U3V�Q�z���0Sl��w���x�����ofyqm(2��z$���0>�K>1ԇӂJ�Xh�!G�3m�\T#ZJyr�'7�H�i�\6��q%�#<�1���hO�h�r�	�W�&��� +)�,p0�i-��dD%�[�H�(�Z�C�S=!��0�9� �a��E"կ.t��
O�-��@ωA��u��^�\�*uK�"ODX�ӁP
V8���$P��9�"O�`Y#�ͪ
4]�ǧH�� A�"OΕ����Bok�<UZ�I2"O\`�e�<!����%�+,���b�"O>\��nC��=R�V%���A�"O��2�M��Ā,��.a��홑"O��*6�A�[�D�r�^',�jH��'��O�(I�(
�}��]�6�]�sɼ�@"Onp�ņ��QA&����,Ģ�I`"O
M`��*)T�&��2"BM��"O��&l�*���	��Ѱ,ν˅"O�I��Ɯ�����dْ��A�E"O6l�P(�*d^��
F�O�� Q�"O���.	�BT�q;��ސ!�z�w"O�@ � 5e	@E9�� �H	8�*Od�0֤[n�L�W �>i��2�'�F���!� ܮ4���2f����'j(x��F�����4$8�C�'��2��Nh��Z�^��A��'Y�����&�r��(��^F��(�'�����'��'���BӌєL�Z%b
�'�t��1�CR�D�I�
98�'�`��c�W�,���DL�������'��eʄ���y%^-���zF ��'��I���,*JQ���Q�w��is�'q����\�n~����X�|�	�')v	��O�C*�T�DA�2M�0��'҄�bG� �0��9�+ɛ=��=��'^�Y�X ^~���Í�-��U�
�'��-��Oexv5��d��&�:]I
�'����U"�����lO`��'��
1Ņ\�l�bX�f�\��
�'61�c�\�UHn����.R},Q�'������}�aS��?B�Ra�	�'l%���UӴň$�V�:��-0	�'�:�Q(	a�t�sK� aDށ��']t	� �٤T���s�U\rԱ
�'N�|���"6	�o͜Xڸ,��'��i�݃=DY�b�C9X�h�'׸H�"��*Cfr�48���9	�'I>ܸqB��4 ���1��&����'��{N�#@����Ȓ ��h{�'C�}S#�ۖ�䫵υ'�@2�'����+�400�õA�Z(k�'r�L�`�C�bE��8ROZK����'@��G� ,��`a�E.@/�<��'^�"��S#NsHH�N�8p )��'�P!J�4b����D�$J�'�����´Y�l�ם?���'GX5�WƎ,.d&=P��4K���)�'*䌙�%6�&�Y�-�F����� �$�W��v8�P)��&R)�"Om��O�p�L���k�##O�})S"O`�����vmR����ÖCD���"O\�jW�O�tdL�h�"�%��qq"Or�&jͫl@I:�ɘ~ژS"OV��<})�4�,�1|��	&"OUJq�O�9x���M�=i�"���"O�Z�k��Jޖ@�eɜd����C"O�<�� S29uf���G�xD�B"O � �t*.$9�a�~.��V"O<������<$�Qf[�
_(��"O���"'�{ɘ�;s%�)R�V�'"OH	��V"�>e9�i )s�"l�w"O�m�T��Tf�kwȀ�W\�Cb"O���)�j�����gSB�y@�"O:tÃ��IiN1i���:}�&!Y�"Olx�"�(|�1��ҋ]]^�a�"OȽ�%]S��� �CI$��"O��p��ծ����1b�oFj��%"O84C�
��"���:3� 1�,}�"O�9î[�b�� -D0������yr��1$�z,��A���q��b�.�y�h�j�=ʧ���%#U-���y�gN����X�>��Hd�N��y�S�Zf�$��T&l014�
7�y ��N�rggY�@�� S�yB�Ш �4KP��wW$@"����y�O��k�����[5i1��
����y�L˾{�x̘�NT�:I����y�#/�Vh:��T��*Qc5����y��%qp�����/"ql�Y�+�yB-7s.��/�|^
G
�yY+�
86��J���5ߤ�y�m���\ 'Ö���\�4o��yr�� ]���jG�eTk�
��y���K�l p���{ TY���R�y���3%��i$�J�(D`,Q0�	�y��^�:��E��͜O��C�� �yr�>��ܸ���(:��zF�ݡ�y����9�ށɅ�b&��0���y�AŻd�L�3�M�Y,��8P��,�y�A� �|�p��AΊ�)��R�y�Ã�]Պ�`��*1��
��D$�y2����42!@ߧ>���W/��y�,���(*#g��5����(�yb�ԯSe$l��hB�:B ���G�y���8 6)sb&
�hyl��$A*�yb��;"��'�b��H2t�݌Ǹ'k:%B��t����8v,L>��^�O�(@h@��-X�d�A���I�<�@�%f�,���ue^(���Mi�<6S ,�mi@M@�IG��k�<���	�=e��ǃ;>����P�����V�HU�)#��<[����D�� ��"B >[��J� �|��n:� Q��3W������;O@.���ɀ��a�����HY2Y�B��ȓ�F��0��z��!�JȰ?X4�ȓ'oܕ#�*H�y,����'��g��m�ȓ\%)��'B#@ƖY!
A��ȓ)=6�*kǄl]�]��aC�
h�]�ȓ8�|Sਕ�;�5Ȑe،�� ���ŧ���uY�
"�*h�ȓRZ�p4m�%b ��O[g5D���O��&�I��>�6ǀA{�Յ�S�? �\�;�<�Q�F>-�y�'"O�53$�(�)f��4�y��UB��6�����i�% ��ȓ^��ٓ��q�p@����-�v���J�h,�E-�H���+Q;@��f��)�F-��jζ���χ�m�m��E�f�A� R��lzt��X�D���ڼ� t���4T2��ۺr:��K��!��:a��)���¶/=R��ȓ}vT|�b�I4g��AV	I�d���q����D�ɴD��b�B�*~���Q�Ik%�³:�|�h[>x���ȓ
V�f���06��` �-o�$؄����JG�I�E��e���Rm
~��ȓx�`�m^+6��pIdk�'i�@��3D�X�6^����"@�8�ч�q]��뵏�*��
`͟��(��ȓ_�|���ȁH�P��S$/=���k�u1���(�<#����X��/3�œ��a�XS'�b�� -�P��N^"5�*��cLX�k�`x�ȓnÎ� ��c�ȣbbK>��Ņȓf<43K�[���p�˅C:���eZ�;������ӡ'�	s��ȓ%rJma��:��1"�P�Zp��c��#6iO�6�Ƥ�.%��B�+�hA*�(߰W����3�?aynB䉲/��85ɕ>l%�\r�o�[JB䉙K�z���H/NΈ�Q�z^B�	xH�-�Ɵ�F;ɑ!�!dB䉳D��D��޾n��  ��M�n`B��!׮ep�Q�'������
�C�ɊYf�|:5�='���+�NơS�C�	&x� %e�6Y�(2��y��C�ɒ Ov��LW�O��e�ѭ ��C��%0�(�cC�#H�q��N���C�ɪ)f����9gW,a	v&�-n*C��6�6#���"���'`@-.��B䉂\a�|ꔃ�0o�f�y��O�C䉳7V�ӳh�z6R4�Eϛ�[MC䉞d��t1S��$*}�c�h����	�3�H���'�*�c3Ƒ�h���d��5��5`��(0��`��n\��Պ ��� =.�:����O�nZ!���;(��	��J1�X�����E=1OZ��䡄G9��2��0�(�ꔫ��,i>(�go���"OB(���Ɂ<��z��,I�y����#Yؔ�soˬV��DX�*.��6]Ry����)x¤��$Ȍ�6/��Ɠ�Q`7��hĜ�����
�"�ju��tR��&�L�	��5��1��{c Ь
��h���<]O`��I�X\�����|���tfP�2^�����F�p"��Űww���3O8d�Æ�-iȨS�u�zXд�x�Ԩ9��� )�r֨
�E�Y�'3'd�P����Y2��/=��]�ȓ"i�h�d�	$���q6(�>S��!b2�s@��x��Zf����`�'��MT&1�)D����E˚0O��*��$D&&v]J7@�*L��G�J�M�RL
���&q	�ؑ�A��<�2�
M񾸲FB�e� y���BS8���j�Yj���	��G�*�"կ8��a$F�Y9�FV�T���N�]�0�3��}��DQ(A����'+<�۲k��U�XŃ'	�N��Q��3��k�Z�9��(jD�M B䉂n���Csȍ�3�q2�S�J T��hO=2��[� �$I@���yJ<YW��8 ����00r�H� *Ma؟V� Q�=�r�H�wL��&Η>0A�)�葢.?�� 7G��o�n�3C�\2�<�w��y�$�y�٤!�\�m_�'�:ݹ'�R�Dx�mRҮ�[����L�@Y�6�gx�p��,mvn$�O� �8b%ǌ�Hla�Ǩ�'�l!W�O~Hb0˛�E%�@��Gi��fG���!�$�(X.pM���	� ����u"O�YB�H$jjp	��Ժ+A@��2̙%L�d��!�� ~@���$ը)��/��&����ʌ+oP�� ǩO�H��S
#�O~�	��P]�R�o��j�t�-J�x)
uX5�Z�0����jޮ0���0<O&��CG�!��T�E���#*~m���I�6y����,��� �$�hV�QB��N�_�]×n6E�Dr�h�c�m2	�'5*���� J_>C�W8^�i:�'�&���R34(`]�#Ŝ�e9<����H\<c?�zE%
 ��8���#���G-D����=�	B7P�(J�0��K�L��a"v�%��J�.���
!�J<A�`�v�<i҇��9d;�8I$��i��,
ԣ�v�b��[�`�H5e�;T͖ ���_�/��-Е��RX��C��ܸ'�νB��u}���*z6�s��U�2$�t�a�P6��O>�z/�!y�ā*���h?V ���*W�詨ш�]������
'��CSJ�Z��vo%�m)@�i�l@.m&����	`�\A�f�����#G��Q&N'k"T�)��@�l'q��0h�B�	A����ϟX�X�f��s&�0�egh�#���t�ʍ1�,��x�P4��W�'5bYz�m� �b��WMq��靵vm0'���գC�*!|@��0i~b+c�9�O��P6�<��F/1�����P�(��	{E�P�xi����L�
�R�=��&D�zH�-�V�9��RqJY�m��y���ɛB�8�؇�߫��5�O��*�\�!� nֱ��cڏ_�*����I�-�6�4�YF�'�1Xˈ�aq��p#D�lc��O����Ě#Nt+S(�&e�8�%��p�O0�S�"ېR��L��K��V�q�'�T�w�L�����(��G�4°�E�s"T�jH�}�v$0DH"��'��'C�i��}F���mߕ|[1����Q�wJ��n��:7�4PS���lY��k�D\(Z�Θ�3#����b?\O̕(��ݝ^PrVO͘FۘĚ��'&6����0��=�E���db@m�!q>��V圮&���A�a4D��S��E9#������U�=��"0�g\ B�*!�H����GR�<#�P�1��8-����KTB�p�N� X�B�$7��|�ȓa��c! ��*}
L��.
/L�6��ȓ]��,����6�TE�w�[/u+�ɄȓP���c�fߵ23�Ƞk�*3��̄�C�݊SN��d���ۜ-�>��ȓ2:-:�ER�;g Y2%�#)h䴄�U�ܩ#G͚3E�  dрB7 ���[/$����O����J��x��?�� �C�\4Ix�	a�:����ȓ1Sҁ��L�7��|Ab��x@�\�ȓ9��Q�Ƃ? |6���J<y��p���%��<ѻ0+��j�>��fبW/��\*�L�V��DS�ɇȓ`�� rb�jp���処I�Z���&%���T�d����H%LU�A�ȓ&����F]#k��T����-��ȓd�H!e ��r&@虂�ԍf�ph�����j0枠S+Y�ĉ�B�5�ȓu�x�t��
�@e��e�2�v��ȓf/�icpg� c�l�ː��j]fa�����E�ʹ�~�K&£uq�5��|oN�T�X�2��ࣂ��pGȓ~Hb͑U C0"C���W�B�K�A�ȓC���$Ύ������G�P̄�ڊE�t`�g�$s�c�7s�`ņȓi:�+1l�<�l}�#��	oP}�ȓm���eߝ7�8h�7H������ȓz*h|�Bfm��]���w(I�ȓ)obl��%֢$�"DH��a���ȓ@�č;d턗O_�ݓf�	%B�p��N���T+I���6&]&����'�h���I�+��l	�J�p��ub�'�Ġp�S).۶<�S�I?i�&�*�'���a�	�R�����̗=�M���� ��X�8z^8��d]��h�T"O��Q�@�7E<I��$��w!�"Onx�Q�ޅWs64�$I��'p�qc'"O�%"$�<B��=*u�1AZ��c�"OF�CW�D���)GBC�M�� "O �JQ6U9
�p��#v��"O�0��ǂ�o����t�Ȝp�V"O��Z��^'���7�G>�D��"O�AxƤ�u5�4�A��Z���2"O浂�hV
1�Α���%(d,�"O����"�*��[FF���xe�4"OL�
T(S�V�ic�GZt �Z�"O}���`�|y��@�+cl~ �v"Oְ���*z6���G/��B��f"O�l3�K����g��!�Dћ@"OX-⑁N�:�+EkI>}���S"O��!*+�t�*aE�)���"OHP8��۶W���g#ɥ�hЀ�"Ob�т��?/���:�Ǩ��A�"O"-i3���E���@��ʜ$����"O8� 2Ջ"��(���"ȐT �"O�8(�,G!q\�4� %úFZ�h8�"O��H��ң��i��'?{(�CS"O}X���R��q�#DRzu"O�����>qL�����)9v���"O���Fɼr��]��c�8la�E�"O����C�P��1�sa�0��"O�ܠ���\� �;«K@���9%"O�"�f�2_!b�(�`��L�"OJ(�Ū_)1ehh�͕�ޅ+�"O�y{2䀾��]��
+o���"O����ɖ����̕��"X��"O6���`���YQE#;%`�s"Ot %�^	$��YRE�,:b"O��)UD1�kG�j���"Oj�a7�L�W��p����.��y"ON���NM��=
5C�f��xC"OLY	��Eh���2FDL5t�2l�F"OX- G�B����LB�"�܈Zt"O���s$�N`ZH��ּe��=��"O^�W�P�5XD��M��e��u�"O��h��ùm���l
G�ԕ! "O��Q���*$���4L�(V���"O9�*
�>�"��ۣ �"�b�"OLHP&�Q�-~��Q�KN�V���"O�FK'/L� 0T
T�^>�]�';��Cl�k2j�";��U�	�'Rȡ���9P�E�SI��e&��	�'.-[��L�b��4+Ģ^^E̱j	�'jd��޼2u,p9c�S�Oo�xx	�' f�h��*u���˲jP����'�U��)�&-/pH򂔦Q���`�'���:�*ك08��s1��A�vD��'mPyJ����E^��Q�IFh(�X�'"��f�3{���2K3Iw���
�'x�၁CP0K�F�(5�e�
�'"��r#��"My�|�V�� {��٫�'�H��W�Z+8'�峥Țzư"�'z*��Qc�1���һbd��"D�$StǄ�i��P�2a���T�a� D�(�^�
� a`R�F�-"6��� D� ��bǲ���ô��Sd�-z�?D� r�	#xt9���¢r����Q#;D�P�U�#`͈U\?R�X���<D�� `��7�UK�!3w���`����B"O*Tg6N���d�&Bf�6D��&����|@tE�3�Bq+�7D���t	��\P�'�)��yC�5D����i��!v��C�N ��f�1D�0 ��(s�|�X�*L�U��X��=D� )E�_,6L!���1%���n;D�P�a�,q��mq���>b=�1:��<D�ؙ��4|��Zfς�)Α�d�!D�Pc6���O
)����(�� D��K��Dl|�j鍡*V����,D�x������@C
D$̨��6D�܀�($HB�|!0���x'�A� !D��p�*N"vEt����%��A[��8D�����,�%�1ͬu�&�!�C&g���bִkζ] 4*ûC�!�$�� Ğ=PM9��!PW#ÓP�!�I�4nȹ�c�ۍA��(c�#��!��i�DX���f���!ղue!��7F����Zz�lQ�II�Tp!���~�v`��`7B5#��S!�DG�$�0S�N<9
�����	 {�!�^�r�ҩ��N���1rƛ��!�$�S�*���ܵf�:�y �U�!���y�,a&P~В'�O��!�$�
_���$��x13�[�s�!��-"g��q�ŎPjf8��HOX!��B��r$����%�F��r�!�dA�f�ܽ�����`l��!�$�JK���"NE�\��\p�g�N!�D+E��%9�#��2��JtgY�4!�$��EM����R�wPM���	!�d�	����e�>X��\y���8~�!�18����qh�`x��(-^)<�!�$�'��!PwnI�R�Z��$�Q.d�!��"f��X�g�f|�x����&!�_�i|�� ��dV޴���P�!�d	�y�T��dR'y�F �F�	�!�I$���`�$=`Z���+�*�!��&=N�K�%�1l��@K�#a!�d_;[6��{�&�J#*	�lǋVb!�D�.^�T�0��L�y"PS��T!��[�
m�U	��C��HS�J:!���	���фIٝ3��MP�ޔ+!�Ā�;*ͱWmA�w�H�P��>\!� Z�Dq�3eQ�ϔȚs��e\!�$��-���'ه�h@S�/݈v�!�DB�h� Tؓ��.��`�.�2a�!�$ΆPꤘ�@�Ȏ\�.��" �)<�!���H�f��?����� �J�!���<���ƙ J�t��!�
P�!򤋿y�Z|��D�euT�)Ʈ�1
�!�ѭHR*)��V����nʔp�!��<<�FT9���<5�y�w�,<D!�$ܧ<��b������	�f,!�d��]�� ��0n9�mZ�G]�!�$��T�Y
Q 9���Ð�V	V�!�d�b����Ҍ�g�� J<P�!�$5�0LF+y����,��?�!�$tP�2d��tٚUhx�!�d��$}ܘ16�X�FQ�7�S/j�C�I/G�$�e�^Z���"5��
��C�I�fJ���[�t0���6��C�I�?��yG�;]
�W��x#@C�)� >�٣nͻ[�0Q���_'A���"O���*B6�-����weA��"O��y�J��4U^������p<�� 1"O`A��]+!Ϻ�I7��<�Q�"O2����9Z=$��A�g��� "O�b0�4Vyf��B�0l��a"O�@Ғ���Ud�,��L��PQd"O���p�P�E��h�DJ�>ud�m
�"OLQ���Ӯ@�r�
��W�h�"O8�Ƀ	g.��j6�B�B�`R�"Oh��퍓e��8c�KQ���3"O$�ӠGɢG��"n���J$��"O�	y��ڮ���@AB}eNܰ�"Or�8 ף<�`;Q��"=^� "OJPt�p����Jz 4�@"O�����/0O��r��Q�N����"O0$��d+�4,J2�L�v'~<2�"O����0B�l�Ǯ,�\ ��"O��;�FŬ�0�!�S9Oި�"Ov4*5.������Q�g�4��"O��G"Λuq��CWɓ'~��!��"ONe㡪�;#tբ`"�V��[�"O(��,�Rx�a�¢?M�0!ل"O�����"P�F0��kH�2���0�"O�u�o��"�ri��1U�%J�"Ox���K���.[u� �y�d@�A"Oj�-@5r�>�"��*v�R	�"O���(�:*��Z�*��l��Aa�"O�eҁ�H2,"Ш�4Aޙ���;D�`C"�3#�&H���E�RYY0�7D�TǣP!e�X�����a#�+'D���p�V�4���$� v04X�8D�ܙUEE�Z#+̈B\�)(��>o�!�S:t-�9Z��8"Sj[� -�!򤅙:R��4��8���.�C�!����e�Ǣ���X9ǕF]!�dr�.����͈]�"�iu�%D�!�d�%�8� ��Ur"�ʱe�
C�!��֐�R)J�i�:)��Z�!Y�!�^���PP4��#�q	�'d0����,l��x�&*'�A�'R-�6KFx���%��E����'��\p'�]�a��a;o�5?BA�'��0�Ǉ�G�����a�!.�H���'�|�	W̓,'�VX�O��Tp�'���1�/�(i( �C#�] �'�4Xqe�R�B�~��3�l��'Gb��
 (@��� U�,(�2`�
�' $�� �F(��Q��²*����	�'2�1�'��7B�������R�p
�'ξ�ic��J~�dq4�ϑ����	�'���P`���qk��#�	*�4u��'��+c$X);��h�-ӏ�8�!�'w8�J!�K�fњ�ȗᕽN8	�	�'3��� 8>{ʉ1�Ǐ8�b��	�'6|8G�KwP�ɜ' ��Y��'lx3f�H @p��W���8+	�'7J��C�׿ �2d���_8Dd�)��'(�ػ� M�89
��A"��C��@��'5v5�r�
is�<���%>@\���'�\(��)S�+��X� 4Q����'^V�����G$@|9�Kڹ!D�T�'�
x��؂)Ԩ4� $+���'8�\�d��2CF��\�a������� \��f�B��8����΂�Q�"O^�X�H�!;\��@ӊ=֘A�A"O�xp�E\#6����&��7�>D�DxF��;q�x3ag�-
��9�t(3D�h�2K��V~Y�U�؀�޷�$1D�`@��$N���;�M;����,D�`
�@�.x�c�Fɉ�@���o*D�HP�!�s*F�z�n��dvXq���<D�\#Ў[�.3$��2I�b�.-;D��!KE�X��d�]y�#�"D�SEM��
t������Y�ѡf�"D�d���O>MBFy����.'���%k>D�<mޣS;�����
|7�t�S�Re�<y+��4$�e�FB���dh;�M3D�$�.�:vn���Ñ �*�`�.D�t�k/.|<)�V���a,�§� D�@A��:�^��l˟NH����"D�Ġc�~b��x
�N߶-�b�?D�H�́�Q ���@�� ����:D�SRM��Nn�U*�m��<�52B';D�xh�I��eZh�5��+j��@�D4D�L�$�5� bDR�^dy��)D�4)�ᓦ��"�"ԒMyN�b8D�@���xC�tq��U�Km���,D�@g�����uÒ�r?�˲�*D��@!g@2Y����ïD*u��$���&D��t
ػP��%B�	3��P!ԧ>D���G��Sp�d8���%Fiلa=D����*P�87�a���#G�H�ˣA.D�8�׆�>��� R!�,'v�A�*D�\8��=�8���tRV0�Ɗ(D�X�VdT=fԚu�a a� ,��($D��b4�Ȃ
�F�3�ݒE��顫%D�D�VA�Pzޕ(@N5J5�!�ah5D�<�W�M"c4���G�;M�^�I��,D���%Q�4����b��:>��ٷ�&D��!�j�piܼ����(W�(!@G1D�,蔠	�)��!ɇ�C-6hI���5D��ae�V�6 b����Nшw(4D�p9V._<EX�A����$b4���`2D�l�U`�`徭����V|��E*D��g��%�Dq[�g��S��XCф>D��'��H�8��^1�x�Vk:D�h#�M
>�r�!���$Xx}��;D���-��j-<�z�_ q��`A��*D����g�]8ͳ�j�(F�*�1�B&D�P�J�M��xs-��!��"%D������.�V�X0o�<8&���+$D����O&k'�=�B(�Z x�D	$D�h�/�F�����
qP�i:gi'D��ʿ,��*rgS.6�\S�%D�tS���=Ϝ���B��PY�/%D�� ��=8�^a�U�� ]��f�#D�,J���m:|�RdJ��N!J(r��%D��9`�C���HE3�b !D�4��kCԑj��#11X�aF5�I#j�HSj�=Pc�`kBN� aw �!�B����2\$�\Фf��
�R�j�I��%�M>Y�JYi>QH�'J
]�L�l��?�&-*��QE��<?�$)"��1���S�ݠt4|�V��?n��LPB��l���L9�ZQ%�"|z@�K�NZ�(6��
�������<�%ϲ`�h���KJ��qP�c�O���h�ŤP�VUB�O׽A�����4Lإ��'�v���'���(F�(��|B�I+�����w��I{�G��t������X(am��p�}���:9V�����}z�[`	�4�6��sE� }.�L�	?��9I#Oc>	��M�s���A-)3&(Vg���JX;qk�8К"C����'9"~z�g�? YEKѢ�B��M�b��	I���X��(O�O��)�ǀ׷t5��!w5&��O<aF�#�S�'6��A�%̈́3p�<U1Pd= �jt�''��Gy��� M��[�k�O=r��$��ԛ��7��<�}篑�j������BZp���KĎ��|����џ@	�J�?D�j�·J<���ħ<X�31( �u'&a��ʕ��v�p��� �DR:�^M��N�O=Z�ې��?^��\#�锂.zZ\�qoJJ�k?�IA	�':D�����5YU����mי �豆ȓ"H.,����K3J\-aB�d���2=���Ώ!�Dd�!
�jp=�ȓ̎)r-��=��Cb���[V����oq0-rViL��DN� J��B�	��T����f�t
s��@��"?Ɉ����p��p�%H�EQ���4F�X!�J��`�X��ͭy<�$p��%�!�ǥO�`(�Q+�-A�h֊��$N!�ď$m̩3��è?����X�KC!�$	��H��fE0E�)�a�C>C!�$I�hD�
�o�$I�a��ްq)!���m�mcE$M�j �Ig^@!򄓵R�|�B7AٷJ�$tzD��?u�!�%A?LKr�� :H�<¦�."�!�D��0�2t(�Q�^B����Y�G�!�d1M M�u��m�J��%�,�!�E�%w:�[�[
뒤�W�T�e�!�Ď�n�lQ�'ID6T�,�!�Ȋs�!�$�
�\��ܩA����Y�!�$H�b{j�*E+�&!�A`ڪ�!��� ]���I!� X�!�߃U�!�8�]Ӗ@�&v�( ���ԗG�!�$�,iE�Dpf@ݘyb���
�!�$[�? I�PfÎ�~)��B�-�!��/!�Q��Fؐ��C��Ts!��^��v���D�K!`��$\Z!�1����V��#4	�=���)2�!��ާ��S4�Oe^5b�ډ
�!��P,v����H"7��q1Ѐ�L�!�dK0�QV��5�jɷa�Gs!�i�VA��mU'z� ���!^�2i!�dS�(	�-�C �cŞE9���f!򤛷�f��%+��i0�ƁY=!�ř9T`��Ğ�G�聛d`-</!��K vE6I��&T�QӪ�!�سPˡ�䂢��12��k&��C��y���=I�"�k��R��NX�&lф�yR�  
H�9V�C��>��� ���y��������<�n�� ���y�N�Q/��y��8N���TNG"�y�\�Va�$��&��)�HJ��yB-�v��H ��ϘpN��'L4�y҉�� ���A�y�jU��dД�yh�&s�������8C�mc�`�;�y��=�l�����m�(���K�y_(W�z����-j^p���I��y%ż8�����gU%g�l ����yB�˝`��[em�vWȵDGK�y�#H����ě�|�4�brL�%�y2�R�?�����mƉ��`M�y�\->���JaPr���Gթ�y�oR�$�XwG�m)Z�	F��yֱ҆H�6�+�Iە16	r���y��U�_7T�`e�� ����"�-�yr"��%�hB0��.n���t,-�yr!E�rS�T)�oɅa`z�� X��y
� ��Ju ճi>|�%K�9!F\17"O򽘕	Li�iH�gň,bR�"O�����=HH9�&��D�p���"O�0"� �)أ��F�!"Ob��2�\[�\���_N|̠�"O��q �rn s��Z+NVQ��"Of�sb�P|��:�⃾k��
�"O^hHa�W67�P��W�[�fS&Q"O� 2�c�!<%���û?�<�U"O�d��mD� )��P��G*�"O6թq��;��`S���)}"�)r"OI�TL�lL( ��J&W��S#"O
��ƤUnP`�����\��8"�"Oj�Kf��l�R���ύG�r���*O��0q" ;j�"�b`˜TŢ���'���R���
4˴�p���^ۦ�9�'�^U����)�؈z�l�U P��
�'6��ϟ8=�	Z�e�|�t��
�'����$)�2�z�����,� e�	�'����P���|u�(di�	�'����jZ�g�8�S�̿��y�'�@p��r�v`h��X�Mv��'R�� _7�|=S�ϟ��F��'x��5'2g��J�BT�)��Z�'`��ǌ�X9xA�L��n�r��	�'�)��e��<憐�7(O3��ܢ	�'���UmST�!�"U�2�d̚	�'�>�f���e�h��v�6�		�'���1�S
y���Ï^�s��k�'S���CMͯH}���HA1dv~��'�d�@�l��WK"ɹ��O�`vb�'z ���74r�"�o^6�s�'a�����Mi:����լ`î���'g�Ճ��>#�j0F�B��I2�'��}�:��L"J��Z&�܃WW!��X�ȝ+���w* ���ޛF�!򄀧l�~��߀@�y80��/G�!�"e3B�З.�?RM>ٺwa�4P^!�T�)��8�`�-I4|(d�ͷ�!�D�7J������J=.-�ABH&�!��l`*lp'��(G�������P�!�$A�\���:KY97@��Q���!�D�"M(�@��胎-���/\��!�΂P�@����#��ӭ
�!��;�����X��:��0� �}�!�݁�Jh��#	��x���~�!���yF��@5��<��ۧC@�[\!�$a�`���D)  �9	7@ʛq!��F��z�F�x�뢎�%V!�DE�%�X��s!����j�*t��"O����'�s4pA�B`��M�Q�v"ODxz�.BK�N4�Vn9)�"�C�"ONܙ
M�[~��؂�� +6���"O�8ۅ4B���K�#艊�"O���3fY'P��,��X�4 �P�"O䘢 o m����g� �i"OMٖ(�wt~�s��LM�$ہ"O�UXB�)� XKW�4Q�P1j�"O�a��"��z&|A���ʻG���"O�Z�&��U�ĵ��G�<� ]� "O�	o	3L���ƶ���AG"O(�Y�E�\O]��f^�]���"O>�`$MN�g'�H�!%f[��]�"O�Yʑ�β�$8zw
y�N��"O� ��R��8(�0ɦ���JwЩ��"O`�y��H�9�z��oP�G�n�
!"O4�!勆�*밑��N��{�Z��"O��;u���$)@e���}H"Oƍ2��N:>���#c�����pt"O9��$]-�\���4o "O�[�)��z#L4�䀀�Qh�!�"O�[�Q�s�1`��!��%�"O�=�r/�$,�n��훃z�ؼ��"O�0�+K!0��|	%�)(��!p"O�="t�J��}�1���&OtH��"Oh��c�#S�
���c֟o6�5�"O�����p3��	���yNՉ�"O��T�)c�1a#�Lܑ"O���I�Z��m�&E�o��]�'"O�hf/�=TأBIM�O�$�""O�\��⓴#�����'�)"�"O�A��
�X�vǜ��\�6"O h�� ��H�aWH^���y!"Ol�˔�H�3�t"6A$plbu��"O��R�9JP�	db��yU"O��">*r���%ƌ&Hj�b"O.q�sF�KD4�вD�n0�h��"O�x�!ë@}��e��\��q��"O���Sa�3wdm�F��1��6"O���A~�Jr$�ף/�J���"O�A�ɐ�"Ȏ	� G��y���"O�קۍg��E2���#|�H�"OZ�kS)���R���aBƨ�%"O�Q�W�À�:$NF.;��!�"O��B�F&} �JV�ض[:v�r�"Od�J�C�D� �ڥ��8�(��"O���2<�|����M%����"OR�C����A�%�TW��q"OESDK֟_�4����VJ��(��"O.�3�Ԕ^���Ru��)d.
!�"O �Cը�`Z��C��V&�)�`"Op@Q3A@�v�5�]�Bk�:�'l��D�O4F݃ f�,�h���'{T����� ��,�B#�)@���'���� ���VCJ-)�����'5��{�#�)c�#�,��1�h�:�'%@����_�9�x
[%-`Q��'-*�4n� �.�3��M3��MQ�')� #夗�i�d���L�|^�j�'&���-ƇA�(��ŏy�PX�'B�|�� dMp�����wb0%"
�'�ȁr���w&����,2<q��H�'���WݮI�p]�P�]�94	@�'?�l��mJ����``G�8W\�'/����(C!�4�8���t��',���D �C"6AzĲ
��%��'���0�l%C���q���I�',`-x3G�4$����Q@5h����'qĠ�TL�	r�TjRG،]����	�'~�2�`$��H"�_�ִ0	�'���z�Ǭoe��;���1�+�G�<��<���C�6��#�@]�<Q�&S4<�@Wl���0��\�<y'O9��K��>8��T�QoDW�<	��4~�|�1����]$(h:pg\�<�"`�-<Tu2�ؔ&�fJ��T�<�� ��f���#�G��r���J�<��*	�?�y��P�k�pe�JV|�<� 25��h0k��#���70ƺ��q"Ob�Ɩ��՘���i�T8��"O*|��h�8���Z(.j)�!"OJ����]=W��� <i.�j�"OT�1"�HPp�1��J p� �e"Op|ɐ�I_J���Ӎ>,��ڀ"O��1��<&�@iR�B���!���`>.}[@�7X��K4!�%J�!�W:�D16�V�rH�c�N$T]!��D8���(w�3S�()�.;{!�$Yv۸�S��O"��S�lE�JY!�d7;Ú`���'v���q�M�.�!��]��Rƽ�����.Y, !"OީjaǤt*x��/I�Z���"O��뒤 �}c|��b���+ۖ8�"O�Ԋw�\qKp�qlFe�~)rW"O0e��ˋ1E���������"Ox����{��H3uKW�QwX]"O�ܑ��φZ��]j0+�!*b�t�p"O4�d;�
e�"햼IL�+�"O�T�CϏv 0jVL��X�$�1�	ş���E��F�i z[�M�c�/����6�T��qOl��u�� �CK(���)@Z-q�p1i��N'ת���L�
?.aCj޿nࠌi��I1��m3���3Y��ЌS�n�D@�-T�`�����$a��x%ASe|(A0�剄Sx*�$��MI�4�?ᬟ������=_�:�*�O�!V -��ƚǟ �?�O��Oƴ	q��!�"�c�
g� ���'�Z6�զ�mڳ%��X�DkFP�AGIe	����k�dS��Οh���`m�pO��#��Ѫ0�x6�W�z����X;T��1��]�e��Q�jPfZ��7������_�!�F� �v=���iJ6-I�ĞA�u�7p" !���Ĕ{`	�T���"�
l �@V.`=�\{ҥ���Ca�Oz�m��M��䈟���џ���E�� )Ν	O�~2�'U��Z���ɗ~��Q����s:����*FhQ�\��4f�6�|b��"\wlĨǋiR`A��Ur�4�0!�<!P��Xe�&�'BT�pgU�B����1�@-S���A�ɑ��B�m�:`�pSV��&BV�I�2s�N,���|��v"ą*"��3�,{��+$<$"�&�`a��(eX-[��ؑ�&B̓+�6%�� ��d�ө �U
���'�8x��0�&�:��O��ķ>�%匱�hmc C���y�f�
E���3'�?�$�t���{���+ �^�h1��
C�"�g�d�mh�	�?���{y��Pj6�}�"�J@zR�IևK�(�h�S/��y��')���_��bT)�I=E�Y!Ӭع,g^x���BZL ⇇��T%�2�H��(Ox�B���{5���HΓJ٠�`��@3Lx@��D<
����*i����4�HOH�AC�')� ��I�BГ��ܘ2j@�i�H�8RQ�6��O�ʓ�?+O�b?�j�l[4|I���ՠ兏Bs�B��?	����i+Z��h��IРD���I	�MD�i�剞d�40۴�?�I|"���6x���Μ��ա��R��?���ML>��P��+w�aG�([�L�Yt�.Ba�Sj
%�v��@B&Rp5Ey2B�.��0l8$�6T�bL&Bڡx!�\��!\�B��C"J*j�����鉽.]�����xK|��4c�(z��	R�H\pE���Z�2��'�O?��KwR �#�l�1q�p��`���E��|��f�T$n��A3�lҐ.h�����66L�h�δ��+�ٞ�M���4����-�dN�@� ��R�я`�)(׮�<�� ���&6�uoa���@ܥ�@`�6�����	O�"�˓�5 D���@���M�3o\�J�]��m��l)1AS�+���]G��+�*X��SV���`�A�ܦ�b��O*�nZ������?7��'8�&���XS�Z+�g�6n�~r��`I0랸!ob�����>61�(S7.(ʓ
��ևrӐ�?!��u�pDA�(�	�0���Xg�|��'KTP�� ���   �  �    �  �*  �2  |=  �C  J  �P  �V  ]  Lc  �i  �o  v  V|  ��  ݈   �  b�  ��  �  '�  ��  �  G�  Z�  *�  l�  ��  ��  ��  ��  ��  �  �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d�O�=�:j_�[����q��Z�|Ӂ��H�<� ���.�:�$Β,�^���\D�<�$��
c�
�sa
��A
#nC����<)��7Q�D�u$8]h�����P}�<���� U��\+ OT�%2��ŋu�<���^ʤ��H�K��U��ASr�<�7.D�(�3��5o��Ձs�I�'�ax��ӊU�$c�H��xF���"��y�Ì�I�4 #1m%��u�������0>i�/.f��4�s��4D��`	�x���'��p;E,PS�U�B��D��<�'��8�I�)NX��a��u��y�`
�&F���4'�ZpbeaX,�y� ��"�f���S�iJ����y����h`h�v�L����D1�B�ȓt�V}*vL�TD@i̯t$h�q��~�	�:zxnt125��1�y� Y`)�щ�nl�5��ޗ�O���4H�Z�F��O$B�jv^��!�d�O2�HWJ�*9]x�ꁷ����@��y/�'(c�,����:�.��r-��yr�ǲl����"6$<z@�%�y"H�I�����V�����?���hOq�XX��g
-Ph@�ݱX&"\#W"OLl;�`B�dxh�o�1^#���i�����H�S�A�4�ę�#� �aL��I���� ���2���,�tlV��s1"O^�`�퐰l��H(2"�|S�"q�'�H#=E��-�>G] }ض�^"DZ0XR���!�$	 k���4��~]&u���y�e���Z�F�:&Q�sȓ���`�(.D�h���G2� %k0iΈX���6�7�Y�ayb�QI(���*پ#�\p������hOq��l���H2����,NRZ,(d"Or�i�P��r�ʣk��
S�D�Ӧ��D-�bO�J����S#��P���D/1XZTi�x��M�rX�'Ka|�m�(f�m�H�?�P���E�y"
BQ����-�gj5��(���0>!��9E���)]�M�ҙ���t�<Ic���X(LȆ�J���v��n�<�-E
Cl �X ,��%k�uې�q�'2����O�R�1w�>'�~A+��U�ghz��1%2D�,��%�.E���*�=t��!˴���'�F=O~��h�'D(�@��nY�	�eB�.�BB剕m��H�a	Nac(-�2f�1Z�,ʓIe���ͮ}�D@8�,�#M�j�!PiGb�����j�'v������Ï�9��`��`O"R�
˓�0?gH��NPr`Ƒ��0"V��\}B�'ӛ�W��E{�'k�m(����`�(TnX�>le��I�<�emaӼ\�'J)q�>��qbR�>+�Q"O��3FA=��)�s�	%6��x��I?�XD�ԩ2S������
[���v)����0>��1V��U�z�u�v2��O�7M<�&
�&X��$/6� ��w���e��� wȞ5��x"F-}����h�1�S�̐��ē�~�b�r~2�=��'�Iٓ%^N*V!�NC�%	�|��'�<I!��Q���%���ی{B�)�I���mIb�~fp��B��i�!��C�2���b7�̦T
\T�qL]K��<�c_i�"����q�s^�$���ȓ��́F��v	hiڱ����n�s(<)�@�1P߬9�5�ыe{ح�ʗc̓�ў����c�a��L��`A"h9�"O؁�7�\��i�b-���"O��@�ܿ_LhK�!��f+@�Y�"O|�K�r.PlΛY�0�s��'�y�C�Sn����� 	���CW	�y"���,�<��4p~���Nм�y"g(g��|2�AObA�AC5^-�yBb�"��L��ȂP������
��yrNٕ h@d����*N1R<b# T��y�ߧW�b���G^�HI�)$$�y�X�A���р�8E�-��L�y�bL�GG��H���B�d<�q����y��T+@����b�Q�(���y�ḽ3�|��t�ĚL#�(E�P��yB�R���C�́)/t��dM>�y"��,���`�����=����y�({Ɇq`�g�'����K��yGֲ4��=�EB��%|�U�q�P3�y��U�yW&�3�Y����O��y" m��eh���~���LY��yr��yf��:c���4����'�y�[�+T�8��K9�*U ��_��yB�V2�8|�҃�Ho@���jJ2�yN�h^��z�o�=�:	X�˅8�y���4KǮa!�돾-މ;��W5�y�� 0��2��Z�)�&tR�]<�y��
�e�������(4������	�y
� �4+�
��T�p�b �X�?3���"O��!ҥ;MN<\`�Œ�zJ��h�"O�5㱫�|l��!��)M��R�"O�i���7���TC	.�hl��"Ot���۶4<C��(�m�*O2�1d�F\X9�Ǥ�po~lK�'�^�#U�B�R)����t6���'� �I�kJ	Nr�a�M�]���[�'�R�VL�'ᐡZ��Ԑ]����	�'#���h=�m 6�5P��'y~�rPـ�BX���y�����'�|!�ȑ�Y���νb�X���'��I�%�^-:%��H1P���j�'xՁ�`���Z���O�C)�'�&3!�G ���YQE	P�(�2�'�*칣�b�4y(���V��Ś�'B��c� 9�h�#�N/Pu���'���p��4M�ZLi��U1L/��z	�'�e�s�� cap�R`BL�)�'�\0`��(mB�Y���F6�X�'8�(����;�\I���>,���k�'Jb4����r2FX�*�e��'`�0P#�L
t_⌰��,%+����'D����V�&��4$��&P�l�'�N18��A���A�B=���	�'پ���퐴C4�!�cgK�4���'�8l Å� �l����^E��'��0�.^7?_��k��֟{ᾡ��'�V��tD�_^&]Kq�K�l�����'�$|�&c�������ת]h20��'��)qiBQ���k��R�X�DXS�'��aA�Pq���S�yZ�'���I�].t)��p�N#�^���'8���Mˇ}�l=B ��&�xx�'���F�N�\�5��������
�'����Vi JJ��BF(\����'ݪED�rɖZ��I:|A���'=��i�ƕW70���#w�"���'H�Z�@�m-@y�Z�%�J<k
�' ��� /zZqp�+]�q5��j�'�X�re��c:	�r��q�� ��':�ЇeԊe�x�b�S��c�''�ᠤ�ǣ�vX2ѯ?Wv�[�'ڹ!tO�+��!;c"�0U�j���'��̊�oα\�؁�"��Jk(��'���� �YKt����G����'�6���Ş?�h�8a�[�3�\P	
�'�Π���S���b0��!{8��	�'���,=b���)\�נ�	�'^���G�I�/�:��g��H}�l��'� [d�R
9i�����܍T@<( 
�'�a!�ە3q�0(pLz �J	�'8�H��E�v-±�nY�H�<��'�`|)�	�D�N8�ש��A�����'`���uPx��ȒP�B�+�'�nH���q$|�c��7(��'�2�K0
���*����w��d �'1��ҕCK�Nor�C� ��Y�Q��'�F}z�>��y���*S1�#�'E�Yi�8>p �R Q5~\�Ԓ�'N-�r�U�7g�`��]�I�~��'�����b�~���A
@���h�'Vy"O&�hQ�ᆗ%*Uf�k�'<�|&.��h��h�p���.�|T���� .�U(
�7�l�+�K8Gj-� "O2L�Wt`��l��6���"OL�"䇸#�b�Z�+ƕR�L(��"OH�d�O�"!	�
��|i�I�"O�<H�IAc��i�C(Z�^Y���a�'���'���'V�'�2�'c�'���c#mʊ ���h��!MlE:��'���'�2�'���'���'T��'�H	B-Ȅ��KZ�B/�����'���'��'�"�'���'��'����+/!$�٘4�	�� �'�"�'���'���'*B�'��'�<8$U��q����+T�ܥc2�'#��'x��'���'���'���'!Ti�`�;YjDi�'S�	�0�'O��'gr�'���'$��'���'A��Z�RSV-�̓d�Vш��'0��'`r�'�R�''��'�b�'>��S�;H�j�( J�"4�'
��'��'���'��'��'*w�-N��Ã��
u/N��P�'�2�'���'���'���'%��'�:��	r'�y��[9."d��'���'���'�b�'1r�'$�'�L1�P�Q�n��dX��VI�t5c�'2�'$r�'���'���'���'��2o�>��K��� �0,{��'�R�'%��'���'��'�r�'��������OW���l\��줡�'��'��'�"�'��G|�j��O��bB��E�ĸ!5.J��H�3�&�oy��'��)�3?ag�i����e�s��"hE��9�*�����ͦ��?�g?��4pC���6R_P0�� ݼ��'�i�"�ݛ���h����-.2�y��~��aB�*�[���&	8�I�r��?	+Oh�}��	�j��}�e �4�&UawC�S��F�����'�񟠭lzޥʡ&@8Cؒ�R��
+S�� @*�?9ܴ�yBZ���jM�B�vӸ�	�$Z��IdHv�Kw�&Y��I�DT���M�v�`hF{�O�B�\
B�F� �&	�3޼5y�I���yr\�|'�TJ�4,Ih��<)Į�)����!E#��cb�&��'Htʓ�?�ش�y�S��4O�2Z���m�{1nm��-;?I� v�^�r5�]a̧\�R�S]w�@��	;�>��fR�yOv!�PO�.0w����d�O?�		D���T8F�1��Jܽ=��I�M��hu~��r�(��ӵxoН���[�\`r�m�h����П�nZ��"�G٦��'��9`Q�ڱ��qA��#�bx�ℝ�	;ʄ9,��9�p�C�o�+!�e��F]Z��L>��F�z�|��L>j�Z�Z6.�W�<�VjU�{P�����
L�w�ͨo�@����R�\���!£u���Z��V"krX1��L�� Z����Ȧs�0uJR
!z�X��O l�Sgɸ)X������X�P� A�65i���7)"D8*tJ*,<���e̶( C�TaȂ	� �B�I�T Z4�Y�N����%K��0,�	&j��U������	�?m �O6�F�a��p4*A�KW.4� �i���'NAXf�'ɧ�OwTPb����b�` ;T��
$0�(�۴F��`�i���'L�O�O���@�̴�~�\=y�)Ӑwв`m�9%��X�Ik�)§�?�Ң�:nJ�٤�O�N���yeI PM�V�'���'K�yp��)��OT���x��꘍��q�u�����W6{3���|�j�I�f�f���O���ձ;��A1S��4�
�.�f���l��0��E����D�O����O�Ok�
h�r|!3��7=�x��S����'�d���'d�'���'MRV�)�w��ǃ�6xaP�l�0|n���d�%�M���?a���?1,O.���O��$�3B�nrO�t-J���d�b�X{q��O��$�O��O4˧�?��վU՛�РM�L�׹��b�eV4�q�q�i#2�'��W�p���0��'dX��I7S���G���<���xc�{�Pmjܴ�?!��?Y��?a��NG�];Ɣ������.��vl�&JP���Lv��7M�O��O�d�O�5��)�O��'U��R�X�Fuqfhϥj���H�4�?����䖿v��%>Q���?�R��Q.��=�4�nUh�뵋Ԣ�ē�?���8�A����S�TiXq�����K�.0 )5���M�)O ��`��1J����������'����-R�>��PD�H�"e�ش�?���EA����S��(�T�(0��� ��%��l%�4<�4�?���?�������)@�,��]�#��+��,�E�f*lZ
Y�q��ٟ������O��'߮qPB��+�zIy����3�D{��~�"�d�OL�d��O�&�oğ�O*2�O&	�Al�``� /R.�,��i�r�'�a�$���?����?��O�r9�f��/u�^�A%5%��x �4�?��a(<>��ǟ<��ܟ�%��X�)IX�r�Bԍo�@\�T�E�v6-�O��C,�O����O��$�Ob�D�ON��X�2�414��� �f4�  t�l���S�Iş�����'b�'���hp�.g����Ñx3pɃ�	�^���I쟌�'bcפ��)�K��=���W0�HLA0�\�4���'����OL���:���3.���QRH�uI�	,��O��d�<����ă*�R�dB���;��GZ���i���4.��=m�q��?�@ �-�<1V�S�Zd �:C���sv��+.0��'K�	ş`��m���'���5����.�~p���#���u��9���?��#L�!�N>�O?� �-�uM5gQ L(�bX�{팸RFY�<�I�O��!�	����I��SryZw(r�Ҧ����X�
^�m1b�"�4�?q�!(�<Y�� �@�Vջ��#<4y#��b��V(�>}���'>R�'��4]��'@�B�cp�M�!����E/�8���ɱ�i��ɑ$�|�c!ҧ�?�pf�1�]��P� Ң�Q'8����'p2�'�|���?�4���D�O:� �>�,0�Nٳ@;(|��%M��5��ş,�I�|����.ʧ�?��'�j�S��U��a���w�.Upߴ�?��a\����{�T��GK��D	��_�+�\9`��Bd��o�۟���:�I۟�	ΟD�'�`����*;uk:Ԣ�2�%�<JO����O*��<����?a2�Ҙ-�r�Q�U!BT <
��M�IN������K6���x��%�ʓ��4&\f��D��̬#�O9�B�	�M����b��-�̔cT%ڌv����2F�[\�L��ϔE`v-9E�& �H�[d�!Wڴ��e ���"]��!I'
h� �Ǟ�Uhx�0�рa�4aKz����6��yu&Fr�$A���azl���;5P��{E��
�۔$�4�ؓ��N:\,�C�� u:�8�$��6TT2�a�<t�8t��O��ړ�8uT�ֆ��2[$�	qi�O��dW�\�+�aM���a��U Bpt���O�S�u�\���Q�#/ֈ�EA	;i5�'�0(B��V�����ќRP�S������O�B�b2�ؾn�pت�n���m�N��U��O�doZ��M�����OT����#:5�H#c"�(7LM���|��'r�'9�	Ο|�i�EjAh�u� ؇��db�;Z �������ߴ�?���i��a
D�<�j��ߧFnX�@OC( �6-�O(��OjiE�$#��D�O���O��0X���{B�7u�a�&Y�(n�����է@�����B�w����%��Ϧ�*��i�h#LA�ONܙI�Ɵ�Eh�(��Y-q����P.峵 AOS�>aoZ�{<��I4�N���Ei{�}aChߙ�$��4<��ɚC���4�j��)�	��+�#	�&��� NH�M*�B�	���%�s!O�`�`��(��i��k>����޴�?�.O�0	���:���i�N(x�*���_�Ƚ����OL�d�O�����c��?�O����
�3!�|" Ȓ9 O(S�h� O��0
cE˼0��!*ÃL.U��#?Yw \5H7�r��l�dT{�CY�F��łtᖻ,��u�,NTr�w�ɥ	��h�1�&Qr��3c^�vҮ�0d�O����NM�Pݨ�\Z�����:)!�)�����mт\�r��p/,r�1O�d�>aʒ? ��'�b��y��Y�7�?W�h͙2�ѥTT��'��I��'NB�'� �*X0j��]�b��mZ�7-�*-��T�ߋ]���ش��x����H�1�4Ô�W�N K�Γ5�TH%Ɔ)@�.	��G�Nr��G�e�PGyb�
5�?ᐷi�6��O��e�:������(_����'�<IW�i��Ib�T��Z�AZ���*� ��M����V��Ӱ�p-��i�(z6�W�f�ʰ��O�������MKQi�>mt����?���:�*�?���N�\&�Yҵ���un���Β�?��U���{�fW�{�"���	���M��~�,��:��J�3~�3�62	<�a�>����8m
��c��k�Z�l�o��nެg�� �c��W<�ȓ��]�<0�'�ph���z<ɧ�O	��qGY�3�8���ڡ!�T���'`�}@#e�	t �Qo�$�!�i>�"��@F������ʐ(C0�_rmZ՟��	ߟ��	.ir�|����������݀Z��8���^� �Se<�М���ZDD�oڟqNzx�v���'A"�'� i:]�����Oȥ�@At���f��j�故�M����������i�$IМ'���r$*�,j�ݰ!����i'.y�P!�'�������͟"�'��	��� i�����y��H�g����˒X�.�Y�^6RΨ{�ND>5����O��'#�)2����A
\��(*�hY4!� �D$;\���ɏ'���D�O��d�O�,���?����t�N?P
&�BՄ��l�0���Wtr�"���u��4ɴ�	L���"Dm�zں�-�B��g�O4q��d+&LO	s~�CS�г"���W	ڰg*�ȡ�'���!��;7&i�6Yâc���yb��	�@t0RAW�
R���d����'�Hc�t�ƪ�M3��?iC�S+6�t��&�)CN%Ӥ��"�?��������?��O���2�K\?����8ӛ6�,�v�+��U����%�p<Q��	'2��
ac�9#��M��40��pn�P����A9�a��	�<3B�d�O��a��z��^�U>B����O/ET|x��?��������̉�o�R>�Ċ`]+M�\m0�O1nں < p�ΐ9u�*�AүV���Yy��
�E�X7��O���|�@\<�?�D��,-f�����IV�ArR��?��eRZ�;�Ð�7d���g�Τ6|HX&W?=�O�Fm��'M�b�b���K@0>E��J��S0KӐYTp�s"��&l蕪Ww�'chH(�eMFȘ`�C1f��O�1C�'�"6MZ[�C��{����v��t浨S�V*Tvc����I��T�S�? >뇧[�T�������=��dۆ�'�<7�ʦ�%��Z�$G�dJ2�\�0�,��΄=�M���?i��&���a�.��?y���?��Ӽ�ŏ'h%���.��=��U���S�V���pᢌ�mT��	H~�<�&�ɧL̠P�f��]l�`4�]�p���NG=^��%�B���}B,ʸX f�	0%�����j��U̮�r���:j[H!������v`����?I��C*b�U=��9uD7qu���}�O�R���4{
��A�}oh�ӛ�|�4_�v�|ʟʓ]��J�c�\�:�
�=�
��@
���p��?!��?�պ��d�O��C�Q<YBD�w�]K ��`��d�l�%rdN)x	��3�2��˓m��R���F�*a;�^�B���� �W0%aa�w>:J5'�'K�B�@3T� �pn�,��5��nת�?q��
����'������?9d蝌��lSb`� �?��?)	ߓ{�A{�E�I�LU��UV
E�O>�Q�i��6��<���U�6����'������m���'N��bPl�t�b�'���"�'���'��s���cUk�k�%C�7�L5�Z\H%a¯P:� a��Z6S��x�Y;��qA�{��պP�O�0���`B�F�@��,E����퍴ȈOHb��'-J7����I�z�0d)r# �2mS^,�|�'\@6�1�	��O_��A�ޞ,&�P�ϊ*C���
�'�x7�O�}A��*�FS;�JP��T� W"n�z�	�@��[�'�@EXf[�f%����rUk�'].�q�肊_)'*��K���yB�BJ���������� ��yB�A�4@^��D�� by�� �y���GD�Ʌ�P;]䁓g�H��y�%�R����bӴ,
i�iCf�<�ʶ?��x� B� �ݳ�Nb�<��JT�t7B�	U���J��!u��a�<�$��h�)�&&a����LC�<��%	�`�dܡ���?,��0�|�<�UE�M_z�B��0W�  �DL�<��ʕ������J/ �9����F�<iD�ؖ&%:����ձ6N¤�%�F�<q�#čc@mH��_�B0����k�<f� � #�*:=��T��y"b�>XNz5�C!_.����p����yR`�##J�����<=Z<990g �y��Հ[,lI���3#�V�Q��L�y�`$�,��4�F��
�����y2��l�h�
�2z��N�y���,��3�A�\��d��y"/�Eʀy�
��Ѡ�[�N�"�y���v<���A��2}ĴAi�ٖ�y�c�od���c�"o��X�1��y��\�&r�(�S���B��y����	�H`R��чL?Ԝ{�o���yF�d�D����$DB�CCJ�'�yr�ڤ��E�g �9{�oϕ�y�g	�5�ba��O�]�^�u�P"�yR/R ��8����`Φ�*�ۄ�y�-ف����V��D�8q����y�*�%s�❓�hZ1m���;Dh�1��'�� ��4y,�9� |l�4�F�N5a*�ͻ��O�(!6B�	�R~�bqE�)�B��֪��2Q+��G
V�$����O�����3?1��³V��qb�6��Ъ�E�D�<�B�u���v�|e$ #��hT ��U��>-G(=�SN2\O����!��9�lJ3>��t�v�'V�k2�	?7�H��h��fr�{V���
�)s+ٰi�<d8
�'�\hx�'ַvۖd�AA��_�6���yBI��6��@���W�b|E������R�Ý����� ��y�- &� L�7obE�f*c[ 2e
��O@�}�pPE��O*�����V!���"���hI'"O����n8B/r\�w?l�|J����?o��!�*ץ<�p��
��~塤j�!�K��X�lY
�鉰@Ҥ�w�A�l�����#�&oN,�P���3��у�(��Z׺C�)� ��!��,&b��d���1wƴjV󄜇q�ƵhR�	;��Î�)áx��(�q���?�v��R ׅ?!�DA>z���q��ˡ�EIE�S���,�\!�v����
tO,�g~��LKaSC�,(�J}����y(� l 0�ڒ�[=�����4��Èmh��k>lO��84F�e�l2#�J.����'�r��DHE?�ME(1�nԳ��\t�ҁ� �Mu�<� ��Ci�萄/ͅ?����l�'�p��	�W�g?��,�Cېي�ύ�6��Q	ȞM���3�Ov��N<&�ܭ燊�~�P �Aca$�a�����c�Q��yg@�6�I��@ܧ1�:��շ�y�i�1/FE(��L,ʠ0l�	��lJ�2T�T��s�q��|��dU>;>d@h�͟�i��D9$�'~Lqb.�A?��Gڇ�^pq����#��E�������'S��UH!ϣ^��3�+�2��ɉ�?�l���"ފa���'��!���F�iaf�5������<��bK�E8 |��GR9cY���D��P���X��'$�1�D��"��"��A��2DJ#]�4��A �<)�����Tl�i�AB�D�k��,"�k�5��%z�0�O� ��֩�Nت$FI�zp��������vAi�㔭��Ħ�T��u��SV�<f�> c".�<�`�/�V-�T��&F�6���&�e�'�y��b�461���%v�,Aܴ���� �:�x��퉤.�j����/���3	�>�h7�ɸG���	�R��DU%S�Q�t�bt�#J��j�� �k̃*d􅔧�s�l�WmV1b(B�Ǻ��L��V�1Uf����r�=�%��a
��"2�K%�ܰ�$�"ތ�'P����D�A��	�<�$c�`R�-<ՠ�`
�H���#4�{ŁD,ty*􆜸Z�;C��W�H�ÆH'��K}��;2bj��P,	n�$��<�Dh፞�l�x%J���&Z���[�-R+/t�d��#A�]D1Ӗ�d��Ӓ/�?�H���$�T�"�0ěx��Y,h�$Eze�ǽ5���ORH�'�`hc�ƀ�L����fK׾0�*	�,O2D�sË{�� D�XZ�3��O��>ɀ��Wk�hZt�ם�
�ZQA\�<q�n����DƪJ"2eBem4�k�$l����؍�a,t?�p��C�Lϊ��C�͸A��@�Ǻ'�d��<���Ы.=dO�.rrĹ�E��j{����O �p>)�.�~o�	�%N&�^aȀ��ay�C�:x�ÒSf�
�z���<;l���4GR��ܘ��ƈ
%>���d��,�<�3#!�1U�|��c��0x~A��KS+sEN�+�E.\��'�
�SU��0|��` ��hPxhha��	5%�	���6"����<�"����-u��h�`�l���&r���Vo��V ���'��i:�}r��J�5ruk8:�-1gF��WN0�F%M7���"����v��
�ўP���ۂ_L|�r��ɁW,j�y�C���C/ax�G �*>��A�Í5�@���e͌JC��?{t��[u�l�'��ͪ0�^� a`��C��<8�r���"���K�.A2A,"?�����Ŗ��W�VUI�fi>\
 ��B�rƝ{Ć�`j����$��-C.- �ۦKI6�s�;.\�'�j�	��1�^Y4�+s
��z�O��#�lw�� Z�JVtB��5�b� saF�o��䈘^/���*�*f�=��B�鎉���?!��`b(�#!(*����4B���ئ��K2i�0]�+A3d�H��eJ �:%���%?p�5D{�e	5#ш"��#O	 �� Ɋ
dܖ�O ����*�(�����f8"��IK~(�a�yB!�`�B_ճ���"1��њ#�1"��8ò
$IȪ ��+T��&Л�@l��A�����TtI_�K2�_������
�Lm�pۮi�D�"��'��S�@�+@�*�0U O�%��l�J<y2��)@&�)��R�{�I
RӤ ���6ϦAӅ��6/���aZ�c4u� ��s#fm�!��d5NCK28�33������<5z��ʘ�A��S ��C���!U����0?���[oƑ���Za�p�TN�~Yp���n�zH�I%���<	��GyR�˩Y`BIa��[\l����ȵ��?�r���3�|H �z��ju���'�Hy{�Lʗ1 1�C&NJy����I�[��<�AR�DCFq�H�k�Ԥ��'��@�1C
N���I�MC���)$a��+����|�!548��@N� ��AS,*�џ�J�b�'v�J��0��@���C�m�>�SBŦ	���H�|`+O�V[ᗀ��� �	RC��p� 0>�(��DN�|~�òɢ`=ۓE�&c5�	���d�Qy�m��<ٗM�<Ѳ(�d�0(�q��h0+�i�N���Ҷ ��Q��Z�O�N��EZWn��%T�ѕ�ԉ�6OJ��K<�S��f�M�*���PM=�5��.2[��'�Q�PM�|�"�D�$\*d��{R*R2n��b?O|Pk�j+��A��D{�]qqO��� n�P/i��|�����X�se��KuR���Ž/��u��遺N��h%B	�ay��#5L�'�� U(͢b��Py� Ԭ1#��4�;D��C�ċBnD=2�^%p�u�@�8��N0����>�����%T�P��
I�XM��9�!D�pA�6:��j�<n����2D���Ф*����@�W�`���N2D���\�l#�8��LD
8����`�.D���a@'� ��֬� ,F���+D�0�k[�vsf�	�J�%m�B)�V�3D�@)U�ݻ|���C-ێO��[P�2D��)֍{5�	�En�0�~�j"2D��9��Dtvp�V"�BpS4�.D�d@��[4-؜��Q�I3S� ��g�(D��CU+�<1H1�VN��3��] Dk&D�4�rlI 5(��5�1�µ��#D�4X��M�b��AcnFeLU� �!D����M	B�@t[��+�ܨxe*!D����I����bG@���H%, D������tuVL�P��g��H1r�>D�tcaˉCe,}Q6�KI��S.'D����&�`�еqVa^'Crv�H2b$D�LѢiݎ^���LZ�)]N��k#D���ԃ�Aw��	"AZ.'�)���"D�\C�1^�
hH�#ͨF;�9aB�;D�xCgDdxI"H��<\A�vj:D��(Q��U�����e�-|�t�Y��9D��Zj���e�4>���� E��!�"�D�� �L���ْ!��>k�!�ĚR���Qw����Č/���Ұ"O����Q��B�#bC,��H��"On�	��Ū��i����j��	��"O���27�ᦀO8 ����"O��j�h\�X�8��M �SR��p"O�@:s�
</�@��k�,_D�r"O�XU��7��;S�ן�6�1�"Oح����c���B�v�.\��"Ov}��fm���R�?�)s"Ox�QBHˢ.��tP�����"O*���H[������)xx�<�"O��Ұ�_�r&�4���˂\��`"Oހ�n�+�� ��J*?D$ ��"O����<Sa���_.9� �"O@@%�L�3dl�A�"R�>��C"O� IbF��Z �L �MbFH��"O>�y� ����XS�_xX�1j"O*<zs%��,r��W�<F���ӷ"O$q���$P��1# �7�� $"O��eֆgZ�(q/S�*���X�"O�94��K���" lŚUZ<=z�"OvY1;�5��`I���A��y�f�\�@��R��g=�����R��y��T�`\�E��,�9��Ê�y��Q9W�4�r.�$"�労��y2��8H˸�@*��ȽУgܯ�y2h��B� t[�'�+� �(���'�y�Ċ�|<�ш@�&��dcR���yb��g�J�b��N�{b�ŋ�y⡘�d��aZ�6&t�qo_�y�+ko�8�愀Q_���E�W��yeGNv��׏�Mq(	[5���y��.�he�ܿK�ո���y¤��nVpٹc+��B�� �U��y��� ���d�n��2�H�6�y
� Nđ¯ۈ7��z��ՠw�}S�"Oޅ�j��[mR�(�$	vh��"Op��e"��A�H��a�K=cb�JP"O|�k�"�)!���i��Гp�`���"O���)�s����P/"�)9�"Oİ��?$�Hsԋݤ$X���%"O�<
0��i�$�	�J�&~:����"OPl��ď�*5�P��L�"*8���"O�c��ћ�0]3èG�	�ڱڥ"O0�1㒴bdP��M��P	�"OJ�Hf�l�,��2~ࠣW"O���(��l�z�n�Ã\k���"Ov4!��
B�c`�;<f��"O�%��a"t9Hu/ґW��M��"Of@�� U$�D�FV{:�X%"O��K�a��y��8�֭AUq���f"O>�{���u����,فa�� �a"O ��5OΕ7�Y�	�&WN$!	�"O�{B�
5h������!0�D���"O�e����	G��a�"���*�"O�h�wm�"s��t`BHƦP��"O��*�˕0��|w��(~�BT"O�����}��(��4J$ Ȋ�"O ec���B=��K�-z�,*�"Oܥ�6���w���Q͜�Co�PA"O�%�B��۬� լ�37���02"O�<P��\\�������)6~�aC"O�p�*TTMBPʡ*�vlD#"O�9Bf�ƿ.�P#rI18vFL��"OL�s��R���E)���u@�"O�� ��)�P�� Q��$q*�"O8�#�L�`jL�HegHz2�S�"O� �D���<�P���(N]�$;�"OF|!J?bu�I!G5S�Lx�"O*D �*�:Og����O�K�b�C�"O�hc'��?d�Ȉ���D/J�&�s�"O �j�G	;.�E���=V��@�"O��+�I��XQ.�sR�/<�%�p"O.��VÌ�F���a�̷���ʷ"O��� R��t��e׊U�$PC�"O,��a�72�0��jN�}��"O�a1@�DZ\ak'�X�H⬝*�"O�S G�@�@H
�E�v�<��"O2p�u�i��)B���"O�m�\�2�i���fm�d"Od� �;ގMS`��
��t"O�8U��>&��P��{����"O��aQ���[����hA){�1�6*O�T�c.�$8U�����$u+����'SH� �X �������a��'H~(��I�Dfv "SÞ����'l�!�gƟn�ѐ��MZ�px	�'_���g�Z�'�<a �`Z'���	�'�qp����O�d�W��6}B�Ъ�'"��Uk�;q8��7ƞ�*ld���'��Z#�ň)��ңE3u�
5�'vbDy��4=�����!� �i
�'9콣��ƝB��X�b�މ+�U�	�'l.�r����E��3	 ���'~���(Q
=݆�`Ҩٳ(�ʜA�'�����5EB���ʿIxZ�9	�'FX� ��O��bլR6=e�d��'��Ԑ�L�����I�"L��ة
�'�\U�QB1fH=�$�Ɨ=�H}�
��� ��-[�pԈ�h�H=�Ԙp"O�[�ƙ�v�j��e�* .9P'"OMr�hՉ><`�;!+utAC��'QqONL;0N��qX^q��*Цlp�F"O~4;��Ȕ�C�*\P��@"O䱸v�ñ>��� в]H(�ɳ"O �"R�JM�t�@�$\+�i.�!��g��ˢ��'q�� a'�B�FL!�$E�t�\��h�C�r���΋�!�$�"'Fxhkʷ�`����=z�a}R�>�T�o�6L�-Zuਢ�.�[�<��ȗ�N�h�*�P.���oH|�<���ܖ�\P��N@  ��%��@�<	g�H:'��C��ي*�X(�'�@yx�$Fxr�Z�o����i�
��Q�Q���y���zw����ۻ18~�r������"�S�Oq�@���_?i&��``�4�xC�'J�dp K�66�^�X�	�.�	�'�p�8�jM�*u�v���uD�	���~rkMp�Ƀ�H
g�&��V�ī�y2L LPfyه!�_�<pXF�Y��yR�2R��1��Z�����iY&�y��H�c\¨:���J�vq���F�yB놽2i�� ��E <G��8$F�J�<q��$c�<0z��ב&S�I� ��o�<�uN���Rӂ��qy��P��E�<ق�ӓc�.��
��f���i�!�C�<i���v�H�h��X,ku�y��W�<i����`����86E9@�O�<���
.fe�t�&}���$��M�<)c#[�zc�q�.Z7w宵`Ј�Kx��DxB
_�W��+��^_�T��n%�y�	0HET����Xn�|�`���y"�R�r#P����1V�,Ey@�N��y򥀣`�iBS���RlT�!���y2�Q�R�Aq�m�`���Wl	��y�M	�x-xU;-��^Ԅ�� ��y"ʌ)Vn�y���W4�����yB@ʳV�����OR�fU�E�ߵ�yB	כ&�V�ؖ&�D,j��H�y�'Y��"ܹ�b'C}Z0q�n	�?q�'�^ r�˗I�xd���ط&�Z�S�'@6$yF䂜t/�aK�IU"<m1	�'s�e����X�0=(D�^@'����'����_�]0$4Г�>��=ˎ�$>�S�$�<p�܂C�7e
�$���I��yR@:��{E�5c�bmS`i��+vў"~Γ/,F�+���	�:3�@�tF��ȓ+r� � �*U�P � ��:�PY��6�37�� 8y�k�M|,��I^�I��%z�"��R�L�M��bb��x��󩀎?<~�P�m7����N��?%!�d�8-��E:��:$���Ƥap!�F*t��ĳ��O��9u�!o!�Q�D'.[�O�>6@iF'˽cP!�D��3�6��ԏ�_%6�yf��:\!�dȩ0�v� l��T�9Z�!�X�}"��g�ؓNvh�	�	@�!򄌇1hH䧗�ewQ�('*�!��\Np ��ܛ^��*��C�b(!��9r��h��z[N��u�Ӭwj!�D:[e`��T�&%{�\���9"�!򄘾[X��aw�Y�ft����l��!�߁+��и�˅�>iQ�&ɌV�!�� H1�q�^^�LT�hʑ-�)�"O��K��(g�N���G�'�T �B"O�����Ť he F��!"Н�S"O"�XL�z�t49�E't��"O�c�E�0l��3�MV�|�l�3"O6��
�v2��MЦG��|�"O.�a�ؒEd��� -@�Q����!"O�`H�&�$=΅qū嘜�"O2�KŇ�,j����*P���T�P"O��!"�
��33�J$O��Ѳ�"O�q ��.
Z��r�5�ڵ��"OPh�b�߰Z�! ѶY��)@�F?D�tƣ�0"�2�ʶ���*�y�E<D��8�	ک ��1�% �@A%D�����;l� ir�A�=��l�cm?D����$�r� ��M�:Qc�*2D�X!���7T�B��s�NCB	S!1D����cƷq���P��]���P�1D���ܻ�`E[5��i��YP��2D��"�!;��ڶ�X�	���r�>D��!���9�H�bu����0D�̹D���.�+�
��δce	;D��3�Ȟ�pgX�`�&Z�%+T1jt�+D��a`��N�01�,�YL@;!4D�x!G+
5DM�QJڏO�R=
��<D�ܚ�ˌTTmR�Y0�j���-D�d�dCͳښ� UǗ!f�z��&>D�X! ?!\��C�F�m۴�KC+9D�,�E �++
r��$#�� ���J7D����"K�n�e��W�"$���3D������`�r&�W9���k1D��9�$�##���IRA��/R�B�"%D��! ��<*3���7��<��ȃ "D�`�� 9W�uq����se#D��k k� M��źTA��4����6�"D�|9Q�N���(��J�~2�!)E�>D��Ì�u@���Ћ�3���L=D�x  ��p��h�D˖%n���R�;D����j#9aƝ� �T�Np��)�B;D������~t�ff:{UXU�7-=D� 
u�	�=�1[S*ڴ2��x�1K=D��Q��q�<�8�f֑O � �e�;D���J�yw�u� ZwOڈb�:D�ȱ��>��{�v�t�#��9D�t ���:VWBq�a%�]�\���5D��1k��T()��T# $j1Ѳ'5D�$�F'8nR�9�Q�&����=D�+���u����"fU�$��+8D�@�"Y�O�TD�#�J7 f܂%�4D���NiÆuȥ#ʞS���ä1D�X�У��V�2	�g�ܐ,�$�!qk.D�$��LYgDd����t���
TC.D�h�bJ�u�+&J�>���RF?D��1�
U��X��%3^P�8��<D�;�ÿ;(�m�/C�J��K��&D�H�ځ02:���ʞ�Z� !�7D��S��i^ġ��"�,�k�`7D�D�b���p�H���=~�a2b'*D�X�Dm֞"UHă'ܚ^te�`a5D��I��Y� 0�Lڵ/q^�r��%D���0-�
	�`W�L�f�j�q�5D�T����9R iS��Sh8�3O5D�l�f�]�옉!���!� !D���`˞��24'ƹP���uc4D�� �E!g芌5�m3��U!u].Mkb"O<�"���f��p)YT=p=��"Ox��.��aٶ(��C�n5�b"O�����90fR�a�g˪3:��"O|���S�������%��j�"O6E�%IE}���cD]�s2"OJŊg+í���	m����ƫ	'�yr%�W���ʂ*�)iژ\���
��y2L0Y�f�1���hC��׈�y�I�XWy��^�]����`N��y��ɬwT�E�Wâcaj�b�R��yR��/d�\3 BAEa� c���y��J�L�r	�)K����b�V��y���*g=�0�F�L�~����E��y��ʉlm8�9uMĚ}� ���΀�y�̊���ʠ��	�Z�S�6�ybiwr���	���������y2�\0/�n�����>&���צ�yR�Y�H���%"�4����V+�yR��f�9uG"��I��L��y��u`�}��H��e�y��W�'��h��/�.+fP9fb֍�yb�B�m��@+R�v(x"�)�y�,F#�X[���2��<Be���yr
̎r�J�8gS�$T�<`"�˅�yb��0qXt��F2"���y2�L!�dɻ�ԧ���s���y���h�Xu�"g�%A�Y*����ye�61&����(w��kU%C�y�K�"kL�� f��P86����y���9%& /$؝蠀�T�L�	�'B���&��$�\X`1�M?J���'���
�'ӵ$ڡ���=�\I�'�ԙ�D��n���c!��/��!�'��E�T>Gp��3@����ph�'x��-D��"�0�bР����'��1%�S� �u�îU�rD,|p�'�L��d�H�A��`�e���%�v�<Q��ֆ1,Xغ�o�:u}���#��M�<�r��9,W���&fL�< �,A���@�<�%^C�x�XL/_��l0&M~�<yvoR�1�p��`U�3)hI�R�y�<�(Ο]����T�ϮQj���`Cu�<1�ꄛbށ��A�h��Ɋ2�7D����a�>l��X4��?�b13r"7D�h
E@�-3������*8\�2�#0D����/�
}9��b!�O�,%0��8D��*SK�6j��SW͒)4v�r0�4D��&����ĨZ��V<k�<s��3D�(3�ES7V
���g�*b�lH��3D�`���0�F� =�B�ǀ{�
C�	 >���{���`q�8�`F�N�B��} nM+���� �|���� ��B�I0�� 8c�$;`���[-�tB�	�w� �8Dhօ,Y2m�TC�)O�tB�IˎIS�$K�Z�B}P�	E�o|�C�ɫFu����A[�@z}1�X�0��C�I��I��a06�Z�`s��@�HC�I� ;�M-w�|X锆%vTC�-<�^Ԫ�k��]-�Tb�
�"g�@C�	� �����)TnD���n4C�
A����]'�>��#��y#�B��3h��ȘCB�O����D�P98�C䉡��� �I�#x�U���!X�.C�)� �[=)kj)�G�3k��(��"OX��Rt8jl�`�E8,)�"O��T&NE�PE�կN|IJ8��"O��ՀB�H���`���"OPy��S�eG�$�l�#]R<�f"O\R�S��jz��BVF̵�a"O<�B�"��7`�P��d��E+�"Oʝ����+N�,��co��'�p!� "O@P;,ٓ[���VoI�F�8��q"O�A���Dh ��A�,ǜa��"O>����/ZN�P��$D�|Lâ"O¬��� #��p������"O^� �A�;�|ͳwl�4uf5`�"O�@aF� �l<���Ń`��Q�"O��F�֑a���/T�|���w"O*L��-^�������S�bԲ�"O^�Ebw9�-�W��*6��M�@"O5����b��U�A��}z1"OH���,��@3TE+���I�"Oa ��ĳa�t���F�w����"O~L��"��>\�9����-0B  "O͛��	�BW��"B����RaI6"O�t��BC�,7Z�QQn���[R"O��ný���1���4���ZA"O`�ٶJQ�^8
m��b�[D��Ё"O�C!�	���x���R/-�D4jv"O<[�%��J��V@X�.�V�Zr"O�5L?lX� k'AO��
�h0"OY�r�� �h��v��F��x�"O:X3X�¦���`�HLu!�DR�X	FM�)6���se_$lb!�$�fk�@r3ϸglj��d��L\!�=$(`���@!	1Z,(p��2jK!�@0��7LR�t��{�c�(U@!�Y�n���d@[���uHS�\)!��?l�Q�b�G�����NH�!�$ׅ�,%�w�.~���Ҡ*Ҵ@�!��ȼ"(�ٷ�]z��8a�̉t1!�9S}#�ˏ�0�@��&�!�d>e��A�A��,�����U�!��%Q��E3W�]�K������j-!�d6�v�aa���8�N�aC2!���pX�L&��
N�8(�"]�O)!��w"V�#(���``�(
!�Dݐr1,U���k�t	���"�!��W��	�&ő�>S���;�!�Dǲ8�"�E≯R�6x��ʗ$]�!�$N�1����b�=2�\��� �-�!���"�h[�ڦ:h�C�b֓4�!��yZȘ��K�SHμ:e�ј{!���;�D�U��S�8I ���-0v!�[)-�&��0��7K��E� H t�!�$�3e����[<��d:3��j�!��7#���!�%� �FCҋ#�!�$D�q/ĭ�d�(�ذ�b��-N!򤊼/�(a��Ԫ�Ul�{0!���(�(�h���l+$��AL�/8�!�DZ-*PPx��,Y�(E����lΣo!�Z�^AҲ�3
,�8ȶ��k!�2@�t|���)+����-%�!�1EЉ)���*�h��On!�$�*k�Q�S#{�$�:��ىia!�U&�}����f�%���ЋU!�DH86��X���Y;���ѕk��+N!�� ��#��q�:��C*T#X	�t"O�����߅A�d��a( �&�)�v"O��@��z�>�: �R�U���"OKǈп(�rHh'�=�pe�p"O��Z���Q�֬8!k2(��{E"OD�9qR\ A��ɛ�1#T�� "O���Ĩy��c����R�z�"O$��:XX�Tر ��zɈ�"O�����}�H�he@̴8��0��"OJe9s��)�,�zB��'>�lՓE"OHS�畭����mO%
��!�"O�-�Slܴr�"܊��I��� ��"O�ԁ��)eR�J!*v|2�"O� �tC�%E>��r��ɠ@�*t��"O�5eG�H���)'nQ:Eg��"Oa�A�^l�˂ `. a"Op�W�+r1�Egj]m���"Oڕ�@d՝M�(�"�o���"O��PENƱz��9[t)��$� ���"O֙	�KG�H���R� �0,��"ODx!�*��Lv �� L�M���� "OV��6��
�����@�4�k�"O����BȤS�V��0ś\�����"O��[��,1��t	��LPu"O�{���Z��+�A n��5"O���c&�=��iQ�`��?ȮMjs"Ot��3�?�0�I�3Z6�[�"O�p�A�z�Fm�H�LA6Ո�"O"��N.������D7���1"OZ Ԁ�H�.� I�4��4"ON`!�
2'?0�Qs��:N-(t"O�x�WJ�j\x���OU�?�D�%"OT��Fmâ@���r��M(=�\�D"O���2@�=0eK���e>��"OĜ`�N�vdXrc�k�0�K�"O�բ���."�YPI��66M��"OQ��k[	r������x.�0�*OR��Tc�=5ΰ��B�B��Hu��'��vD޼58�s/� |M��'�j�RL���&�2&�fzؓ�'���� +ϥ$	����@D<m�d�{�'s�m@g��%\>Pd�'O��Th�$��'X��E�h�a��툲>�Je �'s� �@l�[�Dxh!�K</��0��'x�[�p�И�S�$�
���'F�<��ګ�$�0�&��d�P�9�'� |J3��vU�����)��j�'�z 0��V����htT.l�8qi�']�%)��D"I9�)(�L�r�,#�')��ȶm�d�|�bcY.��-h�'�l��3�^-f^-0�o��P
|�z�'��	9 C��,��!�M�V��
�'Ҍ�0�LŶ^��h���>> =`�'j���BԼI�l�P��9�6�s�'*Zxb�hؑ?����	NV�M*�'��<c��ɝA�b1x�#ȄӚd��'l̠���$l\�Ц��%b�*�[�'��@�Q�q$x�+G�R�"��	�'v>���'�@\[v��v�� �'�j���I����кb��<��'9�h	�+;,H��A�'Z���'#�3��Ӗ?�P�k�Â
MP8Y�'톙���کX�聸s�IБ9�'�v�� �]�1p��9FK�@���� T�s����:����ƈ�
�8�t"OR�sD���7����$ߘhlr�(d"O� "����T�0YbuDBR�$+r"OzȊ�GK������57.��1"Od)x��G�+H�Q��
�0,�~E"�"O �����3f�ph�����-p"O�p[�
	f�]H1��o�z"O~50��J�f���zcM�lr^ͨ""O�}��o6x���T�A6�1d"O �{��D��yw@��0�"O��"�ţ@ � &����x�1b"O�ХI 60�h����Z����B"O(t[��ܶ|*�3%���nq��E"O��`�W�B���E��Q[�t3`"O��x��A�c�B"Ӓ]U�  R"O�mqEb��r�X��Dk 2Ra��k"Oƥڄ�V/`:ƥH�I�V��)�"O�9n�c%��#d.�'^
 ��"O�x�d�ơ��!���Y��	�"O�� �"�||�S�׻:��Q�"O�ᐕiU:ZE��.�
r�8�v"OV�����>��1�8^�a) "Oȁ�H²r9��I��ҟw,$)�T"O�	��� 0�D�҂X7˂ �"O4� ���05��BE�=��}KQ"O��"���YU�衂!K�l�(���"OxD	�_�#������8~R�{g"O
QaD�Ño����><�&�y�G��M^��P���ub!�梃�y���!�^i�2˓*r��M ���y��C(j�6DXvHI_n�|����y�N.e_�8V�DP�P��퇜�y��J�C��$�@(M)�-��,̲�yb�D�J���A�87\DX�I@��y�d�!V^�M*FB)3l�Pu�H.�y���O�QS6l[�*-�1	U��y��,/�F�� 
Z��J^��y�)�J�c���
X����E��y���;�đ{ġ��	�H`�ȑ8�y"%Ϩ_��a��X�1�6���y˟%�>,��Z�.`F��U�\-�yRD��'�p9��٫%��9%�Q�y"+��n��<��H�
ٔ�:#F�3�y2���g;>���
�)���yҭ���yB�ޱ<`�����J�����d߼�y2�ʁ��Hƭm�d�b��/�y��&4��IC�ÒP��+'Û�yK
S;���Ǣ��!x�',��y��@:VH�@ � �|ܾt#�*���y�"��H�t� &u.�R��-�yҩ�'>��!���]	R@s�����y��9wK�<���0H�z�v���y�(���"�õ�F��P����y�6/��q��Ռ�R0([A�'��:&iU�KD��`��آ#,�8�'���� I ��tj��' ���'�nT���ݶwlN�@ڼ9N���"O�m�w��e���	g�+] �M�"OR�)v]>Ernd��	��P�`A"O�(gi��q֐��b�7Ԧ\y�"Om��H�I����aͪWi�"OʐkSm r�C� ���pq"O�᜙a?�\���	S���"O��s�
JxP8��'�4��a"O� :qq��L|�	����d���"O���5�r�b����G�i����"O�-���ʄR Iz&�Z/QP^1��"O�� Tk^�C�X���W�TI��"O���P�K�8�8�a%��!ڴq"O���@@(7����W�<��!�"O~�س*WF�p�	6��d��L�E"O~A��$��?�����!l��X��"O�|j!g��0�yc��g(� h�"O��
d��ke&)��`�<B}��"O��S �#����G`E-I�t"O�l�ӇW��d�ʍ?I�0m��"O(q�&�)q�Ԥ��)D�X�b���"Oz�jӦZ�9>DP�'X� ��d��"O�Y�qdn�R�8��ApT��@"O�AqC Z��cRu����1"O��)�3!0�̲� ��r֮�Kb"O���gG4��D��òu�Ո�"O8\Q�%�>(o�8ӑ�Tj�Y "O�I
����v��(�y�׍�!���hTkЍ�!j�:M9P ���!�´5�X �Ձ"�^1�@	
vD!�?h��c���;B*%���Q�!�d��>�9��Jؚ+%:��%m��!���.�����{!�q3E��4�!����|�P�Tl,�"�HT.�!�D�1�U�DƏ
LΨ��gLR����l��}1e^�s��A��B��h��|t�w�4T��5�
�i(j��ȓ ��bQ�z;8�d�$Ae ��ȓp_Ʃ��EL���ՙ�m	���	��pʐ���ۂ^�Q��jX*�����e������25���u�����lt�s��M070���V�D��؆ȓ~Є���a��!�(T�#炇��ȓD�<B�Al�B!�W5P�MV*,D�����V�zS���`kW�}�XA�*D�h����-���l�/K̤q�vk'D�0V�>,�d��q�H�%�@�R�b%D� �@J'o��᱔��<����� D���cgc��d���J�lj�>D�P�� �2�X�+R�n pЁ=D�,#t&�$��3@�M�m��:D�"���*1ZX�zi� /,�Z�g<D����&Fʽ07��>�"��F�;D� �J���(9�`oM� � L���:D���d,�"G�d�	�>����$D����MJ#.�Hd��*f�*I�$�'D��H�`�5�z�XbN�0)K�pj&D������-�$��l�����D:D���g�\'�t�8t���<�t�;D��J�j�
,�r���z7��j 9D���i6T�Q#H�U~z�a�	-D�Ȳ`�DZ��YQED�t|z�C>D��!�G�^�	&��s͔<�'m8D�P���������C�zT�1 +D��j��]��]�b U	7L��q�<D��·g��p5�8���!�DXQF�:D�@��_�	������ $�8Ԁ�%D��+b,+	GU�錍<��e��e$D�����HX����ǶN̖It�%D��bv�/D��I�i;n��9hơ#D�����V,zx���Vǁ�/T�%��!D��`��N�t�	��F��V\H�� ++D�� �yKP@�7Tal�8�o��k����3"Of��7��/�@dS�LD2|�T�("O�Y#��@Z�E�#b(d*�"O���W�CJ��J#�E[���"O���VE_#F<) +�� �["O��K���4f`9 1�C���I�#"O*1��/B�
����j\�L��'�|�b���.�x�J��\4Ut81{�'����
�A��=�!�*K+�}r�'ҵaѪպM���!i�w�B%��'�Aܢ<����@�7aԴ��
�'U�Q��n:�ȇAU�G�x1
�'g�h	1�¾1
|:d��E�($�	�'CN�2�.M��ïA�Йq	�'p��3��Fh5�b�Ԃ?첈3	�'�.���
�37V
%RC�2<Bl���'Oވ�Ebr$����LM�1D1��'�H����N]���Ѓ	�-���q�'�:�A��1�5�/&�*$��']�x�!-�R_���ↂ�-�N��
�'����H�E�� �`�y�ĸ	�'dU�w�2J���腡���`��	�'��h���ˠ�!5i�$�\9	�'��$�A)V�:d>tH���3�\P�'`�h"�Ŗ!ho�G�D�e"O�p@��,?�ZL�#N��?�� �"Oހ�%�ATp�# 
FXp7"O��A`E��F��@��'��HU��"O�l�4��:-�~���&J�Z4��1"O��2si���UB�8�dR"Or`�#U�;{�p��G��"��r"OL�f�C�mŨq�䖼h�hS"O��PE͑8�	;�,͛7�R���"O������a�.A��6 ۖ�y�"OF��0�̏V�.�paa �"�5"O���"��.}�T[� ܛ~��C�"O�����')�$�h��m���yT"O�����'��v��-�~���"O�rYu�Sv�F���9i"O�LȳB�5�R��2�O ǚ�[�"OP}�C�;]>D�b��I-��ዣ"O"�b"��vj����W͂ B"O(�����&�����B-�`�"O��@�(�r��CC�F>�E"O���5�խ G\ʃ�G!V��yQF"O�p�a��=��hF�,t
b"O�\�G��tk8�X��F�m�<��"Oؽb�O��n�X$kF�ܣm�U#�"O��X�׵d���G%ʸ&���R"O:����#^�@jq���:c��ad"O�RPA�8O�>��C86���c"O,��������c�#ġy*��"O����#�7�|�q��W!G���!s"O�U;��Ǆ,���f!S�	�d\�@"O�J��,�n�*�`��dtk"Ovܙ��b�qʰO�oSP�aC"OLH�b��Ď�8�]��"O �2��=�6���&��]#P��"O�\ō���1[S((D����"O�tcR@\",��S!�χ?H%��"O�j�Rhr���A֏�A�"OXd����w�^���i��F@�""OZY��kJ�RPq���:T�'"ORt
 �F�x�x��'T�[?� q�"O� <���o��1Jf$�Մ��{Ԡ��"Or�J�Ϡ6��`G�A|xN�� "OZ��� l�m�e��?Sd�QC"O���(?UpH���83J�R�"O蔡!���<)b�JY�2�U�Q"O����P��)q��'��Ӡ"O@f��S]^�wBJ�$��"Oΐy�ŏ�yX��o��`g0�ɂ"O�Y���$=�]���Ö/G�ȈU"O6@ W�I ;���� ��l��"O�+s���v��f��
$\�0"O�3˂ .@~0@��TW�T�@"O|��`�ƾvR8�����j��M�"Ony��ѾaG��R%B�*)�y�"O��`+��Uz$�
��l��`"O���oƭ&�vEuj7���	�"OP�� ��n&�ʃ)`�,�y�)D�4U��aI�J#�YO�h�E&D��Y���r (<�H/b<��Y'�%D�re#�	&,�A �&v�P�vn1D�da��63<I f�џODQ��3D��)p�V�w`�q�5�\'7_�c�-2D�\�g�"_�$�����6l�`8�&D� K��ȑ�X � FG�pB��:� D�L���ùq��ق-F�5�h��Q�(D��J2�Y��D�� �čc\h�i%D��Yw$�&Fɂ������c$�P�B?D�`#���M��y1b]�<���-<D��;t�W�_v�̪�J�#�"�G�8D����	˞`r�t �X� !b8D��#�HC�*�a�K�%�Ш�6D� ���H�!`"�⃯�C&��i%�2D�t�\-Xut���!��Ev��i�+D��i��F�P&,Z%�ϝ:(l-���'D���!���A2�-U�j�#b$D��x�HF�?�q8�.�8bch-�H/D�h��KŢX�ꁀ�e��?$r��'D�ܰ���4"�����o���;#k D�����)�v`��\.
�!3�>D�X⤤�/,!����7z�[�$>D��B�e��Uy'�	05D�yd-'D������>!1,0���_<���bm#D�H`gI�X@���V? ��Ao"D�T�1��u䞵��
*k�F���$D���fԡr�"T �9$�6�2��!D��	p+U;I����I*.�)�o?D��b��L�́�enܾV ���1D�0��\1��L�� U�^�yφc�<Qd!��TY�{�Y�elX�Y7�b�<q��DØd+�
�>�2-9��HG�<і���[�q!��G} &�8�ϓJ�<��)3~eåE;kU>��.G�<����%s�N�r����o�F��c��B�<� -s�`C�"G�h8��I���D�<���}���A��(!v0�&�h�<y��E*8 �a�Ŋ%:�d�)�#~�<9�d�V1����CƤb?��р�I@�<�s��}k2Y��E�q+�YYw�{�<A�.�2��M�A��
X�p�GkRl�<����d0��0-ˈG]&��e�d�<Q�ǔ00A8��@-�=d,��T^�<ia�]�g��22��*g0�j%��u�<���,�R�kF(B�jdH���Jo�<A���	���0�E�#Z.�s$Rk�<� *ȳ0	�(-�y�@��e�R��"Ofa�ҡ�����+�]8���"OH���M������/�zK�"OFum�h��qF�V��N�Z "O����A�q��B�J��3�"O�s$��9a���a/�<��Sb"Oh�e#�2n ��2t
���"OE���5a��}����4+�.���"Ol���I\
b���8�j�./�>�#�"O|8��g�H�Xe���
�@"O�L#��-$����F�0��"O`4q��֒sF�mC��[�H�ԭ��"OJ����Ů ifʎdG�D	�"O�u��`���"��2y!��)W"Ol)(E���39Ia�%�!:�@�"ON�2�!��=�I�0�
!���"O$]�k�dF�g/(�.�:�"O�]��+�?����dA�5*��*�"O��C0Nٕc�$q�C�t(���3"O�[$[7Db4�:p�O#�h�"Od5c�g�n����A`V��"O��P�� DL��F,Ԛ����E"O@��tL	h1��bfA�'Ϊa�e"O��K�B3���B�12�"Op��f�՗��AE!F�H�\]�@"OS /ьbҒ�ytO�o���"O����	LKl@�2�˂p�@�V"O�h��nʼ�4�߱k��Bd"O$,QuÊ�:��(b�޿glN�s�"O�����5��1�ʀ4����"On�C�� �j��u�O�^>���6"O8r�6l������ɩ6���(�"OH�kܧ�$���E�w0L��"OK�E�0p�E��\�Ac"O�1`����5]�k����C�����"OŁ�S�Y
������O�$4@�"O�5��M�
-5 ������-�^Y�"O"p��ҳ|�de#�.R�2��� "O�����X7^����2$V�)J���"O���G�lT ��$``jc"Oj%9�NÏr�����+���"Ox�x��V7�����gB�:��9�6"O��z!�h\D��E�j��,k�"O� Z�g��D������̊u{(xh�"OL���~MZ��A\w5s�"O�a;���u>�J��՘]�3"O(%pc�X?8�
a�&  &� 4;�"Oj��fh@�s�Dqb�	�A���B�"O��R`� [�� 'ψ\�� Z�"O ����Vh���5��RA�Q�D"Oj�G�(r�B�*�dS�J�z���"O���AO�f��b7���a%^UYs"OfE��	�!Y` t�W-�<:9��Q"O����N��I�[87#���C"O� 0%%˵q�<�:���	?*�h"O�=����@C��1�EQ�!�T"OFx����:&�D��'˃
�쑂"O��A�j�9A�\P�հx�`���"OnqKe�ݐc��Р��9�f@�F"O�0)�ʑ+t>L�1��;�|Q1�"O^ [�Iȅ�D3B�αqt�`V"O� �E�<���$-�0mjH`(�"O�����ǥo��ȸS��&��a8�"O��B�DR����	S����5"O� e��MX�J�LTQ��T����"O Q�d- 2�FD�e�D��ش�"OqrQD�	Y$])2I0!�:�Ã"OL����]�L֚�ҥ�M� ���"O�\; _�=�T�Ԧ,��'"O��8
_��Ud�)N FB�"O!�F��_�s�b��E	@�5"Oz���&N>�
���	��"O������(�-S2��*�j��f"O�D�d�K+K���P�ܩ�2Q��"O���JF�%o^=$�q�5�T��y��	�2:��	u�.���#5#à�yb��%K=���ԋW�7% c4���y"Ǔ�~��4�0���/7���i���ybF�!X�d��T��S~�Pc2���ybM_�SN���f��?<&u��&���yO�z�hP��%�+h��E���
��yr��o��zPAT�U�4�pO��y2�C*��*�@֊=њ�w.���y�*T�CPX�T��4�Y�I^��y򡓔zy�Lq��ׇ,J�;'�ߖ�y�
�#>C6�r���*�����
�y�˂	[,� (�#���t#�Y=�ybm��/X5i�$X�5�,m���ߧ�yrIWbɡ�IZ舁(Q��y�&�r����.Nx��%��yB�n��I��n�YUa���y��B�2�F۝�V�ڥi�(�y2(V?lfd(	@D��~i���㜔�yr��q�,:�!�q���`5&�,�yBi0<*��Ga%!���s&��y���d F,��$L�&����)�y�DS<�j-�WmN(}��E02E�"�y�� +q���7eW�E��ы!i�)�yd��
T*��
E�Ha�̀�y�{Kh`i��[ Sx:Td�<�y���	r.e��o��I�7�S6j�!�$L8!�l:@/޸;|�U�F���B1!�$� >��*ԬcqFm[2�ǟ;!�$S�4����v�\ ## B�R�!��ɶ���3��+d:��d��$�!�ǄG6���M�a��0A���!�Dşc�4� K�=1~��sD���!�dΧCp��Q���qL@z�`
.J!���-S]6�ڗc��; �X��Z�G>!���{J��c@��	&$mr�F�J+!�C�~a\����3  �S��!�D�4\H|(�M݇s�B�@r3u !��R�s�xJ7	=,Q�Sb��n�!��D,�qx�	�V@|)ag'C� ~!�S��d��W�E_VT%[���>v!�dH���xS@�׀s84�[��_�!�D� <l��hʞ=�	p�!�B�!�@��"K޶|Y�����!�D�
K۲@c�F��C��{�'V�3�!��1j�������4y�aD���!�DN�J����L�%E��!b�"Z�s�!�^>�d����$�R��Q���!��E�/�(�(>r=�A���H�!��	�y������'5�(� jP9�!�dT�u�
hjq��� ��J�!�ɸDO2!㇫
F�9�O�B�!�@��Hs�	EGR�K7��X!򤀤 P��hA�]묜��KC!�� �� �ک(,�ܪM��x���#"Op=�m�H�Ų���V��Ѓ"O<).�"L9`d
ݚ(��UP�"O�U���<|�
)��#�@�dY��"O����	@r2����M�|�g"O\m&<wz,��kF�r"O|h�%Җy��� h�| T�"O�D�Յؙ}i�H`(�4A�H"O>@0C� ��d+2턶=�	:�"Oj�b�H t�p��^�*v�j�"OL@�aDO�:��|cf��n>��iR"Oܵ"��<L�^@0s�пIL�D�"O.ȡ��L��8��B;oA�횲"O>��*����Z���=Àa"Oرa�Dm2$Q2��f��lc�"O��H)~� ��sI�
�RP�"O̬)�NY�@>�-�ȓ�d܌qʢ"Op�;��QF��B���~��"O�1c����s@p�G�]�8�Ɛ	�"O���r_��Q�-�;
�mcS"Ol��$@�  N��9Q-Ӱ	V�mف"O�pw��k�vx;�N+6�d��"O:��pR�`Q�e,�N��P"O~�c�&D&}M��!��5i�� �"O����Bf�ƐX,I�wr�,"�"Oy�։�7r�+�%oU��r�@Ku�<@���9C�=�t�ۦ�l�g�<���; j>���l@�Sy��*�.�y�<��H�!� S:e3�H�"�J�<� �P�Z�b�z1̃+';��kG��D�<`/~���d�ɱ�x�)��L@�<a�� �9Q��(��"A�ȓ'����X�!Ȝh��K�-@��͆ȓ.��$��B�6�J�ZE��.%�<Ԅ�mœeB*(�!�r��T�.��`�ά�f,��t
� ��G�]��ȓ*q�|�&k�Zʾ8��k��7,Єȓt>�r`l�h�ꠂC�ڨ�d�������RGP�b�0��GLO,��܅ȓ)���� n�w��pr��%"d
D�ȓtR,㵩K*,x��b��1m�`��:�݋�f׾|�������eĂم�.j0�x�&�/	��`��<z�ڬ�ȓ��US��'�j� ��y��E��A��|�2�:{|���(�3~��Q�ȓ��r^,S�n�Jᅔ�,��H�ȓ6m8����=�J92W/�: ��U�,��aZ5�@|�%��$����ȓր������7�r��#Y�\*%�ȓ^��Xۖ��2�v4�gB!~�A��Cc*�質A�_�Y� ������ȓY�F�K2��~�hrDC��J�\��u���靼S�ųw��_ݶ�ȓp�|��$U��1��D����ȓw����[-+���
bĸ1��cx|���_B�V�&oL,G��ȓ70��G�Vl:𣧮^K(���ȓS�BmCѣ
W�Ybe	m�v���Ff�=�5HԳ[*�T:Ĭ��N16���uaR`QD"ϚE���[!rE���:=�"��6H�AvZ�
,D�ȓ L&����?TŤ	iF��2��4��+n���ș�-8�X���Q!�$�/�F|z'���5��s&e�.O!�� Ru4�W�-2�q���T�sPzH�"O�y���ZHl�	T,�4>F��"O�h�A������0S�9G���"O��櫓�"kT!�rʝ���P"O�1 �LVC��#�"
���`�"O(43b�[T�`��@M=T8@� �"OB���@�a�ҵe��v.(���"OH�H��éc�)[焞4PMd}�e"O�4��Ě:{�\�� �(�r$�b"Of�zs��J�t	0EJ	
r�6�"O>i;�\�@����Vh�E�&Y+d"O� d�U����CV��]��)B"O&���7�&�/9ή9�%���y��D0���R�ό6Soh<sD@��y���6�P(Z�aT c�򡪣�1�y�nE�h 7�V]*#BͱQ��C䉝 S�)�B�4���qh�(q�bB�I�'b>�Z�7���wDH%]�C�ɡ��A�p!�.t���S���<k�C��t wF�6�>=y�(D�K�XC�I�-�������I,M%X�C�	�5� ������M�������%��C�)d���te��vfr���
�NB�I>�2���Zk>8��HM+C�C�I%ls�(`J-8W�Y5��
  C�I�F0C�Q�v�*&^��/D�� 
մI���R�J�p�ZȺ 9D��!FQ�B�v�J6�
�O���5D� �E55�ہIM�_3>�u�5D��ؕmơ��`ݛx�aD#?D��h�D�(2�D�iG��K��Q��=D�lgq�!�q�ʄ)D�U�Ӆ�~�<áG"� z"oX�-h��QW�}�<���9B]���:u �AE	Wq�<!��<-��[�m�A�q�Ҭ�C�<QNX;.��VlS�O�t�5��@�<�TjA�$��rr&�	��@����}�<�u�E�;.<�S.�<ETD�#u�O{�<9�c�/'Y��`œ1~�beG�s�<���]9�z3��l\B쉵k�k�<)V�bqI;r���*�0{���r�<I�(�+J؜�qeN[a�����c�<YL�
�x�N"��J7�]a�<��#_�<k(1�,��)���h�A�<I`�K�W�
��&i�?T��,a��UU�<��g@4�����	>4W�����G�<�e(z�.��t#X�=_J$�D�<���~x��%߫�^����y�<)ဇ/X�"��2L+GBx�Cu�<D��>� �Ώ���S"EY�<���ϨN�^|��" �ќ�[��}�<��8p�L��pKG�<�t,�E(�x�<��&Y	PL�e�
yE �(6H��<q��ۛ 
�Q�a�A��d�QnF�<��c�?�b���)��L16 �"m�L�<� ���`���*ΰe�p)��a�<�!O�)3lڱ"� �_
xU�G��`�<�D��3 �&��$(c���U��w�<�!��8j��Q� *
:_z��P��x�<y�DOD4d���8FQ��귣�K�<��� �Y#4LȌ@wh�X�D�<�R���{��3EJ�[��5�ǈ�@�<��)g�UA�
W8[������T�<��Ŧ	����	�������i�<� j��5�	�c+��K�KN�n�z��G"O�� v��<�1B5��*l�l�h�"O��B�f�;J��(;VF�f����"O�L�P!G�y`trs�Π����"O��F* �//�|[�TSo���B"O��)���q���᝕�0�!"OLPqGHT6u��o�~�h��"O��iT��M¦��-Y�J���9P"O1�'��������8*�4( 2"O��㜙	�(��-��h0��"O�`�2��P��MѦJ���"O�Ɉ$��X����MR|m@�S3"O ���-7(�ȱ�l�`v pc"O�)Z',���3"���y+,���"OT�2c�X&1@�2��6"F�KV"O�{�JW� oց�C�G
9���"Or�������XH�&I=0�t�X�"Ov�1�ԋY	*�+�nU*�(��B"O��'�K�X�8)6�J��49""OT�7'=���7*�Fv�x0�"O���C�	-�@s�脪l2I�'"O&��aE]%��`	@�E�Ĝ��"O�%@áY�9��������Lq�B"O�# &��n[��ۢ�٧g�|}	�"O��	
�|�*Tjǅ�6 !��:"Ofd�pBιH͈�kU��9	���r"OhU�eK�)S�P�D"T�Ӂ"O>u��%,Zu���Ͳ'�8��"O&�d���)�����!�JC��b�"O�yb���G&��AϞ+,\�|"O�z#��02�H�S�,�i� �e"O"� �C�;�v`b�H��M/jY(�"O�4x��,� )4h�?P8�Ԛ$"O��Aqo�!]M��H^43F�"O^��c�y�D̫$l���D01"O�ի�X���h��.پ�1�"OH���ցw��2E��H��!�"O�}�-Ɛ�FQP.B�A�"OҀ�%�2=��B�Td�"Oj%����E�DI���H=D��m#"O�)�F"	P�`T+���E p"O��c��:)�AQ�,�\)D"O������r�A��5%�	�V"O��
��&��lA�&@U��"O����>#���X9xAR�"O�@��*�,����j�) *]�"Olx:��)
�kVd"�:LZ�"ON�@#�*�Є��̞N���Q"OT�6"�YP��С�I�u��I�c"O~��bI
%`|`p@���.$,� "O�|�t��,E�ZuA��ϣo���kb"Ob\����M�ZUu/�ⶐ�"O�IJ��C0o2"�@��� ����#"O@�ӑ/Vzt��c6��9UhB1�$"Ox�ӱ�!����vi��]_`"�"O8\{�e֚*�|0#P)�4mc`"OF�3�k\�[���%�Z�8��$"O0HÃA
4�!�ׇѻe>�[e"OE��jՋ	+f���& �hpq"O�]h�� `�0�z���@��@V"O�X�bf�DU�|��,ȁ�P"O��:�(��5,��9��s�`���"Oȥ9d
ư��	�M�B�"O��@��B]�3�"D�Vʲ�P�"O� �]P5獷!jj%��b�Z��4��"O\�cf�	4/�䌈��-L�$|"O�-A�l8�P��jS]�����"OBd�D$(Iµ3F��?n��uBs"O��Q�lL��J4b�.�'Rt�H��"O"���≐.,��XmL�h Mѵ"ONi�!�W���C $%��;�"O�ceI� $	����Y^}��"O��f	ͷ" �Y�Ϝ�	�P{�"O|�Fj)?
�A�H�-r�Z�A�"OR��3�Y)>�Z�)��*r�dmzw"O����ϕJ�<4I~�j6���yB'J>G�
<ʅ�Y?A���j�C��yB)փd��	Rs��l ��LC,�yᝍiv��@%��c^��%�׬�yb��H"pT�vJ��s_�*u�I5�y�j�! 6�|�$A\�g$�Z�����y�J�<���@X�I�Qz�ݽ�y��F�0��
%I7��p��I9�y�D���t�� �!_^�(p�^��yr��ffnE�Sj%Q���qb��y�)[N����"�4Wب:�ܭ�yb!ߴk�⌓եB�&a�0k�\��ygO$��̫Ů��!�H����yR�V #�ƕ�ʅ:!�nԐ0�ѻ�y�ԪlBls�-X�@)�P'�9�y��8#d68�c[
$�tC@nY�y�	�/!�|�*��˭�����)2�y�̤h�bI�0�ϐ#�4-b��Z��y2�E�bEX�d	ǋ?܄Ӄ���y"�m؈ݹ�A� ��1���U�y,]�m�<� �r��-��A��ybÒ"~���V�Za�2�+'J��y�e��\��e�O;�@pQ��R��y�&�>J�ٸ&+
iBx� ��y�]e* As��҃3-�ć�;�y�fݞI\-z �n�#2
��zRR��ȓմIQ�E�;�J���b�<X��"L��Fc�hH��,U�r:~���S=���-�3R����d'��h�ȓ;�VM����t�*y!��r���ȓ1Dȳ�ǎ7SVɣfe�� XЄȓCn��:0����K-p�>h�ȓ0t�H֠H>(���%Î�Q�0���P��]�Rf�?%�,��2,[#���3��k� ЄGS0�dg� �jɅ�+K�ېdC�e��\*�H=Xt�	��sOH�7!G�޲�)���5w�>�����X�@n ���յHђa��c����Fg������8�
���3����5l�%Qv<Z�b٘0�E�ȓ3:���t$��*Ĵ| �eR;`���ȓ[��j�B5{S8�d�ضJҀІ������ZB[�M��)�6W-���ȓ�psF�C��J�
&�U9A����ZU�PJCz��A� 3 �~B�ɕm� �a"6F�����c�C�I�dׁ�s�h��)�ex�C�ɠj�(� �	�rh�E� \���lLb�i!Lo�ܸ[�O�
nq��])��A� Q��m��AI1(�ȓVPmJw��4~u��a�Ԁfn�� ̴�eA˻VS���<,	U��7Zx
т %*���+J1�]��S�? �=�e��pa��Bn9Y��x	�"O�w��2�<xƯ�/$�F�Y�"Of=Ac�J�!���o�u��4ؗ"O�a�tL^2,"��� C���;C"OR�/W�y�Ȼ���(I�Dp1�"OBAء�^�<���; χ�F	����"O�\�6��J�Ƞ�쐠 �!`�"O��F�؄R�f�B�kN�Q��,S�"O�i���+=~+�*_!n� m�"O2����tg�=J�¦w���z�"O��RDĘ
�z�����k)^!� "O�|�پ��v�?����"O|93cMR8�x���ՓA�
h��"O��S (V;*ط�θR�Z9��"O�4 Q�V1rƨ�5�����@"O��� �I'g;�)aD\�{�4�´"ORm#B L�7��m�"�N�x(`�"O|�I��+|��hX�G�Whp(�"OP4���Z�XZx$	U'I�{{R�ZE"O���2+�"zY�,�@�Thb.Q�5"O�ȱ��& �j�e�G3n��P�"O� I�iD�+F@	�#/�'��S"O
�QdL�B��1G�\�P�"Ox��?�lH����'G�V�@C"O���'0����َY���.��+ҧ2�"���H��*���1.:���ȓ9ߴ���,��P@A�Z�ʔ�ȓ/��b�>��A�Vb��5�ɇ�[d6�i�D։Mʅ
a��o����ȓKdhƽ/��}��mJbʂц�t�Zm��[���K�aOT(���u��"Z<7@1[��dT��ȓRM���L� U�U��Y�@��ȓ �IrVmI!L�Bu�BcB�<Uh�ȓ��ᙤ�5N���r�GN����ȓ(�r ���ϑ�PкR�.R����k<n��&@Ɖ5x�����6v���ȓT�.}{��'$	�@v���y!�O���'t&ʕ;~q.��V�^�`!�D˾<#�D��ƚ	X��p�B�~INB�xVQB�Kv f���L�5i�nO��=�~2#�]�h������&Jl�v�S�<���'p��a0�D	��be���V�<a�E�,�������C�\u떉Nz�'N?��jw���%�RҸ�᧣;D����
=�!��A�'m~M0�$9D����
��E�@�N�|<�ɒ"o4D��b��Y�nIJ8a�ʋ�x;ru$h-D���p۵=Aԩ(VbJ)�L����'D������dYfA�"
6킹1QC*�	F���'����o�M�\�֧�&^ �ȓ ����	�4fY2��JΆr~ ��C��+dm��ꄙ��~��DzR�~�`��- 4�5ƒ�[��#��o�<�a��A�Ā+�gU&"Zs��k�<��H�=�4���S�1͎���L�f�<1���S��,zW�B5Up}�
_�IY?��{������+.�*��L$y`���ybZ�Bi�!���z��W��y��:�B���B�~]�!�G�Q�yB`�;��Uj��Ćx��IJ�	��yR��!b� ��WD
�C�0��%�?�?��',|�:`"r�^UJc�P<���'�0aY"*�y�vZ)[9Nڲ���� �p�@{t�D�!a/~�����"O�]�d)B<)����b%@<=�Z"O��Z�'�X6%�q��=ZjԐA�IC�'�� �1��4���`�g��o��A�`�L���5+t�QILT'I�]�.ǖ��c���I�:1���c,T�>`�q�,��J����)扦/7N�Ǆ�_�񲳃� VV�ꓐp?��%#�Jt��¦p� �#�b\�'??UCefùw�x�BF�Q�3��Qp�I5�x�!�63Ҡ��D&�*��\�揄�yB'���i@Y+|	I@��tB��	2�މc��S%r~�!6 A )0B�I�!(,�3A 
vX��]�m��C�I�?�T�4���^�|�Zb�kʬC�ɚa~E�Q�� ��٪«O�{�FB�	�a����vFY7$x�Q��C)8�>B䉂k��	Zq�AH4u!!��&�>B�	�#� 髠@W�B�����V):B�I�mw�$��(]� �4��9{P:���2�ɮ����"�KU��� dh���fC�ɚD�zdY�H.C��1Z���
ZC�I�>.�"AM�5z�ƅjြV(�C���<Mk��E�ԥ�©�;4.\C�I�^I��%K
�zL+u��	:jB�		5F�1��N�;n�0X��:B�	A�+p)Z�{R콘'+��B�ɪ{+D���-V1Q���(���<PB�	�a`��4 B�j�u�#']+��B��[�ك �ğ9�����Ϡ&mZB�I:(F�H�&��<a}��2�N��6�@B�	�J:� fΗ^{$m�ӄͿ+�NC�#I���pT���LR"����U�hC�	�E&�(�T�ݒJ�����W�>C�I'j��@�ï�r�)b�%RO�C��6?�6��ԂH@<ÁF*;��C�3�*(j������J������B�	�RM�S
�Kn���ө!pSdB��JT�'��Vh�I( `Q(HyzC�I�0&��)
.l�a�g� `�RC�	
9�U���Y��p���� H0C�	5_ݨ��āG�(Q8��H�+`C�I�?�@ I����ɩ�F�fW�C䉟4[����ɓ[̐��È|�C䉢Z��D2�(<@�H�G��#n�B��1�Q�R��6U��PC�@,X�C�	�F|сGX6|����Ǉ�&d��ȓ�Dxe���jL�x�D�?�z9�ȓMO����{�8`%fε*|$I�� D�j�0���c���&a��%�ȓ�&!���'���h��G">Dj���sƾ���N�(_��

>,���h�mʦ ��%2�U�\"�`�ȓ�>�"�MZp�6�\�F���A<)����l|�8A��	]�>Y�ȓ}��͛�b�2c��8S'�!Gډ�ȓl�&�R���z �A(M��7p: �ȓil\������,���BW̗�L-:5�ȓa��yq�_"9��i�YO�&0�ȓM"xڣ�D	 {��p��Cx&��ȓ7��TC��-.�����H�}q$���j(�{Tc��|�\rS�ԏ�0��ȓ�r�Ô'	|�������\��ȓE�x��P*Q�
�,�p#e�-=J��ȓ'.~�����=��=PA�?;:���S�? FĒ��2���@��'�R4�c"Ov���nI�oJ(�d.	#7l)B"O�����$p�=�'��m��"O��B��Zu��a��-q.��"O������R�3 F�5��5
a"Otͨ0$G;|��ԸFeΏL �C"Op�X3�-X��U���5R�F�*�"O���*ؒ�!Eb)+��4"OP!HqKҤ1&�JP"�,=#꼋$"O���4d��#m���߃f�f0"O�h �KˣŮ��E���F�*]�2"O����,3`�L�g[���h�"O��`DI�d�n-�G�?|�ȭb`"O:L{��,6���ɑ�<	|�mre"O�2���� pD���Z-Qm�x��"O����||DA�CJc�� B"Ov5�Q�Ӆ���$�!���'"OPA2"+
�0�B�"��U�1��Q��"O�ёc n��(�k̸$�8�[�"O�LxW̞;y#z�+3��;��1H0"O�Z�i�'7Y��B�C%}'XȻ"OzUW���0ݞ%�EJ�]2A{�"OP�7,��(p*�d�%H�0Q@"ONE��M���ۢ�y₰��"O���T�J�f~���0t��9�"O@li���6�T@��X6>p��R�"O�!J`�/0�1�t�q]x�#"Or�fJ�G�T˒��+SΝx�"O�
��MR�*���IP���v"O�eX�G�c𭫇j�c4>�S�'�6yK�C�7_+�"�Z��ViH�'X��ʞ
�Hy�k�<X�����'�	bV�Ӹ 
�����' �8�'3ҙ:�-	�������}���'���Qb��J��x��_�p���'+$x��[�}�tl�1�܇�
�`
�'63Q�]0M����N���D��'��գ�.�`�9У�����'��\��d"uÕ?��u��'�����N-;���${Ì���'2,p��@�44�N
����'����X���`F	܌�� ��'cʩ�㢀!@ny�r
[x�$���']X@R�<�����E't"����'Q=���$թք�H�模���`�<�0�Y�y� @I�l@ +$��0��E�<��ጣG.��K�OA��b�HN�9����<-�Iv���<�AE`	J�����
^HAь��<)$A_j�� �T� �K�]O�<�G0X`,*7	CF����$D��k�덉o��P���&2�+��(D����@���=aí���:Y1W�$D��)�1�^0 ��j�\=��N/D� :�m��/�,8�žOZQ��-D�`v��%R�B���.�}I�+D���cF6l��dc����f�T��#�&D�����:}\
傣��b�<:A3D�$0ɞ}�.y�6��>C�m
��4D� T�28�fЈ&c+�Y�F0D��hVAC�H�ݫ��
3|���i$D�����\�-;`�G5���6�0D��Pf�P0v�@X�E���D"D�����X�(P�Y�y�n���d%D��1�\�-�clZ�B��$!D�� ,u�0!��,0���3)�& ��"OЭ��M��T����i��^7:��"O�m�!)�b���� %�)9T"O�A�Q�S�r��!����"OV��	�\Ԝa�g/�h|��#0"O���w�E��zh�䖲c�h�#"OF`QRS.�QsBđf�ب��"O�͘��%:\ [�B�=2�̸3�"O����Tx�f����xI��"O�a��D�@�80F-6i�T!�"Othy�A�l2���#{xE�"O�h�
���c7o��q["O(�����c7Թk��Jy�M�3"O�t1�����,�欇I�| ��"OL��0�.���C���J�"O��Sa �)8�diFo� �d��"O\��Q,�,5%N�Y��U(3�M�c"O��9�B���� (4͜;�ʅ�a"OrI2+˼z��ԌB�%�&|�"O��� cؗNJD�bW���, ��"O2%���أ_��8���2�pؙ�"O���(O�/(*�Y��K�"�vH��"O	�'�P%{:|��Y 2��"O�X��`Õ's�e����G.�P�"O�� R,��5�h�7m��x�"O� {@�@7C��	J�Z	V����"OV5�l%lP��V�	"A:��"O�(��@�*�)[�+
�:R�9XV"O�tK��X�5Ț��7 ȓZ�=��"Ov@���ܶ`� tɣ���Y��(D"O�@��" �F��d�G�)<h��
�"O`�a��@=b2�����/���9"O6E07(؃�|�Ao��k���hE"O�ň0i��6ز!�MH�v����"Opi*���rJ�S�+��!��QR'"O����	+�@C$)3>}BHb"O6�:b`B1$��ԙ��ǬRi��"O�$*Q�
�v�|�P`��m�("O�mHЌ�r �0�d�D���ȓ%��}*�~�N0r୞��ڄ��I�~�L4z�x2)O�{B��*���vqF��^�y�D�3lhcăvІ�Th�����!5�PvBa�$�Gy�M0��i���#���y��0Xsڙ0c��#p���#�� �^�ݴg�S#0p��3@#�`��Gz�����c+��:��9R�M���<�CkH;��	)r��C���A�h�.DH࢓+�0Y~a��==�l�j�d �;��M��ɬ�,!˃W� $�$!��+a��' J�Qr� S�P���\%f}��:c`D�'�6�
X:�N݇i��"(N�x��4�!�W�<�b	�JE���P� �b�D�b)K�r,���d
�0b�&��,��!�"Ix�DL	Q&q�w�>��+ �\��z���3z\��'�8��1�֭j�"`� ǖ�e��a�r�fp٢�NB�ud�x&�޷(��H;fV,i�,xڈ���p������*O�m0�eѾn�џ(h���p8��6��F��Q2�%��]t4��.]�6)��gM��)`%��H��=�u���=�tfq��p@A�Y����ӆ�Ty�a e��:P�ϙ"Z.�qQ�/-F ́���A%�����8-j,Hkq �C�:$j�"O�X۔b^~��	��Aߖ�������ٵτ>b�`�Po�R��}�f�'��I�|^�"�B��KRHM�-�����VbJ�IG�	n؟<����ِe�&M���jE�%j���ġ�ͺ�ti�,�P���!��"!(A0�×H� e�?I�2p�X"�קO~8�F\�'Nrl��KE�4�$E���7�8W$S7|�I$(��u��ȋ���Y��X�c�A�R�s�K�|����?�Ddz�D�*�f�1/�>Y���$�B]�գ�z�Q�V(��q($b	�];h��'����Ex������hC!r$@�R�"O��BQ�ب#v����3u��
,Κ�"`��	v�	3�A�:bT��Zq̸?A�-Y;
��1��w�HIX�#�N�A��I�P��S؟xc"/��� bmx���2l�r�D_�w-p�4"V�qP�	�Af�"H��BW"I)pE g��f��ð�S�z��I�\�b��6�Ew��ꦃ�eC,�@vb՚L��uh$gV!F�\�ÉF�.0��@Q�Q�v5"d/4>�`x���'���*]Red@�V����O@�
c� 4"��z��N��\PՎ��1<<8�b�C�N�Sc>�$�B��
,�)�p#�"U"O.@AV"�5�(=K )q}�!F(Cb.V�b�3�Ґ�f�(HI.��c�\�bK�%λ�h|چ��13��;A��3p�q��	�O͸�-�/R)����
��f2�@r�J�M��Bu���p�BV@C�%Ӥ��tM�,U&�"=�pK�d�5��eA,A�-��w�'Y�4�p��*x1��{j�u���I�M���2��\1t1ԏ�0�����
.R����$�L�ģg-B2���I���N7�I�j0�)�掰�\�J�'qC�ջ�CVc����(�JO����w��P nժ�"O�%��g��L?��SR.R�
�\*�I��Zs�����
>%�$�HѠ���OKqO��C���_���ZfN�
��@���'���ka/��-Ix=�b�)�Ƅ����:�tu�2�V�-���.`F���82aڠ�0@��CјHxTFƙ �џ�y�JL)e#��b�S&����Q�F<z](ə���_4$�%"OT\Y���B�d�C	P�r��Ԝ�x��'ȓ#�����iً)\�G�DȚ�?Wf��a�
�%]R���>�y(w�f�9�aU�&��s��
�x$X���B"jްv+�th���yҊ�3
�В�ٻH�ho��Px�ə	.��u#��֐���L�0�Da��`Ҩ_3���A-z�ԙƮ�߼ �X<(Z�Z�(9<O����)^�R�O����!�1�!�b�ӛ�F��"O�9p�G�yj���ԩ�D�x�@B�$�A�|$)
�'#�X�₃�)�
�2�"|v*��c� 3�7x̑z /�1��9�ȓ{	�IX�C�1@*��vhğK2����|���B�SL�E��IO�q��p��e\�]Q��ƺ}�f��� ��$v��ȓ	ѰyY�L��b�X�"��L�����c�x(�$O4N�2� �E�1����
���{D�7,dUC��@�7��݄�n*��C��N�D��c�5I�����38�Л�K�.Dn�!%�	>!5��X��R�\�L��ȱ#%�D20��ȓr��h
T^5/�偕 0}t��ȓ��ͫ�]7-���	�͕(=pp���$���:6qCƟ~}.���8b���G�9�@	9pf��N2r\��A��JZ��8|�`g;.�ȇ�g��"��ϫtdP#Q͝�%�ja��e���cɡ82���2 �-{����X*�x�̯i�n��7��0[ ��?$��A�A�<�Z䟲_�La�ȓ%}<���C�	C�ʌ��/-��)��N��⃈Ј")�5���[*��e��O����r��WF�X)T��e�֭�ȓT/4q�S�����e
͝Oݲ��ȓ/�Z��/�B�a !��nst݇����H�&�r A���z��9�ȓ$�=���Q'I�P9R��='�bلȓY�l2bJ(r�LU�(����)�� t޴ˇ���#ʔ���L�쥆�,, x;��A�e5�pK#�=�La�ȓ�fd��_L�^���B����ȓs�"%��PGޠ�wB�.ͅȓUb�K���DO�tr���
(Җ��ȓz��ե��8N(2d��d��Շ�="��JK~��YdA·SS�)��WƦ����t���(��� -�ȓni@cDE���Etޅ�ȓ�(��E)�!f���Y ��7T_X��ȓP�LB���@��b��Y��Xq��S�? ���$#�pi@Oߵ��G"O< 1��� S�	JR.ؓF����"O� ���"٣�͋�q�h|"�"Ob�i�i�`��͒��.F�ze1�"O��;Qj��I��!���R�n�E"ObQ�1lY�Ye����9V a�"O�t�!�9/�漣S-\��\�Q"O��c�*�7n"�J�G��ԉ�F"O�(:�֣���H����5��H�"O` Y�d�P�l��m�1�X�x"O��Hs��(Q.��eke��"�� N�<)]�P�&H8��q��J���ȓK?Z�"ȂiklM�W�(B��ȓ*x�`�ƛ5r$�k�-͒ ߴe�ȓ1��P�$��X�AS�ᏓN�\�ȓ�j!6Ӟ j��Y1����l��Gk�,)��5��2w��ȓCM(\Xpf�/Х�B&G/njԆ�ya6䱡�B�}D�d�()𮠆ȓ:��Z�Ꞣ�0���o�3J��a�ȓl��p �Q/�3H���P�ȓyv|�ء!����@2�؅{v�4��a>V��!U�a~@j�)�=.���|���3g��H��	�G�.Ʌȓl��XD�4g��R�ȃ6 �X�ȓ	5�)x�ʒ{U�}Zu捸ub�}��4Q����	(޾UkCd�����U��!y�LP8l�"O�.0|����.ld0t�T.�����X*e���Bْ���&�6c^����(k�ԅ�!�H��սFB�a�B�&{Q$��ȓD�4�a 
� �v�R�D�C�IV��T�D�]yؐh�֬H0EcC�	�xe�o��y��Ƚpt0B�	�.��a���U4o�4h8�Bƚ�B�I� J� ��_�e��!1؎C�I"h�t�ȳᒄ/���⭍r�C�PC\tzFUr�A��,E/�C�	�XxD���`$|��8���7R�C�	 2�Ȧf�U[��a�OP�^C�I-�.=����G��u��L&�B��Yta�'+*(����$$K7��B�	G��92JL�z��صDK�P��B��)7���c�!�鱤
�s5�B�ɼY�pɛ �,>r����� q9�B�@�Sg��8^�.���*AxB�MK@�3��Mee�e#�
	�6	
B�!z�ͳ�n��6�|��/�+�C�I-Dۊ՘Bw<r(KG��&(�C�	�V�ۓ��F0)���k>B䉢T�"e��NG�u���-J�u.B�Io�L8h}|�8�	H'o��C�ɫϒ�s�m�0c�H�Q��I	L1�C�	"z�F�k҃,4\ଡ�E5�C�	�!O�(U��@�!��
��Aa(B�	�P"hY�ב>h���T��C�	�uΎ�b�� T=s��5+��C�I*��Ur�˝OO�CuJ���C䉻��2�˴��u�Q,�_�C�I3{���q�۵	�	�(�M�C䉰)�&�"v�N0���ivvC�	>GB�� ���*���&��,C��28��3��k��i�6�1�C�I.c�xj�MLf�*\�V�U�6�B�)� Fi��,�7��8S��!E�6��"ON���o\6־� vO֊Q��\��"OP���_�P�Ƚ����C�u0A"O@��'[ w��A����j�c"OZY@֧\�/l �1� �g�!�"O0��gbې?:J�H�J�"��� "O��)��3Fl9 BB;m ��"O@8z��@\�����Ț�d	S"O-㍳m�lD���2����"O0�a�l
�:z8�����#J
��""O���3��X�@�'�E�VP�p"O�
Q������-ˈU	R"O���c��q�-	p%�kf�Jb"Oڽ��g�3荑$܉p�s"O@�#E]m���]�?DF�b�"O譛�Cz��ё! �z=��3�"O��
#��>b��/\9mN���"O�	�邰q5�8xP���u"8��"O�u[!
�K4�mp� {:�<"�"O��ciN����!-d/�9�B"Ox����P�Ro`�B���� ;Xh*�"OD�〬Ph@�3��]�u.&݉�"Oh0��E�33w��h�1X,X@;�"O�\Q�̋q�Qr&�.�8J�"O4�@`	�6\�ل�;+隙:r"O ix��PK��%��R���F"O���M�/��Q`�����1@"OA�$�J ����T�a���`"O Y��(H n:t�� ������"O�@R���M���)T)ML �"O���>>�f�#��]V*fi�S"O޸Q��M+yJ\q���<N
�2�"OƉ��h�H{
����"wr���"Oܥ�&�� ^q9�i�G��4"O4-�6JI e:%�1�� "O��#�D�5Q:���)�#&&^}"f"Oн�K@}UjE%��pl�"O��b	�\���J
�R�"OTaC���y����iF7f���C"O,��gFS�%�d,����2�`��"O�q@�*��C�H�r�T�"Op�R�JP��GD�M�F"O\x[b#]7!�5��P�H�D�:�"O0��"+�!���@��ˢ,�li��"OX�0�f �0Jt��KӓlJ��R"OH�0��;�8a)��PU��"Oҁ���߭LX̜Bh�]�<PQ�"O�lS%b`�j����]�@��t"O�#e&����	"$Ғn�ƴA�"Op���NKư��
c�:@�"O]@���b%�Ĺ�#F~B�5a"O!`���PX܀��֡T�(U�"OX��D�	�J�zUj �[F"O2)ٖH)8�p��$�KBj��g"O�����%>���$��TX���t"O<ѳ�@��~�Xg�Ѕ%��$��"O\|�d��=�8���<��$j#"O��*�A��a�)+�$�A�+P�y��PE��� ��"���)s�C��y� 
xi<A����S̶D�%A#�yMM�'��5��8�� P�H\"�y�ε�d���4��#��y��^�CVi�L�q8`v���yB�^��8dK�&h���ڟ�y
� ���%ͷr+agM^�E|���c"O���4gU,YD.DQE��3b��"�"O�ݹ��z�i*
�>A8@�"Or���7��d���C�1OflR�"O~m���̹'->l�i�"O�����ϕLK�hxŁ�|/rh��"OΈZf�[�=�zDY�j�4C��"O��ΐv)P�P��6M��<
q"OR��� �X�˅+��E	"O����lҋm��� C���n�<�R�"O�a����+���4L�[��ۤ"O�=��-�,�x0"'�Z )�L��"O6dYSdGz�r쁣�L�"��1"O���ƌ5������y�JP*�"O�1�"V�lQ�pI_���x"Op��3]0}θ��7	�@aЈQD"O�#�N��8��M�/׭=c�e�"O��"���/� �Z�cO%^X�"O`!�2g
P��1fAY
w"@��Q"Of���k������X$:P�$"O`EP�Yz&@B�	m#�la�"O�l�F˓�HH0ErUA	�#� b"OHUy����*2��hq��>%��[�"OD-����
3�X*��E��i�"Oha�@�׋<�.���.Pd8��"O8a�5�!RN,:��G�F�-�W"O:8�mݧf0����aY��8�"OTd���Ou�" �M�=��"Oʤ�� ʐ;��� �C*"��Aۂ"O���T@ �B�O4����6"O0�
�L3j����3,�:5P���@"ON)0�Gl*@��i57K�8�"OR��6f�.�h���=R|�1!"ODB�f�	L ���șE� �e"O�}�3(X#}2�pM�V�:QY�"Ou��/��<]Xe�06�9�"O !ZG�
�B�>m)�ɓl���jg"O6M�u��1_�X+��"(�.%X�"O��	��+�1a�7�8zV"Ol���Ɯ	<Z�H��J�X�20"OH�&NL�'�:�z�l�.D�"O����K�N�Pq�!�D"O>@1g�_bD����R�*���R"O������V||{f�ܯ�.�[�"OZ��U��~�n �#OV)�* +�"O<���	M��Xⶏ��>Dj"O  ��*�� ����	V�l�+	�'/�����V˂4x�痄#� y��' �����l�a
�+�Y�	�'�:�Ş�E�Z��f��O��Q	�'#؀H�l�R���fO�p��M��'o�=p�=�����5h�a�
�'M>P���#N�\8c'Ui�R�
�'Sxa��DZ����B��k����	�'�4 	TL��4� ��VY�H��	�'ݎ�a��b(R�#��U�258�'Q�{�D�<�V�s#�M�'6� ��'2��G��� [�p�B�ܜ|�q��'��L�B��8t-^��%"cF �
�'��L��J*~kR�`�,, �1�'����w̓4"ߦ'��2�X��'��Q�g���i��'��<��<s
�'�P�	��x��̱u�4�P
�'ʮ���-�6môTH��۽7����	��� ��W˒x�v ��é����"O��SrG\����� G� ���"O���UeL�p� ��EN_�@��"O^��#��.I4��'+L�O�nU�"O6%��E[��X��
_�=���;"O��aP�ݵ4/��;&h"w�L��"Ol����ר8���ϭt�P]��"O��K�S=(Hej��S*]�
�IF"Ol�g �*�0�WI�b0T@��"OHm�G/|nl�;���MY���"O��R���<�|e���"V" \)�"On@YQ�m���L�=#pl�"OP3m�>i<�sw�I�]��5�q"O���7!^
�q�J��oF 5�b"Ony8��U3tXj�Y�+�A��|[1"O��I՘nq�]*&�΃ZR��"O81ee���m�v��
�Fɻ`"O���!�/p*(x�-X1bƜ�(�"O�0;T� T,�z�fT"UX���"O�	��ո4&<(c��	�읻�"O*Y�g�h
q�9���P�<Q��"@60��mY�6����ARZ�<��n�dh�������*k.��QT�<��b�26�"����#Ƅ�G�U�<7�*Ȑ5��,�D؂���P�<Q�@�a9�4q1/�N󄵢t!�P�<�r�H�st�TӀL=A�zћ.�v�<��L�~*�岆�Ҹt���I�O�<1P/�y\t(2q(��*<�{5�F�<��.�3xQ�$�K�r\n�#��A�<Ic� � ��2�#Ǯղũ����<)��
fpT�s� <&z�qK�"Mt�<ڲX{���e�̾d�,tC7Ev�<���!)�~H:v勡G�d8��y�<�B!�5��M×E���Y�i�y�<Q�.��s�����̀Z��	Ū�R�<i�߹'��P�ɇ�(�n��V�<��χ.I��McJ���%H@z�<�j��M:�-��.%.l���w�<��9T�(��'AT�@��c�
^D�<�El�,e����rBΰ�J�BUG�<ѥ�ڌZ팭Aa
�$h�BFZ�<مaшZΘ�����2���N[�<�pG��)3؄��	�{,2P{�ARo�<i�V&#�,ak�B�9������i�<�1hZ�֐�Sɐ
�R�B�a�<A�
� ;�j<�F�؀&V:58��K�<�jX.�l�I:B�pʄ.�j�<�@�0"v��r���$�:M3�ώC�<)F�p�Z�Aq/N�7A���R��z�<ɒ?��K��ކ�E$�t�<a5Ň�,@��x�b���<`㉉w�<�f�S��0P�C��L��qRțK�<��L��l�H� W9r7������\�<a���|����h:M�b��'��A̓J�|���,^A�08��O�-N�8��'	��hK�+�Q���0IA��*� ᡒ|R�څ*a��S�e2F��ԅ�y� IS��F���y�"M[���0|r�ٜ����gJN8?�z4���Juy�Kߩ9������|��	�pU�D�f
ҹ)����U7B�m�"����'1\qxC!��������TlU>���"l��$����_M�T���'����6�'�x�S<Fi��}�"��j�����H�h ̀�k��~*�=�v/H�1���I���M��;Q 
ً3���m	�|X��ʄ.�����=8��d�UڮH�����������I��<<DXc��9N�`�a��:�f]���O�˓u+��}ʞO<RӅ ͘D2�q�F������{��@K���g�? �-�T��oT>�0��8m"�[��>�q�9�S��^��)0�Ӈ<qT{&��>���	�<�<E�TIQ�	ꜽ�R`� d[�4Z�W�[��%�\���O�8����?a*�I	nS�m�f��&c�`S��v�>-��?-��Hz�D�l���&>���D�	R<� 8���?E�`�����?)�c�O���CDM��TP���F�,����(K�:bb����3$���$B	qj��l���$�!��CE/{�&܀R"O��WC�)t/���p����ȕ1"O�ȱ2�Q3 ���U
;-XQ"O�t��g@�IO6EqF�J�s P�A"O��b1�M�bj~0iD
�/L�a"O�e��	(3���c��1���1a�	F�OƢM���,4D��q�<p���P	�'(�pe"��4�4y0	S@n���'b��g�S�'>=s���:��=k�'r�l��ݶD_vѡ4a��)y �S�'-h,
�#� OO���Ĉ��&�F%��'
��8'K�<� @۴jֵ�ReH�'��]#G��#'�,�`�:��D[
�'z֡z��d*�]��Ѩ.+��(�'�(����<�ʝ�ժU,)�0$��'ȦqU#��N����)#���'��A����VФk�ԧH�:4�'
hx,��_����瞯K���k�'%����Ò�,8�[��υLeĪ�'�m�KK91�]�����=��'�:����3���n�x����'���c%�AN�HK2��\p�Y�'��]R&���2���[" �Hh(�'�<���=1b^�#&c�#c���	�')x}�oM�?�У���*N6:���'bV��wk�Ht�4��h>H���'�ⅈu�ÃBz���$��3��+�'��8I ���!Aq�ȣ-�N ��'�� �nØm���Q��Ǥ����
�'e�
A��$W�
\�R,C�[>͈
�'�h�gI�"&ƅB��ǥ����'����W��p�j|P�hg�ё�'מ}� ���h�̈�ʁ�jP����'��	`A��:�H;珁�5���'�����.�w��%��e��1Gzm{�'�U!�$�wߚ�a�+!\����'p�AE���4TD�_��!��'9n����K)�2���1w��(�'����ĤʅT�R���g^��5��'`�,�U ��PH�M�6��V %��'5��
a)��%b�Cz���'�JI�&)��(��ٷ|�.Y�'�6\QF�H=e�$i&�P�_�B53�'��%�BO�O�ʨ�Ԯ�1%'^)��'8��s@��R�x�J͇'J ��'@��93��k*��R�CJ�Mu(�y�'� d�H���3�C� t� ��'��-��-�;������$4��uI�'��\�5��#N��K$�
1F���	�'��LPO�-`!�D���� 	�'Q0=J&�ޯ;1�L����ސ�:�'A�d
[!:�0y�RxI�L��'����� �C��I��fSe|��Q�'��H"�Bٛ+_� qF�"]3����'Y�)bڮ+!vYǦ��O�N�;
�''L4[S�]���p�3*:L�<���'|��0��~���1Fh�&&Y��&��� �n�&dg�-�GD�5ID�p��S�? p O[!q<���-��l��\[�"O�)#c��$p�@��C��V�V�QS"OH�X�	�$���8i�bui�"OJ�಩�<:-L�k - +��{�"O�܋������0�W�8��D�3"OBЫR��%pHQb�J��|S5"O&����-4Bh�l��a�T�2"O��'�&B��Į/eٸ9�"OH�@�V�(&��r��r��`��"OPMCd'Z#���yu���k���2�"O (
��)�`�a�R�|l��v"Od�t%˂.����[�y�8��"O�TK�Ń�\�l1�����: ���&"O�@`�/�0(��� ` �n�2Y��"O��Y���ek5rD�_�>,��"O@ՙ�&-zȾQ���U$|�f��"O�|sr&�O�ʠ:W��8Z%"Of䁢N�
& D#DF�f8	�"OtU!$0T� ��#�->Y!�"O�I����b�|����Q�D��`P�"O�@��eS�9����̐��"O������DH!j 2�0�%"O����%�h.�v�����f"Oj�j�=%r,tX�M0s��lb�"Onl&�p�@��z��-�D"Bc�!�H=u��(�V3o��Ɂ���t�!�DܿZ  �T䓽_<�A�ˢ�!�_�n� 	OY\Jբdk�J�!�d�J����,Z���@�!�!򄔬q"����̌S@0(f*J �!�$9�b@aݸF��{�)�0hU!�d�0	��e Tk8s�.���/^!�Dʌ�RM Ϛ4�:��E!�dƚA�rl�� �"S❡A�G�=!�d�(&ą��Z~.���cbT�3!�I�Q�$N�)�ɧ`ܻ_(!�$��Pn�����X)�a�68!�D]=,RI��X-�~Qx�Q�!���ya Ey!���,{�( �i�!��J%]L�&�O�4�j[v���w�!�d�,+���EQt�$� �B(r�!�:#���JI��3�0 V �n�!�� O��m���W�5&�`cR Q�}�!���L5<�y�ɛ�O!>y#¯L�%1!�d���p��5��f�S
 !��Гp�T(��[��@��C!�dT�[��h�a�\.$�����	X�!���p��pˤѷ'����O"6�!�zɮ�Y"��&>�����d۶q!���i���Y&f̘ܨ|"�B\;!��1^X<8��|ӎ(�=x��;@����*̄R��¥Ln�DQ�ȓqY���0dL,8������=��X��2������N���e;Gi�2@>І�L���鳍��@� �퍯V����Bx�cըi2��gK�- f��ȓ� )�D%
�g�P�*��_�Eؕ��x��L�5滑�b퇸�$��ȓF��1ū�1@��̛��U3L���CM����^=4܋�P�JlnU�ȓ ������ۚh^$E(3Ŷt�68��^���в�ަwE�H�5)X���]X�0Pu���\�|�X�e4y�	�ȓ`۴� �`ˠ{: �CDѴ.��%��S�? l,����mHA����3_����"O.4�a�P<+~�уCG�0Y�h�"O~q0b�|p��3�G'=tb"O�P�ԅ�"��Q�el�2Xr�5�b"O����J&VP�%�&�V�P�"O )�بD�1R'�@.��C"O�4��.F���i�&: �$��"OB�7��%k�EQe��<5�PAu"O��9�n\�M���拵&��XD"O�a��=���"���0}y0"O8!K���YV E�%&�"|��"O6���(	�ld�`J���x��5"O��R��I����m� /���Z�"Oj�c��ڸ0�ٳCl����e"O�c��˴H0���D��'�ir"O�P&h�'/"�t+��U�L�@"O�5�d%��P����dCҘr�}�2"Ol���HF�M+F�s��в2�|�V"O�TA�ԕ�f�h�j�4)��,��"O�E2u�5 ���nۊ�*�"OV ����W�Bu����0%ͬH"Oh�1��оe����"2)��ʲ"O2����#u��%�(�l��""OPq)�/��zD�k��W�$x�"O$Y�`��3��2��\�p�x�"OZ8����8T�$+Da�/��Ѹt"O���\li��d k�j�["O�HK��B5�����ݲlkB�Y�"O�Xz$�ޱB�=+���06g�DI�"O�,J��	Q{b|��%eLJ��2"O�=a�U�V�P����Z kI`TQ�"O�!�t�M=h��48��'7��Pe"OF�h���&LdF�B�G+.H�W"O ���[/�����y���1"O�-[T�J�-ku`���-��2T"O��+q�I&t��Tk��O:(��� "O�ٲ�?k��L��i��p�0�b�"OH!�bǡy(��I�߶G�^���"O��avH�8d4˵FH-{cޤ�"O����M�Q�H��Rd��	V"O||0&,oc.���=[�
"O8���-F�X�ڕ� �Є@4" y�"O:�S��!J~�aw	�J��9j!"O�j&�
��Pq�ш��=7"OvyBՎ#V�6���
Yu�!K�"O@����ժ2<>��Ǚ:N3�"O���n�"���GF��?<�$ӷ"O�|z$	�3<֘]{�d�8n�`�"OL5ƀ�8�"�a� �N)�"OR|��+Z��ĄO��"""O�P8w��u�:������L��iU"O|��`ߙ�ıaǂ�/	��r�"O@�k�ى9��0 �%G�@	Q"OX�����UkdsV�Q�c8,8�"ObT�H'`\,�P�̾�	c"O����*-����]���0"Op��6$	��̃��  �`	"O��񰩜�2|:�)C��7Bօ�U"O��@�>$�}�����h�^��6"O6@"I-=�,��`�3Q��\:�"O
`�!�F8�d��	69��AG"O$���%kg���A�֑R-z5�1"O
%��o���X���!5p���"O�58W*Y�5�xȖHH�eH �v"O� �A�1a���H��bi�3�E�G"O�3��R�6i�3�&N�`�#@"O�y��>���ڏ"j�`�V"Oh���#ƺ]���c��U!p����"O�@4n��2�� �5k�+�"O��T��D"��Q��Ӕ"Om)%��.��'��0lnx�"O���,�!�.HR��Ę�`r"O��STo�6l<XSG�J��Q*�"O��� ��]���fT6U��y�"O�}��H��qz��˕�Q!U��"O
D�Ңd�����@�t&�bG"Oδ�V)tu���&���5D*��u"Oj��A������d4@�A�"OX�b�m�"K.�0p�@�2q��0A"O����	;rkFDhC f^"3"O�tӶa��"���Ф��f1.�x�"O��
P�0cx�x�B�l�I�"O8�R�Q-e= �
d�X�'�Y�&"O�4[��X|G�� �`��{�H��"Oؑ[    ��     �  a     X,  �8  >D  �O  �Z  �b  �m  y  O  ��  ��  =�  ��  ƞ  ;�  ��  �  /�  q�  ��  ��  5�  y�  ��  ]�  @�  ��  p�  � � �! �0 �; C ^I �O �Q  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o�`iF�@A�p �O���D�{^h�����#W�`ł�`�}�:O��d�i����&.K$0A���a�=!�䅙�DЃ�a�>F�����&.Q��2S�"�n`�`�K�u��q����g�jB��ZɢJ"|E����ϟy��C�I;����ES������F�C�	�ݴ<(��3(��$�Ш@'*��B�	�=@�p�D� .X@4�Q�|/�B��w�
���!:f S�Q;L�l��'���Д���,$\�I�c5J�I1��M�I�͉���6f�x��8�y2 �0�4m���%)�p�3ظ'�ў��f�h�˓(,Lѣ#Ӣn��W"O
����3f����fV���2"OR�H�IU-]�@TR"�rX�ɳ"OJ���g
�.���;H͒Q��`T"O�QF�*���1��Pg����IX�O�*b�I��Q6pJ��T��J�'.�p�Ōb|���m�~��1�-O<�=E�� ���V"9W���	�C�,n��x��"OYz0���&l@�B�D�n�K��x��'��US@�����9� ��_(ҭZ�'߮\��$P�E�"됧IF�Y��'c.4��.�#p�������8���hO�a�B�&X�؃�ПY"O�@�JS+*�`�	�Q�z�"O(t( ���@�7?���2*O���!ϝ*���ఀ�	n\<�I>�	�CH��bj<1�B 
 ��I�1��a����<:A�9�RgD�)VNi�5�E!��(V����)?�0�R
I.K4в`�LPgax2�Ɍ^?�G)U�&e�%���	^̾B�I�H���T�P
u�{ �M�I��K�R�Gx���Ɵ��@{�m��A�,|C���/!�!��K�Q��4�h�É�&�1O,7�7LO@5�p�ݖ#��p;�b-+� �"OR��M��~��au�����#��3LO�QB��+3xu�5���H����"O�q7�_=M��0���0��U�5"O�H�o�(s9�}���	"����'��iDx��\<�B�%e�T�p_��y�p�����d�YŲ!I�'й��'�ўb>��GG�5b,"��f��{B���M5D��z��ˁz�k0��"<H�ı��.��j���q���1L���j�w�x��1�,<O�㟼zR��St[�@ܱ77����E���x�ҮN�̒�oT�*�V�g���y2��&M|��H����MO�%����yR���'L� ���/<�=�Ǣ��'k��b�Z7-�<iS�?�@ւ�1Dk�)��G]�sI�Qu�>D���Ue��C�X���/)U�0�34�(ғ�Mˌ��OՊ��e�ɨ 0����I�	j�
�'�d�6 O�
��T'O�{��h�{��'5 |rFkF,o�୨�=r��%�'}0ٺ� H��I���X �}�	�'����a�7J~i �8Vn0�:
���y���Ydb�j���*7�r��j��yr��;��pT>U`H�t�Q�p>�K<����$u��K�>R"Iz��X�<����t2\E��A9 H��2/��'�ўʧfYڽI"J]�M7�1aa��
А��ȓWK���,E>�ՠ%Yr�{��)��ф �)��)akē Q�G����F{�O�l�<���P�s�a�Q� U<~�A��D^�<1v-����ǋF�1���PW���<a����DV�_L�x���OR����Cٙ>� ��	}r��B������P ���'�ў�����#e̯S�dYsW�ՐNUp��t"O�Qp5�>��*��ǥQ�F̸�"O�l*���Q��\:q��_���V"Ol�2gm���%�c*��"�T��f"O�m�&!��]t�a ��)���g�'$�'��@�i4v�8�ó-����	�'u����\�R����Q ���R�b�;�S�)S�j���%Ī
A�8Q4�9UD!�d� �ġs� ީd;v�KC��t�!�d�	D!��#4�Q��A"O�!��×8D�H����&�f�;�!��,��`��L52zȳb��L�a{��D�#o����B��$k�``Aφ8:'!��0T�ژSԏF,Wbt+��N$c�O�=%>�2�o j��A��,K��Q��>�O���4�+��$(lJ���W%�J$Dy���� �B�N�,5�c2?xMSg"O&��@��nkX�uMMW1��s"O��r�-��G��[��% �͒���(lO�i3g&W 
t�[d�/[�,X�"O&l#t�
<Qf�	��J��p��q�"O���R'S�w}X)�R�Q�P���"O8A�v L�������Ԋ.I�@�"OB+U*w6��k�!ڏjAD��"O� H�N�-x�ք���G�\�Z�'5|9���
������V.H�T0���<O��ʔN�
�LD�`͌�xֵ0"O\P
�B����@�µ[z�E�»iš�֗D��}YâY�J7<q�"i�3+�!�$Px�r�0ҦW�640 �H@��!�đ�~�����U�8q-��T��O��GzJ?�bҠؿ^]´�h1r��5a2�!��mڴ��CS�~�� rANSf�G{��9O6�S�l�(c�d�k1�ĵ{�8����'��O4S�Q��Y� i4���V�'8ax���b'��=Z��b�H��y�T�e���!)A�;����AW��?I�'�}��S!(Ƈ_�08�<*MI���'!�h%?�)���2墅��k��He�0y�0�O4�	"1�J��t��l	N��j�ޣ=YÓv�Ru���u�l�ćXMaF~��%(���˞��|���'��`��t!�DBZO���$��5N��˂�Z
Up�ɥ/SQ��|�%E�H͐�"��KF)!�cB�<Q�[0t���0��ܐr��|�<Ѡ�_1(X�Ң&��ј��D�<�S�U��>�c��#Y_8��RK�j�<q��*9F���4=�JX�D�b�<���1���P!-e2��ۅI�X�<1$"
}��xV� oڔ�d�X�<���?j*� ��Z�^-a1MY�<y��Օ]1і�3~<Q@�^�<1�d_�?av�����3��5#G�Yv�<���X%T,����E�
q�5�2!o�<����rW0H㔯�Z�2��`���<�Ā�s�
�C���Qrd`��[`�<�b�,$Rcb��9��X3ã�]�<!!��7��1VeQTy�L�f#S]�<iƥ?dp��՞q��v(�Y�<��O�
���eBR2h�B��R�<1���4DB8%�CR�Uz8R@ćP�<)�"ǙpP���=%wN�QcF�I�<�wE��H�p`�D;Gu^5YP� @�<y®'F�@`��̴(0�����z�<��+��;���gS�hю�eYs�<�G�f_��0ԯ�tf��ȑk�<����\*��P���=�6��OPs�<1�E+9lL����3]�L�{�d�x�<٠�@#X�5�.[�*�4��x�<� ��
CS��ti�1"X��VK�s�<��iC8*�̠JR��;���� /�q�<)t��|݊�[�s+�t���k�<����B���@�Jz���!�Od�<�A.A2~Lb}QWC5�D��B�KV�<Q�	 +Fa�礎>SD��c�S�<I�
�,l)�r���h7��Q�<���W-kre���?R�でSQ�<�f& 8^�0��.U4W��"7��w�<��X�(4$��o��е
��k�<��	�,%��EaD�3� ���h�<� �h5�ĩw����P�_�A.�ۗ"O�ar�A��D����� @���"O��Gm�.� �z�B�.{'�*P"O�@��.��,Z��L��Tb#"O���B~�t�#0�º�$e)��'���'Lr�'�r�'�R�'�B�'�Hˁ��=Y��� UB��)�x�Ѓ�'"�'uR�'�r�'��'�r�'K�1	��g�
�U'Ѻ5�\(G�'O�'-��'�2�'�"�'��'|��P-��(��}�,4G$R�jt�'�2�'��'j��'�2�'e�'�T5kGn	�zp��I�`t2��'�B�'*��'�B�'�b�'�"�'��89�i�[�d�3'��|��Q�'��'yr�'Q�'�b�'�R�'���5M���F �С��R�e{��'���'b"�'Sb�'��'��'�|!��hE�m�T�b$�=y��d���'��'�"�'{��'�b�'b�'�ڌ�UJ�X�akd�Yy�����'R�'�"�'T��'���'p2�'��뇸0��y7��OP%���'���'���'��'�R�'ER�'��A����#�^� �#^t�d�'>2�'���'���'�B�'��'0�����S�1�ԡ���ב|�ۆ�'"2�'G"�'�r�'���'"�',�AH��$`��R�Y�^w�����'���'"�'���'�b-y�n���O{ō�=��q�1J�_��i{�l�py��'�)�3?���i$4d��JQ/I������0���R@AC�������?�g?��4A¢=�7 ���j�@�=��4�i���ׁqD��O�͂v�	�'�-�K?M`��O=,Ns�LU���E��E7�	ʟ@�'@�>�q��)N�R�&�o���u���M���ZY���O�07=��m�Qg8(9#>C
�D�t/HџdoZ�<�/O�O���J'�y�(�'�n�p�#�?_�#@�R��y"�ֽ$j�$Y�%�7�ў��D��)�tO�	��D/��Mq/g���'��'y�7M�v 1O�����SIU"%i��tP��� b(�	����O�6ml�t�'h�5�D��d��Ф������O����T*5�y��I�+6I��� �Od����
j�*���@��Z)l�� o�<�,On��s����M��6 pPئ'����<z�'|�$��4یt�'�x71�i>��u�èZg.YiЯ�{���ԯ����	æ�	�;�x��u� ?�tOƔ��
��g\&@ä��,�l��Vo�6|&j�{N>����?ͧ�?)���?���?Q$��6�`�̑.Z�<�r�E�>������4�u����4�?iK~��'V:���:��#���N����O&�D{�"�N�S�?���$_R� RV��'0��\�ãyo�E2b�Z+fJ�P�'��M�G��0A��U��|b�'�"`ˌ[�>}`�Z�3� )��><2�'*B�'J�O�剷�M��F�<�Q�X<�l!��C�u�n���V��f�'Xџ��4q��v�'s��cqgZ1��� ׃�?�f`*1h��$R�E؛'�h���3�1��I�?�QZc
nl��@?�(��f�F2=�@j��'LR�'��'2�'��xz$�fUR�����b8���=O�pm����4V�*`����>���)p��4ȗJ�6s*2��Te�e�B�D�C}��o�&oZޟ��G l�f�����8���(�$U3�*�8z�L�Q�cI�	 pH��5!�2�&��I����Iџ�	Ο�!�#GK4dqC��
���7��؟��Py�x�&�R>O�m�ȟ��OaT������r5�7��?�$����WЦ���4�?a���D�Oe���@L�5�X�"$B�kfZ4�_�G�&��!H��!���?�Y��M �%����͒� �6��Pn�UY�䚳N�ş0���p���b>	�'3�6��j�(��]���)�E	JY�50O��mZП�GbHjӊx&_A�9�AbÉl��I��
Ŧ�����(�-w��I�~D��!·�@�'��5���О(D0]�
Y�E`AR�'���ꟈ���8�	۟��	R��I�3�� hN�!�:Hó��K��6���D�O,�$���<a���y��ë4�fɰ�e�7*�ڀ6#��? 6���i���4�����Q;W-/>󄀠SX�Wi�3o*������d׬5�9���r�t�O�$�Ov�d�O�`����7M��A�:)j��c-�O��$�O&���<ɧ�i�*�'��7��O�Pz�i�*}Rn9�2 ��@
j5#�(��i��vI{�
�$�s}��bD��2࠽+T�9��Γ�?i �Ÿ%R$d0��+��⟐)��D�7���D���f!�����Q���&g�����OV�D�O���0����l�Ɉ�\|ّ͘�hZ�]Ǝ�$����M�M���?���p.�V�|��y�D�'�Dh:��
1N��UPr+�)�y2�e�T`mZ��M��/��O[ X��?�ulA�{��c` �-L�q��8s ��:��2L>+O���O���OT���O�-ksbPU}bas�C��6"�0�P��<Y��'�m3��?���ZROR7�򉇳4��T����Nf0���X�P<�'d6m��)�ڴ��'�
�'a�,��E�C�>�ڂC�l^��'Ǟ2� 1.O��E��m{�p@���O�ʓ��D�ܴ�Z���(4c��z�!C�:l�D�Or�d�O�YS4O�O>˓ ���'E�R��E�l��W`E}�0��딠�B�c��O(���M}b�b�6�nڦ�Mku#āhޜk3�?ob�JVl� Q�2�9�͉�<)6�L!H�z0p����j�<c��RTLD T6k� ~`����*HVIʂ.�g����4O����O@���O<���OZ����j���!e������/aȊ@S(.H���D�O����̦��hߟ���6�M�����Ę>!�6f�xĎ�s7�' ђ�o��������ܴ���F̵C~�u��?ᦏK +�&���.W�4Q$<��`��~6@���Ǌx��%I���<A��?���?!`@W�e��ː!p��DP�Ըl���������1�jTy�'H���wlv�ZU�|'0P�KOo4�Q�''Bl�>�5�i�T7EϦ�I|��'j��ل3�@�	�NX;+夕��&~�FX��^�����{0W2Pu �OF�Jt���O��d�ƥ�&��1b�O����O����O1��˓��F��gF���e�!�p�� ���(�[�'g6��O �?!Q�i����Fh�~`Za��!��q@5g{� �$�,^!�\��5O��	�x�T��#%r��^�@L�/���s�*ށR�R���f�ܕ'r�'!B�'�R�'`�S#R��c K�y�=����``,\���yB��I� ���?����T~��x����$I:��F}x���J.��nZ�M{b�i=|��|
���B���0.��ϓl�6��6��"=��(�G�#ӛ�'���(P,�7&�h�u�|r���M3��?��"&T�@p	2J>r:��P��?����?9���$��E��#m��cݴ�?٧��I(�|R���w���ñR0��O��lZ �M���	�q�:h�j��l}ʡY�'��b�I��(ݼZ�:\��	�iy��OwZ�B2�F1T�2@I�wz��1�F=���*��_K;�'���'!R�����r䋀];T�:��
�0Ͳ1�f�lpܴK�~L���?qԷi�O�Lm<JQ��hŲX��]SS�
������4Jԛf�˩hlFh+�'k����4+ ���"~����#�$L�h���
��L�0�|��'�"�'|R�'zB�'r�<Ul��A��>i�KF1Ii�b,O��l�\<���.�M����JO~"�a�$9����Õ�R\�"C��N~��e�
5mڟ��H|��'�?��!=�:l��":�L��q��L����\i>6�K��J���O2�D�Ofy��G[>	�p��Ij�[K�O��D�O���O�	�<i��iX���'���QEgM?*G��i�h�;
����m����(�%����n�Z�D�%�:Y�UJM�� &�_�p4�ٰ��_����O���#J#	�2IW
�<��'i�k���N	�&�ә9VvxHঞ!g���OP�D�O����O&��7�SoÜ������z!�4�`�Ǜ)�B,�'��AeӾLaw"�O�����]$��9��Wz�Ǆ��!9lx�rMH��M+�Z����4wH���O`dI� ��y��'d��Q�jc���X�f�!L��(�h�� -�ј쟝-�'.�	K��K�dC�a��}�# AA�Dx��n�,���O����O�'%��l���%���"�柚j��q�'*�z���fӠq�	e�S�?Q9nJ&�����A�]ŲdI�,�Sh��P%#_ZIF��'�Ԅ�Vq`e��'X�ɛx��m����'|�!��7M&l��ޟ��Iʟd�)�����s#˲}Wx���jH��%�<0'�$�Iܟ0�ߴ���|�@]�̒�4%�rI�B��4>��dǗ�6}�!�i{R6�V)�,��u6O��J
z��}����w~��?��;wȊ3 �dE��LP�~��̓��$�O��d�O����O
�$�|�^����S��K$!��H�E�,,4�vd��2�'�R�O>����'A�
k���[�k�,|���ZX $�+:?y��n�-�M;��i���|�����S��9I���͓p���ecO�J�"�Ğ(QPp�W6ʈ�0��DL�O>����?���?��B�
�<-V+�{�H@�u"]��?���?Q���D�����E�g�|Zش�?���X�(|��$A g�"��4�����O�o���M�Ia���
rH�c�P"�ظ�h�*
����D��\�,��)@y��O�@]b�±K�A��P�+�.ꨑ�U=E��'���'mr���b�&^x2�'�bl�����M�T�ķ.+xY	E�'�7��a���$�O@�lğt����w,���.��Mk�!��R'�<	��it�7M��}Y��T
@<���Ο4���<6���0��^#~���C�%�l3�h�z�5'�|�'���'E��'L��'JI�������Hr">l'�ȈcR�L�ڴc��y+���?���2)�@��['XLUaŁ/	�bEJwlǴ%w���'�^7-
�ш޴u��O��t�OvR�s�m_?K�D��C@�
uU�	!5�F�)���z�^�<��eՀ�t����k�I��h�	5[Yʹ����o�i�c��#�Q���\��柸�i>��'��6�	>���8;�Z}��E�8+z��` � �0o�蟰D҅n� Pl��X����+�~�����>V��1/�6<����t���I��UY�K�)�~ݕ'��mz��Y H�t��x3��@�����BٟH��ß��Ο���˟���! ]8�h�TDP3rc�	�2	[�<2�i���j�DI��2O��'��'��Q��D��Zp��Z��Q?G8����hN�ɂ�MSv�iTB��I��d��'����,��@�06���"T��ȵKGMM34�� �e�N��֟���Ο�������ɦ��=Q �
/P�h5ȱ(��i����ݟ��'p�7�^�t�����Z�t$�	ơS��ہ"vΔ1gbS�OL=nڱ�Mk�މOj��H�U��8�G^E�VYK&�Z1x��82L_"S�ɘT[���Sq��@��f��c�0��k �v�d��l�Xz�I۟��	ٟ$�)�SQyF~�*)f�U!!1bM� �Ä�0I����W������E��_�'�6E�����#�C���N��plZڟ)1�?u��	䟼!�*� �����bly
� L�é8M�Tb��k�ź�6O����O���Or���O��$�O$˧*ł�	�J1(%�O3)O�py�iQ���'F�6��M��'��)�|�;r���s�*C�A!�`�H��%��"��inv7��O�֧��O�r�3g0N���'2a�䃘�}D�7
ӍNuؐ@�'&��L�#[�8���|2�'���'-�-��1M,%{r+X-%�B��u͗�U��'�B�'�剚�M3��<	&�i��	�x�a� ��X0�W�"�џ<k�4��'|�_�ݣT (�=���]F����?!�b��ZW�PDD���`<�c%�>=~�d��-��#�>�Q���5��$�O����O���4ڧ�?QS�Q�xpJ�l�4Ӭ�+6��
�?�iy��;�'��7=�D�=�v�Y�#�^X$�0S@J��i��<9q�i�"7��O�L��^f��d�Od�F��?B���,�P
R��0M��*9�U�� u�O"˓�?����?!���?1��,��#��D GF���ĢOK",�+OH�m�&W����IܟP���?Mz�������-$��e�P���D�j(�6A�/
i`�J�O$`n�2�M�e�i��O�4�Ou��[�w{|
�_?h=h]H��0-ڼe��S�����H��xӖ̞^�ICyb\����VJ[�Iz\RQ�L���'���'2Y�g�'��I�?1�+���&]�Y���;�OѸ>:��kA͟��4�?/On���l}"n���o��M�؍�44��i���Ѕ1bkW;�8�K�<����J������4�(O�I\��3�̚#ʎ\)�+��\���b�@8�?1��?����?����?!����K��@Ƞ��O�'Bz��$��y��a���$���&�f���OX1O��(�E�X/F�riK�JId���'X��;J�fht���
K�:�*"4OR���=`I~1��̓`�x�9������r�*0�8/)K�Y�2������@�}�*0�e�mx��� 0��"��J	��#AϱbA4�۔�B:��� �g��n̊U�Ρ{u �#���~aNIˠ�G @��ҖeŵPr�k00�X�R�¬�VL�� ��&���c	7))2��MG f<��rJ��,� 3R�F$��� ��2��ѱօ�)1`��t�;��	���])�9ф��rS�`B�.I$1pU��Y�	���-"�FiIS�I*��.��m����(,��0H���4a�N�Y�*4qE�{��%*Q%s�P���O���Zir��L�@��y���I�#J:9H2�q�ӟp�ɉP���I��������S�z�\)�D��27���ɷ�� ~���ݴ����<QR�o�.��I�O(�)~�^TC��A�=pq�����M�(O�@YS��������6?)���c��$Q@"j�~q��\զ}��������?=�J<�'�xq��C{Pe�fȎ�y�i
Ľi|�+aX���	���3��꟬�oWwDhb@�5&!�ՅO�M����?!�>~�iT�x�O=��'rh5P�73ve��ʝo¢/�>����?9�O�j��?i��?(Α��2r�k�4l��䛑5%��'��2��5�4�����O.��D��eH1P&Z��g*r>H1	��i�rǙ���'�2�'�R^� h�*�D�
)��O@1G\�4��^�vO޹ZL<I��?a�����OR��R�~���r+K�p�FɁbh�#^\c2�$�O���O��C�J�9F=�z 2ph�!<�j�'J���_� �	˟$��Hy�'-�n�����t{�� r�6c���q���ڟ(��ß��'����f,���	����|�����Oýq2o��t�	Vy��'�b��ӘOń|�d�8.b�{�R|���.x�H���OBʓ;rzPr0����'��\c�<�R"h1aohh��c�$z���4��d�O&�DܒN�>��s��+�
V)N�nY��*H�A�t	ַi$��9�>��شJ}���L�S����Ƥz@�!kT�H��Iز΂ 5e�F�'�b�
�%Z�)�g�Il�n-0���S0� R�۬U��6��t���D�O��$�O���<�'�?�t��� �`�)����S$c[�lR�V��: �{�y����O�l�h\�jz�)!1��W���	Ӧ��I�����/
�q���D�'���OX��Ȏ4v@�(�E�]VX[�k
@̓9�Y�V����'A��O��F��L4���?`Jdj��i��/��A��	ɟL�����=)�A=xI@�U0�`5��H}b�LQ�U!�O8��Ojʓ�?�E �5�
��򫂖����
fRx�+O��$�O��D-�	՟(;�!�$8kj]XD虲3Cb��!æ+n��yDI)?����?q*O��:v4��;bs�}w���T�X�i�&]�6M�O��D�O����y���ag�Ru!g�˼�jA[c%݁RG�]��IП�'�� �oj��ʟ�3��߲�1%^)!��(����6�M����'t�$NZZz�M<�B&Κ~P���(#~��5�GbRঽ�	`yR�'9��RW>!����t�S�5\<UBrKN¥�V��S�qi�}��'T �c����i�Y�U�χE�~]+s)=E����c�%˟���Ο����?���u�&��Tȍ:FMO�p�b��#)� ��D�O�(��6>1O����EK�x�c�CƆBz����i���R�'���'=��O��i>����(]�]�igxi�Cn�;3�|!� y����0Ӑ2�1O>���0f�\[�BE�;.u�C��n��lS�4�?���?�TJ���4�8�$�O���%T�,��厗���{w�A����y��05�
�����O�ə� �{�(ڙ6(�rs�Ā ��7M�O�*4��<����?i����'	��hgjX�m֢�˶��}b-��O�u�@o�	"���ş���Iy��'�� @%��Η	2`�xBGLx�"81K�����O����O���I-r���䋞�/%t�C��¤R�I�2�]47A��?!�����On��m�?q���. Eb=je�+�a��bhӊ�D�On�� ��͟����B4^#�7mDl�����q���Ѐ�K5��	ğ��	Iy�8O&Uj1^>��ɢ^.0���9t9�-�����5����ߴ�?����'��8E����SI�xЋʐCu���A�پ&h*�o�џP�'����#g��Uy��Ov<:��%�Zq(/RXи���'�I���
��W�K�hc��'jp�*���:"�sp`M6YU ��'n���X��'���'���T���6u<��2a�Խz���5`��GR듃��p����8�c��
ܝ���F�&�|��i�P�b��'�BT����Fy�OS�lG,r���Y5Eŀ	�ĩ �S�,��V���Gx����'�����*��/�P�A�]�i��\ZĨy�����O(�d�:�:��|���?i�'�r�8F��1h4Z`A�j
�d�`P�@�(�#hN�`O|���?i�'(��'Z
"�`A5�I3iъp޴�?�p؝����O��O�����K�
I7���(Y;e�9�7�>�ӧ?6�%�'���'9�ȟ`�G#ޠ����@΢u���&H�W��I�'���'�"�$�O���u�D�N�nX���<	���dIT�v���Ò�L���D�'5�L�����������W�t�IuI��}���'I��'��O����=8��i�2q�0��,n2��і�K�J�ةO:�D�Oxʓ�?�������O�PX��94(>`��o�G(�#�������C���?Y�HD-r��'��׃_�y�|u�w��8"f�y[G {�0��<9�'6��)�����O����!�J�
�	I�>-�݃b�
��t�>��<,��rċY�S��ϖ����jQə�zͻU���w���7��OJ���Oz�D�Ӻ��Qj�!�.̞x}r� }}�'��z��K�����Oc�9��J͟�v�V\�L�b͊ߴbϜ�����?���?	����4�d��v53я��O�5����"0Po�qH8���!�)�'�?Y���
|�����b��l��C�DE{.��'��'.hr^�������}?1����7�^ӂ���^� 2C	��,�1O�J�^�S蟬��k?ѓ���X�r�@ET0j�@M�%���1�I�̖'LR�'\2� Y���,�$r~�q��!����5��jd(?���?q/O���4>�Ĉ����3���aܳW'޹�� �<���?q���'�2M�!_��d��T/��*���9�������'��'��˟h�ՊN�E%��\�Ȑ�K�,��j"l[ЦA�����	g��?Y"��+���n�v�ΰ�+S�<ܵz�B�e���?�����Or+wg�|j�Ug�Xq��
]0�Sv�ѽ�\�h�i/���e����
9�'ɜ@Z�-��"?j��S��V<N�Q�4�?�����W@��O�2�'*�hqbvm8`f[+L䨼�ӣ`9�ꓳ?)���?�h��<	����D�?A�&���R&��E��,m-)rKx�ʓl����i���'��Oh�Ӻk!e�oN� ��_��)b���)����;��n���	ҟ��Iܧn!lس�, F��KD�R� x| nھ s�I�4�?���?y�'���?�����.X ~��H�E�Q�Khz�s �i� J��'�bY�����'7¹i��]�����'�6��!#G�ڸn��4��柴ïB�����<a��~�ɐl��Ə�V�z�q����Mk���dZ�Z�Vl&>�������l�<i˲�
F���j�$��]�4�?������'!��'��@�~��'4QY4$��Z�V�`4fM,F�(q�O�TxQ1Ol���O��$�O���|Ň��88�	��}����GR�rl� 0^�80���?���?��Z?��'���(V�Tv�ܰ6P�X0ES�/ �p�'>�IΟ������Iԟ�k'
2�M35 ʚER���҂*{ R�C*vY���'�B�':��'��I͟�3�.y>7�Ȕ?��|�B ��iA��[S��!.w���'a"�',��~b5��B���'Ur�Y�g<�hp)�=KXP��H�p3�6��O�D�O�ʓ�?�B����$���J�#
,Y�ы�BS��y��Mi�����O����O*��rĚԦ�������I�?�����uw�Q�&��N�Fe�b�&�MK�����O���=���$�O����Qါ]T,L��=%0q��b� ���O�ŉ���榹�	Ɵt�	�?���˟�;�kڍet:����)�^p�c�����O ��3��O����O�˧��Ә_��]����f{�0 t*ϱl2�6��9��oϟ���Ο��S�?��I֟���0~�܄���K�� ��K�^�B	pٴ5�������?��*.��n��Ο��#bݰsm��P��:r#t���M�<�M;��?�:�r�Zмi���'�R�'Zw����uk�7X���vH���ڴ��z�2H�S���'�۟,�r���+EZ���S"L���tRдi��.�L6��O����O���I�4�O�,�r�����8A�����ȅ�q��f�'�~�ٟ'V"�'���'�rU>U ��%x6d �ц�7�:<!�Q$���ߴ�?��?y��?���Wy��'�$�WCN\ 9��)m����P�R��D�O��O���O6�DЁ�Qn9�ƙ�֫�	$4���B'5����ܴ�?i���?��?a+O ���fT�i�5���#3�P�gg�4)�@�
��m�����	ןl��@yG��4���'�?�q�? N|������H��� ?s8Ƽ;S�i��R����ٟ��	]r�	�����>��
$y2|A�%�W �0n���<���`�I�=�D�ڴ�?���?���B��;��d{.$q��I�d�����i�rS�h��7U��ϟ���P��4:cfX 1�2R��
҆_�_:��n�̟<��8��Pڴ�?����?1�����f�TI��ũ>̉2T�QA�)�X���	'%J��I蟠���$�~�R����:R�ޖ_d]�dD]ۦ%��mX��Mc��?���
���?a���?�る�OO����+.P�%����V���=t���'S�i>&?1�	�'��ȇ l&ޡ��.��u�X�4�?Q��?q�᜽oH���'���'���u��T%�!]�	�I�&�i��'b�'�"�[�����O���O�(��ˁ2Vi\]�щͅ_|H�+`I�ɦ��0�&Q�ش�?a���?��B��\?9�����uХ�	�2o~�ᥜD}�k�y�S�����P�Iϟ��I�V�493dI�[PiE�u��ʔ����MC��?!��?1QT?5�'�RnK�
z�1�p4@��$�M8!)ШA�'����� �Iҟ��'֤@`lm>�g@	*Q��TZ�oƽ	��р$�>i��?AO>a���?i�A��<!��P#)�%���\��Z��C������P����'���0%?�)J&MS��8]��2�#F1@��En���0$��������oy�ФO@�s`�ʻ6IX���E�TV�,[B�i^�'t�,�虫M|j���`K�/�U*&k�7�����L�D��'n��'�HS��'��'����*f5��w�ì7�����.���\�������MC�Z?����?ap�O���j��>�X8P�B�t^���#�i��'V�b��'}�'q�"-�P=�����JD��i��@ls�����O����x`�>�PlI�fu,�3m���� �� 4_�Vo�h�O��?��	�:&���/U�;z���?[� �ߴ�?���?!���'=�'�$
)�RĹf��pj���Z���|�`�#k�������O�d�<Ld�:��/\�#�'P�_���n͟  �K
��ē�?I�������
&1�VE�ekҿ~ʮ���B�f}���}�U�@������	Ty��G(g�*-�I�0��-XR��3xi�&�2�	L$��I�����w�����}����oǓ.����@y��'s��'�I�~j��O`C$l���%K�H������M<A����$�O>�$�O��Ć�O�!w�O�i�:	ЂLD�b�BT�V}��'��'�	�R��)�I|�/KtP�-	`oS�9���3G���'�'g��'���C�'�{��d[�fU"N����� @m0Um�՟�	_y2��X���������d[c.I�#-�Ő�2v�T`�J�M�	����5�Iu��r�v*�r��c�B
Ճ��񦅕'��c�~�P�O;��O���6%��!f�>���·k'���'���|k:�.6����+Y
o�|�#B�B�D�h���i0�8A�'\��'���O���'��S�^�"��/������mZ�	�t!�4fTT�%/�D�S�Oa"�ۧh(���JK�/��<y�	�xuf6-�O|�d�O~��L}�Z>������B��;BTeQ�e+V��2��A�>�>���?Q���?�L�5c,�8�"�-���S �^�!���<:� ���'���|2`̴�Zݹ0�V*"P�|�eL��f�1�P�x��S~��'z"�'���'�At�GC��Ը�BӮ0����˛%C%��'-��'�R�|��'��AJ�i��$ $�7�h����G�s�\��vƑ�����O��D�O�ʓ����2�Z=#gNT&�"���ɉ@'�lq�R�8����D��[�UZ�l�Ou2�P��� !�芴�.>6P�O��$�OJ���Ol�D]abp�$�O �d��m�F@��A��*�5��m�BMn�П�'����П�2��9}�O6��$B9r�~
��I�&��C�iy��'@剨S��-ZJ|r�����߀QU�$S&�A�aJ��W�����'0�'�@ȁ��T?�)��Y@���d�=��!�j~�V�)_
�0��i����?1�'o��I�c),��a�yt��eǍ ��7�O2���t��b?E���. �W�
PpE���M��E�y�6�'UR�'��� <���O����B��b�aNw��t�c����yqs9�S�O���5J�ҭz�iW� ��x��$�6��O>�d�OySe$�T�I����I~?)T��B�Aq�SH������Q��l�|�	ȟ �	)z@C𯚱'NDB�f�<ڴ�?��^�4K�'�2�'yɧ5�Ϝ� O6����NHT�	��C����лQ1O��D�O����<�%恧n':��&��~�p,t�L#���$�'�R�'5�'�B�'��G&#+��c�7%���z&�7ݘ'���'B�R���%�*���e�1��y��^�8= ����ɉ���O8�d7�$�O:�$ыg&���Tm��l�(u�pY#K�!z���?���?�+O���B�n�:U6��T�@n7�r���M�h�r�4�?)H>q���?�0�]d�~K.�A1���ٻ�V8P��l�ɟL�'�bLM�"������?��-^�l��]�` �,w�r[VJ�ē�?!���\��c��I�S����=/�.}��؇h4�|c�l�M�/Ol�+����m����D���槀 ̍�U��4��R$��$�����i��'�d:���IW�p��BT�^��풦��)>ϛ���+)�V6M�O��D�O���J�Iߟx��:wr�� �C9K�:���oK��M�"�t���D�䞻�Z̨Al�F�J9���J�6`��nZߟ��I� X���۟�%?���_?Q ��=��x���t�kR�Ĝz�dcL|���?I��Gc~! �ƚF8�U���J�g�køibKˀ��O���O�Ok�;%�"��sm��NӐ] W�{�����	ٟH�Ixy��U��̀"����dXR.�X �0�$�O��$��O����V���a��$48U#Э�6,��w��O��d�O
ʓ|�Ršd4�\��-۩3��0��f��|�0��pU����͟�'����͟���>b�ʑS�E{�l�(�0��!xy�J�,i6L�{#��!����%]Ⱥ��&�X+NX)����C�ɞ"ib�`n�8w�#'�ߊFt8�	�s��ՑC���@�#�N<�P�WiZ7���{ �F�*���arIO�;C�L۠B�#	D:�F��.���s�˯;F��3#0V�<c�NB�;b�#E�9=,�Q�Ō�8 �|���`R�,�h�9�S�t7�H�c ,��i2�H&��4�C( }� ��hW; Pg�{N�d�O(��1mH�D��#��pY�eāo
 ]�]-��� ���42Te�f�~��
�}j�c>�.�3QF��;�@�*W� h�p2vRyj&��D.*5s�-8G�4���C�	X���!SĎB�l�ƀrda�*sR`��F�(����x��'��(u�}�� �>D�aVlJ�^���HP�܉���!iS�U�*\���Gxr.��|���"&�D��ͪ]�6I�b�Z"3ؼd;���?i���*7v���?����?�b������Oj]�U�>�(�+���!a���p2�����0���j6�w�����	�[A-5GR8�9W����N�"N��:9ǃׅ@Ր=C�?��թ7�ɦt��䔜T�J����ƀ���%���d�O�=�+O���	.�&9AW�W�2��"O�<y�$d��	��l@�Pn�yRw*l�����'��Ɇ_���y�N��*�l^��!o�\�V�����x�I蟈�C�T������|�����]�A�u��q�W�A|h��a)H� 8RA)���tꘁz���M���XI�c\6`�@�#��?b#���pE�$ ,�˙%G��%t�F��b�	�-&N�D�Ox8`fϬ����&�J2-�`	!���O��)e%����Ie�/@�j]�&"O蜛 !ǟ<W�4�c̚�\���Y30O�nZџ<�'"���,pӎ��Ofʧ_1�xa�@�9
�D +�(A�zm��t���?����?)�cS�t�> �G^);�D��nOB�y�J�9��5+��kKx$�'��URrPDy ʞ ��i"$��0\<x��A�#e>r�9���(Rm���F�A�Bթ�O�!~〔Fy.H��?IB�i_p7-�O�˧S�dШ$F�$O\K� ��ٓ��ꟈ�?E��'"�x��q��:��Q�fH����yq�'L�]�5C��\8�9�'�+�xi�'䀴��ӊsy2�'�>E���	䟰�ɘq)��IK-7˄�q �eb́��D

��lC�nA4�������6���Z�)�K9�"��� �9T$���v�E
Srd4�̟yF��Vd6Tn�PD��;l���(I3s͢�cP��~���F@���?���iT�S�S�?՗'{�0�t%�>Ȗ�3W��,rH�	�'%0��J�Dݨ50�V�n(�i���A�'(�7��O2A�g��'-YV]�@�O�q��-+S��O����b�F�jD��O����O���纃��?�W"�d\"%R�Q�;���1EߩLJ�ACv_�7޶e��L���ψOLSS��LPK�#�x�X��ԫH��C�W�Y:Ӭ��A���{,��:�G^�!?&ɠ��/�J��	=��DTզ�J<����?q)O��r��.���g�R)�L+�������U�`��͖|3��k��	.����4Uٛ��|��O{�U�Hb0�Z �M+�K��{]Ha�T�d��)B矰�?!���?���`B"=ϧ�?ٙOIx 0%F�5��|�EB&M��q�5��RArD�F��<��B��S
g&�����o�'d�N^��8ѐ�F@��@f�>,�x���6 ���`�m[�5��Є�m�Q���v��O<�l7\)�E�f
(F������#kP	�ݴ�?Q-O �D5�)��"\0J�&�!+�+&�x�FEt�<a���g��E��Ώ��פ��<qA�^4�?�*O��a�GI�4�'��S�1��]�U΁�Ab���� V�T)��TM���I��ҧD��w��ջV�H�rB���������7��qb:���p4��1OQ��C�.4ep����t�f�~���_$�r�z�-=\�~��'k;�(OX�Á�'�v6��V�0TN ��a҂<X�i�w�Փ-�\���?��o0��A�̂���ႰN�d�P���;��gU����-ٲkeXԲ�.�8��q̓UǤD�6�ip��'���9Bp��	؟��	�'�`	SC&gj|I��ۻ5�8p���X�e���߉H���r-�
���@��f�����ě9�DĐ�� _�5�g�H#V)B�(AI�ݑ&�ާR<)8e◤6Ƙ�>��[%I$$���$�<˄�7"ٰO�E�D�O��d;?�Sd��?� �\z��B�h����˓' P<�?O6�#�O:XJ��L4��͊�ʒ�4��I��HO��O�5e㕋"�:c��=��m��O>��܋'.�\����O����O��XH���'��zD��1oCRU��B%P�jdP��� w,��u�Y
1��BG�J�����D�2/D�;2�P�hԂ@��ʉ8"�H��R�����A�Fυ-j�VB!ݟў��0�[W\Q��Z�b!�6/۟DyU��۟ܨ�4hӛ���$�O��I#8����0~tX���ѫfA>���d��2&�V�k�j��4���>�t��I�g��IhyrE�s��םx�F�'���FYܰ�d�ӄ;���ȟ��	��\�Uɐ����|R��߮l����T�ټ+���0̑�YV\���A}��\��z��i��F�8i#¢<	�@K�v��O)R1�H*��	!�f�j$n�q\�#a¹[]V��OZ4r���<)���ܟl�IJ{ݢ�"�`��H�L1X|$����ܟ�?�Obؤb���1|���
f�� *!���'W���n �|(heπwT�:�'
�7��O|˓-� �пi���'t�Ӹ�0��Tf_.}6�H�o�`;ʼ� ������ٟ8��b�x�
����j�����N����`�׾s���I�,�V�I�CC�>�pEybe ˦����*8V)ѳ�~�0�1D�F�*%��	C�D�X�yD#�&>L�-���[�!�"�'��O�"��
U��is1��E�0qc�6����s� {��d�(9#IN3-����g�#�Od�&�Z�d��>��)r'��yI\ɓ�'������1UmSg)�Yb��G��8ZB�	iؤ��&ĶD�\ r�#��@I^B䉫 b��K�O'#0R�Y���	z�B䉟E�t�	�5s�~9Kbɯ]�B�I�W-��BP�ќ^?N])�"��m2�B��>c�D�C��ݡ2*����P���B䉕t*�@/K�^���F���&C�I(a����=��F'`!V%D�p�$$�q~�AB�7��ڔM7D�$�$��Q�8��gF�"�`{�H5D�P���Z�>� ���#)@���Wa%D��S���w��k�� .b͸ThGD#D��6�ؿKX����J�n&H��;D����A��qԦ(2E�$a ��%�9D�Xpdꓜ��L�Ŧ �mr4f;D��d ��T�^�� ��:��qN9D��W�\�b��m(�-O6/(���R�;D�`�5�U�F�d52S�G.�r�R�4D����)
�z���F̆1��yd/D�|z�*S�P�c��/Y+��Ci(D�(��uz�	�5Y�q��ٛgd,D�d��ɟ&6����{�
6a8D�����ua8���l�W��`���y��7!�nQ8C�fl���J�1�y`�.������T�.<� )�ʸ�y�A�=2/֭�vA� Y8��wII��y«I@�}Z��	l.�7�\��y"l�%(�y�A�����T��y2D%Rܥ���i$�������y"@ӏ^��뒛	��f+�y¢�4(�x$ڳcK�u��(��
W��y�eѸ��[�+U+n*:� ���yOٖ���1�M�p��SPa��y2gÚC?����I��g�B@s,�/�y�O�*����L[�D��cE*�yR+�+$�U��
��\��h�-J��yoZ�Cflͱ���*e� �����y�n<9ɜD WiC>���m4�y���iT�(�'��2%�K���y����4���G,���q�,��y��{�@�Kp-�W�<�"6c��y2�A�AXA�cY
Z�q&�p<a��,IE�.B��'9p�Y��Пd1� ���,\8*�y�A�]�`tBs��xAO�C{>u�	�q2�m�l���$2|cdY�`�*d�"髎���c�? x� oA�d�	֍�{��Z�@����@P�J\X��ZV+��wX� X�׳t`���%5"�z��O���k 8���% Ơ�u$l�f �'4("e�I�5��P)�.PK-���'�) �5��L�f�[ �*�*Q�LB�nX���ڔ-&�$2�ӫm޴a��'?	�����Hě'��P�K��)'H���H���KaX�D���i?VcZ�Z��N߂wl!�@�θe=�u�u��0ҁQ����ēkh:]���y�Đ�l�F����'r�#��epPAs]G�O���x���*c�H K��S�PЂ��S�ᲆQ���>Y�Ƅ�d?�+�*�|e2��!�L9K�k��P��#��St��E��h����'����D�/�b���Ǝ�vj(��
�'���ՏZx�Z=�m�H�2�*�c�-u����ē^[���d(ҫF5&�ч*?���tD�zE��V)�2Ʈ�Xs��:�0<)&�1��s�׺3��6M�.:���C�E���q!��>+e(��@h�>d2��y^�pJs��<y���ē4��2U�Ǔ��I !mMUXD\�'����J˸n"����NH[&J�z�'�����]`3dîI����慣OXP ٱ��2K&̆�	�1�:TbdJ�>a�	f��=.���Zw�Sv���.m���6�+�Ӱ ����'��e�1�)!gAM�O�@�	�'���LU����G�n[P�TG��S!�%���n��L�E�$�8�I�G s ��p2B��#N�����#h0�ѕ��<1Z��"ڴ�-�F�X�J�*�sU�͑�-���+4�4��)4�A��ljz-��
�J ��'X��X � ��R'*�&p��5��'Zय़Pݳ��C�r.�����:�ء�"OVA�cܑ*�����L�-)ļ�m&y���6Jɞ{|�D�	}Y1�εٖJ�)�~��_��Adٮs�j]�$���x���
$���=VQ��炅А�bǫA �L��ih�.Y�Y
6<F}�GږeԄd���
>Z�����K��0<�",��
���8@�@�:6Mʶ%À��!V�2�>��ň��
�L��6Ȭ�b4*��3�O|@h�ķd���I�!�FM󐝟8���\�B���)�/H���h��5,ň)���/Z��t��D�P���3+�!�d�:I	��sD��9�Z@��I�^<6�����?��|��<��V��|І�；á���b'�Ƥ10�X����t<�ǩ�>7  51+ߏ�4�G��RS����48z$��e�2X� Ah2jFަq��g≽ J&��	32��Do�)C2���O/ H��5�:^I��N0e�l)�� ��a*4�Чx���Ȇ�{��0���c|�cA/<O���$HW"����"�H�2�8�C���H�IޱP��p0�,ՇP�hD�4P��	�t_�떀a4j�%`R�*'=���>/"���ߋ���&TА��.�����*i�>���֫�y��]z����	Լ��F�&}~�P��5s6Jʳ �S<��J�#�XP�q&�-�������M��y��)�l��i�J/jE<�Ê�S��m�#V��,�x�)@�7z�@�D�x��݃,��+ԃO5b����H�*�MC�[���tcY�<�6��s�����Ӵ�	
	������'�)����h��88��ԹU���O��rvl	�3+�X
�FE��ܚEG=G�������4%Տ7�2c�&;�Aؤ&�
�y��O�?c|�@� �w��$�2-̹y|��5�O�kT
Qxc�C	���_Y�Ɍ�d�&�;37�� H�mNq@��\�yp�OF#��;N�(i�%8,�@ ��H�6ઘ����x����$r[��j��	
K�h���"*t"��)G�L������uax��.�JD�h̶H�L��5z&H$�������Ő^l��dS���yeI�+����f�L��	�5d��yר�<��гT�D�"���9��4��ǻz��µ�)\o�uN�*v��u���A�ߟ	���X���T?d��Ҋ�O����aK�U�Z�B�K��h-x�E�I�G�^u)d�J�C��jKL�c)ޥy��M�"�*�; ���&qD�y�T�I^t+`�Z�9��,�H~� �$Q벭��	�x9R�i1c@��L�&�j8�8	6M\"|n�Ȗ3P�����D$$�@�U�O�q��9��A馝���H�S
��?�r̩��	5.`��mZ,$x"<�㉛S�T��eK�	q��Qʦ���«2i�]��hܼ���8Ç@�?.�Drփ1s~5س�?�y7,@u~�[��H/-�0�s�B �y¥�.��d�v
Ã =�!#̎�`�ZA�F�Z�.'0=
��OE��O,Y����a-�5��]�i��m�a"O��Г��b8��f�R .|
}x'�i�R�E�2Z�Tč_Ax�L�F@B�l�=�pL[��4!B�"lO��e�Ǵf��\�f��$yՎ�!%捤n�ؙi�?ͦ��&Sɫrܓ_X�x����a��ؕ'V8U��7;,O�pZbkG�aT���#t\���W�`9<m`4 ��l0`��d��+����$��M�A�	�-F��Z=~`��b$�����H�,�<��`�C�����_�hQ�db$�� ��'柃i�)4��,��P�?O�8��)ѽ����5}��#�	�q}����c[�-p���K�;�, �]�:����o]?p;���牠/���i�n��i��q��&	�F!ݼo���d̒M�Q!c�ӾT貕zUF�X����V�`�,��i̅EjB�+cl� mi2Q��jI-4_�z2@K�Զ�XVݷq����nI3|d��"��o���x�+�v�'��,k�ǐҤQ�}��B
4;`P��]O�E�GU�;��1B�o�����J�Td�~&���7NS9R���x4M��0�r����çփ)��t&�"}Ґ��&.��(�G��j��8�C�șgY�l�6c�2}��H��#��~��y��Jf6ɬP{���O@�7c2���I���
�n\�u��ejA H��}�bA�C�����J� &��M�(j،���R#r(�+J�\��OtD+�A�&�ԱÉ-§A֔�Aת�VBT��%�ܿ>0�e���8M���0,m�	��n�>G��o�i�`p��]aW�S��Mc��
A�`�{`��R� �I�KJ Fɐ�P ��G�R ���Q$� �.���y7�	?$$�vB�l����ƴ��$ٖ;��X`���O��0%
��^���s���m}М�6�ߤ}�O����s=�p��.39[��;����ϮYt��`�D�rqB!R���0{�џ0�A*�5Sq���@Y/C��cV��x�RtO�h"p���_��t)��wd�"
�Az^`���L<����<�FUz���K�J6��#fAn~�Ň
��M%Oܢ�ЩHĉP�?7M��M���7J2�!���չA
W�_m@�r��IzDV<Dy_)͘	��ŭC̀���K�:d�� Մ���\�8�h�h)�	���Qv���č�"1����_�̐z�����;�ގ.3R��7�n�Id�Λ#����6�əs>��X� �p�� ��Y��tʘ��?IW��h��Q��!�	���t�0}�!���y���]�4��a2|�׆L3t�ܥ�2B�
��=�Cl��C���c�M7i����(9EऋWcԲ8��k�So�5�WN�8�Vɷ�ߚr�,U���O��jX�M|֕Af��LB��4Zl��9��)���=���O�Q�A!`�T<:RG�-#:����h��CO�H�`���XIQ��'X��E��[�����'> �Ī���B!��Ǭ��N~�'���Y�hĽ0�L��j��xN|k%f�AV�	w�,��ɵ���O�.�@��-|���̻5�V����M0�FH�f��3o"}Z�l��O���C7d�&,n�!u.Å�hO�-�1n�����N*s�F��U�9��`n���dսXm����b.~���_7B�.}!�@�f���()S.؁�.�G��V���`���vm��=	v�όK.��ӧ�$5<<Yj#�M58,U�KϳJ�Q�e�%n1�R��R5a:�Y%d��6}��c�#q�<uQ"[?�����\�֘�j���O�Sx�=j2�s10���O�=y�lbfrA��S�z@��a��<a�V��C��P�<,��e.�~�,uk4)[*lL�6��T�Dtm�ec`@	��b
�Cu	�'�r�`bK��zώ0 ș�:A'.b>Ę���!���O.X�l��<�'�t��$�3[J��b���k�JǬ �"�!]�m�� ��`��/ў�n���s@�°Q-����$Q X��<�:,[�"����5H�%�(P�p!$�K�F�;�BP�A�e�=	/L(I~�)���#F6Ucl� 
��-�h@�!S��|=��Fz"��s�JU�� 6$y�����S�^ZlPz�œ2I �)׾��<I$�&�2�=��{�@�A�fD:6KV I�>��'�����lw�TiRE+=qV��f��7�Bb�i�x�#%'�(:Ԝarq�[�L �Р������S宅�'��m�F2�5! G�>}�����=[j���l=�˓�~"/z���T͒4TD]F \40�RУ��_]<hQIŧ$��dA'�i�يH���;�	Ǒk3f}0PB%�ɕY3>*��F� ���x>��u�A��%R"EM-L���2� R�r�0���E�����	�=���������'c�1���$�ҲWr
�c#��K�4j!ŏ
b,,y!��ߟX���V�쉲��ӰSz�#���N5�O�� crd�
aU���5O������O���c�/��D�!�4$̎-Q%�	�"��@a�C�_E������%T�*6!6��л�Lخ)E�\�@MA�����3�D��j�-p��c�)|j�`:�FT�	.V�B�
�<y/O�i�>{(N�Q�w����{v���o��+�q��A �8��O
x���� �|�џ���ԋ2Ո�*פBC�* �>lO�Ujf���0�A���~f�$�ЭS�6Ě�I���23t���_ ��?!PN�+�*�#CKO9G٘#��^i�� �~�)A�� a֊TzC�����O�c�$	�V���	&�Bd��'yn���)��xX;��N�=��'#�tS�Jv��!�P�1����
�'���C��xֈ�
 N� /4m@
�'H��qH��K��� `!T�Z����'V����Euh%�G��Q�Hy	�'J������%�.�w%Mq�	�'K����#���\���3B���	�'i h#Ԏ^6vx��v�;#����'�����!A]�(ɑckş�Nh�	��� ��If�ǘ���x�( 0F�!�"O@%2mX�?����7��;M�ұ"O��c��F�$�!��	�K@C�"O��j�ʓ$�^��s\�J#>ъ�"Oz���J�M��ʇ�}	�\��"O�5�%[�䀛��Ŭr(��#�"O��df��[�pc�i��m%^h�r"OHqq�'�;`0,%����#*�е"O�@��.|�T���/ux���"O~D���N�Z�1P� B����"O��a5g^��JLr��)�>u3P"Onm蓩?=��D�U� ���"O��Q��t��1��8�(�"O��'	K�n�=��I�$Y�z�Hf"O�QJA�V'Q��@�H�� T�"O�4��N�
I&��{ ��W��	��"O�0؁�����E�;z����"O(�������KAԚ�("O��֨X��Z��1@��2�b=��"O�q1`&�0D&p�g�*���t"O�tr�e� L��8��%�d�a�"O0��G�ػeBϦ:Ք}i�"O�Pq@�g� a$��d���0�*O�m���"8]�q2���P�-��'��@
�3I�;� ד6��!Q�'�|����D�?:pd�c�λ O0��'q�����T�`�3�G;tgT�x�'�*�3d�2_��Z'"Us3P��'q�	0	0%�mX�#шn[��	�'�t�i�����7���4��'X��QE�X�%� }{��	���-�'�p���V�,ܾ���뇂~}��
�'�D�@�L8��0{��{x2�I
�'�*�p��ۚT��b�U�y<mZ	�'�N��m�%¦�ZFOG�D��P	�'�+3��T8�����%zU �x�'�d���j[�9C@���3p�N�k�'����.7{jt�"��k��u��'�\�%�-����bD�I��'���Ơ��ڕ�0�۪
)*�K�'�2���N�&�E!� �� )B8X�'xid��(yL@�y���I
�'�hI�A'��g�8p0WEV�y6xa�	�'#D�xGF��h�d��(M&;IM

�'�|��l�?�z�B��ӄ4�T���' �Xh3��e�ԕ�5	p���	�'3�%ɑ���p�x��ʧ�� �'�����$�}Ij��O*~�،��'�B��S�%]�B���GB�3�'�	�rC�1\�u��F��T����'C�I�UT�&[�|�6���Aht1�'i�]� ��\Z�`2���?���	�'�La�H(G<@�WJ�6q<���' ����'ըRT)�!��2М3�'|��c�^��� E�]����
�'�]�QJ�W:��1㞴Z�D�	�'��qc#�~j����X���y	�'�T��e�_ B�L�f%ϰZn` ��'ل�wȌU�a���� Q�����'�`Hg/X�Ag�E��i��;�$�j�'��0{F�U_����"а1�����'�QI2��#4�C5(��H�'|,�
�$2�zJ,-Y�e(�'���(ˬ'�:�h���"q2��� �iy#ċ*_�԰9$�^�L�Z�"O,�"�Z�9x��(�¥�ސr�"O>!0��
 )�\H�SeK;4м���"O��a�%ŃD��@3#�@°��b�|r�)��
z��]
�Ӛf6���mn� C�,(� �U̗�`,�J�=v��B�	��԰5�@-DX�U1ceTIv�C�IA���J��(�D�"��(ۆC�	f�������%�ҩ���<�<B䉦n�`����ȥ���$���y�C䉦N����M@�6w�}����/E�tC����(c��!����N׍�`C�	�,�D�SAF�O����϶CޒC��'7n���p�ϰ R~�8R���:C�	�*�АaeH�;ub���	�25!4C�I#d���%-!N��|!t�G2A���)?���*	s�l�f���)��G�Y�<��R�)�����$L���#� k�<�e�G�9=ܤ"����A�hp����d�<Qť��Pp��(T%H@�r�F]�<�h��}�4-+2N�:B�t`$M�W�<�Q��u� �M_�5�����U�<a���E��(S��.`[�4	��O�<���;�ĝ�T!ث"
؁�A�t�<�2�ɽi�Zu��)@���P�E%	n�<)B�2O�����NdX%S�dm�<Qr�F6E*��'C��:湲 �b�<q�D\�s���� GUE��b�[�<��n]8N�B����!�yI�V�<qoBB]Sծ;O�,$y k�V�<�!.J�w5`\���P����X!�P�<�v��:{�X���Q
rR��9���A�<���)h��2����5 ��@�<���5#����6V�$컕��E�<��*xBY$	Y:
jd	�b���<Q	��OC.��"S;|�h�n�8SH��'ɢMx�:5��$�
kͤ �ȓp����ʐ;.���pH��7ٺ=���̉�)Q2��
����a�ȓǶ��Z�:V�Q�$O؄""0I�ȓO�t|`c����R�IЄ\i��ȓ7��eq����(aF�rVcǕ^-���ȓ2��p�hM3 9ĕ��I�k��l��8�Z8���L_`��Qf'�T�t�ȓZZ���0g9��r�R.=hqO�x�`�{Dx�j7��M	r=cE"OH�(�ѕh8-�E���q"O|�r�[�����%x,+p"O:t�P�8�0ە	Q:\@���6"O~�����/\� �NE��e"O�8"�K�qF��a]���Lٖ"OF�z�O�]��@ªkCP"O(��]KԌ0�Rl޾=��0"O�I��l�@�Fe����|��9'"O� z��tE*��J�X ���$"O�PId!��(���z����,�"O�<A���nr�1*U	9�F02"O"Px�OҙR~�,��h�!U����"OjT�0b��4�dЅ�x��`�"Ol����EN���2D.�*�x�Q"O�@���=	%�|X�-�T�D��"O�H a��_&jp��늅��`�2"OJsF�@�:���h i�> ~DP�#"O�9pJ\
eNXX�H�T��4"O� ��:v�9f��Ac�B�=����"O�$�V��Hx�5�'/:y�V"OJ�q�J=�0��b���*����"OrE�0NR/�R ��� ��a��"O�d���
��� K�!��,j�"Oމ�`iϲ}����/K��"O�	�FHY�3�h
��bw �@�"OV�G�T��=� 5�Á�#���ȓH�"̀4��P%�� ���m;�ن�sf�����&\X�#J�`�`�ȓ;X��S���ww�y��.�`�$�F{���fɞy�v�)p,�5���.�yB�~2�0)�-0��H��	��y���\��=B��!5���w���y�%��/&2E��"9�LT=�y���(7�� ��.��>�K����y']�q���2Ղp.�����y��3�@����D�^�DԚ��y� 
 ����Sn�2U��������ybAڤ|}�Ɂ5҃=%N��I�
�ē�p>��Q=+�@�j�'��VI�
��C�<�� E�2M��6R7hT�,��( |�<YV��4sI�d�W@�1 �}#���v�<��o�fa@d��p� `��m�<�&��g�X[el�4��ջ�m�r�<1�kXx��2�蜻��x�ckW�<Qr��7	C���r[`$�c�]�<Q��]�v��b�B�<Č
�g_P��hO�m�Z&b=Pw���b��'�0�ȓ��8�!LB)Y�d��NP%�ȓc��� #i�g��X@
ǻ�hĆȓg��mJ֤ضK~��H�A�S| ��ȓr��ж��Z��x`D�=s�D��ȓu�8�أ�^���U��E?�a��c3����x:��¢��
(��q<�U����EA���+�>QQ��D��Ĕ'˨TT��9X�HI�'�>$���R�'�~h���,{ȅ8�Đ�n��
�'{4���!ɰ��t��k�f����'�� f�& 'X���N�GTZE;�'Hq_�\�BV�
��A�	�'k"y)G��a&F\;g�H�0n��	�'�Yۓ�9w>|���PgvQi듋�ɷ~?8��"I�	T�e[R�؏+�C�
"��&�?x���+����G{J?u�aD���Xuc�I�x�U�(D��Q�M؜;�L0� O�kגQb�4D��pc��(��9Bs♞߆�Ѵ)3D�̈��N�K,��lK&`0�B��>�
��`�T1P��#oݢh�� ^$u��D�ȓ)��͢S��-J��I���h����Y����p�`Q�mL�d�Ȇȓta�@83
@.'?t��M�4��(�ȓ^�=B`�W:ք��OZ�f��YbU�q�JHdx*b�
�Rх�I�d�P!Cc�R��T/+�
����|@3�C� 9x���j ��܅�~A~��ch�"_/��-°!9B=�ȓx��[�$j���� ˞|B�CA�<ag[�"�H�@R�u�R��@�<�sł�q�p�2�L�7L���#��T�<�B��>-��X%�]>+��i�Ӭ�T�<wG�>��iXrIT�7lk��@F�<	����dR����բX� ݂e�<� ���1�\�L��i�&�8R���9E"O�x¥�>8���	b&�z@<0Y�"O"��Z)0T�]�G�VB$!�"OZY	 �=Ͷ���K�:�`2"O8ĻC	�P�����$�)N�4P"O�|�#h@ ߴ����m�(S�"Oh0�׈E�d�ĉ0�_3�H�u"Op$۴�
#t�1��.f�"���"O6UaE��l�Ppaݤ5�a�"O(�"���x��	��X�b5�q"O���ӇYwQ��hZV�H4�"O��:�2B���F/.���ia"Ol�7D�1Q����D!uR
L�U"O���a.>q ���Cd0�p�2�"Or�ô�%xzj���͏.���T"O��{���>�&m��_7WB��S"OB݃ ��&U�Ұ���zԬ8��"O�`�%_"A.z@!p�I*{�ȥR�"OrS���3B�n)`�%C
�@��"O���B(ء|$�l+Q� ~�D��F"OBU˰)�%`�qVc�-�T;"OQ�e�e�x�DbU��|h��"OZ��T�,E�>����
4~��"O������yDyK��C�xx �B"O��Dʬ? ك���C�|�d"O��*��HOz�*L�+���#r"O�h'X�X6*䡕�2G��)@�"O��veT�D�0��V�{�����"OX0yt���T���K�7�����"Od��t#ءoĕ:`��=u�@p�*O�������!���<{
�'�`Y!�,�>~8DÀk c�x�y�&������Nֆ>`U��B�7�y��\���Ѥ;	Hb!k���,�y��.0����	�D��U���y2��F����I�!s�Ь"���3�y��Skz���c��BL����C
�y�� H$.�+�eֽ5Ԭm�����y�셦��pơ"�̩�7����y"$`B����j�Q0_~怆�,�z�1T�F,���@���X��O�$3�)N$ q�}���1N���*ũ�� #Q���U,ʆ ����x%�`<df��ѧ̎z#9��k#��x!Ì�GP����R<'I�x��p$!h��<P&���돴o�z	��%Di�­��6Y2�O�6���ȓC��SaiA�lǂ4���_,R�,���4���P��Ċ{Ѱ�HӭI=|�V��j�&@��"]�08�X�O�9h��ȓA��h���Զ!��P��Z>��4Ī,��$B*EP�ǉ�M8T��ȓ`4���`b���9Pbbܐ3�\܆ȓ'�:Ի��)�p]iV+��3pن�{' aڰD-<(�@�3]�D��{����*X�L����4u��U�R�b��=�h��ēR=R��ȓ��8Ҥ�j�~���bJ�^�(�ȓ1���F�41��k�c�#f`!��#��8C�IE�8u�����ވK�<=��l�65�ԯԼLT8p��.N�"O2����>z�$] ���i�z��"Oyp��8yN6ɐƣϐ~���9W"Oԉ��.C8YB�O�V�9g"O� )*�a�R9:4��C�N�F,b�"O� 9f+��!�u�_����+�"O�pI7���SsGO��K�-��"O<a�`�־i����n p�̅�U"O �����p_��u-\[��au"O�����ӡZ0	�<J��0�$"O`ih�%	�Ng��:T, 0c��U)g"OfiY���X�!��M�.0�zu2"O�AH�E��W��"Ӥ|���"O8qR�٣n��)s��Ƿj�*�x�"O��b��I53R ��F��
�ԙ�"Oh�I�!z�ΐ�G�;�l���"O��0@��
SII03p:e�f���y�(�:VK�$��
�[���ݜ�y�ˍ�|�>���%R�A疥.���yb�T�(����|~�a��E>�!�d ���$Ņ�lX����'F�!��6H���1熀 mJ�4�O�U�!�d�*���k%eW64�6|��)�!� Z 󔆞�R4�2HL	G�!�dT>5�H$j7h�*[�\ �&��lJ!�Y*�
Tҷc�:Hj�f��$<Y!�X���RN]�uQZ`�RA!�d
ԕ��H�^Р�CV!��}����O^z���"��
�!�d@+tr=r�i\�g��U�$�1�!򤒂UE �#��Av$ez�D_�f�!�DZ6[��a�D���5b�(D1!�C�%<b���(C;+p�$��!�r.!�ɅKV���4�#�t�B@���&�!�Ć�;'Xcw�e��mr ��$k	!�[(hA�F'��X�Ș�B�t!�d�%YP����ܫ&̉��A��y!�dG�8xbN�4<	9_�L�!���R�j$I��ۇ8��qi&Ҙ.!�dI�d��ycM�/\����f��!��4y!�!A�F�����%h�!�N���|���n�n�6�H��!�^��¸��&M���QL K�!��m��z��"r�3�jC�b�!��d�>m�1��]��S���3t\!�D�, 1�(1��N"U��T��d�!G!�$�)IZ	��4z�v���(R�V'!��	� �4%����P��&B)�!�ظ�p@hW����m�!��x�!�SK��s�d�"A�����c�q�!�̞^p~����S4Tt�k0:O�!�䀼vX�y�(̳~�� dݡ-�!�DQ���
	�eQ� ��j�!��),E	�pf[(O�9��KX&l�!��B:������c���5$ӆ}r!�d�/��e�*@�	b����i��,n!��LJ��S���dg�ܘ�BU7�!�<y"�4�����+\t!�⋇qg!��@,��`(�۔9K�5���	:S!���&`�@r��P4""��I$=!�d �F<r�%�%t$�hWF M%!���cX McE��f}��k�,!�$��@�Z�ɡQ�E׶�:@ˉ�8�!��"�h�y%��O���z$�φ.!�DDe�0��r���
��ɝ�!�dDM�r'љ1�dI�%gLr!�d{����珟:�v��w���kq!�$\	^8Q�%���4ɦ5�!9a!�� ����	��$�q�˔z:��`"O����ɝQ��	�j���^���"Odx�bnDBmlU�5i׺;��hɓ"O��Ru�O�T�Z|�V�6{� ��"O e����c1U��8|�\�t"O�j���N�\T�0�ҜB����"O� ��kC(O+��ʁ�Ǘ3�HyC�"O�y��ĵ:�$d൥ڡ2����"O�1�"S-M��j�eJ&;���"O�� p ٗ� ����1�X�X�"O�y���m����_�E]*�q"O@p!�	�%48�t`�r��d"O���v�	*A�Ik$ ��Z��ɗ"O��r�رv���R��ݻ�r�*�"O�c��{AaL��2�A�"O��z�C��Y�8�G��2�L�YG"OL����N-��,�Ĉ 6Ș�9#"Ojh��OF[n�I҈�?i���"O@ �P,D�_.a���|n0��"OdL�ai�9 �6��4S�yI�5`�"OLM �/В9dc�P�@���"Oh�ᔯ��vpF�W�`ys"O�L�УX�?=R���A�<�Fh	@"Obe�a��Un~ �!�	�ye���e"O&�R�ؐ�j�k�g78<�s"O�8�CEX(L�<���&�
*XT��"O`3�@��M�͈�hZT��Q�"O���.�3,d�ŧ�*�8Q:5"Ot�Ѧ�:Zv��摢c�n!�u"O�����I�o1j����D"h���$"O�	y��9l�:�ÕE��fQ�s'"O�}@	�����$�=J֞xp�"O(EI f��{����	ss�4"O0��� �D����4�3�����"O�0bR.D�(���
�G�,o��aB"O`�h��;����
�Dc�QQ�"Of��"��I�2��FѴGb塑"OP�X�B?$QZ����O4(.�t��"OvQh���=�L��f�#;(���"OP(�b�n��<�bF��u �ڃ"O�	��䕃t���rBӾK P��E"O"1�D�ć�X�gÍ
Y�����"O����$�9yfIڑ�֥X��m�#"O|ɋ�6�n\�BR���@V"O��3�!�|7�1�W��,"�u�"O\�a��Z%t���Z�A�=[��-��"O�%�L��Mm�	0p \�8��$R�"O�L�ѫN�P�Q{'m��J����"Ot��%Fд8�k:A�P���"O0�Z!�85sh�#f*�gd(c"Oԑ��-u,M!�A3dH@��"O�}����n������ j� ��"O.ғ-��5�V�p 	�P�T�"O�{�ɗQ:�L��L�.�)��"O<1�DB�CJ(��X�d���"O>�J��U�� @e��ط0D��[J�^��FF
S��%!dl/�Ov�76�a���u�r<�w˘��C��?Z�,X���V�`NȢ�Ė�V��C�	�_O���ajF�'�(``��nR�C䉫X�2�0�o ���e��4)�B��W�@	N�	��QC��Q'0W�B�I�%���A��:5(p��FW�C�RM���ԉu���Q�b0B�)� ���e�½sל=�"n�'���ڧ"O����Y�A�F�R�,��P�� y7"O`�s�9*0������"Oh�)R*^��$���+|V�usP"O���#N˥]M������_>�$�"OҌx���q�8����Ҿe,�i�"O�����.���s'E�,�-�v"O�\�,���J�ǐU$�r�"O@0�g��~x�3�}�0$�"Oڡ��)ͣ.�Z���+�&X�.��"O��x�eѱK/��9�	��Iޮb"OXl��H�m�oU&Q�|xS`"OB�h��B��m�Pm
��``�"O^���
�2W l\�F,Y>�2�ba"Ol`D�<jȘ�(L	'Ia��!R�D'LO z鑲�pE��)�*(#�A�v"Ol0�$39�`�C+�;�pF"On�	�	K�~�E�jƭD�J8�"OJ�`��9�l��
&m���CG"O։�5�L�R�I�4����W"O@<�����y)1f����� "O�� ��|�D�2VD2t�|���	l�D��!�|��0�%��!�j�4�)D��{S�Éx�6I(�L�����g+D�H�%`�4M�|��ː�J�LDcՅ>D��Y����=��c��9o:�k�"D�|�T*ȈX�P�-������#D������L��Л���:�4�s�!D�ęs���\�vL�d��v*�X���O���G��'�LP+6^���Co���@)Z�'�`���C�l
�'�H����'� =�1�:P�4�:�`Mgh��	�'�t0�e(̐> �, ��SLbp��'���ك�wB*����B��t��'$��À��01����%���<Y !C�'d�к�ʩ]���LF
D�>К-O��D�O�˓��g~r��q�|�S�����B�>�!�dآI� �b�T��0��#����!��$I���E�I)?�E����A�!���GbF�H�OCD!�6+��_�!�d�G��L+$�]`���4hP��!�� "Gr���H�*z><s�邛�񄏀%����� ަ���y�FPG��˓���?����
2��[gV���y`BAY�}�!�׼���E�u��MònC�G�!� �(�+BR���m`F
�FxP�ȓ,Duy�h25`tW�t��]�ȓ0w�A	be g?�$ �aN� W����T�T�Pp�K�%Z�7O�;���)U�U�䉆)Lx@��+��(`�'�Є��~��GۥE���i�m�^K�B䉬~K\��d@��<��ण��yu�C䉻q����Ѐ�(v���Bf �:,o�C�I�D��Avmw��Y#�B0�C�%]�<ytcӛ/m�E��ѭ?T�C�	?y�jY���ނ(�����:�Ob�dZ�_�f�0Fa�((a���b��p!�	y��(��E0#F�fU0A��m��UWF�0�"O(5����~�ΨfHO�\��D"O�1��͈Q��Hg%�>[����"O,��2���R�ڬ�\���"O�\X��$rk�e��F�0.�&�"O>ѣ��U�����%]�.0xP�G�'X��=B��d�Wc~Lhp�ÏH�8��0?� L����E�yT��G�٫	;h�:�"O�(;S��0if���i�SQ:��"Opm��P41��3H7	MJ2�"O����)�"MR�Ź61p�X� �"OV0����E��X���ێi��=�"O���n�3=�l��e�.
��/�hO��D�O�"|ڔ�W{�����Q;�ژ"�^gy��'R��|r�	�n ���J��4A��f��6C�.����u���r�D�61
�B��[��erK�50�<�4�_6zh�B�ɻa�����)�A\�`�v��f-�B�I�a�Pz�B0��候8�HC�ɖ+�	��o��,��K��C�t�B���T��U�
�1��t�� �#/�C�	0[K�(����2Z(ab��v?@B�	���4��cS?m�f1����4F��C�	2ym4�%�**������:��C�c�0%h��ΆG� 4�u��0��C�	�Ze�a)�f�(&�yD�F!�lC�	���A)Э�1�����5�8�=��"�?U �@\n�21P���n�.�1N6D����e)S�Z����Z�,���g�)D��[p씬K��q�D-��q���z��&D�8���B��3����+Dy! )?D��C�تe@�\"u-�$z���E;D��8�ǦK�qX��[�)$��"��8D�X����=6����b��)2�A�h#ړ�0|z1&+I����@l�-�����/l�<��&z��Qڴ �ٸ���@�<��oףa�.%	"*ޯ8��H���<9�g
0I����4��,C�8H�UNS|�<IBI8�ʨ d ����C�U{�<�@C	VϺt�bN�!k(��Jz�<��ka6�*V� ���f�}�'���!��X�͸���#e�IٚB�ɵ_r�e�WN2/��[�m�aM,C�ɘ(������\�U09���ǫ�B�I0n,p�f�!-ᐓ���	��B�	�$L�dy�ɱ6����'�}'*B�	� `(�x���S���á��'t��B�	K���pJˏoݴ�E.T���B�I���Պ��\?�����L�@B�	�M�0!9����f3���J�C�,B�ɋeτH��/Xu��8֟.)B�	N�Py��Ņ����fR"�@B�����!(P"Z����c�c�B�ɰx����k՗;J�9t���W�JC�Ih/�x���ݸ*�]PV'�5yX��D:A�d]r��ļ��xP��,�T��ȓȰ<��#pڔ񑴠��Ňȓ$Ix�:dɀ!a0Kђ(vDD����ѩBAP�r'�1�`��jR��ȓ=ǌ����-/񀱋��r�:]�ȓ�X� b�ČD�~��G�K�f�DU�ȓo����AaD=RЎ�C���M)�$�ȓn�8��U�2Q���fG۶;��|�?����~������"�X�z ��G�<	�mA�n����᭕V_�̒�eUE�<i� +t����G1��2 B�<�UE�40��A`���&������<9�� �28�!��*Jb&�{�<��a��yI�X�N\_N�5Z!hQvx��Fx�J!^AĤ��(���N;�yN�#=T��s�=p����S��y
� L�9�j��3���ԭ�YZ��`�"O !lGi�� ۲�1R��J"O��5�V1;��B%O�$H��a�"Ob)ᧉY4��0Q�܊7)F��W"O<�`�B��z�PЗgE�VH�1"Oh����$lje�eGɒ�l1 "O���H�pJq�Ѕ
�/�DaW"OF�q��U�|� �À�i^H��"O
ذ�@2!�L#�a�//ZN���"O���SH�q��ͣJL���"O\ hWe�d���Ə��5�fqR"O�<Y�CS�X*����ϒ���yHu"O~�2���G8��D�Z�[�h�"On�v��s��-Ӷk͟$���RP"O�8Kᢄ�U�ؐ�t��h�Ā�"O~!�%�
�����)�3.VY23"Ot1X�bR�Uּqb�Ȝ�M���XG"O�e %Y,B��V�X�IN�`�u"OH��-�
��h`�E�5?j���"OT���A���0�6g�<>�J"O�i�%X/}���(恋JY��"OL�p��->(��U;1�R)�b"O$�ŨX��%Ι1��������y2�ɢ��sp���2�GG	�y⯎�@�$��ǁ�-���s�'�y����j9��ˆ�����c��yR�ðb�(B#/�D�D�Df���yBc��0�W��/�*�Y����yR���$C=�L�
Z2Xu���D)�y�A_�H��S�씅%�Z8IP-��y� Y~A
�EZ�- .u�m���y����]��#�R�P 	��'� �y�#O��Fd �W).����ED��y��Z�'�n5��� ����𣔃�yb�<y� �R�Q�5ڬ��F3�y�MM/԰a���!|�>����Y'�y�& �D��M�
z=�-E��yb�5?ʐ��Q8� �ud���y�D	{��1�ag��AA��g�L�yc[���t)�aʗ4�I��%O��y� � V�īW,�B�W���y�F&�*�
2K�28���&�/�y��G�7XD�����_�mseE4�y҇��O'�h���z`�8@��
�y�O�l�����H��j⩚��y�Ko~py�"�]e��s�J���y!�0����gAـ��xp`����yrA�6|������̫Xt�nF7�yR�݅&5���VHr�,��woӊ�yrɜj�"�ipB��9`���Ƌʹ�y�.OZ>3�O�04i�v�Z0�yBl��
����E��/�z"vJ��y"��z8��E��v�>�S4���y"*R�m"�pHg��n|�Z��1�y$�42��)8uƔb��5�WmG��y�ᐯP�� ���%e�H�����y�[�L�1=M;Z!�GM�8�y�`[�l����+	1��\0�@�y�DC��Ρ�,I8^��*��0�y��Ҹ���c$�3jG^dVG���y��@
#�~aJd�K��rl+�[��y� �>5 >��҆�٠��	��y�(қG��(�$
����H��S��y����mY��( �	]��3F.�y
� ��Qg��#�̅AKG3W��@"O4�+'�B?Q&8�[���6J�)""O^�@EB#h���2ɘ�G �Ȩ"O�\���W�~�����Hɼ}�@���"O���FU�I'F,�dbO+�D�h�"O6�����1J|�
�W�jˢP{&"OB�*��P�X�����<�m�u"O��Q��:,ȕ����^.��2�"O�-HF�)�I����$0<C"O4a23T=T&�Փ4h�Y!
q"O2���o�6�l١ǌ$zD��"O
�;�*M�Pg`��7��dI�"OLɒ@��QȾ�#��͋x�n�R�"O��e���6�q5ȐH�hs"OD0�o[a�\���A�bl�"Ofݣa��\�HܢL���	�"Oj�C1��0:��Q�	v���#4"O Q�:ˈ�3�ӊ2Q�`�"OF�1]����2 W�mBz�a�"Ov	�qɂ;1Jr��#�� '���"O��اo��Y��A�i��K"O��#s�=lXZ��"�]�w���A"OBY���E�v<�C�G����q"O4�"��[jY����λ|4�	p"OF%�%L^�S�}�@��h,��"Oh0Ԩ4Md�G�W�[e�t��"O&�j�)�������z6j@"O�k4*�6{�,�K��5T7���"O�e�S�O�Z���&�r&\=��"O��i��6] �!�q��0�Q"Oyڰ� F5�$��f�+���"O!ї�ߺi�j��c�B�aM��c7"O�� УR�TĭQ�Ѵa9�-p$"O�|�e�<Cf���pcEI0��3�"O��f˒�tQI �D
w���T*O!���N�\XT)xӏE��KTu�<��	-��02�� F !kJt�<���ݞod�P�pM]� ���Z�G�o�<���0`Tf�`�ر&&n�*�e�<��	's�@�� _/hۤ�B��b�<i��g0��;��]vW�1*��c�<I�.� 
�k7�[yd�p�ed�I�<�A��uq��;@h�=��=J�)E�<�b�̆K�J�P6�0���j?D��C����;c�l����ntY>D�а�R�r���I�جy,�b6�:D�(�#�ܐ,�6���U�d�ajv�7D�����;`����lU+T�>�I'I5D���d.7�HK aP3C��H��'.D�4(�앴S$�9����-�Π�!M-D��h#�G���҇g�	�����J6D�96hԖ`�1c�&w�vM�&h3D�,�/��z}t����n!j��D6D�P�vLӮ-������V�;o<�b2�7D�d��P&���1B���f7D�0�� G�{��|���ϝu��0V�5D�t�6	�}��J�N#rNt-��K2D�|0�)تn޶:gh:.�0��C3D�x!QiH�,�T@����&Z����`&D���.��}����]� @� D�������X��.{�2��6 D�H�u�ר[zݳE.��p�i:�f3D����n�3I�� $|4l��U %D�(`��̟c�N,�� Cnf03�G#D�� �a��K/$�>+E��&k4ݰ�*O�c ��.lo����E��r�L�I	�'DlU{f�X����6"�����'XX���4=$\a��:*�1R�'��ZqK�`�x����f�JLX	�'g$�0���:l� ����Z[~���'O��jV�>h<#f�ݤvf�h�'o��a��bsXx�D��$���'�p�0̚�zSЙ'��{����'������	n<�Y�ٵu�պ
�'d�����OBB����tp���
�'ҺT�� E3%伨���s@�p
�'�<�	��6~��l����3�Z�K
�'�x�* !�)^���G�W4�$�	�'�����፯<��3$鏊fB�(z
�'��$gòB���i&��<�tHP�'-�M����5����*�B��H�'�}�`lQ�<�е[ ˎs����'���:DW�y�H]JA/ݪ�
���'Ⱦ!Ȑj�V��X�lJuZ
�0�'����E�ܫ+���7M֠A��%��'��% b\'q 
Ls��S8;�X�s�'Hh����w32H��>)\��	�'���Ȑ�$:ژ��Q�݊�'D��R㉿]��	s(�	L<H��2�*���A<\�`��Ó�i�؈�ȓ@<��V
�
MŘ��b� �^��ȓ2��`�� �]H�R�/�ג���Wn�&e�����椌�K_���ȓ8?���œ��M��n�êu�ȓj��� !���x��Hµ+��-���{��M�e�0^s�0��b9*:i��0�
 」�f4�uˢ^6p�ф�r�9r�6Ko��R`��0W��}��C����
�|���!qm�/4����lV����@�2��D`�\��1�ȓ���gܙ%�h�����B����x�*�4K�D���Y��Z�� �ȓS�-���b���	�n�� �hd�ȓ4�zr�K!)���	ѿ[�A�ȓoH�!�'ݖa+�b6�9�<�ȓn��3�n�3�n�B� Bl��PG
)zq��aA��c�T�"��ȓ#�.=1E`��Xt��3�	�P����+�����(t�
Cc/$08H��,�@Z��ߒ-޺�����-	�ф�Dlj�#S�l���$R��Ʉȓ��YA���kv1�e�)WĒ�ȓQ3��@� K���[��^*/��I��`#��$��ZD���A.�0y��W;,T3�Y�MB!�t�I�;܄��5?�(KS.�0�����%u��H��H@X)�F�6|����ϻQG2T��,�^(���=��
,�2���聘0��N�p�H��O�E�����X� � p��>n��`�v<>̄�m��Y� ��h���&�B`�ȓ *~�C��U�(m��y�Ɇȓ� ,f��?W�4H���k.6U��i8�dK�Q N�v�c� �r���ȓk�hB�/�f]��˒�O�Pf��ȓU^���UI�05Ξ�iA�fS�x�ȓ5m0�H��Q4�֞��Q�QE�<I��4>��hȁCH,kT 6���<� ������`	R���Y$��"O 0�T�*A/ ��`�,���� "Od�@W��[�l��GDZzdڦ"O(���� 3'���*��Z�s!"O,M�D!�l�A��]��6��q"Opc�L�@�*�rS���|�\KU"O�T�� X	(��(�"J1��}��"O.�R���Gv�ѓK�)�Ό�1"O��H�O�!b�m �Jߪ�J���"O¥ӥ�]�;�LX+S	סN�Y��"Oi�0�#\M.4r��ȓ`��� "O ,��a�;{�čZ3�ǦqWJԹ�"O��E蚮PMf��P8E
��"O6���NމU�����4*O�@�"Oܐ��<,H���3"��nK4��"Oέ��b�??Ť�r�U�N:�x��"O�ѡ,U�SҼ�c���=tdr�"O(��R W	ZF,9.!����%��y�FD�w�B���g�ld1������y�K�:N���P�g��xSm�8�yb`I�Wy6	J$fԸ� �Ք�y"EP�-j�`�hM�D�Z8�1���y2�A!��+sW�C���A�E��y�k�rX�PS�ű:���K��y
?�@pb� &־]ʇ��"�y��Gv�I�sM�0A�UB�����y���)b����4&���&a/�y���ցCd�ӡ+F��e��yR`R	n���X��������ٰ�y���04%bpC%��銅�֪�yRƐ�n�=j�Jۺ
��m,�y�6�<�RϜfe�m0�o��y��J�s
� ፀLr�A"��̄ȓ�QK��W�Je$�	�F^��P���D���ômH
3��R��<�`,�ȓ~[X f��.�&$+4A0Y�y�ȓ:�5QM�7G��$�e�L�n�jP��@��̉�I�S\l�@��7��ȇ���
�P,5eh��#a�F�^���F��� �Z�ʕZ4Ԇȓ	R�ç	R.qaA�!�E��ԄʓB�,��s/0l;T�K�@�tC�	�@Z*�:댭!ֈ(��ʻD�B�	O��I`�?� Xq���QW~B��}hXc*Fv����Z
h
B�I�F<�YcfOv���+`�V�	c�C䉦
���qL>�xX ��(px�C�	*Y��x�wl��|!@�(���WT�B�ɭ]YJ��#GNȠ�� ϳq�\B��;pT��
�B�%����a��j�C�	�[��mh#�H%�z4p��ΞD;B�	���ȷ��t��&̂a�>B�I
k8ν�|6�59B#�5���!f8drq���z[�������Rr��|�DUQ"�T�C����� >t=�ȓ(�~�	1�։"��œ�`�"4\���ȓ�d�3cט�3�#���%�ȓO8Fh�׈[�� Q��Q��Յ�R�D�s%ƂL��T���GH~\1��f���^�6�,!Q ���~Շ�0�f���	�Q��@h�� Ba�ȓ.&��dj��a�"4@��V�^��ȓg�0�����ܳ$�Y�6�m�ȓ,]��&@�d���ʶ�"-��S�? �D�Q,�<!�6T ��B�`�"�"O훆��1�<� %I����;�"Op��Tg	>Kp�R��O�Ty��D"O������(l삦��.D���"O����8#l<����
fӨM��"O�}�C�a��$��$A=3Ԏ5��'?�	���A�6}y���h�`y�'6�\H���.6��� /3`��H�'��tq�G�
p6�()S.E�VS`���'�08��䔉	�֭���D�J���y�'���8���(ШY�!H�w���'Zv�:��A�_!��3�(˧b: �	�'������"c^�a�DعW{�%K
�'��pD���5��P�SΔT�@p	�'� ��Sΐ�"�D��Jþu��H�	�'~���K@��Hz"��
l���z	�'!<]3��0@��� 㥌:g&��J
�'�,���JK�q*���Ȟ=[Sd��	�'��1'G�'r��u�e�xq�
�'��u#$�_�=^�Ce@Ǻ&�2��	�'�nx#P��kH
 (�G�E�iS	�'��L��ďl]j`��a�8�a{�'S4�D�)P�w͏{� �#�'נ�@�@Y�S��V����� �'"��Ǯ�2;�d]j���v8��+	�'���<ӂ Q���9Xp���'^N�ys�@7h��蕎є,�u�'����䠋+A�0ʔ�]�%���'�`�r��� ĬM`�/�
�j$�
�'���S��ڧY㬑��,F�m���
�'�z���J�"!>yq�LF�h���!	�'�*����ޓ8d&q r��rc �	�'��e'��x!65���;S`���'�i�����<���������'��h PGĿ.�0X#NA��{�'�NS�D�#88�2�nA*C��P�ȓ7�֝	R$	'\^0��������ȓD�8H�&h�.3�Ā��ޖ-㤸�ȓ7�\,�2Dצ0�>��U���z�ĆȓIZܕ1��BWZԵ���NE*��ȓGc������\���� z�:P�ȓyF(�:�g[�_(�|�g�3
<ą�}���!�NWn�<0�J�P�X��Ϡ(����UŔ�k�+,��M��nJ��a�U�9&���0NC
&.��ȓA�&�iDk90�	Ả�;䍆�B�6ʁ��8	Q#^�$�ȓd#j	R��m�~�i�Es�hi�ȓ}�p{��B(�x�s!��'�
���. D�@'��ı� .b���*{Z�0��$-�u)��D�'�j݅�m4&i�h߁Y�81�%�D�9�ȓ^sh��Q�R$j"6L��ȓ4@�J�)�   8�o�,Jfȅȓ~���K��ˍqİ�Q@_{�>1��$l0�Gg�#Y�m{�G�Zf�u��G��(kŀ	*����d�Wpv��(|n�z���I��!��o:6��Q��X���c��e�j�ي���[��I��--�vkF�Q(l���ȓ����C�"{E>d�V�L�,�(h�ȓ%K�U;��?)����]��ȓ7DQ�eߨ��u����� �Pq��	�ޤ� �*N`�{S
�#��S�? yC�.	 3�b����G}Y P"O��r(ߔm���h��\M���"O�����Z4P�"����m�a"O����7q6u:��U���u0!"O*ܱ�f,\@��Z��,��`"OD�8֊)s�Jc�c\U���"O���'Ɔ2V k�A�<���g"O,�z�!IVđ� ���1��"OQ���/>[n��T��LU��"O�̻��ȍ0����'j�>�E�F"O��3� ��"�����BݲQ��"O| ��L�Qt B�P���aW"O깛b� �z ��P!Ҫ��"O�M��R	n�)�i������"O�M��0�ԭ�d�������"O���W�l�L0��J�Kj�(B"O4�匊�/!l���fG5C��y��"O�D� ��� ��x��FަP�� "OV���/L��I���x�$��"OV��DH�)<����؜,F��"OR<�`�Ju�`0��G�+8�tjP"O����6��)�&_��F��"O�a���'ƴ�F�6Xꒁy3"O�!�ŏ�t�m
Zp�YH��;D��B ̇�9+�$+G�ŭC��� � :D�,�BK�<!���d�| s�d6D��K��ls��:�Eߺp�RL���5D��+��L�{�Б �C� A/x�H��1D�PR�]�1��Qp��F�4�CV�#D�,!`��v��ͣp,93��@zRN"D���GDn�t�cj@�k��s?D�\�dɒ�!�H�rl^<B�rAQ��7D�d���� ����-�!^k,�j�L7D�$�b�8%����n$q�ḅ�e3D�X[�h͋)&k��6� ����4D�hR�24��R��-*u�4Kg�4D��CkKE;x={��8.���">D�p�tj�sZ�� �aI<|Up���<D�t;�N����0B¢� �3��:D��WjL�e�L�C�:>�XA�+D��vG��@`�q#!	��X��.D��`W�A8x��u!�O�os�S!�.D��J���쁰 �ϴt���B�*D�� �kZ�~n����p�����H*D��A� W��]�i @J�m:6,D���q�1l4q�E�؍,��Yx�l�<1FH
�je[򢛶Q�t@��GAU�<I	E�bG:���&HJ���j�N�<	FD�WdAG#Dv��qG�K�<�t.�!	�V�Q��ĝ
$��W�@H�<i�f� o	�����g�֨YT�~�<I��{��pZ��R�p�^����S^�<��1j�&��1c���H ���;!��d���+��q0�i�ȓ|�`��4̍�B���΀X����I����fܑ& � ��5�b���h�V�1�B,Kd		6�9��A��f�b�"��s,m� o3"�n���H�(8!	�� Q����"�4j���vn�< ��B	Du0 s���*I+�A�ȓW�L�M��%�y�#�+B1�ȓ<�h���=Fp�{�D1�� �ȓn'8 3�b��[ari���cOl��-�R���`դ�v���L��zStP��S�? d���ǯ������m�t"O�$��E����٤�_�b�P\ؑ"O�iB��Q$	0!jW,�1���;�"O��0pFZ/T$*�
�J� t��b"O��y &�/�;�J�#_묍��"O&��6I�-˘�6�N�l����"O��I�'p�|�1�3oS�܂�"Ot#���"	zP�Qƈ��p<"p`"O���0�ɑx�%��	�1+�0�"O�z��n���⦠$��"O`�s���){B��B�S7f��#"Oh4�24:u���@b�,M��"O���A�tț��Ȩu��q"O" ���-;^�$!��G�MÎ!�"O����I�U��5b��$�B�ٰ"Ox��ծĐ�B��lPs��x�"O�����B��`D3�+�_d6��"O�Șڰ�I3"�ڑ=��B�"O��bl�-`�ҤN 7���l>D��a��g�zEJa�̠e�r=kd,D��jV�s6��#�O	�j��2	+D���#�	Eb���q5t�a��$D���� �T��Z���]cDhJ�h!D�\�)C5a�Pl�`��"z^��g�#D�ء����P�귍جB�@ݣGO"D� ��M�6,Ɖ�d�<r�ĝ�ba D�\Ҳ��p �鶌 �n��@�2D�8Rq���k���9e�f�j�`�$0D�<��BX2\UZMrf��@�%��9D�$��1RJ�i1��Q_��$h�6D�lـQ0w�D�(dI[<.�ĔIe�4D���_�8��W:��0�2D�H�X�j��}��%���c��+D�x"oS�%�@THRMN	g��	K��5D�$��V�b>��8�lX"q�V!�
3D�x�g�O<!������0�Ju��C&D�$@Ah�';��5)c-P+P�h�8�`$D��J�I�A6��VY)@N�X�O5D�`
�oP=
NJ���/��`mi*�C2D���g�(���@T���Up�-D����$H��Q���.d0��bņ*D����/.�u��)&8BF)D�\��!��}�4\�s��?($�
��(D����ϙ&/��mr0��U��R�H&D�H����P�@�Cv�̠T���Ţ8D�LڦkǄ
g@��EH�%`��I��5D� P2�Kg]�-��bF�;����>D���u܀`���t%"9b(QF=D� Y��\u�K��ǰ*��"�'D��`�b]�s�z�`���;nظ��G$D���a���P�Y �@�7������?D��Sdl%-D�{����p���C(D�D V��sh j����0�� :D��Ӯ@.���r�_1��*E6D�����7�2|+֋�VQ�u���7D�
"�U{T�A��"4����r�3D�T�QoP*9B��V���J"j��1D�D2�a�<�
`���a��A���3D��R!f�Z����G�y;:);��0D�l"����=��`�M3d,=��.D��:$K�Q�H�BL<$	@�8D� ���_Q�X�b�����2��6D�r�ƿ!�l��L���X��J4D��p"�
�p��k�i��\1ۆ*4D�� �+���8F��B�]�)�F���"O@]7�� ���[0�Ӎ~�`"OP��ŧ�,����es�9�%"O` �m�5>�zX�D�A�yzH�B"O�8�G-<!V���*"iZpJ�"O֨y��G Nb�S�@�lON�r@"O����ɉ�.\4����}6�EҢ"O���A΀�p��찗�&�v���"OȨX�n^��}�"�B�����!"O�<ˁe��w���D]t�U��"O�%�7�Ơ�X���ד}Y�|!�"O\`{F�U�5�*�7��|�0V"O�Bd/T)8R4��q�[�n���"O��E�X�\;������"O���E�b 0��%*���c�"O�Yy��_�to^�.����"D�l���҆C�����I)7��Dx�!D�{ǅ��X�J�q�@���b�@�H:D�P3UJɃsX�X��ΌOP���C<D��ZE�� �06N�5�R8��9D�����@���dسeB.0m����7D���+�q�L�&��n�FU*�/3D��k��Ҋ>g<tRU$ɓo%2IK��0D����h�7C~
Uz`�ѥHLX��v�.D��2�(:�(;bE�<,�UCd?D����xs���CO�G#���7D�L���D�cQ8i9�I�+�6�3�F6D� X�G�Ԙ[�惴8��S�2D���T��9���W�G���a�<D��p�^����/A�u"��1�<D��P�D�~��A�i�$�Tye8D��K��]�	�&u�FJ\kņ܃�"6D�p�� ]�@���3��x�l,1u�5D�`Uإ0o�=�venpP�Pf�0D���V��
 ,��焁+3��a�(D�V�%:��J�D 2 �À����y��R�43���?ʝҤG��y���I�hՠ�.�ʜ��3�y�B܇<�aEǃ ��gQ��yB/��N��y*�N&C[�Lȷi���y2��A�H����BQ=��$�y"�H
�~�j�	۷970������y/Hd�S��	1���J�IE'�y2MA�,�ԓ���=�����_"�yb�̕;sb r!Ș>��]x��ޢ�y@NIrZ@��lc��<x��/�y�.Vܠ��&T5
u��
�y�kG�ki<m"2$�%,�Ë�y�T������]�(�Z\C��О�y�g
�[��CbL�Ta��+���yb*�M�$̒� mv�@��y�����PZ���Y�֜x,R��y��[2IVء���ėMB�T`wŘ��y2��
�p`��kK?2q��a�&�y�0���ɚ�u"Zĺ�E��yjC#3�2@[��89誽�5Õ��y�EG�zzp���A0�f�HrLU�y�fΧmfq�'�5^��#��
�yᑳw�A�w�O^�l��d���yb�T</4v�b��9m�H\IWG¯�yr
�!M�]p��["&�E�����y⫙�'X��+���Lɓ��yr-]�e��c�#$��Vh�2�yR��xl�͹��9(M���FU+�y
� @d���/ �Cl�9�"O��P��Pf� (��R.N�Ĉ�"Ov WcHm�D@q��\4J�uʒ"O���FD���� �Eb|#G"O�͚G�ĽKT�6.
_.�u��"On�rD�@�
�X<�CJM$G,�͉�"Ov��EIě[(�9j��?�%"O��� 
q��(ע!��"O���2@Y#?�}�e�E+9Ț�"O8�t�ċW������?�ɺ�"OV\���?Oɸ����'>�I�"OTx�өU�n�tPsb�>kV�5�t"OŲ��U4'�j�2K�/GDM�"O�-�AƄ� ���6A  ��"O8�(��8 �����D[3��郲"OJ���F^0&E{����{���R�?O�=E�4k[3|��m���$ي�I�y��ޖJ�Pl3fU&,�颶dē�y���4��#�2|1�!S���0>YH>�G�4��(��$> ���RȔM�<��N��][�1A(5!K�-�l]R�<a�oP3)���,ײW�����J؞0�=��j֮IB��"V⚱H���sop��h8��a��Ąw'���wN�K�@�+�6��q���'�}:a�L+�9熈i��X�!b:���gl�+��,�PaH����Z�C6�I uay�ʘ+�(%)��̈́��Yƈ_���x!%
�
���盃Z�!�+��l�RC�I� AFB.�ũ*�0-��d+<�H�e�,��i``�̤A;�h��o)ཫ�ԭK*������;���=�a(6�S�ӓB�41��&�=���٤���Hw�C�I� Rx1M&t�fph�!�=���D����%>,x��P���w5��b�$8D���4i��J0��5n�)hPft�B�	0Ԃ`+���y�&m��L�1�����>���1I$�p�"ҳ��T@u�ۤ�!�D7W��IJE��!z��$��ȝdb�Or�=%>9#��Xt�QEa�H,1)��<D��!���x�VCJ�3�I�SځQc��-��s�X��̓=3ԜQ�B�%:���A�$D�y�WEp̴a1�أp�X�Q�7D�P��ő�i���CDE��XR���(lO��L��p�L^$�0��D�`�x��Y��M��4��?q�ˏ-H��p �+H�8�! M�G�<�#�<�j ��Q����Yc(�E�<aU�ص���);xnݢҩɜF�&`D{"�'��M���ShhBy���̵ ���' p�P��%�|�+c$�z�X��' T���!ԫ>�B8���>"���
���7h( �ȁ"P qb�(�<C�I#�8���n1"���X�k�8#<�����R1 ���o�2D;�)եL�����IN8��H��d؜e
�KқP�Z���>D������C��p�CP�s�,���J>D��rfF��z-Z$!��])$���8D��A5�/T+�B���:�*]bL7D�� ��8�-��+�����6D�c�(�1B$�I�1Ly�Tj3�O�O�*��[+:1z󊜍]h0ŉ���}x�\��L5Ya��p�S�A��1b0D� �.؃i�1c�ŀS;��d�0D���SF�^�<�C���8):�x��/D�ؚ�`O�Y��Pw��7%��܀��-D�� 6�Y2kk��c�0^����U� ��I%�hD���K)xw�ɉ��\�U����3�ɭt��X��E^�*��B �pB�!T�5����VGlqC�_�}�C�	 y�#�aT�_�|śD]�vs�B�I"v�蚃e�9�Fy�� Jb˓W`���qD$:�˭Z,�A���I��|�i;}"��h޴�ځG�� �X�L����d9�S�O_�L�T��7m��80g�eK&<��':h!�!Z�lڨa��=q`� "�'$D���
�e�������7ڸ��'0��@S45@�U���1.x:�	�'(��A�ˀ �t�b�KĦ"Yf���&�$:�O����ŸhܜX� ԺT��Hu"O��D�ܹL
�A��h��Z|�[T"Oj�/��q��]H(�Ko�\��"O�4�.ծ�P���F{�l�"O���M*vW$!�R�׆K���17"O�в��L()Q y���R�^�n��u"O��k��m�ۡ�Xǲp"O�iѠm�Er#�KPz%�F"O��1��2��H����b��Q�������p=�f��?��ܒ&GE�^5vTʁ!�g�<��˃3d�|3BƇ�{q����_�<A���S� _��k���!=M0\r@(N
X��b��G{J|��Z�x��&,��:=��p �U��<�
ӓh��]+U���k�$�'�X��h�'�ў"}*@o׸��;r�H*�dx��OS��l�'𠬓�Î�eϴ��dg�+a��OX�EyR��%02$�C[`������y�ȅ�^������J032� q���^�=E��O�����@�'�`����<5�l��iJE�3h�F�L1Xp/E��T�ȓP
\��FڐtJ�J��O���Ax 2NL3]�!)r&W�(*��ȓc�����O�+ Ԩ3B��E
<��Ip�',�q"5h��F8�c��TP�0}�'"6!ˣ���z�`{���r��y�'Qў�}��̰g�h!�ђ0ƞ��&ܦ��iݽ�'�'� �s,�����
�e_j�5�K<��s���@�~,�� ֳP;�0����~2d�&!��p�'�y���a�>�yB	E�o,�#�&�!\�ҥ*Q���'��	^��
dOE7�AgZn�L��3�NP�<�`ͅ1Z4���9e�j���]C�<鶊�}�ĵ�s�U�Kg�dI%
�}8�$����q���qWk�+u�e�J�S~B�O���`Ӷ�X�dT�wP���ܪ-=9���OT�=E�D���S��ңT�H8q�S���<a�yR�Ŧ5O}��U��O�*
"�U�Y��hO?�$�2G�́cD��=`f���T�ْ��~2V��d%ƉGߺ��!	<�m���3D��{�A�B
�ꍄ&n찉�&D��[�EZ�b5�4� L	�8��u�%D�ț�P�4��à����IK«��<a �IZ�'x�С�G�00�Ă�c��!K���	�?�A�WjQe���'�2k�2Ov�=�~��/�4%2y�CbR���Q��	D�'5a�deR��t�;B�ɗ��HI���y�k f閌�v�K'h�#�0<�����+���/f���I���
	!��8��` ,*9�&��p��=�	x�'��c���ÍR�;o�1���-  ^�	D!D�|K���u�D�	REԂDN<ғ!�>��'X�$�"}� �̢�!�QR�"q'�6,=�<�0"OV((�b�:Hġ�ׇ2'0�@��v�l("Oԅh>Ek�i˳*�L��`:D���E�A�T`
*P T�Q >D��R���$(,�RPN�60̝pB;D����K[��nŚ5"I�����9D��A�熞!���C��a˄-�^���4�O�e���^?$φ����c��ɻD�d$?Y�O0��|��L�Ҁ�Q�A�/h��[RI��!�dC)`��@s�'�8g�����!�dG�.���+!��g��s!@C�KP�F
OvH�2fۚXdz��ʊ8徭Â"O Us�猉*.�yX@I�S��uc�"O�P7�['AyjfaX��<�##"Oh�Sʒ�2E<�Y�/�	�¸J�"O �	֖>И�p.��*^��J1"Ox���[��se@�&&�a"O�Q�M�C�,h)��׭V����"O�(���
0�!9��
��x��"OB�A�X3-�ݹ4J]Iմ���"OF��G�}#@���0q6�R"Of�{�EO���KaN�./f�H�"O��)�ȩg�@AT���Zv�M��"O� � ��'Gmr5Q��ZmؕQ"O�:�!A�����ߍ`�P&"O�z E?!���e�#4�"O�:r�>]|b��0fW��uS�"O�52�/G�!���P�D��|��(��"O��[fR�;.Ș�S
 T�rz�"Oj��"S2����.��>�5"O�g�[h�1�O�U�
@�"O\XF�T+c!�ZW���N�b"O Mc7��!J�	�R��NS��""O$�iABވT�\�ѧ�%@ 3D"O*IǄ� n�*�X�G� $ 4�f"O
�����V5�u��a#���&"O�H���G�f�2�+@-YâyI "OxQP�^")*D�s�"g�"�"O<�B1gZ=�0�s㍄G�8�"OdQ�eJ�+xI�1�f�(Y��"Ou[sL��S���J&/J-ȘA��"O������m��y(��X| �"OtE²���W9����ؤ ��E�'"O���DM�2��ɐ���w�2u�"OHٳ$�+�LEYV��&݊0��"O�5����E2j�x�D�?��p�#"OLq��ȥ#�vh袄C�|���� "O�X�C62���,0�����?Oz\���P����zC�X�Y�d���ɭ^��T��I��/H�a�%v0�C�	�"`����u� p0j\]	PB䉫?����b�Ѱ:1���F�Rx"B����u�)��a%��ٔ�֭j��C�I�S�t�%aM%E6xp`-R�V,�C�I�TZ�Q# Z[TL�ªQ�89B�I/v��c�,�5���r���""B��L����ʇ4$PȈa0%ړ	�C�	/3-.���']�4�rT�A$C�	5A�	�0�K"[) !������B䉻5�iY��R6��c���@��B䉠-�����LZ�tl:s oW"vC�/�r�:B㍷@�]�)�zNC�	G>�3@	�,�(�`�B�
`�C�	&Py�e�R�|vm��lL�da4C�<r�kb�A�Q��A��l��4C�)� ��ٵ��:T�,m�2!l�zxp'"O����a��}�^����O/�4�B"O�l�U�<8�ZHR�l @��"O � �7�*���(D(�"�"O�s�E�J	,@[S�خL����"O���u�D�{�)w�V�o��$a���Y5J�����O`�Ab�̞A�d��k��Y����0"O�����?&IN"2lӗ#��5�'j�{���#�2y��I3�� ����'i�fqh#M�b<��DT�i��
��gpq��M��E�x�	+ �	|L�֫Mw�<	T��6T?�Y�Ϛn����͈Kܓj����$�!I��WW!���|�g%��5�\��_	�{��'�T��$I�	<j7���gK(p#��j|2؛��8Yy�رRa@7�?����|�G����'�H�d��%����C6�@��L�8�`_m7��P'���6�F��ʔj����5y�> ���C���;1LL #m(t��B }�6T���'Đ��0�@�A&R �W�Y6K�\܊�ɸ	��	�g�$�JN�&�(��!�	��11-S/��0sRN��qBv}B��C�Eb�A���L��ɝH����ֈ�w���1�n�<Kp�y��n��pG�Q������c��p�v�p����{�)�7EsP$0�#�'nn�""N�91�=n.��9��m�q��:ep�ܘ��~
ւ��.V���E��1C	,�gP�d'@��EN/^��0c� BPy��#/R�ܢŏ�3��^���)6E��r1"v+]_Q0�'#X��иp�5���,��b$V>-rL����HXB�?��,�b` '��i3c�<j�����3)|L]46��ػ��'��8�"m� ?���%g��{ь��+�@��ɺ~��t"�(Q���ЂM#8��G�%f��k�l�)�>`׮�af���牭]��@R��'�<� ]�1X)�፝3$�8�E(w��K`a��q��1_�6q1W� <2R Q6A�2&�;�� �B>0�@dA�F�H�NA$�X��O��Qw"
t;�p�
ˡ�v��� �l��P�S�qc���7��2�Wmqr
4Cv��3�{�!�UDZ�F�T��yb@;�� �8���Cr�����T�2�0쁔N_d�xɽ|� �ӸB�IC�&s X��7g�&I�d�s�݋:m@4Z�g�|�t����!;�ұ���'���`hM��uBHA?C�ܳ�.�� ��TL\'U��cM�<*����H�K��A:�h<E���RN�A��K�%;.Z��ʤ蓾��
��B^�|c��k>Z8T�${����oU#^:|%��Õ E�i�ȉ�E�B)ʵ#�o6J% a��z���	\5�z��Ťc�&�����]G¥�@�d��yG�g�Eln-iWf��G����m�>x��w�Ӫ~��Xb�d�9#3~��CK���uj���OĀl��6~fR'�ЧW��#<�Df#j"���f' ,Hr�� !|y�#�f����{�<���hZ�;:���f˒1:T̓;�~3u��3�z�fD�[!�pC�O��Q��5���ZX���ȧY����.ӈG�9����),�\ص�N�X�6�0���!X R���L�X����E�S�A�	�;R��8�G�͑9t�����?[�X��S���s
[
�ʝ`�Ҳh5�8��>���( ��s�>�����m澼��J��޵(��Sp�s����a�6\钨ߙX�q���at6��A��� �:X���Q䄹
����b�	?R���
��ҮM^���iL�.���+�\R59�`U�vO�)���ӓjx��O�(sv�U�"�>�8���( j�:@��0`{FiRBO�P�<> ����u�}Pv��r�<Ɇ��: �$-شE��C^����(��je��c"˓JV܀jT�I��B	ᶦ(�i���Rͻ �ļy�)ƿp
B�Yb�4y����0l���V�1�^X2�,��2n�1BL2m�v�b���F�H�b��כe,��F�,�(O"�# �	}j}�J��<��4�'�0��v�n���_v4�P�E�.:�@ADy#�<[9��ܻE +������g�Ƚr&��G�n�sǊۜ8��'���b��T�<{u�fL��R���
$(�q�Ve�3ן�����;�T$����>s�Ȕ�S�D߹ff��!�)!��hp�ۑev�� foO�pD�q���I���=�'�e���r��۔+"�����"'�(#����EB�}'�H�0*܅s`�F�Z�	Z"��g�'h�H$>$ʾ���R9@�"Q����
CO��;bLʃ.s&�;�*S�/�~�p�$� ®(�b�R�B��	�y�&�
��@+	��B�ܢM���A	˓W8�%�:B���󂛥Ufn��2#��4O����X�FclD9���.;Rk��X]z�EfdH)��O��Y2�(�Ӽu+N��W�1O���!e�Г+�OFQ3�I#"Z��n�0�� ���0��jbU?���hP8��@ j��f����!E�����P�x)���	$.�g�<r`]#�,���S���kz�=���7gI�u��\�~�ٹ�����O��L�m�=���J�啖=n�T�!Eɇ]^�-�c_�PNu�U8�D)��6u�m��d�cx\쪖�Z�>�)��]�jG�,ƇE�kZv<���1t�m�K�etT��'�:�!�
'(����V�-XX����<�p<Y&��1�nq ��Z�c�Tͣ�)�\8����-䬌�ʖ[��Х�	�	�fр�nk��2��1��DD�OM�T���
;�Đ�EƤ�x�_�0�2#���C �%Pl����S j.��%M�N���#��i�%��9[�`A�4)K85N��8P�?�=� J�*��˥{b�S��MT͐�0��-��L�� �K�x`����Q��Mc���?�k���!��d�YVP�sc��=_�t3Q�I3=hy��%%\ON�P��O�"ªe3�T:&�u�aH��l�RL�7 iJ5�S"܇��L{��|B�>.�Y��J4��I� J��d� 1O� !�MޟxQ���d�MA0�T�#M���'R K�)XƁ�x8@pP�ߪ<��{pf��fؑ���䅂���g�#}*�w���#�`SwOt5�� Q��0���'2IP����9ݘ�R���W��O�9����F'@^|2�*�Qk,8@�N_�H+jt"�e����9P5ƃ ���;��4��������EC��HH��hőoc~@��
�8BX8t
���/�@ʧo�u��d>%��:p�xQ,۬M�4���^���W�ƶɆ牆_��s�֍�(��VaM��(�bʀ('Ӕ�P��)i����O��/��BbM��*��;5�t�{b�˨ ��D�O��a�B?[�.�{�홁@@>�{��$^�ސH��^�V��	�F�A�$���X��M���봡��-�����z�,�-ϳHD�� _.9n�ٹ�- ���֝ܲ���N}t�}�'8A��H
X�u����82� ޴(vJ	�� �(�"����$�d0��G����2�S-8vhZ!l�)v�-��@ۂv����hB#F��Q�Ջ[�J�1(�#O�0"TH�\�ax"˖8~Y����5P�2�&�
R�z��'���nvjP8c�Ītf`�`uk�9|\����gǇ1F���G
Q�~�ӷd��|�ڦc��,;��N�gN x�Otx3L�2��'Ć�c懘��X�x�K�%9t|AP��z/��F��s�2l��'�@Ɍ4�7���b��H׋B%8zba(�,�'��v�[p�:��A�O�X�6��(�v��u+��``t�=��ꖱ:,H��2fP���\.]�r-�p��<m��B��O��k��]������\pY��I�5�I/LB��Q�.V)**�Xb �<a�'́b��]*�/��W�dT³M&��6M>Ic��F�U�Or�!�DW�ξ���ޝ�%�$8ҐI�����g��CUOH%,��qwH�L�p� $�9P�@ʢ���M����/���I�-��i!��N�v�(�������ی˦!x"�0Q���´[)J3��0�[�w-�)ke,�-MH���$�	º 碝�U���d��)H9�q1dlB��dR�L��z�έ
���~Ð#eT�[�n�1L��<I���O٨8r�ƅ7]��f��.b�(U�&0tl(c�o���
&�
�P��|
�cƄ5X���檞,f��09Ej�rh#ɂ��p���I�b�,1�1��E�>���W���E�8��pk�+?���V)!;��b�I������A��a<�jF�۶�vh������
ic�F®c8�Q��-�����Q��4e2�z��ڵ�?��gLD�K�� �Ľ�I�)w��'��(�o���*'K�.mX`�`럁!�©�	�z����f��MC0n�qo���Pgݍ:2��*��߶�XPWf�x���S#έ�?y`ID�O��Z `B�5t��A��{��!��!� >�	�AV���`��m�(��2� ��3`���z��-��1�V�c�236�U�r�H6�\t���- 3Bc4)��T�`nDl��3��=��(g��'Zz��uJ�8���e�[��%�֒.9���O\�_��:��Z9�~�b#,U�С���دP߸��aHV�h*u���P�y�IB��eX���f��6:�
#>�O7MH�h�q��4�&xB�&��z��,��lM�].j	�'+��wl�y��II��@�E��"��Jǆ�}��4ɴ�6[!|-��!ui�ixm�S;
���[�5+� `�d\�	�4(� `T��4p���,~��q�MGN�)�m�Aޖ�f�A IX�P��,�)����n����P ���ޟ�)!K\%?�@�γ	0�P@��Ō|���A���0�����M �R��
ə7��1���O18�LpĎx���i�)��p��DA�@R����(Gڑ)�H���	� �XyR�M	G>�g�~����I�^e �㤁ΖHG~�0�
��,����O�pzBk�3P��l�T�ǭ7��U�0�K�"�fc�K�R��o��a�zEdQ� �f�t�L��D{�X�]�P9DI#����MC�X��#&	d��ʔ���]h礐���<J`�z�Z�cq�ZsC�p��ˣ'|����>Zc*rpp�#"�^E`��9}45X��x�_:<z�D`����ZY�	����sG�������H��	4qA���Ѧ�n�pD9�+�
#3�@W�Kn����_�R�q��9!X�O�ʼɁb +�*��p���D�6+�%�5�R��
�%
a�:n�ڔ��OBqP7�Ћ&��q�u�wl�����7����Q�G�.��()�&��(0��T�N6rU1�I`����F>/	L�`�@�',r|�f�\:����B`�%�I7e������L �bR�3.\Iir�MY`J�:h^��%�ۊ?>A�f��iֈ��eQ�hOvE���΍D[��S���1�M����:M�`uC���)ᩘ
uv��a϶U<d}������Y��W8E�Tu׆���Yy`�+��[�
U	GL���eGTi�I�M14ŋ�Ι�W/�Ա�#.醔�t��<.嘥Γ+u�S`�W	hC�����'%{��{%G9�h��&D��>AQn��=�M3`�,ےG	#NI�ԩ�'�����v�҉�3��j&r �3H��0W�\�?�0�f�ǀ;���	�u�¡���ӣm/j��\���9���Gz�P"��k��Ŋ���M�`�gO n��V*].;��E|B�^���S�]?Z�Q3d�K����e�
�6���@e_�@ƶ ��
����)��%r6E�Ey\К�j�&9����q�zUj��/J�@�fC�'�<5:���S����r�O�۳
��¯̶=D{5͋�(d㰪��.��|˓1Wר�� b��4��̷;HSE�xD(��GSA�p-ǜ2�Ĕ�%�P��<�=����(Cn ڒh�m4��V��jt� "+��P���^�PQ�аw�����3ti�M���K���z����(�<F��M�d�<V\��������s�Od��A$S���ɑ�P8�7�F�C<�� )�#��0� ��{�|�����舁1��BD�|�p���d��5x�T���H�R��-j��ŕ-V��㷝h�d��ݠ�J@�"%�N�'Cz��7%hՈ�/�-r��c$W.{/�Y�N���"�)@�pKtݢ�bZ�l���/v��kWD�|]|y�vi�V�N�"4ˈ�j�2���e�6n�t���T ZLDd+5�ݝ)��Q۵'A���yE&�O��+&I�Zu
x�j�RnB����]1b��}��ǁ����iu��M��	F��^}X(ͅL�LA��@�&��M	Ǫ�R�dC�5O��b�T""i�� �\�"-<�I�+�RzrF� T
�`J�Sa��AFY��"E��x��P��$\z��!�P�-WmZ�=�����6?��1jV�s0��43Xy�X����0	fN�#@A��66PaА
ï:X�	���U�jeXsU�>�SZ�	f@� �����KE�	@H�Z���[�Ѻ�����'�&��u�~�'J�-zǡ�/Qd�J��Ӳ���W�
�ϐ$�"%�-#! ��i��M17#�ӦM�ki�!�!K
ߦE)C�&Z���'`�,*�Y2�F1���PD�O�'�-���[�0f�8#�C���w�����8#K�-!v`��w�ћ]�`����1�x�����?�U-V
���SK�/%~p����_�d����*�R�	�M�81��܉���Wh����n�̑Q��O�XՈ�b�/w����I��B}�X�E-	)1�Ht
N"I"Jf��y.��ZG��-H�)�� d�N郧��)vvz���D� J&���>[�T�֧Ñco��ے$Y?M< �e��ny0i&板,I����c½^�@8�F�B`o�՛d�=I68��E�3B5r�Y#B�3}���3ԒG��c�#�6$�5��%�@�cV膎?\�l����hF��*�+y0���%�+R����H�r�L��#O�9V�@���lO��"��� }9�6�)s�m;r�ڌ�xl*�Q�,}����$�=o@�}�A�\H�="��ϼ������L2&�
�i��Y#q�=ѵ�]�S��;��@��R�Z�^*ܭQe��1�?	t%|�	���Q���)N}2�Epe
�#h�`qar��D��U��QP�`�	��	wi��5�m���%x�8��[t�����Æ�_�h��'IL�O�,Z&��0Wjj���h�?�t��a9u�G+]�l�3��1{E�X�T9vd�m�!�۲f5�<� �N�+�F�'�9KF�̲~N�0QM�;td�E��a���⍰xM�����K)���2�+Z@��f�^r��"�;-�x�K�"�h�I,\�u��5;��S؈���eΆ�ęC�ʟ�g�.و�m�	R�D �L]�p��sV*R�zێ��`e�ğ�w�( cdE���3�P/���O�#U��.,��TB�F�mZ���TJ������-� �0���\�:��%�]�����Ӣ H=�	R�g_���)�05���1X�4�8��������!�)�w���aX��O�[�b��=�G�$z�aqGKW[�tX&� }9LL��a�s�b��R��>̤yX�}�bA��!ߓ*I�E��l�O�M��&<��de��}¢�2k��(K=ӂ̠c\�'(�#�Ɛ ,���sm�;��Y{��81l �hK=׈Ԙ��4$/7���>?T���.՝R�3�䚆�\�sCT)�TՅ鉍b���q�ֹ0)^�%�y`\�c�+G�Kqf�3�"�Y��A�U��x@�$'�82(\�E+��{e^�S������cd�5�
m(�ƦcH08R�^z�'��2��� �*��ty�@��\:�d����9#��c�A��[ș�#j����F�Ŀx+0��B�<������R?9˓�Ϋ3�v`�dO�hMȩ��c8}2�I�sӘ��O��ʡ���d�G0f{P�9�G\"x�$e)����i�dŲ'@,r{�!�O���U/� ٸ��e
�U
��!j��u��R/xR��J�^��o԰K��8��N�F&,KE�U�.�D��$����a�{���sF��sz!�DĜU �T���M���co	�q�!����Y���ƙ��(�!q!�X�& ��xg(ˌ)̈IXG�(h!�$QC�5�!��2�`t�p��	&^!�DA%�^�bf�>A����E�0d<!��	�R<XQJ�1�x�;���2.!�$��M^ꈸ�D�*��]��hW?/�!���dD� d��o{�Ĺ�'�q�!�D��}�I��g��2<ʷGC�V�!��Y��AH�#��?zV�K �:j�!�$�30V܀�G\ ^h^�3�"ƍ!�dпY/2��	��rT�MXQG�!���$eZ���B�=[�!�EF>	!�Đp����}Al��G�a�!���e�����n�<97M!��/X�!�t�L$�rlD�_,�T
�i��?�!��A46&� 3% i��	e&ڥ0�!�D
2��d�%!	-[�@aa%�9b-!�d:����p�Xi��5C��l!��E$-���0�
���qD8[!�d��Hd�S3�)s%R���ܒV�!�dG�h�2:
�/�>�0s �gd!�[�*�
��*n��D�%�=�!��\&Z�<@QRI)��@Pa�s�!��E}��1oي.���tK��!�$ �'�*h��
K�1��Y
R���PyB莞I���+W��Bz���稔��y��hgL89�d�#@�����yr�ETT��ⲁ�yЃ���?�y���K <Ձ����@Yt�"�A*�yb��$"����S�75ΐ��DL��y��Q�|8���� �,��`��K׳�y��C2?�@��i"#@ T�2���y��	� ��!� )ΖH�qz�k΂�y
� ��`�BTr��𳯟.T���(�"O���� �nH�A�� P=�X�E"O���1(�I�!���	���XU"Of���h�!(��h�e��2g�|8#"O��ò`�P�"��IE�yk�Y��"O^)��#�G�t$j��Φ2K(�I�"O��w�\oz���i�@"�ň�"O<	��HP��hW��*i~Rq��"O�ax�X�G�j�0&��; ��I"O4��b�?=)ʶ� V Hb�OÙ"�)�����O�	�G�'>��pt�Ë#W�9!�"Oʝ;��P<ƚ��UJߔ{G�tB�'=]�S̙�\��I���cF�x8�͛{�I��@ɽ)����dY��<�g�30Ď�ل@\�����T�E	�PT��W�<�vMX�Q�pa��	�/x4�ï�v�>���7��7hĠ�J�+3�'xn���Z�M�x�sCÇ��	��	9M�|�{S�x���FS��I%�ߞiH:$�� �uO�!����W��陖��O&m{/�P��':�	����C�R���j�1*K��'����!bV�T�}�*�+H��+�)��V�yKc)�3v�(���
*��}xX�0�V3׈�9�䔅��Yٔ&F����
,N�f-1��Uy҇+J�6���� �gS>����� =u����KҸ_F�K����V A'���Z����D�
�/a"��.,x�:��Ã$�$y��j��@�1���.2�>4P�̒�J�b�!Tᚁi�n�Zc/B�u��~z�+~vp����H�õM�h�@Ҏ��V
}�| ��ִΪ!����H���'��-(�UG�8ʷM�2 &Y�0�N�ADjA#~<�Ԃ�&��h��4��͕�\@���Q!
�pF�&	��	� �P1?� U ���@�4������a�/v]@��֮�:�Є%�($�����Ĕ�f�`�����KSV�z�(	x�����[G3�ѯr�r`q�-ϭ;U`�e�'���iƕ!��ܪ���_O̜:S)�,u�vxq�mO-<Xjp�2�Ǒ>W���#��^
��&�Pg���9�Iʢ.z���o[f��%�2�� G�X��V�	���0V�ۀ,)$ D�M�m/t�� �Z�d��-�OԢ��U.Á:�h0uD�N*�lʄ9/�#?q��C�'Ph@*��$g�u��OiƉIC�70����N�+,���01�<�}k�k�&� ��r�	�uF�z������)��4 �*	�A���AE�)�a�8X�s/jr,гn>���� ��鈳G�(���'Cl
pe�(�l:�� #�/h�v�9f�
?&�ll����1E@�6/WZ��x��O��0��c�U�t%
Xѕ��x�� 3�LC�>�Z�{��A�[��Q����3�(����?t(d�Z'}���R�dO�(����F�%E��b�'�O��@��ɜ}��qF͂;�H��kL�n&�A�gn؟vb��Nʖ.�����Zy���1����9�D��̭o'�I�7���&�RL�VhiK6>�F�*Q�3�BA��$��/�*�[��YXE�%w� =�b�&N1>��@�	�]Q~7m�%^<ЃD)8�%9��.J�"QJ��Ɂ;�L�A�o���`�m�0�%9Jx"� �"4���@�u��s�c��F:B�{����x`�֏��;�0(�� D(�YYp�Gv��1�%L���2(�\g��V�
q�t��)g��0ᡢ�u9	EQ$N���"&H/�lq�cq�� C�<�nb�(����@� f!�D�P���!���q��A�Y�b���^0yy1��<�U٥a��u�D��eaS�Q�C�$ϟX� �r.�� ���p�6(�axA_�pn�%�@m^~��iV��.t� ���f���+'���8�K�"sn��ω�s`hU��	��D(g��( sܬرU3��'A�qu�2f�|h;2 ׋躰S�$QH��J�?��+�00| a�V�"�z���8D��wƌ�@R6���g�Z~$ai��W�vh�HY�Œ�|rR	�Gӕ�f�g���'R�j�]�)�B�Iۤ:�p4ru.D-O@��ēf"h��#i���#��K��YP̌*D�8B���9ؾ��d ��,�B�!X�<)��D�	�Ţ��
d�hQ�G�HX���E�2�������i���f�!~p�� l�q�N;Z�y"�A�l�	��I�B��MY'��$h�ą,O��OfA8�d��]�B��׈��,���J2��G����)�?q�PME�((�ĳ�΀��R�ȕ�(F�^�BU�'���P���~W|���E(J)P ��
ق�l����:�#����H:�f���@4�
F C0������%��)c�S,ZCH���0?��K/3ޚ�.�0 A��ގ2��JM�-���I���[y��x� ��7֊�B���6U�-O�PK�S�K24ȣU<	:`�0�BX�lp���}H�R!E}l�h�я��)�3��#z`έ���"�H z(�9�!�w\�#h6�#�'�����ĻF�H��NJ�E��39�'���ʍ?kh�(7 H�h�j��0�ܡ@�����ⱒcoް~��*�m��lL��s���8����m�2D#�����3�I=N3V��S>��B�ǟ+$0���T>��E�C �6�t���b}�'X?�LAAA%���fC"6���[��e*� M�l�0]B3�O��k�j��9>��F�g�@�7 @U���1��k�uP�NԀz A�*=:>��v
a�N���T���� �=*��ڽ!�.�*�j Lej5�'�(��j\yZue]�B�ԝۗ�	� ���I穖�s�r�e]�|�� �Hq�p=a���UY�7m��(��A-3�����9�-��$^��'�!���ڥ]��x# C�o�Ol��a��('C
��Q,6���8u'�ޅb�P
s�
�
�ȏ����D�[�@�@� �/��� ��%�Ր��D�%P˓;v ��|ʢ#9s
�Ч�W�>�v�:ujĵ�nU���A���1��V�W�LP[ۓ&q~��u��d�<�cpG�Y 0\k�D�++�	XV�ÿt�� �5O���a^f�(�#�g\	>Hs�T>�� �ՓS�Z��T)��|�$,z�	)�"^1!�ͅ>O�`���"6���� �U_��@Ӏl֦!EjqC�D��?(d�Х6	�vMZ��5AC���BH�O0�.9&��\*��@��$C��;L�H%S���($KK�5�N���R�$��L2%�:���w�p�Y�	�Y�J��M�vj��Y�
�� x�u�U�jw��+'&hݩҍ�D��[�J���IN�N��� 1E�śEnl���ti�}
.1cT>%h�'�%{��DMd�~�sV�J R��k��^%'h2 ��ӈdR�b��yx�(ӤE�`Z�0�v+H�B(U�#�X-��qX���j���@`D��<��b��چO:y��K	�L4U��aY���a@�T?�:c��넄��W ĨF&>ғ2�
�<�T`Y�'�Ԩ:�f27�n=��ޑƆY�CI�@`��$F+/��	��왖?�xIHd�O�-@d��"/^�uw�%X��c���I(B����.Ó��a�t�ݎGA6M1y��A(B�=I�~��(��U�n1�W�%,p�Ӥ�;��u17�m9B�K3%48��D�ʛb���Q#y��C�X�tAr�0Y�����/hŒ��1��8��%��n��~'
���LX��B��q�ځZ�v��W���j����Q����	��N֚|+��6L��q��PS�P�N���Y"� O%��O����N� ��O�́a�ҋ1���vO��]�Ԁ��
�B[hu{�@l�x�ɕ��Z� �qDW6GNM�v֘[�ʼ�5ʒDQxiS� To�r��U��Di��@A�v�1ǬM?_Vt�r�{��߮(2h���R��46kL�``���"#WBt�3PHS�!Q���3��>6͖�gڲ�?a��<9���[��	Cu�#��']�ċ+Oݡvn؏����`�4%�V�#W郵�M�!�C>}� �d��}� ��P1���|�X{�o�>w�*|��.Y�����`��02�Ś"1��!�0m$�� �mm�ĹP#F��~Rb�b��R�#3맑-, �*���ܰ!��	�m;aЀf�Dx�@�����@_�8	pV�ħ��б�	�m3q�P�\F�U���d]���L\�p�E ��` f+B�ZO�@��Dn�,O�L�¤��t�kBa�"9�89� � 7Ԏ�e�? 4�kBN!X ����*V��K��=!=�y2 Ģ4҄���!:� ��W|�	�W�C���b�x����*?��'�t8�FbF�<��mq�k WƐi��"h"T�#E�[KO�D��	 �v��qC����Q����H'~���+�5pV�;��[�HN�X��I�p��E�P�YYpa«O�$$���$�����?O$��T��J�*�ji
���q����M� (���.!����1��|�xc�Z�UC5�U�)��Q�g��3S��r����^����ҏ[~�E������ye���i��p0�b�,y��ѢL�Sl�x���p)T���A(�ν�&L6l��XpG�-y����}�!vG�*���x�a�l	FN�O��H�A��upVͧ|�<�Q�X9s ��P�0p��J��=]�yKag�	�2A ����Y�E\6s��Ќ҇6}��aaZ=\�u#�
�xm��O�<����`�%���H��V	�~�ۋ�d;z: �cĔ#(��Ɵ�� ��h��>�<�V�8Rn�iP+J3\� �0CM�l �e!����hC�;� ���'d�A�ϧB��e�$A]Z����!�\��'����!N�Y��HrDꚧL��@_�h��5���F��P@��@�\�Q����4)MG�$0n@�.1�����O���C�P�Ґ���O+���Ye-�%&��|�B����2P�ܝP߂DJ�/̧(�2t�Q��)����	$"��\�o��?% (�G�	4@�b���
 G��C�'L�.�L�gā���d�
� �T'�oʤ�ȱ�N�a��L��A�3KwT�3z�!35%˅H�}�3�5`[X�p3g�0WY�T���Y�j�pb,N(�B��5{�(AP.F &ў� �����������;"BkLF�-������sk�t���������ə+O���s�O��N���J�,�����mO�ue�L��OP��1q)�%��	5<"p!A����%�4��:H����Aݬ,���.�&�Y�cT[?�(�1G ���	B���3��U��(��Mn�X� �/
1��d٠k�h3��a��2* :��W#G ��4`�K�д��Br��	 �Hy���Ie�pQY�4�Ī��re4]*C���r�H0�٪
��R�K����E�O?)W'�]"�� ������d<|OX �p� �0�� B'�<���$D���<t.9�g�E�'!�UX�����` ��Ӂy�^���4H�P�+@�oA���h^>d0#	T�ў�@([.���j�e��H�剛,Pl$�%�Ӹ1����M��4Q�������[�(�S�
���d	�剘)X| ��S87����	1]��ђ��l�A��E�(.�����!ŷ�ēQ^����ji�xS�"��t9�%ؼ<<2���'��RdhT�X�b���4-�����#A�v�ie�� (�،��̎_n����6���z�eڙtj\����O½�ղt��Y��d-F��&݉|Y@�M��tj {�b�h̡̓p��yA�!�1b#T5����
zTDŒG��0F>�a���1(��D��yfs���zuUc� C�*MNՊ���
�Z�C���x|�)څ-V�`�8���"��� _���IUˇ���)?9�
ݺ���(X?F��W� V��������D4
�	Q)� �J
��Oډ���"2�n�@U@�T�(Ys���5�� ��U�ގq�@jR4R�i��J�{@}��m��6a%�Z�� � P�նۀQ��ʓ�T�-[@A����'�1NфSU�䘧i���%mX�wz,���Ξ>m��,��WҜ!����9��Y֫�J��%�6̓F]�q �d�ވ��	!l�$@��^�4��v�
N���B?1��F�j����UB��/�����m��Q�`���I�?Z)���J�J��)Ql�i�����b*����4M^V�v����n�Hu�ƛEl�p!�i&��F+4PCb�DF��&,�F��IN4Rtƀ$�T�ıp
���R"Dg8��∶g,HS���JD(!z&�$�h[f�E�q��$��Ut=1֍�8$0�X3��@%H�Rpq�P��0<�1$�j
2ij��)<�� �Ǫʯ �E�����	Ba�3v���bPa�1b1Ja"�;�J
� �I�������1�a�1r�<�C�M�4�ƥZ�ϑ+vtyt�>A�⃞"U �2�u϶�����V(B%�,��p��6s����^���I��>�0C�[�R�ND�@�K!����q��	7S��;�4h�q1$ޞ03,�w�:c��	���G_?g4�K��M�x������������sfS9Glެ�i�|O4d��ϟ�<a8�cf9x���(P1O}����DO���W�A����7O�X��L��O<p�� ~J(�	D�G��B}�Si��dO�����@+d�pLt�&1�,I:�M��Ǒɺ����M�L��|��D���� ?H�X;�*��7�~����OJ��4 �,PQc,Wx��� T�<���H\��A��@�╢
9=��[n�ʟ�y�N.��˳�=D�J�X��S�ˤ�J9�?q�-Ŗ/�V�qӥ�G�fX��'�n?q��-�`J�#4?�|-���K�U�������t:8p��n��i!������df=x�7'��sT�Tz^�AFVf}ZhKB���D�B툧��Q��ӣ��n�' �~�L�ʔ�?��8y AN}��׈1�J�����~��ǀ�z�X4KJ�?��xb �V9�,��T����cƀ�%h|���J�̰<Q�,�&O���CK\JGԑCfd6;7�����(>�Ƶ�Ą�bN\��#^:hR����K�LDн�� �;6潫�o�~�s��A�X����DE����ީՈO���B��)q|��0!��Vp����[�)�n��ŀ<��k��gɻ�W�
�����L	1	���a&?M�~)��Ȟ�@ˀ.mՓ�K���Tc6$�4ؐ<�$װAa�4��9O@k�H�7Cl9{���H��XKF$A6Վ{C$V2Dl� �4i	6`I.|����z2�놢Uvy��2���4Jj���o+P� 7'	�U">`�Ԇ�?c�|��b.B��ch�0?ǜ�kCg͕Z,��:����>��s,I�4u�L�%�[�D��c� 2�%��>b��
�-�&� ]ˑ�ۄ���r��UW�B�S�ްAH	Ǔj	^Ei�$�'k)8 ��^=-.:�O|ت����� L����r�c�j�7�K>m"((�m?(q>!"��xк��B.;�@���x�լ/���G|�%�! �Rc��+�������q[f(z�I?_a�	��n\�4��df�={�гe�زk��AQ��/Kk�����H��(�Vn�1�����<z�4�R�=���Pi�,ۋ�"�(���m:"L"3�4}�	(t�� K&�0��C�5c�t�7�� Cz-�Ԃ�*t����V?^�x<����$	X��'�)+lB�ǂ\Y�L2�+w�g�}��v�ڍ
�@�� ���]�g@�a6����@�`�)ݥ ̔)C���H���N���A��i��$�]�tbd�G��nx6|9��K0)4��j6LO�.MĮ��4��=o,mk�NF �!��f�O����f�7��QD�Z�Ii���d(_>=j&uSaA�F!�=��'��� ��1F^\q�DL��r�٧�ɘ[�ui�)0`�dY�(9�G	�s
R�Yǂn���Y{�x0�`٦�hp��b��RyR&фD�Y��~C��=���d E~n��S)�f��X6���hM���"g�l��*Lȃ����*AzHm��!�{�Lt��C�E���L���B��/�q��'�)A�]���"�>@�P�'$�<�J^�/���C�#�($��q��
I������D͒�:%G�<:�x8��Iə;*PB�	�/�L�H��@k
\�aHG�X�\B䉖3j�X&BQ��X�%ٺ6~C�ɦC�~��2D͓'U�`f�pbNC�q�6�HW��	J�\�t��\C䉐Ƙ����Ffd� ǤibtB�I(Hx�%�a-ҏn/:5 �-ؗ6�6C䉐1�4x�ȷ}+��
��د}\B�	�f^\
�c/l��y#o�'���Dl�x�7�R�N�|�
��?- ����V� ��n��b'd$�2��w�M��'��	�#
%P���ґL�ִ���rL
'���S)P>D�ȓj�t@QIˤ4��m�&�J��F �ȓTyxG�T#QP��[#'�T�%�ȓIp�x�E�)��t�$7�P`�ȓژbQ	�hG�c��ٷ�����	?�yU(�)o������,~��L�ȓI �0�&���>���6�O��!�䞙 S��R�&�����
%�!�Ē�o=��[���w�����Ǖ�!�6p,��si��l��,`�m�	u!�P0��d�g��*dB��@
�5xY��91K���ެqT@������(�x���A&T�$j���.4D�ԩsL_�1���;A�<��i��n:��aK>��N3��i(OJGziz�O�~�t��+�F�~�v���O&�<��R�E$EiM�m8M�@�˪Ә�'��OL�H�h�2RJr����αB7��;G	���B��4_u��aΟ�J�� �O���Y�)>5��A��V�c�t\�C��� ��@c��4j0���[�]N�tP"uc�z�,՛���>�؁��kG�R6�5�	=	Za�td˕Ry�|hE��~�>��`O�"F�X!�g�V�^��S<Q�P"J|�ҏ3�� l}�a��2
��ʥ�ԡszJL�w�'��4 � �(\[N��R�ل�$�����	�a4���#g����$I)Nk���Vc�,<s���G�(��[$��P���bվ~]X�i0/�D�>~\Z�a �O�:�E�Z�|���L�7�v�PO����#\Vn"�O��)�	]�B=�9Kg�?S�@qkP��~���#�O4���I<��o�L08g��S�0�AG�{?�p�������&�x��Ɂ1i���g���g3T�c�����֌_�p'X-rN<E�䪊'�Fac�	~�T-���$�<Q�o�P�T"�h�	�^����Rp�\��J�u�4�3�i�&�z�"�>yw���S�H��H!7Ě%V"4��'n�V��yZ��|2N�O�}R��OyƔ�,,�d�NÔA=�X,O����R�OQ>A��/���T���L��i�,�O��	u�S�?�`�(/�]#!Z,S��k�'������Ӭw�m�7�3aД1c��P�*⟐����~�'FPs�\��ᘊW��˷&XE��
W��Ï}��� ��'6���gϧ@�p�Ja�
Ut�E�@�L~�x�O���"�O�q�d�y'�hA�$�	�'�x���,E�jtzᨑ+%�f5�	�'�eP���1^,�0(�C�>"=��z�'.D@�bԴ!U�d�S΃0����'P��@��w���'���",��
�'F8}� )��gO -H�Ξ�΂��	�'7T3�^4^S��B7�0	 ��	�'Ϣ<D=���W��38�	��'q>�����2���Fe�(+d0��'�p�R������(M��� �'c�h��;a����U,D:�
�'���
�M0�
2)�>Cv��'���R�n\N-�� q-L`�e(�'�L���S¤ ;#n��lx���
�'��s5h�Jd��'!"M�.}��'�`��c��&�LYd�F�?��K�'� pt
��/���;�D��'% }��b|مMJ4�l���'\�0ꆩ�3,���!�>'$r��'Y����&��peE�#%����'H�ԓb������b��Y���в�'$�"goėA��z�Cb��J�'�؀�7�[t��Ņ�\n�]C�'�n���'�56�$��e��2b*D1��' DY5� R�d���l��r�'��l�֪R7{�l���/i}�a�'_���o��~4�� �#U�b �
�'���	�����L1��Ă�@9����'P8x{�GM�]�����9{�%	�'Բ`����6Y��ⓉJ�_�J��'�J��u��	X�6 ��j�!(��[�'_pEx��
DK�-�OD0�Z�J�'�oQ�Hu�Q�$ˍ�N�:�'��ڧ�]�):�(س����%
�'CP��ʈ$J��i��������'0�`zG��ߤ�K�M�,2�P�'h��t�I@H�4
�54��k�'�-J'�Y!FL�I�KW�==:�'w6A�����^l��K16���
�'>�) ��� )�=�2l�1+̖��'A�,�l5|i-���E\����'�%��oЕ`4���"-�,f"�Lq�'a h�Wʱ��yXbbӔ\��)h�'��iq���2Q��M��٭V<�	�'Ȥ���/��|?ؐ
�9;�(�	�'a�l��#�K�za���	8�D���'�����ʍ�ծY�f��&8����'mΘ�"��"F+6��N��(���� �$�a�'0] %-C�m���w"O��z�/ogB$x��;<�6�U"O|�`P*F%%8,\�UKR�Dj"O�����
y@�a*P�<uI0"OμRa�Cav@{�J%�PHk�"O���ׅ��7R�"��H3rs�Q2�"OP��k�0M��8#"_zBa��"O��B��=���(u4��"O ��b�)S��y�RaԹ]px�"O<}(rU��������N8�ȩ "O�9�b�ۃtp}(��_�<�8aU"O��b)Ϛ_���͕SҺ�"O�@ P�o|ΐ*�̒��"OعR6#
F�d萠л1f��'"O���E=kόA��ކ46��bU"O���N&^bEh�>��Q""OD��J�0�p�eN�3|L|��"OHq`�o_�:
�r��@-5i���"OڜjuMG�^Pf����	R\1"O&=ĥY�@Ȉ��]�Z��"�"O�#a��<?�9��˲E�H���"Ox�+���zv�pC��� y��x�"O�]T�Y�1��A���J��#"O�1�c�3���V-�򒁐�"O����T$Iޚ�Cm���E�0"Od��!B^	\f=�D!�8ߤ5Q#"O��U��8wnMʓ�E&;<r���"O.���.B/MŊ��I��q"�,��"Od1�4�U:�h�Bg��Y�"O@�XF���t�E�e�w6�Xx7"O(�6揟f#Lt�tj&@00+�"O����
V���c�*�/-��"O��J������zri�#f���"O���!�"JT��aЙp�IP�"O��c ڻ'��Mʁ"�$"O�\C!l����.����T#�"O���;QL͘s �!u����"O�� E�<����Z���y0�"OF���웶a ��T�O���"O���HG�9�Q��-۲}7D��Q"O�y�����c�m�5D5J��#"O�H8!YE4��!
�5}.�u��"Ou�$DK� FN�A�F)�D�t"O����I��<�v�Ŋ=�e�"O���I]ɾ)������H�����W�@6i�]�R����Dd���ȓG8�x6L#}�:Ĩđ&"R���98���ˇ1���0Qr��ȓJR\�r�G�&JJ��'�Τk>v��ȓ9��б%���{:���!������]߲1���˟�|��q��'D��ȓhL�*���0Oz��)_y��(��"lPi��'XZ��y��!���n�D���σ3ꂈ2Rcƾ.O�Ԅ���ၲ'0}���Q�$X���&��j�A�0Q����,�r9Xq�ȓ{��*��Q�"$�3�]���ȓ�~I;$��D2�В2�U�s�����*���D�w#r��	8yŤ��A��۳Oն���J���2B�j�ȓ5,X��V͈�i��H���R+#K��ȓ�j��lE�xn��K��}��4��3�( ����p�Z�Qb@��M�`<PlQ��4[0J�$�)��S�? �A����(\Pe�ʢf�0
"O^��q�7x#��i$��Ge8�ː"O��S*�(g��}"���&S�٪�"O�l�7T�o��`�4)F�$���'�X��m�0��H*��G�x�N���'�TdR�f	�#�i�MH�wb6���'���cd͑v<��G�y����'��h���$Z�����[T�K�'���y�g���^��WƂ$Z� �'��|��)+D4�A��M��͒�'��Ւ��	+<�HD��+��n����]�.����=.��钂�0:HH�� �,I�����$M95^�R�4��ȓ
�b���P�C�r ���?�6 �ȓ%<W]�z?A�^ZH����"O�}H�k5^���Y%"J�� 81"Ot�'�Y�6�� ��uTlq"O�UZ��Q�!��/��"&��"O����fGv"��3SmS�ZդHxG"O������U��iLN9K�"Ѐ�"Otlb'(�-p���+]3��4�"OX�Yu�Y0V�j(�R�/RӶ�BR"O<�:�Hԯ@=,�z7�Z�r�%"O�ѓ���Z��d�v�<�n!�%"O���e-�A���6#� ���"OȐ��hV�#�8`*�Aˎ.]s�"O�Ր4#��Nx���W���f�hs"O<���U�m����Q��"o����"O��K �!`H��q��D�@�f*O���܎M�hp�S�֙M��Q	�'��!�f�#&pz�ؕ��8A�t��'�"��q�H;�r��P�C����'-jV�G��_�2j��ö�yB�����Y�/�$2J�*��O��yR�גf@P���
��e��D!�yr�ȯt�XC�ဟ`Z (�r�V�y�b�8�$P��T��<��ǵ�y���0
>�q����J'FH�!���yb�6^�v�{��K�������&�y���4R��9to�3A<~$���I�y����J�(�9TA�D@�<�y��k�D�3�ں[�쬉��N��y�.�"��I��1�n@k"�Պ�yb�G?D~�B�CN	�@ڴ��y��r�f�;�e�9���!Ň>�y2F�=Ba�4�RM��~�f	�����y��� -ʉB�o����Fl��y����ZH�*���0k^��F����y��	��т)��c%R-вH��y�-'uh/ h�J`��$@ �ȓ>1>BA*�2���J�g�[���l�� cBlؙ?�l2�c��{��u��w�a:�
�<dKƸ§�;D��}�ȓo�vH�caFo�tn�!%��h�ȓC�L�4�W�?`��Z��L 'Dة����`���_8��H� v�V܇ȓw:��UB�M�9��dΦ't�e�ʓ<��o]�8����`Pj5�C�	&Q���j6&L�4�H;f��O�C�ɲ(�Ը�+�� r�O�|8�C�	��5Bpo�g,l,�Bc���vC�ɴm�A�#�R}P�d	�b�0C��:8�ċ���0���I��MN:B�I%.Z��rO[��z�Ç9�ZC�)� ��������eN+`'�Ui�"O�=��DW�.	�5��  $�"OZm��D�ie��L�%fģ6"O�(��`�9m�a��k�(l���b"OE�#m�h��lB�jj�X�"O,�94EQ�����Q��%*�)�"O �`qBT�j	�shKl%`lr�"On�#K3��iq'�U��=��"Ol�!%�N��&��c A�2i��"O��QHG�kF�ʗaC�ٔ���"O\Ě#G�P
ތ���1}�ĵ c*O\�LφjϦȶeP5E�Fxa�'�.qP�,�_A>�q�MC�1��'%�5�G_`�Jq[���Je� ��'}�4�e�I��������fpX�'n0;B-�#�X�yÌ� �����'������SGPIa"hB-`k�'���c���.+8����A�]'bAz�'�@�R��*_����j��k�'��E�2G�g�K\����N�c�<�D�@� J�ԩ��v���!�UJ�<��,�    ��     �  `  �  �+  �6  �>  �K  �T  �Z  'a  lg  �m  �s  4z  u�  ��  ��  ?�  ��  ş  �  J�  ��  Ҹ  @�  ��  -�  �  �  ]�  ��  z�  � �  a �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P���G{��O�^����0k��	S���$5&bP��'��Ma��/l��ث���*%�u��'��T9@*�'��'/R�!�BI��'u~,3��E�*V����o�&.�PS�'w܌3n��l��2�,��HLj
�'e�踵D��o��aQQ�n�`
�'�:����F�P�z��Xk�Lix��$@�O�lm�d��PF�$���Re�nh��'��	D!^6d`^A��$�)Z�d���'P9k�س����źV�����'�h�ڷ��|ƺ�UMH�N沙��'���sb���8�Dm��m��Ds�T�����L�@�Q�bn�T2B��>�qO,��d�*f/04��BGj+ri���  ѡ�iӺ��F�¨C�@jRˉ^�]�s"O@�Ȅ��� `H��ԫ'M��3��'�,�<	R���X!�hq$��;A�,�ځ��R�<�G�[��8ף״o�|�I��V�ɗi�����>r�a0�C!ߦɚ�@J�
�lC�	֦-��8�4̻O��X���aP�6D�t��X��d��2�@�.$����I5|ON�'V�� pY`�� / Hu��D�U?�ȠE"O6�zS�S M��E�7�:h�X����%�S�ə2��=� Lؖ5�`%� L&o!��[2 zʡð��6:�<`��Ͷe���>�	�=k,�f��D9|-�G�
���H�'�A�U.C�sW��X��ާh"H�{2�'����b�Q� њ�鐠���i�J>���?�Ži��\�wB?� Ia����5d ��'w,�*4a@�^$Z��2L���-�L>�2 �Sܧ9���7a]RE^��o�9j��-���MC�MY"E���Fb�R�f�1���]y"�a��(��������j����F,{�HM��y2,+���c�#a�\��2.��y⠜�}� h�M�Z���r�۰��<���I�qԠ(��N�i����>o+!��ΛR3�u�c��[���̈́�$m�'�1O�}��qp��&��p�,�@�*�W�<�0�/�� b�2T�䘚ËQO��0=�mG����
��.5�|��gTd�'XQ?A]x ��5�Z���Eh<9��
,n@*���g�����#Nv}R�)�ߦ�z�ȍ�ua�W��2U;�A3D���˒]�0MQ��צ#�00�/D�((E��+�B��E��V��#t".D�L�CC��5�&�`��U/(B!�'SM*= P�m�,!�SC/4�!��# J��aTgI�~��0"� U����)�'%�R$Z� ��P��M�<���'YЅa�Y�|��\�ua��K@&E�H�L���7]ҜP�%~Y��Ր7 F����@?q�`K `؄\��L� kt�	�Bf�h�<�G�#Q�Tx�N��% :��H~�<Y�G[2.�:<�dAs�ܱ�]z�<�a�B�K?�U��!M+
(I�g�ty2E���OQ>�W�ɿJ��MQTL��SB��3�F9D���L��$y� )&-J�L�~�+��+��w؞L1�Ě	�D�����H`4s�)�.$uQ���\��k��y��W�V ���G"Ox �u�_���eH���GUVi�Z��lG~R2OHc?�ɡ
��@�bg�#��@�����\����ȓw���
dNT7�*�Q��Hz{X�'��~"'��;/|��[���(F��4�y@#Y+��S�16�(E,Ƒ!>�'�a|B�T!&.E+��I#_?�<���ز��I[�'[񟰉2'n�.�d=�rjN�{�pT��"O�E ��;���(c) *<:L
G�d|�6�=�O�$<k��	s(G��:'p0�'Z�AN2:"R$2�'!���y�'`5�!C�U>��)� N�jEB�!�'0y#�<K.��+ڧi�`���'�a���o|!�U�P�:�>`p�ǔ!�Px�c	>'q�y�UJ�C`�m鑠ַa6�MB�'j�(��Q�1���3�Iǐi=��b	�'
Z��𢈘��M
�.C!g�ܰϓ�O�:](yE�+XQ����L�b��'3��Gy� Gt��`+�)H9ZX;�?^!��U.i�P�Z0-ќuQL�ɓ��1U!�䉊a��5Qv�|"���)2Y!�ę83�RQB�IT�o�!��
'?!��ę+!�Q�d��"����1�B-A1O��=�|�&�N%��Y�S��	 W�M�<�C�G�|�P���P)1#HA�F�<�vGO�Z��-Y5�L�X2rԳc��E�<���Yt����G�~��T��]B�<� �xqe��^K��H�Q 5�^Y�|�0O���=i�y�NK-5��s&�g9yK�nю�yrO������	S4p�xY��Y��M�}��OZ�=I �m���Wo\U� �m��y�C�99��2��]��2�)Z�y�A	�pE��J�T3>/�����$�yҀՔ*�(��o=b�����y��J�G��q�EV%cKu�dj
�y�/<x�txZ ��8kߔ�����yR���t_&��� �P�؍�􂎅�O����wH"c�ݢH�x����&e!�Dװ���E/ħLu���2�V�^b<C�9$/��[u
V�%m��iR���.�C�	�?���)@	�-9��+�K�#�dB䉽n�4BNZO!�Y��ݞX<6M=��h��D%A�b�[�@ N��`Ye�5
d!��ٛa�Č"��O�JC8�#Kay�I�	D-�Bb�:yav�zá7 ���(ʓtI2�%�F��x�&[WG�$��z^�H��"S�2���Ao?dy����-�D&�~h����JQ^��=I�K!LO2U�פ��UŐ
T�(�r�i�ў�S��(O
=�`B�zg��Ya�¶b��
�'�T9������`��\�=����'8�>�	>n�e���p���#R�*C�	.)~Xez�#О>��}@w�S�58�E�հ?��郙S�r�[d��20G��"�b�'�\C�I[S����@(�8$�.HPf0}��'�F@X��G�I�3�U�y���'��(�T�4�\�p��ЋvFR��
�'�J%҂��v����bQ7e���
�'�0h)V(D)"�X�#�Ƌo}~qI	�'����_c3��J���3��c�'Ն3AA�t�l�Ȑ�ϣA⨹�'v�2�Mh��<� ΀�n.��'�z�PGY�u���� �˂H��H��'נ9RbIѫP`�Q@�ׅ6��+�'���0��(8��Q�g�.�عr�'�����\.v�}xRG+!P��'r.��*Ώ&��\�֩�&�X�'���ÒB��h���&�Kݔj�'$��9��܏�(��n�O��X�'2&Y(@�Q;nt"&��Ff"���'�j��b$�W0�L�ū�P���'eȨk�5��j��@��XR�'�n�Á��?&z@�qQ�ج0�6���'�LM� �G,u���!�ܶz�(=�
�'[ډJ�,�&���x�I1	[�08
�'�>ya����_�
�DI/1zHA	�'4�4b��#y�M����$%3�(��'8hHPhT="rMrQ�q�-0�'߆)�o()��ժ�@��b���'�bx ����6�΄�3��V@�	�'Ϊ���h�|O�@1�b�Xn�9:�'<6=)1'��f�Ni�c��U��$1�'zf*��E�� �����#ިy�'�@a��M_�o�i�L�	hR�<)�'��]:�"B
 �d�5��gsNT��'l�����\�Tr8�s��CZ�m�
�' \��&�Ĝ����QvD�j
�'��"Ԅ]�.�$�V�P�Q"���
�'(�x82훷@?T��b��H��}�	�'Y8;p�,4�zlq��TB�h	�'�zY(vD�6~�ə��ǩC������ ���sD�0�@Y���<l\r"O��b���%p�`�2V��QWt��p"O<ɲA T|�����Q/ n���U"Ol�#6��8��{P�:5c:|j�"O>I�g��0=��K�gJ�<U^0�C�',"�'U�'��R>e�Iş0�� X4���Ԃ��IxU���}�IٟX�	ҟ`�	柈�IџX��џh��?z����5e��(� ��p������,��ʟ\��ݟD�����ʟ��I;Mъ�R"�	{n(�p ��p��	�����˟��	П�I̟ �	şX�	����b�
I"k��A�ʞ������@�	ޟ��Iǟ���埰��Пp�ɶ�� �7��<��I� �#����������˟��	͟�������	�x����B�ҡ̐)]7�	�d�-5P�������Iϟ��	̟�����柠�	7_�,�Z3`B
7��G�Ӵe���I�D����l������ş �	���I"Hy�w�2K�� � �ܕ$lb`�I؟����H�������ϟ��IןH�ɛ=Fր)B���De�aeΒt3�U��ߟ��П8������	ҟ<�IП|�IF$�@㟼�(�pBhT�>�1���<�	Ɵ ���<�	�T����	!DT�=#�R< ���'���	�����ٟ,���T������	������;D��F�#1lySb�Ԡ��	���I�������̟�Yڴ�?!�=`8Q�ud�Cؼ{M�f
e�V�h�Iky���O��n�qu���Ƈ�#d  k'ƾwpw�9?�'�i��O��O�7M�NC��1��[�G!�L��a�*���m�����n�)�4�x~�=K�)�>W�OjAH�H8lu��(-�	AaY�y�'@�[�O�t�P��+�<襫��V=j�`��q��2�S=�M�;7�d=1�&Qp��)Cƈ=�l�s��'m�V?O��S�3012��ek|�tR/��l�Vl���µ4!�lIdy���ւ��H�Lk#�V�����'�b��HO�����*��0��'��s�I��M���N����z���<	q�I�k��y+��n�<A��Mۙ'���3<9rerc	F#E��Q���Uj��K��Q�"�ΚP���|@c��R��{���腆K�������
���)OTʓ�?E��'ܖ8If�W��
�0�\'[���1�'�7MP*d��9�Mc��Oҝ �ΫM��$�r�c�(|��'vB�ir�%@KН�O�t!��L�*��@J�vh�\��Δy&(�ꂪ-ex��=ͧ��"���!&e�E�L�8A���R�@�k�	<�MC���M̓��O��}ۑiُB8�p���� fJ֝�,�<����M��'��OZ���'=��3qdա
�q2▗ �J�Y��V-\�2�O��W�+e�f5��	��I(��D�*R
x�D�L��cd �B����<A+OĒO��o.:_��� m��� H���ɚ3d��m+z扇�M������|��?��4�?��F,|���mF�w��ݓ�+K�^N�#e���<����� ��9~���'�Tgy��b�M���ЪrD(��٢�g���ImyBW�"~"�$F`4=ѫ�/G�p�ŗK̓:x���3��$������wy�o&IO�!�ʿ.) ]�GX9��ļ<	ܴl����'��y�)�?�yB�'� ���L�I��9��c�'_2TK'�E�H��L2F+_�>ў�Wy��'_��*��jp@"Ǣ0���8��b��&�@�ش7Ub��<�)�D9sV�رN�J]C�hE�$���)���|�,O���yӢ�f���?�J �_4
�Ҍ#�BP�d�Aႈ[������eB�p����&�c���S�k��.�jt�	$:��� ����8��pB2�>Lm
@��V�O���*����`�F|��޴�~}�t+h8>��d ���O���]�dݸ�-F�]�v9�R	�9`%u҃T�<Ϙ�9Lx�C/ۚ#���I �R�q�,�3�@��6�ݙR��2��DI�'t����)ր�2��i�T��]��������N�% �^a�$I޸|��x��쏅!�(�@kW�x�8KD� �%��ّ�O<4Ɋ}q�+��zI8b`V� \�+&cQ�[\h�I<���?�������O��d��V��p�N�.���Ƅ��T�H�ou�'�R�';2W���mS�M���r�{1���=�� �Ѡ0e�Q�'���'g�\�8��ƟP��&�~jv�)}
�R�ǱpItD���p}��'+b�'��	*l�tP#N|r@�I308��P�0Lhi	B%K����'�'��	C��b?]��拣$2&l���E�cmt�m�z�$�O�ʓp�`�)ĕ���'��\c���%����	�7t.^�i�4���O��d�*>��s�H4*TŌN�`%:@�3=�~u %�i��	-�ݲ�4{b�S�0�ӗ��$�o�J��`FH7A������[a���'�+պ��)b�g�Ij9�r�K��f�q�#�AT�7�� a>|m���	ן����?��	�T�I�G�lk�m�R��1��pf̩�4*�d�����|
O~J�I�r����{�P�0န�0��׽i��'-Rf�'	�7��O���O�$�O�	ŊIi�!īw�u��I"����'/�	�]�h�)���?a���f�@tNOI��@*��(@���i�b-��Oݲ7-�O(�$�On��Yv���Ofؘ��U|����̛�'��uZ�S��#h�4��ʟ(����	S�t%W�|��Hs�kY;IW>������
�T���l�z�$�OD���OR��O^�韘�� ��(��ɞ���cg��5њٳ%��<1��?���?���?y�6����iV{g�,�퉰+�% N�=�4!s�F�d�O����O$���<��uָΧm�̸�FFZ�AD�2���*�^ȂT_���I�H�I�|�ɩn�h9A�4�?���kd�8�FQw�QE*���p�B�i<�'�_���ɍW�x�S��x���O��dk�dɡL����� �"ai�'����I̟,�	�^�p�4�?����?���d-B=YlMV*��ੌ$v�f����i�2U��ϓ}�,�ST��?7[�pt�D��y�>�y���`}���'��n�4Kx7��O����OT�i��
� ��=3t(�Xƺ��Ge��L,�'2#�1Jr�'��i>)��v����՟^XX�YTʌ,"��1�iozр�fkӚ���ON�d�"a�'D剂=P��3,�;�d�s�;N��[�49S��Γ�?y/O��?��	??���4��o[����d��X6tu�ݴ�?��?�'R�r���Byr�'�� YX��ש�?8J:E��Eڑ-��v�'��	)�~�)J��?	��YX�U)��B�x��m��C�CNv�@r�i�R��j
v6��O|���O��D�N��O�l(E�Ÿ��$�qŀU�by8�[���+h���'���'b��'�LҢ�Tu9��L� �{��1��A�P$u�����O(���O���O
����j�@�=)� Lh�i� r�8�d�Řd��Eyr�'[��'��'���Hy��IU��je����&C?h�$��,��A��ڟ�����`��{y��'[ԁ�O�Xha��~؀�	��2cI����Ӟ�$�O��$�O2��O�s��yӐ�$�O���v/©!�H4�D!;^��P�VѦ��	͟���jy�'�����D��_hf!ʧ��=~�x����=4'���'���'<b��4���i�b�'7"�O��l�H��� �o��1c�'e��d�<���/j��'���|n�w����e*��\�}j�/�&HY�7m�ON��"Dho����럄���?�Ik ��Ԁ܍x���C�Ŏ31��Ol����Y>v���O��$��#?�i'���;����C�2Z�����M�7�L:��F�'�r�'����OU��'.bMD�	YD�0g������E��7m�3$����=�4���(l&�ɹa)΋7��[v�ںk)V�m�������DR�Ĵ�M����?y��?�Ӻ#�I��{'J��l�0��0���Fئ���iy2�]2�yʟT�$�O��d�D����V�,�:q����5Yw>qm�����o[��M+���?���?��]?Y��_����!EN�N蚹��]1+$=�'��Y�yr�'���'�2�'Z�ț��Y��
&�ǹ=�x�J5�G>��7��O�D�O��Vs��_���87����P�BP����>T~fq��w�T�IΟ������	E��-M6^4v6��w�j�J���J�.�ʜ�.�N�l�П����������'�b _-����'~��k�+[%NN���._�'��7��O
�$�O����t��	��I�7��O���N>���;E�T�,�b z)�v���n����	̟x�'��BZ��dU��q�l�1)���PKLS������7b38��	蟠��͟+@i���M���?�����&��M�l�0\�$oD
;�\��4�?Q(OP���0��	!�4����6\}&L�C�8a�
�È��M���?�7��`��'���'����O@R��IΝ@3�M�\�j]���ˉ3 ��?��FI;�?1H>�'���2n���*A���4$�&7�6�U-dܨl�Ɵ,��ϟ����?i�I���I": J��#�G�Q~�,�Ճ#�,[�4nt �������	(�i��,ŉ�a
K��Xe��<��Ax���Y����<�	�h�!�ݴ�?a��?I��?��#�]�ք��!ЂnYO�,�nZ��X�'F�`����I�O��d�O�]	��D Y�a
�>ڡ� �����	��RA��4�?1���?)� ��S~?9���8�v�x���B����q)Ss}b��9�y��'��'���'\�S��b��^y�H��ʒ	�00Aύ��M3��?y���?Q�U?m�'l��N�!��K+>:쨐F�8���O~���O����Oʓ:좽��1��H����
s��q�@�(#�ֹ��R�L��ßX%�H��ß�҄�t�PIM�����¦أRQ�mˇ����O`���O����);c���ŷt��Ա�;it���Ǥs�N7��O|�O,���O��� 0O��'�j% ��ȓf�X���'H
�F} �4�?����Ā�
�%>����?e �O�$`��]��"��C�E!���:�ē�?���2P���S�cm)8�&L6b� ����|QUl�dy���O$�6�[E�$�'u���-?y�U� 9��3�!PZj��T�æ��	ӟ���-�S�'(�f�"�탑J��Ĭ�
R`�n�
81�!+ڴ�?a��?��'F�'�rÖ�9Z���vȄ�Gg��&�_>fB7�J���"|��#C.AA#e� ,A��0S��i��'#"��ePOB�d�O�� )L��a�!��)�a�D�[�'��b���F��f��埤����4iB�I'i����aI�1�0"
�M��{jI���Op�Ok,�^�1�G��*���8b嗦a�	�f�6P�IPy��'Cr�'@�I�� ��
;��:��N��� RR�0���?	���䓾?�7e�Dr���a�dijsɑ{#N�b�Ù����?)���?.O�AP��|"լ,\����e�(Xs� ���M}�'�|�'��f^wE��=N�����i�	�n�B��2�p��?��?�-OD�X�M�S��4h�bҲ� %*T�Ȍh�(ٴ�?�N>A��?I�i��<�I�� ��zG��<l���3��3aa��Q��i�2�'�2�'qX��u�pӺ���O������d#��S�� e(���D�G)�u�	֟��	3Ǣl�IY�i>i3�(�;ft�(��K P���@�4��tJAi��p��"N���H|�>����� �+�U"��<Y&��9l!��)R�X(F,T���Ё���&hf���j�d��q�p�=���Ԛ9p�� 'ΐ� ��p�X#�@Y���8�0 ��J �`�H�~�h0�?"3x�`��R����;��݄߀@Cs A,$R����M5H����k
1*�.�˦�O=��\��j^#:�^-YC�M%O��)������?)���?������$�O��k6f�z �5n[x)LIB��P6����ߺk�h=����f���.@���ÙE��Kk�\�T��\�H�� 8W(ġ'���Z&I�?�=�b�@�(�@� h`�x��\?	�G���DJ۴D����G���;_2ڠkc���G��#�@���yr�Z�"D��M}���b�hM��A������<11H�-ԛ�'}1���`��7$L��46�b�'i��'��
��'+�0�4$�!OM� ��Ϝ 216�!��"H��]yV'
�(� ����><OD�襡�8���R�
�
��,97+C�Gf�Е+]�0�b�8C�$<Oh�Ѕ�'�R�g���S1܈8'�c��׳6'��$&��<���ʝS�x�3�)ɭR�(��Da�<!�c�z�X"B�3c����!�[�<��iJ�Y��r�B��D�O��'_F���_
'g��6�9"`�#IΨ�?���?A�曆�BP��S
@kF��	V��t��u J�6q����zQ�x���Z=��!�v �y��ѡ�l�	Ja�����OYX����m�V u��-Q�,���O�n���MK����ja��#���@`�y��ɰ?*��D-�)��<�wo�\%�l�%f��?��m��L�G� �K<-
fIk��a`$��m\C�ɿ�X�r�����n��������'���O�B���A�V, p��vD� �|,S	L�z�EBRA�6X)��T>U�|�	�v`� -?ݼm{%��<m-�!0[H�rc��6�,�r��W��?E��\����0	,T[7�ǊW����EN��?a�����O>��7��yP��΍� b��>?�d�O����W�E0XYRr��>XO2���K�=6-�4@��4�x�$ū?gVx+�ī���S$�OZ�d`�l�Cm�H��O���O����?���>���@V]�:5ˢi�b=Z����Ӱ	F���f����|) �#�AF{B-��cF��^5
�(�"E�B��,25���*՛#�֘4JRa��hOLU[4� �+�vt��#j�;V�O�TI��'�"�|��'�"V�L�d@�'�� ��'�-�"*9D�$[P�Z��
�AgIC(b%�ш����HO��	�Ohʓ �n<㦰i�֨���$,(��#��a�di��'g�',"D��f���' �C�#U)�8j����8��БG�X���`X+c_8���O�w����P�Y=x,��-�N��\���SQc  !0+C'h��hkC��'?����N;��`�M�O���ܸu�����g�8cl�z�kY+`��o�����'���?y�pCZ:>� �K/O�p5j��1D��3�
Wn�"b+=t	2lp�Գ�4OE�W�$S3������O��'�e��*���HI�L�*�1�!#�?I��?I���Zm�}Ö�˳��}r����Ʉ7XQv4�@�%�
	;2��08�Q�@����*H��`B	�����&>A�T@�9�$S�.[�Z��:�u(�A�	�������O;�B�蛮H� �����:�hC�'��O?�	�i�|��!�,��8�t+V�+���$VX��V�t-���#B�᫡(� \���ɇr� ��4�?���)������O��Ǌt]4���EX�Z��L#�_�v�^��$����<��O�ɢ��5���k�$6�r�[<#.2dP�h�o�|����O?��A�8��������A��Ȍ�q��J�#�OL��$?�{��?i�ݽ*����Q *���J��<���>	`��+>��@'Z;R�L �`�m�'��#=�O��Zw�X/k-F����÷^���!�'b�ڣ�м�5�'�r�'���c�!�I���ɁB	k�Ѱ���8G��5b	�?�$�Ԧ�c��L�D����g�'�j��ȁ $Hj2�%�75�&�#��O��!��V: J�z	\������'2�!�Ră|AraBD ����ٔ$B+3lO����ׂY_���_6�.<�d"Ot�GL��Q�y�A$�� ���ை`�����|���Q��6-ܛ8)�Tk�n�7-AB�K�f�6�����O��$�O�z���O"��r>�"�`ݵW��P�Uz�P�QoD�)ڄ�$e�#8 ���D����A�"�3��6�H�^�.i��"W8N����'��qR��?ye@ԻP��)���?z	d������?I������IH�a��8���g�@��2�	�>f!�Ĉ
5Ep�0�RRŮ(���M)pU���p}�|rd8�g�? �`�F���h�h�$�>X<b�"Of= .ہs���@�S�qi�� "O<$0�͚C�  c�8(MJ��T"O�]���Pfz�]jE�� T����"O�d+��K�J�z�C
@},�p"OT�s	�a#(�Ĵ"x�p��"O(�"��W���{S!�"nlRYR"O���&V	�T�G�VR���"O	R얦֦X!�hWzP��i�"O�,K#SG���;7�*G�B(#�"O���� !d��ߑ綄Ӣ"OR � VS�@x�MF�hE8a"O
-�D��	�RI��E�c�Ĥ R"O����	# SX����	!�Th`"OB\�D�ȴH?p���g���{U"O��Z֢V�*֢@�7�V�⁩�"O���^�>º��%;
�ȃ�"Ou�Q�wܽ�p�M4i|P�"O�q�$Bv8Τi�ֺB��4j�"O��0Sc�(c�r���C�����"O<x*�,^be+!e\�mܬ�p"O�0�� ׅNJJ���e���D"ODh1����X�$����V�v��7"O�2��B?T�t)��Y5T�2��"OD,�c���T��e���>{�Bh�"O��@�d�x��`seL�z�Fub�"O��3EN;@��P�9h�X�Z"On{WD@�(�Y�B�w�q�"O�a��lT�5������ۦ��{"O�yB扐z:9 ��� R"=�G"O�`��6S����W?�k`"O��ڥΓ$f�H�ѷ�ObX����'�6m��E��'���т@��F)��E�&�"�s
�')��1d�^���%�r)�5�EN~G��* 2vc*��Ӿq(33��u�<!kPlF�N��B�I'<]fQ�b���F��(����&��u�O<IUhO=m���|�<�T�h��i�.^D������[<�Pt�.J��ԣo�@��C�'b�%I3�R���?���	3><5�s�X�>1p�ruk�N�'L��:���"U�����{�G_4=���L.�Z�bu�˸cv���I#1��C"\�;N�hkdl��D����a���� ]	�'���&�0��,�z)��o��9$���Sf�^�<i���0q�vd:4�0H�F���͘��7��n?��j�?
)�,�Ĉ;�B��e����	�S?6xP���(H��)��;LO<)Q�`�8��$f�)
U�^�9nzmh,�g+j-��~�Ě�OV��e!��%>�vE��2�S�>���P�R��`%����@��a��N�!����'V�v�I��V;bo!)"��ʒ`a�d�`�n�!�r� +$��v�Hݨ�䘚\h�-������ɭ
Ύ�������g���>A�F�l
��!�.(ld�y&�Y]h<Qt��^d�Dm�OcLy�c�7���i��P�>���� �O�M{�k�]��D�����z'`��JDb C��0=��Ib��I�_�
ًA$4�8���!��]��0�^��u8%ҲC͓X���#� �u��Ě-3P�Sᤂ�h�{t�	_�1Oh�yp�-����*g���ش�yÊT�1��J׀DX�o��k�2삖ɑ1S�8Q�pX�u|a|Ҹz�b10�aT1�"�� jV5� ���'�F�'#���dKF�1O�nM<6Q�g�H�)Y4��XzC�'���Yw���K�,����'t5�0 �O�X�1,�W��vB.�s�>����*|̭	bDǒ=P}����7��M�HXo���y����o��I0c��%+�K &@�1�͛�V�N�#�$?a0H�M-ȜlZ:PI����0�O��,�s�tK��V]����|��F(���Ƨ}Ӗ���k��.i�'��-qUG��ܐ��ȟ:ff4��U�3������!����I�.��"���d��#^�j�|r��[G>�l�/Y��Ŋ�Ӽ#��� AE���gD���B.YSH<14��3ʲTȣ��s�I��׹~�ax��R>-��6ϟ�T�|��3��sJ� tmR��\R����ECvF�R��'�R���U?�F�R�I�U>f��W��8�\A��̸��q��X�qe��<	�I�O�Ty3������O̲�4���Q���$)Ę��%��E��u�<��-���t0���>�h�B�J�Y?���M��B�m�(ַ&Pr�qgNJ}Bg 1�d��{�RAp�.�HO�*7`� UD���gL�i/�%�cl��2��VMĘ	��5����5�4%��U��*0e^��6j\fx��U�
�ʨ W�'�Ƶ�Wf�)m<��3b�B�0� Ór+1OT��3���:�d�a�A�%Cd�3�� ,l���剆��c@%A��Uo��wY���Θ�D�Qj#�	�9;��
�O]��>Ov��0mm��I�'�ᛷ#O�َ6MF1r.�����t��c���2g�'i�4x�Y%N �*$N�%�"y�}�MY1�P%C/X�|U��#�9��Đ
Y�x��^�ΠӢ���������F=��"��ÙR��u��8>]�Xb�+�b<�+3O�"?�1\Uj0X��]4CV�驵I�d���Q��U��D1���!E3n��B`�(gV�p�	ǓTM �k�8�
����G����뗳d3ʓ�ɶgH�p���'If9"�/K�-O�	�򠄗:�>Y��f��H�]#�׹d���O<�B���`a�eVF!#۴?8��"�'��<)��N��F0۶���ys�A�~�	{����b��=������(&[v6��'VLL�1���~����P�^��d(�߶B�JDJD�==�T�ԁX�"��l)4�T�t�������e��@"�kX�MT��r�_8#iv,R"C$b8�$��LŘn���sf� !:�a`cI�H�D����~���-��9;����}�9��Y.b- Ӗጓ#�a~rnI�3ل�p��W�=E6���"ڿ	���yM�cjԚ�d��;%��� ����G�|��*ʟI��;��O�E�:�
Q�Q�@y�S蜠6�azbF�! <��I;>�z,��Y)JV�x��� Gʾ-Q�(R<D����ܴgF�SdHص!e�@Ǔ"��un�\&�@��~��nU󇏻M���3�N���'4��7�^䟼S�Aq������x��e���9QKU���!L�����\5pq�-3�P��8��@˹Jy�T�͂q�tS4�Ʌo��4������)�`�\�}��T�W��536����]�OW��+$)O'z�>}s�`B���^�����l�����K�<T|8��j(lPâ�'�<Y)T�G/-���ӇiK3{3�-��̒�F�jԒ�y���#ڠě�����O��x�V�8^V<���3`����!�Ӣ6�����1&@"|	%KVǦE�F��U�2�YUdQz��� ���Y�-�M��/��� �� �</�n݊fr�I���
C41
1�ۧ,����A���K����?)��������R�! �7M��sxRh2ڴP�j( ��D|7�)(5d�,LטȰ�o��-3����ƝVK���.ou�Y�6�K�>�l�k�l�_��t��0d��i�U%ݫ2 ]1�ML�qN~	A�Ŏ��Ҽ(��g�TT[g� R�H��-̉v�7=�����I��8N� �+C7��=����7\�څ�(��>1P�-g�h86�{ ��2� 3�8�3􊇑e~���BY.GX q��|r6d�m��2sE(�@,6�*��"+Cv�r����)-����DF�vl�䪁P��M[�ݓ
���&��y�=5�W�sD\{�X�zk��5�فKl4zAŷ#)��3.��S��I�7�T}9�'�\xb�t&R���=�8bM<)"�:��4r��aӞ��+���M�ぇ=Ō�0`"ѱip���!m[=�BgeČn�؆K-ZF�QK� 4�R�F�-��Ր��$7KԜ�7�ҩY��N&c�p�`H�l�00s�&������J
^��{b�Ƅ7J����\c�DHc�Lz�`Ag_�Ƭ��C�$a�f ʠ�*�Okl�)h�X!�)�I�衈���C,�!� ��҂Q�t��,c�zDb�|"����j�i��`��9zU�vCָ���'�z6햌1��+�A�0B���C[Z� !��^&0� �f�O0�G�*�~� � �vg浙�R,>d� �޴X�A���ܜv�x@P����~^�<�"�D�,Z��Pw��O�mD@�9V���_M����-��E�� ��GM�	�UD̓)t����{���i'�X�A%~�����"��6
��4�СU�U��+@ĉ2i�&����4N�a���p(Q�h&�cƦ��N�pYd�¬$ς�ʴa�:bd��F	�e���Y�\)��\���(؁$$������Ű"ʄ�ub;�O��@7*Z.~��*���)��0qJ P�2��c�Ѫv骨��37������u1-�1bf�)�fr�a��d.E��x�q
U&',����'��:�"�3Vt�ą�B2�T��4�T1��"?o�\�($'F�}2`�qM�J%ѳ�̔�F�ru�#9PW��P* +OL�j��U�B8��7��4��C0�U8$E�'"�A4�Ed�\D* Y��!��-eR jd"SM.��6D��	a���@�.}�ʦ��oKd(ٔ.�J>�0ԯA�,�>��L6ғ��`��OƯ��Y e�@�MkT �~d˓g�-r��X�P����u��4�P�9��r���Z�VKR�j#�^~Gp���G�,&���k�,�v�����ƛH $uSr��,����&N-�j��FZ'�yB��?y����)�Y�xR�]PF�=��K�2���"��K�PX�ד=#��&%V¤�7i�1����^��D�#��	�px���jh� �w�|���*��!�s^y�ΝEw�7�Tsz��B0��l��Dy筂 ?�O�x�$د����'X����Cuyb/�h�Th�n�)2������_����R�4L�30�'Ubm��R�4����Z �dF�r��Y%y�b���	�E2xpBbl@�yB!V/^^����?Y֤��?��O��!Nq�P�f��(5�^1ra��S5�O��V�i�DW���lHM��@�!�\���M�d�Db�7���|֧y��ڐ�J�
�Y�p@���0>y���C�q�S�? 
X��D�!i̸�17�Mmm*�貤�\��bZ�U��'8�f@
n�̌`�Oݖ���3�6����a��=&쟐x��"<GF7�l�'O���O�-!���4��8sf��)|�����W����#�N�1P�6}u���Ee*ғE��a�)O?$�,ٶHC�*�h [�g����'�
T[C(?A�۲-��O��pQfQ=Ŝ}C���
��u��,�W��W��W������tz��1�. ��	�#ΡwW8YK�'?�bW�o�q�{?A��<�s��i�Ҵq��)��	Yl��7O����g�O����h[78��Y>]�"	�@�\8(�H0$jˁ_�����4A��	M	����M��O��v���C4�L�ʞ��׊��9T��(�j�z~2�	)�]�U&�05���J�s�L<i2�^Ҷ�t�_�j1�m�&G}}��x"O�f��%�ɂ�L�3�57��S�ʶh��-��I�x�0XqG�)q�m��}��MK�4���A�'d��!H��e�4�8UIځ9a�zF.�Z؞�<�y%���;y�Ƌn�������'z/D�$�b��:�rd tg>����վ%_6����><��8�C�݋=˾m U�E�L7 ���'�A�Όi��S�hK����O�	`pn\;��I�ɇQ����$t��Lh���M��г���dKd� G�DC�e�R�!�oRD�@�jf$��5��'b�Cej��
�]:�$��K����OK.��'1����*�UFxB���V�wc�
f�j�t��=*T�iuhU�0�֭bҤV���<�K�Tj�iX�Q�$ Vo���%H\�&�$��&JXim�pB0���$pq6L*�'�JYk0�Ή^�ErD���;��˅ď��<���\U��x��?W�&�;�c�Xh:�S�i���R��	�ax�HÁ�L�R�O���*2C�B�<|��B��=��5dM�B�d�)M<i,غ$��W∧/rV	���@Y�Ej�p䯕����Bp�lD�'��h1��:FY��@�4C��0���yDJ|����. ��&��-d�P�C��'/L ����b؞	���f����J��,�h�g�X��en�	(�{Zc`��S掍y�8<�$\���/��<q��)�S�o���Q�ٔ{"�i��ĉ4�T�d�&��<i��ԩtU�`�,A�L{�� O�>��S�P6=�V����IQ�XثQ�-h�})W��;l�x�D�P'o&&��mj�YE�Sn�*��[A�i��'#�l��O8�̓\ļ���ҡ���EK�.IsȘ�'�D��%���3���� ��T8���?%���b��_�5LM���U�~p��I��d�'/�ď2ݛ��O�u���I�<�U�D�5F.���MCl�D|�4�ƞa�L�[g�it�h
�?��,x2n�lXp�ڧ��F#���W�̢gcvp˂�i{4U�شba�>�S!�9�'^4 ����P!eo`u�ȓ?�u�bt�1�^#Q`�4�7���t����iD�ɀ�p<I��'NC�����h�Xء��Gk�<�S"M�*ͮdq�D Q���ٷA�e�<	�h�4K>���AlĔ1R����v�<��σ.N��	��J�s+��0��q�<�筍l�6�x��G�_�H��3!�D�<q�Ď�Zwj�ʷ�V�<�@0�1K�e�<!&	ǍR5J�B`�X�EzRt��`�<I�o�c�V�1����<Z �4g�a�<1�,6�: ѷ�m\����e�Z�<�MU7z�b�Լ\ �-�(KL�<)@����hQ0��9�t�dC�K�<����)�!2�c���	a��D�<�S���d�f�!��V� V��|�<�eI(o��1���tV��(Pgr�<�V�i��"��-z���8�di�<��gL�bb��R-K,=,LP�`��d�<Y.�e���"EJ�8�^��v��g�<y�M�� ��Z��өT�����fFg�<	1�8<�\ ��:Z���bb�<�d@��sߊ�ƀL�#��y��VR�<�f��9��9b�Nդ�X��h�<�rlS�x�P��Ң,K�x��e�<I�d��i<�T��;.����j�a�<y7NF�x��ru*_x��C���]�<YTC�"mj��مh��v+�	�#�Y�<�� �2� I�Z%lX��T�<	cB^�;!�Kp�I)P�
��P�<�d�/0��(�Ґv��\��J�N�<� �m)Qǉ�?�4q�3�V�{���)�"Ot){�ĴM��Q�s�݆x���7"O0҆�\9f~xtp�Ir}�ѧ���<� gR,:�0<�O�W�6��5�KP�<�� g7�1B��r��$�/L�<���*
-�&k�	�U	��ZP�<� 'F=t2`�@a��\A��F�<R�ҚTtfd*�m��05�Ů�k�<�b��-����'�G��H����e�<fl��!��iTC�P���0�Xe�<��.P+8+!��ݽ^%*m���\�<a���Xo�Q�Ӕ2־qSr��n�<Y�)�~|�8�ÚQ^�@;qhg�<�E�ٝ��y��@T�Ԛ�J�<qR�ɄP�t4�է��@w���d�
H�<y�P3'��c��(�:�j�J�y�<�A�=�����. X��x
[<�yr�K�츩��ɚh.�����y2��E������جȶ��-�ybAC�: ��ؠ.{�^Ѻǀ��y�["C��A��a	�H ��kLI�y�dI�L��1	�f�F��uS'�yb�֓7�Y��R�B>(]�	_�y�E��%��%Y�ڞC~Qᖂ@�yBn��`ߨu��3:��ئ`^4�y��Z�[��㎅���LX.۩�yR�_�F-j���S? b
���(п�y�Je��D���L�wV�LI��G�yb��:��=9`��!cu�8g���y�a��0�h�tɔ��%���y"c��>�:t(@���L�R��%(��yR	��^���ÅF��R�X�UBA��yl�& � ��*@��0x���yb	�C�F p0�I#'U�]����yr����	�`��1D�a���R��y���[H�y��*8"U���W��y�̮5�DCcķjZ^x�Ca�)�y�l.h��Ad�3\;ԁ:�C�<�횞H:x�`5�� AD&P��"�B�<�5T�&
��aU"��|�������W�<Q"��4�z�O�Z!�0G]W�<!��\bd᳑�1Ӥ0
F�E^�<���O�	D��! ���Hzv����BS�<�'�Y<�|�K��}�VE`��Q�<q�]�@ l�jQ�Qy2�h���O�<�M-eo��񫔍_2Pa ��Xe�<� �� V�P�n��eZB�:��Nc�<y�E�LAL���m�UZ0C���[�<I�ꗿTp� IL�vu�;��YX�<9b��@"���I [1��]�<)�1&	H}��!np��%��Q�<��-�k��ᢃ��1��i@���O�<�=BĶL��	,97��;��a�<Ag��9�.a�)%Y�����G�'�xBO�U�|)�C&,�F|;��O �y�T0,vL���6tx�6C�:�y"j�F��<���օX�|�Iv�Ø�y�	ٟ+ސH"
��ZVd�tKI�y�C'�p�a�׺S�X]9A�K��y�(�{`��F�=��: �\��y"�ژ	�)�([&/θq���y��W�p8RA�����qB�LU��yR�Ѓ���ئ�L}bQ�͇�y�eN�PS~�2I�; X�t�W����y
� �M"V�^�}�hq��L	�m�����"O�L	Fi�B<*E	�m
]�"O��[��η
��U!�N�q���"O"�X���,�^��d�	
.���"O�l�G�M�f����>D� Y�C"O�)PA� D[�l�!=���d"OH ��)s��`���|�h��g�$0�S��K�kN�$��� ��}p�J6S�!򄎉,���r�I^� |�1�F�6n!�$�7�`���_�wn����<2!�D�9�|2�li�-0��"1�D!�S�Ow��9����Xe���`^�HQ	�'���E(Ҫs�:@�*��^L�'6��a����TH�!�:y�\��'G��Qbe�Kʐd����~�v�I
�'����aT�n��v�-P���	�'�D�'ւ#`~�-q���� ��q�<!�@�	j�i.ރ����\m�<���U�6�E"�������%�r�<��
����g���8���
S�<!G#`�d�梌>em��#Xg�<95;!9�*6K9yB`�T@�z�<��@Ūn\<�5KB6q�t��NUb�'��x���T���ӚeG>�	�Ì��y�S<��������-z�-��y",���z|[�HȞ|�p�����yB�˲Jb��۵ɑ�l&��K�ɛ��y2�ӫz��D#��9!������y��:u8h)�@��f
�#����y"�U�s�$s0$�eZn�Z�ö�yb@ِ)L�a .8`y������yR._8X���93-K"n��[�d��y��S�zV���g͢h�91E�V;�y�-j��	R&�8IY�(䨆>���hOq�α#��I�����!��Vk� i�"O\�x.!M_Z���-�eyBE��'�ў"~
g�
q����bL�`��dI�.�y"B�{�������S:J�c��y2�ʩn�QB֋<9r���r���y2�A-S��9C6��.Q��QNE�ybI��(��Q:c��r�ҍ�$����yҠT{� pi2d֑ihQdQ�x��'�<y�Pn	�GB�)��/p�d(��'5�r�~�����*y�)�5�'����^��)+��	�D����l��,Y!�d�e���[��h�r�8�Z%*U!��Swo��H���g�`%H�i�B>!�d�9`P+ ���p {G(&{M!�D�l��Ȃi4P�̜�e-��qH!�d.�Z��&mT�,��@��&�!���<K�BFBԕO��V֎q!�d݃cr�T:D�V�XlRlaŅ�*nQ!��:S*��b%��a9d�T�!�� Kr��(�J��B)`��`��[y!�$��� �$�ߢD+t�uj-C!��'B��C�K?�U��A�!��"n���D�o�J�$!�%{�!�ʾA��f�����������'��qct�C"}E��"���t�`4(�'$*`)�3^��4ҳ�\�gQY�'�,֛1X�����`l��b�'0d ����I����3|}��'��B&,H�IT�i���RV&�y�̯\���-�x�)��ǓZ���S�? �L#�޶o�D�BwE�5`�U��"OV�o��I��ӂG� ��"ON4��
J���3�Y�4qC"O��3恋"p�p���B��X�k�"O}��䔍`/J��� �Iz�B"O��C���-@,� �[ъ!m�.�!�D�=U�Q��M��|z����Py�ө�� G+�3L�a��V��y�kԷi�� ��F�`�#L��y�B43G��S��A���Kdn�y��ҧ?V`|���Oh�$�8Ԅ�7�y��ǛV��%I�� �x#AN��yBjӤg=0}Ʉa֖87�آ�N��y�D�p����@1�����yB�:5�j<�&Jk_赫�,˨�y�l��f�_����*Ȝ�yR�X1Mr�ID�ۤ*�~��c'��y�� 8��L(�D��#
=1���y���4V���d��k:�a�BD��y�M�j^J�N��q������y�˞
=�ܽ�%%�- �41����<�ybH��J0Pk畧t� ������y�MY"Ƭ�W�˞6s��+��yr	7l�`K42�r���OY��yb��<r��)�S<,:P@P���PyB���H��(ce��U�p���BW�Ij8���u��98�B�hJ<Ъ&�+D�� $c��Pۥ��&��}ꁢ,D�L4��}���B�V�;���14�/D�@3�F�=�^ٳu�߲[�m��?D�����W�7^N�s잁 6����<D����J�W�b��WÇ��t�m>D��bb� 3*T��r
F�QT��ы=D�x�D`�%hQ���D�םQz%�u�7D�pF)v|Q��U� �`���:D�`I�͟�4�^�(7,U�}ex��<D��8� 	&1~�X
��l�f�R7e<D�k�則��50�cԱ+b����'D�d�����CѮ��K�(Jc�ɐb@"D��9�I����ei4�V����M!D�2h��gd��׬�8Q$��E�;D�`��
�Y�t��O9��R��%D�p㣫�YpCY1�t��b "D��{�	V����3&�?^",��O:D�@�ϧG��a��ȫ9v d��7D�$Y�b��v�%�A+Y=*,t8EO+D�+�I�e̢�*eD)QT9��*D�L
p��F�=H��߽!��y�E�'D�������n8^jS��a���:D��Y"�P�� T)��/D�U�`"D�����C�]��M���n8�:�.D��ڂBENK~��#�g�;�B,D��@8yx�͎b�!�)D�ຑ+�%A�l�X��1��(�r�&D����E���AT�V�%J5���7D���Mۚj�X|r��y|	��B:D�(y����R"�3&@%hr��KC=D����ݛ}����7���e�;D�(`(	:-ͬ�h�K�\zrl�dh?D�@�/��/�Ua�K�+D(���=D�dS�?}�(�t��
%��)��&D�PQv(�8kf�b�8���($D���1�r�^��#���PX@�� D�<��'�_�nِ`a���6�"2�=D�� \�M��
�	s놯���(�"O:��tA�"z{�����-�@��"O��z�\6ƭ��K;L�8R�"O��AQl3L$>T�FI��
왃"O�\7�J�������ՙ�"O*I DA�ox�a�!P=Se��k"O>qы�;��y!�\\\|0`"O���abQ���ƶiP����"O�5����}��e��m&G�X�T"O�-��oF6�v�#����K�B�6"O�A�G�	G������אd|�""O�tZ2�3]���с��{m�ei6"Or�(d.
F#p�v-ɦb��&"O���ɲZ� ��k��j5D��"OU����d��q�(��R�o
#�y���)�T��l�7l��"d�Y��y2�M;J*��F�W�- d�C�Z��y���O_��I�jі#�|qbC��y"j�J�<��
"p��"�E��y�$��)	��d�ƈ&xk��y�gJ2}��
gE׃&���;G���y�ʈ�ތ۔�.0C��Z����y��E�^�R ���Ðu2�u�u"ͳ�y�ϖ�:9@I�� ��l9z�E��9�y�#A�i� 0�5'�^^]�s.��y���-ZK�TY�	^���U���
"�y��K0_��=k�$��N!�����y�fę7Z�E8 �!j�2P�IƏ�y�Z3�*���@�/kD������ �yr��cv�!k�&n�Pe��
��y2k��(}���ʌef�I��N;�yr���ܡ��/?a�~	;�E%�y(X
Wİ�,EZF��xu�Q��y-��Όv�ݚI
���D"U8�yr��*'�>�a�Ĉw���q�	^.�y2�M�+pȱ�K��taqC'�y��P!�����ѷ~d2�0�ѭ�y���3#n�+�k�!
6��,���y��]�b"��!H�v�:�I�U��y�	�'l6!*'ID+g�q���x�<�@��TH��+���.�fe�g�|�<Ѡ��2b6�˩w]�Qǃ�w�<q�c��sYz���N�)?�5@�w�<)T��^�
!A��ɩQު�k@�O}�<�L�"5��qB��`�>8���Gz�<��+�"}.P"5��w�rYy@�y�<Y�L�7Mt0� �-#(��Ud{�<!�,���Ě��$��@�C�x�<�霧��x�A�`�u�p'�t�<�4��x�-ac�?A}��k��|�<��FK�`�=HO�8.&x�Qly�<�DJ�% tt�sϷ84�;�#_p�<IT(�+���s����+eX�S#�m�<���p��s���,0l	3���f�<�!"�$F��r��zW��Ce �`�<��׮�؈jQB�8R��k�Z�<A��� �ܔ��#{4�{h�Q�<�ea��J���#�̰2.(��K�<9����T|���L"�0u1��E�<�� -
��T V�BX������I�<A�M�7Z�H ���!k1�I�ॏB�<���	{@�]rW���-��E���x�<9V-�9A�H�e��D�ࠓt��s�<I� �)`1&zۖ(�8c�T�<� ��$(G�����O+>�r@`�"OD$P�'��s�,%����h1��"O�h�5�ޏ7�d x���7I��s�"O����/%V�@�@�7�u��"OX@�!O�*[Qtk��@!�I�"OH�8�$DZm14MW��4p �"O���jA�p���1�擕]��Aҥ*OD)#�@�:i�`�砇5.���'��Y1U 
�7I�-J��:B�l��'Eֽ�7o
$�պ���*�RM��'� 噑R�lM;D�/����'LZ���/��ِ��"�����'��$�C���lB��c���+:��
�'���3�	yn��`����)�'�~�X�J��������9�',,m�&V!uD<Y#t��S$V���'m�H`1-^�; �٣Ё�Q��t��'L�ɓd�ɕ9ppX�
M�
��'����C�&[|d(
6�]�C�����'���8���^����@�QG@�p�'��|��o��=y���$�2I�~-��'��i��-�2����T��]��'b�m9eK�*ex�#�L>�=��'����c�8AJ,�:�D�*=��DQ�'�V��S(�5��� �2���a
�'�lUy��#$�Ҳe���M�	�'�> '&ߣA��H��;Y'4���'q6Q80j\)@fD�hGE'�8�'ݘٸDIV:wWl��D�%Kr�*�'�jP��#H�N��覎�+;�8��'�)�a
��;o��R��W���P�'� K�Ls��a�ѣ xXL:�'è��R	�2g|��va�8��@;�'lZ���d� r�3&4�d
�'�|�p�ڼi�P���-=<L�	�'�v�i��/�D8*����7����''z�)�\�3�V����5(܊�
�'\� ���̞ F�h9AN�8�� �'�� 3�<�j�(P+���'u�U�g�BF,��K��:�'y�|�ÎX�T� *S�D!C����'!`*녞,60��+�V(��'�Pu׉��}�3��O���(�'A��1o�9B)���O�:׶�ʓ����`�ѩ�2�8U���Yl��ȓfrX#�*9��Ɉ�aǑd�>�ȓj�����:!�`��� c��ņ�2H m@2�Ϭ=*ҬA�I��Gra�ȓKo�)A�r��%8�7g����=���D4��# �O�9�� ��T�A��U��L�+�k��	��T�ȓÖ���߶�D+E��qʔI��o�)�S��42_�3��.7L���ȓF�E(@ �e�HiJEA�bv`}�ȓ/*t�p/�� ��L)s=�	��?}&�B �!��P���;k7�	�ȓu�޴U�@�/�,���6In	�ȓxPt�AV�z� ��!@�4l�8���7p�e�'��D˔u#v'�-|��!��I �@B"� ,U�T;q,��\	�ȓF�١u� 8~J�����#�:�ȓ�n�:Rd.Q���
�|L�����D)�����Q�ZJ�C�I?�8�q���(/ �$pA��G�hC�)� �`�V�DT�Zei��K�c�]��"O�Q��8���qf���;�"O�9�d@\�,�������v����$"O����A�b����#��o���"OI��!S<qڗf�%VP�8r"O������F��⒈�>>� I��"OR%ڳk�.H��A�F^e�4��"O
�)��#T���jRF�=�J���"O씺ӈ��b)Z؂`�QOR����"OΤ�dHF�FXj����$aFu""O���tR�]q�1$��$mj^��"OZ�Q�F�=n���	�T����"O�t��[ 9�ֵ�+�i�"O��5cޯ6>��iE�}�h���"O�h��L�d6By)��O�o�	Y�"Oj	����ö��`�� E0\m)"O�lp5�?)�$�k��	@���"Oމ�`n
0+��#�D�s�A "O�	�)�>~���%dQ�.b`H�"O!�J֍i:zi�f��*&�	u"O�����./���Ǟ�~Rq)�"Oʄb`��4\I@�r�h]1j���"Oju	�����F	x�i�.W����"O�]��/��"`���E�V�!R"O��0!��1^]�uqt��D���"O���Ȋ
,�q��J+ax���"O�� ��-wpȒ�F�2V:���"Ox��S�O��j�H�����8c"O�(���	X����޿3u���3"O���H��y��B~r���D"O|5S�a�	Xa86b7�9�"O�e�#2r�H`C�0� �b"O�	b6+ե"$�t�EJ�E6T�"O�)��C%w��U����Z"O�}�"�S?n ����$W콙�"O" �f�(2p�bDS0�DPJ�"OD�0J��H�@8�!ÆiĆ���"O�9��.�
{��;��65��0�"Ola GLCAfd2&��y�P�!�"OtE��MŁ-��	��+w;��qq"O��dς�Oa!;���U9�eQ�"O�A��ɾ:�4��G}%(H�"O8��@��P���*�f�4*��"OHPP��Y%~ޑ���ەe�&�pW"O�e��#a�Hm#n��i��}*"O�|���4��@3ȉ`vx,[S"Ox�D�P�%�����5SR�A�"O���3��� ߲�� @.?Ot��"O�U�0�l08�Ă�k�6xcr"O`l��@R3@I��E�C�A�!"OjDW�ԍl���,z吕B�"Ot�0�/ #z��
��8�"��"O�0A��T l!j�cw�CȊXA�"O�$(�lA<g@�qcB�G<;�B�q"O �z��[�)�B�yB�#�2�r�"O�(���&�:��0E$r�pRU"Or��DeI�X<Kfc��\��U"O���Ǩ��^>�!���U�Q��"O8�"ӎ"}�츖F��8-��	G"O��!Cl�7v@2k5�R�S	�Ř�"OZ��&�Ɍ �
E� #^��&u"OB��eY�K���ە�Ө
œ3"OvT�`@#`�
�taԚ�܁9�"O�{g+��k����`�<��A"O� �]��e��u���`�?l5:�"O���`F
�̅�b@4-&�q��"OjQ�p珈L��181܀;"J�"O��
ģȒh��hANZ�cK�}R&"O�=�%_�5��wm�*��e "O<�ka@��Q�6d�Q�O
_���Cb"Oؠ�K�9t<&a�υy�F�R"O͹uV�d�s��%G�8K"Oh���#��F����� R�B\a�"O9A�#xE��F�V��:�6"O��V�8��tE Iop�D"O�x F��	������AQ�4�T"O<]	�m�E^@�c/P0<� �7"O�E2��H�l�dn�!%��!q"O�<�w/��"�
��K�O��\Q"O�@�T'�}*`-	"m��?�9x�"O����Z�+��$+��~&}�r"O~��C��8� =j#�*QA���"Oά���Aq��䓷�°3OL)p�"O��jqC�="`6��h �*1�y0�"O��Z`O�*X�$�w�!�%+/D���`l׈hf�Ũ�IJ�lM��`&-D���i�^i� �c�.�����)D�p��>pf�)uBӅ�p]H'
'D�t�ohp b��4Il�Ĥ/D��RN�Dpx�'oZ;��s�+D���f�\�V��sKL�"��<�Pb%D��b��@
���D��RDĐ�W"?D�p�ŹlV�	c� ҇MV����J=D�ȣ�lP�`��M�ф!�(B�:D��yv�G�|�$0��E.#��|*��6D��&�LC�`����9�����2D����֩u�9�$H�?����+;D��&��,�nY� ɔ�At���:D�DB�ȧ<� Z䏇8hMH��U�"D�dS�O>�&H#v.��*{jE�Pe<D�$���1$n8:�˓�kL�;A?D�����d��<q���{1&т��?D�|KB�ܡH���22������,s5�C�	�Y���-\�6�!�dO�6�2B�a�pݫgB�4EltJ��@(S�B�	*r�,y�W��7�N���ߊ6�B�	���,;�"ٽ+���I���9x
C䉅n��q[�?` ���*4H C�?H�Y@C�֍n���e�G��C䉔cb����bR4(扁����,A�C䉹n}��hq#�+-ɢ({1�]��rC�ɵ{��`cg���xT���Բ�'@Z8ڂCN�)֨�g���K�'��$C��Ly�us%�f�� �	�'��|��%�18F� DE\�d�i�	�'Ϧ1�� ���-cs�C�_���	�'�6�I#!��4;�@��Q�H��i��'��أB.A8Hf�|��gA�@�@]b�'�`!"��5:v��\��L��'�j�ME����`Իfn\���'˰����0��!`cKڝ^����'
���Cõ��
2��*X�,��'���p�Y����T�ٚ�'x`���3?y����4�)�'�6����ۆ|,�HBF>@��5�
�'tP{�B
02V�y���8�t,�
�'�XlZ���2��$��a5��l��'``�Cgޘ����� )��A��� � (�"?��*q�ɏc�X�C�"OP�E!�. 0�	_��{�"O���HG4;�ؽx��<\N�p��"O�R���	l�dٛs�@?lC����"O"}���˛T���	S��	�ި�v"O�e���V�*\�S�O�w]P��"O�!���W�+1¥���^>3�ȵ!%"Of��g�/ k�� p�;#�ΨIT"O�x*��_�"���d�3{��)t"O�=��f��pg\-�5��49`���"O�x�A�()��g#Y�Ch��'"OB٫��Qj!�Ģ�(g/�r$"O�Y�Pn�N�:m�����$��@�v"Ot���杄z�✢���"��#"ObU���G���ci��h�4��"O@t�tM�km�}{��W�ҭڠ"O�!{ƭ���`X��j٧lg
%�r"O�5y�ˍ:_戕�lA6`. ص"O��� �	�<���KX#~\��j5"OT��B_����"�B��ȸ�"O�b��h�x���c��+y
�P1"O�4����WVt���ǣ~�sr"O�x��n�@d���'h�T\Ca"O�lQ�ʔ�6�1�H�U< p"O��JEd��)�����Ї\G���"OP}���@T������F�* F��r"O��g!��H�4!��؉�h��"O�4�5�I�A�����k��-q�"O �g%א|4h�b	�b�W"OF����l�<ే�0T�6yK�"Oz���� �t�@�F?
7����"O��zD�Xi��x鰏�<-NC"O��a��TWL~Lg�K�TR̺�"OBl�q�H%�L��N���!e"O���lQ�By�� �-��m�F�1U"O
M;�l�KRRܻ�O)p�h���"O�Q+�
#9��Ϋ��L�P"Ol�	C̃;�^]�$���8�� "O(M�NXx;P��)פ}b�[e"O������H	���fgH�W"O�l#N�k�\J2d"CH��R"O��*��#�B�2T��.��}˴"O�M��?PE�� �Xy��+7"OH�J��)$X0�;o�>IftD:t"O0Ռހx7�Ycm,
Z�-��"O�j7L�zv�B�yRHP�"O�T��B8u�ܬ�Ł� r@�!�"Ot��ȕ�;NP*d�Q�'&
�+d"O�YqboD�IgX�9w$� ��v"Oz�x��-y��a��uv��"OVei��Ɗt�����a�X��"O@�pK'E��9u�o�u�G"O6(H$�c�H%��ҷ Ц-��"O�	�I�	:U���7�>�Z5"OX��4%��#����g��Nt��"O�"cǷA��HCGɽn�$��"O����vF��������"O�9Y���+xrihg�:H�@XD"O\�*� P*V��������Q"O~�F�����j�%N�l(���"Op��Q�X�E䈃PDƀK.��"Ot`j�g��q�������b=���"O�)
�j�a  P�1�K.6�yh�"O�h�W.�<��(�ύ��p��"O� ,L�ƯSv޼�ڒn�%{2��A"O"��夕:Wx�;m��mg~��"O$mr`���LtqF��Ie����"O�=;�.K� ��p�G�86GY
t"O<����>C~�	RlB�< |��"O���W�G�2����g�ۭ|�X��"O�0"�NZ(AR�i��[��(��"O�ŲD���dA��	J�D����"O��J�`��n���x��9d
��F"OƩ 4fΫ���*�DX@\ ��@"O"��O��E�v�!���!\:р�"O�g	�)27�ӕ��'���"O0�0v��eC�`�%-�72�"k"O�"$�	cl��TM�?{�[�"OJ8
�n��.���`�̦-����"O�8�S��l��t�U�Q�i�>%[5"OnA7�!=��+7�A/@���ʥ"OH��Kͯr}~H�2�_-j⡐�"O�U�� �2�fUh�	X�QV�p�"Ot4�ŨJ�ن�a�hG�I2�"�"OU:dˠqdx�5p)��1V"O]:�$$Miv��Z@3���"Otă���OWP$+��"5uJı�"O:}jcN
X�A��n�2V$h�P"O�Ez�`�^���M�	yb�찂"O���FhG
RC�l�6kRE`U��"O�}	����l� %j50�-�"O��Q�!7��-H�f^+k���"O25�2E�M�T���+�	)�!򄝿O4�1G��=v�!��&@b�!�$ĝf�n	S/	1b��
aD@<rK!�dI%3;l]�;Ls��{t��! !�D��[�|��h��q<����M��!��:�2Mi6/I4����0r!��;ڠ� g�hN��h�"�+7!�$�,���sL�E�*�k��!�!���z�(����� 8�Uc�.c!�YP�����f� �
��8D!����Jú�4(����]���E?!�D	ȼe0Q� �e���� hM�/>!�*Ċ<xB�N_�Zē�X�"!�d�+ߨ����C�`}���2�!�d�A� �?'O@�����%=�!򤎊���2�G�����ĒX�!��8'M��"�=*�Ru*t�Xq!��}Gx���$�:�4�k_	qa!�$�O�������U\�Mb3�ǨQ�!�֛H��y�1�U�枩Rr#��E!�S\)�$s���1�څ��□3!���!�J��o\��p�lɽ�Py�H	�4���ɖ#�((�5k�-�yB��8�yb��sEf�?�y�n��a|6|�BJT$k�!9�%G�y�f�<���"�l�%9(x����yrF�/�l
G�4z�jtQE��y�˔	zz}0$��]��dq4ȇ��yLI06��,Z��q��k�,�y�g�	0�m�ҍJ�M3n��f�-�yR�]N��,OW3L+�s��Ʌ�y҈I1vdРo�?��x:ҬZ�y�/Ƒ6&�pR�ǍV�(�@�I�:�y�x(Qթ("��3F�K��y�↴��}ٓM9�$��t�*�y2�G*9��ե&��j�.W��y
� ,0���;dt�Q�曼�*�f"OFM��� ����/.�+g"O�lh!��3Z��h�oն�ڽb�"O��ƋJS��� �3~(D��"O A��	%�Ѝ\o�R�"O�h�%mK3b���!�V&l�<�"Oޘ�`ˢ ɂDzAd|f�"O6ًp�߫Y^�����ѓ\J�ˠ"O�9��O\�P�"�D�X'JMd1p�"O� uo�(|ƈ��,�*u׺��"O�ó朌O>X)��
Q�(q�"O^a���;`�1���%~�X9��"O����FRnL4Ka-%(Ѥ�#'"O��a斷 yݢ�Xʹ�"O��
f	%lNR���k�:EB�"O��ք�rE�8��I�V��h��"O����A"
����� �� y��"O ���!�QNEٵ��x�V*0"O�BJ�:*F.����P]eV`�"ORTj0⒴dQX��$%ޯJ~����"O�a�N�+�2A�D��u?�Ă�'�<��%I:'uZ}@�I�0$~ei�'���{��:p\����!z1�=��'�s'��8>h�`KT�{�D!�'��)��H!M �0]�Cf��k
�'`�1��D��@�fHA'ú'@���	�'~���"�B�N(%��C-,3�\��'�� @ �7� ���'+HRD��'�F=�&3K|l���cJ�"E $1�'�y�� ��fP �����!�Ľ�	�'���c���ntz%���Hk
�'�x�`B7�^`�5j��
�']�S$ K:��3'W!,u	�'��|Q��.1{��ps�ǗC�Ƽ8	�'<��4�A�#��Q��:<||+
�'���CB�žW��4�Ql%je�a	�'��A�N�Hh�!��;d�X`k�'�<@�� N�{����&V�U����'� 0XP��G�xp-ǭM��s�'�N��w�Q8J�,�s�gșy� ���'(|�i����BW��S�Aӗj�0(��'eh-�`m�,Ak��x��A;o��|��'p�T��̝�[��!�CkCjl�\��'��)ڦm��D�D0QR�ơl�����'��f'#G���� PS��C�'b�U9R��.0���$�?o��(�'��r�Hևq�`�A��/�k�'����J�źh!��.7�!��'w\uQ`Rc�r g�#�n�!�'�>�#�a�a��(�7�J8��Xz�'��`�D1� �i 䗋TJ�k	�'3p`�.�2N�~	�wm]y3����'�`� ͖�RĀ;0Y�s�$��
�'ւL�P�kcB�)�hݎt6杠�'+TpCE��Ze���/8PƜ��'C���� (�ޱZ�Ɍ�*PpY�''�Mh`&ͅK=��s�(ޕ)�"-!�'���#Q�J��YƬ�$�<�'ܶ\zS���KЬ$��g�6Z���'%�]����|<���@΍�=��'�Za��yz��7��)B�,b�'����Wf$A�q@ʃJ��H��'�����o�3d�M�&�8=��h:�'\\�1���*�� WO�5�<�
��� ��R� 8`���\�M�"O���3�	?d#�Ar�J�j1�9d"O�y�t��	#f�i�)5lIn=cv"Oe+cװn�4�u��Q>z�s�"O�d覯@�*��Ѻ���6s ���"OPE9��ޅb����ф�-p��"O��2#���A��CS "�����"O����'���8��v��~�����"O�@�� �N��b�GLۄ�p�"O�y�g�D�iޖ\�QG�B��X"O�kr��lȜ,�c��`|@�"O:DQ���Ԃ��Z�1��@"Ol�R��D#0���3	e�iz"O�ҍMy���yCGܲd\n 
�"O"�	���]y8@��f�?��$�"O^A)K�<q\���E��V�,�sf"O��VϜ�K��f+����A��"Ot�kC�ļUsĜ�LT�����"O�sI�9�V�AG)G"r`q�e"O4\{R�>N����/(V��˕"O�as���7���A����dT��5"O\=q�
��|��mA$��PA4y"f"O:y��k��/�Ij��
�E>��"O�qb�5!�h8�g6��+�"O�ȳ����+�dE�C�P͈�"O�`�'IĶ?���S� J�P���S"OƜnN5AVT�h��U��pS$-/D�� ����<��C���IG�@#"�!D����oƢ���0�3��uX�>D��cf�|eH���#!o�1�Ο�y�CG�����劖�9~9��# �y��Y73�6D�P���	�,��Ƅ/�y��:t�`�Q�E}��<��m�'�y��W�2�P�C�"@J6UY!�͋�y��Y*q'��Z/M�*����Ȳ�ybnGlS� �'ۦZ�����yR�5������3���L��y����I���6%B(i�E�y@�w��8�sfp�ti�BdC��y��s����p�i@�ѳD��yB.������I	p��xS��>�y"J>x���i�<���1,�y�.��fx�&G�/4ID`	�B��y�# 4T&� ��h��?ȼ(+so�y���;Yv�G�ٚ3{�yRf��y2�K�Y���B��3�����H��y�eH<M���p��תŲq�B��yB��?�R�D��q�j�(Ѧ��y�n�_C�|���=i-� ȵ���y�CM@�6�X��:d�T�AV`�;�yB�� @c��;��A7)j�� f���y��k�x)T卫M��L��M��y�JϫӮu�& �+[����af׋�y���n쐒 5, #!&���y2C_�-�4�#��G+Ev�r��S��y��1Z9&]��7M��	p"��y/ӭi���{7�)�J�� ���y�E��6�K�L��%�r�9QKľ�y�GK~���g#1ڀ�7g��y�B��kj��3,M�E�D���^��yRS�P�F�D!���7'�0�y��ܯO�J�����b���F��yr@D�QXl�ը�|4���Wl���y���Ȕcb
�+I"��g���y
� �)��ڎ&߂�	����Y�}s�"Od�2 ���
���:�kجs�ڙ:e"O��rg���I�da@-L�A(H�'"O��hd�ߛ<�N9p��*/%����"O�����N`�ܚ��V@꼠�"O�`�〭�&B�#���`�a"O\�B�O�_���˵gT uv,��"O��D�ށWƼ`�'�ʩ	ch�H�"O> �OC���Ra��fh��"O@X;�����ܲ�CN�}L��"O(�dAJ��C��\�%G���"O|u��K��O���y���N��ef"O�pI���y1���Cǁ<����"O�eۖֱ��9q@N/H�F���"OP��ccO8�=����:;�<�q�"O�!���6S�-��HQ�]":U�a"OZH��Y�7�И�#'_X� ZD"O�����n*�V旁|T�"O�邴��'4���CМ�À"O��+s�϶|���(�	>Ħ5��"OzE�@�S�,��3�P�+#�P�"O(�r)C�M�شۡ���
��"O|ͺʒ3'rA���J;A���Y�"Oʤ�pm�2J�r� X�Z�^��"O��C3^��qd�f����"O���� Ƥ:z�|�q,^�(�7"OT�2��	-��h[Uk8~#҄	"OR���Eot�q#�J��2"O��w�2/�����'�yΨ��s"O@�旼p�~e�@��' ��"O�4�uf��h{R0����V .��ȓE'h]ڷ�@�c?b4K�	��~���>	d ���ݦV3�m� ,�"Uߘ$�ȓ@r8�A��_ ����̎"s4���~*�Q3���8��1�!��&�Ňȓ1?B`�&e �"�Dl���@"|r����ԉ��d]cx�Ԑ%��]6B�����6F��n�0r��(}K6Ąȓ&�P�!$�S$A!"���@�'��Ą�QzF�6d��� �r����ȓp&tk7��k� �*6�B�ȓY:$�v�T�*�~���[���ȓD�LaS�@V$|5��s�� 3����F��|���K,L���rI�?I�|�ȓll(#a�փ�L����=�le�ȓ�z��c��&�R�a������-��&<(P�2m�}!�Ꮪ"���C���)�,YY&#�<4�D��-w@1�!kZ�����;AVQ��r>&��!�u"N��c�N�aZxD���� k`�K?.8(��2�����,��A�%ǎ�N3�}�d�ŵx����Lx��2�	/[�hK��ܭcU�ȓc ������-Q6F�#1�آ9i�x�ȓ/J�	S��ɂT������!A��ч�|���k��¤J�9vm�����ȓGu�
L�A�L�:Rȕc�f}��f�:��"L*kcX6�]r�܄ȓL��T9qGC	��
l�/c�^фȓ~@+�hLm<��u.������ȓy�4Йj�#��E��kE�#SVd��S@P�0S�ߪC�0-��
J��i�ȓq���17���sҘ�`ƆG�V�<ч�>��٪�	�y��(�J��I��S�? �<�����Fu[aQ=HAr��@"O����^.y.��En�A(� W"O������!� 51LY�H�Ac�"OF!�RCJ�\x)�FKP�
4�HA"Onux��2Lg~A����f�E�U"OiX�T:h�ֈ"�I���A"O�$Z��U�Y���a#�۳,yJ���"O�y;o��e�b9*Qp�ʜx�"O4��G��f�l�X>}S)��yR�WOWx�8BAZ�]�HY�"AF)�yr	�=s>�ЬǮM2T��
��y��
>!$8C�a?�<�bM@��y�eí&_�m3��2=p�A3�׋�yBC�g�Jhz`�
8`��ɖ)�yR�US���z6,�8M����و�y2�^.zc$}P�BSc体��y�Njr<����0��@fF�y�g˾f�n�Ae\�/qՂ��y�È(���Ն4p��a4��'�yB"�7^\�p3�ۜ �|)��FI��y�&�
^��	k���Ķٱ6�W�y"�I4�`}�!!->�4a���+�y����>.�X����&}+a��K��y����*\K'�S�b��L��P�y�аjx��7f=W�L�)�i���y��C�����P�S�	ԉ�.�y�m�54g���`UT���s�iP��yk[�b1������O|�,��hQ��y��Y�}Ȏ����6�L���>�y2�Ț ��Uˏ�-c�<BQ�Ö�y��_3��P�E�	�5r� b����y���5+S�H��I�,�&ٳRC���yB��9_F �W'��q^dR��1�y�(]��i�/P�u�p����yb�ȇn����t�����ܠ�y2�9k�����p�(���U��y�0!.@"�Bџb躍�	�'���jc�/s�m��&$@��	�'`�A;a��><&�����'�	�'��qH$�K6
�Jp�H��^�&��'T ��0o���b�ڦeō@�n��'��5`Db�?/��[.�)*^�IC�'�;GF�Q���rU��$�Q(�'���T�1P�c�����=i
�'=ր`�p-��Qԋ��p9�	�'���R�
Qd��T���(���'m691��WJ,8���{�@�	�'�@y���8j�+�O�������'�)Y� ;�'ԟ�F�k�'�
�#F��e���@0z���'�ɉ�kM9,��iw,ЂB� � �'w"�X����&�:)K ��'ŌM*� �y�$Pb�	ͧ
�="�'�$�u�m�*ܐ��656���'�.$ ��ґ
~�%�à���'���	�hĈ�3	[�6I;�'����D�~�,�&@ǀN b�	�'�t�$aͺu>v��&K�#B�V�;	�'*��J��)���Iŝ�T�I��'�
��!�^���&��{�n��'�<-��%BI)XuvG�#H��S�'Tl!d�ȓ`���C�*��H��'��]Sf��|��aipq�B䉱~����KF�s�N$�a�̪5��B�)� ���m�/pe�Rt!�9'P�!�""O���Ug\�e�0
���Q,�;�"O� ��d(�2%�b/_�8�z!�@"O����fϾ��K|\07"Ob��0���^e4�z'gO�Rl�"O:���$.?�q�P(\$�+�"O:8�UJU$?t8Q(��I]�.1:"Oni¤�J�F��*ׂ[����:g"O��a�L3zg�19� E= ��%��"O�i�����;��4�΀!""OZ�Q��f@j����@~�t�'"O�k�$�0o�6��f�f��]��"O�Ys7̖�sC�����Ps"O&�
@V�<Ԩ��!#S�}�\�(d"O�xB�j@�r�>]�bR����$"O~p)��ʜnɊ�u!��\���"O���D�x�Q�t��=�ڍ��"O��cZg��1�:V�~=;P"O����ǰ�m�t��C�x
�"O<@x�f�=	�E�C��>Ҏ]��"O�0)��֖)1�Đ���l����"OR��(�l����7~|�ei""OR<IC�F]��"Ю!N�l��"O��kϛ�WK�~ܘ�s/ˑ�yR���m���7醕z��SFǡ�y���rQR0�,lTN [��Y*�y_#"t���p/�e<q��g���y��tN���F���� 1u�K��y�e�� {!J��@	Hr�Uk��y�P�x�z �P���,5 =�o���y"�C�YQ��7$X�!�N���>�yңoaUgU�F�
%%z��{�'�~8� ��*}��R�Í0p�ލB�'��Z� �4����c�����'x@T!���; Y�i���C�c3L���'�4T� -ڈj<���f�ʈZRnl��'t�="�3�i��
|�yq�'N��I��9��83����yH�'Y�[$��8Z�0UH]�(5 Q�'�"I��A��{���AgT�PT���'\p��e�A���Fe�0���'˜e)R�΍lR���� *��
�'��Q�� �^�aM��K�z���'��X��⛺\����O��Fg��
�'/:RMw�ji�f�Ҍ75���	�'���*abk��F�1:�nx	�'��Pk"eZ�r�S1B�[r��'v̠J�b��4���U�d��'��0U(0>���YҫPK����'���0��ZAǖ!rDHQ/X�@(K�'&x��u&
i�����(��HfI��'^V�abo�!i�R|��&S2v�+�'��܁V�>F��:���>0xqC
�'�-��,D�j�2�F��3�xHB�'F�%kw�M:,������[+<�R�P�'���P�J߃Ɏ%��5o,�

�'�ܹa�i͟8�Y�G�WA/�YA�'����VB��5�V-�͗3gx�r�'Ѿ�0��ŃS�����/��H�K�'ʲ`rA�!n��#�G��q�py*�'���ȵ��J"��x�cX�dBP��'�0a�Q���;촥���]8����'�(�ӡhԫ w(�������|��'M��5F*J�b��~�8����� ��:�D�9rȜ��cM5B��{�"O�( ��˾o0���آ9���1�"O��7&��G $��d"��[#�bV"OJP�	�f����@��kB��"O ���I����#��"O6 ��@l2�`��]r�DaB"On��a�6Z��y(����^�"q;"O,T�G%��+�����K�3��	�"Op���c�g>�CgX�r,��f"O��ש�!lz�D�S�>�"Q�"O�Py�K��{�.�WeӡZ��ȹ�"O�]q�N�O����P�[�H)[�"OV<[u���f����Pj.@�8�p�"O�A�B%�ؘw�j����"O<�ꕬ:h�� �]�2�#"O>X�0PtsV B��ʒ"Or����4�8�9go��kŮ�04"O��x�P#]��cH_
&[�ݘb"OH<��EK�`VrQ��%�+SO��9�"O��b@�*D�i'�y>j��q"O>-Hd@��-p� r��
sǬ��1"Op�C��!�iX��N�u�J5�w"O�q���k�L91����X�YU"O���(�##������h�B$"&"O�BQ�>g
�����W�`��w"O���+י:����ŗS��s�"OR��`�4����A�ƥ-��e�%"O���f�T>�a�NW%4��p��"O�E!Ӆ>߰��X�l���� "Oj�`�鏻�4+��҄�i	�"O�(��1}N*`Z��� "����"O(��F	
:'x�j�N�m��"OX��/۾=�B+LC�5V�a0"O��#LpA��HS�J�!�Lu��"O"pA���.J�B}�CNKX@Hbf"OX[�5e�8!�cZL<,��"O:�O[�p����[?E2�%�G"O�g�$���#`5*lҨ+D�lc2m�&�f���ŀzxd�z�/(D��ZՂA6mT��Su�<ZBMK�1D�L�S�]�>\�l�NP���.D�4��.�>�r���� S���ch,D� x�-��]z��FWb@ �)D����
�~��AJ�'߿Xw�-1U�%D�4�ďT)�j�aQ�GZ��I:�m&D�г�ֶY.8���#� �����C*D�@{A����
�`�?���q�%D��Cpa�BlvЄI�H���,$D���ϴR�
-���'l���Bl!D�d��͐|�ę��,'|�5��D>D���ťQ&qt]��n]�M�y�Q:D����G�7r>C��:��Q��=D���seO�Jܕa���]t�5�cN)D�4j�A��g$p�-M�,�T�j2J-D��G�S2A~k�mˡ,C�
�)D�X�gAF^����1~3.�G�)D���'����*eg8��L)D�T�fϋt���b鈤\>���Q�*D��z���B�b�G8)-\ݩ�(D�@�@�. ��@b!��*u�b��f�;D�8X� 4�JLSf��,>�遈6D��C5��e��^�B$�2'�.D��B�W2�Q&-q>�9�Qa9D� ���;R�h����Z�f��Y�c5D�� ��`/�nT�2�,�w�,�"O���&@� ���Sۣ7ZY�P"O`$��N :������Y�b�� "O����b�@pק�� ���r�"O C�܆o^$	�l�k�B���"O�z��ۻbO�2�*F%)�:�`"Ox܊�E;r@���kJ 4r ݁"O �+ck�o��5��	ߴsZ`�c"O�QG,�&�je�R�a;�"O��� �.k�^�J�+X7��A6"O p0鑋a�H��E�!,'�0��"O�4���66���k�̣a	΀��"O p��E���Ma���=��0�P"O�E�b�IP6�8�m�,�d-�"OA�$%�<�� ��ʀ*O�M�@"O���r	�K|(9fF΢m�b��w"O�`��r�P��4����"O�H��J�=@^:�	U`M_wX�h"O�	U�ީ[0~Yj���(b�uX"OV K�	���*�IQ�J+EHJm��"O�IC�"
79�\u�oˣ�Re�"O �2��<$�k�k_9/,qSC"O��a�� Xc֐z�jͶT{&�*�"O|�Z$���`4��R#\oU�"O�8� ��Qd�cB�A�N@|�"O��RǑ
-i~H�&c�m8֙ V"O�Yp�Ֆb��rԀ�5_.��q�"O�e��?r�f��G/��_�N�&"O�kAjۥ����Y--�~���"OV�[!�|h�Xv��0���� "O�w��)xD\}:�l��U��y)u"O����R��H�� � (����"O6��ɋ�"H����O9�ݚw"Op�KT�R$5�BPT��I8��%"O���֚#��'˭F���F"O4@���Q������`��T�"Od��q���"U:E�����B�"O��r�\i- oU�-(6��"O�ݛ��<̬4������D��!"Ox�+�d�5\|D⊊ajT���"O�`@4��4jI�9"`+��^&���"Ofhs��@�D�jIS�IYKV40�"Oz`BR����Xt"h9�P;"Ob�
��F�~Z�M��Ց63��8�"OМ���U9��,�*}n�J"O<i+U�S�u"ia��R�fz�I�"O�XI2�6l�Z���/>�r`"Ot��G�R�]E��F�R"/�����"Ol"���:d~�s�,g���ل"O0�[ �/]��Z�aٯzE�H0"O�bU�R>t`0<�!®M����"O1q1c��t��P�a/L�:�,��"O"���"L�8��=� ��?F�$"Oz��1nW�H��&l@�=�g"O�r�CL N�l=.)w�iE��y���jɡ���Rͪ4J*X��yr��2}� vi�4��5BMB4�y"����uR�U�24��UF@��yB ��)���Y�L۹<�j�1eD���yb� i<�4���I<6^����y���1�������~(�M�4��yR#$͢=Ӥ�݉|�p���yb�P���D`QK�E�z(�#�� �yr�Q�S�,�ŕeeDI�R,U��y
� �Q*�(]�)luY6��,g�a"OZ��iUV�>D�f�5w�Ei�"Om�%喺@���P�۔1a,�j�"O����c��;�ʴ�2��2E})5"O���m��9�JpR�N9GD�ģW"OL�� L�+l� �Sb�$4&rlJE"O���&����ڃ!��H#��9�"O\�3C���6�q�JO�}�� ��D �S�:M�DmP�D�)3Zz���.R�?Q,B�I-[ p�cLI�|Z��3�ܤ����ߴ�hO�I*5$X�`m��G�MU��~���D
2fF�=�ǧ�@3|#O@�P���je
O��J�)2�h�8e( 8�����'P�Of��-U���LJ ͇H�
0��"O�u��$��"��٫Il�X�"O0�("f�r�J��B���0u�0"O�d�GӢV�Q�2'^�G���H�"O,�G&,���l�H.5(E"OP�K���^�80J�Mb����"O�1����q���b��+[wbx@"O��y�V���r.A	E]p�"O�Q�2%D�K�\)3��F fhX�r�"O��������5jAȻ*5#�"Oj�C$4p���.sF(�q"Oұ�BE�#J�61��ɇ�<�D���' �'�r(�����&������a�RM��'�ܴ���E�p,Pb�" L�Ѕȓ�\-�@V� S@�����z�bY�ȓ:���	���0�$��e�T���x~rBN������hF�{8pDO��y�^x̨VN�?y��57 ��?����,�¹����/=_D�+6�3e�4��ȓR��9`O�Zj�3�˘�	>6%�ȓq#�ukƠ0b��ٺ%+ǇuWp�ȓJ�,� ΋�Z����՝�~���_ҽ��I. k�c��R0��V=ْ��Kb�I�G��|�H���t�H��Da1\�aĹF4v|�'#ў�|�L�E�(i;p�կѶ�dlJ�<iF+��U��,�E��qZ#�o�<��IV�։8P*�=^p8RW'a�<���3���2��9�����)�^�<9R�]aP�cc/��svЩ��d�<QD͛kb�3p*J��I�/�b�<!�(@�&{j%k�@0t������s�<���Q�d��@�g��r�m�<�@�Sj����^((h�!Q�f�<q&�K�H�D!n�x@CQʀe�<1��� Q2Q#�g�
���_�<���N�'Lx h���\ú�6h^��������4
= �T%���Z��8�� ����)�i�(邷͋����ȓI_���L'>���D�:_(��ȓa�^���A.,�`��CΓQ��!��2@�vъ�X�����%oSR��ȓ-ɂԂ�LӍ3/Ƹ�&/ĝ0�م�.�J�OЀQ��q�a+�m86���Wg�|��eʯ3��< ��<4�t��ȓWJ��w�D�D���#�[IXQ��"��A$Ɉ�e� 8�ƞi��`��r�#&X$��|�2��"��GxB�)b&g��P�U'ȴ!���w�~�<���5:�����#��8���x�<��K]�B, ��i"�@�Ms�<� X���ɒ����#2A�:=sP<�"O���?i��	��2r�i!w"O.��w��l�^�0���ch=8�"O��������t�Ȃ�=g��j0"Oj���5&Hr5HF&C=7Q�Ժ�"O<��q��2��b6�2dޤt�6"O��r�",8�$E����b"O8�s��.?XT��G7Zz��6"O�� ��J�QZ��
�oK��y҄R�e�u`�.� U��9�+���yb�S7�f\��D
�ʵ̋��ya@����KIΪ*��T�����y=�}n�O�n����Q�y2��<.U0EOD"`~Ji�q.L�y2	�}N�4	�%ǃQ��M��,�y���H���:���^$-`�-�6�ў"~ΓZ-v�9n�G2�}�G��	�| �ȓ �ڬJ֋�K�x�	u�J�K����w?�F����ǋ�*��!K�	p�=���<���O\��Q,C"(ؤ�SE̖�e�I��6O���$;f̸E��'���h�쐀Y�Ov�j�O�pHסr����#�uвP
�'�����锹4���Q���\� t	
�'(�]� k:(���ٷ'�P@8!B	�'I���v�/u`��7(Y#M��l�	�'Ѻ�*F'
�@��M�Z,�l�'f�x�AN�j�̐sw#�� ��'Ӑ%�B���6�7��z����'�ў"~�c 
"N����b
A5T�3�Āph<��H��/�ʄ;�N�&>�hhpFi��0<)����7��%)�˟lv�K�'�!�d�)�$E@F�F�8BҁQ�	�&�Py���w���f�6Ly|���G�y�"��A��Y���G�˄σ+�M;���s��ܩV���^X��A�[B�v"O�0�`�}r.� F/�4�"��"O�E��G�"$}\��Ɍ'�p�iv�'��	S�إ���P(/�`p񅕪4	,C䉤3@����R5=~���%ȇ�?�C䉄c��캱�/�|��@�l�����.�	�8�Pd��ꃫx�'J�X��B��y�.��r&x:�� ��#E�B�ɗ^�(����4Ph��B_g�����>�+ƐN^�ѳ�@�XV�{��Ο|��I@�5�R�0W���f+5/zɄ�vJ�R���at��ѳ y	�8�	\���'1����ċ�@bPzR,�&]�h��	p�'��+�AY 5J�K C�h���$5<O��x�[�,I�M�D���T�'�Q�X;S!�l5R�2��h�^IqVE�kh<a�^.HE��V�V�l�RaHj��í]���?�2`�2
l��R���m;��p�j4D�x��O�#b5+���u@��A?���<��� &D�D�d�7,��A���v�<�5��<Y�(H�".+:tx(��B5��x2N��l�Q%K!I���U�p=Y�}R
�N��D��ϩ=)��{b�^*�y2�C�>�i��bս>��"+���y��f\J� pb�ꅲ2	V/�y��#`j�]��O3G���v���y��H8w�$��ٚΪh�����y���yS�Rg��4U��ru���yK�`�Pӫڨ�z��G��y�)@*rѢ�P�핥+3Bqb���y
� �Յ1��h� o�A� "O���R̎L�����M����Zf"O~�rD�U#a= {��5q��Lӱ"O��K�[�\=v�"��`�8b�"O�ᇅN�R@��W��~���k"OB� �V�h>��{d�����-
�"O����
��\	�f�R:{���#"O�;Eᙊ;�l�3)����=�S"O�!�`Ru#���s�'���(#"OvpQ�HG	Rь �oEka,\`�"O��� ��vv���(��G�H�!"O*y����v��g��2D\�a�"O������F�H��^�T̀��s"O>E
���j��Y��k�
� �9�"O�q	ĩ�H	R8@��U�|Kw"O,���Ғ=F�C�C�4N���"O6�H���(8�bX)R�E�W:z��6"O��@�`3Y����śB�Hd2�"OФ�(�`�����8��у""O�IK�i�I����D�J�8 a"Of�Ѓa�W�Є⍰�-c"OJI *�/(�6�rQ��A�xE�"O2��Cc�"R�ÒL̜Ai�"Ox�A�'�;�mڃM�O��Bp"O���)!��1R�,�5��h�	�'T\@jQ	��x,�yp�̯[KP�i�'$*��6d;`d�؈�	��Ot�ɸ
�'В,ʔK�����D�81J���B��\Q�#úEQ���d�ؤAF󄉞.�Z�(��_n�6F��:�!�d�	0j�R6aP�-��Ô�!򄋺^����N
"��%�����!򤖳��q��,A/�E)E[��!�d� �� j�Dgnr�%#��!򄘿\��ĸ��J�]\���8�!��	�B�"ªųPC��r��e�!�$!-ʆ�C�OL�~�vcbQV!�$X�;�6���.V�x>�����*}T!�d�;��XP�!�,X4@y�n�,Uz!�dŏT�1#j� &�X���`�!��_�l��v$Y�x��h��t�!��<��VJ�lP`�e۲gd!�d[[p���*q*(�+`�F�N�!�O�o�pӠ��Q�����4/��C�I/}�Լ��Α�L
�#���3PB�	�e"��(m�2aoR�F��C�	�*��H�*��9o>̀���T6@C�	
:����L����
��p�5f4D�@*�FV�~�1���z��>D��p�JڨF8`8�Ǝ6��Lp��3D�\�DNޘC^p���ŲCBNak0D����%��~AY!�!)�>�S��0D�p�E�I���1���M��=�f�*D��kC��/&Ċ��2I�1�eA�g+D�L9�#/Y?BC$�])uH��"�)D�t;$�K>$m@<k ����&"D�W͜�g%���bв}Z�yZ�k#D�H����3�v�	�D.rŪ �:D��Ӄ)ܟH~���B�M�H�ۡ)"D�B%��!^^�	���b�U
�%#D�`��߷YԶ�0��?+�=��4D�A����2D��фM2�[�/2D��Ps.ʥ!�2I��˘(TNMpCb1D�0�-�p�(�2�е�r��0-D�$#CJqT��HFB��wA0��r�1D�� @��� ��KV����#A�f��p"O� ��=���@7��8+_�[�"OJ���E�X�d� R@V�$q"O��s�TKD��x��ڲ`����"OT�ӡ�	]ʂ�"B&� ?��̻&"O�I�

 T��8��DX"O�)h��Ѭ ��EY4I�+p�H�10"Of�Q�D�r�sr R��r�'3�T���
�Xv��[|��� ��3�:��ad�^��D5L�5i�ߤK�R���Β���@8�I�$i��4�P�r\��K6���b)#D������+�|��ȓ0 b�)E{�z�� �5t����I0�XL�kW,Dsǎ���ȟ�e2(�&6���҉��+q�0ra�5D��Ck��Y`��¡�Gx�d�hи����%M0)��C�g�7S��g�'�0�'��sT�{B���*�2M��ܢ��λm�qY�ٽk����֠H��Y+�
L����_�o�|�g�(��! w���mgPD;Qǆ�(OnT9�gP���x��DhlDd��U��Ƒ36�W(��a��$�B�	�rP��3�!�-�"a��@M����-X��{4����8U��L���	'��ﮥ���.5$���G��A���B"O�Yt<��y
"�̶yA���1�A���#�%%o�P���	����O�؈7�@&y��U�@��J ���p>� ɀ������ѯN�Hp�U?���"��x
���t�ˇ�L�1�#_]����/ԘV�<d1��N5?Q|�Hw�1ʓuC�Ѷ��P�&PYrG�:Zh�p'���?QBv&ō~�B��g�Zd��/D���G"�J�\@�s�p�����L~'8�ԮĖ8��h���]S܀�'��p�ϿqK��P�� q[���7�V�<D�Om?���ԯI0e�o�1����]Lm�W���W�,�)�?��"*3�I',��R#Q5U�L���r����d�(�e��%O&�͈��V�6X�@�g�Ac���"�n�v!3�eK��M#rl��`�VL��X.ed�h��y�͡\�&�cE�.o�k7E�"�hO�pC#��
�JmyD+��D��i)ǈ
77�t}�&G�Y܈�T�0��y
�"iz��@�	N��ӡ/[Qx��kt+��,h>);�֚���X��|��Ҳf��`�r��pK�"�܅+��<��V����h�m��E����.;]U�m��i��LЎ�`�l�-��xBŅ���9����4m��z`.˨MYF�@�i��[T]�IN� ꦬ�4%E��%�ŠU4l��2Ў
+�y�剉��Y�敯4d��"G����?�%I	P&T���O�<*��౦���~q�#�´J��T��Ȉj�}ʧ�V<[<h�T7:&����f'��D83:h@�w �UЉ(�E�(eџ��a�>h9�BA�S�:��t.��v(b4S�@J�}���C4�0�T9_�e �x����A��3�P�ቧ6��%kኘ�)A�y�"BTeP�c6�QVi�	JN�91	�&z�H�j��g���������t��
�H]�= �`�%*,s0B[9�L)��'f�)q���!�ҙ	3��9}$��s�f^� �F)�`J\4����Y?vi��$�	�މ	s,�y/���wH={ՎR-`��Z���r �8S��uB!;Ul�  ,<�����3�I���?B��"���O�u�O�?�&�[�]�%'&��D)��5�}��O�Y9WCƘ����@8Peh�В�	�X8#r�K��Z��բ�nY��@b�ڐ5`��7+�)�|�-u��I���=@��EN�a�����)=O��q���E�Z}@���dq�5�c������Ѩc��3�gO�?�H��@�(��jVL���I���G�ĩ%,}���<)4(9��_�D�����zV��_�Z�b�M������j�? 6��H�q�Ψq)�.o���� � [�T�B�+M� ��Պ�jj�U[��W:$�(U%�H��zٻ!($���u�U>��4т/P��"D2���0O�LM��O(��3Q��Dv�1�4*��:�� �rϑ<�<x�OT�KE+]%|���� �Lz�����'����X�Ku���0��8S�Q
A=n�ҥX��/�ʴ
��&7�v��18���"��kX����)F�)-��P�Ň2Y ��ch/��ņ1^�ۓ�N�+�|��"�2QF@Pc偹>����I��� A�"S�G�����3':���-Ν�C�h�`BG��MR	��?��L�F�A�!{
���E�&܁��H׺ ��>Q)�8����\�+u��À�>�ĭ�6O2(ҡ�X�gf�i�7�]�3�"�oO�b�mHf؄y��S(M+f��8��ƙai�U�Ǳih
�Q���<A׫���P�1��W5̦\quos8��R�GX�]�v�%>
����pb[�w%j�D����A8"픊?���;�B�F�f<��,��MK���5p�T">AB���U�(�*V�	�F��賎�hy��ح'�IZ����l�Ԫ���2IЦ+���P�	�n�ԙ��:g�����4����LZ�t�K�'��p�����c���s��_N1�,�uF�Q���"P��@�E��T��ܺ+��{J4d�a޵�a�V�mb�$ pÆ�q�6\�f�8�O�Kac�l�? j��3.�:Й㷢_�D�a�ʇ�;�\雓!\�y&�A)�@ؤE�f�ңNT<=Υ��4)���t��ȴ�Ȥ�B� ��6��5p�.5����$A��F4�V�9!̙B!	H�~`��N	�<�6�S����M����ǡW)f㊼�3L�;?��8{~�>���;B��Tn�
	�ȻV�⟰�/ѐJ�xp�0@>n����GQ�D�%鄎�6�����#u��sL�|��d���G�4Ac���X�<�O�"G���q��t�a�rf����
dm�-"��
͑7+c�)��o#D����b.w�E��[�t$�a�tmsc,�"q�:I�a�Jx�X��H�BO@h��eL�\�3aR1;� {ceK
_�X�e����:)����20Y�X� �MY�$K��3��$A.^�i��D$c8��W�kJ4�=�@	Q�R}Jy��E�B��% [�
�� ��SM��W��t��HN�|"��D�vx��� G[�� ����{�U�$̦\����L�O,e�Α�L��\��-O�O��=�Dn�$|�i���%[�� �T���H�(�aQO�J�J��c��V�j����<D�hۗ`[��X�CbJ�*�R�
���{����l�;7/���«Ũaz� �35���]f�`��Nü��y������ڌ�p��GkM��Ȼ��<k�Ę`'�E=r#`��Z��0Q�ϝ�w�P�+B�$����a����µ �o��w(
\zQ��D�5�$�*��X�p�N��oE����X�f�]-"=S��W](�`���
2f&�1���y��!$$%Ad��U�Y�U��Q�ΣE~QJ�'��]���/\�a���W��e)�'�z����1���( o�#V�8�f��,�&L
s�K��"%���M��d�?,�r��cb�$,`� �"OD�aJ�:P�p���+�.X��VME+�&�K�+���``�h�J�"Q
s>���M�)H���=���فd�>53��,?�upB�'On�U"O/A-pi�lM�3�Ԉ@�V:&�ΓW�ܸsh���mYՃ®B*~Y��-(��}(edßjv ����rG�$D~���"�@�S���c������P�2|�Ueݲ^��pC�]K�����&XR�1�u��630�ͅH��E+T�a���B��V?	��˓P���#֋;Y�"`:��Ҩ{�F]9�L�?g��U�B�s� ��`kN�0�cɁ/wH�qh�u%pB�/=�bT��4_� ��@F&>��3xy�]˕
		m� ��-9�hX�/�2����	 �yw'��M,H����?(�h���J���x�闹{��Y*Td2s]6�b�-Q�+�f�ۇ��&BD>{GER�R�5т��9{��I$dSp�V?: ��/S/¬D�C�D�G.���	it�(W�ěX�hX�(�k�F��F@�b�~���']��&��h&m�7lO�u��!YPJD�p̘9cb�5����\13��5/
Vh�ꂂ�d��%{�� _���]9A�DA�E����2L�,K,NC��#dr �3�^�PD�#_w\!�gA�`��q��ߩ7]�a'��`u�#I~z�eq�i	���<(�وb�ޑ7`=�W+D�8�%�	/���0���3�~&��BeŗWJle�����>�nM���@)-_B\A��F�Smn�K5 Y�2δ��E�JV���	�1kne!AMR�R����Pc|���^,G�0��a��i�F֜)��9�2$�L؞��AU�crp��.X�+'d��A�9�I����x#l��-��!�Skُp�$uyQ0�L�	υ&dt�a��Ճ,��8�ì�F�!�DS�|H�}2pŎ*&�~areřn�:��W��X�K��"^D��f�S9}Jq��d��w�JX:7�] }X쨄j�T�f���'�>����j��:��G�L�4��M��8�>Y�6-.Dabx���	l�:�ÌE�'���PeY1T�0HR�dT�D��Pr��1Q%��.&��i�B��+���ɗ���X���Sq,��jYN��q~�����L���kO.
M\5���Ћ��8�=q%(��]}��b��Ztle0rJ�%T�Z�'�T��uC�}TF`�w�� ;������򌙢`NW����b��XbN9I@L�/�H	�ꊢ\"4�E&R�O`F�ɧ0W<���oM�R�3� 4vvB䉲��h�vB�x�̰.K!J�0s��Kl-R=��-͈v��I2��2�Q��R�+ɭ/� ��I�7Yn�+�L&\Oqr�������Q�,"�6�����%bf� % &n��!�%+|�P��I*X�j��ԉ;�~]��ۭD�pc�,�6�Q)X'�48�� W,�0�%eR�I��-v����M�\� ɩ߲
r!������6�:��}��ҏM:��k�h����5-�$� ����eN�1������>or(eB �:D���#�2�l��Nʀ;����ƈ�.�MS���nt�U! gܾ]��g�'��ܲըF�Jp�%��Y��U�B`l]�6��3�`}��Y 	����	X�jeV2z������� �x�0�^�RJ�"=AP�rC�a���R 1��!��ȥ)I�A� ˌJ��"g"O���a�dY!Dw�;g�'������J�B�O?u(���%N�x�K�9@�XL���P�<�ǘ
/!d1!w�ƞt��H��Q�<� ʽ#T�=B�����8v�18w"ORU�w��.��05��$Lj�I��"O�$��n�����lv�| �"O�ђ��	JF��s�L��"O�|[��+O �(��
��,O,0Z�"O�3�!ĳ2�d��N�&	*V��4"O(����,��@��I9>�Ԃ�"O�<Qw��%�Y�s��J����"O�q�R��4@��IpPN !���I�"Ori�w�+�}0�-�7)��iHr"O�]xԤ/1��xz�R:Uzܚ0"OH���)�Jf�E&	X]��G"O��hp-� '=�=k&�NB��	�"O�D��`���y�E*D�/���8T"Or�� �P�j�ه'H:u�h"O\�i"�	`;08�ƀ�],��&"O|�H ����X�rƄTr0�1"O�h�PǊ�8Aw�Be�iy�"O|�t��&�����;��'"O�(Ѣ␣zK^�qV��3r%��"O0m[��%(�\;���"��"OҨK����N�	��
Y"�h�U"O����ꊐV�6p��H�/!�=Xt"O��aA腞��Y8��U*$ܹ�"O�yI�d	)p�pQ����ā�&"O����^Q���i2&��=�s"O1��c i�(�
�U�NQL�c"O��0��Y�4]*o�JkƌjB"O����"J!f���"��}J,Ay#"O��Qn��4���ju@�2`4��"O��
�=I���!� ,I8�S@"OrX9"�ƜXb��`0o4-/6a�A"O���b�=a�Y�"Oh|�P܋Q����,��lX-�@"O�St���NrB݃*�:c�����"O�QSW�;
��lhj�l���K�"O�LzD�_�x-i�zO�P7"OAc�fÆh;x}��ٔo��Ts�"O����d?'MJZ��N����PQ"ONA�g�<'�na���	=�ލh�"O�	T�:O�0F��zG�M�"O���%��vf�yH���r8^ � "O ��F~+D�s7�@�|�rܲF"O�0a�������<4d@5��"O"�H-G�?@��%ũ=�4X(�"O�1!�� M�ZE�@�r��9q�"O�d��h�}�\h�#�^��Rv"O~�a�	�	4咡���!w�К�"O:�����8w�$��F

^,*�"OXp�r�� q"œe����r�"O�٣�������J�-�d��w"O�}3%jԛe��a�N�/a�S�"OZe�%d݈��%�7nǯ?���U"O�y9�ESn\�����k��X�Q"O�` qgӤ&xxP��,"�H�� "OZ�G�T��	vfаYX T�"OL=�'J���Qg�u_� �g"O��$�8DR�J���5UF��"O�x m=���)g��7�6i�"O:���≛�^�2ǡW��vջ2"O��S�,�<2���+vϟ !�|QqC"OX9�4.X6B؜AԎz},2��UL�<	V��5I.��9*����aH*D�Ȋ���\�Nm����u�P�y�+D�� V|�s��[xb!�v�k�H��"Od�
�	&P0 8��=kk�p�"O�\Q$G���n��Bc��(2"OTq� ɍ�fɴ��u��'^,��"O>���M�>y���4F�|J`"OД0�$Y:
�1����U0~�a4"O��c�ܼ(' �ʵ&̋`%py	r"O����-+v%�0��t�v*�"O�@(/�|lR�w����A"O��9p�[9S��;�&J$J�B,��"O:4(��Y0���%��Ǫ���"O�(��/����t��
Y.0"0�'�
�҃�ֿ7{�4��'B�6)�(8ӄ�>}��9k�G�#:| ���F��"Pơ��i���@�Z�lK��B�X(�0�Rv�\=�����Y��?F���s�� 	>D��+����a���kkh �Џ�|՜|��������F���d��M	'�ȟ��h#��u�� 4�"D(#�/D�` �,�2�z� ˊ�M�.�9ġȇϺ=9χ�����4@��g�'��mB4A[<L�,�R2*��h�	�dy(����F#j�]���߷/qD!���(Y0���'I��Y�b��<^�|r$F�=4Dj*	 �]�ݐ�(O��$�58?1@�
ۨ+�};��P��l�)��*3��/M8}cc�O�<�1��p�d��5�à��pB�R1�8�,ǫ_^ 8�� �!�<��q�0����WA�51�"i%Z�9hLau�*D��(�+ߕ%w`�I�L_�(D$Y4φ7��Ei�� ��9�p��B�r�S�96��*C�+�����0�B�#�O�lx�+����@���+Vh)�3_6?�l�BH���T�Ȳ�װ;t�u�S�'|�)��DܠyԾ)�'�B3P]+��Dմq{��q�#٤���
;^I3��O���@�p�jh$/�����S�'�ӗV�& �Ǝ~Vm�%/Ȼ^p�8u	Ò5f��80�ԥ[����������0���+�4<�c���<��7"O>@����i�>���%8��q	�Y�L)��k���x��
����	�\��OB�{į¾3ChY��ߺ�E� �'(���Ꭹu��1�˞lYt6�\+Zg�zU�ܘ$I`�{Q��6Fơ��4^�.��d��|-�Q�ᆈ�Ԙ'����,	�Qj�Ny)<����O0y*��2BkÃ~�D���'�`��ע*y�}u�ɝeţ^����w	�&RS���AP�S?+�'ΠD��&�^�\L%	�1v�9r�'iT]��U�%w.ѠBǰX���'�PT#E�0u� !B��
��:H�� ڧq�-�]�&� d��#$�L:7�M�(���#�1t'�� ���'u��(�2�ȑ?�HKwZ5�PG)�+���N�0w ��hCaiޅ��,�%������:Np�c�'�Ox�ȡ-p,%;%gP���#�&"�F��bR�Qv8a�N8cEIjBOş+2S��Q��f0?��c�,�b�
��%@�� B��A�'�p���Kաh��s� �C��`�+:3=�-[��+\�0Y9 (/%v�kc�0@�蜚�nR��<��B�'И-˅!A0Eؠ*���>���0.OeP�ň�zG#Y�`�dE �l�0�P�1 N�v6�uV<2
҉h�H���``�:{j��`=��k`�G�0��m���!^/��F��? �d�pc��_�
!�u?h�x��6��q�E�� ](����ov�����/l����O
< �l2�a7�Ot��Ŋ�_�!�Cʞ%(��%���S60-Z��3�?���݀ls !	��!T�˳*_�/���vG2?���1&�x���X9\����foU\�'�J���h�����h�H���,2e�* V����8�`���[Ǹ)6Lñg��	�`hϰ���[Q��SL#����d�X5w�:����-?��I�0i�U:�K�re�ړ��X��(�6Λ%�M3.�2A4�p���4I�FY�NA�^ɲ�2#���x���2I�P}k��
^6���4 �%����4.ԑ��ژO	�uI"���M�B]Sq"�^6���d��y'��z�4"@5S�>@����xB��gVd\#a
�S�p��ע��gLx�1�����Qz�-Ưy T�6d�dQvpC���$T�n�'�>�A�X�Py8�PքIĊ����.\��y��ْ%r� C�[�p�Q&�D��C�FA�����D�n� �i��2:KpXX ��L���<r88A�P�ڪl�D�S�ܮ���O@�c�$,���[wc�ʰ����E�"F�٢a�=p;>=S�H�#����Ti��F0�]�&�[sh<��EDH�r�btFG�{�̥�b�QZX��Ɇ�Ahj(�)�Z!���qe�K�v��O�t��r6�`RS뒮l�ur���8��%I#On��$��,c�y�&}��C�h"��yA�K�w�l�1g`�C��XR�	��AIY�-�ب�Ps&�3n�n�<���u(�[��i�",��/��ԉ)��ɥ$�y��mD'
�Z!�\%Ѐ`"2�P�k�B��� �D ��2�x�#)�8R���R�|��Q���*򉌇w'J�rs`�4<���[�jϮ!��T��]�16�K�V�hh�ʸ�!�$ˣVIʱ��B�<�,;DI��W�eD݈L!L��W��1E�V�+��
!RNơ�̟,�b��|�E�ag��25���7��B�2�/>4��G͓>�d�2�) ;Є�q`Y�z�,�c��w��T` #����q��;�z�JG�,�	�Q~�\J�b��)*ŉ��V���D�a��B5i[%QإAU�
�&1��q��-r�*�ŭ0�-�j+�̈��ޡ`��z��B�3�L\��kJ|�lC`c����}�`��Pp4�B�j��.����/��; @�!¬3Y0`�J	�� Ik.Y XD��'d� W�^7�`�@\I�T�:V��w��i	#�J���i�`r�87)�U���Q��j�h9��P��N���i�!#�����H�ll�Ɔ�3,�ѐ��N=\�6��dF�-n|,a�؎.��軅��K��ʙMЌ�=���L�p��vz�� �zx��f�G.srd����D�}�v}x�-"w#���B��%H0�p"��;@�|
�ظ.�A�Dc?\OhTk����l��Aj�[�*����9���?X�8Ȓ@c�m"�ɩb�T�O"v��uH-
2�Ɉ���}Qqg+U�N��BW=o C�I�����V)�$X���	zSyZ�I͏l:~|袪C6���藥P&��ؐv�?=!!�
�3t�1�̵"�L�B�n�K��{h<�L��=��<�G�[�h� ��[0h�p��s��~�-����o!�9�&�F�9��ѷ`�R�K��k$�O�0�"w#�O�8���I�N�<�b�C2I�"��$.�:X2p���,#~J<��ew��H��@

FIR���&q�ד R0yKGH�* �,�@Ő3���<�pE���Q�eR5q���Z@�
0_#P!P�n��uS�	Z��e�
�)���[w!�DU�C�J
��S ���6��SX){��"T�*!��N-o�H1��ղA�Nc>�q5�@hÐX�d�*#fE�]�@�(!"O�q��o?�HG���jܚU�\(�L�ئCw��4�`M,Z�-6��DxB��,K�$Q���?@qR̓Vl=��=$��=k���3'	_-H�����`(C�ؘ�3a@<M��Y�i
�$��Ȁ0�'/*��@�m��|�ЍYt�\c��� jhTL:�� �:�vM���Z1�����{�&�	6_�t�#A�g���N�s�<'��(� ��_��|��)q�4���"�� !���uD̽R�(S	)���Nޤ.�r���܈4� qؗL��!�dA8lV@)c�I�I�Ƞ�Q�-t����107K�&Jm���5�����2�ٙEHb���� ыu�Y�F�0Y0�#"*lO��[b�$�Th�W���4�8%��@G�@0���#k'���o�1��(�섢,a{���}�ʒm�42g��cCҸ'�@��Q�A+!Bܳ0�j6��Ac����j´�,$�ËV� yc֧��̆��"OVH�D"�1��`�C�)`���f���I/�,K H�5=?
�zF+�n@l�$�
q�S hs�N�	d'�9G���|�z�����3<|!�d� �@0��#A@��8HpN��y��E�.4ty4+�t��Lxd^�N�� W�~ϒXQvI� _p04����	��]������t�#���P\~P0�-$zS�a�6��heƇ'�R]�wE�x؞����
�C��oH��Z R1�>�ɉn+���o-@ZN ��H{H���������)�31 �S��L�;>��3��]!�DCL�d��1`"�ѡ���D�:0�T!O�F9�!{֢]���RT�C�Mq�X5�w�@�1�,#@uȠI�m��r�'̤E��ڋ~	b�5��1TԔ����J˼��g�G]�La�%H̠U���I�'VK@�E�8�q��#R��9p�O}��R(�,ce1�� (m)��Aæ�?1����a�9�"��"��6h����1�p�-9� ���O6�R �=ɲ�[�D"(p�h�d�f\�q�Y�/|��'s�R4ʔ�� a2�z ��!���(H�q���<<٠1%ޫn����'e�-� R�X��vAx�O����n�2���)/^X :�-�nC�51ch�!�"SQ�~��deͬt��A;#&�v'$�y��IY��蚵1`Q��� �X�g��c��ȿ_��H@�f=\Ox�W.6��1�BdfF��\�E���AW��3�f܉�UBf�݇�I�'��4���*Fn��Y�����c��bå�~�̛c��n��&Ik�I��?ܖ���̌H_��+ ֈc�!����N�	�7J܀1��ϐ7�<{��E��d33�� � qc��9	��`�Lu�Ã��D��,'D�\AS�ZP�[ ��2��U��M�p���y���&&� #��$�g�'��`A�ԇ\�<3�,F�B�B}���;�	�.2^���af�q4�2��l+�@�b�)���(7��y�㉕>n���"b-��'^,#=�R	��x�4�ф�߷Lb1�� X�2B��.Ƙ��%�3W`�"O$��u�9zn=�"�=$#V(��'V#��V�,j�K�O?]�e�B|>��W�Q��qB�z�<�cTrb�z�$Ɔ"�}s��q�<�e���]e(�Z�Y������F�<����� �
��G��;��#` �T�<I��}�t̊��T?�,T��b�~�<��c�"m��|pEI�>�i���G�<i À�B����|����7�y��)�b���uEJPӕᗖ:�����*as��*�;dϐ#�T�ȓBi����"�?=���BĀ�Wvd�ȓZ���F鏣sH�R�N������ȓP�A;�+�/��h6c��W:D��m�9`���A��X�(E/)r,h��V��q��=�F	��n��W�R��02� pi�.|`~1(c&�&J�Ć�S/�	�����|?>3�@��l�Tńȓ(�0��4.)!�\�[V�6�40�ȓ0����	ݨSƒ�: Ő�u�p��E�B(9�MӻO��*`���'lhQ��J�ĥ��ߝ8���Q�o�Q6���;�V�2%W�.��Y��k��*�*)�ȓb���*�� �������L�Ňȓ(*nQhdn�3��YZ��+�^��ȓ9���W�KJj�k�Ν�/u��A.%zg�Q;~��҂�7 A�A�ȓ���T�^|�h�
�|%����k��wF�dPU�J%M:���ȓ>[�!�t@�u��=(7��>H����M��)~����@y'E�ȓH�6��G.��f�n-�e(�	MrH�ȓx�p|��j�Hr�����p��x��i��]R�įC�Z�r1n�X��!���(�&�=^L,���l}{ (m�ȓ;&�T+Z�.@���$��漌F|�g�z�ty �+��XIG#]�y"Ι�?j�L��e�,�����~r�gfc��}�3MD�9Z�*sBĮC��D�v��;�F��5?�R�J���']��m�|�"T�d��a���Z*+�z8)�#՗ +@�I�|h�Ǔr>PyE��25D�����?�l���c��-��,{Acԙ�?�7��;k:��Ӳ�O�� ��B���eXt�L�����L���E��PY��M��u��u��ɡ i���83��i ���Q�� �#��wfP�-&��'�v���'��TC�2���MS
<-)�T���~B��h�P�aQ�|��	��q��	�F�8��pcG�кqk -g� 0i��ϓ�����!��ͨ�W%]����D(6��<����6��"|-����G�-ȕ�m͈<���I˖=���'xJ�k���0|z� ]$@���0��	V��#�E�<	���<�p���b��i>a�B#�T.��(W�#����r���y��r4�$8B�|����Q��M��$_�`�3�O�^���uϚ�(N�Q&�pG��&�X>���9An��#��Im�xH���A�	�[�Q>!�O+�aY�a�+���.� �����[V�ɀ���	L|j#�ڀ����ŨF�RM67	�!��ɯ�M#�D�q���a�~�K?Γ%��	��o����#��,[��mڿa��5j�mQ�~b���U��~�3ʺ��ea��f��F�9⢨�q`q�.��S��%?I�Q?O6��
(���@�a��2i��^%D�t��2-ލ�?a�'�PBdj'
��4G�K��b�� q:`�"f�_��y� ��~#T�;��А�� �\�H�Pj�2�Y�B�26��<�@��pϠ�<�~�sn��2x�CT �
?$�"jV}ң\"8T���y��	�$��;��V�3&j�;w+�_V���B�}ƶ�"f�|J?�������O��́&D�#T�jP��_A���A)��hC<JU�F� K�q�D���^������)��P����:q�C5�!���5��1�%I�1\�=��@�m�!�$ƕ�0H��N7_M`qX1�Y�t�!��ՏOW�P3 ���js�h%!�� d�Cюƽ�yv�	�[4�<��"O�U���7� !���>-
i6"O�\��/�b�aao�|�\��"O
�Hw ���{R���pJ )3"O,N֔pz��*�x9�g"O�����d|h�闭<4之�"O�����J�@}��'�.ƌ���"Ofh�'L�|�QB����س"OH�P�&\PT`CG�ס(�Ī�"O�t� �b勔ϗ�5/z��"O~pBpǔ�3��X���J��A��"O�hz�!Z$� �2J�1��Q9"O0���!��a@Z� c�B
)��#�"O*(� &��D<@��A_����"O
�"R?���J(_P0�*4���y-�u�
��,��Q>���D��y�9!|V%`�bF�H��$�y�f�~RL��C�f�D�g����y��V95K`j�g��.�HT���yB�T	K��)�6�{n�e0��R�y"뎈l�x�AXp�$�`PE�y�υKڤ�Z�z��* �'�y������ a�Z�pҢI��b��y�G9.Z5q�jVi�|
�
η�y,�	�BY2wLV�h��u���ք�yBAWO�v(VP��0y�*���y�H$�J%�֬BL��MP0��	�y2䒬M�<�	�'���b��nҊ�ybF����[`��#��<e!�y��Y�3=�t�Ȳ~�D��L<�yRȒcPh�w�,�h���$�y"���.h�)��¿nf�c��yҪ��W]��䇔+f_xc�.�1�y���d
�,v���d��x3�W��y�� ���q���&/~�("/:�y2	��y�؁�	ަr�29�q�\�yB�ۘw�8��1�ÝY��L��/F��y��^�\舃k�D��8���y��K+,\�����젰P@����y��ȗ+��U���*8���sW��*�y"��	�p8j
Ψ(��1����y2.��ka��Rԅ̀$����"���yB�5�&I�Ef[$� ���y�iI�-u`��Ɯ��<p��N��y�� vR���`Q%c]DE��J��y�`K/y(��iƠX�G����@b@"�y�&O����  ��Er�m	&<�y�)�0W��j�M�1b�M�f �yCH�x�`pA�i��[4d @����y�3�$���VP�#Ɨ�y����_� I�a�T�sN�\�BIA��y�C6^ژhR��/jX& �i�/�y�e���-`Ѓ��Uw�2q햿�y�eП=m�L�Q�ג`��|��@�5�yb��>E�!�3C��Z��-h�m��yGV�3+�	��H�=U�����y��O�bG�� �Q�49���y���l��ʃ����!��y�fܩ8\6����ۀ��x7���yb*�>���k� ��1ˑ�I��y�"��"$| 1Ǩ��(4dA���y�C(uS ]ے��UD<Xr`���y"J��e�iZ����NVF��	��yRa׈y�� ��[Fߚ��� ��y
� �B1�ױ� ؠQ� i��"OB c#F�j�R��܀VMƽ��"O�̉6 �
p��S�$Ïe4��B�"O�З
�#w��(�bÒ.Ph�	�"O&��a��/g>���`'�*F5���"O�Q�A`�\�Z\AǬŁJ0� �&"O�Q��A�8ׄ��M�l2V"O�� �)ڻ�11�P�G�$� �"OR��R	ܼ'�e�p"����7"O@@��kB!"�nly4��rŀMq!"O�:Qo��V��lB�*B�|誁"O�L�v`�0%<����� yT��A"O�m���H����%K�{���"O���AL���´�ӄ_�9W<0��"O��	t$�-.�\9DcC�Xt��8�"O<�r"����ܲ$gf]H"O�����Ձ4J�b �	�NP�(�"O���Ι3B~�JFI��!9�ek�"O��K��ԬtZ&�r	��Ez�y�"O�y`3�B�
 �%%Tv2%��"O,`WA	�;U !�_,y"�� "O�	�rF�2EZј$��(Y��K"O��+AH"\�bl[4hҦ@��̘g"O@�+�-�v
���	��Tf֩��"Ol�kv꛶[���Hӟa(.�B�%��z�Iי�e�% �>��C�GƆѳb�<o�@��`U'�*C�I�v�r�ӳ�6�,	&Jg�B�	�c5R�[s��P�^�Ӏ��CH�B�lZ�h�B��{e.D"�߈T��C�I+ָ@��K#/� �؇ _�xq�C�I/�R�%]�t����	^<�C�	"v_ I���(����4���Ui"C䉫p�h<I��H"�����2e�C�	���Ŏ�6D��@G�a�<��e"O^Yxƭ+���� k��m�!"O�d:iL1O5��ãI Z��"O(���`)JqXE�8󐴲�"O:U�'	Y�h���`�"ۘ�S6"Ov�H��O k�PP���n�D� E"O<TpU	X��HX�dB͓]�Z�"O�be/�	��2��úc�\LK@"O�|�b/Ch�ʔ�ԗKJ&"O����͂a߾��t�N04I,�ks"O������H:<Iz���QZ"A��"O �Z�^'6���`B�˝
1)JC"OH$q�E,}c��Y"l�:G:5�E"O�``Si��=`��"�Q7=�D;#"O�\9��/I|$��q�Q�@� 	�"O�R�aK6�	!e�c�v=��"O��Re#%e�%0A�U�.(�ڐ"O��H7�SE���#a�N) �*]�"O�h�R#�u'�� &��²��"O��bBI�mS� �0�	�"Ox�P#��T<�oO�n�P
G"O>��5EZ�_�l�;q �7'Z��р"O�}P��݊p�<<h3
�#oS��V"OZ���D�L�U�D	�j����"OZ�j��ǎ��!��1{���2"O��{��yjT��גSZ�b"O`���[[�H����p�f"O��*����^����1��9�"O�=��N]�����	��bx��kr"OH�,�Q�s�C�i�,e��_ b
!�� @ ���5z��6HA'{n���"On-�o�b�Z�؆�˶Na��`W"O,t�R�\�tMKd�T(cK,��e"O����p��Z&g�/K렩'"OB��",vİ F��S�r&"O�q	@�=���c1�ϫ�	!�"O���!���j$�*9�@�"OF@�u�V�v��{e�V�D4��r"OR,1rd��܀G  �F� ���"O~$[�$��o�D��MA(�f(��"O��ubǦL���S�`�f�3a"O�Y���7��q����]B"O�����0m�4	z4Ŕ����`"O����)w���Vdɴ!�jCc"O���E ����<h��H�F�Q$"O�Q�QcZ��u�0�9��$"O@�!�8P�
X3���R�.��"O���7��e���c�D�$�\�j�"O@��N��23�z��	lkR�!3"OP����*)P�Lܴ%3�Y˕"O�q`�Q0^8�2��&$��9�"O<,3��@�HȺJ��� z-i�"O0�8�F��O|0P�D�4iq�"OL}�󎖭����c�<e���"OHx�U�=i�H��!S0@7̹ �"O�%.΅�pI�>l���p-�>!�$��J�G�����
~�b-�ȓ�D=Pa%�W| �RR�1E����(�:e8@@L�2?�\J6-��%��هȓ1�0���[�0	����T�u�v��ȓZ�9
cm�R��i�"�2l�ȓWX��`���d�l��Q�w%���ȓQ����1�p8�T���!Vz�<��lw�J�ٲfճb}h̻�H�^�<�ǩ�0>�L�׬ӭq�* �e��V�<��LٳgH�Y�RP"z��iBS��S�<9�Ά�&��97j�*D�	e��I�<!6�H"@�hTzŇG�JN�Cf��C�<��o��l�|	�����]9�L�0��<�Dg�T�LQ��Q==O���j�y�<� Q�V�P�	�!^.&c�Ī���w�<��A�^�f�2B�[�h
��Xw�<A����q��%�.M��X��cK�<�h�Z����΅&E/X�5�_�<��") �&�F��"~�] 
FE�<�o���2�+X��J�C m�G�<q%���V���{���
R�ce`��<�ָ4��H� ��$g|5) iy�<ia4"@)���,����'�}�<yC�U�L�:����<(aIy�<Y�`�$��y�A�
!Q�$�BO�x�<auAƁF�X�K6�OB��s�EXI�<1�-�V(���^�d�ȉc�f�C�<��bH0<r\x�ϥ0	
���JB�<��o�%Y��)�Nއ"�x�p�Qr�<��Ød�2�����+�t]y��h�<��i�*�~a��/F9+�.y��h�<)s��/��l�䩉1P��Y��^�<!�e�>r�#,M$.�qɵ�o�<�FAO1h�X8+Tƍ'-ET��T	�k�<��C�t�*y��O�7I���d�f�<qĦ1v�^0�P�β/�tP�C_�<���*�8=/�&rw�l0kLY�<�6�!� �i���/$�;W��S�<� ��(WN�d�ƥJ�I���CE"OJq�d
 
  ��     �  Z  f   -+  h6  A  �I  �U  �`  g  Tm  �s  �y  6�  y�  ��   �  C�  ��  ʥ  �  P�  ��  Ҿ  �  ��  _�  ��  ��  (�  ~�  ��  �  �  � � 0 �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�	#��$x�R3e 	F�
�Z�Bړjaӕ"O�1RV�GF��УD1�HАa��E�Oԉ�
�]�|5����n��u��'6���½`���!�Ϸ\�~Aۓθ'��I��ܩy>TD�QD��@�0L�
�'#p1��sR��i��̖"n��P�}��)��v���s�_)�y`7Dϛ !���d2��C�(v��S�	/�	r�Q�"|2�M��&U���Y��dy:AD\|�<	#�'�@d�AIڣ��w�<�kc~H"vm&#���硓v�'#Q?u�B.��Z���f��|�  gN:D���RM��C�Ze���H!Z�\h��N,D�li���Mn��!�G�o68�	�)D�@���u\���a�+4�^�˕���M;���>YW�O~�>7�5?�O�eʅʥ,��@��؋�)XP<���t(�X�6f�R��H��9V�N�P,O����+�H�s�&GOCХf˜�
+a}2�>����08B�iZr����F�<��4;�1�L�"\��^D�<IsaA�B�@,�b$�9ۨ��#�D�<�U�\dppR7� SPel�V?9���S	=��H3s�i���6m��<btB�)� ���e�+�h=��M�G��	�'"O \{��G�%��iP��X�7�|%��"O�X@�����i���e�8�"O,\psΛ�L�nE����84% 	��"O��h��A5� ����P��×"Op�qW'՞/�.%�r��V嬰��*lOV�C�̍*x=�a`d -<����;O�=E�t��N��P��hҧf+`e!����y2*�)*�e�fI�[	�T��e���y��,k�,�Q��D+�t�Rp���y�Ȑ(����O���"0���yªA�/����$O*(��`�F��y�!��@�X�r��Tr&�߭�y��Q�.u����! �ö'��yrA�[`͹s`�2d��� �j��yB�>fd$0e��K?X���(��O�#~:�!Q�?��"CO$//b�b\p�<ن���P��a�4��8��KӁUl�<Y&IWX��5�W�/��c� Dl8�lGz�+۟[~��S/��Le�&,ٞ��'���'�>4r��1K�dR���T�
�'}ܹh�k��l\d�eB�?EF�b�m�g�<i��1"VlՋ��Z�=ѐI�ң`�<�ue�9��A��+ Х�"ˌZ�<�V��)�U �K'}�fi�bˀmyr�)ʧh��A����ÂED3B����n��@��;h&��q䐦K���ȓ^��\{�o�%Y���3�I�Qh��ȓ7�.�z��A��^���j@Wz�1��.�����6MY�
��P`ԭ��|�9�-��N�|p��M�Ԃ���.�@���A44���SdgȢ����=PuhW��	]r�:�(��B\l���@��Y�ť�qVLEC�_�b���6�Piӑ�ͣ&�B��a2�0=��n 	Zw ς����Z�}�X���lQ�PRj�:��<��"� ^�zńȓwb�A��FX&hF��Ak��I����W�đ�b��Z���aa�%-tH�ȓk�T�kǨǟS�4xq�G�
_lB�����S��6-��gې���WjH¤ku��.3�!��΢?Ҕ���)�dhp�)��,lazb�$T'=�帀�ضr��(Ǯ��<h!�D�_�lqP��(_H.i���_�DC!�E�r��LtoJp/6�[0,R�+�!�$И�@-��" k��1r()�!���*�8��IN5Zw�́2H�, 6!��J��,�#��Q�G}ԑ���ӞK �1O��ג}2�P��J��`�K����<���$�gY`�S�F�f�����!G�i0!�@�vS�}1����F �̱�a�i�!�Ay�tĉ1Tx�X�r�Ǌ�;�!�D�9'傈@�LC v��ܰ0f	�7�!���>�H�25�=>HH�'��!�$6����WL��D8L�*�$��K�1O�	�����Y�hJ�"dMj�S��I��p�C4D���b&�XR��fc�t�3A>D��I�S`�phF���j���bv�<D�(�7f�,H�v�1`⚅<��@w�:D��:@�"!��� ��'otq�>q���өLz�
�)ߚn ��U�q�C�ɶ|	�pP���R*Q%̒�TR�'�ИDyZ��'d����^�mBf�	1�I�,�hٸ
��~2���2j�q慗�
��b��y
� ��;��B-A;r��7Be>�-�p�����'(�S&\A��a��)�^��D ��^��B�"����%7�����O2�=�gÃ�&�,Ӂшv(r-(�	��y�(�Y���(��g�mJ�ǁ�yb�84��ѳG��4�b�PԮ��0<��d�kH���Eh��U_N�b`E0o�1O���$�&(�v��2�ϧ�z4s��\='�!�$�-n/�y�6����(E�m�!���%���Q�,˦��l
�n�Rn�� ����Ƌ�h�� dZ�M<~����ǪE!�Рw��Ҧ�(>ܫ�V�4[�1�D�a}���OB4�@���x�������0H��8gO�P� (�1}|�lk�@`At��`�4�$/�O�a���[7r1���MAppp�'�F��O6WȤ	3�����S������'@�L1b����cw���:��0Ox5*��Z8p0o�#0H�ZE�'p�'�~��r� �ct��@`NNCrXPxak�<�����. FfЃ4�<����TG��n�$:�$�i���OW>ͨc>�������x"��!�!I�	:��=1@��;(�(�����.f-A,�y��<ə'rZU0H>�'9�M K��r!Ď�eA��x���&O����$LO�=�H��[�	��h^�z��W�U~���$=ꓤ�	O̧ZղhZ���Cf���H�,B���H�I��Mㅨ�$)/��:���~]X��-t�<Ap��5x�j�����"
��j�m�'$ўʧ<h�s'ca% U(�d��m�h�<��K�8Z��� ��T��|����d�<10�W�o(:bŚ�.�H����V�<�G�Е[n<�b���+4`b���LX�<��
g�(z욫����i�W�<)U	��T)�X�/�0�Ub3��P�<���@�5�l�RM�r��R���T�<q�����R�GQ�(}xt���Y�<Yd ̧J���/�\���[g�JW�<�$��SuV�� ��H:�A�hI�<�&K\ {�P�q'�LJ��!v#�D�<��G�V��� p�ٱ<���3�%z�<yV�A�1�J��VJF(=�f� ��^�<)��=,<yp�%����Z�<��^.H�T���9kŎ�#��3T�Hh��;�D`r�,Z�R&�E� C-D���p'*a&��kX�|���D(D��8d��8q(zD Q�6�H��H%D���u �|�Bt�	!&ڨ1U�!D�����)lm��H�C�	r|��Ȅ<D��j#X�J7��� R�.-D�h�GY�)� ��R�_w"J��'D��HD� 3"�+��[s����*D��bÂ��Nj �+r+=r��{�)D��s��� ���w�� �@"D��1�!@]5�w�0����;B�IIô�A���r�`P����F��C�	�0�Ń��\�x����ӏ8H�C䉢1k�$��)�<92ݰ$I f��B�	�� �"Q�Q�����ZIRB�	=@�V\A���2xI�9$� 2 B�	�K�5z���/�h�uSl:�B�I2_��qa��&�b�h�Dևs�B�I�a�N�R��I�6)+�,�,�C�"M^a �#�0S��lVmGs�B�I�!�F���-׿S����bH�(4�ZB�I�=Π��+�5��u�ƨ��zB�)� p�0(�gV�	�c��_<�;0"O:�6��yK5�N�j����"O�������Y��v�R��H�r"O��J����Ŷ�f��a"O �j��nS��#G�L�i��'��'>"�'�b�'|��'���'��Ż�+�{��!�`D5Jp�){s�'���'9B�'�r�'�"�'E�'��4K���K�*�a���|����'���'/��'g��'GB�'�r�'�R8:@��W0�a�bνkH�Is��'�"�'sR�'x�'L��'*��'�b={a����}�!�r/��"�'�r�'z2�'3R�'���'^��'목{W,Фw0�T+!,���B�'���',��'I��'/��'B��'��]�!)�mD�=���#C�){3�'���'��'��',��'K��'�>\H��m�]�d�X�����'��'}��'w��'{�'��'�Ρ�`�Ϫv��A�.y�@1�Q�'Y��'�R�'r��'���'���'W~i���t��ŭ�>3V$�q��'Q��'�2�'.B�'��'\2�'_�8���5rd�����sd&�i��'12�'��'�B�'(��'nR�'?���An5Vv����S.tV�S��'�R�'#��'���'��'"�'����P�u*�ZA�ͷ?er����'!r�'��'9B�'���m�J���OƽA��%B �)��³fQ�)ǝ[y��'��)�3?Q��i���eM	�w�8� �ŉ{��d�m�,����צ�?�g?�޴v^H�!�%��1ڔ)��]�$Mh��iq2�5�a(�O�d��K�50�4[I?}��$M��e��i=��4B�A?�I��0�'��>�Pԍ�)v#�{"��zq��Ї
�M��Tc���Oh�6=�2qQAȗ$�乤b��Eˀ&Sן�l��<�/O�O�,h��@��yBNV)����LՉ$}|�T��y���~�X���G��I4ў�S���:jO$R�V8� c S�� (�me�@�'�'�7��X1OJ�р/�u���K4��yY@����$�I����O�7-b�T�'�~�"PC�"%�i3 �G ��@�O|�S��s�<`�I��pD�,�a��O�B3Ã+?t����_?c/�[V�<�)O���s�D��\�u�ƭ�WJ�9�@t���b�4[޴�L`�'�7�9�i>�q �&���o ��@c.�������	�u����q�$?��B0l��9p�:n�v��'"208��G9�![���p��[�%N"idl��n�_�i���j��r�E3�^��t��vL͛ď��R��j� �8[�H��Fۣs�@�3W��;)0*xk��*SX��+"ʓ�&A��N�E�� ���X�z�,���S�R����W��K�K-��I��J W��@�D�]�n�|`aT��\qg�N�=��I1�!E �T��M"��ʓYDVi��cI0:�B<��E��T�q��+Q���r��^^�A��H+)���\�#��eJ�B:b|Xqe��$2�xn���I͟\�S�?��	t���*���-@������;CN.�ثOn����.���%�4���O,�P���)6O�)!�nٺ,�*j�40k��C�i2�'�B�O����'b�'�h�-Ԧ5	L�bl΋x<x1��m�
 B� �O��O�	!�I�O6�PK���Y�Ûw҂���
YѦ9����X�IN�0ڴ�?����?!��?�;jhY��$��H��AD�0n��,�'Bˏ�<�ONb�' R�
I��i���PgDI�V�@6��O��;#c^æ��Ɵ��	k����	,1Z��7�վ����"͙"i�o:\���?Y���?����?���?��$��U�0TR��J�|ےP"e�O
Dśb�ik��'n��'C������O�K��� �H6�}��/�^@������	����Z�$L�x6�C��pC�|�p�G)�6,���lğ��ٟ$�	🼗'f������.�6�l���*۞R2�)qBa�T/�6�O&��O���E\��GU��7��OL�$�-e�hu�E�:�d��ؐJ�namZ��������'���SΓ�~�fb�$Xdo�&f�Vx�1N��M����?����?�E�%JǛ&�'�r�'��Ć�|�Z���V��P��œ�6��O˓�?�ե�?��Ay��Mk���1sb\!Q��D���C�Ԧ���d�1�V��M���?!���j�'�?�uL�� �NݲrH� a7���E�l���՟$�0&]��|��Py�O�'TWh��1�6���%Bӕ6�(o��S��Z�4�?���?q�'����?��r�X���ς.�n�i�AV�(A�Bùi�t���'$�'�ƠJ�O\�OQ�dj�?8E�E2g���
T
`�ٻq{07�O����Od�H�n��%�	��ԟL�i݉�e-O�?�����:B��EfrӪ�$�<Ѣ���<�O��'/r-Oa�@YS�DH�Xl�ɐ�]�L�B7-�OԜ���ݦ���֟,�����H���,7�`A�(�;1�ш�㏼8��M����?���?����)�tl�`
�0I�3U��Rn>p�"��p��6�'P��'9��~z-Op�D^#^dx�@H��G(�;�L�T�.���2O ���OV���O�$�O.��^�g���m�o�<��q#�LV��z֊�$76P�4�?����?��?�)O���	>��" �AYCH4}�g� G@:]�i��VP���'���V��P�i���'�4�����DX���y�~��KR��Ms���?������O��: 9�,�d���E_�[R�F��~i�A)xӞ�d�O
���O�� ����M�Iß��I�?������'�?��s�D��M+�����O6u�3��$�<��� "��b2U�ʴ!ҏVI�|3%�i"��'~&؃�Ei�.�D�OF�D�N���O������hDpw+��$���0+w}R�'���E�'fɧ�D�~""Z�ֆ� �k�5�*�cT�B����"$-�M;��?�������^�@��q���R!��E�"D.�nZ#!�"<E���'��ӆ/��}q����	��"i��Ht����O<���V[��&�h���!�� ��M�g�^i��o��R9���>!�JJF̓�?���?!�Ź�v�F/�>�^1��J(t�F�'�|Y��O2���O���;��ư¢Dޫ7<��a��w!��iV����/��ߟ��͟��'� s���u�0��w��^0�#�P�\Oj���O�Ohʓ8��H��$E
R�JP�s�VŠ��u��?Q���?)-O<A�惋�|�aG �+S�Հ7N߳u�|e���@X}��'z�|�^���T
�>����B���;PʰJ�JQ�Rg�S}��'`��'�	Wp4�N|b���)i-��4G�,SM�֩؛&�'��'剓d�c�l�͠Q���S��C��)�҃x�,��O(�C��=3����'���M�Q[T�:��߳n}HAx��҉B�2O��,���Fx��`x�$�/;��H��F�"86�q3�i�剂5
9��4##�SݟX����ă7�ZdxF�j� ȗ������P�8٥�$�S�'{ώ��l�rZ�<��T�8`z�oڿ\�����4�?	��?�'r��O���(Oii�Ń���73/���M��mca/�S�O��G�Cij-ɧgI�$N����W.!aT7��O����O��s�$Uj��?I�'T���Ϸ]������tA$X�}���4��'c��'7�F��	M���?��Y�7$�HdB6-�O��Y��q�	ӟ��	P�i�-I���@�
���V�I֩�f��>ᅭ�I��?a���?�(O��A�"�_���o�)N��0���ߙ!��$����ߟ�'��'���Z�y�f�	�FqD�(N�\��yr�'|��'i�I7D<����O�j4PI�Z&�D�t�+�E�O��$�O��O�ʓo�Z��'�\XP I$|����׀� �R-��Ol���O��D�<i �L��O�xQ��>5���#q�\�v����`i�
�$1��<���_��<�#�)آ���E�1�!gӴ�d�O˓Us�P�����'���+"<�>x�e.A�+0��I+Y, OTʓk��Dx������dU�d��:�֔�Mc��i��	�[Ǹ��4:���͟������ay�t��FZ��z5�C��5��&\�4�%<�S�'%�tlXr����!�^�Tn��(<p�Iڴ�?���?���_J�'B"aC:'�����(���l�7B6m
6��"|��v��r��&G�Ҡ�7���G���Jƶi���'�2�W-P�b���IH?�₟�)x,�����4V0h藬�X�6���<���?����}ZU`S�ˊXy�)1�Σ%(-m럀)`̎���'�b�|Zc����4l�ƨPR���<%Jt�O6�K'���Ov���O�o���G��J�x��.c�,���O���#���<y�+�0(z49�W��%&0�"�մW?^��<����?����[�m܎�̧2(�R��κV����n��E�n�$���~�	]y"�ٞ���^*�2M���!q�v�-P��ǟt�	�l�'��i�`A$��ʠt�P0�B[�>���CoT�^R9mʟ��IBy�X�8��=�',F8i�+ک3��IS�L�G&$�	�4�?y����dۛ-,L9&>	���?�iΎ�m�:�)�,Աj��lI�b���M{)O��8��4���4����
�S�c�']AHXj���M+/OxP���ꦡ)������
��'L� ��[�����6H2|��޴��������3��]X��a��T�{X!a��#ћ���
:��6-�OZ���OJ��KZ��ϟ��#H}ξ��#��4s�ՙ#��&�M[���2�����yR�'H�a�֡�1�D!R��2qE��s�ek�`���OB�$�OA*a%���I����I�N�<T�6��1q&ʭ��V 3� ��}� ��?�'�B�'4B�'�Iq3C��Z9np{���H�.-�la�`��@�U��m&���I�'���?@�tb�#ITH)� �2L���6�u�J>���?����򄟙_̩aψ<9�(t�Q�Y\RtxC��\�����k��sy�-kB$Cm�T�Z�AA�x�B�yB�'���'��	�k�=�O �K&��*Ĕ���DMv�V}�O����O��O�˓
�P��'��\9Տ��v������p��ᡫO����O��$�<�2��)��OSN��a�.+�q��N"WX�}��k�,�d!��<I���l�rl�ӴDHS�B�����:�:|n��`�	hy�"^�������,ճ1
�a_����#4r�~�PU�
i�	vy"ǅ�O�I��:2��q�V
*0��ơ�5Bh8n�����	�]�&l��4�?�/���i�u~"AإC��y㰌K�"�RQ7���M�,OP�r�)��8TzI򐄌Lf��W��?d��7͈�~ڝm�ԟ�	�S	�ē�?Q�+V�Qc�y *�[q�+�%3��A��O>�ɺ�� ���`��W�,I3���MX�h��iX��'kr犉
7dO����O.���p����D1n��x�"���YTc�|���*�	����	П�3ȡ&�4KE��0��p. -�M+��V�t�xb�'�B�|ZcD	��i�^������	w�� �O������O���OL�7��`B�J��s�RenF�`� �T��%��'��' �'��I�`1:���&%���"�.�8f2��C�(<�	�����h�'��u��aq>�P)�7�J��(L��$�g�>A��?�N>I-O^��_�pQ��BNZN��"�\�I"�(8��>���?A������oW��'>1����RŖ5���H:l���kb�C��M[������D
7�Oh<s��151~�Q-�l��;��i�r�'7�	*k[���J|���r�#.��ȑM@���@�qfO�:Љ'6剅w1�#<�O�hL:�[�C}b!�d<$��t��4���ȧt�x,mZ����OV��R~���i�x����<h �� �MS(O!IU�)��H�f�	d���(0����a�8kq^6M���nǟx��ܟx�%���?�4�X9n �I��͉e)��� CL�$��?�O>)��7I���L�����	E�=�V�iX��'Pb��-`#�O����Of�$�*op���̞C	��Jc)­%i��>9��Y��?���?�&C\�t�B��C�Y�P�5�E z�'���q�$4��O��d�Oz��S�
4i\�� ��	�Y���ny�O[̓�?���?a.Ox�8���bRy�fnH5]c i�%�Ē�'�$��џt�	jy��'G2��:٣&ᆤs]>��惛�U�(ܡ�y��'���'�4�H���OjL`� �h��ӣE?i0f0ȮO����O����<q��?�G��M�DŃ���հp
N>@��Y ����O��$�O ˓�]������:!�ƙs�ME��(1�7njP�ݴ�?YN>�(O������ם^����I�Wax4�cH,g@���'@�Z�|'Ϸ�ħ�?Y��^^\{я���P�0*V��TY��xb�'�&�:�O��`��Y��%
�!��t�A�1�J6��<	e�&����~�����֐�t���zl9sNP�{Z25���p�����ON	(qk�O^�O���5��H; ���p��di|�V�iS��Ht�t�$�O������&����U���	���I{R� ͼ:(۴Q��	���S�OR$X"aǴ0���0%��c��Bm:��'}��'
lU�&L8��ڟL��r<�:���6 ?��"c�K%�nG��=`Eh4pM|
���?������#l�;:۞$Y�S�i�
x��ia$�#s�b����X�i�Y��Ó ��%���0Y�lm(a+�>�1��<�-Op�$�Oȓ���Ȅ��!�̫vB�,�2��ݹz�
�&�l�I�T&�h�	�t��77�d���V�*&00a#M�u�bc�$�	ȟh�	Vy��������w2�=��@7�VѰ`h��EZ�ꓴ?!�����?)�%��ϓ��\���B;^�AZ䈟0L?*<�wW��������y��ɨOc�0|����ZL ��3�]�e[*=i3%Ϧ}�I@�	�x��Puܵ�	e��HU-\Z��7+����L�~���'�rU�X�B��ħ�?�']-�t�s+@����Q�a�?tq�\��x��'�b��}t"�|���쓓c�]��Dm�1遴is�	�
R��s�4H�S��������"D�0@T�2�U��U{�B�nZ��ɼE`���	I�)��<��B��`�칒ƉK9P7�$e=�Eo���t�	ǟ��S�ē�?I�)�U;9�v޴&E��Ń}A���[C���|����O�PA�ڝ,��u��LP�*�d��C�5�I�����K~�3N<���?��'�8���ʰT�i�eZ{9 H��4��9��H�6����'?�'0�0��8Vߜ8:5+ЮV����*u�n�d�u#�x�'���|Zc�,t�  ո+
nA�s��$6�l�i�O��E/�O"��?����?�,O�$��?�N���灝�� &�ޠn�m%���I�@'���	�p� f��`t,��GH51���j�՞+)t���cy��'@��'�剝y�DM��OE佸tC2?ވ�6�Qp<ؤ��O����O��O����O2���B����R�A3o�	�m��?t��fG�>A���?Q����d�;vMl�&>Mr0Q:HXM� ��#cR�:����MC�����?I��T��Lh���I)�qZ��׮Q�!��B�,
I�!	�	�:^�����U�^U6yo�`��~�08z<����vb�����H��yJO)xV���LsJ\��J]��С�gT~�ؐAW��/W� �!pK$cn�@'bi-��U��p�c5&��1��0x���眃 \>�¡�=���"��7'�i��d /�R�p�&T@x��3♉4tlP@�˽g[r�r�E	_�:t) �ѝx�P	��ɶ-g`� 6(�=U�E��X>R�'�R�'�P�}�D��&}L�Ea�>�*�!MH���#1!x��|ʁ@�$wzc>�o�5}i2执���&��@�6���_0���˅�W���7i�6J�!0�#����y�In���eN��5qr�U�R�0����m�֟��'f��	��|*��D�y���PB�?X���葬 c!���5)�({c	O�1y�4�CK��2���!�HO��O�S�? $�!%V�|�(��U���P�@�r�U�H:�I�t+�O����O|�d뺫��?�ON�!��E�A�n5iFc����MM�O6<b\[����Nޓe�џ��cO�E����$H�g�S�Ϯ':�1'��j(g�0�xGB��$x�4�(T�^$0!�1�,Y#�ċ��o����d�d�t:��D�>H3z�P�LOE��Z����y�Z42��e0t�_&.4��JEI��'���򄞼,���'���p(�����+��R��l6��'�0��'�b5��E#���(=�>%��X8�ѫTEH
tO�HrdJ�|�z�0Si��i4\�?���O�=�b�<E�tiI��ӈ3�r\�#.3>|��$χ<i�0Y��O,4���'��I8:�K'۔u�<��A��=m�c�����*�
קɁx�����Α!\�C�I��M�q!G�iL\ �ՠ"�A��<Y.O�$��Gͦ�����x�O�T�V�'� ��Aǣ*>��s�D�2�@���'p���Ll(�,Z��(�%�K9X��0艆哈:S��Ci�a%��B�&��?ײ�'���,@�b�}����Q���fj	b� \�O;8������(@#���tjDN��A��O��d"��6���[hṔŦFƢ�F�z}����y2�'c�y�T�vJt�G�]ج��V X'�0<���	�� x�O];C��cc�\�]�}(�4�?y��?��ϥPA��!��?a��?)��m6`�u��"jQ��"�q	H��dA.l>���>�h@�C`�v�g�;48��V�Q�b�J�>T���`�O�^�����+�qô��|2l��i���_*B��ʴn��9���'R,��L���,O��d}łb�ԯC~L1�'cC�I� ܈ �ԯ�t�������[<��r���˟p�'\�0�D5P弁��fH�-�Z��'��+���j��'T"�'�re}ݍ�I֟ϧ3���y��̓C2v�#�[6J��h�d݄g��xvE۳Lr���Ш3�(�֪�3��H�o�'4�Dd��Y�*�8����p=��b��a�n�gˋ'<1iC��+&�4����&� �I០�?!����x`�5>�Fk�
8�^E��fvP�� �PɂU�2�8y� �<�źiq�_��ǅ��M���?�ҊF�e�|(�´��������?���@�x����?i�OU^��7�ʤ:��B_�<9�*��\�
��b,j�+C��k8�d[`/\1#Hɂ.A��W��S�
!����	�a�l`��*~���ɬ�M�qR��5��']4a��n?D��]�!n��������?E�d%�Tʲ=��� Pl@p����x��l�b�[�C$<�p��9w���J��O�ʓ5�d�gZ���	c��cN�b<rEY�%����bD8a�TIZR�'0�Ui�f� uLU��cU �X�T>�OhN�P��!I���rE�
�U	���K� v,]D���i�	�Dc�|F�ī�6g���!F.8�@*%��:��	\p��D�O����O<�?��ҍ�$mâ�(�J
e�*eA�2�	ɟ�牔P�V�ār=�h��Қf=�����[�'$�qf��a>��a�(��AK<�8�`Bg���'���*`4>a��'G��'	Ab�Q���e�$i
H$�: k�Q)�FUZF�	�?y�(*PU�|&���ʜ"$�NEW��;�1W	�'�$�C"�P9E��)�MЅE�`�>����<����)C7��"�F6)�8i�$� jԛf�<��	ȟ�>���O��D%?@|�B��d�V]�֪s��B�,O��!0kʉ]WpA�� ��'��lD����S䟼�'��Y������@���
kĝ��ϕ	j,�p��'���'���~���I쟤̧~Kj���<-_�*�YdY,x��e,\�i���U�b�NMyϓ1D�`jɁ	Y��csjM5&B8�J�P�0���c�$6���
ϓP������s�j)�e�?j��TB���?������?�����'�F��o�)��чN�����q�'H������ԇ<q��yr�k���<Y��j^�f�'w�E�S*fY�+_�G6l-�'Kn���'�����'�;���p��  Qk��
�K�Zђ6M	���<�0�I�2u��kfNε��x���6"T�����F�*AᎣe}~��q��$<eNl�CC�4�@@��	�K����Ϧ�;�O ̢A�B�V@�&�{�U��:O��d�O��"|����G㆜{�oܒBtB�8�b�e<IS�i�<1;� �L�)��� ��%۞'J剗VxD;ߴ��|v����?9%�X�y)B43���|��Ę1�M/�?�����U��O���{6L�~N�fQ>ɔOU0��. mͮD��.X����N�ȁIQ�.;��  �G�2����4Qq&?��Ð�v����٧��L���6}�ID3�?i��s�O��O��]�%�_�F��E���*��y��'��yRAV�|$z��;#��Qjr��T6"?��i�67�5�� ���7�ցX0��*��ދO�fEm����I�	6��$"������՟�=� �\إ�֝y�Z���k�(Y�T��ō|5����j֟ �qGP��b>�Oz�S$��]�1������=Ð��74.�H����ȟ���Ի'�q��'���yDI5��룬�0�j{t�m���m͟�����>��?��&!/� X��pa6�"h�
��xb�̄O��x�+4!Bh�hԃ�����_�'�2�'�剌(��AO_~�i	�@B���/�����ş|�Iğ�IZwm��'? ',�`u��jɑN���̱�,�Ы�4�D��BK1LN6�՜uw�q�E�I�e+^�� ���hu�Q�EeP�iP#՟w3R,�͂�b��zWƋ�1T�Y �%����'u��/ʈ$-�q���Z�lI%Ky)��ğ�H<����?���&ї.�LTA&�ק4��	���y��)�W���#̇��!�%�v�,kM>�@�i$7�<���E����'��+�%��A�3��X�!����*�"�'��l���'u�>�0�����m�� ��22���H�!�x=�&��T�zE�BD��+�~����(O.=�	J�g���9ӧ�~E�@�1f��E �R��D�#Px�I G[��(O�y�6�'D�7�AI}�B]�-$�;��bn��!)��Ә'v��'$@-!�g��g;��Ju�؅�~���'۾6�I�0E�J�9vC�Yr`Ϣ_���<q-�0����'TW>=Z�FJП���L,_+��$�0���7�
ݟD�I��JH"�Y2s�*h5""�}�4[>�y�hٓ ��`rJ��^R���r�5}��ڦ�l��C�3<�̕R!#� ��ʄ��F�	]���E���O�zs�>����ޟp�	�d��}��{ƞ�)aB��BƄ#u���|̓�?Iϓ]��4�%'	DE�L	���J4bx��	��HO�a������a���:r��a�bN�O���>�O�$8���!]���a��H4��"O�T��״<Z��q�V"ĉj�"O� J��3z7���ӌ�Y��[�"O���o�#���Pd�A!D�~}�S"O�M�á�&{>���HZ(7�p-�T"O����*��#�r�Y���@�� ��"O���g�)Pt<��F"5}`�؇"O�հg��3Ξ=����B qp"O�}*C����>�ڣ��4g,�h�a"Ob����	蒤���=��T#"O�4�'0���$��4e��h;"O(m!s%���b��"O�1ADB���8����r��p6"O��`�|M��#���/���"O���j>Y����6Aw<��"O�d��J"B, 2ԫ
�j�9�#"O�H��J�?8�#@��LF���P"O6t;pJS.
�8z�F�f/,�p"O�����K�@�R΋�mD�(W"Oؕ:��5���i�&̗+�f"O�x�MF�eR8BE!L�T�G"O��"��A�q�pq�*�b����"O��v�	�TLSg�';t�"O4�9QcÌ>1\����[)/T�S�"O|ነ$��Ve4�XaF.hK�t:�"O$���L.��Pq��8b3|Z"OVmI�K�ix�aO� EB��"O�B�aW�"�FH� ��?%:-8@"O�]����2~<�1�	�fb�z�"OZ9�Ba�'90ph�"��Q�}�"O�C�ڊ=��2�o�?1'��c�"OB|��KԄ��䟪Z�,y3/�7Y�BEH�Z��ǒ�ws�3?����1���o�\�f˗-=�Q;��'(����'��(�rH��;fP���J�Jۖ�i������MXaF)o����e�z�Ĝp�ܴE���:@e�|
��R]�-X.]#B���bj�L�'{fQG���a�	��zx��OcĤ�'��,����¿G�\dzش43⥑��O�ԛ��W�G�ܴ�P,Rf+:�D�`�^��%l�Jl�@#�i�:!b�G�5�r�~nZ		;6a��I���l Qf�6>2���kƦ)3W(��B���DA��򄖍'�))m�;w�X���LA5��{t��\;��>աa��1)�,���kT�+�Eʇ��&`} ����?<F$�fhLD��u��@�!B�w�U9�Ł�w~�I�C��j�A�aH@�c�㟢� vxY� ri��0��������Sh墨��mɢ|�Ȥ#gG�˰�'�Nx�"��f��$QUD�g��K�'�5�p�ԟ��(&�Փ<�$�s�ӴY������)X�F��v)��/�r���� �����aD�-����!�����'�%�P�:7��M���4r�ŦO���� �%�义��P�D�j�C���V��hZ@�ޣy��mkĀ�"N��Dɣ%�v�	�%\T"|ⷌ�*��)Y�Mo�H#.���`h���t����qb���$��`i��5п�ƣ\e�X�)2��|w����>|JDS`��S1OJEQd�-������mB�@��h���Zz�P[A�D6*���ɑ�ˤ`~�6@ɷ_tta�''��Ss�R36֐���j�0L��<�rBS8��5ag��F�?!�Si�!~�{P픆0��0��\�(�Y�ǊI����F�if��imL+=��$�10{efA�<��'HaQ��-a���J������1*��4h1�M?��/�<W��PK@�Q�Vh1�eNE�'IȨ`T�V�=����%Y����8"�DءJ	���$V2�Ū�M�t��<+���]��i$���-_H��a	<Ke�@���
)��\��-#�A0*�t�"M.�P	 tnT9y���Rr�'z@����`�ƕ���=�Pt���䎢3��Eҳ�%>@|�z�� �ZYJ���hONl�f�0?u^�:$[�2^B� ���6LxI+�,��F)�ԛ�U�l�EP"@��r��k�f:扔2
�i�nJ�|Pd��K$e��	�e�4J� �@�D��� � ?����^� �2<�hQ�0��	�`x �X�B*Y�(鶇��~���jөR�1��횲.�X���ߏv*�s4�':p�X�
X��#��6et�P�$޹1P.!Ӈɓ���]�^��p�.l����D�":�l�HE6��a�)U0���2xa���Pl3�O�ق�]4|ͩ"'T/4{��"O�Ih 6���d�o��?��o,��ѕ'�<�*^�-����C�@�����s��ɶc�5&a�x�cX&,N0PR*þeW����(�A޴���'׬5�쨵��,_1��PdIB-:���'Ud������iӕg֪Z�v�XH<A�X�h�� !	Y'yX :��P�	�.�r�r��	@^���"Q�� �,+@G����'$��C BA�����ա	�\�;�HR��"`d@Z^���'H��1�m'*�, P.Y+|�X�(�)#�p��t����ش5Ȳ�3�U��]|RlY�'��؄ Ӆ�Vyu냄m��HѮ�2\�I��!+�<��Ћ��x=��Hz��x�͉- }�0��S}�D��u�sܓC��G�^�Z�p&�A/m
x�r�8����3�_0�v9ר�e�
u:UY�����$�����M�6�v�����?!L�K >�I(x	�c#�5����E��7KB�˚fh
@��D�*�tm�R�E��M[�]!h���Wm��M���q�8?Q��
=���jշiޛ&����I���8WĬ| #&�&��DB5xĸ b�8qQ4(H� �hO��*��i#zlҧJE�00 �G�H��.�
 `bH�e��\�p�'�y� ;z�&�6��@jv|ȴ�̛f��Se�-��x�)�>r��
.���l	w!����bjHS��YP?	%c6�$UG2�L�ԓ���� �l�� ��H%j��D�X:F8:<���d�
[%2��uB�e.)���NO樱W&%4�<Z� ��&Dk���{�PC��۰5Nb�PA��ːu��(�hR�vmN���O{��)���?pL�0�HT�j6��G`l���(sDDȤnè<�ƍ+��� _�́3�DL�l�6�Q?H���]�%Ipp(�j�??,"9�	��ЄY��2+����*���H�>��O�H\����� �Xm��V-9|�9��M�ʦ�"���ѫI<�~"��Z&=H�j|����ːR���i"\O��0`9�l��n�1v�"x���]�	x`�r��n��b���� =�>xy��ŏ��4Ԩ�2`�	�f"��H��\7A�N�G|��
��l=�DT�Y����"��)�y"�Фuᾍ+��Z�D<�j+�M������ք�2�;+�dȃ�I,��D$mT�J����|�0��d�ݻ?���L���x�K������<��i�{o��C��=/$����+-6�lC��̎�H�D�lo�]�(���רO��@W�9�,1ˠ Y$Q֜A�;OtT��P�D[w�58 &��OHJS��nvZ�:�ER+,+�(Q���ex�8��ɪk�T�N��v`�U��m�'�|�����l6Xh�M�K]��O6�'����N��d�>tE��K4O�y)hq���Y�p|Q��AS�L\≓a���Ʉ��x�$��%6mJ�L�?�|����L��TjÆ�yB�פW�'M$��OV�S�lƙ
�Bes��? ����v��
;*��:W�N�,�"��L��[n��"�hsfQ;M�C�ѩHM��"�)^�v��~2gV�k��pv���H���97���~R,��s�E P�ߙ)���7�L���)�)3Y���&'�)|-L�� @�&!�$O�p�`�2�����\��r@�	!s�&��)e��|�v;}"�·>ܞԛ��-��|ʶ%�5�p?�vŔK_�As&f�*T��A��kQ=u4���r��mY�"�_~,���V�? �Y���I�rT ��!"��ȱ�D��X��">)V� �D���6t`���<����;}��X���6)�6��a�L�j��s�>�O�33G=O�$��jXDzub�=OD���B���"֣�.^���O>��"�8�(��Ec5GQ8`Av9r�%ҩ#2���n�E�1���q�dP`�jg��Y�(���P���CJ>)��$���~Bm����,��I�*1�Lcvd���O�r낹��ɱi�l�)� ҽ�Ǎ�-	����k՘6.��ˇ�'\�ِ�i۬?�	�4���'+Ƶs��N^?�f@�yX��[�H�B@ ��O��<��MڝE
��'��
+O8�
 ?��I�PG,��PKA2|x��Hû
���J5�7�>���8�~�c7M�������g�����vS4 Gx>�N�@j�&ԣb�.�pvEB)��M*gh�V�B<(��'�؞w��J���?�=�V��,l$���hO1�����@�A1�\�c��	6���@�AǬ.X�p��9�k��;�N[�4��>.�<8͓�6��M�Y�.0��=�<�'q�'O:-�`�:v�f$�� 43��ei�'����U��֌�'J�@xFh��'�P�dݸ="��o��X���I>�O�!A�)3s ���E�/�Y��'"�:7��Iܔ��VG�e<� C��Ğ=T���J�!���0 O��G���A!!�Ę'0ў�sц�"PAJ�c�+���fE���) %%,O��������-+�ޜ�Ac�
?hչ�bK���`�'��	k?���ɶ6x�c�B�|Q��Yw�X�P��)��K��HOj�p�N�hE��9@$I}��c�O�Ty��Z��鰶�9M��ÁEE�s����+�	s$j���ʆ3f4x�6U���X9,���R�%T;��8�j��M+��S<?�*U��b:Y�Z�c�/�>�֩�?9�'D��ͮK%�x��Ⱥ&���/Q����ˏt��|�4!?	j�a�nǅ�hO���5
T-,^E�aY�M�ԥЁ�Z#@��ZM
��~RS>�$>u;�ǒ�;,�a�4d,h�pD_�#�,�����b8�����E0�yD۹byi�Γ�*�]rU'��?��'��T�xO�����3q�����og� �񫏠_��e�����hO[�4�ѹf�jׇ�z�d���
�<9�N�'a*�9D�ĈZ��Z����`y�D;����'��E;��CTH���K�e)�9�'�&�4�Jt�q��$��+:V�BI<�PcY2U�t���
�$b�Pˇ&�S?��O�)��nƔ*���:s"��- �,`���2InfM��؋s���9<O�j���%KD�9� �MRb*щv�L]�@L��s `��hO�
D�5�
M$☳mԩrL���i�!xc+��85ʥ�שz��̋�m2�?���?ձ�oN�.��x�E/pP�#vE�ܵ)wψWZy��	�s�"i��]�K�F����B���2 CE����8$��d��%�<�+O�e��-Y�j�2�S��^,���A��>�ѬKr�"����~��A���k~rM�n|��������t�E&A��*?��mJ4��^�K� ���!N���ԮT���$�Ph�o�����?.z�Ւ��	f���L+�h�ᦏJ��'~ў���K�h(��Q�
��Q�9	﬩�p��"�(���'2��X�;z�ư*4��2f��c"���Plbm�	K���O�bl�3d�}�e����?D��M�����@6��Gzf͞Jm���s��A&I���T ���5^ht�RD�0����M(U �a�'��b�X�NG�u'~���.�
@a����	*k�@R���0��� �h��7m�7������ك�S��Ix?�g?ihV]4�۴(�'N�c��O?�͆��9sF�?�~�	0i]K�'��P0b P13r��I2�a��-���e���a�䦜��Nl��IіZ���0/֊_�����&
l������iN�U?��!1�D0��Үf�rh��i����a��E�?E��"ע2.���AϗGT�Jw�D���'4� iǫʹ��&}�SI<��ɂ
O0���&_�I�0���C?y��U������҄&���@��]��+�\��R�^�^���瞱18��u�����@κ����N����w"�9�>���j��ʬ�O |���ŜC�ʔ[�ᆲTvN��%�$K�m�\ȢJ�$b�m��탹uⲥ�?1�F,�~I��xk<lSΚ�eu\ �凄k?J����Ӧqe�"=�;'K�%z����E�� a��=���3@�>-< �S���	��!��!D��Y�jXI��)>�� 0��	�rd1F���C2TԲ��;?yt	���;��	O�HlC�c��<���͝+���'R�ڂbגW�|qrHB
L/ܩ1�%R�.UȒ�˳�MK��u��e#D�΅J�2y{2� �禽����0rq����fZX�'��;	�~��+��)c��'���g�' �QC#�-�d�kE�ȁ�Bxcj�8u����E���� ����������qh 9@˄�Oh��Yѱi�|}�4]c8�|@��ߪN��-I�9@0��nß"�N��k��lI�a�!PLj��O����M�Wlĉ�eS>Y�r��3'a��Ann� ,�p־]������i����ɐ0Lལ��	-���"���-^��*�����'2�����_�$ARҏɬ$Ɉ��ab��7
��ȓxjP8�'*��e�y��D��8]h���E�
�(V䅴~ZD���6C�i��}��IS-�	<$��1t���|*a�ȓwx��`ڊXY��	酌Jn}�ȓn<��<�RQq���]�؅��\�F7Ny��)؇2�PD��S�? ^��o	$���DL,O6�`;1"O*ՃU�A�Ub\�;�k�5����"O�U��I>�0��*˪#�A(�"O��,[;e��;���}���*"O<����4}��/�H��$q$"O
m��R�	Ҏ����F05��9X"O&y����T�q��c�0m�<�F"OF��`'/,��=k�a�Zժu"O~�r��V�#�IH0��+3�J�yA"O�u�E�#x�i��H�&� Qd"O��+B��
R�	k�J�V Q"O`9Q��,	(����f����a"O�H���T�B墥�GZ�& �ak�"O�����^�z�jQ�5�&��A�"O֝�R��7H�NQ Ɖ��l{u"O:H��ЁY�ⴊ�*ż!�P���"O�a�DI~jD�It)�{�Z)0�"O��E�1��2')�������"O�̃R��>tވ`�����A�p�t"OT�J矊~N �P,6m��|�4"O:������p@�
ЖC{��z�"O$�u�Yİr�i�;_��U"OHՙ �߄.���cO5en����"Ob(����;F����͒jWL��s"O��0��Fi�{fFD�lp^���"O����&�6%�k�K-]{��� "O�@��K3�p:f%Q��4(� "O�C����x󤆀T��p�R"O�ȣ�MӪq2�ˀ�O!�B�z�"O�أ�I;~�>a�� ��^x�"O@��F���7��4�Yg���w"Ohщq
�<f���c��B�G��V"O�
�C�(^�:L� �_8��)�'"OH�A4q=IV��/_���A"O�U+��B#m�� ���Ǒmu�1��"OVё���?k �{Q�0n}����"OB���/ӡLV
	�d,�l��|d"ODD�2^d6��k�(�6�K"Ol��
�'��('��<�bu�b"O4�1��2}�8�0��
K����w"Od��NFE�V���Z�q�*8�r"OX�Qp!�/Yv�`B�Ċ�h���j�"OV����A5}"2�����,Q���g"O���P��.��Ig�C�8o�,�T"O6��E��T���Y��yT���"O @p���4���;a�|�����"O 0�))7ॢ��ؠ'�"E
�"O�4���X�s��|;c��,2y��S�"O֤��+(���S�,�Y��#"O��2TE�!��t��}Q��"O$�����S�>-2��Hb0UIs"O����:�&
p"�)b8���"Ox�1F[mȺ�B�O�taz���"O�ə�
�-M���!8�с"O���B�ܴ���%�9-Bܚ"O�T��J��ilf̚���%V,���!"OTT"�OҤ+��� 'a5D�	hp"Of�eF�9�0G��AмsD"O���
*��`���#ꨈ�"O���r�m��ʋR�F�I�-�M�!��5��"a�?H� ��k�l�!�۷�4�c�,�-<ޔ�� h�!�$��+��X�p`C�.��6�0(�!򄙜H�:���a� 0�h�Iç};!�� Fy�'ʀ
�Z�k��ܻii$��"O2a�!޴M���bu ���1(�"O�0�Sn}�|���אw�h[�'5^m0�`��c.��K'��L��	�'�b�憥[G�y�eM�*�0�	�'�`�[���O)�tZ�A�Qx��@�'����2�аhL��@�+��D�V ��' 
Ta!(ޥP$0�(!J�:u���'̪�*
\5��
�� EbQ���$&�]�	� A�o	�/=�������-r�Q������$i�
���'
ў"}`.l�<ձgO�N�9��&D���`m�9������A,�m�f'D�L ���"_�%�'�P�l�bM3D�L��eQ��(	ɤg	7R�"!xac-D�(���� W# ��oǺL���r�*D���`��j�EgW�T��(D���hA*Y�Ԛ�,ң#�*���%D�0�'@��rv~UY䣐7
:)�(D������I"gmR��
���*O�0yugS|ܥp焲o��D"O�]�Af�J&Z�ruo�uKt)��"O�j"���hS�2:)^��"O�Ye!�\f	���ԛ\�N�h'"O<2Vn��c߾-[Ŏ�9M>:���"O���D�$�@l��C�;&�ZD"O���Dl"Y��L0�N	8$��d"Oh����P�pr��!/Z[�"ODLYׂ�ƺT0�d�%N��x�"O���I΍�`T�4��cִ��"O�q�P>#y$uAŝh���9!"O��֤S#O	tU@Ԡ�{/���"OT�w�C�l`t��W�h#�5Y�"O��a��%���� M�4 ���u"Ob�X��<��;�/� ���%"O�h`�l��PD�A*`�i�수�"O�Y��O �.�����E�@�� +W"O&��\۴�SB�Lz�Y�$"O�ȫq�K�*`��s�� m�6M�W"Oܰ���ly�y�%kAC5h`��"O�pK7`�9L �Y�6)�Q4윺U"O}�1���^���:ࡔ�,����"O�m�7O�1�M(Í8S�Z�y "O,Ѫb,���zq�p��)��3a"O�`35eŞM�����Ljlx�iU"O�����YJ<dÃ%Q\u����"O@xz���-.�đq�f�#~}��J�"O��!�/��1�NAI0�C�'nr ��"O`�X1�S
�dY!� v`PāF�'�1OH����T-����bu���Ѥ�9D��b��ͽ��l���%��)2�8D����K�b,]zUl�T�-x�"D����kȯM����޿�PȖ) D�,��ϙo��@yp��W�X��84�؊�-��at�	[ԇ˦h��	� ^m�<�"��Q6 U�g%�z���^q�<%�U#/�u���ĩYa�Hs׌�ꦽ���!A'�Mu �V���*k�Ąȓ&?�$�f
M�TF����Q3/":I�ȓ9�*���	�p��y�!���}�ȓz0�I���·rN�b�#M�ޱ��(L5Yp�><Nh�ء.Y���D �E/B��u��I})la�ȓlX���(H���P�s�ͬ�% <D�� n��AC�2N�����	4���0�"O&d�B����qˣ+B�z��"OjT�v�-m�����B�7��=:�"OD�
I	'�* ��(N *���X�"ON��&�2���J�'m�H�´"O�g-J�	i6������\��"O�	:�!�m�T0���.�=��"Ox� � X�G�.����� (���07"O�0�U���}�P�B�V1H ����"OR�X���(G��! ����2��	��<�5�ψ^�Y�t�O�t{��� Gk�<'�_��<Qr�[���EQ�g���xrևHAڬ��Z�n����F/�yҩ��4�z�
���U��1�ADN��y���9I��s�&B�� ���y2L�!`a2p��(N��-C�Ɏ*ÄC�I$m�n��D)�:\�k4�*C䉞I����&��.��UPRj�#5��B�I�>��h��h�C���Z��B�j�B䉔�����논S��1y��A<.��C�I���h���^  �R=0Dy,C�ɌQ.�XYr��:��`���dB�	�6^9�/[�|*]��r���0D������.2����1��� �/X�!�=�\��R,1r�� n"z]!�D�}C(P�l�=�##��1!�D¿�u)Tm/7�.�d��8'!���5�tH�b_-4ʘ�Y�.�	N�ē:��4�3���{|���`,@+c�̡�ȓXwr���K�c�������/(���ȓ�hM�7#ĝi6�[I�/2��݄����#)�%z<@�c�E6��ȓb8���A��M��y�eL'o=L��Ih���#�&!�B1�`�#� �ȓ%jƉ�S/ъd��9��֟a��l�ȓ"49yPB��m҂��Y0zE��o)Ll�tҢg V���k ��ڭ�ȓ.HP�yV	!xˎ�h�RG4�%�E{��4�קP�*�ڴ��>,xȍR���ybb]S'�-�b����R���D%�S�O�"�ⴍR���u ���ZXJ�'Q��9��/r�z���.E�2���'��b*VϺ-;�e�)
�'�H��	zR&񩷌��~q��8	�'�P��AM�B���DLS/x��Ѹ���<�(xj�I�Y��r�I�R�����t�p������I�h�(o�:�8�'�R)��$P-zF8���8�:�R
�'�0A�{l�}�a%�C�8
�'0��HB�]�h�`qo�>,�x�ʓ%zti{�#�3a-�,��)p�z)���?A�K`}8�cǨ�-X��]22f~�<�D�^9��ѡ$��.q7��*@�<�'��Cs�����./����MA�<1��9[���^�	���� A�<ц��9{�
�
��c�0P0�.	g�<��#g�P!fGݴqD�=h G�c�<	U��MFBD�6B/B�Ƀ��NF�<ᆉ[/;>]��FJ'<M`q�g�A�<�`bJ=c��"�F�.<U�D�G��e�<��դ J�<�d�+-?f�q�Y_�<r�wF c��O�:�����'�W�<�s��EX�wnɕe[��p�FS�<q�L��,�E�:}�w[P�<� ���lK�5��Q5�&_�����"OZ�����O�T94��I����"Oz4�&d*\$�i�,Zfp��"O�a���@�>��1c�@�]ұb"O���G��K�i�4AL��P"O��!�˥NY{�)�:r��}��"O�����.�H�A����W�"O�E3�
��~�jG-�5��"Oq Q	�K�� ��l��f��m�"On�B�Mѿhw~��@��w���P"O�,��Cғi�(I�h�?L�|Ы�"O�Y!Q��"���i�e��z���"O����gՅQ�`�������Yk�"Or���&�H�
q"D����"OB��-K��3u@��e�s�"O��[`��7�M��O�7��Բ"Ob8��[�9"�KQ�٨#~2��a"O���i;(G����!up��z"O���p�B�������7J�~Y��"O±����B�Z�(%�[8D�x��"OH�e)�K(��"զE�V�ۇ"Oa�6� 7^O4xk�!цv��!��c�ҵ��:\�Kw䟋!�D��j�t�r�S1AIÒ��:w!��,UJN�A�KG�=FpW>VT!�$^�P���Co�)r���� �me!��'&@�y�kIT�h��Y�K!�+�b(Jb8#�4+P';k!�$�6#�{��q*�.	i��U�<Q��ξO�N�C�f[({�5	QR�<�udY�K��0*
"���z���O�<��(�yN�d��O��Y��mIH�<A3(�����yc����G�<	����N�Zv�+ژ)k�m[�<��kM.y���Q�Fu(,[F�X�<��AB:/�"؋�JҿR���uC�V�<�mV�3�dM��G�v�9���P�<yw�_!{�Z�qT�M�}z~	I�!�w�<	��RF`���D�SKnhK���w�<لK���b%�[�eMڄ��-�X�<)�(�c(��f+$z� �)�n�<�̂
3~�@�!�tpi� $�~�<�ʘ�I��A�J �� b���r�<)�ɐ�0�le�I�K J��&��H�<� hDp�(�pr�*'� ��(�o�<�2��#lİ��$�u��3e��j�<A�i�q�� F
!<6!`���e�<i i�c.P1��C�/��-Pa�RX�<!���F�Q����>���TVP�<�H ��Θq[/MIt��&�I�<a�EQ�C��i�� *Fqk�"XI�<�u�M�+�@u�7b��#�R]+挂}�<	��G)�̀9"��^�`�� _Q�<��T��4�����	!I $�Q�<"+D -��9���.N����,�X�<�"�Ϯb�vD���"[T���AJ�<	�lͼ<)�8㌝f|�e�0Fm�<�å�A�`��G�Y�	W�1��Ml�<ad"�y��m��BC
K�F`@��S^�<q�%L�0/@ԚS�څV�xP�&�X�<1�D�)����Un��7<��e�}�<���^�-�����̴n\,��Fc�<It�U1T	;�a8��X��U�<�0"����uaF�z�ԥ����R�<� �T!'̮��y)��D��Z5"O�jq�W3vS�R��o�y8T"O�,hr�̙~ɒX��ʍ��Պ�"O�@��"��^��M1�)��M��"O�����hW�ɫ��W&H���"O4Ad�
�f� v�<Jj] �"O�c��E?�P0j�R�V4X�
T"O"ܛ ��#	l��v���P"Ή�"O�9Юvh�S�
3(�S"OT��v!ݥIal]�&��	 A�"OP|�D���M��"��*�Z1��"O�@�H��PbB����A�"O&D)E��tnBx3P���}�����"O@�AJ	A������?r��M��"O��ъ���f�oZ���!�"O X�p+�0J�������`e��"O@ ��K���	�ŋ��G��!��"O�ԙd��1Z3�I�2.�RL� "Od�:[9���֎�D�$�b�"OlA4]h<�oU'F�4��P"O0MY���2g��<�f��Q���Qw"O���M�>¾��vi�|t5R6"O��R�+c,�0�Y�Z|�q"O����l�M+�,���M>�Q��"O�0�Ťo����� �4�-�"O2�Z�́o[��z�@����"O�����@vY�l�� ��A�L�Д"Oj�0#<P���ҫ.� �"OJu�� �/� �sa*	QN���"O�	a$ҮY��<��'��>��9�b"O�M��g[7G��g���?�q)a"O^p[ǫ	*�9j�ƙ��P�"O��-��be���H�L�7"Oz�
���8O<��Ad��1^�	'"OԌ	�A �5:��?Nv6��"O�l0s��F���R�煃U`ZD�"O�����N�50��f�J�B�Y4"O4���$�z�0�Z&�T1�"O~��q]d��y��,?{
=��"OjPG6(�걇���K�"O��8�����Oߣ�R!"O �(����2�H-��NϠ,�����"O�9E��7?hf$� �ߧ=��p �"O|�i��i$�*��@'l��h�b"O�$
�!`Z��R��V`}:�3&"O���g�TN\>�ZwO0R��u�U"O�@w�6@���.�%)�p�[t"O����FC�B9��p+��q�8�v"O<�2�+��kxMSA
Z�
���"O:�(q�	(g];r)J�X͸h˴"O�T��G�p,�5ȅ�;��a1�"OJ�ѡOіwIha�gɁ�~ �"O����F�.o��eM]}�@ۄ"O�b��א"�L���P`�"O�X�F狾B4����ݥHV�U"�"O��
E���,+�c��R�v2�<2"O�T��HؾZ8�Rϝ�m���f"O�I��E\0Rp�ѷ��>r$��Q"O.<Ј�[DT������o�EI�"O� ����?�� �ʒh6��hw"O �*�� �[)�ay����qE�4�"O�LB�cU�z�L�U���s�̔"OZ��d̗<C�%�6��/:�z�"O��8�b�1��82�S�J0��K�"O� LmҴm���^�+�n˃.�hc�"OT!�߽k~V�0�g(&q�"O���W-+qp�����6<�k "Oj$�����Ju`0�zu"O� ���N��QKc,��U��*4"O�I�L�&X�P%����`��$��"O"a�cɶ�J�
�-��m��"O���M�,\�@�S�[��r\A"O�ݑ#j���vLh�FۮV6ƀ�"O��u@6v(j��T.g.XI��"O6�
��J�V��}��e=iw
	+ "O`��ëϫo��౔i\V\�͑�"O���rфwV��r�C"5J��4"O����@\�Rq�8%i9'X��sv"O4�8𡙅o�d<w-�2fe��"O�`*E�1Zf�MZd�%{N|Q!�"O^��Aj�?sVa��D�._6HS"OP1�vG�()�T�A��I	��b"O�h �EE�X�T���B��[⡻S"OP}
��N�Sc�a�C*?�@�P"O`D;R-�@> 0�ĂH�:!"Oh��&jϞ[��@�ve�9v<B1"O`�9�cXv��d���9��1"OX�yƬ1��-;�U(�p�P�"O�0��.x��cW��#��:w"O�p!V��4R���0��<1�V��V"O�����!�Ն8���8v�޳�y��y}���NQ���Iu:�y�AZ,_,B� �&$�|��ʍ<�yR�s
�L�v����q����yr(�s�Y21��}V~�1����yF�26Y���z�`CcO�y�ND;b�,���cK�x�͈rl�'�y��3O��!M�L��邡���yr���r��RB��Ķ]�����y2�3J�DM�Fl޲��M�rI��y�
�
��kƁ�~��ӡ����y�hA��9���~F���E��y��X(<x� 8�螅EY�e.��y���J�l2s��m�> ��EU$�y�	�N��Ӈ�5{~����yEH����yB�S�?��(�O��yB��W��ms��R�d�p���ѕ�yC ^,�\��̍�-J��<�y҃_�l���@X�2� h�!�4�y�d�����$��_�ea�ѹ�y�ϑW;\5����*#VX1E��y�O�<T�-b��=&�n���y���p�2(���/$��� ��y�h L�0������ >w�t�ȓC�Fa�*܏R<4xp�A�N�݇ȓ/���ON	f�J�@���{|Π��� t�S��* ��i e��r���������>U������8 H�ȓ�8�
a8j���H1-ߞJ ����|����aJ�]s�t+l@���ȓOHX=z j��jK�8`��R�he�ȓd�$����Q5\�=Q��O�8D�ȓ���g�Q�J��|@N�n���ȓw�vu0���<XH1�ƍS�h	����0gŗ�7_&\{����f���Q8t؆i�7��|a(�5)��ȓf�-�rF��I�q�%M2���ȓ)O2�a��Q�X�rRd^�FAҽ��S�? ���ȅ�!C|��עL�>R�"On��Ԭ
*k�a�4k4b��i�"O��臇P
�Z�iJq}r���"O�-kR��n���0bJ�|�d#"O�hȅ���-40���U>#�$�e"O^�!6��l�ӢՔx���F"O�ڧC�#a��혶�]�@�赙�"Oر�sW�6�T��,�Dp�"O"�Z��F��G�:2����"O2(��ln���<�E�t"OJ��M�u�ա�G$%̼Y3"On�ᧀ��gy:�0%�G-BͰ���"O��Ceې=6̻���/g��""O�1F�\z �,���	N���"On!&��7�R���O9��g"O��X�TF����m�!M>ܴR�"O��Z�D�Pn����/Yr�J�"OPI�u�bi�c���:��@3G�y)�>ds ��t��?�ܙǝ��y��m��,�F��'@x]��MH:�yb@0#.����%{����yI4ˤ��j=e��1�r,��y���.w� 4ж���1�:]��y�h p������$:t��%Q�y�EE-l%t)�R�ȡ9�~]a�P�y`ײ0f�iZg�� 6��)ԨV��y��ˌl t0�_#,v�x{#l�?�y�$BJ�H,�vĊ&8~�����ybCZ����k�*�&&P��n�$�y���''�|�3	&�:�Q�O��y�IH�\�\!����# ��y��(�y�(�=�6,�b葑"�Zd�W`�y��\C���6N,�5�f���y�Ð�(��}�ƄL;a��H���y�k�+/�`�� ��_GXu����y+6<�����玩J)�DKI��ycɰ�j��3)�.F�~��c��yR�ˆ(릡���<i�����yB�̈́c��IS��@�P�P4�/�y�CD��{��	�3�b����y���2N��8hr�(�"�B��)�yb���)Cg�)��E�"����yLWa��q���%��)"j�-�y�FG�r6�!��O��#m���JǨ�y�
�q��`G�ԝG��� !�μ�y2�M4h�`�ʇ@Mm̙�����y҇�CO ��Շ�
=�$mpg���y��̺[�ب����9�� ��@#�y���t�H�si�!"�e�6뛜�y���|aqlZ�&�V�Ss+��y��B(Ҡ���
u��C�V.�yBˎ7x�j����(L����]��yb.�,"��p�l^�{i���Z��yGE"PuJ}�'�,t[F�*d#�$�y�J1[��͙CM;hE�t��X��yB˟e^��Fc�={�-�#KD��yB�\-�L�D�Ĩt�J�ό��y�M��$z��;V��o���r�W!�y¨ ~=��Etv���aY��y���;`*f��.�+p�F 9��Ǯ�yI�6*t�Y����" ����=�ybǦ!ǞxR�#ʕ�E��yR�O4�b-jD&}@�� !O�9�y�ɄfԆ����*r� ���!��y
� H�0��^�<;h5���W�'#|%"OvMR�ƴ���.FAl�(��"O8��w��,���zrρ*vx�|R�"O�p�r,��Kj��"da��'xt�2"O���׋[�C�pAFnQaY��y�"O��h��MuT:��� y���G"Ov$���ĂB.X`�C�7P9�,�P"O�=���#9��=#�=�4��#"O�
��;��ab�ɘ;��<�P"OH҇�߆O�������R��\b�"Of��ѫk8����\���P"O&�r�mL"	�~�sW旯&�Nɒ�"O*�!�g��6r����e�� i�"O숈!!C4*7(�Z%�	߆�j�"O¼Y��E-~ 	Ǥ�@޶e+�"O����_S~ݰw^,Ͱl��"O���V��"��!W���t]Z "O�� Ї��-� �+7�O�N��`��"O�c!�A�5`���(^qv"O��#e��	�~�yP�Ģr�5)�"O���6����p�ځwCB�B"O�ur�/˸Mv��3L��� �"O��%oQw�
���
ҝ?�00 �"O���"�X�w������8��iu"OQ B�1FXZ�k��*����"OfH!���Ba)j�U���1�"O��a�)�C��h7	�A�$i��"O�9t씙w~V������R٩P"O�ty�!G�C�4�(�k�>l.\a@C"Oh@�v-֙h9�Ѩ�.&<�J�"O��Ç�(�\!�Րi-~�(�"O:�a��wO�(ʡ+^�0�Q"OD\��YR�eHD$[�6N�P"O"p� IE>J@T=iS#�+{�]a"Ol �4*�3=���*s��L�"Of�0�A��.��%C�4��p�"O�X�IӖA�¹��c��9�ZE��"O�@��A¾v�18��!?b�$�v"O�%G |���b�"����r"O�`� �faz}A���!"���I"OD����!d`6�{�.7�(��"O���,��7ǈ�VZ�V�jQ�"OBt��ˉ�U���`�f�8<B���"O�'�	�J͑��?;R0�%"O�	c�� �$�e��eV��k�"O�i�	a�b�C�11D�A�'���hҢ6uˤ�(ׄ &����'�!:r��=^g~��ʛ����s�'����c��Pt� �@4����'Ky�c"3'U�p̂*꒽��'��ue�F�i(T:�[	�'N0P����1W�$�����<��'1�i+#�D�r��`��GBћ�'p��SM��O��U��%�sT9b�'Cu��ßEr�Q������'F�ģ�M�e`@t�z	�'�B� "G��w7Xd�����1�l|��'�RHҮP����HC.{����	�'�&�ض�ӷ%�y ��r)�ѫ	�'�.��b��2Gg"�SP,�$kC����'(�P�>�U�v
�2m̔��'��Pq��*8GfuR7k0�\5��'�>��t�[�o�fyyv��m�q��'�V9[r�� !���NW������ �mxq�_Zz������,2��g"O
����.��"4$�>By>�33"OR�FF�3*0�u?m,��"O���� �:����9�f�A�"O,�w�D� �&�� E
0��<�!"O��q�nB�&�`�0�#4?� �ڔ"OF��a�N�`ބ��1�W�l�.�U"O&y��%9j�@pS��!j�z)x$"O�I��,q˒0p�d>R��4Xv"O�ܺ!a�4����Й x�Iq"O,�E]�s��yT*�Z�xx�"OT�:p��A�n�YR�7Xx�rw"O3^|�Q83�΂5�T`٣cV�"8!�dK��=��M�/2h��[3>�!��><S�=ACOy&P
1h�,0�!�$50ή����܅0���S�8<!���'<���B�/��9V�7�!�dݻN�
�U����[%�XqP!�dG< �N�"��[�[�f �͘0#!��O%r�i{I� �r�	��ǃ!�$�Gݨ<`��@I�ZT��iu�!�.�d�Yҭߌ5����aH��D!�$='�@����C�$�Ѕ�q��O!�$T�P�DM����s�p9!��j��tY�k��2�(mH�b&";!���]�PK��-aã�6!��;RN�,��U
I����c�#v�!�D	�
������\��9�$�γ
!��X�K�n�
�kP>�B$� �X�g�!򤗪[�V��UI�R�pd��f�!�$̊{	���4�ъw��s#E�lC!��,h��b�Х���3�$�g1!�\�l�򕪀���]�@�c	�W�!�dN|�>���V+���2B��m!�D���AN~�6���V!�䁷�\A�3AV�|������ְ�!�ޅ��P�,ϧU�1�#�؄]�!�d���Z�X4��;8QY�%�2o�!�d�/qu�	�t�H��܍�d�Ex�!��	�$6x�2�'�|ɱ���n!�d�4;�֐Q�H�$� �!��)1`!��'O����� ���e�[C]!�6@d嫁��m�ε�%��#N8!�$��PH
��� �&j�� x&�� �!���+`�"�˔Å�.|�  �-��i�!�s�*É�Tq�-��Rp&���'f��"C,��H,C���WH���'�>���i��Mr��U�O4Z��d��'3 <��X}"%X�@C=Ry\���'�8���iȔ!�:����#L��	��'�(<��+J8|���E�
5l�T��'w�B��&zNu�Oطj����	�'���j�#�~��ś�Ȅ�L"	�'bc�H�Tt����<�f]Q�'rT���A0~6������oh��'*������6?��
Q	E^}��'��y�"A�e�6<*7`H�R	�HK�'�ĽI�흦q�����>I�0���'J� s��K5 �zu86�V�r�,�'&�)�gb��0�4�������'&L��­�/�r�;4��}� �r�'�� ®�4d����6z0V��'P0̻$g�<\-��ACGY�l��	��'�4�+T�?/����U"x��T��� 5�6a����Em�_�."O�@���9
F��a��>*1�R5"O�2�c�q��}Pe��D����"ObD��&��I��*U���,G>��"O����X�A%���lW�Dkp"O��R�F��怚B	��&D�吓"Op	a�M�9V���t�N�r/�p��"O�x��΃TV���֣"��Cu"O �XSgT�il��"��8!X̃P"O �a�
.�@�4��5P{F���"O�u��KjH��aӲKn��{�"O���Ά*`jx`U��K\h��t"O�Y�J�3j�hQ���R�HW"Ot��6+H�F�:�Z�#�XM�lP3"OL����&W}��aћ>-n�Aq"O�1���G�s�8�;�M�o����"O�=��F�'Q���(�/Rl�e�q"OV<�7M[�IJ�Ǆ0sZ���"O�8y��Q�^�� �IPz��3"Ot�1[9"Z��Gf!xE����"O���K�$|唪�Z�Y%"O�����V���"VD��8�W"OXLI��c��
��Z�h&�9��"O�4��Wm��R�D�����"O�8+��@�L� ��6D�&Y�"O@`B�(ٴ@C�-(�n���p"OvY��FU)3;�¡,�` ���W"O��q3��&���!�t�x� �"O,Ty'�׊M0(���.�|m��"O(�YFK��)�M�R@C7u����"O�=T��>m��ѱ΅(W�X�X�"O�{箇�>rL�D.U�Q��8�P"O��9��?g ��1���o�P��"O�,�rEP��h2P�ǥt�& �"ONygMk�����eCR-j�"Op�)�ϟ������pҲ�(F"O����^>���)؈'�|�e�*D��`t�A*W������r���P�#D��@P/E�`F�	b�jVA_��Q�i!D�,IRX�n�6�1���BL�U�;D���Ti�=Sƨej�	�Wd����:D�������±8��3V�s��8D��[�㜔s֐1Q��$mǔLZL1D��� ��&N����	��{�(h�a�.D�t`mD�d��sp�؃z!xEJ.D����B�PQT��,Y����A4�*D��i��V̦9�K�9��(�>D��`F�7ka�3�U��l��F'/D�$I��V�6����i�#nf����L,D�DK! �)G��!��	�a$D��Ee\="=����4��q�5D�
���3д�0�i8�t�kS5D�d�*�/F|���-ܱ}�V�B��.D�`����%^^�A��,M�:I��+1D���s�+S���@`2y�:�D�:D��12�]
2�$-�1券_L�G-D��Ug�r��x'���_f�4� 8D���g˗��!B�^;)V\��wL5D�H��b�0 Rt��.4�9 2D�q(J����A�bd:�+'/D�,���Ŋ|;�Ȧ�H;  ���*D��D��Y��@M�w!D����5D���Dǅ�b�[W�ǋ� �sA.D�`��c��mS�ݣG �9������7D�� ��87�ӫ9�h��-H��{�"O:�H���*P�wa��q{~�"OV��$͚���2ơڒ1@�L��"O��A�'�lc���>��Q"O$Qafș�|i��3dޡn$h� "O��ţ�?6�0���=(��"Ob��\���tZS�ާj0X��"O慠�N*aQ�A��&�2��"O&���'Y��ƄJ#<`d"O�ɪ�O�bL�H $F�nLX�"O���@��B��Ҋ �ꨪE"O�=Ѵ&�7avq�v+֫BƐ��f"O��Z��R( ��A��U&��0�s"O�� #*F�����I��a�@"Oj���Q;�T�B���Z�"O��� �ÇI�؈�FB�?���5"O�@Y�,<K� ���E����b�"O(|��;	�!�Mk`���"O�<�NQ ff��� �EVH�T"OBE1��B�4���is���n
��#e"O�ă��&kRp�����)�N��F"O�Qñ�ʋr�\J�����%@#�y��T f���sT.ϕ�6�� B9�y��.h����V�r/���`瘡�yBΖ.'��@�R@A���ْ����y"C��;X�]���Jk|Q�QLW��y�F�k�����R(�k�yR.G�M-�(��mL�c)��y�a6�
���&�	e���ڞ�yB�A�E����F��b��`R.���y���E�xe�C�L�N����h��y��I�8�g���Kf�%�yb��� �@#��/A.����.�y�	�'bΈ����A�"y������&�y�sX*4�����9� ���y��̭J/��y��\~H[C'
��y��Y�JdN��4�ˤe�:Uk� �
�yL��{ �[b��P@������y�HȍR!��@�i�2CY�t��B�y"
�8;�ƕ�#�?�	���и�y�΄�Bd"��!�	�rm�u+�+�y��>������F5\ ���j���y�B(dqi��_�
 ܓ�CB��y��sԥ��D�'�@���
��yba9cB5`Vʌ����T*5�yrʚs^\:A�_�3��9�.��y2�۹]��3�H.v��ч�W��y�%�?=4�Xu���$Nj�����9�y�[$tZ�؁���H�E�#�y2K�"0� �`�\�b�j�6����yR͏��ũЗ]��9r����y҅��FH�w#��d�C3�¶�yR����T�"iO;	�Q8�i���y"_�.��j"D������F�y�b��\�����5.TA@�l٤�y�NF=a��)ȡ	��gh2��oD��y��}vQ��I"a�̐����yB�^ �R�F#���"�y�,�=�"��r#
��5B�FF��yb��>S/���
.5ȉ��E��y�=O8~���
ê��c��Т�y�[�OR�����
�081i��yb�",/`�Kd���%�p�#��y�g�\|��+�ϯT�^	��C�2�y
� �$�f��	Tu��4l���"O�U�F�9t*(��뇏R�0�@3"OPD(4�
� �H�!K�>�.�!"OP�B���7L,f��QOƓuC�rc"O^0�o\/ Q��)��C[!p$@"O%���		5��Q�\�pS"ON��i:~g.�b�e] t����"O:Xऋ\Y'��p#%S?�r�Zq"O4���=2Q oK�Q�r`{�"O��Z!���ړ������s�"O��V�1>ފ�B��n�" z�"O25i�,��̜�	ļm5"ON���`���0�FI��Lt�b�"O�Uk҄�_���C^�0F0�"O����kО������cϲ��"Oh����	�v6�=�Â8�$�#�"O" �ևW�2(�����{�*���"O���'Dgp�6ƌ>s�n�z"OF�;�����`A$�Y�1���	�"O�hCQ<�i���q`<1
�"O(I��NA��ݺg��V�{""O�=�r(��J(J���(z;@%�"O0P��j��B��2R+q4<���"O(`�!�
oN��9��o!���"O�"��0{~� ���b
0�br"O�Az�Kۏvt��mX�xz<�"OT|QQ�Է5��ܨA	2c����"O^�[�L�(C��3�@˸?�X��w"O�R��E�[��a�MI��Y��"O�yk���	k����Ì��d�"ONpb�F�"�n��̟x�`T`�"O�0(�iݬrĴ��*�>},\�"O���&i �:���hGJ�4f�\��"Oy� )�!���gm���@(�y��WZ\�ѠҮ8��ѻ�.%�y¥�R��t+EJ)D�2e����y�!�t��HaAڇ!�FQ�h�y�g�2n �p�A��k&�`��i_��yr�ڢuԹ���v�`;vn^��y«�'Ԟ�sу[�h�,�` ���y��h����W��c�%Y �J*�y�G6�eH�͘Y�ذ��d�%�y��Ԩe7,e��I>"������y�c�"��+�%`$T��	�y�K�]�V��CNƚZ�`��z�<�!.KD�u�+����S�bAG�<��b�>̆=���^�)�q��C�x�<A&�N�$˂� ���Y�><�m�v�<Y�BI���"E吻"�X�:+�u�<���)U�.t���9Vl>����s�<�WX�i��|�T�9@vHq(Yl�<Q$��
%�X�Q6�+&��ƏEc�<�%��L��ƈ�V��h�@�Zy�<I��H
���ɕ5LF��F.@��ybi��i�h9R'F�>��)��ˇ��y"��7߀���	�/?�h&bǌ�y�C�OE|��Rcܐ%� pV#N�y�耧Q��|0���;�X5�N��y"B±k����aJ�~j�3�=�y�"�gp�'��.R�1S	���y�����l�Bo̚�4�{AǄ�yr+�18�Zb�Łi�@xR��4�y2��)�bA�'m��WF�txܧ�yF�$S�X|f���$�( u���y
� ��Y�&�=��&��$r���"O!)S(�v�ल�fJTkļ�F"O��෭�	��H���*	?✲B"OL��%�����S"��58X{�"O����H�@��&!T'��h�"O�<��c�<���ώ�7C6�B�"O����\��I@w�E[!�(S6"O���Z�a+���*�`�RtA�^�!��S�m�-r����L�Pa�1t�!��כ5�����X*��Y���F�!�D��
�4�#J�n�Pٳ��Nn�!�L&!�.z�E�;7��dc`�� @X!�d� ��U����L�l� N�>O!���	�r�30@ӑ  ���C�TF!�$_�c�D"u�. �hچ��T!�d�$���2S�؂L%:y�� ��+<!�D'l@ 䡄Kϡ\�!n�<u�!�DF/s���f`�Dd%�`MMW�!�$�'qUB�Sd醵*\�ɘ�� �!��'�V�stmG�Rsk�S�!�X�6S���P�ɞV2�u{���`5!�K�%��S&M��Aa��J!�$�VMdX�Q�4t�,x;6E��J!�N�	���`�(u�H�rB��A!�D�4^`��PV�<�^��E���!�]� �n��*
���D�1�T�:�!�DQ�7Xh��'G�+JD�c��?�!�(T�P��"�="�0�� &�l�!��%h�4)(0�E�8��x��J��!�0"�j���+�2��U��Z�kf!�$�Q|��8V�ؾ%Ӳy�.�7!�e���'�$��e�V�W�!�D��-�tܸ�n��װe�B�'o�!򤆪!���0@m70T\[$�!�d�QE9��-L�Ӄ]�"�!� S=�Q�d����1l�4�!���7��G�8WuX��@*/!�d�AL�LA$��H>�����
�3!��ڒk���t
��>Ny:�IƮi!�D�2��,J'4AC��R i]�0%!�$5�h�EB�r)jرg�_�0!�dԿg5�4	�G�6B��6珸K�!�Ԝ_W��� T�`\�B��=!!��V�J0c�ŀ-hμ9���!�D�����
�O�tl����N�!�d2L:3#Ԋ'�����?~!��&2���#x�F4�Ci"*�!��Z*%���J J/8Pf��G�?�!��Du'��9#GS2|G���#H��!�IP��pY�IC�lQ� #��bz!�DB0t�ꅡ�Q��1)��U�5j!���\Ȋ*�l�,l���`�.O!�D'LjN0��f�13��ݪ��@) E!��\��<�P	\FƠ�IV/&?�!�D��i@��'KD�t�V�C��z�!�8U������0��kc�E�@�!�D�	-P|ɷ�Վc�
��tf!�d;26�O�"��!��E��!��C�}��m�����N�ru�ǏZ�U�!��RR����b�f������a�!�䋋x��2�U:sZ�4�!��(L�!��̏yT�U��	�C��X{ҧ�}�!��!O޾�BM@�O�������<�!�D�
� 13���I�a3aC��MC!�� ���P���Eݤm�壀E*Z� �"Op��(X�E@�	���)���"O>aaq�	�����O	(`S"OlmA�A��6���A�1�l���"O&�#p.M�B<I���a��Z�"OmH��*�Ac's�r��"ODT�NI7+��%�C&�4��"Op;�H�P�4p���	Kܨ��"O$���̍	y �B���	f��<C3"O\M{���s"�8¹2p�ᒇIV�<�w/ ._="�;妚�Y��u�6��R�<�Q%U1����eǿu��kj�<�����w jUҀ���p]QW*�O�<q�8Q*�x"Sʃ69xI��cDf�<��&5(,�P���2)'D�SnKY�<A����Q��r�	���DT�<AV� r�qRs$B�X�(	�P�G�<IǇ��xTn�`��(���(�H�[�<I�ʏ!��!"diӸ:�\�h�$U�<���	Ur4���W�8Z��BP�<�SAVc�4A����%-��JNL�<)U@��H(���%�I12�ְ{`g�N�<I �E�=�`l�֌�4t8����S�<�f���k���!�aHA��)M�<F�ףjHd��N�$c6�__�<1bE�:�"=@��18��H�Ef�[�<y�+�7�V�s(,Y��d��MU�<QC݂ �|����B~� Mz�<��㘼P��R�)��*^�����w�<�toӈ5�\e)w�
�X9@Q��Y�<ɐ�D >�ؒm�"����~�<��	��p[��S�8Z$[�I�E�<Q���=7P����D[٪EK�L�<��[6+�������{aX ���K�<	�IN�x�R�����}�хJJ�<��2ih���c�u����I�I�<����9AH����N�P0p�m�m�<��!B�$����>?}�U����a�<ɑ��v�εb�$@�>՞�gMc�<b�ܞ\:@��oІJEB�d\�<I$�
�;d��ٗ((C�*r#�H`�<�bB�4@�m� K�%+¢��!��X�<1��Ŕj!Ƥ�T!�M@��fO�j�<����0��mf�Gb�$AW�Sf�<��߳Aǜ�ac�&n�ِ��[�<	�B�8��8��R��M�0���y��L�����,7�`:!�
+�y�EF�0��Ar�\��j��@�@��yB��F#��Xa�O��u�p�R��yr�[�I�D�>W~����L��yb �n�>y2���Q�I�B�ɟ+2\d�s�ĳ`XՉ��q΄B䉒�>MB0ό!a�Qg���C�	/G�>����@3ahq���&L�B�I:c��q�����X2�қ$@�C�	7j�~�����l�� 杆_OLC�I�<L�D��߳]��$K^�W�
B��WJ���L�/ꐬ��ߌ��C�I�r�����o��`|��1*R�%_�B�I��Z����J���
7��D,�B�	�Ka6	5� �O*څ��Hš�6C�ɕ���i�>T�w*}�B䉥H��(��f�e��`D�C�[4�B�I�J{�P�G�L#�TJ�@�EB�)� �A�F�+_��Y�%��5�|d"Oı�q���0�xac�Fb{F5�"O��C�"m��J�Cl?����"Oܠ!�ꀄeĺ�"���+|&�u��"O�T���U�k2P�jt݄&�"R"O��6��C�������s���"O ���ډ�8ۇиC�>l�c"O@i��;|��ˤ L)B����"O�q��,�p1&��,Xئ��"OJ��	��"�]K�N�;Ġ���"O:e�x���P3�̷<�,!�"O�Uj`�5(�8��&�5���K�"O��J�G/@a&Ɏ7����"OضІĵ,Y&`�G΀@��$G"OX�1k�:�]Z��*9m�i��"OP�(抅�v���;qgԜwg�q�"O������#|��ط@X8�y#�"OB�D��/�)�q�T�)=~��"O�A�'�.o��D��]'���"O��0��j�F�"��Y�[9� 1�"OL�'��,���*q��3�P"O@d�A�#�f�HS�]�\��3�"O�2PȖ��jX3�� .<v�Z@"OVĚ��z�]��O)���6"O�!�&Y�"�uR�IE�f�ڰ"OB$����H/H I�h��a�4x0�"O��qN�an,]��(��$�"O���d�˜�Ƞ��/as��"O΁��&���6���Vc�${6"O�)�r�	$BH�Xp��-#<|A�"O��ye"�t{2���̈́R�v����.��g^#k�*�(�����~U�#��8,�J�Q��̴}x���:,j�&D���Q�U�A� 	��l�|⧪Q#@���"IfFHA�ȓG�ȳ"+C�D*h����"JjY��71ʽ�G�G�\�d��&�7{��$��/�����!Ǥ|�����GE4C%���ȓG�x@kD(Ն$���Yw�Ѷ8����X�89 ���4��G�1Ú��ȓtO���d�"4��(�T�͒����<��['�&3P�%p�"�+�q�ȓb�x0�PT�ģ�3u��цȓv7T:�L4)��K�e�5Sf���_�q��m�� ���ڗn�/,�9�ȓ z�O9dNp��b�+:�pY���<P�$��p)�#��#7NL�ȓ1����I^\�s�N��5��2I��r׋A���b��x�܆�+kΘ��

(29�4^j��x��cAV��)u�b����]3؊=�ȓQ]X$�E�BQ���rd@�ug"���r�||��%Jm���� �D�>8d؅ʓzĂ��Ë��}c.3f9C�ɯ3d�ݫ�Pے���H�=z��B�iX���C��-%Utm��#V�w��B�	$ES4�f��0%d@�B԰WC�I��\i����VN
,��f��D-�B䉺oW8�A֩�</�-r4b��B�	
K^��y��Hc�� !U�B�I�'Lr�W� � P7e��:X�B�	�*�Z�D�H�P���MPB�{����pioP9q�P�jZC�	����Zj�ȱ�hʁv�0R"O� V9 6f���!��g_;I�j�h�"O2��.�����}����"OE9�Q znHB���2(���HV"O��dDS�J(S�)L)&
�Xg"O��a6	��)�X��#��4�Z@�"O�(�6NҒV��t�nR-���B"OH,s!�q@�]{ Q'D�H	HP"OX�C�A]"q�0��i[.K�j5xb"O��u�S+t�q?s���"OJ�3��Ȑq�|pp�a��z�]��"O�a�X�`��`�JQ�pv�X0�"O`�5.��5��i� ����r"O �L��~��[�_�z݉�"O,��Т½����"gW7'�a�"O��"�
�b\�q��S�Ydd�[V"O4a�u��n���g"J6+�壓*O�`
�h�9��T1ш��
� �7D�X"sBN�W2HQ��O��ɨ 
)D�)3�V�f"�HE��u�B���(D��"���	&1�D�Ve˕0]AU)9D� C���@��*1)H�M>��6�,D��H�i�;>.�I��!ƒ~<�u��*D��q+Y�}����$�1�����-D��p���>a u��!.�y�D,D�(Z�.˅;X�R���A�t�@�)D��"��gIB��������.'D��q�b�5x�1�feQ�y2Ef�&D��Y$AEF6���P�J�.19P�0D�<���5����"����NAB�E-D� ����@Qp��0)v��dY�B�� DAK�.�\�g��M�vB�ɯN�޹�v(��dB���BBȖZ<hB�I:T��x�#̻"���� fS�C6B䉔}C ����G6�x��E?�B�Ib�!BT�Ti:�2���B��B�I>{�Y0���h��5T����>C��"L�U��ͩ-x�}Ѕۘ(�.C�I67sqh2��قҥY�P:C�I�Q��8i��N֨q�fO��W%4C�	�H�Z̡g�� c�1@�G��U��B�I5�2�$_B8D��7f9$C䉜T	�C Ë�'�A�����B�	� >�4�f�˦o���L
Ek$C�m���ȵ�.�f9�ҭT<�C�ɚ��@2�E��7�L�#&](k�:B�ɗH�T��reD'qhF��Va՝�,B�	'���c"ы6D��fǃ��C䉃E�B��R� #DЌ8RI3�C�ɣak�D���_���q�,D"��C�	�b<�4K�TD]��a�J@$y@�C�I�m9j��Ō�<���Bp��;T6^C�+hҸ-
�ջr�Z��Z��B�	/��)``A�9W(�z�eȅA�C�I�WT�`���,,8��Z�.d7�B�	KZ`E!�&Y�0�����C<
�B�	�{4$	���MJ�y�j@�u�`B�	�^腲2�A�j�\��Sf
�4� C�ɬ@\���#�O���Հ�K�C!C�Is� Hウ�6�y�T-�'0�B��*t^����Րl�!A$)�e��B�>o�=밊�k�tM('G�&��B�I,N���c4S�z��С��ESHB�I!
����Í���hm���F�b�B�Ɂ*3��34&�.&�0	�q@� zTB�)� (ReP*@�XHs��Z�Dp "O�4a��N=c�T�`�'�R��yB�"ODX�v��6�M����6Ur�hpD"O����]�JcͰ$F2l6�A"O�<#vlϏW�t)ѡ�V�
�64�p"O,� �Zhԋ`j�֦N��y"�Q�;=2E륥I��L���8�y3��i����d8����y��L<$Z`��Ռɾy��&�͝�yR�ʽjr���CAA'�M��MO��y��ʱcM佱g�	3�p+2�@��y��R�w�]��� ��M=d;�C�
��Fi�vc
��DڼX4�C�	9 M��*���5&����n�	D�C䉬�"�ʗ�L B��\:W<T�HC�	? �@�B��F���yR��E��B�	�'Fxi�b�j'L�8"�<�C�I�E���)�g�V�L@1��l��b�`$���:{�Ű�h�[<�PR�L?��O���s�5'e���ү��|9>�c"O*x�F`׍[����"O�)��;�"Ol9�6��7i>1�񮈣Y�0��A7O"�=��-7�WD�3@h�Z,	�"`�,f�̅�X��#�f��`b�x�
�%��Q��?[n� %	C�vQX�(r��¬Ex"�)��F�,9�ʩ�E/��e���W�<q�'�)��HZ���<>��X�XUx�|Gx��@�}nR-S���\8�PH�8�y2���-iq{ʶk����B@��(Oh��_�( m�B-0Ѵ�ʴ���!������RቬK�\�a@��!�ė�tJ�������8�g��	�!�ԕ_ưQQ���i�ƍ�ס���C㉦��`)	�ы@��;;>C�I�� �AY1t��U٦�H�0C�Ɋ=���9SNS#v��S�JG�FC�Y�`�R���#���A#�&>�0C�	�?��1��}lr�/�[G{��9Ox���T)��K�O��NJ�L�AO��d��b�cAbϟ,��ICA$zŰ��hO���(!C�la��N>W���"O��H��F,8)��k����5�!�"O
�c�נD�>�r�L�<`E6��1"O�h��ϗ��"L�l�\���l���!�Ď$#z�i%��;z@�u-�$Zi!�	�#YUIW���z�ۢ�uk!�q$�л����s|�C�HU^qOd����1|1	DJ:u��E��f��E�!��в\[���V��~��h�CfǇO�!�Ā�#?nX�B�<r��!��|���bx�̫1j��ry��
'�U��hD/�>���^6Ё��hP��8@�Md��1�ȓ;�*RU��y��Uh�e�m�����IĦ��?����N�h+�A����1��F~½i�0�I�N�bv%�8-���q�ʖkT#=���T?Ј�?>��)z�	�a�^ �DE/D�Ph���-
#j����A�(`�a%/��$<�d�<�E�X9ꮕHe���~xYg�>�y�L� ��	��D�H�!X0�y��%�D%)v,]��.Ԩ��ܚ�y��@��&���$��r��G��9�M�'� ��Y�O�Vā"�; �Z��d/��?���s>�����,<d���dnR#ѴC�	�T"�r�e:��2E-���'Hay�_�� Xp�AɜL�,��ƈ�5 �"O�I{�����}�ӄ�1%� b"O���F1b'��J�0�Bi���	�Y~?�+Y�2]2mCOꅠE���_�����M��I{����:�i�,BO�	��HO�>	�$�F��Ӓ�\	\�$	{�@#D��@ �E�64��/�s	V��r"6�O���O�D@���*�L%��N�'yC��S�'F`��ĹJ�H!��ď�r�
�'h�Dc���51 ��H�5
����'�>P � O�+N�=�1
ٿ1���'�����P�Y������kdРϓ�OB�A.���&�Sd0�yy6"O�(�HL� _�ЪB�	�s�2d��"O`}����bC&-�)�!�H`!e"O�0�'�nк�k��:&��F"O����[�e�`��g޽&qN�R�"O %ÂF��]a�����B����D?LO,I�&��s�i9T���(ڬ���"O��t�\�#B��-�X�35��1�y��L�n*1�����*����d���y�r���'% 7M0:ܒ'��y�C�9j�cæ�H�����D���yR�H)Uۧ��Vp:���Μ��xR&@Da�,˂h'S�<�(�ao��֜�|��I� ���JWO^6Br�أ`�;[���hO�>���a����|�!Jp^���1�4D��!��A�P�p0�I
V������,�O��Ot"GT�_Y(�xtC�<��	c"O��a0��hiV�!RL���c"O�9���Y��\px�˟�k���K�"O�rǈ�i���q�B|� �02"O2i3@U�����(A�@?X�[�'���<=�̉�@l��l+"�1��d'ORkWE�4!���3Q悯x�fe��"O��A���]�p�+q�L4KɰdR�"OB��3cܔ<r��F΃+4���ҳ"O���� a�sD�پ��L��'�1O@ȉp&j�L�2���*\�>�س�d'�S�'������ެE@m 0 &z�BmFz��~�Վ�P�����F�tl��i�E�`�<�e��5Y�9[�+&1��[�V�<1PEUR@`J�/.T�t�c`g(�!�$��YPZ��Q��Ҧ���nP��!��,�H���:��r�B\�.z!�D�'e�$TK�hߚ|(����n�Q�Ą�w5��d�H2~I�9���C�hGxC�'9<֩s�8z��sT-�-[�P7�(���R���D^|	��R�7z�ʵ�0\O��A�'���ɝ `��W��F��C`Ni��3�'�V�j���!/�0��g�a�nMx��d�^�P`E!K��z��JZ�� �KzR!�ߓu�%�D	�.4K�H�i��cכG�d������R��[/�!Ӂ�݄~�t �RO2T�p��_jZ<Y4�K�Ww��Q扔r�<�dC�l��i!�A�X���9�̃2Inў"~�I��CH�%��J���fC�ɒ,I^�j�� :9)��`P��/~cJC��
[�2��J�:$6�!���d��B�I3s�^QR#MI	��C�Dݘz����hO>�1Э_$4����g�[� Hn�*�I1D���SC��S0D1S�A���`t��a4D�$��+ Р���,X��,ڲ�2�I���Z������O�� '�S5���*�Ԑ[6"O� >���N=n4��r�HI�Y4<��"O�D��`I=;Y�P�a	�@� ��G"O���P2�+`��&*4�&"O�bv*�0J�Np�`�<t�V�"O��k�ɁP�@�n�"FQn��"O��aGÄb>���lJ�\�HR�$+���!x��脯���hRQ�M�����%�tPGB���� �鋾2}Dy�$#b�YY6	�6/أtT��SLC����?�5Ý�K�a�'U/�5���]F�<9sy��5h��Z�Z�SW�k}�)ҧ)���B
,>V�Cră�"�\��)% ܠ���f��PCO._���'���\��|�R �#r��e�c���Hg����k�Ԇ��oPf1geȳ�P-,!dn���"OnB�,�-�y2A��α0�"O�x�VNB�x�~Q��`,=���U"O��bCK���,��}y��Fn!�d#Kn��L�A�0�FF*;S!��-{1P�2R�P�I�&K4�&J!�$� h�PU�2f0H�J��Td!�DI���(��R�'���"O�Y��={���-���ѣ_��ybl�ILP�u�ƒf��7�4A�ȓpKPQjf^=R��$Iȟ�3�����dRr(U�ϰ.�}	%�([Z��~
�]�6�X:�j]Ձ��B(���R،�R�d�JR���ӎB�\�"���m��Y`��+#��1�$��X�p��b����
_xR��ȭj���ȓi�D؀b��6I�؝y$>p��D��{w i5IϕFd9Q����IXV(��Sv���e	 (����`�*F1L��Z�,Xǭ��w�`dP�NN����L�>-@�J�6G',��O�P�0��%R��2C	�
�X��H�0�M��AGJ��p��5������1V�	��t�lCDD�45Ra����p��e�ȓz �E��M��L�K3	�����<��1���]��՘�E�1 JЅ�P��q0�Aԃu��r�'��^V>��B9��2v��R Q�i�X[��ȓRy.��5-U�g�IU�]� fL݅�9��T��:�4@p3"��C��p�ȓ����
��J�Q�A
�|)�ņ�~f>��a˅:��՛0eŐ3�\C�I�I��i����<(���c�J�na�C�	�Q�u[EZ��`�s!���FC�I�K_,e�&�1'iv$�3%.8 C�I�y�V�X��Z�<AoK�%�B�Ɋ0;�@eN�^�1��ΜK�:�pC�̧V�J���������יS'<����+(l���2e
!�$�L��6lA�0���eF5#�!�dW�:P���բ�p���⃘X�!򤗣n¤��W����*��B�B2F�!����4�ŗ�m�
�(�"*Q�!���
��0����vTyj�c�!����.0�a�#,�pyc�+��(|!�L.P5�8Z Ɨ{Z�D u�I1d!��V��-�o4^q���@!��;��	�ǔ�$:Bӊ!-!�6p�\������i�� w�!�P0��LSD`�-6$Qt&�?N!�$U�A�l�����6��ma��f,!�� ܌;U��G��-��.ѩ@Q�,´"O�ͫ0'K.���4V9LZ�	k�"Od("����H<d�`��L&�dP�E"O��#��Yö�㣧�.�ΌI�"O�"o�r��H2 ��7���"O>��N�@ۚp����d'P�H�"O��ᖌ�# tĳ�m@�E��qB�"O���gT_�ZY��-��{��j#"O"x���;}�H	q��<7l�"Ol�1L˭=��X#�ΉJ.�A��"O��Rp��B��Ġ0L׆,���"O>�9���#]�V�1B
j:�J7"Ou��$зr��Z�C��i��"O�\����A��z�C�S� t�#"O�L�;8��b�#^�NU��"O^�TIB�Z'� %d`O��!%"O��3V��56���j��ʂQ-�ɓ1"OH��'���U�H�@�W^��q�"O&�07#��T%�FɝX�f�s!"O1�w� F��!y%d��`�1Q"O�XkqC��UE~��B�=p�Rx�&"O ��A,h)걈$�:Eʲ ��"On��5K� !��1���
�H�T9�d"O&K��e`�"�)�3N�
"O�� ��)�5��ʕ�G<�#q"O�bp�YB�X`��I�1
t	!�A���㞀��Y���gD[mBd��O�B4]#E�&D�H���?}Ш����F�	T�$!`�"?a�a������Q�N�2{�|pk'd�e���'�$ ��`yR�":P�@�$"K�K�u�����J�i���:,OJV�:GZ��ݠeoL����]�dlJ�	�@Q ��<J$읽?7�x+�f^6wN� ���2O����' ȹ�D��A]B��sH�b�"W �*L�L@,O��Sv*��2Ms�%��Ҹ'� �S��S����SfM��a��O�\�fH�G�� R��F� �DG�2n��$I�+L#dO�qY$��ѳ"��0&?�z�cE�k����eUA[�ie�=,O�"�˨0����PJ�;�?�> b-�SC� PH*)ڒ��r�	�RO$5��'�0xB@�A�Y.���fٛ6F0C(Od�h�fKfg�LHa, ��Xj���k���4fM�eu�!#2%S(=�\M*�O��J��m�����TE�HP���,!C" �m��I:�%Y��a��ϸ'^�IrOE3dKb�K�^(2���aZ�abc
�nѼy÷�2{�<�!p�ə1���mڴy�=�ǎ3lOP�3g	�4�l�{$@�^ؑqr��%4�V�����_s`0�&���뎘^��h�U׀g�ґ�&� �b�!�dǲ{D%������yS���#!��I�v�8`�g�m����1އPˑ>��ЃZ�s5�g�Bcա.D�����T�_3� `�oO/s�L�$���.�Z1�U�ʀv��D��IL�qOX�S���ws�50Be��l.H���'iX� b�����P���$#�E�4^,�� �M�	�x<�0�"0az2I4D},����iv=����ְ<�S�y��$:����?�"�Dʨ&�8��1*Ӭjؽ!ʏ��!�����*C2
oFU���J8�=�M<��E��l�~(C�k�u�P�}�Ҡǃu����յ�I���k�<1CA��@Y0u��L�)�h	��أ1~�*�EGy�e�a���y�$��0��.a{HĢ���:[L�ͅȓ ~���ܗD�:�c��0,�������^�qY��3�O���� ��H����a(�
���J��'=�K���Ry��X�:�c��W�J����Tc��yRn%P��!� ��L�ޕ��H�.��'�ڝ��(�-�UF��M�$XX�IƠ�MP�5����y�$����!�nF{���$OOJ��Р���g�����4txA���Z~Ș�^6^�!�D�< j�s $ɰ.;~��,}!�D7z�Lx
v �l��W8R�aR*Y�o�&� � �%��:pUY���!'D��H�Y7ԩ��a��p>y4
M`h�	w*ʩ��~�'mN<�Q Y;& ԥ0�L�Ċ�l�)R���s�(A�	���yB/3�B�q!�~�. ��gؚ��	$�>QX��O�4�a�d�i<"�Ksh�|E���y�3;?,M ��qhL�c�dM�d!r➴z��r�g�d��.(-���ZI�,$��w�!�d�	$���K©#��+�ʊ G^!��@!��L����PI�&!��B�K��_
_�0Tv�T!�$>fS$�Ȇ��Q�f��V�W!򤗕?^4����\-
�2��d�t!�$Sj�dH6�0)���z�P�xJ!��ŁT8~-2�\�9�X��v,�W�!��S"��P"��7B��	��^ ?!��g�,�Yj���
v*[�!��&׸�S�W�)����)�:9+!��W6Xy灕�\��]Y�0A+!�DK�s��D�vI����ɀ�D�&r�!�!{D���#���sM36�׎b�!�D����Q��K��+.B!���z�@��L�*��\�@̇�I#!�D��� ��f�!j�YD*�	&�!�dӋi�d�����ml&9a��W�A!��ȗ{�T]i���,4�zH�f=!�d\�-�`�v�E��L  5ܖu!�$M2$��X��h�8�,@{�J��`�!�T gx�\qR蝾b�|�5JV�0]!��ٽ2G��Ҕ�J:�z4!I�*)!��/6�0њ���&)q�h`�c"Oԁ�p�	�V;V8W���f*�)�y"�$>"`Q����:$���p�g���y�-�%r�$iQ�ؕ�TYb� �y�Z�s�
PFwo��6۹�y��ĳ.O��#����l�E� �y2��wM�e#ce
�;����䊙�y�΁�uޠ\�qJ�a��TsAg���yr��,9
�4���b̜Ȫ�[3�yB��}[��f+�8r��J��y�DPSQJ"NX�K��鐃Ŏ�yr�Z*?�䡦KͲ7�Lҡ�y򏃑.�l�`*65�H0�5�yb�,a��c�� �����y���l�^!k��6Iq���y��6$���b�Q���� (G:�yrbªB��[�L�V����C�?�y2j��ٸ��2qܺB�Ǎ8�y�cެ4�th�Fl�'~��1#���yҁ>x������i[�YQ1���y���x�¼K��7d��Z0���y�"]c��Ҩ3W����FޡNV�C�I��^T����xH���D��7m��C䉢YL|���țCڌ�0Ec�2,�C��D����Z��8R������qI�"O�E�A�H�x?<��T�$.�Bq0a"O^�b`OOcRđK���9b� �"O
��ABC�H �a���u2�E"O
9�`.�S�]��	ݿyRP��"O��"$IJ|�L��)L�#a�"Ohh"�`�;���PA�2�\��"O|(s�h�[ J�H�`�%�h��u"O`y�(P��x�rE��x��b"O�U�3�w��1ZSM�x��8AT"O0`�1� $Y����+6()j�"O� R �fO�!�}�%M<m-��!"O����\�O"����O~�p��"O��Ɠ�h���b��5zg�Y �"O�ESW��({�*)��Ǭ%y��G"O8�Q ��:����Sd��DR��jA"O$�PsE
J��%��>QO�����'���*��h��N$��R�KU�%���c�`ǣ8�!�d��\�D�E�� ~YyY@�,5qO� ��6�)�	X�eA|۶���x�{�J%!��X)I4����A�xQд��L�|�!�dخW.��bBb]����%�#�!�q�mJ�h�dGι�$M!���)�f���U�m!D��#�P?#)!����D|D��65\�ɐ�Q�N!�$��j�YFҍk�Mh')�" �!��6k��[d�Y�Xz"5"3h�-@8!�d���Ł��\�+�P�1�=?:!�O�q]�⇥��Q��'O!�$v7>e��%�%YQ�a�R.8;�!�d�F�����S�Ή�g�P�"O�����-&���Y�m�L��V"O��!bj��pp���C�84�� ��"O��B/�!C
�Z�nѺH�Zd�$"O�\Je��(nx6l�����| [P"O���6�D:}|8IR��n=��y�"O����T�"�_S��X�d[��y�+��2p|3�ŭU8(��^��y�B�t�
雔a�0C�±�e���y��$s�T8��%�mG�t�m��yI	=8�.#	��h�'苫�y�%�$28��ɵ'K&��a��ꋁ�y2�X�q�P%F	+pO`�!�C]�yB	��@�P�BT3A�pQ`�H�y���2h
���I	8̲) ����yҏV+y��Ĩ�?V�h ���y���{N��	���,BA��	�(I*�y�������t�Ut7�Q��>�y��ɎH�>�c���m�IJ�dǏ�y@Mh�6m��� �tAp�j�L�=�y/��AV�����`�=�v"���y��Q2�Y����a��;#�М�y���_]�pp&�ďr���0��T,�yBi�j0�@�e@� ��XB���yr��<z� ��Ǆ�=���r����y�c$YX\���I�5>Mr��ɀ��y"��e�m:fÞ5��ܻ�B@��y��ۇ%28r����"�
��E-�7�yꌢLܽ��\w�J�ʟ��yLҦ+�(�{����m�H��y�F�8,&�uI")Zr��D�&ۭ�y�O�;>���0�	�k�B$Ö���y򀔠C��Xq닱dC�	A1����yr��.2�ɨ��-\%x���İ�y�-��n,���,LȬt�f\2�y���O����
�^9\5���y�X�@�2Шd%�_`<0�[��y��D�;V�����Qg���'����y2�S%=�|�т��Mj��j7���y��ڒnW�=��
����IC��yb�so6颠JHQ�j�d�=�y��u��sb�8X��󳅞#�y���s(����[
Kr��0@GX��y�M�	�Ԁ�ǗI � y�e��y�MI�X�����\�rM���ҡ�y
� VM����0jRd�)t���"O��c�n1V� a�T9��Ӈ"O((i�g�*q9�s��W�T�z�R"O$U����)}3�蒴 �<��H��"O�L��W >���h!)[�u�Ir�"OB!�#���,,�xà�>�8�W"OX	*0$ԏ�ޙ�r�U��փH�<!�'��t9�`�ޚa�@-�4d�S�<)��U�jb�Q��n�� ��	��L�K�<���4O�j!��&ķX߼�!�EA�<�1��t'��a�b�@��.TJ�<�%���2��%��h �2a�ƣ�r�<�U��6��b���LR��t�<1�*��Z`��F� �3�qE�q�<9f�\�B��c�aE#H0��1�[J�<�a-�tx�OБ4Ȳ��aG�<�!�;��bC&&L����KA�<�F��Gi�1�P��&��shy�<�F��>d�<; d�&{�:��1��u�<�'ȵ5MT,Yĭ�7��8�LRU�<��fԣ8��Հ��FZ��P@FJ�<�g��qX���5n�P�e  D�<��������B�${;�Q��L@�<9�j��`�TQ������I���T�<9SG�?[G���A7%גݘEbx�<��e��#@��VEL��S��x�<��%�H����b�=�N��pl�v�<u>v�͑TI�#$��-Dw�<�޼2'��x��xr����H �yB툹I��I`�EH�F[���C�#�y��)l	ܐ[�f<̢����y���$�N�@6�<"��,B�X��y��>n�]�q��� q���y���})�kl����)�c(R��y���5
B!A��]'
3$��T�1�yr���<�
�bЕ�$��;�y�g�$#��Ǩ��ξT�t'��y2GV�����G
����d(�;�y¨�4(x)�`a���(2$���yRE̦8�$��1N�h�L�&k�$�y� �to|l9I�c�f�(�y�l�2��t�)W��*0!�ؼ3��m�C��](A:b�X�h�!�	 �AE��-l���C�Sc!���:��ԢCh͵D�V=�d#P"!�ޯMp"$�SaΪ9���s�ͽ"Z!�Dܣ*Q�=kf��V�|�#�+ 4!��@���\!"G�,(�ȫ ��i�!�g& p��&7~�B�΁�Jk!�J+{�\���˅h�`2�CC	G!���Z��97Bh�ba["��!��n�$|�3��<Ay<����	��!��I7��Lْ
׿1V��z���x=!�d]a�V% �I�>56��0횘3!�+Z��ƂMF0&!���+~�!�	��H�f�8{�5����?�!�Tb�j�����=Ԉ����o!�#�>	�%m�4��
��4_0!��>���v�;:$l1�iDV�!�$�t�����	U>h�ph�(!�$D
(�N5��F�B��M�ee�D!�dM<[�DK�c��6�(��� H!�DH:*�x�s�Z9j�9tA�|�!��� ��b`��?A��Q�b�!�� �ФT�3�Rбt��.	쀨W"OZ1R�b'Z�8����:X�yw"O<�:���-zU+5$��p^
4"O���oL7C<6��R	B�
0"O���D����B���v��@"O���6B��fD[�R��Q`"O��p��\�ౙ��N��4���"O2��^>z>\���@Gz�xa"O���Q+^+4���� �'L`�"O�a��x+X�� ��)Bv"O�����W���h�6�޵E�3P"O����ۏ]݀L�t�	�?~��A"OV����y8ܠQ�i�>`b��
'"Oz�(R��"e��h7'ξ_x"O~�$͔B��̓�$E:5cF�1"O0[wJ	4_~��C�u�MK�"OL���F��^T��g���u�9�G"O8ia�"E�|��|���V�6,e"O�h�}1H�E�^�/8!�״T��L���/�Ɣ���؋w���	�f��aAn��<��p�,��y2�N"Yb6���C��*��1�Ѫ�y2�J�+���ѡ蒛.ȶ�K3JH"�y�MJ�iR�ބJ[��l���y�M���=�5�]w2��$�#�y���:!rY��I\�n�>�2́�yS�w���C� p��Ejm�0�y��!�n�9Rn�:Q�1��凥�y��F�@�$E#��S=Fi�a���y�R:#0`� NR�=��pa�+�y��4x���*�(�y*|��v���yBm	=M�$ɨ`��h�M��! �y�%[<X̊�B��d�T��"��yR�A�cp�8C�_gj�"����y2
L/� �p�ߊQ�0	k�M6�y�-�4~���"E
M��d͆��y�MІ��B�88��8
�H��y�өd[N�u/�$?��*C���yR�v�lf/��4�j!�����y�au�T���	T�*2�BsϏ��y��N�:��l"�F�/H�
U3u(���y� �]��;@�ݕQ��eĈ�y�-�8fU~��d��:��"E+�y"ʙ"��dz0ha��G�F��yB�\�کS5��]�X���yr+�Af���m�R�p!�0( ��y���fLj�Q�I�F�D��3���y�H�ko�����=��ѓ����y2*��+���C�={_PYr�	���y�m�'�P�JO@���͚eI��y"��k����R'e����Z�y��5X�T1���z��p�b	��y���R����"� wۖ���J�ybbIo\�Y���(X�0��FnP�y��1��)��Y�Y9�B	��yh�9vI+7,ȝ �r) Њ �y"�]�r�u1BTU���pL��y�'�6B�!�c�-�2l	��yN�sOtYy0�	�W��i���y",��7ڄ�(�oQ�+	yB�d� �ybOW�hᰣ*�-�H���	�y�'Z&5
��ӵ��>.	,�� ��yr�@�B�H�Q�%bL!Q3
	�y��M6=��^ע�"(�y
� ^0`Oⰴ��#O�m��|�t"O&�Jd&�57"@�c��^����"Oƭz*�C� D��GFʢ=�4"O�� �kL-�v�0!J�&=2�"O$�k�J��4Z�)[�]����S"O��*Q��Q2�`�Ҕy�M��"O<e��j�wpv9xW�_%>h�5�"O�)
B�R$i$�0r��*\~���P"O���$Z#U�@Q)�)׵��Q��"O,eRA䅘
�4��c9N�~1�"O¬��]D��R�Fϝ~��C�"O�eA唀C>��槒�2�^�ز"O��0��"�v}ZB�����"O��!�̊�x=�Ɇ��:��G"ODYugߞOm�И�
W���-�T"Oؼ[S�VN�J��#Ǎ+���q�"O�����5<�x9b0'Pi��e��"O����! .#E�-ru���St:
�"OFUz��F.AFhЈ��_�8s"O��2'�^�W" ���˲f4t��"O~�#ǅ�=��MZ��6>)��I�"O�1-R�P>�D�Q��:\�}�c"OVPc5Z�U3p!��,~�R�S�"Oj��6cR�Ĺ�._,%� ��"O���q�N�L��Rg.�z�$q)5"O��!6�����`4��92�R�j�"O��س�_�e�a"2Ɠ C���"O��K# ٷb�\�B����"�fQ��"O�x�.C�r:�[��)=aD�ɴ"O�<��<������sP�M��"O�$
f�����cϫ[Wn�i2"O��S+�s�f�����an5�"Od��u��d䞠�@��
xҰ)�"OXA�g�'蒝�'&ˎj�*� �"Ot b��xH��.�����E"O�p�Ξv{Jm��L�T�XM`C"O�@#��s�b,��N�(bii�"OL�ڃ��Ĺ�CJ�!����f"Ov��қV��]�!K3r�&��$"O�� �ܘAƪ),D�]:�-�K\!�$��O��(��Lxt�i�n^	h!�d!D�T��!\!mXhQ�Rm΄@!򄍰#��pG��D�r�Ig�&)!�d�4�*l���մJ� )pl�[!���( X���
���b4J!�$�{�� ���]W4Y�w��V�<�Ra�-� �z1��� L��R�jL�<�cȘ}�N�I`恻=�d��l�w�<9b�2h�z��gF?*rPP�cN�J�<���+!����C��<�@ 7��F�<�����yآ���G��z1��C�<A%��{,AꗭU2S���Z�NS�<�v�S0{k�I�P�����:eVC�<ѵ�ߏ0ԦH��F��໐k|�<���> ��K�K��]дs�jPz�<��^(�8aƆ�ܩr2͈_�<�M�k���*�d�(sEƟq�<��K�:� �8�Z�&�*��B�r�<�C�-R�i��EQ�y8�:��*0��R���NW
��wc�즙Y�"�>�d��X}���xIׯ�6�����$��x�P�OĴ`�'��!�$�+��/�ɲR����ӴK3v䛐�Q�%y�듴p?Y��J�E��mB`�ȱ��<�b	Pa�'$?�;�.۟i�$T�c� t	꘣��~�'���D�ԏ�+ �&�A��Q��dt�H&��'3�2P3��~
���� ���0�#�<jB!'��:�\��p���
:c�"}j�!
 F�X=���Gs6%����<iĬ�38p�O�>]�P�\�b�6��TIU3il,q������1"�����!�,�Q׊�F�~�C�L�,��*�}BKg>{�E�0,e�"DSvV}K��%�	�vTyC���i�*M�XY�ՌGq
1�)!�I,7�j"�=�)��4`�fI3Ck�5c�yi���9TE��3�4\�!��?ޘ�	`�dM��yJ?9��$VY��ʊ�a�~��'˃=�r�I��+�'���֢}������#E�s�
��)�b)�=i��T>!tK�F����2(Ǝf�4P	>�f�0�}���/�bxp��a�͘LlA��.����	1$���?�"�O8@���;�_�RJ��@`?�eM���������O�#�Р�fg�6���ug�5E� 2�)M�jw�b��|RC��<}�
�0i0����Hţc88(���g��d����cN�1��VКlw@O'oL�㞌3��)�B"E1X�ɗȒ�vO�ؚ�ƍ�'Na|J5��Jǃ٣.�`JB�֩�0=���$^�>��=��u�t P&�L�\2��)������ 69����>R��SE��$v8�s�&F�?)1E�|}����ēUeDCr���%șd���-I�	]�"0'��y�(� RM�nT�T��i�+���y�E4
r(���#G���jAo���y�BF�A��R�.2���YB�
��yҧȲv5��œ�(���Fm���y2AJ(g�0� s�^�	�NS����y >`�I{wE�|"P�pE�6�yҌ��j�F퉳d�1zK��A%*���y"�Ω4&̋b*ʆsOƤ�D��y��1��ᒦߤuh��U�S'�y���8I�Oɻy>|�Ң� �y�
_
m���k���E��x�� �;�y҄PTX	�Ğ(���쎫�y���-�R��#� &r�-k�M���yB�V�%�H����& �b�bgd^��y�
Q�ʨŬ@eR���8�yR��8Y��� �W ��Q�/�8�y2`�>��0�¦wf�ui��M��y"��bn��hg�ܶo���@���y�(�$��x��d��B@E��y�Oِ0X�H���P�3����y��G-g|Iz�	b������ybK�6Nd��K*��X�Eꅎ�y�-�o�x�"����v4�+D�н�y�oP	XȔ��7��	q��y�D���y",��4��P�D�P"9M�E�A�� �y�"�5,�X�e&�,$"0����y�œ(gT������^��
��y� R	R��]��ǒ���t�cF��y���^��)SA�A ��ȷ(L��yb�śC��� %I:e��vN��y��I����q�(�%^$F�Ӡ�	�y2o�3��[�B�X�����'�yQ�M�"i�w�S~�	��y�b �-y�;�i��X�Q1Ԇ�y"o�*4pH�0��-�hT�C���y�� v69�E��Y�EsJ��y�K�|�	��kѹL~�[sϗ�ybʀ�f`�<#�".1�	�!E��yR�^	G�^d�$��%1J���q���y�/��T�3�LI�?�@���M*�y�K�#[������1��I0&K&�yA� wp\�
 ���.���AD�Z��y�m�(H����bӪU
����N�y�o %p�� �28L6��,�"�y
� ��"@����]�VM�����"O�( ���a&�h�)��.:�Q�"O��y�E�=���CIֳe���"O�d(F�*ve��Gʐ8v��@"O���e_�X�P�E�K��B"O$uˡG�?����N����"Oh�eL�9L���\%G�P�d"O��@%�/y���p��T
:ұp6"O��
���)I� �*��h.^x)"O�1�'	�07SNxR��:m"��R@"O�S�eM�bufT�to�"w�
��"O�@�ǁľ&��-jg�WF�8ܻ�"O ��P���%������ټ'��5��"O^�0�-�zj��f���0K�"Op��#�s&d�$eP0-���&"O���1JH� ��Rc�E�1"OF����޴Z6�u�D��q�X �"O�5�m�8ut��Ex�UJ�"O�U3��i*<8
�@Z�}K�"O�)��=H�(��"/Sv���"O���
IP�7�)֠pq�'D����K&|���z��3l��s�/&D��!PC��й���:ol�=ҥ� D�`��â'�t݀F�?k�-*��=D�X����V��������ey�M>D�L[r��<�iW-ҋAf����b/D����GW�� g��r�~��v.D���r��F�)@N*pA(D��`m��g���v�i���P�*D�H*��ִxM�ev�Ȍp"��9^�y���8X(z���'#x�RF�Z��yrA_����8�n��B����yB��XnD��DN�m',|K7���y"�ݘu�"	��*�4�:����yR@ۀ�T���ں�+@�]b�؅ȓNS�(�l�K`��r�I/F+t�ȓ9(��ğyD�����!�Ɲ�ȓ�L!��T�/�*����*fX��ȓZ��b��NA*�SMjBꅆȓF���bT
$Id�[Q�ܜ?
Pd�ȓw�ę�w�C8�ѱb��sv���{�4��C�/O���r�;}%���ȓ%�5���x�n1���< �+4D���^L<���	K� �p��d�"D��(�-�������5 mh��4D�苧�[��t�䁞L�})�2D����hC�����!(۪h�iTA0D�Hz���1�`B`�\� `bͩ��-D��Y�Z5=�P��"[�W�h���!D� �GƚsFM1Ci�1h�8B D�B ��lh�#��7� �Ah!D��ҁ^�h��m^"Mؤ+'�<D�˖O	�V��#`���FEp���9D�� �*K/z�Zv�PW�lz�k8D����_�gְ�@eΎ��5D��I�n÷ �h:�.MK��l)��>D�,��R+�8qGG�K�n�)6�>D�LRa"��U怑���W�Qg����:D�$�&�S�Z}�� 	���(Y1C9D�<� �;?Y�c�}���G�8D�0�4�G��pH3Y�*���ǫ"D�D�G�@%���TX/NپMa�?D�pb�Х;+�p�	�#G�Hb�N>D��0���#@sZm�q�¦@9"<kE�=D�� �T���)�`L( �G@�@��"O�#���c���7'����7"Oj]��)^#Nn��v�ͩ>�>�:3"O*m����8�@�ʗ�7�Q"O@"��ġb�TQ��ʶY
-c"O���2b%(�'�:�(Q�f"O�ACB��8UbQu�Y.�d$�"O�@�ˎ#N��캅�g�څ"O�"r'T�B�:��bQ	;�~��r"O�	Ab��Ҧ���A�D���"O&mr��
Vb9����1���r�"OL;6�ux�H�(�!�<q�B"O������iZ���fEP�\��Q"Oh "@�H�����O��&�H��"O"��%#ܜ]Z�	[��/����"OBqr'������
}��aB"O�u!�'��g��)V얈=�P�r"OĄ �G״�� ��ѨM���W"O����'A?Y�� %G��,��
�'�4�r+El^�;��ՍW����'�dx�"Ӟe�|���փ[nBy��'�H �P�Z>:��@0J�c<�Ȓ�'�P����/%XгD��Z��Hq�'�B9�TD&/�vY���Y�Ӝ��'m\xС�$����pH܉q�T�B	�'RV�c���<Nʜ���7;�A
�'$zq:�E>�Jp�ǃ.``��
�'��$Z�¸?l�����;�	r
�'�Z�B�/��R�ۦE<	_�Q0
�'�ZA8*ТY@iH
e<q��'^ި8׍I�)=�ዴ�C�}�$$"	�'R�%q��T�Da�� N�mr�As�'�Ɂ#9nJ�+�b��TQ�'�t�CC�T-A�4�����;R��p
�'h�i�N�BA$����	H��j
�'�&���6u���%��
W�4���'+�8Av�Φ
. ��T�?b��'I�i�1
$�d�C�d�j��
�'Yh��7kK!�r��C�'9�VKF7@|D ��?q|���'u�Ȑ'��"Rs�I1�^"y`��8�'�>ѫ��-!v����HwB:���'�8� �S�p�	�>���'�+5�ʷ"T&hs�k\�̄`3�' ՊhDi6!�ԊI�U
�!�ȓVn��V�G�|�H];Ad�	0:�C�	(oK����J�VaJ��r\C䉠,��t�fK�7 E,Ȼa� <n�dC��&�\�ڲOG86����C��fB�	j��V�e)����KEUnB�I��v��a� r�ȥ[�BB�I�;(��hE@�#~}�]���D�z�B䉈Sל<�Q�џqLvM٣�9FC�Iy|���̓X#vi�ă8}�0C�I1L���pb�B�.D�*�!�B�IPs�T�� 6��-JC�5�B�9W�NQ�g*�[͐U���C/��B�Ʌ\ӪU�T�6Q���kE�]��B�I�DY�۱�[�$*�!H�Ub�B�ɧ�@Px���X�m�B�U&H�jB�ɾa��	`U
�	�Q�Щs�8B�S @9�ƫ���Qz k�kZ
B䉤,�:�x�&�t�t�B)0j~�C�1Y\���1b�N�A�ʇj�B�)� ��ã��
�У��ڵZ7N��"O���ȟ5X�@��AHӮ*!R8��"O
`p�������wF�Xz�XR"O���7֖��0!'K�h,C�"O��FkߩKDX�gȔ.E|8���"OV�Qk& �zH;��m��[�"O��b@53��R2G_7�s�"Ob�su,��#�N4#LM:)� �""O��K�ˈBj�t�򨉚0R�#�"O�<��
��Cg��Q&F[�RF��"O:���_e�|4o�
׸%�4"O�="2�ذ.I mssS�)��i[5"Oܝ"4m#Eƙ���Iy��� "O�%�V��nZj�z�Мh�"O��H����[:��AB���f��|�"O�`�ׇ�[>�˒��R[�x�"OD��ҿ7�Tyc�ܾ�q��d�<��a� x�&���S�c�4�!�Tf�<��@(J�N�ze�;�
 ��*K�<����9RAt��d�Ҍ �Ĥ �GI}�<��C�wM�M���W�&H �U�<"I�<��� �Rg�e���|�<Q��
�r���OA�� �L�L�<��� �F��む�7�d����<�"��
   �O���|t��c��"�� ��'F��1E�Z�`[W(C�O��y�'��þ�Ei��Q�ްa�*�o�<1�o�qhl��ʝw�0���al�< ��,   ���[���$˪͙�y��	�;�Z*��7[&�;u,Ʀ!�tХ����q��x�kM���I2�'s�8%/>����Q�8zS>�9w@����D�q��x(çiTL!f�5n���`�.T�d"����OU���(j�F����
�����˂Č(ce�@0!(�4e���C�OF#%A@�-3�@���yr��O� V #�Ća��%��Q��e�BE�On���K�[s�D���4�t�0`+�Y?��2��&
,H!Pa��PE���'Ȃ��a���B.P��S7G�`�@fJ����)��u�>q{�*F�	e�� (���)�-Wz$H��bZ�f�@ʳ�^���4�����G_=< "~Bv땞W��2�n~��U+U�M6F�6<̓3�$u�l5R��`k$M�C��M�'[��M����E��=#�a�1]�T��阴�hS����S�O��TM��S`���j8�!Fǚ{���3��<��'�nܗO�>UBQ��F����2�3�v�ӄ�e̓�t�۔�=�N	�c#�^�b�÷ꑗ A��RS���_>U��  �>E���۽�09J�ω�T��¡�y/�#��I j!��%�ڀaCq����$@�/P
6m\�C2h@2.;��B�bD�S���Yl\��2I�����>T<P�4�b�Q6	C~]����O��2��%��ӵi=��M���ިs]|�Y��]�]��%mZ=)<a��Jv���(AF�+)��LZ�bJ��քi�/Ke�|>�>����^) �
���Υ
䐑�Ղ��?���Q�x%�a�g'N��1�$�G�<ɤ�ҐP(�)"m��.��pAK�<)�&@�,�r,�����ٗkCI�<Y`J'�F��de��jnI�-�C�<�7NE���(sA�Z�Xݘ�N�x�<w�յH�)�LJ��A��F^k�<q�	'l��!�Ҕ58��OA�<	g+c"xiI�n�IJ�Q�v���<᥇!�jxX��X�6�x���}�<��c�0d5y�ƌ�g0���4��v�<1c��F,>� �'Y�/b� !)Qt�<��,�O�0�k#U��0`�o�<�˜6�XPG=��x5mZi�<u#W�4n����=8�2�����h�<���"9a|0Z���K*�p�jO�<)�n�?cQZ��G�2����ІMH�<1����'��3#H�
�։�U��^�<A�	E�;����>#��b���n�<�Q.B��&��U�������g�<�#+�>%��rQ���[��H҄�X`�<�煈&3��S�B�,2�Q��]�<��Ĕ|�&���q�8P���\�<�G_�O���`���=������q�<�ì@R�`��P
�\srP�6�Cj�<i֤�I���g'D��@#��a�<�� Q���`@GV�>	��C,�`�<1�lW2A Pc���m"tacΉZ�<�%��8>��t���7E���E�T�<A��`��F�-F���L�<�Q@�5nX�$阨�̜Bצ�N�<1d�)<$̑҈��%$�O3=��'
4�ʢAY�?����N_]o���'�lM�ֱGpЊab�,*(����'@N�1E��35`���	�"MbDP�'ٌ��PR�M�D`��[�oZx��'�`�����{�p�.�=m,����'aN�ڤ�ɧt&J y�̖�]���9�'�0��p��?�����[�X(ЀJ�'�z�9&�8�t����r�a�'up<��,QejUS��	,5y����'����#jߪ|�b�
��~�(�'�d0["�΃\Z��qnۻSZtP�'0,1S�:KP�q&�ݔ+H$���'�̝�=�.���
�|-��',D;S�	�SP�qCkQ䀐�
�'��s���%/��BE%�d�
�'���R�%�(1��o�`pY�'X��6.Ŗ]"&��K�)d�H �	�'ˊ��WE�3XB����N�b��@	��� |��$K_ � W/�(JY���"O֍�tEǛpPx�)� $M���e"O$�c�!�+l���s�m� Y3�"O��g�#>�xD��"w����"O��p!�u+v��*Ur���"O����Os2�T+ �ߘu�ġ�"O񁶎�?{$r8�b��8'}$�(�"O�u*g�"X�.]���ʰ|B8�`"O�i���:M�U-Z�{l���"O$��C��J����\�#�t�P"OD壁N�(t@�����s�F��"O��`LE�nE&T�pL��y��A1"Oɶ�S6�p�)�`r�%�"O>�P@��5B>LzuE��Y�@J"ORQ���]2�|��͂P�x�"O�%X��Y��fA3���	�D���"O�Q#�5Y%�aa&���	��1��"Oθ�0D=��9R�]��P��"O�(��!<j�����W-�ܸ�"On1��-ߍr0&� ��8�0��`"OF�#�*.Z��]�T�� o�tx�"O��֏G�(M�5��QFE1�"O<(�tJZ�$l�q�'�i#�j$"O�e+K&"���Z3h�d�(��"O�=8��P�8���Ǌ�i�q�S"O$�Z��U;cSP��)ڰ*Nޜpa"O6��r� ����ℇE1Q��"O�Tt�Z�Ea�})�@��#��(�"O`�k�'�qp�N����0RS"O^�3�n#"ݦ�*E�!s�����"O�<Q���h��IƋ(�%�2"O��"'+ۗ������J*T�"O���u蓆��[��������"O>вҮ�<7p\x���;��9"ONŁA��84"�  �Bd"O����5n{�9��犾 ]l�iQ"OB�H ��.��|;`��%B��1#"O<�#�%ʾa��0�L.;�8��"O� �F�'��X���Y���"Oʤ듬�@D�Zf���-4T��"OT	H����z��{��->�Ѥ"O.��n
5�]�!��c3� ��"O���W�B63����@jǛ_D
`�"O.�v��i0ޱs�H۵0ha��"OD��&&�4!��Yh��@ ��"O8�*ʋ
h( ��e�1�Q�7"O41��I��-�P="ƃ�=3Ҽ̂�"O���
��w<�S�#�]^怡"O�Ls�e��}��⚚l[J�� "O� �Ue�0%\��u!�)�Zq��"O�\тe�2�B���ͲL:*�"O&�!S��6(ˢf�$M4~��"Of,�W�X*��4Ŕ��C�"O$�*��,	h-�Qኮq�X+�"O|Y��M�Nt�" @�O�z��c"O����֩�`eht��R�V��"ON)�W`
<��0�G��_��XR"O�H
E���hL���բ��5(�"O�Xb�[�^߈�Xs�]?1�
��"O��MEC��0Pch�$�z�"O��x�b�l
��n�7j^��W"OXQ�P��*=�j�[�ʝ�?�n`"O���iQj\釪L�����"O\8��l����1�̘����"O� ]��mE�v\�'�Hg*��Q"O<!���0z�yK�'����]�"O�x;*�"ڎ<�æޝw��I�"O(<h�`�=t p#@C)}����"O�1�&ME)u&M��ɋz����"O\ ����4;���2)V��4�bR"O������{n�1q�ǖ�ɒ���"ON�$'Y�S׈�Y�I�P�"O���h�2H,� g�� ��9"O���@D'	f$��� #e�K4"O��d�("�$Bܦp[±qa"O|�6���T��܁.ʵ��"OҐ���*H�9R�Ɗ�e�,)�"Op�9U'W+.�z��.%�X�$"OD̨����K聈��X�$�p]��"Op1�iD�NBjԐj���t��b"O���+�h�d�Zd��zͮؒ�"OX�r��M�b
EC�T��"O؀9f��-l�T�P��2q��7"O�0�B3�x�%D�&'�ۻq"O����%`�9��D�V�(�Sg"O\�Cw�R�7)N	� .I��Xpv"O����e��w.�QA�c\
+�n)c�"O��y���x~,�p��#vZ<��"Om9p�E?K� �Qe�������"O��
��FCX����i#"O�����=Oň��ҧ��#�"���"O�M�qe�1.D1ŨE�J����"OA�֩� �����'Ϥ4<i�"O��!�f�t��C�v���2�"O�,� o@d��gERfe"Oj���#B�@ȜN4>�J "O��Y��O@T��P/�� L,b7"OȔ��ל ��9�M�8$��"O�9��J�2<��ibBO�-ƕ�"O�,#"�ˎ./>�� !!`%<pP'"Ou��/�"DŘ̸۸v4 �!S�%D���f.J�Ry�'nE�E�� I�+9D�H�E��"[.:tc���p�����8D�8��ڄzв�s Џ5娼1�#D�̢4�L�&��(��jM?t,8�х�-D��Q��NT͸@�jM�M�A���*D�@�m�6H8������')�����(D�`��2B�JP���Nh6V�R(!�՗���)E��8I�����:U<!�ڷe]8��Cc�),3N� ��� {5!�DZ�\�� �ү;=\X�s熪,'!�1q0��ID^�w�E�%�E�E!�U�A��́򨋠=��t	���*8�!�d��h�n��p�׃>L^�
�g>9N!���b\X�ʍ(4>�в��7<!�dE�`�$Ŋ�ع4�\��+BY/!��@ix�0��m�����D�
!�$]xh����K���X��d$�(,5!�$*nh&|��Fԕބ$��c�#�!�dO-#�P(��X�P�>0��]7L�!����%�@�O��E�5�Q�Jk�'g�m[d�B��|L� �����y�'�����t��\�&R*����':�EC����j��pB����9�'������M�t�KPʒ�~��y��'T8)9d�M�%MJ�) $�*}̢���'c� �/�##ۚ�����b�L�
�':����A��mN�Ez��S"��
��� �M��!�>(�$���:�(1"O��$G�w�~q�P�V(��H�"O�ȡ �ܳ)��eXs�
�#ƚ���"O�X���~-2�r@�O<͚S�"ODH1�>j;��E'?P�A�6"O�A��K?J�F�z��9F���"O �$�ۗN[�P.�t9�� p"OX`�$�(��wnL�'��t�W"O�xH�j��zX��3�1 �Xc"O���FB�%s.yK�g�:%�J�"O����S�YP�p���/i�~ @�"O�=�e^	���ę�0)�u"O6\�CO��[ǃ��l�T��"O���G Һ	�*M* � �h���!�"O�}�6���&	K��N�Ds"Oj��mWR�lX�J�	���"O��Q���}ư[�S��02"O��1U#ݹ(�Y�/˘5P�1��"O�RK��!
�P҇Εn?�<��"O��Pc	   �� �   �D�8�%.E)pڄ�6ӗs����3D�@
�H�B*���ԛ��@Ȓ'.D�!�J� D�\���IҎ7�D��#*D�<S�m�U�u���2C��P�<D�0�~P�ۂ�T�%R�m��$<D�����L�$��PS����s��=��.D����G�afLbC����~}��&8D��3L�+0ٻ���2��ZE�%D�� �v"�6^ʲ��"g�2J4`s"O���↽B��|[sM�d/��
�"Ot�B�̑h���խ�AzH=d"O���B&$T���C��݅1W�ո�"Or@ǅG�1�A�j_�sI��!�"O��"���y{��i�A�]�XER"O��ғ/ًD�Ѕ	�-a�\ܳ�"O�ɂ!M�';�`�aG@�>��"O���V�
���F^?8ל|�"O�H�L�@0J�9�F�}� \�s"O��ё*X8?� �S�Ԙ'�``��"O�!(�̚�斩��J�9O�Ti�"O�,��oҺ:��Q;�
�%PBA�d"O� ⃫�a�h�zv���F���"O�r�����H(6��$�T�xE"O�H���c�Z�p�O��Ȝ�U"O��vc�#)�2�I@Nۨ�,�*�"O�!����$�M�#�ʓf��E�"OYhA�4t�G�\�(����"O�踳잵4��ˢ�
�[�Bip�"OR�"��Cx:�,:#j�1z�-A"O�4+dM��W��# >� u+�"Oʈr�
�(kX Ya#=��('"O�|zf�A�$y0��;%�1"�"O�����=��+T��>���"OX��a'b���b�&џ?�s�"O�� N2���T��l��l�"O���.��yG��W��Nu�I�"O B���2~[:����:����"O�m�&.����B�ÊŪ��r"O (8t���,P�P��%n�2��p"OfD2R#�;:0�K�$Ҍ���h"Ob� �)ڕuD��dN�!���P��'�d����Fih�
��:K�P@�)Y� ��C�Vo�>�"
�'k\��"�'F�x2�fF9mV�
�'�`u�v*	8P��p�۸`��92�'��}��.��f�k�e��=����"O聙N���6d��6��|��"O���5�Н$O����	�YXP ��"O��Ad��8)���Bʝ�"O�4;�#׈$f �A}�dt"O��I	�\��bʙl]z�b"O`4�4�}��hd��=\�q(%"O���N�g`�jB)M�M��	Xl�#�� ��h��M(L��vI�f�=E�Y�=	�ib>���'l:A��Ϗ�D����J(#~M�+O�$���+�V�$��|�ℹdx��1�F5v�UH'�ڟ�C�G �nPkO<E�DeL:�����1c&9�Ȁ~U����Ϲ���0|��I��z{�(�s`؀�`��$K�f|�<�pşd>���'�$3A
��(Ǉ'xN@+ 2�'yLD# 2����c��CWj��Ԃ�0$�n��C����E�aI�c�"|����MBeS`#ʆz��lf!Eަ}�I (ln@�H<E�o7s�8fgԢR��l��ԟ2�Dt;7� ��?d�>��'M���`R#��P�WF�,3>,a�T.N̓3?.e���b�t���k^�:�
���Q�C@FB䉅2�D��a ��gFc�/§*aBB�B��A*�:T�4dq��[�D."B�I�l��<�vGU�}�T�$�Λ-pTC�	.1p	�1E�Pr���7�K�q[�B�I� ��BT�P�h���H�n�C��B�	��v�3p�J)Y� ��g��ZB�%dP�p���؃% d��`�(n
DB��f�\I4�Q�x���G�U�� B䉌s�QT�
"˨�!��WC�^C�)� ������ꊰkWFY�>���Iv*O������,�M�H�;0	>X��'�m�D�m���ӝ#5.	#	�'�j�r�	�ۮ1b%k!��ؒ�'�����C%�,b�吥%o� ��'բ��w�.�MP+_��\�h�'S��ۧa�;����$I�
�*�'� a���>-Eʰ $Ȃ�LY �'�z��^h�1(p��(��	�'n"��C�؂P�x	��l����0��'&Ց�ĸ�~�{��Ζ��dp�'��8�1|�I�c��9w�i�'�t5A���/$�8j$L�0H�3�'���h���;-
��4 ",}����' ��g
$FKdy��/I�(��l��'�Z�pf�U�ɼ<�3[jB�!��'�p1��1�.]�GM�5��Z�'���­6x����$��3����	�'���Y�N�a�Ѧ{�A	�'�$�T���������:T"O���We� 
e2��CȕK�h]�"O�!��dù�2ѸR�M�$P��z"O8=��E���°I2?45P"O�y�w��y\b�*�IQ�4D���"O�`I�6;�C�F�;E�pÁ"O���
#i�tUq�;b��1J�"O�����+^�V]��H"/m��$"O�U�Ф�<{�Fx�vB��R���"OPD-Y�{D@���!��� �"O�eXq��(vh��Bܦ�|y��"O�+��͎�����L�u"ȔB"O��Q�γ'�~�B@�"r�>9J%"O, 8�IY-o*JS�[Lx�Z�"O8����߀��@iX�[e�	�r"O�q@5�1=������ܔ^j䠫�"O�I��m�\7`ŹFG B$���"O@�"�� �2��U#��]�U��"Ob@�eڸ[��`���M��h�"Or�rv	+Y��D#Ȟ!�Z�X "O��;�DەD��e���/'kjDɐ"O���6�>4:8&�p��up"O��;�k4W`��FĜ���"O����+]�{n��ql�Q�B`cQ"O��"&u�������b�v�8F"O�%�C���qL��2sC@�Y���S�"Oș�ƌ9X�n)��O��S�FQR"O�|�4-
��RTꇮ����!�"O|)®���U��P'#���"O��	v�٧����dD�<npɸ�'^T	dI>*�P�j�Mž)��S�'�D�T��H*� ��	�#�t�9
�'�bձ�hP:c�Ta:r	�� �#
�'�N����F(ʌ�C��V�����'9����\Lx@R=H�y`�'W��b��>I�#W�Ŗ�U��'���q�o�8F@�&F	*Q���*�'��%��	FD��lcW�K�?�Z���'�а�UjY����{��6	��
�'�V��p �"z������!F(ec�'��W)з<S%�$�Z+k�'�����F� |�:$
�e3��x�'ֆ�	'��3L�q�M^���9�'��t��Ɵ� Z����	��-�H�0�'��8�0�׻6<� �n\�V�r"��� F :�aܚn�ܐ�w@JD�)�"O�-��N92���!q5��K�"O")&��T��$D̆ ���f"OIB��@)�M�1��
F((��"O���u�@=;�
��_'(��"O�1D錣52m��,��`��ۦ"O����n[	<-�e�A��Z��s�"O,��ק�2}�pT�&�Տ�h�""O h�"K�1bx���!�M�Dԍ�R"OFah�gE�|���	��ı6CLq�"O��I"�R4j���Q��%��t�R"OZM2b���d�J�(^�&���k�"Oh�1/.�j��*'��3G"Oi a@�� P'
����y�"O�\��?z���uƅ<l:r"O����.wY�dz%����}8"O �vΔ�td̀��ڢ���R�"Oxȩ�%F�YbTZw�S�K�����"O���'�įpq��3�%Q�~y��3"O�D��i�$̒���*l[�"O��s�
$R�
r3h�"O�E&�Y�7�������3(=��"O��2Gֳs�P�J#e��%"�D��"O>�*C��A����&&��"� 0E"Ot�sb�I ��2��5�Ph"O�Ү1R��3DQ&>f�"g"O�ѳ�![g�<pō�'�V��w"O��j�S����C�8o~ȡ"OFA��P�4�(���J��HW"Om{P��bϲ��T��["OP�X�k�%w~��Bh��zV��r"O����K�1~�%��:@p�"O�@ֆ�>���U�+74yZf"O�q��	�v�( ��l�;,  ��"O�<���f�Na�u"àRp~�`1"O4��֦\�~��+� |h�W"O�X�t-�D7��9�^�c���P"O�u@R��CZ��`(ׇ��p�"O���@�:4����P(�v���6"Ov��L�0a���gI}<����"ObmR��P�S�R0���8u0ʹä�'�O ���6%�� ���f�l��'"O�@t��"Bd�y�SFH<[㖉1���'�S�'9�Hd�h] \��x	!Z	'�|\���nH	��}����WEx��>Aד5Č��A�Pw#fd��Fڭ;��x�Ɠk{tx@�n&Z���(��Q��'���ڔ#�7��-�2ɇ8h6"5X�'�l�KK�`L�pӦ�J�(��'�>���	A�5�vT��ߓIӸ���'C���h�3.H�0MrM�'�tM{�*ˇk~]{�DEF��(�'|��0F�Z��2�@�E� *�'}��$m�Y�Ël�2xG��y�	M/N x�@�=d>f��v��8�y��\<Cgj\3�O *X�Z$����yRœ:��IV&L�9�5�1�y"ʟ4{�85���F�?�U��&X��y�.��;�]�3Ǝ?2��� ��Z�y�eV ����#X�0���4����y��S,�A[g�X1�E���B��y�+Q�j���c�-��[�R(�y���6sa��AC��Đ����y��>U5���
i�,&���y
� P�+��
��F�ۇa�,(&��'"O�)S���9�l) �/�^�2	qD"OTbe� s�X���1��I�f"O"I	CDH�A� a)�
b~���"O�ԸrNϤt���b`Z�Hl,]R"ORYq ,Q�Ep4!�N,)�zɒf"O��8�A�Q �ja��Q��hX�"O��[�ASl9R-���*�&|Rr"ONQ��.�Z��$,�f�\m9�"O��{���f��{��ݣW}-�"O:��� �>�d �sf��XjR�X7"O���!Q.���E�BB�Q�"O�ՙP� 3@�����L�R%�0e"O��S���k�~�uG�]����"OD(`�ǜ5Sk���P�D��"Ob̩�ʄ|B��D�'l� MsB"O��8�꜖ %��QUc˱b���k"O� rq'Ž�f��fB��"x�|r�"O���ĕ'��p'M\Y�T�"O��q��|��QP���[Y셣�"O�q3���	Dj㨚2 TV�`b"O�p�SI"n=��`�m�]�1�5"O&!5FҺJ�:�*���t��"O:A�0H+Wm"aZ��[�I�4q�p"O:���I?���QQ�H�2Ҁ"Ox9ˢ��+V�ܔq&EU-;�F�J�"O�z!�y&|�G[�l���Qq"O�%pp���7xq�A��0YB"O��9�!�&Ɔ��ǥ�rH�`�"O"|�@�f���&? 6fl�E"O!��7-:�禉�l?����"OƵ�d=C���$�i�l��"Of�)�E�#FY��å	I-�p�1B"O�Z���]>�В㋧5؂-qd"O8�B���[\��DZ�p�b9��"OdP��	M@ڢ�s`/�b�|��"O��׃�,; i��-�1�.�q�"O�l9��]��d�Y�v �z�"Oֹ]�XE M�x�p����W��!�dF, �*���"�l���0x!�D� h���)��W���b�!�DʠYB���#"��)&��i�Ȑ�<�!�d�jV�p0ğB$
�������!�$�8ot$�S�*��h(�o
�R�!򄇪&�'�8��D���(�!��&ʬu��F?!ԆQS�̞�j�!��E��}�Gգ'Y^Y8�0�!�D�G���4E�1I?�L
7�h�!�D��>4x�Z�^4t\y�P�D�!��#�)iVCǔ+�@��J�~u!��+$Yaŝ)f<�桞=QY!���I�ŀ �I1x���j ��m�!��цt�Kaǜ]^PlI��ڋG�!򤚙WAv�@���z#`���µC�!�$b��ͺ��]�;�n�1�!�D �Z��k�MA���c���%�!�$V��QXM�7[�e��a��G1!�Ŏs���X&���&�:A B�!�D�
�@�@���Gsn<Z����_!�X��v	���ݺG�U��-޿i!�@ؒg�_�B.H\��*�U�!�$�o������X`�4���!��?Q� �  �!�r;���d)7�t�"\'z��b6bl�#g��/;�R�SN�F5�g�(O���2�'����	��� ����щY�b��$H$��3�O��kVȓ�@��0`s�G@�x���'SN��R~�lXƨ��I0H��kQ>D�R��T"�.�Ms��?y-�9����O�j�$�)7(��v�B�_�F��ǀ�O����_�ℋf�0iJb��@�V%��O��ӉS> �����e������^x��<���Z�>-�|�Z��C`z p��J�(A1�O��u,��c�-�5��A0Yp�OȈ[��'�:�O>��&	G�);8���g	�wM���!�=D� b��ŏQ(`��f�ˀZŒ-��;��h��>y	1J���m��E$h�g�	\s�6m�O$���O@�q���'�����OJ��O���$l�т$D�������$W��@�C�0b �#�~� q�0�Y��1q��`:QN�/Ѳ��&Dݺ�ƅ6�û$Ť�aQ
�Y0
�1�^�I�UY>) NN�?��赯�&(�N��*?��k៼�����?���.yj,l��a�,#���y2���5Hj$ r��5[D�� ������B���t�'��ɑO��C�9bz��,�W��2�.Bʟ��	�|�	ey��DȆ�2@dDA� "0�c�Ʒ2i�Q(��˟���Kp$O$�����;�� ��xB _�ED�][G��,Pah�0�#ŗ7k>"�.A�d����7K�A1fڌ\	DQ��i_R���"�'R���N�'y4�X�L�H�"�rt�J1'���
�'����fM�},�B��٤E<J>�c�i�U��R�l���)�O.A���:y ��h�'$�	�+�O���O4�����OR擮9*�00�>4��h�ȝl�FM2_*,�� 4>lf��t #O����.��	�<�s1FJ=7w����ƩC{����㏗hʖI�3��,Laxr̍�?������_.,Z���h�49�1�k�'�a|2j[C��]'b&���c����?y��'�¼�i��,�B�M��'mB<����9h��m���K����"K�G�FpQ�I*E��l���Ω���'8�gO@�hQ&:��
|���tg�q�ɟ(�R��Ȭ[+�4����0@�Ƙ��j� @^�	G(�jڤ�6L����O~c�1��B�ΖD���z�O����'�r�S�<Y���c1�A�hV�p�������<	�Q?∸Y��	9��$"ÎW�'��}RU��S��
�����$�4�Ѻ�M���?��k�&�[�dU�?!��?1���y��Ү0���@��RHa�ۃNh�s藕io��H�K	�L���t�icJ�z�'�jM�VӠ hne�g��9.������1^�썊r�X�I��U:��٩��O��6���~Rh�?~��B��P.v�|��)�?��O
� #�'D��'��O��'�:=��X;��1rl�d�%D�HS!燋�\"�J�s�B ��L�t}�-��|����	9CF��r &��q{��­ �z+�����a������I^yRY>̧2���� * ~b\[��!{����1	򺵡�!�&E7�!	� �f)�c�Y;1�x@���2
�0�M�.�P5`�C�1��0`�З"�(G|�E�`��ɐ'�	��銱� �#'��x��xz�6<��O�,��`D�R��d�B��H���s�'!�զ(:1�����<��s�פ��'7����'���:�Aq�H���O��X�\d�-�c���$G�!Q���O�����KL��O�)kb9���˓$3Z!!��]��M��PxBNIb�.҈��X�g�_��j��dж��u��'	 pQ�qL|��g@�iC
8���7���(�c,�l}�����fǩZU��x��Ӱ�V�1�ȓ���k2"�t�� �sh�,,��	�?Y�#��+2�����@x*m�G�W���t�4�?������$��$�|
�4(�oJ,r5����!�>���O�U0w�_�V�p�.Kx~�a�hN�Đ?� ��
�jGr�	�J�+v�8� 0?)1�R@9&X�r�K�(k�\�ǋF�uG����"3X,��۴9���Q�v���hq0X�'����	�Ct�	�h�Z".�Xr.y3�d=%R�'Z"V� G{�L��!���p�g8r�� wB�)E'� J���?Y�R�̕'!���
i�Q�����	���X���'[��''��35�e��'�r�'�n��<�0��f	�H�jx�個]mι�`H�!S�؀(��B�ki��ؖ���//�DO�}��� �1#��P�E䒑Xn&����6`΄2�ITd��B̧{��'7�t�Glޭ(�H�[�ȉ W�I�@�i��7�O�%z"��O�c>��?q��#s!����!v-�@ǁ>�y�R�r�<@A�c�%z��0(8&�����M���i�'�z|q�O��D�V!����K���hWx0��\�R�I��4�	ן+XwW��'m�	��H��l�4��y.��*�j�%Fh��cjC-]LVA/$��!��'K�9+�	�	�� �l�%W��xY4o��B��S�^�.
w��:��$�"\�HуV�H ���" &�v�'Z�D�'vF�9�L	S�zE�%�\�F�l�{�'��9�4�A���yB��@���IN>���i�]��ʶ�B���I�O��ڂj�$�"���U%I�БC!�OF����%x��O����R@�<Y@2h�@�A��TP�B�`�`y �*RP��<�a*O��:�-��D�� �� �{>�(J"eԘB�8��#�@<�j-���&�Q(���&z}����O���6��!�F�>���`���i���'����ɟ<���AZ��� Ƒ���' �D�/��!P�(#$���Ҍk��^� ��`��MC���?�/�H�����O�`���^R-"G� � �����O�6F��
���^�9F*�ۦ�O���!~�yꑵ .��g��P@~r���0�F�Y�ʁ�!���k��S �2�3c�;3���ӵ��B��vg�5�	��`3�4�?y��Ɉ� IXp��#6<�(	�FqrY�����\%?�d���I��2��OTeT�$�g�vd�Fb>M{ f�.0�ԫ���p�("�D���E������ɷ7) �(C��ǟh�Iٟ<����۠L�)�M�ֵi_�y&���x����?�M��	F��*1(�$a�?f<�z�g����xX�B�*Z�@}�@�ÞF�ƄU>�I!���y
� ��2�˪Uj� �1��cs����`��4m�ڟt�p���,�|�'���B�&��tjV˞�Mx$���ΐ�ўt���K�:�G��8(�}�¡I:���#���kӞ�O¸�����˓2�`a�� �H0Q[�(N%� ����O�Td����?����?���6���Oh�S#	��Iڶ*�GlZx�T��D�	�W���K� =0����jנL��46���T�'��4��R �A�$���r�nN�"�tQ2��31��dCp�G4�M�%F %�<��Q�K/��фhIc�)� S��4�����?1�	Y�vJ+O4cj�0���I�<����N� ����ۊd�TmZa��B�	5�M�L>��-�0k7��':҇VG�,!�2��V�^�v�K�c���'O��	��'��9������'�1O���1�EQ���j�C(8"hˇ�'kL8k��$I�m�����ӝC�p�D�2ruax"�0�?-(�'
� �f��,w`��C�E"�nTB�':&�seGܙ,>a�3M��cp��
�P�� H0a{v��IU*Vʽ������I^:l�Ƹi\��'�S7njm�I�:E��Mީ=�)�LԬ���	̟���g���M�'��u���m�$[>Ũ���D�<˒���AmZ�*�-�w~��/�\���V.IT�HD�d-L�L�R�z�v��9����#Sb~Ӑq'>��|t��Y��{�昍R^,wMzy��'-|2�	�{����/ܔ|�J�kb��{��#<I�O�mZퟜ$���b�6N����H܃Rq�A�V3�M���?I�DiX�[w���?I���?����y�ܡRUr��-�����ұ:����X-��A�͌�.%҈��m��=����w
���'-
�Tn�p�ƛE{0�I�� �M���`f�8dTm`���B�'T�)W���P`dU/B<���D ����D��Oz�Cb��I���F{�������(�� {���Ø3�!�dڳ2*P8���hL������剿�HO�)�O��,,j��è��RPtAiD�vr�}�w��#:m��@���?����?�Ӹ�H�D�O��b�>@ B��-�(Tj�J�
�;��]2 �Qس+�|��牎rD����z8&�Ĺx���TO�+
��t���̛V� :��%w��">Au�Umu xk���"��v��*Z �	��l��L����܁'���|�.4��/R)DE Y�"O�Ձ��0V�Vy��a���A�|b�dӤ��<1aK�-p%�SΟ�Q<3�AZ�*H�j�� ݟ��	�eŘd�	�P̧P&�;��ͭ4$�l1&-WMI1�S�;x+��w�d7D���OH�q�*Y�{M2�R aTDB�%� I~�����f�$��3�
�dJ�?iG�˟8��R~-�3W2�U�W�Ь��ٰ��9���?��8el�%D
~�x����K!:z��<��T>Uz�E�LjR��t�d9����!e|��	vy��'�6��O����|�qi���?AT��mn��#�B�'��`f�\�?��k��Pz�,�T�(p·�MKT��~jΟ����A�$B0�%طP��X1q��0Y`LX�XŪy�a�.(C�6M��ug)���S68Ȭ�c� �sS�A"6�:R6�.�p�I��M������'��0��t"����s.&TC�����|"�'�azB��M)��`chJ)�$�IC�\�hOn���u}��	�#h%���BO����x�0�_3��7��Ox���O@�G�p�R���Or���O\�]�G7�����D��f��T�l4B�y5�ׄ-��8xI
%~��U�E�9�~�I�Fܖ[�K�W�.��w�V�O���j��Ĭ��-�&Ɏ K�����I6�{�Ik�$A+��.�5{Di�"8���0?Qƈ�����֟x�?qr�D�4�8�u�ɿbbP�ac�Ɯ�yR��	8FAj��ܾ^�rL�k^���D�a�����'n�	���Y2dl�=���G�ߟD�z6A�3��x���,�	�P8\w2�'+�T{��i����٢�A�֊2E��9��G�6w��c��e�@B0��6z>`H����j��1a�������G��ۢ�$*}V}�Co����OD�FO����Y8B�!
C͆�ab�'#���&�'s�"��{�9���I�'�Nԇȓg��2��ŕjed��w%��y�0y'�ش�?).O$� C�X@��'�)��h�y
G
J8_}�0ò�' �<v��';���Q�pbf�F0u�³��#q���Ebِu����IȚV��! 6�L 2���f�=K���%�o�Q��BRv�h��!�H0��6��OE���'�B�������
�(p��*"��4`D�8��O����� h�MHUO� bT:M���R�Yc����OH*bлAV�����=h�쳗�'�	
r��B�4�?I����iV�J���dI�X�`ч� �y1�h�I�b���O*|�4D��z�L��a���o7��@Ăx���?�������A��+t$8���!?qC��"J;��A�C�y^\���ڃ��O<����R G����.ۿ20��OtE���'�����`� �!�U�=��Ր�䞢:ׂ�r""OLp�ċؤkَ��!�D�H�$r�ɐ�h�ޥ�I\(*U���n�5"���}�6���O��D�iƨ�K�O���O���k���JH$^���'�.�t}�'�%�N����O�M��۷v�b>�'�"�A�����V�.�|���Pt� ��S/h)��N��&��b>�'��d
�<Eĝ�2 �6s��A ^L�ɧ4s��$*�3扅#����`H�pv���א��B�I�w��Ã��>R�6�+�4F0��Y���F�	�&��a	���
����1���&G���q)�)Ôt������ϟpZw���'��>o7���HY�[\��#��C�Rm"�Y�������c��p=����K� ӂ�O' T�JscRV����f:	�:�Kѧ)\O`����_�p<��@�#� 0��	F��Ц�Kٴ��'�R�?Q���A�R"��#��5ߢ k8LOv㟐;��*-��H	��̇&jd�Q�B5������qyR�"D�7-'��HU����z��#|��ѐ%j��7�9�h�Q:���L"ܩG+�4إ��	0Kk�"<q��A?i�t-�����	�v��Z(]���4?!
t�Ë���X�,��2�!��/m�Pȃ��?�j�����'1t���O�a��I =�2���։x�`�H�|��T$p���	��$�|
��O�"����S&!���� �R�;������?�r��>�e�PLZ��O�_~��I"o�b��"��5���M7O���	��Qꊃ~�J�#wk�u�Oˤ�R��U3FVy�ԫE2% �O� :��'/"���<AT�[�t��-�QAÓ��E�6�Bj�<�сٙ0j���8\*����f�'�<�}r�	�b�G�Y<甌s�i��,q���Hy�#߁n�B�O"�',�	�t�cNلw��9��E:2���*B%U��F�A�"6Z`��v�g̓ɖ�2���Pv��c�߃,T���nP�E�X1�.6����u�g̓IYځ�Ю� �{�T�2��OH�t�L5���TF{b�̈d4��q%��P�����$�.�!���\�J ��7{):@��LY�Q��I��HO�Suy���^�Ș�➏O*\(��P�Xo��

�	��U�3��8=,ΐ�����J�dl�0���fM�.L��аQ��Ԃ��8�u��7%Hb	��>x��'	���k����bA�*���w&�Xֵ%ṇUdjU�"׬�@�3� �!?��+��DˣX������$2��!2�ҡ��8*!��~�МX���J��XB!��9�E���䜴I���'�1���[��T2̠۷JB� ���CS�Є�I�kL&\1�Kן�6Q��/
�r����~yR"�����8Cɚ�VsPe�1��+��$���J�m�̟�	C����1
"��'M��6C��h��k�HԐ��Z��6��n8	��N?����*G�q��!�FZ{�'wN�M+�)RCA��-F�H��D̓
�
�X�Bկ8��P�7�ȐE$�1�f,��>=�PL;F��B�#_�@���t���cd�O<1n���4�?�Re�z9Tr`�p�A��6D�������t�E�ʵ`s��S�B?ړՑ?YA#i��?`�Q1l� ��P{W�}����џl�aH�'���	џ,��D��՟P�(�
*��}�Qh͞ԕJK
1��q�м�>�)p�����4�Om�&���I�B�Z�c��b�"�r��1��I7�^hQ��Q�G�V�r@/5��4|����Oz�pe�;�=��-��S��Lc&�OZ��2ړ�yZ2�TE�R�F���R*�ŖY�ȓn2���p�ݳh�a����(�b,�I�HO���O ˓8b�u���S�U��,�t�ٮ.Ʋ����	�@�����?����?)�'�?������ 8vW�%!6����,x�XJ��*.�3�e�I�a�T��m=�X��<У+�|<�s�#����Ez���'B� �c�#`]��sR�p�
1��$ʓ.L��I�~���ʄ�#��H�ũ�R���b�'��t�3&�]����e�DqZlQ�F9D���E�W�>�z0ã�=bH(�r��<6�i1�S�hk�Ӱ��	�OP��+8�1�A�ϖ;~���#��,T2��^#-�����O�$��2L:���L@�+I���#Z� ��S3aZ�@w Ñ#���n��#>��1%�N�	qFW��1�J��u�͚�dC|�pԧ�\zB����N ko~:����Sd��'H1��T@R�N�s.zt�dGK,�4�Jb\����I(���˃�/�ڠr3�Z�l����RyR坧J��	���?]#*i�J���-e�v�l���	u��K�����'��*`#�?^0,I��7�|���'&"�Xp�N�D��\�c}*�`c>�#񈕵v<%�K46e,���Or��#����*�b���"���S�8!"����	7���C�h�\�&�	�Y�����O��S�Sy~
� �q4`�Zn(�h�#���.|2B"OX��gꐚ'��9��듵�T���퉈�ȟN1��%��z�tH�d��A�j�T�O����O��pԌ֬v�����O����O`ɭ��?�f��4y4�!�d��V�uvh�b��H���hH큥`�V�$!͟����R=�o`z��.<Vp�(�N�e�����5Q�0C���!��aUi�b��4&TTL��+�I�*�)s�C�!O�0���2?1c�Ο$�Ih�'��DS*:{K-_��A�_�����'B&�2�g�rܬ��ۻu���'��#=ͧ�?�)O���҄�?ux��T �����Ĩ >6H����O0��O(�S�'���,B�)�X7�Nr������:��Rn�zd�Ģ���<�SD�Y�:���;P�F�*�mДuˊLr G�b�~-
OY1��<IG؟�2@ΗL���9�֖
��y���V矸E{��'����[�;�6�3ů�Y�B䉭i&��LF\�6��Z���TS�4�4�?*O������A�	ß�ͧD�ZD��M_Q��cGER��I-���������Ig��$Ђ-�{�*	:��
�|;�(��	�+�ݏRꎸ�a�-#�D|B�S.C��)��ъs�t��EI�4�!h���V��$(y�ŧR���O��!D�'>����I��<1f*	����"�$D� ��O2)u�8�����/-��*�/�Oz\�''���4,:dE��d|��*+O��d�O �O�Sr~rœ�T�R�+����/� ���fɃ��OPaF��_�#����AdM%bh������'2�6�x�!R��#�������B9� @��,�4�Z۴�?�r�V��yř&�?���b���y�&UI�މE��\9|ڇ���l(
�$�i��./��=O԰�՟�^w����[�H��2�Ƶ�ă�m.��P���w����O:(��k���?i������y�Ԇ����2�Q-tf� �w�ƗaPJi���?�eH��?�'���!��M��`��F�M����\#��b�G#_X��$���6�O��P$K\�$�'M���yr�Z�[�|�X���Dqx�w��g6��$�e6��'�mQ�'����E����umh��2�$�.D@�	r�j���i���$ �r�'��$Jg(�~���?q��BI�yBO܋ncNe*7�F����2�D��y�U&�?!��JL��O��	$"0@��Ǧ���ë�,[ťڑS=61B��B"!�:����<)c��h����b��?9��~-�%�GYH���	�����U�i7��9O>�ʵ�'�B�O��9Ov�s1;���OB<~��LXlR05�*�Qd&z�D]��O�˓-��D�i���I�<�S���hs�n^2�8��c��*t/�H;�'��h�Q�#]lٸ�E��xLV��ݴ�?���?q��?Y���?A���?���SS�Y9v�6�p��޳1�j�C�+��e�I����	ğܖ'4�'"�O>@*�j��Z�-�q�[< �l��c��\yB�	��$RQG� �f�S��4Q$7-#���O�H�~&���@���3J��s��@�v+��i���>1
��$ZZ�y$kD�Dv�c*�=*,��ȓC���B�C�Pn`ːoǵB�j-�ȓM�6���!NfΔʃ'	m�h�ȓR��@��\��nE:U �s*恇ȓH���`�ڸ�����{עх�<���&����%�>�,4��A���$̇{2��C iưT��hb.U���4�l��#B�J�\E~b�'R�'��'��Q;�I��,��zX�qnĢR�6m�O���Ox���O����O��d�O��Df����Ҹlw�){�����l�|�	����IƟ ��럈��ߟ��ɳw�-�r��d��pk��M����4�?���?����?���?1��?��{R�v����CO*r|�t�i���'���'���'OB�'Y"�'��{���djb�+腉ּ����{�6�D�O
���O��d�OL�$�O ���O��(f��(`o
�xgI�j�@�ʴ(�ަ��������˟��	����IΟ�����pUĕ��P�{�,uM)E�] �M+��?i���?��?9��?����?�R��%��@	e��9����Eꊊ4?���'�R�'�"�'���'��'�r�"4Bp����O�&�H��Q�e�v6-�OH��O0�$�O��d�O�d�O(�d
�>p$,C��	�eɇ��^3��lZƟ����h�I����I����I���Ɉe�8���A��J��<��D��e2����4�?y��?����?���?���?Q�]t��s�,�8���@N�W�v�1'�i���'��'���'@��'���'������R����q �a8.ɣ�KxӞ��?�,O(#~�#oY*��3� >U�hH�RC�!�M�DCC���O�$6-u�H�7A�Q��52�[8�,�u���0l��</O�OdΜ�@���~c��#�\��⃠��q��肌�?�bϏV'2\ˁk��hO�z���5(D}V	a�@F��|�+Tg�O�˓��o$��I���'�� LAHG�B�Y�Z�S�\_T�d p��Myr�'���6Olʓ|�4��ƌ`�~��u��N�[�']����#šv$2���O��͋@�@t�f�h�� ��է$��k�Ë
�"��$�<�/O ��'�g?��)Ӿ%�ȠqBkL��e)V�P��4,#���'֦7�:�i>U#1J[�S�X�0�D��Ss�Ѱ"�W�<1���M��F��Wb�b~B��(za��C���#9z�A����]�c�Xw�'�R^���|*vo$[E���R �%+L�� %RuyZ���n�ј'��ik�/��9L�!P�M	:9�m�QB�fyb�'$��<O2#}�P�jgdybƌC;h�ިJ"�1�0�&&�s~"D247"=Ȱ͌,g�ў0ӣO��X�.��t��\� ���󟜕'2��s�	�M�K�|?`$�Y�ʉ�6�R�1�d)��v2E~���泟�����͓T%t��c	�O�۶E.�0|�r��8�P找m!"��V#ި�Sڟ�^wf�L�Pd��=��b!`p�[D�P'd\$1b�',�Q������@i7K�M�.H�k�^|����|"icӘ������ڴɘ'���)�8y���)�lП'���æx�4�?!��&4x���~B!�gT\��X�-�r
��)����a�L��O����R���69z,���CA���䓥I�����B�	��M�¦@N̓��iil9�3��D{TE��	�|R�	���$�O47�a�,'>��S�a0�Jrk�x^�9(���!pW4�I�C�0Y����2?i�'g�,8ϋ���'c�1�D�̸u��\�nɺ@
L�*O��ľ<�J~�'q�6��Szm�3!P"@��Pa�A����ؤ�� �ش�����'1���:vQT����R$|���&�'�6=#�k���yr�O��#E_�VB|�'�}h���Rʎ$��D_�G��`i��'��IR���� �w�6�9#bF,*�^��&Iզey�o�����蟀�"��if�DЫpJ� `��q.�IZ�&7�ͦ	 �����\�i埶�J�-���9�� ���Сq�xř`���V����"t�%�W�!ĒO�˓��OQ�@dHbI��T�2 pT�R,@�џ���4SҤ����?A��e�m���9ɸ8�d�G� i�L����>�4�i��7�Sɟ��O�< s刟0_Lt�J��پd��;���?��DV�6�@.���D�4�a��D�L�	� ��2�cu�t�iJ�0B�I
�Ha�@H�ha�!���}�B�ąڦɉC'�ퟜ��9�MS���O*l���-���� >�@i6�'�`6�ަ�X�4>{r��p#��<������A���c2�h��#Zn%Y�l�3.����&���.R�{⨙�@�1�1�©we��b��<�y�]�\��`R䊙wP�(�cbN�W�=���/*���Ǵ%42���'�x� XcᏓcx����aI�o��qa-��Qu< ��mX>�&$"��Յ4��ɹ�A�Iˮ�a�A%Ot��(��}-�`;uo]4�v�b1�ҋ(��)yW�>?p�����	6f�"��\
 MD�� &S%ۖ����/(�`��TJ��q��")L�c�[<u�Q�ӌ[k�pQ��: B�i���}�v 
ђ��a�P$.���y�[{+���ϝ3N���Z��ae��D���)p@�F�L��@�^$�����\�,ȁ �Ώm#|AIaP��ei�B�~��xvC�J�<(q.Ȯ,��%�`V^�sB�Ę$�Z�jR�
(WG���&d31�\��+ä8)�P�4'�|n.`�ÉÒ0�
$�Q��>/rz$ ŧ�<ξ���DI�!��	`ѧ�¦���ן8�I�?�IH<�'*
 t��D�(�nA8@H�&�X���ax�Ԃ*O��d�O����O$P
�%}�ʄ�d��fx�hZsL���	ٟ����1�i�L<�'�?ɞ'��	B�>k��Q
�L�!(@�.O��y�ư�<Q��?Y��Dw��u�F�l���_|�y��̂ן��I�<pdH�J<�'�?�����D�WL^\@D_�<��7��)����O���V��O����O�˓I����0r!$D�'*�5jl���!�#l�'��'�R^�X�	ԟ�B�M�C4�	�FⓤlN�HcG�� ?Hb����̟���`y¦�=���iґ/�d�2%��l����HZ�	ԟ���l�'QR�'��S�O����P+{T���Dޏ&�(y�+Oh�d�O�Į<%ۘKH�O����CL Xp����ĳ@b��A�'}��'l�I�������>1���<	Sš k�j�R�sF��O���Od˓ 5 Y3 ����'���5S$�9*g�	{�8�j���RR�,�I쟜0<�'�y7"��c{U׌B�?��8{��ͬ�?1.O�A ��Ʀ��O�B�O�0ʓm}\	Rb�%&�9������������I)R��������f�а�`�1:��	�H��?�vi���G{X���4�?9���?��'G������'��󂭛�D�|�;��0z02�/)��	�����?c�h�I�/���H0�,.�n�aCJͩcC���ڴ�?����?��#F4`_�����'�→&`7ʰK�	�#WZ� �MT%v�����X�	-�jc����˟���+��9Kd���U�h34n�@t���򟘓�������|:��?�/O��%�M�fv�K!�7Wl�9�K�O����w�1O��D�O���<���4/���a3e�y?*a�S��"�}�u�x��'zR�|�W���-G�L�z���ό:��mM�qO����O�ʓ�?I�FP!����G��fp��I�
�Y�S�N��?����?���'A�N��<H@�d� n۵�şU����#>���(�Z���	����'���U�1���҆�G�|�e�X���p�*L�@��s���?y��@�iN�\�O��I�+��Mu���S��4��k�'��V���I"=:��O��I�?�2H�%x�B���9�����(@���?CL�4�x�<��!�ͣ�*A*�q�@P�L�'T�	�2}2�'��	�?��'��P�j�s��e�f盗�!�a^���	4�ܳq�8�)�*~���8q>�(��/�H}���~���O ���Ox���<ͧ�?�&\�HCfQk�H �+}��2!���?��,�!Ys���<E���'�v��t*ק<v潒!�KU�0B��'���'[��_�C��i>M����'��	��$n��Bǫ͑8��h��2��&H�*�'?%�I��4ϓFi�����P3�
�
 *�.
���ϟ$�vK�jy��'9��'�1O�`��Ꚍ6�J%��V�`�h�[�|J,_+AW���?)������O9���C�1�D������Q����ʓ�?����?�B�'fH|9�Y�#V��D�O��hI��ԡ
Od��O&�d�O���?��j�)���˔[�=s�+H.D���L��?����?Y����'JB��+p��b���q�Da��&��OFrEɴ  �rY�П��	Ny"�'3B�tT>A�I9�Zt�ֈۃq�0l�̍;C# ��	ߟ|�?��DW�� ��Gd�D#Y~HHa���@~�9��j�B�'��	���Ʈ�_�Q�<��6ʰ5�u�	
^���Պ�{�nD�?��yhVݓ'd�S�eɌIG�A�V���G�,1�`�gy�'��\a"�'���'��OC�Ɍ\��KoӬ(+�I��1�ހ�'ErJA%�8���y����ęC����ӔR���/ۇ�?a���?���?a���*O��OR���D� ��1	3G��X�X��G�Ov���,O�1O>��\��K#n;B:��9v���ah ��	����Iܟȫ��[y�Oy2�'|�DM�4�����8bX<��:|�*����$/���O��dg��2�A�'{NI�����ȡ��O��d��v�^ʓ�?Y��?��y�$����4i��x�BnI!��M<|�'��'L�Iҟ�z���&'
��F)�$N�Y��-�	7�F)�'���'G����Op�	�@O>{B�t���J����TNA>9
HЛ����ҟ�'�r�0u�I�R��H�����>ti�1d���O���O��X�IS;L@hk26f�����x�̱3�	Yl,��'z��'l�Iɟ`�d+]K�$�''b}{�Ξy��#�/*j�
��'|����O�1�$�ڋ!��9��(��y�B�z_&��	�'�E©"��Sҟd�I�?i�vdI���#@�>�pEoD]���?�fȗK� ��<��O�t���ـg��8�A�'t�葔'�Ʉ����'�B�'p�T\��Z�KT��\i;��?	�����Ny��'��h�������O�a�P�)E�<�@D�X�6a��X4����?���?��'��4�F��z�!�UeJ+P�b$��	� q \�d^�yuXI������� ñ�'�
�R�����ep���L�����I	{�������'Dr9O�8P�;Hrt|�$�@�}�*m��	W���'� s����'!r3OLP2&��/�0�ȶl0;��'�'�k��I�L�	ǟ(�<i*�@R~y�A�Z�:8�F�dyrMR�u����Ol�$�O&��?�d�.A�$�+.E6^.С�KD&d,՚,Oj�D�OR�d0�	�TX�c?sR�(��K/��p�_�A0����3?����?�*Oz�d�[� �ӄ*�l̑6�P"M���ː{�����O���O,㟴���R�+;Ur~H�0G�p.�Y�J�?<5�i�<���?�.O���	�V�'�?�-�#
V�T�K^�JlM�dF�?�����'tBg`j�%aM��"3�W�E�d�����zMN-�Ǐ�O���<1�/�jp�-���D�Od���;xF�J��`ѐ4�'�{�(���05f*p;r�*�?�����>���M��Z�L��$�<���iڪ���?I+O��I�<S�Qs'�+�M� G�r��# G��|�@�3�P�c�qO1��D�r$<��*�O;h��E�q�'6B!�C�'u"�'@��O��i>�����	�	9���-E��م-�O�;�iV#"�1O>���.��i�
�e�=qr�	%.���I��T�'�9�S��ӟ��I�<����,��R"o��vHh	��ǥ/v4c���"�Z�ٟ(��Ο��g.�/i�� W��%'\`eQ����	�@R�iJ<����?�K>���=D/	&,��5�z}���H�?��.��͓�?����?���?a���?a�o6J�,ǖ3�r9i"M&x�M8Q�x��'�r�|��'�b��
�P��R�9�Pݩ��Ȱ,$QB��'�"�'0B�'�RY�4�
��M���H� n$��S�����ʏ�?I*O����<A��?��:�xy�&�. �pk֯M��ؚ������� +OB���O����<�%
E�]Z��۟h��1>`���<QB�3Ι֟���|y��'[B�'ר���'��I0g�d���)	�j�3��F��I����I�ɦm�z� �4�?����?���j{��*e��xJ��2�p���`��?y(O��$N��J��Si�? �rP��I���!鑮<Fx�2�'��'�4a���g�Z���O��d������O�I��.ߙo�bMH����zc����L�<��`�5�*O���|�'��g�%_X�0 #�^�^0����'�؋��i�:��Or�������O���O�t�P�S�W��Q�G��t�.C4n�O�x{��O<�O��(�)�OZ�RrnU*2Ƥ�v��(0�5K�*�馝�	ڟ���&iJE����t��ɟ��I���#Ҏ��dc6�Zv��x��ߟ $���_�Sȟ@�	̟�����:��̫@?_D(lk`�@؟���5c���4�?����?��
���<9�ONjP���ińCq$cLLy�F0�yb�'1�'X��'��S�p�<I��ހ|��Ir��<h���-�M��?����?9�\?m�'z���$h�Ċ�!P�(���bE3ry4��OR�d�O����O8�7>^����O���k�-@jT�C��S����$�O"��?	��?��G��<�u�	*r�ˡ#�s^N8�']�����O����1�'^,Hࠫ~"��rD`��q��%���#�L:?�����?�*O��D�O��D�U	���O`�DG�^�q�g��.����Dπ7`&���OD�Į<qC�[ ���ߟ����?y��B�&�2Y��L��4z��IFh	Hyr�'�B�'ߺ 8�Or˓����]�b�H1%\&G��}#�b�=�?�(O�53�WʦM��ǟ����?Q�O,�ʅ�l3��P���X)��0�O^���O�M��0OēONc>�N�:.�����? e�4r�b�O��3��Ц��Iڟ �	�?y�S��p���d�a$��3Y�8��f�7P��柤�f�ӟ�IPy�OO�O��!�KԘ�U��u�!'%o6��O����Ojxqv���d�O����O���[
�X`��+_�-�!�ƉFh�d�O�*xDX`H~R���?�bL8(qɌ�U�*�h*�2��L����?yD�^�Z��v�',B�'�RJ�~��'*�툁�Y��tx"���mH���?	�iW�<�(O���O��D�OP��)�ԑK�˓�rɔ���R&$����rK���}�	ϟ|��ğ8�����?i��f��)�٤SR��/?�tΓ��$�Oj���O����ON�4Ϧ1%C��Ƭ��!��Bv-Z�`�Iȟ��I���Yy��'��9�Oe:�ڱ�#~�F=�g�͗Y����D�'��'���'U�+^U�h۴�?��hh*hHB)bXt!���!sˊQ���?����?�(OR���>	S��O4��%#� ����`	4��qf��/,��OX�d�<y���:4�O 2�O����ƪ�= ���j4�R�7��8U�|"�'���)i��O��ؠ;GjiӴ`��x�Z(Y�F�+bT�������M�(��d��ȕ't���'�dv�)ȗ�Ǥ,��xx���?I��D�������4���'�y"f��#��C��,;Ьӈǈ�?��jD8i]�v�'b�'"���+���O���%)m\����C�'
�tI2B�O��q�3O6�O>��I#K <a��(S�f�44h�d�����ܴ�?���?Q`ړO��O���q��)u/��O����R	D��~$��c-�	E9Lb����ٟd�	�fy^@�I�x�P��%D�����	��Pz�ć���?�����숽�S����$ܵ,D�,r!B���˰�Ĩ<���?�����d�(I��=�f&��=���f�"�nu��C�	͟X��G�I͟\��� � A�!�Dl����B�J#MJ�Ж'l��'��O4dsAEퟞ�'�V�X�4`g��-n����qX����񟠖'�r�'���՜8�Bo��3��lr��:ib �ACi�rN��̟��	�<�'����h"�)�����`퉷y�PL(@�j�����O��O����O�h��H�O�m؄zE��@%�QУG�,����ퟨ�IEy2`ވ1IX������b�p����f�1е�*6��`'g5�$�O��$�7Br��d;�ԟ�a`���!h��#Ԫd�x�!D�'�	0����4��i�O(�ioyb,�7i&<A#&f�b�*E��2�?����?A�S��?�I>�}��b��o�l���%w�Z}z��Hϟ$��+W�MS��?�����5�x��'�H*�g̨uT���H�jv�A���',���T�'��'���
?�4�IQ)B?1���JZ�f8.�o�ʟ@��ܟب��?���|��OF$i��\�
�B��TD˥&�)���'.R�'D"䘌<�OF�'󄀘Hh��MO�a��q8��'D�Ȱ1�'&�]>���X�I~!�� 
S�>ԢL.Q�0�'��=�dՃ����O����Op˓d���8�^�XT�����AY#���Qj׍_҉'���'��'���'pj��iI�>F-r'�R�0�:�����'���'�Q�|!�����G$�1zB�7��Q�t�;��cy�'�|�'���G��~���8y^�����i��gK�3����O����O�ʓG�����tg�-)Mb{&@G� ���GA�@A��'�'@��'=��R�{2*U�)_~��C��j�\�����?����?���?�g���?����?���b��7L��B�;7T`d��C�9�䓷?��FZ%:�Q_�S�Ec:�|��@	��^�DUg�؟��'ܸ��*t�L���O\�D���'ln�*e������C��ĆB8��`V�|r�ձR.�O��)'?!�`G�\����7�tm�3c�ٟp�B���X��ǟ��	�?���՟h�Oi��Q�瓚b<�䊵�؆V�C��'^���7l�������$+� 0���hl���Ӏh�_����jcӎ�D�O�IN9�`$��S,��1$SB	QK��Xl���ꖿ���'���'צ��yb�'�"�'A6s"��@P&��5��@��Ee�'��JMYk�O��OВO&��2�;i�
���H�R�<٧c�<Q�,d̓�?q��?�,O��3�tt��)�J�I���Dg�lP�$����Ο���Vy��';rFN�%�$S4�H(D����چ|6��y��'\rV��I�[J��',pyp%lѧT���ǂ�u~���şh��⟘�?Q,Oz�z�炊�r8e��~�����
�cl��?q����O��cH�|��_I�MjG����P�RE�L����?��X��RU�!}�̿ �md��8qo1���3�?	����d�O����|Z���?q��(ʈ���ͫ}��i��G�� ����_���	*(����wE\���!(��>���)-OR�D���$�O���O��	�<��!���u�	�S�J�����ķ<Q�hVs���ӽ\S�LP���	�u�b�$.~����}'�d�O��$�O2�	�<�'�?�S�үE{��3JI?�h�����?1�i¯\^j�<E�d�'��\��S�5B<iʰ�  	��p�'���'�҄N�6�i>)�	˟��w
h�ZS��(�ޔ9�ݡ-B=�O^������O��9+0�uI�+��D8L�1(�giJ�D�OZ�桡<a��?a����'��`Q��3�XA�F1I%��KL>�`��N~R�'BRU� �i��>pv����Rl
DRK8@(F��'^��'���p�4�1�K�f��\�ǒ�0AȖf�OF	������ҟ��'9B!"3j�	�6j��F�_B@Pk�iܶZV��'@2�'��ODʓT�n��a�(Ռ�j�� 1?>r�-���D�O�D�<���t��,+)����
`�U󰌐�ª�*.������O��2��by��ʨ��9EY��9���"^��%'��ppj�$�OF��?�ph����O��d��� �4.�dԾ|� ʊ�\>�Y��2�I���� ��`7Vb��Ӱr�=�bLX�d�$�-lp�ʓ�?ɥ X7�?���?)���j-O��w+]6l( �⪌�����̼<�(OZlw�)�� �vE���&-�W\��h�Rn��Ge��f�ڸ�@��S���9�'�ufڴ=9Ta@`סdhP��0>�
�Ѷ�[48@��`��& ���D�<��Md~I�'���'���'�l4���̌Z��Ѧ�!v*"��Żi�b�d�O@�de�|�&?i��ğ�Γ��`��#2����^0�V�"'�<WX�{@.�=i�I C+�m�����'� �@��٫������hL�`��T���A `�/\�{S-Z�!t����Ui��=���i��[��`Q�Z�<{�P;�/_�	@�4�+f�����	ou���	�	s�S����Q��(���/1�h����?$�x4	�C-H�RKf5p0�p��o����n�B^8��P�c�*5쓮<��١S�U9�
�P�'�b�'��p�u�I��8��E$]�<�f% i.N��DΉ*j��cJ�`Kl��%DI q!<�blL��9��\��Hy�@T�H�D(���3��m�+:jLa��$t0��m�|�k�16wМ$��V�O0hGHBeOX/%�@�&��>b���"ٴ ��'�"�'}�ɷW�6��	R�c��1���S]JB�I*)bLT�3�G�U��,s3&\�)��j��	�?���gyb���`WƘ�f��9�>P�eLL�*ՊT�&g��'�R�'��	��'�29�,�Bc�]�0)ޘ Õ�h6��!��נn����m�!0��0e�C8?��?i���.s'��D�A,3��Pj�TwH�3kh ��"��-A� m8�&8�#�f)�	Ԧ=�P��9H�4�/(4�J%X���#�?�����O���'S�X{��>1��uQ4 ɧF�6ԇȓK�¥�SnP$PD�iAt
�M���|�V�'!�I��h|௟����~��-I"h�p@Do��d���cc��҉���'���'&V*���~��� H�P�<Yp�?-�c.J:�<��*�>�L ��.ғh�hH�#Y�p�VbVd��d&�pi_w����"4�pt�ʂ%�,��m�(O8}���'R�i
"���S7#�@�|A�Ȩ'D��>�O�Uc���U�*� D�R�,�Y���'�L�'�1{`c[ �@��EG8�L��'���+TB|�&��O��'�����?1ߴP@��m{Seb��YKu;��h��C\�0�FѰ�C�+`P�T��5���
�b���	�����L�7�i������V�+�ҕ*��X�I�č`���i��0p�	�~�XՁ��ʶpЎyiڴm>]��矘��'�ē�* GLA�^h(FX&�vЄȓY���Qh�D?�����~�X�Eye:��|�޴= �{��V b�H��G�����'��?����'4��'h{݅�IΦE�s�V�(�i��k�NA�CE��:���mÕ4�$a�U�@�.W��S+\ult���6��"I|U(!B�	�Z]a��*#K|�	1b٘-|����=*��,�R?��M�o��'����$�5e�.��&��~P(�X@o�OHU[��O(m���<!���� Vٲ��� �*Mb��QЯ�;i"l�'��'�ʟ�O��+a�@J���0��P�k[�MC��i��'����Od剌�*�#a� 2ѫ�jN�l�r�QЀ�m��čR����̟h�	�9�2��	�HͧD��]��-צi�*�i�O*H�}s�� ���Vi���4 �.Ь�M��x�'{�E.���ɓ_���໕��"�Svo�:(/|AxR-A�m����۴Z�0�FyBjS��?�ᤚ n^���V�O�MU�����mPT2��i��O�}E��KZ��E��\�;"��\%܆�C�V�y1AØqAb��Ũ�z!  �v���'���>(���#�4�?A�����T2&5��Mڊ��	�e�)>uJ5�f�S���؟Ђ�a�
y1�����W��=�F����֪r9��CF*W�b}�EW�
��l)��Y17�d1�뛫\�d�Iɟ8Y@�Bݬ
� �կ��3�R@ D鉡z���d�ĦQ�ݴ�?��j�G�	꼀�a����H���� �?E��'�2P����sP\�@�<>O�Ň���I�@�Nx��J���峄�\�(x�I�~\�) w+�埌�Ig�� @6z���'�$�nզ	�B��Xu��¦h��h@�]�u����ЊT��U㚅��|ʉ�ܴ�6�b��ݜ:�FA��W1d�na^��P�S13�x���N��ȟ���� gLV,R#O���n�p����M#Ԍ�ʟ���~J~���d�mN@�@��Ԋ9)�}27��!'{!��>�@���BY�m
nd�da�5<Q���d�ܦ�o�XN��Q݉�> (�@�� g`p���?@����Xa��?����?yа��$j�����ĜnȠ�璽Z�`�����MM&a�0��<zr�e�����S�u�p�|BFU37�l�b�#7��-�䟰A��r��.�v,j#NW�n.����"� �D� ��p�.��¨)�0�t��.GD���'@M����?�����'��ӓ;D�b�̏?'���JQ�ЪV'�C�'r�¸ �T�+��a��P>9�y���	9�M�����F���IC.[	@��q'�G��x%چ-	1E����O����O�� G�O��d>iåJD�l%ါI6 �P���SvE� g_� �gaʻ:��eF�+U��D�I`J��� $�%b3���Nיs|("oA5((��Cu�I�\g�����S����
��Zd\�B�[�)��6�6�	��H�2�8Ϫ��B�G��Q9�/C��y�J�3(0��H� c�Z�~�ӈ�D�< ���1����'5�_?��T!L�G�<M����
�nP���R%c���?��B��	�q��({���aK̀�����*
�Ѐm� 3���%�_�Zd{�F[�')�%�SM;�ހ��iR,ю�ʷ�\7��*ṕ�ֵvA� �H�Ӥ��p�'�	C���?��i�Y?���I�#���n`) DW5T��	ǟ���ԟ$�I'8�<�'���*���[�F�5->�œU��(AQҔ���g?�ÿi�ў�+���m�b3�_0h�h��sC�a7�8�O0���m�ş�I� �S� 	*D�	oZ+4�d#`�@-�̑�g��eS*���d�d�,2� ��	V�0$c3<r�`������%~j��@Z6;�\M��(�¦]��4����!S�=��!#+�x*p�����6��`��*0]c%�{����iN�j������'E�����'G�im5S2��f��
��2^**���&�O���(�O,በ#R<D�P%;��K1��H�`�I��HO�lZަ����ٿ!@Y��
)�n�I�)��?a�D� 0�󁛙�?Q���?���+��n�O�6͐��6اB�t��cw��d�	*Y�uzg͓�&����Ɋ!u�%s`KϺ����1+�5	(��r�͕�`*��
�Cj��*刘Vg��J󪏻)���3��'Y��i%�'s�6-���Y����]}��\�+r��Sң�=�� ����yRA�=g2i�򄄌+9��k7G�O
$Dz�͞�3�B[�|j!�ƿ{,�L�%�S!_��%T�UD\ �d�O����IΟ��	���D�I�dͧs+�,I�N�f��+�`U�]m6�#ϕ�O=�1�@*ָCd�E���r�L��h�s�.�C`e�;up��4"�%P���_3��" ��N�x��d��Ly��U�8�}��<i�� ab��w�<�3Ep����<!�������]��6	:�@�������L�!��J�`/��Zqo��71X������D	��~�U�@@����u��'��Z?5��ņ�$݁E�Q!*��� C3čX����?��B5�� �dՐ6�Q)2��j�֟<�Zn���p���Z��X���	.@����S0f{�ƶp+n\�'lX�\�F�8��D��l]����EzL��?a�i��6��O�!�K7H�j��p�,��]��i��'~�O?�H��PE�A��C����B�h/�|R�(}�B�z�m"e��]��+��V��~�X9�L:g�'}�_>H�O]������
�K E�H{�-��b��R��� h��u`Á-W��]P���:"k�]>9&?�d�/�A8� �]e|@��BF��?�ӥџj,>���J=yY�p��n�\�E�\cŴ��!E-N�LakRf�(���۴q 8���۟��+O��s���R�	Y�ع�S�u�����O�d�O����<)���O�Z�C�O�L`�em�6\��uK��d��5��4�H�h���!���* ��*}����VDyR���X��)� ���.ѣ2�bH)���9	����ƹi��DO.���P�&�;m8��9�(�4�H��ʚ�Rg����W���ݼ?� 	�Q�I*0!��jf"Jͅ���ը"�P:!�$YY��\y�	Ɨ$�n��g(��Jp!���h��|�w��f�D�3��I�;m!�N����)Ն�28<~,X�& =V!��J0�s�՛ ��Cvd��>D!�d�2O������B�@A�IJAT0�Py2i�x��lؒ#�u��i���yb�ā[�u�X������y��!$��1r�Z]���4�yR�V�+�>�ȡ���u���兗�yr$�2J(�q�d��hR���n�3�y�BJp�dƈ�5��%�V�<�y2�ؑ��|���C%?f>U�F�M��y2· U�]���95aR(�V���y���VR ��o�6���X��(�y��@�n���������y���K&|!�F4b= �w+��yr��gW��`)��-S�)h��\;�yrgѯM*�!�ǎ*�S�%���yr�c�\�+�Ȯ!|ճ'$�y�S�e�P�Y���
������A<�yB#��jQ傣�B�;��y�.����$b�	�s	b$Y�'�=�y�$W֕B�EC�]�3�+D�M�P%ݹ!-剄v�#|�'������ג"��|�3G�y�V���'��4�D�
b�����s@����سAL"�8��˛{O�( �'b⭩�'Ʀk�����&us>�������sƒN����P/�yih��B�RZL!Y'bє�ч:D�|���%|NL@�e�2�,cT�8?����$b4`��0l�RD�į	���Ob����A؅�D8�C�b�V�R�'��;u� ^��i�(J�Y��u:��ٹW���@�%�G�����H^�טO��'\ĩ���D�0�Ѵ���U-R�k	�^̽�w�ƿ�F5jE�9{]���DP!�|��QLU!rZ���W��CH��0`j��ICc��K�")�G�a�џ�Q��A08��M�H#��*��؛I�,,��͠���[�Vp�T���"��NN�J�z�7 L�]���<9AJMl֖�m[,B���s��)��p���-��lg��cO_;^�Z	�IH8�y�	PD�<�ё�݄|�ଊ����!�)��m��*Ϋ}3�lII~ڧ�����EhH��W�ެ�d.ؙ���lؔM2]���90�8�2�&�"Ѯ��bH�|fp�S*�eV�i�
�.�&�?i�` ��5�Ӗ}].9���a�'�3��|�Y��'bu�yaܔd�%@3iΜX�t���R���<aMۃ6��́�W._*��$̾u�^!�d�<[���#A	�8Xe��##O�؛%	9�Ĭ��fM<p�DBdO�Y�ļ3qiM�Yf��S���5|2@H���! �TQڇ/Ԉma�j���iW?�X"�GW���IeΌ5�fU�S
�wun���Q�֌9��W�>�H������	�΍��ii�h��;j6��G�2i���D $�-oAHB'�a���d�z���R&х`��Pi�U3s� �K��N��C��.=U�}S�l]+D�LE�_���Q�ן)ʰ�R�.բ~����^����H.�f�@Po��E�$�D��"�?��֌�r�/�8�MC4�ٓZ8��� �O�](w�@�9�Ճ�	|�h}�B�ڜN}$�3FݯZ	��7J&/���T��;a'��ŀ�~�`eFzbfO��4i�'>��Q�o�,g�0`�%x��x�C�4���Jf�� I��/O'?��mc`���n� 8@o�/"n��0������wm��b �
 �hD"��,7O��+k�N�̱{֬�8d���gI��p��d):d��]�Z;��C��K�ޝ;��Ʀ}'�R<t��	��R���Ҥ��J��v�N�p��Fy�Z,��,�C��@��f�N�x��Zǎ�C�x�f�3�@��K��*��L�Yd�#.D�H�l}���0@�|�&Y3�L���W��,+��<�bԺ&�_o�e&\�l�H�SO�hJ�����]n�1�6� >�lȂF߂��n�6{!�G#�LU8X���"j�v���(ڌ��% �ږ�V�J.��h0"MV2+1� c1K͉@��}�#aT+tj��fP@�؜�]%:\�'FL<a =	KB��E�s�T�wo��S���	�F4�a��T�tu"q�>d�8������Aq)�g�'��{��
�F0Т�@<X�P�h�9���Q'�(b ЛU)U O��\�s�
>}�e��f�?]�^-��N&>���;GZ�|��d��0
Jl��銦u��@�t�J[�'ը��u$D 6P@�	�'t��OӬ��d��*��F^+h��L�c-J�J�d`�A��Jc��f���8Ԧ��L|b%m�(y�� D�����hN<"ěEm��HԺl�F��F���4*P�i��]�~�&-Ȅe�cꙮͺP���Z-Np�px��M�2���:PL'����ħ�`�3��0
�ޕ�HS�"�z��1�S�5d���[�<Q���(�`>������'I&֘����r�(��ݽw�ź@��"V��xk2m  \��C�/�,��O�rv'[�m�
#E�N�N���#�>Z�b�&3T|���/��X���$�Ƙ(8H\����yf�<�IЃ1�I%Zef]`�L3@�t�,�_ґ���R�1� �a�@!^�O�����I�d�����ޞbL��N�+<ے������с��_���O<|��A�,��n�1�Y��/G@���J�f��\%��D�"�D�i��?��¥��5��I�=rd�t䑾N�<����+Ja��#�HH ͳOA2�0�r�P�)32A��dP��HOxј����9|����ᜃ}�zQ��Pss����<���T�!�s�oe�LHg@��E�R����ÑeTI�P4O�d��S���ƙ����2�M��q�`��AD,̈́7	�D�ޕ)�g��T�>� ���Y�qh��u�,�K	 ^�-Õ�A�΍	�'�!V�4��	?��y���_�fw�E�@,K�O�\C�I	>��%1�!з]�����]�Q���p�@S�5}�5�\#�Αx%ˉ�p,1���^������S���(W�r�t�AѰQ���qo=! �T��k7O���F�s�)9a%µ^��� ����Ԍp�O�<)U��KG�B�2�AA-L�#�(ٳ2%��p�:$�@���O����M>�@g�1.����6_��H�],ά�3�K=r�x	RC�G�!���J�t���#g/�!j���av���R��8�v���R����6		�g���$I�
>
�����'a�)RU�7
I"��`�=/k8Pr�#WXfp���S�	?
��FC%d�!Ze�C4���?N���&A�(B�⅙���6w�d����0B�%OL<n��$�'Trd���� ,d�6�A�n�tC�كI�J ��)�w��=��\�9���t"A�a�&�i׮pK�!�'r�gE0V8	���cqH/O^�@��Մ�Q0 �O�Uk�Ą�CQI����Q��ޭ?�F��e��r��D
�+M>ͬ���+�Yޔ]��$ ������'i�ɮ&��]��B�ީ���06���bڴJq^P�S���0�ZEa�柛YD�y۔:�#�m��y�-�@��-p�_�7��ubDƠ߰?	�+�,���C%怣p1�!:���?5-�ܿ�M{$NG�A*����#EBr��7
 D�d<CdB�;|6x 
�$ֺz�Ԥ�D,��vMP��
���'�9�I�J��0IV``B`���9|�����T'@]�K��#�L �sm��""a*ԅI�2z>R���"<�n�PҠӥEV�8��s�(ң�֋$<UJt��aP��K4'Z��ⵃ�V�C0��	"8�ܣ��'��=�����St皃{��˄��8G9��p�EJ�e�<�9� ���%Se�(9�(��B�'�\����O|��ck  `�&�a /�{Nt	I�V��.�S6�E�g�ǱA��6�i���#�jT~����Q�B,2�1:�X�����v ku�ܵNH�����޽O��	:��)Wc�E��D_�{�����	6D�Z��۵?���h�?( ��X�UCWeѴ>����H�9%��ζsZ}�#��:���Ѯ	3�XCg62��Qb&E5M�&�%�Nc���7A2�$eXH�T�[?�X�D�
�?YBF�n�9�m	/^��z��-��śvA�wՌȂu(��b����_<n�<iw�i�
uY$�A9^V�˷��&w��`���f:���c,��]�]��l�r,���GeZ�ɪ�O��y��2e|�i�%\-�:�S��7�b����Q,XL T/,�
yY�׫	B��ղi��Q� Eܣ*g��2���q��OZ��QN���v��C/!��0���T(��l��x5mZ3;F�����f���/'���#�)�:U��n�^l	��A�X`��\�V�u���sl����5�V�2`�2q�e�(�";��"6Ꮤ2�����5E�B i�c�.a�\yí�6w�y+�(��$6��Z�!�4��aHL�Xt�J�#��LT$X�e����O����+�+��}��BA2��DF�7��œuՓ>4U7L׳vQR(A�.ݾ]�@�3���v�l![g��1�����m;&u)G�W1s[\$Q�N(�t�6dʏ @�� &��u���)=$(N�����O�D�A���v�� $�ֺS.�a��C<誰�c#_kN�L�.�;&>�1�
+<2��֤�l� �;��=뢤�3��Br��M�rb��r����߻l�*\(�Od�Q聾u��}�0N0W@i��>�NB�s��ja���c����2�mRGkЩ��iV��L�%��		G�D�"�O� ~r�ժˑ�J��͔(Q�t)���,x�E�Ǆ<�P�j����v���ː'{O��;`T�R���gM>�|)�o3~�j���']�!�6�(F*��s@V���Ъ�%�m� �j��;|�a���[Y�!�fMS)B#đ�@���܊��ݒi=� ��l�(v۶qq�m�>r����m^�h�6��!)�Vݠ�a�B���BP�r̻Ф�s�(	!�(�[&�A�	>J��(�*ґ`�H��E��tɔ����>��D�T\��'Bm)���CN�q��'c��(��	8��X�s3��*!��4@L�X'X��я�"6�A/�V�ʰ�%���0�B#�C�^����7-��u�@�Âo�Ut�Dw�RH��.��<8pp���E�D�@w-��,��q�`h�E TL��/$:��R��'I�Q�ӄ�;Qrm�"+�a�	�	X���H$�J�"�$�����O	lA��Ҩ�,òl�PIɋ\������I��MK��ؗIk��,QA���d �`��H�K޵X����I,r��Vcʶ5�����G�C%|�x1��A���VÞ�lt,r�B��2�i $�m2�piz4�8�%)�$
n6���v�v� ���7��Sd�Y
L�P�>a���7�u�壍H� Ĩ���c"*Y3���7^1<'%R4Ŋ�r'���T� �1qP(Y3�L��p^\�e`�%:�ɞ.B�1SC(H#s�(�r�^#r���B$11��rn��/��)b� �)O�3�H�q�<��(_ t	�Ź�D^
1��\�#@�-�78,�q��4��D�`%�OЙ1��ɨe>���Q�ؠ2�H)e�Fs��O/7�1B�@�R�ıa$��*a6����c�#6�li�wx�l�	:cL:EvAT�x�5���'�&ȋ�A�Sc���� ��a �ʜ!s.����3\�q�o���i�	\xQ#%K�"�)��%y81�0��0Z�01?O��	U�.@I8,)fY�@dn��@��9���1��άFD" y����Dmz���/�RR1Z�*K/k�>MpË�Bg�(9�� q����FS�4�<MC��N�f�
'�	"B�@�� ���M��SV�J�˺�!a���|E����=cH�@K��᠉���V�N���d�����ڈ
�`�S��#Lv6�P3ċ8>U����/��;�:$�TG3�I��<���"M.��O3��$�ɩ	z����D\�6�ZE㞺N�������p��JG�t��i�aN�u�ܨ�@�$]��	a��U�
Q$<�>�zo�30r��RQ�(���yI��S�<$���)�"�%��`�厇�0��Tf�86�Hp��ȶ�?	уA�Hh�C�L���@�en5����::���6J���y1�W�MP� ۼf#�a�T�Oeb ` ��-3q[�I�ڐp��$ �-޳��dV���`bu��6PX�1��ߓH>t�� �ɥP��L�P%��@��%��#���'��@���|�n�1�.��v�F]i�Pd���Q��[���+l�i�K$)�t�	�4~��jR��9.�v���e��2�b�%�R����%��6y�b���VS!*��=Ya+�(�bիĭ�����͟�P1B�V�j�J�����U��]�7A�&\`����(:Z�b�j4�p��!k�J��c��-S��q��1��hy��d��a�!�Q�p��'�,	��f���DXՀM�@����@h(ĺ=��O�$n�H��`�� �Ys���
��%��%	�6DC�hRt �!^�`E�d�4cAB6�'ވ�C�l?z��K�e�{?(��-?�?�����PR u�'�C�,݂�U�}��<c�e�%y54(���?6I��F(���čk?:U0�Ĉ n� ��2�8Aޑ�P�I�#JL$ �W@&�C�  [�A�G��[䒍D<0:�a3@1H� ]<TD$�8T�@�.s�!��u��B�d{f�Lm�*h��N�ўl�B- ҄-A#�6	���oZ�L��A	�j�y�F��g4 y� �'���*�fi�q+^ܮ�
�R<D	�u�5oZ�c>6MiE@[%z�<����96�kq�E=� ݨC %�?YQ#N��J��H��>R
\���@�5�sA����$�ʕ�,�i��DjłeB@��!LK���Ԋ��\q�4��L�$rRڔ�Ov�ǉ7f�"���䖷\�5�1J��{�� iB��7Wl`mӵ+����)�獍�"L�X3e��6_����!}��4)�DϵRd�AHwvl��_�0!ؠ�+Zj��N�lՠd��	�f�1P�S3���� V���zTD'1(��r���.*�V(*�o�BN�L��4	
�∅�W�B$�Ϧ2/��Z��iij��k���m��_&O/�������X`V�B��Gvy����
*>n���f��`[��zB����/u�Ta8�M��v5VD�_2}��BV8q�>��;ړq�|h0uc]By�9�7��P�X��ɆR2ڥh4�� ~)��0e�s�lL`�#�
Gs��G"��Q�T�Qw��7�U���>��V��!��(��Zx����Ɇ7^�Y��E_�<8)b�K�FxX���bNp���B ���0� �5[��D�Y�<A��H�5^o�d��e��.�0{"��.at6��$W08��:Ç��H�C�d���|Q�ǣ�-O^�6mI~O�6�ô]��ݠ�+R>R8Q�o	Z"*l��^h�&��4k����(ٓ_�@I)7@F�8#�">�F��[%9C���(� ܰ�'Eo�&�mܤ/R�kd�M��4i�q
Oܲ}��!T:D��x���S'�����m�g�'�Pēbd0~aS��^�6Ъ�'�m���7�j����y �eY�Y��	���lY�ׂ�g�N�!��B�[���s�E� ;��dY6l�S^a��_�q��H���	i[ĤS�Xtk��0g�������&�M�qڞey���p��P��		iX¨K7���y��ƈRf(��l�9X��▪��x��F�S�� +R~R�����^%j��ؘU��"��g%O8Zv�y�ƪ
]��;�M��g�-:�>�'1��GjE�Cb��ªS�b��9
�wƪ�K�$G�R����)K�z�8��(�kg�B�`n�(I�~��Wb�����V
"8t�(.���tq��H0CM�Ѳ6��?|��^>qj��T�~9�$�¤!D�<�p�6D�����+;\����/��_�Ĕ؁L�O����%��-�(��U�L�6��Ҭ��j�lٕ#NHRv�JV�׋�y)Sn���+u$�!P�y6 �!?�6��#�Ҽ�B3 Z���ODE[0DB2�vg�!ږu8d� �O� 5-A:��l�C\BMpY�ʭ!a䠳C����?����͐��U)g��K��c�<�"�
,*�:vA�:\���"��Z�<��T/+۴�w�Ե0l\H3'AW�<��H�J8�%N /Hb,�E��V�<Y���)m�" ��NL�[t��aNY�<!�1ms�t[@�3�$ْ�(�V�<Y'�
���K|6�x�g�M�<�����Q��T6 �!��+Wa�<�gc��	vTq�c�@tq�C V�<��Re�aK�T�'���3k�P�<��e��u,�j�K]"�p��s��v�<�"@^pf���y��(���<��(O+D�H�Y����"�0��Lw�<q�`�>⸥z�LC"{P�i��n�<AWΙ5v��rOX�	�|4� ��i�<F
���>����9F��C�S�<� RuPŦW�v�̬u�޿m�^a��"O���  �IhXP:�T�8��H�"O^ͪ���2�h��K&�f�0�"OY��Iv�
�!�nt�Xz"O٨c�Z�yX��r�&T1"q0��4"O�䆯m����_<{S.��f)�"YDpĲ �+�O�|�g��F���A�ܼf� �"O���A�c4�8����:9�\�y�"O~:���C )����<gH� �v"OD)+�DODݠ�A��O�g��@(b"O2(鄁�*	�PI�lJQ�L��$"O�l���Oo�Y� �Tkb�h�"OT�Z��+}ZVɑ��F�]^��"O��gº�d�sަIe��"O�����'~���	��C.��W0�y�a	e��̴`" H�C/,�y���V�(��^�W����`m�"�yR.R�Ӕ��Ox�ܰ)"�y)��T�i��H�M���r֩���y�o�' )��1���9>�hy�%-A��yM >��Z��BD|]��Ĺ�y(O ��P�Ξ�3�~MQ�և�yR�\�<�8�#��G�OJL0�G��ybMΊ�ta�cǕ ~�R�[����y���e�X�HC6p���`�^��y�fI�uKԀ���%l����ǣ��ybH���ij�cՇxu���'cP��WQ�6<T�$�9x�����'0��ek�\_��zE� n��Eq�'o4�2A��)�vT 壏h2�LB�'��9�a�$>+Y7Hh,Z��'IZ��T��U<�
WF(!8�z�'?b=:��.�q�Ӻ"ư��'y�I�dl3 �RT�g�BT�)�'<j�KQ�n�!�`%0���'�4����;f �b(*^$
�'�T0��X�@+����(X	�'�z�۠� )�e���S�n��͡�'Dt�'���[s$�@�b+��	�'��K��M�`���`& �a%Z���'J��X�$D�8�J�(�Y���2H<!��A"03DT;aH9���rP3���b�����+B�%��� �
2l���8�߃}��!��`C�	<��`����|�]��j�y'd��jH�I�$�Px¦E*F�9���<+�B�X��Ƹ[*���On���D�17TYQ��LbG�٘c���@@��@T	j�#�%Z!�xR�5�����h�B�g�&g�ݱ���4�Y3�^ a�jv��=kO��tD�usa{2`�/8�(��^�@È�(r����ɝz��U�@=:o�B��Re��֝�:d����(�� ��BV��C�Ɂk���Ȇg��u[��R�g���O�,�6[���K�S���vN9�;$E&i�阎LC(�&�_�%�6����0zjĐ�AI�Ti�
��6��BR��$A�%(��F�%}�bɸ$,5���P�J�(�)�;e.��c�G6U�P��Ȇ o���R�?MPD �&E�V�@���n��D������g�� �ma�Ipgݱ]����D�(��,������q��L�l��Y�V �
�"Y��ц�H�!Y��jP}"D����b�%W��Y�� v�`A�"�h��ʓrh�Ӈ��@����'Xzv�Q(͂�a�đ/9ْ��T�#�
� T$	8B��C�/�Xxr��|r�CUnyrk�c���2��M���R7�2�GM�p>��*v�99#���<�P,�v��I0"�"g���7��	�#� *o`�ـ+�J�D�A����2f�Y�O��f��,(P��"ߞ$�0O�|鷨Q^h}9�B.�����ʙt��u#���*g�b�h��"H���c�>����+��L�Z�p�'&�I��Z�`R$Bo.��db@�,��V^\1`��բH�(rIZ;�`*e�rLʔ� �u7��ss���n�M�Z\!&a[�x��P8�'{mP��I[�ĥ��Ov���D
�^( ��S<F���q�cF(��q�
C�h� �#D4v�Le����� �`�E�	 -�L�ak�iA,V޴pI�Χ�S&L��P�K$N4p#���X�>��i�B*�q�8�?�	#%2ŪLO.K��p�T`V%#3D`��}9,���aB�����J�1*TQ��&/Gc�wZ`лs�X5P�l�V��y?��ν#D�^�С��[�	"^,ٺ.Ľh����ƅ'!��'QH�;"c�+��1E̛W����{Zw[(`� V�lj^�#䵸�R��^�m�0yHS�
��i��L>��g͊pf�U��j�!y�bP��/�֭
c�L�m,f��{*�PĢ d&.����b�^�%�G������%�~�+��E�R~����n�G�"I��а�V2Dx�l�ћx�iՍ$����c�C���'����$D�@?��Kfb��w]B����P|~�x6J�W����*\z��Qj߶_���s��L�-��!�W�%�l�!x>�'��O!��"tM�N_���4J�vmJ-@���Wt\����:#T1hӮ�"T���]�3�p1�B&��o
�T��̉d6%9'�k���>�N"���x��D|؂!��
�7��RL��~�h��#��
 ڬ�sr�,A��P�v�����)N�U*�`*c˄_ Dk�CZ�x�X	�9��4��h�Jej�� �U�7IX
Sn!�
�Ӽs`AҐ��U���]<?����@Px����P0G�$�C�,jA>t*W�@�_$�3'XQ�P	��C�R��� uȏa@�]�%FF:8F���%�:���a�*�?nT��=Q����fm�F�^a��u?!T��\�mY6�I3go��
�XF~�d��&N�Y�&�L��b����O���eG_D�pFd^5jД���'���B�7!��T�E�)A��������{�9u��Q��s���	ZT�<����<�)��IE��Y���H�y{� LfB�S�E��]^P���p��AϜ�`t6b��E���rj<4����$�D:�,pb�Z�k��8��ʌ^�'��MY�E]�9�E%�&��c�O�53U�9g:U����c���2��/A���Ň�]*�����Z�S�#�B��z/
�z1�XmZ 4㤝æJ���DcQ'�?k&$#?u%[�&f�a�fR�	5(X��.ݭQײ4jej:6�&d�T��%(h����$6�vd�"X�T�v��Fa�=�BaQUfWv؟�0�KQ}.�ZS��+|�Iy��-C9ԇ�ɜ.��C�w��H�J��*9�ϲ`Z�p�|KF�kʁ�i��h�B��z���P��Y�`�l���M?�-z5{�JZ �t�y�$S��L�'���Z
Y'�9�r#�N��a����z����J*��8�v+�C�I
^��c��(X0	�&jL�?�����1y�����)"ƥ���Xp�'!�E��芉����%�ZB�K$I��"~��=`�TB�c�[�$�����\�@C�I���8}���h�Mߜk���L;p! ��ͮ6]�̺r�G!P��=yqO��H�M�D��q&�9ztTx��'uD��u.�:�Ty�+�8P9Tܡ$j��_G�ej(jQ ��H�-*b�y�s�A6`ց��'	n�ӕ.��(�<5�CQ�B"0@L>�G	A��0A��i���T�K�YԐ�+"�!���᫒����*�/��q2�!\>>*�kT�'��QH3
?PX��Ֆe���ts�Q��P�U0Q8SiQlXPPK55_��[��SU�dw������#�� RA���dx�'1j�#	�Th�(���ЖKz��T�O�x`b��-�M�$��(,Mj��+��	�6R�`k�;�|%h�A�j��2��/X�b����Gb�Pɳd�#:?h�X�k�Q��;b�~<m��Dʒc�A41d�=�ɕ8[V��R.]�7��	blX��BX��?yE9>���]1$�np��(W�)��1�@�+0�O�0�D�^� 5f��[bD��'k�`��[dn����[�u��{�X=m1��0eʾ>��̓$@�h���'vT�I��Z�g?!�Z!�V�cR#��M��,;F	�9�dRvcDb�b��� נG�0�c2
B4a?V�aV+��E�,9B�ۼ�2��c�, ��q�*�r�`��P9��٠D�Ј��
7�6�EB-��bŜe�┺@����@�+�rIkV�Qdc^�Kt��uD�#�$��"M�DC0ꅘ�yZw��]3"d�8iuLԩU�rA�EA�9�� Fn�s�''V�ȁ'��A	�5FBM����2����oɸs6.��)Ն]��k�b�/Q>�I溛���6�f���'�.��!��sB��D�f������MjQkQC�	(Sy�l(�c@!c�jP`aG����sʔvu�4�7|,.59FÕ���y��C@���I�g<Lhj�V� ��V���O��=Ju�3?�ՎV.q����^�K� �� L�ex���O۪%b�Dy4�N�T�ӂN�?���N�Cˠ �Xw�f���	��D5����	dV�$Z�N�3���HEFD����_�Un��:��	9���2��H(!��Q�X�Z�(a��I�>w�����=�u�E�$�u�˕0'� ��+O8A�ݮb���:$MK�
Q�c$/G�O��)��OL�'�*E�����Xyb[��9{��J�i^;Xf�}�֥��� YX�MϨ0����'��d�'�(헧��Ҳ/�F�ݫ �����(�q��t!ɘ5y��O�u#��H�H� Ϯ	rHS�E^5v�X������p����4Ț5j۴t�Uv��4�H�e"�ɐ;��p����<�j��X�IC*�8�<m��iS�#Ap��Ĉ�ex�(�'�¤Y&$z��*��G�0xz<l�S�c�p�����=�u�'������H�!�@��䢛��������?X��U[F���hT�Ș��O`� ���V��
v�Y!y�|��"�>�| �ꌃ$��5�W�)hJ�ֽ��s�<O�'=�)�p�Og\Aju���T]�w��R�'��p��ċ<n%�I·f���ܣG�����ϱ&�@CS./+p�:�'��4ϓ��OQAAW& Ϻ�1C�% �
KP�޺lȊ���R�ɚ,H�ܒ@ʂ0^��|@D���@������/�<(�ӅP�ʬ�¦H'bct�e�d�^�Ɉ.d�Tb����$)�H�2�VUcW��q���ж�$?Ag�#Td&	���<U=�Q����)0�^ �n��[���Q�'j���Bc��?	�Ȟ��泟���CȺl�A�e͟Ob�l�wJ�O��Y�n
�u��ݻ���9'$�?��)�`Dۺ)�X�8c��9@�8�rGe�V#=޸���Q�l�ÇS�q��pq�@X�+�x�b�ٖ|�8�?���"%��}�A�X2#��С�nU�snX�"�$EiJ�rAj�F�zg��k����$iX3#b�	�h�>(�2LZ�K�����c0�Y�X|��!���$���&҆A1���Eg	F���|׌�`�&�Ҭ�ՇvL8�?���#x�1#*�2��[�?����A�x�8橖�95t9cnվIȨ@Z���'z(��K��u�F�����䡆�y�t8�O����=�Y���Nú=�e�Id��A��)�0�˳���B���	J�$`��,�"&�o�<�2�L
�����/fj���Fɒ�?! h����$� X��ށV�<�b�-̀f�Aj+ %������,��r'C��;��Q/+:����)e�yK �z����"��	_�0�P2��O��cN-o�
��#'��˴�!B�pW���'y�8'�rS���c��9�(���� S�LZ#3=XYz�o��?�9��D2-b��S�'��>z��3���C.L%�&��S�/�@��cc��x�h�5��th�5R�,r�P��s���{,�
nZ!!��ag��h�1��4��)`ޱ�W`*&����Qd��\��*��34�,rR�GC=��f�:��l��� #n�qdaС䶍��̤K7����D"�󤜆$wl���C�w�����D�?I����S�70��@!�U�{��H
�ϗ�))�4J1�Px.z���N<ݰ8��H�+��^/��'����'yp0u��`[�c��Y9�o-�v-�a�vE(1N>�e�12�	sBb��w��p�`ƐX�x0cSL�2�:0Γ i���2�
1\ŒB#�����'E�@'���Zc<���nS���yM�sH �H��0��b럼'X4!y��U)�5y�9+���;E���X�S20��g?�'٪'PY�mT�'�.|`
�1=���x�%^ZF$x6��Wx��zT��?	�Ḡ�I�x��/B�C혼ap#��>L\9�4��x�2����c��䝦y��)c�+���B� �&��d�(?��=�qS�dP6H��(��x�"X����J�k��m@��5?(��*_V��ل
�!+�P��#~�%�^��
޸;T�q��$*�D�%��u��nBT���=.'��WH��UO�L��D�|�+�E}��Qa[N�r�K�e�~1XS�O
>P��4�$'\O��aa̓�OoԼ[���GZ�� �:R^,9�pNܙQ4L�: ��	���ceU>�p��a>�λ>���!�T�c�8[6�3�@��{�J�IE�ك3����@���&�@�O���'� 	���P))�8yt���n"#%�H��[��4k�&$�&�JfOVUx�4i�._&�HbGF�t�Pꅅ�3n��(���a���v�[��8�9���@��Ɏ�$�'-��V+���`��Mqc����h����j�DR�1RRHi���<��/ϲ)�%���e���Fk��Fo�8�ȓ.�+c��rwh�K���F x��ȓA�R�q�h��}��b6#�:[�8Q��
iB�"�?X�J�b0�2	��h��h����וd8虐�0+5�ȓ<(��:eh�Ķc.D��ȓR����e���}q�$3*\=��RmC���+�VQS쓟:��T�ȓ�*0�j�Cm�1��Gpl|�ȓeY`�"OۧG�ݙΉ.
F��ȓZM��k�	R������E�:���h\��[��&q�H�g �l�ȓ]�2	ـ�Ӧe���d��H]~!�ȓxȔ�� H1s��8	U"Y��t�ȓXTޘ�v��B֊QF�PU����a�����
��-h��	k����]�pё�C�@֮����S���ȓB�u��q;��:UMݷ|��B�IJ���QB�$#q��nbF�B�<ciʔ�Ef��0<�t�vD��}�XB��.���4	^����afC�ɽ|]��O;j�x��T
�9�lB�	�Lx9�E�/8z<q�$�B�tF�[aE6HX���mN.WլC�I�zfrа�N�li*;�Ǌ&�C�)� ���Ȗ�o�����Y$���"O��+u��:+&�lj@�2w�#U"O�QR��r��Y^��-�6"O�0�'�`ll�6E�r����"O��BFY
3\ɱ�n�s�@�+"O6�PWFh��Sbk\ ?�VSs"O"\�K4��!-����'2��H��h�^�s���!`WLiJ
�'�vT���\�z�bϫ[�n` 	�'�,�r�˕�z>�\Jɞ�Z���q	�'v�}cVm+AP̹�t!D�)�K�H�<!W �Y�}������4��]�<��-�0<Gd\��iH+;�hc�c�<�բ�;18��(Z�Ųlit �^�<�4E��;�"��r�H9 =X�h��M]�<�F9�t��`�5+�v��'�X�<�R��	X.l0���4i1����oK�<Yd�40JԱc�0�ppB���`�<q���h"�,y���A�/"�B�ɴ>�`�#P���>����E�&��B�I/	�l��V~H�m�vG�)�NB�:I��UCϜ>�����B��3�&uXvm#st���[9BUTB�,^m�y����,t��I�ÃX+��C䉰A��=�,Z���mR7T87��C䉪���1.ʬv[�����"ТC��.?4t1r�ԕ
�T��g�C?~C�	m8(�6��PL�� �� �r�C䉫`�.�صc��w��)����L�C�ɯW��#1���"���_�:B�I2b�r<;�P�P��`����s�4B�I0D��\ҵ˒L��h�� ��YB�I\��D �P.��aڕ[n�B�	�]/���.-S�v��"�v�hB�&\#$��K^@Jݚ�c�(8B�	�%L�	Idc�����$R�hl>C�I:GB��˖�H�g���IѶ*J�C�	���!�0M�,=�z�!�[>��C���
��í���.�ڐC�͔C��u�(	���+?�4�I%�#R�C�	�����	BA �b�N�v�FB�IJ�(�1v�l�"9$ֱ��B�	�`�v��oc>��B��B�B�I��"53rD��h[~� D�ޟK��C��5���	2���+�DxxEқ�C��.h\`�F�*DH�"⎢i\C�	Q^L�"AcXHI�b�#=XC�I;D6�tXEnΙ1 ��k<߈C�I�3��[f���>�*P[A�N�c;�C䉦]����5�
9���V�Kz�vC�I+M��h25��1�p��c)HC��� u��.a�������LB䉧A7�=H�l8v����+�~�LB�I�?� rv�һcʒQs���nC�6jF&M���8o~|{ĉ]�ZC�	;�b���C$HĴ���2C�I&\ʝ��^jk<� %�_�f�BB�II��ؑF
��X/�Yӵ�P0��B��5=B��chNz�"�����sw�B�I$^ܭ@r��o�0a�q/�6b��B䉏d��iX�:h����$:tB䉬J��p��Mu�Ԁh3K�1C�B�A�@X"�R'f����Q�C�I�ul���*��a6b��V�ߧS��C�)� P����!c�� ����Z��hx�"O��#���~���giX�[M|�s�"OxT*2��e� 懏2g�F��"O�����]�)�&��c ��C��ѐ"Of	a$D�wI����3>Ytk�"Ob	��B՝3�nd`��8kN��ID"O���$�U�s�ɘ��H�g6p�ze"O0��t/ք��H1\s(��4"O8�������RCT;5�d���"O(��#U��$=�%I�D����"O,)�׎69��LQֵ0 �]�Q�!�$�t����Cx=����# !�$B8'E:�2�d^"TEXD�ǝW�!�"hi��:���4x�2t-M�H�!�dƨel���s�x�<1�A԰+�!�ĉ�1��#��8��Ayaj�.ad!�dI�jS�}p0� #1���C�K1Jc!�D30)u�����˸0�LJ�'s�ђ���v8����A?z�
�'C.�@�&�=[�v��ӯ�8� �+�'����C4W�,�T�+.��)r�'җ�}�HQI��Uz�(����Q�<�Q'����
F�n �a���J�<aQL
W�d�AƧ
T� &#G�<A���L�`Kf@�7�"�;��A�<����eq�5�a���g� ,AC/VW�<��ˣB8 �w߃E�"�X�aGV�<Y�&PufAx�i�K��K� ^N�<Q�(8U�g��{�̙s�&I�<p�Nr�XyS�[�I���.�F�<� �-{��0HW@Y���"DA�<�fg!d����.^1���c�/�~�<y�.�"C��ം�/j�[�IP_�<�3��V.��C�.bR���SfUs�<����sk|���% �flv4A�,TT�<a�_�B�n�z�P�B�����
g`�����i{~��c��}�Z��ȓv[�����X
T8z��*�m��d�ȓ4�8mr��մsWG�J� ̇�w-��6΍&?2��J6��K�>���4Q��,�:����)��^���ȓ&����KI ����G�S}Lq��Z�pCw	K/Pc���/4�L��9B��$%�`�ݲBA�CbR!���?��d��je���>2� 塣�	��!�dI�-K�eA��b�d[n1E�!��-������)�-�
�!�䒃/"�-Hu@�0EN
���:R�!�D�B���Jb���#h8�en,1d!�$��H|�YPlPC����'X!���//j���?y�t��f�/P!��e�R���T�]�rE��Pn!�$ҝdba�(YE�e�B#m!�Ğk��#ķK>�����*j!��|qL5��Y�l�#�	i!��R0{�K��;N�0�8�"���!��Cx��X3��5���� ��!�Y�fĕ��&E@��H1!�Q�% "�i���My�� �H�L!�D�-@�K�%�>w����Bi�!�$�ZFH���.���ܻ���j!�$]'mlh�kwe�"w�b��F��|�!�d��s��`��8�rq��W�T�!�$I�g\4�R탋lp�%��ǜD�!�� ��2"Q��5r�l�,+�� c"O�L�U�Ϙ�&da��]�ld!�"Oh�e��bz 鎌
\n�p�"O���e�Ӧ,t��#x��h�F"O�p����=z�uр���Y4"O���4o��[B*��I��b�"OPA�G�<U?���.��	�2q��"O	��eaVlM#wA�H�፹>+!�$[�j�Y�aF�u*XDK!��Vsô0���,"J�0�aM�0!�d�2���D�E�a"��7�SuH!�	8z��h􋘌(-z�@��ϱ$�!�䅁'=n`2p�^%L+KجSÄ`��H?L��%�K�Bx؅`�0y��=m2����]:�S�ҩ�����Z��AYڀ"Qb��aZ�@|ćȓ[�����J�8�"Sv��;����ȓ�B�k�4Q�Vh%�řA�&Є�Uƀ�x��
<*I$����� lJu��]��qCB�$ʹ� ��cP���ȓgLư��b\!Td�`��[<	ʄ��d`t+�
Ï�RHB�JV�\��Q�ȓ2��@xd�"G�XM0���:
ټ �ȓc,�ecŋ����/�/y�"`�ȓ"F�1�I~8 TV�+d��݆���y�K�l��s� إ]�B0��CXe���h�Cf����!�ȓ#�0�RcX�Hzn\3d,߈g_��ȓ*d�A8�%�:Kl$�"7�O,��ȓ�T��f��6U|탢�5}�u��?"X�@S�$q��х�`Mƙ�ȓM�"���յqjʤ�a�B�X�H9�ȓvf��!�%U 4A�bRY��@��B��ੑ%ڻ2r\Ő� �#n��z\�'�E�H�J`x��]

x��mC:�`�#��P/MZ�p<��C@|�0��O�"�@��qNF�OI���x�<��	�M�*uS���!35z��ȓ<a[�B[�*��ׇH�Qp�ȅȓ2��5�1C%�f��?��T�ȓ^�RHz�-@�3"��J�CWg�q��@UJLh2Dp#����А!��,�ȓ���J�+����u.��#rh��7YK�t�gH݈:�b�R�M>D��zTf��r��4��z,�V�'D�p���?�<p��	:��]Btk(D��NX(.:��z�h#�eCP�<��X� $2��`<�`CT��R�<��׺\.&�Hp�M:m��j$@O�<��℀I!ޝc��	!P��'�K�<�A�\�go�e�b��#G����K�<i�ԔLf�Pj�le"}��"AC�<Y����c2��jW����$�|�<a�ڣ���p �&�x
B��w�<F�>�~-����!@A�c%A{�<�Z��4XD�:N��k2�\8G�C�2}�$��u�W�.oF!�4ZC�;-U,1��aCL�蒅���lC�	*����Nߎ))�s͈�BFPC�I��B)����7r�|�a�OlXB�I?s���tm�5㪀��5{�xB䉪��к0ض	Ǧ���"\�SK�C�	(��8�HY�j��&	D[�C�"T����S/5FH�����B�)� �T�pi�}q�|���<`ZL��"O�u�5C�A,�|�ȥi:f�32"O�SEь]Sڌɔĕ�</pă!"O���4dV�I�ͩF$I'mt�y�"O��Xql��n�u�V�F�#�Hp"O�oA�+�4�(7���d�{�"O���P��~]j�h	�:�J��"OJEk��0%R8p���!,���K�"OVU���SF9�۠,�6�a4"Od����/T�	��!P�X~=�"O����A
"��#"ӵ	�`�C"O�Hc�i#�\Y��B7 ⸽��"O$M:��[�9:�q�%������"O �&��f��@�%�
wveJg"O<��f@ް&M���D�e]ڨ��"Oj���掷r�X:���zN�͛�"O dz
ߗ5ꑈ�.��M^��#"O� 9el�e��xG@�1]���"O���KЖ_�L
�`�	}@L-�"OV��VOWw��2e 	u��=At"ODD�lA(*`6A1���-L�i"O��C C���n���9t�t��"O�ͪ��H��BiҶ쎽��)�f"ON��	J���PH��
%e���""Opİ���2�� kr
�:Ȇ5��"O�)E�1X��!����E�"O�5�@�Úsl^x�ݻ_��%"O��R!��,*;���0@�u{6"O��ҦcE����+DLB�<*��Hp"O^1�0�3D�|0���2Kb�"Oj,��J]|�=�Ɋ`�r�k"O���b���M?��(K!V��r�'��}����/e���-jm~r�'�P]�Fl��[������]Z �S�'��q�W�UTx"�¤���]�'J|18����.��9�G�;��x��'�j��2��78��*��f����'��LS/��,�^��ƫ�YZ2��
�'y�UrҀM�!���֧ԎV׎m��'7��8��H�*, (Ae�T�S�����'��@� aB�J��%�΂ �h�Q�'�>��A�g�R@!d�G3NwLx�'��1��dO`�{���.�vP��'�(LRڢ8�F�*$��%Ӱ @
�'�l���D$S�~��^�5@�q	�'H������j��s��0�XI��'pN�3V�Q�P5j�,._�Ց�'�8ҁ�	�2��Ei3*\�{�����'O2q�₈�ra���B��s�����'���I`nD3Fh���mdF0T��']�ٛ�C�w����f�kRA2	�'�X5Z���^��P� �$[��Y��'X�U! �Dy����d M"��
�'u4�4��������O�.�3
�'�ik���uA0�1Ŋ˅;6�|�	�'�rI�vA�E���ӏζG�4I�	�'�R���G�0	��� �m��?%�p�	�',BHdg�
c���Y���=б{	�'������M�\C���a⌮.����	�'C���d�(	"P�p��x�
�'tr��S��9t��<�`��H�X�'	
,�զ��F����щ�@�a
�'����'�U���!�@�S�}���$��h�T����wtp�{&�E�p��}�4"O� h�`�V%�0����U LRv"O�a{�쓂g!#�.p =Z�"O$�x1�i"�M�R��_P<�eOR~��';:��:N�ҝ˅�'`�h�'���)'�BV�(��[�Xpr�'�Z�C
�&Q��c%�ֽv�ֵ
�'`�`pZ'?�xx{$��@i~�)�'QJYB䈚��T0�&��$@bb�9�'���`1�Ѭ1B4�%� >7Ih`�'�PG��|ՏV�0}`���'�B�s�A��D�G��"0����'�E�3Q{��;7��7%����'�t���FD�p����Fa���(�ϓ�O��Bb�D�:<~�W̞� ����"O̽�p.̋o依3����Y��"ON�sb�N=0�D,�eݸV\!R"OδsvOA(��$���A`���A"OUx�#;J����
�A���e"O�YRe!I�j��,��$Y �0�"O��i�Z�\ r�[c`�M>xAE"O�h�䮍{ƒP��F�'V�6�'�ў"~rw N�J����e�ژ�d ;C�^=�y��w6��a�Ѻj��xBe�yB�B�n �\#2��I���Z+�y2o\h�&u���=^~<�#�*��y.�	�v5ʓ�ɋMW*������y��Ԟ0�D8�T��
E�LD3�U2�yb��~Y,Y��Y%���@�E���'�a{b��n}Ti�p�^�}�V�Kw��;�y"��+x�țw
N>vi�Y&IS��y�E���EJD��7s�R�E��yB*Sř"��b�L�$e	+�y��E5&\�A �Hp,�"^��y����6q�9aB��4]�!�L3�y��ٍD�X�j�W�2Rm�����'��zr�:�"��ӝ(+����mK��y�AXM�<Y!�.$f���F���y�KW�kz�]ht΍�,9�4d���d3�S�O���"a��}�ґ�B9Z�f�q�'�M��=��I0��N�d]�']Q	4�f���Iv�@�z��Ř�'ZX�7b�}��aou�2�'�b���'猜����u3i��'�����iF X�����R%82��x�'��yʣ��=CK�"��=0�l=@�'�v�9bEPp��I�0/��U
�'*�m��؊z�fl�5iθ!*<���{2�'g�!�-��W)4�'�Jc��̠�'V8h��ٕ_��XC /�_�
IK�'��T"
�:��{�᛿U�l��'#$�e�ܽ^�d�@7G��K����'��t����;iX�HQ���X\h	�'t%��
�%,A�a�
A�R���8	�'j�H�'Dɮm@̍���ŰB����'����!��`D��{���P^Fur�'�.����T*��'�"2���'��Q�0�ZWt�S���>%*b�c�'B:�I��"�]�$�]��8�	�'dHv�
�]�j!HWO�$yj�}"�)�)K3��!K�l�]��1�t�G�D!��U'wA��-�݂AE\�z�!򤘌GZtyN�y @��4%�!� !��5+��
a`��7ɛ5Z�!���/	� �gh3q�����*d�!�� Z�+�-�	:��)�.7?�xW"O��K�F�tR\@Zr�и4:�C1"Opq�bB\+�,e��/�*H�9"ON̳�"
�f۔l��.B	e���c�"O��*�!�'Z��9{��
g����"O2��-�:%Q~�J��31���D"O8T�%��8N��ъ֛NTj��s"O��+�=R2��	@�2%X]��"OT0�B˃[ �r�ώ'E~���'j���f��?�~�ҶG�}~\`��>D�`�&��7��\�U#Q��0#�+>D��S��"R�H����Ζh|��!�<D���h�*�tp&@Ε�~�r��'D�(C�i�F�L|���̦0�dc3D��ȴ�աf�l��!��n��-�� %D�4x3+E�&I.�I�������z��$D���T�G�/��Eɗm�++��rcM0D��A�3WvqH�j_�iu�ݩ�+D�Q1�9V����I�7$k2�*D���w����S���^B����&D�l9s�Ȯ=�m�Pi#dZ!��J&D�8٢�U�X'��!�iWJ=����#D�TB�lI�4oX���VR���A!D��3���'X��E�c$֑D*N��N9D�49��i�Z]2�/<P9�!Q�7?!�6ì$�􉞭-n��*��U3Y�J��ȓO�lA�/ :���`Y��D��s��� U�!�Ν�vF�/NtZ�ȓzz9��B�#`�c��� �r<�ȓp=�x!�䍽������N��=�>��4l���<��h$A�C�I�*J�K��q_ΰ���DJ�C䉰s����нh-�0��'�$��C�I��L�[���L�i���� /x�#<��3�<)�6@B[,N���᛫y�$�ȓE�ʵ�@�A"x{�AP��-��Ī�j1��I��/�q��C�zv6��1�)D���uG�s�L���NΒz���Pũ%D��z���.G�L��@9�@)��1D����d��'�0�2��M\@}J�C"D���2�lp�[r�Ðy}ԉI#,D��X$�\�@��(��D��U�p�)D��:僔&��Pq�V�H��x#$�2D�HxF�ǿu�$Ȕ�T�@]�b��0D��ڗ#� 3��p�Aǣz r�r��*D��8$��-](H�R�F	�k��'D��[Eǋ;�|�B@¡/��ܲ�#D���R�C;vd�]������Ȇ� D��S"��
C`�"���ܪ�@>D��S��<L�ܩ�re̬���b�#*D�����֏9���D�
f����3D�(�9-\�y�
����1�2D�l;F�d��$J6`�0��HY�A=D���O�hŸY��O�cy��Z>D�饊1��0��>Qr�@a�9D�$��A߂]}r��q&!�6�H��6D����c�6i�l��2F"c>J1Fo5D��3�L8 �����ܙ�4�ڐb5D��#�(�5�m1�	�)C"�C�?D��J4��~��Dp��x��)��*D����X��̀!�M�_d��c�e3D��s��*/(L� d	�?�ő'N?D�< ���&��5
��A�
=D�l#���e�z=ⱀG�y�l�F"9D�� xd����c�VXe��=Y�N"O�M�$U��v������H��`(�"OjH�G��.-@���B�#PĒ���"O^XIA��M�B�P���X�@"O�5�n�r���rp��F��%{G"O�4ѵ��Hj(��=%�ܑ�"O�ѳq̑�8m虢��K�d�L,p&"O�SР�X�~�QE�:W�\��"O&�y��B�F���� f���"O<�A��J�l ���*O��Q�"OlU`��(Y��a�S�%H6$dC�"O"��P�&|j���KA({%�
�"O���H

^x��JB<s#�Q�"ONyQ����t���°Z��ȅ"O����FI�PC�1�)�	i8�"O"H�V&҃}�$șB�3o�� �"O*�X��N�Y�D1&���%�d�;"Oޑ8�]�E�����i�H�ɩr"O8D���E�3� ��+�e�xё�"O̵0�M��J�JU!�n�ơ��"O4M��߆Y��ݨ�� &a�Ms�"O�(���rLԘ0P�7�d%��"O�)�ȋjO�yR0/V���%"O��1��iv��E3B��8�6"Or��P�Y�ky�d���^&!�:c�"OR�׆��Cr��(tMR-i��8�"O(�#�B* :a	D�:j0*M�'"O.�a����V"�04��O9� �"O�͊�S	�-�sO�+?ώ�BU"O\A���)t��S�`Q-QkJ��"On��&DV��a�@5	��X`�"Ob-�p�T�!4���S�t����"O�8I�K�%
Z�`�Ѯ=<v`}҂"OvER��̝.����A��nj�a@g"O�H!����Y5�TZ���""OB8C�l���ZM�E�M��8"Oʜ�%#�-:���]D5��"O!DA�-{�Tڷk*]B�"O�1"iFa�����B����"O��/'@YBh�C睖+9 ��"O~�r$Ē0u������+n�1�"O��M��?�8U0�]4^�v8�"O�z�5#6*y�q�7:SS"O(��OY����o��]la+4"O�1�/ǵP�x�+` K�#�,��"O��V�J�c� ��.�m:,}�'"O��Y��5X�|�:G1@`��G"O���cmՠ`|�I�c�%?��c�"O���C��t-ܠ ���$}=�E��"O`��S�ԍ8��M:��hB4I�g"OT�I�O�r�8epᒰn�\�Q"OF웳� 
����f�6J$�P�"O��S4�`wzl TE�(�Ip�"O���&��5�F1H�"ϰs�M��'�\y�g�0D,C����oj<P��'�]��`R5fvF�j�-V	m��L{
�'Bp؋���H��ā�v\,�	�'��H�N@C^X����>C�m�	�'����NY�#3A�m��9���	�'�����CZ�6j������A�"O�xK�jń^����!� NW-��"O(���
�hޚ�+C��p9��0"O�p���]�3#
��tf,64�9��"ORUS��N 7��
�ԫZp��"O� 
��"��)�@8K���lu"OI�Va�	f ��BF@�)-�$u�"O<	p/�&Kn�)��#c*���"O�A�u�u��{�c�a��ہ"OrՊ�!�^ռa��!�^�� "O�U����=&��fA�6m��K"O2��#N!z ���to�"^�s�"OV����2�`����)&Oz-��"O�m � U5Y�eЧ$���i!e"O��*�NM%jN�z���#�R�sP"O�]s7�O�*3��ȒG0We4�V"O*L���ϰ2t��ڣ��$YL"��"O�	Y��:��i����`:}P�"O&,*��.���CSo�#_.�"O�L���O�u�zYY��]MƬ�#"OLD+�!ɷ3b�d����}$�m��"O��2��ɯJ-"�[��3���"Oȸ�Ŭ\�<�,�cj��0�H"O���c��,�[�畿	r�AU"O�Y�4XTZ(9 mG;uk�ظ�"O�k"�
���	��.�{v$�su"O��@�.ff����5NI
I!�"O<�Ǉ\���ȸp�ۏ$/h�""O���'�;N|�cD�^�0#N�"O���EIΔY`����Nd��A�"O��8�ܑi� 8��g�$��"O8PF&�X8�TH�s�L��#"O4y���Q#3x�,c�R D�,���"O~�C76*�F��Wȅ\s���C"O�P�L�ݩ���!
��"Ol��2ɟ�q �8�N�LhD�"Oٸ�(��pѨiv���r�\��T"O�H�o_�L1a�� �v��"O�-˲e��R�t�Z l�'C���"OLj$�øe��)
G��kg�Tg"O�q��g��$���ꋝ@����"O��qU#�A���(ԉ2�T��"O,����*_|���Lm�t�@�"O��!E.�\j2���"9��8Ӣ"Ox��A��� �7
�88( "Ob�Pc�%]�b�Q��,Y�h(ӄ"O��s�韖�h<�G��
� 6"Ob,� מ<�ր��������c"O`�sF#�Vl(����	��l[�"Ot��g�J�z�{ �@ ���"Oj���H"\Q# +��~�R��e"O.�i��
.6"��fj�A�@"O`|�3���TΤɰ%��B����b"O2�ч�
(�0��hR�����"O Q���C&.غ'�x8H�"OX;�@��rV�rE��'��]��"OD��u6nMt8��f�)e4��r"O�|J�G-rx�$&ğ-��"O�s�'�EK����<M�B��"Oĸ���'��\�6�O�y�� 0"O
��h�6߀4[��G/zx��ن"O<��f��ȍs�kMFct�X"O�1A��;}����r�X�6z�`�"O\	P�㪚	?��{�"O�)��휹K�65��g�B����"O�Tc˻kv�E�_�_=%�u"O~��`�P�{9d�s����t���"O`���195:c�@�b��9�"O��f���j(���/�V���"O� �ܺ%M\=Z�d90E,
IL*��"OT��� :�Z�@w+Ѯ=�2��F"O|�J�dUDF�3dV1�b"Oz��P�J!vZvX�4�	h�R�"OPx`5�O;9�r��� �,K�n-�"O����.鸨Su� �4���"Ot}0wn�SͤL�a��!-��x�"Ot��a�=@��1�U(�೥"OX���-�0>&��
�VF*L�z@"O���m
.pRZ�Y$/ή�@��"O��t�҉-in,(g P�
r���"O���Α�;��|����:A{v�s6"O�T��4*�$�*g�B����"O�U�g�YI����+�k���"OPt����,�Ȃ̈́&VT��;G"O��pǄ�"c������\`�<0'"O<X�p�� ^�����k�Q�Vm��"O����[9A�X	�,��T*0"Ox`�1�ƈ�`�A!R�9�a �"O����ўW������i�hx"O��Q&��,k��RORWbLu��"O���m��Y���X���3��e�"O���f�Th��A��A� !�r��"O�PB��/v(.x��/��!�U�u"O�p#�G�*�a�ΐ5r���	r"O�I(�,�z��8�V-9
�;�"Ox���1p�p�s,#�(@"O�+�k��!��� vhI�"O༘���Fu�ϝ�\��"Olq˶��'v�f5������G"O��3 @���m��;�H�"O��K懏7$�y����(p"O�Q&fҬW��U��e�Y�b"O�Yk�D #s� �Q��Wv%9�"OXH�%�Ǉl��	BU�:�, �"O��'���*��rjH<�`��F"O�]��h���Lq��	U�d5"O��r2&@�ࡻ���?Y�����"O2a���'D�*h�<h\�c�"O�5)�nՇj�$���	��:�� "O�(�)Y~Q�nЃ��-{�"O\<���+[��𸃦/��x��"O⬳A�P/@�| �t��
�"� @"OR[�ٸ�����aωGp8l��"O@���I�'�Jy[r˝&Q}��"O:tk�F���,4�P��Na�q�"O�$hVh�=D@+N��d�hᰓ�}�<�h_!K����VM�"�Uh��\N�<I%�J�o"���#�8S�Ճ��AI�<9 %[4�Y��K49���	��n�<�uG�!gL8QC�[����iH�h�<�P N�x�Y`#˾r��Y��#�c�<1��2!�L�aTa�62.h�h`"UF�<ɰ/Q�<�)e ^�W���׈�B�<I ��4XJZ��̥�d�F�@�<�.�f����T�_�q�X�	}�<I���`�qx�hB�D� �&/�y�<y4�
W,�%3�ˉ�h��йw�/D���#&ʇt�,țDl�jӮx�%b.D�$s�K�Pɢ�Q��A�n���Z�+D��y����P�)�7p����7�+D��z�m��0x����/_��<|P'K)D�\1M'Q�@�qvBB5\>vT{0�,D�THgJ
�A��� ǚ*�����%D�� *��EƳ<'�m�U�ݏMvx�""O��sDFɐI���@i��N�����"O�Ez2.��=�^lY�f�6��h��"OT����=6��)���:�A�e"O<Ԁ����vOU
U�f��D˂�!/!�DܳZH��u����
����r�!����Hf�
�� ��O¾z�!��:n�:{W�^�Z�0<g.�B5!�$�#_1���TcJ�7
<��Fd�5!��L���	�C��!�P[���m"!�ď�}��p�m���$���̍?�!��!2Q`U�m�;�lHVƏ�l9!����}C2T� �]�S������^�Y"!��55��`Z��L�[g�)T�!�M��`����ݙ2�Ե�G͝ !�7c���X��ʅ� W�M!򄊮G�^M{�d7���bs� ��!�Ċ>.��0��@+t}������>Y!�䚥E�<c'�2v>��E�!�D]��J@��$E9~tP<���
'�!�$�,O���c�m�:V�a�墝�c�!�$9>�pbA�.D�lr�@��fp!�״
�I� ��Ԡ��JB�le!�DZ@4(1�Ul�h�2l�櫔(6�!�d�,¶�@�kə�R����2 �!�d��:Z��ºt�Hm�#�+78!���40�Iځ�þb�tx��7!���;��(��C�3H�3��x"!�dW�Oq*$�p��=��֬P;V�!�d�N���ʥL�M0D4�'^�W�!�DC�2U�<j&*�:z���^[@!��R���2�P�>���FR�-�!�$�_�����)� c�y2�ƍ
	�!�Ć7ɜ���/�'B������P�!�:[If�	F+EZUp�$���I<!��H�d�q�TC���ǩL�5��B�I)oL�u�7e�-/
r�*#�L�_�C�I�3�� qfB��ZdKS$F�ԒC�I1M�8ӑ	� X��c�+0s*C䉬=hda��CU)jm ����E�\B�	8|�B�1�bF	"���%➥1 �C䉝������ѷAF�X埰`�DB��hT����:e`l����|C�Ii%~�y@�
:j� TQ�&��cB�� $�� 6�Q82�*`ç$��:D�C�ɒ��P+w �E��!KU�X��C�	�1�����M4K��	�!�U	��C�I)����C��Udh�8��Q3�C�	�'����!��Eό�3$��5r4B�+"}XRD6:6Tuc�̪?q B�I�7_4�lג lՉ���2.U
B��-WP�`C��S�6[�NL�l|�C�Ɇ0�$%[��֔-vt�#���%y�C�ɉ�����A��N4��Y.�C�I26kHu�Q�W�lH�RL��۾B�ɊQ��0����q���nY/rrC�ɾ(
ͣ�oŁG7���&�	3�,C����(�
 �]���@%�W�P�RB��&'4h�cU��'yhղ���	Z,B�	�7����a�PL+h)����B�2�6P�/E;>�:!�1˔�C�"�+cȥZ�T���L��ar�C�ɑ,s~�CW+��SVm�8:D�B��'7U"牘�t���!�]�ob�B�)� �Zv���3��Q�ӦD�^�`�"O����Zs������D�R�LZ�"O䙲�� :��1�Y�$����"O�	����-v���դ֎`݌���"Oa[�L��hR�t���JD��d#�"O~���ƒJ�X�i�ٝC��< p"O���rE�e<�c�E��h���`"O̈PŐx~р"�ن"�^8�Q"O|hx�Ϙ��%� ���A�"O�M���6Aap�b�݄<��9�"O\ �)3V�+V+O�1�����"O0��#!L"�X�hԧRg��
�"O~LZ�HH?4�Hb��V:2v�Ͳ"O�ȳ�n��W�&Ū�싱rb�e�G"O:�V�ʖ!>9P��CO�8Ac"O:Q��.ң_Vzq�7�6?IԕA"O��3#m�u�����̇�4)x1"O���3�مQm"�����G�	٤"O�!ⓉHb&�d �g�Q8�d"Or<b@̳��08�� =x϶)�"Oba���&J���&�M,a���4"O�P!�"&�d�񩞠��U`2"On�H7��7$  0Z`���<sB"O�IR���o�։�p(�7J�-�"O�ik7��)2����x愝z�"O��r��";t�v#s�Ҙ��"O��i�	;�TQR���vy���2"O�=�S�ݕPΐ���u"���"O,}cZhH�Vi�2�0L�b ��0�!��7WMN�ۧ�ާ!2�r�!75�!�Č�$[ A���åh�������Pg!��:� ��8L{����g!�D�8��HǤ�1E~Ј
�A�$[<!��W��("W� wfX�� V�-8!�D�nC@Y��E	T`�It.�k!�ԅNr�"��%`Eb!���0�!�#Ov��hf$8�+b�%�!��+X���!�% �Y���F�!�$�/ʄ�a�f�@�ã@�.�!�|PU�%��+�a�aE�k�!�d�,'*Ra���OV�{Q@��!�d�~7@�HՕ
��G�2o!�D�0�xK�K���8Qp![X!��*���yG-���J��� S�QW!��-J�!�շEs��ׯ�qF!�DY:Yt^D��W������.� "!��5CU> [D�R�ܑb���(�!��Z=x���s��-_̀��R&�	?�!�$C�u{���+�&�,Ar�㔛\�!�$}�Is���L���ߔT!���Tv�� DT�~�B�ˑ�AlH!�D�v�4<�A���ys�+C�!�$L6j��S��:��$��,�!�ď�c����?ֺ����Xi!�d�y�*��%�C([V<�!�K�!m!�$0��%U䋒V^��%��(m!��  l�T��1X�\kvf?Y!�ґYqAbtE$1�� ���!��2w=���P�Y[��R�2�!�䝦8�4 �NE�bC��G,V?!�ͯ��Ͱ�"��/��j�ݥ)!����-��e�w�"�	���_!��P����HsryQ�ؕl
!�څV�
�	�f5QgN���BX�~�!�� ���&�D�i:���Ϟ>���"O<$yHC�f02f��?8J�(�"OȥJB�P�Hy<�!3ș����3"O��[B8��|u@G->r��"OX� ���*�@��\�1r�"O�y�
$��"�Y<
AC�"O���yB���:'�z���"O�AB��;'B���[=tX ��"O� ��Sa"aض�� g�b�ʡ"O���6i��%`չ֥��*i�$�"O
q�bԩ[P�]˲�K��fe�S"O2��V�AP�)��`��
�"O�93������;6�:�Q"OFd@�C\)1�A�b���zަ��E"O
 �Ǩ_>���K$E¦�j�"O�*aX=��$�QIʮl����"OD%R7��p54P!O߲Q�.tH�"OZ��w�����%vt��2���y�"*�W	�?{Bl�3 @��y���[�X�(���oER]C�P�y� J#=�(����Ӫ!|1J�e��y�-8o�݀^�[�(K�uE(���'�鳅�, �J�I�j^ p3�'�|� u�- �a����\��9H
�'�0��J\�udll0EV�Rz��' (Ag��<<*5p�#
M�X��'^0%1�
i쮥`�HB	���`�'��-r$BH�Dp ����&۾��'_�c&��3$X%���íQ����'=BY���ZKntPg��D�\T��'�l<ۡO\�|Ibii�p�� �
�'�D	��ă��(չ4�B�\��
�'�t��Ɓ�,D#h�[dNǥPPH
�'en�Q�����XI 5zL�Er	�'�:@�oJ�񂭰�G�w͜��'X���@L<8L���.kFMJ�'Z΁�A��?1p�s�)E�`�F�	�'�n�ã ���	�e\Y�\<��'�L�pp���Z�
y�W���$�6@��'&�� 2D6Z3�h����,e�
�'?�%q��![�h�c)\��`�'t�"�LA�2��2sl�
6��
�'���ȓ�{!s$Z�.��B$H��y"Ǚ�S�:�0ը�<.�\�3Ԇ��y��0 ���E  �t9�����yBo�����P#����Ǫϛ�y�V�Z��9����8���kF��yR���j@���!��9V�<�yS?^s'�²/���6aߗ�y"ɗ;V���W$U"@�M{��5�yR��ڄ��c	�z\
�mE#�y2�ۏm�Р�=	FuJV���y�FVE��X�#�_-H�)Vf 3�yG��I���Љ�<U:谅L���y�N[������GH'��ܩ� �4�y��X�*㺉���E�w������y�ʏ��*��i�~ǀA�����y�k��K��t�w�`�Rw����yrBW�kI$��#��%�~���(��yb�L3~�Z��0���#p���y��@�'cf�:�W�r����(҆�y�D�i�@��B<�B�E�%�y��^���Qi�Wq�l;`Խ�y�"��$ːPE�V-�8���֕�y
� ~ a�DV�({d)���GBBĘ�"O 9k#��mb��s���<2D� "O�a��f��$�������T$a"O(!)��{���5i׌C���"O���Fɺ[�}��iZ\	te#�"O0M�&CJ�L����XЎ}Q"O,U`$1Z̋�H��o��%��"O����Z��\�'iK�h��@�"O�B��	�@V�iQ�M@7	���"O
����be��ƻW�� ""O5��\����͑�o�KA"O0��U,dzZ�� 5-��C"OV�rE��	�ԴB�+��w��s"O���&j�4�����O�,� MC�"O<�U�@�e3�5ї��B�~� �"Oй����&m�X� �δt��D0�"O
��L	�(���bu�\�[��MJ�"O�}Y���yG����Ś�;���""O�'��-_����Q�� "O��R�.J7^1��s�, Y���4"ON䑤G�q���k�,@YV�id"OT���hV�aR6�wˆS/đX�"O��4�O�0X$����6w�,�""OVD#�k�+��"hњB$��"O\�z GY�����R	n��"O\qJ勘�ex(���ȅXc����"O�PZ�f JKf���i	�<^|Y�G"O,	��J/b�����H[�]O�Y0"O�XHt!&4�Ƒ���X�0�"O�<�듊3$�HXD� 8r%��K�"O>��t�ɓ9���9Da��[��A"Oldc�Cސf=��r`H�|)� "O�a{��5O'vP[�H�:�<�Ȇ"OBe
P�@�uw�dG�k�Լ"O��`F�ӌ�(�)ѓF�l���"O։i�gԒK�R�ӰNݠ0��Ms�"O`}Y�ʚ�WШ��P+b�2�w"O�%�
�ul�˕ȁ<v@,tp5"O�����|0�����++��Q"OH���Κ�Qv=�7�P9���U"ONUr$e�)f����Э�R"O�8{tʖ����w�
*H_*�"O��ǯ�(rI�b��-f8ԥ��"Od⅌�;Ĵ0{W��V֝� "O�̀*4}�Υ
D�̘t?��c@"O�)1k�pi8Y��g�L�Z�{"O\���L��bh�&�֦:��)�R"O�-�cA챸��$z9��u"O����z�j��5�X?�z8�"O�Qyg�&J�+w*�|�ּ	v"O>X�2��"��HɐiW=��XҢ"O�m��A�$qD��i�ե&�hu�T"O����L�fp�@�F	�Љ D"O�y�Wɐ�I�a$˹Os��F"O�Y0b)Hh��E#N=}o�a�f"O��� ' 03����L�[@��"O��r��×[��	�g Wl�6X��"OZ�x�J*|n�3�)Ʀmz"O� �<8���)�R���3K�u�<I���H�t��M���$(��H�<�R�J?^���e����E�<9V�L�c6�=����J_$8"�B�<�Akފe���M\x�,m� �@�<ї�լ$�JA�&���GbQ{�<� "If��o#��;�k�ko�2�"OF#�^�Rhn���ϖN[|U�"O�B�@X�Bg���jO$RK��`T"OD� �#<�r}����9~7�\"O���P��g�P��F;'Z}��"O�z3�_��xa"aG�8�|��"O�ȴ��{���f<W��Д"O.����)���+��M��)"Ony��*�/8?��
p�>hZ�"O���Lچ �|Tc�cZ(9>�Zs"O�����¢c�t���(�w�4�"O�D��� 5qÆ&mv��p"O�)��i]�X<a��B%̪�_�<ٷ
�{P������p�����y�<A1Cо-���Q�S���G�M�<��@Uy̸��nL"a0,3��K�<I0�ޗCp(�d��B��b&��H�<�֡@6&;ps��:�]V�G�<12L@3|�Y����5����@�M�<a�EC;i`]����&�ŉ�Co�<I��D�7nu3��ޖ7~�o�<��[�|X�(����0�꠻��O�<�6�U�hQ�E�j���t�T��J�<�V�Q�l��D���P�b�#4�^�<�pΖ��@*>r��X��\�<qP�V�R>T Q@ڿF�eɂMU�<�v�Ρw`$UУ�W�2s�R�O�<Y�	�<<м��R�έ���K�<!��[,v����R�?�4�1a�a�<ѡ Tؔq�+ށb��!`��F�<��@�'~@��F�n�R$�Œ#]!�d@>ǎE0.֦S܌�HC�D>!�P#&�c��\ 5Ϧ��$'�V7!�=4"-Q@�'0�Y w�Ծ7�!��n:�S��b������&�!��5�B|2r��m�r5T��I�!�F�	���F�e��������!�R�U�<���G�]bDQ �5Ny!�D�)`1`��*6�|Q"j�h!�$�>�8s���F���%��`{!��5��L!�J��N�X��ZS[!�D�wt���4I7vB�i�g�Z7J!��N��7� 5Q��c�f��&S!��C8>��h"d��M�H�8gEI�z4!�$.v(��"t�ȗi�|��gd@!3!��)��qk�J#�dYBdj�&~&!��&��-����n�6A�6ÃW�!��?;���� (��))�kR�*<!�ܼ�l���e�!��\�T��,�!�dѲf0,#�S�w�b	���v�!� gk��bd@�+�(��m�Q!��	)B�D�M�]��jm؜N�!��Q�6�4Չ��[%+���Ǧ�:�!�Y�0�
�i���B*��KZ:4�!����� �M0����� -Ki!��ʢ&�V�a�I�.B��DW .�!򤄂O�fͻ�cM�.: H���!�d�2y��qH�7<l ���)�!�$�_��8���L���A��$ �!��z�:��g@Kw���v�"O`M9�L�P�dPs-׉-�,��"O�$��eD2��Y�aS4"�l1U"O( ��=�>�� �ɶ	��ZV"O��1�J�j�x�Q��Q��K"O� �Qkd�R�(K^���Ի�"Ol����6/�I��*M�m�ny�0"Oj�"r��G�1��F�-��4�"O�D2��[;�=kG��;�����"Od����x��Hr��Z=v��2�"O �2gK�m�T���Ëz{��"O|���%��k�`�۳��-.R�'l�%�3��>��U+	�a
�'n������$�ۓ�E�z�D�j�'}=tE��W�xp0�&zhlAx�'�B-{��C��rh���s!d���'�y�!FN<� e[+ˡz�~l��'���q�\z�ey$���k:��9�'�HP�7�� ��=��DUwZ���'�� ˆ`B�C7�Ar���p^����'$PA�s��	����F��s�8��'��}R�,O�`���>x$��H�'0�5�0�,[�$���i��	�'��q��F�
F��iӊS�a,5y�'@�8�!ϕ1_=�$
�\7$<r�'H�	�,N����)��)t ��'�E$�	��V-s
�K|�a��'(�D&�R/v�,x�u,@tI�W@�<�a*]P��@u��r%I�[P�<�"h��I((�k�B������J�<�bޤc~H��"V:>����~�<Y���#
�Q�Ԁ+��M�y�<	�#ׅy�V����TZ�4zb��N�<�G�ғm�Z�i�ƀ�u5�S�t�<�p�R 	_�|�r�,8� �O�l�<��%�'z+|i� ӫPж�k%�j�<ai�����H���P/������O�<��̳0}P�g
���t�P�J�<I�g��9(Z�:F��/|�v�)�f��<��$V&� �_ O%����aBw�<��M�=^��%�����q�fYi�<1�'�+( ��c�Ȏmt$P�Go�<�E�H$%�К� ��+�j0�c�i�<���ۑ/������'�O�<Ie�X�P[Bl
p��0����r�M�<c��Ibd��M �s&�-��	�Q�<�aC��m#<-!��/�"�k��JP�<�Dc�*r��,��D�]4yc%�b�<���b�`Ȩǉ�qs��2gD�<yB+Y�<���r�'E�aĂ�Z��D�<��ӑo��ɨ���:q��s�
W�<"l=R��Z�c�p���0U�<�q*�'�dd�č�7d����Rd�k�<A��T��ej��-��r�.Bn�<q��u�8تG��)GC�љe�@h�<� %W>b`캷c�'3�j��嬅`�<�e�ب��Lb��)���*�f�<)Ƨڶ	���Ձ\�X�*�K�o
{�<��ć�=j����Y��h+WB�t�<aw"_%lb�h�͑2c��lu��H�<CT�]nD�P��w+<�����E�<Y0�]#6�4U��ĥ�%,�i�B�ɴ|j�9�w�޲�$��ܤ!�B��O���vM�+bx!��lC�	�H6J홦�\�`�F�����o��B�	"F���@��5aܽR⪓N&�B�Iq�N�H�i���E��=�nC��1-�h���؛~�ћ���:�B�ɂHl�A��0{p��P�C0{~xB�)� �)��.]%yR���J�5|��S"OPy�q�G2t� L��C��\4�cr"O�c���f�нل鉾8Jp���"O�iȣ!L�g���+�AZ�7�dQQ�"Ol9�%O�^������ʜ�jy��"O�����_%	�� P�++�L"O�I4�K'QH��31'�
^ H�!"O^y㔂ƜT-�h�d��� c��*�"OX��6 �!����,Uh^�iHR"O
�F� �>���k-aDT�:�"O*$h3AJ I&�a)��
$0)6��"OJ0KCGС	Wh�sJ &"�p��"O�@���ə�]"Cf��,&�4�s"O�a��,�/7]Txse�5r�R�"O�`s@@ʶ&�
�:T�S X�<9�"ORQ:eo��d�ȭ@D���^���P"O���d�_����E��r{��h "O`�Z� 0��@0CԡWvB�#�"O��2E��$�l��cB>w��j�"Ov��f�{`�`�(i��("O����C<GU|�A��;G�X�"O�]B�AV� �5؄��qGPD"O�*�nȮG`�k�M�UV���g"O�1��M<=�,��sg��7���o"O��
w�͛u8�������d� "O�����	�KL��[���5�R�3V"O�8I@���gv�tb�$ǓI��
�'�(�Ӧi6\����n�.���2
�'ھ����n�\e��ō!�J��	�'�~�I�J�K���*��jX^T��'e¸(�Ɠ-tVu �C׹j���C�'�(@�#X%��`��
$]�"պ�'G�J�kɷ>�p��@�P{n-	�'w���LS�/a���ƍ(�L���'ɠ�����.�`wHQ?&"�\1�'X,��?�r-�v�A��܄A�'��ʗC�[z)�d`H��� �'�J]X�/�
�6P7��P�;
�'G��s��j1H��f,�;=K�'uD��2ρ�~Q����O�}�ܼ+�'[�tYS�#Q¡8�.G �p)�'_X��](7�l�ǀ2Ko���'KL�#Ek�>Z�V�M�D����'�F5KQ�^���A���=����'�$�ģğ(:�IeEP=24h���' �	S�ƐkR��a�CD�8zX���'5�h�C4d����p@Ш`�A��'�
��4�[�T���P���qBP��'$Q�7��!b5�h�f�f��{�'���r��+!�����ŵ� �:	�'���u��90챛u���,��+�'Z�kr���pv�9��i�'�x���'����I+�����I�%֤�
�'���	��)�L�a(&�y���!Ԉ��p��D�@kϰ�y�˚f�V5I@jH8�F}9� ��y�DF�,�P4�+�hD҆�,�y��?��<���2)x6�g��"�yBm�#�,C�bJ�"��)��n��y�Ѿ׀�A��X4.�	I'oތ�y�̍[7�D�'��%(�j�6����y҉_��FYe�R$U�k���y2�ͳ(�ԡ��X���6G��y�
�4�,���gȽK��+&�Q��y
� ��g�k��	4h٪�Z��""O��`�B�1Btpm@�ĩ�n�3�"O,q`�L�m��i#��D�KqT�H�"O�mK�h z��ݪsd��;O���T"O`�@M�.�T%�%�A>Z"O�����9��8��G���5"O���І�(:�<�qdR�n	�� *O���Ё��]?"��$�(o��l�'�ʐb��W '��-�/ӵ6R��h�'>R���#�0��H��?)���'�.��!N+i���h˞�����'������$t7�`6"_�~�\K�'���gȪm�0,�@[�*8�	��'����O��Y�*gNDx�'C�e��kƤ"M�P��	�(���'v�$r7�hx�!.${�L�q�'p���a�CZ�-H1+�{[���
�'����e]�,�D�q��x�h	
�'4�P�G)�5/���)];�{�'��H��;v<:�Ҕ��Oh���'������ťpׄT�S�]^ �;�'��(��FC�f4�
�N��F,U��'\��C��$:y�R��#���'����F.]7c
PR��_6t�8�)�'�.�V$�c��-0�� |��T�	�'��� �b��Ń�G�+n�����'�J�Ј�
A�@]s�"�})<K�'x.�h���+����ĳp�2p��'#���d"�0�a��5.(�0�'�4��%�< �:yx#�.\�A�'znP#���$�=�R�@� ofJ�'ٺ����N2�f�Z�$��%����']i1��1\�@&�Bʂ�h�'̚�zV��"�a#[�'�p�i�'<\�QgΈ�Z1��yt#��"��H�'Zn ���m&��t�6r��3�'4����>Uø���ܧj�j� �'�x S�aƞ\uPPL�8d��;�'?��X㨜"AL���w	�����'0����#zPF�qG��8/�J4�	�'���3`,����f�"+��P	�'r��yV�D�&�R����E$�	�'�P%�K���H���x
	�'蝋�ƞ�l��`��~��-��'��$�G�ٛl���@7 	�E���P�'
(���� �bf���?\~U��'��X�dJ�\rY��
�M�T@�'5Ȭ#�
ҿ+f=��EA�G���z�'l�d�u �&K�8��Ac��O��L�'����zbH����N�^9�{�'��]Ғ�T.9�H]*�'>Y'�1��'��19����r��t�/U�b,��'�x��1��/t���ԯ��KO) �'<��w��c瀘�rFG�'���'�-���X�q},��DN>�<�
�'A�@h�CL��i2��}�T��'njA ��KBH��T'@AD�;�'$.=K#j��3��uZFF�6�JT��'�zq:uᄆ{�HcUb ]I��B�'t�x�򇚛FV��g��i��P�'�]��ꐿl������8_�b���'l8����;0�I:Gc�%R7Bp��'�(� G����y&�U<[`,��'2���
lx��Qg�]�P������ �4�備�m�6cނc�ؤ!1"O�<�� w�$�נB�P5���""O��#�EYb�������BttBC"O�S�&��H�&nD����Y�"O�Le��&� �>��g"O����G�O�TP�ԌU8~z�53�"O���b�����!����"�|�<�偄�6z�|�C�7���Q7�x�<	��$�CK��"�(����z�<9#؏S��(тF�(P�҄�v�<��`�#�y���Y$�h# ��G�<��MǴE9����߸���n^@�<���byyh4��o������{�<)� F($���K�q��e���Q�<�&�<(�VM"6�V@Tes��ZP�<�M�!��Zc#��{v��f^H�<�DD!�qY��n�:yɓ*�B�<�T��(���OѕOɌ��F,�F�<��^�,�zT;F*R�{�`��  J�<�0A��%��C�7D^ �/�Z�<a`ȑ^ �
��[0�t�qF�z�<�N�+XȨS����~�i���u�<Q��Gf"rA�5��Y�$Fq�<�YL�U�P	x�69:�j�0)��܆ȓn��q$�#yDB6JR�=}�-�ȓx;��+�A4dA�9�RC>@�P�ȓP�3w�![��D�P,K!(5�ȓ�hM#�Y�
s¼@T��<ec ���DdB�
6�LR�6 dı��@0jH#�!�#ζ�Ca �nLB��ȓp@�S`C�C�~1C�ǽ>赆ȓP�j�T�4l�Vd�S<-*<)�ȓ"�2¡��s�i��7O��)�ȓ�l�D�K�+J<!��F�R ��ȓQ�Aav��a>)�h@,c<h���To>�v���)�PI��d�����&t���&�7:��A! �0�|���<�^�IML�WE�A�Gꖐu;���\q�E(eR����0}X<��i{��J�F@:2!�Ȅ1+�9��t��bP`���,����+/ꭄȓ:3ĐqŶe�B�3S�N>{�$�ȓH5���GS,wW2�3��N�$g�X��}���R��p0���R�R���ȓS���儀4WL-{1�׶@<�)�ȓV�ұA��И�ED�-$Ef��ȓ5v�@��ts�<c����;$<���9,��㦊�[���瞃О���5z��F�-^0�pFV�Pe�y��"��9QV�()hP�n��6E��'����7`gP�'��E>b�	�'!�H"����~�`���, REh�'��Įҗ:�db� N>��D�'� ����ݶ���2�j�"���'�(��.�L:P�rC(�s�t��'m>����
�X���"�TH��'�8�� �|�h9�"^T�ȼ�
�'\ޡjPC2*�Z�`�$L|XP�	�'�ֵ���ܮ\j�h�u./AZ`�S
�'��[�A�[�V���օ/zx�
�'Y��ڒ(L$5�����#����	�'Z���U�����7��j7v���'��|�1�v��rg&�#+�l�b�'`�x8p&�2__X�
��H�-�T���� ��{���v���"a�F�/��'"O�`h�i	�C~�y�&��`�s"O���cG}�LӴ�ޅh�bu"OD�q@�H����e�>0����"O"yhc�͓�ĢW����=)�"O<�1��]#_�P�;U�/L,T�c"Ob�p�]�a�PRcK+G"��"O�!c�V�DD�81�BIm`�a6"O�8{3JU?TQ�:%%�y�5"O��KV�SEl �g��!N����"OP��$��!��Y���ȁ�6u�"O�����U=0��8 q��)rZ��T"O��ia�����u낟@n�-j�"O��Q���iK��?9z8k�"OrQ{�OJkņIj�ە<)>���"O�0h�*p~����I�wvT�"O���`��w>�a��Ɇ�jȅ�`"O� �P,T,Ȣ���)F]vdS$"O��i�ԇ]�ހ��1@�d�a�"O�� �j}�`j[���d"Of����+0���c��(ht<l�"O����C��ݺd��%�d��"O��`��wwSd��A��� �"O�Ȣ��U(xw�����*cpYQ�"Oz5��'�I;h��� $_&,=hB"O�@�Ra;�9�&�܅"$�Z�"O��a��#tpj"�Q�,���"O"h�QF�>*
؂���g��00P"O�����46g>��D�&�J	{"Oܰ��Q'C�:e����)m4� ��"O^D�&�Q��k����c����"O��C4
�7?�:PP��\<}���R�"Ox�R���5��8��eԋB�(��w"Ofx��`�!K<�T��`�<Ȉ�"O�a�g!�>B�I�wJ��LR�!+"ODyRQ,X#5�գ�i��kG"O��r�֤�����m�`"O�D�PML�te@c�F��|�X�"O6pC'�� 	����A�Y�X�h�"O=�'�'ǨŹ�i��a�� ��"OL�:e���p��*�)��N�k"O8����U�8ՂAXl��"O����M�HW�Q1�!>�]3�"Oh|��+�5;�4c�&F}�� �"O�ȓf�RP�Z�F;nP��"O�4Wˑ4%��[#F׫�~��d"O�x�Qę92d�MzR�������"O��j�ͳX���̋qּ]� "OF�xQAY"�XC�	+�����"OZ<17L�D`�h##t�2�	�'z�!�m�z�zB�$�Y����'O�@��aƕ�D�yuK��K3���'�^��ѧ#è�{�KɊ4�ȕj
�'�&1RW��+
İ3⩘&0NK
�'��qA0��0�p���=%I&-	�'�"��	�H��x���*uԈ1p�'�$]���������㩃�l�)�
�'��y;��ؿn!ٳ��B!�%�y�b�2N��qb檈=����dH���y�n����Y��V]����b];�yrBD�N&�Ax���T�^��"�W�yR�
� D �� ���Q#.A�y"��0=�ҽ��6��0AR&���y�H�=��x�G�{�j�>�y
� (z�#D8!N6L*f��zT���"O"Akcʁ�,�e3f�lf�83"O6�B�>r�q�ißxRXm�t"O�����#0a�ȫ��>$,T�"O TB��5hr`e�bH�E��|ʢ"Op�30!ΐ"xr�ss�)~~VXY�"O8�Q���r�6X���M=/�q�"O����'#PP��ia�@�(���"O �-��~��U�bm%#���"O͚��Իla6���	8@��!"O�yS�O3^L�����բX��d"O�mI�N9&��u��]�.
>�8�'�Q��8�)D�lP�EX���oȤ��#D�4�� -b�JU��aÍ�.��g=D�LӠ�N�C���`�e��?D�PM� ���-�8Wh��;D�8�uB|a�+U0q� !�0�="��C�	�=h�B��8 5R.�~r�C剦l��@�RX�a+�
@����D��C�NwL�0��&_����ZE�<�ѣ�@G��Ī@ cȨ��A�V~2特E�O>�"�
��j�~���V�Q=8}��g*D�`�$	"a�4��P��/���o��M[�.�ؐ*g	�U�yҕB��B��X��I�'E�qy��Q�0	P=)a��<Q,��'��%�Bۨ5)J�e��I��LQ��hO�O�"�h���E� �M�0a.��	�'ӎ!�h�=R�,��'�$� �
6-4(�Q?�dRp[���ɞ�;�ĸJ0d�#YnE �'Čဤ�K��ac$�"B�
�
�[���<���N�l�80#A�q��J��� B��|�2O ��G`�cW+F0tl��@	˙p�B�'n�D�u�����d�13�||�����0�M����F��~������W�b��A
3敼�yr-яot��c�E��D��pN	#��'��z��Ʉ
��G8?�.9���X��y���Pr1�sGI�:Ǣ=�TA��y�AA�_l�`��4�eD�
��y�Nܤ'�fi*�c:-,�(.)���i�X�e���.�{��0�i��5Ć|�gB�dQQ��I�<
~ ��_&|b��//��+p�A^Fx��d|<�&Iu0
`s��@�����ȓy�|�"�J%��\;�NB$��!��hO�O��	�� h�(r��U!�#�-~�,B�	-A���� jw��rX�>�)F��+LO���U����sdkY�b����x�:9J����}�&a/���"��ش��?����5z��3' �<ty��E{8���=q";Of,K�&�9��x�����'`�C��x"�M"�h"�j�>��$�V��ٸ'�Q�`�O~���Q�������q
x�҅oPM�<yq�ޙJ���H�-X�`��$��b�h���ObƵ*�
�$Z3f	b/�2Ī�	�'�p�링Y�!Z����ȇ�x�eb�r�'���� ��'�0er���bR*t`���=�'S�Z��bܤL���б�+{���ȓ%<���懅L�N�@�l�d���OH�=�j�IƿtY(8��ZS��-9�@�W�<9��;c�D�㦎�K��91�$LX?	��$8��D��kf��3�eo�ȓh�XH�ͺ���z���y,ni�ȓ:/�Ż�-N�:���jWKυn��M��i��ZE#�:3>�|��ş�x�0��S�? v��b�A;v���R�.�Ԡ!�"O��KQ�M�h���.qv5�"On�	��z�Y�w�A!�vY��"O|�P�,�y�ؑ��6�'E*i�	�>�98��$z��'�_�B��	Q��I� i� E�D[	M���D_��(OZ=!��ڸQV%i'���_�ܵQ$"O���'蘹<h�Lc�ɛ�\U@"O�0�f-�{?rm�w�O'�d��0"Oܘ�A ���}��捨B�J�`�"O��"�DQ�n��I��ټG�@x�A"O�!�厳= Ntq�뇭3�"Y�F��PH<ɖ�34�L墖�\.8xإ�B�����>��j31��b��T�2��=���^B�<�e��'����\  t.iȖ̒z̓�hO1��A�F
 4a{ x��
+	gu��'��I�C�� �@���Mz�+ؒO�"<y�! sC��i�\�KF ��%V��G~R�ӱr��R�l�#vX	��-��o�C�ɾ4]Bq{4Q�}�530 ������hO�>�0����6'��r*�	��:D��ʔ/@�;: ��ԡP>�*���9D����+[�WĤ�p(�d�>]��3�O�	c?�5�>u|:U�"�^Nj��f\�<AS���v.�9`㕔��Y�*YoX��͓�MSH����NԦ[ْ�QqS.8��U 3�4D���c@�^r�Zt��/ly�&D��1�ML�JP���ޠh�Th`�?D��� �� e�Ȓ�@�ID.�0�'9�y"�'a�Qqv���ْ2"2s|� ��Al�<!@HH%SC��1WlD1���͑-�!������U"��)�����K3N�!���`q��J�1��<�e�	
8{!���h\b��>9�,H�fL8=!�D�!_��ȩe�o���c���J�!�޾)�V}s��D�<� ��F=
摟�D���)~���F���w���D�Q��y�`_q/��q.f#��� M����;�O8t
�	C�t٧�[8~���ٗ"O(�u,ǜ
��T�0�1��:#1O4�=E��H] v0�B)=G��=C��Q��y�C�
�ٕm�H��������	��p>I�G'P�z�˜=�ƨX�Q���F{��	�Q�j$��I_3o� c�H�jC�ɕ�p��LS�z��F(��D�',fx�'��Io�'���p�d�Zp����J0 ^�t;�'�<�c�߃)9@5�/G�vsve�	�'��M����-ƕ�o� u&��S	�'�*���ɐ��B�^>x(l���'����L��sipg�M6u���
�'�r0��C
���h��)0fŢ��'���i7S�\��9����sF@J���H}���� �XX�!v��z�$�!Lɯ ��XF��dM�NIv�J�H¬^�j�&�UK��;��F�(��Ƀ0v����H�8ٱ#�W�>���7�I=z5�<! �\Dݪ
��q�7m6�@�Qgȶ874�H��&i��IC�+�D;�OLq1b��$.֥+��6~�֍2��'�
,ps`�3KV��WO�(2N�lD{���'S�Ik���/�-��8lȎMI
���,l0�U&0)*X�ƌ�2�V �ȓBD�ppE��*z�!a���d��ȓS�٣g�D�K�L4��	
A���  � ,���S�i����S�? Pi�!ĮY.u#�`*.���"Ox<�8Pi���0$/�y"�"O����Fn���;Ds$��"O����kԮ_���`^�h�8 ��"OJ��:q3�)�U���]�x���"O�Z�dۇ<�4Y�D� ��<�"OF�@�ö+��k.ӫ`��� "O����'Z�����M��^�6"OX���AnѬyqK�X�@�3"O"�����L��#g �1k�"OR��'(�6p�=�p$ֱU�ڴ�e"O�$���,R���J$�CUBp�"Op-�Qh���	J�����"Od 	u��<�<�g'ÿi��C"O-��B��x=`�A���9:�"O0����6�lL�E훥U�$$(P"O�� �<{y�l�4g���H���"O��z�B�j��@AДv�v��C"O�@:��b �c���	�:Q1�"O�$��b��dx)�q�ȶ5�x�#�"O�4�S�:|z�B��}�B|��"O\=��*{�`�gY�#��9Z!"OTuh���]����L�nx@���"O ���
(c_6(H�I�!\l���"O�9Fl�Y�|b5��)	fr��w"OF	���' ��~I8���"O
ܡ�!����y6	ڬA~�h�"O�I�%�>����A��$2@��	�"Ot̀����� ���зY$���"O��s���>c�@d�CIN���"O�����n(��� �ش:62�"O��Ȕ���}��C83�P��"O�i;�i^1%�i��O�Bnތi"O~HS������,c�ψ0%�4� �"O*�(�CL5h�с�g��e,K3"O�)�ÁI�s9��!s��u�`p�"O�؁���c@)��eA�`�6"O��X�+֍%��
0�	&��1�"O�|�@-��8�L�T�Y��8�p"O�D��c���T	V���?!�#"O\)V
*��%�ƌՖ�d�"O,l�#+G�i$�=�SL
�?�4Q�T"O)���Ç42�5!V唠z��:"ORI(���d�D�2F/
>,	�x[F"O�EC�eM3<����$���Q�"O�@X7"�R���Z���_���"O�L�QiY�`�e���W�0�x ��"O��c��W����p�H��V�2�)"Ol����.�V��h �y�p"Ot�*4�U���T�]�@j�Ip"O�kaʟt�ra��7�*c"O򩩷��z�`�"���%M!�c�"Ol h�K�Dj�u�t�-<���r"O�=��.3{`*�SfF&��]b�"OƸ{���>���+BO�n�v� "O�B�̖2��baI�b#�H(V"O:��$��?7x2�{u�W*gra��"O���n��_���b ��Vk�5{"O�ႢG�3:)�!��>_�
M� "O����P�Z%<�x}X6��8�Py���W{Tڣk,Øl�`�"�yQ&��x2�ς�w-j|q���yb�.u����̛m6b8B�:�y�� 
p���Q���P|� �g�V�y
� �<`��٪4(���.��R�,��"O�њ��L�vTqWֲj*̍`"O�U"��׼���b��7X���"O�)��ɀ:�ZY�Ӣ������"O���ԴiÀa%�ɸ��(#r"O��!=A�m���?Ƥp�"ObpY�`	4o����>]���"O|��'��"�68в�N�z�6�Ya"O��� ��i�N종C��4�	�@"O*ݪ$�O	�̩Eb+� �J�"O�t���.n\�I�T`�#lm���"O�0u%�2� ��	�]P��"O��/L�	�D���[��URY���F�O�� F��'�B�{q'��N��[%�'H,��'�Az��ӱ'((e�L%4� 	�'���[L^�PC���8H���'� ��ϡ)Aj�S�ڱw{�ݛ�'3���%��!\0�Q��!��i��'0��u���V����$B5��'@P3�(T�-h^�qsij�0qˠW�hD{��,x��p��uǺ�{f-	3pa|�Y��h61�'hA!F���d�4\�����T2����`��ɵ-N�D��I�<�'Ƒ$�*��f�����q�Cm�|�<9b@EBF�����	2̅a���byr��)�'rr��Pʑ�U��!$��O��1�ȓdf�5�"Օf����ʇ$ L��'�R��9�	!�����M.U���"��_���f����-����A�9��A#c>��(�O��h���y�ųr�A���y��"O��KF�ΰrp�=زa��-X��>��9?`H��M%n����79����zkۃ1K�� ��l!t��hR���M�%OB+|;D<�C�qP��b���b������d�!9��W�IgO�t(��وTU!�9���@�/>GK�Y�CDQ8�!���4`4����+�2f;:��!��9l�1OL�=�|w���&�b�����/b�@a'�p�<��KA�>�4R�+�!:0�V&n�'��x2 ]�<�@���̨P�T\/~|m�ȓe ��!�h�3Kj��Hf�� :w:p��hO�>i!�F;U�4#��G�/���C�&D�T%�P/s��*6�D�{��)K�:D���B(�5xˠ��!��;��9�w#8D�[��X-X��<�/�o0���4��]���� T
7R4�x���	9$�Z5`?����α�W��<7�d0���C3X��m�B"OF(�e�$m0��(�Wt�SF��.�V�',rδy�4N��]#�BޭJ4�#��}!�jZ�|�z5#��p�p�ȓWm������m�:�JG��n�&���aR̢��ʷT�6)���M����ȓDBF����N8�D	���H��	�ȓ0b�Q��øi��I�D�d��l�ȓ|�ҡ�aB�b�.�aᏊ	f�lDx��)T/�W�4��U*�c:��V���<!2���0��^�n_���QEy�<�Å�7��J�©I����Tcy��@�<��)Hd$9+�xMD��Q/�z�<��$L�xJ�Z��^�+K�}�f̄x�<Y�GT�)�Ӎ��7�D�5�|�<�!*��;�H�EȖt���
V� o�'�ax�"�1��)P '���`� Ͽ�yR
�e�0��/W�a��J6�5��'�b��� �Pw��#�e����"4�PA�"On�
BDˌt��(3�Z��E�"O�=��$�$P� ��`	�;��Hw"O�����A���ͲRjB�H�q��"O�P��� ���bZ�.�n�c��KO?	%)�S�'8�TeȲ"�� �����o����؄��J�&�\8$��Q��K�aU޴�@"O\$�SC�9cr��˦ ��}O����'m��	x,�!�2�b�2�!$�]�L�!��B�_ 6d��c*���dL��!�G(2f��h� B�u��
,�!�#X]~%+��ݮ$Z$(0�G�n��|Җx"JV�B	����B�&��<�%��y�u��BG/Yht�m�!A��y��ȈcyPy ʐ�Y�F,�q�	�yrL�+m�Ͳ��L(
�$"�$˔�y2	���p�d��wo���uM��y���(~��tH�v�n�a�Ǻ�yҮ�	$UPၫ��P��jQ�y���YXjp�C��=�0�〄E8�B�	8�����	��Z�l��Ľ*�.B��	cs���i�5)` �b��H,B��b�~�됡~��i�T��n� B�I�y�<�����h��i��7%�C�	�(h�$l�7c�QP�բ%��B䉣`���ѡ��!�ЍsV@�#����M��F.�	i��'�\�OPF��#}�q)��E�x ��'������D�>�#P��OC�M�'��aB6 <o� �(	F<W&I���$x�dG�$�NV�+B�R�]:H�����y�#K�pZ�-C���mI��[�G��y�)� �ne�-�r���A#L1��d0�p>��N��x���H�fP����9�`X��h���'�d�FyZw�����M�O���3��I�W�$��"O�غ#C@�$�`k%�rH�t��"Of��r�Њ<�F�0�	H9�v��"OF��0Nֶ;�-T|
��q���7��'ў�>Vg� A���K���\U$�P��7D�,�C@Ȭ0G��0����]���7D��a��Ё,��Җ!�xF0��ҧ5�d[u�'�1OB�#�bڬ<�=�P��*t���4"O`�p���;<�����ƃwˌ1�v"Op8�L��.l��ig��p��%�'����7i F�`r&�^�T��/�._����Mܓ�0<�"��"Wz�����̅{�$�f�c�']�?Y��,	�H�CE3��Cw���4��	�@fpJ�ʐ�RtႮ� A��	��~b�>�O?�|R!�{�x�F�N>
���qUk�E�<�1+ԩ�M`&��13�!���<	�'��ON�=���6u�yz�GۨQ��I���Q�<�2�GE��Ē$��'(Q�4!�'	ş��	���>�G�C��.D�� �$<�Ό1A�KX���O�d��Z4R'@TÇ&��G�	�O��PǜrHb��h�%I)=���8��Up}B�)8�I��e�hV?P�@�;1aεYn|�ȓ;�.t�m�9K��Cu���2����,���'jȹ;�]+è f��ȓ(0�uy䂍:����w	�9l���DyB�'t�={��R�o@�)k�쟲!u�X��'�D�o�5y� �HRH͵=*��'��=Ҵ�ګFR���Ѩ��hJ� *�|r�|��*��
ė-�@�J��E,W��C��'W��aI��N�<p��C�/��7�7�S��Mk�.�`v��y�O7"}N���n�'E�mE�� ����O:M;�y�Sch�� V"O&����ػu(њ@���
��"O�I����w��9�R`���t�&"O��A�CA�~I�Pb�$����u$INH<)��S+Y����J�.��VN�G����<���B!j���5.�9{�N%�uh@�&X��'R4���þ���r�D@�ui��X�'����ƾ�@q���įty ��'�.�J�`��qt&\P��S�n�@5�'��Y[v)ˡm>��� T�m��=Y�'5Vt��.M(~�I��c�b�����'����
K;R|�P��&c�[�'�Lh#�nL�(�,a𡑛S�T ��'+ ���+)�X)i�j]�J��I�'�����D@�c�H"4N�Wv�lQ
�'�x�aߛ<�¤9t�ʉ<� %0
�'螸�-�:Y��Y�J�`:�l�
�'mLD���:g�cԎK�\��9
�'6F���P!𡃽F~x�Å �9�yRcF(bf�!Ǯ��2Y6lzO¿�yB�UO|{�O�$��x;��R)�y�m��nV�	ٷÉ?�hEHp�ڸ�y"���r������7� ITb�yҢ�l8X�L�84wvѹ�/��yR��-���ˆ,?X9��܁�yRB�y�����1�E@�V�y2m�4C*��[��I'h@�u�	%�y�@�/f8!'��ki�U�N���y���7c��	�!���]�t�S�"��yBK�<*���\ �Q�%ԛ�y"F�54z,��#�����	�-ȉ�y2W/g���$e)?���2�y"I�<�Z� i��j|���X	�y�芖p�=��D�2}��� eI��yR�(������ o{�a �퐟�y�e�O.�����-�<i���y�GA�?�vy�(�
�E)� T��y�g2a��ɻ��ȋ4�vU@� �,�y�O�B�,�HE���.��m�Ү��yr�N'4:��EOulh�����y�OC! ��@�a���%b֓G�
��ȓD� �r�܍{7ThYP�O�JG� 3�쓮@�����쎍z�GG�;���`�Q���؆�d��d A�1DmR�/ԖIbd�Ln�<)�gp��@ ��w#fE���d�<�ClثoD\u`e��n��l���g�<y���@��ei�g֬K&�M]�<!�	.|1Vh�",V�
:Zk�RZ�<Ia`[�h�h)�פ_��ҍR&	o�<i -w#l�Ң�5Lҝ�ֆKi�<m�&04�#�;̖��LYd�<�S�K�p2�pQ�O"L�6jTI�<I7��5]�d�3!��d�B}��A�<�ҧ6HĔ�0k�[K������B�<���)~rZ�#9�:��"�B�<aa�<�x���眝\`���#�{�<q��J"N�h��w�9d8�lw�<�5˔1( x%�Ȗu��8Tgt�<AA��ں��⋋�p�M��gu�<�Ł�p�HX���	�Le��b �l�<y���e7�p�,�	��A�Kh�<q�E��II�P̋$;f4bB�Q}�<yV��?�b9��G����q���r�<�U%�A���E�)�Rآs(�g�<� ��a�U�^\vhG�l��(c"Op�b],4�X+F�I$_�����"O�|[��O$]����Y�pp��K� �7�L��-�<A�n]C����[\ rP�"�X	^3n��Y<	!�$� +��RpL]\��䘓aN�2��У�����9٥O��8������>:\m�D��� ���E̖Xp�x�	өP�(���ߖ3^h�	��ώ-�j�)�l�&���9.��CT����RtTΎ�co��9�(Pa�ܡ�'��#��!'��s[c.6
W��q�'v���w�����0�F�W�U�<Y"$�h�d���EBye�8(�E�!J<���Nǜ}X,��g&1iH��|�O>Ѱh\�|f� �g˂2o	b@��ct��D��Ȝ�<�2 #q�[�.T�ЉP#
��܊�h�0.�T�%��%���'z�RP��RF���@��;`�:��d�A&lI�����yӨ՜a��DC�0ꁹ���8��(��kTpL��dvҮl�Ĕ�!��y;�`D;@��ɐR����WM �$5�e�2�Q����|�C眭9{P`ӕ��6W��y�kBc�<�i�xdh�UO�:xm��;We���rh�gᇕ_���Ǧ��vY�4&?����	|~��^�5���>��ջB)���?�##NZ���C�*�,� P���p��Z-|}��i�	���(@�(�6�џ0�*X06��Dr�f�)&�"	�� +�faP�&�L���ae�Ҧ$�L�23� y�C?���1���%s��$�Q#�w9��Sp�
���=�ǃ�K}��
�ɔ� �d�ٴQɟ쩔��.b�FUI�W�H� ��1��Mp��J�iT��`���l�	{>����B���
O@�6ܱC�ZX؟PCI��g
,M�E@��pt���Y�7�@��2��[�,s� V���R�n�**&Y� L1qz��QY�4�P����w��2��X�[3
�If�%�D����Q�:�C+Ɓ�?1�䞀-U��;%��m,l#�H��6�z7��?��Ƃ61#�,	1�«s*Z@ �c�j"t+S���,�"���<��dREÂ��X�|���f�	�A�4.�b}�uHW�ii� �9�$�����zA�ͲL|�C�t��݈#���L��)1������Y�k\;��$X@��� �w��͸��$�2�zhˤ�R�4��鳗���]�p,!L4J�2Z��?y,�e�<�R4�-$I��@ڦ/��i�d����İ]�\a�@�"\.ܠ)��X�$�5�
�=ڥ�"��5vx���$X\M�v�W�]a����R�Zuhfcեk@p9�ņZXw8}aa/c>De���V�_b�7��)(��ЌF�JԈ����R� #/N�	Y�e蒌%�.�P�V%�X�!s��!	[�}�2�D2j[��iS��6�L�k�
8)�)	,���@��>j�Έ�vH�g���20I�Q��V�:h� (1����߹� )�^�S�ɗ�Q.�h0�����%�qE�<s�h�X��L� 򼬳P�[���`2��e]�KŨ�)��ڷV���I��Kd���C1���7G�I#U�R��dxf������1�DڵS���� H-��@�����@�jQ�L��&��򏏄X<`$Η'Ȑ�(-��T� B�jM����
�4�*��(l�xXc�)ǘLߐiAu�)G`���v�F�T�v�>�ĭYP}v�
�&������Դ<Gr|h�Mf2�+P��!�JA�CDG�N9 �`¿��S���;Hh@tMՃd 6��~ �)�F�9����P��<iaa t�ASoǒ=	���M|b��B� �.��g�Q�l\Ru��*�D�<�Y��S�zQ՚v���)� P-3��P}��J׼�ѫ�_}PQ����O��Q��<��U'��-���4I\�����S�X@� ��PH�-X��Ȝk�$Q�1D�Sf�A� 6����,6�RT�`�\�'�h�� U���bŠ1�`Mj���OHp�O+(*B$R�閥���@ĺˣ�J���d�ɍ�Pn����ʄ4��
�kU�ȹe��4�� �ƍ*�+m��
祐�mmv���G�tq�P(6�ߝQ��e��Ky �dͅ`E��)�%	Rpr��'�q}�x`���W���O�̤Q��tF	��(�9���I���βMbذ���B�8���xL~��ρ�V&��� ���*a�`��*,��C5ڣ*�@�HӕY�����!ZP"�/�0	�w�TT�&�X�H�^����Ć!��ݻ��oP��DO�)�Jd*O�	�P��ИO6|��`��%^8��`'�q�ƍ�0�D��`����~�� .ݻVT0��O�	R.�Gz��x�V���e�|K@�Z �
7���K�}���d��o��7m1Wx�]�q�^T� \����{�qX��OOx�� ң��Z)+ܙ D�cbӞ?4�zb��S�
ǅU�:��)N�&֕�U�+rX^���@�D����_� �"���?�y�NH'
҅�C��M�4i�Ux���Ą�0NBĩ��!�H��V�u�HĂ'�P�_8]"B���f{ҥ1�mE�y��Ձ�'$�F�F��v�Fزw+��^<Q
2�cv�牢>��dY�E.;A���F)���d�/�~�Ib��'70B � �v`JEڒ�\g����W�A%����&)U�m8��_�Z�r%[���:�Xm����A�*��qsOׅ=�.y"#�����=\���t��[�\S�  {�4���t�M\�PS0E��L�����,U��)��l�u~LQ�'i�	=Ύ��D��Dm��y�l�t����U��>A�P4T�Tʀ0a�oO�XH�d�ıGl��Q��Hv��d��E�F[���n��Y�R�t�
�8`���:6���I����eHG'�D�7W�<h�a��o��ik'��?H�ԙh� ������ڷu��ۄ	܋2rA��OZ0j��uCg.>L�Ĺ�'F�	�KO�a}��������i-O��A��R.I�h�:ׇ�O|��ciٝ�8�ڤ(G�pzT9!�Ȇ�3ª�[�	�B@�� ,�!�q��[9�n�	� Ĩ�F�2 �'�Tdۄ+�H�����Eב�P��sȅ�L��6I�03���z"��}q
��6)֞E�T1S�
�%>���7�� ܝ�!e<-|*�k,0�py��'�Ҩ�CKe���@'�:?
$]�r@��1H�A��i�± W瀧,U�s%�(5����	u~H��e�<Qi*�j#LP0(��)����7%�<���L��kO��G}R(��	�]�Ҍ{��9��_>)��5�+�4l,�p��4h�b��w�Ѥk��D�b�Cv h����x}¦KO6i% ��m�x���A'm��d��\I013ѫ��O��MKŃI?A�)�Z<�Q��,�,F���4]J8)Q���K��e���u�`����vW�-�%Xvʐ�fr��w#V_��ę@�d�rf�=2hQ�EK��%���2\�*O(1�%'��g3t�7,��+��9�ڴ�MC�(�g�K�J�u@��tD� ���ȁF]��5&K�%F!j���E����mG�r(^�q2$��b'㏣P������
k�$)�p�%{7d]�z{�L� �G��%�
8Ŋ�kb@�8E�qp3C),������Y:"���C$��1<,��k;� ���ՠHx���O=���D}�nО�N!Q$�8V��+@�'���FD�^av��f��(K�(:2ƃ�jJt���*n�00�d�#a8<�V�Zkn6m�$]�L	�d�#݄�"�yð� 2oY'� t)N%�~��D���ȇ<y�3)F$�yrb��f2�x�ӠQ&>�|d�tߣm��s�h�~К�j�MB>7�4J��:P����i�]�g�� C%���
���O�S��L�����EF�=Hb�'Ȅ��c.8n��7%�32��
I������@��b@�$@�2����r��h�!�Ko�֘�B�+v�HB�L���<��	�[�P�c��
�!���rto\��Ds��� .��8�k_�C�֕ȑ�T0D\%%��Pr�^.D�֝�1�ղ@U�iB��%�Đ`e��%R��K�	�"�<�����*�0���ߋN����O^U�5�Y&��MA�"�`���4]ǔ��`gC<>����IEςm�%��u0��Cm@%� 8$LY4\Œ��aG�<B�K�^��BTsV�<�BL�z L�"�١��d��b���k��֊o�!�E�N�e	2L�{�nѻd�@
Q�V@Є&Ȱ���NV�IU� 5JăA�y)̋�y�O��ӣQ<vr:��aI��MvZi��	�������E�!|t,����84"�*T���ß80��q�]f�}��*^��# @R��	I��g��ЇC\bx�Q��3����¨�.z0`���D�S�?-����q�Xdt �oğ7��ͻ��.}<|�LǪ �^pRQK_�,o@�����yR��-���䗑W�`�
�����}�BIZ-9Ad%	��.!��p��.���ړ��R�p�"�h͆��]��B6={�X��,O.TJ�)�a$9�p=��k�iBz0������d�ųf��a �)�'zܞ|��@�)L@^43�+]�F�BU�M	H���TDE�b��M`$i�%~��]�~=�������k��
�P��>��!B0�`u�%�_Zi,xO}2,+A.&\���8�oH��,	��X�����M؉"�����i�B��,���߹J߆�?�� �5.)<ЈqlCt*��0�T`��r�h6AA;�J��p'L��Y	�!��b�#0�T�z�XpPkZ�Q��,q^R �jA�Q�$q������El�<��	�SU�т��7](D�I �>m{�e/$ny�%!��zR��H6H�Zuі+��]�bA ش6H���Ʈ@ ���(�,�Z�e��{�=�`��]؞h�"@7#���`Yh��R&�g� P�i�(�>T�aʪj�,@��%Q���zA�C��za&�b�|RUiI��<\���m���y1�S�Ӱlt�c�%��\��$���H�n,��MĢU�E.̐.*��D�.~���
�A�l��F��2� G��z�#D^��0$���O�9��E�u�$���GU���@�"HXD��K-�l�h������4v�,劰m��r��^��u���.Y����C�g�
A![s��]�W�ʗ#4<��dɰNf���A�Y>��S�M�#Ș,�T��	�x�EAB�;Xƈ:R,H�Kv��qk@'_ ��Ӆ�'��W���Kf̕|澑���
�Na|��D&SZD0Rk�
w"5�e�������3 d���@gҰ6]x (��
lE�sB��:|6S�eǁ��乆�2#cХ�'��1��G�8�5%G�7㊄��ȸQ��q7�˛A�.��(�̤{�U#7G�}ٷ#B�J��:���!iH�{G��{22�! ̮ OL5�A&U;r>
]�c#�+�fd����P��(�!��Fk�4SЅ�j~D폰>F�tO�[6��!�ƖS�����Ca��Ec݀��%O�?��T�� :x��JE��qg�ܱ��/K��O�48ƫҩo���K~��"X�D�������^��Hb���h-��sD�/���,�FSHYX�	�#�_OaT\��wg���[!����YLBҜ�Vz?1M��6��t:҆D4���d4{��C��=?ШXР�,jʄ!c�an���C�ON}�r&b?]c���7��`� ԕ.o�#5�~2d���>�2�$'����O�� @���Y��5MO�}�Fb�FE�9�������	��<Y�	;�諳�5P�3�ɕa�؄��!��?��Vڌ��hZ�$����'c2�bbLS�t�������|�p� F?����j_-}肕��F�}x��#�	O�����42�:�x��Ou110��?X�D����=d"P`��J�sdJ%�w��8B�~�=�W�\�}7�q���~Q�+˟����*]S,L`���`��1E��+���)��g���q&�T��ۂJ��R,THV�I�m�y�5��h�%LďP�����LT�}v�'�B�8K�$�H����`&񟪴�@��h��1
:z��\� �ع|WRx�� �����+��
Û�OʋL��4Q��յr�vU�@!��r���'�DI7�I�,��U�tē�r�*�A���?��I�Vq�Kƪ�X	��+��}��n�zᡋ�vp�ų����{���tᑰ
��{T'�=/�x)���[�I��\(�Gء?��E9J� '0���⩇ ,J��B'��'%�  P��*�`4�b���q�]b�j$4��ڲ	�/M��jg�P��u��˜2���!��4`�� �ؙ!�ў`�bG�>uj�u[�M�-�m��M]✁��G(J�p�'ڻr��r«�D���A�"D�V}��;��J,#�&�2��xݥ�;�MCW O�ZCbY�5�W16��Up��Z�Z��A�3�� eMD �1�'���Eo�8OH$V�D���]`���[��M��E�eLB4��އ"�paQ��W�,(n��g#�:H�s�V0j���b��~�,+D���1p��W�'�^h@#��h]�) �AD��J�ʒJE5�Zݸ���X�A���)�Tt ����oS� !�E0�XŊ�w���rW�(�<��F�����4^���3e:,OD(�SjΫ��� ��i֥�*͸�)V�|#Tp�f�bWb�r�Z�f\>0��B�'`j��9VEV!+Ͼ�6E$Zl"�Ɖ٦=+� I���I�� ���,ړ2��1�d'�-
R*�F�	r�4xs�݀L�����֐e�6t�V5z.�1K��M,mlAV̓�%�~a/	ʌɥƆ�hOj(���8@"p1��$�q�~���'��3�"�@�Y-9/U`4C�:E(d�Q$�s�x�ے�����QL�XR�aЪ��/B��qĎ��蕀��'Q(��1��G��9���
N��AB:u�� dN�Lɔ̠�d�,R ��ǊB���tL��D��:�w�%�D��1��XQD��+} >�!��`@/��ݺ�a�7� `���8��p��4ZP4p+�4D&���45�j�2kJlc�( �"�*\��LC�'��0�
þP�x���k���F}�l 
�<�3�O��3ߔ��/��^��H��D9=�Vl�$�0;�$'�C�T�R���n�8C��SA��r�4�iuiz�'O�l��J�.~i��
�-a(B:�'U.yѠ닖T�fS1
�8$s����	��P1	ֱ��[��Z�Pǀȹ �h�H#�2�����%ta�!�$�a��Á�Ȃ��b�8p�h�\�J0`̙�-������%�m���A�˄��R���yǡT����g5|�L���-���xҁԈbjY�$�QT�ǥݚlB�Ɇf�4L`�i0�U#zT́iaf�h`h]�;�M��=+���'��D�6
-+0�(R˄:�J�R�tt�z%�v���ԣ(/vIk�M�a���)2m:�N%��"7�O,�2���
Byl�`0f{:t!#�IX�dh6�� ?�N,(� H��S�fn�H�d��1��$2g$5�@C䉘4��Je*� @���q�?hs~���,U��*d�͜E����'�'."P�'ȉ��q�"LW�{�% 	�'jTȖ��&�Ha���y:����E?�����R�����I����䅄n2�:b�FO��[H�a�_�$�s#�;"N�-����)��?85���ɀjK���@�=`�<|��	S�4a*C�	60�Jq�S��:И��N9�C�ɇ�bhH�cF�]�������zӒB��;L7�`K��	\�F*�s��B�	�$ּ�ң��z��,�\ƚB䉀g�8y�U6d(,q��LުH�.B䉲j�@���?A4����k�rC䉦+����7�,t{���%F�C��@fiڇ��`�Yh�@�2�C�	G��ᙄ-�(vP��Y�&T��C�I �6۶nK��2��RuTC�I5	�q�R��vs汁�-U�A�B�I9�zɣ�΀R!���*��<z>C��%[�~��`��5f<���Q[��C�I�r�H51�Cde^I{ՇI�!5�C�I�d'��Å�ќ�����i�B�!v��Y8p+��h����F@�3�tC�I�"WnT`�ە-�6�K�BDNZdB� /v٣C�W���Ѡsj�}(C�	\�bX���u�vTئ���J>�C�I�]న ��څ]Vp��'9k�B�I%At����D	3,t �o�uנB�I�
gEB���t������`C�Ɏ0e�;�˖6Df�QqG�]#@�C��3L��!�۞:b�P��v��B��$t� '�-����r�� L�B䉼e��!�-�Ee���%@:F�,C�	%�ԫtA�rXy�JKn��C�	st|H$��%�)'FA�C�ɺd'B���T7 ������	�:�RB�ɣ0����/�"?��@��EPRY4B�ɤo�z� ��S�w'KQ�@��ay�"O 	U#�����s��}wB��"O���@\	'�r��c��?�J,+R"O���2صQ��R�О#����$"O���H��{+���$�jtZ�2R"O(4�!� +�L��3Í���X`�"Oܕ�SF��Jt���AÊ!3��h!"O ����;��e�U�P[��C�"O0p���B�"VJ�C���"O� �m�Pd�4r���J�G21�\C"O�P��_
c��*�Δ	c
h� �"Ot�q!K\�0��l�X���ӂ"Oe	`�mE��7K��E
�"OV�#fă�pP��Kt�D.��y�"O�,�F�U; k���)�:�P�E"O�I���m�x=bfhQ�O�R����q
Q���<A��{����[eb�R�eD�yL�C�Τp�!���e"8���0<W��%a�}8��B�� B�j �C�� _D��$��E�0�(�"���y#�(U��xҌ��n�V4Z'g�^��)Q>7�q:*�?tE�a�B�\�V��ȓhŌ��텇j^"�{��	)���'ԸH���	�3^|aMXb;���@���S]ڄ;��#;��#vo��Q�!�dȆ(�ni�C�P���H�/K���L��8� ͩ!�����a��)��D `�D�a��Z/OV$E����D�b�>��m\z�hݙ砑!A�d��e��A�w�W�|
58R�vX�$�!��2eT@�^��y�mֿ*џ4@�o��Lٺ�kG��6�����1G1
�&41�n�<i�F�E����-�xq�"��6��Љ���j�
c�@c�C0d;�9ȕ�@�(V��P�Mv̧���+w
�?w5lpKeJ-�ny��xB�a�2�A�:���4`�--�ȴ��%(l $�S
MH��B+�x�K���'�0�)�DEXp0�� =F�����pH�=nD����!R�:���@��<G�틖�+8q�c�� �����O�ib�ے ��4*��(�=ؤ�	�"O(tsr הC��l�C��"�cr��(k�%Qw�4���@O@�g�"�r�fu<�P��l��,"�I�@�t��2K2�W��?���R�	!��}T	h�9y�<9S5�� �(���T��������4�=R�J� D� XGI����?�(�@h��&��s�� c�	���s�nZj�X�[�7{�u��+J7���v%�r��3'����Q�����O��F��5N�w��esG�ɷb���c#]��n��h�Q{6Kџ!_���)��C�İ"����	҅��x�`\K���(%y(]��О"X���Ɇ�F�ބJ��5�
���:h˾=���(}��d�e̵=J��[#�v��7�N�]��6�vڎM����?��k��on�8�-�5H.�8s���9�d�QSdN�<xa�Ԃ��0��(�cOW�6C��s!WL(���)G<]�Ăc�����aL�4���Qd$D6TA�
8x̬qs	 (N(uB���c����w���3���!D�n�� ��:-uB�s��ˆ2-$�6�5��B���.ƨl�x�X �>}?:�� kP�
�|r%  ��������`J%S� �螿|?�6�V�VH��
��jdʠ� >y�`aá�;
�V剞jq`x�0��";p�|I���;����G�����rM��<�����`��o�@i�,K;+���#	�,H��F��s˶��bMь=��캴�A�l�Lq������06��	:�=��ŕ;*�u�VK�bvD�� ��^SN�C�B�i���Fg�8�����\��Ű;~|���r
JH2Ҍ�+��1yfǆxKZmIw@�'%��B�ڑa}x����O����X�$���� c�A9�bK!���x�(��rfl��k� j�%DE�@$Y䆗��`FL�RV	�'��9W!��:�r����1_qȉ�!t����d�zI�4�ŧ�����R�K�1�~@�B&�V oޮG�b���ǔ(g�9S�`�U���*tǍ5�b|���ܱ\�Ol��2�`����Z�d}��i����$k�A�&I�
j��҉:�)�YZTd�5`6W(�qB!�+(C(0�5ĄY
�]X��S!̘��Ă�XX���Z�j�Ѽ� X�0f���TP=�Xл��@�X�q:�ɘO��CKE<*���I��Z��0�)p� :�B���rI�u.��еBw�#`&Dyp�I��X�	�Pnk�'K��(T�H#O�IH#��%\*50��O�L��0x\t:@E��D�Ժ3����L����l2Ց��Y�"�Q4�O%K��`�"�ܟM�:��uɒG��"?񄆓�
��L�V)��r������B�E4S�����p���D%G Vd��ŉ�;w�59�IX�;�t�D�U�S�G+Wm�f�!���;�19Q��^�'-�ԃ�kI7l���լ�]�-wZ�}hc�˟^�� ��-2���:'��4A�Ա��_�%R~�Zc��-v[��<@����f�ؼC�Ě!��z�,� 8|`���۟��Z.���GF\y�O.�
$�O�|r��	43��QF	4|�~T*�M�-08��
e*^�l�d�GO��F�|�zS��T��5a�(ғ\��d��X+Z����@�\�H�<@�'�D#�'�Fu���i��V�W*fo:pk'�R)�f}3C)��>�ⱀ@�-g$ga� A�d`#��	
��d�:#���)�>?!��9E��Y/(�d��L�*��bR�b��%b�UFl���Ҽ;+��a���Z+*0���4ο��T�8�M�f=Z��9;��1��L�LqptO���JAɛ+t��s���8C��d�P��/�獿P��[�O���Ra.I*q��#��<)��K6	0�\�ԯ˒E�� 0,�z�@�'��zU�k�  �%��'Y��AP#ٰR��y0�C �Bi_�RX�	���W��a����態QE>Q�8��6�jc��)�� ��<Q`(͠!�fX`�#�@����A#�0��0r�j�p3����ΏҮ\�"ڴ(Od�b�����qW-�$/ѤI��ɤ/���I�v�ƉB���hoV}[�IY$�N�KW�\9"@PA��&մ���R�T=t�̙R$�lfBQ;1	 �R�3 �G�,�ܙAJX�Y���"	Ó(>�hxQ�S�`牉L,�9� ��1��)K���Ra�j�V��Z���ʎ+@�M@v��#k-��Y�e+Nɮ�2�e�z�U$9UA@ehBb*��nl`��'m�9��(F;���U�'CHA(CFQ���dC[�Z�p��D\J����`(� y������б�o�
��<�'X_HxǓcv\�@�ݰmr�*$��=z���&�U �M���^�����ϔ�8��Z�_�g�� �Ո_*|�P��w�bE)��ưln2da5�Q<~���
��Zb$ݲ�䃺X)�}Q����Q�v�����v18���BߗT�
�su��~6�cW�9]#�eq��8Q�t�� �>s=.��"��B�z̐�MG�Jޔ�Y&^>Q�\;�]�`��tM7��d��c�4@�( �O�Dj�#�$��-���0�0��>&Ș�9"�&FX#@�
C�	�"��yR$� 5�L8Fm���h�+d��l�#SF?Yӡ	��+%
�8`�ش(i4�"AQ1`��t8a�(�ec��I�B��`�"��cǬY:"Ԏ�`�!�/s�%�I=wϒ�M
D��Fxb"��R2�P���I�E# �T�j,Bu �o�~6MQ�>=هk[�P\���)_�#!����|���؆Sn%��O�M��#s�GN;�$ �a�N���H��I=36ax�GA���D�%��0�B1,G�4?��;�FA�^�(;1��4�h�s�dg,�`�3�H	S�G�06��#�f�3]�<[gH�Omҝ4ʓ�6�
<r$E�E�'��%�Tf+G�&9K��FP�i�#b=���7B{!\��V�H�^�9pf}#��K��jO�����g9���"{�R�pI;��3`��?1R�D�RfV�L�z;!�]�en^�K�'��q�V�Y�D��;s
�(}��4^�J j���S�d����{���Cԇ�{�Z��C�kQ�Fާ:���ƅ�禍a�a�7,�����#<о��>a�˳^�H-Q�5$,x�H�8rh�,��'�1� C��"���K���[�\	B1![7<82�:vm�(��N�������c���%7r����莍Z�."��'���#���$6l�� f��`�(b��	�t��i"c��bEN4���N#%o��S�&3f�� D� j�b��p��e2C��(P&D�nܰA��\��.
2n%�"?�A�u�r�E
�wS��'!(5�f�ڛ��\	5��	�U#0hԮ�A�.�PL�U���7)&!�V�Z��D1ED� �]ϻWt`�LבW	��a��RO̘p�'FZ)(B&ͷIL4=s���JM6%K�MU� ��rrJ�:!c8�ۇ�H��1:��^�#�r�2F�9]�(��!ga��bb
F:#f2��>9R�_�#��u��9rM����*�"���'�(�Ǐ�99Ad�s$_1/��e2gnɳz�P��#$�&i�P���_�']�ǈ�:&��PĆ�h���2B�{�J���4A})
Ԣ��R�P"��4���#D%��Q��Ր'v�h�n�Dw:�"Y�\=��"�7� ���Т��ip�%�1�YBD)�0��ȓ,�4�GG��f� �f[R섅��k�8v{�,b�ˀ!j�y8���8.�0�;�� b����P��M��m�1����GE����B0�'��c�Z������*�AC�M*6��Y��*�������A�T�
ӀM~��̫�YD�(0���>�S�Y@<�=�sdB�L0��4*U�zm2����`P٘��H<��W&�+_�4X��>*d�y�14��CDɜ:[�c�"Ƙe5D8c
?0G����e!��p�z��"�>�(����%r�j<�!8�8�0��W�u� lb�
F�'��R�Pp�X���s�p !�H��p��`�  �)K�h!s)D�`�\���'�����gU�R8�@��0_ν��	�JwBA�0%�
@W��"�E�.����$G�6^.�ܴPf��cu���|rǂ�"�2�2"r(�P@��d؞`��� �H�D��F��x1��
:Jf$�u��h���	q	�W�¹���Y�-��\���hu��?A~����j������.������F�*��R�TM%�>���F��C]��,X3�K�O�H1$�*H5����/�q�
�&�X�:�@�4��"K��d�:RɄ�7��  �	�w�����A)S>ٓ5KU���<[gI������?]�X�ZaJJ0p���Y�@A�V4ͫ��T���+�)�($T� ��� L��@��P8����Bԋ�����E!�$��pj��ɔF_ĵ�����������	�G��x$�]�/$��*X��DD(��BU֕��;I ���bՆ2��<sg�0>Z�P�c?^�فʆ( 
X`�+C-0|!���0���9�+.�.�����-<0�M�S�����B/|8n	�b��̤u+�<�/�#(�0�"NbXx�d�Z�'@b��Vϙ!#��OO�a_h�H�$�o��%j��ǎud>�S�+�1������[gl���»v�|]@3��j#�E)!�FL�'$�ܘ�k�f�0 ���%8�7hW�;�t�q���=���"�� �}�z��SK�b�<�Oܭ.ӷ�כ?�`�f�WI��!��/K냞g��������)�}���%u���Ӌ�D�S	�q�UjI$ �D$C�۲,���� ٶX��\�'^V�C��A2j�^�ĠYc�B@3&T��3`nE�qb��+@35��Zv?�%̙Z��Q�ص���d�Zk��Qo
�bZ�T[ve�E�`��
���e�O��9��&����g�2fR�tcŋ�G�X��~򤅭eCh��1 �=w���`mڀL^��{���3�Ɔh�<`�"ְ$?��x �N<zxp����<�C$E;.���PaR��sdQ�8MJ��b���p�)�D`œ�$�ɢ1���9�݉K<��ѥ�W.1����4s ����^�j�rc�\�Q
M8�6�W-Xh ���" `�Z���(�l��%�7^`�����k��H�?X#qO�X!t+.���k�7����Z�	Ǯ�4*0���5YZTd-�N�1�Ή���#�/������Y��{�d�踂*ۯ('���pi��S�� ����gLZ�D�:�<DZ� _��p�Y��%�S�0˔�h�N̕9r�c%bR3?`�S���_o�a�CG��T)8۳'v�>�����x��[�E�by���j���#
 ʥ���I�d�((Ajв~p�-� �'�� qF�C ����٢	(މ�(Ȑa�&( *Q1zz�1�@b�0B!y��Q$g�P��0F�	uy�18�!�s1]RO%�0�D��C��
��Z����P*����i�+��	��$[E��*d`�􈂖k��$˅��0Tpƀr�<O�0@Ɇ(�0�u7�΢���:�T[b�M�O�ў ���,a��̃tE�[��Ioڧat��(hN0cӀ3���Mڱ[��� &D110#���Ӵ=��h���u��27m�&8�}S�k�5eԘ� |�Ӗ�������9���G�'XZy��kߟ@&a�S�� }�~�æ��	���	�D�9�����V�hUVeqD �b���U�,�`VgB�4$�0����~r��3;���aF�'P"�K�ۯ2]z9��!�;�J��t���u�����#~<�c��OS(����,5Sf��ǃ?�X��w!z���2J���H�%4� kܴwچh@V�6,O�ܨ�ЊX���0{2�u'mN�am8�8s��>�|�gCu��Af�2�=ã�ױy1�y1w��bj6� Q��M+wm�<ys�� ��}�T�]k�'����&&Z9"B�03���m<�JW�ݿkb>Ա�ʔ8�bT�2� �"���	�~�@q��J�+{�C��o�.��*4�V>f<��C�\�֝a�-�;+�����6��ܚ3�P��� ��T9v�Q�®Y�¹!�Ժ*��)E� ��h
q�V
~����G�1;u�h�1h��hQ��	�ׂ��e��!q��H�a�X<E�`Z@�؛_�\<R��I$g��[JƠҌ���ʅ�w��|��پA�n�� ���D��/G�p�!% "�.��DБR�tOA:jհT� ���1�F��66�ڗ
��7m��&iX��CDG�M�bAT>xҖ�*f��?Gp�I�w_�8B��ڣZ�\��
�4�@">�Ԏ˛E6EC4+�*P�D���Hऐ���-:��I"A�T�`E���v���"c%�h��5���qg
0�O�0d�B���N"zȣ�fѱa�ʭ���Be:��^7��Cf�M�z�hI���0�y�H0d��h�ׁK�x�&��$l��$-��+hV2.��p�7
ΰ?	V��̀ ks
;�$���O�`$:i�W,�23����PL�>H���F�S~ΆsCj��"���^μ+p�9�<��࢙4AxL�#g��W<!`FC�T�%@�e��Zk�A�C̚&��5mQ%]�ɋ���68�ք9�(]�U��צ�b�.�wj�pX�:�/WL���l� n�`I��I� ���Ґ� P����S
�,d���f�jn�I��Z
9���т�'�l��D�.)@~|�d�k�r���$0O��liR�W�#80A�@�����+k���IT.�<|��gK���!�Q�x� ��rH)eeґ�B��i�"J��+�.�z�],1rM�F�Ө6T<9�K]�ܢ�r<i�ȓMϜ��DX ��t���Y}���쩟��f� *Β���0Fxb/�d�L�W�ܴQR� !2h�İ?9��~9Pv�p��5I�J�.S�X��� 
�>5	w�'�$ �R/��.�r��ĭA�W BY��'�^��5ŗ�7,���#�#1mI�'YȠ��H�Yv\(�S���
�DA�
�'H}j���%wID���ƭ�f�y�'�"���:z�|���\�x�'��=���G�����؊j��''x�:��	�I��+ӎ���N Y�'o�͂Gm݇ 	��x蒢
F �	�'ϊ,P&�D-�bؐ�xe���'�H�`1b�h�y�$D�����'���Cf�����A�{2���'��` p ��ؽx���+D�d�c�'F��AGb��B�R){�(�<;x���'}fy2p�!6�\�b�O*G���'el�ab*ȇH�jB��ڼJ�Ԙ��'��D8�c������$��q��aC�'
�T�S M:9 :�o�U �'�� �*��9i �b1Mߨ[Wz�*�'�,�Ӕ�Ԯz� �*_�R��z�'���*��G�V��ǈG�0��(8�'he{��Qm�x[��T!0p��	�'a���` �\ ��6	�!�c��;	��u�I�m����α>ѢfV8%����S����Xw��r}"�ƦP�ؑ�t̄:[��mY#<�� }b�ʐ�^*QsT)1%�:=oZ$O�Pzc��j�(�(��'�0|"�fC���`#N�U����M�2k4P� ���6ㆹY�a�殮�M��?Ma�Nx�96��p�f���| �k�1Au��*7}��閿	�@��ML;j<��L�~n���(8jћc-��S�(v\�Eꌘ-'�H� 璍<@�"Ag�J�%���ȟ�h�O�i��sb�p��mޙ�4�,_��fn̑���~��'aq��ͭ�VT�I�0��%-M�t��@؂ ��`U<?� ��0 "X�	�'%��ȫg�M=r}.}#��|�N�'����I�<?�I�OQ>�K�� 	�LhP"\$',�� ��O$x���$�Az�O�X��iȭ����9����' \�K�؂�����	8T�0��)�{/H�Ǌ�|�RD�v�À2 \�����p�<§�l�< #�ON�t	�e×l��=;���9��m��p[�'r,�Ӳ�O���K�D��y���F�(e1��H��x��P�`�Ɂ�3?� �a�c�[�1�`|�>{���BR�x��)7�S�O�:�`���EAP�U�@�Ih��� g��Gx���׬*�vTC�%�29�D,SehZ8
~ɢ��D!�p�xT"�&-^�#�+U)k��8� �DP�g��O�l��v�9D��hs��O�0�O>y��P����_��s�S�kE\�P��� Et�#�<y�c�j�kDQ>m�� T��)�'��m��ᒇѶoJj	J%��S�4�DiY0�A�p؎I?M�QCc����0|���H���)[4��
Gd�ǆ@t?��o�"�T<�0�im
�	2�h��P��,�k~���P:x8DQ�BMN������N��p>Q�׭>�0�c	΅c�uh��Z�<i�E�����"V����n��u��]�<����*X���C�	C(Q8#��V�<y��ƭ%�t�W�S)zp1S��j�<�a��?=�H�*�ÞWDYi�f�<�фZ#y����͹$��xI�Z{�<��/�$�KS���m��uC�a�<)��
jM�F�+K� �P%ɝZ�<��X�Z��Շ��_@&��A[Q�<9q&Z&��)r�M�]�P���,�U�<9U�Oi���ʅԴF���@�o�T�<!U�	�	D�g*E;_��h���f�<��EL*�)i��͹^lP�M_�<��hR�w���[�T�^!��Za�<)�C
N7v�p�	?���Zr�PW�<ɔ�!s����� �$-�M�O�<!$�E�܍�3 W����*�K�`�<i�А*�p���> @âJ�`�<)�C�4YcB�f��Vj�r�<��fќU��:���8�n��7cH�<1"�͠.�Y�v��O_���G[j�<�5皑%�N�+��Z� ��Pf�<�O��<=u�i^�ӥT`�<���$�h����Y)�u�r�^�<�E.��FO�m�f)�(U�<)��C��8Z1�M:�rbcJk�<�A(�~��`1��.�D`�&Jm�<9�܄qM6W�;:�!��G7L8!�D	�N�ށ��
��*O�h�^�A"O��a�Ǭn.������V�� "O\�3��σU���A�Ă�>��a��"O�4r��S�U>vغFcMS�da!"O��+�d��;�(���
*[��$C�"OX�'�4.��Tȝ4_�	�"O����HE�{#�%8�ǚ����"O�����J�6$ �Ҋ1�t��"O���e�ҳ5�%���Y�DC"O�1��HS9-��("����f�@���"O�q�cL�-�L�����M��%zB"O�T)`ͺv��D�6�W� v�a��"ON�+��� ���ŀ٣uFqp�"OH`@�.О�`ȣ/�i=�5��"O��ဆ�V�"�9�iф/+�|2"O�����gR>@ؒB
�z���"O�h�����`w<�!У����"O��SoH�(���a�L3��LJ"O��p�a�  �R I�NY���}�<�6F� {��iS�/�#K���f�N�<q�H�*.��A P|2��	L�<I��ɔMF��O7am*��F�QK�<9g�5 �^��pf�7 �lpCL]�<F�1Z52�B`"^�|�����c�O�<yĎ"X/^AA�.��uQc�"]w�<!��	��(7��%3Bd]c#Tq�<� ��cĔ�Gmr)[b(��&�6�0�"O�q�dbJ8�����Q�/�,�2�"O��y�N�)��q6m�n2����"O�h ��;�((�Y�SΈh�p"Opx*�! �4z}�a+O^�0��"O�t��cӳ!�X9�Ԋ͓Y��MZ�"OK�:�b̳w��Eg X����y�fF#X&��A����kԬS䂄�y�Έ�"��1w%`X�1�����y�`T���!&��S���&�y�c�.h���TxRIca���y������f��64�y��C���y⅕7��\�`���E�L*s)_�y�)�26/���S�7���bEg7D��E��TZR��� >���B�)D��0�oS������O�$���'D� @ &*��8��@[�Ln ��/$D��{�jJ�C�b�[ f�.z�HÂi.D�<�b��~8ļ��8ID�Q��-+D� ��#���4-Y1:N���
<D�������@T�M�do8 1�Y�d�8D��"!ˊ;P�e�r�Ԙ|�*D�@Pvm*%7��@�@G1^�b�j<D�lA�O��8
@�k����p�q��.D����ȃ�w~`��ԠCcT�cJ(D�������Mr��`�,��J%D���'��3`�����0
a��V$D��sc�P5z��2�o�D�Ek�F D��*ķ`�8���U�ek~����?D����	Ơ���;3t� !(?D�8�dJ�g�>�rVnY�m���fD=D���%n�6b���暱~x^Eِ�<D�����_�Ea�ٚ5,ݐ��8D��x��0�J|�w,ŧ9w.�0�$D���H�[���3b㏊=���VK!D��� �� �4�Ud�(Q�@�>D�<`��%�ݠPmOU�|����.D�t�qI�;�z��EΊ8c�R����'D��"���M;�踡�H�����'�&D��D,�!>E��8��,��C/D�@5jٙ*h�,(u�VC�N��'-D�p��ŕ.�fQ�æ���P�6D�$� `� v|�z��ڒ4�ZaD4D���t��"�T���+*��4D�L+��	���$@dV�Z�X��!2D��I<PD|SQ�� <I �A.D��+�)�?@!��>:cp�H�7D���?cQڱ8N}Poފ�!���6��B�E�)=;�U{�Q�!�ԅ�%CK0zY��5c���'��%��&ӑ}%е8[� ���٢�yCC�!��凟�"TQxsg��y�H�I��
��ѝ�Pݐ#���yr�L�x�� `�4Z�Yd�ڲ�y��B�"�����D1SQ���yb�?�f���*�"#��,`�F���y򨗭"
����G�E�����yri\�a��3F��:��
����yE)"ԁ4�F'4���Bҧ0�y��� r�feX �9Sg��y�� �[mB���&�)WԪyzuGP��y�l�_�ZMAfǍ�RH)j0�ͧ�yR� 8t�6Գs�Kg^���六�y��	�_fHm*�XC��wI��y
� �m�	R6���� ̹�b��"O��[��7����P���"q"O`�c��	�`9��!�W?9p`"Oh�`@�и8�$u��#(̹�"OrԻ $ݲF	Jв�l0g&�1�"O&�C��R����JU�	1Iq�$	F"O�� �ʟ�ʮ�LʯA|� �"O��僆9�(A�$�_/���"Or�R"NG�@����Мn&-�C"Ox�
4��%�LZ6$��e��		�"O`l�Un�|��֣ڠ�JDsc"O��W�,o�:$��� 6����"O��[g��~Z���t˲A��"O��!�6BLX˒��,([l5�u"O�����H��AhF'� (U8���"O � 
�a��9Qs�ǲwK�T��"O�%�rG�%WH���1�J�|RĬ£"O��i�*Y;�Z(w�L3�Di(s"O � V�$<��M�P���$��b"O�=��@w�?.H�C"O� y�m�H�0�D�Z*px�"O��h�Ƌ0�8&�#0��B"O(x�!�V�M>��[Ą�"8m�$R�"O�a����u���i~��Q"O����ˌF����%�y;蹰"OҠA�
���Q6N�f6�2D�(�׮�f��b�;����1D��n�_�@(e��E8dI���.D�$ˁ�̉�NUsl�0��Q�+D����g�����	�1n&�C�=D��
��ŧ/hh�%Ov��D���8D��j�/?[��� ���]]�`@�"D��y��k��͋)��L\cS�$D��E��\��5�f�¥B=
0H��,D���h�_�y������)�"*D��B擩�L���m��0l$c�'D� �w�1C> �Q���q�X\1�o"D���B09������M6?t�@W# D��
�Ø�I<L[��H�C��'+D��C �ǻzL����@�N�h"�(D�������p��C�bl<+eE(D����}n�����^Qk.�'(D���׌�hw֝xΝ�C+H�%H2D�\���	��1�%�Q%!8Pգ��.D�ȱ�\��=z�P-d,1k�'-D��F³|.�����/��ؑ��(D����	ـ�ѥi��J��Ye$&D�0'dݳgU��!�H@?�����0D�d1ĩߍn�)��B���jq�@� D���l� j�#�.��k�@���=D���C!$}�Τ����:3���'".D�$:��ׄ�.؉n��p:i��8D��#�)H)i��`C��W�5$�!�$D�8St#׺E�������Nk���'D������4�p��!E�z��"D��AnU�ee�z��`���>D�,��}�LAC(!��6 �P�<�����ƨb�f��k!����E�<�s�W&;tzL�\@��CE�/3.VB�	�6 l��Z&�&�kC��4k��B�y@����j0Z���!M�`�0B�I-h1�%A�� C|�\�d�
�+�B��F�\���2F��=k`�	�a�TB��:oK�	в$��Ai�hʀ9\rC�)� ,ݻC�����c�T�Q2"O^	+f���P�Ʀ�!h ��bF"Oı"�oA�J���#έ�2��"O��P`��4��rC#nx�YH�"O�A��c��T����SD7Hiu��"O� i�a�H���G�K���"O"$�4iw��)��"3VJx��w"O l6	��dM�4�ԛ8�&eˆ"O��Ӥb8Rء��	��!��"O���V�%8�	���9,�R��"O�r7� ~ZM�w�X���Y�"O�x��,B���b��'y֕�C"O<@��[�\*�cU�فsOx��&"O8��.ȋ{�5�F�/U���J�"O���	4:�9�+^�8��h	�DO�M�O���;J
1�1O.��t��H! a�1��5R�¨��L[�|�x5�G��+�v��������v� T��݉�8���¢]�̐5)K)e�j��)��k����	a���B��7��7�LqӞ'-T� a�����J-$;,���_צm�.Ol)�1����?!��M�b�BM��T&~L����Z?!�}����?1C� ����Z��ц^�v�x�V������4���������ؒ@L(��6oFxA$::�!c h̤�M�	ϓ�?I��#���+t�?�i�Cf��6����ʓ�~���<V(�B ڍu&��Í�đ�m����%#ѯ=��`xw�\�z��� O��f]�m�rB�w����MS��Ϛ$��lIV!݁$�zh����K!�H2�'��7��Ŧ�IMy��'��	H}"��|Ulၬčt`d�S���y��P1b.���%B�h�bв�#�B��O,m�M;(O�Qo�Ц��i��cJIXX"��)��nRƙ2����!wÌ�両u�0s	���p�͐C��sDĥ3����CDgx4�@���s���<�5��D�@�J�UX�4��e�h�b��6I~}IP
P3ֶ	[F�
��(�FzR����?�7�i$��I�	4,�K`G�#%RD�VI�)j�$�I��,��K�S�'/0�(8�$x.�pP-ݽi%x��gyl�$��(%����hE7t����b��FP��`�@ζ�M��?i.���sdy��" �J�l�����}%�p뢬Q� ���t���f�-���rS �[��i�0燌IJ�R?Y�Ɗ1^=lM�cG��[88���"��6Ǡ�QV���
�ŋʴ�|�qC�o5z�S�q��M�b96.D2%!�\�.OnT�t�'(t7�w��k�K�y����;?dl)r霞��㞴�I@���ē>BJ�����Q�n�+�EL�g :���I �M��iX�'t��ʤ�R�2f�|�6�F8h���JA�\�a��ByBd[/:��T�I�yU��cϟ�'ٚ	B�j�7�7���|8-³�+{�A3`�ö����R��e@��y���3G�H��Q	nkXvZ�j�@�re�	�����F�a�xA)��tĔঅ�|�*9#և��a�����l��'r��<�'�>�8��|:˟�'/�89��G<vZF��Cb�K����ד1�qO��H��P?uѶ�b@&��4���B��>!2�i6�6M7�4���I�>�w�ѢC�baڰ��[�]Kկ} �ܺ.�=�2�'��'�r�]��x�	�p��
�~&��TA_&q9.H��m��'*v�H �|5p٫�#̭=�^|Ad0��<!�0T�0�@��Q��h��NFE_���s%�:!��9����dQu�2��Dx�`tQ�d,��{#G�.�$��@��?�i6��O���?��}"+�m�l*�mA9T���GE�!�d}�	Ο��C؞�2G�C�V�f)�� ��i��dY��+����d��ik�'b��֟�N�� " �  ��   ,  �  _  �  +  �6  ,B  4M  YU  $a  �l  �r  -y  �    �  H�  ��  ʞ  �  Q�  ��  շ  �  Z�  ��  ��  {�  F�  ��  i�    x � C# - �3 : H@ �A  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P���Gy�|bc��@���sb� ~�֙s�PR�<A1�C41Oԙ8��+����"DO�<��J_�l�9
�/ ��|-h�%�G�<���X�,ʠ%�׮K#?䄫%��w�<����:�����j�De�F�Gq�<���]�1B�e�L|D���Kt�<Y�gT�I�� �̓���A�\kܓ�hO�O���UmS�.Cx,Jr�T2|2�	�'L��C�@F' ,ȣ��:�R8a�J���'/�>�	.+z��C�MP�>4hl�)���d$?P膟'$L��UDދQf����<Q�4�0?�� ����9 SLъ	�\��e�f�'�ў�'w��0�&�I�P&l�X��T�\���XFt˃e�*;(� X�e�2�`���hO�>��� /�m�𠉯{�~P��I"D�x��+���hp���ű*F���j }2�i��T���'Jx�bMMK�H�ے�2���?q��
;]�R�xu*�;<�|��r�
z��p=qF��0̎�Q0�ٴDM꤁���w��ΓS�b��%}���4	����#vHƭ{u�s�<�2fն0~t����[�u#����IG�A�.7-'�� f|h�E��49X�@=<���"O8m��Ox�B�#p�ˊ���x�O�����E[P
ڷͲ���E�lW!�d�7_6�X��%��b���	D!�O�J��M��R�ڍ��ˡB+!�$���Īק[��|@��P�M!!���l�\���ԬZ|��H�� !���Z� `�
�I% {�'W+.�!�$W($D��&͒�MRd�%O`�!�Dε��}��m�l�A�,l.!�$=b��5۵OJ	[2�QH���+-�OO|�<YF@�s�
x�V#A$~o���E�FG�<y����#�B6��t�$��"��d(�O�͒fA(}����V@#u����7�'�i�d�z��U9��F�$-P�E�,d!�ϲj7dPa�#N|��c��W��$�=��X?��.(i�1�/�����C�4��I��a�fyy��Ed�M(�ͬ5,HΓ�(O��D��
�,F���ܙm���z�K�$�y�&��p�jR��zd�C�@�iԢ=E��pʔ�g��oB���D�VT�G�M�3i�?��8���͠'��'��~�'�3sI�B�]VqgC؊���hOq��5Rb�ؘ}X�4p��Yh?\p"O�� tm�]��"��nQl=�S��y�I	8��	��lR�0�0c�,�x��'�Td@`AҰI�=�G�
,}�)h�'��ф��'e��B�7m�f#�'ɰ���K�G�tQ�蒛W֮L �'�
=���=\�X���Hd��'G�!3R��l#��Zg�N>:�jL
�'Y�xƅ�B4#w6�b
�'�=��.A\�e�Ӭ8���	�'��|��dSO��Ћ�k��b{����'�:�Sb�P_총�g��žy@ד/� c�L��,��6�%.�
�GM.D���Bkק�be[@Ĝ-r���-�I!Q��O�����NF+��bV�E�DJ��I�'<�@�� �6B#���T�8��ph�'sh�Bd�#$Ⱦp!��D|[�d��'=|�z$� 6B"n@��D�F���'0���v잛�`@ E�
q������E J&i��ᓹ%�2�&�C	S!��ٰC��M��m�=l��5rĊ��E���qyz<:��^�`\�e�GaN
�yR��4PP��Cm�J��рGC�0�?y���t�&����Z���M�5xIn���Iz�%"����'m���I1�0yݰ`�';a~��)&�H�M�6�J�Q%�V�'�ў��Z�Ѣ�ʛ�T��R�V:�`X"O����*M��@2Q�E�=���С�I@X���@���h*%��$+D�ۥ+D��
�A� �X9���.8�ΡR�*D�|a'% �q�0%�`�b5�gl,O��N�[	&�13�U|"�T��l��h�ȓD X!�R��*����-�
FY�$Ey�3O�6M,�'YZ��P���Y˨)T$��U)r)�ȓN� �C�e�)M��������x�걄ȓY0�h��)K�E��D��[�j ��	�<��4BHt�`�\��d	�� x�`P��	���S�4S䪂�
^P�aF?l(�ȓw��U�1L�:f�H��B����ԇ�1L%J�L�%^�R7!T.cB|ɇ�!CB��d��|���oS�efv���S�? �Y�C�'!�@�SV��+U�VЀ"O����K�^0Qc ~�`�J�"Od��R2x8鯤>����PFܓ�hO�OA��r	�wk����&�/VD��"�'T���B��%�}�,��� I7�!򄅯������'9۠��A�_|!�_[|z����(I+����R�2e�O���D[(໴	u��X'�&2U!��z���Rc	1�<�at�^�,N~Q��E'��#�U�?%$�i��]���0�>I
דZ"�4��E�82"|q���P(q��B���Ȫ�B �Q���cφ�@�h2?�O���đ(0����� �P��b^1B�!��؃3��l˴�R|8�(Ă!p!�8EY
|�T+�%:�L�	G*�Le!�ͧD�ּ�E�ՋʒY��%d&!�ϛ�P�s�M��(�n���G[�2!�$�*�pCd��{����e�M�!��Y�<4�۵���v0R���2��I��HO>�1�@�7*�2���
4�6A��;��S���'968#u��I
�<Y0I@�hh�'��6��O����!lK��{P��3tނ��a��5�����>���p���m�#W�qZ�O>Yjš�"Ob(��.גN�.I�N� c<�pC,FKH<��6�Hd��"B���+0Øo؞��=	���(�����HC+q=��#GC�n̓��=A��G6w��"W)XԮ�{$��n�'�?}8�;wx�̚b�E�y ��4D��!���9A�P	c%�͠XH�3D�.D�����Q�ً���/`!Qk8D�$�� ��ʉ !��dq�#�*D�|��ɻ;�9��	].�*�
�!5D��{�Lͣ���Qύ� IpL8D�tQ��K�z�#��M�aFu��a3D�|J��ք{�M�q.$��8&�,D��j��ШN�\��� i�����)D��A�խqĺ�����;D���P�g=D���4��v6���M-�`�V�>D� s$�"t�5MT,�ӂ7D�(�W�9P�$��CE!�ȩK�K'D�����" �4���#F�<>R�6�&D����&� A��rяB�hhN��@c$D�<��N�AiD���*�T1d�5D�ؓ�H̚-q�@���.�J�4�1D�"	D�(�,8 �o�N�p�r3�*D��x����#0֭rBӦkC��
��-D�T)���r�j!�㥐�UӐ(��e&D��G	R��L���@��z��7%2D�0����(��ŀ@I��gy|䙆�/D���R._W9Bq�Q�@=&�>0�G�+D�,���� �BJކO���A*D�,K�;�h<Y�o&zB �Ⰵ$D�̀��5n|��k��Zk��A��/'D���%��J��E�FN��`�$D�ta�%V? �v]�æ�	�%"$D�ܫ� �/Uʄ��g #.~����#D��XM
�y��Zb�^�FaVM�R�,D�L���q��9Q�D�1[�����=D��UhܮY����C�Tj00(<D������J8�
5CV8!�$�Z��.D��i�M(�x#e�:N�����-"D�X���X@F�	P�V�!�-�>D�����+Ņ�,UR�b��Lg�C�	U<��Ku�%i� ;#��|��C�)� 8���L��N�R��6'��z�	�"O��j��;dڙ��F��w��0�"O@qV�PWW���I�^���7"Oޜ��Kg��q���"e�6��V"O���"�ϯF��؋��0[(�5Y��'{��'E��'���'�B�'N��'NP��.�,v�4��% ĺ\��E���'�B�'%�'I��'���'���'����+a�J��S�ل@���'�B�'z�'_r�'���'�r�'�0E�r%�3,�8yS�C�l&jb��'��'���'�"�'�B�' �'����=�F=d̷V����f�'���'e��'�r�'���'���'�Qz%A%G퀤�wh'$>]���'N��'�2�'Ir�'���'��'
�܃�eMcQ��
�<`��ؐ�''��'�R�'���'��'B�'� A1,�7�����O;P�5؞'���'��'=��'���'O�'�$e���N�d�ƨ� ��.�< b��'�r�'���'�R�'|b�'�2�'κ\FB�j^Ͳ BJ�0� p�D�';2�'9r�'���'HB�'��w5n1:�k�'(�SӀʨU�4b��'�R�'6�'J�'��'_r�'�V�8S�	hv������(�r����'
��'���'���'`r�'�2�'H���ϋ'=�8�k G��A���ɧ�'�"�'��'�r�'!�loӺ�d�O����_3,> �Zu�יP�T�w��Jy��'f�)�3?)��i�4ҡ�P/ry���eN�lر�N.�����y�?�g?��4]�z�`�/	�-�i��0O�,��iR��+:6͂�O*CsOA�j^�xL?���G&���/�v7 z�E6�I��'��>%���+-"T$㠲B�3�.D+@��l�'-\b� ��ž�yW.�T0g��.e.}3WdT-��d`�F�IeyJ~�" ��j�ΓG����D�8Fde��@�;M18�̓TNP)�^"�ی�4���ܖD����K� b��Wh؆,��Į<�N>�³im��0�y@4n��	Y�Kٔ.��aZC�j��O��'���i��d�>q�hN	���K����:���"��V~"g_�v��`#����Ö́x��f�JB�v���a"��2Yj��:��E�a���|y�𧈟�D�0��b�,�#dx��A��\ ^��%sD�/?�E�i��O�	�"���(��>���F���A���O7M�OVib`�W���Ib�����1LDب���'��c�\�mn��S��M���dU��'?��Ə�6�J :��Z�8t\!�d�%?q��i�� Q�y�i��;�.|���#c h 3��i4��'��ih�,����� �j��=�`��8�m�f4@}D���%�2�ɕ0�E�s��'��U��>�������K�7$��A¬�+���I��� �'Z�o�	��M3���<�r��!s�`�s�=��!���<��ix�O��O�$cӌ��C�~�D����Nka�|�F��:$�f�[�z(󤯟Ћ���>L�h��O^����[��A�.�� jڒ23��3d��<������<E���W�Y�AM����7d�Ș'.�6m�1��I��M{I>Q3%��TG� �Fi�2)6�M	𩂣�yRT��l��M���
i !Ui�<	�'r];�F+Ă��P'إ<!|4h𮓠pn�Q�r/�_���dY���:�\��5M_�Lή��%S#���n�ɕ�M@��j���I��H��B*&f'�L�偁���	�����ON6�}�l'>���{�x�ˤX�t�aH͢.O�6�
'j���@�k~R�O�D�3�;Vu�'���ƦT�H��IK$�2 `U9�'��6-�&&JpD���e���N��5N�l��O��DSϦ%�?Y�W�DS�4d��yI�#$�8�����0�[�x��i=0}�w�S5�y��'�v�#P#��MS6��T�`��O�@>�Z�ĕ�p��&f�T�'��{�G+-��!2���N��hk�E �eVn6�ò<B��O��d.�Ӳ�M�;`���+q�F= ��芔B�:�r�49+�vo�O ��|����j`�E)K�<-�DWՐ(�$��ۅꘛj
�iΓ"��x�r���_�.��L>�*O2�u�f[���P`���*�:�v��I	�M�� ����OL=�,B+��Y��,��9�G4�I��$�٦I3�4`�'Jf9�&�����[�O�Iʮ0�'����T�AJ3:��?M��)���(��)V���G0��	#��J�V!�_-+;4���˜*��i������.��� ٵ�Cm�\0C6:B��X��<�0��m�Z�T�Q#�	}��(��H��=�@�D/��%��'�H��A&���+U6�R�ڇ�}�R��.�L�
eR���gD��1��Ä�z���*R*���i���)�+�Ң�.�N	��bo�h��03���.�	yRBİ4�~j'l<	������-1l\��m�|֞��#�Ԉ _D�xAH���+�ľ*� ��B���6�pٴ�?9���#,u���d�'Z�X� +0LX�"��;��N)G���^��M���>b�h�<����?y����$/��d�p��mb���rE:G�5�"��F�Iʟ(��k�	Jy�A�	6��f͠U����fМ@�\;�yr�'^��'`�	4=X�"�O6�A����I�M5��@)�O����O��$�<����?I��MJ�4mW����Q�D
aj��������O6�$�O��Mˮ����� � jiR�JD�U�Mi�+ՂF� P*��i�r�'��	ٟ��	>2b>�J�iA%h*����
SFj�:�ͣ�M���?I)O2 XG��t�S蟔�s�9CqG�@
p��3�cB��p� h����?�o����|
���nZ?.��x�n_�Q��Py��O>3[L6�<���T}�v��~b��
◟��u+B�m�n��l��a*����~�l���O��7k�<�O��L<Q��>@ș��� �8]��妭 ����M����?����2f�x�OV��Z3�ݯ
.�8��Θ�u	B���n�`��6�<A���?��g̓�?���S�4��x�0L	>zU�����яIm�v�'�'�
��-�4���$�OL6F�;��I��6���xrBC�����ON��N1O���O����D}+�F=0���&��C��lZ�0c �׺���|j���?�(OF}S��2` ���̴%d �`t�Ҧy�	7"�c�������I@y"��c~q��J��'�q�.DD�T�b��7�d�O(�$�OZ��?���.DLP���]>�+�H��O��c��Cs̓�?q���?�-OD� �D�|Ҳ�l��w͜�s��hw�+}G2��?���?1*O��$�OfYs[?�(�+Ƴ=Z�X��FK� ��t�$��>����?������\.2�
e%>�!��.% �T��Z�����fJ���M��������O ���N�!$�,��n��^�NY��4�?�,O����8o�ʧ�?1����3N�5�`�`�ݎIMU��*ҌMo�O6���%p(�xV�T?i��BS�G~����bI����"ʠ>���0����?	���?!�'����1��B�I� ؂1�RH�P����/u��p
a�=�)��}afeJ�GW$zaj�y�	Y�OE�7-�!b��d�O,���OZ�i�<�'�?a2�D�T] HpԬ��Pʼ�h��ᛶB��6qd��y���O�u�D�+����c�0x��KU���)�I�����$H�������'�B�O(SƂ�Y�>�i�+?���s���J������':2�O�����ug:�P�I�:'v٢��iRr� ���I�T��ٟ��=Y����1@@�� ޟ`{@y��x}��۬. � �O��D�OZ��?Q�NG���H����Slb��p�B�L��,O\���O���1��ПLQr"�W�`��@O�8c|��eˑ�NXPM#��4?��?�/O��d��s���r�2�	�,8�tQ��	"�V6�O��$�O��`���pP(衶Hc�&�a�z#�0�B��A���fP�h�	ϟ\�'�&���(��D�u�.���@�n���qƟ�M����'y���4`'�E�I<��@A�R� ���O�%*��He"M¦��	hyr�'b�3�P>m������FRf,�f�ФJ6ăR̂�"� ��}r�'[�q�@�D������¶8�D�X�Z8N�Y@`�������t�ϟ��	ޟ��I�?���u�D�yGq��˻�yfg�����O��r�+�Dl1O����C�L+j�����B^�r��i���'(B�'=R�O��i>��	?t����X� ����!ݐq����4cf��S�B�S�O��K��&�PYc!��6�V��q�C�D7-�O>�d�O戋��<�'�?���~(��Y�p���AW/a��0��Ѿ9Lc�dI'���'�?i��~� �؞D�g�R�~/:����M���j�lB+O��$�Oh�/�	�oP��eV�=TѺBA9��f�d	Y�g	j~��'�Y��	�Ch��`�-��%��5^޹�򎆐ZF��?I���?��B�OE��C&d�h)�t��7t�<A��i���3�O����OR��?�6h����,A�'�P�y2�׷?���b�!�M����?�����'��	�"5�7햕`��fpa�o�+\OB���Z�h�	ʟ�'��/�4Di�S��[��#<������;-�nX38�Mk���'�bI/JIAN<��h�I�����T8$<LA�f�Φ���Ayr�'��$R>������ӌ=pT��.k������8�}�'RְУ��9����i1E	d]ᥘ���A#bT�S��	ȟ�J�i�ϟ���`y��O.�i�Q1�V�ġ�B�=S�~��T��>��X��	[�S�P�P�/_���a#BJiV	o�0��9�I�L�I�<��wy�O��*��O����)(�|�p�恻�D7�? �R�����C�-+�:�kq�@>^"=�d%ޣ�M��?������,O�	�O��ı���d��%6���kC�I[2����I#��'_���!!6��O�����(Yc��?	��9�6�A�z���Jsӈ�d��oфʓ�?9��?��{���k���G-�~�(Tc�����$�Oa�谞���I񟄖'��I�c��*c��$��]��DQ>�$@&_�H�	ҟ|��x��?� �^�4����f��mI��*�D�O]���D~��'�b\�h�I2#@|���.Ђ���4��јT�(4Un�ǟ����<�?q�M|�)��Ӧ5ҥ�H Y��t�n�GDΉ����>���?�(O��$�	&N��'�?qr�	X�Zyˣ�V~�A������'i�O��䟀]`��w�x�,�j���G�fn)g���M�����O���䢡|�*O��Íg���3p���Y�cO��@��,�>����t�z�!V�S�$*��Y[9F��:DW�t!���9����O��3pF�Ob���O�������Ӻ� ޱ��F\<4N���#f��v 4| Y���ɺ9H�W<�)��	e��4�$��E5v�pS�K
o\7��	���d�O���O`���<ͧ�?�f�ɖ?(>�Þ�{�e*׮)؛��U94��%(�y����O�����˝d�@C&ә�]�4�
��I��@�	�G�X�����'�B�O�{����f���S1s����OܓC0��#O|���?1�'�Z�1�B&>�%;'�^�>��)��4�?!E��3��d�O����O��H�@�+O��A�B��<��ĺ>��ҙ����'�R�'|��ҟ`"��e]�1�p��s$ApԄZ�8�2T�'��'R���O\���y�8�RMS8#�<�"�/�^O�Mbf��X����T��Qy"��4yI����^%�S�]���+�)�BV�ꓠ?�����?���
�r����B��)����O<����� �.s��i���'��'�r�'��t�UMxӈ�D�O&�`��Ŋ5t,M�.� 4B̑ i\Ҧ=��a���8��=z*�1�	͟��ɚ�N�j��<xL0����$��X�ٴ�?����d]
`(�8n�h��ğ<�ӯFN )�.Z&k~Jۯ��%�O0�D�O|�$�F��3�D�?y	��Gy�4xA�ǈf�� p�e��x#�;�i�b�'�B�O��Ӻ��C>B������A&=��[0O�ɦy�	ڟ�hԣa�h�'�����Gd؃�˶��!����B�&� �66�O>���O��i���$�O
��V����J�X H=��U���Ho*����?�g��?�a/��g�Ĺ(T�Tu�2<�`� ����'�"�';敹��w� �d�O��D�O���� 4�i�6l|���)�GH�y�Z�h�'�����O���O$�$�Od���]�Wz�)�)�">�< [W�Bߦ��I�4�&eCܴ�?���?���d��G?���>>�p�y��˔J�5�ԩ�@}b���yRX����ٟ@�	���I�s��JE���J���D�@s䮀�M���?1���?�Z?%�'���ƥ�$!bQMݗ�9Rb��>���C�'���˟��I�H�	ğH	Cc�M�'i%K�fU�/l����l�6|y��'���'���'��	��B�t>i.`��@�C<i	&ЁA�ԶT��4�?A���?���a�S�ck8p��4�?Y��H��r����DU�r�%]��L��i7��'RRT���I<TZM�'���L@v��1���V�h*��)t4�&�'(�Z�T
a@����OH�$�� e�D]p��ɓ%T>{��	�MFa}��'���'<<9�'��	����+�60j0,U�RF�3��Y�:��m�Fy��A�6��O$��O���]T}Zw1Ҽ�Q/�d�yc��  �|���4�?)��ߨ@��?a��?���̊SxNy�K�`Fb�t	Q��M{2K�B����'��'k��Ƿ>1/O�j���1�
�2��+J�i����mʤ$9?.O��?��I��P̪7+S!��sā�	"@(��4�?i���?!b �YP�IayR�'����nĎYA��\k,�!�P�;��|�芘�yʟ���O���U
$٣'��^���AN��vg�	nZƟ+u���M[���?���?17V?��GF����m�L�xaQfOS�r��9�'�
���'���'S��'���'��$D�o��d�$�qZ����I�*۪-��Elӆ���O��D�O���O{���@�8�0�Ԇ�;�DA�������ҟ��Iʟ��I�,�	ݟP���>6mkR�p�6��=�B1Q!g�W�2�mZ�	��	��'�E���䄓�*/�I��� P�d`1!/�#P���?q��?���?�"�+,1�6�'Yb�_�B�����D&;dHc&Еo�p6M�O��D�O<˓�?�hQ�|�L�xcQbѺq̊DB���6<�>�#B�j�0���OZ��Ot$!4��5��韌���?�X4��9t2dM�R�ށv���`J��M3���D�O����1���Ġ<����p��p�cF]��$ȩb@z���$�O��{�CĦU�I������?��՟`@3*ۀ9D�		��|�&�i������d�O�lv`�O��$�<ͧ��
�"L[`�Y�G��	��y�f7�ۋ@,9o�ןp�I�������ē�?��d�R1���X�5R�`F�!U��&�V+!4�O>���4Bl6����=���x	2NQݦ��I����	0>�ɱK<����?�'� 6�P�⚘�� F�o���Y۴����O��p�
�O
ʓ�?q���?�1Tc�\ S剶�P�d��Ƭm�ԟ� �G����?�������U07x��G�/q��Y�LV}�,D�y�\������<�	ry2kN3n3��2ଐ��D�:&IF�<��|��;����h'�L�����ڠa:k��0�����[�)��b���	�(��Oyb�ΜN
��,nuܨ���6�@,1W �H�꓍?)�����?!�p�5��8n���Th;f�Z�`Z�� ��#P���	ԟ���]y�K-F��<bt �*�.x%\���+�K�զ���A��ğ����5�� �IX�䖚�8�s�#�~:�B�m[�	=�V�'h�_�,P�̻��'�?����r�cHI�E~diw"�9+���4\�(�	��\���Q4F5�Icy�O��)W�)JI���9br�T��ܠ0���R���C��M+bX?��I�?���Ob�SfT���
���7X��4Rýia��'�\�&�'nɧ�O�=hV��"�xL�1*FM�H�aٴZ {g�i�B�'z��O�O��A�"�m���	0I�GNàQ�z�lډP�D���c�)§�?)��	�@�t2!���jy�5"µ2�v�''R�'b�}�֩!���O����� J�C�
	�@qr�Z$U������ie�'�j4y3#�)�Ol���O�ЈDC�I�H<���G8�@㦛�y�	4�& XN<����?�H>��|�����g�� �Gh�Jږ��'�(�6�'��	ڟ8��؟��'�6	��Vl�xk[V��C�d�;v��O��!ړ�?��&ݥD�.t�SÍ<Fö��G�
H�"i���?i���?����4�,�BB�ODE"�(Ay5���fD\A�ZT�w���	��ڟ�IO��ڟ�	((6)���nӎPGں��,p���5�.��W���I���IPy��_��@�	�c@�S��U�����|��P��٦��	y���*j�c��q1��27��9w�ЇDK|4��m�B���O�`�d�XG����'\�4�$��ИC,4Z�8z��	�]��O:�D�O�����~��I�2q �����6.�Uy�L�æm�'�8���j�Z8�O���O��Y�T1r�AةfW
T��(Zyl����
]�#<��7g��q!��#�2zz��aG|�Y�Ď�OL���O��D�����O�ʧ=sP���*|��1�L'K0�����i�����Z����V���.J�v���ǒ�f��܁�ߍ&�t�l�ߟp��џ�p��<���|����?�#ʏ�b����Q�q�J1[��=8��O
�@�,�D�O��D�O��:�ES�{���	�f�(	ݤ�ۗLh}�<0�2�'^�I䟄'�l�č -4:�s��˙c*��Y&�
����Ig0ᨖ����I��X��_y�c� Y��`JEaP�<�^0˖�W�u����c/��Oh���O*��?���!�� ��@5��x��(��n�z�k�,�\̓�?y��?Y+O�x���|g�3~���E��%.j�&��z}��'bb�|�[�h�̣>��&�39��)�>j�T�0�	v}"�'���'L�I-^� %�M|j�g�2&5i1lD:<�������(b����'$�W��	ß�KE�4��Fr���1h22FDP�̝6f��7M�O���?�hɠ��i�O�������o��?*#v(�N+�m����{���Dh����SU�����9F�L}I �ßr7�듷?yŁ�?���?Y���*+O�n�qY��!��ٍ��&��dw����D�� 6����*�%V���� ǆ:��(��i�"����']��'��O��i>Y��x$nɀq�Ž#������C�����OP�F�)��ן\�a�W�/��������K�fM��M����?a��Yt�*O�I�O����8�&L�Lv"�+WÁ����s��B<�O�'>m�	���"d�xQJG�)A���p�?2�8o��X# ��Vy��'�r�'KqO�%�tI������ `�I[�t�!	Vg���?������On��&�
zF<�����@��;�kD&Gݎ��?y��?��2�O���gΡ+��` ��E��@sֵi�1��OJ���O�˓�?9��Ƿ��#�b�Dqz�o�"��3��M���?)����'D��[�|6�'z��;���!c*��y���(~ �	����IcyR�'�Z�At\>�������qr��LoHY�cG�<�,��ݴ�?a�"P���p�8�����ȥ)1_�|uY��`���'��򟈹G�MH�t�'���O0���6�D��&Uc�K�5
�h,�!%��gy�.�	�O��0�x��'�ɞ4i�5B�Σh������K��T�	ڟ����?���u�ьx����]�,/t�A��ޔ����<�t��B���'7����C6	Q�������]c�oZ�c���Iɟ��I���Jy�O��T�v���.A�N��yؤ��h7�ݣ�>�S ��S̟�"U�r�\��Z�lv�{���M���?i��R�`��*O�	�O��$���r��.3˼����#�t�;�$^��O`9$>Nth�A�ǰ;�jh� �;D�m��L��9��i"�!��Q��f2�O�IdL3��ADC�u��p��'�ِ��9&��[������B���z4y�b'M���@ώ#n&�I�*7ZꀰENJ4��Hv��nD��" a�\���Ƀ9h� ��c��j�� y���Qu�L�W��!jШh�	�msV�P4�r�� �⇏jh��5��}6��(��(�(l�Mq�x)P�CjՈm����?qJ��?����������=�V�P�9q̏�,*��]����Ր)bʬx�a�1Dy2�ϙm�^���%�,��'�FR����I�|�P�1{t(�w���B,Fy�hĢ�?��if��yي�È�4A�F��ẇ�l�5ϓ�?q�����44H���^#4�a��A�8��`O��oZ�U.4���H�Q��hp�MQ�R��	ny�NARF7-�O����|ZK)�?��F,�c�� �^4IR�C��?a�.���P�hI�)�܋�b�vX���!Y?!�OeL9T�$<�d���p�rb�`�E
:�����@qeȅ�W,�=Z$����Ԍ�1f�\ؘ����QD2*K�(8Uk�OJ���O<��1��.sVȝ�!�P0n�z蚐L��0
�b����~x�\��Z�n��h�$���X**	���)O|�DzBN�*	vִ�R�A�`Q�5�b`>R�6��O����OΕc�N�`��d�Ob���O��ϡ?��`S�
'r��5Jec�O,��"�� lp�#��Q,cB�qp�&/�Sw�Is�䔹�c�&M���GF� *Ը M TT�����fL| ��$�S覭IBDi�� �<Y��6Fͦ��wK�)��CP%�O�P9(��i>�D{�
V�w\y���()>�=�ן�y�f�$Ok�s��9u��,3����J�����'��ɯ@Fy�2�Z�q����� �]+(�Ҩ�L������I��l�^w���'f�逸L~p��a�4vI��j׮* T�Hp�ڰi2���v�HǓC���k%�B wpUy+W�D়+Q�%a�h�1q��@�r�B�H&O�����G:
�"RdU~�ǊO�s���'qў��?��ƙ�1H�xzg�VR\A d�_�<��F�x4hN��g�� @1f
u����'-�	/,��0�4�?a���D���A�|�H��S�D?"'������?)�HY��?I���?�T&��HU�0��.KRMZB	�SYT�8Q��Xj��B�G�%Q��ƃH�)<V�DyG	7x�e��
�5"�I����w�h��֧ıH��|)�MÌ�dpʤM�V��Fyb�,��I �M�ֹi��A����s���(�J1
�?����?���?	��?!���1z�����F�L�``8��O]<٧�in&-��!R�G����tB��n0��@s�*˓
����i��'��S�w�����Z%:�h ��&������4���	ן,�/4+����c��c@�����9�u�lʼE���w,s��.i���[�v"��'���Hs�>s�@jqD=Sb.��f���H�a�?u�j\,=���R��P�T�7�5}rŚ9�?Y1�i1�"}Z�'w
�`p� �z"daKR-	Jp�']%�!��_͙V*Z�"��Ó>��������%i����aO֮:lt��O�M���?���B��Xxr�� �?����?���5A�n�=Nm�S��4��=��lͦ@����"��� �ش!4D1�e�d�g�O�] �Z�ΐi�e^�}�����0,��L[񦅳��ƶ$q��'Ű$b�F�n[� �!�݄J�&�sP�k�p�o�֟�`'����>��?aum�x&���sM��}+`o���x+�u�@�Չ2PT�G�U<��dT�'�^��1�'u�	 *��@���.G(FDc�m��'\.�H��I���������ϟH^w�"�'��I�7��mHP���T�p@��8� ��q��U3Ng�H��'��@����&:�}B�ʆ#���8sCO�)r4���G�3 1L�Ia�'u2���/S�P�)�Oś[� <��i6�?q��?����ڰ r*�q]⸱�b+!�����F��<y�������#1O,LnZ���',��'�?�r	_�Q�X��c��l�0��ʉ�?���:H����?)�O��й2+�(�,�������Qw♆?ژi�E�ΑL�~�� oJBB�Y0km�'����!�{�>؁3	@}%B9�`�J 
x�C�Z��@�G�Q��̞iQ���֡�Oh���<�R�&U\�9A!!�@)�ppQ�s̓�?!	�s=�=��&ݞU�0� �͂�#*������Í #�x�p��"6,��D44;bX��y�B�3�Mϧ�?!-��e�U��O�1w��3#�L�5V�7�t�x���O���ƵjA�����G4:�8t�ԩ��O��S&!x�`ѩ���RP@��ٶ#���'j*m�C��;Z!�]���1D衙��	H�
�9"��XeV*MQ�(:8�ɀ�M���S�?]8q��Zz����۷cH�Y��Gh<�RC�%�a �P�biD$�:���I��HO�%b�͊�8�^�6�U�a��Rǝ�u�	��������'
�֟�	�X�i�5�$c�"8�^�ȃ��Tt�����{T�-���r�p�$�A+&ER0�O4��N7�J�8�'����:�����>ł���,]A��&ɐ$���� �,��O�.�!���<AuHW1f0��v�A(`)��AH�?��i�bHE,%��Ou�4�'�R�'�r��Tl3dː�$3�yX!c�g��ɒ<�l��3o`�	"��g~�)Q�!ÈR��'j$���1�y��'1����d�|j���T��uy`*@mĦ�c��47�a�Ȅ�0����O����O�q�;�?���tS�s,��(ҋ�J	,�@D�����J�������O1Gk��P�0�$X #QF۔%�F��$J:22��	v����@�5��lZ�
�\6�y��)!Ej�<B�V�Rn@eq�Z<5P��B.@Va�I&�M;���?��?)���?������r�8 ��̶��q��E�P׮����JD�u� ��0�_�7�̠�<i'�inRZ��c�

?�Mc���?!%��9p�DѸ�͏�/P���g����?���9h*̘��?Y�O��m	���"��U��ۥ��8>*���	9k&42�� O^I�A��'�H��".�>����3 `�čҗ|��kҧ�y8���v��OJ,lZ$�M���z����W�RnT<�tj�;$�Ic(Ov��5�)§\8����!bj�S#���NB���#Ǜ���#.�T�w'��5��4P2�_�
8�[�̃CM�~�*���Ɵ �O�� �@�'�v�򰆜=O�vx�"OV�P�r�E�'R�N��$����k��-K�`�=y���w��^>9���	&�U�nD*��qlY���I8�F�Zwe֯hزT�P�9���?�zr�qC֨�%�u��qq�1}",K��?��i]�6��O��?� �x�a"�[�.��6m*���C@��O���w��H��]- �h|RB@O%iax2�-ғl��u�c� 1�Ybb;���iVJ[��?���?��,@�qbAi��?a���?9F���)���$M*|���"5o^xYUf��H&�Ӥ��x_8�* �Kl�b>-'�T�� {n�=�3�նcQ�1�R�+�D��Fۧ���B�f	(���>&��HąR	R��Ѡ�֙m�����i��M�c�i7&�)%���,OZ��Z�+U<t%b����h��
�S��C�	$�=#�g��w���Ġ�X
����{'��۟Ȗ'1�U�Q��-���s�Ђ���TG5X���'�2�'e2�a���	��	�e��[ǋ�,a�8�֎��W`R���KO�O� HT)�X�B�o��� 0 �'��	B�b�'J��XJ�	;#^�yCk�9D^��z�CE���xE|R'ċ4�"(��ʅ�S�y�F6�d)	���شՉ'�B�'1�O�Ę�	��c�R�RC^(��C$��O��D�O����&U^@���<�@��#I��2�O��n���Ms��4��� ��CV�ͲqK^�Oh�	%"O�P��� x���ʋ�J� -�"O}k�ɉ"[�TM�&�lBr"O8e:Gd�%m��`l@�L��7"O��&�){n ��4��?rpCC"O�)Hta�
,^�1�h��\]P�)�"OR$C!���2\#B�X�k4��x�"Oz`��˻Yp��ǪS���щ"O	���d�Б"&�&j@=�W"Ovi*"�!2*©��H�2\bŘ�"O� 9c�#Kn.Q�ƅ��̳`"O�)����c�!)�K�=��M��"O��qrO����h0��P��`yE"O�A0��C�+�j�R.XY��[W"O!{�c��F���q�Ɛ��Va�"O�$�0���@�"�D^
52���`"O��[3[2x�������bH���@"O���Q&+��Y��&vB@�aA"O��2 UtK��
	ȐLP�"Olpp�ƥT��b
N6���I"O�0ՉFT&-	u�ڷrJ����"O,��Ql�(a:̈�e ��A1�"OV���j�,;�)i��ˡ8�Y'"O�\"6F�.[��2E��Z��@%"Onc�*Rp���R�)G�����"O`Q#e�5���CCNK�I��"O�싴̞j}��� �_�c�$Z�"O�`���-��a�R������"Or���8.���ig�� T��	�"O�����J6Ms�Yp�f�;{��d�A"Oxq�3:ȖXd��H��P"OP�3˥ ޲Ճ��Q/�����"Oޤ�&��f?�	{�K(���"O��;k�TXѵ �*-@�` "O؍`��gpj	$� -0[�	�"Ov9�k^�4��7��I �� �OB��3E�i�vI ӓ0<v���²E}B�§͋�yjtч�	-�$�Q��N8^;Z���n�6㸠kӂ�#3a��s�Mh<�r�Dtdp
F���G�T9���}�''��s�B�jh�=��Rx��O�M5b�i�'JJ�97�ʃ�аh�!��ָ��`G�/�����B�><x1�d��N������O�	������T>��]P�����Q&�赅@;@;�B䉍'9(k�i">����P�S�;[��z��"�ɽmI�iHc��%�Br�3(�� '@�� ���IC$Ӆk���I:b.]�bH�9T~p풓�E�B�:�që��Gr�,j�L�.y�^�*��8w<*�x �߂&L�D�L^�
]p�@E"~ԕ�G�\8�Oh�	��N<�Vf�
@g��6|x�Ic=OT�PSFS� F���Q��䂥��D�����t"r�au��!����7�4#�J�H#*<G��Fa�<� iq���0�b��'�����yw��3;�1�`U�sJ��������y��3t
���j�6.�ʥ���QPcl#����$�;��'Ed�QA�O�A��g�� �Y�%����.px��!"�;D�'UC`��No��в�gR����.��yW�O#L�2�(T����L��Ba�A��~�B�7EP �0�Oq*�b��j���q/�&��x���$�:/��uh��ݭk\��C�Oq���)^�BӒ� �(H3^�Pa��C?X>>!u�O����u?� �ā$�%N~�'����?[�N���,G�d��� qB���!��*.Fb�	i]-		 �Q��*N���T>�'���vNR�<A�*�@�',g$�� rFB�|��  �z��H�r����|y��AL�c^1� ��+��I��۳
�%�'DL8�O�$y��1H�EC�A�+��,k�Y<<�de�	�wH����#Z,FN��Ӄ遏FT��q�*6	ɴh�@�/9�*�m?S!r@�O �Q��p?��D�~�4���'7��(A��F9qa���-oH�Dx�	]���S� or)�Ɗŝ��$��Q�Z����J�C�U���U�,��V�m�Z��'	��ȣj��֘���,#X�x@歕5.8m���,1;:�0�m�'$^ZXᆫ������T>���$��+��e�x�Q��(~`�I:*1�yZ2�G:U߀���IC���b`*�M\pe��q=��3 �)�ɘ^��)#Qt!j����^`�]�eф7
�!�7C����������H� �JO(6�@�.^	I<�"�����E�FiS+k┒`ȃ�~ʟ剞R�4��ӯ3!���T�ڿc*(�� �5�ģ<Y�Ȅs����P�ʟ#�*)��(Ey��2�X�bm  18�F[d.�`V��D	�<酣�O��?�a�Y�{�>�[�̕0h���q�Vn��j����Yv�T���S�5J\aM~�Y��W�dHfB��'���˔ �X���㉼\�I�7��*t��|:Eᓎ+*4�����4:�ک@��߇�>踦J3�s�ʧbA�D�`W�n�tmۀ��|0,*�:����J�4�H�abƍ���-��,�eKW��8f��YA����d�/}��I\:)g���W��'ڪ!�2F�3zaz��,-U�H'�9}b�H;���G��" �'�l��AA����'�()S�$�Y(xLP$�pؐI����+\N�䀅=��x�D4��+w�����4 @z��Y �O���$�\y��y�d�V=^��e"E�R�t�C"�j��1�H�p<�e
�P�0����5�^�;5l�8&�ma�9�Y��'T$% UK���A����B�2ВEMBb��$ 1�S�+����j�v�e�``H���=iC�AO���*5�C�kQ�]�T��\8�2a�|�P�pϓ?�\9�6i�<AP�r��.u�d�N�u���p�.�4,���}�+#����9z��H���Ś�ē14)Y6�ؿ%ή�8a�ڷZ
>�Dz�ץX�-�W��2'�J��f�K��$»/v*�t��C�\�`&��9c�"��f�R���<3��%|OԹ2Bf� N�Y�d,�I'n-eF�c�ֱ
欉�F����w�f,ie!%lx<�U툲DJ���'wf-k��B�8:D��a�<[�|̱F��p<�KX�]rl$�5�$X���T-���Mh��3i�X���E�=�J���I���J��R,�"�Q����㋟7v�����k�
@��	k��sV�*��	SV�|����5<���?�'BX��Zl���2�r�r~�%��_��"4%}D	I�C��O��Ӧ��n�̉ @�ϪL0�q�-�0��r(@$������B�Pq�O�0��B����YU"�.U��%	w��yGDB�R%9ŠPe������ �xBLR6?z�8w�V+lvir��A�]���pOT )�B�&=���*��
8������2U�J��A_�*"����W!\~��I�e�����(�a��ҡ�PL�$eYI@���?�slІ@[��ZfN��E��IZ/ݦ�`��K�(S��	�ढU����~bB�����[��\��Թ�6 ݚ7�PI�Lq�<�q��bu���lX+ڶX�Rğ�^Gn�"P˂o?ѴQ��;_w��x	2��*-۬@+��a���`��^��	#�OpV�ĘDA �O�)�5���~~-���R�fwD�)e��9��d��@a}"�F9[6�b@/=f"��f�U�{�h��?YR��-.��m���N�A���c�E�'�.-�S�5 O&�����B��ـ7�۠>l�k�!�X�Hc�!@�#$��JD��V��m�1W�#��GZfX��lRXm
Ԗ�t�ȳy�F &*J�3R���B��M{2G��FLTd��N�W�X�e㛣;��i�@M�<�i1u�Dt~.���K�RT�`ƱA�Y�-�|Wș�� U��? &	�X�s���}R�ǎ_C
Qp�o�\���)fbI��hͺ��	S�vp�׮�f.�aF1^�~+D�͟yTb�hC������GV���Y7D؀.��,;Q#E�x�c�ؾ5Ä���T�T�x��ц*q��t[����H+|�QDĭ^��S��N�1 �i�4��������N5��Ok�\��@Ϳz����^/�$��&��:$`��d4�eDz�%��9�^d�f	J�M� �C�M ~�Yڡ퍁��ʦ�@��TUz�BM8&�d8�����y�NT��ԅa6A��;���P�DeTT$?y	���.� �;��73��hJ��h�0����
�2���⮅;	A5����Y�,`+q$�J�Ӑ$Q1���K�kjv���k�<y��p-6M?���n�O�<��N_�a%>c��X����V����H�:$]�=�V���QA����a�)8ń�PAˡ(m��Z��������QH�8 U����u��\�L��-����1h|��Ɋ %����2)h�G�E�d���.2� ���q�\.P�����mBw�(�Xm^���Bj�*KV��p��Z�EP���S�.O�D��x2x"p�Ċ4c������0%p#=)��B�,0��jT�u�p��M	�V0>�`�͊/:< (a�[& ���Y {|,8��`yb�[|y��R�N�a
�����ϒ3O:���s���o��,B���)�V(��i��qp�Ϸ���0�M�(a��$;q�%%j\Z��O��R�M������M����xD�ɵK	��c���<I3�=fW.$:s���v�h�`��R�'TP�;W*γ\�"4Ҋ;$q�����7-���)K�������*]�P�9S"Γ�uWdI)�䩛�u� ���5L��u�4�+tlH0��]��C�iFҦ��aI,��ZH�cìڑ_�x|���p�xa+%�E?2ĺ=�Q��5y�`ŏ��y������?IcU��ԭ�w��U��h�c�M��HO��j�8bF���ǈ�$��`.��^���0	�/Y�+�ĨU��	 ���=OP����K�{F��O�� U�?�q֍�I��b7l]!
��9��� �蔒`�~ӆ�)@I�#^�5C`���|�q@fɘ�D�p`E��
�+!�F��۲�Y�!�"�K��,>���+�	��)���L�����ڴ��@��=O��(Ρ�h˴$���4�Ԕ1������8��l�/P(M+^l[���]�Π��~�j��<�;\���+7��l�2TxaŐ� zh�!�^�6����b%3���A�%=��ي��@�F-r� &��/m�z(!'D��\�4)T"d���<E����~q+�#��bQdE��
"Rv"=ѴK�(7�4��BX�l:�\�	 I�d�B�C̜&�X!U(²bE���g��,SayB�@�%E�Y1� *٦���L@H	�T-1�0(�CMzC,6�	!�Db��$!�H��g��z�:�P��J&"�X���6jt�Y꧸�)rg넽KĄ���\��BD p�xɋ�����D�^nl����	#�85�D���O� Z1Iړ*٠�ՀB1
,�88qD����X84��y��>A�f��g&��P��^<�$�3�&�zb
^/E��?y�l�'F �٤�#
�T9�5CՁ4v��9ѫ�E�L�I�\;D=�G��=�Z��T>q���ȏ����m�.��5�7���HO�Yqg�֧!�DA��T�o
�Y�D�s�~]�f�X?�8����T��G�G�-֎�d8��Wֺ�G����K�*q~(�'���h�었ec�r#�A�^�(mm7Y��P5d �JS��)� P�U��QK�!�S�0=<P�	c��9VB�n 8�(7,�3��3�b�#����_� �l)&$�v��ݑs(F:�脺��ݴfJR (���=r���O�_��mϧr}�����~w�^&|T�8'
L�.
�ce�ڡ��>q��P��~� �z3�!��aK?`�
 y���4~;��'aJ=dn����'�?��
 >���A�閊��I��Ҭ3�a�)MWh���Q-)ێ"=�r,ƥ%��8�4兄o<\`����)�r|���Y#V��� >,X��[2jL������}�� ���ӢE~���'n��k����_S�yj$��2<Stܴ3->ucto��J	�yyS�R#U?����%�����պ�6��YFc���;Q@`EK��_��0�aF_h�F�4|�d�2�5�*��Yr���6�x!����3�,��#�c��L#a� 	�n���9j9�Xp�:������$�w���F*T�48yd��MJ�{�Fٯ��<yl��	��19� ��h��d�4{)�Y-e^=���ox��32h��߼���OqOh�{��OȾ@�u�h�܁ClQ;36*|bQ�"ғr���xk-���c2��;_�.�j�	�S�Μp��1P� w@�{"�mC��'nz0�<A���)��Q(0�T=�#
�V}��V�Ba!��H�Q���녚�M��Ch 1��>F7f���o$ ��F ��"�c�+u���;4�\���%���(rFD�9�qDk�%H(����5CNK��� �ԙ�r�N0LA�앓0R
@pI��*_�%��&u�N��<��'��U+�i��Cq���U�Z1iya}"�T�"Z�=P6b�8�J��3'،L�ޝp�!.!)���G���~{��T��B��Z��K�+B�3�Lq�OT�Q��G�A���[�uZ�i�IP*ΩꃄO�cy�Hx���C���O�$���B8+���ҴnӰ���PD2?��a͖�����^(�Dd�1G�W"ց�E4�M��l��c�B�`����.����)���"����r�$�8D5)!�`3�"OFAzW��V�He	��R8jx�8�4e�7�j�j)O��s��t��D�`�(�%�|[�NE�=cX%�1���Eʁq�e7D���1��
]��d"�nI�S����(D�@�v�١m��`���6�NG"&D�L�!J�,@�)���F�W<���&D���W�ޙ�Vub��Y䘚Pl)D���	�'o�`g�I�ك¤%D� �N%<�|D�
�0n��ջvH'D�4�ዂ�
�t���c[�Lh��#D�La&�Z�LU���q�D�t: �:ǧ D�����x0͛��B�M�H��?D�8{�+����*D B+US���¤;D��� P;R1��H^xT|@��J8D��)�N���Ļ䆖���(��6D�P���
a�P��Ԃr��!�N5D�|����,��Y�"��=�����y�%]�̙���,BE�X��FT��y
� ��ɗʨzyL�2�)��Mj���"O�!{Vc� "�]Z�Ŀ^Q�sw"O��/в4AX��̌�7^�2"O�������T е�У%�\@
�'�������kn�bR'0Pl,��'�R��Մ��:O�S��F|���'6�×F�0����O;J��i�'�x	ʄ*տq�&�i7ˋ&A�&���'�������&E��Pׂ�3��9�'2���C� <g-�iID��:y4�=�	�'vʀ�ĉB���� $lJ'���*	�'o�4;���<q�~�⃎�?���!	�'�ȈQA�ʙ�F�03͘.2�� 	�'a�``=7�L��f�"�B��':��7
�l�h��t�E���	�'��IإNyH�Y�P�ę"	�'�1��O2r�x1��Z���a3�'�P|s+�0dT�|���5�ly�'�"��v��ߐXh�F��#��b�'�x�z��N�9in��0� #`N���'Ab��f�|�����96���"Oi����	��=��ӮZ����"O6���8��г���
Pz>��c"O� ���s�P�d�I
�b��"OP�#�*�0��$�0��ȶ"Oε'��(�a9c�� &��h��"O� v��8_8QG� �n��"O�&�D�8��rW��F0�Q"O�\�� �t���Y�B����"O�!�
�>y�1e��<J2Ug"O�-���D�F���_5{1lUJ�"O�xKףQ�c�2���6C�Ҭ�#"O�U���ܸau�Y�G��?S�6��W"ONm(G�vh8�h�N���4"O2���B6M|�����7O�jhq�"On]K�.G��qhsኝ}���JC"O0e �n��~a�1��NQ'X�*Ⱥ"O�0z��Y�d�����{��b"O	�jZ4$���UowҡZ�"O��c��1���B�)~�tL:F"O��3ժݰ%�����]JBE�'"O}b��<J0�I�5���^D:��2"Oؤ�gN�tb��`U�N�W!�a�"O4h�Vm@1r���K'B��##��"O�:��4n@j踢 �B
�)"OB����?(��8�/�|�D��&"OXb��:*��Tk⭒�/n��+�"OР�.*|g8����[3���5"ODe�a�8g��\1�"]���(�"O��:�
�=c2����x��H2D"O���2�K�o��@�� 8�ָ�"O:Ys'̆�l������a!� t"OȐQ�@�Y�¬��=:Q�*O�1�O�$F)`����2Ht�+�'o$m��/��)���� ]4FrE��I�Q��8��|� �H:h����/pE��oJ
X(`��>B\ ��ȓ���1"�KrhuꞼif��ȓ�����$�=U������5)l���ȓ%�<D�s�������BY�N������kc�>E�lʓ�Ny�T���uOq)5c�� ��l�Ԏ��p���ȓ^�ܩ���Q���2��<H��y�ȓko"X�%`ݝv���@�?Ee��S�? ��`�W�'�r�3R�G-qz�K2"O�lr��΁G\���6��&a�H��"O�t*�f�V@��x��̵U�ȣ7"OR���`S9M@v��"'uL�I ���ax�	ċ��(�Hޤ<����a�9�y�OƝl͂F�:����'B��yBɸ^��16C�,,��hs�M#��O����O=�%Q�2�X@ؑ��!݀�{�'��]�p���i*)p1	�h6`�'A���E@��L1 e��Q�����'(��`��7J����Å�Eʬ��'L4㖣�B��sbcܨ2��

�'e��� �NF�i��-8#�i�';�U)���m�d b����2:�0��'�Rx��_+.Nh���Ȼ+�x��'������0} �R��D� pI�'Q�E!���%M�.� �jL������'��t�Rl�=K0�0�K�tw��ܴ�hO?7�H�F��Ȑg�48��ƭ�yu!�$�@����5yHЪA-�
�!�h9>z��  g1�x%�09�!��'o"�eYT��ID!Ԧ.!�$�&�� �ڡT�N��g�?�!�]�Z���kP���|Sk�j�!�$�d�(Y�F�m)�-Ȕ��_1!񤗼J�&)�&l��tҔ��Ń�%��A�'�X�0# �Z��}�VAg� �'�x����X�`��Ѷꁻ!6����'��@`�U�0q����(�ⶭ��'�`Q)OR�G����u��q�!�ʓYDV��"VG"���:/iĘ��aȁ���%x@b"�Գ�ʐ��IM�0b3�I1%_fE*u�&�Y�O#vC�ɻ]'�Q9d�]����@ҼI`�C�IM#a����2jŸznC�	$:�,�Xd��m��X���ËW)�B�I�2�p�iU<3x<�k��a�B�#�p�ِ�U�L������i�B�	�S(l�2��Û	���S�m%�v��d9񤄦S��|J��w�p\���=!�d�:0�� �=����`Ç><!�Č79v�Pp���L�����<{Q!�dY�)��`#]�R������y\ROn�B`ַXq��:f�)e& p7"Od��mA��
l���&o��s�"O CҎҜG�B-1T�L9Lϴ�p�"O�0#��
4ц�(�CN�8�А�R"Ozd����Xq�����
p�g"O���&\�d�8�%�
'w�0YZ�"O��
�	�>�h䢐�	� #�'�t�f-}E����F��u;r�c���{ y!j�"_�^���ȓ^D�h0���j�|���N,��m�ȓ	R���1`DZ��A�O0*�ȓ2#�P�čũZ�jȑ3*؁}�F1�ȓz�b��@�&
�Myㆻcra��6��ѷ��x���T���لȓa=
d���L�����*]Z��ȓM�	cDI)^���"0��E�ȓC�d	�4��XP�=�v�V���-P��J�"�c�D y�G� )��?��]�D.���f�-���ȓz,�J�&gf��.�n,������A;6��6t�tғJ8��ŦO��� ����mL�Dde� ��ZP%��"O��W�8F�6M�'�'O��Y�"O��J# �3H�̢3�
,U�]�"OfMQs�
�dx��)'�_�Z�`D��"O�30!K�v�2 � P� A�"O��S��	B��Ж@�R���"O�X�MHD1�	x��п5�Le�"O� ���A�(o�Đ�O�1�f�KF"O�(��c��c.ӱ[�,��r"O����`�<H��Ia�
V�&�R'"O��H&��$=�N]@B�*9
�ء2"O���Tu�N�a )gMj`z	�'&��ŮP yR�tR�GMT/8u	�'d��C�"\��	V W�O� ���4�hO?7-Ūz:F���N�����F�h�!��A����@%J����+!�D�:���k�'�7|�X��Ņ�Q&!�Z;S��]���ӲS��s�M�I�!򄄬��Gm����� D�!�$D�fm#�I�3�4��� P�)�!�6
�������@�F�A�!@2O�!���6Ε)B�C(b���B��.�!��R�1��D�V	1p�Aa�O�Ce!�D jG�1Y��9@�X	g�N�P!�D>9�ʜc2�Ӭ(�t��&ՙw�!��K,~��E�$ J\;j���$r�hC��6�j<�,�nd����&K�RC䉧7d8i��9&�I��T�
U>C䉲���x�Iw��Q���γ`��d'9?ZI�P��T�:As6�G�8��9��´��GE�I�I���0�"-�ȓ0�V��0*M�.�$��L�X���T�
�3�CL:�Y(�-ØHȢ���KJ�z��	W�i�*Qy.ⱄ�d i{��6�x}�R��#J��ȓ2�IBR�Bu
�����H捄�3�~a��#H����4� �; 9�ȓ3��Œ�o�,p*��U�:O�h��	j~�
�0�Ҥ��ՕL�q��(T�yB��I���jw��B�ƁsEł�hOR�ۍ��^�*�|�p�.�9xK@|*��
#e�!�D׉���	5�	zJH�Y�#L(x�!�$�	>�=A"�<Nז�ۄ�i�!��BY�ˇ,G'2ò��hɔ=�!�d 	��̓Ѣ��dE�i��ٹD�!�$��d���ݙB�(����!�$��2��eCD�u����C�r�!�F!�b�+���=BV�8���J�!�NtԌ�DA�#Hy�T��P�!�̬wԂ0��@۽94�P@�=�!�$�*� qᬋ,Z�2-H՞�!�$�(]<|�"��Gk��i���*�!�$WUz$�x3H��u�YɁ��=�!�ٝy}�DP����N�C�KN-�!�&1��yc祘m��Pp�/��<!�d ������;R�@m�$�K�m�!��ŸD�tEL�;�6`��ҰZ�!�$�5{s��x�-�U��) �I��!�D�ޜ�ZCoX ��E�u)?:x!�"jX����N� p��@�X�i�!�'�R�8˓��V��b��!�ͼ_c��r�EJjmc���'0�!�dR([���H���WRd4{��ǺI0!��ڨ(9hq B�;|@b�rw��"!�� >-��;,���3��E*~��
"O ����[J;բ@V|Νµ"O���R;p� B��sdh��#"Op�4A�ʹ�`H[� ��%"O�9��i^�H$�G)A�x���"O�8K�'�Q�咆Q=��0�t"O��1�L���rIB�*�z�����"Oh����H�Ӑ	Ї��y��!�g"O�5ɢڧM'�	�ţ) �x8�p"O�U�3�K���t���R%(��pP"O��$$���d�����M��4x�"O|�H���Sk���cHV��$4"Oh9H��M ���1��S��Di�"O��DB�VR����W5���P"O:d�aj׀}�4��'`T7���"O�e�ޤj�6�aEɊ�p�dQG"OB|+"��:���:V�F
q�!�Q"On!���6%��%A�$?�y!"O�p�)՘PG�����']&X�a"O��'FQ�N~��׬�<#V0�B`"O&}	��[���x�� ,Q��(3"O�������=~2�#�(\�c2�uQ�"Oꘛ�@��k�@��4�	p�L��"OB��&��	)�e�vl�+nε�!"O��sFL�70w�m��GORbTI�"O:�{aB�(8�^Ё�g4P�"�C@"O~���aM
q���� Ǿ;��]��"O��ǫ�qV�l2ī�Vq�RA"O܅����q��Pp�G�`\|U��"O��( kZ({�Z(I"�
)OBt��W"O(�HS�Vv�rB�ţ
�:D��"O���*�{,,ad+�Z�TY�"O<!�t�C�f�偂� ����"OxUX��:��!��1
�t���"O�9 ��7�Iz��1��DZ�"O�@�baQ*l0�=�v�ݕyL���"O�ő�,�}�V�xSϬN6����"O<h:�@C��tl8u(�1;Q�{�"Oh�q�KY?q��H(�,��a"O��[�"�'cLʐbl�y�[""OƀB"��#{�n�����Д�/�y�/P,f�~��PH&t)c3`�;�y"�G$4r���C��8�~ը��_�y�Q�Et�a{�h.(�m�I���y�KǀP�:��êI�n��I�����y�
�N{��@Դu����ǋF�yB�ׂSA���ؔi�ڝ�g���ybR>+�*̑6d�8�h!�̒�!���48��]�נ��bL��s#�X�!��l����AI�yx��r��Q�!�d�<T���x���NM�}y�/O ?�!�dF3	l�%��(U3�`e��#�!�D׌oѸ�XhX�,X��4�9:w!�dU�fR� ��T�6+ �R���!�D��lH$ �O P*R�Z�d!�ݤӀ��83��P��F�i!򄋳����aÀ8��h��{!�DƜu�=�A
����]#h�#!�DB�7ґڒJ�A�
��D&� !�$�2tF����FY7�.|��n@7P!�̭�h��N����o�{�fC䉐g?�0��.'x�b���OXZC��;�BT�w��Z^(��EY�^��C��2D�4�*�Ͱ �&��B*G�C�)� ��O��3bR��6�}���"O�Ȃ�Aթ�lp��G�]z���"O�1�KD�tՔ���G�Vװ�#�"O��؆���m�t�*tJ�?[�!ӧ"OD�)��\@S����cP6\�ر�#"O09i��[ؘ�7%ɪqTf�KV"O@��GT�c:�x�Ɇ?\���s�"O���&ѿ(�]��G;/��!��"Od�񕤓�Ziug��!���;P"O�)�#/��H����цԒn{�є"O�aQ%h �J'f�#F6�[G"O$�3V���pkp��v�ϏM[J�"O��࠘�M�l�Sd���xydI"�"O�Ix�+�V��H�){~+"OH-��P$9ǜ�s`J<[�
ɑ�"O(��%B�:_��I!��]:�$9H�"O������5#h�[���?߆E�c"O\��N~��d����M�}�!�$��E/6�H�E� q�P�́4�!��63��8�gʔHg�I��/i!��r�xI�!�R�JJp=2�j#6`!�ĕ�$��	�	F����J/@�!򤛳qh�H��(ȭe���y��؀8!�H=u�l�{�� �0�%�E�8�!��Ô-`�H��.R. ޠ�q�$�?JT!���56������rG�=@!�D�%���Ce���š`!��� ��!�m !C�M��!���Fd��h"R��0T��!���|a����xz�U�G�=|�!�հH*8�pㆎ�o�����\d�!�䓪�4�g�Z�D-m�!�K� �<ĸ'̋h���3�����!򤚧RdGV�{�x0���!��S"BX��*���9��A�E
�g�!�Αpk^9Ѣ�o2,Q��Ȍ�<|!򤖼N�`XT�**J���G��b!�D�;XhLI6����0#����0!�D���(��3o���E&�?x�!���lQ���	{~��YS�?Z�!��:V����f��7L��Jͻ9!�U�m���q�FB ��W��`!�d="$��@��3 Q�6��-~!�D?8_&�
E���Vy��i��L�(s!�L �p)Ӓ$�h����%�
b!�d�
*��#c�$pa	�`G޴VB!�d˦U��,(�͖ �r���7%&!�$�+D��8�so�>�j ���,*�!�/=��9��5�H�XT�WZ�!���$U�~-
`�+W�P}hm�1\!��E,IVu�Ŕ(#�����_9E!���D)&�c�dN���<Hg�H�+M!�đW�4�GaA�+���v���O8!�Dɻ*F�1��"�h(`ū"F�!��-+�x; �J�w�L �2`_�!�DD{�$1��.��  �2,M!�՛VP�89UL	�=�`M$M�!��اOs��邩Ҟ#N�a�#G�-�!��1�1E�^3Q������3�!��Z#!��gi��KОA���E;�!�օU�)��"7n���Kw":�!��;�$����	7]�����ʂ"OĜ� E�nF�`�f�%�Tr4"O�E�r�3C�`HtOL&V*J�b�"O� |M�f����N}K�-c�@��"O"�C�-� ��{tl��ޜ���"O�8� �Şb���:&�P!q|�ò"O�q9��=��(��È��P"O��VO�N[����A��B��u@�"O��h��P�j}׀�����"O~!R�`���/�_�֐��"O�-{���$ Sr�Ǝ��s$�)�$"O�܁�H&�N���T�. LJ�"O����V4�>�mC:)�UZ�"O���"��:id��i�7x��C"O�H�g�bK`
�n�W����"O49���?6�`鑎�)9�2d��"O��S�RTr�cҴT�q�g"O�-b���U�*�p���5Ԑ5"O6%�͗�t��< �B�|S��;"O4͙ŀ��(�ȝ2��лO�RyzS"O֕�r��� E�e�
=��%8"OЀ�$��L�h9A�dU:[t���@"Ot�3A�ɇjڍ�pn�M�� `"O��#F��`�O? ��"O֥�u(U��B,P�"D�r"O�U�g���A�H����W����2"O�AY ��`���ơ:G��q�"O�)�# Y��I��N�9:�<��"O��*1��}b$�1�ᝬi1N�k�"O�qs���4o$���n\�?�Ȱ"b"O���'N�)bVQ;��* ��1�S"OF(�F+�,U|����=���`"O`�S��ڛzz�����	$��t"O��	��p!��k��"[�bx�Q"O���t�Ӫw�&\��a�̝�"O��Xc�ox}�t���$�f�`u"OH�����������#Zˎ$R""O���&(H6u�>mc���;��#"Oi"w��=n��
 �#7����W"O ��c��8�<�I�����"ON�����;a����-^*<��I3�"Of	��ܓBd��-������"OL�c�`%jI@�b,N&���"O�0R�h�;̚Yq�kCg��0"O��	��G��+t@F,|��Q�"O�-�b��l���07"Q#��T(�"O<�+�Kǥ(��ɣ�S�if��"O���E��(%�vKw�`2�"O�p8�y��mJ��_�-HT���"O�$��N% \V���D��6D�(zV"O��s ��r������b�Y""O�1C��Z//��d���[L����"O��)��$�@��s��~;�}�$"O��(�U�k�����˭?��-��"O*�@D�	�?����)g}v3""OP�P&�%Ȇ��@��6
oB�ҳ"O���ʔ�B-�dK�=QV��u"O ܠE%��#�L9����y7�Y�S"O�t#�*�e��l�#Bڈ	�f�k�"O@�D�/t��@�NA�6�t�C�"Ob��5曕|]n�
�b�u�Q��"O�lH5C�"���#��%� �z�"Oi�-خR�
p˂
�$i{�ܳ�"O⑲��æx���+�BW)�"O��(
qz�03 j֏V��a�"O��r�����=�T� �*���"Oa[�gW�E�  tGW�@�!e"O� ���Ue�Z�(x�fA�I�h��'"O�`���K�|
0I�dQ=&:^��2"O�8��`��,���HFb7=��y�"Oy����O�C�AҜa��Xa "O�횑i�:��2ugZ!l�"A�f"Ol�k����v,�v�1 ��C"O@I���\P�XPŀ�'�p���"OR���`�)Ć���D!]KP)P�"O�,	aȀ�y��8(�A�A,��K�"O�,�]�cs���u����%"O���V�� +���׉F�Dzl���"O����a�7Ϩ���)xO�:n��ȓ$8:���X!�&�Z��ߔ����ȓ'��� ��(8�$
EF��d�p��1�����Y�޸\�Lf� ���^e0�(էH$�	�T#I����Vo�1UB�9��I�f�ىfI����9�D]"d��2|��#��[	|��H��oiN�C�_�X<�WǄ	Q*��ȓK'L��LV��P8�g���k,D��ȓ?&`�[RC�d�M8��d�j`�ȓYd�iRլ=o�Eh&��j� `�ȓipp�1����[VO�p��%�ȓf�f��@-���{S�֍PA�݇�Qq4{T�E8̠�0�_7ŌL�ȓ�v��AꇔcȄ���	�h�ȓ}^�K�_��9sG	 Up�ȓa�.��ҮR�xHl�8�AV�0�VY��;�A ���.ޒ����È���=G��tC�@4�[dgą8���^��(3p�Ϫ!"�̓\}X���ȓx같�0M�@�a[�%ƄfWX��ȓCe� �p�yv��F*�U沵�ȓ-ݐ�ʦk�>f,��Y�t��$��'u���c��:\��aǩ;�舅ȓPv��ӌ���Ȩ����Kbd��ȓ�x"�N�&"/��Ɔ	�UhD�ȓl0�����T�m���a�]�<��|��^�&�am^!a��!��d� �ȓ�^��G���b��*'0q�ȓ*�ؑ��+I�*:�f�Z����"9��2O�" G<��c��$-�@8�ȓo�bT�T�3>����0�_�h��8��La�M���H9~\�����%_�D��U~�0"�
h'vt�%IY�4`����s��AI���y�.@��$�6±��
�D1��]>C4E*�+@�u���M�j��r�ÒJ`����	���⠄ȓl�!㵊�1W���a��S9yQ�A�ȓoQ���! ��Oޜy�K^�m�ȓo�Q��� @���(cFAS9 ���T0ʩ���E�Y��%���,����["�UX#�;6 ��3rG�(F�B�	3W.$:D�3LR�d�aS�l��B�	�g�=�d�$P���j�eR�u�nB�	G��	�vL*.�5���#@�`B�IF�
���i�c��x��D���B�
vQ�w���:���rU��.�8B�I�(dP��R�,��Џ��&B��Z	7ɛ�^k 4�B,rs B�I�9Ά�I�n3m�0\3�eM_��C�	.��q�K�-xfi;$��0T�C��$}�% �Gۜb<Ze�℁3�xB�	.2e�:���J�Ђ�#@7XB�)� Q%�ӱ�h8y��#4��Y"OСʀ`���|h����G֞t�B"Ozܰ���]9��sQM���h�6"OM���2n�����
1h�2DK�"O��8eʖd���#�)�.��A"Ox����! ��(�KW�Uyt�,�!�䂒
�Ld���=���Yqaɘb!�D2;7<d�1n�C�q9�/ZP!�d]?lј�B�͚�},	� �2X�!�D"PC��Ê��)R�~�!�dɾL	q����l�vt�"�ާ:!�$�&���P�*��`i�d�!������7�؊^lak��C<"!��uخz�n�~E�)Q���*
!�U���1��+09ȤR1.G+�!��ݖ<��È�[$d�RE��i�!�D���������b��P7�!��Z7i��������< �,��!�d_?D)��3�$':�d��l'3�!�d��$΂X�G��>p"��ská~�!�d
	�HEd $Jĩ��-�!�d��e �P�W��!H�D4�Ԋ�*�!����ڠɃi����!���6+!�D�[`����89oD J�	�!�$��l�n���4]��4�&ϒ�x!�@�I]���B��k���oV�2!�d�b�fP�@L�z��3ŚJ�!�OB��٢V�ݧY���GkJs�!�[�T&|-��&}a�S0N�r�S�"O����]�T�q�)T�Y�.�S"O �"�ҘN�5�)�D�P��B"O`��;'`^R�iV]P
�+f"O伉Уk\ ��G�'���"O�1�c�� ����BN��Y�p�7"O�AG�O5X�QC,ֳ�����"O��#45�<丠���A+�"O��i_�;Tp�a�['(����"O�:Va��&��F��
�j���"O֬����j~Z����2nu,�b�"Ojի������������0"O���� �^#,q��Oºlfq�"O��BU�r�}�ƍB�\�P�q"O<�C���x��4�F��)>"!�q"O�+N�Đ�ܫ_�T���"OR���mG�n !`"-$:�2a��"O�8Zɔ>i�҄,�4ޮ���"O���fZ1). H!j� hd\�b"OV�:�P�ri <H�#��X�4DZr"O����MR�u�NE���łh���"O���tNC,/�`u`��d�^��U"O��{Q�%..��:A�R��f�<Y�����P�g��5W�P�VO_�<���%z�Z���0@�R9�T��t�<�w��?�:�)���$��Im�<�@`'xY�K=>��#�
�]�<I�V�t$`��]~,��wo�V�<	E-Ї~��h���4$���U�<�cĖ�y����W0[�(�)FN�<A�G�%��՛�-�g 2�D�<�w�֦qt�͉6,R8>��e+D
Yd�<�Ň�d���� �%Ԍ��#��e�<ip�X�h�@0
�h�}Yr1��͚]�<!O�54�$i`B�A�!"DLp��`�<yb��F=ܸ2��١�:Q��aF�<� �a����	��P!���D��4�"O^5�7j_�h��ԯ�
���`"O�m�
_*l�漪��RA�*P��"OnT�&��T��Yt��,}�,؃"O☡J.2��(�W�\7sh.�"p"O�p�.D65�v�x���( 5��"O��Fa�@jd��Cd��m:�X��"O���f���C���> R���"O�ݠ����#q*�H��2k����"O
����63~A�ݐ8�T%�$"O���!��<g�
ݣ�'�+Dr��p"O�ph��<u��hy�%�GqL 7"Or*&dA�\ʅ�BE��I�,ҵ"O@��&>ST�ETD��BF�M��"O"��a���w�'D�4~D��)�"O�-pt@[�GNPLSBLE�@R�h��"OPjC���e ����I��@�Y�"OT`���OJh��3�F�\�ub�"O�\����3�%�LU���`b"ODYJ�c(=�N�b��Y>���"O�=�qŔ-�jh�7��q��+v"O�h��ԍe �TS��t�t"O�+���,jFMP�I���"O���G�׊@�BX��x����"Od��(�R��E�E�FJ>�b�"O ��U�S�<
�)�C�]�p*�"O2!"L�L�� E��1p�F��"O���1B���-��Iw�[�"OX�B��6D��\I�-�*`J�k�*Od�䯖T��-jäA�.R0��'��q�Г�psEI�sG�3�'�����C�.u{�a˲�8��ep�'��b�-�1G�����ɖ	(C�E��';��#4A0�l����@/}+�Z�<����#k*�4�Ї�+6x�ؠ��]V�<�7�F�m����7.��O����WR�<���3&�T`CT��>{��|�BG�X�<�ҪE�8��\�c���N�6`�U�<���<
첕k����J��X��m�<i��_�B!���̈e�Vx��A�<�a��$*4�D(F�r�b���T�<��L�2kv���+ ,��d"��L�<�晼6�3��AJr t����H�<1VJ��e� ��
D�9�\qQ�jVK�<���G3��c�;*�Y�D�<���R'W�f�+$!�6;��xRG�x�<!0�8q�
�1��+$Ĉ��0�r�<��h�T/�, 2�P�]���apD�I�<�cB��o*� aE�Cz� )j�L�<Ie�ػg�i[�gLs��h�}�<Y���t� |���H�ɺI#C�w�<ч�R;v��(�!R5{���N�<��.Q�^�����Ɣ�P�GKs�<��O�%v�w ��7@:Lth�n�<q�-�-Sɜ��"�T�'!��Ac(m�<��œ$���$�H� ���r�<�"'����rk�S	ƉA�
�q�<�dk�,툴[���M�B�ـ�m�<��
�8���Vl�h���0��e�<q�Ɗ?]<j@9�C��G$�6�	f�<Q (�z�N��۾�l���J�<����>ߎŹb@K<r��Q�F[H�<9D���m-�5
ClS9x�|��bKK�<�b'�j�붇@�$����(�I�<� �9�u-��=*�pb߲�jؓt"O,��e�$h�H����NDB"Ob}��A^V��D���V�8D!��"O���7�?4�= �����];V"O���r��^AV�k�4༑¡"Ox)s��G1Y��話,���(��R"O���"J�w�<	�U!O.d�A�V"Ol�k�ܸP�0��͠��X��"O$���'a�L�-@�$�(q+4"O�|�TG
HTh�G��9�d��"O̃����q�@�I~A�Hg"O�$���8rP��(D���ܸP�"O�16a� y�u�"��N���x�"Ob��EFǽe�M�"�71+�"O
1c��Q?&��� D ::T���"O�qK����[����e�$'�Q�%"O� K�C��{����2��.�� �"O`�0�%� F�҆ %��p*�"O�\(��!:���{bE���``"O =2�"��b�����=o^ܵ�"O��&D`L�#'$Xi0�:�"O�8���w~��h�G�IV| ��"O�z�+��|s�yQ�lX��B��E"O��O�,^*�8�W������"OT�sA��%�,\��R3OiR�ɗ"O���ۺQ���
V��)^�,��"O��� O%@��ԉ�ǝ���"O��S�Q��(1�	�=�Δ��"Oh S��7����oO=M�-
"OT���P;C�d��Ne�h7"Of�[C�(.��a�j�
��p*�"O��k���srm��G/c����"OxLBBBHJVԑ��[0kѴ�A�"O���7�ݺ)���p�Fi�J`��"O@I:�J"0��q���V65�:H�D"O�����t;���EF	�|�:頓"O��	�e�_6�8���<�(!Q�"O.��V'�L����Ȅnr΍s"O�\��%��T��̑�:Hf�1�"O����ޡ��a���TJ�T0t"O��D�k���s��:+�9U"O��{b�ժ_Z0!cebO0*��"O��p��_c��C��F�j
0Њ�"O��4$�<&ޜb�>�
�"OJ�Z�2���Xӭ #�]�"O��B���T�Dd���л'��٘r"O2�sq��;��,#ޯb�����"O��Y�Y�Z^���H(.И)2�"O�m9@J��z��ܑ߲c��L�"OХA�� 7�$PH�(T�L�#�"O���&�Ǟ]�����G>"^8r"O���0�J="�	ۀ�`p���"O�I������uhݼ?�(�""O�Y�oT)9J.��@A�/�P+�"Od�LF�(��)SS��]ƶeQd"O*$#gl��r��h"��ϙ.��ra"OR �� �:>:�1"�٦1ڼ53�"O>, ��Q2�,m��N�[�H�Y�"Op���){!��A&&5q���P"O���A5�h�r�FӄJ��	"O��s(xJ�x����o��"Oz�;9���7���eʡ"O\�kå�|d�R��n�
��"OV�e���R��531�:	�yR�"O� ����"N�E��̝�pp��"O��d�J�\`zqq�j�U�h��"O�T�P� $?�0	�0�E�g�:5K�"OT�8��X���<����䐃f"O���pW>z���J֫^"b֠Y"OXt!`�)h�0) AJ��f�"b"O�y꓃�]^�Q-O������"O�tH�e^�;��I�B̌ U�>�+c"O���gT�-�4S��U�W��%"OI�Ä�����e���y�!�"O��*1�_�~giĈ�.nJ���"Oze�r��2,Xp��a��&U���"O���_:y���r.�7x-�U�t"OA��M@��4T�c �!J"^�2"O� �TnڻL�,�Fi&q�1� "O����%��ِ���
@��"O�9� o��~��P��%:�A��"O���E_�1.�9
P��+�2��T"O��Þ�u�eK��>�x8��"O����l���5ł-vc�"O4���i�X����b��y>x"OnQ"�  G�.y15A\�2��P"OB��'�ϋE X# >y�RA�"O�%w�$�d�3���D~b<��"O$�I�"^�P�-�6h�):��m��"O�d���I��X#�m�����F�!�1}�Ќ�5b��b�5!�$Y��ް1�P�=dx��Z7}9!���OʾIj�K:3���xV�K64!��e�����'@�j>6�x�CG+!���Q)ޱ��J�:FX��ە�Z5�!�ğ�c��0����lH�I�*=!�䎫�D�@�|Wr��VI�8d�!���F
�;���
A��AI��K!�d(�������c!��NB�a�!��[,dKx�2�E�7
�܊�k�=!�dD;h��yPJ�s(XkbdJ��!��=�Y��` �r@Sz�!�d��nB" p'�S�!��s�aX6�!�d�"�x���(�&]�\��U�ܘ�!��>�lѰ��JS܀t�F��M�!�N�S�Z��WDC�=�Ƅ[կ�v�!򄋓E�B�"3��3'���goR�8�!�.L��� �N�I��PEY�'�0}Ae��x�d (�H�8����'I�P�7gI*�k�88��E�'J�M�w�Y�,� XC�d�"���'�,�Zp�E#J�*D#CYm��X��'�ݚV�>G�0 �cW�v_��k�'���F&οa�F��g��`�Q��'E���C9p��#K/N����']h�#�$�D�����`�6M�=��'"$��7*�A�
���cܜq ��'J��"�Y�^܄i^�)	���y�	L�h4�	1kǓ`����cٕ�y�a�5��)��\���JFg���yҥ�^��e�j̠�%K���y� ?;v�K�-s�D<ieb��y")�d���Ė�uN��D�\"�y����@�f.������Y��y2�(�& !�N� cJĩ8����yr� QT�)�(�TiV,s����y"��u�X��g�B*P$ 	�����y�cZ�&�f+[�Kv0 e	5�y
� ��	t�ʚyi�l�6�ē#� P�G"O�9��e t�ȷ$�}��0�V"O�MP�m_�'�RL��.ưZH�A�"O��;T�ЩZ��0@���=C� 0�"O�x�iJ�|Ph����[=C7L�Q�"OXjB�ɘ4�|ɠ�ĕ�[B�(�"O���
�*��(��B� 0F���"O<t���T�Q`��;E�N�I&�ݸ�"O6Es�@�(�dѸ��Փ9
�I��"O�@������؝pa1`^Ni5"O� iDk��AƲ��Z��f��"O�\ 6�J�M�hA�7*�|����"O!`��O�$a#�(�?0�*�pd"O�Yk��'%��jČ��G��zT"OpU���#]�(�����i9�x�"O �S2
Dl�`@c�fDI�"Oz�#䉹>�P"�P���"O�YxBP�<e�}+��t�N�"O����=*4ZD�Yut�U"OL�;�F1u,%Q��֯^�Xv"O�)�醥74���E�QT,26"O|�Ǎ�1��c��bk&,t"O�4�h\�
�I��̏�D��\��"O�2�ߥ", E�G�*d�0�"O�4S�k<�dR�L�$DJ�!�$��5��QH���m�j��7��zj!��+-Р +�ŏ�:!�Lb��}f!�֜[����vF�,���	U[!��.�8P� �v����A�\<!�R�p�A�g̷q�@�`rM�.L!��5Uf͠B��.EKyps�N"+!�͕^d� �>����,u�!��J�g�lh1��-q��i�'��.R?!�T�E��\�ŀ������;BP!�^��� ��	)dɖ�b�!��
��~D�S�<"�;"CRj�!�D��U��KA-� ^�	k��>!�R��
�i����(����!��q.!��3#�F�p�Q�	�3���$ !� 4(Q�Ef!�~�r�+p!�$A�7���6G��8�T�0Sm�K!�ĝ�p��Ts�熡 �ι*�"
�!�ŗe���*�fNn�@�	Z�P؆�7�$��� EF41 ET�N�<@�ȓ�������"�6���F8趉��u��A)��ļ71����,�)N����BFJ�{�C�tVL�*�f��{B���0���R��;�$u�ьC�3,Ą�A���J��'t;����.6�4!�ȓ^�\ʢ&�3~!�8�Շ��|TD��ȓn�f�f���Veq���UX؝�ȓjR���Ta��攰4��$(=⽆�[:
��F��=z!�Ej�$W�����]�Vm�4j�y�v��v��#H
0�ȓ��q����_'������"����ȓml��Lq�R�A�Mĝ:�$��ȓ�8���ɠ^��b˘�)D.(��9����֮�	]�2��`ԉ?����5嬨�7���)�i��!O.4�ȓ7` heZ���E	��(�L�ȓ6=����a�F/�Kh���B1�z%��y���f��y�f]��X,�HB�A8D�@�7�Ʉ'R��ȓH=�*F�œ��d��.��%P��S�? �cb��2L	��gg�j�1u"O*�7��NEp$�Da	�.a'"O��&�|:��yH�h�"O}�� � u�b�2C?!��8+�"O0����0^m��JpC1',jq�a"O��rr��	0Y0Lj4CS2���"Oд�1"�D\(1H��4"�DY�w"O��ل��z��qxe��r�rj�"O�@�2�M�ou��p`�
a�����"O�B�!~ߪ�;!_�H�XD�r"OL��*I�mw�;��)7�f��e"ORq�B�8�ri��䄢f�h�&"O�1i O@�L�Z���D�H(u+�"O���f��8�2`#%e�F�^��"O>�K��M�,��a��\36��"O�	X�K�$�$�"��B�E��Y1�"O�qQ��%F�zȋ`�MO�"O&��4J����n��pB�"O���&;���ғl؈&�����"O~�jVj��(�"��r��@U"Om�����a1���W5!`j�xT"OFh�2j	� ���tË�[�胆"O��В`\�4ꖄ�`e	s�<�"OlrQɄ�gӬ�@�
0bf��"O� �eJ�!s�UQgCOT0���V"O�ܡ�oB!U�p�����l+"O��jt�Cg��<��&�:
�u�0"O�8���	�8��q%N?H��"OV�(Ve3i���5�I�`��Q"O ��Фڠf}�K����L4�"O �gԏ>�v���?��`If"Ox ��i��%~BTx�!�/�D���"O�U�WnWf�X RBό-%�y�"O�92&]�8I�)s�UR���"O��C�"O�] t�`q�ȥB��S�*O��� �
nN��D�� |i����'$�qqR�J�oۺ��S�� x@t��
�'�4�86��s%.���7F���	�'�ҍH��<���Ӌ'-�x-0�'�T)y�m�!ox���Ï�2X��'��t�5'��B��� %t��'_*=�QMĊ_�����),zYN��'���`�n�:B�l3DV�g�B| �'��(��\�T*y��BG/��c�'�)�f�!<�b ��-��{�'�L�k?D$7�Ѳ32,P�'�^a�c��	dB�<bE�@�8���'���ɒmA�d��4��f,�pr�'7F��珻$ f�����4��ɨ�'��y"jA�ѐ��r�})"��'���d!BX�C�N�*�4�'Ǻds��T�t���1�M�(�� ��'�~<p��U�&�`Ai���4ˠ���'��h�\�`|��@tf�F�x�3�'�Ƭ�F�ީgP��1׎ͧP
Nd�'�.����Z�"'��c��;����'f�y2P̀�#2�	U��&�<�Z�'�­AS�7|�����.��)�v���' hQ��o�6��@���)�l��'?f�Ei��e�)I��X��'f*(ӥn�::X��
t\���'B�`26��nn~0a��F�J�eB�'#.q�Nա&D��څ$�B�0
�'���9�+��N�.@T�]�F[�0���� |D����o�$q��Iը@�0�s"O!���WJR.U���Lw�P�F"O���+�68����q��fj��څ"Ol��N֬/^=r��^X���"O����펈--��cʹ{=L��D"O�Y˕�&jA �#��?I+��+T"O �s�EÑ)�ȕyѭ^#:h 
�"O09z0JضX3��[�_
(Y$hs"O
(Z�k��[-�i��+�,[�	�w"O�)Ї���>���)Td'W�աU"O�+���]/��@��n=|�"O^�{2k* �A�*�P�j�"O�9�։�6u�|��i��z,Ao6D���b AWβ�����*���#D��s�(��xI��s�Ϙ^�����E!D���Vo� gf\{�'�9�ԥ뷣>D�\B�%�q<U����%�u&%1D�d8�+ �f �H��/A�9Sb�0D��R�#��`"V�D�j��2�@58	!�D�P`� d�k�����YK!���u��ˢ��23�99p�/�!�3Q���9U��<Y���ab��9s!�dA2�(<ya��"N�y���m�!��D>)y�d��j_���C��P!�ğ>1 �KSg+[MVur�H �Ud!�dB?R(�`� �>cS��*�bI�II!�ēڢl+� ��P�A(׎-!�d�on��R�E	':�08��FS�X4!��@.xɆ퀧�V�jy�B��"X�!��/���b۴T�֡����!��ҳ5�x��@B�#8���IS��!�ĝ(;�HA`�$�8?�d��oD>u�!�<&z~$�g�ұx��8����2�!򄒬;W���A^�\0��X��E>c�!�d��ƘX��@!=���qpa�%2�!�R�9��"�IC�:yBu��Gz!�$�I&�9�����[%Hʊy!���0ؼ�pf ;X�j��R� ?S[!�d̀�4��G$ج[iB�f�	1!�dF;lQX�����%N�ڔ��	,�!��(��,���Ĩ%/����L� �!��[�v��R���u�� A�}!�J�<�p�h�O��`�@Xb��0i!��{����v!��J2�ȂnB�f!�_>��̲�"�C:R����Q!�䔎�F�Z�ȏ�G�zl2GD!�V�!t���fD%x��s�K�(!�dB/#�� �SgY/E.�
r ��!�d[�^IJI��S��؁�.j�!�d�4�r 
�1|,�jdĈ/^!���� a�	(Qv)K1��0N!�[]�6��HFPlH�nK"W�!�D�Cy΍y4�i�L9����Ɇȓ2Z53�(N"4��گ9�δ��Mo����_��. ��I�|��Y�ȓr|�1g!J�L���+��M'*��Յ�J��l�@�2("9��G�
�ҵ���>�1�	��d\��*�	 h56Ѕ�e���UT�!�M`-ˆ��t��)3�.�Zr��j�*���p��ȓ$*�����Ѥ4��1I�M�F����,��/C^F,9��(����GP�u��#�vq���PD��>H����3��#2#�2V�$��П&F�4��S�? Τ��;j8l�"R��6C��q"O�=1egE$�Z5��"���t-��"OJL��.ΦW��Q��	֊4y�"O�Ĳ�hU<<�(�-]�*1r��"O�p�/�8��H��M7.����W"O����"��1чh��;g���w"O`E˵�K=s��ÅhU����"O"� � \�Qކq�d���@��Q�"O� b���O19�(ܬ8��l9�"O�|0���#t��:�%�0�&�B"O�1�d����(X���>>_��8�"O�0r�L�Ȍ)�b�Q̵1�"O@ �S�'}GVh���E*SCF�;�"O>��BF$�pu�$@��C"O�T5嘒I#����@ǂAj�"Ol)i���[T�q�����P���"O�-���W �ЅhL;4	���"O0�Qf�!3� `� a�>P&���"OzEӱ�H�7?�� 
��f9@�"OB�Z3�D	 e|q�.�0;s"O�Hp����cC��Q�k#Th����"O\e���)'��8R���1F�̑�"O�B1Nռ\E�5(r ��b�
|��"OZ)�f���=H&!L'a���p"O�=�Di>f\-�F`��`u���"OAV'�&6�M�FČ�7Df���"O2�!oӃ7�	�a�[.qސtZ�"OF��+�/0ߪ�ځ�ʷm���"OP����3��՛w�EP0"O8		���0{˼q�����t̐�"O�e��#X�"�>P�0gͫk��%��"OvU+���?,���r&7K�0"O���\�-�x�R�H�3FL�C"O�\��)߲=o���$�)8N���"O�H�r+u��-qS��8?-���"O�X�ѩ�kl0�˗e��҃"O�誃I��ц�	�Q6�d4�"O\�p
��qH����?��`cr"OX	����H$��B�����"O"���A����d�A��01"Oٴ�o��$L�V��)0"O�i�ǘ�E0��Z�+�s��B!"O�32Ł�^$�IZt����	�g"O���@�Q�Ty	���E� �"O�0���)?�L��K/K(���"O�Xԭ+�R�cޏ~'VL0#"Ox��׎$x����'�>t ���"OV��[�L����Q���/U!�D���|��Ν[R���)�!�d߽ +��9%*�&6X��@G"ԩ6!��M'X6^ cc�%SL��Á&ęzI!򤉨��b�#�&|:���1%�	Q!�Z�$����'B$P�$�E�5�!�Ď? ��x𡋲!6
��F�Q�!�䀏�̙uEԤ ���r�ɦ�!�d�V�r֧%�X�p��JE�!�d:[_z�P%E7E��\ �lG$�!�$߾~�!Hd�R�����J�/v!�Ĕ�2~�Y7MRft>���܊-q!�$��Y��ź��U�P[nٲ�IC�pc!�d�wBS���8J"L0X&T!�D�9-�BVJ/ 6����˞�FY!��E6^�+� \���s��
6�!�dR�Nӂ��9R��c�˘>A!�� Z�" ���l����H;]fl) �"O�|Ju����`Eό��Պ"OȌ@��3���4��q��@C�"O�́1�A�1�L*F� Z�Р��"O�A�g�D�ItZ(�!!�+ijT�"O�x��B�����P!Y�5Z��"O�3%�m���W�]'&H��@7"O�l�UM�'RHFljӯ�v�
`�E"O �9�"ƴXyv`x��V0B�Dp۲"OL%2�ļ\h`��#Ǝ�'q�M8�"Oy(Ф� ���K�?[�"O��h���@��࣋ �mRx�"O �H��ެ]m���)u^��("O���hufY���Q)g���Y�"OV-�#Lŏ<��Q�	��y�"O����Z�,9<���	�<,��m0e"O�Uc�A҄M��2���b���"O�}a��T,�N�IQ�v����v"O� H�!��<�r��Υ@���	�"O�t1C�x���&�ҏ8�"O!rT� ;1��A��=ʦ�a�"OT�sC�G$��Sg�e��9�"O��`*�=U�r1�Ӽ�^�`"O�8A���+������+����@"O$�j4��[D���#)Ӝg����"O�� �i)]xT0R��Ǔx��"O��a`��<����غ�>�x4"O�U��.�,���aI$j�<W"OP����F�"PC�*_�8�P�Bs"O��{�  4hy�JR�~�`���"O�$��E�� ]�|Q�NՌH�԰�"O6�����j���8Ī��a"OQ2C���� ������DH�"O�1a�P8���ч�"U��Q�"O�Ё���<w���ój�a�*�z�"O>y���g��	r	�)�����"O"��g[�KQP��0��X�bJT"OZ���K�I*Vl�P���͈�"O��2��/qح���ɍB��۠"OT��b��U�2��E8��P��"O|���J���Vaߥ4�F���"O����D��r�$�C��r���;�"O �e�8P~�M��	;o6$C�"O4Y�f-R6R�a8���uC�0"O�(��E�$60�祟�r,jP2b"Or�)�kC��8��pD��8	"��"O�!� �'k�%�LB�E��ɛ&"O=`�D�s܀����AS�f��`"O��� N��3����T���"O:u�m�&��MpmG��4;R"O,m��E @���0�FH�`ڜHٲ"O������,ѫ��p6:��C"O��H93�YH2K�=Q�l��A"OtI�'�?;�6�
Vi�(���z�"O��y֎�/}F� �W�o�VtX�"O���S*Q�F�5K gO�	{�%q&"O�����H�e�;`FV_jaS0"O6��H��~<�&̣v�\���"O2ذF^=fP*�&P�(����"O*��#��8��ժ���H���I�"O�y��$��t%�eK6ft�!a"O�<j�n��1�.�Q�Ny��!w"O�8���ծ[l�P�	<�S�"O�`:!HB�B>�Ȃ��(r���"O� ,��tl�<2�b�k��F�rn��ۂ"O�-z�L�-O{��a�LE���F"O��xEA]3T׆(kD�[.�2�*O8��K7R&~��bK�'�n�1�Bb���P���t�f��'0���+�;?^���Jƴ��'�� y��6.*nj��'`�Ju��'Y����O~H���I?�Z�0�'���X�H�5k���3�8|�.�q�'����CP&�6�cg_�HU0���'��Y!`h�T���9��X�k~I�	�'^���d�$E��:qχ\1�q��'��Y	�j�$4�꜠� ��Wz����~�MV�y��)�dID(l.���Lҧ|����U,d��d �,�lE� ���"�!�d@<P��Y�� M�ZY�U�?x!��� L�d�rkOC�*�#�b	;�!���:���T#���Jh�!w�!���,�:, ��
�,��a��� x�!��	<�d�I�h�@d��Mў���7+��	�(F%�y@����A��D5��!ef��/���'��Jv��I�
�<	�O�b��| �Q�%�H��!H�H�X{DD�t�<1'HP����D�7(�̬�IE��hO�O'H�2�n�%Ȟ}8"H#Q�!	�'׬eڴ
�=a���pEHV�4'h��ߴ��'?�x¤��3bf�
Ү��٠���咁��=шyr��H��< A���l�A!I��?��'7�Q�J�L��<b#)A9�"�h�}b��8�S�K���&͔f����5#��.�vC�I�v��ib%Ǘ+W@!����H���%�I�\�Ѹ���  ]B�s,_"_"C�I!U����OG�> ���w��B䉂��m�Foڅ:����1��6Pj�"<Y���?E�Tg�2���#���7�"�[&�i�,�`�)�~��Ě���9|�j���|A�I�ȓ)�<�R���^�BA�|M�<��
ڤ�����$��h�T�S"~x�'wa~B+%EEi�3h�9rL�u�����p?��O��Y��,�>��._�i�^���"ONX�u_*4�ؠK1*��1lBA�d"O�yǌdg@�����`���ba?4��z���j�aA�.Wl2}��'(D�tJ��О~�lMb�c��a�	�#(D�`1�HQ��A���r,�tʇ�*�O��'��P�vM�@V�,! ���Q�'�8$٥+ȱ6"�8�,��	pL4���)O�}���X/J(����[�R����"O����f-v �
�(� ;X�3O��	sܓ�hOL]xbDӶ�H'���0��c�"Ov����S|�;�L�?,�(d3�"O��9��¢��|QWkΒ3�yc�"O�"�Nߕh�@��G�a�D0xU"O��L!3�J��m/�~�qd"O6���\Y�0A�Ӭߦ(�$�30"O��#�=[�q�J:�<1 �|�'��]�� �+B�[��б�����'�^L�q(_�0��EjP�A�r!FȀ�'RZ�¢��9K}�x��M� g���O��=E�4'Y�%�l0#�
�fl�䣗-Ӥ�y��А_� ��V%�]��ě�OD�y�σ�r��
�&/Q���J�)V�ư?Y�'�敫U��& �%9��X��8@�'�ri��L� ���'� .j�A��?�觀 @�B��T�4���ɚQ�q�"O(��D%��0��2��1'ꘄ#g"O�`�!�� ���U�%g�P�1 "O
� W�P !�f��acƒnuB�!B"O����N�|x��qUZP���a?��)�?��qM�1��A���j �$3�O �
��J#U���_8H�xy�"O^ػ�n�yJy!�%��ac�|��"O��B3`P;@Ė)#ӄ�3kG��!�d5�S�S�2�ZQ���;Z��1F�<y�<C�	�|wx9�JƦ>�D�I#� �jZlB䉌���j%�!�r���G�<7NB��RN��:��*u�B��E�G5� ��hO>�+�j��nODӃH�"�����1D�D���	�pJё�O�c�T��&1D��1���X�
\a�i�'6Zx`+T&/D�����yn��)AC�4%D���5� D���& 24����UæM��l�Љ=D��Pm�,_j��a3I%�̛&�9D��X@�uZ�\�'kʜ@����6Ⓛ�bIa�
XV,^�q�N�[��"O��8�I;,��y֍SE+`d"O����!!F�m�6u�<)X�"O����c��d��1Bߪe�l`�"O��C���`x��{o��P�"O����V́�C
	;J�4B"�'���8�D�*a� !x�l#w����ƍ[H-T5�'��Inx��1���!)`��*>a�	�a.D����/�>N>��y!��(m:b(�+D�8p��"RkZt�OmOn�+ 펳��'�����{tA�"u
��XedL�Y'zI��0D��z�o l`�s5�"WF>!Z�e*<Ov�}"��8?/���?�F��̐�0=��'�'R&��L�y�ޭ9N�N+Ź���	��hO���&	�<���a��A��� ��`B�	(,o�䂆읯 �b�`RI@�6pB�I�Iw��XG-��;eZб����>B�I#VΖx� �Ƚb!���c���"ꓰp?�S��ɬ`�`ţ9�n2D�f�<y��ܭY"a %��E���`��T�<�p%�W�����y�Bu'��X}��'\p9�K)�L��l��5)~YH�'�d��a���3�=���*�<�y��"o(�11�O7A��57�'1pO��>��?a&�A���)H��B��߬e�����w�m+tN�B�0yk�'3��QFx�R�hG{"�F�1n�3g �2j�le	7k����=)�yr��4P��L'.�i��޸�j��x��1<OL�p� V)L�z�	s�Z/�z�9�'�O�|�lS�|��A"'�y_��a��&D�X�+@66�4(
!M�5��U��$��?I���v0:1�K��� �+Z�niNB�	�aY(I��\�*�rQ;D�W:�'ў�?��p�CuR�����7$}�	��� ғ�'�1�0��@�׈2D�jA&���^��'M�z�f</h̭�J�CJ�1����yr��/�����=<��%�#[��y��>��I���8m���f��0?�(O�)�4�,\�QF&��\m	"O@��(�ycvL�ťV�X6|�qs"Op�{� �
�(1
��Et2��V���)K�s�(	��<��ӥ��)6X��f��F8�8P֯;�u�����[LD�k��)��l�
f�T� 狢B����q�?I��B�)� ���b,��`�KO-`d�Z�n(ʓb�>�uzR�se�)c�40�J_3�5��qg4a1�A�I��S�l��I�6���,gj���HRs���d�E����D|��ӥL2�X4`�3x Q��N�v�&B�I�D6D�ю��}29Q��]�v��)�	�v�8D����!/�H�C �	1kj�d,A�~!�X�ZjP ��㌦.-��a�X�!���(� 9! �O�u��Hp@�K!�dӅDNV�������߾[1 `�ȓb}�F�>�Q � Y�$�Ɇȓ]�P]�!X9;h����J�*�0��ȓk4`��K�-b�<�qpd^�K��ʓ3Ά�A�ƌ�$���򷋕��C䉸i�:��A�&�n����O�"C䉼Hw��� A,)��Y�oP�^�8C�	�A`��a�  / !¹)ц̟B�C�	
��<2� R���]{ejL�=�C�I//��1�l�E����O�q�B�I�M�d�Y�JSv��SD����)ZF�!�9e\`1� ;
	���ȓ	!b`s��)5�:�d�A�(r쵄ȓ^ tUz�ʏ�=��AG�@;h�z�ȓg�.9���/ �20�ᄶ4�Ā�ȓ1Y��샻.6,���Ni���ȓ[{��s�MV����'�A��~`J�렠�O;~5f�3���ȓ^\.��@nݭ8*Q�FH[k��݆ȓm��5ۦ�5;��(�v!�6:.�ȓcR���"ߐ��H��\�BX���`��݉�+E!)%�|h�ܼj�@���R�8���L�j�ec�E��u��
��!��K�f�:�;P��V�`�ȓ�,��o��6������;k�P�ȓ=KVL�q�ة&�����ɷ��|�ȓ*�LR��lu�F�C�k�2̆�O��p�S胎j<�3���_;����V��$�'�K�@�^�bvSz�����
1�=P�g
�c�@]��CI ���)@M����bY�X�	ٯ��݄ȓH��T�H�?���̍7nԁ��rP�Ѣ�ƊPs�A�G�d�N=��+>�0��ͱU� ��s*�+�x0�JMC։�n-:��C�I�9����̉)���{q��,��C䉛v�����M�u{���I�5L�`C�I�%�@�0�M�-.]�-��$R�B�k����KH(r,�I�ԕ0��B�I�n�b�pA�ybZ��F/cLB�o�����%8}m0����Q��C�	)5]B�؁cӌ^����a�4 ��C䉟;uڍ�એ�h���X<�pC�ɏX.��ٱJG0RW�}Jghحrl(C䉤.�,�d@U�	2��w���`�C䉄h��p�v�@�:��f�2d,�B�:50dK$�ʸ3
.�����<{eC�	+f�����ԑ~�r"��)MD�B�I�-��=�5e��G̦L3�c��f7B䉹
Vmʠ�� z�xp#�D� �,C�	
2�T�pǐ�x�CE	G�#�4C�	5�
���!ݮ,�*\ʢi�5D�C�	.2T���(
V~8(��z��B��.D;~��F�T<9�
$�N��B�ɦh�FD���=NYܕ(�.f��B�ɘs��l2bC	�J���'T�e�B�)� (���ϐCy"%8��]�wxp�Z�"O���ţw�$�#��Z�vX�"O�H F�Z�C�L�fO�AIx����'Hz���gτbV�����N�.)as��. Mr,8�&Q9�!�dL�v��cd�5l�Xd�qCT3YQ�@!��&w��{T�ĵm�\`$>M����SB��څ�[(P8`+Uh$D��(�Y�9����N;;�.#DkG�3=�Q��aϊ.�N���jB0C�v"~Γ@Fx��X�Y`��#�P���h%D�T�c���AZgB��g#��B 8viq�.�%v!jqPV���*�I7�X�� QM#Vr�@Rġ>7�ۅD��3sH�\��!H�Z�|)	��ĘD���cQBèP������R��`�ʌ�qB6i*��
��6q��E3���L��e���)6W�-��,._@,��Y>9��G�F��`&Ɯw��� �o-D���NF.6���bM��`?��@S�	 j�v�:�a�(�2�RV�7������Ӽ���!{ɐ\�1% �^N��g�<��ְ4^��Qd�A�
K��J�l�i�n{��M�@����(�Pխ;Y��di��$��4���&�B*����)�DVa{b((rshK*r��L�W��9��K�;2��|�Q,Ͳo"�D9uk�	��|�e��8����3�SY��l#��'T�<#CȎC�������I*@�˳3��擅V6�	2Ea���U�q�Ԉ8f�C�	.W�0�r3�O
Z�BԳ��3��B�(Ҩ2��5OE�.�$M��Ù�U�2�z#��
[�@��1��ݧ"�<�#����b�����ml^C�I/�JT��X
P�<M�
�,�P�a�n��O3��P%Βu��(�2LD�@�@@�Dc�T�(eHwK�)�Fʓ?� cBI�N��QH3c4I��㞠��C$U����'�4�&�M�4����6G��!K�
c�	8'Ӡ3��#�$��PF_�2sjdxa�z{��3�
�d�c�X���|��  P�Q�xF;��K5q�:)���+P9(�x��9}��E�\��ѐ�����Fn�e���GF(�l��%�y���`Ɖ �g��걨F�^ZF��I?ڰ�����9k��*�JW���6mK�?�f���d��`�)j߲��ʝ:m����׊�����<|����@ @�|��w�ͯ8�~���'b���>xjr���#W�>Z�@���[5m��p����5OO�|8���%{�y���˶[�Zy��tS�a�7��7k��t�Ŏ�NK�`xg�\'~�e[�::�@��0 �`��6��E�d�b��P1mU��Z�AG'�K;j�`� Y�B=��J�vΝy�� q�~�в���^�20�� ]�M{�NݎX@��b+�#<
�{s������eTO��)��M� �D�3��S��ȡ<~F�� ��	�J(���;QА �3ge>I�0n�0
��s��� 9r\�� k��2ߘ��W)
1,�\��gIR�@@C�X�|���Ac��'~�1E���5р��/ڹ*T��PN[�"Z�  ��J����⥘3����c�@1���8*R���n�!P�@��L���k���oYI�؃� �I�i�?g�Q�������Қ	 @L�G�@�s���%$���JH	jl�S��?$�f@r��N�+�����a��c�~�c�J& ����k�Ԭ��%�`Lj��I���:�Ĳ1�@�a@�םe��d`���c �,<�XcR�Й�M�,�4Qq��b���%?�C�H�S9����)C�&m�1#��b��x%�L/��r�쓥>�k�HQ���=� �#�E73𤙣�G�M a�8g^|��8tDAG=�Ӛ8pH�]�4��A�aU$Wl��+�,�".�*��iNFYJE&�=Tø�"MO�Q��	q���T��Ȳ��r~ڼ)Vǁ�|�*��
���>Q�Ǎ۟��G/½R������usҘi�� 	y�<�K%�ȩ��lA.��J_�0�4�,�.�2q�����E�d�!O���袯���Q��(8��l	P�3C��m�g���JCp$T���{��N�*<��|@�?��;&��d��;j0I�N3t5�@�O0�@�F�6b�z8�"�$�>���/��Y�N����+rּ@�V�҈-�@}�5��{1��7m��h���O��Z�^=�W�j≦+�B5@����taJL�e؇p �u�B�T����.r�6�3a����_�Ipǂۤ/�H)`t
V�z�8]YR-��|d�%8�+كE�t��(� �L`����0<q��!׀	#b�M�H!Z͛򢘙-�~ z1�X�!��x��),�����Ƣٞ9KB/L+B��""�)�tb�ٕn��X�R���U'�%0PF��6�����	|�HdSP� ��$�1z���DG�p����e�/9�H�[�ڊL{ԄR�k��P0��K��5}���t'�*q��������λg
����Î10tm[׀��F	8��=aP�ȣ�Vc��{pN"�^)s ��/:�l����\���Ѥ㆗t �����z��ȱ%jȵ��݄D��D�a�_�#wj��=��̑O�n��5jݷl;�5s��[�f�>�I�� �R��KT:n�x�;V(��0t��R���{ֈ\Zq�F�`L\R�
* �����I�.~h!���e��PiU�A:*R2��B�X���ԕT����!ģ`Z$��J�]�Vy1����.^�%B�\�%ӕ�ԕ�5�����#B�Y��$��3��y2#	�" ��?HԳ��E-<�ٱ��C'���Y�#�� \���Y�L:XjAI5\��1@,>�ɭ��5A5�̔].r�{4���������I(	z=I%W�8[�`�V}�È�:��qѴ$RuRms��ۃ]-�-���_MH$��'�4CӰ%���m��a��Ē� }�O�����B<KB&�1*IB�,�;]\ �n��<�!R%p����0�D {�H,{2&�9:ilߺZ�U��ٲb��� t:��!"�"x ��E���x�lA
�Aj2Щ��ۭ3��S�
�J���0�#��r,O;&���4+�E`$��a��-3��C�j�J���1v�Ij���}��t��.ڞ||ܩ	��'�(����ߞtmNi��R�? ��c��"06p��tƜ�R`��7��"s�Q�eb��	l�/��NL�l���8�`�el��'�V��U�h��r��gUޤ��{b���)hB�A5"�9t��Mo�-�d�9��L�?�D�1w��;?e�xh���#�6I˅�N�(Ad���f�a���Y*�6_-�|�'B& �5��R̓9�Q�h��~}�u;�"M�)�頓��7U�чg�7c)М�R�=�yK��}u�][F�*/� �����4pG8��M�M��$	8Kjq(G�c��	�ή@�fɑ��'�f ��hhr��T	[-o��� �Ɛ(������J���v�Q�z ���nb����[�o�
��`�)3 ���8@R�`�%�Ƞi��YCq8�@a�!��&���{�'�B�lQyC[M�d��7Y!zN�x�2��1=���Ԉǉ\�����5-��IQs�
O�d��g�٠xK��Q8�5��T�7& �1�O	1����F9G1O����F�;JR��C������/ؕn��Q�ԄxcB�j�����OA8|,��k�3^>`�ƈ�Z����@�k�47�.��3��u�D*�O��$�S+��.d0�㏿5��ZǄR2V!���D�O��c��ϨrG>�"�-A*%ʢ�N=3��2Wd�S���0����d>��r5�'#�rIm�B�� �F�[����$n�'��:�#�3�]�P��?VFf�0#�!A4��YېJ*��Gj	o9d�F;;o9��C������Ƒ0G�ZMq#O�h�X��@�4�%���T�5�֢?ia�^��2�+6H�QP���႒�Ѽ�2a���̤��9$:)�`[,��k@�͸*P���A��#	ެ�ZqN[?�?�2�;��[��܀G���tJ��` ��cAu�\�)����0K�$�gn� o���tV��\�S���P��f)%�& �Ea�0�ę� �k�L�Q�MB�Y�Aӈ Z��Fi���$�2aHH'��2n�5���d��xc@�w�t8�6O��z&�͔6kx(筆6f�)"5��)f��d9#�"`(!��?J]�E��,�����ٻqđ&]�`�Ѫ!���ƥ����n��Ȧ��WSq�Μ� 2���@Ok3.�@e�%�ʽ��v`�qJK�K/��G`S�`�D	�@HpL4A�Y C:A�'��p�3A�pn�G?.�@ƫ	5v�`�b��n!�P��Ӊ`��\���R8�L��BЌC6:��p�r��#΅k+�}�u�wgڌ�6I��!F�<��<�P�Q�a\��/� %be�ѡ̦�Ӕeɪ9)f��i>�ș�iRHV�����������	��6ٱ$%�(:/lȐ�
9���'N�&Ӵp�E�Ce�52�x��dF!j�<zF-�o�$�ۤ��nl�$�O��i�cGg<�fK�_��ce�"5x@Q��c�J���`A
<WaxR͊8]���z&ETJ�Q�go� /Ԩ����(cX��ٷ{���b��9^���"�%��PB�E�W�܁-Ц��e��$  a�Q�"WY� ��f���D2L�������$QG�<�7`�|�N�y�KP�l*i*%č} ���n�G��{A��PD�$�'`ܲ}�Z�1$��8f��Y1z����a/�p��`�k7��|Í�?�4;���+>ɜ0�ȟ�;G�TZ3aު
�,���ȰZ��Պ#I%2�����(:�&[��ݢC䉤1����Nc126���ْW�^�m+0i!%�Ҹ  #=	Qh��]�b����5���*	����Ы��ԇ)Q�p1-�<�f��g�Y�i�\U��Eρ�M˳GQ5����*	X���� ��'$�ٳ��/ƒ��CF2�v��۴{�P܀�X0G�h�P�׬=uBH�iDU�	k��gj��Sg7}�^ 2���)Wp��B��Q9g!5�,�b�V�/����	h�u���phP�2ߢ �P+�o��rg!ܽ�5z�M����l��f_�p�͓��Q"4ݤ,���	i���G��k3ԉ��MхDVŊ��'�O���!����M8�
	�n8XD�E�B�:���L��e��D�� �@ T��iC���MHjH�j6`��DD� ��Q�߆g�B�i$�[R�N�
J�B,Z��$̣p�Ј��.�t�@xb��3D+� �Q/�0�ve T'�<?X��mR��K��ֆCqx=�s�'[�2���O2�|q$�7�	q�d-kgA�=w�f()TE[5&� ˓��!��dP�iߎ�Z�c:Z��qH���1BM�֍�,D<ʝ�k���X�XF씆%T=�� ����h�.�c�ZI� "Uc��0���HN����Iƽ�x�ף�����d�	�p��.p2��^��Mk��~�ɲ���$חe&�rB�!8�u�)�$��O"a1����������e��~�l(��>��c!d� H\&�'�#J���.J<A�<�4e�z�p� ��?��#�dKZ61)��/1� ���,)��Z5�N8�*��2�I@�D����ɀH�*@�/PH�����
�!�^�c$���r��nN���+T��@�L/+�X��^g�n��'��~'���{�	�*[�B��D�<_D��*�p�����/YH���e����t�PWiX(]�F鮻1�p(��G+^7�I:&
b�@K�C��Dcֻ-p��
2}��!�<Z0`��=$"���aP� �9E2T6�̛"�*)1t(߈�)9 �bi܈A��F�� ��P��#��#a�S�&�- ���5v_<�"m�Wm�&RT2x�dn�-��SW:`��n�/(���3m2§7{���D�3cV�`Q���$��rt�)<L�%+f列� R(�!EA虚s䘰d[�L1p�@� ��zD$�(8E|!�O�\��)�!�B
t�v��#㖐l�������?I��*::���]��@��h4J�QKȶ{�����W�r�a�m˫sGƤ!Xs������xNA�R�ݓ2l�[P ڎiNc���v8Xc��[4?�d@I�n-���炶#�a�#�F`�ց��Yp:H"��6=�j\q�]�k'�=�����.���,̟A��@��=+���rᘸA��"<�ٙ;����©�~Q�%H��I�*Vn%�cE)B��}bC�5.��P²�!<[��bԈ'6��I�"j��.^~���C����!aѨ�λWx�2�a�,Aلǝ"A�be&�P���9@�r��4*-Z`���`�YZ������'A���z�N��E��]��� �D@���A��Ԭ]P���E-O!J�H�����f�_Њ�X Aʎr�F��&^�j+�=��M	�F������#������f�X`��Jţ6�^A1��5H�9��
F�lQbi��2Q�ܴ8��Qr��׌!O$����	$&�A���X�9��iG>V@1�V��Ab
=aeہ�|�#E!Հh8�I�&�Q���	~�4S}�����~%XHA��4�ቔ���{�`S=B.�x�i�?.I�'㛨[��	�@o�*8=8 fb��<����L� 	����c�d-Y�W��Y���p/�<qtI>� �1�d�(.�B)�pNؐv�z����x�1"�� q�X0c�B��%T�G�#�Α��%{Ʃ�;3�����֩0�K>^G"���Ag�6 ��a� ��I�%�-�$(ۚD�P��"B$��0���J���Q4��1/'4�9�Q�!�5�H�G�D(�"�Û"��@BY(H'��0��+>��QJ�MħV� B≉I|��B�P��:�Z�I-R%%�eDƺ,
���,/w��B�B�^Fb����=
�(�j�nI�P"��G�)���b�]�3��E��M�K0���pe0���-��r��Sꚹ"[*�:��^���e(��i�4�2�U���s&�W;���0C(�*�uՊ�>c5p�������~:�T�U�:1FT����]Y��'DR��׉\]����C�\�p�K��*|����%�i�r�(BHR�'��	*�O%4+01���� �*;���"a�l\Rۓ"AL5)��Y*�V;p�׋�� b$��q/���!̕�=b����%LTi��O^ CW���9��$�6K;X|�(T�T4
��""O�̈�jׂY���
��CW�E�T���f�J�*L���D%�7I��Ԉ��[���JKAP�m��)L	�$I�a�\�XRL����>S��)4�'�r�y�(z���<Ƕ��a��8��K�8&��AK�L�|�)kQȒ�d�ހk�*�4΢-�g��r�'l�b�.'P���ȭr�0"�B�G�28lZ���� �oQ�&��=cP��_~,b�O	.B�hi�aP�j_�5 �,��-�e�-�a}"i�:g��$�&݈0/��:�U���:eRD��
�<v4���]eY>�3%�xۃ�
� g�}8���K!�D��y�Ne�q
J7>2���*!rT��G���x��#�H�j7��|�/�<2]T�ڔ�~�eC$��Ԑx2�̐uC�����T'��5��@�Lyg_�<B�X�X�^��zJO&I��ыX��q����<�3�Y��V	!^3�y��4c�'���j�m\"+Z��wkɒR�� a�P��H��-0b1�=a�L���Ksh6�'dߨѰ֍�>���l�Y�ȓ+�:�+D��prt)�ュ2���ȓ-$V� �*�Z����0�!$֘�ȓ1����Ұg��pC�+w�8E��|��`��꘺ta��ڳ�͍�Q��<�p�Vo�ENعAr�S	uV��ȓ�!`��)~6�[��9\����c j��d�ɭ��cSmAqO&u��$	��uI̓CQ�%h�L�&=&��ȓ��f�VzFz��+�"9��U�ȓ��@xǁ&���{qb�+uA�i��=DdmC3�ޓ�%c���29��-D���3cVD�R��!�S�M��@2ĩ!D�2�J�'���B-�5S�(�E;D�<:���:NO����B.I����T�9D���
Nb��6 �si�`b�4D�!QjB�pO�xCEL[,�@]X�B3D�l#`�"� ��� xJI�f�3D��Y�B�p��2�c�~�8S�*D��37��8xԺ��c�H�M�&2D�`C�%�h6��4c�0�`���3D�@Q���.r����5�El(��1D��)�-	1'g-"���L�A�qi-T�\W�ǐUR`�����|�"Ob��j�Sj�E*�m[�g&rI��"O�`�Ӭ�5g[��8�jדE���2U"O��b�%o0\X�'��
I�b"O�=� �����BE\6� �"O&P#��	�)�ͣG��C�<��"Ojy�#�^EX)�F�#'��c�"O�< �	��2r��qE\�~��"O&i���UTJɉ'�, ܬjs"O�u�F���R�j��	]��ѓ�"O0a!��"��Q���碘�"O��x�	Ŕ�<,��jBe��I�"O(ܱ�H�=F�5'�2W jg"O��G �SJ�d��� e��}c�"O����$�@8� ���`3�Mr�"O���!�W�=�xC�P����%"O����k�9m�/�O��"O� p�2W�EwnL�v� H!R�2�"O,����)���ذl��0��Pd"OZ13��r~���B�E��"O�Q���	s�5�DU�Bp"On�@��H�N��UÊ�8Z)BiR�"O��CgBG>��H�hF>�,��"O������I��m�r.�A:j����';hɡ��)��\�3�R54A�xB��S�n>\A	p�M5<b!�$J�<Ǵt�"��Y���K��]Dy��Q)���򥗳��Q���� �O�YcSf\�(p(v��?�y�Ě2�.�,?�LS��L18��jB-�~rP�����g���c�o��yBc�(G���{&���i�n5ѵ��y���'.na鵏�3ٰ�#JPo:u⢀\����˟;�z()����O�	����Bƀ&U��
��X�4��{r���u
�h^�Yu*<���G�q���PDW� �&��!�v�7�'��}-�d]kfiF�N���c�G�y���yt�޿*������'-4�Wn�|�ІB�v(���W���T�B�<�� �6nx��,�~��0���U:�T:SF@�Z�&���-O�}R���+�y�eͧ>�n�!0�ڑr��*B�y���)$���2��%&�Qu��J�T�z"�/�Pd�ЂܒS�:��\w��Ļ���+J������G�a�@���
c���dL�od�2����Q�!�eį"�g��:/�>ܛ���76S^�
����}�����LG1$|x@�ݫY�Jt1!��^ƱOH���36H��P�@&q�p�zA�E!*|ϧ[w� #r�m-�t�u�DJf���u=ډ���Z��YӅ^1��x��ܺ4br����_7V�aY�@�v8܍����[��]�0��̻-8 x*V-ٗ-�v��_"ji8�%$�D��l-.���X��Y� '�T�R�
�r�O�P�B�BϧEx>�X��Q�,���U�ؠ.�pJ�ǳ>���,�䗬u���d�0l[�㞈C�6-���3[إ����jʠM��e2]���Q�D � @8�Ϟl5>�ʶrB�Z`d@�2��=�C�n���)7ā�Gb�\�΃�8O"�p�� 5�eK���O�8������Y�#شf*�E�t.:H21��M%?�qs^w2����1~��ЩT�/T���!�#vٞ�9�W��L��r��߰<SFԝh ���T�968x������Vщ�'��[�F<:��Di�딝k!����k�2?t���
���Hݹv⁣9�Ҕ� �	�h�g^�P���&�U�Ц<�t��瀑q$�\�5i�{������2"�QGB�Y���a���;Y��APӂȒr(�|��)Hz����hZ1*�<�b
6Zp����%Ʈ2<���k)Y��cO�p���5V6�����N�W����>�fQ��|��#1eɝx�N�r
S��m�!~���Ӥ$���T%8O�$[t�;&��{�@K0
+FE�Ӕx2�ql�q�.�� �)� k��q��QagV�&�(�����<[�Oph�Q��R&�-�@�3w��y�a�����`c �f��̸�]�m�Ū̜2�e0��
)�ޱG}r��yk@P�ӏ��m�(�**�.0J:�V��<����kҫR�Z���C>haTl-&B|��)+T�b�1!�4 ���s���bD�إ�"Y��f5S��!C�	;!a�}
�ӆ
eR�icŜ2%� +O�5~�@��G�x�X-��سA��D���A
Ad��w�T �k�O6w�X��O�\%�1�3@���� �zz�{�C�a�����7?1��ׇ���qC�,v�(ٴ;����0C8�IO)p�2",X=<��i�Γ!�)���A��:��)aNR$�5�BW�#À��S�ȟ��I"
J"���9����Q$:2YB�dC2XIfU���@́s#�%�Bȍ/�R8�0d�th������~o&90 ��|����Zc$��'�Sh���'��9pd�eJ
�O�9��IY�l��W��^��@��o�1
���Ɏ}樬���I�9�0�Q]�~���n)Z��t�0��43RexwŌ����vL�	�Q��Zs���s^�P��i�
k��d�ɞ\V�����$Ҭ��g��t����%刜~GN�P �+iv�����Y\���w���%��߼�$ĠJ]�v�Ԕ~}�aRAc�U����+��P�$�ǈ(W����I�x^���d�Ѵ5w�x�H�&W@��weY�JIq+�'ш$��t���O\����ж1�$� �G t3I�dM�Cک�W�y�aX���d��տYO�Oװ��`�ܩz���7�[$w�H��H�P}�|����p�
QJw��6���ZU�I�
oz���%���nL��R��(�劐/
�/�PL9�&T.��	.��	+�F|iF�, ��`	�-������b���kX�r�xuK�Ȑ.t�J�'���nQ�X��'mx��jS�&���	& �q@��f���.���Y�bjXA7��flȂ�*S,'���@��u�`ޙI2w	���W�ۇ*��1�@  �	�c�|(��Õb�`P`L�B�]�A��z�����`,�Y�$J��P	�'莹���A���M��]�qOԢ~�䔃�{�'K7v���ѧ�M�YX����!��'�4tC�m�@]����[�$���ȰD?�L��nJ/
	r���K���p3�a���� ƨ�.a�*H��p=q�%��r�Ĉ���'.��{W �f\��iw�A�\Ͳl���8u��#6�Y�w�ܠ�,&*��;'���fZk��m��z m�Mq�1���Hu!�DB�	y����B�`���daJ�Vy.��0���.�.|C��?M�pK��:x��b�õj���4��6W}kLv��,��%��U*��rZ�4Ey�%˓w��(�'����ݻ(T��Å�	= �jHH�CW @⢰JԃX�h�^�3r�FE?~!@�.)G;����oE�!�`PpģWB�S�? *����	D|������K���`��<Bj�X�@�<�+M�<ܸäW@{��㦒�O����؈|�|��%�*H�ɓDDV+pi�0��i �H[F��t�Z<HFf���T�	S�X�d��Q�dy�r�ĀL�F�Ѱ�ͷO�]re�V&/�\$����[�h�d�اS�`y�R΄�M�kLB>���ӊ�8&Ѿa�1��4l����	�n�nQ�!���y4/�'��quJ���(����j5VP)��MQ㢀QN1�%��Cd݉*3$�;-*T��l@�d 7@&��i�2Ko<D�����+qO�A[�-T���9R��M��fõmƬ�� "]�2e��
~L��0�95���"Ս�U����w�H�
J�3c.M�Q�N��'D\@"g�Y̓7:�)@�7�Je �V�A�&I"�R�'
6hI�+Ԗ�n�0t	�'=.�a����b5�A�\,}¤�E�J|��[��G(��PIP0 �|b�)o��#�|�HX a<��DN���0ć�$���!Bg��d&��r��B \!H�%|l� �ϫ�� �� ���R'�	f!�j��8mi�8�	M<hcd�Cdƒ<K����5��oКM�:[`Λ�?� �e�O�(eb��p)�";�-�n�0Z.���Ɨ��Ta�Y�b�Y.|�M	C��Id�����5��؃m�Har&�:SI��bn��71O��n�:�	�V�էe�����1,���` �o�
q��!�<B�F�YC#�0;Ǭ�;���D�a9��D�3�M�D'��t��A��Ǳ�L�v�Ua�#O�5m����@^ �E��G� 3���Fω�?�%"�u�YyЃ��1g��r �	[+�y��_~��-s3J�!�Q��f��t�8<�7�ioB��Rd8��H��.�f�џP�`/T�8 ف�B7}'���aT� ��e�B�2t��B�<<Ru1�@�,R�(�!��'����cU�0!O�Q���,��|�g���RmEb, �ТR��;WJ�[u	Z�i�!�r1;���ƀ��]����&JQ�)r#��lpKp-O��yC%h �?������$fĲ��u���[7 ����8����7Nx��=�KD�$�\�+�_�BH�>=�o
�DG�d
�%�N�:�J���<S�� #�DɦrTp����R-'�L�;��ʰ@O�DJ��:O�<�Z���<9�(ԏH��)y%R� ���d��q�Nᰔ�ߓU�$�� �b�$F����gɏ�z��m2jF�G�x���L�oy �kF�ε/��	��#�:p>Ȍ���B�c�h��K�2|<$�GR/ţ/2i��M@:@�2]+��X�Ms�E�/ڰ@虧i�	���J��i�9�Q/�B(���b�>\�%Jpa	-40l��L��/����B[nl�����M�C��A�
�k���.X�j���a/= %4��T�`��5�VK�����PD��S�K�.Y�`��ԁ�����ֆ}�VzP�S�(a�dA�j�'%Z���͖F�'��l�5��#~"����<
�X���.�\� 	�w �
���� ��9X�rɁ�ɒ!z,���[��T��U��Z�� ^�Z�g�$��Y*C�0�E-h���vTi��h�3�|&t`*�
R@�����B(��'���	�  %(��M�1@�	)� ���ȉX�HZ��̎4�����b��<��d�6cf���mO,ڌ�It��}6��z���jM	�DADК@��8v�A\��!$,��X��]P�f΀\z���Q�\��o�9D�4�B���R3��J�@�:�̅TL�(a��%����P�P���ܸF�8�b&��U<��λx�����(B��j\�+�������}�����!dB����D�F-RTi��$S�
<�&��o(F�x��#�az�	#jT��D*B|	B!Z'U� ځF�w���2+�q�@��f X9%�Q��h�@�(��rO՘m��{�H�r����01�N���
�g,8��!�@8n���4}"�I�V̄�X2�0�MP�cg�ڏ}�@Q�E����#n8X< ��B��~2M��tGY���+C>�``�)
�6`G�P5*�rTa�蘸zVD�A��Q0��R|J��aIqP4�7(�13��'�,y����RYz��oD�I�@ِ�*Bt]����R�T�U|�*Q��UUf��`��>H�D��'�w"�Y'�Ƣ��}k�&^�D:�����\�3.��x��h!�(ں/�ΥrF�?�b��g/ɕT�����l�; `��1lƟx��Di5(�,�ލc���<�r��'O����Ӏ���x<�5
�j������w8� W�P�T�XH��/͋h�$)0�c�^?�M�6��S��%*�L�P8<��Ń��h�x�`%�ܠg�>`5�B\9�Q�=�d�_8���@��7�z�ɠBVy���Ԉ��fBsS(=��x�2<h�쌨]f"��R�|jL�q�D�;�������5EQ��"#Bl���ꊎ;,BQCד��������a����-)�M�a��=���PPlxq��^���㑺i�����,TH���:}�xA���[�As�bU
\*W\����R��F�$e�?k?����־�F��^�V8���㘹s�d��Q,�j�+��a��,�;R���PE"@�"����!M_��z4x2$0Й�F B9@j=ɵˇ&���X�>q�+�~Z2�]�l6�kt��Y�v HB� :\�؊����!>�V�������@.��{�`m����-�;_���P��>��'$����Β�H�ʭP�N�v��[V���+�&�d,\�u��"� 8`/��b�R�#ׂ]�9��520�
x�(�l5�4pHq��6�X|Q"鈐C��3L!��q�{2�B�����"�KD�n��B�AoY�4�2-��@�$7��dAP�վ���	���I�,��F������(k̅Ύ�SQG�>Y���o��'���fo�L4�����O4��pʖ1�JE�ܮ@=�(�Pm�:�ja S`X�W���z���Ѻ���ׄ7	�!��],D5�<�@�;�x B唋c3�` ��a���qi%^Z�xF#���휝u����v,�g��3k�����Ł.�J���%��H�P�Q� ���%�!�4@*���
^�Zr�H?i^Z�-����OT`S�M?&�
���.�%�^IGe�S��>h���I3��0�
+&�����$6Dn���:Ѩ�jRhڞ~���ZA��,u����ǌx���A*����Bg/�3Y�� ��*���#�4S)�1y���� U��(��
�D� ���k���U����n@�R]R�[r[?t��� e�aݭ0�T�y��n!ǀx����$h��󴵻ɑ�7)�8b�aM!��Of8`t�o2Qç˓�&Ec�7C|֕`af�7z� a9� �7�^t#���`(a�g�"	��P� f�ͪ�R��Ҳ(q�}P�T	j�ͱ��zӒURf�N���
Xw���P�mV�b��}��� h�
� �%8+ީ BR��&+�!�6��g��M35�*\�n�C&y�џ����+t+@K�5Q�	X�@�>m��'��7 �u;�Gۂa�=�Cf��t)h3@l7Rz��O�V��0GW,�BF�Г&ܼ�R�%EQ�0�2�0W�� �V� -,��C�W�K�����(~�8�%W�ne��	�+[����ǯQ 2Z��!%kWH������Y|��]$�����q��)�Μ�q�r���i0�]�w�*�
��#uU��R�S 9�҅kGN�/5�2�eI)SҚ1!"�^8E���p�)+-"LU��$_�3�MݎE�Ĺ�
ϓ���@�9PF�ye��VR�#�	����+U�&R�lݲ�%վ��� �۹RA�QJ�l��[R�S1阎J�Q�ևL)wHH� Ψr'ȇēA�t�
��1�T�ɧ+�+�r$*毆�9l ��z��\���"`�j�
Q#��@��ǋK)�|bF��3���#�N�N�J-��@Th*c�'���rƥ�6��,J$f;x��PWLݽ	:�ͱs���d���t��Ƀ#ڞ?ܢ(xp/>9����,�>6������\D��M�%�3��
��T�n�M>�B�"W�~���N��D� ت���7*j"5L�<�Mk�H��.o�ų���wG ��c�4�2Hۂ&Z>O�LH7dRO؞�($I,;�z��r��/:�8kf�VA�ܚs��.�"��h��a�z�&wBr�1��q�r�	@�2s�b��+b��AU����`5�܅Bn���D����T1A��b�C/U`x"���<~IR){Ā_-8����Ň%F���GD�C��r���+_vLJD
ͿL��}���e��R�*�08�r���Ʉf�����ڑӲq��DJ��Ȗ�����g��)*���&��H	�IޚN� �X٢��`J	���h����-�iR���Y�$Y��(�ɤ#ɖ�D�i��h�I̽zqp���$0&��r�LM��$|�Λ`��u���H(Rț���.��}����r�@�-.p:��BZ2�'<Z��\���DR�c¼Bj F�D�U�/$��FbޑK���R5J	�y҈�*l��)�SEol�tڔ �6����#3)6�X��V�K�U1��L>Y�ɸ,m��j�I��]�nD2�jAkH<i�WO^��d��$��EÇ���w�x�y�DIC
�bb�ڴ�p=�`	 ���S7"�&"�ɡ��Izx��CBF�#|�Ź���:����:F�=a�	v�R�b+�ygM�_�*(�l�.0b�Y�r΅ݸ'��H)"�B�9i��F��b�OH�V)�3�(�	���y�]y���
Ր*V�S� U/�y��E-a�4	�˔:5����Ԣð�yr��etFy�%HU{b�kǏ���y���_[�%"�h˗
�8)��K��yr	�M�$��Ӱ)�P죆N��y�D�Т��'wF�� 7�/�y" 	v%�T��J%��S�����y�f��g��IC�E F�J�cMI��y����~9{Uk3���x�)��y�Ņ�bAv˶A�.7��� ��ڛ�y�L�z�I���E#�LӤ&���y"l8,�B���Kw���9���y�9Qr��a��!Q�Nd�EG�Py"IʆN����ʦ9fA�e��Y�<�EX���^�P�� �C���ȓz�I�"@2��u)х�'�:�ȓJ�,����ʵa��9㆔�tцd�ȓq�h�I�d���pU�dNN)K4j���WF�Ԙ�nV1xN���e�p@P��ȓ	N|�S��_<W���ӀQ���ȓ'G���EG�#|����k
�*�r݇�ɽ\�^t��倖X��AnN� ^$��5(؜M�0 �p��.w{��	.A��hJ�!1�)ڧzTx�L'H�B̻�&�.P�P����w��t��	�<kh��
�-�{>Y!sʓ<z&8`Mߗj�h��`ݕ2�>ͫ�A���y���i�����V �
���?������P=	���- ���s�i�Vҧ����	5#�9gR ���bJ/�޵��.�P2�{�43��S>Y	��ۗt6(�;�OD]��-��������&����0|��RIF��+^�:��̕%��A�	�d�$ث9K͇�.InL4�&��XbP�C�T�i����O��Ч�) ��%ɍ�)�D�`\u�֭��{S���t��	(�l���l�Zm>�S�O��ȕ�$��b��7R鞁yݴ�����A�"W\ҧȟ
5�Q��[s�q��h�.�j܉���z�%ǹ>	F���0|����-��QV̖(y����!zx�-P�A�)���l��b[
kW���c.ʸMq�i�,����f���=砈������3��4�[�ʣ6J�hj�'���o��O ��O
�;�q��3� Dx�%�M~/ڍ�4��y\ K�S��s�N$�S�O����!�[L��x��&G�%�f�:ٴ1�tGx����6,T�Ig����H�����}5<iGx��&��h+�@�-Z0����l�<���$������b�H�: �xYV�-;@\��B�x��B��O��� 
$�E�;�V�S���6m:��&\��᧊~�l�I<E��+�<MCF�;1�R�yy��JA�ٔT�`��$D$�)��r�O[�I�*�
%O��b���!��a�(�r����m�a�����D���OwS"c�@������$˕G!F�h��i��Tb)�Ą^z�	�$F?�T��Q֢OM�1m��y��<�s�4M�W?5��,\,�qзB�L5`�Q� <D� ��*�>z�ԣ�j�{�R!"�=D��٘�` �c$$���h<D�H0�mCWe���S�K�2�R&k,D�,�UB��6 ���n�1ҼCPD D���Ɇ�A�@ģ"�A0I���i�c?D��
� �#rOR���߈Ȫp�c)D��%�!{�][��S(VX,�+m&D����H�vԂ�a�	;MZ��C?D�`��
h�&����L�v�:D��j��^�hY����h8*A��7D�� vm�/����
:"����?D�� �1�F̙͍��� W):D�1cE�?c�>�����%׀�Y��9D����`I>ix�CVn���b饄-D�@	&�^f�HB1�ˌh@^��+D�\{f�4z%��a�j`�v�.D��Y�"��-���A�����٧�>D��z�K>y��p�
F.nz���k=D�X�cja�`��ɹyhx����6D�<�rK5��A�D%>I�3D��Hth��QP�1�֑L] ����%D��s�eæbT�cQԈ*���YTK%D�(�1G]?F��!$�r��Չe�'D�����M�|B�	�Ճ�[�J9B3�#D��:��M�P�u��2� � ��#D�`�Ă60���� h8*�9ţ"D�<�f##�h@f��,m D�d*6D�xb�"N 9�T������� 6D�su�S@����Ee	�y���e$5D����E$�ԙ��ejJl�a5D��2v[�;gX� v%�`bF�q�� D�܃��R�R��rE�'8А���=D��CS�N4i�4�gB�@��<�R�<D�X�����
j&x���t���Q�$D��H���g�Dh`���|�r��'D�,�a�D�}XB	"7���u2zj�$D����=IN��3�ȝ�%�$��!�&D��r�U���_Y�J	��%D��*� ��Dd��qub�F�t �5�6D�Th@BH.���1�[�4���(D�(��;K���Ս\�6^B�b`�!D�t��bרBҎY;q�_-�|11�e3D�(�%&�z��	���9���q�"4D��E�J*$A��� 1p4Xp�/D���㐤|��Q���ڕjD\���*D��#7�AC�|�2���@�f� �B,D���v�Ѡq����\�CUb��6**D��{ŁӵEt��D�]i�h�eF)D�d�s@��O�ν�@D��uX�x L*D��Ѓ,�T�mnY�)o��Go=D�@a�\�\���U�֘߈��b(>D��"�) �l>��c�l��u0D�<娛1i�(�	��N���JF;D�� ����yB���M��h�2�"O�D��hG��0���&��-� "O����lP/!�^%�s%O�3����"O�`3�鞾"`2���m�h�j(�"O���W�	<y�왎6q`��r"O����)&aC2�J#B��i$"OD�'l�5���A�)}��j"OxF��ª}��$j�(|�"O5	!�_�t4�EB�N�m��� �"O����b`(�j0�NL���3"O�̔�8�D��",I
'��"ON�"g"�<N�`tSb�݆]�&P�4"O2��w�˔t2 I��M��K�~��"O��#����Z����MB�l��!:�"O�mHW�8mT�U�Z�s�A��"O�Ubc��x��`ӱ�A/6�y�v"O\4�C���>��҂<�""O@ʇ畤N� ���ȹhdB�0"OZ��!��	Z��3�&[�U<�E��"OHMY��0	)2A�PLX����
f"OL i@�J3\~4\���!r�x��"O�X�t�3����2_�	��"O�x։B�3&V1"��L�*���"O�z�� v�2�k�b>G\咓"O4�Ѣ���$�R!DF�`@�"O6h"b�=#��Y���K/W�,�"OJؐ�#� � nJ.u_u"O�������@�"I�g�F�=��"Ov����ԕ>�T}��'��e1��a�"O��K aH�;�����ƏN1����"Ob�"�%?�P���N���&"O��xP��<aUdU	AHZ	��"O��X���`�r��d��,F��u@%"Od���8�Ҽq� ߋv�x��"O�EC���;_+B "��#z�~�8�"O�����ٔ��Nŋ1����"OƔ��j_>h��9�N��&��"O����hŌh:�G �q��"O
)ѧ��r\|�V�̡����"OV��
�5An��  �
�l� �"O��@J^��pk ])8D�lu"O*��0�%	"���w.ɚ48��"O����83^P��ca��`�"On�jdHK}�jU��b��j��v"O"����]&XY�} ���p��ABF"Ol���6$_�ٚ��X?{��(*OBX�韓8
� �$�Jޤ0	
�'2��������ʧP�R}+�'�ʡ��˂(cT��S�[�?{.���'�na�NɠCu�����981����'|�,]���i��Q���l��h�<y&�"��y����Fl�@��f�<���E�`Q�����U��L�`�<	����+-���������"[�<	t���6�`��E��?���BD��U�<���?��(�LM:;��0C�O�<��̇K?:���&�J� 񈵅HF�<�vn�K �����V��D�կ�h�<�1E�MN�(�f�� �6�Y�&�N�<�M�P�r��y�^5YCZJ�<�G�k�4%�Ǝ�doV�p�_j�<���J3���Ȥo�9�8�H׏�g�<ɇO��T��S��*�JX�<	�!�s(�ۑ�4�!�1NQ{�<� �m#`K[�o��ͩG�:W��=�"O��zt!ɇG��t&Z4)�q�1"O~i:D^�wPh���"j���"O���`]_*�Z�C&�` ��"OR\{��7f��x8�)��1D"OT�r�)��y!4�����9�"O"�	T��.��=�r锁3�T��"O������
��PX�
P���$�"O�,��
�)I��k$� �5��9��"ORe��F,>-:Y�A���M�"O�18جL,2�rG�\6y�~P�$"O4\R�ᐒq����D�Z��i�F"O�������	�5M@ _g�Ze"O@I	S,�4�e[dIԏ`< �£"O�|��c�8��-b�)�(JH���"O���7�P2詃�@Y3x��"OFE��`���ӣgL�*+iha"O�0��L��>\�k�ѪA ��i"O^���͈�r�p�Y��E$0��t�R"OJ��� �/UIP�� Q��&�Ȓ"O��p��aF�mCO\�$�v��U"O2�K��C�e���a�,V	2����"O|�G��F48`wmДB$�1�"O�93t!B%a�j����<#�q�P"O��QH^�-f�`� ��C<	��"O�i�BM�G �Tr�H �� �
c"OH�I�`��=��X�sh}_XA�g"O�(���C�fv�+u�|U,	"O�Lɇ #M�T��% ��
1��"O:�	J�?�����$��b��i�"O�
S�פ!����Ƃ

K>�3�"O�z�]�0�@o��%)����"O�`j����x�\����w�~��f"O�	�p �,���'������"O���Dlۼ.��@�Dn�3��1�"O���� �`��,N��4m	c"O��K��?�z�q��Z�$W:�Z`"O`@�b�\CG�95T�ܙP"O��A2�D)K�F�i�,�bk�Db�"O��p�l�=G�����ʗAqp�"O4H!���;e�
p�$�!hXm�$"Ox�C"�ŦO},$����"���"O>U{QDRB�V�B�^�;�،w"O��`��Hm�؊@���)�Nt#�"O
mc�Pb��@�[�f��Yi0"O��rB"�DȺ��	
����W"O�M{u �4���k ��X�V�@�"O6X�4�_�5�E� D"5L2q[""O>\j��+���ɔ߃Z���t"OD��m_�&������ãw�B "O����E�(�- �N��H\�XG"O�QB�oAW�����J��k�"O�*��A�"YP4�IVEP�	�"O*�DN�8cN���O}�&U��"O䙓����srV@��F�n��]��"O�\����|Z��r*�;|�bQJp"O�J���/�4��萷O7 �%"OJ���K�`�\��D�%2���6"OH���W��&hZ		=>Q��s"O����*mZ��T�ְ:\R�Z�"O��ˢG±G�|�[0f]�T�*-�b"O��x G>��,B�ܺ���h�"OF�f��+�Vv��<OD^t(�"O\���Հ3IKD�B��4�q��4�y
� �l�t��4�����P9]Y�"O^šq�^�Z����� \#B�t�"O���2�9f�����.��W�.U�v"O,��ӧ�y�q�"�L�z��i�"O.��gA�	yt�3�̇ rpP1�"O��8��8�����
���z��/D���冗�1��q��ď�vN�so/D����$XR�J��sE��z���8D���v�.E�Dl�' 
�!a3�7D��	���&��9Y��˅fȩ��?D�`
#���$$�g�J#Y��%��!D�l	��)5�I؃LI�{��x҄�?D���"ǌ�@L�|�q��,gɐX��?D�� �%�X)vܒŅ�&T���+�@!D�Ta�G�XP��#�ދ�>1���=D�(#6    ��   �  �  M  �  +  �5  Q>  �I  �R  �X  *_  ~e  �k  r  Jx  �~  ӄ  �  U�  ��  ۝  �  _�  ��  �  i�  ��  �  ��  ��  [�  ��  -�  2 t � � !  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��I4K 4O����F�L��1d�H�P�2�p�"Oʉ����P+�2�
��������L����46k.��āϔ5���тL̩Py!�Ď::Bn�90(�3�l	ӗ û{t!��8L�f�K�Cx�y��J4-!�䗂K��d萲i�h�����!�LpF`���%_�	��m�!�d��.%鑤�;WF� �BW�:�!��"|.:Q�A%�/~KN�"V�Χ}铎hO�Z��&�n�S�� 8Kh� bQ"O�]�"��T�0%���
LH��e"OF�� ����yU�4�y��"O��E��`��Ǒ�:�>|B��O(��S�v���tn�<N^��A��t�!�D�\
J��ԣ��KV�!GZ=R�!�D����	W�C9!O��!��19z!�d��XMB�oҴRI��&&ͯ T!�$I~�-+t�ŧ	`�I㮈�B!�P��} A���Da��Љq�!�DӤdr� SF!M.Sh,��\�`e!�đ�� x��L/g޶���@YG�x�ɥv�DRt�H��n$�`�ޑc(ZB�	 [c~D�q"�%8�b$r�@��HB�*O��Ah�(�Z�a�tň�;��B�Igh��r���4*1� ��4S��B�I��N@�b�5Wq���S%�U��B�)� �9�wkۑoUJ!²dGtl��%"OL�X�S�TCN�Ba�]�Ql����'��F�O��7W"q�BIīWP\}Ȗ�-(�q��"i���M�>I�\�3ABܘ�ȓm�D��f$�:x&D@�%J�+_���ȓ�&8�@�e��vjĄ0��웍��s�hk�C��]u�$�e��� ע9D� cS"�&@�串V��y+��qv�j�`�	[x����P�� ����O��j��,D�d��I�?�$M�)�'�}� +D���aީM����Ê��2�@�X�*ʓ4��ʧ%O��21nM&-d��#��^T��v��j YA�6����X/�	�ȓk[6�KG�&'o�h1�.O�T92I��x?LĹ���g 9	�	,.n ��2�)[c�� ����N�)J�ȓxJ�=PU��BRܵ`gN̟z�T��=��\�TH^�U��<(D'�zPz��?����~�d��<��ivj�)�H)h�K�Z�'Iў�v2P�AG�>W@���
��L%��D{��,N?�~@j���k�j��#���y�A��Gl�LHC�#��	��FJ��?i�O���
�,+x��,V�:�y�#�J�rm�{r��o(8D�ҠP?��X�L]hY!�dR�o�v�x��K�`-�$ba��^S&Yn^��ࠔ�_��u�&	C�h��ᩰ�&�l�	�m-����Tj��W���-8t#=ن�'����,ʸȐ�A��^������hOq���de�@@(O��PP�I 6��oڮeS���U�&�V���oz\�8�f��1O�扷�~�<O�c��xb$j��M�R�͟+˾��r�?D�\H7Ț���Y��o�|b��!�&>}R�)���F� �x�I�����5$�7V���$'扬&�v�Ƞ�
�v�S@F�'�B�I�n�$E���1ml�p	ïE�A6L�'���3�)�S��,��UhUJ���KY&�FC�	0T�aʧA�%���0�8S{6C�	�%\PX��!ֳG���A ׵tV��Ĥ>I���aϼT �JQ�9����r�79����hO>	P�o��,	�O +��Hp#�/D�`���iE${���3���,��9�O�=�N��,(J6i]� ��"O�X�0Oͷ�P,�ȉn�r�r"O���$:�{a��+I���v�	I>����9AM��f	<Ѹ�
�k#D��pm�:9�	�wd��}>�4Bga��D{��I=r�Y���9j@�t�FF�*3
!�Dº>�	��^�I5�'��7�!�L�D�R�8�l�2G�XZ��*Dv!�[3 ~J�a@`�SU.h3Á�:q!�dƶl��A��j���irA\58!�Ď �(�bv) 9��Ёƈ�i�|RR� lZx��j�JU:�VP�!�B��
k��F/M���I���C(�C�	�Jb�L�kÑ9G�-�0���`lC䉔�6��1���{�nu���&�➌D{J~:S�"[Ծ\#1�@,j������z�<!c#ͳO����E�- �N�~�<��I��`4�SF�'Y��a1�HxX���O<���&ޝH��R�Ћ=(l���'��$S��(O���U��;y���.�� b��D+�S��ۡk��][c�׺I�0	@R�$=��',a|�%A =�d�����tD��*��x��'+֥!!�� V��QH�{9ph���x
� P�P��5U� PpIۘ�n<+C"O��Kp�PEl��@�H]�VI�T"O�T pA��ԛ���,������>����)@�a�`A+�jh۷�>%�!�:78���S/<8^�ڕd� �!�䐢I�N���i��s&<���{Y��	l��~Zc\X�32�|�F%#�
҄_�:���'<��1l]�!�0�
+Y�⠫#R��&���4���yG!Ÿk��-P�)��͘T��1�yr�z�$���������Q��!�~S���<���dLDE�1w�R-g-��B"ĉ!!��O|�b�aV��2�o�l]ĐxR�'�쨘b�]�O�̩2n��N����'����bV�zq�R�%Ĕ��'���z��ܲ(��$"b�6u����O^���>m�J�b�jՉP8uIa`��7�t����<ɶ�A�,I�a*�	�m�i���Pm�<�īQ8}��H��T83�V ɔMC`�<q%�՜D����s	��(!�Y�<�V(	e2�}3��(x)Bt�$V?����pA�\��	S"3�XQ�g�
?O��I]؟��6��$^�v��A!	!%��lз�%D�A�x֮AЕ�q!��Kf8�C�I� >�Q�n#6��P&CH�C�	�0:]���Z;r����H/0����-�ɇFP��ˇ���'��4�E�G�4�ȓVUʰA�C��B� @z�N�-�̄��A��57����͝m��4�DjR�,V���%ߨ�@ Lɲ ��a'��K�
u�ȓ/=����-Q"��93�*Y^���ȓ>��QӰmT�2�MR�^�0|�ȓmfh�riKX*�q�T�Q5�Ш�ȓ^n��Ӱ�cO�pzp�Qb5��FS-�Cd�}�Db�!��TA�ȓ)��a��DL�!��U$p��s�Աǫ��TQ���_�nA������PF��\]f�����uG`�ȓߤsg�[���t1���i�Մȓy ��rg�_���wJD�e
,��� P�ڵiW�A�6\��Y�<��|oX`�Q�Ŏl��S �ʎfr���
$8 !�	X�މkҋC�julͅ�S���O���~]#!烆����+W���CfM��4���W@��� ���&��@��U�rI[�W)Z�ȓCD�� �
�.�����MI�І�[q�ř׫�5Un0��!7����ȓ[��Ka���i�\x��Ϛ/�
8��&&z`2�A
?:�L�z��' |$��
��h*��H5:|b��C�܅ȓ,����&F�%��(���L` ��	4:(�Dg�j���e��A���ȓZ�8�g�ȸn�08�ގ쬹��*m��	�.H$y���	�p4��
�Z���fȸM�H�0F�@#\9���.i�aǘ`1ȁr �%"�~8���6�0A���6�(8����g
2��ȓy��A ����6݁$��3
,���4�Jt��0�1�0�^Gt`��P� |�À��'��T2�s;<<��@jw-^�M��=:���9�Le��X�H�#�*�*�0\�fD}EzQ�ȓX�^���k�`�P���ڍ��E߬����6��0@R�̙w�� ��S�? ���J�'&�`��ġ8L�Z"O0���@#n� ����%fKf��a"O6�S� (y��p�P��9H�D2�"O~���ΊY�y��B��6��"O��K������U�L�C7�,�'�'�B�'�r�'
��'�"�'d��'��𦁝�<t \�2K����@�' ��'��'Tb�'P�'�b�'B����ꚯSkF0��+[��4��'���'���';b�'2�'���'�J,Kb�Ƞ&��0B �*9"HT���'�B�'c2�'n�'�b�'r�'��$��e�5T��D�R�3@HX �'r�'_��'n��'p��'H2�'T4c�a�R�O?�n���4�?��?���?���?1��?y��?)W�[85.��{W��U�ņ���?���?���?���?����?����?قJɝ&JY�p̙�R���l�
�?���?9���?����?I��?���?�Ipe^%�`�S"Z0@��?����?y���?���?a��?��?�@&P�!2��N�ڽY�N��?����?1��?���?����?	��?��/�{A@đÁ�M� }�����?I���?��?Y��?!���?���?9v���j�b�I+I5�B �Q�١�?Q��?I���?����?���?����?!�$P=u5�hPt�BBٰ�̊1�?����?����?���?���IC�f�'1rEQ���́���;�h�B�")��?�-O1��ɪ�M�&��N�Hh���:R'�v��x�')�6M(�i>���)d�[�[���a"	�m�8�צ��M��G�D�!ٴ���ȭ"��� �ڷ��ӠR9����^1���3�Q�S*�c���	YyR�S�lEp$�K��2��O��ơ�ٴ�d,�<A��$%o��N�&P2��d��@G.@�g�<�Ty�	ئe�����嗋:��>O��fcK#fɺ�cC,��F�HP�7O�4��Q=5�Z�%!��|��p�8�A��
�
�8��'��g�Γ��d(�U릕��&<�	�=�����}�s�-͞}��4�?!�[�t��ΦAϓ��ɰ{�Q�d�'3�����\�OV�ɰO�����P��b>A!�	ź��'ި" �ˢ��Q�Ϋ"��[�P�$�'���9O���Zo�� �ejˆ'���3O�l� �H���V�4��؈�kƖ,���A��9JI���O��D~����	�UX71?�sN�x�`��"C�/D?�tB'�u�က�>u(mHL>�(O���O��$�O����O ��c�QR��%/0�a���<Aнi	x����'4��'*�O5r`�V��*�a�S�V�"b^�n8��ě&�g�N�	z���?��+/���`���$� �ɂn�;(�$Q���t���yP�|�&曱��J>���?a1��#��<XtD��J�����?����?����?ͧ��d�ʦ�r��x�T�w�Q�2����OX�k����ƕ�M{���O�-oڦ�M3��i!�,���[�re��(�m¹lD��6|�ő�'��E�>C���+�C��r)�	�?��a���hk�1�� �7�A"�U�E)f�hv�p8��� R
��
dK�U&���/r�r(�4�Ӊ��	j���	=�q��� r�t8AS�16���gؚ�jdP�5:9T�#���E��DJ���Tmqɀ$����!֊&��#Ǜ�>rQ��L��b��b�62y	�0 ��D:��  4��(����*Zx�cs�K��2p�����ч�
[�8�d���q�GMК��6��O��D�O�H��AS�I��	G?92&��Zǭ��=�����TT�!�.�M>y��?1�P������
h���Ԏ#	���`�i�@R�Up�O��O�O��ǨX:��c�-j����'� �;����E��c���IП��	y�&x��첶��)3Z��F�̙F'���`.��O����O�˓�?9��Pdɲ�ޅ��@���ib���D̓�?����?Q(O��)����|*V���.r�\;A�>����o}R�'R�'y�	ٟh�� 6���'4A�����v�<]��&G��'�b�'"X�����'%�t|B�����J7-ڹ&��i��i�b�'��I֟��ɴKW�c?��7�;>����(͗:f ��E�q���O˓�x�[՚�$�'��\c.�@�1*�0�Hd���:q�,��۴���O����O>��s��j��0[�tx��I��%�Z�qR�i�II�K�4e���d����Z�X?Zm	�·��$��HO�{��'��l½��)z�g�	�k�Jq�S.
�A�6�a�oQ�hp7�* tBHm�����ܟ��S����|U���5� ��$�W�����N�D�HߎX��Iϟ,�I�?c�����`��Uu�T�E��>w�Taߴ�?q��?9@�H)��'��'f�uGCX�NeQ1��5?~�)���
�M��������?��	�|�	rQ�6��~�~l3s AQ��4�?Q�i
�e�V�'�R�'+2��~��'���-ܡOw.�3�K��� Q�O|x��:ON�$�O��$�O��Ĥ|�M3D�XR�A.-�0A�LÙvG��þiJ��'��'`��'���O��0oL5]���7EK�=q�#���(����O����O4���O�˧y�x�:�ib����
A�����h�f��w�p����O<���O���<��/t��'E�;����:+ Q�6�F#�z�J�X�0��䟐�	��I&�� ߴ�?�w�� �]˄M��5��A�� ,6���i���'�rZ���	?+������m6��w�Y�m��#�Cai<�m�ן��I�p�	�yNr "ش�?q���?!�'8���e֎~#��c��݌EG�I�B�i�"P�(�	�N�@�i>7��&TN�KpG�?m�օ�(̈q��T���5�ռ�M[���?A���Z�X��#(���ľZk�q�e�i�6M�O��C�m��T��'hq�:H�S�(�0t�g���2�,��p�iN�Q�B�|Ӫ���O �D���'e�ɒB�����O�:�ՠQ_�h�4�(x���d��":�?Y���}DJ 0#V�V���d@�z+�4�?���?��ꂬ&�Ity�'(�DZ�IF�*Tᇙ@����"i�4|����'�⧀��w	�<�O��T�'�"���l���p��s0��ږ��Ib7-�O�<��}}�V����vy���5�iC[�P�P�֌y�<���l�����J����O^�d�O����OL˓z���:�WPX�p����- ��Q�ɫ��Iiy�'��	�h�Iԟ�*�C�\����e4z�9d1w%��?���?����$[t�X�ϧ�@q�"�P�8�R&�f"�'��'q�'��'�Q`�O���H�I5f���E�)��JFT�X�I����	ry�ㅆ_ʲ����d@I�B�<L����2�c"�䦭��C�IП��I���r�$	1~�`DDT)V:"�r4F�Wo�6�'��Z��h�>�ħ�?Y�'1i�e�3�	��d�� ��Y4�xb�' B�à<B�|����R��,��G$E�Ȩ�i��I/�|��ش~��֟T���$�ZU��Fٗ/����-v|�V�'�b��;"�|����Lcʶ$/�/;p!F�^�M��mS ���'���'8��e$��O���/�~�pI0�!� !���B�����q�f�p�\%�"|
�> B����2 s0`��&M?�vi�ӽiS�'�"J��c�L�	g?irB9On��"�ŕ�&�22Ð�M�N>��IU!ŉO�R�'s����ie��a�1���`3o�O�7m�O��҃�_�	ş��	G�i�A��ƃ�]ܔ�+�A��T͢>�ɤ���'l��'�R^�X�֦�C��=c��W�%����X�o���!L<	��?�K>���?1(�����s��2H���#�|.ء�<���?�����$�4["�̧G���*Po ���i̶+4�Q�'$"�'s�'%2�'��U3�'�t�;TgԐHaʖ/��Rø��Th�>1��?���򤙅
�"�$>�EB��(�:l�q㔀��8��\�M;����?1�ia������I;�\)*!��2�������`Ȯ7��O�Ķ<�$T���O���O�\�;��Ƙk{2� �J
(A�n����8�$�O$������/�T?a�p"(��<��)����`/a�Lʓ:��Q`Ҹi��'�?��'Z���=^����q�!`5\�fD�++�7��O��D{���O\�O���`�g�O�6B���6HХ"��i�)���q�"�$�O������1&���-+�:�[Ю+%��=XWM	6~2�(�42�h����S�Ow�EcGh/G���XBd*|
���ފF�����>�M�=�O�%"����r L�"�� ��'S�<�(��d���rpmB���#2�S?�h���l*�~*p	X48D�P�p���nE���5c��V5���iDi<-�|��`ͅ-m�. :�J��,�1RKU��h��l�I���PQNĕ9�I�΃#q�~�zDH�	�8����:oU��R��R�;�ղ�͍{}B����?	��?��'��?I������	����U�̤*�LZX^��	ҁ$pP��@"{�v!����4|f쀑eU�5�.(k!�3*����i������)&�x�*�@�'p�3�J���
UO����.��C�����Θ�LXOx���O�����E�@Ú�b��*�H��88��
<���ά ��%8⣍�Nu�lp�	^y��ڮk��꓁?�(����	W�Du>�3Ȇ���jsH )�h�D�O@��_9����!K۹T%�2��	ߟ�'b�H�ha	�#���Z�iޮ ��Ey��U��ag��M+���� ^޵�f*�ZRj)$*O��(O����'�����Z�n��Q*ߑ8Tp3��}3�D�O���dS�WL,X�T$��
ᮅ�F�VU�҉'�dav�M-�b��PeС8D��j�'(�T ,uӢ�$�O�˧0l�d����?��QI � �&}ў&�VB7J�99�T��'��(0B����4z�N���Ͽ{b�c��,�T ?K��(�o@�WjD5j�{ �`�т�9����'��F���Q>�-h�ꃼ#568�ϊ@������?�F�ir���?�D��!���JuJ	Ȓ��#j�3R^h��?�	�cVn} ��R8j����G���<�ha��t��񟴃�Ѝ|W4�� �����}��B�,��!R�=��䟨��՟X��2�u��'���I�]i�ϠMO ���ӏ�~���\��{�B0��X��I�ЈM�%h-W�4M��([�g���	�v,�9��o�>w���j��'��m��Ȼr�ް0��;k EP�'Cؕ�Q$��ir�r�������S��r��I�fT�\���"O������$M��M�CEB�/� ��T��s�'ZB���D�X��l:� �\�Wn�
M��M�rFE�;�TYy�/�O��d�Ot�Ă�_���OV�.���7�ĘJ�R���Οb��0R���5xp��6$�?��Մ��.���$��">���#��Z, P�0жD@p�Iã^�U�I��	�F@x���)k�j�3K�h��o�6rP����$D�$±��5K�B���\�7ԁ�0D����-��>�tlk�L]��0�p�d�4��/�Ƽ�0�i���'��	s'.4M�*)Dt����`�tEß���� I��?I9t�)7O�(��3�4J��>�y�@G�F��Q�I]3*
\){d�I#p�Jy�C���Nd0w���	s]w�����Үb}�Q�	�\5����S��(O0�K��'f�"}"AE)P�`y�QOӭ-dp� ��r�<�W`� t��g�B#L�8� �l��"O<Y#���(ؐ��gS���p$	�<)��X�uW���'E2R>]�!��<����#kH�B�!s6�ü��yzt�R��D�W��+w[�H*#R���CBQ?%�|��9E�X1�����ۃ'�?����F��*Kl��A m��enZC��>�����Jݡ7��\� �5gVo�ၱ	�O��n�ßT�	x�ƟD�I�H�"J���v1� ӽ��[$�ܟ�	\x�`�w ߪ=�B!"C'�&oPX�a4�I柤p��DȦe���8�D��dI�@����΃����ϟ�Qc��)z0���ɟP�	ߟ�\w�2Oȴ��i��Jˬ� ��)�ڸB�g`�>�Dw�y�CXa���<nќ���� r<��+�_?/��c�+�$Q@nU@�Ō�1�IJ�Ƕ?AR�,���:�D#�!�$BN���&���c�|�I1�����Od0'������'��D��oQ�D�T�A�.2��Y�O���dY�gb���`�;z 4����7�7M���!$�����?�'�R��Ny��s��S3���E��)Rc|�Re �O����M��	��-`���?!��B��	 #�W�V���(�JT�`Q�n�JcT`�
Y�A�4E1��'0������r���psb��QP`�0��Vp��p�j�DL��e
8B����D��B�h�<� ���'E2�q��"k'X��R�R��a��vy��'��O�i�O|�z��_'���p��b"O����@�x�<��sk�0U�z��>O��mZ6�M,O�aXw�ަm��ԟp�O�2D�*у)
�h+E��sz���O<�r�'D�f$\L�!��hhKFD�O��2+��������3%������	�[�r�Y�D
M9���ؠ��B�����:��2�������r�g��(O���f�'2�'��W>�
�N� �X�b���|z����쟼�?E��'{B����U���c��-LĤ|��\Q�'QHR�B�+`Zt�3�.�"�؞'|X�vewӶ���O�'?7l�����?���P���j@Œ�R�x7�Qt	�9�5퇵00l�q3��q�����Ѫn���@�����ƣ\r0j��6��2,]�l�Vo�=MU U ��_��-���"_�Lm���P�F_��>��R?c�T�Rf�5v����b�8�.�#ƪ�O�oZ����O�>�d˲t@���P�.�R#Ӛ{����O����\�@Π�# +3;n����!]��(���������>:{�	�����es�)Kw����O�$pr J%I-��d�O���O؅�;�?��`�"�a��B�{V��f�^S�p�(��2���d���Y1�&��[��dٻb�P�b��K�F�̉�dR-|J!*�)٧a����L�X�Q�$ן�;��d�N�x�83�Я~���
�قa��Ę!���'[�A{�,ˢ ��bc�9F���(	�'n�ٷk�]a8�3��F�j�bp�)��|�M>1��ǁ���H�V`�ı�mZx��|��#)�B�'���'�(����'y�8�fܻ���ndR��ɍ?��Ń3l7���=�DH�Ъ<<O@e������H�.��d�J`C���:cG�B2Z�6�p��
�aK�y�KB2�?Q�p���ϯ8����bI��^�����?�+O^��-�)�W� 	���tG,d��B��~�<�ӮƂm�Qs3�G'jf��eOP�<!ѷio�U��۱�F
�M[��?�/�(�Hל	ME&�X�D�b��0	G��h��ON��><��ᨛ;!�EpU�Ҧ��OZ*	�VQ�:ۼDzd�6R�b�Ez"� ��L�S�.M�Y;b�;��V0s����T|�U����3e��-��aS��I6t�\���Ʀ]�O|2���ș!u!�s�z iƁ���d�:��������͌hŶ�	F+6F+�)R#�N{�I���O"TnZ��M[��!���N��;�n!��mȦ�&�͓g��1¹i|��'v�ӹPǊ���ܟ��I�At�)1��3�X̳�,]�i�`xV�Q�Qȼ�j󉌥� ���S����'ΰ{��B'\��E��LŰaE�����ǌU5؂��O?�d�8VsdL����Qwq��0]t�k5��O �oZ�M���͈��\%e�$�'a�+]�
YqD�E)�yr�':�}���äN��T4A$�H;�O:�Fz�W>�
TaZ��R��
��/vh<� ,�4C�>m����+j.�۱"O���ǧ�ɬh�dϜ�ZP��H"O��A�ז�p�Z��e
X��"Orغ��959V1J�l�N�LAf"OL�A�l��%���B�^>hS�`��"Ob�I���W�:�ɀ��Ok� +`"O��.�:k�x Ո������"O>�`��2e����vm�9"1��"O:�2���0ezaZ��U�@e�u"O� e��.cѲ�z�YU�~��"OHU��� ��L��,S�a���i""O���c�ּ12dq%K�%�| ٓ"O:=Ju�@�gj���ꐪ9�`ж"O��a�.�>p��8e�۩�F�	�"O��b�	��.����4�����E �"O�����/A/dd3G嚦�̡��"O�p���B�xA>��!ń����"O�%�v�R���b��ܵC�p��"O�<�&�̰(g�@��
οrL��"O��`��Ҍ�<ɱ	F M:z�"O"�$�� X ��C��f1F�I�"O���癀z]ƽHD�BPd�(0"O��4�6Ǣ�pb(
�s]���"O����S�*��k&'�=>��R3"O�]$h�<�4����O���"Oj`�Q#��eA�:���<a��{�"O�$�A�E�|�@g[; ��h�"O��JD/�$!X�k�)d�.���"O^�35+�skt]��kE�w�Nh��"OX�2W�D�_4,�K�J�%_>5��"O�� ��:K���Є��\8�L"q�i������l*�m31��Jb�����E+�џ��'�(��O~
ş�Ut<����T��H����f�<I�k�71��t !$޸4�&%��M�f}ү(�MK�eB�JX�)ҧ;�r�0����lW���IQ�l\J`�ȓ{��MYSa^3Y��Cc��|�]��cܴ�Mk"cR9Hb����F}B�ڂF��i��9������Ȱ=��(W��=���E��I�$	�U��0֎��M��M�3(O�$ʒ1��I6 ��`�V.���!�#A�E�@b��JeAPY ���K�,�J*�H6�_-d	�,��kD�5�B=�5 %y!���*/>�x��7v�I��,8`����S��xya���LN��>�����0�r�A�0t�
�j5�E�<i�cJ�Tp�C��O�L�AT�G�M���.4��镁�#x��*Ó|�j�Y�)��B׺@��`��0N�}��I7h�rΙ�OyhԀ����.4ZwB�S��D�f��W>܀�'�v�cv*��$�:L���]P� I�{b��h�%������%��iBE.H�²W?M{ �%di�̰֭J��L�h"k2D����S�Q{�^�M��R5c�!���2�	���ؠ�A+Q���R���BŬ�y��˄�|,�# �t��x�����>��'�&�
��*T��B��Zn�=���� ���:O|��ɃY�j�	��
'�b��Kt@Ca�ּslB����3�HO��2��A����wc�v!�P��'��]����(�l騁�UX��Dv���,�&���^^����'
�LA�K�KԀ�#����^~$�ݴiH�|�t�
�:d�0��ß�V!m'��]0h��3Ђ�x�$Y�!�E�`i{�e�<a#� +�TQ�g�O4I��y#�O�v�����
Jp��"�/��hS�w�`$���$9Z�A3�J��&9J�j��� 4RO�5�U�F#,��XA �jf���S˄{��h;b��S�)ev΀�r�!g���T�\1�jb��aa���Ty�x�D��c*����OY
'm�X��`NԱ2R�C�|�<y�SÒU^ a�'؎�!5N�$V}N�5rk�����<c�H`��Q����P�Bƈ���5���僆'���4QX����\~R�xJ?�� l5>����'o@�ZVh1��j] o�a{R��Hf!�*� ��A'�	��(��Z�S�.�s)��`F}�O�vP�hrI��~͢�A��
2^Հ�N�67਴&l��O*�K�u���{S�m������(}�d�c�Z;thP�0%�B�^�b���i;�Dƥ���(E�Ö=�Ti��Y&�O� .m���'
4�V�^�4�,����6+O�q�6MX%�$K��B_J�f��/�&	h���>�'K@�Q�mA9���?����T=%\�0��Hk>*����'&�ș�Ώ�7���$���P2��eʟ���P�*[� �D5�NN�<�s�^扈f���=�D<c�\`}�|���=q2>����7/�l�!�[�]*�=��D#���xcKIĚ D�ԠA<N��l�`��4A�6` �|*���uG�y>7��0��/�mqf�[���R��9�U�>�	G{��`dIG>hb��B��q$�O2tz6aȫ �>M�� K�B$�E�J<�Dc� H����'{L¢i�5֦ 8V�'u��%H�ϜLZ��Xea���pP#`N��H�ם)�X����li2L٧fӦ9Cr�+-~!�d�p
����"�T����N[s�v�	�h��"�J3���<1Ӷ��(�@ꖚH �M'�(�@)��-!fA)�%�EL`	�A]���Z�� @��ՂF�i��\��o�n���R��R�V�Jq��c˥,|����bEL,kI<E��LƋW�B�)2K�f|�j���0��'ܽ"H��wo�� Wl��gL���O�^�Jgŏ6!H������8�j0@ H�4��i�L�~�>̂�#D �@�g�']�ʣK�z�*$��CP�HXR�y�mJ�|:��R��Ԉ�-ռ���S֧����;��`C�L��=��R�Z��7!� v�������~�h�R;��h���]�	=:U�e�'(�E�ᓽ��@X��W(a(�1+Q�m$\t#s�z�A��I�j��i!��M�,��#�)zj��$MW�6�r�x�)��%�r�F����<�A��|j��C>;˄�0aH_�Q����'DB]_��*�!��k�Z��':���Q�S03W��7B�Qv�I��O�9O���-4@ �b	�(b�e���2`��%x#�Hy�$��?9.X)'͂!S!\�:!	�g?�L�犅1R,0�M~��������@�-�G��3]������jlRL�":�=��	⼃�b��- S󯅈-�!h�A��<�V	�u�O���؃�j�%"��hd�#h)X��C���w��G~��U`{@I�B�<2=ԽY����M��O��h�L��Ơ#�꽲�C�pyh��[��'�.DaZ>�ya��"!Q�6�.h��D##�$v��D��9)�	�X��!����R6΀J�M�Ţ�S���r�)%.��<c�E��!X(S4�`�'�sAߧ !L�b�A���J�Ɉ��»v�P����IUv�L��B� 0.�i իJ<���'�`�3��~ڦ�^�.��Y"���ht Y�&��-�����2�Zx��I�y�b�7�P���J,� �!�m���MS�� ��O�>��Yw9��`���Z���eKt8<K����?i���m�:Y���I�\^���'0�I`�/��I��x��)4��D�8��M�H>��V>��@�C,(r���ʚ|3�Y�֤*|Y£O^�Aq���fM�Q��>=rz�m]�Y^,�S�ܴE��C��2�J�	����#��'�´��Jw�"=��R>��1Y����̮K�@䘆�8"�p��eD
����pT�)��m�R�g≖U�L��"�o�JqS`��&�n��b���sF��2�E�nQi���y��ʫ} �l�jV��&a	T﮽x�	�'rM���b]��݉S ]D��j�um"���JZB��y���0<i�_������+���K�o�|2�(F�Y*�"=�V��d���� 4���� �3*UZ<様OH�D�G4k��a�dV
<���)®��|�!+O�Aiǯ�r��2��:x�X!���O�����
ֻ ٦�����&V;�8�T�:��ɇ�M�C=v�腁�&P�)���Fx®J�Z��E�Ӱmڢp���M�ol�%+�m�:T�I�|�|���?�(���'_�)P�	�',D|�"HYf
̴�m���C򌕨�ay�&�����Qj�	l��I�Έ	����ʌ_%��'��ڵ�?9���)2B�5a2�?�'jk �aUO�HƼa#pI�3��1E~H�:*�A0��� �҆��MK5`];~���T(��E�q�ꦭi��q�|(���7�t�"e���dp�����<1�8ҧF�:Q����b�>�!�ub�ыfϏ�T�FX�I���M����/'|�@@#��D%< �#G�p�pƏ$tbx,��I�!�p�3�L�~�2�J��-�B��&7{��U�7%�˟���"Tl~�W>m���. i�a��s N,�fK��_�JT�F�'Q\B֊�%>rٙ�A�<NR �:f	�����t~bQ�,���4Lr�p��O�2��O��aƎHL�]���8�F|���,s��A`V�҇}���#0�,�y�m�6�X�ӓ��}�x���-�����0J�&n^�6͆�-�൓���+Il���� ���C���8Ɯ�F� 4���'��3��v�����kG�*��X�� ��m����0EC�h;v��a�%M�И�28M��xD�$3��DA	Z l���NдL��L0�F_Q�����&}XAt�ީ;t�KФ]i�ak��'R��-��p��$C�u����@�J�7���D�&R�"���ܶ�f�q�dܐ���1Lܷc�2}	����fc��m�	 b�)��[\3�7��z��I��h��p��և2�2�FxR�Lt���l]�5�k�}7>��
�1qb�"2�D�%�'����'���"j�$8غ�/����:�'�v�PH<���
a<d�AtO�c�2��@�;J���K�8 $�9b !=�����	�y��U�GDN5�Э�ւ��iꜱ��cJ58��U�3�i^JP��8�y
� ����s�(@��ڄR��M�5

���|2��ȼգW�ȥ�PA�,VL��6'ƻT5����O�Y3%'˼\gB��+�>�����gR��pE�סz���Aӯ1"Y�A��D�P.��8Po�D�E���kp(V)hs$H�O�>	���J�G\��$���&��Fb��2O2?��H��rT���݄Q&�t�B�<9� W�OK�L�mB��,U��Xz�'G�\z�ҧ,�t�8T�K����q,߅K \�G���t�J��0<!�O�71tu#�+�"t  x@e��#!�zKGWX�`� �A��y�	O+b��C�e_<���hS�Q�v��IE����y���	�*C1HY$蛑
������զ}1V�N�Er0-R'(�1� �2U��-	R�{f�u�'jd�6.�&j��!I�!;O4��'���X�W�u���A��;7C�aB��d�O������~k>�@�ʡ7�1���'k�}5+I6�&��3K�nI�͒�2O�e��f�y3�,㒌�i��|1�ɡy=;��\8B0�Ձ�-V=���0`I�mK�\�� 90G��'���Ex�/u��$(�ߠ_=�GN��[���S3D]�BA�'|џ�S�'_�qVRA�kӷ1���ђ�	��Tc-1?6��$�S�M�Z8����X%�p�8A#m<W�]�Ƙ9�$Ba���{�kV���!D�Lcӈ	!qmγ3J�
QQ"#L�Q�FK@�V(��*X�	�𱺖�-ʓ�~�� ��j$ͤ%xX\KԎ� v�:-� �;q���� D`m,1b�>QEk�|@�Zf�L�%��!�d/�u�r���3�˥D<k�'Y�*oH�"�0O�]HPHГ��D����˺c0J�P�':�s1-e�i�d�^�����K@WS�0R��ɰ�O�ܴ��Ο����H�	욼��j]hX��E��ȈśĦ�y.���4��;�I�KPv��rː�Ȅ���Ā-P3ȅ�Ԯ�cԁ��M��<�ǁS<H�ޙ��o�. ��$��M�@����>�4qkYl���!N�<��MʂLދP�:t�̓��$����ȄlH�
�'P<����I���OȞ��WǢ���GC4�Q�O�����(�.��ɓ?t��Z�X�Dק:��F�5��aQf)�ov�筇{�<Q	SXfD� �g��N���a&a�u0$�aN�(�f�I���~����>zL��>�2�Hř�yc�T᳉��	P��'U d��"ZHZ��u$0"����^o�
���4}6.A� �'-��v�˵k�<tC5ǖs�6�����ˍnW�����L�O�����%�{��pk��bW����'1����������8@C`�RtJ�'oX��W@��Mp��0�C�&�Ph{�'c�SC�I�h���¤ �,�bA`�'3f����.B�<!4�˜	�*�8�'��!Q��Kf-|9��j��}�DE*�'���م�>.�~MxFNM,L�$��'��I#��Q'����6��O���'rlt1���o��q�� J��	�'��[T�M~�E���C�vt����'N���t�T��J`��k�f�8�'�A��G�I���� 3�8s
�'����f�R
J�n��aLLm^��
�' ��9DG�+,��!��kk�4
�'�� �0� 
g���*,p����'��'
�+���Ւq�>�	�'�hL��N��\ ��T )����'�=���N�'�=�wNUEǒl�'ݰ�d��Ňy#Hٻ����y�NX1N����i�1"��=����yҠ���X0� �Ȩ1��"��y��u�@ �U�P�T$��p�A	�yJ�p�����Z'��P'X1�y�DR>`S� ɂAU;@]�0����y�H�3c�-����#'Ц|`�O��y��A�]i�l{����F���T*ǳ�yR��,�u#�?s���W*\��yr�	�� �	�*T��;WHH��yҍ?Xx$<��3k���c�O�>�y��ΡW*��%�F�j��|󵢏��yM��?f�ͻ�'ƀ.���4�Y��yb�ХrK2̂3�I=t�֨rG�\�yrn��y���`��>�Ȁ���4�y
� 4\�d���DA�9 � �>톸�A"O,h�D�9*�J��hߜ�8Y�"OJ�(�$J�9��4p!�_�SԜ=�""O����LüZ�:�3�?*�%A"O0��SfI�&�%(-p���"Oia�O�8��di7F�/<�"O�U�E)L�G����q�ԿGԨ�"O��.�>��]�t:x���a"OXT1�o�"DL�M8	�X0c"O�a��N�x��	�S�[�A�ʙ`"O�X�)�[��Q�H�))Ȭ���"O�p@�͏l��t� ��I����"OVa�DC7Oϖ�*���<#�f]�"OzDx�f�:��(��C~C���"O�lp�`k>AX�#ؠA�p#s"O敻,V��S�B]�=��ң"O��P5�Z�T9�g˓1����A"OJ��&-��V���h��:�"O�:W(��W*��n  �8�{"O�<#��������dL�i֜PZF"O6����"tx�+�ɷl��H�%"ON=5xT@,3�N�������"O��(�C%S�P�8%�J-�9�"O�,@�ӎ^�&��7[�7$��3"O
I ��ȼg�Fu�q ��A+�"O��5 ��>B���O��D;L�"O2�jDNdj�r��Ҳ^(��"O
t82-O R6T��L=���(A"O�|Q"6H�f�*2�Q!�"Oܔ��]�N�J�2Ŭ�q�	��"O���'?\��4����*r���5"O�)R"�N~N"A�]:{R���W"O\�S7
�'�����~'�Yj�"O�Ԃ�#N7T�<r�+>���"O<}D���o�P;��P�_�օ
R"O\��ak� EU$0(2'_�����'D���c��	�YSJ؝Vh����� D���e�!lN���־v	��P@i>D�� �F��0���b��v
L�z��;D��� F�):�&쉰���-c@8��=D�$*rb�,C�
q(bF>�lD
q�7��l��I1�%�E-�ye��aՀF��\C�	?�����C+'X�����=)��?Q��)@�i�J�b$g�����)�=!�4d��xd���	֦�@��E"c�!��;����e���,<�JRu�!���($�%��kE�
� 1�GCt�!�dL��)���-i~8BF� <^�!�DHk�V�R��B�@��nȃ`�!�D��X�*��ēV�$���휙U!�E[�$�r$��{��#A瑻n!�$����igB�"p���To�L!�ԡN�Q��ѫFf^� ���j-!�[�G��i �i��?��}!,.t+!��C��]Y@ē�"���هJ�!�$���}��E�_c ��To�f�!��A;l�д��.�27G$����,0!�d�%_�4���'ܧZ ,��ت; !���?�|��'ˏ?��p��k�!�$����{\I�rIHv@�,}���G�P ��D�  K-����ȓWר��W�6�h88� ��Z���QX�5`�A
-;fdBvN	B, `�"O��@7|�̓@m	*��U��"O� JPyda�� T`��?.�2�"O\�#fFL  x�S+Y6$�I�"Op���o�@��p� �K<i��"O"�ӡ�	�L� ��-�d��"O4�Ɖ��V�GOŦ��(2u"O�H J^:-�QS�� *�}B "O2�@�ś ��[��8�l,�R"O��i�#��%htp�M������2"O��A��t��9�a-�$z�h��S"Oh������]YaM�'�����"O�%�Si�8@���m�-~�M�"OBdsr�_�.�|���os�!�"OL8I� ]1j��ѺU,��o���p"OZ��
l����ciZ�JX�U"ON�B2'��`�A���lAo(D�� te�9@p��0 M�xCf��� D���t�]�Olщ�'��6 �2'$D�6�!B��"�H�#x2l�s
o�<����D��P���R1��%��NC�<��F�	��s�`>2��
���~�<���'6F�Q��tE4A�Wz��D{���6v�N0xdm�V�8� ��y�g�n.�رg	��a`�E���y�h��� �1�,�>�p�.X�y�\%%[PD�D�ݑ䢜�@��y��=J��:j�8�>���bO��y�/[);Y�ܠ��[�biz���.ڻ�yr�<h�z��"�Ǹ$)P����)�y���x���z1@���x�B��)�y�D�7{����h� �㑦��y��Q %7�x�%���~����y"B�'��Hb$g��t@�k��y2�L�����G�q��Q�ܪ��'����'1HA��JP_��tR1ć�9亰��'L<Cu��U�J(B6휼ZA�Q"�'h���ڎ�F�%�ܨ{�Lm	�'���r��lZ���C�x�a�'�-9��O%)����sM�"c:1[�'��q(Ѵ]�2	@)̍':�x�'q�p���KĘ`�J �
�X���'�\!�&f�@���Z���L��'8��@�20�8$8�!9||X�)�'А��m[�E�N��b�\�nw4�Y�'�Zy�C�Fj�ΰ�M]�k��\��'�\Q�Ug٧X���c� ��'3�����7Q����A6�kڴ�Px"#@�Vr�:���?r��C�I��C R���"�+�8�P��$D�h��
J��P0fiK3(��[�l/D��CQ�֞b��|XfɃ9@ԡ��m:D�|�ckJ��*E�d�>�YD�:D��P�R4P�:\�B��Dn�{��8D���͍����-�r\Pbq�8D���s	�3B˲ț$A	ZH�A%N5D������$oD�1���&n�n	Q�(D��K�!?z4h)���;}e\!(��'D��� J�!�|x��c�K��Y��"D�XZ���	���X �����h�f.D�,�F��)]��QJ	0P�1���+D�ȲU��\tő�)B?Jc�}c�%D�����b���`S&B)2��CK�>I��)�'!��|Q�	��<��K���=Sybm���Z��A��D���3 �KT�α�ȓ@�6��^�Ĭܣ򬊴��D��S�? �P�qn� �E��o�,o�0�a"OR<�����=�~`�c�vi"��'"O0��K��{����CE
s'��� �+LOD��s�K�8 �̋%{�
�"O<�9����<����J#�@"O�=����C���"��
X	��ҷ"OڤJP�v"a������"O��ee�R~�$�6�A-#�Z�x�R�pG{���\=�4��G�Cr`'�αZu!���<����)m��VR�g��D�#��U4T]�}���Ιa
h�ȓ5��을$�zE`cl�:Յ�ogP�(�%�f��8 `D�	��F{��'B�5�!�sY��AqA�s�b�;�'F�i��Нv���P��X�l��}��'WʸC�W���q�ăd ����'�@��ǩ� ���,��g��i��'^~�g�ۋ�1����65E<���<,O����H�vA��G��K=(ܨ"O���C�Ŷ0h���!֐X���@"O|	BW�fA�kc`�N��D2"Ol��������`�O
Z�8@�"O��`5c7wv�I�D��2U�yQ"O��p6!�6��!�����jD��"O���%!Z�]P&C�%U��}C4"O�0��E��6ul�r7� 'S�JHCu"O�u⢪S7*�>B3�K5Pw�ɀ�"O8���ч-�<�M>(r"�D"O�i��DT�*E��{�̛8[���"O��{�^}�Pٕ�P@s$��@�'��I3
��X[�π�MǤ���Ȍ6pp�C�	&n�(�ed�3e����@<6W�C�% ���B�� %&���d�_^C�I�'H69Ҧ��.�)��h܆XV�C�ɵN+Z�fQ�]��e�+Z9��C�I�{�Z�Z�k.L�!6X�C�I�/��a��)yL��OÐ,�B��,I<��D9*�<��a��]`6B�I�mzĊ4)�b����i0B�I�IzN�*5�<$2x�R"(�&B�	-��U�0��0g&��q�=.*�B�	#j�t��M�-�XYu��&v�B�ɪZ���Xb*��*іĘF� P�zB�	���d3�N��xx�6o�H~C��$�%��+0B�ە�OD hC�I�w�ve2�i�-~^���FM�YZC�ɵO
�D�glE'nM����/kn2C�	%Pm 2R�R�����ɁH�ZB�I"��m�4C[3q��U*��ӆ$�B�ɑ$���2ϝ�Ta:��';W�C�	�X�´��"�V'x��Ǆ��A0�C�!k��@����O<r�J�
̹n�C�I 280�	3�8?2�X�#�� TC�	"x�� {�j�0f�Y�!,�+��C�ɐco��t�S�6�����CAҮC�I�8�\�CS�
��x%@ߔ!;�C�ɻ>��J�R�S�C�J�fgC�I$D0��-�x�ˠ�<�.B䉓]%�1�+�^h�LZ1UB䉀Q`�qO9tY�E���j��C�	�W���cQ�X�)�҉2�i�
]�C�	���1�'@t/��&e��	o�C�	0T8�a)�'�Q��w��#��C�	5�x�Q�5%1���D\�h��B�)� "@Bu�7>�
U�M'���1"O���8+�90aA�*�����"O�����ø��PÁ�"L�ЊG"O U#�e�s��sç)B�����"O<�� $�-٧�Ê}ڤ�"O<�@e�N?:^�HdHĴ
�|p)�"O|1�Ę
!���Ƃ�*�h4#"O��(�C��q=�s�CY"N�钥"O �k���D�Պ �,�CS"O�i`g��pj�d�GO�V��HQ�"O(P������j���+cD�j"O^�`�0��sueɠGG�"OXDP7D7ܖ)juE�`,l�G"O��8j�"�
�[R��3�!�"Od��PNΈ}Ap�@�שCh���"O�mR��]P%&�k��!x�<l�"O�� ���v�9[A��$V^ܰt"O�5*�ڱ\�p�*�v]���"OJ�a!�U����s�C�&��"O�$�E���H�^~ؤX�CU�<��ԥj,��R���D�~�"��P�<q3��y�Mk���,#�T�ڴ��I�<A�E9Sx9���A�0M�f�P}�<q�h�/b}�E ��@�O�����RO�<QƧ%8���:�P�ְЃ��_�<Yd�A��H�CAE@������\�<y���.[�� Y�쁓r�ܑ�.s�<�@�ǓvZ� �9T�咶DH�<�dAK9a���� M3A��D�^�<�^�2I��/�),����T�<�  �iu
,���M
&E5��,�g�<a)O�'�Ĺ"ÆG�����q��c�<��J<���W�F9j}����f�<Q���k�):
ԇI���K�._�<�Â]W�9s��F�}�p��s�<�F�\<�B���/�h��`�kS{�<��N��W�U��˗�_�����`�<�E��]4؀����944 �g�\�<1ugԠ>��[CɗF3��"$��V�<�6�[+*Fp1�8l0u���V�<�s�4=�SAǵ�&�ʃ"�U�<�B�ǒZ�JI��G4;�I
rh�u�<���U%fqB���.u�5z��Mj�<r�L�Q�聠��M6tA��f�<!s&�UO$�3�ҽ8���4k�x�<���Ė7�,6bW(Pf�[L�<YBGI�!%x}���2@
�@�/QN�<�eD�%J;d҆�8�"h�"�@�<��-/?��rbVŲcD�<�0��.6�&thah�x���V��|�<!u	F�`|=b$�F�>�	sGq�<MIi�I�N�*,z�%p�<S*�O��X���4	w>X�w��w�<q��>:\���W�KN�]�P�o�<�g���qA�O�d]pQ"d�<�(3s&^�h��X/**��1��]�<�T�4^^0y�i�?oCrU�j�P�<��ԡ�`1&�\V\��K�<Y2�[�$�XUQ�C�����e�L�<1P���WèX	c���9�F��I�<is!��_T�`k�`� ��LX'��D�<��e�kk� 8FI^�A$U����|�<��ګjpf$*e��u�^i���w�<�́5v�04�4�Y�nTaH��~�<� �Ԙ����u�0��+2��"OF�����h�b��Q<$�q%"O��P�l�nP���W��`-�XYu"O����
�5锼	B��SuzB"O��Jؓ}�	@e G�c��H4"O��"��-��4  (B?H
�"Or�Q��k\� �,K|5��"OT(�m��c���M�3���۲"O�5j��1r񑷋��H�0�"ONt"�'�%?%\�2���*t&�@P�"O:<�$�&�\�s7#?G��M�D"OqqG�X�`y��
Q���$"O�9�jZ��`�9c�}��2"Oʴ�p(��j��@�5*͢%� �W"O"�jtȻ*����1��q!"O�l�`!�c��H��ˋAn�Yp"O���0Iۣ� ��`+Ƞg����"OZqi�nN�H��A�W���F�N��'"O�,��̨ ��
����yc"O�d:s�a��K�-S��!86"OX�y&J�x����&m ���"OX5�ek
b�� �-M��
�J "O\51`�K'w �`�B�]�F���"O�����V�4	��蕖h^`"O��Q�/>aD0�a�|Jް��"O��kt��5z�Jm�!��04����"O�Q�5}l ��������0�"O���6���͹w��G,����"O.D1�N	 qo�1Q���q"�8�"O~L��C^[E�(�eb8~
b8�e"Ol�����,hS����ʪ .��t"O�`F�Ǌ1b�!�D�P�e��p�6"O�(�e����t�+�_��F��v"O�,y���EWV�9�I)�4H�$"O�ذ� 6���;P��%Zj�8�"OPݡ'%�.�P �c �Sel0"OНy�,n����6����(\�"O~؊@^�Y�¼A��
v�z�b"O�x�Q�׋r���QQ`��ܭ3"OF|HС�U�\���0|�t"O��(�����^�6yC"O��9�g9,v-(�K��ar�j"OLq[%CX�~��p �(�1���C"O���L1
�{��M9�Y��"O}�Pݟ: 4����"?�H-XD"O�M�0��q�|����F'6HݠQ"O�R��۝r�h�T�&���t"O��Bł7�(�gC�*t��"O`���Ə�ct��`��a�Fe8U"O,,����t@T��^�eP�"O�9�/����`�,8@i�0�"O^l#R�A ~��댬VY
�"OF���/T�Rǎ�
���6G�`�"O|	3 �%�tq���$*>��x�"O��{Fe@W���Ԇ�9:'*t�%"O8Y�&�S5m܄t:���S&"�	Q"OX�Bvh̹Db�"�l�'H��YA"O���#W�"�Q�@�֗��h"O.y���̯T7��ѧjD�7��D�u"O���gՐ9�6T��(_����r�"O��Id�
���9�e@�:a�l۷"O�-y4��M-�1g�
J4z�c"O�
�OK�5hMiE&U��X��"O�����K(	�P%�`��<4�1"O� ���@�&>2=ϊ�]��p�"O@�x� >Ed0xq�S�)��[v"O�\rV���T%K����,!"O ��W�8g�p�'k��J�[b"O`i��L	=3�z��$�΃~�2P�g"O�D��*�+9��yY3��6
wԸ��"O��$,`|M���_-~�1��"O��
�G�?H��#SΔ�Ub��%"O��
5��=k��0�k̷p螀JV"O�}�5
_ ��v��q�Dpy�"OR� �)�i�e���F�@�L�ˀ"O:�pb��Yp~`�e�C�>�̐��"Oܵid��P�|aBoW^����"O$@��E�/?�^����V*)�n��"OH�1��_7���#Bq���"O��bU��O�x<ipCʑj6����"Oxs��B:;r1c�GԻ<�����"O܉��	R��4�&GO�z�.�q�"O�`W@�$ 2�C�Ƚ$M��"O������N6��q ؃I�@3�"O �����F*��doČ$���"O�42fXbd�)ֈ�"��u�"O�497��v��Ś�D�� ��e"O�N�}� ���Y:�2�0�"O�X�ѠL	UB�`抅%y��� "OF�Ӎ��J\٦�ł6wN��D"O�`sV�=�TH�C�`�q��"O�E0�M����L/8Y<�"O��;6A�|�X��L�`�&�j"Oȥ;�LÚh�Jܠ2�С�|�Sc"ONL��Ĝ9"p�@��B�da*���"O��i�i�a0LJ����E"O����΃�}*����:
�hS"O8��D���,� kߎ���Y�"O:-�2�[�Z�R���Y�A��)Z�"O�����|̀��!(�5Mx�ȋ�"O��0��^�F�z��I�ONBP��"Of�Ȧ�ڬm�>�1)J�b3��"O�H	F鍮P������B+p/ �k�"O5�$���iqqo�X=�"O��æ�ͣU����NųhpD̛�"O��R�$ѯ)G�(�u�)=M^�V"O|����D�@�a��'�V2 ���"On��p%/m�SҤ�9}?�	"Od��W�'28��H4P�ȋu"OL��� Y���5b@�O@�54"Oą(х��_�0��!v)�Q�d"O��6�C�L	��
�&\�=l���"O�#�U�7E��d@ !�$D��륌Ƣ7�b�����`k�$@(D���,Ǯ.N��$eU��)��%%D��C���-\��AJ�B\Ѕ:��/D�d�Q��0��a�d��Y���,D�̂`b�*��J`}��4�I&D�x�e�8֌}��L���,�(D���&c�%�l���|�x�� .2D�̫jB������JB8�S�.D�Щ�O^#3��a�Ă�U+@����,D��t���b��y�B��hB9�V�*D��3�H��\q��	�8�	d*>D�|��
>l�(7拸N�4��CA(D��x�BW� ���Q��CV���"D����&�9Iw!8VR)!A	#D��g�ʑ~N�8r�i��d���1�n"D�� ���&��*m�ڱ�I;Qrꥻ�"O��������Y eV�!y1"O2p���E�k>�QS7�M�E�q��"O�=#WmL7MHxnR97��3"O*��`G�	_��#%M��pU"O�c���pŲI�5̙�M���s�"O΄V�K��`�8����er���q"Oc��E�Ft*��ܔ9}>��S"O:Ը�߶JdA�R��#`d]��"O~�{j�=W��	3t!��I��X�"O�$�� /�֔ڶ�H���G"O�	kG�E�WQ��#4�T�ce��B�"O�yySk͵�
D�B/S?�`�[�"O��覍�$���YѬ϶<�`�ڢ"O�C��xG̀��Ԃ��"O�`fdYz��(�)�0��i�"O|�J��_�=6Հ�h� O�1"ON�변�'�HL2dgQ�g2��"O�t� ��{���&G�-�l�T"O��WM�;=����eZ��ks"O�}�v�"���j��\�}�p���"O�CA�^/Bx����$^Ys���c"O�i�e/�:�eb���/U��<P"O�h�D ܔBOFiF�Y; ��@B"O��äN7'�AZ��N�WWF�8w"O�ɚŌ)��y7�̂Xڞ�1�"O�8[HE�gk��жL��x��xB�"OPi*>\T�&��"�PQ"ON �Tg�sR*�i�+̈́+��, �"O�	�5���S=����,+��0
�"O4�`"ƽ9r�qE��o��e��"O L��$"���g%�2%@��"OT�"�4`��`��#�6V=1�"O�M� kܖ䬜8 �:\ \��S"O|0�����%��DMn��(�"O@@�d�L�1�>��vĀ�s~�y"�"Ozpƫ��LU������=�"O$�D��&��3���L���"OFū%%أ5���Y��Y�<B�C"O�	� �p�\]�$#�� U"O���%�J�.��1Z�a� ] M+�"O��s���n�BTaD $%��P!"O"lH�W�X�^��bov��c�"O�P[�˄�+`�0�.�~����"ON�"#�X�g���8gm��� R"OT�����/S0���&�+A�0�i�"O�)`�S�JY�`�Ц^�>-����"O�( ���-��5г���[�C%"Ox���A޶m�Oٿ ���#"O�Ĳ��T*�R�����S"O�1uϔFc,ի��Y��p�C"OR��J��A���a4��2(�<�H "O�Y�T��C��X�W��?T��4"O�u�Sg�, 0�6O�(E6�q)6"O����7.kjأ��%G�T�"O=1�ڛL�>�k���(9`lA "O"Ȍ":���b`-��v�LҴ"OZ<�3�]�J�t-k�EZ8iX!��"O��Ô�.����+UT�-1�"OT�!�m��VPX�銵I$"8Y�"OHXefO,&.���K0~�5"O�1H�1�>�Ia�P�!T�b "Ot���?D�hatF�#��ݰ�"O"�C��1���I���bm�\�"O� ��r�_,:9J���TizQ"O���iH(>��=��_�x��q"O�l�q�)�5��aM�p����n?D�tBH�1"�"����8���tb=D�����ɽIE�0�W#O�^Z+�C6D��ȣΙS3|!�w�b~*� �(6D����ߙP_�MC5*�w6�� K7D�D��BX�]��
!h�ҀH+D� �s"D�y���рd!�s)D���R�	mfhГ�h�3H6���#G'D�{Q��2#9E���H�0�R�-0D�á��}�~�3$BD��x��l D���o�p�BPjb�;u��P�%>D��9��H�r@F�P�Dx��<��l�����<�x��
̈v���ȓ[�9Kg�Ϯ!*�T`4A;j+�ZMByjB+�����Svӏ{ �A�ȓF̈́�r��'L8y�f�5�Z���#+Vd�����yx��bᓆzu���ȓ9$�y�Af��h�\0 �B2n���:��kr�Ad�2�c�EO�O(v��ȓ_,nDp�)
80&<bfIS�_e^y��tk������,:*��lhn���K�Z�R�O�����qe�֓h�����/�������*X����T@�M��9Q�Ct��R��� s�ȓhX�H�>R�J��@'��g���?D��2I�*�Vm���ҒAF��ȓ}���%O�!��e��N�7�h��$�p��ϕ�T~IZv�Ƶx��x��b� ��� A�^p��$0-�ȓi�^!�q�q\Ndڄ���mZ���&S���$ώ\^4�
��w����?��I�2K�}�tmAe��r�N��ȓm�V�9�Q��>y���^B����s��9���s�:����h'�e��H(.�	���n��u
 '%��b����G���OBI��$��KL��ȓ	Rr}��Ѱ9j�Q�rLD�@Ȁ�ȓT���WN��_8k ]�oB�ȓbP)�Q-��Dx��8H�͇�e���I:v�Y��BUI*`��_K,�a�&�AUx8ڵ��g����)g^ �cL,>�q�&��O�0�ȓO�(l�#����р5 ��Y��W�hA+g�� ��:Ѐ��fj��ȓ*n&��!�L�#x2���ͣ$T ؆ȓ˨�ap�_�[FS�!k�X��z� ��C�v��Q����"�4��ȓ5�:qI�LH�[�(l���֟jNZ��ȓ�T��t�M���w\|����@�F��
I�5�ʏ/�����|�x�Yf��d��4嘄i�̅�![f(
A߻[�D}x��ށs�\���B1<c�@]���#?m����z4fm�Cn͟!N���P7D���V2����hU����2��Q0�~u�ȓD���y ��7t����e7YZH	�ȓG (f�@�*��p��ሳ'���͸��EH ��U�3%�ǒb�#D�h�ac�`|�M�;�&�En!D�����.b0���!��<SB%D��� �L���jeh�;��$�7 0D��y����Uߪb2�,IC�-D�� ��A�\a��왵N��1T&-u"O�PS�44�����A#Hn� :"O�[`��e��@2�A+ q6%ء"O�I�+� �D�b��^ssn�	"O�L�-ƽv���R�A1FV�I�U"O&i*�Iۢ1�>���M�	Z`�J�"O�@����:1��Y%�4 F\(�"Op�#�S EK�����:^�l�v"O��Awj٠I���2�_�Lp �H�<1����R���E�X���PR�
S�<�$̵�x�-O�\��؁��P�<)�CJ:/ͮ�Jv��,����$K�<5��p*�͡�H�$ebJ5�gBA�<�"l9�cf�\Ot��IV�<q�'Q%sҲ�c'L	�t��hSoI[�<1�HH�a�gû�����P�<��a�9'P4������{|���_K�<ђ��"������E�kc��ȀD�<)�"�x1�� L>%(����X�<�*�U�1��
�8R���WE�T�<C�~^t@:�e��&�J���E�|�<�c�"Eєh��^Gd � �w�<!��څ�,�!P�-0Iy[��C�I�)P>ua��O{+2���
K��C�ɋY�v@R1��^����2����C�� �^d�U��|����Gм��C�I�\���Á�-9�<Â�K�bC�I�b�h�1��P+�b	<t.C�S��e`��H$�\�ꆲ��B�I /.�k!�ԄV��5�an�q0�B䉈fS��FgY �� i�  �B�ɊG d(Xg�ٔj���D�:t��B�%mE8�i�C��E)dJ�+FD��ȓH��kޘ=c��ろ I���ȓi�,A9�b�_�i��c�&}2�C��5^��5h��KP�JLk2	�wq^B䉆+8�]���F�H�,qh��I�C�	,$u@qL-�p�� ��7��C��=���`&��g�F��,�K�B�I�.Bpr,D��$h0���a+�C��;���Y�@X9B!� !Dh�\y "OȈ(c�=IR�3aN�(Ry����"O��� d�3fLB�^t*L�"O���S�ݪ�X����
bdp%8�"O��T�e@�88��E�2_h�p"O�����%"|$�ŤKL�#1"O�	(���?�铷ퟑv7z���"O�HzA�\�%�l(Vm��0"OX\��gV�1$��0�v�hq"O���g�m,�(E��*�X�"O��+��H�� �3�Ƅ{���A"O�|toL�ѭ޶=v���"O>$h�b
4"��Q3Ćn��x2!"O��+a������A7N���#"Ot��Ć�m*�ѳw�ծl����"O��įO�R.�Ea��ڤ:5nܢ%"O^���֮uHzhZEH�(N �M:�"O����_$S��3q&�,{'"Ohz$E���bQ�E���ш�"OZ�A��_b�2�W��n9bY��"O�Hh�^$%��aI�CZ��m��"O���ؗY�p�RB��!C5"O�`�`NH�rLpQ��@
�!�"O,�#�� �����T+-5�a��"O� ���B��M�$8��L��Kr�pa"OJؒ,��Epm��e=O�i��"O ��Tcȓ��U�rD�V���G"O�l�mĆ5�$Z2̝C:2�h`"O�t�%b�����h��[11�f"O�� 5�H�&W5P�"�/I!,�"O��z�#F0,�&�!8��"O�� B�F���B�.����"O�(	g��̽���
h��5"O2]�ŨKn�����:S$@:e"OΤ8�-G�GTJȐ��Q�^���"O�\Y�H�dL�ȓ������{�"O��B�Ύ�ΩrD`�=\��b�"Op�j��F�$� ��Z0� `"O�5h�nh9�9Kv��J�I��"Ox�q��G�@��"~Q�*�"O�����ʄ>���2ʒD�d�#"Or�!؀X�Z"L̞T��"O�@�읟WVx�4\Ǥ)�"O$Hei���� uaǼe���C�"O@��l�v �����u���)�"O��I���AN�	�%�)up�E"On�!eF�@�F@RΛc�l��$"O��� ��
�v�I�*�d.!#�"O p뉶M�z�p��\�;42)	�"O8��G_x��!a%�9#.�L��"O<�P�T�y��+� �qy�"On雇�\+��k���ݴ9P�"O�8DiN�M�n��/5��#��/D���(xp�4�	B7��5pn/D�`�F@��F�.���$^�M
�����+D�x���
[7��?E��xҖ<D��S�F�VE�P��J?gf8Zu�9D�(����6Ȁ��!�w���)�`6D�lr�X�^?����BX/��H:q@6D�DK��S%�jӆ�ԯ���y�A2D����i��|2�,"�b,pR�+D����-���Ҵ�H�x 2�q��%D��a��?,82A�ŐG�p��#D��
g	�Z$�.�j�B��d5D�$ⷫ���$�Eo|M��2D�(� /��i9ځ�!���DA���+D��!�B�=c��E��k %XȂdh)D�L�V����m�;z���Ԋ%D��"�-C<$�Hx� ��*�]p�b0D��;a�*~�Y��B��h}���-D�� �O`�J�+�4V"1��+D�HJ�ֶ+�*Y�`�P/?����<D�`����d�+��7y���{�n D��!F+JI���2j�n�a�=D�D��*
�	^���T��&FLLU{��&D����ͫy<T�YG
[�.
(y�é#D���0+�*J4P�� �6~F+#D�hk3I�8,��D��7}�"d�A�,D��h�W� �j�ĈG�J���/5D�`p���s�
���,G��D��8D��Qj�A�N�(� ?&�4��/*D�,Ì���Y◤�n��	�&�;D�\c�((�@r�Ա[�ձ0$D�\kEf��T=z�Y�o�#K�5X��-D�L���7��t���l����7D�<jCa�9|>Ό�����&Ѭc�'߼i ��ɛ^�.���/�M29�
�'�8�:���<gi8��O3����� ��JV�F# � 	!��V:]\Dř"O���"�1#�ĉƪ��.��"O�����3S�<�[2$Y�6�L�k�"O�ݰ&��dYP��Q�E>)�s"O� !v�P�8����>N��,�"O�X�!�;0�Zr��4��yQ"O���U��L��QxS���.��;F"O��a��ܞ!����)��#� K"O씠&��A|�0ڭ�1Av"O�y���T�4��"���>B��"O�u3����6�Te�ĀZ�;��Q�a"O��x@��e��m�S�SmV���"O!���BE����|`�xB"Od�h�)�#m��,�td�w��ہ"O��(l��Dp�RƠ´OZн� "O�u
��$��e�y�^qag"OpYРƃ�F�m�Pi�9K�Ԁ�"Ol� �rd@֧P�&p�!�"Ox�7�H���X���'
Bx
�"O����q�u�A��0 �p�"O����@S�[+v���	#.�3""O�� 3/G�)� �ȷ��9Q��`��"O�� �$fNlQ�@��&��$"O�����at�7�Je�8�Z�"O�EӅb�-}�D[������0$"O ��!�R/眍���>� �"OB��#��O/�����%g��A�"O2�aW�'�D9�F���<8�5"O�`;�gO $ <���F���"O|�q�&`��Bǔ* ?��Z�"O�x���? 0!?^���B"Of|��K�Nݚ�	� ��o�A�U"O"؀�_$�6�P=�j]!�"O���	��t�QC�� �*���i�"Ot<�g�D��# b T��"O(I����C�m�u.����#4"O6,1ᦓ���5jvn�?L��1"OZh0�
"9i��c�a$�ysr"O�k����0d��Wc|�Q3"O0a�`˥=tY:�ՙ9���V"O6@�֫��c��T��e�a���R�"OT��7��]nF��6E��a�"O�`���O"(I��S�C��+#<-�"O�2��	EJ�3�O��9�"O��z��3jN���pA��j��Ui�"O�HV��/+u<Mi�ʉ�NA��Bb"O�<��=4����։~�T���"Oj��Y�I@~A�u�\�uv@"A"O�t�F�S�d��Y�I6!Z
���"O��iR�5`/hl(a���qR�0��"OX�k������ԇͪ9:�,�"O����
��D1ؐ'�q�f;�"O�{wh��V py��'	@�"�3U"OV�;�O$b�`�`�E��p���"OH2�C�V��!PeV&�F(B�"O�EP4�ՖcҠs�5�f�V"O�@�fM�}b 9ei�%d�Tx�"O2�8`�p��T��hY1�zɛ1"O�y
�kHI�����'_4G�|ɴ"O��1���!����λ Z��Q"Ov�@f�>=�Xd�	F���p"O�;`(;����@�z�ꭲr"O��Ј33�AzU��k��rr"O���W�V$�:���!.��%�"O� ��R�۪C���G��8���"O��i���H14A�A�@5D�:��"OFT��*�xϰū���_9ҍq�"O�8I�*��R��(
1M\�F��B�"O>�'Ń  ��ȁ,�8\_�y�"O2�k���*���w�ږ&Y��p"OD�	Ƿ����P$ox���2�_��yBl�F�Nq�EŐ9\���Ũ���y"B��+��i��a�<��O��yri_:(��S�@�*�ܩ��%J��y�\g&�h�(�-Y��Җf���yr��� ����kF�&29��V��y�N�(��X�c"%�X)��N�y�fD94�d`�v@о!���#p'J��y�A"Fd���gR��*7-���y��F7y�V�	�M�9f�H��o�+�y2*�;�n���� 5j��y&�y��*,L*%;oS�$1F�('�Y��y2D��/ô5�Q�ߖ�d�QF� �y��0hЂ���4�4;F����y���3�܁�v�ڗY���ye&͏�y�	�E����7��Vqr��cU��y"S� �b5:C�JFB�A�^�yB�����N�
g �P؅ȓ'`��
}Ӽ��w���K:����ĭ"��
hw�)�Dd�&nMD���?X��(R�N
��ƌ�#lBm�ȓVH�u��GX=O��)rp
9F�ȓ)pK$R�kfa�1��>r���ȓ=���;ANRM%%f�a �M�ȓ~� ����	'\b�y`�ͮ!�p��,<�7�ۓ���� �+f�t�ȓ[��� �`ӟ"	�� v��n�Ne�ȓJ����E��o�"�3�C�\|T��1�  �.�t.� ���4��ȓs@���^�2��t`��>�����q�R�#y��pU`Ш>n(��ȓ~:�i�悠Ku�O %��x�ȓ��jN�r%�J�0)����B�;��{N�qBV斻V��ȓM�|񩶃��0�ґXF�<R��ȓN<J�Gf~F�y �b�a�.L�ȓU��q�`�,��5���=,*P�ȓ5H�I ���[N:L�'�W�]%�y�ȓ�� F����]���K+��݇ȓ@W�&ǝ%L��c��^�����c͞I�1)۩N��D+��ЖD�0t�ȓ�6�I�n� sR��e��M �d����G��[�:�`��.|���[X\|it�4~� Bi
'���ȓ.^�`���LƖ���@I�a����]hL�+���Б[@�X���ȓ$��E	�j���jE�$�X)��A�ȓ����/K�m��`y��?l˔ �ȓ�8���B�`���様���-�ȓZ/�(S��Z�kJFU�#��9�I��K����/ ������;1�!��I�:�qэ�j�� C�6y���#td��P�R�?��R��.8ڎ�ȓ�j���aօT^�uh���p]��o�p@!W D���۱��r�E��9�$�fGS�jĚaG�U!;y`d��o�DH�T��.x�(A�`[�;��a�ȓO����!�I.2� y��oڦA²���S�? *��#�;"��M��Ů#���"O���H%V�X�i`A�A�N�"P"O�����߰~#"���
%R1:�"O���H�5�R� �B	(���)�"O��Y�`V=�(pvř�غ�[F"O���f��52LFE�������"O<G���R�8Б-3g�u"O�L;�cdY��&��[R����W�{�L3U �S`��΀>!�DfQ�H�4 ��7��)5�X��!�Nx(L�;T�N�l�-��Lv�!�lR\���� w�\�(���,�!�$߂A΄)F�WI�0����UZ!�ڂq��2�` �v>ix"�G?7�!��ϺT:���rI')8�{W"�s�!�dUW��lP%�ta�G�}"!�$H�Li��[� �"K0PU
q��"!�dr9����X-�5+����A�!�	{��x(Q�#u���	�		os!�*���b�h� ��E��FB�I�&�(�#4'�:s���[�8�C�	�-�D��ަ&X䀲!�Z�_��C�	�]���f<#�(ZpkD5M��C�	"W�:�J����f݊�2��K�C䉡E-��"��б8��)*��]+u9tC䉴�0��҆]�6�.�mнL��܆ȓOP��o_�rZ
�K�i�=R�Z܆�KzJ����K�e�E�f� =�ȓ8D�4W��\��]K��� Ks<фȓy��A �D@"+����q�ҲjxI�ȓy6���C�*�����nn�=�ȓN��m"�I�H2 ,��^0uxt��ȓIb��0��]�P~��yL�.D���ȓ,C=���
Tĝ��G���Y��R@b\p �t�����/#/�bĄ�" ��ɂ��eu8���ȓT�>xE��!"���m��L$�Q��)8��;���=�|��'�>no���w��mÄ��n�hi{�e��d+@1�ȓ}Z>���ƌ(2��� t��]��H��I�hI��dn�\�"�Ơ@�r܅�Ā�
o�Xv�M�!ۧy}���ȓw�h0�f�]�B��$�E�[�)���V��I�V�5�Lae��3;�q��u3����'=d=��(@�Z�V����	r���ń�d��X�M�0V���p��+��K,����RV�݅ȓ"*�rsf� q8�cI|~P<�ȓB�pP6�&;98!��_�N0��U6�$�ŋ��D+3�����g���[в*�&$
5�'sa~$��H��s��)yI&�
�,θ�y�Z4fvLy�	 q�)�AG�yb�ZfP�zn��b�N�{����y2�ݏ	�
qO�;id�U����y"F�&� 1�o�O$���(��yf�dh!�MM`x�jT�J��y""�;1\�a��D{aQ�y�Of�G�9),���j!�y����NmΚ�3[$A������y���&y=BȺ������Zե��y2
��3�Ƶ��Y+�d�0�m'�yB�P5p��cs�<r���E���yroC�
�
ݨM�r��|(��y
� nuj!hW�q���f	��E"O$�:6II��8x��&%t�E"O֔�p�#��`�N`��a"OLH02�6<X�:�� �\��@�"Of��rA�R\P�y%N��n���j%"O�Ι�`E�Ss����"Ov�,t�
�H�&V��9#�B�1�!�DC�2P� ��L<��г#բ3�!�ě�`���W9K/¬�6C��!���$#����e�\��l�B��rh!�䛸v�6�CR���ht�p`D�)!�͈&Vb,Q7�����#�"O&!�d�Rw�q�v�ǭ]'����J!�$�.#܈���{.���#@��!�䚣'��V��d��!��#�!�d9����R�`�&}S���'�0ܑ�B&4��R�A�n����'9��w��6�>-!�� 1jm �C�'6��R�l�`����V��$d���'(<��G�O���6�I�d���'��dy¨߾&P�r�*SO,��'9T�P�J΄AFI����y�'h�آ`4�*��%�=
0����'|��s���	iB��1N���);�'cZ��m)���� �vLv-��'��xIFG�G,ܨ�eC� w>�i�'B.���CM��\�U&ٝ{Tl��	�'�z�i�ʚ
'�b���Ҿi� 	�'�.�Zpm�4_�fH�����g���Y�'��+e�Q�l�a�/Ɏe�hػ�'A(��5�ғ$�4�9%�܄e*����'�xj$��w���R(��/�*�+�'� ��$������Tlޟ0���b�'% 9�Ɵ娑c$	Q8s�N�J�'t�s"L�T�$�&�-W�,�"�'��"�RM����&�0\
�4��'�����Չs��)���F2Q;t��'�r�"���G�v�	P,�6Oz�5R�'������5j�(p�i1w���'YIiVfCy"��:�|��j�'��ݡOL�㔵H�� :$�U��'����A҉
�,�{#Z�<v%b�'���@ c�-�dE��)f{���'l����&��6�.��D��3_�œ�'��cZ(l���)��F�����'E�m��H�i��a􈘥M�����'o��Z�NME�D0hV�Ԃ\����'Op,�D#��t4*غ`e�Cۘ�P�'nx� T�@�0�`5"��@�V�ʓe�Li���YUĘs ���t�ȓ^�q�0�D�#�^��$I�@��Q��x���#��օK֌�%ߨ7D�X�ȓG`��XT�I�9�F�v�,���&�d#�(�J�V����J8dɅȓ-W^�h�g�-���đ310�h�ȓD�L�6$�<P���J¤_�`��ȓjN\��R�%�ےGіud���E�ͩd�.o���#��J���N�<"��E�7�@̛�+�k����w�8k��	�Ӳ�����͞h���Ɛ�D�F(jlX�(�̍3�Ґ�ȓD�+�͊�M�� �!W�C���ȓ#/ ��Ю�Rڌ�0�����,�ȓW�����Y�,�4@ Q�\�Pfd��S�? 8L��� d��+���	a���e"Oi�	[(_�ԅ@���nw���"Oz�+�7wخ��%G�"s�(��"O�y`���n���p��;�1U"OZT���uji��h���r"O�d��XQ5f(C�L@�r�%��"O@M�7ɖ�^�a
���&��,D�4��a��.y��0��L 	@����)D�ز�$@1Vm� 30��L�j���N&D��{�K�-X��H�m�,�RЃ��"D�({D��=���#��/fY���%D��cr��U����HU�8��ݛ�
"D��ᦛ
EEry葌��c�U�� D���pm�1gC��6��[1��%=D����'S�1@	R��%-�e;�:D�d�ER9r`Z�Y�B�
eԾy�q+9D����k]�UXx�/W`G��r�K*D�x�l�1d 2���\��|
��3D����G'���"��$G�Z8X��%D�<#w�N�tG�-�C�<%Y���0D���#u���F�t�,���/D���Q`�)q���sf��T�`)�� D��ଢ଼�@�g�^:�`]��c>D�LSe�Jz���1�Z�-x6�1�6D�(��(/�B��'DX>�a��/5D��s�n�*7�p���W�>�@9�+&D�����W%�V@˶���*�s�#D�����T�¨���=:�1��!D��rS
)H�8�@R!�/��1U�#D�T;!'�4�2�� -6H1�'/D������:e���7���a�F��@(8D�Jî�}�ĩ�$�d��ӧ�7D���f�2j�@�x��'d,�hj��7D�H��F��xN�,B�mׅL�{��9D�h0)R6�҃ET33�]b�k8D��ۗd���4\�o��m<,h��6D���`V�d�4"�B'Q.�ba�/D�@B4�H�e�� D,C��e
Ӧ3D��q4/݆Z.�)�k��eJ���0D�ءס��]'LdX���>���*D�X� G�)~ ����0����3B%D��9���a����/����4�?D�D�Ą��+��P��R)/���u�*D�0x���� @Q�C��~�.�p�*O���eo^/^�.��c*ݹ�3�"O������*v_x\����=+��m�S"OJę��^�
fHx��$,R��p�"O޵��ϫA4@�% �=��k�"O�ձ"���X��H	.����"Oh����
�8��ǃX.S�,"O$�KF�o��Q ǁU P��q��"O�0c�Fݜ"�,Ո�E�f�%�5"O.5R6�1,̾���Y1�h���"OX����-��'��E�&��D"O��ˑkR�����1��fQ�-�"O���6�	<V����g�� "OEȁ�M7�l`C���U|�9�"O�!��#�v�Z|!��հA�8x��"O���6눟l�^�ҡ,�6浂�"O���bC�	2А�1N]�Z��)t"O�A�"@@*��Vc�3}�$�P�"O��h�gɆZ�$��UB,�NT��"OF9g�0G*�iq�?xﶬ�!"O����͉-e]\��e ݪ$Mڤ�c"O� nm�'���e9� ����I4hd��"Ot ��ED�C���*$�I�q��["O<m(�
AQ�Q��ꈕު0�V"O\8;���
R�v\�j�%|ˢb�"OD#�OQε��O�!���"O� )Q�ƯM��)���,N�J=J�"O��d[�?�<PH��=�e"O0`�}���ڲ��g��\r"O8�&�\��\��P�ƿ,�Lc#"O��ZBc� 6V��w�A	9̄���"OL��B�,`u{��F�r��Z�"O��G��?k��2D���djq�"O|M5�гt������~��;�"O�H�a#�P0ȫ&����e�"O�J ԝ0`��k��5/s$@is"Oty&��)w���t-�+F�\c1"O��R&ӏOA����I"%F��:�"O&��1��WN�����7<t�[$"Oލ �g�oZ��"�X�5+���"Od5w�N�5؍��n��Ukv��"O�ı�ϋ�"�0��D�OD�)�"O�L:��Rzʬ���_�w�Y��"O����C�8�ؖ��r�(��_!�yB�ܛQC�eB�L�l�4�@��y�#@2��ar�#~����^�y"���b��╙x�HD��ƛ��y��W�^�����j`��;�B��yb!�%+6�i�kYc�:�+a]��y��W�p�4X{�+'T,��(�Ō�yb��5R�&���[.~��[Վ�	�ybH��	�^5)���G�$E!�&P��y���O���K�Z?C�m�F�G��y��<a��(�R�e���1�\��y�FѵjcvY��IDb�h������y�ǉ{����q��1��ls�k=�yb��^j�(0j�9��\�+զ�y��ڀ,I�l!��E���$�0�y��!Ă����t���ġ�(�y*�T�Fa�c�@L!��ו�y�g҄{8�"���$0<�B����yAOE(�5�ס ��C`BK��y�'D.q�D�����>JĶ@8�'% �c
/|��Q�`ѕavt��'I���.�`{��ЇM�~����'��p�͌���)��-O�a+�' ��x�E���sVB��"���'���+h��\�21c��:e�2ɂ�'ߎ!��	�6�&|��"I8�-;�'���TDƥPC*hcD�>E��+�'M�H+6�ZZm�� $',Ph�	
�'w�@�2Ƹ��̹s.P�=WD��
�'&�1�դL
�]�[(T���yR�NI���шJ7���3č[��y��*#���Y-�)Z���KP���yrIK�-�T�D�ðMD2I뗏�9�yRF�����a��@K���W����y�&�]x��z MM�k�J���jE3�y2��:U�
�h�̔�\S�5���X��y��[rxH�-O1P~ j˓0�y���d��`M)>�6	x$W�y�g���E��>MC��k���y�ϝt�ʠ�W�S�/e�t*�H���y�L(9�� � �:���CǓ+�yR�P8:�e˄iR�.X �� ���y
� R(�tjJFQh��.�+tݨQiq�|�)�S���Y���"��Q8��Z�?~0C�ɒZ�����j��Iw��B��W��%ȑ"a�ZxRi�jC���0K4-R*rDPg��W\dC䉫�ҡHU�X+��� ��w�RC�k���G*F0�� �\#X�dB��'n��E#�MA�;��"�\:Z��C�ɻ�L �Gh�D��ʛ/ѪC�ɇ"gp [&/R"_�^����/LF�B�ɟNs�M�ŀ��k.jh�W)�s��B�y��U�SnR(V>H����T�zB�O(H��I'Z�܈J�I5ŜB䉊?x�պ`�$4k�P�w�	��C�IR���:�Ñ�8PE�/N�C��uB;#{d�� 1M�C�	$�(�� S�b�ON%zu�c�l��{;�=���	�*��-�J	z��>�.lְ���49��US�"-����� ��p��Y����cF!ŴX��	�<!�΁�Z����
�BP̱��c�<uJ3)�a��I�O��PY1b�<����M$T���Σ<P��v�<Ał�;|�@�AC�D�$З�2TBў"~��l���L�2D�����$�����5?ٰ&σt����L�>���d�����	
�h*,b������"%O0<,G|B�|r��ԉ��O����/�N�H�SB��yB悥z�����m �7V���r/�y���-#4X�(^	3ﶤ�G���On"~:�����,���zΜ��@�O�<���v����+�h������a�<!�i���~�a���6j/�Z��g�<i1� 7־ȩ��J�TB��Uo�n�<�V��'y��pA�06��P%�Uk�<i 1,t
ƫ�/:�lE�A��[�<)�ʋ�6^�Q���.a]���#�PX�<�!+t��1��U*Ie�l�G�N�<�mޥ	q�K�T�
R���&+GI�<�#�4�~kt��k�Z�0QƉE�<q���`�*���� 4\�h�&�w�'{�T�'�t��禇%1$�U�VP�#
�}��'�&�16EU4j����������'��I��^�BM$$b1�����8�'Z�� 	F�eH>�А%���Q��'��y��`��B8c�� eB����M������ ��Є@�Z�@�O�R�8�hc+D������ #wx����R�jdq��=D���򤊁H+^mʄ�Z>�U��'D��ǥ
���P�X�m�Ԑ+Ǡ%���<�#GR�20����/rZ^p ��{h<�Q酓�����(]$W[��C��;�y@�<Eٞ�:���O�$�R���p<�!�;�b���Fز3W�-�7(��r��L��cځ�도=w,�	���50�P��	C��<��"i��A�-�=/����i�@ؓ)� t��MϏo �d��+�ڼ@�c�y,t1u+O�?����u ����ƀ^J�P�+�4��>I����./�1H�!ōq����:�4!ᇄ�M��  A& N�6��IJ<�)'}�
!y�c�?P�� `'*�K�<I� ��y�B�Qq���Q�6=�+I�� ��ZTFБ)��0���f����S�? ��x��[�w�U8��	�"b`�"O�@��n+h�A(�`Z��a"O���_.^C`�S%��m�u�2"Oj���ѵ4F��E̴J��8Qw"OB\��i)3�������N��Q��"O���A@�YF��1���]�i2�"O���D�;5�e���Y$!t�4
�"O(��'�>�ٷ(Q�eB!�Q"O��C��*jz��e(�1<ā�"ObГϋ��q��
�"|h;g"O:hp��C�`�N��&\2x��C�"O����HokVM�sl�<(%�a"O�X�-W�&>�U:P��N�(�"O4�)�. a��as"�1@��,��"Oz�0iY���D�0�Y�}N��4"OL���Ȍ�!@r�c&�����8�"O��`���B��+���L��4"O$�[D.�<�	�NC-u����B"O����Ї,�����Ā1˂5R��>A���	����(:3-B�#���y�*Ч�!�� o��\+&'�l�V�k𨄍�1OT�=�|��O�2���	�E3$��Zs�p�<�1n��0�ԉ��ĵ˚�
�q�<Q�a��n�Tj�J��*��0�DM�m�<Y�@�E�4��H�2J��Qs��i�<�B�a8���+�����Ar��N��hO�O���q�hG�*��I+2F4:Z�z�'���j�HF>��a{4��y3��H<��W��[aɅ0L�f�$뇮iƲi��J���ԭ��P�iR���(/����=	ۓ1��U�%�tҾ�*����d.�Fx�)�CV<r��&�&�P���-�s�<��mR�5�L�:ׄ�",M���&�Xq�<��DE�h���TOSx�ը��An�<��EZ\wfyqٿp���M]k��!�O�M�V�Z�<)���� �Q�ey�"OD;pL�Hb Rt
��q"O�0V�"	:pFˎ�`�ĂC"OXؚ�Bäu��H	#a9�T
�"O�H�^�B�Rg�Z���"O��s��0O����4��]R�u0B"O��򰈛� %t���M��'C>��"O�U�~�V�ȅCޛ>��I"OF�R��J�@��; ��}���"O��7��-A��ۚ��Ų�"O�L�VE��/U�	#��.v�@!h�"O}�u�
D�b�/��R���"O��b�FK�:��[)���LT:�"O�P2��]��#��C�E݊���"O��c�k�"o�ʐ�toM=x�x�C"O�,2�,*b��S�Y�9C̔C@	 4�\ơY>&��P�d��>4GV�B@+1D��
�H�w̴(R%CPw� p+F .D�|ۡ�-Hw"��bO;B��Qr�,D�����߇#QbܰPOH:"Ј)8�b'D�$��V�VT��ၲbkpQ�.0D�paD���L�pz�g����)D���		}�� E%ޕWM\U�f)D���Ζ6b{��:��)<�`���(D�<��������A˝�5�x��׀%D���C&\~<1G��D�	&d$D����>f����ؐL
D��6D�H�AC^���� E��eD.�3�?D�T(��=q���׬ �y%0�#�h?D�� �9�ĢC�k��F�,L܄,82"Oq0@d�"�"�/��	�ĠZ�"O�aD��%�w .o��Ӳ"O��2̥f���!���(�R<""O��CRB?,?M�W�%_��x�"Op�s��V�`��xQv� "R��xa�"O2h�$"� �ڸ�u��w� �`�"O�A�d�4�|�*�ёX��x��'8���g.�
s(	96��=i��@	�'���{!NS4���Q�s��4��'q�<��4<��X�%(	�U����'���x�{��4�t�.I!�(�	�'��a���Z9�H�c�A.�a�	�'?F�P�BC�ES�m� �I���	�'{r�EjS�MC���R-�9Ty�Q@�'�"Hpi="��KQ�Ud����'H����@S#N
d!S#��/)l��'���Pq�Є\�t##�V�0��
�'��B5���x͚�ȥ"51���'z���ѮL�c������)+9f�)�'���w�ټs��4B�.]!�,1�
�'EVгD� Yv�bmХB68�	�'� Mz&C؉A(Fx��A1�@S�'� t�p�S�H5�4x�g���Y�'/����o �8�
u
�
���1�'jn�K8F%�AJ��B�#�'�NI#��F-f2$R�o�wE�4��'FT	�D�H����c�i�Nh���T��PX��>����!Q5 ����j�,�ȓ�А��K�T[n����L ���ȓsV�e����[��C1k�
`J��_��! �3\J�YcqΛ:0f�t�ȓ9[��S�-�2��`��H7*M��ȓK�Lu:l?v!�{�hҳ^��ȓI��Ӂ��;���
���Ҳ���ؤ�*<l7��8��$�ZH��mI� ��^�Y�*�0`�ї��9��8��%(އ9ir�8 ��*e`��ܔ�r�"��+  HS��<`B�ɚI0�aGME�N���*Y�B䉁'g���Th��4+���!֣�
B�IC#����bI�[&&m��bJ�|��C��X�ұ��W�n���kUlduC䉊|/Ʃ0��ب��ě�J��:�"O4`�+0 ��x�cQ�ݺ�à"O��Uf֑[�td����3��Hd"O�-��J�B���"& O �0a��"O�|��ԺRe�LC�n^nn�H"O��D��|Ɯ���M�ni��"�"O��Yg3�1kvN�BШ��"O��YO�
��ԀP�
�%<�[�"O���P��6xC�ks6H��"O���Q��l3F�9��؟O�W"O6ݡ�-�(�42S�X�>�ڣ"O���
ϦH��&�\s�"O)��_�F��#�dF?��*�"OH��B+]K��zVA?u��Da"O�Ô�}��%��͍-U�9�%"Oޜ��N���}����CO6��`"O�"�k	�%����t��$Y�5"O�8
��L0$���3қaǢ ��"O��ҁ�D.кa��Y(:��W"O��[4��	�NE0dY�N	�t�T"OIS�A��t$|h�����-�"O� ����ٖN�t14/��I�,J�"O ���M��Xf�"�τ���x"OP죗���KvF�����qv@��4"O��Y�%�&"�lx�c�S��ĳ�"O>y+��λ�,D�F�O��� B"O���`�δq7��[���$�	�Q�b@ 퓁/��(��ƚ�R,*��aDô�BB�	�Nd~�h bӷ ���%k��0F��d��#0u�>E��'����������{��|��'���	wN��Ni�!�&�Q+x�h���42���葩M7&�"0zO9<O�1���M#0�����%��c�'a`�b�9-��L�xd�1A-2�P:���$�"��WO�����#�p�@j�7}(���΄�4jC&�6v)��3��K.�Ł�	Y�h�X�JB��'G�qr3�IV!�<�6L
�a@NiB�@%3;�QEB�i¤t	6d4�g~H�1l֮�zNۑ1v�33*N'�y���������R�\,����A�z�S�m�9 <m�� E���Q���*h����#�y�' {��C�&�e�A"~�.ʑJ���T�P�I�a@�����m0��R�l�/��娳��>y��mk<��֨<|�����+�0ز�K�8�jc>�2�B��|y�f�׫Ԃ����;D�Xh��̖V�,$��T�6z���䗇S��X�M��,�D�P��HNr�?�z�	�<y�#(Fr�p�c�FU*�rF�Wjh<	E�<Y�v�H�(��)3���ꭺ�ôm�d����7	<�B�Ξ�}���!ғ���S Ǿ���xC�I��@��>���8��O��p�k��3��Ӂ�[� ��]����/��pO��LҪ>�Oܼ�ORwR��Ɲ�BBDa��|⦝DR`1E̸X��a��n1��Qz!��{�h��'�E�NV��I"O�}S����x��IAB�>M!��R�Cܵ�<5ҷ"����W8�2�	$?��ШM�Y��ˆF[H1��]J�<��ԦE�� J��ҁn��j�&V	�B��^M����A5A}�A3�>���b�&�(R#D�MD��%L�Nazb��$'��R&P#r�t�t��q�[��1	�R�08�A�WT�$���p=��m�%�xѢ��%�6D�b�qܓz*}����o|b� ����'Y���@wE�&�<)�G�A��T�8��J�<1�͕$3+��c��I7Go���&R�r�V]��4]�psĦY.ok&I̧2)�c���7Fm�'�8��Ҋ�9ХH��S�l���@M}���a�&/L�����%y���A�ֵ4Ut���\-�L�o�9`QSse�z�bc�8�˿[F�: a�17Jz�.�;�xQ�/քR�X�P����L�-��p
Vf�%+'P��!�ߗW����o��ag�Y�{�����ɚK8���$��7((f�Сʓ�<6M�q�
�v�=Ze��C�6�xL�@ mTX��#�|z3iG567��-iY*hJԃE�/��ych5D�82Dj��=�~`0�@]��LC�lޡG�F�#���M���7"��1��?�rX���Y��hL��t�?i������rT�F/�Oh�!M��9�:��AG�I^1Tɕ�Az�9�EC�yl��d��D�Z�0�A� Y:���!�)LH7�S��1O�1@e"L ���!p�@6y#Ĥ{��ɺ�����	���I�E5(ր3A�[�P/F�%L��.��5F��$X�9�NU�U��Ғ���_c��Q��'����&醞g�ճ����T�Fh�.l�|ā����,��D(�T-l��Ѫ��Gl���ꎅ�R��/n�Rt��  97��{�d�J�m��'BtW&V� ����H��Y�2hT�Z�ЅB Db�h����_�-�V�5�\%
^�H&,GO��e�u���$)mm�`���;b�a��,]�p>Q�)2p*��􉌊:��P��I��\.�RT���sٖ���O[�:dEéB:TDBg��	<��l��C'S0b��D����ū�3�`����3>Q��#��$_oz�����26�\��FT=41�]ڵfD2`384+6����U����&C X{�#�1ft�!�<IR�d@��T	��3�ǂ�nG�i@FaԞK����lQ�wp:��ޅb^����)�-['�C�mC�i`fA�ePby�7B
 �x��&P�	����ȓY�@I�JE:qj�Ha�Ju��@��oE2�N�����	�Kp��p�OD5�T܁sGV	a�xh�(��Ӂ�̻k��������L~蛧��\x����
�ƤC����yo��Ŏ��zƦ��`��a��p�f�X�%��̋����q��φ|d�1�5n9�	�
�dȁѡ��wF���$��9p">Qf!�;42��.�?Z�ޠ��b��@'�3D�u�ţT{L`j�T�a{�;���_dZ<Z��$\O�a�5,�.$�<�A��2E�A�Ov%��!��	6��@$�S��.�rV$V\U����C�$ݠ .c��� tQ����̚�ɹC�$D�l�FȞ/���C�k�y'����O&a�Ё/�<a������I��`Zwz�O�Q·7�� ��ʇ�Ȅn��a6� k�)�UO������Hrj�9��B <M�t�p�Y�;����g�%u< ���6�������;N}t"<9���d��%7
�rK��O�hx�,+W�[&wF�%�u�]*7΄ (�&�n#�U� ��!rJ� �׾Pj����ڵ
�����E �q!����P)�"�W@�'��HuBXPO��2�!�$t������S,�E�O$NA���J�]�Ye�IG���'C&T3Ɯ��dɂ��)k{J A�ă66lҝ`a�-z�
���G���O���x<O|+� 'y��b�(r�8��OF9�
��c�T��ee��9��I��I��,��P��_[�ܣ#�dx�X(b�׿!<��љ"�"�S�K6<O8ږ.$�<�+`+�!tQ���h�,хqA�`K�uh<aA�S�͈-�#DJ�6P
��GH�	�3�Nq��!L�DA��Gu񟖑�6&ɯZ �:&�&����"O����(�1!�.����l�Ղ��ݲ2��a�$ا:�ڔIv*ڬ[���>�O��PT���_��2"�Q8%@�OĠp4B��nʺ�sA� ���{�D��l�*H��=��P�I_�tMR���	//���C ��h�f��У?a��6-�vZ8W������H�[����D� 􈐢ѩh(<Q�Bӗ���xuoN;G�QCey"��<:�y���̶�J��D�1{4Tѓ�����z�vM��ˊ?w<���e��yr�UF���&I�Q��I��-�4@h@Y4No�B�0�ܥlҚycd��G���iU�P��UΓ�yw�6=F���V�<�$�U�ǧ��?93׷9�6�SQ���w�~������T�����Ȓ=�~�#����N!Hpc%,�ޟ�+�nG>p�`��T��7����8	vn�"P��1oe~q��HџЙ�j �Kʢ���$ħ5pA�nC�&6��A$��5~=`c/�;+p\H�!cӌ�1%`F�j�Je
Kџ����!H��a���#�q�E�<Ʃ`�Z$`6�ע�\L�h��b�.�A�h��b�h:�����If�߫j�����)X��1; �	�fU����5j��2�]�V�T��C�\']Rl���.��	"�	E)>��Q���E�n�4Т�\ U�T��Ӌ�Z�nDc�t̂F��%z�����0q����d!�h�=�8a:�I�tq���U�9�ؑ.�!��{w�ݿZ�ތ���:�&]B�/3r|���%O��~"�єt@�h�5oE/{���Q�
�:��O�)�->�򕂂��.��x+��ݕ(��2�K�ir��OF3�6�B�x-b`��;�h�	pH��(U��>�CE�.������g$*�nEXy��9&�!��H�9n"�(!J29�<7E2�+�O�Ѩ4lEy�V����/��	���N�Z4���
~��tm�Ut�t��'G���G�H��i	�'ͧm,�X��	��lu>���j������/`$]Z%
�tp go(�O�����M��d�@ǂV�d��昛_������v(�7���ciy&���c1Tt���V?���
3r��h레�=_ͤ)���R�'��i�"�B�o�j�v̓�}D�]��6"��|Y�.Y�z�9����x=]kbȉ�Q��Y�G���д��OJ�tA�	y�D�q�-]#v���\�x
�	�pH�D�a�0�,a��b�g�H3�$��o%Z�rTo�*AZ]څ@S���edEϫD����	�BP0�{׃Һ
v��viRv_��b��8p26����Y n�0 wE�.E_.7�'p�0dMR%�tͻ{���2�<"MZ�B�#�~�����t��$a��B��ۃ!�$^T&��А"��ji�2\��K��W��(b��6�NAf�'O��PX�h��<� 
�����
уDU��.,Oq!��U#�����B�X��-�=R��8�eM�n�(��lז�[�Ϡ[[ȈIp��Vvf8�FM9�.�8&F�A`(�Z�ӝ+���&��R�bӜ(����B�ȑdj��(��C-R&.���	��+�qu��$0��e��O+UR
퉂䕂R��Q*c�9�O6�UF]9�~����%/V���ØSbډk�/|��}����W(�i����f���*�$��1�>D�1m�j�,�7�ϯbg��2�"OҵjF��@(<]!��D�OCD�(c�(`��Q⒗5^��$d�6*�d�ڙB.0E�C�MEJ�p�'a���F� �>|�0W@�� @�p��*%��2��D�!)6V�B�<n�ֈ3@b�<����T�)F����L�/��i �z0�)TJ	6��e�$ۣr�t�Gy�l��{4�9D*	5�A��D� t�n�÷�B
dLѸ��˝p�0� ̝^^����ՌX����d.�m Dl�2k��$��-7Q�'�AyV��%j�Ɓ{�Ĺ��}�m��fp�#̴���H�;^A*Z$B���%��mו�n��ө�蔵b�(��d�dy�`�(=������j��4�=��b��� �#}ڡQ�T}��>����5KT�I���2H�<Y%���s�[�J���d�,������9?�΢>)��I�#�*L6���h�`x�G�Yz��H(�GZ����R�N�'$:YB�-���ٙACպ}S6XQ��Q$�$����>f� yBd)&�P�8� �"�n"<A�cՌ�r�fDH'QI�`I~�&iMvT�m�q�w'��`�Ĉq�<� BE8�h�26�H���޾.N	�@)�R%s#�t�K?E��),�s"��%F�ERC��k�h��a��P�/�]��*�+@*��%�X��j+A+���dS�*p�8BG��!������x!��(|�0E!�IO�A-!A�(!��7/���+��D3|j�Jc��K�!�΍<����я�!k�8��Mu.!�$@�P�L�#iş(Y�	����T!򤞉<�����K��o��l�pj�!Jr!��"%�֔#�`J
q��|�� ~j!��4;4i(���|B`B�;h=!�DHP�,���
��<Z@ E�O�!��1,�i���M(}A o3(!�ބk�+����6��'�L�!�"d4�J�B��,�X 8g!�!�ė�.`��jG #9:d�ׅK�i�!�D��+�L�)���$~(0��Ǆ���!���Y��*1�Z643hm���y~!��'But����ݸ5�1����n!�$ɪ�Fa)����R-:A���w,!�$!Ua�A;>d����%F�!��M�j����0e��`)���䨒�U�!�O�Ii(1�oN�d`M���f���'Cfp�(_1eG�u1�#D�jfL���'~j�`⩒�!z�ʣ�K/p��t�'+:q�&nԷwA��x0F�"߄E��'"
T `�Q�VN@�bM��LYh���'��U��/ �A��
M$Ҡ��'XBYr�^Ly�FMU"��'V�90,^	��Y�"��;�TK�'7HȪtb��E�����2T����'j�s�B�*l`��#ئ2��'v�e
c�����	����Ǣ��y��<L�I��@��}"�x�K���yBA/Z�b�:�V
I2Fi��y҈
6v�
���� �cʻ�yB�Q,k�.9Be�M�|	R��@@�yb�ȡGe�=�t��rl�����2�y�,�3�`��ʜ�|��}G�]��y"�_-���J�j�Ԅx��L��y��Y�VG@�[V�,g9��Q	��y�"�
`l�\ó�+�B!��6�y��X�%r��AU)�	@ب�R��yREВA�N�c�(�X�F�$�y��^�r�n!��/S��f�Y��y⧙�.U�pX�cѮ}������y2��YѪm(u�Y�k��0���y���.j�5ۃ��k��<Y�&΃�y�F,.͊m
�N�6y�	�g��+�y��L-+��ەl�y)��a+��y""Q�S4��&���t���U�Y��yƂ�L� ����2S�x\5����y2�7<>�i#3�,T�p�!�-��y� 
l��8��Y�xR)�����y� џP��L�J��<R��G�D�yB�@�W�̽� 咕C8lz�X1�y2n\:4Q
��Q�)�E����y���H��-���Њ�N�JJ�yB�@�V����Ā�=��T2�7�yr��$�Q�+
�5v���KS��y�BF���łB���"^<D�F����y��I��������kj�i��%��y�^A}�a*��D�Z�Px���y����*m!�(B]�jaʗ�Ȕ�y
� �92R=j����ɀ#U�<`!t"O��!Q^3RŠusd��>C(��"OL�J��P�{��ݨ!��*4���"ONP��Q`D@��D<d$P���"O�2Cc�<8�OS����"Oh��e�A =�T���3pz�hr�"O��񪇲S�^� �eT4"O^����2��z�,^r�'"O����
�N���D(ȇ`>�QA"O,��O��"F��
+�(#"OP5��؄��1W��^/�z!"OaKU,]4VQ܁
c�R�/���g"Oj9��_ 
zA��A�M0j�"O(�W�E&l�t�����Q+е��"O~e�4��2/@p����X"O�x@F�ۻ6�%yc���[.�x90"O8����$w� I�O'���s�"O�ţ�@f���bS��L�}{"O�diք��<W��,%�*���"O2�J�U�W���ZL;��i+�"O̼�I�l�D��'�۽#�>q�s"O�\��RG��Q��+43��3"O�5:���5���+Q�})�Y�"O��p�(��i`�l	�g��e"O�#�)��p@$����~����"O�චߛM#Q��He :$R�"O��2��4N  ��GFir�:g"Ov,�R�W&2�|�C�H�<BniSD"O�=2�K�8�J��r�Y9"&D��"OQ�E��p�)8�=�"O����N���p�j�W7,�$5�"O(��BU�ʍ���R6 鄥a2"O��0M��`���o""��4"O�`���8 �zya��K 0y�"OD��gN!�VZ�9���� WF�<�P��u�M�� �-3�i�aM��<�͔� ��]Z��'{�NIS���]�<Q�$5u�܉ⓡ@ E��5͒P�<aP�@�e�|9C�ݜ9c�-)��R�<a���$Y+�$��F.9�q��w�I��'ob�C�1�(E���O�%	R!Q�jːI�t�"��'8Hp7��){qb4���Z@b8��ӪH�22z�SV���9�dP��>Q�,8o�@9�߼i�:��AT�'S�!�`�/S��W�Z�G��j0�����T��A]0���L>����A�N�8���5pH�"�6e{r$Iކ�m7'u3�'oH�8�� >��iKb`��1@8}궄������ƱFi8{&= "���`2V"OQc�-J
���-	����GQ�X0XE�2�ĠG���ja��u�Ӆ,FJ�د ���a7�*ِ@.�����I��S��)�R�'T��&h�O=2�ۦM�h��SN=�#�cN�k��zFټ?B���P/I�Q;�h�-�!c�������ad�Ӌ_C�0[֢=ʓd)ֱ�.��g~0�+�O�F��~�\��l£t뾔�p�	�i��&c��Z�4
�.K���|�̂8t̬�5 �)�"Pbe.��*�(��1��Z\��a�æQ�=�B�C�ڀ��@��6pZ5Nـ�y��7SD(0�fC�im���N'�yR`D�#/$M⃗�y74P��JK
[
XPP"���$4pA�W��i����5��ƺ�t�H�Z]�ᨰ��*&r睝R,*��B3:�ղq �>IN����ƀg�6���F��]��Ct�(����U�Z�D� k�$n0�u8�l�,X�@����7��i�f��G�'lby#�4���t�OcF�*��DD) kr9!��������a HlX�R2��0�>��ԈO7aqd	J��N z�H�>��ÐV8���`e�Ku�U��!�orH�+�?U����G�]�4���QRz��!0��0��˂���<��EVҼ���N�Jn9�S,�!\r��v��H�<�w��؊��Ü�zz�49c�˱~�nгPY�e2���'GJ�6��,�7�矎�#�#\.y}�(��
�l����7�J�q��ix��i��(����9`bW�y���!�*A� �9�
  Yb��	�/j�zD�����0�e6�:�J0�F�T�P@��I��0��XF|b�	$� �J��؋,�$}[��֚Lyй8
� ذ0@��J
x�2exp��f��9 � @'�p>9��P'�4XhC�3����F?�������� N�*�0���]>���țZ���ܟ4�!�/	77�lp0 ��l����"OV���tN}��P!0Y�Ha��M�VL#w�U5n:	:�%͔�P�}��ʉ�y�	�y�($S���;7�u���U<��xO��LP �ӡR8�qӍ.��$���M$)J����4���A�3Z�=)� FO�Qh"��!<��x��qx�XHBH^&$1�� A�3�� �X XAz���!84� g�.P���%�}���BS�د_K^��c�Q (HN��э4��Q!+O\ԡ!m��3�����dU);T���~�W�pq�k4	_K[tx��d�<�TdR�]~d]���ǐq�4���OH8ɡ�K�p	�4~����L���a �"4fz\�ueC/H%���� 4��JW#�G��X��s}2mk�(m���'!]a2�z�h�;=�����	B>Ѡ7�C�5�:�	�B��l�T��C�6�(�a ��H��1(�&!#q*Wc<;3�<���4�Hd 
�'��頓�Y8_�u�GB&a�Z@K<���O�΁��fY9� ;�k=�S;G�)!P��9+p騃LŹǶB�	���ѓq�؀.�&�b�"�'lv쀱
Y�L�-Ђ	/',je�vA&�3�̯	��H��N�:%+��'4!�D���Y5lS�T�B�����g�bp�КP� 1Ո��X��$H�J�WX��	��/�N(؁�I97$m*�i7��X�8!@Ƹ!�"��d	U$Xc�}���4L23�7�h5S�Rĺi�F�X\��՜Zɾ F۝Ky$P�'rl1Â`՚hz0��IP��)E�2��O�īcb�c��5�eA�(���',\���+@!����D� �`5� �Z�~�j��<Z�J �щQ
P-T��OV+A#�蛕,��<	�w��Qc�(E�=!En\�FF1 �S��M+3c6U��Q�ƯF�
Â�@8LT3����|�2� �/7$��ɵR�8��L,A�2�O����H��4L{$'Ω^��	���I&!�\��P?�d��h4g��p�QD��ȱ��Q�L��2eҹ�D6_;���C��tR�\"W�	6I�,SD��(k�Y�!��]��*��Z��F�A�hu`3g��=���RJZ�R�Ú�S�*�ٳ��e�X�a�V�hR4YU�x�r@i�LU�7�aң�� ��2�ɚ1Gz&���I�.2��3�"˭4��=[�'x	���R��8 )��z�[0Ez,��� �(�y'&3���3+���Ԁ� ����?�b�Ӳ��8(��<-�{��e-T�-i��5��쌥z���2-���&��[��] q��(r�4[�"��zs-��S��m���2�D��&��	�BQ
�}9��j��R���x� �P�c#v�����q�tHu���Ms�D�=�.��܍��4���� �OrT�ԏ��g��H��?}�>]��Q�\P��A�%��у�I�2���Ę�M�v_?y�4�>^b�sp-��NER�&۹*��h�S8�v��d\A�r�ӓʛ����"ҝH��yi��F�:��5��)&͹�W�� ː��y�@]�L}LQ�!NWDo�=������?9ŀ�Hi�h�4�X�}��i�c��o�z壕�7JՌ���OŊ�K�k��-�g��*p6T����Z8O�0���F88`�І�{ĸQ�A����n���H��s�%���Ʀ=G�pp�ہx0FP*p�؋]S��c���*�-���E&�����e٬?��U*��:�8�0y ��մ4���S+Py�q�'
D㢄�K�R����KZ�1! �(@&ȋ$ꕝi��Vi¥d�>�A���-@�D6����l���~��Ɓ �:�B��"���߹:)~0`pLB���!���^���"�M�5  =@7 �# ��>pr�ѵD���C�En��+���v�� JĠ��)q�q�� ���4�D��2��ٴ��CpA��cQ�4�!�ǱW.�X����LE1�'������
X�6�����x�b��
��D} ��7v�Z� ��Ӿf�b���L}�]�'�V�J��d�N��L���{�|��D/K2�l4���\Q����f�-�a�3��'�%�!�ۏ7��1	�E�	
��H8F-!���P�k��ZNa���֚KMp��-�\�F�I���=�f����:�<4��d�	i�")�w�ϯ	m���(��?O������}���� �/=�& �SĘ
o�05�7�����;O�6Ԙ1�Z��r��I�SRta��J�z�ZMG
f��%i�!���~�˄֩S�`�(V�c�=� ��?�BU��e��=Yơ"�h�	��n��[;�� ��F h2�Z!g8�OX���;������:?���K7�$$D<�b�{�����=q��p:�$��!��=�7�8��O"�9��O���Е#		6�|P@則�&�)'�R'N���H�3 �H8���tonQ�	[(�����دD�εS�IWR쌠��rt�����TW�
.}"�2��Ю0?@��D�&
�Yy�b�2$���!��%�FV�)c��
x��䆗:�y%N'��W�L��噝tJ�Y@u�N�>�0�0U* nP��a����O���'%6�����d����.]�~�DA�'�(�dA�A}	�2�	>=��V N�0HH#��P-K��@�J�h� D}
� X)�B�,wT�Ŋ�o��U��#&�'���c��6���Z��˼Zr��!��4/��s��
��ŐUG�+Pa�%]&RsHL�e@�<��z�˂�O|UH��K�N�숨��9"z
��`t���L&�����*r�١"O�����X0α����P�n�� �{�q�5�
m5�O?��Y�||6�h0�@�n��M��$�E!򤞎(;��Aw�= �MVd�
N6�'�Ev$܊�p<��'��hu�����|���mV�<�D�
,`y��9m�9D΁c6̓L�<� �R(R�\��G�P;p��3Pg�N�<�LC�CҘ�RPo��9�|a'�V\�<��܋z�)��H�$q�a`�<9��A�R��hv�K�!�4Hr&k_�<�5I^rd��-�`$�aj C�<N�B�D��2,2/~̻A�Td�<9C���8aVXPG�,{��[���e�<)�������	e$�&;�h�/�\�<�H�o�P\�(�e�\[5�S]�<��,�)l��ǃ�9!j0{ ,�Q�<ᒃ��v� e�&	�E�|�r�-�H�<1�g�!!�\,�(\7=��l:�x�<A�iB�Ab�� �لLO�'�Mx�<9��D�f��-y�řESt9u��u�<)R���qp�h`�=,Τ�B" D�<�DOX�@���1�@ 4>�1`��D�<�Fݦrً�Jö-��[�VA�<�!oάE.P4!�O�R)�X/�d�<��3WJ���Ŕd�\�)�je�<q�+G�(q X�K�i�fap��D�<��&��+ H3F��700���PY�<��N_�L>��"�P�(�%�Y�<a'�A8`�ҽ���҅T�椣���T�<	�"S�{yy��C߽r �t�aAW�<��G��?sTHhe�ӿ��@H$�JN�<)�+]�)��K#���޽�� Mw�<�@Q�f��|���:L�T- ��1��H�<�dH�� ��O1�:a���X5 ��p;�D!��a0O�Q��K7�JzH�"~�Ơ���(Xw�9�x�k�)Q�l؈�qo�u&�ӧh���i�x�*jRe$��*G�E������/�yR�.p�Q�,�~
%	)�S�j�*�u��u�Q'"@,;��q�Ǝ� Y7�PW�P�u# ��s	:�B�+���W��0�f0E�2I[6";2�r�p��3m��4e">�m$b�ya�d���+�ώt�xE�U����H�y��)v>q`��1~�����k�x�#&��n��y����OB��	y�LH�&C� ^��P��X�θ�4 �ڴEx�&�Yw~J?˓+�l|�� 8]Z ��@��G/���ƅEؘ�u�%Y�4C!*V-w��xb�i� v�6�Uæ���}��Ɇma"�Y &�=(��,al���$�0�(�b�'YX���R��A|����ɀ.2��>9�D�f�|B�OY$�F�X—QQ��"���O>YA�����O���1���*��㗏G�0�R<?����o?�*ONb>�J�!���H�̀�:�8@�͢F9���޴���E�O�(b����n���~B�� ��Y�i�t���`�nk�D J�0���D�Z�q����Ȃ�W;�>��&R��g�x2�$8'8ҡ�$����@I�&"�+ES�
�� E[��8��"��Q�O<E��h&Qꢼ�A܍�@���3�?���0���H>E�$
��`+�,�$gσ;�� 3u�dͰ��0^�|��}����?]0霭y�ԩ��[8-4A��B�d�6�ɶ���}��<Y��;�Z�����(�b�Cx((��'o��C�%T��}��O`DX�o6Q#�8�狪N�Zh��5�1OXl���Y�㥍�NL�}�T�T70ΑzAE;D�����0M���0�o�{g���9D��iS�'����ăA�p�0�7D����	IV�<��qo^�\�>��i6D��tC�F�Q"�\�,�R� 6D�� 2��P��b߂����� �D9xT"O���&N��=��iGKY�N�ku"O"�K���(5�`hd��j=H��"OFԫCW�?ĺ���g �D�B%"O�5JD�\ ����͑B�0�"Od�Uˉ�N�^A���e{e"O�yd���?=�	�sFӿ]�����"Ov����@H7��j���3�"O�  s�Ws��)�1 �md�@�"O�uؕ�09���䋈�V&�4"O��@w�h�xC4��9P�e2"O�԰b��Tk|�UCV(=@^��w"O��c�ՐK q	�����I@"Oژ���\�d�h�!e >��[�"O��S�� �v� b��5�Q��"O�L!�F�&�L;&!�	8ڸB�"O�9i����e`hMQ�1  ��T"Ohqxp�N��D���H��"z�s�"O���e>ߊ�	mS5P�T�y�"Očz!�έ�N�p��*=�@4�%"O������h�|���љg�
 #W"O�e�f���Q��(X�~��I��"O����v�x������d�̵��"O,DAf-�a䌈G˖��8��"Ot\���B96X���w���A�"O2���ļ7�>(�_� n�HQ�"O�2���f8������QL�A�'nQ0�n�E*2Ř��EL�d}�
�'6�l�W�9L6Fq�Ñ�m94���'<PY"�$'O�TЁǎU��j���'�ش�6���H��w&�z��А�'��pb��xi�#E�2yP�0��'�i��M�t��8�r�y. ���'�
E ��� !gn�2��5Y:��S�'g��C���~�b уh��Ux�Mz
�'z`iӑ-I�:'��C����u��' �h��iA�w�
=#����)�Q�']�� wbA�"GΆ3B��'�����*v�
PB���m�*�	�'М%P�����f\gj�1<��ȓZA$(��E���0�'�T�*t݆�	�mqG�o&,���?n~����8|lQ
�a���Յ��GN,���5�t���k��4�p��BF�7�Շ� �bX0����R�d�J�
�0VL��ȓ|�vX�'f��G;�{�M��F�Ft��/�0����a�+d-N�r� 9��`I� 1��=/����q�KATq��]$��9��Ӹ�a3�c��`�L}��F> ؈7Ǔ43�����1x8���2j������jp� B�Y%E��e�ȓ9�l�0�96�I�A(�"?�Մ�	�����X�o����%AVW�L=�ȓ]�I*S��A�հ0��Y���ȓH��)㥢��{��yx�i�<U*��ȓ
���x��:H��P��a�@����!�ވ���
�|���R��:ng��ȓ������%��ur���Z��-��]�`���ިq*Z��
e���E��l
@�%��i/��P��)D���@�H(U%�T�ܱ�j�	��&D�H9p�K6}���R��������$D�lSՍH�wC.��7�
w`�+�"D���`�	2Thi�E&H�?D�� 8%E(B���H0�Ӷ �@�"O�����8X�r�H,�0ZA�TS#"ON,��R�^�^4��E6D�F���"O��` ڈ�H¼LƂ�)�"OBYQ�jǈx[M¡'I���k�"OTi�j�+u�͑4�5-ER��"O��b��I��a�wh!tE^���"OX�"F�?@�\�҇�D�t�s"O.�	�
�"�lq;�gN�r��h��"O|��H \����bl�k�r�3�"O��I��λ��X ��6b��"OP�x�aA4'�d����D9_Q
��w"O
hP��*x�Վ"L��HA"O�� c�7؎L��_R���k�"O0a��e"sm�	4��@"O^)��E�a���S�N�2��-��"O�-��|W�P2�Q�"�FQ�"O$JbK�	�䰐SH8m�zA�"OX���E�#A�j@�4N�Y���"O6��T��0qj��1t��7DJA"Oh,مB�!&e�T�ͷ8U�U"O�,Cg˷K�Щ`A�'l�L��"O>�ئkR&>Y&����ڤ��H�"O�}PP��5XH[��M�HIP��R"OR-9ǆ� �P�pk��9+Ը��"O�L�ѬN��n�Rvi ��]�"O@�z�29�����ȡR��C�"OYz��J��Rf�_D���"O���G��
j,��rd~!�xC�"OL�24�Y,"��ȅ"\�-l�"O���2�X�w��
qG�t$����"OPؐ���,}�� �ӂ/&T�'"Of��IC�\�k5
�7H`��"O�D���H�~ C�)VT��Y��"O�����*T����S�/�J�R�"O��PF;��p(P�y5�:U"O-�6cO�d�	#����x��C%"O�L�5�k��)s���~��]R�"O"E󶃏��Ɓ �M�&]�0���"O8���;��c-�*�����"O@��2�� �jj����"�  ��"ON�x7O�A���3e+�QE��	7"O0i@S&N6X�0��7��30��"O���D9m�j�#�-���4"O�T��ڛ.�j�*0�΍G�1"OΑRK�yv"��4��4{�I�2"Oش��OU�^��a�؀mG�S"O��k����!f��٤"O"|����,�* �^�$��"Ob(3����-4p������	�h��"OD�֦�6@?j��OA8� @a�"OF�����LH�����h�d"O��D�J85��a��̊7��I""O�1�%4h9 ]��+��*�z�`�"O�DD,�1zI4�y�h�u���"O\���%C$�(��g�R���C�"O&鈢(ڃl:Dh�Ewx��a�"O�\G� �t�'̏+*c<}��"O&�Rw��,^+r�
$*��ӕ"Ob�!��[]h�s��ݒV�!�"O� :$�إ0q �æζh�8PI�"OF��w�@/���$��^��"O���V��D]���ҫc�X$C�"O,,N��%K��^�4]X�"O� J4��醣��]�s���#�Ru��"O�Q0cl��Re�a��.Аc�NI
V"O��I������F�����"O�%{T�@�4j	+���P�`"O�tCb�� 
 �� �k�/0M��)#"OH�ӑ�\�ql$}95�7X��r0"Oܐ	Ǎ��d�xPJtjI.d �"O\�C�G�f�4��7h��ԀD"ORhI��\����h�.T�����"O$�6�!1Xɀ��^�|ŐM�E"OЅ�f�=)�\��OH�db^�(�"O�s�V�*��]2��$V�X��"OҌP�$\�W�0i�U��85��"O�i�&d��Y� �C1��=�l`0�"Oȭ���+2t�9U [28 �؂E"O�%�H��.Ǌ����PBH�@"O��k\�z����cΟ�g���4"O�d	��)g+48�������"O4�ۓ��JH:�����!(��qC�"O�u0��M���rKu~�홱"O�ѱ�C�"O��)��(v����"O2e2tC ��ڲ��na:��F"OXI���=6Al$ &��QV��"O$p�V�� .���G��ȼ�d"Ox�[�@�v88CET�H�n)p"O$8�1ͺqިe���R�
�S"O~����[N�\|��T�D��1�4"O��c�T���1�B�(��4�"O5J7��t��Y�C������ "O�<`���J�`�!'�����ɦ"O-�s,׋9arY`W	X��(��"O�U�����Hpz�7�/b���*R"O̐�5#��2`����`�$8j�"O���ٳk�!p��(�YI"O����oD%	�9�K�na�Iӱ"O �s3&�[͂�"�d�*IX��"Ot=#�(O)��!�'n&'0��#�"O��2�D�#?�e8¢��u�(�z�"O>I��K~v�m��AF�4����f"OT(�kF�p��9���^�J�`G"O�����=v=��9�gB�����"O�U�����.	(�F��%��Sd"O2\A����P㺵��N�.����s"O�I2���4I��%߼��g"O�!kD�Ku���O�3m�\�k�"O�[BMS�cuF�r��ܴ`��""O��84�K#��Ĕ�f�B"O��H��9<f!p��I �(Y��'K'J
�mjt�+�t]1�'����E���V�A�l�=��'�f�j�&�!r^�H�3��%�L��'�*�bK�~�
�q��L�N��'��A7�eՊ���wvJ�)�'|��I�˱p����.W3}%�`��'v`�4F�B��X�D�2z'�c�'��t���-����pa��u�����'����l�_d~	�$b>m�|��'��9	&+B�7{�y�S	�Q��b�'�V|#���T?�\�󈖁Iˆ�P�'�0h��ď����,G��k
�'] �C��A��W.oMJ�h
�'$T�gY	��S1�٘V��r	�'ۢ�*#�ۛw�L�� ���La|Q��'�6e�Ј�.?����'�rU䈳��� Vx��g٧A���rR���O� )bw"Oey�   ��   �  �  M  �  +  �5  L>  �I  ~R  �X  _  qe  �k  �q  8x  |~    �  E�  ��  ̝  �  T�  ��  ܶ  _�  ��  	�  ��  �  ��  X�  ��  � � > � �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��I4K 4O����F�L��1d�H�P�2�p�"Oʉ����P+�2�
��������L����46k.��āϔ5���тL̩Py!�Ď::Bn�90(�3�l	ӗ û{t!��8L�f�K�Cx�y��J4-!�䗂K��d萲i�h�����!�LpF`���%_�	��m�!�d��.%鑤�;WF� �BW�:�!��"|.:Q�A%�/~KN�"V�Χ}铎hO�Z��&�n�S�� 8Kh� bQ"O�]�"��T�0%���
LH��e"OF�� ����yU�4�y��"O��E��`��Ǒ�:�>|B��O(��S�v���tn�<N^��A��t�!�D�\
J��ԣ��KV�!GZ=R�!�D����	W�C9!O��!��19z!�d��XMB�oҴRI��&&ͯ T!�$I~�-+t�ŧ	`�I㮈�B!�P��} A���Da��Љq�!�DӤdr� SF!M.Sh,��\�`e!�đ�� x��L/g޶���@YG�x�ɥv�DRt�H��n$�`�ޑc(ZB�	 [c~D�q"�%8�b$r�@��HB�*O��Ah�(�Z�a�tň�;��B�Igh��r���4*1� ��4S��B�I��N@�b�5Wq���S%�U��B�)� �9�wkۑoUJ!²dGtl��%"OL�X�S�TCN�Ba�]�Ql����'��F�O��7W"q�BIīWP\}Ȗ�-(�q��"i���M�>I�\�3ABܘ�ȓm�D��f$�:x&D@�%J�+_���ȓ�&8�@�e��vjĄ0��웍��s�hk�C��]u�$�e��� ע9D� cS"�&@�串V��y+��qv�j�`�	[x����P�� ����O��j��,D�d��I�?�$M�)�'�}� +D���aީM����Ê��2�@�X�*ʓ4��ʧ%O��21nM&-d��#��^T��v��j YA�6����X/�	�ȓk[6�KG�&'o�h1�.O�T92I��x?LĹ���g 9	�	,.n ��2�)[c�� ����N�)J�ȓxJ�=PU��BRܵ`gN̟z�T��=��\�TH^�U��<(D'�zPz��?����~�d��<��ivj�)�H)h�K�Z�'Iў�v2P�AG�>W@���
��L%��D{��,N?�~@j���k�j��#���y�A��Gl�LHC�#��	��FJ��?i�O���
�,+x��,V�:�y�#�J�rm�{r��o(8D�ҠP?��X�L]hY!�dR�o�v�x��K�`-�$ba��^S&Yn^��ࠔ�_��u�&	C�h��ᩰ�&�l�	�m-����Tj��W���-8t#=ن�'����,ʸȐ�A��^������hOq���de�@@(O��PP�I 6��oڮeS���U�&�V���oz\�8�f��1O�扷�~�<O�c��xb$j��M�R�͟+˾��r�?D�\H7Ț���Y��o�|b��!�&>}R�)���F� �x�I�����5$�7V���$'扬&�v�Ƞ�
�v�S@F�'�B�I�n�$E���1ml�p	ïE�A6L�'���3�)�S��,��UhUJ���KY&�FC�	0T�aʧA�%���0�8S{6C�	�%\PX��!ֳG���A ׵tV��Ĥ>I���aϼT �JQ�9����r�79����hO>	P�o��,	�O +��Hp#�/D�`���iE${���3���,��9�O�=�N��,(J6i]� ��"O�X�0Oͷ�P,�ȉn�r�r"O���$:�{a��+I���v�	I>����9AM��f	<Ѹ�
�k#D��pm�:9�	�wd��}>�4Bga��D{��I=r�Y���9j@�t�FF�*3
!�Dº>�	��^�I5�'��7�!�L�D�R�8�l�2G�XZ��*Dv!�[3 ~J�a@`�SU.h3Á�:q!�dƶl��A��j���irA\58!�Ď �(�bv) 9��Ёƈ�i�|RR� lZx��j�JU:�VP�!�B��
k��F/M���I���C(�C�	�Jb�L�kÑ9G�-�0���`lC䉔�6��1���{�nu���&�➌D{J~:S�"[Ծ\#1�@,j������z�<!c#ͳO����E�- �N�~�<��I��`4�SF�'Y��a1�HxX���O<���&ޝH��R�Ћ=(l���'��$S��(O���U��;y���.�� b��D+�S��ۡk��][c�׺I�0	@R�$=��',a|�%A =�d�����tD��*��x��'+֥!!�� V��QH�{9ph���x
� P�P��5U� PpIۘ�n<+C"O��Kp�PEl��@�H]�VI�T"O�T pA��ԛ���,������>����)@�a�`A+�jh۷�>%�!�:78���S/<8^�ڕd� �!�䐢I�N���i��s&<���{Y��	l��~Zc\X�32�|�F%#�
҄_�:���'<��1l]�!�0�
+Y�⠫#R��&���4���yG!Ÿk��-P�)��͘T��1�yr�z�$���������Q��!�~S���<���dLDE�1w�R-g-��B"ĉ!!��O|�b�aV��2�o�l]ĐxR�'�쨘b�]�O�̩2n��N����'����bV�zq�R�%Ĕ��'���z��ܲ(��$"b�6u����O^���>m�J�b�jՉP8uIa`��7�t����<ɶ�A�,I�a*�	�m�i���Pm�<�īQ8}��H��T83�V ɔMC`�<q%�՜D����s	��(!�Y�<�V(	e2�}3��(x)Bt�$V?����pA�\��	S"3�XQ�g�
?O��I]؟��6��$^�v��A!	!%��lз�%D�A�x֮AЕ�q!��Kf8�C�I� >�Q�n#6��P&CH�C�	�0:]���Z;r����H/0����-�ɇFP��ˇ���'��4�E�G�4�ȓVUʰA�C��B� @z�N�-�̄��A��57����͝m��4�DjR�,V���%ߨ�@ Lɲ ��a'��K�
u�ȓ/=����-Q"��93�*Y^���ȓ>��QӰmT�2�MR�^�0|�ȓmfh�riKX*�q�T�Q5�Ш�ȓ^n��Ӱ�cO�pzp�Qb5��FS-�Cd�}�Db�!��TA�ȓ)��a��DL�!��U$p��s�Աǫ��TQ���_�nA������PF��\]f�����uG`�ȓߤsg�[���t1���i�Մȓy ��rg�_���wJD�e
,��� P�ڵiW�A�6\��Y�<��|oX`�Q�Ŏl��S �ʎfr���
$8 !�	X�މkҋC�julͅ�S���O���~]#!烆����+W���CfM��4���W@��� ���&��@��U�rI[�W)Z�ȓCD�� �
�.�����MI�І�[q�ř׫�5Un0��!7����ȓ[��Ka���i�\x��Ϛ/�
8��&&z`2�A
?:�L�z��' |$��
��h*��H5:|b��C�܅ȓ,����&F�%��(���L` ��	4:(�Dg�j���e��A���ȓZ�8�g�ȸn�08�ގ쬹��*m��	�.H$y���	�p4��
�Z���fȸM�H�0F�@#\9���.i�aǘ`1ȁr �%"�~8���6�0A���6�(8����g
2��ȓy��A ����6݁$��3
,���4�Jt��0�1�0�^Gt`��P� |�À��'��T2�s;<<��@jw-^�M��=:���9�Le��X�H�#�*�*�0\�fD}EzQ�ȓX�^���k�`�P���ڍ��E߬����6��0@R�̙w�� ��S�? ���J�'&�`��ġ8L�Z"O0���@#n� ����%fKf��a"O6�S� (y��p�P��9H�D2�"O~���ΊY�y��B��6��"O��K������U�L�C7�,�'�'�B�'�r�'
��'�"�'d��'��𦁝�<t \�2K����@�' ��'��'Tb�'P�'�b�'B����ꚯSkF0��+[��4��'���'���';b�'2�'���'�J,Kb�Ƞ&��0B �*9"HT���'�B�'c2�'n�'�b�'r�'��$��e�5T��D�R�3@HX �'r�'_��'n��'p��'H2�'T4c�a�R�O?�n���4�?��?���?���?1��?y��?)W�[85.��{W��U�ņ���?���?���?���?����?����?قJɝ&JY�p̙�R���l�
�?���?9���?����?I��?���?�Ipe^%�`�S"Z0@��?����?y���?���?a��?��?�@&P�!2��N�ڽY�N��?����?1��?���?����?	��?��/�{A@đÁ�M� }�����?I���?��?Y��?!���?���?9v���j�b�I+I5�B �Q�١�?Q��?I���?����?���?����?!�$P=u5�hPt�BBٰ�̊1�?����?����?���?���IC�f�'1rEQ���́���;�h�B�")��?�-O1���3�M�U���9�P���A�_1�6�	�J}!�Oh�m�E��|��M3E��VZ�Ґ����s�/S��&�'6��0�i��I
}X=i���T���.�GA��d�F�0@��K�=�<���d<�'����$6�$Xp�ٜ�<p��i��Ua�y2��C���{丢c��3����"@�n��x���M;�'Y�)��.\�6�g���j�i�8YJG�P�L��a��`k���bӰw���뤪_V���4�'���X�ʟV�~�*m��*h�K�'��It�	��MC��q̓^�\�:Cそid�ɢ4'��a�($����<����M�'��	�7��=�1�B[�n��#`�?U���z�� � ���|zB��5�uW��O@E@��+A��i���ť$�vlq�-�<�.Ot��s���mĐ.d�4�g�
[R�@�@x� ۴�'l�7� �i>E�U#�M��yy%�N?���wo��h��릡�	�w�ȭnZk~2O�*��ųW���t�Z���E��v�8���F߱1����|�V��Sܟt��џP�	���M�$4�`Ȓ)X�I����*EYyRl��pv��O��D�O �����B	|�.,
��t��U`�'[5t�:��'̆6���qϓ��'����E�x\JPN��MRh�3��Q���
��ܙ"�@��'9P��k�0oL��q��|�'Krlь�vA���V<*$Zv!�o���'�2�'O�O����M��m��<a��  ����O�%La�a�Dؼ#����'7џ��۴O]���w�(	��J�Ԇ��u�ץX+V�R���bK&PZ9O"�D�-8�`�GJ$:�����gU�C*h�sf���� (�@�v5XX�d�8m2t��HdN<8���/~P��eF�'3L{"��U0���� Y9Ef���p2H[DN�	�� C����\+P��7�DX���!�	5b$�i�Æe4$!�L��������H ���At�<�a�����x�$��	|%���fT���n�g�H:BQ�P"`�����~Q�0'��=,��e�ԿJ��{"���'�r)3��[d��"G���MK���?��
Ǣ5�a�x2�'ur�OtX���T�q�8��b\��z�"��DW�8�B�O8���O
�D����Mӂv�J���n� V����ָi<�V.^��O�)�O*�O�H� 	��JN�vsa��-|�I0�b�h���<�	xy� �&8`���Ď	f���i� ���H/��O��D�O�ʓ�?!��ZY�1��� � ����U��rC�Eq��?	��?Y(OnԳT���|b�����, !�ȑqlX�#Q�[@}��'��'��۟�I�c�>�u$�}QQ� Y�\�W�� �U�'���'��X�T��͊#��'j�R 2�Ď���Բ���~�ip�ig2�'��	ß������c?�%k 6+�V��%�5�h�R�df���d�O�ʓL>�������'E�\ck"�{$#�#mh5�EhP�:�I��4���O`�d�/m�>A�s���$�@�>��%iF�`qr(�e�i��	�O�$��۴x�Sޟ������#g\���bV3~#�1J�këe���'6�a/e��)��g�I{���r�U�PڡV
��6-[�TS�nҟ��I���Ӻ���|"¬B�1b(�p�פdآ�	��'SE�����%�	蟐�I�?c�p�������/�T"1�5+��$9fdi�4�?!���?qF��PΛ6�'���'���u''Бk�}�d,�	��<#b閚�M���C�-��?U��ʟ|���k�q��"��6SD��j�<$ �b�4�?�`Y��&�'J��'#��~��'�`�h OX��IS4j�7|�8)J�O���d=O��d�O���O���|��E0	���Q%YDt���+�
f�v9S�i���'^��'���'���O�1�� ��<)����� w��;7���O��d�O&���O8�'Cg�`p־i�� ��ܜW�"�+�:&��p���w��$�OP���O^��<I��?���'y��%�C*_ H���'�V3T� Z�����(�I����	�8\Zhڴ�?I�=�� ȸ*���Am�,�D�K��i�2�'��_���	$^��������;���;Ç�%%ZM�+��l1o���	� �	�p��a�ߴ�?9���?a�'p��wk�t�"䩖8�16�i�R^�4�	U���y�i>7�ߞ
$����Li�[9ҀU"IF�FQ���h�%�MS��?����z�P���]�88��\�DV�y�Ċ^3֎7M�Ox�����q��'Uq�
�I���,w�$,�=T�3��it2��Dw�H�D�O��d��'z�IgB�I�k�?
��X%E��}���ٴ|������0L^��?I�S�$�xak�M<t�ee��~M�ٴ�?���?q���0�IRy��'8�I����f�T)f�:�)0 �!V�'�2É�G��Ú���������OZD��i�#_D�	�KD�n�T�S�@A�����1Ybi��Oʓ�?I.O���
h�'��Q#ׁG�jL���^�TYar�\�����	Ɵ ��uyr���D������	(H:DS���P¬>q-Od�Ħ<y���?��5��!�qc�� ���;*�4/���zf��t~b�'[��'{T����fՉ����[�`*ʈC��\d����$����O���?���O��DF|$�	�v<��s6�]�!��(b$@���L��?���?.O��#Ĥ�V�Sg��S�^1)���Q��-z����ݴ�?�N>!��?�t��?�M����d��hf�Т�}'�]���t���$�O��I��]��D�'^��e�	qN
� �+��ya��M�Ob�d�O�Yhq��O�O���6ɶM领.Ub��Rl�F��6�<Qt���h�截~J������X���=��)�e$I�!m���#}���D�O��8F��OO��f�+���L�H ,I0R1�iL�1��iw���d�O�����&���I�wsD )A����(9@M(�$mBݴr������S�O�R�	!�4Cl�*3����b�>m�n7�O��$�O�E�R�m��?)�'�Dܺծ�;>�T�0��mK����4��,�4ɕ��T�'{��'�n���ǁy���E�/g�:��E�l���$��|�L'���	��&���B���
�/��a3~��E%����#*��Uy��'Y"�'W�I�����o.>����ǒuG�qӂI3���?���䓦?��#ƴ,H����@�nJ���x��UU̓�?����?�(O�X�P�T�|*f��/s��x1� ���1���R}�'d"�|�'eb	v���$HlL�t�*m��Y#2� "N�*��?���?).Ov��QmOq�ںCѧ�Mf2`���Pۂ�3ܴ�?�K>q��?	ӌ���?�N�xؑ��&e�<�Lյ�L��nӸ�d�O��P������'l����B��EC�IF{&mR�(�m��O����OPl�w-�O��O��O�6����8A��y�Ŏ56�6m�<)��0+�fa�~����ʄ���!��v�м��)L�G����4oe�����O����H�O�O���IU�G�g��t���	 R��<�g�iC���Ɔwӊ���O����(�&�����*�̨�tnˣ~��M�6��.f�F,3ٴ�&�p����S�O��@�0�Ӟ;8p�ZtO�hNq$Dͭb��xP�I7~��� d@9�O�#R�.<���YfAN�S���'i$M�.ȸ;��Ul�4y��9���ŗGA�0[��V�N��n�. �&��Ug	�/!�`�o�:e�������SNP�Q�:�
u�4��/�*y� �����yBs/R"G�x��+��N�yY�(�.�j�
���3�zٻ����aD���5���9�̆�:�j)�'���DXY���?��?�EKʖ�?!�����N6o��X(���M�t=��`U�O�hD��D���Wi۫a������@����@�[�xA:��ފ6���㥈'�B�����?C�J!��C�']�`r����F�	�B@D��C���౨�o���O�d�Ob��'R�y��% ��5*R�S&Q�ȓ`������'�d�˗nV4���̓N���qy�n�?�$��?Q)�ji@&A`[8���Ťv����&/)8i
�$�O����[�!�d�p�$q���ʧu�HT�u���LB��(Ĉ�"|�"\GyrJN)B��Ԁ���x#J@Y�����d��8qڲ�e)����(OP�p��'`��ɀ2X�R]Ч*�Q/�Ar%����O���D�,�T!��!ڼr�8��6f�Jua|2�3��ͪ>���X �P��e�#�_k�Ě�/��pm��l��^�/4I�2�'2N1!;�S��L-~��<7Cv����/q�d��n�k:�£~ʌ��;>bu`�oW�B�zx�o֑d��]�\�4���a7/��m�����k��	�����w�,��5N��I��9c��-	FMmڥ?�$�����Y!.O����O�=ᔊ^~̨����_=VU�t:O���?�OP<�&�7�|�qQ��<-�ID�ɬ�HO��)�Or�8"(_&(�B�Ц�Y.= ��1%(�O��dC�$X�b�O��$�O������?Y���k����J�(sFFe	砕C?�5�,@͈s`G�3�����C{���;@�O�C�jh �ǖ��D�B�;TAJ!�V%!�m�Bi��L�o��I�BD/zVE�d�n �I(�Ms��i��Ol��OQP4�a��$�J2Cn�)�&a
�'o����kҵ�܅K��BE���$ғ7���yyrE3+b�7� Z�n��]؜	C�f���Ն�OD�$�Ol���d`N��OR�ӞQy8(Z@ZX����� Χ�6��U�:�$�;��\�|����ɟ��+�CR�(�u�O�aʴ|PQ��\�w�ܷ8�$������ĕ���� �Ƽv0���m��f�֡Qe�*D�T���W�~=�a0�ڙ��$)D���$Eړb �,J�@�L��h����4��#��굳i��'���O@ؘ2�ɘ	���u�	�A��[�Eϟ���� �-�%QL�1� 9�Ȁ��4"���(C�S��J���������4剫z� bP+��Z��}�C�MŦ�h\w��5؇�\
�*���G��|~6�w��(O�qq��'�("}Beo5V&I���S|��e._f�<�7��R.d]�d�C�.�h��d��CH<����K��	CKF2f��0����<gm�8����'��_>5	5�Ο,�I��H{"�%���p�z�:�(�φ0��0R /zt��kӦ	5R?��|��4+.P���WE�6�`��N�|H+�%Y�Sk��QUȟ�<� �l��Y:�>�N�	v{z,����l�L�:�OڅyO$�h��O��m�ɟP��g�S̟@���Њp$�B�}Ja)ٰZ����ċ埰�	jx�h8Dς�*ȋPoėg���T�(�	ן<p���m��dD�E��`����&�����֟����"jL������ޟX�[w�r�'�^5���7S1|�7�E2&[t]PRy�\<�u��4M�va⇮=#��m�ޤ��,ve`��H�xY�	�1	Z	�d�%���2�F�?EH�->��
[8��K �"��5���0A��t����O���BG�	���ICy���?d�.r�)�.q(�ؒ�*�����2�O�E�#B5,�����Y�ADѪbn�Ц��޴����������<��AmZ
d��AЗG�
a^\)	W��+"Ƹ��֟���֟�2ōȟ\��,��D�68�4�<,Jj�f��';!K%��R��Q���<�g�Ia�>��c�`ƞ�Z���{�)R+B *��95�G�%��%��a�D�'GhE`�S�����C`�X�A�ǗZ h����h�p6��Op��?	��O�R�В|�ΰXgI@�V�-���՘�y�0v���T�K�<�N��OI<�y��zӄ<mZKy�RR�7�O���|zڎ��anW�R(�y��HZ�u)H�(���?)��C�t)�ԅ�%���BiW�bO*�6QbC�>�h�0Ѫ@�%��!�I�%=ҁc'㎇>�41���T�"��~�9d�1�>VR%$� ���Dx�'L��K��?����?�)�PY�ab��.�b)��%�7P�@Y���Oz�"~�kĂ��@_�j�F4	�'�pRܙ���ē8U�ݒvBJrZ�	� ���B��I��i�r�')��k������D��2��!��i]	k�)JէE�8����)�~�va�󡐢cX�P	����.�����c�)�D�sDL��10ՠ�Ƙ NY���ȉ'}�abaY�nT���僌�q�B�+x\%��!��:ā<d 2)���'��7mOFy�'��2�2@(.�1�Q���a�s���y��'��}b��	�]����G�/��8)!a(Xڑ�<��ş���M��N����@�s�`�+�*�Ɵ`��39��)�d���������x����u�'0�̜!�L��c��t�0\; m�+Q_ ̹��Q"8�Av�Ͻ'�$[�Oᑞ����W1\|t�#ס5V��,�l���4�T:rsz�R�G3+���ӿ	�4��@2)۳g�0�Y�g
���ʺ� ��O����E
N`mh4+
=a&TX�l�Y�!�D�?~v����]V@��./�ʵGz�O��'��Awab�d�[e
KPf<0å�'�~���O����O��d�$xm`�$�O��ӕ�Ҙ���U�yX�M�Dx��S5g�"�l�{�'�g�D���	61��-z��Yg�LE��	 "!��%��W�B!��'Y�9�p���W����O��VsCȑ���#��3���Ob�d�<9�����IߪSm��H E<MX��!��)8Z!�D^�o�6�P�/�3���P�1>���!�ItybfDp�7��O����|�'��U�r��'��5���2D�ш)�M1���?Y��K��Q�A��g�`H��B�ћfY>=f�P$_��)W�!�vt	ӣ �Uب`%��?l��"ThN���t!�Ë�uW.�<��P"g��1m���a.O<�(O�̳�'��6�\�S����RN�jRN�s�嗸k����j�ȟ��?E��'�P,���l����ڢ<�T���O�!D~�(yӰ�l����ѕ��KsR �r�
7p[�3It���FA�M����?�*� ����O�d�O�xR�&Z,h��<�+)3F�	k���UlQ��L�*J�(S��P��'���?��EC�|o6�#F��,�H�B*Я��`W�Ę�!�����'О�b���Cͤ
���5��)v2j�l�m��� G���0fr9�H�[?PZ�TP�H�ϓ�?��Yb�[u��h=�W�[�UI�DxB�6ғ��M8��(��ҲrġI����$B�)� �|hċJ+1 ���� �h���"OT8�5�Mn� �ط���i�p"O��b�A8sE�)�,�Y6N�æ"Ol��0��okf8PFm
�JB�s"O:=���܀cNl)W��X��"Ob��Q��#-M*H&$�El<�0"O����	���z��ƶ5^.x�"O�0G ނC�Rpq�B��kD� ��"OH�	�͆㔍k�OY�a.���"OP���L�d�.$K�m
�H�@���"O�d�D�N�p�C�	b���`""O�D!¥^/��R��0�႗"O�0p�Ƒ� pҌ�� q�Hi�"OHT1���_(a8�@��O�0��"O��j����d�⇺M���4"O���ӎة[J��R� K��0"O6а��5^�p���M�"O��Z�� |�Աr�A>���Ғ"O(����M[� ��Gc�"O��A2��J����4��o]��H6"O ��҉̵�b,�ge0H���%"O d����y����p�Țd"O��!���e�PJTcN/"U!f"O�$o�i��)��,@��5�"O}2RL�;M3en�x	:�c"O�]�ǃ0�0A#mf�FY
�"Or�����.>tf��1Lӻ2�m��"O���a�ĉ {`��$zv��"O��� $�!t
����nЇ^�5�%"O\2@(AcC�/��I Ȭ~�!�d^-7"$I�A�eɠ��̀?.�
O��;�*I'^Z�DA5�3Yú�c!�I��yŨ��'*wB�*� L*G�B]��,ݦP���ȓn7�t@�eJ;�,�Zw"&K�h�'�ڨ�۴5��`@���"}�t�M�l�"�e��#c����G�<��A
)[����A$U�zi�M0Gj������ٴ~����S']�IfH���g�'�ʜ���nV�`J�c^/I�"�?lO0$�5��!��ٛrgnѸt��2�If�W�rh�H!�K����+��M�j�B�+�-�칊�a���l4�>Y&�[M68����6�h��"g��-##~X�'��>z�0�0��?yC�C�ɞ\DFT@#�t�)��B���n��AlT%4���D����d��a�6�g}2i�:��5���T�_�8� �@�-�y�M�d&i�&g���ڰbj���M+�d�M_�M�A;�L���'�ba" �p�z�aw�]�Q8)��I>6w�$����d4b` hJ?H4��3����x[G�s����'��݈��S����j���a�N9��{�J�2'L�p�V�Dڝ�$GW �-c�Z?�᳃T�Fu��bF:D4�싓"=D��h'���G��!�`�2#�Hӥnʨ6�y�	?��+7��4Yb��(��$E���ygɚ�1���I�#I������>��'Vl�����a��u@�EK��,�g�<Y:�YV=O^5�� ߂1�V�����!]�t�b
S� 8����A�j�kX+�HOZH1��B�H��� B�T4�1�'����8A~�qEB��ݴ���g��z���`o�9�����'�r]�d�ZFZ^pR6��D�T��`�.d0W�m�8(�����F����j� ���5F���M�Q��*m���#v�.#R!�dO�EYPܠ�ΐ�PM������(��Y��m�'����� 7>��h�!�f?r�����W�N�Eq��1�C ҙǏL9$��B�Lb�9�� Qwk8a٧�B�R��[��[ ^X3v�x��՗@<�b�l{4\�UJ �ا+l>�<�`gX�;	@�H��D��?�fC�!��ĺ�T�T[H�)����K�Jv�O�����G"&<� �)1��'٪N|% e��1Mbޙ��	�1O⩩�ڜY��vk�h^�1��iz��]���E{J|z'��Z�0� p$��Uq=��nȣd�a{�"ނG>�,;�E<A5d,�#��'SO"�p�`&����#5<O"�r�h\G���+�"y�����_0��m�C��w'�)(�.��)-�
9�w��:���Q��'����O�����%I�Rx�j	�:����0H?'O0[�a�8V�N	� �B*�Z,W�� r(j�	��@��0�KB��$�C�&��6��
�f#A=$�heG���^�4��yࠡ߫]�I�чk�Va���5N����A)��>I|�"f�p���zC� ����Gwn�@!FKC�wD�k�(y�O1��1�''Ԝ�0�¬O�p�",�_�rQ�ߓmB���&~�ԝ�t�U ,��uh�])RШM��Þs�Z�I�<!�i�7��I�Ԣ��uGej>7���R�n�R���#.Z�0�i)�I]�0,32D�R]2�:�!���OSH0a�G-@�N}���e����L<�F�IJ!��'��p�m �ب8)��&�F�y��p^Q���cxk�e��H���S>}Y���E@�3�2�#!M]2���ѓ-:����k��sJIV6!j�*���l?V9��p�`d�N�b����O��|�B�do�� �)]�C)ؼ�����{��ݛ9>�b�F�d���
B冡<�ĝ���ʪo�8���`�n�'A̙H����"�x��)�%�PU�썰&�R��X(�O���U:���$
�;!�$M�)����J*[ X��!�)� ���c�%@o�����5X�b=�&�Z��Y �ޟў���1�p�$j��u�j��%��p+Q4�7"&XXs�F*���O�Y��x@��:� 9��k��%S�.�x�K=�����weH�h��c�,)�ʕ1s�<��&���2���I\9R����0^�m�TY�NNf�RY�5@;O*m���ڂ5�b1���ʎAZ�d g�RDv��+E
���U�T<�I�`��b��P�Cg>��3��;v(x#Q�X �0I�,���Jb�O�PWn�X��1�̐�!���I������'��c�.ϷRr(�R�ӊ$l��k�O�)R����U���ӊ˃?���R�A��r��ZFr<Bf�zjrhr�
G�x�a,7?�g��|���]�N���a㥓	~ R)�R��&J)�����;v�:��dc�qJ��9�i�`�0|X��`���W����ا�O�
qH狎_s�#E��Ҡ�FP�G�#?�7g	:Ƙ|�-z 
<xq��Ϧe��^28]P���E�J��ifͽ<A���75��pu���.����Ċ�lߛ���&@���h��p3H�J��ן��ԇ 3T��E�D�}>��X��3`}��|�	$Z� I��F�J��&k��)�@�'znQ�d�[�Mj�: �dz����./,����@F)��g�^'Xg���ƪ��!�
5�'0��3�i>yb�	W�n�JȂ5�	Ҹ "3p^�4�ড়�@Mc�&`��k֩J��䡲�`
�If C��,���J��c��'�M;2�>����0�Nz��Л!O�L@8d��ɤa���y��μH��e �)�gXv7͟�)%����D!N�(e�s)�Q����k��P�A%ӏk� ��E*�S��@�i���I��X ��$	�%Y�P��#o�" �&hJ�'ٲFr� � 
6?��M+�@�(w��B#�i�Z\8DmR�2���	
Xi�h�P��
S���q(S�{�B"<q� X
:]���1�����,�����i��.�vf�g�I#?;�C�NG�U��0;�#V�x��`tJ)	���Z�E�S�bĉ��'zj��֠�[$Rt�!�-6�5�!�*�zкA*U7\">�`'X���,�T�#�=BL5���5ⷪV���DirC�7}вH(��'5Z�R�/Z�[Z�聒MR!lg�YQ��-D	a��BК56���͐��y�� �[���
WoK�
��)�jj�ceA�
m�̑�A�T�0�C�rn��e�Pt9D�LLqʸ{��R;i��`��M����4t_��j� $I�B����%yQ�'6�6xX�jB	ͷ825 �ɈW|	y�� fq�z�Y�fpތZt͇�X��'H��?a*���{7b�%?�h���턟 X�)#�5o;*�ւ�ʦ��ۃr�ayH+:����G$�,j�UYj�������(�Ijy"�X2~�a���0)| s��?y5���:���U+^�(q�fY�'�T*�� g/Z�XSM�#u�Ƚ�ٴ|�>Tp�Y?D�d��f��#J�E�'M� 8�.4t�DSV'JަUr��̧J��]B���c+f������X�h���OY5��lu��HAC5t. �w�<E�� ���H�B5x��2lT�Q@&Q�@��j�&��DF�9k ���L�6����Ra�=䴝��"}B��x�OW���;?hz8�aߣa!��20ˀ�G�"���I����r���< A^� �%#^�pX�ы��~�X�'�� ��m���ӯ���Y��P���cۿ9��T�������F~b�D>X���!�ڿE^L�`@f���!�� ���W$0H�2Ģ>YH�<l>"(���i�,��%���HO��1���Tixx�#V(�*HQX��H���^1B 2SIʨ�ȍ��d	� �<˃*�&����� Ui�1v��|(h`�?P?� R	Ǔ b��� ^+��� d
�/
��
&�~�� ��'�dx ̣��!�,�9�~4QTE���>i�0�8���P���Z�-R�L��YD�'�d80�J jל�YҠ��gH܉0b�8�)h � ���O�<A��^�Q#���TGQ#� �jԺi6HД��1�"�{0Eŝh���:��$ʻ�m��!WH�D��h��{Q��Y�� &�K0;�|�C�6{;��9݂�3���=R����e��t@�G���'�Tag!��4ڬ�צ/�V�H��V56�¸H'��4�*��g��t�j��D��J�<�%f��􉍓
T	�LؓP��Q ܴv�.�1����<� 
���Y�g8�����v&�)P��a��|�H	����!��L�3��?Ό,*�CǺd����O�81���.Yc�{oI5L�ves�-�0K����o�v>�,���Ύ,��Db��q�����w�ԣ��XY|�Z���)	ʨ�ʫ>�#��� �[z&���O��\����*?��Δq]ܑ�u��,	P�E9s��<��	�*Ȑ�H�s�0ع�Ƅe�'U�\9��4��2AƄ�U�.�SSmߵ۰Ag�_W�LIZ����0<1p��3?���jԎ�.���"��\CǺ=�LX���Ŋ���ybo��?Ԃ��ŉY(V�zMXq)�$kv���Ʌt���]�r(!�A�%�@ܨ��PX�����dC:��bf��^�����&^�bȚ��E�'L1y��?0}���N,��|��'o�T�A��HFK=N6�+"�M��O�䝰j5������l��mPSL��0RkďMż����яa��jq�E�S���ۊ���A�V�Z�;!gԯE���O�=Ju���u'�%7�ʰٔ�,?���^��h�c�!9}��ȳC��Q�'eb���	P�v|0:�h�޺X�Q&V $j�|R�I"��QJ��ļ k��i�NS�	
�$����H�	�n;,O�;�J@�@D���WaN�?v�d��K5JAv��f7!#X)$�θ�c�[�'��6�-YAJ �r��?#��	�B�8j2�cqÎ�]�4�*��;@ң<�'����eO̎7�t����Ki(�S�i�>G�=�։^�z��p:f��mK�Ru��p�^[��3��؜gV:��?1֩�4@%h0��e�3S����$��0#�Zߖ91�2���vR �FzR����ި�nZ>6��!*%�H�j�+4�@n��a����MӃ0O�T�I�]N���'Pj���2և�0ED����l�>��"9LO�x4P�c��uQ�E)E	5�1O�D+A=u3:`�C�\���|�_?V%0�F0L(:|Q��F�$Mr���(��`@�離��%k���_+�����DQZusV�Ԥ5&�\�
C:x� II�E'�b*�����������d&��JJ����J���rc�����ٵH�>10��>�̅0WA�����a}��*�0�I��$b
���Zl�.<��p�.�K�J	?�T���йd�0���ҝ$ ���(�>��Y��
T:8��ih�.|�̠bt�\�
0'��k����d ���g�*��dt�=Q��q�%��� mڵ����A#�I��E�6dXV��>F�L}��I��`˧*S�<�ցkB�1 w��/t��t�ȓ4b0�`�ȫsp�*c��ACN�ȓPO��iħ�@t��ս
f|���<���w�ΧL���XD� �ZEI�� X�����ýoq^%��K_3ǰh��{t���j'��M������ц�G �}:"�C:��3
�����a>R��3GU08Isl y�ąȓi�,�x�(C"u���2��Q�3|���ȓs5~�ӄ�K�o��݀cg��Gt��ȓ6łmG�ĕ`�p�XwlՍ|�(y��O,ܸ��ְ���ʰ\�q��H�-�$�Np�ԁ�k�0ow0e�ȓ4̄R�F@� �aD36gX�ȓu��Q����9:j���=��8�ȓ�����M�!JLCՠٮh�h��8n�x�����Ls��*aV�݆�;�Y��䔙czf�)�H�x� C�	9#�jr�Z>H8i�Q&S*U��B��7W�����9R�"��oP�Z~�B�	)1w8�c4�E_'IaaВ$�B�I&�l��e!˶��j�g��y�!� �:^e��F�h�6��"�?~�!�$,U�кW�P��va�����!�$���в	3&Ю���dUR�!��0ZM�����A�b�A�S!�J�\@���>�-��жn�!��5�T};�E�vi�H �+ZT�!�Ĉ?Q����;i�� t�!��P��>W�C V�G!�d�-R8^p�[�F)�f۳uilE��'��	G䇋�.�x�I�1a�����'�4l�d��X}��#AHT�]�*Q����  Ъ �%s�]+�K��$Y	@"Ox<Ф�р��8dm�,m�F�S�"O��҄���E�NA��,_��̅BG"O� �'%r������2N�P01"O>-87G�^_ mcCW2��P&"O��`�	I�8m*mC5&جg
���"O�	�JQ�}��X��o�=
�"O ���(�9xڈc�fV�B2�KA"O�q"�F�7<��y�%�7�֨k�"O�0#H�/^��$i�Ęj�"Odm�D�Ë|t���3��g��%�"Ob����c�J��4aX"����"OLɘ
�<�0ջf�.N�޵0�"O�M��f���-	 lD�j��lK6"O(�j5G��@���ʴK���j3"OƩ�$EB��f��=�p5	�"O�Yw���E6��b*)Z~��H�"O����R�[�`��hE;cʐ��"Od�۵-rpM��F7+R�|��"O8\���^:d�2�a�N
6G81�"O��u��<\�xF�G�}x�"O,�1ĄS0��D_�P�Z���"Ovxe
�(T䃤" 37�ɨ@"OH����5Q�f}��߆@�Ra)�"O��j'��N�����@�(u�s"O|��2�	6a��l�˒Hf�L &"Oh�Wf�n]0�ڡ�Չ\H��"O,(+�#�0vή�2$D�4r����"O�e�ׂ +�h�S5i��e�"Of����s���s�^�k��#"O��IҨ�4�~�HC�H`��I`"O���5�	/	�H8�.]� �j�"O
� D� �xT���c�@� Ac"O����˺yF�UQq�V,(��1�"O~�+�ۅ�E�q�x���"O��x`Iǚ?���gc����C"O8���,�*�"ɻ0����"OL���!��#��+�2�Z�"O�ib󬅃-� Q�A��
��m��"Od�;ټS]-��'��[� ]k�"O��`��upl�����$p����
O�7��n1ZĦ�7hp�57
�2G^!�dY�qފԱC�la���N���I��D5�q�Q�0jC;J�q�NG��)��p�u D _)�ڰP���y��ȓ*�©���sV��� �k�e�ȓ) ���G�
cN"豔�#2���ȓb�uh4O�,��ڣ�͖d��`�ȓh��	��(�%1�x��KؓQFՄȓ�"=	R��#�.� .���h��� �zly��S�$"�	a���@@�ȓ,�X-)�
w?�-Ba�
#���ȓ	i�����`y���+O�V��ȓ�N	����O 1sÌ&1����ȓzJ6�5o&�`!)[&})���z6�}���^�rf`�B�D,7���z$1��%��hD�᭐'ʼT��,ʑc0�^�l���5TM��b8̈���c�u�[A<ԅ�SS���H��b�& �s��gF�A��Ӝ��ä��	�@��AP����>�ֈ�2��1�≅�M9�4�1'�-<���m��TujPX"O�y�u��1�B(��ɮ��"�"O� :P���ŻH��5b���Am�M�v"O��1�a�,H�~��� �&�0�f"OXh�r-� �tZr)�&3J6d:�"O��+D ]4V������%fp�q�"OI�'�i����㫚���AQ"O����Q�Q�h���_�$ĀA�$"O���g�2��U�`�_5���"Oh��wBU�2���j�hܰ�b���"O� �OM�}؊�����C��H5"O�mz0N�6i�h��f���q;���g"Oz�ɰ!Mo��Q*Մښ�.x��"O��3�Z�*V�0�c��6��"O�ԉ��ݱ5Ÿ#A?�@ &"O�D�' �#X��ǧ͏T��i�A"OB��%=mP�G�b���T"OR�5��[;��шV,$D�RE"O
��u�|{zD��᏿fB\�@�"OX�9f��?VҮ-����53 �ZG"O$�+Dʘ�i�0y��>E+^�� "Of�3�����FE�-�d#&�!�"O ��f��x#.�3SmP2|0]y��'�ўT�4O��I��1C�͐o�Y�0B!D��p��1c5>�02Mʵ��o1D�y�-L�_cHt�Ձ�:�ġ��!D�|���;d��Fo��A��A$D�T�%'ȗeݠ\!%-�3qS��X�6D�h�g�o��+k;��r�5D��Q �ܒH�0��N�GDV�҇d'D����ʨb�j��^/$:m1��0D�dJ�C�?��QFɚ�>VX���,D��a�)C #ع��1�L�3d�,D��8gP� i3Ϙ8
�p��H/D����+:�\9r�܁y:����"�IX�'%�	
;�r���F�-�Tӂd
QXB�%X��F�,{&L�T��DB�ɮ3�X��2�X2*,ܸ0�/]J�C��#	�p"���a�y��	y�~B��)7y���B �#^B���"���C�ɿ��6�D����!C�+0�2=�ȓV:��k��>Ub�NZ�*疄��/$,��[�Oֶ!J[�����3D�\�dJ>�rd4�=Y@�d� j1D�pK ��3�d�q��R/~�|��7�.D��� W�$ZdA��7�y��.D�x��ɋ�
8V�땁�3��(��/D�L�d�	?'���aƁ�CP�ܹ�%sӨCተ i ��șu0P*]�s� C�	-$��h�#�ҿmd�����8��B��,-C�dH�Յ:!���J��Re�B�I:��P��;�����"�C�I�g���)��=	T�E�c�E6x�~C�I����b�:�0����LC��?`2d'���`�(ӪQ�C�C��w�'�\tS#��\n�C�	#*2���@ �@ڐɣ�䕞u!�C�5s��4�P�@@Py��g��C�+!8]c��,�$�`օ�b�C�I,Sr!+�!�+s	aH�jz�C�I���z���?}��()u�:��C�	�H���0���':�@j3#.��B��)7+VԢp�P�fo���M�*�`�k���"}��"�1%�pP�&ݣ�,��E�C�<�6�Ę5O��"@GM�;$t�a�y�<qP+�`E�L�T�
�g��1q�(x�<� L R���:"JG�Ŷ"~��"Ox�`Q@��6z�CnA��<Lۧ"O~ī$�D7s{�:#b�8��5#�d6LO�ɢ�@�a>��A�ǂ�U�7"O2���̀�0�0�rE��Cxt"O>��`˧na@�)A�mURmk�"O�P"6eѹ?�*\sb�OT����"O�xKo[������0\p�uZ��E{���K� �1H��n}�$ӂf F3!�DH�]�|pG'E�_�BOHo$!�$U�s���Qׁľo�V��1��?!��@hЩTpq ��@�X�I@�'I�!۶�_�a�D]S�ʭX�<�;���+Oֈ��!�&O�؁x�*Z�W��8�"O$�b$b�5=� D)H�4j�m�"O8XCIݥ�B|�	�#H�,p'"O<�p*@%G�� 
фwAа�"O�ɨ�1
�k�)�<Q=j�� �WX��"6�Ŗ5���@Ə_ubh���4D�,8Β,L��T�10&(����&D�px�/���N��
�f-"D�؈2��>Ds�mp�nO0���C� D����=�jU��c�����)D�����v����Qņ�(�x� �&D� x�JU�r��`���T8)��-%D� ��Ё��y�ս�L٨�?D�,���G�{G4�,��U eC�?D��:�i,��j���8Z"9Q��=D��ٱ�p��)�Ud��+��P���:D�$I���`O����ӖUu��ō4�O��^;���ţʻ[0�w��	.���3��t凿&-���[�cW���ȓ�ĥ�d�]�,y���H�s��`��L�< ��@45��3�cY�F��̈́�,����MNJ�ܽK���+��H��z*�h��Y�t���Xrr��* D����^� Lk�.VRhs��)D����HC�h�� � ��#c'D�D���𽳡gL�@��M��%D�X!so	O#��D�ɟ~�܍���$D���@ '<p��ꙗ��E�G=D�Lk�nJ�oH�Pz�d�9vc �.D��i�+[{u�5���R��2��O0D�hp$h�a�R@
⩏ �Tl�"G-D��R����X�Zu�KB�z@d@�l0D�8*BGT
_{�|ۆ�
�8".�I�#.D����ژo��1�Ӧ[^}�V
.D��Z'�$T�n���� <�����?D�`�3�$5�F�Y�mM$��)Ql"D��Cco��=�d���IJ,J�� !D��"��(J
u���	��p聁 D�@S,�3N�.��raA4Ji��!�?D��bȈ�_D��j]
Q����=D�jd�Y�>7����cI�V%ΰ�go=D�8 ��z�T��K�횈��O6D�@�u�[��@ˎ0h`h�J�h)D����a��t��'�F.�fc)D����%�6���0��9����m(D�,�Y�G'����,�#{<�Y�c�$D�4�$� 1|MZS˝�Vx���(D���A�
�o��䍚�s_v2�'9D��k#��^��)�`��/��!0��6D���q�]m�X�l�Wל�zT�5D�p�7�� Y�ā�'�Z~0b����2D�� l�ӧj^�kߠ�",��X�R�"O�,�kӏ' z���D�W粩�"O����۹��%���
����y��ۧk��	�W�u�x}s�lô�yb��79I�z��em�e"%���yr��-��eG�s��$c�%A�y2��8�������s��!F�ή�y�+�:>t�U�ׂ��n*��[%���y�֧$�$P)2�H�]h9ya�Ð�y�lɉ;��h�e�Ȁe{j�� n���yrlRq3~ q��rdL�G�Ķ�y����1lP�B&�'gW|ua'�8�y�B��B x���5c��p "��y����y2B���H�b!�!�7��/�y�gΩq�^5B�NA�U̥�u(C��yb��!���co}�&W���	�'��S��J��v��+>�|�'p,d�+��GON�F�#D�L�{�'@��'m�G�܉��#*���+�'�Ra�#�/hIx8�5�ڮ�z%8�'�&К���%� ���`O)�� �'0T��/��T�b5��T|Z�01�'����׮* �wFܫ�� �'�^0�TD�u]ZW*H�#�x�b�'P�Trf ��  [�)���21`�'���҅o�CF��v�ߵ]T�q�'Sr�0�G�M�<}#�g����'BrȖo��f��Q[c�>%���
�'��4�jѼ't��B�!kH�8
�'��8��-��S���AjF
M�
�'�*�2J�$�d)��60y��'�d�"�D���ã[54U ��'����#ˋ6 -�L#V� ���'XXl1��Dr��1���JW�A*
�'y��+�e:��ȓS���@��]A�'&�mc��ɸ8|�H�'�(!�A��'VhM�U�ݽ[|Z�K$C��%8��'�t|��h<��C�GT	f�����'��e��/vr\e��O�sm����'b��ض"��TZ���NDl�LU��'rh��B! <N���#Yfv$4�'�~}��1x��Q������'��R�/	�9H���ɗ�	cF|s�'������B�ҭ�S��pj`=�
�'��E��Rժ���+ޚ`dF�
�'s���ʼ Ҁ�R �]7�L#	�'�rh�&LQ��q9�.D0|�$��'�V��vL�3rF���NE�}�����'�60r���c���q�-K�~�lD��'ј|����+��d�Df�>x�#�'�p��aU�/�Yt�4~�l��'��[f�>f���y1�8�'�>����2���S���!��<��'�Hh�Ò&`-hvj&m3���
�'e�Q���s����uE
�0�N���'Xxi��r
2�B"�+R��A��'B��h���*\��e;�I��a�� r�'����� �- EHK�Y�����'I�k$%z��s�)V\����')� ��Loa��I�E��';�U���R�4+�7O�DT�'uD {v��l�n(��gQ6R%&��'v̌bb��~	�V'�;:�X�
�'{ ��`��A0H�dk�#g���
��� �ܠ@�T&@u�|1'�*���se"Oz�F녽+ʼ!`���t�� A�"O��j"��'�r�-Y�_�Ҕ"OJtqA!P= �a���5Ĵ	��"OԴ�g�
6gbи�e�|��"O5��Nx1a��_����"O� �6Ϝ$*��Ă�%J�D�ܭ�"O�$�R�Õ%z\�6dM���"�"O���sA��~'zp"��@2�Фї"O�
��+�jqK�n���kU"O����J*[F�d1-��2���х"O=z$IϕM42�a�?]���i@"O���V�đl���i�J6%|���"O��б��	^��#��3�YҢ"O���cO��r4����=�|�hB"Ol��pW8|�ɲeٙ,�l�E"O��R5�~bJ��Ŭ�P"O"q˷X�A;�tkӤկa�Ez "O|)ZT΃/+O����.hh��"OJp	���0|�
�C�2+�b�"O�|���r28��'��K�fQ �"ORE�#@��TD3���B�L#v"O<h��#�0�|�#b'a�~���"O��ه�M�
`�I� �!\���8"O��@�Kz;�� g�F`N�%��"O
1b׆]6~ ���AANZ�K�"O
�12�n�Z$o�wKR���"OT�8�@��a&ڄ�W(͘.c���e"O6X��lŢ}��D-�	/cP�B"OdQ�3�Y�b3�)��L[�RE�p`$"O��a��j��ȣ����"L���"O<P�#�]
Z��503��XE`��U"O
��fJw<i�
�+^D@@g"O��p��@�`�,�biҹ3KZ)[�"O�5�j��X��x�QH�1@>̭z�"O��S"�$Ma ��w&�*�Ƞ`"O@}[��]W��CT���T�֩Rp"O�����! �!='�θ�"O� B4Ͷb�>p�UFχ�P��0"O�|*bA��.�n�#��\���G"OB( 6l@��sG	/
ڀ{�"O̥B���6b�,`�fcUI#"OJ)`�+�/20��7�Ճz��"Oe(Y4В��Yޡ)�"Ov=�n�0B6�T�baD";���"O���C��7���+��� �P�<1ь�(T�B h7b[>�*��7��g�<�#O= ��%��a��<��@o�<	3&GZt�}A�ޥW���j�F�<�1��H���C,W^�(��|�<�G�\��({a�O�O[ZY��o�<��mp���q��%��M�b	@P�<��MRY�R!� ֤9jƬ�s�<�ʛ�Z�QAΌ16�PR���q�<aD07,0	�j�	�Ni�gn�x�<Q6��4}O��@f��<gk4�pૉ\�<�7M:g�\@푳c�r\�'�U�<A����_F4
�C�+!���!�(VX�<����VO�JЊ��؀�X��p�<)3�1�"�bCJ-[���0��C�<�g �XjPy(צ��X��T���	y�<����D���BhӷJ0f]��g�u�<q�,!��� CC՞aD����Qq�<�ub�t`hy*P�49�1�J�c�<� =���1{H(3�oG����j�"O���IX�;&�M��D+���Q�"O�h��� C�5	�-®E��y��"O �2�г/������$Nx.��"O$�P�Y�[޸`���:m\�\��"O�,+Hm�H��s�F1.L�8v"O�mk�9�9 �Ӽp,tA��"OR,@f����-���	2e��)�"O��x�Cv�Ԭ��@����"O�	Ir��]\za��/�_�[�"O���ٯa���n
4p���"O���D���VZ4p��j7�T��"O�AP��1>��	�=]�La�"Oj��� TW�!P+�(��x�<�2�Nq�ƕ�f牴M�W���!�ć� T�M����R�Z��G#�d�!��R;e�2�*A(J/ֶ�7BD�g�!�MNad5��-F��,��a"��t�!�dT���DDƼG���1�aG=>3!�D
�zn.�0 KѣH>�-�  A'!�$�$$�.�
��'@� �"����!�$?2f���C$O�ݫ����!���j���Ι�oHD�҇a�$I�!��&	��)S��<9�b��[:*!�d�:XF()� mЏ|��P	��L�!��A� &�,0����}�8I �O�<�!���(��5B���9�$�Uk�&H�!�D�+."l���@<\��J�`�Q!�d��0S~�y��ijȉ����%@!���"u�^�Z$�U�^]��&�'Q<!�D��T�D [ҏ�5j��� m-8*!�'i��-��j�)n4��rI�F!�䔤��vf؉LÌ�X5�9G�!�$f�
@�D0}��J�#Q�J�!����y��c�c�J9�T�ߵ"2!�$�3^���#�!�5c��Ұ C>K"!��H$1�Y�fU��C"5!�$Uw��)K׆��NZd�$�	�!�d5-�j=)��ۊN�Tp�dS)r�!��MY�~���R8t ;wi_0v�!���?n��K�a_�g7�]zf�Ӆ^-!��
?d�9b����� 1�,!�DV�onz��Q�r�΅J�jւB!�Zcx���	�,)��5KB�C�r�!��orn�;'��8������6r�!�����"r@�-r9�A�c�!�$�	#�<���� �
ĉU F�!�d��r(�!�!T:|_�����!�Đ�W�plK�,S(a �Ce���!�D�m�DX;d��-Hx��7�
�'�!���Ը-�H[+�r);S�Y&�!򤀎2�āpS"�$%(�C��"�!�	$R)���RDC	9"�P�*/?�!�� m�>,˄�[�q6<;���;S!��_���(z�e�!s�q��Ϋ5M!�d�%��(���= �9�$��/!�D�=Z؀�"&Q=\�,�a�? !�D��E���T�T���Ł�G
{�!�D �p��� �\�|YKT��!���
%�"X���ݟE�����"OL��'� @b4�7& 'l�U��"O�<��0��E�7׉	��0�"O����Oưsxy7��4;D��r�"O��	���Z��C#�jHmx�"O� <H��KwN����,Sv���"O���`	]�k���K4#ǡc<4*�"O<M�@�\B]A�W:D��5"OP���Z(�X���,Z�W"O�H9��R�1��%`�b���r"O�Ss�[6@�f�-d�е�"Ot\���Pv�U��+Fb�[�"OpѨBIΨ"��u��L9��8"O�l�2lR�o������;@-���"O�郢�N�~��%���wH��b�"O�@��i��V\0��Q�	2��rd"O�꒍բ@@�q#�^E=��R�"O�m{3�YW�0���*'��s�"O�|+�䎔IV�t��i�!3`��4"O`��F�Y
�$l��E
L]�"Orl`�G\;b��|��b��r W"Of��E� P���*��x���"O6��E��^L��ɋ6>�Ω��"O��7"�4GU`� н=}\|�"O�Ȳ�?ԥ;�f����Đ�"O��Kf�0q3��p��҄[�Z�2�"O\q���B#Y�Y�0

�q(��e"O*����yp.U�
� 6�t��"O�i��쎌rT�P1�*�'f���"O !GdA�:&(�)J OS���!"O�� 艀iPH���iJ6GI� b4"O����j ��*͋�� 9FJ���"ORm@m�`68h���#-.��"O`y���4�����C��%���@"O@��MJMrY�B �2y�����"O�-K�˖k�����HO�I:�"OF���Oܚ/�$���	�~7����"O�ԥH�)�P�&#�$M�H�:P"O
��HX�Z.(�(Y|p*��"O:P2t�-i|�"$��7O��t:v"O���(�A4(Q��Ԋ.��@��"O��3��È����gܱq�Cv"O��s�K�BtҠ���)bЍ2B"O\����DdHU�&�5l@,0�"O����ɷ_(fT;�.Ă-<)K�"O� !`H�~��{��,*�IXS"O�ys�e�#�:q`7�Q�\ ��h3"Ox�A��B--�����5"O����h��%brL���֮-.\H""Ov�ӷ�'O%,�:�B� )�Q(R"OD�Pȅ/���0�Yvd1�"O\�`˭y��3r�ϰCUH�rs"On(k��ˢ]L
�m�ii�P�"O���o�:�k��TBV"O<��"揨/�2P[7d�?W��t��"O���[1/pb9�l�@4C�"OLp��� Ā�r+Z7� $��"O�I+������P�
C�b{�DA�"O���'!Q6:�Ȏ5d_���"O��:��B�{��4��'G�	$���"O�ԚT홄\����牡v>���"O��Q� d(����[Z�"O*p�#A�d�p)��S2zԭ��"O���Ў�5uF�\q���?X�����"Ofr��ם0��� ��L�.��"ObQ��ݷo܎��`/��v�Yp`"O0�a�`	�2y�sÅ'\9��r"O�<�b��"�8����_�Y#t��"O �H��P�X����#ņz&�J�"O� �u�F���C�z��#ܳ;
���c"Oh�Z�n׳y�f(`�!=bO��R�"Ob� ��I$I�6� Q�ülH�ع "O^���kNN�8)1 �1/e�"O���@ß��j� �oI�Ec�Ay"O0�E�hPt��w/�
K��1Q"O�7�ϳz�<hK�D�f����"OB���G%)6��5N���113"O��ab��|���g+�##�d�"O�@�4*.=1�1�i�)���q"Oً�3Ʌ��#���i�i�	!��ӫ�x��sfE(�ƙ��⇃�!��\�:H���[n���f@��!�d����Y��
b*��uG��v��Ik����rk�2ws��*Q��;|$h�@�%D�|aR���k�&�C�֛-:��I3�7D�PҶ��8a����g�+ %�P�!#4D����"�C]�x8G��9�jP�k6D�d:��
*A8�+@��.�2T �(D���g���&��@r�H���a%D��S�V+"xpȑOư}'��`�7D�8�gO�#d�R}���B�'����B�8D��ڂ���B�zy�W�_+�b9�v�5D�$˓�E6Gd��</��l���4D�p1�E��!n��ς����I@�1D��A��G=z~�	'��J9p!�0D�����@��R/�8Q:"g$D��q�K*�L��p��y�T�j%�#D�ģ�J\=��h�Ɓ)s,$��T� D�t`�A_1i�k���/x��t���(D�����0 �n}�������3D�Љ��4$�4�i��ʧ�2�8r�>D�`��*�$�k-e��̂�;D�4��l�g->}���N�΀���=D��@eiە8d�gM6}��u#�;D�ht�I�AXE
0�ݒZ�Q�!.D�xt���ZD%���ٶbkD�	�@9D���5�M)bT5aU�W %4�rV8D�s�	��t�!OA�A^�R�6D���3��K4H۴iZ<p}0� 75D� 0�hR�.Nbi��A�jI*"��1D��r��� F��r����$Tc��4D���%�:Q8�@�M�eRbҶ 7D�<0�C�>9��P�b)ń!���+�D!D��$ſYkҴ����+U\$��?D��X���9�Kgk��Z%*p�@d!D��rj-B�A��L�H�$-D�PS�أv5`���J[-n�����`)D�L�Ȅ,,Jjx�B���%��E�#)D�p�'��$%�����C�;GZ�qR�k1D�Ԉgj�7���:�� �d�B��4D�|0���&W��a�g��o=8��3D�H�҄�+u*V=�#�K iAZyI��2D�1��݁�D�
 ��/# ��`@>D��#����j��'e��-� �Ċ.D�h��U8b]�Ţ��N<,�Ƞ`#�+D�����N�@����b�K�B�91�'(D�Pz򨅿#����
a;֝��%D�`��	���ۅ"<{ X�+�-"D�H�G�����v�[�;r��7���yB"�qa��*���)7ז4����y��]2��	����~-0���@��y��&蕋�։q���c�'G��y򎟨;�,�a�Ffb`�Q GG��y
� ���$�K���*+hX�5:"O�|�!��
7*��B
�[�.d��"O�ᇏ4f".99��M�(Ѡ�"OT�0��{;ai�A_�(3�u�`"O�M�T�R5-�b�2 H&|��b"O�"t�l$�c�/��lb���"O��DE�0�$�"RbX1 "O\���Ґ_�����0��B�"Ox�a1�&�"���$��B�����"OpM k�6 ����B�{|X�"Oʡ��N��Lq���O�	`h���"Oac@�	���Zb��Ik���P"O�q�Gɯ=X��p�B=uh$jr"O�ݐ5�Ѻ�byzW��u^��P"Or��&�'/�Ơ0�35xrY��"O�����׫q4��5DÝ
�8��"O�m1%���K�I�P���:�H��"O:��A�n��0�$C?<����a"O��#�I�M~r���a�=�й��"O�D��j�3��a��ȉC#l��!"ON	f��
�����H6�J�"O�8�,�4� �'�-��R�"O��J®ŷo�>A1"Ɨ2;]l1@@"O`�!�+��=3�e�gHFm#�"O��`v$��^<�B���j:�#G"O�����dO ����P�v��u"O�Y3fC�]�V�۱'S�@p��"O�@!���AΑ��A7x�DB5"O��#uCGB��\p���*f$M�"On���)��Ls�ʂ�sd�9D"OZ}j  �I����b��`�'լ���蒂@z��8��01�I*�'�\�s��N+7��k.B\�M
�'�25 u��OƄ�ɏz�I�'{�djv���]�qi2x��p�'^&����:̃��W�e��H�'����d����� �H�]�N2�'���3%$ q� ����W}x<a	�'T�!����桂&%BR�`t��'&�So	$-:���a|*q�'��k��LΊ#���GL�@�'�l��r�Y�c6~��Ȟj��0��7��c���&d�K�0��}��WC,�	�ϖH�ji�"�Яno�͆�������
�l� ͭ:na��w���3�B�7h��y�WH)k�d���5���1Qc���Ha���|���ȓ*',	{`b��
"�	���S�j����ȓVP,�`�bV=��.��oD��ȓ 
�AZ�y�~ ɂQ�VG��� ��hjq)�]N$x�G�%6:U��TG)KT'+u�*�#���#����A0����q�F8(���F�v���Fd(,1���G���!�6Q �ȓ;gLP*��_�?��(�DckY>X�ȓ2ᶙ�4 )��9��� ;z!��~d��b��S���В%C��!򄌵n�-�U��<����&���!��6k���8����!��"�!�d_�� \�U.��V��$��ڎq|!�d5o�$SQeN< �Z=8A�@?l�!��	��C��l�(���@ܣO�!�d�UC4u��)L�|#����!�X4dQu�3�����0FG�s�!�� ��h��fgN(#�g�\���H�"O�����z�. ʲ'�!4��Z"O�Kr�@�o���&g��Y����"O���2��4I �[DŚ�kT�ñ"O��P�ń�Q�ADQ*uUI�"O�����z1n�Q)�x���z�"O���	R�!چE90�G/[���1�"O"��'n2)�|m�@�S��)Z�"O��s��^�h|sc)X�mBF"O�ءt��,��C�M�$c��J"O��zG��e��c��+O<��"O��#��������
� 6V��U"Of�S��M	,Ɇڲe�5#�؛F"O��:��I�ƾ!�'�V�s�~(Cc"O�3Ѣ�*8��U�u*IC6��"O�������-�D L0�½�"O�eR���if��@ʂ䀧"O����E�-'�Urf/��p"]'"OZ�s�c(@�.D�u�� 
�.]��"OX5�f'%`d���=h�h�K�'6�mP�gv�=���X�m��1�	�'۪eQ<['��+ƦJ�9���	�'���X�J�Ԋ��ω;;���X�&7D���DI�4��v���\�PH��E'D��'��?4�@��BLҡ<z��%D��a'*�a@R�@�sbT���,#D�Իv��D`��d�O~LH�cj D��P��]d�� � 9"ޕI�K#D��8'��
_lyx���%J&�Q���#D����恰e.��� ��$�~��2a%D�0�@B�ךѦ,T>j<J����>D� �g��fc(�ļw�Sc�:D���럤�6�9D,B7� �*  :D��ua8k�P��&�,���@9D���a�98�����M�F��P�`4D�L��|J H�c��5�|�d0D�P*1�s�y��ɝg3Z��FD1D��åB]?o")k�E�0Vqa�C=D�x)�.��_0��#�![a@d9D�\bC���E=�!�"CĤoEk�3D��ɷ���6TD��B4`И!Q�2D��{PJʜk�"�%@]'ʐy@0D��p���V�6�#C݄7�����A9D�`���\�
��;ǁUD�h�r��6D����m�n ��a�钣ʝ��!�!�4�2:�J��CG�My!��E���t���*C��ae86}!�Ė�w�$�X�-&���v�+j!��P74������4H�\�K�S�!��Zf�	�,Q2& Z�&S	�!��A�| ��iAO�M�OD�v!�d�_3���4�BJ$P�cKB:!�S�)���QaĎ%�^�@Њ]!�:s��r�ғ��� MZ, k!��@�ye�R�,j��q�DW!���
C4�͸�/ZUZ~�"d�ցC�!�$JWA�`�E��H�)��2�!��J�t����bC@&<�$��/��W!�$�6Nd�젣i�d�5�e�\�}!��9M68p�U&�cD�*�l��5�!���
a2����-c,k6L�+s!�$ƩDJ*�Ѕ�RW1h�R6��%g!�D��uk� 1D!ʘwHt��A�&pD!�!=�H�pNޙs���:�/�>;!�� �(��~G��2w/�j@ʘ��"O�2��֖_�Z��1�{�:"O�a0�g��T�4����D�O�0�*v"O,���*�!� B/x�`i��"Op�w��%&��ږo��6"�m�"OܰY"�R�4�X�Ư�oP�c�"O��IW.!*N��Fo]1hhC�"Op��P�.8)2�͏�� 
"O.�%��2[������Nv&(�"O�X�b�]��Ux��
�q��{W"O���͗��\�#O� t~�(h�"O��+���&�v s툿-͖A;�"O.�ДFT���5��K�Z�AW"O���6�� ����F޷2�JQ��"Om��o���8�[����v�"O�,B��;ĐWƑ!��<(D"O�J���i�d�Z+5���"O�p�,�a�F� ���/_�tt��"O2@s���Hz��/<���"O�9��)R��2í�&x��j�"OzK���n5�	1�B�X|�<��"Od��É�1KA�A)�B�	lZ~uZR"Oh��G�<��Q�4+�#BY� "O�y酧�+kR
�*#��'��7"O�$���`�hqS4'B]���k�"O�A�EEđ"z\�j�
����!�"Oq������l�M^�����"O>9��z"\���S��\�"O��y�bB2����]wr<d�@"O�y�6��6c"��F띄s��S�"O&�x�얌Q�~A�5K�
�J�0b"O@<�S/�&9��)I[ v�P1�q"O�r�I�l���kP���x62��"O���E�[�1.I:�Y�>^��q"O��S��  �ƨ1B ۊm����"O����"A���7o�<�>H��"O����T;v�P�i�NB:�9B�"O���$NTQ�+��A���A"O���Qǃ�f񞰠D��B���C3"OH�C%LK:;�6�{F �<O�6)�"OP+�A�@?���N�/�����"OA9�e�4���`���c|X�!"O"t�h��g{��iS�
�J�$��"OF<ZDY���zC��,0���"Ol���)_)f>4�u�΅$4Q#�"O�IT)�X�"�A�0!p��"Oĥ��i�=f��Ő���+
D�"�"O�!L��k�r��&��Hn4D�D�!
I̖\У��������/D�d!%i_1�-K���J��@�5�2D���TO�K+"��
;��`�t�;D� ��͎+f �G+`J�l+�+D���B'Sn8Qc'���Z�4�H�L?D�,YS)�:ĵk�5s��Ҷ�!D���"�<	C�"H+@����>D��6�:/��i���MqLd��M"D���4+S���B3`J4I`-,D�pHfcK^H�3R���s���p�$D��Jbi�]����6	������$D�hjs�ơ#)X���-�":t���I#D�@+g _�	��h�0!Z�^AB�H�l#D��8�
�C��T!��ؽP�.���+D���7f�2.	0lx ��r3��5 (D�8�𡎒_n
H�͖d$ĵB�`"D�� ��g@��(`b�G�2�
�p"Odsͽ8��$1��I�Xe�h�"O���BL�0�N�8$�F�-W��"�"O�C��M<� vn]�E�0�"O�y��KӀ�uCrH�Y��$�"O�h�f͛����V��l�"O^�1w��/^�Z,�]1)[�j7"OlA�@ɇD��a3�m�4M��G"Or�(����g�,�(�l�=p�ذ"O�m�я]4����F@�M$�Z�"O�������q%���?�~P��"O(YqT:f`��`�EB����C�"O� �f� ;(�hģ��s~n�Hv"Or�k���x7t��Ҿ;{�})5"O.-�"IӃ@vB1����i`�ݰ�"O:����J	�dt����QH�9�S"O���v�˘lQR��G��1�f���"O��!�S<k�6$���&��`��'D�ݙ��G�v��� %��'�69c%hJ:?/6�S�/�瘝!�'���gF[�W�#U��-aѮa��'7�dKpjQ<}a�,����g����'��Yc�*�pw��0���1_�UK
�'�j0�n$;��,{S�̉&��'AFp���l̠�KT�2���y
�'BU
'�G%
�x{Ð2��i��'��AT�b2*Y[3��8,De��'{��f�ԁeX���&�P}:�'Ҧ!��h_�4�Bm�Չ�>�=��'�-�D�F����7C �6�'�]���XzRi*�bJ�y�n8��'�@�Q�Q/lp��fb�i��0��'�>�Q��e�t��F��9f �
�'P4L��̋L�(�:�Λs�2�'���Q!�5XCz .�x�6pa�'� 	@�0&K�5��[�gA�T�'�N�8�)J�~Tz�r�#7Y��0�'�&��C�+|�Bs��ɩX�Q�
�'�<R���	IhqUJ�&��qA�'c$�r��(z����(
����'R6z ,�=HM�Fߕ��2
�'�
1����lI�b�>2c�'>2��3�2@�䐔��5w�E��'n�)��O�#��S���%u��`2�'GB�J�k^,s��`����V�N���'HAz�'ݠ.2p0+p)�5�#�'V��0ŋ]�[���A'����'�pЩ�Β�^	(li�e�e�
�'���R��"R�Y/!��5Е+�i�<I��Z�	:�ۆ���=¬tJ��b�<1r�9n������נ!�C�t�<v��)�\�i��D+��I"��i�<I5( *�`��3T'||z���c�<�Ҏ��}��"$��!a��8�w�C�<Y�_axz=��BE�3����@�<��,�:2��C���n���5�^�<��#��k."x*�$�%Y�a��e�~�<��$Ͽ_�̉9���#Z(��`VkR{�<Y �0HX�dA�e�^�� �N�<����z��۳Iāqp�JO�b�<��Dx��pp�=�`�"��\�<��-�,	9�g�8{�=j&'r�<Y#B�Z����`�[ʘpF�F�<���I>5��m���6$!��Y��A�<� ��
 $_\K���􌎥�*(�"O(�G�J݀M��K�6q8\R"O���τ��BH���1w��h�"Ox�BUJ�3���{v�Mk�Tp��"O��@�I�?�t�҃E�]�����"O��!%6p��5������"O�8��iX�?�<�����A�&"O~� �Jkr�@�t�(H�EA�"O@,"tI@7"1d��Tڰy��aA"O�i�+��E 
$:��/�6Qb�"OL�2t(W�S���0΁�4�P�c"O
!j�&�� �>\h@G"R@��P"OЁ� [?@��A�B;ν�"O�5rs/��qt�2-��,�J�[�"O�(��+�(Q���C�Mي,h�"O����bo8��ׂ?_�.X�"O֙k7�F7`��@�N�>���k�"O��dL�u=6��uk�~���6"Ox%�7c]�F�*�V�B�McLI!"O�=B@C��A�F�5>P�P�FGF�<����$�V�Ce�Ϙg94-�Q*N�<9W�I��
��G@�[�&���GJ�<q�L\�h�Ԕ@���Fr虫᥎H�<��8N�M��ĳ=����O\�<�I���@�t�$1�\!�0�Rb�<��䃦cdI �$ءi�F4��_h�<a�-�����*���� 
M^�<�A��3��5���E�)G����L[�<yVc�6E��A1+A7XWƈHE��W�<A�B9+8��F^�QGX`�M]�<��Ö�$��!���/��ajE�V�<)�Ȇ�@����\-i��H�S�[x�<!�T*��(�E�%,u�
Ҋ\p�<�GL�f
�|��-�V(r���v�<!�G�J�N4�#��FQ�I!5�O[�<�E��
=�\u��pCjA��ŏZ�<!� S^��\�ay�� 4c�R�<Yc�mY��2�Kɀ{O�����EF�<a3�W�HL01K��?a01�u �C�<y ݜ �t�G�Lۖh���|�<I��Eb�L�E@;l�6����B�<����}�zH�G��b$P�dlU@�< ���Y��"#������z�<��yԬ��A'ܴѪ01���u�<�s'.Tl���H�c��5 f-f�<q�dS��0�ZW%R�"�\�c��l�<�7.I
2�@��e;�$�Ӱ��B�<a��7(&��3���49�!��A�<�O��nD�9F{��e�'�b�<�t�Ƞ+��;�n�6-�}�R\�<9%��Q�L�6�D�j�y��ImyR�'��Q@ 6tmE�FG��O�ȍs�'&�qL�������G1IҢa �'z����O�=a��[��x@���'>�B��(#��q�B`�?y��} �'���R� C" *��⨆�v�����'���)�-�����32��C�P��'k�����<_�0�a�G���'��Q �E �|��ACXi�p	�'CN��$�I+�(hv �cgެ@	�'=���L��e3�d@	�0@�'j���B6��]�$n�%U&�)�'�<C׏8V�<�c���K���'��թ�윗��k�$Z�=����� �sp�U  4fKR�"Fvh�S"OT��k�=A9�A�WFkv"O8� /J�(�B�	t(V��d0Ã"O~�ɥ���d.��q�q�Ҥ2C"O\�Z0�����Gl�u�E�D"O�� ���C�xT��J�t�V���"O�=��@��q}�<)EgT(�FYQ"O�z�/C&\�H�&	D���@"OXDRd�Y��~���E^:��X�`"OZ=R�Jу�0�����$Qr�,�G"O� ��LA�A0�8�K�>p�l�+ "O"��I�&��5�*�!����"O^�k��(Z�p��Do<�2Y�e"OD��aC�/:O�i3LX�/y杻�"On)FJ�<{��UAw�ߣ@i���"O�d�A�G %HmT��>Pz��w"O&�h �AD��S%�(;l��"O����I�U+H��1D������r"O���)�O�HX�BÚ�C{��F"O�� Lڼm����A� 0�h��"Op+�$G� ���X�@�n̊�`#"O��1U��r=���)�A總�G"Od���o�"x�a�dG�$H����q"O�Ce�OL��	`��-����"O�(1�J�2��D�'d)�|8�"O�!��?C���B@B|
��A�"O��R�Z������a�"O]3��f�&Lf�L=�G"O!��5
!;�X*-���"O���L�9zpe�"�{0
�T"On<���٣}qL�AN/g����"O�+�i�8!�B�F�Y�8-ۥ"O�Q�
T/B� ���
��I�"O|1�񥙠H�Pyj��P���p"OΕ��рV��=�c�] tQ�"O>`c�I�;=�m��m׍a,F�"O���1�wnz�G�ޓsm.ȓ"O�ɪC�&#����/�'�ĥX%"O̕�R��&O��r.��DK��yȐK���hׯ7go�t�a7�y2~���E�8r��k�vI�	�'�ĩ�WN�N�^�;�F�k'��'�B�X#:��ʵ	�d� p��'�fP�ŭ��
�ֱr�(V����'���1%狱O$�a��!C�4�q�'~����Ó72�tL	"
�Q�n͛�'j�"D��+�
��т֏A��	�'R}ҡ��TXZ�C��9�6%�'/b��PL�#fu��s�Ɯ�,P|-
�'8|��E�����A`%���R�'��IЇ��y��ܢ�� �*�K�' ��p����z=xC� �4�	�':h���ŵy)�a��f��	�����'�=����*t�������z�2�8�'D��GgI-_w`��E[�t%���
�'7�̃�B�8Q�dY���f4���'����1�}�0��C靃�v<��'����hK��(�zs�y�'��}#f��&F������ir�a�'`���ĳ_p�钫��7���;�'���xw@��d�ИB�7�����'�h���W�,�@s�e��"H��!�'i�E�⏖�H8Rrh��-��P"�'���[��pˎ�J���1V��
��� �=`W
A'�ι��P����u"O� {�KF3/�1y�)O�p�)�"O��H��*zx��4i�z���*�"O*����~���ZR�D���"OZW�u�H�@a��~�a�g"O����� 1$=��c�p���"O>��؉j¾T[�E: �A;�"O�ɂg���.rࡣ�H����"O2�&.K�O�P�� $S�x)"Ol<P4��	3��!�R�2.pP�r"O�Tj�n"\�qϱZx)f"OH������XX��UɁ"Oꉓ�/��R���� �yմ��"O$=�c�C8_�*���<�ܔk""O���`";?ȌYr%cK�l���"O�q��T�*W���Ө��6��`�"O�H"f2R%��"D��#]��l
�"O�iE(R9?�]�R&͸)�2 ��"O:�a`/����N�+r"O
a۰Kх=��%�S��Y6�h��"O&9!3_�cX(I4�R�L�Aw"O4q����
G�6Hf@����"O�U�1̖�N�(�����	��"O�Gl܈4!�0�q����"OvUc%�!Ww.D�gY{�H�"O�� 6���j��Ի��6b���"O�U�si[�|�鉥BO'zBf�0"OD`���m��`���2N2�I�r"O�!j�h.���&���nQ�"Or�xwGA�n�b�[��B�)���"O�yx0���y�d��9F��Pk�"O8��po�=ب�'jE�y�`P0�"O��ⶄG0-N|A)F�	��q"OX	B�����L{���c��hkU"Or�B�@v�Y�&Zf� a�"O8u(U�ٵC�%�$	�Z���(�"OZĺҌZ?P�09j�P�ps�PQ�"O�a�T�V-��!{`՗$�M0�"Oq�E�Q���8����"O��`�ї����甗h�X�s"O��9�g�q=vA�(R�tZ��)�"O�UȁbX$ t�WIv!S"O����.��
b�^=J�"O�ػuȀ�'k��1`!	?ox���"Of�a�LaƉ��/��t�U"OB�a�aE,-F1�ēw���""O��i�l��:"n��Ҏ�/��$"OL����
$����hD��"OнC5%Ea>ѓ���j~���"O���5�M(Jg�P���H'`b�"Oe*���%��\���U/vN��PD"OlpA�g݋f�l����-0�>8��"O���i]�N6�5'&�A� ��"O0h�Vi��@�BA��:rp-��"O��b��vI8LSj�PP��"O�僅&��0��?� !�"O��4$�Ub�H����`�����"Oe�e�>+^və�HѠ�8�"O`��� �����G�=�Z�IT"O l�aa�v#�J��0:��=z"OZ�u,W)Ϝ�IRk�+Dpx��"ODZ���T�ڌr���U]b�""O��kB�zZ=P`��/_�}#'"OĪ�n�Y3M1I�-5@b�P`"O� ��95�D1H$f͂��͛*�"�%"O��c�Ǟ�9
���3 �5_�v ��"OD�
�'8�t� �0!�"O���o_��(y���#j��"O��r��79�E�đ�A���"OV�k�-Op#��1��c7"O^tzC�ڽMF1ce�;A�Y1"O�5���7m%�YI�cԯD����C"O�4���)
M`)Q"����Ĺr"O���E�6M@}pj��y���ڗ"O��t�>�~��IR�b���	"O���/L .�܍!�� ]GL%%"OΝ��נZ��k�DS5n�s&"O�	���#C $��cд��:�"OD	����Һ��"Fx�	!�"O��r��Y�&�C�h�Fh�9ɱ"O���.�0z�~iKa��7ij��"O�4�n5|�
���cb��%"OD�O������Z�Sj.92"OD��J�$X�Pヤϧ03����"OU�$mH>���BCΰN$�zG"O���bSЙB���l��D"OT�����6��2@���0Dȥ"O�$��.�:� h�bI�|�R��"O|���m�>q�Y��-C��|��"O:��l�#'�@a:��C7/���PF"O�;W��,�m`�� >�r��W"O�U��!�&�[Cb�*ʰ�c�"OҠy�l�%{&lm�QC�l�� "O8�#���u�0��'Csz8QU"ORa��	1^pT�U�ԑv�L�K"O,��i¢/���3�!�
Dt�@"O��g�A�b��G�^=���qc"Oit�2[�`��L��X�S"O�pd)� 	��� 3FĴ`"O�*dJV�]��� ��\""O�m� d>H=f|pp��i�!�7"Of���-�j�d@��nL'i�∢"O���
!P��I	���<.4�&"O�����K	\�9�B����t"O�)��(M1& ��w-���r�`q"OX��#hA�0��4�+�Z�2��p"O�]!RkKnS����<z����"O��������i
ٓS��4�"O��Iҋ.���0'͈.E>U"B"O�諀I�4\xKc&:&P��"O�IJu�X��b��gd�P���"O�s���qA�����J�����"O�aX��g��ə���8���"O���c܂�v�{���1؎��s"One;�� 2%E �(�M�W�bw"OJ�KƎZ"[��rN��*���q"O��	u�V �TmP��3�6�G"O �Z�nW%m��Dh���@q��"O ,����AK�:աS�$�t"O�%�d�i�,����^�,�<0�e"O��SѠ|O��k ��P���X�"O<0�I?+3
�"�.�6H٩4"O8�����Fv@�e��-Gv�	"Ot�h��A�h䂅acQ?R=�5Q6"OāfB��Y���Tl��HGZ�b4"OE�o�(0)�BlC#CD����"Oȍ�0J�?W���E�&#`�z""O2L!���H �
(k���@S"O� �%�n�8���:<-�9��|��)��a�: �Z+Ln�Q�HĶ]�NC䉮 ��[���0O�*�1iϱ"tB�I8{����Ї[�]]��04�$DlB�I�:�H�6n��&�lA��dO9]@B䉘!����n�Q��!`B���C�I!T�RȐF�̅y����AK��B�I�	~����L�1O�(�Џ	=`k.B��'"����	����''o�4C䉌;��-i6T�Z�����Yo C��O�Sg�U�h@�c��:�B�I ��9��'[�N�LH�����B�ɫ���+%���k�^��U�M3bЖB�I9O��Xx�#ɷ�\��PB�5\��C�	1%A�����'w����wgT�3	�'�DQ��L�(�Th���_;����'�f����J�}�l4��%TĀ|��}R�'�i�����zF�U���x��Ó�hO��*ˇ$8��n�Z8�ʔ*O�s�:bx�d�f��	+˂�����y2N50�&�գ\!1����!G��y2�C3o��4��=*4$��g���y�
πkFY�vd��&V�9�S�Q=�y�c$�6��`�C�pQ $( CNc<�=E��z � ���|-+u�:j0~i���f~BFN�8���'K�$XVZI��2�?���'U�(:���~����Dg$]���$$�� ���,%�Xa#%��b�J�	j�!�DX�6:P�R�S��0ڔ��x�!�d�!r-b��4�K���U6�T'�џE�Dhi~�䪆/˄H� �C%Q�yr��~�EV�:&�Ր#���y"�W?v�z�+�N^������&�y�H�*CY^a bE�:P�ֱ�0�_��yR�2j�0���.��u��b�E�y��ޔuod�+ӆ^��4|bw*�/�yB`�8u����(��u��x��i���yr��+F�r���A˿5��q&G���yR���F�jg��"PI��h��y�MӲ{�$IC�7!3 �J����y��;1[�s,C�%�
��G�Ɂ�HO�"<!�O�+�.�z8�d�U"�Y��� "O�y�q��$���qʙ�I��i�5"Ol��.͈y܀�ecZ�r�&I�r"O��;3*��M=�@��S�r�h ��"O��Y��5>�,3BJ�Y+�S��'����)ҧ�M+��V] B­0Ϯ,z��g�<9,��}(�q�#��,8�`U�"�^^�<�GN�O��QQc%] 0��b�[�<)�K�, �Iu�i�&�#�#�[�'x�y�T�?~�L��DP�[ǌ�P�*ښ��x����w�ș@��K��m�M�'h�!򤘫G� ) ���E�
H�`X� u�x���|�'p�(�ޚx;pPb��]sȕ��3�t��뗒@Z�qC��Ӕ���IH�6GN���ѯU,tӦ�I{�l-�ȓk۸U�)����H�E�lT�bi�<a��7@�n4���C���h��g�<Y%�q�<,��W�1���(�g�<�Bd��d(Dq��J���D�afZ`�<���>}�����k�l��B�O����{Z,Q�Ɋ^y��BȟTf$�ȓ�钀'��e��$�$(�lnЅ�	�<a��`�����*<�:�pvF\�<� \ɑ�Ě;�2�	c�Y F(p�j�"O<	bJ�*���n����!µ"O IB����-�YD͔�@�p��&"O>������#]�X��T��N]S�"OX=�-T�$� Dl��fL�( "O:��B�"��u*T���%fޥ9�"O�(x�����qZԣ׻��%;b"O�L���3ќ�ه��GA�
�"O����̄+<*��y���M[�d��"O\�����uw|��s!I�>I����"OМ*��=��<)�~1�\��"O�h0!�_�x�d�jrI�,"$z
�"Oiٶ��a���$��D.(��"O�����l^�� ��I�aRl��"O~]��O�� �&oU�G���'"OxI��
0<���"��Qp��`#Q"O��ќ�T(:�*�$�6�""O��$��|�
��Ézh0U"O�5��L&dl���⇪X�hXT�>)����T�rCP�FmF�t'D�I��O2(V!��9��`�ϝC�� S����'`ўb>�i��S<<dPE���]]�ܵ���:D�Xk�kF	�D��[�j��y�w9D�pa��#U(�c	g��A�Pm,D�x�!�UiU����g
9C�`%(3!*D�2A!��k���'[�fw`)
�$�	j���''�B�ِ�VyF¸��G����1��*�_��TX�u�Z0P'���	�7��x��|uAS����>,tC�	0�̲B�-r�� F���S@���퉬m��1/,	�N�
���,#!"<Q���?����D���2"�_a;Dq�4K)D�L�wJ�7ޑRRa@:q�͚q�%D���,O0>"�H(A�� �1�
/D��ؖgM�yh��E]�8�F�+��7}b�'��y��Z]�@���O4����'�T� ��B(`vl��`�"4q^���'e�+TK06�8�C�M��ZMk�'-����b.���{So�4j���'[��pT���2YL���V���)p�'�T�[5��8�)N�+�I �'�� G��, �p���2�jM��'��8�&� ]0d3�C_�5�dC�'���R�f+�8��!�e��'RF��dS
��p ���&|�'��Y#��5����l��X�'��ez�ʭ#���R������'߄tʗ�L�G�t(Zw�D�L����'�8U2����`���#����'�аE��(2-�e-1w}��#�' �yjt��Qu�|( ��n��#O�pw`�~��t�o^$���0"O,u��Z�T�h�N=f�`W"O��ȑ
M�.�\�-�GΤ�"ODMxƅ�s��h�!lՋg1�"O����W1
�! ���$@�zY�r"O ���P�ёq��?��`�7"OZ�J�B�{���˖*H�%���"Ol���Y2�J�GiI�g< 02�"O&�;B���R�2�� #��pAe�"O�:ԃBu��Yɥ!�/	5lp��"O��;�T1~�R&�ЬS<�!"O�����(53
pk��P/6	&�%"O���@KӢHDq�cMek�6-�U"O� �E����3����E�G�4�u"O1S@FC� �f�0�$(:~�r"O����	A1(d;e�N+H8Xx�U"OYV��E�0��b�A3%���"O�(�d��'��-��\<@�Ȧ"O�ܒF�O�:�bb�ݖY��:�"O�!�E+�-R!�*��Y���`�"Ott փ���B0)r�Wo{�%��"On9
3G�5t�Gh8TG���"O^��C�T�©��ߟ/�=��"O���R*��U�^)n=+�"O�@���U"[,�ʡ��b$��"O~-;�MK# ��+�j)5�~�A�"O
��4���2q bdP��<��"Oq륩�T)�8�$�M)�5�2"O08��N��~9�Y��~!r��y�!��Q9k�}P�V.R�l9�&ZI�!�d���p�K��?��5cW�N0	v!�d߱,>f9���:|�Rp�#Xt^!���<q�3�NY�X� %��4H}!��\�Q��e�&Z�2�����:b!�d��2�P`Cj��D��D��!�D�#=+��yJ��~�N@P�D�!�d��CXv��|`Q����`�IU"O$1R��B�l�f-� I�9@��<��U�~����j��#?N���GJd�<�*�8(�MQ�⁳�X�Ȗ
L\�<Q!��L��p�BT�2�@`�bљ=����ˊB���R�@&t��˱#�	��pkc�(D�*�mѲM�R!@w�H�.ӰԪG)D�@��`B�\k�<�0�ДP��tp�%D�tA)�`G�@���Pp�s��#D�pjSa�=�ҡ
4+W'<�
�` D���'�M�F��Ĉ���@��>D��"�� ���5�ِWI��ࡌ)D� �jZ�V�|E���M�r����-D�d�F@	,��#1�M�Vn2���(D�,PT� D��Q��&	x8-��N0D���T)nE�DK��V�#�5A�1D�`���T�@�Λ����Z!,D���n.l�D���$�;%ʢ�� D���ծ�!:����f��1z`T��3D�<�vL��E�Ň�bMxh��.D�<Z7 �#%n$l�g''j�2���/D�LsJY+e��Db# ^�I�:T	��1D��@hD� S^��l
4XJ>��� .D�8#%�%`r` ��I4�� q!�)D�x��eP�<m�\�U@<Q� ���-D���ʚ�� �$A4;Alh�A�)D��KrN��>��<S��#r��ը)D�8����_�q���	. �P�f'D�Lp�NR�R��G��]V*��d�)D� 8«T�zj�Xa���y��ɴ� D��Zg��*����.�8,�h-D��ڧeV� 1D��ɈX:4s�.?D��8Ҍ�2�a�@�F,8�ڤ>D��qu	�~��@��;��L�7`?D�8K�jS�F<��C�8[f����b'D�|pa ��9�X�d�0`�"�9D���1��/G�(�KG`�?OZ(��"D�H)d�Y�,�����"�P����"D����׃3�l(�5�X�L��"6E'D��Y�D�/N� Ke���!��I#D��bdQKX�Y��A���!D�� p :����U�8(5K��>��) "Ot�1���5���cbS�j�0�s�"O�D����JY��bc�J�-���"O���_0���*C�]:��A"O���b�ŷC��=����Bh���P"O4q��;�biB`�&F�r�"OdI%��<6brb�6wlT� "OL��,��l_�|�1V�#(�sF"O��+��q)Cd�"ټ<��䛝�y�i�>Q���X�nί 窑�sJ���y�.���" �7&\|��?�yR��3bT�C��|������y�h㮄3"/@Y*�M���yb�W�1ǅ�������j_��y���&�Ĥ{��Kq��xvB��yҩ�bFT�b�o�p�`�$�)�y���SL���Ņ�[/4e:.��y2"G�a�A'1Q�>� F�W4�yrh��*�B*�O�0N���e%���y,�(2I�%h�ӑ_ފ	��P��yB�Ү�(L��c��g�bH��eڃ�y���:vcT�)oA�Za#�N�y�ՐI2x�X��Y��,�2bBİ�y�KH�v��̍I��Tr�$���y�h�Z� iA͢JYn �q��1�y�ǚ,=��a�D6rj�TaQ�N��y¨W����еd�:��4A��N�y2�^'|S����ȇ.j��1�k��y����H\��%S�J���`����y�7r}r<����E>� �����y��i犄�2*��D�̙ǥQ��y�%Q8!
����Ƽ9�r���Ԃ�y�lH�K��x"�LTd
fA��_��y�����8����$c��0�v�H�y[�������j}|0���yb�g�"��T�Y�T�,�����9,$��qF:O��X��=O�:��*� #<���Nx�a�m�8������o���[rDWDq�c$��=R�Y��g�y��A��-8D6B��c%\ذ>�e���R��C-Y�o�%�&&�e�'�d�K����H{�(�z����Ai9*�Ji��e����陀o6EIbe@�U�ҼS��O�x!`���Tm��#3`��>�m�����"�JͶpc�k #&1�D�b�����` :����8�C�R�NG0�R*�7PFi�w"O��qL�m0�B��L1'N�@r�m^�sH��^�2WJ�� A�pv>���S,p��0;r�O�c��N��#&P�5��=~����$Q<��|R(�G�x(����b\sWH�81���R t�␌6s��i�c#�/�0�02���tp+���8�Cm�+��0�E5�F�<Q�T�����R,-��X4a� �T]�0AJ%j� ���	9&p�-���^��Dp�6*Q�=͞�s�;�fN�=���$�J��򗤘�oF̉J7� 8���k�yF�5��$]+s�XY��O��!�'�Y"jMةrga��y�i�,lb�� �L�0唱����30=ƘK�⛒��<���Q�Dꔜ���QU&��nJ,w �#Tn�KD�	u%Ұ^����qݡsFSBeXm��L�8,:��I�_ô(#G�:1��ZP��Y)�`�%�'��ғW� �f=��昋��,
�L�#�H�K���;h��qh!��j�m�c�h9�c晉��RٌAb�ޭz�(��+${(b�"�$w@�r�a�8�(O��+v�V�!p><:6BN�qO�$
w�[��ԑ4)��"�<+8���O�0�nd;S��D#�ɻ��ȉ=�<��3&�iTX=(<���y��=X���;7�]�vn�পQ%[�\ݣ��O=w��a���	h� a�eHԾ_���C��x{x���*�%�y�g�=k��ʧ$X#r�>غe�U$�ѓf�+~L�b��/(V��H�g�'�J!s$�יFz�13ᇣ�@��a��0A�d�	�5n��m�B)�SG~�-0s�#�uGgǱW��SA�*J)��g�J/W�jDh=�䬲דҎ*!O�=:���bP�ݤ@�����G��	a��.��ib�JIs��91AN���r@���B��ܹ���a�ψ��歒�(�r$),��q��D���<TU��� '��uY���n���x�z8s3-MAe�z��q�@ ��뇳6��X@��_�T|x|��D�}�l3C�����I��$�n�'_1l���G��|������A�̧u� G�Z�
7�;�`R-?�P�`�!qk����ONv��dZ�W����K��+�d�:�W!9O��9� [�z�.i�H�/�uG�	m|��A_g���6�[.=����6g�?&� �hb����������е7�HQ�u�R�1��<� ���u��Y�j�C�K(m�.�hA*��]��D��pQV�"dEH��(���+
~�9x5Հ.KL(��J��lx����ۃP_L-�rd�J�����*	x�!HU��/����HR���"�3�P$�	�L^��f�D��J�a�P Shpi�jPme�������I��������&߭_�\q��_``I�
���'�~2J�sO:� q��"��p�����#� ��K*t��UagD�|8�� a��]"�2�"`�ԡn�6��2�ܭ!bI�(A\9�V	��,�3�>��Nð}*�"[�"!���5Z!�͘Ĭ%vy41��4e3�(�N~RT�%f4��V�D:�\ �(���@�����ӥ)�P  �h+�ODl�ǂ�|SR���UM��R7i�z+
��Ŕ)I$��h��Z�t�ld�7��~TB���OVK���O	�%zs� �C��]YKHN2"	ϓB��A��πOA,$z�أ5�T�9BM�r�hA�gY��x��/�a%ؼ�@'y��A��'��>�	Z�ڥHU�x�R��?��O�]�PEP�br�K3�ʸD�����$eE�{(��H%_�q+$�]�zS��cm�@�%lP6@V���'��mP 9�@�M-?�&q�"`�'Hҵ���Ӏ����3��*a
 <� �6	 BN�7*��9��n�ؔ��D'tj�����a~b�юt~H,@b��[��eR;@�8���E�!� `�%* �TN.�#��ÁY{\ �m��]� ҧ���Y�p%�`��AO����N���O�����9�``��=5,�)��\�.ڰ���u����a$�ipp�I��C~�S�O�����|�:,x�&8���+O������+��@+C�ϢA�����_/
q�|�Z�$��v;\\��%�!�^�%"O���	!��Ћa��/XV]b�S>�x��?S�%�Ԧ 㼵�E�	 ��ԃAeZ��y">�@)����1l�����$�Ƞ�4�'�H1���.d&J�!�[d���d��Y|����#1T���fJ-J#��I��)k8,2s��\k�غ�����
�@�\���P� �0a��?�D�P��\]C�D�+|͚ahB�֨KD�D�˕�t��t��'W*m���Cd�Ħ����U�m5��z��S�qK��?'���r�q�A����Ay2GU�~%B����i���tOG*vP}����%�:!�6�\�L��r���8�v��@K�(�~<���+T;N����f�"��Fo�o�0�+�Nމ+T�V�Sh��e�&�ӻS��0!B��b�i��~�:\cĩ(u�X� Q2�3��א~��a�քV�4��'����E���뗬UƬ�R7lH�i�Z(3�r�j,�uÀ��ƀB��j#K�/S��G�H�~rE�&uΕP`nL�W���i���O��	'b@;7�@8��%OE�l��f	'1R4�c�A�r����c'���d6�ƋEs�0���=s��rD@[-Jh�>I秔gp`iv���fțb��HyB$Y(	AH��яK:	,��Q�g؞\A�7�	�\4�aY�Or�� �>;nT���(����F�/	�����H~�a�O.9��Q�̉P�Z����1����3�4�М�j�,M�'�ĸPuJ��1닟Yj�Mi��'[j�`�@�o���"Q�i>@��k��e��i@! ��juޘ����s����'��i�MF+<�n9�GlP�
%�Ji}��	0��|3�H  ĉ#�U�{ �?��m@" H�M
P����dM18�q���~M!����Y0(P��G^�gm"��I�u�����C�Zx�]F}��)B� �#���lS|`�T@����7iF�m�	�=�X=[�j��M��`�����,)���u�T%2d&n�楻��E{^9JCD$Emp-�V->�OR s�oDS���b�`�l��p0�E�"�X�I��ͭR`�F��L"�i�إ�E�)�2����t�mk����vFhp���
9go2�<Y��:� ���T,�8�T9�T��J����6 X ���z�!Q)QsN�%^+^�A@���(v�Dˡ�Sʟ�k��A�շh�ay"�T?%�B����)j�,Ei��7N���#M���7��9M�Q*Cd�>��$SA@Oh8����$3EQ��A�بM��($	�<=�<9�SD3�$�<<�4!��d�@����$ �F����+R�>H"�T�Y<7C��$Ȁ�d@F�*@��#�L0I��~B�� *[Z=I�(ޫI?,�h��70R��E7�쥪��C �f}���,V@	!3H�)J9$����y'@�	~j|ۦA�M^�}b�+��y"�U2]j�81ߓ6p� `>?D�e�	�7h�!��_� ţ�'\i��3����s�	����} l��$ץHՐ�XE_�rc*��� 8¯G�3l$�S��WJ��a�O'%����.PJ@:�I��M*�n-X�x]Ie`�ҨOzd��-'Z��Y",J�Y�tPh��I�~l�!Dí&^���6\�nd �O
���#g��3v�U8?�~���}��(b�JEPi�A�5N��t:�!��t�0%'���4 ��h��I��	�/.|���M6���ހ�@�/b~xP
��C8��S�"O��J��
+6���Gg�2X�PC]�`h� "�,v�I16�C�3�hi� �O��ⷌ�/�>`q%FҚ@� =�s"O������])p��G�� ȢDY?l[����◙"Y`�i�) /L��ˎ�dE�d��(���E�.VD��4-����zB��P�.U{�n0��T��"{�6� w��Z�H9+���C�<�7�'�4�z"�W��^	��TX�Y����Q�
�y�� �'%<�2vo4�ɑlV��{��g*r��
��!�� �Ar�ёx
1�.�0q�V|v�Y�$uٰ��o�:��O?�X�~��l�%I��L�*�2T�K!��G� "�qP���B�(A{�'��bN���p<)������(���\���b�S�<	�I	�2s�4��
���ps��Zb�<y�'��o�����%3,|c���c�<�$M�b�.U�t�W<����� ^r�<�5)ݸ�PDI�����h�b��`�<QR@��:�yBF�I,����_X�<�K_�d�Pa���T�~����m�<��X:gQƥH b*X5�RF�e�<)R�&y���V.�*qt\��b�<	#,I�Ch�R��P ` $��%Y�<��K�r�f�4e����X4AU�<��K]�%upd�fLa��}��CIQ�<�w'y.�����=���bNM�<�T�Q9m16�El�3*��H��SN�<i����Y�|�9���$j�
,�g-�J�<�U��:��tz�n@��<	��B�@�<��HV6V�� ����f��T���<�^Z����N�8Z��h�$e��C�I�/}$[�
�� ����SxC�	�h�,���ɃaP��QOΞmv^C�	31>�Rs�H2M�����O��B�	�s3)���7-|� ��Ͼ��B�I�S��t�KF$Ӛ��Aϖ.z�B�I%m�bI����sڴ����>D�lB�ɑ[Q �
�CD;�H8Be*�",6C�� <މ��:�| )C�+*�C�I'~�!���O�?�mX����$3�C� ]��m�UC�5v�1� gC�*�C�ɱx�XQ�%G��WC�e*��e�(C�	�{��e�F�J#cݞersOf+{<C�I�mm�邀A_"�fy�æ��#D�0�3cl��պ���~pNl�o%D��Y�%+:�.����R:_�c�9D�$#��&#<�!��m��8Fa7D�D���9��ڶ�D/��b��+D�,�E���J�q�2��G�����(D����Q�B	�r腉3p|e�)D�� E��`�r吔�@"g��U`#a%D���Қ6�4Y�̓�+�&ܡǉ D���gOs��ps�J�T,�i5%!D�`�&)H�<Hb�AWņ'*|R$M%D��R�+��~�n	�rkX�� @�o D�H�vjV�J��0�JW�h�mP�#D�\A��
=tztDZ%.٦qը�#>D�|�'M�u���''Y e�hS6�2D� �t�h�$p�ʗ1L�8TRb0D�P��T�/��ɉ6.T?�|�0��2D����rs��H7�.GL�C�A1D��F
K�H����A�G�_�#��,D���aς93!��%f��{���{��+D��U�ڱ��mH����A�8v�&D�ర��7d`�30�\�*G�9�$D����/�4�2�A!���^Z�����"D������"r��C�a����k#D�,6�Ф ~�X$��"����W�#D���#��]�j���P�U�Cj%D�Ȓ�d҃d�tM��)_�N�ͺQc7D��B�,_��;Ӣ�r}���Em1D� ���Ѹ�0��H[�h�A�p� D�LJ���0��iX�u�la�`#<D�tғϋ@����̙�!
@�#C.D��   r��ĖpN ��Y������"O@��6b�#m�����^���b"O��)�I�x� �*��G����7"O�1�k�7b�
A��z�$je"Od�f
�v4��F�L�q�&,�W"Op	+�ԩ'L�'��'"�Ƅ�"Oژ�����F����b���"O�	� �O�p�xLi@
ڶE�ؐA�"O88%ɂ5��%+dj��:��ː"O
p��iX�~�j`���@�*�^��"O޵�-�Z�h���$E���cw"O�Y���a#2t��#?q�@�"*O�|K�E
��h�e�IOr\�
�'�jF�1UUډ1@�\~�
�'��h���5[/��B�\�=y��	�'�"@�	�mA�"B�C��
0"�'��pg�,$T��?n�A8�'�ĨH����r����GG�<P����'An@�'`�s�FS���:(Ct�{�'�X�a��
8�>�bq�]-��
�'��Q҃��O��$z�)�Z�d�����&�&Tt�T��G�,���Ҧ�s�<I@�ɔAQn�k�I7.���F�l�<���(|���޸!��;A,Sl�<�#W�3�r @B�JLX���2kP�<q����9'|���[�֢Q��J�<Y ��7 Z���̇�3�)2���J�<ap��"h���ҍ/�:�aPkSD�<���V ���Ã�Q �ᡐCB�<��W8*ԨW�8C��)�d�<	tk����U*�9
�S�aj�<��#Y��釠��ɲE�Z}�<ɶ�u�D���[�]IH���&�V�<�eOE(��6�����1&'�L�<A4"�T���B�>Q��L�r�<�����1���� 5C���裦T�<�e��Q!���b��v��� P�J[�<y����+��� ʜUe��*`gU{�<	 �{	�����dK�i���Y�<yU����4mXp�Y�pIP��CƕV�^��'v�}�DU,-3`T���O�A��*2�Q��!E�"̸�'`�#�(�P�b��Y9T! ĪǈÙ]�r�ےN�!ޖ�[%B �OtyqE��)c-��RcI���D�P��ɗ\ZV�
�
%��@b�� 'S#|�Ņ�=}�>�Z��p��o�;������í02��$S�q6��Y ��u�T���)��F;9�D�O����)F�ç�d��� ��<: �~�1!J�1��:7J)H�Q�x��mی@A�C�N�PI҅����iҞ`y��ìN�Lup"eC)=(I��O?6�ڴ	�$T:�� RԼ��h�t@ ��A�8au.y8���dջ��� �GDb��DE�R���h��45h��$ǸKn@��O
y���q#c�BOt�Gz�	ݾi�,xJ�b�]^���#�׸�(Oz���)�o�6L"�C[S����:����F��.D���m�_X����`L-=��
T��!Bݰ]����@x�3
 ]8�-�SZ ����D&E�0IS�$լ�Hue��VTB��Ñ66qh"͋�R[ 睾DX�My ��?8,2�Hq(Ҕ?IC�
F>)�#��L�MY@N�VΖ�ذDҁ9.��KQ�� �H�lD�Ώ� �:ą��N3D#�w��B�л(܄��C)�/<64t�	���Ę`���,v�@+��߹P/2�s����7:�j���S%�@`���`�"4��tC!l:W Q��*�F�~�s0��F����e%�Y\�j &J�u�+�O�A���aP��/e�\h��J�T�K�e�� �9���'�x���f_�|��0�H��a�&3������y��1m�%�LzsLN�m"0���A��V�`"�N�4��,��"B�y���7��0�5���FJ0)u!�y��-z\�i`��ǋ#�İ�@�x����P@h�x�@LO�8P�n��?ax�d
 �؈����y'�˴D�|w�^��Xǧ�?��>	�'�>T�T{�
�oy�<�W�'q���0���hE�V��}
TLj�
_�e�Y���6ks�Dy�)���dˉo������.��O��a啃:�d!)r���$�Ġ���Y� �5�Lͻ:R������1V���{�䙱��SE���p>y�K�:����U�Z�rl��S?���Tl���B�C�q���q/�&|�X��f�/C>:aw۟�%�T�|
��� f\�C�(� �"O�-�Fj�NCP!�UcP!~�尣a�o�����d��^2	����;�%�}R��G��ywa�`�<�X�k�GZkB��*�B㉰h����GG�|�^4�e�G�-���K�=~yZ|��i�Y^pȷ�Йj�����^��pA���#tQ�B
��3&�y�� be�Ϩ5-�p+W&�^1A��~	2mY�G0tHzEA�oՓ�a~�(��I���	q�޴R��h��ݎ��V�� dO"�<�t�����E[ %�N�i��sU��	�h֮�Ph�+'!� jի�.ÿ~���t��6�>�y�A�><� ��G�hӪi0��6�3}�dG�*�l�!q�ز{t4�f����xr%	8^6��%BD�/��uL�4����%©\-Z�����R�@���W#,<|(����7�^�����*�y�*D�4�H��!�-!n)�#	�'�,k�Hl>����JL��B�I��xx�v��iN�,ha��a��O�$y�肐z�����э+܂�3��$�Q��<"`�ګ9|��3-�C�	�5�*��2ɋ'i�EBB�TF�J�!s
.��d���Ѥ%�F�!d��|�`ݙ_���[&)�M5�MxT�8�x� ݘ\�F`��%]0�QS�V�9��T �m���e��`�0]dͻ#�,,O�9�D�sO�<���ڐf຀�I�@��!�b��mN|�Pk�0i��c�%U�;�/!���1!C�=��B�	XH P�y��;G�O�W.ʓ@��a���9�@Q�0��� :�	�GܧrT�R�+|��)5��.?��ԇȓp-��s'�J�[���F`-�x�s'�غp}���i]߂�\��b���9vp�,�Ui�j����K�O�x�&(��W"]��rWB\S��<iᯟud�YV!5���A����%����c+v9
3���@��,��`�Oz�!�◢2���)4�NB~R�յ0�ٷD��'Z� 0�Y
��OF ��G�/E�T�s ��c&  ��D�z�,H�&iϴnx�rCƽC��E�G�i�"��փCUbЈ'h���O����05��I�]�i�t���P��sĉs �Q�1�S�,ⴸ��l̰>E��x��Z�+(5��N�*-��#歊<�|����J�/p ���K�c�a�'=)�ڵ�g�ަvS�llhF�Ӿ.�ĉ���$tQ8��A��ds0��҉	zO�qJ7e�gvTy�w�(l�U�.i`����P���L��J�$p�����6�clo�6�J"�ǘP
`��9�j9��J��$t�)E  p(-ɳ�W�i� �rB X?9���ᶸ����1(��Gȓ^�'Jr��r��(�np��^�Iw�j�$ո�
�����3f�p]#ȋ,d��`� z;HtLV-m�I�ub̫s
Q���6�u�t���N�5e$��U�<���ں	tΨ�$ꗚ/~�q#��^��O1�L��'VlI�eg��n��E�G�i����&Xp�8��I�^ۢu3�K�y4+�͝)��E͛�4���׃@0"��Y�"�1��#��`m�}	�+��o�j�2b��%HB�L�u�+�O�l9��>S����R�I�	�@٣�H-�~��m��,ǚ�(V�р���xT�	S�.p�"ż���,�qv��#B<&�bH�&�9�'�E�&O�0��$��!Z�a4* ��x��Uj��['1w�� $B�C�%�w�& ĦIj��G/B�t��R�'�6l�b�K�=oDI#>5�|t�+O��15�$��P�a��$
����B��UN��pr�����6�ULf�Z�aףo_\�����>%��U0uDG�r���[�k���xr
K,�8P ��Z����O�	 ���b+��, �%�=l��&�Ք#Plm�P�C��:杄u1�T@�	J�,�Z���E��W�B�I:\H���ĉ�~�v,�@#��6�`)�S�;m@����id�H3&�,`|��w�I�S���0`!G�0d>���O�)�$o��Z"x�	 #�X�����'�B��S���VAQ�1@��K%�v��AB� z��aĝ�Q�Dm�ˀ<(=P'�BFЩ���>=1�u�3�><\��Q�֓O^�&��+R��ɛ��:�-�sc�m.��b�8:�=r#��Y�e*6�8Wy�$�V�!2B����'��Y��!���h���(�f(s7KP&x^ J�kʉEJ�᲍�1q��1"������P� ��?!k�wK��Y��ZK�ȴP3e>*�Ѱ�'��LC�dJ�cW��*B? ��kSɊ�E�r�e��*�>�r.���R��
�`Q в�B>#���} B� c�0,z���#��M��I7&�(a����V,�X��� �%J ���m��lѥ�3-�djQ�A�J!�����I7@��,��p�e�Oأ<����5D�	��/��T��`B�
B¡9��U�IG$D�ӀGTr�K"��^��A��µ>�~�Ɖ ���2R��1M�8G�Ȝ�ēb���n��<�����R�]K�s�)�����3r�)b�
?{O��W�_�C�	�fqVES�LK�I�9�,�$L�yQ�G�Ħ��TaZ!\��Q�D�1�ӾH����<۶AIf�W��x� ��B�I7&h�eC��%LL����T��lc�[77m�E��d�?���
E�η'kQ�� X�h�5�z�BƀZ&f$�|�f�'��9��)�%���Y�"Y�Lu�R��d��͓��Z/+wH5�uT&/�a2E�z�r�ڠL�K� h�f���O�`H��/P��RՁ�'��������W�I�E�[�Ew"O��wF��`��T뇫ћF�����!ze�Q�O�|��q�O?����ӓf�38[@���	��!��Ȇ?x�4��l�4Fv�;��;6��'Gt�+$�Ļ�p<���5��)�X�>4ҡ
�b�<�ă�(4Ȝ���%:���IE^�<�V1<��2�Tij%�� �M�<��N̴`N�5�`� w�� S�A�N�<a���{]��:B'O�$�~S%�I�<!3Ȉ����4i�{ʴ�/l�<�G�I�8Ь4*1�??s"����a�<!���rи��u@�2�tĲb`d�<��Ĺ5)�H��LՍe��)S��|�<��F	%+��Cg��jq�!��y�<!&(�>5�@i�C��-����Jv�<�"]Q虋�B�E ��i[l�<��+E%S�B�y��uR*�c'/�o�<�D#
�btM�����L�k��e�<ce�`�X ��>�~�J��]]�<q�*CV�H�$���Q��^�<�� �yjt�C��C��Q�c��U�<1fa�:5F~�K@�
�t�*܃�\i�<QW�ۻ$�4�R!�L�v06 [�<���M�,h�cH(`�	��Ez�<9biݍ0ĝ��$6l���Gt�<��!߶-J����"��@P���_�<���m�48��F�9N����i�V�<	��;@b`��4d����rXt�<A#��D�"隂���I~`��5��w�<a�U�H�8�:��8!�Y1�q�<1���	V��Ek��J�� ���Bo�<9��5|��Q����B���`戚N�<1�"�����-���^�$����N��<��̰��O1�b��#�E,� a �Z�h�8��C0OZpɲ(R���q�N�"~r��ĺ1bM���3~� ���W�L�s��|��ҧh�J�9N��E���Ǌl#,���2��l��y"⒊�ҕ3  �~��C%�ӓob Q*̬g�����G(9�����r��Q�>�z��1��S}����3Π8SUN�]rJ����t�,ʳU���57O��S�gy�l��B����Ѐ�37_��Pk	�CQ�� hʨ1O�>A�'M� �CFÌ ����1��2���Q��J`y"2O:��&�i9?�SP�U�<�C�OԂ	��K"lUn}�^"}��k}ӆ��-O���D�b�X���D�E�x%b�ʍ)���ߦ�RԨ7�i�5E�g��.��i���	I�P�`�m�	�M�ǵi�c�"�D/K�E�����j�pH��]�L����=��."�'��)�* ��43�䆇N�P ���+8/�O
�$��(���ӕ �%RN � �آj�?6*LO��e�@�S�����r�Rj�SA�]�|b���'��dX3h���姘O�|h�t�֧�άS4�ԨW����%�ZF�z6͕u�����^�Ah䉇'�ȟ���`��℁�6K��F���E�. �S�X��g�(��i�=9 q��N#V.U �� Q�NO^$��ǥ@�4���S��ar��k�D������D�K5\\�5*�/D}��H�v%s�ɂ>X����g�0O���'�.�EΎ�ɧ��:];���}�RQc!@�"�!{���C�DЧ5��~���􁌽/6�)r��L����6�{����d��|�>�OktDy�"V(�)R�`H*<��fG) �̓�M#S�ç����ӻt>�m�������q�s�ܰйK���v�ң|�'�`�:vM�nG <2�N�	fՠY�	�'S>)k����<@ 3`�,8(�'J6����@ HT�5eӠ��'�f%I�*Ɨ:9�y�c��Wf�'w��@���x�j`>H]H0���� n���&V�U��(2 ʂ�P�E"O�x�T�SP<���d��:v"OB�;� �\�J� ���B �-(1"O�-�d�qn�p#��&"��
�"O:B�9'd�t��2���P"O� �Q�K�bq<9�k��� ��"O�H;�a�%Yd�h$J�<ب}"O�<;��Z�Q�ɪ4���o�����"O�P+�њ� Q�t+��P@��"O��k��:ԙ���	5�x�z"O����&��!�5c���|�Գ�"Op��b�>�X	����!�#"O�y��;"���r�鈄p>Tm B"OL!)$S�n���E��]�"I�"O�D��HX|Rg��X.���"O��Y1f������[>W�- "O���X�g�by0�1�EB|�<��D��0(��RԞ�� B�<16d϶6}����JӶ-�pɣ��T�<9%h�����3���gcAh�<q���) =`I���'K�W�uRnB��1[���!�H2t"�fSX�6B�ɽwj0*�EҺ{���VP
@dB䉭{�����'-�J4$�.P�C�I55�I��� 1L � 1h�� zC�I-"�8A:	0|��$[{s`C��3ސ(�ҮOY����SȚ�}fC��4Z�J`�c�"v$8��J�8f��B��3|��+�G+��M2w*�� �B�IxL���N�id�W@ID.TC�	�?.xB���-s#�,���BX[$C��<c Q2"�_�5h8�`�+d6�C�	�%��p�"�8�L� ����C䉗 ���0#�Q#x��9@�;!/�C�I�4 ��3�UXr�Ϫ]-�B�5/	���7ΐ46���2����TB�Ʌ
��Q��8���i�fŋ,��B�I�j�1`� �RZ�d۱e��xzB�*?0*X@!�?%���cd�
;�8C�I�����Ȫ'e�}�� J�mF�B�	�?Ф��4���[ȹ��+E�7!RC�I:[R���`m������4�C�I8��5;��ʯ+��zv��<=�C�!F�4�aT(+$S��ȣ�!��C�I�;.a�� �~	4]���Q�e�8C�	*UT(8:�D\�r� UC�ZC�={�|���G;`��0��&"��B�	�Ҭ���I��z�!�_�&B�	K���FK�P䈃��X�J��B�Ɏzb��a�g��3�|X��(��7��B�I�>�N�*$�̷�f��	W:��B�I�z�X�AhM�H��jG%bB�I8t�T��d�O-�2����%$�NB�Ʉ7����O��|���_�]BB�	���,��böv?����Q5JnlB䉋|����X�P�H�Xp#Q��tC�ɔ�Z�A�G%s���ŌN�P�C�I&p�$�`�9r�"�b�Ȗ�<��C䉚n�țQlO�w'������o3�C�	6	T��Y�%� ]3� 2 �R�!�6C�	� 8�q��K�-� ��B�"C�ɝ!�)Su�^&�уV^#�C�ɆKy���g�[Zp�pu�3c�XB�	;$^H%�$	��rN}9A��/�C�)� ",s�L��ba�a�E�F�P�����"O�L��V�P�A�!O�]@4 �B"OVT�����dJ�e�_�9��"O4m��ȃ�&��	9A$�S�T�[ "O�єF��\��e蠂�"b��hy"O�(J0���f�^��p�s��h�"O�C�/�2g� $X4��7�X�"OBr�k��<b�xa-�w��s�"O��*V#Q��@8�k�N��I1"O�Q�/��F}z�j�d����ks"O��aO	.x�b��#Y,`$0��"O ТFA�#�̘P��ג ��$"O �s$�ÎBƜ|��J�f��`��"O�t�aLFQӖ,��Ȏ��"O9pW��5������CǨ�#"O��3��}�9��I�����"O�h	��>/:�1��H?��;�"O8H+B�uf�L�#"ӴA�Ёe"O�]�Vɛ�	�1��c�e$u��"O,�2	+(<���H���;�"O�	q'W�,X��{@I����hV"O�����M�D�jx� �W�yQ�"Oz�$� BY���ݰoі��"OBX����ɢ�Aˉ:Ɏ�6"O��Ө��]|����M�d��Q�"O&����3i��
� L$��F"O���l<8����$��?5 p��"OP`)�W4Tw��!�N�f-�c"O��°@��`z�Z�� ����0"Ons$�5#�!��|@q2�"OH%z����pZ�$�$r,�q�"O=)�	�J����Q2F[��SA"O^�`���w]���qń4U@L�d"O����G��B�JpNX�_/�!�����8r���F<(� ֧S�!�DP�����A�aK���D��[�!����̐��;� իS�?%!�V�^�hE���x�����1x!�$K�'��:��4���2���7�!��xВ�1牊mIȘq)�K�!�d�\0�����dIӍR��Py�$ҭ�&�kcH�!s�&13g��y�@	mB�EA�L�w `�&jG��y�i�K�t�� A�kd�dц��2�y"�	K���Q6(+gR��^�` �'�|����/8n0����J�f���'�@ѣkX�V��s�Pa�ey�'!J���נ%�j���.Y����'th����W���Fc� X�	�'[ذ�r�R�>��	��,�Xz���'���	ϣl<P�f%	��f��'��+ !9���# ѯd`���
�'�̱K ¸&߬t���İZ�h�
�'��`�bT����U�����'en���AOE�$Ia���F�m2�'�E^�>��b����1�DQw�<�A�H�&+�%�`�Z~60j� �u�<Q��O<9.h��g��x���M�o�<�g� j:t0��o���DA!Nj�<)��Y�����𵲀	qe��0[�!�dD-��B��Y�	�����j�!�F:x��⇂�=,D��aT�,c!�͊TP$�tb^x(�iV�"$!�d�&<��a�ĸm� ��c��!�� 4ؙ'�.Ha��%br�
�"O���$��w�r8� ��h?
aj�"O���EBW<�AZ��Ɗ��0"ON���$]�G-&���"͓ ���C"O��:E��%*���� �'�܁�"O��E��O��K笎�^��Y��"O`�A����yI����H��ը�"O�X���I�Ԩ���Bq��I4"O�,��jC-@ő�G��aY���E"OJ ��aǬS:�����A�Kh<2Q"O �%�HJ�U�!ϯLFlh�"O������3�PÂ��� "O� Y/ؒ�u��oY��!�r"O��:���	Do@���H�"O�)����1?��M �o�o��d��"O[���bx@�R�.
X��qy�"OR���IE"�h*P��"P�����"O�Tsf@y���s�co0"OJ]Z���Od!R�f�;YXp*�"O �aCK�,�1��'M<����"O$4�g�3�.yI� rX�z�"O]�@͊S���`ğ�O�p��"O���s(I!8w��G�2$44K�"O�u�JK�*���pg�h� x)�"OQq���-�L!�p�'��9�c"O�|�%���-�b�1�dĄw�X�JF"O���cF�+��#w�	|�૓"O�U!w3A���0λ)ͼhP�"O��x��E���sFÀ� �"OdPI���g�6��n��5�(�8�"Ob��Ύ _����ލa��9t"O��P� O�	�"���d8	��lS"O�\$)�/�x� $�� @�"h 3"O���eJ]���2 ��2q�"OL���X<K$ �P�.�,[��r2"O�I�ѫͤg%	��-�fYa"O@�qEM��r�6��B<F�F	"O�|����X���:Ѯ6C`x��"Oĺ�ܴs�>�`�m[j�!"O�X�(���Jq4M�13&��8A"O�D��\8]��Q�T$����"OF,���A��$�Cņ��鉤�6D�0��eN�GTRP�D��T�[��)D�L v�W&�=k�I��V�	Sg(D�Tзe�'�BL�$�F�1m�pX'(D� �L� ;�d�ѫ+Ѹ�:Qc0D�t�FGW�Q�u�G��cf>)�s�3D��@3*E.'�ā���#$��S�7D�X��/[f�����[(�Y�Q�3D�v�� 'Dl����! �Pc�1D���g�/0;�q�T0�8�r
2D��˷���1 �d�e<:n^QC��/D��{�
H(*I�y�v$B�z�|����9D��*��%����ը�8KFX�`6D�@�� 3F�
�F,�42�H3D�@��A�?�6t��J*:���sb=D�L�q'�$j:���f�H�4��c.D��	�΂+k�����%֦V��]S��+D�t��Z��1q�ESX�}���*D�$�W��'�D��a�!^ot�)�(D����쌒]��*�$ѝNXY�7�"D�(3�
Ǚ_l�z�Ϸ]�8��ħ$D�� � �Q/~ �K�v�$�[�#D������lAd8`� !F�.�1"D�� �ascG	�9y�k�TX���"O\�k�   �P   �  �  �"  �-  >8  �B  �H  O  mU  �[  �a  Lh  �n  �t  {  Z�  ��  ؍  �   `� u�	����Zv)C�'ll\�0�Jz+>�D:}"a�ئ�Pwas����u��h�ӊtiB)�FQ>�\rMJ`j�UQ�eҐ-�n�X�lX$�|I�Nĺա���z�-M��"v�

iC�)�RA��rT )C���>Y*��U픟��L�Ũt+���5� _wR�T��O�7ЖK�rm8P#7B*�$�%�!L��	B�&#���ɭo�l�8��O!_���9ڴ_{�I���?���?���sN��"�1i�|���2W��]���I��!�Q)kt����Z��MiH����?Q�6!�������т�"�~��ds��?���i��_�h��3<�֝7c�t���n��=�ށ0%��к1�Q��R���I}�>�ΝH�'G�06�ͧ�% ��_��;1����	�<yH>��'g,pA5����Χ-��� A��V��d��_���Iϟ��I����	ʟT����@�O��Λ%$߰�Е�H�3|��q�4/��l�R�m�4�M;sZ�x��4^�1h��i\�e���]7=@�� ���.?�V�Ҩ�&FrD�a�>���'���)��;^���F�;��bDAS#9 嬻�u�k� �,�؇��V�x�QN���b4
Ō��a9.�lӴt�֬wӲ9o��?���&����(X�H��8C�*�,�����N��j�n�8g}LeyӀ٠r��i��#]�PR^�p�nU
7���#�49s�Vt�̝lȆ0}Xe�#%� `z6�ϔFXMc.�# ����4 Λ��d�V��3SA2 �� tΰ�f������A�E� XJ�񚆧���aM�B�4l��M��i��`����V�
�<)x,�E�A�Q��e�PO� E6��
�N�,�6Mǻr���wHZ�el�M`GeY�|�z��&�I
ʞa�4'��Ҧ�Q�f4H���	V���?���?i��i���'�SU�O��y�`$*D�l��`�''��J��'�r N�{�TٳF�v��ك��u���7*�f_j�a����^���Ʉ֦��2*&�ưd�2���cs4)�����M (�!<b�Sħ۱{����P5��@���(O�p��]�l0.O���"��KԊ� j��Sg����'3��'��'��'��	��� ը�H����O!$ی���)HD��*G� �E"�X�I�?���|�g�'H��H���:e�:���H�"=����D´j���l�柠�Ҝwtح�e��)37T]�F����?�SfX�M+�%C�R�* t+x���?eCS��i�!K�}�&��1��K~�f��^�!�dͶBp��$b$L u�׸�( ��$�J�s:*a�	��M���|�QĈ7�XA/z�ֈ(�E�������ǟTG�T�/@��q� ��� � ��O��lڷ�M���t���Wv�س�b�9D�S���?v�&�'�R�'��{W J�3�2�'dB�'a�.�����gCD��p��G�x���ߟ�%Hg��|�5�T�)�,p�AEz)D�/�;l�������M[��țXq8e�|�<1W.�<r9�p�V�B.yS����I��M�Z�܃�(�O2�I=&��s�nS�U.>���N�!�. �����F{���ԕ E|a���4����f%e��Ah��	j�f�O�	�\�?��$s�(��}���r��I
\�^�B�/�5	���ӟ`�I^yb_>�Χ]DD�!C��D�h��(�LSl �kǓD�Tx׊��`���0)���␗N�(!�!�W�H�0V�$nZN��'�~��Y�`Yjձ6�,�8��q$T�2
Z�○ɼ`��d�%J�O"�oڹ�HO��|x��O� m�� �t$�I;w�S��`�I����I��@\iDA�1ɶyp�(˟O���OHl��Ms*OT���N��)�������ʓ�L���ʅF��!p����|��3M��l�Iٟ����-̐��5l�V�4H 05^<���L�7Q�Ab�F��j|Ήѳ��R���aj\�G$\� IH�^�Ndi� �,3�\	�]w�����V�*ٔp��%��D������q�I5D����!Q޴�?yPb�lL�� b������)��$u����l���>9%dT�2��(`�'g	~��� <O���<�iLU����1(.&A2j���D]*5dp����æ�c�H�*U�J�⣮�Xyb�O�D7������A��4Ks���2(�i�O���M&P�aF͈������q��r���	�=g4x����;��+4D�0���0Bb�QD��&HTΥ ��H\_
�t啛G�h�5E��?U��N�/s�ۣ�Y.e`~ha�C$?q�G�ҟ���4Pk�O�1�(]y�� �F�����	N����|��'-�'���'�#0��h�B̐XFrوbI߯>Xl�A��$Z��l�̟y�4�?1���;�x��5 �6`h\ڒ�'����'�2�'Ŷy�@�C�?{��'�R�'P�N� B��$�
H�s�paЀ�K7@H<�!e��x�N6m��6v��i�.�|B�ě�i|J���h�� JՆ�4$�T=���z��ͩ2L�eg"��Iȼe�	�)i�!�d�M>N���,Tuoڦ���(����'�B�'��vOщ���� �$p���Q7�|B�)�'�؁���}l>[��h_bʓC��f�pӤ�O����"˓%8ҵҶG��8��1z���5Ǝ�AT��?kz��'���'��I_��6�ι�K(g'����%W�.`���]}T�e��3 !2�6.<O�t6�J�6E����p�ġ�3at8֮��=���J"��}r,���ɯ��A�p��5�5�e� e� �l�O=m� �HO4"<�挪<��0��,	K>��7jB���&�������F{��DobT�eeZ|�Ā�D4	2�fӪ��Ѧ��޴�� 2��m�ߟ(�C����'�OH����2pȶ���}yb�'�"0�F-����$�^)�E(P��7�<� 5#�E66�l@�\.�$�!��'`b	 g�z��Q��C1B�P�Q�R� }X"�	*>H�VCۨ\V�呋�$�G«g���'�zuy�%[��y�	��oI���K>���$'�I�?�\TZ�_�b�:xY��ΎI������Y�vd�6"� ��O��e�L��fJ�M;*OB�yBA\����	����O<\���'�^�ʲN�<5��`�gTN@\3s�'�"i�o�!@��=�˳� �X맧����Hiq����a�ŏ?U�I�{Uƀ1!ɒ+tL���2TW�����B\�� 3s(�*h1�`1�TK~�P��?y���h�p�D�-r��J$ N,n	`Q24��A�zB��2n�Q$/�p"�QgA^T-B"<�O�aFzrcA(İY+֪H�X�<T(0O5cd6-�Ol�\��T��'�?����?I-O�՛F�ߪ��i«΂D�b�	�äy,6)�S����Βզ�+��i�?	C�C(wpik��Is��h���
d���2��h�K�P�*��|��A�P~�_"5��Q딩�9�pT��g�+򛦏�<Q��������\�L>QC#��Q]Ҝ��6�(��H��?Y����D�O��?a�']8�-�0��z�e��h?�*O,o�+�M��;��T>9�R�T�R>W�D�!t͞e�16�W	H�t�q�`��D��'�r�'��ם������|R�A�4HA�Šd�ٮaz���⎐ HŠ�d�yf9{ea̝��ѩ�*�/ڣ<y$�SrHH�ψ�F�|���	�L� U�N�g� l
��CN��Hآ��dz2�<q�'/��L�%�%x�ֽAS�������2�M�&��s�'�B�(`d^�>a���N�R���{�'��]��B�?�ڸ���|�KH>9G�i;�U�����H��M����?�WʰE2͂����b���@��#�?����J���?���y#"N�3^̀�Q���Zt|�
q�G;zmh��:a��!�����0<�#�M�r��rɝ�^zt�E�?{&�(o[�I���Z���>A�DA�4�v�j�<q���Kܴ=��6�'E��0îL�m��lQ1K?j�^t��]�8��g�S�T��D�˗'��<�B#��[^~���5�O�n�+J{^1��JP�;�.��ə�4���˦A#R�7o�O���|��G�?�?!��L�(�|�� �Č�j���D�OB�b��l�ՑMsT��C�J%Y!�,*@�8mLE�7�ߗO#h,у��W~�
B#�P ���H�U+�48��xZa��V�IǔWZ|�q兛?�aǠ}f�ɶ~|���O\�}���.E��"B�݂+'����&�(=����'>2u�����,]B�K������$v����'9k%�ǐM���O�%Z��y�v�y�&���O~���<=��8j�O��D�O^��|�	�� QΊ��f]!5
�!I�M�>?:�s��!^S<�Z�����c>U+�G׉#����K�F�ʂe�3;�	!�/o�p��&�ٶ<
|���ċ�d��T�i�*��I��'�h�C�(l�!bb`%K�ag�i5xʓ  (��	�?����6�`�B��� �P��F	�U�\���':�YR�	~�D��V#�T��-b(OXDz�O��_�Щ�,G�>]dO m	xĺVk�K.�jG�������	�?u�����'ht���@��!e
��'�<m� !{��F�?�(Q�Y�K>�x�媞/�����=ʓ(}���S��	��J>s�ޕR�n�EO&�p�~\
�HӴ��-�r$��хW�S���[��	+�~��!K�ßph��)A��s�;K����P�e�@���Fy�`)�8$���(dmR�_g�I'�4��4��c�]J�W?���E��zS/H�� ;�@Y#�̤�I韀sg���I�|�aA�#Aڜ�
�b��$�b'J �	k8�����G3���Mސ?�������Bd�}��_�]'4���*�N�8����֔L� ��A�ʭJGѠ.��XP2}�	����'��2�ŀ�D�jY���Hٰ�ZM>Q���0=����Y��y� �A>:�a�D�c���Y��L����g.
s�b�	4�w�����\y��m2\7M�O"�d�|r$-S��?1Q��2�
3�]�0%Y�E�?!��8C����^�B�h��+�^�;`�2z�Pϟj��7�T7jdz�8r ѳ5���Ś���2�͹PK}�P.['���J-&�U�G����6c�U÷E��p��[�����K6$2kx��uF�D;�^x��ޣH0��Иi��M�"O���V�^��V��Ђ��T�j�����h��5A�$@�#: ��W�I�_�v8�B/{Ӟ�d�O2��5H%L�BQD�O����O�Doލ�Ƈ��5�$�H���
)�"��GC!z(ƕ*`NH�JU�1��	Z�b>�%���7���0>&��ԊɼgF@}9Ȁ�oW��x�a��v�Z0cEc���b>�nڳK@�� <���dč�W�l3�D�m�� ?�V��(������?yc� (Z�*��תz-�P�	�4�y�\�P��+R�B�%� ��$��;���.�HO�I�O�����a>Id8l��X%WY Sh&b�����?!��?1±�&���O��4|�R�q@�U >/D� ���x�����(	�ꆝᲧ�uN���צ�� �0�!�� ���T(�3O�"8���F1z��y���nꞸS&��i���h`�
�j6��.g�։���I?`Q�P:C��RE'B�O���O⟈F��ǈ�@���;�� ��P��U��y�">})�$E��
��9�����u�f�'y�U�P�s�4�?���f�pp�A�?�����._I�2���?��ꝸ�?����4��[�:	�d̎=i.
�33G���- �k>b��5�q�ݬNଗ�r��кF�2�H+�������;��A�&�* ,ե|���\'m ��E\0����ڝ��'e�@���^]�'���i��W#��M��O�!j��	�'�z����/W(� I� �~� ���A��E�|�R���L�F{�ȓ�������i�r�'�Ӣu�Δ���Tf�V�0��
�,�1D����ן��ֱp����a �T�yauLO/0tQC��q��Z0'�(�kTnO*�Pp�$�o�ɊbA�Y�cD"mJ0P����i�1H�5 �7i�}�g��X��ࣩʣ&�l	�'��I���/J�&AaӼ��$�'4�8���jش��E{���6�p��	cyR�'��)�=9a$�7_�\1H�	q�V-C�e�w�m+�M;J>����YX8�@%�`n��`D�.0�0����?��hԵ�d�ߪ�?���?��=��n��0�J���j�D 3�&��uF�	S��f��o�C��34jX��1�I�{�z)2'���:v���I����D�$�S>I#�ի#��'�X��N(�S����L���C��_�'�z �u@� e�|�����$V!TR��'Sb�'�2EU,S�p��� D�d�var�'��X�l��^�g��.4B����A�9��$;%	]�?w剸�M�#�i��'>��O��ɇz������-��e�b,�)Έ���­/�L�������ܟ,�֟����|�q.ϛK��=��%�7ʸ�ڔ MW������8N|�$p`��1~	:�Y&
�K�У<����^�Ld�!�"�Ԕ���P������,�^})qk�"0�!#F�ӷ^��<�U� U��Q@��>,�2p�?���I���?10h�9H�qk7LS��8�+�m�L�<yt�K�>���� úȒD��OI�	�M�N>��/�L���ǟX�Dd�#v0q�6� *�`y��BPޟh�	0TF�1���ḑ
Խ"�"����CDT~6���lۙ{���ǀ݃k�d�����OH�Q�f`�,9`��^:�ze�	�O�䃤&S(`�1�"Q�@�?9��ڟ(�I^~�d�QHm���
{rzU;`�U���?ӓ<�2�Ha�x�h�r���<����<y��T>=2��+�����怃6�����;#�M��zyBIO����'��T>MQs֟��a�jx�H�"l��Z��ӟ���w���vNٻF)���G�Y�da&!	�X��O�LA�#ݐs��j=�R���O�� �
� %r%����<���iϋd�2 H?j �D�<a��oZ�^��G+&?���_����J>E���Y�h-R`�b%Md["*⍊��yB�.B���I�)��c1@5H�h���O��E�� 5^�VM0n�
`��m� ���?���?�`Ft���O��?Q��?����yG��.$L�5)O<��b�F��B��r�ď.nt@EC�!
*>�����G2o\H�S���Q��	'
�`
��2�9�LU�(Y�%I�������CVx�'3���ᅻ�t: -�AG����ˬ��h����c�	�����8�3�/A'���!��|���z�ʅ(p0C�I�)�`:e�ޢܨP4&D�O�˓t���SU�h�6i{�	�Rh�C,�W&�IQ·6?. ���?Y���?Q�������O��S�(�F���i�5,/nqa�B�b-"q) "�8[��F ��p{��\�5A�)ʆ�6[���1�̞	U�+l���K�6x���	��	�P��&C\�6�>Պ���(O&�h��!�v�Ya ֹ_9F��c��=Ou�-wӚ�Fz��>U�\@Ӓm˶@4"C�J'�B�	1�ʀ�)�~%ݨgF�(���O� o�ԟ�'���)��~J��@ ���0���Kٗ`����?Q����?�����g�a�4�aM]%�TB� j���`�ޭ>7��A��\���e��|>eGyr^+
XJ��"��(0&c7��G�2����Ɯ#&:��D4Xu��"2�tDyroK�?�ûiR6ʓ[��|Y��27b��� �t|&����Z������.\�[�.�1����N�4��W�=<�©O8E�ᧄ�O��F����?	���I�	LG���֐�M{�J�@�5� 1�I���f�R܅�� b��.��ʧ��>M�R&M�L� L�;2��--~а�F� d�q��̺_��I���IJ̧bt��G���ut����͒X��'��p���Q����~�J��#§S^2�bUD"c|؅��5Q�]'���Iy�i�'�<h�6��.0��CQ�H	4ض����ߦ��ش��dꘉ1!N���EqB�D�`(	����?Y���?��ۊm�*�Q���?���?��'�$���ㅂ�@l(��C�4�d��\0X�	�-w6I����m�3�	�E�b�PB/A�������E�H�M wJ��J۴SV�,	��k�g�S�? ������)d"V�H�-N�;��5�z�"E�'t�������̟�'�H\+d!�/Hi�@l�� �ɕ�J�̃eh֩G����u�?o�Z�N�<�A�is�7m �4�h���<��lO^e�<X��LP�e�~��8 �F���?���?i�V%�N�O`��q>Q�����Ow�(J"f0`шq��B����40l��u*��oZ��C�O�xWQ�D�4"Ϙe�B�C���%N��3c�G�J��Q��=THЈ������W��R��M�?Y`*�:x�N��W�X�=�O���Oz�d4ړ�O�hK����!��aB�'�]!�-��"OR�A%h��r	��Z���"��|fe�&�d�<�4��8+����0��j�:5+p��N��(�ᦎ����I%CD����h�'B��!)�Bď}�8��"���Ms��ɲC��x:a^+5t���+B�B,K�/|�'�\r��S�SXT��FQ1u��hK
J�d[SÄ,T�0�g�ў�h��n�-5�⟰�Š�O���"?�	�d�5�g$�V�^� f�G��w���횕A��5�u$�3b��J�N"�O�m�ɱF��m��W�/\z�{��p��ľ<9U����V�'��X>1(��Pş�K!�@��\z�+�z~��1�@�֟H��!E�P)���zk(|��D��t�:RU��N2��OҦUꆅ?E.����@�4���O������gE�)x�b�+��L�Jw�� h�|�fkX17b��I7l��iv�K~R�<�?I�i��#}�O[ ��c�Js�L3���4e��'	TX0g�*(X�MAɛ�^���$Cj�Oa@x�%J�.�. ���3~�^�+�i�r�'���ҹ@���0�'U2�'�>��`���M��vy<I�( �R�\��D�ֹ=Zx� T�×3�1��|!���~�k_�6e����?;�>��D'��Y�&���� �`�#�S�Ht����h^�r�X�X�S�፹4X��3�J81��-��41���HT��d����g�;�腥�%��qI`�):a��0�R4�`)�	N�ҡzOӽ�X��'��"=ͧ�?-OL�)S�\�~�� �oU��8}s	{f��"�@�O.��OP�������?��Oc2)`�m���L bRa֞q�X��@���w����ʀ�y�m�uΈ73�V��ĭ�v�'����P�{���SΝ�Sʒ sb��5�l�$����jd�B�ɧ���-�q��p2�lR��̺w^�i���#�ǟ��	�&��JE+��	���7MַK���ȓ{,N�� !*$n(��ՉWs81%����$��x�̓�����O�H�B�2�V�"Vc^�;}@%��d�O���Q� 8���Ov��#8��ᚁ�ѡ+9�� �"Ɏ;S�����f�
|�6	�5�L񐰊�<?X�u剈g���:5�Q%��1��I�FX�p��N,5�����T��<�6(p-���剫8 d��I�1�(Oyh�A��j�>4��sJ(���|��'��Y�C��b���P
͠3�����usB��Co�ɰA�
�2��Bf���?�.O*�d�٦��I��O��Z��'�t���bI3>��!�O� 8䙱�'N¢��/T�*��L�	��8�iN���O9��^�d9�f4W6�0J�̓�PZ��BƦ��v�מ��\"2MWۦu�ǻ�j�3u�~�d��T�>�
�9p�Jթ�i~Rj��?	�i���L�d��z�Ӵ�T��n9��iӽC��Ol�$5LO|=��+������W�!�����hO��$�}B�	Q�[!��c���]��H7�J�#�7�O����O���A�U�Z�d�O$���O��݇f�X���[9`���RCĮf�i�k��	�)�ŌT�B�\c�<�S}�I,)����X>�je���D�x��\��.=Vj*Yb���(��t��+'�b�Q�d<2��ϣZP �S�D??� J���ɟ��?�a�U%1�!�P�~�P0M5�yBT
b�eVA�zK�#�.���z���D�'���.�.�C�`֛55Dm�ŖU�nX󇣐�dc|��	П8����IYwn��'n�Ֆ{ �7/�;����FŸ'Ve+�n	n�8��ӷ~?�D�q#<�G\�c��E2���95I�E�8aW�20����h�!�����O��cp
�?^�.U�M��MPv�j7�&�r�' r��"�'4�����d��i�KT��7��ȓT
,��th�5��j�hR7~%|�%���4�?A+O$eCG��T���'��P�IC{����m(��c�'����3	���'F�)�!���� 2��Lb���;��1�O�\s'.�	Sb�e,��mw��I��Y�#�𘣎��p��Ǜ$:h���c �=$�QD��O�!��'��L�2ϔ��M[��Q��$�#>�D�O���D̍t�v�"�Fęw��A�7A�Y��ҧ�O�+%�Y:Vx�iI5�RZP	��'��57�]Hش�?i�����:l���Q�o�*� ĵ�������^~����O`�J�z�褢��X�JM9�'�n���?�'A_, LE�c	K�etdD�F�>?D�܍Z��t����d��ʱ��Ow��ӗO�#h����$�>R���O�d�w�'��S˟�� ���íCSL�S�$W'&�`�"OB�
���c��X��S�l�rq0��	��h�l�h�C�6}�l�[%����@��f�d���O4���0:4�͓l�Op�D�O���yޙp��6OP�qw%�Jj��#Ԅ��%̴�)��C$B<�g�źu+�c>�%� ��r�>8e��zp���
5C���h�Hg�@���AG���b>5&�X	��^�4>4S!��t�^P3���Q�I�v�R��.�3�I.�F|�D�<�Fh��o�B�ɏ ܽ�4Ð��2��P�^4ʓ<����@�I��vy��_�vp���k1��-Hcj��!��1����<��Ɵh�Zw�r�'o�iE2N���H��X�';���h^�P6H(�g-H�'lapq%L��p= ā)��9h�
M��@|H�'E<
�	�#.��2�����(\O脋�GE5.���8�b)���xNҍbӢ�o�i��d�� �H`���La�%�b���o=����'��O��˲`I�i%�,��J g>(X �|'p�~��<���V��V�?�ӡ�ęH�M�򂇠xz� �n?O@�� �	�DX~����F�\�4t�V��?����DURP�(��n� k�����3�ՠs+O
H��'�1O��T��+���JI���% �"Oz�ٶ���eX����	? �D�� �'߄�D�sɰ���h��8�^Uۦ	Y7#�'Vx�Q��'����O�'�B6a�D�� �jӖ3VMٓ�0�?A��g��p���
?*!�&��C���ɚ��@���/��H�`�H	44��I�'q�-��Fx ����Q�O*���2�Q�eT��4 R9��`��OĤ���'@���<����7�� �7��89��hb-E�<q��Ͷ-�:|{H�6;P��H OH�F���=Q�0$���L�3m�L@fe"�?�"眭���B_���D�����O�Q����3�u�5�
9�:���j�S�(|A`�'�bq�Pk�1��Ϙ'%���@7w�����9.E�1�Ϋl�����'��\�p'_<��Ϙ'SF!2�X3u�v��V�� 6�����DΑA��'Gў���0Vc )p%�[/�l��fd\�<y�<Q$�Z¦G)�0�P)�Xy�6�S�tS�$���6C��3��$��a���AƘ�j�'H͚=z���.|�Č��w�H0��4FKHB�c�������Ç*�8(*XE��<i��;���$(I�(�$�O��H68k=�wJ��S�(��d��X���$A"��JF��U�
H�%*�/v�k��I*A8v;E@E���"F��8a�X��ĕNQ>=��A�6��P��7xZ����I�x?t��O�b>���� 7@Kj�)t �8�ʙ{�k�<9	�2&� +P�S��$3Ѱ�8$�V���F{*����'�l�@��[�0��ϛ�z�*B)O�b���-`��Οt�O�*A9E�Oi��+|� �@'�^���IQNU�R���@*XX��I��6��U)��@��Id��i�1��遖�K�-��C����	v:O6TcS��3*V���*R�Z9H�f�52YxMӈ�4�bDP�펶]�����a$�y2dE.�?�Q�i��S�W��`��C�<�3�S�G^����y�K�n�)�m8�0���jݖ�hO(E��M�;d�2�
H[�z�|�yw�J�E���'�R�+b�љ��O��'�r�w���I�Xe�8�\�$P�p��+ҭ
��1���S�"]��J ��a�jVn���Ǎ:U�ŦO� ��D�mhz4 WB��U���X�o �Ay��z8�*ǌO���S1���鶈YFy�!�!�\�S[�|px�ԃ剸m�����Ϧ�����y�'�<{6�˔��.T$��չ��
�'����ԉL��X#P���2��T�����d�'9�m�a�Q�<T3G=E�E�s�K�_g�u�c�ގG��'���yݩ��ҟ��'▉u)�/⺑���2L�(�#��T��!�!lS�80�	pg�P@���3�H�օ��j��s� ��e"K�}�:i�5�:fu��"GȚjJ��i�|*����'�2�J�!��P�b�H&0�L�3tA�^���i(#=I����L��<3�k�-b�80�2M,	�!��B/H�<��6E8I���x��]7��	��Ms���d�=c�x��O�:�bM���[�cz��^��R��'��uR6�'���'���
���<u�FJp,�N��e�֏Z/J�eX��'qfR�q��@Ȧ$�U����(Ohe�C�<a	�y;#m�P�l�s6 ,h%an�6T�e`�nF9�<+P��	A��h+!�OjMo����'i���V�`���c�"K��@�'>a~��V�Mդ�Yc��LѠH�"��>�$]��r�3aZF*'�R��׆�<��[�6�'��Z>������	���09FF�neR� ��D�2�N��	�K���� 3z�`J�� 8:�J��`��Z
���|ZЩ�%f���$KA�"��� ���<ᄋ_�y�T��$<L$ss�T��a�׍L��aŀ�9Ae�
-}������^�<��W�,�	/�Mc�[���N�g�? >Թ���!-��%�̰jA�b`"O���b	�m`�d�!��#1$X҇��%�ȟ.�[V��5��9ƣϘc�
����OD�$�O��9&-�>\����Oh�D�O��O*���&HA�����N 1|&��":M&�AnߵN�\��Lp$��'Y��|��""}V�t��H26"�|ɰb	��hq��J7��t�[7�4Yc�+�րW�&��'��9�0�ؗ0߮њF���Z��SX�`�FK�O�`mZO�L>q�'>b��Q�7؁J�S2���'���2KȚ)��ea��P�S�@����_L���ԟx�'a"MeḐ?2>���FR�Q��Y�5�]�4gDD�#�'D��'�2ml���	՟ �'^�:�b�K�_�\(�O���iSd,MfE�6Ϳh��Ó.�w�$h� =ʓf8��	�r-���ʝ1�:pk5�҄a�KԠ >``���^hT!kdM�Q����O��`FגW�|���580`(�����K��D<�.c�ԓr�. �H��B�g�6����'P159j����̌"VI�	uylx�d��<�A���h��ԟ�ϧz��B����m���%�V��!�ɥB�t]��ϟ0�	2�c'OS�^.Hlf��b�.a Ba�8ƪrƄ�0��q#��9wL��k�j'�Ť�;�I�|���A�C8X�CpLK�#�>�XG �-p��:�bӎ�|�.�Q����O�%m���o�r4�##	;Z?:��I�}���'�a~�W�U�}G&I�5�8�E玬��>�X�L�A�5~Ո-��+�0n\�Y�b�<)���?�����Ĺ|z��y���P�l�e��<A$���T.���p����nyr�>�}r�o]#!������/dt����ZE���MCI<I��7�U�y����#S-Q����%�h�o�ƟXJ�%��<I���ҟp���?5���<�o9t��)�Wi5he�#��i�޴�?A"�F��?Q�'�"0���M����i{�Q�1�?�fe��Ǟ�N	��Ь�K��'r�`�0O���(���?	�I��?�qN
�R���"1#�o��X��E�����d�֡O͟Y��S�����]�F�ԁ�r��w-�KDPt2`n�1����>}o�'�x3N�~���?a���?��t�2��ݘQ��`eɠo��IƮ�?!��4Q�؉������4o��aЉܒ
�&�V��|��x��C��)���O�Y��'��"��	���x���	埤��~"��Yb��8��8q��$d� Y�� �<�1�J��I��u��'_��*sA��	g��(�b���;3�@a3j�s���H��N�*�D��j��Yg*�Ob���	=��ȟ��	.�K�4}��23��@\���ݴe��\Ù'aڙ�S�i��7��n�d؟h���?=�d��M�&���Q�.��s	���(G	A��M���'.�v���R7���?=�O��D���4\D�S��h�Z���l�5#��B�	��Eʥ�^�V��d�`% �v6��O��d�O��$�O,���O��d�Oh���la�p��!PV.���l��K�<�i��'�"�'`����	쟔�Ɉ�4<��EɈ j�\�6'��]ti�ڴ�?!H>i��?�H>!�O���2u�\�!�K�y1��ڴ�?���?a��~A�SU�Ԛ>y�ʝ(X�f�SU� � �H�ٴ��O}�'�	i�'���D�[�`l�U�\��S��Z/�'���'c�'�r[���'.��\ʐʗ,;��I7Ü�CR�p�'���'��I՟`�O��'`m�Q�1FD	�P�Q��9a:���
��`����$���P+I��х�R�P �8:��`���G�A�>]�ȓ
��(�薖d".P tm�-�")�ȓh�, �7`u�Y���� �$���YGFx�u�C�O�@y�C��;d�N��?A��-� dYeL�$�V=�!��U�0�9Bm�[Z��J��h�3u�W ;\�4$���uF�W�G� �X"G$��P�.s��Q��Dye����<� i'n�xV- ���'z�] ψ: �3�'*����vA�0�(A　3T;��I�o�V���keG��D�܈#�˜^䞑�e)�v;�]"vlǤzWn8�v�Uf똹��u�,�aB�D#r�y��%,dMh�/U֎�#K:�M!�<�>U ��T(cF�%�f�Tڍ���Ŧ�u�i'���� ��P슕��Z(���O�➘D��H[$=N��!��ި}����@���y�b��'�� �&C�$� HV�yr�J�	� �9$O�q�Re��A;�y2��dN���G��p� m��DB��yb������X̃�i�&���Z�y2Cڬ�*E4���a���f���y��Ed�� qBՍZ�z��e��y��P�]z���!�@N �J��ylN!Z�2 i��P����ƪ���yr�C))�01�N�`�v� ȟ�y2�C6�b��ۿP��ݰ�f���y2d�)o^�(@F
H%�1R����y
� �����#Y�$2U(S\�0�"O8���,i�H��W$�\<{0"OthQ��?/	�x��菕g��A�E"O4a��PTƲ�1hψNޡR�"OR��6�I'/���a������!V"O؀�a
�b%���ΕU�0�"Ol|IuJ�(�,p���^�6����"O:I: �J�z#V�"/T�GIp<z�"O�92Aͻ�J��#�ߍ1/ʰ*�"O�屆N�	�09���d��!&"Oj�� 
��S�b��EΓ)Op(��"O����N1&��d�����6�%"O�4;&��	�r2�R�_�P|BP"O���R���)h��)��E�_�%2"O���=.sx���ڂ�j��"O.I4����(B&@j���"O����0Mb�0g��~����"Ox� �B��9^z�N�(�&1XA"O�d�腅:蕓r��>Q�� �"O�[�e�d4�0㍁i��Ţ�"O��`mR�x���B_�O�^�HR"Ol��c�?��ð��.�h�p�"O|}r���iGFq��![�?2"Ot|i��Ubn����e�6"O��J�ǽH�+J�	7���h���G�<�dKQ1����н�j4 3C^N�<�7B�,��u���^�<kZT�ΒI�<Y\M���r�j�&�����!�D�2B.\:è$$w�h{�"Z�!�I��� �c�F�3^$5Q��3"J!򄜜���{��� U��E� �%5!��_0 ��ɗ�r����ՈX I�!�q*�ҦR
p���`@H:c�!��*_&d�@�6{RI���$�!�]?<��X�7j˯Tp bw�uKd"O���'��= ,��-SiҀ�"OHd��)2)XXYX׋J�yX�5AF"OLA�&F���3�
�in��"O<i�EAQ�4π�3�'��1.�pG"O�iP��:F
@,3��"@�:�S�"O�dxc�J���P��V�-�����"O�Q�f͛�E9�����!��;e"O�9�v"�*5[n9Z�̆;ctջ"OL Ҕ���]L}�%��Z!�v"O�"�N�P-�q���&��)�"Oj��h�u�E(�D�:� ���"O�8!��v۶p�C��x�V��"Ot����0Jl+En��
��9A�"O�+�d
-Tp�۶L�T��q�6"O���vlN�*Y�bi]�Rn����"O�1�G�!0 <�BNނ!Ro!�$ʚ���2���*N%�ࢵ�B%A!�$]�6W4Hv"]�����2nY�8=!��G��X�$ �$H9"[�o�w !�M�[T99E�(j�� 5/�c�!�3'(�#+G%@8.��vh��!�!����w�E�c)���d��0�'��a��� |���1�H-i傤a�'�j�Ó#�o4�)�Xa���'���K�c��\Sb0���N*!~����'56�Uӝ8^F0(��ƶb� uJ�'圑r�g�UF����n]�'��p�����̐'�ٝU�P���'���RjY�x{Ll`��V�v�x��� �<�V�����X�n�*B�F��a"OL�S��
*J�A"� �N��	W"O~$�E��9@�ɁD�	#)����"O6�(2&�R�A��in*(��"O*�Ѐ#�7ʨ`{f���^(�t"O>M�@���Q���c���E� ��"O���t��
k����$%�M�"O�ቑ���%��FA6�%��"O�`+TD�"� :5m_,^�(d��"O�Ũ�۔Yl����M+��I�Q"O�5ч�
�KE�)����	g��HR�"Od�i��~��f��:�:غ"Oe��(I+u�
�jcd��� A""O	Ha�]�YJ�dp2)W1,�b�kC"O�8B��.�|5@ F�]u|�+�"OR��%�>7��t��%��M�~�"O�ek�u)6<�A��*.WleQ�"O�� �9��P	Q��|H"�+p"O��4c��p���q�o�K)�t�"O*m�sO�>r�hy�֬#7Af�z5"OΨ�u�g> 03�K�$Iv9�!"O�:g�.��P��I� mAL��"Oҝ@@��V�M��)��8�X��c"O� "�N�2��U��nW�X����"Ojt:�<Yh��3"�6�� F"O�P`�ȋ�&C���􏚠A�H��v"O�D����PDʅPH-4zHٹ�"Od�E@��g����F���F��W"O�|q�j��L[uFȱ�"O,��R��]Qp�WK]�xUn�"�"O�<���ۤ#!ҵ;v��S1���"O8|�G�)k�,�#`�Ƥ/��PR"O,�±��P(l8A�,ZI�"OH�� e�69�!��� &��#"O��Q����Y+b���-����"O +�,V>��qCx�r��"O6U� )�5.� _�*Ժ��"O��Dʡ͘�)�#�1g]�5�#"O�"�@�>�m�tl�Xy�a�"O�ɺ"��m���!��1m %z�"O�upOW6�%c� j�\�d"O�a�5�\>M�.�q���/���aF"O��`�'QS!�����ͥ(��U9%"O,�����O�N�(�_"Q&�|�R"O���RB.B�^�J�X<\�Z�"Oܡ���J������9&,�yx�"On=i�J��({�	�)*8ب��"O��0�
"ojLK�%\>��L��"O�t�Ä?�<(i��y|Zh�"O��2�P$�6bcBJ(e�4{u"O�a��֙jt��� õ3V��·"O��s@I\�]0LUqR)�ym,u"O �Q�C	k(����(� L�!"O�e��덙A>N� 슊G.Ѳq"O���W ��D���Y�W\R1�"O�`9%�	%�xCl����"O��ۃ�P�b��I�AS� =��C"O �dT�Y�]Z�@ *����q"O�5�B�%#�>����&I��Z�"O\c3HUO�j�9FoW�(����A"O6�`W�X~r�mTN, �6�1"OJLCRGA��}٣끁0���q"O֩��,��'��L"��
f�^q�P"OH���+��H�phං� D�ɓT"O� ����X5[r%��K��'��Q"OZ��։�7>؎��0�Q4���(�"O�L+3�� x�� &�K
P ���"O��_G1��aiQ/'s��Z "O��(��ÆV%j�(�O
��h�"O��2�I+b]����L4"�d�R�"O���B��	��x�/C�cް2"O��h�E
#	D��(O�u�R�i�"O�ѓf)g�i���)8܆�I`"O�������3�	(1��@�"O���H�7>�� �׊T&���"Ox�q�\6&�niB��� yH��"O w�>zb�=1�*
�w��y'"Otl�$�B�Pz�����PC�)��"O�Q�e��)9U��A��V�M3�$r�"O܅H$-Z�Dx�H�"8��x�"O4��g��5K���1���F���"O����D��TD�'�Y�"O$u{2�ݘ"���d�����!"O�m�1�O����*��=#U"O>S�H�4�&m8���(�tp��"Oj-���1y�z�h$�[�����`"Od�p��{��d���8=�|m)�"O�8�5���s�P�8��$0X�$;�"O\�[3(N)�ղq���*�8�a"O��p��U�|�*�kB:ٖ��"O��"l�3��(CD*��͐Q"O�
&dHh���㇪�+l��Y�4"O�MZAH�=-o�3
Y�����"O���ͣix �CJ��\��!2"OxPsϖ(��YȆ���X;���"OnYku&��j:l����L�S�Ɠ���8��Ѭ~b�DGĆ%J ��ȓ�l8� �>^'6��Gŋx�P�ȓ)�(��q�' ��{ck�=�����E�k3�Y+(�����$!l���ȓ��!�R��R����
O� �R4�������ވp�Z�h�E�
EX������$�C�P�H��6#�*;Xڵ�ȓE P�A�K�|�DX�k��u�ȓl1�r3+In���I�M�.X����ȓ`@�d�Uk
Nj�Y!�W��R��ȓ8�x��&��$U&�A�EJ�M���q� �QVEU�>m)Ө�;�<5�ȓg��1���Hz�4�&���d`��}�z����c�]R��
�Lx���ȓy^lI���C n�8�F�ŵc�)�ȓK�� �-xVv��D��O�.��o� Ȅ_^BxJ0��3�ZH��i����!� K�`J��8h��ȓ&�n��f�y�ݰխ�[nX���K?�	f�W=;8e���V&�rU�ȓ鴔P�̈Vlk<2���ȓx�n�P�ɒ�V�$�{TH9M����ZL$���U(�I�0����]���Hx�c��+�h$���H�OG01��l�JA���0~�p�"d��L;X1�=0�Q�=�a�V�/v� �OA��>OX�r�&�5FV�]la߮x��C�	�N���E�f��D+!�ݒE�!��]5�չwj؂d�0�0��ս;�!�$:��;��
,V�㲪��!�$nH���A�9V�I�ʅ o�!��иg�U��H�'���邧Mw�!�d��zn���#W��J��&&�K�!�� ,�:3�\+���&�1"�����"O:�8Um�
8t��oY(6����"O(U �<��c���c|�p�"O@� 1�4=�d��n�"~�0��w"Oҽ@G��#�:<b��\�?�fp�"O=7$�.����0c�P�򵁷"OX9���/i��y�K�^�<�y"Op�;�#�J�f�5k��dʺ�$"ON��,E�2Vx���c�S�br`"O��#���+�s'!�3N����"O�AطA�}u^�*�E	7S)�!�"O��� x0ũ�<�Ҡ� "O��I�ᕻX�ڽR�)C>��|е"O M��a�bo�R�*P>x-�h�"O�x�	!�� �@)�'z~+G"O$E�6'���~���!Q$6X����*O��x�l��+���0��B�]>�'���,�JP�� �S̶�1�'��SЋ~�Xe��;{>������:M� ���G�����)o�<YV.�=b
n���%i2�}` &BO�<Y��J�<4�P�A�+�z!ck�N�<q#����D�`s�##��y��O(cp�W��V��i�'L�VIC䉵U{�y��[����Z�D 0�BB�I�:Ҷ�Ё�@��$����^C�If�qJ��iZBHE�+Z��B�	6;����Pu�t��3�C�I�i�\�T�|
�e�QDA�dLC�I�'<��J�M�>V.@ͣ�eO�^�8C�Iz�@�2Pg�pR�[���3 C�I�*�4���$P�5Q ��2t��C�I�d��<�cD��LbD�q��Kv�B�	�z�����m:�H��`�B�I5�d���睜b���2iC�	<����='���%.׵4�C��>8- �e���0��P�3h��B�I+
�)� � ����2C�	24>(q�3�T*{̸l�쁊�B�I�(��q���nS�l�d�3Z��B��=� M W@M�o����*"ڒB�S�CRnK7�Դa��%$��C�I�5� t)qi�(�^�8 �)4��C��C��M٥!�g��6
,=�|B�I�Bǔ�+1@P�9#B`�C�B/m�`B�h�l,�`�O!?��X ,ՎXpdC��HAr�����C�R���:b�$C�I
���eK�(O�� PwJ�Ir�C��4V>Q���':��sӎ��0�C�	�I��J#!�-O{*���k[�C�	�4Q��M�`TQr�7��C�IJyu8Ua�5K6,�1U�Vt�C�I�g���ʷ
������%H�,C�IK�PqI1I���A&[�l/C�I.tq����n�4wa~H0v�Ǭ��B�Wa�<��dȑ3xD��RH�|�B�	%���q�I�5�� �l�?��C�I�3Ŧ@�Ү����)}�C�	�C�������GC��3c��d6B�I'Q��� VN͡Ay����.�MEbC�ɰ&�j��QkZv��2�VR��B�	�f����ώ[ȬA:b%���B��j�:|zs!ʺ7�ɰR�R&6�|C�'n)|��ѫ�{]�@1�o�+Z�B�)� ��Jk �^K�<A"Dѫ�t���"OA�d۴x�����-#u떔@!"O�i@q��1Fx�y�F�0�< qV"O@r�(
�?@򭻒��N�JlJ@"O*����[鄽G��	�ԠrW"O�i��"	�(,��Z�5�D :2"O����(/2I�u�ȼxj�!X�"Oxi�&�� ������	DA8P"OT�i1��d�b@���HF"O�y��̂b����O�~��¶"O���e�Z�n+��bO�W�Ra�f"O�g䉒S>}���r�i�Q"O��������K�Ά���h�t"O$%�C�~�4YӬK	j���B"OV����0E�����C��*l[�"O���T�R1Z}u�� W�޼Y�"O,t2 vo�(G��j7z�*�"O��h��Q�a�@CK-���"O�H�)����FB�n$��)0"O�EQ�A?���P�ؚF�,偵"Odhb�@��r%:4�T�n�����"O(�i�jʭ#��HFdJS����"O��s�%ƕ^~%�I	c�`�*�"Oh��B��&9�6�Z�ϔ��<I "O�%����8QKɢ0-G�Y�8h)�"OB��LU3}�$�L#V��c"OX��f�Գ*'*,�P�P�p�"O\嚅IX�Ү���GF�k��G"O�8���7H�n\���&nƐ��"O�-k�F�7Fap���G����"OP(`��k�I01�*��4j�"Ox}3�!
	0!(��N��@�"O �0@+i�b�`c.F�gU`P*F"O �U��[+�`�A��@e �[�"O���"W9��:g�ؗ+`����"O��Q�(��l�ڼ����"O^t�u@F ���@�2q���)a"O�JC� �|��-���ٖ��pX�"On�q�"�(Ĉ�$��9}`�Ö"OJ��A��"�`YX
�V�
H��"Ol����
��P��Rz�$m�q"Otx�d^�d�S&ӗ+����"O���a�ɀ/b@!�kR0[��ݺ�"O�i�/� �hF�߳� �:3"O�X����{]���&eb͔��"O���Gƃb�e����>j��"O�0H�(,���P�
N ��"O$HR�h��$d�oωdJ-;Q"O��k�A�*b:�1 N�^Xu�"O.��I��zF�(�ˀhܱ�C"O0d8�z-��"'D�(s|���"O�	��� C��D�����8c>=A�"Ord����3�,Ҥ�]���F"O�h���p,݃B��[S�t��"OX	`fAn��Y���<sMD53#"O��لh�!!"��:�nG�F_n�ð"O�����Q�r�(;��T�n_ĝʰ"O��4K�,?��m`T�/ND<-�"O�=@!_8n���LP�z�i_�<!q�Z+YN&T��Ae�L<;$�Z�<q�9b�T�S �]dـ]����Q�<A��^s�D��%&�$D��4��A�<�3e�6�j�H�"!.�X�JF�[�<Y�ND�f��XT��>lz��jw(UP�<� pl��B)I���@���-�.m�'"ORe��`Ė(Ϡ��R$۪;��d"OF��
��N�Zuk'䌐:nh3p"O�=�'	�.h����G��
d �"O����Ьn���[G�^��ѩT"O��(���b�B1�H( �@�1�"O$���  �c?"�x�B�%��"Ova7�
�e�D�ժ�K<Q34"O���FՅ�dB+�9�@"O���fP�Li� �w�1b#"Ot8hB��+A�%z� øGP^�ZV"O\Uh��X�4�$��g��6�*(#�"O��b5k�D}N����`���Pc"O��!sAB�`VB��3��&�"O���a��yX|@#!'+�e��"O���&�M�:[΅H���u�|c%"O�me� #�m����7e�bx�""O����k�5d-n���e�;���AC"O���Ѧ�=m�f��Ĝ�?��@��"O��aE�Ayh�Ӣ*�a��Hxp"OhT���`>2�)���	�:q��"O*�JA�\�u3v��xʠDb"O>�C�$',ֺhk�;&�2'"O��1� �K��	���T�>��"O���֮�1K����� �!���v"O~�{'L8qf���� �z� �"O��#��0yR��Ul�1!z�A%"O�գ!�ī5�$� a�=	 d��#"O`�	�(r��m��՗<��d�a"OD��LI�aQ�@���2�"O�U[�IC��:w��(F�(��"O2p�g��{ˬ��$(Cx7��JR"O(��I��{V2}[u�3FJ��S"Oj�����)�S���0%'�q�1"OĤ�f�=�@ '̈́z#�]��"O�Y����,���B�Y�y6I+�"O2�
JM'�"T{���G����"O�Lj��R`�Qag�
(.l`�&"O�uh��Y�n7�0���ͤ5�w"O�QU����Z� ��E.�);�"O��S�E�,K�ڀ��JT�*10t#"O���֭ZX��b��_�x)@�yA"O0�a�L�F!��Y�ş��f���"O\�m�1�@��u.F�`J�x��"O8�AŊ/6�%�C`H�h��y:�"O0pZ6�ϽQ�H9��H�L��(�"ON��B�4j�*!����{�؉��"O=�ćܞI�:ᓷ��$V�=��"O
����RJ}��P' l��@�"O���gW�P�<��P�Ē��I""O| ����>~��X#e�F��RQ�u"OіiQ.Θ8VJU9�LL�D"O��b�K6Q��)�T�Ȇ~`�6"O�Y` d8x��*ؖwi���g"O��R+E�O��������X�0"O�d���ÚD���Y�"�1\=ܭ��"O�ȱ	�G��ⴁ��}�^��R"O����$"?�ミ�F%g"OKE�(G����	DwZ�$��.�y��٭KEtd
�	'޸A�� 0�y�ʑ+c���al��>z �+4G�ȸ'�^���u�ܹ�aC�|��I>9�ǿS��c���J$��q�<y
��-���̙�^�8 ��Œo�<A�L��� ��(�;R���:��c�<� ����kȤ%��AANO�#�`\9�"O4����#��5Q5I��:@�S"Oa�� �<H�$f_Y��x�"OP$�ᅟצ}E��(�l�Ц"O����1&~ݐ5L�f���[C"Oƹ;�3��0�7w�X��f"O�E9�I�C89�p���8�X�`"Oh��W
�"SPp�{�"�[A���v"Oz�����>(\�阆�Ü8(��A"ON���
��I����kʷI	�a"�"O��	��B8,�XYI`�46�(w"O���B�aU�$أ@:\��Y�"O���J�5v�bp _7uܦL;Q"O����B0)|`����Q�b]١"O��7�Syj"T`AL��_Wb8��"O�P�fX��.Y���n70+f"O8�E�׻as��YV�G0p��7H$D�h��i�`� pn
&l����w	$D��)��)f���!jSx��p�Gl D����o��܀1�P,f�)4�;D������j�Vը�`�4������7D�:q���T-�l����&H�l"bi6D�H���İV4�!�M����6D��AT�7K��ٸ�$�P���h�!)D��0�c�i��Q�9
R|��	(D�<�O��b���IRÍ�r�qfg+D�@˦�V�V��
L�}�J0��)?D�$�&g�>�P"4'JJ�x�)s�"D���GjD�v��F������3D������-lo\�8�	�|`"Lsq�7D���(��p u �=�8���4D���R��#H#mz��	7}v�*UA3D�8	��N�|����t`��l�DF&D�@��ǜ�\��y�c��RqhX�S� D�l;S���y�@9Qp�]�SA&�D!D����4�^Db�3P=�E�;D�h8g`�5ג}����	zq�i3��5D���R �&N�8�e�B>8�ڌڔ�)D�H�u邍R�٘��eҼ�W%$D�SlAR��M꒯��7e��c- D��)��2@�����|)�(�#�#D�����Q�k3>�&�ȉ1Dxi���$D��{����b�!r�Y�UFy��d!D����cךT��)@���2Pg�IJ��,D�Љg,Q2&���s�
/&�3�)D�<1�a�2-f�ش��,|ًBi&D��{wh��Mľ���`ǝF��'E9D�� �$=���Q��G �a� �,D�X�K�K�n�r�6��Պ2�&D�83��ǛPd�# -��UƐ塦�)D�x��(�7J΢i
�;�%)`�(D��1Am��&4�yE
ķ)�P���G&D�x�g 
#����S���,_��� D��eF�pC�@c�:tO���s�<D�t�u�I��Z捃#?X����G=D�@+�#���|#G�2�l �'D�,�"2$�Btr�C�&mA��2D�dDG� K� 3��@?X¥��/T��I&�����Ok�|#�"O0x	dχ�EӲ BΊ�s��zG"O����	t���2b�?	��x�"O��Pl��#��'	+Q�Ԁ$"O�q�](-9���W�|e��ϞGK!��P�+�m��G������B,!�� 2�bԠ�v��ӡ�I����"O[Q�GO`�ɢ+�D% �r#"O��*�"�I�ni�U�<���q�"Ov� A
?g�|�*tς�x�yC�"O�`�ɂy�e	��]�@Ӯ���"O�Xʇ�>8���T�ϑ<r�D��"O,y@$��y����E�H��8���"O���e�?	f�0�/c{���6"O8��&��+"a��� }l-:e"O�IS��@	���ʭK�n���"O��*� [�7Np���^���96"O�)r`)(�vܠ!	ϧ8غy�"Od�9PF��
���D�9�d��"O�q0���W�|����,x̐"@"O���F�"=�]*F�� j˞-�w"O��n�@��{�6��M0s"O����Δ̨P"�A�8B����"OazD�ce8|��� ,�� �4"O��8��gҎ��!���q"O@��p
Q�S^9ᆎ�s�@��"Opx3�ނ%~V8�1��N��}�F"O�4���� 3�ѭw���V,�f�<9���W�h=K���d������k�<Q���W���s*�����k�<Iu&�����4͊P0�XC�Gd�<��]��7gp���NGb�<Q'�K���p� �J�f���OR�<1A�7@"I�"��(Q��O�M�<��E��ޔ��
P:�LIA�f�s�<���1 ��I�.��LT��!�x�<Q6 ]��f��FF>6�����Z�<�v(�i�"y0�:`�RPp�<gQ��db��S�a��a��Ep�<)7a�`�u!���Dd	�@k�<a���;~l�BB�	�$D�]�c��o�<���A+fH+�w���W��n�<�%l'@+��@�G��n�	9�n�<���R�)L �Ɓ�>O6$1B�Qi�<��+N\ڜ[�<}�jɘ�o�b�<�0	 7@�\r��	�n�|رDNx�<y�JN}�<} E�^�,���kw �N�<!���y���;TȵKk��ñ,E`�<9/���l�ge�*���p�c�<���3Rs*��5��%8�Az!�Z�<A�J�cQ����+J�Y���IF �W�<�Q�=�<��a钴����W��R�<��eD�r���Q�N�ĵ��^R�<��Ə>���0�,�zss%�P�<y�h�	xJ`���ŀ�(�
�z�aN�<id!4#a��	��_��P(;��b�<��NW��6��a���L�t F�<YVƔ|���c��=2H�J"o�D�<�ԅ �Vh�P	R.Β\z�S���H�<��$ɞu�H0�6�ڋW�X�DQl�<!g�֗N��xZQ,^�b��z�	�O�<�@N��רU1�0C�-AP�<���\c�6�k�V�jl�
ф�f�<�G�ԋ���!�R�1�:� �_�<�,��x�x��aH%P��^�<ё� �J`i�i���X�.�X�<��%ޕICJ��&���B D����I�<AD%�c�2qU�/=5X�AZD�<i��$
�Az6��%Pyl���H�<i�-1�,T�H�D���)`ΏK�<� VmK2�G`^�e W �6Rr�x�"O�Ȁ��F�V�R�쇒Q����"O�˖�ѱ.=���p?�}��"O�p�D#ؖ�J'@ �.>*9��"O��@A �u�R��`h@�o�|�i�"O\�q1�X�I�2y�3�2q"L�c�"OV�K��]:C����A�:/�Bg"O�ݣ#艫,�Ht��漁�"Oڑc3Z�<j�� ��; ��Y�5"O�`�Ťp��h Ȕ#��1�"OЍ�cL��~����E6Jֺmӧ"O6(	Mŏt(�Qm�r�"|�<O�����]͆t�i���~����$�C�ɲe	Z�*D"E�3���K &�yY\C�	cxHYp�ߗ4�$���D�<C�I�	���&�� ��{���=�RB�I9�ZmKաJ*��l#q�
�4��B�		w�����с,�"��Ԋ�J$�B��2 #d��Q;$���˖+<!`�B䉻���()tb��VMϝ/��C�I�U�<��~	N�
��>�nC�	�%�P��Gۇ+� Y f��IuC�� (�rU)�a�,q�9�#�Ps�B䉘�FUz�*Z�:1زmY�TB䉄t������2y��7�8B�I�kX"���Uy��h0�ZB�ɞ%��p�1�A#7��pP�Y�:��C�	(7�v�#�G�K�H�i��|�C�	:u���� (�w؉�30,�C�I�_��,�(Y�m���@N'�C�	>V�ɰ���U�����6�rC�	����!��� \d8��Ť*8C�I�a����P����2XIς"�"C�	7)<TD��oX	j����QI��W#C�	-^v6��c�
?�mAT�I�:2C�	;�V�Æ֪5���ƏE�T�,C�I	(p��� V7�hӌ�+f�B�,"q�u�7-�f/�¶ҫ �B�3B���A_�p_�)�c��=t^B�	9��I���3�s���RB�	E9�8���2P���ňB�,B��|��ᱢ�R�Ӻؠ�G�Y�@C��>e@]#�+�9-�P��&A�+UC��
�^t����D� ����m�B�I�Jh���rOV�R�@f#�*K5|B�	�de���Bs@���ʇ��>B�:.�$MS1�S->V�!	EB�/��25�Ñ `8 l��C�I�%���BVHŊj�^U"�I0~!�DM�#)z�d�ўT9���oJ!�	'}dP��B,c�Y���D4`A!�$��{tD@rM6E�Ȓӆ��<]!�d��.fL�C�a-�Y�GF��aH!�䗭}R6 K�g߮"
���K!=�!�t�ᓬK#Ej��[�\;%	�XQ�'�q����X�X���5%�pIJ�'��L�E�Q�~
D����U!��-Q
�'j��@A�T9��d�6L�n-��)
�'�����C�`	W�m���	�'�x�yAa�8hR"E�s�f�0�J	�'��D�+>�Nj�CٟW����'a0|QV�Z�zd$YS�=Nf�[�'�|�� GϾw��%c��ItJ��	�'왈����#��q��I�t*�ģ��� ��@@��Z.��H��V;�M(E"O`�"Ќ�++�Fyɓ�N2��ض"OB�YaV�$8(�󴊐�\���V"O@]�����+�sgK
�aF��u"O�-Y��d%
^���"O��#�@N�9�����IX��p�"O $�T��<=��� c�&~��@g"O"���ş(�P�Y7K��y?�) d"O�i�BƇiҪ(K�[5H-��"O�	�fH$:�h�*JTs�Xx8�"O�JՋ��Xǲ� `S�"�E��"Ojm��.�N�L)	�3E���2"O�9���:H/d\��
�k�[2"O�x{GI&J}hR�jQ\�`["O`<�*D�8���JF{H�\H�"O4����۹�M�S
�X�F��"O��H�!�#߸E��R
��(�a"OVAq� è��5�{�X!�"OV|K��1�$I���R�o��j"O�u@'/��qX�����T�,�v"O�Dx�C���L�T�1H���P"OL�K��]2< �����z��I�"O>�r '	�p�
�r� �j�1��"O�mG�a�:l��iOҕ�"OF��RW1N��0���O�1�"O^���)�x@� �?Y�b�k�"O�i�`� �R�T�з'���� �"OH=������B�VgU�cx�y��"O�*3�SL*�x�D���hu�p;�"O ��������Ȥ.V�:s�9�"O�q8g�$e�|�֎W"��7"OT ����l־)R�����E�c"O�8K֋�9o����Ш�2!~d]B�"O�t� Rs�nM�Ɠ.|{<��"O�# �ͣC��Ȱ��*~�e��"O���N�|$&@   � 4��"Ov�pcN�W�p�.Ƽ&�pp�q"O�m�Q�݁?��L���v�L�s�"O"ia�/)+Vx{r��q�r�s�"O�,�㕩O R����
ˌ��7"O��b$뙪^�$�Ҕ.�&Ā���"O���5�/������0i���g"O�0�#Е1 ��-��Kت �"Od�3��%�J�k��٬g��e��'�}d�[���q7���?Ѣ��'h����B?9��e`D�O@��y�'�:�������zI[QI�:Q:��
�'o��z�斄/	��Ǌ1�
y��'�Y!�/Y`�᳦�S�Lp��'z��!`�Ͼ�����
�U)���'?�@q�d�/)�d�"�_:Q�Ę�'�� ԈKA @�NV
b�A��'�j�	P�/J������S�X���'*U�7`�:��Y�+E�C
$���'q�	�!͟?E�eB�I���q��'�,<zs�C�����Ěy�;�'����6h�)x9X�3!�\.G�����'��:�fD>��Pj	�<DN]	�'T����d\�h0*�a�,/O�h��'k�� s��6���Cr�D*$N���'(�`�7 �����"��$8u��'�ИZ�˛_����"Ј�	�'L��H�?|�����E�K	�'����J#z)r�V"j�v���� t���[�
R) ��HH�<I�"O�a)�J˕0T0Q�#�ՙj�6��"O�e����+1�<@#�LP���"O���$ :W���Q�7G��|��"O4�`F��M�����/�^�2"O�T�d�)�������V�8��"O���� ��7gDd��J+~|����"O���$�'�v�J�*ʻ@X�XqU"O����'P��!�<���p�"O��T�]?&��R�̵>�b-�v"ON%yP�)%*��E+){X����"Ol��AF X�(cGjQ,HH��q"O��!n�4�l9��k�*�Hk�"O�4�ď��1.$͉`�?0H�u"OV�35���\�H��F�>|�(4"O��"��
�U������/>�\��r"O�\�"�Z�l��l�2@� ���Ic"OR���@�d'��p��_%�\1�7"O��q) 7&�^��K")��e��"O�)��
�k��=��شi�v��"O��zOh�0�S�$.�� ˁ"O�	k�J���1m��P��J!"O��q��<Br��W����c1"Ov��@��1H��7��!��<p$"O؜;&�C�t�Jh��_#H�`""O  (�c����i �T8։��"O@����T<5�zQ�`MϾ )B�$"O
=Uc-f��q�ɘ<�
�R�"O��pF�O�
O���AIP�>�=@w"O��0�m�}�>�#��xf��r"O8�������Z1�5r�0d"On���JS�5���2��Z~9���"O�1�3ǈ'��@M�9(NR���"O��U��h��!&�E:4]�"O��V`܏oT�< p�\�*�=�"Od����db��e��9g2��R"O��p��y%�I�q��+
d��"O<��� +^�.M;bEũ���"O�p��C(`��
 _]�00�<D����C�(0
$�Ǹ"���1n9D���� ����$J��h!��7D�K4�C�y�������D�x}� 7D��#�A�����9tH�x�$�F�/D��Ӳ!�����2B��c�r8Y��,D��B��߉� A�KX�+�D�q�,D��x�l
�&��U�Ƥ�{�L��**D�h�Gn@�h�ȫ��|[��6�'D��D�Z|�0���%^�V�a:T�'D�,I���1&�`����(� �1�&D��B�\�tiD8�ƉY������8D��T&\�]�A���T�l���v�0D�H�T���J�za��Ʊ|�E��*O��*��`~�]�q��?q�Ҡ�"Ot�C��F�j���Ĉ�1�ځ��"O�dp��S�c��Q�"�A�Z!0�.*D�L�B��dU��B��G}p��4D����i�~���)P� ���I'D�$z��T�Y�P%/�)�N8D��@�z R��`hI����re�6D�4`v*S�ZY6xc�g�,m\�3Ƥ3T��نBX�Ei���7��+oF��&"O����`ӌ� ����$`�1��"ORE�nU#���DgK�Q�8��"O�l�F[�M�,AaE�#��<�w"O� P3�"�T�NX���&	.�� "ONx#r��i-��p N��-�P�R6"OB	3u�97s���$MR�l;T"O<H��E�b�ґi,zԊ��&"Oh]���$^�<���*X4J�h���"On�ږn�4Lh~A���A x�^��"O�)@Å��j�D@�$U��	�"ON݀P`�.L����:+̄�x "O����J����#�L,|1"O��2W=!��P(ѯx#�,�2"O�da��Ǫr$��h�� Fq����"O�����8��R�$Ynh�%"O��ɥ~�{fgõRP�"T��3�y�9%��Hx `G�ڹ�r���yR�M`b��ށG���T��yr���oZv���b��Q/zŢ��y�#��7�Z!I��B�d�)�ߊ�yb���_��P�� )~�<C�@R�y"H��.�Ω�m�W���P���y ME$XAd�ã| 2��s���y�R��qU�U�n(v�qf���y��X!�q���Z(�0��2�y��*W��,���_��(k��B��yb��$u]��/׬V��P��㙮�ybJ�qb�r�G��^���9����yrf"�hi����Y�LLI&H��y�IJO:�9�ѭگQ��$�%'��yr�c��ɪ�9C��k���y�$���b'�6��2��>�y�O��c7��P��^�-`��@o���y��Ӱ?���)�[�aÅƆ�y2ˢ#ܤ���
�}W:erTK��y2cW1���y�
W)��,t�_.�yH�T���+Iu
D@���'�y�ώ(h�`��n�+s��R)R%�y҇ØEN�pRN[�*�-�A��5�PyBB�T�\�p�C]��|��B�Z�<�@Ӝ ���JEၳX�
�KU�@�<i&��wtX�2p��m`tٱ�i
W�<�g �qG"`�M�']Sҵ��@OR�<��&�D��宝�K	����L�<���V�^a���[FDD�L�<�90I�}�`f*-{|=�"�G�<��l�N�*��c _n:�b�VA�<	d]�$�n�c�׍e�ʑ�6`Z}�<�E�A�yz:v�bdΊD����"O�8���"��"L�R����"O;ƭ� c4䗴&����+�3�Py�!ć(ta(��T�!�݁ÍS�<�#��j���Bb�S��pUv̙I�<�f�'�.(bO*D� X9�%�D�<�-Y�?����G#�;CϞ��3_B�<a$�H�Aѵ)�M|��H�Ít�<�-�W����D��HggL�<I�����]C�jλX]r���H�<	����,/���!͒W�$L��L�<QRd<�*,���[f��)(�a_@�<!�Kά��h��A��I$>�k�g]{�<	����Dy%��W8�P#�O�<���ҧk�~�q��ջ"U�:˅"Or����U�gL��e+�"3����$"O� Z��O��N]��=N��IS�"O�����ְ<�#��)B^�ᣤ"O��8�/��^��Ѓ�P�DDa�"O� v��g��._� p4�P9fe�&"O�Av��6l�A!9M��=J7"Oz%��
G�WĖ��s*
-���"O����l����$�Ԥ�@��"O
�aG���d�Z�S�����	��I�h�"
,����'���R?�0RMB4W��A�-O�O��m��_
Ye�p���?���f�8!�@H$a��7�1���zQ�Z��4h�+��y�|�[��ИU�:L�EY��(O�R'-[��DI"7��]P��ʹ(V���R�~��K񀖨>��cd�C�"h��ǥ��'�M���y����<���Bղ DZ,{:�Dr��&\��3.T�4�?���?�����wW­Iƅ]�^F1;'CU�)Vy��*^�6f��7�8��!��1(���h%F�D�F�am�̟��IT���5:+��'��!V�`������Oay�2iX1@�p5�~N,��W᝷�N�����W��/r���?���+���:�g�7K �J''3�8lehH��D<e������ʉ79����2gpb>�X�����`bE8eNE�G!v�:6MP�z�Co�d`ȩO���s���i%N�;P��q������O��D#��۟��>��̩^���X�&�7E�|�u��L�'��6m�ۦ	�ɚ�MK����Zw�ܤ�êwX, ��C�4܄԰`��O�$��c�N@8��Ov���Ob�d@ߺ{���MːJ�d�V�HBm1+��Dq8�J�E�S	#�$� /A#�BȀ�O��-91k*��6�Q�f+�=�~!���	��|��L=R߾�2��Ց 	pA�I�����^�P�%�ڳ���z�,y��(C�2�����-�>�V���4��4c���|�'��ei�eY!o�
����Y	de�{]�8�����SR�u3�iU�U���#�T�x�>��ݴ`����'о6��O����ʧUv�0S�J�4+i����eԮ��0��B[!,Ŷ}����?���?���4�?A���?-(j����߬:�Ks�L��bZ�ʇ.C��`*֤$���.ֿUʠls�b�d�'h�����ڬ��0Â��}���a�5��	���ґO0l�T��Gu�yP��:|S�OUZ��'�`��F�}�	U�NO��؉rY�P��6��O^˓�?Q�*��9)�e$�F�R�� )_n,�L�TH<�WL"�`�G(��<~���Xh?�ǇD�"���_��k�N�<:���O*�&�9i��_��� I&E�6�h���
��'q)}�a!���%,��V�>��i҇\i���$^<D�1�픞-�L���޶f-�G��2% ��P��a{���
Kb����-+*��w�W�}t���:��N�h���Ϧ-�ٴ�?���J�������R��$rN�Pr��՟L�?���w�M���]9�~��N& �yP	�E��V�aӆ7mO�"a�7-�5���YֈІv!��u���m۟l��_�DΊ0(h��')��	�KZ=���*EL��{� ��\�r �&؛QM,|{Ǧ&cB��u�|c�����|
�'�5Fk��+b�YZ�A��C�n�Ln��$J�0��[�@>� �+�I��� ��#Fr!'?ט�j���g�_���#6�H�?�<6-M�6d�a�������i��`rM<i~L=��i�1�V��'���'Y�}�b
�&x�քHG��1'�*����DŦQ�ش�䓧j^wM8�:�I��ܹ���O,0���@�D;��)lO����  �      O  �  �  #   f&  �'   Ĵ���	����Zv�������@Q60"���5O�ȑC"J�+^��$E�/�*�˔ɐ�d`BdƄYy�\���S�\��Y8���5OR0�`�0��i���1{����&��a7��ZF"�C۪f��|0�I^v��8U��$[*�݊&��)���jV�Ia��RdAޠr検�cJ3> <i#n
5S��-�fbJ�2� (c\ ��"=E�x�K�J�T8�e�	D�YTL�>C��P"��?O
��$=B�0��n_�|h���O�(|����aX�؂!c�#n+�D��˘[��hpRe-D����S�Tip����G����KЮ,D���5F��,�Xi�B�"Q6���5?D��jץW%��DhMO�{g\)S��8D���H+D��d�N�]�H�Є�&D� �r.� Hl t��N�1;uF:D�H�gݽ��J� @�Q
�	��<D��Q0H�</�yRDN����&I6D��顄E*5�Э�C�ٔy�ҭpw�.D�p�S���p����%�����x�#)D�\��"Q��"d��Nڹ$12�p�)(D��@WD�E�H[��)eX�a��!D�|0��U�Z�)��˻K�<M�P#D��xu��&�x�3��W�Y,�X�o!D��Ac��?o��䢧J!^`!%D���v��=b^�!�6 5-���#�e"D�H{�V�^A����mM����c5D��)�L�0v�&�9g �,�z��r�3D��!��LQ�t���@�;9v��f�<D�|���A�jiPR�V�`$@E<D�x���T�I���zS?v�dc�l9D�8���C/h0(�D��3'����#O&D� �� �$*?�Kf��{� ���%D��0�m�0A�X�І��H���R� %D����CB�B�K3lr�BH=D��A���&I�EF��n>LA���9D���`V[&� ��A�4M"q �K,D�T	3jL$6�jؠ��N�R��c�(D� ȥ䄴4�,�(�2M�p���!D���!��"G�Ը5'�;(�2��W;D���1/A�T���)����2X���;D���	S�/�@Q!�h����4�9D�@1w�ܵ|�N���*�����&D�ȡ4!I{ز[DǙ+A�>D��w'�X��0q��o.�:ա1D���VN]R�(�q�Z�=�����o0D��P�M�kBh9$d��P��1D�\��H�(p*�1�o��lY���6A0D�����H��8�B�aĕߔ�1�,D�\!��G/�܊t퇞?�][��+D��iU%^�4,Y�Ʉ?g���6D�`��DQ�xOj� �@�KT<d`aK*D�I�$�s���յ�`���1�"D�����Q�G��"�V�n���e"D���(��P�����d�x�a�*D�Ds5��!A�b];��@�qS���(D��#���y�M09�hx��B5D���TH]gs8�����"�v���1D�����V�Oz�����%sR�4�+D�,`�*[�q����$)�� ����q�.D��!"��`��P����i�d�q$+D�t�q���hR��f���2�*D�\µo̪4a���^�H�a%,D���u��U�^ͱPA��]�(��*?D�<�e�ץY��u�6J:��7�9D� 1Cg��:y�p7%�,?�NE�VE*D������"B�p��E�0�b1�� *D��� RQA0`{%�N�Je��ï6D�`��Ϫ� D ��ٱi`x	2&4D�� ����ȕQ�R� ���A|���"O�uɆ�I�/�:L���[�o�:��"O����B<_�4�s�w�����"O8��ևJ�wb�E�E�1��I�C"O
�z�-�8Y�B�FY�7���f"O���%J�tE@�
х�"�\|kr"OHA1�cö+�z���ꨪ�"O�\�ч �'��ՑѪE�?�M�R"O:a�g#Z?���'�c1�DX�"O
�+'��(@���r�f�<a�鐡"OP�&Iʎ8E��v%�2�}�#"O
����ȃ�$�bgC�E,��p�"O8x��'�+Pڠ��U�R
(|Დ"Ob� ��X*����d��Ҍ%jP"O(��&�1S�09�M�.j;�:"OL�{�@Ҝ��Β-t �"OfmY�*�!U��$(��<��Qf"O�-��l\/P5���� �hc�Q"O~0�"I�
xvLhc���}�`86"OL����$hw$cׄ�-tX�'"O�}˔$\���8.�\|�|�"OV��֦ ;/�p�A2I=~����"OH`1"K̜!o^�աÉ8k� �F"O����N֎y����6@V�OR0���"O.���mU�&\Ɣ �^m �Af"O�r�(Fj,�#0mSf��"O>�`�C5}�~�a@�Y�bX.D�$"OP=��i��>�0��MN�\Y��� "O�0Jѭ>r�1�@\��Lq
�"O�E�2� �s� z����J���"OةdB7�4�@u����n���"OT��J�2~%�ċAy���;c"O� Zd�Oq�0���M|�A�"O�|�C%�5 2�&/��L�6��2"O\!��n�c� ��׸�V`jc"O�;V���2VlR`�ȘL����"O� F��2Nz�j�D	9<`T�$"O�,�vg�8p�H@D�G��u"O��&�Ӻi�auʜ�y���C"Ol-�Q@О|^�CB	��.k�Mqg"O<q*���-��bc���4x��f"O��lC�A20�����kM:A
�"O2P�u��sNQ��PB%���U"O�E��=�>�!�LJ�l���ӂ"O�E�r]�Ԙ�B^4�X�c"O��в�ߖ9�0�*�/3�,�*�"O�Eٗ��v�QQ�m���	��"Op�)���q�����Ίy�"O����h�+ 픍��d�)����"OB�Ym� �*{r�-bє�q"O��ʵ��f<8i�+2�x�"O��b��\�A��IY�j�X%f�+S"O68��-٫fh�a��ț#Y���6"O$� 4�R�/��Q��7+�0�"O�qaצ�S��)�f�5#K�]�&"O25O�>r�	������"O�ݩ��V4t-st@H����a�"O䤒�J_�=ۺ�1کnp��Ц"O�=��×6�6�Id M8^��H�"Op�zK�,&��5��,?r	z"O����2r����T�VY���"Oxmz4�OUJE[d�Ę�&��"OڜZs+�	BN	hPD]�ά�"O`X0�ߍB�|��U�Q,h�ְ�'"O� ��&�
�_e� �"���.��[�"Oa�a.݅!"�<��iM�>�B|�p"OmBqBد6RH�C��*��h��"O(�"$�_3.�F���;}М)�"Op��9!4L�rMC45D����"O�{���(���Xuキ[ u�4"OꕱC^@��E�W)IH��"O>T���?x]�<���7^R�;"O���0��M��,0QH��9Fp@�"O�<��N�uy��RThD�J �(�	�'	Thз"a��` �3���'\ ��g�N��d��L�,&p���'L~���Ù/{�Fթ�߲\��9�'&��l�e:�@A��Y�Z�<��'�����I7DٞY��c�l;
�'#h,
��Ł@xʍ�5�`h����'���eEaJ�E��2�  ��'~�h�Y=
�
� 憓�Ƶ	�'�邆ޡv�<}�!��20�I�'x��@dp.��pn�x�
���'�4�[7� �-��p�
i�2<p�'��L9〗7ur�2�!E2��'	lz���~�4��H���'D��c�
�a��A��vP���'��9K�o����:��].�:�i�'ܶ�[&�mqL�(� P�!Z���'��ԊH�kJ@�sꋙ	'���'�v�	S+׳2�j���KF`k�'�(�+4,݇&�RD��ݡGNUk�'y���Ƶ%��`�,�Eh���	�'�x<	t�Y��)�@M zƩ�'a �c�	��<&\Ԃ����n!��j�'N�BP卨?0PuF�ɅgNF��'D�9��h-�xyQ*�a�֙��'��9��J$&�����my�'�!�O�t�
�p�IM��-C�'��-#h�ov�5"QbҞ
���
�'�V�۱"6̀� N.<�`�	�'�XMS� Q1x	�ȑE@�:6t< 	�'�p�!�w]b$ZЀX%+�Z��'ƺ�[EL[<D<�i2�V�n��H�'#���k��f���aVl�Ҭ��'�zTْ��_�\�	�i�
�y�'C�p��Ɋ0����_�3�����'Zdy�V֠7J�e9�M���C�'�6ha����ԁ�#�cg���'(�u�O����zC����(��'�8��Q �6��C��G���'��x%�O�Y�J-�s�Ⱥu�$a��'��H�k��+�I�L��:&��'�,M��-la��Z7�!72c�'#Bpp$�*f��y$�-�(-�'͘u��'������-���'���C4�E#L,�Ht��f���'��db�T&�.�������P�'<6��6F��A��< FC��`ݙ�'��Ç'F	j�|�1��uL���'�F�)�*�����a]Sd���'d��!J�+/�L��%�Y�b�#	�'��M��L��"��e#��2�>�S�'�\U�WnLI��8�J�R�	�'](X�C�L�I��"qL 7H����'v�DXw,߫��(��/2��9y�'�h �DGϾQ�����=,�i��� �q:3PH8�)'N	P!���"O.L)�
_/K|����ċ�S�b�8�"O�=��/��d�RI�w�\��@9��"Ov��������0E�༵�A"O�̘&$��@Q��Y�"���"O�]��ʣb�Ե��	E�"B5{�"OR �e[R,�!],��%��"O�|�g����c�ūZ��4E"O q� �X.K-C��[�g���!)
���I`X���'Ί�YQM]5/9UJ" 2D��K%I$z�����![	2c�D[T�<D���u�ٲ2��T�4&ڿ�*��?D�h
�枴5��*6 W�#�:Ѳ�i D�p ʍ�R^��� C�D�X"N)D�Tv�|lva�Em������'D����e��.�~m�c!� Q�d`��:D���w+%���j�R뎸��7D�Pe�\[Xݹ��@
^��5D�lbL��{�ؕy� ف��bQ,3D��Q���~��4$2FjR|�D�1D��5�Ht��ej���
3���R�.D�8��&��2=��Y�mR�X:��z�E(D��"�B;ڐ����ܪQ�^x���8D���6���Pж�	�JCtp�8D����Å0Ͱ��%�W�^�4dXS�4D�|p!���:*z4�"��)H���D4D��x��<Cl����>n#4���$2D�� .��,�v��@&�F{��+�-D�$J�+��^�c��TT��d�=D��� ���2�;�h�Eذ���7D�4�-��F�\(�DY�@��*D��*��U8]��ykFX
n$"$���-D��!%MQ��x�T3�US#-D��9�c��=��@���	��ɩ�	*D��2�G�~��2#�٣��Y��)D�xaC�[;��uy���
h���q��<D�8`cK{�^�
��^�k���21B<D��J�k�8W��`�kB�#_����H6D�T� bZ% ��C��;��*D�3D�
Ʌ�BOv��d��/xrmcJ.D���� K�;4E�b�V�
1R��QD+D� I"<�,u��T�"5>E���+D�Ĩ��Y�x�4�R�5'�)���+D�����Y��/Q����,+D�����3���S0n,�0��*D�$�g`Ϩ?������`�����=D�@B�kͭ�ҡ��!��r�<}���6D��J�ߟd_�Xx�gκ�(Š�$3D�Xb�?`�l�c���$O�����n2D�T!6�̸Y).L�`	��`Lu�6<D��'&�K�̥G��c���J��:D���"h}���-��Mz�SC#D�\��X�������,'m�A�M$D��d��I`0�u��T��Q��6D���%�W�+��9Z�e�0�%���!�D��K�:8"F�)c4mqW���
�!򄒇�4m�&)�4��
`��6�!�D6D��8�wQ-�rP���
�!�Dߚr`������.j� EQ'��C�!�$�7��l �l[8Ff�*ՀV�!�$��'�\��V�-U�V
u!�$ "ض�##I�'"Q`��j�!���+z��� �am< c��5D�!�I
je�� C�`j�L��g��}C!�� Jh0�i�i{��h��kq$��"OD�Q6��9���AA_:!Z�q!C"O��$Q��-�wfT�m�l])"O|D��$ڤ<*ҹbf��'��K"O���q�ם#���W�N��U5"O���F�xm�s�[�:ԭ�"O$A����MBpi��M�ڕ��"O�Hҳ��O�p-���G�@|t<(q"O�K�菸-<4�J�-� ����"OZ)c��ќ#.��1g�4{�DI�"O6�0��
uͩ���_V�$�1*O*�����Dxfy��̸��
�'���,��-��4��*�r�9
�'�l5k�+��]3j��g�˘b*z�I
�'76 ����,}�iI D��&9��
�'cj���	#?^,P�N^b�i�'���zpd�)Hp$C��"ZT	(�'����C�R>�����US� %@�'�%�CKEײ�B�պN�@��'��|3�`::�����?5��P�'�.���V�i�N�@W�1k���'��;&��0�@�Cg���#k�@�'�Ρ���2�ִ궀^�J>�Mi
�'��I��gB�h�2�c"�<�4�Z
�'�~]4�H�GxP�Po�#:V�P�'��cgdE�?��Zq�6'�
���'����G�uٰ`D
N:�0�'�(=a&k�^xd��gFLbjp�'n�ˑf^/C�f'2��y��''t8� ��l�tq$;q����'�nt��₁)Ǫ(h���$J
�'�f\����V���#�4(��R
�'ӈ�s��G6#���蒠��LK
�'��؀�LqWf�*��_6.?��C�'~% �eT�S�&����-@�P!�'���ZFjF�����d��2ڥ��'�0�O�$i�6A@�{�l0�'��h��J=wA���E̄lH���'���������t��(1�]��'Td�wB�,��C� Ƭ�'��-�b�3!��RUK�z�����'h��	�O��^R5K��z0��8	�'�fUQ�$L�CKR�H��C=<TP�'�~-�u��72����O����'Hl���%ۏ>>V�2�9X��e��'��+d�Iw7 m�%��_ќ	��'�������zu�`���B�Th���'���FY�(��y'!�j���'�6�H�B �&�s"7����'̖��V��3\��(��Ɣ-)
�''����c�$>���GO�W6,�	�'���`�M`v�zf	��I.`11	�' ��!ʗH`�Y��ݝ>��1��'���fN�%R1za:��S).֤�
�'� l��A�a�������.�R\�
�'|�餪\�D��c�T�n�*
�':$e�d��sز���'Gk�B	�'3n�� �I @9���͒=�Q��'�V�q�,W�,�~ؙd��T�-j�')&�I*�l�Ka�	<c�t��'Cd����Ty`ri���0v�>ć�=�>���_"#�Hp���+<N=��~0<�&1@��`΍8�䜇��n� �
T(a��h�_4/4Ň�S�? �a�w)��� ܠ�H����g"O��ӡԄm
���/����"OjhXg�r6}��☠)sJ�t"O$�9ԃ%x6�}����{Y���"O�1ֈ�,�|"���!4L�"�"O��Ҳ(N5�,<�l���s'"Of��mܯA.X�T)^�%�N�u"O��Q��rK�S���_�4�ђ"O�\;C��� ��Ҫ�N d�H"O-	�c,B��p����/�#g"O�d6�kY��Jԓ�搫�iZ�<QaW�<4B��6I.�y�ŕY�<�gaߋM��UXbnK0a�����T�<�uJ�%f��Y��h�.c=��k�<YWcȧv�F�tH�_I��@3lFO�<��
^�$�*|;Ť̬$I��hC��C�<�7	^�aɸ5��a1>U`f�W}�<���,�6̡��Zy��҉�D�<A���j 5��g+��sҮIC�<Y�/�W�6��āύI�B�+Bgj�<)!̀�q���P���h�VPCu���<1��M�yʹp"�\�U<f[SHd�<����	N4��"��3�8-�E�Z�<�DF��&GҰ�І�1}����(GY�<!	�	_��Bԅ
0�1���M�<�sM�Qʤ���X�hUc��J�<a`ܢ�iz��ۄD�7��m�<�,��q��J��A,pN�p��^�<Y�:!PYR$�� K�H��QZ�<I'&�
'��! e�Y�iR�`�<id�r���BP�^^x�#�B�q�<�⮑ O�`��n	!X���A�<Q#�G�Sk�����<K�:�{�t�<���Ͻe%�; a�;(��|�&@J�<q@W�)��Qr�S��J�F�<Qq�	� �� `��-J,"��@�<��bN�w%J#�l֬hX0lcF�Jw�<��M�.L�G�Ч�	#p/�s�<Ya7P�|��$�!n(��b�o y�<�Gm�)��5�I�Y��Uj�,�N�<�G+Tx\��X��S�k��e��`�<1A#��rEb��Nʄ
|�iZb�B�	&DDH{�bM"M:����X�B��8��=�7�3-�|k4n�lthB�I/��6�Q��<dr���qHB�	&#�`�S������⤟�imHB�����o��[�T9�l<qD6B�	�T%��҆Z<6M0��R'tpDC�ɣz{z��v�$}�p��1� $�PB�ɉa�ʅ�f��8q���Q���6FDB�/D��&┈gC����SWi.B�ɜ^��	@�?7|����R�g�B�I�tV�w.��wɨ��%�-v0B�I�0����Ë��T�^�3��"�bB�I.;�8�C�m�6XY�O@}�@B�	��2�c�fޚ7�t2qi�naB�ɻq��%�f�g�	b��Q�d��C䉢qJ���Ն�SpΜK�iL�!s�C�>=�\m� ]�늰b��^��hC�=_1�+0��
K�(C�kC䉏S���r�NN�x  q���5@C�	� ����'#�%�pл��`�,C�3d����3��رN�3HC䉹�ց�c��
j�`��F=C�)� N�BTH�D`��G%/�6���"O*H��c�6"$� �!��N��r"OСX.R�U�M��_VF��6"O�L�UɄ�]��� *ܰP�
�"O��D/W�!x�R鐣Hy�r"O�`����/ M���=c�@ 7"O��CRgS@���M�(&M�"O�y�/U1�z����Z.�Xe"O�5ڢA� N��6+�5��c"O��� ��L�VI������\�W"O�[0�ۋ�@
ȞL�\ɪ�"O<��#��c�IY5�H�0�Hd#�"O LI2�U�pohEjA�ȝO��� "O@��t�  �bᶔ���Q(�B��9,P�;�
�9W�ب:@�Yg��?�����Q��uI3(.d�$GF��!�d�+h�B��эb��z��F� ���
�(O�>�J�([Z�&i�#�#fH� ���5D�D'�P����P��"2ȵ���4}��)a{b&S���,�Ы
�Y��H�7�7��?�e&yӰ�	bL�+�<X9��	/T�8g"OR�@���4]W���Ȅ�p�(%[������>�9�a	��Zh�� �m��l��j)D��Hf��T-Q0�̢q�ڠ���'D��
�AW�MS���	�=�Θ��$D���VΆ ,�2�ѕ�C�m]P�ha�!D�#��Ɯh�~x�giM(�&$�F>D�([ԏ�#i�v\�����Q
�"Ac:D�@@�����B��w�فڤ)�W�%D��R�M�M9��I�/_�P���>D�(sʔ,_XI�A�uz�Hk��7D�P��I�?N �	���$G�!Jê'D�hX�&ܔ���{���	����'!D��ꋾ8������֬l�����J D�0u(��bF��EB#+)j��=D����kah|�W��0L�`��(D� ���=*�L����7N���0D�d#�Ԯ[��2�`�
�@$�0D���#�ɖG���bQ��qR� �,$D���'��q_��s��D(?>�s@�7D�`J�/�|94SG�#���I�n4D�p���"?T�(���V5VfI��3D�PJ��I�l���hK�tӄ0�ff'D�̰dd3��|�vO"HXl��$D�T"��E)@���r�/�2m���W�!D�C��6���١#(�Δ:f�4D��sDi�8c$�(x��3K��A`��4D�hI֞2մ�7��}!�B�)1D�@3T��#Y�`0�J>[�U13@.D�*�	�E#��Hq�]%A �	�W�-D���W)�z��}8��ٲ^G��h��(D��3J�?}����gFXC��i�� D�t��-C��U(��Ӣ	���*=D���ЌήFxpA�9F�1XQe�t�<�%�M�-$ ���\yfx�BAq�<QA�Q�""�[5	 �K ����+�o�<�7�Ȓq������|�zS'lOu�<yt�)8�5�S��>p�<A��s�<��	GK.8��� �C@��w�<�
�a~Z��.��� AA
r�<I�N�@�h��/zc,��完q�<	׉ޡs�Ȣ��Z� es�(Ig�<ٗOѣC�P(r�$�
̦��GE�~�<�cf�!t �QnJ!-��a@ȘU�<���C�XyzD
c�fQ ���#�S�<���B@������'��Y���W�<�ϙ*Z�8�B��:����X�<yD��&�Ƅ!\��� �D0dB䉙4ڊ�Ô�_�Q�����$u�C��{Ӟ��Y�����o�&hK�C䉸at�����L1�`�Wm�(��C�<��Dń��"윸��L��0�ZC�n^��c� �s�CaLWK7\B�ɻ`*����̃�m����U�8pPB�I�5�Z�#g�d7`�"��l�B�)� 
����åM�q�+Ӳ4D� ��*O�2o�c!vDJ^��<�	�'G��ږ(�&X�|����0��'_x�����gev�{���o$��'j�X���;=���GÆ�tL���$%s�`@3u��5�K��`���C}�5Q��O""e��s<e�ȓa�>��O�hLX�!�,�C�!�ȓ\h��R�
:�������9nDD��I�D�:̗�,[h�e"�"Zy^U��w��k�AG�t�����:M�C�I#}�BdR�hQ�]( S��_49�fB�-\�Ur�&B�'�(�0,ߛw�����#ci���R�i�)��<��.C2�9�PJc	Wj�* �i��Z�+��i6�Q�B�|i��&�b�2�)^�D�Ͽ���!t������~d���`����z�%�)J�h,҂�AFpb�:�/!pS(���\c�.�
d�KL'�ȐDe�%}����4Q��h����M�WX��I*���"��DM�UbQ�n�첒�� ��PX��# O
;"� �#����;����E~ӂ�O���`��P�%�>f���>>��Is��?�����ycMŚ�?a��?��36��OB6�G�?N�Y���	�2P� �M+�t+�e��w^p�ӂ�C?8^t����?�W���O��G�P�Wc<i��)��osDp��8I��u�w���(��xcb3��?��ġ�b��$@�2�
�E@�H�;Z�"���O����'��7��_�I�����[}��7\�6��!�D	b�؏��I~���O�^-:��?O_H�S�B�:z�=r�ݦ�ݴ�����'���k�h:��@�I�F�S*Ho2��H��G� ���O��!�.
��M��8pʌ��H�E�>@P G"��R�f��y�dP 7��1��<!'�:���c�D˄2��6Ϝ�Z�q����\���T^��H���k�\"=A֢Q�,#�LI��������)�%!p,ƐJp��1��$,�SC��b�ԡ(G�@����1N}F������}ʓ��l�P�4O/'�L�0�R?���i�:7ͥ<Y1�UDW��'�bQ?�#���a����ȭk���)Ufb�(@���?��Z-�HeK�	S|��Hťr�T��>!`}�SMzjN ڔfKN���N˯�Q��cs��M�K� H�'"�,ـ���3�|���.W�VT�jN�@~�h8C끱 �Q�h�O���V���Cׁ-H��J�I��um�L"p�Y0�?q�ʟ�b�P�G���6^MH�M�	`��B��"�O��m���M�ߴmW�8a�B�!_�tq�I�9|�bY��v�v9�t�i�2�'g�S�w3]����l�0��A)g��EJ�mrw'�ol�Q�SU�JY>���BZ�@ bi�%��RA��e�	������֘.e���C
r����e�X�N}66mݺ"�PA 	_%a�摚�o]��{0&�#�1�k���Y��H���T�b�F5�w
K(l�k��?�t�i}7M�O`#~n�_C I�T$ˮ)��1�B��W@��I���	֟��'���Iգ�5s@� C�4���K�9�Q��A۴C���|Bh�:U��ԉp��Q�hG�CP���.�>�@���П �5��'����	�\�	�`�Yw:��ij4< ���6�l)f���U�`�#�$�7� ؘ��o( ,��#Tj6��̔��Ԉe�|���(t����4*R�T�Y���6[#�5CGh�!MeT "5J��,���*����S@Ѳ��i,lb,ƬTǮقׅLFd<�'2b�r��w`�f�*���O\��>ѧ�W�TB�H�w�>A��)�נd�'ay"�&F!��� ���� |�CJ�:��0nځ�M[M>��'�rO>ݴA� � � @�?4   `  �  +   �*  �5  �<  C  KI  �O  �U  �\  �^   Ĵ���	����ZviJ���P��@_zX���4S���1A`N*G<��A,?�����ɐ2��b�ň\g6�I�b
)�6�ك'�hk��
�TVԸ����^��R 1Vp��H)�H�q���)N@�C���qB��1�`(�sc�# �X!�M=�B�#����?L�@���YY�-��B����QP�N��0�VcS�A8|�ypk��$2���	�u^��E@@���i؁����ir�(^D�$k�H�)1�0-�я
�`:Ƽ�G.&�f�$�O��d�O�Ь;�?�`���0��W�A��I�矷J����'?�59�4Y�,|�/�|Fy��R���0#i�lit��lC�L6^�Y���N�˖�
�q���-�Q�l�i@,!�VD�#���T,�<)���ПȰӓu쉃Ŏ��h�r#��Vl���'�P��@	=���֦�?!�n�mک�HO�) �$�v0 Q 1�A�
��d�*R%u�����Q)*���Oj���OV ���?���?��K�(&�̈������ŘR��8�ft{�NX�W�R��aj��)A(���ɪV�M{���3b:)�F�ǷO�`dCA�7\��4���2\�:����
,-qQ�p�E��O�,34D��v��Y��A�Dː�rե����۴�?9(O,� �IC�,GC���샪w�L�k�F؞x�	h�$�3t l��kF�F��d��P8-���$J�0�4��$T�;OU���?y����&�.���z�O�N����&Ι�M�GB��?���?��@�KK(�A��@�2"�A�i� f(�B��[#7�0MQ�$�,
\ў0`w�O=�)��l�:zs��@���r��<����"+NSB��.�T���	N`Q�8���Ob�d>�Ӛ`������)qQ�?����p?�3-b��u��H��A��NX��x�OFd�m��K!���%�P�4&PD�X�쒃n���MC���?�,��U�G�O���~�^� ��O�B.�X  N2�t�m�/;k\Up�DL�)+�ȃ`ڝ�b��O1�L@8�f�3]Bb[fdI�i���)p��O��r��[�u)Z���N҂Z��1��i�#~\LA(�8x���`@B�4���')��	ʟ��䧑�	=;b�:�IB!\o�͂����[ B�I�aH����/v\8;���5��#=!c�� s�H���مkoΡk���J��)ش�?��B�	#EN��?����?�����O�8B���l�up6� �gfzԛ��ȩ��ݺU'�c7ެeDʤI�b,�OMB�`"o�%l(L�qȕ����t�1�TX�F�& �P]�b�Dm�r�'"����'&�܄Ufl�s�O?\~EZ�����	��~��'�ў���awzy �ޱD���8@�2ĆQ��2�tz��^�NR��3�@,}K`]l)�HO���O�˓e����A����dQ%N`�m�k��b��r��?����?	R���d�O��<UTT¦lԵx=��zeO)^���pÎ&m��p��%�`��z�����鈄IW u<P8�k�:�:,a��S.O���3T��X�����O�XpCJ$gx����/{϶��G�ۦ���4��'�$#}n�X����U�O��#��N-Lv�C�ɥY��
� �ڥ"ިlr��,��dԦ��	my��ߓL����?!�OZ�4[ �
>R�ۡ��,1��U�޴$��l���?���"�j��E�>F� S$�FX?��V�xM��N&S"����
 7��F{"O�k�b%�m��~E��&>c�U��L�tlë�8\81ړG�@����M{���2����a	^L����ek�&���ʟh��E�4ˢG�w^.����96u����@T~�`�%u�P�8p!L����Ӫ��$.Ae �nП��	u��@�*M��'����G��#�Ze[g�V
r�����n�� ���X#[��cR��w��T>��|R��Urb��b*T��� r"*�?1�@�3Vξp �C�I��)�'rǠЪaGܥ>8�!�%T9C�M��u��	��MkS�����)��|���E`��$k��^�~%c�l>D��Qq��Q~�c��` `))cJ'ғ,��>Ql�gtp�"-V�T�����I;G�0c޴�?��R�I���?����?!��~���O^eIqŠ�xU�o�3b/�)�"�N�"7���J`�!+��8� ��OE\=�J�C�I`N���Ϯ[��U+��"@�$�7Eذ���U�����2�ʯ|BAmX J��O�|�D��(?�j��f(�n��&W�8����O�nZ'�HO�	�zW>���h�4c��;�a�r��B��) ,w-J�i
l4���*nm�6�����d�'X�	�-C�L ���1T[����f���f���GRۀX�Iӟ����T�Zw���'���s�`Ti���3�|���`]!OlA�����ȑ!H��\]��c�??�� ����r�)	ЎF)S���&.O-UHQr���SN7�F:y�8Ly1"��Z=����/r��F
#�	�cnAk
�F�/Cg6mHp�'PQ�P�����<�x1k��~�.T2�b*D���e��-itR�F@�L�d��o�>�T�imbX���ig�������'jW�zP*E�I��A���@�H�nڐb�P��I����	-t�F�P��Y��1����(	���V� 1b�Æ�t�L
�P�Gn�ܪ��=ʓr�4��B�G���k!�$u�f�� �80&
*�\-�(C�B).�1!X�'d�9�����1擽"�"��izR�↫B/3���p?Ig�G�n�x�F�"-r����vX�؂�Oh��i~!��lF�C[�D
POA��M[��?�+��<�c�OT��&Kr�@�ƨ�7^�)���ϿHC��n� ����ŏ,V�)��o̩m�$�ӫ]&[Y`t�|�P^�;J�i�� %^����)�?	B%�Q�L���.%G��ы���):U�, 5-�S�y��[�'�#Y�D��%K2;���>T|@�D��X.O�OK�?`�����d�Qh�,�E�,r��h�ȓ3ע@� L11ʮ�h"d ���Dz��8�'(Є�z��:P��5�4�:�XL�V�i��'C^��l3o���'�2����'��Yj���c�lhP.��-Ӟ���*��6��ɑUF������+���ʧt�02a/�D��Y�5�ĥX�if���fE�P
,��ã.ri�qq��^�fV>1P�CWU�'���1�Bɹ4\p�Ö)	k���/O�|���'|�7��'���x�� ⊜�$75�6��B�!��?]X����j�DaG����N4��|�����и�$py"�F����)����!s�رҊ�n�D�O��$�O``�;�?����#G0�?��$as�=>	��A���74�}�a�,�~rMǇ`� ���>k�� ;��
���>⤊ӟ\�!&�# �S�g�� ��S7�y�MV�L�1�M
b�N��j�#�y���.�ҐSCC�6[~��e����dC�m'����LE�M����?1�O��,	w@��S���i�K%"���9޴{��\����?���4�$���옧�,T<"����®�=}s��3�!@%�hO�jV�S2P:ʭ���Ԅ	9������=!�ϟ����	�>$i��)S�6���#-�!�䊚|:lȢ�̭i�@��	�=ta}��,?a��,>媱�E��(̨j��[}�F҅1�V7��O��D�|2AD0�?Q�S���b M�hԲ8�f��LS���$�i�0�Ww����b��I̺P�Ƿ~��$��f��T1�C�;�ؐ�F�=r�Q���n��nL��h"�āV��>QZ�
�~�i�e�$T#�t�C�Qԟ�� ��OF�$2?%?1��b?Ƀe�k|��K�lGzu�
S�<aT�.7��02CL�'a����H\W�'D#ʳKF��|��ufV�E��'_�8�bڴ�?����T
R��?I���?������OHH��j�/Q�j�@��͑_wpc3�|��D�F��U���v��.&�,�O`��h㊆�M\n]�`I�l����e�Ғ&��`z��gNd��N��pY��'�O�����u�����.ݤh$�0�b\�|�3��O2���Oh�L�'Ҍ�(%�ۥ4iୣ�(���e��k�\�1�65��ȋ -���:lZ��HO���O�ʓa�	h�=\Q�T��7:�X�FjK�d$t]���?����?������d�O���=w��8���@�9;AE�*F�i�PK�#&d�+T�$td�G
�m�'�HP醂'gߞ혣��YH� DL��J�t���ݖ�;bÚ�p���Ѝ�(OјE�'Ժ��&Up�)���X� 4�H�p�`����.�	z��M{A�-МXʄ,0bQh���l�@�<�tFs�f<��Y.V���6�B}�vӞ�Ī<�1o\<d��ݟ��'m�p����[$� (���?_v`n9�(`��ן��Ɋe�H-��-��ĸ��O&V(��O^�`	�2R;x�K�'ԐT��=0���ڞn���CEJ�t�<]4�%Gn��?X��0%ēӾ�hS�R���=����d��F�'Y�\�jZ(�z����1�ژ�'���'���C�kT��)#�Kܜ_z�y�
�F@�I;Z�HxR��:"��U� �D���*���1�i�r�'哧MKpy��������F�d��+\)&70�	����MC��֚�"�A
�"i[�t��i̧FZ��Wʗ�6�
���֒M�����_ʤ9k�hܘ3۶��mT93 ���	__j�ܡ5��{Y���6/�����Zu-"��(N��#�]%d��3�ʂXz訅ȓ�TȠ�+��@1�
�Zc�mEz�4�2�4����)ǂ���ض�,�10�i�"�'�A wd��?��'3R�'���ß֘93tM��	\`�0#"hU�(�(�ҥ�O�-�F`(2��(�d�|Fy����[�-U!{�5���,炩S�V����q���jj��)�Q�,y��T�#��l"/.r�ኦ<i�k��R	ӓQ%��P����cQt���(MyN�ԇ�Kklp���"�z� CI( ��ToZ��HO��<�ė�i,jtZ�M1N��2`[2N�|!���O�-��$�O���O��;�?�������R���z�cQ�^T�љaR�d���D�I&�!��C�D��LQ��-n�Fup%\�&����ȁU�U��E�~F}�)�|��Iƀ �-�"Iث
��[w�Iq����"ONt�F%��@�ҁʄ�H,u{���5"O�E1��.n�Z�Yp�P�g	�X��@�4��m��:��i b�'W�	E>@aV��}�e���P-&t�ƣ¶[��'��eƑJX*ԺD� �`���˔��O����q
�KQ�ҍ`@��%�r^ўd@3bS�uҌ̱�T�`��U�c�T8O��%�ϵ�,"oݾc�~�+�(Hx�'�v	���D�>ap��V��@���Q3�dy�I:D����D&� �!�5�r�r�9�O��'��q�@���k��a3�F�x�Y�O�4�5aOۦ��	ӟ��O=��A�'e£�w���Y394��R|\6��!,�%EK���뀍��
���Qg)Qjb>YcP`��jpEA �F�6ЂaO����!�3� �`��6.֤ej�F )j��8���1%j� �v��$:$����R��$� iT"�'��)�I }򡓗1�n]�d��51FH%�w��7�y�"�6���c��'���ꀼ�HO�G�����䑣�M�f�c3��)@��7M�O2���"t�%��h�O�D�O.�Lﺃ�G[���P�,a�ȨdQ/+Q�xʗ_����%>�O<MC	Ar�$��! ̠-E@��Q���C�*�O���"
|<�I��М{"^_��('��O�Ą�	@(� 1����!��@�mN�Z�B�'�-!U�C����*���f6[H���D�|�L!�)�c��M�1(Q�N�((r�
��=�r�'���'"�����	�|"�Nd�d��N�F���	�t���.ؙ@J���gn�+(ʦ��#j۔~�^�<i�n�w$��t��%��Z�a\0�R4Q��P1gt�9�M�4wq,��bI�!�֣<!Bl���(q�R�m�	�*E.W�j"�dq9�4Uّ��F}�E�"(@I�Gʃ?R�rГ���y2MI3EҘ���ـG,�e�׉X5��D�Ϧ	��Ry��8s��' bٟ\i�!��ZM��a5'A*^ߊ!А�i��4
��'���'
�S�j1˱�C�f�q��4��į�@���h#b˨\윹���V��hO u:ť\�$~T�2h_#]Zt=��բjA �i�K	6_
���)B�+��#�m�$����M+0�iC2ҟ�P)ᢜ�yh�� E
��7>��1�i��G?	�`�?,�P��@&db12&%�vX��۴%��ߺX���%��&,�V����|�~�~��80���.�?a����:����O
���ēr�<��b�
&���� O��@�h���������;��t0�ș���I1��54���j���ݙ)E� ����	)oǎ�H�k��XA�Ӓe4=��k/� �}g�M�r��4@��R�4�ݑ�+��?'+�T�K>E�Tڞ2ߤȳU(�Zb�P0��X,2!��@�� �amĚ� e�Q+H�_��� ���)P> ���	��� �Y�X���o�˟0�	�vȺ�alY��h��˟p�I3�ug��5�!�	T� ����v Ʊ�1����_�m�|"f��KoH���R�hK6u@�-C��)}U�|"������3L�_!޸��"D1���1db� LO���*�6�ԙ�A+�:��{e"O�9 �$��D`��jȏB�,As�i�h#=ͧ��gK��9���|�P`yd��&�~Hs�_��4����?y��?	����$�O��K��9� �$Lw���q돌J�. ��䞉oh4����S�.�"T�t�ϛhJ=�e�	�oj���Aމr�"�9�g�5%��Q�U�2|*��ZŲ�F���?!��`�>���������?�����ا�U��Gv��t%P�%�8�%�A��$�ȓv0��ᅻ5 X���UBP�'�"6�%�d��l:�Al�ɟ��	X�B|�`c*N�,d�%�Q���Y  '�������@7͈ ��3�ĝ\5�s�SzT`	�p/ؙ��Ε�7�R`�B\�'6��yA�уA�b�Z�m@�#�S;_%��R�h�31�Z���C�	$@Ң=q���ȟ���ɘ�H�z��vY,l�N��a�	a!�d.K��0���:n�a#R�a}2�9?��L�=�FP�	����y��Pt}�i�I��6��O~��|b��M.�?A��	�K�C:CQ�	IdE҅L_��KU�i��ٔ�G-1�`�bŀm��i���D�p�b��)�Z:�M�S��4�����_�������@����`��1`뇁`["M��]��O����֡J�OCVX�E�ݱ:������'����?��O�O`��Oj�;�D���`ay1-I�T�$�#$"O�5����g9��ы� �:E�u���O�`Dz�OV��� cq�N�;�l���ؒHoӲ�D�O@�ʤd )V���O|��O.Я��?y���W�`ف��`a�h�16���wI�&��|;p̌�Q���V>���k��x�'���1�/윊BP92��lSe�ɚ*�$(�Qa�-,!�)��+��)��b8M<��L� ��0���*���Jhy�`���?� ��� v��܄o5`Z����6��`"Oꍠ�$P,b��y8R@Θ+|�s׷iKl#=ͧ��.�>	Ѕ�4~�B��q�_�c� �#���su����?y��?	$������O��-ԉ�d�۠������V?��µ�B z�fibB�4[�z2d�)l�F�å�S&[���*���C�XL��i���F�@u���!��Od�����5�h�,�j�� ���Fʦ�Xٴ��',V"}nڔBB�y"吩t�zm��x�$B����X�B�:���*V(hV>�]a�V�'��� 2)��r��$�D�?9��nFz� 1 &Կ"@	
��dӲ���O��$�O\�	�
F�y�\�ca�@�IefCG�0�Zl@�"F��uX�Đ��|B�Q�sBQ�Ad��:5x�Y�`��9�ؘP-�D#� �6�K���i\r���C6]Q�|�Հ�Ozlڮ��Oe�����"�lE�!J	kU�p#�O2��$-p��h�ٍR�4i�,Ω%�a}"&?!�	E�]�pI�g�hx���ӊ|}b̀6G=6��O(�D�|bD'T�?!�$ݦ�ǉ��x��ŗ.�͙��i���_�n=Ȁ�O�)�>�xV)�0N�����H���rg �kp� a��B�=���D 
���<�d�rK�r�@��1@ܸ͡OE��+�ц����*�p���u�'�mH�h�ɧ���Qr���k+��3��M�� �X��6D���AN�#r׼$b�#L�j����0ғ{y�?��� c 2�: KIpv�� b��M����?���2e�X*��?A���?�������Ɗ̊����F\|�X�d�
���F1jT�i"G�G�m"i�C�̉O�ӆ(]^-)G�x�Q�e��:V��0
�h�����1O����B�ֲw$�L�#K�7�쉢/� )r�B7�ēSM��:�֬V�r9 '�C"z*��'�RM���K�az���]��9 ��aBt�1�y�:7Tj(" �Q�tz� �'@��M��i>-&�X��#G;w�f�K���"��R%i��Jv�������� �I埜�I��u��'�R?��eHUf �I�2�,�9�@Mp�Y�(�ȭ���X(J�&L�"șm�N�����(O������3Z��tkqo�N �8Z�ߐx; qI�*C�?���PW�»("���$݌�(O��8��'�D����F�1s�,�ִ ��+D�0He��E'����΃'���J#&D���Ã��x�UmC�e��9���>) �i��'&�#� rӼ���O��/R�� �[&<�u�Q��9m�7�Ԣx����O
���iȆ-���L@�p��M��M��!�~h�C�,���1tn�"+�n�G{���-�TA�!˳D�z4�J8i�Hຢ�:1��,�G�+[*z�a�&''�ў|C���O�\G�$��+M@I:V�Ȗ�h��u����yBC��u�(��H �BjH�4m�۰>iC����C�ox�C	..h� #�>���O��F�'�S>���lBɟ��I��X!�L
T:��Y�4#�D�BAG/iƠj�%���m0�L�?��|"�K�#95�!�%�['Feb���lP�?���+[��SW�7=�F�iam�#R���� 6�#��L�# �"1�1:�L�e�	5?l�D�g�)�i�N�z�P5i�8�a�ɜ�[�D��'xԒ�\�aΐE���˂&���҉��Kq�O��5y�b�
6�ę��ߧ�b��&�f� ���O��CM�&�D�Ov�d�O���;�?��(���u�O����a��Zg�0��ƀ��MC�a]!>o����M���Ɍ_��hݣag�"�;H�#���Ȣ,&�M�]���"�h��2y�O�T�ql	y�	�z�\�'��I;���g�X� B�	��0=A!e��r���t��t �\�t
K�<�c��_W���f��/~~F؃Ʀ�����4���Ot�0O@�8��x�C�/�8=��Ğ�X�� p��O����O���Ժ���?��O����磃.�bx)��ڝ]l>�V�H�J���$�U(p]Y7� PI�V�2�(Of�B�DŜ@RfK� ^���y O�'�L�v�,O٪���� �=�|6�Q�����O"T�)A=yM$���(�50�$1H���Q�Ie���h���A�7���B�MS �F�ȱ�yҨ�u0t���\�B`������+��D����IMy��˶1�듊?i�O��hh����U�3��w��5C�4c�����?��n*BA��k߱HD(�Ra�1G����e0��:��M��ڠH���\�D: ��<�*�p"/�Z�A�!��0C��XAX�J��F�u�al�3װi����+=`�D\ܟlZ��\��X#l�1��#]�P�I�1{��l�ȟ��?�'�(OL�g��>^���S�7�D����'�F7m������D&M�*a�f��#o�<���O����$�6w�j}o�ɟP��v�@U�I&"�'�41�L��G�ݲ�������~Ӣ�	7N�Obb��g�J��Hb��*B8� �Cp�ք�I�q�#<E�$���-��� ��;P�Z8Q �-��K^�?A�|��Iס�.�rD��0����0��N(DB�)� ��I���-w�f h@�\�LD[��	��ȟ�})��I�H�L�$uFU區�M����X��J�PЦ�	ɟ������^wZc�1b7)wZ&(S���1=��=S�._:AB�53�叶Q���)�*��)U�?���+K<A���LD-q�先��p�6�ۈ>�0p��c٘g6~,1 /�.z�t%�OB�X""g�	�E�@;ԅ��
 #�E��6:�ʓa6d��ɵ�0=a���fW������k��4��O�<�B��V����-ə"�=��Ȧ���4�ƓO�q0��0T�*}��4Dytey�LA�,Ȥ���
�O|��O4�đ������?��O�t�
��� }�V�ʠE�A<�@�b�NJu$b�nA9;-(��6���џ� �o�3�2,I��H���@�U5�
u�%�Ͽd������B6��E�Ŗ��?�U���'�^lq)]<m�ܢ$_#�&�'$�O�}nZx��=����f��t��� �0`B�ɡ-a�&.����Ih)�0�v���'��I�H�9�۴�?�������9���r4o M\R������M�d!��?i���?9��qs��{�*}�` ��i&��R�u�N�B-j�X)����$^ўp�ghٿ`�B,w-�j�l���E�r��.^ޤ�U�,j0�����+Jў �׆�Oґl��M�������
����KZ<1�2#�O��M3�����4�	�d@+tD_�?9����&� a6�����Aش1�ri�R
��h�����Ӆ^��T��]�l����;/�.���ٟh�OFt4��'W��ZS��Z�:
����PnY�,��7M�o�v�SUg��)u�%��BQ'T�D�O���?Aӡ�)0��/ ��=��"�?SER'1d@��\�_� �����u�e���O2rHq�n^C����E�T����'��Y��KR��`�z��(�'v	&�0�֙iu>�`cK<~�L�O��$1ړϸ'�� c�V/]���ZwF��`6�٣���Ҧ]!ٴ��t��	�eU��wF"7��E*r0�Dmȟl��s�rq�F�۟X����	�uw�'B����P�,s�زC��%!*O$�6�V�Q�\)KG�xg�ʧh���;V�4�dG/p}ࢣөc�ju@r��>4*�t��G�8����֔q���`T>���l��m=�'�JMA�e�)l�����	�����)O�����'������x�1�e���b#�y�ω%'!��*�p|ˁ$K*$�
��(L-���(��|�I>�7aُ,��8a�iU�m\���$L&�4���Ɛ�?i���?���T���O��dz>Q�g��nP��h�4r�jg�b��yk6	�:ό�(`bM�C��PE��-Q�Q��k��:&�Ri�Bɒm�z��r��&.v ���5\f~����r4,��I*_�Q���k�OnѨ�e�w �;�lWC.ݫ0Œv�<��k7��Pf�}��2��,�!� #4
���X�6��h�g`� I��I��McK>1�0V2�f�'��ݟ f��.:�*�ꕉ
 a��0��i|�P���'�"�'�:�k�A��k
��viێ;���ԟx�00FQ=JJ���h��q��퉇iLČa׃�aL8"Sh��rc�����Θl� ���:� $��+���D{���:�?1��Ӧ{�d�0�q��Rw�
me�C�	�vB9 �(Z*~�$3�ώ�F�P���@b~�.�,|Cb8 �O�!��s��֙��ă�5v~	m���p��~���F�.���'���EH4�<p�CS9w2Pa8��mӈ�@��Ozb��g�#��}�S�O�G>��&*$6h�	�0"<E��$.�Iz��0y� X��ޚ�@���?у�|��Ɂe�໖bA�E��ix�h��=5B䉹=�����9� ��E�5ni<"=���k���r��HQf�����w-z}cش�?i� �b��,�?���?��(���OklԗNj���F,3|�+�*�0Ğ٘�'���1C	8e΢)(PZ>�<y�?Q���w��!�t�\�7y�u�f�ՂJ�B2��ZS�Ox*mʋ{"Mݙ�$�C���,[fZgG)���� ?LObMS=��1`�\
O�M�&"ORd�B��t�8����0_t�s�i��#=�'��-*SPB�52F&h��J^0_(셛�Gըj&m��?����?������$�O��Da�:=�f(�	+�<�C�%N�@lb�ć�to����dH�N��.	=!L���k�'���)�e��1����&�ƥ��V�1,�;c��4VGj;�mΙi��c�� Fy�j�'�?!���v��/� 	�^ts	�� 2�x��'��T?�*���2>~�2��R�W��|��%��p<	V� >>ꩢ5 �,w,f���Im}�j�"Ln}y�-�� ��7m�O
���?�	�o�D������m!��sӆ�QH�O����Oh����!+�����T!|^`Y��> n�S��&\�J����9�,�`���Q�$S�I &jϔP�5��!2�°�A�ں%�$��ύ�$+D\i�kݳ=�H )���
7���k�}�B�%�?QE�S%
>���/|�lY�ᓛ?B�I�C|�5;��̍+�Zy"u�P�Ī���^~
� L}�W�'u�����&��Y �U�<�!��
�M3��?�-�8�;���O���R�wڙ*�H�Y���J�+/�z�lZ�p��R�mE`R�=y&#ش,��,�L�����|2�!	�H{fZC�H9��+�	�?!`ƃ�g��I�݊J�0%�O3g&�2��W�q��OC��Q��E q����&�?
�j��G�'�TT0��~ɧ���Yђ.�'N=��KE��\Q�防�1D�t����.yhtfD��l�s@�/ғM��?�+�jP�8�T�Y��?��p�k��M[���?���Mږ9s���?)���?9����ƞ��P �?(���w��h�ZX�h�:b@-2��P�w~��󵯁���S�t�6]@�x�$��%����a�٘��ȺD���["��bA�Bw���+B7Jph��.��du�µ?��Q�'�0�↋�7�ҙH��[4i��,OРJ�'Y���� ��9���4C�d�R�k�!�$�p<�A��6^�� �CD=G��a8��|M>q�$�P|Na�V
�9*Ԑ�$`�u|�4��"O�-q�2p"2%{U@/o	���"O���S��ck�X`�ρp�u�"O(p��d|F���o�76���*%"O Z�� �X\���;��E�Q"O&5B�dJ�>��1���[�����C"O0�1K��EW�ST��9!��I�0"O�p�!��S�P�*c��u\tr'"O��tB�@H�L���Ҁ[�4Aٓ"O��A2E�9F$e1&�0�P(B"O�q�!Q::��9�2̌�pL\��"ON�q"�κǀ��5�¨2��L��"O�݃@#Ǭm�p�1��;xp)z"O^�*�D=n%�x:7+��h�$�9`"O��IPj�/D��ڠ(��_�(�"O����m�r�<�#���	6X�D"O��"@ȇ}� X�䀌{v0�2"O���B(C���q��{t�M:"O�ĳا5��蠤L^�{pX�""Ot�ð��'���Y�B�r"O��z���9��	�j˫�d`3�"O���Wǆ�@�]����[�2"OAS�GN�����#w6�(�"Oj����!|���Bf�B'g�P{�"O&����M<����`o6kl�i$"O��1 lW�N�T��m��fw�U��"O���M�J�h�	��rX�t�"O���W`�+*��T�Y�l(��9�"O���֧�>-�����<Z""O�	��%��v��=��"�"O�����}=�4�B9\��"O����!�</�*@T���U;�"Ovy8��)e).���n�8=^���"O�KE'P�|u>@*v-��(Df�2"O��rp"�ЍC��@�7"<��t"O6�#�h�������qn)C"O@��"?k�������~�D�B`"O���k�Z�x�PA�B)d5`@"O�M������8I� ���kLj�A"O�pKU�YV,K",ߐN�0���"O�p��1:���,�����&"O�Ԁ'B�D)��#���s"O����$F`���#c��5"OY����P&�p��	1�<�s�"O��˙�ά5c�c���,U��"OY9��^��Ђ��5͊y@&"O�$+r�óz��Y�fϋq����ȓA�جР
��6/��5E��4��$��s�Y��)	I�iK����?Y|���nL�L��G�;c;�ՌV �~y�ȓ;2��%��-HiB5Z�Kܐ^�*��ȓ��YC�HC�����[�+[�S�? z؊V��L� �#F�E�b�$��"OT$�A�Z�`���7��욠"O@�b3EF,�A��܍t�n���"O���ΦN���� �ɓu���pg"O�0��V�d���BpF� �d���"O����G?�A�ޫQ��w"O�ұ�-}Trɓ�!�%�,��"O�!�7E \�b���(В�#@"O���ᐪX�m��(|�0���"O&��q��90��VN��X�x��"O65��������ƛ!�R0y�"O*5Z�nw{�$K&m!D��m��"O�t���6�YT����4���<�F(�e��L��̔�c��'hF�<!_J@���A�y� P('�B�<	��Iٌl�a&	1G�lA ub�Z�<I�g�S�h��D� �Č���k�<���#C���&CP�<|x(\Q5!�D�'z��B���)mf$|S�˗5!�d�j����҅%��ˢ�ٲs!�LOl�(�5g�<��&���O8!���;/e�๢��NDtūŢ�'j�!�D�,q���L�&~���W��) ?!򤂼S�t�zt��Y���vn 4�!��ҥʛ�Frށ2��W����'���0 �K,G* `��A�+����'�p�vET77g����,�(��(��'� �K  Ň&�E�U��\ʸPp�'�D�� i�\I(Bk�� �&I��'<��B!F�&���r!2�x���'-�8�oDnGV����X?����	�'w =Hq��$�����/rE�E�	�'J.h9p��J�d��bhO�d괘	�'�&5I��Ή^{����I�ϼL��'����c��$AB�NM��P��'��ՁtL��o��@&�N�06|�
�'w�܊�o�/I�5"�k]�ji�q��''*�SC��5pa���ܢ9��M��'�� ��@�v�9��]��XZ�'�\,���.%@X]��b^�U�.]k
�'����ʂ�ohP1˷n�x�Ƅ8
�'��h(�EBd�($�%��^/� ��'�0A��K�>�j%��A�(^�=��'N$\�$�^�|"��e`i�R���'�:|��K�9}.�l��/_�L�*���'�0���2�zp#�MAn�q�'��%@�(�!n�n@��V&��	�'�~i���([`"�A8�
�'�FĹ�@�k�@LQ���$x[&�:
�'���H���Xr���-�&���'|$���H�/1���[B��$�b��'ߜ!C� 4y"j���� �^�Z8�'��	
��ԓ0>:�E�_��@��'����҈ȱV�ܓ��	�j��
�'�4Z�*Ɗ`,T-#�iܛg�M��'�r�C�ˌD��c@�CТ�'�����W��N��@�2CǾ\��'R� &�=��d�qR92�D���Ei�X	%�.��7�)*��e��G֔��m�*�x�P��L;\��ȓ8i$m�Q�DO�Ͱ�FQ�BJ`i��z"�bT��4[�b�?*���ȓU�f5��O�Xc:�����'�y�ȓ\!L$�
�c��(
L�I8Ƞ��S�? :E�HO�-wt)���5�� zQ"ON���j;׮��M-_���SA"Ot�(U�G/��=�C�Q{��i�Q"O��H�k�)��`$�� t�~ `$"O2 ���7j>:l���}��x�"Of�!�훪0�&LCeaѾe�h��"O�A˵Wc���TKQ,nN�"O�(�t�؎axt�#��w{��"O(��0i��j`�u@EC6=^��ʠ"Oô��Yت��àC�u���;a"O(봏��d+�-�c�ב,ᒜS�"OJ�h�D�'j�H ���~��la�"O*���Y�LF�)�L�Fs��C"O�$�Ӥ�v�Y���a���"O��IGi�R!{u�4JN����"O���K�U��q�י��"O,�>G�"-(QT�f=��CI��y��
9��L��(���yA+V�.y�������E�yb�� #����M�9<&(�G��y��l}x�l�2D7<i:�����y����Z8����we<8i0�G��y�d\�
ـ��y��ԡc$M4�y�D�1_�8�$�C[�ޝ �E��y2�B)y��u�тQ�L��U��)ޗ�yb�Y2���I�m�����*F��ym
h-�}�p�+=��ʳK��y2h̭yB\�F)ޮ.�����/���y�$�3Q��e�t/3_)>S���#�y���ɸ�0V�����K��yR"��9���-�R��V���yr.��[b$�XU�&��*M�'���h�bQ��!�I�
�'����ص�z�k���.r����'�6�Ԅ
�a���hϖ0c�ة�'P����E��Lέ8�
��.��i�'I���LQ��n�� �*�VI��'#�0蠯�2K��i�ŕ�&� ��'J,��WA۶u� �L�  �5��'P�A�WiA�q,)�b��f+���'=����8$���Vf�6&Жe �'K����L̕E�n81�*��\<�P�'eR�ׅЖm�!��Q|���	�'*D�a�ƠB2j�$��\��`i	�'P��f��'�V�sf�)�<��'�ԣr��9IV9���6x.V��'�fH��Q�9|$(����t]�T1�'g�,	E�F�������1f��P	�'�$�:#.�y�X�ရ�-�up�'�
X�b���f������T>�@�*�']���q��W�������:��'P �j�KD3D�%�� �?���"�'��ɸD� "&��XQ��#jb`j
�'�>ـ� _�E��m�K" J@�H�'�j�� �G�P�֤�AϪi�.P��'BԘ�j�� L����닮*� ��'c��%��(����&l��M����'�(MQ#��	�����#Kw��,�
�'<���\��`�����6@���
�'�N�3�ŮF~3�ᓒ��|k�' X�#FK�5q��a�+�����'�b]#rA]�M��D:V,�O�jYk�'�>��0Cʹdbච:xrȘ[����aG�O%P���b�)����),D�� �ԛ�@�;�D���l�Y㪠�2"O�*�ژo�:���Z%x�.�CT"O�xCo
�D�ңچSݬ-�5"Om���Z�F���!�l�M�"OdB$/��:3<��a�@�i䂼��"OD�'j��ž-!l �N5.<��"ObI���N�b�� �F#V�=���"O����'��D�\�xA�C�jvupp"O
iD��!0p`ar"x�l�Z�"O��W��`�&0�2(�I���a4"O�r3��?N�Z���H��"O���#(�3w�IQ�H��F���"Op�B�bS21Ќ�:F�w6R!��"O���B/#�&�/�o&���"O�
�K�E�h��4?J8ȓ"O���1,��
�"����.I5�Q�'}jY��gP���P���b����%b݌��C�	,F!�YA�W�p����n\�6C�:��H0��Z���jgi �XC��:I֨2uhZ e�0�D�`XzB�I�#4�:���O$8;��45@�C�(Y���R�#F%��l�%%XC�I&Z |��X�2=�ł�3o~C�ɛ'�ƍůX=X�ЀBg�֭N��B�I	!H��@��r�`�ŬUښB�I�e��-��-_�LQ� G�klB�	:e��ٙ��O:M��M�X=�C�		v�	i����~d���H�{p�C�	�=����
m�-�v�FFC�ɐ� Pl��S�� ��'pLB� q��Tm��+��Ѩ���okNB�K��9#�\,��pv�ܡw�4B��2]�$�I�)Բj�i���E�8*FC�I�$�h����Y�%�)�f�:$>C��.9���CëUP���duhC�	�	e8���H�B��gg_&hS�B�	�ު	�a,J� � ��-+'�bB�I�T`�ƀ˽U� c�A9 �*B�	<,�Ț��Ш�f�_5�B��-�s�F3���o]@x�C��6j��	jӬC�z옅lO1^��C�	(w܈��w��+Fll�(�S&oM�C�#p�l z�Ȫ�(���$�lC�I$IO��F��:n�F�C(\{jC�I(m�<K��Z C��R4N��)�C�IQ�trkzԈ��T���9#C�V4���D�7�(Z$��xC��7%QtQF���� qA�+�C�	1Wc�ꅡ��&Z$[�@<�:C�I�{���!�!E�W�f�S`�
p�jB�	�~��ݑ�@F;͞����IJB�I>|F}�Qa�*P�T+u�F�-n^C䉑^^P�{�R
"����4) C�ɥ]H���ዜ�$¦�r@NB�f�C�	7b�XI��хO�~a�f��(	�vB䉎X"^i�����j]����>B�ɼe��lp%�\��k�T/j��C�I�#�avB�}����'��C�I�V�v�U�F����E�˸>жC�:6C�X���	<8�hf�'�B�I�S"Na��Ĵ?�P
'�Ny��B䉟�\8���1F��jO$"��B�I,O��"S���RNt���.W)�^C�	�g�.c	H�E��$Z��-??"C�)� ىՄ������a�}ǚ�)�"O\�" ,�� ��A&��Z�<h�"OH�A�6I����vȅ1C�~��"O��!n˯V�1�vaŴ-���1"O�X�.K�k�(���x�r,X�"O֬*�R,#���@R��'�`	H&"O�!Fљ#!���v��0�ȸ�"Ot2�TRV�p��r��Ց�"O�H04)E�^�F����¤j$b�"O�X�A+�&�b=��o�9UrT "O�-�S�	�BMj]S&/��2H����"O`����حp�ɠ/�/h@P"O��� ���h�b �ȤA�z%Ad"OZ9�@/ćymd�ɧ��<���
"O<�v���$1�`E�<��F�+D��C5� �`t0b�? �<��A+D���Vm�^�l�� ;��${�;D��v�ܣxክ�c���ɞ�$6D��(B��r\�u`�`��%f9D�\s�M�<>�����9+T�	7�9D���'�"M`�ѳmȣY����$�$D�d`N�h���sC�a��OB�<�A��>�f�ŝ-|i6<�(�@�<�b@�<�񮎮a�FtK�\U�<�g��C���EM�hWB�֭�H�<�(��^(��@LdؤE+��Zz�<�������K�8m������9I�Q��F��'ivp��)������@UR�{G*D�<�!�=g����V��P{�)D��r�"�b��H�h0^�"�k�=|O���N<�6(�6=�"���	$q� �S�Ao�<ٱh�*3�EQ�	��"���葮F�(\���O�"̋&B�-�q�D?���"�'0�M+��.X�B�;�I�|k�]s�'�����)O2;��)���yv��'�2�;T���,��Ԙ&�	���p�'����5��s�Wm��m3�'M6�*��Q&"\ �boY%^-��2�'�,��F��wIv��-^�?v*%��'l� ��_� �`2E�8�Xp�',8ڡc��z(mSJ�}"��'� �y2I�7Ai��Pn'x�s
�'�~yh��=z�(��H��hc����'Ɔ<�vj�67W������#eU����'0uSÆ��6��rPɒ�t�vd �'8���GXG�J����H1$�d�x�'`���q�B�>�:D`"e&k(�z�'�*@�KZ��(���)2���{�'V>4C���������|��)��'���5��n]`�ubs�T��'\�EV�wU��K��_ac$ԋ�'��()���~���A�Sj�e��'b���kW%��4��	�R���'鼽��ē	~<&�āPW�1��'������!�Zp�i�O�|�"�'�����H�M
Ii���1Nܩ�'��ha,�'g����|U:��'Tƀ�5���rD��VD�.B�x|c�'��a� F-{ERD�%#��1Q|Z�'����
ż~��U
�wo�tR�'��|1��Ѧ@lH��.i�v�!�'����k	/#S��)��ݥp�^|��'W�� ����o�`R�+n�ȡS�'X]�eX#2*"�a@�=�6tC��E\P��� p�jdg�Q��bŌ��iyf]he�'�xl&���4��jd�� #�>o��d�A�>D��	�G^�B߶yH�C��]`� [E"*�ɳ
9�3�!�':��r�'7T�IѱJق8�	�ȓ�����,�t����/�-ː��1O�<��4	r����L<�!�8?Ѧ� bmU!A�Y2hOKH<y1.��(���'OɜP�6@yc��+�6CQ�榥��	�L�6,�1�@�l���2ׄ��R`����J��MӴ"ZyBi� ������zծU�%K��y�I*}֨�
w�Y�n_y�����'��	Ӊ���&��'�xEk�S���U��y2L�@�e�u��7v��(,K�ў"~Γ2'|-`D�O8VE��"��jlM�ȓ|"@l�3I��|R�X�5�Ѩ(
�Ln�+�2NA�#��P����G�f$�#�E��=�P����	�.�6�
���1:�Ɍfd�C�	%� �ۀ+�Zb�DB6��AA�#<� ("�S�$j��2T�m�"`Ë*�Q� ��yb� i�:����D�������P|�9Ey��9O����QS:���W�.D7|�B�"O����ɍ�BL��/�?J\���"O<�iW&Äl9*��Q�Y�tS <��"O����Ƌ�{�S�k+00
�Y�"O���Q]��������=����"O�-��@j�L	&"�h�j%!�$�75�.M:T��#`t��k�  �!��]j>�e(�5H
P��䈳~!��ӿpU"M8d���jHS�$!���R?���#[%b̄�z�!
4�!���'���2`i�i���G�^/!�DX>V��1�A�9t�����[�"!�$�o`�GN¿y}8�Z��cs!��06�aPF��-vX��	[�q!�D
�hŀԃ���tL��1�/J4MT!򄐅A����HW,��-�C.Ҟa�!�$D�g�<�P��ؔ��*`M��6�!�
�����4H�U�~1iǋ��Eh!���3KXD8`�ʻH�z�"��t�!��/\��Q���U`����,@�!�D�	q^���NP�N\UC�J�b�!�D�"'f�H )V�`�F�!�ě�f|����9iaB�*�#E9 �!��[�1h��U�T[�]s5�+>�!�ْ/9bi�OBtQ�M+l�H!�D�'u���kfC�=52��E��,S�!򤉦�-�Q�?1~�+���gB!�D��tW�}��`[�&�B��S7!��Q�ږ��V�V�,��)��ɐ%&!�$F�a�}P�J��|�:GA�U!��0���c�Oc�ARb�E�!��Q'jG~����J�j�i��Fh�!�Z�H��1��)%)DMa�K	��!��Q�l�&��m�%n�P
�4�!�N�[8�XƂ�v�ْC
�Wy!�$H �lQE7 �ȥ�F�5c!�Ǻi4H��i-22�[�,�=XH!�d�>�
�!p&�*�mIP�A&9�!�JNs�]���'l92tA6+�Vt!�d9!]^�`��H�%P@LKjt`!�$׭a�աV�X23h}Z�hbX!��ϡ_�z�R�����MT�2�!���l\h	Xo@%o�	����!���GzvI:�oR�i��I���O>7!���5d��TEzj��@ T�E!�� �y� �%E�1�f�
G�.��"OXL�����00��s�EQ	��M��"O���� �DErf�A��d\#T"OFp��c=B=>�#m����ӷ"Oܤ*�%"��bߟ}����"O~����X�.΋X'��R�J�I�<�����re�����T��5)�ėZ�<!��B����CŌ�.��e�I���y��.͆���)$E�]1wg��y���1�f��@n���L��� �y�oӮW����22�X[���7�yR'܋r�X�0�+Z��J��y���Q������0��<c���7�y�`�2v�{%�WY�tI��.�y��(s�U0��G�S�����<�y��if�h��GR��	s"Ҫ�y2�K8hkܶS
9�t ��y2��-bBt�,U���1G�Q����&��D���Ԇ��đ�ۡ]����ȓd8�)��Ӂ8�t�E*J_(���	�& � @�?   H   Ĵ���	��Z0s�)ǈ7U���dC}"�ײK*<ac�ʄ��iZ"w�F$x�Y�	a�6��LMX�{�gY�:��`���O�}*��Ԥ�1g|�\nZ8�M�c����cy�@�ɋw�<��	� � �Q�%�$�SQ+l��ã��-j��Y�]����bW�Eꄥ	K�`���=|�S��iܦ �5+��6O򸒆� Z��ɚ�Ό�
E5��ɋh��2S�1_�S��1CO߷(��%0��2�A��Bڏ5l�p�J��jw� (j����@U��X�.c���A� e4�I�e�t���
�7@!��R�8�_|��$>����>"�B��NR��gF�%]I�Qz��ם��p�\�Lq���<�O��آ���b��Y�'�� ���ޞa�� ��Թ3�h�*rL
 k�F�Yybj��"N.��nX-��G2��X�!�O1D��tj�.b�� ��X�4PI�i?FdJ�ɍ��s��!f�F5�C	�<�N��	z�Mӣ��1+�����<�-�6͛LOs*����,c���nKk�9OЕ*d��2i�=Iʕ�V �B{���Cb_;`��dZ꟠�U������;w���%;���b�D�_�4Ta���!^m ��Z�oQ�d`��i�j8�	^-�-bd\����p�x��׈�w?Q@�i�t��F��P�FT �C�v�!SD

� �J��ǝ|�� k�B�M>Y\c,�Ӷ�QW6���g�
[?ڙP��n�=�,O�ʦxנ=
O>i���sTQ�^>�D���0�r����M����'�bY��NP��~�u� Q��	8w��?k�d.�
qK��Z�)v�C��P�(�`�T��%��%�x2ǚ2��!��*D�A��=AF�N耹*�,Vɦ���C�+$ѫ�i�΂$g�
Ha	O:�^w������ug���P>�|���

��ô	�$6�	�l1��v0�$�h�����x�Ń3f��-L���B�	GwD-q�N��u� �9N>�g�+h����<q�E$`l��K�cQ#/0�*��~��S�"OԄ2Q�  ���Ȭs*��@ȏmuN�[�"O�����ި��L����r,��"O�%��H�D���Q��p��2"OHU���(�d���I��"O��Z���n@ѳ���FP��"O�iБ�y�v��m�]8��"O��kW�Ci S� �\ 6��"O�iq��
�W�X���(����"O��     �  K  �  �+  �6  �?  WK  �S  
Z  S`  �f  �l  (s  ly  �  �  2�  s�  ��  ��  C�  ��  Ʊ  �  ��  �  ��  ��  ]�  ��  ��  ��  ��  � 		 �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4� ��eëF�ڙ��n��R�pA�O��B��M&\׸\�ELHw^��p�'�qO��a��aP�p���
�Uz���"O���	#GP�7I�&=4���G���q���S�x��3Fk ��D@�C�(_�NC�I��b����D�fi3��U0�,O�]�ߓm(��ߔvd\S��*E�X���Iu�H9X��ҪY~K\��'�G�D��� �^=�4'�4�l����& ��A�?ɍ��~2��֨C/��C�H��6D�B��FA�<���4"T����-"�6镣���hO�O�l�$�TA!�ڰcOr|n�j�����l�<���-\��\XSA�k�(4ks"��<ى��&� �@k.��d�q�š�C䉳��I��g�:���q!���D5��H�a}2"�)T�V3��X,�U�Af��y�'ǯb(p�E3wPx*�� }��O��d(
��2M�(\��ꓡ+��}���P�U�7 K�Qp$�|��8�n.D�  �U1�� �'C
˲�"fJ��'�  �O$"��3>&ݹ�`��8k�I��'UĨ�˙^4U�W��:wL��*O�YEz��C�G�IA�MA8D�x�2���pN!�� j,�@�2?M�ݢ�R&��,	��|��'��I��˖�3���P���'n�|(L<��/5J����7`��.<0��ȓ5\�����6�\�;a
?�Z���}�'�8��"�֭R�\X��^���	�'?�i�fG!QN&�!g�&�%!�K�&�Ob�Ũ�(HB����+��)��sX��F{��i��Rv�<S��@p�XP�����Yl!�.X9L�c���47*(��ŷ|���o�`9�4�E+j��y@��K�4l���"O�,�5j��IW��0�ȦYT>@�4O�=E��Ǯh4���U'��Jh�}���yB&��^v4P���ؑ@>��ɣ�yRH�VG|�̇�9�<�I��H���	W���O�fE3掅
�>���A@#��a �{�'�6�
d]�<�^y��O�U�2Pӎy��'�< ��K��=��U;#�
>��P��'���B��;Z*��2(��Hy~P�
Ó�����Ԫ�'8ł����,XE�LB�6D��YU��:����E��&�'?1���7�P=r�㉰m*.r��F�9���hO���>�� \&�&��� |���Y0g}ܓ��=�$��=j%i���2�h��|�<Q�*]�s� ���D�;�&)��~�<�Q&a}�=p%*�N�&����T�<��n�.wf����9�\����{�<���R�J��K��B5���G�Ew�<9��� 2X)7HȪ[l4S�	}�<�@N%!�D(!�Y�J&�I�k\|�<1EK?��H�OT�tHLQZ�@z�<�ƫ�7)��q�t�\�"����y�<����6U$pq���a�4�x�<�W�<�8�s��Y�<���L�]�<�!-7mP�x�8,��k����<�!
O����B@q� ���c�̉��+�OH�J�b=�&Jj�`[,����QB�H�֌# ��rB �R`̌�ȓv��	b�S�	��Zs���Sn�8��5��Y�画n+^YRt+\	��!�ȓf�������
�t��5�mF�ȓ��G�4B�	U�'R�I�2"O�# �D�Қ�H#b�F�"��D��(�S��Κ+24���C�f.t+&H��x�!�u�h�Cn�O��|KgȔ%ў���	�9�&��ũ�'�Nͪe̜�%�C� J�8�Ɏ1l9ҙ*��' �C�ɣt�z�if9O�t��օ7��B�I�x'�K�dAci:�BG�@b�C��;c�s5�W/��O�(t� 㟸D{J?��'�	}1�����ҝ&�qc ))D�(�Q$"��h��K)w�U�#D�\Z7!U+C�B&�Eqۀ��%�!D�;%	[�15L��#G�* zE��?�2��~2vF�	�PQ)�%�-G�I�W	Ax�<�R�U�y�P�SOzz-;�mSs�<�� "A�ZI�!�J^��ʄ�h����'h� �P�O�f�ҐNX�|fp ��'�v<�d&Gf@Yũ�#��dӎ��5�'V�l����NŖ�b��z��xf"Op�ه!Ծ<��dR%GǱ/6�$�`^�h�I*9y�D-?�K<�O�($�g�l��0�	�)A(A��'w����Ʒ$��s��T%�̵�O@�<����E^�:�l��tm\�C��RT��,�'��+p��5�2X1'@J�1i	��� >�1D��*4b�jBej<�U�'��#=E�DmJ����2�
�0�|̸��i!�[�8tF�#�c�^���E��8{<B㉱=�)۰̈́<�NM��D�(����*�	)Q%$����S�*�d��*ᶓO,�=�}ڣ�S�2�dt9�NW3}/��ԍGq�IZ���OW���Ђ�+D��"'ԡ(���'�t*����"��*�;R��ɡ��m�R"<E��4CB�`��ş '\�*��1J����	�':,Ӄ䎐o���a��3ji�᧣j��=�f�i�����%��ȫ�H�#��ɘf�2�O��G�p�J��nQ���e�S�#l|�͓�hO?Q�Ǖ2>o��$���9 P5H�@8D���I��B5� ��	j92E�DFw���Irx������96C�e�S�5�Ze��@#<O���n�������+$XeP�,S�T�B�	����i��$��,k���$6ړd�����Z"sh|�g	�g�PՅ��E})���J= V굣�ޜ��It���O��y80-��"1����+��	Y���)�Q���k4���Q�]�K@�)\ �ȓi�2P��c��`y3��RnY��>��������(�����4�]����P3&�\J��Q�L��$��S�<��Д=�ȹC�gf����	q}rFł�|)�gȆ�QGV8B!�9�y�I�V;�e[��Q�/H���'��\!����e-��+
Wkɮ�j�'r��cV��Xݰ5���|m{
�'Ӳy���I�t��ԺS�4Y3f�`
�'h��ꖶV�"AT�RSD"�0
�'r�x����Ya	CC&�!N���
	�'�����
��e�U��m�+O�l�'+�s%��0'``qwc_�3�����'#*�S�b��dA����&��9a�'��-���!o�<�g�,����'� ��"@
e`�#�]	�J�C	�'N��O_$^
h�a	���i{�'s U��E@c�����!�F���k�' �I���Ca�=��G\�tZ�	y�'$��	 �qɢuP��[ j��	[�'"�����!U`�H �
�0�:l��'k�z�k�7N�`u�g�6�J��'#>t�caH�
�\H`�
����B�',�(�,q�x\A�AW��dP�'��uЁJ[Jt��o��&@�'9�A�f#��L�,�6d�z����'K>!BÀK3[Ԫ(��ъw�Xl!�';�Q�q�F�B����F�}��I�'1����H�,�&�hf��
;0t�	�'yd9f�I	��-�O~��z�@B�	*��}�'Ȇ%d���R#H�cZB�	�n,<5둈A�*��4�%>�JB䉬:8���J�	�����\2B�ə^\�8bA�����]�3 	��jC�I�. R���䈺?��5���A�w�vC�ɛIRvpS�IѰR��%��8q�jC�ɔ���C��ǆ$K�$�!oU�x�hC�I
���,B1����&�\C�I�:�K��ڊ9��ș�jT+)YTC�	)a�y��N�=OP�����O0L&C�I� ~��k��1�*=���;){bB䉍�r=3gmY�`���CD�'�B�	�=j�&��H{�:�̓j$C�)� R���_-mސ@��T1[T�A�"O̪"�9[�H
��̳��<+c"O4��&!ȼS���t��"O�CT�	6ӮّI_R(#"Oz�h��9s8N���"4��tBd�'�2�'
2�'���'B�'�2�'���b'Â!"�<"Cn6q�$B��'+R�'�2�'1��'�"�'�R�';@%�4�ثdA�cDJ#Q� t�',��'���'���'7��'4��'���t���=��|�m���'dR�'�2�'���'$��'O��'(���1A_5;EZ(`���w���T�'��'�r�'���'b�'h�'\:5��Ő�&LL�)F9�\Q�b�'��'��'���'��'���'H�Pb���<��P�H��D��YhW�'���'���'b�'�r�'��'�B��FHh6�K"x�\�+t�'��'�r�'�B�'R�'���'��u�e(5��\k���Zt�P�'y��'5��'"��'E��'P��'wP؁&�D�T�lñ/C8V/|�s��'m��'���'���'B��'%�'c��� �[���#aL�9,cBXA��'���'�b�'�B�'��'i�'�b�s��Z�rx���<Z,�HT�'��'��'�R�'d��'&��'���#�}ݘ!��M6��AJ��']�';r�'���'c��m�D�D�O>M�ԥ�=���I`�2fE�Gŗty��'��)�3?��it�5�ШӅ4������O���SEd�?��D�Φ�?�g?޴A�����-�.Ⱦ%	ǫ��FtfP�i�BD�-z�!�O0hT&�l��J?3��A�x�x�G��
v<,(��1�ʟ(�'(�>Q��m�4�08��D�/V"��K�-�M���F̓��O��6=��}3�̂$NG���&_iV�Z&L���Ln��<�(O�O�@�`&�2�yR,�@��Ș��J���l�����yb̌8zx��!k	
Mў���h�",@ �۷��"w�0��#ju�Ė'��'�z7-ھT�1O���H��,��.��k��@�-�I��d�O�7�o���'`4d��d^�(�A��e�%���Of� �ʈ6�) ��i@�5^�9��'�O�	J�OوU#H�� �3W���r��<))O���s���N,tP��,�B�Ѐhb�@�޴����'�6-2�i>��!�@]� ���!+J~fub�N����I����?K"���!�<?E�-d��1�#�"�[�"9<a~��O&1u�H>�*O<���OR�D�Of�d�O�ۂ�$F�	1�خOk�,�.�<I��ivA0��F�	�r�'��D�O���'�Z쓔�^^��C�O�1"eR�!�>qƳiM�6��� $>I��?��T��z,������"�4Qo^=�R��G��uy�
Dr_����Q�&����n����AD��*J�&%���'	���se�=`zT�)թK�d����a@-y�J��Ԃ��x��ʤM�?9�ў����# ��X2�ܚA,�1� 5�I�b�"��BJp�kP��==�~���,|�)����-{%^��G�:p����Kp��c��r����/�AG��7OM�8�ĭ$L| Z��D-c�n�G؜��Pd�4 }�%
W7Ŏ|��L�Y��&��g�"��r�Św�X �3������2���X3�}-�ổ]�G�6����ߦ��d�O����O4��?)��L�OHj��v,D�O��xc��DJ�ܘ��O����O���<!��M��T>��v�$8�	�ħo��#l�M����?�,O:��O�E2���ǁjr}+A* 5a�,s�һ��V�'2\��˃
A��ħ�?���SdKF04o�D{��E�rκ)�3�͔'-��'V����I䟛F�\�}�~�� Gĥg��I���&�M�-O⤰���Ȧђ�����󟼁�'�TRc*�e�Ɣ�t���B-��4�?	��RPj,O�i�O���x�d5U�졙���Ii�(����M���C>Op��' ��'��dg.�4�>�bf��C�,��e"�
���R�ҦA���Ey��'\r�Ϙ'r�ӌ*��)�BR4J`�P�fS�<��7��OV�$�O ��b�Lu�i>��Y?�q��O�^(���@;�tt�!��o}�R�����-�IӟH�	��PBMCA�TY�∏�%�Ӎ ��M��\�r!�Ɛx�O�R�|�%HӤ:�L	,hlFB-APL�9k���<���?A�����--bbT�үT )\*l�휈À�b�&�U����������'��'��zG�ÑPz���N��\%It�Mژ'�R�'qU�P@��У������hNⱃt��P02��E������O���O���?���zʠy�O=�8{A�@�8y0i�t��7W�Zܠ�O���O4�Ħ<aw��%��O�^��A�ԶW�&�`���Ufn����`�
�D�O�˓�?!�
�`l�~bfRzCV���ɟW�L�J�dK٦e������'�iɆ�%�I�O����:�p�#ÛY=&���/�	3�^��6�i��Iݟ��I�E��"|����z�#�+��c��Um�{��f�rʓdX�:��i9j��?)��'��I0�����"�%14�F�@9D7��OZ�dƣM���S�4��ē+Ix,�1Y�;�t8Z"�ҤDP�-n��v���pش�?����?��'k���dgA)F��$a��?�i��L(�86��R���syb���'��j,�!{��X�5�X�q��_*K�6�Op��O�d�`W�i>Y�	h?�@DYx6�E�iW�]+�ŔO}�Q����'�I����埄H� ��k �[�2�xb[�R
�W�i��)ڣ��7��O���O���Tu��OR�Hq�'� ���M�g�0��[���$(5?���?���?q��?)S�/e���$kܿQ�|,cA���͒A�i�R�'%"�'"�'��d�O�`��Ȯ#2����/|��!I7��!-X�$�<	���?���?q�Zz��"B�iFv�j�f�zbR����->��9�Gz�<�d�O��$�O��$�<��k���'2˘p٦�@�:X�X�Ш̾�z�P�i���'Z�' ��j�e��i"��'�T�8��ƒ4Ǽ8�Յ�U����Dt�<���O���<��kZ6�ϧ�?a�'�.����7�0XX1��2PL8�4�?����?���]�`X�ik��'Wr�O3�)�)O�'���&�A�yꈈ	�b}�0��<Y��6<
y�'�?.O�iجP(�Z~�b��ďo���ٴ�?9�l>���ǽi���'�B�O�t�'�
5�3�يW&B@�� �VV,��>9�<4������|H?�d��
(����S#
�?m�e�B�m����E
Ц���ٟ��	�?��S؟L�Iݟ���	�{�3�A'"FD��$Q�M3�Z��?�����4����P���v-�<����=�2�C!K��Q��l�ȟ��Iğ�Wݟ�M���?����?y�Ӻ��X����9&aD&��I�SnI��	Sy����yʟ4��O<��X,/�ܩ�wH� 8�1+vg��]>0]o���؃a.џ�M���?y���?y�\?E��DքH�����
�쪣���>iB�nZ�6*��B~�P�'{�t�'~R�'�� TG"��چ�ɳ�d�:P�T-��KbӺ���O��D�O^I�O������)!�)]Njف�KW�N�YS�����_y��D���'~B�'e�:$�f�J��.3N8\���T!6�+v%�Ѧ=�Işt����	ly��'�� ʚO����U�0E^�|Iƭ�N�޹kq�xӨ���O����OL�O�$3F�n�2���O��9��i!���Gk�g�4��_����џ�IYyB�'���Of��O�š&T2�F��W!�R�l���i ��'�R�':!��ml�"��OZ���H�Qbe��S���	�cV�H?촱n^̦���jyr�'v�T(�O��'�$����M�7hV�_�T�S�� 5��xB�������ʟ���5�MC��?���z���?a��?=~����K
=H0ո���S��IƟ�0#�͟��	^y�O6�T��,C5-�;�И"�3X�f�m�|>���ݴ�?����?!�'����?���"˺ؖ�%lJ����׸0�P�J�i��h���'S2V��Sv�ܟ��5�:F��
�C�N�R!���R�M���?1�R��a�t�i�'oR�'�Zw����D��k�D�&��	�
���4�?�/O��314O�����ş�ٵ�\|���!�fn�e����M[�"G�A���iR�'AR�'���'�~��2({�|!G��sOl0��d�)��DԅVe��OJ�D�O�D�O���O��ҏ� ^G�`��`ڹdS��@� g��lZߟ�����$�	9��I�<A����k� wH�|�Jֻa[����f�9�y�'��)ĐbO��'A"�'�&TSVy�pBA��Sx0�P�H3����'����IğL����@��Py"�']�
�OA�� 둮L��� M�-���i�b���O����O��,���(�\?�i�A���I�)��q�'I֝
r�����g�6�D�<����?����TΓ�?i�'$��_1c6x��IB�@�ش�?�������Y媁�O��'
��bܝwS��QW�<<l=����qC���?����?����<�,���?�+�-U�'�c@��7r.^�)}Ӹ˓PD��KĲiyB�'��Oq^�Ӻc��W�<~IjTb�w���Q�������។ �}���	oy��P�u\vɧ�ܴc����T�C)^ۛ��M�%^�7��O*���Od�ɔv}�Y�L�R���7 X	�N�_w:��H�M�e���<9����<�SП�z��	�ak� �%U�HB�/�:�M;���?���\�и��xr�'�2�O��	���g�R�j�A_�Z0�G�iB�'w"t;���	�O��d�O��ȴ��2{�`W`��(�z)��M�M�ɻdyL
M<���?L>��J� &\��������;'���'��P�'��	ٟ��I�0�'=�q���6bp�e��/�e�Æs`�e�xb�'�"�|r�'��eF,h��5ұȆr�ʁ��Gנr_��	��'-��ޟt��쟰�'"�XPw�i>U�"��� ��"G�� �r�@#�>���?9M>	��?�pMX�<��`+=}�+P4n�z�A-B�<�	Ο�	ڟX�'a�P�FC7�	G��>�� �p>�Qz��\�X���m�ߟ�%����ߟPte���O"�cѧܧ
�l�
���H��P��i��'��ɼS���K|������g�4%��E�g��bf�;H�����?1��
�v9ϓ���z��3I�-:�
(�j��w̍@}���'�2g�~6�6��O�˧�rv������Hm�=�J9Y��c��m�����O�d@�?Op�O��"�����&g:I�Ci�j� a!�J�M�VH�$Jq���'IR�'���F.��O5�g��8Q�r�h��رtO�)a'�ʦ�3�k|�'����O��H�`�r72hS �]�`~�:Ǻi�B�'	҄�
U^O���O�	q8����7E� �ÍX�Z�N7�'��֯@�z�&>���H�I6�^�2�\,%@d�h�G�d,BE�ܴ�?�a�Z�jN�'���'�ɧ56��lCl�Z�@�7�`�g���d)����<Q���?9���HFTn-�g�@B����-XGXUȰ�	B�	��4��W�I��0��A�"����ٻnK�-� (��I�ϟx�Iߟ �I柔��z���S�MJ�7��M�? ��aD��8D��%
<�!�0P���Iş$���	ş�h1�x�8��%hZjQJ���~��1�1c;��d�O,���O��Ls8����T	ڎ�j�p7��
s��0�w�O
V��7��O��O���O���#o�O �'�f1��[�BV-��� ��<��4�?)����>�ȉ%>��	�?q�g�6t�$�������$�:�ē�?��j�^�����S���gln��߷���fN�M+-O�-�`H��qЪ�����4��'��}Xq�� ���!CVv9^���4�?��A��X����*�		��Њ#K����@G�	�Mc��	r���'3��'@��..�$�OBHh�²Z$�uf	�
�4ъ7.��͑���&��|��IS�%�D�L9i�|��g�/R��j��Ўp9( 2�7�0>)�+E&J���>���C�b�� ˑȌ.�ꔈ��ǃ$�p�='��T��(M�2xT�(C��-K��!���N(s��tHB���8� �R��73��4S4-F� Z����G��pSґ.�$-:�,��[>�9���-�H�	�կ�	�!ߔ^:�\0�כ:�)#"-�<u`4�i6�V�$�v�vd��.lޠ8G�O0���O��dЙK}6��O���!�ץΆv�Z��r��!p2�xrnG�;XPs���0\nZ��M{FIU�'0J�(�P�S1$X��/���Q!�3(e��G+�/�t	�ѸiV�6��uBQ�,@'D�Ol��J#�|"�ć"�p���-�̢=)���īY�45��hG��1BW+�!�+L�l�vM�����@�Qx&�I�M����d�ym�埜��a����TX���X�p����0BC�X(E�',r�'8B��G��r-��!ٜa��7-�|2�B�P-���p��:�n���!\�'Y2T0��kDf��s L<��'MȬ��#hM�8x�G�2ey�Fy���,�?��i��6��O��'G�@�H���1��P[���$u���������O��'�`+׎�ž����BF�	�� ��f�}���DX
C�����o��9��&����Lz(um������|��M�+I�2�'��J5��C���KOnI���ME��1���'$�l�"�H�,G�*A t2���w���;N��Y��PT�M5���(�
����y�t��a��Y�̀v�J�3Qi_��Ͽۓ�Ö D�SԬ�8cX`�{�炒=.8la�iϛ�I�<%?M��ay"Ć��>��7蒬8f��j��y���[�^݃���;O��k��+�O�aDz ~��D_�q�S�L�$Ufި2#�8�d�O��Q�>����OX�d�OȨ�;�?)��B�YQ�,G�k>,A���.��5[�����d�e̚cj��ȱ�iF{B�U�@��`�����7#��sC��|���wO�bĠz�dE5�z����hO��)��'M�䵋��'j����O6e
'�'BB��ay�F��Rupz�C�#"���'���y2)�"_��3	�\j��F(l�"=�'�?Y)O<��ȘI��NI(��۠�¨P3|��"G�П��	����L��Ο�Χx\�����D�/Τ1�i8r���Ԫ&�6iQQ#^��y9
ϓ���(�%��0҄���^��:�&>f.Z�"e� �>�hr���9FuF|��E��?��.p^��&�2��Bv��bq�O[�'nџ�R��B"�� �hՌ�4�1�/D�<
�D7��a5�X�`8R��p�x�ܴ�?�+O^����i��ʟ\�O6��
'B�8
���_�
rlIK�)M4v.R�'�"&(V�:�ku��4Z乫���:b��"�1L��΀�.p�b�<9E��:-�lE�2��(>i<���C���;2(��I�\�b�H��3z5j3&VE<�<qE�S��)�4m:��'B哖-�$��4�_�e8�ӠΔ 3A$��N�S��yR��%!F�BÐP�x�r��Z�0>q3�x�-%~�Z�)��H�JZJ ���y�#ضp]�6��O���|��� &�?i���?	6�ٽYYҡ�w+F#J���T�P�h`^�V��J�"(��BR&}��7]>��|�ɹ�0�*�����#鞁IZ��I�%w͂DZ�ӑ�&��G�1���`��#rr��G$��f��)��hO�U�j��#�M��\���p��<�p� -�B��N��'� ����V�<��O�LXR��7��*o�hs.�R�'�0"=�\��h�oG�t�čX'y)�|�2�I����	�;<NU9���ԟ(�Iϟ0�I�����O���Sa~����mc�Ț�Iۻc��������BDA��vr��hO������-���U�9�L��N�����s�ޟ;L�
�'��m���ɮbV����Ņ"\:分�Ȥdz��	)kZ\�IП���?��?�/O�!�H�F����N㘥R�"O����hŬG��9S���wŘ��	c�'m���'�ɧyǣF�2
 $�X"'�����W�y�JH%#u�4`���5����N?�y�i��R���xb��QT���:�yR	Nx�� 0�
�N;|��TA�y�� x�ht,� X��	��� �y
� 9���zw80�c)��`��j�"O
p�p�_<��ܑ�L&\@X�b4"OnI��l݇`��[e��]��P"Ob]���ѿ_̄����@��i�"O�4�ԧ0s�j}g˙�G8 �� "O�4Wg<�Z��S�ߵU`  %"O\�biox:D!�IF3
6�a�S"O��`�B+^)����T�x.�4�"O� ��Dc�� ���<Sv�H�"O�ݻ���,t�A�Qk�*��"O�0��f�X�#K�)~��"O
@�fB�>7jrx���Z�&����"O,I��h�;oF�+Ԉ�+�
���"Oh9�h×c�68���4m~^a��"O&48��F6���deB_w�T��"OFx�#�U{`�$b�kȼ@6"OX��&).��+��,oVAkF"O�Ū��ͺJ�4���@CK-q�"O��kE 68�0oB*F&as"O^@���2�D�A�N		3n17"O���nF��bx)���A"O���V��p!�q�Vڕu*u��"O��Gu��豵�U�Jy� Q"O�@+�� 4@L�C�E-bd��"O��aD�>�����%bf^��"O��K�%E1ؑѕ	���h���9D�|����_� b����Z�z r�7D�X�'F� �
�E �g�bXB���5<�O����Y��H�������-�D`�� 6D����R�@�R��s�G3����Y�*�@&%�O��P��D��#�K�(AA�']АU����ʤT����h�9$�̋5���S�L��Q���J[�o�─�@^�gD<�!�1�I�'�D=�%��>��4r�N|b�)� Q��5�7c�4-�@T�oCF�����P�DʓQ�s�B�+k�x���Z��B��4"�b]*p=O|YiٴP�FmXD�O֑���O���<jq;��Jd	+
xz^�i*?�	*8�^�k"O���I�fs��a�Τ8�L��uH޾y&)�aJmӌݛO��<�3���L��s���~���K�I�g;���K�*K����s
�`���9��1H?4�'�>���d�>�`�z�0+�m�1���K����5u���F�2Xf���b�pCgW:^�HH1F�1ȰD�O��j=?��x��8$�"��4F|��(w�ŀzc��c҄�=#���I�q��0k�ľUL�wMT&h��hh3f�'U�t#��ϝT���qC>��'h�d��C���M��Jú���^J}��^>��2�N�S�����(��'rd��L��o~���Dg�i���Ӻ���x�r�aE�� �~]����U���Z#�?d����O��[��u�r�?� ���Ӡ%
%pyy̑�I� �S$I�I��R��GA�61O4c���l��	!�ֳ[v�	v��#�4m2��;��s�a���Yzဂ��2 ��'v�DD�O�%U�fdB6j���ʱp}x�O9��UbG�ц%�a{"O��
l�9ش�#��;��;]*�������k�I�>�.O�BWZ���R�ܞw����b M	�Ȝr�V�_�1�P#X�-��Q"�A�{ʱOlR�ώ���|�ÌS� M�!�J�ܹ&�J1;������w5$ Y�@�*��$ojI�Α�e�T}+b��#p؜�>ɰ��,T*����,�^� ς�L�*��F�R*^<�� ݴV���dg�t
E��O*��O�,+5��!w[���e�ގND��޲c�p��H	����?�=�bkĂ.�^�2ՅMx������i�l��։P����Ƌ0f͘����ʼY��1����4��y��ڜ�Mcb�i�ҥ�&�I&|1x��EW�����eh��>�dG[y��&������]�h�bƏ#Q�z �Vˋ�[�:)g��1�JQ&�tP ,�(cT�� �M/$_jxuæ>�'��<k�C�)W�]��b�-3t��H�ű������)�,�#�x)`0횙K��ORQr�V�H�F8ѰEޒ D���� 7�nD�`b�3M��,�nBp̓.V����$�f��J�a�r5�U��;[vxK�c��Z($�b%Gs؞���	�*$YL���-oj���q�(�4O�]�e���}���G�1�WE�O2H	�צ߻A.��D�"�H�Ӯϛ�sI9wf6�k@��x:�tB�)M&X��n����Ka"0�'�����Gװ�,����72n�m�*̦zdTk�-��[��d����u�I7J��2�+�Z��pH��*��扽( 7MD�t� L��G@Сy 왻�_#}O1rt�y~r��z�)`���+2}	80���'��s����_�h$��  +o:8�[����M��c� �c�po�&n,ᕌV#�ħj�0�͔�\e&�:Q7�y��iF���c�������Ƭr9RTSB��:u�X���:~��5mZ�nB�7�^=}��äV���;"��^w�1�'�RU��N��E���0iR�X�NrX��k�i�
z~�)��Z�ر��\0O�h�"�]Y��I F�>�ëh��x(OV�	�>9"	5\�l7�"6��J��\�>�t`ԥĜ(��'���Ġ[�y�T�C(O"�	�j���"[�,L�.^!9f-Q��̀��e��O
�sL�d���Ҵk�"=ya���d�����P9{o���-J�Wv�iIV���<A"�Oe�扗h��!����$����T
o����`��|8��'����cֺ'�(��w �:(���>��Pd�P��f�yւ�o� �M�GiV��%���_tGd\8�PTx�$���O44�d]:/O�xQ��)u�MZm^#e*��^�誷e(sO���'��U r�M1o
\�2�U6��}�
��l��*�D[5|�����)5>��W̓.��0a��K��}y��R
L��.����w~Z���2e��%O�䣀m�y�vu���Ú{�P�Ȧ�^JX�蒋��Ďn�p}Zw'�Ot��ݘY,vT�W&��w.�ո�.Y�mMD��jW8���z��Lm؞�X,DŞ����-4��x #�:U�Oh7��$j�A�'�6��>�y���?�eHN�ȼX��!@�b��%��SX��{��� �.���D�-�b��`C����Xӓ�C�r6���y�/��eliҤM�>Yu�U�=V�xu�r�I�Q���u�Ś|O~43���u����%�>�;$k(t���nx��[փ߮f�RA��R(��M����n#=�펵 ��&d�2NF�Kbg.P�Y	eB�-¦�"��d�F��?��|��{u�9s�L��E��i(6EW���i�UO�JTI[�G����K��h�Q�J�V����ݴv�t�����S�'�l�h����9Q��4VJ��ʦÏd�l���'~jd�����P��Ǚ"g��d�P vR@1�`Ž n�؎��Y6He h#�1c�V�	��V�-y��ټ`�L(X��C�8�:�"���ēt�>q@q�UKi�0���9erp�>������b��F96<�} W�PV}b�-�ʰ�U��J��r�W,�HOJi{6�϶~����ߠa�4�`oG	-O�����?\:i��Oo�&��C�FXb���B��Ș�[FaV ��xb�-��p>Q�KMuh(�1%�=��2��Q-��'�3��9��p�ˤfrV"�I �0�p�q1!��%{azK��Fۢ]k���P�8&.Š�*"�>��jLoP�c��W�'�♺���4@��`�O�@;ڴ���薯Ll������>B�V�<���!F1i�$Ӹ9J%�Ц�Y}��X�QFт��/��h&
3 ���Ad�(���m�P-�Ech�:L�I+�hO���$#BUĩ�a��?,�n��U�i�tdjƬ�U�����-�O��1AV��u'F/?�O��[��¡#� �Q(ϾOQ"�У"Oh�b5��)?xq��s,.��vӆ�8!�=
��@aa��5���y��d���A��!� =*t�|jp����t�	��li�6\"er��Hk�\QJ^"�lP��W���梗���ɏl��n���MsA!ɁM�6)iI?Y��"V51��|p���'	+���3p�1O�
��t�rtP�C�7g
>}��Z���'��H�F8.OΈz�'E �<�#%]�4����9��J�����IX�'Z��AF�K/*-pE�ڝ\�K�J-|� �H��wU��!F�^N}��|������W-{�1��B۰W@����F,�2�cI��y�Q�ؠ焟2��qD�ʈ������*?�爔�qe�q(�ŝu�		cR�;+��8�s�I�m���@,�Gj1�cD���0=	�h��N5��3"HL���lP%ܜe��IQ"�g3 ��a��5r��<Q_w�H�#M�({�����1r��4W�ҜMPu@�(z}L���ź�1OL���՚Sip$��45�d����D?Md!�����}k�c�:Na�D�٣r	L�/M|�[�!�8>��ם�O�H��
+(��d�o�[�ډ	�ę4./0��F�^?p��}��ܺ'��B�3t��1���4*�|P�Pn�=`t9A�g
3/|����ƒ�{L��C�L!ҠI� F�L]�����1W���S�9π���y����B�f� e>,O( կ"q��J�>v�C0K�34q@�"��Z���@�)�3ў�	]<5He��F	k��i� �-NR�
P�^$u�]�8�H���x2��0�(e�G�A��ԃ����'�H��jZ�XG �)"iƵ7�����O�ArWL¬+�^<	�MB#IXL��o�D��0O��f�,>Q��1�N�"zU�#�&3^9��I�:w��U��*��v�՚i�x�wo�>Y%��C��2|O���cP9�0����\�B-4��e�1ʓ�hO뮁�|� p׀�er���w^�)A��#LO�l���og��I�S�F<�́Ɗ�M� �j�,�0c��X���|�'s��`�M 5Z1�7�HD�֠92�i*��KJ�'�1��	���y2��I ��j1L:��xt�P0ޘ'N��{#���-Hx�C�!7�t�O,mC6�C?"��c���g{мC�)� N�q�GÂ3$�A����(vV�����9g�4-:G��H�ډ`ǓW�����E3v��RA$�(;e�8K%޽Z5a�PU�a|ZcG6���N�2?�T�ڗ�(ۂ����$�>)'M�]⓬?�6������_k�aq�-)�q O�ư<��'Ҹ��~�8��#��F��ۗ�ț�5h�A�8{g��'O�DX�O�c��9�.���t�0����o�~�<��LI2{\d0�D�pƴO��bЁ?|`�haЧ��Uw�(Kb�d�32��t�4�FLk�e�0]�2(؁��@�aՖB�v�Ab��FzR���%*!3e͐�}�`^QE8�9T�q������O���?7���I
ny�vV�~��R#n4�$Ɔ�-w`����p>���=f�̀���
��Yr`F�=p�m��<�T�|��;t��O��a�1&M@�
5B�2�(���4���@�\�ɸ�M3%Bء�F����+e��<C~��G6?9��}��Xa
�����>����B<��6m�8y[�:��މW���bIKm��h�e� 1r��t�S/���"?a��U9Q��KB��>b��ЇOPH}��O2"���Swd�<B��Ǣ���HO�|�2��/��͎e���8��ܷmC�	�8P��R��ܬ3��	b}Ҙ��Kw���	�T��Q.���Nۙ4'ZH���X˰>�'G6,Y #M��F	�6G�;�p%�?��D��ˣ�2,��W��B.Y �
�l��v�)Hf���A	�"�� �f��[2��g<"?)��E$�2'β��:�	�3�U%Z1XI$�n��Ò�4�3ؒ�b�W�
4b��@/H\v,�'-�zC#�w`,x�N�K%t����On1�k��\(��T,Fn����	+j�;��E�q�8[ � FP����OZ���)Ȓ@0���'���Z�ቌA,��	cL��8����[�^��J�pF��$C ?�0�#���7^>�@����2�G8��x��#���zu�;a=e�)�5E>��kЦ��J�zm��t����f]
$�$X�Ů�*��=@��x�M�k� �yܴ8��XA�
I։�MK��� �m���.U��XqG�i��<C�CE�j��b�'GX����13��P�h$0h��q���<7k[(U��V��3��|xP�臉'z��� ��ad|�ȓq���#ơ2�d�EKPUx�Ԇ�Ok&5c�	��*\H)��)�q<���d�0�*%i���>�ٴAO�7/,4�ȓ&f!�u�':���"f68>t��K��h3�C�[j�ٳ���:i%@$�ȓ�	�e�޼v��҃`@7a����ȓ�z1 iƥv\3EA�fA�ȓmҺl��O�+@g��ҕ�V�@~��ȓ$�ћUl��h�Z(:1F	,�6H�ȓ	/�B5������g�� c"�|�ȓ:�nu���\�x7RQʒdB2y~��ȓ[�yX� S�G�F�
#��z���ȓ=I8Y�0N��bǍ-}*����Jò,e*I�*��I�хA�&d����nn��Rӵ l���/eHE����i�SG�#F8乣dۡ[�y�<�Gn�t��4��o�KP������h�<��� ���� �MT�v���&i�<����5òH�Q�E�v ]�e�N�<9�e��L9�4�F&X�J���"QmM`�<�p�Ԅ/p�q0��o9�%��H�<��钍2�5BF'W�4�-�D�B�<!��I�h#à�T
� ҈J}�<Qv�7lW�/����4��K�!�+��	�@��|����hQ/0j!��2��I)w)�I�J� nZ�
U!��V5B[~�YR�K�2��Y	���5�!���V��Vd�5}�8�b+̂d!�Z)lv& ��D2k:�p�JI&'�!�D��7��0荫 '��D�D�)�!�Ğ7JNP�C0팔|��sɖ=�!�dG#�x�!��8�RԹ� e�!�d��v]rM�S)ߞj�N|ۦ
U� �!��ʶ@�
0�[����(����5o!򤈒Bf��X �DJ�D�)q��8B�!�� �����&���i�lϓ2�^�`S"O�8�CA� i ��ɷM���<�� "O�d[�(��9D�9DL��S��ٖ"OV=8�LA5�v`0a7,��1��"OT��^�m#<��W�h��$��"Op��ň
# Z�9���F��%rA"O<i�b�Q��fE#�Ì�.��"O8��5���;����c��#F"O�@Iq�6Q��$��lK6Gh؂"O:� I�aA��b��h�"O*&�X�} �@�sdO�l�FY�@"Oj��w��]�PQ��cI�i���"O �W����<!�W��d���"O,2sLI;L� ���#k�tm�7"Od�s��	 �ʕ�B(�Wz��T"O�A&bT B�;XD���"O�u�@ꀉC�T�#�W\����"O����uV�$��'بHT8#��l�<5H�Y�p ���K'@�𸪇�b�<�V�h��q˔�C,y����la�<� DC#\��ʷ@F�1g�����NB�<I5JU7Ba�4�ph�n��Q96�Rv�<i�皕&� �S6�� @@��z�,Br�<a�ǝ2�R��󉌼J/�A�j�<1p╮:Dl����D���_�<Tŏ�j/����lH3Kܒh����D�<q�ϗl<vh¶hL�w���A�D�<Ѧ �)��P0�S>�δ{��~�<ѐ�N5]W�y���l���@�'�q�<AtG��D\�SïZC���E�<ɢ���.iJ��H�b��u��,�<����R㏊�O�(�PפC��*B��o�~]�U-�����3�B�B�I��PIWJ� ��ѣ���FG�B�%{!�7�3~��e����X!(B�I4x��U#ELɸ���i6L�Pk�B�ɗdT\�F��m��A����Hx�B�)�4��钯ZۤH�,�*Bp�B�I�HM����͓�J�p(X4o�JWdB�ɍE�@9�b��+4��D�7&B�	4,�����o��3[�V(��s7B�I1X6�P	
�>�,eۓ��
n�@B��=$�صR�@˳\�����o/bB�	:*|�yՄ։p���IA5d�B�I�.0��q��ŕ�d ���2�C�p�r���	-3��s�D���C䉸d�8q;�>6n��h��U�7��C�ɼZ(�}j���h�l��u&��V��C�I�3b,=���8G�l�(��Զw�C�'(r@A[�DZ�5d,B��I��C��(Xh<T u,]�Km(��	K'7��C�IH,�U�V�<� ��k�g��C�I������]�Y��	F >_ئC�	#:��l����`����@�_�DB�	*6�z���J�6����Ȗ4~�B�I+c��['K�2a+1�F�{�B�I�<��}p���6$�h֣��O�`B�ɦgr�� ��	�А���_@B�3����wſ"&����A�B�I�A�<��@Ӎl|v��$��3�� ��<E�d�5&�E�`��(H	���g�
;�y�ǐ�	Z\a(�$�;�� �`n��y"
�_��yB�B.S���!���y���5Q��t�� \��`�@����y
� z�Ђ��q��y�B�P�Lؠx�c"O�� ��\XC#	1����U"OĘ�VΊi�,�¡�	i�е�"O޴ ��/o�1f!3l�ِ"OҔ:!N� !9�@j]���ii�"O�4��FA/7��c3� ��A�b"O��Ò�\�%T�3*R��Fx�"Ox��c+R�?�����,v�d�&"ORD���
*��@X4 �fo.t��"O�}�gm�Z	�`�rN��BuX�J�"O6���u&ڌٵ�$"�<��6"O���I�Gnف�fI��ra"OR(8uJ�htd@:s��X�y'"Ox8�a(�e��8I��#�B)P�"Or�bh]��M��n[���E"O�����(t�<�'��eo\�X�"O����)Z�rĊ5.�O(��R"O�Qc�*\(`���l��jܞ)�"O�i�"�]/ɚ)� �
x�`�#���YH<q3��..$�V��epX�p"��t�<�WE���y��hA����p}��'wl`��Ab��(�,S0B1�[�'��I�\g����h��>zZ�R�'�$h���
,(����#1�����'w�tZ��/�2a� F_8o|A��'����g� Zi�w*ֵ7��q�'|>��F,јh��F[�(*�(P	�'.���&*\cx��F�-P[j�z�'c�yђC��a�Pe���,L�H��'�M�.�c��պQ��ad�
�'۔\���W�X�6q`H7*Xh�	�'E�P'_1A,8c𥈲�~��'v��e�"Sd;�F��}�$���'�\��ӈx��B�V~�FB�'\��a����qkB�+qJ敐�'p TJ��,KH��tka�l�
�'�Z(���$2�h��	[�B���'�����c:5B�pJ��X�L\�i��'�u�r`F�O�����AP�9����'X���G� %[�H���ȦI�,|�	�'�����2c�ѹ�߶2�Rњ�'(�U��c��W�z yU�Ҹ)!vd��'8�@2��0)��a��Ȩo�$H��'@�8��I�Yu.M�d�8��P�'���a�ӝF,�T��!�	N{�'�\u�v��0y9,5�����t\��'D�P�D[�Z��eZ��n�����'/�U���_�Q<�"�eE�`��ݑ�'G��1�o6�xA"ţF$�	�'\�k��Ό.늝S�M�yJ�R�'�ܩ�3#,�h����Zf�:���'
�m���P\.H�5���a���'=8��EB������V\x`��' e".�QBM�0)��V��E��'�~L�f�����P/On�m��'|M��D��;,�\���I, r	�'"���L<G~DSR��:.B܁�'��p��E0'❪1��%9�0���'8���U���)t��dPz��'j�d��E$"�"=i1�z�;�*�n�<�e��c�8�B��^�8� �@j�<�ֈ�Aq��<z�H#L�f�<�ڋZ�: z�"V:F�,D���Kd�<飍^��12#k�5o���1
FE�<� b�Ȱ�؉Y�����L\�/ڼ�ɒ"O�ĉ �-�J����f���"Oj�xU-ڡ�aKSF��'hD"OT�B⋚�Ri ��U�X%��*4V�T����Ak:�S� ̄k<�@����B��,*�c�V��R :��W�%�pB䉓!�B��E�]�:���ʳ0�xB�IK�t�2F��	j�xE�	l�VB�ɇTHpE�c�+�p�S�)���JB�![(v��*����z�hڽDH�C�$;{���!	�".�E���t%���'�a�'�lβ�8�*�3|T�'���� %�$!�8�r�mTf�D��'��8s��eϠ�+
U�v��Es�'��9��%�֕k��4f�h�'L��c� K�]��q�žE��Y1�'�����-B�����0b>��	�'�6���#$�� �d��i��2�'�b� ,� D�LT�Ei����'�I��0Z�0�UcX�C�H��'���i�l\-r0U:Ѐ� F%B=��'^zLٱ�ԾK�F�Y��9Y|d{
�'%���ʁ�os	�2��7/B�Z
�'�����z�� 9"�U3\d��'���b��Tc�"��M��..xջ�'Z�B����=�$h�9@���0@J>�y�+� d4�-�S�ַ;�!�4�N��y��u>D�D�,B�z��̡��OV" ��e��D
�n[*� �W�O�<ه��(kJ���H ~�HZ��I�<�5�� Brj51�kV��2,���q�<Q5Ṁr:5���	lRޙ1�G�<��
�  �	��·nY�Ay�.QD�<aa�I�z����)8X�L�<i�o�D�Xa��ćk�^ܙ�R�<H�@���Z� τ�^�Alu�<�fc	�3^^@�J7v{�ԙ���J�<	�e ,��y����CcO�<٦a��#pc �!x��� �C�<A�����ӢC�,n�bpcJC�<�W�P�B��a5�	.�N�څ�~�<���2} �,�uə�<&�="��@�<q�L�Y�z��D�_;0X)ra�p�<A��\�-���¦����q��VR�<�QB!�ueb�鴎�v�<�,�-������.	���L��y"��O���R�ٰz�� p`Aѐ�y��R�l�H��.�Z����$�y�LP��ڠH�")v��0�㙰�y�$��Q��9]Q4�!�h�(�y���"��1qI&C��[d���y������ r3�I��<3D̋��y��
3�٫�#�n@����j��yB�@�*!؈�����5@�&���y"I�U�����	�Y���5NS/�y��B�d�h���gF><ڍS��)�y©H�3x\��đ/5>y��W>�yR�W��L!�E�.��\(Aa;�y�͡@H�Co�$�
�������y���[�UK0BԏP�N���V��y2�\��|%#�	�5aD�80�^��y���y
�)$A�(�|�
�m^��yBg��wW���AA�$��}j .څ�y��s�Tpu�C2�ᘧ��y
� xeP�O<�D𙑋@�>R��"OF�e�	z/FZ�%b:F4�3"O(	�EQ�*ۆ�:�3ez�Q"O��!p�H�B��vtX�B"O�ٹ�*�4W�@��R:6�}C�"O��IOP��C�/Ѳ!����"O�tkDK��=����DNH�q� �j�"O`���+�I9��p2$��FI��#E"O ]31�[ /�F�#5����!#"O�pE#R�z^�tr�S�|��)I"O��i�!ȸ�z���N���i"O0��I��6��]� Jؾj�>�� "On�S��Q�� @�H'-��0"On�8���>z���PvG�vx��B�"O�U�s�
�;v|ITm!R@�� c"O���V�/A����l�D�hи�"O�% Ǯ@9TX�,B4+Sqt��"O��84��ƼEs�c��;�t�&"O&�����?6�X<k�њv��Ɋ�"O�	�ԎfqB�&={rг�"O^$q�][�1�w���^6��2"O�0��Q��p��[ܼB�"O6��T	J�6c`yy�߃pQҹyd"Oxř���3r���&G׸%DD��"O�)I�	���vF��A�Ɓ�P"O@Yd��g��I�D,4�J�Ad"OB�p2�˕/x��)T*}��} "ON�*���� )vp���$����P"O4=���N0�X�Xҡߎ%ĘX�"O(P	�>J�H�� NЎ���"O(�8��C�.�`��O�:�@�C�"O���Q?������(%�\�"O.����{�z�{��(�
��&"O.���Q���]� .� k]j�`"O(���9%�h pc@-�\;�"O:�3��.7�*Uj��A6(��P"OJ��"�4G�B���H�\��"O�e��#�H-�H��*�-�0 �"O��3��F)K��3��N�J��Y��"O$��h˳!�T��]�j�~���"O���oSV��̚Wi��Br"O6tq��Y�{΂{�g
�;Bd8r"O6��$l���N��U� �X �p"O8��%h��5��Y�D��\� `"O�`S�)��\z���.U����"Ol�!��z-��P�a^5-v5:$"O�a��A�R��\3v �-��Xf"O,�k7H��& 1UY21'�kb"OhDђg߀�(1�'���ZH�"O"�J�mF*#3���`GLR�z�"O�D�`e@�?a���F�)<��F"Op�Q��;T̒��A�� !�F"O:ɺ�z�� �q\\� �"O��ƊS�ZC��ф
�wZČ�G"O|������$����E�6���"O��r0��1'xR!0'��y~�+�"O*�����TK�b��+{\mcT"Oh��$�;��W��  gp��"O*��\�K�  	� [, ]Б"O���Sr����N�*2BJ��"O���&-D&&��H�&N�5x=���"OjM�`Q�-Y�M��..���"O&Պ��T(��`'#FH�.%a�"O
Ѳс׊g���E5:����"O� �q)��Ў;�`�Վ��j�����"O�`�k�-*t���D"u8���"O�\tN�!���(��m^��"O�8�Մ��O�j˒�0XZ��6"O�I�O�"�`�a��@;.�u�D"O������~��� G�}����"O��ԩ<���K�e�$vd�i�"O(0�ekZ#���Ɗ�$��{�"OL��/��9H&�p�Z�mC>5#�"O�(��P��|X+���CŊ��w"Ot �v!��, AF����9D��@B<���͐�`��6D���X�\�i�e�WLJ�s�E4D�`���ձ�RKPI��p�ܻ�,4D��i�%E�T!X<���@����0D�hw�(*N�9�S�ێ@�H�.D��q֩��B�����Ӌ-D���(|��ٰv�� " �����&D���2��%kJH�¨B#(�p0F/D���scV4����8q�0˲0D��P&�S�(<1H��/J�� C�9D�l�c���4 7ŕ3I���
��4D�����72~���k�MB�s�4D��r�`؛jHM�U��;U9L�`l D����
��8�Z7&;��)�
<D���h!q}��S�D�3���PH4D������WM���I@<_�R�1D�� CY�aZ0�u�
b,0Q�F.D�8Z��K1yh$9��j���8]ؓo D�P cOMd�i�oA���2D�PdÙ)G�P! �	�Sh"��w!,D��J�\� �r�S�eF3^��!�>D�$P���tÖ��𪞴"��6L<D����*<Pɱd��";��3�9D�0��	�E\\���ɴY7�1��3D���V�ʉ o<d�E�&�>0���0D��Y!ET˖�ơ2m,�R�;D�8�Ɠ%fR\;C�ĩt�i�F�=D��ɇ#�f���2�֝/�*pF�;D��c̌*]2�ҁ��?K�$<��N6D���7G�?��M����gS�5��	!D�X;��َx?f�2q�ҦRY�mÈ D�����LѦ�������KK D����z�b�D�9���"�?D�����߭v�H�0��O"0�A��<D��぀�*W�P-�')��Bl�%B��7D�XZUOE�:${�(Wuun���3D�0��ş~�y�)An�$R�+D��s���&uEl����+ol��(D��s%a��^AA�MË�D;t 'D�����H��(�q��@�$���I&D�@9H�>�nP�*Z~$\�s�#D����꛰{:��i��ϔNm�5�!D����@1)Pr㲯� [H-��&!D�t+��	�? @ ��Ǟ�Q�I1ef>D�Db�͕w�����.^:G��	��;D�$�!�UE��+��N�J�5Z��=D��.��l����m��)6�:D�ؘbhͅiB�������)=D���C�1�>�����v[�t��A;D�|E$��h(�r�O0=i�����+D��a!�>�pգ��N4 ����(D�L(���a�j3m�2U@ n'D����F��T�p4:��K??<n��B,)D�� �젳��r���uB��1UpE"W"Oj����V�Kl��h'#כq�� "Op��W��X�b���J�:�$s7"O�@S��^{`�a���@��̋""O�)��
���3&şF^��V"O�Q�B�Il��`�$ʨ��"O�} ���<���zv$� $݄ 0�"OPBuE@>Vp�Z�NȢqaR"O^�!`�Z5ULԺV� )XԾ�C"OZЊ2�Z0d�4F슖���˔"Ozu+�Cl����3K�<5�:`��"OJ�k`�H�L���C�K��AR�"Oze[Vd�6 �6D�Q�1��q3"OR �rΑ��P);��6�����"O����n���`�1RI��)����"Ov�YAЁHH<� 0��,���"OT�YK�j�{��V�0��0(�"O T�ţS?g���#�9(uUHt"O���dU�L����c�](IC찳t"O@K�D��'�&�ZD�T�7bZi��"O:$��1��\���ֺ=dR�{"O(��R�P�@\,+��ν�Ĕ�"O�P��%˞[�E�I�rb��2�"O�ڰ�+"X�sC%J�)U�ܙ�"OB���I�15�f���#(ֱ+""O4<2S��S�P���Ͻ!�[�"O$�D"D�Q��Uc�$L�+!"Oj��4 ������,V���z�"O��*�
�t)0 �	`��5��"O��1�aE*Uk8�Đ?!�T�zq"OH��V��Bv����D�+�V���"O>��gq}��Č��:=t	)`"OI`���i��m��J���Y��"OЙ�2�����$� oo$$s�"Ov��SÙ^N�UȦA�TZb�b"Of,��2��q` ?FH�5"O�A����](�����گᨱ`"OL���� �PE�GӼ`5"O��G�i�"C j;MU�\:�"O���q�ļ.Z5���2$����1"O����8/ y+QR=6��	p"O��`�ЮK�8��C��2�ԉ"�"Ox��2E�-a�d���eG�m�
�Z�"O��pt��.(� �W�D6,�6Y�f"O���6�]�<�P��ȏ�@e"Op�ă�,xu.�S�G��y����`"O��d��(0	��ㅷ$�F�)T"O��F�r  m¤b�%Rb�+�"Ot�f�J�`�A��Π�N�1&"O�E���prؽ�2��5C��|�$"O<H a�
7-�
3�	, v��R�"O��@1( H�����`d$]*E"O<��!۸$Ύ �Ӈ�bk�p�"OԤ�V��5v�R,8c��"O֠8wS�jp`�!�"/S���"O4���f4(�D`�E�P�W"O�ۡ�$v�@T�l�ĔIu"O��ڄ�O�Dq�,�$	�"O��9��H�9�}�C�]��h��"O��[g�ѳh�|�#P�'�D�[�"Oҕ�qc�O lED	�=����"O�pZUiݠVp�q�˽*��@Q"O�1R�,�+d>XըB�S�n��0�"OΜ��ӛt�v��D�v����"O� Z8�*ł� �R �:��=��"O�\[��P�|S��b��ӤXx�$��"O�1[w�ȧlԅ��'O`x���"Or�ԭ՚i�Rـ�i�	{� ;""O��)$��'g�eiV(Ֆrjh��"Oluh2���<Qv����E6*MR1H%"O��	.��0�ʃ!��-S"O�I�e�D�~��	��E$�$D�$"O��!�h�!(� ���8�FE[6"O��q��$oB�(�%F�pN��"Oh�G�[ ��DE��[N�X"O����I>=���2R��;��(r`"O^�q���A� u�"J� A>@���"O�L+�Ü~+4ɐ�Fԗ?�, �"Or�x��ڇ���[Y��c��9'!�> 0A��@�{J�R�!��}r!�Q�r�2bJE�""
(��#B!�$_4��:f�
'2�K��W>!��Dcj
���ꅯ��!b�I� '!�D؄cD�P���x�nh�ZX!��a;-�2�O�(���ѧ�ҏ!�$Zwg:JCH�0q$|����.!�d2� �#��O�f[���H=Cc!���*=ʊP�.�=9��A�w�֪]P!��0Q�Dbfb��uZ<�խͤ)M!�$ӣ)���Q��>�<���-C�_*!�$���H�ڟj�f��X(!���G⺀#�VR�\b����Fr!�Ah`���#��e7��q�9BZ!�d�+�\�����!S"xi�2�CV!�D�@�	J��ܿA�0����Z<!�Q8�|ဆ�D%C�ð-@0h�!�$�8x{�Vg�ٕ�OH�E���ȓz��k����z���UjX����"O8 (�**8D-��oԚ.�j���"O�и�W�WK4 ��Ψ��"O�Is5A��6��7㌚6���i�"O&�	��
M����7������B"O`xQH�(L9�ҁ��pv�"OV�"��;�>(�#��}F4 �"Od��è*{r���b�ɽv�A��"Ov��S�'a��ȂF�':�8a6"O@ы�gȫ#���1���P��<��"O.���M�B�h�Je�W�D
.���"O���%�+qКy���=j(��"O�mAA�َ1���Z2	G�yd"O�pJ� Ʋ@��V#�})���"O*L�q� p��$�	�I�dQ��"O�ݫ�o����$��5=��X�G"O�<��D��|�P�[��;AuK�"O0Q�1��?�������bP8�y2��z2�P�j�+':\Mk�e�yB�S��l��C枢UY(A��ʤ�y
<V�0UN� T)h)�� �y2$r�,4À�V�>�a/���y��CS@x����;�������y2��} *Y�î̵<���`�І�yB�1���B�2��t�!O��y� �$��K��`��H�nV��y�cA�&���"�^i4��fK���y�Ǖ�D�m�fT�V�Pav���yBcX�A��QW�\5$� ��HD�y���9o�ȩ�K�� 9�C�yB��\0	���Y�$V84�!�H8�y
� <�`!JB��@A�T�(<͈5"OP,K2���)�P��P(g�Ą��"OFh�cƌBU�Թgj!6څ�w"O¼xg��������p4d̃P"O ��z�=�â[�+y<�b"O�w�S�h�֬�2���̴��"Olb6n��u�Vu�T$U�pgd%��"ONݣ����|6�zE�!\U��E"O����:N��
��k���"O���B͇	O�BY��AYn����"O�������b� �E��G"O8�7d�) �b���/R>��A�"O��ZU�:����/��,hx�"O�$��U-�~I�F(��:~�A"O�%�bP;�A�D��8p���`"O��"�,�@�v�2���Y�2���"O����&S�z�yHb�ΰA�"��"O�IB�藣(���Y2݆K��A)d"O���3�ȷ���-�27�P�3"O�+��%R���ṙ�r���"O��Hr�Rrp�#b� �`�""O�`+�$�H�lѣB��mU�P��"O�Q��FL�QD����7,�{E"O��N����#�%2 !�"OnM��cP�L[ Q@��eN��v"O�l2��+O�̹���B�]X>���"Or�(t�S���Ej��HcR"O� huX�6���5�S6/�΍h�"O�1y�	��5/|��������"Oڕb�Px,PRe� ,T�xH�"O���F.��7�8�7���_�1[ "O��KV�CTH��V���0$,a;`"OX<���$W��\H����oR�Q�"O�(�w�]*+Sd�!�f��E	<���"O�8��A�f\\`�@Z&���:�"O~�p"囊YƠ�eo��f����"O~���GGۚ�ALIF���Q"O,�3�ė�v��qi�]P+p"Oj�1CM�0A��
TA�´�B"OP�*�A*��0�R�n1yu"O��W�"6��M8��w�8yAF"O��Eb��>�Jmӄ�T�x����P"O����S�E���ZB�©[�Z(�2"OP��#�V�{:�pU$@��D�y�"O�bW#\=8�&ja�Y8r�H�w"O�mh�ңt��Ĉ�D�M�08�"O�E��Z�x�J#-S�\�q�"O�Lb e��L6��#�a��2L���"O��+b�"o��*Pƍ�{�b�w"O�yh�
(�&�� f@�N�`���"O�����J*��U�Ft�$L9�"O�p��&�(X�C�DO)P�v�2�"O�d��n	Ls�pP ə�0�|%��"O���@~~�#�+)Қ�(E"OZ�R&Nw#@ҡ�E�2�.�"O�ɋ����z/�@��F_�)r��"O�*%m{
L3T�ęH��ɲ"O9@$+Ȳ&%-��e\
��4�"O�HBQ,� \�	� ��,U�h��"O�%����X%�/sj�hg"O8@�Q�ȓ*\�i9��?_7~Q�"Oġ��]��d�i��G.t�Z�"O�eZ4`ξC�N���.��X'"O�±�ֶO�R��PE�!9�m�a"O� ���Z!V40a���Q�"i��ӂ"O����M*�L�9wKBtxC"O��a$1w\���aO�FD���"Od=�ޤeEH��⊶E$�q�"O��0�5n�b���Ō2C��
�"Ol���F��r�����-z�1��"O� zĭѫp%f�2��Ǒ_�8��c"Ov)�CB7GCX�h�hN��N��v"O�E�!E�.� � WBơ.� �a"Oj��j�+��5ӵ��+��|�"OzX�;w�Xe.�B��%(�"O&M�t������!m	<s�l�"O����k�n�2A�ↅ�t��'h,���DLs&�+Q/s���
�' .�j#�G;H�@a�W/�)Q��
�'��)�! � q>80W��~1�a�
�'$h����im&\����Q��"O$����v��F�^
�����"O�I��/�!p\dᩒ�U�Rln�0R"O�q�Ĉ�%�����_�#g�%�"O�2-�,_Z!G/�<bJ�"On	h��O�j'�A�)�=Y��9e"O���Ĕ]M�h���I�>.2�I�"Ov5���S�WBTU�S��} I�"O4\
vG�1F�1 ��d��9[@"O`��#T5p0�d�7.FM��E��"Oj�ppJD�nRXD��*$���"O}��-�����,@�N����"O8wA����ѥ��Е�&"O���̶D���e��nC*\�"O�(�$%1,6��de�&AN4"OdH���)*P�y�$�Tܨ��"O����	.�\X	�E��Ld���"Ob���'�$X��,�P�BJ�4\31"OPY���E�E���V�H�^�U��"Of j�"o|x� DfaH�"O����?M��]�Wπ�K��!�"O�H+Fm�.Yx���m�W�)r0"O,|[�A�I��!��ˆ�5H0�9#"O�*�gP�^mR���P0A����"Oz}��f�wh�+C�6C�E"O�2�і)�`iJ�;/�	zu"O�(����=���p�IO�����"O64	5.i[��~ *��i!�E�	�쨚׫@ h��%��MU�nN!��O�@�@=)�VW���b��Ҋg?!�$J�C�X ��$l�|��AK�	|!��>���bģ٦W��aAƤ�k[!�$Q���8�a�@�!s"L��#nN!�$E-]Ɛ���o��zU�	�	 9!�DJ�~�m��*�"I�� ht!��?]��x�w�ԧo7�����V���������B	i�݈'�E�y��>�@����.Z�6@)rZ�yr&W��61�fN�XؾUc�?�y��'!�<��Bm�M):L!��Ӥ�y�`N6E�
���B�9�̑S,���y�oR c!�=�c1=:��BBK��yb�Ȅa��Q�H�&�XHA�V��yBG�Z`�烒�EfE���y���T��݉�J�w��*�j̎�y�ϙtZ��z��L�uѲ,qWG���y���nw�%�f���d����vD��yR� LSؚ2�baA�
�y
� |٢զ�i�$!RƁ�o�J��"O:�����B��ф��gR��z�"O4�`�ؑ\�J�	�z0X�"O`�8�`�p�F�wH+K��,�"O���aA�0�E��'YBi*"O8��M7�Jի��C@�l"`"Op �`*��F3Fe�&	�u,8���"O�5�`�J�G�B��3�ɺ �H�"O����&���E��R�H���"O�э��E����T�/阙�"O\��r��S��e�r˄%�P��7"O\��_� M�����Ϙ��A�"On=�RN[74 ��"���=p�⬪�"O����e�-���sN¿|�H8��"O�s�$.N��q�w�ت �0�`�"O��j�+�#m�9�K��t�Fd��"O�� ��_�r���
�#3�� V"O��)qR֠�į��B>�|��"O>��C����{U�!��i�!�ĆWJ��n��M#x�H�HF�!��y�$���*����w��7�!�$�-J�����9g�~�����Z�!��jcnm
 (T�O��r��U�=�!�dێf��ʗ��L�z�#�P�!�dT=DZ� Tc�>6��cg���[�!�����w��aG��C��!��x<>̛e,9N4�������!�ڟL���i�M�5&t�� Ӕb!�dY����4���uPīE�B$!�d�n��H����	�0u�b��1N�!���|����&kz��1
3͞\�!�Ѫ_#��Y�IעA���:|�!�$�k	��K���*[���M�n�!�dW�e�H,Ї
E3�Dzu��@�!�B+�~Dq���;	�*Aq'�U�!�dZ�N[����-���e�[ !�[H����-��C��#� �V!��_'|�d5��̞.u�����D��!�ėT*b9���bn�	 3FM:d�!�	@
�`@��kYvȢ�nP3B�!�D��w�� ����?*>B	��lC"n!�Mh�t�'#"W5H5��n߁5c!򤝭�Ñ��3w�U��-�1/r!�D�h���CFBx����AAS!�d_�`:}�7��Se�u��C�xH!�d)*(��J�F�bK��,�!�D���}���[�S����	U�A�!�䆻)Z�X �e�d�ze[t_�p�!����M �ƍ.as���F�,l!��(+��h�G��T|�E�1j!�Ā,R�rA
L<��I�R#�#]K!��?u�ș���\���6H��@E!���-T��rҥ�Vw%���#+%!�#L��r�  4t�Ѳ#�לI!��נ���xWhW5�r�cQk���!�d�	���)�g�� xJ�!�!��XFl�da�%ko���(���!�$��Ty)R�""����Py�O-U�ɇe��F\�!6��,�yR�ɗ�dL�aP=Ü���l���yRc�D8�i�n� �K����ȓQE�<z��]5�Yx���G����ȓ	ʜ�	���[�L�J�egL<�ȓ\l�1�2{��q���H!�e��S�? ���1��o�p�H���2@Mx)"Ot� ���4.�*�Qd�3+G
e�@"O �%��zq�,Q'�b�	�"O���Ѯ,rG2�5��3zĐ�G"O��G�~�U����"ֶ5��"O�,k�U2 ǒ|����m䄁�'��H`�x�<%��/�&�����'"
H3L�h���ɧiVh^H��'�*R�ќY;X!�' ��`j[�'�H���b��e�������Z��<�	�'f��ҫF�{�4����i��=	�'&2�v�=@����p��'M�<Ы�'�x(���ά_���gi�L�b;�'
zЫ�oגs�l��#�@�tXz�'�F���a�,m虚`��? b�|�<��F9�l� BNdE0E$ZB�<�uf8~x8ce�VB�Ф�EC�<�EI͸%�,���}|��
��
U�<yC�@*:\�r�D4S�H��O�<Q���Zld̓��.�R����N�<�4��v�:Ls���o�r�	4oEJ�<!)�5O7B����I9�t�'i|�<A'G�[u~h
r��/H�ڍ1s�R�<A��]c��������(T�T(�w�<��IȌV
~��Ve�g(I�w��h�<�#��-��U��p�z!�ڸ�y���',�9�ƈ�
�&�Y"��y�G�u����O
�����X�y��v	�L�w)ƫ�HUA��D �yB����4�g8:��IU��y"!�:�H؃ԧ�9�d����y�C�r�&	Nʨ*X� �%T?�y��A�=~�RUY�.�(�
R���yH�IS�sr�� 3I���ƌ�yr��7@頀jF�R#bg(2�#B��y���Y��!�E/��Q�84K�N��y+�3a�Z���H�G-�����H��y�h�s�%2pK�7����F��.�y���u�࠹�ם/�����MS;�y��D�Jd4A�\6" �%�`f��y�h�P��0J�dU���c��y"/E�9ј0x4o��Y�9w�G�y"v�@ ��>���@���y�$�;_��`�Ĭ܂0���b�yB��-�Y��/ڄ?��@��m��yb`�{�:H"�&�4�*(ۓ��	�y��ߕQ5�\b��_�y�
=�2G��y�ćqx�2��(p�ő��X;�yRG�#����-�LE(��	���y�ż9a
���H�5�D���O��yB�
�^"A�PN��~G�i6!���yB���Nf^U�!�O�}$�]q4�ť�y2a�Ab��'�|����ע�yB�ߟ1,�Xcv����6	3�&���y⎄�R���@'JE�8��#��y��ެ�F��hIHb���y��e�4�Su(�^,�"��yBmK�]�'��>SŲ!�����y2�Xк�IU@�-K6���e�N�y"ڊ'�N4�f�߮B5J9(t���yr�ЎC����5b\ ����y��5추�
.%Mjp����y��7��6&]��Ή=�y���3&�%
 H�C�`��
�y
� �B��^ú�S3���P2.AS�"OHIb�I̭ra���Ҳ	&v�SE"O�����K���0�A3
�!a�"O����N�A�B���*�jhN}�P"O�����!9rX4b��,_x�9�"O�b��v���A ��h,�E؅"O����r�F��A	���g"O"!��0\�~�t�ҺK\2�b"O� ��]�*]�aZW�)WE؅y "OX�p�¦?�d�۴MRXR�s�"O�,��3g�0�x���=Q�;1"O�X�/��FI��厀�h`Ԁ"O=��GB��I�ON,�A�"OraӰ�L�X��'�C�o>��C"O��q �_u&��FC�1�)q�"O����^JT֥S!Z�OH��"O�JT�E>U�"\�1`ư7urR"O�}Ȇn �}eH�XaA��g��Z�"O���`��%β)#��T�-qzl�"O< 95��/i���zC$W*j�+!"O,p��-ݞ5=�|#�Ez>���"Ojl�b� j:�xY$��Gi@�d"O�(u�0��X �%V�����"O�"CO/?i�Ђ3 K�.�L:�"O�}����Sc�!�T�"O�Q;��ޛbiT����A� ~M��"OpT�׭U}8�9�"�^�^�t��W"OD���ʂ��L��I+d���"O��coR.E2|��T�,��\��"O�MB��V�3@MҲA׳G��B�"OtSDJD0�A��\�"�+�"Oh	xנDvTye�Y���@R"Oʀ����#y2d$+a���䥁�"O�y��2��(xï�<�\��5"O�]�3C 5�X̑�n\��h5"Or�u�� �vnպ-@0[d"OE���!Ivx S�I�`�m�@"Od�vHQ�-o��@��7L��V"O"p�WoI,� �K򂂡v-�l#�"O�ܳA�;w�)+ECK(���"O]��X6}� Q�ȉ��ప"O��C��ΚMSܵ����-a��cR"O���E���|�UGL#_�h��u"O.����0��AقkI/�q$"OF �̽(<�ti
�^9hl�5"O�!��O�9߬U�΍.��H�"O�$����j9��p��1�P!ڂ"O��RV��g}[U,]�"�H�"O��P㇐71� k�1a$:t��"O�y�`+�h�+�GS�$:0�q$"O��S�A�4&��"fH^�+)�l�"O
��RM��eؼ�Y�&2u��S�"OR�P��)k���锌?Kjܠi"O�A�a(��Y)���~N\�ړ"O��T$�7�:9@��q/� c�"O��
�M�,�a�H����2"OR��3�&]hl0�$��(23��R�"O� �3i��s��V 
Mr�bs"ObI`"���:��� Xo�u9�"O��W,���dh�;S.iS"O8�y� #;�Q��'�9Q�Lx�"O��D�P�drؠ� N�>��=���'wў"~"s�ԁ;��l�"o��Gzl`��O��yBȒ�D��d��k[�D9��8�fճ�y
� ���K�Vnd8!`��81��6"O�\:�L�G��D�O��l�S"O�	�E9"!����*(�S�"O�Ȼ�Όwh܉6F�;+)�"O`��wlR�=U�ŸB��g �z@"O��G˰�ܙA7�P  ����Q"O������$�B����l�A"O�M�b W���A�"� n�ĥ!�"OJ��.R<?��V� ��� �y�ϞX>�9wHK@�P���y�f�-c	2`Z�n�YE��cQX��yRk9S�HCGJe���(&��y��/����d��k2���#�y�؆�x0�IM��d���6�y�! 'Y>���D���ON���Vܔ�y��1	�1P�?��H�E
3�y���=��%<	]8�ɍ2�y2�P�<yԌ��iW�w7 =qV���y��=V�;�$�p� �ѕ���y�噜���ꃮñkB^����T"�y�
V�Jޒ���c�,�p�:u�N��yR	��D1|���
��^��S�/�y��M���QyD@A�{sp탳ٖ�y��ō7ƌM
�� �zYr I��y�eͲ3�*]wk�P�w�,�y�84��4�:^�QSf Х�y��ӧ>)��!td�+l���u瑩�y�H� � p�p	��:�|"v���y�
�c�>l[��Ҽ+�0;�H
��yB�E3sE�t�w)�>؊�C@"��y*��G��0k�Ԭ�H����yA��)NrI[R��@��y�-x9X���m����ԛ�A���y2�Į$!R����+G�"qA�$�y�D�*�����H
+EO.Yю��y�L�h�0뚞1��I�G��"�y�N��@ �1A��N�tF�ȓgǯ�y��C�(h��уk�r�jH6����y2L��],�(B�ݡ ���pd���y��8)�\�Cцr�pdᵯQ��y"C�Eyh��G&�%fXU�$+��yb�ϤZ�\�	U�ז4~,�[c���yT$Yi�EI&�1+��<��o[$�y\�b�@���ǖm�ԫ)U�y� �-tF
8`���<2��	@2D���yR'Ыoa��;Q)Y�>I�\�B����yB��kx9*�E�&ˎd���y2��0k0�&��+�p��fG��y���7N�`@���D	8rP�4Î	�y� S����Q����E3�y��?N���K��I��%hq�G8�y�I�B����Ο�$d$<� ��y��D�-�~��L*P��� �́�yrE^�&^���%u��&���yB	��g�P�h��e	�`�&��yBO]�h��G�Z����0�yDʵ?^���R��X~�̚b
5�y����k���2�@P� �r��y��:�V$Xe.[�L7�	�db���y(#"��૖L�<�T:���y2�4�*x��\<J���H3�N��yҍF�?]Ԡ�#�2k�B}H�H�yb�ʰ(GD�
�ǅ�.��%Y����y�mN	22i��&S�Mف��(�y
� �EYu)D�@MY5���~���X�"O�)i�')�����	�n�� V"O䔉#kT�`�0$B"v�Hi{�"Oh83�)L#��ڢ@ۡ,ΰ�c"OZTR&l38��w���Xb�"O
�X��I?>@,dc�`̣ �4�0�"Ov驗�ձMX���sm�=5�� '"OT�&lؘ�٠s,�51��}!'"O�A	��ĸ-�x���E�#�̥٤"Oʄ{�*֡���$�G��r�"O2`��D�Se�i ��L|* ��"Ot�� �6	�H�w
�9k�p��"O��׋Y�Y�5�Ȕq��!rG"O����*
rc�juiЉr��(i�"O��h'�E�Y��9��z��q�"O =�A(�|V�S�`�<{�BL�F"O^}�%#16z<�I�eU
T��\��"OhI��B�
Q�T�'�H�v���"O�0�9>���4�$2"O�¢���Ts���Cց'��:�"Oje�v���}M*!y�bƊ��Rg"OX��hY�C LU��� )�^$q�"Op�r畂5�~��ӁX'-���"O�lkK��Fu���ǅ0�ق�"OҘ�S�������D�SMP�"O�L���
W��0h���W-$��"O�]�CQ�C����sJ�!�,%Bu"O���q�O:�4i1@��Yx�"O�����0eb`�he��z�ZDr�"O~�*�O\�s(��`%Jw��R"O i����n��`���F�UXh��"O�T���q���c"�P���9��"O&%У-Yk��y"�."�h�:�"O�1�0�U8���pFg��X٤"O���$��@FH�!Ćܚ}�j
"O�({���=������Ω�r"Oj%�����`>���ǁ��(��!"O�D�Ri	%m��)8á�%��$�q"O��ʲ�[��H�#G�F�[,^Y�"O@��i[56,#5MԷ"x��"OJu!a�� 
!P5�P얃Tyv���"OD!y��ԕ�`��S-�bm��g"Oе{`�
kP�)����x��X�w"Op�1�m1`�he��DV3O��q�"Or)z`Kؖfy�u��o� �@"O���nU�8p�(��d|��"O���n�JZE�g�>K�y��"O�����[~@�z��1@.l8�"O�(t��6")� ��9[1��y�"O��)�Rd��EOE�ff�Qg"On�Ї��T2�.S8-��ѹ�"O�-z�`W0@?�a��(R�� "O B��8� Xb���>̰�f"O�H���j��z� вIn萕"O,�RD��x����o��9<�uB"O���f��r��!
�oİ@��,`V"O�kG�ПHV+?q��8J%AJ��Py2��8&~1Y�W�T�*���i�<ѢH�� �ĸK��<�>)"��Ky�<a���4A� !���[;�JB�-�}�<yP뀃{�N��VM�}_�UA�g�y�<�ׯ֠ ~��h�3|�!�Њ�y2O�0U8hD
�BN=�r��K���yr�OY�� L�Q��BpɆ��y
� S`�I�d�H4I�
Zj��q"O�����p�  B��*P�^m"O@����V8Lkb9����:M���7"O���Q��8;���+�ңA��8�"O�8j���GN�% �G�+��t��'��Y�tØ�oUP��Jk �A�'-4�KA"�w�|(Za`�2:�2-S
�'�0�2���*�Ak�Eᢽ��'���0��J�X�Ra�e�? ��(��'���`С�-iT�ѫ���wنɹ�'5r@Cf��=G��\"_�L�
�'̼=�Q��4L �1 �ٺ 6�
�'�.`a��M6D�$�w�g��1	�'�^4*�i�\�	��f��"	�'`��z%(F#�97�L
[��8�'V`��L�.sN%`񫀞MZ�i2�'����.{p
A�J�ȱ�'�bpW�G"J��}�e UC`�(
�'�.ś�j�B *�xUf��G��@�	�'(��e�Y>C��	�ܡ=kH��'��"��հ![*���߽1�a	�'��Pd@޴o�R��cJ��/�VU��'#�=x��`-�hP�+�"���'ʈ|�k�t|�+��ߌ4� ���'��Cs�'�M�t�� �	�'��)���j�j�k'�_-}5
(�
�'U��#`�7s�:8���KҀ�c
�'�z)��BN08��Y�HO�Zz�#
�'�ֵ���7t�4J��.@���'峴�׌?ZL���M+ai�'�0фbӐ��}�ܩ@K�5��'�D�q��H�Z5+� #@A�	j�'ߜ\!ѭA�dK�P���EM�q�'��e  (E	3����!�B��,�	�'�(`��h�����7PJ��%"D����"�q� lr��ܽ�~$K"i5D�|��Ј�� �셌U���ƅ2D��v���9bSFÀf�>l#�$D��G'�~�K� �3U���s�$D��J�D�o�����۹h���3
$D�� ��ڧ	u6ɺ���:L�5���-D�(2�۶~�<���ԃqnh*�(D���?WD03��8=�ŠwE:D��`ѡ(h �֢׿*��� ��$D�@�@e
v������	mxБ��!D����ώhŀ�eA#]$Ft��e5D������A]<+T�i�>D��&5D�HI��b�A�):��U@��L�C�IKְI��N�C����v�K�6��C�ɻsR��"]�S�F���V���B�ɫ4��4[!�[o6麦"U�A?vB�I�*��ΐ�=��`�7H��	�'º;�.�U�;�X�z�f�	�'?�`S1C\�K�mD������'����͎�����)�,m��'������zÞ1����˖$��'l�D�E�U-��4a����@�"�'�a�p�J�0���y/F�
�'�X)�fE�5n��@/s�R5��'��5;"`����uj�.�-?yF���'=hy�#��+��1s"$�`¾$��'}�	��	�1�H�$�	�@"2T�'�BhhVS��@�;TE@�>�$\��'��{Rn���`)����7�Z���� ��2+�
0Xa !3X\����"O�@�1l�*J�%(���(E���1"OR��$D�*��`΅�E+,{"OL��a���Q���F�6V&Ƭ�"O��SF�H��)R ��!���"O��D"1!��Q ���	�"��"O*�X��չ1q�L�a�Y=2��Ę4"OT\��[�|�v�0�K��y{��3�"O�-�PL/1':�I6��e˖���"Oz�2"'B�zm�T00�H,3��x�"O�q����>H����c�X;n�Bœ�"OV̪럞2�m�畁/ʚU
�"O�y�B��Z�n��B��O�m�c"O&��k��
����+]��d��d"O\$æ$ź6�z���T 
y�	i"O�d��%�t;X4	�I0Kc����"OnY�EEڣ5��*.�7t\�s%"O��i��t:��C��= =v���"OJ�sԩ�~�~��(D'�TT��"O\4�剙�nO�d��@�	iv��!"OmO�ӊᛰ�I�] �؂"O Yقő�w�=���H�J�Z�!��Z0!v��b��|���ӣ z1!�#cVQp�3" `�6�ܬ*5!�d��<c Y`��?-R�'̚>/.!��]�T�w��4�`)�Ez !�DT�o��� bhɍ7�B��#��g�!�^ %� �Η�+�>�C��8!��X&~:С�v����8�7$h!���$F~D����x���'�R� !�DW8-�n��"�A�S�M���\
U�!��F](
\�I��e9�)�-b!�d� ,���sJ\ T򘩶�� �!��U������'�jD#s��7�!�D%RH���o�^������W�I�!����;�"us"�@�A�c�!��Φ&��'�.'�|��ZU�!�DӜk�|�	��]��I�͡
L!���V��:�Qs���&
!��\��)�n�%z�|����>^�!� �0h����&Abt������/�!��(o.�1�H�?unR��8:!�#5߀�������$�ă:"!�D_`~��� �:�T�
�`үd!�DH�5l͡�.�uض��!�&P�!��6D�����fS�eҖ!�3/T�!�$�t� =�ᮎ=��8�-�5�!�@�'��(Zs��P�>�#Q̆�F�!��Գ�P�i[-x|渪��F�+�!��S�4\jd�uEqg����� Z�!�D��J� ���G�RSn�C���x�!�$)��x��Щ0�x��Q�>p!�WE�JW͝"~�:I##��X!�S�k���R���7m�m�% 1&N!�?(,��ϒ�^����..i�!�E.!�n���Θ�}�n��w��\�!���;��R �*�����K�!�DեXi<�"#l�(E���s��9�!�����Qs#�

��P�"�6n!�*X�2�8��ހq�r1�ƭMj!򤎵}R `�*k��A���I�DP!�DT�,�x�hR���4�q�F�J3!�d���UYC�1�V`��Y�}-!�$Z9q�vM0�o�=-����l�'$�O6O�|� THu`C=)�,x�WA�n%��"OhQ{�J
u9��fV�S���;�"O�}��ۍD�L,��F!9�F��"O��{��T�th��;Ud��j'"Ol ��gN�V��d򵨊�P7(k"O�����^;��z��36�+�"O9	�k�(j�B@��FFXH�]q�"Ott�GѸ6hQ�@e B�Ҵ��"O�%z2�F5}?�\���We���T"O%�! �n��0a�)-Vb�P�"O�@��*.��mZ�N�
DJH]�2"O��jC�I�T�օ��͑&aJ>��G"O��aN� 2��m����I 鲵"O:�a`/`����Z�xj�B"O�4��DdS��
ˎ��!pL5D��-��2K�u2d�D����}��lXЮ8��I��,:f}L��P*O2x
���Q�^<6(�4�Pc.D�� SN�F$Z����ɍ`�ʧ�+|Obb��3�-�C蜸�B�HAC�u�S�%D��K")�+�NDc3儨R��xڢ�#D�dBM�'R�V��JU \c��{�� D�,�M"�\8��c�4]����?D�p�i�Z��@�C50Y*��s+D�0A`���0$sG��:UX�� *D���	Q���h���5%4R��(D�LӶ��:�� sU�JS�zm�f�(D��'���a�Ġ�󁞭F�x!5�>ɍy�OwbE ���pW���V�WFnL��'�@
eeW�P�~�A�-�c7�`�M<��.Lv�Hڳ
x��k��H.bض%�<���~Bٴ-ڨq�w͕)Y�� 
%�,�R��ȓ.>Vܫ���]����êT��F~����H�p�Y�7 �}��-Z����r"OR�H ��-Wl�:�dB3%�ԥ��8Op�=E�t�E���R���)G�$]�7eL��y�cY�2��b��#K����&
��y�^ l��c���wf����>IO�P�����j)6�th�
LT���n]z������������v#�@K���!�ɅQ'���l 
������W)'!�d��U��j>~>8��ևw&�	a�0�<��
�29��3�A^z�!�xC�	9@�h���]b"(�h͖��C�J�,������dCL1:��C�Ʉ=����A=7j���S%��}��EzR���$,W�C'BZ��?a�z�"G=D�dr7�H�v�|�s�D�a0���Ojt��5��9)teT`��D`T�{���ȓU�t�.1�\uIҮK�uS>І����~r_Bc��;�(��)�@��6A��y��y���i��W�Sn���tb�:��O&pF��H�W�d��S*��Dl:��K��y�`�6K�f�5������,�)�y¤�5u&����=j��"�ō���!�O48���9Tl*�h�!O�*S�!���'˓|�f�SEzۊ%䆋�"�����6�k0��!~�q��։tX:��'u1O���I]�;�"U���D�2���!\S�a~�Y� n��T5�p�aN-Uh98al�c�<qd@�i����A���]t�<�3�A�Py����8��Ӡ�F�<�Gn����dj�6E`��MŦ}G{���i�0
���.S���0�W�p��ɸ��� ��b��0����s��^�Dq@d"O���n�"=CB0�a 
Ǆ��G"O�<갇��dD����z���r"OL4�$�*l��Z�#E�r�q�8D��X���{�Ԡh�m�>��]j��1D����g8Z`M���B�����)5,Ov�<�" ɐPߦ� ��V�J�Z�)U��hh<�aoGD��}cU�,W�i�fH�y�BemRa˳��=QQ��$��y2)�:m��0��G!6�<j��@(�yR��/)����^a]�%f��#eԱE{bS��F���݊c�X�A�(�B�i�GZ��yb�]�A��h"�$��h�7�O	���l̓��s�S�=�t}9$  \�Nyh�(߂$z�C��d�2��L� e�2���:9B�C��:�hi�큲�hp��C���C�	h	�T�F�J�<|I׋H8O�>B�I-�AA�G�<F+�f�*r��C�	�'u�� ����J��bb y��B�I� e�9���L>]D<iz�G���"˓�0?�i�aeJ�Z���_o�X��I�<	t$��m����PAQ"~��]{#��F�<9U��/$1#Ӡӂ��2d�@�<����p�`�#1�@�iO*;dM�S�<���q��WyڴZ�m�L�<I�ɩ8�I[䥞� T
�ppǈa�<aUD�J�މ��\� ݘ�`�<1�W��j@��?Bf��`S�MC�<1�/C(i[�Y�5cԽeO��Q���|�<�D��-vĜ����<e�8��2�P�'`Q?�{L.�<�R��1W��}``�&D��Pqꋰ\P�\� ƕ��
��c �O�˓XHzɲqa]�Fq��:sdߙ9�΄��O�|�3Yj6�	�I�)Ry0T�xB�'����)�'XT�p�!���$(�'(����M�rM�����W���
�'}�b5��N��Qc ��^ˠ��
ϓ�Ox��c"ަ *.$��H
9��!Pe"O�XG+ *�fа ��+]�iŘ|�d&�SܧC�LhZ�9%nd �[a����'��~R�Ό6`r���%1�dP��D����!?�5�z~ҁƋV~X!�㏀?��D��%�y��0޶	K��jY��[p(���(O4��dFUL�a�ƖA�RE���6Q�!�d�k���cuǂ4��X�d`�#�!��ֺC��!W�2Bqꀲ�I�y�!��/*9���M*AB<�jĩ˄*�!��N2}/���G[�D}��	R'	���D����$m������Jd�}�D��2�y©C�#Z�<�%�%B��K���6�y�Ɂ#.��R��
1r!���֋�y���l�°u�H�1�HU�6��'�y��T����n��@����y���N{.�I0+KgW�h2P��y�+�K�x�"�(Y� }�W τ�y�,G�?'�����M'*��V,��y�l��=l��IW�s?@�����yr*O�;^0|K�+�5i��%�B���y�1_R`�sMүkʮ59��R��y�X�AJ�u�4d��Ű�
Z��yRHH�&ؔQ%F�_����(�y".�=c�V�)�O�j�31IB�y��+���AA�U>\��ݡ�KO��y�[7NQ<Ѡ�"Ui ��T�E&�y
� �H&��\��R����"O�$A>^v��#K��c�Ȁ'"OV����Ƞ~�Q�ЕQM\�Q�"O<����h�(*�z7�,�"O�}�w��Q7z,a%J�(,�(��"O�!dk�!k���I�F���"O69A���x0����4��"O�`f��:Lj�1J� G�ز�"OH"N˞Y5���O�0JR��Á"O��������5n��3��"O�|���
2�`�T��$ �$B�"Oxaxg�ي+���9�"��{Z"xq�"O���hȎ[�8ړ�S>��xz�"O�y�  @{��Y��
]y>$�"O�9�rn͎'�P}"D��#
��9"O��*,�n�j<�mY�8�|3"Ob�A�/���&ǌ	j�f���"OjD�FGZ=h}.QX�LҢ����"OX�镎9S`�u�O5c����"Ohi�Hɘ{�vT��i��}��E��"OPHd�W��R
���L��"O �4�	/�� 2I�����U"O��+��C�=p�unO�^�T���'�Pa�ĞXL�%�e�$�����N�U�D[�'�x�#W�ۧ6&Af��B{̹*�'+^]b�#W	+�4�ef�-a����'P�h�挒� ���7J�qؘ#�'|.tB��j��!`�VZl�
�'�p5�� ��m��@�tiU�e��Z
�'2>�	�f�.��!Jf@�UG���	�'�@T��g.�^�"�A|P3	�'O�}S���d��"��Z�ze�ܡ�'�B�`Eեv%b,iaԕt ��	�'��P8f́�F�91!ם=��hi
�'�j(Y��%d�r1"A�7v���'����Ç�7�!�)/#�l��'�DMK����B��U1 g��A�Rp��'L(�B3	2^�!�'�O/;��(��'Y�}3�h�� z ��h�A��]X	�'��}�@�	ys��I�IDM����',maFMR��v�� <Ǹ��'F<��C]�;��d(���9l͓�'��	b��P��F�a��K�C�ā��'!t�)g�V�f>H@R2eY�Б��'2r ����t_��H�D�6P���ʓΠ�{j\�H�Tu��m�{�ȡ�ȓw��GOT@X��Y�!� ��`
� JC*> !X�
PL��ȓ1B�кR�U�a}
�����34�T��&�j�9�+��.���k�������Ȩ�p��/Bk�!_�[����ȓOV�m�7Mպ��i�Bk��k����x�1��7�|��䛶E�Ąȓ��@��[,Y &QHP�Ȳ�^݄ȓvxd�H'%���HQ�[����t �����1"rJİ�o-8�FTCb��x>D3����)�����Жk���" �(� ei6D��q�㞕u
Z�e�L-C��)�O�]I��PU��*��P~�P���b�ԭ�*�04�����mؾ'�����`��`k��[�A�iK� �4��QF�� �4��D@�u��%��M�#:1���B"O�-�/G�U.���sh�Sa"O<XU�̖n%�L�B`̚J�����"OP��dլW?Vh�a��cC���"O� zQ��i:�\#�ǉ{��u
"O��.�pN�Y���{���!#"OL��!��`~�dK��σB�#U"O�-�!iB���4�%�^>7����R"O��Yq�ʵoKdQ�w�*�H�x�"O�|ro�j�Z���]�q�Aa"O�P1&�.$V۷Фd	��i�"O�=H�E��F,�d[���^���"O�����>4����Q�O�pٰ"OƄa��B�
�|�!W�3�E
d"O�]C��V�`��I��DZ;&�]��"O�T�F�k��Ey)��|��`�U"O>��N�m�4�rCKJ�|s�l��"O����kC���%j��e�,�;E"O��a�!��}無0�j�*v��3D"O�$�Ү�c[��:s�PD� b"O���%!̊yX�����M�7���"O�I$�-Xx�<aR�A4P�!$"O�̈�l�W�l�
'�I+*#��`�"O2)c�%�*3�(��](���'"O�"%A��v�.�8c�D �pC2"O����M/s��z�.@�>� 2"O��r��0n��<ۀ�.|��xW"O��R$�Q��z+�Ə�U�j�+�"OTA�B+�%r"2+G00<t�Q"O��p�k��H��$�qEK<U���"O�ő$n�_m�ܺ҄
�}�i��'�nE�EǑ�rz�l��ԔB�x8�
�'�nu�Ue@�<�j����1�j�i	�'n�a�)�24��EH��'$,�"�'(���T	��!�Cbh<���'��`�Q�D\Q���0+�ѩ�'�8Y570�8a�X9#؊���'�T`IG+��Z�oBL��`�]e�<�S�ɲE���{5���(�Ƽ���d�<�����֑�í� 2��C� i�<qa�*v�ʱ�ѬX)_���c��g�<A!$����)@��[mԔcg��E�<�Bȷ�T�X�CW i~���PB�<��O Y{�-�#�B�%������K�<YU#�?xF��W'�'���h�<Q«�>K��I��mR��DE��P�<)U�0�H�:@�5S����t�<!�f^h@�X(��]I	Sq�<AtCĩ6���VB��yݬ�PFnLq�<AC*�|��IËT���уn�<yàZ�f�t�$#PRpe���TQ�<���I@���F�ـ8�\��c�R�<q$&4l6H�Ka'��vDXȘ`��H�'��x4_t�O:P}§�?Z@p� &L�4�p@	�'[��[���	}6F��+� ��e��E�>t|���GC$}�[Ģ�Ր|y@�/C��![��-D�|kD��A6
uQ���Ps���7��7Fծ�$#P7�q%�?LO}����O���@ Ԛ�N��p�'�i8Pʍ�f"�U�s��n�F�QN[�P����c�!jv��2O,���4M��� _%K������%O����*�nZ�Q�D�1�S�h���·��K��9A@���VC�	#o+n��&�%(�p�h!�^*rn.)�6��Ng�A��h�
��:�F2�3}�'\�i����L�2K��y*�i���Px�O4]�9ӵa����Go~iL�ɕ`�^��ax�<P���'��a)Q֯Jl�ŉ��w���yÓ;�xEBC���cwG��Y���8e-G5ú5��) ?|ۃ�R�pB�ɋA:dй�1FiИi�J�-j�5��qf�+a�� �1�Q}�Yi3�ZܧtC�p���UO)���,���B���S�? �``� װz^M!5Y�A*�i@�Pn9�'�ԖP�!)ԂN5�O� 0[B�>�7�6L���pp�V�K	P����Ty��h"�)C�(�k�0���z�!G�;"�'��>Ri(-��	�f���>�p<a��֫T8�@��'t�y��+�F�'Xl�r�qb�(����E0E��&��ZV㚙.%> ��A�(��K�(�$��Z%�(�B��S�e�� a0l �5#�$�4�_�(/������ 
���$D*,����/�]��@�Q��yr
	
%1ЉzBA�Ud��(`/�31����c*#��CFH�� kK?a�j��6X���j��H�͠ãC�-�t��$��6�!CB6n��w@1[���hج!=8\��!�}o8�e�|������i�!��F3_��'����AR�<�m�8|��P��d�,�{�e	�X�,�C��&��".V��4P�6jƶA�. �D���`7�X�K�N��vh�f_� ��I�����W�]�|>&-K�
_$��>s�\ţ�		A�JԊP�
�xL���n�>���@d�.���bk ���:D(5l4A��M0�'��@b��"n��!���a3$�:�H[�(ۆC�| y���L���v�I�`��e8T�5�����
}�,.:��uFĚS$�v�E�Y�a���v�f�X��8<�YB͇�dIJc�o��PN��s"�`J�0%��0eDZ�2�i"�gOF�'��d8ƣ�6EO��P�իM�ph�����Q��
S�8���A�+�%�Q�Ӻ	�NݢD�-��䰃��3b2�۠��O_v��,N�8�X9Gb&��;!rY��-&�@�懙2��$Q9�� k��ۜc�ڽ��
O�k𫈲J��	v,�b*���6I�6�8y[7�R�U�A2�H��i�L`��	5xJ≡��D)Bq҅����=vSZd�D_�oTZ�z���O���Sw�ŶE���&��Awޝ���
�p\D�]8ɼ���K�;g��u�5�cD��$Q;ή���A�8zq�)D�|CJ٩�ΪO�H��7H�N4���U,������5`E�ԉ1zNP�'�$	R����R�2,s���ƺ����h]XQ�@,@�DV$����N��yCᢂ�R�n(��!_�S���ٴ!4�Q�G1=��@Un��2��EG�$�,�f5���J=F����W�M���$��)�
-��0�d��k�5^�xTҢoг�M�#6O~8��(;�^A������q� r�d�)��?�OT��eJ��RF(�5[x�
���J|��LB�d�0\)�u��O���( 
��"MJ�f��N��.����L����B�|����<-*ĺ���'D0��z�'А|j9x�+�l}2eU"<���C�K�Xxa8�ҡ\H���<��ɳ��]A0L�3"/(�饯��]��?Y6��yĐ�� �=�hPyf��!`�B%�U,��C����a놣m�"�򉕡X�lC��ڪ�t�^�tF"�6yq���@ ��S�@N���䚃C�l`�/�<*`�#���vB�x�(F��� ��ƻb��9sPL
OG�Pb�O��]��̂���Ԅ��(24E,iK�ly��K�{�b���AU��0��$Ot �p�W�Ƹ9X�YP�CfC�tY��K�x�r��1�~i�R��=4'P(�I��r�&5�Oze�2+T)i>p�X3%��3�l��q��sbR��f�1[�	B#���:�A�Ɣ�j9~�`C�]�0�d��ᛟ<P�l��^�K2�F�::P�WE)OZ�ZQ�I�#��p�G^�$�<�a`�@y
1��kQ�	�D3�+��!xdG� \���.
�@�j ��<���%��Q$ H��ѯZ�OL� ���]+�X���>s�
��jŃ���J�|6���˱u�9�g�ܤB�<�f�$r�B�	yu�HxS�ptvbƁ�R���w�7�$=17GF"`СQ��^�y�l8#�ғqu�\�S��� �l�� �� !t,����&��C�I%e�0B5�Co  KíN+?��y
fhB�Q�*4�f�27����C�?�)�2�ē"zHƅʋr�k��A�H]"����:#v@�/�l� �	r/ߪ��_��VSh�2�A��(���ݦ02adL;%m|�D�P� �ɇ�	�"g�5Q�+�y�������lP�E�<`z�x��C�El��҉0D��Vj�. ��I���h��,�Q�0}��}�Li�c  U�F��E$�'�~�y�I�����w*�,����\��h{4#��{�^�1�Z0��u���E7jD�w=O�Y�AcPm�g�I�^�����Γ1����ʁ6�0B��!tal�@�QM���%w���H7FA��PI��K���1�I�1�t#'@.W),P�ȓ"���92�[;#��U0ௐ�I�,!�ȓ7�2�p��h)�HlS&tD���b��4$�BR$���R'`��"O�h��K�p=����$#����p"Oj񡒏�~�!Ò�D�}��4�A"O�-�����H�A�J���(�"O<�������(צ�RqL)3�"O�]#G�8wZ�@�Ȁfv,xh�"O|��O"&�C&C�m�|��"O� Yi׋Y(7붕P��W(��� "O����G�4XL;���Y��W"O���,h�D̩�� <\�p�"O.�i�d�B^��rM��{]��"Ora��HؽZ,��b �P�{�"O��᳃^ g�Y$ˆ� ���"O0�k���+j��g�g�[�"O���j���qLfA �8�"O���e�B�)�d@�[�dB�"O�D�v&7F
��PA��,�!�s"O��c�-�ց��I�D��c"O���f韚8H�4��2֠|`�"O~�� �D�D �"b_�L��q��"O�2�h@�b���
�B�>��t"O$)jRd q\��,��Zыt"O�]�K�>c�p�YDJJbyL�"O���!Nª,������4olt
�"OR�	�(��)��``��-}Q�Ȃ�"O�� �3 ����ԓGd�2�"O��u���q��`�̖rJC�"O:E#���-t�����P�� �m�!�D׉+8��؅EVS�0��$/��o�!���:Dx:���#[+]f���w	��!�Dòi�0�iuD
+^T�T����xf!�dӤq�����F�1n���{F왍3W!�d�,^���Q&O$�.��q*�&M!�dB!`f�Q�KE0k�Z���HV,U.!�$	�_n$�l�$E[8PRРǪ9!�D��GA�B��[>
����]�o!�$N�Ng�Q�l""|2g7�!�6B��U�D!\�g�J�7@O�D�!�$E�k��8�`(È�<���7�!򤙷oݦ��`-X;S���@J3�!򄉰F�q��CQ<X���Ky�!�D��J�L��ɛr]�1-��z�!��<�leX3m�#�����ʯx�!�� �����!�6)Ѵ"O�Ųre���T����<��`3b"O:�&Ȝ4H��+����t����5"O���h^��\�;$.ʿr�	A�"O���	@�<��0j��;+~ �"O*I���C��%�U��X�"O�Yt��>����c�`�\P�"O�����E?A�
���Ч-Ѹ �"O(��0(�=�LIC�Y��"O���ӥe@A�C��1Ku@!)2"O���m��\U�q����`vX�a�"OfU�ā|�bh�vA	�w_�ġ�"Oڜ���ȕhO��yI��*KX};4"O��x�	R������<&:��4"O����aV)p9�dJ���!N*(��a"O�80&�G;�l���p�0}�g"O�DYHf��dy���8O��Xd"O �y�i��scH�A�n�����G"O����:*����n�$�$"O y��Дp�ȄnE�Z�Ҕ"O��e`�$(:N1ӠG%��U�'"O�p#�� +���C%^-.��ᡕ"O��d�S�XT�V�Ė^���`"O�8#7F)Z6�����	J�iC�"O��q��F�]"�QpJ��0�)��"O���t�������R�	�z�c"O��	���&z� 2C@df���"O^�rѝCژ	�B?]k^�٢"O� �Ċ3�\E�%�v�W�lN��U"O2�	��Q�E���X�A�d��|��"O�}*#��^�0���V�� �"OJ��3@<(�D�������1�G"O@�7��h�81R'E�~��C!"OuBPL;BS��wG�t���"O��3�/B*�x��2e	�)x��"O`@�q#Z�}D(:�圷e��@y�"Of�C��#j�4! FD�v��k2"O�����01��H�ߵ�r)��"O� E�ڋ=�4�KB&�&�0"O�=�g*��*t����p�ʵ�"O����]�H@rGU!�\(�'"O����U�Jb������@f6��U"O��h2��Hp�a��&ڀ7�D �T"OZ�q�'� �2S�$]�xH�Ŋw"O�Mh�Q��$�c�፹�xg"O�0!�<�S۫.��i "O5#'ʟ$b2�3��]�:��Y��"O����W�.�T�E�-���"O>M#�'���^�k�BQUhN$p�"O�	��YM��(��V~W��S"O��[���P�!���
J$v"O�|a�N�3�D�p�ٳc7P)9T"O2E�wk;�P`��$�vG��q#"O�(�b��9b@b�1&�(S@"OL4ڲ�(8΍�C �W.X�I "O�ꓪ�>IK̽@կ�%N}�3�"O��)���>��z�-�)�< �"O��gb̓~X���u&хV��p�"OF���O��d9����'2E� �"O@�I�씛d&���B�U�JL�)�"O� 3�\=�|%q�l]6o��sB"O�Z�)P�\<�(0DԣxH.Җ"Ot�`� U�"�0 !F�61�c"O*�I���e�Y�� ��I�̜Y�"O~1���E�&J��cE�Er�PҢ"Op���ʌ�$�@�A���b��a"O|P�\�7��Q ��@7a{�5pf"O��XT���FP6I` �ġ|��#w"O����C��>�}� 肗/�&��"O~��
�9n��j�����"O`��#��]�=z1�^Z�D�A"O��3�JB�]���1F�R?u4�:�"O��ВN>\���F*GRZ���"O����iӑfd��J2]ty�c"OT(j���
��S���b���h�"O0MPv��Pƌ�hR$O��k�"O��r���y;��%��i��в"O��
0����
9���z���@�"O�8���ʨ_d@uQ6�0f����"O���w���!πEc4� 
)��肰"O�Āf�ƛ>�ޔcD�_3�Ԕ8�"O��Т&C�w��(4']�D�a2�"O�Aj1N�{oD�9�L�B��"!�D]�uw�r�fF\b��j�!�D�&�F�c�-�#��С�iR%C@!�$�87�H�+�1L1�qU���!�D=F,	f���v,�@ ��P�L�!���]���@K�m'��!�D�	U����H�� n�{!���%��ڵ�s
�\��T;a`!�$Ѫ?�\�4��<Q��x��bR,¡�D��`���A%P�vMN!S$bĜ����0@Y�V 1��)� ��:�. `��F�P�<�r�'3&!#�G,2����O�؋��ܲ�L��R/�K&|�Q�"O�8���PNv-��yp��T�0��`�1_0�E�.������ak�AA \yjR��p�"O^��S��z��e�����L��ŋ?���x�R��(@����'��i���u;@u24DD!LX�
������'E�!9��ET�"���;t�
I�f8ڳA	�[He2r�'��(�щ�;8̶o��,�d�)���N��ؐ�s�>\)��-�]Zb�ͦh'$0��LX�(�H1�"�k�<�a�S;!X�&g�{8̡���j?��H�=�H髱�'2!X���S(]d��I����+t���U �4�:C�I�Z�U��"Z)~�,�`�&Fx�!�%��$+)���A&Z�4�Nz����Ua.�zrO�+\!R��5'�~��Mh�@�a���;P�\���fӇX~��K!-�1Vd�{e�ĺ
m6y��O��
׊҉t�d&>�3cL�ّBк2P�Yh�f���Q�0�!�%�S�EZBn�j�O���p#�-.3Ta�C�ɤ(�򤰟' ��r�;��\��h/,O��(#�7{+��!�ǝ�9̬���O��s�m�9�.����&e�j����������`ZPZ��Ƙ�� $��o���rh���(����(<9*��th���7Y�<
���e���+� ^z�Qa�%� 'C�(v�K:sf 𥧝4^�RRdMӼ��j��F߾���
p�X��g����3�h��5݉P�����F�#8��a㥎]�ޅ()�Hb��Cl�5X�0���
V���´�[";��Q+O0@�I�l�^�qEƃ<y�`lZ�I'L�"�&Ԛ	��}������a��a�V�NH頭�~u�I�FM�'K�S��E�\}��g6i�nt���ʈQ��Y8$��7vED� �K��pr�	<D��1I�c�/���ɢBU/a�+t��U8���2�ݟ..^�¢��%���nچ����ď�(-t8a	��(�����5 ����c_%u��a���-Ex|[0 ʼ)2�]R'	�/����DǷ��Ӓ�:�ew5�!���>��83��Z.�H�'��9"$(��aT��PI�*`F4�����00�8f��d�����)
E@8k�I�0f[��8��ʩfK.��D�<iӮ�J��h��B°	�ؠ��a�'*"1�2���\ؒc�'0�Ĉ�t�G��PJT�B��l�P� �^�`�x�N�&C�08P-��SB<��H&�'��mj6XK�q��ˈ�`g�]�'$��V���$���-H�f��q{�!�:l�r�n�3�y��5|�|�[�K���Y��
+Ī}��Ox����RתԁrGؕ	z6EX�ΉI��.z�y��!�����*m^�\�C,J�
�	��<�҅9�+G�KR\R�l��ia&��#�'�ڝ6�єd�UHs&+����;t�E�'�P�H^+�ƕ�eȋ1q�4�AC�T�]��-�2\� QE�_��u�R��?( ���'2�Ap�fi
� �r���b�LIF�I�oɜ?��Y6�z�������J���3(_fl��7M�	�0�d�	Q!��!B,wR��7�
�>���U)��#~��tU
a��X��k\!+���pb�.HqR�x��0qS������(/B���bQ
E '�'�M��bQ/)�� ��%*E2��)'�"��
$F�|2 `�%@�q�2--���d�8az�ww�E��K�38�1Q��F0+�R�P�'u�U�0�\�F�2�l)�8,[r`x{@`�UjU.w�ޭZ@��3 < �G��_�H�
׌�(�40�O���v�K�֐�c!��=#�z7�'?(Hk�N=�,��Gh8-9�y��Ɯ
*�l�e�W8<i�@h�"ĺKbҕ�Pb^)b��#Fȅ)F��$،ǎ�(U#���nX�r@�҉''�ѐpe�3|#��a���x�;���\��"��-��ڢ"C�ih�-a?D��uO\�
�\aY	�'DMj�9y��
�#@���� T��rԀ��Z�D�XbT���F^}2Q�:}��Χ@��� �w�Ψb�ޔ.ۨ�ڶO�>e��c	�'ھ�+1 ���h�;��S�5���J:��Qh�8q�6I�����'s�2Of���hϐ9��1��+��)���'�`����Q3h�Dے$�
:m���ˆ@6)@���wGS�=/���>\�:��a�9_~ܲ&���%~ax��`���V�R�0�3��.u�����J�#pn-y�̃<Hp��!�'���i�˫!�Q���HU�Y�J�`�r��,>��؃r��?H�|i��I�* ��c� l5���&.���!�D�=kԾՃq��-���Ôh^�͓m[<�.	�M�� �e��xr��}L`z�?���Y4�,��x����#��@��LQfŒ�ze�ݻ��	;p�0$
LdW.��� �t�U)4�X�,��Q�A�!���vP�$)`��K� ��iP
l^!��\>'""=[�	L�R��а9!��5p۴u��A��{�ʄ��*�!�ІcR��VJ2:|��qT
��h�!���H�<�0�fY�V�f]`�+�'�!�� �]R�>t���F�f|%2!"O�a2�I�Ja$�* LR�ht��"O^+��#d��M����w�@��7"Oƌ��/�=P|�" Mr쀓!"O��Fײ%������) |�0"O��!��<�ȁU)Ei%���'"O�\��_�:�i�ȏ�tf��7"OD�Dn,�JE��Z0;a�)Q"O�A�"(���Ԛ�T�&]��j�"O^����\��+e�5��Rb"O.���C�-��K�i���xM1Q"O<�[b'�'^�0����=���*@"Ohe�6��<U�V��C^�E�J�Y4"O���F���������t�bQ"Op�[��ǋ��3��u�*�%"OJ�J ���)�|AY k@�\�zad"O��Ǜ�t�YtIGJ/\m8'"O��jQ�ʛz���`��ԲеP&"OA�˔,
��1ADC$o��qu"O���䄹���SR��0Az��`"O������A<�zbX�T�y��"O����N]'��ZD��A6�T"O��a�i�5N|q`��$@���"OɐIQ��R<1��JN�R�h�"O��[�jZ0:qD[��.�l\`"O�2�ݸY�,:ŋ�A��l8P"O����s����C+��a�4�!"O<\ڣlŸ}e\u����Z5��"O4<��LɈ=QL}��M�M	��bS"O�!&�A2��ī��X����D"O25����pX ���D�t��g�'�J��dI��G�y��	79ܸ�*�PO��iO>!�L���T�ip؍�޴(^8�fIҍ
}DݱÁ�?'{�PC���k�$٠�gԝ�?y��Lu�OO���'Ee�	+WJ#@B�Tz$�ʹ|�|XD��0r��0
�O��S��#
4�	�O�����rd��KٹH����dP�e^�e� ��ᓮ^ ��*��ܵ_%�ɫ!�]g�OH$�G��̼'��g}R�2>�B���8N6��8�LF0���>k�:ݐ�{��I�0-Z�Y���Y$W�6��îéa���%9Y�A�=E��/�ƄbdCT@�|�!�7[�Х��J�>)�On��ɚ9��W�E<�2���Pe����I|�Z���4b���3��mUJ�!3�hɁ�EɎ�y�蛶Q��:ýi82����?��S�'�����<C�����EKR$wT`�ya�!~����>^�R�O�����O�l�W�G��]
W⛽0>�d�n�(�*�(9K��'�#�Vl�=Uļ)�IE3�l�y��m�T�Ae,�$P5�0|�H��E)8�pgE3p��p�'�P�.�f��:W)H{���O�1�h�SY�*p�$�#"�m���H��8�'F(����bv�O���|��Iچ��a�H��@�j0_�X�� Ǝ[D0b�"}ZƧE�L�L�3�c�'��4�pȗͦ�,W�N�;�C>��ӥQR����"�h�Gz��X��P�5Q�'�����7y��s ���J�P�j�n�#i=�u'��b�N£i<a���VN��F���Ȧ�$��0:�[�mGb�)�$�O6Q��L���ɣi� ��&�O�@�d�M���P���͘O"��r��˸>��PD�N�`�1a'��G�����L@U��S�g~��$+\0���̑�0{�GϮY�d@C��E#*��с�i��ڌ��d�'x������%����)Z���\�9�pi2?��d���O�g̓[�"�0H� ��`	�I	�t��r�:qӗ��:E�C��#p�>���JI���G� F6�\Q��\U�x-�ȓM�j��C��R�(2��\��ȓ|ojh��ږ!2�M���
N��ȓT},��p�_�_|v�*T��Cy����e��P�eF*��ڥ�
& h�ȓB���;�䏉8V���S�J���x�ȓP����əy�r �,�pB����S�? ���E��@��Xv�ԣqz�J3"O��E��8A�H]b��u�.r�"O������9e�%��iґ�����"OfĹw ��g��L�4�Wd���s"O��	s�X�HAi���Ӆ*.:�as"O^��B�\<Tľ�� X#�\��"O�i��d	?���"�f�)�D�"O6I����;1��q�A���K?��S$"O64����:�T����5-����"O"�#[�Bf�m��.^�i�J��"O�i(������k�s����"O&x�O�8΅C��]9u�Y4"OB%�4-�Z&V�H�����6Q��"Ojmn�]����)�ߖ���'D�Tz4�̕o���9b�(�D���*D�4P�M�-cO�xq`*�s�x{�(D�tj�	D,.d�P��T�;�1M'D����kQ�sy�����Q�C�}Z�%D� iFE�$w^�k`�!r����-D�4�qE�"r��d�A�I�|��D��,D�`b��0S_�Kd�\%yS���+D��a��E5ET��p'�N��P���6D�d� ��*f�� AQ�L6+PZa�@ D�Pp��A �E�`���P�J"$�<D���ǈ��|\N���#��tIH8�G`/D��j�i��#4Pc$�5^�P�*O,�q���ks�IPǡ	5O���2"OFԣ��;AQly��H�xY��s"O�[�l�:v�a��c^J�8��"O>����SRF 0B��;\P�"O��0g ɯW?��)���2N\d�"$"OX�t(��S6�L[��+J�z�zQ"O�<�bo�y�!�5�
�
x۳"O����O=7��2E�&V�.��B"O�	cL�4mPD����P-6���0�"O��ڄ��3F=Z�9rp�;D"O��e(�"�l�ӊD*n���"O�x87�I�oG��)��[d^�D �"OL�� J�uU�96,Y{9��"O�m����{^p@��ŀ2x�l�"O1�	C�	��芇��
M��"O�jae[�O�ެ:�I�=U��8�"O���
�M	��؆�^	_�a�"OI�7-^#g��J1�ԊF�a@�"O����F(^u
��W��%x	�@"O� ��0d�yb�]��n-��"O����G�7$8RD��u�ɸ�"OH��e�t~veb�c]�6��"t"O�Ij�lE�eSF��&��orn��`"O}f)�,Ya&b0i�"O�ԋ�V�f�������7cm�1`"O2,:m�<>�!`�%#|���T"O" [��	�8Nd�R!¥-d�K@"OlH�#j
�V3�@;� �-���"O����7P�\lӱo��W,d�Iq"O<�$� P���	X*�$� "OF@�e��`A�D�@h� 	�"O,�K%H�<����[�r�@x��"OxyBDĺO��,�s-�i�*�8g"O�y{	��D]���Ȝ��b"O.9���Uޚ�`RIN�
���$"O6$2 �#���M�0k�����"O�B#eY�y���G��_9��"O���ơ�.˒̉�cФ�5"O� R�൨@,�HI
�(� E�ܠa"O��2�(��E� l�Q��!��Hx"O�9�HT�D� ��ĳ Ü!#"O@��� ��Q�����A�%��"O�]��so6��"�͸yӞ�s"O�m��憱#�JD�E�v����"O�hBp��g<�����T�""1!�"O���X/I����-ě<���"O�mI6��J��4"��U.l����"O��X%�dN�qd�Y�U1�m�"O�Y�J�<�f����}@���"O4��c�3����@���. 	�T"O04�F��9
�jL#f�Y�ڜ�G"O�͠n�;<����$3�ň�"O�̂!-��d�\Rd�E�L-�U"On\���*>�Xd��cM�s���R"O�H�D��v�.-�F�H���{�"Oh]��l�&o��bS�-4�bd��"Oց���N��	�� J�:��"O��T`R�	��CC�P��e �"OzmA*ߊ[�H��#��l�a"O� p���%8��8�`�q؊��r"O���F�-X���p�� Ɗ�R�"O$�j�c��Ez�G\�z8�"OԤ����%� <�CM�.�T��"O���/]8�(�J��8��u"O�1BN;c�4q��@�]H��ҧ"ORl�b�<T=n�"�d-W�B�"O�(!��M>�;E�ˁ�
�8�"O�i`%Ѝ(MdК���
�R�R"O�<($
�у�Uq��R�"OB��ge1W{`�j���ZT��"Oh1�e�J1�y��Ҩ!tL��"O̭�PG��y���y��IY�()�"Ot�p�
ްF���Zf��;@,��"O��!�z�*�k�!c�`��"O�TR kįQXbje۔}W��"O��p��+7;��nR�p�"O:H����nh�E$�
e9^���"O��I�5'�6$8�E�)7�����"O(�sE,Х[D�z���v�|�"OzU"0��ydly��#d�p��"O��xi[T���`��ֽg��Yy�"Or�w�Ыf{z���G۳z��Pc2"O��ҵ(W�[�p�����*��US"ON���A�J�<�K��Ʊ?��LG"O�bԇ���P7��kq���g"Oj��c픛=�.}�K�I��,�"O�����/qU���ѡM:  `�"O0�p�)��+�����+ȦcVZ�`"O�l�V� Q����@�o$tQ'"O�L��T�M(P�R��$6
ȹ�V"O
]�f��F�0P�{��]�"O<�ڷ&�̚�9N��R�"O�(���Пt�@1��e\x�@"O�	���h�8��r*O�_]f"O<�Bৌ`����"�p��"OV�e������ŗm@�D�"Odd��l7"�{Ō~&���"Oru:�Y�E��|k�E�����"O�1)��oEr��`l�|�D:�"O�U��'�
QaLP��C�I��E("O��FQ+E;�����o�p���"OH1U�¨[ђ�qe(�+E�F�X"O� 4aksKG7��� e���l��"OR��T�P���&ρ}�Q��*OJ�(�FH��$��Rl溘��'L�D�#���e�ʟ`�`���'�4��G-�Ѐ(��'�p	�'�v)G̚�0m�ٺ�K���ޕs�'54�Yc�E�mBS	��GB5��'�����`~��#-�u�^���'ˢ8B�)N�
	��aI(:�d��	�'Hbex�E9,Y�bCЛ*DE
�'|ּӢT�9q>Q��/�%)��a�	�'�BU��(K-����ˌ36~�0	�'&�`�Pj�.i����3|Q��0�'&P�!�*�B�Zd����g����'�ܴ3#~���P��
b�ع��'�f���l��7H�'��^��J�'�T��уI=mh�J��2"���'?�`H���:��d��F���(�'�X̨a��^��5
�bC��:���'X��;�xP5�2}�p�I�'s���B�����±j^	qzD!�'!�]z`K���h�aŬ_�4�@�'*I�#�QU00��KM7(��'K��{$ΛA�><{'���T%�	�'�Ƭ�@a�=�F,W3FxC�'���G*��W��4˗��g)$��^�U�q�Ѽ
aZ���5�H���w�	r 쇸�4ነ��$�r9��	m��	a g��1��<v����ՂV�k��qP�l�0���ȓ
Dt�V�M�R���蠅�ȓs�Tt
�"�6-�y�� S/a,ح��n�x�J�i $���N0!zԅȓ^�r��c�D�rS�Cs�U-_7�<�ȓV7��(d	ܜD\�@J��E>`��ȓK}���0��K�$
Ns3���ȓTAL!pq��J�l�@	;G�j�ȓ3�Q�d�W�8�l��>�%��{/�K�D�u:���G�ߨJr��ȓd}q�(�+��*��Q;Z�(M�ȓ\�Z$�/W�(ډ�Q�ѐ^$(u��+4�8��>��H
V�5u���&�f����N>��+1�0]N<��0�`p���in�  rǞ�Q�䙅�"�dL��茳{ﺄ[�/שJ.&��ȓ>�`�#0��B���U�%�^q�ȓT�m{h�v<b1(!�U�&!�ȓl1��/�9%���G�rX��ȓ*E�x�V����4X[E��$p�b��ȓ5�Lzʅ�y�\Y�P�[{�݇�x0�ӱNٺp4��C��5�詇ȓ��� "��=&�]�poF��L�ȓa��|pv����m:1�O�
�h���8�VU���Q9E�z��"��qX�Ɇȓp�@Jf&������WO�h�����?Z0 j�H� yp@;u��ȓ��p��);�H`aZ;��ȓc욙���S+\�L��@�"A:��_JhA3�!��u��*ȫ)�C�	3��8C.�`G�P�pA��%�C�-$6P �  �      Ĵ���	��Z�t		;]���dC}"�ײK*<ac�ʄ��iZ�v?�,x��	��6�^���!xtK݄-ݴe��ג�� r��DG�l����bR��ug��!Y�(��Dݚ�dV�xq:D�RH�~�l����(<�XhS� �2�͠)Od�H�!�OP��O����
�r��)4o�fR|���9o��,�U�ż���L*B��*ˀ��'}|i�O �"HڦWƆ`��p���#U&�H�$Y��V��O2��*�*�P��ϩ`��sDˑeV��fB�B-8�T�M��e�����ē+�q�/�����o��D�c�o<I�r��~�#�_E48�J>5@ŏhU�|'�����J*s�<�%,:��p��߇C8PH�|����zZ04�H>A )�9F
�T�C/�&|�-y��:��m0�K�}�Ɋ-�J �bC>�d�D�8BrV��!Ek|6���JC
�
h�s�O���bW�u��'��4K��\����"��l��YT�ߧ/B��:��҆j���I��y2��f�(4��������P��4t{Ұ�@�2�@�j�L*[b����(�?Ya+C+U�z�'���� }�J�'�6EPŗ!bf�����v.H��	ΟM�!�s�O|̓����䉻<�'�5&���a�$�{qc�	G8Ɯ�©D�=�@�#��²���Z�)�^���|"b7D�Xl
�'�<�j�G�,�i��7q���OB�!�A�VY���<4ħqb�S*�M�D/�(C�I��}S���U��/�VP�m�>�K<Q�*��x?�
�!z��D�&V�*�pec���*��H:w�&mX��nص	^Ԩ"`Jϥ��D��"�X��Pnǟ�)���*L/�L!�,M��b4R���<�1��49�:\&��@�[.1�
O���',Phx�L01E��K=t�� a�)%/��@�|��:UW���y"A�]G�x5�ؕ,� �sE�!
>�� 1"Oj�9`	�  ��D�b@ ����=��a��|��W,��y�/�H.tH����6��2aN�os�zV"O(��  ���q�!��'gT�ـ���L�
�(ͽ�1OH�=�|��K�Fq�+�
Y q���D�<)p��Uk����]�0S��Pv�'��y�ꂯwD��Y��� �����H��yr'��Ux�Ab��"n�l�4��"Sw��'��QEy��$IE:���#�dU��+�� �y�#�
r�c �U�X(   �  i  �  �%  ,  S2  �8  ?  �C   Ĵ���	����Zv�L�3ĴP��@_zԒ��4O��t��#J�+dn�$E�/�*�˔ɐ�d`BdƄYy�D8w'B�{�r�9,�K���&�D�Z6�8�U	�!�� ��(��9K�NT�:.� ��l#H;Z��Q�ްs�dA9���D�n@bt"�/Ѱ�[���)	���un )\*M2Џ�?0Na���3M���I
��A�X�+\6衱�#o��`(`�&I�%k��6A82&������Cg��oϔ��Q?^g�<13�^&A.�]HH�q�VJ_&'� �{�'�R�'���~ݱ�	.X9$��FD#��D[�hE��c/d���I�ur�i��Y�uw��HO44�C$���i��مq�l��DL�v}>�#�h��|��e�4�X4��)���̩�I<ac�XR2Bd�ALP8�RՎ���ɉm0��ɵ�Mc�X>��?	�'�V��SǄ<q�h�8 F�>C����$7Oڄң����(҄-�?f�0�3�i��6M��A&��Q����?]�'�Hp�%K� �����G�����(ͬUI�����'�"�'��.v�U�����	�܊)��(d�3�m��.˔	;f)��~:�(�`�12�8IH��ר��O�DP�@��Y����!��"���_�W��m#v旆k����O7A,MQ��D�6b"\��u��(���z3��H�v7�P��!�Ijy�'��O��Ӭb<�\���ſBa���r�:Q�v���Ob�'o�1���s�!�QF�'�@8i�OV1+�(�ΦU�'ˊ��yݡ���0�'-�uB�!�y�VD �U$�B�n��E�.���Ο8�I,uM�<#�ꆥ.��9���!)�a�V�OV$r�ŽX��h�1RL�X��d_�:���A��کo���U �eW���3��M� �0҂�N����H�����r�'Dq�^աG$M�g�r��쁁$���bsU�4���7`mBi�ƭ�5"`J� FӼ^����SY~r�Z>x��)A�$b�ĳ4�*����
�
o���d�Io��+�=���'��	ӷNsӊ\(�N֒$ ��d����@i��1�Q[R'H�U9��H�G��^>�������̒L�,Q�pǓ��ؐg@�Oh���
9|U�M�Fcb���N�Og��sC��AXz�p�h
�
V
�Ѳ�'5FX��Y��V nӤ�D,�t��@�t�N1;G��1�k@!Oؾhb�!��b:�IǟT������ՍV)�mp���9Db����<�M�S�iE�'�4M��W5���A×@���dO�5�^7�O�����Ye���ef�O\�D�O��Ā^�4�?���S���D�f���"�0D������Тa�v4��MZ�	��:jrݡ���OtЊ�`
��8��t+ýe�B+G�J7xb`��ЊE���k�o�,F��uB�Mˁ�x���2��0��d�#x�HIÇ΅ �M��!������]>��?��'NƁwLS<)�3䚠s�F!ӎ}��''6Y�㘉=>�CH#W��c�4]^�fDn��O������&^�L	�d˲x���8�,.���I��>�|����?����?�װ����O��S�*�$���*�3w�(!��@G�$�&$(��� %�"<[�_�.l�z�2=�ȱÖf¨Ej�0�k�>y���F�� ��;7�U�������O ��ԙqD�)��KQ�V����U!۴��'M�"}nZ�K��e�
o�u��NrdC�ɟS@��Y����'��ih�	�K*�"}���'Q�	1�� ������?A�LE�E	5��}�4�H�}ӖlB� �O<���O����Į#m1�LN��ԟ༪��U�P�a����H-���ɨ����kÕf�A�Ҟ��d�~O�3����p5���hO�4�F�'�7A̧"������X5B�X��Y�|�'�2�'cv4���Ӻ�8T3��Z�l�}
���ɢ&oresfL�IzX���]�C�`�����3�i�B�',哿YA�X�I��<�Jƃ{�(���
!���c�B�nڇZt8)qGY�Nc�eX����ʧ��O��\�c�\{��%��Jd�|!�'�V����M�N: u��`N?E�dm�m>0��Տׅ)Y���v$|��c�=�?٥�i2��S��?��
y�@�GW�q�+�`�\w,�ȓ5g�m��j�*���c䖿m(qEz�f4�'�M�	S�x�L���C�H	���O�F�'�B`�99�<7��O���O(�$�����N�L�c�G��x�E��`բ,��M	���ʷ�ͲR�x5+NR��' ���A7�x�,�D.���c���)�����x��XaGdբ4;�����X�i�֬�,�T�tAK$��V�;'Ƕ$Z�T1")���R��'ܔh9�� ��&�=ғ�~"��H0��-�� ,�A��� �y�ۣ|�fl��'.�p"�Ş�M���i>�	Lyb�N����5��u@���ĵ�:U��&O[���'��'�p֝��4���|j�ȭ+�6�Ð�с ;܌B��*M�.!z�!�#y��is�i!&B	����3G�,�[&�ra]���!9��^���c�#o�bH!�R�E��(�v.����5�+�X����I�D�`�KJ�8�tA��ކW6���43.���E}�b	"6J�	�D�`
�d�d:�y�C��W��B��Y�K��a��剰����ݦ���ry�lW9�y�O�r؟���&̜�(�(DR%i��h���Ce�i`���'��'�,Q�����i.Ѹ���;�Z�lT� �q
F�C��u�g�Lf$�Ic��ռ�(O�q�� � �2��5#Avv(���$Y'g�� ���Oξh�4d)�kP�k�`P�a�AT�'�D��D��և7�0*Ƶ�d �:�\	j�ή��꓊p?��o�N��ӂ��!@8L�����\X�d��Otuz��#L��M9E��;Y]�a��V�ԃ%�K��M���?q,�&�5n�O���Ֆ90�҂�ǫ]����0�~`�-l�y5�\VZ�8�����&���H��5O�1�F]vˠ:���"�$Q�&(B��O�0�3B���"�1F ���G;
�L9S���-��RL�2�X(���Q,r�����?鱼ic�S�J��(�D�t��fX�QΒ���!�D�$8���	K\�V���'؀P���x9��)n�t���LR�g�$ tm�	6�Х2�4�?!�i�D�Ԣ@��?����?��|B��Q_N�:�aJ�1fAQ�σ�=�y��fY�*~r �B@V�;�>�P���c�Sn$��ē9�}��W���0a�"+�@��p��k��y�-�: ]赳#��E�D!�J���$�@ؓ�ْ�r��MQҜY#�æ<�uK؟(b޴;4����&34�Q�+S*`�@1���X�jL蹄ȓ���3��ùM���v�E+^(Jpl �HO��O@�1JB��s��q5�eQ���S�
��c�$͆���?)��?a�������O��S8d���Z���7l�ՠq�:x����5&��rB�,R5��͕!m��I��V�A`�0��ـ!�	Ѳ����g�� aN�.;d1A�PRm	����'\JaC�D�]��G�XX�X��*�<m2t}`"OR�1��7"�x)
�O�	#��
"O�ѱ툂1Pv4 �i�A�$��\�pzݴ��;�$��iR�'�)B�Xq���z�,��C�Wj�֠ dK��'B,��*i��ԟv�"l,/��`#�,��j.��4�	-jj~�~�0�:a��lCG"�t��)Rw�'�(�B��
�>���&7-�t���䎫q���k3�=D�D3�G�#ְ�@�@4�^���&?�O�@�'z�iS@�<.����˅]��]�O6$����Y�I˟ؕO�����'��+Z�$��+;���׮	�6-���� �s�J)A��S�J	np��O:1�Z�`�!��z��\^њu	����?C�}���/���0�S��h�b�H
�)ۈhB���,�V���/�O�R��'Rґ�����������y�<<�p�Հe&�Y��!D�p����`�
sK�.'��DҶ�>�R�?�
Pl����H�6=�h@S˱�M���?��hb TQ���?���?������ 6I��Y8� ׯ^�.�#�����H��W�z}��F"D�T�Z��@Y���I2'����U��36����#��r󪆦cT6������L?������|�����u:�Ϟ/f`	q�ܻ7w剙>{��D�Od�d'��i:$O��p��\ S�ت�$���EU�<���˰x5��B�$7v��Z�!Ѧ���4�z�$�<9�*U�h��D"��2jx�jٱ-�������?��?Y�0��O���u>�U'	��|���� �S�A��Μ�`�@�~T��{c�*\l�qFB/4u"�y�iM�g~�dࢌ��-L�s/Q��@B���1�i<����$i��&�H}�UY�mK�=�p%!��%!f�7�O���F��4g��!�PI"�RL��"V�g���ȓGl�ı��:��M(&ƌ�A�l��':7�O�ʓe�x+�Y?y��_�!K�.<fi���hQF!�ťLƦyɇ#�ϟ�����ْ�[�lW�xhX:���e�O�iɸ�x��n�$���y��d�ў�#����i��r��D�I�O�64�1G��;Ɣ�j\�t=X��h�'��m��'t���1�v��]��=T����e�3%>|��?q�u�~X�P�G\@uy3�(u1�9��ɽ���-<��RQi�,z�� #I�	��|�0�4�?������L�����O��p��!vA7�3k��i�U��צQ����f�CeO��6Ҫ9��CY�u�<iq�OḑCE� !�*%^�Mb�ㄲ�Z���8Q�3!c?U����)74�z"#��1j�>��1�A�p��a����,q
.���i�Ɵh���O���;?%?	�	A?A��;{��`�F�	$K%X�<�����h'%x(�lہj�J��?aV�i>��+��>�LH��g٦;-��jɬ�M����?���ÖV�����?����?�7��d��P����"o�c><�@�iW!)���0#H����(�$r����#*V��I�,� cEC�d11AW�x��0��F�2S(���C|��(U��|�	0��x�i�[���B�-���'4�l��O��,��d�[
0��q˞L��l��[�<)@� �8�:CbRQ��j��Y٦�{��4�8��<�$���l��$��'ɡSl��ٔ�+�`���!�?����?1��8O���O<��O�D+c���1����O���#��z�\�TĀ\p�Gk�dx�@�w�#_�̊�(BM���1n�&/�<���s�b<��cQ�,�M��" �FU�-�I6�� :̠Q7&�n ���ڸ���iެ7��O���?a����5����'6x�h ���0!�xR�'f���r��L� A[��@���үO���h���A�'��܃C�l݉��ɟd��h<
����B}�|��f
 ]61lZ�L4��Iݟ��ɢ/��ب�����Rh@�/ɘ2R�[w-�q�����%��}�蔔;Ų�U3���<��� 
�P[���8h<�T��C�uǡ��^�d��GD��y5#:!b�d���$��i���'|q�٘#���N����XM��S����8��Q��(a~t[��F$�h�"��*�Ov,�'Ud���θ2�!x񀄻<� ��O��0o�˦���ş�O���I!�'!�	  JF�����GlXd(eM�y�7m˚kPVU���-JN�i�I��i�Om��?7_�9�K��9.uF�BR�I#30����G�{�!ʷ�l422��(m�aF�� 	3GL�0ԍJ�/I\�QG� �R��?	��i>&7-�O"~:��V�W�pݲ�D*#�|�A��"��$�O �=	�{b�*f�4��fՒ/1�(��Ή�HO�Yl�:�M�I>�1�J�T̬�a�HM�Gx����-e�!�V�i���'����&��B���'��'������J�#B:r��ʁ 43H8�P�˸6:����5|b��2a	�kdTb(�Q����c�j�$�Ab	�T����+ҿUj�$����8F������g�'aT�:t���XA��A;DY��4�?�B�+�?� �i ��'VB�'(���5��̙Q��<2�n�0;��M�Td2�y���=Y�d���`�0�*���Y��MC��I���D�<!��ˍx�<"�\�X|�)3d�'Je>����"�?���?!��S���O�d>Հ���%x�����N  u>`�b� %�nm�2�L� �aS�I��� h�mQ������{��,�b,	�=�u(� ��ч��=�xк���t5p��J�Q���d��O��r1�)V�4@5�ɳ�~�p"�PҦ�2���7�\��A��O�l�ܠ��I(^�ȓ�^��D�Y�si����L5�d��'0�7��Olʓ���33�is��'��i(:r�ѱV�/�n9�b�B�i���ʣ�'S�'��(V�'��	���5�Z͚�D�7J����ҝtL�F{�OA,d����ՁC�d����G��|�U�� 4�b��B�L8W���0#K�i�'�~U0���?���ir�џ�5��M�2�t$��y,�(x��i�B�4�֢<����M�T@�T(E��5�t��IX�X��4~-��[�m��V@ٗG�6��!ޒ+�x�M�bX3��i��'��/cv\��P:�]B�|��40�}�C���MK��ƌy>Z0���
2i����b�iH�S\�t��M�7gܳQ"��(d��0w_T��T�C͟t��ԇjzx�Z�Ř!t`|�٤��3j"^#|zK�AM֙k�D�U{�%�f�\�?	�d]ܟ���4z�韰#|�O�JٓWB�� ������O*�O�=�;t�&�*3�ߛNw~eڃ�-za֩Fz2�j�4�o�~�I�?I �mQ>��I'�!j��"�������"�A�T�Z��dN&A�4�K���=�(��хYu!�K7DP ���2P9�R�<�!�]�
Ǡ|�AG�R&� ���T�!�d	:&o�"g�����tj�.j�!��$:؀{Q��蛳i!��2刕�wn�	@:����=!�DT�[�4C��Հ�i�M�!n!���' �@jJ�6��R�b[�Sf!���"�܍	@�W,%2�Y��]&j�!��	�/T�I5�0=!5�! O�y�!�$Ʋ/��p��/+��x�G�(^!�䄈,n��a%`^� G���4HG!��̤s�H@�\-�t��+�"K!�D�7x�U���*	���)�
	^a!򤘠#Nn$�%��R�!��N!��l�p#,�+r���P�b\LE!��J#/�$es�N<���҃�/bN!���~P�#�S�]���ap#''�!��"���v_�B��D��7D�!��~a���Q-�7]����� �u�!���>T-���&b�2Q�@m:' �?Bb!�����	��b̦?�d)� �l�!�d�%#rHJ��� j=&������!��JX�$kJ�A��u�P�
-/0!�d��vQf
�9&�)qI$q!�$�~j����0A4�r�͇� �!�� p�� �&-!��Ir�D��:t�w"O�%+bi�;e��X��T��8e"O��gAÀ�`u�B[W��H�"OĨ�giR����"�Sl� �"O4ْ���P��1'���i�ݳ�"OdYY�*���*! [1He
mI4"O^�Cч��y� (JE�!Y\ܬ��"O��*P���H�j�dQ&)B"O̩�qMW$t�� �⣍(dc��!�"O� !��C�}�m�f�8PQ*��"O�E2t��іY��R,_O�<��"On ���K�3�	���R�j�yr�A�7��	T,��1�(����y�(�%~�8�b� Uì�:�y�+՞J�ޑ� %Wey�xC��$�y��T�*&J�³��8�ZL�����yr�;Xw
�s��f�
5L�,�yRQ�C ��p���*ň����L��yB��5.�|�E��d��&��5�y��1z$�(�t�ӊXԆu�aᅄ�y�!\(7@��HȽOܜ$�����y�IҔ ��q��&	H�4���۴�y��$�(���ͼBNtX˕����y�f�o2�t�#��~�P�0�*ׄ�y�
E~� z��˲zM�,`Do��yR��%:�
�G\�l��4-��y2Z�w�8���L̹�h �7�ϵ�ybR�[)�Qүވl�Z�ِ�T��y"#
\M�5��EW8lގ�����y"@Ǝ}�`([�$�h����$I��yr�[�-t�q�π�w��c @��y"�+/���2p�G0d��m�/�y�e
x�ܳ&i� xo(�:E�ل�yrE�,_"uy��� r��j���yR�%':��7o+
�Xs�J��yrd]$72�7�T8wd�ٲ�]��yH]���I�g�vT�m�����y�Ņ�no�,����~��1�r�Ε�ybkÎ f��F�y'�H"�K��y�hX�|_��A�	/p��D�!R�yR�C�м�5�c4RN���y��
(C^�b�HPbzj�f�,�yR�=���ӔJR:�2 �&�y�'װ�7&>�e�V��/�!��҂8�浰�)�䈤T���@�!�$� Na���L];z�8$�p�M&z�!��V<:L�BE���1�/��]�!�D5p��p�B�خL	R�Q`o�O�!�d^�q�����G��i'��@Nͬm?!���R��g'�y:�虈9fęI	�'vn���ς���H�aD�.h�9�'̰�q� �
����7)/��Z
�'�zy��,Z�)&��&�ߧpE����'����u�V!��06�_6/�@h�'�Px��	[!y��юR.2� �'���PƮ�p>F�d��*�8y��'e0)�,��Pd�j��ڄ)hTq�	�'���1���E������:)h,���'� �BeF.�>l@ �G�Y,��#�'m|��@O��3HΜ��j�M�Z��
�'��\(�Ϧ!�����c�2dlA`	�'u؜��g�!�4�:����>و��',�԰E+ҏF�<Ѳ0%�4E0�8�''Ji�WA$5�F��ŌXr
��� �5Q,0j�� PL�=zNH�"O���&�����k#�?w�гd"O�e���ӁL8"d�S� <R���"OR�j���,!�Ly��H��*&�l��"O���b3Blb�BeoC/+��M0�"ON�âhϳ�8@�#M�]�bE�"O63���;v�4��i�0��T"O�|���Q��ĳ�ሔ�N��"O�qr�&̡!��0x�w��0�"O� ˅j�l�ș�Eʩwj8c`"OB�;@	�42=�]�#Ko�����"O���SĚ/�N�����1?�0�j�"O����znA�b#��rAk�"O�Q��t7
Yq��L.O��V"O̝{Ԥ8h�(u�#B�'\�z�rS"Ot1��
��ؑ��Y8�9W"O~L)�D&8rF�+�BG	�Lʕ"O8��3�ٓ(g�m��Ņ4|�9ٲ"O�( fn��%W�j%M�
F��K�"O�<�e�?mۨe(�˜� �j��W"O���1�VI���[+
�p{A"OB%1��̪3$Z�K �Ƶa<�p�"O�1��(�q���[cM.93rAjf"O`��q��?+�.y9��;=<��s"O���5Q�BmBE�8x(���"O��9Ý�QTA�(ݪ�"O�lӁ'��Y��y@d�ǀsi�	 "O���	3H`d+ �d,�1{4"O�	�Sز'q���B
�"u+�"O�]Rgn������ag�&*��M�E"Of���ĩ�\�J��T��Nܒ�"O���ej^�S����C�D0?�^eK�"O8uAЏV6n֚����7��LZP"O2}`�Hձ8��yq�#	W 0V"O�!�"� *U<� w��> ��"Ob%��#N��p���i����"O�5 u�T����C]0C+p�S&"Oi�K�-'�&�āāP)�4hu"O�$&n�>��u±�ZlĤQ4"O��J�ϰ9l�����9a�	�"O^,G�F�Sx�L����:�l�H�"O̡8�$���k�
T	D�a"ObK2��'E��1h"!��i@�"O�2.G�G���0ovz�%�w"O@\
�Cμ{&� h�@ks���"O~�3���k.�!(O�y���F"Oΰ�%`I)�0ˡ�+C����"OBa(f).;�0=��ѱ*b �"�"O�|��哢@��X��\3!X4�`�"O���nǲ;N�k��JPJ�)7"O�A(�?cSȴ{��Zn�u"O�ty熐N&�@"���|8��*O��Cqi��Gޒ��& �&e6nd��'�t,X�G6O�!#�)�(�a�'� �3e��@t�%�G/ӏ3��#�'�Q!� L8�t��D��#~�i�'��s+�$9b�;��Q�4x��'⮡��%~�Tpi�G@#v3@٠�'��A���՛Qq�L��+��uZ�'a@�Co�2`|5��,��:,@}��')��)p��8gܜh��F�7�,a��'�&��ClR�/;�x��� 3�����'�t�Q�� �ȨY�f��Xc�<��'�đ��,�o��SE$=s�L��S�? ���F	\�;X�`�L���y�"O��E/�K¥B#7td�u�"O֙��L��}��5B�!�>Fn8	�"O~5 �Ǝ&Gc��ᇘ(z�u�$"Oΰ@a(I�9H�5h�,�X6�i!�"OD�'�Y�,x$�"��/�BM��"O`��"�5adv����A�P���"O�"\ظ��'�����.:Q!�dA�u�p[�'
,7�������X�!��˟]�Da�OҘi�R) ��՚5�!��R1��dP�2�v=3n]�[!�NoJfE�d�_Dn�u���!��E���R�E�t����0げ%!򄎻l7��R��8@K�d���m�!�$�F��AY�i�.3`�m�W �(r$!��L�E_�(���G�����Su
!���s$r��S�W�n�Xuz�fE�q!��[�-�2"�ܩv��D�̸v!��Z�[�̀�C�҃D�(!����J�!�ď�FtB��-�3)��Y
ŏ&o!�$�]�J���- �p��#A��.S!�D��pJ��%�i0�I�ɔ �!�F
7��HʔRL|��fI��bI!�m+.0��Bg6����*S�!�O:`n��[�K�>���,֯,�!�$�����E9�:dS'C\	F !�ė6X	�d�C����2!�lV!��ȉp��U�e�v����T�E3uH!�=D����Җ%��,�Pd_!�D�,%���u��*��4(�^�An!�D�
:�ȩ�c�˟v?�0�D�B�8i!�$@�D*YF/�� �p�K��=}!�$ȓu�C���;@�ޤ��Igj!�ċZ�U�&�G��ys$��lc!���??&�����4���Uˏ\d!����dy�F���{V�PP��!m!�K2#������ö��*C�!�č�3۔QTO��Fɶ��1��,'O!�ĜLJI#`bȪw%�UIЦ�5�!�D�'/.����S��8��&�1
B!�U�n}�"�Ci�(�$@8!�$Ѱ1��8Ï	��	1a	�qW��Ȝ�p��ɯ{J�,�,�GI8����?ŊB�	x(�0j��H3Q��\�UnZsC�ɤ#kf��"�@)+M��aא,�,C�I���ɳ��
&�4L��*Y;rC��x\j,��`*�����	PJHB��H��u(Q�;4��i�ӎK�o��B䉠{}��£�۶A�,�6 	��B�Iv|M�̈́��h� �+U�C�	�o�����`3G�*��6��zr�C�	<b/�`���{h��Š;s�C䉯%���ز��,_�����*cv�C�	�Ht�� E�_����H	 "�C�ɓGT�5�1�<oj����� h}pC䉖U�R����ݴ<��,�B�P�qHC�IvDP�b):�$9!�ðqlC��9U�e�E�5���3+�y
�B��2)�d!�h(�Qj����C��-zu�TcT�gaa� x`8��)?D��
������7�� �DRs�=D��k�E^�%f`Y���h#>$А�<D��(��nc0 �2E�@-R���D8D�\� ��kin���(]�@^�!׀5D�� ���c#X�L!�B�4p�Ȅ"Os�-8|���EπL�@�8�"Od*�M�?��!JG O����g"O��8�@Ca�v\2PF[�#�TEj�"Oh��h���Ƥ��Ws����"O�H"�͟.s�A��E�'a�(�"O�� 3��5J�^ ���
^��"O`l�K�%����� ܡtSv�V"O49sF�M}~p�N]&T.��I�"OF��@A$�i)fO�"r��	h3"O���K�����vO�p"O$��V$��s���8��"OL�[T�[�n����q�"0�p��"Ol��媋�k)����GM��0+�"Ox��_0n� ;�D.c��<�%"O�!�I6M�@��_�p��"O�����`x&��5#�+'[Rܙ"O�66	��[�ӣ}��諲a%�y���@�,�� @mV����yrʋl�XX޸4�6�2B��M�!��N+.x[����9�H9�aF�U~!��Ĩ@�htu�џv{LZR�ǷPv!�DO��"�qt�F?p�E�Pa��Tj!�$�,'bP[��=?iZA1`�D/{Q!�d�#I����\NI�}�uehl!�D�-wt�%/��o1�(�v$�1D`!򤌬/�<�����!I��%���ǎk�!�dLl.p�#��d�R����^�!�ټ|_.����*{�,\bF�Z�E�!��[�rA��+�j��l��EJvBȮC�!��i�P5�t��f�!2"�(�!�ԠI|��1 � e~p$d�>r�!����T� � \�&���)��7K�!�ƎK��;Tg CVH�1��!��C�_^�j��y7p��c@� e!�D�.HЈ�����|1
(Ap���9�!���Tqf쩃��?9�a��³H�!���u���aP��8��ԨË3�!�F�rc
������q�!���mY�����J�����h�3�!�d�n
������`Y��gm�!�F�TsԘq	�e�F�Y�eA8s!�$ʑIr0�¥���o��s�.Չ�!����m��#�#um������a�!�D�h�)��e[O[(�!���)�!�U�G�ĩ��ު1J�r��?p�!���HI�qBȹO_�����ڟ�!�	^@�E�'Z
L���桝�;�!�䕷h���9s�V'vF`��p
ۺ7�!�$P
W�iR�昅c/TT��kK3M�!��%G6�ŀ��,��C�HE7�!��.tI!�%�]���!*��p�O�=�����O��&�.lZ&@[�9)�p2S"O~�6aD�8P�4��/F9C��W�Ga�������63���h�bҋz�@��J���yIpа�OD�6U�5\��?�D� �Oz���Y?��`�A�C*sM,�۰�'|�'g������Z�@�P��j���'��!��C&l� ��(�� S
�'��А���4@,q�� ?H��P�<!s��K�49�o�t��	�g�I�<9��E2�[6(-L/>|RtǂN�<q#K�?K��QG�� �T(����G�<!�g�ı+&B�#9SH�s�SG�<� ���=daK���vh���"O��2F���{�Z����P�G<L��"O"��J�]HdY�u$�lz)�g"Ox\� C�P�D٢5K���"O�� vh��	Ќ�Rb��Y:�-c"Ov�%B4uL��`��`��q"O
a��#Or,��ERd�5"O�X���6`֜a���7�L��"O��B�H �Ipf��#��}�S"O<��J�&DA��0sh��P�Z�"O��(GN�+t%�ՐR��0i��c"O�|����pXg��,][F�;�"O�c"�1��i�W�oAb�3�"O�=s�@�{����e�1L��y �"O��`��5<d�ԃ��t��[�"O�YQү�R�R��u"[��<zD"O�<����.]j���៬K�.e��'�>��C��$I6�D��1mX� �'|p���O�:\Z�p��&_�<	��'r$`��Q��4}p�.	V�dI��'�t�	�"��3�Đ�2�B�\��B�'C\ *�
��on J�PI�E	�'�T��ۿM>�@hp�J`� 	�'�|�������汋�KP�@����'Y�i��`�MM��c�G�Av�p�'��1����Ap�;�Ά*@�\��'.6����D�+�PDHc�	XID�@�'Y*�D#�=U�"�)�׬m�DZד2qO��)uk�y���⣡�n8�Pc"O��p؝C�&����VL.�3��Dn.��>�|Z2��U����V;rB�����N^�<I�(@�$�� ��ȺᠱpV��T��-}B����I�+�e!��1��U�@ᄄ>� C�h5tXF�LU��%@T� `�6��ޟ���'��i����C�n��n|8FYIד �8&�H��K�-*�a$%��q��1�5D����ӗ1��30.[3�#�!D����d� �Z���i���浲�� D���#&�`z �uA>(k�}�g�<D�D�сDZ��d����7�]��<D�lȥ��8M,Ѧ���fn�M��Op�8C��#��+����a� �䮜�;��B�	�ki8\aP���_��u��$ �C�wX��kb�@�!0Tdۇ^>�C�	8@/L(�ah"D2��[���-]�C�I���H�#a�� ʐ%�t&99�>C䉡o�P���	X������.�C��2#_&U�v��6#������7��B�	e��(���\2'��U�&\/�B䉋&�4��aM�<r�:(����*r�B�I97_�(qd�V�hK,P�D�.q�C��.#�\�� G2���kvAw��C�	z񖭱DΈ<�}#*#�C䉓h6�p e���U�a`�B��	;�2��o��vnp=��b�M�hB�	�)�l(r0ϛ=i7��d��
�B�	�K娀�HXz�
U�Kq��B�I�6�[4(�#8�� S�ǘϰB�	<&�.9ɇ�B���Y��f� �B�INy�ś��O/+��C��H2zB�	�.t��I�e娵�F���w�ZB䉤+�lQq��&��q�U��)��B�<2T�����1KI�8�ri�%;Q�B�	�L��"Z�a����e.N`B�)� ڹ��ʉ=<�1�Rn��L����"OM(6�H��!1T�S�RRXA٧"Ox��� K�P�:��MƼwM`��E"ONL�j9S��:�eD;b�3�"O�L[#�	Rr,#W�SMډ�"O�)����23��}�2�(8��V"O��CJ�	60�H���&�rL��"OZ�c��J�j�j5��S:���v"Ot�����K7(e���[�7��4��"O:DGH7�(A�Sbܼ��!"O����>Ig`���	~�ʘ��"O��sׂU;g� �3����T�k�"O:���H�����FM��I����"O��["	�j��a!���"O�"�nƆU�q`��z���"O���Q+&�tAB�>X�"P"O�=+0D��)U��37�W�
���"O��y���f9�t��@W7�8,!�D�-�xu��m��!�:����B!���x���w.P!���!HX�R�!�� 3�)��S}��Dx��[N!��͕88����E���]K�
�'H(!�D�/`Z0P����6�r��	@!
p!�d5�,�ɥ逰1���0*�!�I88	5��͆�~�����3iv!򤁠OA��"A������W��=r!�Y�C"��p`��)2�l�bU�7Z!�d�*H �Rd˕)��@���+W!���,z�!A��F:HM�*�G�<@!��C$8�d���L�e���@ޝ*:!���6�H�a G�S"F��u�BR!���`Î�k�dD�� X�kF!��>Ρ2֥?�f]�@�5!�Z��<�s�ޛe�!��՜y*!�dA��̑���8@A��r�#H.
�!��vT�yq�K®M9R�#��Ӱ�!��!��U����%�4���e}!򤍗s�E�!^8;��01�`	:Nx!�d�1f�Z�z�i��#��yӒ�H1D!�d�ƎT
1!�$p������R��!�$�_i� 씜e)���O��Pyb��JȢ�v��yz}��Hˢ�y⬞)9���6�������M�y��R�Q����տ*�h��,�yB.8 a�5�"lZ�+E�U�y�Q��bY�wb�7{Le`tF��y�Lȏw   �      Ĵ���	��Z�)	�%���dC}"�ײK*<ac�ʄ��iZ�v?�,x͎	��6���,��@�fD�1X��Ȧ�̾>���l�@m)�M+�o�뎓i�\�I�a���I�$�Ucul^' ���.T-R�U�Uā���)�FP�+m��VZݛO��qp������ߴUC�� �P��! �\�H�4*���9�n�l��x��Dx��ʓ*�$����O�	��G�ޱ"�9aH��k��Ƀ �>����,�D��7�>q*��N �:%c��'�\�D���t���A!1���#��*Ӕ|�k�8#����4O�� d,�%T������]ؐ�O�i��R)wV�'>�MQdI���\�F� �爖+�\�a�C�>f!����ze*�O�(҆�v8�'Z�|��	z����m]0\e�qZ�D83�%!O<�-Y)3�T&�$���1"d�`�ȭ��ۏr���fL��<�z���J^1�󏧟�c�'�@��o�jy�O��lpP���q��8��]�?�bСS�<��� O<��C.du��??Q�O�gS��&��|���W�.$vRЀ ��=�� Tqָ �$.���q@����>�@�Ҹ|%j%� ��E�l��A��
ov��dW��~fj����i����?ݬ13�8;��%{Ƽ���ɺR���`�K�HT��'l(���;���u@�G��<�֪�H:"�� 	^���6�n}M�.4RB���'��I�1�@���T���&�����"X�@:���@\�KMH��v,Z�#��	g≄#,�'��6��,tA��}�fpa6
хdP<���Ö�^�:�&E�l�"�9��ʽY&2|��'{H��&�} �Q��'��Q�b�G�8@��f׈cV6�;-O���!�U�Q;�'���W��ēX��(���I�/q������8����/&T�%��X�>����dE,53x��ƳA�`���,n
bI�$D�<0��   ��(V��^�D��9p8�b�U��EPw�|����:u��U�L~�@�&R܂0;�^�0G˨X+L���E� 2��u"$�w�젴NC����#�'��X3:�H�3�՟$]Γ0���W䙺����S� 9L�����ҽrˬ��Й�|!�
|܈H��?�×�ϱy��*�Ɉ��� �� + ^�Y %�!���s�'�,�� Z}� s>��4c�/ �$�O)6�!`��!R�&8B�NE�E���       �  �   _+  �6  �>  �I  �U  \  fb  �h  �n  0u  r{  ��  ��  9�  {�  ��  �  F�  ��  ʳ  �  ��  N�  ��  ��  D�  z�  ��  ��  @�  ~�  � 	 ,  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P���G���к�ׁM;(�2�b3eR�35pY(aM�w�<a�E�8��h⎗b�h���[�<��aV�RP�����4�P����N�<!s��^��lt	�!�+���Ky��)�'4����G
-T��#EcA+$�ɇ�r���Pd,�!cx&D�C��"D~Ї�x��EcC�O6(�=�c�Q�*p!��\G.=���ݮ]�4з!�T2ȅ�N�1GɊ�� ȗ Ρj����ȓ�.�#¥P0�g��F0
����TH�	B�X�.Ⱦ5�j���ē<k���V�*�Z��U�W�`�Z� 2�}����HÃ/(U��lx��	�O����O����ъ[(����?L�* 80F��I���ǟ�'���ڦI@J��o�,1j���qp�h�$�=D��E��n�Ҽ��cQi������a�N���5Ox�O���IKVl�ТO�e1�$Ч)/}7�C�ɯ��M� E	v���v-C���B�I&׸0�@OElP`P��_�x|p���O ���gkb���l��>��*wZw9!�dT67�칣2��� �a# 6�h��ȟ� "�@1n�O�{�$�"h�D4y4"O�|i0B��l��)�b�V>~b᩶�.�Şw��0�hE&��	��*���H�ȓ*�М�V�ԙAN��[d�`�D��'��A��'g�������( �l@�
)x@	��+D�t:�A
*�������:LjР N5D�$چḽL��c@E�`l�y�"�O��=E�4F�]U�*�5s@��c!��!we�p@CĈ>t/x|jaEG	��'ʓ�hO�h���;[� �QĂ�n�� #G�3�O��'\qY���ezh���Y�7G������'�(	z�@�M ��cv�j����'̊!X�hɐ��`�@�
���F��Q��0=!w�?f��[7
��|^�1$�ȦQD{���i�h�m!+��A�r�
�x�C"O��h�O#F-���(��n,P��<����s��6x���JfԸ���8@g�=��If�I�Na��'�I�J8�\��l�-^�����:�Dθx�d|]��j�~_!��+��h)Q��@���Z'韜U!��E%1�u�7���l�l��&N�=\�F{���'�
A1*,f#�9���yh�5x� �S��?��'�T))pK0��!�H�<���S.viƐ:�L��o��[�,�?Q�m)�	�(Y�9�w�Z�l�L����C�	/{&R�(�΋k��-�%�X�5�n�=��'T�>A��&X�4��yC�/ ]J�i7N!��hO�S ��Y��-]��jRTp B�	�2y���
�19�DҒ�Ζn!�C䉋=y�ڕ�� k�T=�2,©os���p?Q��h�pK�f[ {�T�! �nX���O(T*����X0>��s�
�!��"OZ�*Uk�X���@̾O���"OB9
6#P�[<dS1OI���6"O2-���'yL�#��^�>|,���"O���5�EF�ɥ�K�:eR�"O88��߻Wp*q���7f@x���O����һ`���+��7*J�!Z�:���rx�,{pFϼ
l�Vi�J<R�m4D���U��˪Q[�ܸ=F��o%D��s�O
3sLmJ��ۘ8-��0ʓ�hO��6��� 7塀zP9[�B��+&h�� B]�*�r1�u'��M���r����O�t	P��S�"��B'tSZX�AY�0���
{1�io�� �z�`�(���du�� �7{h�bIv��9$c,D��HΔ�b�Bሆj�z���b?ʓ�hO�iy�,�Aȗ!%"�0j�i_�gR�@ F"O����H5OZy;R�H�i3ZdC!"O̍	��g^�9�B��s4��0"O���I��vT`k�#L�YyU"ObYcK��l�tx�����X ��20O������D2Dϋ�~��1��eM�uz�Y�� �$�~�'I�'p����0_�ZHrCkX� J�I��'�<U��#N�m�L@�B́یy��'e�9;g�N�gA �b#�qZ�	���y��"@ԐS���;. �� Ƣ��?9���P�q��Q%bU�D�� >^h�ONb��D�����H�@��'�77��i#3�:��'�O�uaP2�( Z��H�sO�%�P��\S����,Q++R�ŋQ��"& ��h3�O��={di�ߪy�6M��ޘZ�<���!��P�B��H�l!c�/��dς�Zd"OL	��J��T!�%p�+�׎�)��	`X�� * @��]��#V�Ʊ.Ҫ�#G�'�O�=y�U�uu����<#"he���S?��)�X�c�Ѧ)��q�.�'h&��?��4�hO��;`��y�D�8��kr�׆#B���O(P��h�K�n�� 蒜>�ԅڕ ����M��󩔼�^�1�^]r�S���5n�,�S�O��Q���I�|�dHI�,#5����
�'p�	�▚. >U��Ǝ	.0��	�'�$�*EH�oqȭb�4X���i�'4E�©[
vLP���욷a��q��'ab ��(_�}u��G����R"�yb��,�f��\�|�J0@�n��X���	;�f^�u4z%iR�jפ��W|R@�@��(����!�"m�,n�b�������A#�`A��َZW�����]�y�߸0��XP�E3*���#�����y��bV����A0�l(�7�"�yo]8#0]�b��,?�@]�@ �yR��*���/�*/;f�#�K���c�$;����$I.YS��#gň�$�p�=��=)�y�6@@H����Z�pL��y��B0\�и � �zg���yR��"G��!���߲5���1d���y�Ƴv>��6�W�z,d����'ɛF�'Z
���.�#Ĺ���G�4��$h�'/�%�ǎNݰ�z�F�	���r#�5D���ࣉ .>�@�bH��\��!D�!�Ȟ�jUv0a�_Ȁ�т�#D�آ�ŕ71�d���E,.�JA�&�	k���8y�~�fM�8S|�bE��b�VB�IsL�8�&�_!MEȠ���[�B�I@�||p�lX(_$�h;2`��B�O����Fفs�1����|��B�	6_�I�%? ��%��H�6�B�&n�h��	#nɒ�I@$v�ZB�	�bQ����F&��]�@��&?�DB�	�wК�q"U�@�(� E͝�<�B�I<O��T;"�e> {P���B�I'���S~��;�"ْ)HC�ɮ"
�M�A-[�b̙	B(C�	�2v8���
Q;�<�j���2�C�;I�Jyr�C��r.��֤U>Tk�B�	 n�ȸ�&��J)��_��B��3Kߺ����TT��bJ�KtB�	�Cg֌��Y|��K$�H�4�B�I�~jN����X����z���|��C�	90H��)]�8�vi�E&J�y�C��;M���4NE�E�p50a�[��C�~6� w�M�]��j%��@��B䉜#���xA�*]P8�2�B)�B�	�Ь ����b��X�b
�=��C�	5��Si�-kl���.	-/��C䉛o��̑0**B{l��g��	!�,C䉙Jl��ĴN�fcW�X�	��B�	�}@�����/7A�&�BlB�	�x���0p����uH�k��Hq�򄁮#��ia�8ȶD�Y�6��'�
�C䫔�kɔ��"ԥS!n���'d�ð���y�������P�DH��'����$��].��"�Z)A�M�	�'�h!K�cC�}�&�Z��Y/FDs	�'���+N$xW�e`Ek
�l�H	�'�&Q�w�ܯf����@�0mb�P�'�\�IG��	
�u g6�z9���� �cR&C���	qDG�� P�y"O�U���г����B-�t1�)�"Oi����.��5���3;9,|{�"O���l®c!�L�%%��2�"O���(Яr=v���.)��0�'�r�'�b�'l�'~B�'Z��'��u;eKP�d���S���(\`���'�B�'���'���'�b�'�'�x4�Ӷ �<$j��	6,:�iӔ�'�R�'�B�'�r�'�b�'$��'����� lD�l��]�*Z.!^B���㟔�	��	�$�	ٟh�������3}4�q�X`�򤫄��EB���	������I����	ȟ��I��H�I.y+�p`pL�^���ܿ;��q�Iɟ��蟠�	ӟ�����������D�Pf��!���i��$R���Iݟ���ߟ ���`��ٟ|�I�P�	-����dJ��r��'�X������	��(�������͟��I��I�B��<�S!��&P�����m�f]�	ܟl��ğ��	ğ��	��|�Iɟt��w��,�s@W/ Ҝ1`���e���	՟���ş����D���h��韸���I3�9y��K�fPv0�T*A����Iܟ@����@������������8��P�ͩ!�Q#�)2o�[�"�	۟�I����៤�Iҟp����,��/�Lh#,	q�`X�pj�%����	۟4�I�D�I͟������4�?��WI���p�U���"G	�U��#�T�4��\y���O�<nZ�FFp�C��%o����N��b�����4��Da��@��Z�(X���W��
bz�-�NĦ�ɝq� ZAl9?�/ЗH��A��>��m��s J���
�H4b1C Įߘ'5P�D�D-� d�Q;B��	C9�)�5T�7m�,E1O��?] �����+��~���R6_�!%Gh��iN�<%?x��N�9�r�ɔ9��D#��RG*�L�BM����22x a@��%/�G{�OR"�@;��W�)}<@��eԻ�y�X��$���ٴB�V��<��i�.<�N���:slՃ6l���'Vl��?	۴�yB[����&+3�t���=�P��v�(?1D6 �N����}̧*�BU����=�?A��V����i��^��^}A�����<I�S��y� �� �xE�w� M �B���y��~�Ѭ]~��uӶ���97ub� ���� ���L�IßlZΟ4:�F�	97l�D�q��<&w:���_[2�����tĒ`�s�G4X?��i�]7l��m��7;F4#��ϛp��cG�؋_������B>D�A���0�FEƊG#�ISk�a5�@0�\�A����B���d��èl�@#�jI�X3e�$ț�[^(��6���u��L�aR�F���[�@/c��;���K#^ŋ�ʞ�OfXDR�M� w����8 j��7ↂ<���2�ǭ�d!�@#�w?VX(�@�:%/"l�Q��:@�����( �3�#�ҮɪVU+w_�aXAF�_=�T����W9�M���҅qg���'\r�'����O��J�'>,��'��<�N�2��,�J��?)���?a���4�.�υ�k/�]�R�V3X��݂�Fݟ8���ۗ�Mk���?���:�'�?I��?Yc�׈G����!�B�XΆY!���R�ơ¥9r�'��i>�$?q��+O�A�!��aS4�a䁢��A�ߴ�?����?q�@[=T���'b�'o���u�����M�NY��鈇�Ԭ�MSM>�Qa��<�O ��'��*��p�9ц�!p�r(�K�3�6�O�=��Φ��I���I�<ѩ�t��O�r�(t��'F�3�?j�6��ezl�v<OV�d�OF�)�On�D�O����b��J�����B���$K7�@��������՟@�I�غ��P��?����I܄�	a �M��m�g��*�� ����O4���OF�d�O$U�����I��(�-g&���/�(5�13&��M��?��?����D�O����<�����;�4E���3��*�� ����O����O�$�OR���N٦��I七i��4���1%�~��6!I2�M����?)����O���6�ʓS-N�!���[6`Y	4�]���{���?���?��	�|LbԹi���'�b�Ot<�t3\-��jf&N�fE:toj��D�<��I��;,O���|n��1
&X��D�;44|��PDV=W��6m�O��DL�C��n��� ��П����?y�I�	3B}��c�Qc����cE2X�UX�O"��ǵn(����O���|BN?�*Q�R&�.��r�S)fuPm���hӰX����9�Iߟ��	�?���,������i��X�R�˱k���v 9��M��e[�?QO>�'���?	+��J�.@��"��6

�� :����'���'�<���>�-O �䳟x��C�8P~(A��	�cb��1Mr�r��<i`��<�OD"�'��C�OHV�*&"E�;b�zC� �7�OL�؇g�̦U�I͟$��񟬓�����3�,�b��5B�xr��-w-<�G�(5��?y���?�����O�|�"��Z����^+VT>��Vb̤M�Tnߟ�I��	���I�<�p�R�[��WI�M��oͅB�(�X�g��<����?Bb���?������S�F��m��W(�9� �¤@�����+�2�{�4�?����?����?9*O��D�)r�i�L%ڵLK|/���
L{��o韌�I�(�������/
�@�۴�?���V�����Z)aP���D�,��[g�i��'bZ�\�I�6�Sh��7���󉈄&I�)�د�&�'0��'�"���w�`7m�O����O���Ϭ>xX-�� ��v�&�@���poZ�ܖ'�H����'��i>7� ppA cߤ8��ɐL�8T}���i	�'Đ1�D�b���$�O���X�	�O��`��ݻLP	�A*�h���rb]l}��'O���'��^���v�鉲�Fh���$#�N���:��fo]�J9�6��OT���O��)�����O��d��Ek:��%`	�K�V�� #�`�mZ�{,8(��� ��Dt(�R���?Ś�o�ÊD`�AJ�;޲�WI��M+��?i�PS�5��x��' �OD1)4�ߏKy����eԅ?dp�D�b&1Ox���Op���(i �+�	y*p�� '��l���T�D����ē�?�������+�$h�W+2Y&6�åeKd}RҾ֘'���'�Y����Ґ�@1
��bbv!Hs�G��<KI<Q��?yO>Y(O���V��h�� �)��y��_�b1ON���OJ���<��-��
��t�Y����؝Q��ŗz
�	Ο4��b�INy�I�����d��!���4V偲Eԥ
����<�	ӟP�'xv�*�/�Iٰz�eB(�\��pq��'`jpo�ӟd$�Д'�4,j�}"�S�H�T�/�#���"I�}��4�?���Ĝ�
I&>!���?5�$�.N�5�S��4��2������{��'�H|+��V�s���B/D�(R�lZIy���6-PK�$�'���")?�BѲ6�3�#��Uc�A�i��%�'ӖTa�����A�Ь���L�7�1)%MP�]����2=�7��OH��OJ���r�����n�0u�e�>wS@y����M�Â�b���@��]�b�Nd�1i�K�`+%+G�V�2�oZş��I֟���MR���'��O��s��*rc`Y{���Bi�����$%!�1O����O�����w7@�#�S���l�#/��GcJ�mZɟ��/�ē�?!�����p-�C���H�����R�13'�\}��ј'!��'B�Z�T��n^)FsZ|(��i��JR(�A���yL<)��?iJ>!-Ox�Pf	��̖�
Á�	�v����:�1O8���O�D�<9u��|�A="�^�c�3"��'�S�yn�I��	u�	Byr���Ď Cw��q���� ����.$P�	��	ǟ$�'����>��1��(k�� ��fb�����lZ�$��'w �@�}��,?�| �fM�GF4��R���M3��?	+O4ݹ�dK_����$?�&8��_B�j�8ìR��<��M<1)O���~�U�W��[�
V2f����X���'�i�ad�,e�O���O�@�$|�lR!���YʙаD�gU"�l�]y�䀽�O��d�)2ͤh%Fh��K2K���#U�i�y�T�d�����OJ������>�2I�D4x@
��ۏc�lH�&�q���a�O>���'Rt<��ɀ�x.��6N\�'�v�3�4�?����?)��%�OJ���O�d�n�5%���Tj�%��Uqql�p�`�D�<���?��I�ڙ(�PbblR�bN�bYHk��i����J�^b�������5��&(6�C�.5}J���������s*1O��D�O����<A��8I�EA�,:��}���c��L˥�x2�'F��'��Ty� ǻ{<X	;ҩT\�Ĺ���:U.�:�y2�'m��'��I�F�~���O'�0����1R��2	���9A�O^��O0��<q-ORM)�Z?9��ɔ�l�X]"�ʜ7`6�x�F�>���?����dO�p��'>a2զŵ���P+R�j�B�3�J��M������DM�H��O������6Ҕ� w���<g�i��i�2�'�剓?�fP�L|����i���,�UL���@��0@ˉ'"剀	r#<�OeLyQ� {BT�yD��6F:^m�ܴ��$�	�R<n���i�O��)c~R�Pxd)Ǉ��P�؇�Mk*O  Af�)�S�_PaQ�E�(q�R�sS�k͞6�_�%o��P��� �����?�j��h�m�D��)�jL�+�6cߛv���O>e�I&\j��g�F($�1%iG�	uh���4�?i��?�bh�.=މ'h��'Z���2�h�`�
���2%��-��OP �#��O����Oj��O���848"qB"�W�\tgAH�g���nZ�b�dJ1���?�������"���� xf
��v7��h}�*��t;�'r�'p�S�4��Oȫ��[��	�4eC�ϛ�B���aI<���?9J>�.OL$:����Z���!�,� �$8�aZ��1Of�$�O��$�<1�������<�^���K�Z�|Ȓ���_��'4"�|W�h ��>�FA��8"��g2f��q���V}�'���'��I1;�ҡXN|Za�~���	ц�=6�4�q�	����'�'��8Ahc�����͑A�j��!(��}�~�)U�oӆ��O˓y)��Ֆ���''����eHԬ'V|Ui���v�K<�*O����i>mH��ǒw%<	�u�D��~=��
;�M����?��,$��v�'��'���??�"��J��`%��')��{�DAئ9�'ޝ;���)3�LH�Ή.��q�Q�XP��fе��7m�O�D�Or�iz�	��6�#���q��*s,����F3�M[��\�����D�Q�? ��H��
Ҳ�كC�#!Y�kw�i���'xb��e%hO����O
�	j�.�Pv��
Z[�DJP:b�ܙd@8�Iޟ$��ԟ$����3����R�IJX$;�M���M��B~a��x2�'�R�|Zc���;�n̻Q1���.��b��؋�O� ��d�O����O>�R��Ҥ!��Hn��kvF�$i����@H))�'���'r�'���@|�Qdʕ&�p�؅md��e�&��۟��	ß̕'>5��n>m��~R<���L],� ĭ>���?�K>�+Oy��Q��pŃE=9��#�ѭt��Ycg�>����?a������J˦,&>�`!�5G�쀙hg�u��O��M���?	*O`���Or�h�?�r0�q��	T/��0�	������'װP�qN-��OV��CSsJ(ɂ�ÛS�t����0HnIy��'�R�ö�����s����	+�X��3ǃ��.L�"�i5�ɈEn�y�ݴ=b�ԟ|����D� o����3Wy�=��@��	Q��'3���j�O�xϙ	^�肷EH�-Z<Q��W*�M�����'N��'�$>��^����!�5����q��73���ٴKۦ�Fxr���O�ш ��5���X%���\�P��#�Zզ�������	'0����}��'>�DITdl,�D��m������pF�OhQ�t���O4���OR���Ě�R��3·1��	aw�DӦA���{�KH<����?�N>��J�<9y#G��Xh��F)�
����'�*���'����	�t�'�P�P�̲�� �rK܀n���4�	-�O��D�Oz�O��d�O�:��,u�z݋Q�R���E`�N�>;�1O����ON���<��E�8y��)N�.���Bf�um�t��D!^�T��ȟ�'�P��ȟ�Ƀ|�d��ě(s_PU0t�_�s�&�b�T����O
�$�O�˓ʂ��F��ʜ�WJ�٨B'hr|0p��)m2X7m�O`�Of�D�Oܤ�6 �O�'�(C�]˛������I립��Ο �'W�Չ��,��OV�)B0㬽	F��3{v�:o�>|�%������(�������'��V���`��*tɀ�e*�0���i��ɳhB�Hٴq�S����3����(�|!Y�e�w�a�'�ۭH�6�'�B�Ї�2�|��$*ӝeU�;�a�dx�`p͐��M�d����'��'��� �d�O�,�u�R5V��C -2eȮ�s�,���a�n@֟%�"|:�`�ly�c��.�И0���N ����?���?I@�#d։'��'��ÙX0l�Ɂ���G���5ύA�v�|Bl׼�yʟ�D�O~��$$ԍ��F�+2�ށ��� �[H� lZ��X*��؅�ē�?�������ҥ�%[:*��d	�7�!"%�{}�`�~
RX����ʟ��	ay�_�żq�f�+	���C�#���EPУ;��O���%�$�O����������E5:��%���Ǉ	�����OX��?���?i)O6�9� F�|JcbZ6�-H�,�C���
4�@z�	���%�\�I��|�I|�T˂c�2��`�ԓ*�� %	�����O���O�ʓN��:e��t�L/͔���S�5�ؐ��(Ӣ��7��O��O8���O81٦#�O�'k0T`�
\�i3r�Sf�u����!�M�[�,�J�$W���$ZP�����w��)�lW� P����mZ�_D!�F8� ���I��l�X����>+4f�p�y��i�Fn/!��I�D���17��=|�!���+?64[�H¸(�"��Z�/{�	U�&��\*a����R�Y�@Ϋ]���"M͢��Yp�W�#�lz�^�2��j�(�2�m��/˭O81�)��#Dզ'�(,D���nh��IM�MB��O���O<��LvȌ8���VlP� �(y�`���y�����<Ѱ�S%m���g�Ԫ{
2|b�HGܓ$x�%��#l�(0@r��XK~]����A���A~�#��?�}�	�$�	:"QY�mF��	�U�V�0Bڐ�Ɠ':�q�E�YId��A�F��-�'Ll#=�O��ɀ
��Aw���=ۤ���e���
��7F��a���h����I_w��'�rK�T����&8Ar�BwCC�\��i6*R�
�����)|O��S'��<����7Qм<ҧÈd!3l%SN�./0}B�Ȫ*�xDy��1Vh�b;u�@s"H@9{��;�Nc��igӔ�Ŀ<����'b�;�,��L��+i���O��ZY���	���\pB�l�/V���O�-r�l���'�����Lq�)�������3�V�x#��-but�	��ʟ`�ɸ]&6��	ޟ(�'��E�fbW5QU�u ���M3��Q/ԙ�@g[g�!�'̅y8��YD�M�mG�Ub�Z,-���oZ�	�\T���_������N"P���~n�'#��'��Q+�<j�x�sB��Bpp�E[���I^�S�O�BE���Q;j�N�1R�6�l�'f�6mȖe�Z�Ң�R0U1�� F��PK��D�<1FDM;�v�'�[>]ST̈ӟ,�CLޡg,$���>׸���g�ៜ�I3����k� D���i�|z�I�	Ś���	(�2�`�f�J��N1>�ݙ�FǕ%]05�C�i`�}Y1��9;Z��D���'k�hͺ���`�,�'јu��g��	q��-�3� �풵��V�d�+��Hr���A���O������ٖ�R&)�8H�S[�z�ax�2�D�7J׀�RI���W�`c�i���'`��bf|����'�"�':"�w)�գ��ՙ@L�QQDI��Ơ Zu�U5~J�-@'�u�*E�dt��$?c�؉w˒B-(-�5�9\���G�h���ע^��?i�#�+��>�Oh���S�mԜ�;�X�l��c���O���'.�}@�S�矰�I�\�Ec�M��E���"r=Π�d�f�	���	a�O��`˂7&<��7Dȗu:��C�OZ�mڠ�M�I>�'�b(Oh�t���)x֝Э�=<̀���3O�ŲQ��O"�d�Ox�d��S��?Y�O!
���Fۮ��≒k�nɻ%k�mlm�^�PG\�!$�ۥm�џD���.6�}��|)�� a޶BVP�b!Wyaɔ�V�9w>�F2-�u�����R�ID��`�߄.�|Dx��h�f�i�4�j���&��|>�a`����~�Q�f�U�y2ɉ�>�Z 1�͜�t�Z����'�
�����(8nӟ�I ]}�u2����L���@4�	���-�I�Z5lɟ����|*�eF�b��(q7+ �&��d�pj%0iJ�J@4a��.��x�?{*���C�<Ԏ�I�xd�d�6G�8�$��-;����%�b�'�I,V�d����Hq]�9���#���	�$��i�S�O}�X�;V,�\Y��r�Z�[�'�r7�Ħ_`���A��Ӛ��P�B��<�j,H��	ʟ��O���s��'Xn���odl���FşZ�HW�'�B��7b�L��MX(R9�����|
a�.��s�Ҩ!��т��q��D�h,���a�@M��؉����-Z���X%28��s�`(��Igpp�ɻ�M�3��?� �)
��t��cnE��@��U3����![n�æ�K�9��S���@�ax�D ғ���CcF4mL�a�iǲ��@�itb�' 2O�1pۢ����'�2�'�r�p�		"ǀ.	�� �,ĥ2�:�:R��	� ��
0x���K��]1w��|:��>���%��� řr����*L�6�C�ܩ*7^�Y�K6!����}���>A���/,vYH$�$<h�4C��]>@	��n���N0�"��Y���	���3��L=[�@P�j"����ln.m��J�nb�a��IʣF�2)�'":#=y�'�?�/Or18�o�H����a�>��u"O����.p��q������"O���3��	G��h��L%��!�"O@�Ba T ��D�J:���"O8��/B���QAję�:�S"O*@���B�I���ЀO����Q"O�j��`��C��p�8��"O|L�� �6�I��c�6��"O�Tj�\�֕A����F�`�i�"ODA���
_����:b�d���"O�!Q�������p�W$����"O�IrT���>���KM�:��)�"O�\Ð(��Vv������T�ƕz�"OL��7��*Q�`�R��˛es�l�q"OB��ïŝ<4�y3�Mf^@�"O������K�ԹvvN:�ئ"OXy��ٔb%�c�QK�@"�"Ot`
��S�i � #�[x[v���"O�
g��5�D��g��E�
�{#"OT���C�SN<3�`�1�+�"ODQ@�,ph�����T�Q�.��W"OV�0����<bD$�?H�9V"ODyv�P�u/H�J��r�`��A�!��T�*��a〳J2�*�]�t�!򤈮=P���.E�1b%F�T!�ę�aB1��g�Q֣�f�!�dڊޒm��E�#7r�y* ��z�!�d1 a����m�3��5k���!�!򄀪L�:!v��?�v��@M�< n!��	_��	ٷ錦H��������DB!��N3����M'>:��ذ	!��K_BЉ�e��'�t�Bi	�!�DH&`H��W�����P\�@�<)G�Xo?� �,��pQ�槀 ������V�l!r�㝝^��Ц�'Z�1KE-�)'8��IRI�RnVu��e.}r�r��|?q��K5n{�eQ��O�Fj���v�ңgDb� �k���{�E�ˆ>}����?���C&�:�.
�?���al��h�)���?A0�:���!L�I#��L}��.!��J�@
y?��_yJ~b�#@�Y����9o�p#�O�J8���ƅu�X=l�����(�	7�6Y��#.dwP�� 	L��'H��	r}�HU�`G��`@,��B|ŊF���O0�f遊`A�QM~�'JL$��2Z�� ��"2�@`x��T�_��D����`���
���HK5_�9+��M	2[Dm#d.`�U��/��b��ӧuO��"�'a8�S�-���GLG8}c<D�N�H0�I��,�d�6F�Y�3?Aa`=��\��GW�Q҈����F?AH����'S���OR��O:����E�
����k|Ӧ+�KA*\�$�|�'9�0�3e�����⤂?���AD�_.� Ѣ�$?���*|�		��3}Z�~r��@q�-(�\p�����
��OVX���7�YL~�'XH�Qq����b��f�%���T:Uw�s����^� 1�&�%��D8"�,�VO�{!�Ts��nJ�!��2(u��jYw~@!�=�g}��ȦK
�}(�NƄj4��T����@Y�F�Ӏ�BZ|��2�Ⴂ,�Q����+3glma��m���b �z:r�0 ����O�S�F"��b��6/xlk�+I���j0)m�h�v�	�-Mt$�7�QҼ�d��F�Q�-HV�zD��M<�l��1IS#ɐA�Ę(�gO��-�>�̓  �X��,]�d��g�\��'t�`�����n%�Sj֑^gV���:<�N��(^��z�[��*���G�J�,����|��J� ��q��,�[H����i=,OPt ��ݾ�ԩs�й)������I�z��V���0U' ���e0���*�(H8�lF���j��lP�٩�'��܋��I�r�X���q#��ߝ8�>��� ��u/Q����D�p!�w����X���0{�h�&0� ��A��t:��!&Fa��Ƌ&i�t��ap�i�L7�	< �)�A�I[���[�e��Ov4�+�.,D
a�	u��P�I�=f��l�
	c�65���TkW�<1L�)C�+'>���P*;���� �ĸrT�p��C+�
��7b_JX�lBu��$h9�r\wp�2-�&P�H��ig��rӨ'kS"m@q��6d�8�?)�)$��[ScB5* �P�)ګ"�Q��D{�O��t�A�7m]#��I�L��� GɎ�8W��R	Q���Y�;���w�viYk
I�J]����'R��<���hO�O<,�:��';����$������F����mu��(|F%���1P��&�<$���s�ڤ,Q�l�-�)lU�s��<9��$[�3�<e	eK�=@�E�ޕ++h���Y�{[\I���	�8<��᱊�i~�Ի�ͅ4Y۞ъǫ	}��?˓(Q:բ�%J:)�D�jS��"~z��'�V��Ѯ ����b-Z�4�EK���'>�ڌB�a�($��@7���y���ԧ�u�*�>��C,���3q����C��C*�D���OӨONq˕#���ʼ氱)��)d\q� �^.+��e{�S�O���)W��4�FG�x\�Q��J���T�VB�n�j�k�'��B�l-?Q�JԄ�����	W�Q\���?�\�O8��O&��禍���M-�(z!bҸ|RXũ���%vg�`Z�3I���#�E�Z̈X`s�'�8 3��:�dF�'��1	�J��@�j��*CI&x#)OP� E���$��T�"�­��剭K�	��(F�Ky{��"Nظ'!���N�=���?�N��|��=���Z�긨5ď	���#�΃;a�������@��1ﺰ0�.t+�u�b
=V+�����A����?E������Ő��8 䬫����-����"�҄�%�K9L�@�[S	y�l�'(�j���3�u�Q��q��@��@�ݚ�{���?��T�ֳb �RV�%����(5����)�t{��b�O2Lx(�PU�~b�I�������O�)`~kJ�.�UH����]��+@D�|V �f
#Jكŋ/�ZA��ǡJ��Nģ�ԓ �͓?��'�����\�)Ήg�B#x��(�M�/M q���wɬ9x�b�2_���P�0�O|�{�Ċ�W�����A_�S��+j�� 4��y�<��x�코'(�9��F�ɧu�'�@HsAf�6O����Rpj.q)����b$@IqEn�Z� ���dO�4wD+TdO�u֢1:&�^�R!�DJwo�O�%%�ֽ���+Q�c�N�P��t@��-~�2Jǝ,~�\�#�R��d��f�W�h#t���/�>�3}*�j�S,`�l��!�B>����P�~�@�ɶ(��I�T r��"�2��g��	ö�)u+��~�F<C��2���	�7���3�'���"Y0�['�Tk`oʣ�yZ0�Y#�Dc�'�a��g�C?��&܋7]�h)CLJ/	Df��@��J�H"6c'JE�䋐F;�yi�գ� ؀�E=N<Q����뛰���� D�:�3f�b�+$H�K)� y���6`O��q��1z72��e�U�A_
d2`DU� �s+S*6qO?�I�[�I���Ѧ ��a��d�1n�aĀ�_�qO?�	6㊬��-��
�� +%�D�q�ɺ^�H���'�*<ѧ��^����E?I�$۟'��I���X�'\�Z�=W*=����$�>��&@L�f������i���	A�b��/OϤ�������2S���%�)J>l�f'��A��1�)-$&f8*��[��>9s�W/L���+bOYxܨ��W�3�x����bvɧu�u��*B�nU��#��?��H�g��K�O�(C�2iB���I��y�鈘Tĉ0��O�|�OD��N�
0�@L
D��8�B� �T�^���~�d�C�R�x�C�B�3�I�-�6\ض��R>��kFo2d�ɥ��r�2f3�Ԅ��?���iT]ë�;�����hʐQx�=s!Hŵq<J �'%�M�'�����y�[`����Av�e��(��Y� кA	&�)ҧQ�艣 "d�ZF�:\r��N�O���
�3�D�@��4������D��(�0KV��"�����1f/��X��pܓ$B�I� t�g�N��$���NX C���Jk@\j����6HEP��I��z��z�S�'�4���a�0����2���-O���4��"7dn�js��cͦ}A��	\�pq"eÊ3,�̪��W�Ph�@�1�?��G�P���=�I�?����Rn>��Dl����`�����F�=�7��0�\�N�8V���$�9�	���3|f�a��ߞ��',�tA�E����;EU$������Z�p�f�� Hp��Fx޳
�I������h�
���d�|��u��!�	=��3�oD�)-���M��M�M>`֟�6D��=�zMk5��|��G�6}(�,,ic��q���)���N�T�2�@+wk��1�i��@*f2��<jE p��~p*
�+�����6`����` ̏P�"�-̨���	U���*�@�4I��ԓVcG�|���S�a��"HTH���'u�$ʡ�q�u�O|�I.mN�lڵ"1��#�^�Y��ީ"7�]I%�1zj�3���{��9Q����аx^X��@�0^d���5[N��Q�:L� �A
��$V���'E�
A���҂Ę�)��屳��9Pfc�l;rF���B"�&�h��֦'�A��N�^�� =U̴;��pc��ǋ3,p˓�(O��kw,��@M�W�X�@Y�@���x����4E�/�`�C��Nt�ȊC�	���!��&]Tء�F���qT��0M�Rla�GQ?�Ҥ�P,S�N�c�MY!�˅�z��F\��u�\���a�}b��s�,�	�+�.��TCE/m�����m6����t�-nu���ԭQ�=�f�`a��ħ��q��xuϟk��q%�� @�h�`�^�w���n�?b�|Fy�'`��i�d�N�w�|ux��F����C�D1.���	��K�G��[b�R(��� (�M�<xS��7;��h0� A�O�xli�o5z�OZ�YDL�>N_�1���#D�>|�7��a�T����~PL���Q�j������!=�>�
Ó2Ty�N�_V���6�&<@��[\!�0�40��9���#t�z`K��2iӚA 5���wӸC��d�� �4�p���;��Ҥk挭3*�R1)E�35~p2��>Q�jB��j��` U�4m��iVE��d��J���1j�y3��Ti	�!G�p���!��7Ә�J#E��$P�O/�'�d3r*�F������%�Yc'r��Ei@�Q���>S%��!�A&�2Ax��*�
+M�>��lа/��>��Se��p�R��	Ǔ,�I��B�5mz�(���$P�t�zB�2��8��� !Hֵ�w�wS�lЃ�)R��&����t�CwR�N5L�{�j��p<��55:�2�灊�ļ����z������VK���I�[��٢���>O
�h�ԫ!�E����O����������?��ěD� ��'�Q[3�2?��	V�_�:Y��n�~���z�a�'8bT��ut�D�!jSA��8֍K&�ܑ�'�]"F�`�`H|�	:�:ql�"y�24�R�X�R�4��h�>L�-��"Sj�D(���
- VQ�ǌlޙ�b+�3+_�`���-)��)�񎍩Kv�9��e&����8��{���45HG��!ܠy�l��8y���e�I_;�hh���=b����$��BĪQ�N� �}�K+M��*�&���L��=}��8�Z�j�O)�2Q��:;QR��c��*�$����S����-�i����y��$��|���I$`ְ1���@36��j�J?��>�b��	_�E�M~�'E�,!�BG�+U�A�͝�$i4$0�'�t�'����2�����S�A�������p��|8U@���]�5��,7}pI���9�#��sv��Lm6��E�s?��k�ny"b�^�L�ֽ�DCo�b�<���ۃ*	��P�G.WJ�ɋ��kD*�����2�D ������L�9M���(�ER?	ӕ>�{�dև'��hpR�����1��¨���2��l(����>SI*����O@��^~�mFK?������Qe�߈\TJ+��	 ���OF�O������C|1��Ɂaޠ����!%�<A@c
2Z ��/�(+�:kА��(~.�S�����S2��}\9CӮe�~B�	�^��b�e�$B{!&�!9h1�o�X̖'�r�$>�
E䕸l��ɗo��F
ٮ�E�plXVB ��D�o_p!F�@�oQ�)�mC��XMr`��?b�U��'��Ez�b�#[4�E
� �	��f�p�E��%�0�H�I<$��Hrǭiyi�M�l�(�$�wK|x����#a߶���Ɩ�"�!�C�BqqɆk�1N��ِ�c�IN!�A�)������-M�lIЕt_!�dF 85���BA�Kp�)C�&Y!�� [ʡ�W��J�K�E�sX!�$��EsL�R�nW�+{��{&'"!�	�-��Ѻ����x�v9w��7b!����L��ש0"z�uXD�!Z!��R�s(�i�6m�,R'$P�5!�M8i�����'b����դ�!���F��+6�V�GT��Q#݀9|!���9��(���_%���!����!����ݱp)��h���KDU�!��e���X3�ʛl����`	.�!�$�(딀� ��	w�&eQw��*~�!��I�V��(`GL�=��)e�ڳ{j!��V�f���IX0
��s�"{�!�D��<\Q� Y�u r@i�N�6�!��]%B$@�!Z�5��q�W)!�_4�H]���=�,e
A%ؤ(!�D�/2�Z@P��˘U�p1� �}�!�DR�_Ì��6�V-S�d�
sF�!���I"�8�L��*��G��!�/�%I�i�<x���P�8Ǝ �'�*	����7�ΨP�7[�ԣ�'��[Ṕ;�bu�f)��8�'�(16W�A�&髀BB5.�ZE��'�P�:��7p3�J��̄yJ��P�'���R6-β04n� �Cʍf�.�8	�'�4 �&��>	Z�#�-Z�u!�'cxR�_u`� �+N�b���'dQawe��M���"�Ƽ�Hl9�'�ΐB����K�$0c�a�9	��D��'��y��/F�!�8x�k� �����'3Vd�'�J'h���a�~
`�
�'�z(P��߾r�qc��H�98�

�'�	r���"� }	0�8&����	�'z((�3�V?2!�X�l�M���	�'h|	�������V�"w6�i�	�'@Ա��r�t���ߞr��̐�'�uI�Rh\�0H�"^�o�@�
�'�� 8��*`Y�hr�����}��'tX�P��EK����O?]��I�'&^��)�)8��bF���~a����'8zh*��$ >��J5v�
	��'1N�Q����j&T�J�!

ri��y�'E,I#��M
	S��a%"�
�'�@�D
c��!��RU�d�
�'�4h�F����p�%7`J�	�'�s�\ b: ��}��H	�'S�����ٳFcb����(v��h
�'�`�9x��!��f
�݃�G%D� ��C#+�P�+��K){	����)/D�p����#e�#N�]���-D��ڴB\�OޠX�@NP��PP�4�0D�� G̚�6�\���v�a�C+*D��q���]�P�{"ƍ�6��ȃ��'D� y����jln,[C���p!s��%D�H��*]y�Hq� @�v|��H.D�<:�H� e���#H��HL$)���8D��Zg#�R8�
�`L$(1�Ij�N,D�XH��6�ۧL�]Z�!0D��k%f�&I�p�Ԕ�ɰ�!D�� �h�PA/(j���h����"O�e�C�6w���T(�cҙ��"Ob<zCc��zpx� 2eѰkJ�U{�"OZY��h@�sfmrdj��@)�"O4�A'�B	p�AAX::�0�3"O8uÃ�פ�@�& ���!%"O q���4 �)�r��P���"O��Sȝ�@Y���N͵R�T9AS"Ofp�䐛l2�hV�B��!C"O^��@�~��`��R�!�Z��E"O�ٲ�Q�Z��h�b�!x�lk3"O��dʅ%P�����$�+v����"OBXy�
��OApdR�"	�$$�9e"O��s�ʍ
�`Y�
�8�[""O����H9z�x5`ql���F8#p"O���/F>;�t{��B'5����"O:���
�9�Mӳ���z�8p��"O����C�n�pEY��NT' ��"Or�p����{�&�'f(VК�"Ot�x$��B7 ���W>�B�	4"O(�z�̗�7\8�6�9D��k�"ON�[�	��'���#�b����"O��m�9����Ȩ(�~�{@"OB��2n��@�4!�'�@:���:"O8e��6G1~Q��D���>�37"OڜKb���ez�p�K &�DP�"O@�X��
t28A�ʍ-?�n�)"O���6��(5g��iH���w"O�	�� &�����h�	��"O���c��J��0��O�W�5�%"OZAI�@K9xHpC�45F��""Ozɨ�*�.,�b�!Ƨ�*%1D���"OE�ǉ6Am���̄�R����'�qO�)�!!T�(�t|y��@!�$J�OH<���ҳ
'��[Q��ti�u#��Nd�<Á�	��� �Ӽ0�Zy!U�{�<��
2E�@���ȷ@?�TA�+w�<�VO� 0cB���)6J��dx`�]�<	�ޤ=����a�;���d��N�<�5lG�/�"�b�Ċ�"���CU"KG����R�$��&��T6�8@�,A�x�pm��x@��'�'}�|DzH�<&,e��7q$c�h�U0
i��']�jH�$��#��&�-²=
�޴�4�ȓF�Z<B��(��E8V�IV�����B≍s�JЀV����+���p�nC�9+.z�R�ƛ��>(��+�B)hC��UR9�A�P�J����02TC�	�*QN�"����"��	t�P�&"O���� ��tx�ʧE��"O2i� $�wڦm�5�m��(E�>9�U��a+F�ܶ:�]A�U�ﶍ��a�\�!�7*��`E�s�)��+�����1G<	�PnS�}��ȓu��Q�FO�y����i�+k��y�ȓ j�a�씍6�����$���H��P�`F�/���iV�H�{���ȓ@Vʤ����^:��Q��M���5�ȓ�4��%� 6�a�+����I�<1�'/ʴA!J�!p�{уE�;�A��'�&Aj���Tw� p+X�-^X$��'�l�)�%D/�P�y'L* ���{
�'��hW��x�lP� O�D��K
�'��� '�. y�M
3��D�x�	��� f�j���T��M�e���R���!��̆���9��H��"�Frtdb�C޿MFC�I�$|�;7�d��@���%�,C�	�x���PeC>�rV�ݣ=s�B�`ht8�MM�(Ȫ)��C���2B�I���!{S�Q6~9��S#e!��C�	�>(�|�q�9O����S���@��B�I�'��)H�ͽ#p��D�ɵ[�B䉶.��5 ��]�C�8i �k��1pC��}���h��<<��J �B���C�ɹ@FU��j��8.�Q:a�_Z�DB�I-;�����g	F����a B�ɓ,��R��%���Y� �2<0B�	�g���8H�*:ry��+�=:�.B�ɶb��D@��d�y�HJ�F�XB�	(_�,YD��P���@�	�*�TB䉂�6�f�%HMR����% B�I!�z$�#��+8t���'C�h��B�.Z���.��O�@����%d�C�Ɋ	ʑ�R ���b	;�xB䉋@.M��fY�nͶa����;D�^B䉇&��#7�1Gf����%��C�I� ]���	{tu��˝h�B� ���J��@&J�ܼ�ECJ�<�B䉼<�DlбNN�(��
�.�/S�B�*�� [��ʹ=�~����(t�B䉛-�E�!�S'$
�1q�坕z&C�I/xrJ�w�|�p�Fڕ$/TC�ɨ;��	
3.�%Ș�g�>C�ɉv���CG�;G/�yX�g�;'�C��{n�$f��)K�q�s�� t�B�	��3s��Ok�9��.K��B�$|���C��
�]Pt���B�I3�D�R��ܞ��L�B�nB�IFwtY���,;�9��Č6�,��0?!�"����	B�A�/"�鷧Z~�<�NX�2�M8�$Ն]a0%9"u�<Iri֐x�h@ZR�V>t��Ć�[�<a�`�(|#� �Oɶt��` $��W�<���>8��鈄��m\���p��S�<Q�d�/�:-AD��z��O[[�<ѡ�+B�����C�9#lTkv*"T���$��7�P�KEN��Ȭ���7D�샷�ѽl (r�����ɚ�8D�a3�?L^���J[)kۨ-��f1D��Y�"�>W:���r �_ۂ�S��1D�T ��יE�L�#�n��T�|�!p�<D���3G�<66��)�Kf��Q�C-D�4A�gM�s<2}�P!¯L��$�r�,D���T����a�3�8f�Dʤ- D�\��m2�|x���Gm+�邒�<D���I�?p�l��AA�mP�Es�(D�芲�G�o�:�r#)X\v	"!�!D��a�(�dcle��!�-:�?D�4����\��Ǡ�n�p����;D����^�D��Y���ݠ~�Tu	#"8D��;�gF��&�(��	tXNa��4D��d��'O,�B���jvB��eh'D�ػ`́�(�d�+���-X��@u�8D��ҁ� ��a��7��T(6 1D��3��}}z�I��)/����b�;D�[7$�w�(�FxP��H�5D��B"��C�~0��_�*Ypz C7D�ty$Kӊ&�B�'�2gj�P&0D�� 6%a@��[��P�Ӭ\`�""OZ��l՟zG�|��b�;{g"O�=0eD�"G��tpĠL.7���'"O�(�2�Ƒ3bJx���-^�pekt"O4�r0���X��x�G�F��$�"O�(p��`�x���%fʐ���"On4�+I<2�����
���"O�DK �ɉ@� ��'�J&h�P"OըP�1@p}U�\4sJ���"Op��	��z}$-@,N~�m"OV����9JLX)��B�y��k"O�l+GNbXF�kdk�?`�A"O�Pd%�`Bld��	���Q�"O`D0S#R�>�re�"���;�"OD}떀"���g
�7L��Y"O�l9rb	��|�8ŪL�;��AC�"OA16@��9:H��G��9k��I{s"O�
"�X�'�"\I��L����&"O<�s�@ �.��ؐEW�pX"O�S�i�0ja��Ѧ�����"O�	�V�]�~�x��I�9��	IT"O�0����9�U�A*͓XQrt�"O�!ҖjU�X �	0�P~@J�� "O$E ��5��HJ�ÿ;=�D� "O��K�c��;�zpc�o��&7�\3�"O[�Ӈ�<�F�XƮ�S1zpY3"O�0`W���g�xA�ƙ	��,�`"Oz��C��0S�r@E��� �� "O$z��J-ePH݃C�5G��)`"OLA��%Y�b`35��~3�uCr"ON�Fl.\��u�2�ޤ��"O�� D�L�wDIB�d��m����"OvtK�nW�q�xa�☮F�<d8�"O�D�7�8OE*,��	6�|A"O�j��eTh�oѨ
*��""O�= f��Hި�³N��UBl1�"O�P���oh�\���I�eA��r�"O� !�ߋujt�3Tm�g��AE"O��憜%|I�s1@�P "O$�g�+'h�щI 0�c"O4�A�O�#u���V�U%� *b"OyZ�̚!��&i�:$� ��"O&�YS��5a���A�27x�J "O�}s�k )�dQ�G�+6ɀQ"O��#�n����cC�����"O���I��p�b�ߝ0���R"O�cF(�
9�x�	�⑫w�8Ґ"O�P��B������X��Y�c"O~A��R&�ƴ�`�ɴ&t�"O2�9S�,,�5h�N��	�gI*D��(���C���%�_37��1
�
$D����*]�hX�yڧ������C4�y�Q
*.H��7�J�A�$���)���y�>/{&첷�V9fl]ZRN��y�#�5��.ּ'� �)�AͶ�y2-
sb�0��E�!�E���y2 �I)S�d݃h)1��GX��y�P^��Hc$V�5q�d�1����y�a�"C���bf� .9ʘꑂZ��y�_{̖ݸ�� AFu�` C�ybl�/��chUUr}�,Y=�yB!��x���ce�ǋ~�~��`BX�y���i5h��b#A�>/i�׊���yB�̙h��#�Ґ������T�<� x�ʑ�M�T�XIs�f1u�e	C"O��Yp��a8�+��#pH���"O,8�h�<vr%;v��i,\�9�"O��O07��`��*��Y|6xr"O��PJ�jx��� �Z��0�"O�,�� ��Ԥcfa��m��	��"O���G톌M�hMg%�)5�BU"OZ�I� ϑ?�zlBUB�mi\��"O&��"�;4�ۓ�E!�2���"ODUp��=��ݕ{t�R�"O��
�`�_�l�����;m��DU"O�dBS�G
_g���G��w�L "O���eD"E��5Gr*]v"O�%au��7<�(�H��\t��"Oޭq׉ؤj�FuJpG�TnZ\ �"O���al[	���hW쒋vP���"Ov�������!��,V�n��"O:x�BؓX�)���Ҡ7|�ܐ$"O��bGX��+7��sD.��"O%suk��s�?k�)u	!��N!:  ��7�B?���$�>b�!�d�0�� �G" &�n�!�!�$�R���Q����~��!+�m�,8�!�dD�P'~ ���ӂP��\)�lּ�!���:V4Š�]��B�Sd��!�Ѣv�r�h'#H�t*��Y�M�!��{B��;6B:o�&4łֱ!�˶>�Ea�b�l�������q!��(�ԥ�W ��ʚ]i��I�S�!�� `[��e��s�`���s�!򄗇x�k1N�$� �pG홻.�!�D��L�^����N�@a��i�\s!���x�8&-�=;�$B�ՇM!��%�9��c�/�6�2�ҙa�!�d��|�D,,e�J9qӬT%��l��'��Q=Ū({5+Ϣ��*�'��xY����Q��rXX���b�<񂦒�?���sBdB���4�Хb�<�WŃ$Q=r����Y7y(P���^�<����"&�i��	6t�`1q+F]�<�w���ī�e�\K�lH�k	^�<95��4@l��"�P�w-Z��v�JN�<�p�+sA6�8p�2�r�*�)�F�<!f��
�V���H/+D j�WF�<��jF�v:�Y+g.��(*����AZ�<�FF|��ArO��J�q�A�Y�<�iQ�"���Y�_�%��|�<����'58�@��ԯ�\Q��!O�<!$��\� p�𮍩�
Q Sc�<م�W��"ܲ:�Vģòq&���'Oܑ�i�N�ҡ	$ބ"/ȸ�'ꂝ���o�ČJ1���'tA�
�'��E��J�CG��@��Q:6��R�'�
I`��3}6:��� SfFp��'��$A�n�"�1WiQ;4��a�'܆Pچ�݅,' h����4C�L���'�Mh��,Mfd͚�@U4@�Ȉ��'������tqJ��
�3In��'#0�Cu�د+3��ꥯ��:p���'K�{�G�GgTȴ�4{ߠ���'��L�Dc���e����Dx��S�'T�s�'�/c�å��?mX�Z�'>V�����4SOj8�'";8@ !K�'o�h@%��!Gv(j@�@����S�? v܁��Lo�d��N�_��t�P"O-�dn$���#'|�p��"O m��S5~��pP�N��)m�q#�"O�!`���]��{����Y�4���"O��b�ռ_A��P�͞�]�v�9�"O���&�B1Rm9���	������"O�%%�R�Y���遉E�<��`�"O4�rꑛ<���*Ǹ�L�����"O�;�G�n�H��צ�	l6n��"O���
?1SPl;#4Z1P�"O�5��� �C*�p��a�**1Z�"O�T����/(H���"ʮ~�("OlDA5G��|۬m��P�~��M#�"O`%j�+\w|�T��B��<=1"O�"��U�n�2L[�G�01�ZAS�"O^����;�-p�`�s���"OD	�Wm��C�XI�� o��E�"O���	5�x� 6��t����"O~ �/�Ir������3��	H5"Opu���Fl�5  Έ=���a�"O��wI���D���A�4E	��k�"O��q��+E�q�6�� $]����"ODؐ�8�z�2G�g��3c"O�r�A�-i ��E�����"Or!y���n~�p�4?������\�<A�
����}K661�HR�*@D�<i��%-s(*�"�w�����H�}�<1W��ID$�!1W�{�2�Xu�Nv�<���׋���0�(X�#�&dXe��r�<�D�p���Rŏ[�2�)�`,�p�<QC�?Gt�ywF�@���CsD�f�<�� ��AQ$��#*�t�w�Sa�<�W�]Fj �aLWd��x�(�d�<��/�Gv�M0G͚zB�����a�<�I�(WV]KQK��6A���F�<�G(ׇ�A� FT�VXe��BB�<Ic	K=�\�r�.���dd�<��	�#�l�Z2h�<ت��C�<A��F�<N��1eɒ��B��g�UZ�<y���n�`u㣉T�[��PZ�"�A�<Q҃^�����V�}�|�ADz�<qՠ�7
���5/�,K�ΜQ"cVo�<aJ��\X�(�t����h�<��I
{2�`'��Ia�����m�<т
:�E��LR�:��Q��Fm�<�Ë��R����LH��$����_e�<�FJY�S��E͊!f��L!OH�<� m0�� �%�V��a
���A�<���&?6t�����|��B7��<��b� �zX�� 9JA`�s!]v�<���P2�@1����f9l!� �t�<�s�Е1�=�fb�V,��1V�z�<�'kM4cj��3ҸQ�����Ry�<	7�K$R��k�aj>9����t�<�2��#'���	�$��3�����q�<qC ���(�e��ႈR"�x�<a��_�?�\jVK��y"�j�r�<�(��2��|HVH�,qF��%��w�<�gg�"���{�
�!i�����Yu�<��Ə�@�}ӱ�F8RgP�0#�m�<��㓜$>�eᶇL2u&�����q�<aaA_�xb�Y�¬Q�v:8�+5��q�<�3���".��r�08^ذ'�Cm�<�2#ݳI��sp% O��РvI�M�<� ��;S��9T�� ��j.�Ȱc"O�QLD�& ���ݺm'�""O���'J�;E��: �Ԛp�zaR�"O�l�4B�Ry��s�$�	Ď�q"O����Z9�"U`E�g��q�'"O��a Z �z�� J�$�rxs"O��G��=,�.��D��3��y�"OM��)�����E��t��"O��R�Ƌ�ك�!��m��"OX�2� W� ��e�J��2��{e"O ���Z�%�-a�O�$9	X�`�"O|-8�� vq����Џ���9�"Oސ�!kA�'�,���JU�H�z��p"O�I�(��^uXM	P/`֔���"O̤:U�� .-`Cw焀[(��"Oz)��		4K<�ȺDT$ ,u��"O��p��N�[�Jɸ1�P\yn��"O@���s�0�R��*
��Ɂ"OlQ�f$Ę���Ü�I����"OPe3E	��A�Z�X�&w�l�p"O�5B.�B���:���	rhNHa�"O��'�ֈ2_�J5iA�DGpB�"O�\����+PI��I2�T�h���"OjlA"���P�M낢N>W�(���"O4��U+��z�&�I����"O�l2��#\r��0 �+�$|�c"O���Rh�q���ۺo^H�`�"O��sP�T:j/>���$��	Xrm "OX�A�E[;?����$
�5>�"O6pZD+Z�  `a;��ǈ#�5��"O�C�#N0�pH��\���8�"O$�{Τuj�٤'P�_Y�z�"O�Ԓ�G2�b� b��q�bu�p"O|a�q�&m@�m�8�ԕ�"O,��'�T�u� T��U*[�Ҕ��"O��"�k���"ŨEaOP�|`RS"O���@�W�2h��Tt}����"O�@KdL;��g�	��S"O�kgl�{y9x��޳U��� a"O�4)�k�9<�I�piؚ.�nBF"Ol�qæI�uRZp�@(G�Y�°��"ON�9US3y�:�p��d/�TAs"O��q�ް.�.E`�h^u@�!"OL�(4��?Dl�U+^6�e��"O����J>IJ�	RfՏpR�"O6�{�(�_�a4E)j�J<�"O.HZ�F̋:�0r�i�) ��\Aq"O���ɁMCT��hxV� �"O�Uɗ��=��Ȓr@T!5EB�"On� ��לeM�a�V�U(@%v�[0"Oh�����\�(C�V����"O~9��+��&�Sj	�G�"�!�"O&��bϊ'�p�;So�'@���h@"O�H��-(ǰ)4d@�w����"O�"�
D�\۪=1F�R(v�8!"Or��
ʝ|�XpU![5iҖ%��"O��Ibo�*&�<�@�<3Ɏ��"O�))��|��@�`�G����"Oly�@bY#�`�	 �%�<�y����Ԡ��j`�š�c��yb�IX��%CX�
E��U�E�yR	������]�5\�T8�y2��z���aj-60�cT.C��yb��(G����@њ0�Q�� @ �y
� P�Q#Aܨ nv`(��7�v`�"O�@[DMm�:�S�g�?2�d��"Op�0�BP�"��]K�	�f�� �A"O�}�BA�w/����ӫb�dݒ4"ObjW��Z�VUiq������%"O�Hw"�,.�e*6ᑫw�|�"OR$Bp:�pp3�O�'G�tI"O~��&�B-�}I���8�P��"O��a/Y��t-�a?X���(�"O�dbj�2#N�i��ć�m$v�[3"O>�h#W�U�Hܫ�E�<r(U�b"O��P
%f����fڎMEBA�"O�(���<4�>'�lBL�2"Obi�E"��"|4��F�F���2G"O�1zR�f~PC���*?�3�"O m���.��4`֥��a*2�� "O�)�S�R1WY��뷃��o��"�"OX ����B��C�RB�a�"O��J4C����P"j�4oP4X��"O4�aA��ft�J0)�����T"O����\֐r�j"X��S!"O�M@�e��(&x��T�D�_�K�"O����ꍀ|tb�3 �\�X�t�C�"O(%���܋P������9���AD"O.@�܇<5qR���*A�]+�"O�Ё(ҝ0Xx�x	;,:��0�"Oਁ@�)e֬�k�!� i6axf"Op��p�$>Vn8��ԛC�²"O�\93��n�����W$+,�hP�"O��qADO:��Dj��N�o�v��f"OR�	S�˭uh	2��i�<� "OR`Q�ޘ��BUJ�<ߖ�@"O�rMWo��%Q��+o��|0�"O�L��㏘@����SL�i�6%X�"O�Г�շi��|�0�=r��Th'"O�P��_�~!�"̣WX̩yQ"OT��#��VMx���<A��%"OȝC���vrHT!�%����˗"O©l_�ز$�H#��ո$�*D��0E:>�p���Z8?�Av�*D�Ȕ����h�޽-xH1�r%)D� �QHŽ`N���M%\")p!�9D�䚐�ִ��yf'�%���F�8D�ly6��=D�`eȴ��T�`s��9D���ΥT6�3ֺ��@�5D��p�gS�*���8 �C������5D�`
dm�%1!�`���)��ɠv�9D���i�����R&Sf& 30�4D�ĂG�C�p��\�Q����L�0D��P�_�;���ᩐ%��ac�)D�pj�k^�0?.x�!"t� �Y)D��ˢ�M.7�0Uxv�HbN  )7M,D�DK��T�=�f�
#�  L"�Ii�*D�4 �n\4*5j	ṍ�8�"q��#(D�,�f��g�J���^�Em� 0�J&D�d�V�P6x�L�2��] Z:Pe�%D��i��z�譊������5%D�X!�LA8Z=�Y��n�>w`Z��AC!D�� ���V�Q0s%�" +�q�k D����Dcb�0g��9��%�=D��x��rat��$$��}��C.D���S��!���I"��p���1D��2����ek��ekw�IlW�R�!�D�y)�Q��M[Z�2���
Ԃ�!�� �Ly��1J遄H߇q�f�!W"O�!��eY; ~��eU?�d�9!"OpA)�H �PV�b�nl��3$"OxDC2��)�ڥ˅���4n1#"O�uم��=6�x��!A�H|P��!"O��R��s&4R�τ�Vf�ؐ"OڍAUL��4ߖ욢NiU��3w"OZu���:B�f$�%.õq>��1"O&��u$�IŞ4�tϒ�$+4-��"O�\Hp�B6X�hY��B�a*�m�7"O�cѭ�(	��y����u��X�"O��i��@>yÀJ�-M��u��"Ou���{9�slB*D�D�"OЌC�aP�
��u�S�u�p�!�"O�E�����YC�XUO@ �y���1@ED�0A�4��N��yb��2������.�ڭi)ɿ�y��Ĩ�|\Kq�)w}���0�F�y�j���<�cI�lRd��d�	�y��7~�&�Rł�j���[��<�yBiQ!:��7j�h-�����C�y�(4����Q =a���JUH���y�O"wx���ԐT	�u�O���y��-� �3	��C���Ҷ��y�@^6�)3�DϮ	� �6�7�y"��"<�]`�C��B\�&�ɼ�y"`\�/X��1�z��if&��y"ܲWr�*t+J�;~M� /^4�yB��<K�r񨱣���)s� �y���cf��b$Mt[���'���yRj�Y#�Y���T�l�&5���%�y*J�2�8k�	؀/����bT��y2��a�4���2$��X�h��yb*���d�8uhY-x�{e�V��y�KŞ(�J'&i0�X4���y"�ȟt)� qL�v܆QB����y��@�@h�\�BZ�i�dmҒ���y�OƣM�Ȝ�����L�q)�yr�ֵ^��`��B �����8�yb�����V&�5���@�� �y�口7�,�)���  :=� h���y����O��໵���@wY��L��yᇽ`E�����;j�rd*�)�=�yR�� Yk�hA %C�a8da��%�y�I�Bu	P�S��Yb����yr�@+�v�pDF��]m����b#�yr�ŷ<���r���S���q����y�T�lu���V���bԈ(�'��y�ԽD�,r�bU0$lma�$�y2�L*t�
�:҇�����.)�y�kk����"L�z�@�Y�D�y��y����'I�oZ�q!-[$�y��$RʧDq���a���y���$`��rAYPL���9D� Ƈ�g'��@��T��z���!9D�0�3�+�|���,N� �<(�"8D�Z���k�L86��)U�B�I�~D��S�L�0y�	@��`ܜB䉙\'���e;ơ�4j��B�C�I���ه��	m�Q �J#l�B䉈@:r�!Q ɴU-j)B���y�*�B��HҲ�]�Q�~����ڀ�PyboBZ"I�B�ۦ,�\���x�<��I79���*�	�d)k��u�<� ���B(4����e�b�"���"Oh��㢅.GSh�AtϜ�9�6 8p"O 	+c��
t� ��쌚)	5B�"O���wC��eg���E��wV�j�"O��u�
��cU�W1oK���"O��A��byd% �j�)-E&���"O��B�@_��!:���Q����"O�i��.նM�$��89���A"O��P*&ے�kE'�42���`�"O�@�d�*VXg6F�"i�3"O��"挝(3���3��Q
�1A$"O��c������W�S6<9z�(A"O�Ჱ`��t^����C��ƱJ%$%D��p�_,V�����CƎ�X8zB(D���ոTU&hD�-=P`�O9D� �Q̙�t��� � �b�s`�8D�8I��)g�(��-�*l�N�Y�3D��[�	!*�֠!$��	6���;��7D�X�b#[8O�Ap3�Z� ������4D��ks��4B72Ya�d�$xĈ��\�<����v��	�&�δ*��5��\�<��LR'a Ju�˰1����A��|�<�2a�)2F��u�۫H(hq�~�<)��D� ���)r��[S��y�<�`O7�*����,p%RG�s�<Ѣ "a6�+��Y�&�!;Py�ȓ���[����Y���Lq�$H��4刅k�D�D$=봈I]�x��R�̰���l�p= �i;��u��q�,��\�YƐ��oCg���ȓA���)��1GZջ� ՄP�� �ȓ7�t-ᱪH%v9���e�ʼ�ȓR�J���C�~�E�K�w�҈�ȓS������dw�!��ܖzY�`�ȓ*W�$p&� f~��FMÕ'��A��O�N�ط#�~"�� �7��`��K����q�K�^"d�8֤�1z��p��zg���T�U�8���⇃#O'R���r_�THRcÇ�<�j�O�_� ��ub��"3�UJ���I/F^��ȓBSb�*��E	�h�%I�?��Y��!ԢH��j1$�� �׽?��ȓ@0�丧F�8�B�As��o�H��ȓ*l�d���\�x������{��I��0�`�a��1K�.X ���,8�4���bWHe�%`��{D�IX���ȓu�8����\w���3G�"
�zL��f��B*�7+�HL�VH;����ے�sb�˨h��F�L+qK���ȓfl��a��JpE�ǚ*PN֙�ȓf���{vf ."������P$&�P��H<̐�	�w�l�2��A#L�K*D��IP�� }��@!-��`��؂�	9D�(�d��-��1�����1W�$D�$B�%R�OL�|W�G|��I a#D��p0��4yLL$���g�T���7D��	CL��
\F���拖w,���E0D��� �+6������Pd���-D�|K�K$~���u�ѻ[��Љ@�/D���G( o<|l!�HU�h���.D��іE�"r�Qv�J^�37:D�l)!�\$^�x�/5�l��b%D�0�f��t�X���l^��1��#D�<��Hְe9�a���
�Ekv� D�� N$�����T�fdHK,\wҝC'"O��Zq�J1pg�Dx�G�<OR"���"O�T� l�+fP� z� �r"O�q��*�fO��oX|�H-"�"O&� !Ĉ�*},)Gc@Mߪ�"ORԘ"hN=&�����@���;�"OZI�q��VR�R�/S>9�H<{�"O����OJ�LH��B�{�����"O ���ɯU�^�ˇ�[-E�~m�"O�BAM^��p�t��<l�$��@"O��H��P:��pp*�?N�m��"OL1B�K%z ӅɈ	��c"O�h���/ ����I]!�"OX������j2��)�+�E�p"O�8#�Cq6rg��1��Q�R"O�2E��u���v���j>{P"O����%\�\��`G\�,��h�"Ol4q4B�.Im;�fD:Fx�"O��T�b��aA�FX&-����"OL���j�&)��	8��U�ݸ��b"ON��(E��Ƀ�$הe�� 1"OnC �,��2�d�$m�Y"Q"OȈ���:I4���UM��ײ�p�"O�9P��(8a���ˊ5��y�"Ob��	 `��A bҾ	,=�t"OX��i�Z�I�T���j�Q��"O��2D��� ԭ*�m�$W0QQ"O�� &E(Z�l��͖_VXy��"Oֵjs��ELaQ�F>3�H���"O�M��Q��aQO ~>f��"OtQV�ۘ+�R����IU�l#�"O�͛�녛k�
E��lS�Qz�8�"O�8J�"�6m:�9�eƷ}����g"O�,�|�UIV
~9���UB�!�d�4`�b��W#�9�S'��h!��J$j(H��2O$� h���f!�B(#L����-@���b��6!�$�|��E8Ƅ�+��@����}�!򤁤K89�&d]'	N���a�<e!�$�\p ̉&k�	c�Hq���*a�!����b��?"�T�*����!�$��d1��'R�Z>����V�!�$!?6(��٘N,����ǔ�
�!��1���q�1 {*�[�$�]�!���FX��C���`�J�EJ�<�!�ڔkQ����$l�(ye%��95!�sE��teӛzÜl���'PD!�$�2�-�h\�|��m�MP!��܌;lN9*!�J��~�񉘧?!�d�(�dlrCW
 �4HR�)��D3!򤆄R�ʴOM��(x8V�Z�I!�Dܸ2��H�%�=m���h��K�g?!�$��Ne��g���tі���V'!�$7�v�؀;Ӛh�Q~�!�D�o1.J�`�;;�\M	��*�!��:+���+�DԤ4�8]
��~c!�DRE1�� ��4*����w]!�$�$AңU�h� ��� @!��<���C��<��%���%WF!�M%c�`�R5���p�$b& W2!�d�B�X[�&��b�`ȸ1F��I2!�d�4k�Z����ۯu{d}�Ѥ�)!�䆚�JY��b��OdJP�qcſC!!��Q��Q	D��\W�� "���r!�� � S��T�D��$@ue]l��ڣ"O���7#��=��) aOOV�����"O����#Ċ���xpV�tn��"O�tK�
���3�)�`�kE"O���4Dڪ?����q��x���K�"Oh٫�i�|Yv2���I�4"O\�C�͜2)s4��(E�
�2"O��f �,	�,)1M�{T���"O4����I�����4�F�DT0칣"O���PP�>xH9�f�PK6ܘ�"O��C.�>�EsP�<IH�a"O�����ޣd��,���ؿN�Ѻ"O~!�1A��O'��*����1�"O�%��ՃY�DCpX�E�8���"O���.���s�c�7�d��0"O�<���D	�d�1�!�o|�ԁe"OX��G�.w���W��%v�,�"Oda���QrH9�7W.aj�R�"O��c B�f6a����L[R��&"O�5�� Z7ky�-�QeČw�:�@�"O�\#�#�s}j��&~v�e�G"O刓n̪f)���"h>��F"Oȉа��t8�3�Le꘥�7"O|I��J�� 	"�ҵc�"Olc���?flm腎M���]��"O��3wfEF�D���
LRdP�0"O8�r�J��5p�(S���߂T��"O$1�ۤ!��u�'�ϊ`И��"OhM�"KQ�Dq��ܠ ��"OJq�RA��|��1ڮ~�HzW"Ore����+�Đ�b�|lP"O�L�@+�g�z=��W�fEZ7�1D��`��)x�D̙���fhq�r�0D�"�#
�`8�P����K.D����"W@P�p���4)���6�+D�DX�c��<PD�.Y�j�P̹��.D����Ǚ& m��QPeC�1���+:D��)p,�(�"����[�wF�:�-7D�����0R}�}�-�c]0$r��3D�XH��ݔ@/D-�c�"��=�e0D��{���9�`�'�?V��i�T�/D��1g� t�D%K3-X!u,ƥ�/D�|y��-.x����"y��[M"D���琎	�����yj���>D����ϝ�+~��jE�ɫ!�P��a	;D����);v܀��F�{��x
��=D��פԪ@����F36��[W�:D������
��\��H['d�u�-D��bSOZ��X��F�w�P�w�'D�lq�$T�:��ZB�¡?!�LpQ�0D����*�&� �m�4y�=GH+D�����͙L�H�9� Uo���zqO;D���t��33�d�+Q%��b+9D�T1�!D�[���v-]P���4*2D�۠�#tV���E߳
p����#D��tȓ�KJ���sMZ�	�$$D�����.��đ�C�ZIP�I-D�h��Ŕ�S.]i�)M,Tɳ֨*D�@�)fVB���j -�<��+(D�� ��uW
��H)��H�!D�tSɏ�$�T�aҲR�����
+D�`�' ��	ؘ�$b�@�H�U�#D�H+@�ՙQ)l��7a�#��}�c' D��)��R� �eE!`9�i��<D�� ��sU#U�7e��v�� S>��3"O�12Ģ |S<�[�c�J���d"O,%���M"�t�"���KN*��"O0D�eIɊPR�0J���\�>��V"O�A��ـO��x���%SzHuBw"O6c$�@�U��U�d�N�u:n��b"O�耶��oF�)f��_3j��R"ONtk�$�r+�� �ʘ +��E"O�c@�S4#w���"��@�A"OޑQd'�� ��E��#�<D���"Op�G��;&�tw��fX��&"O���bJݺR�4��W�J����"O�UѲ(��7��֎� ���IB"O��q7f_.� �$n�1��� "OZ���ͯ5�!ٷ�=8�~<�T"OjH1"�	� �)5���&��y�"O� �"��%S�A�H�)'҈�a"O`9g����%�֬&%����"O�pBQ"G9D*�9���P;�m�A"Ox�'�$# �8ċ��.���"O\�8D��U~6U��(=o��p&"Oh� ,�6�
$�PLl�ct"O*x۳�E�A�v�#$1MHe#`"Ov�Z$�
�e
5m��43�C�"O|5R6cs�T�@��Ηe���B"O
	qb��9�4���W���	�'򚸒�_,f)�4�1� O��p	�'�@��7s�  pGO�N�,� 	�'��Q�r�\�������v�콛�'�� ���!l��EHd���{
>�A�'��8�f�`+:Irf�JN��'1*5#���$]��t��h�X�
��'AD���Ʈ7>� S�1<���'?,�$&�꜂�G
@_V�#�'7P�0��{d�5I��4���'0�)1IPk�e�F$Z�`r�'�0$�M#_� E���&���0�'��}�r/K�$dn!Q��P���9�'>=wО)��Y�`c8}� ��'#*��Ũ	�Č�U!F(r�`�J�'����
�re�ċϭ;��x��'U��f,Ҝ~FH�K��F�/��Q�'�@�Q�M�`?@����&�L��')��y�F�s
&i�0������'��\��`�U%v@`���l�- �'9� ��f�&M���������
�'�`js���cd��q&�%��=��'�t�%���[N�11L��:�`�'���k��j�.H��!ކ*��I�'���A�̩nc���/Z1"�,[�'ޘ�c���)�bp��K�: ����'���7���$]C��;re�p��'�z(�c���Ќ�p���0��'�0�y����ƥ�k�,�X�j�'V ��c`R+c�4i�F'�>q����'fd�b+I��sF�Ҧ>�8���'w�t��f�Qu�����.t�|X�'WЩr�kV�I����֠Z'���	�'�,��*�Um���$T���b	�'c 5�l���=X�-�
\�H��	�'�"�
�������c�Ҝc�8C�'zB���,M��5�r_%NpM`�'�re��!F�.�R�ۡ�gV����'`����A�bVpɖ�Rn�Q��� �0�2���d�F-U����"OJ����4v�j8�4mO:1׮%��"ONq*��5����푂OӞ�Z"O������?v�ty򡦑�(�^�8!"O<-�$��Z V��G�W����4"O�<�aC��O3��HGaO���R�"O6X3�T��vjȺWT���1Cɥ�y��]�tc���o�"u������y2��<gU��`�
	4��IC��2�yb�rtV�S���j�԰�C��y�`����0�+[�ZM���I��yB!�3�(a+�DֺfuB��C�y"/A=d���a ��t���Ae�)�y⎈<s������ep,Q�NR��yHל!�Ƹp��ߌe�hp�-�+�yBȂ_�@��	��]0�͚�dO�yBĀsV�[��0���
�t�!�D	�jV��s׃H��.\y�F)#�!�D��#�p�k����$�@KԒM!�č�d�x܃r��"pi� @��ԟ,.!�$�75h��*S�o}����I�!򤕬S��9�7�FcuH$3��!�d-D���r0�Z�d\��;�	� �!�d�-f�$b�Q*R\|���g!���.F� ���A�I���0�"�!�d�!z���[D�H]����t�Fx�!�dÐ0�l�t$C�8xм�Ԫl�!�ǎbj��K�!ɤuT�!q��k!�DP*
ʄ�22mܙWL�书�9!���kU+��#��2+ʵ�!�Ė,:���A��jb�Pc&�	%�!��_�Ga6�#C�xU���3�&/<!�$�6��3!M�6P��$X=�!��O�
�|�uiK�2�h�B��0[�!�d�>�zIQ�fQ<aT=!4+��M!�d3l����(	�%"�!�P�X�b�!��#s������j�,j4��N^!��2~j�k�,��Q1�]I��(I!�ĝ7�Xm�Ëњ�a����!�䖕<�<9�?T��|IU��72�!�Ď
[;�e��ѳF�By�4�I�5�!�Ď�1�u ��>� �Is䓫Q�!��Ƅ1�c��U�h/ Q��lU:\�!�$ܼ91v��#�h��웰%��*�!�ތl}$\XGe�	q�|����!�dY
4� )���ψ"w"�s�D�Q�!��DӓDZ�;}ޭ��h�)u!� �D��%f��;�ș�]�!�� �{���x��be���F�Q!��z�x�hen4pcjE���]�::!�D�?"��:o�k����T!D !�d�=[{H���lB�4���ʷa��!�O�I����
� ��� �I4!��LP���)J6��� OOD1!�ݙ8j&<��E(���.M2"!�D��d��kC  �Y�t=H���!�T����S�DlښR�bQ�!�$6R?2���G�5� ���(Lf�!�d���<!;���'����P%?�!�#w 	��M��^��]��ͰR�!�dT�a�<j��M=t
��Bg�8L�!�$\�yK���fQG�$�8���&f�!��Ζ��@	���Hjw�P�!��*�ځ�E�M%"p����C�%�!�� }�wNL?L}p'��o8PՃ�"OF"�bQ6$B���CY&J3�@�V"OZ�hG 4J��t`'(H'dfl`!"OLx�@���P$�"���#ꜱ3q"O�AAt�@�I&��B��ρe��A�R"Ozy�R�}��AQ���ʲ��	v�<�S� %g
�=�7HS�`m��[��LV�<�5˔�O>�KN�����O�<�uiU�Dp���/��1��fA�<15+�u���K���Ar��`D. H�<�sc�C�<a�tB�;����B�<	�G�r�*�pf�D�I}j����@�<�2��4TP��G'L�x���;6��`�<���I�4ʸ��5,՘.�|�IH`�<yQ%E0AcL͉�	`�u#�q�<a�
*t���q5JϗY��<C&c[t�<	��O�y������;����Kq�<)������h.�T��I\C�<)��G�*Bhj��7|{��� �@�<��#YL��K�
G��Nx�B�[v�<I���nT��Q��F)o��;� �u�<� ��%jt��H�J�zLY��H�<� �
@���.
%IQ�y��lF�<	s�՛,nc��$:�X��f�w�<�U�h�JTI�U&�$@��jZ�<I���54LC��v֌=��MT�<A1E@�Mf P���N��0*rg S�<i08K��R+^�[mXY�����{�8	R�*/p=��H�>Y��ȓp��Pc����
TI�>Qm�\��f��C�Ý>V�,�(�dF�sZR�ȓa�������uG~<� (|2����Z�9�3YjHĸb%�$��Ѕ�p��)���x�&����ȓrv�2�CP��:���}�q�ȓ-�� ; �9)9Q�8e&�T�ȓ{}܌�&UM�F���:\�ȓo�<�"`N�RL�$A���T���Ki��c �	IZl�07
�)) -��v0 ���x�ܤX�d�$k%܇�E�ɚv�DV�A���-v(-�ȓ<�Ơ�!��		�Lx� V�FA@9�ȓ_|������7T�h��NT�n�橇�%|�;E+ǀq���S����k�J���i&�h�R�W�l� �[Ǩ�6~��م�_gx���h��((r��ͅ�gn�)���ߟ���`Ė+YU� ��3�2U)P�άv�����ʰ*L��#n\ k�X$��{��ȓp1Ԝ�c� �2�Q M�>�P�ȓC�8�2�[���I��=�f��ȓa.ļ�A��X]����Ϟ�z"�ȓ�:�k���BL���c�&Jq�ȓ{���c�'��\0����Ϡu/6B剶If���!�� Ɉ�Q�Y�+��C�	cu��IP럏l�с�nX�B�0D�s��2n�К0 Q�	k.7�PZ�<q��F���ݙ"� &����W�<����>�LL�3�P1��V�<!���K���Ye
֑$�)⤋�K�<���N'��
�kL.a�R$�E�<��cL�u����!G(U���Q�<�cN�	�h-�0d	mx�7d�o�<a�NU R)��: ���2 �Sa�<� <!eG۔m�����j�G��u�"Ox�I�E10~�ij�+�38Ĩ��"O"���-WS�`��F��l#`�
D"O�KDg��=� �Y�]�a�7"O�}h���Zְ�L-0�B�R4�yr�Z,�0H�a�˅o�J����y2��Z�D��d b�����Z%�y�HITH�Ȁi�p+�+˃�y�J��oN�b#�U�K:61�v�+�yr�܎B9���'AȜ[6@j�D �yr�8v°�F�%[F�P��"�y*�ru�U���Wv��R����y"�RL��8c�W9���Q]$�y!�M�x�6m^P0�n
��y2 
?IӤ# �ߚ9
�� V�M5�y�]�!kf��<5�N�a�*��y���z2ሓk�.�,�d���yrc�$_�&0��EʏԜQ����y"D�+�T`�ę�ed옡f	��yRe9�1Sԉ�+}z�ñ�H.�y+/��|p#�0p5�T���ލ�y�'xll
%f�S#���^6�yb�,:?&�!§�c��Q���)�y���V�Us
֙Y44tc�A���y2j�<��1�a��zA��r�o
��y�GU!芀�����w��\7�Z6�y�(��eQ$�)}�*d��@��yR�	"��53S喻*�ʐ���I�y�j
,R��¢�t>�y��,���yBL��E!TN�(���r����y"�
[ܮ\� ��&EbL�#gۻ�yB��Mmy*��l4d`:ăE��y��ϭ4���'�B�;�����y"��(��8� �S; �z\z�͖�y��&b:���^t�C��^��yҢ��j���|�а�D��yB��d��l��(C�IR m�s�æ�y���+�|y��=<�ޑ��E4�yb&L�1#f�q!�8n����Ԃ�yri�6@̺�
Ο7�Ҭ��G��yk�]���i7&D7{|3����ybH�w���V�Z�;!��t���y҇;�IH�]*�:�����yrN�r�0K+y��|Y@�:�y�l	�9��]8�i��<�(�*�yL��l�V=��/	m�lҷ)Ȗ�y2�C�` ��c��6�:`���5�y��ul05!ֹ&bJ��ς�yb�"�0�b�"S�P��Ty4���y�F[�q���+���H�����;�y�t�ĉ�e��;c~�зm���yꊷ'f�����և:Q>�Z���y��/@N���=9��t3Bo��yr
�9>��<aF*��0@�zQ�H�y�jF/;:�{G�G�Zh�x��yR�" ���FU�K�`�c�^�[�@B��!u�J壢�Ixj����2�B�	��&��F�~�촂��\�C�	�8A)�#���xA��M�ou�C�ɕڶA��(hG�!�˻;��C�ɓx:�A�D/6ut�갃� !�@B�
�t�:%i֟�RA0�B�!��C䉞R :Đ'D��Hy@1&Uf;�C�	+s2j<6��"�<�X�i�0W�nC�)� ؠ�����V��	��1j�
D�"O��AFI�$�Aף�1�l�hp"OP��$.������"O^�(��E-~�x�t��R�����"O���RiX��	2%*L$^x�\�a"O�1'���6IP� ��L8��"O�P�7�Y�� 8æ��uX�"O��`��[�G�(,g��$ 8IkW"O��K ��7��uA���Qp���"O.�9��,0�����kVl�B�"On��$A�/'Z�5j�̂�,^0��"O�i�#�H(��{�j֐9Vx���"O~l�ѩ�0������Ƅ=P}��"O,2���� ���N�U�<� "OM2%�\�8�����%7&\!�'�41�'M�+Bp��=�ʤ��'����C%N�cSr4����:Ťu	�'�D����_��vI��N 7m��Q	�'���"�ؾq�}���$B����'�Y��*ś,fB9趋�c�Z��'�P *�NQ��Es�֍X�����'�+!M�Z\<�2���NČ� �'�ؙZ!.ݻ����̙0P?�,��'�ri�@�<[�x��c�,B��|�yr�'��e�党rX���E�8�,#
�'�:���h�u����J�+���
�'*��TO� ˬ�*� �r>�`�	�'Ep�s��0:�D��h�J��i	�'
���
�!a�����ԉux�9�'̖�8u�8�cDL�{�5��'���VkQ��i�e#n��%c�l���'�Q���'�hy(t�D;Z^��"\���	�'H�4�k�7���f�K[�`��	�'3]:�kâY)JD�U��~�ֈp����?�u!ˀ=t޽3�NB(b3�s�k�d�'�ay��N�f.$���n�;B��X�f���yb+(SX耠B<#f�+E����>)�O഻d(ƅ3'�ᨔ�X����Y�"O�T`ذ+<<��W�Qc*�3"O�6LڡL�}�4�� ���2�"O�р����֬���N��A���IF����A�Z%������q얡�d�G�]�!��W�@@U�܊]�6`g���!�� �W�&T�
΋"�a�gm	J�"Q!�"O��:r�0#��x&.��"���q��I�<��)^4}�DE�$DU//��芳虌5�a{2��C3e��Q����~�{S��b���hO��lJv��Tu��R�� $@���!�S�n��)(�oB�i�v	����"�����	[����O�rB)��n\�����&p�u&��Aj��G�'�PJ� $>�@�6��yV���	ߓ٘'��Z�ǁ=A��q6�T�xh��!�i7Bb���S�O��Y*�m�b*9Ye![�rrbı	�'ΌaIg$@-"G�% u䜷~���	�'�:!2F_���(*#A�9���'��O��b�G�s����F�7�*h��"O,�JV��>�θ���ƨn{N�b"O4����D/s�h��W.4\��9&O�����	��$`�,[c��吓�X"	��xǖl�'�:�@�L7����`D+`6D�
�'���lS�
�:�Y�R �XM>���iA)d��-��=eB���(G*��IW�'�?!�f�1o�XH�$�JP!"��*�<�O�����E�6������r�Q9E�=U�!�� ���c�]+V��� �F16��"f"Oh��"m��1ᤚ�3��� 0On��dJ!/���3^%�v����ZF�!��T�-h<�� mZ��1�a���Q��F{*��Ԁ�T6�`�kW��8J&*p
�"O���陣B*��-�7���3O�=E�DM-z΄X�J��d�\�:��/�yI�#ژJFd\�\
���j��yBaݑ4\����K
��H��I�0>�O>�7"�2��4x�$G�J4�4�G~�<As'W"B�Ĉ7���r���a�r�<����L�,���c�
�*��Kn�<I���1��؂������BԂt��eE��j�ß� �z؂��>b�<��ȓL��ܘ��̙N2�J�F9=bʕ�Ɠ5���mn6JM�1���j�$�+Ot�䘧(��8:&�,R�Q������ "Ox]��ƾ�6%�֌��:�܈��"O�=(c��ȤC�k˷~D �z�"�Z����r �~Z����o������ڧ�y��^����wFP�i�>(�/Q"�y"�:=�Uೇ��KPt��� 	"�!�(D	@�k�˚������w�ɠ>
�me��-��r�%^�eM(B��$,+���KAf���RB�I�"��lr�];4�d��*Β)�B䉋�|�W�"K�J�r���E�B�	
:�����.m�P�`�kdB�ɟ$E$*sd0U^��4fE.�<B�	�(Flycw �'w-Ҭ�Í��`
0��Ɠcf��!���U62H����.����38�x��->�.X��.�"|���A��@�aΘ-?�.MRǋH�Ҹ�ȓv- ]�a+W�e�@�v唜d.����O�8E��	,�B\:!���OqD{��T"De���'��=��¢R�yr��0a� A�'D��WR���o����D.�O�5��c�t�V6.A�0V�8���:ړ�0|�t���р�ᆌO ��`��K]�<y���$z��[s��s��H�2��A�<��]��i�%fF<V XEM@�<A�h�F�lؓ��3@�J)C�[}�<�%��<���gA�S�2�
&��v�<Y����0L8ȳ�U�iji��q�<ٗ@��/�p�J ��9���� i�<��ȗ�9�fl��� =��;��a�<��B	 w��Jfc�>SR�s��hH<9 `_V����G�jP���'�� �!�dؠ)ܦAk�56��9ku�B�b��'�a|«K�D�R#M��1��5���y2j��JP��I�->a&Y����y��\�� %�ĩ�~���(PCO$�yr��~�(��qh*r�U�W�C��yR�d�X���+Y�.p3����?�f�h���G$��'�?��H���ũ�D(Yu�I��I?D�h:�#�wv��G�S�d]x��ǭ>�d'���~R�j��U	�
L���Px""2��ٱ"O�-eR%�@��(fv\�ӓ�'�ܢ<ikZGsHBb5:ЪX�t'�\�'3ў�0jj��@͎N\���앪l�pA+�'�&a��	osp ���Zx�n0��'l�x07튘St%��C[�oh�	��'_�Ɂ!�����2�N��}�x�K<я��)P P#�Сc��Ex�!����*I!�� ���2ڀ7��������*�JE�)�S�S+8�\s��� 3�&���ډP�B䉪lk(�+��U�*���e�>5ʮB�*$	�t�*�1"���A���B�	,G@l�w%ڪbǒ��d�)h~hB�	�Z�ĈUa(>�>,'W��,B䉐qB ��I��q�� A#��,�B�	$[L��A��
��pp��&XT�C�I�����a+�=�Đ�ɒ�e��C�ək4�H��G��Y�K��Rϒ#=y�$q��j�ς�7/&	�Woߣ/�u�ȓq����k�NB.p�3h���E��/�]$�>�H
r"ӛL	��i0.ec���벰)��[�HK�ć��K���D��)Dsv4�R�E7zxC�	*Fh
A+�S�xyZl)�HE1C�� q9�(T&יL@�
aꝌe�:B�I*V� ���'G�P�QҎW�7�C䉎H��� @O�hc�˓�f󂼅ƓD�A��6��@@�n�V�t��	I�p��Y�r
ݮ|������ $�͇�l!��aW���=P�#�d�Ň�R��̰�F�~�YÅ�J�9K����&``��_�1(8`c�?�8�ȓ5�����Y1xl
t
�d�ȓ/�,{�h^~�H�z�*T�I�`5�ȓq�N��'Ό%���Z0L]9%���Qj�K�
1������	�Z���DZ�[6犹E������ap6���=*l�:�LF��mX�H\�z�*��ȓ#!�LI�ǻEZ���ԏ�@��ȓ|��z��9T<�� ���9�~)�ȓI>i
1�[�2�X �Շ��g/\!�ȓ$xAa�ύ9��Y���Xޕ�ȓh�|ǆ�J��hqt��_�ІȓI	��8T���n��f�))����f>�h��GP�p0�ߧ��k�'� �J�r5^�@����B�xi�':�	ɲ��S��$�G價d���
�'�,���A+6����,.D�-�
�'�Ȕ⤧GA��������'�H��fʘ#G���S@K>~�0C�'�|��K�*|4�+�͏z<uB�'<�����ۻq�8��D��q�|��'�1�!BoT��D�Q�oVR��'�ވ3�Ѱ"&���f�(X�����'��X�- !Q�i�Ư�IҘ�'���!�vkbp���DF5j�'���1ä�U���1�9a�D��'����fH�7���� e��	V��
�';���F��;
�����ŗeLЃ
�'#d���
�Y���F�O�v��4��'�6�8�i�>^�*٩V��z0@�'����C �3s���pE�%�1��'"2!�c>^'@iX���
�q��'7~`I'I
w��y��N1~-����'�@Q�Rf^9�V�_:{h��`�'�2L����{��H梁�z&u��'��YXR��`δt�̣rnYx�'�ؼ�cL�� ��ق��(�i#�'�Și��ܹ�T�Q,���|3�'s��aJ�cC8��q-V�H�@�'bB5j'�ތI��#a̎9i�x��'8&�J��K-o��2tG�+i�
�`��� "�s c���  �S��ξ�zv"O�MC��Z�mk~@ ��(�ԙ�T"Oਲ਼�W9\.l���Q~� �2�"O��挄�H���!ড়n� d�F"Oh�Y��ބA����B��Rz`��G"O�L���G�u�z�xtO��qX�Y��"O�=�Q��xΒ<+��ْ<kl%��"O�̝����!^��@"O��gdУqD8���
7R�,��"O~}a`̑���x�gO�4@Ѐ�a"O��c�%v�U�VF�%?��IB"O���>?"ޡ� �U|�V"O�P�A��XD�a���U��r�"Op��p�=9x4!�+�6:�J)�"O@�å�'U������K���"O�-y��( �1hg�Rʦ�U�<	 f�bMJ����&Y.�a���M�<�-�y��˓%�,j
QA�˄]�<хf�$��h;נީ[Sh��D�WX�<��ǅ#5�9B�3x1�q1V 
O�<	wmK����g�. ��YRD�<��S&~zȲ�O�0H�m�T'��<Qp�2U�j��%�,q2�����v�<A�E2u6����2�4i ���j�<y�cc.a����&b���%�g�<���Z�c�1x�~5��R��c�<������$��M\02�p
�Y�<A�j� h0<�qG#�
z_ptCLOT�<�&�^O�i�֧�������T~<���M�p��V�
��~Ř���<[�(��[�N�SCG
C9�� ��)M��YG~b�S??�n80Ą΅2FԸ��T�F��C�g}�]��*fe���$A�,B䉎�И+�m�8,$�	{�iΈq3�C�'X_��ж�EOL�U�Ek��,50C�IR#�m�B�q����!� �C��/�\r௚��X�q�B�ɳbd �n��{���*�4\"�C䉼F]�]S3�I3<�8��'��96�C�	I���h��h���Y�R�DC�ɷ,B���e�
�P�ؼ�u��B�	Md�QC���5��\�R���C�	R3�m�$
$<���2�"5m�6C�	�R���Z�'߶H̞�01oQh� C��,o�� �(O��h�8F
�P�B䉑e����~׆ K���>>�TC䉳Q�ihP��5J�p��	��qv�B�	{�ܵZuk0�R<�%l^�<�B�*]2 Ar/."���QCQv{�B�!�<(I4�h��ag�PQ�'D��B��Œ+������ͮ��q3c#D��(pM���(��p��A�e� D�`(�z��ԋ��I6Sf��u�%D�P3o�<|���n�4eF���'D���4�&U���G�_AB�!�'c7D���b�νd�pᣠ]b1`��qm5D�(�c*k ���tO�X\H��5D�x�'�In��R�ͬ&(�0!a�g�<1#�	�q���cq�֫x��c��y�<�ɕ�"\����äl0���c�z�<a�`N/-�X�ؕ�A8@�������r�<��AF���q4.^7;g�t�cu�<a�����l�ʓ�ۻ^q�ł���d�<17�׹8BI��G�� f� A��Yi�<� ��t�]�M�b�@C��5l����"OTY��O���]<Poޘؗ"O�A��gL'���	ϦX����w"O����A	
B��P��h٭o��xh "O�L��#iRX��@S���1c"Ob h���h����-���Q"O���l�)��b-�C��U9w"OL}˴��fp�-E&��a�"O�TB�C;[0ƩY6k�'3s.��7�	�KʖmH��	^M!�0�A�T���W�A�*�!�Ą�]\Pi�GK���%���D*q��ʻ?X$⟢}��^]rj�F�33�@���"�`�<a�LW7�&����[�F�@�c#�X��7.������0Z�&!JR
�)v4NtkWŀwd!𤙰Z�Z<``�e�����@��#y�q��E�R�Rfk)�O�1�T
(<� �bD��VS�{�"O���R(E�%"��9LtZ�"O�1�Ń�%�\���>�� �"O&���CD!j�U[��?D��"O�Z�[$3p�2�l͏#hi�"O���@��':
t���;*`��"O>�3�OQ(r^��`��$b���"OFh�wCJ�(��[��Ĺ;P!"O�$(!�!�*��k�T�8;�"O�T�ש�U�Œ�H�POb\�B"Ofi:CE�BVt��*�!P��)�"O���"�(_H���[�i�SK��`&!��W9L2	�&K-<=hz��$�!��N/{�"e�5/	�z?��� I�\!��Y�7-�)����@����$�Y�.R!��̈N��[&%ˢ�L�R��&�!���]E�hJ0�� &�d�1�
�`�!���w�b`c�.�;g�]�d�!��C!�҄��6^V�"1h׌E�!�D^�b�Fq+E!�l!A��
!�D��"q�����a��(���!�D������X��&�@v晇h�!��׿y��@�ݼO��=�p�Yr�!�DK:]�&�q�)t/�D�d/D��!�0���a��[,t�*x�C���F�!��7���c6,�}�n�q�M�.t!�D͠x�^D�rJ�Vu���+R���'K��˅XVF	0���UL"��'��Qb �{\j0���R�%z����'�����Z�(�8�1��� 2ڡ)�'���k�J(~};���_G/�9V�➄G��'Sʜ�1ȑ���hQ��b��E��'�&x�4B�/sv�q!�'_#jD$O�N ��*�!W��0>�(T�%g��` �R�^��D���ux��h 撀\��T���x���A #^a����U���HpD���y��:Q7b:���r�|�X�(N��ēQ�P���$�Z�q���(�4�AA���%�R)`4"ܕt��\Cu"O����-?~���*s>=�xb�9,޾��G�.�?�s
ǡF���'��k H�@Y~��fy�VI�'��9B�̤E� 	ɱNJ�MT��6��#��P����p�����6�E�Hq�M���˿F��m��e*O&�yg���+��'��*s��i���u��ʕ�����hʬ�y�dL�"����$�$������V����ɤ	LjUa���/3���i!Dߒ U��?Ѩ �R�e%=,�� ��dN:D�0��f��I�����&T�8�e�a�ّc��Ȅ(Y�kDU���ߗ�c>Q$�в��T:Xk�ARĥ��!e�5��*�Ԫ�A705V���Bϫs�&�+b패R�lC��+\&�b7j�; �Ȍ�OH�9�.4�IQ�ec3%X��R��A#V�8��ۛ+��d�'��m� �ZDA�)�ʸRT���y��p� �@�N��8�0�,?�$� s�.��?� @u{7�U4XQ+1�7K=��KR�����<k�lLYw+k�����Fk��p�����Z}IB��`� ��u�=) F��@Ӽ��O�D`n� bM*Z;,-���9F��4+ĆW�$�������	�+��t��s�&��
6�`w�?vjM"�`�F���� �'WNE���]�Y1�`x�aO=5p#@KC	�uҵC���kc'1��I
.2����d�� �I�M�v ,,�6b��x�F�֡��Z�\�r��-CHF��d�-��S�؁�
h�O�1�'G�����O����ǩN8E��\�v$	0p�Z(J���mc���x�d�9\�0����,r&
�y��yL�h�ƚ��bb���&E�j8��JgN��̸{����l9H�)w!��ZpN�:F���V�Q�xb?OИz��Q��������Pq�O�HY��K�]�D"�'SDSN1�Q!�1$�����픡`x:yY�4\O ��G"���:��
�~����'���"�g��v���,�̦�Y%�B��P���b�>,�Di � 8D�$ڄ��p�h�AV�ԁyM�}�7'ȸ��KQ&_?��[3T�8h(���.a�1Ƨ&D�s��p�脑�if�}H�� 0��T�{��(��F����W���`��5�5D�����=s&u�VEݰ�dIA��2D����-'����]=�%&]��!��[��u�"�D@ؒ�!�>�!��
���E�5ve�� �N��!��M�z�:rI�- ��E,L�{�!�䚳&���K2�8��x��D8!�ٖWdtMs"�ޚEcF��5)B=h$!�$�}��n�GP�\QG�9w!�$�y����g���BÉ�!򄜽~�T Qo��s�D�G��V!�$(`'��r%J�}�>i�猯=�!��œ-vlB��G"0��Dr@F�I�!�䐤7����H5<_Dsu�P�g�!��!z�,̀#�X�|�t���lN�!�J�\&�MX��3zuJq�V����!��[�Ș��Z�Bf����2j�!��
ps0��E�S��sM��B�!���@m"�Ӧ.�$~&�˳Mٴ^!�Ą�Lն|�QJ< ���(��5LF!�����|��.QC���kԻI!���I�������*�6ĩj�}!�$�y��)�q,�.�ֵQ2I!�dM aZE�	Y|^��ʇK�!�dȉ@��,c�,O�R�d�q�)�!u�!� �7
���m�!NL��c��6�!�$�(^��W"Ժx+g��_'!�d�.<�&,Ҁ�ׁ���Y�GU. !�dX�{,��0��
3�X�kw�I�\!�R�^Ԡ)�b��Q�� ���q�!��-&t#%�[2XVԣ0&F�5�!�d��3�j�ѶeC)Y��10�D�!��%L"P�2��&@ y��d�^!�Dٗj*Ȉ���| 1� !��x�����b޵�̆�2�T��?�.���H^�X�)���:����2!�Ց$ǀ�װ+�Z2tVt͇�dh"p �h���Y��D�dPZ���b
5��V&b13h��WrF���O2�$HOϣe�|�ja$��2hR���SC��H!��AP\#�g\20�I�ȓzֲ0(��5���.YmJ���ȓXz>�Aց
8p�^t#0&��%HR5��o�(�7kD1��ZP�@�`vpC�Ʉҕm�P�m�호L���h�'\p�zBǎE�T�Z��D�@e
���'�B|�aO8~
���`��3m楛��� ��x��M�kH�{� �T��H��"OlUr�>�HX 3@�Oy��e"O䍐�G5-�l�`,Cb�ȳ�"O�(�5�;�f\+g�Ӆ$l6�+�"O�q�+�r�3KC�`#���p"O�̉��־T*�H�1�9��"O�!��I(J�p���S{.�C6"O�9���g���W��(���"Od��
�*��� 83��A"O�a�����Hj�Ǚqj@5��"O�q*1e��ƈ]V���W"O�X����N�FD����L���r"O�3��ֲim$��F�U�Q�ș�"O�m	r���`עY��#q��V"OQ���Ś6��Qv�mb����"OP�qAI��6�S���3xBX1i�"O��c@���-��Ż%�):ʠi�"O�]b��P��R��E�i;�h�g"Oᘇˎ�D��Q��� '$P�"O�e���P�v@a�㍬2X��#"OVt�!!��,h+/����M#"O�h�r�B*^'����OE,wV�z&"O��R�N�]b���I����c"O ��ìH� 7�ih�G��~vP0k�"O�͸2a�����S$�G�wO2�p�"O�|��JWWj�l�#,�5998�"Oʀ[oK
 �N�Z�N�/%Z@ZC"O��ۆK��a鈐J[�Hv��j�"O@�äVfƒA�≞�]�@s"O�dy���\3��֧h��mzc"Oٲ�lS�	uj�ٲeM�i�q�"O����#����ń��y�A"O6��o:H�~��B��F��Y("O$H����%� 8�T�U�%���P�"O���ᒍi`�1 �X�Z��i��"O�8��$�9X˶�0���#Q�N`C�"O�c�N���C��"\�P��p"OL�P��?'����@��h��pp"O����a �lPE�:r:Hk�"O�x��՘D�T@-чqƘ�9�"O��"`KB�D���3i̙+�R-��"Od1��dA5�𝩷.������"O
���K�T��9��BF}3�"O�)����L� 2,۳c��MkR"O4|�beӐ0FDM`ҬJ�D�f���"O�@��K[tX]���G0=tΥX�"ODـ6��
:8�/qݦ���Β�ybMO�y�&��-ߔ]�~s�,�y2���I]|�k�i�,x'DDڲ���y�gنdJ��؅��s���3.��y�˄� ���mߗn д4=�yB�	/s���$nE�bt�x[sDO��y2���p9B2M�K�(��Gė��y �����)6}��ڧ��:#t��'c��DǛ�y0��BPa�8)y|�'�x���
� ܚDa�\�az�'�x�*��#�2L��nZR�z���'�>U�� ��uify�c��6U%� [�'�ڄ�H3s�����G3�	A�'��q12n�8�-0p3��3I�
�''�Tj&��@#R�*��J �ū�'�&\q���58Kr�W"a�^�	�'�T��C��%���?[y�i��'��(���#إ�ԧQǞ�
��� ��5�֥B�t��"/�2>���"OR��1fO�4�|e�l�ˢ�)a"O�!(%��j� �Kc�'|��mX�"O���&C��x��ƢH�9��(P"O±�����B z���&8�J|h"O" i��z��B� S�:��ESP"O�u	�(͞{)�,;���w(���"O S�K��T�Aa�	�7X�e"O��4G~� ���ޫr�p�@"O�dBcXN@AI^��p��"O��xe�g���0�P4����s"O0Ls������`�P<;��Z�"O��Ssl��zX��?Ez��a"Oe��	�Y6|�z�XBC�!�%"O0|�ԍ���hUI�	k��/�y�j�,jd�(D�j��.@%�y�␋D��sF1ad�Y3	ַ�y���*�(
�m��`SƝ��y�-6g:��� $s
[��M��y��$ΜAK'��`��Ĩg*��yr�V�o�����#i6X`w��y��8y�t�
��Ȏnۈa��_4�y� J% z I�c�΀S!��UkJ��yA�s`-j���22A�d�K��y���1b�����3�\8A�[��ym�|��u�И"�i���yR���"�\�g�J3#h.��Ү���y��1A �ВE5 �pظ���y�����R�ot}��@��yb��81�̕%k
�{L��g!�y�,�/0�$Q�����T*E(�y�!�\\��(ڔ��EF��y���-*��c�j$�L���k@��yRc�h�p�n��-���`�aB��y��@-J�ҩ{�H��@���3�K1�y���#���m+N.FX��0w��;�y�bH�B��6E�8!��:7A�y"��2�����"FqK&��\��y2��2��Eg\6v <�E.L��yr������dP_���ڒ�˼�y�'��t͒����X�y�A ���y2/�(fR��.��{#($��]4�yR�	X�B���#{]N��2ň��y�'G*�x�z���w�bĠdd^�y�T8nת�ٰnP�t��9�#V:�y�M�
r�"��o�~��Jޮ�yr-�b�P�
`$�:^�(x�bR�yR�RE(h���C�Phq"n�*�yZ%�h�03Nŉn�<E�;9��C��&�d���Y#�,Yk�D%E�C�'j8���$ׄ��z��$BX@C�.e����Lǻ���#��M\�B䉐3A�0�5��t$>���g�B�I[a�Ճ��U�B��*Q eC�2x�3c�/q��9Ye
�^�XC�ɀM�\Z��3��mpԩD�P
C�	�Wj�ؘ����zt�ÑHy\�B�>^��t�@�\�3��mC� n�B��E�$p����>T��"A�~�xC�I��V� ��
�8��ܽRGC䉊t�jT���2F������\�&�C�fD���2���0Ԉ�c�g�hB�	���d�<X�$`�@mY�I��C�I�L��	#�W&4�Z@��D  Z�NC�)� 2cP͝HV�����F�	�r� �"O��:5
W�#�m�>zs"OV+!�ڲy�pU���S��X�U"O��9$�Ŀ"�2����.b�����"O�8�q�9���X���%��� !"O0-`g! ;<�i$�M��y�"O����n)�(�\1M>l��t"O��8�lʔ8��S׃�+<yx�"O�1x,�r��D��I��c>�x`"O��"���n������w
z��"O�p���Ӭ�L@ig��	b��"OR��� �8R��M0��X����q"Oެѓ�M��9�EJ�qվ�#�"O6 RC��{����eܐZ�N�q"O��A 	V�H��#FBU:2�l��"O�i���U&b�N4S�!�i��5s�"OиIg�D�mf���d�&6�e#"O�8�d�%~`�kO� U�t"OT�˒� NH\a0eo�>^Ұ<a"O�ԣ偈�-�,q0�F���"Ox�0��ϑX��䫡�W�p2"O�L�%K՘,� �[VCT�A��A��"O�)� ݾ[��Tڦ)"���"O�� JTv��h��{�l� u"Ora��C"0�$��q&�9!�j�s�"O��hs����q�[lM�U��"OL� �)]fv Cr�V��켚�"O��BJl�hT��DP��Q��"O��j��U�-.�4# �hؔ"O.|���fA��B�MT?}c�ұ"O|d�m�ʜ�#�AOh���s"Op�"�A�'����F@/)��[�"O��PbN]�t ��eX�Ux�(z"OJi�/OG�.A��	P"5d!*V"Ob�+�2#j�� R
�}n6	H�"O8̸��*i۔��h^�dC���"Oj�ɐ�'����Q� "��9�"O��r�";ztXd��!��"O���i�-�Ƅc�O�>Z�x�d"O�ig��yqV,���[. �t���"O��9���,H�k�(X�R�S�"O�T�-B���9s�^#7�����"O�X"����D��6�S��ea�"O��G22~���E@�[/j�X"Or��)���P����9����"O�M)�fͼo:Ա����2�,�y�"Ot��wC��	�� E*C&��e�"O~�pweS]Zh	�/Λ ��p��"OU3��E	���C�Eh���I"O�-	�#ÜjT��N�a1BL��"O~��&I�5@�"<,��"Ox�H5��A�@	!ļY�tH�"O�M��L�5�4@�k�pT�"OHr�G�v��)�A��m����"OF���A��x�t�:� �9M'r�y�"O�ݐ5�H4>d���� J��y�K�U u�ǌĵo�q��]��y"M-,���q��]H��t���y�@ݭ?�0�(�H]Y�"�#�b��y@!?h���	�Y�B��Z��y���_���I`�V, _Ftbb�.�yrjW�3� ]s���wx����O��ybk��e}p)# )3g|���/=�y��-2D�+�mY	7��j����y
� �@�W�B���aD�I�h'"O�� �,Q�$����C�e���b"Oj����Ɏi5F̹��C<�ܕZ"O�%�.�&=�����o��������� l�'�v��}ӑ>�����ܠR��\�rn�)oz��'�0Ŝ.S߉'s���dE�qx� ۉ^�L2�Ƽ �BT��r7U�����<pa�B�Y?W���`e�%���b���<!��U<}��y�P&�"�H�4D[�)㛶O5�S�O�T����"}p0�`XDN��c9��0|� �1"a�0�k]�p���2f�@m���hO�'X�j�����Ga��2G!+X�Z�$��:���I�0�����g{0������E�'�Q>=�������N�f����5�v�4x����/$���8��β.�T@��G�]�@�Fy�	4���]�'M�]��N2�I��6{� ����L�� [�'��i��F���
�(���Ql�*l���m�Y���	b�T���l"��2$'�O�˓�~�'(��$�q�A2iʐ��
��k�.�p�L�>AS��>�p�	��H���(T���q�ٽ���Ni�@7͓��(O�?��beQ�tx��B�\Ĥ���Sk�'�8���/V� �%��
�Z�Ҏ:q��O��GzJ|��L�"I8�I�bQ>Np��{�	~���OY���Y,e*���:à=/O��=E�4�Ӷd�h��l1K:Ț�)��?A����x܌�2L�c|Xt�A��5{B�Dz��|Z��>0�zS�@ެL�F$�$��<	���p}""	e}���(���4(aK:	K +C�I�e���'��	X���[�O��]��!_��y���õea�С�U��X���=�)��srp�����n��r&�����FԼEGJ����ƻ�M뢁��6�|�"�YJ����R,_\����.���y��Ƈ@���!��@�q$*�!�y��&#���#��2y�F|@d�ê�y�Q4p�`j���>#�Djs�^��yҫ�"�uHE	6�Y{Uj���y�% �'L�*�
F�YxT�Ç�y�ˋa��9 $��L�s/���yR�52|1pm
�n�k�����yB�Y23zf�bw�@o62�M��y"$�*	�YY�[�0��Qb���y�E�'QT��b�]�#�tx�!ɚ��y���0�Q
V�ۨN�n9��j��y¨ζ"�m�tJ�/1q�������y��B/!w�B� �90v�y�����y"�W�f9�&K�U3��*��T��yr�	�R⼳,ƩQ�x��� ��y"��`�f����@EX������y���Q�FѠ��)>�l��d�=�y��j���s'��;r���dP�y�(��B�`������4�����y��z�x�b"�ƾ %�!�A\��yB�(IOɹ��;�a���Ѓ�y��ܧoFTQ˗)B��HA�0�yR!P9���B�ԏ{�p� ���yRcT'���bh�x�ؐ�w��y2gŪ?�Xѷ�E�вg$ɢ�yB#�!G�cp�
�"�!kƛ0�y�ޅ�ґG�>S��h ����y"�K�Yd,p��+AJ���q�)�yN�@��%@Z��Ĺ�����yb���T��ʥ]���x���ߗ�y��/a#b`����r����E��y"+,N����!�[�����b�'�ֵ됈P�,�p'h�1j��(�'�  *���a;�Xw!G�Lj�!�'^�t3fK�9~���#8N������� l� �7��� �G�p�ؕ�W"OD`f*@Pa8�A�:6W�H3"O�xӦ�!#����� &}=�5""O*8Po�\J6/�9~�-�w"O�q��zBbT�u�ȝ_��"Oz��uL+j/*l���	v�jp�2"O4=���Y�0���S�P�v�V��P"O�`)c�ֹU�2h��ʍ+�ĤYg"O�H` �Mxp=D��!�����"O� �WC��J5�䰧��><`"O
���şu�}X��7$,�C"O ��rmM�f������BZ��"ONX�$��x�2�Ӯ'��y��"O����O7�	��
�[��9�"O��r�O�%zD�qwig��yQ�"O�{���=�P0hU�O%����"O"��,��55 B�5�a"O �`�*�R�[r�+z���ر"O��qa�?7�r��tK�;Ǟ��"O��'� �P�	���@�:"Ov��ǆ�w���r�N8���"OJ@����m �*q�^xL�{�"O���ƎC	?�xl���\�,YV!!V"O��p��0P�`��h�@(%c�"O��	!I���	s�G�2O�p��*O�]Z'�����f��K�&C�'i>,H�mL(uwX�s&i��J��I	�'�Z���Hdkd5�&+�P�	�'7z�+��0��e1�B+{�ɳ	�'����l�/%f��4"69\8�'~��2�˰%�p��/[��L�'�L1�	q�0 ����bTU��'�h{�"�\�}���".X�S�'���:�`�4;`ab�K��,(� �',h�)��i���O@~�h�'��iȦπnvhb��A�]
H�`�'���0��3�V�ڶ��j�h���'��Xp�����80�K0!�4��'6l�����FH���u�5�h`K�'OH<�H�;�4C���u�R�'��������5���8��A	�'��Ǐ�|��<Q��X�D<��'�d�ӳ�D�w�1b0߶i̙�
�'X0���%y �������'6��ʍ0m ��e%��e`	�'�:̙f�e�0�x�蔥}~<x�'������\4c���?~N�H��'� �:V�?SV)90n�#�� �
�'ߖ��I]�g��� P��.!�"	"
�'��Dҡʕp6��0�2z�ջ�'��0I񣟅ZC��v�&�v��'Q
�6�%4ز�aG��-
HH���'�� ���@�f�#7�[�~3 C�'��D����%h�mɅY ulB�h�'���Ʀ���vA �A-n��#�' .�Iv�	P�0�Ýd���'H� 8Ed��%Q��@&�W[j���'�*�R����9�CG\\���'K4��0I��BO׋��4��y�a̍� pȶU=	`.8�����y����Z�z���N�3rf$P���˶�y���t�~���H��4��+Ņ�y�/ש7�+�A�=w��haS��y��|��[p�
5�����P��y
� Jx�G���l5�CӁ$GrP��"O����ݑ;<� J`��ڌ�aQ"Od��6d'3�����W-e�B�"O�pK1��$A� m��F��O�ȺV"O�`{��VF6��h�dM�JjlP��"OV�����1�����R�g?@db"OJy	���^T�-K�.Q�:,�<p�"O&�a���n�
�kF��:4.���"O$�I��Q�.l3��QT ���R"O0pJ��L�fx 4��8E#�@�e+D�t� �Z-|ۜ����*#���*O��ZE�%D��!I�<M�2���"Oh�KW����$��N�4�8Ԩ�"O��0@&��0�����&�x���"OR��	^�TA����v�p�"O����),��`�0������"O��e@I%06����Q2 "Oh�����MU���%z�,�Z�"O�,��E��(���뇣�4�:#"O�܊eGC���4�s���*#"O.���dة!;bD�!(�\����6"O5g$�^�Rax �_��5��"O`�`GG43��27�X=�V��"O���&L8R#�A*@�t�"��"Oj�X� ̜"T��f�\�dBX��"O�]� �<�x Q�̊8�HjE"O� �֯K!3eF��������|�<馫�b�d��E틢�%��{�C�IgbPOU:� �bB��W�PC�I��2X��+��<��<�E�_�~fB�	47����A1�\ї���dB�	8�QT/� ,".�ȑ'Z�A�C��*hA��A!{�4=S �6CH�B���!��I	��t� $�9t�B�	�Q2��j$I�7�XtJC�H6Z�0C�:Q�j� U�P"	T�ق�X�C�	�36���r��1
6H��I-5~,B�	�[e�@:�Nҋ�Q�s	|�C�ɟ /�ش푯2	܁3g/�7��C��({ǎg�W�����B���B�	&�f��4Aʜk����S�3t^C�Io������	��2�]�d��B�I.,BL�d
�4�ɱm��tB䉨� i!"+�4�
9�si�38�B�I\ڼ��k�3T8��3cǵ0��B�I�Ѵ��1�1�T��L�o�JC�əi��-b��i�ܐ#D���!&C�	�����4���9�I_�DC�	�W���q�N�]F�����z]8C��/p�<yҰ�r�T,8te[�U�C�	������ B�6�+���	��B�ɉ\'b�K����{?D�`�E50B�I��8�ц�1`� )jt
7 ��C�6p�r�'�[52L3e��0<̐C�	�ic�5)��һTs"�@%#�7h�C�/�܌xA�n�� ��& �XB�	>lB�(�U	=ĽqC��*WD4B�I&&���nT�WND��̌iB�I�t�f���E�8b�6HS�1 &�B��',���n��![Z��u�ԇsJB�I3<�����2Zi@�� >EXC�ɘK���[T�(H�ք�0'D���B䉎{�D�3��W�����?J�B�Iy%r� 1�H )ش�p5��B�)� P�{�c�He�<�k�Y`���"O�]�͐!���K�>C���W"O\!�3��&b��2�-��"O��"&#�&��c�/| �� "O��(H�me�$H$�Ȕvo�!�"O��5��?]�乃��+b��y#"O,���۝�t|K¡uH.�J�"O��U��<
ݮ�q�ڰ�(B�<�s+@�K����2��7KX|X��]A�<a0�M��N�Fe�HPW��e�<A�!�]|�8C[�,�pU�Wa�<�W�\:BKŻ�k�D�� ��c�<)E�E4d�����:��A�fI�w�<i�?�(]��-�9j-V)ȁ	�q�<�%O�,t�<�cO�̡dhOj�<�W�Q+M*>4[cJ�#�v�v�A_�<AG\����y1�pb���$X�<�m��AY.��*
}~�� "��k�<��'Ξ+%"YKь�<E�v��s�<1��^�%��^�J�r��1ACl�<�A�� ��Sύ.k�ju��MGi�<� GV�/x0l:��_�?"�X��|�<�D�G%Q�6��#�+|���`��b�<q5��n����3�uRU�L_[�<!���;����E���%H����<AP)ЉM���"��V+^��JPp܇�J����ùA��)�숬X��B�'8�A�¤�U��i1��_H�;�'�6�Q��>>z����vP&U��'Sh�����;H�Ƶ+)_�t��'~�87�u}:����Ӌ �:J
�'��m�1��7Z ��c,݆ ��!��'��  ��   (   Ĵ���	��Z�:tID;U���dC}"�ײK*<ac�ʄ��iZ"v-�(xrğ	"�6��������ϱmwN����"(.�tc����}oZ��M���

<�����a���4!(0�����0Ài��'��E,�  n�	^�6x�S�(�am�/.�H4�H�,)��	#P�N�p���
S��p2��=5z��0�\=��I��D9s�%#(O�E�Ā�2���-O43�M]��ܨؠ��P�M�TN.7�T��դMJ�D�bf䒅��[�$K;T9f�rӪNo<,���;Z��リY�{���'v^y8c �� m�'Sp8v�K�F��)S�!�����m�[�(�S�A#a��d��n���Rf�|2$F�G۸��N>q�lB6+¶��s��]�h ��N��l�9�)1��� I����"�|�D�E���3��ү=��}J��N�?�<0lٕb*T�d�埈yt�ڔ|�P)�²<IQ͛�FI��r�x��@��	Rs��ط��L���	�?��K�tW+�O�M�6FR�{@^� �OB� ���H�y#~����Pf��Η}�\'���Z��P�� �Ӂ�?�z��%$z������hϚ<3U�N��$��.̐u�t�|�`W6�0!xL��KN��R���2âZ0U<p�ؤ�?qO��C��x?9 3O��p'�P���ԟ�֘��K�./`�����Q,ff�dCb����� tř�M
_�>;��(i����� ts���q.���,�>��' �Պ4��p��dJ p��-O�	އc"΄�@�T�u�	p���aJB"�a�����%���_9vA�C�C<��5d�(j�dyRk[�$�d8�CC!'�FI�֩��,Xu0A#>  2"�'�`����dd�	�_���p�m�46
š���(T�t�AZ��Q��B�	(!P"Y�4�&��T�(æ��"H 64��Ѐ���?VzhS��|R'^�20x y�┕?6�AaT�'mh�Qgf�-�.ݓ�"O	c��  �?��Wm�g�Q�p ��trY)�	�(u�>}��J;���!�,����鍠9vr\����)�Q�����O��$�>�B*H�{K��[���=kܬd��[ܓ��=�S���0��ԋ�A"zTȍ�倍L(<Q�A�)9���a�' ��$��˒��@�����ȒR�"(nޟ���P���S�UV��2��� ���!a\p��;o��L�Iҟ��P�Q�-�gJC�P   }  �  �"  �-  8  iB  �H  �N  KU  �[  �a  )h  ln  �t  �z  4�  u�  ��  �   `� u�	����Zv)C�'ll\�0Kz+��D:}"a�ئ�Q2�}����u��h�ӊ-$�iq�L	���2&�T�4m�5�=�c���*Tr�)�Ǻ�f����W.��z��\�WXVш��׮DD�)�"���g�0���Dk�ͣ�%�6=i��$z�΂�P*@�	�Oa��LG!*��Q�4i��R#�Q� "܈\0�b�������9t݌L
0bW��M�R���?���?��?��A6@\�y7E��]�8�df��?��bW�hc�|��?��	�����?邮�6�8�רd�tP۔��?�����'��՟4#w�k�������(����p%��
��Ԁ!�!w�"�hS!W��5�'��S��!Ey�G�:��[��W<��D�TL�2zt$��\��͓�䓎~�i��N�8u��'��|�!	�J�4	iEk�!O����Iݟ�IԟX��П���s��8�׈+mH�䎘�����Ԍ�՟8J�4L���`�.��'/*6���C� dlqDJ���S�`��
�A�k��;ů��~��s��D݃0zB��0�		5M����H?p	�.lݍ4	�8,v^$z�
��a��6��8	�p�S���.��|����WsӀ�o��?��'
ʍ��	K���#��],�c�͑R��Al0ADx�1�΁�xoܔ0bF_���A$-F�x��ߴfG�� bӈ) !�ǧAd���sKR��D�T���]ny��>r���m�4�Mk��i�>�HS`�7]��|2��r� �pB^ !�Q��$��oX*�*��+n���ڔ4d���b�`�oڥ�M�G����H#S�*p��p[7���L��Pҍ��Ex�� Ô�a�`�Q��iٺ��O�`h۴��:������'K�O�� �J�|�~����X�P����O��l������7�MK���?���~�j@X�.4!���P�6�?a��v��!��?����cE҂"r^���P,Iɛ�	/��L��M+�$�5睐l�F7��~�Q�p�T��+
������ !�xoZ"h
(ib&�.O�h�q�AM����4$�Dyb�	���wy�jS�A���Z6�فChu� �@�?����?�I>i��?1(O��d�.u���`�Dj�F]�ǁ��`���D�OЙZ�f�� �ԓO,�i����S�?ч.Ȳc[��@�����wd!o�B\���^�M����O���=}jT���P�(bp��h x���'����Q�i�5�K_�M��4mZj�'R��aȶ䉘�l�
�͛�O�lbBI'=5�(�4KL�"O֢}�d�3:X��M5�¬B�!�g~�F���?��i��#}:�O:����.-M�:��J�NJh
L>����?Q�����D��_�J�L�����u�'N�7-_ۦ�|2$ؠ{��)ǉJ�+�h��-ߨ�Ms��?��J�������?9���?!���yGCǀ����ۓP�lт K�$���O@����.LO�␺T��T1b��*r�<� �rG�%���Φ�H�0r b>c������3��	��M���Ycc��y2,O��(@�'��t�?�O�x[�
�=(���K�kY;�Ht��O��=E��eB�=`AH!��9]����%��I'�M3�i{ɧ�t�O��I?S�d0#��K~){�-�gH�)�#K���d�O&�d�<	/���*,Ҭ:�E�:���c�"a���S.��I\jE�M�O\����#)��g��h���㆞�f�Tx`��+Zȁ�N��"}�E�H;$�">)QEK2q:���eM�dB���5m�t|�	"�M��IN�C>J%�cK��������U,����?���0>�e��9C�m�#crPPU��LM�ɡ�M#·i��ɰeQ�e��4�?���QV���D�jg@ �D�J�}����?�#�H��?!���?�֠�9"&�G���)����W�l>"q�c�-�Db�g�	��aÓ8���@�����p�
߃+�P����V�HA����d�Dhͻ�A�K㴙����u#�qO>���Tޟ�J�4ܛ&�'��(q�gD�e��t�%��"u���SU�o.�?�H>�nܧ|���á���I�<��+՘p�f�����0�'<�7��S��̓3.�\Z�� ���l�؟��4=4��BȻ ܰ$�/OP��	ߦ����E.pXF��!7$%8億Yq�a�Iߟ����jn��Fa�)n�pUjT�Pq��L�$Ń>1��]��H�=;w���¥,?���߮I,���l��D@V�_�^�¤!0 $f$��'���X���zD	+�@�n�2��'��2��*ߛ�C0�):�S�c�v����.*�:U�w�?R�*�O^��)�D�O�d�<�U�Qj�$�����$'�v�0B�]�5-��|K���MS�]f���'��y��耤�rH �2��'@u�7��O��d�Oft���ɞ1���OP�d�O��bR|��r��N�xP���6y���%g�7{��mZ)ւ��'*�L�E �I�b9�l@��R]iX��bȌ�yY@��Å~�n�� H�+���U#(�S>�>�r�N�q&g�&}�e@��}�y�ߴ�ɚ!�:�D'��OF��OPl(6gB1�t���M�k�$���'�$+�S�'�Х7��W�81�"�䱔'6�6ئ	$����?�'���
��&�BX[���n�<Q�B(�6��OT���Oz���`>��c�'h^��I�:&E��MA�T�,0�@�ɧS�)*��Qx�4�cf�
+JTM!ٰZ��� u$�(}��`��aX�"BN��$oŔd&���� �.u0<s�2F
�!���I�QŦ@ȧ�����xܴ!���hEx�K��ް#DBG'Z��D��$��?AI>	���?���d����p$��Gp 	�e�$n����ZϦ��&�M�C�iX�ST�.$*�4�?y�'$^i[��7UZ���X/x���ryb�'�2<�� ��K��VQ9/R&^¾6m;� �< ��Q�pN��#��_%�Z�#��'��=JqL��M�֌`lQ!P<Ԑ�!j�K����TP�Z�
lb��ҁj���)��D_���erӨ��'�(A�#Hm8�H��Eߌ:�<	M>1��$5�/�e������Aj��_�X���'pV7��l�^9���#$	(-�U˘�}zPml�Ly��΅CD�6-�O"���|�D���?1Un�?WѦ����O�L��欆��?q��<0�wH��]�*��&��7O�B!I�_?Q�O��u�&ƛ~yN��ߴa�f��OT�&��y��M���|;R���"�f<��`gY��Z	�0Η:S�:&���ݟE���'�����œ�n�%˒M�ܵ1q"O��)��S�X�����>7�v��U�n}2�/�N�hMɓ� {���Cօo�v@�ĺitRS�P�i�?��	͟��IAy���\L���Y�v~R��d�>܉�戣�R7�Ͼ.�N6��\���9�	*{��(m� ����
��Mm���閑��K�L�+�����\̧��l�'��xZ�Q�8�0��C���y�vA�U�i��ʓxv���	�?����5b�R���38т�*�Ýv�J���?�+O��5�y~��=W
��`��j�%�9kq�-�'`�6��Ц��ɺ�M�+�X�ɯ|�gC��#��Q����V{�5Ha�׫7����
J��?)���?���+����O*��m>)[$�>y���tE�[���RN1�B��W$@]�IѶH����$`���%N+Q�����,ppf��v�9�	#6F� 1!��w0P8c�՚E|�p�D�$Q��PH [��e��PN�f|��c	l?p�D�Ʀ5����;�5�n��'�����7��h�� �ȓ(�H,c7$���t�Q�ʰ�|�'�X��4�?�-O(�" �����I�� �1Wvmf��最:P���k����	�b�9��쟄�	�W�?��HѠ��9]KZai��Ϟ ���J���+@�Ѷ+�&6�����D0t,���"9�*��! �<�Х!��]����B�	M��$� +��(OP��'��6���u�	-��9�a�K+$�$i��6xp�'�r��?��'�mX�H|���U$A��|3���&k�.g���⓻S��)���N�j�6m�<��gv*T#��?i(�4%��-�O��@��"=�>e��Ѣ[����f�O��䑲k�6K�"4�9�C�9����G�8l���`�h3MԲ..0�9E
�@��=�'����W�T)c�PEIFYS�E�Ζ���Y#H�^��'ӟU��釖�� �G�O��4ڧ�?)4OU�pڨ@��..br��TJ��y�gE�3�ڭ1��3&��Y������O27��O0eEzr��(��]��h�WA�M�%G[�^A�6��O����O��Ků\\���OB���O��ݖ��}�&dG�\p~��ʃ+od����<\b�`�V ��m����;�ӴZ�����O|�!CK 9#�Q�3�̼b�֍s� AEl��ǔ�U�ȃ&��8 f1�hp�e�P#�~���	��x�S�0�h�8��=����<�w+��p�@�L>� � �f�I-�m�R
ߝ[~��C	�'Q�q�Wf$O�t82����"��)�/O� Dz�OGrQ��� ��2��E�� s,���$I��@���ן��	͟t�	*�u�';B5��̒vL� -�0��`���R�\EA�P�]㜽ѣ�� )�*�)�~?У?�� A=/��C�'�2��BQ�	D�ؒQgtPL��-�|S��������9Qz�"4g��~J���AȸHy�	x��'�r�'�O#|�E@�H�`�@�Ƅ-{zT�����$5�ɭ	b�Y� ��;P�!p7��udz�OP�o����'1@��¾~Z�C��!���A�zZ���ӟ
�н����?)B ��?�������hH��>�m�L/�:i���[/$�����W3�����	�vڰ�'�M�g�YAad�"rA��qp��5|��L�d�!'�eR��E�'��u����?9�O��㕦̍D�\��!�6Hh���E�|��'mazbƍ(B����̫
w��Y�T���?���'v��( ɛ�p@D�C#��.�b!����Ɇ7��doZ՟���u��T�X� ��z� ���9����N�2Y��'��M8`��1�جS�ݰT���	�pk��?�`@hA	�5�7U'��%xe)?��H0	 J�z�P,`H�H���,T��p�b�5��i�9$8��p�'>Oq*�u��g3���}�����妭���	d>UI�N�`5���I�(bV��#D�����u'
 3E��-���	�o ����>� �Qy���W
şh�����k
̦5�I���*�zRb����	ҟ��I����O��J֎�PW��0D�2�L�z��5�댚B�Ƅ�B�2%���|�I>i1��]8�b�_���I�%Ӓ�a�G�T�� ��L���|b�4h�����X��j�����c3j��)��w~R ǚ�?���?	�ba�7¨���'X�m:A� �߳b!�d̠8 ��I���M+���*΂E��*����ʟĖ'8l%�O���O� ����Ŋc�\�	��IΟ�Yw	�'����Z)��
T&|���PS$]�n�J�h�D�
Ό�b��V%mH�,y�zX��	D	B� �	��*�=�| �j�]~`����X�}��x��DB���{��{�T�rU�	�V���p,�'��1ئ��~���@I�Or���O.��D����(C`��ホ�@M�P����yD�
\���fS�Z)@tq���%֛��'k�	�w���I� ��>_[�(�����`�^	�f�!76a��֟�EKTҟ8�	�|�D��Z���e�ʺb�Yʶ� p��TeB<T��p��U��!K�x:��<�U%B%Tc䰠s�ʅe��i2�Ů%l�I_����#�!=,��w�0�" ���!BN���c�I�^u��K��>t3�)�� ث B䉁Y���r��'X��!Q!T�,���D@����J}�v1B�I�����>��\|� �l������~��≔2���J8d�ؕ��`
�/:����Q��'>ڂ�W+X�Yr�
"R�]��;*[�ɢW>�#�7T<dI�`�ň@t�T-�x~�D��+j\<KG뒗J{���k���u�Ʌ,S�Ή����}z$���N��������D�ܦYڴ�?���$7n�&o3�9F'����� �����On�S��{�dߦVy5���mD�0 �A�'����}Ӣ�O y��$�fn�h	4]�z�x	��N����OP��<d��h2��O���O��D��KG̩��(W�_�`=xY�2�J�c����"oER�lO2]=&x �Z>����d
�n@Hc�Y�QX��O�:�5�qjH�E��&Ǝ�+�.�������D���bT�d�d�]5xz�1�Z��v}L��;��OB���O�l�c��iyH�맅�Dh�-��O��ĵ<������	�	'�tb�2HV-�^LP�jћ� d���O�I���˓)>T�f�f��IC��D7K;jy����+3�vh��?����?��'�?������O�0_U�(�SO'"�p�ҕR.0t������H?4w@Q1m�~@����D4&ndIPA��9_�P�-�=Xr�8eo[���1!:,����&.�`1&H��(Oj�Q��� "8@�V$�L� �!���e��!�Oʹ�W��.*`�bt��=�����"O�kc��}�tS$�E7�����|�Hz�ēO�xiW)�t�D�':-;E�>H.k���-By�Tqu�'A"�)PpB�''�)&q4!��%h�ptG^�)0� uJ�j4b��\�f��LP�&��HtLm�"�C�2I��G4-v������mp@ة$��7> �<9�Ń���O��q�'r��<°
�2�F񡰎b��!h�`%�$�O����� W&6�j���g�H��Feޱ` 1OJ�=�O�r��M�l\
p��#���I2���[��[�N�ן4���D�O�0����'�P�Ye�I�N�X�Y"B�A%��%�'�i��F�L�D}g�T�GEt�Paev$�S(!.X ���}�:�FB���<f"�ѵ�I)��M��02@H��r��i(�O�ܨ�c� h����BO�<B����O����'�O>IxK*)� G�����4H��5D����ѫ��Y��R[��<�`j3��8P�>գ��ӁqZ��p��+-v�����O*���O���A�t��%��O����O>�$l�IS��J�:%���=�R�-U� $�Gm�0���C�˫ ��b>�P'�1���<l��L���
b�L�3�J�I<lM�dN�+�2��C���8�x��6�i/��T��'R���sÙB��i�Ee�R�<���|2���?����y�C�����j�aC?%�>�TC��y2��}	�,"�Z�p��ɚ���d�G�����|bo˱Q(٩�n
A˂��f@�r܌ R�><�2�'#"�'A��]������|���j��Hi�⟰͸aQB.Ǎ�=�6�G�5rݪ�����a3K�.]̢�<Q7�90QPqn�<8�d٪�lH޼hÀ��&�J�I9����뇫8Wp�<�C��)2�@�Un�~B� �%ك~�8�	��MC���^�'7�����[0WZ�AU�nV:�A�'�~Q6�Za�4:�.�?9&���I>�$�is�V� A��"��	�O�9��T�oGȱK�!�%����G�Ol�J�#����O�S&X3rKq�V<	� A��[�&��������Ұɡ�n�%�r��]�����ɿ�bu�Ռ�B<��q˄
hln�;��$ڌ�'��?�q�ULN�Dߘ�#�剾3J��$Ԧ��,O^5C�癍t�P6��P瞴���|�'��ɱ F!HSnD�@Γ�k��c��9�")XauB<A�%\��2�����?�,O� ��	�O�d�O��'|L8��gK���U�ف8,�hS7NS%I�����?f�Fð�;W�	.Q�&�ia��d��M58�>�"��	�]�Z���(����8�t!�TǙ"B�E �<e�T�8��4��KS�H�t��;%j�q�AO�◑���PB�O$ioڼ�M;�����#�Μ�M����@/_y�ô�|��'K�'��T�T��f.� xD�x�t��p�>�Ӗ�d�\�O�p��_.ՠ�ɀK��XZ̊�lb���O��Ē�|����a�O��D�O����M8p�N� �jF� `��K�m8�,�'n��B4�ݞ\�ϸ'A��J'I�:���C��*@�pA�&�3E����Q�sӌ1+vN�5[�1�1O� \�pˋq�^�J��k?�P��u�R͕'�]���r͟�'��SanHV�0��Ğ�s���H�H*�)+:1���.�hp�/�<��iҜ6�!�4�*�)�<�#�Z�,���5�4k@��[���)6�T�?y��?i��l�.�O���`>e�$H��� ��ɨc��01��R4��,��쇻j�Z$�Չ��s��I0P̂�;�Q���P�ʼ"����zB��8���B��#�, �� D#C3��Q,PlpZq�u��M(��_U��ۑjP�A�s���ȟ��If�'����d��[�,"t)��9L9	��#D���Vn�Ҏ���)��O�n���`7��ZȦ���zy���S�B�'�?i�b] 8��л o�'d�;�	Ѐ�?��}�.H����?��O�> �$-��[aZ�揝�O���L��.�� �N�aF�]�CI�!	ο�(O@@�r�Ԃ%!�Qw'�6m_�Z�j�x�D[�	�P� ��.:�(�Fj��@*��?�"H���h��A~R���(�� �3N���ː�ϖ���0>�a1�r�,$HÌ���.w��� ��U�z��K��{#iY_���	fyrG�(DU�7-�O��$�|
3Mɢ�?��� hb��t�>8��e���?��������(9f�BE��Ȍ�#�N����ɟX��%@/+�m@��	1��Rf�����V�*���h
5h���B6f��:)tuA%�C�t�U)P��@�@Z�$�I����d�0��s�RE��2�bc�@�b���T�a����"O`,�Ȋ:x�Qj�Q�d��&�ɜ�h�D�!�a��\o�1��S�m)@��Kl�<��O��D[*A*=!���OT�$�O��$v��9�PH2yBE�ȈJ>0�2�D�S��<��b�=n=�$��g3$}�b>����L���\;�-�2�C�"�"��!��QX 5S2�ԯ��t�j(��hw�3`0`�'(����o�r�8upw픿/�[��i���h������?����;+H��E�H�|5�X(�7� 
�'%��5OC�e�6P[�(F� 8��.O�$��|R����!��m`��]�м��bAv�	�6���j�"���O^���O�i�;�?�����T�׫V�ʵs7-��?���A�R_yp��ܨ@���S�k�!W|0ؐ�C�]�5GyB�\�r���Zp��>uܐ}Z�Ө_�Hٸ���;2�
���ԯ\��YK�OٕQ�& FyB��0Vd��C��V�"�֣_�c
����#l�Bf��<�p4ڂ���ZK��x2��'�y2`Ȃv�:iz��6�����+���� ���|璶x�ꧨ?�6)	-v�h�@ə�y� yzE�Π�?���������?�O���	)�F�`i��M��(�z4cWK�+3�I���P$>��p���	ژ�r�eO�'�UYP�^�	¼`�1LH0�pXs�۱�|��2��c/��Dΐ.o`k�,�e�'ͤ]���'<���<����Sޢ��"*ͨ[�n<���Qi��k����@S�L� I�''�zpjx*��/�O1���E��@Q� �&�~%@�M�f'��ġ<���Q�6�'2S>�
&JEڟXP�D�w�%�u�O��ά��F^����ɦw4��h��:�ق�E�ᦥ�w]?��O�<�Gnޙ\7d͘��8	ۮ��O�h�2��Cwt����\��6�ֺ;�Bc�	ӍT��H'��S/|Ѻ#��T���*e���D����N|:��z�O�l#'��y�xDB@g��ɒJ>���0=a�K
b��r���<O����Q�'G�i�>������"?��]�gԝ��AZ�^,O;���'K��'�L�;�I�6Cr��'k��'����\W ��̐-p��A���~M`1j��L�L����� -4(	�&�i ��\#H��Xi�ϛ�_�^�0&	�0|�"6� �&�bA[v	B8J@2�/�$>J\ZZ�\P�t8;r�ϱ4B���hv��O��$�OR�p�G��X5��iE.vx�����k�<��C��bX�h�O�*��	��jyM:��|R����1����M����a��n�w�F��5�������O�d�O�����?����4*Z�Z��4mأ��- A�h�������m���
:+�|�B���."��Ã� �ШB�!D �|�@Aǚy�`
Q�@7S?��B��L�'l�}�S�T&�1�C�ʔ_=t]9�Ǎ)�?��?��R�_)����	hVP�����y76B�n�� "��9 �"t�e D�9p0�O܉mZȟ�'}:�n�~��5ͼ��ٰ���"b+�b��Y���?9�%S.�?�����4�U,41�e2-�
?r�"�m#ܥy����}*��с,Z
\����I
L(�e���x}֬xN�I��i�h��,a5�i*|r�	�O�'ߤz���?��O�9��D
D��M�f��cTiQ4�|B�'daz��7U��ɠ��|����BI���?�!�'"��!m̈́#��U#��W�X��������$�\jUn�ǟ��	\�T��>�bB�rR���)�6[���RR��7n"�'�4�"v�45kv�C�̦bbp9@��~"ȟ�x �LU'e#��ґK� �X�ğ��چĚ "���lR8d8{�K�`�'/�p�j]�)����Ud9�$H�'T Q���?ь���O6� �H ��c���BBكd��i��"O�I6b�+2��0�!JI��A���	7�h��AIG�ӠG�	p@�o|$�Q֍x�|���O8��W����A��O ���OX�${޵���A'�dP�ƅ���Y��*[HPԘ8���.\�P�̔�{��c>%�l��e
��𓍀���I�Dޣ2����]��$2�WS)�c>�'���#�I�s��Q4J�rC�Q��l�pC���5�3�	7��)����4
��a4�]��.C䉭bv����hS��^��0�* ��2����K�ɾH����Q.Ni�d#�߾nr0�g�s���	��	ן��_w��'��)�VI�0���>B��cjG��\�rF˸��y*���p=����:�|A��.�?�BA��L̕۔�!��h��I*#�8\OF(�^e�\�(�a�ޥ���	<f�=�	0�M��i��O����C�+
�p�� �"��|{aBO��\�?I�[>,�2	ɦ��]'TY�d�_G���M����dB�lS^mZw��4��Hr�A�$�L�%F��0<���KK�'�*����"�+��|��-2Ó#�^�ExR��*Ɉ�x�iܸop<u�A5�0<q��ҟ��<���:D�&ā2�3�v����h�<A�E���rIQ;�6!�F	<��?�v�'}����߯a��qY#U)d���K>��-�?q$H�p~�V>�ݤM�t�v&U�;W����KR/���Iߟ�:��D_�dIs�� !*L��S�O�Z����&���C��X�rM��O�-j�a�/�8e���T)l�}��J<:�A���lD��r@�JF~�*�?����h�4�ɓL��-����L$r�kdmST0�B�	,iZ�y ��I�q�Z��"$\R��?�퓢1��lp�
�vيf@�_p�����j�D@���r���?).O� ��� \�X��ۨř�-� �F�`SF�88󪗇>�<b>c�@��Uj~�2\	��6���,f�m16 
���y��^�b>c������=$5r���c_�=�ш���O��Ox&�����pE{�ԣ3��i�Ǎ ��9���8�!�V0&!��F�=�&)���&Q~剓�HO�Syy�`P�v\.�T@�H ���0A�7+b� a�џx���s��6M�"!��U�r��Ʀ��cH��M��;SJN`(��̝Q�
�*߃V�6�;��X�����?i��+���r�py���b��꤇��I0��E,9�m2�@V-f��|�TG��^��<)��f���4S�.��G��-0��b�O��	r�`�il.Qb'bT�~N��<�פJ�����J̧�ʌB �H!���뎡d��'a~��\<���Zg��VQ�c������.�S�T(�<�C�L�4�hmVJ�`��2�BSy���7��O���|�Ŋ	��?a��&d4*�j�khe�01�n���J�(Y9C �g�I:0M��nH���W��=�����/κP�ʵ���9:At5����y�IQ�}p��pBӇH�z`�7	�'d��3g�": ��:xЇ@�1zFu����� ���9O�c��'r����:�S���X���~��� vlP� �FŅ�&�`�E��6]f��H�/u3�E{�i6�l�$��&nƧx\������/�ҭ"���?!�h�(mY��)�?����?��'���OrTƚ�y�=�AJ��g^��Rʺ}f����^�����<�j�OS�m��(}r"�jD�����Q ��\�q� M�ብ���Te���K)�DH+ʟv�ː��R�1�'U�))��������٠)��ա�O8\�e�'+��	�<)*<�5u�ݻ=%\��#��~!�Dޖy<�$��J�Rق���TV2,5��|r����ߕu�X x�HD�Uo�V{Z�PAbC� �d�d�O����O~ ���?���d�+/B�j�Jl��1C�OΊZ�*%�ũ��d(�����6�&|�fl_2e�ĸEyR��/����&Lc��T�d�UX�AE�)Ũ�UO�8|8`)�Cn](�@J'����v�dۀ~S�h�U�ć\8Px	�)[�" ��&���O���͢x����+��*�.���"O�Hd�K|������^�vq]���4�?�,O�pWH
��'��)DAT ��ĥ^���؅�L�?q��L�?����?���I�#4ѧ��b�P=H��e8���!P�����m@�R�v@+&�P�Ty�MDy�"�5��.�FL���
�K�ܱ����;\�\x2O:H~d��E��TD�HR�C�'��Odp���',�6͙W�I�,��G�:���$]R�)
)O����E s ����BO>:",#L�<(��}�<�%c�4d��+L f��*�Iy�n -1 6-�O��d�|j�G 7�?��F����#�4��E
Q�N�Hd"����)j��U�'#��"��ߑ4�2 )��^��X���T�����Á�?�,yӲ���y�ʅ
s�`�p��8(J�8�^|HPg��?��O$,��ed�3��#̯&�qP�'A@�1�� �V��<%?y�π ��a��C�Q�i����(\�"Opp�͊2^.4�P�@'�.��퉥�ȟ�MN�S*�1X�P�l�O���Od@�5���7ņ��O��D�O�I�O�� �;:�c��\��Т��	^.�U�𤏳f����1˅4*.v�U�X=�b�;}2�@��i:�D[�~��=��$��"_҄�"�ܻ{���h\�+R��ɟ<�jF����I���M&H_Z�[�h��V��<�'|a����N?�O8扳a�|��,�zx�;�߼%HB�I�>�����]�����!�#B�J���u�����'9�	�Jqa6�R�r�"5�+y���F�F�4��	��	���j^wd��'b�ɜw�Du���@�2�\T�BdP9��$ɢMMĴ�LH�=��8pF
Z;@����΢@$0JǙ}��ҰL�:n�)�EK/[���5iW6�N J�F�R/fHÎ�F4l���_9p�S5ER)E���g��7-W�'��h�b��yӺqS�"4\%�s`&D�`y򮝧z@Z�S�`D�o@>e��(�<���i"�\�x�����M#��?��O��m�"�
1�<T8���}���	��Z|&�p��?���v���e���<ty�+�	z��3����O�{��ѾN�}��~�'O$���ER�`yi��ݪv�T��JȮ 0���[i�D+�h����O�U9��'�BC$�i��l��5#@��,���B`�C�t��$�Ov�@��ğT��Ey���G|؋ʋ�G�8	&!�8��}�Nn�Hl|��Q�>0�6}h��Pr,��'�"�']�_���	ϟ4�	�<Yp��80	��
S�@�ɻ�	�i}�9O���<�GR��>M�)�� 	��ջ@T�b�F/�I��U&��c֚��-%B�����>Q2]bP���y�,7��O�'�j�p4O�O�$����$l�H�D�(���)E��-�zl�C�2T�
PnZğ��c�̟��NR0���ם��T9��놭�0A��8bEG�/~���{�hN��?9��QtL�˟'��N�O ������d�\��%���h�ȤyB���%c�"hX\�$�OL����O�,�I�b�s���V�y"O�]E0��Fג5w�M�������?q��YI�YC�Z?�Iڟ�����*"��/�I�ǟ#-j�93�O��?��[��$�I�3+M�ɑ�?�"�_\n�N�v�b��#j ����DU5&T&�����MST�'Ԍ�j��?��	F���$�d�OL�)P�U"�.u�����;\�^�"(f�D��,�b�'d�������v���'�M[�j��'�*����
<T%�Q��k�u�H
���yr�%�?y�'�0%�O���'T9�Q�73P  2g �f3"1G"~Ӵ(�V�j�x�,F�!ݴ�����I����lU�a�Li�-��%�02�P�V��f�T�f8�7�	��tm�:�Bߴ���^?���0R��H"�䇯O_�m�fʃ�%��Q�
�'ƕ����}#H�s�@�r�L4��4�?����?y��?����?���?i��{ ��:.�dk�-X5�p�]���I�I�ė'82�'�B�'#�=�'9�桺d̓��,\�){���:���OH��9���?���d��8ټ@Ɫ�/c�|@�GzӜ�D�O��O�H�O��SF��##�d`�M��@��eF�/���П\�'Nў���]���ra*� ,wt\�e>@���%�d�	�P��ӟ,�	My"՟N�r�B�*�^�)��[>�l9�U������H�'��T>���na��ϙ).L��.�/zq��"O@ȡP+�:��lA捖<`�l!�"O2�P��Jz��SઊOLTA��"O��(ɔ[���@�R�f4|P�"O�5(��۬Gۀ]�p�٬v*d��"OJ-��#V�~,\�s�
@���v��D�Zpc���2�򔁂��:n��V	ư'J�H��H�j��e�nŘ #�L��,!pI��'���?�f$���è���;�!�T�E�AIO�
_@t�'36p��c�H�܀c���p�*���}�2(r��@�Kt8�
��+V\�y@�D
 ��`ڔo_�1)�,��$+'^-�a��[�޵�Sc�5G\d�s0���?��3V	�V��.	�]���5g�H��3�K�"��`��E ŮAdϒ�!�T�1�Q�4ȩq+s�a?_>��vMN��l�=r5���X!��*`?/Vuz�@����5�IP�OD<Eq�J�	B������&�H�R�'����qİ��A�I�z�@\ �'c�RF�/i�j1i�k݈�"�'Q���[�P�t�P��c�} �'�v����Ϊ]�ʡ�֪F�`c����'x<ЗaC���t�f,�=d�Q�'\R���j��AV�����I:5��'�"P����b���ؤN��0L��'��4,�vJR ��āX�H|��'�v�+�ގ�e���J�<��
�'P�����gW��`P�[	)��'Z���D��`3h��]���� v�Z`�HD:��B��@���ir"O�����՚�TRԛ�~�"O�<8W럿�\5��ܥ����"O�L� ��{�d�h$��<f�Z�"O����*�7s�Z�1��A�S�U�P"O^Xm�RT�]��c	.�b��"O��3q�ںp96����%p�X/�yr,�1iX��U�	hƈ����y�!W�nr�E��.����)��y��ƇH�b5bu�Ϡ}��mn'�y�,�H��؈�ʍ7ogV,  KN��y"�(�6ĩ���~�0 )lN=�y���::ػ�ɓ�H�(7�yBl�lư�*P��6C����FeW��y��0d�h��Ǐ=_4��>�y���s���9�����x ���y"�sl|@YP���0E��N���yRDѭqΪ��E�'	Uj'/�4�y��12�8�!�Ŕ �@S�(�9�yB��;)���@��}�!��P�y2�]2���1���,Nd�!��9�y��ܫ
V�AY��}jiщ��y��Qs�TH��Qr�.��`��-�yrKBy�|��� <����H��y�,���ve��.D�6�.l��#Z�y�.�f���j� �-p���w���y2$ս9��`0��,�t�A�G�y�L�Z��9g��	)���G�Y��y��..�n�� ��%�0�v���y���P���7De*"p�EM��y���'��eK����'ŗ�?�vC�	�m��2�M�iR�SᔥN�jC��'>��ЅJַ/�*��
D�.C�	�^H�ب�Yq��R�g��`�C�	��f��� �_� R�C䉵'TU�LУ����`_�{�C�8 ��u��d�d$��j�_�UݜC�I�x�V`� �O��l��@�"bC�I<xQ�$)��X)T���. 1B䉬wrx �v���~( `Vi�C䉿>�i0�%�?]�)�P�ȉC�NB��?q��ӡ���&Bzq��B;4�$B䉧�2��N�L�x�`dK �J�B䉾_���ʣσ2�0��d��$~��C��@pL�2a���&n���C�$E�����"�r���߾C�I�8a���ID�0E��ec�B����Y�Aį����CL��B䉔/�rh�F��?��M�EgCOh�B���`�!ʆ<M�ђ2gL,��B�I)oN*)*-�*,I�x�
FxW�B�	+G��+v�Q�z:��KC(p��B䉭-
`���z��-(��]Z��B�I�LB����Ȝ}�R��'�8C䉻{�zF�4hyy�H0GGtB��ZJR�qd��������8B�	�G3�����ܔ3���y#F�:5��C䉟S�T�`EȒ�6P�т"�٥%|�C�4eK�1��Ȍ$� ��Ve�g��C�I:c��K��W���8��C�IY���L\�Fݤ��ٌNԺC�IfR�C�%�)Z�]��a�>�lC�Ɉ_���#ਏ�uh�sa�O��NC�I�����D':H���w�P�j�tC�)� �����iQ��3� >��d�C"O��A�R:����!f^o�\�z�"O�,a0K,l\�e)�Č/�:h�G"O&�*�Kߘ.R(< ���yf���"O�bD!�=�P ��T�zZ&��@"OF�p��H��k�nڿYD�ؕ"O@��R��+c�Yj� �)%�a�"O<E�!�S�bV
�2C�D 9�:�"Oj-#s��)��\�1n�G��1�"O�D ����%����	�`�"O���BL$�x�Gk[6\��p"b"O��xcU��=ģw_@y��"O:ycI�#�"���!��rrm �"Oh���B�0-ڌ���!��Zu��"O�Y�G�H�pOLM�5 ¹)�*��"OX�3p��R���⇚.�lI� "O�만����2�J�pE޵�"OR��5�2#�]�1�@�0=���"O��6�	�eT����HQ=@H4��G"OBd�܉Mi�-�B5<f0�s�"OVa�C�ZdJ�9��=G����"O ���kG1n㖥��< dp�"OVD:U�ݥR��a7Zr8b"O��8����P�>L+��?/ts�"O�:f��+.j:}��Ň-Kf|��"O��q�ɗ]�d��嗰NԍQ�"OV�OԩF����Q�Z^�NHK�"O�Y��ʹ *!2cٸ{��T��"Op���8V��#Cto"త"OԔ�d�Y�`�R��&���Lyi"O�̛�`�>N�((���^c�u�F"O��3.׵Q�L�t+EK���E"O�T�%)O�P:m��%R��5��"OJ\��K�T�@D�f*�)<�JAˢ"O#��]1����F���D�@�"O�87zYfXP�Ӧ��+"O�"0���4� �Z��бf"O"t"��B�J��g)}��8�"O����ꃬ_ �{$Ièi�B0)�"O� ��~`�5hU:�1R"O*�@��c�M�4Hޕ\���"O��;��P�2
����Õ�z�ȓU�2=zf�.+�$�fG	V�ȅȓ7�*�!�\-d�h �n҇G����l���UgX^���S4K
�XC�h�ȓ^ (���,�*{̝SQ&A>E}�`�ȓ'T���5JT�l�Ȁ�L�{t�	�ȓs��4�Ђ�6�)��m}�� ��Z�p��P'aӔ-P��W�J\�ȓ#��	�@�L?����b[�=i�ȓ���"���K����l/z��be؈b�.[�?h�d,C$x����ȓ`^L�kͫYzH���Ӣ^������P�Ι�5QLŲ��"��|��#�� Q�D"l�hD��8�&t��Tt��	5&������w ��$3��ȓ?.!��:�TQ4���)4`�ȓ,xf� ��=X�
�	!� 9S4蔆ȓk|l��@M�w���R������3D��Q�ϒtv8W��.�v�f=D���j��`��i�&oE�`z�`��(D��J`��-0E���>i�b��
*D���0X�B�K4J��?�Z IA$D�(s$%�Nt4|�  KmU�`�#D�� Xp�ؒ|����ℐ�D���"O��:�+U���
��]$1=� "O������v���p3�9�(�yt"O\ j�G^6;� m��b�
�~%�5"O(�b�j�)W�)	�A�t*u��"Of9�OC
W�hE�5ʐ-�B8`"O�T�%9d��t���K� �zl�"O��p��ԏ!�L�q�넁b��U"OUYEU$M�5��kC�e�$�`�"OJ� �&���	@d��W��R "O��62gA`W�]8F�����"O~�q&�I.�Z�����0w�hx�"Oށ�׊�b��tj�l΄u�f�qw"O�衋�$-s��X���[xfeSe"O�<+�+��CЦ<b�+αM�T�V"O8�����N�K�I�(%���X�"O@�ӱ�e��#�(���B"O��������赯Qyv���"O��qEŹx�@d�A���ĸ;w"O�)I5�E�
 jF�7�lР�"O��`�f��?�� �a�r�"O��� ���qKX�`��^�0l����"O�dR%����G�L�:�2H�"O��r�`C.}.P�B�h��;�"O�a �b0w��d�%���RFj���"O�( /P�M�P�� _�!4���"O���9!&�)7���3D���"O�\�t��;z�԰Z��+�\�Q�"O �!aV�C�$9���#6���"O��B���
�c�#	*�x�:C"O���3��
(�h2C[�(�����"O92`h�4 6ja1�!��IJr�ؑ"O.�:�@C>o���G���YL���"O�,Z��%% ����=#��6"O�0 4㊃\H�Z�KH�u�n��F"O �!N�~p��c���;��x)�"OT�YcJ��G^
}�t��)d�^e��"OL�4c9~x(c��Ě"�!��"O-C�I��2.��	��)p (�"Oj�j�ω+'� ț��ʳHLn��"O�D��m�,H�\�z��+՞�G"O"�3¡U�b��Pթʨ�p���"O�z�'C�����o�(2���"O&
G/� ut4z�
�o���v"O�	�q��j��:�lJ~{�P�S"O�`��3!����!����%""O|d���PU�F��2*\�z�"O��;5I� t+>�ڤn��i���(�"O`�!�)E��*��/@�>x(�"O��P�F�\R�"ד/��p��"O�Q�	�W��K֠O:��@!�"O��ȓLE����>/�LZ���:�!�8���qB[�^�E����5!�L)U�a$&��'C2��ǅz"!�$��M��*E�׿N��Iu�Մ!�ĕ I(�b� ��Y	Z\(���i!��X�#� �+��i oא&qO� ��o@�%�h��b�QG�\�Ś|BF�-��,�2���%c���Ѩ�y��� �,��BQ�V�pd���y�a��m%1�&��Np (����yRk
z�$p�+�Net�Q���*�y2K^/
�� Q��F�62�-�ř��y���$n�D���!�Z��I#b[��y��'}����ѣ)~�d��,K��y
�  p)��IFl\bք��L4jZ�"O�}�����h�ˇ�:��Ȃ�"OZe�p�IbPz(Z����0"Oj���aU<e��e�߈M�"�h�"O����"�8���g�!i��!B�"O��a2FʮLel��E��8}��:q"O��!��n��u�1fR6u�Ѐ:"O�}rT��5�&$K5�Ll�М�"O������,!࠹������T���"Op��M��9I���j�=� !u"O$ȃ�/�;"�v�[��D'J̛3"O������n��r/׺F���"O6��`M�':��ȹ���,@�tls3"O�p(�.�4( T�9d�Y4"O�ukt� ���Aļoaz)��"O�xB  �Tj�ŕ�5R��"O.(��$�_<��eA�{���s�"Ordؖ╴��Pd���4�E"OBA�C�S �"챲a�?�
h"OTl	�fʞHQ��f�0a���)�"O�!�3Ȟ<p��y��ٯP�B�bc"O�d�G��#c�<��*^*p�,� �"O>=��eP+3d�%A��O�TD�%�d"O��+A�ɦO�p$���
9#0@�"O��y0CZ7t���#� t�(H�"O4����"/<$�W�Ai���`d"O�и��֟ka`�86(�:5+���"O*Y"���21�qZ�/��h�Y�"OP��gNx�0L4�s�"Oh����	C����PC��<A�p)�"O����޾sZ��gH�T%�f"O�%ZEF��`�d�N�~L��"O,��W�?���1��8od��E"OL��E�Ļu�D�0daR3gL��"O�,��@�&q�0�'�pR 0PW"O���4���re�]B���T*O�yb�8�y�J[U�8���'\9���J�w�y�E�;#*|��'�y��-ҿPT�C�A�G1��h�'�n�sfJ�1�b�uiz���@�'��HӁ�uk�ސq@�m�`�*�'�d����l儉��M39���R�'J��A����Y��c�k�1dôԡ�'P����L�d)�d�j����'���J���>��� ��@HtEX�'J��ߊ8ؒ��!*T�	�'�Zɂ"�7`�U)���Tj
 ;�'�^}b��|�VJ��F�=�V�p�'t���$Z�=�`���C ��ȓn�6 ��4S�� �e�Ē|�A�ȓ*'�<yӧM��4՚NP)5��8��[�@���nw���"��%nh ��+�d���\�S�(��Bf�*1	�مȓs��� �ި[x&U�4��pZ�]�ȓxAƉ���M{�D�B�"YT<�ȓ
�Z�;7�0��i�7��4TX̆�`�d` �֧7N�=B	P	;"j\�ȓu�
�@�!6�,5J�lm�H��ȓJԁAbCƫ4!Z�c�L�-\����j$xBNe��a��N�-1��ȓ}�6��2e��m����	U�l�|A��
@6=�4_�U��x�e������D�4A��	QZ��5@@�_�m�ȓ��H���)i`��QmD:`̍��S�? ���Pq+�� �J��F��ɳW"O���D�<Zѐ@�Ek�@S �I�"OT-�`cMtI��p�V:D)���"OT�$(�7X� �a�n�H�`"O(���,ީ6����"�Z!�b1�"O�X��"F��T�Ql���+S"OX��iF�&Dsb�#|Ğ��D"O���q�>q��X��f 	MƦ�� "O�9�6cܫZJ~���dY9�ʐ"O���f@\�`L�x��Aܙ!�"OV�� oT�gy�	�����Z�R"O��pR�^6oD�9w���&�j�"Od�	;�BI��N	+o�4��"O~�0 �lX*�Q5(�`�2(w"OjԨP%QN�*=�ӯͻD>$YBA"O���Dhڐ*;Z�q��ǟ9)<�p"O�!q�g�1m`�uY�G #T�@r�"O@`áLD�!�8��D��7x0�6"O*�1S���ػ��̂*jP��1"O�a��e]��Ұ��*�&K�ds"O�%�,�x�&<��J�#����"OF�������74�Nl�6����!�DG��d!4@����aG
�*�!��D��)��3�$������!�R�=�	J׭Q��� D�زy�!��	r����?$ʹ�+���9d�!�DK�e�v���R=C�f��eH"�!��Y��l�`� �'2�����V�!�(~rtU��'T,%+�GH�H?!�dO�[�ܬ�sdV�wt$xq&��<!��A�a��� ��[r��� �#�!��R#��X�R1AUf%R���,�!�$Ԩy(p���8Bc5@E/M��!�ɂ-�X�zCm��~����F��!�$N�r��������ӥT�B�!�D��pe�a�s#!4�� �-ɋb!��I�?%�������LQ��*F�62x!���Gs��ca���> Z�%d�[!�B��@̞#Y{L��ԋ>�!�D�Fn��чk�iIHp�!�Ě�v��Q�k�8.�0�0i��Kj!�DM)����+:ڮAB�.� E!��E2(H���C3��"�
�
]�!�!W1l�R�C AJy���)@�!��Šjà���g܁^�fI�Q/,�!�K }�%�4��^6j�q@i��!��#���ȵaF�'N �+!���_!��Z=9�{���If�E�s�!���s��Yi����j��-	4!��>w�LA�A��Urw�\�!�$�2t*�� ��B�Z��&lՒ\�!�D�9(Dh"�!�%Q��c腾"0!�*8����Co��r��`m�2)!��AiJj�(�a=���%i!�T�<����3�s��J�_b!��yQ����F�P��mjҺ5W!�D������-��yq�]!��F����1���#�� �&�2!�Ď>}S�01E�ݟ �H*�厎B-!�$���<��XS�~�#�A/'!��4x��i�%Vj
QP�傧9!�$@�2�2�0��^�y��,B�K�4am!��,�y�Qnہ@�R
ClV!���uOҙXPLM�;zL<��	^4`�!�� �P:�\�T��#v䅤S�49S"OX�K��!^Ӿi�2dЍY����"O\L�gA�^�Ĥ���J�Ū"O8�z�E��y�ǥlU�5"O\����R��Q;�R�T.zL��"O\���I���ɡ��2=�bYK�"O$�Ғ/�0d#�ɂɜINXp�"O:Y�F@[�-'����%W�]��@3%"O,�h�MH!U
	
�%U�4�*m�Q"ORQ���	D�ѳ��1K�<Af"O̐��B�$GV��D_��a5"O��"cZ}I�yH#
�����"O�5��A��AJm�3	�����"O��A� �Rߖ8s���l�:I1D"O��T���b_Ҹ8elO�[��I8�"O����K�-H���RF���
$B"O��3���uܔ��Wi�e��i�&"OZ���'"x��NG;���KA"O�$a���P�x;Q˗ 1]
�"O6�s�)R;]�` �F�U�	�"O���mR�4Ѩ]`��!e>��"O "��E�X0ܘ�k�1����"Oʜ!G��tU�X+�X�p���"O&��V��u��r��qǆ��"Od<
�(5n�y��!Z.��*�*Oe����pE�A��1�'�B�"�?w��A�aBA~.D��'�q`���0!jӜ/�,|!�'�������:`��50rV��<���'��3��=!���۝��c�'} ��˽\e(8bDC6hB�'P8=��L	�]���Q+��8�'W��Xq� �I#.��W�4�i	�'��5�b�Îu���ٷ
�;D�� 
�'�,���ˇ/}�]��֒IDl���'��K1c˄��u&��R�|��
�'�,���oXߚo�Ju�La
�'��)��Rr�h�q0pD�=�
�'�`�3�\̘�q�g��}�V��'6��'�ݠ"`�e���T}T@�
�'>2�ժ��V����UnMm(9��'m�y��Y�y���bTG #{P���'M����^�&�"�%��'��I`�*��`+m�A�  �\<�	�'�b�
�$'}<�f��S���s	�'אY٧�>dG����DW!M#t���'�,9��a�4S.��sQgO��,���'�vt���[hg�"�)�L����'R2��?�Dm��
��@Cn�A�';n�E� 3VN��)�L՝+XD��'	1�D�9"6�|Ks&�#^6��0	�'%L���q�bD�s���(���(�'ˈ�	v�{��d�I�]в���'�0�c��Ϸ�K
�L�HR���c�<ɤ�� ?�q �D˻CÈ�sl^}�<�3�Y�r|x�� �N�7�,�6��u�<�!7v_� QQ�?jʈ p
�[�<�D�^������f�JEɚU�<��H�]�R]B�ԣ$�RpRULO[�<)sK];D����I��S����G_�<qP��wx(�Áe��$3B4��%�dܓ9a�l�A��"�@��A%3T%$�p�7�Z�+sdQ�a�Ԇ�@�D�<D�|��)��ů]�\h����9D��``Iw`�	�c�=�x�"� 7D�� x0����\�B@8aϝ 4�N<��"O�MB�� C�x����̞[W�|aq"O�} ����!�9�Ԅ�>OD4q�"O���k��%�d�r䇖c�2�I"O"�
�ڹG;x�3�"B�8��SC"O� K���-�J0d!�>@��0�f"O��R�o-N�8�@ԘR�`��'"O>ix��`S^azS`�#}w���S"Oj��N��#X�첅�;#lx'"O���6D�
�d�����ZQ>�;W"O��)��@3'��	kw��%}T���"OB-;�0�P$����uvE�C�!��O�u��£�8�F�U�!�D��tPдȏ�_xSA� A^!��颀��˓W�L���$S!�6��j������1�K�qD!�$"�ıZw� ��A��E��!��ɿ�jİ�\'Z��TC��:d�!�$_�e>�����	��ux@
�!�ğ� f+r!���f-)�!�$L�������1D�Pc��9!�N`���qqƐb8�T覅U-+'!��G3")r\�,�
YL�.K�=!�d�W�~��t�H( ��,�P"Ƈ=!�d�C (t��'�=j=H�sb�� 2�!���;Utt�U�W8/=X�9�.K�!�ċ/
���"nɋ2����H�M|!���,LQ9��g�Uo!�$ �a�6ds�O��=H�L��+[� V!��
r>�Pq2	G�89�k��ѳk�!�D�y�x��$�=�-pv��-�!�U����XB��^�i!��J'��BqƜ -V\X�G�A�zc!��f�mЂ��$RP��y jH!�!�D�(y��ɉ��̰+P�HzC��`�!�$T@ä1���ZL�U�r,�2�!�]�Hθ�*'�>L�ail�<&�!�P�uڀ���8�p�;WA�!��$-F�#�I	(��Z�]*!�$��8dJb/ݹ�ұ+�L�#9!��C9j��AZ��,����J�
!�dE.J��2G�Q�V�����R!��ؔP�P��u���l��i��5<�!��M>qŮ�����5>.Z<��m��;�!�Ą�:Q�����s*��*V8�!��u�MXE�;�r���+B,S!�»"�HEb�$isĴ,^�Ψ��'���(���&��0���:���'d`��ʀ\��]�7מ�J$�'Z�y�gԈ2(�"�H#�3�'L6Xk��70��)���֣H!$ !�'&%CvNU�#$Lݒ5�\.o�UR�'�m�v�E�kM.I��C%-��'�n�qE�%(���t�*V�	�'N�NS5J�$����їWd�eI
�'qjE��- ,;�)QC+� LÞA0
�'�"t�4���%��=J�F�Sb��
�'o�x�"e�>q$$��i

-bi�	�'`�	3r�۲w��yg)�<>��	�'���
��$čj� �PHj�J
�'�#k٬D|p%8���.Ya	�'9��2B�(~:����Ǐ.����'��<�v,�6Q��� �:�D �
�'�F�@�C4*�FMi�#Z(,��8
��� |�B��+~F�"��L XL|� "OL�ҴD�+r�̽�çU]P�"On	����g&���坳m?\5S�"O�Ik�j�Ni(��%ٍr"r1*"O�=Z��0.0���Q-mP��3"O���ļq��9б��'��A��"O�5`-G� 8���SMǯ�V�ږ"O�1#MG0mob�����nـ�"O,��Z�;`����p�0���	Z�O����Kزj���t�	�Q���;�'4����O��"@;���(:�
u�<Y"�(%��E�� J>`�Z�KVm�<����!Ŷ 3埄�X0p��s�<ɀ��Pl�s�����Phw�k�<���I�J.��SH6z#<����A�<���$�R�K��a��0C�əz�<�֍A:"�Z(��`]"Pz�axd��L�<A��� �����A!\�4�E+�`�<�@�n���$� j�6�3Ư�t�<�����cZb��A�@�C���۶ONw�<)��@�H��裢L�|�]	 Ju�<iR �?t����@/f�%��
u�<a�H���>�3A�W�~%� �Ms�<�2���|fLP����

S� �3NAn�<�dG��U�bV�[y=u
�H[l�<q�J�q%֥��&=�|���hAh�<�7&�֧!���*a�d�<qWJ)�B��QF]����q��c�<���ڈaw��a��2Q�L�P���\�<��o��fTȽC�h�}�II��Y�<Q�fN�>i� h5�N$�p�[r��<!'],Wt��%�AA�F�����S�<!�3N�PM��=�hUG�<QVH�9*$���-�K���v+�Y�<p�2��e	S�F�>�pAa�~�<�0�M��j��S���;����![x�<�qZ9��s3�ٺ?�4���Dv�<�AJ�S,��HQ�ċ-!X�cB�o�<���I��ų����e{dC��o�<	����g�Z��S�d�nI+E�d�<!���	N���B�/V�ȂF$�U�<Q�a�?B30��FX/hk�6�,�y�G�/jr5�"�7^�Y�'��y�b���0��4��/@qNh�p�B�y���J�!�0�Y67������2�y���VF���QɃ�1 �H��ѱ�yB�	gӨŉ�FM�w���6"���y�i_) #fm)cQ1Y) ��gL��yR�WX�40�׌�>U-�lѱ���y�OYf6�9v�˦�0�a�Rl!�䋋BG�Y�f��T:<!2���3;�!�$�,-��4X��W4(�P�S�"	�c�!��� F�T�V@��~�.-��޳CD!�D�/�8��F��e� y)� �g�!�Dԡ%�&�����$�$ĉw!� �9�������1{�d���k�!�d��E��p�����A\��7�G�iB!��i-�lh���('��x�g!��	22݂� ��.䠱%R�Q!�{�Na��hĐ_���dD�iO!��K'=)��4�^>`�(	S��/o�!�E0c��PHd�éU��0BW�b�!���ӧ!��+���+b���-0!�������oə:���K�E�u!�� �,��X#v��ź�Î{K���*OP�����xh0l��,.R�d��'�&���N�/S�U� 0z�i�'���r'�s6,@��48;�'�����Ĵ.�8Qs*�t�^���'@"���cI�z\X���.nB,X�'`����iO�����R�E�<O`T3�'|`5����[� 4�A���k�Tl��'&�q�ƨ�>��� �kV�f�����'��H2��Y,T��q0�\�4����'�݁e͜-l�(��M�\��2
�'e,��/�K�\�ѡn�k�L�
�'�����Iӟ �.� By����	�'C�\ �M�1R��yWfN�m1t%��'�D����	W2�:�Ą�V����'����4b�[���S�X�{)�5@	�'., 1��TMn�C5b�>��	�'�ԙ�/ɕ��C�H�\s����'�z��Q�R�Z���W�$��'�ջ�k�nZ2}萧
�S�(���'��8G�q6�K#�ӉID����'�6 ��.T�}���Rt�� ��'�����Q1L�����K�"�0`��'��ِփT&oQ
lA`.�hT|;�'�u��ÞA5�,ڤ�[^z�l8�'o�j��ͦM��(�#N��'�V��-��[�(hc X#N��{
�'a~防00�8��{���
�'�,iaFZL�H�x����
kBw�<�q�A�� Ux��4@2'6P��-�%s�J4v�� 2d�.��]��*O�E:�
��_8��aׅVp�z̈́�r	x<HU��7dB��e���P�m�ȓV`�q��X>O�dY�
J!U�굇ȓ$��lh"�K��4Q� ܞ$�=��y}�����dE|����|p�ȓ4.T�{��.��Y�a�Дz��̅ȓ%�>\�0"�$P��_q�`�ȓF�T�(�#�>k������ ��	��������~(C���6�P���(��@e�*o�¼�i�2�t�ȓ%���B2lZ�2�(uz�N)��ȓ��!�uo>)*P.Ð�܄����j� )לؑ��\�&d���ȓA?�̻��ҁ}���q�m����Y��h����1�A0 R����K�OVE��i�dq9�]O$��"؟��A��Y�T�q�0�nݸ���֘U�ȓ���D��D�,��dσ�7 Z���8[�H
�I�-���O4O�"��ȓ
�1;4C�~PHYS�	Uq�ȼ������b�vL�L����up�ȓ�����.�LEn�c5�F�uܐ��	n���E���g��sP,�(n' ]�ȓ:R�]P��[�
�t$�ǎQ�`��\��&n����*ډ[G�:��Q=lL����B �����$xN�"��_�_�:C��2l�C��26@��ڲC�ɴM�n��X�,M�#��B�ɣ`bX�ZD�^���#��&�B�I�|��@@���V:�c"׫g>�B�I�-�Ԁ*䤖%x�r���Պt~B�I�*xT�T%E\�s�#Q�LH^B�	�EԮ�6jW�{D�S�ԧ$�C�)� ��!���9�PD�`B�"G���#"Ov�Ҡl�B�ѐ�әV@Ly�A"Oh�q�(M�e9#�����B"O*5�G���J1���o팑��^\�<���ݙ?<�9q�>u�j���A�<�C�5}��ibH�M��j2C~�<���	d��5����G/���㫎}�<a%bŒ_�
AH�,^�x�V�6"C�<12�9�6, �%݌Tl8XI�N�{�<���ZAT��e^k	���j�l�<qf/�y��(������j�<��:�Y�f��r�>ܠ4L�l�<㪂�������Iv����B��f�<iTȐ�	J����ޅu��0��c�<�G��r�θlc9\�@����Tv�<9�H��5���h�d5�\\h7RK�<	ЊV\-@�af�.�v	 �*�G�<9rꋤ}d���5?t���[o�<9efd��]��D�V�æ+\��yb�¶tzxU�Ž�0j���,�y��� &�H6g)uv �d���y,!�v�b��$u&($���y�%�4V�{+�ǒ� ���y�`�\����7p���!5��!�y"�L�nL9@� 2xª�tJ�
�yr��^m�Ň|�\sӌֵ�y��R)yi^ʕŻ��zb%�/�yr�4^�lu3���C���ȇ��yRjҵG�ɪ�/�-frY��J�y®��޵����c-H����5�yrbZal�q:�� )ZԒ���<�y��.l�ѵ��v<��A��y�FVv�80���0$✱fN	�y"gU&@���]�w"���\��y"M#4_�
 盎w8�J�@ɵ�ymH7+��U[�Hq�$4���Օ�yb � �E��Õ'jg�A`n9�y��ц8c� �4c�+u�DiaW�C	�y"ʗ5c<Q�ŭ�c��x�����y�O8Lm\�&��$`1ksC��yr��%BZE�P�� ��i�Mި�y�`�(xIB�ݲcȀ�p�`T��yb��y���"��:`벝J&��yBß�zݦ��PgR$X��S%���y�֨uD����n�6>���k�F��y2ʉ|+H�R�J�=S`̹vB���y�#�p�Q�����в/ى�yB��mi|a��"ڈg�^M�E���yr%�~�*���G�n��WN��y��/�1�UG�=*��Bp�U>�yBf��� [��/=�,�����yb��%l�MpUm��C��%X@]��y2_s�tY6e�K���Hܞ�yRMғ(~��!S�B"S�z�� ����y�hV�qf�!���F�ܨ���y��ͯR�@}� S��@ʶ�!�y�BX7���	f���Ll<��J��y�h���Z�DZG� \���N��yh�<G�^0h� �0�r�*G�B�y���j�`�#�l�� m26�I.�y�� �N����b��"�J���0�y2�Q)xZ�h'���Ȕc���y� &��e(5�^�uQ`��3"3�ybGo�B-����Z-c.��y
� ���ѣ��	����A�R���\iA"O�D�J�.��Ս��d��	��"O�<��e@5�|�uM^"a��q u"O.��7 �98���m�|�l�rD"O��dɄ<J�)
elC�R���"Or�[����s��I�LÇ
����A"O���<�޽�5&ƞ��"O�)
�F����Ũ��'�6��"OD���T	N�*�C��(��q"O�e���؆lVx�CR�Xi�"O��"L� uRH�I�jz�k�c=D��8�]~���;�F_�8r���!/D���¨ƅO�(����/hq����(D�<�ӬK�?Ԃ��]����*O�}�玘�'<j�J'B���� "On ��@R�z���O�n	`�"OD"́7�L�i@��0l����"O���Kԫ;�F,�$a�OF�A��"O��9�g^V�j�Z �,7PPkC"O��3E�NkXe#�叙#&�,�B"Od���� ���P�s"��%"O|��B�=,ތ�a�������"O�vHE9Au0�*�E�$�q�"O�	Q/�#H��a��g�(O��%��"O�%�"C�|G�	eS�j��uu"O���f���saD�z��:� 2"O��;���!
�pl��Z�<9B"O��� dsK
�	%��z�d]Z�"O�"�f0&�d�H�+җ	�R��f"O���c��H�1��
LNږQ�"O��+�)nQVs�h�1ٜ�r�"O��e�?m�K��-��U�v�U	�y�B '�l����X4{V�RC(J��y���'>`�,��iR�2޶�-���y�I�[���Hі&C)����ye�$oV�-�uj�%�6T�� 2�y��� d�p��n#>�z����y"lD/���B��;.˺��m̟�y2��B+XLsU��+s.��ł��y�k\�>o�%���ʾ�ԋ�@���yc
W��AA�A8�@T
`(>�y��D>d�(`0q�Ɩ�~�wj=�y2�W.�zl!���m*hВ�h��y2�ٍB��pҧA�6iz���#F��yC��4!��R�&L/�6�Ӑ��y"�ڨ'�n�ʒ+_>�Ɣ;�(�(�y'ÓJ ʌh����O� ��+�y�Kѳ&t@��q��>j0�D����yb�$
��|*�e��a�t�Pk���y��?�� �,T>	��9���y"$D�V�D�i5B�|HI�)�&�yB��ܬ��f
U1i���I'�Y��y�ij1R�I�nd!*0AQ�y��S70��%�Ԡ��h�(��$6�y�%B�Y[�$���'���$k��y舖8@z�@ M�r7�`A��a�<)��ݠ����,�G��y�Kt�< ��P_Ա� �S2r�v($�Cn�<��J%��`J��+h��[քIl�<��$��]*\�c�(\�'��8@h�B�<����� ���e�"aBaXf��U�<A���JYV Q�GH󰴑��QN�<i������i��ї/ ��RdFI�<�IO�j��r���UZz$J4JAH�<� P��T��tUc�3O��p�"O��(
PV*�#� ��[��`�"O���1/�"��$S4���0��s�"OB����e�v�b�-\s����"O�(3��QV�Ջ��>Kx�E�"O��A�ʔ-P ���"�U3�"Oּ�s�G�yֈ�bE]���b"O`ڱ��Xɠ��Q�Y����"O�5��K�	&z�A��ֵ$�8"O(	c��͸M1v��84�h�x"O$�st#G�``�Z���d{�"Ot����0wʎYbw��'=���"O���5@ۄi:*�6��9`�Ԋ�"O��s��%!x���Ѕ�E�4�f"O����([I��0I���"O��q�CŮ5~�"q톜`?r)��"O�������o���rEχ�����"O�P�KC�# ��*iR?�R(��"OHp��%z�� 	���5"O�IxD݈+f(x���c��飗"O�Ma�� Z�JE�0�ÃD�l@��"OFH�uٱju>$�F��F�$���"O4�*3�ڟ}Ex�:कT���)�"O�%��m�^����`C�8�H�p%"O$��e�~��)�#�� Eʑ"O�ˆ)���
�a���	K�r4�D"O*��E��;`%&hS0�*xU�"O4� �H�o�\邆'�5���"O��Cc��E-BG�s2��p"O =@2��+����-ьi��� "O��!�g��h"kJ>b�PB"O�l�w��_R�HS�*� j�l��c"O|�v*-i��ث��(M�����"O^\�<'p�:S� }t���"O�tj+��f���p���i�!(�"O����͙�%7����Iۏ��"O8�* ��w�<�)���6���"O<�Õ^��E���X-n���"Oڰ11g�-��ؑw��HVpA�"O�dY"�Dxgd ��R>U��ȪF"O��Z�ېCO��b4
\�����"O ŉ6�X�'H �R�� ��"O��@EĆ��,jAur2�"OV����K�zz}��l;Hs���!"O �B�Bȡ1��|��N��oU���"O���2 C�B.XR"KИ/�0 8�"O���doK�md�`���Ch��E"O$1bς&
��`�̉���Y"O։�aȌ�P'0P KT-3��ŋ�"Op�)  �`ț��R
Q�xT�7"O�x� �	DI*K<x�� ��"O��B�O�
���Z��!BؾH��"O�9��蝖RX�	IsH�e�I�e"OlY� X1J�x���+��g���"O2��@GU�
@Ƞ,Z\Ui�d"O�ݙ�3N�@��G;8a��"O�@ᰧяv��9�k�}H�}�s"OR	��� H�0i��r:��*�"O���-	�(�#�E݇8("!�"O�+���h��!��,��"Ony�nأW�"%h��H��P�*�"O@��Ԅ��� �E4.����f"O<� "b��x��KdgG�LP�d��"OhqCT��F �MRC�(5C���d"O� �y���} �C'	�#��d�D"O�4��$_�
��jD��+ ��'*O�xF��h߸-ɖ�ߌblE��'���yU�	��6yIf�أ_�0P��'/�!
���:����"]��=ʈ���O`xbB�.�M����⭟�Pɥ$�cf�� n���% �:���	���	�xa@0c�!ƕWo�����*��� ֌Mj`�<ZreN�q�z}r�L�[=x$a�@x�'�� :q�ùa��CA�bNx���M��%>8T���7 T>Y1Q��2}�,;'Ҏ����=�3i�ӟ���4A`�O*�6�N�z@tX��a�� c�I0e�"x���� ��ߟ��	�<����'�!7',���юI^��l�{8���޴-��iˮ�r�Ȗ�2t9A�P5�=��'��F�j����O2�'k�$!���?�ٴc�&�R���*`�V��*"|�0�:v�
1?�� W�&�B�sT�^�Y��SЩ1W���?�� Q�uΉ'��U�*��4lZ2q�*�0�a�0Y ���� 6_�̣���4:�c>�X�
�8��mW����@K�%��6-�G�gr�d�O�T�s�PL�"DE�ܸl*狓Df
�9��O���?�I֟h�>�⃅�s�&!�d/XT�2`�3�VO�'YL7�Ȧ����Mk����Yw'(Uxԣɍ������}�8r��O��d3(��,���O����O��ĉ������M�D�&��uΓ,c0  �*{[N����
]���
V��T�O��ȓ��r�h�Zt��2�mp�GBg���D,ڠ� �! �)�(p��i�tπ �v�$�<�r�1Tjm�ň���"Tf�>�bk��{ܴo7���'ؠ��5?>.8Q�'B�x��{b[�@P��I�f0x�'��<�ذG��Zġ��4a����' 6��O����h�'\2
��Cl�V�F"Ȍ4�0d�s��rB4���?����?I����?i���?�� �1^xI�2�XP�5�6�/&�Ƥp�OK��ґ �>ntcR�m�jEyrM����ʓ&S'�����m��ȁ`_ Q��F�+.��X�h �Zc���O��0�`�Ɋ#/40R�o��SF�Ր�.�$ٺp�BL��M;������O��ʧ(�l-�D��>CP	;��L5U��`�RO��V��.j8��#P���:�O���Q�	�-�'ifyЧ%�@?i�����]�Cp��i!��&�i���[�AFa�۟���Ο��g�S�Tf^9�S$O��}���2ly���0f�x�@↺Qs��々�g�l�<�t-�,T�	 1�ˢfN���]�PԊ #�L�WQ~�����yj�@�7�_ ���B����?I��i��7��O��'��͛�kE���D�K J����'��O��}�]�	�]��O�*_Vv<���̊l�������EA�4�Mk�)� ��`F$�2�
Ƞc�U?���)4��V�'f�Z>i+�&M��D�I����ը��I<x;A�/?�F�Y��U�@�H�Ɖ�#d.}��O�%�pX�n׍8 ��2)���iu�-ڷ�ڨ��9B�o[i���H��q���dܲp.���q˜�)L�5Z�h�A\�9��3��Ƅ���HK�ژa`-��(�s�iWi����²<��X��M�WӷqB�R$G��<�δ3�^_?q��ư>IP��*���ks)�6>��}� �_�'�X7����!'�D�պ��G�}"L�Q����}�`-
�I|�'�a{�h��   �   '   Ĵ���	��Z�:ti��:G���dC}"�ײK*<ac�ʄ��iZ"v-�(xrğ	"�6��++ 8�p�5L�����K��$�P�'�1o��M{��6��NP#�-�	��ZD���4H��R�Ws�BqK\�w5����ȀYg,���T�챷��-�V��L���1`u��L�Bh �K�;�vX���P��I�'��`���"r�Pq�'�� �a$+`v|�'H�UcI����`g�?g���f��]u�dR��,}��Ձ^�p��;}��U�}���C�(m���J�@ɤ|�$a�@
�8�(ʮ�# ��/*�{/�8���9������`����2+$\C���/�~�c_	(����K>Y�۝%D�$���v"�>���"�o�PU� l��Z�h�81�|�F7Gtv��I>!BD1s�t�HF��S�P��N�H�ܴr��բvhb��O���D�,n�X�RGU��.@�i@1띳W�k�ʿ0�H(p��Q�F�	��ۨX����Ɋ6Ǝ�qa��䰜'@�}���<Y!:�:�7 �Z``B�2�#��0R�zK>q`�OB��c�F ?���*A�!���X'5(V\�Eۆ/�W�K0�l�'��� ,����g-�\���m�Dӹ`�xx1b��ZXjS��%;�41x3��c�����yB���l������$��dԛ�/hH@Z�lކA�
�UJ�6V��U��1�U�c`�O��)�B��M�DF�kab�Ŝ[���3���4 �I%b�Ԕ�%�����'�Nd�$\uy�O�``iFJ�:{�Z90��7�hpW��xx�T�'`�'���'�t��n� p�e�^�Ld�sv�ޚGi���X@
 c�iޜ�#�i�|��#�ȃh����>5�̂3�M�?���ܸ`��5���ʶC��ic���TyBj�
����M>!D&��%ʊ�'�D�#�/K�5��F��6!�@�2L�M02T�:�dš
W��v�DN4M�X�&h�@o�e؀AL`+�`
��,D�L��   �  �E`��3�	��\
��4���AD	L�U����_��  q"Dᦵ�I��؇f�,6@T���Ɵ���ɟ\HXw#r�����y2���:z�hȑK'k��y`��sK��n�(��Aa@@r�-�3ғ1�D]sE�J61�A�6��'>Q���0�Y.WN�Cc�5jm\�sp�G���A�U�v$�(���W8e�f�Ä7XO�dв�g����_,vc���Ц�(��ΟX�      O  �  �  #   f&  �'   Ĵ���	����Zv�������@Q60"���5O�ȑC"J�+^��$E�/�*�˔ɐ�d`BdƄYy�\���S�\��Y8���5OR0�`�0��i���1{����&��a7��ZF"�C۪f��|0�I^v��8U��$[*�݊&��)���jV�Ia��RdAޠr検�cJ3> <i#n
5S��-�fbJ�2� (c\ ��"=E�x�K�J�T8�e�	D�YTL�>C��P"��?O
��$=B�0��n_�|h���O�(|����aX�؂!c�#n+�D��˘[��hpRe-D����S�Tip����G����KЮ,D���5F��,�Xi�B�"Q6���5?D��jץW%��DhMO�{g\)S��8D���H+D��d�N�]�H�Є�&D� �r.� Hl t��N�1;uF:D�H�gݽ��J� @�Q
�	��<D��Q0H�</�yRDN����&I6D��顄E*5�Э�C�ٔy�ҭpw�.D�p�S���p����%�����x�#)D�\��"Q��"d��Nڹ$12�p�)(D��@WD�E�H[��)eX�a��!D�|0��U�Z�)��˻K�<M�P#D��xu��&�x�3��W�Y,�X�o!D��Ac��?o��䢧J!^`!%D���v��=b^�!�6 5-���#�e"D�H{�V�^A����mM����c5D��)�L�0v�&�9g �,�z��r�3D��!��LQ�t���@�;9v��f�<D�|���A�jiPR�V�`$@E<D�x���T�I���zS?v�dc�l9D�8���C/h0(�D��3'����#O&D� �� �$*?�Kf��{� ���%D��0�m�0A�X�І��H���R� %D����CB�B�K3lr�BH=D��A���&I�EF��n>LA���9D���`V[&� ��A�4M"q �K,D�T	3jL$6�jؠ��N�R��c�(D� ȥ䄴4�,�(�2M�p���!D���!��"G�Ը5'�;(�2��W;D���1/A�T���)����2X���;D���	S�/�@Q!�h����4�9D�@1w�ܵ|�N���*�����&D�ȡ4!I{ز[DǙ+A�>D��w'�X��0q��o.�:ա1D���VN]R�(�q�Z�=�����o0D��P�M�kBh9$d��P��1D�\��H�(p*�1�o��lY���6A0D�����H��8�B�aĕߔ�1�,D�\!��G/�܊t퇞?�][��+D��iU%^�4,Y�Ʉ?g���6D�`��DQ�xOj� �@�KT<d`aK*D�I�$�s���յ�`���1�"D�����Q�G��"�V�n���e"D���(��P�����d�x�a�*D�Ds5��!A�b];��@�qS���(D��#���y�M09�hx��B5D���TH]gs8�����"�v���1D�����V�Oz�����%sR�4�+D�,`�*[�q����$)�� ����q�.D��!"��`��P����i�d�q$+D�t�q���hR��f���2�*D�\µo̪4a���^�H�a%,D���u��U�^ͱPA��]�(��*?D�<�e�ץY��u�6J:��7�9D� 1Cg��:y�p7%�,?�NE�VE*D������"B�p��E�0�b1�� *D��� RQA0`{%�N�Je��ï6D�`��Ϫ� D ��ٱi`x	2&4D�� ����ȕQ�R� ���A|���"O�uɆ�I�/�:L���[�o�:��"O����B<_�4�s�w�����"O8��ևJ�wb�E�E�1��I�C"O
�z�-�8Y�B�FY�7���f"O���%J�tE@�
х�"�\|kr"OHA1�cö+�z���ꨪ�"O�\�ч �'��ՑѪE�?�M�R"O:a�g#Z?���'�c1�DX�"O
�+'��(@���r�f�<a�鐡"OP�&Iʎ8E��v%�2�}�#"O
����ȃ�$�bgC�E,��p�"O8x��'�+Pڠ��U�R
(|Დ"Ob� ��X*����d��Ҍ%jP"O(��&�1S�09�M�.j;�:"OL�{�@Ҝ��Β-t �"OfmY�*�!U��$(��<��Qf"O�-��l\/P5���� �hc�Q"O~0�"I�
xvLhc���}�`86"OL����$hw$cׄ�-tX�'"O�}˔$\���8.�\|�|�"OV��֦ ;/�p�A2I=~����"OH`1"K̜!o^�աÉ8k� �F"O����N֎y����6@V�OR0���"O.���mU�&\Ɣ �^m �Af"O�r�(Fj,�#0mSf��"O>�`�C5}�~�a@�Y�bX.D�$"OP=��i��>�0��MN�\Y��� "O�0Jѭ>r�1�@\��Lq
�"O�E�2� �s� z����J���"OةdB7�4�@u����n���"OT��J�2~%�ċAy���;c"O� Zd�Oq�0���M|�A�"O�|�C%�5 2�&/��L�6��2"O\!��n�c� ��׸�V`jc"O�;V���2VlR`�ȘL����"O� F��2Nz�j�D	9<`T�$"O�,�vg�8p�H@D�G��u"O��&�Ӻi�auʜ�y���C"Ol-�Q@О|^�CB	��.k�Mqg"O<q*���-��bc���4x��f"O��lC�A20�����kM:A
�"O2P�u��sNQ��PB%���U"O�E��=�>�!�LJ�l���ӂ"O�E�r]�Ԙ�B^4�X�c"O��в�ߖ9�0�*�/3�,�*�"O�Eٗ��v�QQ�m���	��"Op�)���q�����Ίy�"O����h�+ 픍��d�)����"OB�Ym� �*{r�-bє�q"O��ʵ��f<8i�+2�x�"O��b��\�A��IY�j�X%f�+S"O68��-٫fh�a��ț#Y���6"O$� 4�R�/��Q��7+�0�"O�qaצ�S��)�f�5#K�]�&"O25O�>r�	������"O�ݩ��V4t-st@H����a�"O䤒�J_�=ۺ�1کnp��Ц"O�=��×6�6�Id M8^��H�"Op�zK�,&��5��,?r	z"O����2r����T�VY���"Oxmz4�OUJE[d�Ę�&��"OڜZs+�	BN	hPD]�ά�"O`X0�ߍB�|��U�Q,h�ְ�'"O� ��&�
�_e� �"���.��[�"Oa�a.݅!"�<��iM�>�B|�p"OmBqBد6RH�C��*��h��"O(�"$�_3.�F���;}М)�"Op��9!4L�rMC45D����"O�{���(���Xuキ[ u�4"OꕱC^@��E�W)IH��"O>T���?x]�<���7^R�;"O���0��M��,0QH��9Fp@�"O�<��N�uy��RThD�J �(�	�'	Thз"a��` �3���'\ ��g�N��d��L�,&p���'L~���Ù/{�Fթ�߲\��9�'&��l�e:�@A��Y�Z�<��'�����I7DٞY��c�l;
�'#h,
��Ł@xʍ�5�`h����'���eEaJ�E��2�  ��'~�h�Y=
�
� 憓�Ƶ	�'�邆ޡv�<}�!��20�I�'x��@dp.��pn�x�
���'�4�[7� �-��p�
i�2<p�'��L9〗7ur�2�!E2��'	lz���~�4��H���'D��c�
�a��A��vP���'��9K�o����:��].�:�i�'ܶ�[&�mqL�(� P�!Z���'��ԊH�kJ@�sꋙ	'���'�v�	S+׳2�j���KF`k�'�(�+4,݇&�RD��ݡGNUk�'y���Ƶ%��`�,�Eh���	�'�x<	t�Y��)�@M zƩ�'a �c�	��<&\Ԃ����n!��j�'N�BP卨?0PuF�ɅgNF��'D�9��h-�xyQ*�a�֙��'��9��J$&�����my�'�!�O�t�
�p�IM��-C�'��-#h�ov�5"QbҞ
���
�'�V�۱"6̀� N.<�`�	�'�XMS� Q1x	�ȑE@�:6t< 	�'�p�!�w]b$ZЀX%+�Z��'ƺ�[EL[<D<�i2�V�n��H�'#���k��f���aVl�Ҭ��'�zTْ��_�\�	�i�
�y�'C�p��Ɋ0����_�3�����'Zdy�V֠7J�e9�M���C�'�6ha����ԁ�#�cg���'(�u�O����zC����(��'�8��Q �6��C��G���'��x%�O�Y�J-�s�Ⱥu�$a��'��H�k��+�I�L��:&��'�,M��-la��Z7�!72c�'#Bpp$�*f��y$�-�(-�'͘u��'������-���'���C4�E#L,�Ht��f���'��db�T&�.�������P�'<6��6F��A��< FC��`ݙ�'��Ç'F	j�|�1��uL���'�F�)�*�����a]Sd���'d��!J�+/�L��%�Y�b�#	�'��M��L��"��e#��2�>�S�'�\U�WnLI��8�J�R�	�'](X�C�L�I��"qL 7H����'v�DXw,߫��(��/2��9y�'�h �DGϾQ�����=,�i��� �q:3PH8�)'N	P!���"O.L)�
_/K|����ċ�S�b�8�"O�=��/��d�RI�w�\��@9��"Ov��������0E�༵�A"O�̘&$��@Q��Y�"���"O�]��ʣb�Ե��	E�"B5{�"OR �e[R,�!],��%��"O�|�g����c�ūZ��4E"O q� �X.K-C��[�g���!)
���I`X���'Ί�YQM]5/9UJ" 2D��K%I$z�����![	2c�D[T�<D���u�ٲ2��T�4&ڿ�*��?D�h
�枴5��*6 W�#�:Ѳ�i D�p ʍ�R^��� C�D�X"N)D�Tv�|lva�Em������'D����e��.�~m�c!� Q�d`��:D���w+%���j�R뎸��7D�Pe�\[Xݹ��@
^��5D�lbL��{�ؕy� ف��bQ,3D��Q���~��4$2FjR|�D�1D��5�Ht��ej���
3���R�.D�8��&��2=��Y�mR�X:��z�E(D��"�B;ڐ����ܪQ�^x���8D���6���Pж�	�JCtp�8D����Å0Ͱ��%�W�^�4dXS�4D�|p!���:*z4�"��)H���D4D��x��<Cl����>n#4���$2D�� .��,�v��@&�F{��+�-D�$J�+��^�c��TT��d�=D��� ���2�;�h�Eذ���7D�4�-��F�\(�DY�@��*D��*��U8]��ykFX
n$"$���-D��!%MQ��x�T3�US#-D��9�c��=��@���	��ɩ�	*D��2�G�~��2#�٣��Y��)D�xaC�[;��uy���
h���q��<D�8`cK{�^�
��^�k���21B<D��J�k�8W��`�kB�#_����H6D�T� bZ% ��C��;��*D�3D�
Ʌ�BOv��d��/xrmcJ.D���� K�;4E�b�V�
1R��QD+D� I"<�,u��T�"5>E���+D�Ĩ��Y�x�4�R�5'�)���+D�����Y��/Q����,+D�����3���S0n,�0��*D�$�g`Ϩ?������`�����=D�@B�kͭ�ҡ��!��r�<}���6D��J�ߟd_�Xx�gκ�(Š�$3D�Xb�?`�l�c���$O�����n2D�T!6�̸Y).L�`	��`Lu�6<D��'&�K�̥G��c���J��:D���"h}���-��Mz�SC#D�\��X�������,'m�A�M$D��d��I`0�u��T��Q��6D���%�W�+��9Z�e�0�%���!�D��K�:8"F�)c4mqW���
�!򄒇�4m�&)�4��
`��6�!�D6D��8�wQ-�rP���
�!�Dߚr`������.j� EQ'��C�!�$�7��l �l[8Ff�*ՀV�!�$��'�\��V�-U�V
u!�$ "ض�##I�'"Q`��j�!���+z��� �am< c��5D�!�I
je�� C�`j�L��g��}C!�� Jh0�i�i{��h��kq$��"OD�Q6��9���AA_:!Z�q!C"O��$Q��-�wfT�m�l])"O|D��$ڤ<*ҹbf��'��K"O���q�ם#���W�N��U5"O���F�xm�s�[�:ԭ�"O$A����MBpi��M�ڕ��"O�Hҳ��O�p-���G�@|t<(q"O�K�菸-<4�J�-� ����"OZ)c��ќ#.��1g�4{�DI�"O6�0��
uͩ���_V�$�1*O*�����Dxfy��̸��
�'���,��-��4��*�r�9
�'�l5k�+��]3j��g�˘b*z�I
�'76 ����,}�iI D��&9��
�'cj���	#?^,P�N^b�i�'���zpd�)Hp$C��"ZT	(�'����C�R>�����US� %@�'�%�CKEײ�B�պN�@��'��|3�`::�����?5��P�'�.���V�i�N�@W�1k���'��;&��0�@�Cg���#k�@�'�Ρ���2�ִ궀^�J>�Mi
�'��I��gB�h�2�c"�<�4�Z
�'�~]4�H�GxP�Po�#:V�P�'��cgdE�?��Zq�6'�
���'����G�uٰ`D
N:�0�'�(=a&k�^xd��gFLbjp�'n�ˑf^/C�f'2��y��''t8� ��l�tq$;q����'�nt��₁)Ǫ(h���$J
�'�f\����V���#�4(��R
�'ӈ�s��G6#���蒠��LK
�'��؀�LqWf�*��_6.?��C�'~% �eT�S�&����-@�P!�'���ZFjF�����d��2ڥ��'�0�O�$i�6A@�{�l0�'��h��J=wA���E̄lH���'���������t��(1�]��'Td�wB�,��C� Ƭ�'��-�b�3!��RUK�z�����'h��	�O��^R5K��z0��8	�'�fUQ�$L�CKR�H��C=<TP�'�~-�u��72����O����'Hl���%ۏ>>V�2�9X��e��'��+d�Iw7 m�%��_ќ	��'�������zu�`���B�Th���'���FY�(��y'!�j���'�6�H�B �&�s"7����'̖��V��3\��(��Ɣ-)
�''����c�$>���GO�W6,�	�'���`�M`v�zf	��I.`11	�' ��!ʗH`�Y��ݝ>��1��'���fN�%R1za:��S).֤�
�'� l��A�a�������.�R\�
�'|�餪\�D��c�T�n�*
�':$e�d��sز���'Gk�B	�'3n�� �I @9���͒=�Q��'�V�q�,W�,�~ؙd��T�-j�')&�I*�l�Ka�	<c�t��'Cd����Ty`ri���0v�>ć�=�>���_"#�Hp���+<N=��~0<�&1@��`΍8�䜇��n� �
T(a��h�_4/4Ň�S�? �a�w)��� ܠ�H����g"O��ӡԄm
���/����"OjhXg�r6}��☠)sJ�t"O$�9ԃ%x6�}����{Y���"O�1ֈ�,�|"���!4L�"�"O��Ҳ(N5�,<�l���s'"Of��mܯA.X�T)^�%�N�u"O��Q��rK�S���_�4�ђ"O�\;C��� ��Ҫ�N d�H"O-	�c,B��p����/�#g"O�d6�kY��Jԓ�搫�iZ�<QaW�<4B��6I.�y�ŕY�<�gaߋM��UXbnK0a�����T�<�uJ�%f��Y��h�.c=��k�<YWcȧv�F�tH�_I��@3lFO�<��
^�$�*|;Ť̬$I��hC��C�<�7	^�aɸ5��a1>U`f�W}�<���,�6̡��Zy��҉�D�<A���j 5��g+��sҮIC�<Y�/�W�6��āύI�B�+Bgj�<)!̀�q���P���h�VPCu���<1��M�yʹp"�\�U<f[SHd�<����	N4��"��3�8-�E�Z�<�DF��&GҰ�І�1}����(GY�<!	�	_��Bԅ
0�1���M�<�sM�Qʤ���X�hUc��J�<a`ܢ�iz��ۄD�7��m�<�,��q��J��A,pN�p��^�<Y�:!PYR$�� K�H��QZ�<I'&�
'��! e�Y�iR�`�<id�r���BP�^^x�#�B�q�<�⮑ O�`��n	!X���A�<Q#�G�Sk�����<K�:�{�t�<���Ͻe%�; a�;(��|�&@J�<q@W�)��Qr�S��J�F�<Qq�	� �� `��-J,"��@�<��bN�w%J#�l֬hX0lcF�Jw�<��M�.L�G�Ч�	#p/�s�<Ya7P�|��$�!n(��b�o y�<�Gm�)��5�I�Y��Uj�,�N�<�G+Tx\��X��S�k��e��`�<1A#��rEb��Nʄ
|�iZb�B�	&DDH{�bM"M:����X�B��8��=�7�3-�|k4n�lthB�I/��6�Q��<dr���qHB�	&#�`�S������⤟�imHB�����o��[�T9�l<qD6B�	�T%��҆Z<6M0��R'tpDC�ɣz{z��v�$}�p��1� $�PB�ɉa�ʅ�f��8q���Q���6FDB�/D��&┈gC����SWi.B�ɜ^��	@�?7|����R�g�B�I�tV�w.��wɨ��%�-v0B�I�0����Ë��T�^�3��"�bB�I.;�8�C�m�6XY�O@}�@B�	��2�c�fޚ7�t2qi�naB�ɻq��%�f�g�	b��Q�d��C䉢qJ���Ն�SpΜK�iL�!s�C�>=�\m� ]�늰b��^��hC�=_1�+0��
K�(C�kC䉏S���r�NN�x  q���5@C�	� ����'#�%�pл��`�,C�3d����3��رN�3HC䉹�ց�c��
j�`��F=C�)� N�BTH�D`��G%/�6���"O*H��c�6"$� �!��N��r"OСX.R�U�M��_VF��6"O�L�UɄ�]��� *ܰP�
�"O��D/W�!x�R鐣Hy�r"O�`����/ M���=c�@ 7"O��CRgS@���M�(&M�"O�y�/U1�z����Z.�Xe"O�5ڢA� N��6+�5��c"O��� ��L�VI������\�W"O�[0�ۋ�@
ȞL�\ɪ�"O<��#��c�IY5�H�0�Hd#�"O LI2�U�pohEjA�ȝO��� "O@��t�  �   &   Ĵ���	����tH:9���dC}"�ײK*<ac�ʄ��iZ"v-�(x�A�	"�6�	M��r4G�g�R�YP��X�p��� M�Gmڥ�M+���&1�NM&C	�������͟xb5�^�y�,�Q��ϙg���+G�$��@F_�d��F\9�O�<�v!P;�"�jd�U"4E8��+&{ D���'�I���ҳ��($剏lW�,:��Ё��	@����K�@03"@	�~��g�y�L��R�(�7� -+L���Κ5����^5�p�^'k������Y�d��s�"�sSI��dJ�:>4)�5�l>%�����A�
�&=�}��)���8� S1_�Oڔ#�es��'��x��;8&����L��]�u3��&E�h�&�B$m��^�Ope9�l:�Ƙ
���T�B�[ n��(+�Ɵ�s�5���P���'���M�)[J̭��E�6��;5�	�
U�5�ݛk�L�Nᆵ��'f��	�ib/OV�ϧ5Y �z/��2�z0�G�ݪu�D�\�~��N>�gf �k����F�*?I�"�	���5ML3a��I����e�Jd���%5�I,.�ډH�3�À�ᖛ>�Zu2
�n[|�����#���ʇ�8��	��y�	BΔ���4�ƾ��E��M�Q��NU,ZޑYC5t��JU]�t�"��?�j�O�{�Lݙ��d�70��H �O:8�-)�FЂ_��I20��� �Ȣ����'��`�N����4�]��#���i&��Ѣ@L$��X��O}r�x��p�	�M�F6Z�{$��$g�2^@H��JF%����AL�3��V甊n�<�գ~�6���f�O\��l�f8�$h�E|��'����	2#H�|^ٖ'�NY[W#���iZm�Tf�\�I \�1��EX!n,�i�0�.dZ���b�֍O �O2]��g��+1O�zb�+G�[�h��l����I�`C�ɐn�� �  �Mh�eD�jf�,���R��u�F��y2H�	T�5Y�JL�Up�%aϬ�y�Xc�Vu���dS~�Di��0=�q�2��z>�yr!��^ˢ�Y�+�,İфȓ[4yȐ�Q:����cѾ&!  �=)0�)�I?\���9�A�'�$����=N�!�Q��Q,��!s��ߪUw舲�ቀj6Q>�0Ȅ� �k)@[�i��@�*F1�'�V�W	Q�[���Ib��cl��ڴ4�!�� r�X����mb�̾K;a)�'P�2`� [���3H��G���	�'����5R�	��!��C�Ȱ9���)�d!�j�K3�Z���t`t�̛�yrEQ�o�>hr@�N�	L��%�y�_�(>�M+U���2	�"��y�7լ�E���IH�1Nۅ�yb��=n�۳��X���f���yBK �B�R�z�dA0�(��y"�Bj� ؤ �`��}�3"��yBm�M2X��E"6T����K��y2ԁK �L@�&2#���h��y�Ǘ5`<�j�n��@��� �#�yR��֠���c݆bX�HfNҡ�yR��<��V&�V��%;@��,�y⎗��|��qȊK�ԍP� ���y��L�Qw�s7���G{!�F��yr,ޟ'"�c�@�>b��Ƞ
X��y���<�1t&H�3�6؃�@�.�yRj��?R�=�w��^D�\)e���y
� ��2#뚏A���_=9�ȁh"O��idJ5u�޽��lL�pG����"O촺�
0@���gś(AR t"O֘	��M� %<��8P�¸1�"O
�/5<�lq��κ�Tu��"O�	����6���V�Y�d�)t"O8�*wo�
c�2ȱ�D�8����"O0�`!��MнB�D��U��R�"O�H���];�Y,e��ᱬ�y��Лx�>����1��죡�
��y�]�v�LR�l	'4�A�F��y��A�,h�7�B� ��5��ޭ�y�&7]���A��~�H���ʓ�y2)۽/�� Z"�&.�đQ�G�y�/�]e��S�� �b��sd^�y�T2>�:�i� �&��Ǌ<�yR	��t��dT8J�p�&�L��yσ�}��%ِ��$`��@&H��y�/��VQV���� ����E$Z��yHH�JTX�

"��Q��Θ��y2ą�	D��W��u��u�ś,�y2� :\�j��VL�iIB�@v��1�y"c�QsB�+�g�$N��( 7�Q��y�ޣ>!�}��� M>��#�>�yBc�*54�	��;?�L ���C��y£@�2�Ҵ!'H�5'�G$�y�nƈua����/\�#����c��yM^)�f]�b�1�~�p2���y�	�0+�l�1��4��H	7
��yb }���bK�0��E��dծ�y�-S%FDlE����v��IQ���ybL_$N��Ъ���Z��-�0 M��y�mJ�vh��ԎN��0A��y�ꔚN�F1�Ǉ �H$�6⍐�y+�01e�qq��F!u[z��6H.�y�DI�3�"�1/��v��0#Wa��y��Ө\Y��k
�5h��Ă�y"ޱTb̒j�BѰ�N��y�J�%�J5"��Ği8^�`�)��y2'�t��� ��@�l���(ݪ�y����J��H��Ҕfu ��$C���y¤�e��B�ӄr7�dK���y2K��%�
a`������j����y�)�.�F!2�i�:~d ��Q��y�21���׉K�F�Bը�I��<)��E68�JL�F��r�j�	�P�<i��m�5��I���e���C�<��\*E0�����5i<�£N�Z�<��d�5#�H��-��tkt�Ͼ�y��^�ؐ!Ҁ埰<m�̛��y�
Ͻq�@ѤH�&��M����y�i�x��x����&�����yb�޹4 T  �   )   Ĵ���	��Z�:t�==���dC}"�ײK*<ac�ʄ��iZ"v!�(xrğ	�t6��<q'��F��)�t����,v\Qw∈/`j�m��M3CK�U�뮈+eh��	�l������x{3����U�M8J��TA��z],�P�Z�@��k��[F�x�H�P�ƀ�T,���R�;[�쐈�ǯ��,Eа9�'�؈����E��<y�G��$[d`�<95L\C�)y"�O�D,�2ʁ�j�T��H7&��>�u	7�
�nO�bZܸ#�)&�0�i�O�#��H�b�2k��zJ��
��P�mT�Q$���&��)e�,��'-_���!�H�C�,��"��ebvU��z�Q�eH�@?��9O2�����ԟ�e�����HL*�̏�-!U�G-��s����J>i��_���%�Pc�H�J�H����.n|��a��)p�>k ��-�?���'��<3P<N����*OȈ��NG�@�8ɲ[c'�ash�_&�QQ�L'')��k�O�O����"����d��<������9��F�/w%��CU�S��E)���@����U��_�	�R�y��HX��3}���t�?��b�H�M*�(b���a��O�h"�%pb�'�E�Q'L��	�m�Ճ�fc�`1U$��A�0��J��.b���?1�D��d@�)O�	k��#���(Ik�	���]��NT ug�!a ˴<�c�>;��$��kpm�zX��	-r��Ƀg��$@�d���=v���c�vdZuCp?�F:O��"����ԟ�eZHQ�;b���!e�}�:��	R��XC�O|ORY�K<y4L�z�d���ݑ �P�m̑-���A�F0{<���N	5��\I2ᇣu�E��B/x墐�;7F�l9r	E�>?2� 0Zx����c��xf)�#��'�T�$� �E��CP�T�Oh��A�R`i��

��@�6d�I��a �|�Aܟ/д��y2��)��S3�QT����[N7��1"Of)B��  ���r�N�*��dr"OH@ö�Nlj�q�(X0zb���"O��Pcڛ\���T�Y���f"Oڠ#���>X�S	D�0�b�"O01��+�}�\A%�t�p4Z"O`��kѴ���CԦ��lĴ��"OQ
҃x~���K� �`	ɱ"O���י�\@扛�1�0��0"O�����ct�4z���u�>�U"O�9�
�8a�H��F�      O  �  �  #   f&  �'   Ĵ���	����Zv�������@Q60"���5O�ȑC"J�+^��$E�/�*�˔ɐ�d`BdƄYy�\���S�\��Y8���5OR0�`�0��i���1{����&��a7��ZF"�C۪f��|0�I^v��8U��$[*�݊&��)���jV�Ia��RdAޠr検�cJ3> <i#n
5S��-�fbJ�2� (c\ ��"=E�x�K�J�T8�e�	D�YTL�>C��P"��?O
��$=B�0��n_�|h���O�(|����aX�؂!c�#n+�D��˘[��hpRe-D����S�Tip����G����KЮ,D���5F��,�Xi�B�"Q6���5?D��jץW%��DhMO�{g\)S��8D���H+D��d�N�]�H�Є�&D� �r.� Hl t��N�1;uF:D�H�gݽ��J� @�Q
�	��<D��Q0H�</�yRDN����&I6D��顄E*5�Э�C�ٔy�ҭpw�.D�p�S���p����%�����x�#)D�\��"Q��"d��Nڹ$12�p�)(D��@WD�E�H[��)eX�a��!D�|0��U�Z�)��˻K�<M�P#D��xu��&�x�3��W�Y,�X�o!D��Ac��?o��䢧J!^`!%D���v��=b^�!�6 5-���#�e"D�H{�V�^A����mM����c5D��)�L�0v�&�9g �,�z��r�3D��!��LQ�t���@�;9v��f�<D�|���A�jiPR�V�`$@E<D�x���T�I���zS?v�dc�l9D�8���C/h0(�D��3'����#O&D� �� �$*?�Kf��{� ���%D��0�m�0A�X�І��H���R� %D����CB�B�K3lr�BH=D��A���&I�EF��n>LA���9D���`V[&� ��A�4M"q �K,D�T	3jL$6�jؠ��N�R��c�(D� ȥ䄴4�,�(�2M�p���!D���!��"G�Ը5'�;(�2��W;D���1/A�T���)����2X���;D���	S�/�@Q!�h����4�9D�@1w�ܵ|�N���*�����&D�ȡ4!I{ز[DǙ+A�>D��w'�X��0q��o.�:ա1D���VN]R�(�q�Z�=�����o0D��P�M�kBh9$d��P��1D�\��H�(p*�1�o��lY���6A0D�����H��8�B�aĕߔ�1�,D�\!��G/�܊t퇞?�][��+D��iU%^�4,Y�Ʉ?g���6D�`��DQ�xOj� �@�KT<d`aK*D�I�$�s���յ�`���1�"D�����Q�G��"�V�n���e"D���(��P�����d�x�a�*D�Ds5��!A�b];��@�qS���(D��#���y�M09�hx��B5D���TH]gs8�����"�v���1D�����V�Oz�����%sR�4�+D�,`�*[�q����$)�� ����q�.D��!"��`��P����i�d�q$+D�t�q���hR��f���2�*D�\µo̪4a���^�H�a%,D���u��U�^ͱPA��]�(��*?D�<�e�ץY��u�6J:��7�9D� 1Cg��:y�p7%�,?�NE�VE*D������"B�p��E�0�b1�� *D��� RQA0`{%�N�Je��ï6D�`��Ϫ� D ��ٱi`x	2&4D�� ����ȕQ�R� ���A|���"O�uɆ�I�/�:L���[�o�:��"O����B<_�4�s�w�����"O8��ևJ�wb�E�E�1��I�C"O
�z�-�8Y�B�FY�7���f"O���%J�tE@�
х�"�\|kr"OHA1�cö+�z���ꨪ�"O�\�ч �'��ՑѪE�?�M�R"O:a�g#Z?���'�c1�DX�"O
�+'��(@���r�f�<a�鐡"OP�&Iʎ8E��v%�2�}�#"O
����ȃ�$�bgC�E,��p�"O8x��'�+Pڠ��U�R
(|Დ"Ob� ��X*����d��Ҍ%jP"O(��&�1S�09�M�.j;�:"OL�{�@Ҝ��Β-t �"OfmY�*�!U��$(��<��Qf"O�-��l\/P5���� �hc�Q"O~0�"I�
xvLhc���}�`86"OL����$hw$cׄ�-tX�'"O�}˔$\���8.�\|�|�"OV��֦ ;/�p�A2I=~����"OH`1"K̜!o^�աÉ8k� �F"O����N֎y����6@V�OR0���"O.���mU�&\Ɣ �^m �Af"O�r�(Fj,�#0mSf��"O>�`�C5}�~�a@�Y�bX.D�$"OP=��i��>�0��MN�\Y��� "O�0Jѭ>r�1�@\��Lq
�"O�E�2� �s� z����J���"OةdB7�4�@u����n���"OT��J�2~%�ċAy���;c"O� Zd�Oq�0���M|�A�"O�|�C%�5 2�&/��L�6��2"O\!��n�c� ��׸�V`jc"O�;V���2VlR`�ȘL����"O� F��2Nz�j�D	9<`T�$"O�,�vg�8p�H@D�G��u"O��&�Ӻi�auʜ�y���C"Ol-�Q@О|^�CB	��.k�Mqg"O<q*���-��bc���4x��f"O��lC�A20�����kM:A
�"O2P�u��sNQ��PB%���U"O�E��=�>�!�LJ�l���ӂ"O�E�r]�Ԙ�B^4�X�c"O��в�ߖ9�0�*�/3�,�*�"O�Eٗ��v�QQ�m���	��"Op�)���q�����Ίy�"O����h�+ 픍��d�)����"OB�Ym� �*{r�-bє�q"O��ʵ��f<8i�+2�x�"O��b��\�A��IY�j�X%f�+S"O68��-٫fh�a��ț#Y���6"O$� 4�R�/��Q��7+�0�"O�qaצ�S��)�f�5#K�]�&"O25O�>r�	������"O�ݩ��V4t-st@H����a�"O䤒�J_�=ۺ�1کnp��Ц"O�=��×6�6�Id M8^��H�"Op�zK�,&��5��,?r	z"O����2r����T�VY���"Oxmz4�OUJE[d�Ę�&��"OڜZs+�	BN	hPD]�ά�"O`X0�ߍB�|��U�Q,h�ְ�'"O� ��&�
�_e� �"���.��[�"Oa�a.݅!"�<��iM�>�B|�p"OmBqBد6RH�C��*��h��"O(�"$�_3.�F���;}М)�"Op��9!4L�rMC45D����"O�{���(���Xuキ[ u�4"OꕱC^@��E�W)IH��"O>T���?x]�<���7^R�;"O���0��M��,0QH��9Fp@�"O�<��N�uy��RThD�J �(�	�'	Thз"a��` �3���'\ ��g�N��d��L�,&p���'L~���Ù/{�Fթ�߲\��9�'&��l�e:�@A��Y�Z�<��'�����I7DٞY��c�l;
�'#h,
��Ł@xʍ�5�`h����'���eEaJ�E��2�  ��'~�h�Y=
�
� 憓�Ƶ	�'�邆ޡv�<}�!��20�I�'x��@dp.��pn�x�
���'�4�[7� �-��p�
i�2<p�'��L9〗7ur�2�!E2��'	lz���~�4��H���'D��c�
�a��A��vP���'��9K�o����:��].�:�i�'ܶ�[&�mqL�(� P�!Z���'��ԊH�kJ@�sꋙ	'���'�v�	S+׳2�j���KF`k�'�(�+4,݇&�RD��ݡGNUk�'y���Ƶ%��`�,�Eh���	�'�x<	t�Y��)�@M zƩ�'a �c�	��<&\Ԃ����n!��j�'N�BP卨?0PuF�ɅgNF��'D�9��h-�xyQ*�a�֙��'��9��J$&�����my�'�!�O�t�
�p�IM��-C�'��-#h�ov�5"QbҞ
���
�'�V�۱"6̀� N.<�`�	�'�XMS� Q1x	�ȑE@�:6t< 	�'�p�!�w]b$ZЀX%+�Z��'ƺ�[EL[<D<�i2�V�n��H�'#���k��f���aVl�Ҭ��'�zTْ��_�\�	�i�
�y�'C�p��Ɋ0����_�3�����'Zdy�V֠7J�e9�M���C�'�6ha����ԁ�#�cg���'(�u�O����zC����(��'�8��Q �6��C��G���'��x%�O�Y�J-�s�Ⱥu�$a��'��H�k��+�I�L��:&��'�,M��-la��Z7�!72c�'#Bpp$�*f��y$�-�(-�'͘u��'������-���'���C4�E#L,�Ht��f���'��db�T&�.�������P�'<6��6F��A��< FC��`ݙ�'��Ç'F	j�|�1��uL���'�F�)�*�����a]Sd���'d��!J�+/�L��%�Y�b�#	�'��M��L��"��e#��2�>�S�'�\U�WnLI��8�J�R�	�'](X�C�L�I��"qL 7H����'v�DXw,߫��(��/2��9y�'�h �DGϾQ�����=,�i��� �q:3PH8�)'N	P!���"O.L)�
_/K|����ċ�S�b�8�"O�=��/��d�RI�w�\��@9��"Ov��������0E�༵�A"O�̘&$��@Q��Y�"���"O�]��ʣb�Ե��	E�"B5{�"OR �e[R,�!],��%��"O�|�g����c�ūZ��4E"O q� �X.K-C��[�g���!)
���I`X���'Ί�YQM]5/9UJ" 2D��K%I$z�����![	2c�D[T�<D���u�ٲ2��T�4&ڿ�*��?D�h
�枴5��*6 W�#�:Ѳ�i D�p ʍ�R^��� C�D�X"N)D�Tv�|lva�Em������'D����e��.�~m�c!� Q�d`��:D���w+%���j�R뎸��7D�Pe�\[Xݹ��@
^��5D�lbL��{�ؕy� ف��bQ,3D��Q���~��4$2FjR|�D�1D��5�Ht��ej���
3���R�.D�8��&��2=��Y�mR�X:��z�E(D��"�B;ڐ����ܪQ�^x���8D���6���Pж�	�JCtp�8D����Å0Ͱ��%�W�^�4dXS�4D�|p!���:*z4�"��)H���D4D��x��<Cl����>n#4���$2D�� .��,�v��@&�F{��+�-D�$J�+��^�c��TT��d�=D��� ���2�;�h�Eذ���7D�4�-��F�\(�DY�@��*D��*��U8]��ykFX
n$"$���-D��!%MQ��x�T3�US#-D��9�c��=��@���	��ɩ�	*D��2�G�~��2#�٣��Y��)D�xaC�[;��uy���
h���q��<D�8`cK{�^�
��^�k���21B<D��J�k�8W��`�kB�#_����H6D�T� bZ% ��C��;��*D�3D�
Ʌ�BOv��d��/xrmcJ.D���� K�;4E�b�V�
1R��QD+D� I"<�,u��T�"5>E���+D�Ĩ��Y�x�4�R�5'�)���+D�����Y��/Q����,+D�����3���S0n,�0��*D�$�g`Ϩ?������`�����=D�@B�kͭ�ҡ��!��r�<}���6D��J�ߟd_�Xx�gκ�(Š�$3D�Xb�?`�l�c���$O�����n2D�T!6�̸Y).L�`	��`Lu�6<D��'&�K�̥G��c���J��:D���"h}���-��Mz�SC#D�\��X�������,'m�A�M$D��d��I`0�u��T��Q��6D���%�W�+��9Z�e�0�%���!�D��K�:8"F�)c4mqW���
�!򄒇�4m�&)�4��
`��6�!�D6D��8�wQ-�rP���
�!�Dߚr`������.j� EQ'��C�!�$�7��l �l[8Ff�*ՀV�!�$��'�\��V�-U�V
u!�$ "ض�##I�'"Q`��j�!���+z��� �am< c��5D�!�I
je�� C�`j�L��g��}C!�� Jh0�i�i{��h��kq$��"OD�Q6��9���AA_:!Z�q!C"O��$Q��-�wfT�m�l])"O|D��$ڤ<*ҹbf��'��K"O���q�ם#���W�N��U5"O���F�xm�s�[�:ԭ�"O$A����MBpi��M�ڕ��"O�Hҳ��O�p-���G�@|t<(q"O�K�菸-<4�J�-� ����"OZ)c��ќ#.��1g�4{�DI�"O6�0��
uͩ���_V�$�1*O*�����Dxfy��̸��
�'���,��-��4��*�r�9
�'�l5k�+��]3j��g�˘b*z�I
�'76 ����,}�iI D��&9��
�'cj���	#?^,P�N^b�i�'���zpd�)Hp$C��"ZT	(�'����C�R>�����US� %@�'�%�CKEײ�B�պN�@��'��|3�`::�����?5��P�'�.���V�i�N�@W�1k���'��;&��0�@�Cg���#k�@�'�Ρ���2�ִ궀^�J>�Mi
�'��I��gB�h�2�c"�<�4�Z
�'�~]4�H�GxP�Po�#:V�P�'��cgdE�?��Zq�6'�
���'����G�uٰ`D
N:�0�'�(=a&k�^xd��gFLbjp�'n�ˑf^/C�f'2��y��''t8� ��l�tq$;q����'�nt��₁)Ǫ(h���$J
�'�f\����V���#�4(��R
�'ӈ�s��G6#���蒠��LK
�'��؀�LqWf�*��_6.?��C�'~% �eT�S�&����-@�P!�'���ZFjF�����d��2ڥ��'�0�O�$i�6A@�{�l0�'��h��J=wA���E̄lH���'���������t��(1�]��'Td�wB�,��C� Ƭ�'��-�b�3!��RUK�z�����'h��	�O��^R5K��z0��8	�'�fUQ�$L�CKR�H��C=<TP�'�~-�u��72����O����'Hl���%ۏ>>V�2�9X��e��'��+d�Iw7 m�%��_ќ	��'�������zu�`���B�Th���'���FY�(��y'!�j���'�6�H�B �&�s"7����'̖��V��3\��(��Ɣ-)
�''����c�$>���GO�W6,�	�'���`�M`v�zf	��I.`11	�' ��!ʗH`�Y��ݝ>��1��'���fN�%R1za:��S).֤�
�'� l��A�a�������.�R\�
�'|�餪\�D��c�T�n�*
�':$e�d��sز���'Gk�B	�'3n�� �I @9���͒=�Q��'�V�q�,W�,�~ؙd��T�-j�')&�I*�l�Ka�	<c�t��'Cd����Ty`ri���0v�>ć�=�>���_"#�Hp���+<N=��~0<�&1@��`΍8�䜇��n� �
T(a��h�_4/4Ň�S�? �a�w)��� ܠ�H����g"O��ӡԄm
���/����"OjhXg�r6}��☠)sJ�t"O$�9ԃ%x6�}����{Y���"O�1ֈ�,�|"���!4L�"�"O��Ҳ(N5�,<�l���s'"Of��mܯA.X�T)^�%�N�u"O��Q��rK�S���_�4�ђ"O�\;C��� ��Ҫ�N d�H"O-	�c,B��p����/�#g"O�d6�kY��Jԓ�搫�iZ�<QaW�<4B��6I.�y�ŕY�<�gaߋM��UXbnK0a�����T�<�uJ�%f��Y��h�.c=��k�<YWcȧv�F�tH�_I��@3lFO�<��
^�$�*|;Ť̬$I��hC��C�<�7	^�aɸ5��a1>U`f�W}�<���,�6̡��Zy��҉�D�<A���j 5��g+��sҮIC�<Y�/�W�6��āύI�B�+Bgj�<)!̀�q���P���h�VPCu���<1��M�yʹp"�\�U<f[SHd�<����	N4��"��3�8-�E�Z�<�DF��&GҰ�І�1}����(GY�<!	�	_��Bԅ
0�1���M�<�sM�Qʤ���X�hUc��J�<a`ܢ�iz��ۄD�7��m�<�,��q��J��A,pN�p��^�<Y�:!PYR$�� K�H��QZ�<I'&�
'��! e�Y�iR�`�<id�r���BP�^^x�#�B�q�<�⮑ O�`��n	!X���A�<Q#�G�Sk�����<K�:�{�t�<���Ͻe%�; a�;(��|�&@J�<q@W�)��Qr�S��J�F�<Qq�	� �� `��-J,"��@�<��bN�w%J#�l֬hX0lcF�Jw�<��M�.L�G�Ч�	#p/�s�<Ya7P�|��$�!n(��b�o y�<�Gm�)��5�I�Y��Uj�,�N�<�G+Tx\��X��S�k��e��`�<1A#��rEb��Nʄ
|�iZb�B�	&DDH{�bM"M:����X�B��8��=�7�3-�|k4n�lthB�I/��6�Q��<dr���qHB�	&#�`�S������⤟�imHB�����o��[�T9�l<qD6B�	�T%��҆Z<6M0��R'tpDC�ɣz{z��v�$}�p��1� $�PB�ɉa�ʅ�f��8q���Q���6FDB�/D��&┈gC����SWi.B�ɜ^��	@�?7|����R�g�B�I�tV�w.��wɨ��%�-v0B�I�0����Ë��T�^�3��"�bB�I.;�8�C�m�6XY�O@}�@B�	��2�c�fޚ7�t2qi�naB�ɻq��%�f�g�	b��Q�d��C䉢qJ���Ն�SpΜK�iL�!s�C�>=�\m� ]�늰b��^��hC�=_1�+0��
K�(C�kC䉏S���r�NN�x  q���5@C�	� ����'#�%�pл��`�,C�3d����3��رN�3HC䉹�ց�c��
j�`��F=C�)� N�BTH�D`��G%/�6���"O*H��c�6"$� �!��N��r"OСX.R�U�M��_VF��6"O�L�UɄ�]��� *ܰP�
�"O��D/W�!x�R鐣Hy�r"O�`����/ M���=c�@ 7"O��CRgS@���M�(&M�"O�y�/U1�z����Z.�Xe"O�5ڢA� N��6+�5��c"O��� ��L�VI������\�W"O�[0�ۋ�@
ȞL�\ɪ�"O<��#��c�IY5�H�0�Hd#�"O LI2�U�pohEjA�ȝO��� "O@��t�  �   (   Ĵ���	��Z�:t�0=���dC}"�ײK*<ac�ʄ��iZ"v �(xrğ	"N6�V�:�p| `b_�d�vp�f�K�I�>���� &�4mZ!�M�b�R����#�(�I*e^x�	럤@P�M�B��$x-M���H�-�	IK+L����_<\S�� �[��,#p�d"�7Sl2�dN�>��9*��>%�N�Q�ODi7��JJ�m*O&|(�`� S��@�,O�1�dJ@�W/�Ц��MJ�k���.��`��K�X�d�B*�D�
W^���3x $��F��H�y�R��A�$mbR'�!n"�'AJ��a�	@���'�~X�ѡ�T���g�Y%�O�]Bx$رBC�-�D
�H�j���Od�S�2��K�<�'!����mE1Jo�u�W.Zd-�'.%��O��(�����'�8TJ!J��]�	�C�̟�6!p�P�V>lYᖧ�Oޱ��dXYNT��'�<1�(S/[f�8a�{�)Y�hF.D�f�B��;!2J�	`��?��N�"-����Dh󤑚.�]�')&�FlP�kw��Q%����D2!cX�ɠ)����'0��E&M�V�^I�'��q�DW<s�
Y(�d_��8(3p��wm*�k�5?��^��A�|b�G����jI�\r�ʔ�8�n��&��TL`5�ҥ2x���k?q&2OR�"e(S���ԟ.�UZ�k�ƛr��NPJ�Q�EŸtY�˓��@ �A�	�<!rXX�aq��2W�T;�=��&�?���`�ã>��鄡����_��DBa<<�.O�)F�)S�#H4�E*Z'CJ�@� Ln9��O`O�8hK<QQ^�`���I�K��<������6��DQ���u � �{�t��s�G�/�N�(�D�,��^/�< ��0l�I�B�F-iE!ٔ^Lݨ��9Q�t�(P��x�?` ̕�W�>I��A 󼭘KϤ������'7l�`+1�Y^�ɱOO��"�3执dx��j戙2�V�#ε2�H0d�e�<��
�6 2  �7�<�vVi�A��9
Ā(H��m��Hw��7���`,(?��+�;N��K� !?*	�t!]�	�������<'	H1	��Hܝ���ٹJ��r�T#=(��]������ӥ$�6�¤�T�Ј)�a��.mBL¬Olz!xu�`��ɉ�DS tYd��po�e�� �M���z��
�H	H�O��"0���@�踓�����+qD�,
�aY$.��#��U*��,6�FL����������Od��7B�?������l�"�؇BŹ �`,if��n�l��@�N�-\�pic�@膈V8��w���ti�@�h�v���I	~/Xx� ų�&l+%)�1;l�
 B,��&0;n�"@B�%nH{�oôV��|*��(*�H���ĽL�a�1��9���Z��7
��ôM����[1*�.TzI� `;I�u��Y����%W���d��q"�U�U�@�G&��A��_	XU�-#�"��Z��)���Ꙩ%�Y�u(�am��=�B K�B�?��#��ŀ@8(�$��r	�4�r���,H� B jL�<q7��+�����*�ŨO$������ş� ҢH�j
1|Sθ��`��b��2Xb�S�Eٽ,lJ�y �òR��F�
�WV��FE�	v�y���^&����I1���%F4��E}��8K������n]x�3j�
RƄ+��v]<��в4б�dC�5�҅�ݴF[
r�&C;s��L�B�8v����Q"cb$�[goH�,����3@VA��m��Qn�U9K>�&�%Qm�My#+�<p-qT/P��u�It_��2OLP԰EoJ�>d�	���������dĎ_�������g�\��1�HD^��eo
�?g�9�mU�����+�`XxAœ��ī���]�����KGY&5���?,�쑀Um�-.�vllZ%&���we_�����%�V�3�L8�A�Z�Lr�����1��
c��޼݂����>����A�.��OZ*7i Ґ�K�'��"8�)k�Ň"v�DYA�m?Wx���c1!Pd
'iU#֊�kՇ�"9�!KReǣt�B]��-�#�:d��DG�cg�A�5���d�E~�A�'8�SM-?Ⱥ�#�#6�ʢ!� W�y���֨#�l�A�C#*�9 uA��f�j�*�&?�,�!P�Q�a��* �f�Y���S���Hq��#���2(��'��#���3+���bU�5&�Hyk��R�I��W�����@��IVJ ��~B�P�ą˺+d�ED�r�x��g��LP���2�KWJ(
��?G�ɧL�j�ٗHسE0A�&�A�du�TOVy����R�n�dti�.�J�~��hY�O"a�vL@�f}�4V���A�
�E��a�Tl���R��0�X��Ԩ T��O��q���A!�ֹm����7�O��; A�Q��Yz� >�ȱѶ���e`���F�퓑)]�mW$�#XwB�Kw�1�䀄y��@�C��J�eqJ�m_�!ⵈIdy�))G�iY�b���~�J1Ҡ�K;E�!�$��<@�F ؑ�ǀo��\׍�t��{����`<��H�p�fV�*��J��'�!����T̅2���/(������ �����5�ٹ�	�?���f�H���L�TMߘGd0`���`͌jy�H�^F���S(5Y��S�]b��XSHY�<��\�%Kh��9`\�1��٩��̶_��$*3&��~"�N�c��I���)Y\i9�,�b���m�:t�m!�C�,C��"�<1�z���ǞV5����d�� ��'8�*�����Z�*E��b�k��3B?/t�5�E�S�H$������?�bg"X�,��x�Tu:g���O�H�ņ_��ꉻ�k�%vJ��$��&Ya�%�`�8y���N�T������;m��(�慮}���z�lۆh��Ő�N"�?ч]�c��A�mN���$ۉj<�58�F
>7�v��U��k����߂Gg��3�JF]����^{"���,�Ȥ�Q�/f��E�Ƃ[�h�	c�:(״����*z��5�n7L��*O��s��x��%$�F�G� 5qĀ�`G)H�Bdvy(w�Bn4*�8"=?�`�is����#Hp<�erb/�Z�)�[�I9��$c���F-�lD�Ѐ�70����7&�	k������a�|cJ�ޢr&Ĵi�|�X��Rк�1U��=0dFH�`���FA�q��
~,4u�&�(�+�D��A�`�'BR+�e���CK�U[�@J|/2})��j���s��Q����DDP)@�t��LG4
��ea���7��J��
p��u�0/AN<`cɀ�])�B��Md�rp흅i@r\��Ó�1,�|�	���yЦD�&_7.Y��O乚�	�8XP��2�ͳ��5Y�*z�̙[��U;.�����ؐ����\9XR������1-�L�dEٜU�=�0�0O�0\��5��8!`�x�(B<<�x	�G�$\�B`�1cA� .͗'�܌�Ђ-�$C6DO;��P�K�;#X��ON�s�.��P �*'��yV�߇GVu��Q3\�yB��@FQ�1�1[�PB�)�upʱ:�)~?2=![����Ws}ҁB�M�*x1,��: ^�](E�ܼ�g#1u��OA��AS���acC/�@�H>�Q��+�T �dP3_$���h�;.h��H	�5O�DQ����!=:�z���f�I�8Ԍ�s!*%���ap/�S�'���9PN�Lu{C��{ ��bY[���52�DQQ���p���a�N�6
Jq�;^H�0 �??r�A���&aj�m����qq^а,�/�`�:�s�EPv����[�&�({č@3$^ q@7���m۬��"��C�bQ�s�4����-�t�A0#�ܹ"�N@�V��0&ڒ	�l�ZϓU���F��z�E-��f�x��F%
�J=t��6/&X�~�؇��,hY�`���k�tt�u��}�lݲ�E4L3nŁ�/�g�� �@��*�4�>�� � �ftIx��|�@�efa F�&��Q�Q�x(3���bҪ`���F�V�X�8f�>Arr�i��P��dH`%�EqgF�C�gV�� �� �'O�5أ�1�,L����0G)��PvD݁8p� SL��+nC4cD��#�3�(H��A�C"��F$�9`r����ʻ�B����(�e���x��M�?�<���۞.�d���RQ^�𚃌?|_���"iVjH,�`5�.:�:�oZ�?Y"�
bm�$�����gȖ-^�a�	�:t��ݑa��baz ݺV��Ԉ&��3@�d�#)����эK������<:�����Z02�������`hٓC��1[��H����O�<�!"��mw �1#�,��)��d�s�� I�EَCi�#���lh!G��5Z�7�3�>�!nDo68�Z"N�TFr6m'c9ԥ�0mGRAԕ0��(O�)����$qƢ[�N0vU��Zh*j%1�i�O���4�J:�=��BV��y���M8d}�4# m!:EXM�C�8� ��e��kD�!�����s�MI��48'`R;A�Ll� ��8ٖHK��'"�3��E����#ѭ	5�yZw���;:���;�A7���0�J_�BtQ��H�4aG�S&�TI�#�ɼ%���r���t>*I9�̕�<���韘���I�a� ��>���SL��=`�A 
�bqP��o8� ��a�G�󄈵#�00
6&J1%�İ�-Ëj��$�#ag�kb���9�4����
�S~����i�:<��Rc�Ià��@;���'�D�T��ͅ:|g��A��H<�'+G�@\0��O��2Eb�'c	�#�U#N"*��J�S�Tj �jзmꀩ[!�v�<�M\=;m��B1#тlÒ���<�ì[�.,6�"~ 鐛XQ��֬'�|�:uFr�<�A���~��dQ��B3a�l�i�<Y�M�)�j�;%(Ƌ|��Y�B�q�<9Љ�M�2	�拀t�A 3��r�<�pL�"C�hձ�GS XF����l�<��@R�6�u��M� ݢ�0oMG�<!�D�Q��)QǤ��Rp�<X�}�<�G��c[�d���16�p�fu�<	&˞~ޠ�1��c��y+D��n�<i���*���J�bڐ[��5ӵ)�C�<١�Z��5���]�נ�2�o�C�<��.ʊ/�(�1�A�r�4i��'s�<Y��>	��)pD��~��pnn�<�#��&��8�)��N�9a�V�<�Â��T%� K&oV�e��T�<��J�u)�ӓ�A��l�*�D�y�<��/�)0�AaB�,/�`�Q�)Ew�<A�	�1�y���(�����Tn�<yA�Y.\�f� &C"��8�mLj�<�6aܯ�	��N�+T�l�B�e�<9�'�z�9#���s^S�[N�<9�!��4_���'�!1��`X�@H�<���� *Y<�j�ៜS��[�CM�<!$��I� E%"��RSЀ�n�I�<	��O��\u���En|���So�<A7Ⓗ���X�$����A��NDd�<9�'�](�q�ŧT%]ܐJ��ȓA�<���FQ�G�X�/Hb��ȓ��&���89����!E���l��S��3]��iP����^Y��Q �d�g�z	�h V�S�f�~D�� �!Z1 K"ޜ�Ktȁ:$��Ɇ�>��E�������dlm��/���4	�6T���!*�.전ȓ	�l���A�_�X�#�Ⱦp��Ԅ�u���ᶊ �	n]sM�2cu�i��S�.)��H�6�
�@��ޤ'��@���I�Q�xA `� iN����9@,�Z�FL�V"�*�k��tJpp��E�����Hٶ1nd�rd�T	�܆ȓvn�uTjµ'~��c�Q$r���ȓ9(D�����SDA��]����W�x���9������.`%���W�|� ���R�8�J��c(���7-�	�Pxrh�%�T5���G$`J]��O.�����<4�H~J��'g��� �1Y=��t�<Q@���JNƽE.�1,�.̻&�����$�S�	�l�j����9O�6& �L�ٰAB[j��E�0�>D�h��O�G���R&�,�
�)��@��`t,ίb��R�J��aL�`�'>�ʕ�ٹN�|*���	����+��ie�B�a���8�('�1���_�i��C�?F�@�B@��~2��b�R���N]��ű�����'��ɑ�K�	$�45v�)��t�Hݜ��鑵{K�(A"�"A�@�
v���4	!�D�l:�`��Y�C�� �n^JD�L�&C��e�c�(N�T�Om8�$>�sIh�ѐ6c���l�7j��&a����'4��cw	�IV����&n��J��T�t�l���A2缨1RFN(Bc^%s7�֘MB,�P��Z�sǮ<��h�)a��)�g�p\H�Γ.�����[�y����T����t����E4?�Yi��2-� �cj
<�x��1�ߑb��A��9#���{�.�V��@6<O�4P�nw0IT���/�@�"V�L�����VGSE4x�Ѳ�-f�� p�H	hx.9��-�D�2v���1%D�(k�P�+��@���c��YC�����̱$��! E�60$RP����5>��iU��%F�RMS�b����3�R��mDiյ7+LTؐl���O��MZ�iԷ3#�Ba�Y<r�k�M�W
�A�	�  �I�"Ĳ{��{v�*� z�ܺ#Q
��Jȹ��>9,}�Aa�'m��hpQ�Dxx�kp��X�f��\����<38U�O�*Q�	&0
�=��-T�*�
%b�m��S�@B#��N�Ze�r,� ּ
a�i�-0��5T��s4Ȁ�j�Rd��K"v�@1��LDu��u�a��m��*k�>�\� W�ul����k��d"`�׊u�V=9�Ú;�v��v
�&�j��h�%6�Q���G�n��DrЫW	s�V5���;�x���
��=y�Ѧゕ?I���B	
ir�4��$��:1DD6?~����ሏ&?
<b�Rf��8�L�a��H�#��#s Y�Ƙ���0R��H&?0c��S�e��ݸ3��IX"##46!��#E��C2���Gp㟜�",CrX*FeF�C�BVė;(��z$���)F.�1UI��d���i���C�e��05D��Nk���&JP�O8��1�M�VN������I�;�Hc��u���w���W�(�����6{�E;W��;�B=�Iè<�D�'u���'�!U�"���g(Xؚ�`^�n�`H(Ā�|�~�Y�į|����jF�e���'Ҿ	0wUW����%�#��u��M��w.�I8�K�R��k��MѸ��SY����%�?!��u����p���HG�Āg��@��㘡���f��OX�đBi��@7*�a�mY���P��G��
��b6E�(��M�w��yʁ�z,6qkġ$��@��'��8��Sv�Ԇˇ:�`���ʟ2$���x!l5<z:��y2,�5>6��j���RL��y�#GC��b��8
�9J͑1,"�v�S����k�f�� 1�Bj'���.�3}�n����fK2ߖ���A0�੡��|g� ����;]43`˟�o��Os��n~��C�Q=H�tb��T�jM���й>�� 	%b)�X�'|�`�t�Gt~.�0�l� �c��ȖI�bPg��
��X@0)����p��qu>�H0,��,��K�*v�Ћp	�-.c������0��<A���&b���4��281�r(	Ef�@�SS*X(���-*Q��� �ֈ�F9ł�A/��⒥بDj��ŞL���i�+�%S�tJ�h�,�I%�|Rƈ�)�}�D
�`��|�`ŉ'e��T���M���B.͢(HDps�G�+(4`��+��0��'D�6�x�I��"|�'��u�r�7/��;�i�$ղQ�.�L#��'�i��,��y�B�6.��+��h�.��w0� !���b2P�"2��r(j,K�!��f"�v���#�N��d��vM�7��yH`J�7S2�� �+O`�N=
S��� ��AK���r��t&��2��M ��[t̓_����P���hP4����"Z�G�σ)p��U)P�,v\�XpNV�:�H\H�m@?`�
�qv
Ŵt%�H���7� ��	@�d�^Tc��BLX�M�≓0ꍐ����b��P�'=�ty�WFB��:�=�Q��+K<1"��t	��Cd��a^^���C�ÏO�$5k���7i�ֵRf��s�z���Ѿ7PFa���ݪgRZ�3�\rH����C
��ŭY���!�ED�p�Pd��)^ߒ��ܑX{\�A��@��%�ټ��	�5���i)��5~ك�HA�tu�'\B��ץ�1*4�	�w��QK��q�`Q75HdI貃؀y�20���u};C$ׅ-;�9�'m�T@��g P�6MbA��C�r���t�܅r%�I��Jи.��G}�,��M�up�B�<����a�w�ݹC�ϮfQ��[t��pb�2=�����`�6i��U)��#���O.
hq�VU�7U�i@&� iv�)4MCo-1�H�
U�#-�#olP+Qh�.� �D��59ڐ�֡������N�Z�6�hw��C4��[aC�[L)����s���j�ɿ24��dĲC8@P�J��#Fd�@!�9�RsPda�z�.���*0N"l V
 �)Rt��rQ��1��C�3t� Ν�	\��S�퉒�p?i��oLT�Di�,k���*e�ޕ7vj����K�@Ţ�ܭTH�i㇇L:]�d���l���D�4sb̘�!�I�P�Y�%Ӣ&P�PS ��_���*@�3�Z85*�e�3���ja
S]4�Hצߘp�&�[���V�tdJqg�I���2��8!uNf9��E�6��E��yw1O�-Q����2�xŧ[8���O村`�ũ:ό��A�ءw�$Y�!��
qP��s�,K�)WnH�Wڥ9�L��.��	�"ѭ��[��ܘ6��ȸ����5%͚�<n1�4 blj	!�i�lT$�	�CV�I zt	�F2�����%��:`-�T���ad~%A3i�.k[:���V��Aa�3SH�ȓ��*l�bT��	�+
�+
� �=Xԁ��S�͛�Cʸ�PM�DXG��+���<I?����IU4M�5H��ٸP�ݳ��
9�Z]�dFh1��A�:)����␹n�`x������@B�O�G��AW^�]����I�5aS/	/=Č�G��9���q���:��p��e�a�4�P=z��>�IfL��Ff�*u�F��A��-V�U� �£��/]'N�h����X����ҩ?<�.�)4k��rhЬy�A U�2<y�����8�f�&����'(X������`��{aS�F��M�"e�[�ӡf�=e<q!$�?5�7C��*t�O�AP$Чw�����˗ j���
O�, b�̜4
�HZ���N�DC7�	$E"��s��'`@, �4�U�p�Xz­>	rA��p���Kp䲟���噦�0��_r8*��/O�s��â45bQ�A���8jhA��]�B��k�P�,\D�H�eѣ)��Qt!j�`��%�]1�Rɜ%@ў��%�@0t�X��v T�b'&}B� �9 ����V��1`V�щ3� и��O����� "�Bt!����z��=�rm#&bbmR��`�R���'c��"���#�X�Bਕ�j)(����+w���ib.T+ �H]�ƢûmbĐ_�� Q�*T�E��Qc����0bJ��g���NGF� Q!�%f(|y�kL��p>��mT.0��U���ȫR�\����N(Z��KG��4<ˀ�j�Ȕ-����	��u��pӓ�ȪW�N����^��9��
�>τ��;2wN�Pf88���Ǧ��D\*�Fy���/0rD�+ ��8:���HG��)GZ$�b���>*x��%�
��t��=*��CBƬNV�1�`o�
G������:-t��4%[���P��H~2U4
�8���S� p��ٙC�TI��*@��2����B&;���	d��5��!�	$t�3+Y�G�Di��-!.D�i2f�=p� �ks@�HԖmqR՞"d��3g�R�5\��T��4v-h�8��×5Z�q+���@bXK�"A�$HA�E�7�E�С6��/(n<2d�
�/Բ��'�<��+��U�m�Z��viKk��KQ)���P���%,Or;�BR���rp-S������#�]4��!�Y~�,y�J;��8��	�HX�������dc�P(���k�\v�8a�H�e.@��(F�F����N���D⟌iB���0�J�(!Q�z��"��]�%&�� c,D�	���J6I���T���^�:A��Po��c�r�kqn�5)��Eٳ�͒���b	;� t�2n<J���l�-�fߍ1�vZP�U�6E�FY o���@3O� �ΰi��� d���4i����؛3��E����3n�m� �Rk��m�iՒg
�ܡ&+�	�6Aئ��W�L)&���k����õg�I~,�{�BU�C/d�"��9X|n��B?t(\���G�U
8����FOs(�S�╫C(n�" ¸[vz@j���Ԗ�c�eP��V��Q!��}f|�Ǔ@�(l!Gr���фJ�9�L�{'�ʆq� �p��aE���C��p-���FL�ʐ��_sV�*�D
��1(��+
Ād��'��Y�[C̉�9д�PFY�@��O�$tH`�z=Hِ j�9��G�p59ƋW:PD�HRQ��H�y���6d�ud�N>��!J�����R�@W9UL�\Jq�B�@�I�	ά��D�-)����&��y��	тf��ɪ���*`h��w�ؓ+d`��Q(ڮ,��)m�,Z�v9�����`�M֕s�d�Q���Y�v-H0k�"(�R\P�@K��a��O�  ���BɅG�"?�����¤J��U�m=X,��#ߘ\�&%�h��T~X���ő84콭�O@d<*C�T�Td��h��Ϗyfxݲ�DF�8̴a�C� 9gNb��E��&Ij��;,O�Ț��-,A��@��X @��4���ɣ<%�F�~�s��^�@� DgE 9b���� �@��59�!��CrV��J�z�[Ĩޒhd�l�B$��N%֢��~�V�?y�/T�f�ܰ� �	�4�"���R�p��͛	)��eE 
��u2�	����Ţ�1^[8���qE(�� ���
�f�(�
UPt�ӹ �NL�'�~�'��1}o��z������.n��S`��2ln�E��<z�lq4�:���+�Z����g��B�����c�o���
5�_>ܩ;BK�/5bЙ&�X�T����ɺ#���R�v��"@�tEl�<R4�+��͓\�I�7	\�e���R8vt���K4{��1�A�=S��\�5Lp�&�@���4y*`�m��(�95EۂH�JHk)O� F��o(y3I?7͂�PR�!��-���)�޽:��)��$-JJ�(#�"kl�?����',HD�A\!jm���ɱ/�fm�U5�����/^Q�'C�SnH85i�=kB����ѕ{3�{Д���")�nRj�>��7�+Z�"�a"�U-#�Z �UA��z�↪ʚ%T�BrjE��y�ϗ+m���	��T�$�@,�աA�x�ɐ���&'O
��Z �R!zA�i>���Ԅ�b��E�P`�+@%~La"�Y�ID� P��޷
��R���� �ڊ��d� -,[�8�Aۏ"����a�J�
����Ek�#��D��t� ,�i؅HR�X0tc/B,%�'J�L��}��叆F;r�zD��y�����|:d�/A+5�W���L���x̠�Q���W�t�[���^٩�,�O�}R%OƼ �&���?#<�DK0�:�z�DV7]2N�2���!L�Z ۑ�R/rAtQ��CE��0$�k�1��Vn�k�v���`�D�~�H6`�2sl��^�m�r���?8Lz�'p:Q��6�W�TL��c��3�8̈1A��tѤL2UH�Q���cH�L�t�P>3�p�AG@�>8�p��O��CJ�O�QؑWv���k'�ո���)D/B^��OٓP'��_R�%jf�T�DL���=	r|��%"M�@,U!�2"�������m"���� U�#�J���4������?A�a�0&�������d ��n���0q�eb��hF��`H�Cd�;7��=�6����b�Q���2t�I2��jB�
uR���	�
H���[�`we���o��m��U	-FxB�#����-,������Q�9��%ʡ
�xǸ�2�x }���^����'l�-���ؗ�9���ao��m�� �,P�W>�萗��/���
�F�C��x�c�&o��C#��>��qˍ��X(0w�X|  @�B����k�Nw�����AF��:�O�Z(P���,H��(����%��6�hHr0S�zV�y2�ٷ�xl"�B�~Q�pТ)@RX�@C`�@V8�A[pHU��3�ā!�ł|<��5O�%(� EP0$>M�$�� ?L�6�C�fj���:�ă,d
z��0�L�z�JPC�-l� �
v���A�\w�,1�Ă�>@�b�S��ޙ�����R��$I���䉁��	���	dT�\(�l\�P�V�r�ة��Y�e�G�֙I�	Ԭ,��J���gQ�T ,�^� ��eY�A)� �:Si
jEHekF�$i�F+!2�R���I%7q�+FL	�I)������>�j`1�':dΆ@�T�.|���c�4r�o��+�N0˝'-���҆ p`j���V���5iE�tLn�
ϓW����	rAx�KrF��4X 0��;AD��Tn<��-qE��L�k�D�O��h�)	���\� �P`"/��d�* �d�R�=�A)�'Q�%��'<�U2� �P��!�L:�Q#!}�H�=� ��agT�*��G#�de2����'wB��@�{>t&�S�^�axh�!e��5��->��T�Ȧl��@�Ɖ�S&0��#�_�1�l�&(�C���?"l<(�$MQ8J�ы�(�{2�j�:_A�Ը�Y<	�!��UXLYb1'�� �� �����.���Q�e�'{�Y3��Ͳ=>&��b��QSXUr1�ߴ���,���q�%�/xm�Z�����y���az���n��`�,��
z�s�T�n ����Y>mWnT:���ZqBe���+��͓E���?�%��7o�����'�P��*J�TK`$��2j.X��{�A�5����*'QPh�J"c�q��O��1���Q�>��H��◢�hUK�Z	�#/�7\!hz1/���0<Yq�܀LC�q3��2&=`��p�ޑ���䚷��I���dOp�@C���$ ��[P�Z\H���ƨ�p=�F��m=�M���%��ч���HHlPŅUV4Ќ�sj}�����D�U]�$M�8��͙'�J�LBpx��5�S�?�ԙv#]�{&���^rC�I'&u��Z`b�=FJ�����=��}z'��.��#�$�~��s�L!H���n�Q���%��P��i3D��:LX�m��.�lH�Ao��[D��	�l���*F�t�U�'�HYks��wG^� %�?x5Z������@�
[�P��8����>;-R8� 
 !��)8��3ސx��\"��:+ҏH� ���V-�HOh1aGNQ�qC ���$ G�D�N�q�8C묈�����yjH�'�4�����4f�����y2h�=����=E�$CQZ>�I�lF90]��r��X�y�Y�md��k�9�v�H 
ԥ�y�aϨr��=�ᢓ�.�F�{@���y�O�Hh�I@�!	&�����V�y2l�9=&��c↋d�0i�wn��yR�K�8]�7�đ,˖U�g��yb�5T:���B�՛�<��bU�y"�� ,}�,�Gd*O
��j��y�mI�%�&i��OJ��1�v�ŀ�y��=h�=�FO/s�ز����y�GP%=�
����:B4�F���y��p����d(K8���1'�.�y��WYɺ���+3	4�JV�ʋ�yR]2l�]X6F�3��  % \��yRl��C��`8�k��R�����.�y2�l@u��l]~�Ks���yB��2�����B<vyZP�W$�y�B   	���9j��A�HҞ�yr�9��9�t�O�5�\���kQ�y�ؤW�� {V�� 3�:`���y�Z�s����K�r��)�r	���p>IW��1�<�f�2�4��4J���Z�lE�F��=Y����L��J1��릩J����~b�њV�i�!i�v�P� �� ~F�ae �Ʀ�Ǯ]����S�o���p��#o���a^� ��!�f�io�Ep���>rH;�.�:â��ޥ��mSJ8�!B�B)3-�e�O��Z�IMѦ�&���nY
��4j�Q��.Q��Y���>�T�Y�\��v�|���E��a���bŢ[(_�$uC�mP��~B�V��@7m2�ԟ@�>a��;I��b�,�6`J�U�V�`�Ű�����S�O"�u���1�|�%+Q�Y[�*0b�NO�"ç*Zq1��e����L�%߄أ2P���w(ֲq�2xr�O��}�&愐EN긂'ߏQ��� �'&�(zB�U�8�|���]��>��o��i��s�/�
m��J��j�FθG�@ͨ���:0�������0|* c�R�p�����3T�J��33�)'�ă��ȟ�x�
�%,���UgE/)ХVm$�bO4�C����0|��핷D��$شo�o���tCb~�I��@�&,���DF��+d�|�a�o�? �*'�d��扙f����Q(r3Q�b>I"P�Q����
�MO�{�T�kU�O�� ��O��OQ?�9� &YNX�;'e	�>O�ZU�M3"��%��-�L5���X<6�4�k�bT�7��H?O��kl3�>�� ���1Jݙ
��@&a��.�t���l��֓Ov����O�`�`�̸j�y A�h��4㤑|a�h��0�çaU�M��!Cr�-�&n�	̤�'�>!Z`m�<3ɧR����	�R̵�v��19d���ɐ�yr��l�\��|J?�J�!�0�Dĳk"�9����X�@P� e�\F8�6B�3H˨u�e+D�S���O<�F��07ْK��9���P�c��n��{�	0���]�ոOo�}��|b����Y�8q*Qh	 2�&\�6���S'�����	(i���
�Oܛt��	^ 1�C�I1`��}26 ��.�����k��f��B�I'P�a ����A�X,<C�	,*B(Z�u^�c@�2a� B䉠 �d�fO��i�H��vnЍ �C�ɀy 	��//jDIr��--�C�	;#r�2�j�3L�f�"�LJ�B�I����{��X�=N�r��ˁC<B䉒U|4� B�"d��U�T"B�	:/>�4��`�6N�T@$I�A�2B�ɐpZX|����"�����e�B�	�$���-
�ȵJ�	��9#0C�ɠ(�b ���jm���ԋ�6h���D�#� �X'�X&6�"MK�o��H�!�Ie?�e�5�?j�\u�Pm֘Oa!�d�I���IKth1��ϫ`B!��{���dMT�I@�XaR,��k?!�[�p�)�"��8���ʐu�!��[���r ���0�6��/E�!�D��Ve���`H(T���A��ix!򤅰P�^@�Λ#+�����@�3!�$�5"�%�A�]�v�Z���g!�d�0�,��LҼ}u��x։�%!�dG�	���7C+vĘ�JF��!��8�ա�邝[����(��!�>V��l�� �0ѲG�V�!�\�c��PD�k�@$qѠE�\�!�d0��5j�IP%����4m�!򤀎B�Rc��$���7�1-!�$Z-'4�!�@��$R^a���
�0�!�DO�tr mFJ���0m!���.j(�-�P�2(M�$�݄q]!��A*a��R�FˈU�D(�D�S!���J-V��!��/|�f퐂�I�k�!�dV����oM�C���3*B�,�!��s��C��F8SD�ڔ��;�!�ę�hR�4*BO��b�*����2m�!򤕴}Rem�+}nM�B`�!�ā|��!��nB'[�������!�d��)äYŋ�9��	
�i8G|!�X| �Wо=(Uҳ��Y�!�$�m�%sck�"-!��NI�!򤚿.�t�rO�2%����[�A�!��ߠ/��<:��݄>�|��n t�!�Ė�It���r�؆r�0uX'-��!��L�t��Q�ً_�DQfK�g�!�$L�B�*�O��%����T
K�/�!�$E���`p�� ��&j6�!�dH%mN�E'��U�]I$��?�!��ʀU�⁚F��P�xI�b�!(�!��^�+��I�O��;�ޅRa�!�T�k�(2- �#7�\���W�!�D��=�H�B�DЩ
�f�3��s>!򤍎3���S�O��r�A�˥J�!�V"�Ik3���&�����
�C�!�Df����7�����Ռu+X9��'�䜒���ag `r��F�?jB�*��� �U�����<��c�ˀ.,���B"O0��$Dz�<eZ��%i��ٱ"OX�� �N_�"��A�'d`�;@"O�\R��l��XBq�W�2��"Oʜ@EYc��58�b)&(�%�"O@ ���B�]�B�y㯞�r�8 K�"Opcp��Iښp[u�3�4h�"O Y!�ުJ�X��.s�Z;�"OРb#��`2XHbqn�,� ��"O$���M9X�4�H'#G$I�e"O�����=h�`��/8"��"O���g'��NnJt K��M#4�9�"OM�D�*-r�y&k��JFh˕"O��b�3r�}�3��g����f"O� �%�7T[�mj �p�VՐD"O���f"$؅)Ɇ^P��"O�z�E]:&(��@'DNj1"OzDa�h�?�"�k�.G�s�-v"O�t��B�,�^T�s�%}�|�E"O�A����"+��������"O��z���4?��̐���8��([�"O,�!V\6��e(�Ѭ�Aq"O44
�2J�E�gI�)� �
�"O����O�F�4y�w	��~���{2"O>���ӎz�0� �'�^uX��R"O��CD		mΘ)ʠF^�g�-��"O@a��H��\e~8a�Ӝ[\����"O��@"�§�6 ��W��P�"O@@#���)̎ٹ�M+U.��P"O�p󲁊�A�`)QrK;3R8(�"O�؃�J��YhhD��D!0���'"O�\��^�׮��ڞsv��"OHɲ�DT�!+b`[u�]7$I��Y�"O�,K�q�Eab�>YҾ�#*O�ݰ���0v�@h�`�4?4m�
�'����]��J� Y�#�5;�'����`�*.D$A� �ר)j	�'��\Ƞ-��Hv޼��@T.�f�#�'��1 ��PFd���5b��A�'�Fi��"��"@�^�&=��'��:`��e|T�1KFT����'�nX��nD&��m�Щ��w]-s�'�D����#��+Pk�	hg4 �'�ޑ�o�>��aQW�bۖu�'}�����)�6�(����p��;�'��kE$�3 �Ԝ��ʾT�:�
�'r>\�J�6�����n�L[����'��M��&��b�Jd�E�ǆ>����'���SE�&�R�;5��<��%��'}̑�w��i��Xq܌2�pi��'���	3銔kѦ�9�������'��!����dդ�
#���rϨĪ�'9�	�F�!�X�g�x��\��'1>�z��ϛ�&�f�Ѥ}Ό��'tdPxөж2���ӣ`�!r�<���'�.uJ���:�P//8�f���'\����C�jo��G�5?��b�'�@��7�I8+b,�)�?-���
�'�����M=sL��+�5/<�Q
�'mDq�"�E�Ci.�����@(���	�'zj�Ѯ�0~�aJ[�0�Ԝ��'��i�,���0oE#���'���3iKA�h����E/����'��	*&�(e�Rxx�Ȓ?_����� ��y�
}��L��,	(n�p�"O �&�Ğ[(��
@ ZB�	�S"O�(ZfAԩ�J����o�R��F"O�9V���*' 4Y"i�p�����"O"���2���x�"E��c�"O�E��k�)�6E)�f
}�Dx#""O  �u
�e� �H!��(Y�z��&"O�t;a@�35�U��FQ�&e�I+�"O��)d�чA &��&�n?.%CB"O�l ���Y�d�Q�ˁ1/
1"O��ǨĲ�4!��{2٣"On��LKb�e�G�
`x���"O�� 88|xr�=%LM�r"O2�P���W\�a�0�"8F҅!�"Oa)% C�vzA{Eʔ9*XR"O�����E-s�n,�b�H(��CW"O~D�4$R
4$X�$&�q�"O�yA?���% �G)<M�"Ok�jߚ[I�������L�W"O�L��n���6��5���"O����"��D����q���`"Oq��b�_�0��aL�O�Ƽ0�"Opp{�964�������hH�"O:�S,�G~T[2FE#\:N�h�"O�l��O�=28])�e�@7����"O��[&/^��Rj��v0��"O�Ԑ��ιL�����Ƌr=b�"O@IZ���+��H3%�ݴ5醴� "O���#�@�2F&ƾl��1�"O�lr�F�0d����V��6d6܉"O�88�lS)�N4�e��UV�  "O�x�4oT@��SBK�{$h=�"O|lj�-Cv��17�4>�!"O
�GděGnLӠj�[Z(�"On�Y�iߥP��l��� LZЁ�c"O�q�e�J���	if��
vN���E"OM9�
۫QP��_�[5.�"2"ObQ�N�ru(�䃎\(z�"O��Ň2a�j�cV#E L���"O�q�åE�yJ��8Q��:~`@9V"O�����U5hl=�èŲ!BF���"Ovb����7	�8N�]Ku"OйHߜL�X�(��|I�  "O>%��$2��RE�<mR
x��"OP`a�N	*[2�Lc�E�}�%��"Ot�`
��E�F�X�Lq���"O@�`�Hi��Q���iE8�1q"OR�`a$�~w�Qy0��<*���"Om��܌0�Q��h�*kZ]��"O��  �ߵ)���'Ɖ3Jf"OzI6.ǰb�!{6*�;#�$yA"O*S�H��,Z!JI-FXma�"O�x�&GD��p��._����"O�EЦd�P��As#�Ρ�"Ob-�+ �t<ȐE�� �"OzX�#�Q=:�*�b��T��l�"O����\ d��8V�Ag��H�"O�D�BN�lZ���t��]�^-j�"O�a�N�)1r<0�ˏ�\]~��t"OR�X�F*�E�g�	�qMzب�"O�� w*��)�v�i ��F����"ON)��S(e��	3�kF�
<>ɤ"O���4�
�u#\��k��5:�p�"O�����$�Q�Tk��%h�Z�"O� �e9A$��IdH��c'G0M�@(%"O�l�c�8#�.L�&�%��`��"O�H�� �h\ B#�a�2���"O���HD��,`��\�4���D"O�����-"��b��ۆ!��)Xe"O�􃦈I�x�)�$@^H�̂d"O��:A%�1٤�4�ťX~Niig"O2�����&$Ȑ�"��`���v"O����'�RE���T�2I�XB�"O��r�ŗ�s����`.\�~-ʌY"O� �7i\%{��(���8
,s%�'���G�j�|*0e�F	JY��͔8I-q�4B��͇���0z�O�y%L���F�� _��r�Z(`�r�@6,$�X��&���f�+�֢<ɓN@-<l�A�R��%���*C�� n�\����x��7��A�/�P����b�KhӲe�gD�%W>�	�AԨCvU��![��M˰�x"�'�R��O�<�;�G�*nV`�U *F����[%q�?��f��w1��8�(�e���S��3}��r��oZIy�F�8�<7��O��2�Q�\�[� �c�� N��`Fy��'�4](ƎP9{v6m�{��!ӭ�2���ޞ"*�#UGG�)�jE��M�j1Q�H�ՅҖ|�VeO*�����,X� �C�J�?���
&�J*(���8��i���@E�Ol�n��M����u,�9�"����N�p��$�%�~2�'E�	my��	�U8��`��T�T�F�B�M�aB�i�FA(CD�^q�ic��Z�Q�� �%�Ƹ2���0k���4�?iJ~������@N�"�eI*1<��(&^>����?z~0/[��!Щ��cq0�sU��3H�-�R�?��@���5*�b����	�c�+Lw��=!2&�3o������BƏ�p�Zk�@���O6I	$�Y��!�d��L�B���η>��GП,��4u�|�Oȱ�ڑhF��&t�m��[�b��>!���=�h�6ze�����FZ�@ɳ���'u�7����'�خ�WQ�<���ÔTWf!Q@�ۉT�{U�'rr�'�����&Q]��'7"�'N�ϻEex ���S�/D>)���7���xW�J4h��Z�bW#$?ҍ�Rj��"��!Y�\yR��0	��2a�Ș��!r�Ö=�iЦɴ!�@��PI0^0 @I|�aǜ pgr���'D-�V��9`X�j��I:0 NsA��FyBꍆ�?�%�%��'>��'����A�E�<��4O�<UM���'Oў���d�r�
��ts���_�����OBo���M�K>��'��)O������V�4t��.�8QHhի�kZ;L�o�Ex�����8ٜ(+��1#���!蓴�����L�=�{�,Q/���j�)Q
|d�����$ʓ)��R�K��%� ��fb©OܮE�c�l(��iы\�Y�8�'�-T 6�)�oO�QmZl��I�Ή�8�.�bbAƕ-���@s�i�h#=i��$������.`0и��PQ�<���?)I��V�ld�w.ԅb��qS(}� �`�n�y�F��T�7M�O@�$s���;�����6J��(����������,�����ٟ(��<bѐ1�,@�[�0 0�o���%D:h�`<��K+�:0���K$�����)*0Q���q�00�Ґ��'{R2�9�.�!8HhI��ՇRv�Ѷ�?(p=)ХF��#<q�Ȑ֟ ڴBG���'C�Ά9+��;a�!J���2&���'���d�O��$�O��K3Q;ը���Ԃ��b�:�����MU��Efؐ����9)LI:gůO1f`�H>ag�/�?�L>�M<�� "  ��   +    u     D+  ]7  |B  nM  �W  v`  Ml  Bw  �}  ��  B�  ��  ʖ  �  L�  ��  ү  �  U�  ��  ��  �  ^�  ��  ��  n�  ��  ��  � � 5" �0 :: A CG �M �N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�'&�IK�)ʧ�X��)N�T��mkq�����u�ȓ1tu���W�7r�u��084�1��3��y��i$[:T�8��OH�F�����)yF.dJ�,� I(e�d"ٞ;>�b*^L�'Nў�'~B�����Ɗ�VT�^'/���	j��X�գ7N����# �zi.��p�z����I�T�<y�%Y�0cȩy�f��:�a������ODt����k��B4������!D٠g����ȓx�D����B�l����!�*M���ɩ����d�)�$��6F�0�3І!j[�@��p>�H<1�7BӒH''F�'�,!X$e�zyr��M��(�8�CǍW��J�[�YV8 ��"O�  a9�L�;U��Ǭ�%}A���;O����=I�P:P*�:r�c�fX15"W�o�L~��K��X2� N}\�J��֤�y���dzjysUeр?��õHN1\�J�"�i>}G{���c��Uh���v�����yB%E88���0b�**QrăUD�-�~b	4�Op<�o�N��,����zw�����'��I��, �DZz���N�Hf C�ɽ;�,1YQ$�(K�P�r�l��2B�I4"�l G�0�nU�(�1&�C��
C˒��Ѐ�:$I�MP�	āH�tC�I3G>&遳�L:wJn1���^4�C��v�X��ؔ<e8��D;2���y���8�	�$˲�M�F�㴈�d��ȓmz��cZ�"��L�a�S>���gd��ɦ��7��B$�r��e"O�9�����Pp�l��,�=��"Ob�K#Fe~�AI�%�d���"O�p��eܾ���H��[�@��"O����	�jP+$��|AEq�R��F{��	e�� G�=c�d���C�_M��$v��k�j�(�^�H�HQ!=TL��"O��c�A a�d� �Hk-����'"��	2���mL�]쨁�D�
�C�I�h�p����D4zr� �:��"?A��S�:+x����$��TсmY$XB�;5D����nP�#t(�.K�
�ɝe Q��}"���\HYW�U/8�,����a�<��I&1eʴ���$N�,��f�G�<a�Ι�Q���&��0�A��DX����S���Gn�
�D����֧Q�%���=D���'��@��-�.֔11ғ�M�G(�'D�9�Cn��pfB����43��B�I3
T����ճY�&9 1��g\vB�ɋ>F@��A֯kd^��P哟FN!�d�")P�HD�a��iE	*L!��U򐫴�#M���cS�U�Iꦑ�=ً�i�x�@s�ȋ)�Z��"��0�!�Ć�)�Сɳ�?�e�r�:5�l$$�l��O1��'�kpm����+�J��-v�
�'�� �&��	G���x�D�l5@��	�'<~���%�3�H@��#�u��
�'�.Ԙ�6G�`�,��m�'���(E��-��I�d�d��-Z�'@��hB�E,q�hETLʥQ}�Y�
�'?�)PL�g^�����J�赘�O�tb���C�2h�6�u�ԝ��'�� p�J"��h���?��UYT�&D�@R�]�^v�t�F*�=W�ȡf #��"�S�'O�e�%[�?�,���^�]�@Y��KFT�s��1,�¸�`b8%����';�I��(O�K�\�8C$���^�S.N%f�t���;�O>Е'B�X��
��R��X�D�Y���d�O�h�vg�5$~��t����R��dG$s�Q?93�n�y����G���D�J5�n�G{�����S�<��cA�*^=ZB}�剤�HOQ>��G%βy����f�o�Ѣ *D��p���$<�9�/��-���!Q�%\�'��)�3�� �t钰���9d�rLڡd�!\!��*���$�� Ig~�:E�χ&�h���)j_��v�V�.��%�Ǒ	8l�ȓ)����4(ȥ �J����(
�nh��E;�S��?գK�F5�a8&h_6]͎��L�y�<q4�ӠX��e�FW�`���sFb�r�<� �d��(ߕ��Ҳ��'�$���
O~6�ӽTCF!Q���g�<�:GER���:�\D@'nc��xA�͜Ͱ<���ą���A"fݞN�@�Z7�O0��|��x���!<�lI@�b!��(���<�HO>�iϯIf��kT),� �+��'���Eyb-O0<��l#��ɷ^#ΰ�u�� �y�.?�p{�O4j�:�YuK���M���s�f�cd��>:dP�lR6�� �"O�᳓FC.u��h�%����(�"O6(�t�N�y:�� �]��h+d"Obp
R,�`�����S���+�"Oj\3��#I��6F����Ӟ&�!�dS'`<� ����$Ġ*�E�!�D�7>�����k �-x6b�0�!�d��i��(8�b" D�} "�ղd�!�DOVY�QQ�e�)0Če+d'RC�=�O��c�,�M�&`D��Ŕ;\����-'D�ԡ$��-mb͚���--ܮ@Qe�%D���UI��������6늠:��#�OЙ�'t0��WL7=] �P	�(CO؄��'��$���N�9���@���8r��B�'���8�ղC�1� &��,�0
�'o��������3�!�)��t{�'j:"=E�t��!�`X�T�Y�yƄ�A��y�W>[�|M*�R�ɞ�!��#�� �OR��fA�m�<���9zuhQ��'H�'Ӵ��[/'t)�
�",	��
�'��d�D�б����&BU�/(��C
�'����L��,�	\�=p�	�'�،�ѤK>7�
���$6�v���'"ޜ1�.K�nZ("� �)�L��'���SF�N�$���;4@;v��	�'�dqᅈ�!"����V+e��}q�'�ȈG�J�,;8��6(b&@\�'d@��'�.Wx
�X6Ëh�$�
�'OX0xgŉ�����Y�r��M�',�S'-�J�&��CGC�gz����'ؖX�횙=�a2�U^��u	�'a��	�1ctT�R��T��a�',E�-`�Lٛ ң�|z
�':��H�L�������`��'��pɅ�'S~X;�C��x�'o�, �A��f@���(A$k_ڄq	�'���3��ވI��t�T^T��Y
�'˶�[#���r}82S%��,��'Lx�
ޏ ���������@9��'���W�̉$/��I��?z�ܥQ�'��*��-�0Tp3��(w����'��A2�ӄ[�n�Q��[�iH��A�'3D��A-M;������ j1t�'��XH"˂>A���q䂏���	�'(�Uj�J�*Ϻ0�AI (pu��'�bh�V�K��RR��.�H� 	�'����g�G�O
�h���651	�'�"8+S�L�!����0�T���A��'�#�C��|����uR> �d
�';`j�C�7k>ʀ���"$}ȉI�'ٰ����S&t{B�ٶ�_V�\A�'SL(c��P>�&r������'>���r >{��-!���lol��'H���� 9�0S�N��Q=`��'q�A��	$b� X0�@�;y�Q��'_�}� m�f��xY�͐�}�Ld��� ��ց�8~L���Z�&~�HJq"O��b׌S��\ �A�ϷAF0��"OրSP�_�O���v�ڋ1a
�"O��#M3h7���v#\6�A�"O�gm8D�8r���"�.�
�'�B�' ��'���'}��'���'��-r%G�?:�� c��ǯ$�����'w��'!�'>�'�"�'���'$���#�K�Q1
)6�BF������'N��'���'z��'6��'�2�'s���&�<���ڶ�"���b�'���'�2�'�2�'7��'���'&�eig�A�1V�iÕƏm�L����'���'a�'u��'yb�'���'�x��QeQB���b�Ϸ3����'^�'92�':B�'	B�'���'_�aTB�ZDLXk��H�{�Z0 ��'$b�'�B�'��'M��'�B�'�lX���v ��	�BF��#�'B�'I��'�'��'�b�'���qҡ(#�]�ơ3E�(��F�'�'��'��'"�'���'@��#����I�׋S>[�h\���'��'�2�'���'�b�'�r�'1䩠��i|�h�j6:F��$�'�"�'c��'�B�'���'���'ߔ�%A8_*�s�A�	]����'N"�'R�'���'I��'�R�'@*e`B$:^��q#��c�9��';2�'�b�':��'��'q�F���O�E��A@+;	A�/A1�e��Dy2�'0�)�3?�´i�йx��Fm��`2�Ps��Ś��������?�g?IߴV������B�f/>ɰ�԰\��j��if��7N�F���Yd��&txC�~��T-fT*�Xp�F
v��:���~̓�?1)O��}B��
�}���§k@�d,ʈ�A"�//����٘'i񟀈mz��:�c�+x)Ll�K�H/�ճ�K�/�?��4�y2Y���J���u��扏E�fܪU�Ӷ�D�,1t�`9OXժ��Q�Hw~��a7��|��=��<���3�|�d���d.�D�Ŧ1 go-�O��Ceۉ1ʰ��I��,m���?i�Q����ئ�ϓ���X,G|4z���zEh!	��D8p?��7B%�����zy���I�>t�����?�M'g�2|Ҥcْ8w�������d�<��S��y��I jO��rt��j�0I�"�y�@a���q���Sش����$��;L��9i�.R� QW}��'r���'(RC��i_�	�ѸPi�%��0�����Z���B�l �L�#�G�Y���V��$?�V@�>.0p�N�5o�$�'?�R�i��tH�y��O��O�bm���L�B�,�T�,H�a�<1���M��'��Oi���'�Hei���F�͠�O�>=�dmeP8872uX�O���&KI��Ε�YwK��'K�y�Fa��U"��\I���1��Փ�����<�O>q��i���'K^��T́1�֭����(�؜��'��6��O��O��O���mӼ��^b���(Q8�HI�N�[��0� pӎ�	⟠�V�K�)�n`U0?��'Uk쇹z�n��"�,x��U7�	8����O0ʓ���ӬP�:���D,�Z����T�M�qOl m�M�4�ar�v�'��ɇmp��@a�,6q�郶�1�)���$z� �mZ��@�%�����?!�Էy�@���u�BC��l9~A1��T8b���P��4��ʓ�?9chGt|�9C@c�	18������<IO>��iW%Y�yY>�f�I!a�����)V|���0?Y�S�����A���'�*@d�b�`���3+6:͠�lBD�<�u�+a��$�'���Q�B�$���#p�)`G�?�����dQ,p�P;���AH�A|~��,D:�V8�M��$�aZ:\��t��芜�P��	G�}>X��)Dd��+�.�?Vؔ��" B"o�*��*[�$���E�
�"pBƫ�t���k��A:^μ��B��#o�t 8d"Ӧ9v���A�RQ|��5� �YZ��2�B�)6D��D�R�$���'ذW�t�S�L�f9� I���e��M)S��L���CQ%4�D3_���`�`����S :�|x��j��l�=��%`\��cP�H)G�:��b�����R���&�@;�� >���cI<����?����D�Op�dM�?B�9w�Kz��7#C����f:�D�O����O��&L���5V!��6�m�JC,e�4�C���O����O�ʓ�?���G2(��O&��r)W�+}�Ցq�_�1$����OP�$�O��Ŀ<�U�N1�O�8�e����c��X�EMTp
��p�N���O��?1�\HT�|"e�>�����\�,�«(g�F�'��S�8)�����'�?���OE �,x����2\eLI(dQ����'Gr�'ҍ�T�'���4:���IT$w0[%P�EܰlByB��� #�7�K�d�'`��,;?��C\t)����G�o֢9kuf�æ����|�W�tyʟ��x�y����	ĝ9�� W
:�M	[�W��V�'<��'7�td<�4���C��P�|�^�@��A�XS�������Ky��'�b�Ϙ'���ְ`���e�B2>*��k@ �t
7��O��$�Oꀉ���a�i>������ 2�gB�ȫbF��v�<�XWŜ*��d�O`����1O0���O��$�3Z�f��EI�3,d�K�bQH9l��!������|���?�*Od�AT�À%2e�f��q<%)&#Eʦ}�	f�b����Ο��'(���a��5�&>&�RHiw G�K����Z���	��T�Il��?iG� �S4�Z����+M<#N|��"O�:�PH�'>��'c�	ߟ��S�f�� aq�d�ɘ-Q眠���
̦���ڟ���W��?A��U�>xo�'?���@�]�0U@E �GW�B�\��?9������O �z��|
��|�:��uDI�\5D����2$Lcr�i���d�O:�+��|,�'+�\K�IU�Q� �c1�eW(u��4�?y/OB���-`��'�?���:�B�0 7"�{�Λ�J���ơ�9R	�O����f�~!s�T?y1��A�T��u�Q�Ӳq:}Q硠>���7ò����?��?��'���6�&��`��0�i�Z�\<	�T����v�0(�6�)�S)��`RQ*�_�f��ҧ��Mm,7mE;(���O���O����<�'�?1t�F@�y�R67'���-Q����B]�[�T];�y��i�OT11�9~�}��Oí�T�#�!U���	��t��/^�������'���O����aԴ{0�M�$J�\���U@̓�*}qV����'i�OnT�)"�,Wy����ד%���'�>��[��I�T��k�5�����D�����D�� :�i�'����J�����OF���<9���|m���+<�"��L���RW��2���Oz�d�O��(�	�kE�h��̓�j� �Uc�`:��{�NDd1���?�����$�O�yBo�?%�%��ZqD���1�$�gaӖ���O`�D:�I̟8�G,V�{v�6M�#�d�XSA]&I��}bc��jd�Iџ���Ryr�����h�|���"��se��}-�L�THݯ7Sr xu�i����O�,
0,��
@�'~ �j�)�� �D��k�>�xߴ�?,O��,6�P˧���r�����.r��)o���!�('�O$��Ƙ&{T�z�T?Q�gN/�����Bþ.�d�w��>���zE�1����?���?	�����)z�P�%�FA5�)Q�V���I4\��Q��6�)���X��I�"|�h���C:�6���QL���O���O2��<ͧ�?�gO��*�	�d��5��͡�V�f[�V* #f+�y��i�O�b�'o@�mR�uV�D�Ԧ��	��T�	Т����$�'2�O�)��P�2��t{�	�Xn��IF}̓i��e���'���O�au*�Z�鷇N���]�T����k{yb�'���'�qOЃ4�^R|��UiWE���h�S�$� d�5Dl��?	�����O(C�ñ��͸"a�*t�& @]P��?���?��'�����!��W�b�q� x�&T��B\%r�<Ń�O���O���?�KQ��Ĩ�&�@�����(�]�7N�!�M���?i����'��	�Es�7	� � �jqe�4z
�DE�S:_i�	��8�Igy�'ѮV_>��g�r���`��@$C�0�xm֟��?�*O�Ӝx.�*r�i�fŔ�,ހ(5�D��M�������O�kA�|��?���=T��Xv�(8v�����邬*A���O�C'��_1O�S�z�8��3�ñ:���(��M6���?�bK��?	��?Q��b*O�֒|ؠ}ň�)�(��B�%���蟘1D▨U#�b�b?	e�.z�J�9���0N7�����v�z9IU.�O����O��$� ��|b�x�qS� �&'2��N͠��A�i�,aq&��Ϙ����D��i�B�l��	S/�,Q
�n������Tȣey�O�B�'��$īb!ѱK � P$�E'z�A�<y��X��O/2�'���H�#��]���O�����F$F��'�>���Q���џt��Cܓx��3�ꏀ.���v�a�'{�Hf��7����O����<���G@�D����*�����ŐGb�Ѱu ����O���O`�X��3<��3ej7C-j,�g�F,Y �
�)�,Y8��?q���D�O��!�?�@C(�"@S@���홶,����{����Op� �I��4�D��.7��''L�M�Rƚ�� H�,�������Wy��'~���SZ>A�I�����eޕ(a V)�:<���ڴ�?9�B�'�|��wn���C��ɂQ�.]ʢ)]���(�i�BU���	�_�l��OP��'(�TO�O������,|"!%�5+}6b���ɺ�T]���%�~�A��70���@:t����b�Y}��'���(��'���'��OJ�i��� J�e�
�8��ust�Q��>�K�4c�O�q�S�'d�*-0�f_�C�F�â�>!V�l�*4���IٟX��˟l��jy�O*�k��2H����"ȅ�������:o,6mڣBC��B��������ǂS�R|z	���kdx� V���M{���?���`���(O���O@�$��L�4(����i �> ��Ū�i+��'M�,�Q�1��O��䥟����
s�p��La&Q:@}���Ĉ�H��˓�?i���?��{2^!aòQBc�\Μ�sT�Ǿ��D־\��Ĉ�OT���Oj��?	@�D��Y�6l�e��	K%XI^U�,O�$�O��$1�	���)��ZȀH�,5����
�O�X\P�.>?���?�*Od��5Z9d�Ӄt����b�A��M�3��D�47��OJ���OF�<�		u�֭(�bӔ<�u�0b���M�>P�PBX���	Ο��'�#˿Sy��ПغDB3Se��XD`Q#]$��"cU��Mk����'�R�G�qr�l+L<� ,��#Ʉ;}�거�o����lJ��iB��'"剰d�������	Ο���I�@���
@;���K��K��e��}��'w�8�F�7Ę��4�r�Z\����s]Ż�EL�8����?��k�!�?����?����+O�.Δ&�T,R`�>���K6�ÞFg�IП-�l�G��i�((��a�o(�$i�I �92���Ʉ-��'$�'�DQ��ܟ��Ю��<h�������7
��M�f㕝CgF�<E��'���SN�*NR$�0�b�+R��Krb�|�d�OR���2dX��|r���?��'@�`����E�L����
��8��2�?Zs�8M|2���?i��l�¼+$dB ��	MԻ1��A��i����07٦O���O��Ok�ӡy;n��"�:P!�R"!|�V�'3�U!��'�R�'���'��R�hB��ARd��0j��T#x���'K�kwL��4�?���?��t���OyR�'�\��'IĨKàG,MH�m�b�؎�y"�'�'?��'��'�@���x���HG,�4H����	Y��F��]��ğ������	jy��'t�P:�O�H�y���6��$��8���ʹ>a���?���?I�y۬0R��i�b�'��!�$+]+:��ՈdလF&�2`�wӦ�$�O.�$�<���`#f�ϧ��ɿz��f	H05�J�E8R:6M�Oj���O���n&$!n���������E���rhƔQ��!!c����4�?a-O��D �w\��5�4��F ���LuQu�*Ze;�hG��M���?�E/	$�v�'�r�'����O6Rf�ʔ���p�7m�i1v�Yg��>A�;_ ������|�I?EI�'Qv�e�'�5�t$ ��m�`�z2K��������	�?	�ϟ�	����թF[~$s���^0zL��M�Z6��D�O��|BN~��A�FL:ӫ\�Z ��I�m��bլ�#�i"��'b&U��6m�O���O ��O�NA���x@fG(Ơk6�F�M���'��1��)b���?9�Oɘm�1�ƐW�� �q"t� �4�?9�%ν���'���'�Ң�~��'`��mI?y���;p.E�f�$Y�O<5r0OF��O����O��D�|d�Y.ZvT��7c�x� �����ԡbR�i�B�'�b�'\������O	u���- �m+ �4O�I�U
���$�<ъ���?a��?!��n��,A�i44�S��m��A�H��m�H��B�i�>�d�O���O*��<i���>��'1o���u�#"G�,��8�L!ղi���'���'�Z�'X1�h�#�i%��'�nt���پR�1#!bѨd׶	��d�t��OF��<����8̧�?��b1���υ5=P0|C��ދL��4i1AC�?���?��per���i{�'�B�O���x��S*6 �{�dT�x���r��`�p��<!��z6��'���|n�$&��2w�Yc�v�is�J�.K�7��O�dnBW�&�'/��'����Os���i�x�BҢI�^u:u�.:�듔?�F)C-�?�����4���Ot2�� �T�JaZUIL��2olZ޴fb�b�icb�'�2�O��$�' ��'� @ʰ���r�d�[��CM~���OxӬu[��O����<�'��'�?�P"�s�ܸ���3j�f�P,�(����'���'�fɒ�u�|�$�O����O����,��%
�s;�1��I�	���s�iu�'���2�����O����O�hц�V�z?�H ЎR"s!ܬ;i����I;2#��Qܴ�?���?a�>���J?�ӄ�%/V�mسH[J0ak��Qh}Z�����?q��?����?����? ��P�]�թݍOD8TAM�i�`16�i���'("�'֦���d�O";&�ʊv>���E�h'\A3ç *���<���?a��?y�-���i5�iTVZ&.2=�p�S&ا�T-�e�y�����O���On�d�<)��TȆ	ΧG� ��DF]=_&�H��~�
(�d�i�r�'r�'���'J��`�c���d�O,�Aq.H�>��}{����_���Ғm�妁�������Ly�'eH���O2�#|�� �oZ����r�K�5�En�՟����x�I�se�@��4�?9��?i�'46�lYr�	�^��s���̤�ºiJ�\���I�j���Sr�i>7-�WldL�u��?8����?,����'����
Vr�6m�ON�d�O��I���$
��>�Bd��
�VL�R��%��'
�	�$t5�'��i>դ��Xrf��
O�)���jPH|���i@pj�i�����Oz���P�I�OV���O�Y�CJȬo�P��Ƀ���lc���˦IK5�ßX�Iڟ��hk>9$?��ӛY��UD	�N5&i����C@�Hٴ�?���?�oL5#���'���'����uH3E��tj�k��A&�Ua ���Ms�����6��?��I֟8�I3E�T]Y�j�o,�-��ܤ���ش�?�ꁷ9r�&�'�b�']2F�~��'�jm+��ѴΎ�)C	�%�8�+�O��qd���������	ȟX�'�-�A�t��b3EJ�-(F�;acБ%�BOT���O�OV���O�Y려�*�M���l��C�!�Z��O�d�O��ľ<a6��g�I�)f�|)���ަ!i�A��DؕG�	柈��k�I柌�	=,���2iY�(��)R�0x����G[�Q�OX���O�D�<i���m;�O�(�R��j�$�It�D�@Ä�pӨ��9�$�O��d"w���1}b�K$N[~a��H"�,�f����M����?�*O�0P�$�g�S��S N����E�X<;Vi@_��AO<!��?�0j��<�K>�O�&��g	��}��j$�:��4���	S�t,lZ>����O��IB~Ҍ�+`�<Q'�ϨO'�	"�۶�Ms��?�����<�N>�~� j4��C�Qu�׺9@Rt���iUD��r�a���D�O��$��>9$���	�5n8%��4&� x���m����	�^�#<E���'y@�!wJ�R�����bS)�>0�b�>�$�OP����(M$���Iڟ�q���Sʖ�n��5Z�I�4�ElP������H|r���?��!$����GL.jyF�q ܔB\}J�i_��>��b���yy���5V�[1M�D�f]�1rL��(���Ĕ�$��<���?a���$ʜ`�.<ñ�NZ<���X=_G�ɣ��s�	����I���"s-t\�ׯ����@�F�9k˦Q���Eu�	��������'r>yƯn>��K�	��"]h�)ԣ�4����?����䓀?��1@���_�2��g/�Y���!�[����qS���IƟ��	Oyr�JV�B������	q������:t�:�b�e�5�Is�ȟ0�	�~,u�	F���>3�$�%���JیLB���U����'�BY�d��%��'�?i�'63N��%�K�$�vUbQ��"�h1��x��'"���O�S�#@�"6Oک�08�R�A�7�
6-�<���_�欠~�����Ґ��rP �_p�Xs�A
	�����>a�R�H-���?(O��|�xtkSw-Z�1�M�0q�i&5�C�e���d�O��D����$��Ӯ[6e!Fތi���Q�%��[�d��޴y������?9�2֑>M��b.1��.;D*���JJlЊ�4�?����?���	.҉��T�>��N�;�	����f[�L
C��������8��fD���M|2��?)�:y�4
��� $Y����T��`����'��P��'�R��~b���F
 \Ч.�4MsI率*�F��VY�8b��5G����?���?�*O\,����镎2�J�e�L�io&��CD}2�'i2�';����=%�>D�4�P/|X-�DVTH�ɡ�#�d�O���O���O�����?�zm*?l>YEk_ }ެ.��F�'iR�'��'h�~Ӫ��jT� 0[�'Ȼ���Kר�sf�3��p}�'R��'��'����t�'�2�'E����S>��rSܣU-�A��*z�\�d �D�O^�d�lt|�C�xb(O�pP���u��[_*�A�L���M+���?�-O�TЄ��x��؟��S�p�Vy�f�L�Y3�`u�)}Hv��ݴ��'��)���i�f�q�+C�����3|Wr��ݴ�?y�qc�} ��?����?��'�?)��{V���K������WhX�&T���	sy2�?�O�O���S)�
4r\xeL܉?����4&r��g�ib�'��O*Oz�$�L�&�r�)�) &��RŦG��xnZ�z��#<E���'^n��A�,Ԝ���S�q�F�pӼ��O����"Aɘ&�����p�lм�D��4_��Pu`�
�N��>�2�S{̓�?����?I�&J�V鬙�Ңݮ&3�@�e�e���'IH�SU&��OP��4������"�R���"��A $��_�D�i,�	ϟ`��󟨔' P|R�bN�{l�Lq�D �.���P�m��O6�D�O��O4�d�O&��넭]0Z�`6_�P<��D�L�1O��$�Ov�$�<�b���f���B�/��R2/B�Q^ja��A���	ҟ�IY�Iҟ�I�%H|�E�(���G�?uh0񗏘+r��'b�'�rP���G/�ħKb���c-�-ޘD�U,�?��EAԹi�|��'R���'�D�`7.ֿT�^X1u+�]�Y[ܴ�?����D� \���'>e���?�`׀ѹs�0�i�@ơP�xl�0�M4���?���Gj!Fx���٫A��>�L3VH�8!S��i4�.D���8ݴ[��ߟ��S2���+h
�b(�(�dt#a��(1���'C���	�O���(���4S� s�(�(��A�ie�dV�b���$�Ov�$��]$���	?�@��@��!�� P��)S��x�ܴ{hUEx����O�y؀HZ�+�pIT��! �j���H�̦1��ҟ|�I�|+:	�I<���?��'.�s&B_"nY���Vn���}�Ꮭ��'r�'�"�Y-Fi���&�@�c}��pXg%p�s�4�?q����BI�'h��'�ɧ5�!�)Y���g`ެ0�HI+� S��DL�m�1O��D�O&�d�<і㓔&Ɉ�9e�^Kv}��N����x�'MR�|�'L��n2zMpv�Y�`�~�b4h۪c��%@�y2�'�"�'���?i�����Ol�G�F�t1���D8dHf���O����O�O����O�X��1�π�[x"T��jB$Kxј���>���?Y���� ���@$>�3@��X|ʐq���3_�m��*���M�����?���~��>�Wň)D�D��KOr`�Iܦ!����,�'t��#�4��O��Ɋ)%ǲaBR��E4 ,�!�b6�1%��Iޟ��g2�S�d�v� �Z�˔)/��eA֧A	�M*O4]u.��p��x���2 �'N�ȇ�P�m���H��Kh"Y�ߴ�?a�6�F�Gx��t��$Ry4��5��0%���'D��M{��̂A���'1"�'����6��O����d@�P�.�S���y?�yIt�ʦQ�Y��"|���$���c�@Ѫu�T�a�+�"X�гin��'`��܃�|O��D�O��ɞb�Q��U�T/�PQ�˩F`b����.;��۟���П P� �y�f�ԓ,�´h��i������i�R����O����OʓOk��;m����� ��ua�h�5QN��7c��b�h��㟈�IKybj�#&6�X��E�[�"Ax�����N���3���4'� ��埀��.�=v
���+�Ax>�{ �I�I:�b�����h�I۟��		͸���=_$�H$/g��h昣|(Xܴ�?���?�L>������P���L�w���wB�$U>!(go̲����Op���O�˓ v������]�(���vˑ#���ak��H�7�ON�$3�	�N'�b?�H��}�p�(E�ɦi:�!&rӈ�$�O��d�O�5��m�|����?��H��;�iܚ3�mp�b�)�`8�Ǚx��'R"�n��p��y���t�s-̞)������f�< y�i~剸ᢄ��4  ��ʟ��S���DIw���Rd�^	�x�U�J�3n�6�'^ҍψ�O���@B0��Bd�q/܂y����i448
Ѫp�&�D�O��埪&���I�	'vm�*
�g�~(���`��zڴ�TLDx����O��r +�/KB���N�� 6����Lɦ��	�$�	�侩;I<Y���?��'.���e����lp�cǯy�J�H0�]�<-1O\���Op��U�j5(ALEn������y8Pn����!B�����?�����31���@��A�&�G=I8��RDd}bm�9ߘ']�'�Q��y�@�w|��E��5d�] EL�r (�AI<����?�K>���?I��7]�p]"� L�Y�ʀa�J�z��0�<a��?A����&%l:�'y̔@ʄ4U�B��E��#!w6��'$�'l�'%�'S�=�O�-)3J	�66���Q�>)6��7]���Iҟ ������I(|j&X�O�"f8>B�Q�5�^?B���⃅x��7m�O��O��D�Oڭi���_6D�zc�U��v���`]�1n�F�'%"R��a���ħ�?I�����7�q�Aʬ�.	�L�ܦq�'Qb�'��"}�'����O�0��KBaˉubX�ڴ��$݊J>�o���)�O:���z~��W#��ݫQ��+������ �Mc��?i����4��<	��{���,F,s=Ω�w�O��i;�fM�6����DR�O&$����$��Ԃ�Ɯ)u�jFX={M�Em#D��%��
�0-�q����A�f5e�r�PЎе�b� 
�ZY~����� �`��� ���HUd?q�"ej��C(��ŬF[*
U�&�K�\
D`B��Z�B��d U�vf�<SDb��9����Do��Gj����N�H"F�H��l���+1��2_�%x� �q����X�I���	�ug�'��<�6\x0BN�p��*�)X6�sO��w>�0X"ƛ$H�^���:9�<7MI�1%Q�4a�Z�n ��p�ӾRލC��-p쐽����
�UR#��#2YtAo/�@�<	 D���`�V�X%R�j�a��j���ڟ�F{r����GUF�IP�6^�8q�c�!�$��&�%����-cny ��;V�1O��o�� �'_�m""�>��x�b��@���uXpq�f0\�&�����?��K�?�����D@�z�8��8s��`����%���}���7@�ԆٚǓ\�Z,��!
$3�P�-�۟�v�ײ��u膈5\%qÊ0Oj\���'*D6-Hڦ-��4$��H�$� a�L|BkY	�$�'#B��S���(�1/\�0�`�qt�S�:y$C���MkB�8b[z����9��������<�-O�Qs�VG}��'��91�^�I)K�j)��.20�Z�,_�P,���ʟ��E����;f��{���S��X>��P�Вu�Z4cwS"!�1��4}�:s.�XG�<Gt�+���J�4�Z%v���[� @�q *�'�"�����?q��i�O`(Xf?]�1�d&�8�p�I'4�D�q��ת����)Q+��(wc1O� Gz����14*=��S�4�B�;&�!x,��?��K��]����?y��?1��?���\fb�A�!�<Pn������	j���
 "v�T��F?-�����,�3���JS�Hk�ɍ�>= -�"�g�Ȫ��Ĭ0� ���ж6�4���|2oK�FGi�� �i�D�A�1[�R��\�`��O�(�ze����τxy�ԁ��G�*L��61���h�:^x��c�/-�H�'C#=ͧ�?*O�؃@��f��q��p�J�K�HW d��F�O.�D�O���Ϻs��?ќOC��iV��hx*�����2=!�!3��l��aAա�<�f��A��7���a��M�'��M�AE�����Jt�����0K��NIz�IK�=~��j3�(`p"t�B�G�'"�}��DP�~�rM
��#EѴR��[�?ɑ�i�N6��O���?q��_
�t3�A��=�|�3����y"fXFʤ�C�>8�L�g�)��'G�6��O���&����iT��'RM���Y!Ŋ1��p��7�'��&�6���'s�i8qc�*>�DK�xS04y���3���Q�(��x�M�� �`�x�"Dc��'�X$P�U�E+�,�p<ArK�����4-c���'��ݐ�EK,j�N4@ '��02! 2^�t��V�S�O}64 ��p��lZ���լQ�	�'��7� �����<����tb��\P�3O��:���b�i���'���SZ`��I�%��JU(�yY m�tg�1���I��q��Y0���b�|�)���I7@�JܒiEg�.F�l�#a�>i$���y��m#d�x���$�
	��!.0�*�B-Ϝ��	�\`"���ަU��4�?�������5�bx�0/R& @H�@����'��'���K�(P '�P��D�C	쪴��9~�����$5l\�1��{��Q2'g	��M����?��.���P !B��?���?a�ÿ���סT�����ٴ$yd��C���OTI��S1��'e>BWd
�{����p�:K:x���:���1L��HQR��|��إJ��r��}�)p�ߠPk�7͔Ty�H�?�}��� ϓF��f�]2��l���5|�U�ƓeNp�p���8`8(8AVcB;B+&��'?�#=A/���Kr�a��S	iyb��5�5%�0)��W;�С����?����?�����O��S�i�؍�/�C*Ƅ+�&߱R�r� c�0/���Z�d�(5��ɣ��x,yc�5r��"�l�"d9���d�*�(Y�S��0�r����!�?�\�� A�BN4m��f�1��H��d3ܴy��&�'����?�㡑T��B�EF6;���C�<���]�ib��Pf	�	�aR��~̓y��i����5Ƚ���?��s��i�/
�`Ǝ�X����г���?�v�֍�?������[˦1��U�/�PP+ti��\�Hm������`�g�o�|���$h��[��y-|��b��f~2}9�焛Cᔤ��ԂgL���q��N�'o
�����?�.O�8�! �m�l�� ?n)�p?O����O �"|
�fH�{����W:d�,����|<�W�i� �@�i㮐p&Hʈo�U��'���tU�;�O����|����7�?�geB�,�5�@�Zt�9;Ub���?�R��\҆A��dC��CN�	�ĸBv\?��Oj�X�4n��n5\�N�t��z�d
S�Z-��.�=S��kOC��b?�QE�	*2��ȫ�׀A�����m?}".�?�ĵi�\#}Z�')C��1���D��y��Aڢd�F	�
�'6nD���U�
|�(Ʉn�I��hÓ{S��@ZE��v���pW�P�EP6���M��F��O$��O�C$�Y�"i�D�OZ���O�(e�Zy�1�P�~�`F�fo�Swo�)!�)���G����5�3�$������n�S�Dr�&��n���P��M���	�v�9�5��|�� �?�&�K�@8W��T��@W�
�(���O��O>�!e��ZlV�x�A�(~���"..D�@פ��(.��B��(���0�'2?� �8��$�<�KP�_U`�Wʌ"S����ە=ƒ�H#�?)��?Y��ZT���p���J��83�E^m�ĉ�)�"Qt�YtAɨ'.&��@`G�R�	�Y�B��(]N�����A����X�������@�#k�D��ב��(gF�N��di�� Q?B�&A�U���t�����4�'�����X+2� !��B��f�����D�7�|�ʠbQ�FN�YcȰ��'���Y��~��IL�L��Zw.��'��$c��U�D]v����[�j��Ppw�'��J߇.%r�'�� w�B�|r$ u�V���\S�b㉁#�p<�%�s��}X�u;����7��\qbM=XL�4��IV��d�Oj˓�f�BQ�C9}�
����95�<��?�������c��2��iŋ�����#Oel�=��9�ԃ��\]󀭌�C!��I~yҤF�+ ��?�*���bd�O.�۶D���T���_7;Ir��C�Ot�d�!h�"�Ґ�Qr�=ҭO�N�e��q.q�P(�5(A�� ��Zh��1���Q�~4����=n�J�ҥ��31�����d �da�	��M�#���?����y�Q����-F>`�g`[h<�58�\�	b��%jyD̩3�v�<��K�z��� g���ep�GfV3V����'��'�:Y��![��'Xr�'\`ם�.���92/�-�=��l�
T�1ځ)Ӄ��T���i�Re)B������8f"�h �
L�1�Ң�	D���  �bs(��s��x�r�rY�}&��Ca�6��@5E�4O͈�[5W��M��V�drFd�O��~�DpdO��nh>Uh��ƹ[��%�v�8D�h� @�yAf9��i#��{�1?���3��d�<i#�'��	�kJ�Դq'���Ybf�:U,��?��?����n�O��u>��F-T@��y�bG�i��l���5i>�5 �DE�B�D��o$LO� k�[12�c�-��Y��ϒ5�ι��!0����b�'�^л�E���|	dD��&��	�?�G�io�6��OH��?���8$h��K�G$yS���m��yR���O] Xʇj��B��ѓF�)ʘ'�*����D�..��Q���?��S�? ��:�!��$v2�JE,y��b��O���{�L���O:�S�wZ�,�,&x�3O,i8qk�).���h3/�/s0����'�`D"�C����$����h\�'8�H	Q��h��7O��0�'��'�2�#8inY��̕�}F����L�7S��I�H�?E���ί|cD��FZ�| ��(����xEq��q�k�7p��Q˧T1i�d̛���O��b52,�!�i�"�'�哱!à��	��ƥ�CM��?;@ə�̍�?��U�I��a�$YK��@�@*Q*����4��i�|�BE� ^���
&�'j�L�7�p�$P�t�����
X&nر�2d�ls��D$�1��D۷�8H PqgR2��I�p�����OT�n�4�R Ã>֠��3��JiR�;��XB̓�?�ϓPf*!��F�vb,�$�5K�ȁ���0�M�p�i��'7��83�٥|��9��R>*����W�'��'1�m�"�Q�M�P8E��MT�-��'�t�
1I���&�
�1ȵ��'mX�c�A���T�OP��'�P�:��C�m�u��!X)l8\!�'��h {7������>0'�C�ɶ>k���&�[�e{�g :��C�oA��X�jɕn�r����3ǺB�	8He�U��S�E4U0�*+P��B�*�YFi������d���8fB�I�3|��f�K�R �A�`O��wjZB�	�h�bQN�-�@Y�1돫e^\B�I;��`P��"p�{���>}��B�	"y,>I9�N�+kH�� ɢ�lB�	/B(fz�F�Par��ڀ/HB��Ҡ��K��~t�ӅZ��C�rn�DX6F����(x<�� �=D�ȳeiB�x�"�
�g���s�<D��#�Bѕ�Fdz��G1O~����;D�8�IOc>l�G+��+�n({A�.D�$��㙟
���ʅ>�p��PH0D���r떏jx���Lw��s��1D����DJ -C$����[�j��"�0D�`�`�
7L�,J��^�9\���(-D���#��W����mW4&�� ��"*D���6(��U�B	{���e_�&&D�H��e�
���D���)�@b#D��C	�a�L�b��(���r�A!D�$HPE��7h骱�@5vu��z��>D�<���8���i�D��{6�Բ�l?D��@�D,[#H�s���M���Ђ�(D�@��eJ$����1,�>1��1D� �P���xN�<��cO:|�;D�x����.1��i�`���H��E#D���0���-���G�@��H��!D�|X'!�k�&4�P	��h��?�O�i��ϧ5�r�0;S#�����q@S�"��	W�8���ƥ\��`cb�#3�g?����L�*�Q�@�P�Z�р�I|�'���b�@=�[�o�-�i��ܟhhc�44����a�Fܪ��⅖P�LA��K�[�n5�å��h��$�Y�m@��Y`E���'��9o��Mh1��X�3�%bFjO'2 I�ϸ'�8�g���e�����	,�I����8�z�Y
���h�&N����F(UzބBE��&���$���n[qO�S�ޅ̻{��`*wX\0��m��x�p���
w������ƹ%lܑb��
���`��L�&2r8��4V��y��!�H���A�LV.gع!���5����(���I
)�9���T�pȥ	4ö"=�-���$�eZ$j�8�Ѕ
���$噆b[��X��Qj^��u���oҞh(�-��d��D��)�Zw�Q�A%�Ihz�b�]Pnda��m���%���D�B�ڭl,�3�B�|R��i�~E#��3���KU�F�,��y�Oŵ%��B2/L��ju�f�'q�Q���f~x;�L <��Y�p8ʑk2闕C� ��4&��=�F;v�6ܰ�j�8��#�2�h���W�N"�`�B��#�H���'Ƕ��[�I�t#�q��R�D\����&�ȧw���n�U�������s^����Oib&��������[?9�W�� �[-A���%�Q�'���C��#��ݚ(Ah	�aeG�m��i��)�f�� ݢ.`I�RY�"b��������X��$�>� �l`�MY�X6hآA�ȿ �4��V�i�(���/����)5�mb/�hQoZ`�pl�Qm9(�r�z��*a>���1 (&�^�2�#��^:���ɮ�5� B'm�W+�4(��YV�A?�?�2� �15rm�&���M� @�JR=`��W�mX�}�3���>�E�͖"[��p��5�L���(Nax��6H��a��U8D82�C �i����ad�q��E�y����v�X,��
���Х�L V�6�Р�ԀM�k�S_���O�-��c�U���a�� �Z�����(Q� *����!IӞhMӇ������j�LXR�D(�剢8P\{�A�&L�Dc�C��؎	ȇmЗw�9�Zg*� ��= ���@��3B�q�(0�n�AT�	S?	j?�Ѧ���&A�9<�u@%HL�H"�0��ՌVE�]*��5u
�ŉ �C8�(R[c�@�����*!���6�2v�!D���yt�R3fD�A�4F�0a @}>u,�x��VF�	NƂ��1��7&�>��1	�35ax$�)��0����	`v���'H�8��1^�Zq��,���[�O
�H��G��\S�Y8b��&����O�0��˺Z�p�%˚l�F��0�����C�uYЌ��iP@� Tӣ1}*�V��m]Y��hD�7�f�vd�Y�T��͈�V���ygdF*!��n0� ���BC7+BdR����f�
��=A�4ur�*TF��|�>I���[�L��#�M�@_HL2���T���a�$�O��x��96��,�vtf%��'xvEy�O禀R&��8���q���0T@�xq��IՄ����'`���իKn�I�"�TF�9��������C>$6�P��K��HO���Dd�7�p�{ǩ?R�D)C�]����
�:H�2�pWK��K��,?q妆p�
)���9S�Z�S�NF�'k����/U/B�n)���
U�.�{���
yR� `�"9�H���	(<�x�B�Y�������I{Ԁ�a^�Qp����=R�1�ִ��W�t�C�aO�xR�YD$mYaE&�^��1A0#�� ��U�V�I($!�<�U�E^�$ 1���$l[�l 0J��B�F
\��t������0<Q�M�u"P���Du�-228
������	`P�A
-�h��[��D�*�Ri+1H�u��X��K'qO��w�قR�& A��+k�j� Q��LB�  VB��3s��B���s��vA�(�LP��X(�H]����S���,r.���($.��ب9��Ps���J�KCxYnڼ7��� ����d0?q�� /���P�������ѡ(����+
%5 a���P5�!�d���\ �@a���cN`�F�'%9B%�� ���r�+�+d(�cR
��l�KDnީpd�A8��`�ì�7+��i1��*�O��f,�5Ul8�&�
�D� 4�uF���D-еf�l*�P
�P��i��A�"�Q�"����$���D���j�>s��1S$a�푞�j��)���b�O�i�'�&=�� ӽkU.H�P��  |]�&b�1z�"���퓤M�h���ɡ?2A���ײ@�q�����2�$$^�|,	�'������$N *ƽ��kB�~e��K3&���u)������([�<w)3J��0#��I�?��[F �[}��	��yH�0F�̩��	�>���,�?	�,�O���A`��]�F�)h���t�,0`���H?��q���'�ąs)W�:(����<'[��z�FL8pr�2Ԧ3���d��0!F/�^S�QxG��������:1�G��nZ�k���6��g��Y��c�(Y�:�.�:/��`z �5.��z�����8P$�VD|����@��H�S%�n}���-�R]�3���b�.qƀ�d����hI�ܓ�a}� ̙g����-�5~����κD�����F7�X��Ppn�I(O�B.�R�������O�$��<z�ĳ�I?kKb�Ј�䔦*�� ���>}��X�����e1�	�R��A@���W=�L2iJ ?�DOz��0l´ ��� W��H�\�;������d�xqlGv���q�E�u�6�,Y�����N x������1��OH�Af������"T@T� � ��qc��H��p>��*��(hcTʐN�T�*T�� ^&�Ȉ�:Oy�dJ��F])���¼�@0p�&(Hr�ι(�t͐��AX��%-\G� �C���/��[�!�=i��\� C�]� ��-&�d�<a�DV�^��<k��L�@ê\�$��f��AK�$c�rAz�L 6
D�`a���Mu��!@��10(�%b��D*_�Q�S`]93�@4	Нq�B0�'��#�`�{c��b��F
�
�)����g}
Q�!"��8m|h�%	�*m���_
�T����-i24���%jO��KT�+���ҦC��~�KVe �;A���0'(����cQЛS�t�h�G |OH�fF�+HF�0���_8�8�x������1etɻ��� 
$Ό ��O���x�;ʲu�I�[=�
��=p�����;��ѓ�KH�j�x�� H:<��i��KE�a�6���J
���'�vy���4Z�*(�=�O��e!ѡH���-���;T��B��de���ԬZ�;\�y����3�f��)9���z�L�)� 1�baպ��7�؉WN�P�& #�����OB�tͻ9�Ŷv�踳�� �X�`��i��`��3Y��4A�(	Wl�ͻT�s���C���^��|�T�M�d�:bA7}���rI�t8����(����ò��'���s��\�&hj�V�G=j��پ�����a��v�`d{ЫV����E�� ^���ĝ�!R�bRf�(Vr������(z*Uf��>a�)טQL�nY�e%jL�%�3�h,����NY�$XR�քZ�3�֒Y���ꐝ��>���9h�L�b~�ޡ��D���#=���<t�&���!o�Ih��J)���� -,u@����R��)���!8� �FJA%px���Y�f�<��4 �X���X; ?�1��Q9����������i��5�%�"2qX=�ũ��A?(`@�s��zn�7hK6��$X"��A2�]�S�6mȄ}��%	 �M�~�����̶+X�Mڋ�Ή8������S�G�"�:�@:m���g�oB��ȉ �L8Bid˧���/�wi��QƘ:|cv�{�(�#�~B��tU��n�"�s&�V Ta�{rJ�A~0
�o�K�r}���!��'9r|�g�	]/�`���v	�3�ȇ1��oY'�Dg˦F~���e�ps��)��R��yb)�j���Ai۲�e�>z! �������0eH̲e��6���':� �ϻBŞ��,	>dQr�J��s�6��ȓ�@�F���|�b#Ж�*�ۦ��󁐶K�|%�Vȉ����"�.�y��O�%�4h�X䤹����b����gH"�y�AF�+x������i�����0�,	$a��4<�T��A)^����!����G�]�L�Ա���_��t�F	�;,�Z��0'���u��)cw�Ղ�X��%����+�2H�5��9dF�1l��DE׈';��"�'�� �ңmհ=Q�P���,,C�t�z�Y��p�C�I����!�A�6���A=`u��U;vD���?�⃤r��I�3Z����E��,�T�!��ԂB��P`'�X���'���"�6Ĳ)Pq����
�h����Xc���U��������.�*i��4P�z00�ξ[��D�(Hi0�eQ�7�I�.G0XB�$c
��x���8�v�dy�A0��߭w)�R���'�΅�Jp5����'Z�B���r����쑊�੸��D
`�0xh��Y����嗒� �`����9°����~A�whdu�!��i]|�rK�Y�D8N_�;�����~��reѕ,���n�(]��8Bw�7lOҬ��6hN�G�ڂp�phvb�<od��9&�~�������b/���&Y�'ڞ	�%Ȧ���9^��'Z0����9�` ���]�N��B���`�d �>�d+�Y��e���ת����9m$�ԟ�x��D�̰�����( ���ȞCy�h�2��܃Ѩ' \d4�� ^���?��d�W��)�C+�	�V����N8���s����|42�b�aE�]�ԟr��f���.T��=�V]Aӎ��M¼ɡ"�)zA�X{�i�7pe���Ċ>j�~���N;��Y����1y��b �0���'w��1��Hv���+��f���8��>gx�e����+X 1��I�^hA���qܘ��
�]��PÅ	�n,b7���)
�aU�S�t������"�Y�¡	
r��E'�3,Q|�j����?�cQ�C�4
�����BWkl�x�q��G�D`�I�a�C50�i���i��t�B�M1l<f"��&Ժ⠅Y�T)5��.w��Z7AR�/F��҃�S��j����\�1�4��f�<��>w����%��a�n��R�Ԁ��c��)1��?{�ؙC��4����bS�6��m�1�l����e����`��À<��<(�Ι��P+��k�����+e�A���;��,q�N2HX��P�� �}����a�"'Ip���A`�g�	��3 _�?������pu���Є���!�Xr<XL�Ɵ]��T�����t��cE�̦()lɑU�L�(�UI�?M�Ώ>}�U�Ł��Mk�/r철�wh�>r���N�♅�Iw�"���Msd�dCE� 5(ya���6>�&)�fcl)����|M��f� �&rB�UѸX"4��ϊ ��(pMS�"���>?�Op����W�U�$\!T�HfD@/X���ZH��e�pa�EJS�q"��H���;P�)Zb�$4�#
�i������	5�����O�I�!�	�/�H�Y�>�Q`6ę!�A��d��qA��(	�FxɦFL�&Tn�3�Ǎ�
B�� ]�m��N5~�]qd�ɷ��m�mƶ�hU ���5v�}Y���6@���>-�B1�|A�@e��#�XAB�lٷ �93"O�ѡR��/�`A�;Q��tK�"Or�#��\?O�\�a�,u�Fd��"OT��vNWv�
8�B�8�0mq�"O�m��=%ފ�Q�AA��y�s"O�m�#���Q�!����'I̎8��"O����Q,hT6ә�4�b"O�U�L>Xp�	�bB ���C�"O�m�z�di�!�Sݦx�h,D���B�B Y���l@�m p���e5D��a���8hʼ�1`b!#j^�Z!�4D�������"�bC�W	*)P�Z-3D�x���� [�z�P4�=R�n��%$2D��qFr��С�׌����M2D��S�eǅ Z(�@Q7:���	�k0D������@����>iH�e�.D��cp�Ġ{A@���(g50�B&-D��  E�\5 L�� Q��y���*D�� P�!��tі��v��U�*���"Of�	S(RIr��яP%T���5"O̕���1j9YAdL��L�P�"O���b�R�*�+D.�x�pU��;�y"��Y��
���h��{4�R$�y2-Om5�`�7^>R�$�ȟ�yR�R�y��)�!(Y
M�J�+���1�yr��WrM8a�ęF�8!�ڪ�y�ҜHL"�9S`P!A�H�0b�� �yR'Z���-��H�Z)H2M[�yR��5!IT�Fc�7s_bT�`�B��y���D�`��u���wBtt�!h9�y��ԑM�aj�cU)8�Ȝ�P�7�y��@�v��1�i=#�X�v��%�y�����tAH��()�f����y���'h�8�r	?�j}�E͋=�y2�܃i�`�Ru�80|P���y"��
V� Ț���/,� T��ƅ�y�ʝK�qH�!+�$��t�Q��y"k�<"攡�V兑#��$��2�y�J
�O�B��p�_�G���@���y����T(j�j�T�����0�y�
�3a/I�ڹ��% <IU��ȓ ��u���ɌmQ�l��; 3����Py�8�VE:�P�h�	�I�8�ȓm�D� ��ɵ:^�2�Nޞ��up����Z�A�R �A씒4�*��y�X�jF�B�&R��$�
O4��ȓP�@d�P�J!^�̚�G�)/z�ȓuL��/ͩ)LRu2Oζ-R��ȓxh���-��t�v��n�b��u�$A	��$��2���n%���sÎ\ۓ���X��I��ȶX<�l��(��p4��Hu�p��F$��ȓmL��{��Gl(P�I��3�1�ȓ{rhјC��6�h��E�� �v��L3���'��I4�H�BK^����ȓP�<�i�5)9�Ӭ=�v��ȓK�QBAL�5N�Y�a�Փlz�؅�l�E�c�CW����G\��ȓw�ʸ��%�6#&t$ ���q&���ȓ/��z�)�u/���&�7k[�<��d����U�e�dM0��7t��܄�|5|��KïkyL�� ��5؄�X�b�ȕlE�jŘ��.8�؆�9�Pa��?I��X��L9<O�<�ȓU�L��b� t����S�6hψ��ȓRA�Ex��_5���-��MSClTD�<Y5B�4���Ed�>T
��u�F}�<a��ܞf������/r�=�$
�A�<Y.V\�L���J�'2H�C�E��<�L�8K|j��S-U���yf��~�<1s�P�XJ�f�ʭ<��`A�a�U�<Yq萗y���
4MÕE����˕T�<�PK����X	����<԰�&UL�<�`�H�8X�p�?�1c�J�<A��ړ��:��<X�d��AN[k�<� ��`W�(��U�]�4�񑥁l�<)�jA;>�	r����܉� �g�<)��M4Ys�H[���bf���g�<�����{����ڂD��Q�e��M�<i�CƛZQ@��[7c��(��G�<��l]</X����#�/R��@%-BY�<��-an��"-�	@8�YV�i�<� �1��M��0$�5oF�7"O*�!�J&A�	TCʸ2\�Sd"O�ԉ��h�P��X/�d����5D��*Jn,��8��yzg2�	j����EG,Y� ����
BBt���1��9�S�'\:���IR7�f�oI)KR��ȓD"H���/u|L� ��RL��k_
�srEG�#e.h��	ȳ%����G0�� Ս�x�6��N/A��(�ȓB�A���	`�p�Z�F�u�|eG{"Z�G�T�Y7,p�C��<D ���y��!J� �C�O�MHH�D���?���'���p6�̠u�ʘ�p��R\�)�'�ʤ���S+�6X����>�X$˓�(O��6f�#8�����!^p�}c�"O�!2�-6%�����!%{E�"OfI9TK6cu��)�΁�P`��b"O04:4�\��9)s��)Fv9"�d;lO���O�~�#.X&'� �$"OT�B�"�4c����Z�#b8i"OV����FX)�,(+���1""O|�0��$#c��d)�#<��]��"O��q�k ���E(� pr��3�"O���dH�/@�A�xm�2��'���>~p�0�&���i���ʜP��B䉭HE:ʁ�
�^�>)���Ǉp�tB�I(q�(�5��x���,P�Y��C�	����h�?$����	A�6��C䉾|xtT c�3���k�2
��C�	< ܨ�o_<5�`��E�C�V�fB�	t��q���؜�1�
�iP�C�I�6��	P"ĿM�uw��9=rC�I�^]��:�gܢK��2S&B�=	T���#��<V�^�I ��f=D�Y�o�X�!�DԮo��(�� �1Ar�ܳ�!��K)+/ZЊt�^1���;mG<%�!�Đ`�f���������w��h���(�S�O��!�-�&���
H֢���'�*��%���;�)��=�j��
�'9���N���{��ڜ=T�4�
�'��@H�N�e�m��'�=>�B�
�'3r��&I�8�+�<6����
��hO�4(N!cz� *�|8CciB8�y��ēC�v-; 	�L�\{����yr�H�EJ̡���w��T���yr���G� ui%?g`���� �y"'A/8�4π�n�JX)d�Ħ�y�	=+��r��وk�L��ƺ�yr�ĢgBܬ3QJٷ[�Y&���y"*C��0�PO\\Z�`[!�0�x�'����'�ğ�0��˞+Q�h)��'���D�īw���t�ث@	��'�|,���Q���D&��,�	�'� z�K��]t4,��`I� 9����'�d�X��w��p2Ń��OiR��'r�DSê��e$
x�%G�:��N<��k�8��V�	+vj�5r�Ӣo�
��3b���2C��/���m�6N�E�ȓe�N=8��/� ����}h�I��	p�`�����k@�����^)C�RC�	_r�a��G3s���䝃6H�B�Iv\.��jT�o��X1� N83 �B�I�K����®��P����E�c¨Q��'6� �nB�?I�I� �B'N%@(���>��� 8���%}BB�hc�,:zL\t"O� V�Q�T�1z��+%���k�"O�5��\4q�6mQ�R�q���"Od�k��_�
����Ӕ�.}C�"O:x;��<b*��څ���O�|0(&"O���N7��8)�Oц\T�|�4"OR�J��	v�8X�NP5+'��B�"OLʥ����i��̘>Pz`�F"O���a��Ix��G�̏t�d��0"O�T�o</$�a���!$��E"O>�s�F6�BdA�k׽z&-��"O��ţ �Li������$�<i#"Onl9�BL�u�4�!��!r�<���"O�YbTJD>n�pQjB�͓ �
�"O�u�h`�q�G�1�F���C��y"O�+qQl�����B�m�qƞ��yb�v��aR��4E$����h�y����x��\�d`�Ns񉡏N%�y�.Jً5��K�hT��gM&�y�"�"\tHj��׷?mTdzA쀒�y��ަIgZy��D<9��:�I�	�yR�M�[뤭��Bm����#U��y"#{2�S�ϲITL0C`�y"+E2Y�����1�pʷ�]��y��EFR����L�$�0��OҦ�y �|w������4�[��y�%�ԙx �ЂHp��E�>�y���nøu�2��*�L�ʔ/���ybA[&(6,hu��9!"�K$�O<�y"��06�>aP1&�Hg�ɳ�y�)F�wbD�ce�[ O��9V��?�(O����N0\D@h����)(�ٻ�<D�!�DK4@L�@�ҕ*69�+�o;!�$@0��de��
`͸g
�S!!�Y��\Dj��d����$,ֺ!�ć�s�j�'ן3FnI��+��!�D��\���ĄκJ�6�B@�Ԩ	O!�$ǹh�8����c�Z�8�%O��!�īJ��e���R�N�,�k$DҝA�!�dW�GZ�\����Af��ؔ��9W!��"�fU�c�5]O�m����%+�!��� W�$,؇�Ն_(��a
"s�!���Q��W���Z*g]!���"	Z��VI	�@J(���ހd%!�$�p���`�V4IA�TGH5�!��%� ��HV6!�U�b��<�!�$�%R+��T��!JY�o^�u�!��G�*Ę@��� /�I�� E$Z�!�˧Sˤi�U,T:[=�	��o�5S!�dǤeABi����)f̾�W��r�!��]Z���@��Z�4�{7�#Ex!�ě�g�����!T)��p0�Ur!��9z���Z ����B6!�ߪ[`�e�L�1?е�c��I$!�d^����t-� O�r�!ׯ��!��-F*싔҇����j+vtPC�	�)S萘7P&n�T�*Bf�7!B�	!)�b�EB�����cO�1~2 B䉭��ĂDe E@��Ы��0�C�	:ɨ�8�j@W��IC�FX�C��<*�v�Qh��ּ8�a�>�C�Ʉ2�6��*��\�n�@0�T,~�B�I
A�
��B��=J�٦�_[�B�	�Q��)���_��c�����C�)� x��4�̨T��qѮN'2�>�x"O����	K��n���
�T��0�"OT���ʜ�Uئ Q��:	� %"O)�`D�2RBqW�K�8�R�"O��2!;(�t�cKF�D�xu"O�4{C�͜zW䘣ࠅ%��E"O �!oH _�2%�,L6�h�8�"O�s$H?E>Iy�A�=`�\ F"O�� n�KU`��@���Z�"O��!&��9`�\,)0Y�}�$`0�"O�h��.�߸:%N˶D�3v"OH&��'��9k�l�.����"O�D��K̖x�ث�˖��ek�"O���$H�*Q^8�����9�ּj""O$�����
�0� !�Z�Q�����"O�`��:=l����\����s"OP�
��Wq�di2ꉋt���Jq"O��b�?BQ��P�o��C�"O�=�h�,>P J6B�KVzț6"O����MU�T4(��3kӋ{����"Otٱ��	%!�г%H:o(\�;""Ob,XH�D�ހ
�Ė<92��!r"OX��@}�H��f^�!���B"Od�Z�+MLP�i�Jȁr���+�"Ofy!�M�Z�j�BvÝ� T8�{�"O8W�K #KJ��GY�eF�$��"Oƅc��R�bDP1��`<�`�"Ohr��u�$l��&[7�9ؒ"O.��#��[>�@�^�zH�"O�)���0r6��vh�D,���"O� ���Fs���xH~��s!"O�ܳ� Ofˈ��C�L��+"O%J��C�|����$l�iU�P �"O։Z��[>���:�+Ï%E���"O���H�xi���H�=SC��H"O��Q�ŎQ(�X`��ɨv�J�:�"O���c�3<��|[�l��NV�{c"OT��e�R�:y�L�J?̌�"O�����ڧ:��9u�2�Bx�"O�|"W@�U6q �;c` y��"O��5f�U;�0U��EPl�U"O��;-ʝ3��l�hB�=�X��"O`��IĩDd��Y�H`P"O�X��A�8�Z$4�6$�u"OnEz���
-rV<����L���e"O�U��g̎%,�d���7�X-�#"OJ�!���n
��$R$=K>y�"O���U�E�5�\�����
{/��k�"O�0!�Űt���� J)Ze"O<X{����M\�$s�*ZU��4"O�ĪՊe��Щ���wpn�BC"O�`+d�ňf�T��o�%.jP�1"O�C�k3@�����Y� 	&���"O�I ��ۥh�=2',��$�.��`"O|jed���Az5jI''e��t"O2�qS�b���(F�Gl�9�"O@��u*zI��q�FP�Qy�0"O"Q�iJ��؜B�O֧W�q�f"OrY�6��w�"�(f�X�}�0Y�"O0����	RJ�9Ƨ{���W"OVPلo/yx�M�wǜ�p��"O��b�bR������*  d"O�%�7���~�R�aʚt^��"OVAb�G�uX�B&�ߴy"�"O� |hkP��W��(�����5з"O���!�h+Bًሃ-6�b"O:u{N�4,�1@ �{%4�q�"Oh1cc�F����T�J�|{F"Ov�kg��L4�ӨGe�T�W"ON%��cճ�x��Ӊύ^;,4pV"O�(��fƊ �¡{���"��T@�"O�ٱ�*W��ě�B/����"O*�aO	�P`�a�r��e��"O�ء*?)��ܨ���5PgNh��"O�P� Ɗ@�NI
aNqf\�U"O8�� M�,��5aC�D:g�,h�"OT�B'I�\�X�sE"��~~���"O����e�L�ї� 5��q�"O�]Q��S�8��A�/?��M��"Oh��AB��vh�%K0$J�II"O<m���Ֆ.���M�<�:a0"Obc�IR=:�� C�ͅ\����%"O��!���3������zzmQ�"Or��	B$ЖM7*��X���e"O��
r˝�T��t�p�N����"Oh���R;c�8(��R�<ݛT"O��d"�Xyhq�wƨ��"O&Ѓ��n�m��*�'�"(5"On# ���X܁ъ�W���2�"O$�RubG��&��R'�p�,l�Q"O�t`ǝ;���ǥF-�B���"O ���̟2�����ڞH��4"O,�C�/��$=v�3$���	+\��7"OVl�f��5-2�,H���}x�a�"Ov����R���a�	E�pcr"O(Es"6j���կ�-B��0�"O���3&�P �.ڶ)t|�@�"O�����%]~� +��%]��!"O�J��_�R�dPR)F�GU\tv"O Eɴ��0~rY�0/��p<��p"O	�.�+��-��ݿ/0t$2�"O�`�ǈ�W� ��wEУy6v���"O����%��tC��{���K!ȫ�"O�t{t�\��Dq(e`�"u�ps�"Ozq±��W���Ҵ�T9Xh�8�"O�D˷��#�z�r������r�"O�9q��b������*�\���"O6P���_,x4���$�8! "O:$!t�րx��a#d�;*b(��"Ox�1pDY.pb�(��wL�"O�ԙ�$��"ʬ
ӡhr�P��"Ou���kI�ygC�v����"Ox �E ��!4��RŁ�u��Tp�"O�a��͍�wvޑ�2AѴ�~��"O�)�&�6,Kb<"��Ń	��	�"O�C`�ë.ƴ�6
:v9����"O�H��M�m"F�S��wVĴ�"O�L�v�h* %�ՖM��2"Ox���P���2,�
Ѻ$�"Oq���H�8 ��j��!�JI�S"O�9)�� PH���=�4qy�"O��C�d��m�UcWKE� ��}��"O*�Ön2i$�#R�_%
�\�8�"O&�
��������'�=m�>��"O��2ң��]Aʩ����7FA`�!"O��+c�	���Bbӡ"�黱"O� ��)R��[�J��m��"OH � FX��.daE�;^Ƃs�"O� ���v�T��H��!�P�L���d"O,dp� T�}��;�c��S�����"O� �:4���7mM�n��p7"O�Qq��Cy����}Xv���"O8Ek��ؗ%@�Ɓ�4?ቱ"O�<V��	��������&�P�"ObD4⋴]\r1��]�O��u�c"O,-)@)��r٩Эٙ]�$��#"O��k�#\�R�X�Y��҂m��|ir"O�c��&Quh�S6h�fش�x�"O(�0��ՎN8��"���:+�T�g"O�Lsf��4Z�&�;`��. �ؑe"O<�2�	<K) ՛��V(���J�"O��@ �ɛ[`��`�!�|�V�SC"O��#$��u�^M���@p�0�"O2�h��L�v�@���`!#e��P"O��SBo7^ʷ��VH �D"O6���*@�k��Zs�I;yj6̹"OZ�رȒEW�]���6]E p"OT�S�+�k��Ur.R�7CP"�"O��vGN�j�Ұ#�fY7<�u��"O��'+���K�+��<BE�A"O,��e�,2 ���q�W5.�JC"Op�9aM�el�j�$	/�V<�"O��c@��<m�ݡ�c��t �"O�{AkM$�A�aX�y "O�( 6���b��1gNFZ�Pp��"O�AI�C�Ys8�ǫޥCژB@"OҀ���Y'i�$%��)"���"O��
�gǘR�$�iE��vfn��"O*l�7�˰&�h9 ��L D�]�"O*�i���?B�R�� �3�aF"O���&�NTB`��r��@��"Ol�zfᓋ�j��Uc�<�^���"OX���H@��kA��6g��t!s"O�Pr��4~���2�J�n��d�"OZq���)�`�"	<at����"O��
4Ȑ���u��Gǚd[��p"Op���V0_���z a��_7�a�V"Ox�S�^*g#���G�J|t��"O�+�fM�"�.�j�o�-c6y��"OJ1�S��::0���4�6��1"O������^�+�GɳM)�A�"O�$ItK�5i�=�w�O��=z"O\(@�c8#Œl����;j���'"O� ��N�=k��E�s�A�P�k "O^��'�U�~�,ѳ���E���"O���C��G�A�`ED���k�"OԤrV�I���q�j,l���C"O���އ3���.���#a�&�!���0�
tS��-2rXcpE˦>�!�D�pq�k�N"@`���e��<�!�D��/�,�Sr�"G_��+�e��MX!�ҋf�~x�TM��E Ԙ�P�!9A!�DY�Y���BE�p@9�J[�5!�DR "��	��D��$> �&�^1!��ƞsޤ�x�.Qm�(��eQ�?�!�dA%�t��g@=)! �Rb̞v!�X /����Z#
*]�&j�A�!���Cgx8c�'�V�<=h#	.~�!�$�4/���d��b�B]B#)R�i�!��F?pz����Z�%�&yP�ғ�!�$
'
X,q�rm� M�	�*�g!��']�Z��.AB����6S!�� ��ı��(X� Q%2�"O��d��_�Լc�	<g����!"O�Kf��#b�NE�w!��g�.���"Op<�Չ��fZ�}8�� '��E��"O�����(Z�8QY�mԨ��[�"O�X($CÿW�D��լY�k�j�s�"O(�X��^�p�2@Q`Z�4��,�7"O��c��9dm���C��{c�!�5"OL�"F�ӄ_Q�d�˝G�)�"O�u��)�1�Ѣ��M�0:ᡣ"O��A^�a�*}#� �*{�F�(d"O�X�/I�v�v�wO��DXlmz�"O|�)��&6b�����>���"O���#�B��C�B�!5sX��1e-D���)N�Ky�Q�p��=�bT�B�7D��bW<"�h��lϖB�&����!D�<���C8�����Z�oC��x�o D��#6bF�k�!xu��X���f�<D���B�?bec��%MXh1S�.D��@�ɂ2߼�[�#Դx&$:��,D��x1�QDz��w��q $TB�*=D��A. �^Y�iX$�08:i�d;D�pa"$�����L�>6��8Ղ:D��3�J�o��xal��xT��SH:D��1	��e?RX�-�
'[D|�6D��ٰ(������!!n�3��7D��ӫ��t���w�/>�.��E@4D��t��3,��Гu��r
�A��J-D��ABKJ� ���a�/V	hg��z�"-D���� �`p�Y�*�R�`!X@*O��Z�	�,lF\  �F4;��"O�lVD�6x�0�D�S�����"Op�d��?L�|�8�$�[�^�[@"Ou����|8N�S�B�$m�Z`�S"O^ ����$l�c�A�#v�F�"OLL�ȗ.jjH��֠��l�"OX;��g�	��L2W�@	� "O�sVM',��9r����0ISU"O�Xk��mh��P%��7O��xv"Or4��ɟrd�xFΒ:p�@8�"O$pc���%-LL]ÇnٺE��LCB"O�]Ȅə"�*���ˉ�:/�#"O��`� �b������&�	�a"O�8aԯ�<F��넥�&v�\�d"OL��0m�)vB��gĂ�jr�%j6"O����P�C���BP?=q6|��"O*�j��˝@.�i�9+S�< �"O~���j����2ɕ�_k@`�"O�@R�j�hS�Žd_��"O����8?��ӂ�]��3�"O��)�/�'�#�ZPQ�P�G"O�xt��ۀ�Ѭ~�s"OL�#cl�?2ւ�!`�p�"O�*�HP [�<��c!֍k��1Ƞ"OJݨ���8�A�_�d|�W"ON\r�E��Mx���&�ƿ�
ݭk�<ёg�=\�����/���b�m�<� �m�ȱLI�k�1����!�$̤zK�l��DˏDCc��8�!���(�XcR\r��P�>�l��80n��Ekڅ0.��rn� �̆�
$�h����^ڂ����/zr��ȓ(��E�U�	 z��w��!&)��\��9�HgŸ+0&�}r>��"O� 4�k�㚳��d�f�J�cHbf"O����лw��g��!p���E"O�S`aE�4~4�xBmǩr����"O�Ͱ֌V�r��Z.�b�#�"O�PS�6 ҈�0׫�C��Mj�"Oz��Ɗ�N��B�K��/�H�	�"O��x�a�`�BLs�K�|+�jE"ORD9'��K^�T�ܞo!�(�"O��Qӎ̋Z�0<C���h ؆"O� Tcı�V�y%D	��UH`"O�(�&�
K�BD��Âv��Q�"O�p�"�#$�`�%@����"O�]x��W��8`+B�z����"O<9ס� /��yA�
Is(�
"O �h���zb� P��l�U��"O~�y7 ÌeM�L+ BڭwN0$s�"O\]�3�*Y^t�j�!c:N12�"O.)w���l��Ȥ��y!
��G"OL�Iv�@D->t�O�.���"O�k$�
P���	�=�N�"O���F��J¬������T"O��@v����@j�
 �Z���"O��ɳ�ƚ#ux=�s��>m��D�"Opa��l!2�$��d8B�Fy��"OPY�S�1�M)��[��@�"Ol] A����U���O�tm��"O�����Q�:%�%���A%�~]��'�T�G���"���
P�HN��hh�'z�MC��8$+��^-v�j9�
�'���cA��`
4@���s��y�'�����Iڮ5�Rd��bAx���'�P�$#ض@]�,�6��*�S�'�ɒ!��E���.���B0y�'��Q#GF�´�1�˕�4q�
�'n�5IS�F�8��e���׮��S�'�6�
A(�3*S|�ЩSv�ι��'0��YGo̲�¼� G۷|}-0�'��tz�F6?���p �ձv�qy�'�\����_�be`�A
�?o#����'er��1 ��m�\�j��دE��i�'َ�@���Q}�����D"j|��'�*5�"V��YsAǈ����"�'р5�t�Y�Xx�Ɂ��JD��	�'�-��) 1S�d��a��n�z���'�����)'��1Qu�ڞf;~u3�'����+ă"%��5nP�W��E{�'����r,s.��E��*N]��H�'�,�g.��Ew�4�/��1�'W����J(3�����&w�+�'�Ll�%���� Hx��<aN�{
�')�Aq�a�(��d�2	��K���'`f�9e��6�B�+�֜���	�'��(��Lۄ ��΋>w����'�>���N+S'pѣ�V�m��L9�'�h骦��g���hȾ[&�P(�'��X7B�+�G�]�6��''
�5o�*���kd��T���'X`�p+_�yf�`��/IF�%�'}��@��B+�0���I]���'(A��eO+
k�q�@ K��D���'���6��T`~��d���R��
�'��:d��n�<=��b�~`�	�'�t�ʓ�����`�EN�	�iQ	�'�fT��O>(�h���� Jz�	��� Z��c(��+eȑb�*�v��"O2��-�$8jq���'g�b��"O�
��V�M�~�swH�XZU��"OB���&k|��s'TsQf� D"O�K���`�Ф�0F�8{�"Oд��C�&*�5��c�'BR�e"Ond�U�$�̣fa�8�A��"Of�
5C�*o���q�M�Q��"O܋��X��(2�T$IB%��"OT��0*��2��@����-�F"OpI�����+���!��EIc"Or`�Ю�eo���D�K�A�@	
�"OLM)'�̯V���+�8�,�"O��@D,�r���A!�Fs{h��"O�y8dN�6M�õ�����X�"Oj�f�+E���4EA�7�H@�"O6X�Q�V)�=���F	[����"Oʡ��G�6�r�"$ҙ:����d"O ��U�;c�H��"o)|�,�q�"OZ����J�H�o�N���@�"O�P���{'�1�7O�9����"O���d#��~�!�-ݩC*��A"O�	Q���.@S~�i�i�6[�u�2"O�x�Ab�M�D�)
#�A�s"O�����A�]�� IB�ڋ�jɛa"O�0�\J�}��B[�5t�fL[�y���UAT�)�AKFU�`K��y2�H�%u�/FH`+g:�yb����@d�W�oEF�aS���ya

G4h1T�jE������y�-P/�|,��@�y�<{�����yr�UAzr���\�����yR�L0[��+��"<�������yҍ�[td����#����͸�yC�|k��S)�{�"�""G��y��+y���1,H�JD�� ����y���VV��S�)��.͸�{【��y�A9::Ȑ�B�Z�8c����y��ݝ+�|I�.�U Ei����y���{���x%ر[hU��
�y���_i �CЋ���
C�ݣ�yj�>e��Y�AHQ�ȹ�l��y2ȃ	}��ȇ �SR:��g�ؠ�y�A4]<@�w�.P-�����Y��yb�^�V�6p0���.X$ZA�B�yb�]�Z)h�4n�W����g]��yR��b�ZD`cFY�N��H�I[�y�On�����t댌3��&�y�,�2=3P�ӣ���j�Ȅ[�j�8�yb�;x=�E�E/gt)�\6�y"�P.v�93.ԉZۉ�y2�ծu�JEb2i�3/�dX�lG��y��"�`�AD��74n����	��y�	��|� ��G��=�$��nû�y��1�N(�$�-2��<+4����y���M�Z k�k*" ,K��ۛ�y���3����J�.e�$ӑH�>�y2�S2� ��*ؑpAX���N�y2�B�GW�9��NF*Y�d���-Ʉ�y2��UE,�Qu�"J'^��E!��y�K�t�P�
�L�'H�� ���P��y�҃{U���a
"<��y�Q�]�y"��	�C��;l�`� ����C��������J#�@��#�a(�T��S�? ��x@���O�v�iv�K=JuB�c�"Or��OW�;l�A��)D�h��"O^����#ANd�@'VD(
l��"O,��Uo��8����([�:	r���"O� 6�'�^a��G^eJnP��"Ox��b��	9M��0�ES(��"O8����Z�%$��vDαj���R"Oƥ�'�<������@�,7N  �"O�MK$�����[bm�
�!k�"Oҵ8�.m|1SB�H�*��p�"O�8G!&����I7;"�ag"OxQ��79�
u
A\�숡"O�Vj
�}&�k@�Y0$�}#�"O����FW�E�9I�̾j]��f"Or<9G)C 3Sk�xV�ҥ"O �!&�J��"�j :��8:�"O �c���j	�tÄiW�w��;"O�@JW�@q8n��A��LP$"O�\��	�9�ҩx&/��k�v<C�"O>`8a遌Ee�� G}�<�$"O��k���	����.�{��4"Ol̢�M��sn]��O]8)r���"OR���nI+M�r��a+�l �"OnL�W���! �0`���Dm8�"OT�`�,Զ�F��$��.�����"O�U��E�`���J���'�r�e"O�U{W�N�9)5X
�� �F�"O(�����	�H��.��_��Y2�"OFQ�Dn�fE&�.S�p�`"Op�0��I���;�C��+v��`"O�&Z!uI�Yfc��f��"d"OĠ���0$누�"��;ZF�"O�L��Q.#���׫ ;�~�c�"OL�����d�f��jٲkv�͈"ON4��&»LR�9ŊI�7����"O�	T�f�e���_��"O,P���+t,A�G�B����"O<-����X���Ԡ��Z�04�1"O~��c�J�p�ĸm�v����?D�bM7/�1se�h�|�JFM7D���ȁva�@8w�\�3�Qs�O5D�8�O<��)x3���ax<U�H3D�`
H�! ��a
�v��|��E4D�hZ�@ߞ]��Y��A�^~��8D�3D�|��#T6�&���o�
Hi��J0!2D�8�vo�9�42����GNu)2l"D��q�ЇC���z�/E*�q�$4D��j"i�hD!j�@O;
X�iы1D��Pt
��q�����䒶N3�86�.D�`�Eo��)�&4
�H�����J�f,D��(g'�/���:sO�8���Z5,.D�܁E�W?"qr���7��U�#�-D�x3U�n@p�+C���f\��sV�0D��kR�I�����F/)��i�U�#D���q�V�T���q��9ڦ�� )7D�|����A�T�؄4(<i�!7D��;���iC�\hd�חO � O4D��c;�r̃�B60B2A��6D�$*��j��(5���1��&D��Ȧ	�4�b(�-@}�!�2�:D���AN��D\0��N��o�,���9D��bG$�.*[���t��G_X����7D���G!Pgv��3��ٱ ��X��(D��H-��Ha"�r�
�=�E��`%D�� �Iqdфo}��sI��n��F"OR���k��y�*劦���(Y:h[�"Ox�I��F�;��p갯ٙ#<
́�"O<�ᆅR�3I i��k�5:4$e"O��E�\�W�:ux7�:V0���"O�5#D�3p?D�#	0g7ʸ�"O��Zr�X�;�H��R��9UW<��a"O:48�؀l�6��GRH���"O"����Ǝ|������UM���"O�}`��	r�L�p��NQ���p"OX���@����@�q��Lؽ�"OLY��Ϟ��9�	��9�De��"O0�lOE��0̲�K� �)�P"O(���"�B�^�W��	�XA$"O��1�N�
@��p���4\�"O\  SFW=M�Ь�5E��D�P"O.b��ܨZ���D�#w2-zW"OT�k���=y;Xir��)�R�"O��S� MQ���@v/�"D �#"O��鑁>^���ç�9�����"OX�JԠ3���bc�ƕtLx��"O�Lx$#�0+j�@&�>*h<Q��"O�,��XnU�u�0`��Y"O��j[����!�oE7΄5"O�Cb�'i�x8@�FD�@��"OB��T���\�cf���:(H|�F"Od��N�#Dc�)b��#%"r���"O�bg!Cm������_����"O�l0�ϐ?�Ų�`�*g�X#c"O:=�`�&<g(�;�o��f�"O��33ŁXS���\�i�bp��"Obp�Ф�E�μa��¦K=�ɕ"O^Ix�J�;��85��U�@"O�:���)��H�A�|aj�X�"O� ၦˆ;��b�7V|0(�"O�̲�뙔p�Xt��m�5T�|J�"O��)˗z��I�f��0;��"Ot�yA��g��lp ��Qİ�"O$�p��	l��p��-td!@"O�%@¨�i��(��l]f�V�g"O�y��B�[��ؖ�R(딩��"O���̝Fs��KsDݑP{�yb"On�`boD+ ��]��b�;]�dPV"OF��$��3��-(ԁ�5�H��#"O���o@=���S��*0�^��''.]�fFX�E�q��'>08��	�'��٠�bf y�%�"EW���	�'�t���-;"b,��b��=���	�'�4Ѓ��[$<����ӡC;���"�'G^�IGlCF�[!��$%B "O�y釣�������R�RTc�"O�� �*`a�d��G��z)5�B�<���	0���c��?#S�h�%�|�<�2#��A
U�aJ�MXh|����q�<�C���y�|���	56N0�4�b�<��lA$f7D�c`�H���`�U�<y`�A�a�j1���gP�Q
�M�<i�G�,X����BF�)�~Y���.T���(�-
B�]t����g^C�ɍ|:ıq� �ZԔ�B�kް0\C�I�jI 5���њl�V���P*Q..C�I6|�Bd��g��$T�"��
�e� C�ɰUj�m�e���&��K�B
1D�D��e�����Ƃ�v��ǥ.D�� Vt����KIz�y��?�1x�"O� &���>�������l��8"O\�Q6�/! �����2WW��"O�AB��'h�1�D�5h���"O�m91)O�����.��{yl�5"Ox��Dn��;=B,9���*#G�hb�"OI 5�*}�� c�Ms)6L3�"O��S�aM	�^��(|r�Q�%"O��e��}����ȹ,b����"Od�X��=��qH7���&"O\l���3<�L�Z!X�_����"O���"�n=C��^4bfda�Q"O[�	�,3��e���ÔU�h� "O�$`R�I�{yrPC-�`;Rqӑ"O����"d�&�H4�M;i �M��"OR��F��]y��)�ɮ!�R�+v"O��" �V�l�@��#(����"OF��#!�&R�v,�%Oōd��Ca"O:����H�r5Z	�'Z�j�yQ"O��� S�C����LH�8E��"Op0�̓�n��h��)F֒��"O���F�T-N�@��NJ�&!� e"O&�3q�X&TW�	Ҁc�%y��	�"O��	GGգ�F�MI�_sN,��"O$��D��9	���󭟾c�9A"Oƌ��j#B�A�G�EY,���"O�в�,��+�=*�eof���2"O�R�.x�@p�Sr>�Q7"O�*�kK#hM*`!v#�v�De�"O���5��j�j��2aH�H�;�"OL���Q��v�����E�����"O\%�j�1 稕xe��Q��5Bc"O�h�̏�r�f�2B'ܬp��w"Ot�z��(�+mޚs͘��ӏg�<	��'S�����M�Pd~��3e�i�<�֪ț�Y���ۅtK���e�e�<q!��p"x�PG�1��h�#a�<9 ď�@���Ss�[�yJt9�6 �S�<��ϝ�m�<@
U�V n�M��b�h�<	��W9l��a@�Tm��2p+Ic�<9�BڌW��(�@%��qd\16#�S�<Y�"�;[L�œ����ԁw� {�<1����Y�P�Of٬��6v�<ʇ�x	������h�v�Co�<ɑDM��X�&��"<l�ԏUl�<�G��k�4�J��P�Q�<QWɐ��n�����'�dd�SDR�<	�f�"W7H�C���5���X6��J�<i�!F����^$��t���D�<Ib�׺b���"�k"|"�5�w�XH�<� �F>t(��u��'�2)SCZA�<�wk��X��1��W�F�l�c�h�<ISLK7Mr��׊�D��1&^a�<��՘(�u�u��;xƴ�&kZ_�<)���5e�ԭȑ�jɻ�+�t�<y�&��y�8`"a�^'�p#��p�<�Jҷ�+�!Qw}��q�e�k�<��/!D,{���s�$�)5fh�<9���$>3҄E$`6� ��ɕI�<�2�D�h�ٶ�V]_��C�<��!`a��kfϷf;֭@��A�<��Ȓ�Kb��f刴%�6q8�	y�<)����t�Z����1�������\�<��hK&��k�i3&H������y
� ��z�j��T��G�6>�-"Oq@H��oȚ��L��>~x�"O�ئ`	�AM��p�A�U��r"Ob�f��YI�L�/��]F��Е"O�\��#�&D&�����0fZ-Q�"OVA`�B�k�t��@Md`�"O<�0&b��F��q�ƛ
�桓Q"Oj(q�Q%��I(֥�/>�!)G"O6 13eՋD����2���L}\�3"O�u�Uc��8������-j�D�f"OF�a�; �`�!Q��]��,Js"O&��.�Z�4IWk�j�0U�w"O�qQ'K�5Jw��R�_�UKD���"O�=�� -bgf�(��@ CV�R�"ODY�AI�$��t�k֊W����A"O�	I��Q�Ԁj�k�
RO$YX&"Oؙ�5@�ac������!Jg"O��Q ,�L���Ҷ�P$}�N|�"O~�:c�H�#�DBW/�W�,t��"O�u"�ɢ)S���0oC���L��"O�e���	3���b��N� �:"O�@9�&\�Z Q��C�b�0"Oh�
���jL���� �v�
t"OD���H� 6�!Q��`��q��"O(A�.�e�$�"QJ֕���ɠ"O|���gָd�>x�A'� o��s"OЕ�򂙋"P*�K���Q��1"O|�p2�Q���N�V�0Q5� D��:�X^��9� ÖL��|q��>D�
�C�0 2&_5S�� a�7D���$��\۠ձ�;B�\��6D�������|�\8\%����/D���t�Ҵ"0�)iV%��x���),D����Z;E���؄�Wo�θbbc+D��"���������*��hצ)D�,��%�4�`�N�G��8f�3D���a(�:ю�ԡB<�Y�C�%D��ؗ/\�As�� �.C�����#D� ������ƹ�� T�l�"��!D�[re���(:t'�C�.Q)bn$D��%��8hXw�G�5�ZɈ�%?D����s�E� I9"v`�@$3D�����Q>��4)Qd8��Df/D�x{���U�����(�ڇJ#D����K¾A��|��R�Y6����?D�$�����Y�z8bP*C%"=H�"?D�dЩ�P3DlK��B&O�>m���?D��b@�J9r"D�H�$�Z��F�)D�4c��5%�6�����Р�"D�����AQ��y���`��8B�!D�XrkU�^$r	�f�n���K\�!��w���O�"�  �V��!N'!��U!�|rA�& ��0[��G!3�!�$�7"h���h����P䋄'�!�$ԀJ���¢Y�k�, s�S�)�!�C-��4�v眞��(�1c�uR!�$�l��d;B��g"0���b�!�ߌ{P���B�u�\�w��%�!򤌓j���瀋�\�b ��Q�!�d�W��p@�"���H�.S�>p!��>���0h[�M�rQh �@�R�!�P1-�T
UȔ�8I��܀�!򤏇z*���ɵ1���rC���'�!��h�4��SL�0����	�!�� ��	%��J�4|��L
%���@"O <aF�1j}�\H�H6�J�Q�"OLDN֤�p1�dCЌr�ؙ�"O&��EU���	6�$@c�hR#"O�R�Hӓ*�8������/G��"Ov��Ĺ�<�C�I�.`eJ4Xb"O`��V���E� ���yN:�;�"O��
ScQ�n�^!ahčFH�p�"O~k�HYT��e��g�7i7���"O�t�' �!R`���.��"O�����s��Q�R��a�0�"O��#�$������41����"O��&���L�h��臓z$��l"O���*�={5đ�(�8O
D��'"O�u�*L�T��-�!^d���"O��h�"ǌLSZ�h4����BL��"O�1�u�O���i�:���q"Onp�G"@(wt��ʚe�)be"O�+�@��he�D���r{R�rD"OLpR)����%�6�Ǐ-��"O�e�ՎB �$�pF�%rv8b"O�xKv"޺F!j`�WEƶ%�
#"O�2m���!�I�o��,
�"O��0�NݴQZ �󁂾N鲘��"O���S��5J��w*�T��"Or���f�J��-�� �*�b��$"O�D#��*y�z4��g�&�Y�"On�wX�1��8�$ȉA��"O��bDd	�L�j��P#:��{�"O���B�WS����7`�eF�,q�"O(�IÏ߄S��� ���]E�l�f"O�:��[�H��i�2
L$��"O>����;nQ��0 ���i�"O�=�S��~E�B"h�2w�.8�""O�9*T���`G�z�P�5"O������<"� �۵/�[�(��7"Ohx��W��(�O�5y���`"O��B�&����J�N�Eh<]��"OHm���.�,)� ˆ@h�4��"O���쉹q7p���MK���"Op�"�)�8S^�8k�"O�_\h��"O�\[D��J%8 ��M_���"O�T	r��G���V�GP���.�y�߶,Ft�K
�*�lxJ%�Z�y��^�1{9+��ޖo���q�J���y2�߳6�Y�  ��j�ިk!�E�y��)��;T̀�c$�UY���+�y��H��C���\��t�P��y�	S�w���E'=1�e��l׌�y��F1#dX�^<�h�4 ���y�D۱.g�I�@<G��{d�>�yҪ��fYC�B3�M�/ϣ�y�+N�a�|Qɰ�M�	'X� ����yR���z�j��pkØ@� �R�8�y��I-+�Ȭӂ㓣~Y��J����y��͂q0����sn�A:Q��y��H�Z)� `�݊A��p�A��y��Ʊ'a��iV89�)��yb�@L5�u�qΕ�t@��Q��J��y�֩E�(����ړV$"�`X�r%��T,�S�Z]�7��?8� ��\��,�oV�	Q��ѥ�ˤ�p|��:�(5O.yJ�eJ���:���Aq���듰
�>�i`4[Wnh��S�? ���jݧw^��)T�O4\�N���"O��뒂�'u������X��y�u"O̠1%/V
+��x�8C��"O�|��ćn4���5hW�%�,La"OH�iQ�
(��2��d����"O�� po94�Z5@*Օy�� I@"OXi�W�B�/���*vhHr�2�"O�իuT�G�tUG�<�m�"O&;�%�>��9{T��Q�����"OL<�ES=����%@�\����"O
�;��׶:���{��Y�?�r9*�"O I��H!I��S�R-_����"O��b�JH1U�ܺ��z�m�"O���7fO8XT�ʄ��(}fn)��"O�	���7iB���厓c���@"O0Đ�[�q����F!70޸�f"O�����ͱ�tySZ�D+���"O,�37�WEL��b�'+�9@�"OvPuڳ�.-s0#ͺ;���W"O���r M�,��u�G瑮����"O�]PNȳ[�4!�")5�j1�5"O~E�u��2�0) H�
d� D@�"O, c�/�ž��W�����[v"O��p��R�$�J�9�	 *m��"O�ɑ�
=0��d�2;��-8��T�<9��Fjp��J��4 >���g��w�<tʏh���BEL��иK�d�u�<�Đ$>�l!;*6qδ�����L�<yD${�:q��g�
9Wb�qԧZL�<	i����DH܅}�X�;��^�<�!��-�E�A�Y����p�<���;i�i��FXİp�C�Yh�<�D,è����`��7��ЯJk�<��,ųH�l9xd�#{kQ�+i�<y�)R7�:p�g���꤀�GNh�<irh�0 	z�Kg��S���$�Jd�<��i�'t��]�Q j9�Pئ��u�<�����v�����=hk6�Lp�<����u�,A2H�O�ƴ���[m�<�0�	�@q&��t.�c��Q@�<Y4)M�U{��Ruh��W����F�<��#�(_���P��Ld�-���AF�<QO��(i�uA0�W�3<Tyש|�<	��5x 1a�1~�n��v�<�⭋�3f� 9��(Elܸ�`Qs�<!q����NB!G����Ru�<�� ��\R�JB �%;Z]�D�n�<9vȌT�@�	���!V�$��n�<i#���?�LX���5*8ph �ej�<qg��:D� 1��0������i�<ѧ#fi�lx��f�h� ! 	z�<���"}���hT4~vB�<a�ȓ+��jª���	0B�ȳh�0���f0�SKF��N�  @47�r��'��	q&���!ٌ�1'������'�V���"R�8�.A2փHm��D8
�'���(7�Z+7/ܜ�$'�n��	�'PD�Dmɾ?{��g��7M�Bh�ȓJU��@�S�6�RG�:s=�D�ȓ Z$р�,B)b�.���n�`�숅�bY�0�f
ejv��1g[ a��+d��S��Q`��T�eML �ȓT}��� �B��0��<�ȓkk�$��.��b��!�ҁγb✅�S�? F]�Ň�H����/,�<���"OV�"�;��68X ���"O<�0�O�J���B!��.9�ЍRQ"Ox��eh�{�Z�b� ȶp ���"OD(���HAdZ�����X���"OzA�W��'�09�.� 
�	�E"O���� �0��a#+��ޭ��"O0����Z��ua �S�Y�h܈T"O���G�:i��3�P��9p�"O����Ba.H�'X�U����"O�-r�I�z���&�4���0�"O�(B�܍e��D,q�U�d�Ҏ�y���LD�d�O!YƼ��A�-�y���'/.pc$IA�O�fT(��H�yB�Q� vP��ĞU�\�{#�\�yBが@��Q�΍S�=�C-٣�y��
\�^�їg9a
���"��,�yb�"K�.��q	9�8���G�yb�� [����D~�*�)��H��y��(>��� �C9g��Bv���yb�* ?Nb���)b@T��&k���y`H�O��p΄�\�eȆ#ݼ�y��'R,�#�(��HmJ0��[��y�o>π@���K�COفf���y�Kܖ3|��%P"U�����yBHɫjTBX��'ž��}�7" ��y�ɞ1H�W�AP�6%�GK1�y�*	�4�8E	�hYT>�JעA��yb�.ܠ��f��4O�@���B)�y��2�J���b[-��Rf���y"��k`8��"J��H��@Q)��y���F��d��M�jwz����y�C�$�\05�����4&�$K
C�ɇ��A�pW$��eA]�x��C�I4*�PU{��Rl�}R䭍�t 6B䉀�X�B�BB1V�Ŋt�-;DtB�Ife����(o�<����LJHB�	J(δQ#Ĳa� 9æmD>!�&B�	 W5�|#��� I����C�ynB�f�~�d읱I��hb���C��<"��(6h���I��X�U|C�I�N�<8[W��>j`n	��*_|�B�	F�,�J����pf`�R����F�`B�	�e�b�#�#,sFmke���zB�I.&Ȑq�eN2S��<��M�!jjB䉻o��Z���l�� ��s�VB�ɭrW~!2ǉ�x�԰��N��z�FB�I\Ќ�"_;%^ �Ƈ?1"B䉓���cD�ѩ?@�X�O�=�BB�	;�ҥ�P �
\���v���JC��o.!�"�	 B�G�/�!��'{����g�/I�ٲ��љjc!�>��82CO��2䒴R�D�Q�!�d�&��)tAM�e�~+��X�$�!�D�	FЁ�f� %��9�E��$�!�$N/K\pA1��<B�J�1"%��!��ME��A�D$�"�Y'�Ͽ{#!�$�(k-���COQ.��9f��Ru!�d��m���"a�M2q�`}Y���*[!�DOL��
��@���|r�!��2M!��=p�|]�4\�Jiv�׼K!��ЋO�xq���	%z��(�FD�!���	A� agCE����b吾�!�ĉ�j4@�3L�X���k�P�%�!�� �(�tI�c���W#
t*̹�"OZ�ʓ�Q�?!�=�D��jQ�I��"OR-jQ(�'Q��5�e��3C2��"O��V晿xw@����7=$}�"Ox@����El�ȥ��q0NA[s"O�0��PT�1����Z�"O�I{�e�B����W_�>���v"O���t�SY�J�,γL��sZ�(G{�����u�സE�Lf��mz�ȴ"�!�d:r&�d�E[ ��m���%�!���/�D����ܢU���ꀀ�
-�a{���-U8��!��7,tɗi#�!�Ą�?(����#q@,9�6)��eɱO�M�����KN2Eh'\dsS�ԇ�y�b�ǚ�C$��?$�2H�bN�<��D7�O���f��u?I��,L?x;bu� �'�,0ϓ��'��'�J�K�H�&���-OB�i
�k��X"�M�+t5���Po�ن�I%k����!��r��S*�mS��`�Læ!l�o؟$�'�Й1J���s�L�p�jyӕl ��ȟ�)�WFW}��t
��J�����'��f�\sQÔ�$�
��P+F�d����OFX��	�A�S�OH���t��:���5�۳=�N��'ٌ�`Uɖ8 �A�U(��D��BO�L��	� �0(sw�ՙ8�*Dh��ѽH+�6m5�S�Ow�l�@� "FJ!j4l&�{%��:!��VOx=�Ջ��).Ա�(Y�.D�5��'@��DD ��WDS-�$�
�'�� +�Y�t�1��u�HI�C�'����L�Wɧ��J�S�
�3X��'<GΡ�"O��SwE�S�4�4�	�Le$�1"OHtj��A �qv���#]�}�&�i�X�9�����7�Mc�4vz�sP�ȁNn�\#��Tq����'LD�4A�<��@�5N������O�	��I�2��Y��kE
s�CK^�Nx��d�O��'�$5�����Ix��H�v��)��OԢ=E��fY�{V�fȱMF@Gh��y�Ɯ����4�	F�@�1���4�y/=I0*��L3�x�Ҷ�8�Mӌ{b�O?7m�UI���G��ya�E���=p�!�D� *~�k��i&ʥ��!��{J����e�%�P�J:�a}�W�8S����`)�`rfJ*]Q�l�㨑�y�V�^�T�qr�A�b<i`G3��O����i""d}���Y�Y���b͗d�!���(�@�'�
8�(��4H4�L\�<�*�L[�vl���R�D �uG�h�<����""�ҍ���"O�Y�1#禑�<A�Oq��-�	p��
O�T+3\�
��I[�'��c��ϮF��i(�	7W����}b�'�4�*�-�V�Z�H���Y�@$q
�'g�Q�LU�]kޤ���'N(���b�N����&�V �([�Z�@j0O�LY!�$V,6�!3�F3=���U-�#l_!��;[��rԁDN���Xg݌����A@�Z�O�I{�l܇9� k�R�E)��'��E �΄p����
,i�
�'^��x �D3[��tH�O��L@�
�'W��z6O33�H�����.<��'qaB�v�����;,hqЀW���>1�`�>ٰHV4H����E��ӈH��BX|�<�ӋC)Ztt���f��X��DRv�<q�h] �a`EI\�����O�J�<YDA�W �k�$�q����� �B�'��y
� ���``YD���u`�&��P�r"O ����M�!3AF<"�|��""O�iS4�܏l�B����D�r��p7?O�Ot�S�g~ۜ@�5�4OQ&#�e�2[��y����ҕ��l��ԉq	����p>�t��gN�a�AƉz��I��	m؟(��'��z��\��ժ�'@���#�'!�4@��I�F^콱�T�5��}���DR�OӠ��ϕ�;1Y�HY��S�':�ĩuR���k�|�25Y�'�Q�4D�DB��@� 6�_������yb�̘h=�p{'��*M��CWΌ��y2n�*��j@��v�<�s�"���y�� �~���0)T�<���FM��y��u^"Y{�`�>.�di�B�>��I���矄X�"Mp��()/fLI#͓�y�T�03"U2�aל$�~�RhZ��~b�)ڧT���Kݮx��P�@�mY������}24�S> {�ݰ	Y�"`���ȓ3��l
�M�'��M:ƅ�J���Ez��~2���6��_%~�.I�p(U�<�c�<�DYQ���D�@�H��e^7xb��QA�	k�!�ʹZ4�4��,g\���IҺZ!�Rv�p`:7G^ J>(��B�p��>�����3� ��ˆ�:�N��#)�đ�ȓ~$�[�W<U!�()�)^��H��+��?!�K�.�&�An�N@T3�k�'�qO�Q%>�PŗV�����R	��a�  3D�*%*�1A��r��C�V��=)��.�@�?��{��$	�()a�]kŌ������yb�π5�����1u�Y�T���0=��3>ьZV#�9i��т˫�ye�%p�!@@&�h	y��I*�yb�
.N"��90�CX�Ȓ7����yb��65����M��Bຠ�����y"lJ�q�4�s.D�-ӺpC�L�yb ��{2��K��,��Z6���y��c��QГ�J1T�0�*
�v#�5�(�ɧ����$�h�! P�� /�2�̝.�!�
�mE��Q�d@���h�p����!��9D�l�K��Ae�v���NI�!�D/}?��3"�\)J���"�`C����'% ���C<W�<�����u �4��}2�>�����ٓ��D�9UQ�[�!�d:q��c��T*��!Ad�2inўX�ᓶ(9<<ᅍF5iS��0�!H"�ޓO8��� 93\���b�V�Ҍy��'&a|��/Pz��iC�U����q�l��y��`�X��)A6~#�̪�	@
�yk�Pu��A~V�� U�ۗ�0<1��$� 6���V�ٜ@=!Z��-5g!�D� ���w�ß.*��R"ީ=�az��$R&0�ؕ:�
�.-5쀑���X�*C�	�N|�m�vO��<p`��*vV�8�D,?E���_���@��%(�A#C�ܣ}r!�d�TFR}��fш1�!��ŴJ1O!Y
�
�U1p
K-�z����O��ȓC�2�1Ɇ>�R 	
�\�
�ȓgL��X炜�tn����B�l�E�>I�{��
dN��O��
 �@��/ B�!򄟓=nkf̬,�]��ܸx��d0�S�O-��B� ߣ_B��w��l��P��'��$P
��h膌�iƽS�O�ԅ�I�H�t�v�8���)������>� (��d��@`�4�;S�P�Z!"O���r��6_�$�nǹL�e"a"O�1���D5=�(Q­O�B�Lk�"OFhB�[f���ѫǒN?BcF�'��Z��a�kǠ�(2*܈�R�ȓP��}�`f� 3�LQ�qJ݄}����>�y{t+�fвխ]7���4��{0JJW/�!�3.ĳU��p�ȓb �U��0(RuP�*�T_����{y�4@e
�+F�.��3i e����=`Zd��/=���"%OX(��V��=�`��E�M�b�޾T�ȓ0R�X��ذ@��pRw�S${}��ȓT L�2(Q<<���ʧ�(�ȓ	����2��9�(��� ɠVrq�ȓ8и`�F�1+̆
W��Q�$D��#I~(`���@�iHb�i +"D�<H��&6�����2�$y�$D�t���D�L�!ڧ��b�� �&D�����d�X����O�J��;5�#D����_!L�дk�3+&Qc�k#D���f�
(*���B-Q�(t�@ר;D��4�2g*�u/��>f@�$,d!��>$����K�6z�`T L�xc!�dR�/�~\8ׄ����1w�E!�DЏ?"����T�9��ë5!�W:.���Xꎛ=l�DP�mR3v�!�$��)@��U�Nt��e{�ʝ3�!�H�`h;4
��p��M��*'x�!���	�\��S�o�P��_J!�
˞�S��׶q��HڒO׳�!�Ć�(�&���1l\�8���il!�ě� ��X����@��&��Jh!��	Or�#̘�hWr@8���7 �!��Rs��6���*6��'+�<�!�I�Q~
`zԍ�	��p�Q/�8&!�[�����k�X
t�����u!��..�ˣn	�t�:���R�6A!�C�mHdT⢧	6 ��H���|�!���t�$|�E.N
.�j�[Bm��$�@�8��[����rL9"�az$�?7NN,
Ŏ� ���"�y"�¯̔|�coԝV_�Q����y���`�Bi���I�ށ1T ��y��a¹����sd4�3ԣ۫�yR���uR@�P�f��쾙�L1�y�jõKB4�:�e|��%�Sc��y�E�"F�1�cJ�N��8�
W1�y��b�T��C#8'@��H���yrԢA���[�N��g�h�"��B�y2�E?(�܈g��[��<BCÊ��y���	"{� �E� V�E!�k�8�y�*�����N�4OС��M��y"�I�>�̙��=<q ]�[��y�\s�}K�Fޝ(Z��b#l��y��� EG�`�g�A�C�0AZ	q�C��n����S���2gG���C�	#\��q�%g�5"�l�OQ5D&�C�	��*��s��򘁚s"DC�	/. �c2(���8�Q�/�*C�	�n�Ve����d�$a�%�?�ZB�I�KQ0uXă�n�B@�0g���B�	+ȼ堳.JJ�4���Ő9����;馰��{���[�HW�Q'���R�A�.�*"O�tj�IZ\�:�`;hs�(*��O����B!�I��S�? ���2�u]�M�r�W%%E��u�'\�E�R�ץ$A��%K��.�,�E�ȴJ�6���pi�Q�+4�+3`[�H��<D��%
�܂��>}"� �J��5�]�abp�F��F���&e!��pH�����7h�:A�"O(�*8
ɞ�Z���!���$� H�r����FN�
q�ȜoD1��&�pC"	ؕ��q@3��MY�9�f)�O�x[b�6�PH�A�N3?.���,�mD@Y��������C:�P�V�'���cJ��a�F
�Z�P����3&�B��+�,0U"'|���A���eؚ�hO:*�Sc�J�ʹ�+q��mx��0���#���q0�=F�^]��ʪ>Y���d��V�CP\~�1 �EQ��4����#i�*\H�O���7����:�U| ��
�S�Z-�!��)��	�(�r,�c�HɈ�+�d��&���I�gS)7�@!��غtEj��[_��e3a���!�H�mFd!��5N���{%f�<���ڇh-�I�z�H�[�F��e���0)���'Eh��P�Ϳnx`}�@O�$��i9��Ԥk�Ի6�W4�py�AO�'�@QB�ƌ<huvU��/7�	�{$ᐐ`�+S��吷��S3Dd�G�R�x�
%�ُ{�:�d�M�ԣB�X�V�+V߸l�\�ha�_�J~섲���:o���e�W���(ya�O*_�J��V�M Y�a{��,'Ox=���]��(���_	Er�B�D:?�qmZ�v�Ca(��\@���Ƹ(/�q�%:�K�%<$��,�P�5�6��9�~�ϓS�-Ҷ��;�p<��c�����z����!EB(A,Ј �O�Q]��W*�U6�j��R��p�Ex�����	�� �.8�R]�S��D��\!���v1.��E�Nd�'�fL8����΅�7�ד-�(1P.�3��I���{�r�iԈ��q���4-ų0Ҡp�(�E�:����J�F 3�MK�!���9t�ҍt� ���}�BD��d��,5[!�����'b'R4��k2m�j`�ՂZ�-�MrƲ�~̲A,���|�����9e���(�솊�^X�."2w��hQ,��Yٚ��wIDR��	b'���0=�bםY��q��K�)s����#�l��u�_�,����[�D<�2B���X��Y���	+t��)�DR�%�z��E� ��a�Qm�*1q�y� �߰<A��Qh�ċT�
��hR%.qE�iؘ`6��E��K�2y��'P4Z����
&V���t�$+~
]�%)��4� ���I�8a��U�k,�K $uY��0��Y��H贴;2!	�"�6��0���tb��n
�#���'
�9�H׋{���T�=Cl��%a�G�`��7�_N�h̋���	[!�(�y���}�M�4+|쵙D",�l��]L-�v��8��P×bДh�\�j�i� ��IZ<��֝�Zg>���6.�" ��3-͌ɚ��UT�|������,����-�aybA�E�$��6[�źB�D���(��eʂJ�]�%�ۮ/�F��1O	R�8�d@�Yx�ْ��=������H��k�^;�����.S�^����I�yM�|�r�ӄ~�T�+�k

 �
ݱFRG�~в��U����fo|0y@��G�	�x8 ��J�c&H��G�Ǧ��);�9�4o��;E�����۷��dR�Z�4�B�k�N6�܌a�Q�� K PZX�͟�Q�RC̄Jl��cH�4r�qzT��-0�D���8��\Wj��B���'k���5�5D� 	��Q8O�^� ��[�q�D�����ԏ�ħ$(Jwi)i��1�+��T�j�L��;ǩV�9bə!!�8�@ȇ�I����`�Z�����l�������I��n�(\�Y����8z�aP�a�y���E _l����Ǽ�ȳ�C�#�xU��a�2�)��G�K�'9�0z���^X���ѡ[v���H�Z�E#Rρ���u�3f
�A#�a��ڴ#��@)&>d��9d���D�%y��bF�H���	yaR�����
+f��G%R �?�7f�"�A�����A9HE��#�*^�}Epa+Ͼ(�����H�Kj�L{Q�:X���4'���=��$��k4M�#>���4�t��GD��A�tqB��)K,v�!Cl�+C
�#T��&���D��6�|��G� �C�dU[�Q����"��)vK�\@FO=o�,�B�.�j�j��'� +���-�d�ڳ홙?��!D'F8Z/d�r��=ٚ��si�Gy|�����'�p��:��J�'��X,`�jR\�d�#/�\q�+G�3m	�+ʓ1<�|�-�RQ�5kF(5]Ys��<�th��D5j���,�D�*r$I�JHPq��u�~��bI�/!A�x��DUw�'�RY����9d(���ЫCz�R�I�n�Iڽ&�٫�4d��T�Fy����e-���p�B��@�	n�NNM��#���(
M^)o9����x<i�!�)�O�����8J��qh��Ȑ��\!��I.:��ˤJ��r��<Y��� Ϙ���̑�N��qxw����Li <��	#���TND�S�@��y�¸3��'�#��\�[E����B�o���y$�#'Th�d���%�8d��J�wB�xy�B�$H�АHR��k���)��L���qb\���5{�"5��M�� �lP�d� >=v�Gx�Ǉ�u��uP	�+j	�� BȾEtt�@W��$�j�4��): 2�M�,�Ѕy��G�@�5��"vԮ��H\�a�d�[���c�'$�չ�g�t��C��ir��"e"xqB5��<a'�Y�F�˯Q"�š�GՁq��Vbۇlx��r��}o�upG�� ��*�&X�h3E�[�ph~��A��^8�P��ft"�3#ծ��i��U�.l�x����:@�Z��نm�Lu�F�pv8�+q��.��U��u�Ŋ���.c(E�,S�ы�?�O��h^�2�vm��o&�D���S?�^���.��� �(U�,�S��Y�ؒ�ON%�B��!듌>�Z��%�/���@Hʑ@h�ͻ�O Ւps�O��Q�Q� ��j%�	��W7?H�DS�mA��L��RP�"�Ă��*�Bt���1���a�>H)DĚ�넶>�<�꟱! �b$ʓn�0[�@	.,����̇]�P�f�ϳw��(�?>��h��A�m�${7� �,*��H�_�D�!ϲ紜�ciҜnZt��E�{� ]x �(<�,����'�@�:��j��4�w�Ud��Q@�D�w������"x�Pƀ��D��)�i�2ku�<K�0�� ~�`M]����\�?�YY��'�Qy� G	<�h��=w��C�N�e���ȑ�Jc���g�;q��h��}ӰXY@,Ѣ�`kΜ�V�>\���֩!+��b�텢=��D|���X�(�{����Z��tǁ�t�@�U]<�@ȥ�-dD�ITFZ5B$�'Ɋt+���tX�b��1d�)E�ֹvԄ}��!k��(@��Wr��ٵ<�8
Q�Ԋ 4b��Oü���E�&�B�����)] H"a��.gaa�KH<�V�6g�n��cŠr��$�!͇�mϐU&m��H4VzG�	�`8�f�ضf�h���E��y�MӼ�'+��B+P8��[�D��P"�V�� 	��?\��,��oMy/�qa�C��R�V�-�1����b6��3L���/L |$�E	6�?Q�P��'W*2K�3-�u�@F�Čʉ��P;� 4dמb
2끃�Z�I� BFL�h�25l$���jyr����	6,�%{����+�z��W
+�Nם�{�ܤEx�m�4��bi^�>��s�韭]��A;���
#�����23����E-�6��r���`w,${�bY����Q5�ɮв��.�g���	��ڥP��1m��p<�f�'���� 	�}[�q���2�)Wi�
�:D����&^n���u�������zW�a��eƱ�91�M�3�Xk��I���ASRN�:X��[���Ӧ�ďړq��R�L�F����+���!���D�k���� !GH��#0ϝ�jNB̨v�)|��'���V��o������J��5�4�7F�	��속~���Zsm�P}2�զ���+Ϩ1߆,�D�G5C���Lƌ}���H�O+�ք/_�p1�$R�I�����;Fd��"%
�EG0�a �L,>����ᤖ�.Z�Pa���',��ɷ���-ly`�+[�,�B��VBJ�y�ಆQ�u����҉�h!����i^�$�Ў�7^Q,�JqD2�����Pp����f�}
��.
g�IWA����A?����@���6��л�)\�c��e`$K��R,�{#�<{�C���C�tseAS=4��ȳ�	ܹa��ap�A4V2�Ӌ�7lɈ|�ъ;?���D�5�
�>Ѧ��⬳SJ\M��@���h�v���
ü\_;p�V�[�)]`"r��@��__NL	gO���%Q�"+�.�u��v�B�c�Iݐ`!x���*�n�hPq2�R4|L�x�Jٷf��	0��a�3J�!SƤ	[T�5l8�Q���=�J2l�1F�h���MR�88�),�R�Y��;7��ȐeH�"~��Bl��0���ٳ�
V�$xbG�+)��'�6	��,�%O�:��� zu$�J��҃�Fp��
R;+ 0���C)4��ֱ�@�D�9/( �ߴSk�MR�AN/l�Xy5��Gby"��Y������ RRdR�$W�pآ>���,j���jtdC�@0۴b]P�Hy'd��GB8@84�3H#>�e�qM����A�@4���^Q�La$�,@M��s�A��R�"ԡee��38�V,�a���)"T)2�F�4>��]Wf2�zF�I�tYP0�&��{�T̨��.c����EAskH���nD?g4�"�(�rT|`��.z��N�	��T,��}���s� ��,���qT��C$�\zD�ņY%P>!ZV�=C[�@冔_k��hR��b�L���L��R$���Ve@$��oD�((ڼ�0��#z@�p9�fŀl�H䭻2'6�S��>�I�,�^�����|�=�e�.9�~١rH�q�a1vWj����ם)�Lݙ�!}�-�%/;�dՙH)KU��k�`�'���W�ĲF�(��䅞8u	� H-Q�}J"?�dIզ/���տ|&Z\3�&F-/$����H��pST��W�5sbx����ߏ���{�E��| PL�F�/+,��`�Y�uYR]�d�D���EA�]�o�e����ȃ�H�:d��'
$�� f�J#)�Q��-.��M��
8(J����!��\Di@ŧW����BdN�(Fa󰥄�+Txr�K�,D⠲b!մ	VP09�柠�"N�Lvj=:4�Σ~�29;�d\���Q��M���2pA�Q���GH~j��O!{�$	c7D��Y�b ���ȉ/w:��t��;�����K��yB�S(Jf�́�K�<����ȉ,s0��D�<�2 "�t@,�S�u�E�ε>ܤ�#�6�,�hQ�_�Z<�t�3A��=K`XK��ÏX�U���ި�[w�4� �ʭ���7�S>*4��yB���|��oz�0�r�[?A��W�~̓N|§�'
�(��J���Xbh���(�bG��1=����Ģ����Q�ép��
�1�@<r���DH�;ޘM@Q�nm�!g���[�V$n�\����v^
|�e�Eps��z���r��j.��Cg[2/4�����:X'���B��s%��A�B;(�D����AY!P0R�BK�~$批^*Рu�ţt(��9P9,�
\S̓.�p����*d��+R�4��'
��;r%�4�:�ه�I�_��"�Y�'^`��*W�"��׫�+�
�ѣoؠ6H�R�b��2Ȁ�?�� �)P�6��Wk�*��Ϙ!2N�Z�+�
U�m�G�ƊavL(qΑ"��I�)��	!HE;Bl�,���×jQ�1�����ug��#º�� e�2���ig@�1R�R��,�� ہɊq
�@�����r�H3���yw`�B�9O"�{��!���f���8=:� ��"�.8��J٬o^��hQJ� ��K�O`��&E���߇rt��-HDB��Fh�".������n܌�!��E�i����_~R"�����5O�ਃ�qs�u ���6x�s��3� �1�� �0�iA�B<4��	�,ҟsu�i3@��2|���
4�2�i��ĻNy4�J�# Qp!ȃ�Ɣg-D��L<I�'�(�^�I�u;ʄ)@�W>�dXQ��D�M2�I�YAnD�#V�_���Uψ���%<�rE����\��\�ю�9ozt�kğ<��ɧ�АR@�e�<�G����`�4�G���l��O�('(A��|s��O�H��P��b����;��m�\��aE�*��ӱK��C��e�&i�!V��I<���{�*�n�V��Q"EX~�"N�h�x��Í�9�Q�B��.w(欛��W�?�`)�C�-0�R'�8m�n��3-���$�9렁�pM�/<����C��x�QR�|��������t�Ir�'�"���%P�2
	h�ˆ$`��($+SLV	��!�|x.O2m)��e�p�+�%f��@��ҏM�
L)6Gп*��$0QC��h �I*2�Tx�L2b)�f"���֑:}�c�%b� ��޴�~��;ȨiZf�(n>���,ג8M����d��.I���'��3��Q`v��Yz႒�l�'ʌ�d��1����R��q�~��g�-gj(Ț�ղR�BȎ�Vx�
f��-Dc���F��z�/bc<��� �W�&� sFܛ\T�p����L������>�*E�I��QRG�%<��i�n�,	�L��d�i�fI�CfƄt��%��1W��c������'AԒH"p��2rPd*�N,\O� �8��ֶh��&$P� ���;�n%m`Mö+�dK�̌�b��@"��j� �+f��� ���cn���@��*�H��CKg��pv؟��Vρ�=t��)���@(�%
��K�lu!'gߙAˤq!!N��_����ĎV�rw��Y4l��N�
��O�|]y��^G�p!#[�\��q2N��<�d=�����܌��w�tr���u+ٵA�����
g��m�S�\�B�^paqc՜6rĩx�^:|�5Tiŗ1F�9��]�b��]��=�	�&GT iK�$0D�Kq��*N���`��!�,ĳ�6��3/��M�:F�e�D0����<��I��
�@9Z��a�v� �G��*:D-��� 3�H(&WK��s&E�g��A�@��%��`#��eV�)hvk�4��A�1��0�@=3V�0X޴jX1��c��aZ����v�֕҃)W�.vlkqឋ%T�4��v�Ѕ�vC[L�n0�`�Z,͢�:��T�h:���LƒԬ��l�,T�\��������	ר�2�lZ�Q�F��&��0*`}�D��ќ�r�4��Ȇ�I@�4HkҫE9�I,.���#d�AXxT�Uh�{8N��&�I�M�L�%G�[�����#�n���p��B^t@�=!���9a`�I'��$��0�4& g���8�$��Ě�.�*K+��I��L�O��Y+w�9Y�������LGZ\�ʏ=� ���-�(_3�}�4�e�����S>p3D��𦍍w�b-r�!7��͍v�d=R��W�^�>�7��i��87+נtz��]w���5�Q�-^�QB�KP'`�x�',�q�B#����}����N��S��ߗ(7�a2��x���� I�W*�a�b>��<�y'���/�1ÇAF^	h���#�y	ݾq���&�K�f���K����;����\o��V]�-��8?
��r��k^�h��fo����Q��ߜ�y��".��Y���R�|-0H�.�"<ݜ)�2i^5|(M��qnh|8��[u�"��5�$݅��1~�P[^�8[��zi�#�"+8�͡� (D�d�FEČh ��fD�,r?�� )D� [fٱ0c��AD'W��l��� D�j���)*(:�)s�ˋ`Aly��;D���@�>x�CA��#j�X��E8D�T�%�Q�N|�i�ׯз^,���5D���S�<�Di�c�\*���E�1D��Q�L��FZfe;r��8s�|5�vK)D����Az��! �c��j���4�2D��a��0�q����7��ѱ�0D��GB.���K֪T�~����'f+D��`X�q���	�22�@�B�H$D�8x��(BZT����
N�-:�D%D���É �9�%[*���Ī#D�Ȃ���H����1�Z�x�F+D��ʐ��OL���'brd�an+D��.˚DLx[�"��_����6�$D�h��@-	762 ���Ih����%D�`b�T�!�&�H���R�r�C&D�� cV�GR~�c��.%sdc�&9D���%B� ��mh��Z�����2D��y�'4Z �AS�J�R8�k$D�0I�ۉ.;�9��Ɣ7�<� S!D���2��2F�� �rND0�<D���@:?[�u��eU�d� �Q�,D�DV�P�d��y_�5
�c9D�$�D��1�R�a�KümJ���9D�z�l
M� ���/A�o\��`�6D��6iC�.h(�-_�3�B��Df:D������F���4�ݝ09���3�%D�"3� �NI�]��e�;1$ԭHA�6D�8Iâ;H�t0[Ԉ"M(�	r�"(D��Pqcߢq!n��P�4
&�* -0D�hX� R�9����P�@�hr���:D��� �QF�~�i�ڙ;Z�x�E,D�8 !��+2ٞP*�Κ�%"ĭ�R�-D�$J2��Px�4�'�1h3�
��&D��qbF�b+�� \�L�4Ѣ�'%D�#0E�/oRaP�O�v�)��&D��V�܏;�HS/G�+�?!���d����W)(��) 1%˛#!�d�t`�C�Ѳ' ��C��ٸ7!�� $Ո���$�hl�碎�w02�3"O�j�GK�J�}���P �$i$�'z�L��+�g�S�O{��0g�
�����-ʃm&*�H�"O�t�A��-������}:v�O�e��G �]��ӓY�����_�~� r�&�*�^���	~�$z�F���T鲥�ϩ,�j�����K	@t0�'�&0��0�
�'���mM&(�PC@��Bnn4�I�<�����>���H��ÛZd���4e�C�'k���1��?>G`�S�	!I�<�ȓ �)ʠǓ���a -��O<!� Y�r,Y�!���0�d�Ŗ҉'VI��邟�����H<�V��	�
PY��Tnnhc5�H3O(
���:F�ن&@7R:���A��u��'��  ��2=�PJӂ��W�	K��D�?=��H�)L�I� ta�L.&���Xp�[��7\��0I�kK�2;T��`���*�u��ɑE������V�X�S.�~Q��n�p��EJ�w;��"���n�)��*w���ǜA����rE������<�{�B
����ӽ6.p�����sG��8&JC �"Ir��E	P�<�2�Of�"�i"��'bP��NB-���0Z>-x��Z��ب�Z0;���{)&��æ>r��T��{BC�9Fa����w�~�ki�74��ZR*��8TN�&Q��5捁;��)���ӢE��`�%_�Zn�,��\8�61b�#[�=���C�! 1�X����?{a�(
�f��6?�*BC+��w�̣ro��H[w�����a}���I#�q=�����
W���E�rf���hI������*KRHh'ƚZ؞X�={���P�G5E=`Ts��`l���L��H�i�(0��#��}���{�!C�|�^w�z�C#�O� ӥ|��pH�j�2�����~��Pj1���h��. V Kވ�;EU�kE*����ŗr��d��?'ZJA�v�B<Zti ���J���ȔW�1�P�U\�� ��-�z%A¡T$
��ƢJ�	�L.2S�����GE��"B,�J��B 6�X�Q�i��*��d^�]1��� ��#�@��H�JU�I��C�>
w��!�Ų�>���E_Z=�b��{�	��&�\�N��\��c�J>"��Qp���L��q%O;<�ȯ;u���B8Qn~D�N��+��DwL��,����x���
`�.Qc��E1*�h�`����'Ǯ��'�8�40��`_(v�FT���9�}�#�B�x�
�)�7"[�����=�:0�����u�JH#bE	�}�M	V��U��`�# 40�^`�#,O �{�j�nm���χ-˒a;5땨6E���p?�Q�g�|��Eꕘ	�(aI���:�6���@([�Z��0HR�?��B�Y���5
U=*���A�1�^H
c��n���'cJ��d$G�����U27�`K�U	MFh���OUD1�e��2�ZTӧ�܇?|��f�<P4�q��~��X{�YQ�ɿZ �1�	���O>�k�L T�����N�{�4��!mB>A��, ��g����
�<�{��p[w�fur�c��y��UpW@�BC2��u�	�2Lt���V�q
�Q{�$�:\��X�剭���L���dY��K�gJt�j�%�(N�ܩ
���&~��@&d��SP����ݪ�nE��됊aHv�Ee*M�ԡ�R�ȟS��W�5)!�v+�$�џ�!O�&avĀ,F�x���`�IO�H��
�"`�r1�D
� r|�H�ɑ6H��5"v
W2I�"$xgo�}�t�{�L�F�td��}� ��d���x3�����T%a]:UhgQ%Ǹ�q���?FA
��p? ��O$���fg��,�÷�ƀc*�\+��orbt�I?}�bx6�N���g�6���͘m��9Pҫ�)Ѽ19㏎�]՜A���%�@�z�m�Q⓾Ov�r�B��"n��q�d��!bm@�_�6�*\�w�!'G�X��P�W����P!d9�4m ���a�κ@`ݣ�f�w1F}�� �	���#�a�;i`u`7#�i����j�:Anݫ��O��2�W�<����pJ�q,�H�'!� �xa��^�
�npq7��:s��יPp�Qk�W7i��<���F#��%G�5W|}��i�2	�`Tr�Yy�ڧ/�.���~bMך}|p	Y�r*̡d����	��"���pwb]	E�j�;�M~xp��Yp/Ƶ $mG�g�r�IТ�z��:ө� ~j��%�]qܓ5c�
�Θ�7�#>�����nʤ Y�zl]I[ݓ�aS�lX��V-� u�Υ��P?$a�ƅ�o��J�LܛLW ��R� ˨Ā������]{v4�@�bH2+0����5qr>�x���3/PVe�WI�R����PC�T��%Ն�P�hŌ�Z�m9���-YBM���UT������B�\��(�4!� |)�q�a� I��Gy���8�88�!R!x!�Y���#O�����!{h�b>���2L��`沴k�'��%|$H���P�.���I�K:~f�R���Ҽ'tF��B��&S�bhb�R�%qH��⇚�$�V|r�M�5&�>�;2��/w��@��$U�vLK�S�"~�h!�T�dr>9�u�*U̚U��鏔�Bqbf��SX���0%Y�}}�	���\�@��å�:_����+�̵�mT:=Y"�۰��yt��JܫZ�^��S�s��� o�U4���A/+b*9"q�%�O|U9#ɐ> d@ȗ�N�4jȠ+�SR�r�)�˜�,
�<�&�cY4�pe����ڂ`�6bڈ{6%R�Q�z�9�k\�( �p#�A�S��!�!��'�ؐۓ/�I�Ks����5"��B�&I�a7'^�6�<�W�^�lK\Mv��:Q�U��^�m������'e�4�C��Q&=#�ŋ6<oCHaz��ɾA��9���P�`�$���	L���i��-a��M�	˖��d�A?C��1��h�� ���H��s$)��f���lZ�Y�R��󊃍_>��dǾ��j%�Ob��-JP�^��N/{.r	򄏆�3ݪ�1u�D�W������H�p�RMK�T�Z� ���.x-l��?�V����A>g�Xh#��#lX��'el	�`��!^�:j	�vF�qcvkїi��q��\24��p:�D�c�Y�v�yW�;J��wE�}{F�h��q��ܳ7��Pz��
�I6d-#vK��~j@ĸ�Â��(O(4[�C
�M>t�­|iHА��x�q%�d�? �X@ w��H�,�j���zW�4w�B/�̒��6��-tR�T+�ߡ�(O
5�	F
��qsd� ��e�3x�h��J4@��hQB�/YQ)�W��
��i3�X%���5e��z��Xf�Da?�9)�F�s�LaԄ
gCB@9���SX��9��Y>Hs���Aj�7�Й&� ���ägN/��XH���l��)�o�Jw���	�M�M��S`������"� |����bx��藄D��b�V	0d����{O(����d�f)s��@�IF|t��D�M���S,dϐX�H/�@P�O����ݤ���&d��Q/��͈O ���Ꜧz��<��dȥT$�Hs$)+M�4��v��V֨Ti���V-ƕ�0j#�d�^�#	��L���A�H�4��%B�[�D��]��$+ )T4<�E*��Z��Ů������-V�N��G�L�^���q��eق����oL���'PP�ySMW�`z
��� /�!y�E�1�n�Y'�N�!�¡��3SV�ac-�a{��D0O�)�w��43�N�f�8�,5��a�]�,rt�ؚ>�`�D���+L�Y�P��D�B�f�;�JֽAu���+؟�yh1!�n�3�Q+Z�V��'��= pb��6�qЂ��8C|����r����S`��&8f.��0��t��t��<>�J��1])�܁��ڼ~�Q"�S*B���
�]��c�'\$p�<��w�|�Dx��ɝB��:k@!7W8��"��s���1���/!�0"��B:5) T{'ψ�F��*���P�`��	 ���#�V����f�e���v���vk�0X��I+j��I@���=�_h0R�\�tTi��N�E�R��'�&�БZ�E�>�,9D�ę}�	c�J��r\q�cC�H��w!2-
!ᢄ�G6�ɘ0�U�H�	��I�F5�ݨ@H��M��`Гx%L��0�nY��m	�Ir.�&�#�J]�_sv���-��Nt��r>]��'ֈ	ք��ԠG�C� �j\>;�
�n�!�nI� ��
L���&�@�`EH������\��� M֥
Z
���K�,x~�6�M)LJ�Ȃ��G�| X��#j8Լ��@�*U~�	mF:���6�6�cʔvc�`�C�C�>)�eBh�!& �]K�X�;�,���B��#��<�Q#&dX%8�.�l:-B��$�o���gUoi�l+�+�f�bh��<
���6�M4v���9�
eK����6�f��&��S�P�1@��8�q��'�j��10��I�T��`�*pz��f��S�X� ��9�M�2Ǘ*m��}8�c�);�Lس���v��5y@�>O�`�CaN *���;vĀ~ɸD�Z�f�@9 t�X�X�� L��JG�u͔�C�ՃE�	�pa��$�'a�^x�o��]���� lVHA�Q*�NbD9�#C�M�������L�	�D��F�H豁 �Czj��N����@�HF&��xG�� X�+���
��E�5I�%p�5ڥ1BG^�� ��&]��hbW� Z�9cD?��Y]�q���Z���m"#J�q�e_�\ �!#m^4%:�����]'�M��K�4`
����F��Mk�iW��(�
�_�"i1u�DUO��Ô��d�&(�ŌӕV�^�yń;O���4萰w��Q�h4�-�&�P:J�
C�ˎ%��`ӱ@0h;��$�q��Q�h�� �)�6�:K�!���F�7W8T���G]6^�Bل�	�R^Qx��Y�s�lAc�#�M����1�գ\Uԑ*��	a�@ �Ĉ*D���(2a(�h�LE�K���сBT XYΥr������Y;#c\�KA�)�GPV�JU��)M=�'�����[�U�`���I�'�U�B��)]���P醺h���Cʊ�/�F��!�̂-(�ă;����B��lJ�yaL�g�Z�S��p
��ۇӘ'q"@P���Q���aҭ&d#"T���C�c���I��]� �0Y2�bC<{6h�KS���iZw������N�����ҺI����  y�W��<����+ꆱq "2,O,tB�AJ�z�BgG[:N�`�B�E@��Ȑ� )uw���$ɗ')H`y��ˈ{�j'�[�O�p�Y�"G��h�T�z��p(޴On��a3/�V~*p3:�qN>i�!z�(�!�̾lRN�`�k}���0�	>nb��𠎺+Q��3C�'D��S��V�	��2W��`DH< gv��p�ϻ(Vb��7>�@q�u�߃M�`��<:o2x'�����/||�D����j���+� j�,��ק�iwҥ���Χ2f��c�*R.z��6L��<1CY�&�(��2'��n�5���N�0c��{�Z� C䀗*9�"i��X�&L�B���<�R(S��R'<���.0������1�4A��,\�j�o�S���,I�s.8T��R�NG3BO�����)���@��x,��_,�~�H](}N�`����'���y'mJ��L�r��9j�h!�qos��E�D�ͦ/Yj��6�!��-_�L��|�rŖ�h���ߜu�\a���=A��h�NDidjx��'2��#T��4.�Tȡ�W�Ih^ԥ�sm�/ܭ�v���&�h�����	H8)f�ť~��2r,9���8 ��d�@L��n���`�I� D&1Y��E&y��rl���H��g-�D7��w��a|Ș�|b�Bc~̈1�z�b$��	�{�<���FF��
b �݋����Õ4X���s�Ñ !��I[9ZY�e�ȼF7)Ђ\	�����'���[���!������Z����56h�Syr���(~���P�\D���u���T���"g��`V�:;n� �%/�tqd��q2�0vhp��e�2 L�A�|l(w�ßX��_$-�p%?�I�iŦ���
�H��4n� �
���l��od���A`T�N�
8�끘k���&�0��aީ�D�!� d�?8r��P��O]8�"G+���gN����>�d�P�k)�3)�/HX� ��C� $�J�GR�]����TeL�-=�	�`��F}(��iJ.JZ�4�2�_
-� :F Ƌ 9��AQ��q宬�"E?`d�D~��Ίx��'�U+��#p#*�F���(�e7p�*��X�<F��R��*�:�h�F-vD�)����-�T��a��d<b��Y9L�5��-z���g��?�I�s��([N��O�A�C��ZM�ݲ�'ˮy� T���;�D��uĘ/q�l�0�1��y��<R�4}k�-	=
�jC`c���Un�OPY��C /2��%>�ɀK��Y=>�2IK�c�<x]��R!^F���5g3��G4^<5��dX�8�(y6�͂=zYӝwt������
��߳���'���� �+[i�!����o8�4�3A�44<��8#F��]ƴh#�O�8zhs#N5n
���˶$�V<���$x�K�kH�P�ǂ"ƙ#e�
'x9�Ԭίb�xu8@<�Ozyr@ݻi�ZP�H��Ċ]P�K�������0��EY�,��b��(0�٪n�H((cȚ��� 
���-�C�? �Uwk��"I��� 9l�	��I8Z�j5�.��%��ˌ�S簸ӵ�35&��LN�.6,�q!�[6G�^�YsC��A���r�'C�iSM�72,��\>�le��
&��U��=)g��x����'�r�r�H�]�4�c��O46�p5K�+(PА��U��|���K<n�m!rB�1G�N�XWCC�J�D���!!�k�I��8�N��,7�ੱ��j�l��3�^!T�+Lm��������b���̞��F��;��5ݴ:���Ο�
��ɷ,D/Ox�����6upS@i�8W���Ӗ9:Zx%̈́!k���+5K�)#'>I�cĂW�V(�v	
:P����ɔ=2J08�- i���+� Rp���!�4?�.�b�
���O``�S���u���I��U*V���A`�F�p�X� ��-OQ���lU#!��ti��\��$��OT9:���s�P� 0�?OP�J2ۤr��2�F��VT��0V�< b
\�Jq�#LU����f	#�ʱYH?-�WJƎ2�l=
����"0j��c���j�xSm� Fa~HR�K��<�'A��z̈@#2HC�H��`*7�SyRA���ȴ#�0 �4	�'q�4�'gG�Y��'OT$���I	=��8႒�܈�c���1(I��O� ���^�����H�;�xl��I�t�d4���?<�ƽ�n��8��!W(�1X�������|d�!�	X�ԧ�	$�Jp����<r2r}+qAϬ�p<!�E��O����Ս$?�� B�zA�D	5u���[�\8��񡖵N�����>���~&���C"TG*�[f)�N�|�p�8�]�O�x��{J~*1���V��Re��x-��#��f�b=P����/_DM��W�p=Y�
Rl|���T�D����e�@x���$��@����s��$���`�p5"T(�����S�"l
B�	�|� )3L@�I4) �0�O6	1`G��	��h��H�F�{ �U8V�Q��)Q����"O���GO=/�X�Q��|tԩ���ͱx���2Ƞ<Y�F�b���DX*	~8SVf�uJP�fԀ/t!�d�G��<�F+8,4��:%��+J��ht��j�d��R�'�(��4�
Qj��I�˒�<]�%�
�D�(a�Å�>91F�6��0�X>���,�[�<q�d�X����׋I ��uw$�T�<!���zG�l�`C�$y^���Lk�<cH�-X�T:4����f�<���(@�Xm�e�=@:�HV��[�<�Ӥ':�a���5&�6И�ZM�<�`�O�J�֑Pu�ֳq ܄�%�f�<��)�1V����m� �*��+�n�<�����3�B�	W��e�t��unZi�<�A�O�\��bJ���1PgAy�<��,�I��U�(���/�w�<��*��p
$��������c��z�<Q��Ԓ1}4Ȕ�^G�St �~�<	���9
RLƎ G@�
�M\y�<BE�*��1����z�B�
�p�<�ЅAI�&�c�J�|Uzf�Pl�<�a�"O�ei�*v�n8´� F�<�!Ɛ�Hl*pfJ�T�LP:W�@�<I� �G�)*�IP�o֮��Gd�j�<�2�Ï?˘��G�* 24��7�Z`�<�v�T�[���y�N!]���&G^�<At	V D�`$�3�R�L����CȎC�~98T釁=�6�.Pj��4r��>&8��w̏
9�.9jBe���d?cV�m�#&U���
q'��GkM�jz8���j:�� .�� oZ�3XZ�I�O?� c���E�8q0��B��2�
�Pܴ.�٩3P���i��N	��㳤�^�q g �Ml�V�>N��	�R������-[�Ha�`	�@��O�Li�@I٦��D� JA�!�V�AL����OJ��	-B����I^�?���?B'e�-=�P����{8t�cry�l��cH5z\\�&�"~rV�F�s
"h����1~�Ȥ�%�D�g4l�0� ��S�O���@�O2nqsFL�7��� D�A��$�0�V�Wa�I�E�z��#�'��dm�:Lv�`R: ��KӍ��$��t�~�HB`Ѓti�5sr�O0��2b\,p(P�y�#Y�+V8ip s�D��.E�:�| '���O1���ċ�j����O�s#���T�ZA���FJ�@�)�\��� $yJZ��%T����E(0
D&�06�=�`��N�h}^��D+�7�<T Sa�;t���'=2}����w�a�4F�93�B��L�>��RG>�ē" ~ 1����S�S�.%r�N�0�D�SЫ;�ʓ:4�d���S�π |Q���N5c',��6��$c��5�i׺ءv�'�ɧ�)�8
��	�'���	a�Y6�
��8[3P5�ڴ�y2�&_��' YG�t�B0k�f��I;a�� rhH:6�(��J� �䓶0|"��9n����MJ0+�~�W�M�2-��'��G�W>�+&g�06Y�ir���^�'+�$U�\�7/+�Z��L	�V蜳B��#A� b��� �r���+��D3�J�!Ga���`�@WbľAH,�f_��?	V��t$D��� lG�q
�'XӶ({��K#��RJ]�i�4���2i8��$B��.����k�I�O��ErÑ$W�"��3gU%��y�"O5c��\�D+�1x��z����A"O^� �
�^:X�у���4؍�"O�Q cDچ{����'�=`8��"O���슺!�JH�փT
l��B�"OZ��$��>(2�@�b�)F��"O$H��#AP51wo[�O$4�"O�����_-��Zd�Ʉ�qC�"O8p�'��,�|!��L����G"O2}�c��5K6�ŨA�l�{�"O���v�	6h�6�i�!	D>�!�D"O�\�'.A���ap�T,���"O&5�0@�(S�X�����<G+0A�W"OdI�Qg�'/��a%$Z&0ɾ�"�"O ��̒
�b���7N􉱒"OM"��5��ePҪ�/]XI8�"Ob���P�xa5�Ѫ)]���@"O~��"H9�&0�@
 ,S]�	+"O �:U��΂�`Q��X[��	�"O7#
~�j�a�L��2E@��A"On�a��2�F����K
<<���G"OZ�Ä�iE��k���	LŢ�"O踁ğ2_ �8� Оe���r�"O�e�RL�|�Q�P�,#�R�Zf"O�9q񬐙{ϼ�s`��#�¤��"O�qB$�J�B�M;�C׮lx:�"O�|��jR#'D���·[>,��"O���S"ɇ|`����"M��:�"O:$�%́�"�����6z0V�K�"O�Y�qNn�fd���ȷb����"Oh�J�#/l����\�i̜ERT"O�E�wEE�;�T|pCLR�'��F"O<�p�	���*���[�7�"���"Oi�a#�����0�F�*�A!"OEQ�KG�9�^�k��+ؐ%9q"O(ܹv$Ԓ|�~51��O5{��A�3"O��@��&�R1����)3�~�X6"O����nѴY%&��/�G�.a;�"O�����[�<��Rm+x��]�"O�!dB�=>�5�D��6!"�PR&"Oby�������9j�h�&E8�j�"O��T� �.!`��e�ܡT�&���"Ob}A���9���ڔ��K���RW"Ot��J�����(��Aת}sc"O0[�F�0:*�t�	�~��` �"OܸBÔ/z�޽)�++�<�3�"O������(&&���Ɯ�[z�|�p"O(���E��[J�h�tFV�g����"O�urv��'6j9�D�-KB��W"Ox�Ҧe�?[B�ͳ`�;�n�d"O�hȴH�,-�	Q���z�1�"Ovu �Ý4P��L��υ�Gef@a�"OH��g%Bb;v�m�+9WJ%��"O�B�c���H�W,��x@
"O�|*gJ��D��dcS��2X���	�"O�
T�Wpҁ�#L��hG"O� T��C 8*��!��Mf"OFl`�@?��,Z�n�|�Q�v"O��Y%�� b��AA��2H�^�W"On9�G��d���Vk^�v��P �"O��ڌ
��ph@�/T,�Bd"O�ɔ��5iLຆǫAG�!�"O����fòAO!��fPϲ���"O�Y�!�1�R%i��/I�h��"O���s�����R�H��@�!"O��	��JOgꕨ'⊻e5�T1�"O|�3�b�!�@iA �'>)'"O��J���$/�N�	׮r�� �G"O��ԇ	)\�:��JT3#��(`T"O������/<V8i��$o����'"OPm���9:K�Up4��;P�!�P�\��eq�"��N��	��S\n!�ʤ[�V�
EO��>�:ҍWZ!�+Dh5Y ��<q��u�$�Æu;!��n�T�	�;Y�>Y�"�!���?�Ȕ�%M�"l�
���;c�!�Ź=`R�2�#@6��L�")�*7�!�d�'�$�������;Q*ĆL�!�D�u����a͝a4C��T�F�!��԰'9L9k�,i� ���&y!�Xr�3MM�(�v S�k0?:!��I��u�'J�Dm<�QSk�}�!���'G �����0`�;D�мD�!���Y�`1���$L4@�Rğ�-�!��U%-BR�̜o��rDC٪�!� %�p�3�UjԅbF�ǆ�!�P(b����T
yW����b!�d�,E���0k��K%H�8Ō��w_!��ͦӆ����1�PA�]�T'!�~� P�^�4��P���C�!�d �Jlԑ��&�/8X�]���?�!����\H����A�^11q�ݕ^!��^�݂C�G���0 'BLI!�>��E�aL�����Ѱa/!��DnqJ���A�7f����&�G!�H�w��!`箌�;τ�"�_=3!�^+ZZxlC���AȎ46kJ�S&!�D�<g"QK�I�
�`�����uo��U�>�X�!hC�P�^,�m�yBJ� ?n���qc�#:�2�YD�S��yr��,NX���jX-=C|���H��y"��k��a!ǁ� D|2����'�yeV�|�@�8t���0K.�:%#�+�y�B9N�81+I�"3L0��� �y�@��"��]�M�P�ZF �1�y���,t�Xxq�"�}��ҵ�Ϣ�yB�L�.��$a�������y2[-�����K�%*Ա�dW��y2+SihB�K ������cg�"�y�k��g!��q���9aY$=�֣��yrf��Y��YPR�a�U�r ��y�jך`2fls�b��g.�E����y�D�`詒e�`Q 9)�J��yr%�?�"�8�V{x��QO�y�@���X����5w��a���ش�y�剖?���R$�8��j����y���`��9����z���͌?�y��Ǎk{z��aǏ�t�*P��N���y�Y	�n���T�hI���p���yRʑ�[���Y��L\�RQpeB��y
� �=&D�JP�+��Š<� ��$"Ol��Ee[�P��DP�Xx��%C"O&��� HF~Lx����A�S"O�A�E�@�6���Y����Y��"O�m�u-Z�E��NC-L��H0 "O>�ڄeP�#~��{-��$u�P �"O�݃#�����q���yt�$"O0X���ս7|Baе�D1iF�
"O0t�S)[�I=+p@�+Nk�48"O`���R�|�fՂC���&Ĩh&"O�I1&�I�Fl�2��V�L��]J�"O��,�� �p#�E�.\0F"O>���RM�z�Q@kL�p�r"ODjc���GV�m;��8��"O�	�Al�6N��Aq�� P�"O�5	3��>Lj�i��Ewh�"O.Ds�,ل$Z� �s��:fְИ�"O���sl����0&R'U���G"O���
�Y����å@0uN�<ۦ"O&U	E+S:L�L�s%� )H�\�1"Or�����]��UK�LޏnS�|��"O8-Uޒ%�,L����N�L��c"O��h�Z�>$�1"^-^}� �"Od\��M�O���ǈ�D�!�"O<X
F����u8��ӕH0�h�"ObJ�I)y0Ej��ڧ9(v	�"O���f�<X�pw'ݨ'  ��"O6��g�K0C�z�! �e�Xb"O����àHj�p��W3�츨�"O�Z�E�� �
�����@��"OZA���)�UC����F�����"O�P��b��bJhE�CG	�b>�!"OМ�be�0e��6iP�1��L�"O����fQ�4�`��@g� 7��m9�"O>-i�$P�p���ƆI�M����"O�0
��	b�����7+J��"O�Apq�k������JH$ŀ�"O ��a�J�A���h�n��D=�(ؗ"O.@�R�J��Q���$\Պ�K�"O�Ax4/�0@ψ������p��'"O>QwՔ#��%�s�O��X%�U"O����މ,}����d�&��4��"Oz���IL�1�����4/��u��"Ox��ЉH,Iò��S"Ǹ
V�$C�"OP+d䌲#��Tc� �6����"O����X2{�Xlg�܆�d��A"O�$p�iX;8H�9�ߴD�H%�"O��2�`�_�0�2*�r�z�r"Ob4�C
 y*��cgJ	X�^�k""O�D8ej(t9�a˚V��%�"O>	�H�#J�<�`�9�45"O��D�җO�^<AB��+T�y��"O�%B��ބ1s���� �"O�)!𧟰 -p���ִ�b�aD"O�U�ąՠf8j%��ـ ٶQ��"O�Y�D隰{B,���^�'���v"O�#�9yߚ�!�N֥s�B�k3"OB�Z@� �Pyӧ��i�РyC"Ol��$,#$�
T��-WP/��P"O�0���b�x�B�5t>�PF"O��q�š%��M���>HȚ�J�"Oy@$�B�"��#�q�7"O`а�	�<��5CdsZ��$"O"�� ����9�1o�8?�Z���"O� �la�%԰k�0u�!
�l钐�"O�Rq/Z���@S/Y�#�!a�"O
ɺ��-E����O�#j��E
�"Ol���˞/�� hf(G���T"OL��daM�W�@����|��a"O �ȑ.20p�<8�m!(
 ��"Ov�+�D�!դx�Q�G�$%��{�"O��٥E�Um�#i�;@
��"O�@�1E_>cD��iȭVt 0"OQ��W�#Z�q��P�j"O�Q��5q��X����M:��"O��h&��h�
�ط JI�<	k@"O�}	�CM��NT�@�6�N��S"Oz {�
   ��     �  ="  �,  �6  �A  �M  �Y  f  6q  �|  ҇  �  ��  �  8�  ��  ��  z�  ��   �  f�  ��  �  d�  � � 7 { � �! i( �. 5 c; �A H WN �T  [ �a �g �n �u g| ,� 3� A� b� �� E� �� �� � =�  `� u�	����Zv)B�'lh\�0�Iz+��D��}�2T����OĴ����?YV̒'�?��]O+�a�ڦj�ำ5Iݞuv����bMs���&+W��Q��D�l��A"����ֶf�����/��Q��`K�p���J�E��PI��
��H5 ����pp�#����M�����lZ9�$٢W+�||!�7B5a� ��ƢX�j+�{�#�ʬ�c�M�t�Z��i�����'��'��'%
�"��D#���!$�0U��
�GO�mò�I'�V�no�"�'����O:� y��O���'?�i�c.�7U�X��֭bw(<�2�'���'f2�'$r�'P�HYw��ɹ�$��b���W�A�y��Xu�K()�1�I~2�Ij�DG~7Q�H2�����!�o��z�acˀ��n8�'��'�$����f�17;�h��6�b\[&��P�IԴE#@IkA�'�r�'�b�'��'2Z>��;%�6���� :��Y�H���¹�I��Mŷi�6��¦M���M��n�8��b���5�(�9 ��#ݠc>�q�Z+@��L�O� �	�_+^�D�������=N`�� GA�	T�^qsRD��R�|֏�|�p<�ŌW8���d���ɭ�M��iM�ݟL��n�=�"�ǜZ��-˵E��&����@�Ӧ}�s���eˬ��rm!u�H�x�Lȓ9/p9P6b���Mc��i/�6m�aO��(�
��{�4t���g���
x����OǦ!8�4G�����?S���=��g/_� ��|!��I0 �~|�e猰X���ҷ"ȳb�K_ G<��f�i2�6m�Ц-{�́��p)9�ė�-�����c�0��$oF&��`�$�_l���P,c����Ѓ	�N�L�cw�L�R�a���OX��锤�2vdZPc%�ڜH�P
w�]��,�?)���?�C��,0��f�?Mw�<r�\�T<_'* �B�O,��?��������|h�v�ӛ8a�aD�i�vHJ䄃�q(0�ǋ�\\6Q��'_�0�b'�$m4�D˱+�%oU�ʖ�1��t�M�. o��F��3�0<����� ������,��i����˦�iGg�#�r�'$2���O���O�牟�H�ˇ�U�?�F@k�nP����G٦�1�%�85B�bh�m�����P!�Ms,Op�bsަ!��ny�R>%�ɮ������Y����h�?��8��ן��CDæm��'ڋud�q���if�0��Zh�R�a��� ���8#�+?�QBJ�����J�?%<���I_�|�E��k	,�2I�sj�2.2���X���	�)���ie>�F�:���� M�88:"���1�$�O4�d�O�"~�0ٛUM��CcG�/C��ѱ��W�'�`7m�Ѧ��|B�휟Q�L���Ǫ#��b� ��M�����	Sh�I�Ok�i��W����� 50��t��-(;;��e���H���
����MEB
��M;�Y>q��n%?5BmrgNPw�h��h�:������.M�Иd�"C�-��DC���Z �D�Ơ�/B����lţX��7MBMy��W��?9�����|"ȑ4��,B�h�g��1i6
Z�qK��'��I��Z�O�eP�G˕GbTSW�V	Z����gS���شz��&�'V�7�|��'��	�#`4����ï]��}�%�!/�,8R��M}��'rP�@�Of��ٱ/�Rq�� �(0I���qK��m�<E1���=cB���)�
��Q�th�
CG����R06�H�(�@C�F��d��M��5���Jp��{z�pP�]� �� P�+� �:E�wBXd��$��m��$(��9*+z h√�
�0�I���6g�0���ß��	\�he�-;���O%`������3����	#ٴ���֬e�8n�$�a�lp���H#�DQ��+U���Icy��'�8��Ȫ0��(D�lMt�F���!Lz-���F rn�Hg��(Aax�\wY��@�ΣIv������A���CP����I�%fozu`�ԬV��YFy�(�%�?ǹiL�6��OV�B�V�W��%+�m80a�Ad�<������0?ᅀH7-�m�C�^.6��L´ǐP���Zݴ$=~�I���:;[�9S�퀝N7����in�I>�h���@�r@6��'��D�f�f�IܜS/����D)��×*�r�x���Oh葊�&l��4˜e�f�ˎ��O4&]8b4D��]QP`��������9�����o��=#,����&9$�+ajR�X�l��7
������)�]1�c��K]B�QQt�I��M!����|��1�`ɫe�r�8��' ��'�"�|��'�r\��7N*A9̱1G���u�{C����OFu�Iئm����M;�J�6����,��}B�KQk��@�&�ip��'��$��D��1A�'��'X"<������
�W8�1AM�U�* ��L�6(�lD�'m�$��p�Z,�^�'?�OaQ��,�,��	�,a���0�^��X��m u���K>1��土l�e��7&�P\)4@O:~�
1���%�(O��c��'31�"�'b�Óf=�93R���\�� �$��'�ў�>!��
S�BUR�!�n�5!\X��A.�<	��iZ 7-5�d����I�<�q�����@�@�ccH���MH�bڦɹ�ib�'�B]�d�O��	�.PR,�2Ϛ?:�jlP"��	RGt$��*Ŗ�Dm����R�����(�����7W��a4BQ�X�d���@W��r���xB�Q���}>���h��*#��ͅ�>:t��"��G���𦕻��?�*J0I7��10~k��RG"���W�ßT�	R�'LحR��D+GT�����%V\�Ӣ�'cD6��Of�nڶ�M�*�LXXg'�Y�I�<IScLl�^50�mZ3��4���
� �'���'��I�`j�1��="�6����a� � �a��ώ3Vy�*bkůk�
9*��'$N	���KI����H�z��t�_�\{�["��U��1���Z't0uP��ď�pG2$|�ҝ�'����t�N	>Q��dJ� [�<�O>Ɍ��2扌D��ؒ$�H1k���WE�N���d�ɦɻ�AF��:��8|	8mPE(��M/O4�{U+��	�I^y^>=�	y�>�U�OKH�)��9���	��)�Ǌ�dA�a�K�օ*ƺ���aꆭ����jK�r�0T���L����"�H�����'{�bmx�`�(imfc>Y�6Ɛ6"j����]�=�`H#?1���<��_�O2�9�%�� ����i�Pǝ�h!��O�d�����7�űǥȧ>�џ@�����S&���nL�~��SBU�p:6��O����O���aE��7�T��O<���O�杗+�Nu�bf�D��� �.M�ba��Sid	�ߴ5g4��*H@�g̓T9cUm�+x`��W$܂'�P�xB��d��̀�i�LL"3���Ϙ'�w �6i��h���
�!�xd �����>BB�'�r�d�-��Xāj:��Öu�dB�	$~���+f@�#w��0��{�6ʓ>쑞����'J:�;�ϒ\���͜�Q��Va�'I�i���'��'R�r�I�I����'nFD��*��`���ʤ�ބ}cܘ�+�J<�g���&����%�ݳh�$��(*P5~І�%����eH�1��2���:c��0���`[���ħ��M���+���Q���ԡ-V��(!�>$4<L&���޴��'� ���]?	�	�B�ĭ�"Ή�Ks��;F�#�p@��������K���	�|�G�q�l
�U��0�Rʒ�A��9 �̮:Bx5X���=,���{7 7�<��'�.8�i�c�����[�zZ�$���G�0^���[<q�d�<)'IV䟬��B~g�J٬��B�o�)�UL����?�ӓ_�����L�yp��!!�p2(%���=�?�Q=�腺�A���naj�N����'z~��$�u���$�O�'�<J��r�fy d��Gw�XI�$CY�ٱ��?�t�P'������I猡)��{��M��m��Ur���լE���хͱ���űc�� �d�J�jy�F �~"*��v��}P���e�LtP3�z~��ǭ�?)��h���I&g��C��N�f>Ȼ0����C�	ab��-��)
S@@�C0d)%��!�h��8HE��i�@�h��
0C'Zc��k�*���O��D��~n��C
�O���O$�${ޅ���ɩZ�t�&ʙ.X�2cՁH�VK���S�^�fX*�c>��<Q��&c(8�'X5�5P��X0Uu��C��|@�{gW#KPc>&��*W��[�����IKm�nŁ�g�O�%��������	]��v\�챃E�r��(��]�Y&@1#�'�T�gʓ_Hi�u���i=�	�HO��O�˓F�n��!��I|��	{[�3���Zݩ��?Y��?q1��2���O��f2�8��)&0Ӣ����̅*���q�:
��Ba�$;6�/��Ov���fy��$�a�,��3���B�Y`��n,
�k��i�dE2�Κ6�hm�B��P�<\��ŷ"!��j��1��v�'���'��'�B�'I�����
�e��T���ȁCD93$>��D8�ɷ�Hb�G�<�vN���Ƭ �̦5�	dy���b�����Ǖ�-$Z7��-u��䑂�'a������	������E�r�1Rp	פHtz]Mʡ{q��P1d�:�ىy���7D���qq���]X�(;KՁPp5[d�ܹ-ztHٰ���KLr��,��yb�Ku�
�Ϩȏ�d��|i��'f�	"z}�LY"��,!�M���օ.�D�O����4b;[�L�}���v�Ơ6��b�O�!Ô�GV0��td̲������'��I�*��<��4�?������p����$Z��Xr�"�:8�!LLG�����On�Y�K�;8�.4w�Z�m��Y2�S�4�?5Qϯ/	T<*�)Õ��l�S >?��ߚ-��`���,�JP��gI�u�Ƈ����q0� r�O̔�ޡ��N�S>��(a��'�Må�ie��ӣ	�^��R�K)V��a���O��D*����H�(	\�)UbB�<�&�!���=Yџ��4Y�V�|rA�_��<���	S�-��ɗAfI��'�r�'��uS��D�Y���'3��'_d��>m��d�]#v8D��iM�@�e��+?<�����4ᄁ�O�'"���wG��,�v����(э��AY��F�V��l`����%�����P�v��(�|rr�PB�,�	���i�Мc�x"�(��k�H�0?�t@�p��z��5F��{�����J�{���j�eUl�<!dBC�o�ĩ��⋹.�j-0)�dyRE-��|:���dV�&�X�)�`�ht`��B����8u./E��D�O����OZ�I�O��Dp>yr6��Jzpip�ㄧ
c��J�����ا�q���3��c��H����
%�� �
T U�6����Þ~��PY��Ё7�8׮ސN �Tब��E]ء	��dݚ ��Q)'�Υ}>lXa&���@�R��' ��	C�'�F��I�>7��"+\,��1:�'�6��jӓK@������)@�e�K>Y2�iRV�<"�ɓ��I�O�X�d�E"|�l[���+h��(�Oz�D�R����O�)�%1�(�v�(|hDit#��#-��D�p+�-g:�u�Q�186����d	���*��Ao��#];8^��. p̈���d��T́�cX+)��s���;G���'f�I�G�*���9U�(+�
ݥ䀒O���$�%��)�0J=YCL���J��CM�"��O���W*�R|`� �X�l����F�'���ݶi"޴�?!������J���7��(���Qe>1�A�֨�.���O�(b�ި+��[�MN�6�֐�U+B���t�?��Ԥg�Ȱ���?�t|  � ?�q�Q�Hd�U�M�2��J_�����=�6O�oʠ�Yc%M6�\ŃB��\1�f�O���3�'�yb��EJ]��(ʔ0<Z��FT��y��"R���&C(@d-��Ā ��Ov�F�돳Q�$\QG�V�0*���O�C����'���'YBƒ��yb�'w��' ���N�z�x��Hn��F$� K�����FBt��RT-4������?�$�9@x��ǎW7W�P��'��(*��N��u���_I��q��5�d�� ���R�E��\�3��3CJ�7͐Jy�����?�����|�Ú|����ă�9�>e�I��m��O��7�ə�H��I�ȹs0�U��))1�O7����I���p�O����i�O�˓+אI���:�qF|`���T�Vc-�����?Q���?ѓ��(���OT�l}<D���3`�Z������찅BU� ��g�l�|��'lz�q����ؤgڔs�S��H�$�&� �m��]lɈ�+L-e~h">��\���IB6-��]��<�b�W'�5�I���?�b�D�W��,ٖ����ԑ�*�k�<�f�I�2o У�B�1a�>$���{�	��MCJ>Q�[X<����C��P�XK��Is�"U$�p �������Iϟx�'q(Z٣F�:f/�I�㩈���q�F���M4:��S��>A*0�����O�Ɂ#n��^6��Z�ON'��وs�Z�8�����I��iU.,q�Z�?�ve��ɓT�<���On�.�r-�PD��|Dɦ%�J:�q'���Y������02����DǃY���S:�O^X�I:-.�1hׂ��Q>�=[U��S�����<�r�_1R!�6�'�RQ>{s�П�+��^��` !&��7lv� B͌ӟD�	:Z�  `�\� c���?�O7��b�։hW� q��R�a�% �\�hG
(�F"�x`�-ɔ�S��h����\X��`��1���������O�d%�'�y�����1F^<+��8xb
�
�y�O�	�s�BO�y�·���O��E��J+u	�&4Z5�u8��G�.!���'���'Ò�Y��-P��'�2�'����^P�C��pQ|����L5	�<9b��X�8z���F���9־�6�]Q�4�#�S�h�F��q+�l=�Ā���}����D������[�Vɱ3G�!hfB����c��O��6�[:e	=��rGL��#+�<D�Q�� k��(�'��I��<��@�<���i>a��RyB�ǭP�d�K��@�n��􀊏H�"�����$2�"�'t��'6f�]�H�	�|
�`�FU���+D9U
;W�\?E2���
+*�� ���M+��<�E�p)�)��k��-�ѥ�	Pp�a!�u�b��	�(1�ɠC"!w5D|�N^�lJ�Q���)~�`HR��0IG��Q��?i���9�X��X9/΃j%�%��̐�c�$%�ȓ8�6=���8Zj�qG���LL&�,��4�?Y,O�D�1mPD���'Sڹ��ȇk�����fC��!E�'�G�2�'t��MQ�`� F�B6`h�A�ODHڇbMq"�	��T/:����';dXZ�Հ1��X��n��HE$mS�@��pV��:��X��Q�Q�ýgbJH���$J�^�R�'��5�Mz֋�I|�Ѣ�E{H|�O�����) x��B"�':���;$�ɕQU��j�O��0�b�=^T�0Jsc]��)9��'3�Ij�`ߴ�?i���ɤ
����S���͞�#x28�@��+����O̕#���(9)�4�#�Љ)s�a���v�4�?�J�D����'jB�>��Ix5�=?y�	zA�W-:���v���U������!f���9��P�m�iQ�҇���ݡB�"�'I�>Q��2W�v\��AP?C�\s���#�&��ȓ�+T�r�A'޳+�)AT�+���>�0b�?C�Ṱ�[�G�0[3���	��� zBSp��ɟ\���L�IѼ���[�����Z=��=X6j�*x�u�V+C�Ba�R
�u�J��|�I>i�O[u�P8C�p��<�a��E�P1@�(Th�P8��O9�� ���F�$j2�$��� H
r���Nن\��� 7�m�b�NI�'�� �������'�.)3Ќ�:RBa�vC�{� �k"O�"+�9�$��N� �J�Ʌ\������ݦ)��ly".� ���jG�R�$Z�����_�-�L�h�l�2p���'�R�'���]�P���|�w�G?;��A�(��P`�aR���m��Ґ���P���Xay�D' ��u�F>��չ�+ �l
����S�Z�� �S �����ۧ~��`�H:s�̠���'�+V�'���'��O�"|�BB�5e,-��o�3:H�Hx���}�<�c�AAǖh���9h-<)8��z�Ɇ�M[���$�8k�8��O�B"^?V-���h��+(�j�r���'b��R�'��:��ah�`'={�5*�)�F�,���ҽ�`������Q�Rp�䍝8���?��@8H	zڮF2`�t/�5w�fpS@.��2�oW8f��%�4TcDyB��?Q����dI	qX��u�D_��m����a��'�a|���<ł��1E�;{b͚S���?�s�'��6�.�]a�����[�����֑NZ`DnZ`y�W>"(��$�\Y�0��g �WB��h$�B�o���'j�f�'#1O�3}��ʕF$Ft@��^I�����ޓ��ɦ��"|
�R+f�b����70�qH�R~RMY�?���|��	B.`s\��@4m�$2�KWj!��C#{��h�&ϙ�IY:��wh��26џ�����������BXPX�̌:w�Z6M�O4���O,��!
��W�4�d�OD���O�ݑ@�-1���	;���!�b��tA҅�I�	E��	�@-T6ZQB��0�ӌZ��;�O2!YlP
�.`�0���<�25����u��ON9��Qx�	�)t�1�h�y�.2�~�)Ь?<gnT.���:F"ҫ�?I�O��E�'����hX�]�%Q�Q��\��I9cb\�ȓM��`;��I�y�*%�3��0U[�U�'2"=�'�?a,Od�yag��Ij`/5L�#&�ʜ^[$X��k�O��$�O��Ăݺ{��?��O ��ȳ�7?a4$�W���Y'Ј�wf��P7 �p@G�H�Ƙ��'d�9�C�K�e�ا[�BF�	H��P3��]�\X�˶/�9@K�����jg�}0%�O�o�F���M�q�*�@g�'���'��O#|Bgꖫr6�q���(j��ͪ�l�<�dL�/���`!X�9+
�[ k�}�#�M����M5�5�O���Ѝd <M���ɥ;�v�`�M��g��'�X�ӓ�'�R>���;0X%-�\����w����C'{0�!� Ӏ_���lD�o�?���Mzo>�9�	])*�N���NP�v���!4�I.����G�0}�q	��d'�b�'��0J��1iSf��!̢�����x�l�O��;LOD`��ͅ�/k�8h�D�/�`���$$�S�$��OZ��`�@�3(,p��8}�^`
��'K�	ҟ�b�4�?����i/{��d]�Ђ�E�~D���
e� ���O�H��;�d4q%l��jb�6�T���*B �2;s�a��I�p����`~r*���8�A�az��0�4Ty>ם�D��O\L*2��F��� 0X�O$�3�'
6-LG�Sş`��|27T:Bh<�e	A��4��h�[�ş���	Q-2��� 
dd�CL��=)�z}��@̧_hVqA�eږ4��mcH�Cxy�ݴ�?���?	�̈:o_�����?����?ўw�I{aa�7[�� y��
d���D��! a��3��bjh8u&���O�'fD� 4��*���a&W5}1��`@Оu��-�S1-Y����eU��O5�'���E&B[*2����Bx`lJ���$�(Z��'���W2p1�qk$&����M��a[��C�Ɋ<�J�2c�54�Q�P��e��˓Kő��S🄖'"�#���?X�T�1��e��ؐ��+\�E���'��'���b�M��ß(�'Hܸe��<�N*v)�Yhf�
�]<������Z���Н��O�}I��_$S����Ǡy����@��	Q"�3���&���vD"4u�?����j0*��s&GT�t1PXL��۟d��t���N�X��ׄ2�L<�ЫY�/�y��"O*�9��ȩ;� ��N6?�h]k�|R*q���D�<!B�ٲP����`Ȓ�#d,`v)��GDpF͟��� ��	ßPͧ
ȱR��t6���@Kb�Q�!%��rs�ݨE1�0�'���O2d��M�g��E�&ބ8l��f�N/HH��Ҷ-8N��P�)�_�6�?9�J��� �IV~���wN�`���WI"�};���?���?ӓQJ`aa�T0	���PJ�t[����	5�yB

�d1�2������EʟԔ'���J�o�P���O�˧��(��2ڂс Ō/J�m��T�a@|���?y��S
h���s ��l�^�Qpf�&��C�����rP,����VL�d[�N���$�-%�@�G����m�W��_���?qꐏ6`���q��S����2?��
���	V�O��� ���0��\=j@2�-��%I�}C"ObqR �&�xf�.�2����I��h��a���N� xk��-�E��|�J���O���?!=F��Տ�O���O���s������j�\j�dH+/t���j�9FL���9R<����<�c>�'���c�ϠEt�А5�H+� ��ŉ�0��!Ƒm��ʃF�+b>�'��	���,�B��F������Z�ɫD����1�3�	4[��pSM�o����$�E�{�NC�)'�x�D�":�ds�J�!qʌʓVu���@�	�_Q�E����D��33"�B�0�h��V�2�F�������	ɟT�[w���'P��m>�%j�k͠&��3��dI<��sϘ��F�c1�:�p=!��̽,4�᪒"��w`��
�̊pC�ɳ%�Lp80�$\O�`I���l�������8��D����n�ҢpӘ|og�*��2J����bP#ď_�R��:0�'0�O*�@�X!�ͺ�':@F�x�1d'��@Φ��Uyr
�"�.6M)� cK7�D0ۖ��<&���@��H���59Z��Gǂ=hDj͛�`�
%�=�ቮz$#<!f�8E4DQD�й	er���UG�4����O�c��(%��WEֽ�fD�:r��T	�g%D�X ��L�HP����W�b
H�R+$�O����#�U�%�H!��2Պ��t	�H>��KL��?�j~rZ>5��l���ŌHt�U�A�s�X��韨q�
�h�^�	���\�d!;�S�O� $�Ն��V�8(��h�n�8���OZ��a\|���R�cP��}�uh�,S�XjYTδhT�.T����џG�d?O,���G�%P��pe�8^^� !"O�eX���6t�J�(�[_J�98���<�h���*��C?�hd�ȊQx���`�'^�L�sR��"�ş���ɟX��my
	�1ܖ�H��gc�qb!C\�Y�KE �P��������­[Җ����9{-At�M���\�wK�z���$	~�|9�����Z�x�ЏJ�-g�P�p���+1��O(��?�/�ݨ�h��cX����m5oC��3�'E�X�GGP�8�
�#�jg �-O��Ezʟ��>��D�͐cXLfk["`���w%��`���ɖNI�B��\`d��(�zFk�G玘+�;uH4���	=�\����:����|^����?���	��#B�=��K���"��C�Oɲ�ڱ�G�WdL��CB�n�
��$��lRh@� ��oܢ�)�%\�f`J��eE2��ׇ�Pw"�҅@F�B����>�R)�%��ϟh�|J�-�!id�C�-�D2�D�M]}y"�'W��
T�]�l���%��6\ HI�|��	@��mi��q fz�+޽��ʓE�vР��?������˳O����O4�c⇂(FK���5`�*Xn�����O���l#z1�d��	{%�mb���s�$�E Ƣ�B种M�:������$P5N�ЕmO�OH���KI <�zם)��>�('�Q?b��9�CطN��2hx���#F�O��$??%?!�'��%�CIhO�!B��_��u)�'Z��C�k�:I����Y�P�3��$�{�O~ �pA�#���ȓH�+�H;��'<�I0f������	�@���Ċ���exÂ�9\�������p�����J�+5OV�H�#̟�,�Mх��a2A�Wn�=��|@�J#5��Lp5��}����*�رN�;��IA`���J��R��?x��;�H�1^u t��:?9G�Ɵ��Iy�'��;;m�%�F�+�
h���ԅ �!�^����Z�N��-&�2A�Yla�G"��|r����Ĝ�ev$qr +�5Z}Z=`����:�0W��Ob���Oh���<�|�&Q���Hr\#�"J� ȧ&���#�A�&���ï�#h�y����"�\��pA_^�*`��LC�"�4����8q���(O�[��y����?Y�d�;�8�:p.�> HI`�].�?9���(�w{ �p�ˇ��R�ռ/���@CNȓ�+���t�@��E�X`�'��7��O$˓*����_?��I�|��+�n���牥I���T�[ȟ`�/������5�W<	�����8y� $���|�!W�b|�� #E�k�h���o�'2�4àJ�7*��eV�H= 4��@O�$Xl��m�q��ʕ#Z4uȠ蓌�dċ-42�'�1��VO]��^̈!��G�m�Y�T����a;�MzfU#4�)��\*0W&��d�Uy�m�.6�q����w�X�C�W����&)j����O��D�|R�bĦ�?9��������X�< A¨U�/�r��yZ�V��q��:҄A�4X��H�����U�`l���Q�,��"���y���+9��Eã�N�`��!���b����PM�gܧN�x��f�lnL`��[%%��̓hu�a�Iȟ���'��� � �#�^��a��<A��-��"O��b���750D�Wcހ��HH�퉄�ȟ�i)��50��m��	5e�G�OJ���Ole!I�P���O���O
�)�O|��u &o.m:��w6��qG� k�̝a�!�(#��s�g�g���e(*��"}�T�(-LxR�9�@=FO K��q��Ą:|B�+�*T�F�$�ϟ*<�T䘳��K�<�Qq�\-&�d�0"V8��YO�������E{�7O�l�ƅaܜ86:�2i"2"O࡚Gb��~����u�$���'ۨ#=�'�?�)O�%�R��)9���%�X�`mrQ��R3_H�d�O��$�O�ŞH���i���2
Nݰ�C KB���F#9\Hu���ПIZ����'���3 �~�@e!�Y��	0t�ߜ7W�M� &J�fw��&�'P�M������d�)"2�LA�g��y�����hO#>���	�g^�{B���:��d�� RG�<1��&S�PT�ND�Ĩ'�iy���L�$�<T�V}����'R8�����Gɗ��'�W��}rb�'�|� ��'(��'�<U�`�i̴���I�lRȁ�i>��gMO+b���M�VF�h�7A/�y�tyhE��:���`)2ДOܤ�p$#ʓo�2�X V�y��`��d�����Ӗe��!��_�7��g@�K��C�,(>HP�$Y�r$�a���<���$�nyb �X�,$/�L���!cz�A�.O��O�O��q~H�1b�($%)<=�8��o���O�5D�d��g�,�%�J� ��0
�iЉ��'����xR"�P�S�rR4J��ܲk<�!)֤9��4�?iV@���y�⚴8���?����<�'ŉ$�`Yz6cO")B	:5�N0`�<p޴�?�FbE�?�'�z�J��M�;P����A��G�@�a�o�z��i��F��?��t��'���|����?y�'t��E1S�z8��WR4��4k@?�?��Tؔ�A���y"�۱������4�s�DIQ!RՃc�߮<@�y�dhğ ���OT�ĝ�K��@�O����?��� B�U)`��l�Ψ�A�)n9p���.*��������\�n��T�������բ�BL2��i�4Oz���4�����?1�?�0p�[?��O+��Bהq:Z�����O~�`"&x�`i�3O`���'s"�a�����<��.�����4�FQ!�c�
6:@�(@��IE�� �U��?q�'6, ��?)\T���	��6҆��2a�8��Ez���(��lZ�uW���K�;�4,f��O�R��O|i��'��U��*0h���e�-F
�Aa��j��1zv,�O��>M��i���<��*FC�������1H4����0w^���'�����P:(i*�*Ց�:	��4�?���?����?q��?!��?��;�ʝ�E��HBD]$,3���Ӧ��I��4��͟��'���'5��'�Lxq��>�3@oKv�x҇eiӆ�D2���O��1�i��$�0R���k�j=.�4�tӊ���O8���OD��~&�h���a��$	��N�
U��D̿>���n���Q�o�by�,�Kh�y'����	ǀ��(O�b\��ӍK�L"?1��i�$X��a����u��	iIݲ94!�$� $Z��p�S�%�B���|~!�$ͦDU��CE�j�@�Z��	`!���48��S��A�P��X�X9<!�䂪#4b�I4Ȁ�
�	q@�_G!�D��P���#�oݡCӚ���-J$ W�������	�H�I?QW��1P�)��],N���!۴�?���?���?���?I���?A��4��Q6jςl�5�U��<v�=�q�i�2�'�r�'`�'��'{��'�F��mO*��F���N�t)Hmi�f�d�Ox���O2���OF�$�O����O�i@/h�|]!�H�c4x��é�禩�I㟘��͟��I̟ �I�T�	�|��a�+Gn��H���z޲��T�ɐ�M���?����?����?A���?����?�稓�P*�C�]5\���D+7���'qB�'�b�'��'�b�'X���
@�$�ěJ�j���噔D2�7m�O.�D�O��$�O��On�D�OX�$P5��)���'*֥��D��S��o�� �	���������D�	�8�IE�&Hi�.��k��a�@�P�FO�| ܴ�?����?a��?!��?���?	��!��ШD���A(q��~n(ua�i��'���'W2�'?��'�"�'�����U
/^�q��K�/t)��xb�h��d�O|���OZ�d�O��d�On��O8�" M�.edքR�e֘s1z92��˦���۟��	Ο<�	՟D�I���L��e�Q��&U�>�q�6�Ð�M�O���<��I7����Db�vDh�'/�q�7?C�1O@�?��۴�y�C*n�T�ٔ��"I�)���&A�i��d�<%?�
�iK�1�b��R4((�$H�Ԉ�)�<�I)ES�c�鈅I�XD{�ON�d�Y�z�A���V���3��TNBY�$���ܴ6���<�� ����fձ/ݶ�i�O�;������\Sy��'Z��>O�ʓBܐUR��4��h�LJ�7�m�'oИ���$>l֤��O�#J)����y2��30���W.͂~��iAUB7��$�<I���h����8F����Ӗe�tq�(#E���o��yJ���0��4�����&L�x/bT0�!��bqQPG��M��Op7M�O�Di@*q���T�5 ���e�֝���f(�>'FCe	�=:�(�=�����D4� %D&��5R��i�e鉹�ʓD�L�2ʘ'��!k���IZv��N>��q����yyB�'�V<O�#}��ݪ_�>2�f�>2ĸ�&D��t���ږ�ED~"L��|�PU����"&��'���K��6F��Q'��>O���d�'|��'�b�'�"S���4'�$`z��d�����8͑�g0YXu(� ϛ��'s�'���yE�f(l�H����7�F �k�*hڰ��nջBQ����Nm�^�ןHz�a�#K�b1�Xy��O���.�F���7�]�U+�%£	�<��'d2�'���'��ᓋ@#^�82�9`�H9�	Iw���d�O.��ݦa*��Tyy��b��ك/ĴAm�J��!K2�pk�)HߟH�'�x7������	�Ԙo��<���/Ʃ��\�V�z9��$S���'�cD�!�̙#�����O��D�O��dѽR�H��.�<g�f��S��%#/X���OVʓd����� x��';B�?MI��#g
��%O�wN��2#θ<�&T�ؓ�4sk�ƀ�O�����E5h^��7!��WȤt��o�H�Ts��+���E�<���H���Xw_��O&��Ùi0��r��T��M` G�O���OR���OB���˓FL�fF�i� ��w+�$�~u8p�̥I�d(��^���4��'�~�b��ʙ%,�R*�������S-X��7�ꦝ��l Φ�Γ�?���Å��y6-����ٻk˦����*r��JY������'P�I۟�����H�I�����O��.�Yit� M�(	PEsB�,˛�IA��yr�'k"���'�6�n�\�kF�ǋ�YBh����#QI86m�Ҧ������$����I�E�w�j�Ɍt����+ޏ�{�k�>[�4�	����`@��6m'���'�"�'Id��ĦI�8
�+q�A� �xP���'s��'�B\�|Y۴gȍ����?��8���p@ֻS��и��4��b�>�i�d7�ӟ$�O��I#/ 
n��M���_�&�>���?	'�O *� k�]�������a��+w���'ٜ���ǘ!���š�OsT�����?q��?����h��扠+���I5��k�b�)�mQ�G ��D�֦AjQ�7?Y��ix�O��	�?�ԝ;��$$&I��ˇV��D���M�ܴVQ�6B^�3��7O*��P�cz�I�0���a`�Q�?��0�Q�%o�� D�9���<a��?����?����?�d�t>�Z��>!�u���B���Φ!�m[ǟX�I��4%?�ɍ|�,+"c�-�y��g<zz���O��l�/�M���'։O�T�O[^�)�#�/�<ԡgN��J)�%�%(���C�Y�TY$���E�Z��;d��'�剥*�j�Z��S�uB	�N�tX�	�� ��ҟ������'g�6�X�D+���@X����_0:	��� A��LpӔ�D`-O���ҙ��#,��]Cf�ۆk���prg+F�!�g����ß� b�.A|�=���^yb�O=�NFԨ8a��P ��9���R�'jR�' ��'�2�:d��lv�(M���W�B�T�d��?9w�i%<:eS�i�4�?!�O"�QǶ�H��1DE�Q�Deq�`�Or�a��Gs����WD$6t���$��obx�d	7L8�y����Cnpԣ�ʁG�
 ����e��������ON��O<����A|�0[��R�y�pq�&��Z� ���O��-\�MS)=h�'�r�O�iH�%��ۑ�	�A�����_��ɑ��D�󦭠�4Zv��d�O�
���o��c\½�JI�+?Ȁ�î��W+Z5�e�����?�ʕ��#�|�h4�RC��)��|ȕ(*�r�'O2�'����Z��s�4�}��U0@ �$�	�`P���`\6�?I�"L�v�'��'���~5�f�	A>��V�-~�u�F�η{�6mK�ىg&E��=��?a���37��P��6��d�)g�<��B�!>��اdU%�$���<���?1���?!���?�ϟft�"��A�NI9�&Ф��,�c�b��qW�O����O����d�֦�ϓRvH��nB��EI��O��ܴB �O�����"��7�MÚ'E��3�KˎDQ�(�e(���1��'���ڔ,�;>O~��|�\�4�I����Io-���G�5}���������	՟T��ky� ��\Z36O^�$�OH�z�)��T�2��r��5����1�	(��$V��e3۴M�T>y��$�#�B(2��,~ѫ���O|��O�
(��3$�<P�x���cO��uǏs�4A倝;BrH�k��_�$��4
���O��$�O����O2�}B�'0"E8s���D[�Ř�b߭"��1���&1�b˵���M[�����Z�m�)g6���צyj5�b�\�?q�iO�6�ڦ�9�� Ц���?i�F÷g�q�e�)�x�Bs,Z�ɲ��"D(%S2�pL>�.O��O0�d�O����O�,u@_LڠQ���]�0\��<�'�i�hp���'~"�'��t��Db��M�|}�GWP������
rZ�~����z��H�	K���?��S��e��_?-�|Œ�'R7>�Z�[� OX[�ԗ'�����揋a�.��[y��ų��0�" ��	x$T�0k��'��'l��'��I!�Mcj��?�� �pc�z��ɒj�"ke\�A&�'.�7�OP�O�]�'�\7���M��R�^!A�94I���P#�q����ϓ�?Ij67�HI�B �������+� �Yoź/JH�0�BI"Ir�$�O���O����OB�D#�'` �=+w��7���U��.[����I�\�I��Mb�R3�?Q�� 6��<xT�Q(�#de�8�1흃3���d�>)�i�7���H�
F�mӾ��̟j�F�3O�ag�[��a�lT Pt�R�Ɓ ��'��'�B�'P2�'B�d�
� �H8De�x�����'��]��JݴFä Γ�?�����i��tH�`�ЎS*���,i�	>��$_Ħ%��4S9�������P�E���Y&@˝EJpA1��N�S��s'@�gW�Y�'e�TG��*�뮙]�s��(R�	n�q�ujW l��L����T�	˟`��~��]ybxӌ�:ME<Y7��	b͓Km��� ��2z��ɯ�MÎ�<�t�eǮ�-�\�qm�`���ߴ)��fn@���F3O���8^v�]H�cJA���	�@kF�jA$hXB	�&�hH���D�O��d�O~���O��� Z�`ڧFa27�]�aVᘄ�ɺ�M���H"�?!��?N~2�s��v<O�����)k#��ӂ`�0���djjӾ}o���?Q�O��i��&�i'V�7`�|rg�/D^&kp�^�y��0B�A���Bd,P�Cu�vGIL��Wy�'��.	 �jE۔$Q�e��� �f�f��' r�'"�	��M��hE�����O�͐�/	34����G��-:��{��7�	��$����ߴ5�]>)8'+��+[����O�l�jT��O����?�0��J]#r���
�"^4�u'�j���v��T�D�C[�^���sg(�OH���O��d�O�}"�'6~����i�2��Ù3�&����,���h�/W���MÊ�OX	b����>̋v�=]av%�����oZ)�M�!�i��M�ҳi��Λ�F�T�\�9�-T<��1m� ;�x��I��D`L�b�|"Y���I��������џ�ˢ)�#t���pFa��FYaᄋVy� }�@VJ�O����OB���|��(�ҒB��P�3]w"E��Ɩ.��I �M�ĴiS��3�)��,�	��`�V��`,�<�I�6f
:q;(C�H�7QR�&����$!H�u4���<	%���yl� ��5��)h*�?9���?1���?����D��%
T�U��<���#%��Ep��"	s���˟h!�4�?YL>!�T�,8ٴ*�ւ�O2���(��0ə /4`k'a՛Y��8O@�Ă ��15dh�˓���w6|aB���MP&�hTjT&|M��p���?���?����?9���N���T�|�H������'�r�'��7͈S�˓ �v�$Ƙ5SVa��	�?:T��'�;?�f�D�>�P�is7m��j����f��	ן�/�&��� `�G�u<��Y��*��$ˢ�ez�%�,�'ar�'�"�'w"��D�Uז1`Ol>�Er2�'=X�H�ߴA��h����?	���	H	\��4�'�Z�I2��:�'��˓�?�۴Yor��T�O��l�2b�,�	C솧FR�(OͰ!j�pȓ�\�z����?�ۃ�@뺫W�|o^�]�X "��$X���;��P1i���'jb�'���d[��޴
f܁a4ꇘ߶�	�����v��?���Kr��$	W}2ajӐ�b��8\��Q�!OZ��u�o�⦙�4��D*ܴ�y��'��4'@�G>���^�|cdϙ0����b�?�z�3������')�'���'�B�'���C]�p�T�S��l,bl�*XO���k�����Ο&?�I;�M�'~��i�j�S�@@ ���mĴi�87���<�'c�D�O�����:ԛ�8Oڠ+��?�p�&�sc��he�O�S�O}�఩4F=�$�<Y���?i�g<}e�����؝/,�a�._4�?	��?�����Ц��r�l��I��U�ބ:�U�'o�3
�Y1 �f�S��4�M���i�����|z@^%&��x��%V�5Z���%�H蟼�I�tEr 	%_���'I�DA�����<�3��e�tD���U�<����`�����쟔����F�D8O=�A�,\v���@j<����'~P6�@�~����'��'"���.>��i"XQ�6���_�a��y���o���Mc����M��'��.S=t�E�5�A2v�`(f'5<4p$��.��!�>�3��|�^�,�I۟����t�	ğ�E���3G�$�%�6L9(�����zyR�lӶ`� 	�O��D�O�I�|J�z"�8��eX�<	^���g �s���I�P�d�ٴo@�f��O�H�i���\�o'r�eq���]�V�PN�-a�@���H�<���ѽ5���v�-O>I+O�-##�=5��i4W�s�T"��O��$�O:�d�OT��<���i*����'�Rl�!�B�l���hP;�m5�'�p7m;��
����Of7M�ʟ�+F� "R`(���-g<4S':!�7�x��	�fr�=C.�$7���'/�t��� a�ݢ4�^`�F!Lf4�<:��'!��':b�'2�'�>驇�P7H>,㷣��V��P%�O���O�n�	Q��`囖��]�ƴ�$�ҔW#���t/ Z���D�>Ӽi�7���&�Y�d�p��ퟬ#�!��	L��Lv�T$���׳B�����c�;Rd��%�З'|r�'���'��H(��.�$zԢ��g�����'��U�D"޴<,�Γ�?!���O.����_Ɉa�e�FM{,��.O�'z�6m�ɦ!��ħ�t*!�.��uE�)U,�pGl�6�r=��)߅SN�8)O���_�nB�]���~d1K#�S�d��,y�D&tih����?Q��?��������ʦ� l䓡�AL�n	�%͔S�%�T�������Ѧ!�	i�����֦iJ���(���ReHSwX�5S䀜�M�"�i��<���i^���O�H�V��)Qς�k���<�C��?��呦�R' Q��2�eK<�?�+O��D�OV��O���O*�'23��&� �0�l��Bֵa��ڴS��]��?������<Iоi�ĉ%fo  �b�/!T}�BX�2y�6�¦�@����$��V�i��� ������V�:����@��C.T��	�c��5���K 
�%�<�'q��'�XH.옵��j�1�hD����- �R�'�B�'d�I&�M��"�?9��?�e�-1rX���b��t�d��h����'|@��?��4t�Z�l�'۽I�^i1���/Ji#��O��Ē��a��^˓����Î�uW�t�dA���U� �A��ː��A(bC�O����O��$�O(�}:�'4@�k@j���1풰C�-���V��FF��}0��'�b6�5�	�?�R#� H�8s��82v�b�J�ӟ���4=S��`n���p�tӠ�IןȘ�*����m1��+��p5cVa�d��i	Gp��$�ܔ'<Z����'��'ҡ���$DzvO_�G�\��� ��6�M�� 4�?��?������qL�Ҥ�K�RmK��A��m�gZ�hR۴>�&��ON���)��ʠP�-Ԧ8�RYX�H��d(�"�,Ȑ� $�<a��GhC���^wBP�O�˓T
X��$̙u��+�(R��y��?��?���?�(OT`n�)����J�ey2%.l�H ��H
��ɣ�MӍ�>!'�i�L6���P0�_��f���'ڜ*< �#Ɉ+ �6-k���	�X���h��'[�����`�t�S�Qx.<�v�,@�t:��'���'�"�'�B�'8>�hb\�"d �1BGH�<���xwI�O���OެoZ��"9�	��8��4��'�,z�)U6�f�OK7�R�E�'���,�M#p�i��D�G)ћ�2O����z����ǅ�8R �B�J�($�t\��Q:k!p8�f!3���<����?)��?90�I�&�!SŎ�j���փ��?������Ʀ͛���ğd�IƟ\�O܂	zRB�aL0�ǉ�d��!*O�=�'��7m���99��ħ��`.��&\`䞍>��x�Ն^5�Bx�$��Cm��+Oj�I��u$�](�� "�r�懀C����D 1���?��?���������̦���'�h���t�F� E*p�� �Zm�'3^6+�I����¦m��&��A�d�9/�\�KfC(�M���i?� ���i���O�`�sl� 2���!䢼<qҏJ�A_T	� l _>�,��(���?��b�<6���[��E>Y��y��Jlp�Ӱ�X�Y�bE�ŅD��y�MH2�$�Q���H�z�J��ǈ�����ʁKZ��)�,�B,\� HM&�t(e��T�
@����$�2HJ�Yh|�R�&�aj���aC
`���8EGT/+{zݰf��̰��JO�M@,%s���y_�Dx !N�s�&$hD��z��b�dȐK�m'o��bPJ�-_%l[޼�5�޻k��Qz�� �n��wgϞW'��[�m���0��O�d�d��d͎i���bV�1�����T�\�ע۠g��b�J�p�!X�gʀu1�e�� �9%���W�����!�]�z�6�҆�)�$��N�.����$w��p������`��Z�f�f9��=�Y�j^�B�|�0��.O�@ßF����$ʲO�l���^�H�h[�V���[���2g�� �	�F�l���Ƈo1J��b�p/�eST�2O���'S"�'�L�:�)�$�O��dz�йc�S�M�59#�]@�b�C��j��mZ����	�O$�I%?���������0@��fɭV��WME'|�F�I�,���C|y"T>��Ix�I�#�0jMǎtl��H��F![���'��lp�����d�O8��O�d�O����[*��8�gX�i��񥇇Cߚ�d�O���?�N>���?����@$�Щv�K*]�2y �A�%�(����b~r�'\��'���'\zI@��'��8�OW'j���� Tgr�Ȗ�'���'�r�|��'�"¿IdxÆ�HR��P
@lL�R��Ѳ!��>D���� ������I�`�C��f�$>Orpb��O��2�Ғ����(e�'�B�|r�'�2&� rl�O���g��1E��sՇV6)2���O��O��D�O<�bw��O���<�' �@��e��,���B��}5D١M>I���?y$j�u��T�<�'B� v%DdEH9*��=F���	ɟ0�IԼ��	П���ß����ͻ1��ـR%ԑ���
vf6q���͟�ɓ$j���h7�)�56�8)b�j� e����/ ���D�$��n�埰�Iݟ��S����|�����B5!E�I�G�2HI���?wK����O�D�1OD��?j�A�3@(�\������v�<�o����I럤A�������|B��?	'.E�j5�}A��I�LT@����$�O&����W
1Op��O���1����/����˃@1G&���O���p*�~�i>��ȟ�'��'�Ұw=�,��Y�D�:!�'�����'�R�'$rQ�؊ /!=Kp�q�I8�T��$��9����K<I���?q����O��>OL��!��:B�,�R�,;�(�%�d�O@���O ʓ �����Oh���%E���i?4h(O���O�d�<A���?aƅ�~z��^<�*��>T*(�4�hy��'���'�剭C�zMXM|jd n��x"�S�!�hi����?���䓿�dX�q���S�Ŋ8R��b��8�@!b��'���'��<S�ĴiI|���y�l�m� ��A�Z�D�b�cK7�?�.Oh���Ot������O4�c9�a������!���-�X�D�<���ìeq�&Q>=���?��+O� �ҳH])SǍ5mY ��'���'�r�(�P���ß��3}ªL(J��,P6�\����E���?Yt� �f�'�R�'��Dm �4�~����
+|�F�K�c�v� 4�bM�O�lh5��D�'W��y�'cN�JQJډ.�\����K�ʔ��t�����Ot���`Pĝ&��������'f�}K3��Le��geѼty*D�'�B�'��L;�y��'���'�\�iB̟n���wD�j�$R��'!��S�w�FO���O�˓����<zF- 6'��n3�pӪ���$G1O��D�O"��<a�@�1:�DEF2]�谅�
�_LҜ��.'�$�O��=��<)b���: H��ek˂o�����Ѥv0���<����?�������V�
��?F4� d�A�7AD陳.߽AV���?���d�|�Au����1!�qa�I̐wͦYE�A?�ƌ�'i��'�"R��i�N��ħ.�h�p�,	�SmƬ��c��nr����?!M>�(O��i��i�V��X�s͘`�BݣK�r�'#�\�`J�W��'�?a�w�zX醡 �>e"��u��T'dI�L>�-O��e��|���3��d��gY5(��V�Ο�'˄4�bx���'�?��'a��	�S(qb�n��!;���; U����<���XT~ʟ�(��t��y3�#���krr%�G�On�&��O���O�d����|�}���#d�}�Ȗ�L�g����t�$�"�^r�S�O�BkF'Q�}j"���8�Xd�5&��'��'
��sS��������<��ӖI���c�6�"�jҁ׼!��b�؀"�C�����	�<ɡg
?	z�}��T~�$�f��ǟ��ɬ$Mhѕ'��'�B�$^�mN~�Cޙ)���듉�*l��'>X�O����OH��?ѕ(�
�䵑�ЅFI��j4C�f�֩((O���OX��"�I�<)���q{b�\�vA���1�@e��D�X��I֟4��Gy��'�.H��7��<��f��^`  R��)~BIZf�'fR�'���Of�z�/�/X�h����Y��5�& �
��7J�<��?!.O��B�(p ʧ�?!���HT�}�a�%��iQF��?����'��D�?j���8L� c$=��j���`h�Җj�O��D�<���(W�P)�X���O��iG�+.���c�	+��E'T6㟸�I�yΠ{�
&�?���,G�0m pF�sܰX`���<��|s�5k���?A��?a�'��$�X��x�c�+A.xR4S�N��?��l��3����<�}��a��
�� �ծF��AZ�����,#��ȟ��I柰���?Ŕ����'xI�ahO�#H���Th�v�Q��'�Xd{p�P�����Z�X,tĉ�"H��� �ӧ�ac��$�O����Or��&�<�'�?���y�G%~��U LG,2��Cf�PN�:��<�u�Y��䧤?���y��7^:���G%pn�B�c�	�?1��D��*O��d�O��d)�	��:�F�1?�RbZ�}>�ʓ,�4�a�v~"�'bS�,�I�̑��� �z�2��֋	8��V�^]y�'&��'e�O���&(���"FPw�R5���C�o� ���JàV��I̟p��My��'R���0�l���ؤ؞��64>�;��'X�'�B�$�Od��'B�İ�ӱE��qD&!Q��N54�<0iW+�<����?�)OV��('���'�?�H>�a0�挭H�^��'��'�?i���'L2���Hn�@�H�|y��$�UB��ˆ*P�5�r��O���<���J�A(-�����Or���$<�9P'�M,[��݈F蚂|��X��p��\�W�3�?�{���mנ(�e_�Q.z��I��`�aA����\�	�?A�'�l$j��׊?��ԍ˷w��9��V����l�Y��$�)�S.Y�|(0�i�����'�ѡn����\Z�����O
���O����<ͧ�?�P(X
?��=Ӡ��[�$�V����yb�A�rղ��=����+00p�R�[��8CVjϋ�\Q*��?���?y�ET!��4�����OH�ɻ�0\����*�D� ��ʠA��@�&�d�
� �����OH�	�����L\)2�z�����d����O��c��<i��?��ޘ'�d�5NY�k$| �&ۀ88)O�c���$g����X�Ijyb�'�^���;}�dcf�UO�BJ���Y����ҟ��	c��?ab��#6(���s���c��z��-�l���?9���?����?�*O� `���Or=�D�n���%dR�)<��@�O���O���!�������CDx)|-�"d�+Ɔ��.J�_�V 2��yy"�'��S���I�Ā0��������^HJ���$Y3��Y3/�|)�P�	���?	��\��QD��e������u��z},��-���'����|���G�D�'���O��� �	h,�����Z��7�d�O����͞�p�1O����Ir0"�F���1mA��ȟ,���\��������?}�'�p�uCL��I%B z���X�H�	�n*����#�)��;7�R��=v�S��V�E ����7k����O~���O��	�<�'�?�K�j��sV'��$�>�n�%5�B@Am1٨�y�O����'�R�'�J�����^(�X�d�6!ε�d�'��'KҠA�E��i>!�	۟��S�? �x6O���4	����>4x% wQ���'g$�����'*�<ONL@�(F�z��@���,3��'����%�	�����ҟ��<�r��y%0i2bE�8l��Y���^yBP�hN�!�O��D�O�ʓ�?�����:�@D"���b��t�P�BX#+O*�$�O���.�Iԟ	f$�x��))C�H�3�`�4�����q�&?���?�)O8�$�h��瓭E݄��¢B�8��Ul��d�O����O�����E�hdHBG�2.�|I0f�t��m�hJE�F��'�R�'��ğ@��
�f��'F%2)ǵq�D�2iz��:��'���O���"��K��
���ݲ7�FٹB�2U�0��ʟd�'�b)6
��ߟ4���?Uht��m�P4���L2T��U���?IUHD%�\�<��[y@Iv��+�"EP��D)��'c���CI�'Hb�'_��U����Q�W�9u�Gi�t����Iy�'��Q!f�5����O�Ph���S�<q�QZ�̂�M��+��a��?����?�����4�F�d�
B.X���S�>a8�HW4����	�hOб����Sҟ�q4ؽ?abH���O0��`�؟���֟��ɾ�ȕ����'�"6O:����[�r�"y�nB��A�K�$��'��-�w��4�'�b�'���ŋ�7�`�h�ލT�t��u�'�ª�n��7-�O����O��Ě}��0OT�.I�oh�)�͉{%���_�T)��-?����?���?!��?�A�'{n虊寜<~.p���D0Bb8rжi���'yR�'�����OD�!�~h���$g����Un�(��D�O��$�O���OvʧK.8�[ �i�D#�G��Y�8D&�7K���z��'���'B�'�BW��I)m	d�ӝ��h�!ː"�[g�Y
�4��	Ɵ��	����	ny�dA�4��'�?��K�'.|X�Q�,~��B�M �?�����$�O����O|<�T;OX�$x���q�+Jh0�Xai��V�ۻ�.�O^���O��F�H���Z?	�IƟ������:TkV�|��8Zb�Z�>���'���'Ҁ�Ov瓯u� 9:G�h~rA�4!�{� �$�<�V!�� =���'��'���ϧ>���΅�yE��5�.*VhE9�?��?��o]�<9��?��aG���On�Y�`��	`VtZQgU:O�Q�g
P]�5�igb�'K"�OC����d�	R�XlFg��;���a� t��X��lڢ�'���K���?A )_����:��՝!!�L��n����',"�'�2�zWB�>9)O��f�d�WD��=Bwa�1\Xԍ�`b�<q,O�h�u����X���,��ℷ.ɔ����ޡI�\�%���X���:�����4�?����?���7��s�}�DdK9����w�FmTLB��ҟh(�"@"K�J���,�	�?]�	ܟh�O�8=B@i�[���Q"�K2~�Mw$�lP6��O����OL��J��S����*Ѩ�7K	6Ig@!�Ek�3\9�`a`�d�I���	Ɵ,$?M�b���MKǏ��hЇ
	*hsNx)��V��?����?����?����Of�C�<�H�+V�I7zcX���-(N��r�!�O����O|�D�O����O���,�覽�	��qC!6;� 8q�,�"c4l�'Ȉ����ן,�	yy��'�F�ȚO��'G�4�f@��X/��F�<J?���b����'o��'L\���.j�\���Ol��,�!AL
,�4)$��D�F�c�O���<��p#��'�?�*O�	L+�H�[R�T�(B����D�v7����ON��E�,��o�����L���?)�ɶ6��IX�J��p@�G̊�1X��'2b�3;�'�i>��O:D"2�
��Z) �H�bg�����F���ֽiG��'���O �d�';��'|&�����f��(D�	�+�b�� �'��p:'�'\��6^D�`�S�?�X�mӝm%z����FY�.�S��&�M����?i��m/���?���?���?�E��6���ǖ�~\��!����d�<Q�AD~�O"�'��f˝)�����e̞q��Zak��B�'�nt��E�>y-O6�D�<q�w��|QC�pH}�aD�24"*O�!��7O���O���O���<��$Ęv%��'��:P��CLP�.Mdȩ`R���'<bP���	ݟ���7y���b�*V�L4�j��p�7?����?��?�.O`��Gb��?�اַ�,�C� ��X���Op��?A+Or���O>���-"�DW�=6\��),f|�X���ʜtR����O��$�O����<i�X�OU�O�����O^དྷB�_�}���:U�'��|B�'�E��y2��L�uoR3g7�T��Z�gL�����O����O�˓&�t�����'��4h=OK��@"��٣���O��'���'�I9��'"�)�O�h�0��m��Xњy#�b��?�.O�(	�,�ʦ	�OWB�OAP�}QrH�ħ ?ij��p�J]A�M�����I�*Tp �IU�)�9�x�q`�G9^|�,K@(G�T\2��?wޙo͟��	Ɵd�Ӆ��'8^ ��Y�lE� ��7q������'����'+�'!���$�,�@P�9q�"juNJ�"	^�l�쟄�Iş�s��5���?���y�j�S)&���ǈsߛ�X3Ad2�|�.��Td�O��'*b*D�f�t9h#C�!�-1do��"�'ƖH��>��� �'��
��ŉ1 �u��a
�-�:�'[��Y�'��������l�'D0��B�>9�d�޺{´B& Z.#��O��d�O�O��D�O�� Z4K�J��oh�+R-��M���d�Z��y�V�x�	ş�&?1pf#�/�:���0*�Xxb��� i���1�PUy��'�җ|��'���zW�d��Nn}��h���2���<�� �	ߟ`�'4�r!C3�		�X0��0mي8�t�[0�H5v(��$�O��O���O�y��m�O��W���/3t���Dƣ{"��Iٟ�	ny"˜�z����蟨�	� �7�\�0`��8x���C�'���O��D֝{�d5��g>��@[�|̀�`"�F��К�@�O��@6AJt�i���П��S��䈠��|�`QL�����P�C�B�'wr��!%/�Oq��E�V�.p�$�a���;=ɔ�RD�'&���"r�^��O �D꟪I&�T��-3 !Y n��r��DǯN��P�� R�=�Ih�IR��O&��/p%t��qˁ4�ڬ�& Ӂ*���n���<�	۟4##�\'��'��8O�C1eɀN��Z�녈3Z��$�'V�'����&����'��'R2H�b�P� �hlAA��5+����'��B��lO��%�5k�$��ET�ed�H>R�y�	⟈��(���ן�����`�	qyR���b�J�g�̙��e%C�����$�$�O��=��i72HS��\0nİ�@��"f��r�M.�?A���?����?a�����m2R���c� -�r+Vp�nU!d�F�r~��?�����O�� ĥ�O�E�-�m`�iڅ�~$ѐ��O���O��D�O�ʓ4?4)�A���
�*�0�@���-�\�	3�I�fEb��uy"�'�I�;����N!d��AI7-K�#4<�d�O����O��d+5����O����O~���DY�T�X�,ʽA��0Ww��O����O�� 6�N�6�1O�ɝ?$���ce�O���TlU	�bY������M�.�����歖'8�X�AO��U�]
Ѳ�iN>)��C�����L������kE~[u�N�<" ��O��QFE�O��$�<��'��<�� ��tL�t���-ޔ�Gd��?�`!�0h�A�<E�d�'�\�gՌu � (��.*�L+��i���$�O��Dًm��1%�$�����&2�ݠ�*]�6*hQ%\�7����?��CT��?����?��O<)�2�J��6BP�K�4�?���:Qf%#�x2�'B�|"%�;G¦8#3BUv�еHV ����I�R+c��I��8�	Ay���D�bDF�H�Ah��C��Q�"����F&���O*�.���O(�d������M0���1S�G'�n��A�+�Iϟ �	ӟ �'��35$�HYA0�[#`�np�p�V3E�{�[����џ\'����џ0ⵅ��l[�ɋJh�i5�G Fƽ: ��<���?�����ٝY��	$>ua��aEV�J�,�xx��(������T������(u/���QK�)V@��jGD�P�T�ئ@�O�d�OB�O�V��F����'���b> ��� ��Ј9�����'��'b�i��ԟ@�g)�>6b�"$�לZ�f��'��;ZmH��ݴ����O��	�ly�L Ep�:�
\؎A��l���?	��?9�g�b���O��	z�L�#�Х��
��F�����Y��y�f�i)B�'y��O"
O���i��F�!{���)s�]-M�t�ٛ|�"|���fXp�C+ �Of�B!��)K%��{w�il��'+���yOR�d�O扥A�|�h���P�D̑bI)�����2�؟��IƟ�j��$��8K !ػfTv�C�NK��D��4 �]pN<����?9H>�a�+����#�Ӱ|Y���E���ĝ�b�1O����O(�D�<QR헽Il�cug�v�@��Q���X�B�[�xB�'���|R�'��J��M��Cտ\� 5s��~� �J�yr�'�r�'?�Ɏ��]��Y����'J��$��cX)vlq�'���'E�'���'����':��YA�ȹvyB��Y2��3.O���Or��<���# �O(���m�0:N$t�
�3�  ��'���|��'�rχ�'��E#̊�a�^I�ê�Nj1����?����%l�'>�I�?��e�_3[��Ų0��y�4CKN�Iݟ��	&B�#<��E�.	s̚a�$����[}�|���py�ۅf��7͡|���ڢ_�T0O�U4py�^+UV��u��O��$�O�x�)�ӐM��y[Wܬ�J�ܖ
�a���$i�a��iB�'R�O�O4��ƈ4cX��0 ��77���/U���نX�"|"�N]�@�˗�\M��AB<-p���i���'Kb$�1To�O����O��ɬiN�][r/��85@M@u��8S����Ұ
5�����	ҟ`���� <[^��q&_?���jt�ӟ�ɻd��}�I� �On|"hג|��D��G"u�SK�S,削	�c�p��͟��	ퟴ�I2Bx��C$Vg>pjцYh�Va�D�U۟P�	��IΟ�%��	Ο(���@,M(d�27*��T��<iT&�7Z8)s�9?����?�����dX�x�,��"��CҎ&�@�e΂�R��D�O��$�Oj��(��"H)�	�t���S�B9Xv��I�Bq"P��'�2�'L��'9��՚6��Ο�`7��ZLҭJ���#��T�Iϟ���n�i>���6>v q�ƍ1}
� �y91l�|,�asq$B�p�>��!�'���'F�	;]xl��������O��il��e�`E
�Q���A��:Y�V˓�?)��?Y#�D�<�*��Th� u>�y	1x�#!;� M�q��Or˓Р���i�"�'���O�&�\�2�H���	;b|i�0��@N�Ds��?��T�lϓ����O�ʭ�`B1x���B�.6Nr'l97�U#'��:A<���SET'��Yw���OS	%�� �%h|��B����z�dP?p��| Q�O��D�O*��,���O��O���ʄ����@'!��� ��J�6��7�T������Pm�4���?���y�k�'A�n�*A���Ì�J�Z����4%���2����=h/�H�Sb�I�Qj��Y��׫^4��C-��C�I�tҼ)Y��)$�R5��Y��.�2xȄQ��K��O���J}/UH�P7��i��yh���j��	 ¥D�z=;�u�$i�	�;nòD`�*ٮU"Ra�͐����Cv�I0��]�d�a�v��UF���&H��0��ɦD���؁h�$��+CƜ�����8ة�qI�O8���O���ẛ��Mc��I+����I�ed��s��,6D����� ���!����A۔D�OS����[Y��%(�Z��+ܬ��5�g�q7��#Ai��Mr��K�D�i��`K>�`[�4�rQ�����HӾ��ҋ�G}��J��?	���hO�]�
��9B����d�1'�b���n�u��)�9F��e� ��R2��!�$��|�����_�~�l�pni�^&e_fHzB�
�|k�=���'���'�r×�kqB�'l����EX�I����[�Jы'l��f:�q�흤vV��*Y$N�x��W�Oy���v�U�[	�X�A�_��|���ˆH�|�g��s���$�H���"o��e������K��A�<E)RcoӦ⟌؋��'�4�Q2)��;��p!	ɖz�L�	�'�xQ3cG� ���Q�
B�'��7��O�˓T���xfU?��U���^/R����'T�8�sw����k^�?a��?�d���F	��鋄D��Œ�����WW�vM"E�ĨlA�M�6��� ��D0A����#JDT=j����
?�P�݆�h	G��F���$/���*#=1di�ǟL��G�+�|�Ä 4Ѯ�hgf��j�������?1S��*t��P$@��7R�ˢ�a8��JM�<h2��9r�.��0bM4 �&� �$��85A��M��?�(�p8Y�-�O��e�
�F�N.9{N�z��T�km�5�P�B� @�P���TMԁ���ͺc3�E�O�1���DQ ��ţ���$2�T%����M�r$#O:%�Gղ3ټY���%��	�$�O�9�\}��'� v>!���n�J��@�'&�����<O�<��P�޶���c�0���`"O2 ��]�xFN�Y��#J��ܱ��	��HO�)qӨ��A�:�&���͇�*-�����l�� j�8LcW�џ����L�����|Ӥi��J8�UK�	�e���Q�����V�+"4��D�?�@���	:O^�[0&�%)�I�!ٻ�5lO�l�£Rn䨃Dhړ_B>̱p�������F����I���<�����dH�#�$�ʀ�,srа1bֱe/!�Ě!T����߳-�zl(�JI�婏��|�-O�=[G��*'Pl#@A��t#f��v�S�]
Z�B�O<���O�$L�m'\�d�O\�&,-�Թu H/��Q���;v\8�;�ʭ� ��R_���D�^�'���*w쎤qT1гm���)F��5C�B���G�
�Z�`��Rx����҈>���i�.xh&��)^��90D�_��f#�d�O��i$�i�?���1H�3
���^�!�d�	/�]���	�����"O�M���ry��[Px�7m�O��d�~�cB�[$ q���b���U�Ï>���Ѕ�'��'D�XI �i@���6Ϛ�V�46��~�(�YV`�i��úY�T���v�'�d])�¤V��J��P�cކ����Օw���돜����ۑn��[v$,�#cе�I'�MK���i����E�M��ZV��%`������O��"~��1ith�۳@�W8TA:RI�7z��Dx"��O�'\[���pӰ7M�(�f��B%E�L�`�bO�?��\�L,n�Ο��I\��ɉ�2��'4����.>@�Y`�O�?��QT�3����`���*�� ��wL,�n�W�ԗ��};�8W쓗^(	P��I�$�nڱ/�P��1��15#v�H�Aޞi��bR�6��C���� ��;_Z���R���2���Op�dhy������5>���b�xC@�h�0�~��'�'�ў�IƟhb^�y�½#�N��̅�f�Q�x�ٴ1ݛ��|��O~��2�� "ꋺ)~1��Z7�x�������->h!�M����I�p�]w�"�i!��0�F��r]*Eas�V�(�ְ:d��֟�Q4C^�R�H�iKܡ��HO�['6.�d�1#ȓ�@G��p�+�>�?�`�� #��)���6��3�6�N��F��BE�1�����46��ߝ#�dk�$�����	ӟ��'9`d�%�J!q�R�EC�?�{�'��Pv�I.|��e+��)��Qq�'it�;��'j�	�[�@�١�>F��D3�)��HT����#]�D�������I������E����	�|���߃I��pk�� �H�&_%oA#ԮV m���ۅ�E�QR(U*
�K�V���K7q F�⵨Ű)�R�f)��h�
�%��0g������i��D|"�Q��?y�lg�P�P*��"ز#s$��#�aAa�x��'J��T>y ��¨<�+3	�!!lT�s�(5D����%OL��)97嗻�J<��(�����4�?q(Ob{F��V�T�'�SG�"%�A���r����B�� zDE���?!��?��"ؘ^���"�ɲ"L5(vdɸ>�)d���E΂��ġ���>������� )TW&͈�CM�mND�3�
�I�8�ZEIE=�x��(D�Z��0�ڲC�Q�0#�o�O�imZ��On��J͡_�m��$u��)�'�'�ta@3k���b�Uh��P)�)��ͺ5�Bc�$K�B=jm�2����v�����i��'��ӭo��p��埴n2F� ��A5G�� � �!
z�S!ܓuT��Ǌ�n���2�Y�(��c������=�8R)�qk�O?!țV�E6ĩ����|X�b�1�$����ȜS����(�H�[�ȅ1$T�i0��im�����^���I�<%?M��D}A�	qH�y�m
t����y�.�P1�yԀIU��L3�G�(O,Fz"ol�7-�lޒ��2 ��B	��0%��6����ʟ�
�h��!h]��ҟT��쟘8[w[r�if<�D���ye�9:�� x6��{g��)�t�t���E����'$��)?�Y�8墠��6J:&اg��rE� �$��8���2W�ߚm��BE�@x�T�I�<�)Y��_#~�U��cN�J�4���ɩ�M�q�ir�OX��73|틗���9)Jd	b������Lt��D��FR��RB�Ĕ'��Yő����B�yx��H���* E�9�b"Y�S�N�2��������Ol���O���O���z>�+��190ゅ�Z;<1����V���d�P�Rz����$����<I���ɴ� �U2&��mcd�ͮI�TuQ"��X����-�ayR�D��?��"� 	�ej��=�n��)��JΦ�i'�i��O�	D��;2r�
⧂�c�.�"��)P�jɆ�\��tH1?bY'-�9~bf���InyrGғi8|��?᫟p�7�<u���)$ݬF��� �O����I؟L�	�am�,��o�$F�R 梓�u�����LP�[ (8� T� �-ar��J����ϝ�Ք��êY����K5�ND@�']�[	�U� kK=瑞�!��O��$4�T42�(���k����	�f�	�L��ɿ0.h%�E��:M�Wiǃpp����Z�d�%lN$�@�;g+��r��Z.��X7j��=�'�X>�����������A�Ȑ)�]p@߁F��.�:�P�@� T�7B$����� ���*��b>7�Ue���A@�5��C����NA��P���иCo8M�d9�����@��b���YiŃ&�Vm(�jJ'�M�`˟cش!�)�i������C0� M)���P
Գ4�~ńȓO��ы�iژ=�45��C�b�Dy�)6�1&�֟r�X��G��)v����-Ѷ4C`���͟�zD���M�	ǟ(��럐����DlZ08ܶs$O�&{�<c"�U�S�ʅ1+�-wՆ��l˩��9�i�?=ʍ�$*o�������^��У�����ei�>F�K5M5f��hZ?U�p��3[�	���>A�n+\�9WFA .xbP;�d�a}��	��?A�i�4O(�$�O�"ɴE�ƈ��k�i�A)�<�,���'	��~�PL03�Z��"���Z�`"��ŷ��6M�ȦA�I��M�����'��陚N��	�#���L�%�HQ:�A� ߿ 4.���O����O�h��c�O��Dq>�8cf��X�Yx����`
���	%lF�a�'LM�� r��'�2�j��ο���DVB�5k$�G�=� �F7k���	�D����G�' �d8"G�����o�J^Ƭq�Ʀm�	Xy��'��O�,~LȻ���{�Qa֘�<B�I�6P��R�5X�%@E�io8��*S$��<�7
׶R��n�O��d�~JB� &���ɠD�_Kt���ښ$��p�'G��'�. ���6mق����M�n���G�ꎜ�1ɿ[���ȓ%�|�'�8Y�ŗO"������Ah�شg�����'�<d욳	_�Q��d%`��x`U:��$���Rfӆ�oZ���O�UJ�ң.!�4����D!3�:��7�)�矈���˖Kd��i�#y��M[b)�O̥Oؤ:�i͆!5�P�	)tp�$�O4�ѦYY��D�<�矠&�bӡ� B%��(4Ɵ�\`��C1"1��p<�G̊��5���I9k��#��We?�N�'a@�e'�"*�4M�ӆB�':��x��ɚT�:M�Mǅ\�P���']^���ıNND��O���"�'2��VZ&C�'A�-C-�'G8с�7t�$
��D�H�8�'�3�dכ��1��&/A��+
��� �!�$kVF��pQw���~G�� F"O�\���X]��1I�9$z�0�"O��f̒3�	�NH�+K����"O~��W�D�)R�H����&>�u�"OBY��$� D�t"1J�&?�|Q�"Op�;���9|��9v`�'�}s"Oh���.TЂY��e -Y���"O8U��OI�Q���
B4a8���"O `��E�0,3�P��k�4Te��rs"O�YKǯT�(��|P�	9P%���"O&��i 9�\���0l,�+g"O����&I��X�9@I�-U���"O�X���;�t����*��\�"O�]#e��D�i���H/�Z�a$"O�+Bl�\�����IV�R0�y��5.�<" ʂ�uk��C��4�xR�KS�Й�g���m��i�&�&rI�� %.�	{g���Z[��<�7H�(9t���G	X�:G�8O>Hّ�֯i�20Z��;Ś��4N����U�v���{��$%�$C�M����KT�gl)I7�
!*˓Q�1�����(�fp�4�/76�����$9
�
�! a��p�Ee��N !�C"�p�ԪP�`"��B���(D��L� E&"Z�67��a���t�ɒ5]�u�UB4'F��c	C�J�������'m��3�ѐ?r~DjrO�|>����#G;9)�cG&"�D�󇣞��~bh	:82�?���R�_n���v�_4c�0��&Qt�'m(5Е&H�m��as&aL!da�fRn��a Ao�K�F���S%�i�Ƹi%�8Ai(`V�D��I$���d�����d���$#�p�I�0P=�6;49�&K{b` ����u7. KC���d�T��ʗ��9TI���ؾV�D9��	+}���5��0m�͙!+t�.��h`(�v���xG�R![P�� �Ǳo�ٹkOu�$��@�ev �։�7U
����Q�wy:�b�q��=Aԭ_ !peYT���~�#l��$h�
X/@�U�ڞ�A��B����� �^��	��P�P����Y*pХ۝��)4ؙ�_s&���E��8S1�l�:0��{.D�4��xw:OVd�C�<�V,#��ϵt�x<k�!D�9�"(�u(��d����);c����iX�|�ˎ,y���&�!,O�Hpl�P�c��A=w�0M���o��ŭ�2Y�k��R�, �,�L�R� 	C`%@�w�(e��΃ªT��-�*�����EU��YA�
E��$K%ؙ�x@7G \����G�OR�|2�C
)כ�d�	5�
���	J�K�b|1e��%;H�@s+�l��СԎW�i�SD���Ex�eM�p�=iF���1%��<cbY��ig%�v�1a��0 ��q� lee�V�W�e��Uq�D��_F-�V�дi�t�X6���bH�u�%�Tjoy�&�V�a��u1��q� �b�*T�83�"w�8�U�T�(mt��b��0�:�.I!Z-Bѓ�6O�h��p�$�b��,d`�����230�Ag�^�l|���o�9>��+#әv��١'�O�h����;078�y��ɖ��V,H,P^�j�i�MÌa�'Æ��`�E+��u�4l��z��5���	�\H�R��[�OϒI�G��?�zY��� {(vE)�iհ�h��cNW������əO��� ���u�����G]b��sO�1V�zdRul�>GN���?�*%%�G&T���sĠD/E[l���O�P�f@,<Bx�i"���[�M�Q�l�8����3i-t�!�ˑ^�m�oF�<�޴>Jj���`ە>gh)�rn�'��1����h�]�s�V�)��m0�^�+4����9lxۢ��$��-�1�C�m����Ɛ-1ʠU8�H�+A��!�@^�{j�*#�<44�T�E Ԕ���4�d�yV��G�H%"�@̻�����
6�����ғZ�*��Uo��P븝hS��#}b6	�e���u�Aչk-�4�(�X�'�r�q���3t���d^F��o�O
4��\T��0�ŋ_�f�3��j鋥%gZH���/3�b�(ba̅FNp0�͇�I$����M$�txD�ҨOx�4�_j�n����~��6T�_���Ѧ\�#�ߚi�R��uj��EiI�eO@2s�����X��JTF'_�Kـ)��hr옟6m�e�&$\52��Dy��J!�� �L�1f�I�VD�|�cΞ5JT�a~� �Gؒ	�m0L��BX�ph��Gt�)� ^ʒ)r$%Hdt���X� �Ah�8K�Hk���@l�` �Ɠ����jԳS��Ua4Fމ=����+DɺZ�?��@p��$Tt�t��O �6ԩ��7��1;��/� Y�-�?7�lk_�q�h�����M�ç�l.��;� �OЙYwI�vv���c�� L� �n\��M#�n�Zt��p��!҅s�.J���D�g�#(N�H1b�;0절wa�p����`,�uG�;v�}a�� =b�(�Qmƃ[r��KױH���uwC,=���� ���,�0�j
�	nIPБ	�j��ٴ-\U��`�	M�!^44m�"�n���䅡!����	�4��s� O��u��M��� ���	<�  �Z�(d��*���áM��i��m ����Ŏ\�k�s;X�R6�ەn#�Px�I�(�p� �Å-c-�q��BΘx��+�r:X�:"�n"�DP���AYt(��&�#�2�9b��6�������ĝA���9w�Җ:���@�/�_R�Q��Zt�:A�s�k�Q�)�6��BN��1�(*�*ҚN2=��k�.��#��!r�$����1(�0����5�>4rWJ�K8�uj�z u�Ĝ9��Qj[�����W �?�ӊO�p���K�i�r8EMĝ;��ia
V�\��I��]�5RR�:Q��/��1$��'�Ё�)P�����Z�WK��!",:3YF��'�� 	s$��u����s!��'�J)reEH7/��c6�ȏ9:|
��T�UR�d�2�йb��ذ�A&#�\:�Eɴ)� ��S�? J	k��G.I>^��T���:���U2@�d��dŮK��'�b�����^�>Q05B�}H0�zF�V8���PD�ʖ]x"m3	  W�~=��*�AO�h�Ň4$�0(��?���I/>��=����X��4F�*=�," �k����#�Z�XJ� �=�ag�3���'�CE�;��u�q#��	�Wy��"��@�4�p��񏚳3v�����.W��q�g��QkfƂ�SU����?帗#�cm6�P�e�ؿ����4R&�qsw�3F�آ��W�h�d{����sO�%C����-�z5�^=�B� �=�� �0Y@����P�ȳ�B'8��)F�!qΠi�'��>:<T�CНa��1J'l4zZ��뱓x�X�i����"��
=���/����1���-) ���`�Mf��T@a�ٟa����� 
�:�	C�M��,[􌗗PbT9���$nx]x�l�%z��q[� ��(��&ׄv��./@A�A����y���S�i�̠���D2��Q��r���N����R�����ш�(��N��@��\/�P��q��Z�iW�,��S<�)�CQ3"�k�ό/��ɒ)0P E�Ҽ2��,�!�	�ɲ'Å�M���ߘ=V������	h���长f��Y�j�0⼌�@ G(L�P�s޴K3\y��&�6�R?6��lTڼ��6��*�KK�a�-b6�:[Sa �#g��DB� gb`��V�2�k���Y\�|mY!����6�%W[zY��㊚�j�8��ׇ'Qbt
%�ֶx6��y��ֈ2�viPB��RQli�OT���d
�H���NC�IW���?4-;3�֪q��q���Оq?
��3C��69|�R���A
�8���ɱH��@�����!�H��@
,+pЭ�dMQ-����A
�Oj]�P�7`��E�3��� ��4�ǂW44��!b�̼y_�d �#�;�x��͙#�Nx�u���S<�s,��c�ȸqJ?Uy�΂<��ԈN2��|�3M�O(�{A��=�n��k΄;��d)�.������۴a6~�Ѱ'z>Y(�ǎ�y�P麔�/�,��VQ~�в�k.K���i� Z.n�%>c��b����	�xa@�K6W�2���m+� �j�
�(�|{�l�*{�ܔz�8��tI0��4Q�,��7���2�zĥʋ7J����ʚha�ON)EY���!�)Y:�6 -���!�}"(˿z{\��喌/}��0g5v�:P� �Jyb��"G
yBx3��ݶ���AW�*u��P�GD�r�(p��-�v�b�o������=<���\�V�膬P9��'�P���ѻzg��m�4��%x�/Dh�B�rĳk`8-C���y6�����,�T�f&2d�(ȋw
� �Z7m�b��pj�l���M�OUб�3�@e��q�d&�t<���9� @iv�Nl�a�'�0IXʅ˓��c��7�M�+.� p�Ort�b��ɏ26�;�(
j$��DX�����EV�L�p��&C;�?������@�j�R��O�s��}#@d/ �s�,�qV�D+7�i���U?�J���w��]c0d}�aZ��N�.�$����KW�U��ŧ������DD���
0$����K�1 :5�%�1l� 2�-�)<���x����?;R�s��EԘ���Z�b�����)2d�,&����CU(6mX�����!]��9���/vv����,�l ��� [�I�-�d��@� �H�F�V^����h l��ГT���� ��W�@��v�§=
�OB��&`�%9	���<9V<�O�`}ˁ��ՠ���o��t�B���O��6��渳��/R������N i����z��l�;��@�`I�1v�	1���M;B�)")��fO0*r�±dYx��M�X2.�NY[�k_�Y����&ϐsՐ���7&���e�kl��|�5K�jm���~:Hٛ�({J�1@B�|NA��#T=�tax��.|hg�?IDzҦ´A��!��'h����¡Vm.@;�*ޚai�m@�&X�o	*zŖ|�f��m&B��6Fp���C8E�(}�p�C!a�&p��G�:%t*�{$�2ړK L� ��)�6剖	?n�Ω��n�u��|�g�:.j���D�7��UK�NL�r�������>!�u�O~�Ȁ5�?��hc&!��/|P �y2a,,z\8��L�Y!���=�sf,��S�m̅&L�I�G�ՉM���1P-�>Q��t0r��|MJ��D��'�"�;�D�q}��'��tX�ߪ\�$��V�Ã��m��N$���F{��	R�O� �e
[3Z��y']��&!�TaO�_�����s�%Z0���N�<�D���5�hAvN�=� 8��f�a|"�  �� � �~N���q˓;�$H&�Iu��Ё��	*�4��s�ɘ;�8��Hq������'�D�IRkΑNQX����`A�k�b��`Ev��S�W%��� SA*#Æ�S%# ͛���T�.t�@��Q�>iHH�X�B�Ai��U� `�!{7~Fz���m}l��q��7�d=)%K�
��ش;<�����S�����%Ѱ%�t��i����+-_��&gr�i k��qa�AJ��(U�A���6�E�/�L�pi�
g�t����-�(��R���8&,V�3����R���O��:�nZ���� W�L��p��+����=�T����4]�Nڌ5�����G/n�� keH94�IC
<��Ox���l��\��#��F3�6<g|��r�c�:�Y��+h��OHq�q��!u��i���J' �����U���$����]p�䍁�*�k'"T'�V�O�Y��N�*Ch�rc�>	M�"=�V$иu�2������ ֝C�m�&iJ��K�9����;!�A�v�O�4���_9��'�8!���C�N(&�S����k�^$�	��.lôB"���޶�iR�Ǯ'[Ʊ���C����`mJ� �`�e�:|�� ��ɵ(}�4`�--"�h�Q�A�E �A)%�D�eRH�Opl3��P�a[^�P4D�=h���4G��!�pu�&�U}��� ��t�U��S�)�R�O2p#�q���l+.f�0{@�C�!gB�'P��1�ǄjNȄ�S.�&ˌQS��̟fn֘1X$;B%H�(��T���]c^-pN<��K�T�Ƞb���bE��=ᔂ�-�vՀ��ƁG�fy���6J!�9��h׍Y�b@4��#��M��1/�xɸ�&�)T-*�@�&]�{�����P���j���ui�#>�B/�;@��L��j��<Q�$N�E��z���7��pKK3M��x�dH���1a��'��񑍃�l�)�1o�,�:�����o�$�C�Z�BeB�l�1�!�͇m�"��)�1P�6��V��J�R�{%�8NP�AB��_�0<Y��\�"d�Q�b�v���)� �t��M�<O�XsHɕfQ6�yNlT����D��7��XaF��f��h���M�8G�`�	�gP0�I�n��iX�4P��˴PHh}Q��"STX� t\�$��̈́�.�Xy1%��9	P�E{�f�;a�!�h�	jh�`�#�!b�ơ3��Y0Z�,e� f�;b2v
ܺi���ቌ܍:��@�,S�y�o  �h��\)19�=! �y�d�#@�FD5@`���\� �a���q"
�����?��J�>g���OXb];�*�,H��p��Z\�|���O.�� �0�8��h'^����^�k�U��V����Ƣ�wx ��Ǉ����dꙄ5�X�E��ܟ
ܢ����b��z�6O
�k�i�;�N0au��M&Լ�3�ѻ ����EQL�E�⍊<��Sb)���T 1�D�I�R����"m^�*x*�A�i��˓x>��@�]�"�I�&�:�O��
g�N�%%x��nŋ&�5�����,r"��(k�B�(R�ߒ�f1��0�
�+�!��)�U�=2�p[�/��S����I¦u�w�/bm�);��֒>KX�kP�ze&����1T�T ��)��Q�b4B�&߷h��%,�B�����A�(U��ᢁ�0��9*��@���)�rEK�,<zM\!fQ�KahXa��q, ���F�:��rL:|�� R�˰})��JÓb���w�`P��k��w�Taf��/ۚ��,U������e����m8#����ѥ�-��y6荲*׀�kblޟX���';��(
�(���É1Y�D�R�O.��a��`�\��G�y2��>jfY��T�W�l P�I�H<��p��K`�}A���? p��ԠC�/����q�$�[!�'⨁�b�Ԡ�����d׳T;���p�-�����%������t�VTY�
�a`r7��S2�у��
Q���p�D@�N0�8�d&Ob�((E��O؟4�A'^�n+�������A���B�l�G~�!�&��x%��K�i/v�DY �'߃i%����"Y��J��TDv�	�dH#>���pE��o����OP��0=)���6���'�P�ڕ)�>�Y�C�ϓ����G��Z��Jу�;��y��[�~�V���)�6�y��N���Ԓk�\%��L�0j�m�+M(J0azR�7ٺ�����$��|��n�|Ͱ%hE�+$��ze	�j���U�L��"�/$T���W�$̒��6P���qƗ:����=1�+��l���u�V.Ѽ���ń2���Fϟ�Xj��� �2�f1sI�2���@�.^��A<<%	�&��4��A-���	����rk��@��=.L����B;2=!�F��i���s��'��h�7�=nP��t�<Q�/�5'PhIq 9b��S�m@5U�6Ax3�E ,�+&�Z=�Tϧ5&T`YQ@ҹc�'���c�*����ǚ{FZB�B�EI&" p�ìjf��9�U HG`��+Q`Y+ÏM�.��y"
�^ǚ��`nϪ=��!1@ʘ�0?0%�P	���PJв6Q�����%�`0��M�<Iի��j舑�J+A�(�qF��J�<��͑�����U,�l e)T��G�<9f.�����E	�L�f��h�}�<�G�j�&40#"v��`�"� �<�`l[�\� �a�EM@-1W��n�<����O�&ŋ�jߔ{� (��%�k�<)���8���iQ�<�]0�dl�<Y$g��f0��ʋ0��u�w*_n�<yu!��zq�,
e�8���o�<q� 1Vg��:s��*�r� �e�o�<�Q��t�n�pL^���0��\p�<��-�+�P��
�w�0��fm]r�<Y�"��9�\��geU�[lY��e�l�<a���&
x�Q��A�^�ʭh�e�n�<Y��^xB�0�ϖ8�α`g�i�<�񄀡^?�]�g��	z���sM�r�<���0=�a��!J�`2F�l�<	�k�$���-�^�>����o�<����F���
�a���tΕw�<)sdV�,@"ق玭���	e�W�<��L�o�N}�ufU��>�	�O�N�<y���4G��y����AO�ay��K�<�
�ҵB�cI�-6�Ԑa,�{�<!���4��Q�c� Ar���ƐO�<	wh%D��u/��P2h�0GnQI�<I'o¸\�����㗡l�D��Q��x�<�t�^MѦiGN�h�1؀An�<E(@�r1��ה_SBE��!YS�<��b#94ѓ�J\@\�U��M�<�g�7\r�aՆP��|-3u'�>�b�(1�dx �X*<����	NX�'C@��1��/w��S�#E�"q�l�	��� y;���^�N|�WfǀF>Ҁ�F"O`�K�� 8tH��Ǝ W�M�"O.��$N�\���T�R�|:�	��"O��ّ#�
&6+��� Q��-��"OP�")P�
x|�3띊���v"O���R�Y�(v���9�4L� "O��p� A�Ԝ2��n
$�s"OT����B�'�<]s��j��j�"O�aAu�A*c� �UBĉf��x�"O�̩��Om!����ǈ.j@j�"Oȩ���͆Ej�i�)�` �"Or�Ӄ;`t��)�ȗ�M���
�"O$X�wFv�<�9���L���U"O�9Q�f��g�$�[�Ɯ5�p]؆"O�U�(ĻF�z	�$�պ+G1��"O�<{���9S]ڕ�dIǚ93�䘄"OPM;@��8��p�5�(��(p"Or	��͚�g�<�I���w�؀ p"O<�J�95dl�����ֈ�6"Ox �6	�̞l0��3e�X9�&"OP A`��8l[�e�%��	�q"O��
�H[��p�
%I��(��"O�$�b���a�M�$�M�z��"O@�yg����
ܺF�!Ej�)�"O�9�.֔t^�8Z��
6.	�Q"O9�i�����2/Q�g�2�"ON� �)��M;��qǍ�0D^d�"O���Q��L�&!
��66$���"O���,"or����	����"O�t�S�~f4���=&݉'"Or	`U�	�2T�࢞�!&z��"O�A֣�?%ע���Ǜ�}I�"O�x��)�V!�CFB�#�y"O�y��+Z��1�Ĥ�;4\
��'4Z�ar�Y]�i���/�)���ߒ[p4�5�֭b�e"�ʙ"kZ�,�W�#j�(��'�@qj�'��;D��0�lV_WRLHK�de�Ɍl>����.-���u�8���t:�=��i�@-�*�;@�B䉲)���[3�L���R�A�bH)�D��us�ł���\�S�V�Q�Q�H杭:d�бFˬ%�D�/f�B�I=r���nB[ip��eł	1���@�Ē)qj���D�pl&Ų��1O&�2��)9I�݈��?�zm´�'&�%�r+ޗO���þI$ܔ�7�Y!C�U �n�+I�����F�x��5p�PT`v�� �,+�j����H tB����:*��P��B�	넥�Ć����(d��I��=)�<\XC6N��i��P����'�"�����>pt����>Ш(�A"�K̈��OQ7*X����@�K��h����ގ ��[
U� a�&�Zrd�y���I�/�:|�'�y9N?��X��f�+�~uxe듟�(C�IC��i�����p��L0w���@��2Q����� �"�$3�����-�(�.�F^�qb� \�l�:0m@�=�>m���<��4Qq�'q�A��A؞sd1�WL�7#���&̐2U� ̰e
T�f(u@I/d�	
�_�Pc��..P�Eb�����@�āN[��b4*��D~@!	�%V�q���O��@�[�f��Q#Ea��V���
`��(�*7V�y�
�Ͳd!�26�vY�"m�& ��%�|찤Mʼ� 0��	�\,#<���/MN��FD� ��:v�A5��ؐ`,�-!̤`H�@^�gt�Q����BL��:��|��� �!A�J��R��4H���ԋ9����D0�(���w�P��MV� �*y�T�F�W��zp��t�Jp��5HzT9ρ�?�3�	�]�E��OB�r�\C�-��	&����'Q��pt�$�%�$f�&Y<�q3 @�0	,��a�Ɣ	CN!��J�73�I�ӫ>|b��o���|��6i�	sT��bnQ�|�81�c@�(�t�����&��O��r��0Lp�gf�`-ʐM�,sx�=!P��~�^�	3���6Lˡr��[���b����4Kϫ�0?��遡vmN�QT��=]f�A��͈h���>�H�AUeG`Bʬ�l�'�X�M~2�j�1z�q�#]���h�$c(V��|�����1,O�(ʠY��q��9Gf̙�n�'��,ڥ���<�qlǞ�]���L>�5`�/K���:rQ6tZ�2��D8��a��Y�xj��L�f�rZ��!A%q&"^�f��s��Na6Ygbb5i$��//*�Ob4k ��G�*!��!�FPYկ�?��R��-p�r�b�>��K`�����(j+�Ԁ��8�0���G�@�̍���'� �|h��L�.ܡC�*0m��X�	=��
p��Z�ͧ������=z41O�A����va37�Έ`M�H7F	�:�`!;ee�l�	ԀT�T#@���sV���,��'s�N�	��Flv���"D
p�R�0C�D�0�n�R�n-|�B�����re�EO�Y�ؚ����*u@L�/_�~pT����Y�Y�T�i�1��X�P�<)�(=D���1�OF�*�\���#SX� �gF���踐�Wf���#���	��UE[�[��ܨ�N�$�,ɚ����q4���OΝiT	C&�"�D�}�$c�udR�s�
�l
��� ��*EF�B�	?k�a�0�ݺv���s#ԛM��$ &J�ڬi��B��览�e��D*� Q�e:~Ny�S�1D�px�M@ ylr"KT�O4�$���~�h�3"R}�E.�8V`�3ʓ��h��D��8����6nc�Մ��.���*4&^�Uj�H�`.t9�G ϵ4M(�p�-K��a�c?�����&N��Ш�A���'�Ѫ�Q�\��A��_?x��i��t�m2��kwę�^�ڝ��E(p�6B�y���#�K�5�(�ǒ�<�8����"<� /+R��K��,�ɯOx�`E�k�A	g���C����Oy�H��?����� ?f`��H�_.&��v�2_����U�������
��O¤B�Ӎ]Evm�cN��	� �p��7�v۱��Y�&���A�t!�X3�l�nE0�ӷ.c��*UH_'N���R�'ת��C�U#y)��'�J0x�)�.,|��J�aC�I;���g#�M�pu�<:B�����'=��Q[�H�	$�^�	��٪]q°�?5+O2r֙�6�x�Of\�ٲ�G5PL�)���Z��,ɳe��m�|UAA��l��D�M��W�<j`Q�tR�d&�z��Ӥ*q�(��$G%!G�� ���9E�IL�O�:({6�	"�6ɚ4�f����c��F��Ɓb��Ѓs���q3��O
Y�*�:���z��Y������'����
�C��Ea�OP$�/�~�[�8=
Xۆb
/w�$���0q4dH橘�;���v/^R8��!��f������=,��<����$?T�²��$�`=�'�qRa�r?y���'����<�'0�b��Ǡ��d
��BG+h!�Q_�REr��FX�1�4E�4� &P��afJA�
)LD�@*��?aM�>&&�<�O�R��V�DR}�G�3dq�9D�d��R�ϕ�0=9q��~�i)��\ �x��9/n�,4d�`peK ����7w�B�N1��- ��rx���u��	��?G�h�$����Hh���� `��RÓ~�U&U�~`A�*�p�B!�bО`s	�'��� ����yP֕���	3"��$;�D]/�?�mMj��1#��]��"�������)�	W�P��&�]�%\��$��Eh<9!U"�`�A�KEaA��3LB��R�"F �9t9T�L�#A$�'h�$��V�v b��TA�'vZv��D	K�h�yRI�6�v��@�iQ.݈��9,���Ž^|�gE������M���3ƚa����dʅIz6Hzw�FYl�Ƀ��'�l���(Gr�\��o��7�I���L��.}}<�[�o��gaj\:DbϞi0�����3��H'Z��R	pү�&��*����4r��%!� �y�CN�R)��>Ѡ�>��M0�Τ�1�,:`0:����p?i&�<v����É��6"�Ux����(��H�z�i'�>9T�>YR�U:��i�O��3�N	50������p�H��g�	m�Q�0�X}S���?����ߣx���j䦏�-2|��a@�
�<�Od�07ː$G���d�(�xpCYl�d$ڔf^�>���ԣ[J�ai +��tsr��2 �.T��~��Z��%��G�.L������RS�|	�aHb<	r%��!�\��2+5jhڰ�Վ`���6Ņ��y⩖�M^��3}B�x��݄~
P 6jH�!��zD�R�~�D�7�F�kh	8m�i
pEC b�:`A�+A� ���"ɏ�@׻�鄝|��S>-�d�5� x��e��>���P�pXQ5�7\��'��(�!�78����]�|q$�����M�Z�|p��� YF��0"'	���2A҈Lcf��1yYHArA�I�S��d����Q2qh�a ]��hC�˗U@�H	�'C@��r�6"�ڠ����Y�H�D�I�=h���d�'�n��B���'_H�dΧ%����֧���� w�'���Y$ŋ�y��d�q�	�ٲ-AT����\Ɵ��%�2�H�'��|���1{O��@W��5�b	����{�'"v�;b癸^h*A�}b3`��W�� ���}R��Zԅv̓=Ҙ�XЍ.O�<���k�H�g��>J/�����' LP�B���:����Z�"~��rK�Q���U�W�̤�0�ҽ�y�&ڋJ Nx ����$��So��;_pZu���_�u�L��3-�|�i�MzI"�N�}�晦���F$�
z���j���j$�zR`�y�����O� ȼ[���a�9P��5L����	?roVA��bI���|
�)����v��<�й���Q�<A��'H.���)PY������EΟx��*�Ut�!`K~y��ɓ�Tl��1�݌����¤Y��*C�Ims�@�G� 7�t�@	�=�$�ql�RV)� a�����d�x�8:� }᥁ݫ|V���ɋL�V���E-%�3V�z�:0�V�E0p@b�,�eBT��_%�}x��X	)Z(E"&C�,ؠ=D{��G)>���;RJ�6
��R��?a��3���F�#!�T�A�!D���0FB��µ�a;uz�kP��O$��%!L;^6 ��T�W�F�����-��f؀@��%�H�O���>	d�N�(�bLq`���ML��S[<C� ��2�����z�0t�A�D��y(/�Q��gH<e�l�'C)î�hb�&ړ���BN[~reU3[�l���ģ&f�C�J�>o�\I��3H=hf�\$-a~bkM"�X���D)D��!l���?-V��d"&?ybc]3biX���L.i����OD���Ga�2�J@a���`��(��"O�}c�;[��LJ�;D�Ƭ���'�\���cކpx��PU�擯9���{f0�c�@<f���Ǚx�Z�{��ر��>9v�ٳ@��A d�����PJ��8�|{kP���dS	eB��U������$���=���/����7c��n�ўKg� d��Y��ta��/D�n���� �<H'I� �x�	��V��x2)��8��*���5A���iDN��ڈO&D�OD���������RB��#̤;e��PM�,�y� R9�1s� �7̊������y�n�%ܘ�
o��^{��vN��yBLY�5Sf=�����9�Q��,�y�Qwb3#ay,
���/�y���/n���[�v["�+�n�)�y�D �U�֩;�&�m�H��䑰�yR�>��(#1b�`�FQY�m��j���$/Kv��t�T6Ht�ȓl�8���D��4j�I5��ȓ[O���*-�Ȝ��S�h���{�(؋siP\����6`��s� DJO3^��
2��Xc�<�ȓ�&ĳiL��x��Wj�a���
j������Rg��zl�
t�>D����@�N&Jt�e�L�.�Z�b��6D�,�mO�#����VG̉R��zq)?D�����$~Z�"�1,���
E& D�T)�`W� ���9HT�رb(3D�PQ�捊5����`�@w�ࠈ1D�Xb�^��<(���S
� �%#2D�Ԙ䪃k� �u���:D���.D����H���&,���ʶ2�H5 �J-D�؈$�v�D�"ȑp"�Qun.D�<Y�M�B
�e��mE5��p�Ah?D��@�n�'L��`��A�8����1D�V�P�[ "_5��D��k+D��x�C���@-c	�z�h���3D�0��B	m�$y�í��A����A3D�@CM��a0�m���ϙ+y��	5D�$ҦK��=� n΂Tq�H�4D�pٵ��%N>xhk�Ë�=�!ʡI7D�0�$�K"o=��K&XV"�A�� D�h3��F*L�1 NI�c'�U��l D��q n3cu�"a�-t�qq71D���H�,"�MkS��7H6��v*O�@�3Ŋ�w�00t��&���"O��s��51m8a��#k��i�"O�QX�/�Wd���d+
�>P���"O�Q�J
+	f���ʗ�<F�
"O�}�&�Q�ش ���.=���"O��i��5�t�'�F�[.��"O� r�.�`��0���cD��ٰ"O28�*�5*t�9Zq=@�{"O��X�0���%D�7-��hc"O��F
�\�4a�s�3Y!X(�"O� �\VX �1��p9��*O�����Mz����M�T}K�'�8)3�T� �
�+pd�N� 0�'��`跡\�o3�A��OH�>t-��'1�	�%D�yQ����J§UM��;�'��DA���y���[G��	T��i��'l���զM'wo���M�S�6i�'�Ҩ;tb���3��L�.Մʓ)q�襫�x2D���TD0y��@�d�է�a���Xg�.�,ĄȓC����CBMf���i	"%�d�� �t@�TK���Ƶ�ŋ 9.�p���H0�O���L�*�;4N͇�o�L��(S�S����hǟ%5\���L$=#�#Ih��3�B �{�~��ȓ?6R\K�K�6����F�4��ȓg�D̘��D��"!k�  �N���F)�0��2�Lmµ��%����ȓd�����Z�i���3��CCl0����D�Ɍ�Dz�M���%���ȓeQ� ��	Q8�#��B�EZ@I��+	䤐�/�q	8�s����bC��[.�u�P�6:�ұ�P̗��r��ȓ��p#�֭FT�d��&+~��ȓ] �!pD*@���a�C
�#����x}"�wa#����š4������0b6���c�tY�&�lal��ȓ_�b��@-��d�& �$ٻT5���w�(��E�6�h�P6H�3]��̈́�3��y�f�4	�H @*S.+�e��T�8�G-����#�툥o�r��ȓ�J��.&1*�ۢ�7G�ه�e9���3O�P1����싪Z�<̇ȓ	f0��W|�zu��!��E��)�8��"�V�Op�8��S�J�Ą�A& 8dC�Pw޴�ġ�pn�̈́�;�P�������A� _���ȓP@�K��8�,a��5����� c`m!яV�2L���AHݪF�jP�ȓ�hg��"�Ҁ�e�'	���ȓ����v'�E�R� ��$Y�L��ȓ���Ul�A�:�;�m�W{r���yp��gJ�'L�8��eP�[
h�ȓ[����B�<�niQ'@�M�"��X@�i 7�܋l�Q�fn��4��)��E�B��'%]?h\Pu���t� ��|�VP��ζU��Tӄ�ɇK@����(�� r�F)����:S1<��%d��e��M^0�ā�:���ȓD��8����L2��:ea�t��(��{#EȢ�F�X��ϻ.`��� M�u ��� r�"�I=<�dY�ȓΒ�`3J��0<TdS#�i��p�ȓ^A��{���6�T��cϞE�,�ȓ��iA��΃H�Z�����V�������1�i�-vҊ�� B�!�ن�vF��ai���B�A�"WNv��{�d�rSB��C�P�9L����ȓN�&q2�;E��EA��>)-̬�ȓ|<p���D���eBO2QS�1��S�? �Â��;�|IÁ֑���1"Oni�	.�y7�� wHX6"O�H�j˫� �ؠB�@���b"O.ZU(M-i,䋀A�8KF�Xp�"O(��M�@6���� >0~��"O�,�Vi�/����Β J���s�剀�HO哓+h��xB�ȯ2Y�	qo�3E�TB�s�Fh�3 ��0��U �)vC�	�P�@;�IT)l�9�KJ�?hC�ɲN�z�2�@M+0�0}��ɝi� C䉎~��,��N@�M|­�� �9i�B䉱G�,��S'DȪɡdKX6߼B�I#8*�V^�!��P �f�=m�B�		[�a(G.
>}����f!Q�bS>B��~�0`V�>�d��9 �vC�
/��Ys4��@H�dx#NM�X bC��4ED�к�@Z�]ް������Ly&C�I
QQDxPF��z@v��<WC�ɼ������O0<u��˵��?�&C�	!Y��`�@����0��m�7{�>C䉗aQ �ӓi΅w�
�c�'	\) C�	C��Bq���irdA���B�	�AN�5ZA%V1A!60��"S�ZI�C�I���e��蟚���'Z�C��5���i@mħJD��ғu��C�	�%��|J���	ln Y��O��B�	 ��h���c`��%L�1�B�9]� �R��N6.'80����!#PB�	�VE�d�@a��cv|B�K�FS<B�	8l����IS0Lk��[,B䉺<^:�+�E�\t�QSe���(#�B�ɑV$\�"E��4�����5z��B�I�>U(�i���Qw�]�sO/��B�	8hvX9)�ܺ|X@)âL@D�zB�ɫCiNiaӊ�>r�0�+�^�(�<B��b+�i�4E�3�:����B�I�8|�y�c�5_ �15��E��B��%^и#� W�Ei�R��Q�E��B�ɦo�Z�%��~��O� b�)D�t�ѡۑ/i�Ԓ�'�-Y���z��(D�Ty��N
J&N�Ґ���a��è(D�`�7��VpĘ��R	a�4C�8D��B�EE��iDBPW��8�o6D�X�anR��j���捿 ��y"D���a� `���!c���TJ>D����O݉Q>��!�)��V?"�#K8T�4�g��*@tł�TB�p̊'"O �3 �P��@�Ad��x�q"O,��/K�U����� B�$���'\�,@&+]�:� �
ԇu�r<!�':m�c�.-�-k"d�[�����'��D@�,�3A����aj�' M�I�
�'ܰ8�@"�F�a��3.K�Q��'1��kR&��{��A��8(���I�'g�LP�O�b=�ـ F�� 궩+�'+�3砀��qBpiϕgX�R
�'� �0�� J�h W�ƿ=D<Ȇ�((lugH�2Sh<˖�>����ȓ!G�4�`*V!<xe�g���,F	�ȓ�l�s���8FRxx�>uHu�ȓ\đ��J;B�Ӑ(��2�\���.lV�R���z����ƚ+<� ݆ȓ\��1���&!��J3��Ն�<2,����1,~-�FD�5`�\5��S�? .�Kˆ;xBh��kѭg�N�{�"O޴���YN�x퐒*�b�4��b"O�⇂Z�>TL��	͑~�>�e"OtГQT)��\��IZ4GJ<�"Ox�[CҐ'������8~Ϧ�+S"O���a���X`}[�7(Y̒�"O<QA�#�1��4hD�mNR��6"OH����O�k!�t�V!lE�"Oh@����?!��Q�����8`"O~��'"M֮D:��T�W41ɀ"O��҂R̹&�D B���e"O�
'��L���)E+/8��P"O2���Η,3�bxу(L%2։��"ON@S�
�t�X�"�K�k��5{�"O�1��f* 9E��$�n��"O"ɂ��Jh��q�qNը]
��P�"Oⴘ �Ԙx*���N,\#*�i"O�ms��4�h�#bҨ6iI�"O�C��$=|���'>�Tp�"O��s7�&���7F�A���"O:��e��F�#���%Y�F���"O�l8!���E^nirE�^�|���3�"Or<����=:w��:���uҡ[�"O�C��_�?�Q��y��4��"Oƅ��&3�̕��'\=3��"O(l��>	�<�e�<
X�=�"O�Q`!�A�$j24ONm
��"O�G�/�h��u�@��a#�"O^q�P�^�[e6\a��"G"`��&"On�t�o%TQa�gW_@�a�"O�EQ�<�H�j�R&<m��"O����¶�P|��Xb�P�"O2�B�iQ�v��#�,��,�f1��"O�0�QN#g4�p- V�d��@"O�P��Ʉ@:t��u��0����""O X�q˖Dc��buk\.��!��"O�u��
\�06�=�%�@4j����"O���s�ՙ3�*5�,��6m����"O"�@M�	� (KS;<MJ��"O��˵�_$m����1<��2D"O>�O	g0d����59�	"OUӆ�� R�:�����2�1�e"O8���ᕑn$:maG�K�)E��Q"Ot�jH8�\�1�E=�U��"O\+���G���*��>(0=PB"Of��1�@1.~����	n���'"O`�B©N�NRQ�"Y/ g�=X"O��#���O�(9{V"܉R@}�r"O��9��Ѩ0�B�K'bߴp9Z��"Ofy#1��DB^�+�@	D1J4��"OXaԫI.v����R(uM�I�F"O�8���H���bf�ĔJ��c'"O�`�N��\��RȎ�Y2�S�"O.A���̽/�J� �Q�^�P�"O��"'��W�����7>���"O�T�J��.N:�(�˛z�PT"Oe���ͤ}Ҹ�I�L��/�hu�#"O�-ڥ�T�M+�1��E"r��	؁"O���EfT�0�̰T�Bo�d�A"O8�(2�ۘFu��@��K Ar���"O��J��ăG<l�1LY�Z�`��6"O��&a�0Y>�d�m�Z��T�s"O��!���&�`K�K�;~��1�"O��(үF� T��J��;��M��"O� Bl3�L*-fY�bK�|����"O����j�j���%S�8g"O舘U�P�c0�4�T+QA=�"O.����E.0��@ē�]#��Y"O��J��s��p��#��I��"OM�W�����S�"��`b�"O�����Y�=��JS�K3jP�c�"O�V�I%��,�!��f2S�"OTP#���L�R�D���)"O�$�@�L<��2�9 ����"O�����=-��ᰀ�L"^���r"Ot��/k&��4�	�Pt���f"O2�BLλj\���5 	6n�TPQ"O������5KQ���B��I�"O�L��m+9��8S�#�Wi��q%"O��;%AR&_�R�����y�2"O��ʒ"6%����R9Z�# "O��7��u���#Q��O%�"Oܘ:uEU�<�1���(H��"O`��� .�<�r�M�K̱;C"O&]�DNZ4H&�(2��ڦU�"���"OZY�7�ȜN]��	�|�>��"O4�";;Q����&_��1"O�Z&���^i��C��E�q��jC"O���"*G��z]YA��`����0"O�M��M�*A�mh0���C��ae"O(	 ®�]�b5�� 6b��"O�%J,[�kɆ�a� � Ha@"O����ҾH{��Q��؈A�^��!"O���D��*yv�	V�һ��AJ"O�h1ՠ�2w�}ؖ��yP`�"ON5) ��n$Ysm�%o�^u!'"O\��6i��#4\�Y����Z,�D"O���@F�#��P�*�,Y���+ "O� 8a��d��[���"O s�둜!�LE�4�IJ��B�"O$��c�~n�TÀ�ԧ<<�9�"OH1�"@޺�$yر�#RR���"OPd�U�H"8�f����-qޞd�B"O�TpD�"jqB'=e�	�B"O0 �ͤvF�Q���S*a"E�u"O��gF�r�J�#�Q ��"O���T� �v/HH��3d�;���T�<y��ai�< �hXb��P�@�N�<	�%�ZqdUF/4�|��QV�<�gL	xN��w�K�&�X��i�V�<A"�Qq烛�&��!B��K�<���Yvup�K�wȘu"�[�<yE�Ú5|�]�`�7t4%ڷ�}�<�"͕:W� �T��WP���l�u�<�AȺ�j��
��&Y�=���n�<��!�`s���s T�d�<!�_�<yjQ�l��k,v����o�<�+D�k�mЕE_#6-�ps�j�<	�A��x��M01�σ_n��葢L� j����Od,�"�2���[�a��!'ح@&"OT�Iӳ����1J�Y8%BF�'�!�$�4�ڀBrI�V��� 3�S�O8�<�H~
��$H��0��A��NWd�;SH�Z�<T�;^+�� e.
�֒}�Ҏ�V��?A�J|����am���ٝC�x�z!-CR�<���vh���/�Y� �JA�Yd�'�axRa�M"�ʃ
�n����O�yR��?9�Dy AO��d�V�Hd���y
� �9Juo36DX��C�ݟn�D��#"O�-i��Z����(�kϐi�P�`b"O���uƟ�>OZL�Q��n�.�[q"O�|�#�P@pJ��~�҄��"O�a�MPS���B�G�i��QH�"O�Xje��	r��4CĩI�B����'��	�r�0a�,�7�BS@V3RC�+dO8�r�J �V�.0ië�m�N�<��;����BY�Vw�h�1��ca6"O�@��`I�c���#��@V�U+��$�S�����ƨ����z�Cͳ.�!�V�j���Àܻ6�q2�噰X!�Ǫ"dT�Pf2/��$�ģ�!�dH%`{xu�ԉ8	I�f�çV�!�d^,T�����mSe�A􀛒|q!��=?$ʼ  ��+�$@�� �9l8!�Ӝ<��}`��%�y"@�`F!��P=4��D�2)W2q}\��-
:�!�ܐO� �qeb���Ԝ�wn}�!�Dz[�8�����$�4ك��!u�!�Ğ�E#��I1f�K��<HE�.YT!���F�ܼ���1�):�鞬=L!�dH�⎨�����V��IQ.!���2j�X�3���gq�<�Ch�8�!�O0V�hW.R�0=���G�W�!�ìn�~��_3N.z1��hW�!�D��{ȶ��C�B"+lE��GF�W!�d�\���Q)�$< 
ѧL�cG!�d��@�U�d�t�It�:7!��J;�4!� �,���]5#'��'�S�O3�A���>*ڮ!� �Ŧ,�
4C�'&�=[b�ٴZi���"��ZT��'�"8��xi*��a�{�4�Y���$ψ~zh5�M�uK}S�-�:m!�ZGd�p1��q�|U1�Иh4!�dX!h�Z _( ��*\*O(��"Oxac�X�̍�5ɚ$�)�"OX	b2E�%�d���au,���"OJA�ѪN�mR���mܙ<��4�v"O���!��D>L��Q9y�>Uc�"Obe �W i!xE8JU�b3.I e"O�͋��4�f���!�4p&"O`QB1�M~<���ύO]X��"Od�)`�T�FD�<P4��"OR�R��;za(р�M,����"O�PX�`�.+�$y��H�X4zc"O�a肼��P㣦y��(�0"O��#�ʏc;6�ӆ��tp ���"O��K�RN��I�.AZPZ%"O�(��EۨH	㈵q]Z�S�"O�t*V�T�{��H�6oT�YF��"O�Y���y�  `-�-c�)�"O敉�l�>u>" FA�Ebr�b"O
XSv��Y4��േY�ZZ@5@�
Op7-�U-*�ql��w�1�#�
 7&!�D�x�D��ЪЉ"k8����$�ay��	>���F�N�Z+�+B,�;|F�B�	K#�j�D�%L�4#d�Ϗn�(C��:�H�C��|�0(�AI�C�ɑx��v
M� <06GN�t��B䉢.�,|�Ԁ�M�����(Л`C�I�A��bWgVX4�DR2�H�*�B䉉.R$r�R�3��C3$�(^'�C�I�EҬ�&	y2��5��tC�)� LMdⓒ��R�*2g�ȵRR"O�� �ˍ��"c�ǕmPI�"O��* J�	Y}����)J�,t4��"O�d���	�h�0�`i���!{v"O���C�)C���ڑ(P0a.yit"O�)�FߛR1��G�؃2��y�R"O���G�9_)��"%���#��T�"O�hK�rSPĸ��ܶu��p0�"O�¡C՗o� �Ed�#%�=�"O�l��ѼiD�ɷ"�%f�{�"OڝٓK�v�ּ B�y���ӥ"O q�a��n��ѡ�+U���!"O
UZa��4Lw  �����Q�b�  "O�	3c	Uq������#S�4�Pw"O
�)�dF'vɶ���s=H�q�"O(D�䞌E����*	;
L���"O�Ȩ'�M_"�x5��\��)�"O�=!��m�zQ�f��t�~�K�"O�(�,L�"�t�ґ�+kAQ"O2 �aa	 a�<%Q���5�T4"O"�R��	�U��ua$�#�Nx0�"O>h��$U
�,�h�HE0N�|��"Oڹ�w ǌ=V�us� ��Y�l�Y�"O�P�$ �]�a*��.ԶY�7"O�]��� ̂�Q�Q&#I���'�'W�Ig��/v����+�����i�<a�A�5_˒��*׸e�ޑq�a�]�<�' ��
J�i�T2zL�j��O�<��a%(�0�(��A�$EiR�<�p%�b����H�H����F�<A�� �^����Ȕ9��D}��'��B���E?ĭ3��D9^$|1���'��y���!X���]�=/rL;
�'K����E�J�  ��(j��TY	�'����+��o��p���hh�� 	�'�֠C5ɠ8	��g䇣_��)��'�\U��(�&_�"����֮QB���'�2�+�dգtT��F*טHyJ)��'�b���.Vs���;&�B<9�� k�'\nDU�ْ8� au-�����y�'�TS�g��!���(��a�'�2�2�Y?)��%X �ҹ&����'n��K�̃�HY�4�6�Q�=�
�'C�A3��ҲkFjX����b��'Ɔ�BRnȃPS&����-o(�	�'�ckJ�O8X1�3"9}%�x	�'�ɋ2�U�Z7��1��8wh��I	�'�x�yՎL ^!(�3х��c�L��'�������'>}6a�6`��Z�'p�,�q��W��/P5��		�'�v���Ͳ�,�tǞ0-=�{�'Dy[� ˭��
�)8���'�f���e��~:b�qS͈�}l@�'��8��C	$��E�H+4�,���'��ܸ�M§Ia$5�K�.}�JiP�'g����b6z eOY&��h��'����Ȓ��й���q��'�|0����3:������?-H9�'UrQ��D�$I��9R�-�:>�8���'�hPyPC�L���be]/9Bجi�'̜гU��r�h��b�gd���'O�8 P$õ|��U1!�a���'����C�Q��R�p'ܶF���k�'�ʩ2��ͽ\ƞ��!��9Þ���� ����խ$V~UK#ENXk����"O楁�o��b!Ҽ�f,\��bD"O$���G��[��A� �~Y-{�"O2]�Wb_��0��Y�e��"O�|)�N]�\mЅ�E��OtfP�g"Od8�4 ˼x�~���޼�m"O��˒��g�r��#��./%��Zu"OB��Љ�>8����M a#�!�1"O:�z& �Q�$�2���V�aÕ"O"�Z��E����+� ��²"O�E��/�?)T3��ңXdPyW"O��x)��40��'�0�v"O�z҉��E,	c�N ��L�"O`I�tiU?]�1�A�2}��bT"O|�Z�$T�^�lS6I�#-��!�7"O��� m�. (�	(UZ��;"O2u�d&͡*�HV!n�����A�<�5"�WM*)@��>k��80��~�<�7ڹ&0��S#%��K`�0�T�<Y���=i���F㈷�0�����Q�<i@	!~(ּ�S��{�r ����U�<��O�'"�4��o]��$���a�E�<�Pf�=�X�sgϣ2Jv��W{�<�� 8J<&PSu� $h�l���v�<�1�ǩ%z���©�3W��1Ĥ�H�<A0C�/6w�hR˗t�&�Q��]�<a�'�'!ZU��%T� �I�-SA�<A�x�嫓jC�L�e�|�<"-ős�%ie�̲� 9�P�<�0a��W�E��"�5�ց���q�<��P%F�t��@��68ȋ'��o�<q��<m7�� �/P'* 4���kDn�<���F�m�2䀤Ⅸ"�:T{�LO�<A����|=�E/�!M�y@�B�<�u��8s�±�����h��h�Q��<��E�'Sn�;�H�vrȌ3D��S�<I�I
f�(a!��r��
��X�<�į�܆�p��?jf��"��VV�<���J]��1�IU9���Z�<N�#s��e�U#��6�dձ�S�<IE'�7M.(�l�#4mQ@�Q�<)R�O��*�aT��6fL嫓A�P�<�7��}�~�h�E�'Z3B�Ĥ�K�<)�)�uE���E�#$бД�BD�<y��J8؋v皢=eݲA�G|�<a3@�7��Y��%�$>6-�4f[|�<IS�S�-�v]pǈ��)��d1q�w�<!�dK,��𶊝�|��A�w�<� ��9�HI "�	�a�~��W#�w�<�����=����0X���(���^�<�4e	

[|a
BP�kG�ihgW�<�����?�\`g��P��I� "�U�<�K,S��}� �"�±�7�[N�<AǮ3<$�9(��A�c�4�`��H�<�4�"v�\��BNA�@�K�j�<��,"�(K�L #�|9P`��[�<yt� V���nI�)����KT[�<1�*X�Zv�� ��Sr̳�(�V�<iD�qd&EK��K���YB*�R�<Q� 	�T�z�
"���G�ݳ$(O�<A��F�*)*��4G�kp�{�)^v�<q�.�(`�*T`�&B�f�n�0�Tp�<94#�/�~�YS�VR���
V��W�<a�A=_N��qe�36��X�<� |�P/��$#d�ٸB�~�� "O�}����;��� h��|ev"O,��rՎo�M�dM�����v"O�(����:��"���Q��"O@|���Q�i�*u�q�����A�"O�u1"!7�t������r"O�Xb���Z��d�;OzH���"O��ćݒ:�l�asNI�Lg��r�"O`�h��Ë/nd�&Ǌ�f8��"O��0\	SX�Ha2��1�Z�I�"O�%�'z�@�	*r@�x�"O~��D)��wV`1!p%Nۖ)�D"O��1F4�֩�6Ąp�0�:V"O i��-v)pq�ԟk�Pk�"O��ZE�)�0aє���f�����"O@�Pf��Uƞ�37e+�
��"O�!�� Q�Se,�9Ui��b%�Z�"Oа�,K*h�BeKT�J(q��բW"OV0��9/��m�M�]��"O��h߃LĊ8v�G�x�@h`"O����

t�r���J�Aڙ�S"Oƕ[���20�C&�N+s��Yj�"O�,ѧ�!��m{t�#;�8��$"O,ԁ�i��Q�R���e0���"O��?��e���V(`�X�"O`1i4'��P�dH�`��2Ԙk"O�p�4�]�p��)��c� ?�0��"O��7K#W^����cr�`�&"Onh�0Q5S���@��5ma�Ѥ"Oruq7���wϺ���K#G8.�+t"O�+%�_X$Š&M[�%��R"Ob} �机R��
�L�,�m��"OҰ�A�&*\����K�X�K�"O�] �U
F�1c&lʽ'ƪ1�""O�U�S MMl�A�Kն	��A�"O��K%�;q�AP����s��)�"O`c��47�*�Z��Gxx��"O�x��&��A���8u�G?`�� �"O���d���7d�s��ӜTW�}`"Ov���'�*��ӫ#��,"�"Of��d��H�$�bS�0n��`zW"O�}����2����u&Z�Q�"O4��V��_�H���jֱ|�V�c�"O���I�S�]����^�jP�"Op��2�����QZ�nP�"O
YqbK�׶�p!�y���"Ol�˧�>nq��o��&q��"O�`1R邅�ִ�@m�-A�!��"O5��B(H(�CBl�4xոc"O�mC�	A�,q��+C�J!�"O�]1�a��Uz�\�d' $k�쐁�"O�!�$��RM��FA�?x�Ĥ�"O�)!Ub��F�n���͟�h�	Jp"O-�����*�� Ѡ��cQ����"O�=���Ҡ���UBj�vQ�S"O�9C`V6�,��o�T�z�"O,�#���`�Jd��$�%�h�iu"O.h3C#Q�E*�m(C#_>l�l�Kp"O�����k����2&���"O���A-�H��b,� ��ڀ"O\�f�ݖJa�h�dD<nKv�"ORppǂ����Q�0�6P�"O"}��"�OSVQke�G�f�
�"Oz�ȷ�77�A�v�ήe�*�˴"O� ^�`�H
V^��`��{}���"O��`�̂!xj���
yd�3�"OޡT`�8`�Ryx��UR`Q�"O��Id�E����[�ΐ7dOH�Y�"OJ\[�#��`҅���*3��q�"O�Z�C$ n6��#�N�Tǘ�b�"O8�#�e��SckH�y�.l`T"O�i��Å�x�m@G���� "Oi��҉~�`�[�k��Uu���#"O�\�P.
K^�Y��) cod\�"O4�➼�0)PK�a�m{�"O�|���K7[^u��iI�b�6(�"O������4��l��tج��P"OZ�:0��%�R̓A(D��t�#�"OtHq�$A<e��һK�P�z�"O ��b��55�9E@_�&�T��"O�'¾$�=�QϏ(d"�"Oڈ�"�9NVt�H̭UDే"O�L��)"��؁g �I��H�2"OJ����2����Ƅ�1P���"O4��v�ڋe��q��bw,�BB"Or�ɆcҪWfVq;ՈT�`?h4��"O|�Ӣ�W)R,�E��fT�"�`�"O��0FL�A}p�c2� �y����"O��t��r����8Q��=
!�J2`~m��-ʇg:6�P'�N�Q�!�IM@0D@�/�
	�V��/�!�I3]F�BW֠���r _|�!�D�O�j�KG'@��$�/ھ�!�/&�*HI<�Bd��d�-�!�d�>:v� Jr�ֻej�l��C�B�!�$�)E��#��.h��ȳ� *t�!�W>��3'O�"Z�l�2 h�5Jx!��#�RS�&��I��f��!��kc^�@p���Ph��ͫH�!�,c���!�E�<����$�ǂb�!򤀣D���>s7 �1婙�<�!�$W�Q_zP)�`�6h|�� �JC�!�DگP�
��@�m��"�'n!�dDk|R��1�U1E	$I�t��m!��c����i��i ]����=]!�/B�.��,V%�|�h0/�4V2!��X+2�]
Db��4�:�D_�X,!�Ě�p6�ȀU�ЁC�웳�A�%!�$P��*�����܂��U`��!o!򤎝l��J2/�8M�t��2/�.w!��Y"y��)��!ğ"������-b!��_9���I�\+
�bB�Е7g!�$��E(��SP`"u����0Q!��Ǥz�@�AY3"���00��P�!�$�9�>�Di�Xj�i����0N�!�$�48���D�F
_�q���;O�!�D�=9Vȉą�c�:I��e�N!���)z��l�ẃ#P�� ��,�!�$ս
��|S�^�~�&�X�˟+�!�$�� 8@�G�5�$T�k�]!�$���l���'�@�򤚈:�!�$�
������8N`� �؆�!�d[%F��d ���dL��{�!�5[-!� U��{�d�?91�3˘+u!���<��p����$�h�F�ĩB!��}N��B�-1XH�i�K�!�D՞{�Ds�̓��
�Y����3�!�Dǡl�)����2+��r7d�?u�!�� ZqR�M�q,���t���$"OFab��V�v���1�FT��"O\12�*W��Q��@\�^�w"O0�:`,8q5>m�p�$oi�h�"O>�c�9N8�%kE�9a�ӓ"OΘX�q�}#e��6H9��C&"O��#��G�a�6Y�4-�)&5�ŠU"O��*t�	�
�0�H#��a��L��"Ol��m<�����̅	��$�s*_��yn��X]\̀�CR�{��0dB1�y��$[i"@p�]$��VmE�yr*� �Jt;�ES''B<�6�F�yr.�>�p0��mK!]�8��dK�y�m�������$��u�r+	%�y�]J�F� �����ؒCЃ�y�ɘ9!�!1 �0�f�A�o���y�f4�@���דn (I R�U>�y2�ıe��2��I�f�d0�p�,�y��
�Sa�	K�nG�t�@�Ӈ�=�y""T �,3�C9{��0�.�"�y�h[1N�L��� ��4+�����y2�>" #���]O��j�'9�y
)=p���"�X���p����y2IL55�,��/�R�� *@��yb��$:���	G�I��5��܅ȓjZ`�WK�%_�Е�_6
��ȓh���f�@�ǔ2Rtԇȓ8�R�'nB�[���Z�Q�+x�)�ȓN+K�'K�eq�Y¤�0T1�ȓ&�u�D8�aن���2�d���2�H������@F�cVfՌ3q��ȓu��+P�P2���d;88�ȓ]�Xd�7ř.Pn�г#��3��,�ȓA��a�����ܙ"!�H��ȓ$ME�!D�^ڤ�A�bR���x%&��a쟄�ް�O>�2�ȓ1�d�2)8Ҁ&4����d�����;XP��2�E�(�fA�ȓ;�$3���G`p:f�T�`؄ȓN�x��ENEҼ��ӕ|� ��O��Y�e���|�x1�aL�Ha(���N���F��=�h�G��9�xu�ȓt�|�hW�D9bA�!)ʹ]�:�ȓ0'�0�.�=K�T�D�@�I�`p��nXȸ��![w'xQce!B	M����B �ܱ@�Ls�����Յ�O��<�ǎ({��(� 	�2���ȓKVҭ���y).m��?�����:�m�AQ�Bɬ8"Q 	�e��\4��A�.�T��&&�2��ȓ;��C��2� 䓖.�9}����ȓA]*�ɒ�  �����@�5$�ͅ�R�,��W S�$��x��F�o $��%h$��OZ)��1C"&� ���ȓoK̕[�T"%�<�����
���~WT�it!̓n����b��oɾ4��aP<����^
9)�tZ�U�D�Ƒ�ȓ e���we����	�vj��	J
���l�Z�����~��P�Х�u����D��	��G�D����@)2*�V����n�Vg�%Fy�1	n�<P���x��A�f\`�,XC]�u.�Ćȓ5��9Ѧ!m>e�DE���ȓR䶕�s+�2a*�Q�q�W���S�? ���c	� ��#���q4"O��¶�J%��ja�é,\�T�
�'e����iZG1��E!nl3	�'���7�S<q�������!Њы�'z���q�Ŗ~|:2L*Kg�8�'5�5�%�C-6]j�Za呲>���0�'Y֡���3:�a�c �*�a��'���r�R�(A��!��ˤ(�X)�	�'ʹ U�S�Z
^R��2`Q	�'�D�8�i��#�,�9��ڦl��K�'�Db�63�j)i�Ȓh��%p�'/t�ӷ�*�B!�v� c�'��t���V�$d���ҿ?8�%	�'V���0(A�mD2aR�EI�m����'�M؀�]�7��p�l_Q]4��'��$E��k��D*I�R�'�P�@���> ��� �H�x�:}��'�je�S#��g)���t�������'X�snToaT%�fQ	76dY�'��d)K�T0����Z�t9�'�p����N;661+�!�$="�{�',Xp��9�0i� @՚��P �'yFP�-�Omz�P�]"uW�4��'��R!�$ EҶ@��i#x���'@��!�̀9T�yQ#\\r=�'H@��ȟ<�,�Q���k��m��'����� Ӟh��,�f�3nT�H��'�$34-�e��D
Q�bx
�h�'�z�q4��6�>��j�$cC�� �'(�5p�%�*^�x9	��(V�0�)�'���{U�t�jM[�` �%��e�<a�z��Y�v�3L"�c� W�<'$��?Y:�Q�㖚�@6Q\�<!1B�b*�G��o,~�+u\�<Y��,�������j�{�ƆO�<���X��@��	��L�dR�<�q��?OxZՐ�%Br��sCR�<yu
�m��x�h=KaS�m�L�<!S+���\� /�Q��aBl�L�<1G��k�b���GZ�{r��t�LE�<)p������;K���Z�A�@�<���6� p2a�Z�,tĉ2lXd�<yC���+e��a��ҭgĐ��7�N`�<a���.�d��& V?4�x�i�B^[�<ن��F
���ꌔ6΄�ѳ��B�<����d/t��6�z5�aQ��s�<9�!H��|B�錰 �v���h�k�<�R�د|Ҫ���IE�J֪%�Bc�n�<yE$ӡ=�􉑂�χC�E��kCC�<���V�C��!�q%�D�$���I�<��
��� ��Q7��ISj�<ygڀ_lB�za߉^(�����q�<�
\#<����3��{%��
�N�g�<၇3S��C!&p�:�Hc�<�AN��m�-B�hY?P0��hB@�U�<9�+U1�|���Wd�&��w�<�dX��.K ٹ!|^�[�n�r�<��DX\��떄�2w(��۴��n�<��F�Nu�P�ĦͭA٦���Ov�<��-�\PɆυ%=M�ebc�Y�<��ٛ],�3AM��X<p:r	VK�<��.J9���@ā,��Y���J�<!�� �&l��N�-��Yq��o�<E�Y�UI�L!1�&_X����l�<� 2��"ŗ_�v@[.�h*t�4"O̤���c8T��GO˿R���"O$���J�0oofq�A/C�^hr<�C"O�0���	'v�Q(��yUn��"O2-�!�0[\=��V�2�*8�"O*�K��\�G�^i��=���4"OT�1�GV(k�(�ǣ��?�V �"Opl��;6z`+��ژ:���j�"O�pI@�(�ש+]�N���"OtL��n�[=�q��'вA�e��"OFAQ���]F���SE^��9`"O���()rV=y�b�>@� �$"O�U(S��a�tD*!��q\M�T"O~��&�ͦxA�-�Ut)X�"Od��7�S�E�@њ���K9h�%�d����ڸ2 ��S�ˤr��E� -�+C8!�֗90�0b@�ȘJ�b���.J.X1!�d�qo|��=6���%g
;!��:7+ �2�+%w���f��^�!�Ȅ_O��e�:�ԫp%P�c�!�D�2,��pz@"ӛ%zb��[�Ko!�d8nVIr[:I�@-��HN�Ad!���&<�r	�GOЈ)����E2dM!��c�N4jr�O&P�[fdդSL!��#DD�� �I���a�@,�!�$��g���LA
h�]��2�!���7 ֦��eD�(%��Yւ��!��_�V�2��'g�f� S�ZT�!�Bmxp�(1d�Gp�=ze�H��!��<o�����-~�앹�/�i�!�d�`Ǧ �r�S�tP����30!���<���v��������?o�!�=.K�ly�l 4@��*Am\m�!�$�����E+jD���>g�`��'�As�'�l�-QVK�*	$TA�'��,Р(�3'$8��Ô�9�OH�=E����<V�2�a6E�)l�Z�# $�;�y�N�:�\�˱(A<`],��恚�y���V7��FCY�Sd�"�G&�y� yz���C�6]pũ�hɆ���@yS�H������hˢ��&IR,{�h��P�hurs&
�L����~y�<��%W {�<���Y6)�v��<���?-O��O󩇶P���V�V]�`ڳ�V;NL!�$T2`��ٲ��4LM�x�2�ПbG!� /.f0M��Q6k�u�êJF>!�Ć$&
�F\�sX���Iͻ&I!��X;5a2$@,%=X�0&��a�!��7��0;��
i'�%����!�� ����G��}�l�"�	�L���l��hO4ј")�(7�f9�%B��i��Y�!"OJy�e�*~���A{x��"O�y�cɋ�\*����LYy��+�"O2��`E
�c�bx�S;pt�e��"O`�j��:R�ɀMY��F��T"On-Y�J�5(�	SS��	|��!�e"OL{�ŕ���l�Jˋ
ʄ����<).OJ�?�8������ȕ	��ԙ1�.D�d9%��Х���Ǽ6J�-Qt
,D����f҇�L�1X���9d�5D�t��$%-̀�1���1�d�Jp�/D����nQ�T��yz��Ǒ
*m��� D�xb�D.Ͱ@���W� R
m�>D�,p�ߔ�F�çFV,(�	q�z�ؔ'�ɧ��� &�w�s]�=ɖ�E<Gjq�"O���@���x��cd��V走�"O�a�BJ��L��X�&@'�����'-�0$��A3�9�B~ɣ�'��|�5�;2j�H�b$�3sQ���'|��A�Fm4Z����o��C�'�6Dd�Y
';z����z6��i�'�����:k:	f́�vx���'�h���)�/@��D��D�0!��'0B�A#��K���s޽::���'�ʩˇH�f#ĽQc疎)��m��'~��k��`�d��cǗ&���J�':�0"���:d�ݱC�7��I
�'yv��s��(�������>�	�'�"p��.4V��0
S�T�bܪ��:D���e���!�D-K�$A6<�`k+D��I�`ݛ5�Hq�P�ѿ;�$�: �(D��0Wj�I� �aQ�\�43�G!D��sfj� }8@�b��M�d������*D��@K�Oz ��F�Ioޡ�j'D��@��E��3�ˊ]�H�k:D����9j�P !C�w�p� ��3D�,"%�q��@��H�>]|� �j5D��s�AP�c���h�)ȍ"���9D��BE�E�����!0q���S�6D�l1��Ȇf?퉖�B)�~M	3f9D�$��#�N�J
ޜZz�b�7D�t�U��`0�U+.x�d}�ǅ6D���"�V
���k�ꖏq�h@pP�2D���������ժ�\b� ��1D�p�B��?#�J\(t hX���/D�����8jJ��`�T:�(���:D�8Sr$�3�&��nBUY�5D���f��C���83K<Uu����3D�t�d�E<��a�D�WeJ�1D����Ė�=�^�IRHA�2CLܳ�k$D��b�X�f>5���*(Q�?D��a'Á;?��٫C�=}D �F;D�(yCK�h�zA�]�Tц�9D�� ��̲o8i��	 1��Y�8D�h��eƹ9��yrB�>���:�/ D��5)�ۂ�9�hr |���<D�������21��&��^jTU��*O�$+�*�&G�b�1�K	�n+����"OJ�Z$�aI�u	�Zp�is��,�y��(|5�\;w&_�Yj��Rؾ�y�`��J��`�b��1M˨H�2��?�y�Z���X9�
�5�y�tj�y"�X�� ��8&���Y�"H��y�FX�f�� +��[R�J�$K-�y��{�6Q�D�<4H�"�S��y��>	�N�[�Z1��h���y"&G�o4\�'��'�x�K���yB)��y՚���gϯ��@3��Z��y�)H<e��=����:"R|Q����y"�C')��1��W�	��S#O&��$9�S�O�@Q�t�[�P����EA�,ܠ	��'�8���* �'�V���)�#sS�@��'A`�EТ{nR�z`kF�^?*I�	�'l� &dL gFpC��ERZ&T��'謄�$A&$"���j���0	�'j���w��,	^mh�(� ^���j�'#���U�І`�����ݬUnT��y��'^�O1��yp��ƲP��i���E8Bt��"O� r-��L�5�j���Ձ
+���"O� �5��,���^$r�ѳ�"O��IpJ=:c���R�Su��p"O�C�\(`(��H�ꕜH���R4"O�t3��Љ�8$��
^�;�Xt��"Ot�����1���Ө؈1�Ie�O�̰�F�� ۨ��԰ID��' �Eӧa�q�L���� �H�L���'����#�(�x�a0���W>�U�'Q҄c���2�����=�<��'�P5�a�n4t����-0�lq��'�j)0@���C4�MB,I-t9R���'��;��0w��l@���	�� ���D6�S�dE�@9"�:�CXbX�4���yR���N)Q���� ?G�U��G-�y���3&�JEj H��!1�AR'FI�y�mD)o�n�`���k����JL��y�\%`�(a��/c�� ����y��(*8�����_)Z*��:�.���y��Æ4^,H�oM�d���'kT�y�m�ieƤ�d@>0�Q
���y���a6¡р���%�$d+f蕑�y�e£X�bD9e��S�d�� .�y���2h ���W�� [.\�z�b�:�y�)�%> v<�)K�MY�Y ��y���@�HU�ҥwƽ��٬�y©�/�|ehԬZ�$��� �yҠA��FE9�!(X�Z oS+�y��R�eH"KB�u�|1+��.�y�o�*IRԢ'N�u�������yL,
��d�2XrQj&��y��O8`=,d�D�?�X�8� ���y��G ��� -	״ AE���yr�@�|�,��`��|5����y���^1�%�h�lj�	2��yc��e��R@䏭qZ<�4bM�yB��,25 D�����!S�î�yr��9Q)��	$���rȕY�0�y⃒�0Rl���� ��p��:�y��M=z5c6���pK�H�KO��y��>t_N1󣏐�k"LBT6'ў"~ΓSrx��e'X�r��!�O�_�Jl�ȓX0�����̶K=�<�$��ARԇ�Ak��A�)��fI,�"�PL$<��'V�ٲD�N�EXF5�W�Q�.(u��.Wd���!Ɯqf䱧癇]��ɇȓ��k��O�'t�YP��V�?7F���Uج;��O�*��H S.ȽXwƬ��J��I�l_/q��T���4wjVŅȓ4D|�c��e;��K�/t�4�ȓ��I�(nr���4L̋{�$���"OX FG��fP�����!�B h�"Ob9��SHV@*�DGl�  "O
A���Z���RD77R��X`"O��c�W�l���䄼��x"O>!	F��'p��IH�#��]��B"O�D l��/P����+�̍��"OT�+Y�\~���G�w�;2"O�9Ã
����ҒG�5s��8"O�m
�,�N�@�d  ��l�"O����E'��]��K$U�:Hz0"O��)�+��+j|2NM�b�T��"Or����875p�_�{��%)1"O�R"*P
U�D�&V30�$��a"O� ��D�šEB���d@��$� �������O�t��f�]�v�$̑b�>~C�I�9�����k�
\�=H"a�<�^C��(F��L!#'�Q�y��^T��C�I! "�A�%q�\8�̖:=`���$�<���Rx�6QY�H� �����w�<�QMK_�	�������Cov�<�Z�k׊��͌�#ڰY�\k�<y�ƀ3gXE�oJ rm�(��j�<i��Flq���OIw�6,h��[h�<��Bɥ)$�A�¡
�oAm���a�<��-.������)��
�ʏf�<q)I)r���V띹(}��^��?��Nb�CdĜ��n�2f�Ƚy�z��.#t4hs��"�(���(�:b;ƅ��/�Y ��GH<��Y=����ȓ2O��t�z�T�@u�9{�f��q��aH�?������7.
Dͅ�K� 5��N��ȼ�7��4Oh<�ȓ r�;��i�d���N�o��Exr�'V�[D��rf�h��o��/Ü���O���D�bQ�QR�N� ���O]K!�D��Vp��x���wO]�%>!�$�9W"`"��rL��8I�!�d�rHC�DC��!�-��^�!�ƪ\�Й�+�>HȘ-�R�C�1�!�Dβ���F�V�RqyV�F�E����	=o�-���_� �:�b�5c�2C�	|H�� �,H���&i�T,C�	�[֮T8#�Y:����'��+C�	�H���Ǣ�7=�а��}&C��/AvI�b&�1a�h���:�&B�	1)����'C�b�0�HG$%��C�I�bzpk����x%�3��
 +�C�ɫA�.�B�-JЮB2��<#��C�	� h����A�>ONpH��E}�B䉢�^�2��U�������#!�B�ID�������@ u�d�x��"O��+��97��*��߇tF$8"ON�22!��zҌ�!�͊t@�h�"Ol݊ gQ�/{r���.9^(B�@�"OThAb�L����G��,��@�"O��K��i�
�tF�\\*�BE"O��v#=P�h;�eI�*ܼI�"O�X�"�F0(m雷�E�/ޅsV"O�*s���
{�4	#'�2Y��m��"O������'�"��dc݉t�D����XG{��	�%Cb��.��3x��o�!�%9f^��*̙~��Y�+��@b!�Y����g�
�J��drek�//!�D04�;#��
y䡁���.|!���C�j����[�Rr�(�d��!\!�d\3O��@�`*�Sm�w/B!�Α�}ӱ&/-R��Z��O�bBa~2U���C#��7���BW*�]�h� ��&D�d�g�,2܁P �X=h]m8�j1D�(�6�D4K�Z`��!�o�
U��.D��`���&O�����J�c���07*,D������ �X��Î	�WG�,�%D�d{�/I��q��� ͓g�!D��k MU9��a	�C
Au��)"D��
U�;=�v����BSk�L��  D��Bb���f1T\���:�t�hg�!D�0ܩ[���� mO����d�9D�� Xҧ�	� ��&�,��"Oz!1��-����*4s�va"�"O&��w��-bh�JV���1�%"O����у�	J�N�*�y�����	N�S�O��d*��'�y!��D�8*���$<O(�W�p"TH�5��Uɠi����O�b>u UJؤ<	~0�2*�5Z�h��=D������ !"�Ӟ8Z�A�@I>D�p�u�/&�uP�#�3&�A��(D�л"�R�zs�o�|��*:D��K$��$=H�aBȹA>�P	3D�����*�y`!��� ���#�1D��	ȓzE�+�O�x�����,���+�!V�l52���go��iDR�<Y�c������_�<�-�ǧ�N�<!m��A�h� P� c$H�f�GL�<5��x��C_6�x㕾�B䉡x�������S3�\�aO�:$�����>q!�0a�� EM�"Y���q�HT�<y��\0`jC$���\�*��N��G{2bB=&�T�!�*�;Y)ĀJ��y��6Q0�8 �HS`��Q0��6�y�˻~��U�\	K�V��e�=�y��J�E�L-!V�F@�=����yrL�-,�4-�g�1.uR��Pᚋ���8�O�Y��_�Sq D���D1mR�b�"O �ţ�>kR�{��ҿ.�>�����)�'J��+���;�>}�t��5y,<��ȓ6s�����A�wY�	��0=���ȓv_.���� �r�U5nB"X�ȓmy���a��z�����;@G�)�ȓV���Q����24s��Н|����'�'��IpS�
�}������Z�4tT��'��t���%[<��#Ń�"1��'H(;�G�gRm&��ʤq�'������sxCt�S�u����'�&Ȫ�,F�@�P�!t�Ђh���
�'�����YS�H�x����]�"8q
�'�X�F��K��x�,�/$!nic
�'�%�3��9Qc���� (�,h0�'���Ď����	q�f�I�'�@H��F:D����u�Ul4HR�'b�4��B��{:޹r�Cw�$)�'Z����� R��ɹ�U�q��tH
�'�P\��O�G1�qaˣf���3	�'Qj]r��\$� � n�Y�$`�'�̉�%iF4�	� d�(?��ـ�'�%9�F>��!s[I����b�,���	�]%v�s+�|zr�����/�l��x��,)$Ĕ�Wm��0Pd�04�W�=D��eg��Rq~t�T@��~� �#�n D�\�!@�9�䓒\ŲT��=D�`3��6
.�3vCİTk����*O���`�-"�P]� �\�H��16"Ob�IfN�2dn��"2��4mPL�"OZ�����};qҮ�!Dh��ڦ"O����Ƿcs�����I�(��"O��%��zo�
��%XM��"O�}�C,F�D
�|R�Nۦ9�<�U"O�K�YE:�D
�I�$n�;�"O��(��6�24�+��<�:�:4� �f��"�X�h$3URL�F/D� �2���X��K<,� L,D��i�Bu�6uE�L�B:<��Ճ6D�� �9�WէQv8���֪S�\@�"ODU��<������x^��w"O��z2�߿;�sÂ�U�*y��"O~���%-�=bW�\
Z����"O���憅D���1��$o��a��"O�H��kè)�<�:RDئd,���"OH	� ���(`�"�9hQ���"O����ܸw~~尷�[�/� �"O�k�C{�nhp��j>}K�"O`-a��<\�Ȥ�i�/b±�t"OԡS�8>o$Ї�Ɨ2���%"Ox��Ĉ�3l&�uX�IG��x9�"O��R���N��h�cCj�h؂q"O��C,�2
D���!��W5d���"OH�F��Y���(�oD S���"O��QsM�7�����Oͩn��20"O���j�7���p/�\
��#�"O8��*=<d5�D�'"O$�3q�J4Xy��'�u݄б�"OH`(F͜�X��q+��[���9S�"OP���"��H4��CRĔk"O<�q��#�L�Ↄ�<��I""OVm+�eC8D�l	� �[nT<��"O�aRG`Ѓ�X�Q� ڇ[|E��"Oڬ�GI�68�Y� ���>1�r"O��#��$�$EB�˼6�f�q�"O���%@,��a�4ϗ�,��-�&"Or�9�J�H?�`vM�*��I��"O~͘B��xI�@�T��]x$�`1"O�m��KZ	BB0J��X�>Y�"O|]�F��coh�;@+�x���"O}�D�q>�a��SM|�yp"O���AB��#�  aB�ĶD�M��"OD��e�7=����=#+x#�"OtA7�]*A"��;����pHb "On�;@Lƍ@M����ǁ:��D"Oz1[��J�����y�d4 "O�衳�K7pT��vď�H��x� "OP��Γf�^,�����=v�(��"O<��	t�� F$N34�,�"O^xC@��F�h�G�:D����"Odq�b�N�XA%��x� 
�"OPD[SgM�7o��:V"@�z�\1"ON�:�Z"H���-$a0�"O���H\rCfk��	1c���"O�2�,N^��(�C�*!T��5"Obk�J��@e�X� ��O���"O����R�!�Dз ����"OY��/D)����5fôw_�ay&"O �k�M��E.�[�kP�a#��"O@p��@�(+c2���2�8u"O�|	��H�C��h1��A8�!&"OP|R���b?j!�c)���)�"O��TO��E՜�k>0\��e"O��2�M��'�F,ZP��H��""O��C��P���H;j(��@"O`p��C2c�h+P$R�re�HG"OZK�	Z"�tm��[1T�g"OV�;���4��FҼS���p"Oȝ2���]m��.K>ex
�� "O�Ya��r�ؤXW 1WYb��`"O����v��I��� o=N�"O���p��P	$��+��Xbds�"O��+� ���	  Iîo��9�"O� LA�B�՘7�=#�b��=���w"O�}Ө�V���?����""Ox��h�B_N��"D<����"O�]�®/�����@V4	���3"O�)�Ä���`�3OK�1��IIs"O^����,Q��X �&�����"ỎB��(!�DD���-a���w"On�1�#�&�n4��앦e�T	Z "O��b�
V:� �
��x�ER"OhA�䀕�s���󉖝5q�8h�"O�l
�a:!�B8G�CW�X��"OD��DB'4FQ�3�?3L&A7"O��3��a*P�RAO	Uixt�a"O��B��Hr�!�K�G� p5"O�9�VHR�ElH���g\!?*cB"O�- ��S��:��<D���W"O�p��νBO$�*��-I$�i��"O���Z�����$�U� R�
�"OBqÍ�U������ͲJ>L��"OB)ؐK�Y������0�H��"O"�K���#D�9B�	O�$��Y@e"O'G�#���R�)��	���"O�5�7�S�^%^�����|�VX�"O�����޷7��!��B�/�pˣ"O����͊-f؆��r�X��xR"O�<X���0w�^�HFA��5�V8`�"On���C '�llsd�X<w�R�c�"O*��E�	M�A�g�Y��Y�V"O.,bX�	j�Ay E;n����"O�UɒAַ�$����5^H���"O��B��J5�tIR��-����&"Od�$���y���A�o΋Zp�s�"O1J����,)�=i�hL� j�v"Oȱ��B�R�nQ��%H�y�"�K�"OJ��Wn�`��Hcu�ьJ;~�"�"O�(�5��`�a��EJ Y7JU��"O�u��JE�C�b�I`D�![@��a"O����ݑ�`耂c�'q2�0 �"OL�s�/�78\K4#H$'�(y�"O���,�s�*�C#�#$��d"O��B��2\sx���"��o8b��%"OZ|���P�R+�H�u�)p)��+�"O��v�A�
4�Ua?=�#p"O����E��#�D���#>��f"O��TE9(N��(u�d�&���"O⍡j4hWt9�ψ�S���F"O�`p I�o��u��`U *�4]r�"O$ y1_�C�ļH4�<W��щ"O��2�	�7��1Qv�Шj��A4"O���`]�9�Q���.��i{�"O���)��o�g�;�AC�"O��XӨ��p[̍�tj2��qA"O�i%�����H
�*<�`=Q�"O��#��k����Vψ/$���F"O(����^�:��!P��lԅ��"OJ����*0E�`�'�RE��"O��* ���)�U�|���r�Ǔ�y��}��9��Εy�Re �n���y��G4�P���A�����A��y�Z�P� \X�X��@T�A,��yr
Φ3�̬x¦�24�2��y�fF�F� I	�#������?�yb	L>"���t�ښx[�lZ�ù�y�ك-dl�iqʝ�v>�Ă��*�y
� 8a�'�["3`��V9ny�X�w"O�Q��*ɿ
��)�W,��?c�H:�"O҉���Ž#  x��9`S��#"O ����	�',�ʕ�:eP�Yj�"O��Ӓ�͆X�F-��N7c��`e"O���2)��N�$�� 
�<��4"O@���O1k��%�
��:1"O�����W$H՘��Øq���"O��!����e�țя��(ڜ�C�"O�����!��E�c���n\�"O6h�cO\�"婗d�%a����"O�R-(3	�8�WD�#7;n`�"O�
�V,.�I�#�#�yE"Ot��e8gg�`���u	H!��"O@Xgf���lk���p�$"O�Y�a�hl��h�I�l"�b�"O������*@���UF�'�q�"OX���E�?
��8�& �J����"O������)�L<�RA���`"O�X�3d�/n:Ce�2w�rQ�"O���l�7��}��[�p]���yP΢ٲ��a���aю�"3!�ą�|pq!w��t
�r5�g!�č4u!��E�UWp�U��Q!�$[�!Q�$�էX�J��}���� H>!��T�|Ԕh:��Ռ?���$̆`�!��-:��2q�����h���w!��*3���Rϋ�~\0P��oߟ_�!��
�ה�@bN��^�cfn��`!�d�	�Ju���M��� �΂M�!�Ċ��������"~��Y�'�v!�,�0��a'ڎ2Ĥ�� 
	x�!�Ċ<8��-�G$�*?Ô�h���vo!��r ۃ�)D���g�J�JP!�$�0:z�ҧe���	�����s^!�d�6v2|���
3j��p��7n!�d]q�MF�\��0`�
ߵe�!��O-0�!�&��C�΄>
!�DȒd�:�����38$�����!��� pq�0�B;.�<�A�C�N�!�؞-I&���%N>�)���J!�dդz�ĭ�QB ?T������.!�׷���q��'y��̈��F�;!�d��-��y�GI�-��u�T�U%!�D��fDXhE��Zg����O��o!�$� �ұ��l��&��4��M��x�!�D��Y6����k$�,L���8rV!�׉A����w����*	¬W�!�Ĕ+j{0��IG?)i�L A�+Y|!�$�^(����RQ�=��#$l�!���Q& �)4]�;7 ш2��h!�D˛?NH���&M 7��P @�(.�!��$v&A��NF�uX����N4w�!�dXER���ʢ^|c�.ĸ�!�D�:F͘D��[;"�:q�m�7*!�$ٻi�@)�7l�<C�Td)S�	�n$!�!>�J �'&�:��U	Co!��Ϭ����rqQ��b��%x!�F�H�F�B�M�
�ʢ�Mf!�O�d�4�C!D� �t���:2!��|�"�xtj�=
$-҆�-�!��˚|0�-��{x� i����Νu�<���eNvE��ˌ'?��E����Y�<ɡ�Z7&��a�G&OQ4�1��R�<� <$�s]��1����
~ZŻ�"O$�4�_�t�rGL�YP�X�"O\U1�¥]}�҃�_�2���Ze"O��Wh��X��"�?�Bp�"O�l�g��>w��5�6��[��L "O�j��#p&���o�r��Yr"O>UK ��$G> Bn�sSzX��"O^u�1�M�c�`��F푹I@��"O�q��K;IZ�)�`�(B2��q"O�,j��g�v)�0��Oxـ�"O�y�����M	��Sc#8��h3D�H�4��e"�3�&S'��K��$D��1EL�*c��26�,J��c#��H���"@���0g�H�Y�|�X���6x��B�v��XB�� m]~	�B\nG�B�I�0�.U*�M�!JՊ�	�٥}�`B䉔^.����`T0d����7V6�^B�	�:�T�祎%y��HR"@�@O�C�	"_4y0,����vi�`�C�I��\���W�}`Ѓ �4g��=��D���BE���K�� ��l^�I�I�ȓh4,"ī�xK���B@�#���������R�L�>���z ���\@�Ie��F���iΙ"�ͽ*��q���%�����W̓p'"4��)0t�l=�e�FT0��w�j�s�L�Z�
��Tj���O�8k%��{�S�'_���+�F��I<�
S�/�F��ȓO:Hu��� Y��y�!)��w(ۉ��s�T�f���x5��j��{����6��\���'Al(��َQ0���-J�QA�%��X�$T�3̒*L��\]��Dz��'&�՚aY=��<*'�N�Uf� �	�'P�0��e�Y�4X!ʄ9=��p	�'� �#
��k��0�ɺ3Ц��'z��ΛtV�k��%�ȭ�'��E�G��%Gܠpw�/.�"`{�'o�P/U>���P�eɢ<����'[>x�B'գ0N��E�[r�#�' ���UB��|�Dk��j���yҫH/n���@� }H�uxVG�y��Y�m���NS p_~��%�y�B��o����-�^r���0�T(�yF�(!�"\p'ͩ$��4���E�<�!�_b[VZbJ�
(m��q�Hj�<�g�j3�iVjƛ%�4���jRP(<�4}Q�t�7L;1���c�:	�p�%(�(��cG/CE� ���±-E|�{r�5⓴y"�H,��O(�L��B�Rb&�xe	L���Z�'h4�����&�´�t�0D9�'���H�)�b����K�"I`#j�Hl8��J�h�1p��.9� F@�*"=�O�8��	�	��H[�ٌ`��U@�I^3b������B�LˇH|��)���8u��d�O�C�ɼm�9���٘b�i��(�1"�C�ɨ2효���G�AP�K+6iLC�	'
�X�a#�4�taA�^��B�ɕ^:���'��nx�'A܉�C�I�sk��uៃ=��{W�\r��X�'��EcV��4T�a�N>v��'a��Y�&P�M%�UI�O���	�'P  ��f@f3���d�0�A��O �=E�T�� ��-�G�ۣ=���)��y2a0%����폳1����$ɍ��'^a{
� �٢�f=�":P�@62���[f"O����B��'W��!�� 伥��"ON4�T*W'X-h�H,i&���u"O��4#Џ'���5�b��"O��`!�PQ�
$���[�P��'����R7EZ	O�b}�@@?|z&tu�,D��p&�t,�q��8|�<�u#0�D�;��=��5T��q9���J����-C`x�� �O"����O�l�%�6f�i� ��(w�d�H؞�	%"��S&�|x�_e^yx�8��(O���-~��-��c�4Œ�cY�#�!�D"va\�tBϜ	�&�6BI�J�xB��h�'���I�Oj���b��I�Mc�'Λ�͜=��ɀGB�J�t[vOë�䓈hOq�&dk5�����q'@-v߬hR"O�@��L	!61A&aJ�<��+'�D;\On ����\�d$�"�J0A�:��"O����/�o��a	��:\u��NH<鰊+S���P�K67�Ʊ��(�i�<y�QoU�L���K+�#Ղ�i�<��ŉ�o_@����S�X�Lc˔f�<y���L�^hÞetb0C��i�<g���o�jٓ%d�XZ0��-Jh�<�G�ʈ�a�v�Ɏ@��aIpG�d�<��� �ڰ_%��K"�y�Ѹ`YzPx��K�X�
]:�*�yg�)��l@�˭IMLY�A�F��y-p�ؕS5b��Pޔqn	�yr9|\p�#j�?JF���@���y�anX���6��Ĩ�M�*�y2AGF���R��3�8�Pw͜!�yb�޷Z � ��.:<�˖��y�䌴4Ʊ`�߱[���#6'�y����-��'��M@��1 ��y�K���$����Q��$�f
��y2�V�DQ�7�E�v"� �&��y�nK2�$X��_=Dn����9�y�IX}hD�饅O,+$�=����y�`N��H@�v�W���3��?�yn�QrM���&g����	�y"�D�Z�R	�S�U1+ e8@J��yb)��"Y�Rǈ��H�{'���y2�,2x}s��&&d1z�'��yr��7at u*'_5�� �k	7�y�H{�M���?O�Z)f�e�(C�əb���1�*	;��Ԫ  ��m�.B��`{R|�E�(���k���-}@JB�I�u8Mc�,ҞG=�1�C��(�B�ɂ?-��S2G1vA�ui�1��B�	�z�ji��gC�"T$U;�	T�B��y�ʁ1�웰s���@oZ;^;$B�I,u���32��&q���Ї�J��C�
w�������_��-$�E�֤;D��8tϗ6�}���K�p:w5D����1tl ��%�nٰ�F5D�PPCJ��':nd�1�R/�� XA*4D�<ӷ�I��
 :��ҝwM��dn2D�HтF�<4�t���I�+D��В�L�I�X �0)�?�H�")D��j�*�.TO�IK'I]�KXĩ�!�&D�(Y�#�6\��BGJ+u���`-#D�����L��j��{|~YQ�h5D�(�1�	��qI�u0��[�!��P�@q
�O�:I�c�h8w�!�� `YBPΊ�t�����[��kr"Od5�s+ߨc��c�L]�x<�D"O�Y@G�C��ĠK�,��P��} "ONQ�I\�thP"I�S���
"O�8�u��<|U�e[�d�ʱKT"Oڕ�ATdW\�+cЫ/	�8Q$"O�y�G጗^�v,#"F��M�
���"O�:�b�v��g&�?Z�u"O���$fE�"a�H��%Ύ�J���"OVQQA��E�$@3�O� J�\�"r"O�8�f��2U���$-7��tR"OI
��  s4 [��¡4�00jw"Oܱ����))�6�RA��;|f�@�"O	b�j���� *]�"O�Q#2eQ���8��J&o=V��f"O�ɵ@˰=��� �I���� �"O������U
�p��I{H��#"O24� @ٗ0.L� �C1v�MsC"Oԩ���P�h�p c	h[l��"O�T�1A�Yz��*�À�=��Q�$"O�pa�2T�JYYC��V��a"O���!R�']�pY�A�%t���`d"O�P�$���r�C�4LL�g�<QS'�=8{�= Vʐ� P�Q�u�M�<QU�}��4@�L!���ׂ�T�<y�#�lMɥ&��!IDp�S!JW�<yWO��`��Aէ
$���$�VS�<�Qi�4l�p�mP?�!Ka�VT�<��0(�@�"V&8@F�yzC	YP�<A�釭F��I��׳~���˓t�<!d�͚k�Ι�6��n��T�Y�<��큦}t1`��ەXdޭ╮IT�<��!�.����S�|����P�<�P��_D�mz���G,|�����M�<q���XGn�k���aZ��i�$�K�</��B�*P����H�0�ZM�<Y�ku��1�5d�)++|��.�I�<�fb�3��<XPAU:W.��6&�o�<��`�t"�CS$����d�<a��x�&�5��">�F,��)b�<�f�1�Pu��I�"|X1���Z�<vk�-���p��vU����Y�<q�ꆰ��XA��3��A��FAW�<񰎋�=��%	���.��)���W�<	cNB\8Z\���=6ƪ 3D�w�<�BC�)6�����CL�QXse!�s�<�@��K��)vD�|B��ZF�<q�.��EK*l�ɒ��I����~�<q�1� ��RoG?��qP�}�<��ʜ�O�b(�Ѐ�4wy����*N�<��LQ.Ny�&�G�/�&���CO�<Q0a�$r@,��d/�mٸ����^A�<���i׎��!b�3z�"2F�@�<����}ԢR�jR4��\�3��{�<I]��1G*cm���҈YEd�4�ȓ35r(!�_�HS<�9���?l�ص�ȓ3��Q�@]��i�Q��)7���$w:�7,Z[Z, b���
x8���s.8��Ah�0i�t���B<O۲�ȓsx�E#A�	Kf�I�g_�,54��ȓ"M4�Y&��%y�E9��E�z�A��F
�i�l�";S邊�&����T�B���,��j�H�%N8Z��m��t���EL�j[�ɨ�g �*��х�S�? ޭi#MB*�ʹ��ʦfw��a"O��q�ɇ�r���V@��	a@!�"O(���W�Z�ʨ  
JM��8"��xy"�'nl��SX�$\R��
�����'���8�h�fF��A0��^�'a�dr��3:�h'��sH �'.�,y%��%�¸���@�����'؊�	��ּH�Б6AI�x$r�p�'	�����
�M@���	M,c�`4C�'	0UzT\+��izeOѩH�.k�'�ў�}���E4l�!l2u��1�7h�WX�T��B�tJ0I�6�"�� 1��ͨrX!�DJ0��4r�*�$`��Ĩ&%V�eFqO�6-�O�b�����|��D\�\�H"�� ���Xs�<U
^�6@�(+`���p� ���7�O���Č�HK�Yk��H%�ΐ�GЋw�!�d�U��AՀ����i�q�ϓqFh7m��0>���W s�-��d�F��HaT���'R��2DQV(�_��!iw�޲% 0�"O�hF*(�`��%J��00�!��$�Od�#�$m�e�S�S0E�5I�MRS�� | ����E�Z�<�3��!v�r���̇�-�b���O!=��>��K�O�O1OlT��h� n�^@A�M#�5�7�'��&
]�B�(}���,�V��^�O7�)�'_a~�D�5{c.��W��~�|E�R�
���A�~E!I>qߴ��O��|��ř,�ԭ��-E0/����"O��	��#{&���̭KY4������O��9�' �O��bKp�� �kh��S��y�k��)��H1�&�#v̒�5A��d3�O�4AG�7I�� �:�nt��^x��/Ol�FƖ5K�aa�!@���`:�"OĹ����	�J�5y)��Y��	|�����f4p9I �]�]�B��G�C^�Q�t��ɟ�4Ez���=	�l�X��=Dv����(O?iB`��#[�p8cv 4}�w,�D�<�C#3�� 5� ����v�|��(ʓ�Z�y���|3ơK���-�V�Y�$ �y"-�z~��y�.6X���[`�����=q�yB�U.ߊ����C� ����yrH�Y�&Ѥ�F!3��Dj��U��yR���{ّ&ɺ,�VT2��*�y�oK�x"���FO�5"֩z����y���\ݸ��C@J�Q3G>�yb��[g����� <�:aɃ'���p>�����@�SҀ1�A��/m�.� ��.�qO��$$�)���^�dp�@˗b����"�ʹ\�!�d�����t���=���:��5(�!�d)
�p ��
S�z�  j7,[�M�!��s�I q�؏?�`�j�K�5��Id��|"G�֤^���"�ӽq���5\O�b�,�52L\)�g�\�0���(T쒿�yb�ìYʞ���O��'����c���ORb�\�~B�	�d��\�q�Ū"�F-���z�'Є����-�|cR��.U6	��A�\zC䉯\���1�T
&e�I�F�0�O�7�E��|�O��e��H�LPH��ɡe�	�w��=\O�x+g����uHF�	bV;B"O��H��5s���I�"Ťk�*�C�O�I��98dt� ���&[����h3D����*���#*�"����-D�SF�!,��a`'غ�h5#��,D�����3]�E����8o�n9S��O�1{/OЍ秈�8}�v�ѝ6P4�b���}B�KO)D�t�4�MTGHis	O)l�yr�"���	d��� TQ��BY�Ed���$@9x�����'���*��H3P#�=c6PU��%�E�!��H*	�0%Â�
u�,@�צ��P�!�䑡!{-
d� DX���f��nr!򄝌����	��	�!���+��gLĽ��	`f
�G�Q����9z��d�+�������C�I<,6f�k�Ŗ�v�P�aҥ��d�$C��$ΐ�I��We�l���L����=ʓ1���PB�N�&16��͕0f��p�ȓ[t ���e���}`�'�ԇ�R�Fѻ���Q	�Y�� �I�E��	Fy➟���5.�p�[%ル;��X��@7D�@3p��ˌL����V������5D���C�1cf��`��*aA��+Ff5D� �V��4t!VEۅ(@5F1�qBK3�������)���``�$�v�Lԣ#"O�`��bϟIP�+��.-ޮa��"O��k�k��z�I������c�"O���T�^�f��C
D�R�t'"OD���Ǚ ��e�s�A�(�,���"O|�2c@ߘOs�a�fءy|re��'����0��I�[h������5�L$�=}�Ih�'w�)�%A.)��2�!��GӮ݆ȓ���37�B���cj_yn)�ȓt5�P`��98D��� �O����II��ug�ɪ��u���m?hm���"_�:��p?yp�+	Dp��.&5��h�,�w�<��/Q���љ��\�x>��AnL8�`$�00iS���zv���7�f����E���xҪ�-,�HTT�=�Z� ����y��� �c��D'�|����"�y��L��a��
�$n���Cm^/�y��^�1Ƙ-����?k,H
s+��y���	��	�J(�ĥ��D� ÈO~���6	~r�ȕf� pV�!Ѥ�T�<s��>�B��SO�G*��s���M��5�S�O;�M���Ap!���L;w�l� �"OdqJ�l�`p�����L`8	1#�>Q��0��3��;J�p(Ta�.3:XI�?�����'�r3Oh�C�LnBC?���xF�'�!�D�s�𽲱$I$x�$�q�& !�$�v�$[5瞞x��:��ڔk�{b��(4�⭩/֗M�r�!m�Io�	W�`
F�\6����ĉ�l���.D����F��ev�a��B�Y��$,D� ��Z�(�e�T8=��@3�)���<9�'(�>������b�]�X}dT[WA#D��10ł�z���A���j� l��!?�#�'�	��&]�G���F�Z�f�Z\�'��ܨ�(X�L���I��HG��/O����74�h`v�� ,0�1bJS��y2��j�I妙SShе@&�L`Њ_��?D��qE���E	����$E$L�س�*�	F����1OD�9��;Hz��� 'qof|*�"Oh"E�%�8-pa�&HhF��"Op�%C�9�^��<�t8�"O�@b�E��	6��jt)��}�҃"OD�!���朱��å.�ʱx�"O1���=��X9TH�'KZ�9��"Op���	]�'��q�� �	�� ��"Oh�3��i� az�@7�T� "O
�T��j�xш0 ]�8.��3"O ,) ��((�P�g.E�x��it"O� h`�̐gY�H+���+l�L��""OV@�ڂW��yՌ��̐"O>xqr�
!h^�U��*�B¦q3�"O,�"c�T�M(p"SA.jE*a�ȓ6��y*Q�*�
����*�لȓX@���%H�&vr3f̡e�:a��:▐r�	��i�����OM�gD�u��V1 Y�& �p��@���ȓ8�]��T.C���R�D�a�ȓ6%�a�O��1ۓ\�H��ȓK.��Ch�z`b�N��p�̈́�~��}�!ܼg˸Q�� �ir��ȓ ��=b���-,BXW+�	Wd`���{�����_9f :ǊX	KX���ȓ����3���Z�q��>7�5��G\��/�.2~е`;|cԀ��`�L�����<ۚ�S�OE90�@��ȓ�ܑ�蘊Ze��+fLU��6�ȓx�Ҭ"T��&h���C�,�ȓN��ԉWA��IF��A���"8�ȓs-x�ۡ�ע2j����9��@z�'L^�`Q FS��(�@�V�d�����'�ʌ���B�.@x`���� e2��i�'2� d�߭w�4� �р'�N9a�'�$P��D�U3"m&Ț�#�ڠ{�'��%����AhJY��J�*��А
�'j���b�m��pS�N��
�'����4gت$�Ń��xH�	�'�ua7"](e�б�P0]kL���'P`�W��49ڵCRb� N�pI�'4Y8s�Y�kBX�0��AGb���'�v�����\^��rq��"5Z��'�H1��?E�0�0..'p��`�'��2t �$,A���W)q��P�
�'\vH���,L}��P��e.�}i�'Jz]�S�U%��1��)4��;��ˣu�\
cAƓ&�S�>jM!�D��Ql�Q���61�bHYS�]�`)!�D�!�~���ۛ�x��c��6D,!�$��>�̠0��\�y6���q-!�$-C>\��lo�4&ˢf�!��G!6E��! �L	asf�;3!�D�� �$њ�)�`�`LR��0jg!��7V��a����ۆ%�8{!�
�9ݦ��C�X
X�zP��ٵSc!��P�>���K��z���V�-!�Ć2���ۄ�]�%x��E`�7u�!�$���n0QvjҬzUNH��9a�!�#,ƹ�L�" \2�[Qǜ&{.!�DXwbi�fJ�m�-�t��8
�!�$!&ް�6ț�QF�)7��M�!�$҉9�@�M���)�&b!�d�,KZ.�bE��h�XR�iP�	M!�d�Rir�R��t 9�d�Āb3!�D���8aU( �h� ��g�Y�!�%W|�q3󨓽WmVz�G�$�!�D@j�&�F�Q�f�����&���!�ڣfY��y4!R(>�<@RP���z�EG ��s�C���=y�]�Ip�a[ԏC.� i���
j�H�o"lx�&(˜]TV5���$�,	c�/7�v��D�=a�C䉿����t%�=�L(
�G��^w��(�d�L��|��OF�;q0U����](�0��cXN)����I\3!��\�'���%���Pƌz��e(��S"���^d�H� �)5�~-a��JX�I)p ����Ў8�q�BO/zs
��$��8T�`X���Va��:���7�2F��a�jDBUƍ,0jX끮	��~B��3lf��?� �{�!��]�dE��Z-�l `��	�fHe�
׶uļ�Љ�3��S��J�;����$�X�g�$�
�K�J��0mڱ��3�]��z��Q�TE���OG�8�B����~�J�4.�TrR� ]�u�|��M�`l��A� �c�^9���_�~�X��!�	~
Ib��� )�a~b.�a�L�;�C��y��u�&�"e8��43 0���$$`�q�l�'��i+��A�z��y
�fٖ�2M`2Lܷ9�w��CLR��b@%�d�8�ň��hO<��"ePVk�Hd饟i�.�`�AN��}���s �Y������ "�p�ȧ(X��E���_,z8����x�����8�$�.0��m�`��	��ЫD^���ڹo�,HR�~�̓\c�����O�!�-/�P��Eo۬3д���ͺ&�tpcM
5(��=Ӆ-� >J԰+��2ߴL��m�sX�H�Ǫ�03(̨UZ�.�^E[e��<�'CB�]{�Y��շRJd�w��2{7$А�ۦ.�Zu���6~��y��JM�m�`�J�]V�$� �]���=�EE�J�]�Fj�Xl�-#�f�#۞��S�O�l�x6-��ao��04B[�Tv���6e>T�"�lX46��U7w�MV�ĭ4��4��31� x���N%HbFmр剖-���b��4�X�Ђ�d���L0=,&�KW�ћo�j��u"�Nm@p��t��V�,]*d����T�'8<��AQl�z���"֞MkHh���OV��3�Q1-�^�.6���E0 +D�1��t"B����R �I��UyԨ8��!�e�2!R�!�S�D��qe�b����Uy�)ڣ\�!���ϳq��Eh��%��1�5�I<�D��¯53�D�Z����T`�Л'��dcL�,kެ1��9�\��bM�5�R�b�F̙V~��3�D1's��	 �ʈ^�l���ކE�j CBGZ�G����I��8��Y�<٪�{5I�>��C�Ai�`�Z���9Q�F����3S����o�4G���)ԛ<��1#���o�|�
��;T�Ha˕�+�ܙK���*�����ɟ[�DA�5���ι{��E�<�ݴo����(ӴE�J�#�����l;����.�*MCt��>@�P��q�5T����R�6B�Z�CT�Ռ��p%�+�<��W��(aξuX��L���Z��~wP�*f�څp��Dؐ�I*�?�G�ũc˴ap�+̄����jV�{H���h\�l���K;P�2(7�Ӛ,����@�.���Ce*� t�$��r(؁Z�"<���pS�,��BT�eP�%	�~�"E�#bWh`i�E�T�,��m�&uX�&��AU�yp�e�#y�y�g�V'+>�y_	&<��!D�^���iK`�ZG�	�mLT:QeZ�b1�SEG�_\�H3�[�Ih�%�װ9XjT�Q�D�0������1DHn-�C�%WH� �+Z>Lb�=3tD�1;_�hB$mDH�P	� *��q��@��I�UM�H�ͅ�N�N%°jK��)Q�(>��p�ϖ	�Tc��J�����һ��XY� O%05���Dȁ))2�� n� �|B�c�(H���"@�B���BV��`5�`@^���S�TWR=k�i3Y��>�>�!K�� �H2$��p�IP�(�,L91�����a.��q��D(���\0O��0g��3H�&X�/����]��
j&	�ğ�Ð�H4r1H�yb���ADX�f���VNF�5EX����A	
ٮhS�j�l�@3$E�>�����
6rI�,�]�\h�����P�bKB�N)�U�D'~���O�G)��	dlTX��i�	X��J�E�R	!�O��W�)"�a�A��s�`��V6�ԠF�:��(����#�b߉�L��>h�T�[�bA�1/���!��==ed���m�~怤���3|w���#�ֻ�r͕'��ͭ�:jx�����}ኬ�6�X�|v���C�߹='��wi�wւU3�.�& �䭣���t��@`��ٶW�T@rm;8.��A�)�wؘY��&"�����&�Ɛej�# @$/���lZ��Y�"��@�̀J]������	G���0�͏r�8�$E[��b�p�%�3f�HMܐf�٣g��mS�!!a�F���&a�>{ �օې0`�P!�\�b�9�'Q�kX�a��D�R2�ᚢH�c��m��d�o�@�uX�+��	�/G�`�V�ŚV5��(�a��q����i�\�AE��-Jt��2��+���9� �-r�Ɋ�G��wfb�"a���w&����߮Ly��r�OD*�N?\�h���+W�(6�%R�!E1�%�"g�)�d5��ڢt5�	rD�[�.{h�����-?�	��#B<%�~R�
^ ͐��F�FY1Ć�6֜��aQMif�YI<1�C���Ԉ3�I '#��pWC��8P��c��<��]�!���)���BC'l06,�S͞���Ѳ�ߍ.<:h��O"ȨumLW�rP��'����
t�!�#H�:5PE�I��S�ˇ� |~��c��K&izѮ�9@�b(��G�,>�5  �c���PH��){�P�kO'��YjVL�7��&eO�jDx���#��Lļ�)P�wU���$�K5e��Y.�{�c\�]��M�PQ<id
]�!���!0ҁ�e��
��v�P�^"�[�#|>I�`�Q��ADIǔNi���&g��b�X�C75�8P;�f�ns����v@Z���·Eb�ԫ��Q���o��H�m-r	D��*L�\�,���O;���2����M��\����?�̕�s��/uP��O�̙Ǯ�igp�+���kФ�B��e*����b�"���m[�W�4�SN��q�͛7P�� <c'��'��!y�����ILN'rq�SɎ+R����v� o�����8���bu��k��<��͎O"z}�۴Q�dM��m����  /C�Ԍ�櫒W���I�%��y�	�m�&�HuH�QH%P�A�F�ĐцKr�ݫ�"+ b�e�KWvn�إ�٣<t
!��+-.r� է�^/�7��!c�b��E�����S#=q�e�N�(y��^�|�%J2jM�fs��2���b����iP!!��hz&|���F�}�!��4���A��Q*n��W'�4d` Ñ�i�d����& ը�p���=
����� 8�\e" -J��"L8��>�d�#�mȠ�Z�c����I�L�J��皘y��Y�ᎬH�Pف�H=Dr��I��e��ʜO�P��G[�����,D-(nu!�oU�:cXY�h�$FJFؚR��3�TO���U�A/*m�Z�'�-���DH	_[<����&M٘�$���A��� �!J1je�D�4-J��Z��T���ʤIє���+A��'F��]B)L�vyʹ!�>4��I�E��T:'ݘ$���*@��A�i�%st��d޷6z`ΧK�DJBI��P0b�	F��F��Aa��'�l�0E#'�h�ɗ�D��g�w{1P��5�`�P&^��V�w� #�l���f���C�,Ռux�;4�n� 歟?�B�`��Q�K�z`Q�-Ԇ"�]X�#�:`����G�G�Hy2/�ŦR'l����O�3 &y5�T��
�J�~���͆>���S�����4���%��D�S���6$`���ˡN�l�C팄:���{�AB���@`͆~l��6&�$��:3�� �d����;�@�g�܌oj������5�^�k��̴2�F��Ge��Ȣ��C�4PLxK��y\HÁ��8fbAP#�����
�k=�QC���	�-+��lC0X+h;��P
����̷Đ���Jq��Ѫ߮-��@+ଙ�]�Ѯv,��9� �XrF�>(�<��i*~�8\`�P�DYF`�.M�^��a�L�?���hHy�4#�ꊩY� ��3�����`�@�I�������is�-0�S?=;�*J�]���C�aލ���'&�6Lj�e�3����",�*tNu��-��Ahd��eI�����dM�U�3
�"�,�`��M�:��\c�M�Q�P92ȃ�ppƠ�#��7U���`�J�!�8�$��� E��%�!�0��!;�H���G��E�1p'ʐ�
H���Dl�ɠ	@��l-Hr&����r�)� ��%,� �w ��ʷC��x�" 3z%�O�|�r��~/��X�� ]$�x�OE��c�T�0�Ʃ"�Q�^��#�O��.��@����眛'^�q0J��{�^	�ho��Ǘ�^���-W�o����l���M�B�;E��ZF-�9�����o��MC���L���PO�"o�# N��Wd\@�+޳�E
�FP8�l �|"�Ɛ8��	{�0��uݏS������F�N������Z�����ўx��h�?�Fz�i�4�f+5�8>�rDJ�X6I���j���0Q$���#��$%��m���|2�G$'��q��)O.3�Q�7L1���O$�b�K�!^�z��m�$� ���҃�I,�Xe���Y�r�'�W�؂�.ɓt*�����:���:��>}4��'��tL���OĈ{�A�
U�(��Cȏ~%"�y�Hx):q��1v��=1f��;U�0P�/^w������֧k֥@������(�L�+|U��T��;{hht�@�S5�P杯/@(�B�8NJ�E
�e�T�Ғ��3P/�G{��iF�u�Ľ���D9u/�����Z�(` h�o�*h!\�7ؚ��������t�£<A�ڼM(��0jA!"!�30G
�W�a|�`]�=Xƌ�䍟�!4 �W�ZaFp�/I�h��1}Ј̹�IZdJlӁ/ N�xڴ�'�hQt&^�)�x��A�^� �r�b��C��b��>S���㎼I0��D��$��������!^I�L����0= V�¦ɀ9�8�Ez�Ŧ[+b�'�?*>H�/�N5Tp�b4x���s�X��4��`�(S�˜; *  `�U?9�*�4"�T2���kAb�<V�Td�ႼA�a}��`#���"N�{�0�ȅ�C%X�2���/%#���g.G�V2D�P�Ƶ��%��Uq$�	6
��Qp�'ߎ@��(��ܱ�ԠH'�y��h*f�j��И`~�4a"�	�z�8�2�
�
J�1�g�Ӧ�;�O��Z �U�6�D�rC+.�	:W����C�	�D�!:@�NPȀ;Պ퟊��C��d �
�
E/BҤ��8��
_��)i��wynH)�̀`�'�T䘧ǂ�7N䌑c�I-A���C�q<�k��>��J��<�P��B=5I��ɳNn�䁻	ͼES�JZ�!|𨒂�iM��p�Z6F��QF~��|����z��V��=��EzA@ъ.2�X�1V�h����I[%�?aB���2�Qb�'p@�����ŪH��b�8`�je�I-+�Jӧ3�Jȓt'��.��`xW�R,T-2`*���xv�x��]�I�@�� ��#u�����"|X�[��б$.f ��K
b㾝�G�x�����]K��N�qn>8z�Ď �uYQ,���D3t����C����]�f�ѿF��'6. �r"|�n�H�.T�'<�)�"֏i��`A ږf��M�E�ПU ~���E�qY�k5[=�	��j��t�=	�H�%�,���<P�(Kg�D"b�.HbыRo�'�T��w�Ü`�6�P�'�8�ऌ�� �k���,/<��ڃF��ː�P�dH��$������ák����`�4$V�ģF�| ��&Q����Y">j:�vϞ\�T{剽ic���&\XUH����G1VT��hb�LYaxb�_�E8���"n�([h��!G4�yF��xD�����UP.hA⤒�a��`PǄ�)��h��"@:�I���pJ����MTU"H	BēN<$�S"Ɂ6I�]�4���2^Pp�'�4)���'��\�%H�ўȓ2���,
�������X�*_7�T��� -|�,k�+�$��U�U#�)~����	�]~R�#F�y�0[�C]� �0L�u'ĻPbf�=���^!�D�h�� <�|�Y�[~���R�� u����'b�?�G��*D������mz꽑i�}�,���Ɲ�#N����>�DM:%B��c�R<4�,��S�U]ް��<C�0�+����|�Lt����jF��	R#D�*?&�G�a�;i^�)�R�I�٤�0>Ofqģ�[�|���+޺%y�-�/�A8XH������c�g���`ID�6]�f� �{�	 Ut����H{7 ��g��1��˓"Z��x `B��|�w���O��"� hٶԱ�☨)��t��?�D��m
~$����ˆ:m����1,"��I��{ۊ����{�N�KcCi�R-�I���Q�_�~o@l`��a����c����Ч���!E�M��ʒ�q\���ݢWT,
�Yt�� ���([��+ceͦ%y��۟R�B����81T�X*�3���E*DZ��>�D�p�E��v9��!i�J�(D�1$���Q�H�M�!�5�.)0�l��`�D�ِ�ᴁV�^J\����UM�p��	MnY��`E�>8D�{���ՊЉt��X	Pp�'�|�bQ5c�dIQ�,Tf��YJ�Ol���B�)�<ћ���yB�֭*"����R>Ne �0�CZ��	� P��� ��8oT��E�3�-j�
'Ҵ���'(���3&�*[踦+q������+?a0���\- �k�ME�HD�qC�T/zHoZ�tξ��W�:��9a��0����AK�F�ߐ��?rB_�z�$��2<|�6����ߖ����wm��-���J��~��i頻�Ɓ�Dn��C����h��υ�ny8��ao��2��1��yl� ӓR�y��,}�c]�0I�SA�,��pZ�C;0:��(AAS9`��r�M�a0�#�]� i��A(��X�Ou��g�42�=������0���'�uZ���\OA ��;���������q쁳�v�+R� t��a!	����G=�0<� \�
c��f�$��È}�D�����x�Lh"��H�)ku�G�n��Wjť&t��$+]�Ga� g�+����Ʃ�F�Խ��6��A�j�7%6��A�P��s��@���m{�����l�[�4��y�ʘ�$4ʧm��e���g��q�j0��o�+�!��
4�$��jX�>玌�Ѭ�\��$QC�II����s�H(ΎX�8�� ��*ػ?䈀&��ؓ̍1D~U3�@Z-��#"�Ot@ȑgO-ڄ9w\�-E��J&h�8,��}��'�d1�-��@y�e��� 9�0�N�s} �A�H�3����	��iƋ�
 ����i��ase�f�!�čK��rϝ*��q��&��E�!� n���A0d��w 1� D�!�H�r����G� )���+��W"{'!���><�1KV@I
�d
=>�!�dKe���!%Q2e���R�"�!��^�!�L���M��	� O�z�!��8@)�u��X�<����4��$!�!���~5(4��,Bj)
ӯ��!�d��T�VH;��:2���'O��!�$&`��	��A;2(�R�S�e�!��K�]O�Yz#G�.&<!ɳJ9R�!�D�".��s��"F,Y��o�!�d����0�L`kqMF�QW!���K���	K:cj$�MD9N�!򄚉5��r�#o�@�3%,�!�P�{�4�
`��l��F���
�!�˰Q��u�󢟟&h���A�F@!�K�.`����.rLXJ���T�<q���7��`a7E�m�<@9�(\N�<���Mp}aC@�B����>T��I3�_C��p�#D7c�!y�($D��`3�M�h�ج
��K��5�0D�Hi�D�JP�݁���	h��An,D��kl+-�ɵ�B�E��x�L&D���w _�=b�,b+�"[����%D�l[q��+I�Y �MB�: ��&D�H��m�t�4DC�?j6���%D�,2w	�W?� ap �/ �밉.D��qG��~p��H7@�)kȑSf/D����P>|�t�g�2╻"�-D�,���Ϝe*����bR� �𡓁�5D���!N��6��$�P)n����T�3D��s����\eu�'�|ȩ0D�����@v7dX�(K�%01�T\�<y�bڮ��aT�X o�T;�
 f�<�El�4b�p�Sb� Q~�2b�<ɂ��;����͂UĎպT�a�<��dQ�
�#2����[]�<	�J�ny�d�	�g�4�1��DW�<)��X���C�
(�>dA@�Rj�<� j� #a��Q�R�$�Z�i$*�`�<���ʨ)B�|�Q�G�J��@1���J�<�֢UQ�tMD���;�NI@�<9��H7�Śs"�L�����|�<A�GK�%�|(%��F�6(J�`�}�<��l����肪$mb:x�o�s�<Q���l%IU�Zv�[SYn�<��䍙D���RP�J�k|4�#P�o�<!b・By��I����,d�u;���M�<)")D�Dr�!�%������0�I�<!1!ݓ����M^,szT9�+yH<A焜�1g�8�͞ -��aX��Q\�̡	c��1����k;|O��+G�JP�Xq�'��5h���'T����Pv�I���P�<�Α�&�D�1���zb�UJ�Vx	dP�y�"�F�9Y6L��J��<����#��DY�L� ���`>�ơ`��oL�#|� �$�m�;�P	G�:"ٚ��a"O�L�C]�2��`"E�G�xʸ}�5kϵ=�ީ�'Sd|��l&\��O���$�0
�e�?�ԡ��K~ ��'/4�O��BtL˒"�I���^%e����!� �j��ݖ��q�!�j�h�'��`��p��6�Xs� �BXj��`��=OB�F}2���U$z$��A��Sd�2�H����M��@�!y��i��F�J�b@3�d!o�{��D:G��A|�]z$)��)�� )�l����/�!MjNuY4Hb�4�{�@�"=�(9�\wRqa��J�LX���O�q���AJ��z�#_��8ڱ��}�v��EN�!q�\Q��:U�YI�g��Y�(z7�KP�L��%p|��%�� s�XA5- >_�m!Q�]� �v�nA�Д��-����>ړx����&�D$2-(�'�v�{$�"��l��+;p�>HpdO���;�͗I���S��BC�ڝI!���\�tk	�v�$x L>iB��=?c�9����> 	Y����Q���:$���w�@" 
�Ē5yy֔+)�*x Jb`lG8I�Ǌ�)�.T��!v�f ;���:���rAB'oD�8*��F�!�.��� ;r���'��0�&�٢)��i�牯~�az�B,�>�� �<1`ܒ��X�2�:�т�+`��;�N';5.��!D�Uɪ�C#� t�p��00("�'�%><RM"����!:����l�-U;����i����d��2��!�5�7#T����*�/D~�	Y2^�bls�eJ(J������ W�[��֍)Pd cVo*ʓf���B4�Q�
8�J�?q�J)F�vE����0��ic�O6�n��w"�JVI�Kِ6��H��OV	}&�q�d�D3��%)�N4�b��G�\ǟ0bB��-�H'��Ab���a#'W2](q�r�޸[TfI0�ye��"�(�lL�Cg�(�c!��"\6�����%M��aF^�3�PT)"���_���rȟ0l�=z3�E Gp�ҕk	
�HO�e�2e�
U�9Wh+>0)�J��<�p倞0�rI�B"��M���X�Y���j-< I"
Z.VRuyㄈ3gj1�*�j�����4I� [榑���O�  �M�y���bhВ3:�:�L��VXx�ȁr�-Q�)E��u��P=�Hg(��50�
���QXLz�I�q�1C�9I0K��$Cl ���"�(O�'�U;L	P匥Ao"�Ц�W)J� �i(󧓛b�raӁœT��Y@�Є4}<�q�W7Z&E@�a���}s�d�hQ�%P��9�ꓹS���2k�Pw��Z �(�>�;qE
�,�ҸZ�',&ڄ��9Q���b�L�Ru��b��̪�$�{���;�D�Si8@aA�2��@�H�<���9!���.N@I$K:�p҃�I%v
�XL�9m�P�)W�D��dA���L����u|\L ��'}� ��Źj�P�!GD�r}��K���-,I��D�z�(`���~҂ݺ4�!�"\���K$i���h��/�*5��b��D�ѫ �T��I�"�_%�<Q�� �� $V��i���[+�9N���c�Ӣjb~�(���Y:6�<���S��ٳ!omh�6�~��	�ni� �����m�	�b��b�>\�.� jI�ZՖ����&؛��â���Ʌ���_}
p���M��d��Le���I�G |1ڄ��τz/��q���Ά~$��i�lߚy~I���l�=�Q��&x2tV�Z��yq�Z���x�����G�t]ᕭf���N�64H�h�� [�V	ck̔��^����0V[�v͘q&h++�:G���b�JK-�؀��B�6���3�oͭg��܂�
&+T��%���G&p����<DR1B\6N}{�!�7��`J�$"�i�m���2	� d�p��	�n�"�_S�<����1����P�֨C��]!LÙn۾�pJL-�x�b��^W�2���M۱����M��Y7ZIi��.4H̸Q~�U��g���UG��]'^9@yI�
گ7MȨqDU��rҨ��I����Y$F���h�扒%��\�����Jg�e"�3g�$Y��̄	J��d��&C��@�ƉӼ;���-=��$0�d�Tf���'�Ŧݪ��ڞ�����J���XԢ�G�_����MS~Tt������g\`�IQ�K�"�'EW�n~N�PA�'�YȴM��Wr���G�mJP�)PN�0-�hOW�P�)��a��*��E����YE�՘a@�0&̞�p�V�Of�ك�0z�ĩcA� ;t8�8EEJ%	]x8G������#I��QQ�l�@e�r�<�ȟ�?�"�P��'U��?}:IX�J��\�u�� 4nJ�VM�g[���5��&{n\�Va�b���nZ=�|�� m�0�h����[ʰ��� 7"�'8>a� 1�hYjv�ՙ��\1I�';:4�Gݸ?e� qRɤ	Şc��-dئ$Hg��:F��)E�M�sh��nZ,�́�gɘ9��;1Of9��O�,	3'��3�ĭ)��)iBe2�"��{�H�C�HٸY�<M�I��h�.Q�u��Q��c̪I�Nx�4/RI�'��-*�Ýr�
����O#�pHAo��6j:�m�VyZ8+�I�%�IK�';�(5��0T�R ��w	��I��,3����ѽ~���� @�A;��Ҡ�	H����	;��O���'*I�����ԕ>1�%ӢC�8�� CLļ�@U��Z�(3�y��3p�P�+0N�;:�	�J<�w \�/rƍ�Uc�=O��4�ȃ
rkT�\*[?��[@��Nx��pg1G�̡��#����D�>�%�w�U�$�����
q�Aa�H�?4
`(+��<x�<�('�����Ix��m(�V!,�G���c�L�W�}X��0mJ���3��T������(�J!�d.O=ob�"�+N|T��p�i���q ��[���H�D�j��b�
�*=#��~��)(�`)�@L�1W�ň�	<B�~��2o�¦MR*�����:fTH *21/�|3EOW�~`��� !&�7�ŝh���r�#��t���*�\c��u�n�?@l`ja
Q;�� 6�N
Z]��[df�#�v� �{���5H�$녩�| ���/)E�%2��� E�=�+�8:���j��5*5��~�Rѩ�c�/�,� R"@��'?RIP1G�A��x�P�۰cy̘81eL(~u���5��'ɤ-c6��Z֘���[)�X�l��bz�)�xt���բ�%���c6�	&�Tm���p\X�+w�_�g���pRl5��N?x�P]iQ$�H�H(c�
�u����w,�]`�A�>�P�zgʩe���ņ��0e��K�T�sy���@[h�	sf�?�T�r�~:�&��$��*�*Χ5'8��e�@���S���W��H2��B_��[S�R� ��8r�i`ZP s��|�7o�.te�Î�Fn�� rcƥ.�p��?�)q�F�!0h@�J|�>�6F�tq�ƃɜM�
t�' :M�Q�I�j3������{5�#D~>y�cɞH�H��@�=B�u�Uh�nx�#n���3��_����F G:@��m�3ubY����Z�d�Z��'� �42S	�B+4D���A;���6 #2���a¶Zbx�a�H�h�b�i�F"&`��@5����@	!7��X��K?btF=k#�>d03�M��`�+�y�l��r�s�U12�" 	!#�F��d�a��zJ�����|�� !�W��,���
� 5aA��=�P`%KhӀ8Z�Y!$(@��t���<%FYB�#��AJ��J��?�s�Ԥ'� `bl� ���d�@=9/Pm*"�jӊɻ� C����M!*[6���S1O����F�k(�����H�oϜ42�QS���*6,z��&e<vڑ�	����Bւ+fjA6#��h�F��=Tn���d8z�������6|t��k�N�2oHh�e�K;Z p�G�y?is�˭`W:������O8������9N�K����L`����"j����aO8E'>�y�lE%N�(x�	�-��sD�[�I�,��3Ԣ7G)ԑ�Ġ��Y�&@E�`��Y#Bܸi�D&�\349k�N�A�oBSvϚ7F(��3E  ά=(�(_�i�	�`�O=3U���:���2P�P`�� ��%�F��@�a<Y�L��$[�/LR��F���D&ڌpy�
�7.A�x�C_�(`(�@�Ȗ'�^`�O�H�w��V[0��̈́���Zݴi��Y����1P��Q���[�E�ܴ5�&1w,ޞ[��PH G`��bClSw��́5JH�t(���i�'q ��Q�ul�X�� �.��~�Z����T�U��\�JL�0��5��.�.hTV�l�'�F4b�CW<�t
j�8��4+�#d;xi�#��s��lА�N��'��`��!S�M�R�Ȍ;thJl�&K-u^����*
k�֌'���-�-��i���^+n-�B.��$@"���?s��a�t��3!��(1��@�cv�ؤT졛�B�@���O�:�i�KU̤�&j4ay����y2*��`z�����S���=i�iN�oU�PB� �./b]��N0ioZq�J !�سBbW�(�,æ&U�nT���(uaG�6���]6V6 BFE�2�H9���W�P)~pK5�R�e�RPD{�����p��	�6΀;�%b��8Y��:	�m��`�Ѡb�����N�q���<)�f�(q����m����(�)
a|�)A�X�(�a��B� �g�ON6I�`�>:k�H!B��~������	�N:U�`�<>l�X9b�'�0�Z �aTm*T�)&�TTX���	C�Q�u`��7,ܜ��ȄPN�-�Xu��M�=	���RK[ �:I�4)GV�I �I��*,��mFzR�Yg��-�lP��8�z�*I���0�I����k«"��t�p����%�T�P�,�2Zz8�IZ2�`%��":e#!��K!P)!e�P���	�R�2�RD�	�L�"Ċۍo�`�k��C*aH���p�ŪG����m�=ֈO�q`���䨅�!ˈ�U�\�k��]��=1�̔�1́�U�W. �'΅;f�`1	у��ZzD��a�"��OX�KV��0,���%:"6MK�^�*�&��~��؆��P��O��(�U'L:��
�0j��v�[�w*���?="X ��K>=��Y�B�y:���OjR�<�nl�����	#�#=A��S?�=2WىB:li�E�`��bu#\#sˎ�XTc�sU�5X&�O=�)
�LD7�'���`�SlʢY9plǊ���Xw�Z�*-�:���D�܀7j��.����0B��(��dO~��u���/�3�I�<9�TS&�4��%(LT�
¢}ˇ���i��O9[U
�3m����)� �8e�Ac�4_O,����زO^�1
Ǔt�t%�$f�9g�0a��`�O\y�݇ny����^�D�^���O���'�\��7�	&��Ӱ-N55���{��T��Xi_��$��+"�"�]9H1�{N<�%\:p�l)�L�:��=�U�P; j踩P��za���EY-�cB�ф��g���]a�a�u�P�"l椑0m(�I~j��bHD/V��P�ë�<�|1����*�F">���U�	rly�QgS�<� Ka�Ԡ�!��Z�`�R�Eӱ~�xQ�K:�h���'�tѢ�ӎ�b�2�	d�D��Յ���d�L��E�P�Zu$�8�h�@�\�h�=_ZM��G �r�jk�S2n[;�KId����T�Ɇ!A���8-���ͦ8����a�0{�L�t	S��H�c�މF=��l Kb<�(�.';�����䐲x�D	�dfSP��`��/ҹ[��M��c�1��iGϔ�H��I�h4��rT�?V�2}�4�f�'�L����%J�`�2�*@�>�ڥ�A�)&�x�`ȴ/�2����\�X�R��	G��K��T�{-������0���`�k��Q@X���B?�|���a��/a>��z%��S�L�y�'_M����P*�X�W|�M�O=\Oǔ#V,�+�E�%C�~dy�^�O ���̫�PH�j�=sˢ �4�R�?�����B�B��Ѡ�)2�&�����0�B%�}�'����B�~0�d��1.������s��.VNF|�
���n`�>0X�U�D�o��jˇ�����C�-SFH`&�$ ����J� c�k��z0R�(�<d,��<.��(�P�����$ 3��h��Q�32��7���L%��b��Y�X�c��}$ ���Y��p<	č;���"�@� hBK��Qd�
9����ަժ`�I9��Y)�b�0R
�S���
��`����u� ��qiK�u�ؔ=�$�� ��Aca~���!32 PxMѥmH|�2��e��ͨ#G�$�U�V֯w�̈af��:}�f�!G�E��td�l��U���WN\�bb.O�i�NҾ�>�J�J��y�[.f�Vp���S�!�����n��b߾�j��&J0} �-^�h�m�e�B@�`dR�$���p�����H�/PŪ\�l�I�L��r�/?�Nٵ�����E�X���
�m#�Iߊ:TZ��%i�/Nw��+a�~̑5	Ք:-nT��ქ?�Zd:��F�\�Jy�s�$:����52(�D�5_K�$��b���G�L��t?��F�J
����k��B'�O$�M��h٨C�hs"	�����Y����A@'__�T���'���䤇�tKJ��׊��Z	�D�iHGhl�խz����� �I����d�pC^������L�T��LM|� T��b�M܀hrɯ,D� �'A6����V�d�..:�`� �X�p�W&��a�4��B@�G	���u��4ym2�0�(.,<� T �\�X�ǖ��v�$+��(�G�[&0�h��*LO��;����T ,i�eV�g��e���9Cj�Ѱ��f�*����'hì���@�̄*�
91ax�&ƞ}�NL���LԚ
@d-�k'�	!�����?�P���OU&f��X B���Y3�����>�x�vj\�%�N\0JAF��3	�'�:��S	ͲI���dϒ�^�q�S�?��<�D��)J�*a�����6��#ɍ�K���OAt�X�.t�7]H��4�t��e�tC�	, ��6��6S.�,�"mV��^��bP�k�t�⊢(�`=X��u>���
6R,� �J<��jlT��gőLlr�B��JI؟X!��Ý�X%y�L��jXڶ)A&�p�O�}�f�6L
F �ϓ $�Q
2S�Hd;`
�g~������?��)�`�k��}�6c�^�\��LӘ�C�5b��A�6'A�Dy0�
U�Gk0C�	�O�!Y��b��+C _�~*C�ɅWu2hX7BL6�4�P]�(�C��d��(���,�(1x��ڝDQ�C�I�G���� K�H1k�̒z0�C��Q�0:Co54Y!�M�{H�C�� S�T�1H�J���G֊L�dC�I2_,)h6/�9i��hP�aÐ�XC�	�H��5ҤN�����k�C䉊fBe�!C�?s'��� �\��C䉅"��[R��l|���%�M��C�	��"�Gϳa�L�u�E9-�hC�	�>	��`��"T�L�?st�C䉟xI� @�ңh ��'��PC�	2T5Ji��I	(P��
U�G n�<C�	3u����JӃw!����/lFZB䉅wynɊV�T�%�H"�g�$I�0B���J�"eE�4�]@��ƒQbB�I :t`�Db��<G�`��n�C䉃U�Ĉ�R��i	�l�Ď*!�C�I./L�Y�ç@6��+w"���C�I,Db�t�
n��;�m��`C�I�	jr����a���r�n�0=2B�	�C�*��a�X Z�q���<j�B�v�c�aȋ_2*�ka@��VފB�ɗe��[3�
�?�2�i�	�B�I�<M�qV)^9aT�v�E�h�bB��tc�&(�'D����J_?t�<B䉠Qs@@u.ح0@ �i���w)�C�ɰV�u�g�Ă$�=YcY�u��ɾ*AT�t�̐󀌙�w�$�=�#dz�I�Teݣ=��dd����4J�gܔNT�9�.�@�����dقF���`���+mx���l�-if��P!K&Q�����O?!ѡM΄�51��	�(���j�D���Hа��S�����O?��19��(0�ML�r���S����z��ς3��  �{��	χ 5�]c�ٷ � 9*�3�x @#�u��h����	vz���
)8`�Z�����p�dӰ�0|J�KN�K�q��AT�{�29�s��]ܓD�豈��?��v��8��W���'���<��-_'��¥��R-�<�a�Jy�Oy��`���2�6u�F�2_�́�G؉vZl(�'���BMNt>}r'����`K�"U�<�8U���wh�	
���	։� ia��J��n�A��D�6X�a�#��~b�N&��ɂ/˗���G�$Oն)+|���`�	W��}���`2
�G�d�p�Νyy"I�C!@�a�$��w�"ܫ�H���@����SN��=
p���Q+K4
+~�ɟ���엮M �mJ��8`��� �gҜ"�|���tkvȘ�{$��S�A�BQ�Ϛl�|�h�n��V:�T���M��W�?aU�3��]��!,��E��`&5p�Q�G�5zOb�Lk�d/�''��H3�lP��\�
p-Ep�1�N����'���kH<�R'>t��XX���#���V��Z~��xF���=E�D+3D�^��2D�
[�Ԙ���@�ybɅ�/Bf��=E��d�L��9�Q@�i����pI�T�tI�ɧ0|ZW���.���f� ����`#I1u��l�<�p	q�O� �ƤA!4����A����S��U�����{��t��3'�KA*	$��BD%���4�O� Aq�T&l��R�!�=C�f` "O��a�.�ڔ��A�d�<dy�"O��!iY��x�
5�ȠO���
�"Or�
F
��|�dk��X�68I�"OҀ���.{���Dh��*m�8s""Oęҳņ���}�C�4w����"O���J\�M����3�J�$L�$��"O��@$ϊ�X�µcF�D�2����"O�y�taޏu� ҆k�@��"O�U�G�����gFݙ:��);�"O��J ��tOB���BZ�xHP"O�K�F�jళ���R��l��"O$�x�D�f�Z$��@ޝ"��T�7"O
�Sb��X�6�0��� �@a"O�y�2��\rn�%cƪU�ц=D��Ah�X�L�P��UB��M �o=D�(��	�Z�X�hT�-8N�%<D�\���W7 T���*�,�����	&D��q� �2	���Z #�7P�BM���8D�� ��;�ذz2�C^�� �1D�lk�תT�� RtU=��}{�0D��i�㍓R�BlYG� ��}V�.D�ܺ�ˋM��hq�D�G劵�7 7D�܋ �P$}�jtiG[�:X��9�h4D�,z�����@��1azD���@'D��7�Y\����F ք (;D��I�Dخz�! D.Cr)t�1T-D�q��Q+a����{�$Q�W�%D�tZ"���q`����#Z���@#D��X�H�$N3ԸKv�xJxl+#D��p0/A>5�y�#�/U�REK�-D���W�\td��D*��)��T��D0D��`�oV8|�`��Fo��	FG1D���EOZ�zța�W�����c9D����F0I�����M�p�xy8�%9D��@��� s��ԗ �TqHv�6D��{��\O�`Q�
��a��X{$�0D�@�D��}z*�A�Xg�#��,D��Ǖ#[bI�5bN*��ر��&D��T�
��|B�D˳aМPbL/D�@�R*P[fEI�j²����(D����3��S�F�8��Q tl%D�P(�e��u�\�J�慫v��B�A$D����D)]�.��Bؒ]_vU a!D�K"Y�s��t���֥5�XA��� D���)R�F,$C稕�&4n��ԇ,D���#��[���Ԁ2�4)�B%/D��SP�$!���Z%�ݧX&(9(u�+D���Î`��l��)$\�<ts�*&D����m�F��Bo � �IQ�9D�Г��1o��h0�	8+�bl5D�,bP��[(���E�,�ҵ4D�xIe�˺A8P�(J%�x� 1D�T1��T⤙z�CIH��:D����(�3�lX��H(�04cFg*D���Nơ 3|�`�F���90;D��@�U3m����Ţ��"��3D�Ț��8nC���mz^}Y��6D���@�vW�����OgR}���"D�8��& ���8
��;w(�Y���!D�|���i�f�ڰ�J�-�x���@=D��2V΂�HT h���	�&q�<D�� �8�T�F1d��%�p��9D��Ȅ"O��3�.�!f��t�K4p��ks"O�"C5%;�q7�Y�6G@���"OHpّK�!�P��@��9_av]A�"O����F�S����K��J �+�"O�A�P šE�nQ�b�3mJ��c"O0�SF倕)�eq�厩@`9��"Op�Y�Iœ2�؍.�<�Se"O����V1�����,�lT��x�"O�A��ܘX��͂$+�-�!�"OX��d6vXHdjui_%Sc��J&"O�AZVbZ.�~��͕�mOHd�"OΩ��, �
���g�3[>ҽ��"O<�
�A��awq���X3����"O�d�D��n��9��>��$�%"O�(���/z�\��5%�p@c�"O����[�U��iq
��C^�"Ot��&q�Da��"`��]�e"O���ǊG�g/�pIB�O-}($X"OX��+R���1 �I^@��0"O@e��މu��M�3ϔ0RDtPR"O6!�C¯G`BTG�1b@p26"O.h�ѡ*[���cg恪^x� �"Oh���z���Ò%ϧ�>��A"O�\���*!�[	~����"O�ȳ��9>2�rԠɒ&I^<!w"O�a�@��m� ���H>hud"O` �5��g�4���mA�l=P�r"Oڈ�v��QV��,��E3�e��"Oؠ:��G
cl|�1K�D&�t[V"O,�YE�@�y,@�g
#;:���"O |�"�<V�0M2��Q�f� �u"OP�E��%Z(�$ǋ�\gJM�%"OH�t"_�zL�����_!qN��X�"OB(��X>@]*$aP#�BjJuS�"O�E�tAJ��,���NO���"Of$c�����Hթ��� Y4���!"Oz��Mߘ��5ѷ�51��$"O�وCi��J�J!�t �,���3"O���I��KbMQa�J-���Y�"Od|�����%a��&)�&%h&"O�;�"ߏf��y��Gq� -��"Ovx�B'3�b��*z��IY#"O�D◁�9G\ e��%|z<��"O��i=�@��GG��A�s"O�	��iX�L�L�a1I	`[�={�"O(�Q`�S]FY��AVT��"O���X�� z�c�>O��"ORect��n�00W_�h@�i��"O�{w����L3��ŵt2\ `�"O�$��< �)Zt��6T"�"ON�����g���j���	Bf�`�"O��@`�N
1S�p�f�̘�"O�#����WT0�������s�"O����@[/��h�b2I8�-��"Op��F)�K��Jq��w�A@"O����J�$�8����U*��"O�<�fM�NK���w`\}��J#"O��Pdh܌]��p��,ʿU��q�"O�l��h��@��+�>�t)3�"O�E#eJ�fs�t�W+ߛZ�����"O^څ�V)/� �2�	R4Pv,P90"O�=���`UTmA��-i	l��"O
9{�̎6[�%�1K��6��Q"O� 2}��ʓV����Ԁ�u3�\�w"O��a�.�0�k��f�r� �"O��
��V �b��0d�| "O|[p�=����@�R�Dn|x�"O.p�%52���̍RZzpv"O �PB��Zg���F�? �pc"O��S"H�5Ą�ʷ�F/,B5kC"O|��R�R.�Fqh�%ܿ~Dl�6"OP1�޻*;���1F�X�Y�7"Oz�z�ի	��� lҵZ���P"O�U��oY� H�DX�˂(h�a"Ob,��AW�%�8Jt��10p�H5"O0ђ�5ne�����O%C�3�"O�h0 �]]���G&Ϳ^����"O�Բ+ݙPf µf�B���0�"O4�sd��@ξ�kG��P0�"O|lZ���-g,���UŌy8��"O|X��ˁ6���8�"��Ж"O0	 cea���A�?W���pu"OЍ��#)u�t�k���Yh"�"O�i�Q����28�'a��6)^\�7"O�@je��9O�$�'�h$�#'"O���!��.U��I������R�"O(e2�#�)V���שŨ�ZQ��"O��`�jA8�PB�)��K����"O^��s�ޘkL��#���K7���"O�L����	���Z�DG�M�d �"ON��WE��`��!a�j����#"O䐨w
N"1?�-��i �(�"O��ԥ5h��I�7r��L+F"Oڠh0d�z��R�$>C��"O����9*�xXsǔF��!!�Хm�	�bn�3P���+\�Nv!���)_l�*�N�H&"��Ƭ��;<!�d����XB�Q�B�L�1�W4V�!�~�tIG�_�Zڄ� [!+�!��<C;)�@5�@�!�� �Tɡ@CY<fց�e�0i�!� �Fp�0�UJ
[M�H&.W:H�!�$Mk����@��5K���$� 0�!��8F(xMw�0E��w�ں[�!��
�^��A��N�-%HI1`�J�x|!�DM�fL������$F
ȁi� ��ZB!�������C���ˡn�C�!�d
|n8�D�-������J�!�kgx���(�GD�bt�&)�!��X �8,�v�(��5ve!�D���@����s�dѲ��a�!򤂀b,��i���.�Z�犘` !�d�,J���0���^u�${��s!�$`z�ԋeile��
�4!��K]�T�)��U�q�8�
P�!�H�m�́�'�>}�؋�B�K!�$#DBm�A_�rĄI!��i!���	d��NL�dR��iW�.�!�Ĕ>�[�+B&ER��	�!򄙱=)�sUEYb����@�	�!�$��:�jX �)�ki8���L�!�	;���w����A��>&�!�$�Y�-��i
1n{�0W�N��!��($�ʜ�%��GE�ѡ3K�N�!�dC�S��Y6f	2=zhX�*G1P�!�D��T�q�kW|ؙ�)�=�!� r�1��`�UH�jW�	!m�!�� `89���5���A�7yB0	c�"O�d��?=&�"�C�LH�u�""O�=�C���&+$D�BfA-"����&"ORQ���	ÎL{��.9q�L��"O�̩���$vճ3Ŵ:"�ð"O�<ze�Q)w(٢��-դ�RB"O�p�C��~���4�,�V��"O&� �*��f��`�#�"����l��T��� �i5�?��`l �~8� ���ƾ?0�0J�O����ɄmV4M��&2J���aeG&+��9�e߂,$�˧��Ć�+#\���,��$�d&��Q�T�X/B���F�g�
�Ru�!xL�͟�Y�
ؿ/��u��W#:#�]	3�x"�A��?Y��iζ�4��AXSjW'v���o�3Ρ!W��O���D�}zt��5=��DB0N�Fc��v4�<�ûi�7�3�L�(���#��/5�u�@-��Jl
�4�?�,OV�HF��"=Q��Q�\���Y�+S
f�)S�����7��/���C�k�3k@��B�?��� P�PK�3��`�tD� !AR�R�ch�K!�}#1��l���f��4��p1lV�y"ɉ/��@%X�Gx	!��ļO�L�n �MC�T@J$@�S�gy·ivH-�삄J}F�(4�(�0eǲ<�	�u��h�d@e ��B�|���$�4nڢ�M�O>��'�ʫO����
�$�v`�Hp'�q31��/v�X
ڴ��<���&2���@�H�D\j�N��\��)��G�z��W�Ⱦt���&���.ߤ$��G�p�',t]����*.�*�Аc�=�R�)��צ@�,�a��9\�YN��"����W` �ʜBlCIȼ-���W�xa��`��˟��ܴ<��'#��'��Ou��'H�IȺ�i�i�@�<�)�"O��3��U�?�UzŇ�8Z���#�X{�I��M�e�i���|����4�?iݴ8o8p�*���j��Ǯ_����'���5 ��'^J�*tB�F˵m�^�;�CN?Lq�5�҃�j�"���-m���a�A�pJ��	���U�ĺx���9Y�h=@�a�s�4�qҭ�#qi\�
7Eҡ/�0Q�IS��ڼ+Ġ+�	�v���d���A�'�$\yՊ��38����e�(��'Mb�'��O�d�[�	W�숢(�g�UXE�O8�����S�C��s�8�P��N�3¤��3��,p��Z�+eL���M��䧦j�46�@��QeF�Z��3�kO�V�p��?��҄h27�6Ҕ%j��43U2�L�����{�na�G��B��A����({�'�6��A!�-f�Pl�0�Ӷ����!n���͟�iH�^��#�m��g�|Ik7�x"ۚ�?��i�"}Xwȉ���[-Y�$��Oln����'(���5��0�zA�&iV�a�4�1�Z�'��7-���&��9�!�:�̲�ř��@�B�L�]�v�'hr�'�L`�3�ߵDy�'Gr����6Jh~A+eG�+Ek���&O�D%��v �i=�7��Z���qU>���j	�X|��@�6f `�6Ȓ���y`�ѵk:��B`O�Z��!a$o�E9�F�.��q�\ኝw������C��$y&ė>l��8Be��秊{޴�?��/۽�?�}�'ڛvo�i�"�8�a5P�XI����!J� ���O�ʓ�?��,O<���̘~,�uA��[�6�	aW�>5�imR6�*��X����>��(�&a�	$��l��Ec?�	��[�
=`  @�?�   �  �  �  �  �+  =8  tC  DO  gZ  we  ?p  By  8�  ��  J�  ��  ��  A�  ��  ı  �  I�  ��  ��  F�  ��  �  X�  ��  ��   �  ��  w � %"  ) 28 tE N ]T �Z �` �a  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	���y�'H�5���T���B`�T�m^2���'Q8lI��ȵ�|,JwI+����'���0!JҶ~(��	k��W�4(	�'!���.���v͍|�BQ�	�'Y�0�W����M��\��x�'nуdE�du���>V����'����	��%ἘPu\P�p|���~���@ȵ�P� OC��鑪��y��
+YN1
��tL̝ pM�-�y��ޭ$L�0�uC߷kI0Q8��&�y��W	-�]��#a =�c�ۦ�y"o�t��"�4�
ԇ=�ybC��JTD��+J�\�ykrGN���D*�S�O{�L�W��4v\�`�L���I��� �Ȳ!@�;s�l�G�S+T��<O�00�@JAX� �V@�d�v����X� ���.4�O
扈;��X	�׋,t�Pb
%b�&C�IcEV�#�l�|�a1�� Vp �'Xa}o_�jL�%��ͦL+"�����p?!�ON��D��4F%�U�'�g����"OIr"LM�]$���X�3�lx��"O��`�Nޔ`����C^���}�"O�4 �'�@�8�b]<Rr�XRd"OL(1�ꒃN.ְ�2OH�V.�C "OB���/�i�P.��p�s"OΝ��f܍ �tC�
z�Y��"O�U�Ώ�ZvP�Fqd����"OL��EDU/$粘kwd�9D�0"OPYƤۨo�T�Wě�^3��"O��J%-¦N������9�jt��"O�]�4j)9+|	�eB0+]�zu"O�� #�v�P���I�,A@t%ے"O���cV��<���(_&A����"O�8g��W�ʑʐ�ܚw#Z�9��IҦ���� 6��� �^݈m�ABBu|�C䉖#ņ�j���7U�b���əh[��:�4��}��?�'A݊����^�)e�i�@�
�'5L�R�Ғ<*|z�(�"�r)*[����ɑ^0|5aV�6k�01 ��
YN��D�{�}�>�I���8(�Pb�]�^���r�0Ag.�	9f��E�(E���=9�O��~z4���	�rl�d��%�$bD�N�<!�gS)��v��?0GN�2��M�<�v�R�Q�T\@�%ļD�t���E�<��g��h�R�(�8bd��NC�<���\	�`·� �Y���Yѭ�u�'�ў�'#�.��6�Q�`C4��Ɩ]Bb]��D/�|Y��b�F�R�AI19B�y��Dx����	I���#(�3n�L�ȓ$���w%�=s	�Pc�*��T��	W<I3BIE����vȝ6O�N� F�x��&��sd-S��VC��4S��
B<D��hA!X�1�D���%0�s!�-D�tP'N��5!dU[����rz��%�,D�x�
�g.�q�ѭ��gl��â(D�X0��n߀����	�@HZeBB�(D�,�FCևf72E�WjƛhX5��z�����Nh �"#�"CQ6�;����;*�z��PM�-�j�afe��4w���� 6J�|%��-��yjp��`��SR��� �nڬ����%%Q�)�t%=�ܴ?��hҎP�\���e��Jn��ȓge�8AF�Y�Pj��^)�^�k2�$��(O��W#n�S�#&��ġ�^Z� u�ȓ*~�j�h�=2Nm����a��ѳ�<�S��yBT�Rˠ�PSiީ,����g9�O�=�Ox�i��c�N��ő�n%�0�O.��$�"u4��Bڂ7jz��,�5	��|r�xbD�?4i���CFVd��<@����y��,cE�f�A�M|��(��S���O�:�cQ�y�0RF�ʤnBq+V�z�<�b�8<�X���EQ�{�&Jz�<i��ӊ,�F��3]6��g�Ku�<�
��1r���Бj���s�<!ak��q_zy� �\���B�AJs�<q1��*԰��ↀ:Ny"�A�i[m�<9�ˀU��x�!��'���&�O�<1g�J;�
6+�&��Q��_c�<�e�Һ{洽�4�U=	
$�q̟T�<� &I��W�U�H�H$��M�4Z�"O,AÍ�}>�hP�B�P,D�a3"O��!H��'F@���DD�A� ��"O8uj�@�1�r� 󣈦m��c�"O�q)7*�$�ap��D�7���ʵ"O����^���,�ꑨ���"OLH�u-��]�2eA��5�B0��"O�0'W��d�YaMҬO��}��"O6�p�����@6�&yj��"O-Vb�8vp��	lǧI�"Ob��&*9.y�HL+ah�K3"O��X��ҥT���4�WR�(�"O��r�bКZ1ȍ��M��uUrl�3"O$����'������BU�
G"Of�2�$C}l�Y��ԿjD���"O@����ѵw�t��˔�p}y�"O�I91�ʹ\id��᭏�d����"O �E	�9�L4��L�" Β`:�"O�M�#%ͳ ��"�K:O��)�G"O.��3��UP�8����v�^�;�"O0�j����("ܘ��8߸\��"OȐE�_�	d�,���@�\�B�"O�D�׉ۺC�N�hQ���y�	�g"O��9��Z3G4���'E�=d���"OĬ�Q�ʒ|�B�HG����$ �U"OF5��c�:W
�i��I�Y�N��"OT���8e����5B�/$j��J�"O�����S{ș�d�\���c�"OXM�B��?�()�E���� 95"O�49�9g>�ps�R��"O��`�&B��b�8'2�L��"O ՛�L�	0P��h��A*hفd"OF��tC��%��� �;r����"O�	���T�ZM���H�{��PA�"O�YX��$�{��ՈF���^�!�Y�ꄃA�
��i����%2!��|�� Ҡ�H�5Lѻ��6x!�$λ�N�9�!�)@84a�bƜ�`i!�$5��B�V�w4D/iv��
�'�B�h�!B<�ܻ5L�;Y����'�N�:���YsU+T�dh�$b�'����cG4�t��L� \��  �'Ҳr��6n>p�0c��"�pH	�'bJ���$#��<���܁�d�[�'�6�;�)��~@��6��!�����'
D���P+[�\M���K  ���'f6�"o�����	�`�'D$�����3mS�3u�J�3� <��'��qXO�E�&��i\�(,v��
�'?:�i�G���RAq3G��k��I�
�'��D��WV����fփi;Ґ{�'�B9A�d�	j#& G�i����	�'w�-�'�3�$	z�l��p^�P��'4��a��^vV�ʒk�>��'�@@ ���Z�V�聨Á,] �'�FxP�JR4 7z����J�7�d��'�����H*Mn�X�e�V3��[�'\dY#���#J�`���$�\�����'7�AsĂ��8����A\�,�i
�'(сƥL!{�I0 �85�ld�	�'�+A�^��|�+Y�}���9	�'��$B�L�(b���[��͏zD����'VشK
�<����иw�^�J
�'|f����Y3�.cU�Xj���
��� �� �L,^Iɔ*��g$XA�"O����$F-�H��
�_(�90"O�(PDo&f�� �H�!D,�"OZ�P��P60 T�J2H%n�`y�e"O�T#���>,2.�0#�%������'|"�'}��'B��'q�'���'��򇢎�S}�PR!(R[%H��'{"�'���'S��'DR�'U2�'�pzDң� �yg�&0��`A�'�B�'���'�b�'���'Q��'��A�W�#8 ��*�v `��'MR�'}��'f�'7��'���'j����K!�v!��Ĉ?h HI"�'���',R�',R�'�"�'j��'������i��+�@׬�1Y��ߟ$������	П��	��I����I՟���B!Y^l�o��r�>�˕՟���������������	ԟx��ß���"6�*Lr�B�+h����ϟ���h�	͟�����]��Ο��I�q9���%Ւ��5���q����ϟ�������������	�8�	�� �(#�YL���QJ�?:�x�	˟����d�IƟ��	���՟P��D.�R�#_2*��С�j�~G�}������ӟ��	��|�����I؟T�	�Mgr�2�E�=���ɣ)��&�$$�I�	ٟ<�����	����	���ɬfI����m��`ak���L��	�����������D��蟜�4�?	��td	¯��n� (��m�9P��HR[���Iwy���O(�lZ��y��)��}��<2#Γ�Uqѫ<?	��i#�O��O^6M �칡���S���ȗ��h�Tl���dc�L�צ��'�ܐJQAH�h�\(�����T���(g:�)b���3�)���O�ʓ�h��̓��L�{V�H��ǝ��B�I�i���U�P�*�v��'^��w̽�6��C��T%_&eM¼���O�7`�엧�!g���޴�y��(��S9z��ƫ��yr��&�<}�#ǥn�ў�؟H�G+���=2�z�|���F|���'7�'MP6헹/t1O�`!���إ���=���p�-�I���$�OP7mo�\�'��Qg�Nn�}���)h��tC�O�0{�G� A���q���!B���ݫ�?�6�ͯr�2�c`�B5m��QER1��<Y�S��y�̈ ��)"�q��Ԡ�9�yb({�")��<Qڴ�������bF&@� _?�\��№�~"�'���']����i��I)Ǡ����5��z���#(�F�P��u��o��]y�O���'ZB�'�2�|(|d�Lت5�ɸ�m��m=�	��M���B,�?���?I�'��I�O�
�lB{�΍�f:� ����f}rf{��@o��?�L|���B �C7,�*�
7M>"�0�� ͙8Eܐ2��L���D4+�&EQ�Mr�UO>�,O0�(2 �'3��E��b��D?���P��O>���O��d�O�i�<!�i�����'UF@��)L�If����&�I�A�'��6�,�I����]Ԧ%��4*!���N��B�Æ�n�${0�]7���t�i/��OR�+ǧB�7���� �<��'F�k��<z��!��k˯t�~�cD�к.����O����O0���O��$-�3I�H=@�XUTЃ�*YMo�!�	ßx�I��MK�)�w���sӨ�OX]e뗵Q���8����;�A(��U՟\�'/n6�ʦ9�ӀT.�]n��<Y��YWp���'IV:9�ph�W�(�ѷ$�,V�3�ǝ��䓭���O����O �d0�ֵ(�.�K��#g�<۸��OJʓ�F���d�b�'�BR>��gŐ�����/��BE9?��U��j۴+�&$�O���)z��"\Amf��M�.-X�$��	����ЂÝ�N��F�I�Z�8@��6*,�0�����ן@�	����Iǟb>��'=P7�Z'��#�.��r� E�o���Ha���s۴��'���?1�vO�L9�g�>r4�`�A�h3�7m���z ����̓�?����"~&���c ����G�*��D�+}y ���m[
���<���?Q��?���?q/��!�V�01"�{b�+_����J[����F�t�	֟�'?y���Mϻ~K�Y���K�U�Տ�C�,L�շi��6�r�m}�O��D�Oe�p�2�i����4}d�q&� ����V"^� ��+�:����X%�O<˓�?y�t����2#0\���O��~����?���?*O�Ml�,)=���џ��	=?���p�L�\��1�'.D��?�7W��ܴ)����O����-�wa_�N뢽��B�� �����?��.9D�D����ԥ����34�v�]���2���CY��lӦ�Y�D�����?����?���h�2�ę�/W\��ʜv�&��V�\S��D��ِ��ey�w�P���C�0�W>�H�ŀ
NӸ��M�B�ij7-Q*27d�d�I�Z���Kt/�Uw�8g�t�*'i�Z�nkb�GJ��ly��'"�'�R�'	򤖩H�f�˰@�����Ae��Ɋ�Ms�f�J~r�'�h�ę:�8�a9&��ӵL}yB�'z���O�������tU�Ƽ V�y�@C?e��9�A˿*W�ݣ'�<ɗ�V�o��h^wq��O��P��)SA�H7^tZ��]J���?)���?y��|�+O��mڟ.���w�&YZ�-�p�j�hCgD�"���	<�M+����Ok�I��M+ӷi"�7M���r䂱-�|�|)�"E�Ұ���t����/�"l[$�X�wj��4d[�<��E����_� ���@�V�J ������;lq��<Oj���O`���Oj���O �?U{��U��p�I$�3z��2�E��h��ڟ�K�4?Fr�̧�?i`�i��W�<�a��\��}�s�Z4�I�CE�3�?��On��M��	S�Iڴ�y"�'�D�P��T#��@�^d�t��7. /�8h�vÝdG�'��џ@�	���	�c�B�Rv��P2�F�ܱY,�I�4�'�\7m�1N�Z���O�������I�T�Th�U$C�x���yf������������= ۴r����OLΕ�Q��w3N]��G&m��<ʰ�\��wh�B��	�?р���+��|r��J:�Ȫ��77t��c����'��'d���R���ش'q*��@b��ta� �@nҁ@xgV���d���?�@^�<(ڴWh�
V4C,<kBCq��S��i��6�ϥ4��7Md���ɷ;�̳"CVk
��'�`3ō�H)�D`Fb�+N�̀�'P�Iɟ4���L�Iߟ���F�$�^�TD���1o]�2��+ዋ�cR�7�LZ#��On��.�9O��mz�m����	��(�O��m�41����M�D�i�D�>ͧ�Z��1&N���4�y�@_����_37��=�c��9�y2�J4Mo��H��<�'m��������v�P���VJ�d���Y�`L��	ȟL�I����'  7m%k4�d�O�Ċ�?�ii�@ƾz �6���:Ш�d8�D\r}2 l��oZ�?A�O�Y�^�����

��2s�·�y��'��2�e� <���e\�l���W&���;Y��E���S�Jgz�Ѯ����'%��'��s�u�ƭ˯y�vX�&�7 20���I՟lrߴ3��%����?�Q�i�b�|�w����R/�hU�{�K_�v��{�'u$7MX����ߴdq> �ڴ�yR�'����n
6��q���Y��X5[GB�r��U0�A�l&�'���ɟ���ӟt�I��������Ie��!�m��0�Y�':�6m�0$����O���4��<�dQ�7����R��e��D牆�V`���M[��i�8�$,���F��p��E��6��Ѭ�� `�3�(G�N����h�<y�ϓ&P�r�r_w�4�OD�Х'��T���5��J�y�h��H�	П�����Iy� qӮ`Շ�O,x��f�<�k�ƩG���I��Of�m�g��n\��5�M��i86F.s2hMxa�_$Ɔm_�|�F�k�"��ʟ� ��*V����by��O3p���lX1��9+j]j��I0�x��՟���� �IޟX��m�'�b�sP��1������Hdf͓�?Q�X�� �������&��jE^%=�i���� u6R��!�*�?٩OD�o���M#�'9STl�ٴ�y"�'��g�ȉQ��Zp�AdZ0�T�HBB�S%���'A���4�	ß��I�b�̄�d�:Be�k6Ҕ*�8��	�Ė's�6ͩhw�d�O����|�u���>�h�*˰z�`��7cJg~2$�<����M���'��O���$���jc!��^?��� )�Nr����K%�z|��Q�(���(1>h�;M>�'����hZ�]�
��eޕ�%cE�?)��?���?�|�+Ov,mZ�iȰ�PebJ5t��(Toөgh����[ɟ\�I�M3�r��>	 �ic���3V�/����˙
s�r���!{�D�n�3�6�mZ�<����4aB�@ UⲘk,Obqy���4Qc �Bg�B�P�8]��6O˓�?���?Y���?����򉖟?Bırf�%MS|����-X(�m�46d�<�'(���I��]6<���'-u��t�7�V�t�n���4+�V�O���|��'�1��6�M��'��i@'���.Q�H`B �F��y�'�Xz��:2\jt�|�\�X�I��xTg�%:��0G	[g��aRE�̟x����IQy��jӦ����O��D�O���	�Y8�Z��@��/2���̘�O��m�'�M�#�'����?|v�Ѧύ�����ʎJ�"�I۟�!pG��<B�x�5ʆby��Owژ����l��$y���M�H���n�$!������x������i�O��F�&���;�N�(F��g�Y3\g�ki�x�)�(�O�$@Ѧ��IO�i�M��BF�ul84���P�E،�q�"o����4���!q�v0Sc%t�*�I˟I�
�}�E
�~��A�D�h8� %|V��$�(�'$�'
r�'G��'on46H�91���s��(t�d�$R���۴s�
A����?Y��2.�H�$�h��01H
+u� PC �E+���'�27P�����ħ�J�'r0�t�ۊx{
����_�K>�y�Њ�!{\1�/O� �LP.`{������D�>��2�K�%x�gk��l �d�Oz��O��4�z�4�FB�?^��p=����6 ��!�E��y��r�p⟘íOx�mZ�M��i� �
�E���� FƖ����C:��:OL�ܲ�
�a�0ʓ�� ��ҁ�1DPh<�I��İ3^�M�u>OV���O���O|�D�O��?�r� H����d�-�ܻ1��ꟼ����PZشc7�A�O��6�2�Ā�N�Z��4X�(¬�iR��$�P��XyR�isv6���(��m���	ןd�P�ӺY�$0�g�R	 ��0��L�� ��9���o5(�$���'-B�'y��'��@r.�.��97
T���8��'��_��j۴AEl!i���?Y����)ׯ-=���b$�\z�O�'0�Ɍ��D���YܴC����d�O�J��q��#e�0�bA�$Ir �;��������8�I�?��4.�꺃s�|�[��:Ƭ��:L��Ԅ�D�b�'���'���S���4'�R#W�~�x�v�ٜ
�JX��.�!��$�A�?�vZ���޴#S�U�v!_�TE����?�Fx��i�*6�H<�7mi�����
	씸��KV�ܕ�� Ę��_2\��)�$X?
����R<O���?I��?��?����)��(iy����97F���@ω9�l6<2�Iȟ��	I�s�P@�����J�	\��b�m�?`�J(p�cW�ZY�6mk�Nd�Im}�O)���O����¹i>�D�#,�I��M� �ò	Ba��<�Z��ŉ½���O^ʓ�?	�S�`0��E�?�ʥAT,�'�j����?Q���?�+O�m�8K�޼��ޟh�ɾxmPM�qo��k5�<��mO�e*,���t��"��D����
�4gVR^�|+v-O(|���t��"�X�d&k���	�N~@��AB�[�\�'���dď7e�Ώ���Ko��Z0�];����M�lPʵ����	� ���@G��'Fh��5�V%��u�g��!e��T@��'�P7��=�d�$�OPln����$�杤{�u[kʯR%��Jw�B����I��M#��i��7Z�"��6�|�|���u?
ؓ�*��mi�	�aLϲyv<��C��	ZT��G
�r�	Py��'�R�'e"�'��!B� �~���E�MR@�x$�.�	6�MS �A"�?a���?�O~z�&���P(��>L$����	Uu^�����z���'�z�'K�VX��ʔ>ެ�P��	;>0 ��ݔ@NЩ+O���@�ȯe.*��䓢�$K7;v^@uLV/;�X�Ȗσ#|��d�O8���O`�4��W%�ƌB��y�ԉoeHU��(+G�T]Æ@���y"`q�㟰!�OJ�n��M�2�i�@����ˉI��pU���fD��nմt�F;O>��ތ 4V����9��˓�z���9Z�n�>Px4l�!�+3	h�c8O���O�D�OR���O��?I�Cf˂~�<K�D_&&a��x�<�����ڴ~�&]�'�L6-�O�˓Y��`��W0>�2=[w�]�
7� ��'?�ɂ�M���i���爝U˛�>O��� ������L.v�t9��R�\�B���
����ʥO3�d�<����?���?vn[�w�D�qg-�V�T�Po�#�?a�������"��m���	�\���?�2��Y90�ؔ��j2�q�@-?Y�U��aڴh˛�n�O������<EG�����9�x�zQ
��Ƥڝ:�$�I���<���({���\w�Ob�8!D�C��u`]?��er���O�$�O��d�O1�Z˓?�f�Y9�������O�`�Y���.[
\��O\}n�J�`���"�M�r�� s�x���U�9����O�O���n�"���u������X�㢊�x����@yb��2adF�f�f>�Aq-G�ybV������ ��џ ��ǟd�O�dp�6����q �N�~�`�a��e��@�"��O����O\�?������6���xmH���d��Qʧ�Oj7b�i�$�<���?���(� �l��<Qk��Cv��臦U@��!���<�d'�}�6���N�����D�O��$NN�}r��7
��E�ƀW�C����O>���O˓zB�věx���'KÓi�h�c"O�k�0DIpN�fu�OU�'� 6M�Ϧ)�����Ыp���1d��8DX��PTq���O��ADMZ�G���f��<���%-VYK[wV
�D�V�.��ꛁU��e�KI�5>���O��d�O��D"�缣b���F�jPD�3w���1�
�?QU�i��@��';�#u�Z���_�e��b�z��;���I�M[��i�7��'8�D7�{�0�	p��)���,��8��#)B��(@�$S,�\k���H�dy"�'��'���'!�Y>���eK�8�|
#B��P^���M�$��?���?�J~��1�`(�uI#y&fD�P-@�>�a�[�H�ش|��O~�b���|�j��C�%r���+:�tIb`医Oju�Q��<)%��v�	]wU��O��X�8��" r4X�e\X����?!���?���|�.O m�+.����	<%4�2��B>`��� �0y]ظ�I��MC�rʬ>iT�i�7�ަI�Ud]�] .�p@B�N�H5begM�xmm�<���i���I�*��x��\�)O��	��sQ��(|�^@�cE�24�� b�I�<���?����?���?q������m�0����Wٖ�Sa�
�"�'���z�z�s61�����ʦ�'���m_*b�3!Ȗ'_��:��?��O|nZ-�Mk�� ��ڴ�y��'ez!I��A�X�̐r3�<P�"� 4�O�y�6`vN�57J�'���ҟ��I�� ��/lI��P0�C��p&���8��	�'w�6-�7N�D�Od��|"��O$�,�z��l�c�s~��>aаiD7-���<$>��Ӑ+m�bc�72����i�$'�����i�I:(@�iLMy��O���P��J\����5Qr�)'C�:q��B�� ������E����.*q��yA�Z�uT±��A
��s$G��-hTu���qv| B��/ '���b�7u8�zq��3ih��3���7����L�XS���%0�A��@
#c��L6mn��#O9b��x�N�5�V�h%j�^n�d��L��|��t�C�W�X�^�A�J3N�\k�E���E)�l�bx�B��P�>R\���n�"/�~-�/�wt�HbFS�	��R�oէO��������=���;��ǰC}�i���J�u{�5s���@f��� Ϸd?�@O<��?�H>���?A�h�*Q.�\����V]�L؆i�*�'����'���'���'��%�7�Ŋ"M��(��I�~�<P�4Ȋ�7��6-�O>�$�O&�O<��OD�K4L+j��Ve��f�r�Aӭ��	��r��M���d�O�d�OX�d�O@�F�Ov�$���x"Õ!h�� r��6��4{��cӦ�#��O���n	��#��x�%��7g�0h���)�.(r�B�MK��?���?�T��?i���?	��r��$�K��_"���#�'B�'k,�Vl��������$o��,Bƪ6\ClAХ���%���'�2�˪ ���'����?͖�5�H�&�2�Aʇ���bwĻ�Mk��?i,C?P}�<�~� 8����Bo\]*�*�,r 9��i�ZD[��'�R������IIyB �$H�~�H�oT�~u��A 2�^7MU�@9p�'��S��,��H�}��G�ċCi�u�0cؽ�MC���?a��P
\H+���?)(������\ aIV��^��ϭ3��b ��'B����1�I�O��d�O.�*dgY�hw�q��bD�d�jq���ަ!�	/p,3N<ͧ�?I���DYw��� ����(�����P;7wymZ��\��N0������ğ�'�x�Q�[�$F�(�un�$;af��&�}�O����O���<���?	�d "V�z!�#¡#�@�	�Q�kD��<Q���?����
T�~ͧUU(����%80|H��M v[��'w��'o"X���	֟��SM�~��n�8 �X}[�FD_x��}r�'lb�'y�I�^.�(sK|�"Θ L���X��gIF�BP��+���'I�\�X�	���I��#�SqU4HJ��Z9���L
�6��O���<���¼^�O����5�MY�\u2�ؖc��fA�OH��MC*O��$�O�e0���柛F$B�q����`��J�Mc+O,@q�������D�D쟺��'�"�b�(RL��L(������s�4�򄓔Y��)�H~n0_^B�@��J �J�̓�}�h6�0`Ըlݟd�I���������|�J �_9��B�\�]2�CQ �ƛ�a҅oI�Iʟ��I�?c��ɠ���ӂɀ�l=�D���S�O4��Jܴ�?���?��/B�-����D�'Y�MK��H}	Ì��V���#h��h���?�� �0��<���?q�m�� &�wX�"�Ă]���ؕ�i��iO�S,�O�I�O^�O���g[�TR�����Y�qM�U}Gė��'�B�'��X����	̵[v�8��Nȃ�5Jv	����M<I���?������O���F�nܰ��t�D0t�K��/�le����O<��O�˓M�
x�=��dñI�&0���/�$����U������'9�s�xw��~J@�P:fy���ǘ9�rD1D V}r�'�R�'�ID7Ը(O|"���C�`��C���FX�"�"'<�v�'q�'O��6Q�c?�{E˖�.ddBڴ�j xjb�����ONʓ_q��˕����'��\cPP��#d��jH�ٶb���z� �O��Į<Ib�V�O2�	9q��i@��K�t�Ȁ�t�޿K��6^���$��M��X?%���?�:�O��k�NG%u��͙�i�<z�ǽi��*O��S���ܴw��Vm\�����@O�D�ґl�$爵0�4�?���?9��b���tB�+w<�_�Nwfa�ì�0t�E�ӻi�� K�O�˓���<���
ڪ�B`"h�l�q��T�l���i^�'��J0vIzO��O��ɒ1X\Ar��3�pR �J�D���$F<91O8�$�O��I3����a��PD�D�A'��!�z7��O�����<����?�����'�����!iQ�,�4��:Y�	��O���"��v+�	ʟh�	xy2�'K�I�&�߶��L,�>�'-��	~�IꟐ��쟸�?���y䐈W'k"�=�f�Na.�)c��~ގ��'�R�'��I��D[4cY�v��;��q�kR\����IǦ��I՟���p�����8țv!�~�����W�F,�)��$�O��$�<���+Px�+�"��+g�件��G���$A��d}�Hl�ϟ��?�)O~qAӞx���dx7��:��LJFj��M3���D�O*�cw��|��?	�'Bv�2�J�Q������2S��9q����O�T2 (ە*�1O�S�c�@AХ/V��U� h�)Y���?12'�?����?I��j-O��Z�dl��fm�����bj�&L��	��qvo�,\�b�b?����A*
T���7�xu�%�t�*@�U��O��$�O��$���|����{@��xR隖��7}x�:UJ��M�ʳ",,��<E���'D�I�׊��]�<�{���H`PQ5){��d�O���#���|B���?��'�� �a �i�="�bɫx&�)se0�-��u�L|��?�'66�K�38�1+�/^�%w��ܴ�?�M���D�Ol�d�O�㞨1U	|��	�a�%F��st��>q��[�|1n��'���'���$�d�$_���a)��Č��e�Q	�'���'?���O�=�tȏiF �iE�3�H��"Ι$m�k��$�	៘�'*���y��i�R\�`� 8������#���'�'��O ��ƝPFp����i�r���B�C�~��������O,�d�O�ʓ�?�Ӧ���)�O�;�	�"i�
<�b\+T@d��t*Aզ��IE��?�B�R��&��;���L�*)�0㔮1K���Mi�z���<Q��\���-�t�D�O*�)V1� � ��;�������0C�j��>!���z��_c�S�T�H�J���#����]��0�O
�d	�N����O����O���<�;MT�z�aC�(n�qt�����'"�>Xj~���y����	=/��t�웖@�Txe@�;�M�D˛�?����?9���*,O���O�y��J<H<\*$RLl\B �ܦE�#?4Z|c�"|��C��wm@G����D�!�]��i�r�'���8#�i>a��ßL�S'd�㕨�9~�.M7�#s��ɂ��8B&>��I��L�S�?  ū2
j�]Q��#$����e�iV��F=#{���P�I����=� j� r=xЉ����¨]Byrحm�%�'gr�'��	�����k\���xp��'4��*B�����'�"�'u���O�-3�
(�`�3bĆ2("y��D��89Tz�����	˟x�'"R&�+.�i͗s,ht��;?L�V�K�ԛf�'���'��O<�d�Q����i��i�O�3D��dβR<�h�O��d�O�˓�?$$����O<i2��D����E@>7̤y�4l����]���?�Ոڌ~"�$��B6B��
��r�X���A*V�a����O��;�6e���?Q��?���2v���*[�q����P�
�zE����O����B1O�	_�Q	4�t&ОS8����L5d����'��'IE=b�'2�'S��R��]'A��� �À;/�yi�����?� &֔[N��<�~J���H>\��b�gxfAS�m����*5�Eߟ ���D���?����$�'K�գ��)���)t��#Z�BypCӀ9�!�.Az1O>��ɰ#J։a�F�gD�u���C W�t�)�4�?���?���
��4�8���O���;w|T
�셷7�&m���a�(E��ybH�QX������O8��9����f	%���)M�pl�6�O��E�<)��?��Ѹ'G��B��B�aVF\��O�%�p��W����O$���Ot���<�'
U�(�ta)E���4Ωqg���! *Op���O��*�Iޟh��F�;C�t�׋?5���V�V���B��4?	��?�/O��$�X������t*F�ޤ����26�FI)s�i�r�'�����O$ѠG�dٛ�#و3ꜽs&�S,l��*�LM��$�O��<��� 4�-����l�D�� o4DS@�y&|}m�ПL�?��1�tm�碞�I?5�z1����2bgf1ɴ�Ѷd_�6��O���?)��ݞ����O��$�X�".�=z��RO��L�(��P��?��@.+���<�OѮ��4!��s�^�!tϒ(��)��O��׶r��D�O����OV���<�;O�z�2&O�dr�A�Q#��t��m�'y�[v�X��y����0"e*,��*' ��xA�.�M˰��?����?�����)O�i�O��!&P"P���5R�/� �N�O���,� &<1O>1�ɫD�l�� �"XKGO��p��iAٴ�?����?��^���4�����O����-���W�"�ұ��Y�`"U#�y�-�<:���2���O����~�����1�X��� �{{h7��O���b�<����?�����'B0��D� ;�Dl"��f�P���O�$a0�� �I�����Ly��'3�u �(%�\�T�B�e���'փj��	㟰��Ɵ��?���SXYа	9MlvTc����~�GLÙr�nm�'b�'���'�"��=�7�!P+�5�_��1�����wڴH��i	r�'���'�b_���	�e���s���ML6rTQ�% �w�xy�u�i9��'���'���'��*�%`���$�O`@�r'Vj�DG	ƻ�%�Vh��6�O��$�Odʓ�?13��|����~�k�!}fAHA�^�kpZ9s��A��M����?����?�R�� @��'B�'���oHO=�aZ7)L:?dmr�GU��6��O�ʓ�?� ���|z����4�����&.qdų�DA�K��Y�����M�,O@I��/�]�����	�?���O�.�; "�ɇ��
�VU#�0}7�f�'�2 ��y��'t��Aܧ0�� C�ё���wɃ9�N�lZ&s
e!ڴ�?���?)��PG��GyB�F�M2Ё���V�z�3�욓 �7�P0Rs������8�Q�$��<-Nr�cՠ?z7i
õi�"�'��LƥE�����$�O��J�� ��Ρ/�̝1M (8�6��O��$GL�Щ��6O���?��	ݟ<���R�x��(�����m͢�xp��M�;�:\Q�]���'�_���i��+���z/Jt����<Q��B��>�F��R~��'3��'��X�4W��M�jE[�k
�?�iЀ�<�(�ʬO�˓�?)-O��d�O��$�e�P��@'&;a@-yd�AE��1�����I�x�	� ���`��J/�MK5��I�̽��O �C�A�cE�0��F�'��'b�'��Iԟ(�$�>MztA�^��*A�c��!�S�M���b�������?�Y?�25�\�M#��?�!BQ�lJ�8p��� �nE3��K	+ᛆ�'���'9�I�$�5�z>���U?)u�E�Ww `�B'�$$����΂�����ȟ �	ߟ�g�N1�M��?������ԔQ|�M�E%�,Y(<�e�C�?�����O���12����<��5ʀ��}�EZ���	J��)�7/zӲ���O�ȣQ����Y�Iԟ����?������"D#�*�v�hT��Ae<H"M����D�O@���b�O<���O���51�&�O�}yӦ��(2z��B�>��4j���#�i��'=b�O����''B�'gބ� �h����p�O'����~�f����O��Ļ<ͧ��'�?��GZ	,�(�Y�KR�]e��)&/1Q���'2�'���K�Ij�����Ot��O���^���U33t��w�ɗ!�d��i�rV��ض,u���?i����T��OX�0��	MO��8Q���M��h`P���i'��'�'�2��~��19$�1ਔ�|&R����9�M�1�X�k��<���������O����O4%Xe��%��逧�7	� �#��4\�Qn�ӟ���џ��	5����<����E*���(~9#,��{T��A�A g~�'��'2U�� 0����� ,��E
� sà��Ջ�-=�����i�������'�r�'�b���yҋTX��ʂ����	6 ��1\6-�O����Oj���<��D�;��S՟�X,~����hr�x��+p��7��O�˓�?���?)��Lb~��M��)Q����c�i�~L8B"������ڟh�'��!pơ~���?A��L �a��i�$ XU���P�B/q��������şx�2�n�D�	jyޟ����\��FUط��3�D�¿i��H(��ٴ1���ßx�Ӗ��DE)���8��-�za*�+7�6�'FB�č�y��|��)�:�D�I���BK�*˂9ϛ���+:i�7M�O8���O<�)Rw�ܟ�yEFW�z��	�
�$�N�9E�.�Mc�kȆ�?))Or�D���'����P�	< ��+� \�C~H��Le��$�O��)O�j�$�<��។���D�q�M�{cVd�
�9X�x�lI�ɛWC��2I|r���?i��y���e�8k�	�Q̏�2r�,@��i�R^�	Ōc���	u�i�Ac��U�J�q�������R�>ٰ���<�.O��d�O�d�<Yp/[�o\!�7@�б��培d���ǖx��'�|��'��)	�+�@�r.^y��`�?:?h�'��	Ɵ��	����'��+s�v>��+
:�R��`��J��݇�ē�?i/Or�D�O���'t��dWL�taA�K�9����h��2��}�'r�'!_�<r�����'^XD�BՊ���$2v'�&v��pP���?yH>Y��?����<iO�p�-H�t� �'��Q�25���c�&���O��?W��!����'��,�o�An&�(X2���O����O��
�
 ��~z�� k������3�����Ք'%�̑��g�j��O[�O�x�{���@�'�������3�$o�����I� ��IW�)��cH���ǆ�4���
���q��6-^�Pih�lZ����	����'dH� �N��>�
��$9E�C�c��'!�OВO �?M�ɥ;���g@³q�0	@�S�K�Ⱥش�?q���?���K%�'��'Z���Ah��{$�'T9t�!t#��*c�Ob����*���O2�D�O���(�u q��Ɛ�Fi@�т�ئ��	�?j��	H<����?y+OR���l���)B#XҊ���dG��
�U���#k�p��h���� �'��e�ኖ;)[F�QTf�>o� ���E�3Vnc����Q�����ɴf��\x'��'`@i)$��;���(u-g��'V��'%�W�0��.I5��4�H�f=��j�QG�� ������Or�=���P�*���͈�� ��	Y��-�vhG��(�"�ib�'���'T�ɇL�4� L|�1_�h��0" ���E� ʕ~��lZ]�'t�t���'���ձm�V0dJ
vq겂W�7��'hRQ��˱�ڌ��'�?����r
B={�L�{��ӄB+^Mp� M��?��M_"�?A����T?��tlݤZ���6~��x��Epӌ˓ٜ��ѵi맋?)�'h^���O2܉�����r!�%�ʣ9�<�����OJ����h�KK�t^�p;��E7ZGz���i�JA��'?�'���O���'��S\����噴h$�$�'-�0�Sܴ$B^�j�b�g�S�O� �Y��,���רkҦ�Є�!Jg6��Oz��O<�T�C�i>����XCC`ş*&T�橇�r�̰p�L���'���y��'��'~f��kم����4,�(Y��H��>ɑԣ��<�����]�R���ʜ�+�����9[n~��SX��q��;Y�0��?A���?�-O�*$l�=Jo�� ��é���HK��M���'�l��Ο�%�h��ΟXXᬍ.,�@8�3U�~�p8��+I�
�b�8��ӟ���cy"zs�'S�lѠ&��s�T��eC7;�T�'Z��'�'[��'ݤ���O�ᐄ�0�1��;�ޕ^�x��矄��hy"��_Z�>$�r%�+cφM���J�k����cH�ߦ!��t���$�	�I�|b�xb�;�H4ءo��x����l�����O�˓^i uB5��4�'��R0�2҇� ��	0lSp��O �D�O\����~:ag� -��dX�����d��ܦ	�'����5�~�B��O��Ok��5���赉�8��Ň�,�P�oZ��T�I�t3r"<�~��,E3����#-O�.�\e��N��U �b�'�M+���?����:�x��'h�!�Dl)�|�u"�B�!Ythn�:(���)§�?�g╆(���i��L��z��hP�H���'L��'� u ��O��$���jǮܟ*��i��J�5ݮ]��(�	�9�Bc����矀�I�rD���"�oH�zw+ư.B��Zٴ�?AfMA�(�'���'Aɧ5�jϊ~�R�km,{�E�B��,����|1O��D�O\��<�B��'�( uh��8�	gJ
�LD)���x2�'�b�|"�'�®כC�PlS���4.�q�C�ME5T��yB�'��'��	3?6u;�O��#C��$�X���..�n�	�O����OP�O����Ot`1U�p�훵n�f�
0C��hz0�q�>9���?	���d��R��&>u�VB]*��IP`(	�O7�t*cܒ�MC����?I��2��P�>q�*��>�@����$A(th�7(T�u��ڟ�'�@����3�)�O�)�g�? �T�`g�NLi��h�$yy8��x��'��Ҍ�O���*ܬ�!�P�G��$��F�6�P6m�<1$�ʻ[y�F�~���z����2�@�-@�r$8T��=,���Px��$�Op� S�)��v�H@ad�Pd�`�N�U]�6�U'��mџ���ן�������?�F⃃k�z5��:����ck�lJ�fG��O>a�I�k�84�D*�(^>MAq���Ϥ�Mc���?��^YZ�x"�'i��OZ�1��ho��H�
�+��t��đ=>i1OR���O&��P�/(x!�ↀ(�`�C��7R^�l�ş�X�2�ē�?Q�����p�?+`D�K�hlЬ��A_I}"e����'�"�'~�V�p�W!�犛��h��qᤉ�;T,�s�+��O���.�$�O��DW�����,�!T���B�C�Yw�x�0���O��O ���O�:�'�O�Xq���O�T��F�Ilxxy�GĦ!���8��G��<��$x(�T�)�@a�:XPzUQ�g��Cx�'��'
��'���^� ���'8�HѢ[��<�b�F�Y��ct�-'U�7M�O̒O��d�O���Ô�s�'����A��ctt �#V�~T�4�?����$� D
��O��'���l�}�Zl)��BL6������7�1�	�#��)�?������5N0�4JM�$�*׋�����I����#�ß�Iȟp���?q��5E�'�䙘w��[`��ID,�
�M���?	&�Fvv8�<�~2w�/�]7(��bU�h�P/Φ�S���M��?���rt]��'+|��q�ܑ��4`�I�"-~�֠d��ȅ3O(���O�i��&���?Q0wOA�q
�H�rm$U���*Ԍ���Ms���?������cW�H�'nR�O�Z�A�,_$y�W'27��y��i.�'ڂ������"LB���ĂzѰ��r��))�FT{r��3\e�Ժ�D�-H�)��o��|��h[�O��8w��J$l+ա6\O8��
�ZQ�E��j DarA�[�V�� 0��Wh]Z��+���4���P��Ԡ8�2��^�B�t|����"��B�19&���cND�.H���T�I�:8��ܠ[����hĮ8����.A�D�aZEaKP�4 
�L�f����Gb��h�T%��臂e= ���d�,X���� �'���M�|\2�'���M�_p��&���~�j!�0�X(��Q��D=-�Zq��Acz����qӈ=�D�ɇz@�	�ՉP&�L����8<6��ٟ����k�,[df��#���� =ʓAЍ�I��'���se��;��cb�.����yb�'~x �f�5+�&$��zѰ�eC@<	4�i� �?�
�¡�ϡa��(���'�I�X�2�"��|����	݆$�dG�`�8��&B�pEJ�K�E8Hl���O�tCI�|���$KR��4��|�)�6ѱr�߿D���#50�\��A�>�G�\�a2a=3�����I
 ���#c�D4M�P�5OB�fL�k�|5����M�@��?�`dϊrj��1(=*��x�Quh<	�C���d a�)>��ĀX�H{��$P�W��̩��	�-�k��M9nZݟ�����SCJ� �ڕ�I͟����rXw���X�D!}\@�+�/�mP
�dI��qu���$��O"�p�C� Q�1��'B��3��[(M_j��ː�?� (�Ղ�2g�~5�CʝJ�D���2�q��E[�]�l 懝/�DQ��b�	q��1&�Mʟ0�'�l-(��|��D�3g`.L*�-����ݹ�@�
d!�dĖj��:�⛓T��˧��|�	��HO���Oj�$����O�W�9�楖�m8ap*�s:!����?���?���\���O��<3��l��L;K��4��ܐV�p�Je� �gZ,����i��hu�'$@�H���Ot�PE�����|x#fPd��'A��ez�|J��_8�@�qFL�@��T���W�o�l��#������O�=y��,^�a����$g��Z��yb@�9��h�͔�+# ��$�+��'��7��O>����`V_�X�I� ��-��[>en�	�҅ 	�P��Ɵ�pVA�۟h�	�|ʂ��S|�$�GL "&?z�F���x8|���4Ox�RU�0��'Ij�xW&J%
C��7�;�8m;�(�(��I��H�Iӟ$�!iKu�< x�O�JI�b�dMPyR�'��O>�wAO�'�RiQf:u����,�(��4&�,5H%�[�B�bt�X�f�����򄁦nw��o�ҟ��	f�t�M~A�4	����fƴP#��:ק�9xm��'{�Ȋ6"��c�#%�B/�:Xa��~�+��ћ�
�	j ��H�k(�1��>Y������a��A]��w�r���%?!P�mZ/���uᎢ^nꕀ7}��?q������'�x�#BΔw�<sE?+�2��<)����<����X�%#�KK�v��;.f�8ي�D�ht)��F�4u�p�s���!i�Yl����	�dJ����ij����ٟ`�I���C�hT�>c��%���Vbh�'�p�LY
�4$Ӧ �!"���g�<��ˣ%>^��,�EDʵ�Zȹ`��))b��m�\A.�Tܧ:|9Q�O�dxS�K;V�X"��
�Rh��ƦY�/ORȸF����?����?� �`�&dZ3|�� ���h'�� �,�O^1��=O���v�WsQ�k"���E	���F�� ��4.��V�|��O��T[��Ȗ̅��dU���H�x��kp��I���җ�W����I�����u�'���'b�ы`À�?I���� ��1Pƨ���7Q��b�צyn�R�� <O@+�Čam
H��ހ�t���K�;�pi�Ċ�I�4�I�l��� ( �/���Z�h�)U�B'�6H�^�p��O��di��ݟ,��b�F��}��a�h{Pn�~e>(Gx"�'�vMW/�:3�&��F�ԇX��'�D6-��5�'h:l2od����O���P*������N�Y��L�O���_Pa����OD�ӞgD4���x�HQ��K�ƦU�� Ԋ��.[�/O�Q�J
�p<I���||�d�]#7�Ui޴V��!J�^��e�%��W\,���()��dK���4�?y�A�'�\Q'�
���I�Oƃ����O�"|"+��c��	�/UWB�����W<��i�R ���	Pܨ�X��6À �E�'�	;5�4�K������~��"@�[�"���a�Aj�dʶ�:� �B�#���'^>��r��	��X腆Wx`�T>��O�Y��I d�|QAD�(-�, �L��б�c(2]ѕQ<K�|}�*n����2�GZ;jID����H~B�(3�>	G��Y޴(��OO�O04A��ܿ�d�&�!"44"�y��'�y�✶SI(�& --`�����0<���	>�:�ЀaR�+z�4�3`�\x���4�?q��?�`��RbZA���?i��?�;]ܬ�SaN�JT~���4�ε���^�{$1���X��0�nQ�ݘO�'��Y3c�N6@B�!� �ĳ5k�;򭓽�6��T8?N ��޻��OtXe �	��<iS䌣L�����c��`��S�nA��b�<�GhD���?Y�?�#�&V��"�
i]����M�<�!j����PޑC��eY��~~�O;��|2���%i+rP���N&v3�Ļ�*�@�x�R4��*W����Oz���ORT�;�?����T/] ���O�,|l ��q2%0�<{���(���@\�!~��*��I2Cd� �2��}Jƌ�L��Y�h�R��
�D�6�A1I��H �h�15�J">Ysc�1�(Q���l�^|)�ºW�*���MS��iV�O�h�~���
�d�Հʉ&ܠ��h�!�d�h�m3�+Q��0�#��V�b�1O�Tl�p�'�j��wg�~r�}W�YAg��X�d�J&���!���?ihX��?����t
A�^uZd Z�/��@���\i(PX� Ϙtִ9�`HX�"�rd��ɖ���e˝p�h���%τ2}�����@=�e�� \�b��5���U���O�8��'�7�GD}�㎺&���7`C"��&gZ�И'V��'�
��Ԅ�7
H8���mO>W(|5a�'@�7�8�~�r6iR;Yr)k�Lڰb@�ī<qKJ/a��Iş0�O�z�j��'�����dì_qT�X���]i�����'(&_�Lo���t�U1d�Bqp$���'���#�.� �#W	 �r���$��;#^Y+bP-h�-�3��"pQ>�+��[�А����#X���U�<}�AC1�?���i^�"}��'Q-���#�!��XR�jT&o�$0��'�D�!���$��!��.Q�G��Ó ��԰r.O>5��Y�N#C�1�`S	����O&������D��O4���O������s�^�1�����jЕMU����� p�!8�.U���7�@�#�����|�N��,@����Ű���'�(�Hݹ�h��bG��lڢ,.�z���|�.:VĀrR��9���W�#a�"���ᗏ�O�i�O@⟸��Ǐ�}P=����-��E�+D���`G ��co�"0z�(�a>?���)
+O0d��ɞW���"���<�&�ꗎ��ZS�-�V��O���O���޺[���?A�O��vd�1q.��� ��x�a�Õ2Ugh�"�_'j�I�����0<)��I"��Es�GȤUؙ;�(�� v*�#��P�vF����R�ڈ��ɀM���	��k��É	AT�(�"�ݺ�B�j���l�R�:7����׬S[^�Չea^�P�l�"O�iV���nq%P6!��#@@IS���g}�^�LR����M+���?��ѣu�����k�=�ą(����?���F���?Y�u�Jq����A�-�=N��fD�c�>$	1�Ղ�\��4#C�X*џ�j�	�aeFP3v�ߗ>��1Q�,���F�R�%<����JK V��|)�OY���˓e6�	�|�d����O�]	UI���`��F%܍/B�6O��$�O��"|b" T�)��p���E��L� ���'�r#?ӱi�D�Z� �(St LI3�� ���B�uӎ��R̦9�&�H�M3���?I���$B��?!���x�t�{f��G��X�a���?���o*��H�Ɲ%B�H�K?�O?�ӓ{�FA a떩�r��t��'�l�'k]Qt�Th;&M{Sku�O!l�QA�y��%
�W�&P�L�ď�O�@lZ��M�����OWF�*�k�(E�Vl�rM������y��'��y
� �m���N�H�\�����x�|�2�'�,"=Q �3#���A�T�l��T�V�1+���?��f���u(V��?���?��
��N�:�0�G:C��Y��c[�#?�E0 H�S>�FO�����C��ḩ��s>���J�L�Y@͊x%� ���W9ڴ�l�cD����E������?;`$�i�.����קe����DW���	��iB7�O��:f�Oq��I�H�ȏ*G:D#7���49����Dh<	'ъ H�5 ,�����E�W~�?ғ\��I|yb�W3x�*%�� ��h`L��y����zp١lF�n�2j���y2�%zģ��K�i}y@�Q��y�đ�R��`��M\	4�'#Ĥ�y�/.���DcK�X�\�;�o��y��C��K���K�X`��'���yҪW/t�"�#L+S̪�#��W��y2�[!VfZDRq&�uN��d
��y��2X=��)���fD�Y���=�yrI�>4ᦰ��`���!���yR ��F�@sd�AVZ�p�ɜ�ybl_�(�֝)�24�0ݪ��7�y�B�&F!�dӢ\�<P�v,U2�yR*�� ���R(� ��E#�y��;vҚ(8��L�\�qvn�#�yNJ�1��ja�B	e�������y(^�'��i��kD��P����y��C�>�����%Y�&%2 ��3�ybj�<o�@��6mIi�2��'��yF4}
�0�QF%/��ԹDn�-�y��X�r��Y�D��(G��B��y���
�����	�| b���y��'ԃ` �;*J��(Գ�y��W#u8;"�-���7Ґ�yB$�*V
x��W$Θq����#@��y"�O�hA'BZ�6�+���2�y"H�(� H�KR�S�*@ qH��y�3	����3��H�ܘ��j�D�<)D��uz=R�Ɉ�oBڔ���S�<�%�j���u�H�R��`�&DKL�<y��QP�Dy��2x^� �ECE�<�e��.��)j����X�^d�э�~�<)�HΩ����GU��`	�x�<�e"T�e0���f�"A�1�5D� �A�,$\R�H(h�����'D�0{��3 ���P+�2/�X���w1�84 �*O5R-1���5*�0�=�Ͽ.�P	<�)$������F�n�<�����M���W��&}�i�1~���'��'G�iP�c����Θ���A��'u6��g�%.�t��Y�1q6�	�}N����i��Z���-+q� ��#(�
e�v�ń%�B�DZ1 �N<���@�-7\MZ� �W�Q�t)��>M��s1� ov����"�Z}�U�Tf�Z	I�j� ^�ϓn%V�:@%��"�SW	_�8\#�mJ�C�"	C�'"�O��c���6lV�Ä�j�fm��nYV�~}b�j� x�� �"a�$f��!E��5r�F)�)36Ip[w,-	�N]O,�Ăc��5,�y�g�ݲ o�B���7�� 7���I���d�;�����t�89�F
V�l��ʐ�L������i�p�b�/{,��@p����Z]&�"�.}����ŠP���6	X�b�
���fɅ:�f���N��Ynͺ4�i�Z����U��0�K��fz��ՠO�.�"U͌,c;��'�
jV�Z� l�����4%�ʈ��8�9Ҡ����I��i�Z�	H�EvX�F��9X��D
����m���a�.�ʝ��^� ��;Ԯ�a�f�?���$��
��By:
�����>�j�Jd�֛0߸��#���ĺ���`~��Hq�R89�
�����޺����@�0m��h���~`��Y"Y����o&Y�u�� vȚ$��	�,d�RR�=?tR��kw,�EJ�.!���#�(U������
�_�d�]��|�H�J4񤞖212��a�"Ys,�B��W���h+�K/P}���[�ZZ�cvI�.\򇢒:mr����6B��A�6��'{ :���gЋ�O���j�$'Z< ����fB6nY,����)w���$閹Q>> ���:2=2���M���Zg�ʝK�05�p�A"�Q�#�vr����}��<;�>���`ҥF	Di�B%�X��RN�}�6�rC��ꕥ�^e�	G>p��I�A���TQ�vX��0f�
�UP���F�l �(�'�� 쭒v ��QF5��D��<к!����
)�B�qiDI�4���RX�|z�ƕ�V���(�1@B�ys�Cەs�Lh)��ɂ8B&��'Wz4}x���>��$� �\xp�Oc�5�5 ��a� �I�dQ6=8Ho!�O��{ĩX������~%,HZEc�r�$j
�z@h�UƋ�Q<�! .��N���Gx�A�66u.��ң\
,E�E���� )c�]k�ĴZ:#<�RCW�t�
Ɉ0KG�a�F��P$�-=d��V���uAVn`֠�B�_"*��M u�Oj�O&�8Q,H�K2jp�4
}P�s�OB��U@иu0Ya!��,�v#�'�/��Y��%v��-�tcb���N����k�{;�ɍU?��q�ZP��a54�D�Pw� �m@:Z�Q�E����Q��TS���s�	�+|���Y�CBA�@�l���
�@�*<�ўH�+G�eIB�	26�a䠇)AIzH�v�I�dt��񄁣^&$�%�F��c�_�f�x�׊V X�h\{�D/f�p"=i��x֕�T�`�ꄻA��Yʱmː<��i�[��`i���)76,��oæA�|��;?e���O2x5cS�H7}�Nc��GJy҄]�b]�I*6j	� ��?�q�����O:`�F��F�����b�u<54��>��ii�"[�I���Rs�C#:���1Y$�@�t�豲p�6WTv�ԛ��aa�,.���#��f�J��/�-4�Y�sf�g~!(�eɱ%��`�ē+��##o�=��y��'�Pᙆ�rr6����w����@�o�@�c(��
��؆�Ъ\�ay"�@C�,X�Á9F ��8JS0�8����NB(����AF�B��m欩B��*uhT�B�� q��OЩ$��b|t��Ō�h�ީ��&�.5�V�xlZ(g�D�i�"O��B!�SB\��7#�#"�X�OP8�"ش;yfEx�IT^�&�'B.�O�T��C,wp��k秅k��I��'V
8x����J_Ab��V&.tX�ˋ+��
 	
V�xD�eJV�Q����ə?Ү��lݮgQ�m�q�B�y>l�\j0Ǘ�s��\FKɚO�E�D��g?��}�{�	*󖩪G��S�dB�	S�b�:��E�C�e:u�?GHq2�#V�C*Xu8 �J�ߞ�1@����>q"�w�e���Y��Y�1��U���@�O6���S�EM��f��"}R�I�2�m��j�O%�婵�#Q��K�}(e%_�=�֝�g�d��T�D��=u��f��T���?P���'0���	��{�J�`!���7wP�P$o_�_���K�� @���2@�=N�ZE��@]� �0( `G^,�p<)�� qy�)
3$�1;�Ѓ^0>���ħ��4K�<�'�|mk�_�e{b�C����-O�@�n�CC Y�H� �٧��Ox0�H�ƚ�����{�R�{�֜p�@.��;x�C�O�!��S%21O����y���J�׌!@�eB�C� _�(�b4!�/�R��H��`BE�V�EXx���:�t�QNF̓zKt�U��PP�Q�W1��'��`��e�z���$]���₩0?A��H�V=
ܫE���Λ�0-z��c��	�S-�Wh�@�󬐯<4�q�1D��{U�Pz�n}O
���K�����*e�P�$��
_#�h��+^��̓BX��1��~���J�(�Ӽ�J ޞ�[�N�,;1C�MJA�<q4['Z��gP�y�α�I6��TCt��m�d�3�+~a�d����쟐�ɔr"%��:Ҟ� G�j�P���
�CUڠ�VR�Xb�@�Ϟ]���#G�B-�
9�!n�!}�x�I�p\w�Q��0������U�TZ�U��*3ғT��D��'�?)��@
mk*˧e�83\r:�0���$��q�q��91��7�OL'�V00�pq���G~��}0�ib��N.1�։�8�̄L?�H��O�i�^�"&���RN�݀���1t��H��'�Hy	��V~,��P���?��T�₄�0)�0c���>L���/O��O�Y"���Ç�*}8|5����np�2w��h�q�<}����{(��Q�/W�F}����'�RP�T�tI�kF-�?9��Fy�*�4|�a7��+V�t�����'��p���G+��Jǯ	1Ê�`��i�Wg\5�v&@��z��P���✋Z���'�L��F���&7R��  @�]P���Ô�,H�jv+E�M�5���3}"<�ұ�A�۸yN�
�⛋~���R"O~��J̠N�$\d�Ӂ0�`IH&�Oth!�� c�'-��'����D�/1�ZT�f#_!}�f���n�qt8��=LOz�x3B�x�X�Ԧ[y��eC0y�vKԎ^�8t±V��%��Zw � o���EyrjM�=e��IP�*hQH8vO�+�'�I:rG�.'�u�W���OѸ�i�y�&����4H����4s� �&'��p>!3BY<i�Jܘ���+z^4��f�r��đ�ԭy�	cx\�l���M��?��ex���0��=��A�]1���I
�'.,�!@�d�,hP���O�:���ʂ>Bt��C�Ò柘�Ч�
�&���8S��L�Q�D��0b&Gf"p��'�~e��s�8	�C���͔�@�H��U-�i���2p&��l^L�O��D��O� ƨ`���<>$î��H�ia󤍉N��kef�*���r�����MŒ�lR;������}�.|k fC�d����ċ+%vd�+g�ƙ%캤�ւ(]�PfOV\��:⒟�tK���DA5r*�e��>J��9����! !񄌪{�ʠy��#^��Hb%���c�<}����g�9��a8�O�Az��`�~4�����2����R�'@��jd�E5�N�G�OR!�D5U���1�4`���"O����@$t����'����p�x��!i����5Q?=1�"د���"c�Ɋz���Pl*D�$�g	�`�p����I��"XSME�;�0
"W���dE\���ē%dl�s�\�j<\�(�B�[I�ՆēF�����n�y}��j₃�Y�HB�ɏ�me�I��OJ��p>��a� `���B-֫c��ys-�mX�@#��J�O0���Jz?1 c� jiq���.�XIS��P�<A%K©p]��A!D�r����A��c�I�0e: �A�W)(dHF�Tȇ�Y�f�1�'�"nx��R%���y"M��n�8��GN�[$ :�[Rz�.��X����ɁC�`����L<��g؇_��1�&bȯP�8��-HH<�	?H&�q3Aā�	4�0��G�&fP��`jS���D��p=�3M۝@����A,f��2�EI�6\�*i��4?Q�')0�t@V��V��M�r'��
�����e�x�̸kw'� x�!�$X0VC�b�JBf��
�`�Q�%�'LTp�
�u*�	�b���S
 �Ԩw�8$��
�9��p�$��K�X�K�'~�+��Z^���G[�m�(Ш�FM�f�zq����y��:���k����xc$!��h5Ǒ<i��J��F��<yQj�!%p��'����k��I�a:hl
�(d�W�M1���������|��S(k8p o�.�����g���ZUJu�с�b~\�9<�������DȦ%�Xst�	�=VJܺG�"v8!�ğ�h��F�z�ba�֠Z'H�y�'u�����P�
��������@�J"��2n�Xh�T�=�֡�#L��B�I"x�as�&�[Ŝ-7�4k!�%�����)VB��O������a�<|H�k�}��[b"O�̱%�X����Je`F�/�>��"Ov�z���.�R�i�/N�k�"D�c"O�Mˡ':�T��F �K�J�e"Opm��J�#=x��b*
 ����"O���$��'�B��%B�
�y�A����@V��"9D�iț��y�"� 1p�XG�/��H��@��yrA6jf,A����Š�O,�y�H6/�6q��Q���b����y�.H.E�l�h�"аJ�
�2Aа�y�a�)�q藏��HX�E�q��y���9dI� Y� G�|�Ð���y�,�1y[Yؗ� t�Hy�@�>�Py2�9UD!� ���;���eRK�<��eAp�%�Ν�@6F�2P�F�<��l�7��2���3%D�@UC�@�<��ـb�`q�"y�2�P��I@�<)��T�;6�A3R���y�4x�V�<IGM�~̸�娎ʼ���@z�<���<;6LwH�7�4��&mR�<1uЏ|8�s�J4�Ql�O�<A'�����Ut�����d�<����5/���U�B &r�[5�w�<A�[�J���nƺ.c1�`%\W�<I�@E$]��b�mގq�H�31�CP�<�!�C%Q�DV�Q
�ҭ��P�<�Q��aVYC!^֜�d�L�<	 �z�i���j^d%+���L�<�E��vSx��	*_d�r0�o�<�#�ƭ:�j�k�A��;��<ʒ�A�<��c�X�j)E�2Pr��#��EU�<Q�����p��DM�DI����[�<� ^}sq��E���kн~�xѺP"O=#�׀|��K�<'�L�7"O��*p�&X%2�k ��n|�z�"O��"�(�R�8b友:�r�cc"O��'B	�sx%�dD#&����"O�\��`����=z���Wͪ�"O����:`�d_*�Di�"O,<��n	3��	��vu�C"O6���$t})s����hv"O�=��D;]/"�*�֐AJlEң"O��S�=~V �ro�l<j5��"O:��6�ß8=�e����{�X� #"OjEC�� NƨSg�^ >ل=8�"O�t� ���4f5�#�E�M0}&"O��z�/��.\�J�(��q+�I�"O��8�� 7si�Y�'�"�zQ��"OX���JF�+������#D2���"O����ǜ�W�gfR�kFNb "O�ѐ!-�ca�% �F"629@#"O�����w���ԣ�#$hxY�"O�0"��,0��\1���y d�Ұ"O&��C.ƌ�bb�H (I064YC"O�p�b�ݼ=�������zxم"O�����F��ɋ�"�"��bV"Oh��ðK�x�s��O /����"O��91�G�O�t�(P�Ħ2s�8�"OA
�Q#mSB���%Q<ZE����"O�4��ՒM`t� 7��n<����"O*�ǌиm*պQ�Q6N/&5�U"O�������Τ�O��g � "Of��@˹wVJQH1�	�����"O�@�@�2B�ļ�$�<�.Bc"O�L@��V(��C�
�]��[�"O\����'���g#VOQ�93"Oz�B$�9B�"*0B�Ld�"O��#C�"�LD` �ԟ8Ad�p�"OL���eD3~��,�1F��r%"O"�	��ףwE:���S ��)H�"O���@�K>dM|�Ӂ"i�",�`"O¸*��8n?�x
U�T/9ZD�8"O��[��4�Ta�#�S�H�C"O���$�A�TM��J�/��x� "Ob�*����p`j��V�l�<��2"O�eseRJ�
B�I;5ؐd"O��r$��.$2b��@RH>x��"O
��uA�7.4�c�)�lʃ"On��L�*g�, 4�ܧ
���H"O^�Zg	X$>Z�ݑ4�F����x"OB�����)9<b����d,�U�"O��������Xi!`N�K"�-˒"OtRQD�(�\$B�H��34P�"OT����*"�}�&U��@0�"O4u�UjW1R�vAꅏ�U�ѣ�"OД��i�89��L�d���#F�(1T"OR�6�Șk�"��G-�'�����"Ol��ծֲ1w������"Jy$	G"O �!p�vz8�Q�btX�j�"ObQ*�L#? �`R'W�T=�,91"O��a���D=����5[\P�O�dM')7:C �Ǌl�>��j�=�8B�	�{uԤ:�M2N�
.B�"?��	°8L�훎/�6�IG�P&T�!�ډ0�$(qs��'�J-(VG�V��	.b�Q�\Gx�M^�RR��ڣ.�5�r�2�	ӑ�y
� �h��E�$Nyd`R% =�� Jǚ>Q���=�瘶&juK1�8Lt�����]؟���~�n��DU�fm��P�ά8�ܰ��<N��1Ѕ��*=d�T�Ҩa�[��N��=z`�\�~s3�ڏ��X�ȓc�Zu���\3.���EN�6.ňa��PҪy�4��iPa���ȌŇȓ�&��_�5�niz%�\�\�zq�ȓyb❰C�N3!��Q>
���ȓN�*Xa���"2Bd���@�6QUN��ȓBѼ!�t	ۢf���$�"�%%� F{����R�<�N�J"�%+P�3�ʙ�y�D
4I��̢#����"�,�'��T��I��pUX�m[��h�y@��u�JC����%r�S�NaN��e�O:XBO.��V�Y{͒ j��§[�-%!���={aV�ܰJ����g�	Q!��εq~Q)�nً��H�FQ�!��/�x0���1�n��"g��Us!�P'cB��+��#-��Q٢/�Qj!�D׈2���˵�X$<�y���S!򤉁|�r���U2n0 c��+9!�˚G�fL����f�b�a��e�!���qBup�n-|�.u��EV&!�A0&%��@����]�V%!�D�y?�a �#<� �u/֋/u!�$X΀|��!҇?q�Y�r/Ҁ:�!�ߖ ���c쒀bp��0�%.�!�P�T* ���-z$]��c^�!�$�\������ݴ{u�i fC['_!���-$� ��6�����AٙW!�	U(�0'��=
�4E�3[!������ؑ�ѝt�
a��@��04!��$�X��ߢn,��� !�$_c|J���I�1��@��Z=<
C�2jJ^)�0dL%OF��A��'&�B��w`�03�)[�M�r�q�j�<TsC�ɇ"����],X��YpԮ�>V���OX�=�}*QL���sua5G���t�Md�<���N�D�l�3�M�$�09��Kj�<A�$X�y2U�0L�*B|��!�P�<	��'mޱ��դ F��A獉P�<�2��&A���"��#�ڕq`�e�<i3/-j�5�bE[�`Y���#"`�<�P�BLUB��V�Ys��(%�Z^�<YTN5�B����|��US�<�@��\�D��T��V��b �R�<��"۸.H�(�b_�t�`�JwOYQ�<I�
&��t�S�	�i\���F�X�<� �L�K�4;d\4-ߪ��,R�<�S�ʯz֍���S�`#�h{b�Xr�<	�@��n� �� ��H&X��r$v�<p��8R�v�`��	Ԯ$[%\n�<�4��l�H��.��2D�:���k�<���(u+�lg�H|J�D�i�<0�Ԑ5G�蒗�%`�Sa�f�<��!E��^y�!��uF�L3m�{�<IteY�:2Lax��y�����J��yB'�
z�hM� �y3N������OD�=�ORT�j���%qAn�#�J�`�K	�'���(���:N�!�f�Sf\�� �7�S��?A4g�E����K�Ħ�z2Bu�<A�Èe��d����(H�$ɻw�j�<q�)ۙJ{�`j�^ݜ�S�!i�<� �)�Mb�~p���&`x��s"OV��]
]Ğ�M���v"OШ�����\X��h�.)bQ��"O� QnѠL"L1��Z�DjN��"O0�����1���SPi60{�U�&"OZ�j4��5J�b���%5p"P�"O���6���aN489��^]<Pb�"O>��+�*�$q[G`�:]PN�!D"O��
�'��P48�"�e<C�HT�Q"O�����D:��:P��&�J��"OȀ�C�Q"c0����	60�fQR�"Oj<+O�/��b���	a"O�E���Z�
���T�6�*�X#"O\d���S�Oڊ�Y�ҕBZt�[�"O������,kJ,9��؀=P*��g"OH��%��zG�,:w�[�;���#"O`�3�&�h��Yd(��=�,A��"O��S���Y:*lRdn��8����"OFh�Í?r�*	��"O�}�#�C�1/|݋R�C
w��R"Oހ�1��"x8(Q���?D� |1t"OD��K��	]|%IFԅ}ul�J�"Op����K��
-å�0#Y���"O��w��2\�L�a���=~Mmٱ"OFa�FH�� �С��d�7��yF"Of�iώ)g���u�Ҵ�D{T"O��ZG�A#>�j�9��`
�	�"O6�Pa�Pg��I��K�p!"OT� ��9Hl�5
H�u��Py�"O�Ij�nH���铦`Иp����XD{��S9RdK��1�d���Y�Xú��'j� "S$A'��4���զ��'=��8p�28�|up�C��zd��'J�):�'�<z�]���Z�y�4�y�'n�\x1�O�r������s���Ǔ�HOx,��1'�:@��F�8��<Y��'�D����˱:C��x&�O�pOʈ��S?N�P��� �B�,�<i��"O�t�"����2"&�t����a"O:�@�ҲA��Ğ�[<���"O�H�g �����֌[=?,��"O��@���5�
��i�`"!"Oz�Hc�ק'��;1) ](0�7"O��C�2 � ����֧J�`�G"O �4�Ǖ*�)�w,�W��V"O�|H-��Ϝ����[���"Ob����$=е�^��LK�"Ob����MK�h
0���{7��D"O�����R<\��eV�O�\�A"ON��WE�bTpU�]$��=-�y�L�&T>��&��r���#�=�yRb�-6�X2d#��R��!�����y�D����T;r��*T��4�K���y�LG�Ji(Q�4E�i�7�y҈M$e��h��7TҘ�*�H���yr��b����쉮{@�y�#d��y¬#'���4j�+����/(C�Ik�
Uz$��XG��X��>v��B�ɷL�N-����_z�������B�I�̪�e/s�<z�NK�|�B�ɘ$cԈR�͆U��=�#˷/��C䉎V
,i��I������� s�vC�	fj�:��Ѿ7T�<�G+R�`C�ɔ�!�$ �*��!PXfC�)� F��h٭~+0\�	�K"�᪂"O���ѭ@
��lڶ�N>m��S�"O�5c\*E�$�9$��u.re��"Oڜ�@	��ј�r5f��+H�q�"O�!�Ǹi<
� �䚤���1F"O��#,�<'t|��-�b�"OU
aI�@2��%�U�C��Uh�"O����#,& 5[��
�N�Z�iq"Op��q�4P� ��#�l9�"O�}A������3f��$P�V"O��EY���){ �S2�p�/�y"BI�z����	��h��v�Ә�yr̊F�JŁj�5^���/D=�y�`�3Y�!�D�Y������η�yҊ��q,ay"�E�����\-�y��*g�:M�IS�Kİ-󐨐��y�q�䴋�́@l�h� ���y�Ł�̶d(bCU�L�Xy��j���y�j��mQ�	�@��<Z�u�R�3�y��p�B-�S:*���"ݨ�y"B�)O��	�+�"k�Ҙ��MU��y�m�5΢�c��\2�b�Ф�G+�yr���D����X�#���3�䚺�y"�,`���X�D�X�A㊚�ybǖ�m��"#� r�0�1�X�y��X68����BW� &(�5,���y�%�B�h|��ݢc
�m�yb�V"e=z	r��*�:T�V�E��y2�Ú�P���^��ޱ&*�%�yR���D�*1�c�X0(�V�Z�o��y�ܛ&)��+�+&�A��y҃T8?\=�1A�� �$ɖ�;�yR��}�.����U��y��7���'�		F\��U�.�y"-B9)���h%����%��(�yRH�	&q��9��̔ ������y�d{�&�{u�v`���#@��y�AZruB���7Z$ ��
�.�yrǂ�y��8��(�O*R]	e����y����,rb	�
NZ�L�)��y�JȗM4�R�jIp��bg+��yB�Ą�թ�3p<��zv�+�y�<)��-��F�i?l��ee��y®۾�mV`Q%
+44 �i��y�S�:���� K�|=���P�ձ�y�Dͮ������I�@�$���D�y�L	70��P��Ό.b�(@���yB��5d��C�/j\ ̑2.@��y2�M.��P��DdM~�X`���y∜�[O��0oZ�P�͈�b�!�y2J=L�2�"� �d$��%�y"�.h[F��ǃ6q��Q�@�&�yHA�5�4��a�iX������y�J�|j�s���$P��q���E;�y�L��:M�H����]�༁��W��y�I_+� ,���,�NȰR¹�y�M�Q�F�K�+��M�t*�i��yR���VH��"�?}d� �G���y��)����&G�5�fL�S��y�KS3u��}�+���s�×�yB��:�}�u큶$�xD����yr�0(�i Q�W�k�^i��X��y�H��jF�HCӏڴ_o�����+�y��T�{�~���JC�xx�jU+�y
� �}@V��J���:�(7Q.z�S"O$8��'Tu3 �P��/��x0"O�ajP�ڋ�X�3�+J�+°�k�"O�t�6L�yjnA!#�\ [VФ�"O�lG%�9(�a� ��	N�,
w"O~�Z���Q� đ}2�u�"O��q%��P��h�g �:�j�ȧ"O(	82d\.X �܋FO�	nx�Ųt"O``X-���0�{"��1GPH9T"O�`*�,mT�y	��)Y	6�
s"OLI�Ӎ��o��!�L6M���"O�ᡦʠg�.
զ�6�*�`"OR}96Gi!((�M5\�"$)u"ORУ��	[[�t��/3�е2�"Ob-�DK�&�*���bD�dx��+�"O��@�h� T�����:bt���"O����>�n(�@��$WVq`�"O�#SÔ�}��䊐Z.^�|���"O��aqŒ�?�@Ș@�}3�+�"O�qȡeB�VT��ВdFm0,,Z�"O$�acH�P%�y��� ��(�"O�� J�+
d��QkJ".D�(	p"O���bo^���|���Ո	�2���"O���b�(&r��IT�.wP|�""O�Ȃ�R��Q� �3	l>,��"O�Y�l�:�|�"ČH MY$1��"Ov�Y� *Zx �
��L�[��ͩE"O����*YKn͐U�\
��i�"O�,@�
\��;ס��`�C"O"ઐY	!P��&���!�"O�����R��q�L�	I��a4"Ox5z d���2����Z�#H�	A"O�%C_�0��.-�`�C��T�!�(����r�V�d)Ƽ"���){�!�$#Mi�q�R@�r5����!�!��y���36�^K�բ�C�y�!�d����c YQ!<42D��G!�$� �2��P��J��FJ�	!�O�`H��!eI�Z�]a�đ�!�$Ҧ9b̨a%��x��h���7�!�C�D�b�q�TA����T�4m�!�DD�u�'R/�(�.�
i!��F�e�n����3�H���1N!���f�`�3��F�[��<�_�1!���x�$0wg�4��	 $%7!�Q�"R���ȍ 8�9���Ơ�!��W<e�7Lȋ-�4b��n�!��%'���j2���4�0 j"jО �!��S�=����A � ��yaa��(f�!��*=���� @��"��}I���u�!�$�r`�Pڡ!�7HeW���:;!��On#b�"u��2|�FE��J�a0!�dO:vB0	��<�.8��J5E!�ݾ==.�CѡX<��!� Q�d'!���ȉqG��"ddu�S�W�?�!�dG�6�쩺�)�FJ�8D<Q�!�d�i����V#%�vJg�;#�!�$Wg�4�Ѫʨ|ۄ)�r�l�!�N�f	4i��CA{��j���7�!�F�!� ��I[(FVء
6D �]�!�䁾8�BT1g�N�9!��҅ƴp�!�D��$����iG�(�eD��}�!�d֨#�䝫U���4B�ڞ�!򤒠Ll����-�N�{� Qx!�� rl�#OQ�Gƚ��.1m*L�W"OD�Y�� s���E�F�F����`"Oh˕�{-9qG�ǤM��I�R"O�%bC���#������9mt��"OT�!i�#e�슐i�YU�q�"O�=b�FS\�R��</�]�c"OJa!�����",���M';*ZuC "Ol��"�\!Y" �^'`Ic"O`���S#9�bЁEA?,R�4��"O�t��њ��ы����f�#  #D�Pc�aդS ,��Kp��	�r=D��Y�!47���G����k�g;D�P�gh��2Xe�Ä�K�tQ�<D�,�Rk�i�-#�lҘO"6�Bd>D�Ы%��*NYn� V����I�!D��`��!��C1+�����e�=D�<�eD�$3�	��N;���2$=D����E�(J�H��"`))��L�!��D�oD�;��ͷ7���0�;t���d�8 �D{���cMH	���E,�y�-[=%�N�S�`)�hPpNN��y҉�2	��#&d�|,`K�4�y←|�*eJ�]�\(��Ó)�y��HXRaiL�\�$H҇&�y�
<&�0!�q,� ��$ǚ�y�*^�~k���R� {Y����y���4c�����*
�M�(C3ʛ�y��*;�,�H���-�0d���[�y���8G��u�?���!5hQ
�y�!�.O�캷*��r�\K����y2��0T$��Ѡ(�6ql*�kC��8�y��.UE�U!��X�j�� ��8�y�-RaaBA�!P8t#�9���U��yg��Vk�\[�т[� %Z���0�y�D8�4�0�)�<Z�(Q2S���y"�	�pB�I�v��Q1��s2f�y�G	"�#�Y$AI$��1dH�yr@د8��a3D�&35���Q$ؙ�y��uo>ģW@=,��������yR%.Z��� B�N%� Aq�����yr��8zfH�s�%N�sw _&�y`�#�@46m�o�I�񭀹�yr���-�,�dԬ�d��y",.S�|Sf�	22~�i����y�ʟk"�U�_k��%�H+�y@T*-���2W�]9fK
x�����y"E��pa|��H\8]��$� �y�Sy�hm+'8$� �F�ybO�����aG�BlY@V���'h�a�B��^�D"�j;����	�'ٰ��6-7��l������'7�A�e.��=���C��6�:�'��8���"�~����'�tc	�'�q����z��A�R�R~b.���'���C&F��`��MWgB���'��Hi�@�n���K�f|�=��'^��C�A�A�ā`��P"_hd{�'�$}���2W�d2��.R���'��d*r$ xK�dз��^Y�Q�'	�P#��KAj=�`�[�Ldx
�'?j� "nM�st=�E@�T�.���'D��ic���\a&��b%�G`��Q�'�=��i�L��a�"TQ]�D�
�'��d�Pl<����L�H������� `����ŹT>��@���Y�X��C"O �䢊�Mp� bo�^t�ر�"Om�M�,�x��!/��Zl�j�"OZy���r%3�M�!]~� c4"OB�H��@�	z���֢���IU"O��@V���Se�#��ΑZ�Ѡ6"O
�4Aʴ x���ݒO�<�J�"O�q;W*�����a�k��{y>��"O�:Wg�#E�)�2��n�ԑB"Oh*��ݳt.�:f���Ĉ�zM!�d��`V�	��iN8<����@?C"!�x��� EV*@4��bN)'�!��^�ՐpC��;2��%$2!������c+.XL}���(T�!�D��o����:��@��*	R�!���
����S���\v����^�F�!�䔗z5h3�XSt�8��+s!�dѥ�6u� M�Hs��
��L�Lz!�߅����
�b\j1����F[!�ą��4D��D�9c�HSg�..!�$�\�pv�C����2��Z%!�$
)cgd\�ƍ,_v\�b���!�䆤�X4&�[ԅ�Ē�6^!�d��-�Ve�S� <�	��L�"@P!򄓘{mR���M�B��xr+=l!�$ר}�X9 ȋ:�u�Fj�+|N!򄆳�\�=sL�W0N6��	�'�P���g�[D�	�-X
�4��'R�l���ؖ����Q������'� �p	��C�ER�xЊђ�'��(�e%L�a�*U3R ҥu	)��'}8�YU�oqp��Q@3d���b�'���Q�g��D���`aE�:ba|���'a���S��/՞�Y���bbr���'F�M����܁�p��-G�չ�'��T���E�p�P����!��'�$��d˪2�"i��J~��[�'�BDB!ԅe�)�O�>
�Q�'�$�B�M�,��MQ"Q�u�'k��F�q�0LA��O�6���'���r��+Kn��kS��S�8��'Xذ�H�H�Lp
��V�?��t�
�'l�8C A�!-��*D�X4hB K
�'�H�S�F	T���+�G�0T���	�'L)���a	PI��K,C�Q�'3��*Ƨ����`cIR�H� t@�'b(�J�$�	Wn<��BiĴV��i�'F� ҕlȟu��Y2��Ӑ#5����'DA��.Y�� �J# 62r,���'w��0)'2B<����-{��'6�yz *^��t=�­� -�y	
�'�܄��
������&����'�f�x�CͲ8���ԁ��'Ҡ�0f�J=f7��@�ܤ�j��
�'X>Q���b<��� L�{�( 
�'d(�¦���t����L�i
�'�z\��K	�����Kh�^�`�'��sT��4:���W� ����'δ���č*+䴕�RBE�D�Z�'�p��Gͺu��w��Iق�!�'q���N18NѣA��2��	i�'ӌhp�`�d����E�T���#�'��������9x�j�x��'�����a��6C8S�Ww��j��� �����W�B��tb�"ˌ܊�"O�5����M����B�_��5�"O���V@�+	��#�N?�ȝ(b"O����ƋU�V���,��M���X�"O
�&�Q�N�H;�M\
8��|�s"OJ̙E	�9(L��k�� �Ν{�"O�Ȣ����t�1�ꛑh�����"Olh��0z~ �3)	"(�D��"OFY��iDc7F�Ԫԑ"!BhP"O�1�R��v�~qS�"��kʹz"O>�8��լ+Jvq� �X�b��+"Oh�YT �>xUF���_�r��2"O~BUkǋZ͖	���ƃ�X���"ONDY�i��R�Z���̋=X��X14"O��p)��~d8S�K�;����f"O�(�3@��� ��DY�(�pU"O����bG�x��b���@��Q�4"O@���(L�R}�AdA��*z^@�"O΀JeA��{�*=[a��_d2�B�"O����;
��ӏZ�5H���"O,K4�E.'�P�Aő>o�@ۦ"O�(k�C>K|�	B$�wl�yC"O�bf�'uV��� n�m-��"O�@��K�8��qy�̍[�i�"O*-��_)XZ2Q���B�f���"O���v�Z��9�1�J<�,��"O�P�#xa,��O�\3N��"O���`�ˮ.�������G�N-2q"O��hS �0e��=� ���p�"O�(��m��@J�=���C<Z�����"O��0���,bEB5�H�!���`e"O�`��
�=?�ވs��30��"Ob��A��5҂�ذ�
2'��œ%"OT)ա�P�����;!p�б�"O�)vN�e��I	˟�{|�U"O��W��i����3�Ul8�� "Oư�Q�R�,�ԩQ8[��q"O�(��f�#��5ZB�R)5�E��"O�`�舖M���$�Jd ��"O�=PR���[���Ks�3���"O�@
HK(U#bu�ŋ�6e<�"O�%:�! 7&e�Ъ��v7N:�"O���"��|{�*2JL��^���"Ofh�"�8��Q(E�4�yѣ"O����(i����E�pR��q"O����[��D� ������"O2q���GJ6Y�p��z��"O�Q�b ��y��/�6)�0"O.�IQm�_��k�)MU�r�b3"O��xԥM��1��Ԛ?�h�;"OZ�s�@  K��-zF��&: b�#�'���#ߚ��1&�%k�x	�'�� âheȼiZ�/��P��@��',����߾B�t�S�	C�h��']x+ '�X:b��Y�m�8��'VVd
�)A#Y|ԁ9�(Щb��e{�')@�[��B����@0��J����'_Fx�nT�Sp8\���=pb]*�'����GY�H��	�AK�:����'��=B�%@�0vف�&ݑ}1��'	���1!��i�@�7@���	�'���!5ˋp�����7����']^"�@;e`�CG+�
4熤
�'�h
7��D�Mq/�*:��Z��� ��C4IK�  @raBS!Z�Ti�"O����k��ik��S"��[L60P�"O�����^!̌��&�5�����"O�<�fk¯_ uY %"D�E�%"O
1[C�[����������"O:	��S�wt�P��F�}���#"O���2*� 4�X��u���i��c�"O�p�P��:��4�ǎ�&�Z
�"O�ڵ�]I�ŀu+��I�Ht:�"O$`w,ڂ/騌���\���x��"O0<�EL&#�]I�kW��P��"O�֡'JEP'��'��p�"Ob�f7r�M��KA(MD@���"Od]8��B^Z#"hR�+N�a�F"Oܭ��֘�jaǇ^!b�1K6"O�����yZFŒ�g$\����"OX)2k�X� �s�V1
��=�#"Oh�x��E�J�����h �2��y��"O�-����m�=ɀ"�ź*P"Oε;�CX7?��Jg.��~)�Q�|�'敛�%
	������"c����'�`���n�w��y�!� ��ٚ�'��a��L�;@3 �R�õLR5�'.0�Ѡ�۫B�
��Hp6��
�'���8r!e����;
�'����?;����S�d�$y�'+��hb
����0�$
�p�
�'�����$'hP��K����	�'	�e�a��&�R�o���`c	�'l����2l���ܞM�)��'q態T$��2"�a
��D2�]��'Z9JPM�9�2IR2�ї0�D�'N� ����00��>�K�'����D���-ŒK.�R�?D�$��fK�:Md :$������?D�d�s��{!��sf��V�PF+>D�@9��Q�0�@a�6i��'
9D����cˮG;T<�1��I�`8*��$D��b'O������z��R�'8D�t����(���@�E�5��WO D��zGC��gPC�3l�+0��O"B�	��2�S孂N�~������!��_��թ��$U�9#B��&a�!���p;��w�@�R5�!���=]�!���(~�9�"��2��YG�R
?�!�D�#s��v�Y�<��� u�!��K�<�QW����|hr �_��{��'\�Ʉk^��D 7Ke�Q��r<���*�Ŀ<�|�OZp�N� �t�#�T�s�@��"O,��Q熰]���xD��?ߚ0�"Of��$m�l��MR$l&4��;�"O�)��!	�njIA!B�X2�((�"Ont; '-�Fu�u��)!49$"Oĩq2�j!�9a�l�kh9 &�'A��pӎ�H�L88�'px,Q�`$��0<��G�
���Dɡ2��Pֲ�B�IzA�?���YV�W�sWdB�	G�����%�]�'��-�4B�	�jۀu��D3�q��I�.�C�I�]��40`mU�vB��bA�R�z��C�I��$(kE�ʧ.��}���>�fC�I&{'�!"iG�Gɺa�1b���d�O�����!�6�H�`_�q$�@#D˻gm!�ȓh�9�SĊ�F�e0w`]<vɾ1��S�? �����&�Ġ�ψ7&褸�"O�A��k�j�u�PΊ?A@L��"O�hcƐB�8�8N*^%�p3�"O�] cڻ|��8�Қ1h4YZQO�1�R�T��Y���S:Q�ri17��<q�e}�a�6�	�༚���#�Y��p\���u�8H��]����6BQ�ȓJMt��ᒓP�lHAnJr� 1�ȓ|@�5���:(kD��5m	�팈�ȓ�R�b$��T�كQ��F����ȓMR���'��(��[��\�4��ȓy�����A�_����h)�9��q\a�G�J��x�D6%@��ȓ
2�$ieLĠZj�⥧��Uk|��W�2��yP�\BA��,����ȓ`�"�q\�8���/�#�6؆�uhf��0��c�Z}���_)|t���ȓr��*B�_9=��T�G	�v��܅�|��y9���L̺e�&aW�h�����m
��Pk��:.阤��
Hc��ȓq
(ؚ�`"{�F}�6��M�Ԅ��P}j	�F��?H��4 w�{Č��a `1v*��Vq�Hh��e:����iu��;��>Y;�}��&���ȓa��U��-$�tJ"��T�bчȓ&���2�|�!�A�=f>�ȓ~;
�r�h��T��if��D�(�������B'��ݩb�Z=b�ȓK�Fђ%��v
Ba�g+ٽ2��e��ma���c�!Y�~�{cd]J��%�ȓa� �A��:~jY�GEA�6؆ȓ
���#G�ȦH�Zt�E���&zZD�ȓuA���6��-<T ӖO0bl����3H(��ᘾx�ZL
�&ā���ȓ�`��O[��,�0�"I�ć�"R����?����K�"/>���>���{3M��H��t	%g %�ȓ^VI�w�'q��*HE����9�⬐�i�?�P�
���
s�2@��Ks�8 �"
#���A����tnh�����E=gH�@2HT�]8��gHew%��95���,I�^�����<mJ�'qCL�A�ļ^_�؇�D&�qE�'[��=X4@
>D��`�ȓ�Q�U�E?0b�\i�:EF u�ȓ_."Ujc�P,�p�� T5.-&��8�Թ`$�Q�3�h� ���l�e�ȓbdZ���.k(*���+�^��ȓ �f��#F� A�p
�Kн�ȓ0�����ϟT�F�/�>dr��ȓrE����kA+���a��LHH�ȓ%}vq�F�o4*ـ��<j� ��n��eE�	�e϶!H�E�ȓdy�� ��޾�d��LM�2jU�ȓ\�r���cA;@�<2G��kp�ه�x84:W�:��1��l��Q��RZ����s�L����J�9FNy����]��lV;u9Tlb��?-�]��D�xH�b��-�P�����%����ȓ+'||�Q�Ϗ5B�x��Q[��Q��U��2�"G:�l��C�-�&���l<�3�ŽQ9~!H�c��
�x�KĦEG�<��kI=>����*=�b&+HI�<)DȆZvH���.b����O�<� 0��W�M9mȴ��CU�{dT)R"O&�	�hY�^v���t�K�HCnE�1"O�̂D儗x�0��&ςX'�1"O(p��ƕE�����.x�!�_�$��z�D:$�,�l��#G'i����=D�|��L�d_z
L�y����ƪ7D�B$���|���bI��7�fKs5D��ɕ!E]Ё胪��i"*�"*O�:u�z�!�H\ xR"O�1Yc�	C��)�&��L��"OH�P�S�4�&�a���l�C$�d(LO�u:r@��E�� b��a?ve�e"O(�,�	S.l�c�P�eT�D91"OD��W�K�l�jd�H)zIR�a�"O����İH֌t)������"O^��e�U�Q ��B�6��	��"O=	�(?a�� � �
T��"O>������)֌D[\�9���|2�'I���G�90f��"�����ݱ�'��'Ɍ����S^�X��)�'�����b��	q�is� �{�|���'�@"�� (*d�Cs�ȼlj���'IV��F͘u���rc��fIʡ��'�ő���/Sv��"%H:\S6u��'����扄�[����K%T �{�'7��"V�W�ti &�	,w�l���'�j���*��_��)f�B�h�8���'1ZM�pJN	>�p�)׎۱Wlč��'
�XQ����eJ���&*�I��'[du�]�R0@Ȋ�-ך!�B	��'�ƍR��D0��\��^�&��0�'J��%B��"W� �T�\ z0�X�'����Z\�N0	tj@�K�,R�'�*��SkΙz������{�'�Ԉ@�"���#1bE�vfRx�
�'ϼ��EF݈J��mʧ��u1���	�'Tj՚�%*�B-2��� p���	�'Q@�Ca�2I`�	g��p�l0�	�'J�];Q.0\\㖏F�m�����'l��5�I)~v�A�(�Vm��'��xUgԞ<Ҍ�գ��'�:��
�'�|����u1���pD�ڱ�
�'�^mR@��7� ��w	2���	�'�D�r�‿3��P���='�<��'�,x���6e���f�˅	A�ͩ��y��j%��� Q�zM����s8�B�Ip�6% �#y�F}{��[��B�I�5@9�@�O�gLR)x6 þT<B�I�1�j���&��Ih�]2RB�" �~0���O�*� V��Y[�B�� f��1�c���&}����%}fB�	>��1��	ޗW��M���׍'s$C�	��=�v�tj�u��e��_�C�I>��l2u*ɛy�|}XDX
]B�	�E�.��F�$Q�Fe�3��6+# B�I�X�
�s��F�P�b�F�;�JB�	G? �r�H3�B��EZ"mMfB�	.yJ�Ќz��'R�Z��\�W�/D�$a�`�xB��#���<��$�-D���2����r�A?-Ш���k&T�H"�޲A���{0/��&ڐ�@"O>)C�ǎ;����n�&��"OD���C�P�fU��l�=	-��s�"O�y��感h�B��f�P�"O� ~�*SV�ma!R"��s"O�P��˵CD*]c3�U�f����"OJ�� ۢ�6u�cZ�>r���G"O�`Ҏ��sYa0��Co�<+"O~i��`Ā4�|ɐ�Cơ{Y����'��0�©�8��Y��.f����3D����/���8P�D�L P��N/D�\Adjɂ!�5���)�*Y�e�8D�$��D��.�b'��!�pi�**D�`��D�`�T��.
�>����!>�D �S�'t2(S5�A3F��Y��
�?��`��,�ݚd	�VXx���i:t��ن�MG���G��v���Sv�[<���ȓ?���IeOGDހm���x_����P4�F&Z�2���� �7\����-�t�{�j�"7�IыT��u�ȓ?p��!� ��­h�f��N�=��ğ��'�V���L�,bt�a��8t ����'�l�:!�T	\n�x��� �Z���'\�� P�j!py�bEM�x�R�I	�'��ŉ��W�h���́n�~���'R�3�) ����
G�k�h���'0���d��k���e�=b#إ��'-6�V�� [����3�˅[�2}b�����2J��¢��	o�y���=O�y��	�Yp6�Q'L�7,���iWo�B~�C�	=U(`��F.+b �k�Szc$B�I�A��;j2S��MxB��G@^C䉟dn�h؄E^nvd C`�"�8C�	+-���#�Ľj
��D_i�rC�	'.�Y�.M '~���\H[l���:?qaD�`��2f^�S]��gUg�<R׺H�f0hC-�1]gv �֤�i�<����}��Y�#`P��"9� g�i�<ɰB��8p �J�Vu��S��i�<y!57���aB,;�d!g��N�<qEO�fn:-K��(�D�e�_�<��h��^����B'.b��$���D�<1���Me��ac�؁�ti�f�Dw�<��\=I������5] �@�WJ�<����\���S^șˁa�<7�G?���f�C} ([R��\�<a`(�:[gd=P�3MY�<��ַ���g�?��-��T�<�5ɘ:`��3�"��@�f�M�<�@�򌤹`��`�(����G�<E�(�`lAoʬ>:���BD�<yU��c����f�%G� z�τ{�<Iw�a~�xh�-��T�Dy��eS�<!���6(���b�%)g�P3�z�<y�AB�q�ꬂ�nY#Rz`�Af�w�<1�$?+Z�0�W�S
� +�����:�xI���P�)i���3�j����-����)�zba��K<نȓ]H���P�D���Ǩ�#N\y�ȓ<��L�5"��%x��+D�B�r8�ȓm*�YuD
.SF��&�&�ȓVD�)�g�[�)����Ri�Y(Rq�ȓL��,��hkW���&���,�%�E{����=* ����*a���A#�M �y��R�)��0@��Ybԡ�RjQ��y�~��ن�"Wb�$뱀��y�R�Es�����\�Z2 �� E���yr�H!j_|�p�Z�_�29�F��y
� ��y C�Z5L�y�+��w��\�""O�]Y@+�ج�T,PoD��"O.$���u�r��S�:���"O^�BW�ۜip$��G�:�L�	f"Or8pD#��gRZ�1�H̵�R���"O�} SJ��s˺����Hy���:D�Ģ$���Mr`�y��T�,�!i7D��2��H�M��d@�@�*����6D��U���8����H>��ey�K�O0��><O��udE��b�)��	�Ą��p�͇ȓf,��k"�`("e!ue@�x�~��'>��'�T(��hM�x,�A�Dd=�'�����aC���#`R�48�B�'Y^�J���f.Q�cN)%؜Y�'�њ&b��V�#�O�j���'vN��dL�'fZ�)�
W1�6�	�'0����ѩ5z*���D!k'0�B�'t�����Y#Fn�@jG%�3>�i���'���Q̇�.XD�)�$o8@�'7��� Fxr[��Ϫe�b���'8!p,��;Y~hX�#���(�Q
�'���B�*ΪH��S�����O�x(%�PPF�"F@Ύz���b"OR���C��g��9�So\� ���"O�ԩD�>r��*���:�pH�2�	w�h92B�/o6p���Եu�vu�g�:D���/�39���c��im�ѣ��6D�xK�)�QW�������e:�6T��q'c��1�ҐZł�����'��ؘ��a01�"�1	.|���4D���f*�v<�����@>�7J<D�|A7i^�F!��ae"�:Wb����/��_���a�����QעĲT�����.D��.L�D�b���/�7(�ZY�co.D� �ч�����+M�N����E D�XQ�� �����6&�Iʇ�*<O���*��4+��t���+&,��pCCE�1m�C�I]֬�QB��5G�\,�B	v��C�$;���y�+O���]���D }��C䉩5�^|i��1��R��R|C䉥g]`�[s��.ڀ}@%�XWZC�ɇM��I�a)P�v�\�"Gt��C�I�C� �#�PN�l�BÚ�c&B�ɂW�x�IӦ�.iϴD"@*Z��B�I6
AX���;#!r$�Pbע"�C�	�6��	���b88��W/��B�ɔX�����#O�F�҅��x�dB�,:�9P�R(l�88z�"��H�JB�ɠ4`�)�Ղq*�!���7�B�	�)��قrm��$F`�u��p.B�9�4PF�[)�����J[�C�ɡg�r
�= �L�`�oi�C�	?:b� �ɕ?:��=!%-.���d�	��@E�4��*O�u ���u�D-S�O��yR��k�(�3D��i���l�yE�
$-����d��� �Ҷ�yR�˦?!�]�EI�Zc`�k7N���y�R�R��IG��'�V��V*�y�Bߊ�z=#���&i~(
��"�y�lѿ@$���"���>���_��ybō)�DPr�R��% �6Q�΍��)���eѮG�pH� ���[�<��ˎ��ܨ�V�|Z�1e/S[�<�c��T�^,�#h��*S���B��S�<� :i�br�a���jg@��	i>a�cnO�\_J���՝��tc�b3D��цC�5v�Llr�ˀ4+����&1D��( $�QQe�ڇ4z�2j/D��� �җl!^|�3DX�O�v��֧-D��Z'��X�,P�2)�x-3r�*D�<��KD�<-]H�/�a�"%��M(D�8b!�Ix�!"�-?%�M@�.(D��v�� MȻ���<v���K��+D�H���׽=ǎ�s7�T"�.�n-D�|�혭3x4'. �l�
r'-D�$b�	Y
)��Q
��t:.�6j+D��I$�aQ�A2���l�.E�h*D�ʠnI�R#�ȩѭ��F��<D����!�B#~ыv τz�: ��H.D������.h�̵��l��u��J��y�i�3c�t����ٛrN�4���y©OR�|� J=��e�c�B��y�LI"��݊cJǁJ�� ���4�y�Zy
Rm 99�HA!�G"�y�� �l�T�c���'x0P���y��Qܜ�*I̖!I"��y�@M81�\���K� J�-Y��y�挋i�L�g}i"41�J.�y2S�.��y�DX�D���(��Ͻ�yBC��;� ���;E�(2Ї�yR$L�9襤��ȁB��pYVl�y��L:g��eX���'t4=��� ��y���91L�1b�T�&��y�U�
��y��$q2��B���[X%����y2.X��9 ����&-��,��y��R��3v葎@L�Q�Eo�5�y�A6h�2�']�>���
5���yR�X� N(Y�p�A�L;j͑S�1�y�	�d��kwɒ�D�`�s�5�y�eNИ�C`��5���NE��yrL�	|vT�� ��`ix;"�3�yR�ܬt���Q��c��Tc��]�y"��Tbx����c������yB��N~��Y�腏\�( �`c���yRQ�l��9@��jt����C��y"� 5����C�x%�%	`Z��yr�۪wA�I�����&4�tX�)���y�Y q|���V�i]�ǌQ��yB��H��'�G+[:�e���D��ybM �oL�T+�CEN� �HW��yb��\L�vEH8\����N5^oB��9wJԲq��<����K;�B�ɏ
7�%X�" �d��Y�MI=j�\B�	�4 x��Ȗv��� #
��<�"B�3�<�W��`���e�
=�B䉧*zz�Af�؄,���¦t��C�&e�����,n��4�DA_0�|B�ɘO��|�b��R~���Rꙶb�PB䉳pz^1��'�(�qԞF�C�0S��fǖ�,M���U�A�C�ɏi�)kQdڜm7�� ���TyvC��3'��+p舕)ʴ� &��lC�	�P���I&���\X�#���C�	�7 t9@�(S#��hr�T���C�:Ye$҂�Q�7�0��")��E��C�	;4<��`O����q�N�C�'���\�ST����)�xC䉡}�� k�Km����q"`C�)� ����bB�dW|`��F/�\�1�"O>��D'�v?v�K ��)s;��"O�����;T���K�V\�!�"Od=bF�!F���L�>GHqrq"O^\���H�,!A3"N�MA���"Of���lC4qpE{���Ao0D�� #-�0>�� �cA�X���Q�+D�h�uoE����rZ)>����)D��R�玣<Ԕ8���!��Ң�<D�� ��D=FJ�9r��_+U0��-D�@��H/b���R臬>޾���?D�h�D`^@{��y�G��G����2D�<��Gҟ�mm���=v��I�@�0D�x*C�M�Rt��a�^Fp=Z�,-D�����^PȀ�(ݖdY0�J�O+D�d�����6_�IY�#=;6�!I�*D�P�����N%�Y��̃DHn�p7O'D��1����j����A

6'�NU�T�$D�0J½p�F����p ���!D�PJ4f^w�1�CM$+�@b�$ D�����>�x�Eά)�x�0)*D�d��!��u�ɋV4���<D�� �/ɴmk�;��J�~�؝�c9D��V
C_�f�`�@ɏm���cgN6D�H(�t9n@�4�*�Ƭ�0�?D�@jG�R� 'L��uA�0�h�5�"D���%�&#2�y8&���,�N�� �!D���!�*n���w(i���ñG?D�x5Kʜv��x�j�-��jq�>D��t�;(�� JDT�u�J�2p�;D��f �s , �GҺ�,A�#;D�0�o�ED��:r��a�D�y��+D���`��/A<��҆w7.��U?D��r-B�gi���CdϖH|8��K:D�4JVg�.b�Za�tH�&�r� ��6D��3W��Gk�s�メ,z����6D����F�Un�pk�@��Q!�}�W�/D�H�&�cb�S�h5X���8DE+D�,�fa��e��Q��%I��y�b5D��`g/�?������(��=2T�2D�0�g��.w���'��B ��s#2D�tB�Ҍ��ԈU��
3��lej0D� �����_Z�xc�T_�>��/,D�0 @d�N�x#Q�TWq�e(D� �c��0�><X�턖j���!�9D�ٶĖ�
iV�(Fˁ� +��y����*�,��͔�$P蠡�#�y��6%|Ac��%<�܋@i�%�y���T�|����n$Ӕ ��y"+�#=�ԕH��'��a-�*�yb�(,��p�f��ն���F��y�)Y�4hD'��$yb��Pi>�y�&�����N�����.��yb�ɪ�����n�,ːq�A���yR��:\����v ��,�lk�i�y����U+�P��
�)��M�2�Q�y"�I;&�4ۡO��*J���-N�yr

5�1d���n���c]��ynG�)���J��^��h;B-���y2.��${�蒊N����@��y�-V�>�f�Kp𔙐LF��yrℱMz	[t%QFC&�!Q��y�`�2P��#S7r�D��D���yb�{��L�B�ި!�j8D��5�y
� F|�p��9/�(��d"ƂfX��E"Op�� H<�px���'d l��"O�8��K �J�p@��	'RC5"O,-jp��(s��D��#�
&⬘��"O���j\FpڅʃA�^y�"OP|+��OJV59�+�9��i�F"O4�P�C.�,Ȩ"�ޒs��dj�"O4����32�DO�?<r"O�œ���YZv`&/&:,u@�"O�x���B5g����R��0H��C�"O�p@ˈ�ZD$Kw�
�i]�1�2"O��с�K�j��$�%��~����"O"��w�T21�p��5�l��"Ov)P�"�Kw�eH��ٜ��h1F"O��4�Ó`���{�	�<
��	�"O(ձ� R�x4��
Y�(�����"OD@D@��!�y�����z�&媁"O�U��NB�V@V��hܬ=��T��"Ol �'��:^O������7����@"O̅q���9Qm����IN�r0��"O�l`��:�~�O��1��1"O6����=�H��`� g{��0"O"5�a�ĸTE��xV �#{f���"O�q��Ѥ/UA���M"EjD��a"Ot�ce��Vs�$�b�f�$��"O�!R�b��^HΥ+�DW5Q�4��u"OZ�!6��<�0�Æcݘ^ج=�F"O� �1��'3xАі��.�ZR�"O�DAa��z�(�)u�M�W�<4Ӡ"O���m��d��8�g���Ey�"O�am�L��w�J}�(�D"O�sâ۞Hg$���f֋9�Xi*�"O�� 6m���i���`� D�""O��[�I:-6A(r�V�KQ���u"O�=("H��i��hK��	�"O |
V��&5ܸ��3Q���Ѐ"O��ɡ脀C6�%�5=ΰtR�"Oؙ3��I�Gz�=j�lF-[�<�"O�9
6AI2�ȝ��,ls4"O0����\�&�� Br+R5d��Q�"OhT�$D��:�r�+0	]6o�����"OP!��� 7=; �ec���"O���p*n�1$ �)*H��S�"O(�0%+�E�8�1NI�R[,��"O:����(fr�s��^<	�v��"O��CP�J�3b^�0lȹ9�n�� "O0@K��),J)�U�
[Oc�"O�xd&F�5��� 6�586�5"OLx��M4B�Z��⋧q`�Ђ"O2 �7 0GrTI�У_h$�J�"O���f�	**�!C៞j<�)�"O��`F�5�Yz� \8c̀��"OȪC��D.�m��OF>V��(	d"O�!�a�ߩ}�lȦn���vu��"O���1���ؓ$?��qu"Oƽဝ���,`��Z!�Y�"O�}9���\иLKv�LB�v�S2"O��;����d(fd��d�$	�"OdIs��_��n�*���.`��"Ojxp��� �$���`�%z��3"O�qSHS:R`M	�-Q:*�t���"OH���^ ,N.]�V��ᬈB2"O*�06�
dGD}�R�L�Hе"O|�Ãm��CW��cb�L�`� �:3"O� �y�V(�{=��z�i��l�� ��"O�T:w!��7�5 P����"O�M#�υ'>Ґ��W�^�F.�0�Igy���C����$%hҼ� ̲ o!�$A!���8�Y{X^m���;A[!�dH�̛�b 	t��H��I�!�C�i�b= 
H�&k�pä(T7:R!�DW�|�Z�G��)0F��vi]"2�!�[>����ФR )9x䛴��Xk!�d�Du�dkA��21LD92�2.X!�S�=}`a ���wj�R��W<�C��+U�t�`F�	e�܀���N���J�o#�S��?Qc�
juh=�g,����	q�8%�����ti��+���)k\���4�D���}��'k���h�Q�nG<���ǀ��tF{r�IO�ԡ�;�$<J6ċ�~a(��$���y�L*L,p�@�(��(f�(�ƭ<��O
� �4I�F�>Q�� V8'�d�g�w0J ��('D����`X�C�p��#�eBhX$�c�����'�ў���K�E�� �+� <��L D�,��.F2�4�ră]`r�>}�Ë� ���%�/��k��i��	Y���"C�W��)��@�i9���d��?	��VQ����/|{��u�'�M��'�ў"}��ſ]a��Pt�ץy��� ���M��#��~��ʭ]?���$;:̈櫔�!�D�!'���b�1KM��Ŕ����i����u#�<��Z?c��s��Uˊ5EW򘛖Ä!7��S��'=�OP�0��W�/�p�@&.ž���_쓧y���O��т��F*b[�$S%F�Q���(O�;���H_|<�T�x7�"Ov����	��n~ � aU�x��:�S�'E~5�
G�i�Re�S)8{p-��1GZ����S��:���<���=���$�<Rg�'L�dra͟�B���4�PpH<�u�P$^�z�)F#�$-�r����X�tzC㉂t��^��(�(H�U鰹��"O*���E�"G����gB����"��i=��б���~�|nZ!?���@��Kz���o�nVBB䉛I��)qPA#^b�c��Y�듥hO�>��@I�^0���-T)0>�a�$>D�\�g�m�q"e��+	Ҥ[S 7D�����k��l� n4����*D�H�C�	�!xX�+1�&G�b�3��'D��"BiJ�x7LA��+��R�A�'D�<!����˔�M�\\yP�(?������H����A�E��>5�@��L�	_��P(&و0p2`�S��(-�b�Rw�6D�d3��qڀ0�dڒ�.�QgH3D�tYDX�,L�1�FD8�E0,O��<Qqe0g��cu	,�2�q�<�t&�k3��I5*Eqf�I#E��<)�y�U�"~�Q���M���AB�	�"��ɩw�Qo�<�!gňz��$놮ۮxN�d9TO��<�Oc��G{�(H+kT=xB [�M���UoO�Ә'����ɂ�M`���2C���3㟇K�:��D-}B���C��ܰ�#^Ѣ2���dh�R�?�K<A��1U��ċRiW�g�R��g��b�<�T��-B�+�I��W��U,U�<I� �J�n0js$ӈs��@ V!�L�'Nў�'xy̐ 
L"���Aƥ�%!����~k(� �e�4.����/ӕ[�>�ȓC��%� *b\ �&нi_��ēR����Vi�nU�gc9Q����"�<	�'/����$$�`6(�&W61Y��� b�%m]*SI����Ms���C�i�ў"~nڞeR�B��(h
dQ"2	T�<R➰E{J~���Ð'I���� �pQ�G:�y�c�78�4��vg��,��B��y�ѝ�RP�SHR�QN��q"Ѳ�yR�� Ԃ�b�/t}^a�pʂ�0?�/O���B�&p�ʽy�&Y���:�"O(`�)Ն:�`p0A� �.��((�"O�8I�޷5p�H��J>Y�𥫔"O6�����T�D����
eK�eC����BJ�3�2� [+.]�1���;�yr��'���Fg�* ��5����7�y�R3])<�2�hC>�M�-Ot�O?7�Ө�~�#���D4M����!�!�DĦuL�����8b�`���0g�!�I!�q!t��/Ml0�wc~�k�'+��dQ�gD]��*�-0�5���3O\L��m׹e�uK���X��-`r"Oe;���z�Q����I���"O�tRg��9-=b0�0�W��ք�P"O���'C^�moR}��A�}�2��"O��+d'.A^�Tp�b\�zv4�4"O���HD\}��u~ڔ�����Γ��'��	��lŕ�#d�Q$`lek�:O����ؽw!Th�fb�L���Ť�5d�!�Č�H�x���H5>�^Y�V��:/�!��l��h�����jV��� oE�3�QJ��ԟ "=A�m��hT�܂C�ܰ;P=����`�<�2�31-"P'P'����o�X�<���s�����
9�<yS ��y~�|��Ӟ�2�(��ev�@k�@��C�Ih�]�t@߸E��Ĉְ^�tC�	XF�*d�%Oء��&�:W�^C�I;Y�D��%�"D���"��dB䉯Rg�jw!X�>���`nD��|C�n^V���!W������I�s�:�$��I�};4� tC�i�=�.�6-��=����JA��ݻ$�bM^ �N�h���'����b(&a҂l!n�V,����'�t���'U�W`�a��p��	:���~���
[�ꀥ�j%��Q��
�ē�?q(O0ʓ��Ӻ�#-�?n����
/a�Vq���I�<���fP ���#3���p�-A�<Q��Ӳ]�Ƙ�`c��_Ȗ}P�-I~}���K�	^?)Ǌ@�=N:|B��*��x��
_y�<���s6�8�jK�XDM8'�x�<��*�81�E�#7�v�xteAr�<�͘�FXv	A���xL�|ȡ�{}]�T��0<�4ǖ@��B ��@8Pd)�Sx���BY)#�Q1Gϕ#*]�) E�W��y"`�"V,���&>fA4�U#��<	��dƽ�{��@
tH�t�c!9!�$TS��S�׼D_~��vdB�3��&��J�V?E�ܴ�)���?��J���d>RQ�ȓ]>�=�a�ڇ`K��B"͈�x�V�$����C���'U[*��uD�9d������.����� �Z������gϟF��T��?���T��>B�b(r�Κ��ȓA;���ɏ�r9(��S?�)�ȓ~���SC�5s��)0���w�nP�ȓ7<�`��X�gNDi�@!�>�b���
�UX��Ƈd�mb����w��	��iNd�f�u�6���ؑ����D��(���;_5���r�؆�S�? �tk�
M��Y�(^7V�����"Om��99b.1��g�*�,H�"O��X���u��q)���#�N�`E"Oa@e��D\����b�����"OV�B�'\И�卉�(��"O`!��5WY� ��BH�)�(2"O��0&�.uj�(�g�QT�r#"O h��=M��rƅ
K"M��"O�I��&�;�Z0寁#rYu"O*���+��4��g
�3>n�r "OVd�0�ʡ/(�P�CΓ�cD��1�"Od� ��?6`� �l�8W��P"ON�0��d�>���iP���j"O�����п�0��f�M���zE"OݺL�n3@rfE�B�̓S!�ӧjN�e���ϼ!ۮ\Ӓ"�?V�!��Qj� ��`�ZM�RaH`��򤗡D��1�5M�i�(�2#O.�y��K�0����	��ag�y����yR%\;6�$�`8_ ��hr���y�BU�,2�A���b���A��y�B� Z �2��H*D<������y"���0�d�<�>�@����y�ކhi���ݔ.�0�(�$�y Y�U�dJ��G���xJ�J���y2�M�I����v���f�I��y��O%=	v�H� ��0z����y����Ԙ�%~�ɢ���y��U ؜4�c ��ak�^/�y��C,�`���b�?�"��ˁ�y�K@89hT�%�E�[<Hu%E��y���M�v}C�H�C �	Rg�	�yB��0uo�7	PC����y�)�4.�&4��I�!��5-���y��C�e&��D]�"{fuq��!�y��ۅ7��` ��	��B䜌�PyR�Tt�t��"�ѣ,�ju8�K�\�<��$��(����S�!'xi��Ef�<1�鈖e�*Aa�<bX�z��S]�<�4IV�U�v�C7��\`X��dCZ�<�!Ń$M�6�r�m�>��8��W�<a�h~	����BY ЋF��M�<Ѥ���q>@��I��5���-�B�<YV)GNP��U�M�@�V�k��Jr�<�FbOe=&�9�ą7䐨3w�]a�<$hDk�A�!@ B&q�ׇ�P�<1�`?x�썸R#�f��e�.�y��H��DkW�],X/(�P��<�y�A�2F��V �.�J�D�	�yr疕Gu8�q@�.��!Y�6�y��U�h�Y� N�$����m���y���?�,8��OK|,q��
�y£���,	�˞0
�h���H��y�ޜ,�H	Q�ܼ�h)�&G�y��U�l)@mA�kS'��a����y"�R=)j����&[k� ��ˇ�y�I�6wxx����Z'z�@h���
��(O�4��	��wxz�������O��K�C�
^Gri��Ʌ'S��hy
�'::K@*�I9�;F��>=�Ä�S1�T=��C1b��d����h��$K�o�B,"�Q�(A@����n�!�$�+7�LT2U* YS�)�b��J��r�D�Q��u%�l,|����ޢ>� �T>V�jYc�aCG�5�A �P��h��E� @Jb0t��=P��hY5 � ꖜ�f�Q��h�'M�V� `��'�v������ʙB@��3�H$Ɉ{R��y#�D�4��u,�0���1C���'�d� h�*G�v�L�3#���{w)r!�d��-�z� �ԽC�X�daM�8���֋6�F�s�. Iz0�Do���u⌰S��Kp��t�4�8M��V��~����y�#�'� �c�@i~���
$ ܓ�M0g�5h��%����"���< � !0����A�	,��A-��c�02�[[?�e�΢=�ge�b�,}�נ�`��c�*q��� ^W���pU�d`Ƭ�� | ���!J���l��o4�1��H?o�hI�$鍲*ǌ�6 �q^����M֕L��,G|�*�!��h�ƈJ�=Y��'�����R�ζh���ã���zI&m�@��"��X�6(K�8Q��7d5��82A�Z,5���sg��7{%l�8�$���j�)�;�p>�ˍ'�!b�J�j�aK0!Ng"H��� C�Z(�fh����t���!D��n�q{0�LLb,h�A�MĘ1���19����!D8��� �F��k�;ra�Xq���[��б�%��/P��err�A"7�¡���?[`�����&'�
S�;o���e&\-U��A"�(� 2����ܥaP$���D���*�J��-A�z��lI6� ��t�� Z�:���[���'eZ
��$$��fl�{V��=dL�8���иIIH%Y��;e�����]�����Ԓdh��>i�GR��i4U������O
�0pP�`E��7C@�RQ�Y���G�
Q��IC��'��ͨA��2q\��p΍u��Q�tkY?;��@��̺��pWk�I����s!]L�LHwf�)C�(m�k\W�]9�$B� ~��͒���EaU`^�BL"��*D�<y١�R	�aA4�/'s`�B4m�4�VYQPd���k��cIGB%8:��['�w��m�:P]D��ǫ�<<����u�Qwl΁p��x�����
�[L =p�F]
PP\��g�ξ;����dQ�sfر(e%�{���x�O�I��e�Cl;�8b�O�
W˕9�l\)d,S=��Q����w�XY�#-��D�4��Q��5���y2�Vt�6�Ҏ�D�x����'�re0�K�",��8$�����9B)�p�"%&����b�zP$�T�Ckh�j�mT�J��f���@NTyI$&wٰ��&}{�<�u���&��82S�+l��I���Z{$fD�ᎇ�3���bJ[]�����b�%�j�hÊH�%��ٍ�d|(Ή0�&�,��+��S��G�a�����?�,�2u �cw��#+f���/��
�F�r�O#��ULI>�V��@)	�v���&IџYƖ�>�cϕ���|	'�J#n������R7��rg
�LFШ[��;mR<	5#O�q��5���Q@����P7��zG�LF޴cŁE9	fJY�#�,v� `HPN�}NM� l��A�T(�'�����q�L�bN� ��y!�l��Xw�$�]��D�]���hcB��U�R]H�d�n(Z��\�2-00:��bC�}�BŢX���@B!P�Hi�O����A?Z�A��V�~���k[*]u����ϲ�e��~�����gA>]�9P�L�+W�b�����^qlt�0,�+���i�ꄵkl�gJ�������[0�Xp���y�,ܿ/���%�ਠ��&�bi	��5l�H�Z��
=�� �	'�}��N/Bg����nُ �ju1��еl�N�*���=��xbI׹8��쫳�&P�"a�;$�^����itr������Z ��'���7��P�|Han�;R��L����V�xL�O�$J& Q��ɋLv�Ke���&h��Bч9̜���G9P�b@�q/�d�'T�Ap�@� �\��奃�48h�Q�Db��W�
��H8P�P�]��ȥT?xm�`NM�|�'��-b����$����Ku��������EH�ҩy���q��O�/f����݆(���	��v�����_.��Iq�SDR���c��e"p4�ht��>=�8��`�R��	�"(��Q����d��Z��"h%�,2w��) ��"���T�",��bL"rUܩbp(�1��!A]l]k�&�.�Z)$α<qTͅ]�l��	T�VT���$("V�5��	���J�r�!E	HL�"�ݓ^�d�0��*T@��Đ�%^��e�s�8�ӨR<p��p��. ���(�.3�:�S'nC���R_�,����9g1q+��<j"�ڔ��9�L���.�U�lX����&Z��T�����)�v�I5,��*�FY�u�=�\���N�O`x�B�ԥ_��t�!F<��4�h�V���{b��Nd0�'��A�Ǥ֋y� �P�P�E����
_�{N�S�}��Ay�lD�\�ʡ��!��E���A�\ĚUL\+��Ă=MǶ*F����թHu���'2�}��� �*���K�x�Z�hb�=R�A��S<)��8�哂x�$��23�$�(�*iJ���1�.扃;�ҵ���Y3t$a9��1;��È\�oG�![g�>�4$G�<����T$]|1@�IJFz\��˩b3Rmr�A��T�'<���V#�$\x1P/��LI`t�lП;���V��
���X�K��1��^.hH����"�c��1 ��&�)���R�lH(f�I�79�x�@�K���UB��ǆf��(i�CK�ѰT�����?A�lȐ2=�p� �
���y5�f�Ceo���	�BLA+�"��!J�U��'5VM�d��L��9�2��'U�(5���u�2)u�jm�XZxp���:�v	!��c�ld��ĄQ"����IW�p4:�-F�\Ph`�2�r#A f�U8�g�b�,��2㒝_z�Xv�QyH]phӫ)?4�%��gA��Ԇc�.�'Ɉ(���\��!2�C���rB �'DD�E�r���#�,EZ�A�	i���{�(��96��rt�%}�(\�By�a�`;�����,��5"��x� �G#ÃZ��&��8E�����@�r28��O��Rd'�y6m��M�)�����
�X�R�2�'�mبݡ����D�O�]�#�@y*x���S)P,�b/�����Հ_*�V��썛$�0��@�:^�-��˕.���i������(�X�2�L͚&�4�)�EXz�B$3�[/o�&���#	]��\ےm���Ɛ>-� ��o݊a,Yӕ͘��M�GDcC,�Ї��5�N�C��dJb�S�w��Ka�A#Y$��(T*�''B(��ǚ?����NL�\��Y���[$�}��ꕽ&V�2�G�zH�!���)�F�+B�.�v������R�q��OP�!+f�)�oZ�n���J1��~r8��Aʆ���	��+��x��g>�h��� m���
�y��Z�C	T�A��"B8�U�rL��KB:�Q�`�ئ�Rd����9x��T�( 7�����1OR���wi��9��`���m3��oשo�D�t�L4S�}E~¦��~�ZMK@�[�&m��"mJ�OTx�PqH�?z�8U����x� \�ĥƎ��ۗҗoքɺ7��4IY`� �H�|؛�i����O8\���a�P�'B�+Z�0ŸO<��D#S�U�o	v���h``M�n�R��p���01�yv�!+���<�IH"4����Wg�2C	.<3�C$�<1Y3	�yu�)#�����sӀپ`�*�§aϰ�`$ң�12��[F�(y� ��l�9QT �X��6�վ��C�.%����,�a�$�e2H/��e�F�	�&�A��զm�֧��U��O��,���!��E�? .d!�`&WrxJ@A�H���;Cr7��Ht��	��y,M�2@�,I�<���� �� ^
,�%�K�d�أ���gY�<�� ]7��q&��<Y�5&��ifN
=Q�:�eN!RQPVv|�8Vzx���	��(h1�GF�f�nH���[�ۘ'�hX���Z�_i�|��:A��I��s.�y�Wb�0J��u&�|�g�1I��i�c�ˋ��P75/�%�d�ݦ8E�����
��k�� '�]����#�� %�I�@�^!ļ��N�:��O�d�H�ƚ���x���.*���f��
&
d���ɚ	"�ɡ2�Ij�j�`��F��iE�8��.R�ܤ@EH�<2.�@"������rL�Q���"x�ftI��9�3}�b65�]�!�J��Ԡ��I�Q,�u{#�Ԥ���N����X�B�64�Q�a�X���dM�r˂�N�P)���]crl�AW*�*�<P���1*�9�&��sL�͹�Ɲ�\غ���hfR9 �j�8��īO�EQ�d�6�ՂP�6��N>���R�<���B�M��d��\��hjs�L�s�옴�N[�8Ѝ���Ya>����~|\���ͧ,O��3q���%J� �L4�`����<�2DH��*ĺ�N�"��`���)C񟆀�& �*�>��4"�12'�='3O"�z�KS;H&�3�\p0������:��$�i��]ŊcG!+,���o��C=�ـ�l�sB��Ђ�c��xxTc�]ǎkW�O.�Op�4'��r���і��X�f�RE�h�h�B���� Ux�*��E5�&��X� jt��&P"6L|��O`�-A �!Xm �<��fP� 3Fh˱�M&pV�CW�iEl� "��z���hO�§�,ޘ�"*I>����$��%1��[���)[B��Rm���D�<� /Ĥ3��cf'�(Y@b��C��'Y�X,h)��7X�]�'ȹ<q�@U��\��c~���h�6M�d�ΈHP�N�^d�����D���F �*�����E$/s�����0=!R��AB�#5�_�X�Ā��'���y�U�Pe�ᠵ/�~��"��ER�uF?�I'}�vps�.
T�;$�	�np��I�����Ag��d��K�#�4�cf܄�I9�ךr��� ��(�E�l�2 �S�Q�Q8��
v���� �Qzd�G~��_ڜ�����c����+�.���W�RP�r�a�@ƾ�*2,^F̝��Z-@��p��
��^]��K�!�	y5��J3�bU�i�'<X��AM�]hf��M
-)tƅ�@��?��%&�/ܮ��Rg�R۲�5�z �7nת��Δ7/6��9��x�x����'^dݱc�![��6������W�_=�,�UAP��(};�N��Vp����(�4��b��ю�l5愘'�P���I@�<4�ΩJ!�ŚG�2S%n^
RP�s+^�q���X�s�B��0�ޚv���!�G�>5.H��J2P(���Q���=a֣�gprpȦ�էb�dP�OBb7b�Hi�z��"�&��U����2� Y.p&S.4���i�͜��~`�9a��U�$�i���.I�R�0 ���:�F��)�=5�,c�jBz����Dj�0�{�x=��O�MǊ�z��»8�WWJ�l��L���,">qW�����1��%T!�ɰ�l�yX\ah4�ڗ(}��]X��0�G��B�i�A��(Dk��+Ƨ��%gx��B]�X��#>��7t��*O`����0�|]�q%θGl����^��t�S戇��ȩIƬ�5�
��:�4*�#��q�|j��R��?�C�C!A4v5zG� g?YłY�W5�Q+9_4!�0	۝W*�Ձ�K7I�,zvA��x� }y���\�/�|l�c�m��AA��"�ɷ_Ųݱ¬� ����ȼ/�t�%��)�b��(OyҐ�2�L6]��չ��=���M�~y��M�Y��@Y{0�rU��!4S P�Tk�7.i��G3�]� ms4F��h�X2/�A��Z���>�3wǇ�!��p��D�ޕT�����م�I�C`-)Ą(H���%D�"=9�� ��42N����RH�O�RKގ&�!��֫r��婳��5��`
�ӊ
����:ob���H��6�A�hٸe����ND�C��QlZ&5�	S'�V�Qڙh�h�3	&mB���p�r9r���5���4I<D�6���-@�$��J�̹Ј}��Ҹp& ���6?���V�D�[;:��&�{��Ez�- �A����ú\o��'��X�/��_<���� �(/f}��HϽ{���qpEߝY@���4��ȣ��	<x���A��
]���샒��m�6��J���r��.<�2<	��Fx����[�Ɖ8���l6��'#8�	�r�ps蛵$8�!����|x�柰yㄨQ�X�F���K��h>@s��s؞��A�%b�*f)P����dJHK
�E�nD�~��hP%.^�J���t�]4�L��w	JR���ӏJ�eS1΅
x��L ]�v��]sv R��85�I'd����'l���뗋�b��虓6��F�z�z�@�V'.0�P��CU�B�`�[�I6^�T}���
�z2F���;V��E���%+:�`�7�F��e�&� �1��+��D
�B�A$�^$kJ� �ʑ��y"	ԟE��U��d�4��C�E��N�Q�*ߣ�����Ȉ7E�� @�'f�J�@l^�	d��l4�O2A
�l�'w��	QDX/w��-�S�iC��7�88+�<�e��cyD�D�|"N�dw��ٻM�|#�k_/��D1���,7<���
��n��QL�'vZX)�`J&T��`Q��;<���B"�W�xbݴ,J�`R�'P� Q\��r�O����"��st�Y�%�ߝ���R?���!K���90�%�\���Ò?��Hy��@�]�j�9`߯%
TebRמV@��ʅᆘ��2@ԧ$Vz�)��/Zx�i����(O �*
�J^~R���Q�̫��'��@���`���^LA���ʭD�d�p�J�{�<T�� ՚T���0���!r(�%�A�@���L�'$,���'8M�C�_D;(�FHY��v�x�?v��i�c�b���y�id0A�g�@2<�@�H��r�̧�� �1����,BP��-S�zV"O98���v8M� DC.Y���7�P� ����A�S%C.��BE��{�1�O�"i �L.B�ţ�w5r����ʙE��Q�[�/����v;���u+��q���qD�NA�!Q���_ĄMc��B5�䞒$ހ��5�X�t�����d�a�(=1��Ơ'��ћ�$��-Bџ�Ԅ����[wʒ-盦A0�2 �Ѩ�O�����L�f�@׈C����D�'�����ԗR0�[����6!��{�/B�i��T�S]N�0��'H&���.\�3=zk��ݧR�n��ȓaz�
�0�i��V-f���I0��S�	�f���A ���C. ��\�r��rO�YA&�Y1!򄜵W��`T`��&XX���j3!���#h	��W�r���sEa�!�䉆 ��(���F�W49YwN�"P!�dՔK	�,����	!�h 0/3!�D9=�� �N��L�ʢܗ?�!�D�4��x�3a�$Ԟ�"eW�EY!�d�)i��t�u�B�$i*��r�!�d��,W`�ІE?��M#���`�!�D��T�eg�Y.��hT9>z!��_2�i���BC`D��f�<�!�D$���i�B��&M�*���Q�!�"~>�P�k@5: ZA� 8��	�'�r@���ɽ/yJ�� �Z'jst��	�'Ϫ,�Ƌ�Y2��@KP	k?�q��'����䊏Z�! t/'7V��y
�'-��Ӗ�Z��Z<�s�Ћ?����'0.-�w#�7#Iq#i��<]\�k�'P�P�߽z~؀Ib����A�'�<us��r��1;v%����A �'�(;'2E�����	�.A"�'����ǔY'��J�6L��'�
�#��ǃ3�ơr���Phj��'��	��£*>)��@0_���
�'���E����8���ȰL���
�'B�(�C�
;��1�1Q���'2�U���V.O����!��|��%
�'��]"1��ioH)q[iDݩ	�'�z�N	3^$i�0OT�~��I
�'=\���N�<�<�GoQ�v"���	�'��i����W}p��樐�GG�H��'�F���A��V8�B6 \,5�v���'Ɔ��B���x `t� 1T�
�'�؝�3��S l�	H�7#��R
�'/�I���v����7@���'��A�j��M�r�)��A��'�����Q'Һ�(B��/����'�L!3��%�p-:�j�>X!���	�'��aQd8Т�6�ti��'| (��5��X�@�Ϩ[�����'��9� g�$0WRI dF%cP���'�NE:E �y�hm�G$��D��'��0q��5
�hMSG!ߩaw$���'w���o�gL�I!b�t�4���'��81"�3�q�5/�5`�,��'H�;��tM$�2�
!z�}�'���Q�e	�<Jt�Ɨ����'ײp+�@�'3n�K��(�ѱ
�'٘�Rǯ��VX='�I �!�	�'�4�Q� �)o]�@�ٗ)�0d
�'N��Vm�/.�JM��W�##���'���7$+`��i@��2j�򄆁a���7Y+b��a���C�#B�j2ݏ��ܸm��y���E����C�� f�|l�rϑZ�z<BD�?=v�x�*��6�g?i3l� 2�l ��b�LUr\��d�<� ơ��k���
��GO\��Q��:M�P�1��z�!ٔ%Z�w��n3�1m@��V/	����"�Zq8����I�|~�\���+g̠1q��2T��١��)�~X8���m2�EϘ�a~�&�'����@�F�JI��4��'�"��#@3�,�x7�_2�(�*�OB�Ʉ,��} hրnr�X����a.��r�?��kBoO9O����/<�P�����"�⼣�
YU����)? ��;=�8�V'Ծ1�>�ݨ;睙7+ZX1#)@/t|BU&G�dR6��$��T���O�xR�#@�w�V�x7+I9(4+�g�&%9P!ǎ�p���q��37r�tz�#�r�N�(�+;#,5{�'����ğ�-w���$!١�p� K>�a!�v��O�>�#��'�Q(T���x��͓#M zi��$T?v�~mh7Η=��,��FMAF�CG/ud�h��-�B�'���b�G��b��� ��Y��B���-e|`��da�R�C�Uqc���D��Q3�O,}`%yԠ�x1Z� 4̵1�d͢"�%�6a�D
A�T��	�*r=�fOɊt,�]U(��>���J��0n��� 7"�7U���(��$-~!�FO		s#�yC����<���b⢗�k��]��IV "5&�8�bёr�����'�Ĩ��AO�0G���<A��V:6x�-Z�es�p3���p^j�+�`�-HҢ�{��5��A��;2l�´m�az�9��٘�?�rA� +���BրI���S�W~��ac*U�� �;T�H� ��O�%P ӥ����D|�r�#�:r�f���$
~<�'��B=|�+�+ƪ}��e�p@�5v�2�ǻs�`b��Z��QuFp��^��jtBO*Pb�!��d�5ˏ!D!��
�W�R}V40B�ܴ\��$:��N�Pjy	�$ƽ(�X)R$ذc��Pc"F&Gv����#F�+/O�<�c^4x�"�;�e�"Xĺ�$õ/:�Q��	ºV. ���Z�tJ$h�R��7�(�;�� _ͮ�1G�õ.5�}�'���d���p!٣�B�eõ+�(�?q��`�j�ruˉ�	Фx���]T0��)H������`�6�&��5��=���;p/���,qcI��_T�S)�������`�3�>�ɥ���4SB!������!b *x���'!~�{D ������
�#��>@P���?l��.�FM�A��r,Ec�LI�0�<��U����Aw�ƀ�X�蒓(�\y���p<a3A�xBHo�Y��G	L!�W�߈*U��@'ΧwZ�s�'���eK�������|��*���<[�����N�ZY˷	�$W�H�@�#	�4ٱ��7x��<
��] !� �]�'�Ha��A\���0J�<u�]�BE]�ޕ��N�!Q�$�W��._�1Xw�p�/
�na�'Ύ�oY��;���8t5t=`�)\��~Ě�;J����As�'�Ā�v��gA�5A�,� ���G�R/��A�(lG`}��FE�l��B���dצOoL�9LF;U& ��1�ΨmBl]�t&D��5�Ծ�$�gJ��!��w�4�<�.L�4�8E�g`�F�1�,a���^�L�����
A�F8C#)&��X��/M s�H�(�00�|�	R�H��,R@��B�R+�7}�E��Y�v-	v�G:N������uR>H�e��ep|6���}���f�O�|�jb�O�p�ju����l�x��k�+�H�§DF�Wvf����T�S�Ε2�-yBp�GLBy(�'�Xق$A�I9S#���§^���  �W�;��}*'D��+w�Q�1J��d��c_&pF����'�'��(`�W�:��Ur�$;/�esbI�^���(GK�q��E����&����P��ne9n�}~��נ#9����L;~����-i�T��B�-k����vc�r��]y���9p(,��i}���#��sU��.]�M��q:�K:�S�hh�
Rk��}��ya�o�Z�H�.O�uJ�e�<M�~A0�ᚃ_����*`֍EC�ڶ+�+Z�xP���*9��� �D��h�������M֠�����GG��ֻ�X�tL�d-�:���@D,� 5p��]#�d���ʔ�����1�ЂDk��!�֋i�F��q�|r��.X,����ǰ~�j�*�&��B�J1����>D���
0uj��P��#j�V�3�o���TC��K�F�^�&�E<A��˓./u�smA_n�m`.R�
F
<����8�Hȅ�ܷ �$	�P� #�`�3�A]k�i;�n�I�@���<��`�N/6ź�/]Z���"��6#�n�aWaU��#(CDP9�!�Qy2��<A٪9e@�nB(�P���<=��d�u�
2��8���72
.���l�&^��0Ӈ vTKs@?9��D������?	`� �78��S��0p���,�0f��"W��/8r;��`Qe�޽^s0�&⎵au�9 �V����OC���ÏP u��X����i�ؤ2�K�>�9:
��H���$XN���(Q;Tq���4dkB1ϻsJJ�1nݛ�b`��3Yq4+��ġ�Ɲ��/�hyJ-�E�@s�Op
<o�	@��8�B.&-ć�7U�4�9�'���*���DrJQk��R��hvO�/D%<xtǔu��B�I��̎B�ఆ��� la�˥C�(�@QdLn�hP�I���t���@�䨆����xy�a��F�6����@*R��i%��b8-�3ϓ�{<�rEi�5Vi��Bp�Sb̓Vh��r��� ;�*��W/�	�X�q��;r}$,2��4^�dؐ�ȄeN�;��#Ja��'��d��&:sy(n)o���j���6b�+� �i`6¸K�
��H<��,�p�R5���G�j�y0�ݳ��7�R�C:klB-@�҄��g
�4ݤq�&�^�7�6�ZԌ+mq�sM�h���rCH�/E������2���^�4��S�+(�iA�dO&�~as��դz:���brD�� �V5A�NYZ��'-�eQ��?������RX �A����h�0:8>a����"�v�)z��F%(?�}:���2(�= ���#fy�/��[P�W|�TuԍKW���T�L8��/�J��E1�B˝[�Z�!�`�.1�L����V���;
4嚠h��^�Q��� (@XX$�/��XxA�v�b)�"$}��5�.��@
�X���m��������i��`P�Y�v��@�I��XI��ۇkQ���Oo�ث���y���[�|��`ˌ8�X�Q��<zߪH����yj��'��E�ࣚ�,��@ف�Sn5=��
1��oژ(4�D�E��$y�:�N/W�`�2�/�kXQ2���V���J�F/C��u�6%Q'%{
��O����j����@V�CD�$0�,�yN)�TI��Or�p�$N�jT�g�I�b��T �GB�(8�OxH=��igޑ�WN]�:�p@b�D3�~]y6F)~��逳�O� �X�1W�e`@���9�P �yB��1Cp���Ǐ7k,�d��'i:�y$�Φ��F�C�Rd�T��3%e�ȲQ!Μj� ��'I�v$k"�ɭ���#D�=�T�S-�%��A�L�'h �!��Kl��1T�֎
n|x��%C����f��<t���H5W0�`��[j��g.K�l��E�!��D������i������ �S�k�/Б����n�0	�B�xB�ݲM�FMz�%]�fBl�����8w����T妽#�I.9f��iP�\���8RbF¥k���cƘ�ȹ1��#$g$X�&�I:9g��y@�I]�5�Aɤtn���@E�9�:�!eD
3�|G��/F�����VO�,#Q��qg���p!e>�95�
��yI�:+���HBIZ.6�|8kTM��l����͎'����g��֮�?���4��uT������{ x%�U,1��Q��Aۣ?
H6m@/c��D��f���&D$��`��
��ɤ��6̘����\7v� ��Y'7��q`��Ɍ=��i���
��q&�`��g���Q2C)�0����C�ؗ0�`"��x�Jm�#%ԇ<)�U鱣�%�\@��/���'�ZP��/�;ZR��ɮ���'Y������$f����5�ā�g���+�f�v� �I�(

d2o�=eiT��gY7�p|X�eX�#A�����18G,q'���'0<N8Y� \�!��b��[XNY�⟮s�ܘz� .#p���Շ4!��Zw��+C6&0�bW�Y[J]�O�|l �w*F�Z��Ƀ��)�N�1Z �"#B-0&����
S�6f�Ub��
����3�֎?N�u�BM��dt��
X<5b�ȓD[%*�Ё�aG
������=K�OW�BjO�� ��XF�����<,v(��v�ˌ6���1��!J[�O��C��I���� b/mW^aD`͓kuB2���f�В�U�D�(���g�	�E�<��F%!5 F��jZV�#�EN�eʠt���HT��D�x�'$��rg �fW4��B�%��y2D2���1�x�L,�S��o��-��Q�x#���QR̓�A�~$B@�7��O-����[.A)[�b�*H���Y�'N��24A�3,<��4���,��).@-S����ܺU�BaW���Q��e�%A؁��um��y ��4}V�xB����T�Fe�'�'���t"��
u:u����r5Lx(�O!�iq!��$��O8���@D�r��P�h��pt6�Yg�0e�N��Ȉ�DaZ�Gft� [��Ċ0d�D���'�	n}�,
�b�$ear�P/_��8�	P�'C� �R��OP�(Ik�$���q$�y����Y�zKJ��	 uQ��b�K�z��*���{J1O��:��?N�����J��&i�@X��*�ǩPz��1�@#?�Ow��i@ ?�B��q�592�1 � J-F���@��.@�S�V��RDK�I��`�&�M�XԨ�Pf��Z1�I(BK��m�� ��fV���C�$��x���L�\ܦ�p&��ؑ8wp��̙t��\[6�'+7����ʌa@��ٰ-
� \���+&�&5F�ָdSb LH�rR��s��!�B��nV�)B�a�e������ X╠0�P��"h�����-����3Dx�Eh0MY7f�ZI
�햩	��*%��%c���` �0m��&���"�$f:���@�U�SإQS��>����G�<��LH�21OӲ�\��+��T�����D�i��y�#˚(-�jhM�8M^�����>������&<O� �1�P=_.���J[�k.�x�MK��P�S��E�Fb�%zӤ(��a~�'B`E��o(
6����_
���'�-{ҋ�n���tH��r8zT(�I@�6����g�O�%:��	)MV�����6�b��G�8���*�C&0!`��F��<��{2o�-d���n�JmP�J3�<�����ы=�0�R�(q����s�'�tPHF˒�q9 �"Q��'����t(�2B�!:֧W[���'��pB�3:>^��D�szP]D���!��c�*.C]��}�e��v�&H#q�Z�_(PL`0�і]��*gkC5ê�E|�KŊ	�)�ba�.)r:�c"O�2Kj͸#��<t��Ң�B�%���{$�>[(�k�-�k���D#$|��BQyG|R-��C�ΕHS���Z7LtE�6�1l��쳥j\06�h���Ul����`n��bae*�kL�	<��:2�G"O��ٳ���b���� �l��l��~R@�`=Y��Q�`������0@�L�a�D�2a�q`�NG�*�=9v'�1��'�����b� ����N�O�b��%^�YFLd�PEsxI����,\W�e�E��WU�gץL�j��5%އ[CBDXEс��Ć.{cl10�F�Sk�X����K�j��G�WKz���U�'޵���X�М"�-�DyR��-���M�N�F�~�Y��`۸�b!j٥ S���䜒H!�S Y2H@�`F�]5l��tx#�	�ז�����",j$��'�L!E�6�*�����sXu ��SP@ȅ��vTUH��0VZR�QAN0��A��HE�9��J+�M�0�Z�Lk�1��H9eF�2%�B�a����Y�:�,�v��*�?� &�\�8��$߿���΀�}رO���c�4�he�B@Z~���:�b��%��D��R���~�d9*�h��w��h�S�P�q�X(��V����XN�?"$�,�2�Ab|����WV���K��,{n�	�	�Bdv�a��P��x12��E��DpQ*�k ^y� �';�x��Dx��"Q␞dW0`8惐��%��e%�� B���#;Ī`� ���= �%r�I�N�6]{�Q�� �&n�U0���B؞@�� 3,� PM� 12U�VmM`Yr�!�;u�p��7/!W�d���%F��oD?��j��=ِ��DH5p����c/��k�O,HW�$��g�1ir��	6� �ɜ<p��s�씞;�0A���ߟ����:�@��s��8�v [e��)9q@́U�<U�U��L�0Qn���s�\|��C���=�`Gy��P#�r��i��6�=!e��s|-�a.FN�hA9P�|��2�P!�h���)W;�q�(D�pz��,C;=0�G ͖wy� m�$$�s#³y�h��I�\Q��(�Ɔt���i�!o�7m
=��X"�ܝ1BL@Z�a�>���ODh
D�ퟢ�CE/S18hR�-�3�:���Sl�(��͞4�h��������� �.]���Θ$z�"��I�	n
��k�7���D��&030���6_�P��]3L��q*��r�
�NQ%.�]k�N[-u��EyB
	t��e}�� 8U�`X0�5� �M�∴`�X�턛q��ź$p!�hK��+�D�Y'�/L�iAgbI��(O@�D�hn&��Q��t8�S�'A���F�J���y'�Z��̆9�]Ӳ�P�%|L���"�>5�<�{&$S�5��}Q�O"8�ӫB=cJ>QA��'��ĉ3Á#	@r��U��5jP�+�81(�`�ל]�B#8��șscA"If�����7nT�ϧ8�!���T�s�!M� �1�'yh�!�h�7i���BМ!�g��`��p��n8�z���D͙#zl�'wߌ�)W+�#m�ͻv�B���M
r��DQ�+�(�&���I�:ܱ�k�T���i��ߡV�(�ӊɻ'\$@�/���bU�B�2��� V���Ez¯
>�^ [�H�L���gL����Ortj!,�"D16!���M�we�a�.}�D�� D�<��Ґp�ڰ0�J�6O ��	�Z.V�Q�$�!e`�1p)�,yʔ�=�����=dH���5����Ѧ@�U7�Ӥ3��i@'�;se�P(�.�z<4B�,?"�X���� �AH\4E�ГO"�a�Ÿ��O	^q�T�^x}
(re���te���'�9���S,�މ�E��=i'��k�'vl���.Y�AL�$Ť
W܈��'y����m�2� "r�C:D��0r
�'�|���J��:����(�IH���'"��r���C�ܟ]�ؘ��"O�u3�� A�l�U"̄;���"O)��"M�0��w"�f��!;v"O���c��z�*yGn\�^=P�P"O����g��6���k�ʕ],Jс�"O���bN�"�@��P1N,��"O��+j3(�ҙ�JD,>�v�R"O�L3w�S�-��4c�ZE���� "O�P�懍[pu@�O����d�1"O�4���̋ �ڐ�Щ��.��%"O]ۀ�Կb�T�u�0|X��ct"Oj�y�(ٯR��mz���<IA��X�"O0hKB�_� �'�8(�
�"O*��%��k|�&�<=4|�e"O.Py��J*O`<�ʔ�#���id"OP�@�ŕ���|����G�ȄYQ"O�٢0@�6����hJ�s�M�"O�kpC1X�8��hɇ�"O�Ѐ�;i�ĉK1eZ�i���"Oԅ���a��9�7E[;_�nP�0"O$�j���rJ�uX�
+n��ѫ�'���W���Ba�x�1ǉ/JER��	�'o� �����Q�}�1�ȍC�.d��'����RI�	k3� "#�;Dl��'$X�����
�Eݚxv[�'��t#b�B�o�$򑉜�s �����D
�"w,@�6	 ��ʝ3�Y����l�u�J�XG�8Y�����>d���Y׎u5���e_o�j�KçT�t���9� ��L
�@`��Q����d��+�����4� ��ӯ�^`8y�2�S>X$�1*@+:����3�)�'tȊ4�⤈PoT2��Lf8�H�����'r��i��!A�<�І�;�\5+��I�}-��8���%�F��sjQ�q&��J�b�<Ntj���DɼNuh�b>�
��[,��<�e���k��4���-���\�'1O����i�- ���!MO�mK4J(���
*Ot(��X>�HӍ�� �lI��i�
�����G4��d��O�P�� �%4=a�4�Elӎ��"�ʚYDb]��B��y"�Ȯ/ì��U�yp(��	çS@�B%���z�*U��AyP�0d�TcZEp@�G,R����'�N��iD4"%�@�Ι]��1s�M�KIDD+BJ�$A��u�\�'�����sӊ��Ig�,�w�N��I����?�g���&���1o�Oa���
B��	��� /ߛ�MK��8�6�he��O��s�O�lQ�JB�$��	�f��  ^�# ʁ�U�&�PP�'n4|�ɿ�0|:G�T�d1�%�� �Ze��Zb~Bk�ɟ��6`7���(�P#L�J��	c��Y���ɋE1�ڰ��S�O�2�S2KQ>m�2�(�c3\A ��%���v#�)�'9����̈́N�X9�T�=R��c�ΰ)�qO|�7>eIÁA<"^���φ�K���6,4�O���&7�'�� rY*�k_a5v����C�HDJ�0��|��.HEH��=�}�$ ֹ6|�"&�ǋHG�f��jyb��(. �=����V/R,�A�#N T(%ku�!��l�|�YTL@�BD�	pɌ(?�!��-�Q��/A��<Zs���!�D����2��]9��	¨��x�!�D<��pb�LF�'�FP�'fY��!�E]Wl�3���!�b\릂U��!�Ŗ1t��
�gf80fBO!�!�D����LPw냘lU�I�G"�1[h!���eD��"D� �08���L�!��;a��I��Y{�`@(ŧ��!�$@o�E�􄛥l�X�fG�&�!��\�_�9��F�����b�� �!򤏪zp����c�c��y��D��!�D��"P�C5�b�DL15d�!�d�<�T;�iJ6:�f}���J�1�!�9��8�d"	>#�֘��`u	�'��&��9N2Ńt[&uD���'R��!�ߍ)�����撑W_��	�'D�� l���^,C�d��\�\��'�&E!��Ŕq��h��@�|��'r0M"�Ĉ.s^��զ��j�<�9�'56,�L:H��z�b_6E��'�>��5!L���%����.l��z�'���:R�P�3t�;��[��a	�'@�X�6�]P�5�'��{��s�'˲=��$�xv�q����7F�����'�ڕ�%��]�z�ڶ��<�6���'s�03V��
JN�W �:
p$��'��p�ۙq��\3���/?J�r�'&��J�]�v���)(����'!�-���">���q�
#�K"�yR��3���Rc`�R�C�L��y��C����d���
a�DJ�,��y�'0$"�T����  h@hA��y�g�}���a7h�vKx���@T��y���CXL��/ǷV�(��6/�2�yG�$���`����r�xV�O��y�b�*\k:`�أ'hp���[��y��ً4ܵ
�Ɖ&p�IJ��N��y2�P�s�����N�f���5��yB�6|�ʝ��+\%	�h-Iā^��yB�ާn�<�P��������yR"��&��]��0��X�"X�y����#�hԁN�/�0����y�a�|�x}K$�9xC�Q�ŕ��y⯅L1��J6s�<���I�+�yb"V�m����o��g�r(H��]�y�cű�*D*uBa��s��ܸ�yRc�qk.pI�,PPs�bK�yȚ�O�=��o�3�ͫ��/�y(M�?jT�AK%����յ�ym�� ���7��">j�����'zQ��hވd(2A�Q,L�[�j�[�'��GF��3��YKa�-S��0�'�b���I�x(�
6�՝<F�uk�'j��[4$�,b��&N�32��H�'�N9��&BY��-9�OQ�.��M 
�'�@�u�̈́c�CcĔ����	�'9t������)�E�>Ȭ3�'knm�
I~1�@X��X.p'�y��'����d��g�t�!�@2R�b	�'�mc@�P7#��cPE�.@*R	(��� ��S���p��4� ѯ4�VE3�"O"���Eh��A����p"O�1c�3J�� �@K|��9��"O�wC�{.t��Fu��i��"O����/~��8r�"g�rM��"O�eA��]mP��2��U&�U"O쩘n�V���T�
�\e��"O� �#NΒ}�<an�Y��0D"O��KY��=+䊖;�n�j"I��<ђj�<yS ` &K�x�\]H�<���8Tr�{  �s�&m,��C�I +QҘQ��I�wKP�1��!O�C�ɂH|�2��տ��+�ǋ�PhB�	�W��1`U�[0sJ��
��
�x�JB�	�=�$�TO�T�,�`�ɚ:�@B��'1�d=���!K���pA.��R�fB�I�/�!p�M�C�����*~C䉊m�z�`�bD����B2�v_�B�2[�u$�y�8��p�Lk��B��JhN�B�F�B,�@!f�ɪXنB��,#m�Y��@��d����-G$�fB�	"Z���#��M�͠`yr�	C�I�+E��;2�ٖCF�����@�3"OP����um����fկ8b� 7"OXH#iAl�f�%S0��ٶ"Ol����4� ��3Kî,K"O6ղ��J5��ͪ�ñM�8;"O�%H��ذH�@0#��9hD�@r@"O�����_�[��((vG�MV8 �"O��:g�� =y�E:f�MJHŉ�"O|$y���R
�cU�@a�}��"O0A�tjؑfݾB�$՚"��X0"O@���΋�ix)��d�I��0�U"O���F��;c|��񠔉9ؐ���"O*��NbR�@ؕ��K�^8�"ON�+��Ɯ�Nl�4��<�!�"O�ի2�H���5C7dI�.�D�"O(�k���f�N	� �
�9(�"O��/�-?=�S�׹��%#�"Or���\=����*��i��"O��[��׋Wl�I�g$/k`y�"O8��u�wG�Y���L�
X�"OLEc-��.���@I�1�j��"O�I��P�
�0Q�
���"O����`Ǉ=��l��h�*n�h<Jg"O���ד1.�|p@��fE��ȓ d�ժi�D�gkPDf�̈́�<�%H�/� n�ph���g\��ȓK��J�¸u�\p���Na�e��|S�]%o�v]�	Pǌ8�de��c��8�`�!C:DS���2�ՇȓfVD�2 ��@>��ؗ�>U����O�p� �SFN�h��X�vD������z�CT�Q5���nO4HB��ȓw x�b��R2vQX��B�$��\��B�p͈��z�(*f,�" �8Q��:�XA��+3�  �0��%Yܭ�ȓ+$�DI" �=F���!�a?Ksf��ȓ<9`|y��W�X�
�$;[����3V���D!|n�2���tK:D����L�^Zp��V.tMN%X�4D��{@�Y�/�x� ���[�p�Bk.D�`��ߗvbf�b5`�*/�>t���,D�D��	\�GA6[b	�v��@�*D�� l� "E'	J\p�!�L��"O!�cE# ��q�ʄ;�D�@6"O����
R58(ر���D�"t��"O�+��0x��d#��2F6��f"O.Xb)��(�b-iE�>$da)�"OQ�$������KU��_z��A�"O3�#�7��hIp�70a�}��"O��q`�L�\�l0! BN��-xG"O�m㧢ɂ%��H!�a��h�j�+�"O�Q�t�O&r���b�.�&���"O`m
�B�~M�v�� /���"O��z�l��d:! �+
8
��G"Op��B�; tV�`��X�܁2r"O:��!@>w�60Z��(h$�"O\�C�,�,��	��9q���q"On0����U��ŨaT�i+�"Op���q���'g��h4��k"OYi��6
���E�=w�d(5"OI�w.�1��e�3A�@4�B"O����P>����]X�8"O`���
ơ	*Jɻ6o��F�
���"O��� n]�_~�p�m��q�"O�}R�eX�Ei�8����
r��0�"On�+��0$i��h#��xk"O0�ڒ+�
@+B �@D�`��W"O�m��:y)�J�(0]�d�Q�"OH��U�7� �Ȇ�"&I"w"O�V�9=�h�Sń8H@�p"O�ͣ�J��%.yӃ:F[�r�"O�����Ϳ|���u-�)|) ��"Oةp�]�L�MYd�шC�]�1"O���	) ��s��� 	T$Cd"O ���[����rK�k8H�"O ࣥ�$�u�GI]�-��"O�5��Ѽ\�.�V�N�y�!"Oqx����)�beG=A���T"Oޭ�]! ���K���4�\ж"O�\�珤]���2r�� ��qcS"O���g�=���G�8��ܫ�"O\�4=|�A�@wd4��"OZ�Ȳ���C=�Y+��,S>AI�"OH�ƃ�(���B�)j�*�g"O���"�I������W�n��"O�9Pq��% N��R%�W�h�,�"OX���ѥe�" �"���j�n*�"O^��6o�*+;���ՇL�o��)��"O>`�%ւ[m��j�MI�Vm�X�"O�4��u2N�d��c\���R"O>Ec5�SdL!kǫP�ZTZi"�"Ob`S����e�=�ՌݟXO��m$D���RN	%�����ٞu=ʬ���(D�D1�6��h�D�תc*���:D��R�݊f�D颁eֲ1�4ű�F7D� ck��x(ܼRSTF0i��2D��#��_�j�+�K�N��H��A0D�j@�i;��'��:/����!D�I��n q�t��|9P�Rd D���`��n��E����&�p����+D���
r��P�M�6���o� M�!��I�l8��s�n�~�wL�j�!�No®�i�� }�ԕ��جi@!�T�c$R�+<ňz���d-!�d2I�V�ʲh��q�4YC��ۅ;!�&2J��𨈀��y)�I��!�� P�v��,+�`��D�9�T�"Ob��3m�7D�<��#��/�|�
�"OV(�Vݟ8�j-+���$	��I"O��i􍐘.�H]����J^le!�"OTi�hH,S���!�ap"��"O�y!"FUf��R�BM�nRոw"O�	�	`I(-Za���qh�!�"Oȝ�
'W��Ɂ֊� X~�:P"O"�U   ��   �  �  �"  t-  �7  �B  �N  �Y  Fa  �k  qu  �|  �  ֒  �  Z�  ��  �  /�  ��  Ǿ  �  L�  ��  ��  �  \�  ��  ��  $�  g�  � �	 ^  ] �# =* �0 �7 �C K �Q �] Ye >m �s �y � %�  `� u�	����Zv�B�'lj\�0"Oz+�D�/g�2T0���OĴ��� �?YV̒'�?��]O+z]I'������Q�tO�eÃ��m@�I� �1���W�Y�N�.�I�T��I��4iBh��%�fybÑ�(�Z�v	�	0���E	�6�q���90���;:a�����Dh���I$����h��FLݓ��9�8Y
�F�>]��d�fp,�bT$L���oZ�h�r	�Iߟ��	����I�S���ac�J&&��(i���O^�5���I�P}��#S��M+���?��CLh���'�?��3R��E�_8]["���fO�C��8���?q��i<2�'��'UH��\w|VzT��%(���֣ۀ40�LbTřn+��q'j:��c�Pj?Q�Xsv���h���]�J<vL��!E�cJ��'��d �伟��e�� �<�b1��|+�[�it����@.Z�����'�2�'���'t��'+r\>�ϻi�~�F�*ڂl��É�`M��I��n�����4כ��'j�ם�z���ߴ
N��5�X�b�L�S�.Q�C�>`��A
�3Y��@t]�p�޴n�Z}͓D�N�[��N�<d��'3Y���'&f!&���~�����ұ��@b ��a��o
�^�4=�	��M"�i��D۟\��j��хL�.����mæCE����ƒߦi�EE�Ce�M�ԡH�0����]�Y8�(�*�MK�if�6�[�3�<9��k�$]h����25fJ�S�� �(Mze���H޴f�����Z�$)���򖬌�Z���3��$XH��
��00��U�X�zNlDD̬<����i%�6�ӦI��W�n������V�:�օq�c
1��i�2�ާd=|%��BB2dLT۴ Y����׬VrX}v#܊b.T3����'R�Dr�E�.i��(�I�ND�h��'��O2���O��$n����O�f�H��Q9i�$ߡ�T$����Op�d`>�����E�����'# �Lo�:���2��A��3D�H����I�p�h�6*�)8DR�:��M֟$�׮[b�@�v/۹]�~���:O[��'�<�BM	G��LEc��P�Ę�*�ٟ��I͟��?���?����y2���#��| En�X�u2V`T���?���i�Z1P�Ŭ>,R�[ �U�>�RI�7�w�h�)�B�X��i^X��O_Ȋ�Gr����J�O� �T��.SH2�'��$��i�-���K��\lZo�'	ަ|�F�4Nφ ��^^Э��O:�jc�7R�T r��	H$�}r�/S��x�֢�8�T�G@�O~r�E��?Q��iF�"}:�OI�X+4Oݩ-�4 ҖlW�<UU�L>���?��ǈ����ق�N!�N�sj��A�ɯ�M둸i�1��5� �\��6	r�,տ`9`�XD�z����<��
6�b���?Q����$�y�@��T�~���1��4�hԑ&��+��l���,mZ����TU�B�X�b/B�"��QƏTL���imɩ�b�i	J�~�h��n�ḨD����'1B�{�O;?�̼��Jd � �i_��W����	�?Y���g���Iu".(�H��Y)������?�*O$�d=�H~��V�-?̨6cC�4e��;�J-��dʦ%Z�4�?ѕ�iT��?y�O�BT`׀S�F��|ё��1��u�b�y:��?�����|�Oa$�S��7XnDs���{~�x���W�ry+��B�uʄy��'���J EU�7 �
��Q�����H�(\5�� `	�4o\�в�N�TE[��dF�-�墳�G�|	p��0*���;��'�p6MG�'��O�1�u4ҜsOLȕ(����'��'����bC�Kq� ������N>٦�i��7-�<�,�@����'�"�Y0 ب�!A1 ��]�S�j���'���jb�'x��'^��l�1�(ݘq��z�Z�
�`03�]��%�?'����ˋFLax	�9>&0�9��O<��ыA� �(#L>lajćV�q�l�4(^�;�Ey�����?��ic�7�O"4H�A8r�p��M�δ8Al�<q������)/?9����4�ʦ)�w��)�M�w�����4'�"�Q��F��*Y���Ҳk\Q�i��	?�����
%�e�<��'sk�f�OAV`��%�=N����t�Vti��';�b��G;�x�L� ;Vл"�Q�2D��}�a��ic�$i�&Y�#ܺA�������*Q.pъu�7'��6���4���cV,[��aI#�>���Sk��8I c_�'���釖��a���O�o���ħ��O��[���Z��Y<
М�R��S/���?�N>q���?�/Onlj��G+T�Dx�M����`CD�d�'5d��r�,�$Ȧ����.	 å�K\�X(8qN�N����4�?���?!�O�5�� `���?Q��?Q�w�$Y��($� Yf%��uJzQ���@!H��i� ��!5����OI��X gg�\�&8k�6@������Bv��k6i� 68)dK^C��c>)�g+0?y⋲Jj����5f0<���7�M�U�<��i�Oq�R�'��l
z-[ +�6ư����C#D>�'�ў�>�2�U�~�|����H����<�u�iI�7�+�������<I K�- e0!Kӈ�F�D�
oΟq=H�cB�ih��'!"_���O@��M3E+Z�2d%�� �, ����J`����U=u7�
#�N
�0��&DRB������B�^�0��Z�{l�p�`7G��u*%/	
b!R�JW{�X��H�2w�e���ƍ | [(y^���������<$��"��_�9|(�"�L;H)���Ij������o�'��R�(e��kBȎ>�e���'S�6��OAm�"�M�.�� n�SԦ�	�<9Wi2��]$�݇@��z�I�ҟd�'b�'+󉋰@��4�޺b���3�pӒ� (q�6�Q��8�k�/!~�����'��T�ǫ�o�U���Y�8��}��?�-@�I�t9�d�磒�t����DºD@g�N��'x�X���j� (*mG$o�XP�J>��d.�	H�!�#Ϙx���Fx�����̦)7Y Ka�`��!E�����oJ�M�(O�Kc��Ϧ��I��Ol�4��'�� ի�
D�M�P��%f�@1P�'�B��5
0�cg)J��H��056M��C>Q�S"jz�JÅ�
�V@ʷc�7d��v��Wi�\�z��gGI�`P�Q�ߗ|���O�t!�1I�/0$�������n$4�OF���'�R�ʟ��7���^v���2�Hj]`7ǋR�<y�C�N�r�1S�()V���Q	�N�'�Ģ}���#As
x�5��6�Q���Ms���?���q��c�冨�?q��?���y�Kӹ5�Z�Ƒm�*�Cu�#�t�Zœ7Q�i�5�N�c{(C����|���x���C-��.��Eb��P.,��$iW���	��иau����d�|"�IHx���&�R��	��ƈ�?��O�!�'GR�'��O !J�F#Y���D��nЫE&D�3��*<!�A��7p�H�Ke*�<�G�i>5�I_yr ���Њ��Q� ԚX8Ut�ᐊ�����'A��'����I�|R#�B��``"� �K"�B󀞘ǲ��+���r"ֽeQ�
u՞�<ѥk��0>hժ#炷K��Be&�D�L�9�C��	R���ǎE�f�icw�P(�<I0��>(1
��ViV(e�ek���V���I��M�!�IH�'Z~� $�h��91����e&n4`
�'�r ����T���FMD\t65I>	��i�W���Ӭ��M���?�ub�!r=`�
� BhJ�N��?���^�L�S���?	�O@č�&I22$FH3M�'@�᛬f.�(��a�"h����J��0<Ic���!B	�d9ht���(�:��D�=F�l��Fٸk�����&(��$t�ɴXl���
�?I���ٓH�C䉻F:"lV�٧h�����k�K/F���KğhAt��7vy���b/��W�Z����2��� �F���O��D�|�!��?���E�tq�d�YT��A�a>�?A���ض��|V����t�cТ�c=h%Hʟ����,=����]�3D@A���pӖ.�GV���ܩ餥�e�T8h��9�!�H0^����j �̓4�?x��;"�O'6m�ɜ+~���O��}r�'� �[��E�w�8���ۄb7:���'��1��jѹwQ�|��K��]��X@����T�O�L�c��4���j&��RC�|#��?Y���ybI+/�x���?i���?Q�w�`�C�*��r⁡��e�持��Jl[$'^J�:Ĳ�IN�ϘO��@%��P?	&,Š ��EB���@��S��3'M�b��P�u	F	�Z4�(�DM7s4!i�wi|h�  �qq�x�N7VզAY����͜n���'ўx��W:��JB�ØZ��y��C�<������c$z��8�������&o����ן��'�6|�
~� ��&
,!JT�u�;"�Ё�0�'ZR�''Bk����՟��'�`4�tL�=;*��eH�.G��^I�\8���k)j��a��.��ؗ(ʓU�h����TY"��&"N�&!@ꆡ����U�Dj]�QEޯsa�<�!ϊ�
���{�Y���98�I�`����R�Ï&zr�x���?Y��$79��1��Z�t�t3��ڋ-��ȓf�����p�H� [DT&�T�ڴ�?�.O�D�h�E���'�v��9��*7�%d
�H1�'nR%�=t�r�'S�	�""<LeB��-MbF��b���ڹ@�ݡ}6<��g��6C�`��C$;
����ڡp_���`�>j�ʴ�]RPU�s�	�a��L3��؏1�d�h��؎8�N|h�*�/ո' 8�z���?��Oތ�M5=唈�U��)'Ԫu�V�|r�'��,"�]�Q۞���M1rߘAx�xbF˺BЂ�zD�ͥ	�^�q�/��?�.O���0D���,�Oڒr��'�@� ���D+� �55'H��')��c��R�D�iՔa��$�
6�~�*�.&�S	0��p�΃�\d93�����E�쀱�`�'�mxR�U o<ݩuM@�U�F�?!c���NP,�R���~
��E.?�jKȟ��)�'�y���:M�&��2��,l�6Qk�!��yrB˿D��������Vf���O�0E�to�8�Z�I�������돊}���'���'��u�Ȅ|b�'K��'���O$>�q�I-_#P�El��(j0�"�� ,�FPS��Bkٺ�P�	�k�h���'U�!�bψ2i�*	!���f��4�&�f�ŉ��$Z�����w4(�����Cj^:e��.=O%�z�n�yzTxq&���mLҕ������Oh��&ړ�tyJ�%E}4d�k#�ԨA�' 큐������7Oհ	�.H,O��Dz�O�"T�\�PH@�R� �ЃݫdEx���F6(D6���Ο��	�� ���u�'��9�.���%͑s^ 	 �*M6����i[(Q� IÜ��(��D�g�|=�,͊�(O\YU� ���+�,����*�%ܺؐī�_���
��3y�`�
�y��A���v�y�]0��#���� �4l��t�� ��H�
�'��%8��Z�C�y�@�9$�9��I"�[�D�w6f�Fg�'���%�`��4��-�qƳi�r�'�-;a�T �B�BK�2t��H
��'�R D�&���'jrɞ�0i���m�)t���CV()�,�q2��c,|�ZC��C㲙e���@��DR�`@<Ik@��<z�VY�������Yj�](
�g�^�d� yZv��?aw�9Ӌ�d3=h���@t�'8�3ǃ� $>ٸ������ �O��D�OV㟢|B���*�  ��d}��k�������WM �S�O,6�ޜ�"a����%��)p�����m�vy�#)N��6��O\��|���*�?���@�W T�� �[8SP��E韩�?y�0h��0��i򾹃�c�PgTl�s`:�q�͟<�˗�U�H���#�.8Ԍ�`����#K�j��J��P;L�VW�7gA6�P���j�����:`�	fH�����H�l��'��Z��{����,�'��d��I����	!ƍ��o��䓈?����?a��i�y�8)dM	6F��4j3O�t�џ�9�4+l�F�i��#6uX%Ŕ/�Ra�'�C<(�7M�O��$�O�	��F�kJ��O���O�杠j� �
�1R���q��;]bt��D[����f�ѱ(ut�&�*��j�* �WX�i�ɑ7��,��y��ߝL� i��Q�H�Fx�3�,�SH�I#!���%�0ܤ(�(]� �:��(?qa&��T�I� �?atퟟ>E�������x�������y⧔3\UV��f�D�����m����D^�����'��I "�`�{���<Plpa�h*O���ƈ8?�T��ܟP�����qXw��'��i�x��P�i��V��,�t���
3:\�jc`D�z�V�"�:����T�Ф�V� j�2=S��Ϊ:!�-p�菇:�&y��+��O䈨�@�)�a@�$C�J��
Ci����'��d0�'0�`H �M�Q	 ��#բxHV͆ȓ[N!8��R��0ԉP"-�f�&����4�?�-O>̐�ަ	�I��l�«55�%�"KW>&�$z����I��n����0Χ��EZa�'Ѵ�s҄�8�?q���W�l]����8:V�
��
_���mΔG�F\���u<2<���I;�f����#\����hW��xR�8�P5������}��Pa,Y�!P�3m��o��ȅ�}����� �H�`e���R��"ȅ�I��?1��$J>�*%&A�<��Y�@�s�	8E�HIQ�4�?!����I��>����3q����T��X�p��Kj�0���O�P!6��`�p�є�M+q��]��|�ʟt���Q�X�Z��� ��h?ZX ����[b��73��4����2�~�G��摊a6Э��/��@�*�̛���x�F}���d�Oʓ���$Zj�rQ�r�ס3L�����ˢ�����OB��O,���1ۼ��M�/C����aʜ{�џ������#Z؜Qr	"Srht�GOB �oڟ��	şx0T'O�&7������P��ßt�_wm��W ��LUJ��oo<u���|��ˈ^
az�D��83P���G���hp�7N����× 8�Pߴ=l(�7/MT�g��: {�$��=I��Ӓ�T�o�.q�	��M���[p���ʘ���OЩ��"�*,�%"�g�I�F�1�=��0<i��4��Ȉi�7�F��a�GryҌl��m�H��?��Siy��T�6�`չPӫdCE0dG��`8P`�X�b�'s��'�b���0���|�ƌ',�����Φ&��ţ�+վ�\m�2��&�z�/&�>̈́��v��Mb�+C?Y|���D_� �j]��$��l���ʱ?'>��n�!J�">�ă�N�^2&㑐7��XJ�ȇ�N���,��?A�i�4����ǂF�`����#�q�<��Jƃ&؂�JEE'}�l��p�Lp򉘂M;I>������'����0$j0���ڷ	�!,Q ��k��?i�ŕ�?!��?)1�Ą@=9�t��<jZ	B��X�&�܅�C�7Xܸ�ѢA2}��\�R
P�gX��Dy��E�,��'*G���A��g`���<g,r����r�NU���� p�VxFy+���?Y��'��mnVq��R�2����"C�B�D�O���&�)ʧ8.\<��ҝȓ36:R]�'^�{��q���Q
��&�ڸr-\�����=�'[����u�*�D�Orʧ%�����C�(|�#Ls�`Yc��F'FK��2��?����U<����ñh����c�i��Sc���	�uix��c	�7۪���'X�O��ɉ^���i��v�v���l��H����łN3��J���o����ە��O~1lZ��M�����鲁Կ>�Y@�̛)k��S�|B�'Wўh�'���G`�>�x#�*@D���$�>���i]6<�$�.cv�b�KćK�fU BKZ��&��2&�O����Or�-���p�'�2�')�aw�풷WG�*�;RO�'7`N��2c�J���ǯV.���cF2Ju�|J�`�,]��I�Ge|�΁ 7?�2Պ�qP��y5�Ό.���!�D�S�ht�4�S�d���i�O� �����T�#	�I`.P�P.x���F(��P�P*���C"��ؔ�ʱ7��0��"wn!���U���%)��F��m����v��I�HO��3��^,v��X$�ֺ:��!Qt��03���R�ו}/n��O����O��;�?�����$�-0�D���3m�t����@.J �G̗:Y�%z��Z'Gz��P!gI�j�DyREL�yB�@쁰/$�AkZ�x�ԅ��6�^"2�8�KסB� ���+�?K���M�!�n= '��\�gPߟ�8
�g*�i�A>xJ2У�Ě�)bl����\D2�&����2G�R�	U��%����4��T�LlѓQ?��	+�|����͒�ꗲ<ɼ!��"�O|�䔟]�����O��39�E��M@�,�V��%�A}ʞU�
�8"n=�s�W�c�D�H�"H^�'��X�J�h��;r�ȑ:|��鎊>,;-ԛ*F��	!��@M��(O�٫�?9����DD�X�����E{P2,��X�
��'Sa|�Ą�gf옡�M
�1{*���_���?��'YT�PK��H����X�������,�@��'z�&r�h��	�|��3G��	��i�I	�6�����ԟ8�"�ɟ��<����t�P�ʅ�6Ԗd�Q��/���(p�Dx��I��h����	WJv	�a�K�1#�ɯ ,����W�)�'*���%�O=��}���NM�D��ȓ3�(��7%H��Q��o��G8�dFB ڧ�F�Նߩ0���jBb١c��bش�?1���?��(/Sg������?����?�w�Q�q �!���5�S�/�`H ��&kکQ �3e�.�Q����O����N?	U\�+yn(x2D
#"�X��S�܌c5L��Q�"|��3�?�Rq�|�@ۖێ���l��v'm+��	!_��4?�fb�۟p�	M�'6��!֕)N�={ԁӛ
��ɩS"O��S�
�Qꁠ�&��`}b�Z Y��R��4���d�<Q�ěn�cg���R4Xs�H�tR�������?��?���l��O\��o>�,[c��Bqi�+�m8�k�J!X� �#�v1�a搜��y�E�=?��y��Ϳ\Z	��j�.b��(6��Pɞ��v'غM����� ۈO��2ꘋ vJ����Ήv�4P�c� B�'���9�'�l��eE��V쐑d�I����ȓP� Dj�(�"0��i�����^D&��j�4�?1.O>�'hC���'�@����	�1�>0P�	�:Hq�m��'�ퟘc���'��Ø�&98�ϙ2bPՓ�Ƀ� ��U(�	<�D+�IK9[�][��/�Q�L�ѫ�=�ĥ��kQ�	W��[��')�ZQA5	�!
(n�#�.����O��kU�'Nғ��� JO�R�����L��//$i�5���O*���ə'���!�>�����G�~�1OĢ=�O8b�D �0Z��`刏�D]>A��Y�rP�p��#�M���?�-�l�����O�,Z'�U<&������`^�����O��D
,M��q�c�]���#Tntӈ�@����6�����[,g6�X��ȚVN��'��0���T�2��$�MCMt��S#%�T�N�	�p�3 ��~����� ����W��d{ӈ�&>����?U�'o�T����5�[g��L�$����O������'7�LH5m�dpD�/&��?9V���|�	�)6U�	��%���)�M;���?��\�*��_�?����?I��y�f�o������J�`���}v��5m�w��o����M���t�|b,�#(8�@C ��-F������)C�"i��d<,}�k�P<x��J��ԟ|r��	��cF�9��)H'�å�?��O�S��'���'��Oz$B�ͅT�Ф<Jʔ]:��:D���E$I
��i��W�Hla�<���i>	�IByr��O�=sq)��m:��#A6S�dHR��C��r�'&"�'��ם�(���|
��xvd���'�N �m�C,��rw"��A \jQ�d߲�-H���Y0�PX��-����E�?GxNh�ug�%WLay����L�f8җa)�{�XY�cݜT�-A-ŷgF�	"�Ο����`�?��)�#��) �g�Ք@�d�ǂ"O"r�
�X��U��[θ	 p�|�+eӞ���<�v�N8_(�ڟ@B��Q�y$�x�!�>������ڟ$�Ɉr8����(�'PG0⁇��h0b�搖C��ငcÖ^��Q*���i��p�å���O�U;�/�(wcj�Z0끌V:&)y��^�C~B��� RS��R����qh6�?1q�VßT��@~2ϒrM��e'eP�|å�ǃ���?�ӓ~�b\cѫ�5��{׏\�}��q���(�?)d�$�BR��ZU����ПD�'�����kӄ�d�Oh˧h�L{�� '�Iz�$�9O26`�4�e�>`{���?q��y_�q(u�# P8��qb��w^��r��J%c�����-K�T+	ip�ˌ�����3Ǝ�#&ʟ3~�Q�ei�If�?�ـ`̽O�� h���$4ȝ���"?9�O韰�Iw�O B� .���mE#/^+ӉI�G��qk�"O`ICR� �T��(��V-4��e�1��:�h��dX�H�V��M��Eƍ�FX���j�t�$�O����B��M�cb�O���O���y�a�� ����y���-;�ڽ!R`\R�m��p� (ћ c>�'�P�#C.T�ԂuG\�"ތU���^�Mf���l�)P!KT5=c>�%�8�2$̟t�uh�Y<���e�g�=���d3�3�ɿHa���E�h&���N�+ ��C�	-g�,t����@��E�����z��˓9����}�I+[�,Az� TI><\�UƆ�u�l}#��>dZ��������Pr[w��'���гX�"���D͠��� M�,E�-�{mD�s���p=�&�V������?�2�;#4�HcT���K>ʁ��?\O*�]3�<�p�LK7G�H�ڐ�#§s�xdm�u�Y���qe�4�Vh���d��	[�'��O��&F�;o�t�$L�:F8d�֙|�vӎ��<ebH1��֔?yqrk7�*�4ϒ��hP�'K'O&X�I�B4�}�$F(<�$zq(P y=��S<OT���c	�~�1FԈ�"D5O�������<�DF�xv4��fC��l�i��f�<�"e��|0�U1k�<�����Y��l��I�L�BQ��o� HQ /��.t%� �@���b�&;?�*���	V� *��S�!X��T/�(-A����O`ph���z�|ӓ��6C�H�)�'#:ps�j%>,��u��0Y8��'��s4-IV^�PYr�Y	�>a��D+Z����?"v�3�g$?!g�Y���ID�O ��j�N@�@�ą\}\80���_!�dE������Ū:i �jOG�џH��	�<�h�'�??D��$Ù4O��b�15i�	�\O0��I�?��	ɟ��'�X��7�1V[H��A�4��GH	\���*���O����^�h�1�1O��6nS���H��D�㘘K1���%#���®�i^R	����yR�ѽM}B���a��5�:�(����?I�O�y�Q�'����&Lu��F��;-��a7�G�&���ȓ6����C�G4VU�A��9[ڎ�'.�"=�O��/Y6�b�7d,���E\�l<=��q��_9B0t�Ď\:�� #�[�<����?�ͻ��5(5�:S�N�ku	η]�Z8�I8uC���������%�6!*�BE%`��Ib�/C4n��ܡC�]�w7��A��e��@-��nf�2��'�k7� 8�V�0��6]�%Kg��:ަŃ�iSlL؅Q�Ϩ!��q��j���O��E�'+2�)�*|��.�9�e���0��{���g�	�.�{d�Bu�P=�O���'�̔�Q,M��@�A��S�[�0�/O<�[��O|���O��'N��A���?�Re��*�x�)oĨvӮ}��܇�?)m���T�ޕY`�Y$c��"�<���I3��O�X���-B!I~�b�):_��0�'����b"�!�R��v�AX�X�0�N�3(�Ec��a�	�Q���	�}�) SkU�k�󄈀9/��'��)��6?���*�Q���� ���GC�<ƭW�B���eJ �?<X8C�%D�'�z"�vB�E������T0f��E��4�?I���?y�� '�yK��?����?����?��ꖢ}�����ſf�����Mɶ���Φi[Z��V�Y)
(���ϟ|YD�����A:8\�G	F���p�i@����y7E,LV�1�l���H9�-#B0��'@|������8IBN�l� �B�e#����'?)  ͟���C�'��J75�ΐ��i�	!���( ��r�!�D
�`&f �oE7C�����;De��9��|�����@�N�V�	� ��US�hAa���x(ҝh0���O��d�O�଻�?1�����D]�
W��8��Q�o�2�
���D(�oZ8cNZMе��6�Y��BO�%�x=Fy�lھW!�ͨ6�V Q��� ڿB�A�v�D U��M;V�A�9|b-��b�Sn��SU�2�I�$���W�&9`��֮IWV,h֭�����<���Ovq�B��������!�!�(a�"O@��e۩EK8#1`]�3c�P�EQ�Ђ�4�?�)Ov��*l���'C�i�r�@Y�v�!~�
)�t�-�2�	mV��'W�oęH* !ч��)W���B'�T��8�)wT�(鈵ȕB�E��*�4�0��$
Y��Q�D�k�H�y��,!j�d1&i]<}K$)pU�]<�x���S�~�y���[�B�(��I˟��|���:_����ao@��Ȉ� ��Ty��'Le�Soۉ#i�`6�+:�y
�e��	�6�RȠ&�'�z�
r��*^I��r�d��i�b�'~�S�1q��ʟ$�ת�%O��i#-(%��JQCTȟ"�P�8co��!@���,Ż-!� ��Ih�'-
��೯_2�X�����;,�l���X���|�<)���kPD�P�_�݄��ǘ�$��;l�hŨA
G
-�eЏN �y��V�?��������� �eH�/%t�qC����`�"OƘW��ab\�*�I�Y�N4j��,�ȟ��`�����+�jͤ���l�OT���O�hqc�;�F���O\�$�O���;�?1����z��H�`*���0�`@f�6"�B��4��:���@���1 
ɟ��>a�nױ��afC�l\{��S���
Rf��g~Ig��4�L$�Ohb�*�(v���G���5�3?!!�Ο`��}�'��D�>\��a��	�CzK%���<�!�$�
���I�v�
 Jz�r�7��|������8+5q�cH<*�tt*�n�~�h��LTæM��Ο��IIy��T�MZ�� ����512"�����t�D={t
��|�R݃qe�jjbL�d�Y�G�E���$��q�e��\�~N�Zê�<�����&A�b�Y����ɖI��섷)�8ʊ��L�,G2�9FJ�	�B��32ʞ$y��ނFy�L�'�:�{W&L(������	�΅!
�'B,�X�DR�d����1�L3�|��.Ol�mΟܔ'�q��bn��~ӂ�Dy>Mx�`Y�G H!�ÌE� ��O��Ga�O.�D�O^PSf�O4b��S.SW������\�2@J�L
�!|>">�lc�O]B$A+D-+��JCJ�:0��Yˏ�DK�D'��?�S�{*���q61�
8�G
�#.�B�I+|��l��EG#]~�]CeıVB���Ny�E�(<�`A��	�hk�m���d�O*��(��?1�'�X�z4�\)����$k  �Z�(���U�OʰuJ#-� ��d����s��yI�"�i��'2E&>!K#�M�8%P��&3�~�e�M[��J�М'��`W?i���:p>���
S�s��K6���,N
��dȘ�M��U������y��&�����kٟ��]/pZ2fz�^	Sb'ϊdyQ�'6bꕱt�di��O��$�'���F�]��52҈��t��Q��l�%��Ӆ�'�ҏ^�F�r2O�-*"ן�^w8>��b�0,Q����C3E@���*�x��g���	џ�2����ɱ|��'�?I��I)yo�-�$˔6ER�i�a�={��f��?��l	��xhr�U���ܴ{҈D����<2��Q*�EB�l)�t�a�?ƛf�O�`02�'Ab��!Uf��k�1�OC�$�28�1�FR� )N̘�ߞa�y3O>i	b�'���q�����<!�^4���4��E@�#��\�bO+W���	�?��'+�����?��Bj��_>�#�H�w4���b�;)l]�PdR�M��N���y��D�JD��#l��i�Oڱ��%����;bU�Сs� �,`�#�)�6��Em��8{���ly�*쟴6� �?��\*�>y"s-���ꤺ�-Q'L!���?:x��K4԰��L�]>���'a��'>b�'2�'��'�Zc��Ɗȡnc�M���EQTP8B޴�?����?�����OF�D�O*�DH4%�q�R2�ڱ�� T�%���n���&�\�����&�x��J`]d�<=��8QBB^}��nZퟴ�I����?��I�|�H��da_*X��L9�MH�5�f�B�M�>����$9��~R-�cQ�XAB­d&^��Y����?�*Otʓ��Ӻ#FEY�4����ë����DMu�'+Q?�Z4��=nI�cR=';�
3@:D�P�r��N �r��
�����;�y�%ɂQ>Mq��/pt&�	e�I��y��U�e�L��(i�"8qT�ÿ�y�@��oKF�AˎaJ.!S�C%�y��<(�B�c�ĕY��)5��8��O��D�O����O@��4�h�iCF�!(#\-0֨ƣOehxl�Ο�������I̟��������� ��	9�X8�D��AP���
 �OiV��۴�?���?����?���?Y��?i���|U 5��#j= �lYT�|x�i���'���'���'fR�'�"�'⦴�k��>�S�a�j���5+v�����O:���O����Ov�$�O,�D�ODM�뛜.b ����� $�|�)�\�1�I�X��ٟ��	��Iʟ��I��ñqDN%��;����3
Ș�M���?���?����?���?9���?A5�2s̊�r`��"dn0@�����7����'��'3B�'�B�'���'qr�c�|{�	Y�5�mZ�S�V7M�O8�D�O>���O��d�O����O��Mh\�U��I�~yl��u��$4�Zem���<�I������	����I���	�J�)�wK��$Ā�/�B�v��ٴ�?Y��?i���?���?Y��?Q�����#+��Du6͘�$Ï[u\�{��iy��'�"�'�B�'���'��'cdi���m�����%Z�MIn��}ӊ�D�O����O���O����On���O~؛�d��%���5gN�o�p�`!D��Q�'lBR��D�$�BI�X��,X�:"��+��� t˛f ��'��V�l��<�aSl>0(beV�N�z��S�Ⱥ�?�ٴ�y�Y���̔�Ag����G�x�I;��Ҧqv���B̭D�2F� `�"u�%/%ў��<Qૈ#���$�M=Ot�(�ޟ<�'��'6MZ$0n1O� �iz��Ͼ`Mp:C��k椤�$�Fy��'9�0O4�D��0�c���g[c�a�>-�L�'՞-r� �i�x8�O��7Sf��iqJj� ���K�4��kC�K�li(�ɼ<�.O��<�g?Yr�!8"X�`�V#,2<�&��p�ٴH��'�6�3�i>uMǁ��8��L�j�j��ԪX�<���M#��(���'�}~�ZYo6��T����c�-_�8��0�Ȁ�?�e�e�'�BP�\�|��`I��X�Hp��3;� �y!��Ly�h���!$�$&�Ӝ��-�jt�ԫwK~�*O��$r���IU�O�l\!��%Z�1cNR1������(�֡1�O�����>���bh+���<��癘N*��E�F2����r�Ϛ�?���?���?q���L������c)J,RR���bv��[��ΟH��4��'\(��?ش�yrH�fH�0�ʅ�W�g@Y���b�R���O��Ə�$Np�Q6ù<��'j���q�h�XSc�
0J�$�B��OP&�Xe��5ll���<P�cw)��,�&,� �"J�a~�"��O��X�GY�=w y 3��,���XAI۬wd��{���$'`C(\���چD^�!Op�ಣ�8��e�Lк[<��A��j�l`p��C�|`���Z�v�K�
sT��I �%�(u�T��
q��ɨ�&V����N�K�"�X��:��� E��#Q�9��I�4Z&.�f���s�����8C��f�'ٚ��3)�&2��뀄 \�4*�
�5��f��h��Ź��>u��d���S@$���W�-ƠQs�OWj`ɘ�B�Y#k�4b�$t�B�R&�	��ؕs=f��ū§x^�}�F΋(WF��� ��"Ǭnr�����Ʉ6k.0��[&Z�JfٽB��ceO(]WP�s"#��_RQ�"��<^�ZTa4/�f���?� �@j�x�'a�|�*��0���"����C�>\R�'�2�A��'u�7��O@�$�Od��O��dK�8AE��,lP�Q0����h�b��<Y���?������?��w$;�EE&T\=�VA�R����jO-l����'�B�'���'��	?7���%�(��ÓI�x9P��sR�P�Ie�	ϟT�	�+M\���Yn��3�K+�4�a@��<=>��'Nb�'���'?R��Jf��'���!Om�m*�j�H�Nܣ�M�1@��'��'A��'ݔ�٦���	4��$�LMOЀ��[w�����OX�$�O���+y���'��d���¥e	/o��"Fȏ��bl+�.���O`�d��	h	��ԟޠ`Q�٥��ʕ!��S��&�'b�'rf��A�'TQ������T�;N�\�ҁ��Ipr�afb��H���ٟL��8U�|��f+�)�;X,��&��(b-�܉�lW�W�\�$Ҡ#�r�$�O|���O��i�O�D�|b�F�k\�XId���QE���?A�Ǉ�X�<E���'�r�7��N3�I���<IJt�y�NgӞ�D�O����#`��$�������Qi��R�@�}����+R�J��'N��'�$���yB�'��'�T8hc��#T�B�C������'�2�(�>O�I�O��Ķ<�f�	�N��`�N21�`2D�ؠ�?A��1(��<���?����򤘽-���1��1q�(��͸J��'�j�۟���T�'o"�'��SE��+�|���
_J-�����٘'B�'�_�Ă�B8��nS�	뀨�!D'7�0�Z�|y��'�|�V���B��|�M���1���W�!�J��º<���?a�����@.:U��$>���e؁|�b�z���(L�^�ZD���	쟈�'�r4�t���ɚ�2�>���¾==�@��gS2�'��W��Ya'T��ħ�?�w�)��@�/w�֑Y���K6 S����D�O,��@9|1�(�}�i�3�ٸ0֢��£��}J�F�O�˓X:Zy�ùi�����t�ӥ��D��O���R�Ш&t�H��Ʀ.R[� s��4?�Ow�O��]�Ф͞79��i7 �s�����'�mcIyӶ�D�O4����$'���5g�;��O�'�L��Ȃ�[�ε�Ɍ ��0�'[��'���yB�'��IP�����QB	'�P�}���$�OZ��H�YW��)�O.���OJ��O�,��N�xD�i�M�'z�|��H�O��d�O�YЁ³{����f�	�O����5j62���D	(M�.�P�ŀ4;L�$�O���˦�	ԟ`��ٟ�c��^�	� CT�&�?j"��J@�%s�r˓��d̓�?����?	���'���;��5q�b}�F��:��E���ܼ��6�'(��'��N�~�.Of��֧0$�AiF�L4OX����v����2O�ʓ�?�����O���'ئM+b'�=G�ђ�J=��u��Pğ��I�Iӟ@��Gy��'��8�O<q�%���>0ƘCό�=V���U�' ��'���'��'@9��lӮ���O�C�ф��d��P_Xը�A�O��d�O�d�<q�v�ϧ�?��'ڑ�u��t��d�s�_�������?���?��ʞ��B�i���'5��O���U`�9f\\1WcDR,�֓ş��hy��'��h�O�B�'�0���O@aH�F�7�6@cs��3R6�j��'l�I�mV#�4�?9��?�����	�u�N�i%�CEِ����/il�	ڟ@�	�l��Iv��';1�����OǑY+r�Q�F��4���'�̕�Nw�L��O�����"��'��1
�aS�Y���.�8�l-�Ɋl�<���H�'����� 9tc�s���Iɚ_j�=n�Οh�����@g��ē�?9��y
� v����؜X[�18㭞/eܤ 9&�'=�'&u�6����'9�3�����Tu01�D�M�uJe�'B&��JO ���O��O"Q�/�j�&��ujX1o։24I�<	�"�<I/O��D�O���<����C��TZf�U]�ǂ. ~���C�x�'!�|�' �̒�OE,�s3��9'���Q��AJ� k�y��'O��'B��F�6�#��h�T��[+~z��M��*�B�:�]���	�'���I����"�����G��&_����a�C(}Aj���_^yR�'�B�'x�	�^�$$�O|�䣏<"�9�PM�D��a�T�)�?)���䓰?!���B�y��6���Y5�ʎ/���H��?���?�*O�X�q��S�����Pժ�rciIʦ� ������$����ΟD1�&_��%��8-�偔�ź� �8g�.ud�İ<��H69l��Q>����?)z+O�Yk��.�!��Nނ*iR02��'��'n����'hɧ�O��t)��;;	~����3X!Ը���S`ޅ���i<�'\2�OOO��D�2�<��N*�x�c�O�Q0��d�+ ���'��S��T	�%T�	�.�1g�b�`���M[��?���c��Ă�xR�'�>O`P"'f�/[�8��"ͼ\d�+w�'`�'�l��d����'���'c��)�4ey���>��lS��'��>`2�O:���OD�O8	1�ȋ��!#F��K},Q(C��<��?�,O���O��D�<I�LL
=˰|�F��x��M�T�Ę[2����x2�'�"�|"�'����<g�d���)}�QX H�L���R�'�'���A�ō�(Z2�[uOۣ mJ�h�F��'�Q�E�rH�tA�8v��k�L�|9 ��4J�O����OR�D�<Y�a����i$$�L���*Ѳ�d��p��bs��o�)�?���?q��䓱?�0�A!E8��tGO�mM�m�0)�#�JQr2Mܻy(����ժ;��}��eeN�q��1 E�B����i0����� �r���L�nx1+b  =Ɇ�)��x���A��l~�r��Ζt�H O�z2(�k�`*�6�脨�L�,4���''�]ơ¢A��[L@'34��S��8 Rܺ�+�20�D���)3�R�SG�u�Ԡ�ЉKR�l�2!X�q�"��0���������ݟ��0KO�@�	�|JE���iy�B�z=>���
�4.�52�G�$�b�C���K��y⣈�}�6cȽ[���9��Úp�:MӴi�p�J�QÁ�I�,�t�_��O8} S>Oh��4c�PQbb��5�*q�a&&*C�I���M�1I=�*����@�PC�I�z\4��%�F $q0����͟I�>%R0�i��'=�u�%At�h���O��'C�Ԝ�5�%l���)���7<Vy1`�
�?����?IC��0f�-���Z>P�l}X׿ih�S4,�0w�{2H��\k���Z� ���W �8G$(SIG�'��y�1�?Ń�c��Cd�̑$e!��a �n=��.h����Ϧ�bK|����01��Q�b��Ǉ�u����	X��?E�,Of�b([5 �����ǧdޞ�0��'t7m���'ZntZA����03O>i�v�j���0�Xm�����	ܟ�S�Lo8�	��l��ɦm8�b�*�h�D�_�U�FX+���GZ�1��"x�$�(�i�(r���U�'�~��|��H6�ҝ&���p�OP9�����"cҭ�g!ĥSF<��(ҧ�~�B׋KJ����m 	G�jeC�%*4�D�Ob�H+�'��'����f��ch����k�P4R��'����s( �D��3(�tC$�:�{��9�S���i
ִ3b�"�6�	Ԇ
`N�X�`�O
�����x`����O���O����?����1IBL�(h���v$M2���I��T	h$|#R&��T"� "���of�ם	�`0����H>����&�y�q��GL$B�Xh����?'!��o�<[�k���|,j����'XI:�]�j�� 㤈*}�zEZ2$S�����Yݴ�?a-O��(��P�E��	��j����1�!��շO8z�Ȁ��,X�.*Q����4�?1-O�릧��eo�!�vq���[�^��5#2U�QB����?i�X��1x���?!�^�R�"���G`( `l��rS�=�E��2�ҽA���<i�A%�k8�C�!�k�HAX�J��3�\*|$Yv@Ԑm1�1H��
�a�x�$ف�?ְi#�\pVG�54vq�­1ڠ�o�k�D�O�D:�)�	�7g��[AA��\��}W��*�铄�>�GA�v���S�!���mbFy�6�����'9ڶ�l�����O˧t$RTA�ǆw���={t0���?��?1��_) �v�(���F�ѥ���G��S��5�͛Y�0�2�]�0�2m��P�j��`�R�ٸ�=RSĵD����&//����?���J�\N�SU-*;/�OR]K��'�f6-Z��h��+
H�&0sB�8^MH���#�����)�gy�����aF#W�Ȉ2-
��p=�6�D�5���D��\�V�p��U�2�!�闧�M����?���|R����?����?q�4~*0i���!�8�t�S#C�n�q�`��)�lOp���O����Q;�d�����7����$Z�c��-r�K��Xp-�/*�FI?�g}��#�<)����<����N�m���D�æ�ش�?Q�a�|���>֧� ]CSK�0"zlQFeN80A6 �$�Q󟜄�	�o�0�q�\:d:<B��ǎ����ڴ7�v�|bY>%mZ�250p��a��n-2���Z1`��%��^/���)]�?����?i��e,��O���wv�U��i׌G��Pq�GM.��`g+�Fiq��g��ʻ&��7�֦]��0�I>0D$�e���>I�5�׈0�Ā�a�R?�8���ݾj_�	�3�`��mZ4+;@�H�$'�<4������h�>�)�Ϝ�Bp�ȓ��K.��i�Y�`��x�2ᔼR�*
T~-$���Ad�'�a}rɄT ���[�X��Eױ^��mZA��M;�'���˼.g�LoZɦ!�w��4	��F��
e���B�?q���?q�H�"�?�����U��p�;��T��������j؀�E��EU�E"�h�2l�J��b�Ʌ|�����o��S�M�2�L��N
��G	z��Ⱥ`��o�'~8��h&�F(օep��8��ܥ?���xp�3C�[�'"�	����?%?-p5i4.M�q��D��3 9D��:��/M���`�+�MiLt�c@(C"f��������m�0�x�k3��O�P�$��RD��1��)i@ ��F�x��)���&nA,^�V/q����82Ģ<�ӣM=!p}s�̟Q M�#�CylĮ\ɚ�A2]&a��CI<�y$�)c����S�Ѳ
>�y�n�
fo��H��ߧw��$��3�y�D��,�(V�̮e��IX����y"	
�p��[T�+\���.���y�<At@"$��*Q�aC�,�y�X=.��V��,S0�X25���y��5cޟO��(s%���y��Bb��*�H��?��i��A��y2�5j�@��w��`��Ԯ���y��8+���G�ݑb�D��I��y��
�_O�`�&�"d*�œAF��y"a�d��p���>�j!�5�y���
/Z���F1s�R$�+�9�y�d�r�
���W�jt�I�oH��ybM�RPX9Vi��m�0����&�y���4��r��5g��t�0'���y��X?&����Ƅ�x������y2M��21T�r�\��ՀP��yr��R�j!��h]s d�ir����yRDB8W�~eHe��|�P�DGH�y�Ø�J����E�o�d{!�\�y�i��H޽�e	�5�Ej0���yB�^����2�*>|�M��yb��v,�k�$�j������y�J�YAHI�H�2��jDn���y��Z�`�n�;��1�>a�0����yRLο,x`#Pd�!��z��M��yҍ�l@�E	�H�3'9̘H5m\:�y�,��3����O\�9Y��L��y��S,~,�}�Q�+��� �E�yRMR"�4Pa�����y�ph��y�5:[b�1d[�|���aʑ4�yb��W̺h�U�!O?uɵ���y��, �#���3;qV�IU)��y�C�#L�\I6���2W,$��X��y�H��Ȁ*+^<����r��yT�9�؃hE0m���x5(�2�yb��o�=
����\%N��W"Ob��ˏ6!�ɪ���+6�(`S�"O��	rB�1�6<�'B�Վ��"OqW!H�D��!Y�f��z�T�U"Od�!e���Z��`�� 5�ba�"OpxjsO�?I���S5���6*�`b�"O�e`�v�da#��*�1p�"O�G�W�|��@�[7��=9A"OT����@7T�:-�P�P�aDx��"O8��K��Y���1��M<��H�"O� �%��oG����;�@SP���"Op�PA�]s��3��}��lbp"O���J?���T+���6"O�`�q��X鰕0������q�"O41h��Gu��D�TMڮV���"O���)��D���d����~x�"O�A+FdJ+OB��r/ͼӦ���"O(u��K���@���Ƙ14�1�"O��D��C�$� ��:?�j�"O��q$&�_�`��ueU �0"OP�#����"�υ>�{�U�X赏�},�5��	�'M2<�a�I,1o��@���>����D3^�<�S����4�܋ �0�zY*����WX��p�'W��˰/٥;q��9g�N�J�>���d�aע����It��?�WA:4y��A���.�
�b�n9D�X�"ϛ�M���_���y��ʬ
]�e��d��i��<-�~���BJ�p�<ƌJ2�
E	�L(D�����̋a�ޔ�A�!	�V `�"xӰ�YQ��4�Yy�aT�\���Z]9�D��v[af�]�\��z"�Fߒ�;�N9nd�����,���iE��:w�c��B�I(��|�B�ɲ�֍�T"��eFO�����	��Zt�f&J����D��B��Bc:^ �)��
��y�DKNa��q� �W5��#Q��"[O�и�O�$A5cX�Ѳ4���t�?}b,�w>�s��5@q�@�֣�0?)G�Qb�����"�p�u(	6��&�EM}@Y�Bυ^��CA(k�^�񤈾E �w���g��U�&���-'ў�0��F�D�Ж�X-i��e����$�pA�e�<a�$KV%%h��]���
\2B�IJ
P����o"\��Q�=c�7�1���Co��gǍ=(� �����6��k��4����L٦Gю��!J�`�!�4k>�J`
L�:�9ad��w�r|�� ���|��,��J �"'ڟF)eƂ�f����O漹b	<Hb��#K�=GV���'(��	�j�z�x��g V(��D�UX��y�"��
dp�	�a�HkFY�hZ�*&��򤆱8e@ؗ�ˬ
�ȳ�'���O�hp�bBfz�� OP^*
��Ŏ�B&2�xfg.n8�h�9u?νB��!�X�b�'��H��%,׶di��_!%2���M�xU����
� ��)*�#_Y��t�w�-Ӳ�'!��.��AB�c��� >�"T��dÍ.�!�ϐo$ ��+
�f=K��I���0�0f��p���0b7�x���0�a�����2���8}"�b4) U1Y��!��X���=9f���8O (��ן+pu�&dA�;{� ���I#	L�$�W���nO��C'O\�ҰDO#}tax�@� n�YD@�p�x��͗��'7�$@cE��r9"��Q�Ђ~CZP�� 0P� ��B+'��1(U�s�J�#�L�#$�Z�,����+�˒���l��}@4�Ć�	�D�YA�ȝj� R 煐iDz��@������,�~Z"3��S˝�X�A���nyx0�"O����뜖�H�E��X�KF�Y���I��� �"X�|��h�?c�뎆�p]pS��I�2Y"(�'+�5����ra6�y�A�33� �8K<t���#�HT��o�]'_�3PD���F<Lo���a�+w왁��|T`����'�x1���hl���_*�6�}��&N��ț5�ǿ=r�A)�yR�@��l�X�v�C�d��XT�<�pa4�����97H�B�	*k�$�.��:�DXEN">?:���)�~�\���R��#�B)m�:$�U�9�@���ۂ'���l^�,���r�LA,%�!���@�rg�M�]⦔{��\�e��iT!�#u��|�En;B�!&��i�2�\/0Rh��@~�a4[�.a���<aȶ!	��=�g��&(>]1��o���[���qJ��Q�LU4�����*�8D�iW���s�J��X:
���?�$i��W-r�����e*��k�x��yCJS'
�``YD( ��$��gIQ�5�0}���J�+~���N�k�|}Ң�98���Gz؟���Zǈ?V���"����A�`�(���&r����M���$bm��7� a2w�]=R���:��O�h�&
ߺ�1S
�O[��Z��&(*C�<0���+�2b�.�����E���Ӄ�*k��%3�(�;<��%qt�NF�S�b	3��p��AC�8B��$Ȝ �"�kGM�sP8��.
�~�a{R��d��qY �p�1y�dY�gt╀�.}�H+Y!kF�����ƢX^�"G�7D�1���y�')�l�΄�S	�����B&MT��N�ح�?6y�Њ7u��Y�*zt@����%
��a3�4>�(�����:��hR�X%: N4r���8hI �����y/"�3��W3X����%3O�N�gBC�d5`�`3%[(ZU���|"<�o�,m�Tc����g���;?�|Ӄ�d�k��]	�z�cV�>�O����'҂� �\3"�*�5�F�L�% ���7.�ȩ�B�#k��<��$��L2s�L�!�	ږ�!,29Q�'V0z!@]T��UI�#��4���䊆C,��
�)�x�Pa�!}�D��>�|=Y�H��_�RMK�G�b�t���+����N61
jkF����O�9(!�R)>���'
~,�6Oȍ �BS89x�|ٷ�k�P��]�Q/27-�/�Th�#��,��ф�N���L�!b
�n���PGKI�tR��'��`�MWo?�@
2��'<��U�h�S�jɐf�$!�M�ë�/�
�X���l:�HbA%:��}Țw����U�/$_*pJe���8:���	�99��ˁk��Z���*ԅ�P���l�4+�%P .H�4�^i�`-��O�~%hӂ���{cJ	�N��4LW7/�-@ n�=5(>�3�٣!�ڴ�S��6ٔm"��D��l�Yb�H`�����Bj�(%a��9�(�WI��_��B�C�n8����M�~� 8�U�-?\M��C��;�)���'�jik
<xQБ+�G�&��x(޴"�hY����w��1D��V�Xh��{����O��p8fꆑG���1NW  q���)s�劥���`����5N�����\%�Te�tH�s��ʝ�;���)��5N�J�@�G
���£X?M"�bŋ?Q�P�Nם@��6�X�:�XH�Ê�i���j��^Wa}�U�&��8S҃>D��hB�nC#.�}"bDS0��;�kͥ"�,X2�&B�y�#<F��@
J��HCZ?��@>A�.U1�O�#e(�A5��c�`^�k��$�w	E7x-���26 UA�����6�+��	��0�e9m��Y�>A�*�g?�h�]F�1��Q�G+^����I��kH;6��&�(���+�)��9���C�#,�s��!Bȓ�=�J�����v��O8m���;���Q	ۓ+�^YY�Fȝ-��`2���=k���rUFj�����'�j��@~�4��T[>10�_6��U�I�����[	4���8�Nw���D�u��X��_�-�T�w�O݌��"�v쐐���t��
�m@�x	#�'h s�i�����N.������ۅ̖|b'��5�(���E�
km�Y���I�=4� 0�H_1\����֦�lz�C��:JK�L3��3%��� �GʇW4�扴;�)kΉ5p�P05#�;KI�H;��	JY���ND�B[vݛu��!=!򄑰]��P@F�'t4>�U� �W)-�jϦm�F&�| ��$Fx��Q��"�)3&��غ�ց��p?)�*B�E�DD��añGޖ�#@.ɩV�UB��,03���:��>q���
Y� ��+���`�k�'��H�2�Q�s�t	�f��)��VS ,�4f�?o��YD� ?'&!����R�N���Y���P��r�	�_�pq`b�=*�?��5���R�H�`]�t�r��g'>D��z��U�X�c#F��uX�;L-C.d�@�'`� `%P>D����Ol��H�2&�P"��B�y� ���'9��x���FD�����I�"ZM���ɀ��5��Z((K��9
�B�8�!�.�}V�ԸvGC�{k�F~�	��v ^���7?.�K��N-�� �;^�:�h�,���f"O����EX�f��!z��X�k�հ�[�<�%�!�4�0S�G$]SP"�UC:q�"����(2#Z�
�'C|�<)�mޖT��ՠW,D=��k�%G��ui�;OF�1���9��i&>c��j4�ܨ�p��rMFX-.	���5�Ov��h�;q�1�K۶I|Ur�I�!2]����
��y���''�[A��#M�X���Դs���z���
XRI"W"�3����e\?u� �ʪ`�6��!�C#���=D���V��tu��s��!-`�h��<y�O��]È���cU-��?����MBB���C�6m�����#D��*"�׬G@�0��bѱ7����ĕ� �~�bl}�c$	j�g�Y&�mC��\>l[j̫.����ܰ����X�7���(���b��l2�&�::�ic��'2&ĩC��$5���/�<z�
�In(�R�ɯ,�:d�SC÷Nƶ�i��Q8k�B䉼p�@�Z����ltPW��#I�HB��(�v5�v)�0��:򀌋q�4B�ɻ�tq��-=[�P��)tC�Ƀ	�!�7��"fo�\A0�˾l�2C�ɍeh��pV�V6R�ht�"�FQ�C��e�b%��pv\�`��A&�C��
2G��(p�C��!����TB䉥��5�&'1i�Z�	b�T.o�B䉩�X$i2���&���+��*L�PB�(T�V�	6+*w)�,���E}< B�ɵ_�޽��P�Hb�z�q�B�I�|4ℚ��U�zG�0��I�x�C�)� \l����:DL0	s�Ʀ2��k�"Ofu��)ƮHzh�bÄ6�"O2���^'}hxUjC���v=b��a"Ol�+lϵ	��� +*�<i2"O�ie �,�P}	�e��%*���"O�p�A7]�M��d�t��y�"O�fC�?r�e��bߍk�ʑ��"O��i�J���4:���8~�f�"O�P�k�*�`U��v"ą"O�t�ah�<�� ��\�&��k�"OD��o@�#�,�*��S�6��"O����2&�걁�I	����"O䌀���Ḡ�Je/�<\���U"OXtz��$6"�����|�> ,!�D.���i�L�>�8pbmF�d+!�DR�)3�l�qAZ4���We�$]!�ǾA�t�R(�7Q��5B.�}@!��4�l@��7RxL�"mC*~�!�DJϚ���{ȶ�A�6:!�#��b��_�i�,ہ�J�Q����@C���!�n�24�q �<�3�ܐb����wi�M�t\��z�<%�I�6�T�C�V�@(��[Q�<Qf�W�JaI��_ܒi�
�s�<��*�0%�6��-�:V�B�PE�s�<��IٝV��*tFR7h[�t���q�<�+�5������%�A7Fz~C䉍\���{ƌ�*E�dE)gH��zTC�I�U�4���Ϭ!�p�1k�#C��C�	�<kJ�R�`B�^10�aC�G�fC�I3rl�Q�ܪVV�����B�I�P���#F��&��#@B�$�XC�	���y"��־u�`��	�7�C�D8|�.��)���g��	�B䉑`�E��F���ɢ`�
�B�ɊK��e��bɑ��y;�M
1^S B�I�6�[GOW�	
���[r,C��< \pyg�ZI���'��le,C�	�(D� %a��.Ѐ����$l!C��&O�`�#�fF%���"0�6$��B�ISIȑ�Ӌ�;�vT����E[B䉑#��0ѵ�Ϙp��@�]05��C䉋o޶�����Q<�p�Ձ6f�C䉚�v����	��DQd�^�dH�C�	*(ƶu� �&B3&��ɺ<��B�	�y3�i���^3%d�BuJ�5W��B䉼_�DLy�)[��u����I��B䉜As�E��Q�(!J�B&�P��B�w���E�Sx���*Gn���^���Z7���2�A�%CX���,�2r�@.�8��k�0����ȓ�pU؂o�h ���#dצI7tY�ȓz���&����
9Ҵ+��A�z�Fz�cE���Uۦi�ٴ�-'����FR<'v�d�]<m5`qnZ��xr��0�$;��2.�9B�N�H��Y�<)��½c�\@�c}r��M�Ͽ�'BG�~a��냎YTN����+�_�<r`Y�|ׄH�&oK/kf��9�冗a��dȋy��w�"L
9�zX1���qy��'P*�U e��K��P������p>�F��6��`��D2�L�#�k(~E�!S�%�s߸� g�2<v��SE��:�[o�'j.��s��Q�j��
ʩ�&�ȉ�d��\�.��w��-`j��ډDw�I�N����D��"X��j1��q�b�"�K����W.P��|�0��J�҅��P�H6�L�^����e�C�*%5!��"�L`~J|�1+
=��'	Ę�@��qƭ�ȓ!�l�:���8~Ⱦq{���L,Df�F�#1O,E�~"�(�a}rCC�<0�; ��;+g�)�������	E��x0nij�� �Qf��h���@���_��̈D�'�&H��|BOQ��~�DD'*��0nVD?�")^��XHP�M�v�jTi�*Kv�'.�e�&!N�J6HIR�E�36jUk�O�����*rf�:��Y�[@��S��O ��&oV�3��4�L�5a�����I�^�	��K���\���I��0��q'�0{��5(��ܥ8�� Co}��@+��$�>q�Eɕ3Z��+�'�}H݈�%)'ܔ];��=�$��q��v��ȹt���J�`�$����(�
`��WGRV>��R�PD��S�BC�����I+C�Q�JS�Y-�"a��.%0ې�>]�5��щ:���':1OJ!b�)	=:�Pi�	�S�����'�ՠRH�*�D��ͥ|�Ri�I>��݅<oRh��iJ-j�i�6F_}�V����k���	�@ӑD�P�%���\9q_0�MK���B:��E�'��AB���N[��ȋ@)q�T;�1갭̡-�yB�'%Q�8���ޖ�c�M��[$�\)%���eYv����	5Z��s��/.Q�!�;p+r�	N�'q1�ހY��:mqXm�e�Z�L�w�9M����w�'f�M�s
�A���s�Ŷ^�*��U��)c����H�*
���R�m_��:�j�0��K8����^��*�$4|��ѨWL 7Q��� G���'р��$O�]�@��&�:E� p�O��;H\<�R� h�(�B�e�Jh��ϓo��	�ڴ(��zDM�;���z��	S6�l��!��T�T�Y6�Éq`�q2a��&,��9K�Aջ%#��,oک1��d��|l*���X/#zP@d)��d�v��î��o �}�&M��6�#5KIaD�!$�C+3�'��'�qO8��6+]�S!���\�;�Q�	�^�ܒ��'�)�a�&�n�A�fߔH�XeJQ��Wi����H��X?��R-O^�dc�|��R�+E�E�8�61�^w���P��'8<8��'����c����� �}�K�'�T���ăK��&n����4���s0ߵ�~��ĕ.4�(�s�n�\�u���MӁ�
%7����h^�'�yQ���S���L�'s<z�E�7%� h8Q��0I� x6��A}���ɡ'���rl�"� �9�A1n:[p�K%�VR��}b��d�21+ $�,JB��v��]&:q�`�dP�O�.	Y�'Sv�.	��d�+��+��9*��z�P�����2<<�#�MK	��Ɠ#	 ���.V�9+�M��K�}��`a��Oy�g�y�tc�{>�"0O���td�L�rQ�#�Nd(ѣG��:t��y���8X�$��O�M�����b]�x�p�V垇y�|1�D��\��ĉ��צ��4����1��$I�l� TB�N=xa��	Œ��2�p�Ћ�?� ��T�O��$ŜV�F�3LH:&>�\��	#"R�k�`��p?Y�MI�*x���� z=������Y�E�'��Ey�O����0�hP�BE1-oxE���&��a��'�~i���;&*hQ�F��0/��5�g��&-���6gH
J�O�oڠ~B�]���&������kݥ��'�2lyg'(�V�ԋM8/",��MԠe�<d���^f�ĬF������*���ڥ=�Բ���I�p�oZ�V�@��o��tTQ$�.4��>��Fj3�E�v�F�&=0�a��+J�� �2�N$)7l�i�:6�0�ԧ��}re[Bʐ#�@l�"ٲ���Bl7����D�v�Jx�l�$o���W�R�aj#W� {w�=��?��G�����"�y�;L0l��/X10��{��~�7��U���Hǋ�&�Y����Ƌ��'֔�z���,a	t�jUcB�+2� 8b�����7ݢ�vdBT�����1}��ؤj(�!G�X�44a�K���'_����g^?rL�Q`�N i�@<���ڬ���!Ì%lD�B��0<QV'�M:��Hs�ŀlN͢c��!%��Ӡ똩t�X:���,�D�OndY���_Ĺá�׏=��#��V�h������1�Iǩ6��
r�Z>v�N!�c�$[~�|B��{�0���3G�,:�ڥ��	�LU"B��x��X(V�"l	Li��A�8�¥A� �i�d]$�FN���0�I�xu¤C�穞$�$�
�O�8qf�2t7�)�Æ�=*D�r�0l7�9sb�4��(�˖�}�D�U���9� � 8��4�3��%r��I�#�`�I}��\@�'��`y���Z��+��A*a�΃�M��@���0���P�X�GQ����u�O��O�H���,M�D��G���h�G
��Pxb�I�6��P��h��6ղQK� ��ei��<�B�I��MK���yw�M�$�(P������
	��p>qĮ�dD�hW�P�e~�(`σAK85s,J<oE`�<�RF�%��*dǓ!�84w$Z�?�	�%0pj���J�yNT�5("<I��%<�Ja���G#�"��� �H~�E�C����I������ 	v�X�9���XD�HTL� ��Ab�ψObu�d�3)c҈�59}�F��,V'68�6.���P�ѣd��9Hb��?�O<و$H!#	�)�UL&>�C�ؖ�0������>aP5_2�h*�������� F��'��Gy�O_
��1D�
E�j�%y<(��@�w�jĳ@�'��<����Zq,�(��tki�C�y���rdl \��-Fy��ɂ4�h�K�9$��p`d ��S�? �6 �C���a�1+J԰A�K�JղE ��!�R�8�Ǒ�_f��N��3W�V���BuB��u�����<)�� ���Uo�h@��G��aܤ2ׇلGn�I���Y
��E�3��L�u��4�O��3�$ɢ>�h�.* 4+D�ۻd�-��'[�a���أ|��g�ST׸�6y���M�2@<�IW�Y��4�C+̸~�j��k�#C��B�'���c���F_y4Z�H�,�[�
�x�NF��p7�Ũ$M1O�p3��O"9��@���b�i}rÐ�`]�I�D�U4�Pڷ�A���Yj����|np��"{	�����>
{v0�'�J�[���OҨi�`� U֥p��e[�&Hv��TmM*W)J�E}�Z�E#<��v�GR�Ҷ� k�tX0΃.���{�(U:Mp� ��'��46˓2��2�l�>WČ��o��I(XU+'Ɓ3Lv��D�3}(���͡y&��R�6tRy�Ճ��{z^�Ud*�ɉg���z)<��E��5R6���&ʘZ�y�w�D�H�㉻h���Ǒk�4�&M��M�
��q�Uf�F�J�
K�w���@�>��T~�#��p#Il���0����?QW�
Q�`�	0Nw	���gc\i�d�n.��Hw�ވ2*�X�%��r��^��Iu��غ+`�V�b�,�!eMS�"�Y�����9�b�		+z����60%���+B���=��e�cE��Yf$.U�udٚh��P;PHѻ��@�޴B�,Z)�ʺ+�\�T�'�Fpµ�V�'$ �b6��q�z�2��(+nDyF
��p>����8� c�WhIP��� �Jq�㈇3*pƀy���>QP�i�q�瀗a!������X
�d�rJ:�*���	�g��(��u�h�&BH�l~Ƶ��)슒���A6�a��cL+.���]B�
	�-;lu�P/w����êt��-P���>}a0-is0}�j=:BaY���C�4xZ��CZ�òv7 ��œ7)�:��u
���r���|���k�н22�<�\�aƋ43���DzRƘ�+"� �+��=x�c%��I���$�N8�i؇oB6r��VΈ�k��7��2�;y�����d��R!^79��0�Nqb���4C�i��t��I�yrX�k���eb�4Ϝ9'������6�\��S"�0s̘q���x}�be���OQ ��Ѯ��
��q��V�j隰aK����$��nŸ��3m۶N�*�SPi�)}��*� l���X@
ŕpGM�ֿi�`���OH��昂��ٴCаtkCk1��Gf� #��͘rf�q`
�V_PO��s��$zm>�je�\=$DڼW�i�قF�����IO2H���n�

T�;2Ɍ��%� �@��~�bϱ	椹�[w�`��dY[��	��I�m��hR�9�$n�A�~!k�EM2�M3@JN�%�l,8�O���U��!���P�t#�@F+'˰mc'O[� 8�J3�!�P�p���Nۛw$4}8�GU�s���0�
�Q�4�xEBç�T9�7��`$��'$F���ꅵ62R����P�RK[�sM:��-J��y�D5O�4�d����Be���^��f8��GT�a��Q��-Ed��ӆ �Ʃε�)�Sk��Y�����p�w���	17a�j&�i9��H�T~ �aWK>}�(B�Xa|Aҟ'f&�RŔm�2˗���Ԑ#�'�@i筋�_����V�'O�űݴ$e�T���^\�]����O�H��dK�)����� ]�MGR9 voV=@���<>�Ф�p,�d�v��I�i��CH�<��� �ZP��E�Ӥ 18�x�'dO(b����Dɜ9hI�e���<JFi�/r��9��O�X5�'d|�w(	2����eG�`ay��>8��K��'A��K`a�*|{�$�r=&h�ri�?������V�aZ����PWy��xb�������g�l5"������dF;.j:|8��G�6���Y��P�r��'{��[��@ky��Ю_��˓2Kf��Μ=b�l��G'ˤ&�PX��C"���!B�V�?��Mh��E�:% ��,�����g%��#Ƈ̥$7�1�䖟�B��In��_s�͠`�$?�(����<�W<n���*�7Lf�0��!�x��D��1�|�Bb����E,o�	�) �`�KZ4E0d��$�O�}_�7��O�O�X��ڃa�2���-�4+��p�'*�(PAB&(o�i`��� 'itH���"5�$e���&ɘ	r�FP����˓p&u+R`Cd�Ω���9���ȓ��&-Hnrq�t&Z�\z�5�)�zqa����sQ*�з�'	�H#I�g( �BiH��N��:��F�S�4��]c�h݋)V�BsM����}b��6��$�Vl���ɀ�H�l=��ׯ;!���t�9UȌ)I]��ѐ�Z%!��> ���b,ůhS4�b�U!��T�f}r��;����̷*!�(+٠4���Mq���!���7n!���8b�|�J�iN�t�H���H��+�!�:�{t�óh��x"G&s)!�$($mLl{D,��-i�t#�#�	&!�	�b�1���4�2�",S�!�$�*7����@�6�pU�I5i�!�S$nPV�"�C�P0���� ��!�� d�s���K�ʸ0G�R T-,��"O�m wG@8��R�Z�CJ&��1"Oڌ:R�6I|�0I��ʙKI(�"d"Oib�k%����dF�V2xՑ1"O�k%bL�#�\y�6�>����"Oĥ�q"Y$_�^��$��4#$��"Ol��ҪT�l<H�����y~��8�"O�يW�@�yU�p"b��~�Y8�"On|җG�8�dh��A,5�"O���ƜD�t�`��n���3�"Oɘ�/J�T��ӍK 2�V���"ODh0 ��6vv��1�O��qԸ)�!"O�]��n�6W٨<�J�i�:�J"O� ��o�34��][���"Z%@"O�а��6��t#��4(F�1D� �hP�f��4p���85̸��`3D��*���ԡA �N�`�N0�7D��	�o
&H0�@dJ7f�X8�L4D�p:#�`����EA<�0D���`�</H@�%N�PM0؊f�.D��(��ٌ;?bq�L�j���Ei+D�܈�Ш ��Y(�"I$-OHu[R�,D�u�,Y��=�wl�-�J��sl,D�ԋ��+@t����*],8_<�cg�+D�T`��k����5E�!�T��i*D�d��G�7(���L�=Vq�'D�ȓ"��!"{
(�%JJY{�qp�$D���s��R�6)\� ��eX�B"D�Xr��٧u��tA���(����gk>D�H��Ŕ7���y5>S���0�<D�������Wٓ �e�FG��y��C�eɞy��'&�4��׆�;�y"( ?1�vQ�2�ì#����!MQ��y�F8CV��J�=1�� �+�y��vn�Ak��ʺ`�(�Ɯ��y�᏾'U�����.Ɂ��=�yR�<L/�+� l�x�-K8�yR�Q�@y�SeBb疬8Co��y"�ʜJD���0���Rqv���A8�yҧ�Up~@Q��[�=7��NK1�yr$�*���w��'��YA�����y"�I 6+l�i�G�?o�^໖≰�y��?�z���'�f������y��2Z@(��(g�B�)sID��y2�ƣ@0P6oO
c�����S��y�F���A�M�p��u�A�>�yrA��	��E{ViGm��0QȚ��y�d^�=.�a�4R����� �y" M�3$��3"�y�R���.�y�)D/M��C����}#��fU��y�E�CA>�[,��#(�S�-�y¦��'$�d2Ҥ�ݼ 3]��y�,'β�`D�LD:U{��?�y򎒐�\L"#-ʱ5opP��.��y�iH�|*@Õ��1+��l�ѩP��y��چUR@e��P�*y��b�*�yB��=T��R��4&��������y���c9���+K$"� �Pe���y"�	�W�8��b�
��EM �y��J/�&��Ŏê��@����yRkܚgn� b鏬~
j(*TBF��yr��"�T"3�S$o[��6Bȉ�y�D�/�	����{��HZa��9�yr���.+��1B�*$��s�b��y
� ��0#'ʈ_xё7䊦Z븭"�"O�4A��[8tnX�d�\2J�+�"O�}`�-'.����!s�N3"OҹjU��$0�ȑa��+`��"OPiZ��-hn�R�m�; N�Y�"O2`���
�a� L36��f�	�"O��rc�I���ĉ�e�~��"3"O������-]Ea�*P��Ea`k0D��8���h�6DV� Av�(P�f/D�i���|�j����FX��.D�p�c�� rA��ʁ�$}��5Q��(D�D(c�(*"��"�,̓yʘ!��$D�X*6��/`��F�=f����B5D�d��/P�g��`���(7D�l�#�I�qՀ<x�jC�x��-{
7D�����&z8�L���23�����F4D�T�e�=4}0��[oPt�#K4D�0���W"K&4�J�jLm=�@x�'D�H3Ǌ�6"F��rH�7>>	D*O�푱���t@����*M��"Ol�g�G�����DBːB�HiB"Or�K�g�f�`��d�0M��8p�"OtX9� X7h�<��,���:��"OM�� h#| ;W�r���"O��xL�7'����T�d�xw"O\�:@�S�`$�a�WE�ua�"OfY����:�t}�%�%;:�8"�"O�� s���0�����"e"�Q��"O�P�ꊧm���;��®8{�@c"Of�����!���1���>^Ir�"O<`q�ȐG��c1HU E����"O:]cD��T8��d �$?j�)�"Ob����,UhS���w�@LS�"O,��B'o�(��No�)Ig"O��X#�r�ݐ���=xR��w"O�XJ�c ds&U���D	^{h(�P"O�][2b�,+˄ȇ&�Z���"O�e����8�$�ȧ{c�lY�"O�ʅ�D�6�h1HņG^4B"O��x�G��Jv&�L��b�"O�Җ˚�;9��z�e�"M�l(@"O�#ᣔ�"�4�ċ�NOP�`"O�i0�KbH���w���Ei�4z�"O4���De�Q�7(O! �Z�Q"OD�Ẃ�^�"�璢
��w"O�z��B>@ &������C"O<���H֟y2lq�犂����"O� �E:> ��x��װsą1�"O<��a�m�$����D6i@aS�"OQ��j�
E�Үɓ]h���"O```D  �&��d��L<3���V"O����a�"p�z �L׾*v��"Od��oZ7���i��[�RV"OD4�q)��0�m�i��e�u"O�@Ж��|��iq����1�#"O�1k`F��@�5J��ٶC"O*�{T%V�U(�|���Y�`��x��"O8-@��ތ����f[I�8���"OP��iY�_>�}��R�K��uj"ON���64�H����{�f��"O�� ���� (m�j0Hs�"OL9k�&�N႑ȧ	T� ���"O����L�':��z$��5����"ON��&lTO�u#����D�s"O� �`�P.M6s��E�7;s,�J""Oڅ�T�<�0Pa ��O����"Oj�x�)�+�ȉSa��$H�ȭp"OB@k7)�>���V3k�ܪ�"O�5Z���/��6�R�y>��;�"O�Z4hͫ.����e�X�a9�"O\�°�ǿD/�*dW�e�\� �"O�hQ�6h�����Ð&�X�"O2�b�O\j�l�)"��,et���"Ohx��-B�,��(�U�"h�Ur"O:<�T�T-;e>�Sa	S�0���)%"O
�S�)��D��V����"Ov����8[�0}k����`��"O��۷���Rf���Š��C��{�"O��Ɯ�V�6�ŀ�mHVV\q�<A�h�;5������r�蒍�k�<�sk'B�DK�*ܗy`�9pq�	|�<ySc�S8��
J/"5��[��C�<	�ǚM�~��M�-�:�k/�H�<i�J����Ζ�Tր�{�`KF�<	�OC�r��'�BJ��m�$�z�<!��["vb:!��L1a9��j�i�q�<���;k�^�� O'i���*�����x�Ė�U��HA�OM'|� "Fm�=�0=я⭂
sv��Ё`)��Õ!��y�l��
b��ǯS0�����JP?�yB$"S����	�2�hv�C�y���"�ە�.�^�� ��y��y�p�r�O-j`q�oX��y�.�⬥��8)6�Ť�y�!������:iB����@��y�L[�7G��� y8�3F�	�y�	Թgz~9���	}�dh��ϯ�y©T]F� (��I�&!eȋ��y�I(@��"KnP�A����y�-L��,�BflSn䶀KT��y�LJ 2�@ f2��Ңb��yRc�'(ب�wÑ6c)��.4�y�O
6�]�$-��H`�aD_�y)��tt1`�
GRl`��8�y�/�8]���� �68� ��-�yR�ծ+iP�E� 1�0��J���yү*+��[�0�����Z��y-@?R��4�0�Z0)֥�����y��ѯW��{�	3P�䂓���y����
���(&��*9\�­ �yR�Pa�i2���)��ZR�S��yrD"`�Nb�	S%I�l㴈��y"E�;t���S�)7�Y�sF��y�&ǩ}עL@Cf�'(�6�3��N�y���=�
UR2'?1h ��Rɭ�y"�ϓ$ �R���r:�m�J��y�g�]Q��A�o��<cq
	��yb⁀)uHa0 +$� �;�H֑�yBa�0c-�	�Šݱ�F1�u^��y�@J&K@R���c����Ä�0�y"���T�hI"DAƪp�4����y�M��V�1B뗪�(TIļ���f���0��,N�B|��m&0�͆�lWnZ�ĈogTM�Ɗ�)�r��ȓO��#I���]c5������~�u0�B+6�2$��P�'7�-��E'�|H6�F�o'�dᗠӷ+	F؅�z��1��T�T�@5�E��v���S�? �#m�pgͲ�j�D�~��U"O�hJ4�4G�td��M��[�"O�� @̩w�\a����mo$��D"O,���m^�.�b)�*
�x�'"OpU���B��AIG�F�z\�#"O
����CKi
�Gː`����"O�\�3�Y<���ʃ� >�M�t"Of	�pN�Lo���gm�[!��B"Oҁ�4��:]���`�B;v
��+c"O.qQaV%��a��ƚ _��g"Oj�`r�Y�j0q��&I�%P�A�U"O���uŇ�t���k$�ïԆQR@"O4��r�R�ST�A�iۤj󆩲"OKF�W.B���)�).����`��=�yr�A�Pk�YJ�n��)7��@�A��y�!�	Y5��Ps��!����kB��y�$R�n�� +��"���A%�y��-*�x��O�(�� ����yB
6�8xpu�OSi6��gP��y��i��J� �yH��x��J)�y�`G&����%���|Ul��.�y��ՔJʺ� �,���u;�E %�yb�؊;�P�� 琍��P����=�y"��$�hm{s��Q���"%5�yR�7r���2��Z�v��	�=�yR�*Ul4ԩ�,T���d�9�y$W.h�8���g`�J��F�F$"=!�ۂ7�D��:B�U"e@]�q!�$�-
�jD���\N�ȁ.�[)!�$͔'���P1�|t��Tǜ��!�Ǔd�ZA"P"�� C'&N�K!�ċ�PS0�z�L�V},���U�Py��+�rqh֣�9g�ZtB�	�y�!ߺ@��Z�%Ȋ6�j��'0�yΛ�^�h�.�ڐQ���yB��#	*� �o�+I�ѳ����y����a���	�-�I	Cɱ�y"&�2k�%Hh�,1b�C7�ò�yU�Ć���ߝp�:q�B�<�yEF�-�P-	S��xo���ƃ�y��VRd�Yс'E=���(��y,ǷE�4��H
D�v�#$�y�f˱=�2jȓ6�J��S��y�
Qq�����,����I��y��TY���%H� �p=2��I�y2��"4.u0��]>�����g���Pyb�۱z�,8" n�I1&�Fe�<qc�V��4|x�`�Y������d�<��h�\�I�6�2����H�<	Q��$�V����dȊ�:�,�~�<�C�>*LL�#b!�`��d���D�<�7E� a���Z>W đ��Y|�<Ib
E�fRF�!�� 6��;)IQ�<yV��k�\@���͝
�T�UΏP�<�HC�'���I�΅CY`� ��K�<���R�.�H�e[�j�Z'��G�<�UN#U+&�2B��r8����BVZ�<QfDGiE�����o�V�jP�<�RQ!��bU�,-�t)��N�<yCh�*��e�"�<Y�$)�)K�<����0����!/��4)P,�q��C�<� K�cJE�t�Ɓ'�q��A�<a�g�;�6��n�f���-Ip�<��	'�r��Ĉ��GF0xRa'n�<� (p��W'L��m!�� ���@P"O�����"T�A��>*�HF"Oƀ��?���Y��C�(�Ҡ"O�����T
gL����"O�
!�èmѸUU5s9��Q"O�%��&ȫa.4�!��ؠ��"O��`�R�To�Y����:#��"O���ďȒB��T	r�K��ժ&"O��"�@�1!̰4y�A����1�"Oj)�gl��.���r�C�s�k2"O��zA:a�ثŃ@�`Ar��6"O�!��!�<2 ����I�p#�ɐA"O�U��j+��̫�%�X�}s1"O��o+fH�&D$�r�Ĝx��'�j%b�
٤0j����#m����'\�E���RZ4�P��ʖ{����'r
�Z� ��	��Z�(Ć^�Dp
�'�ht㣆U�P%��ңa�jv��	�'ƲHI� �xtA	�[Cl�i�'�����I^bՠ���,_�	����'\jR��9MD��re�! �,K�}b�'�ԹY���%�F�p�g��b�`k�'
��z��2TBz=H�EX�)�����'� �透H�:JD�Ҧ�"�XȈ�'eu�UD�/0+�����(�'���)'�_�ԤiQ'I(�Nщ�'���V#�!eh�jC����R�'Q�ݨcD [�6|A��.|���Q�'O)�c�^cSbpKRF�*y��m
�'�$aa�eK�M��}(w�_�[L�i��'!�My֏��m9�!��Ǐ+M~	p�'h��*�Ο!�����Ca�Œ�'�a�1j�;rlap�HP	J���P�'=�Xб�M�!ٶp@q�ص=F��
�'*b�W�o����Gtz�'�P��U@)%�~ųO]�x�
UJ�'� �L %@QȄ�\-z�LU��'�RysE��3e�Za@�f>��'�u�W*|%����M�F0��Z�'���p���	O2 ��M)F���c�'k�<�'�7�	��B �`�
�'Έx�2�M���H�|𨕂�'�֜BSG�w�������$%��	�'��h�AmQ�Aޢq��i	2d����	�'	�X�� ՞l��ֲ[J6xa	�'C��{����^�C�b#S����'�Rec֣O� ��ڃ�̨My�C�'�н�cE�+��ʣ�KG.�H�'!��a�g�X̜��c咬Rv0E��5Od-HCSH0���8m\䚆"Oʄ��耇�L�07,�]��j�"O�1+!�ŷA� ��F	5^�["O�ȠW�ſNC��"�	�<8�pa"OH�ަ"~Ja�a"�<9��*�"O�4��V���6�8M0p�"O�%�	PXx R�ʇ>d����"O�`���Ƨf�4�Po�}Ef ;�"O|i�p�
?�5s�c\z<�ґ"O�aF*_��&�xց���x�"O&$����z��/ч��k"O��3&m�XA��{S�B�zݚ��w"O 1�� �!e�@͐�S�z sC"O� �,�
hD�+�3� �D"O��kp�\$`� ��9ۺX+P"O� ��GB��4�0(�+0T���"O^�N� '=���_R��2G"OV`��cգOF��Ӊ'~9r"O��dKB:1I8��D�Z\^�!�"O�t�� W�/���d��n�*���"O� D��+�T��d�7x:�}k"Oޔ�'���܃Ga�R��p�"O��S i��π/:���"O\( Q�����"����5��"O9�r�?C�z]���A#�Xm�`"O�5��H��$h����@�N��"O�-�r�L�X����즠p�"O�ЛU���7SJ��vI�H9� :�"O�P��� #@�C�GQ=�(Ñ"O��S��Z�\�t�[��ڧ"$�1�R"O��V(�$\ŁA$ �w�܈RW�'31Oj����F3,"F��@�b�@�C�"O��g��Y
2��GڷgEl���"O���e�Յj� �[��	eL(��"OJ�/H�)�L;�I��6hmن�|��)�2O�9��j� UiT���L��v��C�?�Pd��R[vn=��ȑ$Z�B��r�`��#88��D;�,C䉣�X���$Q�m����X�㟴���K�.���#����痻Di�B��q;xy�@��T9�d8�T	p�B�IIfn}`F�]f���6Ð�P�'�a}�"��ǂP����\,� �!;�yI�ȑ�ņ��Q�h4K���y�?�� �T̄��`�1�Ͽ�y"�	
܉�P��c�b��E��y�#V�=.�`��M\"ZRq*b�4�y�4I�$�%��?p�͡čK���#�O:���%U�<j&����ӂ/�����"OBa�c R1��"�r6\!��"O h�c��6�J���˂1~�`B"O L;bg
��iB��@7,�鱆"Oj�s ϔ�w��1�0M�;$r��t"O�P9"aE�n#��
�ˇ
h��*!"Oܽ��/�@�a�+P.n�(h�"OF�Yu��/g����M�_��B2�'��O�U���=J�����W�|P�b�"ON��nP�quL8т��w3��k�"O�ͺV.`E�(p�锩F�#"O�L3#�S�~`�� c$��"O��f@�a�Qu�I�(�^]�$"OЁ(7A��Ac0�;���-_ײ�D"Oz9��,��B$VEc6>s3�2"O|����󰐡���#*2��{"OEP�%K�Y@���Ν�a��}�d"O4q+�.O�J�r�bA�W����"O��@�E��j�矀&�Jݓw"O��*؊4�=�`ҖY��Q��"O�W�!#N�l�c�R}$�m"OR�2`"ؾ-�`c��U�(j�"O������"�jԋW�x���a"O�� $�x�
�X�N,��"O8  �3�����ۨ&�z �"O������5�r����'7v�8C�"O����o�y����M�mN��f"Oi��	�K!��k��*W<�"O*����E�}'�	��ۦ*F�<؄"O�tPgjL1?/zX��DL/1�q;�"O�U `��|�dy��b�<��|�C"O� ���e	�O�@H�tA !v��x�"OR�0�"��*���7.J�y���t"O�XR��֩;z�q�
Zwv�	�"O��T�V�S��8*�*��}�"O��cS�ͧL.6p� ��2.���#"Of<�r�G�'�:)h歘�U�2H�"O~�T �"�P���X��I;'"O�đ#4&r�{��ڏU<4|�"Oz�;�&�E^> �"�
6���"O�Y���E��%Ά: _�$� ��4�y"�Q�����EG�$�g̛��yr����Q�0B��?����V����y2�݆&�
����/�6��e�	�y"�TeN�Q���
���!����4�yҫ�nF��C�õ��x�"�.�y�JխJT�z`��
��a����y⋐�U�v���њX&4�dӖ�y"EΔNSm�r��sD���L��y"(H>L�LhS���&U�y ����yBOh�,,�f'�9Fu��ȓ���y��F�Is��<1ä��'��yBNK�E�>�� T@"��7���y/��a�䨄�C�1;d[6�2�y��^?����b%�%��0�`��<�yRk��C�� !f��G߶`S�A��yB�))-��JEhE&F�"0k��	�y�݋g4Ҕ"ӯ��Am�5���y�J�&����H�?t���DL��y��1��,�dɖ"t!�Ai�w!�d�	%ȕ��ʟI]��iC!�	,�^\pU悭KJ4�d�U�!��mV � �-_&6X�1CkF� !�Ċ6n��09��+H���:*��S!�ԗ:�\�鴀�.l�d"c�W?�!����S�PlR���G &�!�Ă�8wZ��f�H^�=	eG��!��E���xe�q�x9��$�6^�!�D�:'�pa" d@0x��Ⱥ�D_�!�$��kݦ��+��7������{$!��$g� �a��
 �H���0!�$�2&��@O ,4��(^�m4!�F=E�
�����	th��E�'!�ķ$8�BV�E�h�H��A�]�!�;)����
~zH��Cy	!�$Ս]'v�`� xl6t�WM9cJ!�dI23��`� Z^�t+��!��_�x�R�(@D�#0j:Q�!򄛥z�����[�g6�0�A���c!�ĊC��4J`ݿ�%)V�VX��'
&��ԢN1i�͚��<q�'Vy��.��.8x�c�:+d|��'�$$�@ƭq�^,�Q�Ó\�4Hi�'nFid���H�q���)U�V�
�'�b���� ��Rփ��\�E�	�'�,
�`ʺ�<}@��"ƀ-"	�'�l�`cK{.D��{��A!�'O�����-k�6�'Q��G"O�9�$Q�h:l �b-�M@"O@4YΑ\R0���V�,�α2�"O�0�N�`�tB��D�
���"O��8� ʩY��E��^�^�
"O�!�C�6 ��yӠͼU�N�*w"O�y��֘~�r�!��y�J(x�"O�p�aI̮w���)Y�s�����"O� �iD�.z�.mZ䇁%<YtE�T"O��¢'�F�2�+Ǎ�]��u�P"O9�6�F 5��8�P�~���A3"O.y��,� 'Gځ@fbў}l@822"O��� �	�3L(�qt�;2�
x�r"O02���zXRu̗?u�\,k"O�Ց5&ǒf�`mr2+��d�P�"OtuQ��e�҄�j�A`Z`"O*����f@.\E	�n.~x��"O<\Ys�E�
d�����q `��"O:XkP'ń'��\���A�?����R"O6��k�� d�j�7k�d�g"O| x"�c���6�R��Ma�"O" ��Ŏ�j���Q� M�%k "O�]@A�7m�ָPbh��83Q�s"OD�;�:E��8� ����)C"O^�2��Ջ�R��E�ڤ�\�i4"O4�0���&
f��a"T�j����&"O�� ��Ii%��ᇠΒ)D��&"O:	 �g��z��Q���-��J�"ON�W�8?��Yj�����3"Orm;���M��Ai�������GV�<ɲC�";vn1A�a5�������U�<����f1TX�S��
:i�LQ�<�F�b{>E�EL��nn�X��s�<f��	�"�Cf"��$�n႕f�m�<�l��7�����ԁ{m����*�f�<�2�9]��`Q2Fחh���V�C�ɵ)I�ђ̀{��L@ЇݦB��B�ɣYQ�QⅦ�0��T���<�B�3���3�c�1Q�
�؆��U��B�";�t�����(U�ʥ`[�B�	]�X(*vgT��Ҽ"K8�NB�7V�l $LI���H	�o&�0B�	f�[�E��r�8���AB�ɡ!�ظs.Ъ�d؃g�L�%R*C�I�duX�����!WY��:юΆe�C䉍*�Y�[:Q�x��E� ~C�ə"#�M�A�AJ�4"'D�?/��B�ɲx�8�H2**��a�!	�*�~C�0 ���mP�,F a1!k��:1ZC�� \$ԝP��k|P1�"�?~�C�Ɋ�\��fIİ�����M&S?�B�	�7�\�d��(m��ۦ�I
�C��7"����7g��#QmE�/�C䉐W�ra)Qiʢ5=�� �+�.��C�I4Tl,e��)P�:�r z�BA>@̚C�I����D�N� fR��c���nn�B�*�x8p4��� �ӏڃd�B䉧&���K�
����R�X�B�	Yٴ8��R+C��m�F�U�d_|B�I�l��a����>LZ�PC3���XB�Inc�ź��Y 7��Q��P�!F$B�	�j�ȁ�)�����!B�(���D�IT*��F,nfz��/_.0�!�$ůveP�;�#�� �R�˴I��!��[�h��waި:��<�iv!�dF�F:�M�����~i�Eg	�yB!�dχCԜ�7�	�l�`,��3Y!� }�EZ3�L��lY��@(P!����ģ�~��h7�)!�d��l�X����D)~��a�"�G�<iB�Viڔ8���g��m ��D�<���$�I)���(়['bQ}�<� ���E�9ș)�	M8%�h	`b"O�]�
ۥ#��h$�(4�z�8�"O�Xy�
YF�I)ͪ����G"O �a�]�lǺsC���V���"OVX�SKI�X��Uy�Ҹ#z
@T"O��Y�d�+:5
��a$��,[���"O"��@�l�uۡ�<)KEx�"O����Y�kJ �&"X�-F�=��"O@��w�BD�s�+ػ.4���"OR�b��#�M��ʙ�04 ��"O��Xԋ��F�H�� ,��"Oz�`v�*Aܔ B�m��&�x3�"Ol(�S�[��8 io?cتmYc"O��U�+$�1�D ���å"O@H�e/��R��q�=FR� iq"Öɀ ��T�����V'��x7"O�gM+����t�+B{�<V"Oh�Ĭ!Sf���i��av4��"O� �A�����u8�KS�tNQ!�"O�5  ��=H6X f�L!OT�52"O쬰qH��!��y����>@�	��"Op�V�-
B���M��@H��U"O��9q���o�HCR�I-/:�1"O�U`!�X.qg��CG�H� q�"O��S��]�y��I8U��:0Z��"O�d�A��D^��C�&V���@"O�M�7@ԥ����I�)`��"O\)����!��@
�?=�I@"O�-�s�ĂZ�-�`@H�3���{""OD��Q
ˢ3H^�[��A�4�"�S�"O��f�;(:�D��Tqۨ�R"O m���P��1��b��2̰��d"O����^6G��1
�Y)��a��"OZYI'��S��)�#HR4��s"O
�ې��=&h��th[�
�\Ȱ�"Oإ�f�[n�C��HLڕ��"ON���B�"gf��Hq��%L�H`�"O��QfGBz���cfʰ\�2���"O�%��Nުf8�5c�.-��T:�"Or*��*l����TB��4�sB"OF��r�� i(�!+rK��iZ�"O��
�dЯ��(���,kqӀ�y�K�p�����īw	.�h1��y�m8-(��) ,�q��`���'�yR���Z�D��'�7�tA�D�9�y�Ǎ�2�����[O���oQ��y��T�hX�A��D<{�J���Y��y��'�|���+�����@���yblB:0���_$\����s�8�y�K�
�^� �ё)d��h�O%�yRiF<��Ă���O������y�H�(1\���E��Y�`;BI�y�@�fspPkvC�1�� A:�y�˲/l�\
tb��7��ȉ�O��y��SZ"`r��M;6D�@I ��,�y�8m��I1��L/�NI�ā��y��!Ј���*��y�3���y�	*;��U'#ÑQ{z���H��y��4l���cʂ�F�ذ����y���1aO�xP)�8#a��kG��y�
��|��+���	+&��ⓍA��y��]%~���a1�k��A)#ǚ��yb@��AW���d$�=hI�`�����yB��J\�WM@h]���ܷ�y
� 3���?W�\��V1[$�`e"O�p��ňCq*�@�K���,9!"Oޡ�A���2Mh�r��'<Z~�Ґ"O$@x%��P�D�JG��WҴP�"O�����J,%h��y��;Jx��C"O,|R�G!D)�����uF��k"Ob
��?�鋖O�7.���"OX��$��/����čǊ>�l�"O~�A�˦p\LP $��;9
V��"O�����48�:���C�3j{ "O^��bő ����d'&a�"OT�)a��$h]�h ae3h<��e"O��H�j�
�l$�/-uG���G"O���ˈ-P���D2n��1"Or9��db��McRCѐy/�ai�"O|���R�d���������R�"Oj%!&gH�'�,���Ƃ0p�n�q"O��Kń�w��	�Z]Ͱ�"OT�yg��	A�Ѭ��Z���'�Ya��ޠ]�\uf�ƣmK���'|�-�1��1)֜ ����"b�ڰ�	�'+xS3�րk��0�@��Y�XX��'�Č�pjڣ9)����!�P�����'����������Vꅤ;��I�'B�q�ɒc,��� �9��-�	�'��sB*T��aI�,H�V9��'��,5��>\���3��;�E��'��a���+R*>�ZB䜞 ��u�'��\2 �ba�cR�R���Ȏ��yҊ��tf��Hb+�4K(����Q��y��̔r�f #p�E zT��Z�Z��yJ2t���7�^�a���x����y@�o!�B�J��G�����yr��R$�t�>	3:Q
��͒�yb�KV'`ݪ#��	�@3��^:�yR��u:�r4B�ua ��vς<�y�Gʝ>1Zy�IX:��G�(�yb��/Aڜ&�X55~�,�&,8�yr#+>((x��2<L�E[vd��y�%�^�7o�"
ع�'�y�aIa���9A`�( ��1hT���yb��+��y[�E��������ybŊ;U�(#a!C��J���W6�y�=C��=�딋���K�Y�y����b�xL�!׶�*h���ˉ�y��Ǵ$�����ȟ�P��u�\��yrn�";h^ha	���m�F�yb"�G�V�	�-Q
-��Y1�ћ�y2E7I�����#ވm��Ҁ�ğ�ybl�#�F�9ף�
f� b0�ʖ�y��)*�xy(�Q���g���yRlS(Y�j\�u�:5#�m���y�U
5�J�(0��lt �"g��l��4�(�j�
D�7���PAP0:��ȓkd(ʳk�	��I��E�j"��ȓq��Ӡ,�=��	X��[�d*Q��E8�@�ɉ^�����&M�c�,���#��M	���d�<Z��2�y�ȓoV <⢒��-�8Z��L��(�T���o�i�a�
E�`ͅȓQXH��-��
hz��ү�	_�܅�op��X���''��B�׺P[�4�ȓ4X�1��HR%"��
qHF�&>�4�ȓ,�2�HE�O[J�`2@۽r.���S�? Dh�o :`՜�򆇁���+�"O��cr��8y��@+faߓwpz�q�"OHx�S�Zw�
��8A��"OƘh��W-�FaQ4���""OL]�B�]�����QTO P�"OXa���E�^ʪ�Q۬V=�YBAH+D�<X��qь�r.�&��D���*D���to��>SܐHWEψ|���l(D�8�ןz�B���μL����9D�$�3nJ*�,��D#�!H��=x��3D���6%�=h�`r�D��
���2D���%�K�s��-�C���I�����1D��P��>}��1��.���2@/D�H���<���J����P3�4�"�,D�,@�'פ?|dr�l�"v�t���+D�D*���(�eƭ7��/5D���bf���z�g�pf��r�4D�XS�Y�/s�eC��r9�c@L�<1�f)8eB%��ϟ16R�X�J�<Y ��	a�rǭ�4PhXWi |�<��K�_O,��@╚p,z���J\�<AS*��hpII��|���h,P�<���U 9�j�9�kF	R$�����^a�<�K4\��kk�;�X��&�\�<ٳ��.	�l�C�G���d�\�<�0@KG��m�P
v(@����Y�<��O˃:VV�p����o�mc�@q�<Y��B(&�R`��\,郤� G�<��2g�,)���+V�����{�<��śf]p )�ɉ7θI�EON�<Y��U?%XQ
��y���ڀ#c�<�獂2D�vt蕂�icFᒒ��]�<�3g�	o��ij��K�;�" +��a�<���3�Rl0�"֊X�d���HXa�<����8U&<�����9�v�<�w�F*l�"l�I����qՍu�<�w��;1	�%*$'ʺm����4�q�<	�g��1q̝��ȞڈIis�m�<I�X$a�J5�Ц�D�n�F\h�<	�K%1���X� �^�򇎟j�<��P>�9��*D�r���G�}�<�S��vƪ��u捈�,��@�	d�<#l�zZ1r�G�Ln��%&�Y�<��hU�:�J�a"�#	���rD&U�<�cd��"�@(3�Ѡ�!�O�<W�76t�a��G�[�t�A�(�M�<%�] mič�k 6G�m�Gd�N�<Q�'����֮n��QY�]J�<Q��˭H1�a���L�zn��c��\I�<i��ܝ����mˋx��h��I�<��ϧMO�S6C��ѕE�C�<�cȑ!A. °�ߕ\�r\Q�|�<���F	gJ��=��Q��u�<y%�Ϝp�8�B�O���(�{�w�<ɦ�ܨ�h%鄦[?��H�u��s�<�;O�ls��E�`��	C��J�<��L��H�Ʃ��CFRt��JCF�<���N�d����n��Bz�����EA�<g(^�8آ斔'{��:�]~�<���f�� �ā��o1���[o�<�"�P!R�{"K	ko*��tf�i�<	��2�-�`#�`(��7�z�<a
�َ�AĎ#;?J�IcJ�O�<!6�&-�,mA�máK���H��IE�<� �%��O�:�1񦆵(.�ِ�"O8�� ����<��F�v��"O������VQ�;�c] iH5��"O�L�'`��}�p�BM�t�����"O��Bcˁ ��;���y�~��4"O�S���C|d�"�΀YҀ�ZU"OQ:5m������(F$8�.=� "O"T(r&���ѣB��8{&X��u"O��U ��V���� ! �7"O�-Ka(%f����*{\��"O���-�o��eVȟS���y�"O��b瘲z��Eђ'F=k��C!"O� �%$K�,8�6�ѷ@K��I"O̚A�C�!�x䲇���b;t��"Oҭ���	U��8�ɓ% 2(9�"O~Q��	 +.��Ka�Ŭ@�z�j"O���t�&���Ś�>��s�"O� 3���am���p�ų/�����"O�蓕��hHP9�"L� ��x�V"Ob@:&hW�D�P%;��&"ȅ�d"O��R���&+�(H�cǈ!W24*"Odu�0�|�R(h�� j�d��"O&� c�bh��wjҾSO�݁�"OɁ���anJ������Lĵ�D"O�c@I��.�8�KS�O�B�̓�"O4M�b-�4w �`NP)^Ґ�"O���å
(MM��!"���`�>�*�"OL�[q�Z�r|��6&^�>���"O�$�˓;�uZ��^�hE"O��СL,P� т���L��IS"O�JB�>;t���$� 9�@�)�"O>��G��2lo��¢�S�$[Ƞ�"ORtz�-�>�6��e�T�~1�(��"O伓��1�IbT*�h9=�"O���?[ 0���& ���"O �����Z��A膉h֮�!�"O>Y�a֌t�\�
�`�0a����1"OiX�OC�]!lq���/�B=8B"Ot�;Q���Tp�5�`� �np��&"O~��F�׮@h`�{��X�Zj��I"O�!�oO3Y���Öǜ�pKx�0"O�ik1���RxY���yA�E�"O�S��G55�d��Һ=.QS�"O����6#+N���+:�j���"O`��qÙ�q�q�w��<�p�r"O��m_35��% 7��sX&��"OR�U険2~���΁uK�<�"O:� ��"
�Tl
?�}��"O�]�1N0O0�1����G,�=*"Oș���˽.�T�2��+ %hB"O �`���O��je��W���"O~)�㭇V���o�*W ���"O�ۃc^�!�M	����*�(�"O~$��(�8dwt� �LQ;�F�h@"O�M0���@D:T��%� "Oƥb�!^�B�+� \jd!C"OD1��癫Z�r��fh�(hT.���"O�m�C � z�PUe�(E;6,+�"O���2a�:^���DD�� �޴�"O�D�N��L�������.�3 �	O�<I���n�͢��	Hľ52�v�<�����&�B��5v����@�t�<%bˌ�P�u���X���&�t�<���X�09VŚ=d�x�v�q�<� � �F�J��h41@ч�vpa�"O�X�ҏ$ ��<�v��9:$$Kr"O���U!A")��d���v�0"�"O���D�6�ʝ���\,i$�p�"O��	�)F !�h�3�b�Z�("O����
�J�6�r����jA��"O��A�?4v��	Mjl1"O�t��(��p�n�A2t��"O���Cj�
|��C.M�w�8��T"O�A���!���3mҟ{�����"O$=��O�ltyc .^jԨe"O^��*_kJ��k��L&R�f�Y�"O�h���V/Z~8��:N���Y6"O���P
AY1�p�H"e���"O�	���%�pC#�I�[���"O�8#��'cԴ�%&�4X�����"O9�g�u���b���8�M
�"O���&�R,8eR�`�͂'���4"OX����:%�a) �37��1g"OfI�ݩۘ� ǋ�О(�"O�;v
#(�������qh���"OʕJFg�6h��c�E�]k M� "O�k��q(Z�2áY$Ce&�4"O�kB��9e�DKv���pGd�"�"O�\j�-�"IH�� �oA(A>���"O�Ep���������Uǖ�J�"O���+�#t��k�h�
Ʈ���"O��9�޽h˲2'\2La:ȘU"O�D"6.�=�\m1��*YP�D"O1�t
%^K� �&�sJ,x(�"O~�PC,�<X�� �qE�7}�k3"O<ự�@�P��E�%�q��"O )��H�E��ץT��̢Q"Otb1'F?qkY���'�Y`R"O��;���a"T� �DM�#l2�S��y�g��6s�@c����x�a�����yBϝ,F�)�u�O(�(�ǈ��y"���v@)�&l�4	6BPA�N���y��*v:����ˋ˘��A�_��y�	� ��R�!����э���yBD����Y*q��x����E��y��C o��ÇNO�$�xt�����y��U�F�H��E�U(�,t1�E �y�`Y�Y� �kE��G�Q��Ե�yBŞ@]"�b��)Z��0Sf�N��y���N�ٖ鎦Vِq�T��ybB�*� ��C�Y�!�֍;Q�֨�y"
�va���S�,ה�����y� Ҁ�P���Vl� h� �y�%=l�rcɅ.9�����yª@y�ȉb֠~-.���۩�y�	�?�ltAD��~ �F+Ж�y�`ޮ%a4]K�ÅFg��"���yo�{n��@!,>���D+��y�.�&9�xqP£�64��	7���'��e���	"��# �l=R8ö"O �KP�J5cP����?(F�x�"O��c�(6"��$��9�"O�]06.�t�0�2R�F]�`٢"O�U� I��8�V�bp�T0�E�"Opɑ�]8G��ᆊ�N��0(w"OR [6H$�V+���V�K"O��{`J�'!�B�E�֜?�u�"O�����S.��f��D�0"O� �d����1g�d�G�%�V�j'"O�MJ�Ɏk�`��<t�|��Q"O> ��I%C��ȘWV׶���"O�s��k��:5��=,F���"O*� �@�p�����+�>h HT��"O2��w�,w�~��U*�b�J�JS"Ob���͆�V�V�2��OjG@d��"O]J��$Gcf�S�)P�b���B"OTmkS����b�X+ǶK4�u�"O ��6��`�𸨅��RĮ勆"O,�B% �J-Z�	�E3Q����"O�A��K.{�j5��J�?h��`"O��Q�>�����R�^�%��"OЂ�
O�VS�<�gA:E,2�"O��KQ*��ew�����^� !"O�(���C-�F�@$���p1d"Od �"�Ur�)ᵯ�b{00�"O, 4�yX6����]_���""O������T��MB�,WB)��"O�iC fݑm� |C���6����"O�� �儠���E��&Ҿ�)�"O�萃��lzmS`,*(�u�"Ou��2��&�C�J�!�"O���A%ߞ��W+�"�`�"OLPb$5`d��AGIq��pu"OZ ��M�����(ܱ@�<�#$"O�8K�E�M6��A���"��"O��*���j$D��R:S�`��6"Ou� B����b&�+:��K6"OJ}��Á�&LT�ӣ1�yZ"O$����3�L�S�G|��"O&���&��99��AD� 1����$"O�#c�\1$�d�T�ȳ:�x��"O���u�
+�`!�r�Y=V��ݩu"O�I8��׬U�|\�E+�9��Ѱ"Oyz���"�vHj�$C�8����"O���PNPX��֢��l��e�P"O�	P�A�8�HD��!@�2�2ݐ�"O(īaD_GHy��5B]���"O��i� �fh��h��E�v�|R�"O��"ӬX'}�a�ͰW�1q"O6��Q�ԩٺ��!J�==HY1"O����@�$k`�����+:-И��"Oh��ԣ̙fL͹��>9��J�"O�ݩ��$;�\��bQ��@{"O��re P-.s�Y�# V<���'"O�)x���	��5K��T	^+��W"O�xc�m� ;�rHQ����	����"O�Qbp͎/s<�p�L��q!��A"O��2�D
Y��4�삫% ��"O�Б��_9\t|�R)|E�S"O,��䚨2�<K�P��#"O�@B��:��%�)0�jyQ"OT8y�03�����-��dҝ[$!�$��JF$�gI�0Br�I�Aʝ�1!�9my��Т̙D��h`��`�!��
�Yj��@�B�M�����c	T�!��V*$��"�a��앉աP#/�!�d	�Y��qR#&�/�
���Ʈ!�!�dX�!�"a�c-ز]�|Q�ᐌH!�$AR��KEm�	or�8b%N�G#!��74��� %�l��z��B�,!�����~XW.DΔ(&�L�c�!�d�0�f\!Ǐ�̜�4��*k�!�� �`0%�bH`�[w��#]��DK�"O���:2Έ%�%Ah�LlI "O����t|���%I�gqf���"O�Z0��$k����IN�J_��:�"O�J�悽Q�I�PI�,Q2(�"O���ר̳f�T�3�gB��Ĩ�"Of�%/E�/05cVGʢw٪ [v"O�P��ޒVxma��^�L�:�P`"O�%�b�J�F� ��@
I�"X�7"O頶�Q�3y���]DjT��"O��#'N�*�;RM_�|_�"O��; �0fv�x@��2v�	e"OlIvb�	0|���#k]4��Ȁ�"O���؂0r�<:�)Yjr��@�"O���'��r���a��Z�R�*��c"O�u-v=����A��r�|l D�l�'+30��!�a�?�X��`-D��BF��͐(���لz����
-D���4��Ao ��˄2	�����*D��8�E�7�Ѷ���[���.D�P8�,E�)>J��!�������)D�0"� U���!!ײ�R�1�$D����Kشbl��،(}Bu�!�'D�DAfG%
�2ɓ��T�s��*1�8D�\�Ԇ�24�vefL�by y��/6D�T��m�I?<p�'wļ0��'D�ز��K1<��bDɄ9F������)D�2ӨII�콨 b�SP�3Qf(D�p0T)̮:�0�ӣT�z���sS�9D��C��k%n�b�E�̬�RD8D���Ň�@}��E�L=0f�5D�|R�B���� 
�Fz���9��8D���S�x�ybqˇ�ܫ��*D�p�ߚR��$�P�0"�ђ/;D�8"�ȍ'}F-��� �ZE���+D�8��K�Z� ��A�K�hi
���.D���T�IV ��F��n�����a:D��⤬�� ��J�z�x�,D�A��9�%�Pm�)>6���*D���臝l�j�EՖk�||���'D�X���?dl���&'�	7�H���0D��P2F�*;D,U(u�*@p)a��+D��A-�$8��uD9E
J��(D�����6�$���BP�ŸP%'D�(�E�	7(`���T41�<`��%D��B ���&��0�dΔ68Y�����.D���lNJ�$� �r�,��B䉣@�#$��y>�m�f�D�7�B�I���X�J�
�¥��/D���C�I;C�\�@������k���)ԢB䉵^tR�*]�N������:_%�C�I�|�m��K��S�z�)�
�<��C�	�T��b��ɚf�p�b7��C�I"K�b��`��
`����:lrfC�ɀ�q�C�I�F1bL(�@Ņ"�4C�	�{�4����N"	����t�Ȝ3M,C��.+�)�Az�������i�
C�I�<C��Eh��h�IE��c��B䉆E�8`8��&�B9�+�O/�B�ɝ0S\XY�L���ض��hغB��,h4�6�T�ll����j�B�	28�5���'è�ȡe^&DB�ɷ�E;��W&��\+B�ۭ5��B�s4(݋s����5�F)�IG�B�)� A��
k�@x[`�+>"���W"O�4:�c�.*VN�;������TU�<����By��R���&4jȣw�
M�<�e��7��=	P��"伫���C��h�� 8�S=M%���,4U��C�#'�:���#��_jl��D�%��C�ɪH-�4�g����`�"eLD�} B�ɍIRX=��G${:6��v�]�e;�C��?@c`&�4?�}��\�nݶC�}��!��{����隂4�C�7��2ҋ�)��1B iXq2�C�I�{*�����
 �]K���g�C�	3#	�P��ÊG�|�97��rC䉠b������v���kZ�7KDC�ɞyB|���փK�H���%"�C�	8e��0E�ьb�Q:���fi�B䉨.�؀� ^�-�"mYW,I�:h�C�	$�e��!d��Q�cBC��+���᢯4UM�8(�&&J��B��#[ц4�B	�d b+ /YB�I�H����UNI�e5���'��ED�C�3v����%�wN���D�[�*D�C�	ђ"c�4X`.�#� ,�B��Q"O��f�ӛ3N�xQ 9��\J`"O,0Wo�iSLt�֮� O���"O�b�W�-���߯1,H2"O���i�	�^�0t$U�2*�"O@�h�E�Kwx;��9\(i'"O���Dč�:{(���58P��ZD*Oj�"b��%g���(R�!"���'1�9kg��(R{�@��#���]��'�$�p�dA�hV��b��ѱ}�d��'�699��� ����6$	�p8�'.��:�� ����F�V�.?�m�'|桰4bɫIt�� C��3��)��'�q&FH�W<�j"�6����'�p@i�"h|P<p!�M�<�8
�'�.�"�˚�r;La����~�B�c
�'���L�+m��m�R��EI��	�'� ��ɘ�? �Pq�5?U�̀�'�j�16R�$$�@CV�2 I�
�'�ʙ���¬���e.N�����	�'D
\�p�P#�e��R ��'��-B2�̲��BU �%��s�'������N��T�7'�d�D�[�'��3��6ͦ�(`�(�ī�'=�s?1D0!�Q�Q2���'1 m��H2�T��0�
=	a8�s�'�|Ah�,\ȶ�aWa��o>J�
�'��$[�C�bjҌ��Θ<7:&P��'	xcߪY�X#���@�P$��'b�I��$o���j�6��C�'Ȩx��	�,��HQ!P�A�� :�'�<e����$b(�;�[�Sd�Z
�'~�uBa�������K=/@ڑ�,D�$����_26jQ'� ��=D�8ꏏ6�6'�;bz��Q�<D�P	�lE�-=�J���}]B��bF7D��h���@Q��]P��9�9D��V	R*>b���u�E�x����8D�hhb6$���B�L���.#D�hY3�J0N�(�!�� ^�	C�j,D��� C9Lfuc�d� A�A�`�+D��{�$Q:,��RՈXv��C)D�� n=z�%�[Լ�v��0�<$�"O�%3�L2?,P (�[��P�"O�tcwn��L�3���	"�^X�%"O�U�����O*�qS�/ �FA�4�"O�AS�ا0k$�����M ����"OX�E�YP�HM�e�R͐1"O��Q4�$ne�&ȏ
#y:T�"Of�Z��7��� �8cd9Ju"O�m�!���D� �r�	/Z� �"Oʡy����A±�d�����m�<����dk���nTA5�h���
i�<	D�R�Y��)ƀ�+wlDp�'�z�<� A7H����l#V�)dkw�<i�O]�U~�S�n"=#X��"�q�<��� ���]���q�q�<����MI�I�r���rw@	p�o�<QBD[�S. # @�h��[$+�m�<a�L�Wʤ�:�+Κ��Yc��E�<	� Md^&�˥疔@y��F�B�<Y�ʈ,u�\ (�	�*H�Z�C��y�<�C-�)9T�D��0y#�E�g�r�<�� (G�� J"c���m�!�H�<����?Zb��"ߨ\�Z�$ �<��إa�hH�ڦqx��z�.s�<�#�T�qu�%A�=O+��!��h�<q5ō:L���0�D01��V�Bo�<yB%] _�0��[o�(�8�� V�<ї��*��x��mp�pq��T�<9�b���@0!��>8ZHQs
)D�����~��MS�+`BP(�n4D�t�֪��Q��4ʀeV%X��D-2D�`�!�W�c9f�I���%�H��l2D��;NV�I�`��	V�>�m�r�.D� ���ʌI5\�"�Ƣr��e���1D��xeOB�1���P De����A.D���ј����� �/h�ai1`0D�ܲ� J�f��j����"�3D����01���$ϊ�X���(@A7D� pt'ČF�8}�g�(`���{�2D����nA�J�K<"����t�.D��H��6k����q�w�q�	.D��b$aX$S$1;�_/��mk�j,D��Z�F["��R0WLt��)&D�x�7�P2��M�!a��Ei�&D���3oE�o�����ĭ��ՠP #D�,�����4��MĖI�<�Ug?D��B3GS�U����g�c+�s%#D��X� ����u�O�3%���&D�\ht�@6`���5��a���)8D��Z!&�=un�j !WpÐl���7D��H��<��؉gV t~,�$7D��A�U�քy3�I�K�h�f�0D�ܡ�M��t�ҭsW!�1tZ���l/D�xA.�:pA��B�w�x�Re#,D��a�&E�-��"S+=���� +D�@�7J�#bp9��ÕUX�	P�<D���&	#]��$��ʀe�
P��.D�@��
Ǫ,Y&��� ���+D���gȏ�	���F�F��;$�(D�\��KW�JJ�,8b�C������(D��s�D�om��j�3w���h��:D���u�ΐ:w�ˤ�P4���TL3D��B5��-{�e+tI�u{a�2D�H���B�G6��K�;�f����1D�� �tHP#6f�,̢&��r�[U"OV��F��� q�2c֢j��9�"O6ʠ�+�
�X��S�*_dT��"Or@v�حP��)���]"Aب�1"OR)[E�	�b��u��
 "����"O�E�@"�ophq�n�124(�"O��%P[w�L뵬ƋJ�5"O�d�A/X�4��&��$X��%�"O�U�℆�a^<���̆A���ѕ"O�xе�_qLMȃB��w�l��"O`����v��ej� 2�԰g"ON����Ww��$1Vi�'m̠�D"O8��u��Mx:��	�gM44QE"O��q'B
vAdx���c���"O���uǂBc��hڷ):��"O~\�&%� #lf[$E��e�(�0�"OTM��F��̠c0BP9��(A�"OEs��Y.�����ʈ��Q"Ou#�Oʪ!��m��1���"ON�����?+�Ҵ�b�.+��{p"OJj'���i�����>%�`�H�"O�(�%�B�m�ŭI�s_<}��"O��F��4���@u"ԻW�b�d"Oč�H���Ⴠ�0?.-ˇ"O,���kY�s�Θ��iaR��;l�!�϶f�5�Bg��hS���!�QUS4Qї⍔;Ȉ-�A5E�!��xR,�a�֨e�:|�vOFi�!���2Gz�A4aG���hBf%�U�!�d�~�E�Ι�^��u	f����!�[
��"2Mˬ%x����@�!�J&P����� ���X��B��	�B䉱c-M��նE���*uD��	�"C�I�s�x�3� �qt�@��H�	�C�I�{_�]˅����@zR
W/��B�RWt����.y���X�gSVe C�ɧX:�}�9^�P�H�/��B䉅l;>�4eQ	s�d��t��B�!�R��p$V
��21F��z�pB�Ɋ(�r0pG��+|"����g]�!�B�	.FXc�L�"J��X�R$ؘp;�C�	�jt�Ąc������,�2C䉂a5"9����N�p�
 �DC䉝v��3P��%�$��0k C�Ɋt:�����5���G�N�'��B䉜Ɗ|X�#��"�rm���%_`�B�I}f�XGbP�U���b�ο$��B�	�I����L	т����	B�B䉳Ch�8��	[�l$Jp8�J��mk�C�>�<C"�V9F� ���η�C�O����!��i�9� BLq��C�ɀ7>��)ɿNtdK�B��S2C䉻R.�V,A�-�Ht��	`��C�I+g�%;��.ov<�aL�Gq�C�
��Ay�A�aEB{ō�yA�C�I3].ʀ��۲l,x��M�c��C��|ΰ��Sޑ8���4ƚA�&C�(|����C
9T���6HUI(C�SDp�B�#��:��F5�C�ɯ,�Ԙ�#�˂u	wg¥b�>C��5��,�/�33`m��R�A C�ɽ/�f�`�K�"�f@{w�[''�C�	��ٖh�k� ���ڑ��B�I�tBA��MA"a"b��>�C�)� �aUd_�{�%sSf�3d���w"O���So�H�a!Tğn?�\��"O��S���TE�$��7#�٤"O򴉤�C�$�F��!�]�!"HԀ"O� 4�ՏaHz!���		$4 *O�ț�bSv������D(֜��'��$BN�u�l��P�ܢ�Lc�'�P�I���~���y��<y����'��$���ژw-�]S ���z�����'4�+�	�*.�he�'��t�gr�<I��#��`���W�s̗�^LC�#*ݹ4�@Lp�	B�Z�[��C䉋�Zm���'$�	[W�C�	�0,� ��	���Qe��J,B�Ie�xE��8%�^8)!
_���C�	 =BD�XElģV�8��[�8E�B�	�
�P�z �4Fځb�#\?"B�I�@�܊�f��6�©sä�T��C�ɩp*�0�a��&��T8�h�;բB�I*�Ω�s	�w!�	፛.M�XC�I�
���ÛL!Ġ��JV3\S�C��Z�R��&�1%�(3e咻
��C�I6_���B��8�$���BNB��@�BT����1.$���-OUw<B䉊ux�`����U�>E#�3I�8B��=[�zXQ�O��{��a+N�'�C�	�j�Ƽ��� U�DĬˋ0��C䉻U.��5 �K�B]�2�,H�B�	�y�!�ں8�D�&�$��B�I�w�du"�ZS���GD�4`2�B�ɺ#+|9o��!�\���V#
�~B�	�-A�M�+V�n�ܳģ@!&qTB�I�I}���`V��İ �C�lC�I�Y�~�2�U�E�r�QG-<`<C�	��X��U���@���K9L�2C�b�6h���
_�+�@=]Q(C��(\G(�B`�=0_P�Q�\J��B�I9X��=�L�<'�������)Z܆B�=l `6H��}25F߿E,:B�	�!����n,|�n�S�0�"B�	J�Ԭ�2K�Z�2Т��aP&C�	1k���ˀ�^��h��3�C�I�>����,K*NY��Q�$�xC�I�@�u2��?|I�ʍ�c�vC� }�� ��ʬh�00���7 B�	 �D�q(Ԉ^��H .,6�&B䉔(�R�wŋu�ͱ�Â�O�DB�ɿ>�� ��9!�H5Q��@�fC��?����A{
�z��55,C�	�0T���BR7ڀCfΠR�C�I�__`5zgB4=%��Z���K��B�	�C��ɤ%	�p��,9刕*4��C䉙�浣�^�i7Դ`%�Q�4Z�C䉾��	k��Q�U���%%Q&f�C�	�"�L��b�v����7���d��C�	'8�-���U�=|����3\�zC䉡6��ӑ��*�Z�@�eʐ�pC�	+]r�mco�9mFX��S)�\�6C䉮V��J��Z�6�"H�!ix6C�"(n�qf(�"��9fC�	�al���ae:�4á��%��C�ɚ(�}�J�{@zT���� f�C�	�xH�;7G@�nN���`�aj�C�I�Yj~Ip��'�S/i�C�)� �E�A�X'50��AG�G���;1"Od0&
��H��5ɉ���"O�@8���#���8@hٻ'- T��"O�E��*pTH��g��h��i"OL�F�U�e�5 �D�?\zg"O��MP�m#0%�֓,��Pt"ON�:�iѻW ��Â�,�Z�z7"O�!ZG�X���CN�.���"O�)��	/�)��ʙ����X�"OHP��M�r��	�1����\	G"O2�:B��%Mt�"%���b}��"O.ْ1�E�m�&�-ur�<�!��0�y���C�%�4��?� ���К�y�CC:X�PA����7d��#q��yA�0����fFI�-"H�SA>�yn2�@�"���F�l	��^��y���4cW҉X �#��"A�y倵\�Ɛ��8����R�D��yr��E� �V+}l���1GV��y2"0)�aJo{��������yr�͸y���Ӵ��*	���N��ybb�s?�[ �
1&�0���/�y����/q!sV�3wxx{wD��yr�ѦfS`]�
�YF�ʦFO��y�����ر%�!W.��֠���yb��3�~A"CK�}#�B֢ �y2D��0Al�1�B�:�mU��7�yr	I���1�SDI7zƬr��J��y"��"h�!�{����"Q��y��01�&��TF$J3"�q���y�+��_�
��߰+�Q��!W!�d�3:�`g���H��.�5b�!�d:o ��C9N����ս�z�"O��Y2�������S.ָw�� ��$�6�(O��	�-ڵ�ܠF~8�5��0?�T���<��w�Av�]��-�X�`�" �)���!�,;t�ђ�H���u�-O�#=4I��V��Yp�lψ����G�b�<I׭��H�0�X�,R�
��9r�^�$-�	S?A��T��*s+���
2::����y��'�t* 盌
�f9�7�����M>�2�#ړ�ē`�� �bZ$^��%� &�z����ȓ֍h����}�^`�!�riZD�ȓ&$����)�r:��A�;*Lمȓ)��gj�qH-���++F���ʓ}{8ᗮ��CL��c�IT�0ޞB��m��"\�]S��zg��&h�B�8i���x��ۛ:�,-��L�4w��B�	�P�|=�p���� ����B�S�*B�	�? ���D�K�=��b'��v�0��p?�e�w���h�`y9�C�~X�H�O�����D� ����'b��:/�8�"O� bT
��W��,���S,$`)zcOܔ�B
�,]��آ��D�Dx�u��x�<�S�4!�L�� �	e�� �
Z�<V�( �$�� ��Q�j2�W�<Q�$�F=4i�J
!@���)N�I�<i ��	5 �����6�x\C��^؞P�=c>!-Q7���"�,D���S�<���R�S���ӵ�]�8ZL���O̓�hO1�,��Ư
��b]�P"`����"O�q�Eiح*I|رU �/����"O�,�m,+{�Xj��L�
��TI�"O~�@ĉ^�aB����ׄD�d3�"O� 
ѩ�e�xü�YK�5CV�'j�F�|2�@?B�5i�'jy�{��y���]������k|�K`iD��'�ў��II���T�9`�"�*`�.	�B"O��&b^9w���)H��V�I�?�����4-���8)�(;#N�.g�0\��"O��I0ˁ�z+�t�c�Fw�K��y���B��t�LI/b�N�C�H�yrm�axRUS���qv(M#���y�Q�U�Z�:��F�V@�R��F�y�t�� �e�B�M��U 
��y��k�Ji@��vz�}qDR;�y�Fʸ_�m�s��	n8�W���y�L�l*<1�U-�U��
�y����C�9PM`�Beb#�y�L2����pJΩ�q������y����#e���T��h���ꦤ:�p<�O��"EN	�&�X7A�� �L�b�J ��'�(�Á���r?d����>Z�(���)?9��iԂ#�^2�B@�%lЪ�
�9`!�dG	\�BD�p��,1Vl��IK�o!!�1f�x4�@�ѵqs@��ś�v!�Dˋǐ���w`p4�E�H(!��{��	⮈@�ڊX�!���!������<�eDE�v�!�dP!0~тGN\�3�"����n�!�DI�E�� �ݻ�dx��D�)�!��b~���K�5ƚ�Yv�H=$��ٰ>�P ��N���"cn[�`V���r�<��d �2���r���rvԫÍl}�'C��j�lñtK�<	�l)z5nyZ���$��a����
{��q�J?4�!�ӧ�6��d�n�<��BA�I!򤂾X
��*B��o�!�߅,!�$��W'��W���Ud(件E�;9�d-�O���K��d�<z3H!�BI���'��'����@�)�_�( �'.rDcuM�:2���3-������'1��C��i[X���mB�*�'����N	`X� ��Lg��H��'��y��T>u�|Γ'1z��ʝ�(�:T��:,u��o� �#�3"�΁�DHE+S� ��ȓr#%��N�����FmW�}�VՇƓuS(���ݒJ����㏰s,a��'na"
M/K�D�� �
�@%��p=�}Z��=�����5�a�*�y��P��^;4o\*{m x*"�Ҹ'���>!�	ɰoi�lJ��`�F�V(.�!�Čs�<�K�fe�r���'�!��ub`���s��$Kv��$!�D�2�~��ތt� ��,#qO�x��'�0E�4�E� �p�F�M�B1I�'��e�"o@T�{r��&�
�j�<�F�'�\˗I� �  b��J��G{���&zLa�̛,+$�X�����y�㛀(L�,���υoƚK��A��y�H�GK���cl�?i�6d�K�y"�6U��3�/B�^�Ti ၩ�y2卩>TE�V%H`?��X@ʋ��Px²i���`�F#?s���u`ܾ%��L	�'�qS�,OB8lӇ�˂S�B��Ǔgp#<Q�&��R/E�M�0�g�T�0��dw�h� �����e�uŔC�Vy�b�T��Fx��9O��[�b�+�:�[W��$K����'�"=� ��qE�]�i����H��(;~��w:O�	p8�PJUEZ3�X���"Rg$,e���?}��/��'~f�r�&�?pH	5I�6a��'���a�.qb�����&�4i�'�X<�	���8�ueL(ZTh�'׆�Fm�<J��%.��rFr�)�'�� �\�\:��c�#`��y�'��|���Օ��@�� |�f9�'���
�j����%N�lL�@
�'�0�i%�B2xq@�yt���\��y	�'�$S��PG?���S�D��,I	�'$*��f��;_�,\
���0ՀT	�'�T���Ɠm��,SQ����*9	
�'���A��f<VQ��Z3�ȣ	�'q�T W-P>^x�r�@ǓSgpa	�'���g��(N�n��ѼЙ4&�yc��I��qpR�� �x����y�����9ё*À�0T�Ԧ�y�C��)J�hڳcת6Ʊ� ˋ�y�MY2oD��h�#_�0��m��Y��y�N�*-r]Z�F+������y��BA�=��΍�' ������y2dB�Y���r��°)�}{c�K�y��޿N�:�I"E�v�P����.�yR�D �*(����_J���jF��y"��W�Z�B�@�I;J�c�@O��y2b��b�	yF�CF ��!�7�y�`U��
��L�t9�_�y�h�h�pB7cT�>���C�k���y"f�r�>���	�:sԩ��a޺�yR�T h�r1Δ..���j�g�)�y��I1���X@�$�t]"`(�yB�91��YR���@@�O��y���\��!k�JW�uhX\0��ѧ�yR�X���8P)-��	A��y�L<O�`R�ꊺe�,�P�J��yRA��j
~m�ꂚJe�!n]��y��]�Q��A��#߿ �lIbqD�yR͞j����gEC&��Y��k/�y"*X�$�ݚ�l�4w�d�2�n��y"��9}���Z=��(h%�y�إذ�����;+�Tx��^;�y2'\�4eb�HYBB6�ꗨ��y�,m!"�^A��Y�WÅ7�ybA-^xE�ש�6d~}�V%��y�l�=.x�cScZB"�)�F�'�y�׀xM֜�)>��9�c+���y��ʰ]���r�ʇ6AYX�js
�yr�(z�:�8Q��9N��kb�*�yb%�'Ȧ���8}Z� ԙ�y��#m�r�C�R�M�U;�����y
*9d�Z$��?t���ع�y�'T�DZE�ޔ2_�Բ��-�y��=��Б�d	',�MYR ���ybj��M��퐣��'�V�Ju.��y�$��;���N�R�z�.���y�
_�:R�LI���"h�L�%���y�M�L�b  �_9b��1*#���y��ӗZŜh���a|<� ԥ�y��ҟ��Tb��W5Jv&����̸�y��Z�X�xRs�I�F�v�!�\��yrj�����cN�P�nm��BN��y�Um�0�p�U5K�)x�*��y�*	�2a���elE�D���CDgۘ�y
� ��3V͔� ����'4o�T v"Ol�J ��,�r��Gf��J���g"O���呜A$��C$��3s����"OԂW�� �[ /���Y�"O��i��L,u���[�Ǉ�l��eQ�"Oy�H_�0G�����٠5�P�"OVa�4���8���p7�=��Z�"O �RA.]�2�xh�R�;�\̉�"On@&_6\�d���o�t�$U�p"O<x�6F��Y��I�����$"O��bu	�/�%1�n'�zA� "OV�"��ݚ,�6r��Y�e�J�"O0p#��ǩ�� "�m7���q"O\ IB�H�& �`E ��(t"O�Uc�-�.% �\�A��g �C1"O�]ѧ�f�F�����q
���"Oxx�a�|(P��OD'{�P���"O����AK&0�v�ؓ�\���ݸ6"O�#+�����-B���;U�!��?=R�i�nM�F�@��Ñ�/(!�	O��`ӏJ���3��hE!�D�&P�x�{���	 ܔ`�uA�!�Dg�R����U9j�2��qf	�@�!�_���)�td�<<D406%�3-!��Y,�+��!x2���?�L�ȓ7�`�p #��J�'%H�F���1�� �e�H�Yk�i�=t��Io�'<���!��%$}E�ár"np1�'�{�I��sD��B��ȑd����'kZ8bU�ޭ��P2���`X��'.t�B'_:e����d�
{8h�'�9�`)�#bH���ȥw��A���~"m^���F����h����y��Pk~h+F,�����$

بO�#Z!J${�h�����T�~p�T�U@�<i��0oK�1)��ڨ�m�5�r?!���jdQdE�r\ҡ	R�L�g�B�I3����Bˮ��w�8c���'�J�If�����U�P�H7B�b�IV��>Ba��O�TY�Ç�G�d�$kK%p>(�ڦ"O:�ꊩ`�}
��^OLɡ�s���)J�X�pm�w�ȓe��+c�7$�l�<�	�VR(�I/#��qP�� v^���E?Y�{��I�R����%I#���R�y��B�	#��T%F�#v�=v��/�NB�	��Z��IeT���L1x�bB≨��X��#�U�����H�Sd����'E����7����Z�O^, �'@V��
Z�E븄�*I��0���'�)��N0�+�雵 ې�[�':5K��4 I(�*pL��k�.��'Zx��`�3|^$�WnՒe��ջ�'�N}��W:$r� ��J!g�ʬP�'�������<���E��L �QI�'j�P��Iڎs�u��E�=�!�
�'6�y1 ߬`T$�a�"=����'�&qx펨B����0��
k�ju�'	���#'�7�����Vk���
�'A�PBu�@�J���Ȉ[HV�A�'~�%sn��X6H͏QB������$�o� X�E�Ŭv��xǋ�A�!��2!�Ē�(T�uY��z��!�!�D��]q��R�IV.8P�Q��!�$ٻ}E&��S��kxE�t&��/�!�� �qX�ɓ�Eަ���.�Z�C�"Ol]��b\�%TTh�g�b�@���"O4�aE��1�[���8T/y{�"O��A���,zk�%Ief[,4z�Ir"Ot�����=Z��������J�"O���w	�	8��!#��Ҵ>�2Lu"O���Q��7]�Ub�*�sY�8���'��T���b��9����%�.&����t�|ӑF"b8y���"B����;岝+�ƧA������$�ȓ& D�6*XKA���B.A@������a0Nΰ��ٲ�K�J�X�ȓ1�����!�W�"�q���%>0��ȓ ����	%����ÉJ�~�l��b���A�A9��X@
�C?y��
[LЙq�вb����%��,l���m�����@�,F����Cs�6,�ȓ�¸C$��nU1K�#�*u�ȓE�:��W�!LBd	����"�ȓ7bP� ��I�0���H�����C��ia%'M���sC�!����|�N(�B�O0����HV�9l��ȓ*uz�$��7J�2�QD�گz�,�ȓ(y)��;d
�����j �Q�ȓR5:琿Q3䰃���*!�I��9%�U��F��ZJ�ŀ��]65�6�ȓM bY��^�a����LU�?*u�'n�}b��:vR�`�mE�h�(�i�3�y/�v����� Ě��gaH�y�� ��
�lւJ�Bq#��M��y򥀒T���a�BC`D:&�M��yR.��JP{`�	?8�$pq4���y�c�0Z������(�B���b(�y"�@I���ztk����ʐ(���yR���� F�� �
	�p"N��yR� ����Ӥ�fh��-��y�f5q�9� �O֚�0�>�y�C� �xp&�?
��/{������T����-i9R��H���ȓJ� �h˒�AӰ]�I�����_��,��g�|���`�ł8Fi�ȓ/��:� �+I��KAOז:�u�?!���~jV	T;��Qe��'?z8E1�UQ�<Ir�"RΌr2��!i��	Sl�C�<� @�g��q �I�o�Eq�C�<�c�F@� G�O:`{G�B�<�'V�v�\Kpύ_�s�[B�<�e��LY�����[V��IV@y��MX��Y�Os=����.�$�bP(>�O
I�������րY�xq`�E�
�I�0D�ܪ���1T	r8��O#b��B9ғ�?����ߘT9FL" ���~t�́���(�a��O��D�7���1�Ѹ�Rׅd�y���O;	���_��xCԯɔ4���9�'�*��Nڒ!Tn���C�]��:�'0�����L.�q��-��\<��K>����	�56M� �K���JI�ra!�$� }�vc��ѩ9�$h�L�9�ȓ@&>!���nBr���ʻ%���ȓ7��YZ��Xv�\IE��1��X��
V�Ш.�g�܍���M9$�
���4zV�i�N�.�v�Ӄ�ɒW�?Y	��M*5/��,���9����H	�'�\u���KxQҦ�X(�`���� ��@�.ʼN��|j�U��ո�"O��a���T)
tk�8j�1��'��\h��$�"k�d��c�;fG!�dՔz ,����xM�S���=�!�$[f��Dȗ�՛J���D�j�!��ُr����f#k�	A�S")�!���H(�TEV�`Y&@h�K�p�!��ğ=%���ٝPP�Z�oZ*\�az���\�4J�DA4��8*��-R�s!�B�R����I�%�<!����?c�!���!��[� �*�ƥ:�i��E�!���[r$ت�FO?��f�^��!�d�	R~Z��W*�r?��C 3U!�D�:&�a��,S�3á�)F!��e^ͨ��@� aQǎP,B�ax��	-W"<H�
�1ڤlZ�y�C�	��%�C�m��Y�2FI�A��99�"O�uR��](Z��0�B��y�Tp3�"O�٢)S8#�4�J��)��HC`"O���q��>$����@L���Bg"OL�M�����TJ�3���s"O4Ī��"b�� jG�J�8��C"O�-a5ŝ�;�B��D��aF"O1�%֭�Jq �g���@�"O�� �i��*�`3b噎9!�y��"O0y�a/X�^��BCWp�eP
�'e���D��)D<��րWn��q�'�4���ۊQ��B��z�d$@�'��l��n��i$���I� �`9�'�xx�Ra�/
p>w��0(����'e��H�A��)`<`�a����'D8m+%��jw$m�����yB͚3+��X�M�:`"�]G���y2ES���#'�#�Ʃ3`Ќ�y�N�fC��s���q�2�`��
�yC�9 FQ@��DAke�ꞩ�yrN��^	�F�0� �SF���y�gɶC�Va�c��(�ԩ:��&�yR�B7�@;���+JA�O%�yb;)V�H�`N�A��@�y��)+`|�q'G#2���X��yRa����M3	,��xS�O�2�y�C�O�>ݛ�1~�pu"�����y"��(w	�q��A<�8-��y�dؐX�2��"q��I��Ю�y�G.��P'$Ms����\���G�7D�l��aߋY~��6���X+�f2D�8a-3]X̃���B=�1���#D��b���k�l�J|\���"$D�(+�D��H㈤k�C$AM2�R'%D��"��9f�	@*�,C��ek0#D�l�Df�e��=�%�΍L��Y��"D��#���0hM V�ߑ_Fv�!�(!D�ĳD�G�<�d��"a<5�`i�@$D�t�Y�����ܒ8+v��E�ԆH�C��~-�� �`]#�� �W�-$��<��b�y"��X���$��X�"�sy�/��3vLX�!�O�(���,.�yRLA�ZF"tk��O<0�\��f�B�ICeq����^��`h�#K�O�@B�1��z�H i�`�W��w�lC䉼�d�K�BM�h��i¥���C�I�˄��0]��4�ݾx6�C�	&fR���`��7F�	��嚯�:B��@�ҝe�Ǫw��]ؑkT8�B�)� >ũ0B�Z�T1饋�A���P"O2H�'�<L�1�\�h3pha�"O*-Ch�u|�a���6N��("O� ��DV�*h���+�2��"O��p6G\�X0����\���C"O�y�V@M?P*��C�
��4"O������8AU.����P�D��D"O\\ڒ�mB���Ab�q����"Oz��4o��`]jP�v'1�t�K�"O�I�7��n��-�ԬF�F#�A��"OA�M�[���S5#H����"O���Z��y�f�T�h�tL	S"O�l�faYP9��hǇ�	X��v"O@���Ѣz�����(И�"O�L�d�E"H�|�I�H�`�:x��"O�M�5!�?�������)	��|�2"OV�У�!" 
uQ��K�/��a+�"O��R�	���5��*M��!�G"ON�F�;I�p�iD� 7n�" �'"O��hq��n����B�2 -�v"O�	2\�L�ȝ�p�ّ�&	�"O��x��\=�6���^�$1�5"O�4"�(L�^	^劲��)�ְR�"O�� ��S�Q����G(��"O*�A4g�sp ��I�l6��"Orؓ�J�)0L���%��f<���"O����#E}��x�D��m�,X3�"O��EB�j,�y�Ô���U��"O]
q��a�"����'4��9�"O������E��xw�T9AA"O��ᒃ��[�޽��'#,'��AC"OJe�g�*z�8��돣|/H�"O:����ŷX��-�J�)C	�u��"OPqY`/F1��8y!i,B��R#"O�D@S%UF1ƍH։�d
6���"O�˔�WJt����ޫ-�́c"O E���֫@]\����~��� "O����3\LA��V�4�Su"O>Ń��E��j9�MN)&c�"Ov٩�G�y�I�] b�0��7"OZ�4K\�E��}��늑5)P�9&"O4dsr�3e��a	����oV�1"O��ק�>���ڣ�BU��;�"Ob�Q��z|�w�1$K�p:�"O��E/] /�F�A�ƍl5��+"O ��EԝOO<P�U�2~�Q�!"OT�)��Y�X���f��)��B"OT5B�B�B��c��:�$b"O�����F�+L�ӱC00�j���"O��)�!T=���2k	 Z����"Omp`G&,�x����D@M�]�4i!�[�^� ��	*:��@�
	j\i��K\U+�����pa\�@ƪE>�ƕ��iȎc��DD��>\ \k�'����F�Q����p%�Ѣ)XN��D	@�V���M
�X�
�?U�0mZ�R�0��%PP���kB�=D��/K[ܐsG)��(Iy��.[��8�%͸t�����'��>�Ƀ~2Ѣ���=[�� T�N�!L�B��Jltb��͆Z���'�^6mI�LjܱH�EX��T�7Od�sl�/T���v�R(s��90�'{�Q�d�]5t`�e�0b�N�	׎�	
 �j��* �	�4�d	��
�$a�C��L�v5�P-�+s���Z�ɘ*Lft��^%/{�>�a�EӋ'�k����-D�T{��@p���COJ�RɎ4d7�Љ'��\8 '&�D���S�$
<�
}21fAM�����*ja~rA�4�V��� ni��%�&�:K�Y��Q�.R�� ��2CP��x!��p<A#��:eH�ȹT�M� ��.Aq�'�ք��$u �+��ĺEz�3��L�W��CpI��;P���gC؄����<�Px2�֯W���a+�+a���F�J��M��
�3#3`}i�S�ma��.X�C"c�����C��_������̖o|�к���j�<i�O00�>��7++��]���^"@'�8{oB�~�R��h]�|S�	���٣�bL�A��VX`[��/zϬ1#V��=K�.��1��E"�IQ)%�!�`�֙�|�[3LL-�f��Ņ1
Kv�� .�92���
���ٰ<qC"h���b5͞�	w.=��O�`�����*dL�A�PQ�[��` ^�G�r|x$�_&[�`�C���R�$� H��C�ɟ.^����f;�NyX�`ڀ	n�ْ%\ma,�Qj�r�1q`)Q�����:��	�ӓ@��"�D���Q�V�t��$#�h�<��$];c�X��Ī�`�@$�v�WF΅cV*E;M�^\Y���h�fѬ;t".�)Q��{I�������R�F0sSl�6_L�[�$lO�=��J�{�����N&O��}FI��A��-@ O�(��ɛ�Ο�g���`�OہK��2��|�$;��xeȗ�޴,?�z�0�I�"��cD��Gm�)0d���|ܬ�p��?E�،AD�O�`��# b�|�Z9���(>c�� �'�pS���
o(�����E2Fx�Z�	@�W���vL�kP@Y�d( �L;q%�k/��Ү�^=�;|��@������%1n��v�b�<IM]�3��!��Xjڨ DR!�Ι��Ϩ��e�5�̩O:)�;t�6и��E7|~�S���q`��1ߘ�Y1���z�����#lOB%�#o��1��EH �(���̒:�3���2����Ҁ�"N�2	aAҿ�z����}�D�+�0Z���ॄ�/���X�i6�I4w2�T��m�/c�vU��cV�!�zp;��H$^�b��*�D�8�w��5��}� Ɗe���Q�'d`tJb�Zu� ��<���%�%!봙)iу�~�A[ix@2���q�0�����;JÒ�b��

�1�R��\��U� �O��$��IZ2.�x����%��F�i[rj�!��\�'���s�BоEՈ��׉;;�	"Ӡ�*d*�4kD&	}����$��@��LHQo��K�}s�D:0��,�ªZ%;�@��7hP�{�i.��i�èЃw�H�i���C�T�>�J�r�e�ŎJ��O|����Ġ	RL��@�P�k&��fmָ- F� Eԫ��ذE�~�>�	A�K. %���Ya���n�΅��bX3����$�N�2�V	�N"�)I#��*B�L�DjRi�ԩ�Db�0����yG)X"?$�P���B,1{&�	�AF%�yªL�!&VT�^J2�s��Y>l��� �M���:4�%a!� պ;qn��nLaNR� �'���X7��=I@y�ˆ�� 2
�"�e� �R�CKRUA��IŶİ�R�L**�RB[>��򤌊�,6	�TBC<&(�	���X*ΨO6QQ��\�0 6�
*꬀��>iPL��
a�lQ,m)��Z�H�GK�,���V�r�<���
ƌ�~l��b�C]��i��8M�nԘ��'_P���ËR^u�b`N,a��@Z���,%.�,&��Ly�'�2^d0�2�U��M���/��
v�ͤ�y�+�kc�-b�l#��q����p?����.A��
��˽5��)�G*p���ǃ*���;����c|�� ͯy7څ*�K<6��-Q�a��t��W�O���p+�9f��!{�	��v�]�P�I�9h��L�5gI0��E.�1,p���֬D#�T�H�S�(%�ԫdK"�jTB�Ǝh�� K�l6�-G$Q��y`.�l�|A:ow^D1�bj����I�c*����0%����E�h�pl%w�⤰⦄;ޡ(�G�:N�X9p�lʥ�n�h&e�fw���T�5�O����a ��`� ,�=��d�"`D\��&�� ���@���Ňg*��p^� �	�`4�@a�[��Z�9OS�3.���'(��#
�rk�uyG�\-I`� Įߍr݀����s����aǉF���0��=>;�E�ᝯLz�XΞqۈ��Ã�rnSe��^���Qq]?oZ����ɮ4���gӭD}��Q޴+�l��cY+h40p�0ǉ u�v�z�.�&"jDZP��5y� zH��뚹Ab�04��B��O}�wē��ȝ!�oޅNe�i��hz[�6�����@*- �VOI�q��+��La ��Q7|E$�d	�seC�ÀA-�� �O��h����!3�������ږ�m���! ۖ�!9�L.jg���6����UQ�a�~B3m�7
FB���K 	Ѐ�lZ
}h��'bI�ZV6 �#�ԑcoh��dJ�!���z�!��H��5�QLK�D}��e�-?9�P���Ȯ�q �Ք:Wx���ȧL��-���>��g�~ڔd�'G���pĕ6��ݒ��Wa�'�}b��!OV�9@�ʙY�xe�A�Q� �4��e͎E
�h	3Ȥ:~*��צ����(@�.b�7�&�|���2�R*8�6��C�!EܼPmZC�H
��$,`tY�ڕ.%a����Vsc>�ؠ�x0D��bt�Z��U�>X���ʆ@�h�Q�����=9`+[�"y��1��+�z�ce�;��Y�G_q�dX�놽P���O���Sg��Y3�R�O\���q�hF�!�>\�����33=�O�c��p���
NC����5G��$SE#�yUZ��D��)PDS4�.LO��U�%�
������b�퉊xz��5EH%D?<�#�&�'@�P��W`W�>����%�SV���-��VC8E��S�? �h�s%M�+L��M�A��� >O�����!
��c���`�SP�O���ȱ�Ă \�}{F�ߐz�xp@
�'�\�u.�T6�8
�kWv���o�[�7�ƙF�r�qN��{L�3��Qi��+=� �b�	�*� ��	$A�r����P�k�	z��D8r���jr�ƅd����"D�F���I�]�4ٰ�d�&������,A�#?��	F�#0r��ܯ9l�O���1T,��DXL*@$5��%�'x�Q�4%�SB��0�
'�.�	�Oԍ"lE8_&M�a�>��?%��!8b�,`a���048ZQ(<D�h���Z���܀u%��-D�-�U�P�	�E��'U� ��$�Y:��O�1kF����H�B�"�:�@P�v�'��([F�	^谥�U�7U����I�7s}���u���Y�``C� (����I�h�t�#���>x�z�E~��ƙ&F\pCU�޻���������.D\��=�sMR2j4R�3�"O��F��/uV:	��ʉy(��X�����P�SC"�+!��C��#�.[�	2s$l�%%v`X��H�<�P��M�H���愊��@B�Ȁ	l�e��>OJ���Y"ْ<$>c�D�db[z�Ac�`��O?��dC �On�F�E4F�&@Ivd�� iv�⁫�Y9TÖaO���'MfљFnU(�2��+Z5������4p�L��A�Z֦���T?"  ����x3n�R6ʕib%)D��f�@�R
i�ơ�59�U��G�<9�ɛ���p'�ޞ)�?���N�� ���w��ґh&D����J�>��!�P+�9������j� �p�-�AF�U�g�,������.>ԀO�G���T�$i�#�B��Z`�:wH�sf]�d<�Q�'G�s�[a��u�`I�>R��c�$�������R�I--�3b�IS"��!I�RYDB�ɀ@�nl6)F�H2d ��$P�LB�ɛ>R����NS(KT�Q�5o4B剱u�Ε��J-;.�������W!�dA*V
 u8�dJ�[�����!�d�-�֕� �S�0�R���ÃA�!��\�];j��O��&�T��v��)�!򄓕�@��e&��QȪ9�M�~�!�DɁ����w��0C�X�Y���6�!�Q=n��!T-����۱R�!���d��Yb�Y� �2��"���d�!�D�"�� ��Ze��Qk��`�!��^$
3PC���=}Dd�g�D!��=P�򗇘o7�TR5�O�F�!��>;�8a營0��X��7~!�dR.�#ʄ�r�P#���3a!��>��(q��l��W�Q*~�!�L09+ݡ�E�?���t� .`�!��TK�z@ �+*�z�*#E�o�!�:Nt�A���ݤZn��'�3�!�X#�v�q�B@.`��80���!��
/G�z4Kc�P�CsjEC�ؔu�!�DD�Y�i����JPn�(7��Z?!�Q#F/JUP"�JHX�c,!�$�|�D�;�&P1�"Z��!��ڥr(\� 檜�h���[v���!�$��`VP�7��v����&�W�j>!�d��4ĸa$�21C��R-?*!�Sz�N��	��"a3T���'�!�D+r����<3�� �@��<�!�]	F��A���2��}[���K�!�$�7;�@0Iq̀�z:Z�96L�6�!��W8K��$��U��Y%d��Ī�"O*���*$z��U3R!ȁ ��t��"O����G;e��)�c!�*e�6LHD"O.!)��51!p���N�����[w"Ofi"��v�X�qƌ� c�~ �"O� <���A-|T�Q��/�"��6"O	PR�PN�sQbP�f����T"OF��`��}0� M�,y�Y��"O|�����B�:UA��H�5H��"O*��fϙIJLi�AS�I#���"O��q�#�2!4\�`>}*:3e"O0�  ��e���yU��6<wJ�K�"O��B�kL7L+E#Ηn����"Oԍ0��6�fEa�͏�rC�m��"O8P���?�* +�3y"��bV"O�h
����I0J]�u7�:0"Op����K���B����0��"OH�A��5M�b��F�lI�"O؍x2�_��6�g/�(/hH��"O�Hq�/�-�8d9 �ߢh�~0��"O��:��_V����p���"O��R�C)��4�$�-sUqR�"O�չ�*7X��.��5�$�+U"O�Y�i�<G��#~�0(;"O˶�Ԇ;�� �"(	�e����"O�hRD�ԸNf�%p�GV�ڊ���"OL8h@J%)s����`�Ҙ�"O�)2����JN�0h�_� ޥ��"O,Y��A�����"6�Y��.��"O<��5�\�,�bز��e�vBa"O��b�ۮp�z ��hJ�}w�\ �"O±x�G؃5q�����o<�c�"O�}�JΝl���Wgǻ,���"Oz�"��Q/4X9XT��>��k�"O�T�$0L<�כ��"O���hɉt�J9wX��'"O�mw�KL��h�.s�0�9B"O2Hy�kL�olK��b\*Q*F#���y��[@:ɫХE�I-���U�O<�yr�:H��фd�!Q� �K��J��Py"��/Jל�6AD�EE0	�El�<����4h�̰U �����e�<Y�84���+�E��=�F�K��b�<9����}&��$�[�<�! D�S. ����+��PGR�<y�FK	uĵ9Ꝺ���x�cL�<�b�]\�i��E:a�\���$�L�<�#S�����E��|@hè�K�<��C	�3��"T�Y�As�C�<�B�T;t��x��Z�|I�����^x�<�q��N�f��c\%���3Ҭ�a�<))U23$6���)�#S��{DdPJ�<Ѡ��_�E��㎘:��ѢB�F�<ك��D-�1���vH�ODG�<a��*������ݙ>h����G�<	PbG�5�����<�r��WʜA�<�1�Ŭ[=�U�GK�bL"|
u���j���݅Ub�sT�P�K�хȓ28�q�5՟*�P��jM�s����e�,5(௖^�L)[GJ��K�`�'���:F
Y�RK�z�l��4Zʝ�$TC��$���p>TƓ�Q�f,Vmͳ'�4(Z"� =���a�鍬TTB�	s�z�ʣ��܌�;��	�$"�#<1��9�b�b��U��OպY��ƃA4,���[��c�'@�y� �E5�Q��)�22^$�5����a$#��J�6��m����QR����XOQT���!��y��<t���3LI6G!8��p)�.�M��.� ^v��v�&	�Ǔb��(1�җz�-�5�B����뉆a�p�అ1Bg���� ZY�ٻ#��As��'��{@L���� �`�WŅ>;Jt\�w��9d���$�xό�/w�D�3)ɝj𰈈��	�i�q���kqMA?W��h� ķ3Y�x��"O @�[	׀��2���oH����뀱/��h��Y)/�����l�q��q'� {6➛}$Ld#���xA^%c��'��9��m�2�nQ��%A�x��[C��9s��,i1(ִT `���?2�޸7�MR8�����H����)M�4r�	;u#����c��dC�I�KLv�P!�pg9x�����4`���5=����Q(<񖣌�"��18�
�.�
�Ц��D�2a^��ՠq#��d�5��#�@������C��^����بc�jP��B�M�<	Q+�l�
 Cac�L�f��$�����/A�8��DI�K��%��x����`��K������@	)b�$�&��@ᒥ��	�1} J� ]}9���UIuƉ#��W�E�ʇ nTB�餇]�5�9� \�<v�T�l�����AQ�8 ���D���좠�+�~-	��B�7�H	���,�\�� ���V�xQP�JO#>�2<� k�|D>B�	/wp�sf�[.��`:%)
�,7��� �bڢQ��lM%T������ɬxj�;M[���м���#�0 �7� ���A��H�<a�GV�6�؄
��?I�e�u��pqx�:�*ͩ �>�{Q5^xE��Y�Д"�J�5L�VO����H��<$�ՉG䜩xE�!� lO��e��3��-����;4|���
L=�@���$A�`(�!�=���;@�
�Y��mxRDLF�LX�bK���䯕�|�tt�&��B�����1Td�F�R<Q����!a[+M0 1��;�,�3�zNF�� ��0T�sO���� `�����?-
^� !9˲=��f�?	2��R ԊF���,�i����S?	��w�ɻ���>Xd@Q�$�~���'M��@��J�t���{�'�z���� �Z�a���h���u -�W�Y��u'�Y#)(�QR2�KO��JB��I�i/= �fF3I9
Ї�	���0�Ɇ�},� `$Ƒ�q����Q3�D�u�Ǩm�c�.Qm�	[��ս_�p��Ó�t��Ė�L�6%xV��Z�Ra�>y�@:P�Ī1�ё\�,��d �"!r�#u���e|l#�)��+R�9����U�(h�q.G7@�!�	m)!����l���2�����&b�1V�4��A�,�2M ��k&Ce!�n����y�������ڛseաw^��yR���Ċ�QTK��l� I�(Z$���G�@��f,S�X��YXw�^�'����a6?�� R�"�
�(ăM�?h�2 _G؞�����UKؓpE�'Y��uK��1;yL�@�/�/�$eSw�4� %�cgE�c��z��R�t�џ�$��x�P�D��?M����d�)���}g4=8r��` �Q���
e�*���҂!�^,PD��*D@)T�.�J�oi�N��?�O��t�#T,������s��Ԛë��KLR��%<>�deA7O�.?�Ԛ�dU�]>ܣ�*W���;��i#0ПV����Iݤ7�J��"O
H`î��I�����m NA�0���� �^}�̙��ޕ����9+*���ᖝ%y6��G����Ӳ�@��
٩w��%����%lOJ͑¤\ 1r��>R�r�L ;I1ꔙ�C�5�ѣs�����ˤ�6��9���<9L�>�t�I�dBDx�b�X�nZ�@���䅚W0D�aI\L��Hc@�1��C��M3��ȹj�Fb�Gs$LA����������a��("�IN�n� YH�/	��LM��Q���Q�Q�,�ን���z%��ʦ=� ʞ#?N��$b������8\��ɹ���6VݸP�YU(<�������L�.g���paBѰki^x�`�ٻ&�x�b�/X&1�^]����9#�b�
�Y�/)��O��*A�dAvLp���db�	���'`�0#ң�RK��9rv���MU�d�Л�f֓.4��"ͭ�\]p��<j`r�B�����ˁ�VQ�p"��E�	g:�0�a�Ejy҄��<�@B�8-���S����E�!@l�����Y�$��W���j�-��nԡNȅ��+C � �7��>�@��I�W�T���
�u���D��)�11�-9n��<7M\�K���A�T�Z�����0v��	�J�#�睜x��܂A�ûr�b���L�;���D�;�V�k&��Q�Kގa
Pɠ$��Z��A� �]�p���p��@�M�܃e뛥��9��dH�d	�[��Mr�m��U��/�˦��AeH{�'�|���S�x�f�0�M�-L��F�G%Xi�\j�eH(.��t����P�5H'R������Os���qM$��D�T�O�Y�A���l+p��5�*���'V4}ccN/FBl�T�_�Ӷ�h6S�����$D�8A�F�I�5�� `F�F?�A�D�ܨ[���Q�a�i",0T�t؞ EI:~�x�(�"C�J�� ��oҡV���w/�*6\��jO#j�8�Zd����C��]zd�i�p��
y������>Y��B}���g�h�L�zUmԓb:��]HD3��o�V��͕n,�ʥ��7h2Q�ƍ�m�ā���)p�j|�^��8�%ȕ��]ڊ�D\�����@d�:*J�X0Ə�1T���U��?1f9ʡ��5p^��C�X�_����!i�3�h�|��g��$H����,��U%�I&�>i@�¼�4�Ra-S,0X��s ̯T$��~��M�<E�e�����@�ڍ+�����{�!��<�e#�'���>Om � 㘙l�\�!!!J��ˤ��
4����(D���'"h[-��<*6�� �C �0 ��Q�,M�����'Q�%x ��Y�Xb�8�es�%G�`,Q`EK�Bj���A�3D���Dծ(⼈���{���s�����L1��̾C+��s&���0Q,H8�
�q U�+��R ]����9>|8B	�'.�L0r.Πq6�� ��')=X@��O���e�+I&}�Q�
I"1��ٰ�xP��.G��L8G��!�C�	b�SG^�c�N����5����a��?�y�jD�l�*T(�)*��V'^;xlѤ�Q�B�B�sr�Uv8a⎇-M�`��i� d�=
���n&��V�9�lqH2�ܢ�>9�NѢS���`I\�TWj�'����ōL�x<8 ,С����;Fy������J�6q��g��!���"�a��F�ifr1����s}��7D�ikCk�2�ځ�#K,�'YC�U�!BO8��T�l�8#��A�ȓ~�~�31�E�:6ƙ3q%[�u����W;1�$�8P�ك�gy�3���/�h\`�愺"���RB�!����$�00Xl����ܱI�k3Æ�[�t��D��;��)�Ѿ41a}�K�E��<CVꇽG �i��!A��O�=����0T0�	Z�����[	hɪ��b"�`�Dj�2\(�C�I�ZnƤ�&ɏ�_��j�y���Hz(����a �S���m�O��ј󋝅:z��KVk�iA�'�B]"�l�.Kz,c�B�4��@�$a���1t-�c���g��6u15�Ψ4߆�K5i޽���;v	~M��	O�F�í�Rc��� n��(Qn�2���D�M�|�S����s�pPY�C�%ő�l*�\+y,��cJ����(RyR@�T�eFNX[k]m����ȓg#�Y��6����c�%�t�',N�X���z_���5�9�'!��F2��9��)�:M����9S��QF�
�P���%��'�l)�s�\~�+ָdI��b���y��6V�A�1N� ERh�Tf��Px�"ۄtI�CLP�Ba����1j�;���83�����(��zC�7�9�vo�9ay⦂<m(%zN<�sA�p���6�ؠ_�<�[�K�<4HL�67��ÁG}��Ǣ{�<Q��C����&O\��Ӵ�]w�<Y�K��n�#�J��i��t�sGo�<9cdY�OL2*�@&�r	K��j�<�S�A:+
y.̬��p�L�o#p���O~T�0�E�= "���&�X]�ȓ1r�����+gR=I���
jw.��e%�
�OhO��8u�Y9�� ��RL�颬хQ]�A(shΈu�\���U�L g��O�8Yå�t�f�ȓḽ#DEH qN.1X��ʍ!S�i�ȓ
D:0Q�V.���;�b�+����ȓ
��%q��| nы@��=U�&�ȓ5�$�b�RPf����)w����iN�Ő�AĊ"�F# i@�_�t���#n���+�5�U��چi�ڥ�ȓ�F����O�\�&�
=5<����`���KgH�F���4K��QI�<�ȓU6%q�İv�,�qd�-d�(��ȓJ!��y�ôH���S�6���ȓ%-z�%L
��B@mE�H� ��(u�}�wE0fȩ�!�,�Lq��.^��Ȃ���q��1���X6�=�!�91��v�L�-����'�!�D1>i�e��"@��Ph���"�!�L)�R��V���,pX�ґɞ�t!�D?��|�c�4~�Z �R�ֵg!�T0�2hC��b������D4[w!�D�v��񑋅�/�B<S1Mщ*j!��Z6\y�v�Μw��R��^o!�D��@��@���[�x��!�¬Q�V�!��P�#E�b�G���i�g�Q�t&�,$J�)T�@����+`��� (���L�)^���\�Y�p�3q�ҹQ��b������(�Oa����EZ��Z�g�X�4�	%S_�ȵP���-u~t��U�'P01����'����R�P�Gˇy�Vɫ�	 q�(!(q�A1~�x�/O�妟�6�i]'Y.��򤦖Q|�!;(�AV�q���>}b$�.��b?���آ�Z&&���"�
bN9��D �O� ƘzB�)�J��p�:j�4m�V�\03�ɻ4T��ڤ)r|��HN<%>��'��q�$
�0g(�U;#�R=	��LB��O�2{��53c*����:��uMRM�"Mk�<P��[�iՄ�Y���:!� �������&���Ȅ��}�qBO� ��hrP�K	L��	�i�2�;��!�_���92EA�r�m�Ԅ�1=]|m�˪<	���v��p���O|�%�gl�	��@sp���W��q��':�Ip'�k�����O�>q�灗	]0İa-ߐT ���k�yz��cL���	�P%���}���O� ��@"�Gט,s�
�&�L��/P%��sd��r}rj7��'L��p@��1�:�rd($Y,ĉ��M��ēH�Z������"|��״�# <�X�V"?�f �x���0}���is��b��O�>M�7L
O6^1
%�OB|��I�=YaP|�S��y����$�j$�)w�^ �� ��?��hB+F����S�O��	����j�0�V!�!$�@��� YP8�M�N>���o>ѲDg�'������.$���&[�KuDc����ퟌD��n	5z��l1��Zd>9X`� 9�yR���@�1�>O�h%?��'SVN�0G�|B�<Y14x0uU�\���S4���S��Ɋ�`ƢV��9J~�H��n����شB��3WɁ��4XϓW�#~�Zw7�L�v��~� mS.�
b��A��'�Z�'*��e�`�(VZ�"~�ŧ�90�;��N#/�h����t?���dt��d�Q�ȳ$I#$�a�O(f!�dS��D9h��!���o݁0_!�A�Bi�1�@9!
6ذ���,/�!�D֯:��%pF͗�?��"�<�!�D	�h� ӳ�W-l�lI�eL�A�!�䁛&R����Y��ռ��j
�'~d!���-JL�t����Ug�Q�	�'�4��s��oS<�6�P;FPzy�'j��S��*�g/�8w� ��'�y�fgM4<er��\#x�����'�&��%��<� �S���n�j%�'�����l%���EC�^�*���'=���hF�s�H��]<'_f��'ޖ��r��,2m�I,Ύ!D�[�'�J�����tq<my�Ԑ(tD�'�<Q��y�D��1'�8���H�'���㢈�T�@D O�y�Eh
�'u�e�U�)�t#4�R�k�@b
�'.^��$M�[�­(��]3�Q�
�'J@q���6'�ɺ�J�W-p���'A�D��׀�cA�I��Y2�'��dK]"?��%&
�=� @��'��� ���c	�)9�n�8�'_p���
�d^��C)W�/v�m��'��e��� e��8��IB
/<�J�'=��"�=$Ep��Bn�5Mdi�	�'�����֢"�ݰ"!�A͔}��'ArIZeK%2�ȍϗ�?(B9s�'?j@9W��Qc4x�e�C�xU��'�	�I�7{b�1Ġ�;)�.X�	�'Ӧ�ZB�PZy�c�M�1�	�':�S�$�=Cp4����-:L��' �:�ڔuJµ�s�	�� tY�'LV=`��X�`&�d�p
�8��a
�'��Rf�S;%�>ت���+�d	
�'�=ZT�1���1�BɁ'b�0
�'E��R��44J��c�X=��؉
�'�n�b�	� Q���
�#N
C���'|�-��K� LAR�>�R��'� (*3��?���VH�"�-�	��� $AuHöc��c�LЅ[9��`�"OV\b���P�<QAL���Pc"O�;ӊ��4� �b���"OX}�g��H�m[G�]-��1@�"O���cZ�HA�g�`��<��"O|�R�G%0G�-H`�A�=�Ր�"O4Xu"�=h�V��I�&�"4"'"Or8`�ʞo�f�is&�%_��"Oy`�� "J��@C(
a@�YZ�"OР�e�'�B��ݟ'��ʃ"O�<� ,�:u.b�f���= �k�"O�Rd�	�le(CB���"Ot=*��D
@���)���1����"OR��V���,(�aǖ@Rv��s"O��&&�`Y�b��6�p�rE"O��vm�5>t��P�N���7"OB���J��X�D�rO��l�����"O���%�C�U
�ȱ )��'�Ճ�"O$�Y��FJ
�pBr(ŉ1�X�"O~�1v��6_�R���G;"���"O��!�
�])��Pl��;�����"O�NX��nT�R�/@�T�y�"O!��1-,���U� �\K!"O0!�qU�T���	��F��"O&�Q�P2	-�C(B�N��3"O�!����B. ���2n0t��@"O� ������0�DPљ�"O�+q��z���`��_'R��v"O�iA��U�"vh���w�ޥ0"OIy&��6lL�:�N��"OV%򰎋~��Qa�"}gҁu"OP�JF/�l ԰(��! H�y�G"O0�
L�2�2�	�K�[@>\� "ONUhF�0�|��K��l��
"O���f�$�ָ��+
aGPh*�"O�RS�	-����!O�OАq{D"O8q�6�259N�C�%��k���a"O��d��>wV�&�>cʂ1�D"OrU�2�@C)�dĉ�<Z"U��"O����&D������n8�)5"O�U�F�5?�0	��P0r`"O��qZz��"�ݾO&�К"Or���Cʏ{���3rg@| b@� "O���Ѱ9�HZrFĖ;��8��"O��"�C��H>���t�:x�='"O�)�ң�䈴��.�6��|�"O��3$Ld`o�h�`�W"OP 0�GV99��
� (gۂ0 �"O6�i�l\�nLg�J�HXc�"O��J#�N�l#��p"�\���ѷ"O���"��i_�!�"h�r�^-�`"O"�BD������g��Ĺ��"O� !��o��y��f�b����F"OP��B埁[��
��8];^䩴"O�D��9\`0��5�F�'(Fx��"O��͞4J�uB�T#Q%�AS�"ON�C�B�#3��,�#@f�#�"O���ÁT�x�"U�с�n t�"O�)�C�ȹ�J��KM+n��%"O:��f�g倬�BK� $�VQ�"OT�Eܝ\~����5a��m �"O��!Ɉ;n��đE$Υwа]""O�u�'�
�>�룩�UU� �"OV���*��Ap�AY�h�����"O� �Di����O�$q�X��@�A�"OpQd�oĜa�@E��w��,��"O�<yǫYX���D��J]��"O��sf�]�B��!gJ^*%��i�a"O��9�&֎:
N�&�=�<�f"O��Xw-nk$1�A:>����"OT�z�(Y"�;�j��>���z&"O*�Y5o^6;�ٰ�	��|L��"O�P��&��C5��EO�9/Z�1�T"O:���M�{��h�m�!4@P���"Oܜ�����dI��ҏgxݢ�"O�-�����E���yl�b�B�"OH�ԞB�Z)�MܑI���3�"O,r ��.Z�0as��F�B����"O&��U$μB8F5*�#C�lg�e¥"O| ���,q�{�K�ra���"O�0R$+��0���*B	OW��T"O�������X��*
ܔXS�"Odc�/A(ɬ�0��	)}�~ŉ�"O���p�@?,��@E&o�.�ۓ"OR����,�%��aw�M0�"O|��q@�-L�rh*� ��̀b"O깫Q��G�ȶ�d{�Q"O^=i�nF�n��dH��%e&�;�"O���hԔ;dvܒ-�KJL)�"OBYR��Z�vj���%�A�"-����"Ob�T��̶��1��5�`rP"O>A�tk�c�]�2�߯d�l��"O�d�t��5.f�"6,��Pۘ���"O�P�!D	м݉#W/�.�2P"O�e�GGݒ�h�C�*�*	f��C"O(�r -�����[9!"O�� �&*���I�HB+Z!�"OT�{�ԾYX��HIXK��QT"O�[��`��ȩ�ME{?�]"O ��H�*�a F��4]`HhD"OT���Z�s�R��ak@V.T��2"Oj� �'�v�sc�E'-�!(V"O�YZ 
��{� e{�I�L+V���"O��H�o�"Bt��K�Hֵ�rრ"O��i��܉m����>H�XL�U"O��3B*��(.ez��|�]�%"O� ���A�+q�IA��I8(g\� �"O��	u(��G���
��F�BR��he"O:ؖ@<1�ig"�;DD��U"O1�3%�5l(Q�SC>�2!"O��)`j,_�I*� ��f|��"O��Ԯ�u*A� J:��"�"O�9�!�ߥVp`o���]i!"Op�z�e/��k��А�9�"O���G��iL�|:GHǵ!"r���"O�@�Fn�3)��Q�理.�0+�"OrL�֧_�E|�8sA�	M|TA�"O���I���|�nB�7'�|��"O$L9�@�[֬	'M	<G� ]*�"OlۅdSD~��K��A�<üI��"O&8b���`M��!M
�*m�&"Opp�O�^�Y�&
�;&���c�"O:�r�OƳ�>��$X�k�p�xA"O��C�NÉ}��&*�Z��X8�"OB�:7e ��M goE*B�؄	q"OƼ˴L	|�ˑ-�n���c"O�AJ� Q�5�Y d��݃!"O�|Q�.��X:H���EC��j$�d"O� B}
WJ��["Ja��Q�em�a�"O�	��`ب<��	b�D�2k���"O�8i���,�}1��	pk.`K"Ojq@��//��	�r��Z^8�0"O�$�3Ih5�]��6K ��5"O�i5�A
2>B�1��z��k�"O4��GJ>*`4�:fnM����*"Oy:qf�@殨i���8c��=V"O��"5���2j�q+����1 F"O^m�udѬl�<��UK��'�X���"O�4���3Z<)�J�
l� uA�"O�����<튦i�"�R�"ORay��*ע�h���*� R"O�@c� 
�F���)W��2'"O0�� K�A��AS�z�pH�"O�i�"c_#;�B�KNT�u".8�"O8Pq5���	ѱ�Nu, �"O��Gի`���h%���FM:�"Ox�g�r$�1�@N���ԹT"O�eEW�,D~�JP&�U�:���"Ov=�I�c\l�*a��oȂ�"O)�%�~"d���*c���"O�ɒ��g�6���J��\""O�M;�`�+B�����f
D�D5(q"O&4ڳ�!�ZɻF^����"O���!�ٺT*dd�4�1〈HG"Oby�
$F �4�ZQB�)
"O� y��%'�@�!U��8�\ئ"O,�!eC5Pp�YW"�����@q���� ׀�9㛶�����&�M��k_�~@r�uJ]9�(O���]���`�4��pip-ڣE��3����G��s�����S32�0��C2���M8�@[�@$B	��h��0D���+L����@f�*w��]����2�6�>�O�����M���~*`K`��A82��;�}�t��t�$9�O � �l� ���֌ԟ"}�F��WR�'��7��e.b`2`a��
I���(0��R�"�<�v�I,N����'zbZ>��՟�l�Xn$���)�C�T�'��5k�����6�hMY7�'F��p �A�PӠ�yڊI/���Jň8@�c��留o��5�FX�p�3��	Ɍ��U�{��"��N�9.�����$̄�M�>�@ c��9��|��gB+��ć	�'�~Q���b?�at�O(}���s̦uTĜ��4}��'���|jRmI�`��p����:��1/�z�'*�6ܦ�&�0��?>(���ƕR\��4/H�fz�����'r�'4Fu�'�192�'gB�'f���;-�QzV�P/�,�l�:=u�R#d�\᢬�v䈒�����i"�'(H��� �Dy2dU������l��� ş=hc�Q9ӎF2����ꐉq�y�M|�`˙9(��(�'�����_ r���s�7G�I UnA¦���;>yn��� ������O�6M؂2n���quΡb'E��[���Byb�'@��L>��n�,3���IR��_?4�i�26�+���q�����<�'������Hޟ0˞��L�d����wA�?����?�������O����O�m����2�@!�g��y��LE����B��C��a2dF����C/��30Q�PZ�N�.�@u�� �����(,�K��LYR���ٴ.@��Af�����'�ɠ3A�7-�= `����>�2x��A�f�شtϛ��'��ɟ4�?��U}Qc$��( �3���#s���'.a}rgּ	Ӣ���n�~-32�^��I��M�q�iz�	VDȫڴ�?���M;��N!X����U��2~l����dо�򣂐X.b�'.��D=nV�؈$��(Hf8M���\$9�"�Cc�O>恫@e��,9
���iݺ"����D��LR�=�Cg+Z��!��:5K�8A�%T�Ǩ!c�
1^98�UCǶC6B���D�.O2gk�2쥟��{f�#H�R\���5�Y�J���4��U�S�ԘxR��?�qR�j���ɸ��ۇ�p?	��i����"� �ix�,�f
b�b�# �ͧ)��I�KA���ݴ�?�����A�H	|�}�\����#�L	٧*;@���v�E��|b�O��1Jg�i��`�]����ɔIŞ��O��1�taq��@�J�\XХcV$��e8�S�&'ۨ�����S�Vh�`�P�QA����|���l�ڡ�ƲF�F� ���]���,6���	��M�@�>���Ʌ$z8`���+|<<@ĉ�G���?����?�,O&�d&���pcl]��GRM�`c��A>'�Q�L�ߴ~��|��B���EG,d��MP�\��(��-��4$����)���\   �   �  �    �  +  �3  �>  *J  lP  �V  ]  Qc  �i  �o  v  Y|  ��  ߈  #�  e�  ��  �  )�  m�  ݴ  R�  ��  {�  c�  )�  ��  ��  m�  S�  � �
 �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	F~2������4*�	p ���H�:�R�v�$4�H��� .�2�QNS�1"�/LOD⟬�aI�Y҂��v�ɨ/���9�G!D����U�LFQPs��r�eW�)?��g��qGI�'��-��:c��M��	Yy���8{�������rG�������o�#���<�I/î4���3E����@"کf��#=)1�#��EJ^��vE��<�"��ׁ�(�Gx"�'��9Ae�߁cI���M*SP4%��'�ִ��]A��h���QHj}Q�'�%yW�t���ѨYPI��Q�'�
i�'��4@⸅QAF�1O�JM��'r 2�LR�ʩ�#�1yaʱ�'\��cG��(�K�jGx��QH��� �LK�W�	���g�\;k�R�b3"O���4F��QQ�Ce��~���D#�S��x���a0^�A�cǒDl�B䉦|�@H��)^*����Y�j�<��Q>��P�U�(�d��O� a� ��E�D<8E>G����.G<(��hO�>�C�j ������ϛ�9�ʤ�4d'D�(p�E�9@�(q5�F l���Ǎ#D��	��I�P�x��̂gtt��4�4D�d�� �;M��������#3D�rN�7X�����߭$�N!;��2��j؞ȳ�ǂuq>e��ތY��isd0�O�扥G�z�C��-&ܵ���!B�B�I)w|�1�吅.�֥psn-�B�I�)Ĉ�+AƔ\k��i�Nz&�B䉐94ڌ�$�G�B�{�f88�B��^��4)uN�W=��	X�fC�C�I�dW~K&M[�>v�ҷ�ђIlrc��n�k��8�/�G��;WB�'(D!G ����$6F�p�LT8a�h�����5u�B�	�7?��)�f��k2���T�Z���A�'�4�+�y%�� ��=.̃�'�a�����L�F�M�,uPrM9�yᑪ=Q���� �E�B<!�gJ��y��ͨB֤�ɶA�E7ȉsdb�#�y2�-G
� Q��ƀ>wN�&�̉�y����LR��7u�$hF� �yǖ?gj��@�E�����OC��yr�E�u�<�y��W
�Zisؿ�yRD�Y�nDڧ�<�հPaL-�y��$Q,�`�2蟝|>Pܱ���y�E^�'Q�8p�8zg,Y6�J)�y2�Dk4-�O؛u?����OT��yBN>7���G��g(�\PL�������1?���Μm���	W抲r�6�j��R�!��P� d���M�e�4����')�|�O�� #�i�IY��l�q���y�I�7t���&��.����hY��y©�$����CO(t��@h$C�'�y���1���K̃�� $�cMT��y�Şb�(��5�v�R�P�ɏ�y2f�����h��r�j�Ѣ��y�Đ�uE�P� �Ir�\Xc����y��ҖFo���emT*o*|�SK?�O,�=�O�v�C��%@I��@�bB�2:ʡk�'�jy%Z�iL��{�k�"0�jMY�{�)�釆B�Q��Hʔ&G��б�9I�!�E5QD0�j�e6���ꃨ3xFў����'j�ti�/̙U�bD��8jB�I���-(�OQ(4���k���jDB�I�|��䁑�\�"�{g©0��Of�=�}
A���')P�ҏ�r�L�CC(�Y�<q	L��p,:��Շ#��(�jQ[��0=eҖO����+��� kCX�<�À�6_��1�� ��)�l��u�n�	b�LyR��~���N�i20���6<O��D"}���'��%ڑR>z�D��D��q�0<&���	�4�Dm�Hܠ6�x��oG�|��B䉢�&���!�8U~�1Q$�ZQ�B��9:r���`́�n{d���kBb#���~���"9"08Bǉ#:�DY��#`��B�ɹ*{��Sv.
����ՉVb�<��Iz�t�bg�ߚu�r`���$BB�����KZ�?�NH�t$N�U��Q�C p���L�� ���JX4 ��9��	 ����"O^�w� �xك���(g�4�(6"O�X#e	 `]|p�ȝ9n�T����	
�*"~�扜�s�Hj0�!�$Ź��v�<9����%%�DCXG���<Q@�)�}��@�iܥl���  �:u�ȓqS�d�ת��u0|�EoW�e-
X�' a~B��(��=Ad"S9G���z3CK+�yb�T��:�CR��&0꒹�%����y#��o��-��M0z��2m_�yb��k�@t�ŋҝ/�̒Ϗ��y���<$�Hx4. ����U��y��)��]�/_�g�F}���]��mه� �8�-��L4��	$Q;BƂ��'��ȇ�	'�rP��7	r��C��$��7M,�S:�4��'�&�KVBO?��x���{����'�, �ϖ96�0�˓;qiH�(O�Unq?1�{�����B��H�K
�H�Zqb6�Z��0?�(O��2���y��7��."�����$/lO┙�=@D�(��\<r����"O�k�P%'\a������
��5"O\8I��y��4#�g�XY�r"O�����y���j�P
�0�J1"OH�2R�P&��ɑe�^r�պE"O.	�⃁ �����d��c`HR"O�D8��?��L97䜤NP����"OȘ�A�?{�,�v�PeI"O��z��޾Jh�R����lf���"OlH�m�5>����s�K/Q��3q"O���q�1���d.��)�u+�"O �0�G�/�d@sP�^���aF"O�hƃkP�����9jp�p��"O�}����u;z�Â睬WR��"O0P�Ë8!�,A�P����p"O�I��v�F� �E0�`"O�s`��T�s�ݞ  YD"O�%y��zx��a"D6	u �"O4�BcI�)^���`7H�0h�>�A"O�eP�����#��Ŀ3Ty�a"Ofdi�-�%�u*�e *.��PR"O�<�DJ��4���J��F��e�U"O܅�g"�3 Ɣ��HpN���"O�غV��!~���'� 	�l`p�"O�m�b��[Fq:��@�����"O����*�15y�D�af>����"O���pDN4:3�آ�n�T��EP1"O��*�-DH���,����"OJ-�� ��d�����+P-(�9"O� H�K�I�CA�d�rY��F1D���V�A�� ��W#R	{G�0D�<{�@�$L��	�e���:+6=:� 1D��R6E@�>���5��*��Xx�#.D�qsN�<N*�!D߀DR���� D�P��R8o]�p�e��Lj�PH�m4D��A@dD$O��jqlёI��B�d&D���qN�Zˠ�� ��(m�p;�J&D�(��F�^YBu���B��[aG1D�|IS%\MK�M�'Z�%��'�-D��!��vxH@RO��� �G�*D���ROҢm熕3���?-�:! �4D���D���D Hĳ��آ_>m��b3D��D�	�&�S�I�Fv QP�;D�Ԓd�?>�����ҳ#�rP��>D�<H5�)$eR��O�v�dP�f�6D�� ����;a��A	��G>nAAp"O��b�e��,&D0#�O[=��b"O�uH�OX�L�ĥ�@��!6�yg"O�h��9:W���f��=X~��"ONl��㍉/��*��=5��습�'=��'l��'�b�'�B�'�R�'���F,�U��K��� a��=x�'�B�'W��'�"�'*��'���'�jA &b�Y�>5@EbۢӰ03��'��'A��'���'���'���'In #�'�4{��#V�S�4�`����'$��'���'���'�"�'���'*�uɅ�!��S!O����R��'2�'���'�2�'�R�'���'p��j5�[F>�sQ�� ,�-Ye�'���'��'���'��'$��'�$�2s��.yD��.Y�T�M���'XB�'���'���'Ob�'�R�'V�*�BI�2B&�R#�`�����'1��'.r�'�B�'T2�'"�'?�0!�b�p�}Dd=�����'�"�'���'G2�'I"�'���'��MX2�S=XP�Y{Q�צ���`�'��'���'!��'F2�'���'D�2�/�?#,ƌR�HH�i�����'��'���'�B�'��'���'��9��o�d����X0o�����'���'E��'�2�'r��'�r�'�v�Ҩ�R���B��r����'�"�'*r�'r�'�.x�d�$�O`|15�� v�Y�A�η%cZ\�G%�Wyr�'��)�3?)R�i���&��4��y{�$F�a�pXQ���{��4���jӜ�p �ͭ	�<�� �ݖ?��2���Φ��I,�6P���&?sk�e�>X��)��B�*G�R)�F�`��# �F�Ϙ'aR�xF��%؟?���4!I�]���O\�A$7�A�)�1O��?B���;e�a�B�)vիR�dIZb���S�"�i��<%?�h���B�R�I�Z�g�Q�ZnLQy�IT9/1��	�y����f�u�D�G{�O�a�Wm��*1�M�la�Yʃ�޹�y�V��%���ش9l�m�<�1�S� ^�yK��UI��m���D���'�
ʓ�?�ڴ�yrP���F)�����?(Z�dq�" ?�%�K.N�| ���Ņd�pI!��?A5�ьq���WǦ ����������d�<��S��yr�A�������J4N�JtQ�y2�q�B�sq���)�4�����O��Ȉ�D��U����5�~R�'G���'Lj@��HЇ�����yrI�v�!(�Qz� 
�A���["H�U{d�g�=��<�'�?q���?)��?�u�:�Z�K�ћ��|�Ҏ���d���}�'K֟�	ޟ $?�I;�j�h�óy%�2��ǔ7t�@+O���iӖ��X��?9�	�mPQ�D��w����ɉ\ܰ�U �c&B��'r+�Mdp�Ȓ!�������ڪ��a��Tˆ�	dӨE?�Da2��U"1S�`!����ɬ�bġ@>JN1�'�Yd���H"��1[5:���g��z����.�68� aS�"P�^�X����xD2Ajw�	�)u����;.��k���|��p��Aƽr��QY ��L,⡫���L��g�M1&I8\��4�BH�<	h4ᘣaf��e`ҭOx"�d蜁*��t�1�؛Er�K ݏq�4��2��N@��LN'v;�8@3Ǆ]�����L�2nV��?9���䓸?1��#��`�P��q�G�P��1�.�2��a0�i�B�'���' r�'��lC�'`R�'��Hb��&e1��ąݶA�Vy��g�N�$$���OL�x�FM ��xbf�mt��a!�u�2� %oS��\��˟<�Iȟ�)ďU��T����miVU�����)�U	�D4��H<Y���?A�8U����<�Ol�]�W#ҭy3D�0�e&��J�4�?��-�Q���?����?1�'��Ɔ�cD�$�5�EE^0�(��ia��'��0qQ'�9�O�ԣC����i� ʝ$��02�4O�\l����?����?�'�?���i9S�Yb���6j�@-mʐ~n�?G��)�b)�)�'�?�d	GT�Hذ�5����w鋲����'��	�Ŋ��'��I���aт�qH�m�(*5���Z����_k��m'>�I�h�	�1����h�W$��bcG��0�ࠒ�4�?q������|���'��'�6}d�\%~���
M�7����C�>��[e@�'���'2B[�h�6ko�c׀y�^	�RB�f����N<1��?�������O��d�8O�f=pU�LA�Va�E)~�$�����OZ���O�ʓ�����|��ƃ{�N��ML�dA��C�w}2�'#��'��蟈�I�z��'>��a��;
8��
��ԣ!�(�';R�'��T�t�B�F��ħ�M����6��ZD-T��P�Qr�p���O�˓�?��]�RI�|�E&ļk�@��,n�b�\� ��Jܴ�?������@�~@'>a���?�X�CMT�WAې�`�#�#�Kc���<-W��#|:�O�n4�N�2D0|��iP�~�ޙ��4���:�N�o�+��)�Od��I~"i�5;���,u��TIwɂ��M��?�&��?	�3�dŢ0�H�`B)3xYÂ`��!_�֨��n��7��O���OB�	�}�i>����ķa�B�X�C�0|ah�G�#�M��Bͅ����O����1O����0%1�0V�P,/�ͳf�#)�uo�͟�I���d΄
���|b���~2��:P"����L����W����<II�v��?q���?Y�� r8�c!֫qG�-@�a�|2�+�ix�D^@<O���O���<�cAD�"S�d��  Έ�W�]�T��F�'M��ȏy��'h��'���'i �5���F湫`�R'A'*�$�V^��6-�O����O��d�]��[�H�I�^F�X:6-��4.�e�@� A��(дNm���	�����˟0��Z�Ň�Q�27��1Df�R.G7N��1�F�{�"�nZ��������	ğ�'�"`�����^�:F��lK��H/�z�(��aӎ���OD�d�O�8�O�����oӂ���O��C��K$v�m����WTc��O~���O��D�<���f��ͧ��ɦ.��@NP��1��0e��6��O����Or�$�Rp�m��T�I�T��:Ur�q3�_Qb��J��"b4�4�?�-O��D�=Q�I�O���|nڈ5����CN�FSlГ�+�	`��7��O���H�)]�(l��\�I��(���?��I5�`�Ydd�qB��K�o��S�O��BXrj�d�O���|�M?�*R�â�e N�/&*Z�"F�g�K�"�����Iȟ<���?�����P�I��@�"y48��&�Z{��X��'�"�MC`��?I���?�So��|RM~���H���iR����h��χk�(l#�iq"�'F���-j�B7�O����O���O�n@�R��L ��.x�&�&X�v�'�d�)j��?��R������3Up�����A�^���нiTb�U���꓊���O���?�1� 0��C#�Iǣһ2���'�2ђ�'���'��'5"Y�0x��	7�M�Q����%���$���O �+���O"�D�E�X��4k1x�(u�ʋaꀀ���O���?�����-���C5>�Τ*� ��+`I�4��W\��	ٟ�$��Iٟ�I�s�	��>�D%��D�m�D����$�OZ���O��$�9���OF)BT�ݛ���K8}�g'�;R7��O:�O4���O~�CS�D�Pp�� ��;�b!@DaM8~;��'/bW��õ� ���'�?��'Xph��aS�nk��P�0䲗�x��'$����`|�|��j�P�Ş5d��t���ȅQa�i�剄Vd���ش������� ��d���s�X�j���!PV���'y�aH��O������N�wx�� ��g��UX�i�J��"bo�Z���O��d����%�(���u��	����Rp��"��v�4	��4F.`{����S�O�$?6&~E�1�@ Ar��s�)q
�7��O����Of�#�N�r�	ПH��x?	�$YU�jգ�ɓ�'U<݁s�Ʀ-'�t�f�b��'�?����?A�B�h9l�x'C�y�I9��X^��v�'�����#��O��d#���\��U�P;�f�Bdܧ'v�ACY���DB\�,�'���'��T�XZ�.�-m����
� ���#
�<I8�O<A���?�J>I��?)��6j���.۬G��i#Մ� b�������d�O�d�O���
`@6��5"�M��=���  �(J��Y�U���I؟ %���	؟�[� J���@�z���%�%>��� a+�2��$�Or�$�O��	<�Y���d��4r�t� n�
���/��,7��O�O����O�p���O��'�Z�rC��04�N�ZBΗ��^�AU�K3=�������+۴ޑ>�kN��T ۣ9���pv�C�8��L�ȓ�^�։��w��ذ蛟a� ��M��j�
�#w(�<�����B(�l�I(9x��P�BJr�Pt��O�l�4�5��#c6�}pW!�-F���D`���%$�MyzA���>*v�ථ�9Wn*��$�-CC��e��I�q��"F�r������)<u|`����?>����/������?a���?Q���Ve��Țt�J1��ӳ_��y	��دO�f=!�h�� �v�t�v��|&��� i��`��<cK,LR�/P:g����@�"Z^�W!5�B�>"��<Y�ˈ�e��P�
	Qt�ةd�w�|�O攱9O1��'+�1�⚤mB���w=3�P)a�'Q��ɖ� I�E�u��,#�ؔ��Ol�Dz�O��'���c��V��iu�Z9:��A�թ%�t�e�'6��'4�Bw���IΟd�I�~�J0 �fܳ�6����[�]�0�aA�"#�z3��1~�n}�ϓB֡;�l��yn�ѣA�^{p��F��c����!W�+����-U1��+U��7�T��
A�{��q30MJe����ئ�I<����?���m�'t��9A܋v��Q2#i��y�h�!YX�զU�#a�ES5��'�Z7���Ֆ'�P$��e���D�OP�!B��2��I6L��8I(\��d�O��dǎ\Ά���O��
��P���(�����BT��[3�$y�n���,�0#Ct�1Vb�'�:����:��,�A	o��\�c�\E�ms'��ES�� w��]џ����Or�D�<���6sC��� ��$�b�s��F���=Rk��p��q�7��)RW̴�-H]<ᥴik���`�D��LS�l�22��;�'剚I��ߴ�?������S1G���$�$i�*���@8>,��E��2����O*�r�����+cN]=P�!P�A�#>p�xiSc�|r���F��� ��߶nNPe�A �`��S#Z�T � $�e@|\����!O`�ӕ�ı���C�,r�!)�*�x��츣�^�:����M�'�i����F�Fbt8�p�B�G�=���zc1O���<<O^� �Ɠ��=S���#��(���'a�#=� ��IB��$�\��V���Z�|XA��ܦ!������ə]�4��#�����I����I��1��R�=-.	z�I��D��6�O���iK���3��d��n��_f4'?c��9T��=Xaf1�5Cs�R��Ǭ�uJ��D�?i\��Q�*˗D��>�O�X!7!!_Mte�*��;D愰S��զ�P,OJ�!�����?����?A񨟋[� ��B���S>��⧚���'Eў�Sբs�εO~�%��\�Iؒ�'�7m�ͦE&���?��'�JPӤ��9KT9�t��0V�Tp(���YH��?��?��^5��O���q>�8"-[�8f�]8T�O���0�K�Z��@!��zX$<Y`
���h����$U�:Y��f��>K�b�0��=D$�a)��PbV� ڗk�S@�T"פԏR-�YQ���U��k"�G ��m��#K�i���at�'�x6��{�	ǟ��Ii��N�Z�Ӣ��va�Q̈�:���hS~�;��,d�$�aaeƒB��l�<���i��^�\� �"�M{��?�EFW�e�(�A�X`h0���I��?��2en�`���?��e�� bcX�U�'��s��/4*=�`�P~m��I9eS��{N�njh�S*^;/v��A�-�,�H@�!O�\@�@R�'�
L���Rp� lӂ��F�n���c4���6+�Jʓ
:zH0�Z�MkH>��f̲8X��4�T�z�;Lp<g�ioF�Ȁ��H��t�wg��kT�$��g�Lʓ���r�i+��'��/k�,��I"B!@GП)���X�5��	ڟ����U���ia �X95zBxߴ7뮉�J�j�'?8�G��2!�rPcԨ	�?����O�a	��a_��H"a̘7�ΥX�b~��#'B9�DȠz#�MC1�Y^�x"��$�����O�6m�Ox�?��ď>i�j`��bhH���;�I՟�F{Z�(Ya��)�����eL����9Obl��M{H>�bO��FS5#�C8�����f��:����'���'�ltK�l��O��'��'m' �8?����C�~��1�i½yw�<ڐ��s8��ADF�T�fԒ4��2� D�T�0׍�x����G8d�2�#�IќD��U	�i��S4�i!���u,�C�]�Z�	:a}��m���Mc�f+iz�S�gy��'�t���'�S����L!C<]�OZ@r�B�:}��]������!Iv��(@��dݵw_8���<�/�U��3��]=���FVX�<�ǅG��~M�W��o��eb�z�<�R�T�`������Qt�T	��Gy�<y�ʑ��Uh�dY�(L�HyU�n�<94�N9��肁�!��0�ƕf�<��h�P���oy�~���'P_�<q��,\	: �fb�&V��f'g�<��Ý
]>��rb\�-f�6�Aa�<� �C�8�k���2�0᎟b�<��iډ��]rFK]�](Df�F�<!r 
7u��P�h��1��I�$]�<�G`��9kd��9��}��&\c�<�)Y/\��pq�c�F��p��Hc�<��Kz�E�ڝ6b�i��J�<�d�[(YF�#AIИvd(�y�#�F�<�*D.��#���Vx����i�<�0
.Nb�X�����RA�g�<A֦�Ky���A��骅aTc�<�� .�$)i/D2����u�<)aHQ $ qks&[3N�*E��W�<���F2��ŧ��ZT8irt��n�<y��V�-���s h����<��@;d�x�pǇO��t����J}�<aw�=An�M��, ^Va�/_v�<1@C�+>fY�@`F@
`�U#h�<�����1l�8L�,6�� M�b�<��D?�8BÒI��̑�`�<	����o��&�'Hq��P�<��j]����
QH�!`Ax���P�<���X���t3 f�!G�nTX���N�<����<�<jtڝJ�z����R�<A�
^�k������O��s��WM�<	�*��*��X�6�
~��aa	W��y� |��Rŷi�6�D�<U�ϸ'_��!��H��ȭ"PJ��u�B���&dV*!?O�T����L@�iQ��,8l%��2z$� l�6U �ɀg�F�0J� ��)� 6%��N�j�D4QD_�T�:D���DO�:E��mC2m~襫�CT3%�1O��"�BI�N0�y�a� 	��QsF"O�e��Ӛ �ha���G{x�dK:�0�V�Y�8�y��?�(��j���"P�j|,��  A��tD(D�l�e
(`�*�� �1R�*L�'�8�*M�#�ȶ��� ���L@Nb����ʟx�Թ��⃽nY��{�O&\O���d�K63|��U"
?�i�'㘏C���%Zu�p1Ƅ��?���8`f��4��#J�@ܘE��,M @H�Q��H>���*G�Q_OP���z�dh J"��
QV�	�3�ƿ{��I��H(t�.�?w0����qx�����W�f��j�Ύ�ltn9lֆ�4��Ԅ��m�����M�S�O�����=�AL�!��9{N\H<���s�ޅH��$
�F���I�{}r.E���OpM�$bD�?�����tG�� ����U)4�!�*̞l�|M��ɊTؑk�n^�5>��9v׻ �8���S�E��`e��`���%��ba�� <����!�<�[�a>�IP̰�!�
Y�v��;���#hBx�$Q��cB��?:�(��l��$��Ud�>=� ���[�Iׄ~v�lRQ��J������UtL�c���p<�qG�+�����(^]� [��[���f�ˌM�1O���>A�O�����x�f!� g��*�N���L=La}B's�	'�֙t>bdH ]�O'<�1��p�'#�b>��p���M F��L
^���B�W�v5�p@�e�iE�kN+}x^0��L�!��4�-������
X�+�Jp�q��<O���r�i�P &��0��,*�� �5�8ܺA@�G��:{��L�6���,�⁋���<� ��L�'n�hQh��ΌnӠ�	d�ɿRB�I��/�`4�Ub��)�6�)!L�$���BKM�Θ@��'*�+Hl5
9!��*nf�L�jϐb�@�R��>1�� �ɗpЂ��qGג;V8$S��eO|(�'J���<F4�K�#��ew�e�íԎ Xp�&�P͓]���Ok�S�x\J6�9��i5�	�����KGP�Ft��$�U�'Nqj�����h2��e�޴snz�#3�L�T����&=�LX9��D��ң�q�)����8�W*���s�!76��	����'��� �H 5��̗U�X�;�y��On�a�l�v��cm>%���2���9vJ�0eOQ�}V��Q���p<Q���-]z*<�6d�%n�T�a�%5J8�С�ҳ+�fʓ�M�{�J�i޲����S�L$�3��	g��,i�#�dZ��D���5�X���	��Т!��L�3��O�ju�r�}�H0�C�L�G�
 i���A��`/IRtay҈?r��c%�n�#A�\�=F-���Øk/�� �M�@��aenԂ��d)` �d�1fF��Ӹ+��]� @���.�ؠP��uC$	bPL
�O�I���&T� �Ӎ;t�����O�9O U�5�\*�jೕ�O?t�@�0	@s�y��A��,Saxb����j����	)��x��i�5i����ԥ(���`D!�>�g~Zw�`�2b�s2K�aO4�kr��!�<)G(6�Ob�iA�N!Nx�%�� �V��&��<�ꔷY��I�t��O��ұb妹hE��-[Q����2Z0�Y��]?�����	�r�0�[��MZ}��ڶ��`��K2B�7��X������'����4/�X�`�"�<D�M�3���'��A�	�2DVxܰ�d]�`x��9�($�dM� ���;� >4�-A`��-K����V:~����V��*�I�*2`��FZ1.}.`e�܌R4����Y԰�EgS+ZD�94%�:[��ܒ�I�6��A������]�N�9�>�zՃ��Ҕ,����'���1�L-:��dnX�2�ص��ĩ>)��i>���\6�)sv�\E����mݵ{+�$Y�+� ��!B	ϓ;��%[�#�@A� @�_�A ���rɀ�:��H[�d��$ �(@M������e� �S��s�.�W�m>�O�� �@��J&��1�+ �L5�V�|2�`+L4�Rk
+B��h�`�џ��4���@-4��Z���s� R1ALb8%�F�Ȍ5��:�� �0=q@J�6r��H3��-P�!�G$Ti!�tS���E���=�U�*,K�E�V����7�Y�i{@A[��' ���RiI�W*xbK�Hj���!kčp�J�R*O ">Qפ�-�n�Pb��k��3a�R�~|��:R.H�r"��±��m�'�LT(ׇ_���kQF�9�v���'V.Y��Ʊ�!*0̅
����	�`�	���@t��6�1O.��GG؀G�B%�$�ƹ|��d˗�O=�"a�����/K�,�Bɡ'����� UCub���>^��� o�+c1�R1�@'F�h��a@��0=)�*�e�Bd8D�O�*m>18��F�r)b8S�"Tf��?˓��P����p��,]��	��6��1��g�$PP�R�(q�G�̹����'�i��3�XʓBB�KR����
 ����R- ��$�Ón���$G9\O"�����"�S2�G8P��t����#	�2�j���?v{��G>?�Ѱi��7�r�:UxS큤(�O0Aqc��04��y��F�NkPAI�$J�u(�����;C���K2ƃ,8��i�7� he�D݊u����rF�,oU��
c�F �ԬZ�f�?k�4Ȅ��> �R}�B�����F \�
h$��!�@�Ĉ)�A ,����?�<نL�$CƆ���(���
uk1��-H��DB6T�n�0���lb�I[Ƨʹc���uXģ<�;qL�,�W�̑x��`q���Y�40r�F�Wܨ�i��J�az���.T�5��S��͸ъZ[�T͙�շc�&Y8�Kƹ�~��O�H��4��ThA%��(*�͈���,�'�~5�@f٢^{X�.�M_�H��r#L[�="�ȏf��-Y�c?���M3���v�,��֍R����{��C�`xi��,](��T@Z��8݇���l�8�l��,��3��^�4�̲��֪N�����!��Q��QԠU�g�1����R�T�V�;�a~��w-��4��='!�E�7��t ��Q��2��`���y�+.� ����ƀ	� ``ʄ�0{8�SC�F9w�^�h��#�Ԅ��)�:�ʸ��bW�D曦f
� �b8�P��2D� I`�Ⅺ���~�JE4u�x�ˑ�
���X�0�Kt|
Q�ĳF�`D�,�>���C�b'�4� +��'I�I�R�E?9�O�6��<
��HlN�|;��B=/�-s�4EEN��ř�/�Y��5<Op�҂����H�"�^�!�mP�BT���<)��>A��u'�A�:4��&މ>�E{ul��%�Z���ɲ+�J�o��2@�T�3�>̙�@L�$�|�7�`��$Al��"YfH�d[�� 
	Za��fZ�9�$)���M;�JҠ�d���g�<�$�)0�(u8�$�!0	:13�d����ò &�š��P�8�%&�4pu�V#n�����K�F(�m@�`z�4�B��?/��h���&T��4rq�&�x��BflȎ$���ؗF�>6�c@
$F��
ݫ=����g+,O���f�
?5J1Z �ߦC�T�$H)Ʈ�Q��'~:��'0�+� X	�6,����<3�5]��0>���м+GN$7Eb�y��΄@o聋/�Ǧ����3<��I�wt�D��S�uWe�)�J�! g���PA!�c�ިO�����>B���t4r�f��'+���Eڔ�Ɖ�$�4a�,I�'l�m{�O�X2�h:?�A�;>cDY�M�P~��мk�yqG�*28�P U��~r��{
��Q���B(2�SF`�պGz�/�<q8�M��0@L9�i�!��ˤz��	Դ6��^"�	�ߵ��ѫ��{�l��a(�@�\�':��|q �
�oͪ��Gޙ~_��@E�'/0���(��S�GA�Z�LB)k��	t]�A��'븠p��Ф��C��0�Sca�>!��@�U����Z��	>�,�#�eD�E�\v��X�:���-�yT�X��,HkH�0�� �D�˟�8e�qM��׮|�d��;����,T��c�ˁ+I��F��<��$f?��A��Y�!���S$���~��N?]�f�˖#y��C�֓'�R��0'�)��m;�/K�`<{�&�;O�������y�<���+��5TE��	�t�	�#ƃ	X=��I�A�Am:���ʟ4���43��͜Z���I�	[�jy�<�$�Pc��͇�ɳ�42�@��r��f�~ۘ�)ԭ��8dD�$�^�v@�3��]�	���?!'�Ϣ�x9-�la�@n7%���F�׈O��p��L��6M%?0��c�E��tA � �P�\��E�WT�+�mV7�����7����$�L�<dJ���Q��|ؠ�(Oғ7+�0��A�ϓBq$<{��W�<�Th�<X�����[�/��u���l�|�������hǀ�)�Y@�Ö�!���)Tc��6���v�%�l�F~rO�0%Q2�\>%�Ш$�#w��
WJ �a[��`.	�jb���iݕR�m�4���|:���;[�^-���\'^�� �K���,��	ߓ
��{���+cɲɺ@�҆3_�����Ҫt��92�$�L?�����ēK�.��ڋY�(�H���ü�EI�I+$�q�H܆{,�A�G"�}�'���e�]�6��#���Jb��U��nU�ު�x���(B�z"\c�P'���@��qNy�v��nj�&�02ah*HĨ��C�X36���~���Ą=[ټE��4!�x�a`��6�P�e/��(1fm�'���P�&G��~�j_p�j�ǰk4��R�.W�\Q~�h#�B��~����`����V�/�*�K����� 9��/<~��r���T�@�d�=�IJ���Q�4�!"�)S6�`GL�/c,����8+8�\��"�1v�^]�p�-$"��U��hhRaS��U�	)Q�ɧ#�hx"A̍�?A_c r	�� *�\���/@S����$C(��'i|���Xk0x����?��m2ר\�>qʭ�v��'����e��Wf�պc�d-�r�وyb�7_B�ɘ1�؁8��n�Lm���-p�Θ�d����Ub��g1��bd�X�S�ְ2�'μ�V�y��V�T9	ӓq](e�fQ�XQ!�+z� ]G���8� E�gM�4X/��peL7
$����)~=�Pa6�
F��!�"OCP&7�F�P��ec>=�3���%�>=�7��D�qE�4�@&%�Q0�ܩ�<up��D=�y2`ްOl�H��	˥�n|�V,U�z������?��˓%�|�'F�%��h<E�~�P�d�3Zd`M:�'��)v�V�ԡi5L�T��I��� h��b�j��y�#��=V��)�"O��i����
1h�@�%Xf"ON�p�_�6$����Ã.ډI�"O
�r�G�?9�%,� ,@ə�"O����J�=��ph���Hva"O$� �@SJ��uڠO��c���i�"O�5
ui��?�a�펢Uׂ��A"O0�A�1R:�9Z�<ό)�t"O A�dΊ ���3A�Ѧ\�����"O0�k⪖��d���?E���i3"O8$�vKx�jx��O�b!��"Ob�H�o%��w�L�o�<X�PDx�<yR��!U^�5d�3�҄�Ul�<�� O�����ჭvW~	��[^�<qu���6=R�1o[)/�*L�UaPW�<q��˯y�<�9WI�'R֐<�5i�O�<��+�s�
!@�*ֿjҪ�1�Ot�<ɰM�p�j�A�#R:yoܬ�F��l�<�&�V��p9yÂ��f�uB��f�<I�l�!@���h�؝-1��B��}-H�H��?PNƼ��Gˋb��B�I�K2��s�ɜ�oY����w�C�	���%�������O�u��C�	>-�_�
A��B-�C�I�I�m��h(aJȘ�#̣o��B�	%�Xс�e�RYGT���B�	0`�F8Jg�/*z���%s�b
�'�)�$�h���R�Rzt�+�'��b�,�=Z�� UOT8I����'����3-K�2Kz�H$!�����	�'��E@�iC%B���`�� <L���'dU)� �m)P��W+2/��3�'�|� M�V��k�
N�0�	��'�@M��h]�S��m&�Η9f���'����3*�\1�/��Up�'�� 
�!�?X�y �Ř�*��j�'k~yڄ�K�:La�h�l�N@��'[~�# ��<@�����۳`�*�a�'w)�4B��
	���eI�:Q�q@�'��$q�]K���u��'86���'��uQ�nʆH�T��JE�1�H�'�H��d��$w���b�'ݙ0!` P�'����`oI
^�����%���c�'���0��L����^��$��'NpP c��!�Ԡ�@ú���'2|b���1s^��B�Βul ��'���0޼%}"��#����'�P�S�
��V�!G�ޛK�y�
�'�J����J5 <�ff���<�
�'4��VL:9� j�'~�|
�'!���G��Z�T��BJK%||S�'��L� ��?]}�P⧇F�Tz�'*8h"��E#,���[�OC�PxC�'ΰ�A��K�O}r���	�I�p�i�'Y���XY[�8� ]�q�Pe3�'��a
Al�8kR���a!Tt
���'c��z�#Y[���W�![q*��':^]2���c�̨0a��VSzTh�'�2�Cia�ZQ��:��!�'�`�af�̠hx t��	,ؙ�'#v!A�dQ�o�\`v-��B��
�'�L4p��"Q����݈u��E�
���F'+��d���L�J�Xcj��y����r�@�uA�kb)0j�>�y
� (�c�L83��H@!C)zJq@�"O�I�1� ��DB�/�q�!A�"O��6�ɖ��U�g-��W�
g"O8���J(z�v  �öZ���R"O���L�/U� KV Ӳ(�(؁"OxT�fL�UeJ��Z{�0��3"O�h�sN�>A립1F� !{�h�@�"O��	� �<��5�P�A���� "O�e�G��,�6�xW��CҴ�*C"O���0+X5H6*��!�3��-�b"O����Hά.=�K��>�N��"O�y������dt)A?8�4�(�"O8q�kA3aD��ѣdkz�"O�� 2� 3p&4!�f]!s[4�"O%;�Cɜdy�(2��C�@�"O񪷇�(ZН��,�;�"O2(���D�%��p��e׆n��A�"Ov٣6�Z�[z���"������"Ox(���8��!R��n�Z��	v���ɉ5x�ʙ"�j�3�Rt�gM�$s!�Ą�R}�T���R7g��-aF�@�[]!�E�_��mq5���W����*�9�!��b�ʽ��E̖b'2�)W�١(�!�D��*;����L�2'J�x!����!�ϣP�P��wL��:��Q#�-�70i!򤀩V[�d�`O�m�$�	���K1Q�\G��HY�z�OEe�a)T�5�y�)\�E�Z�1�
̃Sf������y�i��D�ґ�
,MXH�U&N�y����I��dy���r�t�#4���yB
U���k-p��cS����y��+K.���Ι�X��lJ��y҅��k0�E��L����!���yb��(B�1d⏔9��"E핧�y�đ6#��%���Ӻ4D�$�T�¿�y@��t�.l!G!F�u��e��'ת��'`�="���q$�C�z1��'��s�d�,�������4D~dk�'VMY%��t�D���B�.��x��'�D�	-D ���Q��U�s�Ș�'K��	���!b��P��܅�Ȳ�'��}�ץL�x�}���#vE����'�ƥ��#�N��[�
������'�J�i���PH�Q�C����	�'�t�sg�^&`��xH�� @O�P��'il�c!τ�;�cK8&�Y!�N%D�`������Y���r�`@���G��yB�לmI|mA6)1Z���H���y�@E�h�A���PM�!2u��#�y�����T=kW� U#����S��y�i��g.lP$��9U��T�Щ�y�N��2F���⋳5�m"$J�y���1G+��A��B�(vt�P#I���y��T�O�B])6(X�w[�$*C�į�p<��DΘ'�ы�۫y��s��@
q�!��ż�T ��2B\Mi#���!�DW )��t�FG�I6�L���U	e}!�D����z��ࣇb�p�ft��"O"�0�"�Ct� 1�n
��h���"O��ҷ��/.����ŤQ�g��8S"Ox��EK�-$�qA�C^��	��"O�*r� �.��@��jĒl�"OΈh�d9$ %��Kح��5R�"Oh�`h�/<��Q�A.���`"O� ��s���/�����o���""O�ӢeZM��X�#U�D�`�"O�(� `�0
��(��D�u҅�!"O�Y�`�H^��6͒&0� r%"Odȣ��Q�ᤨ���O�}4ca"O�I���@�3��Uȁ��eVe��"O��:���=��i�Ƈwa^���"OnT�1�V�WD�t	"'T�+�&5"O���aT}3l�æ&ۘ!��5�5"O���G�N���p�ɥ)�v!y"O����iF���:���X�6���"Oz����+PL8XqkS�
���b"O\0hgL�- >N�+2*�2I�|<X�"Ox��5! =9��=��IY�B̠�H�"O��r�-�F��5	Y)[j]��"Ov��!��yx���,Yi�"O��R䅭l�`]��Y#w��X�"O�����!_*�j��{%��� �N�<9�!�j	��n�:;ڐITDK�<!��+;������DV�y��VJ�<�a0i���Q7ZƆ١RC�G�<��[�Q���qiD�|����t��l��p=AO_+BN,�e�c�,���l��<A���p���B�Y�R��h�P�<a���X.\����<�t0�挙M؟4��>����df��}�֌1Gd��yR��ȓ0�d}1���Ҁ����̑��>q�Tz&�S�`j�m	vlH8k�(�ȓH) �	�M#~�D<YP��i�D~��ӗ0IQ���C�- n��
[5��B䉖o��8��T#�pP!�N
*F�C�\+х+H�m�.y5Ō�Ks�#<����?}�̂)�FҌKj�P��c9D�p�Ԍ] )��R#�-{����H6D��Z0���~��x3�Mϋ�0�A �!D���p�SH� Y����.R=�P(4D�(�F =�iSd冫KZ��Z��1D��34+�;�"T b��|z�q��/�a���\D��h�4U,����e�3G�"���]�x���P���hܨ��P��Cv|5�0"Gp�&p���:ä�ȓ�` ƃX���GN$*!�ȓ_��`�0�k��`
�����ȓ>z�(bX�$�9jvI�MC����3
���.�>����  	�]�ȓ4��C�Y/&3�Eq��Zf��ȓ3�� ̖8E~�1�P+4;�$���ɂm�� 0����v�4lVA�6�B�	9X	(���WY��ح�C�I�cL�Ā�4Xf@4c֞{u���O���#ٯT��0�LE!�D�2�"9��n�����aaؠ!�$�y[�eA���'�l�+��ܝ0]!��fX3�dE�GA�xc �5T!���s��=A�k�0΀�0ԉmP!�d��jP�I�V�4m�n�1��]!�>:t@�3��b��찲&�
�!�$ڨmE��T�A<�ܨ��}�!�!Q�^�P�NT�G)��C���!�
�l�@����O<U�>P���!��F?-��ǪL�]�]#�!�>%�!�=�Р���%{\8b�.�.3�!��	P�zpSF�"E�iq�"�!�D]!�pxf�� Y�]���9W�!�� ��CM�|K~,�v���3N���"O|����Sk��#熘 n����"O�)�)
�!#�а��c�@��"O�(��JvM�梓�t�*���"OZ��DL�u<��j���7�e�T"O.]!�kE�kS4<�a,,���"OytkZ(Nl���M�G�tx#"OB b�	�'sF`��T�
O���+�"O��D���'��u�����ۦaze"OL�& ��c�D4U$ј.�f)�"O�D�H��\X�4� ���8s"O�Y�v�3�*��c�X+}�Q�B"OT�@�?:4|�s�o��ܠ��"O<|�aʛ�"����C�K5r�ȑ`"O��X�Tm4A9�n�^q`�"O$|rW�I�_�ri�"@�y(2��"O�HT��x���	B�ۃ4Ɯ���"O��&ѓ>�țɆ�*�h���"O��(TE�f=�qց̖�x�"O���@�fB9�TaO�#t���w"Ot$
���uhB1�R�+(]�@d"O�U�V.!�@�	4E�;`B���"O@��iM! `��ӓE7���P"OH�`��ڸ.��6��-&N-�"O�A�@�۬�����F�T�JW"O��JBo+2N��k���"O�x�V��OBZ<c�l0"���q`"O�<�� ܰ`�5��\a��+�"OtE�zF�r���hM={�"Oڼ�q��'W�:�JM�͸u"O�Q���9v�	��5V��&"OX=(��	a7,y�ef�-����"O���4��?���3E���" m��"O:h`D���y�`죇�^)_<�T��"O��{�h֕o
nJr� ]Jz��*O`M���G &�|��[ig�$��'u��2�^>08D@�� \�w�$9X�'�"Lr@�-h� �ƈ/C���
�'Hb�1��J���H�)7��D;
�'��s2M�����0��� "�*��	�'��Qr�ٶL$h���B.�4�!	�'�n��qDϫTP00�KS�rp��' p���#&���g��2`� ��'��W�\($d"	x.� ���'�ؠIP?-�[��pJ�AS�'�Y0��K~0ݒ���.].x�
�'R�Œ�JT[9<�GE� /r�2�'���B�L7eᆙb�GR/�����'�vE	5`C�>��ࡷȝ�z���{�'���o�,:>$�g��~IY�'j���)ǅ5�Y[�)FM���k�'5�u �	5�t�wES�K��<z�'�@�&�[0U5�8BDa?H�&4��';���pOȜ�N��cG�@Ȁ���'6�l�L�QC"���J�k��`H�'܄1��ό �<��NF�T��c
�'KJ�����uDA���GyP����'J�ccD�)3�H��]'q�Q[�'C�E��
^.HQh �ܺl$�q��'�X#�嚈>)&Q�nۗf�`} �'���q�����b�a����
�'d�`[A^/?IV���[�
Y�(
�'���8�*bj&}� ���	:�	�'q�0�!僽 ���@��5u��p	��� �Ŋ 惃qZ�p*�i��!P�"O�x�'Ҝ�F�A6 �g�r��6"O�a�`E
���R�Y�'��%@�"O����Xp�	�@ʹq�.���"O�h�Q�
gH(J�O i�p��V"O���t(@4�^ufl�������"O�Y�o�56 �+���G�$9b�"O��iT-.(�iы�: �yrA"OȜ�f*܀-�x�!("e�l�S"OR�r���N,�ͱ��!�R��S"Ox@����0�aHT�sCj�#5"O��k��0e ��+���(I?��s"O(���ݷ~��Cw憸o>�H��"O�Y)t��j�օy�����pv"Op�3��'*<��j�AņD��`@"O��qb(D�dY��Q�B�]�*}BQ"O��r%(,$te��B9$�X8k"O�(�� ĂR0�0SD�C7[��cT"O��ࣁ�U`��*`"��CG|e 1"O�pv��?xp����1�]s�"O8P�!T�t3P�)�J�	� 0�"O��2�5WR���C/A~��"O��F�j���Q�H�"O�軑ʌ=ck��@	�:u�����"OV<@!�ǬX;�TH/?k�|�@"O�}�ǉ��p�ї�0��K�"OD�(�j�54��CJp�A�'3D��H,�a��@��T�^�hu;Ae0D���!�ԝ
��ۡ�й��$A$0D�RE�J6B�⽡!��)��Xy�f,D�d�rH_�B��ӒK�:1�D�11)D��sG�\���܀p�*)��|��m;D�dK�/<ې�j�%AHL  !:D�pB��_��L�#�j�3|����5D�$�RD b�xE�0EA)u�x�,0D�|�geZ6�p1:4&@�.�X�Sׇ1D����B���*���/Ȏ�[ĉ.D�\CC��L@D��uH��{R���T'-D�|7�7O��Ԡ�噳_~$0��7D�p�C
�L
��:"$E<4U���GH!D�d��M�N(9��G�}|�0���4D���� �
uku�B4Zk�M�#�2D�ػ��� )p��SVd��:�a8�b/D� �ns�U`uJQ�H�
X:V�S[�<тƁ�vL��C�iݠ�b L�<!2��1�,%����Y�l�c��b�<y� �v�ܡH�N�2�l�§]�<)�
̅1o<q0��y�	j 'M\�<YB&N�#4zC�$&��yrm�X�<	�*I�jl�t㗶zj)��Z�<9ϝ�q"tbc�6�V��b�p�<�p�՗D]�t�"ʳYz�@�# j�<!�˕W2�g�ů$��0*l�<�p-��Q����E�h��(���q�<	'�3H�^�����U��|��D�<Yv��
%JJ!j ���~tU5E�C�<ApIԪzU�A��Z%y�`xg���<ab�F�-_�u���9G0��[G�Fw�<A���
w�@P�DD�>�D��"q�<�Wb"(2�B@+I���aG	�k�<y��i��)�n� <�����f�<)��5m8��갌Żq��4�/Y�<�P.�*)Y�R��S�%�Y�\M�<�V԰��)x�j��7f�ɰD�E�<� �Y�Bc���̠�ϮSs���"O�5��D�@�ڝ�pJI�
�-3�"O�-��B�N R�(��"� � "Oh���D�""b�S���m����!"On8s�j�3>���4����"O~�ӊ��\��u���Ii�ݠ�"O���G�%G��e[�IPH�IE"OȽHV�N�N6�Ix �k38�q�"O�P�s䟜Vr�l#�i��~,�M�"O��)a�U�zw��⳨_6=$\1kT"Ox���\�~lV�Kg�!<�`��"O$͙�+��\���S�M:�����"O�Q2���0Mv�`���H�"T�u"O~R�J�7.钙8e�G}T��"O\@{C �Da��F�.k"DH`"O�p��>7��I��ǠZa��A"OVU�E/�u�d`(� �^ب�"O,BU�F�\�J�H��]��L�3�"O�萅׸�BQ�@�����`"O@���=7
v�� ʅxZ��G"O����*�&��	�:vv��"O��r��l��Q�f"aKy�`�"O(X��A�^a�m�g��!e� "OP��O�H����F	lJ��A""OV��P'��R��spA��y2ڐR�"OJ��$6��P��`�.
����"O����Ͽ�zؒ�)}�H��e"O4���N�	G(�r�_�ڡq�"O�Y�̻C��d��0t"OR̓1��,0�����>W�0U�&"O��beaڛ0�D�y�ŉ(޸�(�"O� fݮ&u�|I@����ܝ9c"Oj��f��{�6��ѣ�'�J�b�"O�i
��Ñc���!�zʒe��"O�a1&�A�A��J��կ� �"O�	3n��:�A�P(�6�
m�W"O\eBs#�SSz}��Z�&��,X�"O��2O=f��eB���nQ	�"O�͠a,��~���r���13�"Ö¦*`La�7�]J�¼*C"ON<ZG�Z�og" r�[C���h"O�@�v�՗A6�(�^7Nf�u�!"O����O
k��8fЌLL�e��"Oh����JJ�X�_8Bŀ�"O�@� �ԕ l�۔#��$�ٲ�"O�,�
B7�r���A߇f�f��"O�U�#X�L�@h˶a(J�*Q�q"Opo!f<��1j�Tc�V�!�d1y�����?�0!.M�!�dT,��+Ɲ6 ���/��!�I�S�KӍX���r(I=����'�L�����놭� "�'���`BO ���6��Y����'?,��� �1lF�V�����'Ѫ��SA�7����#����@�'�2���!��E�0��`=���
�'J��j"Ο2#jU���ӧ��!�'��@��	����@r�W�s��
�'�\��@h�1���K	� 5@
�'W<�gk�y���F�Y"m���'�P=���_�`Z=&�2����'>v��`ʙKT�!d�}8�'��8�SD	MT��R&Q#*9��
�'�@�t�*&����	^� g$����� ���pKS(e6Y8�����T��"O`U��0J���E䖳1����"O�9�!/� ��!5��m���A�"O`9B�nG���ږ�W6%��:s"On$�q�[�(��*�Hf�TH�yB���(�r��3���Lӟ�yR�������Y�:�;�*Z�y�a��3��S�J�|�؇�/�y�Q�L���*&�>U�q�'����y#�4.������-kp���F���y�ե�e���A?8.vM�F���y�,Đf~��Ϟ� ��H0�-K*�y�`��+�\�"�,&n�y2m=$�v��B�gh��m���y�D\�����X�$�*դ��y�Β��.H E8HX24(�`N��y� ��1�D��*�.=�u��m���y��Ǯ^�@��1S
�	Q�X��y҇����f�	.��a�H��yboMy��w��1��=#�P��y"蘨P8J�f�-8��q�P�"�y� ��rAp!>(���G��yA�.�����tX|5��E��y�L�# `]C�	{�d�ʧ�y�۸d�e�(z�2i���U��yR�ۅ~�%�E��, K1&_�y�LQ+^P�4,Z<	 N�X�㖭�y�Y�b��dS�8ʼ@e���Py�ᓬx���r� ̶{k�+���J�<i2�Q�k�	۱"��Zq6lSE'ME�<ir�ʾ��0��hR-vh�TS�dJD�<q`W�iF�qqѦЁB���J�fR~�<AqKC�	�\��W.̂�L�"Rf�<ye� 2HtE�����6���ەl]`�<i�.�3<��uAς$B���E�<A�ɓaA��h�G�T���XG�<��s%�TH��db�E��JB�<�&g5"�z��H�#gӠ���hh�<1&f�b;��j��[�m�����NI�<y%��4%���U�%'��1�B�<Y�\�\��Ki�<m��v�<�4BY�^F�9d�^Fl|X�ÀY�<�Ud ?Dp�h�㌗U(p��@o�<���B�v�@B��8v[�Pd�o�<& ��EU�ͨ�%��iD����B�<	�!uj����h�-?켌�ըDA�<�Ӈќu얄�G%ְ~
~p�§�c�<Qd#�1N���f�N"Uҡ� d�]�<�bE�����/Z�.o���R�<Y�N�-;��ӯ�4T�����G�<���,�E5��,�:��UcG�<)�$IL�s���)�vP��h�<)��V��J�T@�H�٨�yB�p0�r띳Jl�������yR�E*'�Hs��'xM�9�@�,�y�CR�B|�`v+�l>�I���1�y�J�-)
��b"a�e�.�AT&��y"CP`�(b��,������y"��Gưk3�ʩ6�<Ҳ!�y�&�i�|�"q��\�H���	���y��Xy��S��N/��K��۩�yB.���8�T E�Fqd��`] �y�IɊt�!���7p�@�I�-K��yrj� ��T� �Y�h�l���)�y
� �e��D�a�9Wk�d44���"O�0 ��ZO�N��).��*`"O�M�b?+�p
�$֏ ���"O��w,��ܭA%J�8\	d��"O D0�$�"1����ACU�y&�Q�"Oڠj��B �PU˴��3/`S�"O)
0�ޫ;���
� Ә�	a�"O�I���$�DXzf"��T\�R"OV�+Z�2�C�
U�	�J�;�"O��R5� *���"�J�xt�|!"Ox9��/��}�G �H{�}��'�^���A	�2r��00�G8J�l��'C�qk��D�`�&9���Fr� ��'m����.i� !��N�>F�m�	�'}FP�#�J�!�rU��ᆎf��3�'|�1ĭH�Z1 i�J�E�'D��[r�^�qw�}k�� �'��A��!$���l%	��8�'�Ш��!�YX�4����*��	J	�'讑#��fBF!Fʉ,0��`�'A\l��KM�&WZ���	Z�J�'I��	7�Ͷ+�� ���I3tTPB�'%�8�5A�! �!��/��%6��`�'�2�xb̂�g�����)UL��'��l+�F� 4\�!�I8�%��f�<y���5!�Yy$≊n�8�P��`�<��"��1�U9b��x>f�ĂH`�<��O�5�6�9�:h�!v�]�<�#)�S$Pp��EHf����X�<Q���zh�|��Ő�*㐭��BQ�<!�i�E&�Y����6�VLKpi�<��O NLZ̓GC��J��+�`Xz�<Q�@az@A3m��1������Ot�<�U�J�Dh7 H�#���C��m�<Yu�d6X�aI�A�aG�f�<�t��'��ժw
�V\R�q�_�<9��R�#�_�U�"�i�a�`�<a2'�& �@���B-l�1�J[�<A OIU�Z��!#����` �S�<���#�$�9s�!����CLZ�<AV�ӻ>�p��w�$�:E��k$T�h�MM�|%x@1�� �#"?D�����~L�꧂�nhHLz��/D�lc�/ɴo�$�&N�2L-&�x�!D�d�fM N�$<:��ūw��8Y" ;D�dZ����P�h �j�M�بZk6D��"EQY�p��� 3CB�l9%�0D�̒�	N�L��f�� i��$�tf4D��1�fNP�Qiوv�����L&D����
��~M�t���Ĩ\�l��Ѯ'D��q
b������v��I��&D���bV>o�N�jshH�^
�d�eG%D�d���M+��K���N�LXǯ5D���#共%�
��	�7,�P��2D�8ʗH��d��r��'M����vO2D����G� I��P�aCEHE�hQ��3D�p� �#1N�I�@�F�V��TM0D�8�gL��E�t #EH'T( �#0D���bX�,� �d�؏`���$�+D���Нq�M	��Vw�M蕂*D�D��*��,� ��Al_���rk*D���+yJF4ڢ��'nڭ���&D��@��1Se~�+fȐ	u T#�&D�HI��I2+������C����A?D�� 
�P��U5,gfж��o�$"O.@��f��	`Rp�����HuR7"O�%�ͷB�b��A��}�"O��B펽X�az��~3D�S"O�*��� 8����d��UD�#�"O����٬w.ޘa4	�<2��X�"O�k��L�l)��H���Q�8|��"OȑC6#Jb��8���>�$��"OL���dxF8Kp�B�B�B���"OШy�F
</|ƼZrB1a�d��	�'>�����p��$"P�Yf�<�DK�gb��sq��bqՁ�@a�<��,n�m�萁N�9PB0D�8����N�� �p��f%�@�Ń,D��p����_i8�{����nB����"*D�`cG�p�� ��N�H�HW5)TB�l/�����֘B�>��CK	<E9�C��Ò!$L��re�f�Ƨf�C�I."�Z����I	l������vC�	�#�8y���5@L�!��7s�hC�	�{P� ��B;f�
�Y� .R�B�I|M� cf�h9"!i��I;6�nB��_y2ؓ���E�	7
+6B�	?N/TУ���r��x+��B�C���ˈ(xAL�9t+ˋ���`CJ=D�\8G�D�x-[G�G<.~.dڢ!D���D)X�X1��/Z(X���G>D�h���)L2���QYN-`��)D��[��V����Sm�")�(�S�,)D��Ed��?�հ� P^���4D��q�τ
Ype෩����a��/<D�`)���g�6	Q3�/�8hqe�8D������{F�%�gM��R�C��$D��as/ųJ����\aH`��.8D�pZ�c�*[��A��R���ݐ��7D��T��9�:YK���}F�����5D���"[$�99U�S<V`����e2D�)Z�2��YU��o������2D�[񇎩0�Pm���h9f�0D�`���Ԝ+�Ҙ`b*�5d|���/D�T t�=CP�����	1�ty�"J/D�̀�I9`�qH��^*�&yb#j,D�4��*A�c -�SFR
]�DuR��>D��pa���:��6K�O��d��(D����k �-�(I*�b�H���h�f<D� H��adF%���4�h��.D� �C*�w(^1� ���&�Y�&+D�H�cD�:�Ù ~�}�a@*D�4;�mV%GC��"�;���נ&D��Z�'���<�9��ءUԒ@���%D��	B킧=�rXYϗ<n�����!D�[����mDX�q�mR�*ښ�[En>D�����M`��K悑O�^�Hr&9D��)����l�c�N
L56|r�8D��x ��$j�Ȭ�"$�%]�*�1`6D�dpE/ݨ!U	Qw�;�`�B�3D�t�S�N�.�^��%����5�V$.D�LHRɀ�T�Ҕ� h�u8Ν���,D��]	�<<����8&Rp�F�ɼ�yb���݈��S�7T�aCB��y����k.��@x������5�yBo�/U�d��p�ښt�%�dR��ye�S����ՠ���L��@��yb�(c������E���}z5�9�y
� �D�K�N(rt{�#KG��{6"O8��D�~�B@��d׆+dL��"Oz�ː�)t����
5��a"�"O8\�a-Πu��pQ��n��8�"O��t�H�k�ΠS�"^����"O:hp�MF�z�0���!ŜM�F�:f"O������-b�3D��s'��"OpY�!J�&`x�.�5|x��3"O^���Q�:|^)i�2WHuÔ"O� 7��F�mY�lT+R0���`"O8���EI�oȞ����PR"O����E�>#�EѠ.��2�5:�"O�� ���Su@l���R#���"O�i��P�"Pt��N���ɺQ"O�-q���ZP+�.��q 
9F"O����ʹRm��Z�n�2Q�i�&"O~�3fÁ����DK�,�ت�"O�1��#^������h�y��ɂu"O,� �'9��h�U�H�0�@"O*k����(8�8�@/����"O�����TN�����d��"O�I1�ƼU ����ͤH�%F"On� å�iJy��T�=g���&"OuC'$O>Ix�cU
�9N\`��"O��@�E�L8�EJeB��<�^!�"O��V	�Nƨ��ABB����u"O����-2�(tB�E\��Ҧ"O 4,	9Tq�eʄ%���3
��y"��;n�-Av%�  !���ޓ�y��չ&�z�s	���>D�uG���y2�zA�T+c�µ�`U	�h�%�y��"_��be*TX ԑ�K� �yb,[:Tr\�ԅV�Q�hTa�Y��y���'_����B�~5�˖��yR'F�4���P���Ar6� �ʋ�yRǘ�	�"���N9/�*ڗ���y�%޾e.}��
]�q��P��A
��y�KЬV~��6nUr�������yB�т5��܁���Ɇ�P$��'#(��aML�|Yy�n�b�1���O ��`�Q�l�L�Bɺw�`}P�"O, ���u�p�c�M�Z {R"O&��E��H@Ҝ:�É�_Tu"O���J�MY������Cp����"O.�	R(B3�|P����21�^d��"O���!���!1�\��)��-�"O���s%�T�V�@�U���"O.�S@"x�R��Α2���"O�$ʶƚ�W�����%o�Ѝ��"O�a)A�)W�(�V�M C�t��"O� ��h''8�D�/.�~�1e"O��@d�#���0�U�w�Z<cr"OR��`��6d)�N�5.���"O���%f��F=�K"��S�"O��	C��v��$�/��1f"Oz���H�M0���jɜcp8�2"OҘ��a\�쉳��)k�\��"O�����8��pr)�BF||!�"OF!rÂ�1xL �!4��1"Ot�з�R����&	�7?��	"O���c�
(ȵR L�'4<qp�"O��Ljd���P�����"Ov)���L+�t�8��*V�z��""OԹRm[*0�}8����-��u9B"O� h]
0�A�1���с�$�X��5"Oj�zQ!�?�-3fA��(p����"O���'A��a��<���_�e��[�"O,|S��9�H����^�J�p��"O(�PI��hV\b��ݣ�|q`"O*�ZM	zr����+=j�m #"Or�����5<��S���'��s"O�U+�&T�$�PT0b�àu<Ȕ"O��R D8^*�Y�'P�b�hxk"OlyƁ ;	l�UH��. 4N5��"On�h�)߀VS���ŭ]�a��T"O�iJ����6�޵��됻O�����"Ovp�5B�q�dz�*��"��ͣ#"O�<��C0TJxݘ��6Y���`"O�)�怄!aJ|U��(��E��I"O���B�4Fl�L�G��E�05�7"O���q㋑#iH����8��#"O`!qg��8]S�X"�_!E�G"Ox��e�
I�|R��ڮQ��zw"O@�e�N�q-���w��JIl|@�"O� kv��?JT7OC>Lм�"O�Ӡ�]k���s㑽���Z�"O���-�)�V؃#�ׁU(�1(�"Ox5�PO�	����er��x�o"D��{��\�"���S<ȆPy%
=D� Q��P� 2�� ��}�����/D�P� �O9A����Y o$T�Ci0D��xf���Z0+F&W�q���s�/D�$1#���Y�)&�!!���� D��	�.� ��Ш��Q2�p���>D��YR���np����N�\V���<D���W+�-a�peӁG'np8
!h9D���������tZ��W%�bd��O$D��#C�ňv'��3��T�V�v��$D�d��!Z�W*lJQ�QcT^x('j0D��V�U�(�m�D�
��N�Y�o,D�p���<_
0�ŀȵa*����+D�8;�M/����@�2)�&o+D��+�+�^��h��\_/�u(�N+D���`� '.ŚDsBa\�cm ٧�'D�py�%�;[�Ԃ4@τK��Z�&D���R�P��U;t%��N�� ��/*D��ؔ��*Xʝv�X��D�T`(D�T��b��\����ҍq����#�'D�����ι8�xe�%�hb1��g(D�t��ǚ�B��]X�m�78e9g$'D�$G#G2�`�f�;{�<�H7�0D�H 㐅<vA�"*��$�fEb�� D�лQaR�e��᠆
�d�~�{5�=D��i N�s�r��@��;E=��o(D�tB��H�~}r�1M�X<�m���&D�؛b���
iLA �N�-e�]�Ь?D��`�Z/F

�Pch�x]��j#D�< W��~C�ۧ�'.�X����.D����)B�e>~,�Љ6_�L);1H"D�sp*�O��0��E�/�N�!�	 D�<��S�]�6u�R@�4R� 1é>D�P���͡&��A������O/D�����]���=C�<�I"i+D�L��Ը'V���N��0�S�)D��@��V�>W�=K7������R �9D�P v��<�H���ޤ������3D���G�&�i�b�Z�'���y��/D�,ڣ���n�*�uKD7u�rdP��.D�� �J���,&���!/Z�	&��"�"OP؀ȋbt��;�`�5bv��U"O*���� |R6@ȕZ��Y"O�q"�c�(��"��>(��-q�"O����$V�JF&AR>�B"O`�2BČ5|���@��
*{��U�5"O�0ʠ���v��x�	�
$���BB"O(qɃ��"��=���%!F��"O<A�.F��ۓ�:8R�ISF"O��Rh	/9��)[��ѺK%8���"OJ}����k�b̻�H��=z/�y�W?HV��p�\�U�dRq�Ƴ�yRM�E�0T�׆�S�.!�G�6�y���5V�Iɳ�@�Pv^,ʇ�%�y��5^�Z�ꆁ�9K��p�EG$�y�AW8\�� �wl��C{�U9�FŜ�yBM�9%��ԡ٬��� U
���yR�E�|��L�v�^��D2���y"m�(]����fІtE,@�P����y��z�lU�$�	/U��+ 0���'`1mS�&��1���98��2�'�b�2UF�k����AS5 ��}��'$��Xq	 	��C/�D�Q��'dv���H:"v%
@��K3��c�'N�аQ	�'NX�c#,)X�L��ȓGX*���(^�&1��&�'
�����>�)%)K�F�t���̟$-"�A�ȓN��X�%��G�sv&@(�!�ȓ�0|��ª\PB	�d!oo���[�X�r*X�8:a0��kv�ȓwv��R#R��HX �3��X��!�4Rg�<g���vB֘%� ̆�W;:�xe$�{�f�2�����f��t��	�#Ck>l����&��ȓP��(���ڸ	߆�:���6�@���%���V	:9{��@�]�1���Z��ӵ�ϳO���d��>G�,���)3������$ZP���W��Z̅� ��5I8?^�jsʟ�v�5��lG2Բ��,[D<٨g����ȓ���q�O�� ���h������N�a���|�����gH;D�8���&�p� �Qذ8H�AZ�}��-�q�IKlD�����d��ȓ���s%�\�B�٣�ŐY�J���`�V�3���N�����QY|���1�ޱcs @�Ei =Sv����Q��J{�Q��� 5�!��CIP^��ȓ0ڄp�=w���˄pt�@��+�L̂�ê;sؤ� e�(%6d��@0�¤��9�l0�T A�f�:��H
)jiߝH���kK���A��i�ne�EN��T�.A�%J^���j�ԅ��|aD�R��r\,�ȓuQ�� �`�ȹ���X�� ��(R��Df�%t���b��!�Ε�ȓsL�pD�ܚ{�l@�*@� $05��1��ݒb�^yI�%xv)IA��.��P�F�֝�p=�G������ȓ5�ҹ�A��f���Q$պ<��L�ȓCU��٭"0���-C�_�xD��jw8p!w�@6{v�����wZ���>Nt���B�"2��;PJA K�$�����ƕ�j����5d��9��S�? DP�mL�"6�4a���L���[�"O^̙b�&L���c蒺[�Z�!�"O:l�e&�(�"%�W��1ʾd��"O���JG�K(1j�B���<"O�t�2@�K��� V�A���ڗ"O���F�r�>pg���9��!��"O�l�'ўr��z�n�Đ�!"O "E��;���CՋԒ�Aȅ"O����Ń�P����ާm4I�"O�۳�8*?ʀ�󪟏	ԃ�"O4!�U!-ہ˓1�0�*u"OZ��A�"C�Ҹ[Kޤ�Z�2�"O
<�`�Z� G�YH�gν��d��"O6]S��?&>����#BҦ�(%*OBh��e;G{�U�Pm	�[#@���''*��#�O�66�u8ЩD+i`�ً�'������[W�0�_H����';��mE�&�qÅ�P�$ȁ�'*���⏹B��<Z�m�Q�hYx�'w��!�%mdvțf�:G�\X��'����p���\�@e��İ95!S�'� �f�O�8�,Ģ阗	w �P�<	�'ݡ4�\8��\��xc�[d�<����";J�1G��2{`R��Q^�<Q�c�41(] U�2���)�Z�<��D��E�\�
���I░�D(�@�<A��+zrD����cÂ��/�f�<A&�GH^:ꅤ2F�	��W�<���W� ��qoD!0n�C@� S�<�0� %��]Cb� A�N��DR�<�ge'T۠p	E��"DqY�UP�<Y��x���qWL�!Z 8q��Zc�<��e�9�2Aa�� C�� 3�^W�<����V�`h��P��Z$�^�<!QD܅WJv���_Q��IB�TW�<�fH�p!8�9�OЎ�\��Rm�<�3"J2�|��#�Q
�jͲ�i�<9g��1�6\c�I�J�F)u��p�<qA
[�]��0Pf�.�Dss��k�<Y��S� v$1G�Q��+ F�f�<	č_�~}���ܔZ�`<��M�<�!���E�:=Qa-��o: �b��T�<1�Ф-�8L{��;�ԡ"g�Y�<����lu�9 �ͫN�Dlb"f�T�<IT��"!�Hp�Rƞ-;�<�p�/	N�<���#CD�"\f��#��J�<�!�m���Ԅ�R�>x��BF�<i5�E�u�<u0f߽na�(��DB�<9!�	dz��
3��)ad/A�<���.g�������+�R��&I�@�<��(�3J�8�{��K��DTDD�f�<	-$dtHqҤ��-7�j���m�<�G�2qz�,�Њ�4+�\@FK�a�<� �M-b�@C�o����V]�<���_-q��H�׌B#Nf����W�<I�+�h��e���N(*Be��o�T�<�§ɥi���cQjm����R�<�aD@3G��F���j#�36����[f�X���w$!����B�|���!���*��J�{B�ɉg�@�i�t�ȓd�L�@���/����B��64�L��E��`�"��,�"UbFF0R0�ȓ=����`ɐ�r�Q@��R��N���-&k&�����6&(��S�? �@y��r��J&�πѴJ�"OR��(�H��k�
��s�,�["O���d��\��@��k�;���3A"O �0%�?E�]$��?��y32"Oy��ƪD.�8T�'|2Ve��'�)6ĕ�pR����F75�	j
�'d���I	�f�]!�Ν0����'{x�2E��b7�� 
Z�.F����'n�= �퇠2��x �*�D*�'�xE�p���`��x�/�".	B�'J|Ċ��ϟU�|W�^ ș�'M`�J!���w"lГ�
�)l�(�K
�'\�0ɀ�r�. ���G��@�a"OD�S�х@ �aQ�lV��0�Q"O.����G=�h�"IT�q���"O�c"急����`L;?��ذE"O�Ȑ���.��<At&*Vi�,�r"O>4CQ�^F.��K[�!@�"O�(�i_�S��<C`*-�^С"O��Kݒ$��`�d�)��-�C"OZl�/��p(��&i�gf^��"OL07]�̩�	�Z5{�*O:z0��NU�����(S���	�'8bCO�%f2�p��> r�H�	�'�d�ѠS�#����5�Zy���	�'��-B�(,غ9���o��e	�'p�|�B��9\�u�$��8�1��'jx9����jK��SiM*�=P
�'��xH�G%N��1�>tQ�0��'�Ÿ�3��e��@�p����'{<����)�m��.��f�@:�'���tmZ��J�@U��'~����'�X����>Z6ly�b�,�I{�'�dA ��v^�����&��`�'sBp��0W̐P�g8[�&��'z~�"D+\�>l�ү�*T����'�����+��P��d�R}t�@�'�.)`����&*f8i��Q�%�]�<iv��{��e��P7��E��Y�<y���|�t&�
��`0hPT�<�Ǌ.�6�OS�m����x�<q���p<Q%�؇&���[㣜~�<9� FG�X�@�O+n7��K�|�<��(\>M��u"O��
��@mw�<�vd��L�,�B��7 �L�<��B����;�H'_����Q�]�<�um�(��庰@ g����kIo�<i`,ЭMR@����A��9�aB�o�<����1c�����ˀ�3�yR��Q�IՊ˼Y�ːD��y���>|��ç���`���p ��y智e��q���:XF�v&��y���B�0W6ظ�+���yңI�䄰�(�Tf�j��3�y�W�!�@92�'F#X��(e����yR��
��ʀNQ�H�V]ɤȈ1�yB��7p`A�Ӥϱ	Ȋ$�®K��y��FJX��)	���R&���y�FO��&(�*~�h)��A�yB'�k��Yⶄ�}lb|C�̞�y�%�
x���� ��n�p�;��y��-T�1J�X	�dS�*��y2I�<9w�͂� ;��+wص�yb�0|̸� \$��
n��y
� \\�Vcy ~Y`�`ĕ#o�"O�,SW�jG����҂gY�ŋ�"O)SE�ZG
�2�ؔdܢdqV"O���I��d�ZQ���a�0a9"OX0�	482�
�@��t�:�k�"Od���)�޸Ȇ�>C�.u"O�T�<�1:�o�)a7���V"OLK5a�6p��E3QaJG*D�"O�͠%Ȇ90y�pB��d��"O��X��	.���,9qy""O�ɐ1fުC��R4�Q<]���"O@pc�ښf~�J�O�� $hBg"O$ J%*@;C����3E���Fհ�"O4�;�ɲ�`('EE8Z���SS"O�h�s�ŦQ"�p`�Y�(���"OD�c�R�8褸�V�&�ڌ��"OF����f��)p芢U�v�s"O���"CV��噁aL/W�L!��"Oh���7N�B0���r�3"O��q���*�u�A��j�Ð"O��Z��(,���CBiK�� =i�"O^Ic�i>+a�5)���g�n�R"Oh�#��K	RI�@���[���X1"O�$����C�{�j��aG���"O�-@���7'T3�o:)�1T"O\��G=V�L�3b�Ÿdݼ�B "OvaJ�<p��H�m�\�03�"O̡�A��P�
$K��Y
8	RP"O�Z����8|���<���"O�tJT�X'e���J�Z�M�hd�0"O����٪8��U����W��y"��cB�Ȓ�'@]s"��t�N��yR�)��URր�R�2�r$����yR�S�L�t)򅔂P^���r��y2��
5���@�D=(|�a���yr%߭]:����"G��*�8'4�y�Aoz���7c�V,��C`X��yB뙷5*�rWCŠN_Μ:�N��y2.T	N� �0���	s�PJ�'��$�C%�%ru�aC)dP�X�'�vY�g�I#
(lP0�@�_����' ��p$,�E�{�,;�	ԖXC�I-HE0�ڦ!�,\�L�0$�w`HC�n�f��ׇ	�K�4CH�0�
C�	7[�ly
��A2���:�#ͽ]��B䉉s>��7&[�=�M��W+w��B�I"b���	¡O�v�69�I�+!�B�I�3�~��I�![_,��r F #|\C䉛�t� D(�_;��2���q��B��.����Nu��)VqB�	w���d�9%X�Qa��sR�C�t�ʄ8�e@uVz�H(�4uǚB��/J��-��J�]�n]��=d"LC��F߰X�Rׄg?2�sa�Й^tDC�ɣ%$:�+�"�'J�e�M�7%�C��[|
.�R�@�J�)�[��B�	�[�{�c]:}�B��eT)?M�B�	$3R�1��$��A��맯P(g�vB��=�y!W.�t�Q�L�xHB�I�`�J}�e�\>��zW��$6(B�6y~�`��)0���!a��B�	: ���lΕ��@S�@U-�0C�IZ,��x$�Z�r��Q8|`(C䉱�����.�
u��p��UU�B�)� ���O�
��W��2P hP�"O�DH��R�>͸驵�@'2�Д1�"O���'̼��$���@]��"OD��g� 9C? 	�TD��'J�I�"OTB���a��ip��ֹB�@j "OP��uh-R��"�I(H�dIH"O�q���7��%iI/:q��"O��seaڢ0��1E.�Z�)c�"Opò�ڟm�H�H6��s����u"O�4��FД/�-Q%!����"O�l*�6`�ͲP&ߕ$� ��e"Od�'�J�t�>d�p��
�>� "O��h��s�yc
T	2��`[#"O:@�Q��2�*�sg�*'��Y�F"O�l��J9R���N ��ѳ�"ON�!!���oW��c����Q"O��p���O�T��aÚ6b\i�"O���wC�QY<`r'��F����"O�(�����d�ٱ/@	KE�ݲ�"O�����i0�M�qڣJ'x���"O����g��rFE�]}��"O��B��J�z���0��]�Y�"Or� ��Ph�0��*[hz)x�"Ob����J�g	pE���F�z���F"O�I�Ӌ� |U*=apA��+
�3�"OҐ�W {�`�* 'Y�VlL�"O��2�퇻SY.:Qy�qI���!�dR	�����IU;i�Xa���S5K�!�B�=Bj�Y@�	v�aU&V�=�!���#eIbe����:��0x2�
� �!��W0�(�s�Ͽ+ܔ�񆌃!p0!���0o}��b$HBp�,�Zw�Л!!�P (p
؂R鐪w��l`�
Y?�!�d��M��)���ֈ������4�!�$�K� Q�*ƙ_��.˘-�!�ʩb+�	"#@λ:�5��E�G_!�K!L8	�!Hѣi��"�&!򄎩s 0�a��G���k0�̻e!�68�VEr%
yJ�)CbO�g�!�Dܵ;�� �Ξ�`7|4���M�!�O�7@� Sm�,/��PQ��!�ďu�Zis��%!hq����E!���4K��IJvg�lj)P���0h�!��	8cb��D��脵���1=�!�T����BI�<f4�������R�!�$��^H!"���jZ$�Df�v�!�dٜ) �"㝏�l1qӯ.2N!��8s��A��e�dc��� @!�d��k{���U�xb(QQ!MC*X!�@$|Ό�`�I7%+ ����N�!�$'i�@0��,<t�9�fw!�;<91�F�P)"����P�!�DG�:,�W�H�k�hs���!�$u,��v�Z1Ք���.Y�?`!�˟>�v ���p��q���QM!��ڑ(�±a�������[B!�5u��Q;f�!L���2)	}6!򄟄e��Y���-Zb"=�fʟ�G5!��V-Bh�F����A4��G�!���<�h�����%��O�!�dS*Df�i5-�,2� 0Oښfw!�dبb���*��R�dZ�l�.q!�$��2в���B�M<8�K LX!�DH�.��,�M�<R`��C�A-V!�� �A	����W>��X�e�4>A4u�%"O��{u)�y��`RդH�5���ӥ"O,��h߹RQ��B/$n(A"OX���
M�uc6b��O��Q%"O�[����)
���D�ޥ��"O�+5��.V�0 `@Q��|�Pa"OBd���2v0����/&U��}��"O���@�DTb`��2!Qܴ�w"O>�Y�+�Rp(<�B��=b��pa�"O:��E�\KǺ���C�ު���"O�
�����EIB�$`�X�Q6"OɊ�����%�1�� M,cD"O��W JW/ |�B�V>S'�p#�"O���n�,�\i���G��&"O�9��j�����u�W�s�E�"O���F�ip�|��K)w��G"O��Y�S�+���cq�Ǻ���hA"Oj�x`�t�\�cu��s�*�rf"O��-������d����7	�!�D�ب�G�^���U�E�Gn!򤖿4���b��95�>��2��(b>!�[!W���1ł)��)h�n�T!��V�L�|�7o��5�<�Rrn�71_!�d�8P����>�U��δ����]P' s�(M��խx<����,'���W89V�t�*�+wtY�ȓp�(���:��H��N%l@p��-찢�M6�Bm ���-�����+����P�S�X�p8(3�^�d\vH�'�a~2-�
^Xk���B���I��yr QC�͂pGŗ(��I�n��y�nK)D:L����caP}:� ?�yrO�	Zz�=�!O	�U�lt��D�y2��"��@�@�_�?����1$4Y�(�=E��Y$2�z��R�&p���c@ D�Ćȓ,G��d��.7)ȥ	��SN����?٥����R��.*�$Th0MM��$�`�poG�a0�hV"d�m�7D�tЂkf��$z��($�A�v.7�^����'}����h�(>	�e�D���j�Q��'��z���?:
�i�dF�ilZ��)-�S��?�Ue�&p�x9��I�� �C�~h<�WdͲ�A�a�^��Y�q�%���-ʓ�H�՛c�3:1fUx1�e(��*��'J��<!���8T�D��&¢�Q��INl�<�*Km�$̩$K�:�p��p�<i�f5n��4	����АC��c�<�C ¸*����7G�`��i�J?A���<o��< �h�q |�("�724B�ɫTz492�˵g�R��w�ʒ<��C�I|��"H:�&�zp$G�F]�C䉏m��AiM�R�iW��g�C��,ٚD	#D#�Y�BD!o��C�	D+>@0a���Eb���m��B�7l&�=���"J@1�!�)?E�B�Vtt ��!�8-�8lأ`a�B�I	[�Q���<F��PU���)F�B�I�c���vf""�Ɓ�u�K�=�C�	y\L)W�ɜbH�-�jHd��C�I�G���hՈQ1V?��"H�OP�C䉝l���� �G�N2�K�E�i4�C�	�s��#i�Te�H��@#=	���p�ҪT�S4�:0Nٵ?����ȓu)[��
	~Lёu��1��L��S�? vX�����i��eK�s��Q*B"O(x���8+6����?G�0��u"O��3"��2�NpEe��#t��9�"O����cB�����a*s"O2\�6L"C(T	Je̅+���"O�E#T�À�܀s���'Z:�e��"O�TnU�9�.-A-�4)| �"O�!
U�Q&I� �pf�F&�YXp"O0|��ā�/~��	�*z���	hX���ByblAi�Q�OaR��g<D��P�C ��T��,0�����$D���g�7���CC�	�k+�18�l!D������Iʮ��I�:n��t�$D��3@�M/\���B���m����e�"D�\�v�]Vgv5��*��r=y!p�<D�hQ�m:s�8�2�d�e��qz�*'D��XԈ	�?�XK���#�-�2�$D�d�TI�$Np��2��=�p�۰N(D���Ā�h
` �Ą��2r@��tj0D�@2�+�>����	5v{>���-D�8Q��œ7J�J3ɉ3�4��f�7D���`ߐ?���Z�c�(g�&E(w6D��z��\�Y:.�bW�G����X�M0D�ȐgF@�F�!�%cD�e�AUe+D�ȁ�f�U�}y�斵���*�n*D���a߰�n�J1.�C@�ѱ��4D�ܚc���;����c�Á+�4�)�A1D�:�e�0\a�ACH�4,�3��\����1j���O�.�)��@,UJB�����P-P�h���ܥS�B��b�d�H��
(F��$h\A{�C�	�/ ����4��U��b=�C�I9�j��元�}�1h�8U,bB�Ɇ,34pړ�� �ƨb��B�0*B�	�(!�aP��Is��X`�� !�C�Ɍ ��93�g�({���b��#j��B��u�,8а���銘��. F�C��<n/Vْ"AZ�\n�iFO?2^C�I�<X����)[V@t-��5�C�I�]�ma�A�M<2� ��(?��c�\��I -Rp@�@ȐX�
��f�2"b~C�i[��T�t,�wq�u��@�
{R0C��;��1&�ĚT�C��V�`�(C�ɶE��ȀP�q���I�T�rMa	�'!,;e9&0[2�! �H��	�'�, ��Ň5H(ny�BK_q Zq��'�� ;�
��EdJ=���S�d�V�a
�'���I��� 4��x��I�2�x}R
�'ml��B9� ]���U��k�}2G�w��ħC��a��ˑZ�`���c����	f�a�I�
��M¦@L�U1�u�����?�(��	X���AB��v�<+ӎ#��B�>"�fXKg�1Az��F�ֆl|b����ɰ?� ���rM9@��1*@p��FZ�	4ў�|:�'����.�M͒c���8RvD:�'��-�����|���bm3�'�Ar�Om4���)?y�!��~��U3Jߺ������O���O:�y¦��9�>���<����.ɯ�~B�)�'Q�2����J�҈�!��)^�fy�ȓ#����ǩ�&�Y!�c��Qԥ�ȓZ�ͻ�@��O}tةcN� � ��ȓF�P�MD/���7�L$B��F~r���
��3�	#S�@�s��[�C�)� J�C�c�<= ��`�#�Kau� "O��s�-LŊ�qgB�F[� �"O�!�"�>Tk
��`U�0"O���BԦ_��F�R� -{�iTў"~n�x�(�xb�ךL�X`c�ҎV0B�I'+~��%c�"J^����Od�C��Q��=�a�FF8[&FP5`�C�ɳ%�R���ܾ%�,�	��˅k.�C�	P��Qe�Ӱ�\t���3y�B�	�Cj�q$�I�n���QӤs�
�O2�����*=J�r��yl(���HA��!�ƻ
Le���5HX�u�HȬn�!�$\�3�6u����D�$!�-��!�
�h�� -��-�0"�:5�!�^�{5�81�	%+~�;1�C��!�\������� <M�!�AP�Z1)��%�Vĉ��(���F��8�T˜�x1+䮓��,�pK:D����G��f}�볫R~�a{�8D�H����8J&0����yC�0D�`0ģ�,'䬉p��J	6���(B/D�@"�kƿ2�v!B���1*Eb�
U*D��X��Tq��Y�1h[�+�L�i�,D���$� �<�CtԹ 0���$*D���a� 4?�*p�b��"\����.#D� ֩�;b�P!
E"�Ex����=D�H��U�3<��C���8��ի�a!D��*���iT������1=&ƕ��-D��;��ۥYD@�*�L
�K�'D�����_�l�-���W���a8��2D���w"8,z#�ҟL�����e0D��zr��b2ڈ�ӎ�*h\C��.D��� ��`:J��!�;�޹%�,D�Tp1��!{�MAT� |�\Q �6D�H�t��/tWn��$B�~K ���� D��*��7��TQq�B��S6l#D�lЀ��=]Kx\���U�}�~�2V�,D�|{�'e��]��D��B"hx�)D��+ۈ`G(��L��5~Q�	y�<��nW�c���'� ���؂�@m�<Y@�ܻ*��)�Pńo�C �e�<I�\�2Y��z�����dL^�<Q5�Y�3gRL��U�q�ZA�<�����T�&tH&�ļ!l���y�<��E-9ތ��� ��	8�c�t�<���%q�A�W`PZ	B�W�<�C�>������|�ZY����O�<)�ʇ1xn`����5m�ES��L�<A��J�jy:t�(A��j���r�<Iq�."; !�(O9$|Z�Əp�<���E+̖�+�E+k�v(�)X�<�!��I����I��9��B���R�<)���~w�y�6��8C
C�<a���J�� �0i	�ō8I���y�؃z%Z���L�_��^��y�a'*F �@J
I���Q�ӌ�y�Ǎ�=����R�t|ε�aiH��yr�"|8�ٹ"I�n�\h��@��y��تFn����+D:a�R�k֏ٯ�yB�ԳC����K��d�޸x3@��y" A�
F��Y�,5P.��B�O�yB�X��	�f(fj,�6�O��yR/��vr���K�-��L��y�`�0fR��/^�F`�Å Q��y
� 86�B�c6��⨋$}��1z�"O�E�qA60XA)Rǖ��hR"OrqR
U��<����Q���#"O�͙�o��# ��Ģ��U�3"O��Q�c��5����WN2 �"O"�ᓋ��m�>���d���s"O.��� 5��	0AŶ(�J5�t"OT�E"��ꝕ)!��"Oi�B�V 3��񚲣T 7�qa�"O�t�vb�"(���/�X���"O"�����Y�VJ�O�"4�4��"OĀ��ǗAD<�-F'o�4�q�"OpCpd�80����;j�ʓ"OԕsХ�	v�8j�.C&���J"O�	2�
D<=j��8ċ> Y��I�"OH���j��
��q�1�Wl#���"O�	t�
�P�-+�����"O����Ʌ9>���emR>w"]Kb"O���+޺:�r�T�� ��ȃ�"O��i�$��7VX3`,��+�xxAt"O�����D�X�b`ѕ��0\I��"Ot}�d�D&dS�!��Y�X*z��!"OT���߲;�9��Z�Y �J�"O�ɑ䆄o�Afi�-��}C�"OM��F��.F5j���fͲ��p"O^���F+^��1e+�	����"O�e��쁵T:�u���< ���"O����B�h�l�	���
�r˅"O0<�#�^V��THA�쌳"O��|xĨ
[��i�/��3�!�Q�r��i�9\��m��oL�!�$�&"�T �ը��Rv��$ܼ}i	�'m�M#�H$"��hqvbG�7]�q�'�ޥ�󤕱e���낦�-/U���
�'Rh9��A�:����s�V�nu8��
�'>��[�F��&���(�3t��� 
�'��<���
.*w���!`�y��q	�'�8��ŧKgR����yw�a��'Jd�cu*�)ҶĲR���q��Y�'��=� �r�M!C�С3���'��<�G@�'���!�H�nI��'�|� �
�:H %���.4?�hp
�'��x	#�G�,�&�)`�Z��:�;	�'D	��D�*Ky�DN[{�*��'�`�C� X�y��X�6D� ~��	�'�8a�3& =�֬s��A��p,��'?��iU"]�!e��H�#^���''�܋�ʁ�p\�� ��l/����'Ֆ,��+/:!d��Z>�	9�'�h�i��'0�M��K�?�~�!�'1����,�(I���B�j� �'���C�ɫw�"X�V��/}��`�{B�>]m��{��Ӽ1B��A� 8",��ڬ��B����Q�1�U�O� �D��*_��`pmܵ��T�T5F��O��A�W�2�В�{�� $5��x��&AȦ\)"�Y'zݜU��kɔh�q:�J�!��e���'����g�:��*��#���T�6mAꕥ4@!��O2�9p�\._Z|I[v�L ��]A�"O�|�-��+$��GR�(` i�>��%?Y�$��Hl�雏�)�Q�>8�A�p�v؀T�J!��ԙ���{#c�&��� �&&Z��`��9470%lZw�yb�%�3扔yF�oJ�b�|���gKd��ęXQ�Q(!iԬ�Ƙ�֊.r�� 5ύ2�T�z���*l�z��`/lOr�#A�O�th2�ÈW9�!�`�ɎrG(X�p�
F�I`�ƶ`�� _�� ��
���*6�8�P��7I�ڔ'"O���%\�If&T���Ȕ-p$�Ad��.R�e����]ўh��ǁH���b��gܧ�yg�T�e�e:��#m�����#�y���4p��Q�V�Dvi��[�	�@0p{�nٵn%@Y熘9 �6t�Yw�ƍm[��'V��ւ�,�孟+^J��F%\O��1V-
�2��	�eQ*lWȐGȌ5`\��X#����h �����l[f�7Q����ǅAQ:�`�G��$F���t��9b1O��� 	�:ep|H���cq�50��^�K�p�c��ź�楟�`�2�W�L�)���4
�n�<�fH��n�[�HԽ�y�C��n�����;C�^�q�Ѵ>�΁������'nr �[�w�!"�=3d�Ms�(��Ь���'��!HfJVP��(ê�:Y�6`Q� `�b�a��7����E��>0xJםU���?��Ɓ?x�4n��.����Qz8��$�ˬ��FVA�Iȁ���C�B����+Q�`3Ù��4@�ɕ�,�z�"u |O⌚��w).��EJزd+�5��>)�+T�a�@��xa楁�*�H`Xk�3c�@ SF����u��\;na�D�_�&X�@	�5�y"�:QX�p��&K?���?B���kuE��Q�\�C�z������;R\�	�O���e�����;]��H2����-�d��1��b(<ɵ+��epF�aFh֣K
N�:��[WU�Hif��d�v�D �*D��	��Na{\��� LqOn��t�H+B�Ɯ{�a��%��	ST�'� �#�@m��׬�\�,�鐌��jr�ɗ%l��NX	Ʀ��,@� �`i�6\O�#�a�(a����P�?�j���>AQ� ptH�ժ�}� c�l�~<)2�.Y�z5�g��)
�S���J���ҝF�B��':;h\��lضv�N��c��2$�A�Cc�;ØQ���9���?2fD��\?񑅈ٌ��n݃,ۢ��t��]��h�+0���A&��G߆[��a��#�>�Ѐ�ˡJs�u��\�n3\AlIJ�n!� ��\��]�=d%�)r2�M(����34v���O���� �A�!9�����	����r���`BN�3B���O"%蟯AfV�y��� �PA��I�yy8�1<�0�����E4�'z�y�Q��!�v 2�O���Yv��1�	��W�.<��Bԥd��q��KD�4
x�9'�^�<�t���Xo�ᘒ��%�ք�e���K�5��.��q)�
Y��Ā]�[k���'So��z�ef�q�@�և0Br�FJr�BX�@�$�Z�|���䅃
��p�1���E ,X���}IZ(� �I�O$ ��:ˑ��4�C2%��Rv��e*_��μ�C�S����	�~OPb#�"UR�sPbUp����"\O�LK���
H��ðтN���6P���t�X�0镄Ò0�v�@z��z�/}rmB +�(���I� ��L ���y�4(��X���1R�I�!-��"Qwp��k	�3OpQ �
#4�m�$��*F�Q�+����:���J͢��R��D9��K�7�e���(H�	 ;�\IP�H¿V�؅�PB�*?]x��
O 8iF�x,�DJ�k�	�DK"O�h�ht�ߴI�p�I��W�dD��A��Pi�Fd�$j�'t�$�D2AC�-8�����Lp�� ��=�!0��£ʏ�Z]�ԧʈe�iB�!B��l�K��
1�<�JVg�j��H  ��9"�hcn�*`r�P��$r�����>Y�샰 ��M��	mz���N�T� dњ v`��p憚:P���p��	@�bǇ����D�\��,��C�~OEQ0O�e��/� V5D�GO�i��y����y�XC�{���H�Z�I�go��U2P���ψj��]S5�Ĳ�`��\���GC�Db⼃��'���Iw�[q�3�H��`,����`��]#=a�<�K�-�& �/���+4PU�t��h�'����]Aze F%F�������o�'���tnĬQhAh�E ����K��J�^����� b���¢f+� J�-N�Z]�fʞ�/m�����Ȣ5��X��%8����j�d���F��QOha�����R��f��j���a$�$�� �*��e���&��RIdy���O�2KHر�/�()���� V�j��dD��8��I�R \<(��Zeϼ$BUCD�,�2�Sՠ�@�AFL
�R:XL��B�PT0 ġZ�dϰ<z�C�4*�(杨k�d�B)�B��B�D�:����	� a��
[��<�B� �kM���M�
Pzx[�mҩB� �V��?9ʈ�����"�:T���nD��3S?�����	��ܰ?�4���[�Q#�Fyb����qw 38�*�{Vk�+U$�r��tP��"gH��-־�s�N�90k���e)��9pk�HK��L<���ժ-�����3Y]jL��d̪{	V��A"f ���7Aހ�� ի���b�'ʶR���#�>V>��y�蜧Iu�@�N�=<�}�掜y���B���G��9�H�7`���kݯ9<��I�0$��H �O�r��QA�Iɒ=�/Oα���7��H�H¡7\�C�'�^�H�oLt#\��QfR4e���Wl�R!�f͙�l4aƠY��r���Ulђ��I��R���D��h���닐=Q<��R#����'Uh�Q�d��=!t�r5��"|�d 1eF�VM�	ܙ�F�	�� "X��4y���Zƍѝ|��+X��0�)����qnb��ЋP�mJv��<�a�G���Ƅ��2��?��wR,���]�j���S�Zq�VL*
��� ������̊��[,!1�D�!c�SrqáL�3e��z���6�n]ޑ�$�a��Bن���b'K�`�B��%\Oh���i��[��TadS�L#���_9(��"�:$ �$��)�0@�$p��'�Z=��)����-����1��{�h؎c�y�u��H�^8(����p��J.p�20Ӆ��ȓ'`@�ĄKή%H�@[`)I�G�ZJZ��L� P葨�`�S�O�剐D=T(��P'kN�	r�N"C䉥!��0�5��4��I�C	�CVTb��_ʜ� �]'8��� ���e�'�X�3��|p$
A�|:xY�P�'Y8(:��μ��h�@kD�5�R Js��dq�4�E@�:�h ͅ�6U���v�8d`QI�2~ߖ���e��'ސ���eP�tE�-�o��z4�ם�TF�q�u���تFg��j��ڼ�y��8�R1����1@�
_��� �ӌ� Ha�EB�įR3�����)�<��H��_��PE� �0&h^I�<��8X�LpbZa���-N�gvx\�B��-}/,�$&ɟi��`CGu�'QV�֥�JF 
Q�����)
ӓ%!� ��w� �B
Y7YlA�g�L*0�����?`�L:�5��?�[�.V�(i���	��]�%�[�Dæ���ό�eӺ@ق%���D$?k���;�䳷 v�Α��i(D�X���k�ƨRI�2]F��)�)��� ��vM�%�@�5�"���|�'Fl�Ơ�x�LI�P�X42��%�	�'D1��T/�ʖ�D\)tA@T3y:H�R`o�*h�^���@�џpp��s-�I�C��A�;�j#lOt �]�`�ZqؐƂ$)�\U��*^�dAm�>0�BKu<㯌�Y���0.�?���8'��x��� �	GF �V)��z�'j�Ι����nX���� ֖��\&V傃"zF8!
1c�B5���u"U Q->8�'�"1�)��d �7G�4��ώ�,�`��@/D����W�<�R���o|&ͯ<A��BnP�9��'6ёr���/�, ��^�*���x�'vNmT�1!U�c8+n2��v"O�պ!���t��d�L^^�K�"OV�3`�.~��h�PjZ3U�}"O`7h��]�~e�F��EG�Y�S"O��35�^̆9�'됒@PB鐂"O4�cE�Y$"=�	BDNu�"Ob]j���8�tt��kr;��	"O���BM�AE���*$h9��"O�K�,¨t�E�1����W"Oڀ�teZ�E��p7hQ�(���f"O:�KF�ުrM��Ĩ��k�8��3"O��� �_	T3aɋ�+�
�x"OƁ�T�߶.�Y�։�
H���8"O�2�P�#>�3Tg0r�p�Ie"OlH�j�<=g~Y�@��?~��!1"O��8!�Q
#bDS�e�)xz���"Ob�J�]�N�8�M�wVj(Ku"O x���Y͎�{�g�
1H�"O�d�2[�0���Q���ATn ��"O4Uc ���P)<D�5/YU���"O=��O�~�@�*�n��j��`"O.���ko':(r*��X&5z�"OH��s��,K� ����+.
�X�"O�L��i�1�<i��bG���2"O��,@�t����d��>����"O �c]�K����5厷Iꜰ�U"O���d)/Hs��`��IW���"O�9z��8$kD�� d�n�G"O0�Zď#a�v��AD�[� q�"Ov�u�qv�����T��p�A�'D���T����l�P�7Aʐ��@ D�� 4燑3n���'N�C�ԣ�*#D�\;�%V�2�����Eϡ�y+V�>D��Ѡ��"���\~��"�d0D�� Lx�D�X��xd���ǫ5�H���"O��(#��y�ڍ�P�� �@�"O���u�ti�m�'�T BW"O��;�C�3!���K�G1s��kv"O���+¤ ^� 7��z*�C�"O��贊�+�LdA��Ǫ��Q�t"O]���^�oCr�+�fRd� Rs"O���pl�?;�D���
Tz�9�s"O¼�Ӧ��Y!���f4��"OV�9ңD�PF���@�>T�"Olՠ�I�u���q%�_�$E���"O�� P*C=pV�Db�i
�T8�u+�"O(h�k��D����ċW�E��x�"O�� t/X/�nyZ'if@*0J�"O��
c ՙC��"�G��AM� �"OT��ͦI�,���&קH�0��"O��
f!C2?u�XG% �c�\�*�"OB� ��b��ر���%�虰4"O^� =9��u#d3 i$�@3"O6D'(� 	����\�z� 3"O�q�$F���s���:�
sq"OP�����
d�!#P��$!S���"OlH[�Q&���-+S�A	�"OF�Xt��%~)��#�(@�"���"O@	CC���@��L��J�"%��"O��*��9$Ԍ]Z���<��"O�%g��5*ZV5��I^�(�4i�#"Oj�A)�>~�
%�ΉbS�P�""O,!D`�d��{G����ې�y��,@#�@�.�,83��R��yBh�>X��#N]�1�i�F�
��yb炡���㇃09��9x�ɔ��y([�Bcf��u̔"IhP�@M=�y�G�]���b�Z���B2N�#�y��τF� �g
ҔC��"�����y��78D��-��D'ȉk!OV��y�^' v���%H�oApi��'ڙ�y��L�kFus�&^'t������y�,�(X���P��&d� �y�N�#�y���B� M�d��]b�MŠ�yb�A;ς	��NF<;GLa��aI��yR�ŏJ�8�дOĜ�r<S�E߯�yb�Ѩ���`e�|Dvu���y�\pm��0%��s��Ȉ��C��yb�YM^
�b�B�8Z��4�S��yR��Yi����	ԋ`�Y"#D��yR��)J���;ă�ZZb������y"̑�f�h0nC8.�J��$�!�y�M�����T�Ŕ��pر��y2M�2(ި��Ѥ
�T��(-�y�,9�������������y�D�=*��8դU�pn�T���y�j�Hc ��3�U	j�٨�A�;�y�U ��9J6.l6�I��a��y�mP�6����g�/0\2�[�a��y�'R6kt~��S+	�,-t�@V�C���';~(;��E�>��?5��j��h�sh�� Tb���`<D���r�����	5�P����� V�� �>Q/p���$�b��!h�g��!.�(�ꇈt���d 1jʄ��K�6qIƨ��F0�f�)��p0�*3�Oj9�T�,i��	4DpK7�'Z,�4��o�����l`vfN�VI��`���R��$�%d7D�\2$gD9u�X8"��ġ8l#6B4}Rd��@42T��LŪO��0�� �,$��\7@������C� g C�)� ���������;���29�b�؃�>�N	bq����HG��q�c>c�:ƨ�9r�Ms�ؐz��9�;�OD��fhX��z�	a��Zʸ�5JI�pyV�֚&�\���1]� ��ą�5i6@��l��v���P�����臦�K��aU�e�󰃕
�u7��m#�H�F0̪�1�y�@�h� k$έ(t���B�̙V�K�G��bV(�2�����k��>��;�j2��V(%7�k��[}B�ȓq<pkei?Fl0�3��$���S�'´R�P�c��üP�lm������͕�W���>)��F>7i�����D4P�"M��&�z���!Q�ԿK���5���&5#��
d ��V
V+<����6�P�(��ݓn�f����!D�@$��(\ VU�Rg�v�lc�\���u�b�k� 
�4������*x`8X�H��u�C�,x@��h8�:�PAGR�y��ҝ{��Qa4i2��Jf$D�c:��(�@��{���/bJT�I fR�y��Oˊ�x#0��)Q��]g�j��1,��(�OP%x"]<6ȍkb�'6\�����=(ƹأ#;"�x�	�#T<	 ��[p�]	9=ޡ3�2��	pۚ ���ZE$l4[$�&�p<a2HƧh9����'<��q ��]�n%��A��С!��҄@{��	����3�9"�� ^��Z}2\ʷ̓e�Bp��
VC��'�t-������L��M*P�V�D�}���:��.G,be�����^�u�^h1uB14�!�R7<Hݹ��h︥ ��R��:A;0cm<R��&n�e�:U @.S�:@ѱ��Vc	��y'-��O����⇹_��5*���Px�O]&B��0�bo,h�vm���®U��a�ʊ(�H�Ҷ�%�2�"5a�A��ؒ�ůo�h�(+� �4T5�d9E�:tA㐪1OT�p���;M[RԨ�m�)A��8���F��6iԌIV�mQ��[f~t�ψj�P��^V���q���	�^�R��с#}��$/0*����=a�l��!(d�<l�b#R�<��}��F�@��1�H�2�1B�.��'0��r4(t�+J,$TɱPO��d�4Y�c�9���:2�T��2lf�˓��N˞ZS��=���4�6��G��
����L�A�3
O�����iJ��A�ӆ%��rʉu�8��d�a&Y  ,������H�oE��9q�E�H��������`4�Tu�nQ��ID�4X�`7TR��µ�)v��*�c��*$�K�� !H9��kwG +46�<@Q��> + �דX�����4:���CK�IvzզO����W>�����+�W�lh��gA�~qr����"�K(T�x(P׀�6ިm�i@�iMTP�ȓ*�p��E�!�H��'�ϵA��p�H�4hoB�b2j��y��xKDύ7,�l�F��h��'�|a���}��� ��+l����?%a�B�I�X�*�� L�u��騔!j�"�@d��	�@�k
�O�J,ڶ˓�Cy$����>r����d�$���	}9�Ph2�[̬(�H�,��xb!I5lDb��@��_��R����-�5z�^�"4h�R�„>n�b�� !�9B�.!/����'�Bt2�ʍi��r�b��+�ikJ�+����VZ�5�II�a��3F�L�J��Z�hF>��4�æJ�b����#�P� �� 6:h�ēr������1�hT2`��D�@QP��?�Dlam��+�� ���t���qO��3��DBH�G�Ve�;�b͡���F2��e�	C�"`�c��`��cb׆:��xT�
e�nāD%���M�0��J���)qL��>�����A_~����Z��t�8��-Ǯj��Y�a��b0J�>I���[�~��v��@!s���q�.RC*�OҰ�Rw��$.Ո�	�0��m���ڨr����0"R���<��˓<Y�x�O-� $�D��<٣�ވ$���bi�M��䘃��8P��0���(�:ʔ���8�$	�+�#�֯U
]�� �P�n1��'�4x;��K�r��%9�)�@�x�A��4V6���o��px��D�7�"TcU��/q��1	��GG�Tۙw�4�BX�|0Òk� іȊ� /�5�e�[�!������`M��J�d\�
k���8)n�� �D{Ӟ�Ss�c��[��̞͌H[�lI���~j����	=��YI1�̅dU��GyBE�<yz���U�9��m1�`R��c�'		 D��D(܋��a�,��a7�u�p��8O�̡@���U�J�F��'L�>��"T������|����N�+.<z���)KBx���o�=W�~t��A�#U������~��;���). ��G��-��p��Ijz@�𯙙jz`�2m�I���°��1d�X:B�	�}���SG��VJI9cf�$'�d���q-N���E�1b�X"B �~���;�bd��5�H�rM�I���g��!�BO.�O���H˿���$����� ��TՂ�ҡԦk��)�Dh��Z
��툩�VQ��o H����u��Q܌��_?]*��F&�0�H-y40y��T,p�6�Gy��:O0�H2�îv*)��t�:�[�'=C�x�P�CE<��a�J�f��e��$L��	Q�N���L<!r#�?LN`�rw�a�^��F\?"5��td�p��$y�Hoc��k�>��n4��	�5x}!��S%`�@��$'i�^,�c�!�}B�J%'F�}�ā�l�RL���Xb��x"⤛�L:���˄k��y�O�0t�`�̴Z-�D;/O�a���"���
$L�N	���'�8����$u�H��Q����UD�1V4���@�
� ��(YC؁!E̲�L��+3��� �H�/XF0�1�qDBAt�+�I� V�%Bϙ�@;�-��ӞAFx�3"5�(1��`N���H�0( \ȳ��%D7�OX胫+�3}r�E�g������њ�
d�$�i�Z$I��٭����L�K �6��S�Ͽ�'�\�1�8]��!�.bd(��ah�<�ʚ8`���υ�;�H��FS>s�����L�|�J���,�Hg8��'�HO���e��S h��A�E�\��I���'�z�J��ڰ�2P�%�޼e��$)��\����7�R�]e��K�
��>�'��gT��B�/#�fi� �I�':��G�`[1ۂ��.��'���q�瞐R�>�pS�J*/Cu�ȓ��8@/�$'�v(�b�޼{M����L�w�ty
��F�*�ݫ����b�Q6]p#���$&���׋�1�y��B@0�s�R
� C�`[/��D�9�:�8qM@��55@f�'�����̛8��4pBP�0ê$��@���"`S4?˦!e��1+�����"t�܈��M�Q 4���(j�z�R��5 �h�v�ۢ�<��
�n�`������#�`'?Pk1=����ELY>@����1F5D��'G��S8E�-��,�]ɤ(qv�$r�!��4��MP�<E���Q˾ȡ�Z�,��� "��`�ȓubt���\�~I���W���K�'�!�u�VC���1�/O���OEqT�D6 $DC�<N����b�'�0	�sF�:G^��S��+�2�Qa��6�>�'G�?�6Ъ
�MVv��n�>�Z�Y�aY!!Gy2⑳N_`����oM�Za&9���NuԖ*p{,�cB��,�l��'�� Z��]�70>ɱOJ�"$2��­�"�̭"�����1R2O?��Ի]�<i�L�(~'�ZG��7o!�ǘ:gLi��(O)��zA�CKx�ɦ����l�,s�1��'�3����U�V Y�<�u�ق\¸Ȅ�I3��m�攑,e3e	ή4p�zr�)uO��h�A�6�xb���UҤ�w��WM��A#�?�hO�±�5*�����IO�m���
���p1B��ĉp:!�'ܑ����-l����f	����9_�@��毙}�)�'V�xt)	�,b	���2H�V}@͆ȓ�T��v��o��X;��7Y �@�O��VF��o��y�,�1p٠r�,Ida���%�[ �y�O{�bݙ�Mݸ�}Z�DZ��y�O�|5$82!H�&r����c�yB�_3F��wq��!#Hԫ�y���K<���oɩm=��0d"�ybʢm��T+'�$g�����y��y�ܢa�ވH�v��n��y�M�ݔ����\L����Ҳ�ybd��H��Y7�9B��$٢L���y2 ��6���F-�=0)T��CB*�y"�B�i�S,:~Ipt:��X!�y�e̛a�*��LU���5�EI�y2/�:��C ���N8�&"�;�y���@%H�#��^�'f;3���yb�wF((8��Ԋ���͐%�y��		-��B�B��	������y�,:'�0�p%<�@(�kJ�y"��<�D@wJ�����J�%�yr��&o�-a�KY�Me[C��y�#��\�q��M-Vn���,Ƴ�yb������TCK!@D����o�y2�]�Y��|z ��>B>��Bb¢�y���Ӓ�!�%9g�ى�bվnA���ȓT�&��.K�~�V�	5�'I����s-d%��FI76�0A)f��)����Fh4 �I�+�ȍ�W���ޔ�ȓ(悙3��I1O?���&�J�A�V��|��Ƞ�E+iR�|��E3X�DՄ�i ��<�)���-t�> �ȓ;��#s�D0b)z5A"�;���ȓ ���z4������{�v��S�? �%9P���)\�ib�"�=I���T"OJ�����31|��'A�AE��h&��*�y�g�ަ%� �Ⱦ̆��M$?�ۖMF�b����?��0������#F�	|_��� ,L#)�(	��QޱZ@ϗ6X�2��6�Z7��V
�����C�v�է�O�"�#l@}��o�Dg�a�tǏ�VM:�&��M�T\Hd�^F����&�%�6�!a�ڕjͣd�&\q��h"�OTI���ꨓ��E�2&�\��PB�Lذ�.�D�!�!��ӵO0��u�� f����퀥O��X�O�!CᛁK�ZAE��iv- g�!N:�a��dX?{�� ��Ou��,�&���KŖ�"}���#�e:�.):��p������Kf�Y!LG�A*UG�<Q���}g�y���K�#��|�g�; �*��gfاL���'�4������xu��%+��;W[�z��i`.���D�9Z�h��V>��)�*{���wI\CS��C � 1��>����9��	C:�U��c�+1D�ޤ� J�=��
�˟K���	����N* �X�D�D�Ы	@��Q���%��y3�'��Dɝ5��Xo=}J|&�֝f�HKE�1���1	� P� �i�!�4T�~OE�O��'����!��Mr0A�=L+`�S%Ҕd6��d~r�
$)�n�O>i��	ΝP�\ ƄT�5'��#$�2}�I)jLT�Wh>��	 /���;O9�⠀ƵA���'��}�P�51OQ>�$Gv|�	[�'��QӐe����Op�i�'�0%}1OQ?�0���z|Ȝ�e��e��ŉį^�C[8��,��~>-���ԟ�qJ0�E�$КEK�@׹z��@!'r�t?	f&�(��Y���u��E
S(<xDC_� �r�����~R�'�0 �ܬP�ڡG���'U3u�"��܃m>��ӳ��>U�u� ��!�m?��ۣ���T�,Oq�<i����Hݢ�L|�Y��dW�~�Q�{��D�\��V��2KH�V�jD�0c�9�y��;5�N�d��C]����
'�yB�#[��!��H�/NP��W��+�yb$ź0�l�g*�)(rD�b6f��y2�E�+nP�!�:4�2b�����yg��J��I)��80r>�pT�P��y���m*��8pFW
"-�A�����y�~ PbU�	8��mA�(�y���6�ɻ��7���33È�yZ?{��DC%�T#��a��=�yEBE�ڸC��������y�,�<d��E9w#�
�@�qKC�yRJѪ`�����`L�B�AYq�@�y�L�>=A�T��8����0���y�J	���wU� ������
��y2�ێ2Ո�$MÒj�n Q�! �y�j�3z$��aЗ[�^1)�C՟�yb`B�od���T��=O�|�2E�R�y"H(��Y����>�F b��7�yl�uR�`!+O�=��$:�]��yR�C�'F<��bԁ��yQ3(ͫ�y"��x@�dhV6��s���y�(�9C�T�@�m�-}��)����y�o	V|+b��3 �x��!���yb��!s�x��V��&e�*�Q�B,�yª:}Tp�����j�!2�)L�yB	]�T�	5�iv�h�J_6�y�)��/-J��'N/�|@�ϗ��y�N��4�he3�[�g�|i`lٹ�yBmà�^�p��u�z�)���yRP�h��	����m�0ظ��Z��y�DȄkHXI	�_&V�H$a�ٜ�y���)>���m�y��2�y��Ѕr�����6yO����yr,�}Ƃ�q5J�BniB.8��'j�x�B���e	��U$��[�'ϊ(*`��'�������#F� ���'W��Han��9�.�:O�f���8�'B�ِ��'@�2���#ѭd4������ ��(c�;F(Q���;d��S�*O��".ߢ�`9։qOH8�':�p��KR9q�@yQ��F!;I�!r�'��i��a
,2�5Z����5q&8��'we9abL�	'&�(2��h�'"8	WÏ~["��H   �(k�'[�������#���4l"�ܑ�'Ǵ�a0�\?~����KS,a  ��'�h��¦�i\���𢖭R
 k�'���i�䘗�V����I�_)pqZ�'Sl��Ъ8�H�I�eW&��'<P@0$�T�'�ڨ2��(�'�ޕ�v�]<es.}��IV�)l��'���p�]8cN8u��kR�q��b�'5���.]&a�A��P"dX�)
�'�����G�L]2Q�u"3�4j	�'�v)DkF%�*!Z�E��Q���;
�'s�|�go��k�����o�Nd:�
�'-p�ABXY��0/ZQP	�'D�a1t��+#�6\0���`щ�'Ĩ��v�މz,Fy�	�=L@�l�'���7�T�j`-�����Z��
�'�R�!���8t|͹��T�ʥ�	�'�N]��L"�D �vH�9uhb�	�'��3q��=;���+�,�.h�$x�'����գ&9�9Q���j����'�F5�
�ϒ���@\`�B�$�\�<i��V&ѐ=B��=����R��D�<16n��o�N�f@=�ez�H�X�<ɒ�^�q|8�"@�a)�Z�C�W�<i����n"�l�Uj����}�0�RU�<��C^�;
��B ��9g�r�#��HQ�<y���D�uq�H�2<�\�5	�O�<��+�(V#~X��m�P��5a��c�<6��Snhq��L(��|'��[�<)1���l
���� �ލA�F�k�<9��Ύ=��(#!ŏ�a��ٲ怑_�<�A����up�J��c)ȥ��o�<1!�G)<G���Ԏ68�2�B��E�<Aro]�yV��`��y�6	���@�<��-́'Ų�C�ݖq�l�"�,�x�<1B,�AC����i�\��x�!a�}�<q��=$$Pc�_:g@�I�	�{�<I��#UӒ-�ju�B��q�<��f���� �ߏ'�+�F*�!�P0\���{��w��H�"K�!�ĥR� �&��u�t)�/��!�� �a5J��tXD�R%�9�!򄒌#KjLh�CN?3@�aa�ݚ+!�D��p{����C%P�03Dܠ&�!�D��G����"[��I+��!���+_��a
���]!������n�!��-F�MbG-0`#�&=�!��\�5�h	��A	���`��/9~!�d�9;OPU��ֲY�b-	"�!�
�WnyW`�6�2Ip��{!��G�9�Ƀ�m�&,�#��H!�D0)��JA��<8����P�! H!�Q�0��Y�e@JZ���Q �8qE!�D�}�X�H�/N�DE�n�!�D��@y��y�S�x��jV�#;�!�O`�h�s��N�k�P$Ƀ�Ĭi�' ʉ���� 7���;�F<l+j-�	�'-XA률�`+"��fH�r&1���� <)!aO�'k.�H�kT�V老�f"Ol�����0������ ��t�`"O|ĩ��
!�0��E�;k҂d@�"O�T�a��s���X���(�A"ON��E�� k�\�
 �3V��bT"O:Y�Pcڂ5I*a�F���2l�S"O∈���#?A0,2�!�Ar\�ig"O\=@���WM��	��Q
p<� "O(K������q�ۯ}` j�"O��QH_9|�,x �Jļ:�"O�;�ûV�jQ�u�إ��]y!"O��C�3r%�y�@}��("O�ہĔ8`? �[���nx�K�"O�L��,�(2¶�[Aa_��P"O����k�nu��F41��Ҁ"O�p !#�8g�&�s$�K� ���"O�x���7#{H��4ė� T|A��"O�8�e�aG Y�䎛*^�$+"O��t ݤD@�k��?R�=Z"O�tg��7� ���L��{H�qb"O�ɇ|V|U��W'8��Q�"O�蠱�ޮ66��
�_Ю�7"On�WJ��S���Z�	�1~����"O
<��)ЕQ~D�1隷~|���"O܈�� R#	<��ɑ)[�e��"OD�����7�h�v���3L��3"O
��Ɖ0b� ��[���p�"O��R��P*3��Ai6���!�"O��#d�� 4�<�JI�4�t "ONe��S����)��%���"O�L�B�P9uCX"���j��Č�!�Y\�D,��>l|ʲk�T�!��� �$��2JVQ��*"O!�T�j�
�eITAK��� y~��?D����PZ�$�3��E��H'�;D�D��)B&�T�11hG2={�����:D�t0�#��V���w=�����6D��#��#a������/Ƙ�d�6D��1�@�+E&�`3q� f�@I#'4D�p�uA�t���$D,Y��1D�V[�h��M����?���-�6�y��!Ot� V��G��Qz����y�c}��@g�܃F.9��G��yb"ƾ��Sb <?��8s�k��yr�]�g�PL�A Ԑ+@��
7�y�� ��LyF��uw�b��S!�y��ڞ>o�	�"4p��)w#X��y���i�AT�i�\$�%M�y���%��8�&�&^JHхjP��y�$���3���E*�Ѹ�Ο-�y��P�'皬�f#�
+������y�m�2s�����'����+��y�I4�l�Zg�
�%��|�E䚞�y�ߢh�A��FC
�p�ґD���y�@�!Vpظ��m��͂C@�"
!�YdZ&*u�)j)��(t�ظ}�!��|�2�V�ٽ!��$  �_�d�!���L���a��@�,��ʟ=�!�� * N��$�U')�>Dc�k�0X�!�È?W@uR��;Äu��h�In!�DB&s���S&$Q�w�]�aN!��0�j���2k���Q�o1!�ėu8\dpG�D�-�Y$�?^�!�$��Y��x��,?P`t�F�ؼ �!�� �xYq!�=�P�aF�'`	9r"O�4�?}c8�*'���.z!��"O�8����,l��(e\�
�<��"ONqۂ�ʉM�ղ��/����"OTS��IJ�D�Ђ����&�`"ONM�#+Y�7�2`����O�̸xV"Ol�x�hTD�$`*��Q>%Y�"O��@T�Y{^!h&bN�EgZ�`V"O�(F���[ �"hC9TH��BG"O�(����6�^0��F�*Jj)C�"O ��p�R�	�ޭ�6�ݷg�T2"O�C��gs�=�Ck5i�qr�"O�4J���(�H�Jg��;j( ���"Ov��Ոߺo�@ԋe�^{܁�4"O�s����f�P�RnD`�"O��)���[���R�4����"O,D�@Cޖ[�5�0oK�c�1�"O,qH�3^�A�N����"Oj$HI�Zf�zC-��b�Z��5"Oz��e�D�G�@5�Q��-��$�e"O|Yy�ċ�a�����a�M�}R�"OdM8"�G�^D��1�z�H��E"O�Q(�BD�S�	�ԎQ�D�Z<��"O��K"߻\�	 � &�16"O�y���3L��+�,,
�fl�"O^�0"�K�_�&-҇n�/9�.�Z�"Ode�D�D8wz�j�M�'�Mґ*Or�b�kN�$�.�#�Mm�N�
�'��Wa��l���ERl'p��'�TyT$�=ԨTц�ʖfآ5��'.~,1   ���     �  Z  f   .+  k6  A  �I  �U  �`  	g  ]m  �s  �y  <�  ��  ��  �  I�  ��  ϥ  �  T�  ��  پ  �  ��  i�  ��  ��  6�  ��  ��  �  �  � � < �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�	#��$x�R3e 	F�
�Z�Bړjaӕ"O�1RV�GF��УD1�HАa��E�Oԉ�
�]�|5����n��u��'6���½`���!�Ϸ\�~Aۓθ'��I��ܩy>TD�QD��@�0L�
�'#p1��sR��i��̖"n��P�}��)��v���s�_)�y`7Dϛ !���d2��C�(v��S�	/�	r�Q�"|2�M��&U���Y��dy:AD\|�<	#�'�@d�AIڣ��w�<�kc~H"vm&#���硓v�'#Q?u�B.��Z���f��|�  gN:D���RM��C�Ze���H!Z�\h��N,D�li���Mn��!�G�o68�	�)D�@���u\���a�+4�^�˕���M;���>YW�O~�>7�5?�O�eʅʥ,��@��؋�)XP<���t(�X�6f�R��H��9V�N�P,O����+�H�s�&GOCХf˜�
+a}2�>����08B�iZr����F�<��4;�1�L�"\��^D�<IsaA�B�@,�b$�9ۨ��#�D�<�U�\dppR7� SPel�V?9���S	=��H3s�i���6m��<btB�)� ���e�+�h=��M�G��	�'"O \{��G�%��iP��X�7�|%��"O�X@�����i���e�8�"O,\psΛ�L�nE����84% 	��"O��h��A5� ����P��×"Op�qW'՞/�.%�r��V嬰��*lOV�C�̍*x=�a`d -<����;O�=E�t��N��P��hҧf+`e!����y2*�)*�e�fI�[	�T��e���y��,k�,�Q��D+�t�Rp���y�Ȑ(����O���"0���yªA�/����$O*(��`�F��y�!��@�X�r��Tr&�߭�y��Q�.u����! �ö'��yrA�[`͹s`�2d��� �j��yB�>fd$0e��K?X���(��O�#~:�!Q�?��"CO$//b�b\p�<ن���P��a�4��8��KӁUl�<Y&IWX��5�W�/��c� Dl8�lGz�+۟[~��S/��Le�&,ٞ��'���'�>4r��1K�dR���T�
�'}ܹh�k��l\d�eB�?EF�b�m�g�<i��1"VlՋ��Z�=ѐI�ң`�<�ue�9��A��+ Х�"ˌZ�<�V��)�U �K'}�fi�bˀmyr�)ʧh��A����ÂED3B����n��@��;h&��q䐦K���ȓ^��\{�o�%Y���3�I�Qh��ȓ7�.�z��A��^���j@Wz�1��.�����6MY�
��P`ԭ��|�9�-��N�|p��M�Ԃ���.�@���A44���SdgȢ����=PuhW��	]r�:�(��B\l���@��Y�ť�qVLEC�_�b���6�Piӑ�ͣ&�B��a2�0=��n 	Zw ς����Z�}�X���lQ�PRj�:��<��"� ^�zńȓwb�A��FX&hF��Ak��I����W�đ�b��Z���aa�%-tH�ȓk�T�kǨǟS�4xq�G�
_lB�����S��6-��gې���WjH¤ku��.3�!��΢?Ҕ���)�dhp�)��,lazb�$T'=�帀�ضr��(Ǯ��<h!�D�_�lqP��(_H.i���_�DC!�E�r��LtoJp/6�[0,R�+�!�$И�@-��" k��1r()�!���*�8��IN5Zw�́2H�, 6!��J��,�#��Q�G}ԑ���ӞK �1O��ג}2�P��J��`�K����<���$�gY`�S�F�f�����!G�i0!�@�vS�}1����F �̱�a�i�!�Ay�tĉ1Tx�X�r�Ǌ�;�!�D�9'傈@�LC v��ܰ0f	�7�!���>�H�25�=>HH�'��!�$6����WL��D8L�*�$��K�1O�	�����Y�hJ�"dMj�S��I��p�C4D���b&�XR��fc�t�3A>D��I�S`�phF���j���bv�<D�(�7f�,H�v�1`⚅<��@w�:D��:@�"!��� ��'otq�>q���өLz�
�)ߚn ��U�q�C�ɶ|	�pP���R*Q%̒�TR�'�ИDyZ��'d����^�mBf�	1�I�,�hٸ
��~2���2j�q慗�
��b��y
� ��;��B-A;r��7Be>�-�p�����'(�S&\A��a��)�^��D ��^��B�"����%7�����O2�=�gÃ�&�,Ӂшv(r-(�	��y�(�Y���(��g�mJ�ǁ�yb�84��ѳG��4�b�PԮ��0<��d�kH���Eh��U_N�b`E0o�1O���$�&(�v��2�ϧ�z4s��\='�!�$�-n/�y�6����(E�m�!���%���Q�,˦��l
�n�Rn�� ����Ƌ�h�� dZ�M<~����ǪE!�Рw��Ҧ�(>ܫ�V�4[�1�D�a}���OB4�@���x�������0H��8gO�P� (�1}|�lk�@`At��`�4�$/�O�a���[7r1���MAppp�'�F��O6WȤ	3�����S������'@�L1b����cw���:��0Ox5*��Z8p0o�#0H�ZE�'p�'�~��r� �ct��@`NNCrXPxak�<�����. FfЃ4�<����TG��n�$:�$�i���OW>ͨc>�������x"��!�!I�	:��=1@��;(�(�����.f-A,�y��<ə'rZU0H>�'9�M K��r!Ď�eA��x���&O����$LO�=�H��[�	��h^�z��W�U~���$=ꓤ�	O̧ZղhZ���Cf���H�,B���H�I��Mㅨ�$)/��:���~]X��-t�<Ap��5x�j�����"
��j�m�'$ўʧ<h�s'ca% U(�d��m�h�<��K�8Z��� ��T��|����d�<10�W�o(:bŚ�.�H����V�<�G�Е[n<�b���+4`b���LX�<��
g�(z욫����i�W�<)U	��T)�X�/�0�Ub3��P�<���@�5�l�RM�r��R���T�<q�����R�GQ�(}xt���Y�<Yd ̧J���/�\���[g�JW�<�$��SuV�� ��H:�A�hI�<�&K\ {�P�q'�LJ��!v#�D�<��G�V��� p�ٱ<���3�%z�<yV�A�1�J��VJF(=�f� ��^�<)��=,<yp�%����Z�<��^.H�T���9kŎ�#��3T�Hh��;�D`r�,Z�R&�E� C-D���p'*a&��kX�|���D(D��8d��8q(zD Q�6�H��H%D���u �|�Bt�	!&ڨ1U�!D�����)lm��H�C�	r|��Ȅ<D��j#X�J7��� R�.-D�h�GY�)� ��R�_w"J��'D��HD� 3"�+��[s����*D��bÂ��Nj �+r+=r��{�)D��s��� ���w�� �@"D��1�!@]5�w�0����;B�IIô�A���r�`P����F��C�	�0�Ń��\�x����ӏ8H�C䉢1k�$��)�<92ݰ$I f��B�	�� �"Q�Q�����ZIRB�	=@�V\A���2xI�9$� 2 B�	�K�5z���/�h�uSl:�B�I2_��qa��&�b�h�Dևs�B�I�a�N�R��I�6)+�,�,�C�"M^a �#�0S��lVmGs�B�I�!�F���-׿S����bH�(4�ZB�I�=Π��+�5��u�ƨ��zB�)� p�0(�gV�	�c��_<�;0"O:�6��yK5�N�j����"O�������Y��v�R��H�r"O��J����Ŷ�f��a"O �j��nS��#G�L�i��'��'>"�'�b�'|��'���'��Ż�+�{��!�`D5Jp�){s�'���'9B�'�r�'�"�'E�'��4K���K�*�a���|����'���'/��'g��'GB�'�r�'�R8:@��W0�a�bνkH�Is��'�"�'sR�'x�'L��'*��'�b={a����}�!�r/��"�'�r�'z2�'3R�'���'^��'목{W,Фw0�T+!,���B�'���',��'I��'/��'B��'��]�!)�mD�=���#C�){3�'���'��'��',��'K��'�>\H��m�]�d�X�����'��'}��'w��'{�'��'�Ρ�`�Ϫv��A�.y�@1�Q�'Y��'�R�'r��'���'���'W~i���t��ŭ�>3V$�q��'Q��'�2�'.B�'��'\2�'_�8���5rd�����sd&�i��'12�'��'�B�'(��'nR�'?���An5Vv����S.tV�S��'�R�'#��'���'��'"�'����P�u*�ZA�ͷ?er����'!r�'��'9B�'���m�J���OƽA��%B �)��³fQ�)ǝ[y��'��)�3?Q��i���eM	�w�8� �ŉ{��d�m�,��$�צ�?�g?��4CV�x�@�)Ri1��;��2��i:�m�=�X��OB���ȀFQ)O?E��D_?嚼	�J܋^��F	9�˟�'��>! 1��?������9Cz����U�M��']̓��O`�7=�`pSBZ�{�@�"��)=�J�d@ƟoZ�<�*O�O�f``�T*�y�@�y1���6�� � ���F��y�B���5%�	/{�=D{�O
"���P����0>pʄ��y"^�($�Cش�~��<��E�[/�|���ED�IJ��Z���'�z��?ش�y�[���pc��@��EKʢhz�z�L4?���L����ģ-����h��?��8u��
�+�6)/�uӁ����<�S��y҂̉C��x�AfWb�8:5�\��y�kӨ��f����ش�����ЩK2tTY�鎃T@�t��NԵ�~��'v�V�'�B��CЩ���ɟ&:r���	!J��P��J��y���X�I ΰ�!�3�"���B"]�Z%9DcnHؐ��WSD�rt-R�]����/��Ѱo�/#fLyj��G�~S*yR-�.(�!�7f�|��E;�L������(O�4�T���<�t�&)�ue.���d�!M��pc�"�a�
|�gZ�LrT�< �챧(�aM~ �ag�/Q�^(@�
N�l��qY�L
1&֡*m�*��h���#ڌ@����,Ď�2E�@�D�cN;28�j�n�6箼 Q���e�>]���1NA,@"�Xi��L>m��#��M;���?�����'�?A�_�ފ,��Bڜn��y䄈n�	���*U����$���b��R�(/\M��NH�,�2�	3#��OG���2.��7��O����O������O<�$�`1R�+�1:&1�TAM��mڕV�a�	d�i>a%?��I2F)ը0�Ӹ&D�P�E�8Ej(�ߴ�?Y���?�i�9��&�'��'�"��u�kEg|�ؓFFX�	�)Ȱ�ס�MS����H���?�����D�	g����vMԡ��I����4�?a$NF9���'�B�'�@�~��'φ�s`�!Q2`�0��*�� �Or�8C9O����O��D�O��D�O
�$ M��C)տG�6�	��	�Ku:�+kP���۟�	ߟL*��"˓�?)1n�W�d�B��� q��������'?��'cR�')員�h(�4W�LL���1<�&�c&�&!�9��ij"�'��'�RY�d�I�Xp��.� ���rm>D1�O�b�޴�?	���?����� �*�4�?q� ]`�З����M�P�)��ia�'!R^����
t��9ON�Ƀk�49C��Y��yS,s|7��O��D�O���ŗ4ظdn�ß�	��)Mψ��/^�7P��N�t* �A�4�?�-Ox�$��$�'8�i>7��,�rD�kE?`�6LV�%5����'��"n�7�O���O4�	��B�$ /.�>���
,,,��DB�`��'���Q�?�2�'�i>����@�ųX}J�`C��(�h}P�i�A��o�B�d�O��d�$�	�O\�d�ODr����V�~@�%�E �X�	�$�	��d�ϟ��I˟8��b>�$?!��	;��u�� G��$(��j �$�����4�?���?�*�c���'o��'�r��u����\3QG
�����c���M����_!:v�?M���4��`1J7
Z�2�Rm�'����}�۴�?I�&��Q��f�'���'�2��~��'�h�"Eĕ,D��dѳ�
) �]��OHe�5OJ���O���OҒ��`�ܯf滋z0%S7� 2AN� 2Y>�n�����џ�����	�<��p(�!@?��0�ݩX��E���<��?A���?����?)��j|y�ǽi�8���׿]�v�dJȍb:e���wӰ�D�O��D�Ox��<1�x����+��X�B��C(˴I4tb@��u��9i����ʟ,�t�0G'��m��ПP3�	0����r#��a�^ �T�Ų�M���?������O����?�v�$����0M
7����2f��,��5�fӐ�d�O����O|Y�paGĦ���ڟ���?��c]cR��F��:F����� @,�M������O>`�>����<��� �,Zwg]�k�֨�Ń	x,!�i�b�'�"9�La�*�D�O��d��b���O(�	C�� �b��C/�>/��iC��C}�'�x��f�'Oɧ�d�~r��~ДY��	�y��@�K������[��M����?�����g�$�l�zQ�sM¸s��9*#(�:Ul�94f�#<E�T�'�(�xs���{���:֬�6tP���
����O����*���'�0�I���0���zTᚬdZ��CIC�%00`�>)'�D̓�?���?�s�H6M�2hۥhT�h�X!�B�yכ��'��Q�2o-�d�ON�d:���p�R�M�}Š�#V���	t�0S[��y%<�I۟@����H�'�*�2�d��.�e�8x�b#�HFOd���OВOf�t7�]�5�������$&�Pg��aA��d̓�?����?�(Oz������|�� ��IF$
��Р���k}��'yҗ|�^��� >Y��5\�XȦBY�hPx�Y�m�}��'��'��0.�J�O|2D�K:<�}��no�D��1G�%⛆�'�'J�ɸ+A�b�(�7È����s�uAE"ҳn��7m�O,��<R�W�mE�O ��O� k&�P�W�3 �!�p/;�<i�[T���	�>:t����%`�-�,�0���W��S񈘰�M3�[?��	�?)P�O<�@AҘ=�<,*CD+�y`�i)�ɍJL&"<�~:�ԨPy���ףd�\r�.��uHg��3�M;���?����:��$ШCX!&AI��<]X�酉���m��<  "<E���'� �6e�������ܰ3׎k�\���O����M�J|�>����~�;9��!�ơ��i��P`o���'h"�)�yR�',��'�伉@���4�B#��ld�U�%HgӀ��Z_�)'���˟p'�֘�Ȥy��0~�6���b��;�R�<���?!������J$�ŭ\�2��+ �ib�a�	�4��E�Ipybf��-��!KA�W)HY���3Γ�[�l@��yR�'���'u��j�pU��OA�t��� M�4xt Y�s�N�C�O���O�O �I��'
8��	�X`���aG+(�ٯO����O���<�g��HQ�Oxf�R�kӯ7���`���F��%	��{�v�$<���<�.�]�\��a�MH�P��p�k�-���o��@�Iyy敳_&6�n����aB�ǂ��٘c�	gऀ��[�IyrLݻ�O��	�D�!��Pi���/�(
�6��<�&���&�~z���Y�Pp��E]��%��%V�^m�� kӐ�7�� Fx��d�ՈY��\�K	>=����ԅ?�M���ٛ&�'8��'���N;��O�zť<F]��"���1OL�1�@�Ӧ�{�.�S�O��ޚ{�4�JB�M&p̆5�-i�67�O*���Ohp+�-	f��?I�'��YbIB�51�Q�Ճ��>XJ�S�}��ڝ��'IB�'��gI�e	��aT/��Ybya�ه�.7�O"p� !�l��?�M>�1f��;qŞ�j��:�*��dR�'# 髍y"�'��'��ɮB���Q$@�~e���]3�z @@��*��'���|�\�h����radD9�M^&6�x���vt&c��	���	Ty������S�(nJ�`Sْz���Յ��^:hO*��/���<��I�m}H2/0���K��W
 �������OJ���O�ʓf��Us�����L�l����$C9fg� ��߸t^�7��O��Ĭ<�*O,�#�?�3͖��d.�S��<)�mo���,��@y���a�`��������%
A !�4uR�mO5}�����F��%�'z剭  2�g~��M+R��Z�H����H8�ӡh�%�'j���ӊp�O���O����E��N�� .0Z�(�?R�	n�vy���{P�O�x"�X�Q�֩��@π5d�d��i���M;a�99ћ6�'���'���K:�D�O���5�P�8�4�X���������զ	� i�F��|�<���P�Vѱ�J�0L�����@<T�x%���i���'\�$Y5c9PO����O2�D�*ey�9ʇWD8�@qI�I�,��>!��
��?����?���?Q��Drxy���@С��\X�)��i�R&N�=�0O0���O8�Ok씐qS�ub2%�=g�&�@$c�D�I(�p5'������<�IbyrȄHђ�IЈ]�M�����O4.��A9�$�Oh�$'��<��E�S~D{��9o:��cA�`�j��<���?����d�1�R��'x��xq��=;�҄	"BW�
���'9��'��'8�<%�4�o`}r��ҪS��КPc�oB�'�b�'�Z����ר��'Z�(�:��M-(�4d�m.2�Z�iG��|�R�dv�8������C�)HT�	r��@ܴ�?9���$͡:�,&>U�I�?�B4�����1 AS�XhX���B�����D�{W��S�~�,b�h���]2 �1Gz��ٴ�?Q�m	ޥS�i��W>������Nb���[t/v��L��d	=1�V\�Cv�;�S�u��3.��H؀|�b�ߥy�ylZ);ص�4�?����?I��2C�'��,/n��� ���*Νx�*R\~6���"|��w�� ����얊G���wHyZ��i��'�⡊�e�DO����Od����
���B)��E���^*<c�P���&�I���	ƟP*��X������I�+�M�
����x�'�B�|Zcˮu{���z��G�����[�O�Zp���O2���O�ʓX@�,�2#�[n
�z�.D%\�kS�H0�'#��'��'"�I�T��-*a��2�DYa�@�t>'�7��<�I�(�'�̭��.|>A���ϲ)����@D�O u���>����?yK>�.O !B�Y� 1�(�>bx�xt'ēV҈�aű>	���?��������"�>�$>1�Ǡ 6J��	�RZh0ಎH��M#������_��OH0�U���Buء�/�4@�xG�i���'U�I�K}1H|�����T@C3
	z!c�ҶO P�q�Z2W��'��I��8#<�O��D�p�H�`I�5��j�FXa�4��D�`d�ql����O��	�G~5j0����NF<�ť�5�6�n�uy�*��O��<R��G�x��(U�NQ{Ѹi%~,�@�p�&�d�OX�$��8&���Is�Q�C_c���� +ޑqS(Dj۴cļ�Fx��I�O�U��-:PԚ��E$�0[d�Ԧ-�Iʟ��I�k�R8�J<���?��%k�њ6'��bsJ�z��U~HhȠ���1O���OJ�Dڜaf�#D�2�l�毜�D��o����)�AB.���?����?!/OkC#�|4���4wu���2C���7h�1O
��O����<C����P�m[ˮ �Y\��`#dO2�ē�?����?Y(O`���O���1��0z ��7��,\�؊G΋:1O\��O�$�<IҊ�M,�	JI�@]sA�X(S�Vpk0����Iʟ�Iǟ �'(b�'*�@��<�Η;B��(@^�T�tZ�P�Iß���ey`����B���B��F3�AEc_�7�zzT�KߦI�IF�Wy����'f`�3 �*�R�l��2/�%��4�?����S?0<`�%>Q�	�?!��D�;e���$�F�^����2�W����?	��wGEGx���PS­ؠ�تK�);J�1�d�iK�	�	RJڴd��S̟@����$گ.��Us���/&��X��P�q���'O k�|��d��1�d��%T�KN��z��@��M+��h>���'�"�'����'��O`�i!�μB؉EM�etxp��릙�f�A��<&�"|�� ��y�#����(AG�-	,Z�&�i���'ib�Q�$/�c���O?��K&� -����b�xddO��u%��办�ħ�?���?��YM�A�3l�p��	�N�K_���'M�|���?�	˟ $�֘�T�11�͐��Iic�>'��7UR=͓����O|�+��I�]*�+ (X���c�Ϡt�ꜹF��{�ޟP�I��ޟT�I��j�͟:H���+ΝG��8bB �ܟL�����'#ZH3Ѝh>]�e�*nf�1�##i����%�>Y��?qL>Q���?I��J�<�2�a<vy3Ҏ�8輊���)K>��П����\�'� [�	 ��|�h%��)��f��y�%�E�0*�}lZ�� &�T�	�������O������5L�T)BshF�$#b�Q��i(��'i�ɞ-�J�{K|z���B�&��9���*�1x�H�q6B(1�'���'�eA&�'�ɧ��عg$0����T��s��!Da��\��c4ʙ&�M+V?����?���O���o�4�����ܠ~�|�6�i���'9����'�ɧ�O��){PiT�%��U�S暷>�����4@α���ii��'&��O.�OB���L�����Y/P����J���Lo8�=�	c�)�'�?�'n��G��р�©A�xh��9��V�'R�'�p{�7�D�O��d����.�H&D0b�8[9���a�ޓOdH�Tb�C��ɟ������B��
}��5� b/˪e�B�Mk���0�ԕx��'@B�|Zc��]r�ט$���[A���L0�O�|�c�Op��?����?�)O�x�2L�X�Z�����o!�(���S��\'�P�I���%�T�	����t��\��k��Fz�\m��@�(����qy��'v��'��ɣ Y���OD�CŦ.���vl��"p�O8���O\�O:���O�Ŋ壟�A4��5Ę0A�ωv�f�P�ζ>���?Q������l�%>U����:vXC��jx(�z�B��MS����?Y��������I�P����M(�| ��B�z(���6(��r�!�����n�M��~��y���`��D1������#�y�,��L����؞-�:�
!��@$k�ⓤy�r�If�
��fD�"�F�(79:ǭ��rZ�����@	7�+3�V9`@�;'B�_�괰�&�E��$�]�u�ԠM�e�d�C�
�O��tB�Y�G��;��E'0��ՋN�NB��i���R�)#���6�P�e#�j��6��~��� e�̨	�۟��I�L���u�a�:c����I^�H������lrZ-[�k
�*7���G a�r�#�˦��a#�,:R���*" �IR�\%4�Òd�U�1 pʥ@��]9/H�>1mZ�'��I�9�j\ZC�V%[���C׀�;*�L�Ii~���?ͧ�hOJ�Q�� P2�Z ���a!7g!�dݣ b$��JY�=2�mX���:J�I�HO�I�O*�S�? 4��NLG ,��G��$��[7�TT�H�X�`�Oz���Ol�Ժ���?��On���! [A�x�;-�;f��mQ)nh�i��Y�nɱR���џ��6� ?���E��
 hAg�'G�0�`L�0I�v颦�,@E�$��!�P8�D�55d�%1�NւL�ɀ��cI���l�\�(9��� ��m�*�p7� �E� �ʢ�y�G�<�2�!��!�r�0�`A���'����2V�'G�Ƌ�� ��o�ud!�T��
 �'8y8��'e"7����g�ca����ˑ4rȸLCs�H��Xc� E�thYu��?����)U�M2�8UM9��F�-Ű�q1��}�v�r�0#�义�$�;/b�'N剬�2�ɖ(��I�feӳ,��v�Fb�h��I�!j�Bl�0Qb&D��C�:n�C���M�K���5	��r\|�����<i)O�Q��Ʀ��Işl�Ov��3�'�0KRIF,g��jJK�>|%��'�R.�� ʹ��"�]�j��Js�ʶ]�h�c@m��	}�
'������[�:�Y�,���'��sv:M?"���e	3�nh� M��kNb��O�1cj�%t�8��p�^�p�"��O�`���Ol�D%�)0�ɎA��t3��A/B����mہ!�1O���8<O ��T��9� �A3m�<�D���'�2"=�s(�Mj��L���{Ǯ�>F���'�r�'�L�C1L�V�"�'GB�'g�]�]�!s�U�D��TAVΝ�/`6Ӗ�W��~��ǩK��ux��L>A'B�2�`�4o��h�l��QOĖCU��@ˋi?y�%��@2�>�O�� �4\i�9�s�Dcpؓ�O�O��OB�8�Oq��	ş�:�h�T�B�`�`�-.JRC�I�}D���n���H90.X�P��4���㟬�'B-�B��L���AqDMG�� 1*'�Da��'{��'��g����ݟ�ͧ`���B
ƈBI 0S���N���]�!ˬh�"��K���d�+ex8��$p���8��,����!|�ĉP�p=��&�,����vE]�L�����l%�`�	�t%�t����?���14���'JT!�����[z�<�&$|�Q���ܾG��QȻ�<I��ix�^�(9u���M����?��nK:!9�}����4U(bZ�?��
��+��?Q�Oi�#&�<� ����<!���*�a,]3]��J5��:��x�˩N�@�E��<����q�h,�1�Ǖ��	T �7̋2O��"�'y(6Yw}r���t��=[`�+�#�"�yR�'2���F�,x���~p�!���&,�B��"�M�/B 5��@��n×gӒ���;�?I)O\��N�V}R�'���Gk���I�L&DLC��G��|ͳ� ]�N��A���$#욧z��JT=|J�t{�S�DU>�$L>"� X��P���W�<}�);.n�HBT�� 
�Xt�S<>~�rn��	��Tk���"d�'<�����?����?i���i�#�TX�6ါ2 h��Q� ��'-��'�!���2�	������
�s��Ը6'ǝ�L��a�1�x�$#kdr��	ş��	;j����ޟ���������u�NS)M�L��#!~"�ռP����"̟lU��;��A
��|R��]�z�[u)ʙy�x��$��{���E�r��I"ʔ@��d!���X���) �՞^����7��>VZ-m�&���������?Y�e����E�z��w�9E�	q�'C��i5Gך1�����kl�u2�O�Fz�O��R��R7J�����
�-ڕ\�����iK*$�IrM��,�����I�u��'�:�64b��E'$pCu�kH ��A�<#�4y�dO.b�
1�e�><O$�p�
�(y����.n�����ޙ(�h	
�Q�_} X���<<Oj
ea*񂅫fBޱ@���q�[�{��'|�'��'d�OP�De�38��$	_�";a�"OT�3qȘ�{F�����5!$$�P��$�ʦM��xyb���T6m�O*�$�/t�����Fh��#�4���O2rB��O���}>c��=���Ȥ$�� eo���Q���>S]���"���$�H� u(�$.������C��(�4I�x�\0z$MмXǓd����MAU� Ҕ� �aNQp�γnH�AF{�4�	͟|�?E��J �k�	x$��0���W�S
�x�Ӹ�+��[�[Q����`� �3U=O8�_�iU�iY�	O�D��0lQB$.a
dx�".@hzf�]I�'`j8Q�ɿ^7�����o�6-�|�)�d\1EE6)u�4h!�Y((V4��B�>�Rd�f4��#R���ͦ�i�7��L�`H�p�N\���DG�	1�&���	ɟ�`J|bM~�Ak�xd�'a�M	z�pA��l̓�?�	ϓ#O��x#�����T�A`ԊD�P;b�	��M���i6�'��[鍋^��I�U��]�����z�$��O*��]�h�v�*e��O\���O��4�� �-C扚�w �E�E=~e��'��:E�F��$���䚴��U��c>�OhUBvl�7)
��S�G�i�a���X-E�8|�Q���x�r �W|q��'����W�G���C�D߂U� �{���n����V/��>˓�?�!'΄0
�A�r#��	�rc/���xҩȡ�Q�M��}i����*���EW�'�Dyۇ�'<�ɬq�"H��ײ��XAFƙ�w[� ��I�$�f��Ɵ�	�D@Yw�r�'�h@�-��X�HP%��9���oeYQ#�+����BMM
��7-úJ����I�;W�L�v���|Dn�9f�	�2P�A�cːOz�9Çb��WTp�[cY^��G��*��'+�Q��Ey�)���m0���A�?���Yl�']��'��O�}9�Jb9gCΏw�"��43O�=E�TC��GʎEt�
}
���A�D7�'�7-�$�+O�������ƟWBŖ~j1�G�ݙbQ|5	��,�	�!aĭ�	П@ϧ ��【�A8��Ո�qO��3C�U�l��u@5'լݸ��1�
�5��h3�y���A��٤ �\@�"��o��Ŧ��O>�43$�>�D����҃kX���#ʓxR8h�	��Ms�\�L���\�0����.m4P�@f2�	蟀��	1.��A�u�Q�(�伃�'&K�C�Ɏ�M����9$��� <j���D��?�)O=:��ߦ��	՟ؖO"��Y��'&���d�*��x��$*
�eӲ�'+R��CS�У�d++TYc�����맅�i�({l�ŉ��н�C���#NXRF*CF^��K�I�(�&p���4����J&bŮ
�����OQ3�'�U��?���?��D��J�R�� �^�*%XB��'��'"�i�R�߾-QzxP�*� �|C
�5��@�k�~10"��0h��&�П���Bx��s�d˜f����.�"c��iRl%D�� �ՠv����6燕_c�����$D�����4~*�!��%�L}��!D�|K6nЬV�T�0C$G�*	!�=D�P�W��ND�,�Ui)�0�/D���W�K��
#�˷��̫�$-D�l���_�o4ָPv��eg��㕃7D���T��-<��ݨF�a��H0�"D�����Ӯw�~M2s�N@>! D����I�wd�� �Rn��f2D�� %��i���]�?����.D���7c�u!֠�g�ab��!�',D�Xc�͏2=h�l+������,D�d�F�Z9?�X����8�P�4D���7-���������5>I��N3D� *%#	���8��M�ycDL$D�2�h 0"�v�%� :����S�"D������u^��ӁV5D����B%D�|���D�D �Pc˓�4Dα{�a!D�| ���xtN����t��i@p�$D�d2#�H+ ��5zQ��+u���B"D��sMʁG�8����1F5�	ې�>D�t�RJ�>1�%�hU�
ݾ����:D��Rd�Y���`�-k4�8�#�;D�l��M ]��� ��8Z��芐�8D��#���]�B�8@ R3+�r��4D�4��i
�2�ջ��B�U�L�v�0D��[@!��1*�j"�A	;4���m/D���#�H�n�x�+`"�~�jK�&,D�m�"B�Y FkE�%��h�5D�x D�<:��! f�/e�`�s�1D������ Q�4#悝:9�C� ߚ�n��Z"����t���g~J?yab���鋖 �%���,0#��.9ľ��d��F!���@~~X�2LN�#2\ s���0�u��hC��9N�<�ȟ��
�+����O�ba�1'À$U��R��dxI��D<1�՚�aP�j�r������)\i�6����B�*�@�L�ś&��P�<\�R�f�|% �jW�������L�m.nQ���U5RZZ���@���M���*�Z6�����-�%�B��M�Ň���]��I��GVU9���>�|9�ܴK�<�����ʟ�Z/�Q��yb��d
��Q��7T�6���GƘc�� �<ڧ2��b��ɠ!d��F#t�i�葞SȜF��(��C����n< �@�}'�.B ���褆���8�G���L9"���l�S�π HBt�ȏu(p�*,�XX[%��	VVV$�c����͓�rh0��'VF-HuKX>[�,�E�vI�ha�'B��Pc�ԟv� e�S�d��6bQ�<+B��ᡉ�!m,�ȳK��%ȷ*D�X�����B�|۰��8����<%?�Q���*ig�%��NM��"��3}��xq�AHOtj��R!�ܔ��'p���k�x�BX8�K�z��4�G�N�O�!j"�S2�D���4�b�xG���	�vY��ސmgXx`�%�7ԊX��b�5�(O���ΰ-�Xy�'��`H��,u|�y2��%�N�p�G�@:�S�y�O �T��O�4+�$-Y�0��/N� �jPȟ��'�
��oF>	ڲ�cBOG�T�: �Ӭ�<�	��_�t顩N�3=��ɠq� 	���Z���'�>�IC��z�G��c�@D�Ǧ/��s�&�/}�������M��>#ҥ��C~���E�����I�<�嫇�{d6�ۜ%(�m2�� �����E� ΰ��Wli�d4��q�m�2TY6�=9��v��%��L.4��<��.��GX��h�U2����'ΎA0��@���ǃk�r8�-B\a ԡ��p͸��O��D�&�&��H:Ǔ~�~aI� wX"xac���6����3�I�B�����'�ʈ(�j���(d�����x`��Dǭ�<��fAih�9���1A����"��hO��[�H
���x�v \�A�`�KC���e�$�(��P%�.a�6%Ӳ;J�h���ƍ"|�uP��"�ɭb��tR���/�2,���Hhj�	+¬ ��≦*	Dd�F�N��R�-���˖�@�zߢ�a�N�%$�P=ҨO����!UB�masg�u�����9�Kc��6v���So	I���wgѐt�x�dWqjj�0��,{E����Ɨ�h��R���8�z��QP�dp���u5D�����N�c�OP�<YSjGd�����߹8�E��K�u%v��dE�=��-B���$�DQ���Ҩt
�h��~Ӡ���������F|���Ty��ʈ\��+b���Zm�TJ)�|�Ĩ�R�VT�g�'Ť���I
��hXW���*T�C�դ:ժ��mHd_D	�a9<�m�Q�A}"BX.HX��efK�
��2,���h&�!��N�8�ġ'"�A4�'��EC\�iB�ik�T$`�k�/�\<�	8ij�'��Bs��[������N� hF%�
tGh0��(+ɾq���'H,�#� R�!qpuڢ�[�MBn}S���"	"��9�"MS�45�,�!�X��]�M�}R�'�HE��#��`Z0�#�6u�PY�D�)��

�:��M��2�ްՅ�5k�� Ĝ�4���; ��Q��X�I@}B/��u7�sܓg�ޱ�ɂuT*}�6I�)��U���97����eɜj>q� �4)�Px�]��0�����3����&J�P$�3��{r.?�I�.p���C�įFv�)K R������h߆ϲ]�s�� ~���4#�b�ٔ�I�K��P"̗�x��n]�"D�?;x��i+�$0��0;�b��6c86zi��O���+��Y�����C�U��Ë�D�DV�x��6�,��W�Y�l�ԍ�Gl%?���ģZ����i��O�'"��ك2a�0JT5`Q�}x ʎ:ې<*�'U�D��q�I�"�Q� �Q��4��c�m�$�����p�x£+Ls�g��<)�D< ��_-ܦ�#sL�V|T �/�w�'_H��L�il��?UH������L�Q���H��A���
@�Ŝj����Č+E���º���sɐ�G��`ϓ*+� �4�V�<�Sf/�$_<9ϓ	nT�wc%vRMC�̓�j���2�N�\w�P`#�T~�(��s-E{'.����ҢȐ�?9�*A�7b�Y�5�^�i���� �B�'M18����v�؊�͉1��E�l �#���j�4{q<�83B[�h����O�$#�g�iO��%�׏R	�hJ��^R��Ѕ�I�iR�!6�tI�TiQ�؀�"�Iؘo�N��01�B�J
F�=Ё�U.T�P5��O9��(�F.��OP�ȁ��&1��+��?^��bg?O2D)OE�iÎ9� +ƥ^*�%閰i%�$��Uɦ9���Xz�j�����q2�̜���n��W� ��"�{�̋�I[�ik�{�f��'�� `N6]��iE Y	 Mߎ��|*���yUR����s���%�I8)��b3�S6~�2<�m͸b���Iv�>ʓuc��0FP*��S�Ɂ�;���pt$H�_↜jR��VK	���H)�p=A`�������M�@�䤰 �)�D���7L��5pG^j��W�dY�D���s�?E�<!'jX//���+�0��QH<A��6�?�ڨ%��9���L}c�A�ʟ�X�C�# ��2�2O���*���V��� ;!r�ǚ~9��$�ʓ:*#>�h� .��Z�'�#DX{V�Q�<V�:tP��&�(	�0��C"!� �A�9�O4 9RC��nLAՇE"kܚٵ�Od�qk�~�X��,؎M�����>%>yz�NP.N�`�WL�"iZ<h��<D� Y�f�Y��X�t�U�Dǈ}�C�=?���F˟�6�,}�O��ODu��I�	qm
��UL�9I4:�'�@�)��;�^LY���j���(�撪o�08mګi��XG���\�]P�&g��"?���	k��ӄ��		*��c�	l�'��u�4i�18P\�&)Q>�=��'~J4h�p:l3�k�4���/���܇��0ec$AW�Nm�XJa��l3 �I04>0�KT�a�`��qɧ�S�X�
��� �'��U0怔Bîd������=1F`ȵ�5V蓻uLE÷Ą<R�8/�/M�>�Y��D<��'<������O�I�U皦P��T+
!H���b��	8�]��>�'��<� TU�G`۴*bԝ�t�Y0�i8f�'��L�&N͹�	��'�>ɀ%E�Q?�劜�f�����F;+1zPJbJ�<ir�OH�h�':\�1(O�X�ՋB2���,6�8����B�� 7n�
���dC�sk�U������0�4&yK㉈�:����1"X�cl�8{Dk��4��Dx��>	J�$끫�J���L�/p�,2Q�I�^8�,���'Lk�w��� �9<�̑���+������hO1�|az�+ڃvp���&K�8X�(s!�C!Rވ�Y�f%�Qdq4%��x*@��s�ԭΓ)���Cpj�=�v���cV�p�'��'�"щ}�i����S4�X��'ih8�U���S��w��ND��'�h�:�F��88 s��T�8�h9�I>q�O x(�h�'u抰��E�5���!�'vyPc�;X��Y��/[� y*��ɾX�M��I�I����Β$,����ʤ��'xў�S�nM:H���"��K�@�\n���Ҭ��;�����9ܙϻq�P �ߟh�~�Q�I��0ZB�	��y�Q�h�S�L��*6ƒ1J݌���Ö�wPT�sCf���zH���DR�.�T]�e��h��#7L]����[:���
�j���kS�ѰZ��S���O�b����"H�ehNxB�]9Cj���'�*T�����X�1��zQ��۴* ��6*G8+�F=�G'"W���U1�y���~R�i(���ǇW�Rf4��� ֎5��la�O��0�	�$F1v��@nTV�����z�~,�`QH��S4���E�ph���>��`���?q�'���X�+S���[��%v���"�-"�b�0��5K~Y��I�X䈙��wo8-�ƧǺG�A��A�s|���~r�O�qt-5�L�\I�Â/@�FoA�z��LS�5&��(���0t����M��^�l�k��7��DI&`QrF�H	zh��蝽p8REB��Ob�D@�1e�!����&+��	�+e��JQT'RM���ڿj���҆%�䁕?Up#������ 	Q�)���+?�-z��G�!3��X7m�37%ʠ�%�<C8p�6X�5S<q�"����cƗ&l�����.E�|"&���}�|h�)	���#�SpiŒb�ΐ U�H,uv�	Ɍ�AaZc��Ch��a2 #�"=�hРK�Of�=�Oq�B��Ҏ 0�"���`�g]}�p�ό_�ax"�~� A�����f���*�B��R�ˣ�:�!�+K!N�$z)On���%x$��kպ=��;R9��O@���k\�1`�	�����ҙ��aĦU�h�3ѭ(7Tx@D��<��O�hA�B�IԊ��!��������V4.e�@�H1i��Qkt�?�p<�rI�7�ke�ڀOX|�g�� hd`zf0��`����l"Y2
�va^#7x� �%��9OV!�!�  ��<AZe��.C�pͶ8�l_9�����_�m���)�S�-n2�D_����$�7��sT��98��0¥�������ϧ[��8�U��>�e��:�hBD��d����TyR 9扱�襠]w���H'9�~A��y1�,!R��l���F��vRV�m��e���󕅟7AVh���F�*wrb��~��~"ظe�ZxWgԍD,��n���~�ʓ�z#n%p�hQ�7+dT�d��hO��	G��+�Vѳ$�ЩZ�������'�p��ɛ3A�kw�&BX4,p��I�x2��6��i ��i�iZ�(F7s2�,r��Y��Y�H|�h�# 6r��$2�㟢��G0�H�1c̶ ��)*���o�0
�,��B>��y1$�׬q[��$�����X╂�ቱL�)Wm�����T�S����/fk����K�60�������6z�D����cFQ��O�z�l�sG`�8#4ne�S�S�
	�d�a�K<[���:rN�z`��'6:�q�
�du�U�R)Ѻl��y����({�sS!Q����zX��Q�O>����+W��`����\���@.QJ��v�.VБ���4�"?8v��.A�� �����4͙��#����?E�d��>@WL8(�"�\�����O|����^;= ��rTHU�Q�2�b����Z ��"�R��偓�G�tU�x�,0�!���qO�1��4��$u��( �Ca4(���D'�A��FĦbs �&E:}s��ThU���4�sӾ�:���:q/H⌖-h3��B6�ˏ#�:��Đ`Nh؀�$��3ғ0m�|{�o�A��j0���J���ޗ'�F�  ��F��y�p��`��O�O���H��J�F��P�=yj۴YivX���!O�!���C;���&OE�>T0CvNYN!, �Ub*rTE��K���<���iJ�qe	O���F�9+��xU��6A|�:@Ƒ��hO�1��`�O^���W0%�'.�\�e���~ 4)�G�t�ɵf�Y{e��PyF�p�OWr��Nƽm����e.(���
1"O��{�b���j�0a�G�U�4���"OT�YT藪@�8��� 1`(�*t"OX	i$��R�ı� ��*i��"O@ع$f�B���pKĆ$a��c7"Ot�������E7͞	<Yȴ5"Oܑ��-�Y��+�MDT�E"O� ��!�c�$q!�z$h�y<H\�"O� I���>9�v���T<43^���"O&�3q�B'-� �H�`XIc"O�@�!�I�`e'P���W"Op�Q cº\�jQ���
�
��""Oޝ�Ҍ�3Og�A�g�Ԇ;��@��"O�u(UJ
}�E�2i���I�"O&����"�:��Ti�I��5j�"O�DyD�ax�ɠh_4~}�ؒ�"O�0Q��If�E��D�T{>�)W"O�=��I��F�
�*ޫrb0��c"O0�BR���!=p��HF?hNB��"OfϘ�Lv٨ǎ&O�2�"OP���$g��ݢSň�.=l�J�"O~@j��Y�V���v��YJ��d"O�X��J�9 �����+F&��JW"O������c\.�Q�
 P�pB"O2hAi�.�����Ћl[&%AV"O�y!N�в ٳ��4H.]��"O�L�QM�4ڍ����$4v�"Ozա4��;*^�ZdbK�=��"O�C�o��4���h��,/&5��"Oq��B!U7��+�˻
hC�"OjDp`�-2�����F�7��Ii%"OXZ�IT|�8A��D�� ��0+�"O�"��ѳ(����Gi�C��t"OF�����Dx�'ˀ6����q"O2�R
"(Iv�Jcl�"|߬Q7"Ol�%��)��m	��-谩;�"OjP�u��!�l��
Ź2b}(�"O E�倂1B��H{�˃�I�I�"O�9sDE�]iN���@�VqZ�"OV����B�eVq�VL	����{�"O����b�/{
���+W�W*L�"Op�0��RR�,y��i�Cr@"O؁�R�Ֆk4�����?	����"O��*G���
Q�e��?��0��"O�HfC�'�R�Ra�A�\I�"OܠjD�?Vj��@�)FL���"O���qi��*:�����%B֚�yR�ؐw*�aբ��")hPK�)�y�b��F���Ǵ�&��䋀�N�pB�`�@��M�/�.�K%�^#oJB�	)}��\��݈r��3�@�nC�	HU=�w��17�V	���t�8C�I4i�0x��0�P]��`��,�2C�	-f{�I�̂2'��2!�é02�B�	��\dp!��4~� ��tā�SΰB䉛8	@E{Nۘ����a�*&�|B�	�T���L>/#��h��; ��C�	fvڔz�%���R�q�Μ?�C�I��l�2e��~�|�bL�T�`C�I("���#�OF,,�$���9*C��.T5r�����d� ��H���B�|TJ��A�HlNԁWgF7N�C��(B�8�1��BT���r㎤g��C�I�<L��R�٦IG��Z�CH��C�	�f���١��>\�6aq�N�[m�C�I�I�Y��!��3Q/��P�RC�	;I�‒�Ǆq����͕&D�4C�ɚf�,��!����hqC̈%XF:C�	�X���9A�����\� k?hC�ɧY���kr�R�=y��{5E�$w[6C�ɚcz��J#eW�1gpX��o[�� C�)� ��R���~i������96��$Z�"OZ��W� ����	�%̊���"O\��l]I�Ĵ��&�'0���Z�"O�j"�A�_��X�6�O�wP��Q"O֘���D�"yr�رu��˱"O��F:����Z6y��Jg"O��1��Ж!�%���
ai��j�"On�ԑ�����(�{���rp"O8���ߢm�B
'ŀ�����	I���'E��c$Dۘs�� A�n��/Ɍ1��'U��JW�ǖ^�ޡ�p��)j�HI-O��=E��hW��=S��K�N
�R�7�ykC&X���b2���NN���aT��y�Dj�MJ!n��G�~�*4H��y�e��*�0� N)G�H	5`��yҍ	:l� �R�9���T��;�y�[9>%�baL��-  )����y�DZ�&�j0#A�ι2��t�R��y�.�O"�e-�cJ~�9�X��y!ӟ[��A�5aD�a�ތ��D�y�S�m\:��T�ןT�ٻ!/���y��v^��(S�� ]�HL1����y�L	;b8���D�U��[�,\��yR/G�kwR	�#�U�,p�;�y��Y�f9�aA�|��Yr0�D��y��*�T�X-�3x��q �Y��yR�ƒ;t��w�&wn��Ӗ���y"�֫]�CFn�=l��Yb6�J>�y�ʠbz��R�d�(.����m '�y�� <v~	�L"Z�HEi�+�y���BaBs�Ϙ�ZL3EG��y��I6˸��D� �t!�PXD�D��yBm�0��KtN.=^p�n��yrLֆv���&� }�\s��П�y"��Ќ1�kE���9�N��y��
!_��q��ƨ2	���$a��y����<�C�D30��(T�S��ybG�U(R���#(�a d	�>�y��ā	��J�WO!ެ���Z��y��}g���ϢG�,��ȸ�yb� �X��d�E�#����C]�y"����,��%�ԋ��MhEd-�y��ً:��% �žFR��$����yb.�25 �������$ C��yB�,S��tq���*"�L�$Y��y�ΟI�-��t�X���٢�yrL�S(rH�4 ]'��yK���y���\MQ@s��n���f�	��yb#��7Q���a�Y�q�*D*Ɔ��=��yJ�b�~�B��ؒRnTe��DK��y��Z:r(xd P�JĒ2/���y�-�`��g��4>�����E'�y2�Q;�U%3��p�*T7�yRK��X���杦/~6��W�����x�Ŏ';rt��b	�&A^�A�D 9!�8g޺-�$�X�<��l�3���M!�C�n��e��J�3hV�L���-]��O���tmY�H�c#� 6���'9�V�Z8)�Ybƽm,�
�'�\@R�ЩW��l��'
&n��C	�'�2�83c��i�8Ր&L�i�.���'
|�Hb-�6L֎$��jK�`M���'0"��E�='V�=	u�,z��
�'( 0p�KM���C�L�/ <z	��� *4(���%lk󢘏`;T�Ce"O�Sb`�'Qpd��V�+z~�`�"Oh��Gn��	��p!�̘	 ��Y�"O*�kpoG�I��-k*Q�5ꊉ�"O���d	�&qR���Y̔� �"Od�灂[�9���m	������y҉�hq@�A�b�&RD`��]��ybHհ��0�$� �����]-�y��콻(ߤ7N(q��.j�|B�I3x�&����/F۳ڽ[��"<��'-����ӃyL���^�1�(�
�'4�;�H([�����n�-�݁�OR�z0�5d;
����eښ�[ "OT9+��YOd&d`RKݜWtD!�u"O�� qH��Z�H-�q	��}#�"O��kF/ܙ:�"�0� 3��h0�jZcH<9����8IA��ř8�C���j�<	BJjN:X�#�?F�2t��n�<� �J;�!� kR�"���R��k�<!ԇ	�8���B�$\0`��%f�<������|�D΀��*9�7K�}�<I�
T�Gb��ig��|�yH��u�<Q��ϰY�R1���jv��#��Wk�<I!��$��%��ہ`ܸt��!�f�<��J	?A�T���� 	]����w�<��g�#K�X�ԦY|Ӧ�b�p�<y�ER+�@aȦl�=5��phl�<��l� ~����5c�Z,�q��Ȇ ,�!��;,����$DF.pIRN�+�!�Dӛ/tL"1��k`,��D���qt!�dBY�T�7i��3W<�crI� fm!�� �=�b�$�V�;�gt���ȓk�2�%�R&eސmñ-���ȓPdV	*d�݉/��i;��H"��y���͒Gg�/x\�'�Y+⼇ȓEO��� j���0��"�]�G��a�ȓ��3�&Ʋ �(�c�gR&;�P`��e9~��1�G0.-4�S�����'��F{����r��R��R�j�cL��y2�ƚx~t1�# ��%!c�0���6�S�O���0���twԙ�B[/zZ���'�~�  Z�j��L��ضM;9��'��I�b�:(8�KQJԮ>���'���K�\�Fv�b F�3�����'��I��JPgy����*3\ً�$<�=�V��4��}� ]K�F�&)����J��i�@� JxT�؆%R�b	r�'gI�p�ƏA�j���.Dv;8�b�'Z����i`����Ǩqn�A��'�&�&�j�8Y���5���0�'S��H{��x%��E�f��'>R�A�*۰�Ñ�M�ME�\�C��4�y� ���qGI�N2zI��"�y"(��)4�цv��ug�U"�y�V/Q*(*f��6��e�ɇ�yr�R�R�<��ꗎ9^y�!��y�����H ��PQ@�,�y��+ U�qi��.Ɇȴ���ybF�&Q�}X�*R9v��)�DNX&�y���`�,�3q"ư��W�P��y���F�HI1B�W�������yb�d8�|X�FN����Jǂ؆�y���9b$�y�a�B��ܴ�yR
�꡹�P�&����O��y
� ������A�(8�␳< � Y�"O�dQ0D�&��d`G�5?X82�"O@�z�cϖV�1 I0oT\T3�"O�a��C	�a;@�9'�ѩ/5(I��"O֥��� n-rO��P��i�"OR�+�.ɗMX��Mj��y�"O�,;�g� vx�*�c�N	�"O��*��÷d�A���4��"O�\1��J�	�Dð")��Ȥ"OdU�B[*�z59�������"O�9 �`�<��0cE�V�N�HĒ1"O@�ѵ�ƊN"��6!��)� �K�*O~L�Pm�O?앺�@�R���'�����*:ݖ��um�K�"Yy�'L&]!#��'�>�B���-�zd@�'��|�&A�(�f���N�*���9�'��� ᕾ�Hը�-	m�t ��'6��_�'��j����͐�'�H�2 I�3�����S[�hl
�'�(k��"}	�B@#d��	�'�2a2En< ��cB�K
�'�ڔ)��٪XF�#1���W7�P��'�@d����<(��Ӆ�1N�E1�'s ���j��T�,#�*�N Y�'V]�+N�p>��t��0�����'��4����vg*U�WE�|ے���'��e���2F�f@�I�f�n���'b�� �4Is9�6.�*`�U��'��qrkΛII���N�eL�`X�'\�i����:gQ����H�R�����'!��kD�ӿ��� �2�Q
�'W�H�Q �t�@H��Տ`�2�	�'�ڬ��cS78����������'�@!q���E�ؘSbU�'��I�'��	q�
/��@JR�^K��'���B�Jx�ER�B�-
����'�
�peLn �@�we�	 TXQ�'�py����=.lJ5�w���PE���'�M0f&�6LZ�j���Wj�D
�'������;���b�%&�uq
�'F��aQ�E%8����J�.�24s	�'� �[�p�EJ�J�8���G��y���?zt���)��0�^���
 ��y2��2%1҅�ʝ"N��I�&ͯ�yb�@�?٘�	�с�U�(#�y�m�97�X�P�㎫:a��D��yR)ޠU����焮/<�Ay��U�ya]�j!ܼӃ��+�h��ĎO��y��,�0| �lH�Yz�7��y2�ٸ�2)f/�	�n=�f���yRŘ=>n��3�N���)�Uk�<���V�*��q;ӦʅʂPf��~�<i�e< K�H�fS��v��Bk]{�<���=:)LXkÃӅ6��\�q�<��[���i��˄^O��R�/�j�<�� %I'*�*���(?���#K\q�<�Y��2d�m	(C|��"Abg�<�' �:��� L�=t��Ju�[z�<a���<V�|4��퐲%$Z�dt�<��b�$��Y#$���#����rn�Y�<�6�UF�8��nF�G֮���cU�<Q�ô?ܼ���?)�L`��h�<	gg�-KC��PA]�\mH|�c�{�<	���#�:�`Ѭ7�t�֍�a�<� �#i"� ����
�K;�E�"O��!�%� K�$�� �V�`��"O�2$��yEL̈��܄NӲLaU"O��I2_ ��Q�Q/�H�r�!�"O�:W�!+�h��R� V�dU0�"OH��s�()�ʅ��L	�
б)�"OR�z1��e2Z|8aBP�d�0!S"OX$�4Ҧj�~X�ǦU�(.���"Oh4�R&)�h����ϝ��H �"O��HGa׌l;f��	PO�IY�"O
1�a#_��������&U���"O`Q�1o;LoJ�C�#U�z�"O(�0���F� ��'�98�E�b"O
��P�G����˓F_ZP��"OP۲Fo���%ƅ\ӦqPg���y��s[J��".��ZB�ih3�
��y��Y)yw������f3�u2n���yRF�k��Fյc�
E ��G1�yR��	Kk0Y� M�X;F�`�؜�y�O 8��)H�ğ!T�Y��D�)�y2��J�^�3&L0�t�R�m̠�y�)�*�aR�R� ��`T2�y@�>���kJ0 Ԏ^#�y�+G=�|��򣊂Ld���U�y�FV�{���y�(%3	��y".
)v�ʽ�fBŗF5����F�y�b��
��-��G�S�������y�E�U4�i��9T" ���H�2�yr���}cĥӲI�>|:<03NW�y���r#n02u�84ɀ�b
��yR��c�z򦜴/���(����yB���S1N9K��L�'����v9�yBa\�U�ΖuAj|��YV�PB��Pڈ��Ä�>�@�FFW(**B�	0u.�	�c�e�6PS����"B�	�Rk�ax���j�j���n��C䉛%X�Q�$��Gn�<BGP�/��C䉤'��	06g��0�ht2h�C|JC��<n:�3C�*�<�!�Æ%FklC�ɩd�80�k�*3x$�h����C�	�v8t��%�X��u��/��:�C�	�&\!�����5��) �bՔk��B�	7?�)���g �(e˒Q��B��#AI,=	�+�#K���/P�2��B䉲�x��5J#�1��h$ڤB�	� &v�:�� �l� �#k	�I\<B�	��GH� ��")J-A�C�c4�e�Y&��̸��B0B�I�^��!A��:d7<�d떥#w@C�	�6�~�Sq�F�>8$�[6#U:?��B�	,.� 
�K�
��Ī���NN�B�	,��[ó�"�R��E�BJ;�'��a*�$��c�~��6N�<���!�'�X���'w#��
f;.?$)��'0��G�"#�$�TȖ�3��Y
�'��|���&]dXQS�P�+���2�'6�ۆk��e�-�G�ݨ2�<�	�'�ԡ�f̎U���� &�|I��''
�ȅ�I�0晻�j�5�����'�TD˰�AD� -P��~�(�'.��@�W�l N���f�0!��P�'΂}���1Au�j���*B�9��'���E-W; I�a��*;d��\��'	TA�B�	#��h�Q*
����� �����ͣPq
G&�n�|��"O���CE:V� �DI�gI��"ON���hțv�����B�6;8���"Oؼ0h̿id�F&��K&M��"O�1��,��]���_m���"OH���ݝn��%�u���v�(F"O�Q����E� m!Qb�'-��X�3"O� &(^�5~��� Ůyw�h�4"OtM�JQ�6�������6jo&��"O&	t��o]��ɜt�2�i�"O\��űs?\��G�>?tŋ"OȤ3���4ވ�@Ɗ�:鐑"O`���ۭ�,,x��L&_X��B"OTC�ꍎ�( �S�A�V����"O2�%g(s������Yخ���"Od�@�\!>
,�`��O�~�H�"O2��%�`:��G�%��h�"O����Uk�ڭ�$õi�&]Y""O�m	��[1p�JpFQ���d�"OE�V
ښ?jB�S�6a��"O�3��f/��:�I�6X~���"O�����#�����Ŕj�(�Y�"O<P	A��'T��Z�����yR"O�=��h������w���j�"O �{��r�6P�#[W�4�a"O"���\�-�|� �`�{��"O̹�2��-\<P�d��@7"O� ;�`�$�F��րG04K�M{""O،"� R��x��9y�"O�b��&x��Ei�W86�F��c"ON�Dl��-�䨻�c�`(�"O�I�o�����̋'�6�
�"O����ꔍlL�T0 �D��XIP�"O���0�.z߆�pb�=�@��"O�Ւ�FN#f������E2�!"O�9��.�<`�,	��M�L�c"O��å��c��PP��I���"D"O4 [ �G�]��:f�L#RlM�""O<9�/�fysV�Ѳ��� "O��Մ��Q��ݒ��L䉆"OHȣqc��<�(����;����"O�l���̶,��H�k��8��� "OV��L^���w��)V�
a3�"O|Y���W"J��%iYh�"O\q���U����r3�.a�(�"O�@8�̂�Nt�F\�*X ��"O4�(���?5�T�v�Ã.�rf"Ol�@�y���	�$J.\�I"O�eP���i���D��Am�̓t"O�l��*(�Pj��R�`Y,Pb"O��H`� s����t�C�|F�-hr"O�#�8��x�C�S4�9P0"O��3u�ÔNmr�AUkۗx�$�4"O�*��� �	�(֍FT��"O��s⌓G��Qh�eJ&zz�U"O�+�dV�oZ�lhFI�w]��%"Ob$ԝN����ȹdhJ��"Oay5�*T��S��˛-�(��s"O���wN�*������� ��P"O�����G�I�P���}�D0Y�"O���.��8*��1 N%����"O.�b���J��*O�W� ��"O*4�"Po�z7�7p��"O tSw˔<}����@0b���"O�  ʔ�F0�N�X�/G;�d�s4"O��P�Q�����Y�FK8��"O2њ���B�p1c��V�P�8"OЄ)������AN]�5�r��"O����%�hH�̋�w؊Ic5"O��iʬz�`$�.�:�
���"O�H��P#n#�h;0���:�U�<Y��C�Y"v��!����Z(�2�N�<Y��'�ƕ�u�MD)��1��Q�<���^�J݊q�M8!����,�O�<�+���n�F�)�(�֬WO�<�T��nEJj�㖹2i�$9F��K�<aT"ڬmZd��䓷>�� �u��J�<���+4�L����aOԐB�Q�<	���-��1*5�Y8g`�UB!�N�<Y��Ё_�(�Jp�N9K#*Y!���G�<9��ߏVu*�0*&8�w(EM�<��A3/�t0����)u� 0�w�E�<�W�M�q�$كP��%P���8R��H�<-��Cc'D!�|�eQ�9 I�ȓ2�����P�е$�%	1�t�ȓ#���b.q�,e8ӣN�6�VA��|��(G�w:�k%[�7���{�y���$Eј�����0\�ZQ�ȓ-h@�`JS�0�y���{L����8�s�BW�eQ�5�Ō�|%�ȓZ�� r�!Y�)RV� 7�M��%����f\!R�l��+��I|����;���B�3CC�)u�G�E�0��OGt%!i�{m��z�n�6\\L,�ȓ����A����bF��C�:1�ȓ�W
'���RGхr��0Sf"O� ��J՞&��� 2)�W�<J1"OijvF6m&X���B&sgP31"OH�ȶ�@q��I�æɌmKd�G"O4-d�ԟ!+n���#�q�*�3 "O���b�~I��I��24p�L7�yR��?�J��Ї^��`42n���y�	G �ʉR��
��BIRC�M�y��*|�b�Q�	u�`�
 ��9�y�ăi	,1��,6}�B�Q����yB&�l�:fj�x0�X�S�K"�y�L�/��hGS�v��%�#�F(�yR'Ʃ[�Rr�]v�Y���	��yR%�ᔠ�p�f�#�n���y"�R�t�m�t��X���JD��y¯�5����p���BT�`�)�yr��<,]H8��J,8��u���\<�y".�z*�бvE���Dp�G�Ϥ�y��L!!zD�1�ͨdM�p����yR�;tMdUc��G�]~�X����y�o��p�R��R��a�Ϝ�hx�UB�'�N�j'l�|�U�T�([a���'-������L��i��]T�M��'�*M�� ��^t�lP��H�OH��'� �J�	�H>F��@d�/3� �'}t�P��!4>�5ìP���4	�'���`��:v'lY �-��1\z
�'M���E�ŏ~�Z�c��E,wh�Z
�'�d���@G*��{ �ݕC{.�q
�'�0u�׾6l�z��J�<.B��	�'X�\���ĩB�f�{�+�=&P���'c(����J�_����v#��8�� ��'R�a3��,ת�P����8�A���� ��G"J�B|(I��P�LHL4
�"O��ҩ<��I�&�� - ��"Ot���f�p�NA�̊!wl��b"O��"�$q��Xrf	 \�ApV"OP5sG�������⟘|��Aw"O�}��H���P蓿YnD@�"Ox!��c�`�r͐��:�Xe"O^�C��]����l\��qF"O��B��	*j���#ɛ+CX~Ё�"Oy���@�(���2=�m��"O6�qF�X�0&�d�!d[ o���"Ov�cGͪF���F�Q�F-r"O0Uy�%OK:���@;yS�{g"O~E�-Rz�ICj��h� A��"O�\; ��,�����V�ъ�X�"O,������Z?�T�&O�Dƀ��6"O�U�g�--��Ek�%\�0��%ۣ"O�C!#̄:.���?�I�"O:mK��ܲ*�IX0�N�Gz�T+�"O�,��Hӎ���('��p�|��"O&�p� �}�p�eb��i"OTm���*�8;`�֏S��Zw"OZ�K�D�%'G�=1�D�n�y�#� _RQ{� ū:�}걮��yrjB�q�h�#g��#2�@�!QN�+�yR��oϴ	Jky=�m�aՌ�y�"��k�l��5�ip�� Oš�y�O�|��)�[�����,	��y�
Q?u�v�.VFN�Q���yB�_�<�Vi٢�	E:�15)��yb�'=�U��l
'nVh	 FK�y�oY |�ᰵ���e�V�;w��y"�H.S}����ȆTzV���J�yb�U�p5`!Ł�@�L)�A��y��ѼZo6�� hG�>�i��,���yBC#&�l4�V�&��L�kÕ�ybI8z4�)�E�0'��\���yr��2�`��#U�%�i��+X�y�N�"N��e�eD��!`l���j��y�h�4^`$֌Ŝ�2,��h��y�N>)ց��iͯ#d��cфS��y2)�R�tD��a@PX�ʠ�M��y�H�Nb�����X����� �y�=�IC/M<u��`����yҌJ�`6\,�5���|�C`͋��y��Ӆ	���9�珜��{v&U��y"n�:E�*tZ�!�G����� 8�y��HݾY��C�,9�6������yr�W&��Ԩ/>6!cV���yR$L/"뒰�@�>�tpy%�Ĉ�y2'�37)��`A�M�8|�P( aC�y��.��$��c�#4��Q��O��y�13�}a���?y�����ٙ�y��	~G�� ��!;��Xc&��y�jMҴek5�V�:�,[s T��yb)�(]ߒ����_38Ь�"H_��y�C���qo֖w;Jظ�A�5�y2�з<Q���bD�~	��D��yba�>$�\�f�x����,�;�y��~���;rK�l*2���ؙ�y�c�,ej��l��4PJ	�r�S��y�LH"T��s�X�b�U2��=�y"�G� E��c�ȿ]���rt��<�y�DR����:w/�[g`D2�LU��y
� Z� ���)X}���$`�
���Z�"O,)�'H����H�@E"%���"O�x��>~z(5���@�,�XB"O88pEeT��P�ǃ)�b4�"O4!ۏYE�IE� ���i0"O>�8V�ѾC�|�+�W�X#8�@"O8L�4CS	�Z��
�@�HD"OL��w
T8h#�	/X�)*"O�%�ĭS�Kh�A4�Y�fU��"O�Ћ��D�;ܒ���뎮$�F�J'"O|�"��_����@��\�B,��HE"O<�R�/ªY&�Y�3��,X��0"O��zE��kB��!b��]�L�8U"O��cBǴf\��;$@��Z�t �"OvM�p양<N���B�Y��#w"O���N�[�*<acBH+�hxJa"O���V�L>R���.�C����"O>mkf�D]���瑕n�y"Ol���U�~dp�/Ә~l�h"O����C]9f��`�&��s�"O��37�Uz��1��E^*��"Oҝ�T#C?�b܊@���T;��"O*ej�˞/�� T��v4�Mh�"OD`t%�?�Rx�� -!x M�"ObQc�mq�(p�ϥY.��"O`%�wiՏx��)%�H1bjl)"OnE�$4S=�9�� ܃ZQl��"O�H�d�N� T�~+<��"O�{g�8e^���jW7'`q�6"O�	1v��%x���P�O�%�D���"O����82����4�Y"2�<@xr"O�Y��Bӷs}r��X�a���(#"O��Z9-�1�M۫B��e{ "O�p邥Ǟm���{�M���"O
yJ6L��T�	�[)H*�-*�"O��n^�S���2�Ȅ5��R�"O�9�iȆ'��)�5��4b��B2"O.��S�)tw2�gIRV�d�r�"O��:cV��cEN�[�Pm��"O2@@v��;9�1�S_,��Q�"O呑�]3{2y���+���s"Oj%�CȚ_�>]���!��y�"O��$	�1*����=~����"O�j�GA�o)��� + w�$�&"O���bOO�FPj0AQHî;�Rta"O6,�`�C�#shiA(�'b��A&"O2c�*��mI%'��'���c�"Oy:SZ>������0}&U)�"O�X#�аpjM��E�_\D� "O�@:w���kۺ��w�U(|$�S"O^��#�ڒC�Z� ��-,pL��5"O�PJb��Q��t��N��<H$�""OJ�)�F�<�hiQUC�/D"O�3��@Zk�B[�x����"O^��!ݟL�
�ơ�(J���j�"OB��B���DH�+`� �l��r"O�L+�$�,�c�.��v�~ �"O���c�)>(�LQ᎚�\���k2"O��!��TZMLi�MΰQ��|��"OJX�c��K��l��˂}��5`�"O 􋥇�5Ժ��Æ&8�"O���A�5d x6�4,Ӱm�"O���GP�M�bL#�@9W�PlH�"O@� Fˉ-���R`�D<�"O� r=Rq+��y��I�Da�',�$)F"O�pѥ�D�ݪd�
-v)�"Ox�s%�Ԑ�w�ɶTԜi"OJu �B�9|s
�ö(��.�fp�&"O��3�)��4����ǺD����G"O6�S@��
���h<$*�A�"OHઐҲ@�D�!6�H�`j�T�"O8X,5�Aٷ�ص1Z�4I1"O^��c��J�)�G�L8�xA��"O ![�BA�tB�����4W� ���"O<d��ȥG�*�`�G�J�dd�H�<��GT�������Y�B����TO�D�<�qNP$&�t�"t�;f>����k�<��Փ<� 0��ζ> J�sF%�j�<���E�1xN���0?�Lc&�e�<9AمЉp�#f�(�˧/�e�<����I/� CeÝYՎ9S�ij�<!D�ͩq�Q�"�(� I*�k
[�<�o��6����Th�r�(�����X�<��oJ o�� ��&z�Ҝ�u�UQ�<H�{z����S�q��i7��K�<�����/H�QB�Q��IK�<�U�Y{��<�g"4XHuKC$Na�<�
�N8J��6���!�H�<�2�63XAe�ڽR���r*{�<��C��FdDL=L�(�w��M�<�����:�q��CE��h� ͇F�<�&m��{VL4���JIhP�b��x�<I�ֶx��0��̐�
:��u��p�<1t��'1�0]`@�B���a�n�<a�d�>Fb���0�j�|�� h�D�<�0�D��0��Ɛ1f��t��I�<�"�A?�jXb�����U;R�G�<i���QZ�Ͱ2M���H\��K�<�A.��k}��qG��t�(iLN�<	��Q4@&е*��m`� �J�<1g�<��x8b�f^L�)p�<��
O��*'F3KՂ���Sc�<1��T�Gb����6x\�!�f(�h�<�Ŏ[`�&�(��3��hid�<!PߟVr�[`h�^VD�pda�y�<	&A�@鄐ф��o��x��w�<�RH"x���I������Ja��r�<�$^4�Rtb�͈Xb���1��r�<1QSv/�9hd��q��݁BM�j�<٧W4Z2��c���-y$\#��f�<�v�ˀU��P�Zo�P�*b�<�w�]��}��c�P�vș�]�<�@�C{g ���T!e�@��L�M�<I�ǂq�"���)�����;��(T�x�'��{'�Պ�,ɧ���2�,D����@�=<*Q��Ȍ7g�	��j)D�<�7DR?P u��çm�����-#D���R唘3���a���$�)c?D�`�DǺJbh��L��VW���O(D�೧MK:f�`�*|'\���j$D�|�`c�V\[��[�r���C!D�,�+ �u4�C�k�b�[Ҍ>D�p��B� ,���9k�>1�sn<D�x�$@YB���s2
P48i�q�;D��� Җ%8BMD����F$D�Xs�B�EF�t�OHkjA�A=D��;�әz�J�х��]�Z�k�<D�pŨ٪!j��eJ�y�����%D�� r���K�xߐu�a�@�H#��A�"O*���Mߠ@{�tU`<JJ͂�"O�*S&Վ	P�2f1L���5"O�Ɋ��� �&h���5�p�I1"O�uR��O.}6Q�e�ʪ߲��B"O�!��.��5�x7$�j���2"O���$@A
qS�솃\�Z��F"O )"2w�@ �c��9�xej�"O0���¸ Ո2��"��,B"O�
BHT�%�ب�j�"���"O��cȞTV��P̘���W"O�x�v�Q�e��d+���@�p�3u"Or�p�E��p����ܑ�w"OR�e�Ε�$��#H�s�<��"O�e�V���1�����^4��"O<���L�c�l���D�n,��"O"X�B<F:�
Ń~V���"OLS�
M�^�vM3 ��%��A"OڔT�I,}" �K��=Z���"OҌA�C��b1�AP
7q`�ht"O�P ��X�2��E�%�Ô)��H*0"OҤ��ǐ�4��h�G�J��,@P�"O���ǵ�W�D� MR�R��p��"O�*t ��FE^�J��%��@�"O�yp�Ck�a�V`�v#� �0"OD�&�K�k'(5*D�ڲM�4}B�"OX�����;Ǝ\5n�!f�p,�a"OD,Qa΍�&�R��w*�u6�TC7"Oj����U�z�@=��Q(�=�""O`�k��Z^�bG��Y��"O.��$�j^��"��M.�y
�'=Bup���;Bjt�z�nR#v� �	�'P����� �8b�B�b���	�'0���v2��(�HǛ*i���'���(��$O��$c1��%ð�#�'1�q��F���Ճ�%�F��b
�'K�cG�yv@�*�LmL�
�'���z$�Ѡd��C��Td0�'�^���E������vF�:Ͱ��'���h���$b[�y3nD��'%"8�FFBeU y�L��[ ԣ	�'��! W��'�`���]�pȑS
�'ȔY���n���v-%[V:!(�'��xrBOMmݼ �ՍJ�j�虑�'{ ȠW&@�?}\��_�j̸u��'?��CW�N6O�4�ԅ�4d'���'Z�!�`��2CD��B�dD���'�2���K�W� �P��W��P
�'��m`p#@�w!�Kf(��L�(z	�'�*���P�4>��bǊ7��h
�'��A��	�Bn��1&��
�'o��;�o��x��ڢ�;9�v�y
�'�l5�Qg��{��A2��0�8�!�'D�M�j1��m�q�0yQ�Ց�'���coD�$[�٫wq��'�¨Yt�L�9%��`�p�X\a	�'�	험nvf��`@�c�KI�<��o�9|�����^
v2f,#`)F�<�vg�=���P%D� Y�#��C�<�'Qo�����L�XR)�@Z@�<q�Z?|
�)���Z�2���⣠�p�<Y0H��߂�Ђ玲+9�AV��j�<�v�/a�Pd�U�­r���X���c�<��̋'}�����J$ra0�$]�<� ͪ�L\<F��B�0|����f"O"�
��QcuQB���)'01�"O�� ��+�DuA�a��6��3�"O�(I�ʂ.�H�d G�,T(��w"OH�B��0��/D@���'"O� ��'d��2�O7G/���"O��i���nm�բSH*"Q �"O|@84�>CR� 7�߿R�� !"O����jȴ@pB�/R���"OJ�E��7Fq����"`U��Q$"OF�2G+��A.��T,�>D�x}��"OV����T��9īZ�LZr"O��2K�Xo���߬-�x�$"O�!�V�6}�`di�hL#߼PPe"OD���	�J�Z��W(I�H�"Op����b�5�E��"�p�8�"O: ����W?� `FӬiP�2�"O���C'�9C�DA�Ň:p�U��"O��9�兿m������UklhB6*O�}��ۑ<y��H"h_+B����'�3��áA�l����L�����'g�����́' N�a�B�9Hd!�
�'����� T��Q���)_S:T:�'�x����$z*(�3�/#��t�	�'`��sl;ѢT��Ƒ��8�s
�'���W"9OK,�p$^�n��' �}B
�6_�	�TO�:��E��'-�\WK�*��53��!
U�y3�'��Sa�g����_1T��	��'mD���A���c�.XZ��¤6D����7|��L�k�7�(���2D�l�"JF�X��#�@60]
��N1D��X6���\�B1��G����֭4D� �Z�Yk8�gE ����:%�2D���e�N�<�yB��+a>��3�4D�����ϴ���:��F|�0q*6D���w�
)j��#@L
Z�2�(D�Z���</Ǡ�`C�I�a�<���(D��t�+W��9��NR%x(��f�#D���3*�[.Ut R;:9�e�%D��ÄKX(%@����iL-j�XI`�/D�(Ѷ�C�	,�{�@ֆH��Р5A:D�4KVΌT��h�񅐌plH��6D�Lk��ĉY��եR�:(��G4D�ɲE�7�P�)R�N-Bp��0D����b�;A(2�ʌ3WO6|5�,D�<��F$p�U9A�Q��xg�)D� RR��3���X�#�)>>��3`<D�Tpa��w^Ԝ��/H�D
�J;D��P����΁!3CG�O10�8׭&D�����ӕw�Tk�L�J�ڜ�e*D�D3�H�RL�xP��]r�s�-D����B_~��9��9-���#6D��`F��^X���@�3&x)��?D�x8�n^3"4$��P�.f�2�U�<D��:�^6WZ@!�%��=��!�%D�X&'�]!b�E��?���G�#D��[�( �h����bŹ#��HA��/D�pp!D�y\�ɐ�A�g��饎9D��S�ƍa��0a�b_�nG�1R�6D��R�H_z�D=�� ӭI%,%�3D���S��e��i+5&���}p�)4D���0H�-3��̊46��u��2D�\�TA�:e�à�M�_V,m��%2D��  �"dmh����E�a��5"O���7�٨#�]�Q�W���i��"O܉	��YY�
0y����X"O�X�W�դN@�����ų���"O(2��w����  ��-w>a��"O�U0��]�Q}L��Sn@^9d���"O>�T��.�j�.$��Y#�U(3Y!��2MЭJ$h�-"��9��!Дv�!�d����l�C���4
#/��O�!�d�Ӡ���O1j|A���f�!���S|.���R�nLR�@��)28!�ēB#��V�C6hhh�ࢍ;i6!�D�_c.8PV@�'�����i0!�d��0��D"`"�J���$  D�!��	P�1hv��	L̌k"�#V!��?"���J��qi��لV*%=!�ާ�=�t����=%qČ�H�<�L
��d�P�����%�z�<a�JC�m�������"&@1p���w�<1-�)w�^�At̋�&��L2+�v�<a���9�D�R�T �,�C�OW�<!g!���% S�^�x��8��L�<�S��_�����D�-�G��E�<9U��	���3"#�
4�гC��~�<	�"�2uV���d_�zf"����z�<�Gk�9?�V���*I�N�T,#bH]�<�0$�%|��C�y��*T�\`�<QG/۸7�v�ˆ�L��ԁo�w�<��b2�>4j�<.XUy �|�<�!oB #\�1���Sb.%��ITy�<!4F8� � &�%�c
v�<Iu�S�t���(2� J'yh��Yn�<Iva
�U���s�ȋ~�F5 �U�<��O
y@pā1���ك�Q�<iv副G����2� -[��؁.v�<�#*
�hU ��7@�=Q�ت4$�n�<�!���7��Id }����+�n�<94�=a��@�%H:�(�KVa�<�q�Ě{UP2���e�D�[�<��@PY��Ԃpd�9@��Qc�S�<��ƽk�XH�J��S�(P���.T�܀E�R��ز�B!r�����"D��A��V�[
xԲ�FG��`��?D���$ &jb�Xځ��6�)��=D��Q���QP�R���5G�a�7�=D�ly�G"X��Ґ7|s�݁�>D��2�I��m&̔�eY�!: )"D���c�M�t��ғjt�!Â3D�<����A�\�A�� ����0D��; �=~W��P�B�>�`e�6�.D������N�Io�%"��e�,D��Y�Q�0а�,��{��#g,D�hc�G����3�I�D��l�3d*D��@V�GN.�U+�l��P;v�)D��z���"uj�)�o-	�,"�$D���E�Q����� V~`C&"D���D���)zx���G=(�X��h D� ���D2��`a�E�cҪh86�(D��b@�֠(��z����`Npx��'D�P�0���BM:���C�}�����+3D�0!�ψ�)=�`T��5~��0D�(�CC�>4@�)�<  bo-D�(`���*-K,@
����;v虴�&D�H%!P�_�0���i5��HҴ�&D�� :D�fb� ;P8m��L�-N.�!6"O�`�"Ǚ���0��Q�j�"UYQ"O��
�J����x$��7u�B�z�"O�To��h7��'��� ���"Oh]yI�.ׂ�SD�
����;7"OV(k�n("�ܠZ��\ ["O�*�g�1<���ڀO_�Q�X
�"O���n��z�+gǙ28�B "O��[����~�U��D/�Eۡ"Oԥ�R�ۖ`�nm�%�5r��x�"O�l2ʏ-KJ�ɵĚ9WL�"O���� �7N 0ѓWMR���"O^31��>94��ReK4 ��Er"O���6��9	��6e�C�� �"O��	�M��3�9�#�[���w"O�L�e�x:�e��(٩F�蹡"O&�Q"�4�����;Y�txc�"O��p�"'C(����M��"O8��@�]����m�
���"O�␇�b��y[@l_<�l�"O��Kp�X�rL-�s-B:6�@�S"O�=Zq�2\�xj�jZ�j0`��f"O*���F�G�������l�"O0D�tK��5C$nq	�C_��yB�NI���ʕA	;7J!ԫ�+�y�i͌1�ܬ��GR�7��,��Ǚ�y�͈�I�4�eX��Q"_��y�*��{�!�,�A �Ś�y�n�!9%T��&/�*��ZXR0���p��!��d�:�г��K�Z��q�q@ՅP�y���T��=7A�Ɇ�Y�f��R/ݹyeF@��^2%G<4�ȓ���"��?��ّ�H.�����`��m�j�3\�^�y �Z��4����DL ��\� Jni�7 
/	��ȓ6vv\��+ޯ	�� �a��
P����#���im�M��퐇�߈l���ȓ2D�93-
�?�8r�.w D��,j��C� 1QJ5�´�H%D����f��m|�"�On�T�[c#"D��	FO�$@d�/O�_A���?D�:�KL�m�A�cN��Y��*D�0Z�,�6$� cDK+}���5D��~J't�(9��DA�f�ȓH8�xr�H�C^���f�%3D�ȓZ���a㔾��$�a[�p�\�ȓ�}�tn��:�����J��gl��ȓXV`�dFՖ'�@9�.�>�����E��a�V�\)l(�uhV�N>s��d��tL����oHl(� �;#'l��%j�3VaG �dе��=~yČ�ȓ6��$�]=/�B%h�GG8��ȓ=�B����MJ �d�@�&l�ȓ4�f 8���_��]�0N"9�(��s(�`rē�p�Q��J�ȓ`��I ª̠7��0! 6զ$��@�L�cM��]�@h�钘m��	��M���#W���D�:|/�/Sׄ���e��@�����R*����J�K����f�H�l�(�F̢d"k^��ȓt!����"F ,́���@�����R
��L��OB��C�L�&(�ȓ����'��+,�f�̪x���L��C	0!��q(VaN6��)��S�? ĥ"!NX�W{⨛���:���"O�k�b�4t�Z�{��!;����"O�yX̎P}��ᧉ�d�8"O��DM[p�,X97���v�����"Of4A��'b�4��5��a�r�w"OTBG�C 6���!�9=��"P"O���$x�r%�ᯑ�n�b���"Ol��Rk��1�#�>&����"O�	���.#(�#�^���[�"O�L��/�i{2Aˇ�I��a3�"O(-b�68�*3��9�|���"O�@Ah�/s��[�N_6��"OR4�`��P��ä�� #@ja"O��!P��(�i�r�;�"O�Ț�Cmbt"$L��z{�a��"O��h��%��P���'\.���"O��zc��.���;%���w0���"O�Pth���F���>�A�u"O"8���X.��R��N:��\y3"O�|hqhL�G�����8f��� �"O�T�&&��;v؀�h[�2��"O��b"��H�X@��`K9b&ĝ��"O��B���l�����4?}�H�"O���v��7K�`5����bfP���"O
����6�s���n:���5"O�Ɋ儝4{:R�YbĎE̰�Q"O�Rj�� g�%wڱ&2�)"O��s%�r��!���ݚ:6���"O�cfi�"�!I���}rШ�"O.	���yC��b6+!���*�"O�X� �T���I�0�P���"O�eJF�U�\>D�V	W�"�j�`"OX�2o���.<�A�
�6I�8;"O ����E�ȅF&[Gx]�r"O�	�D^}(j�?3z���"Op}��ÖT���x��]3)n��p"O�Ej�i9NcT@p��M�E�r"O̡
�L9E��y��%I�z�)"O��qp8�e���>y���"O��7	W��Cs��v���"O�K���/�@���g��
^R�!P"O�P	��H� U)�F�@�Q"O�k���5!
P�s�G־��"O�Jb��+[%T��䅞F��ղ%"O�ī2��)'<4����%����6"O�8�q-��P���S�	'yr�!�"O�hJ��J��4۳I?w�L`�"Oȹ��⍔zz	��gg�2��"O(]r�\#};>,�AG(k�����"O>���;L�$�ă��.��"O�1��5bRJİ5Â�r�s"O `���Ce��B��&S�p�B"O0E�^�-�0Ph`��*Z����"O��Ҷ
]�X���5hO����"O�J/\;u,F��B�� ;��+u"O��[1��
0�Q�Y4kԛ<D��@�M]��T��wŵ`fIh�J:D��X�V���9`���o:94�=D��Z�N�z��dBt*�v�XHK��?D�,JA�<c2>�{0�Z� h��<D���4jЙ�.��$�?D�y�+.D���̿56����ɀ(Ab~X@�+'D�dL*��6MB�(JJ���%D�������`���JV}�a �*$D�� �!W,]+5Gj�3�Z":N8� "O�e���H� l�=A*-S&"O2��%:Rձ �րo>8�b�"OBD� �?_q���3d˖\�>u��"O>�@��S���'$Id���"O��B����y�!�J�\���ؤ"O(=�%Oަt��5.�C����e"O Ypq�D�c�^�PE�O�(߶��"O��
̉!��ϑ"��=t"O0����E�Z��t�'��R�ya$"O����cΟ+�@rw'�>z����e"O��c�\4Tb<�ÏT�fS��"O�L�o0�q��T���#"OM��A�J�$ٛ�)�{��tړ"O��ae�W�E)��k��*��%Ó"O��e�\�{�Bd{��K>���9�"Oh�p�e_���:1�K�`����P"ON��l�I�Ј9�l�I~�E�"O�����^�?�f����֟u� Q�"Ob�9�GSbLQ�*E�6gTmd"O�E9�!N�*8��k���n�H��"OP1���P�U��!�E��$VR�R"O@ux�!�p��'kK�iHD"O���#w��·l��
0|93`"OD�� lO� �	ǅF�VDXcu"O����%oD�����#",�5"On�����<���Q�f�1?谥h�"Oڸ�� �5�"��
���M!t"O<tA��$	��k�d�X��l�P"O�i��$W�Z���eɰ�~)y�"O��D��C�T�ՂSrx 0"O��ƪ1d�b�pQ��<|>�!E"O�x�R�L>4|���h�	ƀ=i�"O� R%Α�<�7�țE��(�""O���D4�)q-͂. ţU"O��(�n�)���"偃>6�@B�"OHy�g�:q�᠅1g�"O������"��Ec��,i��<*C"ORj�d��	@����X�Sf�0��"Ovh�K�s����"�O�s���""Odi���4�. �5h[�l¬zA"O|�bŪ?;�UB���~@(��"O���s�0<dHA�ǐ��D�E"O|� �"	>���`MH���u�"O��B%.�.B����A� �����"O��sń����h��%�L�)E"Ox�����i��y��Y�:��f"O�E�$�[�:��aŀ}�H"O��
VDɇE�} �<~�"�h�"O����m�,`���3Z�r�r��"OlQK��ھ62a	�c������y�ѫ}�l�E�ŕtR��Z�[��y��K:�A�Ã�r~&|AƮ�2�y�"�u�ĉ��3/�K�)��y�EK�0GziY /ʳ SPA���&�yR`�ua�TS'�֍g����#n[��y��ǹk�r4��F�'f��PČD��y2h��p�t5�C��]�~�CG��y"��*I̥�rn,Mi��ꦎ�y�I�aB�+���:7�� �Z��y�k���E2&�y����BE��y�+�\r�+ŤG��q��$���yRi�cxH
 dګB���y4�ǟ�y�ǔvK��x7c��7-ܽ�	���y
� �ň�'�3/+ŋG��o� t ""O��dC"0� ��6%I�}�IA�"Oޤ2��׉cX2�ÄUu�6e�"O~�s��Q?�(�`�c�UJZ��D"O�����c�Ĕ�h�p#�"O8��w$�4wЕ��)�E�B�e"O���G2"�fp"�@%Ʉ��"O �Ag�.�t(�!h�%6h�x��"O�H��sHư��I��1�b �e"O�]��H��~�h��#VK~y�b"Ob-����^��A�@�1�Mx$"O
E���Flh|k��[ T%���"O¸��Ί �49 cA�
v�>l��"O��Qv+\1/�$��b�-۰��S"OB<ʗ'� �� �#����h��"O�%�����A�f��$�6"OaK�.�;RB6i�4 #��	�'"O����刬DD"`yCaעU-��h&�'+�d>�D�$�vY�):NQ2`�4L��Oڢ=���г`X(=Y�Y�.�@��3"OZ�	O��>��Lb�M/s��"O�D!Ҋ��B_����L��Q�P7O��=)e�=ʓ)n>!pD�ǆ=d�	I�Ű.���\d6S1n�
s�p��S�\�ȓ��p$Q�.S,H:��;X	laGx��)�A���rSU"5�>����PaI�<!�`Q�DE�'��"���� ��[x�pDxR*�.<���H��𞔒 ��y �HSN�O X�BA�A=�(Op��$�ϒ�P4`џ<�(�T07I!�>Wo�ēTfӡ����@�^:!�A�)H����N$����xB!��"?6v��M1)M��b� #�B��'�"�ӥkA L���Ѐ���*^nB�	�2�.�*G�]�9���r��|%B䉇[e�s�@VR�C��?��B�	 
\�q���͇>oZ��l�Oh�B�6lst�Ff��,����r�� @}X�G{��9O�q��K��co�����C�6aˁO8��(K� ��� ͭ��|@�.�����hO���h.M*g�Ω���ܲ�t5+T"O�4�#U
E%E؄_��{�"O�;��ΝWl�;���(��"�"O�� ri�f�]ˆց%q`|�"O2�$!�?C���W�μ(ZXY�R"ObU(AE��6��=1H;	<h�S�"O���`�@�$G��9��Y +�։�=iۓc�����c��	s���G�xv���&.���`��<��PH�e�LiB�	Ȣ�͏�	���c�O�t���������ɀB�i��o��jp����<���ʰ?Awoܘf?n�[SEӉ֐
�E;D�4#EC�-gKlbD�()z��x��9O7m;�ɲ^Q��G�E�}�TeiB�F��B��M����'��O a���|o.�{�P�lJ^\���H���	f�;����y�TT����"�!�D؍	L��h���g]��5mı4M�p�'�'��	!�(�jЁ{����F��~@`��ȓ7���aE�(;Tj1S%!�N[�M��]�l�;C�W�F��-C���g�<��ȓO����іF0�{R����mZ@(<�c��x�x$�Q(�1I���8�NU�'Nў�i�O�ǀG�;���2��/P9v���"O* b����D0�q#��+L6�3��>	˓��� �z��I�oB̓��w�j)��"O��U*��F�J|�@�U�t�<��v"OFM� l�F�f1Aj�.p�$h@�ɩ4�?�p�ͺ'u 9@d ����#X[h<�� W�h��ےI�p��M�T}b�0�S�O� �CBԳ�"���L����'��	��^�;�`z��	&2�hա�yb�)�S����ǥ��p��|歆�l�B�$n�Ac���h)
!��&}�B�=v`ı���=V{X��^.�B�	�TZ��eqb�[����n�hB䉼�t� T�̛8ʌe񧮚�*���*�U(�����6ـz⤈�3J�0��Y�<Tc��РGg�!�'T0^�h��ȓV(��(U��n��pǃѨ<��+����bo#�~	���ů@�V�ȓ������v���@E��6H[����9��@B����`�@cB[[���?�
�4�h�cp��I�I�W���ȓ#��=r�NC%{Ӟ��V��	��m��/^�5M��B.�D료�BP�	�ȓ=D��X�� ����ے`��'	�̆����;&��(AZ�9�
�'e�V��ȓ]�ai7�&D� ãY�j��Ɠ7Q�ER9Q�Fp��ی@)ٴ��$)�O�0��"I�ː��:4�$3R�D{��)٩"M|��ҧ�2O�,�Q/]2U?!�H6		r�w.�<d\v��.Lka|�|��t������6b	�y�F]�D��ib�aȠ8U!'��y�ܘ�$]{�G�}V���%����y��s0!x��/d����L�y��ݙv�hb�G��)С���ʳ�y���$ᘀ3�iǶ�J-��$V7�HO�񤜊(���i-r �d��̮Z�!�DѨ?1���gᔽA7	i��ؑM!�$�
~��p���f!����/3!�����$��֐K���V��X��{����(,(>L�%MX	��A�Rl1Ol�=�|"QjD,M��&��x:$��b�T�'pў�'U���A�? �#G����Ʉȓ$	��gM8&�<=[��=Hr8Ʉ��ʱ1*O�8���a����xMۂ�jH<�Ĉ98�2`2�j�e���iC�<1��ߣU*�9C��4��@�&�Z�<)���n�|LA��H�2���j�\�'�ay��}rt��4Y8:b���R�y�Č�\�u�f���B�M#�'�
��CV�X�� L�^$0��
ד8B����<���1|�����Gjd�"-�
z!�Ç�.� �@#Q�v쓒W���	Ó;���H,`3����"�V��ȓ)GH�W'g�th�P�y(n�>9Kў"~��ܚ��H���#fX�Hrg�^H<I�F�i����EC"��T��Ó� m!�͢F�ȈcS��
J$`	�ɟ�-k�LG{���'�h���Α0
+��1�o�?�9�'�`q;�F���������!Dɬ�
�'�8����N!β�2T��s����	�'��0�<;x+ș1��Q��^e~r�)�'ldШ`"ڙmt����?V�&\��o�`��*�|��H��n�8�ȓ"���PjTǬA wd�����<t�O&ʓ�~R؟�	�H��	ڤO@��"%�􍒸
�B�)� 0�3r�_��h�P+<@�f�A"Oȼ1�D�=�n�R�'R ���"O����A�~�U�4GG�d2q�"O�qH�]�o�z��P��"h�f� �"O�p��F� �֑��4D���"O^����п"[��j3��մ�Ï}��|�(iU�d���L�b���6b��<ZC�	� �9�p �
(��Ҡi]!!X<�<�q�i@�?5���85�9:��؃~H:2LO���yf�/A�" �ЦRg,\Br�.D�,�!`\�.w��:��7Bj��jq��>ى��.S��y0��1D3��[R��O:C�	85��,����D�쉁��5W���D7LO�	�+�(A��ENF�?�����=O���d�ju�]Y­�b��҉
n�!��
k�
��gʦ�0��i!� ���Rq$�6eP�!���?j!�ѥ�\	����).?p@*s
P��!�\�%�C�l�5)F�2�"U�}�!��z����TL��d%d$��`\L~!��@&_�RDR�*�?l,1��S�@H!�ܮin$����e��D�R㒮.�!�d��`���x0��l�ҝC�=g�!�$�arz�T�ƍxI�I��>g�!�$ބI��z]����`�d
\�!��ʨ4(Ѥ��v�x��S*:�!�D�#f��8Q5�@�w��c��"�!�d�'f�X��A�X�Y�\x)b��5�!�����S�,�'`L0U!4���y�!�d
Ry�q�����'!xQjV�?O^!�$Äd�i�� ڣ �|��A	W!��Rkq����&�i݄�ДkD64C!��X��0=r �ܰY�n �iT�[:!�d�,u��1E�Kw�����뇩2!�P���+V��0MQ�ͩ%�߾2!�ę)�u��ө��͑�Ș�d!���H\;\�c����I��9�!�#-N�,�e�;\nC��) �!�R�S�X&	Y_�X�'�C�&�!�$ڟx0�C���`H*�HwdM�d�!��?N�(�CI��`/��[9�	�'FxY`����:�Pp���� >�b	�'u� �E�Wǎ�Jc�����K�'��x��ۥ	�ԗ$V1�eDi�<9p�º&��h��6&����f�<�6ƑC��ԉRoA�%����XJ�<���%N:XTh�J��d�a���I�<a��^<+l���O��+���a��MH�<A#@3]}:9�U�iD��6�h�<yR�-d�.	�����\��K�<�fF������F��<�1��oi�M����"� �$�	P��Le�F!m�l��Θe��4S�j0D��XmC=HG~�Voֽ���)�%D�X"��z��,ӧ
�c5@��«>D���E�7G���ԲyX��©(D�s�m�#B�Ԁ���z����h*D�0y����qC�\,J�z��T�(D��(C	�)il��K��t�~THp�+D�82&�K�~J��Eϼ@�Z�;0
(D�T�n�$?9�y�G����d1�M)D�L��/��3��$�ݯ+ʄ�8��$D�\�)��̈B��bT,��� D�pC�oNlD�'��Yl�`!E-D���ӫϟX)k�F^	7�L�1�6D�� f�Ұ���~h�7�ʤ Y��ѥ"O$��h�&4ʈu3�a�>>N>�X�"Ou`Ǝ�Mwꨣ�o@1�IB"O: b�c\$\�����E�l��"O�-��e$\U���I._���"O�M��@0X1���,=]6 ��E"O�瓔7��b+T�>ؕi�"O~l8� �`0��A& ;��"'"O2*�(Z=tH���/(���"O�@ �i��)�L�F�֨T���J$"O�� s-� cv�� �2t���"O x�냶F�� �%��+3�3�"O�i�&�N;p"n-�p�R�P��"O��Å)?��0B蛢	ެ:0"OB	��i�2y�UZ樎�]�m�%"Op�(��]2p�,�Ze�V?�D�t"O�XI���H?��'�MHv�`1"O���+R�%�(��)�*h;�H�"O�mq����8`�g�X	N�It"O>���x�8ebJ�Y���"O�MV���9{���C�+�,�4"O�(�AgV	b��r�N���ق"O��D&ٙ|m¡#F-�2��I�"OR����e�ȼ5��Cל*"O�|b�*�3#+TH�s
G@����4"O�-�˖g�Pl#��̄_ت̠&Ϝ"1��T���Y��b2���_��� �� �c)j]�U� D�|bu�W?�S�dy
��=?�3&�����-[�<J_���-$XfHS��'4<��$�Lyb#ߜnA���OQ0\h�,Z���NT>@P�l:,OԍY�K��B��A�BH3D�D ��d�3E�H8�]��:�K��3��\��uv�$R�C$u6 ��'SDe���D_��5l
}�4��`�(�<9B,O�����㟢�4H��'U
lHB�۸.f�� j�h�!O���&.׀$�d�8��B�/�4����:o�xpҭ�2�<���d�|�$?�����Dm����!�29D�%�d9,O�1g�C>az�sbIڲ�?��%-F1�#���P�h�	����p�'�EQЮV�3�ؐ�C�N����+O̬jc�N�*m+篎�uT������]�D�d���ٶa�D0A��Ƙ<�x� fOƙ����)h�XĀU&ĖSm*{���}Q*��f�XdBh!�f�2��ϸ'6�5cc'Ħ.�|��g� � �@��T6�9KG�9 n��F�]�w�B,����WvDx��B�hn�)S�n$lO�}yF�]�. �+ �/�E��I%v�P8���vC\����'c]�)��HR��\ۚE�a�6�!�dQ& ��IR�D� Q��t���C��� B�
PG�T�]��>{��>��gh��)]�|y�'@�o�4����/D�PģG�����z�p%Zt��G7n�qP���'�ףA����qO" �� �.�V���f�)p �Q��'N"����~��8�cHENG�|h��T5�'��>�DH�4ď�&az"� � ���7�4)��	W���<��B8l6IrO��
����2pF´�s -CV9�͑�;�!�D8C����Ô��� �$,��R',:�a2���B���#WH�b�O��P��D�;%K�ԘS6��'�	1]��� ���L�Ҭ[��ؠN�F�-O0R��9�3}���@!��E�|�j�#F���y����!���iBko$H�����|�A�
(p�"���Is�:���dĒT邽��2�j���6�&�Q.O�z�ǇAy�anR�g�NE8"Op1kf�^(���a��C.��q����.��}��B�3樟t�h⤕	Z�C�C��rt"O*-�taM�<�B��DƔ@�,�
����M�� [��Y�ē`�EI�ls���6p�VY�7	$D�k`�L
	N\r�M�b�K5%/D���c	�>� Ux�کD���B�f-�Oؤ� �S�? ��
�)�#r�E�2'�FӺU�d/"��,7Aۤ�p>�d�&$i�ra�W1V�5���i�'����FH��\Q�T�,�~��N��2��J̉_7�q��lF�yR���q�qY'�\ ��U�Ѥ��' F���Ha�D!;8*�uAa��̒h�3��>�y"OC�=��a�s M(�0��Ӭ�X�6��a�#l�g�D�R� a@�ɨ""�P�G! �!�$��	��YE�ڔe6 P�#E�,}�!��Ҭv���HL�@/>@deU��!��KX��(�`� wd㓣�)�!򤃶EB�9��ipt��ׂ�$y�!�ʮ17�9�vNR� �(�ʴ͘&�!��.	��+dP�ߔ���N�'t�!�d�!f�z�FZ%9��%)��	eE!�N5q�ъ�k��lL~���ڥ!�:�l�s@��
V8�S�b�oV!��ǯl��qt�BKĔC ضK�!�d
�	V�,>�, P��pa!��#e��X#a��M~"�M�>=l!�d$hw�c&kɬ"n�y� �:c{!��_�U�$ɻ3GW3���+P~f!�d��=9`Y;��A�<,�<6cΑI]!�dA=<�n�h���/<EY�B�1<!�K�:����曈5	H���ϝ�!�J6g�``b��D�X�E�'��+�!�D��
�\�K
i���g�̭E�!�(T,���MɵZ�b1�1k~!���F��*�k
4��ЋZ�3!�
�:�Nu��CR�|Ĳ�"	� )!��:b�#�	�|�� ���d�!�$�UD�#j��y�^�(cG��P�!�D� �1R�1����qmC.f�!�d��}����Z=1�2]�`L˓u�!�=V�F��$�sw0�����4<X!��T�0a�!�QK�h{J^�hA!�3m�D9����]�(� ,3&!�$I�/���q)�Nd�Q�cG�(!�A�H'��s̓+}f�\C�D��]h!�}�j|[A�V�$A���%�ʖ2!�_&_<t���xO�0��'�!��$��q��a�9\)�l��n�x�!�B�;@e*��DD֜�E,�7K�!�$�3n�zf���'�"�l��$�!�$�WȞ��t́��Y!$���X�!��%��ҡ�I>-<��EO�I�!�dV�GKJ�9`�Q^uxs�Ƙs�!�D��n���C��%���0,I0C�əv9�fO�-���0�M��B�I�0��Y�Ó�9�R1(��G+lvC��8J�ds5�38����A�j.�B�	|�9BUL�	�@���4ZB�ɇ���rMԕz�����t@B䉡U:q[�B�^���	Y�,f:B�I�R�С`��<#�իAւ%��C�I?1tqs��΍6� ��m�?9>B䉸E��fG�hD u�AXN�B䉧@���"�P��Mۗh��xq�B�ɵ<�d /�:[5��hb �Pq�C�Iz�8ŨO4[h�%@L�}�C�/� �SF�tD�ܲ&�ϟU:@C�	� 0�T:p�X�#�� ��l
��B�ɐ�
�j���)G^B�� �?H�B�ɀ����Aˊt�X�C�`~B�ɼ )0�#5	��&�.�Kt�́c�HB�)� �Y�U	UI���y��5=�� "O��� &=-����E���~�,i(�"O�T��g�$f�P�q&�_Ȁ��"O�8�ɕ?�ۧ/�}L^D�a"O��ʵ�_�&���Ӂ�ΰ\;����"O���K�)M�Ur֮��(\b1�'� %S'��T�	$1�dC�N�"���`B��&�!�$��.�
�0R����*���E�qOnsWG<�)�)ֲNR�����4d�䃡�!�Py�� $A����,R�u,
ڷ���y2i��/��" gM�jXl0AΆ�yb�	r/��ó�D�" DypI�6�y�� �*�z1��y���]8�y�/��b�4s���
��}@'e���y�e�/h��E��yc����*���y2�[)pB�ٳe�
8:\i�N�6�yҭU;$ɬY����(�#'���y��$[�:;RIN�q�B����2�yb�~��@iA�t����bΖ �y�MϥY2��1���kĴ��1��y��K1V p� Y���q.��y�l�2Y����
�j�`�]��yBw���! �n?yH� ��yBF�LbTvɗ�neFm����=�y2 �7k�B4"���*�8�mD9�yrď,���s��E�+�8��R��yRϕo��y�a��"L�a�E@��y�߀qM cv��$#Ca��3�y�(�������ΖN��*ͫ�y��R�-��ţq/-R8�t�2�y$�'@%l�B��%U��Z5jF�y���	z7Q@�_���<*��;�y�C�D+d�k�f�;X�Rt�	�y�,�Q}@m�"d��h�)#`�yB��[N>�0��h5ځ�� ��yR.҉����ӝ\Z0� ��U��yr�?@:�X��#�N��`�3�y����R��� `c�9*��GbR��yf�G�(�7cZl`��* �y"��o�,UzD���Tol@�� �G�<1#*�n���h�(c��}��Z�<�⊰��A� ^R�����W�<y��:��!�G�\�Fִ��OI�<Y��<R��X���´n������@�<���Y���I�	�)�"�)@/��<�U�U_�dQq��@)sw� �g�S�<y�7H�-8g�J�Hc���a�<�f�7&i:%��`<�ѩ$#�y�<I�'�j\ɂG!�6����Uq�<i�׾A~��j�Rl�Ĳ�	e�<�TC�go�sk������f�<�B$OWt�y"�U,2��L�3 DZ�<�S Շ��26n�+��(��� _�<iM�=l����cI;[��݁R��R�<ak�9wu��t�7j�|�;�H�`�<!�"��Q�|yvN��8v(c� �\�<	��Y��q��FێR���P�G[�<�2�+t6�8!�%��D���[�<є��.O�J����iIl��bF�U�<�U̧,=�=�� �p�|50%�WJ�<��J>5j�����˃1��� O�<)##Q9����ĸG��U�c�XF�<���E.Tprk��"�3��RC�<���ʪ���1R�#i��0"��g�<� ��iS�O:����!�E�0��TJ "O.Q3��	���й�f�%yi�h�"O �2����R�8Ttd�gȈX�"O���>[�*�����g��|�"Oz ���\f��7Ē�7o�|��"O��:�� ^��]
7mI6(!jLh�"O�L 娜'�^tb�,��r����"OV��B�ŀI������ a��Q��"O8\9V&j4�5��p�rAX6"OVu�Ō���/��'u`}��"O
u��N��D8�	���Ua���"O�$�Rƙ�d�b,�"ʌdf~���"OP�3�T?�`��"E,��"O�Z���l�5X1�X�=6 H�"O� x@��d�RQ�V��9HF"Oz�$�A�w��8q��$-Hj�!7"O\ AR ܇!�B 93c��t��"O�3�.�=�"@3T�F0=�$l�"O���
�
�Ix'Ĭv�i��"O6��̯OS���F�
�^X�"O$ C7�\l�W��._�[P"O���v�_�?���+ȹ:>V4ɑ"O(��m@�("<郗�BG����@"O�A+�-��A�T9ytEU�#�F0��"O�9�!�R.m93.�����F"O|<#$k<d��@�n�<� $;�"O��
���;b��=��١"O��Y�%T��H��-�8u���""O��XF^/�Y���D�u�l�*�"O����?lp���B_74r@�"O*��cg*S��]�A/�w�b���"O�`Y���z|�R_5�6,�"O�0�s	��C@�X����+ ʔK�"OlA2�E�st`QAd�
u�X"O(�K7�\6���fC֣91��
�"O� wŒ8N^@3��Z$|5��r"O�c.��{S-:��ʉT�pv"O*p��@�,�D�T�W�i��0�v"OZ`�N�@ ���2��B"O&�8��δ��!�18�|X�"O���p�G752q��甇h��H��"O�U�\$y,`'׵+��D�"O��:Q*�- X=Zf�M�'�h
�"OR�SE�aR1�W�Ɉt�8٠�"O@�
p&�Q0��q�٦��(Kg"O(�z���71F%3J�#�4]Ʌ"O@!z��%M@�f�V��4=��"Oh�P��ղ	ZP����.oP(�e"Ot��n��W@�!��(�zA����"O�N���&�GD��p���y򋕔N%~t�&�/�X(�`���y� �C-��QQ�2���X�D�yr&�c����O�<�,���η�y�'��P�L�b� �"(f�9� �X0�yR���^HR1K�W�"�&��qoW�y�9c(4��7bE�$�b0�Ǥ˳�y�	�jd���ek�BD25x�G���y2 ɛj�r���kW�E������B5�ȓO�bu%� �N��$����6�ȓ����tG� p��!��,+L�ȓ���)2�Ȃh���
�K̨
��0��p�Tx����D�*��� ڐ��>PP���<�(0���Zh��]�8�x%̏�R���J0C�)� �A	�7G�|���Y�XT��"g"O��Ib7z����R�I��4"O���'��`]�d�8#	p���"O0q�4n�,豅c��%Ƭ��a"OH�yꂎx���	�09�zQ�%"O�,[!b�tÜh��y�<��"O��2��8&\�;!-"�n�)�"Ol��4��#�h�;qG06�%�"O<�RQ�C4EО���F@6�΍qU"O|� ��Q:�v�JsOE=<�y�"O��0���V!���	�V@(b"O��(�+�	0�xJ�*	5�("O��;��Ğ�<�螗uI`-j"O�m�0�Q$/�����h�:F,Q�""OpAQ�K�7%0���eNo����!"O�0���J��Ź"�}�ju��"O��9A�ڵU�ޭ��#E�V�H�+�"O�,���߀/2���!����C�"O���婎/��`�� !� A�"O��aQ��ZpQ�.�����"OJ����,g+�MQwn��=:@ȑ"O�Y���6p����mB,0�-Y�"O�p��M�-q�XP�L=A�N4Br"O�(�1&9D�D�[��#�L��"O�$�I��,$�i@TAv���v"O����o_�)�Wʌ;{��a�"Ob�(7�W
>�deqt�
6�!��"O���BV�"cG�F���1��"O*`j�)�����T � ����"O@��
!�pٚ� Tm��tR�"O6}r ��I 
�O��ș+c"OT�3 ��q"��b�^7!�D��"O��BzQf��D�Z5wy��2�"O̰���[)-�:���G0@J��3!"O��jR��uup�#c�T�U.�Q��"O�4��cͻe�6�X���a� �!�B:6?����-F��a��Ʌm�!��3���r.��jP�iGD4�!�$_�Hr�� IQ(�H�ʏ/:�!��C�2�"wLނQK.�P��^n!�yA���$�Ħ[��@��(}N!�.-n���&��W����H�,P)!�dS�L�����-�(U���/J!򤅕%GF�j"kP��>U���H5s!�D�-g�v���,�Q�SA
�'�!�T��q �MtyNa0Ӧ�=`�!��� &�� �eѴW������J�!�-&p�H!&����=C'���!�d �ngz�{���/s�T���F�!�D�P��CeN�r�T"�"�!��6�2�3+N�}�؁��!^]�!��t��q��� ��O�*ue!���mV�0xƯY8��U�#�J�X!�D�PxP8��=x�;eG�(�!��]�^ì,IV��lʺ��%&�x�!�d٧ M�r�:n��0�7OD�'�!�$ف;�J�91!�bˢ��g˖"�!���9U͘t2�@:v�0�+�FX��!�D�[��p�3��tZ�E�����r�!�V��XQq�I:FEb��� �!��ƭ:�� �c#���:���/W�!�I�3�y����q�$���W<Q�!�d�`
�z��Y��j���Ɏ6"�!�Dŀ� )1�B�_��(�DA0�!�� �mP4Ȏؔp�Ì�>j�
	�"O���/ۛ D(��*]*ά��g"O~ I4kܯi`� cg\1R���c"O\�A�G�#Zq�yCɍ�5���0f"O@��@2\Z\�V�ۄUR"=��"OL�zQ�H�S�� kU�x`�ESP"O�}�3
N H�~��XWT�T{�"O��KC��z���ۅ�43�h7"O.pX0Cª]����BH$TD��"O�`c5g�(X&$���֤),��S "O
��VAؒM���CI�]�Ό��"OT���l�,_�z1�fl´)|E""OP�B7� �mo�I��V���܃"O�\(��#Y'�����z,�5�"O�,c��� �"#��9z���"O�+���0#��� ��[p�8�"O9{@�2'EHs�F2pL9d"O��6o�O�ƍQS�	���$"O���"P�<Y�]�Q�ƝD�H0��"On|�4ə,�&,ᡤ�O1$"Ov0!��L�DC�ȕ5/���p"OX�rѧMKd���E_�'��"Olpr�����H�"VK6�	�"O�� Q�A58�P��:�8ٛ�"O�2�A9Ka"�H##�t�
Z�"O�`�0g�.#��Rbᖉkq�"O0�0A�]$DEܐBwk�+[#���3"O8���D��E�t�S�q���S�"O`�z2L"^$bՐt��+4
��"O*��c�ܣP��}��w���Jr"O~�B!�����pH���Hs�"O�\��
��D}�����)mvh��"O��h2n��Xjh�j�e�B�Y+�"O�|9
IM�諰cU�{jV� w"O�D�D�47�0���qC, {"O���q��=Bt�{Q@Ę`=�@��"O����"Zb���Y����x:�i��"OTd�6
�~���-&=+�`�"O����F(n��x�@l��g7���V"ONI������b�Kƪ؁"O�;���@-���)A�m-Z�@�"O�L�#%�
ꆩ�G	O3K�����"O��ɴ)��N"�Jũ�2QbjM�"Ov�v��>12r(10�4tg2*�"O�L�EY(Z(æ��R�]) "O���+�V�8��8�����"O��{��(u�Tx�g�׽*�^��C"O�Q�6�r1Ѱ��p�(�"O�8���7&C�x�`f�>Gz�Mҁ"O�L�C�_�D9��d�)ez�1�"O�=���) ��1�ɖ�G?���T"O:D�@._)nʭC��C�q>����"O�q��h_N���q,�ȗ"O:X{�MXL�ؕ��
j�Y)0"O� �#L�#"��b İ-�e��"O$�C�D�������UTy0�"O\�;�Ga���b���9��)ك"Op\��Ȑ�=��M���4}�pb"O����&�������G��h�j
	]/\�"
��\�$�i�BI)�O���P��'x�2آ�Hɕe&9p�n]�M�9�GK�(��3w� 8`J>!�}�i�=8j��-�1{Ĭ�7A����-�O�X�v!U������#������E�OD	a'b�N���Jٺ>�V�z@鉃
��?���B� 
�]+�NEUi�v� �ɪ	�6`��}����)� h��D4W1&�X��زc�4�ÔY���!��Ɣc�"}�wc��V9: Ir�pIsT�\�<9�N�#��O�>9)�<y���)|���bc c� xȋ���L1���h����3�+�h��0�}��|>�r!BL�
wv�ڄ�D�"�\��(�	"�^����	��Beo��f
5�P
��a���]�4b�4�)�E+|��O�=%��Y�ߌ{��[��L���[bo܅!o���	?E*x��yJ?�	��'�B��H]�^�.��'� ��}J���<ڧ��D�+��i��bJ��Z��zb��=��aF}>Ր�c��Η;@wzH�4c<�ɻ@vxL،}���K�A�x�d�7T���j '���o����?���'�1"K�����	�p2��j?Q"�'�������z� 	��ʑ47��=Zu��~zPM��(а8�c��|�'��B�ʢW�:��u"�8d�+�i�Y����D?��K���W=I�ƅ9��� j��)�逻gf�Ir�U$mXyi��ɢ2f�'la|��o�QE��#Ez�Blaӓ2�O�p+�M��T�j0���
6+���c�OV�O��9W�ɟ��F�9��'τ��"��	zY����hX�%�O�LivR����ēzX�������i��Q:�nl��(�l�|��B�	>��Z����}B�!'�ȇUq�B�;6�s��"�~�[��2=N�B�Iw�J�3�`@21�Ra��@!_�B��>q������L(m<E*r)@�~�C�� ����r`�I���Q�'I���C�I�38��4A�	�
0�g+��8�C�	�+1��1�EB�S 0�*E�xE�B�&_��sp(���8,��ZT�B��!��۱N�3j��,x*���H$D��ڀ�։Z�vaT�=$���ɑ�.D��� NЏ0�HpI�؅��ȩV�*D�|
W��#P�R����;0m�#D��`5�	l%jAQ�T���]kǩ?D��$�puНx�m�2NU��b�2D��ʢm�t�z��PC��i�D�1D��`�MC�`��F�$P�a�N2D�T�Q�νXR �3U��:��gG5D��b8
@�Q�\y@���0D���'ٛ�<a�7�Z��>�I�*O���Ѓ[�F7�  ��Z�H���"O�E[��Y7����W�Ns�K@"O�x�Q዁U��Q��<Tnx<�Q"O����Ոe��4�'�}�(�""O���� )X�PTr��Ǣ.��] �"O�Y�c�FY�̵	�lѧMOʄj3"Op�[d�S�t �P�D�4M�ek"O��A��\� ����"#}VD��s"OvY�]�An���ZVu�@"O�m5G	����M�+t.��"O��B$&4f�\H�Fҫ#��Ô"O���'&�ܠ�����xmYC"O�<�W	�c��X���ӯ^�V=��"Of�ंߡ0� ��`�J�J��d��"O�ԁܷy��X��m̲a���'"O����^I�(qз�!���y���r
\���C2d�"J5��y�S�/�	�r+�5_|Y�'���y¬�'h ��RGF�b}�)[RX �y�n�) ������+~��r2����yb���YP\hq�ᓑ"*Z��aÁ6�y��_�)+��h_�mH#ض�yB�M�I&�cQ&�"7~�P��A$�y2刲*;�Ex$.U�9p�{����yb&�#��U�6*[��"}a7
Ҫ�y
� ~�PŌ;&f�l8���XD�$�!"O�}��aվGc�0Y�ށGB}�"O��3M�&z7�h��`/�`�"O��tm߈B�,�RO���0�"OjL�6�!7jP����� �u"O���tɊ�b&`8b
�����""OT�+�%�j��]I2j��=B��1"O
\`���s, ɲ�Ʌ4h.��Y"O&:¡�%uLp1D�D����"O��A�(J�r�D�� ����e"O����`k�|I�,�w��S�"O|���B F��y�
�c�na�"O���+E-����k0l�(d3w"O���AX��ҩ�j](r �p"O�͋�(վ~-bQ�'oƩKq�"�"O*���{ä(!`ǨP����W"OFY�&h��g����I9N�(���"O�l�@��:���o�}�|�(v"OJ�qC��((� 0ۗ+�	��E��"O�Q��u�d�;K؈�␚�"O�YaD�0���b��ȹd����"O�{�o�z3��d)
���1"O|�t�*o�����ӀH�<��"O�����iR�R��T�p��<k�"O��Ӫ�9&wL,��E�k/��"�"O� ҄��0%�}��&.&A�"O8 ��>>֔ec����$�(�"OJ}�$�_�o�h�Р �5B"OH�Y��EYr�a����T��"Or�xġ��n�z%��q�p��"O$�j�	�.?|&x�����X�*C"O$-��P��X��)n��`�"O�A)��2�f�@�M݌z:>���"O��4ɕR���c�ˌ�1�`�( "O���e���D�^�b`�r��5av"O|<��n��*����픽}�V�0�"O��pdJ�>A}Q�U�jV!B3"O2a0t�	-I�2\˟�~Q�9*T"ON��+�[J<R�k�	��k%"O�h9a�ѓl��Ca+ǒBt|�@"Oxu�T���d�tT�ZF�Ar "Or-Q���;����7��bUB"O>���(�kv�} pf�j���X�"O�Mx�
������ ��@�7"OZ�9���X��\�%�""OD�Y�� 1�f�~ e""OƑ�uG&L���A��y�`�ʃ"O�1�˚�P?�<*�#\��>\)p"O>��Zb_Mb�<ׄ�Ҵ"O� IE�ǜ\���:Abe!����!��ɹ3n p��-��$�\sˉv�!�=3��V��3("`�e	T�!��R�i�M/��P
��U�^�!��^�m� ���D��n��0��ϐ��!�$B�*;\�����Rx{�/��m�!��%1�r� rn��8dث���< �!��
3m-V=VE�vp�V��k�!�č>A����*��p���@d�,P&!�[�l0�b�������I�7Dg!�DŹQ�$}{�g�;Cx���D���B!�ğ=%zbIsF��=E�~��v&�gQ!�_�J����w�����!G 1W=!�DL�] ��w���d�6��u��V�!�d�&z�� P �ʰ����'�!�� �Q&�ߖ'E���A+$9�0�b�"O���&�6c\�烙9p�A�"O�����r������t"O�1��'v��R����+��${"O�,�"�W|ԭBp�,#��,�F"O�D+�D��$�<H�� �2YI�"On		�j�=E��ڂ����ؓ�"O�5�`��l�� '�_��}ɲ"O&)�!ψ=�814��Fņ�p�"O�=�I�#(����Í�%��C"O��*��
Yȓ�X�T&x9�W"O� I��#��Ԙ��j�	�)��y��N��K��(�lA�CMq�!�$�/#$p���/��xT��-m�!��]-*Ȩ�1�MH��scO�O�!򄕢wA��A�b�;-���h��!�D��B�xI0��U��,b�!��!��|�2����!=� �Q��Ŋ!���Ur��0��o��!y���E !�D�:8V��>H>���8�E��'4zl8׏,���jcn
�-&���'��j���9]/򤹒�[�(x}�'N�[��ׇ&,is Te���'Z��A���3�A�!� %%L��''0u�P��vy
�Ҫ#��	�'��@ ��PĔ�17���I7��+
�'|�	� băI��8�C�ߣEk���'�p�dJQ�=��1�#�ŗKo�ĸ�'�^)a��IҨU�썰H�x}��'a�Yr�/�E��Rtk� =�4P�
�'&���(L)l�ι��)�/�v�		�'F�	`u�1V�AZg��eB4)�	�'���$��0	29���7'J2�'r�(�t���8��J�۰5�x��'�����̑�%?�M�m�f�H��'���;�MӰmX����̃�^(�H�'����>�l)�J�Q�LI�
�'Di�'LG�R�,��I�L��,0
�'C���hS��jЀ�-90 b�'�Php	�9~x��y�Ω��'�P(��]�.���cI`��
�'/|i"fd� b�����ͩUr�Q�'�T�H�oQ%m�bQa�fޒTi�k
�'̺�+e��#t��*P J3K_�ݹ	�'=X��7��� 0���Ũ��'m�5�[�m���S�� <�Vh��'��T!ԑzGJ���j�4#��i�'/�}�Q��W��xç�$q�;�'����K�Mlx���2VK�	�'��}�F��M)�I��]Rߨp �'5~�sAǓ�w2� J�!<J�� 
�'��K�FH/�`p�=:��H	�'��a �ϻ	���VE3,@R�a�'L< ���f��*M�3�`�'�ƈ�Gˊ�>:�Z�e�ʐ�z�'�ĭK�$L�=��2�@��8��'��m;�bM����z�腩���'�\;T ߆c��� M��B9;
�'w��ZԌ+qg�p�ճ7Bn!2�'�P])���:P��͈�
��/^X��'z���n�.6��L�[96��'+�1a�A��`|�bt��}]0�c�'����i@D��UY�M:}�T#�'�V�Ҷ���\��`R���	p+ژ���� $	�a��.z�M`���8r�D�`"O"Xp�A:-t]� �H6s�č�"O0Q��e��n �@떢���t}�"O�@��M�t���ʬy�Pd"O��d�̓,��|#��"�( s"O���7�B2
��d���>���q"O^�9P��;6T�1F�?��"OM p�\�@#L�뱫�S��1"Oh����B0Zx��$!�b��=�0"O$h�4쀓(}���F�L(P��<�q"O��K�A��ܽ��J�#y���v"O����ց���g���DF�H�"O�VFeTTɧ� T^,�ŇS�<�D�*Hs9� �R:a�9�%E�<y&EY�7�*,�Ǣ�5o�����}�<A��d5��`@�_X�,�a(�P�<��gǻ]�0Q4�E4O���A]K�<y�.�4�ASc�M�Z�M��%~�<�3 T�KĂ<�Bo܈qrM#���D�<�q(�8�9I��Jd����~�<�����q�"�L� U1�{�<Q�]���1���q�`���L�<Y4�4;΢�90��";<W+O�<�$J���p��f�B�0#��N�<�a�S)   ��   	    $#  .  �8  �C  �O  �Y  _`  �f  �n  Kw  ؁  I�  ��  ϗ  �  [�  ��  
�  N�  ��  ��  �  X�  ��  ��  #�  d�  ��  ��  /�  v |	 � � 5 # �) W0 8 �> �D .K :R �X �^  e �l  `� u�	����Zv)A�'ld\�0�Kz+6�D�/g�2T ���OĴ���[��?YV̒'�?��]O+�e@�`�L�w���|f�����}*@����"<��T9�e�nY�MA��޳	3��	��:Xv=��gP 8�:<H��cQ��4t�6��0~�k$׬ 0���{������mڋUO&Q���$j�)�%�'�>UT�S"*�� �V)�.R��	e��?:��Q��i��'�B�'�2�'�^�f	�XVV��3&��3V
ep�'�2�eӰ\ꀩ�<I��A*������?���W7�ѵEͦ�t���p�����?��i�R�'���'�$�]wA���ǭ ����F1q$ε���&m:�3��*Aj��w���+AoQ� �tFA�H@ZI@�D@�X��iS�^6n�BX�'
�D1�d���[��@�O�z""?������6� �#����:�z �'r�'8��'�R�'�S>	�;/�d���];E�f��CD�"_�ة�	��Mkv�i7�6M�=�I��MJ��$U�%؈v_ج���!B=:`	a��c؉s�a��5���?Y*Oh�+T��, t��qLI�q/8�y��
� ]E:̳�.���Ҕ��]�T� B���<B��h��X	&SJ��G�U�ߴ���On�����׫R,�`��@������/q�:T�P[v��z���Q�. ��Y%EX�� �'��Qi޴���aەiIiw�{udH4-C-AC�1�&�P2p�b\��mfӖ`lڪ�MSuH8\0X�+$#��Qי�{��V'��>��0f!�'M��ɪ�>hu��S���`}n���M��iiNtC����<��dJ��(�-��V�\�t�b�� �rS�M�1h7��0YL|���lc:�I¡C����(�	�S1Za�G��1qb�j���($\�=�	v���?���?I��i�R�'�B�c�@������
�����r�'R�&y�"�'�Ք!�ݣh>�\К��h���:$�U�z�P�N��|�4������5(@�7ʓ)��E�P���F��{b�:�M�χ�@V��k��T���Q%C�m��V���(O�i�V�HZ.O,R�R�<��b䈗$!�\�i��'�B�'��'��'�����B"`��*��%��I�,�ᥥ�$��?#��]Z�'\�	�?]R��|�q�'bL�TLL�)��� ���/"��J���򤒛ɂ�l�\�*�w��\�ÏV�����)�℺��?y�)"�M��O�tҊm�gs���?}pv�ܗO�r�3DJ�Ќ$AF$�e~B��/=~�HË1[��j��#>dԔ�G/Q�v��ͣT�d�2%���pW��O��n���H��S�u,�1Z�%�.m�ޘ9�E�ZB�O��$�O�D8�'U��ˇ�ؑ*F�l��Oܱ �V�E@|�N�mU̧3������#����&3��E1�4�?a��?��́�A@=
���?9���?y�w��S#ɧ��[Q+�<P��pR/Op�D�9`����D�#��1El�KHv�X?oԩ�R�ыk���m��7������%�3�iEG
��T�l�J��ݾ+�x+��i1��^��m�I�?����pE�Ő"%�5�����.������hO?I���	yS��2�$I�8Z��/�Dy�$v�2Lm�J�i>a��myr��,M6����G���̺
]Za#�@�>���?a*O$ʧ��ĮV<3Y^�X�N6g��؆��XMz�cR�d@c���Z��y��Fdf�@R���M�n2���/s��mx2@��Z��G��![�iC$�]��O
�A� ����	���$[�N�-�bAj�uGz���N5d�1`��k>�<�%`�{Ҏ���O��$.�O���"�5{^nPg�#3��K��|�lp��xn�`yb�f�7m�OF����3�hP �@?#��5�r-V�M:���O@a���Ox���Oj`x���:�H�рkY�-(�����LzP(/&"gZ�q4�S�y���$�A�����F8��ɲ�I���WCD$au�u��I�+��%@aN�IRD�+Ձ׌�z�O@�+��'$t7M�զ��	7�
� ����I
F3<PJ�'ϛ��OX�O��iوnI\DH��
�Lu�x�2��D�y��'�I�M3�o��:&�ąWe}�����}����'6���t^�$c��� ~�\ʓ���i���	�;2*%�0�Ĝ4ȲcԾt2�'B`}i�GS�y*�	��?*]�}� V�N�N �t��0T���@2j�����/X��1�bb(|�p��+_�~���\"*Hʗ��L�0#�$n� �90�8X-n�ƒ�D�s��O��l�+��'ИOވ�a F�bj�Y�$�B�'���H>	�����?!���3_�(���JٛU^�8#��efG~��O�7�O�5m͟���ʗ�y������G����F�ӹ�M����?����4��G�,�?Y���?Y���y����a{�`2�E#J��!�V��n���p�����V��,r�*aP�[>p��L$�|-��BҶ:����Ʈ�.�^Q QN�Xa��ʐ�[l��q���U����Uʠ��!��hmBXiR�`-
6�VEy"�J�?I����?��HQ��n_�7�.��%d�0�H�J>a������Xi�	�7�
2���bv/�XR�ɲ�Mc"�i��'��D�O�剳Q�Duqv��#1t*&		���!q�^��MS��?A�����|J�O|&y�a�WEs����(˥M1.�#w��q��Xw �O�`��d�'��q���<w��knN�j��`�� �]m��:�f�4!��ܢ]~re{SODr�'h��Z4�̰H\؁ɳ�ދV\�H�P�!�?��i�T"=Y���K�̱��4]�ȫ��Z�Vor�|��'|�	�)v%�$@.oV*�"Lb߀Q�I��M��E���|Ӏ˧e�T0�$�i�r5O�u(fM�?�ؑ��*��P��'��	ݟ��I�|+BFj�T�Q�N)LO�!ݴ� ,�b�D�|3VX
��' ��'r�\�� ߑ$�إ����/��1���2u�H'·�={��@�E����Y���Μ�2	o�`�'���C�+|a6A�M�X�l4�H>9��9�I�K�R��O�~\�]�`RV���d ѦE�V!�%�89b��79 -��O��M�*O�0c%*����������O�8����'ɨ�Y�B-�m�4͛�u�vxt�'H��s�d�[v�ˈm�F,X����F�'��iF����Y�.E����2�էD��+V�����A�_iV��`ޮ?�2�+�=n�0(��E�4���F�M~"l̥�?���h�F�/k`
�.0قM����:d@�C�sM D��U�C�D	�`�G*D#<�O޹DzR�	�NA��K��<�n�
�mA�Y�"7��OB�	�����'�?��?(OV��W�>W��E�WO��{l6�ACHmmpd��D�����'��F��|:�d�O�<���φu��鱵����D�ɇCC�:l.�Y��S�Rxi��)Vj���:w� �A2�R4N9�ٺ�R?a٪�o���d�X���O	�3�+f��m`%Z�j#����ڣyˈ�d�O���?a��䝟l�f�@�$�	@�].�����<i��i.7��O��mB���OM�S�{+5�Ue\)��`'ѢS���RjU�]�ܵ��ԟ��I��t�_w|"�'��i��o4�D��FҴ0x>(�5�VFk�dp�����;�`��La�-���ǝ�l������kش��I��"�LF�U�lr�8aB�(���)�qf�aE`�T��� �����G�Uɲ�R�F�bd�U�'v|6M�v�'��<Г�O�8ǎL	�@�F]����%D����I
�H K��F��Z�E6�D�����	xyb.�`�7m�O����2� �Z��b�"R�����$�O� 9S��O���O0�j�F����{��� ��	�d��,�f�W�~A�A�cݪS�@�Q��'�$(
��:$���5D�K�"���/�t���@�B�s�T���xb$�L�'D ̠�(����v�z�$	;$�y�T�2FV�	�G>�bʓ�?�ʟL�}��:�FѶ{�x���-�����I�M�4JU>jiP��6��hc��z���o��6U����Ɩ�xt,x�	��ؗO�E�0�'�.�q&EƁMc �j�M��n��ahP�'22g��/�\��h�,��(p'�K�w��b�jE�Y��ӰG�f�p�̷Go��"h��	���F�:�*�,d3H��n�8*c����(`���O����ǛXV|��A4�u�O�� �'�����@Y�o��J��PP��B�$�k%Mi�<ٶA6�J%�<q)R��b�'D�6�'ߒ#=�G�EN�q�1hҪ(�~\��ցu=���'UB�'52P1��$���'1R�'��n��v�< �iζtK�@�r��z��<Z�H�>�,����L�&ʬ<�%�i��~���'��|�2�͖U �y�2CD�f]����O ��W�ӪF���E�ޘOc�t %��X?��I̧K��[�	��x�t����M;VY�� �c�O<��1&�|*E�&M���~I�|�!'m�<��
�z��h���U]�� ���jy�O*��|�����!x���T�(�M�S���
%>i��@�#�Z���O����O�̮��?����l�� �#F�Y�!�θ'���H]r!�d��U���b�*�#Y����I�G�k����"UNE�c�,��)D�&hH�n��e��$���~�џ|��M�dU�,C��H��F�Z���>5����O0��4�Ic�O��еEĬk	h1�k���'$����G9�x"�M�xo�*M>��i��[�\��ߏ��i�O�q�A|F5:�� F���"���O8���<!�v���OZ瓋! }r�
V�fQSԎ��k��h��E=c��f'�(n���2"�]�'�JUJE�+��]��Ad|Y��F��#�*�;��QX���SAџ����O4��-?�"��@6.��n�4P�����d������ I���C��Q����9 o}!��$������*�r`a4m��#�����O��W� � R�i]��'��,��A�I�L���]Y��u�qfӧq*
�z��'���&��FdL�d(��:�&�`��2A�F+�ST�l��ǈ��u��B"��)���mL��fB�``�(A��#���{ׄB�n'�4.�(0{���5\x�8��$גgf�W��i4O�O~�lZ�H�L�ӗc���W�D�]�%��k>�FB�ɂV2��j���ڭ����+/��?1�퓄g��4Y�,C�*���s�.�3�MlZџ������ �FS6��!��џ���͟$�; �E�w*Þ #RI�T��1���"��G�r�p�۬Tv���"�\@̧��\�t	��+���yBjA<0%H��]@ҒP0��׿;��+cB�z̧�M�� 	A?a��̽w$�����)I��,bs$�ݟ��'��Q��?���'�^8����{�� ��9O�jQ�"O��0柎Q�,uh %;��`�'ù>i��i>M��fy£D�!�� S���^�,�kקE>^,*d0AeF�c5�'7��'��]Ο����|2���f������M�/����
�?��II6*�NnvA!�L��Y��4���Ey2�U��� t;F��.�]!@�� 88C��W�D���j�P�fȫQn��YSu�I�T�4�Q�ЀKkR	91�ϹK�U���O����O�⟄E�TaΊ �F�;�ڃˊ��r���y�	�=��t����0s�"u(����J��'��	-�TQ�����	7�~�y�B�4G\�� bRU]� �Iڟ�Q4b۟��	�|B ěEO�`��e1K�M���y��� ]��h���F{�0�­�����<�O�9]�Ԁ���# ����6I2���D[�IQ�+Ҽ-�B�B g��w£<A!�ɟLM>�f�AF�����GV�@�@Ӧ�f�<Q�$R�9|�r���9���UJ�f�����*�l�%�Q_T����;Pa$�%�D�`���M����?)��+�i�O�蠧.û	�ҕ���@�tE��0!k�O��_
M�Ƥ�E"G2�X��d(�0�0%��8C+�ʧ<~*�H�fc����tJ�Q��tR�O2��Η"������O�2�<L�YY���+�� ңV��,���ڃ4g:r�J���$ѵ��u�n�m�tD����j��Q�X�PY�	H�Rs ��Iy"�'��)�=1Cc� y֨�"���=�2���f�n�4l�McJ>y�Þk�f�' #�@�Qb�Ѹ^:L����?1��<�
�RJ��?���?I��S;���c�|%���Ǫ|\q���}L��1i�_`�0oڋ{l,�7+�e��c5��(��m���(8�$hQ��P5VYS�*a��D�ou�Ax6e1擄'u&�=�ti����)3\�#���I}�	�� 
j�R��'�b�'��M��nW<�}J��;�"�C1�'�bS���IZ�g��%^�d���$,Hh=Z��+dY��MC�i�'����O2�	Ei������2UW��!W��pzȀs`��d��)��ӟ��	����S����|J����Y��=���bү).|��B�؅�<��@TK!�%����R�<�C��5/fhব���4<�0��O]�z5�D�
mp����.5C&�<isd�1�R�IR�ÏX�A��������	;��?�ņ�N�x�P��c �@P�<y���P�(WA
�2Z��8�\`��4�MI>ّ�D�/����A-����U�Ƥ�.�����ğ��I"T)���Iß��'.�P�#VI6.0�1B�܈(��lk�ץG��3�ڬe9�D��
K���O���3I�{�Ze���1<\mbf��.y �"���	�H1@4��hS��?9t��ӟ���^~bA�4S�(�`�.£o�ҙQ��Z���?iӓz�����o�ob������b� �<���T>�P��H�dA%EC-X=�$�&p~��PybG�5Q{��'`2P>)�AAFLY���0(�|�cd�_��a2e����Ƀ)����GsfRC�W���䙀Bk~h��Ov�k�����Mq�D��>���9�ONQ��d�9��!��C~4ѥP%ZDt�I?	c���3f���j@F�1��R�o5?ᕀ񟈋L>E�t�4+��m��	>GUB��Ҩ�y�ށF�����@<�a�㘁��O��F�$���/��Ԉv�Q�m�,`31Jǆ�?����?��	A�հf��?����?��y��pa��C���i��Sm�枽( C��8(�3���P����A	�N��I0��@d.R
;Q�\�4F�.�L�A�t����G8\b���A	]j̧nlL�ϰ���Ug����O
Bt���'j�@x�$3�3�I�aܲ�{�!D�[��hBb恽>�TC�I�
-A��ٓ�h� � m�˓�����W�	�q(M�wD�=e�*2$H�.H�^ ��l�{���I�|�	Ɵ�]w���'���Ш[���`d�%kS�q*�L�?��ȲF.&)�قd��b���S`��[�"\��$.+@b�s-_<��\�6��W� X����1�>�����yq ��v��lx�����$�*+�$�i�'RD �恒-�����'!&7m
H�'@�|�6��J��ǌV�+@���)D��C���*�-q�K<�(t�-�D�æ1��OyR�\�c���'�?�4kU3C(��b�*s��ŀUa�,�?���waʜ���?�OE�X3�`��L̈ݩ��$wւႷ&�V��u����x�@�1*�Z����\�'���A τO� ݘǬ�skz�p%�X&5��r�s/=Y�T��!&�x�'eč�2⛦��<��Y�{DN�)2�I�J�||�ץ�l�J���`�<������S�����5�O���IW/,�i�oW�#U�9B�K.dP���<��"W$�?Q���?�/��qc���O6�T���5����Cb��d�O��DYX'0�(6@�}���`'L̦-�ON��iͰ�z��-������jL]�'��U¤�O-Y:����n�*���޹O����Q%M%�c����O�,J@�'��7�K�M�	J�O�zyICؓ���N� U%��#H>q��䓅O����d�T��݋a�ݢV�N)���I�M���iU�'ST�h�RF�p�в#�d0R��rIE�6m��'s��D�-���'��'���O`��F�I2�j��#N%9��нY�T�#���b(����gܓ1#$X��Y,μ\�2�!8�����L�le��i�(��Ϙ�� &�1!�u������3v��Dpb���'՚�;���Rȟ�'����@�0v�p�CW+~��a�@��y�h# �׫&�Nd+��l}V���f�<�Ƽi^26�5�4�2�i�<��͋>u�`|(sb��,ئ��o���������?����?q�}���OD��r>��i�P;���V&�w��g�QmB�UǗ�7H��Z�ZQ�p�-ղ8ۈ�$A�7�Ș�3	�!=���0��ߢ7/�!y�B����B1�8� ��`ē�WX ���5�	�X��:���A2h��V=`^�!W �Ol��+��O�)��j�4LH�k�/��]��$"O@ 	�*n!��Q
�=B��|ay����<�BO� ��S����� 	px�R�J�23��cG L؟��ɒr�>i�����'3��PD�- ��Mj���Mk���3~5P�� �^l.��V�R'(Pr<�$�t�'�����i
n��E"=7����1f��0�횣7�@A�0��@� S�`�`�|���O �d"?	��ʴF��f��#�D]�(E��Q����B���ٹ�	�B�
t�d�!�O�}���g��h���5����q
!<�X�Ģ<aWl 9ě��'L�Y>Hg�Vϟx����5[����f
����w�ӟ���z�P�cOK�Ob�(�)� /z͠f@	�>�(��O󢴫C��!�dEbSH�s̝Z�OPy�G���X���bQ	D:h37x8��w��|�s�V�Y|�����GӼ@c�/�N~����?��i��"}��O�dtQ�Cebܲ�^!b��!y	�'*qI�d�
r�qq \mdy2����l�OgL홂mY B��' ��'oB�kp�iR��'���L:@&��#�'_r�'�"0���fD!S�V��t#G�q�~|`�Ɇ.��fL�r7&�SD� 1�1��TR�J�~"��PjW�/
��P��ף~Hѡ�؝`�X,@t0f=�d9�C0��{�Oȅ1e��B	ڦr��ũdH��L�7�GyRLN%�?!�'���|b�@�6�(Q��<h��#����l�!�D�APR��
D����Vr�I��HO�	�O\ʓ]�@�K��N�vw�,idM��y��k�"L]Z�c���?1��?!�����d�O��>n怬S�+N�wǪ<s�B�W������5�<x�(q�!�IO5i`�#��	�5����S�'������ܙQ�B��!'�5<;$�C�o��<~l	H���/
��P�	�	U.�jP
��D�K���|��c��O����ɂv�����j�"��x�,�92{NB�ɱI紹")�"��RG�QS*�O�am�^�I����è����]�aKz��b_�\ ����hK�D�OT�	"��O.�D}>I
�r2��LΜR.0��%C`����/B@�Zf��=B�@C(ZxMS��$߯A82a[�̡u�,i`(�fDȉR�V�h�J�'N�7a��B��	�(��	���[�_��&j���'���`���<�l�6d� ��+O>��3�B|[T��4H���A#S�Y�����I �?����6	|8P7�ٛj~T�kbI_8�'n��i��$�Ovʧ)���+�k(浫	F�z�Pl���������?9�
��N���r��Z8i�ߴf�*�'��i�BҶ]��O@�t�8pB��rF���"{*�[2F��
�z"�wӈ`r[w��)IK?)��	�#k�j%�DځR��@)#(?i&���P��4%ˉO�b�O[�A�"p�aB���m$�Ť�6���?�	�d{H����02�|�·�R��hD{��'8�ԘO4^�k�bD�!�t��tk�]:!�P�i,��'�"�&O�A�'I��'R�1�(����"r+r��R(H$�;WLcPN�#�Ǌ�伬`t�Ϥc�1�d�Ox�#I�-��[�cJ0���E�'�*tp�g�G�٨U���51��O�yypD��l����&�9P+��A��'��I�s�T���O��$6��Byph��jG�=��\Ц^�7\�<�ȓB-��;�C F@�i�%�Q�� �'�#=�'�?9)O� �M56O�
��CҶ���I�'��� D�O����O��N��3��?y�O�X��0HΝO��� g�=z�؜�O�c�<\��ɏ�w�X#E��<�џ��S�S�+�DI��Gۍt��8���H�p%�!��*j9�S�zŪ(E� �$f��H��o��<�t /S�����?����'>!	2,<? �S�'O�8�9y��6D��ʰ�̒gm��hqLk.�����.������	[y���Hd�'�?� �.'�|9tB5��ȓR��?��B��e����?�Oغ�Z�
S>?����!� �n68{a!�?S�V���RNČJ���vzџ�C��IAԔ�r�DzU��ؘAR���s�H� �@���GH5	��=D��ϱ�?A����I�	P�ɦ�X�"�.E*� �

��'���'�4���ƨ%�T<H�M�"�XY�~o�F%E�� �kμt�����$(�?�.OXe���Ҧ]�I�\�O�R�i��'�t�cҤٱ8�!7��N�<H���'-R��*I����u
��Q�Pb�GT����'��)ߪ#�!>�D�ia� 4
4�ɂMX�9{� x@�8*�aN&=���zAa�<Eڂ�HfH�'s��XB�o}~⬐��?���h����>� ^�ر�ESX�śÉ*cX�0C�"O�QRR��.��	�GWl4
��"�h���[�o
�=�z��G��H���ǎ|����O����먁�dh�Ol���O��}��Yc��~q�a�&h�#��C���3Nۻ*��4��Z�E�|b>�$��CBm��F 1AN�1@��� @��\�#��̎'���{�&W?Wm@b>&��E�� W6��9@@��;�du�c��d�I�9�h�� �3扁Tݐ0����#\%�$��R,#�C�!f�~h��
P�EX�"�({�˓Oԑ��`�	�}�4#�N��$$��c|�|uK�'A9�	�	ן��I�$+Xw�'O�i�3��H��̋���k�H�!�
�"�L�H�,�$%�p=)!�_ U��[G�Q9N�>����&
&����Q��%�7?\O��(�H�-7�j�:���\�@��
�6��np������dJTg|��re�\s[���c�&�0=���� ,q�"]r5-� �
ps�:��yp�&�'U�ɿ'r~���4���2"E���rSn��`�fG�O<axB⃏�O�`��K�7	�p�"�Z%Q�p�D�'-�h���3<P���4�������D�ax�BU��?q�y��P�Lc.�Y����_~$��t+��y"��{Ε#��KdJE��(���?a��'���a��@�S�Ѓ�G�4��*H>Q��]��?�Gd�a~W>U�SX�� Ɂȗ�kBD���TZC"=�	ȟ�8��W�	�6&��h�v8��S�O0�ô��1��b䌎)fq��O�u�V.�C�긢�)�A�أ}j��A�C�L�0mC�Q����b�x~�چ�?���h���ɹ,�Ra1"�Ǌ>��҆�WXpZB�W}TdI�,ˣ#�.u�� ��_�B�?�f�c�$4��iʭ(t�{q��{\(����Gg���h!��R��?�(O$ �a�.Mڬ�;CMB.H4�!Xpi�PV�h�7�柤��ә2��c>c�� �#�q�$��n߱H��a)�mV`q��pԪ��\��kӍ%��c>c��+��.y�P���䫔@�Oj�$;���	��F{r�Ƨy0qaB*F�qP��C�W L�!���C⁤ZSPM��BG|��-�HO��my�Oo2N�#�;C�4����'@O������`2�$ID��7�˪5� �� "�=ir���M��;d��$ W��[�Ɛ��X�ypX1��(��)8��?��!�@�ɱ���d���Y�o�{��Z�.D�Y��o�
�����8;:��`!'~�'"�1�#���=�\�9bL�	T4)���76 1���`�8P� �
j&����h�'X؉����?���!P�V龴�l�	x��*箊���d4�Old�F�0O��(2 @�S��(%��E{*�"`�'�>ġt$E�H�N Xb��Xah.O@�`Cf���������Oov%z3�'�B�6����U�K�ʄBw+`��JA+G�=��o@ ]�V���/��j�¢%��|�1��!*0��;Z�y;'���
�,՛E9O��h�c�Fh;���b�(���g Z���J$�e�S1G���J�f�ġҢ�I2��=p�^���O��S��o~��޺W���Ժ�]���P;!CB�	!R.9`uU�*���jg/���ܣ=����%a���e�Y�^�P�@��k�@5�I���	O��ؗ�Uǟ�I韠�� �u��'׊1��P�A��@�A^1W��s��U�g�֡��NL+���2��S�?V�tZ�>A�"�������ᕚ*02���\�(�m �R�ݙ�|I��.)Rg� ^r��Q��i�O�6;@�n��`\t���}~"*���?)��hO�	�zoT��������@G	�%c<C�I�>���:�L�|%�A���n/����W�����'���7r�Z�#2J��}�0��Ǌ��6���`�)Y�4-�H�������͟!Xw�2�'�󉗼^,�4��
�1�^�b���<^`�2� ��!�Q��3]�LB6�2{���� r�2���� .����i/0��a�J�����P�RѫЍIV+pH*u�
?"�ODQx��'���A��E �8�6�Ȯtp0pP�'zў�E|b�

Yw���Ue��x9%�"N	&�y��ªw�v9�W���\C&��fȫ���¦���cyi�y���?A�Oz��*��0ղ9�-�,�Di�����a��?��3*j	��������5������ֵ.��1i-Ѱ;�������B��%��H�'��Y!���8)]��i���5�UvJݐ,���J�
B�Pf�R�5���R��I��OD1�0�'L�6M]�ShW���� ��#�x%a���ixt��0?�$P�Y���TJ(e���ɄKx��/O܉��P!W�ސ��R/<���]�И�)Y��MC���?y*�z��V��O�Óg%�IC���&g��T�g�L`<,����S���EÜm �`Ł��RP�2�)߼P��b>�J�N�=�Ե��I��J#lb� ��o��VQ��%,���t��O�
�<`��BA��N6p�1�<����ō/cE��Ɇò��ߦ��-O�O}�3� ���&���T��0��$��ತ"O<�Q��阄�RBE${ԭ	��	��ȟb��*�GJ��ÇE׍$ �h���OH���O:�H�ٖ*���d�OR���O���O&qs�N�.5�Qz�ʌ^� ��#,��y��W(��`�uO�	H~��'b`�=�!-3}�J(���OR�;DV�y���dƌ��-]�"�&!P#DU`]8�͟V�K�aE���I�8�ze꠫�  �j8�p��<}�'����B�V�?�O�牝21ޙ��L3�x��\�hC䉻�X�i�M*ܹ"�H�3]P���v���$�'G�I<\�QVA�/���"$�_lRJ�o�
E����	����ԟ|Z^w�B�'�IZ�k�H���BH�����S�Ur0�8jG%D��փ� X����F��Ԥ�3��D@%I�Ra'E�T��M JE,�l*Ɯ8�{���b�l�3�@=B��p���ˇ #RJ_�d�Xi����u��\P��A	9��7��k�'��!�������w��Pę���8D�hI�)��DR�,˱j���3D�<1�iX�X�H��`��M���?y�OX|=���O�q�L`�aM�o�h(B�hF2x���?���L���e&JA�l!�� �hߛ�9��x3��-o48k��߾K�*ASE�I2 \�ˆ��S�<zd�9h��ͳ����)k�
�{zB1�Ϣ\�#>�� ��4��6��'}QXECԍCY�9Rv�^�<z�!���?I�"�' �'s�	�Nw&��EB�'6����$�}��	'�M�s�i'$�XG�$��*�Z@�ɐ_���	ן,��jyR�'R��'��N�u�����	�o�:�@qC��b���<A����$VU}���N�C��H �HO�������'3�Ɲxr�
gⓧC�@z��,PJ4�	ĎŹ ���ڴ�?�j���y#@�?���r���y�/JŚ��	8�Ī�'W�(PS��i�G��R5O��֟�^w�����+��L��@B'�A�	+8 ppn�� ����O习'c����?�����;�2F�.����AO�<5s�̨W�Z%sj���?y1��
�?q"�'�����M�;ij��=~9���6��QU囁5�2���2R�����O�`#�_���'�R�O���YXUK�������$OfV��I g
���Or�4��O� ��=��s�T��C�
�(Xt����*��I#�˓fIJ�m���?��ܟh��
3[ �����u��']��O5��#��a mEE@4\��!�ņ�LF�Q���'l�]ҟ�̓ �t����M3�]���`S��2U�( �쌧d"�A���y�/"�?a���OG��'��g��;�(�3�bQ"�ܕcf�n�]�S�0�q���4�����RKݳd�4)D �$��ԋ�kJ\ѵ�X�5���P'�x7M�E}�B䟒7M�?M���P�"Y��p挆_�$���7�!�ę-�hĨtF?%��	2��%B���'���'}��'�'4��'�ZcC� ÔU�_�Fa��)X�0Cܴ�?��?	���D�O��d�O��D&[��3&�	��yga���ش�?yO>a��?�O>)�O�f	���*�P�H�%�HQ:ݴ�?����?���J���W���>y*�KC���B+d�$B�g}��'��j�'��d��W����u��'V葑 �,,��'lb�'��'�T�d�'6t��8��$f��C�S z����'���'������O��bh���`�ő(���a��;p������8�uK��U�p��V��e�ȓʍ�B+bfFai�]�X�v���O0h"G����Q�dU.v�¡�ȓq�:�1�� %/���	�c�樇�};�x�&A�)Aw 9a���3K!� D~B�'�2�'��'5���EK�\�ȹ�3�G0C��q�a�T�D�OF���O����O�d�O���O^h9�Ɖ<B���C�k#�b���D�����	ϟ�������Iğ����<�	🠐7�Ċ#2}[P HY?��ɖ.�*�Mk���?���?���?y���?����?�A�Q��b�F�i��x8��'v���'k��'���'7��'^��'B���-F�؜9�jˇ[%	3��,��6-�O���O��$�O����OD���O���QN����H����$��nk׳i��'�R�'���'�b�'���'6|�ҥ1�ꨘ@�)z�FEsªd�l��O����O���O���O ���O�t��g� }(b5����"J�����	柄�	ן����@��������(�#Z�� ��2�6X�B�M#���?����?	���?���?����?����."�~�����{"��������'��';��'��'�B�'���
0{8A[�DP[ܭ��#/��7M�O����O����Ol�d�O���O��$'Y�����dZ:O��E�Q��4 [�n�쟴�	ß0��� �I������Ɂq��ZA��1�H�e�Y2\�b��ܴ�y�'���)��R)�*�0l�/Uu�צ_%Z���*�)����O�i�|��~��8�f (�� N*()3�X.R�R��G�O�6�g����'`- 0z�"WN?)���$�(!��L�oߠY�Un� ��`R)Ff,���u���?ͧ�y��ɏ��(����q�BL F����OpoZ�?z�?	� ����-ߺd$��R�>s�r����'��I�Ԛ)O��$k�p�ILyBN.��x�!6Nx���ł7��Z��&%�A_��i>{6��.6��Q��[��
3=�L�LH�Z'��E{��'���Is'�h����SNݴ���b�("�����y"�'�V6M�OX��|�')\<	@��[�i䅁���q!�'��i��îüx:�Oy�V��l	�`i]w�$F��7]�8��3�[�g�|����'6�I�?�`�d,����Uc�Q�`�')�6�+C��	՟@�S_�T�'^�(��$�j�40�R2�^�` �<���M+�'�>i���A19�`�U���y�U�3A�WWrᣃ"2?q�g܃]����gC����?��L�}���?fs,����C�F�=����?���?	�� ��d�
-O>�n��# ���(}"�#��Ʃ77����&ԧ4�������z��'9��v��O���Ӱ�M۳$6`�Sb8�� B�FY>s_���"&@�<YڴD��3�A����!FS� ���21�X �A�O�Lm+���Դ��E!S��B�I��@ölҸZ}М���@�.y(����=��I(@FW?�@��X�I�!YHFձ��U5���ޝ/�a��RQ��0r��9ح	1#\\<��pF�^��-b��![#L�:�!ɀ� )�ĩ�',���@R�I(��x0���T��͢#�/Alaj�����hM;v,�0AT�����)�:��C�6q7"O�xZv�܎PLR�䗀D�*��"�'�,j�M.� �ˎj
�H���b'�X�J�L�\��C�>ǆ<�7��8��q��̀v"\P3��v8""O�=$2���%� �l�6m�,r�B�B�cp�}��+r�=�҇JQG&���2߾I�^��'[�;0tA`ՃIu�m��؁� �+�#�,��O�D]z����	~�;T�q�OX��Z�QwK�zS����՟����ޟ����l�	̟t��ϟ|���޹�A�Ӂi�6�y�gA�o�
E��
�����?���䓟?��u:`����D�ml��	R��l�c���?��?���?���?q����P�2�Oh��&#N���b�֊H��#-O
��O�O�$�O�u��O�e��KZ�#,h.X� GH��O��D�O��$�O"��O$Q�.�e⓼9��q�(Ṵ�1jM�{"$h��'=|�'<���" ���'��a>;�µ��㜬+�Ie�1ΛVG�W:t����E�$����ƛue�ۥ��?Tnt�b��6�N��V<삀 ����:�N�J� �d�O��Ov�$�O���!���JP��b�V��p���?v˓�?Y���?�M>���?��>^J:bIñ�l��芤|�H�4CK�f��O�$�O�i)�I�O��dHb>���_;F��8	�&��(��ra�%�y�	k��B�=��d݉t���'(�_H���¯V*D!��e�A���O��%����.2ƍ�,ЖnRL�zԩ��	�T�r��߯k�*=��G��]��yQ��$�-�w��-@�W�kE���',�oL `9�[�F1V�Е�Ƴs�zh��u���� G�ۦ.�{dP���H����%L!C E9�n�{T�U�I����-:.&@i� �u8F���Op�d�OR����M��V5p������i�Y�a@!T��JD�m�n�3k��,�\#L?m;ڴ[�lĕ'�|M���$ܬ�!d -�r���N�{R��D�,, �3�M��'�M#3)�lyR"a�`\(p��?(r :%d�6%n�n�̟|�E�ܟ4�)�,O��$|�d|����(:�Y[Ä;�
e�`LFޟH��ɸ:�d! fL��c�~\z�J�([��	��Mk��i	ɧ�d�OR�I,6Ϩe��k�3te��[��*�M��<w�\�	�0��П�Zw���'l���+fin\c#)X�v��x��&	�UK�䖿2�$u�B���G��Q���.T=�EZ��d��<����-#��W(�=�Z�*uŘ�Ά��P�C��E��+b#^�;����3�Fm�*\渁Ȕ&���܄:E���B����4�?!+O@�;�韾4 !�Jf�&��'.��= \��"O^Т(V;r�2��� � �>钷io�T���\�M+��?��49�Н�l�%vĸr���p��'u>�'�'db�'�^!z�i��pd(@�5s���i�U�r��R�z �S�Ҽ@l�Ԁ-�@y��&�ĖP�,��CEW9���mQ7D�e��\[�N9�S����O�� r�'���>�sb�ݤa<�"��U�fqԬ� %D��[��@��,���a�(:ݾ��@=�O���'�.�)��(�nΥ4���O�x0���M����?	*��h �O�7m,���S0&зr�H$;K��E~�@�	�#��*'�����S'A��(�Lz� �*F� '>�k�-Y�'O�Qq��
:M�|� c�>0I�τ\h��/{ �E�xq �(��D�dk��L�~iy�ꍦ�ʐ��O�aV�'�27m�ͦ-��r�O�8`�Ȟ`������^z��Y�*�<�����?� C��T�b!�Q�:�ir�/��M�t�i5�'��N�^N���f���N�:�g��#�����ß���*S��$��ޟ���ğ��I�#��^�fon�1��3'���8�h6���"�zp��)�*��r����H ;��'bH�
�h۲(s�<��ID�N#|�+� ��V�j��b���[�bt����;�ħA������E��ԑ~�h̩`F0V�D��+�)tjJ=�'�Ɖ"��?���'{r�ivD	�BɌd�r�*c�Ȓ�'��@������6�tgp��'W�"=�'�?�-OƉ�	� B�g���p��ND�Wۦ0��� I����I�|�	ן��_w,�'�i��0�K��M�7��%���֫�\ [��՚E�6� �"8�az�o 9Lo����G��Tx��9v��������n	�I�3M,�0=��ņަE�
,��c��U|^u���I�F]�f�|�^���<��������S�c��19cgп6�0��B#YI�<���ȕE��IV�8QK�욥�L���
i�����<�'N22*���O���u�n�� �D!bdnt��+ʳk��]AV�Fϟġ@G���͟� 쉆d4Lۧl�0X�H�xݴ-v�����N�*��eƘY�l1�A�[y�+*��'�X�'�8������n9,!�!�N"`����e�۶�X��Ϛ7}�蠣�_crc��3`)�O<���O��Dv�y0�̅�
 ��9BQ#�	��ʧ�h��T�S�O��y�vǖ?�~J��i�0�Y	��3��dLA�� �Rł(q�!���H��<�'G�2D`tӞ���O��'[�v	��M)��$�tɘ���)-:��A��ߔC����Ӧ�O��5�Ⱦq���ޝ,�O�"q�׀�� cr��L�@e^���O耹�d�h'Z�+�M l�rl�#`�M\��L~ڣ揕
?ftypd�p�A�MM}���?�гi^6�OL"}z�O�2HWF�p� �R>B���CLP���O���<"�xpZgJJ�s��8b��?7!Q�<؍�$v�as�$A"���Pe��	e#D	�6�?����?�!�\�A��T+���?Q��?��e�1.$�Uӄ��D�zD*�21:(s� P=dM*�o�D��A"��JO�S=)�Α�������/B����7'K�}�<z�c�����L�jr���4���O�8�ȶ�J~Bey���sg��A+'��N�	).2�$VQ8���TM�-0 ��$��&�	,&D�� �G6M��̰3쑺?`5�u!������4��O� �$;��0ar�ԶuJ��3d3`�]��.C��?I���?�4��n�O�df>�t�A+	lv�K�R'-1�L`G`W�@ln��"�Z�4X�ųa�Cq��z�`LQ�\��#V�R��ҧ��!�d� ��� :�td�����cLR�$�b�9`�	�'Q���p~��EJ'O��UO5A��[�J؊��2��柀'����䟰�?��q-�pykLl�L�B
�mA�C�ɥ���W�W	{P�(��Ԥ=�P�'�7��O��h�p�hV�i!��'�v�	�@
ƒ@58��
R'��d-F�x�$�O���M�*|��zר�	pA�œ'̓�y�M$�Pr��,���Mϳ��O�Q)�T _𨝱%�9Ni��\z��Bꄾj���k���e�p�2��I;AU��d�O��l������&��:��LEz@k��ԢL����?�����
QW�T��kۃm�|1҆�"�Q�F{�g`�̺" �� �جreO`���*�"	��#��h���iK��'!哾fF)������sHC�hZT1��k��)�H�:�?	��M�?��y*��'�h� ���DE��&LǎoS�ѯOf�K��)�'.�p��㌓���rei*��L�'`��;�����H��-+2L��I/́)&���9mT-*@"O����%�1Bt"Yѕ�U�MX�t����6Ѩ�
��5�C,:Z�(  I�b,lr ��ڟx��ޟ(�%D�=����ğ`����zXwa���XG'�)èZ�8L��s1��8�Hx�O�y qA�A!*@%>c�p0u :@�.��5,�	AJ�bM�ciR�{��Ұe����4�K�GF��yXbNɌ���A�d���靖B&�}H��#ED�'�D,���e��xҬ��i�~��'O�Z�U�Ǡ�y��N�r� RJ�+��a)ĀE��~��6�S�OBZ�0I��^�F�5�� $��e2�CY�1��'
��'-�hp���	���ϧF��o�;�mHQᇾ"<")d�E#`��Dȗ~�v���T �85G[�2��2 gޙ��?S�X��-��	I.;��p�Ɂ�d�6$�?���ę�)���ȧ.�0e@$�x�.�1(!��'EU����<1#�[`������O2a�/�9�IٟLo��_���J�i�F,�q\
6g��{��z�޴0���?a��_�`���Ø�u�[�f	
�&×S����j�4��O�d�v�ӵ�|0��dR�tR@�ƈ�
�8#?ɦ�Q��웊���Bzh` �%ҿC�@�b&'�<�y��^���� F����p?I��O0�B���&}��#B�Ѧy7F��>�W�
��a�|�����(|��d��K$>f�������M�{��O?7mS�Zjt�z� �,+���F(x��^Y$!�#�L�W��Q���L�[���?�*x�3�]���ѕ��z+���ȓ?�b8k#��<�����D�/H��9��co1�Y�� �:)��ȓy�>\�C�� ���1$�xq����S�? �a�2`��K�!��K��|�:"O��p2	�0����A�-�"h�"O��)i�B+.�*��m�|ͨ�"O^�Ѓ͞�8�pzAF@7)�F)��"O*}��������+���B"O �P��ӹG�ٸ�/�+�ZA9"O�%�ցA�6�*�q�oٞ|�4�"O���V�(��k~�Ĩ%"OFx�ӌ�K�xۆ	*Y�J�a�"O��%b�<~��}���h~&H�"O<#��2ԠM�`��X�x�"O, Pˮ,Z���J�@8��"O�����8pn1@+�UeT���"O���GA�:�8h�k�Z;�)�"OLXЧ�ܖT�$z㪅b���6"O4(�GK�
}J�i\?G� m�c"O޸���|u,!`�Q0[��|	�"O�����g�0Q�F�	�|�
4"O*䊗Dup�y�CAd�ܴ�"O�5 �/F�rV�X@'A��U�1"O��!���#f�UK�4h`5"O����lI�-�B��D�ȥ&0�U"O�Ur�d0!f�h�h�Hj�xc"O���X�Q���K%D�5w���"p"Or�SF���c\��,�c"O�T�O
)���b�Ƥ ����"O��@�="H����CU�"O.�Hg�,�R�����nT�"O���΃�^��E�TJ���qT"O)ѵ	\�l���]2r���Jc"O�m��IS�_a���#
2F	.�� "OΠs�W?{fd��)����%�J}�<�
�B�p�*�N&Mn�4����f�<����6,pxpQGew���A �E�<I�k�Xjᢥ`��Т�bG�<��֕V`���C�BS���G�<�aG��)�����M&Q�Zy�W(Ff�<q*�e�2�t*Z�_H�H2&�a�<�P7r����FA*$�|U��Y�'����P��C���jƕM�1 �ޡ*�B�	!*�v�0��J�J6�d3$˘;�j�	�]S\H���퓗Yr��)ЪǱ���9P�/�C�ɠ#���I�l!'E�!�э
�O}��'M�x�CT��HyU-	�����Ę5��4��I5�O"y
�eT�&�Zd�u�A�EcZ�Yf����e�	�'�* ������+Uπ;Q|� ����'�����iك'vt�r@@1J�,s F@�YH!�d>xOV�q���V!j�{���+]7���2d����{���%j����q$�3c̸ 0A�(!�86�҉�O�,��Y3����4�'Zn9�F�'��;��]�1�����N?�J���'���i�� +y>��Q���9.e����'��8�#��Y����2�C�&���'��(R}�$�2jJ��uH�'x�ȳ'J�o'�0��,#���
�'�zQ����_̡p*׬���"�'�V���C�<w@��.ľy����'�@Uzgj/d4dIC�X�yΈ	�'�h`q�	�4)! \�Q傁p�(-��'*��&N��MW�:1�J�h����'�
�����0�<,
&V�x��C�I�z�8:�bS5����d#�	'��C�IZNV�pDh�7I�)Sq��6�B�	/s[d�+T�Ԡ^-������Y�ZB�)� >���O��'p0MC�m�~�E"OR	I��7W�
l2�Lݮb�Z%�d"O���7
s}eQ4�J�q�K�"O���1�6��e�V`P�����C"O�Q�3Aʰ3P�6d�be�6"O��Q���;8>ѣ�E�4д���"O�{�K!TG��k���7� �"O��3�G,@u��虙��t"O��ɖ�A�~�RH���RJ��"O��"4G?��1��^�eW(8@r"O؉	�7t�L����Op]��"O�0𥢅$M�m�7I�j �y��"O�X�v�Q17P��NEL��"O���3C��1�dt�� ���]��"OPh#ŇÐJ��� �N�.J�$=��"OR���*(F�.7��0"O�� G@V5lꄳ�O�?�Z���"OHd�%�	��P���)v|t8�"OdTc�
$I��� �`���a"O����H>s9�!������P%"O>�p���ޕ���Pj����C"O$i
��`���d���ʱj�"O�)򲅓,5
�\�D�T?�J`%"O�}�["v�e$�0b���"O�\�`�p���cR��t���"O0��U�ұX0p�ɐ'�<�2�
�"O \��gO�gQb��vc	an�Y�"OIZ��@�5 ]
�cO4N��h�"O����n���G
8���"ON� 3ő�8�Ei!��p$��g"O� ���>$��]�
����#D�|p��ƃ�L(��K	�i4��3�&?T����R�!�^]�bm�oR(h;F"O�+���P=jUa����H��"O̩�싳l�pK֌޲%3���"O>��@��Z�Դ�QJ]�LG��b"O�TR�ߧWR�1A�@H%9$ٲ�"O|q����_�� K!/����"O��VL�3����BO�J���"O�i1�N����?>�BL��"O:�'"B�8TCY'U�(�c�"O�5c�e[;1δd�����D�4"ODP����S�ܼ�s��%_&�(+�"OdU�6�<S�J,�@!f��Ҵ"O�s�̍�>8��b
��_�D�r"Of�Q��L3���k�����'��I	
�*@1�`�M$���B��W8B䉓N|h�x��Կ+{�}�"��z��#>y���h�FX��F^"{*Ts�.G�M�C䉹�4�!�'��� 8b��$l��dC�(O?i �o��v�^t���?��jt��E�<�d���IK��I`	1��II}�ٰ̊>YG,J�x�� �2ۻ2Д@�Ti XX�,�4)�>��$�6;�T�f,N7���*�,�S�<���z)�H*�L+�5�MH�'�`��B�#;M(��5j�e~�����8c�C�ɐr.БQ�
ð
V]#�C�J�d!�b��������ԴtL��B���pla
N�(�y2K�!��gL��y����8�~BO�8?fa}R늝�4�����L���P
��p>�b�C����%%�R ���ͭ)(�`!�ړ�!��	"�L��	�p��9��5�Q��IN�N�O�-�S�^�i�d�k�g�4=fq�'���X3BΣEG`�B��]�|�ȝЦ*��7&��"~�)� �c�	5�d���LԊ銴
0"O� `&ۊ�h�*�kZJ��P;�OR��4�O�QC�3,�lP4`Q��A�'��"rT��X&ǋ� �0R�_�&b���ȧ��`���S������<�<���)L�@���i?Q����X���	8D9 ��3x�튰�
&��6��{�"qw�>D��zG$�7&rĕ�UǕ84!�]��jw�޶���ƣe�@�{�.�mO���}�(]>ؑAΚ9W	*u*�!��C�I"j�H1��9m[D�0h��[.�5��FM��2�ۆ��<���?��A�w�,O�h ������r1��Z�2�Q �'#l��W�xY��d�T�PDDL��=ɶ���t��y�NAL���NZSx��EKF�xRC)�pL�u�!%4ʓPF�2�O>���+�"ޮ����U�X��tJ�����aa��ȼN���w�gH<a7ᖂzdX��@V�-"0�ɔҦ�B`�>����t�X�� ~lT������b��$����մo�0M��"OF��&C�V�H�0���3w�$A�h��8c(�
e�� on1o�%-�'V�L����D¥X�D@�'DȖ|C�����>ji�}�A~}���d�4��j�b�a�L7/H.�y�@0X�p��&*W�t�����7*��XE�cE��0.�T��O���aaѲS��=���64/�4���G�T�>��7a�
0�(�IS�SH<ad.<@��j�J� ������t?	�O`���k� ���&�l���~�b�܁q��5S3ϔmjᡕEp�<v�\�#Lr= `�Y0R�t%�b�ޭkbd�A����i��Tp�𙟼��>U��5��N�k�(}#��*D�\���Q�	��kM39���ϵ.�&��%����(��.�jx����#O��i�?���y4�*\Ox�BB�.kQ��/_�-�B�Ka�1w9j�r!�H�IV��O� )&���B�b�v�Xq���P��Ɯa�0 ��9di�F�4n�0}��+��D�|o8h����,�yr_t�V"a���NF�t�=�u'� "d!�'��>�I/sPZxrD�G�xo�)��O�	*bC�ɱ*�D��tLT	y�X�W(Ėa�t�I'c�F@�c�:|Oa�) z�b����H�q$���U"O���vi�!.�>̣�¢jr�ii�"O\���'�,/n�!!fe�o(E��"OkKE4dh8cr�rB�];"O.�!%�άH��`�'Կ
��Pq"OD|�0�߹�f�A���#S�u	F"O�,)��
2\4-���,R��"O�  � /+�2+�-_+.����"OƘ��dIXm�i�a�{�"O�tcC�	M��t9��P*��c"ODi	V�D�/	�`��O7�c�"O��j1F@�Eq⋊<���F"OZ��!��4�F���*�h����s"OD�G��)��s�P/0�5@�"Ov���*�)���uf��V"Ol]�cg_�(���bG��-D�����"OB�B���9������"rjѩ"Ot�Wj�R ��S��T�y��"O��rt
�[�l���#Q�)�T��"Oz �v+��>��,�C#04� ���"O2x�UK&j��,0RLY ����"O8vĕ�z~囲��'+�@Й�"O*%��Ïc}���q�]�l�����"O�a	�=0�
�� '�,�b�"O+��C����a��:P�@�C�<�snL'3�k��U?m�����Yg�<�iܻD�V@����(����M`�<Q�eRa@BMR�h؛���2�[�<fҫ!~��C����8#��F|�<q��W�$�`2qd�*��Р�S�<���9������.��]ʒ�P�<y`�۾���KP���;g�O�DV#U���.�@
�����O� �	I�H��aw�O�3o����"O��"�-�R�p�/Ɲ_�@+R"O�X�p+
�>�x�An�Sޕ�"O0(�ĎI+huH�"D�36:�"O�������Nђ4s��3�@�11"O�
Cf���Q�S�CL�U�T"OXAS#(V!x�>�Qr��-GlA��"Oh!����0q6�R��J�4�"�Q"O���F�G^ܑK��Ҋ|ul���"O �@֦��\�X�C��g����"O ]8C�^����$G�d���"O�x��]�a����N��&�|kC"O���r��$��!��g�HF����"ORE��H�h�Gǭ�����"O�l(b������K���1��i��"O�(㦅ظeBru �<PzXTc�"O����j�-�X��;i�.8�'"O�;���{(��r$,�h��t[ "OD![�NB3Q�Ш�/b��A�"OH<[#�I$^��{d��w��`ѱ"O�i2^30ȍ �lsL҄��"O��)cL߬3���c.!���p"Ol�k1�_E&P�m��� Q�0D�Ӧ%�.u�8��&�t�
DJ�!D���q�_��i7K�"f������!D�p�#��P��m�a'�<B��5A�=D�\z�Lԟ� �vK�0�@Y���;D�0
"a1QӪ���&�46��<h5B:D���a�	>JB��W)B4+Vl�c�<D��H�*8L������p0p���;D�����^�ؙj*X%"�`�("
8D��kfgN)L��8����B`���i7D���GN:sr${  �6i�x����5D�*'��!L�
��̚�J�:�
2D���� �p�0C��!W���"�0lO`��1�Z��`e�!bZ`d���1�Ҕ���O�@``��I� �`a#�V�/��틥�W�=� �Ѻ�R�=��`M�+)�|3�eO%ȹh��	d�	�u�>��#�J�;����Ƒn�#>����'r��Y�w�3A���:օ�<�C(B2��:A��S�੢D�]�!��  ���S$8�:��
��<ٕ��J�����I�`����OK�<����y��U�ؼ�Uؑ�A�'�f`�u��;K DS�n۝g��x�OF������y�Ax�@݅o�e�giD9.o͛��	�w��\���A�;󮃊�P��4I�$�"����:a~��T=C�T-z�C̲N(�ŁF�80u������'r�� �O�$\�t@%&B����O>���Q(S½a�DK518�Ц��z��0Q)�;ϴU�-
�I�=�`4'D��!O2�ۖ
P�O>X�%D!0¤��,ӟ-) �� ���<���ík
��5C_�~,�����vEQ#Z>f�	���EQ�\w�n">��I9S ��#��fBBD�
R ��<�"�O�IĴ��d�dXH1r�A�3l��� I\��OfAJ��g�$=��w>b�Z�d��4L���̝ts�(s�y��i>�c�ę�:�]��@X#[� X���ڮZ�h ;��2�I���`�JDB�hȚ'6Tv�O��0��	��aj���-���8Bቕ�M�w�;�&�����
޶y��c��$� /D4p�!�T�:� ��;Y�	�fIT#G�"=2�Iŏs���󤅄w+��fB�~(Z$&�Tn5Z��^(>�&u胪U� �N��R���7��D{R�)v�˃f���lЂ&FTx�����6iC+ڳR'6t��χ�_>>aZp���8�	�jC7|x|i���	�E�9��I�!.6���X۰��a�M���r��P(1O��	��$�b��{�� �����(�k!ÓR��,�2j5qO�TY�M	�Z����A�M+9������|�a֍MZ^L��a1g�x�����M�M��ݴ�?�4��m�&Y㴏�Ӧ�����y��Q���A)Ė"$��G��,=�x�'�;dBm+&H:T�y2��X�n��v"�9_����.Ә+���֋-�2��ŝ H�2��6����O2��"ː�| ��V��Ly"#<O�Ik��A�Xd�|a���&��MXeΛ�]%�A�7 Q��jv�ʤf�X�Q���FW�Q���"랑v�J��FD�f̓�~"�>�.����aİ?0� ��Ú�dMj��ؚs�z�0&�d�5=j��@/]V��!cB�MG�'@��i� R�iSD@�E@�Hܴ��	� s�4`�HڰF	FM�( $�º��0O��H`C�'\��bC�|vt+��D�d}�1&�v�̈�3h7<O����I&#б2$ �4U�|��D�O�el�a�����	S5�]�Ű�'\�&�R}�Z8��	ϓ�~BD�H�䔘1���SS-��	��<jbH��<N��!�uUQ��D�܃fd�[����ڑ[�M�Gݎ�{[إ��O��1O���Oj��jц̢-T8�1NB�@j��ɜ/qB=:�{bF��x!��!��1���T�U.��f��x�@DEB�����1i��|�<���?aB��7`�D�S �N Lh�����<��Eu��I���3sPP|/�P�ZPo��T{�=1���<�3�I�l��c,��6p�����?�"I�F����e'Jɨ��3�Yu�'�0{��=6Uh(��j�WƠ���'��O@=86,խ!�x����JRI3ҹiG���1�,� �8dHY
)�:�x\ckP�I��T�+�  J�,Y5l���y�L̓k,��i�l���U�DA�; �P�V��̪�3a.%@�{B�	�p���!X��AmF��ɻC�R�S��H�'�H�m��Q�f�(%Ee?��yFAQ�d_�gƩ�'[��O�Y�7̌�IrI��N&8�$�x ��?C̩�0(�k��e���>Q��$N�P���[S��$�đ�BH¨ ��$�u�HKfB)j$��'^�>���� x�J���j轁���),��hO���aZ��F���kp�ȧg�h��e�E8ju˕�ɛF��}xR�6�nRn�`� @)�^�B���!F2c<qO~YD}+�^�q��@ag$h�M��J�9�T:�'\�x�G"�Fr	9'I��,�Ux,O�$��H�1��$�cޔ���&�6sC�����v��Arċ2Y��e�bfx��pU�) 
ĥun\�<��@�.�0� �HL�gƤ��ȉ��4��S��I��xw9!��-)���k�c��?�s���Q�ݐBZ�v��1��A�c�'�9ɔ�Iw a�v�˃v�&�M>�r�ۣ6"&���+�l�)ӣ�
��������9=�Z-�ȓ=�N��q Ȍ-v�8Ck\�J������[��r���L��b��%&$*�vY\a�-/4�\qTÄ�T���K	+e x��A�L�I��0a}�%K�Tز`�vGy  �W7��<�rOҶD� �S�>A#�g14< B_H����d�<9¦V)XL��z�H=T��4�"��H�IS�5�&���c�?s��J���I©�J��@#�
"D����W&�mA���h��	�C#��~|��rI�\ЏVZ�g�d�T�� Y�nv�Dt�d�C���Ȁ.�z6"J$�����F�$2�6	�'��uB�X�ڵ�V�vS�5�@�(�]��I�6��4�D�!h���M�B��1D\A�d%�u=iB䉅y�����h�2c�d �G���O��`�5?�X���I"{j�!.ێ1T�tK�(y�a{)�
Cn!��
v"����	3�.�È	�>�8������Oҧ�]��k���zi&+�kx[g�6���=���[;_�"�X�Y�ī�Z�	�_���� �n?|S7�M�">���4���r��/"j������<I3j�&� =k�+��y����5��t#V�cV��f<�٘c�?��<Queͼ �rܑ�E�?h85�3BO�<	&$�=I�T����C�z���Pqm�\�'��(�q�?k|���w蟏p��+%`>$��k3�J�g��q8�m� $?�L�Q@O�v��5xB�-�#Z�	@��Y���]/_�n���c|��3��2����91�z��qKA>uդ�x�j���Uڵeý�qO*�ض�έ��"ճ��t� �|�E�E�v%���G.��!�,����O��� Î$�v���m;a����p9O؀�����8Ab� |��{��8+X��E��a&� ��-<O���͞�.ȈȢC�������=O�h�Ɖ��l�T�;g�Y����	�~��E&V�V8(���9N^��I�U��\}Z�C,»a2D��7l�jB>���3d@"�"K�h�'C&��"�S� ��1�;�]hEmAC<��m�T���<�e&}҂�b�)�,�8a�siá�c6��W�,�a�@|�qO�1 Q(�|�t��Q> ��b�|2"�.6�u�V�'S6�h[������ �~���1�"��eJ��?1a������'C�ٓ��S.��z�A�1�	�7̎y[8�@��΀w�t���'��](s�ϰ���V�Q/htb�3�'������1)U�B/3�\*����~��Ёg�U*)�:�Y���!��C�	�2�i�F�U3q$��
gO�0��z$+�.�^�>C��0vt	a�#p�q
��؆ndL(���2F�B)�*���'ʄA��!Ц"̦Xx��	E������ԷiR���{r�K�t)�Ha2��#^gR���S�? �����>�Ay�Y),�
E:4:O��D��A�=��������p`d���N\74g�=��R�L��I�L�`�tAwϳ�?���}ܓxZ�O�Ic�G6���@���M��9OD0bߴV�@Ղ��N�	8<�¤?�r�8�3u.@�,b��8���x!�{�Aax���R��3ht�G,; 0�q�8n��:�6�=�@pö3X�^���Ċ�9E�d  I�"�v��d��;�ق���\܈�����f�FS���a�qO������%<���B�?xt5�0�|��L1t,��0)�.�xa�"�>��d�i��'��A���*lS"�0���:��葝'�8tp*\�(��t�Pe�1[��Xt�S''!�$���X'L�����2p�6˓H�2I�W/�<�3C��c�Γ;u���D��s4N1)4N��22HF|Μ�Y�P��%`*�A*�
��c`�OJ����ȟ �DD�W�'pf,͒K�N��;��"f<��f�Y1$9��L�^�'�X�"f� ;��λ-l�i�)W��X�2�*�!U�,�@Ğ��?)㌝8,����|j�!'�4���E�ٰ��k�D�Iӂ�#	TؔȦ���'�JeQ�ȗ;(�]�!j^�VtH�N>�&GP 4~��pkƩ4��A&���	�Ο���:�Y�H���EE�� ������3������yrꆝ
\�@�,J�`*@{�ɜL'n٫�M�!DK�e���G1O"e
���gZL��v枭j��)�֛+O$� `j�*?j� �'�`���LR.B&v���+ !�+��dҶ�\�K�F�z�|x`��"�&�O�xa����lJ�ɝ�*���~Z�O6'�)�5�Z�Tyn�H���E��e!uJ�B�'�$K��F�d}�yλr@����0/�p@�A`ɭQdf�j5��N��@	:D�6�Ĝ��Ɛ�7��&P�<5�)�,�hHp��O�� �0��$�*!h�@��Ae�BK����'%(��f�7^���I# J,BV�ڎ(� 9q�
y>4��z��Qٕ	�8d���Q%�W�&�Y�4O��A�ЅͰt �E��>�zls5l�9d� \:�[' �D�ꗢ7�S7 �Ը���&w��B�j��+��`��ɦ�ڄ��\[�nZ= �T��+ɔ0y��c�"��">��%xt�c��D3K6(���Z_�'��P���
98�>�q� ��\��c?���`��d^ �y�������Yh���I�"�g뎡�4�Y[��]�W�ʔ( �M5
��}�@�
*�&t9�E�"�\T��,��<A"h*�'�L��"E9O�޼CÉ�w}ؘȗ�T�.-\��=It�G�V�|x8��:nv��OD@���Nh�Ů�!�2����i�����:�X52fes���6HOy\P	�'�E#�6d`Ack��qn�}��8ga��Onrq��?Qg�aك�I�3�F9��.��'��9��*_�
�wb�10�@A�t��=xF-QE�v̀�4�j]҇o�2D^Qb��pSQ�� 1ʌ*w&��.M�0z��#P� D�8��[�y�"aZ���a[���=D��b��B�8&Q��

n<��Q2�<D��[� D[���F
8m:�� �@>D�����O�*� i�"�T�\؃5N;D�@�ԉ�F�^|����D���*Q�6D���2+ɸBS���@�ے5�&졤�3D��p�*nZ��a�<���B/D�̡ I�b��]zU�W#4��m+D� �BD>:�t�+T'h�YX��*D��rA�T�j̑R�Ewj h $(D�웶h�2U~v��RI�>:�f(�-)D�h���?�2;�b�	8�a&D�<��$9R�v�ӀA�%��ɠ%/D�pb4�A�8� �����;'Rd��"D����W"ֱ��I�U� h��!D�0���m�$�l��`�8�A4D�8Џ]� �j,�A��;�H�	?D�Ha���3&߶�sR�A'^��逵�!D� ��I
�:�m�@�
�}ĬQ�f� D����@��%?<���,�9*8���o?D�d3�
M�e�4����E"�&�K��<D�(y4%��wI
�@��/� )r��<D�"�e��=p\!�c,�W����U9D���wV�0�FHR�Kޔc`�%�,D�h0d��=+aD�hbA�S�>4!&*D�x"SH��`���SIw�J��:D��bbN}2��ߕ!��E���7D�DbulH8���ڡJ�
i�쁑�G2D���MA�"�*���a�'Mw���u`0D��yǠ�+up>M�F5� �č/D�h�Q�x�z��s+M/dٺ��rD/D��� i��rF�]�DL�O� ��G)D�� ʽ�T��3bH`��	/!����C"Oظ;r�D4Р`����]Jq"O��r(��bܴ���n�.'�� [d"O�M���>!QV�8=\b�9�*B#�y�g�(l���+��H�-Sh-yS�9�yB/\gÒ0C���sҦ��Oד�yRaM	z�LB%�R:c�A����y2@���Ĳ���)�6t!�eN9�y�@�?�t���E���إ�\�y"��'n^@TB5�M�� �1vȜ8�yRΘ,+�j�̈́'�f�:5!���y���*z��VD?p9���B��Od�C�I�m$�YS#�ƸXQȁ0D�C䉃}�D����H��(��̆<@�B�	�G��Щ%����ȉ��� n�B�0.�ơ�C��7�24K�A���VB�	�dP��5"*j;fL'�6a�ZB�	��x7�I�0�za�ƌeh.B䉙l�](T�D�F�(�Yd���*B�ɚ&���7��0� e�9c�B�ɛE۪���+>�&���!#�B�I� ��\H0���Vk ����?h:B�	/?.�L���N�e�+Q�
B��K�n��$�64�j�ة��B�;\:�� �5��dڇ���B�	2���1���f��p����ǶB�	*W����EJ�d�0p�Ъ0�@C��(8)J�S~��8�.NH6C��:R#�I�Sb�!K�x����̫n�"C�I����x1oE,n�:��ˈ�$�C�	?�bI �ׇlq�!13b�)>�
C�	�q��PS'ŋ,h��"�	���B�I�) 85
C�?�.4`%� �B䉨/��H��S�d���B�X\B�I~T�e�tū/@���[,k�DB�Ʉp}(�Q@(\�G��1%��B�	�c�\��#�N(�}�Sɉ=s��B�	=iumX#E
r�`�I'W��B�I�D�*� ���rw�ᩱ5�B�I���M:�ãn�b񠷄?ݞB�I��ص�dB�.�LsE�x&pB�	�noމ����#N���/]�B�� ����*a0��$��=c$�B䉬-����ԩ�:9����x�B�I X0�p�ė�M�mU�X2|�B�	�3y.8�1��j\��Tb�j\B�	H�0T�j�;k~hpů�_g$B�	u��L��CS�F�^8����	��C�	���m)��R1�J�8Ԍ�2C�ɈY�H�U��u�Lq�@'> C䉧S�h�)�$��j��E&x�*B�4	Q�d�A`�'!�h@��fX'�C�ɿ	�.�b�6����j��D8�C�I�2[H�T+6�L���ʀ*�C�	��Y2���%�.ŪG(I�Y��C�3+����"�.^GT�8s�ȶזC䉒/�^�;' C?�@`&H']��C�A��4�W
�<����s��d�C�I$LO~L��� (̱���*3��C�	] P)'�ݟK7PT�IN�I��B䉜}����k"|�ԩ����M�B�I^��ui�ÁS©���8�6B䉫�B8�4cV�(�9&� �P�BC�9Q"��a]�ݜY���y��B�)� �҅��9���D�.)kD�	""O�8@Ο4�B��g�κdd~���"O�]�ğ-p��y:�́�x�ۅ"O�g.�����`�l2{nH=[s"O��ď^�E9&A��"�?N\Hb"O$�A�\�d]��� J*0�R"O:�S��:m$L�!�����&"O��k�f���e\�|��!"�"O�����X�*��e!��G7;�taq�"O̔(�	��6B� ���&n���QU"O���($=
��bbI!�
���"O��j�%�}�Ꝙc�V�CW����"O��wJ�QB�#�oU��쩚�"O*�b�'×T?4(��LH6�(���"O�"w�7p�����b"O �ņO?n�d$9q_��,[a"O<أs�k���F��4����"O�0��*"'q��
`�]��H"O�l�aFS�9�,�mJ����"O���aٳk�T���F��,�Z%��"OT���C�7o4�"��@�Z���"OBU�3:�Q+gE־!��:Q"O��q��ɊXq�<	�C� �8��"O�tK#/H(4�i�� �F�(��"OJh�� @�m?T���/��0���""O��Y0&E�~s���-��wu�8ȑ"Oʥy%Or��C,�	5��)�"Ol��C�m��C�+�:n�<��V"OvȲq�Ç��V��?��xG"O���L�^⺑����]Rr5rg"O`��3a����W9F
�p�"O�@�7�O�<�*��� %[��S"O�hX��H��1���� fS�`��"O ��f�!,�l3��]��"d"O��
��¶!��{E+R�#q�(I�"O�`�wG�5F,�#�	�%k��r�"Ol!�e؊PR�befW`U��7"O���`���;�~�K��	�!q��!"O��ˁ�W�p��3[.YY"���"O�,�e*9n��d�H71���hR"OhpSgiT1fڂ;f,�=K��(��"O���Ț;e�u��\6 ��u"O4��0�S�*���k7&Y�X�q�1"O0����a2��ω%%s.1�S"Ob=��J1���#�� �uV&�k�"O��� UH"�"�%��q:�"OʍK��V�H�B0�3��'1Rs"O�TJa�̆ xl��VBS!&5�!"Oȱb.�=2�V4qu� ��!�"O�l�ε]�T��j�I��C"O48I�@�<��`@��#Z��@2"Op9h��ŸH�&ءȚJ�` "O,y;7�Qy�xL�w��lϮE��"O�<ÔHY�{4:]�l&�X� �"O8�	_	HZn����<g����"O"�q���2�t�#֑g�T ��"Oh6f�ޡXş�H�@�"Od��ÀC�:����%u|rv"O�X9�/J�� ��!
P#�"OR!�A�ʟW�ȭ��߈'��mAw"Ot4i"*�>ݴ�)@�����@�"O�-pRbD���3 E�c��l��"OT�xԢ̦�B �b��(2!�(H"O�D֋H�$C,u	J@�	�"O� <,��)>:<���GO�0ɩ�"O��0�@�Mn����@�t	��"O���%��z��I���� x�򡑕"O�t��� �<q��i�d���*&"O����Ƃ�^�����(�~���"O`�Z��S-�9Aק�vP�i�"O�8��RAAC�� tP!��"OZ,x�f���:�!��ln �"O�m�.O	/�rs ��Rȩ��"O� /ܺq�AF'U�h�{�c�Z�!򤅄=�L�0�a��1���(Z�!�$P�L@��Ǣ~V�e�7�I�?{!�$ܷo�΍���@-sV����D޼v�!�A�C\q� !�;T�5��ʆ%v�!�L�?�p�;�NѰ?��[��׋a�!�I#e�:�@��O�i��	�deN�'�!�ď�!x����GL��Jt��o;!��$u�ؽ��f˳*�<��,�
=!�$�;�$����9!���A��O�!�$S�\��X��`�9H�b�9@�D�!���>@�NT��T�w��4	J��!� 6]2|h
�ƻ|y�1�%�+�!��?N�lqs���o�����ʏh�!�E]`
	���8J��PP�4�!��8Ia�Tbc��;���x6C�!�F����у�K\��)'�֮wL��Wx����:x��9�')��n<�&j=D�Իd0�tđ%BX�Y*(8��=D��r5d�.�5��fI"r*��e� D����b�&d���ٱnp���Ђ;D���2j`���sm�c��yE�8D�xÆi�;4*�S��X4iL���d(*D�0���IA�{�NV�S:����&D���d釅:�QO�:r��a��.(D�,�ܟ"�ڹ۵@N4YL��sa*D�<��k�/���emY�#l�Erc�3D�|����j��)���1z�R����0D��)��E�C��-ڕ/�B��Ap2
0D��[A�
>�m2��� ��ѣ+)D��r"H�t��p�V�-��<{'#-D��ygeG
[���\:\��4�,D�|y�g��#ʘlK���o1^tj��+D��a1H@A�&p�G/�Kj�bc�'D���5C�y�����D�t�N1�+2D� ��b��|\�rIW�:}Q9�/D����g��|�JUZ��(�u�9D�0�bM،Y�-��ҵg��l:��;D��r��>(!ޔ��`Ϡn�xH1�9D���띤$r��uLM	5(82t�9D����u�Fa
t�M�GC"�4�3D�tR���!�y���$<��fk1D�4+�MѬMLh�c��K)@S2���o/D�`�6���H�9g�
v��;`.D�|˱G^"k����g���:�Δ�e�*D��"G)ïz�=� ��JĶL�%�,D�����P�BfꑏOxTv?D��ZeaB�<Wb-�W��t�2i<D��@Rj�����x���U�;D���t�^�L���¬O�A�e�2�.D�4��JlV�ӂ�άI����2D�@A�,E�`���;_�|ѐ�/D��R�YGvZ\�e/2!���J#�,D���3�&P��2�N��\2�*D��؆��(���9m(G\p��$D�� ��:WO0wޖ���Bۯ.���"On�3��!>�M0���7��XȐ"O֙B#B���ب��=Q�RuQ�"O���-�eM��sT,zt�*!"O�����@	K%�Č��)9t"Onk�`k|$��QCɤ6�R�1&"O����6�N�c�b�!98��i�<q�j]B.��B�?�УN�<9s�K4��E*0��X�Xx�O�I�<IV�	 �\	��Ď���á��H�<��I�q(�It���T�����!�F�<q0Đ�pJ���NB�Ť��F��<�P�3i+�r��-���n�S�<a'��7/Æ��K Ns�Õ)�z�<)�B�>:[ʄ�DV�*����"P�<�'�R-wGn�;Weӟ&��`��H�<y&	��fo�岠��e���v`B�<9"�V2)�������Z���E�}�<A�%M)-Y�j��V����'Qn�<�F+�nQkRM�]��7+���y&(H�:��D�[��5�wΕ��y�P5j����M
 @h� d(��y�ɕA�R�2�lA#"�d�����y2�����jᆟ=�&�x���yr
"�ƈu�+Jﰴۦ,�$�yRȕ��|Eȇ`�4p��4�yr�+>�d���N�/T,�R@�@��y�`
=􄴨�A�*-�%!0fW��yr�B$�2�Ӗ*��XˈL;���<�Py��	 }g��㰂ԃgL�8��y�$X�>"fX"����V�R�˚��yb?wX�۲OQ^�P��$B�y�l� ����&����술�Ԑ�y�厍9b �A�@m�@�Iʾ�y�c�,������ia�Ų�f��y��!� ���ҲgvT�Ж����yb,Y:%�� �Cm�Yp��x�CP �y-T�_��d��*ȹH#2�U��ye
e&ţ�&˞S(L�9�LF��y���6E��b�Jtʬb/˷�y��g��z��� �J�Q �y¯o�4�s������1J���y2ֈ�r0�"��R�Rahɳ�y�B�2t(0SU��t����i���y��k��Y{�,P�zAv4�@aѶ�y���V�j�i�gU`(�Z@´�y�A��%����JV�c���"�-�yrG/rKF�RO�j��e0WS�y�/�*��d��Uî���&��yR�Z��X�a�8ŖrV
�(�y�N�8Ä)[�\�01���5�&�yI&!2���I
�2U�@�Pxr�i�=A��[�T\ ����I^!�	�'��ɺ���n��3$�Z)��'�l�t:��R�T�@4 , "O�@&�#�f=a���5&�A"OT����"92p��NLP�"O��;qē�j��2�jM�'�L����'=!����$n�9C
0t�Ԍ��T�&�!�$@+-E���2	Z�tIGV,`!�$�&Ql��J�� ��Aq��ɣ{P!�آE�j�zq	K�T1bf�J�	6!�ċ*��S��Xɕ+� }4!�D��Jt���D0w��j倍[+!�� @�J��]	yu��I%	�0f�����"O�I����B�Dm�r!Ҩ{�0D��"O�����(w+�(u��#BVR"Oĕ1�AЫjt�����ԅ��C�伟lD���ʴ_�p��#���N�>�Qt���y�;�t��j�@��	r����D,�O�܊$
�/w��1:���of	�"OXx[a�� v��E	�WX��q"Of�IeM�d����T�s�|d�Q"O"�wk��� �C^:{�(��"O��kp���րP���@�N��"O����׸����Ę.��(�"OPe�wb�(baQs�B�D�.��p"O�8�
YA�R�i��Gdhh��"OJ����^�|X�mc�HʭD���u"O��i���u��9��FV��>��&"O��eb�"1#��h��M�*�"O�I�aݘ]���z�iK� ^�hg"O"�T
|p���Jr؄�ӝ� ��I#<lD݉Q/���:��7�C�+Bn����P'T�$a���ύ4:C��>�.=�F(زJk8@2���C�I�m����g������(2B�ɿn �ƨ
+s���!D�Dw�C��;�����9&;v4	��&�B�I> i���Th�<#���Re�O�h�^B䉧L��L�N_�0�jQ�=�*B�	.XWf̋.ZtP���\�s��D;���0�K=W�d�����$I��YG?D�$)3퐮d�(�����v�1�0D��+%FIr�[̟�?&t���,D�X�4@�3�;���[��[%�+D���6 Fi˂#M�>��A`>D�D��ᄋr�{U�3Nz�k�?D�,@-Ҟ5���J��%H��}Z�8D��`Bg�e�8�0�CI0l�~�eG7D�d@�D"K��BuGŉdtL�!�5D���`��E�z���iã^6�[Ѫ=D�ؘf�ɼI[,ٸ�c�$-���P�<D�$�Ǭk�X��J3&5�= �	:D��������%�F��'T v�Bl,��0|Red�I8�5b�D��v�mJ3�Z�<�G�[&
��W.�s�x��#L�<�T�Β��X�ao^10�^�"�hQ�<�b�9<q�l ��F.d����7+�M�<y`�E�1��i릌��1o����lG�<ARaP�D"�E��~Pd�#�`G�<	�Ꮷ.~�҂�ח99�]`�HOD�<1�kډp͔�j��_~����	}�<!ϧ*N�jP�Q�0b���'y�<)r���E��O�3��10�c�^H<A�@؋arJ�� ���<I�R66m!�䖁 � t %��'���J+���qO��=%?RRAݨp�څ( �D�٧�.D�h ���RY�m�4�'!����CD9D��h��̧{��Ւ!�?/v�h:�d6D�āe��B�)Ν�~0�p!!D�`�*[ˎ���h8��&2D��c�C��ٰ�V�5�8��G4D���F-`�\m� �B��25
%D���.�4G�� q� �D���20D����2$�!!�
6��q��0>YJ>�Q�\�>�C�C���3��t�<��k�^3� �F_�6�贃��s�<� HH��_�ZN h��ݴh{<<{�"O�ôX�7.��ѭ�5p��5"O��X!@B*K���c�yT\���"O�ٲo	�v���Q��¸^":�B�"O��"�@���Q��רim���"O�����w��s��̪PvI�$"O&L0�
�X��	�%A�_�N8�"OV̰�	^�@Q2dh6��$� d�W"O��bK�Kh��n� �� "O����~AJ�Gd� en �C"O*!��*�"x �QnM�,��A"O�A�ѯ�-!��ە��k��c����D{��I�i_�8�G�3g~x(`>	�!��h؊�*t�G�(��UgDλ&��F�t:mnx���!ap����N��y"#�#r�D ��X�EC5үr2 b��S�g~�+�%i�M�7 �Ws:�Q�@�y�K�*��;`⎡G��� d'Չ�y�Q2`�١�
��A<9u&N��yb��J9��ʵC�42�14b�3�y�X-v��=a��u �yTӽ�yR斫g	��c�N�Y��4��%ʇ�yb�_��	��&��!F�8�-��y��U"ObT�ȶ��rPP��߃�y"�O+C�f��#eҲ00	�B��;�y"O͡[vd
��L0[��!���ǲ�y⏙$6tF� 5-׎|��}9�KL.�y�BH=�B0C��_�z:��������y�d
�b�@Ȑ�u=D��&����y򏝱f�t���Ɨ�k���)����y�	�+����`ǋK�
��E��y�J�����ګFw�!��eQ��yr�Cu�lj��߿w�][����y���k�dkt�������y���+r4� 1� X�f|�d:�덟�yR-�1���[1�c�"�S'�@��y�.\�&�|� 5�̃U���hV��"�y�&�3Y�X�Q�� ]�	�I�(�y���\�C���3cT�ٕ�Ґ�yBkXB`]q��D0K&��4l׬�y����o�����&�;����-���L�AdP/X�F9�3�*'�x9�ȓ0ݜ������+bH��W�Q�4��G�~l"��#� y���?Kj���ȓF>�,�e�Ģ
�r&K>9�0Ѕȓ�(�5�􈳨5	�ȓT8@s��A63Z}���ʲ܅�l�U��*�>��� �3h���ȓ 2��xR���Z¤�&\^z���ȓ~cj�O�
a�*Ep�.������bl�����! v~HCF�6 �I��/<��zҁ�(�>U��`ثYO&I�ȓ ��D2cķ0@& � 
,#±�ȓ#i�PC�QN�QB��a��}��'� ]�RE�4V�(���.�\��'�\h�!��B���%�.{���		�'lVi���P�(#�Ђǅ�*]�N��	�'Ǻ�Q�B�
E>��@'&�
$�^͈	�'�����iΌ0����� ��;���	�'�@AI0�ƩC�����E��ք�	�'���[���>�M+-��Z,Ɂ"O�mb�݇>Jy�1-ɐ��%�c"O�`���6�L�1��S�"O��AL��ʕ34�+l���"O� T(2Qj� ,�E�wʃ%7�Ω�0"O�)�wl	�a�89����ml2�+3"O�-Y�ST�(���B� e���"O@��*5#��BX=+_(x�F"O^%��^8�I�6���"�����"Oν"PBc�nx{�OI��]h�"O�i�'�؃x��0�� ����$�u"O���_�1᦮׽lQJ��6"OЉ#��L3�����,�r[��ʄ"O��Bh��Qb���յUKzhpT"O���f4�� !���3�^���"Ob�B��
?	8�Q��8f�8��F"O\�h�*�F�Y Ɛ�Zmp��"O�]����7����@o�(Kj4"O�-�F��&4+W-Ä~5&�qp"O0���^�!30��e�N�V)6�`g"OD�ɧ�E2fl��ce��>'�,�u"O�E8�`ơhy����|`�i"O�-p�A sU�uf�.�"O~�;�e�S�d!���s� �"O�,:��wh5a�ď?����"O����h�3T]�����=�t\��"O$��� �2��-��~��,J�"O\�Z�O݈3�P4��� fv9�s"O�����E�ڍ{aō�fU��S�"O"Dd	�4
����(�@�I�"O��{���f.�m;#8	�$ "O���Z�&�h������6"O
$�Df�z��)���/+�U��"O~��Fɜ3G�)�'�����P"OT!�0 �%8�*���o9l��Bt"OXL�F*R���9y"�C%1���j�"O��'��3/�Ihծ5��X�#"O�
r�_z2�!yd�݃q�Je�"OvI�T�]?��I��ոw�0���"Ot*��&l���6'�Ɋ��4"O�LQBD�b���j�K̐QI^!!�"O�=�+l��6�L�=H�5�"OLH[���!䘲r� ,j�T�S"Ov�z�/sjh���(�5h�"O�$��猘psl�gU�@��`�"O���Td�8-j@�鍛z�ĕ��"Op�1�ڠ}�.E��P�=�b��"OT���%B�����"ũɄ7h0D�����ȯ&8�Hbc�.<XL�Q�+4D�XҔ�QI�r$)!DA+M>��3D��8��+{��$��hʔv�NP �?D� �t$J9EP~HK2oF�X��yTj<D�\!���;kX���
CJU��$:D����C�=䎑�ũJ�T��-8D�����U���;��tI���l4D�܀�����2��B>:V�5R�=D���2͇vpx�H!�aBz�E�=D�����!2Jyۦ�ZQy���b;D��tG�>6&�cf�T�?^����9D�XX�o�$�*Q�.5�B8�� 8D��$.��'���D�hR� $ 5D���!&$�Ya���`�-D�ܣ��"���@%D��-���ʧ .D����c��j�B7f��|ȁM)D�h��[&fDYC�, |/�8�&�*D�t1�!S$�2u[J��4p~x��G)D�4�3��D��\���Q�z�X�7�:D�x ��p�Q;��8[	Dp"�e3D�� P��Aς%;МCq!�&aK�"Oāص�D�E# �f.8&�!�"O)U/de���{�"O�xRA�q��a�A�5�h��P"O�E���
S��٠�O�B�fdۦ"O�Ljp�� ���N�D-H�"O~ق��2��0h�n�'j�4d�"O���#�G�G��<�m��G�1x$"O��2�`�
N;�<�$lЯ~��Q�"O�|��
�G�ҀH�+B�lVTrS"O�١B  �=�t�E�US`�Zv"O�M�˒j<�|�t�2x�B$Jb"OR�h�FC�E�6I03g�1��Q�"O>(�B%��8 �&� ����"Odd�r
L�s��J�����<�E"O콫#�H6W{��b��3R��'"O�̡p	�1	C�1$%�8Vk ճ7"O�AJ�D͡��)��WX�8iC"O��b�3Lݲ��,��Nja:�"O�[s����	X&j��=��-"O���N��!GL,i#�x8�lY�"O>y�vd�TBҕ���#���"O�[�DD/i�q�&N�q�,�"OȈ+�e�/*��iSMM�i�h�"O��{ŏ4&!�HFk 9����"O^�K�Q+p�!���[�޸q��"OR�04��c��XdH��/�
��#"O<��@�c*,�F� &��0"O��R��{�	����Q턭�R"O��Y��"����C�*�V	�"O2i���.r���$l
�az*�q"O��	wV��;���"[te��"OnlЀ��|V�ѓ,@�X���"O��x���1p��JEĲz����2"O�E;�
H�1C��hc���ޤ�:V"O�` �ʛ�"��|a��F^d"�`�"O�0SCK�a�����N�64�"OJd�J
7l���D�F�k�=�5"O|l���	3�����9DC�H[V"O����\;��K7,�I�QQe"O>���ꞨW�m*%��LR�ȁR"O�!�H�P
��7)�9c�4�#a"O�A�1�ֹ�$���++��;V"O��F�J�`t\����*o�rd�U"O��ҴkO�r�XP��c�g(l�C3"O
�J��6���;�c

f���b"O�	`7��AK
9�͜YWD1�"O���wLH	��H���]r�"O�D㦁��e�>%�0�V�W�2��"Ot��7��jAb�`ʹU�2�`V"O`�xS/m��街�Z�`��!`"O�c���?�v�/� )$�La�"O`�J�r� P��!T�h���"O�ݙ�d��D1��ʅ^O�7"O~�X� Ϩq����LǄk�ֱi�"O���k�6<l	����(��!#&"O��P0I��%�F���-F`�9'"Oj�)G�� b��ģ�!�!�Tѩ�"O0�A���-_�.!R�&O�~�޼;"O�:qg�%�J�!��	�k�̚�"O��3�!Z4-�tL:E�*�(e�d"Om�w�� yȦ@(�"�!�"O�2䕮&D����9�B�z�"OQ[��$�X ��u���j%"O� �Z�[��lL���
�.��"O0I��D�4��#�@��l+F"O�ae��,����`t;�"O@�`0!׹bކYB+��gxh�1""Ol$���l�
X�W�opr�q�"OT��R�>,��ڃhE !����"Op�$��o�Hh����@��<b�"O"�rK�z>.H�¥P)?hXx8�"Oq�wO4Y���ؠ��,3�TY"O�s�m�"K��x���W�%�85�4"O"U�c��YP��ze�Z)$ŤH�7"O��F�0������¨|����"O�hR럻������p�z�#1"OdP b��&�Z؈���T���"OF��SM�C�a��B�9~2H`1"O���� P�\ӧBT ���R"OD�(���2NiX�"�?'�*��"O�yq6��Q`�hzw��Z�Z�)5"O��*�.?�V�Qa�5	�\`3!"O0�UΕ���*�eWj��""O��WO�������/�*\މI�"Oj�rl��2;@ @g
�@Cj#w"OL�� �$��`�V���Y�>4�1"O��	!ҤZ��q��N�l�x%@d"O(4��Ũ3jAi�'��i!"O�1����#c���QP�E3<��E"O"�ЂG�)à�3K�C3�Q�`"O^�8�J�o7�@���GP,P��"O��8� Z����6	İ��"O�@�A� \���$�[�� a�"OJ,P�Ν\"�� ��h�s"O6��)JdȵY�-� /�|;"O���PAP�J��u+��+�샴"O�Y�Z�B�d�&�5 ���Qd"O�M�b
j|�P���Q�ZHd"O�����g�R(��^���'"O��EF�� ����w�x�3"O�)�b�#'H2�1�a�>G��<�4"O�e(�g�#y�0d9���]n|Ec"O2D3%�(>���K��@2Sr��"Oe�	�#v,��hǤE{|S"O����LR7>Q~��L,kTQ�"O"��,60���؅��;V�x�"O�� ֏�/�:!�c�"����^o�<���9z��XXEÖ��(|�ȓi�lQ�
&$;2���e۽v6,q�ȓ��-�4fɺv�&�J�Ӵ1����ȓI��z��Ê.:��r��ƴ"��ȓ5�Ă2LY `L��6�ԇȓ|h��J�/#AӜ��Vl��1d8��9�8����ŐVV��v����j��[
l�H�"�vӐ̻'BCs�Q�ȓ��3�\vT8m˷�����u�ȓ!
\�P[�aP��W$R�J=��!�8<#�'G��>�zUn�\�����C��qQg����0P���ȓQ:n�[��Q�Jx�Ј���Q���ȓ^݂D�Q�;��X�m�.��u��O>�`�4�"9d8؁�n]�4����ȓ2U��qcO	Q�(sV���6�I�ȓM��!�j�YH������M�4��\�����)swnq(�_ ���ȓm�dA90a�Z�P��쇹x�6q�ȓ��Ղ�F �g��!����_�dم�S�? *(@����$��݀F��$���9"O>�9�H��]k��
��E<�Y�"O(8�	�.2�|X ��~���
"O
h��ׂj9�a�2� �N��"Or`3`'Aw�ݨ0*�*&g�I�"O�Qr���4�>�{`�7๋"O��Y�aS�%�>�C�M%b֘�7"O
	�%�~eN<�`!�!rM��"Op���M��p���E��/Qb�]r"O$�E.��%)FO�9��iJ"O�z#�]!M~]�7��C��x�@"O�c��ƌ2�4�Wf��D�q��"Ox��	إ
"8[S�ݏ�la"OB��RK�-7X��ӊ��y�8�z7"O0�'Ȉ-t�A�)��H-`=�!"O�A	�fO���t��n�	!N�R�"O�E�5�Եk���@��U�T�:u"O��A�F;g���!`Bp_z��"OPq�$�A�+�4�X'nX*E�4�t"Or�:0;�y��62�{C"O���'�<=R��qå�/���� "O6����@Q���-p�T�"O�x���f&J@S��-s���%"O){�#�3&&��T	I�%
�'��kDj܉a�Uk�ělײ��
�'\���%�WX4.ݒS��ed�r
�'�&���z�YHd$B8c�L���'춐xu�M(4�@�X�g]27�ؓ�'��3r,��؋1۲�ک�y"�$>�`TA�� H��"ф�yr �\��9"!f�<f��5����y�I�]�PQK��V4a��������yǁ�V� f�W���4ͺ�Py�j�*��h�+�\�BB�LQd�<� �H�KMz4
�a$}�0��a�<A��?�ҽd�W5��(����b�<��e�������2B����  �\�<)4#_�mD�%���ï90.-�cTt�<)�9�b��$(��m7z�+�E�<�*�C/�]�W�@t�� '��D�<QtMٌ2
I�C�׻e ��kEAS|�<��a߸e��A���Aj��0���y�<����"�1@e7��2A�@w�<��
Ɉ#�6�:���"p�Dhr�<�E`���m��b�u���0�n�<��@E�亜�2W�;OTt!��j�<�b/߼d��sg��;O���p�f�<٠�ռ_~AKE��6q���R7�K�<S��+�����2J��X+���G�<�QE����2�e]B��a�w%G�<�a͏7} 
6eC�'�~#�	�Z�<!�J��3Nlp���6<$(@v��U�<!6��,"���S�(dN|0�$Y�<Q��K�J�t {@�&[t��XQh!��	S_��Ӵ�S*v6pd���K5�!�$�*t�r�K �2~�X�*�<�!���S�u[�@�V��a�Z�8�!�D"33t,a��ޔF�z@3�g�L�!�ğ�F������?]�q0!�䒺:��}r�A�-�� �dC�A*!�D�;�R����-V�^�#� !���2R�,�J<Xm��e�g!���{��=�q`X0MW �r$��!�䉐v��I���X��RuAm��\�!�� d���Ą�^7m���>	�tK"Oz��u+	/d1�Gl/B`���"OH��T���h,R��,]!fE�"OLq��I�L���GBZ"`�g"O&���f,$ycM�8@�"OV�Hr">z\|@��ǁ����"OT	W��>WZ�1���&aK6"O"�3��ʱ
R0Q�f�Ja�-��"O��� �:8�h��=T���"O.��K]GJ�L`cʄ9Q@�S�"O<p��N�N����#��$��{"Op%�rAX�v�Р��	�.�ې"O��@��%v����b܀P���z"O E��n՗L ;�>+[R�3"O:��g�K� Q\i"�� H�bѢ�"O^�Q�L�`�!�oO<!�vYw"O��E�T�
Pk�E���"O���\�Z�0H���;��ٕ"OV��s!=4ejY���V4"3�	��"O��1�[�K�x�s���7�A��"O,tIdD�Xd��P$J#a3�"O.q+�Cˮ�2}�5#��,�f"O�aq3IE #���j���	�QӤ"O�7�Ò>�!���h���g"O�L�@ׅ:��T��� .��5R�"O0�ôJƟ\���I�`�.U(�40W"OȬ)E��64���둈���m�F"O�4�3)�&'��ŀƍ"yxd���"O``PF�W#3$�͸ �O��F�X�"O� ��i˅���rC��G��C3"O���HL������~��w"O �����=J@� ��A3's:��"O�I��\�E�69!.�&X�D�Q"O�l)F,V�8�dtjB�U�)~jC"O�j���]_*�s��)\=؇"Od�hq��&@��,V�\5��e��"Ov�'��x}�%��lQ���"O�e1E՟23�s�/uI�*%"O<%z3K#3|���
_D24"O��:�cV4#�Lᓱ�ؽo�R���"OV	���	xf
@��BSu�⼃�"O��;n�(;�|A�z�-""O"�R3f�T���f�Z�*U�e�"O�H��ɹ|6���W�%���#�"O�L!���83(Z&�99��Ɂ"O��$�L��xb���z�F��"O9����=;$�9ёI�q�~P��"O�4��E��X��ʜ3-p�!�"O�Ё�&JC^X��5DP\"O������J�����;b�b}��"OI�"L��I{dX�$n�=N�L1#�"O��Ka�:� (`���t�h@�"Ova۶�TJb����N� Du"O�1Ѐ�(��1t7�I"OT��w��8'��!��sNQ�"O6m)t ��z���E[ 򰰁G"OL�V��>�9)�-�ʩh�"O��37�Q(�b��Wh$�1e"O�9�d��0h�Z����te�0s�"O�srB�(v {�G[wR�!��"O���a'ɥ�T1���*Ն	�"OP �Ug�u:�d�A`�c�p��"OΉ�AO =��l���h����"O����L�"y�T�efϟyvH��"O� <e�A�?r�'M�p�"OJ�p��O�$�$��0x	H"O�|�T+�{� T85��V@��"O����	 ��e�0F�"S򰱠W"OqrR��^� �zD��&s����c"O$txp�Լd�
`��vt,�A"Oz!)PcE�;C �2�`
��t"O���E��`�GNJ�""O ꒊ�I^R�D�Y�T.x�0�"O��9w��f�x�Ac�dƲ��"O�q �'W+�p�SMB�5���s3"O�,hS D&HK��W��|�|M	�"O ,8ơ��/%�3�"�.�h�*R"OB���+��vF�x#�C ��B��"O�,jPl��#�D)��_�����"O�,� KX."�d�C��K��92"O�a��0PZh�b+�2����!"Ob��2�Õ[��y	�*"CvP���"O���5��bo��Yco�C�y�q"O��[gV-��%+ �P��Z0"O.�vn�1*
��\�a}�L��"O����J�`�p�# \gH��"Oz���l�:l��5k%.֨K��1"O�,X'�bt(F������"O��U�ؚ#���č�4���أ"O�]�DJS����Ꝺ�Pd
v"Ol�聏�.0z@�'j!6t$��"On]�qiÎL+xh���APN�9�"On$��85�����K;h�9"O�;��YB�����@!hp*�"O�]"6#�8L*xS`ν��"Oh�PQ�_$$@SB ��-�$@:�"O4��5�L9���
�~%��"O��C�_m��W(Y9�����"OZ�:'�	3x�(�P�'X )2�G"O�;�CLtC\�J��B6�D"Of�@�EJ	.�Ie⋉T|��6"OBm��-�sTFM�w��4
PlX�"O���'��l�F�9eC0� �r"O¹〃��!88���X g�r�"O\Ya��]�,�����<T�"��"OF+�%Y�KUډ@0NN���p�r"O�x#Q��~���B�-�Lm1�"OxI�����)�R��a�<���*6"OViB��V|J�:B�t�d� "O��a����NC�@Qu�5�p�
�"O����0����� �'����"O���gG�%SN&��J�OV� ��"O�QZ㠂�����g��UMl`IG"OJ��D�B
]�����%�z�,���"O��C�F�_j���Ŏ�!��!��"O0��eӚ	|����u�� �6"O6h�&Nǌ�����Ɋ�Cl��"O���Jʨ0д��R�֌�=A�"O�� gjS|��ѧAW/Y���"O��T��.�>����R����"O�%�����(���i�v�H"OD��B�o�0�kc��jf�S�"O����ɥE���xe�Wvi�-��"O�I�凜yN�P��cȿFQ����"O0��Ө4N��`q0�^{<�p9�"O�}��,��}�\��G`�=U2��"O 	c	O�:�R���v�3�"O:������	��[�k(��m!�"O� �=��įDq܄���L2~�^-��"OR�$o�-S�RU��63�$p�F"Od(	�́h�\���t�,��R"O!�IUbN-��fX�Z���$"Op\ ��I%�rLؠ`봠`"O��kT��a͚�z�厭SH��"O�0�+1��)"��:R�D;�"OB� �˫�d�	^�VQ��1"O2��a`P�*��L��n?a�	`""OzɠS儒 I�)bB"8#��{�"O�p[t��J���B���p��S�"O�SP�oP(�O�1G	��ӧ"O�;�"� fּ�#b� `�B(��"OB�Q�@F8_/�ti�MɆ&�T	b�"O��v	
!pбb�-�-"�Pq�G"O�A��kC�a��9�sKX���&"O����˜ ^�a�&�N�眕2'"O�9[F	'~�l�fC=uJ���"O2)��"ʄ~�A{Ì��'�� �6"Oڑ镂�/�b 3��v[Z�[�"O$=b�-ҩj�P��@�ןs�jT"O�}R�gJ[æ@�%i�e��J�"Oԥ�qn��7z�c��֢]��Ȥ"Of!:r�F��2%+rg0]B�Y��"O<��@��5���2�c*(.P�2"Oإ��iQ"ho�R��M�RpK�"O�i����'۲0�OP-�l���"O��R���A<�9�w.��ԕ�"O����Ƈ$����UI!2{&�j�"Oj%��n�?�}���	0~eJ�+�"O�ر��ÀE���(��9C���"O�h���F-����c�W|xF"O�P�"��;U��A��[�8T�,�C"ORE��.�g!���#��!Q���"OlPy&�IRي���눈?��cC"OW��d��a�J��`L|�F"O(���MY�c0�Y�&�2[��L�"O>�����K6$9���:V��̰�"O���1�T 1_� �F��+��e:b"O Ő��\�x ��1F�i�Qr�"O�i��IP�Xy��	X�&���"O
���o���� rͨQ�BM �"O��a���+�ޅ��ض�B�9�"O�9��`̭A+^��T�i�� E"O `˦��j�%r�G^1�p���"O�$����il�E�L�P/�T�"OZ� g��i����'%� RD�U8�"O0��O_U���B�N�8"O���̱�iB(Q;%$i�"O����K�;J	��sU�ӆK�4���"O�Hs`�"� �߂Xt�"O��H#��#4j����14C�"O0�)�#�Q�V��Sf�nY�Ӱ"O>�y0a���˗)�u�"OPp p��%?A�!��T�h=ʇ"O���f�	��(iR��`|e"Oʅ)��A�qFؘJA���qe�1Q"O,5�r�@6qx^��Ծ>���1V"O�%��`�('�6�!UgJ�R��,P5"Oz$���)*�n`Y���w�"O�|�"K�_��Q��/}�,h�"OT�`��1Q-b�J�d�rH�0�"O(�"�=�h���BĲ}�<��Q"O��K7M\9��u;gT��*x`�"O� V��c���6j$R� ����ɣ"OVl��a\�#��L��/�T|l(P"O
E�w*�0���.�0Fj,L��"O��͐�d�Z�@Ӥ��7r !�"OjpA�fߨ.?��qb�ī~?�P�"O<����O8-�soܯT*�!*"O2�AaoAj���W�N' ��"O�<�eNȱ��M����37����u"O��:#�H�2��%؀Yy¼"Ox����Y�}�$���"_�ȴ�"O�x�"ú5�x�-�h�"O@���#K�1,(e��%B����"O>�bG	YS���ցj"4,d"O&ݒ�Ηq�b��bO	�V��"O�Ys��-B�́=�̋�"OpYb�G����{8=��"O��C�/f� 
�3*#�Dr�"O0�Q��ey��)��"J6`y
�"OBYkз����0 ��U��CPGl�<�O�IĀл�	�"7�Nq����]�<QaM� ��`*_8���
gNO�<	���9s�P�#�su�m" ��K�<��M���J��J�jSG�<����/��Qf��@y�y�<90���o��a7!��O�bI��Er�<��c�0Ap狌Ū�qmGD�<A��ܙDB�� ���j}�2͛u�<!TǓU�֡p� �<�ؐ����j�<aD��u`�e����v��k@g�<�f�4�v0R�W-N��p�,f�<1��NFpȅ'A�l���d,�`�<)���"�Y1S.+o߲*��R]�<9S�M%^��`��#
>2��MW�<IB$��	�A ��>Q�yK��W�<��H� ������ W����t�P�<Y��ѕb��Y��_6H�P��ਔq�<�'1R�x��`.�1G�^�*a��l�<i��!""��1w��)܊�)���e�<)p��I��pv�։u��9�1�\h�<�4aPLa17�=$�>�*���b�<y !�
nh	��R�G�M���Z�<q����0+�M
� I��0A�C䉴XR�d�U�̘]<�E9����z��C�I�X���/�w���	7铹<��C�	 V�\�cS��NՆ�j�j��O}�C�ɺ���V�Ι$�A����e:�C�	�K�z<���� m��dF9"�C�	�m�"5R��# ��@7B�71Y�C䉒'i�%�FF�9'�-ңL*C�I�af�r�/G;K���Ebm��B�:<�0YQ��r�� ۡ�*mR�B�p�I	��>Y��K�p��B䉟2X��2�;���bf�.
nB䉠S�|Q$&(BvѺAP�XhB��)t���P���<� �	�7�VB�jW����ՓU�@���ƻ1x�B�Ʌz�����ҋiw8y˅��TNC�I�
Wp�z�X���q�eAC�B�I�C\�\�"�S'i 걒R%�52NC�I5Z,�E�	|޵q�)
K�>C�
��h@#	�f�ĽK��#G�C�I?��X��\
H�R�C'B��=�HB�	�{�0TxBo�#?��U�F�6l�rB�	B�T̓B(A���)A�I�JB�)� rIF掁(�v��39�l�v"O(��q(��?��/�x�L���"O�S�@jBma�_����"OP`�%O�0 �4���݊5�Ddz�"O@1���n��HAԎ�,���'�x��¬�)*?�Q
�b܊p�©
�'����
'f��S��0�6I��'�$�0m[�n�4e�ꕛ �f���'#�e��`�R��?y�}q�'� SR Z!�4!�C!� >��#�'k��*�ӇP�j�X#Ǳ3�vl9
�'����'��5����w��;;���(
�'�]���� U�N�xTj�!9�T,��'�0����!�����&S�$xj\y�'V�E%W�{6�Q�[�G�*��'B�2�/�	N�����`�0p%r�'��Y���x�k󈋒cT���'."\!�'��
<��˳��<�$�i�'"px�1B����[�߂]���1�'�| @��0�k*��\�i�')��"�Ɗw���C��W�����'�0p��ih���@�Tn��x�'|�a��N�:�t�9rԚO$@0�'�4�0�H֨~�ș��C�}2b�C�'V��H5I��XK�qS�����;�'�!"�e��iyΗ�a��4p�.t�<G��#W��:q&�<|D�R6�F�<�7��$�|�q�)�z�R����<��&��D�\8c3�72VB}��^z�<�䍝ey��P`EG0E�RdMy�<q��.X��ٰ�M�P:a���q�<�$��sDBa���-rr<4���Ze�<9F�Éx�LM	���3d �i$j�c�<A�dX&`��Y�d�D��R�[b�<�"厇8��Iv��$��=�e+@g�<Y3kA�H�T@A��D�($��c�<Y7j	�~���mRx�������`�<!FO�KP��:c�V�]h�(�_�<ɣ$�/C}�I�� 2I���SC��<�$HWTĜ��␸o��Y���~�<AQ�@��)�c⊮;B�\�H{�<��ȏ4'�X �cc+*��@����N�<��-U��)�uO%!� ���*�F�<p��7*վ�`G[���iWT|�<I"fXUK 	Q�j��o�Fy��`�<�D�{��	?&~)ů�c�<��M*)���q N��+~W�<!���g�4
�Hٳs,���V�1!�d0i� 츢O�6�V5��fӥ !�$�$p����I�2�v��d敚w+!��\�\u�a
��eN,8��*O�!�P�jb��"2ȃ�[
�����64�!�	n`�b�*��%b2��9�'���#����]�Z�`��G��t���'�\	���5:�64��@}u:�j�'�d`*��J�Z��%���ؼ	-*I�'&�|�#eL;Ѕn,�@�yB��::�Ѝ�S�t��h�-���y��\?"�8�bjU&������y�U{͢aX��ԱzH��'�y��O��t���'yc|���f��yr��=b�$t�S.D�:k��;����yr.�R�PA�W��.����$	�yBg�C	�)�A�<&��q��y
� &A+	���4�G��ؠP"O�4�A�VT�2BAR!Z�3S"O�@)@��w̸��M�345��"O�dqbFW 29v�{�)ʵk���c"O��bȃ�=ƹ6H
�
HX4r�"Ofdp�`�� �!�C�2gA6m0�"O�ec�E��1�T(fH�y)@ܨ�"O��#�GD�D��E�"��0u"O�,C$��F�4Xطg�%��s�"O�]B��2f���ד2���"O
�P��i"&aR��\�NŜL�"O� :"c©z�^��a �($�¹��"O�1��H_(-�e��h��O�bh"O@���M�'N��`b�nH]x��"O|� ���8}�-qCP>fE�"O�9W�[% ��ѵ`��A�XL��"O������\` sO�O���t"OP����F�9��蓇@�8�P"O��
�>^�Qp��Q)���"O�і��e8:Z���k܊0�"O�4�`(B�pNL�Г��;��0��"O�Y�E����BG����"O�IA4슝 �j�����vڤ�B�"O�,Pc"X�x2^Գe��%R��أ�"O���a�C�Q�4�7	��=��g"OL��p��X/��)/e����"O��f	B>h2���Z�<�N���"O|�M�f|�X�o��#��s"O�x:�&cu�|{3�&}~��C"O�U��nޡQ�4Q7P�>D�"OXI!�����e� cէ�*d�d"O\@Z�ߩ`-P8�Bk!{��d�c"O�A�	�#W��(�	�-���"O���l�7z(Dzdg�
!"Ӗ"O���я$��)9��]�$�������Cx�����L+�.k��9�T�F+D����DN0L�,�
��U�,0�5D������8^	��`Úf�`z�(D�p���|=x��@����*Qn%D�I@ȪkX�rth_9c$I�3'D����0D�Da٤��]Y����!D�T�G��56��`[u�Z����ö$$D�p	��2s�ti��%�%�%F%D��Q�"�=Bع�'��nm��$D�����_�H����f��2J$D�8�q��'r� h8	�X�:U�rJ<D�LA#�=U���"*Uj�$k5k>D�hWoE=�`�x&CX^ԲT�Bg"D���eEɁb$h��&qn��;0e4T�`�f�D��ٙT�؏"Ƥ�ч"Oh�H���-Y0"�bJ� [YBaP�"Ohtj��ڔ��Q9T���"ONyK5��5F=ve�)*�d��S"OV z��ޘ%qRx�5���f���!"O����$g��hk"hS�(x�b�"O��CV�k;�x�g�+]� �"O����� �f.8��嚡C"D�"OT8�S?^v�y2���k��d"O��Z�gww���d��.��z�"O��D�0	��!��-T>݀�"O�㥎� B���֠Ї@����"O�B ��dȮ� $�M�T��AR2"O����N�eB�g�7󌰸"O�A���#dT�AT�*��-�"O� a
�݊F?��5��32�L���"O�Ic�n\������݋b�@���"O�<2�C�v�]3���;��A�"O�9#�X�������T�b�0�"O��!��)]������\`}C"OjYR� ��G�:���#+�Zm�s"O��"7��5[��J҂_)����P"O����G�(�ޅ���E�(`| 	#"O
�""��1Qc&ș6[gH�`�"O�I#�!�)Y�[!�J`"O��bD���9P�q��O�y+!�D��	� ��n�5����rOE�u�!���&�h���h�6e`��� �!��VYLS��%u4=Z����!�	�s"h��k�*2k ��\��,�'���h��K䬕H6�O�.���'�,����\U�M�t�6�~QK�'�ƩA�HS�n��9�7*���'�D��֨��Pev\At#&�`h��'��T���I�_	6��3��K��H�'��k��"U�N:�f��D��h�'�4�"���^�~�!�MW-�4�
�'�py'�EUL���$}]b��
�'�@e`�͕�1�Te�qW*����'�:�8a\46��d����$K�t�{�'�8�h�*�4p�v��AAߏxFq�'�ʱ��$C?�xzၜ�x�f��'ۆ|�w�) �D�C1Eٷc�6�+	�'9�M����O��q��0KF̝Y�'
��6n�6nt���UɎF��9I�'NL�!D];i{z� ��M62�@��'��!�BM(����5e=?�0=��'�ЀS��p�\m:�Θ�6!�M+�']2��4#�Z�$z��|��U��'@�s1�B�f��� eS�t���;�'��PG���i����J(n�|!�'���(�$�"��[EC�X�$[�'��*�oެ9ka��O;	��|��'�j����#�Z Q�Eͷzd�e��'�y��	�6��  ��7s�B�x	�'1ح�s�ؽg�t���nv�����y���bj�95K��Zn�a��̳�y���4X�t�Ѯ2��2e�7�y��3B��t�ք�c�R���y2�h�L]� ΀ �8�CWK��y��BJ��3%�*ͼ�/ڀ�yB��>}.��9�M�]`���y	hмk0�( RЈ�U���yR��Q�Q��z|�U�4�J,�yb�M"q4$��J7m&
�"�8�y"�� ���"AZ]#8�)c��-�yb,՘]�����ݱfQx��ý�y��Иd�̅�R��(-��i#�Ǔ�yb
*�:]x��_	(���8a&Z�y⤂�T�~�e�M�Pn	�w���y��WP�]𵆘"E�1!"�� �y��X�(��Y���7*��!hӕ�yB��(gǮ�� B��*3��j�BR��y��E�	� �иg���yB"��c���y7��`	x�@ٶ�y������P �͠X��AW)=�y��VTDQW�9<����fO]=�y2͌5~ԛw/��:+�\��gB1�y2[�3�y��S���#��y
� �@���Ĺ�"mZ����h��"O\IToH�Y�&	�C#�+)q
��"O� 0�/(G]p��1cG-q\�a��"O>���O;D:9{W!�!) <�"Oz�q�!āJ���AK�/�`#g"O�\	w��X� �!WL�9!C"O^]�����O�r�Q��
nkV�c "O�y
�6��[�P;cBu&"O��p%���6�L��A�QR�-�V"O��S4�;�2@��'n�M�1"O�1B.�*�H��d[8$A�(�t"O�r�@��E�TKFd�P|Ru"O������$p\]�2ܭo����"O��"p���F$	v�_<�&�jA"Onv,F�Y
=r#��~��r"O�Ez5+�.<���Ο�g�p$��"O.	:$Ά��|^�oϰ]�"O�rt���3�h���6D����"O����G�&��{uG��o�Nᪧ"Ou�K<N�AK;�x��"O
�s�A�|,lA��ly�<�t"OT����]�,��_�=\h��"O�Q�S�P� mx
޸'[�M��"O�	ja"�fH(��t�iV��[�"OJx� &Q�I�����#1Y�@"Or� C��&��]�҈�W6�0iP"O��`�j��IS� ���;Vf@�"O|�@��W9Z��e��'U�X$0��5"O�yYG��Bݚ鈇���z9 9Hw"O\�	[�P�N)x0�x��ܒ�"O����o]�WB��1g��;��\��"Or��#iȣR�����E �:�T"O6�'��#w��y��ʘ�Q�� ��"O�mjō�"���Qw'6n���W"O�i�2�[�$ P�c@�5:"@�4"Oa�i�6��s#�\ qp"O�q�t��^X��Ƀ�U�U���@"O�������4�\=���7�4�:�"Oj͹��Ŗ�"�Ū��if,`�"O�Q#��؛E�P0{�iP�/��8�"O�-
b��?(:����c|H��"O|�K@�ż)4^t:'�U��P�s�"O.=��@�2o�����?)r��'@(+��B�ޭj&?cP ��'����W���t��S�Y�
����'?ظU�r,*eRIZ<P2���'o�Ԉt�ۊdeDb�C��-�'��!V$I�#�T�����l�����'F���K�"+��x�%�a�J��'�6 Z�o��I�䙅f�g����'J�e
2fN4�����-�4`��,y�'�p�?j�}y��S;V�z�B�'�t��Ċy���`'��%�L���'���m^6kg�y�H��4j�'a�8�&ʚ�z��PSB�3LQz�'0Qנ�##��i{gGɧ�z��'���"Pmڀ}�V`�\~!��
�'�j��h�"����a`�=z�zͱ	�'��
��I&�|\�Q(Ĳ p��
	�'�D�Y!�k�h�5��V ��C�IC" �P�9@���XĨ�4Li�C�	2[�kD���
xԨ�}ilC�<=��Z���;'�	���S9nB�	�Q�X���܏p�Mh�ǁ*)0B�)� F$JV�Z.V��0��9y�$d�p"Of���Ē''(i��U����"O��b��]ە��xCV���"O(4C�W�S��}ɓ�+T-�"O�����-I�1:#L#*f�(c"O�yZ�bY�7�(pH���>�PH0"O
��2k�~���b,ˎu�(PR"O,@o2֬i���1X}�7"OAB�G�)�D�P&��HG"xj�"O(y�!��f���V���|�Ȑ"OR�D\#t�U#��Ǩs�,�s�"O�P"bρ��4��	�#T�T��$"O��pS����cƆ%V�$A�"Ot��Bٵ\�j�1�,N�u��|�S"O�E� ���Q�a��Rq����"O�<����49º�j�'	>zn �2'"Oܵ
�jI�.!p���@aA�p�(�ȓ �]"���pq�Y�d�F��ȓӎ��a�ԹY���"�����:D�@0��ޘylq �#	�yu�ٻ�6D�@1���a���
�O�Ju�.2D�x��J�P����%�H� ��QK=D�t��h�,�4��lF(�4��&;D��k���M3��J�����qd<D�Xɕ��8~�8��l�α�:D����8%�����'���O7D�̳�=C�&|�wCܺ~f��k��5D��c�͖?ɦ�V���LCn���+(�$�S�'4|��Cr$�D"vL0/]-%޲Y�ȓ_��ȡ+?Lx����E��фȓ%���фQ6��h8��`�V��ȓ��D)"N��,���J�b�d��y��v_�h8��Φ+�0�$�X5{Rل�	Z�,r��'�`̱�G"X�����}���4M�	e+��S��0�ȓT�L0+�	>��(Łۇd���V���1�HT�7�t��!�vT�ȓe}*�XXm��,�#�2� �&�p�<�V̏�7}DEzE+B+���̎k�<)�a�8fx��7��
$
l�
&#Uh�<9䡙'U\jհq螉�zs���d�<a�-��2Y��hA���!�Ya'_�<`��7��@aG�ӽ2����W�QO�<!!	��ԅ����L�A���N�<a�Ȕ�M���x�'��w��| ��I�<�p w����l�w�>�ۅ!Y_�<�e*ѱ�֙�GU�����kBc�<���S� �z1�� %�")��L^�<�q�I�
*�[�mڒN�$�sa�o�<�Fn��= p+�p�CSB�i�<��N�i�t���]W*L��X]�<!�Q0i�k5��[��"�o�<�7C^�l��8��%�Qq� ��E�<	�@� a`���L��hߎyC�jB�<	v-�,#
9�DZ�k)��}�<y������X�?0l�¦�Q�<i�+^ ���N��JDx�g�v�<)�bU�i�`%���ԖmP.��Qo�v�<�vjL0Yx�wEN%|h���p�<�A&0��0�P�_q���7��g�<�F�ʼe)�1�r�.1PL�So�<9�*��� �͟"8d*���A�j�<V�k����K 7�4J���f�<Y�#W�=��Qd`�@�*���Ŗf�<� @����"p�5M+c�|[��' ���,B*uk�l�-U^{�;�ı<��	x?a$>k"mᅗ�K\lT��hb�'��~���Ͽ9���: T�XÄs���:�<�	pyB�i�]EaE�qhV89���4L��(���#Ԙ'�$#<���p�� 7V�@v��.�ƙ��(� ^l����@2̄��̂����,0��<����8��<��*Ua�����Z�G}��SfP���]�?�U�MN*ъ㍻c2|B�I3B�ՠ��҂r�}i��L3؂�8D{ZwD>ʓS�Y{�@G*?AnE!�l���AD{"�'D*���'Kg��1(7z@���,}��>a�UT�a��9�\��hZ�L�م�k��b��=,��=�F�B�^���iN�Ik��hOΥh3&��`aT���88�R���B���i'0tp���˧p��][�5S C��q��8�g�5d�ڨ��g�QD��<	��T>� �D��r>�1��2�p�9D�b�W�_<I��W|��n#���>AǓ5ۊ܀�-'I���U��(��l����?Y�E�[��"6�<��X�6f
K�'\�Lq��Y�t �(��.�Jxq�G��~��p��`:O���~�*j��8�B�G�z`hL�-6$t�)U���<i��'��u8��Q\�)H7n�jT%��g����:s@�K�Z�Xɰ`b�%&�HE)6D���CH ����f
��3��5D� S��&	m�3W��>2͒��`fs�B� (i�UJ�"2Z]ɩ�Ɖ'*v
#<�a�gy�9����Ɉ;C� 3���yb�O6l�Z�b�,�
���ԕtў"~ΓT94]q"�>m+�L^��`��yX���UjL�@�B��ǃV2n���x�k�KѤ��h_+d�@�"0�"�O @Ǔl^����A9B�5`�A;O�hH��M�x+��R+o��i�!2X*�Ey��'��H�SCHL�2̆�k���
�'���Q�W6��@���iʝ'��-�S��'��y�'�O`� ��,��*�F��D$�$Ɩ>�Jyh��К^�&�ۀR����>9S�3�������8VY�&E�]쓴hO��'���p�'۶�hx�
7s����
�'6���(|���g�-d�>�;���:Or%(q�%P��B�K��(�5"O@��a��U�����#f"O��ɲD�j�j�zφr"t`Q�"O���� �v��P�vcA?S� �+t"O4�)򉗳-��p�2��4j�T�b�
O06-���|Sf#7m6�$��ı8rr]�
��y"��lY�����6��뗵P��"OX��)ްa��`���V/<��P�A�'��O��%Ȏ�
t�0f!I�F�t�z�"ODPj��SS���@ꈷO�9�Q"O������m;�r�ɍ�=E��[�"O�A�NҦw*L�HC�3ǔ8b#"O�3���/�:��?/��@"O �9�ݖs/R)�ओ�:
n��"O5�ƉvH�D A���Lij�9�"Oܢb�t�d�)$�1�������@��I'��L:P�-κb������3?92X: sb$S��YV�a�N|�<A�C��+ﴁIf엜U� x)��x�'��?M���8y��iŢ�7蘸P�#<D�LZ@��C�XQ��e����f�t��D{���	&
z1 �dy�K�*I�A�:���� �GM֧,ׄ�Z�kK4v��9wW�ԇ��')��"��E\��ej�4ވC�	b Z��F�@dy���)1aPC�	3���C���miҘJG�P �~C䉹3���ke�Im �|s���gDTC�	/'W�P�M�>;��б��;C�G�����:R$"Lz#��#6*��?�'G�H�u?a^w#tR�E�fT��색`����hO?),�J��B�m_ ���/Yc��7�S�� ����P�<=X��C�F�����'0`y�'h�҆�`S�	i�@]�8��a�f<��|�g`=�AH}�u��8??��CW+L!!���9<r\Y��D�Ut�L�#
ǟ /ve��i��P(3 �9a7�MbtD�!1RT��4�ĥ_ʆ��gM��:����hO?���$�� ����D/mb��Aծ%D�li�0V��a�_=�X}q0Ce���I1.��0��C�/����&5�PO��=�~r5��w˒���Ɵ_n�Qv�YC�<Y�C�7=~�b��!�N�ɱ�~�'{ў�'y$4��`&��G���xÊ�.#\�G{r�>��'�8�ʆ�ك"I�3�J��Bm4S�,͓�ا��iJ2d�9���&!����]�(Dy�鿟X����$2�� bR ����V)8D�����z��偰M�F)|k�7��p<I0�da�i"5�@�f��Ua�K�g�<Yf"�_i\ d�:\��1��g�'؊�[F��Y���)�I��j���l��nm���>Y�'J�Y�����2,�
�U/O�P���'�&�¶k�W?�p�#��?Hъ�*��$�>���m��:&[,D"E	�\���m!�'�aE,�,�����Hm`{扆�~B�)�'/��e�A��!������I�N��ȓ���SC�����8�eB�8�LE�'���n�`�ı~�E�|�'H���Ӥ-ܭ7+�����ȓ,/�u˷��>y��1�1��6.�%��oܓ�~��,O <G��x�Zi�A߃m�J��v�O��=E���A�*�2f`E�m��PB��;�y���d����iD9R��+�"[�-��ػ�¼<a�'2�Oq��Qhֲl�3��<������v���?O� �a�.(��"��b�=���&�$<�O��cM��D)���˒R�<
���0}�6O�b?Q�qI�1|��|���͢����� �Ij���O���k¤�zu36��7l�X�O>!���D��.H�/�nt�Q��$n*tR#F
�O���D��x`��� u�aP$��6��'��m�OL�D��R���1 �[<,�R���n�Tx��a�r�<�W+��{��!��8�X\��e�bܓ�M��3O����ɷ|���M�~QJ�2-��"��6��\�'���%+ғ~� U.�(4� C�x%���ԧX��y�]�D%
0cܮl�(9����=��>��Oa!���9��E�ԋ��	6�`�"O�U � c�B����~�z �!�Ia�O%�谆���`�����v�����'�,b�@Y&1͔�Y�Bǀq���'��SBGN>}`j-y�GMh�|R���'�D ���{�m�'�)L���K>��Odc���<Ѥ��(���@1L�T�`�j�V�<a���2e���Z=n"�t���S�<�2i^,)�x��D̙9`����bCZQ�<9�iƜ7�x���<s�Z����T�<a3��	���ڑ-D r<��iPW�<���ƚ�d{��=A�-���i�<��ő\������x�Pe�<� � ��Ø�����Aݴ(�I�2"OJq��&K�#u�`qϏ3��"Ov��M(Ap<��GK�0�2HC%"O���G���sM��8?��c"O����E�,v��3�a�%�q��"Ob�ŋ�+!xș �D?d,�W"Oh�Z4}<u��!��D/����"O�� a�17Y��Bd Z�]l�Ё"O���)7^i�}p�\�Q��%�0"O>�ãR�
��IY�u* J8V!�D����D!u�
�o�����
"O�TsA��nV<��@!�?2���S�"O�Ls`R�TXcW�ި-td��"O*e���T�j�9(��Z��[&"O�*@	=�pt��C�%B2"O>����,Wzexr萕:�<S�"O<���엁I�lm���E�x$%�'"O�J6�ۣT�m@�eF�-��i��"Op���^�r�a�#��JUj�"O*`c��4|�`�q6���P�̉G"O��j҈ØSA*�K� �p����"OM��H�8xv)I���c��y�"O\�� �L/$(�UC����(�"O��{���	Z^� a��*zJ����"O(KEB��j�D�����;�Faa�"O�Q8��؄h��EB%�n��yQS"OTp³�S�Lx��S�&�2��p"O����DK�V��'#M�c�XY�3"O�}� @I�E�܋���m)�Y	A"O&4pş�Sr��S��>�씒�"OJ����
"���V �&�|�cp"O"��c��)�h���Ϛ�vG��)�"O*t3�	 ��T#殍
h)�)H&"O��l�:�QQ�.֛B�|�"On�T"�Y�X�����oK�5ia"O֌��j��i��Q@���(8��a�"O�Ѹ ��	o����KB+��}�"O"����ϑN�P�j���+$�R��"Oҭːʏ#��@��
#ܺ��d"O�5��R�i`�ᎉ�N�Y�"O����@7Z�Q#!���l��"O	r��0�0bJ��B�I�"O���㝉sf��qJ��8 ���"Ox�GO�l�ʑ��*X(���"Oz�&�2�h� ��GQL�`"O|���T�U��P���� R�"O@5 jV07�0�
ƯS2[�|��"O���
F�̔)�@�"1H�"O>H��ҥ��!�n�+���I�"ON�!�+�����;i
�q��"OL�T/t�$vD� w��Jt"O2ܱf��g���2�T(Y����"O2�2���P&�݇}�V�� "O��k螠[���(0�� �lh�"OZ�K6덝�d�ڃ��'b�$�`"O�呕,��S�LI0��".��h�s"O"��#i��~���N��=@"O��hCR.Y<XwZ�Lm��i�"OV�R蝜@V)Б���L�έ�E"O ��%o�%}�� ����rp�"O��6h��;Z����%��la"O��B锳2� S�ڹM����0"O�X�*��|�(���?Q�Y�"O��K��ԧE�%jĬ��s"O� `� u0Rh������2Gv�ɤ"O<CŠ#J߼��cČ@+Pp:�"O.����B/}c��[�A�=)N<�"O���]S6,Ô�Vi�x9C"O���D��	�X1�c�_���*O@yY��L����2�ӷH�h�Y�'�Ba�U.�TX�H�b�C,<l�C	�'�2����zH��A׶BPh�b�'WZ��)�И��Q_j� *D"O�Mʕ�.R�dx��A�mK�u"O�ѣS�@	��Ъ"F��|]+�"ORe;P�B}t��������p�RC"O�d�RGϓv�DeB�ɛ�O�2�h�"O܈YG�
�R�� ��^�j�"O^�+IU���*�d��>|ze��"OV��7'V�:W�Ih��@���q�"O���.���˧eB O�JAr�"O��Y��Y;kWĔ:sJ@�,�e"O�p��lE�F�`�
��M� 䈔X�"O�H�PG��M�̐f���"O�P#RE��ThIB	�*ْUZ�"O���i��=9m:S��p�	q"O���W�B���S�{�J5@V"OtQ�"�-}��$	�2'-��F"O
遦�׍3Z �1�M�D���"O��O�RI>��0hG>7Xm�"O�!�Qn�,A��iѥ��@�B`"O��xb���n]�刯�s"ONxYT-�T��y��W�v�Ӛx�'Ԍ��ҩǍ^�	�E�>4a���"<O|�`����ͳDC�e��pA"O��q��0ג0��R�'����"O�=@���%����l���"O�mi&���o�֤���;1*�"O�3e!�e�"@��ƕ�a��k�"Op���_�p@e��R"�R�"O,��l�9:��QIB�!`A��A%"O�Թ��۾��akǹI-���Q"O�P*�g�?h��h��b���3"O��1���2߸�ɒ�� �ܴ!�"O����_�3�ti�����$U� ��"O�P	��3w�T�S@�� �(4"O��s�P<7���ۜ?/x3"O�����Q9߂P�SjA#dV`@�"O�Y4��lR�<����*�apf"O
���������Wb�U��! �"OD(�MT��l �#Z��T�y1"O�Mq1����~H5��y��;�"O^��W�ߋ<��	���K�6�.�A"O��H���>[t$�������4"OA��H�ղ�ͩn�^e�"Oȩ�%��3�j2�J,1h<��"O��ҷ��=���K�<�x�P"O��ũ�Q1jX` ��"���"O �@J,���)��Rm���#"Oh��  4"��Y���١$Yh���"ON]�Fb�Q���t�. \� �"O�c� 9n������"O��B�o
�4�a�ĭS�h�P�	�"O�� �D͚B�RP��.��D�$�x�"Op�ta�&~$�is�܋y�����"OҬ�5�Bp�V�9X͈"Oha����E�t��a�Zz��"O��2ER�<�n\��Q�B�2"O� �ٱ�,_=w����uJ��+�"On�Rp�2V��ixvM͋!*taI"O I���U�(��d!��4�R�h�"OX�Y�Z?��ɱv	'\T�zp"O3�$� ,~�1�JO�@IȐ�D"O�`�� Q�8��]j�Ɍ�.*�Pt"O�A�"�.^�1F(��K�<�"O8ĻC���7I.��1.#Z��A�"O�xH�)�_C�X�1�N'C����"O,ib��%f�	R�D(� <h�"Or`ra�حs%�y ��j�̅"5"O0<ae���]�e@�G�y��H@�"O����nI�v/:9g�H>F�z��S"O�xY��a>�|�v��!x��x�'"O�"���?;�I��&P�%���"Oࡈu!Ֆ4i�02R�@-L���b"O�Ir�"�,Z�*�*�4�"O,�1��
�(� ���¿o�
��"Oh�k�)W�j{܀u��(�V, @"O�<��#u=����D. a�Ӟ>i���iJF-�M+�G�0��7b�*x2!��K�%: a�Ȕ�=���Ia� W!���tġ�a�A�Z�`��T�X!�L5%�D�)QM u��tMRm+!�d�FQE�,O�ΐ�1�P��!򄊖GlX�c�`���Yi��1i`!��Y�m����f� Mr��6���=R!��D ����,K"�8�\64!��>Bʽxeh}����-!��5@�j�"�'6�: �#nM9o!���¶(D[E��17F�9i!�$F5-��,`���|�jR�ǁ?t�!�DR!1���8��@.�V�¢G��]��$W3Qn�0����-��P��/O��y��Z;\���hS)'��R�K��y �#Y���#�$�J
 ad�>�yRJ�oTTP0�р%�jfޅ�y��1 �N�c�.����a� Gܷ�y��K<2c"	��U�����(E�yB�[36p�a� ǇM'�a�P��y�m@s�K HBIH�"HN!���[���O�1�F6?
�[��Ԧ8�u�	�'Ţ� "K�R��BV8b��xQ�'r�����E�4�ġc"���YB�x�'Mm;��*s��XB�B&� ��'��D��d��2��1,�3|,)
�'Ș��O��L�/��
�9�	�'(��󡉮K+�8 �`��c
�'8$H�`
N/���(�r0qX�'�椛���� I!�B���k�'���j��A�.��͓�MW�t�9��'���1�J\[�q��K��r_����'�B�q�ؕmR����b5j�'�BK��\�a�Ճ���`I�'��C&�~�|�
d����~�x�'I�hR�`�nk�!33a@�H�$���'c�x�u��GT^���X�>�N���'F�-�w�� ��X���K��D��74Ƚ)���6� (r��G���ȓ���:co��JԼQ5�3�Q�ȓƴ�[�G�0):
��e�,������:[��G5rB��OJ?C��%���°�$��&M'�T�3�� ����ȓ��b'`_2g`����eG(+���S�? :X��C��DS�m+�)3�|�j�"O��LÒZ*2�D)J�Wq,��$"O�u؆BB�c�F�IHP�T[(��w"O���PiK9$�J���ǁ.vw��K�"O�E*�����A'�}�2�G"O�ݘb��4��Pp�5�T3D"O֘A�E�դ�7KӒx���s�"Of�z�-]U�j1*�D�pF"Oдc�/ݞc���a�K��e~.�;�"O�j��W-0��U��E=H�Ee"O2�K��Ư.
V��؁)$)"O^Y��*�k,,aᕇ�4"j�9!"O�����P��h GF�x�$��"O*|HG��\�Y�$>���"Oj5�3�Qo�&i�Cӹz*�pi�"O����N�5Mz�s��ٻ&�da�$"O���M��]>(�dԵl��j"OҔ�&��?x��gÝ�o�txR�"O����
 ˚5`C�*s""O2|�c�@�g���+^�,�J�#5"OD�'96��u�D)��$Ǹ�X'"Ol�ʴ�P�1�
ŚX��(�"O�#4$��B�Mk�U>x4��q"O�8��+�X�[��ǿOsrd0'"Ot�'E_�cS@8�o<
Y2�"Oڰ1s�ӝx��p#�˿  �`�#D�09�m
�]����Q�Z2W����7D�h��1|x�y��A���3���l�<���H1p����Rb�vmӑ�q�<1a���:��Dnd~H����l�<��^J��4 "g�*"��n�<��
��1��@����1�i�<��ڱ ưH�āN	58�$�vKHc�<�c�G*lk��V!�mJ�,C#o�b�<�#�D�*J����$�ц�[�<��͏i_�
��[9���6���'�)�aCzYcw�7iq�t�R�s��\ۈ�ǥG�>۸�3���8�|؆�}D�mc�B,�Q�%�ʧbt恆�xL�0�!�!#*�Ź`�T�~�D8��&2�%���˺t�������9�C�I�	7b�2-��J��Ĉ Ү|�C�	�~,X��P�F<"",�;v,�2��C䉕FV��1�ځP@⒌��(��C��,h����'H�k�XQ���@H�C�	=s��!�,�˳�K?~C�Ʉ6+���mHF���	�u�(B�I�v"@bP�]?Q�Ġ"FB��6��H���Έ׸�{��5	��C�I�#����C!E%jd$A *��A�C���,Z2d�<n�D��BJ�tC�I�(v�eY3�.(h�7�aʞC�o#2�Kra4%���kd"^�*"�B�'5�d'��I#�Ũv�ݘ-iDB�I�S�ry��F�*�X]�H�9�0B�&$o�y0�ݿ]��8Y��L�S. B�0f�n��f�R��(,
�c�2B��&f8��r@�JN���o�c�vB�Ʌ,CȠ�qE����I�K�y�RB��)Z�d80���{�t�J��0v�B�I��*Yc�D�<�dyZ�O
�OW:C�I5% |ABB�?�h1UF����B��(%#��yw�P�C�p�:�ԸG>�B�	%\E�Њ�`ʊ/�p���ө=i�B�I?x��k�� 9[:Z����N9�C�)� 4Q�ڵW�,$��'-t�6�R�"O�lQ��U0[�8U�vŞuӜ��"Ole��ǜ�T)6�P,�>�Z�"O���Q��:dY��bv��7Ǟ�:T"OVX��⒝�|�7I�&��<�!�䁯<d��Q��1:P aŇ�7�!�dIx:hJt(�/2�<�J�ę'Q�!�dJ� ��r��f�)�@dς1*!�$� �4-�E�k����5��A�'��i�ƋΝo�(��'�Z�(�9�'���zVN�:y� �R�F�6[Sj���'��y�d��7!��P�`P'� �*�'�Z����9!A��鵫�T��'� R��)b��e�����'=5ñ��)&sbEH��[�$������َ7�H�|��-_�Ήj���!>E�}��ny�<�t+�Ja�\+��$<%x�PF���\"��d|qO�>����)2ji�F�ήaȄqط�;D���*�df�]c�B@�mx}��F9}�H�&���	�Yn��(2��-;����b�E�J����"W�~��j�A� ��&�Ĝ-�fE!�ύ#�ye�?&�\�钫�+W����ͮ��OP�3ҊT����Ա�"�?96 !�*�yu��(7"OV����&"���O�0J�����O�	aI�����h���ئBèY���&=�d9��"O�L��ߐg�"��%mF�t�&���x�+���z�AB�B�b����qi��5�y"ٹ@� [֋�%n*^Ź�FQ��y�G^,g;���@�w��\;"BǇ�y��P������7:r�m8r!���y2��h�A�$J�#3�@��ǌ�y�F����)aA i��3�E��y�Ɵ0].�bT3= \���lߗ�y��/j�5(���6�B�PB*F$�y��G�B=A�$&7$��s�����yB`Q�li�x��͟/�D��"掻�y�/A�0��h�L� 	2��Cؔ�y��ܲ��\xF`^(�����ּ�y���(5QRlRʗ'����h߁�y�#ӧ�
}��	LRȠ� �U<�yLq8�#M1����׭��y�BP�4�M{l=3��1@�O��y�)�����0��+d�$Ӥ�U�<�sf�j��B�I-m%Li�2�
W�<y0��l? L� �̩�c�o�<�c�I'e�F����ψb��H�skLA�<q6 �-=#�je��z�6�Z�f]B�<���@��	����s�z��C�<�3+�yӊ��F�It�z��{�<!�aY�{Y��rF�P�HHUgPt�<�SJ�60�]�_�J� C5��C�I��\9ae�FS�qE� A��C�I�-T�D*���Y���Fj[�xC�q6���8��*@-M<[xPC䉢=̾qhG㏆Rڹ#4m�0�XC�Q�Xy2WO��4��4a:�.C�I�<��Z�A�A�����BB�ɰ%j��Ԅc��M�D��E.6B�I.B� `���5�H���m��C��	y��=�f�,��l"Ț69�C䉖9(|y�� -"��Q3l(�XB�8B��d#�n�!2��� T ` �C�I%\�n���	]:S�h9���� �6C�	�4"� �S�J2I^�0��MEC�)� &��Wh�����ȗA*��"O&8��� �H��A�
f�"O����ȓ�������		8�^���"OA�s�NLƼp�qz����"O�yk�J�&iF�s�dX�U�*h�D"O�(���و�`��'�2�j]��"O�u0��Џc���P�r�B� �"O6P��� >�Z=�򣆹
v�	�ȓ"|YZg��r���!AϞ�����tTh���ܾ+d.�9��F?to*�ȓIV �NC
�nH	ԇL[BJ�ȓn������K��S�l���ȓbu$��e��u�l�צ�9������T�bK�1o��%S �F4W8ć��T�1!V�6�Jƍ�56����?�B��g����j�H�0q�a�ȓC6���D�=�ޱjV��(�2��ȓm[d`�@��uz�� Nܷr���# UH��>�Tb�ÙS�ͅ�Iu���b�*Ff�P�AǉD�v��ȓ*� ���,�w��+��,�ȓq�̭�R�Tg��ѳN@<7)l|��	J}�gö1b��i�+ף�"H��
D�yr�$i��Z����� ���3��ǪG��OSt\�	F*̔���m[��y��
�*�t���:Q��@��?�1�2�S�O<�jb�ĕU>�
rg��2%9V"O,���rI���c�d0������� _�a}K{(���B��"���*"�N?��>iu$B\}B10�X|�t�K�TW|�a�K+�yr�r/|��%�/Ut�JV�R�(O.��F"�'~��1ÕoV�g�x(x�-w���Z��zv��-':pbw�ϭe,�Р�eB�O?�$��R ��9v�Ą$�L8�D/%!��M�a��Y
6�	9�ZXAV�y����0 H���D�!gu !B���.t�y!�%��p>1������=�c��a��A�'�!^!�*n8%���;O�N�����J�Q���D.k�O��g��"�\�5�[�0��X��'�B��S��2��(��Z:vU��o�?=PV�"~��4p<L�qf��M�T��-T�&�
C�	�U(��C���5U`T.!'����n0��I�f7��!M�g#�=+¤�$M����ȓL�8�;ԁ&�!i���!�
����A�AkG�M���J���(]�DHpƥʡlϾ8��4ʓB<D�zK�P)�� �x����;gu�L*��Żn��a��F�
)�ȓo'f=�Æ�aR��%�2dpH��Vֲ:i�I�d��B�M�-eu�XP�����r\��e����`NϡY�,��K?�z�H�T�<��W+ܛX�$��#�*d��iIխS��y���rZ�����Y����,��6�� �R�pf�q)��(�O��9��>	q2��ȳ�(�rv��!Ư����0��J�>o���GJ��<I!���j�@0-�V��tb�lž�GyB��9V�I�6�Vhz!�˴gU؅��ML�t���G����j�(�U���A�'��Бg�G�FT��Nq,ά�ܴ:�*��'o��!G�M�I������Ɛ�Db>�6|�4��q����\�ϖL<C�	�V�ȱAB�.[`]"�״C���8�j��(vѲ¥%�M�F�v�T�/������$�5J��u�fC
-]�pJ09�OxZ�O �r���"1�hã吖"���ATJ��e��I��I�:VI/_X��y��*7.*q T7��1:#j&�7-��!L�!Sm^ 5�p�9q
�=JD\�f�_.fMD+��h�Z�s�'��܀r��n�O?j,��;�'��I�?���@���6<�82fE���O�Z�Sc�T�ed�bb��b�J,;�'Ԁ4�N*'yr�@1#�6^���5	�u��:�W1�7��05�>��Ⱐ�J�%egܠ�`-ٸ*�ԁ��S�? 61�tJ
**�B$0��\�Gޒ�xi��O�����*E 'Z�m)<O�DX!�H68���jo�D���'�b�:��2�.=�R������a�8gpr��Ea��c��E�	�'<�juϖ+g*6�c���w�A��}R���j�*�H6ռZ��#|�$LM5j�AIr	�:�xy[�@�@�<9�F��1���c��S;+��l8 �X�n�u ���>�8��h����^�Y�w��<RN�h9B��D�!���o��P��F�/3�!i�`-���Z�m2�u���'TZ9z�*Z?�����=}h����'�[ǃЊ������k�F��'�b�� C��+��l�ŧ�?��9��'�J��Q�Z�[D.Th���?�@z�'oh���a����t�^��\$�
�'~^jAY�/v�9@��Ƈ8Ÿ�'�����(�oKpt�V��1]�.X9�'�D)�EQH���'�
cD��'-�a9��P8������K���''���������NI�Q�\��'�<��N����PR��D��'��|���[�|��H�e��8��'TM�R	�X0�LHD��9�'O"+�20�v��F�X�?���J
�'��̀CE�9(F~T�@`�6i.�B	�'� -���&4{�W� !y��, �'���:��[�h���3�˼)���
�'1�� ��^�\��X���+��qY	�'��m���G�]p�	�ń� 7T���'%(�P�b� �������\`)�'�t�F��LS�aYu&�t��Pq�'|��(䊘�sd�Z�/�6\ɨ�k�'���1��2pr�9�͞@�`٨�'e�	�Z	yo�]� �ˎ@0��R	�'��cň�,w;RU�0n�<Ɣ�	�'Q�xF�V�4�)��Í(S����'�H}SV�wV4 �# [�#m"�#�'���V�M22x��!��7%����'qTٺD�j���r"�,S�̳��(D�x��n�1���pwK;�0
��&D�tʦEپp>��:�鏁p�R��"f"D�4�0ǋS�d`ئFk��X���@�<��\A�(�j4��Oܞ@!K�A�<Y����DQd�B�J��>m���p�<ѦdR$=D�|���W����&Po�<�7Ӆ/4vM���U�E:�)�'�A�<CD��R�b��!���!�$�C#C�<��O��0� S��X��:1���G�<!�%�1<�H�2�ɉQq6���~�<!f�S�^,�b���U�����{�<!�\9��-��
I?k� q��(�O�<����,'2d�C��:]&��i�r�<��.)\�ֈ� �>y��	i�.�d�<)G�]%(LJ��6�ž2�v�۔��f�<)&�%r�XZ��EbT��i�a�<�3 ��rD�T�$�fE��j�X�<)�]_Zz�(�FI .(�����~�<Qf���K��L)@.X�e8�tP��m�<)Ԉ� P���"��D�$�CU��k�<vi�*4I����	".�,�S��b�<���[�p�Hū��b�����O�^�<�
P��A��l��@��Q�DU�<�A�͒]��E�ğ�7�t�a��CR�<�!���b��QUJ�"%���)�M�d�<)�V�J�`�uO�#��!�!af�<!�9�T�� ��%W�FU����j�<� �Z���t�� n�)\%�ܐe"Odpʦ��_A��2���r|ʆ"Ob4Rׁ�D.�}�L����c�"O�-�w�-J�ٸu�6R�T��e"O����C�\��}A0���S��؈"O
d� 9
i+�F �PXE"O�T	¥̠�fe�W��l\'"O�Q ���/�\Ȑ'�Лv���"Ov0`����47=�0$N#��m��"O�)�HT,!�jŁ^����"O�-*��ǷM����%�U.O���""O0��v鏣 ��c"Gκ5�x�P"O>Y�ToT\*	��8�rt�U"O�0pWdT!)�q� ?(]6�&"Ol(
����)kr$��)A�4��"O�*Bg؇$Ѻ��M2	�51"OPU�E#������2� 1R"O��(/�h>p���H;,ލ£"O�q�P���+����%�= T��ɗ"O��H�.�o�����R�RX~(1�"O�壔X05��,���D($�p�#C"O����!�����Ht�<��"O~aJE!^�[��hnh��"Ot��rK.03�ؗ�?B���"O<�j�e�
EҕRbj�1-6:��s"O0	 �8	���*������"O���3+�{3չ�D(u���i�"Onl���%q�t6g�F�
�zf"O�(��ߢjZ0�eh�2���"OB�¤���Sv	�ow���"Oi�F�,p0�`ѩ�%�"X1�"O��+��U�)�|%�s�]��젶"O�%p��, ȁ�h��`�P�"O|�Y7��A. Q`�ޅo��`�"O��,O(H�v��`��W~�S�"O�s!�V��V��@Q�>ƀ=�"O��	��˳�1��O�.H�.A)�"Ov�#�A�a���� °.�����"OR��Д7VX�as�G��T%�"O.t�W�6R\��@���@�$��W"O�Y�p�=��+�Dٜ��"O��h��ݳl�<�zS�@S�8� W"OT;��@�&�x�	CKź���H�"O��h��34�pf���m�"0�6"O����@K>�I���ۘ4��(�"OĸȠ�;[�*A�A.s괵��"O:Q	�N-huн1u�!O���E"Ox,�'2Xq�@��Β�Mn�T"O&�J -{xV T�V�( ��w"O�E�'����3TM�- L�3"O�PqdC�>7$4y�Mo�ZE"O*��u�P6��Q8��Ѝp����"OX��F�̷T�J���!Ԧz��Œ!"O��h��^g�ak�]�f���"Obe^8X�k�+��a���N�H !�Ӌv�*�A�`�G�Y�L !��ޑy��)АA�48\=ӗ���3�!�䈌����!I{I���ظ@�!�$R�}úuQ��2A7��$ĈE�!�$�.@v
,S&��C;�� Uc�y!�D�(8�A�#�خY/J�����!���tJ�{T/��-����3/!��K܆���*sҪ4���DF'!��2-e���2P<`xA���Z>!�� rx�P%	$D2g���L샵"Oz��/o52={�S(d�X��"O����Ɲ�1Vf�� ʘ���qq"O6%��n�_���!�a�U��"O:\���m�Lݲv ��L�, �"Of��p�T�?�N�Rf�T�\��"O��A$c�
/�uI�OR0�����"O��
�牠C`D��bm	�u����`"O�|�l��7#H��B&L�&i��D"Of�3��HP��r�E�5j�"Ol���@�@4�}�5�՚~[p��7"O�ɒv���<�F(	L��PC̡#V"Oj��iނH���(�eA�!F���"Oj�ۆ�U�t~�r5��[��ya"O��]�EAp���^�>�p�"O:�R��δ���cUI��� �"O�)� �;B��&�� aq�Д"O:�mO�%V�yHOԽVed�;"O��i�	�4ǐ��d/B0U�-r�"OX	xQ%��R
�̃�Z�&��Ht"OLJ�K�'YPU
!�D9)��Њ�"O���.0p��	�w�˃5�
pj�"Oؔ5�9;�]X%h�%��P`"O �C����v�-�ҡ{1"Ol�$ (q�ɂ�'��6���!"O65�e�ƉO4���'mODL�s"O��x��J0��S\�;�[`"OLi�C�-8�py��*81""O2�;�l�[�.�"B�Y>F�|�Z�"Oh�ʅk�?]�5�V.�l�nI"�"O�H#�K>3�t�1�S�l-RlS"O<���/=VH��,� `{"OD�`�k^3KZ�2J�T8��"ORL21�;$/���"خɓ"O�Aʄ@K�D����9l��1��"O��r��5,�1P���!"!r1Z"OPh��w��Żc�3\,�� 0"O�l:���3eZT��O2; �y��"OTћ��Y:9EXM�Ǯ�Yv�s�"O� �ĄpF�)ŭQdH��"O�L�UN["D20�L�c�6)�a"Oh�����5lL0�!hM�v�L(x�"O"�I�&�36�p:�HU .c�+&"O�9���ʝ|i�)C��5<��5�R"O�X�6̉�-7�%���Y!q2`0�"O�Q�PFݜeM&�*C�2�5�"O��p"W3ʥ��nE+���"O�A�G��DS��ڧ�V6R�hZ�"O:m��C�B���1��B�^�us�"O����!��yv�m[u,Ǯo��	�"O��"jFkF���K%?��ajD"OB�CgV�H6�BI/ �(0�"Od�Pg*7 $�R��=9�^���"O�Pk*��]�^	"��Zy��m�"O*�9���Ǟ�{���i!23"O�2&��E�0���n�8���(!"O.(��%���2�'~�x�"OD�B�AJ$<k:���N�wu�m�V"O�M��#�,����Ύ�=q�x0�"O:�#���cHFͫ���+
�z1�"O�d�6�k*���F�m{ �Y�"OBXI�j�'e�Q[�eD�BƤ��"Oh�Ah%��p N6J�P1P"O�a`�L��4�0�js��*-
��"O� "�����l7ҽ( �� D�B�"O�04�M�DC�t���!D+,�r�"O�Uq+ۥw� �����p!"O��'�]��|I�.��Y��"O���mT<HZ�ر-Ւ.
��(6"O��h��O���:E���jU��"O����cA`#�e�U��7'h�:"O>�u�FJ�%k\-n��"O*�9E�~5�d� ��i�Q�"O�a萠G8����`-M�mj4 p"O��Ҭ�"n����,O�7�T��"O�w�J�3\܍�m.��130"O���G��m~��M��Od��Yg"O0,�3���G�Jt�F�QJ	S�"O�UB��vu�;�-�Vt ���"O���'���~h��aw��B"O�7 /�d�hUn�9[�<X���8D�(��nK���	���'3�uc�h7D��!��J�I7�M�Ka����)4D�<+'畝��)�&M��愐�4D�b�#�?H]�EiFF��@7�9D��"1�Z,ِɓB��%d:�Xsg7D�<�戣�a)�+�r��#�&D���1�قZd\��V��jHHLBG+!D���܈J�8�L�F�PLx�/(D�T����R�j��I��8�*t-D��Ѐ�7�����"��i��=Q�7D�b�&��5����g�m�̵�b�4D�X��a�9��ةqGZ0,��*��'D�$ � �&zճ��}E�Uh�B#D��Y6
��R>�2"�M1�\"B D��2p�(�4�q��0�ؼx%)!D�4��I�>J�X���H�C�H<D�T'�[��p�!p 
�LQG)7D���qㅯi�TH#J�D�����/)D��.  �IR�s�q�T�&D��`�$�N@��)1e��w�t}�e�#D�d��̵pV��tF�D�a�� D�T14)�*;lYC�B�,LQF|�� D�0g��
>�����k��V_j�8� D�X8� ވj�:%��[7J�(� �>D�ĚsE٭����!Cu(�c?D��ʀ:�4X��l�0�rd�0D����"�n��2���G�9��o-}��ā���E�D8�"mA���'^�\�a.U$4��d��D�3n�b�����P#<E�Ԍ�/<j��$��s���U�P����V>�Eo[W���C4'F�vm�����=�I6uQ��O)DѺa
ԑ2���b�O�gIx�rN>r�/�Sܧ ��p��!�to���͇g���'%йEy��r�p�-$2(}��
	��AG����P	+�+�p&�"����2�a�-�p�'�a�4e.(a�e��!Z�-��%M���'3��EyJ?y�2oX8J�����W z�a�5�����(Oq��Ԉ��Q�4�p\Q7�Ex�I0DZ��a��7�'"6�Ԛ��O�](���U�]�J�,��	-y�"<�'D�R A���;��]�U�O�<��b�u�r�:B脟
f`����
��'��A��%_2��OJxѶ+"���lӅ�KѦ�X��^�*B�C��W��'٤�+��<��!�Y#��K<�Qcs���OjHt2eG������U"�vQ[*O|ts��哯'�&賧b�;&�ĽD�Q�W�z�D¾�(OQ?�	�n�<wp")ɐ�#.�04ACO�~�|2R>c����@�Xԩqϊv�f�Q�-yYf��(0�)�d���xc�^�:�����5��:�¢<�}�6a^��,S>a�(exq.NVy+p��(�� hœ!NͤG%"�Yw���[�0Q��'��HFy��	4�b�B�m�3{3&��� 0�DGy�O�
!�sHA�� l2A!��k���؏b->�O�']8�@T�T�V9��S	X�(���
 F�C�L5�O`�"�Vs2*�C��Axx��"O�	j��\*!_����J�r-9�"OT�#(Y�u�I�`G@*}���
@"On\P�9<�.e�,H?dꕒ�"O05�t�	�+��C�M�JSЬ�5"O �Zg�މ?��Ҩ	�g F�@�"Om
RWOk�-�Q-�t@��"O��Ȑ�5��e�SK�?*��ܠ"O��3R�L:��v
�mD<��"O:�F
ʹp��@"*G�uX$�z�"O"|9g��9QD�8�Ň	|�ZZS"OF=��.�% �%���VN�^D2�"Oм�fIC(4�%�IдR���V"O�\s	QA�y�(�.�Z�`D"O�T�W��L��ɱ�D3��d@�"On���>��U��%�8���x"O�58�a�7&�Ȁ�P�F�bg,xS�"O��s�/[�-��`�4���tR ��"O���`P�Ǝ�HEK[.��,t"O����'{N�2���K�ܠ�"O4ӕ�K�v�X!+�5KZ���#"Ox]�k��~��VIP�A(	p#"OB� *\�QPP.��!S"O�1�o@h)�y���צ@�Xi�"O^��)�0�L����?J��[�"Oj�j�Tj��2R��q�F��R"OB�MO1�	(��G-e��д"O$)!e��j°Ċ��T�P�8�"O��HS��}���虗^1H�*O��K��P�"� @Ԫ��,�1	�'r̨T��N�}��+�P�[�'K8t(��ǰ3Q�Afnۇh����'�R1�U�N�"�~`+F�X�[v�u�'�B�����D��_����'����@I

.D�@4�T0��'h�ڱ��W�p�G��q
�'�$	��`�3J�x�gjW���I�	�'2JS�M�[R�Z��Z5�-[	�'Lj�+bC��xJh�1�T�l�p	�'��� e��x��ыʏLI0S�'!����S�Qp��0�'ծ@�f��'��S��X�vw�iAw�4���z�',�z�HL�:i��,�'��+
�'  :R ��v��Fk����'��Y�lC�� �J~c�l��'_�z�	��5"�]��9p����'�8��v�!��8E�>\N%J�'��)3l
�fa���d�
QHS	�'4��)���g���oʠC~����'C��;�F0b�*h��+������'���볡��V�Ե��H�*�����'�8� V=�d�Q �;0|P|p�'�ZŠDM�~
���W�"��)y�'�|�3�DX%M�4�y��ՠ;��p�'̰�	��ZXV5˔�N0�
���'���Xǉϖh;4bR�}QIR�'
y���0m>���V8b��Mr�'T�	S�Z�M��(�m�`�Z�8�'`6���\�l�<��a��7/1����'Z���V�u�6tK�\�)�)���� ��Ù�G�,L�V�{1@�;�"O���FK���j�A�9v0`Q�"Oj��7���F�� RV~x"O��z�$��,�``6*FI�"O8!ktΕ37kb4���>b�P�W"O�@j2�O#JS�E�a��5�>�"O��[�`�+" 	p����|��"O�-���8UWP	�fM/�,��'"O	�K�E�>���M[�4�D]x�"Ou!�Z�x	��R^����"O�m$K�h� P��������"O�("l�	^~�[3�ɰ#Xb��7"O�\"�� �/�xR��=(/b@[2"O���O�`n�����
=����"Oa����0p���u/�lvV �"Ot�pD p)���a�2<e�5C�"O�MqP�A�i?0\���?`f:!:�"O���$��p|{�c��@G^�� "Oz�qDeK���U��1^/@�:�"O4�
��?��4CP�VW���"O杲��U-��S�Ώe6��"O�x8i�#O�.${�:;�j�:�"O<iq�06\V\�`K�$�x�k�"O0h����*v�
��s�L���Ӏ"O��j��P�$�E�T�m��(�3"O�5�&L�	4��z҃T��Ʉ"O��Qe%#{������@m���"Or��ĥM�{�80����-��"OT�sVɘ�E�
��/ُ�y"O*P%��p�Y��
/�ذ[�"OD� 
�$]̵	�g�:?}81�"ORL;b��# �t}���%F[���b"O�]�dEb�k3I��w���q"O<���A�o�*T{��M$S-ܜ!�"O��brMʿH�8�B�=j�hr�"O l���?����e�H߲�2�"O�����t��`�����.�qW"OYj�.�2Iі���N�E�&��0"O|$b4dߗgp ��O�BI#"OZm�S�Рk����3�{�j9Q�"O�|H1����عw,P�c�py
""O$�b�i����4�L�9&���#"O��F���L��͑6��ɘ�q�"O`ؒ�+*k�&IZ�A+xea�
�'���ᑆj�`�h�f[�[�t81�'O���R��v�@4bb�6U}J�'�b!�X$�����YO�&ia�'B��b+�u��u�q�ҙX*��
�'��kA,��vb�]YV���R1���	�'l:M��F��	�e��#Z.��r	�'�DHˀ�h�����O
����'�&a���B	W�*��Oɻ2Iĝ��'E��"�$��o0�z9n!(����yk80r<����/x�d��+^��y��U�^-6�x� �9nְё" í�y�!s��̉c��$!���C���y���~p���셥�-�4 G��y2E+zp����S7!��H@uKJ�y����s����`��IRԱ�d��yr\�e�8���XH����H#�y��
�n��!�I@�B�
�Y��6�y�*^tX)�փC
L�1J����y�˗I���֏�-X�b���LA��y��6:�$p�6`$�unL5~r!�� �5;b	ĉ{Bl��K���"O�,�E�3��e+�΂ͱ"O���c��9�ܔ�6	O\�<��
�'6>%P��0�"A��"A�>yY
�'5^��PgW�#�dd���7
��EI�'���c���M�B�C�ދm�>���'���L �x�r܀�`�0^uV�	�'�4�ٖM %�&�qRdD�U��m 	�'/8A 6(G�yj�l��� �>4��'���SGʁp���IȢw�d�a�'���Pb�>73�Ԣ� �F͐���'�"e�dO�,�Vt:u���q�' j5�d/,%�̀�e�	?౓�'5��Y���}"�đP&M; ��R�'�h �tL�ƒLxP��#Ip��:�'`p
�dzvEa#�B�j�
E"�'$j�r� �1m�$�c�F�,�N��
�'+���A�
�8	.�!�� K
�'^�i��j�d�&�r�F�.@e)�'
T��X(SH��G�
*�X��'��\�%�)^�4C��O�<�J�'	*�cTmՁv Z��c� |�H`��'��E�SH 3mN��(Ch^�!0D%�
�'G�tۦ-ͪ9n8i�"EF HʬQ�' ���ѻ]q���$Ô`,�؆ʓDi"���@�MjU!L�lV��_*����K�|椛��ػR�f�ʓ�R!k�^�IH'���&�B�I�u���&%O�b����F\�6r�C䉔�& ;JO�J?�-���|nC�	������}�t���O$C䉒ijE��!W?YHQiԌ��C�ɯWaV�y�D�Q��x{�Kǒ�B䉏Pt��Z��M�;2��4lB�J�C�	"z�������H��$���ĸ/|*B�	�-�rx�6��)x��ġ��@$Q��C�	 $bl�t�O�3͢�R�C��C�#x��A�D��*צ� �C�3IߖC�ɽn ʑ�NV@Ut�`���>�^C�	��f�
��2$���T-Eo:B��:	f�%�gc�=���u*B+~��B�� #�tm�VgY�YweW���1p�B�ɨP�E"���=^ЪU�lމ�jB�+j������~rt�T���?�.B�ɡ/���YP!^�c��Ո��0|�\C�I%7�B�Y���x�HE�-+PC��7Z�k��Iw`�X���&�FC�� U�* 𤨊�����S�$4C�	�D<I)e�-n7Lr�V�8C�I�)���0���v2�Q{�c@�2��B�ɑ1�"����נ�Y����Z�B��T�����&l�]&I���~B䉕9�rA㊛�3�Y¡i�RPB�	$r����61bR�hCbA�i^hC�	>[�XLz�F�9�@uۖ��,)"�C�	�j�^�z��	OC*���B^�:�B�	Fp"�6���*���"]�b�nB�I�"����ǜ^�� �sk\4w��C�G����F#�u��ԓ&)ܒ ��C�I-x��yAP"�Es���S��>d^B�(v���;4�J�nI�cM
}�TB�Ig�.����1Q�6YB�M/HY4B�ɳf��B�P<[�b�a��J�}v�C�	4!�lTKv茜1�FE�fǛD��C�)� 6q{s�F
��u�v�%IǬP��"Oji���B8�n����/0�:@�c"O�ї=;[�k��F!�0� �"O��e��A��PX���5sЀ�´"O�\���"~��X�Wgޓ:���b"Oy{�J�V��(��F�F��"O�9��+޻`�<`@א.	��	�'�F}�"Y4&���ҡ��b`�'���ޑOp�-�͎�����y��'�V t,������?ɔO�f!q��S>j�i���� �xe�#`�2�'B�n��!���ʦ}��㏴au�M�ǎ�G�:��$YQ�2Ye���%���b�|cR��v�p{�b�a��Y��,ؼ/�b���N�$9��F�_C���� 	�\u�&�$Y���pӌ5$>��O�h���� �)��
�]X46�'��Ɵ$��l�'��8�d4[�ďJ���C&i<g�Tt��	��M�ӱi���0n�A���Cul5��Ȁ�V���5�ǖD�&�'�2������:���'��i�iS%�B�=�=�����NN�E�AIܬdR�t��I�#`߰��V>���*Ɓ�|���o���9�m�f�7O,2)y`�=G�d4��ܢ\����5�4�,h�W�H��P�2��d�h��Tm�.~m����A:�8�����?� �ia�X�'��(�����S5 �j����e�H�R���w<U�����O�#=1���+�9�Q�J�~L5��w�#��6�uӔ��E�I�	�?q�Sæesc烶i���A��N�e��K�GD��?�6��I�������?q��?������O�6�V�g��#tŨ�vݙ��L�~��G�v��0;l�9��Ԯ�N�rq"�!��"��Q�F~��;s�[eW�\h���)~-)a�7���%�h�q�ei
h%�O�Y���J=� ��eF�U�L-�ѳi��Y���I��&%?ғ�ēn12��#F�[n��c� � I*��O�ʓD����O�zh+F&[�r�$�Ag�M�/�v� @)���m�	��M;��&���OA� Ơ�p�4�Mk� �6J~n����Z��<¢���V8��'b�˺*�R�'H� ��mA���1�	d��2�dߓG����vʝp�"5����L8=�G,��]#r`x��d�|�����L��+)��`nF7��	��$��7�^t��d��"���p��z,��0�)(�	���d�}�Ú�&mrUS��Q.F�up@������wy��'��O������de!)��DI�<��1�T)9D���G�}������U.�tek�%��I��q�i�剧r�M���Od�D�|
�OHt�eH�P$:��GhV�?o<ei���?��sƤ�Z��]���&N�+RJ�m{��[���`Yw��z�i��4& �RT��}2-��-�`�kc	Lz�TK�һўI�vnOv(蝙�N.g�Űr�:��>D1�����10ش�?	N|��G� !t����Zl@�@hq��.�O����~}H���2�[e�2dK��6���p=���id6m�>!0�2p 8�	�C6Zá��/���S�a�&���O��4���P3��O��D�O�7��p���W+F˞��)*h�P �(�|8�k'j"�*��3'�&�t�O|�TJBǼ���r������6P$�B�Im4B�StiĤ4,\(SP�O<P�p�bT*K�̒�:��;%�j(��+|"�8�(�r� Pr�'�6�syD����; �d�p��G�o3�BC+�,- P�'�a"�̬N��=���Qx2Q��K2��'fb6��%��S�?�l8*�^����|2�Q�@�+? ��'�a}2���w   ��'��5�褑G��g�'Mb�{�,��kz|8��!Ġ��t�4F�-�"2K_�n���
c��h��A�z�'al�C����6�(�D.�&̐�1�\�Z6��$���X�L;�ֶ)�
(�GbD�^���@���0�'}"?᰺i��*�=i��D�P$�/�n�O��r��mh�D9;Q������ȟ��	�?�Yt����Pl�,U&8��'�@�~t��A��1�0�Z�r.�|hC��Rn�]��1eA8y*w`?��̉.���ݼP��A��͛ON��3(�K��	0��$�s�4�c�H�3z�`<��!��9S�`hO?%A�j���S�)oҚI`A��>�W�^�؈�4~����'$�>��y��C��D��p8�&�
2��ş(�	R���	G	�<dmJ�8#F��TNThQ�h��4c��6�|�� �[_����+-qn��p��I��1���?��Ӣ���[(t9����D�	͟���O����Q �3L��R�<f׾ ).�s��8����R�0��������O\�-��.����DX�Pn\�U���{�nuXũ��V�XC��Hz�R�j՛S���ز��D*�7�x	���Or�@�o/_�Li��mO4��ۃ,W6�M���
���x���ʟlړ%�ȉ5
:���*5�E�.��Ć��9S<��� H�Y�B�		1\�I �MK��iP�'L��O-�IP�z�GL�'�Z�*����_�$�Ӫ��f�Nh�	�0�I��h�_w�R����4d:���Ұ\p0)���5�d�[!�K�V��F@DY��Y#O���f�Ȇ��k�'(�9cF��>��{"�_�]���\H�(	���'�]��٭q������C�0�OXt�a�� UhgOF�*��]b/����Q�M+B�x2�'����O�8�{թ^�C�|�^�`�y(�'�ر�`ED����Ɔ?j���K�$�ڴ7����|�'n�W�|��*   �M�`���"D��bg�� 	_����
Ʊib6�p"=D���h4�= ��@��TI;�0D��J\�1WJ�~��w�ٜjf!�$��xLԚ�h٭1��0*�[�!��X9(8�L��Z]��2pcB�`�!�Dl��9Dm8;V�*�b�-!��L�S��iY�i�.�#O�S!�Ēi�"�%��� �����!�d�8���Pc���8p���b��!򄚼J`��r�6U��i�A�RG!�O�K+n�ЁoE�O�t!�AU�b6!�ؒ*�p����
\}��)Vi�=J/!�� nP���&ٵ"x�=�U�S=@!�DԷ0�,���������
X�	�!��F�0A�,��Bz��d��!�d�K�(���U=i@���ѣNm!�� 8ف���*w̅sd����d[p"O蘉�%���c�G0����"O��#Q"-2�����&r��{�"OR]k$	�c.��j4�* ����"O|h2�ڶf/\������"OhQ�vM�-��d[GeB�BuR��u"O�	�D	4l� �4��v��e"O���v�V�Ψc�  �y0�1�"O�P�D�#�.]�TN�7X隌!�"O�}�H�cv���M��"��"O�uȂ�p�� ȓ�
*��0ã"O���3�	�A�����'4��A�"O�-�`�)X��ݫ+��|J4"O�`�	�U��`ŲDYPY(%"O
Q��nU��*D�˯rV���A"O^Q�1
XM>���h�����C"OH!! �ոW�v�ccfO,Ơ�"O佊�/\u��c�nP�	�6�ѓ"OV ��Jёm�����S?J�f}[r"Oh��lV0u\R�@�̧@��*�"OF����
bR � ���!���9`"Ox�sa�-!�� 	רhf�u�"Of �Ǐ�3���s�˟wSR�Y"O(�X��-&b�sU X�^H��B�"O��p#�.�}�T �VHz��a"O D���0C�B���Ȗ&.)!"O����_�X<�3k�NF"��C"O�za�~����D$Ú@SP��s"O<��C�u���A�$EO���"O�&���������T+��*`"O(@�䟃wnrxB���!EXu"O�����٢uӜ�8����;�@*�"Oz�ҁ�"Yk���IH�VD�z%"OXtj���Y#�<�gE9Y���d"Ob�j¤ȒG4�<;��\9bH ��q"OL4s���+ǲ��FM�	0AP�s�"O��2��� :�0�̆�+*���"O`К��4�4I`���:�XTC�"OTA���K 9���:�C�"�U@�"O@u�U�D�r��Ⱥ���b���d"O�u�A*C��÷�õ{�zur�"O Ӧ�=f ��4꒝>���ZR"O�͐!��,����+*!�쓤"O61eD>��q"���T^���"Ob�!@�Jݶd�v���sb��1�S�	F�w��Yp!f�]݌$8t`N�G�!�ē�!�h:U�ƌ4ev,���[��D<�S�Oz���T	G6.5��l�Yf���'ҼEz��/�Vq���L �^�p��'��4"0^�)�vQ�+�,5��B�'뾭)VF-�V��	�: ��x��'1a"�:s�f�@ϊ�>���b�/�?Y�'��<��,ω;�T�#�%�\Z�K�'t��ٌp�H�Ib�  W�5q
�'����ʇg��""L�F���`
�'gl���y�J���L�(o4��"�'y0�8�ʛDz%���	aP���'IT�q$b�:�p��ۘR�H���'��] �ǉ��B�#�CM9�I��'W�P�Nŵm��!扅�:����'�
iƋ6Tp,��O�6X��2�'�.��B�Z?����u%Ͽ� ؃�'	 ��w$�/
C�ö���-���
�'�
���nt�fEi��S���R
��� ���5���/&���,�TY�"O8U��FBhr�@7��`P"O����a֋
fF}��⃁8�6�ie"O |���
]�M8�!������c"O�H*���\���9�Oܳ��:�"O�P�`d��~!f��7Oܴ1�4XT"O:�h�g���
����cИ}F"OHp���Rn�"����X�Դ�"OB�@&��	{@Ѱ)S-@�0��"O>Bu�fH �5��5\��x�"O��'cº	P��>��pb�"O��#���2P����-*"�)�3"O|a˓��=K���
R�2���"O����5M�d�:�.?t���"O:a{Unȸ2�f��b��:6���"OF�4�;��<�%�6k�����"O~��� _���&�>٬0�"O�X
�m�.�&��GM� �6��A"O�� �*�X6�QIë�)]���"Ou���)'�&H�7�p�"Ox��C���|BT�ȟk���T"OV���E]V�D�a�KjDm""O*���L�#�&�Š�+\9��"O>��f#>�X\�e���<�&��2"OTH���h�v�)��P<��ٺ'"O�u0AcΓ {�=IP�������"O&����iHbQ��oژ�3A"O�x@n�:p�ܙ�oD11�䀐�"Oi��L�q�b� ��"f�n���"O̬�s�	��1�roZ�-�� J2"Ou���M�1�n���ъ�* j�"O.m+%��<!�\����"�`dHe"O��爇9<�y��@%7T��"O��Y��42��扱�DE��"O�q�v�C�]j�[s�I--��<r�"ONJ��#%b�q�J��Z��4��"O�}[�V
tk8H���Hv8\��"O��.� t�~+SJ�l�q0"O̘ʵFږ~�4�RR���\i
Tr@"Od�yV睘;���@��"O�X��mD����81����"Ox���r��F�=�F��Q"O�Db�c�#1p���d�7K��A�"O�hzD�XHAl��$�,%MD� !"Oh(���@�%ތ�c�]��t"Of��F�M�Ls��W�V��4K�"O<|�4��:��M��	A�hQ �C����4b��i�bKǪ\"�'���'B�]ǟ��P$\,�Qn37l�9 ��0�1xVDˈ�4Q3�D��7m�Xi���!M�0YJ>1%K�дy&j�2�T�âl˞sR�X*w���j�t j��G�(�P<�O%�r6�� t^
��'����N�46���o�Q��O�i�Q�'O�7]����	G}�/B:���2IL�i�vi��,7�4ʓ�?���?���'��|�uF5P��uЅ(ߡ;)�Ы2*Ѧ	�ߴ�䓦�'��]�H��\�5j�}�>��f�ɁMĠqçAC����O���O��q3j�Ol�D�O�m���Ӆ�����gմ#�����Q�th�E�+]
�M���ܕ>ʙ;�X*n�Q��SUN�5MZD�2aOd�88�A��:$>0��D�t�Xp�oϹ.����3�Nm8�"<q���lH��F�rL��b@E~{��,v`hL��>����?��Z?�y�JL�'6j�3�i2O� ,tg(ʓӰ<Y�%��A�4H�3퓉) ��3sL��5Z�*a�xEn�ٟ��4(dp��'n������O(j����υ�bE�`.O� ����'�2�'�Ɣ�7|�$��G��<��Ec����� ��K%ZlTH�5�N��K�͞ �(O+#��i�� RO5(ЍZ7�ϬHg����+����F��'
���p��ͣ�0�<�Q	��|�޴nFq��E A�^0F�b���pg0����O���dX"9��Z$a�(2\���ꟙqL�Y�'b�"?a�iz�7�rӢk&А<�̑YT�Ҫ*���p$
:�M#�N-=����'@��'J���V�L�r�'��� ���J�&*\~�3�C�59ƬR�,�������#IR�x@a���FA��l��3��O��Է��!#@�?Y�J8�Ü�ApHZ6�iF����mV_6� : �M�~�F ���L�B1	Փ�\c���$�W�/NZt ��QC�-�ݴV�)��3�M��i�B�s�r`�EM�N�0�G�$afD,���O����O�=%?�¨�=�f�7�AX��M��k3ʓC��F�u���O��:E�j������&Q4 m*,�B�jsF��?a�[�T8��.
��?��?1��M���Ԧ	����B]�Qk�[.���9�)�<t�h�0�N5�l T>T�B�?� �T�_���O\*�!ڤ �^�3!��SWt*�Υ"p���kF�:3������d@�u�a��a�D��.edȀ@�۔Kb(��A�$X˄��I�5������M��i�~�'��T�h��#m-����A�8�q�#}��'�q٬)a��&�7/��I���M��i��'����O��I�h��&"�U#T%
�%� H����� A�����T�	ݟ��Q"���	͟��)uj�fċ)�zB�H���8 �	̏i"�ܘ�.ʡ���1S���T��<����["D��)�%���qg��.\5� ��JY��ȣP��N�(8��O�]�JD����[	�?�ԠL?
�jc��mjx�A%g؁h�.��x��'.��T>!:����f6���Œ�]$$�wb<D�trC풕7��z��Έ(��⥌��(��4^�&�|"�'7B�x" L$9 \  ��XZ���A�Zy��'����`ƒ��V������~���:#j���k��S�JD����n���E}a�������مl]?�B�F{��Oev�I�#�?�F�)AJWvɐ0B���)�
 � ��%(�l !:wV���EC�䓺hOq�4%iWOαm�M�7���bm�%Z� D{`>�I03Z���W�@�c��
�䕉E8��JH?�y��t�O�@�c̙�Et���'�N�����y�'�����X�iKyx5A�
j����v
�5Q��OL�=���T:���TEҡ�'��l�і|��)�3={�l�)X�V��K1�$����hOQ>��I�XΚ�h���(l�R(�"�O�B�	%/ξ��E0TQ��B��eAN�>��̋�a\VKQ-L!VQ�O�IPAm��4�×刎h�s"O|D�!�F?3��mh��J+|舺6"OZ����eKlp��֋�U*"O��2�$_�>���#�Ѕ"r�R"O.� _%��0�ъǬ7��3"O�`j��Bl��$���+�6�@�"On����aLP��J�^�~X`�"O����R��@�X.t�f=:�"O(��4A�Hc��gS��ֽ��"O�l9�j����NdH�"Ot�A�i�Y�V x�4I:`Bg"O@h�kH�K���	�)%+!�9�"O���kש<}r�z6� 
k\�Õ"O� hqÀ�H�Ա����!��4�"O��)���<fH-P䈚�3�8Di�"OD���Q$y�)@�g�+>�`�X�"O��k�i�6�d��P�P8�"OƸB�O_��I�A�҉
G�\�"O���O�4�&�b�=U=h���"O�` �d�>��8�B�(9.�S�"Ot���(1p�)�3*N8y����"OJIYVR!K�lz��ē
 `��"O��a���+k�M
cM�5�̀��"O��ArI �{eH\s���3L��У�"O��UA�5<>*��l��e��80"O2P��=O�؀���	CX�"OT���k.<�p��8j?�p)S"O����'�6�,���-?F�/�y��/,(-`VE�%��e�p�2�y�H�P$����N�����y�ǋ:\���J�h��s���y�.B�R����wj�&�~��"@7�y�C�&a]b�f����|<�E��;�y�+êI{��sEHT�|Đ�D`Ɏ�y�؊t�$="%O�
)���m��yb��H*����ɬ2�0��u.E�y�IΙx�$���vCX�:TM��yR&�23��I��Kj�B�d�"�y��\�U���%�ft&����Ϻ�y��=B-�ybb@�[$�!!=�y�d�y�P�j���~�� �yR�L�4
h����w�8�a�!�6�y2�³u-x�KgDV7o�&�ƬH��y���,҈Y��"o��Պ)�5�y���k�|AUa�;`��XA�/�yrjYZB�� ��hv�E���y�EQ�Y��{fl���홧k��yRĊ�8W���V��
���F�y�G��z^�� ˒
	s A�����y�Hb�b9����*�(�PdY7�yRh+����G��"$(���Ķ�yZ�e�4�!���j����eY��y����%8��˽s[����?�y����HL����i��y�3̉�y�C!ʂ�(�U
g_ܕȲ�O��y��5/��',�b��(�N��y��N?Z@p`���݄R��i9����y�GJ� �<h���HTH�m7�y��@�D�&\�`X>Z�g����y��dV�4ʂ�"r �VC��y2.S*H$����1/*���!���y���c�) C�.���S��yR�Ҧ�Z��'ϝ 2EB[��yB�+Z��ȒK�	�&������y2@�3'��@�/��|�zQ["+W2�yRcS
{���RE�@�:E"R��yrǛ�t�]R�jDj�"�c`芤�y�3:� �!`��do�xIP�:�y��ڱ�Q��i��
�������ybei�<}J��<Y�Pi��9�yB��@�o˾K!x�H��M��y�!��>q�S� pX���"�ξ�y�	3q���B̘6or.|�b���y�#L�����)�5j��5�CN!�yB@�� ^��9wGʔX�tUPQϚ�y��N�5MWL��쉨�y2�׶H��I*�f�#yyAQ�9�y
� 0-��MѝIJ�k�k�D",�a"OV�r�H˃�Ð���`P��"O�b툀S��jQJ̸�>��!"OB��$T�9 �	�IB�T �r"Opɀ�c�?v��Ao���bȑ"OZ�vcO�S!����[3}YB���"O����.O�P����sAH�yP�y�t"O��XtoL�iX�K&؉TC��"O����xW�KFLsKl�`	��t��� �:��2�X�3CPd��T��0���WzZ��1��y:���C��y���?Ĩ��Y
 ^^��ȓ7���ˣ)��~�k�hߍ�d��%k�yS�!X�:#,��P��	>�.t�ȓ;^���#
�)���^�4Q�ȓ<n
H*��Y��
�I�� l��ȓ6H��Aƚ�����e�c�r�ȓ<EJ��C��.i{��g���4�t��ȓ@6�Ѵ���^aR��Q�kBNх�KF��F�S�vBZ�(3�OCtX��ȓ��A�&�O%b@I`S,H	3w���u4��-���#&M�w��ȓ!�-�%,-?B uW��MA�'� ��(�K|yg��v����'�N� J>T�'��"m�څ��'j*l��/+�����,�]����'���(�!�/
��q�#c��{�'�DQ#�R9C�J�yd["{��1�'vH�c��ۛ	Ʋ	�##��
�N���'�u��������#M�|*pi�'6xQ�vؾ�~ūB� ��I�'� @��7�L�����&Z����'�V�����%�ǩ�.���B�'2@QB�CO�}H:��FC��\e��'���&�G���@�Gh�hI��'� �r�K@��4 '�Y.$����'jfX�#a@��f��6‎'QX9�	�'Wh�a7�Áx��p�f�
�nB�c	�'\��z\'P��	h�$�3��U#
�'��P�Y��I�&��Fʈ�
	�'��j���I�TQ�	ʊ1��T��'�HU'�����K51��xP�'.h �CF-��j���$r�p���'�"�
� :-�D�B)Z�Z�0�K�'` �M9v�|,1R��A�^q��'�fi#rk�9&���⪙�@��	�	�':.�R��S##(~y8���=�(l�	듛�Ɇn���`	B�����69;�C䉊�L]��L.�혤'�~RC�ɶ�� 0�(P��	KD�L�
�&C�ɰ.�f��a�Hr6���E+8TB䉤0��8s��N�%���)�*'KC�	�}��k���:�V0pCϧs��B䉯U����b*V:����,�rB�ɈL�J1���9{;nEx ��:;FB䉠/�(x�cgY�9���ꓥ6"�B䉷 �F��䀜�MzP�)B~�B��7wN�UI�!�pT2�;,�.C�I9n# �	сUbr!��'�8T�@C��y�NQH�mB������ZtC�I��� �2C��FΈQzDmY;�!�䊙kR�P0���'mfI����G�!��޵V*�H�L&1jbui!��)J!�D�&c�<� GK0D2�\)�ß�Y!�� �ؔ�}�T��#M֨��"O�d��CgNL��6�y��ك�"O�M+S�K�,BjY���K�.�C"O25���^�L�\�p���P��E"OD<r�	#�b	��=ø�1"O��RVjM�7��}C.���L��"O������0=}Zl�f�A�pP�p"O��[Q�HCg�H���#r"O�xKå�` �`�ĸ2�2Py�"O��9��Ot��U������"O� ��O�a1T`[�X� ��"O>칲��`��Ӏc>&�9p"Oֈ�C_�T�	�c(�.�z9�"O�����;�E�'��"�l���"O^�j��T4���ဇO�<EPv"O�p�"�Z���1"��L
�f�_�!���ot9��g�,��	aO��v�!���(qC��c�PH��A�Q�!�d4J�FQ(`�	�;xy��
�	�!�䊐b���������Wf�(�!�ޞ�$��BG�b;������?�!�D^�0�0���=:,��yԁC�L�!�U�RX̋���:��P5GZ��!���hHȈ��L�虊V�Ԛj�!�d�-�vx[�j�&����Ui!�D�.�Ҙ{���>�-RF��
�!�Z]�0��4$ *�>�U��2�!�$�X��p�� #�d��+ϴY�!���uT5ڥ)9b���R
�*X�!�ЂV��IE�V�"�Fx��+Di?!�GyN(��(x{��J��c�!�N8
l�X�,
?Fm�=�!�A�Z�!��	�r�k&N�vR�dYc��"�!�K�D��uKG�B&$8�Uj���8�!��"��#dn��B$�2� M!�!�$�I�<p��*5��l3�@[g"!�D���hbH�j�J���f!�d�;?�Q��,Ѹ7�E�#��%@�!�d���#��̤\(�A�Hڟ'!�D͓_�l�S�\��ic�gD!!�D�
V��2�����Yq���5!�ΧP)-h椘��,h ��)W]!�d�G��� M"V¸ݱ�jL�~t!�ƳAl} l�WC"ik��S�d!�$�#ݎ�(��"$�<�0'^�YS!��3(C�p��iM7jny3��X�!���D�����F0	����i�=�!�D��96Hpc��V:,�B CBR�!�d�KY.�[�iB$ �bD�d �TZ!��PjX�+�z��EQE`֤7G!��M�?0��z%������	W�� l:!�BKPs�	߳g�@, �	�F!��2<^�9���&0 ޔ!����^�!�ox����=����O�=q!�$I$¾Mp�͙�?��s6��7i!�$ȫi�X�6`׍Q���֊˪2!�d;7 @  ��     -  /#  !.  �8  �C  �O  X  �c  �i  4p  �y  ɀ  �  R�  ��  ؙ  '�  n�  ��  �  6�  y�  ��  ��  @�  ��  ��  	�  L�  ��  ��  >�  � �
 I � � -& �/ %6 g< �B �H kP �V �\ (e �g  `� u�	����Zv�B�'ln\�0Hz+��D��g�2TP��ƕ#Ĵ!�5�?YV̒'�?��]O+0���֖i��X4�^_cZE�Wh�~T���.6�4y��P5H��x��	Ѷi�J���-D���.K4n�$�!�.b�Q�NϝnY����끁x��A����5���;/������k���H�
�r��P
C�8b,��􋋲G�	��K�d�d��ӵ0@ՀS!N�2@\l��:)���P�	ş���<O��8针ͱ���*�m�;Wn�
CA'Qv&y{ٴFg��'G���O�T {��O���'l��Z�+n�$A�N<�c��'���'�r�'
��'�ٺ�N�=�k� A�h��Ա�z,8y��B�`��=˄��\}B�>�Ԅ�]�'����F4!t��Σ0��{D�!A0���<1N>��'��T�@�\o��Q�'c��q�ELr@.t�Q>p\$����<����x�����	՟d�OU�.�,<��ː
�X����?r��{�1oZ �M��ik��z�"���𦥈��ϑ=��(-u�FU��������O1 dV,�'���L�x�BA%|�(�.?�tp�׻<ł���9 j�sZ�"���G�eW`��)�Y8�8��!�8qڼ���O��m���M�����D�Ou��L6D��V,L �bˁ!}�j6͒�4�ꄡ��IC �=(����e2"�߷`����i6�LͦI*���`s|�XV%	�)$�a��r���nFeΈ�ڴ{m�f�|Ӯ�6#˲zDHM�@�Ce ����+�1�Ŕ�f��4V��v��e��+��TPF�Ӧ9۴���I<lF(�I��I��`�U���AS%�[EfF�3�fXk����M�g+Ǡ�4�r�o�,�B &�?�bNT( Y�t�$l_(<"�$ ��19�����Or���OZXmZ����^Ɣ�	Q��A|��hT���N���ܟ���Jȟ���������7w` �!�*�����4�bU���7 �~��0A� R�2��D�i#�#�	�:����f�q˴���=��l�bPs��) � �@� �!�M#k�W�'��}	,O<D�'[
X�$�M�]�xx��U8\������?9����?�����Oj��M��?���BfG
8�V�'��OP�d�����{Ԥ5��쟤�oz>���Ge��S�ƧBt�I�DW*(.���|y���|��6��O��?�̻?�jaJ��O&L��1у�=)O���I�� Rf��¦��D�
tq��i��������Y$o��hϾ�;g�>?I!�7�R���hJ5 �i���	�/w؜�WI���aH%�	
C��I%)��D�ӦaJ��)>�[��2a���<:۔}��<���O����O#~:qILNl4���e]#rlz�'�7�����|�gH4��d!f�A��a3���M����?�Ky��*Ӈ���?a���?1���y�d��Uq�O(JL�y���@����O*y K>LO∃�ӜYt4#P錾�� )�!q�A8f���՘��+&`c>c�\�����ܻT	Q!?�T	o��9*OH��'��t�?�O����c	8�:�ʺ<z��Y���O��=E��$�Et>XGM�P��«ƨ}�ɺ�M{!�i�ɧ���O+�	�!&����h%h������p�~�	���$�O���<I+�^�Ӏ98�0�H:�L��U�Y�f^�h^�2�P<B1h��n<Fi��	7��hY�Lܚh�p�ɝ{ N���ӏ�5��o�W�VXT&I�ls�#>����iOR ��A��J��DH���6k���	.�Mcs�]�[e�q3� å+0� 3�Ri��)��?)��0>!�"�3 ��sw���_q
�@*�}�I�M��ix�ɘ+�)�4�?���E����o^�'N�$3�gM�L��|����?Y��1�?���?�׋�1F����%��q�.�xo��z=(�hpa�,?E�"�.@VmZ���-��5`a�!Vn�0�l�<*�䡑�
	)4�VhLi4� �)P-�L5� ��+W���M>����ܓݴf���'C�x r+ےh^$!��]#����\��l��?J>��Qܧ`�ꈘWi��kN��*�E�d0����ܟ�'n�7�Y���䇈�>S�L1��G���m�(�4�N sP�U���(O��	Bצa� m;M:�+��<��4�@H�<2Q����k�4��lʂ�mWD���ի�q��WJ!@.����Ev�(C�C]����!��Xe(C�
U6�� �E�B�� ��ɎV�2t� �,<�ln	X����!"j]7as&��'J����G��&5�i,�ӳ+8���S?l��9�B��5z�O���-��O��d�<�Mܢ,உc�;,?0P�2n�ؑ�H����M��Q��'e�tx�熷S��,��`��,�f�6-�OB�D�O�LC)�5<b����O��D�O���I<�%A
l�k����0*^�f�6m~�=mZ�]xJÈS��%�	�0h�+�G�L4�ԏ�>!#��ѩH,0��'�N*A�|hsr�<�S�z���+�f�Y��r~&1(�L��4w^Arڴ��)d*���>��O����O`�����)���P5�T2Y&�ܲw>�2�Sܧp��Ӕ5T8zdʃ(���'[(7�@��$�$���?�'�*��[�,�=�톬)����[�[��7��O��$�O����	e>="�m\�;�x�K��T�a���"r@�	t�r�9Q�[&F�ԑR�vx��Pr
 dV�wI45\eO�&j��QaC��H�:�Rq�Y?��% %�;)l8��f ,Nl� С������Bʟ`�ܴe{��HGx�	�g���vF	0g.~�� -�?�I>9���?�����0ߚ�BDQ��B��2	Nhi��$R�%����M�ײiy�>)@���4�?q�'�X]S#ƍ�d�B�l�I,uyh3������O���|>�8@�U�xThX��3��)o�Z�? :��a�:��e s�O��lQ��'�aqF̎�;��q����Z~D���d"05R���֣'�P�Şq,\!����*3�r�w�J�'��8�
˓�`� �B�%v��<�O>��D&�	7�t�[�&Σ D�1C��~{���DBҦ	X@MX���UX�L�i�h���N<�Mc-Ord�r�B����	ş��O�b���'%i�Q#K1�ܭ�v�E���9��'U��Vn��plœP��قp�ǫ-��5� ��S�	�*��0*��:+�A�bņ�<���A����N Y�q(��iq��n�N�rट�d:ܦ���V��%	���G������O�(o��H���St�ɺf�9{����K��D�B�	;w�
��ꖧ]�h���
C�n�?����Y7"�{"d�,�
6�Q�x�lğh����p��|�t �Iܟ���˟��;%0�Q�L�?1��I� �Z�*T�S��s$����e��;z��&��Ņa�'<��fO�MQ:%c!=�d��E�T����c�0h��c���Ov�hX!�EN?yC�D�^L��O+:�T�dJ�˟��'s�IG{RNFN`HX4k	��6�����pP!����@�Rd¯@��|�!�G�4�.�HO���O��q��ੑ��#;�NYpf�׸���AD���ؠ	����?9��?�������O�ӕh��`Ʉ*:J��7B18�ԼJ�ð7!Hԩ3'�&IW�J�l�p�'�LY����N�SG�q�1{d��"����+GA�8P$�3wJџh��g
J��� ���7���;t$Ζ1_&��O��$.�	Q�O�#���1]�t	� ޕET@���'(�
��ǟ9��Z�k�AC�� O>�2�i��[�Ȳ���8��������ћ%����c���p�K������)#p��Iԟ8���Z��qGL�ɛL,��G&BH6�4��%VB��І�I�a���M��ؠ㗂6���g+ �BU{�_3<��PAP�K���!G:�9G���I�M�#R��wf��X�(x��V����dh.�D>�	ǟ���ܟ�͓G��D�K�G�= ���U�a�	Ix�D��47���*U�<SܹÄ`dH�i:b�d�N�bT�Ħ�	hy�V>�I(VS��P@Q
������O�+�m�����-���u���&?�~h"��i9�Yy�K�6)R�J�4�h��"?I���Z�c�([�����:? ��|��(�K� �i!��(jQ��"ခE~�"ޓ�?ir�i��"}z�Oh�Y05��.&3:@{�悝T9B[O>9���?���7�k3N��&�H G2�"Qː�#N��?q�i�^7M�O�n��|�B#�#�ɲeK)A�`�A>�M{���?���3�FPa�C��?���?���y�����ipTd��D_�)Sѯ�[׈`�l�n �L��߷�H�Ȏ�����!����v�<T:���y�~�y��"�H�Z$�&ީ�DO�MQ�h2IMţ?�X����\ђ��"i���b+S���Cn_զ�I,O�0��'����?�OX���B!��V#ӝO���)5D�\R���7�V$�@;0��y�B"�<�f�i>m��ly2�W�u&��P$_�m��̻o�
LF�`�f"��IR�'�b�'���h���hu�f��&i�r���AЂf\nfc��Z�FT�\DhuXWFu�V�n��r�<aj[�2�UtaΪHza#�I�D�Lb�b��xs���C�-{:�80��ͤ"AJ�<!��!1YDu`�K/{[@��Ҩe�,%�ɐ�M�V�i��Z�@��~��!�~�P��K7Jz B�*?Y����"���O�I� �h&&L|���;Ə�����-�M��u�����i��S�$�`��[w���'pF��0�GM^�H�m�=����e�'S
�B���'��)�;��� ��51�D�D�445M��Ɉh2:�3kL�?��Ȉ�*\?I�^����iV:��­@��x��Хs� e�Pl�l���c�쑱��a�w��=<������ə[���3�D�4�$��%*N�A��-i���-�!�D�F���Hwk9���r�fը6����O�Q�7$����	undq��|��V_rf��?�/�d�91h�O����(_1�t��D�V���r"�O*�J|)�uIc��Ȝ�S��3fE`����[:8��`ɤ�u,ܥ_x�uF��$�4��'CTxc"hĀ.B���ꕜ(�La��� �0����P�Ƈ�<c�l�����C�,��Č6*��'Y7��O�"|*S��a�P�#T�Q �;S��D��ǟ�'��Gx2�E�o�ҹR�*ưu/���Cǆ�?�����5�4�?qv�i�8;�`�a+�	����Ƙc�7�O����OR�� I˨B{��D�O��$�O�ݿ8`dӲ��{q��z�̀��<e�B�K,KzT!T '6��x��*>�|��F����(ϡt�mTH��O2(�aՉ��V�R�۔�p���'a/�R�	0R9.a5�:A 
1Þ��+?!�@ԟ������?�4�\8
*Z��eA0HL��K����yr�ߖQ�D`Ԩ�$FU��Z�%W��d�\�����'�	�����G�Tv�	A�V)J`Z��$,�.L��ߟ��IΟ��^w_"�'���[�
ض�ိ̳s��hB�S%o�]�C����6W��ۅ�5��:|��� �r�*�HA U�"� � 8g�p=��� W�Q0�2�� ��X�k�*e��PBω5�|b�'[̟ �ڴo�' �'��O�]����"_R*� �"�%9hm9�( D��c�hߢ:��e�7��4�$!���;�$���M��dy�*�'+��7-�O����� ��!����&�>!�R	� 3�H��O ��B��OD��x>=���;��������TU�I�1m,@�� �9R���Ǡ�3	Yl����<0��A{�H�7<�TɈ1UxLsv�\�3涜ig�V%D��h�`��4^T���uF�O��&���!�V`��]�Eۻq�f`!�!.D�\�U!K�>l�\�pF"pU$�A,�O>����R�
p@%�A�F� � K3��O����O��D�OB�'yQ�� �Q�)) K	��3��ߘ��9����?`$#a,d�n�q �@�FE��I �!�	E��eh���wx������y~��E�@��HX$�A�����2;k�2���LSܵ��P��)��eޓ7� D{F�T�ART��'l.p�����=��;�ӠL������	�Rk:�1eӐHQҒO4��O��d�<�����)X�?�ؕx����!x�Z�
7џ��ߴG���� �4�p���:tŒ���״<���'���'�KRFD)�y��'���'�nS%S<��@��p� PgoܠR��'�������}X�\��M)kk"ă���.L�(�0k�(��!��!�';ZD ��፵�
c>���(>��牥%P�(6�N�h+8��򅓭��Hn�0��$�/���O��3���O8�� cK�ukh�ר�F4p���O���?���ԓ���UW$�J� Zw�%���<�Ļi�7��O�lZh�4�OH��	N��4:D��vx��ɢ~�v�҆Jʉ�Z��I�`���L2[w���'��I�1��1 di>J9v�sCOI��2�@�Ze��a����#'�^|��1�x�!��]h�޵ХԼ4'�`��ƶX�~}h�%z��M{!6���"�H[&( ь��M�j�,,����ٓ��P�3HR(a�"�o�*(Gzb�I�G��!r��'"���+"k��B�8A7�8��ʫ-Fv�`TD����O� o�����'�ҹѣ%�~j��eԄp����9~y���B�V8����?A�@��?������ͤWܤ:s��5p���jE�Ϯ8K!L?� ��΀,7B�}��*ǫ.�jIFy�O��!���d��.`�"�l����D��O��'���wHO�,?�l��� ��QEyr��?yU�izʓ+��<j񉟼YO�x�U�:D�v`&�4��&��}ED
���.ZT�Z��DJ���yk�?i]��t`�F��-�TN�Ob�Q��H���?	����鞙	��d��'����4�_�/�y�ل1%&��O؅��Q�D���޽��oZ�?E�3C^s��0J�(�@�p�"$��̑����^���I�̛�~I�On����R:?��'g�B�/O?�\l+!oâ'�(m�'-f�����?I��	k�\Zb�0�ܸ1��Xe���+��*D������!�U�T�8"&*�	�>E{7�x�T͒�m�A�b��p W�U���4��T4 ��Cៈ���,�I꼻�$UEq~��bmK+J/Z��4�P�hm�qG �4�^[�"�L"�y�|"$xMN�ɜ�U�F��6g\�7�8I�U`L�W�Qh0a�z'j��DeE�ӁM'�0�cq޵���I�����ޯt�f����O�\��Y��ݟ�E{�疽<���ȵ�Πd �m�&㚙~t!�D�P����a�,j�T`�tg�6�8�HO�i�OLʓ��)K�, ��FS<� 2􂌁zw�hR�ON!�?	��?)������?A�O'�{���/�)��R����!L\d� ��D��Y2�iQZQ�`m��(O�ĐV#H�O�4�ɍ7=�h��/����6GJ�\��90�f�b��A��E����?I���!�tP9&G%t� �eG��c�@��ٟ�F{r�ɀg���ת^�:��a��	��8�jC䉚a�m���1/��:�O�:��O~1m��0�'Bz��y�2���O�Y ��4d8`��L���xK�;���'�����'��:�B�Y�i�Z�@MHE͋ ��8�äݯ��ȲTX�o���z�g__�E��HG7�(O�Ȣ
ض�jJ��R
O���*���L�J��u���F
�l��	ÂC���(Oʨk��'J��O�PB�I!SV�q��Z^DmP�"O��c��� ��e"`���wU�5�S�'JV�$Ec�P��(ԏR��蛠���&��'"PRB�q�t�d�O��'� ���[�\�3G�%�䭐2O l)�Ջ���?���Ӥ���S5.��T24�i4�Sv�d�hK�$�Q�D9>�4��l��R��� ���D�՟y��"Rk�4_R� �)擷O9�q'�G�m�4UQ'� i,�;٨5�	��M[���D�IS>`d- �t�̍�F�^?��'��|��I [�����ϛ}5R�B��l ڢ?Ab�i�R6�%�DÁCH�R�LP��< �)���$�O&���O�tx'FqP�$�ON�D�O��ݟO ���GI#Wj��V��*B/��}r-��Ƅ	��gܓ	� �;W���~�1{�F;��� I�'A�L�T�i=rd�aŚ���Ϙ�� ���2�B#q���K�@�a z���'��x��R˟�'s�<��l�gbZX6�٘-_fpRT�u�\�t/���T2�G�!)�X�ń�<Y�i,�7M+�4�����<�dO�?Qiv$(�M�&k
���F����b���?y��?��Y)��O���j>���iۢ-�qs���r e�2����51�.G���C���XjRI�'Q���'� 	��h��KՔe/�qC��U�eW6��Ǧ8��𕅖�$���)u�M>�p��?Q��T5�N�Qb�2.��A$��<�b������F{"�	�R�j��#n�� � ��<#hB�	�o!���F�-0
�s4c��}~Z�O�l�ʟ�'y�h�F�~"�a�>p٢��?�zU�0%N�qv�Y����?��.��?������g��}�n�S#J>K��3�i2��;#�h2��U�ӓ_�V(�u��3�$� ��D�
�!��fߛ{����GyӪU��M (�j���G1h]�!CR�+���A�F��w=U�	��'���%�#I|�8
$cɗ
j�	H>��ViZ�ҏg2ֱIVFU�k�e�����?�n֕6=�`2���JqIc&�<�'"� Y&�q�2���OZ�'{�4K��#S,�7b�FԪ����S�QM�4���?�)�p��Eh��O"+��j��S�N�vjw���I��.�;�Cݫy�s2�*1F�ɫa���6D&Fh����?B�v<
&i_V &E�OgL����c�H|x�bXB<���O�����'^6]�O�)�1�8��\/2#ƀB�Ǔ^
!�^�Mn�б(ց.�e#��,�џD"�����~���ደ�	�G=t=86��O���O����B�-����O����Od�OO$u���ơ�@��` !\����^�%�����oJ*�$$�Ӽ:o��S�O� �ӁV��m� ^�W�@��#���A���+5p�=3�
DF?1�j�2�-��~2O�7z�"A92/΂4?nE����Q��Ƨ�<�A+Bܟ��~�L>��9R�X�SЯB�y��8 �DE�ya�px�� �N^�p���څ��dGE���$�'-�6iy �'b?v<{�k���p����O==��t������	��$qXw���'���N�	-Ԥ�R��xM m�"��
K-N�Äd ���Ͱ��ݍ>��EH�|<�������(!U�Z�tw���C
�"M�P�� ��u�d%z%`P,�J�{���28�� ��$B���I�(S 0���p�o_�XЦ�ؤ�'�"���".먁�P�r�<���F��!��2F ��ʔ<%0����7P��'�07M?��C'c�a�O�R���>���ѳ=ԊU8�o�4*"�'�)�S�'��7�>	Y�g+�F��hɩ^! �Faϔ�s7L'O������Z�L��k!�(O̠K�k�;_�zy���U!9>f�l�`"���@ Ǥ3�8-0�N��8X{%�� 8jQ�����O(`l�����ؖs|@���t1�Ci�
���M>��C��!8`�S�.�0���#G�Jr������?��&E�>�8	 I�}\hD#�GVߟ��'`B�x�����O�ʧ6W,���|�֔1��H*m��)#L�86�j��?A�ϝ�2dԩpEB"g�H@ڴn���'�����X��V+��x8d���/��I='�0�ـρm�=�'�f�RQk^wL�h�O?�)'f�1d�*�:e(A�&��`j%?�U�џ\�ش3�OR�O0�	��t�D�YU
WN�,�Ad`d�'�B�'R�(���rߦm�WH;Af؊���O8�'�1�>"��(3�p��`c�?p�,��s�V���O�dU.g�z�Y���O*���Ov�$g�a���C�fzF0�(%e9��Ǌ�L�8�e�8V��JE��^_rb>'�+���} (`kѢ�^�Bb,��r� L��ȭ/Y�A��BQ:�\b>�$��,W>�03��B]��9K��&\�b��4k�b�Ob�d�O���(]�<�	���j8�82�ʁ�7�(B�3]X�e)�,2K��� ��,	�77�������'\
@h0aӣ$��Ȁ�h��Jꮉ3�$^���#b�'���']Is�)������'Q�����텈fGB��`�٧Tv���T��,�4Yu��7��=3F����OP�#�� YʔD���>)riP�Q7�A
cc@1k֩H���ޣ?�7)�TcZ�ZѧQ�o6��H��B�nM�I۟@��O�������n=N��[��[?L�Ft�5"Ob�+� ���(	wʂ�$͢�֓|�%}Ә�Ĥ<����-.���ܟ��08m�ֈ(��?Iv��J��՟����"������̧D�2$I!('zV\1�t��j`hR!l���"���0P:��	^"!���?��ʐ$����ĽC��p�t��0D����2%�hM��"��؜5���!��D�L{B�'��I��-@����
��a���fø�O �d0LO��̞%>�6e"G��#g����'����݋plN���nv@��ą�0OS���R�Z��Ms���?I,��8��f�O�`�������#)�H{�ԡ/�O��Ċ-� 뷅�j�\�����/�n$�OK�S�ysP�	���%jP�
j�#F�V�b0I�.�t����i
�sYڏ�4��%9>-Z��A0Ҵ�G�!����,F�B�'��>e�IS�? R[�A�#��b�FT�< ��"OV���)�5^���夜��̑����h�����b@���[�d��ɼ��nx�L��O��$A:>l��4��O���O2��|�)��ڌC/0բ��Fd@ #c+�`daq���N�n9ł����b>�$�8K�n�;],�� ��8�*͸&��&6�<��f�=p��)�\��b>&� ѣ��]ߪ����T�����kt���d,�3��6K�Š�!B/�B�L\wEhB�5��ؑN"��J�۸,�˓����b�L*rUᢡK8����\=b��DY$^'u�e�Iޟ��IПD�ZwUB�'��)�O:ށ*%�B��]������q��ٳaR���]��p=i�U�|/*����,.�H�4�7)u�9�dβ�uǭ��p=�6dN�,Qȹz#�:���$�4)Y����M�P�ia�OT�J�T��^<�B���b����5JA��H�?��hY�`�8\��%��f��)Y�@�I�M[�������|*�lZP�t�I�����W�F�!�����H��0<��b�f�'Sɘ�D�K�����"ʸ���CÓ�8�Gxb���5x�������L���<�0<ـ�ǟh�<A��6Mq�,�C���૆�V�<��(�3���@��p���R������}eF5�� ��*��Ъ&O�.g��$��1Fd�� #��+?�-�N��ɤsż�2�#��y?��E�7{R���O"��Dܑ^q��慉�E��P�)�'f �	�`�/V�D9�N��yǮ��'drp��z��}jҊ�&�>9r �
� �B��voC9^A�  ?Y���Ο���L�O��Y���
�� 3SJ�v��!���=s�.�kB���$뺄�g���Pџ�@���<*D^�h�L
�6����g�܈h��0y��	�I��9�	�?E�	����'D�����Si���I��Z6{T2P�9j�%�Ō�O
�2"��>�1�1O�ͅ�U[�	����>5m�X!�-�U��(V��O.P�@@R�1�1O4)�p�M�<̼aP�_�u���V�'���>c)����Oh�=��� &b�N�[�Ҝc�>혷����y��('8P��+��eCb�!g���QQ�����<��ń4H��\ �"
)\�D��4�Q_BL+A��y��14P�@�q���^S�����'�R5�����+�bQ;6�r]Ig �_	މ�&�հ�?A���?q���?9ч\� Ʋ�&G�me	�w��+'Cص㲫Ϫ[5�u8&$L":kT8YpfȪ�$Gy"�O,oZ�@E"ȳ ��"@�16���Ʌ�|B�@��><WV��w+M�y�GybO8�?	���O�����]�9T`YZrL^�r|��X/O�����9�6�B�KK�OLڂ��%��}r"�<A�U+@B
�0F�N��ś6�Ky2�8�'��Y>��� ����I3a]*�q@ޤg�
�����.Fzz��I�3h�ŭ��	��xkg�
��Mc��s���������Ky~���ެz��Z����y�
�E�0M��H�3g*`5��i��d)T��O�
m��\^���ɳnǹJ�n�@�'��5����?9�O�O��I�).j��' /U��TqtA\X�~B� [�6Z����Io��&��f�=a����o9J�Jcd�#(�J�h�莀Z�np�	����I�h5\���Cß�����4���?u��*:�6`A1a#3��1ۦ�[�m-�<� N���MKg�ܭh��A�׫A���'�hQ�O�L�n	%��)�ш��u�l�{�ˑ^�J�o�/U�eȢ�Z�O���?i��n��\Pf���HHC 9ä�����5����O��=A�'Rl���%`F����_	m=@�`�'x����(�=��=k���3k#T�"��6t���ޟԕ'��j&�Y�"�@�O,,>��V�>pn����͵[A"�'��	o�%�Iԟ�ͧ//Ի bҙ\�p�ԉ-�80r`�~9�T�FI]Te�	��M�o���d!ʓb9����O�c�����j����J�Μ�mJ#^X<���ʓ�$PS+!�2��I=})^8*�#\,W;`�y��Cl��	y�'����B��B�q,�Q���ڥI0D��I����;�d�[
=��	���<i��iQrZ��*wEP�����O|�D�8�q��{7 e$��1�@��U�(�X��O����80����JXke����Բt�C$[&��-���.���ª�.U�����	(�F��
U>�E��X�e�N|j��׭w�2C7"�� 1�Š�'��x�+i��l�z��I��P�|�ҩ�$����uD6���Q���Qy��'aR5�E#S�&�1��D�j�x�2
�t�I	Nht�T��]��+2�E>0h<���� 릹�I����O����4�'�B%�i���ddɎ]H腚���"�w/HT�dBR�PK�$)b�S�4�$C�jI1�b�	� -s�d���Z!�Z58O�l�D���9B`�@���n�p���6sɶM���V����d�맋�,:2Q!�8�I8�b���O�S��z~
� �鐖�w��#�H?&O����"OJ�7�"w��I�WK�/NR}!b�I�ȟ=:#�Q( ���5i؈-�p<�W��O<���O>)��j������Ot���On<���?�F�-/�VQ�d٦j���L��4 �QJ�s����Jܣ^���˟8�zǫ����I2U����X���Ę�� ER"-��o�`)����!=������=5���'8,z�*e1}R��5�I��gѤE�>�*rH���D�I���'Kўd�:�0'�Ō
��ȣҁZ�Q�pͅ�2��ۦfW7��2���x�@��	�HO��O�˓ ��l�w��4����*I�l��i��
Ȥ��E9��?����?�w��l���O.�ӿ�8�
�KD�4�e�L�*����<�r�@�ߺc��P��_ $$�`�I�<��a1	R,��ic�h˓b(�������<��l�,�|� u��i��LB��u�*Ah��ɰo���/K�]c�a�ʙ>EZ��	f�'��2s$�T�6yӅ��#��(D�8�`,^o��K�ƛ�U�pƥ<�q�i��Y�X��l���`����̧'Gĝ3��־{�d#����,d�Ʉ�t��	����	�& �9 �ۥA�̘"���3/^$̧x5ʱ�ˈĒ�� F�M� D|��L4qK��(�V@3&����3Oj +g�ЅC\�՘p+^�nz�6�� �J���c�Q�`��0�I4�M�����1wf��+�< �j��"-���'��O��$�O��İ<�3n^$_[pX2��YU�Ɣ�C�����>9��i��7-V6C��0�wBY ;�����:C�˓�?����?Q-O�˧�?Y�'i��꣭�)i�j���'z�a�OJ��П�'z��S�'B)�<aP(ĳ)&��Є�Еp���?�ڴ�ē*IN�H<�A�ֽ������D2��L˦��	0tTb�ΓQ����������1�=�Í&k����!��M�Eб

��M��:������yR`F������sbן材O�|�m�q�LX Q�-{^�4�'�rȄ�:��d`ݱ�������h�#5��!�>v�(��qɄ?W��#�����ɹ�p�I�<�uAAnz�EG8Ob5���L>T�
����<�x���O��[��'_���>���?�������Tf���f�`Ed���D׺s�L�q��'i�����?�ȕ'�?��'@v�q��M{�oN�=h��ȃ�ڐ��	�[mv80G�i�0�әS�"�'����K�O&�Ο��	�?��@�Ǥ2��E�����r�S ?�]ΓH��L���qXw�R9O|x@@.쟺6��A�&i�d�Y�`BgL��Iy��O��ɍ tN���O$y��?����\Ӥ�C�S9��rĘ�k�z�(���M�V��ym�ћV`k�.�)�OLE���q��t�S8#��L�rC@)A��+�!B0�08m�X@(0�4c�����ڴ��\��i��z C�iX�\�H������;��ȓy�X9� h�z�^}���)U�*hoZ韰�I���	Ɵ����D����T�i��h­�5�, �-Q��3�yӒ���O����O�˓�?Y��?A�w�$�VoM0j$l�4�B�$v^ v�i�2�|r�'�|�ٟt��0ސW����M��!j��g�iB�']2�'����I(}2þj�������	t'���B�C�����O|��hO��	"AN=���P1�U`�뉇`gfO$���O@���O���<�O��,!q��:3���&D��*��"�O����O���?�*�P�O�
�bp+��8�x��O
�)4L��'�H
�GJ`9f1�k�&t����'b�,���-c��`p� !�\��'�ha8E(�pT2�O�DmN��'|�@��E� �S�%_�<�L���'.M��$!tL�a��d�	ߜ����D�O�d�O���O�us'.щ<Qcq [+��`
����`���������I�����ן�:1%�.4�m֢ĢW�E�wd��Mc���?!��?���?����?����?i¥��=�!`��\?�Bir�G�2��F�'���'f��'B�'��'{�#f��i�K�70�.��R��UH�6m�O|���O@�d�O��$�OD�d�Ol�$��{�Z��ǣQ<���D�ʮn�韀�I柼�	������	��$�	/Rm��7m��H`�Ś0��Y��4�?��?���?)��?Y���?��!�P��ÓY ҵ�A�ϧJlv��iVb�':�'Z��'�r�'���'LB����Y����wH�q@�ls�K|ӂ�d�O ���O����Oh���O|��Ov ���}��kv$�)����%������8�������Ɵ$������ɟp`Ï��D9�l�%�;n��ك�޳�M���?A��?���?	���?)���?y��0_�t�/��d��Qg�6��V�'D��'5r�'��'��'r��O��A����>:X�FK0|��6��O���O���OD�d�O
���O��Ը[��5�� �XQXA� �s���m�J~R�'y�	s�O�03t�ˣup�E9w�[$-�Xe b�i�!k�yb�)����͓ &�86�E�Pθ���M�U9V���MC�'P�)�	�.=$��A�O1�I+�,07gt�p�'�4��O�Yw�\!A�i>�͓h*���e�e��7��"�O����f��v+���'�� vp04B�3"����ӊ1ep�����Fy2�'���4O2�Y �YF�@a��s���(�L�'V�-00��)l��O���=@1Oz�Dr�+�Lt��
�4-3�7,�<i(O�&�g?٥�߸4pa�fa�4s\x��bT���44���'�078�i>s���4aܐ� ��ݨV���$���<���M���rVh���dSV~ҪU�/�6Q@4G	�C�@V?� $�1�J'IZR�kV�X�'c�Q�p�|�6�U"/NȲ��ԣ+�&͓\ʓHϛ��
�Ș'��Y:ņ��h̨c�ī:��=	�L_my"�'���<On#}�gb� ��h!(�1b{n�Ke�4�eHV��a~"˂�7L�tr�j�{t捪j5E��X�QI���0xG����0p�4�,h����b�τ+Šr��o�B�UBߓ[lҹ����)f$h��g_�_XX�<��'��ZTD�Uf\�MVĠ� @2DjڙKa�F�Uq��sd���Ei���S+D$D~MxD�Mx�T_7�j$!�bz�@���:"�`�E@�,p�p%6,�m)�A�P��h�� �|8�Y1�U<*�]c�.Nc�xD�܌(F��2AF֬}�"�!	
�!b�u�d�D�Ln�=ΰaA��8	0بr��g��S)On��P:O����Ox�d�^�d�O6ԠC�hrCnW�NKdŢr(�>\qO`���<q���d�OZ7�C!����A��t� 	 t'�?>�&�<�'j>���qy2�O���;`]�� m����CC-�T8����'�R�'��%8��'Qr_>�i>qm�����4�D(��C1�<t|�(O���<E�T Ѥ#4����7A<�*� 5Z�y�Q\R�R��׆����=y��&��������RbB<��٦@~��(g��Ub����E�H�,��$f��xrF0;�D_6�jN��TV�h����IZ�`�1�@�\�|+�c��ЈT四,"�h���	�b���BA���؋l6L��mO/�TpH�朕0��( ������b�&��%M����0!fV�4-6�;޴�?����?IcA	�ĉ����'�F������I�� 2h�G���:q�O<4�D��l>���OX��Ѧp1vU�0A^?�@d,�O��
:H%��ןh�IH~�(�\Q����(�Y"���+OR��G��O��Od�z-읲�%F�/Z���[�S|�3 %*Y�'�r�'>�|b�'��sQm��h�I��w�����C� ���'�B�'!��'�r�'�7-�l���ٚN�*�r���Z��RsP� ��Ꟁ'�$���Dɶl���@�W��5'+� C��	�x�ZveC��|���H�������������ħnDXE�%#�ȩ�g �A�LX��?1����?!@#�Ģi�(�B gY�^l2��� �Ai�����?�����A�9���%>	�	�?����^. �x��GJ.����b�TH�	ߟ��ɭC�#<��XF�%`�78� ��E;!�T��	qyR�&�6͢|�����&T��3&�"�Rz�)��H�
��<A�'N�+����m�\ ���I*kJ�ڑmC)F�$�d�;��l�h��ş\���ē�?���KOH z3̘�����Eݝ�?����?�?Q��?ُ�d�'��k[�0�V<�B�
%
ڄ2�-��9Ѱ7��O��$�O����'�v�i>��IΟ��@���ix��m�B�r�۰n�I�����<���?���䆌SeE�lF��0g��1G�؝Y��?)�
���D�'�X��ā�g 5r�(O��]A���l�I,AC"9��^y�O�bZ�����4��I�$MK1����ݞ���X ��Ty��'j��d�O���ֵ[�50��_&�$��Ȱr2I(��1�I럘�'�!t��O
Z��v�ށ�zP�P@�P�z�̓�?����'!2�'���Z�8O����Ȝ�T%��s�CՆ$�8-{EW���	ʟp�I]y�̧ �R��i���[%(�����m(D1!�2O����Oʓ�?���Y�����	�1m�n��a)���"�SUh�'��Y�ز���'�?Q�w�
 ��d(��������5��*����$�O��$ӛarl�$#��`ޥ�w�:�0���]ZݾE��H�O��פI# �i��ԟ�����D��O�mu�"a}���e���;�b�'&���v�X>����?]�O9a���x@Х�2f(#�����'e0���i}Ӟ�D�Ov�$���'���dI���'̂�9�����(ZȽ��z����ş��˟���P�\?1�iI��Պb��!F�z�G�����a)$�������t�l��)�>���r	۝�?9���?13� ��A��mR
{�2�+�.�/�?������?���?������y�B����B�G@<l�������ӟ��I~y�#�k}�'��S�LR���PI�!aZ}j'�'���'��I
�y�'4R�'n�S0y�����E�m���7%\�l5�%���I՟ �	s�IП��	6L�^T�g�в^E��� �Sy�Q�I����IX�ȟ�Iӟl���<I��+-���ƯG�n�+B�G�	ןP�	ß4�Iz��|��	�Zv�h�iY:� !٦)����?����?�����?� �M�y#qހbx���@�Aq����Q�/=��&�)����Q>{����l���?AQ��W�N�^��)�L��=B�m�u��kj�$�4웹�l�:��)BcX��g�I�Bז�[QNŮ)j��B� ��G2h��G%	`�p֩�;/7����:_R�P��}�2m� �{�8}30�@+:�0��б;DԠ���;� �:�ש%)B8�4lN�&`h9������ß����N����⟼�'	��l:��9��f��Y���԰Q��E���R� ��m��I�Ge�9#��3@�He3��C=�Zt��ŉQu�E���T�!2�˞y��8a���gT���!TXX$MR:(��*R2d:JuA�E�������d�S�D�N�5��ЮQ78�fǌ��y��̝)?NIB��v|s�'#����$K/F`mZ�p�	I��&�:>�Y�S�ɣnQӗ$E@iZ=�0#�O����Or�`g��A�]a��Ey*��=��șU0D��g�vR����$.��X��nwF�>�S��M�]S����**)*����'ғ=������%?�l����� x��as��[b )�������G;٘YJ��}���p썅�p>	��>1TK# �aQ������C?��$؀e՛V�'�BX>�`�Cǟ��I����V�
 +�v�wd�,/ȝ�G��gp��1
K�V/Y�AW�<�O���?�<+2�;Q�_3z���$� ������,R�ej��n�V��)B?�쒍�\cv����d�&b2�j�+P�p��`شS���ɜ�MSR��I4���!��=@�(�� &�m�]x�忟x�	I��P�R!��xŎ�k���0�h�z��GyR�z�\�mZy�J�ԅ_*D�@s�Ƚ-�YZI�o]
�d�OTp�P:'�����O��d�O�]���?�ݴS�:M�6K��*I"S+դ_�,��̛�W��8*�-�?"ڞ�b�-�p���I�-������ �m*
��T�w=�C�n-^��"����t����-F!���;ʓQ��BA*��xn0(s$�"0�0a�'^j�{�iޛ�ks��㟠��O9���)��~A�m�o�57����'��i֡ݲ0t��Z��2���!�FY�'�v듘��P���mY�H@�ä@�Y1>pY2ϋ"����O����O�� A�O���d>A ѩӄ;qr՛����\�U���o�Vu��-��Զx���צ�kkP1�b�<���;@j��A�[&�� QF�̕o�H����$�b9`�o���M��	B=�t�����mɿ:vPu���ؗC��p�&#��q�c�u��d�<������iȅwZ��F^xb&�끯B*`�!�ğ�d� ��<8W^Pqv�\�Q���E3�����<���^�͞����DOWi�B�h!�z0��a��:��'/qO&�?����̮a��9�@R I�i��7����b���:9�$�P�'�`����?�-�3b]Q�����6:�B�	,�jUHP.ƾ.%�y��L9i:B��(��]#ď�:N�����h�K�"O���͑����&�Y%����"O�
�F�����bn�Xv1a�"O����܊4�NF�Vn�B���"O���uf́?��c� :|�~�P"O,8�"��8K�p��Y��v���"O��)W ]�1� AZ���0�TUI"O� �S"� -$�ʄ2u��F"O�P@��ԋjx(ԃ$ ܡdͪY:�"O:Q��͗9Z:Z��f@�D�0�T"O�E�Ek=@Oh�(�e�2y8U9t"O��+Qe=gF�����%iz�˦"O�l�Fn��rL&ڐ�A)X-�b"O� ��d�.��Ɂ�O�NȈ �"O\�dS�&��� �=35��+S"O�	#F7d����S-�Q�\���"Ot��"nzKj�Cl�=��Sv"O���̈́$Z�����p�@��"O=#Ć�"D��Q�|
�h�"O��J5c�(&�WK�X����"O,�x��V�N�v��Q��?D�<���"Oq`# I��a+�)#qFܼ�"O�\�4�oWd��RmM'pG@��a"Ol9#ւ��s� 9`rK�'eҴE(�"Ox�Ѐ˻y}$)B���7H�U��"O�Y8j�=5hPI�5藲K_�m�"Oܡ��F�r%8+Gq���"O�|�����X�N�(F��1z��YA�'�椰Ǜ�E3���0k��1a<(A@n��+E�i!�'���q&A1)Ҁ
G�Q4h��Y����ʔBa�4����i� �>1�Վ\���EH�g�=��9��$+D�� 4�7��!�&H�A�ʹ��x;�cS1|��:�����1L�O?�I�3�E�WK�+\J�p�
!��B��/��������V��ť4V���P)٘XJ�E����YY�M{5`�Q������1W������,h$%�s�.lOR����%Gz��!SiA0���I��>钝0&*6�4]�1hJ�e]��D�P"��9����m����+[qO4��Ȁ.��B��Γ.꜐-����iQ�.ԆR�d�/0�.|��ȣ(]!��F�j�6$�o�M���	���7k�f`�vK 
�ј��2"x���&�S�n�^��46p�x�Cc�t��-3��I�.C㉚3�z$1V��q�9S�e���	��`14���۰C�4�c&�O�2�|4�	�Cצ�k�֎*Y�9���;Ӏ���V+]�	����=ޞ�Y�m�b�X��C�R�!�0�L��.Q����6́���Hr�o�&z�rݚЭ�Bf�&���[*���C�"R�O����X���a��}��N�5>��i# #C�zo� U��H�<Q�BϠ�j�[�.��Na$IH�B�f,�,"`�G>@�ࠔf�.��I�b/�i+���;2�V*��U��xq���</����U�Dq���X�9��<��&D�	�<vŔ7y]�a��L1ydThc0@��dPBa��%���(O:$j�ć���`��#�^��a�'Zqɑ��+C+�zACU�B�4i���� �"��o5�y���j� ��P�ѭy�|�b� i��1 �Ź+�ꅛ5�߫��Dρ0-�Qi�\-:�L� �BO2v�(Xc��W��ٺï"�!�$=��̈���9`dp��nɳ��x2��e�Ma#�^.Ij�K5N��i��M ��1���관;Q��(�v��d��Ay힮H l�Su�3�y�'C�N"Jh0"`�M���5N5�>�+\�k��t�	|���&AW���=�S,��o�����oj�"�韀:��1���P ��5�!V( ����L�<�0a�!*��u�˟@I����DR�'�H(�p�R#/��;%DCA�4�Flő<a�"V)�5��.�n�,���ާ*i��Y�2���ɶm�=%�q���	�c"�H �o�F`�Cʌ`}�p1�b��4��V�f6��HF�ϕe.�|h�K Op�sf��b{�lV�� VH(�Cp
d�vy�ggI�R)�J����?	���)6G&`XЂ��6M�Ǜ	sg*�:�'.�I�@s�� �fë2M0PH�$m�dgȼ��䇖#�Y�΋����H� 8'�ā/(V�Rc
�`�d C�-Q�4X���g4H< �+Fr?����I$�1��_4����
r ����1�~"�B�vb����e��p����'�]jw�H5��pԭ��m��9�/�'q�|xP���p�J��Ꭻ	��	Xp��0s��Z�i�2��ҠJ] �h(����t��LKu�I�)� � �}Y��+a�V▴��@�dF���X�!m�-�`���;\��c�BзR댠 U���~ʦ=��,P�ԁP�k��T]��ȗL:�O�YA�]�DV��c7�W�#�.�b�E]���%"���wj�c"-�� ]�%�ܣ@]��{��ּ$�8�"�w��T��Yyʚm�r�܄v�P�s�'��]@�'<��hs3䖾yHL	�fM$�\Z�[�u�p��!Fa�d����&"y�=p7��}BX9Ԇ���@b��ۂv���Q!���f��C�V�;EZ
y��O�LkqoX	�Z���ME����'*��􆩘Q��[y(�3E�Ĉ-��Q�.K�|n��'�?QF��2�r�h���0Y| ">у�_�{��j�eC4�<q���<����g�`Q.h!�#O�%Z����j߾x��B��C�0�$1rE+;���K�e�l��M���^�K ���6E�!W�0�f	�D����Fξ��hs�+�"b�`H�V�L -l���A��q�^Z6*G�j���b&����Psw�E!f�vl�&M���
6�åx��qT ƊcJh1u�(�OR� �K�L^-�@��/U!FC%5N�0@�)tz@[��Qg:`:#��#A �6�i/T$�b,F�Im��AD�@R��dх������j�6;��B�4(�T�����vQyr�5�a8F��c^ �� ��%ot��èP�� -�䈚�/�[�fW�?��z*�M����� �$mQ��S �S�����F��^��@�啼�6q�(ؽk�0����tYP�+�S���ŋV��zm�v��T� äϖN�88���\q2Z�J��C��fY��#�O��+�ёJ���@�+C�A��DX���<S5锉͏F�8�3��u��EaQH���p��C��T@�0�PlHf#�#B��@��3X�V��'��j5���d�[���bKp�9��̮rj"u� ]8$J�2�$Gb���2�W?Yb'U�$=� �'&7�ܴFGv	�Ӏ�H�H��Z'y��G|¨H�`��6�P�<��������rq��&+��z�Ή!����(W!p1x�h��p<ѳ/�OD��S��a�XI S|}��"D6"�=�|�o�>\k� �n��\mp�q2jH�FBb�h�/*4��J��I�vi|��AľR�RI�B�:D�dC�'<`��c0��53:�Qi�6D��	�� Y9<�8A��-|ȌT�C8D���BHX�`�(Q*��.	�| �#�6D�����Ap��\?�r(�GT�y��H�V��Lyu�Y�bay4�̨�yBaԋ	��HX$!!T��I�)J��y�f�+)��,�:=.�`SLI��y
� ���	Q�����ц	0u ys�"OpUȕl��K�J�pc�[!d�����"O"��u 	7Q�B)!��R��)�Q"O� ��W� �*A�RE�PԾY3�"O� ���eܨq0:�4��"O��ٳ+�6q�i����oE`�J�"OQƋP"������Q�S>���'"OI��\;5R��UM�	3��<�3"OHdC�ɗ*	,��ߞ�d1"O�@WG�4�$#SC[�s����"O� q��,47�m�!�ԞO�@t2�"ON�u��F_x��çGtȈh7"O2z��E�BG��u`Ga	l|�"Ol����!G6�1�v΂���YS"OQ�BC��Z^d!R�>n�R �"OB�1��q@J��$��7+�΅��"OV��a�ͣ>�x�d�Є6'zd�"Oѱ��S��`�I����y�"ON�r"$_13�X�ʕ�t^�[ "O���r�ÚQ��TBF���W�-[W"O���UΗ	^�� �F�,��Q"O��C���8G>���`�*ub���&"O�ة'��P/�I�N�%Xf���"O�%T+Ki�F
�L�A^,*T"O�qJ�H)v8��!�ګhO���F"OH5��U/	8Π�P*��t)rg"O��9r�ӟ)y��5�!l}1�"O`4��ΐ�$��-�Ӊ�� ��%"Ov����6 2(��W�(�P"O�$�T���p%���Zx�^�˄"O�(��+�Y��1xV�"Y� �8C"O`e2�aS'9�֌�ӌN�ܜ0""O����%;
��p� �:�VHq"O�:`�ߴ�@����\*^��k�"O 1�č�87B�B�G��x��"O4���֭K��k�����b"O ����|��$M�
9�$S"OF|+��B+y�rB$-Վ(���R"O�Yz MJ�F���yt�Y�OU:lJW"O�d�'hX�Wr�&ꍼt�n�s�"O��yT �4cdι�PO�'��"O��Qw/ƇC{�̺�a�?_��`@"O�(0��T��S��%}��z"O�̹��E@@z�v�Y��� w"O.���c��1�V�K)�p��Ӳ"O��	!���9ꐫܾMa���"O� 	�A�/!j��G)++_�=��"O�M���8�ęz�hY�hC�Ds�"O(9�e�8�8X�g�[�@pȃ"OD5��̜* �d+�o\�=����C"O�y���:��(Y'��>�@
F"O���GX
=y(a°#
J��h�"O�5E.B�z"(%�ta�"O�KukS�ͪ����;Q����"O�u�� T// Z�3��6T[�"O�t#���,0:��L~(
=�W"O��r�� ;�q��E��0���"O���L*|�Q�ǯ4&�H34"Oԭc`(M�)"5��N��w&�3"O��rRGѰID��rb6��z7"O$5Z��\?g�Љ� Y�K	�a�b"O:,I�`���)R���Ie"OF ��S�y���.�',�
YJ�"Oh�I$*W�dI+���^�\��"O� �E�DlR�L%`c/UÎ�	c"O��X�9%3�]v�R �0%�"O,�!H��gz)�&k�3Z9.y7"O���n*F���@�N���"O� ����8�Dt!��h%Z���'秊��iI�!�Dx	@�C=�fT�	�'��5;��M��|IE �P
E��'�)��D�o�PTꔄ��`�pL��'Ͼ����Z+H�Ź�"8da2�{�'��])2�U�k6���f��kD��'fHz��ͯY�*P6(�ʑ	�'��Ł�K�$�$s�
�H�X��'�F�J�]+t���窊�@�t�'�0�!�k�gC��5�#D�pC�'�N4�5��6zF^�p�0���'SrW:�Pq�B�Ɔ��Ӗ�6D��BD�j�@A�6 Mֹ�:D�����P�0F(��΅�P���r'A6D������*�:�@�H�4�pC��6D�<���ƣ	��!c-�7�`t��k5D��$��X(�˦���^ɺa��g3D��gՈ=H:�'�L�����4D��wh� s��p���)ێ�j�*O���JQz�^䒀d$�lD��"O���ׁ�+5��]�����Š1"OR@8��b{��
�B83�(��"OlmXWF�E8�P�
�.�� ��"ON;��P:
�Ԁ� ޙm`�}��"O���Uǘ�n�Z�a���
̰"O���2��d���4�HTx�"O�����^�:!�N��Y�ʥ�"O�娳�̝U��h�0̝%z��iB�"O����!�<����@|�U�g"O��v͂�EovmKE�U	�uQ"O�1z�A��%��\)#ό4/��W�� `��!�H5��tKbLv���d��J�$��GN�-r��%�!�d�g��P�&L��E�l`��/� �!�D�E�^�dÒ�n��N�� !�ƠZj���ϛ�T`�Y:�N�=!�Ĕ�_ ��B����M�PD�<xc!�dD e�ls!L��*�Ơi��7�!�$�9L{�#F!�9~����BN�G�!���W_�Tj�F�#c��#�%4!�$["&|C'�Ͳ%�NP(��ݽy,!�$�8i-\HX�I�~�
��#�`!��䂡�%N�|g\m!3�K /!�Ć�
"Qq�O�#K`�;�!>.!��ҠO-�&#�@1�j�]-!��	e�d��� w�x����'!��M ���^�av\�	�^�@!��C����p�U&js���3EE$S�!�\co�ڷH�\@Pa�\�6�!�DY�|�̬��͆6NF��J (E!�d�b!���OC�=��m�3��\!�Y�i
�_�4�9ć��^B䉴N�`�"�*�b�!�`-Y*C�	�)���CߪC�$�2��A�(C�Na��j���p}���B��
t�B䉘l���б(��d������ЙBQ>C�	35���3Wϝn�r�z�$�&8�C䉴c�(<��ϛ�mR��2ÏR| C䉪�a;�.���r7(��\@�C�	hP�C��"C5�� 4-V�y��C�I3h�"8��+���,׃S�C�)� �@�p��9hK]!�B�3����"Oʡ��H�E<j����˯���"O`K���'EyL����!��[r"O���B�/*�,X"A��cX욳"O�sC�7lǸ�k�@�J���B�"O!�&�A��|:�喩n��܉�"O�-��b�!M�����JMަY�3�x"h˥\Z�z�G�<��$�Ԏ[�&͚��qjI��p?YT).�py�Y�] �s �>76bDP��4D����hH�8�l0b�S+9B� P�1�J���>�'}�^���"�4`"&H�����ȓH���֧��"�:��^v�là,�)�'&'t\�
��d��R�@�-Ҥ��]ל%����bt���iϏD�h8@��'Bk��NXv�KR��#t�$��	���(O�QTBT�=L屇�"^J����'��!2���'J�y*CF�����4ņ/f�J���/S�����..���a��ԡ:����	�a�V�QD`J qخ�E��/T6�'b�\	&�X���m!4��*UJ�M
ش�?�����$�Ę
��[��2\��d3U���y"i�7#l�Ѓ�� b��yY����8�r7�V/}��#�{ʟ�x[�����y�LG�+{��P'I��#e���fK�Px���5Z�Q`*�oH��p��+wu���O<���7��5yA��Jl@��$��#Rn�DD>#�a�e����'�Ӏ��'�z��eӟ\BI2�$X, �Ќ*Qm��x�b�Z�O�>Ĉ� 4݈RU����I�Ch���WC�>�	�+U�+��'�|�Y
G�:�V-�w 89}�	�=��(�%2�۰��D���C�	�r�Dx��Ww"����M��� �(�GԁgZzs#."�)��E��C6 �]�I9�����~�r}Y"���v\B�Ʉ\�ƨ���IX��`g�-U?�tz�>����#*~���$�8t9K';`��ܣ�M�)S�EХ_+#�t��I&,MI�:<-��Х/��mw>%�!M��hR�7���%�S1��а%�u�a|jӱQ"�{H]�o��u��C���8_Z4�d�/Bm8�(Z6qO�T��i���k��\�W�0�ce#�yҏV�Q��t���ϊPY��B�7X}hd�]�x�����{ʟPX��J��yG�^||(yp�6�x�nU��PxB'�):7~��F�,�Y��id�u�'3XH`��2P��v��[�b�
'd6�j>& �q+8Ԟ����&r����ɍH��Q�'����k t�����E�@�F��'�tC�'���D@�7(�NxuN�� �Z�O�:��j~�+ !)_�ӦB,J��W�!��h�q�� v��"�D�@U� �ȓw�ر�,����p�B�_�`'��t�R���`y��A2�&���/7�a#ЄָB8+7e=wG6��d�Q���˧��	��)B�#��ybX����<�<�T��T���O?Q����(�Bi�UB��D�Ji0���?a�A-2Jc?Ũv�Ӕ�b�a"�߻B�
EYA$�<�����?o
P)ӓ9�|(H壛�w� ���U� ~��'�޼ `nTJ}2��/E)|u��|����yb�8o�I"4'�=,s"�+Ge�<�y�눙fR�-�À ���Cї�?i"M�2kQ0��^
���q̼��)(��4����K�?;-�ei��
���%�9�O���CQ�>�x4�$�Ë	%��ɀn�l����b�]&4[@
a�ix5�;O�&���y� ]���M>�=z���?��Ot�G`GG�4���&/~T�(HǍ��P���]�H�q��bpdܺ�����@�A���PgP��D�fkj�ڠ�ȰM��)��(2剾cC6�O�Hh��ɺ!6��w?�'Jdi�f@!&^p�Qsm�U�85�'5��`C_b��f/�/T�R��N�� �q(�O?��'���O\����>r��U�H� 4S���zJ�]z�拍"R�"�E�tN�G݁\| zr�|TR�*�9h��$����

Rd9�Ԑq������g�1Ot�sN@�>�$��E�E�9$f�)$��A�����'�Va搚U��,���u�N/d���*��8ӊH"����I�1?*�ДF�k����ul�4H�9Ӭ.,�:�
b�!?q �Iتt��4G�`"��yZ�?	f6O��B$H_5'|���ₘim.U��2D�\ҳ�O>e-V�0�(��f�*���e�O��Q�j(sr��	��&\з���I��?��w��婕�P�^%��ړ8���'��P	�_���åM�1�̌k�\�fH�9J"�A��018�b����&sK2�R��>Č�)"O�,˔BAx�1b�X,H�D�� \d����[�m�g�Z6��@K��U����AF�6>&�ԇ�I,��и��7'h4UG�.|X�'�N�j���x��!��0Z��x��{Zw+�9P3�I�@Y��Ab "+��m
�'�� �Wɖ�%�A.�2e�S�0>�m��II�\dqO�S %J�#�0��F�E�c�LԹEl
�_rP�q
OJ!0 �3��Bi�� ����∿��E� ����1?��k�Z�(�>iq�ױz ��s�N�3ص[�&CN8����z��]�\���8�N�H���X!�rV�A�����d��>��[	ۓ�h�NL���)��?Rr�'�0xW&�Y}�l�%�O��倳�O��' ��5F�0���8 ��'bt
#�y��b������c��^?q!�6�㞢}� i��~�!W�X;�*�#Ha�<G�5l�X3���!��d���\�I�g�H��7"a(��ˈlZ��(�D��B䉼 <���ĝ��@aB-�E�B�	
/!�!w.�v�z,�T/q!�B�I3y�b<"ҢB��J��2i88B�ɳ$�Ђ6 �	z�ɶ	�:IB�I�H�B鉴mU�� x#�j/D<B�I�L᪑����G�ɋ@%��7gpC�I��J�ڱ�P�Rϸ��vn�6r|$B�"��D�bǗ�N��#/^�[��C�0 �Ԭ R)��*Q�C��]7��B��Y�d�!�y��ec&��?.�B䉓6]��VL���5�@��:Q7xB�I�s	�0s	ˬ	���GB��HB�	6*"���6�� c��"� Z4SDB䉮kV\|ɔ΅2@5�=pB�[��C��6IU���t����\�a��-%�C�ɇs:h��K�b<A�"�(bm�C�I�gHx���"F��@��"(�C䉥>/n(2C>[h$�P�B2.2B�I�W���y��t��t"�m��O�C�+l��!Ғ �y�T��I޻(�!��%)c<��X%W|Ȕ�fĨm�!���)}$i��/��@tA�˓	�!�D_�8�b�Ȗj�$T"\�(�)�!��,n�������ސ؂�F�T!��͆_h\�4�N�D��|��$[1|�!�$ٱ4?n�RD��>�>�����m�!��f�t,D���C�[�!��$?a�2�#E7P`��**�!��8I��4��CI����8�ȯI`!�D������aN§|�}�5G��X�!��(6�.�چ'וn�	�3ŎY�!�d��ny��aY�y�~���#̑H!�d��	O� �'P$��T��"\?=�!�J�S#$�922�ćv�h�ȓG����2Ɖ5��&M�O�V��ȓy4��ad^�X�j�92��=.�y�ȓ~�r���O�d
���r#ń�XClq٤��&֤�iA*��HR�%�ȓ�=:���r@�x֏�i�'W
h�E�m���2vC<����'8
V��FE~Ix&���/_TT��'j��sB�$p����\�T��'��s#Ǖ<N��u�q��	},���'��+�O�W/����π'V8�+�'j|풴�)��u��+�t9��'�Lx���õ!�ҍ�k���x�'���@���r+X!�ϟ"nb�P�	�'h>� ���0h���D�_�e��	�'�"�9���X䭱d�D�p$6��	�'ٔqw �	�u3$�7�l�	��� LHcE��P�$�7��lP8��v"O����6>npA�)MNTq��"Oh� �%Q�Ld^��b�\�X��3�"O�!�aȐ�]t`$ȳNՍ/�r�"OP��+�7z��(�Rk����j�"O�0��1"ftҁ�P3q^�Mч"ȎHU$�H�P�2$�_�$\�0"O��1��$wX�"ą06J��"Oh����^ʽ���Q�y8�m��"O����k,ȍy�!4��r"O��{��$vax�)���Z��9�"O2E�DÂMf,]	�țp{*DC�"Od�����?�����5�:""O�԰p�ǂ8���HeLI Z�!�$�+@(��ÐHި�fN�z�!��%��m�'�R�dЊ�#�(�!�¼�z�`�ɝ'K�JYQG�q�!� q� ��Ђ-���٠���wP!�$�$i�����g�&.��� �ED�!�O2f`���w���v�
!d�!��R3`e�`s�Z�a �<���ת�!��n�������Q[��m�q�!�ă$4���B�WZ*�`���,v*��D�q�,X�$�V{<�:1�M6�y��T`�`@�G,[1m�d�J���y�K�4���+̐W�
��O1�y���3�X��g׽"4��� �K�yr�11�lm��FF����kU"��y���&PF�
n��`�A�N��yr����=H�%ԝz�tIq��yBN���(�r�_/vI.��
�7�y�-Կu�������>��l�J��y!�'m���� 	)�@���A�?�ybhР]S��À+�/'PHJ�%�7�y��ytZ��'CD=����	�3�y�aӢ ��T��dM	â9��+O��y��;�^��T�̐ ����y��!k�L�R'( E�fH0�H��y2F,c~&4�Tk:��<��'��y� F���񣶧�1+��(R�H9�yR�U�>@K�E/�Ƶ��R+�y��S' 4Bu����W�	2D+�*�y�ę��MKsFR�W���F�?�yҢ�B��R�_ Kޜ�����yb 	�V��)�����.R��yҬR�	���F�D���4I�%���yBC�^��t�U���[�A]�y�¾^E0�'����[a��y�nD�Q�����$(�䩏�y�mۋN4�=� ���������y�J��W�J�P��4�&�cs��7�y�@u:��)�$[��q#��� �yBIX K��p���T��	3���y�̐(�~ԈAD�y��8b� �"�yb ԉ#��%	W$o݈5�aH���y"募&�(�zB�S�m������J��y��SkVّ��?e�,�!�2�y�j*W��pr2l��dIY�V��y��?,cX,J�3'�*����y��> �b��V��3%x�=p�m��y��bx��'g���E�%�[�yROI-O8ȔCR� &�h��6-���ybk�@F<��G�.��
���y��|����2e߃0���z�a���y
� V쐑ŏ	s��@���)5.�:�"ON[����=�a�ş9�>�@"Op�0���P^గ��v��M��"O(�p��͗̊�QF�L�
m�zt"Ohi8�&��LH�}�СASv�`a"O����ʐ<s~јj͚SR���"O
	s���t���T�JzBVhR�"O(e#�L݅=���� �[#
�v"O<���i�2��m�����0"OT!6 1���cb��%8F�*�"O*Q#��S7~��)���!y :��R"O0 h��3n^����e���!�DWM�P	��H1Z9����Z!���V�h CG�6�"D�C�.5!���V9�e��ú%����ׂ�O/!�Q�}:�h����9��T1#�;M"!�D5G�~���Sx*�Q E��-r!�d�%v���k�R�,)�X�Ql�D!�DS_㴁���� i>pɒ���h2��l�O�=Y��J�|��Z��84&~-�"O@(�A�>d}^��N&G02\a�"OV��������#'M̱9�ȥ� "O�0��@4b�،��%J9	�0�!A"Of�4B�[�T	&�I7Ch"�P�"OJX��N�2��p�d��5���y�h��P�-��Z$�#r �!�y�+ .��[$�]0%<�1�lޛ�y"Hۇ1H0rJ7{Pd�ŀ'�y��_�-b��X� ָ@�P���y�	�;/����#9�(�X>�,�ȓ
����" �\�3�� H��(�IgN�.�
h���(5��ȓ$�} �jܪ�c��# �Bh�ȓPz��`�>/�|��	�#;z��ȓ
K\���Ο��@s�Ӹ,�h���wa
��֩��$�@D�7��:Z@U��Ҫ��Vc�)vT�fD�QCd�ȓN��C��j ��Ăݪ�,�ȓ,j���
�DT ���U�&'хȓm���#�NӫF�pU�3�\%�T��ȓv��t��2.ji�.�03����ܦX3"
|=��"Lșo�����T6]���
�TB�� ��n��	�d�u�d1@)�� �T�x���Q�B� Ġ��Y�,��d����p�ȓa�y��E��~ ���6,A��F�ȓNt�Y���/.�l�2��[2��ȓ"�6��U�zz�J3�X	ؐ��ȓ.��S"�]�c� #dDmT9�ȓUkXs7B��i@ԆT��zਈʔ�r-����b̃x��ȓ��uf!`��	�p�ݔA�>���,�Ơ��E�0+q��h���*m���� 5uk�f8 5���&8��l��u�J�y��"��Qr3��Jp�݇�ZX�`A�j"*�aS�_Z<H��4��mp�S�N�� J6lS+X5�t�ȓ50%����mL(Qec؟7�u��W�(��-@!�ѧ*ԝ�5��2lD,�7��H������GT��ȓUT��Pp�g+�0��-FR��ȓv��UA���<�x��̆[Pb��ȓL_��{a΅�|������Tja�Їȓ���� �'��D*D'�?B`�x��S�? ����#Ʉ�i�<d�nШ�"Ox��v�N�j�#�g��^���U"O�Z��Ab��]{%��3d����"OB}0 �ՑK*�L BX�i�zX�a"O�@�j��iT骀G��.��E*�"O4}a����Uua��G:����"OD�k�ȃj6�aR�@*��"O|�X&��-"��Yj�`�2|�@y�b"O��Y�(��|W>���#�.}��"Oޭ��5y稕�6����=��"O�� �W���/,�^s "O�H`C�>�B��s�	Gh�4"O�Kvb�0p��UJa��>�u��"O����@"���a��14WHq��"O2\+�:Ɗ��!d��nDj��"Oh\�G`M�$Hx@��M@ /J`�3"O��G\s��j�jL�4�0��2"O�-���R�Ful4P`��5�j�"O���K-"QX"��~L��3"O�hE��B4�D���˜Xft�7"O����&Ww�HkU�K+u)�y�q"O�(Rl����8qF�s�}ч"OV�wJI8g��e�c�%�E��"O^��&Q�g�0��$ ���zp"O���un8YB͉U�� r
���"O�H$dW<r0����ɯu�\��R"O"T��&͛mo.9�2䍓F����"OZ���Iы%�z�t�IRՊ�Q"O�`{�g�|�.8��aІlӢ���"O��"�.��)>�A��*ߺj���C"O��`���C��5ڡ�S�w���"Ol�{"`K A�����P)k���P""O�P[Qj;T�Q�_*|��"O�&;_�{W��qo���fF��yG��,HY�r$I�j7.٘E�߁�y�!_?��,1�J�z�5�t� �y2K��u��q�O��;۠i��	�y�����$mX�8^t�Ó.T?�y�C��]��0�abƙԬq�ٖ�yR�ܸs�L�@��4K5b�R�眒�y҉�8�ސ�����MPJ}z���:�y�i��<Þ���;B�Q�0���y�G� �Z��S��,�΅2�D���y2��`�z�E�ϛ�,����6�yBЭ5�<��Kثx)��[Eǆ�y�ɐ=P�.)�����r�x5JŪ
��y�nˠ/�X4G��lc�1�ӯ�y�(�9z�����G��\4�ݘ���yb˅�D�
嬟�V��9�#���yBcX3Y��H��'��H��lp�Ξ/�y"�	:��`�(�;���)3�ԇ�yB[� �⭱rj��	@�t3����y�)U5?�0��ʶN�NI(Hڇ�yr�ޯdMF-�v�@�9���(%���y��GB>��z"��<n��ä���yҤӴM\�(�'IR�2@����I2�y�KA��uI�/�R%�D�ɛ�y2�P8�	q��\I�3��7�y"�� �JT(0@IT�ݙC"�
�yr׼�l|���6՜8��i��y2iP�#�R���@�{ �Ya�9�y2 J(|m8�+��o}|�s(V
�y"�]yi��Z�K�5tL��<�PyC�vE���ڗ(D�@bK�N�<� �4��P���J�+&<�����"O~ j�-#>���!�C� �TD�v"O^=3�@��y����H.'��0��"Oޱ�d��uQ��2�(azu��"Ov�xF!^�cgP@+5,؍*Q�*�"O.�����
�L���![CvUs�"O��X4�Ӄ�N���Jۍ�ZQ�"O�$K��x��P�ek��1�"OR��`�>�ʠ�MO�6� "On8)�D�@�	"�4;�x�85"O^�0bJ�x�L {a�șJ���;�"Ox��B�67�����Oa��"O�-	�KF?-�dt(�&�8Z��H"O�|��痏����3�۫.C΍
�"O�q�_$�vU��c�o8nE��"O��[C��"50)<�ȫ�M�6!򄍋3%��䁚o2b�_h�!�"OH���D�^�B	�@����Հ�"Oj)u�<OhA{�b�s��Q�"O�ՠ��� c�t�f��_�,���"Oʐ��-��b��KV�Q�J}��"O��U��=N)�C J��u�\pd"Ont���HR���R��+���"O�`hFF��$�"emB�Ɛ��"O�)a	�!~�`F&�=z�x��"O��҃@U%tTف���s��T*q"OT{6	X.&���I�>OA��9"O���"n�4�n�(HX<���b"O4yb �#0Bt��S ˦44�`#�"Or�9�MJ����A�I����"Of��rGT-�1�tl۵h��,YV"O����F�s�����K� /�z���"O���$�V�g92(�w��(B�FY8"O2�W��/ǦYV�x��z2"O�S`Ȟ/��Q$Ȓ#ռ���"Ox�j�&T�h���rg��S�>q�0"Oހ(q&J">]�yҋޚ[�\E�f"O|ੲa�J|c�*�:#��l��"O����HЇ>�ꍺ�Z�U�1"O	R�]=C]Lf�K@;�"O�aI�"�|s�<s��
�j�$Xz"O�E:`��54((� �Y�h{�"O��� ;b4{DΫ3����t"O HU-�~ Hi'�Ȝ��AЅ"O��Z�n@4�$�y�I��بE"O����N�X�@5ɳ/+�9�r"O�xy
U;J�H(��C�lm���"Oސ��"�dC긚Ł�pa�XQ"O�`ѣPR���@�D�N"�"O�Kǉ�(]�L����X@A԰�"O�%X�I�]X���J�t&t���"OV}c�)�
mh���1)TI-��Qv"O��"�E��\r����Y &e9"O�1��Ŗy�
!a���N|��p"O� X�艔@�D�bQC].�e�&"O©�$�3)q��Q���*.h�0"O���#φ�yt0Q�J� L�i�"O��QኻD���G�f���$D�pC�"�rFH�PL-�H�i��%D��{�f�"l�P�4�J)�!���"D��ȡ)]��4D���ʐä%ф
?D��s��
 �t��d�
</��8V�"D�T;&\�%N�� M��~Π1)@.?D� �TjZ�|�E	��&�=Qq�1D�� ^�xT��Y6����m�`���V"O��XF�:�(\�6v:Dt"O�����#���q-E�\��c�"O�9ҍ�">�8��,;����"O���2��Q"e@�'^36��5"OXd�$�!�v�`@ԓP&0�R�"Oza��]�A��)1
^�"%&�I"Oh��2�N�$���o�Y��2"Ox��#t:0h��_v��h"OR�@7E��T�J ��D�W�T�"O�S�ʗ9=�`�	95�h4;�"O虁��Z���1��
�B"O���� ,&�"�E�{M\�e"O��;� ȄZT��jG����S"O�=�t��
�.�����_����"O����H�V��h�@Q1�5"O Z"���M$>uǝ��F�	�"O�X��R�-�"-QS��y;q"O��@��ϟE�����ъ@��Y"O�QbjL�}J�L[C��9;�"yq�"O`�#wMh���k𣟃h�29��"O��:S�F*�l(�T��V�v���"O�"�	�~�z K�.�r{"O�����!�Ƌ_�R�ly؃"O�-Q�H�&�3a�I���QR"Oȝ�`��O>x�Z��ʸ;�VhQ�"O�9������0����$���K"OhYQ'�ЙiX���$�~A�e�"O�1 �%��@�Bؿc+�ը4"O��pr%�),Zd�B���'�]Au"O����J��ؑ�ꇢf>�#C"O����<h���$'��2�"�	6"O.� ���'��x_,i;���g�<��F�@� �wƂ1^�rhc&�]|�'�ў�']7"�yr	Z����Q�=�|��ȓqㄍK�ˀ�s2|��'�H�@!������p�gI�p�b�h1eY!'�b��ȓZ��T'��h�)�V�F�h]����?�&l���v|Cþ2rn�a4 �w�'�ў�'�&L��!-�v(�3��+vlȅȓ,s$�Ò��%^�zI���ڗ�JP��+�"")��$�D٧��
$&0��vl���	K��$��i��q���ȓN��]	��&9���x1hQ�bh��˜�H'K^�D����M�㨱��d���"�=?�|��bY�:XR���_9�lZ�呆$Sl8E�t\9�ȓc���b7�ڪDr��Ss�T�}΄	���D�9���q%���QFʎ:ΐ�ȓJ�<��֧I�'���YBj	)�����	�H���R3�(��΂�5V�Q�ȓ]�q	f�6 U$�e&�_瞴�ȓaш�y7�F�`��%��=��ȓ5`E���!>� �)�,Χy��h�ȓ�9�CJZX1	d!A l�Fp��C��АA��~`� yV��i}X �ȓ6�P	��bԎ%�"��G .!|�H�ȓ~�1�p�3tE4�p���V1�)Kv�ޯ6����J�&%����h�"���|�BxCaƣ�pŅ�uBwc_�Te|e��j�E����ȓ[�|�K b�������&�ጄ��8躵R��Zl�FX#�d_0*�R݅ȓJ)",0���E鄥�R/�y�f0��S�? ��a!~��@��шo]Ω�D"O�I�'��@�,sea��0�A�T�ď��p=�"c�CҼ�f�*/����Ho�<)�ٙR30��>7�\ AD�d�<a4
�f�xTj���V�p#.`�<9����z�����=��`���_�<���݄;)J��S��W�X=:�ʏ]�<�V�H�~Z�P��ǰ
= l�KY�<q�Mȉ+�4(h'� -'�]J�T�<���[�$�I�dA�j���y�UM�<A����]�2m�H
&OL�BD5�ȓ"�䅋��Z?F�V]9"Ȍg�n	��dJ̸�L�`z� ����{3�(��zH�pfO�J��T�#ܔP��Ņȓ>�2��� ���1I�8'	�8�ȓSjʙBG�Ԅ-0ziucT
:����U���4�>!s��1�e��#R�i�F�<=��H�O��`\�(��!4,M��f�k���'�#i�T��ȓXZ]E 	6AϤa��Ƨ5���ȓd��SP�]�8���%��ȓ���#tĜF~\����`%F���aa�Az��?Hd<J�IW���ȓ�t0R�H嘍;���B1���|���ˁ�I�}�&$��Y�9��`���|�'bH��c��[�l������:a�;'=��wA����x���H��d��r1,��Č�6}L���)�H���
�L�U�&/�C����S��k�OA�V}�!qW�P�j�ȓ����,���*�p�cߌM��3���NY�-!�LЂLÉ-�f��b���%EQ;r��2A�XY����\�^a���*�G����ȓ%r^%`��?w�x=�v�]?\�<݅ȓ^Һ���,�?����![;c���E�&"��	0O;��
�O�i�je��L���W�+�F5���ĳ�Y��k����n��l�BIk"�-�(x�ȓ!���i�+XUU6�Y�MY�
"�!D��kF�I,l�ԑ�J@�G�Q2ń%D��r0j¡!p"ɩ�k'f��Ȩ�-'D���s�ȑ7���2b��f&� *�k%D��)�����~���&�T2U��h7D�\�C-�����I�Q�,Q��0D�̛�n�ꪬ�D�4?I@j*O�y`s�.�0�	�D�h���"Olu16�D�V��G候R��P��"O̜q��\����j�T�Lc�"O�p�C Q�f�n����JF��[�"O$�R`�4&Sx<�H� hb��c�"OV���9:�@��@%.<����"O�������\� -<[���k"O�ekR`�3-���cw�
1f�"�k�"O��xD�޿]�\R'��π�S�"O�S'�ĥ54��8�ȑ5-Ů`"O��mN�Tg�dx�(�O`\�E"O&�R��5�Ҭ��@�hHB���"O6� H-��Q� ��.2�쨠"O�uw뚋M�����)BO��1"OZ� ���V�9��?n�Hx�"OV��$��ؑe�O�t�ݣ�"O�*P��B�bc�:S�Ҩ�S"O�L31�^�8���a�W�l�:�"O� n���b@�
��3��#��x�f"OB��b��i=�T��*M}2lH�"Oi�r� |�� ש�	�j��"O %��%
+D�*D[fɑ8�޴;�"O6$�Q/-�G�9{��}R�"O�} q�Z��n9�S�ճ=�&�I�"O^�J�e��br]�AC�|P�(i"O���ˁj�Je�W�%)7����*O���� 03��r-[�cj�T�	�'�Б�o��2ē��U�(�R
�'�ʴA�LZ��ԍ��/܂L�&�[�'1�"eLO/�B,;��+D.���'<��
���"�1�V�Ң6�1j�'efU�wS'n��4�b]� �:,�'�ޕA�, Q:|�H$J��'�EX�'��4��LbE��t-�/u��Y��c1D��\� XG�,]�xX	sf �R�!�T9j� I��F��E�QfY��!򄝼.3��1��m����%Ŗ;X!�dN�oC0l�bȟ�#��r�T� �!�DT�,�`dK�+�"lV�eG!��*�6d'�,u�t�[��]�t8!�J5K�y@D6��}���e!!�K�|��	�nեW ��a�Ӡ{!�D�,{> 	S�R�f��8i��!���j�f(J=�޹q���3{�!�3��@���P&㾉�J�4�!���*&�(x�g�.�8]�����!�ħ-��������R����!�$үg����wȵ�th�1�!��bh^ݨ`�ׇM�Hd��i@�u!��ڸ��Dc$f�
�v��@���JW!�D��"��E��
l̮	����!�D����H��:b��9C��W�!�1'��4'V�c����"\|�!���!���E�\�M��'�T{!��@�T�b�Dr��(0?x!�D�WL�i�h #b��q�,
6vZ!�䇼#b���O�-���O�t��3�x�:P�
�H��"Ꮝ�\�책�RMJ�h!�"O���9E T�)�vA�ȓR"���*F*������[��]�ȓn����B%�� :�]�@Fכ>�hH�ȓX�M�GLL�a���c�0-��|匨�HD�I�~)�Y?b���a5ީ���L�&69*���<	���2�PrbO�u�șUCW:BZX��2�J��N&�>4SPap�|L�ȓ���턉W�h��K�BX,�ȓp$��FJǀ�T���b�n��._�����1I�В�㍙;�����i�R �? #T��Y�~(�ن�Z@n�k�i�1?:upE)Ǆ7��E�ȓ�4���jg�4��́�IE܅�9����7��@~d��C��+8Ԝ��}@�e��H��%��kV��Cp��ȓ��]b��߈E����C�}T��ȓP:μa#��6��"ю��
��]��C*����G�7]��kS������ȡ��EL7��]�) 5G*e�ȓ ����
�d�a� �8R0)�ȓM@t�2'�=��%����k��ȓ;�Ȣ��9`¬I;��ʸ}xFņ�b9�P2�CW�qo�i��e�;�t���S�? еa��v���ď�`�>싓"Or@2���X�v��@-�1	2���"Oj-Cf+S� 5.��W��7XD�H�"O��YFn�wM�<�����H
*DР"O�hzcxZ�:"�=OtT�"Od��qF��-RP�8I�G"O�8akI,�؜��Zt8ř"O�]��g�_r����-��E�1�@"O��6jT��8b�N��3|&Q'"Or0����. ���mD�y��#B"O4�`d�M�}9��&�۩rz�u�"O�<����J�zU�6b�	$iδ��"O ���C( }��%`_�v��dSe"O�9 ��h̠1�޵�Th�S"O��(��ڀ5���yPl�2���$"O�{B[�lTy�$�
�=��$�"O��!K �� #�]�E�d�A"O
M)���bk��8e��X�ܼ�"O��{�&��{,�]�v�V1W�����"O��
􀂩K4�G���C�"O2���@�,F!+�
#'
��:�"O�4[�Q�jI�\� ��]�DtKR"O��q�ZFLj�&L� ���3�"O�( +R4@�@� @�|ʾ�Xa"O��0��͝8Yr+!m�����6"O�P���T�✠U��(O�l['"Ol�S��$p��X#�G�D���t"O�M+HR�N�N�3AL]�4��"O�ezb�|��8aR%Ϣ�F� "O��q�J�i&��aҞ^��x�"O����ā_����6�G�C�f-��"O�Q�,C�!4/A�_�lM�`"O�6�0ѐq�Z�h���@: !��6V�ztV�΅e�v��P-G
f!��7d�ډ+3!�a�r�g�4o!�D��^�zš�Ģ/�Li�E�`!�ɏ7<��!
����S��<R��)�J�S��_ܾTp�kE�y��B+���qE���%3�����9�y�B��5��6+��F���k�l��yª�PYd�T!�8=�@��B�2�y��1d=$����83lX�0Q��yrM�'����F�_: i8@"���y�-�!"
�����Si:�Z��	�y�#��.�tT�$��`Ѻ�[!o�1�y"��=���
�#�N��PӰ,�y"aķ>`�`���1��`�w���y�Cƻq�q��!�4W�Q�D@�?�y9�f8CW�?\�,yN�yB��=x�P��O9���Co��y�9��q8T�#�쉃!ۓ�y�(.��	�3#E�s-($����y�
�.�҆m;s7p�[���y�&�O7`�YW���v�c�nɷ�y2oEk�l��S(K^���*���yB���9�:��gC,|�b��B��,�y���O��q��JC¥be�M��yrdN�cp�%"�z��x���.�yb��8
�zw"��n8ب2N��y�AI���]S�ᅎ�y�H1wWB� ����V��@D��y�j���H��1��1t����W��y������iSD&c{` �����y"I
�,�D��E�a[��IbBN��y
� r8JvE8+ EK���n�>�95"Ot}��K��Ho��'�$^4�%��"O����	]b��A�C�U4�p �"OP�%�ڏ��U2����T��Q"O��q�'�8=��-��@�R��C%"Oxq��̈v���B ��=Rz���"O�x�&ř//ɞD��m��"OZĺ�ύ��h�X��w����"O�5���U<f�A�K�9_Fr,j"O@(��ˉ�;,P��)"*P�Eb2"O����E�}H
�bsLh�-�"O(1���u�����!�2\SXu��"O��狖�9$��j�f�d8��3"O��
�,/� R�,fE(ۄ"O4պ�͞(�x�s�W'?2,5�a"OlZ��(?t\�j�M�u�Xh�"Oɓ���>#􀂄.�{`�h2"O��sb�ȋb���,mF�q�"O�ɨd#��W����4Xl@�"O`h)���-0�a��[���c"O ��%Q���¢�9�渂�"O~)3��+=lH�ܑE�H1"O�l{"Ǧgej	�D�a"O ��RB��n%2ޏ8j��qe"O z�G^�k#V��,�{T�@R�"O�Pb�İ5��T��O"^��"O���a�Q3lcFɲDH�,2�]�v"Of( qX����auf���R"O<=yG�i�����O��q�F�b�"O �qU䆵S�F��H�z�Zͣs"OFy�m�!s��A�-A(#]���"O���I����RFZ�H�"d"OZh�5+�f�*�!r��"0`젢�"O�a"�FPo�I�	ϨB"t���"ORy��GP�B)١i�
Yb�"O�yys��3nd�,>
��"O�q�F��XJ&TEA3H�"�"O@hy��L>����Ro�&Q��@�""O@�٧B]�t
�̂��>�.B�"Oƀ�`��kZ���á�7���"O	04�S
ZŪ��*����%"O�}� h�-�^Xۃ
՞f�p�"O���F�F�Ց�OZ8��pa�"O�ػ ��g��]� m[_}z-�t"O@a�u���h�L6jH��"O��q�O$K  -R
A[�LB%"O�}��
��(�j�h_�ddhI�"OV	y��� qP���U:Of��S"O|����B4rk��	7'7yMn݃�"O�d���T*���&HC�wFj!"O������#N�h]s-�
/����"O���T%ƚW���E��.���"O�̙�>
�:�X�+��WL���%"Od�`f�:3��=� MI�eJ�,�#"O�)A��;}v��CL�.f:��g"O&I����
�H��'��"�PB"O�yp���3=EN%ِ`��4�b"OȵZ�a#�ҵX��3�-be"O����T1{\���2a�����"Oq#nµ"j~ňF�U�*`�B�"Ox1x�F�(�!s����?����"O��6D)����BS"O�x5��T0�m�?��2�"O\�c�X�B]�M�,M��QӴ"O� jP�B#Ǜ ̜pص�ќ(�@�"Ozu���8�r�R��5!y��"Oڬ�W�	�vhJ�䒵D}�"O�a0u�X:ty`=�0C�*2��"Ol����_�xE{gH�,�I9V"O2ZUR���T#��ݖU��("O\l�H�+f�zV� wښ@a"O:!�n8,��E�,�><�p� S"OT��*0r�el�/	�U�!"O}K��]�m*�0!� ��t�9�"Op,�#+5��L����<���"e"OV�P$��/��wK�q`���"O سh�8~���`$�7~MC�"O �j�*�?ר����%&�ʦ"O��@�
x��Q�CQ� "�9�"O؛C����Q�Fb��#a�"O�����FB��hf V���"ON�֫�)�~�2sO� �нm"O���K���4񃭉�z�3"O���ĭ�A�nLSv��;��S�"O5��K��K<.)8��|�Bؘ$"O�l+qB �����1��\�N�"O4�{�&ڼ`�����a�zuI�"O���s�Ë �,�CF���<QB"O�h��d�/O�Vm��D\'z�LKS"O�d���ȴe�	�" Y� E"O�#���0� �� !��Z]��Y�"O(,R7ˇ2��ɑ�o2i�n|Q�"O���V;�,� ��o���s�"O�̓dc��J<%�SfڀK�h�
�"O.�9�& ���Ч��p �Q1"O�h��^�	~�I��Ֆ/<���"O䰁�c�j�$��C�G'����"O����8W�� N�.H	�I��"Ox��^?5�҅�g�����.�y��Z�2��PH+���5�yBʉ&9Y��P��'+dd�2���y�%Ԏ9B�8�ra�X��ȓ�ybAԡtҥ �-h����$�N�y�
!q$a�p� �V{��@� ؋�y���Q��ɘ��K�
	��۶�y���E�ɢr'��Jd�:��%�y�׈8��G0JHp�i'C�)�y�`��[~�|�R��!J��2'/��y"c��z&^��-
6P,	�nI��y�M�zs
y����|��P%�L$�y2���Q-�Pß�
��\�4 Z��yr��T`R��Ն� �T�2d��yR���:z�+c#��I_�����
9�y�L�uu�p��W�H;���y��7:�`��J,D�����탻�y��$ ����W�1�m��\0�ybݙl�F�#�AEW@�ɊGȞ�y"��(�h�gM����-�y2��:s1<��3kҀ��X�
�y��,S�*D�?�ܪw����yr處y�|p�c
� �͑����y��:i������j�v�1�.�:�y�'��c�1�K�e���Y��N�y�c�%1�P`�g�/U�
;t`���ybo�M朡C����Md��c�N��y��+2�
�q��2HAh��Q�(�yҬׂ
{PQ*�C˪�����]��y�`vn������`���HTN�y
� Py�!�M�`��W�l��đ�"O�y���˦Zլ�h���Q�>!�"O�Mp�%əN��t¡�َu�حs�"O�\�G&L�G-��2o01�
�&"O��bs	 <d�����4~6H�"O��a'�X�u�pj�G5ff����"O��a��-,�����
f }0c"O��5��4*�N�"��̤`e�� �"O��A�Ė|�6Mk�ؽ.�j���"OJ���"P�1K�0NBl��"OL)x���.AO��ؔ?'d�G"Ox�jTJ
?4I��Ty-��x"O,����ߍ��� ʇ��Za"OL�۲��#`&[D �-O��%��"OP���I	�,���OY3�:*g!�d�5�>uy1�$�$�@߿ Q!�D��`I�R��\挔㓡2�!�D�`�m�4����*q�Q.�:,�!��g@�y��
B���ؖFՐr�!�$r���`�GY�x��r��!�D�T�0��ԣ@�k��U$ݡ�!�D_�+��LP�����5��a��#�!��i�1J-�(a��K�a@�!�d���z�*�M�F�a��I�!�D�)7:�i�F�s��5
�YD>!�!.�����94�1I���;!��.7
n��QL�c��]�"���Py�K�}MX�҄,O�=&�PE���y2E�[�h��d�75�2��lX+�y��?4�A��[�&�4�#tm��y�㑓p�hpGֽ�|��F����y�ʘ�IO�=� ��p�s���y��:4 ��ƙ$  ��yӨF��y"MJ0|v�Y�C�zw M�	��y2�ʄT����6�Nt h(Jda��y�� h�d!��ޭ7gL�(񥆐�y2��+{�b y#��40Rh���y�Ȍ�l����#�<�3�ƥ�yҦ�.}�ձ'�G�c�:@�r�%�y�k.�pY:6h_1THp��	�y"ȇ/IU�U���^">���!���y��ґ|Պ���l��8�rA@�m�<�y�(J�kY��!֎޳3dĉ����	�y�&�:_��5��G�48�bP 0�C2�y��+D��1�ᤚ5���y'e݊�yb �1�*��7/�����yRc�KaBA�e�F�#�<��Pf�:�y�㜱�LD�G�Ԑۗ���yb�HD����V�D f?�`�ץ��y�n�?�-����+{�U�ۊ��y���2a D��s+��z�Ӧ�y���Dr�=�`��h�@�qSf_4�y��ݮI����cA�YH��S-J?�y��B.8�$��J��b+���yR�>z=xa˘�(�!�H��y�٭L��3bnW�BX�1����y�GA%<�Zܐ� [�R6굁`�]�y2���w��Rv�u�p5��Q��y�@B�t�@���M��V�� 4��,�yr�Z�?@��%�f�{rE�1�y�_����q@�;pz�k�ybO,xB � ��eA��1DB��y�D	�.�N�)&��(�D�1!����y���d����G&	�`���у�y
� r�C���;����Eoӌ�j�c"O:���G�2Ō�q��3����"O��K� �:!;x�1&K=�"4t"O��`�^�P�JMjS�8I�}p"O��(OG�t��C�$Ō)R6"O(���&	$����h�C��+�"O�e��8]���^�i,�� "OdT��@�/���r��6��Bp"O�e�򧟯G-
8C��k��ar"O�E*�j�L�.EZA'ˇE��!�a"O�l�Ņ12W�C�&X�c$���"O&͢$��x��$/T>w�.e*g"O$�(���N�q9��B
��xE"O�����#N
b�׮�n�J\�"O������,P�, �$�:�>��6"O.!����]��LF�~ kt"O�-[�H �3�V�� bκq����'"O�}Rv�R�6K����
�JU{6"O�;T%�=z����!�E�k���z�"O�aȷ��.d+xm�ƃ�Gf��"OvT���16��0Y1�@.P� �Q"O��� ��C
=x��ŧQ_���"O~�j$dT8v5@�0clL�G_nu��"O���G�T����G"D�BR.�z�*O�᳆�P\T#Q4:q��'�H1�D�XH8��_�	^f�	�'מ�A3,FJ\2�; Ǹ�l1	�'�5"��ڤO�Z����u��'M�؂��N�:��$A#O���ܲ�'p40g��X�2`���KYl���'���s��Ѹ���С��<�2�'��%z��@"�~H�p�����9�'d�M��葨c�=+��#ِ���'upѡB��P���K�����t��'�8�{gk�y�0]��G��<�8�a
�'����GG(=�P�Q.B�d� ѡ�'�Rqp1��>37�p�1��Ve�R�'� tY''��E�l�p�T!H���',m�a�ϔy�B��F���uD��'��ݺ���C�:�q�n��\��'j@�f��4����3��c�T$��'����$�!n�>�c�������'t�yʧ+A/����|��)�
�'{°���>zP�3`�=sM�my�'L:���	�K���뎶d�}*�'��T"!�E��0RU�C�W��H
�'��5��fb"ȘW�լ"�^��	�'��Pp%I0@W޴ZE׌m�,��'2(���@�[$��v�R+bhʩ��'/$���ꄣv���bG�ZV��d�
�'��!y�	�JXD�VhQ ����
�'���Cç�D�<`���/x�te�	�'���p�MB?�l(��Y�u�f�9	�'1��I �,byZ�0�q���'�����{��4�A�!nX)��'�:���"%�u�Щe6mq�'��0f��B�@�2P�H�&w����'M�k���'�h�J`�S$���'3^(�2d�Be����30����'�P��·X��z�&�*2��AC�'qP��e��Z]x7J\�VYq�'r�MS,	��QA]h��'�(�d�R{�Ne���82�<c�'|����� $4 �ԈL�-O.����� �u�¯��	���6�A�w@���"OĴI�ê`+\��iA69:�Lu"O,�r'NoD-e+Ŕ?��"Ox��⇗5A��tʙ�f�"���"OlT�e��'?�����Z�y�vP�"O��C�nŽC�j�K��R3�8�R"O�u�L��*���&��b,�7"OX�Bv��"PA.)s�*C
u>��E"O`�J�l3}��#��D��xSa"O�$��T$"� ���"�x�"O���Tl�T}��:�TP���R�"O����Fp1�C�'�n�H "O֬(D
,����(ޑD괥��"O���v���%��$�T���yռ�:V"OZ���ޛO̜:ce٧t����"O�����ÛHk�+��X�i�tF"O
��H�V�|[�`�'�L"�"OPI��c­i{ڴ����Ds�1�d"O�����;x�&=��!̿x
�\�"O��T�R�0h���3:Pn5i�"O0�8�Iޫ_
¥#`j�(VAN�Cb"O>T�������!�6]�1��"O��@DМt�}� ��,�3�"Oz�2��$CIl�A���N���"O����7�fD)q'A�#p5��"O$(s�$V4<�P�q�ř�,��UC"OT��V̐"9�vV��o9��RO�<�%C�C��LÊ�!0�|*�
�J�<ق����)0�dz���ul^�<q�.]�
��sul �\��h�§�W�<I���Nx��"/a���0���~�<�4JAJL�#�T)SU0Y@���q�< �C�1�hXp*U�yE!f�k�<�3�Y�X�ĘP��D�fa��HW �c�<�ff@�%����ɿG�:�p`�<qVR�xl�6�9��D��$�X�<y�W=T���Q��4C��0��[P�<)4aO�v��q)2�B�[�j4S×M�<���SA0�sa�
����gF*D��IU�[�]���8��V�-4N�S�(D��*ű^U�*��U� ,���-%D�q�-E�?p��YDT�R|E1p�?D�tREH���t��P�zJ��ǩ=D�\�C3��Es$���pRU�%D���T�s�	:$�[����5 #D�Tc�,�}y�A u�O |�<E�&�<D��2�-Sg4L�b����OB29��:D�8����Mh�bQ�X�
����%D��Rv�D��Heȥ�� j�޸�b& D��I�7
:n�+�(���b�0D�,�4� *��0��X=)S�h(��!D� 3��0~3�p��LW>Ub�\���!D�P���T�ڵ9Pl��j�p0�?D���0�;Ds�Q��^+B�JP��$#D�����[�:xȁ{1�X�@�@��"-$D���`ލZ�dQ��L{;�1�#D�drde�A=�x(�@L<V_"�3�?D�h���f�v`����sS�!��I0D�<�6�ŗj)0�87`��Q_�m�0D���e�T:��)�,�de��3D�$��.T��t,ѣ�Z�°�0D���G���L���j�A�)��Q��2D���`��)�0x4$J�5;�\bs�2D�p*�/M~�LXT�ýQ��jG!/D�� ��R�.o����!�HHP"O��c���0'���\�7��`y"O�%�� Ԃfud��&�A8/����"O��AZ¢!� �K��xY�"Od�9`�@X�\��>�0q�"O| �s���]��M�w�кe�杺a"OpVK�44N�$�0O;m��]�v"OV�Z���pX��CP��N�� i�"ODԳV��"#�Þ }HUY�"O��x�)�e���"��N�D~�\3�"O"a�tC	Z^�D��H�,Dip��"Oƽ#s-�2M\P�)Vg�sf�eX"OJ]Fm�G�`e��� I¹��"O2�hq��&��D��'�
j.�tC"O$�7��i�f�;�fc��2"O���4}�(�2��L�,ͮ� c"O6��d�j�b	����'� H�"Oj$X�/W�4׺<І����"O���V
�y��Y�����I��%A"O�W�2@>p��J�?�,��B��f�<�2�N�f�z@��$�!z��p��A_�<Y�
R|������͙���HE��b�<�b�  v"M@�CAT�!
�O�a�<9`NL�"�4M��E����)�ɛw�<�U��>z�V���m��&9���C��w�<i��G�rU�	���e��Q�C�<QR%ڈ���9����q���{�<Y%Bă'���"�<>�)��AD{�<�`i�&Q�v�1�N��knD9�E�N�<���د֔=� "M?Z`|��e��K�<q/�|c1��OӺ.I�8��l�<񭙣\ �0I�O�?bDx��D�f�<A�̧zAu �ľd�L�Rē}�<a'C��$�pG�~���}�<Q��V�r��yQI��RI���v�<A�ˋm�Dd�o��r��`��r�<��N7 ��EY!+'U�,�IF�n�<	��(qI�,E����!		O�<y� Q�0�8p'd�B6� VfHO�<	AiH3L��P����1@`u��gWK�<�5.Gr��s���+��i����J�<�/�!�J��d�� b��#0�J�<q*��uY���23��m��D�G�<qQ�ٚ-��$���/p������[�<�2�Ŵ%��AG�[��=�p��L�<A@aӐX����*�M3�(�J�<�F+��*VzE�0厤^b@e;FnDH�<Q�7'eb���N�iv��rq�z�<w/֘$o(�s0�Wv~�p�Jo�<Qs�%E���Rf&W�~8��N�D�<q���DĚ��"E �~���Zj�<�ŏ�pUk��Q
��D�E_�<1��T<}0uσT�-	CDY�<��o��-���C�Dٗ�UB�Z�<��$�e7�0qv ܍@<L���`�P�<!cB��V���p(؊D4"q�OAA�<��(#y��Kq�{��:�/IU�<)7�X'$8�3�i�,]$1$Cy�<	2D΀H^<�@�D������{�<�K�-/�\9����U��=@W/]�<I�/fs����h�f��$�f�T~�<�@
Ι8�����!Sx���/Gz�<Q��ֲ	�d�ৌ�6�ਠWd\r�<Aŋ�c
n��$��8T�����͌j�<� ��FJI�l/�xK1���f89�"O�1�oW�VK��B�M':t�IC"Or1������05gX��"Ob�j�D�^n���$K�dZ^�S"O��#��E?G�H���]Y|�"�"O�=IՎɅ���(RL�"O@�s ��r�\�X�LM7>H ��"Ov�CJ͎'�b�8��Z	�f�Є"O���3N�&!6ZU� �4W�� � "OV`�t�D�[�4���,T�:��J�"ODU���Ҡ͸���)tlx�a"O&GbU�j�)�Ќ�8RT�]�d"O`5H�aWDP;C�اVȱ�2"OP�t��q��;��G�i��"O�Y�!�&	N�\;I0H��"OFH���3%ʌ���p�$If"O 94Ge�d]y��ːF�X�2�"O���?*49���0d��tbp"O�I�Y�K��U�Ua� Vf�5��"O�X0���?xDjfo��l�ܰ�"O�l!ǅN\Y8
��l8T�@�"Ov9y��x�a�̀�7.	1�"O�����ĥs?�d���)f5F�8�"O�%4/��7���k���t9(q"O�$���8Ic�aѲ���p��R�"OęAD -3J��юJ�R���"O|�E�Ш0�f@�5��&^�X��"On�K���Z]�ǋ��IJѸ�"O@rv/шG;��7!�@�z���"O�uɡ���A̴07��:I��X8�"OB@���a (6O�9;��ԊV"Or�)�g�|,���ǤIk����"O�] ���ws�,�c��c;n���"O�+	��z�� 90��D"O�l�tM�4�~���*�)֪Y��"O�qyG)@�*sbEX��N8S�`�<!k��&��ˇeI�a#�dac�D_�<Q6*� 1,x$P�K�NQ�!�Ee�<QDJ�X��x1d��o[ބ5�d�<I��dRČ
�Y�BP	��I�<��`G	)�0!�cĉ,.~X�s�A�\�<��(�iE�x�o԰:�����d^�<q�_�9��KQ�Wx��0
Z�<�S�V�&�Դڑ�YL�� ��A�<��l�4�����GT�n�P�ar�<a'��CK�$ئ���b�"�#@m�k�<��	�d����T#Wު,�Mi�<q�Y8�BE�&.��ne�A�LO�<y�i�C� UJ� J0 4��H�<A`�P�:���V���<����ˆJ�<ysfA�H3��e���<���gi]~�<qUΓ�o��@�L\2Ws֠�@Mo�<)V$�2&z)��*{���{�Hh�<y�<OA�����%,�&]S`��L�<a��N/P| �J��"a�$|���D�<)�(��b�^,����b��lB�i�f�<I�(��E�|��r�-6���i�<�$�`�Ȉ2�@�sV��g×a�<q���.o� ��W��P �bv�<@@<]Bb��~Ap�*��u�<gB�=r:M a+��M�����T{�<I2��<h�gG�'\��qP,�z�<QE��BD�0Y���6��i���
a�<yb-[�]IV@8�o0.�Bչ�BFG�<� : 2�-	�-�q�3���+_B�õ"O4]Q`��o�i� �^�N��I"O�}+��U�_>�� У�4��f"O� {7L��;9����W�B�YG"O��v'�L%����^�<2���"O�`�+�<#KA)c?P݂�i���yR��:#��{��äc$�l�@FB��yr�
1����ʡ]P0DR�� ��yoZ�&ր1"*R8 p����FT��yb��E$rl���.^���*֦�ybԩ.y>��WbY�?�Б�B��ybg�>M���@ꁀ2�Z9:��J��yr�\=o<�ycR�O~��6�/�yR�3%8`��΢A����f
\��yb)�OT� 
�F�#E
 xnT��yW�s�u�aD�*'0HlHa���y��ѐ^$m(�h�OF<<�@����y2�P��D�o�:D �QJ
��y�a� G�6@B��B�N���yҡO��"i���r�)��;�y�#�_ sT �[̼����^��yZ:iQwJȽX`���Bh�M��ՇȓJF�җ�N	^vLq��̇R�B��ȓ X\X�-
}+p�a��܂H�,�����%!Ac�&(����a�*�fЇȓl�"A�M�;?ڝZ,�,����ȓ!���ņܢd�80BE��5|����ȓ �D�5d��}��"�/;�d�ȓq���{�E)z�*��RcY�3)(��+�:���NY0o(���Q/�lw�����(�2cā#q���e��d!��%"�s��)Td)��=fȩ��st����݌B)~ �	;j6bŇ�W���H�C�Yh�y�֌#�B�	N4t|��,Y'�<�ӄBE?�C��>mǪ�g�F7s��)O��i�B� D��`�o-Fs��h�ӻ:[PB�	/C��kW�G�V"){+�"�B�I�p=�°o�j{ڜH���/G�B�ɸ,ՀL�"�!hg��1zB�	�K��Ak�͇)K����C)^(5.C�	)HK���c�]���`ȯ/s�C�,:���`��+W��!Gl��?��C� �0\ppַJUr�b�Ϡx�pC�I�AL*������^)8)"D��lyhC��/Pqt�q��>L�Z�rB��g�B�ɍ<���v��z��Ś�-E��B�I*�) vgGm�]2�gR�W=�B��<E.�4�V�]��X6��Q?�B�	A��"	���
�G�/<`~B�	�NQ�x0c��0��te�խr	bB�ɢZ��y��F��P�k�ZB�I1&/^�)beѨGi�y����2ǊB�	K���'	�F���
9I�C䉊
]�XP7o�z��kw��T��B�IR�u:T�r�����,e��C�a�f`S�A�3�F���	�[J^C�I}�L\y1@N`�[3!���# hB�Ɂ8Xv�����@�L�!�By�C�I�i dȀ�i��x���qv B�]ۖB��7���!Z�&X��B�)<��B�I5P�ؓ�+�20b@P%͟���C�ɽ'���S3,�m1�S�CRVC�	�g����FA,l�ٸ�#�hC�)� 6d���̪xY�%�Ů+p�����"O:u�č���$���DC"OX���0�r�k�\�QOn-*$"OZH�vfSO�\(@G6w�ƴSc*O|�9��>��M�H�st��'�P�"�JP-tY:d.1yz��'g�hyt��Ŧ=#��.H�r �'3X]� �[���� g�9�$T��'����''`��(R�H�{�'7�q�F���H���&AZ��'��`����0���pXKjn���'�r �I�(���=�@�q�'N�mZ4��N	94��aj����'G*]p1��@��Pz�	�`V�'��a�fan�0�Hh�
�'�J�H���<˂��-�ؐ�	�'
P� g(Y�.4V5��cW�n�F$i�'���Nײ�H��xú<��'�*�R�χI��0ⓧxb�+�'��+�a�"��k� �.)�	�'��Uq�)�a/�LZ�#�k�Z��'�V]3�T�%5P�M=W'Z���'�H�����a�\@�`�M`�!0�'�B�c�M�gX�<��6OȺ�#	�'��` �O�n��a:�8�����'ٌ�k�n��$����q	C���M�
�'���B�σG��I@�Tw' ��	�'�z�y�yH�kf�Vu�L�R
�'C�� �� �S6���q-(p�	�'�����%�h`hv�� ǰ�Y	�'K�m�瀛:�H�V)��|��'{�@�C�5N��`c�إs�&���'=���e��?�~铇�� z�y��'{�y2�'"_��PPl��*�H�'� �"f���qhH�BPcͫ-	^Q��'�
%�
+E&h�f�	$�(��'3��#K
'BE��ɐ����'���q��ZBaQu�.[0B�s�'Vj�)�OD�U��ȇ�C�d
�U1
�'��L*�[���hw�
�Y�� �'Ҡ�ᅪE22����ϭS�t���'{��[�J�,x8��x�A�|���'�+�,�4nh�5�׮n��QQ
�'�T�3'�"L^�{h��S�21�	�'�j�� �: bN�q�D�K���	�'�*�#΍`J�#C(�=➜��'��:�
J�O% U0"#K�dD���'�Tu�m�7�-�Ȓh��9x�'�h5,݃(6�����T �l�A�'�A2�iUfލ�1�"� �'Vx�b5J�{�T��T��N- �'�:ة�M^6{�!�のr�Т�'<�!�Nv�ZuY���b�d��'],l[P!(�����%�	L�"�'.��c�̙)�
ͻ��	���0��'H�PEd�55����OM�RI���'�@�S��:^yƙ�#�@�C8��1�'i�����M?�˲�C;0��'�H� U#t^�x��J0�xP�' @�p�V�V�v�h�"�9/s��'1d������L|#a�?O��	�'c`,�uD	%L�Piծ�`[	�'`j�5�M:yx�x`/A����'6�Y�!�3n�(8�c	57��Ѻ��� Ea&!�(��Y�����W ���"Od��f[�j/�=r􏓇9BX�2"Od�jRD�
Q�`��۩H��س�"O��zՠ�y�X�+�A�+H��2"O0�*��	��`�A� )Z{��U"Or%��NK�_=��Bp
�����"O�h2 딱?B�֨�v���W"O�Ib2�6��Ӱ( ���d2"Oؐ�g��o2��r�`^���)�"O�0��I�-����^<[�ҁ2�"O���Wh��g����<�,tC�"O����ی������ί@�B��b"O ��%�R=i�0�q� ć`��	0"O��S��߮J�9�H��,`�"OHxjҬ̀�Ji07�K!&�e�"O<�"u
/P��� �L�D�B5"O�0��i�/P�p5ʅO���`"O���J�+�|�CAG���3�"Ox�K�lG�Z�|���ìJ��ж"O�k�kJ9����v�W�jt&9��"O��� ˔Wߨ�r�C�FQ�3�"O��i%��7z-P���pи�"O�������cJܺ���4Dg� �"O�]W˩.�I�4a� |�P"O��b%�	FR�8ZATae̸�"OP��ԃ�U|��5ō�(�%�"OT�.޽s�Rx�aD�/3��dj"O,�i�����Y�hU�$|��;"O6iI�&3u��=��3'q���e"O�0���S��Jm��(��r���t"OR\I_�+�iXUNJ%�0!z�"O��I�e
�F!2Q�DL�L��[�"O�1Qp �2a��$���ݗz�\�s�"O�}���s	D�)M�V�4�&"O$@%�9�
�rl
!�� "O�L�p� �bZ���F=�80c�"OP�����=�B<�Bk�'>�L؊"O~�e��2<��!Y�h�csd-��"O��)gň�r�k���]C@"O������2"�E�7ŝ�hA��X�"O�(5/�U���2��$
)��"O6���S%�t��qᄆF/:��"O(8��f��oՌ�U�I�/�dXk�"O�ѣf�_��$�!t �+ݾ	Z�"O��{�̀.m�lx�`�-z��`[�"O�Pf��r�%11�qۤ4�b"O,(�wE�P��M*@�@4wi8��"OvQ���"��ـlJ�[L���"O��R��0K+5P�
w9�蛑"O�!-��-�\�6 K^)��*"O�U32!̚
���CE��,EC�"OzMї�ӕl�i�`��Dl� �"OQ����,�r�Q��ڒR�$��"O��+aC��/LN��d�M�B�<B�"O�hq����!�2���,He�����"O4Ġ���8����K��Qr��8C"O$Z6/�!.�H��U7�(�B"Od�1u(	J���#&o�Sv��0"OP����9l6�-�?A��kU"OhD;�[�[ā�lG86�=�e"OީJ�D��8��m}�t��"O����0�z��G�48��*�"OnL��
P�[��KA�?!��Ma�"OpJ���h*�`�##�� �"O� �Hs�L܇Ci�a���A��T4`�"OL,���A<=�����+���"OB"1A��C;�A���x� ��"OB�@���T
�F���ii��YV"O��:f�[�Z��I�S痸4��"OJ�#�����Ć�0G&ѻ�"O�� �<jhqgԀ��`"O:�1ՠSqyjh�g��� �"O��P��#}���E�*^�X�g"O�@(s�9h�L����/kD�@w"Oʐ�f�,h��9�bØ{����V"O��hC�-gո-�gL����;A"O�QA�P	r�p�au뗬Zqz�
�"Od�(�gJ1�4��
�{5�� '"OD�r#�.Np��eJF�#��Kt"O�t��<+�� A�ӊɃ�"O�1� $F"$�Pڥ���4!�A6"O��rc@�Mς�K#�� ̍I"O����-�@4���[�Z��k�"Or��B�^�-�\�E�?)� ��"OXl�Po�;W�2�ꑠ�r���&"O6���M�7Gn��4-�.��(�0"O�M�PG�z�l�Kӌ�ܤ�"O���V�3o'@�� X1Ic����"O���F�̂nU�L�Y��lpPR"O�d���3ZN~hE�y@>@�"Ode��!D�#�\ Kd�SV0Eu"O��PB�j��t8��&>�l��"O=1��E�;S�� �[a(@���"O���$k�){�	�Q�����W�<I�MI6X-k�22h��B�CT�<A 
�9g����N�(J.yQg�Q�<��,�	A5,E�+b��!�s�<����S:��g��jF�@���e�<�g`EN�:уO��N�x��Pk�<U�>C�����*,98ǘe�<i���1	�$���+�(|�FH��b�<�e�@�dQ��c��q����d�<�� Q�6���+��@)�x�ISDQ_�<Y��̡3�rY���
,|�&���W�<��囤�%��n� 4d�!�S�<y��A1T��e���c��arq�O�<�ċY"=�� �v���T�Tr�jGd�<��DXn/��s2�B�*t\�	@K�<���..��t���������H�<�e�2)~1�ϊ�c-��C�<��_�z�(��Ɍ.l�����@�<A&�^�f$�t��<�L(W�}�<A �!�$.Vj��qE�v�<�kWGBΰٱR9�"�[�-�G�<�ԧ&#]�uB6�J!>-ftk���C�<iE��J+d�)��F���th`ŇC�<� �B��^q��E��OY����AV�<Y�����A`򮟘~r�|*��z�<aQ���rQ  �C�u��Hr���u�<ɲE@�Z}Xr!	�l	�(�RV�<�q��{`ucS�� Zbj����y�<��[ �
�Ռ�<�d(:��
]�<15�\�U�Ҭ0O�6=�H@3hZ�<y��]�`@2�R�)*?��x`�X�<��Gxe��jbJ&b5�A�)�R�<�4�J�	��4�4�Y�X�4�Z��AH�<ц��3QH�����s�^�í�@�<QF�D_�!�'�<�p����g�<� ⠉T�Q�.]�-��НS��pc"O�]��B�VJ�4P� -g�1�A"O�!�ɝ�\J�XK�-Ԭ`�d(v"OT;U*Ʋu랴�i��a��5�u"O�)2�jۗ=(�(c�g�!|��1"O��B� @4'T\�'ޝ[Ԋ<�"O��cs��NSL$�� �FȲI��"O�,��*C
�b6��qk�nZ�}!��\82��"�π%&ڀA�j��I!�D��1�Ld�DD�t���Y��!�9Bt)��<wȰ�;�A�/w�!�@��Ԩl����}�Tb�7�!�$��3?X�IN�/t�ڱ�A,�d|!�döX��X(2I@���y��Md_!�đ2E1��Q��Q�Lk��R+Q�R�!��_iJx�I�"������˷�!�$V8�$��,���Za�O�-#!�D��Nh��v*�G�n�@҅��C!�D�ZN�!��+݆��5�b�şh-!�dP"s�d���,y�����!��CB�Pի��A�j9��)�o�V!�D_9Z�x)r���6����.^b!�"*�%IS�N$=#R��L�8�!��	�	��awO_%w��,K�K<?�!�䎀F@t!a!�nz���c�O6Y!��֤T	|���Υx���Z�ssB��FH�ḗ�F7]���2�)�BB��.	��=c�釕K�t��G�;B�m��+2�5_	@c%NK�C䉕#X�Tї�L0�6��S�˃:}`C�I5�X��$N�2wtQR��yU�B�I�w�Z�{ΕT��X���}K&B�I�B�,�E�{���aݦc,�C�I�l�h�K�Ei��qc���C�ɴ-��7/�?hg����]�C�	,?d�h:棃Ұݨ�O'L�xC���8��ǯ^������WJID*D�`[�L�[����'S,Y׮�z��)D�Ѓ���:Kv���WP�y�,"7�'D��󦁃fa>���&��k�Z�*aN+D����#ɛ�T0RE�ɶ
�R��(D��[A�?g��c�m�s�>��H"D����>{����K�@ypO2D��ǳZuN� �&|s"�q#D��F.ʈ
�\̺�fK��2�y�I D�@CvN�7mnaR���L�µz�>D��Jv�-Fh,X��:���أ�}��b��K��>���+H�. �.�3l����r�<i�gS�]LB�jӤj�ҔZ��v�<QLиΰ|K�ɺV��R��p؞4�=	���.x�"�h�4j�r!l��<��~�U���y8���'}��q���l�ɝ8P0��U"q� p��J� d8C�	i����D��g@慘&L�O�4C�I'l`��%�xڑ��C� 5C��7&J�ಳ*/����p��c��E{��9O��ۣc�,=������4h�:���'��'I��U@(L�@��7��pk�僟'���D�^��]���D�VJ�\�t��(T��O���}b��bĶO'x��̮2"$�x劙��y��	D��!���06� ; �ܨ�ybƙ�p���>-�d9 iK
�y�pi�8�U��,��u�F��y�M	p���jU�3F����y
� бY3��D6*k��E.-�@}�"O�������6=�$B�B�H����'��I>uUT�iI$�
��˒�1��B�I�>'d�a@Q�@��PR��u�xB�'��&={�x	듾;�C䉋Y9���G�/�xL�*Ъ��C�s.�� 썬.��AEώY��xr�		2��A+���%�EF� xj(�O�������HK��J��a�!Go!򤝼n���vC�W8pHB'V-kz!�U��D�U#Ѻo.�	D�KvqOB��R &l1M`��y�UdPbd!�dW�ִ�LT��B<���@�Y�IH���j]�֨Z��p%#��%x(��[�<��I�YɈ���"� $���n�u�̰=qլ/�UJ)S Q�ve�
o����,�d�-�Uk��n)q����,�ॆ�g��sƆ�oXP}�ѧ%J��܄ȓq��][&�+*�p����J�?�	����?���d��B@�Y�6M�ѩ�#Gc�ČS���O8��ի>)*��@	� mq��'[��R,N��ι��E����'��tA</V@1I�"�F���'�~��	��z�f��q0���'˂������h���f/�5��Y�'6Z�{wŚ-d�@���:.�(R	�'����%ūI����Δ��	�'�11'�i0`Q�h�� hi�ϓ�O���b��7:��ctjE8���6[����1|�P5Ge|Y*dߞed���	.4����cjB�u�6I6�x���QgzB�	�0�J�	Hԝ2��,#E���O.�$�O�O��S�t!˩:�>@h�+7H����h^��y��[;;�ks+R�X�b���ꍂ���=�S�O��I�2�ǫz Y`Vo���6��'�"�S�� F:��Ơ��+	�'���PLF*,� �	��{<�3�'Q�蓰)�6+��yG�]�mu�و�'Z
�i-L�w���1�Ad��z�'��H�Yj�m��f\���Z�{�<a`(
�hd��BYU$1�GA�B�<���÷^$V��pa��RG6�9�@�<�!���>���#�$�1K��$��/y�<�RKL
�x�*��0A~\��f�t�<� E�~0�Qz!Ȣ� �rn�<	���  �50Ň*���@���h�<!ᮉ8l�t��nԔ %L���Xe�<Av�Ϲ���G
�	^�H�CQ}�<y�����d���h�����`�v�<1"jT�%��{����tr�BdDOp�<�ШΈ	�؉À�3hb�*���g�<�cƔ+6f@��!G�3&��z&��M�<�a]Tg�����د�]� '�o�<���Rζ�g��g�	bpHk�<��F��^�V�ߑ�qVn�<��G	H$�QA�'R��11ԉMc�<)V�"@�I�R�ܾ�d-y�Eh�<)�,���G� :u�lᘵ��<�ׇP3?�B�X�W�.��l�aKw�<���I=�3�5.�0���Zn�<�$K}#�Y�k١8�9��$6D����nC9u�FD�t�m	 �{b6D��Y�AP�e(��2�W#(&(	Qg2D��B����h���"9K ��r�0D�� �|��'B"W�>E����#*���$"O~tZ�eˮ���G@�A R"OzH!���n\4���uI�H�d"O��86A֡c�����G+1Z1�"OԌ8v�/F�xx�mԼ^ ��Br"O�UȐ�#� �9B�.4��f"O8�DC5�P�!�S#/ ��*""O���
�0�*�93�
{���0"Olպ6�H\�PT����+ Xa��"O&d��d� �n �և�

P�"O&�ɧ��~�Ԓ&1��#�"O쓳m�%8B~�*g����pp&"O¸��h�9P�	�ᣜ&}R��1"O�i����#TV�*@�qW�ĉ1"O�E@�ށ(�e�v�ѭO���h�"O����.4D�8�f ��q���P"O��$Ë	?����,^0Jx)�R"O(�Ze�&+4`K�Q�*��c"O�ś0�˲b�h%��D�VX��a"O��(פ��T	;Dݴ�S�"O���g2V����A�L�xE��"O���͕	D86��˂���"Ob� ��F�\XBmT�����f"O��� ��I�l�eK{���jf"O���Ҋ҃IW|X���4x���!�"ONP�#E/0��9o}��YH�"O��@��E�}X�h�9L�h"O\��%N�/+GڈI�GG�[����"O
�1�n�+�X|�el�=�*`k"Oܭ*�I�>]���'hp�z�"O�0A�I�G�.�����,s(�(Y�"O�ɓshU�m>�:t ��B�BH��"O}�%�Xa�5AF��V�JhiA"O4�
ӈ�`b� ��[�� <�"O�a�#�X���T(O� :�� "O:�ˆ.:�����y�.�:�"O����GK�5����g�,}��2�"O���b�W
����taV;F�n���"O`�)p���e���#�/�����"OR�G$ܜ@��غ�E�P�@{�"OxԁC��=�~ ���r���"U"OD�Rwf�G=���M5'�*My�"OX�)B���4��s�ϒ6L��a{�"ODy��k�"D.l���dNO�q07"O&��aрCW�d�H���z�"O�4��W�P��\@�'�'W��I��"OHD����v�މ��$�*K+�	0s"OTA3�OU�K��H �n�#��%"O��#��B�GM.y�҇I-Ue��ٗ"O�I1��ΟZs�@p��Q] �d�A"O&�兎��� �C;&up�"O�)�Xi��`c�+<
���"O��K�&re�M�� ��g�L\*"O<lC%#� ��x�u�űIw��Ȅ"Ov�K��B�Z�B���G�gi�IZ "O�]Ѵ�2|).�`�W
�#"O���PO��٘��+!E��"O�p�	D�0�<�E�0+�츁p"O��8U���Z{p)�kD2��t8"O�q���sr�x��	R)C�.��a"O:q�Į�F���+�iTl���S"O�e�%lOgB@�y��M�G� �b"O�9�'�Duo&`�&��#��DR�*O�y(��Y�|b������!��A	��� ��+!Y/R7��e1"�
�:F"O�0R�gW��Sd��uѲ���"O��2�Kփ0@x�p΁�-�J�.�yRk��LB���w_�n �(�����y�	!d^���eA`�򌻦�5�y��]6� �!�[+��I@F����y��-��qy��ܩ��Ń�z!���0�L�#S@ 3b��|����7!�f��4;3��>�4苁�W&�!�dՆpv���ӳ���JȻfu!��N�p,H�TOX '�@�6(J aV!��Z�baQO�w � S�B�:K!�$  Ϻl(��Z�f��4�@�!�Ēl(�@sW.�������)u!��J�&>��f�.��EW H�C�!�d�+o8�Ar���<�x��4�,*�!�d�(L������.>�zD�@6�!�dS�ר���.@�h���Z��
O�!�dN+����.��Aƍ�,f�!�ę�`,�O�9o�Z�a��ԘX�!�䎆j�%�c(ɐ�8��M�e�!�dC<@��}�W�
�m�dEq!����!�V	��,���J�h8����!�K�LR�'�(hcaT	m�!򄖝_�������4:]
�3�fH�
�!�E�n�@�����4>��A�+�/g!�䕿>44� p��$'�.q��	���!�D�ٚ��ЫD����0hU�!�}�>�Б�'u�&�y%FuE8��<|�;�i¨z�,�p�Aޑe����m�L�s�ȏ�f����%����r#Xm�PdT�K�ܩ�J�wO����r��YB����D�&��2��r����dY3FɁ%m8dY��i����\������|.�<Q���y4	�ȓL�yӅ�X)�����7D"�m��h�8i`�P#E���S�?���ȓ^��9�G�ĐVٖ�HQ�A�n��ȇȓ���v��+��A�U -����ȓ)�q;�g�F��@�h[6��l�ȓBs�Ly��ҏI�A����Uf���Ȏ +����G��%���ܐ2�*	��=m���paBEϚ)�V&ڍc�Q�ȓ~X)��B�|)̤�Q�Ɋ����._��26d�� Q��1����;��2�.i$��#��)!���,:n݄ȓ]/���'ŃsY	�BS�"�̄�G��[AW �� �c��<&f̈́�:��Ze��'Cl�؀���f�q��	w�'V����D�05�w��;N"�A8�'�,؛�HC�+`Hp��(�@��X�'$�i��-X�6+�����%@�e��'�eJ �
�U'&7)Cw���P@"O�����K�n\Г�%)����'	�'olh��)�t�qe�_=9�>Q�'���&�$L�X��V��O���hã]��y2��
x�[��N�8@��B�yb U�o�H2�a�9E��q;�C�y��\�P��ݙw�SM��y�!�'�y	c1��#A��	L�� !��J��y�e�!O�uе�T,=�d�0`Ą	�y� ^>gJ��2J�1��1��Ƹ�y"��
Vt&�Q����1{(����)�y�	�
�d�S��/ LA����y
� �ě��h�^�#e\�}H��9A"O��J���2Q\:,PUǡ8j���"O�u*���;p���F��/c-����$ |O�M�d����9Y�&�huD�۔"Ol���;"ɓ�c�10h PKs"O�#�a��(��Q��J\X���"OQXj&"�p�J��@7ȥ��"O�e�k��I�D���p"O&��� �	a,I�r̞����H�
O"7��`(6��JV� ��x ��T3x��hO����w�Y#>��V!lS�	W"O����2e!\���B�>4��C"OęxEE�	"�(���,P��h:c"O�݃�C2$X��R��ƷL}�cc"O�e@��W>G
u*v��qf��bW"O���� _�&0ycn��Y��4h O��P�Öf� 8��NõR��]��+k��	�k�Q�"|b,�92.T�A��A�ܴ���]��X�<�#l؞%i�!�	�M5���ġZW�<����J���R�/wa�"Xx���d����|�)�}�	�RL�
�Fd���ձ�Py��
�A�V1��H5\�̔q�k+�HO��=�OI��+�Ȑtj�t#d��&P��̒�'��"c�Cƺ(�K�y�f9��'��}�kK	s�&���-|�@��'zਓ��ͺP��p�\({O�=��'?�(���˳Ni䴠g���	��'�����B�֡�!�Y�N^ͺ�'����؈�M�B� ��'_�%K ����  ֩H�� !
�'����S��$�J�� gǭ>g��1�'��c��_: t,��"ݍ+JR�h
�'8<�`d�jږ|#�I::���	�'��p� �G)j	�E��h|4�	�'�|�`
�r	ؐ*�lU�/%�4��'��y��"
~*�A3uM[=Y2�'�d�ǏZ�X\3�eк;<��'H�m����!.P`�2NR\�p�1�'uƅ���Y6�F�PeF�G#pU��'��,���%�B����F�.�P��
�'JB�ٱOU3a��0a���*�$��'3�P'�0=xLڒ���X�X�'BR�#��Uߤ�*g�
=���'�F8yKB���$�6�V�+�YJ
�'Ez9jG�A�rމ���;v�
�'"����z���R���8%�đ�'kT�{Q" ��|z��Jb�t�
�'�^�[s�P��<A��_~�
�'ff�FDãUp�\ �H�F��
�'��pÅg(,�tq�B'L���
�'����d�9_ʱ'	�T6\�
�'�4%Dߊu�p8'M�t�Č��'�8��2��#H]ڽ ���r�����'�ZeQ���
.}�P
�l+
!�
�'�.��#Iƌ�6})�J�7c�B�S�'ꐩ��#��-�M��#Ї� ��'�J��0
6� Q��� �1
�'b<�0&ϗg�PE���A�u`��A�'��dㆍ+��|�W/Bi��S�'�TB� ��q`�6*8�(��'�J$ҒN˴Tktd:Sδ�L���'�~�z�IS (�ģ@�0�P�'�d���&(.���b��L $�+�'��܃�ŏ)G~��tMں<$Ȅ��� �d��+�-yb�S�(S5w�pQ{"O.̉$�  G�q��Ƌ�I�r�!�"O�E����T&<���#[�$z���C"O����MB���y�M��j,1"O>y�c�	8C�u��6ql,,�7"OBQZ�`Ʈ5��4+�? i1"O^)��OԐzQ��[ %���"O�H�#(E>YXr霡
�ؑ�"O�8 ɱEa(��âM2�L��"O�e�G18L�v��k�.��F"Ob=�4�;/Wm��k^`l��	V"O��0���7n�h�[Rk�e���U"Ȏ�/J�1�2ybGW;6�ec1"O�x��A	8^���_Gf�"O<��e�Q8j�4�p��,x��5��"OP񗩓�!�a qc�(_L6ؕ"O���ǎ`'j�VH�P�(�c"OPp)���� ��(`GB5c�M;q"O>� �Eu \�R4gηJ)n��`"O�ʣ�˭eUJ 1	J*7�q�"O� J�<EX�P�DX
�4�� "O�1�	Q+��pЃ�R�w]�q24"O،i�(�E���
0�?i�Z�C2"OV �!]�3Ӳ�KUOJ�
�zM�"O�P�	�+J���v�[��A*�"Oe�F սK���i^�>Cd!ۤ"O,xG�Y�8�h�0I�?GXH`c"O�8!#AӋ?���#�S+08Ia"O�5;�G mS�tq��O�LD��v"O(]��T�?{ pP���;n���"OD�3�k�_���� �ɳ�"OD���� E��E��Hh��-�
�y�D��xD��)f��S�5�󡔿�y"��!��	�R�Lx�L�y2( �x�Z�NѝK�n�rc���y�H�8;f0��T�B���R �:�y�,Ԙ*՘��I��:��$Y�eʋ�y�c�l Ȧ��F�.i
1���y��X7.OƜKҧ�;1���@JL��y�=\�q�ӤΚ��� �y��=K����DL2t�2���E��yrŝz���A�J�d�h�G��y�KV�n�$�$�@�J6|Yc$���y�K[�C��9���5=-\�҈���y��)h�ȅx�l,M�>�a��+�y�c��fb$lq.L�W�\��,��Py�mD�/q�1"d����H�#+d�<�oQ%t��Ը6�[�c�j|KwKb�<9TBG-�hQ�s�К�R@#���c�<i�̓&i�Nx�Q�U�=uP�����y�<���cdtJӏԼs�F4Rb�Lv�<ٶ�ظJ���� V6G�@�Yv,�H�<qU��'^>�	��ׯ<��y��@k�<�E ޖB:6��*K� �[2lY�ybCGl���b��,Cu���R��yB�Z�gm�}²��R�!�;X��p�'��/��,�~��4Ke�]��'k����/W�l����(<�Bт�'S^�IB�	�U���u�� 8�t�+�'�(���� \9�����O4�f���' �9�#�Ѭ3��ȢfIO�XM�0s�'ʐ��ҀL�Vu����#�Lɲ
�'eHȺd$� B��ɆIA8O�P��'�8YsR�N8����I#1���� x6�^
�p������"O��bqnȲv�PIC��U<Lu�"ON�p�١{g|ب�&	�a�P"OڵY��.i�����T���"OB1��i;K�<;ӯ�Fq�"O�`�@�޳Q�Ɂ�_�R_xv"Oj�� �P�s�h�Ib.�rm��K4���B�j#��`X'F�?C�t��-2?l��FZ�o����⁪U�!�B���K�����ą
���;�!�DK�:l`%�����u�C���L�!򤔦C����!�t>��bf�M�@p!�$��(��d�o�-K)*��[&C�!��5Ypx,��a��T �`i �ז*!�@ ��Y2c�g��!�wlD�N!�d�9<���bŗemCq��.!���A�V� d/�	>%��C��!���H�r�s��"+R�Ԣ�;�!�Éa��B2`���!���?�(�cR�o�b���F�YW!�d�72$���V�4��4����$d"!�͋'=�q�Ԫ^�V���)��5!��U=�����LN�
��
�+ !�D��lO�!�l¯B!����GW!�D%oj����97,ޘ�w>j\!�����'hфK�QK�b�"NN!��):�9ӳ$��k�J8���(`�!�"[%0Pa�i׈m*a`ь�!�Q�^PEc���D����!��m�!��؂W36)��R�2�x	�$�9�!�L�W�e�1iD�=�l�nۇ*�!��P�Z�0�م�\>+��]����Q�!����H� �!�b!�S�D�W/!�D�UW � �5d������(w6!��τj���'�K����a�x"!�^�8O�S"�:!�6��d�5H�!��M�!��<�3Œ�Ν��O߯�!��)8�jA �Z�`!2M��Ƭ�a~C֋Y]N��
E�:{����ï�z�AgH��y�f��>	h7 W�|�*&���HO�h(Cf� ���6�Ә��)�ᖋ,"z��Ģ @�C䉄|���)��h��r �%V�M�WJ�@�����A	-"�Y�)��<Qcǒ'�i#�*RGH�	�b�[q�<!A!!�lE�p< ��bu���� b�V��.L�c�˭W��T�3�F3�хǈ@g`�k!�(�x��I�x/b�+��+�vr�&���9!-�|&VU*�o�3� Pq�*�Y���Pu�U;d@{:$�����tzm��{B	Ϻ�<a�1�ݩs��<+��Ѷ4���O���yWmJ$z�Ȉs�.O�e8r�'���K�,U:4�Y¥�=��KK�0�FI��#O�!Z0��p��ث��4���y�D�L.�4�6mpg��x���*}����Z#9����=�2���Z�Lɸ��H�+|Hv�C0�� +y��Ez2N	�|���#D�B�HQё�ɵ��<)d�B�DM�1C�6G�X��*%�I�-O/x�*f��o�t����m����Ą0I�]AB/��d���/�b��x���{4�ݨU�d��%�"�_._����G#ڌXC�IM:eM��p�Ë!�<�#�M��<�!��"m����Ǆ3��U!��7�T�jR�*K�fdh�J[�Wq�+��PYS8ﲌz�a�z_
,`v	ŧR(�q��O\u�5K_��ܤ	G��)7��A�&)I�Y��M�!��u�N�*���j����u��5�̢<q�DF�k#*�B"�A&O�P�Z��ZMX�\���H�O���"�ζB���B3�xh@C��2M�� �C�*[8�PI�6��!��@K&�3���wM��e�ϕo�.�g�t�{"G .8x�\�ա\�#���9"y삳g
7Z�R"��	V����U�(H����3�ZC�	v�6l�"�O4��`���	!�� �(+_�� �눂"������w�0`��4��xҌ:'��);9(XX?W����Dq����
�>�t=S!���IP �M�}�4���m�ڄ��%`��G�A�*�DX�F��lV�]`P&M0y���/D�k���S�? f����E�#���9b����剚_`���b>&���n�f���!�G:_"�����#W"����-��`cD�-�v$BE�B�
���
A���7E�8D~b�7|6�W(Ԕ;����#�7M�\�P��C
r�LQ�#� _8�]��m�1q,�p�h��?��	赃6N�P�@�bǩy6��bƓ�6Rr�Td�@/|���A#�O䜰ǯQ�>�1����p��M風΋��a�1I]�)�'�G��12�1�$�� t��U��8��|x��˿�j��.�F�(p���'3� *$��UjS� �&lp�l׾
�<���!���f���~�Z��h��G�5�\96K~S*0�3�#��	�-)���v��#��p�V"N�N
��������sS@�[a�ߧC,����E<� �QeD<2ᢅB�fkhq��IN�phC�n�)W��Y6���M�����6鲙F|�@�Y���Y2鋖f(���9q<@�U* ��X1��C�|*p�[w#]�����J�e"��G�;t3d�E�ޚj�8�a�" LX��H�}.��� H3�0?YCc׻Tf�P���g�r��"�A 72z�k�����(vK:-l���Sl�0	P�K�c�n������߹���	r��l��L��A9x �F�e��� �#�1;c2h���
	�dس"U,lV�c4 �-s����q N;$H�*AF�:@l�"�
���x���խkX�[D��p����v�0P��_�U��-��)�ܮY�?����(�M� '�,�\�c e�^�E����	C�p�X�>�c4��JP���#6��e�<@�f�4@T�_E�#���אb=���f
6m~Y¨��h�~��K�ik�� c�Ɠ!����*��a;���V�H4ixq��آm�`=If�ɶz�p���a�<B44P%G��?�H�Ǭ/Xa~"�L_������'˰��ٝ=��x�e�Q-���B�
3Ҏ��S��Z��'����h�����/v�Ÿ�V�BS6$�1��>���Xx����9L�p�
s�2����E� )���v���2��$s��=7W|����ܦ��e&\�g	f��W��>EZ��ӭ��@���ؖ2�X�Ąi�zԣ�"�z�ZP����)D:Ѧ	�f����ą)Zks�W (wFI��p���k� 6(ly�`�sa� ёi��xS�"�s1޵q2J�ԥ"g���h�;�]%�HYѠ��+qst����=v>ȩQ
���ݝ^(n��e���rj�q�^z6�"�k�tx9PLT;)�2d�@A#�O��8f)�
Z3���É�}�j���b�&��uc��>���	_0��6�S�X5����#���53��i�.k�����@�M� q��'��	� ��@9>����ωv�=@$W�c&\ktM�	K��p�L�uCp��F�u?���D;f��;��,�ܴS�xj�fK�zs0����HL��E|b*�@��`r/N�<y����t&��DWH����6D�����ȝ)��ĕ+m�>!�����p<�E���
nTaJ�]����'�I}�*�l����=�|rU�Wg2Ԋ��S	��p��%V� ���#4��ـ)�y�-"���+��%��>D���꜔GX�h�ā��D��S�<D�TC�/�8��"��2x�^��m8D�P�g��p�4C2@_~�YY�"D��%e�� ��Š2m�9 �����&D���B&\��J�j�
"�*C�+D�p���%C��0
ԂP
dn@�Q�'D���1F���8|x0��9k�"��!�9D����ړV7~A����`�>�
��+D�X�D҃G
J�&��>Խ���)D����F:-��ys�ƵhR��2�$D�,ؖD��~\tl��
�b.X{@7D�l�tR�*����7E�yB�&D���CNw|� ¡��A�F��uN!D� ����[�f:Q �Xx��A�%D����0
(��-P�d.���0"D�,�d���L�j�KT��*H��y1� D��y�EMP�0���5Ut�hr*O���ANG+w�e�PI�X$�g"OR��eD(<h(:Q�KR���"O`5�v�*qr)��&*7T��;d"O�I��e����,�`Ҹ"OtE�T��a����3L�>��g"O��2� ã���8c�3����"O�<�5�ݾ(!�A.�	n�\II"OMc�T�L��A�g�Nl�"O8Đ��k	� ��f(hX�xۖ"OR=�!A�~8�1��l�-C'@�"3"OP��}��

~�&�؁"Op1��ժ_�`�(Bi�
�^@�"O.��tޏ<��m���30�*�!"O0����>F|�u�5,��	���"�"O� �t",ʶ��d� �0�AP"O��h�S���1�Q.�o璸�`"O)[� C6����.�_��A��"O��9U���
�9���ؤ \�"O�%p�7o�(8�m�5hY>1"O�9��,�b����J�S6V���"O~����(A ���ʀ"8��s"O$��V�wgT J��Pb^ʼ�r"O�(�W�7,�t ���w_L���"O� � �!��("��`1�`	�"O�U
�<�`�!34�Ę9�"OD%���F#W��{��Cr�P�"O��+�դYuB�j�o�ss")Q�"O�U0�']�(A��;aZtQ"O�0���kF���� D3V(9%"O6=�`�F7n���\)\�P��"Ori�需�r�H�hЏ-&z�B"O��w�+�r]�qLN�P�` "O"t�#��s0�����ɡ9�j���"O���V� j��j��2��H��"O,HҐM_�� �.��]u�Y"O��1�Z��0�glY+,�
� "O<��aƥ{��4KT�~���{F"OHh覈�!o���7�>�­�v"O��w�]�{jj��ٓXH2���"O��	�_�T D5��@=M�т$"O�����B3C� 0K�%"ؠ"O�A#�$jF�aj���;0��q"Oʸ���W�A�lP+�)���A{�"O����l� iYЩsX7{��Y"O�yrb,�%M�X,��˪	A$���"O��DF	���X���IG�0��"O0I�,��s|݊@:9ح��"O��0*A�8���p� B�!j��R"O̛jD��x��(\�S|l`�"O`Փ�cD<QH69P�'�i�(�"O��g��Mn����N�DB=ѕ"O�%����=3�+���6(����"O�1��\#MFT�X�۞i�`��!"OB�	���0���$�N͠���"O���CDȃL,����4���1�"OR�p ��Z��i���?w��3�"O.K`�A�4�Z7�_�6d�ʤ"O:��� 
g�V���dg(��"O��[tf��_Ze)�����~�ɶ"O�%�D�
�b6�|Z! �9�V�J"Oꕚ�ϗ�Yq:Tг�آD��"O�-q�l̵Yl ���H��_Âd$"O��0�k�'u,�:�AΣ�V���"OV�B@����ip������
"O��hpݩ�����`�.���BE"O`����k��L�!_,�vX��"O��!a!��YX@�_2��a��"OB�y��]W�9v'����g"O4Xs����@��!�Ж��=3�"OZrTi <z�x8*/���F"O�	
���"P�r����CA�W�<�7A�R�F`�0�6�
A�)�z�<���! ���3(� ܀�a�ML�<�c��;L���@E]��*�s�K�<1��C(:v������_���{�h�Y�<y3l��b�Wq���S���]�<�-�N7���A�&$mKb��M�<Y��B83pb�!�Di�Ё
�ËJ�<� ��GIʏ5�yh��Ͼ3���"OL�˱�(Z���[4O���jHy�"O�y�gl@/ �|!���}ͺe5"O��7%�TfI���Ko��	ч"O��!gȚ�1
�Z����w"O��í���� &��G���X�"O�h���W1)0��x���r���j�"O%c�N��LC�P�l�=4���I�"Ou����1o�T˄d �5�-�"O��yA��	'������%p8&�۳"O6�)���1��Q�c,!5z�S"O|J4�H
�qI&��iV��)%"O���d
� ����S�ǟH�Lē�"O���w�M}�l�
�@ �&��"O^��V�E(<<D�v-̜@�^5B"OJq\6
��3���,ƈQ""O�����B$7��E:D��f+H��"Ol�H�J�	x�%�$c�3�!�"O����-�:���C"-�%U���"O(��񣄜q!P��3��X�t��"O�Y�EgB2��c���M�QbT"O} T+N%Z��p�
#�r�"OfmX�,%_&X�5G-b/؍t"Of��U�J?v��� ��ߎ_��"D"ON��Ť@��,�`'�Z�)��)d"O��RFA�*T��j� *��#�"O� ��)Q5nj`Z�TF�3�"O&�h��E�w7j�Q�a�.=��z�"OJ��_e���xV+�-�0�w)�o�<��լ�$iۑ&�p9i��_�<y��y������@[(4i�#�q�<�!�.�j ��.��
�F)VJ�Z�<+R�$*$���
8ۀ}��m�<1C��D�pm#nb0��a�<�$�NۚD���{ |��EX�<1���=O�Iۡ��_�D�b�[�<�s댋N����2>�P�J�<��CكF�1J$���G'��U��A�<I��R��<aT�Џ<i\�;Ǐ�<a�a�7��a��'Uv%(��m�<I�e��r�ܸ��#�~��2�Fm�<���T_�Щ;�b��R�h��Ԭj�<q.�!.=Nݙ��ȫ'�Աu��B�<�A�\k�n�CC���4,���`�~�<��֏oO�h���	XȍHg(Ss�<����"����wd_����ѓ��Q�<Qu+�	9vv��BmSRbHa�H�v�<�C������P'ND����U�<Y�ʐ�XCj@ 1��
�\�rd��L�<a ��!��l���!�Z�Zu�K�<q��8N)NI�"/�\�ږ��X�<!#�9��(�Z\(�f��Y�<yf�
�y,n��֯�&T�H�lZ�<���	\�Ԩ���G����N�<	�o��!�h��ŌY�Q��8�|�<�H1M\�:�"��U�AL!��+Q�da�ԡG����@Ө^�!��T�a��)��P���8�h	�h!�$[�0��H�����^�J�ח]�!���'(�Zł��E��	TD��8!�ԧWuР��*� +Y����;7�!�[�g���JE�4<���(Ԙ;�!�$�<3���x l��'#�x��'ʻ*�!��O�D�G��Т���NR0��
��� h4
3)ǑW8p����.�&9�"O�첥̉B2��'�U;S*,�8"OT C*ƥNn������<���"Oj "�jI�*�i��6�T՚s"O�M[aeF�}M��y�j��7 lXK�"O��b⑑/�F}pa@�/%(8�"O�b��<xjjm�CK?/n�)"O�����3�q��)+lqr�"ON���32��I���L��h0"O���㉌�S��5`$�Y�]WD�[p"O�"p"U�i�b<� DAWz��"O������d'J18��N�p�t%��"OvM�0�ֆ?���B�[�{��HH�"O(Q볡Q��e�lQ�ew~�	�"OP�w�H��]pWD��.��P�`"O�LJ5LZ69� )��Q�+:�Q�"Oƨۗ&��J��|Y�L�9j)��@"O�M��G[Z pP��\>��J�"OT�(���(2��i��*C
b� �F"O��1dD�
�:XP�/��|�4��"O�]�uhˈQsz$��m�{l�$��"O2T��ƚOX�*���=�n�p�"OD鈡��7A�BU�M)q몐�"Oִ�!�7d�8M��>M���G"O��F)��qT�( GE	Y,f<�B"O��I'�͏`�h� V$ܩ*VU�"O�PRW�X�Y�r8���7�.e �"O�)��D��0��:o�2��V"O��bJM���a��d6g3ڼ�"O�y��%�x����3�k��f"O2\Iҧ��5 �"M u%�DD"O"�颩��Ni�z C�$!���"O�����K���x�g�ȾS%U��'�a�l�4=�Dh91�			�.�*�'mF�+���?�[��t�
�'�l��P.G sܘt .X{�0�J�'��e��e{�	'�?qfa�	�'o��J�!4t�jV�^�n����'�V�%��H�ĥ���^�����'�ܸ6����݈2�ƀVDu��'��k��,��U��̙�t��]�
�'�H)��M��2�5%̑�i1
���'^���Ru�r%[���)Ad��ȓw6 �Q�Ð�\z��e+R�Q�Pu�ȓW�ʈ��H1���
�F��<��ȓ]V���5n�(\���Hs	�*z���ȓ<,\h8a�["��^Gt�ȓHhu�UL�-���1k��9P��ȓ*��q���m�@i �2V�̇ȓ2��0T���i�F���!m&9��95D�slS�@�\XX1�	q�,x��:|�dJA�(}/0i �g�A�.��ȓ�~5���a�p��@��'��ȓG���!Qs�q�1!ĝmST�ȓJ`1�g"��s9��{��I�����|���L��c�n��BD�ȓ����P�ek�.D
�لȓI�zK��<h!+b��ڨ��cJ ��ܦI{�@�i߸L�,��ȓW�t��ԍ�;%�Q���Z.G�썆��rز%'O�I?��" «M`)�ȓ�8p��$�J���p _�g�TІȓAE���h9�v�C��Z�Fn�%�ȓ1_��HA�2XP03�*�T��8��S�? ��PUj"#F��1A�/f6���"Ofr�BM1V]�y
��!��a��"O�E7�\�{���%o���L��"O������#wR  k�/!D{R��"O$��V��l�6��4�7���A"O� !ul����-�"}�.��"OH�SQ�!t�-�f��<2���AC"O�� �a��1T� ��M�8y��Iq�"O� �	N9^������� �P"Ox�`��S��MralŪV�U��"O\�Ig�s ��Fj�&�Rp��"O^���E�M�z���G� 	��`"O:	��ڼ˄ �$S����u"On) '� &�̤J��k�N�8"Ofm+�`�'~��v����G"O��� �ɁH$�ЧL�	`&�2f"O~}2��C�h	`�ˑ�߱r�f|kr"O4�QS܂,1֌a3�@��@b�"Oؒ�@�t0����A�a��I "OZ5(r�����6�͵,�`"�"O
h	�)K<��Q�t˔���Q�"O��0�`S�h	���Q��"O2�r�͔ ��5c݁?�H9�"O���s��$����"O�?�$$�"OF��Qe��p�P�aJ��,���"O�H�'X�C:	T/����"O�����y�ء�'�6|��Q��"Od��  ��}10c����<!C"O]��*پ0�� #�J ��+""O\5�Se߱��Y௚����б"Opّ�,�^W\�I��D� ��t��"O������Q���A�� �,IRP"O���)�C� ��E��&�� �"O�t���ҔZ�j� �)[o�"5�e"O:���_-/��ǀ5��R�"O�-�6$M#f'�m9��ż�D(�1"On�x	P#P�%2�jM�$d�y�"O��Y�������0%�x��"O4ih��$�Z(9�ߖx�N�P""OѪ�%*�.��S�\�D9 �"O(�bE0/E|&��&�([#"O4m��GF�<9�	@nZ)z��"O.����H�R��x���'0�acu"O"-����_��!��M���J�"O�8��o�*)��5��
?��7"O�l�@eT������:�:]�#"O�@�CZ2O"�ȳ"�!D�����"Op�@Gé&N��cp!��LXhq��"O�A��҈wOK	7]+#���y£ޠz���u�W�~�f��Bb��y"�PJ�THbV�u�1#���yb-\�4���2�承s�.�"D���y"I\l0���1XȂ�����y�I�.�f�WF��R��̹ �H�y���cVh��c���8�Q1���y�N�Yn�%��ʃ�D���҆�y�GF��8T��D����g@��y��ׂ~�
�$/Xޕ3�ݣ�y���,B ����&n� ��Ό4�yRlL�
���jD-P�	�ȉ�(��yR	�>�
(�-TK9R��V�Z�y���'.v���i�py� q�
1�y�J�D���@WeRX���Ä��y҆���D�X���_��5�F�%�y
� x�"ɞ<�~��2�(v�P��"Ox��O�j����Q�k�@9�D"O�m@��U��1'��4����"O� �s�ú��C ɐ-(^Eh�"O�Q��
t �a�2&O��4"O�}k��蛔 W5<�a��"OI�󃔔=�I�T+SJ�P��"O�	���Q�ak�,F,p5A�"O����9��ó�Ug���#t"O�c��t�R�e
ߔHl�QT"O�l�GI�)KĊ�����A��80"O\�h⥂NxZ�ࡏ؏B`��"O�t���u��9ǮS��\be"Ox!��6jƬ�h��Д"�d
"O�Hs�` g@(P�5J�./�����[�{�a[/V%hE�����72�/�ZP���7K'�������y�E�;��O?���S�9�� �ՍP=A/@�Sf�	_a:��O\�J���}��O�Z�q�
)ϔ�	C(�@5F�o�8M�f��"1�Nm���Tb&U�v��$h�a��
�[�.7����G à^�2��*]��Xx�ޯz2�U	�(�0|��Vp� 1j�H�3сͦ�M�� �@�X$Uǌ����F�j>=ɔ1 0���ԩo�U�p����NC�H���f�'&j�|�����c�S+L�b�D�-x�Vi��jJ�6�2��$��vJf܊7H�֦�s�Q>�#���A������[Έ�ѨV�b��X	dN�d�����hc?i���ئ�M s���B�L.�')m;��	 ��,UL}�����a�		�3tĂ���L�@d8��t1�a�8�8=��$Et�[	�'?��Y����7��w@Q?��$�S�5y>�yk k�q� �B�O��ӝv`b��$؞X�r�0��]�o�(�aV�`N��g�ԴC�UE>U��)Q�e
`D�Vk���Ġ�_ܝ5�yӎ̨�J��p����Ms'�!?���3�
N��d��,H5SR��O�����9�)擫H��Q�.i�p�����#�.B�I),��;��.#en������B䉨<���3杤l�2�ҡ�؄wf�B�Pܜ`�����i�y&�vJnC�	K���t�@0q��Z�-S
B�	6'0��x���;���:@g��^�C�	�'�D�:���>dv~T����3.8B�I�{ܢQ�TT
1U�D���	%mB䉃7�`EQ'�,,������a��B�ɷY���ŭ��k���{�cۃ5��B�I���pH��Ym�� DM��$N�B䉥�4��n�1����QhX�X�jB�I�6�ؠ6؂^oxe���TNQ&C�ɪn`0����Y�Jr�ݨ&���*��B��, �J,Z��N	sL�Q��I7$��B䉬 ����D�� ���Re��L�C�	�^��8�vJ�}�����x�B�I�.شY d�ۜS�D؉�¬$�B��.���y0$�2
�"�`��R6�B�I�W,):be�d������fI�B�c��c�ZW�ങ��KTҶB��"��,���c5щt�G{�>B�	f��b�R���L��,/"B�	�_:ᘅ&�$B�@;e��3�4B�	?4����Hq:z꧊X.=b"B�
 �K+F�b�V|�,��TB�	D�з"�K�xL��#�+�:B��ZW���'��JK�(
 J
���'�����P`
X�*���&��-R�'|d�D
IA���q��5(�	�'Hb�ʤ,_�[�`bb���ڜc�'��D�cR���kN��X��'5d%jsIݳ9��Ic�a1�X�'6"|��CS=l�	�B.^, ��'r�u��E�q�Rp��o�8��y
��� �i���4֔AV��%�|Ac"O��7(� lJTP�Nʦ;���w"O>�A'҈/F<e{��K��:�"O�[ËV��6�4V���"O��S�Z�\��$�/��t�ȡ�"O`l��f�
��1qM[��d�#"OmR�'ǃK���2��\�a����"Oj�{�N�$�5@�F�� �"�"O�H�Q
�};ڽ�/C���{P"Oj9
�.	�pH���(kG.x"�"O���N�uӸw'�|����"O��ã�zά��ܳC-�l� "O����D�:#p4BHۄ�骖"O���k��e6�`�h��{�pa"Oږ`EDyn-9�i�,����"OR�a����̅;1('�&�9�'�6�nڷi�Y�Xmް<��'ǆ�qj��~x�"�nw���'+�M�L@�� |qWn��.���)�'���K��il���VG.Q y��'R�A�qO� _���*O$4�&E�
�'A�@�Ӂ�h����̍W�Tl��'Er���N�k�	��F=<�T��'�p`���\�lB�P�k��2�y��_�3f� (���i���N��y�-]��6(Ʋe���i����y�=4z9� �̴O�P�EO��yr%�:�\@"7a�2p���Ǝ	
�yr���Ա�v�I0A Pfe��y�玉8�!����%p��)�%�y�A�9��eA���S�@!�)\ �y�b�2a��8Ic�]$DKlk�ʁ��y�KÔ#Ԛ=�ЬP�@��Yh��	���'�{r.��`��#pOW&L���'
��yBb��C�aA�('T��);��R)�yr��~�ap-ʨ6�E�1K3�yR�ƿQ��\�G�Z29�а��*@;�y��S�$�:����
;��@�h5D���٣bK�\�Q@ld��I�
)D�@�^�,�҈+䩁n�v��S�'D��6	Q�7(@����ʚ]�N�Sa� D�L�Q�W Yn��A*��$�@��<D��B���:"U{$J[�n������6D����%��p�AZ�l��-P��5D���0/ޗ)o�E�K�&t<y�&D�ȱ��=Ka2H�����T�}��.%D��R"���Ԍ�0GѺJ+	�G�"D���J�yt��g,N���qӭ!D�t�cN�jh��zg�1Dv �he	*D���l�Iq$�������A�3D��8HF?N�Ľ�q͝�/�����3D��KU#��V~�9�%���=�����5D� ��*�>b���[��R*�D�d�8D��Ӵ�F=�!���E9�`TX4H8D���jAyJ�1�5��)���8�o5D���aԉ4e��r��"�����#5D��1�J��2�*%��"`��8s�2D��`e�l"(��T��`�@�/D���T'ѥ<��� C�"�
�y'�-D�,#��ٴP�#kG���U��N6D���D�:nL�ᪧ'�!����4. D�H@�Ix��#���8vyp��+D���ū�&���㖈]8�b�Q��,D� i�@@�H|�1@uf �t�+D�� ��� �G
'� q� ]��!`"OH�0ƉR�
�΅���W�*WXY��"O	`P�K�슄�`���[q %�D"O*U��Ri.���u�J�U�h�"O`j��G��i����E�"O��s��ͺj��(x5'1sT���"O��;F��a_h<jWf��Q�8�"OPiXr��YܔU�d+]�8Π2"OZ�
�ʄ.��l�4!]#.��ۗ"O�x��%��s"G���!3�"O����I�&t��L:_����#D����E�
��4 �Й#�"D�`x�H��'XI��0/�J��1� D�p����c�*1���B�	%H��   D���1�I*Cհm�&�A}։�AA0D���qB��c���A��D/�U �G+D�|�4�Ş1a�MY� �,-(��c)D�X�7`D� Wڡ�7�BEQ��8ԥ*D���-�Z��L7mذ5�b�%D�4R�YN�J@�Ͼ@���%c'D����'
�O"(�A#��?��s&
"D�̐*��d�3��$�����!D��e'йnĬ|k�a��rj���D?D���#�>��}�pb��{�X2g:D��ڑA�U.L�M�#Lxpq��8D��0�#�y<&�z@h>{j��u�$D�8h�� T��٪s�R~�&�P��.D��3��\�XLT��u�E7<*6u g9D�x�Ċ�!�h�X1�A0Pͱ��,D�ԂF��,�����*A)\4��P��*D��
%�Y�Ɣ���A!,�J�)D��PD(ߣ
HbD��{�j�[5�&D�@���zk$�X�C3	�TБ�� D�ЀíL>?�Ay�G-Q0:��3�<D�\���Ȕ-����e��k�HC9D����E�Y�*a �ʜ]�p��a7D���cJ�"4�1	�=,��}�6b D���G#-A���m�;=���=D�4�dO%�f�gcL,J�vəW�<D�d D5fl� ����,(^����-D�0)��:W�����[���D�>D�4��5����^�c��� u�:D�����[��<�%�Y'<��,�@�2D�T��B�}V�i���B�c������0D�`�W�Y��,�+AD��f�r�PeB#D��9�l�]���!��B(7 b��$D��)6��e��h��_�
�;�+5D��P�k��B�n��S/�͑vK7D��qG�M�b�0��^�N1�%P"#D��R�D��H+G��.+���ի D�����IXԌ��&T8d��}��b*D�T�f"�E,,��i�k��P��4D�j!˪B�,Pb�NIjTy�2D�d�%@&=J)k�͞�{����-T�	CKUb�ݡ��G���3"O�a���}�&܀�G@�`$T��"O�y23��-vyr�2W�n�A�"O
�(V�χ"�,Uj�ʪ�H�C7"O\̡�J�e�¹iWCs���"OH,�`IWA% Ô�.�Z3�"Ot��c�S�L�<й���TmrU!u"O�Rq(">"�{�+^RL�)�"Oɑ��E�F����qa��M62�`"O큅 �����cK����bf"O� �P;�L��.f�ԲaBƼ}���"OJ]ر����t8_��5��"O\S�\8yW���%�Z�M*��"O� C_ F��9�\8D��y�"O"��e��Mn�=P����y�C"Of1��Oٖ-b�\��m�B �!�D͊��L�%L���0Հ�C��Y�!��O1HEZ�ȇ{�Hh Cx�!��OU|�"�)<MQ�wA!�$�	i��l��f�G8h��o2Q!�Y;0��ْ�	(@	sv�ҚH_!�$F���A%'a� ӐW� ^!�@	��Y7� w���$�_!�d��D�����@Д.m�=JW��!��"��+��;sj�|� `��@_!�$�z��҄�E�	�cB _�Z�!�ė;X@�x�C����;ņ�U�!���VCJ��.�?*©����.�!�d�D�<��Fm�a�S*#�!�Ě�|@�a�o��Kj��f�R�Y'!�7R�R��4fŹ}�*p2�@F}!��.Z��(��<E�%�Э1q�!�S<]���YF��e��p�
N��!�K7��P���%�����b~!�d�u����0�Ly���Ɍf!���P� XKa��'��%�O��"�!�$Ԡ=�H����%���5$��jq!�$	a-<!��M^�8�IP4�7UU!�DL?o-����6�0��W�M(;�!�d�XB�m���V?�($�B	h�!��ʭ.=T��<WL����R92�!�d�=u��ys*��(�\��g�pb!�$C�T�ʙP�@�pi�. U!��!-D�0V��&Z�ޜ�� =J!�" �$a�4L�9bv��:!�DG�&[�E!7`:�Э�&��!�؟}#XT	���u�ܱSR�փt�!�d�7yɴ$�Rf�p�ڙ���,}n!�'f���v��:Bͳ��":a!���&��MЋD?r7�9�u�?P=!�؈9x�+c�Ң����բa1!�Ğ�B�L)Xtl�.,����CI!�Z�V
�12�͗�e8&���E��s�!�$�(p���QЧٸz1��DĒ�V�ax��'�L�V ��i�������lA�K�Z �������G����?9�q9�Mx��?�K���[teь!�H�%��)��H�U�
a���;5�܍;4N�!��9`�rd���e�'���[6#Q�+D�y�����W�r[c�^�N� P�CI����)�<)���^�'�������-������	�i{'�Y5�ܼ�1௟���러�?�O!�Ix8h �D(t�l�GKq�B�Ƀ���T'XO)t�f�R�=f�R�#Z��M�)O@I��������͟`�O�����i�5v�Զb�h�kqA�:DE0���O���T�/x�Q��sF6�x�'�b�Hb�Ѡ+{F�'(Mf�DV5�r�P����e�'��R�_��ڵ��Ť9ZP���7'����RZ>A2�G�2W�N�p��/q��q�(�d\�=��'�����n��V��
"��" �wN<kG��O���\qdI��s�� ��!i��X���ͦ	�ߴ��=�`�P�F؀_0p��!��Y;�g�����O���AzJ �r��O�D�OP��w2Yf��F3ʄ�K��E�l��$_��M��H�g��IPf���;|�`�Od���:R�<L�l�5�2�W��z����/|�<�ebV)��bR"�..��5)a�[L��I?E�a��yw�\P&��W��*I���jݸg6Dl���D�U������?��4O��0��Y��,���ʉ$��u�4�'�RY���	v�gy��]�G�*(y뎠F��!hQ$����	��Mk`�i��'T���O��I�2�,�@�
٭�L=��K�4i�����D��X���?����?�w��J���O:��^�Rڑ�b�ɐE�����H����f"�*:�P�M�R8J	�7KQ�Z&
5�a�	&%b�ٰ❧N��!��-�Y�P��BE�*��KNڹ�̍��gĩJ� رg09� l��%V)�>�d�̀Y�#������+شf�n�'��'��OnI+0���,Xpe��o�/1�d�S��LD{��)�*�l{�`X&@��S͛�:�"��I��M���U��oo���'J�|)�i���i31{�n�v���@��$Zj6ɫ7��O���I5h�d�O:�D�B�TTQSA�=J"�MʤEު'����Z�Xc�H� ��-�x
�-��@!���ITb"����LX��*��,X�٠=��4 ��~L"����O㚩� �ɻ����ӦM��'��є��D�;C�<u&T��{2�'5��p1���h���1�Zh;`M�@�'p#?��Evʴșu;�Ĳa-\Q���(Q�iRd�X�R1��d}"�'���ON�mbA�iΈ�T�LS�����"�.XS� ���O��̎,^�iv�՘9�L4	̄c�X�Ң��o=�V��Wg�,�<i���8M��'�4kc
 XV��d���,��<7-B0����O��Q��LQ�e���9���F≰	:����¦��4�?����)у�,e�e��9��J$��'��'����?�d��}��%�	c,(7jV�u��x�eu�(Uo�@�ɍIzٰa���a3�C�"����͟�&��D~"遙 ,  ��     }  �    �'  �1  s8  �>  E  KK  �Q  �W  ^  Td  �j  �p  w  `}  ��  ��  #�  f�  ��  ��  \�  ��  ޸  j�  ��  ��  /�  q�  ��  ,�  o�  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6�F{��'O��V���&�;�+0:��x	�'%��"J�[�]�R�K2r��"
�'Oe#W烹�R}aC��z��
�'��;��7�������L	�'�:<*b&K"4����M����9	�'نx!c̓>�D �,ݻ2zX�R�'��@ �F�9<�m�7I�"+�a�'ր����>��Y�
�%&���'��0��3L�r5��M/� HJ�'U����J08fx����I$p:<����O*b�X�S�!��G ��s��PDd�o,TC�IlߢE���5Tvf�����}�LC�&�L[f�R%'�Y+$�@�	�2C�I*zX�ic���%|���g��d�ʓS�v�<!����
/����县)�B�ٲ�ITl!�d	�N�(4$Q?a*FL{��[6M1O ���_�V�� ���C�!ږ͒?!�ͭ~��M ��<
ݪ��5lN�!�D[�$��BAĚ�0e6���Z�q�џpG��ч	�fh�ǈ2���
-�y"�M�s*ZT[�IU�sԢ[��D��Φ�?�g�Nj�yc�Q�����QÏ/u>����-?BM�X�A�!Y0I¸��u�Δ�䓘0>�D/��>� ��E�=N�U�G��t�<��( F�qb�5 *,:�� q�<�B鐨>spU�Ў�i������Bi�<� �k�CՀH�)�.u�r�#u"Ox��^ƴ��񊓚mHX0�"O~�0��)[���#��0 ���"O��i&i	?f��t#��"9^����D3LOf}�լq��CC@��Bo��"O>8��%°�t�)u��]j��Ҷ"O�8BR��#`�(��lN�1�l�å"O.�ґ逜!�I��B̦H�Q�3"O����Ƀ]6`����5e6��?O��'iў��X��Q�W8|x��(%� {"O\|⥭�9DT���\$�8�"O%��iy�1�-�� ��S���I�����C0�!B8t���ӎ�MR!�$��Q4m26(߯�V�� �K	LP�{��	�Pt�!�"���>��a��I�A1!�G%R��p�Х$�l,z�M:W"��G{ʟ ��R:*P��x�I�	p�n�#'�'��I�YDT �刚:E7�(ڵ	�fB����kk*tH&�F=	�F-[���-�t��p�\8��,�f�t!�kY-a�"D�ȓ@�}���T3O���i�4Rs�G{B�NF�I�_�5���n&N�)�g�5^B�ɋZ{�uí��N�T��Ԙ��C�I�r�l@�C�:}���cCC�G�"C�I�
d0�a��	E&����rK�B�	�E�̍)�L6g�FqY��Sns�B�IM�.��TN�x3a��}�B䉇_^`p�1ֻq���p�E�#a^�B�I�q����l�jhr���_ �@C�	�D["����L�#Ǆըl��듎?!�)��),�� �KO:dQ��*�h��H�BC��_��t�ī�P,����
�{�8c�����'j�Tisn]1�	�gƼrh,��>��|���i6EQČ��3���ɗ꓋W�ā�'��Q U�0,��4��90,[ۓ��',Z���.H����$��70Ѽ��'l�4�e+]"
"���"$�&	��'
(p�ϋ�R��#��l�R`*�'6 �3�$�S�pB�B^4f���X�'֩·�+g����7�Y�Y��\�')�)҃f�=��Q{7��)UЮ���'�H��d�z\�#�#vth��'�b�Cq�ѷ)���í@>� ��'�����G�?|�H5���<�P�@�'�h�e�Ò%��ȫ�B���e�V"OL�Z��̆:���#�
IT6�"Oʜ�K��Z&�
&�R�Fd��"Ov=��۾7f�ECF��w�(r"O����CI7C���ɲsA�r"O8(f��4���0V�|4�p"O����'JD�Z��ڍV�q"O�QWL�ZX�C��W<7�j��"O4� R�[?d�t�+��> �2���"O6����8kx���n�F�6E0e"O�|#�N�0�n9�D�I�.�
�"O�$Xs㊑qԈ����1�N��"O�t����Un�va��/v��K�"Obm�5C���� ��V�z_��p"OD)�b��8��"fM=|N�r"O&�0����kj��Eʢd99 �"O�-�s
�{@v5c�/2��pG"O��G��5�v1��l
�o�I�"OJ���"�*Ǭ*(zĩ&"O&�Sԉ��S,��X���]ؕ"O� 8��GN:30(�m��x9�"OƉ[u��	X,�T�K�(	w80�"O���3+������[5dr4l��"On�hG�M0�j�2Ȋ�)%"O([�ׯI,Ќ"qG�0� �"O޼z�Ì)�D�D��4�"!C�"O* xt
L�w*P����"9��q�"O`�����.�v���Jh�� �"O��3��B�?}���vYHL	 "OH���1���['�O�e�e"O��;�(�����bHA�:u��"O^��2��w�P�jQS�[�(y�s"O�e�f��W"���A�=�ɱ�"O^�:���{MVTb*
0�H�2"O<��͇�x�p�jtnN7'42�"OJ0�b<=P����c�2N�D��E"O��(���!jf�J�C�)B�0�W"O S'�/��q��S�L�L �"O�Pq@I�7%��p
��T�B9҄"O�)�� E�b�d�`V�(3��4��"OH<�Ѯ����ՍB�h����"O�� �] I_�)8�FH�;���C�"O�YX&�#8kV �d��)�Q�"O�	�'C�E,��(��=#��W"O,�8��`�Ѻ�h�:)I�"O"��!��U������&��M��"O� 2S�ݸA����&�&����"Ob`ժ@5Jw�P�R��W�^��	�''�ѓvG�#U���&�79�<B	�'H�a�M��!�rȑ 9���C�'�����<�6ۢ��4aC��'^9!� OH9x�*ԅB
e��'�HH��Ƙ;`)s�h��fbr0��'ml��E��s�j���� R�ha��'�Z!� &�-$S�q� �4KX^l��'e��Z�nP^ZtX�F�@� �'�6�P'�3U���X���5�,�@	�'�V��3f�@r�vN�
z.�|Q�'r�y8t�I;,'�ă >�x��'Q��J�,�
N�m�E�@�e@PI�'he��	Ż ℉�8���'��i�d��f����$��!8�'dB�(_�odU�� �S��' �k`��(blY
�a�Qt���'(=����s<:4��㞣�PI�'��U���6Ĭ���ڑ ��
�'�F�`A��>�ɺ�Σ58�c
�'�d����2FX�4�c���'� dr�'5���蕨6R@(�V��/j�ޕk�'`}avO�8S}6x�e�R*v����
�'�2a"���0���6a�t�.�
�'�Mk�M� s�*�֠He�B`+	�'��s	M�k",�ŭL	5ܼ�	�'��Kw`�3A�S$nP�$�,��	�'������_����c@
Fk�H1
�'Q�P���[��,�A]�KH�B�'W��Qm�Z�@C[�|hh
�')P��^Rt��c�M
�(���G�<�1
ׂW�(A���
!v��(�G�Gg�< m��IPi�Q$�q�Jl���a�<���U7"��e�f��-Gm��+�LS�<��A�P���3��W \�峕�w�<��6������q��9�P��|�<y'/3��ui2�Z47�<��R�`�<� 6�SK_��%�6��v���"OZ��9g[�01f��E��%��"O��g���8xmiU͘�t�6"O���ld�R�K]�J���"ON+�z~D�P� �s�u�'���'�r�'_2�'X��'Y2�'��aꀋ�8	�9�cK��Ox����'��'�R�'���'#b�'L��'��Ժ���(����c�klTxJ��'���'���'���'���'uB�'�ڍ:$�;&����w��Uq���'-R�'�B�'���'��'{�w#�� �*��/���"V!RW�P�4�'�2�'�"�'4B�'�B�']��'߈���h �D�̑�vg؇hQ�����'�R�'lB�']b�'��'[�'��=PA��(��^�o������'*��'S��'{��'"��'�b�'$L�
"EB�~�����+;��E��'MR�'D��'g��'���'���'Cv�AAG�'�j(�4���f-�dc��'���'���'���'CR�''"�'�ʌ�t��Zy�+G�l(sA�'�B�'���'���'o��'��'���5$�%T��(���+sA
�B��'|��'�B�'K��'���'Kb�'r�|����
h��EË�;ud�X�V�'���'��'�r�'���'n��'�r��WM�?O)�I���	QN�Y��'�B�'���'���'�r&gӐ���O�ܑ�
���q
�%��8ty[W
�]y��'c�)�3?�"�ib�#tƗgV�� ԣ=O�!%���Ĉ�9�?�g?Aشfz]���&"��a@���f��ih�i���J�$�Pp�O�q��)�.sM��xO?�
����o�U�C,_/�,���?�	�'��>Ak2���.�r%�mw��YwE��i��6�^�1O��?aH���� ��L� �QK
`�VD�VK�.!��i(�Ķ<%?�!gNZzr��3��и�1Q����E�2`�ɋK1^I"hV�"j��E{�OB[+_~|�"�]D��H���y�W��&�p��4 �)�<IGI��o�r��J�{�l���%�%��'8�ʓ�?��4�y�W��C0-��,d~I�p���iTtX�72?I��޺�1���d�'9�e��o�$�?��@�q�V=��8Q�Tъ3���D�<��S��~��� 1H�!�#[�N���p���<a�itv4��OXymZK��|R�Ƀ��TF0A���x�&W?���M���J�h��CM~¨��Z޼H�LSS>���͝�J$5����4.�Q�F"]!6�8}[�'iJU��i�g�I�4�;q%�F�$1Q�¾VHC�H��:�ń-L0�Ɵ'5M���DT�xH�F�Y~�	�e�G�VI*$��>X��p$Ě-!e�|��W.w(��P6\8R�<h��bA�u��D�B_g5B�M�31>.���X4C@pԑ�W.~�l��"`D�]��SņE�uJ<�(��F���q`�=	.���Ü�{v��7"��07-�Oz�D�ON���f~��[-���$Î�*����������O�9�q,.���?OrQ�e����L�%���0�� &�i ��l{�L��O����f`'��S9��Jd�@-+샠+;T��lZ�t8�p�?��g̓�?��D�-��C���
���$t����'�2�'�f��0�4�r��O�H(dJL'���SȟoOB|�ŤS覥������I�Ұh
������O����O�t*f!R�_���S੕�8TQp �Q�ɉl"U�J<���?)J>�1 ��p� &	��y�b�9���m���`3�e�ҟ��	֟���🔕OY�O6,w�󷫌0b��ez76Ig"���/��O���Ot�O��WnB�ر&�'������;X�Z�*���O���O|�y���#�:�n���Gǜ+��L�I�&x��ęx�'m�'V�'��	�Oh�P���;Wf�	qÑ�� �+�Q������,�	Qy"	;�h����6�B�d��M���\AԼ2�ۦ������'���ɿ1jhc>7[��!"Ņ|� \�j�W}���'��_����fƗ��'�?���S�­�#,ʤF�����0+���)b�x��'W"�$N{��'�ҕ~���^#VY2Kc柵E*�"u�Dצ����8IŮ/�MK�U?a���?	�O�� �b�P, JP�T�d�B�!U���I5=
, �?A�g�W��x�c] U�qq5,T�9Ҿ7-Q='��o�ӟ����T������|�2%ľ+��p�H
�m+�d�)	83ۛ��p�b�'5r�'U�TY>ՔOAy[��ϯpc�P)-�hZT�w���$�O,� 	~�(�S��>�7�V�U}����l�-,	�Ԁ�aVl��ܟȂ'H�l��?��'�F�"O�g��m�t�N�n�
�2�4�?���;���a���D�3$�{��--BU�����mb0]oZƟ���h��Ɵ��	���'ń8�b&546����x�H<�(�-�dOT�d�O���<Y��?�HͿK�~�*�[�0XL��KZ0Ed������$�O"���O˓wh9cg4�1���&'D��	ѯ��}I���Y�(�	؟���hy��'aR���h���6s��ܫ��R�RW,�z�A�&����?!���?�-OJ����We�S�:6�d���j�4���d0c\�9�4�?�����D�O2��˄)����|�d�6C�����șrk�̓�Kν.כ6�'�B^��3ꚛ��'�?����d%�U�ġ�	Y"���"th����'���'W�yi��'p�O��\� �Hh%.�+`Sɑƣ
;7�9���xR�H�& ���n8O���A�m��������8I�"O1�L�"N�X"I��*����� h�
lj$�>h�IH�Ad{6��7.ū\��c�K��>.�q w�t��}27�+*J]��m�64�ẕ�c�:I����a$� PΞ��+�1-�
�r���$o�< �*,q`ԴPɖeӗ� �x$J0��n]�<����S�G��4aD"��D��p;��Oz���OB��ƺ���?�g���xqB�( �l�J�M�H?!U]�V��x��Y�X/����8x�%K��97%4H��݈gVҡ�R^��2b���=Q�ӟC��X���'ļ��hX64������v�|��'�Q��>��f�,��O��Ĺ<ɗ@�T)lL���T������H�<a�@P�:����\%Ꝩ�遭i�x�Ov�	�=،�pشt^���AB2t*<��aBJA�~@��?���?�CLK'�?�����TƇ����{��5�0��e��9�ȱȃ���D:B�"`�'�ĐA%�0'����k���%�K�N#^q:��?��{�'�?!��Q����q���P��^�Z��TYL>q��?ɌʟLYeHP�+��x�4�Vhj1	f"O���xQ|�X��?t�EhD3O\�'�剏��d�ܴ�?�����	X�R=B�IJ1 N�i:�J�^�؄���O��d�O����� !��oFh}BT>��\s��Akt*J,Ǹ�p��9ʓ^�L����@��Bw��>�\�p�Ȕ�O�!`d�Q�!.�J��c~���9�hB�q�I��M�֝���'Z%�B�� ����Y"`(���E�'h�O?�	�D��i���]h$т�j�@�'���,yٴA9���'^8� E�+,�ʡ s�	&܎}8�'�Ћ���>)����Iݦ&m����O|��Qrf����ƨ+F5�����2պ�	�ۧO�+�皸]�E�p�UU�t��wj���݉y� 5�ǤΡ�bXɥ��5vU-���\�T84���LΈeТ}�ݳI�dł�	P� b�um��$�:=�4M��ش>��)�i���{��3�JA�<}���@�M!0�ȓ>X�2$���[�(�HQfمA'��Ex�;ғA�I�#��ĺB��'��� 0��V����䟌;�+� 2g�a�	��D�����XwTR�']҄@ŁDsVƝ3��Y(��5�a�� ��)mR��)��	�D1���y��� ��A2���:6����2�N7=6m��H��ܒ��ІP9�݉5џj�C�����Ov��gi�	T
h��U	V��e�
ft���T
�����-a�t�'{rW���MϮ��ٓ*d�T���!D� �!`G @�@�(��,7Z���t�9ғ0�� ����ӼS���"՘ !�>a��x1(�`�<1E.�"*a�}ש�:���6�x�<y���/X��j3c��c���P4PI�<�G*Фq�	+�)
b�%�f��E�<1'o[�w�њ5	_�io���E��j�<�t��J9��H'���O\&H2�%�g�<y��I>��C`雀	���I.�z�<��:>�lQ�c�50�]��g�L�<y�KH�hʙP	�2'jJH�Ǥ�M�<�)@�F#`���cY57�zEADk�F�<���#
��ј�A�%@��� �HA�<y4i�<fșR�!��(�G|�<1��
�^� ��p瘑~��*5JUx�<Qi�=$H��B �r���bHJs�<�ʴUMi��KB�f7ȽRĥ�p�<����3��I� "G�H:�@Gl�<9��=��ŏCX��)��f�<9kF<%8��#�܎ȡ9�n�_�<��#Ʌxì @�����"p��[�<�ݷIȐ �8=( �'��W�<�s��94�PC����4��ii�V\�<Ѵ̈́A�8r�k�2r%��O\�<�[�#��yv�ڙ��5�P�<!��;M�tڳ�/>n��0� ]O�<�4oO��.�G�R(	 JH�<Y$C�,N�p�3$%]8jXP�h`CQF�<i��V�[�)Ȣ���R��1(AC�<鲩^�Ѫ�S��4e;��1�[�<�V@,;���F�5/�dx���A�<1���	2�Xd�T4u��uY�D�<�4I	�d�<1C�b��[I�uXA�<� ~�r �31�Ҹq��ʲ-dn�s�"O��;�	��R]>1j���H+W"OL���I0��c�cޗ&�(x�`"O�M�L�\�����K�؂%"OR����zw�=�š͈tB�`A�Onѹ'�)�)�'C�0�T8���	�C� *�8X�ȓ]� P!��3H*�D㒉�.��%�'Tɋ�-S��ؒ�Vug2��@��=G)�۷;�O��هEж\�(\�ЋZ���=����i��dc"O�����r�p��ɍQ�𬑦��0[y���7��g$t���F^-Ą���'��q��C䉧N��4
��B�&�P�*v)���y��d]�0ʬi�N���T�B|�B�ͻy1B(��R.Y ��{T��R�f5���9�B)��W29�:]#.O	 �Y�s��hyr�P�|�a�bA�-#`���D��(Op�@d�[#}>Fu��+d,�4�'^��5�˭�!�d�_�q��!0(łos21[��G&����' R-�2/�E{xe���"u"uz����扙�@���pt:��5,���cB�.d���k������h��Y�J({z,C�ɗ'Q�0��dϻH��c��CF|{M3/�v�8���?�g��0P�F��>(>L�r�V�Un�Y��,��.C��h������0W:غ�h߇%B�IDB"?�sAɎo�	�2��$�!�:ʓ2d ���d�(���'�j�����I'Np�!�A��~I�T� #\)R����Wl$u�Af�C�y�� �/�.>E�@�Uo?$��|2I��sC`��a�̴��glã��Ěd��hq��Ȧ��qb������p�����5���q��T,�yҧU�lK����F��V�����j�Z�ȶ,�)�u�=�OXV�	�����y�h �@�f����� ��I�օ��x�`� �x�Y -{W��*Q��17��0��O.��S���nllc2�/q�����DJ{n��է�!�����f�;�axr��~��	�QG$5��٪#)��=����Ŋ�R���$[� ��d���
�a߬)*��O8��
�W�!Θ��&m%M���qQ�6?��E�

^���-8a���1�!�i>)4�قs!Lq`��y
K�I�!��̣}�������u�V9�K5��=lZX�r�b�J�d/��ؑgت��w�8�i5��1|�ҧ@g!NX��'\8�k�\)yشd�Q�@��E�r ʕ�S�]�Af�Ԣ�yy�����D��59I<�㈜,+*Z�Q��>��oW�%�`����D�Ժ�2�ۍX�^���HB��d82�n�{}�j��j,�ۓP%�(Q���z�nL3'%՝"�H��'\pԑrk�Y�S���^1�h�(uMɥtp�ixd�ȝ2��	a�/C�VB��&4�t�[p%�[�4HVΞ�(��O�h���yQb�ۀ6���O���K�����D&^=0�{�&LE�����B89&LK�FR��GfȤ1_e���d�`E"a(<䆓O?7�ܙyW�eB�MU�Fz\e�B�Z⑟̹�$�.*�	5D�h�!s�icb#t/�.8�fE��&��T�3.v� 膉�/�$��	�c�,�'�������d_��!���Ͽ�|����v����`���O�� �킯XhC&#B-g�|}���$D�� 6��o����PȎXhp�PW,qӦ����OZ������*`O�MSS$a�u�i	s�0�둄޻B<Fu�L>�O���$�æ&����D����1l;h��~�P�I�R��ى9��8�����'�4ikF���}B��J�Go4	P��DKz�,��EG�6�=x�A�*��ᕒ_ʠ���#qH�@�c��8�^(�u��]!<���i��H�2͎�'oR�фoː9dF�Q!c�>y�"�<ۆ�#7
Y{$Y�b��s?��'����6�Ի�/�'�ԙ��C &o�B�I�<8ԓ��R���c�����3�S9*��'��$���IL7;�r����+�.�*S1�����\��&�q؟�2R,M�fB!�c� $�y����|ڌ2�'��$�&��8j7�H�!�qOL�H��=M���= j8���	�_v4�krk���S�I�&r�a��>~��� W�^�C^�Hz#LV�Kp�m�UdJݩp�{؞�� V��8�e� �}.��S�"+?9V�!v{\�$U6����K���U�9���6!����N7;iL�6a�I�0���,�ܸ ��,�2�{�bP�@�����ƝA��˖!SZ�S��Հrx��wC�M�Ve��tO��h���=LX��'ÐL��+�x���k�2w$�̓ J%��	$nH�#I�$
v�AgI=�r�P
f�W)0��b��$�+b�-�0<)!V�sv\�l��N�n��O�? 椲��آQr. �W���fSi^
+�,!��;u����-tͺGR�Y[
�sa�_�F��	�"3�*�ʞ�T�ó���wh��i �zZ�lq�%wx�J�жiu!���h�����:_o� �ԫP�d�݉��;������T>���G�vI������H� >h7�xa���B�	�Tȅs��� b?8P#&l����,0sF]wj"�5"B�H��R���'��'�@�2B�����4���I���	�Y�خO|���=T$`i��Vr��H;���)��0�E\���&�n�ث¦�2��@�L��j�4� @4�;�ؕXb�"������[��HX�AG��ڵɃ`�^�<&3-lP4�C$sc����e�c?i�h�����h�,�;��Ƽ~ͫ��P9"�yU"O�jb'�"�x�'�0s�(I�c"O�h���'#�Hm!��X�P�4@ "O��k��6�J��ж�xD!$"O��E*եpr�)��$Y�=Pa�"O�T���F)5���c��6�&L"�"OR�� fBVST��e�0:�t��"O�����=q˖E�t
�:���"Olq( �N~\��dI�,�I+"OP���j�)(L8L�SC�!-���"O���B��#*ڽ��@�L �"O��pN:`�K����8���"O�)�!̂_��x�T�	0W���14"Ox}s�ԕ9���0��X�UB��2�"O�� 烮[�$H��O�5>78%#"Op�%a�6� �k�h��^͉3"O����F����h�f��.�(���"O��ȳæ&�P��a
 5� `��"O��`�)ߙGXh R"�hƊ�sC"O�h��<(��V@Ԑ���E"On  ��$C
�Y�1�`}�I��"Oh,y�!�7�0��!�
>�d��"O�d���Cд�B�Ēn�8�3�"O�y�'O�� �(�BF5
=�McG"O���d�64k�HQ#�N�j �YCG"O6|��_7#*��7��@E���a"O�q��o�" S\�j�� �-|m`"O���֭m;HYuI "�i"Op�87O�nZ�z��
 �`��"O�(��j�)�n;ǮK�%d���"O�5��%��h!�᎒,UY�"O�<bD+�r����V��%�e"O|h;T�D y�$8
B##n�}��"O΍+� �L.⡊���4"�{�"O�Md���y;�0� �X[�Ћp"O��+��A�NӴ�)fOڷ�*�y�"OZ�iGbT�E*~)��M��>Ԟ4��"Ov�0E�E�x���qǪ�� �90"OH��OE �+�� �Gj*��DlS5�y2I�.s�8# '�=�L�XW$�y�o2d���g͏�4R����`R��yb�[�o�,Ub��^�\�X�2�[��y�L�6��3�DJ�#�p�)��ѧ�y�-Z�L@��I ��*dȩSTA��y�L��[BZUQE��*��`�#���y�(����A�.�(�# ��y�(рN�4+#���@�7���yRBʌF(�A��I5���  �y�D'����H�$dR[♤�yr.χk¦�����F�u�5���y2/ݢ*�� �נ2?�&�6� �yr�U�=Ur	�2�N D���h���y��V"0��a�FE#>����āԹ�y
� f���胗a`�bB"Z���*O���q)˔�v0)c��Ұ��'�f�b�HI�#i�2�k��!�l��
�'�p���=eLY1�!��!���)�'$�ϭrѓ�K��$_���'�v�	5�֞%�����h#��!�
�'z����5~�
D��T!	�ؒ	�'�@���$Z���g&��
�'nP���'x�,"���	}�Z	0�'�*�r1�	�@@�%�!q p�'�^����^�P���(B�SS�2`�	�'�r8��Ĝ�\��1�9Gf�`p	�'�,��D�X�c�(��e��6�D���'�����&ab��$ǰ3@��'���D`$8�ȔP/�!�f��'�Vt�#�J�ݜ-��(�N�,q8�'��	!�V��@���O3Vl�0�'�x}��ZH:�!p��*q�@��'u~� ahŰÄ!'*��Vp�u�	�'t��w�͵6*b�:֪ANm�I0	�'H���q@X3M�6@{FK�� 9��'�H	��B�d��#��H�^��
�'���%-ޔ�t�T�םS((�	�'oV}�ƃG��8���%{����'~�%�%�͸K�b���A@*l�1�'��$�Fӕk����%òaZ���'��P��E���T�^SRܹ��'���B��#1� �#l�}�V�r�'M�C@�
j�p��A�u����'U�	�ԡZaaP%A��`���'g��83�Q�$N��kׅr`���'�@a���(֨����p�(8�'3ڀ���٩(Μ��#��`��<�
�'eX�brK��h�:]���ߏ�%a�'Ϝ5Q������d�.rA ��'�
)�'nY4A� u9 �,cox�1�'�r�5�>h�.m3 �/I�N�j�'�[3b˭^?�d�"�ͻ0��D��'�v�!�D�L���Ѫ�)rS�'8>��#�A�Za� ����w+:��
�'3"���I��g�����[��J
�'Z>����6�rd�6M�X��,��'B�	j$�42i�C�M:x0��'�8��G�,���!V0K�B8��'&n���	$Vzh��T�K*;�<
�'/\��퉱~��,��&P1���	�'��ʑ��+T\���Ӯόx�d`	�'�Fu��y�P��ECjI"�{�'S �JQ�j������d�`\��'��,cu�¯{��t��_+̠��'I��F��b���T�Z��k�'�R�kk"-SÉ�(��I�
�'���C�ҝ@q��i݀+B�9�'�J��vb�18�u�SՀ[��Ԉ	�'SP� ��G��l�׻'+�@��'p,��E-�%0E�L��g�;&!� S�'E�t�QE�{��S�E��l}��8	�'t��đvT����F�gY�t�	�'�X�kG�]8a��KG�a����'�� rm�X�9g��Mdi��'�JQ�eC�s<4,������!��'��=Ac��!c V��9�,�(�'Y(���Y"}��Ca^?M�n���'��1Q�gV�����ÌY6������� ���A`	'3r����R��d�G"O
�ӂ�ʜO��3�@01z}�g"O�)�3�V+	��1C�0  �M��"OlP�E0}��c(B�w��p �"OܰBgM��p�B���f&=�$*Q"O���(C�Q���G�L'S[��"O�5J%* �g�r@�����$�H�"O�I�uI�i���.l�5yV"Oh�s�(k�(��bP�}16=�3"Oh�#�N�=9�����"3 �3�"OƐ��']	G�[0`S�c�X�"O@�c(V4:/)H%!���!�"OfݢD-ܠ}y�X�@.#�t�"O�`(P���U|�+�"O��;5��u�P|JfM�E�!�`"OL��Ʌ�@5�L{���-n/̔
�"O)��IϨ�I��tS��3��;D���4&��28�X�uN_=�H)4-;D���3f��~M��� (��2��@T�<D�p{%�WV}JU��Z�VovCFb9D�а�Я+����9Ahz�H-D�@Y7��o\J�B��zBj���)D�lѣ�L�eU���S)�&Qb���k-D������L�P�P�Ƭ4
hr+D���'�kt �g��Z9(��G *D��Д�_�p P�p�ӧaH�g�'D�ت�B�V86Iy�I{�س��%D��PC��o��A�dΣc�lb�$!|Ob��)P"��K<%�S"B+ 㒌�p#D��2`�A2\ bT'��]1��JP%-D� ���R�:n�)2��b����8D�����^,m����U��)�%�_-=�=E��'��W�:?�`��D_Oh�����'���
0$A�=b�1�#O@ጥ��'��������z�
�+�c��T�
�'�6�9�oA#!nP�A��^�t�j
�'
��8�LʹW�� ��U�UvP���'s�țug�x��@	r�ÿE����'��I���$4t@4��f�@W^eK
�'en�iM�<����<�\Ɉ�'f�Ч��y�� �E�G�t��'�\L*���< � �k'g�1@��3
�'��Xu,X�j\��  c�D�	�'
~���t|��Z�"<XNy*	�'4>�נT;/�D����S�1
�'�ȔB��0�c��	*�0T���A��y" �'��`#��.�p���E1�yb�P+j�HҭN�u��c���yr`�t�V�r!H�?�������=�y�*�86��=@:�0�!� �y2�G>���a�&i8N�Jpkа�y�˪s2d �+
Z��z��/�yR��hl618V�	T��S0%���y#��m�e��6O� 0���V~�<��KO�P��@RF� cM`ɳ�GTo�<�� 	�y:�ds�K'rȜL���q�<wB��e2l�k���;�Bɡ�Ɇg�<���il�Y�G�	��Yj�<Y��� ���bI��^Qᨁ�b�<�Ce�Z����U�c� iXAL�wy��_a��(�:Y��GL4$ y�o�0_����"O~��Ɓ��v��b'������c"O��p'�σQ�t����ґ 5"O�E��"�78�(�Cb֟��p�"O� �՛�'صY`%��Q�D�"O��!#E,�tST� (V�����"OT�s���) `�A�@&<;z,�T"OXX�>��h��"��)�v0He"O\ă�AϴN�N(�ǫ�)9l���"O(�HŃ�
^n��d꓆v�,��"O�!qt$LZ�x�[T*ѽ��	�"Oz�@aI+C��	��^�t��&"OL�R���R�S�ɠ'+:`��"O��x'I�#r�Z����I�F��"O
]vCX���P	�m�=�)y�"Or��1�_�\X^p��M^�e��A;�"O� �!�"q�TY�3v$�:�"O�%f� ��ђ �G��<�E"O25���,,D�R��0&yc"O��t	�t3^�!��t(��"OΜ�T>K:Lt��/T�}��@��"OL016n<+"����%X$���*�"O�*p��*�Tа3B�E�V��"O�����i�� �N�i����"OB�0�IY4yDL�AG�<��-��"O��1vm�~G`e�2`&���Q"O�	�AD�T�FLJ X�p�e�w"O�����3�lP+Ӥ�S_����"OR-��ܹq����!�ӏ9ԹJ"O���EĤ_�=�Q)D2��Q�"O>��EdM�#�P=���M-} ���"OJUp7bCW�ԊTf)P��""OX�j�kǒo�j�2����E(.hPG"O"�@�
�ch��X�l�8��"OI�B�����rGΏ']�\�IP"O��A�zȦ�c���
��E��"OJ1bY�Il�ܓ���	e����"O6�1r�S6L�H��$Y&n��@aA"O�@��M�5eI� S��B�Xyy""O��hE��(�ru2�	�c�D���"O��x�m��.��f�$��p��"O��ڄ&��>8�D_�t�1"O�H;@Ě)[Lp���ɛC�0��A"Oм��M��554`@���1�Xd�@"O�1; ,�$+˜0RD��e����"Ox���@�x�
\c�+�5�2��U"O�H�A 
�1�Y0d�@1��H�"O~���'	�4�r4a�
x�*��"O,�D�Ĝ"P�
#�ۅy,hqV"O Ց���D���p�`�Y���s"Oj���B�oHV��C�+ݢ(�G"On���c�"Z�������MńTj�"O A��C!�����%ҡ��%�"O !
�J�r]}�Ċ3�D�5"Ov�1��Π'H���c�9�ع1�"Oܭ!���:y6!
$�$w�f�"O̬ ��*cD�SVEO4_l "O0��&%T�nn����ݴ!^|h �"O����A�B�
(*�b޶YɳR"Od��e��zf��Z�n�$ �!�$��{|+���h�k[@�!��.�I���)��s��Ó6�!�֝]T@��tKӆXƦ@�c╯�!�D��v�p��ѿ0�ȍB����!�DϻU��C%���x�[��$�!�D�Q�������j'�\��!�Ӗ�4�i��!p�Q��c�!�$ɾ/�6���#ې$4A%�Pz�!�� �E����z^��� �Z5�5"ODqg�S*���q��T�i�4"Oȉ�s�_D�.q�WF1a�2�!�"O�Q�LX]
l#d��V���!"O�|t�E�����%��:�|d��"OVa;��@�`�ƙ�Ĕ�!��(�b"Obpt	�&p��[W"W�0����U"O�y��C>@V,�b�j��8�����"O���bT#@��|��IP�bE,0S"O�(&%�;X��񧄆$'"���"OtL� K�4]Ry���12}����"ORԛ&�o�Z�q�K`TD��"O�L��AH�T%�$���O6EH"O����,(r�>�#Qg�3Vlqt"O:������S|��H�\(�	(�"OH� H
�7!Έ��a[�0 �%��"O���`�=&92!2���b�"OV�1�Z 	&��GA���b�9"O�}����L�@� I��<9"O�P�+�'DHP��c�F�Z9qW"Ol�`�!��N��I�d��.]�&��a"O�Y�to��l�LL:k��q"O��!�N�n�r�ڐD��+R�$�$"O^P��ڲ8�Mq��@�:M��"O��IƖ�1!��z6���WW��"O��;�.B1��Pz4��s9�Y��"O�p"��3J��͙�ā<9�Ċ�"O�<HQjC@��<سb�>lzّ$"O����H�4Ao�$b߆<v�xt"O܍9�nJ�Wvpx�N�,,xi�"O~����/Q����d�
��C"OP@#�e<Cؾ��r��-�i�"O���0��� �2�sb˜��H��"O,8�d, ?������02!"O|aׯ�!�h���I��x��"O�dI���0j��ǁ2�ȼHp"O0�"A_Dd�<��矴d�F�J�"O���Se�3"0�s�������r"O��R�ȇooT����[�*�!��hA*��Wg������v9���"O@5B��'3����'ϔ,H3��r�"O�eK�K�4*C��ѵ�=$���#"O��!Iؓ]r*y2�� 
p l�yB"O�U����6ں����,��"OB3��״<��J�K�I!�W"O��2lS�|�k�c��5�ȅA"O���f���x����Z,U�pй�'ϾaX�&��zhJ-��_NTԱ�
�'Y�E�6G]<tpp�k���4a�1�	�'U�Q��>J8(c�֚D����'*ʐ�E��rV
�gφ���
�'�ޙ�" ��K'�}��$U�2���
�'���Î4)
��"�3|��:
�'�ء1V�r�(���2��I�	�'���;!��EX3d�C)���'w��b�Ë�`X�|��ʃ�O�p�#�'I~�jS�r�� ,ό�9�'��9�ğ3G���AII$ ��' �쑀��@o���~Ȱt�'4�t��.Ƚ1��$���`� D0�'�`�K'N��a� )4
(�����'��㵃^�.n0���	ܬV"�(s�'��%&��}�|��ƭ\�)��'��BU�B�er9��-:	2�iX��� da"��w69�Tc�2���q"O���BO�D�MqUG�4;�"�rF"OR� �EיH�( ���I�UZ͹�"O�)�
�T}��c�$U�*�d�U"O�a0VD��5��L ��f3>XH�"O�Tc�lO�@��:CA�a2$��"OX!i�&˗wg��K�К)�驅"O�At$?��i�� (��T"O���g��Ke�����0����"O���pN�=GQ"c*�=hdk@"OHA��(B=6�`�J%��b�"OHh�O��:�)�����p��"OtB�M�4x乖��:+MN�p"O썛�bߒ7��$�E�/{G�=��"O,��c�o2v|m�#2�x4"O*��5m�%Ը�m��l<�r"OXa;6��KP���ÕzJ����"O$�[w���Lx��\,`�3C"O$�3��	B\zj�d5ǊE�A"O�j�	�n)��Ƀ.^�P֘$"OM*&H׈���D.�7�"�`'"O\2�M1�~�s��U�s��e��"Oz�r�(ƈ$��j ._�0P3"O����D��Y��<s@�#-!Ã"O��'lH2 m�i�1`͈0�be"O~�2AX�b@H�oƅ#���"O��%J��b���"c�± Ѹs"O�h�g萸6�`i�g5.� �p"O����CٞiJ�؆VBl�4"O���gj�qФ��d%��T9F"OP���F�a�z���� IۨDq@"O��2N
g���gH�4(ʐ��r"O�Ӄ��PE������S�2��S"OV�ۣ)ʋW�j�b���7�>��s"O��YA'?B2n���B���F87�!�D̥\�L��%A']����uIG� m!�d��D��0צ!��,0�F\G]!��B�NV �9A��L2�c�sN!�$��8��)��Wמ�3���3Q�!�$� !Bb�C0�E�H�H�Dd�!�$�^G�}�B�R^���!�$�m�p9å��_
b�!Í1J!򤞥w貄1a�GM�r��!̡G@!�$�8� �q�NB��5j�o�!��ʥ3�స�ќV��7��;!�ĝ�u��e`�l�������B�!�$bS����'�X@`fh�s�!��=r��ar�D�q�B=J2eX.Z�!�:���%C�#M��S�J�<�!�Ė4��`X�Gʪ�L�94�ЂF�!��������M0jb������;O!��sĈX;�'I�,,@���I�E>!�H�A�:}��%�%�Z|�@lW�G�!��T�c	^�
F�Z#M;�ͪGk� �!��A�9�뀈%@��kH�!�_�3�����-	�(��ǚ�i�!�$�r�F`ٗ���0N ���ˠj�!�G8�yy% �>0�UE��!�D�
H�������R��x��bf!�ڊJP����Kl,I��'!���|���C��b^����Җ*!�D(a5�,y�ڻi#�!��T]�!���!���6oލ � ���.�!򄓸z��L���4��uѷ��&[�!�� ��3UdRV��Y	��Ηqv��6"O���F�  ��i�s�ț�8"O�t��IX	�l%�TIC�xvNmb�"ON��O� "`�"�iٗi�H���"OtԩgNF�D_���'��R�X�"Oj ����Xi��'&;6l��"O���D��-g5�t�D
��d\�""O�h`�Ñ�7���A���%��2"On@VB"�L�C�6W�b��"Ot#���
T�f� �	�!�� A"O�1�i�~ߪ(������S"O�I�@��3q7��8�j��P�"O �X�JA=eF����w�Й)B"O
���+����-�Q
8K���P�"O��� �HeD�PE(�6�F4j�"Oɡ0�V4lx�����M�jz@"O��2ԁR�r� 2$�q�"�Q"O��ځ+�>����3�� �$""OL�X5 �=Rhr�	�����:p"O� ��J��	�#�d}B�"O�@�p�6�Btr� r� �"O,=c�目&b0���,B��|R6"OL�q�>3r�;cWw�d�*O��ɳ
��!!�Dy�����'_.�`��*Y0�x�gd�I�$��'@����@�o��a�E� 3]��y���i��0$۶l`A��(_,�y���,vEȗ��XN����R)�y��΀)��Aj�!fP����a���y��~��|��ދ\�L�f����y�H^,BYt��蘈g���n[&�y% {�d �L�H��@Y,�y���(R��G	7��ʆɚ��y��D+XXZ�d�3��xu���y���%ӒqY�cĵ+�H��Մ���yBI*s�@wJ19�byh��B��y�(E��iFk4�`����'�y��G�5�H}�UG+輐;N�!�yR�
��\��̜#Jp�t I��yB�A�C�l����(kڄ)c��§�y�I�6k������w�8Y!tA[��y"�@;?F�4Qhƃ�"m��R=�y�'҂Q�2�� S��t1���J�y2�V$`���bg�	��,C���yb� �R��9��H�fO��˖	���y"/E@x��aꃙW9�������yr�ʐwI�qI���Oi�9v�2�y�J"X��a(��Zs��	xub*�y��4-l� �. #�H`S�H��y�%��x�F�Cl���8t�S���y"ݯ5��Q/C	z�E�'�,�yb�1{�u]�~���h��yr�FP�u�$��g�5B�ŏ7�y���5$˒��ბc'�Q���O�y�� M(P��a�l��A�2 @��y��Ħ
�zQ�G�	dL<�Pр��yr+�0U�Xȱu,cn��Q�E��y���_���p���*L]!P�P�y���x���̤�&�	�y�&I�	_�T��0� ��R�2��	�'�<Ī�N	my	�+K�I�z�X
�'z�LbG��J~��k"�׼?�F�	�'��9*D��V?��)���I�.e!	�'Ɣl!��3Y&�]�C�%2������ J����#m?00�X����"ON��b�O�<��n�(A��](E"Ob���L�5Mn�@P�0 eD){�"O� �OԵ��AB瘬���Xp"O6LX�%�1n�`��Bǋ80氌;�"O`ȩ��< �����&ۇc=��+f"O������n�Α��F�5�&y:d"O�q ��U�
 :��������Y�"O�|�V�ƳP�\�"����q��"OV�k�f
�)�0h�E����r�K�"OlP'��>\`i�o�-]Ⱁ�"O���C�L�a�W�^�u֤��"O@5k�Nl�P���X�v�l��"O�9�5!ޔ��D{���	�2"O����RN˚8h�,�
5��ɐ"O@�!2���:�]�R��;`�ypu"O 0�!��)R�D�)B н,�B��c"O���g���0i�a	5�ŏ(�F�I�"OTL�e��8��+E-vׂ@��"Ol4E�L�\�DXrʀ*o�h��r"O�D�ED�r�ؤ;���*�ɷ"O��§��''Vl�@��$E>0MQ�"O�8�A&��4.j�*b�)1%z���"Oxe V��2NU��-I	��9�"O>��5AT�/Z�\Y���|-XF"O^U *PY�����?��S"OT�s�jE�Y��� lR
h�<�c"Ov�Y�͎�Lա��J�vXR"O�:"�K���(C�-K�o���6"O\Ma����:j���E>	���Y�"O�2w�	�Jij}��E��ߜEh�"O�Yr��]L&�� ��A�-�@�R�"O���VEmK� �2��TʤE��"O0��Ѡ�(َ��cN�b���"O����T�d&�KU�QN֠Ÿ�"O �pUa��U�xyt&�O�\�"Omrs�ς%����W&?V� �s"O�u�U(� r�h�y�dQ�yV�0"OP)+ʃ;����CХ[K|��"O ���\k��â��>Es�"O���W�]�PK����(P�8���"Ol���*�ޖȀ���]x�	j"O�U��
C�?��� ����r�F���"O�Q�- ���t"�6�HY*G"Ofe�p��@bv�!�ƈ<t_�չ0"O��R��:pY��J����w"O>��EM9LD6a�5N��z8��"O�ݑiЋ��Ћ"MGV8�"O����+uc�Ta0�ݤ���"Oj`�􋉏0�9�m�'\ڢ�R�"Ox��u)O�ƌ��)�.̦���"OBa3`ⓂVъ�Id����w"O�4�6J�,n�ٷi��P����"O�%[q�ߤ)�L��u#ɛ
Q��Z�"OV��Ɓ�,_�ah�_Pb5��"O��[�AJ��`�Q��@�^ ��"O�wcZ�m �T�u�S�^�V4�s"O�"�/��'`ĵ@�IWg`Q�"O �$d����b���6�5�!"OH1��4"�,�(�ᄇW9ؽS"O�P#�%�	m���Ua�.:�"O�|��'�1'��M�U"�9���2S"O A1Bog\����:Y���"O,�Ə�-zzL���zD�f"O� �E;qED���;�JK82>E8p"O^d�����a�s��K0���0"O�Q�q @<&L�a.͈,����"O�,j�Y�,ҤX�D͔�+^���"O��7_��a�L�;fFȊb"O�a��A�}�����J"Rd吀"O��B�)��`����v�Q�5>$��@"O�9��Д(���"h��S��"O!a��Ċ_����Xs/,H�b"O�)��Ai���#F�:��ɴ"O��2�V�ON,,���F	֚y�"O����ȧwC����> �p�"O�ݺt	&��l0����r%"O���怆-f�)A�Q#0��ZU"Op�u��g��Xұ_(O�f!�q"O8��uNS7S
T�iCDu���%"OdQ	K�r�ó�ƃ.٢ zS"O8�Q�M��qd�13��2}ڀ��r"O(�	�G��E���@�k��"@"O*�QrCƇ3���b�Q<Lֹ�"O䌒�lQ�{�y�m er�p�"O�`V"��d4`i#E���`Zт2"ORexUB׈U���Ţ7/*���"O
UYr��ku04�/V+\dV"O��OZ�uc�@2�`�%��	f"O41Z�m�%� |���O%GL�@"O$ؤJ��.���7�QS v�9�"OV�;�E�jb�:v�͟(LQ5"O������6�d����S�l��"O�(x��,F��
c�5t�X<ˆ"OR�ʢ�
!b�bt�5������"O�%c�i��S�V���l�!B۠)�"O$l��F�SH,%��,�u����"O��+C�I~L ��+� C�rm��"O8}x���06l��+rD�{��$#"O:h�� ��߸r�=G��*�"O\� �'ˤN�\���&��Y�}��"O��PfB�>x� ĤAmOx��3"OJY!�,�f>t�n��bY���"O���0*��,��A9QF�MnA�"O^��0"�!o�鰴F̒fHpP�1"O,`Xth�P�����ӣ"O��gb�+LI�d9�V�dr�,�v"O�����[51J�x� ��ho>���"O�S�Q�]�����`ڶf��l3�"O(u�"�I@���F��"O�1���~���Hg,J;`�i��"OLlA��� 2�Y[ �ʟ)�mPC"O$I����5zT�z�Q�f�Q0v"OhD��ĩZ�y5�K���@Kw�<�K�	F8M����:f�A�A�o�<yƢQ<S�<��'��[�(aH`q�<��N�*Yb���ٴS����	�r�<aWiT�lQ�b�C��H���k�<�#�1\u�%����E�\u�rP[�<���0 X��q�� p�=���TS�<�A|���s��V��aW�LN�<�C�Ԣ5��A�%��Ȇ�X	v�ȓ��l�'@M�>�|���[='$|%��v�,@��a8��Pw+P7H�1��|��c�ۥt���1��'�-��X�H�k�ņ�6�f��U��(-8�����8#6!/�v����0M��|��'`P��ER?oqbT2c$@�hek
��� �4����%��P�ǩ�:Q�&���"O���*�"�8|���S$�|
D"O0�e('6K"��g&�`#��"O��F�� (��b���%F!�!�g"O�c�J�5+��� 7e��z�M9�"O�tc(��U^.[�6Ae�u�$"OD���gϴ@JՃBI\�!I4�*�"O�\��y��<0B�Q4w8nY�e"OPC�B҆q�%(�%X��Q�"O�1�6/�k��i��f~ȔXZ�"O�`�b��%!�4A��X�����"Op�E���'3̉���P�4��h0f"OhPyW���h��;]�R���H\��y�ꂫX��!Bŉ��ք����yRe�<.��i�OP��ꘪ�O�y�/��
}�ikp��y��px�@��y��;^-d��3���o	�x{q�S�yr���M�X@�rA��k������y�&�4�� ���2W�4���-�yb�B�s�
�0«SbH,;q�W��y¨�S�~a��H�q���S��y2�@�H�2ջV�I�Ţ���	�y���]��E����]��)VlƋ�yI��R��	c��	��D��y��W>:s������vv�0S�ߡ�y�J�%�n��%i�$�v�ɉ�yR�7f`���0��&x�d�������y�B�`��1B�O�t|��%� �y���G���iE�]�W�Ь���_/�y�rdmr�M�:K}���h2�y�ƐQ���a�H�2�a��Z��y���?b$,a��LW�QB� R M��y"���{�\1�0逳*JݑT�ͧ�y�O�|`L�m��% ��[��y��N�ܰX�4�܆V�Ld	F�E��yBiX;@s�X*M�}p�p�坞�y��@�3boR�s�>P����:�y�M�!wI�L��g_�e�J}�dj�+�yB��D��p)�Un|��GL���y�F�V��[ ,if�|�&��yRn]�* ��wv��� �!�y��� h��٦�-t�$�p��L��yb�ԒY��Ѐ��T�Xm+��y�K�^7j�����@���(E��y�F��Q����d֣(���A*�y�MP�Gj���h�'|���y��$�Nq0g��ml�e��y���������y�����y�A��@5$��"#42nF�����y�b�x��g�J�%9�bA�I��y2��h��Uz�˕)/vb�"��ï�y���0�R4a�#	@L���[��y�m�,!�re0u���&�P����y�&J�*�z;��\=1h9�����yR�!4|d`)E��0Zwr��7�y�'S8e�x��!�O�0p��)5�y2!̪}�*$�%�Mr�i���6�yr$���`� a]@v���qś1�yr��E[���H�D;���dc��y����$��M Y"��� Ā�y�*Ś"~�ha�!��:�*DT��y"hĦ�̌��
�.
�mr`���y���<�6�H�䏔8�8	H$ܢ�y�a�$D�4��)0Z�����5�y
� ��X�Z��T��b�<];�"O�Q�cۧD�^ aejC� ��d��"OFX�7'!^�u�j��w\Q��"Ot�Kӣ[�Z?���uK��L�Z�z�"O��Ǧ�Cr�:Wʞ==ϔ�"O�鐲��drx�j�*����@"O ��IT�f�pDJI�J�jYS"Oj��J	�hJ�h�+-� �b�"O�@���C��P����>�:�"O0���/ӓAL<�2�˗d ���V"O���T0KI:c�P�nɢ"O
�2��[�f�:XqFI&j��0K�"O2,�a�/{��#�n�/��eC"O�9�U�O�og����$�mɬ}��"O@������T���ܻL�H���"OقԪ<9��9I�j��!c"O~�K�{�DLq�C�?�f���"O��iR&F�)��q��5Mo&,h�"OP9��Ċ?4  (�T��(L�"OXZU(ɒ���ش|�0H�$"O@��2䪙�vA,'�5Z3"OD�pΟ$*��´� H��J�"O��R�B?~�Ψ���X#bj�8�G"O~���ˏ��b���@�	|[���"O������a�1l1���T"O�]� J�;^ڸS��ދJh9��"O:��QeB�F��T�v*K�{�L��"O.���:(�����&<���+"O�p��-ݮ���pL�9 �Y"O��SE^�E|�0�pM�  ��"OdAr��]���;��� z�t�"O��3�B#6juk�`��;�"O>��$']�1h49��Gvȩ� "Ov�اꋠ�֝"3*D�Qh�"O�@a2���y�!ɞ*i8�5#d"O����ؤ3�i���J��"O�)A �)a|�q7�W��E2�"O�$�נ5&r�I��<�z={�"OK�ň�wW��1,�CQ�ds"O���掣s�(�0bj �g=F]y@"O��;V��m**D�sIG�z9tA��"O��� �X�*]�3�:m!�
U"O���	�j$YjK�xD"O�Cڸp��x$�#:�p��2"O�챵�ȅ1�$�(�؂�d;@"O�h���QAҍ����"2�HА�"O�u�� ��m���� (F}���a"O�q��O�_��2��ǅ	hX�b"OlPR���i7��PƈĬ)K��@�"O5�-=��I��B����P#"OJP�)�1{b��T�KxP��"OZ��%��� �:e	��g��:�"O6 ��=nL3SHA�/]�1"O���G �hu�dxb�	OB�m�b"OH<�!+2�eڶ�ɱ3���"Oh���O:`ʨ�V��3	-$e��"O�!� �W _R�QW�?0&.	��"O�밨M&q��3#�%z$��C"O���T�ٝ&(�a��AH~���Rd"Oh-97�.a���Y#�j �
�"O���4��7�Z�x�+��X	0�0�"Ot��ւ?n�6 xak�)�t@D"O��20�����Q�)J�By�"O@��@֘����N�9k&0�"O� I@T��=|x<C��O:B�Ї"O�) h��4k�L����"On�2�AOs�5�B!U!(�нe"O؝y�A�t�w�H�DZe"O�JqID3Cdi��
K��] u"O2�k��	`��q�3�@x׺@ �"Oz�9���s���
��9��=3"O���'D ^����ˡ>��1��"Ov����C<�ԍq���o+>x�"On�d*7{]��F��0�4"OtR�"�h�H�!dg_5r��H��"OPe�gG�7}��TJ�F�P� �@V"OJ�X�����Y�+�?��� "OV�Ƭ�-���*Rj�<,�!2"O�8�g���Q���="J(Z�"Od�C��3>�E-Ƀ<��p�"O !� ĬCA�E�7m�!!����"OL�y���8�L�y���0u8
�"Oj���X�-^6���Գa2��"O��J��]�A$�-�bjA?*��"O0�G΂�x�y@��7j@��i�"O.��3
�FP�Y'�^�a7���p"O�(e@�o�z�fڙ>1��c@"O�h��#Jgd
 � �4 '� ;p"O��z�
��d.��3fo޴��R"O��z�YZ��0g��<�n�JR"Oڙ� A�[uZ|"lN��Vh3r"O���⫈�i��
� �_�܍)�"Ob�Y���A�ֺ�t��d��!���-zX��s$�+0���[7�E�!�d�Ep��d��?cdM�5φ?{!�dX�`����*RЀ����A�!�dH ƍj'�;J4�	h�J*�!��N�sh���e%��2Fj=:���p�!���G�����̗�w�x�y�G�%!�D4I���Bf�*��+�%d�!�ĕ�f�BPv&�lq�و��ʢt�!��P%6>2�A=�$��N�i�!�D�=�e3�#�5	_�� Ν�!�D�-s�l��E#L�>DY�cg�g�!�$���>�s���k������!���':�h�j�
�x�,���E�
I�!�D9W�EHVD��n(�pb��U�!��eTP��E�W�>Ę7���e!�*8�
�S��� ��C�'7!��9�ZdSp�2���ǆ0!򄙹F��ya�E�XH�& ��Ql!�^E���哳$qN�"���w�!��Uvc~���. �u{� >4J!��8xb��H��P�u�T�*D�8!��͎ T�ma��:y�Bب%�18|!��v��X`����z�;�H�!�!��9"��M�'��H�Fo�B���dk��4f�9 �<��P �N�ą��)�tb�M�=�:�`E��Uդ�ȓ��I�a���a��)�b=|jI�ȓf�Q�C�љY��@Z��B�$���Tn��14-�G`T�a�J/jU�ȓz(R�S�D��c
n=����B���ȓQ܌����]�m	d-]Q�����+J������bձ#�>45e��D�2D ��ʽ&B�Lc�;I�(`��w�fE�e�Q�p*��Ύ4�de��*���T�n�$���G���\��S�? �@E����IZ�3h�h @�"OpD���-PD��ꝗO����"O|���jJ^ٚ8�Q`��"({�"O(�9���*m, �2��!`	�'.>4�g
�;Ȝh�C��	Yt����'����!5��rb$_�l���'�,�2���^8��a�`؅Ug� �'v���G2%r�¡���n�0�'�(�W�+-
�q�͒1B� �'�<��憅�W�vtq4'ـ0k�ݢ�'�A���k��3d�U�P	�'B!K%MM0�>���
�O�2�b�'��M�V˕�yv���,Y�9&Ƶr	�'���*�.$N����F	�.]���	�'��Qk�&�m &�Yף�����'��u(�e���y�w!�5oP!��'��i3N9l��7�P��Z�'����͙w|����K�5Q�m��' �K֋�`zr��c.ƾ@�4��	�'�fXB�(F�l��	bm 3C`�z	�'ݰ���BĜ_����!BO7z�,1	�'���%�s�t̓��"8�^ѱ�'-L@@�$^(U�w�~���'ݖ}��(JW@�`ȶ��~.z��'��}3�lV�^�򴂶�M;q����	�'$z=��B�Y>��e$�2v`��'ʾtR�.�"ko2<)��Ս(�v�"�'�&���둠1ġ.� O2��''��gD�oE��Z��.0���'gH��)�ɿ!z��򅊌/X0�C�Iw;ޠ�B�%-��Y��D�0VΖC�Ɍ3�9D��'R���$J�SOZC�ɮ*�	��b�,G�5r��ę�B�I��R�ֈu����OB�Kp�C�I2�훔��
��G�*f*JC�I�9�D*�l��] �R�$@z!�C�	������x3,("C/ҾC�ɩ�j%sv� =/,�cL59��C�I� ��G�'5���0A ��z�bC䉩vy I�Gm�;��q��ʖw�C�J*b��%��u*���b@�O�zC�	�)8h�NΜ�xҡ���!�����̩f��Cr  ��a��z�!�dՔ@�4]ȅ�G>nV&y�e`��!�])���F�V$-S.�"�ɒ�+�!��ЀMH� ��L�}��H�o�=�!�$E�! �KdGa`N���ȯh�!򄌉H��I@2�V;�*h!��2r|!򤌶z��j�救_��T��`!�D/-)1�g�x=��AӚ&X!�D�).�N`� ����e��R4g^!��I)ngh�c���P��iW!����Bd��\w�v�YȐ*SC!�Dυ7R~i�ҁ&����GR1&4!�D�O2�C�h/]i� Rv&̓�!򄐞&D���	�<]4	�T@�+�!�,`��ݻJ�#%/�bM!�D�� ����O6���r�S$~@!�>V�lD�K��u��"���k�!�$C+�)8a�<qlh�B�\0T�!�d[k�ZDL`�h8���!�dجR���*Te�-�	�e�!�ڦ^��8�`��~*��"��̈́W�!��]]Zv}#�"^<�=��ʳo�!�� ����([?v��Hz�.H�U���"O���5oH�Y�� JC-�eJzi��"O�����2�^\9�L��NS�ȱ�"O�����
e;4�"��=B�N���"O��#��/w�x��r��N<(��"O��iFÓ�(�N��p�V|��x��"On��`���%�.`�0�ƽQ�H��v"O�d E�ݨ�n����D�8ނ9!C"O``I�㍉Y�Ṇ��Έ`�6H�c"Ox��q�T*3�D�B�Փ��œ1"Of-0f�:d��)��L��9�Q"O6�����I�>!��.�5B�<��%"OP0�S�%��I�ęmM����+D����x��e��/J�r��*D�x!�	 MĬ0t�֒	vrH@*O���5)��``�eӷ �/S2�q�"O�ˑ�,+�y[��=�K�"O^��獌~Z�8p� GN���"O����@$���Q#o�*�H�"O�|���3<�p9���\�N�<{v"O�l(eQ�W8�@#FME�\����"OD�-�,R�p��ˊ�|y�+B"O��a�U2
��5�4`��p"OTdK��<�6��w�V����u"O�t�a��c��D�`�3A��#c"O�ᑌM^N�8�1%@[	�'F�A(%��&n6��i���-x
d"�'hd4�u�G�?i$-Ʉ�����4+
�'of�B⺤qہa�}�u��Sd�<��yЈ����m��8!�AV�<Q���:>R�g˙J�(2gM�H�<Yea�;�L��V�_�Gr�y�D�<q�;H�����Cf��1��\B�<�� %�&4)�Y�xļ0�N�b�<���H�=T��:��I]��U���^�<y�/p�>|"CB��,9�y�e
p�<�!!��6IZ�C���#��=��h�<�V�T
C���ڡ�P��H,Ӥ�L�<��b�.U�$���I$T�HlB�i�N�<�ر[Y��""9z3X�ԃ[H�<����$()x}Vጲ{��H��A�<) $�C�Dܠ���3��0�d�g�<�ucX�p�N}�"A��T��ScBg�<y�ע3RxU�&C<
���sdz�<	vDM NN��2���X�d�#�
w�<y��'Z�|k�o�%0H����NCL�<Qp��	1�& �!�)��qddM^�<�B\��l����%�ॱ�@NW�<9Gn����X0�厤
�F|�I�<���[�@�pe��.�( ��"$�F�<ɡ�Q:�r�耽L���`j�Y�<�4�̸BgXRuΘ6\1����Q�<�2��2�L�TH��6�k�$�Q�<9�	��B2�o4z��d�EB�<��
�,���ԑ|�`i��o��^��C� k�9
�D��Y���uN@�B0�B�I�[����q.92Ȑ���C�M�B�(U
I܈BԐ��W����B��q�b��lԄb���U�ަlB�I��6"	�p+�DJ֑��'~P�ȁ�"GA6�� mM�;F��B�'G0}yR��en�����8A,=�'�����l�v�P�#e�!.P�e��'&|��h�>�xHj��܀-4������ X�q6�"�,�hUX��E"O�P�f�Ó(Z*$�N+sE�\�"O���L��Wwf��D�� R4@4�"O�TP �sІt �1K(�)�P"O��A�M���Cr��r
��"O�L8`F�2�lU!,��UT��"O$�6���q��Xu@E�S��89b"O|�
���&�F�=k�:���"O�T�/]�Qd挫�eӌ˘\j3"O�@f�C���@��ֹafr�x�"OD%ڱ�x�D�` '�_8B#�"On���+��i����	)f̰s"OR�8��:h���R2&��bx3�"O��`�)anb�$�ȱ6��œ"O�t���$DKIyEM��!�ZqA�"O� p�z�U��&Ҫb�ذ*w"O�1cQ �3w�h���șo�\�T"O&�PĄ^<7�8za%W
.æ���"O������V�>H��䋵!�dk�"O�T(Ҡ�??�SwfQ�}�v�A�"Oj�Iѧ��q�|E����pL(q(�"O���3�6ܘ�A�d.l�"O�� �=s$ȋ4�(H ����"O�K��Tl�UO�r�$YW"OR�05f_�.<��;��ØI��"O�@�S`��#T ��ጂv����"O`!�a�FŊ�)$��)W,�b�"OnкR��q��`1`�;� �"O��r����=��֬
'@ܢ]�u"O��!�UJ��k�Pe L��"O
E2�΁�:BN-��I�a�D� "OTlZ���!j��sǘ0� a��"O�l�g!~mzv��!F�L���J�<�cسj'�9���#XW��ÎKC�<Q&Z�I@�;�F�Z|!ӉT�<���#|^�A1��+�^�9��S�<���˦H���;�^��N�9�bP�<!��:N����N�r�ݨ�@AM�<�v�P!���T��	�d)zPJ_F�<	�Y0-�����R��đp�B�<�c��j4Xt���J	a�Rɢu��|�<Y�J���\�����N�`:���|�<�3�W�S�p����3Y�yf�Lx�<�����7L`I�O,w3����Lx�<��6�z��s���b׀��@�q�<Q���vc��@F�A&��C�y�<I��%��)�$�25��ASr�<�+V)�^�J(����@�D�<a�GP�2\Z����Y�J���DC�<q�E��-@%���ˊ*X�P%
|�<!���/݈<`#�ݭ_�T03�	�z�<	��L�r��O5[�����_|�<��4r��Y(�60F����B@�<�u界8�BD�FKM1Q��ّ�KYp�<!��Q�f����G�ޮ(QS6�GU�<���QB�\����ڱ)�TW�;T�`���O2E���s�⃫n*hQ��$D�����Bc	�%@���'e�2�)P%<D�sF�]
m�Z]h�BW���$D� �DM&Ub��\5Y��p$D�� �"��d�,؜5	�{E�-D�@8Ah�!���SHZ.X��d�*D�DY�n
.:���	�g�k��h۰M4D��``��`�jy �#o���U3D�� ����gM�k�jI��`�V�`}��"O�M�G-�NV@��w�ʥ�.�RW"O.���[7b�j׫π@q>���"O|M��fHg���N�IYl�A"O�q�儌�oA���M9HU|��"O轑����Eof�ar���X�"O֨x���N���k3��3x5�QR"O����_)a�� DG8��Ӗ"O��kT)�7j���ۧmE.Z�z|�"OF &K\5�h)�"FE�a_�5"O���Rh7L���8�V:N t�"O��rJҙO��Urt���FD�h�"O�H�D�Z�kܸ�ᎈ�\Fby`4"O��UB�P厭�d�[3p@��"O������dX�r�(�Kd`��"O0����3�������zgH��r"Ot�dL�u̸52A�A��A	�"OH1rBHL�M���S�?RĨ壱"O������r�����Z��h)�"Of����F_��	H�B܌1	�"O��CD	�J�P	���l\ZP"OR���O�lȈ�gPyl4���"O8���0~�݊��6�}�"O��-�A�H�ʖ%�8#� ("O��3�zS@a�%��@�$A6"O~��p��i<=bU�.$���"O@���&�Y�X�1�A�#�bB�"O\��O	C2L�w�S�-6
�q"O�Ѫ�M�[S&�����
}�5Z�"O��daU<W<���՜6��Ȫ�"OrX���3uO|4��B4,��9�"O�1�$xv S����8r�$!%"O�ij�_�C���2��m$��T"O^3�,��M�n���U4�|���"O��ZG�\�^��`�]�X��"O�|3�F�g\�5��.A%>T���"O�0h�(�Y�p��k�W:�,�r"OT\&O�(?;��h��ҳ~6 ��A"O�0q��#Fw�}��c�t':�ڐ"O��s'��<j�^�PҡK�5!���#"O6���Yh�v��S�@-ap@�"O��S,U�T�����\�{T�:p"O4�⧈эpLH(K$��_;N<Z�"O��U�Y�AB�����63�\���"O���	���1�C��*�|���"O@�
��X,^U�T�򆨡�"Ov�q���)Y~�8�@�l��b�"O��@��H*U���q����"O�a�b+�8k�H��R���sָE��*O���B�5I�4�
`Kƴ-ݸ���'!*$"B���l��xw	_��N4�	�'�l�:�o�@��$�������	�'lX)�����@�Dć�6��
�'�ܹ1�k	�( ȁ����@]�	�'� �S���6�չC�|���'�p�ÄR�:|����xc����'��xF/.'�TP�QFkf�D��'�����B�Oͤ��mH�T%���'@�X2`jӎ�:d�	MF
��'l���p��,'����Q�S�(T��'�J���2<����+��v"Y��'Y��	6�������0��$���
�'��p�� R�VaCe�̴���S
�'`�-��L
�ȣT��!c�.2��� ��S�f�!?�(�hG.UL��R�"O�xS���,lh����31���`"O�T�!�M�`R50P`�T�be"O�쫕I٬�liW��?�H�3R"O�0G�!t�0���!gƴK�"O0�Y� �5]���Y��ԔWBʉ�"O^��D`�p���ec2Tt"O�D��V��D��D�	�,`�"O>��L;(��Q��!>rU{�"O����hϝ[�������<$E"OʐqT��?!`����]�F��Yk�"O(�n�%uV�r���%sܡ"Of5�e�S;Z�I��hn��3"O�i�6D��1~�1"V!O`����"O��"$�8%�^ur��|Fة�"Oh|��B�1=��P�/'q,�1��"O�=��o��O��h�EO49�6"O��صF]P�\��僉�&7H��"Ox$�AbO��(z�B��z��P2"O�-���-T^����	rp0�yg"O֡�TP'Xi���k�d;C"O���CjHl��ၵl�!m��9�"O����n��r�Z���D����"OH}�f@.~B����A]9ZOT�:�"OJ$3F�,?�F�0cǟ�DJN��"O�9��i��I��������f@U�%"O�Т�Ĵ2R��a�$q�)�"OPY�Q"�"\W��Y���<~5R<
"O��9!i��2OV���Ån5؉{�"O��J��	�|�3D��(g�zD0�"Ov����>TA�M^;6>Q"O�!F��	�d�(z���"O��ʇ��+�^)p�LB,���0�"O�|9�O3yl���˛�C�� �f"O�2@��\#.��ʈ�0��U�"O��+�����h2	�%y��%�G"O���BMё.I�T��\
 �I�%"O
Hr�MD�?[�e�O0���e"O��@�&@�⥎.�%"'"Ot��VH�6.d$�Ef/FA� �%"O�jE�iW4�E�T;��{c"Oz4 F�>xD�SbN�3��ۓ"Oƨ��g�Z�nTf��"?	n�SG"O�Z6+ŭ�L�A��ך%�@L�"O& ��H�a��p�T�\;����"O �QdP�k��Y�"AF�=�$�0"O��h�M˱/!�Yª����@�"O���%�#�Dlqg�	�@U�2"O@��K6`�NK�2%�0x"O��2i�J�RDy��D��t"O���F�N���ui��B�[�[G"O��P�oT�S,إ��"I�,ID�`"O�}9��L�h��1���>jHtt�%"O:\5MBT��ā3 Їr���y�$^�
$�d�0P���ɇ��y�k�(u��J�l3Ua��[�f���yX�8l��$N�N.��:p���<�ŮVb�j��"��.����@��u�<�,�#!0��� �ŞѲ|��Fi�<q�&�T�JKf�`��� f�<ѧ�F
&6˒���:ڒtg�Ly�<!�hW75�lĸ�K�7�<5k�*k�<q%H�1G��D�č�}�N�J1�j�<y�$4q�����7�x�:��l�<� n1b��;g*:0z3͊(����"Oإ��+��D�,���J�
)��U �"O�*�ʛAJ��V��G�@	H�"O�c���%J�TĻ#o��/|z!��"O0����6f��DV�L��"O0`��@�7vb��ڑ�`��U"O��۳�X�B��`H��I�{���`q"OȜ�u.��YH�i�d�W E��5B�"OИ���o�L�"Ɖ�93���"O��sB�*W�X���'Y�Z�ĔaV"O�)s%�)A.Y�qM0r����"O�i[��D�T����e��Vt�pr"Ox�8��XpzAJ�ѠJX4�ؠ"O�"ˀ�`�`<KW ^�V�^8:�"O1��� !A���t���~�A"OꉺU��S$������.�"O"�X5�j{D\�S.,��Q�"OF�P��-,�֔Q"C]�|k�9#b"O*��$��
P�@_"y���"Oh�ҩ��Y!�Ja�N)
�"O���fm��S ��� ȍ3lzH��"O��2�5h�Pq�܎Y`�X�c"O�A���+�
��r盱b&l)�"O��!"�+��8��[/", 1D"O�US��51�.����&#u`�Z0"O&��2Eق����H�Of�ɋ�"Ob������Ȕ��<mJ��C5"Ol��oÇQ5>� "�R@�Q"Of�1AIJ�`|cb���Y&�u��"O�(x@i�0��yk g�-L4���"O4�(è�&��U� �y�Z��6"O�L��ha���V�٧7��$��"O~�� �� ���eөd�,c�"O���w.�
��5S�Z�R~���"O��: W��	�4nnƂ}0R"Oz��C�{8%8ujL�d��u�"O��Y�B�H�|H���G"k���"O*��"U+0^L�)��Pc�P��"O2aT;<���beQf��5)W�'��J^��d`��I<	BPHE <�!��T�(��P�l*ơ��R�A!�d�<D2��C���t��Չ�bL�"!��A)zP��[��b����-�!򤜈�r��
P. r<��]%|�!�E)2�t��u�E�@���Q�b�R�8O��g�)*��p$l ;�ƕ�S"O��°/��UBcX6`ޝ��L�<�����,� �Gܻ5-v��3�A�<�eB�Il�};!�@9"�h8��[A�<!g���К�o�2
@�;Q��F�<%�B1@���C)����HB�<Y�����Y�C�4��TʒT�<�W�B������$�:��ƅO�<٠�W�9W�A{K�
)�Ҕ)��BO�<e��_�|m�Ek�U�$�M�G�<�!�ϖ0����n�O��) ��C�<)�ҍ)�r���O�k�p�l�dyr�)�'c�lŀV	�%&ȋ
R�=:|`�ȓ6�� ���sw�qɑ+��ȓe�xdN� g�P�d�B&a����ȓX���`�=E4p{W��� ���]I�Ua�;Cq�`�p��~��$��p�l��MB'ߠxAB!�G����ȓq����q�"_��1y��ô ��E�<�M>9��� �`�CNؘ� r�)Zl��"O,�!��ԅV`�`�Ƃ�=I�9(S"O���Ӄ�b������=hv R�"O>�ٓF� m6�)�1@��XW�'"O��
րIN��1��~;��PQ"O:�u�p�Ӎ�
� �K�9�!�2a��砐A�Lrj�E��'o���O�=���$R�$D*�qt��<$fA�$�i�C�ɑ�Z4
 ��Ġ��
HȊ7�=���b
�%hh`)q)�J��<h���d�>1�&w��2�#ș��D�aoU�?��i�F����I�3�Vh�1O�<Bq����8����D%�߂V;��k�%���!��?*!��N$R{��ȁΐ�Y��ď� t!򤅰����#c8�<bs2U !���J�f�/BZ��$c�)-�!��S�1O����O@��D�D0��'�ީ�aʝ�)L�pb"�B�Z��!Q�'�H�C��wN~��$��JdZ���'�� ��bTx!��'x�}�
�'!�p�Ì"?���p �i�`�"	�'�� B'֡6��X���0����'ܼ�@�D���N��A�-q�$@�'�RtrvJ1M3�4�VK�2[���'����q'ϝ9	bd	�^7dt��'C�9
5�[>P��s��ȻFĢEy�'�.H�P���6��S�� ?G�3�'Zy
���1v��0�� ߜ/�f �'X�9A�A,(03Qm�1"%����'�|z$V�ty�怞��}��'1��p-�4-�ZmE�&~����'޼�"4a��M�e�ݑtQ���'V1k�FO�b)R����\!p!X!S�'���&��O֔�D��=�S�' ͱ���>	���\�p�R��
�'� 8`B�_w���fFʊb�L`
�'�
���O'J���ŧ�&`����'pH)IԢ	:`�����8	N�P�'��u@5� ;��!��L% ���'�R��!߷	o���c��@і	1
�'0rѨ�2���c8]�9��'1~D�aI�_X�fձ/N�0�'�r�[�LƖ7���&}����'^(s���r7D4zF�r��=c�'�2$��FN����2(A�i���'�~��#Ɇx�5b��R�ih��2	�'�:��$߈>T�[���Woڙ�	�'�`	��܏D��Dc�E���jX	�'������
;���G�m�p|��'a��d�Z]�����6;4�A��'�¨K���@O��*5+ӏCl����'C��9�-�`�$�q��:<n@���'T�A�rAkTPj��X;�����'�]�Da�*$y�Y��6=�a!�'~���=��\�c�ݨ3�M��'n�ajU'[�K��!;�G7_�`��'F�)z�$�n���w��4d��Q
�'�-��GB)J@y�v��2}:Ԉ��'�j���
���JQ	t�����'����aE�;i��b��ҍx.X���'@� o� c�"�0�`�fR�A�'��yK2!Dd�P𡰬�k��r
�'���3c_�Eb� Xd������	�'�L�Heo̗YU��#m�(��M�
��� ��Tb�fX�
�	��Dl\��"OB�s3� �@yaE����@��"OL��N�A,.�Z��9j�6���"O��%GГj"����,݇Nɔ �	�'�4X)�q�\ 8�"�F�bi��' �@q���7?�*�!Ӄ�0
��)�'���o�).B����e�/���'žP��+7�tL"ֆB-L��p�'��JE�0[�qX�O-'�I�'ڢ��а^�Pa����"�"�*
�'���AL�)F�2�R�%#"��
�'��@��Գg�2U�b\�$�@��'�Ųp/�`��#�ա��\a
�'�\YakC�S	�i��BF��H
�'��0�g"@4:]|�B*�9���*�'��3�D�	ޠ{N�+1�$A �'4��J�.���I�$xZ��'����Ҥ�+K�F5����$1 Ȳ�'ν0FhՏV���3�NX%(5���	�'::� � F �r�Ō��(	�'BА��M���0�i3��5 �\�	�'b���թ�0D@F({��V��0z	�'���S �l2B���Q�Ry	�'u��뒡����Ë߆��*�'�dy���
�lI0,Ef��$�Rn�<!�eH�?v�b��u���E�_B�<u�ڰV�2H�I*2�l@�A��y�<	t%B �~ik#ĝ�bT�)�!�a�<�檑�H��`qwƋ:h8 2�_x�<	��J�aH�;�lJ�hÞ� �K�I�<Q�E�'}���ǧq��
F�<��*�=5������	d`I&C�|�<�G�P�������}��} s�v�<!����)⨖�%�F�Ht"�f�<A��˩T頕��[׮�P5l�e�<�p���w����K�'fN��r@Dw�<)�n	'0h�U� I�&kRJ���e�J�<��JR�>Z�up3�Ǹp0N�C�<Y��z� ��a�ѷ,� ��{�<�ca��X��Z�&z�e���t�<IЏ��Ḙ
F��d= ��n�<���Q"1�$Q�����<@�.�l�<�-�G�F��B� �V�ʤ��b�<13OE�W�p�R������ -�T�<�D�Ch���(C+{��e�G�i�<9����pu�t(ޣ	�|���z�<� c�a�P@wC&��DQѮv�<Q��̫m�jZ4e�&B�2�S�I�<��"E
8�3a�Xpz�rw!�G�<aRO�L��8�s@�1O���Kx�<QP�^ mLTpp(ޞ;J�$�~�<���ΈxV�M�%^�*����f��v�<����v�
�@��Lw���l\o�<R�@$x�(�H�P���c�<i�Ï�Fv�9P�\�Mf�XZ�<A�M��Y��M�ql�Ll�lc�U�<�b��bc�}���O�q�)��m�<w	^6|�\t�ǥ54#���_�<�D��T�|�9���\��1y�a�B�<�' �e�%��埜�`�P�]�<C��*��X�Њ��r>d}B��SR���3�H���D�0�A�9�e��Q�5��GC#D�+�$W�ziFy+s��_�}H�G;D��ƌ�
_�:@���d�X0��4D�� �)R`��-��a2� ojp��"O��Q+W.0(f-��D�;�"O̕"7��P��A��\A�"O���"�,n�b����X{���"OT�)��E.1���Fj[����2"O��qIh�+ClS�%�V9��"O�ph��y�L}MҔ�8+�"O����0���Ps섮*6�+�"O�V-�kFT؃ծ[�8疼y�"Ory��)+T�Œv���T�j,��"O8�� �� d\Z�HW V�ܽ�$"O6�fhNx���G(��y�*�I�V�
Ee��9��A�'��yB�D�?�p�Ef�ށҷ�K��y⅞9�t���I'[�� ��y�@�b^�� e�ԁC�9�$�8�y��X)�$+�E�7��l�J�!�y2�ٗEX�XAg�,ڽ������ybKJ�7���1�_�.WV0s�l!�ȓB�Ȧ�Nb(�M�!���n�8p�ȓ|�t!��]B �ZP]D�@��K�Hu;v�:H4����B8~����5�H�eD
/Q^��`o��a 4�ȓ'�b%� cB���j�.z�
y��T�قF�U"p�4Cw�+C5�ȓU����C�*�~y��";D���ȓS0BP#���+�鑣�Ý]^@��qێ�h��Y5&0n|+%�P|/�d��~�j@۵A�6c��5kc��I����ɉfZ ��&���D��D�(J�
6ݴ.�̅*�l�AH<)S(ѬBN�񐄊�_'��pIRR��C*AZbƐ"X� �x�aI�ݘO�b�ԣC	݅ͅ]�rx����yR�[�Ĩ�B(;J�� ��Ӯ	�d�%ˌ(���Tl�<銈�Y��"��T!v��h��OSha�9q��#D����gƸqVP�՛T9���!��>b����s[R�aՃ؊q8���DS�C�rx���R�v�ؔ��Ł{azRi�;@h�С�"@�>��	z����0d��;P��9ę��x���M��@�q%^$M�j��6�-#u\���J2�$J-"vT�����P�Y�j�j��"r�%.9ٶ\[��K���|��E�!�tB�;.}%�O��t�PS�c.�Ӳ���j����q��6Q�1���{�'*n�SQ7�$D���B�]�T]��"�:C"�h�Oj((�x�����?��ɰ�LA�N����e���jX����0�T�hOL`ŅW-����bN��+=���c�'P�(�C"8Ծ�(�γTQA2双z.$Hr���2El��T T��0��%va}rG�4��!���� _4�,zՏ;��I�@�`�q�Jr3�`+!f�6ap#�+F�G��u�O���WƓ�-��@U���y��*	�'����&U%L|�S��T�h-�PJgDy�t�]2PpZѨ�P��֓�J͐f@P3�yG���`��H�ǋ��L�ڵ�hҾ�Pxb�L1n�^�K��׎V}lm�@�}^M��< h�0Gו82a�@�%l�R� ��\&x���	�&�\0,*G�Ƣ>�u���ic��YB.�d���ʍZ*nh��V�M�Ez�@BIl�Lz���4�f���
��&����(LO�<�"E�$z�
� c��!F"�Ѱ�'SPD���P�1�`ZTb� ���'|��@K�D&�ɀ��*Pl�[ūV^�>A����2��=:āF}H<��bL8�F��4��+
ڭC!��7&���Ê�H}��Ґ :�lt���L:�L��$g�* ҽkAoF��r&��O/v�:u�M��~����Im�`��CO�=K`�@� g�ዖ��e�!o\�b�	PF�n6ĥ�A�����V�`���6�;c!���^y�M�-�C$B�?\*�*S����O���D �(!j'ȅ'x�p8�&�{�Z,�I��[{���pᏋR8\�r��[�22��Ňݯ���#�.tɶ��#�K0���}<&��p��4c��O�P�W� "b�JGΚ�N<<�����x�$Y�s�!��� �H����*=Q��`��s�z���o@��a�j�M�ZmZf�5���F�c��}�KT%c�ƑQ#a^�7l�0�'�.3�n����3c��aR�)&pyj��Dam���gW؞��͑"�섻�Ұ 4f��vA~���i!�ŀ1�#ƪhX,�n��@<�#� /<h��@�z���9��D9���/�~txO�=��1#�T�6�(�>!% �)B��aP�`��P�L��V	���2�J!� ��3��]}'�0��,�/�l8�!Y� ��!��⌱n�
	�r@̄ ����$@�mըP�'kϵ�R蛲 J�o�
0����7{��h;Pk�<*���/A�iݸp�W�O��Z��2@�i�����4@e�L���ܼt�$͘u'N*l;$�p?14.�"��ڶ, *U�fLCdǗA�\�3�O#k��M7LvHa��D;'��چL��P�|`����C1N�U�4�T�ɼ"dܱ��kV�d�a{B䌺Th�T#�����՚k����MF�<��M���U�/�D��&�ʫ�|��3���[T��bN�i���"𭆨?��Yá�O8Cc�cj�\b6!�,�z���ÂA��M��l�.Jk��1�I��n�24�*]'M���
f!�Wz��b�� u����$`�<Y!eW*<������.A�Y"&�+�� �ٖƚ*AOX��� �5x�@t�@� �i`��JD��Z�M����&
�
���F�+��d�/΢ᛴ�m
�逯��Y������G�g����N�����'�@���-It䱠�8JF\�RO�\��r���S��3�$�-�P��5..Ih��شt�����w�T0"�0}�2����L}�K� )|O�ٔ�8G �� Ĥ�	&� �s�%�Nѐ,��P�/�B��!9G��S��b�K�$�d��v�)�Q����D��=xr�:O�d�0���"8�X@$�G�gv��$��ӄh��Pt0 ���Ĳ��<����\�Ё�EB9U0,�7a�Ӧ5����9w�d�PgJ�G� (Eb�O&� �E���w���wǺ��$�J!\]��q_�p��d)׬J���IP��fق.��*���ۇ3�کqÃ_?P�|0�-`;����߅Q�2	D�N$x�#)S0��U0u��B4�#B�>q"i� ��?
�(uB��H#&�ɇ0���K�yb�18����6 I�n(P�}�.��Q����
'�,� AN�uԌ@���'�tr@nI���Pg�Ht��O"ؑ���1ݦ	��# ��dC�[+/4��>�M�0{;�"|��%ͬ���RLu�H����>!�)�:o�����Op"��qJS�i5�A���_�Q�!�DN�m�乺��C�t-�x����k!��B�+��<c�� ��cփ�sW!�$Y�����Mx+V�{���v�!��]�~��\Rt	ޏN$�$
��!�5q7j�jt�����{���o/!���[609KU�cn����=!򄉒5��� �צ>f*��D�ͽ)o!�d�X
l�Ӵ%��vJ�����#%V!�ݥ#��xf�EI�e�R�U�'1!�D�� �,M e��0�<q9��5Y0!�$�>0<�!Z4*ȔoL���CN�v7!�ċ!P�)#s�۰<&�b�g�8!�=��X��L<1��D�y�!�d��2D��
��#�رp�̛�p�!�DO ��m� Or���C� �b�!��.1�0�6�P�z&9rą�O�!�G�B��e��Fl��j�!�$߾Q��M� ɑuqa%�%w�!����׀˱]m����l�-/�!�$�#w�0�v!G�n��kN�f�!�$�1���!�[�r(���9�!�$��r��Tvf�)C1��҂�E�:�!�d�k�t�����.���o�72s!�䈼D����#�T�Pk�5K!��WӔ|:YYzu�R�Av�~�ȓ`n4�!��"�VI�R���ȓw�0����I9m4���N �V���ȓj�`���.kf(9�o�#P�	��-v�šT������p�I�<4'�I��1�L�&%D�E�P�hs
Ӆ{G m�ȓ-sV��P��4G	TD�5�٨v�
 �ȓy�\�굤�5�� �A����P�8D��)�b��p*&H�$V��1�n6D� �D)	[q膮$f�Q(3D�T���G�y(1`�'�\m����H5T�c�_�l�BA�uD�[�0MC"O�E��ͽ#۶u;4�F�t��{�"OFU��
Tt'��+$,C#;TJ�R&"O�1& ��R��fk߬G7�"O��Qē�8@�A��6�J��"O�ui��^��	H0l�.�i!"O� �LjW�Զwv�	�	]��DyH�"O����CFY��GgՃY���p�"O�I�M !�X��R>A:���"OP��'#޹Dv�"�e� ��!s"O���'c�@I5�(�Q��"OZ ʇ$�+z䈹A�;ccp��G"O:��7��#T�zh� �9.p>�1�"O�*�)�jH���w͂2��-Е"O@� p�Z�M��ȩ��I!w�\kG"O�(�c@
|��X�u�7sf��""O�Q�D
A,h���`��CQn)��"O𨇉I�p��I1%�&\B� !"O�ј�/֥~Dm��R�HK�G"O"()��˚:��=���GV�4J�"OD�	U)ۻo�\��a ^1�Br"ONi�Rc�)��u��jH2H2F��""O.�1�l\A��Ua�CEvM�""O8���"�7�^e %�Q=f"�� e"OJ=[���72�
ݙeY�4 ����"Oœ N�0�΁vDVp� yZ�"O��B�[*i���� >�Ƒ�5"O� 9�dةU�l�PT�я8S8�U"O�!(ӧ_�D��*��C��\�D"Ov���C�95��+�]J405"Ozx�"��&i
t#VI๣"O
�Z�	%'X0��BF�V^�ұ"Or(��F��,�u�߃r�&=ZC"O�$���Z���|9�/�zFy"OZ�@�d�(�pLH
=Q�8��"Oz���J"Bx�a�k��nV��He"O��ʗ��w&��"�W+���i�"O��+G��&e���7ɞ'p�2;�"O2�R��5$�pf�M۸�c�"O`LA��?mBm{��J�h��ĨF"OH	�@��5�4bE֏"����"O�i�l�bnsC�N�C���"O*Y#���"�Na8У�X^v�#s"O��1� i_rܙ��74 �"O���fA�ّ�ō�R����"O��B.KZz*��EFր<(�DJ�"O����.�Z}��g�\��p"O��8�&��Gɒ���E�*~���9�"Oh����q;��ȃc�x��xZ"Obhs���1��e� �*1}V�h�<�5
�B�XM�#�5:ȁ���x�<7��?bE��-Ҕ0Z�%I7Wy�<�@",�X1�!���3��w�<Q�˻�JT��ݚic���pJW�<Q�(_�x��+F�' ���Mj�<�Pd�a6��� 勒 �:���_�<9p"V�,��t��C�t�@�ARZ�<9t�)8�f�W$
Pf��#-H�<QA(q����e׽2����B��]�<���X�_�t�'N�4*>�¤ _}�<P��]\L�K�44�ԡ�'�z�<�#�C�~k�	�FF���d��<�@��l� AWbO?5��A�q�$T����m���r�NڋDV���n+D���V�G�_������a~,07#&D����/�f�<�P���c�l��(D��ۆ���}X4���H
 �H���'D��5�حJ�M05�77[r�8@�&D���6�E�{H��f$X�q�H,y'!�B�8G���ڏr&�SS$@�!�� :� ���6]��`b��H�w(�mc�"O��`EM�)���#���(�M!"O�[",�%$VE
�G�;�����"Oni( -ŰCjp��䉛ܨ��"O@�H�%��qxx�Y�b�j�,Tc�"O�x��T:V�� s��XP�ր��"OZ�	���!�+�z��X�2"O`�����=in:�;)�yR�`�U"O��@�h��u�X�@��&�vY��"O���$�̦DGJ���g@�]�b8�"O>��Q�$*��ÒoN*F���ٔ"OX�q�`��X�RрJ��#�"O����Nބ�l����ܙo���ps"O�@2��2dMJ�*�0O
��r�Q]�<�E�.����B/
����r�S�<��!��:��qUk�*�
��P�<Y��܉Mv85��D�+/����,�D�<��
��smǧ%��10�]�<�$B |�R-Y�nA�X�f48��Z�<a�L]��ܩ��Ɣxx�tbsg�U�<�����b��
?|�����n�<a��lm�8(� ������!���,yk%R���Cf�2@fA�I�!�4��ݓ�	 =j�r�P���i�!�$�aN����D}S�ك����d!򄈺R��
a��E�8hQ��
4U!���]�,��r�ԁV��hi�C��DX!�D�:F��DX`߿���@Q�ӱVG!��ě�D��c�'	�B$*�ǈ-[8!򤕩�p%Y6��^�4��F+B
{3!�I�=ǜ�Sd�I�d� ҥ�ʴ{S!�,�PX�$��eUn���%E(!�DX�c���`Sh�3)^�Q�c�W:@�!�DZ"��1�D��F9�Ʉ%S�!��_e�*%���MA�Je��%J!�z��;Q�ǁNK��8�I�-�!�d�K_�aYԮ�=��S�ɾ3!�Ē[����g��j�y�KT%?�!�d��A}��z����%��S�.�X�'I.��H[�&d鰧G�Ad��
�'�NY�j�/\B%�gg9<�
�'LL��МLr�a1�i 2-�T���'ԄH0H�Pv��#6h�RODm��'[�ISL̤22�lӒ��:z�,<��'��ॎ9�
�KbG�!}1�9�'!�I$��@θ�ч�kDڰ��'�p��̓"?�� �@��m�����'לTh.��4�N�9���m��B�'+b�x�e�9z�$�%Y�+0!!
�'��M�Q��<q,=ōʥ-Dlb�'{�љ3@�{�(E���)g��
�'�,䃲,D.t��A�GH�[���;�'�����o�ѱ'cۜl��p1�'`��3��<'��r�)$i6(	��'>y���h�� ��`�:6H!��'4<V�7�A��
O�{B*$��'��	�ӝk$l��u!÷z#ʴ��'Z6-o��A��zEN[�{�}��'^>�r�
���ҍ��!;�u��'�D��diH�}�	q�Cϡ��q�'� y��&S�"��dSS��3�41
�'^��+q(R�yFA�]�X� �s
�'�R523�ٯC|�2��'"���'v����/�hiA�j�3n;P8�
��� ��sUl��R� �����#�"O���W�ݦm�%�Z��U"OB8btӊ3��6*Y�y�l�"O��	�ō�!0F���B�>�N�#�"O��D	F?Wi��2͖3T��U�g"O��cF�A	v'�,3E��p��B�'#�;���k26L�F�͉.� @�'�,Qp�L��0��ʐNB�i|j�8�'SZ���C'3��k�ae>p0�'N��9���Eh��'�\����'p.58m��i0���k������'��|cV`���$Lo$y�:���'���@�7Y����#�;gV��'��੷�ؘQ˴�k�~$��Q�'��)����8�#�hf63�'Ȏ�ҥmP>��l l�<j����
�'Z6��V@
�y2���m��jD��
�'�^��5
T�}��;��*f���
�'�t _Ņ۶1��@���H��B䉛���V6}|1A/&֨B�	�	<������#�L��cX C�I:C $]���_�>���΁T}^C�+�ܑ���& @<eΚ�wC�I�*�x�9dM�~��P��0H�B䉃,�%s*�W{"\�+��%�dB�	):��P�#��KD�Ytd��TR�C�	6Pޅ��d��8l�sj�>&@C�ɯ`�`���[(h8$P�E�7N�rB�I�7�V�PR�z��E!j�#�C䉘!z��� h[�]���+��C�ɞ7䄸�([�1	�����S�,��C�I4]��:��BA�hH�FЅeO�C�I��)Kf�&��v�[*(ӰC�	{�mP��-F�؛�H��9ެC�Ɂ`�@ç#�p��M��ٙK��C�ɣAg�]@unM�maT)
�mW; BC��.��#�Y5�.q�5��+t�B��7|���lI�jY[B L�'�dB�ɱ8���` �/0v$�CE
T�NB�I(��+��ޑM��%�#��0�&B�I4S�+�AN܎Y���/	B�	�o0�9��M�PA~��%S�c��C�'v{b,m 	5E�T�ui�#l��ȓF���@�S9d�2l26IP�[5(���a`�\ʥ`�@ΡX�E��u)"ɇȓFk�r�@�T��l�0� ��$�H��RO�Z����G.��X$��L(���@��˷$e�%�ȓ(�} ��v"�1
�i��uO���ȓVY����ȏ�@����f(ò9#`لȓ|>�/YU�<Ȳ����G"��@�QoM����"	(�P�ȓG��8J�aڍ]��z��������ȓǔQ�ªߍ�Az�g\�9���Z�!p RO�d
׭���쩄ȓ� a�jʘG��	��� ����H`��J,b9`��v��Q�$�ȓp�Z\P��T�|NYBK��R< ,��f�@�ruꘛf� ��W!D�x��d�e����x���U�sIp��v�IQS�b��[S�B�/��X��
*�{��9j����UA����!,�[�L6,o�\�bM�#B����ȓp��]��EV�=�hY��@!zl�M��S�? B���>6�戙�F*7.��1�"O`�I��K�~� i����=��2"O�r��:eI�K�.b]��"O���Ӊ��(����	C�{,�{�"O��9Eˎ�SJ���4 8"O��I0�ڶ{bL1�EU�`hȺ�"O.�s�-��kod���eA`	��"O�`�@D��i�©o46�j�"O�����I&!�Nؙp���eY�!.�y�M�1&��#,t%I!%��y2kF�h%��
P>�1P�T�y�NK�5��f1c	YU���y����M�IvFB(X�%ۧ��y��T��Eݢ\)�w�C�y���Mzj�@��݈`� \7�а�y��E�Dp}
�̍�"-B�����yR���9
��� &��*�U.���yRFW�vf�d)a�V�EaE���y�m�4��B��mH�Ԫ�Aό�yR�C�|(� �-p.1	*��y���E#>L��ĉ��&��R��yBaֆO�a�ER�	T�/I:�y���r$	�A [�	�ʩ����8�y�%�#�� ���� �`�J��yR�ʂ/�h� Δs�d+P�A+�y2Aj5���t�LqB��y��:E1L�؃��v"���kY1�yr*��GŴq�5�Հ[��8��ӱ�y�X	~r剣�r���֭��6� C�	�R�HU��o���zx9�l\�S�:C�I4g8f�Ȇݤ\N@C@��?kvZB�	�L5��)%�T^�H�e/��B�ɫ~	��s������w�$*�B��?l	�Y!6)	�D1��;��\�]�B��&dLri��H�)x��N\$xJ�B�2b�|�F�J�༑�V$}��B��	,� m9V���x�hN�L�JB�ɡ-L���4a��L�P�M�\��B�	 Z��S'D�I�>ȡ�@K_�B�I��<lר�Zq�R�n�`B�	fǸP���Y��Z�O�.�<C�	�{�����dL&�Z8��*{�C�	9�PXr��-�J5�&C�M~�B�I����t��3o�,�*�X$&ORB�I�xd<*��X��E�3�?F9�B�ɠ7�l�ī�t���p�ԿE��B�I3-=���s�L5C	쑁�mތJa�B�	�P6���&+���10�#�NB�1�ZX�Q曌l*`ڕI���TB�:MJ\d��v��f]�Y� *�L#D��8���5 �$'۬Y��c�B#D�t���Ԛl<������W��0!D�\�e�9Z�\}�O��N��Й��:D�������=ˢaS�(u���ʴf8D�(R��
Hd98TE��6
��0�7D�@"�^�r\r���OW�e�v d�(D�@R�DB
��#�۬`��=	3�$D��@Kڛ`�u���M.6�ܝX2m#D��Bq�Q4}ZV�!Tl�2�	"D� @B��$O���$ɉ1 ��Yg?D��yǪ�O�R�Hcf����%�1D��!Ѕ7P��}	d��y�^ݛЯ9D�zG�%�*N��%�WɼC�ɗY$X�y��΁-
ʘ��-����C�)� "����H3P*��e&_�M�N��"O���Q���I�b]��뜪W����E"O�����`Ƹ�x�*�{��`�"O��#/@"NMP�"!H��p1:DȤ"O��A�*D܌pK�'�<"��"��'f-���		�
��UAߧ+�ո!π�OvС���D1B�t#~�5��K�t���T�"kPlJ� @W�Mh�J�l9�������K �Z騩�Q�D�Q�Lh�D��94�
����OL����6L�l�K���1�0|��!T �PxkPJ!c��UY�M::@�(�7$�:6)%���	� )��P�5�������D�qѲ��kH�XB�b�)�ȟ��Oࠜ��#Q�<�:����Ѥi3��.��h8�����OI�&̀�0|Bg.�8^8����T�2�0�R1�^�t�p���۞l|BQ"S(�R�Q�}n�?7��H ��(S��yr͛>
��âI˄��:�!�'־�L��,�a�TC�z(x��a��d�>��@�46٨��§[$�@6��\O �	ç`���#c"W�����OB/?�� �)N�2'p�R�(/1�&���J^H>�z��]�b���(����L�BW(Iޑ"��"KhI� 픞
*v��hc>��3�ȯ{�4#+)�t��:���'�i�d��r�.������aH�1��R!s@����Al��4��i�T"t.ȣR�9��m�_>U�%�Y(�"���M�L��`O�Z�*��.>�7��)ZY �S�L<�F�E!d�ܔ;��^>z�j4�R�<�G��<)_��k Ӟ#��X` ��J�<aՈ�^�\���	kc��L�<	��8$�st�]�P�N�-J�<���V��a��L�j��gg�C�<�t�ď]��= ��J\���.�C�<i�dR=>iV܀�H�~��0���~�<�F�ʼkԞ��^h��$��x�<�[��8@,��UH1�C���ݰD�ȓl�扂��=B2����j �hJ����[�4�
@���B��8�.]+�$��3�.��'CC�vi h	�]��S6��K�Ňm�$M��!A'x	`���+-Z2�I�Jb���散N��������� !㔼�7�#|�`���W,��m�N��@�kI�[7*��ȓa?Vh��*A� ����5X�2����C~�Y�mЁ>�N¤d�<P���ȓ%�$��B-ٹ16�M�ա٠w0��e�`�:��&6�B����5��؇�d�fd%*B�� ]jg�Q�YE������h:f*á5~Qґ�Z�N͇�/� ��\!hq�Ӡ>/kh0��"/�4��	�6j����Ud�6<o4���Mt�0�W�<x�<�E�W�sL���!Q���͢F����7��W$����2�����ˋn��T&�
C�N��ȓ���e�P<
��Ҡ�9Q� �ȓV�����ٕ���"`Cƅ�ȓbW�ISM]�J�0@��Ӂ_��Ї�	$R��Щ��zY�Ѹ��=�d��@/����b�JA�Y��!��,�ȓeK<e9�AK>L��0)�J4s-���ȓ-�d5��B����I3&H��GH�%�&�3#?�#WI�	�����6��Q�o�.Ĭ�ۆ��o�Ʌ�5�D��-Y�q���@e�)e�>�ȓ)���A�#��[���%;��m�ȓ)�qA�H�(	if�+��#2(܄�)�L�8���x��b�Z����F���%��d|��3 |�,������2��0S�`�b���cl,`�ȓDĄD�%j��hr:1�a�	<d�q�ȓ8��LSg��A[:�C O���~�ȓl�bP��&W���C��
���S�? �X���31���zf�A�)��[�"Oj�p�k�&jΤ�����tYA"O~q�D�zd`tGĿ���`�"O,lk!���:���[��4D!��""OX @B��%K6G�=��d*�"OtC�ѝ=�E0agϧ5�0�@"O��3��CPx��fL4}��p�"O��STo�5V�mȷ�ݲS� 8��"OvM�d*�3^��B�P�4�<1d"O���Qǔ17@@DA3Hγ'�.��V"O�Uϙ y����[�	����7"O ����FU�����YX㐴�"O2��t䞘\w��RrH����qS"O& (�$?G��{��LX�x�"OrP:���+/���;�F��:�����"O�胵��	z신��/p�K�"O���:)P���
\��P��"OP܁�قzpA��85 H��"OV-
QၓE1 !*�@�{Lܩ�"Oxx��G̼!
q.�hDQ�"O:x����QѶ0�1�JCI���5"O��B� �6lN�pHQ�O�G� ��"O����үQ��ɫ��[�����fT��E{��7 B"e�	ι,q)7�W�e�!�L�]���ҥ_�2$j�j�0�!�D�*C�h�G��wOHQ��*��J�!��α$M0|"�hK�|> j%�L�&_!���t��4�Fюmɀ�Q�zA!�$ �=�@AZ )�!m&���GP�j�!�$��wz�1�
ĕx�.T���\�!�!��c�Y"�f�.�Y�w��)|�!�$�4sr�"R �$��y�ë(T�!��B;p$Xq@�^�	O���jB�'�!�dX�̔�٧b��F��s��]!�2�t��!@ذ��vNۜge!�dO��-/}�9rC��5[D �Jp"O1R��*8�B�� �gV
A�C"O.�BfO8�D�P��U*4nJ�q"OtH�������EhΆjް��"Oz��6˦OCȐ*r�.u����T"O�1i������E�?4״�ʗ"O��C�,��15\py�$�?����"O޵�u�ǟ9�����;0�֍�D"Ol����e,���.t~�h2"OČ��B%�j(����a~���"O8��^"&j���K^�
�y"O��c3՗���
QL�l��"O�mF�L;V���jd"X�tl�R"O�Ó*˿7�B!Y����;�,��"Ox�jr&N�t�Vp�í�>N �1"O`���O?�i*q�a�Y��"O��3CF����hE��ؐ�'"O�u��ʯ&�&���j�-�h(S"O�=��F܄n!B�C�kO[��|��"O��(��j���� d@.Ġ�#�"O�X�&IߠH�8s�.I��aU"O�<�L��5)�P
i{R�D"O0�q��	�^�DX)�eP20��m�"O���#��7�"�ڶ˃%5_���u"O<-C�#Ԯ,"�5USENT�v"Ol�a;�@Գ�\�@O��"O����M�U*��R�6E@��"O�B"�Y2�΍B�-[<���"O��"�(��(���ê;8�2q"O� ����ĝJ켘��EѡPjR��"O�	�ސ����ą(Fc���`"OΝ�5@.rb�l(N)Jfp�"O0 8E�	Q"jy����&0D|��"O��F��j"�D�Ү�i�x��"O�����%^Hx��|\N%�%"O�}bqOF>������39�}A"OF���DR�"�M��΢m3Rh[&"Ol��oL�}�-�c� e� h#�"O�����-V�V�a�䗥D���Q"OVp06��i0\��ID8<m\���"O�A1���]`���v(��1�aib"O�����X�7�������N��b"O�͙�-�}�`+B��A���D"O<0`6��A.��tሔ��DR�"OB��N._#r�b�.�>O�1r"O ���ThJ���Q.Υz�؉��"OМ2� �7Q�I+3�Nx�@��!"O�@��ß�`�,����N� ��}(�"Oe�1'U�v6��pB�=Oֈ��"O�T�$	�	}ؤ,�áG�A�x4p"O�YX�,]�\aR�=D~<��"O���gLA��\3��P�|q�e"O����aC��q���%�Z"O\ܡ���#\,}K�HU	X��\{�"O���jǢ4�%��!O���G"O(ܪ���!]����UJ��@"O���f��\Y��Ɉ{@�}�3"O�� W��;��򏊗'���e"O�@�d�ʮHIB��Phƪd��`�"OLdH��ǔP����F�ϒɸ"Oj��5�[�����@�&���p�"O�q۪
�Ҭ��$ѕO���"O����� ����!��ڃ~��"ORA���B�XZQ䏠!輜y�"O6�{EB�&
���Y6�7�v�pA"O���ш�?cL�Z$%B�A�Bո7"O�U�`d'�XD�7b�< ٠0��"O���2b�$�Ԣ�D��2�"Op:2+E<g>$�p`Q�<�^�c�"O�l���%7�hc'�0xu8�"O�A��D�k�HY�r�� ���"O�e[��U�e[��!CL\�	N�,q"O�m��B�.��	�:P;d=�"O6��W�o����V�"*3Ёô"O5�G��ra��G��t�0�0`"O���B9:K��,�/�<��D"Op�1��.n��3m�5z���e"O�ɹ�
]�s.�2��݇p�ppI�"O|u�e@2{~��J��?���"O�-"�	�lh��d��n���d"Of����M[��hKLwZ�2�"OY�'�[
J�4-��L�V{�M`"O|�0 ��gEp�F,��v�E	"O\�:pE�fS��l��wFl�Y�"O��p�ɛ>��}r�jN@. B�"Obu��jT�.�Z�)I1M�\�d"O�� "a��E������
�v8""O�u�Q��;o��1�@jv:���"Of}j�"F���ۗ��S�T1u"OHP��3R�Z�uϋ;Gߪ-S*O$)j�g��y�&x@�!ǐ8���'0�����:_�5�%�]|.�"�'lX8���� <�c��;˄y��� |����1X`�")Św\�`{`"OL��`:Cor�*�?l&j��V"O���Ď�[���p �^�����"O�Y�P�X�%�`JN��|��3"O�!��K7W\�;2	ۥ6�JU"O��@&@!Y����4�R,��Ib"O�ų2��f�1hM-*Ϻ��"O~�0�G�+B$�BFL>�D}!�"O`ѡ2��<7�D�QwDنq��\�"O�,h���R�k�C�ZH�s2"Oh9#E$v�` G� dT��E"Oj��&gКottJq�	�Cb�,0�"O!"B
Z�\�ɺ�h��4�(�a`"OZe��X��K �֦a��u)�"O�H���	�c2�����!x�|(�"O,�����J���Ge��z���aA"O����2}�Qxv�Z00����"O��X%g��U�d�Ǐ"S��-I6"O��P,��c~�xk��Me��3�"O�(�Ċ[�d��l���[
��a"O�e�F�[r�8:��U�B⵩"O���N7*ߖY#&ֶM�r�E"OJ؈vf��kֺ1��$�(�xf"O$Q��U�g�P���ٰ_���"1"O�@�u$�-Iޥc���-b��B$"O��x�.��?�4�M�=��m�D"O� K�'�X�b4��\�B� �ʕ"Ob�wd[9^� �X>�x|�A"Oʁ 7-�7}j`��#����0"O�Q)���aެ#��i�+���yr&��Do4	j�&[y�!��&���y�Ð,�A���-aFj�t���y��g��ɂ�PPKPh!<�2���'o��ctX!a��#�Ǆ*=_^*�'�z��   ���        �  d   �+  q6  wA  �K  U  �`  �h  o  qu  �{  ��  @�  ��  Ɣ  �  J�  ��  Э  �  Q�  ��  ��  ;�  ��  ��  	�  <�  ��  /�  o�  + $ g � 1  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b��<�ߓ#d��t	H*"F��9S�U�ȓO�����0U���6�*hU��zЀ�L^4�z�׈�/Ae��?�-O,�=�Q�A�
�b��҆��Й�I���yR��)'��S��ı>v&�c �&�y��ܞߌ )0Ֆh�]�G	$�hOb��I!k��̹�0Q�A��
��u"Ovm�� ��q��&@?1�,B!�'�ў��s�\�=����M�2��l�$g1D�L��םC���@#
\��0�$G;��hO�Ӕ���N�\�jpT���{-�C�	�3Ľac�tX<1צ;f�c����I	)��p�C�w�l�:�ʄWg�B� /-��b]�c$���bD=_��ʓ�0?	�#])m̕H��S��20Q�X�<1a�D9�%���ѽipfH�Ѩ�<���9{���2���2r&�#��G2��''`"=��g�����P2�Q�eB�yrGäw7��b��"A��$��Φ�yB��$����F��h�t,�=g��!C�NP37$6Ʌ�M����;�|�3E�s�4$��W�<9@됻0� �S�%@�=>��g�Wx��FxR�
r���K�w�X}���m�J��\؟�k�U�W�� �$!��J$D�X5�f��x%�)�T�Jtf�4Lڴ����
�\>@�ȓ<,�dKNO*�$Kr�ֳUY(�'�<!���#X�j�K2��4W:�"P�Y�\7�C�7*M���]7���$��,m�B�I6�$QC��N�s�ڄ
�+G�r	tB�)� Nu���\.N��cHF�y��![�"OV��E�R6L��-�!�� �"O�HX����mZ%/�R4��P`"Oֽ
w��4B������~�x��D�>I���P&P��4SC�@�l��ɪf��*�~���OD�ԨKX	�U P��fV� g]j�<��&L�8Y�� G����f�f�<)@��C��г�+�����rN�j�' �y/�9&ߠ��e��2EE��pv�����e��(����Ej�;Z̹�g�N��-d"O� 9P�+V�d�B��P�6v�K%�'X�R��?�"(��gć[G�m�@C��S�!�O��кצ�c+�|XG�� ��
����Bu�ӺK�yBʗ)`ZD|�b��	�Ą����&��ޟ �?�B�Hի-�9�%K�:��/�)���O<,��I�:�n�[f��8J2��L'd�(M$� nZN*��O����V=Z�� 3ac��,�Ex�MN*	9����'��5@��j�D�FA���y�g˼<q��d�(61O"�P��7?c�3U%�,�:'"Oj�XW�0Z��*掃%ub�Xƞ|¼ii��>���lF�<Y��"]�9����:D���W��21��Z��s\�A{���O<�Iʦu�'�axfP�P����)D+3�>�16H�y2�	X�1r$ֳ&VJH:�/��y����h��,M���)�y�0������?�2��f���y�ߝRtn�I���8;�i�(��y��T=���C�*a�TrT��y�`������֏��5���rb�N1�O*U��IEh:��g��6:���J�,h�*C�	� g�()Ar�����EndjB�I�Bf|��� �&	�����ך@�
C�ɲq���M׮T~�l�!��L��B�	a�Ŋg�ɻ~��4�lQ�)��O��=�}
qD
�#LRHC��JL����HJ�<��-�C��@���jG�]ҁ�QH�<ٓ� ��P�{c��D��R�-�G�<�J!>�4�槛-l��	�!�K�<�tj����΃,y��Q1l�M����?wN��d~��4G_(����B�r�'�ўʧyN���@f��S��Qzw^Ѡ<��%�b�:3�K�m[�E��O�V	�ȓX�֨k3KFQ	z������K����?!�Z+ta�aJ��1hN؋m/�h��!x<5�D�Y�O���z�fճJ���ow؞�&�x����5^�J��&�_�0g|q�s�%D� �S	 �+D�	�E�H'�R9�R�!�~����a]�	ʢ	�%ސ�����5Y߉'(ўb?��6j_�>(N8�����lU@�H:D��(��� �|� �ʧ�pX�� 5D�����ҿ]�j�(�ɌQ����`4D����d��Z��Y��	A�>����0D�г���o�ȁBB��6� V�,�����'�B���U�X�X8�s'ʡ�m�ȓzp�L饆%WLJ� t�Z�a���Dy��#�S��G����E��E��I($�W��y�B���6�J`퐁"
���� �y���(I5�x�c֊/B��跥�"��It���O�ȫ�-O%O�nD�q���4t�O,���8d:,
�8Hwj�q��Ì4�!򤐘�6�BƁ=`��d�X��a|=O>�+n���ЁR�MI|�YR��A�*ғStax�jПm�UXM("��p�+ğ�'*�I�<��I\�1|dݑwo	�%,����+�!�� n@����� x����
&'N� �]��'�`��Id�N��U �u��i���O�~C��(��a#4 ��]��"J��	ey"�Il�ɋo7pI
Fc��mz�$A!#��B䉡[�h�rw��&�h�BŅ:��B䉋r4�3U��.���ǹłC�	!%5X�5�9�@���#w42C�	>?H�a��f�4�X��#p��=q�A[r�kS"�}��
�%�N�)�ȓ:�օ1T-X�ǀ �1���P&��'��}䘶ZN@������vqp�L2�O�#*QG
-� �Ɓƺ`/B�7�:T�<
 �� �H�X5O� ~\�Dh�0D��j��'^�f��(9=&�x�)b��G{��)�)��D�46Ba��E�qO6���y��i�,ɚv�pmq��{��Jx�$�vlZ� ȍ`��0Wl\A��/���E{���^�G�ڬK�dZ;��H�4&k ���S�t���aD�9F�t��׊ۀ0v�$�dE{����D�'d$\ui_�'"��-F�'�ўb>�C��<X��[��ٽ�`H��*�	az��E�f�牜�Qg�I���$�O�\�剾)��t0D�����H.O8���Φ1�6�� �x�#!��RA�E��-�HOh�G{�w>4�����9J
���!�X��
���yb;an���t�K�I�(� m��y�d�>X`�8C��^BB������y�J�E���5�ڟ��� �.^r�r��%�)��t1T�X�s�ڱ��� �;z�
�(;D�L�ЈJ;8d2�p�Y(�f��w&y���<�O�$�$�V;:�H�u�L�(�!���'��+�l�`hS+ �t��#*Иu	����	H≚(��av��<U����D�?VC�ɋ��q�	j"���<E�B��$%��P�1aJ5#�>ɀbퟴZE�B�� �p�C��
}�([?��B�ɴuKڠ��-�	g��P���%7@C䉔�V�?�a M�_W,DX�'�6ٙ��6�����Ȏe�0`3	�'/��0n�=?�Z�C��N(�vt��'��	�k�0s�X���W�QJX��'@d��i��[����a�ӰB�V��'���uG�9\t�L+B.�)Z�ŀ�'m�a�4� �<Yq�B�<&��M!
�'2L��Y$w Q ��I��&��'�v�$l��*�����':�i���x�� ����\�@8�
�'r���Ђ\>$����f��Q���
�''�H��	H�Q���a�� ;
�'ږ��m̀Uk��2�ǒYl(I	�'�8��*��0<����B:he����'т`�V��d>�e���([֘�'Kl��c���ZL�`c`@�9vG����'2
���K��L��!��8K�'X.�c,�pF�%�e� ���q�'&�#O&��lJ`�D�~0�AJ
�'��X���<8�FH��Y���
�':"$J1�O�}{$9�R
�+m,��'7D��bM�'�*b��[Y���'�D�J�a@�8x�؂�کNe�=@�'�n1�Ԇ� qx���F� Hr��A�'��q�/�*x�T�Z�Uz���'�����kf)q푴<�f,��'�4X���;�����\#7J��
��� ���n�?>�H	�J�as@Y(�"O�arA�\�,&yc��Xб�"O�I�h��+�pi�"�l~Z�H�"OԜCgi�9��pE��0~Ab�"O�3��^t�1葊�.p����'�b�'���'E��'VB�'/�'�:��Ga�0i3r0y��]<Y��C�'3��'���'A�'��'t��'f6YRV��+�)a�)N���k��'��'�r�'p"�'w2�'Z2�'�����G0F�8tLݨn� ��'$��'�2�'S�'r��'�B�'ZPK[i��dp#�P	REFTȟ���ߟ�����ޟ��	П8�I˟$H��Η�q�E�V� ��P��h�ȟ�����H�I���ß�����	ğ<�e�V�����`� �h��#��͟d��֟�������	�X�I�d�	ڟ���Y�d#v�Ic�ZY��Xş��I�t�IğL�	��Ɵ���ȟt��Xg"���� O�PL3#�ɟ��	����Iɟ�����������I��p�E�H�1�0�~EPq(���H��ٟ��	şp��������l�I��p3Dឿ/�<�k#�W�ke�u+fW�����h�	����	�0����\����<�'��J�:�RSX�Z��aC������I�(�I����џ����H�I�4I��8J�
�8*I���Y3f�Οp�	֟��	ݟ��I�l���M���?����g��=�g+�-8k6��$p��ퟨ�����$I���i[iD��Z�DԹgzѷ��hA�\��Of�o�F��|��M�� �dz^��r�O1ph�5���P���'�=3G$����䘞mL�����_<�XA��"2N��] �c��	@y"�S=T,$�3a�@?~������u��r�4h&��<���T�r��.�Q��cl�>Z�ȱK�/`؂-����������'�0u�|S�'���j�%��(7 8Y�`��9�����'A2ɰ"�O^ՙ��i>a��g��Da��s�d��l�:,�l�	Ty�|bA}�T�S�J�?ۺ(�1�ؗX����t�ښw��t�(O��kӲ�	E}B��,F���� ��A��H�a�� ���BS�5���J� 1��-��J' j�DԵ=J�SA_=7�FAӥ���}�F˓���O?牕<��ٰ.� 'fF�!4�[��版�M��^H~�`�F���*#���)5��B6�k��	ܟLmZ��`�#�x�]�F�0 ��WB�9�ٴ,J�4(ޘ	�B2eų*Fv�RQ��{�8=����$*OnL"��,Y�a��"�B��g��6~}:�%ؖ�<l�� ��1k�	\�M z�X2Mͻnd(8��g	���zd�<�|��$�.Ud0Ȱ*['�?T�؍&8��zp�c��(�▵E��� bc�-5���p�X�|6V	��)�6�R K�%h&���Y���3�Дr�����a��
� �CA�� ������D�Ms.�`O08���݂^��{ud�������C����}�S )l�H��W.��o��	�%���p���-�$(ګN(6m�O����O�	�@~R��V�,�ɗ�@�m�T������M.O
�j��i>A�O"�خ~�jd�Q�ʶ~�/�M[QI-��'�b�'����<��O�@Ȕ��&(p�8��k�̍�@즁��CKn��|�<��U��e���:%�(�@F#úc��ث��i��'�2G��|'r�'K�ğ��m���cf��F��x��$ʴc�\�I'����� &>)�Iܟ�ɵ(jHY�Ń�͉B�D�OHU�3�iQ�jP�C��O��D�Or�Ok�"*|��`P��u;��9A\���Z��b�������ay��$���K�|+�p ǈ3f9��3�L;�I'�4�'"`@�ӌN�k%1`B�k��Q+e����'��'���''��)UTΊm��Iq#U16�$q�gH��6��<�����?����Xja�ɦ�@���	T�x��^:2��9�q��>���?�����<W���'>��t4����5$���P�WF���M����������nݱOH�3��!1S�E�/ʶ2�x�v�i_�'?B�'W�\S��'c��'f2�OkfaQT��[HH#�\�_I�H�s
3�$�O��D؃�����T?Ѻ]#L��!h���[�P���pӀ�gȀ��ix
�'�?Q��/S���)���Θ*�H�k3�\�6��<Y�,�[���O����E�>�v�+��i���Iզ� i�՟����4�	�?�'��S}y� ���E$�-c�♡s'���4^�M`Tg�L�S�O���ޮd��6�����z�@�u3`6��O���O��Dn�̦q�I�������V�|���Y/0;�+���,����	ß;�����):���?	��f� !S󍔨|	d��c������h�ib�'�9��6��O6�d�O8��RY�D�O�5�����`L����O����S�i��m�fl �yr�'w��O�r�'�b�'�����ٸ..I�ӌI�,TP�� )Q�7��Ov���Ob�$Hs�D\���	3y�~�I��Ë;��@����'X`�I�l����ğ���ޟ���Jy���r��瓤|�"��#�co2��EjS!�^7ͺ<q������O����O�n�<�a,����q쓢Rr��ƶj����'�'�B]��Iw�P�����O���T$��7j�`!�6{I��  ���!��Iy��'f��'�5��'RB�'�rš CJu��t�gA��3kܵq"���u ��'�ɣ��i���>�D�O�I���@��3.��/ֈ��E5P���'�R�')"ް�y\�XS��S�  ���	CO�ҡɺkǄ9aսi���9%"�9 ޴�?����?�'{��i�5:P�غcWء����D�J�Dx�����O`1��2O��O��>�c�Ae�9���ɴo �hgw�� �ȗ����	����?�O ʓ	(B�Ǚ�$p*P�]A���iY}�'rQ��*��	�Գ��<P`��0&�S#[���s��i ��'�"C�.u7-�O����O����O�NT�h� ���Y���6�^�Wx���'q�n݀�,�������R�$�O�Ѳ�G@�
s2l	�kؼ<�8"�(���)�I�M+f�ߴ�?y���?�����t?��C>�I����Lz*}xe�Z�K���#&d��Ijy��'���'�b�'c���$�ҩV��`HB�6<���*���K�*7��O��$�O��DYe��R�����l�:�u��<R�@l2��'A�tr�Lu����柔���4�	}����
-u�7��O��	!Q�T.6܈7�7k�|�m�����ޟ������'{�^���OH�bw�� %�	�7�5��ٮk�6��O����O�D�U�d��07m�O��䏹�k"�VqM��I勊� �.\nɟ���ߟ��'%�c-����'��n/"��s]�7_Xi�gj�W����':��'�"ǋ�4X6��O����O���ً\�������.n(]��IP%�Z�l�����'��#�2���ߴ��4���C��`��@;m.`��`V��M#��?����/]���'�b�'����O��eůx�	��C��	�i
"Dp��?Qc$J��?J>ͧ������ G��F�i�@�ɈP��7�2/�tEn�֟p�������?m������I���� 4���\U��c�M�z*��4{���{���?I*O��)�)�O��YP����ҡl�@�Z�(�-ĪToZΟ\�	���`dY'�ē�?����~���GvZ�!�f��Wj5�6A��'�V�y��'�B�'k18�儨U^l�4ꑷ�B,�� vӺ�d��X��0&�d��֟,%���/l���*�=~��h:Ы3F�*�C�<�<���?�����'.L��, D�`��Ô�̄���T�Ɵ�����Fy���a�وdG�^A��	�$'P��y��yr�'�2�'w��p�^Y��O0��!�f�0� D�Lt�%��O����OO��q��Y�'�H��jвgM�aK�!��Q��O��$�O����<���D?
�O�,�&�%����@(r���� �x���D:�d�<��b�.p��v�zmC�&~_�o�ʟ\�	oy₌��r� �D��0谐n�|�h1H�'��h<�`�N]m�	py!F�O�Ӗ%a��Β5q��=��V�27�<��ģ��f,�~"����v������G��;�Z�K}�8�#�qӢ�&��Fx����� �0�C�$h#:e@`��1�M��+��y���'"�'���� ���OJhh��v��!I0���<���#vl�٦��3�S�O�R���I$(�sHЩi��U��"*Aä6�O���O���hAT������J?�&AO3����_Јc��Q�7��Y�>Ѵ��d��?���?�ӌN�G��1
c���~̋��5;#���'��|4;���Oj�d>��Ɣ���ʅpI��rt-�>I�|]�Q�T�bF8�I��	�L�'�{R Qnh��".�yxcG+`�&OX���O�OZʓ6�~�a���,qZ�@�U}���4.MK��?i��?i)O�qӅg�|z*�����HC�}�� a'��P}��'�b�|�\�AQŧ>����S��L8@���lh,��EMB}�'�"�'i�	Ym�IH|:��	3���B �I ��!�B�M��f�'(�'��	�[o~b�$�3��$\¾Hy�k
&6��|�T�D�O|�DF�����t�'��4�M�`�u�Ǔ||*	BE�L�T�|O����Dx�� �!cۋh��:0��˄��M++O�Ȱ�]���Ȩ������J��',v\� �\-���+��8e,��b�4���@�b?�K7F�^�n�Af����"��s�$�
1�ͦi����,���?�I<A�#��Y҆�M��A0b޽dc��#�iM�5ۊ����`i�ț.�|���*�\��`J���M����?���T��u0e�x��')b�OB��#�X�B�����`�z))���	0<O �D�Ob�d�O����O>����	!Lmc%��+؊tzRDӦi��=���bM<���?�L>�133J�!t(�-5@���5��F���'\��y��|�'R�'��I�h|�y;���%DXj$A�9V��`���ē�?q������J &�ZR�P�D��z�ᗉs6�!���d�O���O
˓u����0���7HW08��@�t)t\���x��'6�'q剗
��<[�
��žX���h�,�TrV|�'2��'G�R�l�����'8�-�@�ۮ7(\؋���U���i��|�[��:ւ6��d��;3�53���'�ɂl)z6-�O�D�<�+CFD�O�B�OD�8���΋�h��Hbf��$�#�<�dIK��������3G���e}���BM'mn7m�O���B�MP4dl�ȟ�O��$M#?��mG�P��Yp���`��g�@��'�Jdʌ��IW���"�$2�q ��^��F�R9p�^6��O��$�O`�)
K�	���@`)n�Pm�#��K��+�����M�`Do��?�g��?�� nkaŏ�ARE��B�d~��;�i:��'��c_$q�Oh���O��d��x�4pQ��Փ�J�$�ڰ�>!ą{��?����?A�@
�Gll��Uk��T���!%����'J`���/=���O����O$��C��ʾ8���CoW4p�epw�E}ΐ�'K�'��\����OV�ɚK�ށ;d]���+�z��H<����?IL>�(O��c��������;�LIB��r�1O.���O���<�cm�:kK��F*���#
5L�|aRraփ�Iğ`��Z�	DyR�!���d�R��Ա^O*1ţ�'���îO����Oh��<����&r��O��-���;j�
�(�2� ��e�2�D&�ĳ<��ns�Y>�0�
ߠ~ 	2(Ź �z�o�̟h�Idybe+�d�T�D��~��
��'���yC#V,r��`�ƅ~�	ly2�΀�O�S�/�F�X�kB�mݖИ��n��7�<���>����~����ד�T;���%Ÿ�	7F�A��(�h}���ʱEx����7$�����+%g��RU��9�MSԬ�<��F�'�"�'~��3���O�!AW- �b% �E'R:r#�%��n���8E #�S�OS��]츍�3�A�F�u{���G�"7-�O��D�O@� �d��џ��G?�T�Tӊ�WaҹU�tаnAi�y��<����?	��d�×�B�x�~���ɴj�Ja ��i�R��3ZRc����M�i����qp0�PF�� 7I�ø>i�lX��?����?�)O���)M�Y��y��oԉm���Y����)�B��>��������/~����ɀd"�
K0IO����d�O���O��s��:��a;R@S�#ژ*��SREl�Pb�xR�'��'�	�b��N@�Y�K�$jX}:��Ɔ_��'y�'o�\�p����ħPu��A�K���eu��`�����B�|yR���'�~-�JCMN�)"� Z!P�1�4�?!����H�f��Q&>�	�?��O����AGo�;qÔ<�Ç��ē���*V��_��x�E�
�DTöf^cb�l�ryB�*24�6��I���'��į-?��J�9�XL"�ٰt�BPQ �ݦQ�'dD��������+j]R�D�*$�^��WY/
�� S1L��6-�O����O�)KS��ן<X����R�6��cH1C�I"���M[ũ�E������G)f)��1E�kF�JC'[�ffIn������t��$͞�ē�?����~2�кGMX`Z�H�>c&��g!ɡ��'�v-�y��'�b�'�M��
E2���Pd�=5ut��f&b�R�d�1$��&����⟸$���*�蘉��
2bd˓HV6�2��F��<��?y����1_g�	@���#�:�0��1
�9p��A@�I���K�	qy�`Cz�)���-<P��wdC�uTȤ�yB�'��'���T��:�OGФc���Z`�[%�8`�O����Oj�O�ʓ#�bu�'3L컀�_�<&$Ai�+9�)!�O���OF�d�<�Ƅ	�P�O�.��g�+R�nI�L�)V9~([�q�L��9�$�<�4.v�s���a�铟D-R!F�G�A�:�mZן,�	Jy��zp�K|����b'��\�>��'�2,/�91�lP�'Y�I�
�"<�O�hD#�J��&�l�ف Q''�`]K�4��$"<�B4m���)�O��)�S~�ȡh������
�ꨱ��Б�M3,O�-jU�)��ڔ����J�v)$ y��3Ef6�9m�~Um�̟���ǟ������?�����W��[t �;)6Lh�EV�
�VH�j��O���O�\�a�8]��QSa�W�n7 LA�,���������	�~p�e�O<����?I�9��r��X��FQ�%��� T0d��Y�C1O��d�Ol���;�ɡ֪�b�JP�TI�T��Xl��D��kV��ē�?����?I*OkҲR�V��r���U+r\����]���: c���I֟T�	fy���.:R���(U�{�"��W�a��"L%���OD�D�O˓�?�U��������,��A�w�ۇS�p�VGf̓�?����?�*O^e�0i�?�0'�qw�ii�Ø�P�D�>����?�O>�+OΤ�U*���]����'R�'2��C�@A���Iԟt�	�p�'�n�����gJ �&MbS�?z�԰"�hm&7-�OJ�O�ʓf���{r��	_�:�����(+\I���M���?y.O<�� �Yo��h��_](�k׮�Ls��A�	h�0�cK<1���?9���?N>�O�pMش�����D�cO�(	�4��D�5Akvo����	�O,�i�q~�Ό�$d�u���Ef8���O��M���?!Àކ�?1K>	��ĭ�2�d�����Bi*�#gl��M[��_�e����'���'��4�3��O���̅�u�8H�Z!eQR  �.�̦5�"�3�S�OD�X?^�Q�	E�4��JҥQ�46-�O����OXm��*NF���4�IX?��BW�%~@:���p��y+�Fئ�&����,{��'�?!���?��hτ.�<���������:L����'&���U�1��O���<��ƈH��/�*^Wb�	r��7[��2VZ�d�bBП��'���'Z�V���� �%��:6�,�b�(Y.����#c�'2"�'W�'32�'��D 	R<���.^D6ĪT⁬{�S�x��ϟ��	Ny�B�5M��ӎP���y"̡��٢��5��듪?�����?��wN���lz�-!��Յ=�>�a�?R���\���	@�Imy��R�ʪ�p���<$���h�� �.d�wF�Ǧ��I{��ڟ��� Ms�c�Thv��3'4�ܠ� �@��u�`���D�Oʓ
��f���'A�t��fJl��$��.򐐷�5U5�O2�D�OXL���	M�dm�HI�#�`���%�Ӧ��'rڜ��"d�^1�O�b�O�D�,��S#�TDQÈ	E���g�
���O������O�O��
�(C�_':x*p�"$C(�j,:F�i��1��mo�:�$�O��D��H�%���R��8�*�#�&\�Q��X��1ݴ4�:����S�Oar�P�S�d-П�L�[w	J���7m�O����O(�G{���IK?)��ف3�J<�5��5�57�u�&�P]�N>���?��g\�r��o����B��h���b�i�2��'^�nO��D�Ob�OkLP1�,��sكD
6��#��G��	��(��fy��'rB�'�� }
���b	���`C��¬L�R��[�ē�?	�����?�Uwr�8����S���e�X�AFar�H��?)�Od�#�Kރ���L����&?��f�:Lp�U�Я� �v|a��<D��X�c��
��)�r����?�ɝs;|IÕ�ǐ��(#d U�w}ja��B�3R�@\� IN����)Ab�jo 0�5c ;52�In[�8N��� 8n_�`�`DE�*�Nh�d�V��C�d!Zl��HM�g_�1qE)ݎqIb���eL�����6D��Y�꽸��J |8�+�F'W=Z�X&�E#�=�3�� �J�dS�gȴhL�=�Y2���0����Od���FQ>D8摢 ��Qf�(m�7�uw�_";��S'v����&c|#��ή
d�'ȱ�ČjyT���HO-m$��eݭjr#v-�%���!9-�ᳱG�)Qj�'u\D���?���i�O�J!)̳��Ļ�)Y�\2�-��"O:���M�[�MZ1)[��Ȁ��'��#=Is�r<��c/�H,���޺9ƛV�'���'�d�W#�����'�R��y��R�R���ZB�
�j��[��
tG������n�nA��;�%�3�DB*��`@�j�Z:��*2��<��,E=�����ߩ�DC0����|��	��$t���r2ჵA��e�WF$6�JyB��!�?�'���r/�jj@�e[4��i���6�y�&t��e�S	�d`��/˼��D�y�'�n6��O0��V���!P�7�F4A�eD�y���	��V��ߟ$����h�I�u��'b6��P��^�Z>q�!�N�:�����>��!�:*���K/<O���L06�6��Ɗל
A��&l��
�bb�7Jɺ}��B5<O�b�B�1@��TH�K�C���៘k��'0ў��?!A��9U1Ze�#h��Z�J7	�r�<U��+:\� ��}�.�3�oe�5�	ny��Qj��?�m-x\�0 �@1(�	��HТ�?�Q���?�O�Y"��N�=xn����S
8�v�r�Ȅ)�@�`2�3O@TzF-�9Ɍ8k7E��N�8�����5p'�[C?hҔҮ0b��9ӏ��(O&�T�'�\����B�v�,13"ρ"��m��+�I@��pB�	��5S/�TN��рj)����4���!K؜Z��9V��<e9�͓��D�� ����'i2_>Y:r�Iϟ�PI�f�xY[�@ǽ%)�z����D��1Lo�`:Q^�D��%{����'��I׷k`rTCY-P6�3+��0��sÈ�P�`�JA�U�%��Ob�V�ʉ7��y�W�: ��23�I�r�
L�>�UfRӟ$�ܴ.}�>�ӬUl�$��
�9���3�ᖒbsИ��,I���C���3���!b��&�t��ቡ�HO!X�k���X�$ա��40�m�ΦU�I͟h�	<b N��� �ǟ��I��ɣ�u�Ә �2��c��!|Z��g A2C��E`�i�<	�i��0����|&�ܛ֏��<�y��ȝW��2�5I��M[*O���D����� ����V�`e�u�%A��Ȗh��i:�˓��P�)��O0�$�Oa�K�0q���`��\�@�wJ84��k� ނP���k�@@�q3f) ��3?� �)�)O�����٭0ܨw钮)8��R�	����ș���O��d�O��D��S��?��Ou���dq=�}�P#�R���S��3n@�Y��՞T��iĥ�0<)��@�)(L��b&��aRi�`C��q�z���Ǚ 
ʬ%��8Sy��P�'r�8;ӧ�Kd�-��L6��́D�G��?1P�i�|O,�d�O���2EF�I�a���9h�15O(D����N�(�0q��'@�	[��*�I�M���D	/r�F�nZ��L! ��@�JVH�A�^�v��ߟ4 `Ƅן ���|�bI�7f���B�W)'j� �ߴ��d���L�]<�9�&$�r.^x���&
�I��枍(��u��Ѭ5m�Iz�^�<�D�:G�v<ᡧ8.��#>A�kS�\��|y
� ��"�j��A-2�KE�Π0�js=O����O��"|����ʀ�*=�T�Xэ]<Q�i�^�)q'Dg���d��

� !��'C�I�*��C�4�?9������i��d[`Ŕ���I�L�Q�j˕\`��D�O�j��<p�xܡ p��\*EO�|�*����D���Պ'�|�f��V�>1W©جU�T�Fa0��%Pc��_f��Тe�3.��q1�I�:�ѥOtX3�'�7��O��+�	�Or�f,ք)C�9�V�ƨ]V岐K�Oj���Oz�D6<O~@B�L͓/�qSD�Db�abG�'�`#=Q �O�����ՎZYq�ՈCJ�V�'B��'�� ���X:�'�b�'
�֝?d���S���9)���1�-X��ty�Elܬ�r��!��v����C��'@�ZE��z��г,�d�A�T-��<�%� �r4@�'\�c�1��I���>q�4`�%ij󤀖F^���u
�==����Ŏ�1K�mڤ��D�/������?�6�F]�s��~�D͑2���T��`�	�'=�]JR͙�a����Q�
�h����O��Fz��O�T���B��8B�<X�T���|��Hr���8�n��Go�Ɵ<��ӟ��I��uw�'�2�D�+f!ȣrr-3@ ��8̚G���0
��ۺ q��X�O�yr$ 蒧Ÿ�(O� ����)F�Rp���϶%��@(7���,ub-&�	�~K<�z�n�ߦAx�°e�Q�C�jɔq�l�&��2 �I{5�E;������C޴��'�c?!u�S�^�`���C76y�{t)'D� (ǋ�U�8��Q��+b%n9J� (�	�M{���<����'+���3̌�P��h)$��-����'c���V�'��:�L�t��\���&��>�慊�m�y4�L�|�!���F8�:צ�8�]u�+Klp���(I�?�s��[3sW��s7�X6��x����?a�i,�7��O�AW�B#k�q��D�=�ye�<������&q�%�Q�V���:8��˲O،oz�!�����2*j �I�a��ly��,d�7��O����|�f*͛�?q��Q*(n^p(��@�B��p	����?���J��ਗ,AjX�a��0/	*�@�'6�Q�fL�*]hT@�Z�h8vA�OV���+�)Z��l�0�S">�N�{Fm��3��Oz��`���
�q��lKxY�H���@�O&�n���M����O���d�%G<�k@lN�fE�ӊy"�'h�y��F�w�88��D"p��"N�0�0<93�I�S� 	3��
��D�f.ֱW8�1u���I����e�l�9�	��`�	ȟ�9]w���G%�ԩ�LL�l3�A;!Ӆ8�#�OЀ���ZŅ�~1�bOH�Ȣ�ɟ[��<�hY4I�\j�lI�<\D����)d�N�X����0�q��O�@�"ɷV9�)"���(*�͢�I����.O�IQ!�����O��O *n�(C*�Dfեy� ³"O|�kr�� ��<��E�잱[撟,����?��'k0�1���TTe���8~�T���#�)P"(�(E�'��'.b�OB�'��ֱj
p�i�ጒk	^����]'gG�qcO��V�B�I�ydND (+�r3J�<X�hx����q��ȅ퉍O��}� $�}Ԝ�ඊ�!�6y�4'�OZ1l+�M������O<�Ш�#֤,�`�����x7��#��Ih<�*\=#�&ݩV�Mb���^���v^�vdy�n�A�p��U�H�I `�Q�`ڎ%�^���Eۏ3���	���J�����I�|J&V%}�p���Ҕ�^YBuh��w��P�UA�Y�, ��S��I[���!5���A�X�6�uBhܼ���H�E�!R	X��ោzn�z��#��]�H)���I󟴻aE�k������ЄCuu�eKyy��'>�O>�`'��(J�\�)��N<Aۦ�+�l<�4��4v}�Ԉr�u���Ss!�4�����D�i�ztl��<��o�4�U+s�R	Ͱ,�
�{��ڌ}��X�5Ôs���'i$}Ѥ
�%lT�8$.A,�
Yڑ �~�)������˓��1K�nͮ�]z��>1����Muڠ�7*��X�P��دTq���҅jL7y.)I.��ym���>Y��̟��ش���'��l<)�]� �J�̂S��b�$�O�O����O&�}�9�1B�".����t��tؼD����M#5�i�K{���D�+^��#��4kCb8Ю��
���d�O���³`r �ЂTE]X�'��F�!���q*n\��GX*���P"+�!��9O~�Y0�T':%n�9�閚G�!�Q�58��+f3�L9Q��,!�]z"��q��:z�"��'1!��*x��TSt ؒpN��4�.�!��;&��uhG�L'��ujq�M�{�!���+Ա�'_#
� A�/J�!��T!A߰�9T��B�������)�!�� �D�U���Zw<�K�DQ���B�"O�����2�R,zf��L����"O5Jʗ�#N
���+�4q7"OH"�N7G����0 �lb$E��"Oi$��FB��!��O�N` �a�"O�=[���|6�۔�R�Y_�(�"O�]��1�f ��Z/��`�"O��Շ�STp��%v���i�"O��e.�5$�|]�o��-��iu"O���O�k��q2�0d�5��"O:��$/
"/��퓕��]o|���"O�	�&��T�v\x�� R�m�T"O*i�&Ŋ4$�Դ
B�rԹ{p"O���Ҁ?g�Jɳ$f_�����"O�5�M�7�n��.D�`�fM#"O������%#�q�\=����"O:�[&��P3�i�bQ�m�i#a"O��Y���1n6f���bJ��潩�"OҠ`5H��kL�IC+]$uʱ�R"OD�7Κ-H��y'Kצ!�ȉf"O Lq5�O�$�,�A��5�<� "O���oɄ#4,Z���vl8P��"OL���-�/5h`�{��I�}��A9��D>���>�v�/�)���sӨ�����I=x}
4I�=l�n�B��J�+0�ЋǇ ��֝�;X���@a�Y�_�^����E�!��X���%?k�����)ӎ#�T�AGB�\�(���VV��O�A�������1T=I�r`�p�x�k$p��8F$�f鑈��~�L� ��O������J�
N�k �AĆ�3�>͒r"��6lT������:7��i�2�h��V�8�O�OL��1������B	�"냉��i�SHJ!�d|2�Ǒ�S�FtP��'�	�s�}��I@|��I՟@ܡ:���(O�ӎUs�4�cy��$�� �1���Z1/]yF ��CXB�����q^��ݳ(o�$�Sm�_�z���x�Y��'�ў"}��.�$
����`E�IUl��OV�^�Ȩ��ˋ	�n�ɚ<b�٨�/}"e�(v�,��ЮG4K ly� J����$2�9HEh�+�@6�T!��%i[F��UJ�R��%w�*��e���<)qDO�1G,A���N68�ꁳQBo�IV~��W��yE��A�z���H�'�?q�D�$8�@��+4x0� �r�'C�H�����!�� ]�G^Ap5,�t(<���Bk�HU0��&X�ҕ�C�L�i�.���D%s��iDzZw0��)��P��y���^��2KY�?|�$R�`���Pxr�-:NI��.B�P ��'�Q'I�H5�>i�A�9C B�H�B�:���|�ɷb�.��c�&OߴL����JF��{<|�6�J"K�*H����
�a:�b��N^�S%L�5�d!���c�v����B�(RWD&,O@a�6⎄w�(�@b��b�PL�&�>Q���#E����ElTFݓ�&�z�%�(qW���V�j 0�W
:��S�O���L܂?�:����i��H�u�]�iM�,���,���<��?)�I�q>Q�B�u�D��BУ����
O�)"�/?BN�+�3.# ���I���'�� ku,T�����1V('�FZO<��V:�b�+ص)��ݣf�$�'�I;_��`�#ȕiY�ܡb˔m~h<P�+I�(�t �ㆲv�T-��<扒6T,���#E;�U��gQ'R�n�D5?���AK@�c�s 8(r����P(�V�@�8�3\OP� `�8-:@yb��)x�
�U.B�젃ת�g�h�ʕ�'Nў擁%�:�a�!;�ƱkS��u���L���+���d�6J"n8K!	5\ �Z���$zT"�i>I�GKwyBm�
��LbS�Qn<rX�p�9HE~|0��	6a�I.+��@;�دO�®\�UvDՓ��=/���D�ȼ�˓�?q�k���DDy�Za���O�\�t��
{"H���撦B��J��0o��!�!�T(I�.h�'��xIa	/i$��@�j9��i���(�`o*|����f�% ��l�'(�hp��O��~�����Gy��W�)G(`VJ~���10��3�xĚv��<�S�ǭP?R�r�#�=b΀(3��S1<\
�1�)Ug�2�E|B�	0%�^q(�w9RmI@OܪM0���6)$B^p ���hO�>�ؖh�c�$�cb��i@�dK�M��X���0C�$"GpH��*�S�˒�+?�T8؊��W�,.?�Ha� n}R��]�'X�T�n��Ic�(@�
Q&AGx~����8D^HC$J�P�Ur�>��|�G�"$�S�'�y�	���,�K5�Ypъ��I�OjE���y��!e
ɢ=���� ��z�E�=4x�ʍ!f'�eї@N���'z�Gy��������+(DR]�IK�h(��'Ȋ-�ȸ�F,�q�"=�;DD�RD��HS��?#���Ң�	� x�E�O��=E���Hk"Ha8�#U 1�,J�#_#~((Fy�J�+�H`:�+E q[-H�+O>���+v�&��l��B��Š��,`A�˓�OX�@��_.qbQ�ag�`n\�)2a�8G�����&�ci�̹'�\/61��>N�209��ڼ;���`k�9�'r�	2���SCA���˥�ٳf3^��Q�|��������<i2�YpQ���+B�!l�\�$���(����0��D{�O�4Ѫ(�3o&B$k'��)f%��D�j=�b*T��HO�N
�L9H�7ﰔ)Ed�W�MX�/Գa5q�0�'�ў"}*W���7#��1�E��4���Y-K�c��kRÂ�-ލ:$
�(;�$)�@:񤎁`�^0�C���ު�����+^��I>:��0���B^������i�
��҈;l,�υ$E.��v
�ik.�����!x\I U��,'�@�?%?����Ư�hHb\k�:×�)}2� �\V^t*�'M37x���-��'�|�
a���Àڴ��
�G�>�O�i�㓗4��8#MH4FGf�h��ψH�pyKg�ީsR�Eapl�k��j��ߨp��F3:��E�p���9�)�5� �i0�C�����%�F���H���m��G���Y#�dD���HЅڵY�������'�I����"3h	�IG�4@�4�ck��y2���tU���T>���A=[k }�b@���Bi�ToT��G;7��p�'�Xy�ր�w�S�O~r�����=���Q%)7p������[���~&�x��.�rٺ�,� �i��%�dIA�6��
�6�08!c�%�Kt@�
T8� �3B������[�j �B��S��Y":�{�D���p<	A�_9Hrf�O䰻&j��Mk6�ғN:	�pI����lX����hO�p�!@��Mx��[��' ������S�%˞y�b�S�c���Q85�Zp�'�ɔ%�_�S�O. ��7�D'~Q�Q�n�z=�a���G�^f0X�~&�$[�ǚX(4	�u(W�/@�u���A?Qa'`�$���3r��K�.	-<��3��"$e\=!#�dj�1���i�5�c�=���]�<^dl!���.Im��Ⳬٵ4�E��M�6����@�3/�u%��CZ�P)t�C7�$D*]n��raߜx֔J$J,)��'Kd���\j�l��C�H�*�"�'`�QQb�ԟ@��W�tZ&�$*�晪��=���Ơ��T�]��`��Z������-�Z�IQ� ��?�G��� &��A�H���ɑ�m���O���M�w[�	D�X7p���24��ؘ}VA偏�0`�ib�L�2[��GxRn�q��$��O %���!�J�r)�%��@v	@�AZJ����aQ��)�e8�B�wsdm���W�d�b��Su��es���U�her3C>�'�D�9&���<�x Ȇd+-��H҅�(�I4	:cwD�u���B���4�'�H#�(�� $��.\�H`��J�$B�2A�I���T;�d����x�Ё�95�h�B��>��8rD	�;k3���S�Ŧs3���2��,~�Zm83� �~-�'5�I�cx��@p� # X�4�J	�*;��?dwp�6��
#��2�B��Q�+ԥHJ�0�k!�!���*�S���`�'�ڈ�b�O�犸��'������}U�1���`�4U�wA!Z;�i�S�#�HO�}@�h��7�}�U�ޅaH�@ �-8u���'E�	�����ڋg��u��ێ"+E+";\\��HO-)����}R�P*7`��F��<�qsE��%��r6nIy�\5P�a��t�ȩ /T2C���QȽ���FJ�?��S�Tq�\ޠ�P�LG� բ��jՓn�8�aD�]� �P�P%Z..V<�B�>D�D	� %}J~
�9�����hսq�"Q�櫕_vf��	Ǯ^���Z5+{��SF�{3��؀kG�'c~����d� H'f�Z��49� I� d�nevFx¥�n~2I,lڶ(���R�9ʛ���mR2k2퓯t�~�	��Hh�n��"-C�fS>�HC��~���X,�yg��E4���sf�̀�P1�?Y�O��2a`��1���0>6�b?�@�`Z:?pA�E	[�a���e�`�t�?1r���.S���B
XB
G��O���jl�QH��B�>p�L��׳J��D"� t����^;�=��4��PJīR�~��M��σz����N�9/�:Y�`�E>9�N�Pb�����񖤃5�~r�2C~�**O̽�#O�OʓJi����(a�n�#pn��H�����6z��S��f/f���`e�йRo-�2�`�s	�d�%��ٽ1�v� 7'Vy��$w��� r�,� ~��6o�=���1ta�.d�I9v�"-���өu��@�)��#�Q�(�6���x�$�2e|���o��M:��!E�b�Ҙ�xxA�0`���$���_>�LR�A�|�o��Fc�q(S��+���bVK��`�,��ڒ ���@0���]��~©ܪk�t����/At�h��H�gC:��4O.cn�RTA���Uy4�{��Ѕ�Ҫ<T�'uYq�id��vU+�&�ˠ��)� ��y��
�i6!�C��<-�PD�VeR��?��O���UT��S���M��ѣ�i��vы�NJ�*�g��6w���dH� {b�iV�֊$|>�s�H��u_�U
�{"���(W̤�i�� �����
�y��V2"�@�L�0� �鑞֝�$�R�0�Io�!�P�(���&J.#:l�s..�p`�8}������2#��EI�Ä7رOR�2��Ec�<r��SK����x�*��o��""n���*�bȽ�p<�G����L����awֹH#�>6��Wܶ}s���h�f������el˞y���	�B+3ay2�0�0j���<����ȓ���	|�����	�;�F�0��>M����p���k"�1�P+5��!Ȥ��,ϐx�gD$y����eA�fR�.��D��oT9`���uA���&����]��yW�9�De���0�Tda1����Pxʌ'h�� 1*��?�a�㔥uq�`�?��&�8l��i�EjD4]�~��r�I�$	 .)aÚ'�� �aP%2Ò �b.�Z��?eWʖ~N8"E,Ӏ
�$��M~6�9YIe��9��E�J���'�D��rL�����VI���VS�b~B$ �D8�� Y)Q��:�0�?Q�@��m���P�ȍS[� �A,n�'����٨�����,ّ:XfUu��p�' qO�=�e�~J2O�eP����A*a�ՁM�ds�S�;�ĠDzZwB
ͩ)�"�yǉ�!s.��ĮG���-	�?1�{���"J��>�9`&�&vE�y!�_��,��7�k��O��Cp�ʅD���L&<�R��@�x�.u(��c��
� ��!J	P���"�{�1O�)��y��R�,����5�h9��a?_ibuItkӽ "�QԂ�>����.F�76�	&
,�)���f��Ҁ�{�.t�]ˣ�w��&B�蝹�O�-.^��2��yX��H�Q��8{��"�"zf�������'8�U��%��تD�%�f��t!�EŎP �e��
��!Sfg�j���p)�<E��]i�ԥp�	�4b��ze�ԗ~&T��BM*����`y3�yܐ�R�� �Zi:��O'���b �#Nr&�!������!@:0=`rʜ�`� ���L�Q^���''�b�>�.O�Ӕ'B����]1��n#.�JmB��Ѥ'	�	��$�@�<!V���R���Θ$^r� �Re�<��ME�9zȌ�B$#C��0�ǅx�<!��=hn�����C��h��H�<)�� w���z5	�_�R0�EhC�<w�5[��rAFS�ĺ��Ǩ~�<q�`ؕ^4��b��5O�!7��N�<�L�k9JQ��J�l��P�B�R�<a�&K&?���	CM֢]d@���̙Y�<I�M�)(�,+��g:�XPg%o�<�2܏R�tI�u �G!�	��m�<����6{�@X��"621f�n�<чk� C*h:���%
 ���D�<��n�`���L�ёU
ED�<�4!\!!��d,�2,B�-H�}�B�2V%A�C�o�8s�ҵR�B�I�zF�Pc��؞D�fʌY�B䉅T`���π0�����T#fB�I4 �d�"$gܫ�0���ϖa�B��3U����R�E���r��̎��B�	)[�nTYE̟�\��� 
V��B�		:w*�p��}�U�d+K(i�C�I����畿���Q��N�,l�B�'M�6A;���7PpI*�A2g
�B䉬$O�E��a#,u� �p�B��	z�M��&� d�V���@�$VL�C�ɽ]��I�Q	3Ӕ��#^�&��C䉖L�d�j�C��
�X����S��C䉗=�dX1↉����m��	�zC�	�[p���͞�L$�0�ꝇ
{nC�I%=OP�X� S�y��)����C8�C�I�<РH6�Z�I�R���!˃8�LC�ɓ6�`Lq��1%i)Vaǌ�LC�I>/T��`��F8O���b�j��|B�I������ &7�j��ϗqFBB�r�H�2�HB6|�E��[(XB�I/<�oƌ2�A���ɕ� P��c��(���n�*��4e�Z=���ȓ �|� �@��	s��`��S�? |!���o�e!W���h@1"O�=���8����gO�c,4�""O����I�μd0��uz��"O~=s���b��cd��e�\�"O�����S��Պ���s�U�"O�&��p ��6m��"O
���LY���A4��Nv�c "OnD!�� )\Z
���m�= [��y�"O$�S�E�F�=�W�\S�A"O:��2�Unc���ݡ6>e2�"Oz<0.w�t�HaG_V#0=`�"O0 �U0S�$�ԣ�#�y��"O��+ì�(hs"�l�h�""O4H��*N�'�� 9�`��>�j�+�"O��b5E�<t&6l����/0����`"O���&hǾ<���B���$�p`"O��g%D.Q�: �f����A��"OX��#;YE��w��8��}"u"OF=����
��z2ĉ�\�2��"O�! �@��S����,N�~��ٰ"OT "R�Z�G,T�ᓷ
�"Ģb"O4�{�a��u����! ^�+t"O`�QlX����e�&���E"Op��畴v{^��-�A�N�� "O��#�/��'.` Rm�YV��z"O|(s@��[�ޜ �T{�b���"O�����޵Bʘ��"��R����"O���4�Jx ��j�&޳�Z%"O�ɋ��X,�X��%��*-V���"O�ej\�z媄k�,�*���"O�C��]/x��K��L~\"��"O�	�W�P�P�2ت�BR|�"��r"O>����{�Q�2b",����"O�ؒ�+�ʰB3�<L��3"O $Hco�6������3y�k�"O&��`�ӄw~�m3g��8�U�"O�Z(3V<��[�DŅv�,B"O~L�V�ܯR��5�dU4d��1�c"O�l�"�: �̕��/��:f"O�$`��N6,��T�'��Q�^��"O��)өC#V~��"�%U��}�"OFy���W@n�B�HЄ+���j�"OD���eZ�`-.�:7�R�w�Ă"OΉ�Q���>�q���-aV�s""O�9[�+�~�H�;���<gCR�Kw"O���H�S�he� �ߓD`�H�s�'�ў�`���5F��h�S^堈���4D���NX9��YK�j'h����D�1D�@Y7�D�q�h� �h���p�"D��R�F�'�f-�F�K3C����@>D�|Bao�i�x��%��
;�n�J�N8D��x��M/F��My�`�0"f��5D�����S�q#��b@��?Xn6i�E4D���������H3n�r8��%D��Z���҄��4A�j�:�դ0D���d@�V����$��IHƭ�9�O��9��l�&b	�y��3��fL���Y�y�NC�����aDQ�9��(�ȓ?�H@
C�:�v��u�I�}�|y�ȓ5�T�)="d�!$
��E��ȓ��Hq��i�d�#B��T7�q�ȓm`�T���1W�Z��Ei^W*Ȕ'�ў�|��@JД�kP�U�[ ���aAF�<�`��0�陣Mt�"��0�E�<� �!�3�HP��E��#�9J���"O.Q�և�9�U�`C�1Z�""O�P�ÑV�,Q0�#��t�"O*���/۲��G�֙M��q "O�a�®x��R�n
F�J���/D�X`� G� ����k̽0nF\�i*4�0q�5eu���N���,0�b@w�'��&���%�,�cSOѹ@����eߴV�C�IM���b�jM*Y�\�؅�ޓ"��B�I?=XQ�bϭO/t�����ƬB䉄r瘵"0�\�0�Z�苐CQ6⟀��	<a�εI�%��Dy$�r��G�C�z^�*��?y�
��.�$"�|��r�ȱ��V
%����I�J}�ȓ,�" �łM�}ex1"1'�o�N`��)����U�M�w\�!��-�& �������B ��1%pj1[�m�j��T��v��m�&[�n���� K�d�ȓ2���i!f�3p�8슱@�΄�ȓG��KU-E_�6��5LB�d�n����f���W�=��\Z2@�x�D��MܓjvV�ыu:�	����0����l��n�Tb�,x6�T�D��ͅȓ)<F�pvd��8Y����Ad��ȓz�]�H.4�1yǅH�
�5��:�<H*���V�b]� ��E�f�ȓnЉh��ް-��]zS䕕T�R ��.���JD��4�����'$�}��U+��x��� ��EͣAȔD�ȓb�d�@��p�����̠J�2�ȓR���3��d=�����T ��@��v��
�#C�>�Q�Em�uji�ȓ9�r�"dƄ6�"�R'H����ȓ^��8C%l��U�!�P&,a�)�ȓq�!�v��<Nl��Ȓ�v�x��� ���#�E&[��ݓ��W�	��WYL=3�S�w�J���n��蜰��6nJ11�i�!=���a�^1d���"��L�4J" lc�"�Ua8�ȓ@Eb	��HR9S�J$� F�O�!Ey�'#����k!Sp�3�h�҈:
�'��Q��%�������TH�'��y[��V�<��y��@�;oȘ�S�'���j`�";�D����;�"�'nP�B�Iїu:
�T���"<��'md���U$��Q�nCl4 ��'?`8X��ʪKf� �WAD:d�I�'qy	�`H�!�ۖ�V�xii�'���Q��6bD�f��x*�SL<	�xwR���I۫%��=�@Ȉ&+c^Յ��?��D��q��mpd�E�Pd�j�Y�<d�U�c鸅�I�/zT�HqL�<��I�D�2�����xG,t�E�GJ�<��o�L���	�	��+Z�r���[�<�W+�0>������h�V�P�f@m?	�:�T��M�X�z̈�nR�w��E��D���+7���6c��-U�ތ�ȓ�R5i"ɖvBPqqWb�'(�����q��H�o��I�Pq���+�xGx��)��*�i@T�� F�[w���W�s�<���%T.�Do�]u�����o�<q�I�ot�Q�� �(K2��A%�d�<���
CN�B`,��>p�l �h�u�<ɷA6}W��P��ؠ[�d��TGNt�<� ��rE#mW����/����"O$EI�"��wL"�j��52����"O�|��.+��gO߲�YS"OvX�í�����B��({>�D�O΢=E�d�W�%Ȫ�ࡔ�V�0��7'V��yRCՕ'�yѣ��c�����&�yB���|�X( ��CM�xs1ˑ-�y���'6���'�~�Q�U�ɥ%��B�&$D�����T݈��ˌ5!�B�I� ��rmI<w���i0mK�Y�B䉥`�z�I���n.J�zEO	�,�B�ɒT��2�O�$X�l��H�Ҡ��s�- �h�[�hЉ4h�=ty����A������DY���o������1:���3�]�r�\9C�F��v���1M��:󤆰/����$g�2F5&��F{��t��Z��CR�_�[Z���u��.�y��K.��$ O�@�nB�'!�d�^5R�ҬIU&�F���'�F	;�.�"2`�<+f��Mh��S�'�r��҃�&Z[vy)��=:���'0�,y���#)Yz� �,�0לq��'�>̫%.��I���v�Ž%�h��'� %��!_�:�l$ Չ��Q�Ȼ
�' �Q2#����еO���'«f�(Y\����ո�,q��f8D�4��I)A�mk��5�fu�7\O�b���0!�|A��'%3�,Y�4D����h�6� ��'}��Ja�2D�ة'J[�$d����
+ ��3�a/D��	�"��d�\R����L��x!�TC�^�����]D�m�U�?!�DC�I��d�$n�TP���!�$W�2�fE� ��"�q�S�D<7�!�đ"fО���Gk�N�����(L:!򤚭&���v�V
}���� &!!�$D��dM��Geո���֭0!�D)bٰ��$�G
vל,�f�!ut!���#3�����
�5Cv�؀E�!z!�4W�pq;�\LV
���J1 \!��  ���#�U$| cS��b!�Y�Q �@�Ӿ1�����2[~!�dQ'���1f��m�u�(S'3�!��C� �hQѲ��.<�x@�w�њ!�H?m����Z�?݌Q���`�!򄒓D�(GN�@|"x�E��!�!� �ȑ�B�LP½���޾]�!�dʷp(�����A�IY�v$���!�İU0F,T�v0b����	�5�!��@�PL�ڔ���`Z i���Y�!�$�[���2�g�tmt�z`4j�!���
"[���䃔�R�جYC�G��!��)L0�K��&V���	W@��Cp!�$U�!`t�����*Ĭ^�7n!�� ]��:��A�&�0aK��?!��ڿ6�� �N�:H�P�j�!�&�r��n��� ���E!��Q�}~�طnڠs��e��M!��9p���	�3Ȝ��Z�v�!�D��W�V��WÇ�z�HPZ!�P`\����=���В�ə�!��D8��HѤ���1�rahd���Py�,MX�h��5�Z;P��� ŏ�y�E�|�]Yӫ�4�Za���*�y
� �Q� *KJ�����=4C40 W"OD��4��5%0��'��{�����'6�5�AD�'t ȱP�������'Z�`f(ތo�a�!R�v�4���'����!Q�������gX½��'��Ô��7�>��L�Z��1�'�E��M�A���&�!�ԝ�	�'Ϙ0 i�0hⴓ5�Ӕy���	�'=Z�qC��9!nD�4D~C
H�' ��T��K�tHT@�#Q LZ�'O�)����h���R���.���'����o
%x�u��MW�O��:�'s��i L�;E�0a+�#G�D�,U�
�'��$[�'�%
p���>0����'Mt$��矫Lr}5�:|����'�(y���1 m� S4M�o���H
�'{�H�`S�}.�Q�V�7j����'j(i�5%��Q� ZG*�J�<)b�'�y#&��*q�Q�&��J����'����2oO;k�e��o�(p�"��
�'2��bL�`|�٠+N?Y
�'��*p��;.X&x�C�ʺ�d��'������!���&�]�9����'IΈyӏ�� �:ecp�ǅF��3�'����5,)~�����C�4��'������A`	A�`�����ã�y����%�0tz�'ML h��ͻ�y�o
�j�x��Q��]��)%/A"�y댸IV����ˈG
�D	���y��H(Ĭŋ� �-�^�I%)R�y��_#��S�M�*��(��J$�y�c� d�L[�� �\��I����y"`+vg䩇����A� ݉�yrbX-��0��
W��p���	��y�jKP*��L�b�<pZ�[��y�� 9�n�Ҁ�'b�����$Q;�y��%[�|�q璘a��C�% �y�e�+D�r�X.�v	G_��ybE��qZH��M� ���H���yr@S�Kk�#g)L��u�����ybm��ɣ�U�F,Lݰd�@��y-[S#x	�/F#@�^�2��:�y�G�C��:�(��g��rӌG�yBF�R�&�Ч�Q-����b.ͳ�ybh���:���!���H넢�y�.�;[�lUʇ
��c-<I�%G��y�G�?�f�dO UY$�b5���yr��wV,P�� Pj�=ZE� �yb!ŗ�Ji:�K���2l�����y圞}�,��m��"ӂ�pc���y�A��RS�Ԋc��� ��b`(ȅȓU��zaʔX�hx�Q	][��������b
8
Zx�#u$R���ȓ7��P��L&{�"�Z�?8���ȓ}��rD�/$��j#��!>���ȓ�@!A@�����.6L�R��ȓ@�H��W.�w�0�!KG�1�"��ȓ�v��b�8���fª�,�ȓ^6p�Q'@�k���I� ��%�,D�ao�%9���6��q��`�I+D�4��З�Fd8��A�-���2�4D��S�Ѻ�x��b� gW�䨧2D����Q��]@��9	��-�34D��a���o@&0B�A�y���aF3D�� �8���� IJ�j�j^�YϼYR"O����,	�}�h;���S��$"OL���A�-��t"��ߚT�n���"ODİ6��\��k�D:i�� �"O�� �O�\���X�6�0P@"Oj\��̶1�5´�Zx��G�D�<9u�ñ~�V���7
�Zg"IA�<�Oա(%`����3.HAʅ���<�Kҋf>�-*�j��6�P;�a�G�<A�,M��I�f�	�3�N���A�<ه'W�k�������$$	�D[|�<�4�ݫFl���IP�&i�Ȩ���t�<�C@
����ī�6j�4Ds�+�n�<� e="���SA53��-3�B�o�<a��)*WvA��+�'Hk挋�eEk�<	E�ԵOo�|RBL��)������f�<	%���E�)q��[�K
�(r�J�W�<9��5�0�@)ԃ	h��#BT�<���[�~��lCWK:���q`ϏY�<�B�DQ���`l�: bn&�n�<)E �>,z�E{�H��l�D�<ѓ��;H��t��3<\p�J��<�PI3[7b��4*E${�� �FP�<V�E-	�0�S�T�&��٘��H�<���ޮJ4�)H��Y9Wh(��A�<�� �#��Ah�5.�]�,h�<��N��� 	�s�D1��K�O�<y���}�^���A�/^����Alg�<�h�uQ���6a�+qz�Q�b�<ٰ��a��T�@��Pl��%�\�<��E�tUh�p�J�O��B�$_A�<�S%W *b����%�$Ը���+@�<���Ɇ��#0�F�Zʸ˖K>T���H6������H��q�D,D�` �/��q����/ÝF4�c,D���*Z�b�ȡŋ�*�dA��+D�|y��֨�r(2D�p\�Q2 �+D���G`F�^�<񂃉�)�^�q��4D��!Re8����n�=x\��q)2D�PX2��Bu� ��)H�m0D����dɥp�r%�Ƌ��N��t R�-D��Wlі^������֐C7��3�/D�#�@�i�1��ҳG�����7D�����\<�үTF�r�{�E7D���ԁlm:�K]��!ؓf4D�p0��ϘI�����)x*�i�2D��pe�7z�,(�!]�M����B�$D��#�c� ��T�G-��*ɰ�2w�$D�h��mW'얕�L��o���!c�0D�Ti7�_;2��e�����ڬ`�b�3D�@i�@ܠ�
)�σ�!�n Q�	&D�X�w#����d���d2P&D����nBv��}��d��4��6O$D�0)W̊�;s~�*�]$��'�"D�pۣ
�l� ��N��5�O?D�@k �9T��4q�
�Oij����*D��2n�6X�!��"K�W�.˰�:D�x C�"�m`FKݥ-*m
��:D����54\в�_j.�:D�X�3�I�X#ĝ���\<�F�6D���Άg��� ��c/��F*OJ�"�
��v���Y�%E 	nз"OX�R,�%{E�T@�K�u����"O�Q���ʮd&y��!cI��E��y
� .�Q �8bX�6�H"]����D"O�u�����Y8���j´,�0u"OB`	��E�~�����E	�M0"O@���/�V �e��
;�T��"O
�b��(,$b�A�S�V���"O��0Ƌ�x�Xy备m�l4��"OJ�J��"���M
���3"O���bOqCP\�D�� �H�zr"OdP��iA-I��p(MD+��1�"O<�C�.�K�N8BqJD�s$rhh"O (�SCPq�u2�(5w�@�"O<躴��!�~0 �&����з"O�Hh�ށ�,`Z7��/+LX�"OF��8@��d���.�pEB"O�a��M?U��X�w��S8���"Oz|b�K�E=��d��+,q�-"O� �$����A���8!��;�"O"=���H ���'����Z�B"Oʜ�%}kT�k�(�$pB�"Ovd���K8rBbBn�Pq"a�"OB�����y�-𦬈�ci��0"ORE$Æ'�Z�c!�B,��xr"O�`T�; В����e\�Q�s"O2���oO�IK~Qx���nK�ʗ"OL��LZbfN{ �_�8��p�"O>�x�bT7i@� � �vȚ<��"Of�P���	6���T�/u!���A"OT̑%H @�h�寁��m(�"O\��ǈݓg����AF�9`t�b�"O��0�޻
]������u�>H$"ON@;2l�q���T�z��"O�=P�Z�;�ҝ��	AB��F"O�Uh�KˑKz�8S⫅>w)ĥ��"O�8A���' .i��iӮ(0�ݹA"O:\�C�!q��P�#ÔU(n��"O�q"eH��;����ՌD�t骰"O�H���Z9����B�n|Z"O��H�#�"E�R+��II�<xʴ"OH%)��E�e��@�|z~S"O�D�FX8>%��qr��*1^�|�W"O\X� �Z�#��)��b>t7"O(�
��'�&��e�&3�5Y�"O:�1am�Q���pL��>%fi�7"O���gU.fTj� ��M�)�`��"O�����&�t!��L
�Ȑ�"O(��g�p4C�΀f��Ub�"OA��ː>	N�\( H;p�qC"O�8j�	P":��̒��T�c���v"OD$'��"$r�[��� �9g"O�(����64�Fy:��L8b� kr"O$@C@��b�r�4���*��"O����瘣w�ڌ�1o]�Z�¹�u"O�,Y�^��xH��ٍ��h��"O.HXr�N�c�(9���*d��u�"O���c�D�Q��s4�����G"OFLAEߤ`��ȼM��(�G"O6�)@gB~L�H#ۅ{�4-"O���Ă�"=Z!k",)�ZQ��"O4�2a�E�]�|PS�̋Q���3v"O��� B�k�d�r7fۥn�u"O�ÃE�6� L��Cњ\p@L��"O�D�1k�Ht*�r�5ecv�KA"OBX�Ę#tA� ,�x�@�
�"OF��`�Y^8 �`Ƈ0�6mA"O� `Aʧֿ��baI��W�F���"O�$�$x�	3%
˺}�2��0"O���e��iظJ�G�h*X��"O@9X7̎+'��Y�I3YT�h�"O�a2a���a�䊢'�4��6"O~�3@�}A����6"+C"O�Є $�@i�c��8���c"O�i�s��H�Q��@i	��"Oj�!��K�r�4)�I/n����"O�r�M?�hCϞ�e��
"O$�7�Y"J- �M�Jz�x��"O:8Ǥ˷w�hU�o˺Z�x�G"O�TI��B�pY �O)Z0 �"OFte��}t��Af�+k�}��"Ol$��KZ�^Φ��GE+&i\({�"O�(Cg�Q�:�R��ő6*��v"Oc��	 �*���N�=҅8�"O��c��C+М��F ;�s�"O�a!�*��6!`y$"R�L�]	�"O��o��n-8�`F!}�4Y��"Of@bq�-V��X��%ʄJ�t�"�"O�4�F +qq.LRǯ��a"OrT��H�A�A�C�BtcD�;�"O�YW�H�0�|`���N\�b�"O^�[�d^���A	�&	�"<%�"OP� ��K�t��F�� ͸'"O���E囟\�Q�P�:*��r"Ol ��d�'5���c?HhQɑ"OJ��fCT:9����ÅL_��U*OX�J �+/�����
$��)(�'��(�BӜM��<�%H�-O�0Չ�'�:cG�3pe�\�7��d�1�"O�M��o�.d)�0�V=q봐y�"O�<�̀�10�-R����FB���"O�L�� R�mH��ʤAD&�"O���b��Y����\�%2�t"OJ@˵�*i��-I7��3#8Z5"O���Kߐ����
E+!��"O*t@��ɺ#������@���"O6h��M�9odH.V�]O��"Ou�T-�i��Ӣ�3~`I5"O(,�b&B�����]�G�%2`"O&������(���c�E˳I+(��"O��[�	P�
ݙF�65{R��"O渒�GHH%�A��Cۤ	��P"O> ��_�#Ԑ� e"�D`I:6"O.��#kr ,���նC��`�r"O\��5�ڶZoZ���O�7eO� QV"OT�adܰ2�2��p��JR��"Otb��
3&���988��"O���A@yLQs��4����"ON��N�SLٔ��=0q��"Ot0��A;P��$K�.�$W�}�'"O��x�c����@�\ V�10"O�q�C�@�~p^�0�H8?Q���"Oĭ��'�
y�F��k�8�%"O(��e�QEv��3'��^g+a�T�<��LثbP���c���Ta��LM�<1���{~��HU�Ծa]$�o�T�<���A1(6��H��*ZYD�^P�<! #"1��
6�����8���v�<9Q+��حHTF�0z:l��'��r�<���׳0H�,`T@H�}�Tx�ICI�<��!�����d�� ń]�<� R�#7 Y2d��<+��[:,0P E"O��'�9{�{��"P��<j�"Op�MXqG�t�7~v�(�4"O�-	��K�#$�	+w��L�n8��"O]�efϛShfQ酭�7#p��!"O*�Zao	"���,�!Yl�Y�"O�4h�'T8�Qh���v�0�4"O�@�%�(y�&����0٧"O�h�g-��#2��2����u�F"O�`�^�|�N���j��0�\ES"O
����L�kH*��		�o2j]ap"O���7g˔x*t��ӥ�Mʚ8��"O�ذd���[�X�%��z9a�"O�9�%��?���Ee��G����"O���r��;w�N��F׎s�H}j�"O�9ĬFʒR��+4`@ظmQ4�y�%�$>��}�0��V�H��kR��yj�5	m��Yr�S�졠cdZ�yR��7�>袡'F�Rx�Ub�3�y�iι5� -Q����R[�	�`F��y"Ŗ\���0�
�:C<���)�y��b� 8ڳ �3��;Cٝ�yҫ� "lPԪ�'���а���yR/ɵU��tؠ)��a��"���yr�_�v��!�*�L9���y2����) �7'v�2B!�y)ľ��R+	0�Eh�
��%�P-��'D�ZKهH%�$���!�����'4b:M�T�}��V3���	�'�<�ԡ��r'��e��L� a�'��8(�'��6�ڔ�I�7�>q��'�.}��l���)Х+ް�j�-4D�$���,OS� C��X5n�|�9��1D�X�CgH1V�Ի`�աy�0�c%D���k���3R�?ڮ��#"D��J�I��*9�೅�41[�b��?D�\B#-�1*>��e"��X�b�`<D��j��7:�l{�hM6q�@UK��;D���0H�)�j�Z5�3Gp��c��;D���EN�|��0zcj-_1��r�<D�4� W�7�c ƕ)b5�N;D�L�rn�i���#��ӅF���T$D��yA�:(�m��̑+)A���-D����;���Yg���0[T��s�6D�T
Ӌ��T_�H�A!t�a(��3D�Xi��ׁ�rE��$�Ƭ�p�/D���I;{�i+��\,���8�B.D�|b����p�%Vryx���L9D��Ӷ�V;/��aY��V�jXbd�%�5D�DQ��,XO��a�ŕ�:ZPдl9D�\��� %8��Գ�`<Y"t��4D�h�ρn�x��Ή#1�L���%D���(O3�MB�(.���"]F�<!��]>m���S�D		F�Pk��|�<���˰,�����܃$���<)31��И�܀n�Pc�P�<A�^UB������QR�����x�<!�ǔ>��EA���w��|�0�q�<�2WE��R�A3>aҐȴ�l�<!��I�z���`��ԉq/dQ�D�i�<A�d��z�T�_3D����m�<�d��pʾ1��/��Gs�d��K�i�<aV�Y�,n<� U�E�̐� e�<�j΀K�tP�ʊh��`^�<� 
$��A��PF�ٹ0cRo��ms�"O��*T`Dl�f�ܹ"�`I��"O�2GcU�~�c����su0Hi�"O��ij��J���1�EL+;u���"Od� I�,���:aD�:���S�"O��b�M�0`�ċ���"O*�]|�X�ۡCݳA�P�#q"Ot�YR!F�D�BBC�x�4Q0�"O�=��KU �8�b@9+�꜁"O�IGL�;m��1��%2��a*5"OZ(YG�N�9̠���|�Dy
D"O܁�hP$ �����	ΛI�6d��"O�L�%�
eld��S��7='� W"O��8�K�רT�IA4dܻ"O�A�QKO�d�P�󴮈�+
��ss"O\q*֩΅)��p��kέ	�@�2"OH����ܦ7�t���iB$�
���"O�`��@Z1fG
u˄N��D���"O��P��,g�	w�$ ��G"Oz�SG�!H�e�n
�w(�a�p"O���;ʅ:E��jzv�)�"O ��@��y8�qp�X�rr�`Q�"O��U��N�1e��w���Q�(�Y�<��O�+`z&��'�M+���� \W�<�䨈�L�Z�)F���x����X�<9�j�1������R���3DY�<7�l<��B/Ֆ���"B��O�<)E�1bȝ9�I/xH�A&�U�<'C��%z@�Ȇwz�8y1� Q�<AEڍo}D ���"Ո����DO�<Q@F_�N�Dc�A	�2,�vn�G�<qB�I-�Ճpk�=(�x�ƃ�X�<1�l�u�>(�%�ԎKp�z�j�<ip�z�,�$��n�$l�T�g�<�K]]	:Y�#�"<�ar�`�<	r螞� �CW�E�EF�1���_�<��h�-o���떡�^��I���U�<ie/��fJ�2�L#�hA�$jQ�<i�Ò�T��	��G�~�"���j�K�<!F��3���c�S6W�d���jPG�<��#�lDrD�6�"ﺗ8� B��="�",k��O&q��x��M�2O,�C����J�h�q �΂6j�C䉊+%��Z@��Z|8�(( -|C��!�|��3����'�o�jC�I�U8�e�S�@�a"�@2=TC䉟L�Dd����N��P�r�xC�M���1Ѳ8�%;�b"*�(C��Z>��@�+V|�9�-_�\gHB�I�7s�9H!��W8�s��Le^B�I�0Ϧ��u�s# ����7^B�6KV�Q�E^C�e���Z���B�I�/P�C��ץ}�u0�B�;� B�	5;�dt�V��W_���%�=�ZB�	�"��&	��B2_<B�I<�D`������yyQ�K )J�C�I-a�0S�W&�"}����}s�C�I�1kfaW��4�ss���x�B�ɤ0YH,1�nC,Z�[F�D�T�B�	MT��[$��y��A0$��C�	�)y~��5#Rh��t蟛q��C�I�1��L�V�XrM�0A\w��C�	�m��r$.S�e�V��3��}n�C�)"8y�'M�pI8D�B@��,B�)� �0wH��!ܖ��@��j�l��"ONy9cLz�䍁�oN�:�X|�E"Ōh��ڨ$��"/��	�p���"O�Y�$
=��J�nӜ �XiX�"O����Ċ�TPh��̞Z���p�"O<%��$E'D��8 ��H���
��+D��[p/�;)K8y�C<
�&��׍.D�\��S�Ա���"Gj΀�w�*D����JU/F�ia1���z��$��&D�xI3n�/WDp�M��U1Rx0e�"D�,"��2p�Ua��˓1����"D�Ѓ��I(��Q�ʛI�~�iB�!D��0��0����	�|���kTa4D��+Q�M���xg���_���˴�,D����$HW�P��Ȝ�����m D���`��W�4u����j��b%�?D��r��"2���Re�X���\Xv�<D����H>j�4��-y������;D�p�UF2{���Qs��9����t*9D�����H�<=8�c&�?X�.t�B�*D�����V�$��0� rp
&D���$M ��p�g��Ki�H&o%D�ԫĩ�}��nX;|�,��"D��sH	?YK&��(�1I�t��$!D�d��EG�<ІTq�ԿEAzJD D��"B։���2c�+d5��C�?D���D�	����yEP�T�Z���8D�YP�NG�R@:P��'�Hq��-;D���B�Q&�Yr�^�(�@�e-D�d0#�o6�|j"��6@��X��"'D�,XpIW)I��I ���yܨH�e*D���)yk�IH5���b8�L�F�)D��bqa\}`�D`��Rs��,���&D�@ZejG�6���cb�R=#��sd�%D�41e۪s=�`x��T�t��4�#D����LB���\9�ƒ=zܡc�#D���#�D�.�ђ-	�2���?D��m�1��g�P�| ��C�b�y�<�#.��e"uJ¿L��a�L�<Bȋq�$�8��V2}0�[�KD�<ab�N�+����V%,���*���h�<��aG�;��0A3a%���E�h�<1����N�9c�ɢNl�rf�y�<����O����	�c�B��AL�x�<)Q�8i@h�D��_�h�aRʟ^�<�o���` C%�Β���A�MRD�<�-�Q�N��޴1hl�~�<Aw��)Z�6.�J�hc�{�<i�-!l�l��#\%T��@N�<��K2��+G/&	��:@��A�<�߾l�N��ρ�+%��ҳA�<٠D^��P�e�����
e��<���Y�z]L����&��-��l�P�<�҅E�4�~ ���I�6
��T�u�<نUw����#��D�ī�i�<�`,Ʀi.�PH�bX�l�F��b�]`�<�uE�Qt:��}[h�����^�<�ϫ<6�ʥ���?`ЅR�*Z�<����3h�ԅuFòof0���V�<A$�L�n�Fh���//\�c��T�<�j��ēAkJ�.�xq$nXT�<q�D
*%e���%�)�8"˚S�<����g"$����I"h�d����K�<i5�H�U.N��w�YhJ����P�<� �$S���!'Ҟ�����R�� A3"O� 1.�*�5y�㋽4����"O4 :W傕[��|�Lʵap8�ye"O��̴|�J���J�1_h��"O�9���H`JXH�+��Uw�pBQ"O�q҄��Z�&9q�ʍ(x��0"O��윌oЎ\�v�F6{̉h5"OL�r�		����D�I	Ev�y�w"O�ѣ��(���`Hs6�#u"Oq"��JYL� ���/Bf�YP "O\3���,P5(�$DX�6<��"O��S������������2�sV"O
��dM^��Z���,LR�TH!"O�m��b:�l�;g��\��P�"O��X Ym�\���U��Te@�"O
�֪�Rݴ�k*�*��y*U"O�I�� Lc������ Tvt"O�X{�\�����Ȝ�c�>��"O����Q�ABRr��%��Y[R"O�������{�qp�\�b�v5Q�"OT+�� >{j�8&B��z�*}[`"O�xy�+_'r6幆�$�n���"O�������@��-����"OV1�$�H�sw�9�AO��� �T"Or<����?QJA�3��?��L�"Oz��%!�%\!,���,<30�8�"O� ���՝
7*���� $|%�"O4r��w&T�'M�4Yf�p�"Oh�e���2��a�K4^�t0�"O`H��̓c�]�S�Q䪐j�"O*T �%Kv� �-]'+nҘh7"O��p��}�{�-�k �"OE���)St��l��@��!�"O�,�'�@�!J�lpq����Q:�"O��A��6:^�\g�ȑ��{�"Od��7�YMJzd@�Ľm� �"Oh�8A,�((���Ӗ͍��|Z�"O8�P���lr �!􂘆2k�q�"O�hq�B�EXڽ!�-%U6��$"O4RB��р@��ID|�z
A��yi��!���@��C'��@
�y�Ȉe��L���H�:�RPZ��yX2x��%�b�ʘ�����y�o��H�)��^��Ś�l�"�y�g�[�V4	�I�Y��0�\�y�)v���AE�5V�v$B��F��yr�N7(E蕂�RH�tS�\��y2�C46[�s�1F7�A���Б�yZ��1wh�(W�:E���/N���
�'Yެ�ůJ�#y��c��9U���"
�'�gH�T����MH�# @	�'oB%k5�Gh�؃�3�`�	�'�V�9%��-^�0�!J&>0S	�'�D�`҇�4��H�rꂝ$J�1
�'�\i[�'� a��C2Cްl��)
�'{��Ӕe�$y�R��C���2أ	�'�%k�,l X�BP�>i�i+
�'i^t�W&G��BаA�W�*%���'Sj��!*��dYH��H�rex�Q�'`谘eFgIqp��e�ƴ��'v���W�V�x[xL�
=��!��'΄�[%D�7\��NZ}��1��'�@�3�	�j��X	4�M�?1���'�<ɠ6�Ƕ(s �c��
����
��� ��	��{)��*��ɨY�5�4"O:M�vIG�r��HL�H�g"Or �G.5X�>�S@�O���� �"O�� ӡYlr�A���Lc��hѦ"O�XgGҚpʼ����^�9����"O�Ղ� H=!ˊA��L�58RŲ"O
������l���U E%4X"O6�@3��'n\�30��3�X�A�"Odm�3�ΰb�I��d´���"O��Z�bC+4D:�ؒ���6_h���"O�|15�^x���[�a��B��D��"O�ـ򀂹SX�q�W���l�(\kW"O�U�Q��7L�D�*��2c��j�"O^\���'��d��/��?�Xź�"O�!Z�%ĝ+>�D4�=H��%)�"O����fXD�L�sk�\��"Oܼh�	L>@C�\���� 9B"O��Xd�D
@�F��%u�Ha�"ORT���G>9k2!K�$QR�~8�"O����F�Nq��n��HJuc�"O  ش,W�SK�S�ez��W"Oc���^����ՠ�D��U "O~D�u��)�*4�mI�V
��Ȗ"O��P����)g��w����"O������9�z�Kg�1�j�
$"O:��.�&� ��ף�p���"O>�b�)�� ᓬ)�~�@�"OޅS� �89�X{��j由��"OH�E�:Q|p���В"O:H��]�p�pE�^�K��3"OF,�AM� }xx�&�!ꖅ/�y�Ȇ ���k��W%{� �U(��y�NM<:��=����&#P\����yR�$D�����@ޅ�r	��� �yLP#��I��/�>�  b1��
�y�Ꝝ{���ѵ�>/}J�S���9�yr��6%�"���"1�$*����yb��8��8jT�������y�O:<3XS��[�d�!rAjI��y2D��t�R���l�(��yRoG'#'4e8�F�28���y�g�d�R@7��-S�|���̱�y�N��E=x����Qh�u{ �ا�y���p�P�X��5 �EH��%D�x��I@�"!:]9t� d}��pse)D��PhΖ@�5J����9�v%0��:D� ��/��edX��.}���YG�\�<I$$S6o?ĘreOV4	U���Ɨ~�<y�����p GΎ�r�&i1A]~�<A!`N���2#��'5,!2�w�<хU!a��Q��&n)��@"�Gq�<qw��.bs����ʝ�@Vt�"l�<�G&��f�8Qq����@�#�e�<���J	2� �94�U}���4��_�<9��xz4���K�Q@|�#��X�<��B��2�:��'#N�H�q���T�<� �ެ@�闁��A�CR�<y�bY�#�����D: 3�U��ȇy�<����k�pF!�7P0vH�P�<Ic*9)�~Q�D��N �+%�O�<y"@ӳWZtyB�ˌq6�9����P�<q��ߏqtr&�X$v`�O�K�<ҬE��i���O�B��a�,�K�<�d
���uX-�2WJ�]@�MF�<� FA '�:�6���|��@"O�)D���#�>5{p�G^�0���"O6̘�Lϧn����T6G�x�"O���6ƟF�����R�z�i�"O@��@@�����?(]�"O8@�,�)@�L���;3 V8��"O�0�5H_�/J���˕2>���sF"O�P��
�1"��E��K�L	0�"O��qDL�=�V�5Þ>°�Q�"OR��iȺ" xKgH̓M2�+%"O�8���ġc�:���	M�0х"O4���<@�^1P3b
�u^��"On8�̒G���@b�F��@�"O�	�F���W�|đd�#a붩Q�"O����Q�X(0!eLLN�p�`�"O��a��5�h!pcLԊ$�>$�R"On�5L��vY{�ME�~�Lp�'���h�NO�|��AJĩbBJ���'LVubA�,ِqq�'�9IFH)��'9��@�j�c,T��p"�;�� `�'�\P�'�G�=ۢ���$�:���y
�'�hq��}�`5
v��*�։1�'#�(�Sϊ3�l�)� ΌU��P
�'�Z�IU�E�R�x���S�G��`P�'	x������fn�XA'�*l����'�:����2^�������3��,!�'4��G���/���P"M�x��<@�'[�Ԁ��	T���A ���s�&�q�'r��
#IT�rt9f)l��1�'��L��o�Nl� Q���cUJ�B�'�9u�_1ӄX��	ִ+x��'��JfLѢl{��z�N�!�,���'��L�G>t�@M����'x0C�'�h�0�*Z�vVi`�H�
�����'�8���F�( l�ZDřtF�9�
�'3�u�{����MֹH�b�("O�ux�ʕ���36��3�"�{�"O�V�/>���bt�^-m�U�"ǪS�˩I~�DK�ܙ	���"O�l(�nF�lpxH��N5{�^��"O8��*��D(&}$EW�����"O�	kG� �F�_+5�Y!R"O�A2wE�9T��5!���
��R�"O����*M���m�.��Qr*O^�J�C�ܦ�FM	f���Q�'�����ߤV<��霓]֊,��'�Ce�ٝhEΘ�V-�<Gh�K�'Y� �P}�5A�-_2+y|�
�'t����gC	~L��c�G�OМ�
�'n��K��B+pt��=oFZ�!�8p5 �(�
�*�+E�\ *!�ϟ�~���@�D�l5��F-MP!�Dܝx���!�� ����A��^h��Dͯ���r�$Y!BǸL2�҉�y��*1�(�R�),��D;"�Y&�ygZ%������0���၃�y2	^�n���VnJ�:��咥�y����`	�<Su��q0�G��y�ưmߖ�ᱥ��_)���vjו�y�M�k��A ���L�d�ã���y�B&h;�@r���ru\hD>�yR��!�kd�3Tєp�� � �yaDtx�H2�F
:O(}�S͓��yb�ԫ|���z��&D(���N�!�y
� ±�fφTb��S�D7x�Ӕ"Od]E��ʊh*Ф@�'I���"O�5�4&v��1�M .H,+"O� ��!�#08L��H�@e���"O��eF%Yj�1K�e��sK0t��"OY��&�v,�b��28�˅"O~�!t�
�)Ԑ*C��<
 ��"O�u[g��$�8}RuC_(׌y[C"O ���2W�����ǟv��:�"O@e����D�.��bg�3Z��l��"Or���%��$@��3'JX���"O�L�q��:9�-��Ł�]�I+3"O�dA�/p�%%�=uf0Lrt"O4��#I�L( 8��Y�6IJ�#�"Ol�����8�Δ��G�h��I14"O"�H���(�A	����&/h�Y$"O�-�&�1m�|@�[6�h�$"O$��B�Ͷ���S���L�њ�"O��	��q<E���7+�,��"O��#�#����#��6rI��"Oε��Fe�Y5M��6,*�K�"O$�sE��x��t��688�w"O�p�ꅐf4a@5���dWnP��"O��4�3�KK#]k6�s�j�<�Q䙉!�R��GiP�({��#gIk�<����`�p+��Gf��iÆk�h�<y�d�p]Б�`�G>��DjRo�<1aR�����&5�!Ӧ�V�<�2**)9��rK�-8,I��S�<�Z^��CA�RU�!�hXR�<1����+	
����ȡ>d�d�C��M�<q�$�.R=6����o������Ze�<Y�ᔸ2<.q(񥃽+C�0�5/U{�<��	�@J���7X���8��OC�<q%�$�R��6���`B�PS�<A�ʆ:#DBA��)�Z�����w�<y'J�4�Ua4�n	��Mp�<��d��H�����X">����ƍq�<9�ιd�n��p�@�d]:D	j�<)��݇T5 �-�
MB��
3c�@�<餅��Y����N���x2s�<�b�V�f���AۅMW�YJ5�[n�<��琏\�,�G���j[�tI6�Lk�<��g,B�|)�E��'�NL��l�<	S�й5�sC,�~�Z��B�e�<9�	A''v�@�F	��l�����_�<1gFR43�q�"�1�X���]\�<�lJ4aEAݠlL4�.Y��B�I�%2))�* ��ۆ�Նy��B�ɜ|Df�wF�>aʝ��M���C�ɂ"�
#E�C��M���4F�C�I�PR�E�e�ـ°�K �K��B�A2
%A򯙅OBN����F�k��C�	(VM�P�B�O�4@�-��C�Ɍ+�p�-�K����C BE��C�I�J�P��m��l�Ĵ�vӮ�LC䉩;e��`����x
�S�ʏTxB�ɕ#����h�P�hYPO�{f�B�ɹ^{��J ��!n�0ꀟ58B�.B����5ϊ�t*���g�K9`��B�I�L�\�B��3D6�tjǤ�F"�B䉞/�>}�e&�J��8BA�,;��B�9G���:�`ؘK�(P�#:��B�ɖ���ej��r%"ܴJ�B�)� r9Xp�٪c���$�՘S�h�5"O�Z�B�iC`ͩ7O?@�ν)�"O��`b�[��Sb��K��E�s"O*Y�Ό)UɡSE�Fބ{S"O���o��ts��e��D�t�p�"O��g��H��8�D��u�RUb`"OZ��Ǝ��p�IHĤ]�:�4X�&"OL,� ���k��R$��4L�r�R�"O��)�IT�3���b��,NQ�4�D"O�����(;����p!��/��-�"O$ؑU�1*llC#���;Gp1h�"OVqD`�#p���C�˂D(0E�"OX�ȤZ)։�R\�d�b�"O�1ȷR9��vG+�ĝiA"O��I�F��"I�s�\��(� �'q�q!��b�b*J�l��'�(���Ğ-Kj3��]�?�>��'Y�H����Vô%!#��:����'�BRU�$�*U;�K�;�P��'`��!GE	�|���h�H�^���'� 5�̄�a�ey��_
>9�)�'bXd�R�%$���Ѩ�8
�s�'���I�L�Vܜ���F��E��`�
�'�fq���}�����I&U�X��	�'�ޥ(�g+|����e��T�!�	�'I������:�a���-E��	�'����@sy`eIX�D�ꉩ�'�"|C"�N����
�7`xX;�'<= t��7����DL�6�0I��'{���@���k���P��	�'�˱���!|���7`�	���ȓ'��2BI[�l(��3���.!J��ȓ/lXr5�ߝ_�l	���'��4�ȓN�8�"'}8�! ��g��Յ�9��pB�ZX�q�b8z{Ұ��Rw�!"c'Ń�D���5 &쭅�[)$��ULDtM��2�d��1K��k���%�شT.�Rr)�?zĆȓA��90�"Ŕkp�!q��J�,X~E��fN��:�枒U�.�h��I:�*-�ȓIn�ig�7�Ըa�$��y��)��y�o�h6����љn&P��ȓ5[�$H2��37�$3���e;���Aq���-V�T���fI8"͆ȓoY���Vl�*N�0h|e���ȓj�V �Fƿ!����$Q�l����E���b�Kдag>�A6�`ń�"3܅���؃	}�4�7��I�~i�ȓQX�v��4da�Ѕœ�N�>���n�܍��͐��)��l�87���ȓt���P�GP0����'�f�~ �ȓ<��@�$;��eԁ>�jĆ�7U�P7$G]FL�$@�&�2%��8��,A��;d�32f	��"%�ȓ� ȣe��P�>!��"����ȓ4��.̒ �"�R���H�*���zV�*u �<#r��R�ș)Ƕ��ȓNv���9c���3�X�yٰІ�r�l �Ąn��i�M=�)��8�K4 ��8�<�8g��&x*ͅ�.���Ԧߙ�6�		)�⼅�"?�8�2�\�k���[��z��̅� ��ǙV��,��$���М�FLP"e�,S@@\�'����S�? �܉�g*@�x]����`�U��"O~ذ�FK�\|��P��o^z��f"O��4L�)vW���T���(`)3�"OV,j�V[>~أ���>; 2�Qg"O������=D*�Pp�-h���"O�0$kJ5�)sEL2oE�q�d"Op�Fg �}RP�L6�!r�"O�*^#*�B�N�c�$�#"O X�v�1�0#�'j���h "O6p��@�):5�s�ɹk�r�1`"OR�����nJT  �/g��HS"Olu�!f�].p	�7Ew���c"O~�)¦Y�%h��)]1_]��R1"Op����]!�� �Ϛ3�F��"O�l�Ci�98#xLJ!L�0td�B�"O�,p�N��/2ؒ�
ҊI�;f"O�CǧT(i���	6�["T=����"O���� zX�UL�0x��s"O��C)M__:�
Jk 0�Y�"O^`���%&��l �#q���S�"O�<%k�.
�L�RU56x���"Oּ3p�	�Aޥ����a���r"O
�3쐤Y(\�	��� hP"O� ��kW�W|]��{��LV"O�XЗ��|��c�M�	O�l�#�"Oy����n"R�V&1(�a"P"ON|�����4	�Qחm�j��b"O"��&80���7�m�2 �#"O��3@FR#�Ԫ����3�$Ak�"OL���`\�+_̨#�	:v�И�"O�	����{��h�X�: *֯��yb�[#Q8�i����&;A@����\��yr�A,^�����5��P�Xg��X�'[&�dJʠ��	� �Od|��
�'�D��7O��Xպ&,[I�x�	
�'�
���`t^�v��1ۚ��	�'D �����]}��赹YljP��"O��9e/�.x3	����z�d���"O���`\1A� ��i�a�:�)�"O��Sea��sP��n�?k�BH��"O���Š�#<�΁E���c��Z�"ON}��W�p��n�346(!�v"OX�D�'I��m�M�D*4��q"O�pS�R8a��>Fp���"O�5Yu)J-%�FU�f��A(����"O�՛����B���|��[�"O����Q���2!!��NT�Bs�'@qOf���BE)��i� ��(hl��"OJ��P�?.�hQ[ad܋3N+I�J�<)C�Ԃ`^�l�D�P�4q�.�F��X�'N�q�wO�e^�31G،I$Դ����!,O�D��-m<\1q�q��0R5"O,�@� ��Nײ��w��*t>l�F"O� ��O\�I묬XO��2�,��$�x�'K�z���1�}a��ܢm`d���	�y�$M�3�b���b��1C��H�O��=�OX@�
S ����t���G�`p=�	�'�J�".�t�v����D��Ś
�'V��3at��]��A�t�2�x
�'�ʤCG��S��]a�р��RS�<�g�q��I�dP�U�@*�c��<�v�$ʓ�~����rV~��ƭ	%w��(���C;!�$�!nB4Ԙe��%moh����:%�	a����!��Z�I���h�!�7q�P+�i�/8!�� ظ ���*��d��Z��s�"O01XO��/ �(���C'�$ۢ�	L�O�Ey1�ũX��=d�'��d7O"6�7�OjP��'~�6�`iC�l����"O�1��C�`��u `�@:i�:�
c�i�2�'��4��J�OM�-��Gҋe=,� �'�M��ǝ�7Nr<���_2h�'��d���>?X�٠5F�g�.!`
�'2����I�&V؀��-\"tU�'��d �͇$Th���E=N�~9Z
�'Ƽ�3(V�,�X-�JזA�n1�枟��'ԛ��Y�8�5f�1o��m��'ڬx��8D�t�΂zL������zO��[�o:D�p��U?�$d�P�-kp�ؓ�#\O�b�L��J?r�4�EQ�F�8��*7D� �3A�s8�W#N<R�pYbR�5ʓ�hO�S�5�����V�D�u�'��ko<C�I0}��1��#��y:0�pfF����pE{J?��-��E/��Z��2� 8�4�(D�@Z�%_��@�1���0�^�{4��x�'���D�,O:Q뤍���h��E��>���B���8��?	�$�RX�'L��$&�㡁�0z�ԇȓ;#�����W�Z�B�cRg�6 L�ȓy��#�4lq"�;5�ś{�⨅ȓie���`�z���u���L#܀Ex��>aK~"�'c|,�U`��9���]F��$�*O�����2K�|�q�%S���L U�>��O�'��2�	�|�>ū�GA�sF�	��ψ�B�ɂKZ�q���w�>,ӷ�̣'-��	��?���{��G�6���"���y�o\`TM�$$�2"����n]>�yҧӟ/���a�/��`Y0��4�ēψO b��ᖂ�h�N����jA�y��2D��rD�LҀY�0b�4���� �/D���B�ǳfN����L�0w�+ʓ�hO���)���PGԎ<� 1��'�q%�tD{��Ĭ	&�ii�K1y�X���y��8k$��d&y���aď��y"�ʮ6�L��'��r:TQ��N��~��'�R\�U�-#V��6'�0ꈤ��'�kF@M�1Z6����Q1�'�v`��*�|x-�G׿![|(K�'����HoǾ58��E�g4���}��)�ɟW�.D#�B�H1��J�� Z�!��/qq����Õ�@8�C1!�5!�!�L�8[b���e�� <�tː�S$-�!����(� @
G�E��^�fn!�dľe@�ͪBܝ?��-[��W�Y!�$U�\��Ô)��7�V� $s���	t�'Fj����K��4�TfJ�n��8�'�^�h�gQ!H��e����S� c�'c�T��E�&���s+^=�9H�'�`�(��۶2#$�3��i�B		�'u�2b�\Ȯ��,	>!.�a�������/�O���#�J�>];��Q���ٱ3"O���H�i6X���z^�m!�"O8=�A��.<�"�y5�P:^�<p�;4�����%9|j��(�K{���ta;$��r%��;[)��T�J!���� ��y"@��)e4�� ќ���Y+�HO���}j8 D�RM���D�F��
O�LQ���C�t�{�@�76�� �pX��2#G�/Z��BO�� ��C3�0D�T:�@�x��Q�@�?h|�E(�/D�� �|S爡cX|�iᮊ(+���4�	j̓�O�qR��LrVL��B'���	�'��uj���56GTq���׉��\qӓ��'�1�q��S��|cW�6�� !�'�6 ��4�#vʌ�x��$h�'�½�c�17��Ea�D�vՓ�'M�蟱kx���KڗK�l��L>�����Aj�r
�
M�����̈́�!��?8�N�(�쉞;�2a��/xm!�Č:���&G�)����&��w@!���9J�$���g�x� Fg�E#!���	�
ܘP�K;��L$�K�'	!���`}�S�L�/��i�΃:!��F�q�aP��:x�ܡ�.I�J�铌��-<O��#��"�Μ��յZs��1"�	W��?�'(���P�]�U`4����U�Z�@�ȓP(ڕI�DH�y.�[6ڐFzb�ipў�	 �L�|��6��*E�z���I��!򤗋x<�i��C��� �ÕE��z��1�\m��|"µ��U+E�J���ɒp
��M+G��lp`�Ȁ�Nc�1秊E��;�O�X����0nZ��$ȁ76�@��,�S�d��a�5��n����7+����'dU0��ƻ>ڙ�eڅ�ܜ2�'����D�Lq���=����'�,��7���j���@@A�zej-OF-Gz��	ݸ;�N�����;%�������#�!�$�����+ƟIkD�2��:_��'��9�S����1*���IrÉ��N)�*R)�y�C�c����c�>ey��L���y"�t7<h���ɶUhY2T��D� ���|#>q����ʆ	]-S�]���J[�<+��i�l�P&�ʓ�\AFG�<Q�y��'��e2�c��}!�R0j��
�s��'z�2Q'
>-Ʋ�Y�/	�piȊ"�'�<�j4���������.��	��$+�S�$Kd�A�D��
ž�p�!�6�y����?2��z�*S(U� AEG=(������O�pRόx�J���q�ΐ3O̅���M�t�$C:"����O� ����6�DP8y<9��ן#�dlzFg�D��d˚#������zT�Z��M�Y��b��ϓ�<9����Ri�ӰM��#1�O|�<)��וhbe[d��0 �8@2�AUQ�<A4����`��(ՕO��٧�K�'5?- �@�-�`1`�`�6]� ���J7D��k���8�`�9P�N�x��!��4D�(�ᬇ�h��(�7+ȪfD�%�C-D���S-�:A%T��$�ƇF랕҇�,D���էE�_�8}��ꐥ;���rD�?D����ۇ69
!k ⍨Č��N?D��y�d(z�y���1"լ��#D���$�h���ۂ�U�BPX�R� D�(���
k.p+�D�n���,>D����+��9�f��j*�%z�#=D� a��v��(�.R<H���6/?D�x�'�Oz:P�3�bQ�DjQ��i D��0pH�`��p�hܿ@�1���#D�Z���0#�+`��U
:���F D�L)�ԸP�" ")Y��
��;D�p��Ŗ,qZѰ�e]7|�ꥱ�a&D��'�1NF���)}���#�'D��F��6��g�ܤj�a�q�*D���HY�Z�H�ѳ/@�F$�ʆ�(D�� �D�'�dٓ�I�3�dUG"O<A��!U�s��"fѠ��`IF"O����+Cx	j�H�M�t�{"O����"-�h
33t�.��D"O�A��*ؗ�*h�ƥ.\�&D�"OB���m�&�(�����2 ���$"O��"#��e���#�.�##�T���"O¤��E�$u���!��EK(��"O�l���njb�Ib�hhA"O��9@���Z˂��w<�4�&"O�	�޲b���Ҵ��ȐmS"O�`Ф��_��$�E��(A"O��:�(^5��YC$ �"�<Acf"O((�5���8�D��`�(�ha��"O��Xb�le�h#�@E7A����"O 8ږBF�~9J���Hu ��T"O-j�@��Y~Ҕ���c^H��"OB�(�JǴP�
D��/�cK.���"O�i�2��""�`؊`�� 
����[5.�Z��G.��A���'=��1`M%)|�u!E�����	�'#�2��`��H�N���^���'t�{Sl8u��	�����'l��-�
�G�N(�����Ci�<�+J�L�4[ө�(z\���n�<�Gi_+F�R�iV*<��N�q�<��"9��-�5mw�Z��m�s�<�p΋u�F�𲂕�]{�L:g��[�<y�D�/^��H1qiV�5��|��Շȓ!(,�y��.�`��C����Hs� ��ȸT	��`0�ՄR"���ȓ5'�`b�-i�* K��؂d�\!�ȓo���s#^2~���eMԿ`����ȓq���S�E�FL�1���88E��M3>
�TK��M�Ǧ7� Նȓ��墵�\�>���.,~V�̆�k,�񠂆 9��RT-s_�ȓ;�x�7n��O�F�ñD���نȓ]�1H��9CaB���ɉn]�t��`8��0���}_�Eۓ&%Y.y�ȓWLT�)ǒ�+�!�׍�R����ȓC���Md�(��u�Q')@r�ȓ3)tP{��ۛvY��Zgc��qG6��ȓo��{�W<c	���DR��9��ywTM@ �D�p,�0�+�#����:Ɩ�!���ͣs��$b�A3
�'��$�A�<@�2�2�j�!���	�'�z��f�J��|����|	�d��']Hp�!��^w^���j�6�&�C�'y��@�*J�?�V�V�O���Q�'4����1�t,ȅ*���Z�'��b2��$<��#�W,l��Z�'�B����9�q�o�*W����'��e�g��"JL��i��B[<�z�'���7D(=S�Hcsg\�-i�j
�'��7 ¡S)�ł���66���'�f�:ɟUq:�"�%I��'V�j&�xdT2�
�o�d���'�&ᘧ�GZ��i;�6q��e8�'�49�PIJ�Ԏ$���X:����'Q8�.ߐjzD�BD�!"Y
$��'�h(�eɋ�do��D�ź���'0diha$U~���c?
te�
�'���Z )*t�Q5���7;�m�
�'MvR�U2O��Y&~10 :�'�T5����3� �H�"��"|r�
$�<i1n]p�"O ��A�^(����1%!8*调�Q�\�Cb�a{��ľY��T�dG�!��qr�,���>Q���m�J6���]�4q�W�Du���X�!�$�i��S���v(�Q;r�E�C�ў��f�{3��Iם)n8����o�:��Ϛ�MK!򄄳+�`7��
��X3`�6p���L�s��=E���1�ް[U�#�(@��)�%u�!��O2�V������rgHQ�_��E�<���'�DirgZA�n����L�2(ܙ����v"j���9?`�܀6A�![i���(C�8C䉭C'��:�E���!���d~�B�I��IQ�#�6���iR�{��C�IU���3:�M��Q~˖C�I	m |�k���hX���Х^krC� -"RhÉ�"U�<���`�E�vC�	�g��-Ѧ�L���)�C���1�B�	�K���(��H"ց��� _C�I��8l��)��6l`�A%d^>�B䉍ꬼX�$Ph��F?�B�	-uI"��C���p�Dph�e��C��
?�9"�jV,^�<$��a�y�tC�ɏPj��/�dKİ��hљ�0C䉭|�.���ʥvb�Jq�� )�C�I:]�ܭ�'"��&*Ra0J/F��C䉥d��:�σ!FȞq�
X��C�	�Z��@A�ȓ-����s��zrB�	9"�F�I��\w�E�E&��{��B䉵Jk�`u���S���r�G�>:��B�I�Q� ���ؓ!�n�!���/S�dB�I�ph�[(��`Bzlzd�!S��C䉺1v�ě2����\Xh���H*�C�	 W�ȑ"c�H'[#N ��T1x�C�{^�0;�C����`#��V�PC�I�Y�uS��%k�����M��C�	�
>`$���Ui��������C�I�hp�@�5M���*�ȗ
RC�C�	�<�bD�BmA!/�bѡ��Fm�C䉱-�~����o�P�c��]�dC�I�_�ɹan�"6����^�pC�I6���i�e��e�
`�f�Q?$� C�jn��b��
0P��P�O*c��B�I��T��)�Pj��Jd)L�l}�B�IBE&�:�MSL�m9҃M��B��y����tn�v�L�ÄFȉ1]�B䉻���$�?7�)@cM�_͚C�Ɂh�
T��e���~ж��%�!�$2� ��*�j�R�ӼN�!�dF�lo�x���Q=fҔm�@9o�!�S?0�2�1�&A�0��mr���|]!�--��D��ʪu-�`{��T�k�!���i�|��6�
��AT�ɖf�!��3��
J ��9�!�D�,/J@�#D�<"��M�0�2��=�2˓b6}F��OB!�F͂��@�I�ՠY�h��0O�U���܊A4僂�I�T�6����ڭ}Oʡ �!��)+�lZ�I3\OL#hO�z�����?=����'d�݃�N��[��p& +R�L�te��:4Cw�0��MpFC]e�<y��$#��Q+@ʘ��u��Y~B���0	Iː�F�1
X��T�9k�N�B�Sc9`T��
A�����kj���ƚc8`గ$� qPdB��� x��-Z�ěxO^�#B�E'F��Ǫ�#wJ���� �O<�����YЈ����D���B �t�آf4�$���X�$-_��Q:�%^��X�����N����@ߤ ]�a�ALKY(��ĐJC&�3Ǫ�t�.�1`d3���Y�@Y�'7,��N\�1�ܕ�d�fW�� 4�Q�? ȣ7�
�{�ċ�ɔ��X1�  <{B!���7�$Zp�]��؍s0,E8�Pj�QX��\�e!�A�`��9������^?-��B�Wo��(0O->�,"D����+�T�&/��C;����@�Z���"NȤl�.)�C� +��џ(}�'ə��ʓ?U�ub�}�N�g*H�Q�ک��I��y"�;wz�����:(lQ���A�~���5��muc!��Y"��W-ߎSf�A�F<�>�hQj��Ӌ#i���P=�|,�?��'}�݂�,�&O��Go�"��F'�,I8�а#jƔ+�(�(�aI�������:�d��$0�f�CG!O��9�ԀB%V�$�!<p~��KL0d"���5�t0�#� M��1�L?�)��ǯT�"�1��U&h8��3�=D��&JC���3�N�9z���G�؍m�~�P􍞽V���ݬ~^�����'���X���	�_���JP�]�V!�m���X.hV��d�4)�z��F���h��~�L�Фk,�z�P!�v��y�g�U�N���2�Ǎ��O2� ��9��nĎM:6xy��Ɇ`(`�SG�{�ƹ�A��)ĎA 1Ƃ�⡪qmƿ$�Ƥ�¹_�p L�*��~2��/w��ms&��\+.��gG*�y�)ܷe�@�%��+yuj���.-r��qKF ̔])(����a�����@E�]��Ȩ"OF����l�)��T�zsM��,I����FKA/L���琖e7�Ӏ"R�'oO�,����-	�l���.�I��C�6a~��BBbU�V:'2��h^�3�𘶫Y*�r�+�A7��=js!̎j�����L�x�'��EpS#'��T�#�S3Y�%i���>	j`\��dӓO|�U2����!D>����N8��2��ǱI6�
R ��j��x���-�p?���0D����y
�(t,B�<I4�@�,�D��'` D�6\�F%�2@��R�y	��O�J�!���2��"Ts���:�'v@0���:��a"��R��AR�'E1? b���-'a��ae͞���i�?M�r5�6�Z=�~��K�{>@��0/	#�Ƹa�"X.�p?�k�-����S�Z���ӎ��wqc�a� *G,���3?�f ( G�gD�b�	7��	�B�F-0�f.�>y#�X�-��yQ��2C�}�&��5�Ub��}�d�2�_3.��Y�$D�%G�J�Q��'�0-8�(v.<`�֧e��e�'�$�a�7hxиal�'�<5���8d��7i�'T\M��HD3C޴�R��ˤ0dD���	�WZ`�DƬ>���\��X11b"nܰ�u�K%��-� +�'P-�F��]�@&?%�V�'��	t�!kG�+ ��ڣ�j�,��y邷d�>TD����s� \�NֱKv��+Dk�NP�~�n	�4矸@����41O("?�V�A:�꽪1&�� ޸zC� i����|r-�b�w��0�ц�Кi�m;� 6=�:��'�_�P-���K*�B�	0Or�$yg��
&1I��O��Tg�r��xC�I�"4�! ѰLw�)����O�ljv�`�ڬ��f��*�7츁IA&A����W�b:��xt�ޠ/��K��~�:�\GV�˓x�xD��Oα��	��2�\�ԌO� ¬\B��$��dY8�� �=�M��2��1^�. ��ǆ1f��k	�"��õl�Xyjs�1,OZI��#S<\;G+�UF�D	'�T&N0<�'�H1��?�2V�֨��x�Rn�+H�t4!���#�X"����t�Sh<1�(A�52DY�*c\�b��)c�xa�#S��՝!dh�"���69P�S��=�֏�x���
V[�&���\�L�C[�<J�I�6b�X�{r.���^ �f1D�p8Ҁ[4ZU�����"�la���.��|����Bx� L�тA:bD��j�U!��Ժy��e�uG�7����%��?6V!�$ҠO��d��B�i|�)yԇ� 8!�DJ+qX�)�2�īv�������!��,�^@�5�N
h� �Rw!�<KJ�}�F [J� n�;�!�������U�&Q:DM�"�!���Ϫ�ZG_�aelP�^!�Ԛ'�t�xwl- 9B *C!�ą)v�8d�L;g-f��!��9H(#� &z���p�!���(p`}��aI4����J.{�!�ըvX��p�}6p��q!��H��U��A�J��Ð�3T!򄊎*��-�&�Z�$�C�·b!�d�Y���� ���A�0�3����!�D�\��y���I���6�\�!�� ���V�L�1ɧ�LfgH���"O���6 C��
Ь��Z���"O�|)V刾-b��dI�)3J��"O��4%N�]��e��>8���+f"O,P��CM&h��0C�ʅ/ �����"O�	C���T�ʈrV�ݪBU�i��"O�Yu��q.�49c��<���cp"O��Y��"YI��҆)༴��"O$���f��BDE�{C��Z!"O��Q0-����&P�E 2�"O>Ș&��B#��+`� ����"O<[ *ѽh;�$�u��=8yz�A"O�Ԩ��dj��nƹz�T�e"O�@P�g�	�� 3��[/����"O
�)�6K�rM��*
�Dt#�"Oԙ	��C�	P�XZ�hA�W�$���"OΕ��,Q����á�D�F�ƅ,$!�$L-�ܩ��Y�_7�Ѱ��M�JT!�
�CH�e/�+��cQ�;<V!��Qz���"^�Q��cժ�FE!��:Pظ���'ȶ��]h���k!�6w/l��$�}�NP	�k�#U^!��O
��`�Ƒq����l��|C!�1cH~��K���0���̄�M!��5s��0��[*��q���0Z+!�dӖ\��}�.�0j��X�a		�C!�1��s��=���̛D�5��+�vD��播/�ȉ�6A�Z�b	�ȓ$�X�b���&�q Iܴ�D��`*�����6s�����Z*8��ȓ[z�Qp�-^Tݑ��6�x9��9�T{�aY.=��-� A�3In-�ȓB�u���٪o6�Iqh��XAh�ȓu�bpB��K�c����R�ݳ�^�ȓ^�a#ũnz@j�`ܖ}�|��[�@Ds���4	�jM�#��wXV���f[�8����|El�;3��O��P�ȓ+����D	=?�)��o����|�-3��
4�gb�.0���ȓ(5��@s*Ū7Ju;q]^e����	�8�Q�B�p�Dx��᛿f�d0�ȓ6�`PG�	W�����Q�B��RH4�0���Ue�(�8~�T�ȓv0�@��c�\%����ݾ:���ȓGDPKO 9��1�O�x���U.��_�Є#��Zֶf��B"O([E�7!�=���
V��(q"O� S�IJ�*gv������3O�U��"O��r�䉼%+5閈��$��'"O�lHG"=I��U��$| IC"O&�{nA*|�,�*s�^�S_R��&"O���sI^2}�\Ԣ�Ȭt58p�4"O>�S�F׻
�iA�Γ9��!�"O��Z���).Z���-ޞB�8aV"OA�$�Y�6đf�VҼM"O�<p���:;�*�ǥS[΂)J"O���g��w}H�f.�����"O�<kF
k@�d�jB�z����2"O�ԫ���gO�48�/�
�f@*�"OL}��e΢N�!�7G2g��4�d"O�"��Hi���s��)C��H3"O�Ęr$͓/�U�6O��#�T��"O" ���b������
 �t�$"O|I�`�)wF�5k�mLM!"O� �=qG
��'Xl���$��<"�-S"OdȈ ���!T�����y/��("OX�{��D:&a)$+�0��J�"O�|�ׇQ�X���K�.Y���"O���Š�'|��x!
� j�x5"O����o��"��Ks��06�!�1;2��¢�FÆ�{�ʘ!�JAv��@@Lu��D��@�5l!��i��@��b���6�I!�G�!�$�%�xq�2l5��ݷ	�R�<�e�F���"T�
1��D�KJ�<�A�FzT$( �!L_�(0��@�<YP�h���!��q�H@:�n��<��� V���A�%�S:6�BgJn�<Y$��|h�`M��V�J�)Io�<Ag�к<����/�H]
va|�<��b��R�=x�ҌPl�J�z�<y�"�{�L��Ed�o �b4�{�<�Rl�7���B�ҊVDDx��B�v�<�B.=�>��foA<
� y�CH�<ab�zI�A!�� ��=�WJ�<�r'N�jO����m7w�2�j�IA�<i�`��a_>4��7&����Â~�<Q�,��1E��di��)�.1�#�W�<a� ��+�H�%j��|�^�@�N�<���|o,V�	�F�|�%��I�<�իT� \�HȈc�����D�<)Î �y��3lD�T墩�-TE�<A��E	tzi���Ti��G�QC�<��m�v�7G>w�VH+f�g�<�L�7cGN���Ѹ{gD�`"�]�<�!傼Y�5c���/��X��P�<���ØB���R�ȸ:�h� n^I�<a�Z�6�
�"dΞ3��!d��x�<16G�D("���bז8��5��M�<�MA��(<#bE4RPY�	�H�<��"QG���@���(n��Gj�G�<�3sz)�teV�8?n4�t���<IGC'z��E��l�*,�f��%�@�<`��4:�����!;��u�g�P�<�s�����O΁�q�O�< ���-�hY eDI���+�GF�<	F�Q�~�jBr�ك��N�<�2��&ojv��SD� nēW�O�<�� G��|�R�A$$���XD�<9�V3v\�+��� -DU�#&�Y�<�%L�9X��	���1t~
�b6��W�<��.$���RdKƲg�F���șu�<��/8 (��B[L����c��s�<�өY�CB5*��
�-*�h�n�<�@˅�5i�@��� ]�6���,m�<!�	J�f��У� ��}�c�d�<9Q�њ3��8R�X7��[C��c�<�5��n��li�Ηi��9*�f�Y�<��@�"��͙���'�4�'/�N�<��c��
P�����9Z��U�BȃI�<!�G	�&���ؽ��Q!��n�<A�/E8;Ǹ�Q	>z|�e�G�i�<�A�!.X�Y��B�T4�a��^�<yFG�ДtP'�Ȕv�J��OCc�<i�,t��DR��T�r���Mc�<ٴ�O[
��)���dˆf�<iA_���L�w+�em�q�$��<�ծ�0} &ތ~��dqA��`�<� R�10O�0(6�����* ���Y�"O�y�
�!t���Q����c�H��g"On�vn�fV�����!x�Q�"OR�ҧ�7h�0�!�КGT���"O��I�BTZ1ȢΊ�Z��]�"O��R��P�x��XW�r���9�"O �@�Ƣ&]�����ys�=�F"O� �P%؆N�<�cL@{mȩ�"O$���$ō����.�����"O$��s��@��Y���H���x�"O6T2T#�87�)���&(ϸY5"O�!Sp�� !+�8��AŜ_��U"O�-b��֋4S���Y�́�S"O
���[(n^� ��h(0c"O�xԪ�3�jD�D�@��m*"O�i(0nY�[`���I��z7|-K"ODԙ�d�-���[�Ȕ�@/�1S"OX�i����)O4i��"O��VIS,d���S�J�|A�)�"O�t��cĂ �Ĝ@ѩ�� Y&�"O:<8t"�:T���D�R�0�ݣ�"Oz�@�+\oB�CS�Z�o;l�h�"O�p�&��1c�\��t(�@)%[�"O(���A�D�����+K��	�"O�!@���%8��X֥L���	F"O�$e�����6�<䑳"O���Wl�&�ha�a&ěZi:��q"Oj�ˁB  ��T�7�\ i�V�2�"O�(R���>n���زE�=�x��"O����cF�����U�X5WH�"O�5(0��5Q1��03��Y��A��"O��*q(ӥ>� [W+K�^۰"O`�X�9E�&��N���p"O�1@c�'y8#��ǄE6�X�6>O�u2�'!�Ot��v�Pi�}ѧ�H�F�	��'�2�#�3����x �#�޸u���b"�-�!򄁾��%�`cE��ы�'�Y�qO�Q��E�[�#r�7\2\���՛���DMi�<)e�M�Y��Q�]
:�VFHW-ĸ�e�|b��N���S�l��k@&xKb'%�;p�!�$V�#�<�j�K� b�X��Ge�5�b5�)�+C�z��I��Qh�k��%�xMy3���"����([X�P�2��>����0~��͠��\3'-��� l�<��]� >���-���ɏkܓu�T�T�T�ȟ�x��M��A�b�S=];��Z"O�}��(p��G��|����R)*u�&�����<!W�'0'��r/ӽ.�I���`�<i� ����|�&i�:m� ��%P�p ��N�j�a}b�_?&Ŕ����O(w�d�8�P4Ű=�R���')��]�`�v��jX��{�'�pISelR�p\*�P�F-n�r\��䗎I��,X<mWZ���N��X@a�FY�<Av�.sE� ꃁ��{�di)5E}�<�3�RR]�9a�\b?Y��b�<�@U x�X��M`�F�i#
Vz�<�p���"�%�" ,X����r�<!RI�"����*��+S.Wm�<	��d�P=��)B�s���#���n�<ye!�4�8Q���<��ɪ�|�<f�}�0��L����%�x�<�u��0�c(
)D��x2!��]�<�a ',`��R�)k6��qS�GU�<y��M�QK
��e+H�1�ȁcM�^�<���ۛQ	Ј�o1%1B�A�l�X�<� d�K@"؉;*�%@��Z#`�t�#�"Ot���%Ti��-Ȃ�)J�#�"Ot���M0Ȣ!�l�-vqBS"O(�x%�8
b@�Z�)����"O���q��~��Ac��3;?��kf"O�%#���f�z���J�2Px��"O���v��w"N���	�M
�[5"Oj`S2��,N�S��T jt�V"O�,+��+(f���M�5v||��"O<���(D�Pp������"XI�"O�4��A4
q<��$�~jP�4"O<��`�'4���q�b�2y�|�s�"ObT@�]�hr�l���֦eq�a��"O�T)��_$0�\��*�jl�t��"Oq��l��?��!�*�kXp��W"O��:���9���)6't͐�"O�xpS���@C@hwՃR"Od��gI/mTԂS�ԾO�\��"O`hLƛN���瀜�1�ȅ��"OX��2��7��!���j�)��"O�E��ɕ ;�pcL�00�U"O��qgV�z���� 6e^4�"O����V�H
\�XD�ĩ*W@���"O��ۓ��m&MC�Q(7����"O��h�	��d(�C+�?p T�e"OtHz���o�x� @���"�S"O��Ж�;8�E� {4���E^j�R����7w�4ʷ�'��&���Al�@��šk���	ߓ��'L�PA"L	z7 ؀���62���*O�=E���'BJj�dk��@{��S��,�?)����MK��3�3	#��*G ��N�=1	ç��xr��y�8P����IW\!�?9$�i�Yy�@A)"��	���V<0�rKЍH�I�6OH�I�bL>E�Dc��!B@@�D�=G�&H ��+��$ʈ&�Q��Dx�Ǌ�q;ZY`��-Y^��7�U�?���[pT#�I�"Uйz���F�h�=�	ç'Xs��މ'�~����=h[���?����~�CLE�>�\��lH�~��C��|���=YV*<v�����M0PK��	�7e���kW(���RB��@����O`xܟ �	�SƖ�۔�G
\&�����[�txF~��I�hz ��ŉ[�2qY&�«a�d�=�	ç(�paC��9���)b�{���?i���~�e�pcP�Ŀ&��ݻ�D����O0mZ�b�!s���ޠ\��i+O��="��I�X�c���C������(Vb«���<�}��'�x]8F[$M/&��w��#Q��*��,ғga��ޘ*t tv�֤j�Ĩ�m.��'tў�ON]�$G�6_F�cf�]+�Z�(L>i�����n�萔�щ��lQv*���	f��(��pB�CS\itQ��k��M���:��';!��Q�X�O�1��M�D;b�(�2�����,c=r���4#���
�d������IG��@q��)�!�D¯{�X��pnT%UI �U%�-�!�d	��c׉0S5�E
$E��Q!�DG"z�4�B�H1(��֤R�y�!�DT+�hx'�	 w Q�w��!�$�RzIEjֿMA���՝�!� (ָ���DH u1���ƍ	X!��M�}]"�('B�3���	<K!�d��4B*���h̠	ʌ�pd2IC!��#{p��F�J 6](�A�ۛ4�!�=fT����6�,��$m�c�!�D�2%�����L-r��a�v�<!��׉R��5�@NɃ�����L}�!�� �9���lN`͑�h��\��P�"Oz�Y�DxYP����:���xF"Oh�k��ӈ-�� f'��z ��"O�e:��D�#QƱ� 4����""OX���77���qf��D�!�R"O��X"���8P�%KJ2|m>�d"OB�Bgg�f��;4�"Jj�+�"O��	�ʫe
����I�i`��AU"OtI��ԅ/7~PȄ��uO��SQ"O��S�
(�ݐ�a��W�VԱ�"O�	���,{� �y`g�~.<��"O ��tϚj�p9EH4d�#r"O�Իd�ΗR���ҀI-/�\�S"O�IJ�'ǌ5x����ʺ$�5B�"OveHC+
4���ǚf  ���"O(C0`:�2ʓM��:&��"O���s�� E�!�uM� >p�a"O�ic��@���#���\n��3"O�}����-c=���0���CFN��"O�<�᝻��L�G�Y�%��c�"Oj|� �U������^�a��	�"OL�CQ�!R�{���ԁ����S2Ep��պ� I��	�<\��}�ȓ�(q��#�*ؼI[ ���p*(U��z� 3o�3K]�HSê�*6����GK�#b�2#pdEOڦ)�����l`�Дo�܈9Aũ�
~b 	�ȓh�j��0i*�P2bZw�R��_�F賃�N�^܄����9Np̄ȓ1�T�'o<C{�����:����ȓ _:��A*�Wȅ06*��jyZ���8��i��O5��Y�E��bp��ȓ^��� �FYEL�̟�SZ�ȓ��8JՋ|��7�]1f��}��b[��ې�_�>���4M;X\���m���0�Q<!$|�87K��^l�ȓK'� De@��@U��;3�r4�ȓ#�>U�n�>s|�i��6N���r,�h�0?XF,�r��2.����+�Z�6���k�J�'!T$�ȓZ��2��^L�S�����tu���޸R�f);H��ц�`��ȓ7
|,R� ��0e`����іF��D��;5�Ӧ�Å,N���4 E�`�фȓ EX{E�;T+�xwN͙c�h�ȓ`�F�%�d���p4x�ȓS~�@ �Ǫ3�^����}Y,���F��e!Ӭ��7�E�!!���dp��[<������l��bW'}|�Մ�	 в"�֥Ř�B����xu�d��t���r�� \5TewÒ4I��\�ȓn��(Q�ӎBI��
�d�E���uF.e�Q�ىR\r�
e띃S�D���:2˴���CL�<^�:��� "�!(��ԻJ��0�e!�"�ง� 0R�m�"_�Dp�X!��9��h�k��t2�	��cW�g�T��ȓ7s�qY�+�B@�[� ,M>���/Ә@���T�|���F�q�Ն�R�� � *\p�9��
#u� ��ȓ5#0��hE�O��Z%�W�rz܌�ȓ/I� �c��4�^�kui��Gۂ��u�,X��&R��,ǒ͆�F�\[T-V�'C���Ĝ�4�<��S�?  @ڔ�ab � mނN����"O@,��hJ!E��Iq��+b4�` Q"O��sE��/�J='*��"O�<2v�ߕ�j���#.I� �"O:LA���c$�x�t�FM��D"O�	ԥ��*��05^�H�����*O�E�P#�6W���G���y-�� �'��p��K&v�\�Ԭ�
w��8�'�l0�q�	=O ��f'Ț[ӆ��
�'���z��H�qǌ�(��P�
�'m�\�AE�)pq���0.�q
�'��}{�熽BS$sv���^&�I	�'���C�ٹ�I���$s��	�'c6`�'/�}l�9�/�'>E��	�'(� ���-]ӈ ���J�7fa��'��ݡA�Ds��x*��2��i8�' D�kүfy��Rj�?	$�	�'��2B*#��%a3
�)i\�"
�'���#%лv�P�J���k�'�U�ҩ
x\^1��jYhd^�h�'�!�v꘽F^tU� /b��9)�'�Z���+d����ea�Y����'�eR�ŋ&(���t�YY��
�'V���D�p\KS�W!M �pR�'��ȧB�.���*`�Ҿ=~�`�'7j ��E�ng\Q��B�2���	�'���&M�JsJ}��D5U�@!��'���w�}%��c냫P���p�'۶q�
�i��젦F��WȈ�[�'����"ީ8�u��+�6(��'=а+���J��;��(�B�P�',�uJԉA+*�FPKf��LƼ��'�`(�ul�)c6t�v��7Ӻ���'�� ����DB��R�2l�l��'��j�Gܢh(����K�|p�-9�'~ ���A�>>��\rRE�x[T���'�V0�d��H[3�M(1`��'Ҁ=�rF8@�00�E��HԜ��'u�M���<w��R�k�6i�*0��'��F��	S�����aϟb�����'$��v"�
C
�Hku�ɭJ�E��'$V=٣ ��Y_Ld��R;.�\��'u �s1���<��x)�5�(��'Și��g�
(� �я@����
�'��e4�IR�k�J	�8�Q
�'ޗ�sm�dP"g��0�x6�M�<��@�j&�R��S/�飔��mX���Oz�#���8�J'� ^���ؤ"O0�{ժ��H�ltI#��7�1�"O���oݰMl Q�I�(!"OLi�֭�.��` �	�Ĵz�"Op0P�&�1��A�O�Z�E�2"OI���S�a�6=b76�=
Q"On:d�K'0a0'@"9�P��e"Of5Ku�AL���cŃz�Ԭ��"O �ˠ�'2�
��sB�$v uKR"O����nYKt���`�]KZ���"O��B!ͻ?�y�0 �]N&l"�"O�A��h�<�f@��$v��s"O��*v'7�XhaX")���b"O$ ��Mͥ#vF�aZ�$Q�"OF]��F&cd����لy촐��"O�ur�FlG�i���e��["O�h��C�Ȇ2�<��0`�"O� x�+����Q��-J�f���"O�M!��� ���K�!7����"O�L$c��+T�ѢE�c),��"Oȼ�v'ǒOR�&��lz�p""O�QG��>X���fWL\1(2"O�t�� E���#h��C;��s�"O��r�Ħ|!�`"��	�u+&9!�"O�23f�:�Q2Q�ɉj��W"O�e�ӄ�-8�Ѣ#ߊl	l�!"O*�B����'1������;*����"O��� ɑ1cv(�Q��d�:�
G"O�hy&� �Y��	eC�6z��[g"OdȀ�K�)I�dtKc��;m��90P"OD���f� &�R@9�o]1�X�E"OH�@��_&!����Ê3�H��"O�<"q��F����vd�ջ�"O�*�喴qϴ`�FN�sĬ��p"O���C�,x�q�M�c����"Ol��t��\� y�tI�<�p|�B"O����C�4�����˃�f߼L8�"O��s�[}��R3%B;��!�"OXm��ń�0�Q*��,/!��p"O��Q ŵ)�h��`�Z?Pb���"O�X�e�Ǯ��}"g�S':�詉�"O.�A��G�J�*DA��:�2%"O&�umͣ#<1q������"O(���aG):W�X�+�5�"�0"O���@"]QB��f
ë�l@a"O�񉰌�-&��Hҿ[�p�  "O����L:>qV�s�`D�B'f�P�"O��pӆD,l"��	�Mw�mY�"O�]�v(��]�&e���V;�H�U"O4!a�ɝ=��%:E�	�K��x�R"O��c��v6��j�N�:;�@A�"O���]�Z��D�w-޹+~����"O����׺��4��B94d �6"ON4P#�q�XUY��2�$4�p"Od���M$xz(�2B�.fr��"O�9���xX\�����&I�pa"OL��w#W�H�t�5ɘ&t-�Დ"O�p�'Lص�ll9��4����"OL�@E��@�T���+�ftz$[""O�P�+=n�j����[�|0�"Oz�u��G9�82�U;μ�"�"OΘ��I_!>����m�!b���"O��) �k�p�p�-зw�3F"O�U�e�5\�l�䬏1C�Ba��"O�Q��EY��� M�l��ٹ�"O�U˂,C:�(�F�0$w�Ea"OB �K֖`�N�&'ɉY�83"O�i3P�A<(E�e��_�
b2�c�"O�%˧�N'	"h(t�S(~6�Ej�"O�4�0A�z}�0{ �D-4H�3"O �'	�jh܀���(n?���"O(<��@ m�X�X`��)g/>�(V"O0(�W���\7�Q#䑒5�P���"O4�	�   ��     }  �    �'  �1  o8  �>  E  EK  �Q  �W  ^  Kd  �j  �p  w  W}  ��  ۉ  �  `�  ��  ��  X�  ��  ��  ��  �  S�  ��  ��  L�  ��  ��  2�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6�F{��'O��V���&�;�+0:��x	�'%��"J�[�]�R�K2r��"
�'Oe#W烹�R}aC��z��
�'��;��7�������L	�'�:<*b&K"4����M����9	�'نx!c̓>�D �,ݻ2zX�R�'��@ �F�9<�m�7I�"+�a�'ր����>��Y�
�%&���'��0��3L�r5��M/� HJ�'U����J08fx����I$p:<����O*b�X�S�!��G ��s��PDd�o,TC�IlߢE���5Tvf�����}�LC�&�L[f�R%'�Y+$�@�	�2C�I*zX�ic���%|���g��d�ʓS�v�<!����
/����县)�B�ٲ�ITl!�d	�N�(4$Q?a*FL{��[6M1O ���_�V�� ���C�!ږ͒?!�ͭ~��M ��<
ݪ��5lN�!�D[�$��BAĚ�0e6���Z�q�џpG��ч	�fh�ǈ2���
-�y"�M�s*ZT[�IU�sԢ[��D��Φ�?�g�Nj�yc�Q�����QÏ/u>����-?BM�X�A�!Y0I¸��u�Δ�䓘0>�D/��>� ��E�=N�U�G��t�<��( F�qb�5 *,:�� q�<�B鐨>spU�Ў�i������Bi�<� �k�CՀH�)�.u�r�#u"Ox��^ƴ��񊓚mHX0�"O~�0��)[���#��0 ���"O��i&i	?f��t#��"9^����D3LOf}�լq��CC@��Bo��"O>8��%°�t�)u��]j��Ҷ"O�8BR��#`�(��lN�1�l�å"O.�ґ逜!�I��B̦H�Q�3"O����Ƀ]6`����5e6��?O��'iў��X��Q�W8|x��(%� {"O\|⥭�9DT���\$�8�"O%��iy�1�-�� ��S���I�����C0�!B8t���ӎ�MR!�$��Q4m26(߯�V�� �K	LP�{��	�Pt�!�"���>��a��I�A1!�G%R��p�Х$�l,z�M:W"��G{ʟ ��R:*P��x�I�	p�n�#'�'��I�YDT �刚:E7�(ڵ	�fB����kk*tH&�F=	�F-[���-�t��p�\8��,�f�t!�kY-a�"D�ȓ@�}���T3O���i�4Rs�G{B�NF�I�_�5���n&N�)�g�5^B�ɋZ{�uí��N�T��Ԙ��C�I�r�l@�C�:}���cCC�G�"C�I�
d0�a��	E&����rK�B�	�E�̍)�L6g�FqY��Sns�B�IM�.��TN�x3a��}�B䉇_^`p�1ֻq���p�E�#a^�B�I�q����l�jhr���_ �@C�	�D["����L�#Ǆըl��듎?!�)��),�� �KO:dQ��*�h��H�BC��_��t�ī�P,����
�{�8c�����'j�Tisn]1�	�gƼrh,��>��|���i6EQČ��3���ɗ꓋W�ā�'��Q U�0,��4��90,[ۓ��',Z���.H����$��70Ѽ��'l�4�e+]"
"���"$�&	��'
(p�ϋ�R��#��l�R`*�'6 �3�$�S�pB�B^4f���X�'֩·�+g����7�Y�Y��\�')�)҃f�=��Q{7��)UЮ���'�H��d�z\�#�#vth��'�b�Cq�ѷ)���í@>� ��'�����G�?|�H5���<�P�@�'�h�e�Ò%��ȫ�B���e�V"OL�Z��̆:���#�
IT6�"Oʜ�K��Z&�
&�R�Fd��"Ov=��۾7f�ECF��w�(r"O����CI7C���ɲsA�r"O8(f��4���0V�|4�p"O����'JD�Z��ڍV�q"O�QWL�ZX�C��W<7�j��"O4� R�[?d�t�+��> �2���"O6����8kx���n�F�6E0e"O�|#�N�0�n9�D�I�.�
�"O�$Xs㊑qԈ����1�N��"O�t����Un�va��/v��K�"Obm�5C���� ��V�z_��p"OD)�b��8��"fM=|N�r"O&�0����kj��Eʢd99 �"O�-�s
�{@v5c�/2��pG"O��G��5�v1��l
�o�I�"OJ���"�*Ǭ*(zĩ&"O&�Sԉ��S,��X���]ؕ"O� 8��GN:30(�m��x9�"OƉ[u��	X,�T�K�(	w80�"O���3+������[5dr4l��"On�hG�M0�j�2Ȋ�)%"O([�ׯI,Ќ"qG�0� �"O޼z�Ì)�D�D��4�"!C�"O* xt
L�w*P����"9��q�"O`�����.�v���Jh�� �"O��3��B�?}���vYHL	 "OH���1���['�O�e�e"O��;�(�����bHA�:u��"O^��2��w�P�jQS�[�(y�s"O�e�f��W"���A�=�ɱ�"O^�:���{MVTb*
0�H�2"O<��͇�x�p�jtnN7'42�"OJ0�b<=P����c�2N�D��E"O��(���!jf�J�C�)B�0�W"O S'�/��q��S�L�L �"O�Pq@I�7%��p
��T�B9҄"O�)�� E�b�d�`V�(3��4��"OH<�Ѯ����ՍB�h����"O�� �] I_�)8�FH�;���C�"O�YX&�#8kV �d��)�Q�"O�	�'C�E,��(��=#��W"O,�8��`�Ѻ�h�:)I�"O"��!��U������&��M��"O� 2S�ݸA����&�&����"Ob`ժ@5Jw�P�R��W�^��	�''�ѓvG�#U���&�79�<B	�'H�a�M��!�rȑ 9���C�'�����<�6ۢ��4aC��'^9!� OH9x�*ԅB
e��'�HH��Ƙ;`)s�h��fbr0��'ml��E��s�j���� R�ha��'�Z!� &�-$S�q� �4KX^l��'e��Z�nP^ZtX�F�@� �'�6�P'�3U���X���5�,�@	�'�V��3f�@r�vN�
z.�|Q�'r�y8t�I;,'�ă >�x��'Q��J�,�
N�m�E�@�e@PI�'he��	Ż ℉�8���'��i�d��f����$��!8�'dB�(_�odU�� �S��' �k`��(blY
�a�Qt���'(=����s<:4��㞣�PI�'��U���6Ĭ���ڑ ��
�'�F�`A��>�ɺ�Σ58�c
�'�d����2FX�4�c���'� dr�'5���蕨6R@(�V��/j�ޕk�'`}avO�8S}6x�e�R*v����
�'�2a"���0���6a�t�.�
�'�Mk�M� s�*�֠He�B`+	�'��s	M�k",�ŭL	5ܼ�	�'��Kw`�3A�S$nP�$�,��	�'������_����c@
Fk�H1
�'Q�P���[��,�A]�KH�B�'W��Qm�Z�@C[�|hh
�')P��^Rt��c�M
�(���G�<�1
ׂW�(A���
!v��(�G�Gg�< m��IPi�Q$�q�Jl���a�<���U7"��e�f��-Gm��+�LS�<��A�P���3��W \�峕�w�<��6������q��9�P��|�<y'/3��ui2�Z47�<��R�`�<� 6�SK_��%�6��v���"OZ��9g[�01f��E��%��"O��g���8xmiU͘�t�6"O���ld�R�K]�J���"ON+�z~D�P� �s�u�'���'�r�'_2�'X��'Y2�'��aꀋ�8	�9�cK��Ox����'��'�R�'���'#b�'L��'��Ժ���(����c�klTxJ��'���'���'���'���'uB�'�ڍ:$�;&����w��Uq���'-R�'�B�'���'��'{�w#�� �*��/���"V!RW�P�4�'�2�'�"�'4B�'�B�']��'߈���h �D�̑�vg؇hQ�����'�R�'lB�']b�'��'[�'��=PA��(��^�o������'*��'S��'{��'"��'�b�'$L�
"EB�~�����+;��E��'MR�'D��'g��'���'���'Cv�AAG�'�j(�4���f-�dc��'���'���'���'CR�''"�'�ʌ�t��Zy�+G�l(sA�'�B�'���'���'o��'��'���5$�%T��(���+sA
�B��'|��'�B�'K��'���'Kb�'r�|����
h��EË�;ud�X�V�'���'��'�r�'���'n��'�r��WM�?O)�I���	QN�Y��'�B�'���'���'�r&gӐ���O�ܑ�
���q
�%��8ty[W
�]y��'c�)�3?�"�ib�#tƗgV�� ԣ=O�!%�����9�?�g?A�4iN���ʢA�Nr�!W?S��c��iH�ć�k�:���O�;����T`PL?�3A :�^��oA�B�=
v�-�	؟8�'��>�V`=b����8Kԁ�Ԡ̈�M#F�FQ̓��O�j7=�R,��jP'l"��c�
.Q?�M� %�pnZ�<�-O�O�нa�D��yr�R��PAcD�([��Af^�yb�7��`�aў���L���ؾ7$.���X�h2L���x��'0�'ٞ6-�S�1O�I�!�V\�J ��x���Af=�	����OB7Ms�,�'����LN�5�*l�4逝i��O�UX�ɚ2k��<���i3h��,)���O� j��ۏL���0�®N�ʔp�<*O���s��4c��"���c�j�LA�!{E`d��*۴c,Ld�'�~7�5�i>UBCˋ� �)�ƍ=�̋ҋ�� ��Ϧ���<`1��HC+;?ɱ�SUv����1Pb��&�ȺM�B� �s=�=�`�X$R�nl��:Hq:b�6�3��܋:��a)I�Q!N0 '*�;�!��(�@4�R��$�2gJ_\��X����F�ݱ���,y��U!�M��',��
uh��t=r�HZH���$.<�s�č�X	 �J"*�h��d&M&��ցЯ.�z��p�>d�Ѳ%���t!p
�(�]� �|�4
�"V�&@@"T�A5������W=lS����#�z��YoZ��������������Hv 0jD��*�De�5�رp�	��Y%Mm��&��p�D�eyH��&��&�� � �k���@L�ɦ}������	�?	!I<ͧ @�zR�H�]u��0F(7e0Dt`A�iW�躥���1O���M	dڐ1���0�x��Wk;��lZҟ��	���w�F����|���?AژJ2��ˆ�$T��<�7-�Oh���O��ra�{���'���'�$�G|����	H�"@{��Ȗ|�7-�O��2��D�Iߟ���O�i�CCß#8Y���'�ߖx����'�l,��'���'a2�'���������n���[�!§,i8 Dޱt����N<���?a�����?qv@"Oєuh� W�#�����	�=�2��<Q���?����V��$ϧhE����8 eX�Z��ɓ+X�%���I[�	ß���>:Z�J'Z<i%��׎��g�;3����'uB�'��^��3f���'OF��F��  �-��DB&#��u�b�i�B�'��'��B���M;��̥
	���S���Ȑ�-���ؔ'�Zt��2���O����%}7��f'N����0э�-��E%�P�IݟT2��ݟ��	������j�/N�D	I��x��A�i���' p���mo�,P�O���O!��$��1�ƫl�����i��K����'6҉ʬ|��O���x�Җ���d�]������M�C��6z����',"�'��3�4��t�"!�]�y��E�?m�jI�U�K����e#�<�	�x���?��O��ӕ-�&�b�'�
A� 9�O|@�x޴�?Q��?!R�F>��?�OȂ+F�����Au1z7�x��'g`�{��d�O��	�6~�A�G��\��82�dT��ߴ�?Y�G�-��D�s�����'�th	�CǼ2�V��T�T�%�d�n�ϟ����j�Iϟ���័�'�q3A������-��m��n��7��O����O��D�<9��?�c��78��$J���oK�Tia펹O��������O�D�O�� o0���=��,2��
f\=�Ձ��64����]���������fyR�'�2[@����t��q'ӂ8�&�A�gRE����?���?!,O�� �D�S0|��Jԋ�/���ˠ�Щ3V|��4�?�����d�O���F&0>��D�|
�HRzX��z4X{T ���7x
��'�r_�x�����ħ�?����4*F6o+�}��Oɿ,�X���G���'K��'��u���'��O<�\� x�X����>��whS(H+"%�Ӝx���9n漤���6Ot���BB�!���F�O	gd6L��"O+I�<e^(���֗]U�@	1�C">��S���D-y���gt!a[�-A����ӝI}��I��D,��#
W2M��e���aϲ �6�б֘�r��T�V���6��g�"M�\$a� ���u��ط�׿�u1ς.B̅R�F�IRH���#Lo��I���Km���f"ӥ$^��O����OjL���?i��E���GL,�	J�؉.����pM�J��tA��+OQ��/��CR9Xuk��s|��'��=X בK��8)r��S��)��1�\���y���w����2Y��Q�ء�~�����?)#�i�O@��ORʓ�Ɨ�y� }�b�9{����".D� 2�D��/G���,Y2q�Xx`��ȟ�HOd˧���ٻ48m�2O��0ʧ)ĉbH���@ɖ&���`������#���	�|�!���rص�F�x��Ʉ���
��`*�LC2r_Pm�c��z�E۞a�MB5�2^�B�&�.u��ڄ�?��=I���͟P��? �ڽ���"lL���̅Ao�\'�\�	ǟ�?�O�t�gď�C����J�)[��P�'\lT�&���B)�D������h�'=����d�=f�F�o����`����s�H�kt^�y+N� ��87��R��'���'�1��E�7e��Bg��>i/��Q�K��ih^h��(X��0J�ɷ`� 8p���y�����бj�Ұ�L�|��LSeeEn�mi�+B�a�-2T�"B����ǦizI|:��urd�Y#dɉoQ�}��+ 8n�����������D�jR6�S�@	-P��ɑP핚S6���OP�m��MK��EO�[Ԫ��)�l���&_0pɘ8�f�Z� [�d��n����4r��'�脣0���`5��CT<�9T�� �贛0��F���-o�:�+��qB��x��ߥ��#�4��0G���@C�^�bI$�PqK�;S�1��n��i����wQ|�1
��6~\)��L�t�5�E��b�g�|����'�z(O�����πUg^`f͊L����v"O��ua���x��Ӌ��^�$��P�I;�HO$�'�&�8��_"A���Y�"�d2H\���'��P���"��'���'`"p���	�PXAˎ�`0搇@��|� ��M��㘷an b�	t\��+���1p�<�ɚy�*�q/�W�ȑ�gI{�P��4i�=)g� v�pcOSpb��ɢG�h �K<��-X]�V=s!g
h��4�����?��Jճ�?@�ig,6ݟ��Ɵl�'^BS��A!O�����|�4�:	�'߈��q*!�]� ��!n��y� b7�yD��0���Ӽ$���&~8([��^FB�r�@�<��)����)2�@�0�ҡ��w�<�p�Ո<B�t�2��>mq�R���^�<a�9,��C��޻{!���Ŋ	Z�<� ��li�}�v�K�T�ENNS�<���ǌGQDa#v��-w�P˅��c�<��9�*�����&.���jf"�V�<i`��!� �fǙ\���c/�h�<ir#\b�b��j�D߶�ꠍ`�<ѥ�ϑ �#��uJth&�p�<AQ�_9�T�ʕ�-#Q�b�b�o�<!��ڕ"x��ߩ
�<���j�<�����uޒ0���#}xLW'k�<A�E�-�`!�@�x��5�g�<q2�_?y�`�y�W�2P0ÊT{�<q�-S5v�*p!��C�4����p�<���  �9��C�Y t��T�<!`!�� �I��h���!�iBN�<�0K_2j��YA %A
Z�T`�@ɔK�<a���<W�N9c�*ؚ#����� YK�<�F���a{z�6��*b*��1�TK�<	0�S\� 0�+IƽJRFI�<�������)���[����j@H�<)6��B�誖 ̛-��,ʴ�VY�<9"�ZJ�u� �N�=�Xb��P�<2*P�\,�0�SC>IA�D�0�O�<YB�Ԩ:�1�7`�5V��0DN�H�<�ԁT >ƭ�J��K�vPyq΄G�<y'bׯ^:ܱwoȹ����f�YE�<!2CN�j5|�Pٰp�<2��3�y����aBP��jwTtZ���y
� �X�wkSU<�ťZ��0-�Q"O�(*פD�<���B�\�.`�"OVĠ��{gĸ�d�w�P�"OޕFk�D��D%����p"O��c��9>+$H�3�Z�t%�w�O��[%I2�)�'lr�O�B�D���2sr�0�ȓ{5�S���w�}:��O�D^lp�'n0	�p&���$��aZa&�b�mA�l�\x !>�O.=�'�N��ԙ1��5b4E٥���@e8�"O>���N[�.X�lrCNE&+�8��'\��h���ӄ���Q�J	2�T	PT�X�kzB�����ٕ#�&S�ft�#EG�f��C���2m11aVg����)V�^6�̻��OQ�C�� u,�:�(���Vb��5�� a����ش!T] ���sy�+\<"�QRq�
GOd̪!@H�(Oޭ����:5�0�*@��vk�i���'VԨۃ)E�@*ĵY�G[6/VHx����F|��yv��ba+(���bԧ!�����϶�uaP0S�U��j���v� &�ԣ�W������Bv���ӆ��� K�1�-��/N3F9!�DEO�`T�s�]l;�[t�!n�Tu�`	^�^'XÈ{ʟ�Yp�.�N��b&����ϳ3"Z@)�G�
Q!�D��"�TA�bң�xhp�͌H]\�Cr����怃)mP��j��
�@Mx�剘_7r��蟜X�V�;%�ž����� ��h���	A/v��Bԟ{9(!9�$B���m��'ʔ"-����C�"��$��6�p>��
 �4�`e�?'&`V�L\~��t��,�$AL���S) J��h�=�';|�G���/^	Qq̅�eW���ȓL���`O8\�α@WNܕakF�IŬ�m�v��3�,�)BSF̵!�F��;.b�a�0)�J���ǀ�����n�b�C&G_�Xd�	;��M�>�Ě&N{~r
ϫD��Ɋ5E�6H���\Z�'�а�u�YJ7j�R"��y�1�
Ó3O�Q�Uc�2)U�#���%����a�~�bU"o�fʠAy�d=O��=�&F"q����F?}T$��f0%�,�!�n�<��� ʰX�G�;9���롃�4:�qO��x|�`� �� t������� �!�䚃^�p���R�|� "�hH�8n�`?@�zEf�O��'��#Py�AA�w$>����G�r��B�f[6|��	�'�>���CB�	;B��6��'4���Ecުj�$䘴++n��}A5'�ay���8�V�*~�2��π�L��-�[(���D��T	��YǺ�`�=��5�0�7t�iwG�R}��A�y~���ۓP�kV͊�|@J@`�LV=*+�u�'�d�V
k�S�$��UW:��X�YyX��#ַ����MRo�C�ɯ4�µ��*���ѧ�C�f��O( ��G�x͚����f���|��F��ݧQ���놃�
9h$���'4����#�-6}���aee�������`�ϊ�X�p!RR�|���i@�	)O672>$K��)[�:�����X������Ol,� 
��MK�#S�6GB(�(ѪB��=�#,��4��$�+ �(��/\ON|� +>=�:x ���6O>!�\��K���M���_�S0�H��O���W�~+�
>��)�G�RY;aM��!�$ð	$����CߣH��i&n՟7�6��8�~�y�'bV�$�P?�S�6��5mڿW��� �5g�I�z5�5���I+�ab�
8�2�
TdSik���R>}��a��
��H��y��؂
\=��Oں{���=��N8g����-�9iի�P�'J�8!�Ȏ.o���ja�Y��EH�4+Вڤ� ���@
B -�%ɠj�bta�L$ ��dV[B��%LP��$(��Bg�I�ق&M_��87���m���	T?1�'[��j`A��� "֗v���H�"O�9��`F�l�a�/�E��j�f�c��`?Y�'���O�,T�!h�(à�]+Go��P	�� ��2��@oZ���D[��9+5�/
��P���*��p��+�u?�'���1��ۏ8�J��r�rbS���'e,z�ޮT��d�`�Y�P�\ ���:8;R|��Ar�r���
��r��y����gN�cqb��K=`�dP�Gl*7��!�N��t�7lO�m�فQ�2%�c/^�h���2%��dHT�N�vQbBB�mb 994B�O����?��9 -\�bq$̃wT��IϢ5�XB�	�Q6����òi8l�p���[�P���qY��{*�V�� ���p��WoQ0��0xX#"!��:00�idI@�`���P�]�d�0zB�>I�
P�PI�c��&t,����`��I�(��z��%�E��v��ቤ �����%�g�q�`"a�� �5��E̮q@M�@Hht�b�/L����cĔMT����)O&}���*�M����U��	��� �$��h+ƀQ7�ل/u������MA�#��'��Ԯ�2C7!�����m��l�m�Hx�KV$Z�� �CˆO6�2�T>��&&��4d杷=!>�財��(M2��òU�BB���}�>8"���H�:@�&�^��q��B��!��� �"m�TP� �'��'�&=���9B������bk�	Ǔf�ɪO�-�!�Ȅ'���@f��W�Lٶň�S����%Q�,�6m�v�T����*��Am\�B<��e�?�J2���&*/ʧx��ͻd,���R���� b%&)��fn��)]�`��@�U獚�E�i�������Q�jX�E����b�Py"쟑j�`��j�T=ҡꜽ�y҇$"������fpDt��y�T��Ԣ��_2l�ٳ���yb�_<�F	��c8$�
-����y�)O
Ɓ{�
2�Bٚ�B���y�O0|��2s�͎�~�#�ص�y¢H<J�-"j�>k�љ�8�yr��vi�=X�`W�d:�@ �ͽ�y�U�F�PHc6��Z�*���#��y,P8j����냁UXf)�&Ė��y���k�h)S���J>(�@FS��y��8t�X�����Jh���@�M�y�e��hObXG���A�4�g���y��ׂ?���Ph��l?���F���y��Z,U�1o4�҆kّ�y�'S+Wy긳�A�
&j��Ʋ�y�gE+P��`z�l�iʢ�������ykăm�J*-�R�=z����y���$�䍋.V�zW���m�y��\�?�ʤ1���<p����BK��y2Hː*g� �ʑ�p��.��y�͚�xCٰ���#+��0�D��y��1ϰ\���C��y�b�2�y�I*U*(p�g�ȟ:6�Վ9�y�+^�c�l��@�v�\H��%٭�y	Z������|��HD���ybk�?s󔔛��_�t�"�2���yr�N�}-� ���^�sQ��q�U��y�ĥqK:�"��93�i�A�8�y�mG�j�mi���"��=����yR.ȾCE.��� �%6Ի7��/�y2f�u����0�A��v8 �� ��y�#��(���ݸ����*�y�Gȱ9�H��̀TlE3a��"�y�j�i[�e�M)qk Ѡ�K���yB'�j����!T!�H)�w��y"�� R����X������@�/�y�A �d�C��9�f�� Z>�y����ث��S�v��-EN�"�y�,R���R�M_�gj��ᮉ��y��Rb�>�4�]�dAѭ@�yb`�Oz���G�3XA�A
�`��y��5�]aQƃj�hb&���yR���P�p$���^#�hP`�C܈�yR��-&��/0�������$�y⅄3�y3���;����L_?�y2��2u�ș`W*�,�����O0�y�*�X�$ ��Ԝ �l"p(���y�/� ^&��	��د{vq���\��yB���$K��CV*��Pr�@��y�m�
(�YM��:��f��ym��Z�Bt��� r@�d�A�y
�  Q�Ŏ/�$�0"O�21��C�"O� ���e9b���8c "OF��iX�ob �*�-BX�Ma�"OX ��M��(S�gӕ*MXѐ�"O���(]*\���915|LAa"OH�Q^Jά�qꉨ-*p-+�Kۡ�y��L�
b��C�'��Aʐ(Ѓ�y�F��2T��%'oj�P��E��y��0rj�	��+|ܥ��&���yb�נkp�]��*\8:&|i��%�y�k[�@�v		�>-rhM��y�f��Z�깪�A��赚@�	�y��7�0��w����0W�!��l�=RA��� y(7��1
!�D�&�*���.N�z��#倈's!�D�8E�X$Ys�W�E� ɩ�Mř
!򤈦*j����\,�JV��"�!��0r��-�l�<$1���;�!�DWy� �᎖U���a�.|�!�d�,F� `95(܋9�L��pf&�Py�C��L�ȥ��]����-^��y"��;��hE��;\k
])�)��yZ���:aa��n	♺��5-jf<��x]�� e�%Mm�q�'¼��ȓM�ԃfD�8gi���I;3^�Ѕȓ~'�9i�*�w��R�B:(X�ȓ\�`��)� 5nN �'^�)��-���C_�{���y�CɑP���`(A�^�h�	d�-@��ȓF�� �GH�K��J�Y�b��ȓ8H|3"�9va�u1F�)<*�|�ȓH
���6���k@�
�kȤ+NU�ȓq�`)ɚJ����G�J!=ob���K��vW�FG����S3P�J4�ȓ5� ������ �2"�<��^�]H�I\*����10u����� ��7h�(��A� �.
҈�ȓH�R�1�I�}��P�֏I5+9�Ȇ��Щ����Z�!�-^�&�U�ȓ��D[e��q�4QEd-Y��u�ȓ6��VIHV�
q�OF�uv��ȓ/��E�!
5�\p����Ԩ��}�Py���;�2d* +х���	�B��$V�#��;��ȅȓb��1U���RQ9Љ��Uc�q�ȓB!~=�D��;w��2fǱF �=��Q�H�ӥ���=k��O5PL�ȓZ�BQ�u�D.j\M�r�ʳ4�d��ȓN��U
0n.����'�_�WI<���5��l���l�*�"+H5a�m�ȓz ���U�ZKR=[��ݭ<�8��%z��L�y���Sm�*Xp��ȓY���â�A����r뀨E%؉��v�L��������i�q�޵k$"O!�uм���	P�
���p�"O�j��D�3��i#��(�>��3"O���� �.>n�e�2��jl��;'"O�M�S�ҿo
��z�eM�!kR@�"OD����z�|�"�c��m��cq"O�����$$4��eɍ�ē�"O��JE
��t��i��L�:��r"O��P��^[�a��e��Ӳ0:2"Oj=��+���d��JR�Y��Q��"O:���웞iL�%���L!�6��"O� � �5K���*8G$MA�T���"O2�*'�0E�0��V��Yܒ��g"O�� �L�m��h<��z�"O~-�aM�0�q��*�<i�#"O�S���l�$婓H��+h�I�"O�anŷ�:MP0��|���k�"OR�Z�H�� ��T��eY#/��"O��KemP.��i#�DB3h�e+�"Ob!�sm܆ �%Ғ��5�0y�"O�������8A� ��n��A�"O<%2��u�Bdg$P��-�%"OMhӃF���ܾ���"OXXD��M��A���P��ъ�"OR�9 �D�EXd�zsI��
g"ؙ�y�T/K,1$`T� � ����y��ފHD R(Ύ9���P�ӯ�ybOӳjg΀+�R�1��@#��yR�صMt����.0Ԙ�; �ڳ�y�mݯ`D���D�+�$pR�̒�y�M	�D���*"�Rq�}�<I�/Y�T�>QC�I�A����
W�<i�eF('�p�:eeOn��97�[�<��"K�M�|"�"E�Pp�m##m�}�<�ԌӅ>����E+�y��	�Ιz�<A$���XSF�#j�`����p�O�<�E=V�ȣ�(6�*p�oKD�<�(�������Ũ]b��S��e�<���N��8�#��M��!S��[����<�F�UB�ܱ�B��$����]~�<��a�/b�Ĩ���t��2�%�v�<��EH���!@�˞7y
0)o�<1��$�X�0쌘(/�
Ҏ�1�hO?�N��M3�.Er���Qw��6w�\���2�I�G�xy 灇Fn��5�Q�:C�I��~�!h�&]�X��c�"O�9`i��x�&0�F��?���B"O@MQ��]�o����P�E�����"O"� �\'�,+#e��9V,Q"Op-��BOe4�Dxuꆕ}R��"O�s�j�e�IP�'ń	�Xr"O^4��BK|!�j��	:i�m��"O��p�J�(��1�1��0T�R�"O�`���2�*zpgZ���"O@\�mF5|Ln=�F��&(Έ\	q"O������:Y��E�%�)]�F�A4"OF}��R'\H����k�xe��"O�}� Ɖ!��d��Dߖ4�z��"O؄�ƍs ���4�� i����"O�IS�Pd����E�}�F(F"O��)�'D#o�P4�ŭ+�P5Z�"O�q��b���EU0�`�C"O SA�\1U���0"C��G����"OXT�&T�2�kB�߉�6�Ҥ"O�i�2��]�^q�sG-ʼ�sE"O��p���;��}iRiYi�\���"OP ��.C�S����bhZ�X��%c�"O�q�X�Q�h��-ӆO��"ObX�a�ff�,�Ǣ�
H���a"O�����
W��V�EM��"Oн#� ��v�2]�V+�8D�U�W��˔�)�'k_XHqE�(&�Z��q@�~�l���fx�ջC(c���`��g7�4�ȓu�����
���(>&���A  ��I�+��;]%��S�? ]��H>+�Ո����7�r�4"OԜ9��S�E�~�I�hC�~�N,��"O�g�?Yn��2wEnfhpcw"O(iۄ�S�`>�D%C�>J8�۠"O̠I���.A�|X�"ώ?G3�M�"O
����o2�娒*0�,ܲ�"On�k�A����u�'��
��h"O>�"Gr�D� ���s��xr"Ox9��4�ĥb��ļ���"O���¨�<0YHe�C��a��)�"OP@�%�g��<kʌ4�.�"O�@�e�F�k��<I��D��^���"Oh�+�Dޗ<���8F�A�#���w"O���1�-2�p@Y��	��<8&"O(�w�G�"����W���Z���Z�"O�<�6�-47쑀�F� �V�s"O4�Pd�R	� ����~�>�zc"O�ò`˾$�VuZ�gԩz�0ȁD"OP�v���jL2ux�ٔh�e5"O����+H��@���B���(q�"Ox�f��7puQr��>Q��\r"O�)�%cBr���	A=?G0�U"O^XY5$O�>6e ���
4�Q�g"O�Ա��!@�(���r�0�%"O.����I1@�㕍���p"W"O��PH]�R��i�e�_�v� E"O�<�-�!Fe���Q�uW��b�"O��(_#l?��eE������"O���D`O*[�HY�"�N�(q��"O�PrDF� ~��Z2!H�)�T=0#"O��{��*E����I\�	oƝH�"OP�3�n=S{~$Q�h��WǨE�%"O��V�C	�����B�S�\%��"Oh؃FK�-I�,eqׄ�/X�:0�"O����.�7|�!`!�ΫW���� "O(��4��%|��Q��X�}k����"O�X9H��?�xE�Rk�W�}:C"OX@��ڕR���e�_;f��I0"O�x3�V�g���D [�M���Ұ"O������ % 0��^�와�"OrÀ*��/��Țs�Bg x�(�"O*�@D=yV�Y�@�[12g\<�F"O�=R�*�1H@ �1+��-M�x�"O �a��	"�|A�dJ&_>�)�`"OB�k'}rh���Z�6�Q��"O0PA� -p:��ЁJ&^�B!��"O��JdZ�qʠu�#ϩ|��7"O�T����(*:�=�A�&A���4"O�$ʖk��D�x@ Q�0R�"OX���lQ?@�V����Q[x���"OD�S7_
��a��/H=T�I�U"O��h��+�&���,?��U�"O�M��ƏS���q�C\r��Q�"Ob��ׂ�5l��T��#�)Ⱥ�� "O��(W��1��b�E
-��(�"O����$��gaפ$��	�u"OHu�����x�2�yV��$����c"O��2F	��O��9R2��`v"O���%b� Y+L���A.	�R��	�'�D����*���RC�KV�I;�'���P���]�l1��%A8�(��'P��� *�=����D&����'��l)3W0Oq�X�\:Om�$`�'�+4V-i�^M�6ę{� I���  qy3J=2H�yU�'3��"O�t[��`a��Z;}�=��"O�Q2��z�2�i�h����"O�X3,�K�Tu��(� I�Z�"O�)�Sh�%��ś�gQ�y�1)"O�Q+S�yCL�z(��h����p"O<����ɯk��!�l���k�"O>u˷L@�r	v�`P��E��÷"O�=�0-_=K�N9� !^�dX5�R"O��kD)�.�Lł� r�d�e"O0�c�K_)��]#����&pk�"O*(��Fߘ(�R�	��Y��P�"O@�Y I	)�tL�3�Q�\'"Ot�4LH�B��u2'��7`Z�%�V"O���H��t�"��e��
�~M�"O���E*��~:-I��
)eJ�"OB��էJd�x�k̘qr���"O�̨�� �J�T��b	$Gp�A"O,���F:Y�!6��.a��:�"OR�8׎� Sn�h�۟{`ˁ"O���pdF�c5li�WeݳQW��p"O*�*Q�B�7��`b�#3����"ON�ᚈ&������}��v"Oڂ�5̐!����$�K�"O��2S�M�_!���,�1�5Y�"OtHB� �<9L��+%0"�U�"OP��@e�%9l��Z��xp9�"OnE��#f�8A�nG�v�D"O� zv��kb�EcGΔ|�
�"OTMy$�]�_�lk���X"O4	5c׋[����wm]�,^X��"O�4:��,�%�Ȝ2�z���"O���hE#O����O��s4"OT��� 	"�T�iȂ��P "O��#���'7��kVh/
:H��"OTuq��$XrQZ�H	5� 2�"O�]���l�ʵ�q�H�	3 ,�"O��Va��K���Q�u?����"O�A�Bwad�݀GY���CƉw%!���sԄ�9�ω�R�Ų���8�'L<-Iv`[�u�t}p�@*	��e�
�'������+q��\�7Ύ
}@N��	�'ҰI$��4U+�=`�@�;��H�<���4_S-��ʉ$J	��Õ��O�<�Uf[���@���"H>!O�H�<q���C ��/V��,#�j�<SBU�3��r�ep���m�q�<�w%���	�c��d�X�k*X�<�6��ZW��3ՠ�"Bh6��\�<���_x@�%�g�x���B @�<9%cѲD��h��`�{	`�Ж�w�<!R�<^K�E��É"h ��	p�<�̚K�����;G'�3�F�<�mµqeB$�� VH�!	�	~�<qtO'MB	�£�<shfY�Uk�}�<Yf�	�
��TIf^�Fe�|����{�<1a!��vztS�KH�j�R	+T�
u�<�ToR�AWl8�����B�����m�<��Q'# �=�U@�XG�@�vGo�<���M\\����ъ9�:���i�<��ꁦQ��)IUM�/;!���P�Ia�<	F�	*@VK�fH�/6P����JC�<	ABù=�$ȀW���9����R|�<q��
"�nͳ�-~1&����y�<� h!Q�S{��a0�Ô7��P"O̲��J&6rX#C�R�p��"O�Y�S'��5���/n�J�v"O��0�E?Q��@B�Aص]�茊E"OV���%܏Tv�ke�ߥN	޸
'"O�T
@l�d��h���G_����"O�M�SJ�7BX)s�K�3=�<���"OD��0a��U�vQ��_L� }9�"O���#G-� ��,ȅ
����"O�በ���-�����y��drd"O�y��5�Vآ%�U0d�k�"O���Sf�jL|@OU��zr"Oi�&���H!��K'a��Y;�"O�iFR:zEꥃ���J�p}��"O���[p ��u��'߮D�"O.�kD�R)H�(ge�Ln��"O�}�GH�6!���7�DX����y��X��X���hO.W&H9�aY�yB��0��9��,�x�I�2�õ�y2���P�02рc�!�G�'�"�;�'�ȉ �A�2�v5�ƪ������'��tC��%Z�f��E���� 	�'f�@p�~yNub�>&��;�'�X����W�
M@ �(S�"w
�	�'��3re�7Py�PId�-�q	�'� x�OˮNK�ǴGR�#	�'�d9
R+9ˠ�ñ��!����	�'[�����@���Ԣ�+L�����'�TLeݽN�Ԑ�����x�'�<!�)�(R�&:���+��'��`�G.#Vl���S�l��@�'|��y�B>��McG�hZ�'L��+r�ŮK/Y�Q�4����'�����SP�6擑1�䌐
�'\�<��+�GC��S��җ-���
�'	��q��	+��,��m���Q�
�'M0!E�D�>Q2�F�D��
�'dD�Q
$"D4�j\�Ǝ\�	�'�NH2��IT^F����ۉ>-��h	�'�x�Wd�^ \!s�]$#la�'V�;b�A��$Hp���\(z
�'�~`c��E h�:Tq�ʿ����'l�A�T/�8p2P�pB�-���'�՚eዬ#�2�S�J;t�h��'�b]R�A.�n��2�÷24*5a�'H���C�3��1� Z'�u��'j��4��:�T8+�oJ�%!�M��'y�}��"8:鉔�V11g5��'�����C�-�	P5���=����']��BȁGK�=��i��3�DY��'�$8�f��K�J98a!�3�%CQT�<�2k	�G�t��h-*j�@���[�<����'
S`1׍^>z�h`�K�A�<���Y~xyV�7����&�ZG�<�fE@$Z���9W�L�]i�l�Vh�L�<1B+X\6,�v.�qKZ�2�RB�I6.{h�	B�r!R�2jA�v\(B�I�]�!����3;�����jYApB�	�w;��Yc��w1��K�h��P�C�INp����됯?��	�wh���C�I����+����w�z!�fMP��4B�3��9�"�-�@Q����%�*B��68GHd����B��jq���m:$B�	ir�B���>�AR�	�^B�)� "�:DO�S�I����$%��K�"O��̓S� @�v鋽(�ݨ�"O��Ǫ�==�QX�L�Dy�v"O�͙�#_�^t�P���K8 ����"O��4}��ܙ|r���dG��y���?�J��GҰu��qU*��y�B3�A�+u����n�>�y2�]$Rx�	�b�)@
�k��1�y�l[;V��*��1ǐ�qh�m�!�d˵��t�!��)T^H+ ��
�!�DE�q�����ڬ�SR����!�$_H���!"�L0H���{t!�D!(�y����g��!��3N!�dۊ
s��R���Qa*�S���bX!�Q58 ����1*�����K@^!�$kTr��$���T�`a@�ۭ!>!��X�\G�������:�ʃe�
q�!��S�%�Q�A�4���::�X��'�ν#F˔�`���%f|n�`
�'�|�QD�>�qB�
Yt�r�'+�E�;x���S�e���W"O ���5�P�*�� h.�\S"Of��e�*%��p���A��Z�"OYz@k�Ag�
�MB� �L�Ce"OT-���4!���ㄖ}��(s"O�]x[rD#bZ:V�p���y��"x�H�Af���\7ʀa@$�>�y�r`�
����� ��y��C�%�T��aND�HaBիď�y��E�p2������2�x���x�<�􊃴 ���)��Ēa�r��t�<Y���dl�5�P+�:UuD����n�<�F)q+�T��#U0��=��`�p�<Y�K�L3��1���>e*H��v%�j�<6 f�>��G)�o<RH��Jc�<��mz/"�*����$��t�%�E�<&��K��K�,	z~�8c@�<��IS��U�u��]mn��Ц|�<q���E���V�צ_�`;�Ox�<����:u�l,bbW�����'l�<�b�������4��ABU��<�y�	�7}/�$;c�'3P��R��F�y"#�.>��h��`��.�88Ô����yb,��y%��uj@��8�"�E���y2�D��ͩ��D�(��&$�y�k��ъ�f��b&��9�y���M^��kէ
� �j]�VC�		{b�l�9�� �`���Q�2C�	��v� �n�r���0�2%W�C�I9;̀M�%'��m�Rܹ���i��C�	�0�( �!@����v��'!�B�I�3di�L-$(J��J�vq�B�	�#�4�A�4N�F�K��Ћ`�fB�ɘ^+.�Swn�	:��R���B�I�Z�`@2�N���@�c�34�B�ɩ=�`٦��{��{t&I&�B䉓�ɩ�@!��SӍ��.�C�	�նU Gꁢ,�|�$�����C�I��ꥢf�@TfP!!'��&��B�ɠXqc$��Z�F�
��	��B�I�H���B�0+$~+0̍t��C� 6�Be7�ZRbZå�܄s�C�BFы��4#I&lj�YG��B��2�M2�c\^�ppFM��u��B�)� ���t�%�x��ԏOШaJ�"O*���:,a؉��n�&C��tK'"O�X�l�+M؆\���S�&Lv��"O0�tL��d� �9�LO,I�~q�"O*`It��!!ƀ����8[  � �"Oh��(<(��ZTT���"O����={4,����̇R�>�`�"O�����Q([A�r���O���1"O�p�e�/g�b8q�py:$[C"O��!�*cC��d��cZB|h1"O��Ѷ�!�3�c�!A���"O���@�&��p[C!�"(��8r"O��@wE�ܹxq�t�-�"O���G��}`��0��>�bq�0"O��p�%�
d�>��ɴ)D��3�"O�ы��� ��så��{V�ɀ"O��U)L���rg" q� �`"O��R��$Z�F���T(#D���@"O:9r�Ύ .K��
K, ��U"O�#� 6I)\8�׉��zn���"O�� ��"����b�H�N�� "O�-���6<�zp١a$��9�"O&���iQ3l���ub�5��E��"Or����W���Р�9h�HQ!�"O�=еǛ9`� ��J_�i{�A�&"OB��SH��[�.xqQ4c.hZ""O����A?s� �ZH=	�ŉ.c!򄅦�ܲ��6w�4��椓�X!�$O_�ِ�@"!y�%��c��-7!�d*fL���q�MBf"�!۝K/!�$�<�"Lj���>������.�!��I�W�<�#F��5O�l��k_�K�!��)�e���K��:T�ɐ�!�dB�-lYQbI ?4����$g�!�DԀ���f�O��(C`P�*{!�D�1xZ��Ʃ�b��p[���a!�d��8m8�n�:�P�A��?!򤙐H��4�0�N�M	�L��⎠&\!��F�F�
7�͵~�p�2�K��n�!���&J���c��O/<�jp	��	�!�$��d��������_�;�-�H!��t�����M8�Qx6LJ�Rm!��Z�YQ�-\8�~��:1e!����h2KV�/�xI+S�ެ6O!���VXt,��RMs������/n!���u2L��m߰e8J��=oR!���쌺Ў�>��C�Kĵ7�!��-7~) �N^�MѴ�[�i}!�d#�l��b��B��=�AL��zm!�քsI"��C�ԋ/|�db���mQ!�Ѫg=z�0��8']4 '�&?P!��&��R���:J?���ҏ25G!�d,P��h�4t���"O/j�!�إJ�@����8l�.9��۟>�!�������|��ЂT�SV�!�$�#3\h����o�p=�`��&\�!�Ć`�rek��#�XSQ�q!���Y��8z�!�)q::J� [�	�!�dϮ,ƺ`��NӅ_���1a�t�!�䝃WT��*nҤ-��A��*�!�E2�#%���D��n�!�D�~�H8�*]�1����(F#�!�Ĕ�rav���Q)Y����.�!��A��]���y����J�5\�!�� Q
'���l��i`�£g~u�a"O���C�%w�l�Ƙv|�c"O��C�X�8��е���	ˆX[�"O.I��ώF�M�0�T���0��"O^�#�JT��؁�T�B�\�V|R�"O��T.� \� �p�=B��Ȥ"O���T��	`Ⰱ��,	-:��J"O�HcD��	>h�J���"X����&"O�5)R�Q �ʄB�=&�a�"O��H1� 0��)�I�+�I�"O�t`��ŎMޠڵȑT�x���"O�i iO�:2j|�h��%�A �"On@kuk�1`td<�S,�=�V��"Od��"K:�� �4�ۤ���I�"O�H��HU?��ژ9�`��0"O�+�F^<-iԎ�:�d5��"O�@��%1oϒ��an��y ��"O����S_�@x�r��Q{�zQ"O&ܺ@KK2�Jx�D�,q>��b"O�XH5�*c���S-�S����S"O����B�:�]� b�m
2��"O�!�3�V��^��$j� �P��"O��2�*lVX!j1�@0�i��"O�:��uPl���MïRz��"O���GW������^s@8
g"O|	�%ĕ?�~`�c�]+5�4m*�"O����E%R�� JM�0���g"O���U �	�1b���<N
B�a�"O@�8vCƀ �z��픚�KW"OA�g9z��-���ie�ͦu>!�d����i�PO�5I:4	�	\v]!�䐖�B�:�-�7/�����:�Pyb͌8B-��9��ӻp�p�����y�H1)@p��ɑ!p�}p3����y�o���`�3�l�2��QJ㩀��y�Ţ�Nr�o��]<4���H��y�d�6U{tu��
����Xw�J��y!�6+�E���$��vk�y����J�+V)(։�%bS>�yb#ӏ�2���ę�	ؕ��j
�y��Sm��]BAiE�S
���Y��yR��?b@����1%b#�y�O%
�⭓+� ��	�4#U�yr� �3��9p"�_Ḙ�$�T�ybj #����_��p�L��y:2�"�)�.�e�<�*��y�YR���Qa�Ƅ_�F�1Fk�:�y2 7ܝ��b���M��y�Ef�D9b	�!	$(�d)���y�hA�k���(�|Τԩs�5�y�+Jg�p�Ӌ6uO��r��y�X6 � L`�r|b�##�³�yR,���m�`�l_��c�	�y2�<j�` {PƋ�1Z��:� �y��� �4<��ٔ/=t%���Š�y�Mu<���� �'�1zS�G��y�B2c(ɹ #]�m�V�� ��y"�9C�)K��͚c󾤉�BI��yb([��.�d�W�)�i���ǚ�yYP��1A:7y~�Z����y�뇇ee���;�bppq`���y��##���iZ9B�0��
C�y�HQ����{UDK)8��=R��Ľ�y�I�����DE�`ŉ���y
� ,�� K�%�.B�T='��(�"O����$r��r�'G	@��"On!	*Hg��U(A��(T�4U�"O���Y�T]�@+�i�<%��(�"O>Ia� �{� WIH1K�$���"O
iA���+�D��'��'�\@@"OҠ��'K���3�,F�H�t:"O*Tc���=k�z#s�$_�l�u"O��yA��<m�Z�kʡ%ڢ�:s"OĐ�flϏz�h�K:�б�$"O
@��֐.8Mr��J5 | �"O
`�5e�+���ߞ��"O�ણ$��[&Yh�M��t�j�"Ot��I��88��B�Q3���D"Oz�##��?+p0p�*�$�pI��"O�)���;%��i��w:\�"O�ᘴ�B09jljÃ#h�a��"O��U@U(gR!�DaU8���"O\(�S��&t`"`F�4?<���"OL���'\���Umߤ]�9B�"O �#��ѕ V����W�V�6p�$"O�\』-}W��E
�6��u"2"O�t�àT�8SDt���6��I:"OF�J�nջ���`�$�6�z�"OBq��	�g^x��"�.����"O��Z#�\��Zu�+���p�"Oք�冕�[�X�1' �.qo��"O������8Q�� ��[<Y#Q"O�q�P ��?���[v+K&&]E"O\��g�>%�f���<����B"O�x�J�#!�A�ą	(�x���"O��z5�� 7��[3��d��+�"O�!�&f���C�+Pb�P�!"O�4#�������e��w�(0�@"O��#�![?h�1��,pxX�"O49���۝� �:ÂC�)S"O����oS-��6+K�%���"O �q�M�.��uP0��"a.�
�"Oĕ(�ۛIHT|
G.�`�x\��"O�sfm�u��l9�_
p��iS"O�4�u���	Fȭ���w�T�hw"O����_��R�8GO�7d�]{"OfD֣w�>�k7*Z�k*Z�9�"O҄����:����'B�,@"O"�`�÷jdI0E���*\��"O�A�E��3L|U��Y�(�"O�j#��)P�!z��;h�}2�"O�Fj-g����&]�k�\�#�"O"��F$Q�P��mHʘg��h��"Oʄ�V��h���(6�?s��� �"O&Y���^�-����`י�t���"O��k0�¦w������/z��;P"O�lr��>G$t����4��TS"OΡ�c��HDΈ놇�s�p��"O�(��)�!T6`\����6��x;V"O +�����%H�6��5[`"O�`BQo�/Ԗ�ˀ�Ia�2}��"O���[�<��e�Ԥ� �J�X"OF�Y"+��M>ll��(�/_��1�"O��z�G�%#`P���gٕ,K��r"OB��5���e?��R����#�"O�4AV��a����ׄ��Mp�q�"O8����4h����o@��"O@Tr�]+i�$�r�J�ޚ�@�"O� f��#HA�0۶iŉ7Ĝ`2"O@��q��7F;zp�a�Ϣ!��̋C"O�y�QB'F�@��5\���V"OX��Nߤ����n=P5sA"Oz�¢H,\�̡4왯/ˀ�R�"O�� ��ǿ�N�9����,�S"O��0�9|�Tmv�[�w8��4"O~����N<)��s���v����"O��s�Q����2�H7���"O���5��~�*�cVs�.١3"Of�SP6{�v��СZ�&Y�<�"O�A�wK�)��Xa'a/&Gj��"O&5��G5�x����7"��p�"OzIU 7_�`�&�J.c�"O"�(��ިbԊ\�p��T�P�"O��@�� �[b�+u��J|��"Ol��DKI�>y�cI�|��� f"Ob��(�?�����_�2���"O��SD'<�RhcT�
Q�,�s"O<�isM\�|8��!sk�:�"Ov4�1)\7R���Z���"'�1�"Oxh�gN��T�c���/2Z��*OPi�MQ0ְQdF�
�vx��'3T���ʖtR��΋���P�'�����Sʑ�G@Ư����'�2�I��ȚH�L��Ø�-;�'����I"~�{DTJ���4�B�	g�Б"i /qV\�fB�>B䉄:���H&iо"���Ġ�fC�ɱSuP�� [(1 *��ß@%�C�?�h�Hv�W�GԞ��#�b#xC䉿
<�R!�78�LJс�t�C��$D��y� I�t��P5"�MK�C�	C�|U�`�R(J!:��oY! pC�ɠ
;�y@$B� u �ycM��TC�ɭK���1#��e��8S�,C䉸{��IAT�͗3�d�6O�2K�0B�I'{6^�E��t�ٛ���+�C䉆HkZP�b�Ww����� O�C�	&;՞ ��*
3�G�@��C�ɨ?&j�C�7Sv]��;�pC�I��y���#�Lx�啗:ÐB��<ka�D��M	50�|Q�Ȇ4��B䉰*�Bh�!*Al�T���
Q.+�|B� A�^(���ܖU�`%�K�2$�B�I�����7_mr>Eq���%%��B���9�`��>G������B��	�����@��,������2n��C�	�7
��Bj���΍i7Y�%lB�I�����h^ް�3եZ�e��B�W�4S�!R=j�|��`�ڬ��B�1NI�dpg'A�/�}kG��ߪC�Iͨ�3�O3o���hVcD��C�I#*���!-�i�u
-�C䉴'I��s��2�V��1ʚ�L�C�IO��xI�FV�.zv���=d
�C��0۲�0e�A�jͦ` ���C�5M���r�I�+=���[�G�\C�I95��͋p�_#,tp8�(ىZC�ɘ�)q�>ix(l�� T��C�	�\�jp�U�W�Fa�⑉��C�ɽ��8vXbKZ�̩R�"O��;F�ɋqz]�ǂ�p���sS"O�4����3� �ժ�MfT��"O� pT�E��-`�A�)��H!"O<kB k�8L��h @�:��"O"I���6��$�r��N����"O���1jӒ=�X�RćB�0���� "O|�K��;!��	���Hx�<xjS"O���BP�?H�5�D2yz��1"OP�ۓ� �}_�j�C=lZUX�"O�ɸ�I����
7�;T�r0Q@"O�myGBƮ6�� �#IڝA�"O�d�!�T�H���CMd@�!"O8��Σ:+0�A���#�j�h�"O |1$�ʄ8�p�s��O���J�"O�9�K�uw(L���7VM�y�"O�IJ�S�W�$ɑ���wG~QA�"O� 1Aƞ��@��h�>Mv��"O\e:���#~o<���&Y���"O^�#٤����v��a�&��5"O*L�/ծ7`8(Z�MJ:�d�ȇ"O� �G�
J�T�C΅C�Ȳa"OP�pN"`ںI#���+%�,8�W"Ohyɷ�@<�l��$՘AQ0��"O�S�g�+~�<)墋"Z?��v"OȐc,�h���w�β��}Y7"OȰ��"�A䬜����(J�"O�ݻ�$Y� 9���wH�js�ط"Or����D�<�0�ch�)���"O�$�e�V�Ͳ(H��.mQB���"OL��C�D
mKT�@C��"O�Y���X�+�����i[ c?0e"O�k�)�<D��`��U+v�h�"Oz����X|\���MN�&�刓"O��0S��<6���>=��P�"O�h��)�?_�|U"���KӲ�Xg"OR�[��ςD=&L�1ퟸH�x��"O0I��B%���l߆Y����p"Oؼ*a)@�]� 35&�1~�jV"O��z���,`J���y�%�"O������.��	j�Cd���ɴ"O��S����!ӖCȬ$,��ض"Op�iv)\=CŦ-�R�P%n D"O,�F&D_�}I�C&T$����"O�A��NN��+�Cτ@����!"O2Ԣa'C:}���zS��f�z�"O�B��ÄUʈ@�����B�a"O�y�.ӌX�0M
�ΨC��=k�"O�([��M
��;�H�ʤ��"O ݻUD�7Zh�`oA�����e"OX���X2��P��,�0<���"O�݀��� ��$K���M��5"O&\а!�JO���.��3��%"E"O�\����6ec.Ӑ{H�c3"O�@�#LD�ĵ�rF�p��)'"O$�z�GT7h��4p�ۄBj
0"�"OXAJMW; ?���&FoS␣�"O���7a��@���Ƭܩ?GV�Q"O���,S�4���A��֓8r�#�"OrL@&�"0�L�tI;o��h""O2u�E2����d��9L�*�&"O�9d�͢s�L����J�X�^���"O���ō�s�,���t�~i��"Oڱ@3� *ZR�r�lH���a"Ox*�"W�I	8���iӍ���U"O<�0Ò�Y²|I3��(!�nAI "Or)W�s�es%҂n-��
�"O� ŸS� �E=�u �j�&/0܀C"O �q�2u��Q*IH't]"O���q/_-T��a�d���8��"O�DK5`��I<��� ϒ+�r�0r"O�}�m�$Рai��u���@"O�L9p��;Lέ�'"E�fp��"O8D�ʀ=Ƞ}�0��8'�y+"O�`8&G }�(M�ӥX���+$"OzUPQ�Vi`T�X�Yy`9��"Oص"֥�!=��Ê ,Z�ֱ�"O.U����9|��c�7>�$�g"OJ�H�J>7F2���(Q�Td��"O�aa�監*���#~�<iУ"OH��Ң��vrf���B��?Ta�@"O:�K˛aH#�š	��mh"OZ-���Ƀ<3
eCv�I5e�Jh	#"Ovs��-0����Iؽ@�~HR"OVdX5\*
Fm	b�ѭq��y�"O�z���P0�3�ϛ-Tܙ�$"O��:u(��s����A�ɥ'�J!3�"O2��7����*8��.R+{Ҿ� U"Ox����X��5��0iX��	�'y��g���݃V� �<F���6���#vg.ov�dJ�Se�L��8�~!j�Fڣq��52F��%��l���r��ΥB ����M�����{���KҦ�,�`t&
W,�x�ȓLV��!Oe�݂���!T>m��_���C�9fy2#���7��Ąȓ%�=i���d�� �G~F���ȓp�r"M�-���� �q��Ȅ�z�� lC�4�.���޽!�l�ȓA@�sW�<A�ċ�_7<$��	]�y����N#�dߜ7u���ȓ|�L,� (C&+ֆ�R��E�XqF���E��h'�I�/�\���Ũ4����foY���I�~4�\�G͡r4,���d����*��R�y��Q�ȓT���B�
1�&��v�כ��!�ȓ^qbԀH'F��!c�䓳f1��ȓ`�]r&Á
�N����5����ȓ+��tkaɚ#�A�j���x��ȓ>�ڑ��:�T�3��݅DC�̇�1j��V��~]�B,Ѕ/�m�ȓr�2xR�JDV\���,%��Y�ȓ�^U�M^72I B����p��ȓ)�F�{բ�+�P���J��C����ȓ$�t���D�b��AgIҶn�$��ȓ|�r%)�BW�~����v�i��drm�L�!�	��地ɸU�ȓtQ�Y
 ��#��X�J0-;P�ȓ�(�1*�<��b�� -Oja�ȓQRм���){�M����#}����SDʩ�1-�$(t9q�+�
d�ȓ3�ԅ�EnU�y^��@7
�v��4�ȓL�r��C�	? ����:V���ȓX��с-�� \f�� mR�^��}��k��M�aߕtr��i�d,� �F�
h"t�˯>S��rA!��Ѕ�D,$�U$4m�8�K���"g���9Z4���C��8c4�Շ�f9��/j�q5�B�y��01e[�J	�d��l�p@��A�2-XR�@��jK����(�L�@,�z�Y�7#TZ[�-��S�? �9���9/G���b����A"O��c�O�t�2�!�#�.u�t"OL-j��z�):���\Բ`Hf"O6�eB�4�� ��Hɝ��`k�"O(�3��	�y�N5SF�]Z�xj�"O<�K�W� ���F8f���"O�ԓ��7��D@kY)+�*�"Ol��)F�Yh�X"��#Z (i�"O�%$ԓ	�s0�X!MDTYb�"O����H(H�	���Y[Ј��"O�d3 k�16�a�f�-Y:�%��"O^�%��9q�&ћu�^�k��x��"O��	 ��;@ղ�%��$���"O<��u
�>�2<�U.�&�Q$"O�����
]�"M�2`_�TR"O�ػ�L�+�:��� AZL��"O��x���>G|ض/�q�ҭ��"Ob�:���,J-�1�8���s"O���.X�� aREI�6wt)h�"O���rLN�C��ܰ�A��^2���"O�|���� 7��k� �6��S"O|�;E��J����Z:!(5q�"O*E���XRl�[ƤBwb$#4"O��ԧT3B2` ��C_�n�"O��͇%<x4 �W�f㈔��"O��9À	p��B�
�|q�"O�iy�$�;�
�y�ir� dƕ��yreL�\Ut���띘u�
3J4�y��@�Y H��g-S�B��M�y2�V!w�q��Ô"�\J"υ�yBa�)�LڔB��]6h1�FE.�y"��TѮ;��P���H�J:�yR�`��Pk��|�
.	��ybC�9�$1��O�*�A ��y��04�@xB'�<P��� �mJ=�y�F�y^|I'�NbA9�+�yR
!X5x���
�	�.U:��͈�y2 4Ke��Y�aR��.A(���y�N"́E��� 4�nݪ�y��V�
YR'��w�xx��.��yr�]�6�����NiS�i�pEF��y)]��4C�Ć�l�>T8p/�D�<ąH����U	�5d����bM}�<����a�V�ۤ,D(�0K��O�<�B�>�S��θE.4D����`�<�s�Օ*T��s��"V%k0/V�<i#�V$161��.s,��
�%Rg�<� b��5�NMifϖ)b�:"���b�<�'cXu�2���%
�0�����T�<9P�@��r�r���i���a��D�<�����<AcS��Ur�ac�k�<A7e�6�h�7(������e�<a��$q�E�s��`��e�<�w��#]:��#��.w)��ȅȓ. ]B&�R�aIf�D,RyrP�ȓ_�����f#Gn�h��M(IÚI�ȓVҀ}qW�ƀfc���oŢ����X3��H�l�1�̜KeȆ3:ǄĄ�>��u
G���3�ƹc􅊈Ir���_ � I�/W	7`�����͇�L5�	�ъ�*M�~h	$��+\l`��i@�r��\�M٦��e�C���ȓM�D�
�W�?HҢS>eV�!�ȓk ��� vM��[��8FM���S�? dc��Ŧ�被	,<)J7"O&}��n�s�H�#K�Fn�˳"O�����?>8-�
�D	 ��"O���� 3���7	ǘ)JH�"O����ᛟ]�`�s��έ7Z���"OJ��#@�
��G��1-�#�"O��K%��NEZ囧���u$<��q"O6��%�Q:��֬����ڕ"O��ס��$�"����ڧ.�}�"O	B�
����H(4}c"O�$*U�F�3�rYkcM߸.��)�"OĨ�ᜏ<U�6킌0@�ɢ�"OB$�u'�#LN��륬V6L[<��"OՂ��ޠ �lA�%L��^̼"O��r��V�MS��4hT2DJ�9�"OZ݊5�A;��k�-�6v$"""O��	���?#R��'M�W����Q"OR��S�L&J.!t*�t2�aY�"O%��ǜt-��r0d֥���"O���d�,\��5"Y!+����"O-�#��!4�0��s�/`YN8�W"O����<R<�Uk��AᜈrE"OR�n�,m�ᄐ+5� `x"Oҩ6��l10-Ą2~:���"Ox��"J�]2X�4��t�� �"O��i�9y�����޹�DM&"O>	JCKI�Q"�"�M�0x���"Ol�q0�Q�q��kB�Ȃqe�i2�"ON�Ս�8D�B�'�<z0f
"O
%�ĭ/�*�C2L��	�vmY�"Of����
e �B�iڬW���d"O�e�7��4-M���I�d���/�yb'�,0D8C�X�rPցp!��y���A��D��
J�r�� �R��yB疆Ww�jo_ w����D.�y�^4F,] '�{~����� �y� ����mI�" �b�$ɹ3��7�yr�EC�a��ݭ*m( �И�y��B�1�TD����.D�C�FA"�y�V�9��{��4�<���?�yF�xۀ��E�x5j�A�<�y,�!���S���o������y� �:L:�US5JO(jp�01�L��y�lL2� ��cX�bmi��f���y��M<M�᫄��-^j���/X��y�E͇��I�&+׻]~�٪��ڔ�yb�/! A�ƳOꈑ��m�a�<y�j.Ō�a�#l���{�M�I�<Y1	�r�$�:���~\��Ф�I�<�� ֈf�@ ���)4hㅄG�<���ג6�e�4��)��ݻ��Y@�<1ƌ�ej���H���ȇeMy�<!�oL���]S�d�1��� ���u�<q�+_�F���a�r�U��n�<ف/�X�| tI��k:�8�H�N�<�o^.9���օ^��1�#M�O�<���c��pz��E�F��5�f�<�&�
)du�#��i� h���
b�<�����@�w"�#Y<�q��]�<y��ҫ"�t���X�a�*|R�k�q�<�aA�/�T���ƕ'l��	:3�j�<�p���S�"<�#�c�	�`�f�<A�ˇ+p�R�,�����c�<Qff]�`hݘ6D�(�$l�Q�c�<� �IY3�r���u���C�`+�"O��B'o�9!�B�1\�B��"O����2>R<�8T��)~��P%"O~��0 e������o��3�"O����)��OҼ�ɇ�A�<|i�"O��fk �Qq<�!S��
�.T+#"O~pgHd��б�����$�`"OL1V�^�&�R�PuL�d����c"O����m�Ef����}~>�BT"O��*M���:���H_�3�4��"OVy!�"i)$d��I�+^ꤰ�"O�d�'�ͻ4��ѱ�H�SZ�|�c"O0�c0ʘ=�u�q�׾HG��3�"O��j�f�<�a�Fѷ0<b���"O�t#F�B=��h�e��!X<L�#"O����¡.[by�-�1lJ��D"Ol�� �8I,��"]9S �Q�"O��ذ$\�~[�:F�ܮf�"uj�"O ���Ȗ�53�d��O@Y�>mЖ"O��v��>T:�<�|	��5�yR@0V��jW�ǒ"����s���y�Mi�T�2�M=(��!�$�yR
GK���񬙈�L�ȳ��9�y� �.^k Y��zA�&��4�y�\��y��� 0�B�ka�@ �ybhp�D3cA�yvB89J���y�F?VEhI��N�o=��3���y"���FmU R��=z�j`�q� #�yB�L�]�z�rф��߀�za��yb@�N�&d B��.�B����yr�X�.f���#e�.�Q ��<�y�οz�������A� ��.�RB䉣r�,5)�j�@���ѐ��$}� B�ɵH�����X#����E��_]�C�I�)3e��I�5J�� ֌�<"�C�I�C�h,a��	�4���Bd��~C䉽�P0����N��x�7,S3>��B�	�X�ԙ���$�td�c��R-hB�	�.<����3�h���*�6B�	}�.����8QЊ8Po4��C�	'NR
���X�Y��󉍩C�C� v�)�FۖZ�`Ta�bд>oHB�	�MM�@���)�8XpPa]��C�	����d�2#Pg���C�
wB���ʂ(ؕ21e\�hy�C�X����-@0%�8�s��t�`C�I	z��C�I�^�	��T��DC�	%H���8�
�<2��}��A�&C�2F�H��&�
5�@ɡ-ξ$ C�Im>�]	P2C%2��$K�E[�B�	0st������'>D50r*��2�B��]� UA�ˁ�*ۧp����@P�<�/Λm׌M��� �-H1�x�<F/���l���؋^��{�i�s�<	@ꏛi� �Y���!>a��$�g�<�N�}�����Z��YK�(�J�<���!N�b�Z �N���"�N�<�r�J�Й�"Y�	I���� M�<��	�<́h�3vgB�z�L�<9�i �>�2��
,(�M�T��I�<ـ�L�V���I��g8�P�"f�q�<���8.��Ze�ŖK�` v�r�<�$�B4O"���Q���&l�<qr$L+-X�#6	�f�)R��Ki�<� ru@�k��������ٶXkFdȖ"O�m���%���"mH,� @�"O�xH���J��[s�M~�f���"O�X�n^9A02ub �Nsࢂ"O�)�3"&��2�mU5sN��"O�B��#\AE��W��	B"O��ⶊY�g4 ۄ+![�&|�"Oj�pC*��~��C'kۀQ�晀�"O�i	�g� �X�Xv��p1z���"O���r␀#񶅋w��+r*#�"O\�@q��>�$�+f,X�0�t"O���te�'C�Dm��kا,�n�"OJ`P�a����3*��DQs"O�}Z�ጉI),��(�g�\S�"OV��BƜ'�����j�R�R@"O�@���FR1'�	J6!%"O�Uz���7���	��M�3���C"OR��`�
���)t��ɲ��"O�m���6X\XR@g��x��"O���!iO(8�1��� �����"O�,�5*^���Ek]$�p� g"OЍ�u���
���/�,.̍(�"O�����"(�0���+g�0�Q"O�A%eۋv�.��r�@-%6(�bT"O��1��Vx����Ј>��9��"O�Uj��Ba{$m`v#�t�,�8�"O��E �@L�Y���1GB�	H�"O�!��
�O4�����&+B�Ѣ"O��Ib�X�Ab$pj�	��yf5h�"O0xG��\:HF���T"O4��eˈ s�I�$�j��[V"O��!*�c�HK�CM�[�MzR"Od@�T�ۄo�$��Ʒ8{�"O|9C��
�h�A��2Ĵp��"O���EO�g8��Cf��t��"O@��u���^�F���͑6���"�"O�1�)�<�͙0A�!��Q3�"O~����G˼,x��T�օ{�"O�yKR �R#�H���Y36C�4!�"O�t;S�O+f�񔩟((�R�[$"O�\00��M̴�q��?(":���"O"�qR��&ZnP��¥�zp�!"OPAr��C;hA%�vJ�&��b�"O 5	"��%G>�ܙ���*kώ���"O���$�\���W���K�"OfX rO�[�M����:�%.ء�y�.5.�"�0+�)�0x*5ǎ�yF��x��rҮٌ.i P�׀
��ybǚ�w,	(1�7$��б��W0�y�K�~�n�0���l�Y��@	�y��5h�����;��y���y2���l��tQg��4
�mґNF��y"�Y���4K2$W��U�;�y�Sh�j�!� �0* Đk2G��yR
/��������"����yRA�;Xxd]����;EŴ�y⤎�%U���k��jP.L�y��]Ym������!�y���˫�y҉N�1����v	�vv����\4�y�)˞^�f��_Ī��C.��y�
	.U`%J��DR�B����Ƌ�y�"R.=@�ٳF��AH�nU��y�����D]�sn��-8�Y�Q]5�y�/�"C:T�aU|�(��Q���y
� z$!d+�X�Νi �]&���c"Oj��q.�#d�����c&��Y��"O�+�J��H+�%H�h�k�"O`y�a-��@u  ��a��|���{�"O�����/�EK�m�.5�&��"OnD�KK"H�~ј���V>�H�"O>���aжkl�r�,�7 ����"Oqa�i]O����K@�~�VEB"Oȑ[��ۺK�}�K	7+��R"O�⡪Dct���D��*Q�]r�*ODE{0��G��hꖋ�"��x;�'8�P��߳G~��Qa��e�hz�'F���� �2`t�[��9g��I�'���DG��X~酅��Y��Y	�'��
cc�p��+��K�;�!��'z�x�e��S�x�T��}v���
�'�P�@s�A1hj�z�'@��x�@
�'L��2�M�D�²�оS�����'�(E��C\4$=J9�BY/G�f��'ST��$KRc�=y��!D�t-0�'�Tx)�M�Q�)(��*߀#�'�>h@��^�!���ߜ����'�d��%B�H9h���%�-���h�'E����j�:�#��{y*�p
�'��dI,S>���tTH�[
�'��h���w��r7oˢTX�}�
�'� ��@P*/�Xa��	F�8x
�'c>-���i���$���?P�|k
�'�@���lA9%s�%�$H�x��	�'e <)àց>��d����yP�a�	�'�9��$��9^5��)�+tp��:	�'�R�����w���Z0!Z/Y�$0��'��=���1ry0�0�i���`�{�'+�u��JM�_?������&�|X�'+�X#�K
�]L"\����=(pp��'����� ��� K�<^�K�'�̡���M7���{w��.b��r
�'����S�p����=�+=D�$򡠔�c�`tX���z��K@I;�OZ�	�J(��$ɐ�>-���'ʌ� �C��@RX����
u\Q�,E \�C�Is��T�Ї��0�X��7K���B��<OY�����^tpB.J�L$�C�	�	���	��ݩP�&�C&��({��C��>�Ry��O ��ԝH�)�,<2��5�I@����CJ
o�~��B�9#�.M��!D�t�6�ӦlN��x1HS	0�d��`<D�${�S3ok�X��lҨF )с�8D�D�`�O�#�����̇[̼sc-6D�(�c��h�B�dl�S��)�9D��7&
�q�J��#+������5D�ЊG!ƄW¾��ᡘ���}�W�4D��h� W5P�"p��!ɔ��$�3D�,V$Ǔw� A��R��r��PD3D����mޱm�<p`��>���IQ�2D��!�Q�s"��`p-�:Y䄠@q>D�t��H�%�,���)M�N�I����<A����]¬��7"G#{���/�;~ڮC�xy��9S�I�<	��"��jƀC�	.El�K0넪#s��c��Q{��C�	�	�t #�B?bxZX
� P>|7�C�	��l�@À1H���bON�rC�
\����cD�N�8�Ki��s0C�I�b��)��oO�	���� "�Klb�8'��D{
� �ps�jW����k��_�y]��B"O��$oW(�4�2b-BC���yE"O~�aw��B��}�Ŭ�m)�1�"O����\i$^��QJ(3��k�"Oj|)DB��<�V�A�F��"O� ��\[np`��V�[���r"O�p�5F�+g<�se%E����+��|""�\�$���(O����G͊��mF�w��v�+D��QOa�T���*^(�A ��j�C�&D�W@�I��Z�K�� ���d�>�Oe��8��ESP5XgIҟ��y��#��|��I'8��iCA!��:���" ��:B����$�K`�Qtj�I/�,��KX��!�	Y�- q,ׅWM�Ip� |h!�Dےx�jM[�h�3�TY���!�nZ�{���@���i	?D�!�Я5��8� �vm���g�0{�!��/Ӳ���m�4�����-Z�!�ʒ9niyai�2��tʥE,px!���k� ���J&䋽7s!���,\k*�`V��Gx�eI����A!�č�LlQ��ji�1�ũ�2w�!������PӪ@9KY��ksIY�!�G�3��lSEI��m?�p4(DE�!�dPhƱ�E	�c,�Xx����!��V�'vhB�!U/x�'g��[,!�D
�K�f`�	�x!"�k�@�8H!��C�x�C*�7�l��-V&e'!�$X��n�8����ULT-(�Tr�!��
�
|�d�tB������t!��BZ�h}!L�)�ա���=�!�d�O�r Ԥ�@��dh7(ݏ>�!�d[�Y1^�°���мo�!�U7rވH��� u����c��c�!�Χ)�P�"��ˈa}����,ݥ=9!�$�T"vD�ď;-b���܁a$!��͠#~f"f'�.N�����1]l!�d�`�*A��"�T�@y��JŌXM!� N��(2��h/,�ʅI�8dY!��'*�8Br��%nɄ�a#Ǘ?C!���4�2L���
B�>c׫L"F!�O�(�Q�bM^�lof�c���r)!��:a�%*��\-qh���B.I/!���r}>��%�%UV�p��^:p(!�
#5U�XE��Z8�RQAߊ<!������a3��*"�p��D!�d� N� �'��=$쑩TaӔ6�!�4O�~�Dm�
N P%����1�!�$Z��9�˄'ᶼ��+�!򤊲H�L��!iā{�|x*�I�,�!�d�P�Q��G���"�'R�f�!�Dԭ{O�	 ��Pv�&�pgǏ'�!�d�FR"h����-�⥉�-�!�D�M!�`+����AɆ%��|�!������k_6���ҸL�!��u��}R�/��B�d����7{v!򤎽4u`����d�DI�'��*�!��Tq@�U%J�S]dx�p��!�$�".4$����^2l��c �U�!�d�%o������̞Uܤ�+r�.�!�CP
6��DեT�`Ĳg�D+r�!�D	!Ap�SwN�%'깓BI�>�!�J sh"ɹ1!X-"@+3b� 2!�D�7�Nee�G�M��g�:/!�� :i����'�a��Iϖ[�e��"O��g�\J"���G�(Ny�4"O<�S�� �/��j�&H�4"O�ʖJD>&��H�e�]u~$"Oĝ���0U�ܽ#UB�j� P�$"OڅBb��$ �I�A��3��8��"O� R�[9I�x4�d�_'o����"OP%�%��K���'��|�:�u"Ol5���Ҳyظ� ����I��U�<A��){�-�RjV�U2f�M�<	�醻B)d8Z�,��uo�!���XH�<Qv�P��ᚷclq��!V}�<���N4����kKLDbD�e��c�<�Q �$�;��F�>�&!�`�<	�%B�)-:}��L��ULY
Q#[�<��g�L5D��SȎ�n���ծ�X�<)V�߹}
���(�0b0EQ�<yw��!q��'lϮN�j Q�`@h�<���ؐ�f�)�m®q��) H�d�<A��C�S4Kۿ�L57��\�<I���Y�4����}#lXVI�c�<�s�X�7��"�%B�~,��Ӵ�_g�<	��_�x�\��U�@�U��,8�\�<��P$d��M+ƻI> �c�T�<��&X�2��1��8br�D��T�<���)�fh8�fA=/vt�D�Fz�<�B �*� A��o�UO�1*�Lt�<G�0z����w�ٻ圍 ��H�<y�ץjۨ�9�aN�gqx�)�BA�<ц��G	�\� ӌ4��+W~�<����}Kp@$ߓ[@�<�A/�t�<)�S�O8�MxF�^�+�yP�e�r�<��<~I�6M�Z&�����o�<񢌑";�����ğ(vf$ņj�<�g�L�21��❄-���;Ggg�<	ě�R�A�mZ�0ж`�F._�<!�CU'ey��i�M�\�M��k�Z�<��/*��*"b�~ �}�Gn�<��gH�ZѼxE��7�(�V Ff�<��A�6 ��I3�G�=�xӆ��c�<i�)Z�d�z�����eV�q���g�<�`�	 @��@c�i��y0�J�!�^�<I4DeH����,vy�S�\S�<��"J{���e^/G���;�Ōu�<��i�0I��2���b�0ptD�z�<�b΁Y��p���,a(V�i�PM�<#b�u|B}����qj�}A(EA�<��ԫP҄\���'j�x@�4�F{�<ia/	
�9P �!n�2�(BKB�<�b�����!�f�Z�x����f�<!��B�1e8e��J�O�聀+�k�<�&���+-�%an������}�<	�W�	V�{%�0?� PG�KQ�<	A �)���"��M�`�q���L�<���J/i�IC��E�ڔ� K F�<����A���WB��8ju��@�<��¦�D��d#+WpDj�&Da�<ieեNTbp�`��b3I�е�ȓ�R��g	��~Ֆ��ByD
P��"�d�A���J���X��J�ⴄȓ}e.�V)X�PX��Z3Y��H��I�P`:�S���Gq���ǏϮ��`Y�E/B�I	hֺ���HQm���pӉХ?!�C�	%m����`���[�S���R�B�)� 4����E`z8���P�\}x�yC"OH�ytN�%=b2,��m��fB�P�"O��؂.�B���0̅>�UhD"O\L�U_�3���R��L6q�Rd�P"O���Bh�`�`�wj�#��D�"O&��EɊ�z*��񧋓�)�&"O�a+�r�~У�Ӂ+"0�"O����ʔ%�VQ�gR����D"O2����^����Ā�;��܀S"O��h���  ��M�4JJ�q��"O������=Kj.�TK�#P<l��"O.����ظjռ�:�$ܺj��5r�"O>�q�.�#zuFI��Ĝ<}��3"OܩviDw��yU��2K]��X�"O4��Smʗ2�\�Cƥ�?70r�"O�8Z�I�%��EP���DI}i�"O�Mg%Y9�x�P�X#36E��"Oe����o�T  ţ�,�#F"O 9���ַ[,��V�
vEb "O�9���;C�z��aJ�2)���"O�y�Tʍ$/{,��#	�����"Ot���O�KS@4+��ߒw謤s�"O�u#�
ˀ'4 ��k�:	�dI�"O
e���3F܀���ķu���*�"Ob9� $г
��E�!�%U�D3"O2e� Qxw�ٚ��	cJك�"Oڝ:�b
 3F8F�[�̀��"O�T��N�W T#Q�OR�傴"O��Sh�� �1$*�7id���'�ܠq���v�:C-@�X�j�aө�%6;r��m�+3�!�DK�
��i��݃4r�4�vE;�O��q�#G/~!�⯏�h�b>m1�nQ�"dD���O�n?bl�f�!D�h�V�ڵc�� XѠ9\�<ABC��o&�MF��	���ŌS$4��#}�'��!��>!�~�!��ՙ=�	Q�'��Q�+�H�:�� [36?\`�Ɗ� �D\�t�/
�%C��Ŗo��#?�G,A�3^4��f�Y�"-"��D��L#p쁭V�����>a`��`�P3l�2`�1\�8�ΐ�g���=�V�'�%XgN�V`lr�D�1-�~a�L>y�O1/�tu�A�v�(Q1��'%L��ʟ�4�u^�0ߨ�	��\�-8h,J"O�0�EDUD�A�b�0�y���]�N�h5d܅|,��!C�7~w��>�������y'��s���3�X�0y�@���xҤ�46d9�5��$�@��SL
0��@�V2^tmr1���녙QF
��q9���4(ԺE�r�r2�C�\����㉠Q����	�`EK'&��C���ےn�7qlq''�������.�|i3'�VX�Ps�%�\h�����%"������?}�	IAh�c��=o�̰6K̒W8�d����4��-q�4|0�i�6j$�`ɢ� �
{�B�I�T^��U�����`���]P�	U�T�Z�jPi�
���%�����f�pޅ�5V.^��PѢ��G��Z��%��A�Ev ���]�\�\�%��nX�APg��tr�u��]�$�Aq�Ez�,M�5\!X�cL=`��X�KZ��p<a����2;�����,o�P+SL�?����W$0d�<���`�P\p�� 	xtISF�m ���ި~o�Ms� �/l�1��o� ]�S&�߼(�s5/L=o�L[be�1e����p�C=P��� #LY�����?6��������x��ÌHk��)'+��2�aFj�*��tFZu�(͙H�$`����ÍJo��1k���6�"1��yǮL�`N�m8�'@5c�du��$,�Pxr�S�4�\�CZ��{��X�f��]"���A���4ٳŘ��I�f�v�!�jL��) ,�?`��u�'�T�A��^��y�����cK�Q�+Tpm↡r��ɣ�T�+�|x���"����'����H��R�dx6��o�.vͰ�ʙ�V.QF�T�U��)�接@���H�����I�J���;��%"�4�
vJ�`����d([��<d2�(�b�~Yq�n�T���!fb]�r��l��(�e�r5���]2��Ӈ��4M�p�9����Q8���Ͻx�`��K�g-�%������'Y��SaO����nB�'UhEbUʑ�N�69�K/��B+�td�Iץ>�����͢uy��+�N�&~�vU��hH�:��:'�ȼq�~p��I�':��<�c�L qq������p��6�PMA&"9\	�݇�	�
޼jU�Y�l�b��σ>9�� N���=�ղ`�_>����nE�<Ϊ)�C/Я���KAn[��^�����M�����cᨼ"'ʯ׉'��]YE�Ε\���!i��u�d�UG�l��@[����i��=o��2��2٦��`Z�B������'�H�5��7���H�:�p<� �\$��I�P�x��#��f�x��BȜ2���P(�;�v,(�w �8�)чxhU*�k�=��D��'���VB\-x�t�B���mW��"��l)���wO�!%$��Fe �,Ʀ���z�x�z���nQ���'v��!��,ܘ-s@���)�TӓnΒ5��g�v&�+��l8���*�5�mj�,�Q�^4���Z/Z�.H�Oۥ`�dY�)n<��>�m�+!G�y;b�U�9��A�S��KܓJ���13b��j�T�Oېz�.��\j��i�ڶ\��(��B�dU�%z�C	�*�ta���O�(/�4I��B0�3Ӄ��/��ӲL|-��;$�M�0:<ْJ�,�0Xٗ�?A8�$ks��,��oz>aӟwg
Ȕ��)�HQ�D�Y V��'�V���)`"���ꕊW�biz3�0�t�B�:�R�pM�&���,k6����U�V�f�wU��@r�ъA��K�OT*I���ɿR�:][���#<N<`� ؓ\7\ah1Z)p�L1���æc�k�**�m{u.�(Dd�Df�;#�D��@��i��2��6�(Ojt�&�:&�X�� s�x�U���o3ΰh g2<#Z��e����NS�.,��%�OKђ{T�I���6j�1+V�IP8�7E�e>>E��OL���!œyP�Q��Ҷ����*�"���3b䨪dm@$����G"Odh��č�:��aB��B�����'J�0��
��&^0P
@?��U�� Ѣ!��<y�E�4���U#�A�C7aB�d�9s¤��`�5yr�r��%��U�Ìjyb��-K5�h�鉂u.���@�B.vl!Qs�B�%u&�?A���,	��c?�iF)��H`$ࢴ-I*4!4�P3�#D�l!q߂,���c��P� �s�4?	2G^������8�n�F��1cY�p�H��w"O [RΗ.q����7b�%֨�!�"O�0���`Q֐yWAN�n+�]�"O�`�UHۏ]��q㣯�u"�{�"O<\avo�$EtE��M�An�3�"OD`�U�>��cGM M���"O�r��!f�&�X2F�W$y�"O$�ȓB�D`}��S;8��ڇ"Op]�榘�sH���AD�86�Yp�"O���(���b@U`[�J�J�"OZ* C(/Af$�� �,m����"O5� DإB} �SL�1�}��"O.X��-�|.4:���G_�`�"O��Z���J�>ub���	B�<�F"O���#����(;P�݅eP<�1"Odhٔˤ89\�)ㄗ�LnTt"O:�u.E">��M�Rm��Y���X�"O��c��E%`4飯F @q��A�"Op-9���dpU.ęN�F�Y�"Oh��lǧl��`�G�/V�p"O�x�a/$��º.�H�t"Ov�ɒJ�rX�I�Q��,I�h �"O~t���R��q�1�H�>���"Or���g�#(+�(Js��&>��r"O2qH��eg�]+& `{�"O��Q���V�Z)ffO�;0�8�"OZ�K��ˡT-\�t�CפY�"Ot��s厴;���P�X+�
I��"OXm��jgz�8Bo�V�4��"O&��5fn��Prn��k���S"O(�҂�%���0g.��[cR!�"Od���$4/IZ���m�?rB��:P"Od\���S=��j�B&;��ѱ"O�Q3!�� |8�r�ÞS�dq!"OF��W`�u�d��;
�a��"O�m�e� �b(r�<n�f��"O�H��KՋ &������Dܺ�R�"Op�(v`�{��E���Èc?:m��"O���/5�踰��/��2!"O� ��k�e�<Fw����ٻz���`g"O�����cD�L����;p���A"O`A.f���Q�̣=c҈�p"O��*���L�ҥRF�����"O(�9j	��b�pDC��8�����"O��"C	�|e>�Cv@��z�P��"O6�I0KˇO���ɝ��Ե��"O�T�0 ��S#\�ʢ�J�F���"O�!P閎s�0�0D�lܼY"O�pzoƭ�ڸ㦤��s��i�w"O�m;�K֣~C�����H��R��D"O4v��N�����L��@"Of���m6J�2DC��R�u28��w"On(`7�:��v�L-�ej�"O
!��G	3jyr��͚�H���s"O�L�p��GRT����e��Ѫ�"O����4�c2J�&��<Ж"O��ca��?G��J�U�3	F@�3"O:�ۧփ*�|$ 5gà^�6q�'"O��õ���%񬑛D�� ���(�"O�����2%�z���d˶l8�A"O�,�lNY�,I#iE�HA�"O��1��%+t��ū@��[�"O��Pk�A�^LJV�e;�2"Oށ�U#U�L�V��"-���"O�i�Ԥ�#.ר�������#�"O�� �H�^{Y���ā|�Ĕ+D"Ob�: �"H�+a���@v���`"O��砆�o�N���ǚN�ح�"O`��u��_]��aًCv�	�"O�(KF�9NZ$E0��U�Ylp��"O�1�� �z a_�Gh�$��"O.x� KJ5�>`r��%Z 8#�"O���t��7b��qˀ�Y4����"Oz�TCj���I��t{ハ�`�!���_oF�ᯋ$�n��F�2�!�>K�2i�����t�P�$��'z�!�$�b�	b\D�v�"��!�d<�K� �
�U��MD�!��
y豠�,�]溝�֭�0{!�Ėe��Sƀ�laB�K��kZ!��/0X�x��P*w�����W
z�!�ĝ%si��	Cn���>)�w"�?�!�d��x�c#��4x�&)
'��*�!�����)32OʍV�켂t _
]!�K�S�~�����؆K��9*!�D'��@��,��%2cB�fe!�Dߊ3��x�EN�`���&BKa!�$ȧ\��ݣC��b��"��؍�!�DN��Q3���UR��bOZ�.�!��̸g�v�Ȅ���r5�ӮY�Q�!�Ėc�A"di�v}��W�D.)!��[%
U�Ba۠b�jPJ[/!�d�"]�ڬ5�=�|$P6��Y"!�ā�pL]�S��u��]����:o!�d^�R��T#��:���+u���Lm!���!�j���d�X��&�=uG!���x[f:r`��{DN��Äȣy=!�EAsv��L� N&����"Y�E+!��U-��Y�*h�q�AU`!��P���4�L�u+Ό���<x!�d�z�aJ!`:7bAf�6K!�E�P����	N8�PiF��7)!�������+ڲi����!�� H%�B�+(��ˣ����'"O`���ϊ~�u��	=�-�P"O1#��E�H��h���]�:H�"O��)��:g���WJG"_�L)�"O�!:��T-k��)� _K٘p"Oȵ�g#��.�"Q�1c�x��"O��9�M �iªT��f}	� ��y� խ0��R�c��"����̈́*�y�(Ԯ�n�HT	�5�-���y�/J�@QVt���L���"��+�y	�ql���"hծM^��@׳�y�#�.lR��j�
U�������yr�V�C��́���	W�8Ā�d��y��< ����Jv}
��c!�yREH�9�\�*�љSw2��$�N�y"f�$��T2V�P�6<��a˞�y��=7����'f��s"M0�y"�+���j����JYɳE��yr���O��ѫ�Wx˒�#����y2�,P�ūPH¢zh@ec�ϱ�yr�Z"�,�!7�Z�a@t0gE��y҇��idR)���u�ؘyW��	�y2e�$@0����6<��'�9�yR*/<p(㇊T�L�6���y���ri>�cuNGVYTK6��y��R�sy�H0s쉡'��K�O��y����9`���G������y����F`��!L�k���9ǜ��y� P���A��X�`���	��y�M�#xb��B]�YJ^p�r�Q��y�ND�e�b`��ގS'���+��y2	�$LѾ�ȣ�ĳUYq�6��y�咭=Z ���@�Bm���W3�yb�@y��U�F`P>;RL�������yB�^�d����C�7���p`�F��y���7cæ0O4|j��G���y�#J����͟(����u�L��y��/?�)8����a����y�f �~�YJF��>�Ĩ��LB�y��q��H@gFY"���@
�y��Z�
'V��ġ.*�����G �y�bD�0��E(�nG*o�Hw�P��y�B5�e��	��&0�:���-�yR(ɴ/�R\1�ۆ�Z�J��ڒ�y����`�l�&`�`a爼�y"
Ъm��u��
<��ka��y�,�v�Nq��GN8�2V�6��C�ɈN��I`'@͒X���%��i�C�I�o	���2�04	�a����HC�	�r��X�w�0�흂HS�B�ɤ2I����ޮ,�H()���!-�B�I�>�t�p�#E?$��+X�se�C䉌j��1S���^v`
0
˕&�C�	|{�4��i<l Q�2ӺC�`@x�Z��D��h�¡����C�I84^1���SeH���B_̮C�I�:�\�x���<�}H%���avB�*j�z��f\�e |9c0��@m,B�I�hFH�� 'P����u炕b��C�I�>��(b'i�t���{��;�C䉀:5����
�-ꪑˡh�b��C��>QXPk���:k��b�?B�C�	�L�$e��Y$H�i�a.%��B�I� +<sB�	ZJF�ρ<\,fC�)� ��3� 1q�h8�ݍ/t�#U"O�!F̠I�l	�§Ej����"ON�90gݍi�H��&N`�8�J�"O2�I���d�ĝd�\����C"O�8k�n�4���qŎ��Xԑ�"O�Xv��t�8�3����4B�q"O0��p��qU�+4;G���"OX�0���z���Ӥ�׌�ST"O��a�(�W�H-���RVE_��yb@BN��SVMZ�[��,#�L��y,يt�4��gY�W��;T�E��y"#��A���8櫁<G���8���yBaP�+��33̅�  pz7I���yrI�O���f*�d:��'���y���?)�����x����
;�y��X��~LbA
ˑq�ؤ�aL;�y����@(��w��!~slXp��'�yBKE�
^(THs�Ǜs���9�*��y�T�b�h�Cf�;;ABQȷ�y2�3>4��
�ǒ�#�LÆ�yr�R/3G����dӎ�6-��'��yr�S�hO �#�NN�.yc���y�Ɔ	k��4Ҡ聬Z�e[eBڻ�y��R'䁱c�TqLLY)e&��y�V�	7�Шr��` � Z�IV��y����r��"&��Qh�9$b��y��PH�XfL�q��Q�n�3�y�G�[2xSCQ0"�
qҦ�y�){�N���S# �-�eK��yBe�����X�-*pl4]�E'���yB�N�*�4�qOu?� �E���y�
�o޵�2�
\m�E�$���y��=�����ܝV��8����yHR�5t|��K�K��Ræ�'�y��P>J(�2�D�M� ���n[��y��&=^���C̶Mra7�yBmG�jN- +� �T�7O3�y��֩m� 0;��ٯO�T�1����y�19ޢDz�2>T��Co�7�y��ut����7epH�m<�yR�Ƭ���9g��+�G��y���U�l|��J>ź����ybJ
�`ZNa#uG؎K@d+6#I��y����H֑"�$�tM�Z$�(b�'�pD�e��
tQ�L���[$����
�'��PjDH��豩f.S�@L��	�'ܮq�l��1DhI�Dg�<G�����'(��C��8�z5�d�Ϲ6C���
�'����ub�/NH�ƶ$���
�'�d3d��B���ː�v���	�'ь�i��7@QZ8����!I
�'}R0t��z� hbg	:H�th��'�����Q	���0-խD��(�' ��0U��% s���b�����R�'���S��FfX.�.P�"�'�0�&g/Q��`3qmڝl����'E*���Ϻ9��؃��C�H�Z�'OZT��)ת>��x���vЊ��
�'7������~��0��߲d��0
�')n�����JĂi	�i�S 6��'�0�C��~�M3��	�I\X�Z	�'�L��!MW� /PI#u�G
؅X	�'�jA�P��:?�\�D���0�^� �'>rPр�,Nj �0���#*d^����� �җ��"�d#��V����"O���a޺����� �9f
�Ĩ�"O�4��_�d����ؤk,�J�"O��C�(�v�Hh�ȓ:\;�="O�=C��E�s��k��>r��P�"Ot �f��y���j��)Q���F"O�p��ƀ28ib�@G%�  +"�#�"O �W�ʾ&��Z`�B�h� { "Oq;T�.V\[&�5�.X��"Ox�{�_c����Z�{pq"O�`��O�K�2�9�dN�K�(��"O�ʓk� VR�����(҆H�f"O�Lr��
E_�	#c�<���2B"O��*J�MVd��C�
s�|P"�"O:�`e�\�a���h+��`R"OZ-q`^'2�t$b�U�@6x���"O��j������D	W���wJ���%"O6PP���\�e�s+	�[7��"O����L��K<����ܹAض�{�"O�X��K�TC�]��i�;~�E��"O�	r'��Bq�Dx��O16S�"O��f�P3?��}m�#+{h%��"O��)�HN F�xTj!X���e"Oz娑�-w"I� ��T
g"O��Kte�S�v�Y�e���� "O�Qc���":,U&e�%���s"O���PSAN$qan�x�B8H"ORm�aʑ1z�I �ȭG�I��"O$�Bt������

?1��!"O�ൡ�0!� m;�i��a`yw"O�h��IY+@�v�8P��<��Y��"O���������Ɂx@�x�"OސK���5�(/ݒ|MάB%"Ox�SA,^��s���6��V"O�<�C+8�PD�ϒT�E("Oy�@��h$*ƁtQaV"OpU#�48��	X���*zx*L(C"O����\�c���1�(^ܮL!&"O~$��
��ꬤ��N�Q��Ua"ObI�1OH��ʵc߭|Z8�6"OB܀AI�G�<�(C�2+��zw"OxYs\ ԬI`$�=�t<��h�<qu��9�>��`�S�.|�s�i�@�<��N�k�}�Bo����Q �C{�<��n�%g�X=	d��<�!�de�r�<�Î��Zƴ:w���s�$�1a�Nn�<��K�?\MSԣgj
l1�NHV�<A2�Ͽ-9�QQ�S@XR��\P�<AQ��e����3M�g�I���[�<@�͇;S��Q��	t6��bx�<�rA�)$Θb'���Xu!���o�<	p�͵:lB%#�m>U_NA��S`�<A a�"�f�9����14N	�l@�<IV�f#���AK;���p���v�<)R�<1M~�5�����9+��z�<�C)C�+h]f Ǫ;�N@�Уn�<9���o}�iaQТ ��%i�<I��Ȱ3����B��r8�j`�<�F��b�Qӥ�ŵ�ZA��I�<��"-�Vh9��m|D���\�<�qϘ� �e�3eQ�C��m��KZ�<�ƅ p�y����>+�.��F�Q�<a��3v]v�ȓ��9FCb���AR�<)���U4�����(�$����M�<� ����ߝ�L�r��>rMʇ"O����"���q��"H�8`6"O�����׍t��1����4]_�a
�*O��V�Ι�����%$jb$9
�'��BQ(�2��')��&��J
�q�\��Dԫ��I!Wd�?h��)�tE�@o�MF{"	�hS?���^�r̀�p��E{�`�6���-�ĦOހk1e�^���=a����ӻO��]`Bmò)����'�2��i��&�4(��a�i>]�T��b�.e"1 D	G�d���5JDB"���B�xoV��?E�T�k}��	6Cـ�[a��V1B��Z_���h���`�T���0|�w�ƣF�
��G@K�ײ}HQᒽ}vn8bd�~b�,݇��+��I7	C3,<��Q���"G�Y�⠟t�2@9��S9�h bd;�s����u7�Ƈ4.��S�jV����F�ڷ9�jx@��E�f4i�h��m�y�ç0�bhDZ� j��*]�XaЁ,�DЩ�.!F�,�z���U>���1#�����I�Lwzdb��	�x��;��
L����d��h���&D�ZlHů�:x���fc?8lJč�T�8|����n7�U������ 2|V��� y���A�R��*�G��MR�`8L�Qj=���{0 A8CF�(ጙ
�ܺQ��=�Mw(�( �9CA�[6�����7A����7*��[e�<�>x��N�t��i�������g��(��@s f?
���'���+��B�= D :��%\#���8��B��03~n��q�V���А�+M�B�I C��X ��7+��d#A%
Q�B��o��[�ćaL,J��F�R5�B�	>E����B�<h���bB���C�	%/��m������dhv��0x�xC�I�|�k:z����F.J�WJ.B�ɂ-^�&cٍB��壆�@��C�ɑg��U��(M
X��	b��ؘC��8>	��BKU�L����	t6VC�Qyly��Bױ*�dboM�%YTC�	&I�Z��ۛ��L9⢋� �C�	) �����kF)$!�w�
8�B��k�V!����<�@+e�]4j7�C���J9�7�	�`���A��B�I�ur����;{�^�k$h\> "�B�I{(=Y�B�I׌u�Eښ'�fC䉃k�>L��FJ$8
Lբ��X�K�VC�	�����'��{�.��1	�P�2C䉚/�~�-� �Ѷ�ϗ%�L=�Ri/D�pA�J���6fA�,�&��G.D�¦�Y�N�h|� �̴��l���/D��R5�T�Z���jP��np8v�-D��(ƥ�4��|�B�ͦ$4(��c7D��Y��֚�4,X�\���&6D�,��a�-���&�TE���K��.D��R&��])�c�.Z��� �(D�P�B�R;:�y��I]O߼#&D�D�K�j�,!��-�3\Rp,�8D��h$�)V8Ft#J�d2���Pj*D���-�^��سNO�)Z�]9g(D�X2蚃kF�8h�`��M��b,D������ܘ���'i� ��C0D�8�c��A��U �
�&�l�R� -D�h��Ǌb8\�K��A�83RE>D��ҶfI6&ds�����غ%E>D�D����Q�B��t%	�u䢄�C�=D�d���7"v�x��:9p�$0D����c6�=E�I���h/D�<1u/��@��Tj��ɄW���HW�.D�$��K��j��FfHFA�J-D����P�W'�,ʥjZ/>dʔ *D�0x���>Xp��+�8�&��&D���6�Ë4�v	��M
�?UR�hc�.D�� = �bė`���A��ѓf�Rqٷ"OZA�ugԾ7���+���*7~�Z�"O��J��Q=dd@ "��8r�8��"O�Xc�,�Q��P�$鏹6`�i�"OjI1�E�m������&���"O�a�ӡE�'J�гf���hK�"O�h6K�4d�h����if���"O� �p��@Dޭ3�O���T;�"OlLbcN��G�pe����)O���z"O�	�'!J�J�]���
G��%;�"O�h'�5�xA31@]���m g"Oޅ�F�ѝ6T��
T�؝=�*Q2�"O��v��S F/�4��1�C"Oִ�"�t�B|{EOC�(�<E)"O&��q�XH!0����2|�
U8�"O����μc�X����.�)�C"O*���Q�_0A��M�"%Ϻ!9�"O4۷o�14��r@<R�~$ #"Ov z�Ń#HBB0���J���"O��&L�?Ƃ�����8�ʝ�A"O2�(E�{�dY��V��0��F"O�
"'�M(`c'F5�,M�"O�|r
<_y�����M�S���*D^�D{���\f�������jd
���+�R�!���,��pW�M�jS
��;�!��
t��$���s�V99!gg�!�-Q@�;��`9P�5fm!��/o&�K��)\�0��1� Ve!�$۱W��$�Q�Q�f���Yd!��)G$Y$���"�p���+._!��_h��TjˋZ.�J�oԈj]!�䗪 f�h��ͯz����B.]@!�$��Cܡ�Jր]�X�a'�8!�$�I�U�g�ܼck����Ԑb1!�$��\9��@nZ�]Y�ϙ"z!��	�HH�	Aw��;uF�X�u���}�!�N4,��`��c'�� (�'Y�!���~�a� � �y�p!�$�7 � �I���j�؁��%@Q�!��ͼ���M7 �	P�X�!�S�m��*sR@��HQ7�E3r�!�]�k�4ԓ&��!�@�A�bT�[>!�����2�X��ԩY���#X!�W'A˂���efA��U*H�!��;0v����M���q���xw!�d�jޔ0A�+z~�[&[)x8!�D×h���!�_buY��6!���0@��J�Ej�Yv�%~Q!�Q'WĜ��_F��kr�*K!�ĔY0�U[���/'g��*O!��&sc����\�,�t��&��'d!�U �Cg�C��;S`B
)`!��9�`Ŋ��Q&�B�;�oI�!���@���kӓY�f��p��9=�!���j�Db��w:���CO�l!�W��\<B�d�p�r��NR!�a)��05mX�V��X�� S��!�dA_����AH�P�Uk�@�Y�!�$��C�:��	7{z�11ņ��!�$��ҤpB��T�I��ĕ�Q�!�p�^��a�um�k�C1AR!�/I^ ���Cs�1S���	)!�$� o�|h��z�F][�BǦ/!�$G"25���g͸0�.`PR�X�Gj!�� 򝳶(T�u��ci�*n��E"O�c�$�&��4꧈I2D��Xf"O�i9ba`��Ex�gX7� �b"O�`��x�L0u!L�cİ���"O��âD�/z�ĥ�s��.H�(`!#"O�4 ��]�6�ԕ����eR�I �"O0�r'�ҭh�X�l��j=���%"O~���S1C^��
��ҿ�|��P"O��Yp�K���a���"O<mA&(,LJ�mt
�6���:"Or��O+n`��Ո��X�|��"O��{��Z�)��bƋ9"�8$h�"O�䑕F�g��a�1� ��1�"O�q�5eV�T'�t�� ���ɵ"O�9��ʥc��l�e�4�84"O�ܠ�ـ?��TbE+	���h"O�=0�_7��q�e������"O��͕#J���a�K	a&�PP"O�	���8I1�PH'�1@!�d�(��$Ek+"�(�-�8�!�dY0;���u�^	�i�$f�L�!�$�^�H�(U�XN�|U�C����!���1��g� U9����s�!�� L~$h�ę�4�Nk�(V��!�d��!֐�C��0�l�i�Ѿ!���:)�4�X�-O8C�0��QT�!�D��"����%Lx���U	W�FC䉜z��\���������S�U�C�I5w{PM�eS�u0�W� 7TB�Iu���P�+U2i�׽D�6B�Iզ�I���{��Ѓ�(�@C�� <�xc���2���SW<C䉬`�8"!�х v	�JxR�a�'Xq$ǆ$A��%ӵ`�M��5q�'�ԭi3��;_6���E�%JR,��'�
m��a�<PC��e�Z <Lʼ�
�'<���$92��!�"�8/b~)[�'���JAɮ^��y���;*�څ��'����A�˦�c�ON&���'�0DK��x� �Iҍ�I����'+�E��M�6I�1 ���9	�t��'�J]���O�_��@h�h�1Y 8�'��`��!=���G`П
��Q��'װ-�� ̲8�VI��Hn�0��'�f�"&��7a�f�AG�<a�Qr	�'	� �O��kq$r$F�GE�M��' �I�dԢ-�`#G��$��'����e�=`5"�6c@N�ŉ�'<C��9��v@@(	� Ph�'Ԓ�)��M672�����8����'�<���m��h-�e��F����'�r��P�ϒ_X��5
�
�s�'��)sf��s'DT�G%ד3~�4��'��h@"��0��c���"t�ȱ�'�T��`۾SL��a������'.ļ�G�0ⱻ�dŰ~^��S�'G:!��bD=L٬|@l$q���z�'���S)�!��,K%�!\�<,b�'�<�x�f!Aɷ*1b�@%���yHH�µJ���6%e�0JD���y����k�7e�j �s Լ�y�IJ!e�>��3��-XgFi���y"��Dm���Z�Q���ӵ�y"�T�c6H����(H�X2�
�y
� ��B��w�4R�(�$�d��"OԜ �*�>@[���)t $ �"O0�!d-��O,J��iA�,��a("O���a�vt����0f�p�Q"O�=h���[gVQ����L�21�4"O��x��۱Ef )��͐(#ƀIu"O���U����Kwl��K��,��"O@�K�n��Q)�L��+��c�|��"OF��Bd̞m3ЭЕkJ��85�'"O��[ta�t�̸`��B`�W"Oh�#�I�1J�<���,�l��"O����3N�pc���(m>$å"O�d��'���#n��X#C@�z!�d�-���
����J�w�!򤝺��ě��¯:r��I�oܢr_!򄉔c� ��J�O��q�5o��&!�4;X��%bϡ lDp���H�J�!�dQ1R�n�2NP�[Xൌ�D�!�dR+��q $�H�����W�T�!�Ds,��@�Բ9��)qQ��W���L�7U�xġ �B�\�8v�M��y�D�	�̈W/�;0�<X�eR��y��4a��4��i8$�n�Zq��yN-B��D`���9��"���yr�#��e]0~�Mi��(�y�I�K6�뷈�.M ��p�Ĳ�yB 
��x�Uǐ ���B�OQ�y2���/��A���ϋu������!�yR�0|�ޕc��O'@b��{'=�y��˰8KE�F5�ة�gù4� ��ȓ:�J!N'��dQ��Wƞ؆ȓn�1т
ȟP� !��PZ]�ȓx�l����]��h:�ْc��i��'��h���$j:j<:$l�ivT�ȓ��� @�?�     +  �"  �-  ?8  %C  �N  �Z  af  tn  �t  �}  U�  ��  D�  ��  �  <�  |�  й  *�  n�  ��  ��  2�  u�  ��  ��  9�  ��  ��   c � o >  & D, �2 �8 r? �F �N U D[ �a �h �n Bu �} 1�  `� u�	����Zv)A�'ld\�0�Kz+
�D�/j�2T���#Ĵ���+�?YV̒'�?��]O+��yk��P)�T�pH(�����8��)L/	����'�� m�E�e���S7X����1"���r��=�ʝ�A;E��8��/ xS�'S��pH N؜3��<���:`��:�f�ǰ����(4lc��˻Wn�1���X3_�����i��A���,D�r0o��a��9�I����	ݟ���/|�^Adpv$����\Ӑ<��>�e��h޽�Ms���?Y�� �F�����	�1IR��t��-��聂0K�����O<���O����O���Rk�N�}�,u�BLҔ7�Rh�#��pɠ����xL Г7ͥ>YN��7m%�,�F�SB5sO���B�|���a"�+���~��&���!j�)[��� T�瓏.Y��X�O� A�Ձ�*^`�$�O���O��$�O��d�O�˧�y7+��6���Ŭ�j���♂�?�s�i��7M��QQ�4�?���iF�	Dx��|1�@B p��x1*Fyn*u(�&�=rH eHUJ�F}��bӔ(�p��OVip!
�yoTq �fɽrI��sYw(��!Օo�d��a�ϧ-�N��
vh���KV�I���&)��-bӮ��?��SԺ���%&k|	J��<�c��>* il�&>f�HR�Ł'����K���c�ʗ$c@�q�4tV�Gc�d���E�A�PU�1c�H�� �EQ4��С���o��MC��i"�����d׈�[�g��g�r����۽L�C�,Q$
�ه�ő\	���$O1t��@2�pӠ�lZ��MS7fL�C�29Qh�= ,8���mE�/�6;Oq�⟾ ��-P�<tH��ؙQ��.�<0�o��F�%�;���'S�&��H&, Q���|�����'�O|�D�O@���Ŧi�	��D���є<�A�<@v4�oD�X�ɺn~N��	��	�7�F�!ط64���O�0�MS� M�D�♁e��t�U��@�/Qi��O�'�(OH��͆
ȠX�����k�6-���6cT#��)[d"ē0��mZ!���<Q᫋}y���<�d�&��
a$�-'l�!�,�ܟd�I�D&���	럴�'|�"�"��9��#kʜ�A'N�^��'�|Kq��cr�'�t�s��)��|ҵ�ӐI���7e�K����a��O"�I$Њ��i���	t�mC"��O�����һjά\3�
�O��N˂M~���e\	]$����4��O�F�Q�-�'*��$�D_b� �@��`���؄�@Ӈ��R�E��`��$�� ��G�
]�­����2{���{�ΔE�d0�*E�7��$( (��E莘��|��'�B�'X?E��*�� ~��d�0-:�y`0�;����r��b>�i�-`4�!��ʧc���[ᬎহ��ɟ��Ɇ.�=(E��˟<��͟,��ڼ�qk�}Xx��O���!s�y��'S��au�'`������I@����~�hQ�!�|�,���b|�0�I�I�69�1�1O�)��/X�>S�5q4��pXBB�V �'�]H��ϟ�'���A�捁t�|MS4�P+�㘝8r�)�5�\��i]o7���_;&��{.OB�l���M3J>ͧ��.O�,"�/�l��=}a����(�"w��T�'��' �	[�4��
A�cH�(d���h(02�1~)1�G؂f��!�m*<O���Ȕk���nˆ\V�({r� 3|J����QZ�|�6�/�@�����D%CD aX�hu+E(�����Opnځ�HO:�ب�/�	V�]��h��V1h�ӟ��IƟ$���Y��yx��W����AӦY	B��Od�m��M�.OJ`@���ۦy��ܟ�����)T�	6��?.Ve)�kӟx��9Rg2��	՟���;B"ߔ/l��(�̇�;�z9�r`R����a���V���r��CF�x� �1�E$0L� 3�J9<�ĕQ��*ۮ|ZrퟸTZ-���P�!.�Q�!+~��!.0�$���H�4�?Ydeχ	0��f�A�E8����ۘ��y���	e���>������$X����m<���U�2<O&���<�4�i1�����
 �N�#Q�_*u�T@��gz�h����I�j2�,b�i]Iy�O�T6-�HX��Kb:`�s�+D�W��b�d�O|�$T�PɈ܊@ �4%X����RV�=J���Ô�,B �*�a�F
��HU�9K�	-y���؂l�Ds�C̿i�L�תO/ϊ�����?mE�P�h/r�H&�)>�|1:RD3?q�Lݟ�{�4��O�1�⁒�AP���1��ݧ$������|��'��'���'��I'#P ��^y����% ��q��ҟ�m�����4�?9�ϒ1P�|��k�0w� Ճ�Q>g����'
��'���E�μe���'���'���]x����PCH�u�*(�d�S$w6���,�84J6۔_�T��B¢|�!�$>F��L"�����Z�X�
ub�Ĺk0Db�+�v�,�v�)ư���V�J��҉DC@9��+����o��]����'�B�'��$bĨop�I��[���֝|��)�E�@9��D����	 e�ʓ���nӶ�O��)�0˓׬����N�.Z�m� ��7��݊��.|����'��'��IT��6�D���S=q̠�l�V���u���:�rtFB�J�T	&�"<O�!c' ޕ�!�R	j�|�pK�7��Fֻ	��0EO�1���"��!:C��&��.L����aꝠ
N�ы��OH�n�'�HO#<U睤=mVA��6L�����̟&���	ȟXF{"�L�?�h���@.��Q#� ̨&�"v��ė��%"�4��O�;X�o���@�T$ A
]<�Ȱ�c��N�(Q�	Fy��'sR;��43$ ^u��/|��7!� ʔ1�kV��r��aS���'z��AnՎ3�,����]�w ��F�wC���#H��L5r�;	�a����<w�x�40�'���P��ɶ&���M� �b��I>y��4�ɱw܌	0@+�k�F@`�	� ��	�M�3\yL���ae BR~TY� @�Wh��V�P�c�G�Mc���?1(��� j�O��ˡLF�䬱B'�B�m�J�Z�o�O���X;H��VK֒f+zٛTE ,e"�Jfh,����O�j\���˘n+�q�W��=c ���O�l�È�AG�D�P��xT�0�!�M��~Z��<t"�H
1��=(h�a�j4}2B�9�?�&�i�.6��O<#|¡Ʉ=�ŰR��*)�({2��ǟ\�'��^��ߘ'���"%E�Q+�}���&<̺��Ó�Mr�i�{���H�&xDrBD�|nha��v��nZ̟p�'��	%�O0��'��^����H
aG��6bʱ#�ni8�cЈn0-��n��
���m�(��	Mw�Ae��	�I�ip䌘�� nj!Z�`�W:���UA
rD�I����v�'H%*��'͖	[��[/po>!��{E�3䌄�m�.O\p���'��$�?�O�$�Y� ۰$R㯖�oG�<�C�O���<)���Ow�ɩ< �����Ge4�I�L(��ᛦk���]�}�O���_>����S� �d�XRN���@[l��L�֬���������?=��ȟ�ͧO�T,P��I1�<{@�K&f�f��\�!�8�0�B��A��*z�l�F(�
YoQ���6@�;{�F`�@L�q}he�W��(ؤ��������xDA��{�,��˄;M�Q���dM� @r��B��I>�x��3�O}X��Jh���x!�Q�.�F�R�,T�
�����j5LOj�$�rf��ep\����m��ɹP�8�$���'�d�%A������� �6�_U1|�ɥmӔ~:r��4��R�'�
����'�"�'�Aa���k&0���,ާE zeX4gS-i�\�ۅ���NJ���1�	V�m���H��(O���C�^>v � �ܐ4V���M���ꝈSgO�4'±�&"��l�9����(O<%���'��7�[����	"s�)V�#9/����T!-8E�'s2���#�\P�����n�Tڃ�N)�8��d���	�#T�8����>�r9��c���M�+O=B�ϙ䦍�	ϟ�O�je1&�'0����>^(�1�&ٯ6�̐kQ�'��cT�}�EkB �5@�X�jP�dN(��W���Sk%� ���P�}#Rя^�n�^|��b�%�D]��KH]|x�k�%$[+6�O��@�4J�:)aL���,A��@s�OȔ��'j67m�l�O��i���iP��C�c�t��'M�@S1�Oe��X��kO,R�H����*�Na�fIl�nc>�@.�:s�pJ P!mrD1���������X�	; K:�s'�蟬�	�����Ѽ;�㌺G� IB4��2A'�j@��*I<�,��M;
	�IdH�x��T�i�,�'���*uGY
L�e!H2\��\zюR3`�b�i�j�(��ݗO1��6�[!��$߾=����J�9>�F(:�lEB�ԓOH8:��'�1�1O~�P�T�D��r���dv�J�"OНJ�jT-�@��C�ip1���'�2�;��|*K>��ʜ�G}�`3'�H�7z��!QON�g(8mh� @��?���?���H|��O��$n>��w��T�@ȊwU�_/XA�u.�>Y�"�1�	�h�U���\o� P����D*~+��`��g<����B�1r��f�q>� �"A^�N�����J�ir�ma��D�F8n��2�F3#Z��#Kׄ&S"}K`�'J����	7aj��䠗��h�ȑ���2!��[�O)��7�Gkyr@�V�)?�'��7�4���2~��OR��wJ$�G�^�a�yZ�g�<R��'�����'r"3��at�l��ЁH'b��ؤ��M�!9G��	�5������t�?9��Ҧedf@ ��ȥ}
 ���l��pB0/��U��@iu���SHD����� ���'&��&$�
�۰���bǈ4|�h�Is�|��'�az�CVkĤP�D�J��N� ��?�S�'�$8�Q��!>�@)qҠ =)�����@�W��l���8��A��a���RÕʂ=2��Ǉ2�SD�i���'-��\&%/8��Tj 4�N�3�D�~ʟ�|x�bI6{�X�œ�Z&��W��h���<)��h0S+N�8��� eo_Y��kOD��g��1Q`��ᰄJD��'������?�����Oj���D��Y�&��wrf��
 D������h������-Q�dRC�:��/�>���'^���*��0H�bަ�����4�	�$H(��b/��H�I�������'��$e֭���]�NJ�P9 �3X��(�`Y�+69Pդ�7 �\'?�y6�ƌo2��7% 	�w�	�`� ��%\
�Qf�-N T�
Q!�/u�t�@�4�654����ORU���I b1�3�م���DFu�@5�'�(\���"ϟ�'�+bK-~,H�e�"�E;P�Mfx�,�b��#!]�˲��\²�I���ɦM8ߴ���|:�����_]��� ��4gLQ��C�q_�+Î�?=|�d�OT���O�����?	���tJW���p1*A֐�2j�'s�v9�Ӌ�� �R�ȣ���Ƅ�{d�;�}KĔ� N�jp���o�pmiR��5Ꞩ�$�I�!�����ڍ6Ͱ�;0(D�JNk������=b�(ݓ2���q�x��hI��'�����R+= Hr���4-�:��mh�!��'G����Iׯ+fH����p��'��77���(lC:i�O�R@5Z8���.�6�� �R���'�Ny+`�'��=�9@����X�r��B����E˃z�
Ń���:!jLx���<oh�E~R�)z�
�Q3eFd�e9%A�O������a��9b�1� #���a��Gy"j�9�?������M<!�D�D� �+֣
�(D�'�a|�nX�`|t�%&
�7�4��A��6��?�!�'�@�j�0���W���<Q���$R;4~l��@�	H�TɈ8!��Z�t@��E���O��"�'��EJ�'�*['I�4r��k��W�drn� &0��IS��?us���P%�T� b�L�U�b)?)DǊ�Kg؀�s匏XB�)���Xu�|�dF$�d�(VDzS�� H�����I���D΁A'�s��F��2�d��l����#'��6�Ba��"O0��fZ�g��$��-
)=�Yq���%�h�b`3�ű\b�T�ƫJ*'�ʴf���d�O@�$P71��İ��O@���O"��~�E�Ǆ�T��BJ����ݣ��ӭk�fgN¦����ܿ{�B��|���"O����0$�t(�bL"W$�ӫ!y�ʑB#lK�*KƔsr%N�:�2zwI�)��'F��i(��3�I��J�f!�0�\�j��Tʂ�M3dX�(H3L�O�� &�8`U��6�2E���U=P���Y�<�3��x�)�(S ���p�̒`yRI'��|���d�>����ۈ7�P����Jq��a�X�sE����O��d�O���;�?�����t J�\
5�Y-f�*M��i&o |
�Gݚ>cZQ5oM���(D��Dere8RA�d
�G��(97 S4�qb�'M�x�V�>~��p�݋Pՙ� �;�?�Էi��6-'��)��O�����Z/d@&���zs��ӓ��'��1[s���h0
ӃL�x��AK>�ľi�RP��ٲ��$�M���?��ήV���F����x�<�I����͟P���|r^}�I#��\�� }*��g�Z@��k�]08,�#M�]��0�a�Mɔࠎ��\T8��ҋ�y����䅏w�6x����p�V�P׮G
]�吇�<_�x�z��dG�G�r�䇾�V�I�'��>�xujs`�;2�!��Mk�Ju��ʪ0�� ����6����O���]f�@U��l�d1�xI�|���t?�6��O��Ŀ|�eo�?ar.�4�1�M�]D�ݣ@m��?A��:�FfU��<����@T?�O�S�%$0��#��bW`��b.��{��h�pl�P$o���Sb(�'Gو"5*�?/��0PS+�%8DZy�'Yd���?s�f�1�'�2TƼZn��F틕t���ѓě�y�� r��c��n;p�hSf�,�O��_���)U�Ny"��ԩB�^#���A�M���?1�}k��R��?)���?Q��g)�j��ٚ����ge*�`�Bؔ�H���Qt?9����j�|�<!�U��d��Y[��K�+�75�R���ģ��Qh_�c>c�4�! ֯ ����h�
�qE͜�e�-O�L5�'���O�Ob�q鈪�>	2�+ӛ&~�-{�F!D���sOC$($��+s�\�0Ҳ�V-TO}�"�/ěv�'������ �6��C@
|�9"4�M�U%�Y����(��矤�Xw�2�'j�����Hf�Y's�Tz2�Q�hLH4��W�
�;j�:�p=)4 X;)Y���3s�x��E(_�_�đ���=N\*�zj+\O�i��-m�Eڱ@�6{�x��@CſV2RH~��%l�n��q	񟖘�rL#�%k�囡��G�f���2�ɋ<�(���B�a�$(�a�?+%X�O�ml���'���4��~���X$ $��Jk��pG�]g:����?���
�?����j�=��0ƪ^m�m�'��z��8�v%�sJ��3Vꔅ�I�+�!x�-asD9�!�O�@P�h�� �j�����X��	#d�'�2!��3웦�<	3�.u�5��$R��h�"�U�I۟��	�,��M�%́cJr�Zv��Q*�c��F{*�����!��0����� 5��D_a���$�<�nk�&�'^�_>yq`J���顇[5Y��mh��P%*7�T1p�[����� ��ɣS 9pE�SaU��M[(��ʧZ�����t'�ų4��o��`�O�L���Be 4����O�� C�
I�x�1�H2m�-z��� s��=	p� Y7��,9A�O0mZ��M���� ���	���ޕwCReKa�|"�'q�'�� �P��3s�Ҡ1�C�B���(�z0��x�<�O�u�#:2�� �N�J���G 1��$�O`��ӜDh�(ã�O6��O�����Ǘ<5. Ba�����Va���y�'���C��8k�ϸ'�*D� .,�� L�ڱ��L�(>����v�Typ�� %S1�1O� �`Yub�	$.RL�B��RX��m�rx�'��x�����ɟ�''� O�,��6m�:9z��Q�q�4�w��iBv]@@���bԦ,c3ɶ<!"�i.6�*�4���i�<���8B�����z�ir�`U4%<m`w�X+�?a��?�� x�n�O��t>Q��&�<v#`��?���I#���x�� �
)$�$X�W蜈�
I';.Q�4ˠ��/:��`4�� y:T�)��!˖�c��VQ�9��I ��pa��48la�?���$"!�\��#$y��6	T^�������E{�)iYM�gNT������5�<B䉽)$J� �W3޴�1���?SjT�OJ(n�˟�'�n�WC�~��u����EK�;�V4��Ή ��!����?��	��?����ԠF5y�B�+���:�j����i�0�	c��iq:l��)CSV0)t�΃0H�Q��Dվd���O!g6��`�b�B�����q�n��c��U�(�'
}�k�@�c��]�IꟌ�'w,�6�E	񄡰4C�#J�}iO>��w'�E�?�r$�R��dq�ȅ�I��?�@���q$!��'�b?��Ku��֟(�'N`8h�.}Ӵ��O��'oĲ)S�a?fġ���L�쑖-���d�����I""$����N�/��L:r��!��%"�@�)Xp�O���'�U�2�!Qb�S���OZ����I F�.7�W�L$�XCU�;�0�$�Tg�tBI8p �Q���Z3h`����2�'՚��I�M�D�S�|Z�	W)�H�[��ց:���!biXE�<��I��\�V8�NB)DKx��	y�'팢}:7��cA�@th\��ib�l��M���?)��4e왠Ȝ,�?���?����y�A-^��bg΋f; �H�튫2XZ�KcBU�XiA��bڔ�S��䇟�X�J8��BD�̳��X&Y�K�nA�4��]G��%\D��f�v�k'�P�L��c>�$& {��ē�t�,��N�0sFC�S�7�Cay����?!�'���|B��4y�څra�H�L2�<�L�Q+!�A�
��K�0T,���#g��(O�Dz�O-�V��[��/�QQ�$�
��!�7 ;���Z!�[՟X�	۟@����u��'�0�b�~9	��ڦq��"dL�;��ayc� '��u���W�'�	��V���Ey�ŗ �s�U�
������Sf� �R���`��s�Ĉp�
ŋ6�F�0Gy��3b_����֨(H�����u8��q8�b�F�Iv<E�-�>Wۄ�2�"���y���	$�t�R��7E��@r�`ߕ��:���|�Η.{z�ꧥ?���0
.�0T�8��Q��&\��?!�Q�	��?i�Ok�q�旙��A��W�� N��w�H�S�jӂ8� �3��=��I��h�b�'�N��,�
g�0��C[��`�شBK�B����E3�钲ѦDh�H��EQ�',\��w���<��G�*
bA2���.E��ɓ@��S���`IǥM �D탨qc4��f;�OHl�	�d�F� �u|.$c$QTCH�Į<���FR�&�'a�X>�f�	ꟸ���sSHI�cN̼V8ZUb��D���	 �L�g%Y�*X#C�֦ACQ?Q�Oa�)����Hi��)\D0z�OH1�Q-٣6�dj¦>>���T��Y�i��h"V4<�&m���G-R��	�ix@�$Ʀ��M|*���*�O ع�D�q-��h@Ė�5A6xKN>����0=���R`'z��@m	�TB�����s�'�b�>	��4�̗���3�-A�9'�apƈ��YR�F�'�B�'��d�6k�)	��'��'��n��7�tz`HݮbTqA`KZ�S�j��a�ɺ�
%�u��=�|;��)?���3� h����%`G |�El]���ؐ��=>.�e��e�% �i*��O*X�4h�Y~.���f�!5�r������O��D�O��<�&l�g��l�&)�I�t`�F�N�<�2D&x�v�� �R�Vv��F�HyR<��|�����8��@IULR�V+xX�C�A���wZ�c�>���Ox���O�E���?Q�����S�]��-Y�mْ 92�1��J�TT��N�"��}p��^+&N�C��ɯtV��`�:P (h��B;S�| fA�7/�04�M�q���s�\�'ؼ�2��>5D�����6��T��.��?��?	�R�ӝlٸzu��)}l�@儆{��C�I+5�|��j�)>\fԩ�(N羓O�)nޟ�'κ�Q�l�~��;8�!��/���-�B�<D���?�Rb@,�?A����G�I�D�q+�s���14����@�GမC��D�"`��E7��-u�9b��Ժ=2c�ӂjw��:n   
�A��M�@�V 0�ӌ��O�$��'-����o�-2{����e� 8�xY���&���Ov��2#U�4C�H�
r�0D�ʖF��k�O8lQ�eS<�x��Ɏ�c�Q��'�	�F�"UR�4�?������:�b��J5�&�)T�#>Y���45Z�d�O@\@�:A�R�B��F8�*J�T�?q�t*�4��ģ�О���r�H(?u�׺q��[�5�e�ᜇ��O��(�둘��!�S���i'��h�O��C��'R�Ɵ�� T4��lM�|��r &�cǢ��"O��B�NX�B��@�ݥL�B�2�	��h����De�,+5ڙo�+M�(��}Ӽ���O���Q�L������O���O:��{ޑ��Ț6��h6-ܳ"<A��9�fu(�K�R����&b�c>!&�D;�$��H��`��Y0'h�b�cS!Q'xD��n�b9��A@̬A[vc>&�@ʂDPb�PR�K�bӜ�ه�`�I`Ӑ��:�3�I�2Ӣ�a��ˆ(қA��C�!;L9���)Y�|�B5cZ<�˓X����O�I�1HR�+#�.+l`�H3F�v�]� "ܳ;-*���˟\���#[w�2�'��iJG��`0eN�4ym�-�ѣ�%j>|	Z�k�`�Dؚ P�p=Ɂ�U+uҾyBf�?Rƞ��P���)S�+���Mj�
5\O����&F�UA�d�0{~�9�a�%$��|�p�m_�Px����7��B�t�s�g�?o�"�he�';�O<4���+d�1�v���tȜ �|��z�����<���A8Z����?�@g�ӳ_�Z%���#S� ݨ�o=OA[��	��J����2{�l�JL#zk|���?n���r�@C{���#Ah��~����H2O<��f�'�1Ot"��L(y��)R%0�J��"O��ܷX���H0ElR�v�'���d��]XIh����>v`he��-n��'�F��e�'U���O��'�����:HF]��AX~К�j$��?���NZU��k%&"0 �M�=/��� rx�\0Z`� ����	-Wjf|1Bh6J���ŉW�O]�����/%j��]�Eیq!�OD�2�'�b���<���|�V��J�������X�<�$���!�����I�F�vL�Ō]T�'!��}V�ј&����	Y���˦��ȟp��`�hy���!q22�O�R�',�ɘ�T���K�6�K��c �,	�J̙+��h���l_�DC�I�g̓g�r���MG *�S�e�pP KE-^M�����7�ub��i�g�ٜ������~m�<:T�ie����e~�2�?����hOH5�5N˚��Q��1pc8e���1D�ܠ�m�>a��(s R}t���<YT�)-O`�!��>8��q�X���	��yӦ ���O��ҧ�C��v�L��4AEh*�ǿs�'�m[B�9A�5<H 	��Ģ�?q���?A��?٢�u�X�"�$�� �D��>�Р���x�̨��+�<�`��p-ގ"�@Gy2�)L�(��-@� Ҹ0`"k�����*TbʜdѬ� b���9`/�"LxtDy��G�?�@�ioғ�����C�Rl�h��|�J��R���	���p�U�6*$��p�Z�/��$�xy��@�;�z�`UJ��l>�ɻ�KD����N�4��$őnF$�Ħ|j�G�?����檀S��L�~����B\m��1��Ԡ�΃��My5H�z�~Tb��D�>0������e[�	s֨�Z���1��X=�y����S��Q�&���)�TU���ǃ^>��EN�V�'R[��yOT�J_�Q�A���0(H��$�DQ�	��M3V���R�'	�nP�`
��`�Zf�M�.`��2!�#�_�E���VO��KAD{�n3�{r�3��մ+Qʭ�r,J�F�80�ֈA�?��^T5��O������?i��N��.�Oh�&�ږ(�bYarÛ�*��`�
*V`Հ�	[�&C�!��k6b�'#��
��:}B�W(o�
i���BӀ$H�!фR~�]�e��;|�(�Q-�#xRΟ��)p�����I�x���%%�$L���R��7<��J���Iӟ�F{�:O�){��'������-.2M��"O�h5F3{���
�F&�I���'�:#=�'�?�)O��X�.�!8���Ƣ��b��VVb�b�8���O ���к��?y�OX����K �Ʊ���rip�)�h�x���ۣl�
p�1A����r�"?�ע��R�<����e���h���<E���b��\��|:�IKb.�#L�	��<��O����!(��Q��%��	$��O��=����X���:Ђ��8O�)���;h�!��Ƭ0Z��D�ԕ`�����˼]~�Ɇ�M[���K�U���Bk��$i>%�B���^�Ɛ;���^S\ͻ�B�O`���Ot���O�d�.K�[�:�[�h:@Q�����������JZ~`�PƖ>R$�{c)K�}EQ�$��}z����b�&3;�dz3��J$�c�V�.2�M �sͤ�"��C�Q�Q�X���O���3���a�Tː3I;*)�ve�@ʓ�0?ɥ��){M�Y���'lĬ�N�fx��
+O�L�C��^7Č 
�:)�!Q�^�p`���\Cq�V�L�O�	�S�O�B��PJ�E	.�:p:�p�_7a����j��X��a߸(B<�Z+	j,:� V	˵q1�p����)	��#ֈH�tH�y$7O�$�#r�D4��s����2},4R��t��\@@��Qn�5C���QQk���yrdD<�?���������� ���D���"�"��&~�K#"OZ=����8��PI�Ҡ�r�	"�ȟxu�c'�`2�9�[`"(�����F�v���Ox�U՜���O����O�I�O!�sg֐r-��"�Ǹ}���6�N:
��(�� '@�����|"�6.�PaTi>}��0l��*��=,�6ẰL7_!���˽)Zb�+�M�=<��P�Ο~|�V=��IN�@$K`�_�0͢�.�" ���������G{�?O�!r���S�����q��-	�"O��w��o#�m�G($soQ�V�'��#=�'�?�,O�D�������KB��0<��0��= >� ;2[+��D�O��D��x���O���JMj�J�,��}���=����Bk�"�q�s�K�eУ��ծ���I�8XͰp	��1F���Z�
��r$X}������'rr�������6�?n���ǉu��	�Ȼ?,���� `��?���O�l�L^2A0�ass/�4X��d��"O:p8��^�FM��A�^��P�P����4�?�.O�U�!�Mצ��	���'	��f��q�J�w�)j�$�	?Wr���	��I�*aa��l��|B�%��Q�8���$̃g�h��m�z�'�f�R��I�I�0��=�4��N^�|��4��O����h�yF��蓛Y
�`+�[[�<a������P�D�|�huoZUx�0�*O����k�d *�(��R����џ��ISyV>��O��
��Tz��G�>�jͪ�O�П�'��S�'d*���%� =�(���C1d��?�ش�ēh�d����F�2An��'� a�`����٦}�	��MϓW\`�	������͓1@ҀQ6��V��؉�o�s�aP�N!�M���Q�����y"
�������7џV�]�[N�!�p�˾i@ �p!��mģe�'B���?�$`�%�I��(�S��xyt��"�%P��7*D�& � ���?Y��}�L�P���2�������/?�ش|p�]Yw쉅3��b�
�$:Z�dtb�'��Q��Š~���?!���?��,_Jq��F<M�,u*�% 7N����'�?��`X���XR�����ܴN��y����ҹ�$C
M6�B�"�,O���A�O�LP�'�	\��$hݽ���P��E�4����5�
	CH�8���@��^�<iQ�������u��'��D�!���is�j�(f�Y�6� l�S$ȓ;7���B��dw���b�4�sC�OP��Y0��Sğ��I�8g��N��2 ���=r��4g��e"�'8�̰4�i�6m�V��HΟp�����?Ur��Y�'����U+�T�A��V٦-� 4�MS�P�ț�'�M���O�韜�,H�P�s�#K�B��h�q@�X�<٥��1	pP�W8Wv��E�증���x�������ߟ`���X��˟����<qR<g����L�-o 6��O����O��$�<���?Q��?�ֆH� ܞt�5��@��zf��x��V�'��'���'��'���6kJ�mPW뛀7�Ő�)K��6�'���'�r)�~r-�f�'7���F̈�~0E,��3�̱�O����<������2� ʐU��!��ЈO}\�3%�3��O����OR���O�ʓ����>%����)Y�>>�%s`�
��$�O��d�<����5�T��u� ���gq����׊�y�ϘxI�Y�!��/3��l+�Ε��y��O讍�qO�~~pU����l�<�#F�u��!��Ȇ{S,Y�0�w�<Iw/˶e8�: ��?)���"e%q�<��@�-�P���	D8cK�=��,�o�'��'#b�'2�ϻd�  �EтO�Ѝ����Ab7��O^��OB�D�O����O��D�O��$2L"�`#F�1N&��v�q� =m��P�������՟\��ן(���������|J���-u0��S~�rU3ڴ�?����?���?���?I���?��{I�9��5{�rD	�qڄ���i(��'"�'2r�'82�'���')�Y����Od�eK�� 
�"�(c�@���O��d�OD���O��$�O���O��F杼Wyؔ����w�(��6���u��؟��I۟��I����	�������nFfp��T*p�5�� W��M���?q���?I��?9��?I��?y�o��m�Y�]���ٕ$��m��T��ǟ���֟��I�P��˟�ɏB������*P?��b��%�4E޴�?y��?����?����?a��?���09����".����*�_<: �i���''��'��'k��'��'76����Y�Ar���d*�A�$�pӶ���O����O����O,�D�O��$�O`utH��Q� ��m�* ��8�Ԧ��	��@�I͟p�I��0�I˟8�I���mf�d�C��G!��`g��	m�`~��'��Is�O>I�dX,\�Z��t+-Z}�\R��i��I��yR�IW����w�T���JQ50�$ ��B/Mu��x���M�'��)�)�H��a���O�$�)��sBM,���zS�'��`��0#����i>̓"�$̋���<S�4�+JG ���|y��|¬oӆ�"��d>� .�a�@E9p��[S�L[ژ��3��ry��'
�?O�˓+$p�jf ��n2݈���_mL��'��U��R�34ry��O��Q2`�j��t�|Y���7t��u�s�5^�@l�2I�<y/OB�d&�g?�g�V<z:(�lK��Xl@�`�ǟ8��4]�d�'�6�9�i>=+�C�6��'+ʎyn� ��0O���fӂ�$S+2Vڜ����h���ގ'� Ѱ�=�BKÖ� D�Q3 W4��C�I��Ԗ'1�&hYc��z�c�7MI$�4Q�d��4[��`�<1���×'?�n�j�N�7_z�����{�tʓ�?�ڴ�y�铞R����$+Q:md*���A�F��<�1A.N�n�9���"��1^�d�@��$��l��8��,I�$ ,�r\����D�<)(O��Ovo�f�n���*�L��"��v��6-Ą<���ɦ��?�g?!��M��'��I��_$��\@��L.�~E�nL%-��̓t/�䊐�Ś��
�����S�����J�3�e��l�o]��{� ݝ�?1���Ľ<E�tU���E�x����<����F. 9�������<��m
/U����K� VY���VG�<A-OZ7�X��	���0��e��q�֝a��%��.�
#J�D�v{�ȱ%.�5�n�	r"�1Ae�'j�i>�'��\2e(LX�1���$z�⒬_�`m��|r/vӺ�ۂ�9���&p!��Dܶ%�#�|y"��<���M��'��O���n+4��̐�j���fGT�ߠ���H�)^� X�'�
� ^wްQ�n!k�O�a��OP��t���5]׫��5��	ǟ\�'������̦���/�^7j�h��0Uu��<mF�f.���4��$�O�hbq�μx7��.&��(�r�7�MC��C��L�����<���D~��ҳ�̰_H��'���KWꜘ(�0v�U�3n�Cu�'���'�B�'�2�'_�'w�ӻ`:�8��8M�h)B��C> )ލnZ?��\�P���,�	�?q�����O��̭^�Lm ���-dC�QQ$+�ch�6m�A�޴ ϛF�'��$�O��$`ӛa6��'��X�Ά�n`�t�f�J+L�Z]k��'�l(��*�
G��|�t��`�Y<.��7A�+n�Z$G�7i  �Iny"�|r�v�<qK�$a*r(����Q���
a�'k&�'�dey��'A��5O,�v�s�9:�)r��ː3hb��I��(�ӀP�6����1?���`�Qͣ�y��:jz�MywN� ����V��?����?������<!����;?��2�'jQ�A�!8��4@,���?�����|�'�% Sg�\���8s��b�bC�f�Ӧ�m�|���p��v�`�	�6R��$�(����
$�SU ֨C�@8��b�'��R���|��S<C��lT�i
�a��\y��s�L�$�(�ӿR��M���S5"n>�H�ϯh�4)O��y�T��H��?-�	�ul�M{��=Μ1m��y�����jѯ$}��H����+��]M� ����ޞ��C�����ab文O����<1,O��Op�l�!*�I�[a�	@ D؞9W��JD���W�\����?�g?	���Mۙ'�D����Z	J�H!�#�A5��� 
דTZ�m��?���!�H����\I~r�O����"1�$uZs�B*J)�y�pH�%0��'�ay��)���!֐A����3�_��hT�A�|�"vӶ�8���t�ڴ��'���u��b�Nذ��n�:9��'���æ�ߴ�?)�
)�N Γ�?��I {^@x5GߧS:vT�	�+f���3r E�Pw�}2M>9���?�'�?1���?	'��9��ݢ7盻x��TYϐ��?�����^��0�h���I��`�O1�A�!�V]��=�W+�(]t�� ��?A,O4m��M[�'���Q>��%{(uP ���T�+6���$]Z�S�MW-�8�ɠ�Bb}�������Ll�c�t
��.�Ta�N/�I��<9���$6���<��4#ۺ��0Q�@u��Q��<�@�����k~#f���$>�4��D�On���*[6%)1�٘T��V�fӮ��B�16�4S8O��D
==|z��2(;�I^88�D�_�_�lL:���)��'�H��Qy��S
X}�y��^=�@8�'+>d�|�mZ�4�zc��~��5�M�w�����B� �X�[���lgܰ���'-�V5O~��?Q��ן�B�ĭ2n$�?V:^�``j�D�y&/��`�4�IvȄ� 鎙e���E{�O�D�u�ҽʐ�eY�BDI.ע�����d*��\�esh?扶/�H��@=�Hl��cT�P��IA�Ɋ���O.6�q���'Ph)�/�!CM���ᗦv�@��?��.��݋�c~��Oa`�U�G��#(�R�F��{�~h�(��
I�IAy��'H�>�ɠ&�RBJ�Vլ=���
:���R����:?�v�i��O���4Cz-��H���X�0�N#���Ҧ��ݴ�?Iס��l���?%���r�`ݹ@�`�#U�ā�ԧ�R�$hA�<�����O8���O����O���E��0�JҮ8DN�$s)��V��vi�&X"��?��O�����?!c	DU�Hd"��QM�R}�sh���	��M��ia�$2����b�i r�豱��/_3R�����Ttъ�,˓HDb�c�@jxlT�O>�+O���&�Hb���G3+6x����<���?1��?Y(O�n��/[*�C�? X����ş9^����E�fǴ���'�T7M+��#��dWͦ�XsC�˦9`#�<g1��aG�v�����j�<8lDaCy���I��8Dz�I�=eI茔'�����$}�]]I�	�6%�Y�6��!�'qR�'��'��S��Ol���s �#TҊ�#�O[�2P�1��!F9<���'��c��|>OF�$���m%��ڂれ��4��j03�ƈ���P�?Y�O�@m���M���a�J�H]�
���؂)ǿ:w��H�Ë�D����(Q&z2İ����6��$���'0r�'�r�'s<d��D;��ä�(	��%�O��.�bT��R�4e���'��8�/�+Ӵ�U��_��a�ş<���'�F�țF�kӄe�IH��?!jMc@�=Ӕg�( ydlYE̍�6�2�d�NKz%�'�����Gg0��%�䓡{j��Q*�=P��IQ�$B,D��	� �'��������i	�._���yaD���D�����f˂ {��b���4���O8����ԏ"�fa���I%��	`�c���L�܆���2O��D�wB����[���I2	�p���LY�܊��T��b4�	ꟴ����Iៈ�Iɟ��IQ��DҮ"�vTr��Y�xi�G_%,��g��y�'9B���[>��tЙ�� ��탔O�@M�4jś��c��In�����?!���ʔ�tf���I[�h���t��:z�t��6�W؟��Ϭ_q�wK�p�Ilyr�'5L�b�v��Aؔ^��rD��I�'��'��ɣ�M,��?����?ɕN�r�����W����O��?!/O���b}B�p�d���՟(�O����J)`٢"�����Y��?�J&Aɐ@��j����dz>�P��*r�T�yL��䝫's���K�(q����O@�$�Oj�S�O�Ā(Z��i����<�v�� ��r�wӖԁӗ�x�4��'��$�|H1�E	��{��0EeY�;��Mr�h8n�%�M��G
�5�PM�'���B�i�/�XijaK *p?쐧1��Ԩ��'N��'��������,����h�ɝ%$��d���r�ހ����/�d�'XR7Ky���O���-�i�O�(��g�2h�&�1@��}+ ̨S�YR}2ki�ΔmZ�?YJ|����ҁL�e�`J�k��v���k�;��(5F����$ү��	;�&� &�=I���$�@!�+�,u�N1ZW���?�(O�˓��j�������~B���yz8�C���kN�uz!���?��i��O��O��dv�,�I,��,�nL7n�
d"��
9:$��DM^��O�9!�cY-��<H������ٿ��EY�j�rs �	���27����py�[��~z�զ"t쐢D�	d�8�j�' m�	�M�D�@~�
b�2b�����6yV�*F�B�D��v�O���M+a�i�M�<>`S�'RI��\�
��Q�+q�	ua �N����2f� uU9��i>Y�'b�P�P[B�� ��bl��f�#Y]��|�d|��Z4��.�
�m��t:+�>bk0)E�Kxy2i�<!��M��'�O��4�F�{� \�eQ�ɔ�فLޱ�nt���Y���KUn~R�Ox�r��_&`�|�OF�A�K3Mf����˅X� �A"O��R��F9DԤ��4,���}*��\�R� �h��|��ՒÀ�6G���iŭ��Hm���D3F��)X��U�D�2h(�%�w�d��Ȟ�K�d��T���d5����O)r��W�X�x��"H9`Ճ!���F�D���#:�\0��P6>,����&Y$A� �XD֥*�d�4|p T��V/bX�7!�.���RDE_�P`{E��+�����?q3F�	+&�!bv���<����?1���۴[D��b�I$~20����8
��!���'���'�П0�Or_����Ǝ1)>Z��-N����!m��?9���?���/\�0P�9��aH���?aF���ꘘa�]3h��ٻ�̾
�B��H�C8	��?1��?ͧ�?������'S`H�B@�-B���>6:i��'���'�B�'w�I����g���q�.t�7(-2�q��N|վ���V|�\�4>O�I:�b�~���Ǉ�^�$�O&ט3I�2\����M�|Z�k̾6��8�� &������?a���4����O&7�Z7Y6��uL�z>��!O�j)��Izyr�'=��I�Oh7mN�#~�1��I��
Ϥ�P��
F)�p�(C8A��sFO��v���՟�Q�@$D<Z�f��`m���ܥ#�D��,�40��4h��?�*O��d�O����O`��?�ݴ?����ƩJAo�(p��F4L�����'�RR�H����@��5A�b@Z���� ��6�5g����+�=
��!Bp�M�5�q�	؟X�/<� ��S�q����ٟ��	�?un��8D$3׮B!@;� �2�G�ʹ��?	����O�˧�?1�O�Y�$�P/Q�b  �I�
<MڣN��u_��Gx�g�'�<Q�!�=9I��i�L��b1��'ؼՀ��z8ZY�C/l�X1�ۍY�Z9���98
����̖�8e/�w$`!9C!��>HH=` �އM�p�!SA��}��H �?KMX��a�Za(x����:Ɛ!X.Ҁu��G��I@8	��)g��@�_JX}1s�L�@�U���=w��Ag"X�,l�CC�c-�����ldL�G�iTr�'B�O��'M�6�.;'aֵmM�0SP�|2�'LR��#O��'0�U>]�Q��NaęS�`�-mC��A5�K�,�����Db���M�-���D��D��'�Є�&]$|�@ȃ!.@���b��?9��j�(#��?����Ozd��G� 4b Ջ�GC#2f�$���'�đ9�jp�~���O|���� &���I*C<�:Ĉ'h}"� ��N ����I�1����Ο���w�'�?	�C(|xɂdO�[��m�� �1$�a��ib�'��5PO.���O�)� ����c�L\� �)'�Ȱ���'���'(C�G��~��$ƶw���A�ZS���ǆJ3s�1���5.)�Љ`$�{cp�Z&f'�<3"�I�Y����O��$�O��/s`Y�	2Z%H�B�[�n��	/Z�d�O��$�O�d)���O�x��L����I0@��h�+ç�O���O���O��jB3O����O>�$e>�1GgI/=� �㎁2wЕ�g�O��{�6!����?a����9O�9L��=��$��#4�Q �E&G���Oh��OH�O��D�O���O�y�f�I���Q0)�|:ژx��Ox� �<A���?����?I��j٠��Z Z�J���3r����TJN)�$`���Mk�����'�2�'��'���,?���@�'�t��O9�d8#�@K��h�q)ID؞<	B	[�}��a���T�Qv�����8$���f�U���xW�_�TC(�+�H��W�pe��Y�}�օ)��8����P��e���X�H{XPk3J��C� qC��'t4|�PÓ�Gr��k�Iח!p�q����!��EO�\������3\d� ��Z@�u�R5X(�:r��
kC�4y���Zq\�Rcn��9�(X��$�O��$�O���ʺ���?��-Y<��fĞ	SX1�1k�X�6��I�Ar$�b�.Ү�6�iL�6�+gQ���� F�o�<�Y�'ŃӺ�Y$$C��pAԩIU��p�
�O�lڌ��<�an^Ϧ	��d��X,L}�陾TN��R�`���?�#�i�2Z����ٟ�����,fpd8(aH�,s�L����NI�"B�ɑ:(��ӡ�,w/\\����e���'�7�ЦE�'�2��F/z�6���O6-�	z�l�Gn_�sfTQr�11S����;%��e�	֟����\�T�.Zz��P����9A��(�7Q"�ه��(���za�?J5��Z��/�Q�d7�<{Y�hQ���.0���+7El����a��Y�A�W:�(Oz��1�'in7��ݦ���Ӻ���9�� c�&��)��z�Tv?	�����h�T�85J�+h�v����8s�ސ�s�'��	������#�S���xG咧v���-OjԳ�d]զ���Ɵh�OI@̛d�'=�V�S�ژ�SR��
m��D#���%����۬� 6�X�;A4��q�$�?�Or�OȾQ;�l�1z���o]�.�d�O�4�m��Nˊ� #EU�T�N�~��Bż�񫃍�\��]šFA}�_�?�'�|��)�$<����"��BK�9�
��!��X�O#��b� W
��8@I?�Q�����^�Z�2]2�@�G,XNĘw�����韘���$�J_ߟh��ǟ��Iw��nđ�u� �+QtX���T�DMֈ���ќ<`S�W6]�ҹ{ז~r��B�V���'�H��Q��V��á�MA,-*�*Z7�@a�C�������*��'^]��xn�"BlL��wsLY:�&��|���HĦe��,J�ڬ���YU���D�O\6MT�	��lk'�H�3�>L��%��Q]��3�O"�ҦL?4�	!BJ�R;�ᨅ[�\n�MH>Q���:,O
x����~���Q�,��P�&4J��$���T.�O����OP����k���?y�O޶({4�[?\{<١�lDe�.59��yc� �&a�ɞ� ��x� D9���k�'F�p�ug�
G@���'�u��ɑ5w�(X0�$D B��U��S�����o#.�b��˃�zӔYs�Q|h�m�eNI��$�2sI�ǟ�'�����?���L����1����j"��=g��C�	�u~�4p �1}��!S�B 3�v�'-�6m�O^ʓY�p�ۀ�i��'ɛ�l�"Ͳ�N�t����OB�˦���5y�|�D�O��d�)����f��N�.T�U�`�֝�*��rM�B���R&X5;*"?t�?R����)R�"�t�O�r	Bv�H�8xp��b�_�8�b��P�K�bet�z�m�ǟ��;|K��ڥ@W��ԃ�B���Ȝ���?����)K# �d�c�l��m�)�g�˘)��~���;� 	�a��
q��Fg`�j�����һ{V�
�O|��|2s�\��?Q�4 ��sd۟�Ud�HUfVU*���\A�@�
I��l16!Y%Q��X۴�"H��)�
��'Z*�����"�`$�3�f���'}�PT�8sR�z�C�5f�xq��B�JY�y��'z�#�.|J���/7]^���$"�l}Bb�?����?���H�����o���b��N�2P�(}��'�a{r��y�m�������gbŌ��O�,Dz»��T1�g̈́tP`��L�\��E(�՟�	��RE΅O��d�	�\����E8���q+۽�іgI�(��H�Fn�,��s(E�~v��K�$V��O�0����Wy�oJ�*�챹3�XM������L���T�d�����9^�z��K|Z�O� G�˓	��Qsd��#&�2�3�nB�6�,|� D|���dѦz��dτ��gy��'��f���$Q�)R���-���'ǂ�y2�q\dۄ��:��S�k�� ~��Y�'����'z�ɩe��9��iв}{0@��4�(Avc�)��͟4�I՟@�]w���'-��^�d����-�bDjWc >ъ���F���0��@�K�fg�Cp
��I���򄇂�0xb��S�s1`[_�̱ՄT
���1�Ǘ*�Mٱ�Q��r43��2!LF7��1�T�AcŞ��d�@Ҕ]�U�'����T��iC�Ppa �'NV�z�'�v"��Ao���`Mv��O�R޴��]�0aٴ�iDB�'p�� ���V���B���/�}��	���j7L�����ϟ��F�v��4s�)�17u����I�,.OP1fJ��\@���6$3�@r-.Tɨ�<Y���~`�A���/4\B�J_7ָ�#��dc�dZU���~NY1#
91�hQ0���S���'t�O��u�ɊqB
�U���'�^�0���O�i��O�>���D�C6���A�!�npa�E;�O&���r�%��1r�6`��Hu:�`+�S�T�����M���?1/����r��O6�P�z�Ve���W�p����H�{�
E�	�y��p%	Ú;�d ����/�MK(�v��EP�N%;.���-N!Z����\�$�"�YJ��T��CŃ-e�c?͡��X)��Q��I8�| "d�>ه����I��M���H�"<y���#:�5I�*�%��9"�>���=)��^x69	�"\�=�q�M�R�ў�I޴��V��� [��Aڱ �#D�lS��AO�j%��ן���zqjl[t������əO����a܎�4���N�|)2�Y��'ڪIsۓl��@2�E�V��j�J��&��{#9lO����Q�d������6��x2'�;�?�˓X�0�9�"G�5��¤g�$7Ph����Х
�'(@r}��"�X���*'��"|��hC8m�\��M�v4��
5��A^\Y�a���?��?��pl��OT�D|>e�������+�,Q��<9'$�:MQ����^� u�#��i�2�@*^�J�uN
!�z�ySa�����l��aQ˂p q��$ʓ,�Ho��Q?,$`4lA�%��a�q�%k�1�
OFHygk:T�$`%n�U\��"O&���aͅP����Rmѝ#"�=�B�>B�DD�hi��nߟ0�	ަ��D
] __�����(u�r��Pm��?�b���?��?�4�P;�?��yZw��#4�ӃN�J�s���B�ܰ ���׺_��>�WaC���`V�_�<EΜr�;�	*��IڸO�^�K�	!N)֐��{�l��'�h�Ů�X�����g��)�����U�������{2/ʘ���DX�L��4;�5o��aɧ�O=���䇐C���U'�4Qz�U��4��'{��s��E�7���/�N�H�>�P��>qa�׵r hP�9O�8��EJ��h�Z�Y��L%v�`�I��@�ȓ}͸�е��.'��[����%6�Ԇ�x� �3���"e{wa*6�4Q�ȓ5�L5�2�ѕR�@�qf�@�%�F���Dފ��0g�/lsT(q2���{N��ȓ�N�2a�ͽk� ۡ�'2¬�ȓ}c�p1�W�Qs�]HŃ��*�D���]<8�r���F�Qj�d�+4���Z��\+�a;0v�!��Y���E����FܽJ�$�a�m�<4���ȓt;�'�5mjL����4M��ȓk��j�)�/[րYr��[i�5��'��]��-
�/H��HoS�o�l܆ȓ=DpC�AۺH%
����{'\�ȓ^����X
=�� j�i�����*���Y �T
�Pm��]��["��⏍)},���ӛ_@&�ȓai�`q1���#P�Q�t�0}��u�>����E�l�a��G��L��q�ȓDZuq���'�|t��K�&J�ц�,Qh�����r��r!|�	�ȓ	���Ʌ�!]�ԃ��^2������3/�,��k%ȉ�}��9��&]򃅝=	 x��\�P�U��(������	X0�u��ML�g��͇�f^�|���X?��-T��ȇ�1I4UXh�wTୃ���vZ��ȓ1� -sl^= Cؑ�E�L)�}�ȓ2�Ac`���!)�њ����8F�������v�@s�`u�>K�0��ȓt��i�׉ӻ/~z�J��4!k4���Q&��yw�ȯ<bJ��f%݊K�A�ȓme.�у"�
+8��������S�? Ω�bG��sƵ��ψ*,(Sc"OV���Cr���D�Jr��S"O���M�l�t,`!)Z,P�z"O"����� Y~20+��ϵc�(���"O� �AG6DUˆ6�A��"O �U[9�EPG$�,��Mӆ"O�|�`�	z��a��7#B�q�a"O�3�E6��Y��-5�U��"O���5�H�*�@���(��q	�"O���p��- � �ID.Ar: ��	r�jQD���&,�.Icd�4Y����'٨���J^�mg��q��؀�'�Pp�hEL�S�O:�LHC�_(�]��@':{�l�	�'���N����I�?6�}�I�!3D͓}haz��0/���z�T�
_�����#�p?�h�d˴<z��\xT�`m�X^��� D� ���U5"��1H�3��Г�<�(ȊU%�2�'L��}@V�F�,X-3E0���ȓz��$�ΐ~ZHxRa��?\R��r��ȃ"�)�'8\�T�P�w��Z4.�1c&�%�ȓ/,\3�NC�h|%���B8�(%� R6�E����1aB�gu���䗯5�D���,(D�4Y�L:@ׄ���o�S���(#D� +u㔆#�)���:9�����>D��x�fR�������"z�l �E�:D�Ȃ��ؚR^M�#�A� �@��k*D�@ˤJ0c�v���
^	)��8���&D�x�B�@2Ė�: �C�UN��q^B䉌�P��GA(-��1��,6�nB�u;�D*4܂%,��,g�TB�ɻ !�)��7�p�;�ɀLϘB��#���gL޿hɸ��1&�1�C��F���ŋ2-�t5J��%"�B�I+�m{т		$�F�N��n�|B�ɖg#XL��b�Xa�(z#O��fC�ɼT���ֆ\�8�,�R#d��>B�I2$��X��X�	#��PDB�I,�Yʂ˽ T���tֹ��B�	�p�6�J O�~!�̂�k_�oL!���k�V)Xr���[�EzR�@%+!� �VҐ�@Č	)5�<d�7��)O!!��!N��2�$Ҧ]fR �t���7*!��1r�%��NhR�.��D/!��e{���3tSJ��G�3'�!��ϳz5�j#�S�y%\l�`��=IN!��X�?d~4`�X�R�ܜ���N�|�!�Y�:���� E�o���a�-f!�DU�6����fɱ/�Fd1��
+v�!�dX8�q���=[����b�!��(�@鲥"�h)���3z�!�dH�f�8��q%R�����ʫK�!�d՞;|d�Fj���H�87�R��!�$A59#ܠ3�ǎ� l�5Z�K^!�d�!qD�m�,A���!0'�[C!�DJ'�T�ّ�/��UjѦ�v�!�@
NwFl�㏅ vSb\�t!��&�T�G瞾`Y2�tD�&j�!�����pP�pBD�R��R�!�$N�:���6`զKC�1���3S�!�d�0�����T�מp���ۊ!�DArKpa���,1�`�'�$�!�d�t9�j��R+/���3w�
��!�d�3�@p+6�5�8�&�WZ�!򄎹t��˱FC�V�"(�L�!�� �lz��P��ȧ�7TQF�jA"O���O�G<�a�E�k`����"O��ra 4䀸J� ��;] �H�"O�������z��p*Rχ�e�N���"Oh�/"�jdq᠈��"��'�M)T���ܱV�܂y�P�$Dܲj����e�9D�P�e
�FO1`*�1VcBوA�#0�}�T��=���|Z�J0P�~�!�&���\1��,T�<� �!]|��,H�3�8�)�j� 
4� �G�@Ɇ�3�'�"}�'��ԫ%�,rT���D��f�X
�'��9�ʌN8���*����X�șR�����#Y+C�����(,O��P��ǯ,��)2�)�$#D���'���'v�p冫d�^yY��N3O��W�M��yd��W(<�% ٫�p�P� �N�ƹ��A�w�O���ഁM6Z��
�����|�l#� 9z`I�&�-(� �e�<��NV�MX�
��D�c��'"�N`��eff��;�:7yvm�J�O����o�а�qN�i����O��C�$̥#|�8�Lܩ-#P��J�D�G�F'�ֹ*��� !�PY��	�S<�LsD���	����!Ԡn�~���1+|�eªD��*�jG=inb�e��g��|[a�P"N����fF�gY��׽ZRv�2�;��	���I��v"h�;�#C�^�����+KvI�@KWB�;c;8�'f���Uo�B-f�
`�Ř����o�"� ��P2 ༼�Q��P$��I�	T�[���)R���0�O\!� @�kG�E2����T �)��|a� �s(<��BY�)�H@k6+�}1���IX=���6c����  c���X�Uq�"�q�'�
���(ԙ`��� S'����Pe�izs��YTH�30�͢G-�t��4,D��ઊ�_�Zt�e�D���y��T:��>��΅"c�ZU$���'�th��l�d��V0B �@n	<_8ā8�,�/���)������' �H�vJ��O�d(��en�ȓ4�a[biڨr�c��?+x�0��5#����� �6Z$���aƌ7���|�'��y(��y��/�?a�ؕi6hH�Px∍�!e��3�.`~�POc� `�F�%��b@V��ƼQVj@�#`��{�L �?b���Fj�����nF� �ȇ�I�M:|��
Q��l0��ONv��d�Q�[�r�ʐ�H#J����o�����kס �p>��j�#~Ԑ�C�Κ-n�̐���v≝4X�ĩQe\�i�LY �0e��9�̜V�u�'SI�pJ���P�>�Jp(��
G$t��k�j��"�B�Ԡ�vI���-���G!� Id	̨m��=��NѲj�1���a���s02*c��SN��
-9�Ojh<IV"*/V~��p���VPA@fŬF.����
-���`�6n@�:tB�-Sr"=�# T�f�Ԍ��'^��f]������	G
�[���*�3�ę�4u��Fz-�,b'ͽW@�yG�а>S�@� Eά3&e�_��m�H�_���P�5��A���`U�]ʥ@���Ϡ ��q��%ć`��U���'M!򄘄,4R��S�( ���P�E����%�*��O��>��u�SP�$ۮG�1ke׹C��������M!�DG|!��E��@�d��*�r��
�Y@�y`��C�"���ϨO��3�/�e��-GvE{⃍U��|�I4v^a��O�~����+�&ka�����>4�� �m8N�a�dP�)�V`���A����&煒�hO�(	�J��� "��	�T�MA�� VpXɨ����T�!�àa��ի�A�{.�Q&l��+�����⟢}*��	O�x���֛B ���_�<���-v�4⁨����SN�T�<)'I+m�![�%�<B�h�Q�V�<a!��¨� 7JـNMj)�U�P�<I�i�&��o�lh���
R�I^���Oo�t�ѼЫ��.(0SB�*�yr��.bXh�'Dŏ@p���;��'��z��u�\ؚ���wZ01q�E��xG9(���a�,T�	+�G���C�I4=WX!�n� g;j��6탷;zC��,=�
\���I4tE�+U [+�B䉞l��x�C	Y��%�ӷ#�B����1��J�g�|�+μ_o�B�)� |�Ӧ�X�%.ũ�FZ4U{���$"O���ڌ�� 3��Ҥa}"�b@"O�PP�0vI<ݒ�)�8D�ܴ+�"Ote���� �ĹQ"����໕"Ol�A�'� |���Ȓ�d�rmp'"Oʽ��/�=R��GX69�be��"Oy��=�lp�E�&R�Z�Jq"Oh����1f��I��ۚ��0��"O�)�tnG�7�t�"��0u��#d"O�@�s���;R`�I�!2~���"O�j�-}Ơy�ơ ���!�"O��{Ӈ��f�xbK��[�`���"O�� ��߁��%i4
�vB�B�"O�Ó���$�T%�é�|>��"O�`�G�
'�:�HuGE�W^�p*O�ɠD�Cy���U&����'#�1a��<M
Zɨ�*���|j�'>RA�w�_�;l<X��gH+;�V�C�'oڠ�ġ�8w���!�Nl^��I�'Y��9�B��k��؀7��l�Tp�'�&8���-;�~�hp�^���>D��Z���:&��A��ß/'Ƚ�2:D�,J��S�[�<K0�t	���3M:D��2-T�Od1P�!C�����;D�� �aW�1�QrE��R�� $7D�Ě���4o������o�Jt�e�;D�l+pfҧtʈzԎg�����I*D�,��$L3��ӠcG8�̸`2�)D���KIZV8e, �;t˥7o!�d��*����5r�� #Vk�^:!��R�%��Й1�4�f�� ���Py2dGI���fK�LtM�Wٙ�y��!P�t,��*O�M�N1��Y��yR����p�:W��]+B+���y�C�-tQ�ۦB�8F��h������I�v��թBc�Q�`�u��d�J����#�8�x@[�A&�t9aנ<D��H-[P�
��/172�(�  D����H&k4�(P}%�YW��y�j�}����elϦhH�90fk��y�ON'o����h9KS
�yr�e�A�i��XNX��%�T8�y�dʝ}��!aEA�ED��4`��yb/15��U�񌖚@��T��Kч�yr�=?hz)�s�ؿ3����2��)�y�NխG���f�M�+�֑j����yrB¹9?�J� -Z��|�A��yj�`w\s���Q�H�1#���y�ݕ BDH�΋F��Xa�C�(�y��Y9sE��c��..�(p���yM�'�Թ�u���&�Ĝ��R��y"�A�.X1РNY"x�C�yR�uQ��f��v����B��y�d�Q1����˴���zF�S��yb �`U8i���824�Cg���y���lx���
,/d�z���y���U���vH�8pu���Ĉ��y�O�*a��A�R!Q�z����֫�yBIؾ8t���W�o=��S��y�.I��ݱ�!U3e�����@�8�y2a"�����Q�LJ��6���yb�׮�(�B02<҂b�!Q
ZM��f�R��s��� J����挆ȓz�rс��	7���1a��P�ȓ�≘�J�+^�5Bg������S�? l�I��E
NxF�&YZ�ks*Od� ��}�ܸQ%A��-��С�'�f��u�Q��c��I�R��]�'ui����)7l�����@��'r8� ���}��i���R����l�j$��F -}.LH����y����)I�Tar4��"X�JV!�]N�1J����<͎��-F���>��%V�W�"�ّ�̦�l�A�EP��<�����'��QFD�T�6|c��l�=�J>��ꄑ*ִ�D)!�%!���I�'Y^�2V͊ `��!!́d��Q1�'l��q�g�)��!��^�
tP��X<w����|\bG���<��c�/.2�!@�Z�~C�8��J�<��*C<B��t�3�lp���k��'�p���,�?�)p���,��]�PO�uG��	����i >1ٳ�L�1���3����YF����}��nG<� 9!�Ù784X9DJ�$k�a~"j���z����Ƃ[HT���
L��a(`㊃��'K0�u�Q!G��@��ܐ?Pa J>)�� ��wݷe$�-	�����K�NtX�����ҟ�/~qO$I�ϟ�Q����ݢX�3�|������zN���%�z�@-�s�9<O��03mٞ����b�_���x�qOK�-�)B�P�l�)6�M8o��֝���O
��T��*>�B��2(�*n�Q�� <OB��
Ј4	�̋�-�h���� � �J�;�(ؐ�V�<	�x��5u��Ƞ�bA�*��8Ќ��%E`b��F{�OF��uE��c>�рF��^�8`yvΑe
�4H�{�@�E�%�ZG����	ۓ��v��	0ǕfH�+q���QDxb�d��x	p/�<��#E�ԕs��N�<��)�3H����T����q1��k�9���O+�������<��bC"�HL��
"�"e��$�>�?!v�Ԥ@(�a#V"B�,�2���jSl�'攍��G�_q^�r�旐� 1P`�'��DX())2�dL>�ك7� P�u�c��Qsv8�&�8�D}O7}��1o����cW:-:��;��Y2PJxiXF([g��~���<�s\>-!ش~fp�A7��c>U��ˌ*g����JAܓs���b��Y%P9��ʬ@�fU'�$���^wҕ�wʔ%�X� @b�~ҧ���?I���^��)��ɦ�fA �y����Ebѐ��3m.cE`���
��U,-Y�*�:����y��ܣ\�@��`T�lԲ]s�C3O��D�;�F�B%�G�>5��̃��OVq��n		v��"��N���c%<O�Ia��HpMX"W���O��j��E#���ӌ� 2�Q���� �&�\5p����yh��Z�P��܀0JR�'�LY��D����O�˧x�V�"�Y2~4z���" �d�뢢�����=Q�J׬5������W� �� KNw�I�No�	"o�� ʹ`s�!7[�7�=}B�'�7�X�wҎ���E�&��;в͓"S�b�wH�a���_��+6-�<���s�X�x�����t��8X#�X��QqN�����c�ZV=H'�"6n����P�Z��y���[�S ��0��9J��䫟�x��|?Y����o�P$ir@\K�T�{��Ĺ��h��Ur�'�Ĵ��FU�w�N�Y��Vx�]	��U�g�~�
�D/
C���<	��T>QO|U��ʷ/B�kf%��Ph`�B�`+�	t�| y�F�=�*Z7#��n��O�Y�Gȃ�|�v��*����XT�$�O��=<���eG�,2	���Q�U��\���i�
��Y*&�BG�۪;�xP�a�\�v/�y��j�4�����8����sm�
<���P�c�1^����W����@,e�v���?x+�Rc��:R�,|S�� z�=��#Ax�|�?�c\9&�ã
g�������Ϧ�)&ϔ"��OxU@�4_�R���Ow�ѹc��/ov�e��GZ7�
� #�	3�1O�d�����{n �ֆO�Q��q2�EYA�8�Va1� <�X�� �v�J�p@���lJ��'m�
� �T"j�F�
�k:�dk��Ӂ`���B!���-D�1�I�v�>�\�ş?9�cG2g�@1�3m�&�R&�|�� q"�{SV�e��@�D>ʓh�t3��:x�un�<-��-̓q�
0Ie���g�ц�΢(^uE|�E�G�D�$�4q<�E�	���hO���@9A�І+@L� �Ѓ*z�
��S�l��	, < <�֨׍P��n�J(�-�E�پ[*"LA(�5~�qO��F}��
���T@Uo�Stis7A;T�@1��.��'������:��ᚦC��I�ؠ�*O��kȼm<�M{$��?~�F��`͹?������)d����(T�̠;�oe�� !��;a�M�q�
�C�͍.P�n�(���16NХ�����4��S�$P�X��SG,ǞaJ��c�(���?��@5Dr���	2�&@g�'�j�Cǎ�51�;�S�z���SN>9�C�֠�Q��&�'&&���HƏ����*QQˌ�ȓG��<p[?��<�K*>�"�x�ޓAw��VD ��L�,�sՖ[F��`�A?C�ր�	-4��� F$���5`�-�W��<22*,�dT�j�phR��BX�ܐ树7��PPg��Pbtm�o$<O�RTo���tl�O6��̃P��q�ɑ���"O� `ȦGz����O[�Фȣ�|��_/Хʧ	_I�O�(�g�\zmBS�/5kV��'����Fh��.N���͒��:�'��,&�'��t�C��>�E�W'$"��Ȣl����@-Cbh<��+�>b����^�QQ��]�;<2�!2"O�	1���ԍo�T�P%țE�4��^�t�ϓj��- ����"']�|�^�	@>��c�
,m��P#�&D���c�<p ıZc'H8%�4*�#�$Xe��5(���ȟT]����X��8�"��Re\d�v�'GR�V���\Ψ�Ë�:y|�k��/չQC	�g����V�D9}J~b�d 4���:�-
���tk� %Y.$�+Awܓl��鉑��9}HhPr�G�C)'���#T�epN����"�x��'��`��މ^X|}C`�F#o�"�ΓU�8�$Ջu���&�	m�|X!��>�R�Zi�:)����
�c���
�0�5KV��l��?��a	�I�$��!��9#1�F|B�O�S>��'nؔJݚ|ҀKݷ+$�C�=�@3č��.����HЩ]�8ف�D\(�>��E�X�ء�c�yʖ%H�|xꄅ�[t,�p+,�O�A��C�l�P��l�'M{�	y�N��3��8��D^�Y�p��"��&k<h�'Fػ4��'|��b�/S�������!��-����ߟ��@�a�F�]�r�8&��%���P9R����?
��j�]�!�F�9Y���d�P�a(�����*���fAs@���%A�pW�;��2,̞�4�s��4L
�RPl=5��Q���{k.�8���@�'J
����iT�$�O)*�&��.8[$̀�*B+ꘊ{ �Y�"��#EHE}�����tD�Ph,�8C�+�.cR���OK��x����J���	�90�`\4c �"](*��@�S��魨+�b�q����5<��z�U���s"}=�'`f�"��[s�:�	�����n�I�ORt9[?-_>���ܬ��u�g�'�����O��䞾#��z��Ӯ:�RH8��Z�f���9��W�:�_$��u�I�F�n�8�!*�Q�iL���jY ��`mZ�?��|C$�BZ,�h�;l�"#>vǁb��*'A\��ݠ4%�2��On8qBhȄt��b?��П5:��U�81\�h��^; �[��3�������Fq>�ݒ(>�	C���|���I�x�"��Zר���~��	N ��E�u��e͌9�7B�	�@+�Ht�qO�Z ��1�)ib��Ox�J��|b�$U�i�"DhJboL��yR=O4�ᢅ���FTJb �dղh�&L>n��	IdcT��y2 <d$��v耼NJ҈��E"�б�GN�.�$���qO�tP�'�X���!>��R�"S8L�N����*�v��;u�26�͉>�`�FM�]��u`���0r���F�Cb�J�(��� 7����OHU!b/-�&�֝|��ja�ى%<�<���=�bS�O��V֜�>YƋ�#Z�Z��7"f����L�v|��8y�>�����`+���}�D�B��>%?����0Q���s�&˴I�H�X��ӀQ���f�&�ɈHv�l1EK�3v٦L�C�՚&�OXd� ̈́2�2Qx楃QyD��Ք>���C/�r�9���l�d��TNFj<u�&&��3x�I�C�2�"�H+BrYJ�nԚ��; 'Þ`��  tmF�G|2$��PGdd9��7�.!��S'*0� `Ҷ��q��k0t�k��&l9� �{�'$���c�R�i��`�(�{���E�4�Y�6�L:��		}?�#��Z*=Ht�W�ل����"��ЇL7�8u�E_�0�]���L�A�
t9��*}h�ɐ,�Ԡ��F���ɴA��'y��ъ�I����k#�J'l6 P�&C-p��=Q���V�b42FO;A՚9c�	�B�+�P[�oQE�J8���Ii���*㤞��0�c��EV�Y��r�����ɵe$�L��%R�@���L��E��]YB�ٔ	�"D	�&ON��E}��ԅ䞩�`,	*$\�gi�	^�@�	y����H�%>���$�!$���d$"�7�ր�E�& p�酮ԇz���z���
P�h"}�!�I5v����%��ZZUQdOq�'=`82 A0��Tϻ[���:��H6>R䉣aM�d"���E�	�����������c<J5���KN������:�x���D���V��V���\p�,͵��'�p�;gǨq$Lʇ+i��[����<1�����:���0��B�}��nϛE����Q~\Y`�P �P�ؖ��`Ü��ѵE&���-�8��2%xI�ɣ6��t�	~ i"版`)8�	8	׸��#�2����Ã?�6">�D��w: @��J̡F��\��L#Y��O0$xSH7�)�t��H)�9���#M�`��e�='���JQz�'�j<Ѐ���\��;,]ܭ��ӛK"�'�W�ԀR�ܸ�����V[77k*�����914HT`�D�z�tL�F�$Y� ��L!ViW�Έ�E��x��'КE���X	FTx�7ǥvGh���J�s<)ŀ�~b�����w��� ���0$�Z�ڨ	�%R9:{�<��IâP�Ѣ��`�"����CX�l��E�&!�z��Ҋ�66b�t�)�O�h�m-�ha'nX~Bm����*6��@&�4q]���3��&>�C�I��\�B�	08B ZK��`�B�	�%����/d�hlP����e�B�I�#Z��j���=�
�3f
V6�B�I�Kd�
�k@�aa���@	�m��B䉩o���7�	H=��������B�	=f��ء����>�"��c==ɶB�ɽ@���H��Jq��0)�J�Rt�B�I�E��Y�&	,BǨXr����l]�B�3;�d.H�P��. ����"O�D9Jo��PE8%`ā@"O���P
�6��B���>G"�`�0"O>�SǬeޔ���͗8u}l�"O�%�À�:;�����՗t]	�"O6iS�t�,x�%��zb"O�A�G���f'.�y�%y�(��"O e�˙�M��:��ԀK�'�|�U'�h�v=�E����'G��#��ut�ݑ�&ג�N!��'	��
AM�i:�0��{^4��'�|pz�N*s	H����V�E���'���X�/�$�:UH%�U�؂Z�'�h�A��G��ya�����p��'I`��J�Y�����$�3հ!P�'��ŪQ8�p�"�&{�|x�
�')�x��(�?<�)�b�D  y�`
�'��d@T����*�#]C p�;�'�.�Ze+��R"$��B�;t6ps�'�d2fH�%.6�٠#��@\(��'$@��$��>��ъ��8��u��'�@��S��LPB02t�=��'8�I�f˨/� �x jD$#6h�`�'!�EH!��! QД�ޡ#�m�'����,"Ya���c�%-D��'p@%f��M��@�
�Q�'/���MҺ
F���s�H<d�rI�'ӊ ӱ	]�Y-^�b��8Յ�y�Ï�7
���MեN|�R  �=�y�"M�i� 9+B�����'A���y�자vD��f�*T?�����Ĺ�y�$	�>1�PX���;X���ȓ�+�y2�8oIj�1�)<���i�˲�y���7�8�)�[3ʹZ!JJ�y↎3lj�(y'�\A���� I�)�y�9䜤�Bf� -X����'�y��ȰTp$�k�!�z0���y \�yM�p
� �0�S�h�<�1�\w�� �!숎u�vL�ʈL�<�B� )�i$$��`'d���RC�<�ԉاn�V�zCA�L&dU2p�OC�<ys�q������Z�����u�<�#��F��:e�ԇ�N����F�<A�E�;zWLr�!ˋ*-�9��G�<�G ߃PX���KfV X�7�~�<Q8�RJ�$1�b��o�-��x
�'�%r�.�"mr��+ �\�&�Ԓ	�'4�����ޏ%���$L��*�Uy�'s�EJ (V�
���Ч��K3l3�'�Б� �995t����E���"	�'���ٳ$U-m��C��ތCɊ��	�'�Xp���jw�͊�f
<�	�'yX�zV��;���u��0\P"Q!��� �����zlL�������+S"O�9�Q���MIe��1��|��"O�,!A/Q��ir���<���Xa"O�y�$^��|�ӖT�.b�2�"O֍����1�xt�
6@a
`9s"O�u*�C\����s�䃌K- !3"O2�hWcE1�B�a��z�y�"O�X�R@ʜ;��<Za�S�	] Y(�"O�AB�O�cQ8P�VXDx�٧"O����h�� jBGY�Ma"O:1�&⌐57
(�@	̓W�"�3�"O����N�5|8���Q�8w�޵"�"Op���A`弉�(�+f��hB"O�Y1���{�:���G�.+���h�"O��;C/Y$R,�r��)4�NK�"O\�yD$H�pzQ��Fi a"O��ZEd�����׆bJ�X+�"O(U"!�B6d-@c23z4�"O�!a���ةk�A"n��"O�bǘ��L�P��E�d�˲"O����dMFm��+fAҹ+�4D�c"OY�q��#S|�H����C�8�Z5"OT�qB�U�E��0ar`�"O$,����3���4N�b.E�"Of��T���h�F��.I❉"O����
$`/��Q�*B~*ps�"OȤ�Ħ��Sf�����F�
l�Jr"O���ć�;=��1FF#tMT�r�"O�u��	))���+1%��f��M��"Or%RVꄑ.��-ڗ�@Z�"O�YB���-���O�J����"O�Z� �$�d�j2E��k�| �u"Ot*���:D|��G�ܫP�δ��"Ot�s�ZY��� #�ކP���@"O|	�N�.T��1�>a��""O��ְ5N� ��/'��@$"O��'�F� ]�H��/5X4"O�}�׮��CqR<x�x�z��"O�Y ����L;^@�B��f��lX�"O.й�lBL%�UQU�F<y�]�"Ov���T5,0�8���_@�NԹ"O����%X<Tp����A|]¦"Ot���F5����t��m*l-P"O�qY��˷>L �O�R����"O�	R@�Y)k��tА�д\	�yI�"O��i"��'ìPx��ϼd�`"OD��F�pK 혳B���g"O�`A��;�v  TlX�Yq���P"O��dC�)�晘�aEC[���""O�8��I��>d
� ���Y��!���N�r=X�捠_������ЀM�!��M8h�P�ӥC�+i�������#j!���B�y��b�0\��9���?M!��]�JxD|q���R�
Ti�^8�'0h��D!x|�a�W:f J�@
�'�)Q�H�yfp�3�]Y��	�'p�	hq�Y	#X��2�B�`)��'����Iޚ\ ڀ�@�m�z
�'=.x`c�[;&�-�qnA�k#>lP	�'��#��
�� �t��u��'cL�`�ǮU�lX�":q�'�>BRF��*�Lm���)+��J�'��Hȗ�[�(|��ۛ҆��'�V@O�5�Vݰ ��;!z��r��� ���� �	�$�1�aJ�R���P"O2�b�!U�L�J���84��� �"O(�x�,�]���&l��${��	0"O�=�N���TѢ�k��_s�j�"O�!�ӪR]�K�'/j�y�h[�y�"�*M�8ు�.�Ȑ��M��y� L�%�&͑!��n�ՊR���yB�ܡȬ��7���	��c@��y�%Ӄ}�����צv@X�Iƣ�y"� 9~j4\2Ƀ�}ɴLZd���y��XEDH҆BT7@R�D�c���y���w+l0aQ���K� i$Ŕ.�yR�#��[4�@�+�P0���y�b�=Zn�`�AHջ&�8�GN�<�y�@�~�b	����q��x�6��yң�)�^I�5���9YxQ).���yn�:P������+������ya�-�BDB�)K*K�Бg���y2�ў5z�\�
����	4�V��y����i���3���B@�Y�� ��y�Gͤa�H����(%�Ћ�̘��yR��1hp���N���$k��[%�y2� X�윪��bA6��杅�yr�R�(0pgM�_ƞ���$���y-=KZ��u�G*D���z�C��yB�A�r�+�HK&��	0@"��y�X�t��x
�aY,>r�`�*�y����kC༐s�Tbtݒ��@��y`_�&�x@����\gd����y�
�]1*X`T��?�r�J���yR�LbT�{���$@����l֌�y�l�.��oQ	�PTb����yB)�ET�=���#�0E*��N��y"�� p���a���$�}�7ā=�y2�(��)�B�å~�p|�UcE<�yb�Hn1����w�)B2�5�y⥒�nNx�aT�( �`��!�W0�y�M.������{��������yB�J>z��ʰ?y]���`��y�Q�0ӄ��E) #t8��*`Gè�yB$��*��S  HҔ��cQ>�yj_)��)�E���!3$A>�yhB�܄y��٢N�s4A���O�"~�W��"ri��g����d��C�<�èZ-Z�����JT8N�n����BAy��)ʧ	{8��n�:8�<+�&
�(x��cP��Pk�%���d�M
E�����~>����6��*â�f���ȓ:Tڥ����,R��,S[�0e��g� �"7�G�� pfMB���1MJdY� G01��=���X$����R��	����@2D�3���=G����ȓX@=x���Ln�PK�-��F�4����V��`%dT8���չw���ȓU�< ��$9�qGB3B�e�ȓ]���v�N�o�����+�_.�h�ȓA4���C��4m��,j��)Jj���C膥�4ƒ)iĮ�ѥ`�f�؆ȓQ�� �.��(����A���8T���V�L�J!�ݜ�N��%$U;T Nȅȓh��1� ��|�b��f(�P\D�ȓL���AE �#_���rb��/��(��M�.���,$���8�I�(����ȓf�kR�T�N@TN����M��S�? >|h�ka���%-�%hd�w"O X��BĔH���W������d"O��b/�%�v�� �t�N$i�"O@��V����]jiU�
m�C�"O�H�fo�U�x;�F��O�8�G"O�|ҀE�EiH��k�>K�Hx`�"O��.��I��ȃ��mx�"ON]�q���;>��Z�X)�"Or�S�Ή m&�y	�M�Ti��q"O��#O	9�g�XbO�u�&"Oΰc�I��,ha�k�ED����"O����T&#���D*�!G*�h�&"O��!J�7n�����4=J���"O� Y��Gy��( ̀�P��Mr�"O@u�v�6c쮥�a��E�$hj�"Oٲ������@���ac�!��"O8,� X�i��f�_Q�9r�"OB�2Ɍ�(	��B�X]���"OX�P`�S����R��wOv�a7"O
i��o�2#K.C7�!*�Kq"OH�ɗ˒%]P&�e
�g�P�ɑ"O����NE�űb(5�h���"OH���G�}���d��p�T�W"O!����`a3�f[�#֐}IT"OQ/Nbd�1�	*���P�"O���tBH�K<dq�'ɢ��P9�"Ov0SS�[`O�8�K�"O���Ud�;k��4b!��]�P��"O(���6�����ĩ'��E�"O�q)ӯ`.�D�L��z�p�1�"O��l(YGX��J�6R�4���"O��۵��p���%���Y�"Ot�(�$�	Q8Hb��l�M"�"OFiB��%"�4�0-�B$>�91"Ob����
Ns��.y�zL�Ň��yb�ھ1l�YlN�^���Yb���!�D���p���x ��j!L#�!�dE%E��	w�5_�Zڧ O�<�!�dG�Xtƍ���220S�ȑb-!�X�!��}�Yu�V�@l��H�*���|��G�M
k�XA�Rk����=W
lh�+OF�GB�je�����ԅu��^.ӭ��A�ل�B��X�`CE�u(��(`��=D.Մȓcd�)��,u��}��D�;$*0���tLǃ\���4��#RLkF]��7T����P(.?@]B'.��@�ȓ���K6�6|�&}��O�.؅�����
�N���[��T�nC��	����	�L�P\���roB�ɱK��AX&� $
���ƨV0A�
B� A���#N�h2�-�gDҐ�B䉢'P]@WKJ48�Y��Оs54B�I"#n�J5'ވ Q֩˕�,.�lC�	[n�`�U���Fԉh���6MۜB�I�!yؽR��L�"�f�5��-��B��+��h���Q9h���I'hW?p��C��1(��	P*�d^�S\!��Z3"O氺s�
86��,²�_,d�"�"OVE2�� tJ�8�@9C���+�"O�;Ѭ�Q�0Ĳ�� Q���V"O�IA��� �� ��E�"��Q	"O���-�/L�t�rbG��Ht��۠"O����g7_�J���c6�(��"O� pD{�d֝c�X0����73�U�T"O��F� -��K*h����"O0L�T�]�*A�a�&ʑ��"OHyɰc��_�N��#	�DѠpp�"O<��J �S�D�pÇ�>;�xh�"O҄b%��m��x�g�qƶ���"O�İ�.�>`@�`
F�.D]}Ѷ"O�����n� '�M�7f�T�1"O�L:4�>��-s��8���[�"O��z�Č�cBjP`:��M!�"OT�͋96��@��U�L��P"O:�J�K�B� �V�ݡ1k���"O��P�ǒM,i�ND*od܋�"O��s	��m{�� 5͇�u��|�"Obɒ��Q)|�ѻ�fY�<U@�[E"O�5�,A�U��Qs�eЫcM:�A"O�EX�nE��2�����K��!�D�)jx4��A�ŬK$ k"JAL!�d��V�C�,�=0:����V/!�D�6m} 񁑉Ɖ:T(17A��!��.Z���c�)ˣ.���)9P!��P$}F&��I��~�\i��O];!�$ɮ�(B��7x�hPrk]<.��xӐY�'�ߖMx�@�s���]�L��C"O2V���ns���)[2�=	"O>�	T3{�@ۇ*Չ(���"O�S28DaP� ��!L�y��"O��%�)'BI�&i�M�,��v"OHl	�O�}��@"�H]<}��'�!��Y,�m�@H�����h_!�䆧'���RRCǂSy\8:���do!�!.Q�=��E�;d�3��8KH!�dÚ5��i�Ej\R�5�pMj�!�R2�2e�*�����#�V�|$!�,�j�!�K�4F� x�`L@	!���1pe���5aZG斩ce!��F��,�5��z( �{��(eT!򄘀)񶡸��	�&��s l@!�)�(�4%H�c
6h؀�T��O��	]�O��a�d��5H�F����B� �'"�%1��6*qPIK�Y�W�4���OH��DT)0��E�!��P��C��Pyb�G�p���Ս"�tᑔjU�y�dA'A\ 	;`	�KZ� ��bK��y�mF<K�Ÿ�FȢDSM�����yR։M���;%h�ТkS��y��
<xM �Bɉ>���"'N��y2)@6+ Fͫ�G�<J.�k�Ɋ��yr���8��� /,QR�D�u�V#�y�/�;>��xq$ďPFY����'�y�mK�(��X�@��!�8��$E@�yBH_��X���>o>\Ѵ�ȶ�yB.K'E�EӢ�	p��	����*�y�k��/�r4:R��d{��g�����)�O�f@��7�:��Ы����"O���SD����H �^�D����"O<��ƙ[&��3��7^��c"O�p���(z��G\���"O�q
V ܙ"T 8��/1�P��"Oj�ѡ�6H�r�PВ3�� *U"OnM!A��:�OD/�2c"O|�SEE�{��]���ܳ7���ۑ"O�X��#_Y�f(2�
jp��'J!�K�Z-5�c��u��I9<!�� �l0 M ��KR�@&�0���"O&�aM7& �Veԗ)y|��"Of4!� O�#�q�%��0~� �� "ONL�w��};�����ˡ z�x+"O� s�<#��<��J�8Ch�"Or���� �!2�H6kw����"O0�ÁCI}������s��'"O�LᤧUc(���F����x"O$Ћv�ɎI�4�"�^CS�̙�"OԢr�W�|��'*A+;�Zm1"ON��+ŋt� �v��!YjR�(�"Op�#6E20ڲ��oɱWF,���IJ>�mк^A�m�pO��;�A��y®��nf�S��j�n	ó��1�y��|� ���F��Vb(� ��y�Ń�n|�i��GЕQ�t0�w�(�y�& 4QXk��<��L��Ę>�y�,����Q�ӎJ4�v�
���4�y�V�%�|M�V��10���#5��y��.\n0����&B90�M��y��C.oN����НR2 �"�b�,�yb���{UJ8��ϵ^��q�aҐx2�ަq<�(:oU+ ��0	�8��C� l{p���"�()��:�N�
��D{J~:�fU�=��p�n�N���16�R\�<� LI*�t]��N_/�i�B�U�<a"Ұ@*Ly�A�B۠u���Q�<�0 C6:2�È�'��c�!�E�<��(>6�΋+_ �6�v�<тAx���#��#�ɊL�<!���,�`�� "`e��GF�<�g���h�y:�gK��� ���W�<I�]qh!��a�n��bd�M��&�@�����D��!�'Z�&U2���n#D���cܱ�8\�oE�M?�=��� D��:3��4N�z��#�V�)����;D����kB��t��C��`����6�6D�<QQ� k�T� 'G
�d��R�b5D���qc$J)�CsCM�Hp,4�ĭ0D�b�n�HN�"�,�g���ʰ�+D�xZ2
�j�P���m[�:�����,5D�����ҠL�����׻t�=3��2D�(��L�O�f�Ѧ��h��a1D�$�6�56(ȹ�feV�>��v0D����ʦkO����剉v2�:�O1D�$P�@�h���qtc�9&���$1D�4Ham���y'��)s���p�#?I���'�
lR�#ɛ{X�H�0O;�4B�I�G�h�T�X14��0"B�G:C�ɌcL0q�(��Ҙ2D���G��B䉚(���(G!O�q�n��7���6����}�5O��ɘ^] ��Խ$�z��!
I}ȈB��-X�F��Q�_���󬉁o��C�	�8Dqt�L����(���W�`C�J=Td���:��X�W�W�8C�	�8}�-��#*?�ܐ��O�5�C䉶�@�8U ~�p��3�-[D"ORаŌ�9F�����k�ov��2"O�Dj£Td�.]������U�d"OD�&k�{�H�eòF�NP�T"O�u����_�X�B��]y���R"O,�P݉ZE�̉�%[��bQ"O
��ӏ�>&J��qwg�Ϯ�*OP	c1�]�٫BO��m����
��� ��pQe� z�=�D"�Ovp��"O�ݒ��I�P|���M��<)��"O|ؘ!
_�>�b�J�!�9n(�hb"O
�� �K�7��ɺ��\�4��<x "O�@q��ٕ-��h�@+����C"O��J4�\!W�t����|��p"OB{��D�WI�̛րP���"O���g�4x�|����4&����"O�]9�d��#`����Zm�Jћ�"O*܁���u�xTP��/@�P�"O�a�CK0`�(8�Hٝ.ţ�"O�[筙&dB���
	�i2"O��"╲i���eȲ\�2���"O������|H��d�!4�R�c"O"����
g�e�EV�	�̣u"O(�Z0�
�f��5��B�`�v���"O�${ՋѺ2��5���̴CӸ���"OЀ� ):9rt`
�B���s�"Oܐ`��J%U� � J�u��B""O��3��X�h��(Xb�ʛV�]�"O:�h�`	(%�A��`��@��<"O�4�T鑟A~j�toT�z��R�"O*�c��~Д����j4�˱"O�� �,H=\c�8�`Ӥ	c �pW"OL�sq%5��p*���� K�"O�Ljd�H�4 ��b���2�$���"O��쎪"��yQ�L(d��哕"O�QPeΠ`����;�����"O�|�uk�=_��"fEˢY��Ȋ�"O�0���i�<�2���6Eu��e"O9�G'ٿZ�5#G$ؚ+�ʩ�2"O��"$A�;{^$SӠ�i����"O,��F��J�\�q��sy��2d"Ov])��[s� �i��4&`,��"O�t0�!K�I�J�C5��RG:Z�"O4�cF�'ScrE��c�I�e�"O�X���CQ�.	���:FBp���"O0��e ]o�����4����"O�0V�R�Ah�X�V �[,��+�"O��Q�3PL���T#jtT�b"OՋ��S��r\IaK'x�:� s"O���c��C��"�aA�I�Ti�"O^�A@��;�V�"�O@Y�.�{5"O<X��nW�0�<�T.�u���F"O���D����1ۅ^3�:��"OP8p�عx�TH��t�M�"OPqI���,o�x��4��<Z��c"O�lXu�}�
���
eF�Z�"OZ�UrI�]���Q�&_@�Г"O*|Ȅ{�t�K%�mS�,�d"O~H���ȫ%Ja�L��&<��a "O䨚�(�"]7�Y���V0G5�]��"O��[��b 䪰�Ǳ<�Е9�"Op�� Y��KA����S"O��S�m�8�f��6�'�bJ�"O�X�@á��!��M�_Q��R#"O��*2�]�	:p;��~3��qR"O@�P�E�9g�Tm������{�"ONE��D��~{�_�>w�*R"OZ��v�Վ  �YR!�dgl�H�"O^��â�6z��1����4�b��"Of͛B/��l���(A�E�I���"O�0���K3n:�9R��A��v"O���^�4��Z���k7��r"O� F A���K���⚃NȤM)0"O�(�����y��� �^��r"O��c��^�k�H40����Ӓ�#�"O��X�%AC�8CU��#Y�(
2"OX���n�1"��-����29�i:"O�I��$}<)�*G n��"O����E_lҜ�:�)�6���"O��I�,O�g���Ȏy�麧"O�a@�͚4�^�a*]"nAW"O��;Q&Tk`��krC�'L���"OT%�ӈ$���)�&�kT��k"O�����I��6Gb\�b�"O4�s"T	���ב5K\8��"O&�z%�',���[�a׫Фl �"O�����Ԕ�� @���E"O|���BԐB��a+!�O9����"OR�ѡh��Ţ�! ߾K���RR"O*����� A:�E���Ռ�y"	Sj�=��mϰ]>Z jd�H3�y��ĭ�Ƚ��.Y�W:�0$*X*�y�ͧnp���M^e�@)�%��y����TW�݆J�&^#�C�I�0�x]3�ɇ4Pt���W?d��C�5CDT�+F3JJ���k�C�ɵ�ҬANN�j�1�͇��B�I:9�|�Z��/N���ѧD��B��P�V!����B ����
PC�	g��y�[$,�h�j�N̊F�FC䉗h�B�*��uDf,)��DZ� C��'.�-���@�~��°G�JC�	���8��-�� A��3��!*C�ɝX����&Ղ�DȒuݐa���d���#bC�81��w`��WV!�DF3$%b%BT"HG"�PU���]�!�Η��#�OS�B�}��.�U�!���H�pH���Zp�#w@�M�!��xtT���Q'G)$��㌝"v�!�D�*��	�"J�>'��p�T�t�!�ܼ$Z��䇚�7V|!`E-,�!�Z=X�x0���;a5�8�N��q!�d��g�^I�R�M����'�s�!�U9m��p��E {����#!���(kR4xg�D#�����&��B�!��E�p��ZDk
�6�H����	"o�!��N�T��$��
s�U�E��0t!�MR �,�uIgC��s���5 J!�d�	��`�X<
Q���IB!�DCI��M+�ߖn�&�61!��l��@ׯ�;ԊA���%"!�$X�oӘ�W�V	`��a��&�!�D�&�~M)����!�<�h���7V3!���`*ԵJRIȔ�Ը�R��.�!��E�h��hp ���Z����o�(�!�t�<�!  �RBl�/&�!�d"v<�0�ȐQ=��JЍ���!�$F�7shKg$�8B"p����S�!���$lG ��Ȅ�^���h��=S�!򤋿y ֨�Wl��h�$����V$$!�Ε]��u���[�`U�)y(!���`i�@,���%　��W$!�d�D!2�9s�$CՎ�C M�!��J�u��Ez7H�?��њ@ҏY�!���.��` t�I.a�Ri�o��W�!�DZ�w��	X�C�6G��iA����!�� `��dV�a��4Z@D��My
ٰe"O��1�-!ar�cA�Q�:��"O�h����`'H8ӵ_�V��t��"O��G�@,bT��&J��Ʃ3"O`�h	;��(F'F��F\2�"OFdPqO�`�H�A��+q�H�"O��qc���}�
Pa N�x`j��"O�q���R�f�l��ř�\M>@C�"Ox�x��L*m���� 9,P]�"O�eH@�'_��*a#pX�"O��r�#���l�Wcɋ>��@v"OL]��X3��7脽n,���"O��'@9�x N��)|1J�"O���E�{�tRǝ��I��"O�����9��9�6F�0]2VQ�@"O؉Fn�n�9�W�[�Q*�1$"ORB	<d
��@�ђ*mt|�S"O"5����+d��⠜�q^ D:""O���a[��x�$�ZIL���"O�e+��!v��5 g���!#�@)�"OP�ʆ��8-�ʝ���Zo0I0A"O���,´sC@O�f�"O��5
�^�$�U�́5��$��"O�b,ˎo�p���n�$#�"O����iԽiMΘb�ĴZ��<�f"O6ed+[=y;�xB$R)g$��(�"O���@
(tcFL�~���"O� �s*�N��D��k��,��P��"O������7Těb�J�K�`�A"O4y`��Q�Yܪ�� �o.�9c�"OJ0	�P&��hѰ.�*B`��"O�ؑ�ғXd���$} �	�s"OH�K3��QΜ�A��1 \��'"O(���H�/������!�9!"O����œ+�P��!��Z��X'"O�p�VB�HAt0��COI��*O� �`e�<j��Y����`�'?z���e!az\�0A� G�*�'�¨Ype�QxRH�'
�6*�)�'v�(&)��QS���Wj]���`H�'�`�2&ɴdPn #7`
�N>LR�'$�%��ʜ�8/�S�k]�~�P�'	|����/d)�V��|�5)
�'a��WF���kE@$c���	�'}��H�C��1D�Zb��l��'���V(V4Zќ�x��P\$���'���9�a
8'�
H�gdE��H=c�'K(y����^�:���Eݢ��'$~(�g�+���Q�9B�8Ě�'�5��9�e�G�$0ڵ��'Eޭ�e��[�� �a@ֻsȈ`�'�l�y���)����ө�1c�^)��'�2`3�C
��L�x&`׼MY����'V<(�Y�A[�d":�aR�'�:(hƍĻH��)�T�2���'�X}ҷ Ԡ.�\�����1&�2�'�Ɓ�C@�w5Ԋ�(�r�d��'�\@{�,�P͌M( #�&ᖝc�'@0�ڵ�X�W(.��gE�P����'t�q��Ƙ��p!׀�*A),�Y�'R	�Q#�3��IWK��b�
�'�>)iD�X@��V(�shLt�	�'G$*�ٛWb+��N敛a �d�<1D��{źыક!A���g�^�<� �HC�(\:V_�)՗L��%a�"O�M*	ל�RE��KL]"E��"O���@y�0Țg.ڏ_8l%�"O��sV�W�|3�V���� "O�
�ܫ:Y�F��z�q˝z�<�b��"1�mٲ-Y�KTl� �y�<!�
�1E}�IJ'�!nt`�f�q�<�1��y��aՃ �D2dXŁv�<�q��Z�x�)?�h�!`�Zo�<!DGM�e[�0�Y�(���8c�NE�<�vE�F� �ťhQLXHV�I�<a���z�����áFF0���H�<	�ذ�Nt[`o:3����N@�<1gi�8]\��ٱ��J��m���D�<�E��"^��xPj��M�ud��<q��<��A�c���c��9:����<��W#|��$z��7�A�ARG�<��9<$#�Ì�-"�e�B�~�<��+I�,��l�KP3��u�[{�<1��#��K�1Q�|����w�<� f�,[�ج��dĮ+����7��H�<�dJ߃�D�C3�H�)��<z .�@�<�P�>U���e/�_�hZ��H�<qt*Q-�����]�F]i7����y"�2R:=h�i��2��	;`��y�^�⡋��ߌ(g�4�gM�0�yrHS� � ,�'�`��	�yB�V,dR0�"f�#��Z�Fغ�yBD�L1��RM��M,<�v����y�az$��
ٿG� �k�/���y"'�-?O�L��睠pH���6��/�y2����Q9qO��T�������	�yR�R	3�.�u�tN�%x8Rx�'Z��!��ݮ?���G�7D�-��'-1P�܀Lˀ��TɃ�w��'�Pu�D��/�d�C�+A(wy��'��8)6��7 �X��3%�o����'���S �';:3-�'x\~���'�����-�7~ɸ8C�GvLnT)�'�pY#��_�WK����늄:�B���'r���]�f�$A�e.��̲�'"T�#.ʇ_�b��W��>+��y	�']04X�܂@�f����ՍVk2Ԡ�'�8���G �2�<�A� �P��p{�'{����"׵Z�{��O/S@z��'���R�
5���cd�ۊYs-)�'j4u(挊�^�,���L��ea�'ߊ�!��	��F��4y0�	�',�bm�Yp���`�Q�t��1"
�'x��V�\�FK������.i=B4
�'��Isi<V�B��섬d��!��'_���7 ��
���T��`6f���'-<�׮�3+	�Tu`N�Jt�+�'���Y�)Y��yzTL�Ji��i	�'fLl��N�:Sp�xhġ@"/Q����'��!�A͇,7yV)�c�R�.հ�P�'��x�1���h3��MK��� ��|�<!��+)L��:PlPe�ŋa��q�<y��J�>���d�	c�TՓ$�\m�<1B`
Bņ�q�.Z�l�)*�(#T�X)u-C?/V8�%Õ�;�P�f�3D�$���N�K�Fš�!��nZ$�+��-D��+�K)uV��d�$x�&T��[�1ƴ�*� ���~��"O� ��Pƍە6�th�,�+d~M��"O2��V%5:���cN�Ta��� "On�K�jT�"�l�H�lͱt�d�`"Op٣�ˇ�/¡�%��/w]B\K�"OB�'�]�{D��8���NV<��"O8�rQj�1.O����X�\z�"O,���"H�shbDZ'��4����"OP8!�D$f�f)��&ߥ�Bu��"O�M�.K89����C�H0b!�""O�hchU�^8�ucb R�B�"O�xB�G�n��cM*�"O���T�U�X!��g��e(����"O���`� ���r%��qj�y2 [mVN�0��;gruc��ی�yB*��d�>]2�&H�G6e� �yr��� �^A�W�<����X��y(�4�,�%BW�,g�t ׈D��y�O�{���3�I�S�&̓ƅ���yR�[0�ĨX�DD�.Y����y�L�*����F<4�b%��!V��y�͗�s�T�21؃{��6Ȍ��y"�ķ{ϪP0��Wz��	���	:�y�Άz8��D�S#[�[E��y�# �*���Ŧ�)Q��ԁ$c��yRN�3-��<y��:� x��yRjR6@营�CkZ�H�.���y�CQ��k� Ĥ�D|�¡�	�y�@Y'^��2L�,[l�� 2���y�mF�L�RA�U��Z�xb� �y�&��pk�YcFI0��@J)�y��3c�Lp�C�&��p�WgK�y��&����+(h�
�SG��	�y���/H���/Ȅ�붂R��y����o~�����1H2���@��yiZ�����"R0�hI1d�/�yҪQ�)Mf��v���,��2�%��yBiE���@�����R��Y5�y��=�](#���j6� �y�f��v�ԡ+Ud��)Q4�"&ǀ��yB/V#E����@�ZX�s��^�y����S�-������S0BfB䉚r{�#g��+��}{��ԉsc|C䉢Q� �ƬS=q������02�XC䉴����ھq�U� �B�:�L� �/s�@��T��o�2B�	-8�H2�e�B�~�h��$�C䉳7X|�1b�y�r�B�*�T�C�IRC*)06d�3Pd���ll�B�I�J���aŏ>+�\��&���rB�I8�b0�ĊW1]+|ŋ�)W<)z�B䉻XUBl��0m�p��LR�=~B䉴:��!6�rgJ=frnB䉸a���u��'&���5≹#ZjB�I�^P\����d��$؃���D2B䉹Y3ʠ�3E	?ƀ�'�=uR�C䉝a;��c�*�b����I� *Z\C�	���۰	_�=���J��@|bC䉪N��0�f�~�t ��ߣx��B�	��iq�ݛaL@����u<pB䉀Vnĵ����I�R����D��B�	�T؉��.���2������d:�B�#�dxa	1p�̹2ě9H�B�I 9\�$Q�N�C&���B�	=:k�	��н6'�}2���/"��B�)� ���qcҡU��Qh��/%�,L��"O�;�-䚄ـL ����*"O6�jp��v}�@3�L<D�"Oژ+�/e���@`oH S����2"O���'%ʉ4�IX��N ��e�A"O�mj�ĝ� �'C�*l�FE�7"O��B1�R�Lz����Og��a5"O�y�R�N9A��*cᔬu 2x@�"O�-�� �8��i���S�:��p(�"O���!�W��a:q�ö�n��"O���$�wz��D�܅q3�`�3"O8��6K�m���
5'D�<`�!d"O�%Z!`Q�o�*��[�뾠�#"O��EʩW@�[�Cb����"OB�c�  U&bhm�h���"O�;a�V:Fd�P��!�)x�"O4�S2M�����$�QA"O�|��`_�+��� �|�V���"O�����)m�8�B�R��ԥ��"OR�B0��v��RT�Ɋqp�|q7"O����ʲB�`�`UH�oe���w"O& �#���U L<j�j�)	GѲC"OŰ�jV�{�>������A���`"O�c��ilȢĀ��� 8c"O�Ѹ!O
,�z�C`�)x�P�x�"ON ���۳���*��H2g2n�cw"O�#q-����L;u'�݊�C�x�<�!�Jf��6�V3i���4"Fr�<�ы���DRBJ�=:p9 �h�x�<�4�ߌjpf�0��F�|Θ�e`Jl�<�"�f};Ubö�4�ː��f�<��ai��9�J\�]��Ö�x�<!�� E��V��_�xuSS��}�<�F�E�v���I*U�ČhBCW_�<AvA��!g���,�Jx�yQ�Lc�<a2'�"
�`pe�a�
�� Xc�<��B��B�X8
�¹��͐GX��ȓT#,����%�Pe��)]���Թ��@����L* M�9F���Q�*�9�b^����˅MLq��Y�ȓW.T"�N2a�� t녥1ҾY��l��I�"#�,�@�䇤Z*��ȓ��@1�.�7B�Dp�G�X�;�@��ì��Th
g��ȓ��G�,WZB�	�z��I����Y<���׭��0FB�ɾe��`��GM�K^b�֨gf�B�$>a¬H%���9-��eL�k��B�OTȹ�fh��� �0Tu�B�ɒ{�n����ϠQ����b�t��C�	�@2��z�l°x�ʱ��C1o�C�	4]� PXTNM�JͺhC*?�C�I�n��Q$�	�e:m�v���C䉪&3D����{ld��Ç��X��B�I�Ğ� $�ğ2Vqz�Kn��B�ɲ�x �W ɞI `��ēg$�B��T�`Ua`m�.]�}C3��;&�>C��'h�BwS(9v�A�b��BJB�I��r�����9-�i��I�R�hC�IpS��Jʴ\������81FC�	-`|��'����E���euTB�	�{��= �o:Ll���L��BB�7ja�"��ӆL�j͢&�TjhC䉗]�2ۄE�J�r8�`� �C�	4N6��灈1�@�ѧ�f�C�)� �]	P%�$(i��t�$�̸Hg"O�m�g��LE��	^��,�&"O��rhʿ���`aǩ�R���"OV�(���>hTX% އ3���%"O���"�K ��Pe��Y)���"O�H;uk�*�H,���!'��c�"O�\�����#>~�R0,�<M�`�a�"Oj��Վ��Vi!%"�6)���I�"O��
ei^���z�`̑U|�g"O�u+U	V�Q��U���G�bH��"O XA���)�49X'G"b;��9B"O* za	��p�ةb�+�	~^��"O��� ov�a�aJ@ ���"Oj�B���{X�nC�w_�`��"O6��:�J1x4/Q�hJ�['"OL�IէT6��=P�N	5�����"O@L��LބAP�H�NN:�9s�"O@��J_�n��q;�͜���Qs"O
�	��	�]$8�`Tk���X���"O|ȧ!ߥ	�))sl��j�(�"O:]c�S��5ck�f����"O"����T��GI)R��Y�e"Oȕ���.]D8����pB��Q"O*)	�ǟC�P����8*�$"O����gS#��Q�EB̲~��T"O�t~Q�VΕF	<�cB�[�j<!��E�4U��+#�Q?W��!�@/��&!�ϭGn�� ��%k��T�w��q !�$�Cj���MS Rp����MM.&!�� {9$�ч�Ǝ�0���!�=sKp�k�D:s���aȿ?�!�ǁE,Ќ��ַ`�yxQ�V�-�!�䛭MU�ѹÆ�Rh �`@��g�!��Iti���c%�~ ����R+�PyR�^�k������	D^���i�6�y��ǗL]�}��H�WS��@�ϟ��y��/y��:�K�H0�fcȝ�yrhC�r�y�DHD�\�A��6�y���)�FI���G<�T��E���yϙ�k��ۓ�P�4�������y�Ŕ�2ڬr\��9c�P"d���'��!�%!��FH4E�Rdŭ�y2�'#��*���*x��bM�	sNI��'F])�c��\j�Z��2*����'�%Ч��1�r���Dx�'�B,qF���tn���q�p0�'��ڔ"�7w�VxZ@��94����'�f�6��tC)�d!O0`��xS�'�.�A��@\}�������'\� � !�z:HE�AŇ��
Y��' `���D�0�Vy�"BGj�	�'�0�c�31̔A���c�� J�'��d8��ݠ%	
*�aP�'�@����a�J-�!�[�X�� ��'Nˇ��oÆu3�䊚^���"�'�&�`��$YTh��K�Uj���
�'�$1��BY� R�1�$ �w�j9)
�'..�����	5��S��S�a'�B�'�B�⯁�e7���3���^�0*�'/R�0U��4�pZ�M����Z�'T�q�-�8s�D�1�֫R��@a�'px�{d�-����O�����'t�;�fIW�J4�$'�%6
�E3�'��%���˂-dQ4��?5g�8���� ��������- �FA#FÐ�i'"O��A�7Swڅ�c�F��@S"O.l
 HmJ�S��A�<����0"Ov�8�憹tԀ�%�,o�Ty"O���U��Nev�)�N�1r�\�"OZh��a�\y|倲���1E��"Ot�� �,d 0�R�3A�^��G"O��5��L<�H�e��a�,�c"O��Y�e�tKF�k ��@? $��"OepglM��u�k0a#��p�"Ox�$!0b[н�g �t����F"O������9Y���3��.ז9��"O|��ǆ)$�@I��#
�l�)r�"O�iS�-L��sb�^ʚС"O4��Y�rpLh	� �?ɘ���"O���UY+^JeK��a�,9C"Od�q5�	XXl��ʉo�`�4"O�x	Q�ߘZ��u(�'��4��\�"O�4��E)!�E���7~���H"O~9A2��-p<N�q���[mxK`"O�EP#O�	���#2�%Ydp�$"OD{�� )LeR'�[�B��A�3"O��9R����8�sl&6v�b�"O����Ӊ228<��KE>[c��:�"OF���$^�.����%K>�#�"O^=����g,(�'�x��h�"O�JD�
v�ti1 N,l��h�F"O�U��n��i����1�p@�"O�AJ�q�b��g�����#"O$@�@�6+iDi��Η+�z]�G"Ohx`1�H7>�BL3�H.P��E
A"O� �
�S.��k��QJ��]��"O����o�+e�	"�KɑT��@t"O8�J�� �~�8z�DD-|SvH�1"O,1 �ٓ��5(W2���"O^4�t͔�/
e�Ŭ XFƩq"OP�a�'6�hu����;C��0�"O�83��@crUs��$lڢyI�"O� �惕5��hC��U����D"ON`���	:�j�cb���-��R"OJ��O97{媷�C8n̎�3�"O����OW)oݱ��T�v"OL�{��^��F�{�,_�cP�+q"OVQȀʒ�)Ru�2��I|�zB"O�e���J�b�K'Ϛ�^Ң|��"O��F��(E��ˀ.G%��q)�"O�4�'�F�Pٖa����)�� !"O��Xu�&+кݩ3�[�P�`"O�mi��@�M��xb���Y���ӓ*On	:���8T'���@�3C�ڍ��'Ĳ��n�3�p(x���N:����'*�pA�h/G�2y���Q�D,�x�':���#�$(����b��hmV�1�'��	��į=�a�э�Wx6dA�'��d����m	f�`��Q���'.���g��t2��­@V���P�'j>��U^!�J�s�Ɓ?�h�r�'7�e�3��%gnup�dX0
�L�'z�A$�]&D0�Mҹ|��h�'Y���O�)g�zE�6��GZ0�s�'Waٶ�G�Ѐ�h�Yt�D��'`=�t) &$3|Dц���g�~�0�'ۮ���f^�z
�xv� �dp����'Q��R�%�  W&D^�M���� ��{�.I(l���c�Π7���e"OB�E�
�=?t��͛>J�x<@p"O����&/�&�8�+��E�����"O���℄=R�=����4���q7"Oޑ1p6��� [�#vQ�"O��Q`g�Q�8�����Hx�$"O���,�F,bi� yE����"On�cw�͘;xH���!ȥ�Dap"O�hp��`Q6���o�^�B�"O����i4uۢ���o؃I���&"O��� *ju�q#O ��r�($"O���g΀"g��� T�n�z=�w"O��J��L�*R*��W �A�X�"�"O�0�:M����gO<���"�"O@��F�u�������+��	WO����[!��9!��$<�Ek�XE!�ѱOKp�bEȢhi�6\�'!���Rtr�G>��"@�\�Ew!�d֥@9�<�6̏�%F2�X���7 !�ԋ+SZ���*d#bp��L�!��Z9EW hի�5�%Zpk�}!�D��ASRXH2�p�pMs�(M�uQ!��O�jp��1��Y�*��ah�Z@�	U�'��O��ȁꓗ=����-ǵb��C�y�	�0tXZ�tÄ�<<�Ө��yRT�}#�)P��w<)hA�̪�y�@��Jr�����}������9�y��Ɯb'��[s�6*�n�AP��yb!�K<���BY���T�E�y�iLQ��a�̛�Y*$���	� �y2!0Zŀ�xS�^(N6 ����&�yB�ND*�[f�A+ ���k�yri�M
DH�&��5]ve����yr��g��H��7er5 R
��yR��t�5{��=�`�9�&�y��I"$)���ɚ�6fx�!���y��ζ\v�&��8����FA��y��R�?DJ��	+�عӤ�L��y����2��!��l��)��5���Y)�y��S�NR�x-��%�>�
����yR*�
pC��C�X�*(Y;F�֐�y2F�(��%��0K���y�A�.lڐ�g��+�XU×o\��yb�lb.4�ōL�3����\O�Igy��'�T��R���T́B�W1 Uy�'a��!�e�T�<��m1R��	�'����Gb�R�<4B.ŉrz���	�'.�X�cT;t�X�'�|�*(����[��^P�Xv��8��լ�y2oé7��qg**;�uP�ǟ �yBJ�(H�.qd#K�2H�1�C��y⁾*�8����Z�P�*���)�yrj7_���	�j�Z�0<�D��y2�(Tuq���$V�P9�"З�y�aZ�8�8!�2�J-��4���y�Gߕ8�2�Z��%K5�]�&U��y�BTK��9�,Y�O<I�p!���y2�܇dAl0�Tg��~g�ԡ�ۍj7�	Lx�|�t�!�`§]0&���Y�!򄌗"2��xh����qe�<B�!���66�Xe�6�̿D-���UH!D�!�Hu��i��˅Y���&��:�!���(L��k�O:3�W�!�d]<a��qse��r��cܥV�!�� \�����J�*"_��xK�"Ou�a`T	�` ��恭&{��`"O&yrv�F+)�݃�Bnw X(6"O�Y��#,����-��A��"O���fF�7����B�A_�yJ�"O	2���>Y�����jQ�-:�"O�ep�)��W֐����Um�4�"O�I���՘dO�.JT�q�T�	jx�Lz�eפ)Q.��2 |�kVn'D���iX�:_�x�v�;9�4���%D�D� �Z�D1Pe@�mۺ�+b�#D�`�mѱ��
�d����24b!D���(�m�h�cp�K���$`D�<D��{V�]l� ��I�]�f4Ҧn6D�x��Jʐ:+����F�g`Z�Kg�3?��n�����<,��xs.Z�4�����Q+@;��M8]���;R�ϽN�}�ȓ%�`S6�T:	�=��LU�>.M�ȓR# !V�
&D̡3�B���y��e�ꍐ3����N����3M
L�ȓ(�pXS	7+в�2�ѱKf�<�ȓe~>Yq O@�P�b�@%5"r��NC�}+�-D6��"��� Y�H��K��{u�̹p���x� ��Tp��ȓ!�t4�g�CD���g�T�j[(��ȓ@���AW�K��ׂD� ^p ��d'")�&�c��dIF��h�!�(D�i��H*�1��h��qU����*"D��1��$
�1�B�}�2??Ɉ�ᓒF�у�k�	���Q�۸	V*C�	�O�5�����Xi��Wi�. 
C�I:
s��fcX+#~�iס_X
�B�ɂzf`�X3BG�7u���reS�7��B�	0L�|�0(˵L��P�d(60dB��?Cϊ��B@�A*ܓ���l�B�Ik���E�ء'(��ĉ��YצC䉣c��CƓz腃�c�/{y(C�I1��A@�`��)A�P�P�*B�I��$cD�N0�т%��N��C䉂e|,��F��uXĂ���`.�C�ɦBl��K��S�:�8�3���>}�nC�	�yƒi�P.��V��Qa'F3)bC�	
W
\C�!7c\B�'�5v�B䉑�H�f��,�<
qOߍ	vPB�I>C��e�k��a=�$���±,�B��V����ɲD�b`��Ճ��C�I)V���d�Z��qAd�Z�C�X��@���_+�b��K�E^�C�ɾcx챳L�*?�(\�r��e=�C�"!U ܻU�Y�UUF��&Ň��(B�I�Y�(�%B�m5f��E�df�C�ɿyv��)@�ݙ^(�R�I@�+͢C�	�<�q[cm�{L�0sC@�MC�C䉔i�f���öPR.M@u��&dxC�I7r����q	R_F,3�흣,-"C�ɳi�l��1�jLk��1 ]C䉀j�������4z& �� [�rZ�B�I7Pn���gR�`"��!���C�I=Mۖ�Y ��ҹ`�MĊZ�*B�	}
���?*��B� 4r�B�6;^HK�$�u[\+RI@�!ɚC�I�9�.����Q�������޹YC*B�I�jwҩ@VnOL����<,B�ɌJJF �V�3�\p[�`�0?�C�)� "1ӌO�*6L5��ܳ{Ȋ\�A"Ovy�t	�j��R
>��)�'"Of��3@��x�b�;|y@��"O�۵�P�9�nѡ$�Ώ:o�v"O����l��;�PH{���<v��`�F"O�B��t-��@��]6&)�e�0D����	7����7d���Awh)D��Z"� U!��ǥ[{l���B�4D�\)���0Q$cI�v�����B2D�$�oѝx�\�[�BJ<Ed$�rh,D�Pd�Ʒ,h=�6̆�t�4���M?D��
Q3���!��':�SqL*D��KBh��-c�L�Pl�\z�T�&'D���4.�=� ���J��u꤆?D��6�w�f%�cF�-�	`#�>D� ��GN/XC6��!*҆n=ZP��8D�x���@�@ϊ@`ty*D�P���«NH����φ.M�^L�u$(D��1���{���6�3/�.�R�%D�8���ݙR#|HKҡ��	�D,��%D�qU%E�T�����8�@�&"D����b���Rg&��� D�,	��D>G�TUq��
F �5���=D��u���3xNA���w��Ѱs@0D���.V�/�Ő1�� t�IC#-D�����K�o��s�`U.�TY�8D�X���=và�Xc�UMY�a�5	7D��AOߊ(F.���	Պ��A�K(D�@��lU4� �a�0y��$�3D�<1� �,8o�t��D��%y��;D�\�5��1)����&/��d�$"$D����5ZPM��` �Q�� � � D��R��Z�)��?	�`y�2D�����+k��q�J�8 hDb0�-D��uΆ+ͪ�����K7j���n'D��3��@c"jPQN��J&x`��$D����e��CB���1n�q��� �e"D��j�S�%�(��34b��f*"D�(��R�ss�[��\�T�HX4n!D�x��VD�P��Wg�*Љ@�4D���S��̨��F(8bF�?D�8�w º͠�����U7^ 8Ua:D�X����O�ԍ��
�C�7D��H���$�b����]�U1pg#D�L��e���\���犇q���o3D���$m��22�m��(���`��0D����I�?�@e���+
hla��4D��Z%�fx�ς� �P`�1D�h�b�I�T�Nlx�,�Ct}���3D�c�H�?�P�V_�>9S`�2D�`z�n�v!��x��:�j�(`�/D��0dÞQ��8�a�{�=sF!D�h!$�ڥZ���ԩ(�kd�>D��Hv���$�d���[��=D��kc� y<bT����@�ư�3�;D��ۗ�Ry�t���"r^�Q��9D���GלG��ɤM�H�򭃣�7D�DKbi��R������L �䈒I5D�|�w@�؂7A�r�
�2D�
ՎU�#���}�.�5(!�2&�n���M�.mAR�X�!λj�!�d���8���p4B��b�8ti!�dĤZ�-�4%�ZȖy�p�\^[!��H2)c�iHl���P��0S!�� t4�v�@���x@�ꇮps(��0"Ot1C��ߜ{��ܫ���J]���"O���7O��.���pj��DY�"O�<+SE;&KZ �P� �D���"O�u@�,L~�1)u��,:�i�`"Op�˖ �P,�s��"O���e�$�t�XUj�5d�|P�"OPp�6��0{&���� r�����"O�E��F'������Y"O�=�7jݸ-�*5�S���'Q
�"O��;��'k�8�Ä�Z�D1��`"O��`g$'�y�#��� �Q�"O��Pd��~F���GG|d��Z�"Oh-�%����d)#F &3]h��"Of��� 9i.<�Я�8Xԭ �"O��q��7�B`OaH�K�"OV����D�{ ��P/�(<���"Ov��,E�� ��M�E0�-k�"O, ���9U\y���?R��$"O���V�� b]�']M   �"O�1��Ǩ0�J�Z2偿8B�2"OZ]��f4G�P#�4i� �"O> s�� t�`�`!���X�as"O�� ��͕i�L���4{W�m��"O����Ài�"�ӣ�W�V����"O�TЧ$�8=(��0e,MO�U+`"O 麢��>����N?Cd8D��"O��'� �4�*�!э��ER<H�"Oz��5a����[�]4X�X�"O�����ς��\3 ƃ�Kxx�3"O�	�3"�/-���1Ŕ�Ol	��"O���$�K�~�iX2�W)~԰��"O��)�J%W�>�	փ^�w����e"Ox��,u��,�Т�bnxP��"O�����X!K$��#`��._�LZ�"OP0"l^�%|#F͸Pb4e��"O~���,�"� ű�g�o��x�"O�h�bl���1�q��I���u"OJ!��İZ�y���>�hx�t"ORlH���
22# D6zi��03"Op��ᄓ$4�{5�׍;2఩'"O<�8�'K�>� Њa��#C�dy�"O��#D*	%����C���6��qK�"O�堧��!b��� ���N�"�"O"a('�,<T���$J��@9B"O�T�g���D|"�'ƭAt�E�g"OPr�'������c��.Xl	��"O$y�̜*K��R�\�q`�i�"O �FĘ��T�ab�+��xba"O��s�.�����	!T"OHݢt�Ee�@�k�'�  ���$"O���u�#���K��3����"O�\��ʉ5DX�9��M�YB"O="�(��t#DH�,=2��D"O�UI�-��tk�xP��<�a8�"O��/U�"t�AweE�^�l
�"O�r �[�9�R�O|�d"OX!��O�J��k�b�k:�)�"O��!dD�l:�M��BX�HY�@�"O䙠ւ�G���t�H�,���"O�i�gܜvk��*��A�ڇ"O��&�Q�!�v� �P/6v��&"Ol��'�9uZ�óg��]�>HX�"O��H�
2HQ��$�<~G���"O� څu��"��w��=�e�t"Ov��sbźS��\cb��]��d1G"OV�3�G�T�+qa]2yB(� �"OTRC�N�;+���׀�*c1��H�"OB�f�[35���s۬v-B"O`E�T���K���!�;(�� �%"O��KRKL$�0�{���?GH�"O��&G�* 6n<)!�(@9f"Ovy���(wR5��#%��<C!�+y����t�t@���!b�!��s�`=A�N�su� ���^5�!��Ĉ6�T�RTIP8Ԁ��LO#!��߯k�8��	�]`@ZԌJ: !�F�V76ybС�|�T<��,�p!��Z�D��X۶f��0��$�%���!�$ J��W�b�tP1O�)�!�D��^Rb��;sG���HE!��_��xX;2�X  ���I +dG!�Q/j�*�7OT5�JI&	4!��Ԓ'����"�B����1�5 $!����� �
�h��E��1xv!�D@$t3D�zQ�v�ܾ-8�`@"O�E2-�jnh���6v}� s"O8XR���xޒ,P7�_�l���"Ob+��	7�.�e���f�\�
6"O� ��76:]@d��*Nn%PT"O�mcuc�B�8ȱq'�WV�x��"O�e2D��E%z0B���`?����"O�mB�dȧ*��œS��n���s�"O�qsa�V���Ё$
�m�܃"O>ԓg��~�v 3�U�\2���"O�0C�.Ҽph��)Jd!!�"ODt�%ܝ��f�;Y$v�07��W�<�f�D<7aʥY`ǃ�P ݒ&�CR�<aqL��j�4�mƱO�N$�D�PE�<�cG�:ߨ\��w,�)ь�C�<	5ꘒV���*��%�
���|�<��A�sZ����1x�8�1�A{�<�.��3^��4��'>!���Em^n�<ABkB�2�Hj�g�'-c4�sF�<q�#Αr�y��'~�� .�z�<!��C&Ҵ%0& ?Ble��s�<�$�ݷO��h��l�.V^kCD�K�<Qḡ�P�W̓5���W�JO�<��*��P���G�z1�<J��M�<ق�PeP���5�s���C��^�<Q��Ւ`Y��h���pA��1 r�<针
0Yz.ł��_N��Ă!!�j�<I��آ� �����Bl�"��n�<A! �>{�{�o�@X�!4aa�<2�S�}�b j��R�zO��2�F#D���Vo��zZbXhҀ��x�$� D�����'x��vnM�|��Zu� D�H�Iӿc҉H �0SL.����?D�� "k�|;�q����;F�+c�>D��b�I�)[���-D;�&�b��=D�L���@�c�A��#E�:D�x��f�c�.|c�M\(��ؑ5"7D���6�E"��up&L�0���"�E5D����9�H�1ɝ�r��$��J?D��#�L�X�ٱi��5p~�
�	<D��i�&��y�	��U�R���c �:D���Oڪ`  I��X+�N-D�,� �P>D_.�;b�S�y��A�,D�� �-�cѶL��T���]�"t��"O���`A�c*�0W�V���"O�myw��4D���qjćA 1!"O��'�#F�S���S�@a"Oި"bʇ�_2!)�~���{T"O�y���Ιe���r5�O�媥QA"O����Jr���K����z��9��"O�(��I�..o����+w�:]�'"O�٢�
�>j�WgH�hv~R�"O�5YU����$G�,\TTAf"Odi@�/OCv�pǈғy$�5"O�$�3L�/�����,\h| ��"O`��e�_�r�X��2G5_r$��"OR�[�J�7��a�6b�@��S�"Oh10T�F�h�� �bG3eUl��Q"O��S�����c���x_�jU"O� ��Ǫlp��m��{N���"O�����R�ke���F�O)rZ�1�"O�u�c�?K���`�b@$��"O�05�P����Ʒ&[ $�4"O �&l�&4H��I	�j���E"O�Ms���2s
�Be�܊��A!"O0���ō;*���Bu�@�92�AXr"Ozi#b�4*��k� �k#^��a"OH�.
 B=��5 �>G�Q�6"O��{gI�'Z���Q
� |�5"OF�S%��/w��y�3ÜD�"O@�UC
�3U
��-�Z�H�"O�I��@�0�0�k�LWB}�Y�"O*��nA1<����((Bw@�`�"O@ԀfWn�����S�a"O��{GE�|B�CO�A9���"O�����7Tݺ��%��05`���"O��1,ʢ�M1�	��(h��"O
tyrZ"o��	��I�w�Tp�`"O�X[������Er�VD��'$��K���M$& �F*�3me��*��?�ļ<�J~�'x�d$k���s��_�)V�E4j�Q�ȡ��	Y�h�����2C�B���Z�8HԽ��'}����MA���9"�"f��n P#q���cSXb��;��ď�M��O:e���+�P�+dώ�ȴ!#"Op�����-*�l�i�hQ�Q��	Q���6�����f@�6�!!*�o��R;O�E��y�������n�.yi�"O�1%��A�hC�R�/�
 y��3�Ӻ�wR�1���!��8��Qp��@�-ړ�0<ɒk5nh�6/2��hF�S�'{铡�I쟀!$��\Tli*Eg��*� 9G�*D�� `�I fG�P��I�,zf��7"�	�M�O@c�D{ª��rq��gY�;�.���(P�O\�=�O9V=t�;v
I��7�L ¡O4!�E`\#��S�� �z>q���O����P�� Y!���^7y8��O=L�!�ĄKv�l��	A�v���`�\�,t�'3��^8���ć�"�,Ks.�4ZR���.����zZ�T�I&&dX!cQ�SWo�"<���[���d
Eb��ҬiA��S�HC)%8ax2Y���t��V�}ǚ��p+˽6R������z�.�D؟�[�54�&|itĆO� ��׋�OJ�=E�t�**�~�#�,.����so̶8*!��X�`����_���.Вb�!�d�]x�D���E9y}��,�.���
O~5pA�-_�-[��B�n�	)7�
�HO�*�*ݸ��Kz8ISNU,!xh��S�? ^�X� �%�"���$J���C�1�S��y�*�;���W��򅫧ʁ��yRh��wpA���/��Q���N�M��Ob$��O�H���C��Ĵ���p2�2��xr#Y�6��d Z�4j�5BF��/�y���>q�<�CdP<�b;%��/�(O����+kFmIp�Y/i	P�ʐ�Py��!6Ύ���ƙ�.�V��B
�yҊ��O?�a�O|��a5�lz,]�p�8�O��O�`�G�n}��z�
"Ti�u�>!	�M �y�S�پR�=`�D-��E�>���D:}B�(2�bi�q��{8���ǁZ��y�M�_òD)��,{H9(����HO���;�P0�3HP�M��\�FP,�!�$�10����.�/t�p`�C3�!�ę�Rnh�"T �P�9Xu&ގ:R!�F�[�6�����o�x�rb��#C!�$�:2\���2�
�Vv�����C�jA��qӔ�G��<60� �ݡ��Z%L�&�0?�'��I��������a
@D�'\�9���f��!Ju"ps�lד��'�����m��w��aô��k�6$Q�'W��h,�Wh]:#	,ުi�'�p���@�j���ڎ6�B]�'����`�3T�n��f���hi�'�:��'oC�j� �vKK�[�~�
�'(���U&�V�������W�"�1
�'���u��z ��$ ����	�'O�1Z��	�#O�Q1D����j�O���L �|��ӆ�+j�"`+�b�'5�}�����N��7h�`��N7:j,!��A�f��"I�F7Hв�	�`
��D��J��%���k����yB�C�~��cʧ`|V�����y��)��NH7aƇ	�x-Z �ҲV".�����w�(@�LB��2����'ja~"%]�e�dXK�38p����6�yҍ��`�$�H�O���ab��V�yr��CM���(}���)ҧM�y�iK�}����Ǧ�@�:�Ba� �yb�Ԏ Z�LJ���.��]1���y��֡4�a�ȎS���I����O���韈E�O��]�y.�z��ۥSa8�hQ�S�v}x��*�S�OFP�ӆ�
d���H6'��^��@��>	���)N6Z�ղ�aL�Ddr�3�&C��	� �����l������lC��<t�G{�O�t�Dyb��'�th+@� 6 Iy�MD��yR�X�,���+|�fa�a���yrsv�(�)�� ����g�<�y�B@�E��EW�+���jGd�y�)�'@��m7IT�3`��a���:i�扄�#���:	�pj���̞������?)��Ԉ�ƩS����95�A�_u��o���O���6Ib�\�A�lB--V�4��':q W�G�6������#:Z<j�'Өi���S�zK�2� ܌tT}���?�Ic}�=Oz���`��C�z���]Ұ� �#4��;F�ӪFK�E����?@θ���>I��$!�S?1���D��z�B�&h6����B�b�<I�D[!�D@�B�T<dyz��F�'��x�# h�)���:������y"��C,);��<[� ��݊�y��?q��J�dL���4x䎤����df���f5[��a9TN�c��w�!D�� ��f�Z�jX��s�"W�2 S��	P}���ۉ.��,����_�t �7��*�!�D;1����!�vM��Ǯ���4�S�O�.	�֩P	f�H��F�%��'��MHP�Ա&q��E�3b�|��O
��ݴ�اu�6��=�B1j�c]�<}�`�@�#T�B�	�zQ4djtGZ�zA�5#5��:�<�˓s��:'�;+Q8# ƒ[`���hO�>Ej�㔬&��"7�[%�Z(���f�@j�'y.�Q`�K&�J� �I�eenq�/O��N�S�O-��h`H�32��yg��)�d#��yd�)Os�(��(n��"�|�'3a|�,�
V
�h���ڒ|u)�֍@���'���yb����T`�(q�!�t[�!��1O0�=�|
u���(YY���U� \ �Ǎs����$�`c.���l�1�<M#��R�i �Fx�'ےu� �g=������|R:��H>���%}�S�x������σԂA�C��e���^>~~dC�I���dag.#��Y�\�+�~㞀n��y�\���ON�ӒQ��uSWA� 
�'߈">A*O�7����d�nĺw����3��-X[�Y�ȓ?��W�.\j����)c���2�'��ɍ'���jƽ���)�L�W�nC䉷WK؄���[{���u�ۉT�\#>���T6fܒ�p�Q>I�&ܢ�Tx�!�D,?�^!�T���?�lIs'A3R�!�D�)/��Y��C�#n��!"�M�2o�az���8;p�� �T���"L�$R�'}��w̓ߘ'n�[���HG���+�pJpq�
�'�����ʎd:��ek��b�	�' ���"[$�L8IO
��R�'*LYg���U�9�R�0�Ȕ��'��� �F$cPh3�� n�	��'���Ղ׃>P�s��
r����'��p�!g��D���Q�̩����'V�	(#㖁�!)F��[���	�'�@�A���*�8��uƙ�'���'�H��&��z^��pM��t��[�'�bz����ڠb۲>T&�1�'���bRA�Q+�|2`�,:���(�';D} bY��5��f�e]h`a�'����a��VPP���U�+�'��Da��QB(H|*���O",��'���(�mH�Lh�ͱ�4e�]J�'`�\BA*Фl����ΚY[���'�rq6��)tq����#��M$�c�'/,�r�/yu���Ť\�7Ӿ�H�'��٠� �A�PL�/���H	�'�:0�l o���r��^�����'J��_3"��Q�A��^��,`	�'�ܬ��g1M�����1W��9	�'Ͳ1��'�O�V�S0a�&R� ��'񊙱to���4�[7O���!�'����w�^�FaV��s��5~l���'^��d��2c�X8.��Ԇʓ(/�uY�N��L��u���X<��6��d8`��sehāF�Y�aa4�ȓ}����"O�)%t�M1�LE"$��Ćȓ@Lȩ��^�$��	��a��1��g�蘐w��3v�Y��N��aIf���8$��`ڀW�R�2ȼ	\�=��+�^��!gEG�$�W9�)��^F(���K\�`��ETA�\�ȓK��9!�Kمt�1r�ډ[uH��S�? ���3
Ÿu��-��oċ3�xI"O�a:�M��jPA������"O��W��'/��eX�/����"O��y�/�S�҄: �ʶ*w�	�"O���Û 4x�*/T���w"OL�sĀ^�ps�P�.L�,aR��"O�|���@/ pblRf�A�!`�"Oz��3(�X<9��$:4�}R�"O@ء1ȅ��=9%�/r��*O�a��.ͷ/�e�^�R���'��� �N)�tt�Ğ*P�p4�
�'���p��!lKf��Ҋ��1� H
�'���2��	!���� �!�&��	�'��A;aÐ�E�!뙄oh��	�'�i2 �=`\x���(���/D����- U��$"�};�3��"D�����@����[Fb�-�#�.D��J[��lՠW-��6��mcS�'D�8�2���<1v�"�@��(,��b�#D��RD��6S�������N�v�96�,D���f�ȐQa�E���Y��3?D����+� �2e�1���:~�q�=D��fbC7~���I��C�H�b�V.0D�l8%D���%R�����РD.0D����+�VAh�m��PF�5rF�9D�h�G�D�[6Tظ��53j��g*D�(pK�Ter�
R���kYĉ�eH2D��&��fW`�X%�I�nÚ���
=D����B�$޼A*�H<�~� F�&D��xE�W d����$pjY�&9D�Īr(�#�Υ�Ba� bm���*D��ۆ���T�e�pkK�"��,D�Lz&Aˌd�L�zdȽl4���%D�(YaA�]_:ti���HĨd�"D���ˍ�<dȽbr�Z�z�8�J�l D�pcQ�\)B�:�qQ��4)־|pb�>D��j�EM�_�E��_��B�G1D���e挊b�jt��_
p�8�H0,4D����e�6l�]�#�[�E��ݒve5D�|*�Z?���JQʗ���M�#�-D��p��/���:#�׊'�ű#�(D�L:��[
P޴���c� ���T4D���g�4^7��1g�'�m��2D���&aA0_��2�e�m�H��7�$D�8Z��w��0�CY�ʤ�O$D�k�E�5���çX`��\�a� D�X�đ�y�+E��>T��\06�!D���.��XD�tb���0#P�!g�3D���eo^4D����*Ҕ>����/D����L*�e�$o��B�ݶ0�B䉸&b<L#v"Ab$��噧�xB��<r.�ua@M�z�p������n.JB�ɕ4V�3`j�u`x�2 %��zv0B�,"�@ˢ�7r	t9�1E�:B�I�4@�ԯ V�fed�7��C�	�c����P�'�����!��*D�L�I��e���J��T�?�$,�WC'D����ᄐx���z"�O..��i(��$D�<��OD$r�XU`'�<t�[�E#D��@��&g�P�r�z���Do5D�0��P���ˀ擸{�v�!�'D��C���;UNN�c�P�R�`Ul:D��R��by4P!���-^Q�b�,D��a�D1X����D�36]��P�)�d+�O� ƀ�q��1D��j�bP�XNb���	lx�Ē��-�	���f�.%D����ȅ2%��1����"\4�a!D�`�%�K+zHT��d�<�$��5�$D���7GV#.	�M��O�:�*� D� D�lV��#W��!��'ۜE�&p�'>D��c� ��� �҂�,G��")D��S6DPv<�@ǆ�!���0s�&D�P���>*��J��Ƶ:��s��8D�����-`n�)X�m�� ���(-8D� �kH�'��者��
���[�K5D��h�O�6\Cp"�5m�`ĨP�1D�4��A�Y �rS��D$��0D����۰_�ur��C�(`d�-D���W�l����1�S ���P@O*D�$ؓ� �"M�c�D�4
K�͡��'D��1���4Y{�պ���m�rq���%D�X�t�Î@X���'�Of ���6D�,�Ѥ�K6�pRփ�8(��a)D���Cǖ�z���k��ԯa/�����'D�\X0(�)u�^5��ҿF���+*D�{Ѣ�PIPa�n��[�`S�"6D�d��^�*�@XP��*"��ly�A7D�P���*�\�fiU/?������'D�`�f'YI4�$���WĀ�)$D�xKt�ɹ%8<[�
�DP��%$D�0���Z)v'u� ,�9&]8��"D�x��tk�	��C�9RU�0�� D��릂Ud�(��-K�`%PeK;D��	�F�e���U�ɬo���,;D�4Sa�̥
�ԁ��WF xA�#D�T�����`gh��,Ż4H=D��ʖM٥UW�����8hW�T�9D� �r%�:R�1@CG�]�
-�T�5D���燅w9p�J",�$sL��.4D��1G�@|iR ������%?D��1eG�&�m:���Nm��3��)D�,`q� 6R*��1Q�v��
��2D��8� ԁ`j��ÞC���e.D��(碂�qv��D�$5&>�CÃ9D��(�	Oô�����&}��:D���gO��#��}�'.A)b����5D�@�U&
a��<�p��TŲ(���&D�t�[-+���hrl�yS����)D��ID���B�e!ƍ��[1�$"q�"D�h��h�D�hJ��T�+B�qq?D���䪃�Fs�=zR��(:p>��1�>D��C�#.���gK�\?( ���?D�P��ٛS#���[��=� &��y��3 ����Q�*�-� N�,�y�E�}����r��ZX��e\��y�dX�.8��Zg�Ǳ7I��B��;�y�)B�2��)[����tn]x�.�y�lA K��h�FL�h%�-�m�;�yr�V�Dh��͙j�2��!���	l���O���(�o�m�
\#vM����+�'��K�L�.8�L�:�,���D��'��ӋSuޗ�a�d�z�N�B�<��غnx~-�W�LS� =k|�<i�k�-!;��b��
'2iX�/w�<���ֵHt�e���e��w��u�<�¯1�q�Y�(���ۄ�[s�<	��K>�N��k�)0��c`�Rs�<Ӆ�E��8�-�z��VLAd�<� "$[����. p0�Y�|�fi�V"O^h��e�<J���i��;��Cp"O�M�$n�
��� �B;Z��x�"O���h--�0!�2�@�<B.��*O�a�rǂ�r��2$�	!0PY
�'�J�#F�#RΕ��D��zձ�'�h�8���4U\��@�EC�@�P�9�'�6�q"�4S_�����0��t�	�'���JQ	��������.'�����'ז��� @�Ҹ��Ս*{L�0�'{�|�����sZ��� Ӊ:��tY�'?��#iB�1�Z�f�f^� N��D{����^�~�̥����t� !L��yi�:�< ��n��Yu����y%@*�t��'�"`�Z]�����yr��Q3�q)�	��n~�iR4E��y�
N�X��Q���w�࡫&�B��y����2�;g�B8r���v$P!�y��5,Ò�� ��>b�\)��P�y"�ΒF��� ).))�|��A��y�{G �Q�:ITVAeZ��yb,�X4�9Wg��@*������yR(
RB�D�_#�=��
�y���`d�͡4��<O^�B%D��y��@�7�xx00������-��y���ָ0G ��j���a��yR���6�I�CC��}�P��MS��yR(]+\�v��lZ�"���*��_��yBÀF�ؘS�I8��|{����y��E��PH��`֒$�\	@w� �y҈Q�$9�82d���0`wf�.�y��RXh�����ؚ`(�h�y�~��Q�q���	�'��y�.�9[����n�&28e��5�y�+T��]KCf�&tP���EJ��yr�ܩ�re��ɟ�l��ua����y�&5D6}��Ɣ�2\]`1����y�H�|b�D�Pș|�ԝ�QW��yR�pL̐��F�X�ibv�W �y�)�X6(��@���� :�KC�y2ڳs�A��y2R��%̀��y�'�P�)xЬ�3w,P�E���y�)�6?8�!���\�rO"aI���y�D�U�H���B[�|(��@5���yB͆�of@�z�GӢo�H�Eݠ�y¨YC�G�S+k��@��iL��y�ǚ�~��@E��7gF�"T���y�3L����醊�FP񆦉�yR�K�pK�0R�/���<���y��������%	\�!�nѩ�y�ڪj���K��L% ,Ƀ�ӗ�y��W9v@	�!��Z��\)�
ʤ�y���"C�H��еM�e����.�y��\��G�Ւ�r����y���D�P���N�� ۴�И�ybh��[�� �#�W�<�s��y��(VR�ZsD�U�)dD�y��B����K�`�J,S��H�y�ǂ:�8�sS�͢5ْIP'�yBm�Lh$�1�[}����O��y2��mq"��tC���SD_��y�NP�a5�p�7B��pb�!B3���y���;�VY�4��#ԌfjJ��ybK�Ou���w,���|��e!�y
� V�s3h�/X������X/g��c%"O��s��U~<�SV��:~Ҝ0"O����&\EA��ɜ	���"O�UТ���W�����8�h��"O��B+��q�d0x#�%n�2�@�"Ozh2I٤�d�de�/�l= �"O��H5�T�At�鲗��=c�N�`�>����
|�� � U4����h�s��sl@�*FN�<mt:)""[��q��nZ�]c��oOb��E�[2U�ȓT�V<�u�iu,�pE�.4!��|�fxƤ�UhP�Ã���ȓ8��eK7i��^��`J���nM$d�ȓ)��&lҴ{эЯg�6��7Ӽ�IS)��ZѢ�o�����'Ry����<.��xAV
 +����Ej�I��J$��{�m�<ft�ȓ ��d����jj�G��2�$ą�3f��
?a�
�A(ϳF�����}��I�dF�4��kãN�^�\��_f!��`&���Ҡ훂`�t �ȓ2���#�'1T�*� ƶ8uV���e�Ѝ��EL3�l��q��1@��)��Q��⃬]  �����V2X��ȓh�p���dѹd-d*���Ke�a�ȓI�DP�3/�80�µSԱ�ȓ[�\���Ə7p�u2$"C�>4
���i�&�T%ȸB� �W#G�(�zA��n�й6a�<İ�"��#�l��ȓ 
�Ir$	-\T0)��uBVm��`whYU�t� �P0�O��H��� =9�T�����t���L݀�ȓ]O> WI��&@�����Yӈ��ȓsc|��7)��1�ԽH��T+Xvņȓ�ҵ:�@ �R�%p!i����ȓN!�e�7 ��S�����	 �>Ub���}�<����?�4xƩS��`|��_<��"��J�|$�0�秕�[<$p�ȓu��I!�PI��[V�]�Jfh��ȓX1 ���0n�lD�����4U����~�FL�lS>�؝��*%I�`�ȓE���2��T ��)2Q�� j�`��e/bQiUa�<Ka�����H�Ly�ȓᎴ�)Y\Bn�Su!�Jc"|��?mX܈ ��s�KE#˒>]�H�ȓ�@����7.����f��	E�V���7U���C��")��m벩ӽGxx�ȓ0X`x�D�B>	�r,k������ȓ0�X�h�,|dR�@P�E'�$�� c���Q��h3��J ��Q&���}.��`�W�P嚕�d�ӛQ��E~2(Ɔ2�Q>�Q�����5J�H<��Є#(D���ј^8 ���a	20�Y�/����q@L�IqO�>�p�܍*+�q��-��A2�#3D�ڷN�5s<3�����Q�*}2���$0N���P
@�@�=��͈��_�x:����^�{LX	 �F�-������-d�e�6 Ñ�y�N�,��i�,��� ����O��q`ٜ����b�Hpd�����#�(�y&�vw`%�`�7z�.��!���~"�A�����=E�dB�=�rm�bJ��$IFl�
�y��Ѻf�pj�	�<T�������ēx�$		�9s�qk4�B"��L<j��Y�ȓh�9�'$�����9T����ވ�ȓ3�<�q��̇K���{���S�? V���C�l�\!����{K��7"O�l
�M3�,��#]!8���7"OȜp@h�=[lvp#P��,L�6�3�"OР3���/�`�q�.��5�v��"O"���Ӧe�ֹ:��X��M��"O�T�֯K�M�|�b�����з"OĠ2��2�Ȑ�6�]�Tc�$��"O�,H�����Kd�>V���"O��P��ˠf��S�ǕW_�Y�"O$�1��H�����ωs%(A�A"O8�c�ǛE&
���&�w/@`�5"O������9�� ��d޴e�z�+7"O�1�1�B�O>��C��s����"OvA�#�H�0&>�rE�D�.qJ"O�TKFD)uW)a`��9�Tl�"Ot=r��BV�ll��Cߗ$�<��"O���Q8n��1�r��l3a"Ol�+�0�v͘)�+s��M��"O���iAl4���I�y�V��&"O&��`W�]�$)*�Л1�(�!"O�@�V��'�p�Lޓ/�	2"O�=�ь�6nRh��R$n��lң"O��a��4Y1nu �OX�}� �ѱ"OP�I��*� i�����P5��"O�����l�h�7��K�i�"OXY���J�~Q��F%M7���"O�@���y�;����k<�a�"O ,[g��7��poY<w�I�g"O-���
v2������R1��I�"O�Hd�׶c:���Q�:��pF"O��;q(��LqJB�	�o�ЃF"O��z�یe����Ʊ�ޜ�A"O��Zp�74Z��3�'B�LY`�"Olh�!䛒-���0���k��ŢG"Ot���&7�,�X��P�2��H�4"O��r�������#E�xf�B�"Ox�kR�
�PF~UӠdU+'�Ԭ�c"OV8#	�  Pd��&V�]��s4"O,���+t�fPoL�6��pp""O$���$��y�	Ѵ� �nD
1"Opݩ�l�I
�)
�s�Z)�D"O\��JŇ�^��Rf�,q�h9q�"Op=��˂+ EP$)VdP�e0r"O8 ��w#l�ѳ$4t
X�#"OF`�� B�@�(����Ƿ+��%Q�'VX�C�(�ȟ��w���t �/��}= a�!4D�p�lƵj��3D�\�Ib<=zà7�Gn���Y�j֢|2d*޴q[�]Qs��lRZ=�A�<�� D�z�^yq��A4h"8(�N�-F����U�vx@��'�"}�'�V��`/�f`��į@�x�X݃
�'�4�bN�H?NL���q֤x��`ˣ-�"Q��cĥy��m Gm*,O")�"G@�1�t,AwnW�?ЊՑP�';��#�+��j��\�E�ٕ8��򧔕z}h$���dT�Z�ʑ(<���3.�TH�e��6IL��vM�P�6HJ��&��+$$��^u�h�|B��T��U�5]p4��L�<ɡ��&ѡ��]�u�BL�\�`!kӜ	����%]�.�<���O��r�C��?].�����q'�'$���ѭ<�DO /|����)P�n���#��P�O�ԊG��>\�
���->�<,){�lbtqҏ��/����剷 ��4В�^5"Up-Q���f/N�0"M�:Ty(S�̽#�xa�BT�b"������GU`񻀢U�R2�h��C/i��'�`��T�G?8W�X@��.{@�:�O�p��O���10AE��Y�1�#�P��'�
G�Q D��h!��(LS�}#ր�v(`��؍�t����g1�z��t%6�y��ʱ:<��F�F�zO
�(DM���PxB�M�? "�*�f
;ڒ�R��;}�	��i�Sg���c�H�C͌��w��z�(�5F�Y�'Y�p���>^���A�Ξ�����~�Zb�8~bNpӃ�R�,�T�r�/��c�R$�eg�+.�Q�S/�- F��ݰ>g-����ٔ��
~V���GU���<� ��,�]z¢?�
�a/U����'5i�|�ፘ�J��p���޹�ȓro�MQ�[��| a%��h	ȉ`W�ޗC���cA�P�5�f`�pl��PB��8�y7g�5��}Ӑ̟�u8�����Px�H�A0�{�A��P벍�C`=`�c�>q�h���+�*�Q����C5�3�� �xT���W�
5��QxB�N����	�N+���7�H'?cV��__�� N��C��ɨ J�	��I�Ɔ��ha������Yj���s��f�8�!h;+��'�K��p����H��l��<�ì`�,�g蘻��T�]�1��mڔ��p@�hPD�S�yR���U>!�%$t����ݾ=36��eR�]�8hg�Q�;v���c�#�S9>|���w�D���gЫPu�1@�9��Q�'ܚ�a'ńL�>���Ԅu	�I� �X'p^P���Ҋ}�Ta�YX��AB�EE�'��10B
��1���9����a� �	ӓPK�k�4��֮�A����C;�b�� �O~�����Jk�4���'�.���
�8w�<� bf�3?��z�yrF�>��J$�S
Y�B�K'.�!`L)��_>y{�l� �,�����.d�f4�T�3D�(�wkL�-�p@Q�Q�m$D$d2{��,�R��S�)���C@��|4$|��z��ɹ_�d�$�8f���+)D���G��}vx|K'L�7��|�F9|%�9�W��Ww�lH��ʆ�h��	l>޵8E�P�|�L�`T�	)����ѩ&�<����v�us��^���QʐMƎ��w��7VȘ��D�L��I�d�;Y*�P���ў�VdӱG|�0��.��H`�E��r�آ'Ͻc�B�ɱ^�@�F��.�L=]�����Z��4�?E�d�U�:� E�D����n������y"mG�Z~Ÿ��7(�p꟯�y� P< I[��@4B
�I j��ybI�=yBЩ��'�@�r�X �y��G�v��z�/��&佒�+�����hO���@Kt,ڊ<;�HR��|Jh���"O9�b�l`���O�"&a��D!\O2���R%T۞���El���O.8�%���#'��:�J7{�dX`��E�<��V�[��3�.SQެ���fYA�<!�j\�Gĩy2	Y.�)Qcj�P�<�FI�& � �1��%3�r�i�t�<yAi_��:��w"�pr��l�<��@^1i��A�늦��%�c�s�<9��FC��@9�K��wnI8�ʉv�<�@=c�YX#���=U�1@��^�<����1c��S&����p���r�<���$> ��[��dh�5
�,�P�<1�/��� ���N�QE֌!r�Kp�<c� M.Rp0gA��>H�e�m�x�<a�˜'S�@��I`!Hm�<IWBÃ%���*�Aً� �s��d�<��造0a��ä�M�L�)�G'_�<U�\��!K#b�=[��Q�<�'�ӼϺP��n�&�����Uj�<�S,�/*����'b�er�rgy�<��G�J{hm�5�R.^f$HҢ`�N�<�um�8{�
0'�ĶH�ɩ�VK�<�5�\�d�>*5�:3���Fl�K�<y�π6$�DY���;u�&����WE�<yD)N�G��ه�F�E�$l�|�<��I��u	��,��-y	�u�<��R�/ Ԓ@דc��hb��m�<i�E&e�8c��<��0VA�<���e@6��g
-FK<a ��	B�<��@
.V����`�(O�������e�<!֏ϿVp�8j�E*$p����Tb�<� (���E�9l�ȅh L� ([�"O�b���5|��&��h�S�"O���G�Q�vz�CD�ay��8�"O`I�"�!䠘��=l��7"O�:'#G�Pw�yZb�OP0�@"O"a��k���ɆςLHdQU"O:�	��Y�)�^�S	���y "O�̫��O8��a�jW?$�d2"O:�@�ܿ0���t�S0�ΰ��"O���a�(=�̼@�'^3`�2�c�"O:i�@Ur�r�"������"Oj�(���YZ1�v��'n�`��"O6M�u���O|2��&�8��"Ob�!MM��Bu��=����"O*̺s��+}^��
���</���� "O@IC�E�D�xv6�|11"O(�Hւɑs��Pӆe�u"O)�`&�ĵ�cJI"���i7"O&K&��+x
���\�4�fp�q"OYj�S�P���(�jƱyVa*�"O,�*Q��*|������[nEi2"OjW$<34x
� :Nr�d"O�l�eC�h��i�� �6��`"O2����T2�Ib�iD̔k�"O2]h���y*�J����� Y�"ON@�+
�1�B�R�Øz{����"O�	G��ba:�r�"�:4�h�@"Om�R	Y G��`���I��EiB"O|�*�L�-e2��â�mx�\�"O���*ĽZ=*�@ƃ�$'a�<��"O��@Qa��T���ՃDMn���'"O�Ej��]���0`�
1]H1ɷ"O41�a.�wz�3�MJh"�'� |�f��9t|zpjL�`�
�'�.�ѣ��Du�x����Z㔥y�'ш���.��N=���'^J4d��'�d�`�o�
I$��)غRt���'g�1󐅘���0�� &��'@�5�3�2ZŎ�;���++K�\��'�^��
$&3"�Q�-�� p���'[���0��	K��SF͚
����'GTE�p/N ��AfУ]P@�;�'o���G/����`�:T�ш�'���i_�\�I����WR|��'����H{jPˢ�M�E%�%x�'��%���5���
B�C�+,�@�'J|��XM$����J1p�,Ԣ�'e��gi�9��
f�lrd���'��	�"������9`�P�\�	�'ޜ p�圥!�����E3WLdL��'HTJ�'�2���� ��H�J��'�2�S6EK�"@T:�]�C'f��'�5`Q'S:W"�Y)B��<0�(2�'#��Y��nK�h���B=t�2�'�����<v���Ԁ˭�,Y#�'�h!�@��>>ou����L��0�'p��v�P�+����Bg0kw���'�85��U
ت�'U�h��5��'��)��h�5#�؈p��4l����'� C�$�[����u(M�Y�(�I�'�,��"AD����$S�W��e�
�'+
��k�~�X��jI�N6t	a
�'� y�O��Y���w�^�W�|�`�'���:�"6E�r��(F�LT3	��� ����Ok���c�� x����"Oz�� N�8(8�qfə�3DDdp�"OT88bNP%0�@p!�4X�2f"O\i�/ܺ9�P���q6�0S�"O|ɋ�(�h6N`���ޢw���˖"O�$10	�, Z�Ȳ\tNPA"O-Z�aW-%@���
*.h �c"O��` �ɹ-�b͚f,�f��9b"O��[�b��
Z�9qf��>�:���"OF!y&fПO�����Aѧ:�Y��"O����@�5*dc ��~p���"OD\8����K���FǇfv�C�"O��A���fk e˶�ҩ5\!B"O���ꗀZh�I���qa��7"O�pZ�dE~fE�(΄z`�(�"Ojt�׫ۙ�q27�V9m"!J�"O��uM�>�Y���4x"m�e"O$�;U#Q�~��Q�҃nk,�h!"O������v�i�撲3IP��#"O����R�0�h�G��b����"OfpA5�D2-<���+�'&��X�"O8yF�]@�$h�@*P�y���r"O�i��D��IS����j�"OT�96�(u�J%���ĽX�,�#q"O�E1�&�>1�>%���?[y����"O�ƙ
�@�0:�+�F�r��a�ȓH�h�ȂT`�B�.$!~Ą�xb$<�Ώ�w�d]�QA�������Q��)ই�5jy�Ň�zH��*~��� ��~X�T�RM_=L�m�ȓO���Q$W�rF�7MK�#E�Ň�I����w&��.Y��rb�8�����9Z@i��F�%����F�4ɺ���V���YǠȼKuFD������ą�e�I�#M:�m��DP�MZ�l�� �P���/����5��sID	����i���(�"ɛ�b��"�
���(��tHdA��5:��W�3Y8ن�^�j�����^h�����Y���(��;Y�A&�x(�3�W'�h�ȓLΜݨ�+�S�l�j��1]�����"0�5��\��r�(]�>�졆ȓt$����GM-@=Z�O���I�ȓ$@B��U�ȋ9z�N��+�!��B|�las��#_�x���M
ZI�ȓ#��	cN��ք�b �- ���ȓn��1��Ʃ
��
3BG&GK���ȓk�Υ�iF�񆸀M:/TPy��y��5 ֫cJ�X`�Y�@Q���ȓ�Eڑ��I��E�f�
�:)؇ȓ`����RQD`�N��>�ȓ�2$��FM�%n�XA냯
xq��mH�+7'
�*��pV�N H��a�ȓH� ��m�!4��7�
�İ�ȓV�ⵊ� "r��!S�����Hф�.,�l�K'�LȪ�H[:�!��[՚x8�f$7��B�Ȅ7��t�ȓt+^uF��2�|Ȫg�P06n����N�^4j��4�r�Y��}=��ȓ+�p��̐m�J��� �U�`}�ȓk�hY��&	&3�Z�;v�(��܆�K� Q�IGoE�M�#��~IF@�ȓF�y[��]7������Ï|_ �ȓ$�j�3׎^�x8f�C��]�;����S�? �!��I�N*�l�y�LpX�"O�D��F 2�F顂�9�vփj�<)CjO}n$�B�/��R%�(jgH�x�<���܅$�R��4��:Q8�(��	u�<A�
ۮ\=��zN�$�d�Р˂N�<��lǇ\�M�#��6/jlQ�p�<��|��@�	"�A �� t�<Ǎ�6A.�ђ&�j����q�<�c�H�l������
�T�,�Q�h�<Y�.Q��n]��k����4GVB�<���\2|\x抹{���Я
}�<-=���f�� #��q��� I��B䉮FnE!�c
mG��"GN��6�B�I�	��C��΂f䂝sS�In�B�I@x�۶� abi�U��:iB��@LU�� i���ʎ�ivC䉴P]���B�-(���X�"� ��B䉻|��M��@?-AziCp�H�G>�B�I�`����Q�Ϭ�ZͲD�F�&��B�	*l�P$qPB� 8��E�d�pC�I+ ́�2`��C�k(C�I
rIH�)TD��xy�d�%(1aPC��e�X,�$�M�А�e�R�>C�� ��9 Vm��I���sB"�#TC�I�����+Q�T����	vЄB�;b��-��S�)	�����V7w�B�I
Z�<�����p޾��K	�5��C�I,1�8�A�K�bj����F%uN�C䉨s��A�O�5����-'�B��R�S���I`�]���	V"Of���嗍s^h\�3AGc	șKS"O0 �(5��"�&[�k��Y�v"O�Z#%K��P5Qs�Y�=a�lIG"O ��Rd�0.J��r�C�HW��7"Oht�-�=s���(���xE�e3""Op}r�ٰ���@@��r]I"O"$���Er��yE�ʼ^�%K""O0�+rk΃x�i�'�Y�I�-�"O�(�f�TcH��hF�;D��i�"OBȺ3G��6B���֕���t"OZDz�dKT��6��c�J��R"O�� ��YY�Uh�	]՜��"O6���d<V	
uC��b���C"OH��K�6dD��g���z$R�"OL�c�N< H�L	��T��"O�T�A�7>�`��Q�[b�P�"O�}��퍚Nҝ���kd4D��"O���aL�%0�@A"
mv���"O�i:e�\�7Y��+B���:_���V"Ozuc�J5d�H��~���"O`�[��U +
�|���_<qx�٠6"OP C�^C
�l�!)J%����"O��pa�W�`��*����l�&�9�"O� ��,f3���'��uٔ4��"O�5�P�W4Z�@go��jT�� d"O8T��9,�*%Ir��^�P���"O�0 4 $Om m��Q�vLE"O
`�e��/E`I�� �eH��"O$l�ԎEn�@���xV
4D�8�#�q�EҤ.м$뜄ӂ 2D�TX�e�� ��P".�-\&1�ց-D�| �J ��귡�/sB��3�1D�,�B	�w>�� �M� ����m,D�\�TN� N|�
�*���/D�� �=��7��D+P�A*2qh�"O������Q8� ��C�r4@4"O�Dk��h�q	��	.G"O���X"]�D�x�a�$�#"O��[�韤%��]R�ڀiȉ#"Oh#�����%�τY�,��g"OtxEGq����� *}���� "O,Uȥ��,��J�!ʆE�"T0�"On���c��Jmk�Px�Fbr"O =�"DO�N���{6�S%E�p�Q�"O�Lbt�V�^)J��Bm4U��x4"O m�D�L�p5���p&^ ʐ�E"O����2H���F�~2Z� P"OJ�h7"]uɄ�9g(иi&"O,����#��EځÌ���Ȁ�>�D�F�V484�a�^U8�}����U���CM0&�(*2$�d���S5쑝=��"�'���ho��5¢"�f���yCQ���S�j�Mb.��}$$���o�6DH��ۖ�)�tlRV�BY�����0�ඬ�"��0��<�}�ЦQA�R$����pܐY���ay�$�Z��(�h��j�!�z�$&s\ ��'�ĽEy��i�[����'��x��D���� s�eEy2�OljP�e��f�h���ٚ'M�ݩ�℉w����9<����>��d�A,�%�0���)�5c͎l�ʤ؁ �&�.˓4:�㟌E��&X��ɷD�0��IAň��?��kP����Oɤ`4����Q�)����]�A[P$��a_:eRN��Uy����$�*�0|�"g B�P�O'�`���"�Zܓz1D�iٴ)sDI�����pJ(���A�X�9 �͢f� ���놴]d�'�*�����5%2�D2(Z'>��	S���Jc�	 h�Q��|j#mP�#+R}�q��2u
�kǋ�ퟠ1��)�'�6��GdW��H0p$ϮHN����O�O@�g�S:�(��\P�ҽk�5#��Jf�fE��<�����C���Q�p-s#D�O�fUS0�|2dHI���O?dH1���	��[���3Հ�r,O Ȋ��S(g" jBc�82&ey���h.�B �(OQ?�����D'l%!�!4l�A�ٙ�(O���I�|1@l@Qd��gF�r�n@���O�	���)�ĥP�)�z�W�_!�N�y��A�j]q�"�!zd�х�?,�����?*��"�1��C�ɡ7eP�7d�%B��#뇏j�C�I�L$\D�Èċ;��	�5��@�!�d�rR���4�
 풵�6a@�~Z!�DJ9fʺ0�a�%L��H�@��$�!��M�l�\LR�DS��LX)��R�!�� ���0��cd�I(��%�!�$L�dn�	���>j@L+��Z�R�!�ɈH�
�;�A�mQ`�@U�X�!��W,!�N�үS�$�9��j�!�DE;tؼ��
WG�T5�tK��y�!�d�]�r�z�(A�U�f�ժ�x!��Ó!ڼ�
�Ʌ�2%��$F�N!��1T$iu�Y�K� �3.ǆ['!�Dn#��0�΋5�B��a,��z!�d�0�ܰՋ��O��t�� �!��;�U�ש�%��y�&&�n�!��D�T�v���N8�B�u�!�D�+/B\l@�"����0A��F�!�DUtLP�d��[��\��iҢ�!��V/W��}�al�*$��ѹ��d�!�d_3t��6�_�z���9�E-=�!�D �H�Y�.�_o�|ȧ���!�dV�A]شiW�L�M=�yJˀu�!�$ۍ~�R`��A�f7�1x��G�cS!�� ��pT�Z�K�2�FmǗo�
�q�"O8d�F͞� ]¥pƫPx�"O��v��TSc+��o[�4��"O��rFųs�zdYK������"Ozx��H#�X�;u/��i��2C"O�T�����$���*A(��y�"OZ)��Q���5z��G�\��|�"Opđ���,�%��O7܉0"Ov��c���Vr֩�%o�'4��q�"O.8��/�*Qц�D�[�4E`�"O�ܪ���2>��$����?���("O<�8�b� 
��q	3���P6�H"O�=��߰v`J��@0V���U"O�سD�0R�x���H��h��"O^�Z4JB�Lh�7�M�@��P�d"OP���b���t3ee��Q"O$�tH�m��kƣ[#�����"O�u �LH74ڜ�
@c��S�����"Orp"�R	;!J����-[���"�"O���`N�i����&�\-CN�0R�"O ��ǔo�\,CwOPXG�	K�"O�m�
p�F\��D f.\��$"OB�de��B+��X��[�7(���"O8��p̃�`�t�rٳ2��#"O�A�eN'�H�SĐ#N��D��"O�@���]>4�ޅs���<S��"�"O. �pkN�{Ǯt�Tb��!<�ٶ"O�1tN��\bd�q ���"O�%���7oLeZ'��	'��8�w"ON��͈�5�XCR�@�4��L�A"O��إ�9r�R-���""O��RɜD!N��Q�8��(T"O<����2wJɢ���71Dt�"O���e�4�(�a�,�_�$Jv"O:���CY#j!������\��w"O� ���X+jp:Tc�̒$9T��CE"O���'�K �@ 
��B����W"O64Kb��%��,��A�R��Y�q"Ox�[���}߀�E$@	0���y "O��-HBM�d�W���SvP0"O~]�4�K�Utd�f�
�a���g"O	C���<@�ءA��wM̩�E"O
��Bθ<=@ 'a��~�ѣ"O>������� �c�@R����"OP����A�8��N�?����"O��k�6~��4t��A��"O���1a6�0�saI?7��	�1"O��� �V?�y��OUa�&�`�"O}P��H#<�15O+?��y�"O��2 J�F$��")��)Q�"OH�� ��G��;b-��� rr"O�%F��vY�1�Fm_�P�.���"O�;7�C;5ݮ�P�6<�t��"OX�+�iM$/�E�R��)$����"O���r={>"�"���:+��u"O���A�,��x4�:$h"O.��F�L�.��Y�OH�j���V"O���<"�@�@35�:�C�"O�X�v�j,ȉgBD=)�"]"O`�����|:J�I@�ʢeup�3�"Od� �䈺�蕃���\tR�Z�"O�1po��Hl��\_~(X�'DRZ�<�W K"!Gr-B�k��j�`LPZ�<��+F%��<H�#A�'ذ�!f@W�<� ��s�� �;��!k�"O�|�$�_w3�X��4`y��r�"O��@� @�t)dE#%vN�#�"Oxt�ӥQ�nMĵ���SU���"O��S���)e7�XpA'
LR�p�"Ob����R�T#*�qE�3	��"OJI���ԼP� ��2#Ul����"O �� k��s�N���Bʑ���8�"O�違�^�Yd�a8� �Y{漸�"O��% ?8��S�O�+i�|H�"O�cc@,�@�fdE;Cgt0�S"O��zq��^��`��GI
��"O8ik��_�N2�U� Dˍ	D�|��"O��# �qf:��Q�U �6�%"Oe�fF4p�qB��l,��sg"Ob� 5�F�e��P���·c 4��"Ol92b�t��ysT�ڈy%��xV"O�� f����1�!�	L�T1u"O���@�Siȱ��Ά�Va�"O�5�$�ըY��p� /2~ $��"O�-K�eO h#e��}�j`�U"Op�z�*�G�؛���O�Υ��"OD��@�5*�����Ɣ	d�D�f"O�-��횀M�<����A���ڳ"O��X��ׇ~g��&��8g�\�B"Oʁ�a@ޔ>� ś�*{!��Ўi�!��]D��V(I9i�^E*Cc�5O�!��:w� ����g�HX#�$@�	�!�˾QE<�����Mm tK.�!�ԂtlnA�riX�i�="��]�4�!��B
x��4(�́��u��Һ�!�$�S,��&��$�Q"!��6s!��3|X��7���t���C.'O!��j����DGc�	+!�K��!��ܖD���K�aI&Q��m�V�/4w!�dJI5x��5)�#��#��{k!�,e�\�С��-^ f���# 9;h!���� ��R7;��-s&���!���q+F�c��E�~e�ظ��y��|��H�hIS�JJ�>t6	`$����"OteP�eQe�D�G)R���:���D8�\�d�]1zK�j�c؊`S� =D�Yr�z���@E!�>z0�a��y�8C�� ��ĺ/Пr�%h+ː V�C�%הe�1kV�|>Ұ��)K0�`C�	%sx���C��#4�0�Gc	W��B�I�t�<c�Tdע���E�a�B䉒B�V�S��5.$� 0��P5��B�I0�*��+SX��R��0H�C�	�RH~�*� G�����O	���ȓe�fEBFI�r�Ƶ!PlT�K�\l���@�[�<�F��P	�<�����$�U�p�<g��`1�H�A7J��ȓW����拥g�0'��%Z��ȓlH�1+�cP���m��nК
����Zy����A]Ε���[;����>v��ȝ�s�<�kC�"���ȓ`�VM��b�j�X31��q6̄ȓn��YY)��E]��㐥S<nz �ȓM�0��QH�6qk4�ͺqd����3h���V=���Z�G̭xL`$�ȓj������_ht�2cA�+M�	�ȓX��P�	�4s,�����M
	��g$�,г�H�%���$S5N���S�? z�1��r렅B��=	����!"O���V��Ȝe��JM�_�b�x0"Or,"�܏�B�#A�a>aR�"On�i�ߒ�1k�IT*d~���W"O�1)2HI�A�|�*b�r�1�g"O�jTB�jJ�L�1�αl�1ʗ"O��R
L�V� =JQcR�R�`x��"Ovr�-X�M� �q�Aݼt���k�"O�$��H�+Ǹ��v��"���15"O(�rn�E��T�֊/~����"ONA��@>r��hsBi]�@���"O��s�EJ��dH�ƂL��9��"O���2`�\s�9h厰R���z�"O��ՠ�:���f���:$"O��X���k��@U��\�=P�"O
�A��1W�Wc	"�6��u"O�ĺ$�^#RĪ�W,f&� 
U"O� Y�
$;�8-pF��E����"O�Q9�@��"�ds1DJ�E2,���"Oj؇�V0��]���m!pM�"O�|���� ������e)�#�y�K�&K���RVė9O8zQb�ޚ�y��_,���)�'ְA�p�d.�1�y������I`L :ozbu�ɮ�yRܥ�]��C�db��J��yBh"2�l�9�j�+	��8�e]��y�(��B�P��'�!O|������y��,5B�8��DX'A�fF��y�BD�q���a�*�0%1!��
�y���0L���A�z���3�!�=�y"��E(���ϓ
c�e��̕��y�@�%8�lkG���x�NIP��yr�W����c�r=zI"�W�y�`�,� yI�h��<���\��y"�ք
�N�_.y�!O˨�y� R�����!ΐg2��tᗛ�yB�YT�HCu,ݺad �C�A'�y�j*[@��y��ԄD>0��L��y"ʌ&f4"�ԃt��I@� D��yҥ۲Kުy��i�s�Ddه.K��yr��S��L�X�lɰ[��^��y�� �9Tfщ0Q�3�"t�ݑ�y��+��p;7��17�����(�y�	[6��I�����(��f =ј'.b�� ��Eo�����o�D��@�с੐����h�b�C[p9b$�'�B�'8��Y'Ú>V^du�C)���P,��ěs/��7����9v�Ъj�8����W:D{��č:�^X���V�p�x9���Ǐ>�����끅���J@	<w:�
�C�bH�6��n�P�m���M����$S?����[قMY���\)q����'c�O���pp��V�Dܠ���2U�B�;�i3\OV|n:�M�O�A�a�ŮJy�
�U=�@�f^�NQ8��4�?����?ͧ[��h���?���MKT�Ä{l�JfƢB��iiJs��L�&�B�@��c7�m��@��Lm�S�?A��4�a`&�s)L�;�${`�L����Q�@1��Y����F�4�`�)�$,�S�y�Jհd�S��6:��}�J]�[�����O��'�j�2�����3sk׆>z�(!m��!�F�Ђ�G+3�b�'�T�'Y�,{���R6�%�5a�=<IhR�{B}�|<nQ�����4x�*	�p"�g�&\B�Ȗ"oO�|�g�'~j$��gչ���'���'�6��������s���AClР��;o����M #7���$υ*�f7���*[�<��˻x�LXȋ"�E��v���M	���;�ϒ}Ѵ�R���|i��P	O��u�c�1���Z7K�dѓ�|��A�F���k�n�7�޽���MS�W\.u��h$�x����%�<����%�����E�T�K�Ǹ� �I֟��XX��Zq��@u@�����mL
03T���e���|��g�T�)�<I)ء36�&�i��P�1�]>���v`D!I3$���O��$�O�)����O��$�O��5�ԨJ���Dj�$.X]�,�<L˜�������r�%Y���t��LGhQ�P1�F��N ��#��8v�)�Rb"�m��6ˋ���qd�ԸK^���\�V"<a���쟠"۴�d� ����II*":�
��ޯ=&qx��>q���?��Қ�ĭ�318��Q$��K�x�h��<��'a{�-]7Gd~����֔P$��֦ف1�f9o4�M��K��vL C��7��O��$�O����( ��! b�$Hp.��C�9��\C	�OV���OV%��n��|��Ɖ<~2QD��0�i�/z��9'	=��+��?p@4m&���<s������0*��ҩY�#*�`Q��..�D@�<��l���u4x�	?��'úh"�C��#1�'G���%G=g�>4Sa�r��,��?��4f�z7�A>L�]0���N~���	�����4:����'+.�RQ��W@��I�Y ��%������>����?���vK����?���M��	�)ڑ�0H6[E�,ڲ��3��*4>��҃�ݨbuD��SM9=��-�O��D��UAMz�<d��97Wp���O]�fg$ٴ��(tGbL�p�&��ًVA@M��r	λM��AB�mT7Gh���Cˈ�������'0@7Q������,z�>� ,*�&dۄiS�M��`	��
R�'�Ob"?A�&Z�L�z�ꒀ$�J���+iܓ.��Cv�ڒO �)�� 6흕�����b	d)���B�����>��� 
  ��   e  4       �+  f7  O?  �I  (U  j[  �a  h  ]n  �t  �z  &�  i�  ��  �  2�  ��  צ  �  Z�  ��  �  -�  ��  �  8�  ��  �  X�  ��  ��  � B	 �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�rdFz�Q�`�'�@o�	�*�)�D���	�%��	�OP���,�2��AK�}fԠ�2�Sp1O)l��y�S�`l
)��S��fE �6�����B|*����;�	�D����&�!3��ѐ���c�� Y�~�b��}��?a�bW�W����q嚱xNCb/�Mx��A�Zy�X��A90��
P�T� H���4 ��ԥ�4H��`y� �+	B0�*G#*�D-�S�'q
:-�b�� @٥�'Wǂ1�ȓc�8�y0�n�&���@,t�^��vC��Ezʟ��'�(���,�B�qE�|���'�`��R��D �uN�i/�51�M*}b�>%>y�<��( :l.��1p��
T��CR(^�'���OZ��ڂl+�Y�͟�xd��a�?oI!�T*D,�=�.����� �Py"�)��m�f {� �!�\�t.<�y�I�$�b���ҧqED�X����d9�O0|�1�_����c�>n�����'��Iv��/|��  �ۃ/��d�@:X��B�I#c��Q;�½��2G.ԫ
��OZ�=yʜq���6���惕{¤����B+/;�	o��,&`��t�d�9��(5$���!�O�I��y21ORc?��Oô�i�O^�L(*Q�M�J��9�U�'8�d�[��M���ׂ |`�	p��<0�!���k��\�#i�/o
��v�ٰEr!�ę���4�����8AX'�eQ��E{*���r�m��F)��I���R��	C��'�ɧ� ��h��~�
 ��	M�Z��LkET�̅�	I���X�I�~�ր���8y2����8?�Íe6�@���j��yq*T�h0�@��EPN8�J�9%��<r�e(�F����'(
8 ҏH����@Ќ]�$�Х��	O�':�5��!:w\��ҕ�I�<!gB�<]xT�v%�
�\}��WF��$���"J m,B"-�V	�q-!D�Hh�d�J<U�uh�� ��:�J;�Or�q�" ?�1���G)Y�¥�ꉳ�BB�I�Ly���&U��T���ƀ5�t�D+�|�ў�)���؝�b����S�O5\Opb�PQʗ��\!h�{s6pd(���F{��	�-_z�śv���L���s�1��|b�xb藟qMCfO°wk:h㓣N3�yO�>.~��V�y�|���!Z��yb�+ �
rTh�p�p�S�9�y��H�Fp8�(��k=6������yBH�]�X#�Æ]EfD�`����yB*H�`D��ᓋ�*km�8�V���'�k:�)�)%N����A
q�İ�v�.s��Oʢ=�~J�J\G��yb�>Vr�P���s�<��AY�oBTA�a� І�Z�����hO?�	&��!�$Ɯ:& �iU�B�	.H���q5 ͡M��8sY7w;�C�Ɏ�J��4�Զ;X�AWꗚ�NC�%�
HgL<D�ipP@�-%NC�I.Nb졂ӡ��;���q�
יByC�I/^�L�p�_�	
�y�!`FC�Inڠ�:E�7.X��mqm�?���I�.�b��C��j�^���i(~|!�$ß{���˒&�2��Erԡ��-���^��H�����]�v������zB(�"O�x�֠�/~B���%�1�:Y��|�'ffD�&�z ���C<O�T�Q	��y�N��M�F��H�����)�#�y���FN:d�5%حv��@� ��Oj�~����0,8���61�:i�"��`�<�%������
5b�����SE�<�W*_4h0Ɯc�C�\�pHQ7�]@�<�ԃI*<��#3��E3�5��M|�<	��[ J]0��@	J!&�~�<ّ`_�`t&A�2�[AdLC�	C�<��D�FBJ���
b��\j�!])�?q#Ĩ�bT�O���d��lj S�
�z�2�+�7w���' D�܁�'&�Z����AΌ��KYE�'��aڷ哠D��r�/�Y�����!	�2�&��d5?y'�M^8��%JR8QhIp$�G�h�D���K�mE�� !���X��F�F�w!�D��l|x�� }��d��/R2e!�������"I��\�s��TW�R9Oδ�G�	�Z\��GܼR�p�iv"O�dAӈ�#)`����_)J�b�C��Is>��K<�m��BX0"��|�a�(D���Z8'N��H&ŀ�A
b�zT����x��]+ϼ(@Щ�� ꞡ�����y��J�)������:q��u�N��y�R�6X��p�Jo`��+�8�?y�O���]y*��b>�yEgP�mt"-�J�� ��E��H(<��4X��@kD^��#Qi�}Zq�O��	r���'�l�S�Y7�(�mح\>�\�瓐�b7��h��H�> j�!$BOȾ��$&Nqxí�N:$��.�=/@�ȓz��	�#4-��b�S�R>���S�? 4h��j��"�r��0"��!�'�IC�S�O�d�a� G�Q��R5�fǦ��"OH,�b�O3�D�@e�D-�`�2�>	�tD}���˦}5�m3a�ѥX :]���?q%�̆#���X�O�3�9j�b}�<�ǨĲ�r(j�I�?��0QaGx�'i����i���S���-�̘�f��<]򄙳&Vg�����΀5� b���Bb�9YS���J>a|r�|rI�=>lʱ��/u��Y1l�=�xR�'`��4O�Q�潫�@��@0� �����ȟ�mS�^�.��ć�4���O�)��ʆ�$Ԕѻf�W�>Hj�QpE�ܟ���2���`�� -�R�*Fc��GČ%����ē�(��Y�M�='�|��J&NH�f"O�i��e_24 �"Q���`k�04��D=}�1O��?�cJ�;IҰt��L=�<h�ڟ4���+�|h��g� �r�r�JU<��l���1��'�*ub��B/(����d
��C-�,�˓�(Oh�C&bsD0����x�|!T�$d !,O���yʟ,�'��a�EoD)2�
��L�(�dߓ�'(�P��P�8�0OĆSH]���'"<O����O� ��
�HP��*0��'��w�i�V��'`��>O����g?٥�C�:!H )�.��"�m��U�<�"��й�񨞂p���r���P}��)ҧN��[�E�lde��̇+[�L)��#P,�U�6�b����c�@%�4����%�qG�<��,�����i�`B�I�N8�)8�\�G������;8B�IOa6=�B-֧D![��Lx���=Y�{��x�-�C��xp��T�J�������M3�'O����Ӷ{eT��cM�
�4��'�T3P� :�B�/Ɲz��'�zuH �E(f� �;�0`�'sʉE�$4��:7 �,4ڽ��'�^�C�(�"DbT��l̲L�^,��'΄)zäT-m"h4�%�!?P`��'6��VA�<b,~D���"m��a�'�1[�*��GN�a�X��H�'0(�����4h���H�' Q�
�'�h%�r�]�,cl����rɒ։�d�<i����q�P����9O!RLh��Fb�<�F*�';�^	8` +�N1�E.�c�<��f���(c�.'B�4�ӣ��\�<�`�A=��HS/��Yx���&V\�<�1 T!�����jǈ~�lx�7`MN�<���=t�d���|/�ɂ���c�<�qȋ�m`�5S��&w�v*d(x�<�Ch ��R-���$n����b��x�<��B�:�*��,נ*��q��w�<QO�9"g�<����>�(g'Hu�<9�'�[�D�	S��cd]��IOq�<ٰ��4�kU�Q.�ʤ�w�<����,z �&&�i"f���*�v�<A�EӦ>�Bv!�Y�6�S��v�<�d�G�i֬�Z�J,ql�qK�[�<��m��^�@q+.yܢE9��V�<�GcO�"�~���4d�Й[�QR�<I��ϵ(�d\0���2r[d\���y�<����Z�j�
P0L-��"wDq�<𦑒
ʁb�FG�K1�Q���c�<i�L����	�(|���9w�S�<���-~�2`��Jp�4��E�<���&1�<R��$5z��B!�D�<���2Tqy%�^H�����j~�<� ��'�ε$�b�Gs~���"Oz-���L�]�"�Z�;v�3b"O�8`����0�"L{�bخqpP��"O������TKI2f4XZ�"O�hC�M�3 ��b�ɀ�c��&�'��P���Iٟ��џ��	���=M,ʓ�8[,C� �I��I���I����ǟ�I��T�	۟\�	�ǾI�d�Y`�<��"�� ���������	ޟ����h��������.<xs*�&�A8�a�7u�����I��������I��������I�0D�t8�J��S����P��`�	����ٟ���џP�������ߟ0�ɋJ���4���9Z�ͪ3�:��	ȟ�	����џ��	����۟P�I�Q*@p�UnR'�Fi���N�;����ß �	�$��۟��؟��	ܟ�	���=�r��(T0�e+���J�j,��ß��I����	���	����Iݟ<��)�h�h��K\|�0��B�������͟��Iɟ,������П���"o�"4J��"������!^4u��������l��ȟ\��ӟ�I˟��	/�qA�õrD4:�ҳ]M�)�Iٟ$��ԟ�����X������̟���!{�m�hT�|$��0�K;n����Ɵ�	���	<�Iӟ��	͟����;�v�
�m#�s��(�d����������\�	������4�?��b�V!����VP��� 2Z��#^�\��Cy���O��m�Cv���&��X�\ P��L�n�1Dn<}�i���'���/�9r잴Q�g�4 R}���Pi��7-�O4�R� ̪O����'���xR-�V��^X.��j����5@�Z����<I���7ڧqn����g��J����N��9r$Y�&�i��#�y"�����* {U	��3����&�j��
��M��'3�)�I,r�l]C7O|}����+OH*�ؐK�;-�8��0O��r�X��l�KO*��|���a�� b���f��$�5N���ϓ��6�d����s�m)�		�&%!僕m"���`��-%��Dx�\�������̓����:���;u��^^1�+�/�	�5l4p7�-(�c>aAW��,	���I�/����ƚ���1gĖ�sW&�'s����"~�yL���C�o�4�#�.��Γ7p��N"��ᦹEx��E��Q���Ym�0��7d�<_�Lp���?9ܴ�?�"ċw����'��쩷n�$����fح�D����]�k_h|IY�zjў�`y����6|��x�BXfv��6J̎������C8�J��P4��JB�K�=��Բ�Hc�z�[���	�Mϓ�ħ���.��@*q.V�ML�9��]�6�"�[��:"��'�2����7W�z)�f�$Hy~�"�M ⼰4�O�h�ҒU)R�8�'(�'x�6�Y�l��B/.�*(;��H�K6>�� �<���iӎ"<Q.O��D~�
�D��
�0t��N�]2 �剽K�@��%��m��ǿRQ��;R蛻	�8dI�O?����)B_c ┣ǈ� t��P4�Qؔ�*�'��]�d�����8zq��(Z��c흁1砅a���Ҧ��c?}�i��'�)S0oH>mK`�z�+S�dv����?O���M�r�i���E,d̒�'v���to��ZT��$g<���M�U�1�����W5��rF�x���{y��'�$�R4�6.�L���l˝����'�'�
6���1O�'�|��Ȣy��F���S �i�Odʓ�?�4�y����O�X��O[V���f������k��Jn����������Ĳ��9$$�O��׮��D#(�qW@�n	�U���OR�d�O2�D�O�	��0E��]��zٴ<��Jp�C���#�"��!����(��<Y��?�����4�ʓ<���C�~E��Dy�`{G���7m�)p�dW��$�����!=FNqJ��gy�kVO���j�x��U`g,K���'�r\��G�ĨD
j��ֶ��vh��l[����+m�|��E��b>]mz޽r�ML�{�=S� Y �Ez�A«�?!�4�y"T��	����� M� 4��>O�Mj!I؂v 0Y I�1?n���1O�-�၊��\k�;���<ͧ�?��f�nS ��Elr�!Z�b���O��d�O�Y���IV9�y��'=��q2� G!?�<�P��¬sh�'��Y��ݴW���O*�1X��r/�&f"8���#� &����?Y%�W4P��� ��3������"��v����?b�����6.�(�R5���?�˓���O?�I�*o�d���� ��A�"��r��牫�M�`�u�z�^#<�ӗK6:@H#�;S�͋��BdF�	ڦ���4�?�%̘�n�l���?��4���2�@�,��� E�$-(@���ܤ��4�B˓��'V��	��\�G	S�%J���!?�ֺi�(:�y��)��L¤ʥѫ�H�S"
"<�'���iD�)�	����a�Dy*��o,��H�˰Er�8FE�\�ɑa[0��,��)��E{��O�{tx`��LQf�jL��KgRW�d�'�'��6͑�U��\�T\���R�,�R�L��
��Db�#<�,ON�Dp�����I�dy��-�,^��$��:UĹ�nI'��ON�)%e�J�li	������3�5� �="��Զ*��9[&
�ZfQ�2OL��O��d�Oh���OD�?�ڑN��O����N�Q��	F��y�'R�}����7O2���O��OT3QI\�v9x8wːo˔�@�f�l�'&x6��Ʀ��ӊW��` pNi��mڛC��:���>��%�W�V�?."�¶�+��LY2�hO>�į<Y��/��.�2!R���!Y���*3/��<IO>��io&u��yB�O^���t���A��/Ř�"˟����`y��'1��<O�d�)�,�*����+m�(p�A��' E����}��JW��\��66�2h��DE�2Qr��I�HRIf��7j,�'�2Q�b>�~���J����{s$�;J͞�a �g���H�(m���l�<y.O6��4�.�r0�,KlJi2(V�}��EnǟP�F+5A�����d`�P;[�r�� g0?&i"Q��:w��nD����Bi̓�?�*O^�}b�@S�`f2I������r�f�;mE�����'���I}��צ��q@i� {l�Dӱ�W�6�pi�	ڦ͓���O����'a�����S��y�N��\"*�w���YJ�ZŨ5�y��x�� �%ĦU�ў����v�ۻT�|���4N78�v���'��'��6�LU1O�Q6���czn��T�٘r}m��'/���d�OD7m{�p�'���R�@_�L`�Q-P��V0��'� ��F*Xq���/���⟜L��_
Fb���	d�ظ��N�JKu�{q��$�O2��O&�$�O��������4L��rs��a�n�K�\�Z����?���i�Œ�'fr�xӦ�O�9��If�.id�!i E^)8���
�:O�0n��Me�iOBLR�N��y��'�LASĈ�-|M��j�E��0`���( Ϯ,1d��W��'����Iџ�	˟ �ɭ�$`�pc�xo���q�C�:�N�'�z7M���O���?�9O8h����/b"����퀵(�Ձ���gy�)g�NM1��n�8q&>Q��?�C�Dս���1����j�6�,A���J�5����0a�*)�&�;J>9-Of	sB&�J�����W���1eŢ��D�O��dV+jtfo�jyr,{�fH��8�$qX���y�f���G�W�s��O1oM�i>�@�O��l���M[��i\�z%�83X�c~�1MV�C�j�@F���y"�'�d�JE�Q"}V�I3�W�l��5F�1�j�↨E<7�*���R�y��'���'���'�R�)٠N�� ���U�)M�9p�k�.|�I��O�����1��w�����M{L>i0�7$���jW&�5vfB]1đ
��]�0��4[v���O0�y�v�L�yb�' f�GF�9�.� С��Y�f��݊�p@�h vў���ay��'�l�!��T!L{ϖ0xQ���'��'g�7���r1O�ʧ``�{�	��yJ^Q �������O���?	�4�yҜ���O'Z�w�
�"]ˤ���D�"8�!�՜s��5���9��$���["`ѤkdV�O��f�D�Hۆ�AeE��v�BTI�O��$�O��d�O1�&�'"�F�	���ReU���H� Ӄ>,���'���'ɧ�\�0��4�2�E&��n����3~�u�i��6�/o0��:OD��ҙ� ��r���sW�$���hc ԝ,�6Pb󏁕b;H�Γ��$�O"���Ov���Or��|R� �.f��x����c^Њ��A��OV"M��'9��O��d�'"�i���1��4B@�Χou�\�f#@(�4n�M���'��i>���?���g�PZ��	Qj�2r�+\�\�Hb�PBh�%#��q�n��&!l|%��'^��'�<Dbq��I�a��H��ϤY�4�'hB�'�"X�x�4z�A��?y�MZ�c�cֲ(`j�c���d�>Y��ig�7�C�D�'N)�WBɁ���ʴ(�+z��O.�pk /k �횑�,��'pU��
���O�z�n
"�
�"rrEr̘�D�O6�$�OP���O��}
��\���1�-_�O욄��nõa�Hh�����v�݇�y��',�7"�4������q��B��brLE�m�����Rٴ(���M��E��p��'��C�t�"�[EËvlb�ڗ���
�͘gf��d�(e�w��� �'g�Oƨ�� �f�tis��>]��@�O��o��Ojpc����@�Q<΍`t��x.�-�P�F(��џ�l��<yL|���?�u/����4Y!���&%�榙#"t�hkl~B�M�DuH𐓈X*ў8 ul
>B`�Xp�Er�-�g'�ß�'<�C��M����<�C,
+7XqHW�G���a���I?��4�O,ʓ�?iٴ�?��\u[ذ��	�y�����E0m�p�蓅M�<��
j���@w_���'�$a�AR�Нdgdɹ��+/"�$�7$u����\y�T�"~JGb1Pf @fL�,\l��C�^k̓7�ք�����Ц�%�P�W��s���Z1 �����CdR�<)/O6�ߦ��	��1K1����Ƀ|��`+���#M����+
H\�@�?���(��Sn�A\2">If+Ըgu��y3f�AN��wgZ�<6�á ��h�`P	:�p��#f��`!>"  �"����6pp$�Vc�'���S�*�6�B�A�t	n�"cd�9'��%�%◷F2=�֣G*�I�aMTd^���g��YQ���c�#�|��䚡jZ�]0T�L���BT�|�:�B.�����(FܕA��Q=)_h��(��P����٦��I���	�?u+3�V8G���;b&��g���1�a��ē�?��0ц,����?�����#c�֑��Z9.a�4)�4�l������)-�����4?������S7��� ���G=~�%��)�+��� ��i9��'s&I �'�b�'��v|�F �>4�`����^P����_ɦE�����Mk���?������x��'��u��I�h'��H��=]B�$Bd����O����O ��~���?��DV=RH0��DF0}�P����R��F�'���'�����e<�d�O������Bl�z�*yXD��� `��@%�lӺ�d�O��$�72���O��iʜ=�Li �oB�� �a�͈�.�� �n��b�dl�&��@h<�b�,�RE��KN�6�lPbiHK�� ���:�xRr�^	E���#"8.M����^�Q
�z��]�$�q'K�EO��yd���M�e�� 2:e�d97�U�}RB�;w�P�~��@��8�,�a�v�H�����#��g*�6J0W��,	C�¹��dц��h�R��O@���dң�mR��P\(X�D f�:- ��'BrJ�M��'
2E��u�,I��΀B���iCF}����ǧ�8h�ʰ2#b߱*m	�̒Ʀ�R�1ʓ`��	XTA *U4��������C�#Ղ]��IC��G�����o�!�M�#�e�'�|Q���?��i��o۲�"���Ā���13h[�K��ҟ@�Iɟ�F�/�F�,@ڧ.N%�n��b T>�xR�zӮ@2U�E-_���R6ni�
5j2��o�]y���+N�7-�O��Į|"E��?���Ͽ!� �� ʓ�Mp�H�����?���1���
t�r�y�$·8��P�S޷wj�dA.����5�<p����a�De�Vd��>AS�,��-PvB+6��a�H�+:nH�RJ<�N @V5�COA�\ 6b�T���&$��NdӜ�oZ����J`�T�L8���7�	� �X���h��?Yϓ'�ؕb%P��8� N�<,(��ɯ�HO���Oξ .R1��"x�Ъc������Iȟ��I�PX9sD/^ޟ��͟������1�+\Rڠ� eN;Kf�;DJ �R��⃀��?������ы�L>чΒH���
��[��ވ1�� m�����Iз)���QΔ�}&�p����	�H|����Z0�E2iK���Y4�U�)�3�DS7�1�g�/:�}�0�Ǯ{Y!�]��p�W�8J":��pN@3&M�ɩ�HO�#�$12���@�B��G��0��H�]�n #���#V!��d�O~���O�����?q���?�Ѩ�"t��ܪ���n�DXւ��&W�I�w�M>]���J�RJx��!c�B�\Fy2��8i��)&"�&�.y���O�=K�Sx�+B�ҝ������ `DyB` J�4�p-�\��A�����r�Cԛ�D{ӊ���<����$�<Q@���n� `V� '�d��F�R�<�"=8�v����ToF�Q�R���t��lӮ˓}��,6�i���'K��j@�&h�.�9D�%30�sq�'d�M��'W���>Q'l��Bb�<��Q�H���mɟp�j����ɷhM�@Y�ьKd>�I�n;ʓb�RE襭�-\(r�X֫\xd��ó.8$V~p�A���$=r`A�L����Q
�#
�.��O@���'Y�@!�ԵL4)Y�@�"g��ʰ�`�H��ן��?E�$&L�QXR��0��?u��M��x��s��|A�2H���S�8�i��g�Oʓ �,\H��iq��'��Ӕ����ɒc(Xe�5d�9'yJѡ�A��v���I���A�p:�(�t���sj�9�S��^>u�@K2F�@�D��Jzr�+}��h�)��������I��a�q�g�[d�����	?�"�4����M#��i�����9d�,qL�4������l-1O��d8<OX����W}��2�hP�Sʨ�'��#=�Ӏ����	�v
�;M��p���8�X����?��S�����Kǖ�?����?���7�N�(�$`:�?R�g��Z��D#	���ⲹi���s�
{1�*!zV)�y�_�s@E�� ��D�����7 q�2��L��K��ܺU1h� %Sc�ӠBʊtY�4��$�#��E�|Hb�"^+]T� ����O`���O��EE�Oq��ܟ�q�����{��~����AG�gq��D���<1E��`����v͕�B��ɐ�HO\�)�OPʓM� ��qdCQ���
u�J�t�b!��7Bz��h��?1��?Aa��B���O�瓖,�PQ�Cl�½��S`�paU$t5�d�U�� 	q��hVaC>'���;��.s/2jRE0c~!�v�֪ b���� ����K�1��ݺb�ٚ/�Hp�N��(OХ��cZwd��p��پ9@Uj�S�Y^��h��,o�̟D�'����Z�#@P����/ʸ�*R��<	!�I�;`�z�ׄx�� k�� %�1O��l�$�'K$\��f�|�$�O�lJ�I$��B�* ��yrM�O���I5�4���O�擄�TTs��9�DDq��T �"�R ��-�wbI�2�H8�2�3ơ)s���x-�t�ľ"����1�V )F��[G�]N`4��oȎ]��`!t��B�2!X�Ƀ7 h�HN�Ƀc���qOȱ��m�!kΜd�&C�	2v��jf �4���#��̍Ny0C�ɍ�M;�l�^�QR� D5�.�AI#��F625iQ�i�"�'��ӱj���ɌV����BFYL̝7�����I��p���p-��q�	Ē`�������k"MA�TG��ȁ�Z�	.�>w�JA�d���:M���X�AĴ/Թ�ě�
 uC����}���:4��.UKm걋�I�z�'��,j���?AJ~�L~� ��q5F͸)�N�4��Q��!����O��D݄-�N�r��'cP���&ax�%7ғ;��0Z%d� 3�ȅ�VΙ�\�|Hs�i�B�'�	���Tt�']"�'��w$vX���d��+��X4NND�hP�ʍ'��@5l��ꕎ��--J��1O�e�r/��X<�pf�d�@(S�/�X)�G�U���(�)��"&q���b'T���tK�=�$;pڳ�Z���ϟ�X�4�?I& [��?�}�'&I[�T�#'햾\�L��fӋ��{"�|2C_�rڒ�saA@ZW�J�.��$�Ϧ��4���|�����Ĕ�~1`� I�f��D`%��v�d��@�,=�6�$�Ot�d�O\�;�?�����E�Acf��˄z�dɲ�b	6v(�0�'$��d@7-�h����F� 2'��x�7@��3g�J��= ����������?A��E�AYf�1�͇w�B1��Ar�<YP�١0k�thv�V�W}�M*�)Lt�(��O)1d���9�	ӟ҃(��~�^�"`�3Z�H��Ў��H�	�f�����']��aZ���*i��l���O��h�㑃��D�w�É]ux�4�'I��ҕ8A6���aܬ[\�tц�$G&�BR(�g/�@��4T�
���q�')�c�E.�'�f�B!ʓt�(�0g����Ţ�'U�)��
\��`e��MΣ�nP
�'�x6M)4]����N'2q���
�N1OXq�lIϦ����O�L�''�U�r�ԡ8>�ċ�LP�wj�u���'��"��>���T>�u�]�anY18��XE�:k���O��H��)�8\4�@qg��"X*8x��`=_1��'�\p����ɧ�Ox8T3V�N�jܬ�s�(p���[�'�<a���%,X�@ԆZ.,|��
c����=VHL�S�Œ&�p2�7D��(fC��d�.u���L*~� 1"D��J���q?�I##.D-^)� �#D�P����c����d�)X�@#"D�t���ޚy�^yK'�.��=�E)-D���Ǉ:R�=�F����)+D�h�����\��Yhh��0���h_<!��ψp��(�ę5W������e�!򄌚*d�S�"4D�T�!���5�!��/%;*MCE&�nxP��p�!��O�F� YK��D�)�p�k���Z�!��6�ʒk�=X��J�n�a!��P���HiB�(��u�'�?	�!��2~�PQ���P��������f�!���m����+�D���_<Y!�[��P�@ˇ�,:��- �!�5pbj5Yw��\	~����F�!���q:ŧ_�E�*cC��$8�!�_�u5��H�܉7�p	4��r�!��Ωs����jK1_����T!�{�!�䌋�>�Ãj

���h��E2�!򄃂 ��p�vk�@oN-��E�*]�!�sC�	�̙QZبq %A�m!�D@���9��:Bz�X�c��!�d�S�~���E'2�����f�!��QB���eU�'H-�Si���!��Y�?�Raӄm�6&�K��B�!��C�^���梗�����M(v�!���F�<� )�![W$yQ"+�3)�!�$ &����DQ� CP}`QC!�!��C�nճ��g����Ä�H!�ė�w�@Qr�U�ijz�Y�L-!�DS0[�ȳ��YH�x����^�@D!�DD$qFiއ:����1C!�:zצ�)o��2 =���)4!���4@�MrS�Ɋ�Yåm��Q��3��� j�LpW�٪UqX��e�<���K*x��ǆ�K�D]1!*Io�'��YP�cȔ��]H"�zJ�CK�i1�N��`�3�!aV�0� �6Snꕓ$&{3�|n*C������f0�5����v�0�G+ݬ7��>�|��l�43ޕ᳎	�6���<� B���Ӛ0�z5
��E� }�-1K�!�܇�kVGԚ\�ԑ�b�̅E��|�b��&�D�ˉ�D9hf�]Zp5��hctӄj I@�_�|Pt8y��'��iap�Q1�:�	��^'"��Q.�
��$:FiŃ"��t���Ĕ�1�,?)��͋E��͚Ԋ�	��E1�-VI�'���2cBr�&M�̈́���5x�
��G�>1���W	Q��h�Kٲ!���zp��z�|�q�[�V;�,V�'.�R �F<<P,��W����Erh��=q�@&��<��O�}&4Wo�T�(A�a��e��	>��F8RDҒ�3QT���%��]��a�+Umy�2M5�	ނ��ԭ����L�!V�1�'�Za� J�!e��hO��%4ڗKW
��Hp��2pw����#v�|j�'��T�r���B�%`�%�'#VH��G�l~�DY����{/T\S��D�O��ӥ��~�V��d��+UWT�Z%I���q�`�T<El@�bG�)�A��'L&H�aT��o����c ON��L�,:�	2DC�+˜�B&�'It7MWAijpm�H$��ó�dXFy�	��?4X�ӥؠ��0ՆQ�z��ϓҘ'��0C�� �E	J,�)$q�TFtkZ��A�'@�|��J��y�=*�m�n׎�r��c�9��'Z��jl�fǮ��	�dZc��}K�) �?B�LK�&1))�%ȰΔ+^{��V�?����'���a J�VP����i��8�'���Sr�'�:7�B�UԼ��ܴOcv�I�ϕ-w,��%L	sJD|@�,�z�H�p���P�2�L�'TO�=���o�xxr�N�{VI�'U�@�}�������
)|���M�/�7�ى;z�Gy�X*r�d�B�G�E�2����Ta�� ϓ�~�S���uI�Ks�@�� �����7��t�0/{PQ��;ea��;���Y+��HH�@�xT�e��$�<����W�$���#�䅲�N��jʨI�"�1�	�	�c!��	a#�
U<�S��U2K��QL�����M�"�|�.��2w��I^���O��D��<�K��d���D���`6M���0�{Q��H5T�����CQ��t ØWكPK�=m\.m3�*O�Ų���?]^�5�AK��~�n8��'97͛�F�hH��'�-c� �a����Dy�nI��h�3G�gH�YԊůjh�U���~�꧟�l��8Z��b�ܥAa�0��E��QM�h���U�o�Q�\��ߔ�nZ�6Xu;$�_�^`��˙ �2�p��j`�堟��O����5W�y+c�[.x�V (�,Q)�$H'5m��R΄�pf�T)?�u.��*`
i�� �Iz�Ey�n�C���?q�s��а�Q�c��(�&7K���<(���F2P�lQ�*Y�MxZ���œ2Y�l%��a+�ـ�E]�0(��~�dH�q�Af����wk�O\�D�$]��bR�Y?7�1*��1>UQ���.B.Up�ŋ�ժ`#h C�	A	m"��%�I>��Q��[�����M���1�g0�Jܲ���.H �Ґ����Q�G]�n�Zi��+� E�ؐ��*�	s��|��z*��y���$�
	�t-�=�`�Z�ÆI�'kp�2������J�;����O�\�#ǈ;n���)�Õ�W�9�G�E̓�B	m��s�%�tex���49N��ݥ|�b�%c.{rf �Ek�~�n��C%��6�#o�4���c��8{����'�H�.��s�PTG�S�6i���tk�	�=�tl0��<t	��(J���7j@*{�X] d�pȧOj�=%?qP��7Ɋ8b����}.4U	w�A�|ᕤ��Q����JC�0���M���h��L�Rl���Mԅ�ڢ<i����u�Lb�c̞J���DD���9��5�G<b����׸}�<X���K�V��'v�l�s!��s-�C��.~!2��e�=�~���9�J�np��*Ӝ�5����5����*]�g�����a'{���UI�.��z"�H�:��q�c�<�3�Ʉ�	��\�q7"0����gc �3a�܊���"Ğ��4i֙"B��GyB.�o�ʘ���c0)a ��|dB��rV�<�A)}����R��X��1o|`x �:W���#��� �X���ɫ.�aEA�g���eO�N<���H�1��`�Ox	F��O���f�K�\\�'�))U>�K�"O�ݫ�O5,�90p���G;H}�P�i��ৎUG�.����@��EȖ�-d���lُ!�����r�,�5Lӕ�yb`�Bj�kS�Gi6�Ͳ���s�<IQ�)��񇥏�z�&A��[�	ƥ��.U����}�V �� �z���P K��qr*A|�<�IƐ! PQ�둓ow�jD�d;
5��	�H��I Cp�@�e!P3�n��W�@�wĶC�	,P����ٴ���"S̙�o�t7MG"=�0<���O���=�Uj.�ab�c�R�E���l؞L8F�H�z@��'�l�x�Ć���{�%�N��$��'Z�� QLD"8ҘP����?і���}�_�%��ic�TQ�π �h C�m��K��/�V��"O^�[v��#��a�l
lk\�Yv�U�%'X�5�?}��"�g}��'s2@I����Z�\��R����(Oh8��3�@H����|\��VV�����k/2ɪ�㗤aM��+fMk���'�p�]y�AF5_?$i�N+��qnZ.�BU��4yw��	d�~�`'D%!\A�sOI� ��C��'O��ڄ��=�X��÷v����R�Pa�fL0O_ڨ�+%)6`�sG4ʓ]{��õA �!����獧1Z��۱�Y<�����c�.�`G#5М�82ږ[9r�@p#?��ױaP��&�e���~�P��#S����d
Bv �RGA�$�4�p"�@\ؤ%3��($�C6���N�Nh8�LN�l8�H�'��L�B�,$����P��`ٌ��1R0��0�&ߧ�@��mu�y�`�f<j���~  �q�I�'I� P�egփF�(�R:����
>)i�Ye'[>ZV��p�4k剽,��i[a�Ӆ'�Э��GZ�"VB�<����G�2;eAԺ)ƹx�^�+�^����Q��S�Dx�%9�E�tM> �M_u	@��C�!�3�\eH��м;�	�%L��쎯IB�xD�UK�OH�'#D)��Z�ۀ��4��CG�D�O����i�j��"<WE�;,�%���~|L���D~"[�@�ȹ�ta�Z2ѱ'�̘22�6-)7ۮ6�ƣ�~R�O�p���$�?�gG��� ņK�6nG�'!؀@�+��Rm���Q)cv�z�(D;qzD�|�8d{�q�'� &!A#N�!0�RA�J�� �5��"A*��	>Qq��SC�'V�t	`-�+&/��@�3tm�ir`�X���G�Z���Ē�N�?arq�����ɗC�SE���U�W�|��5A�<�Q�;Q��
����-1D����M7j��4LAi��G\�(�Xt�OR�F��B�m�Dl01���F<��B��9?��(�h&Y���dj�x}a���2�� �'��*p�ىL&޹R"!G�=�X�Cݴ~E.5:���+w
�O�]hp.��nI˕n�VzPH�ӧ؃3t)3OϬٶ�R��^��&<:�I��rs��X�e�ȟ���b2�$�1�X�Hw�ʹ�?	7,F_�,�b�-7�*\٧�wyr����h)�tm��*\����G�(OpM�����!,�h�DG??ڑ��)��'J��"�)�Y�|"��n4z��݄m ^h` ��Y��:7�V�h�L��&ƨO�����3��nJ�r�"Q`b���n�Q�&#'3�&�)!#���'&<M�QF.��	�g��,up�xp�r��T��/�Ov���D?j6���
7\dj����P�$"�'n~�藬�5J�>����O"Hp��ߚ^���O"Ir��Ϻ	�]�@�ӏa8P� *�!?{��� gl`M)A��Kk��OM�N�v��ƴRD<����-��I�x!ueU��?9��&w����AǞ4�LCqyR�'�@y�h@MExB���=�(O�ų$�V0m�6��Vc$>��m@��N��'<J�ڂ���V��G�D�Ɉ	�-A􋞅(w3��ҩ$4���TI�2?�XF}rO�3m,�H�weޱ���ϔjNr!�k�5� �CU�;+8~L��P���Az�T�YN�$M�7,,�pөL�N��+ fD�o漩W$,wu����C�*����SHܨ����':2��Ŕ�W�@�c���o��$/�2�����wPj@�e�������:���Z-�?Q����:T�`)VL��۲
�p���	/1�PL�jմ޺,��סi���גxR�c��9�#�ڟf�(r��8��L� �k`��O� ����c���@�'v� �O*Q�����#�JM�.H�W��qB5#��@K�OZ��nN(��D�$OG�i�FU��f �T"bi�s��'rt���`D�-��G}"*��{'��z�w�dB+Џ-��Ri���xT�A6��G��^�®D[D�^���(S�::����� 7Ҡ]����	N<�ēU�R4�t�(p{bk	��}�aV���'�- �$���.��,"�,�5"��kgyՈ6~X�ڃ�@3X� ������`��}(5�� (����`�m�z�l��'Y���ď�1q�
�)�P9"m�M�,OĬ(��: e���3�C�-�0�e�I5�����Y��|@�S��Sgi>���x�<�G��N٠�ܡV�� dGN�pAƗ�qn�����=*e�D~r��+r>�ͻv�.�9��ȴwZ��g�*r����'��l�?E����� |���-��q��,A�xȉp�	/y�n ���I�Z���I(p��#dଚR�]�H� a�-��w���'=2��|�bZ�6�2 ��E�(��q�9x+z�0bl9-<a�Lֳ��I����*cF&���-Ad<9� ��o�ax���T�s`cǧobܛ �5��đ�]F��ugPW8�&n�;DQ����*@>TF|�5d�� ���q�;-��ɐu�B})��Q�i�m��KL6'�X[�&ķ"��y�@Ȅ�5�D>p%*�sA
Вf0x���ܬKAK�
7p���ߊTP�0�ȓ��h(@�$p�\0IƊuz"I��p����Q�Y�Nq�5XՆ��G�P�ȓ#:p@��aM�U�����E	A�
̄�ev�{����c�\�8'C�#bR��ȓ$�
�k���Bi�Ё�=S� e��S�? ��k�#0�uC�A�1>�<�"O��d�Krz�-�s�}�t�3"O�٩���+$�*����B����"O��t�ë=�4y;��ԝ2A��"O��!�n(��!��$0 ��"O�����V���U��P`��y��Ʀ*L�L���W�P}s�$��y�͟"mwY�@�&}@8Aq�JS��yB������O�!'vE�e*N��yr\�B��K ����`�$8r�'��!`�.^!%ܱ12��3k�~@�
�'B��D+U ���☎6�\�C�'���@����j��ѣa��D�A�'�hy12���Pe�c��atS�'�@@�H�3v��R�-s���0�' ����΄���!�BT0li�j�'��%�/Bh���b�Sj�x�'1>ܒf�@�q��R�Y� ��'��Q"�<�,�1�ΐ~�2$��'j$���
"�)� +"��uq�'z" ���FzMc�A�*Di�I�':�$7D/9n��f^?;���J�'f�*f�*l)��#�gכH���'� %���'D��XUE�^,`�'�j$��'��H��M�4�U�r�Y�'�P��LI4z
���aˆU�0l�'� `��d��]�N}�ӥ�;�����'_�	kQCH�&&���7�� �����'H (�+]�E��U��B�0;r��	�'�,�bצ[S�BM	F�ڵ"'J�'4��00�{����V�="��R
�'/�̛C�G6ߢ�1��&H,��'��}�R�ؤ@lZ�A����']Z����C�ia`aH֫LV%��'�d���N����{w��:Lm��'�н��%Y�q�����:wǤ�'��2b�kGZ`��+i���0	�'�2��ăE	!��B6!Z9��I`	�'�x���� �&-�*T�7���:	�'-��Ӭ	8|8�0E 3O��q�'�9*��:�6 ���Ǎ.�(���'|�{c���H�d$�"D��
�'D<i�6A��+ap��G¶^��
�'f��ƃ�1�Ũ�O]$	$�b
�'���	�ߖ��]��U8�< 	
�'t�r�lA4hY��� ���I��'�B�@�B6���g
��'�H��5�&��"�"hV����'��!w�_�76�
�bŊ[��r�'��m�ԯFRB^�)�CT��:�J�'%pA���D�zu�I�%�([�'���B\�0A´ ��)|��
�'>��(&�ן#����H$�N(	�'dNh@dNѢ'T��Ґ#��q�'?��*� &c }�0�fR8�
�'���ᏉN����G�[�.���'1J�r ŗ�^��l	�O���',�u� W�}�� c��r����'�N��f�,\��q@"�Ey� R�'#���JD�ٲu+���nN
���'<��3��;�(u
�c޼i�Z4�'�	b��S#Q� ���c�����'�%ad�_�}ݼ��k�8a}�D��'b��C�/%<�"J�$'������ �����p���j��<�U��"O�M�1&��J���#ri�9$N���"O6����6�\xb��o"�Pw"O``�-Ԃl�i��F_�J�;0"O�ѺG@�]y��(�IP����"O�<����t�p�t�ѽ?��P�"Ol�B+Q�L	�A��Q��"O(}���3tސ�u!�=�p��"O�Bv�	,�Yh�O	%4�ěs"O�e³����Q[�.;��2�'��O$ԛă��%Ȭ1'@�r��Ek#"O��E�-am�	H�l@A\T��"O��E�D�M#pmZ;*���"ONcFl_�3,ġ;2
��z(H+�"O�T�W��Ii>��/�c	$��&�'��*>�)I�M�)h�)@��r��ȓb�
���j&�"wh�M���ȓH<����
+�6	Г�Io��m��X�=�!$-+;��K0^�Ld<���m��5I�!�34����y-�Ɇ�J}Qh7,51�r1*̍C ���1�P��wr���Y�OC"���C�<!��־b�9!��&W+~·�]~�<)&�F��)���V R,�E �LQa�<i�IΪ�"�7���#�ppÔIP^�<餈ֺ|��
נrp[�l���5��ϸ�����,ȷ�jȬ�@��� ���8����ġ>�5c�('rd�gD�H��`�g�y�<9���~0�Mb�煆N�>P
�nt�<!�bƖHk�h�揜~nT"R͖r�<	%�������=�����F�<���Y-	02y��\�e�tt!h�<�w���W�6u�3��#t�M!uM�b�<Q�#Noj���L�1�j�e�]W�<��N^�*Z5��U�R�ub�B��%�"��a`8cVR	:�
�+~��B�I�&Kv͹�	�7!$-�7M��*M�B�_�l@��GS����8��B�I�B�4�GD��r����IPs�B䉭`*��bǭ��V\�|31��MP����e��Ӱ�_�.h$�k�$��@Q3��&D��p-�m�4`� �%�8���%D�P�$� �̱a��\?KF���s�0D�lS��H�2Zm�@c>9-�l9��.D�X�Dc�0l���҇�&A �<��i/D���g��.6X0�eˍ]�Z�1�1D�,z�%�u/$�9ƃ
X� ])�B;D���/R(�f��@'a�!�S�9D��A�W�����C��kS�� $�OJ�'�5�PiT'"�8�)�
F��"�'�>YYv�M�v	>y��'^�9+�|��'�ĘJ��}�Ph��N�#�\�'Lh$,��HQ�%�JT�R�'���r%\=1v�Q���%@�pU �'�$��E)y(�,!�!��2���'�MR� �dV�9�T卌r��\C�'��� Κ=Z*���П4�� ��'���"`A�}���$ND:&Z]2�'ސ�Eo���p�gcY5vht0!�'@�⤇��3-���	n�����'��}�r�H�� \CDJ�Nt��'/���!@בk ��G�ȷE��T��'rL��g�H�75$"w�S�)q���O �=E�d���="�"q��k�pM��E_(�y
� ��s�o;9n9�����9����"O�9��z��h�F]I�.�(�"O�D���O�� 4�ѣ	
H#�tZ�"OZxxЊX����"�#�.~�`��"O�PAB��TbP�Ԉ�7!h��&"O�� G	�7�P����2��P�E"O 隤�
z��#��6ob���"O<} &k��t�#HfD�x"O �+��K>\2Ľْ�]���U�t�'�O��z�)�N�y�(	.$�p��"O ��'v�x�P�\g���*��-�S��yB�	7!�A��17��i f�B$�yҍ�X�4!�a��c$A@���=�y�	���C���6aR �I�'�y򢌌Bάxs��o���P��ybJѷ �&@;톡��ӆg\��y��b���!�Iª&��q�u�E!�y�Eͨc���틦(�]���ͅ�y���"[��G��@�P�g*�y2��Q7j��A�����p΅��hO|��	�t�Q�ɒ71�U�T/:�!�D��9`�)�[�1v�`E�B�d!��^���L�⇕�jf((�K��!�$L<�Z�b��R8�PWk���!�dJ >�����E�x�(�� �h�!�dW�2�l9(`e���@��k�!�ۊ/��Ś��ǂP�vɻB�ۉ�!�dD#r�~!��_�`�zp+�!�E\��,Ac�^�5�d*�*��nT!�G)����m�3?����?U�!�d�
�:�C���X�P�DQ�t�!��P�"Zd�B�4�L�J�a��Q�!��Ny�d{@�O�p�I� 
:��� ����c�  Ȁ�ӈ���'
az��#%#�@��"�抝�2�Ё�y��«h�
���(��F��G�"�yR����r 
T�ű �"�q)��y2GY�T����W�����a�!�?�'��}�O�~�
�!�!�9�"����*�yBf[.i��H���SiVd����+�yoO�����M*6��LZ�$��yM,$��|��ʄ|�D���EϮ�y���*4�� �r!I$sg���ꊮ�y�@�tp���//rV���dm �y�(�0Zw��E��m��A���y��-�Tm�E�L�_�ޭ�ԥ���yR2)B�ȘgN�"iĨ��֐�yR-  ,�%���l��J�y�_?5�@�tk�"t���b�!�yR�ĉLt�J��_ vV�Yg�8�y"��΄��C��i�hs%%��yR�P��	���ã`bĈv�yrH�Ly��Q)Ʊ\m
HJ�FL�y2)8/`����FL�U7�`%��yҢR;%�$Y�⌵EMڡHBM���yr'S+.�^9�c��:s��4���y�A�tkh�Q4b�9t�̙���y� �V`t�Cu`�����S�K��yBD�,_@���S����Flı�y���9�}q�胾(�L��bLÄ�y�D�
s<��]$��]iRO��y�E.sN S���"��0��#��y�^�p��j <v8{! B��y"�/s\X�W�X f��ER��y
� X� e��**�⋾r�� �'"Ov�Qg�	��(0����9���J�"OV0���l+����K=6����U"OA�
�^!z��9E��`8�"O|�#�X�2 �8`T�إa�0�6"O 	��&��]��� BI�
�(8F"O�`�ҋ��m}(�J�����z5�D"Or�s���'l��2e\�,�ڦ"O��G�{A�A
�,t%['"O&�!� ��$��i̥��3�"O�y���<��b��Ý+�$4�"O�yPu�F� q���C3z�<���"O��[DF�\x�"H}�8Dʂ"O��HeE��+���b��� &�Aآ"O��1���n1z`o�#@	~p�"O�A�bCP�*!X�A�M�A�N�z1"O���� 4$"52�&^*@8�ӂ"O�s�Ô�f��5ɗI�{�e�!"O0���o683A��16��y�"O�\��h0)#�͇bA^m��"OT��p@<2eг@�4*�8`"O�<�DI:�X�B� 9p��i�"O����Oπ%���T��<i��8�"OEyfJ�e��4����-mT�}{�"OdZp��,�V%�Bo
����"O�=�gdF�k�4(��OU%:�,p"OtLs�* �Ld�AJ��f�\��"OZԹ ĵ [�)��(�Isg"Op5�τ�͠	�$�K<V�X�k�"O$���k�?nXH��뉤)�މH�"O@���lHo��+'��?�te�e*Oj}��i��M�v��&I>Z(�'k�H��!	�S	���
̺6`�U
�'��0��@����ԏ,�n�Z�'��@��/��9�����.2+l��'�V�*�$�*<��HSt�V&����'�6-3O�-�Y��K1�P!Y�'Ξ9�M�#=:(��BǕr~�,��'�R h�´xf�ђ���e��|�
�'�U�G��4+U�)IR�A�\Iճ�'�$�pK[� Ҽ0�Ҧ�/Xl���'��Hj� 
�0�27�L�U^����'��|��D��M����L�\�B�'���U0i���V��$Ii���'k&����r��y+��� lH���'���g�X	Z�ްK0HS$e�Y��'�p����pi3�b�{¹��'=01���(tL��B����k�'o��8wi��BM!�!J=
]"t`�'R�`BqFѼ@��E�lR9�� �'.�#��F�~X4T+���21A� Q�'b`� #�q87oŁ,����'� e�C,ޕM�)��**����
�'�P�j��bW�U㴯�,x�A
�'4��Cv��!�,�t�bA#�'�`���HͧU�~����A�d# \��'!�����O�)�nQ�Dl��Za8�b�'IhQcǒ�\34�YM`H�''r�C�*b�T�2n��Tr:��
�']p%�ƿIJ�=��m��w:y8
�'��]���Q�+������ȇc�`���'�,Ȩ���&��a�W�]�6��':�0��X(�����MۻK4�}x�'2�h�LJ��z��F#X�8���  DCg�@�0��5�GX��E g"O"h�D��\� �� lضw���"Oư�p�[�:����K^4kb���"OޙY4\�qoz)p҉��Xj��"O��X��͝/2����%�� �t"O�Ђ陼D!ظI��4M<��"O����Ĕ:{����&��4��\K"O�i2&СWæ	�.B�m>�)��"O ,#î��jv��{�B͎'
r���"OH	%h�:1���Z!]4�<�j�"ON�Jf�
Z�6A��F�C��w"OJ��e�c�L9 s�_�D��Q�U"O\���3��rQ��1y1@"Ob�wjH�Z����N�\I���*OV\�2�I(��{��PL��	�'��	�DA%%=�(�F �;� l��'�p3�cW;(�J|��Y.@����'�PT� #�* ���A�$���`	�'� 1�㌊w�� ������	�'=B�0%E�<],b� �C�;����'38\��NR<�.L3$�fD^��'Ҟ9�D ��u�e��c�m��'_i���I�d�8��R�ʤ^ඍ��'���z�Γ��*	2���]%j$
�'Ϯ�K�KS�~�d����ҝT�.���'�^�$J�qp]�$��G����'0���)	�N��%�smW8
h�'zp��m<#F��S֧C��:�'ܪ���bϤ@S��"�I�8��`#
�'LBTxW%ɰa�@�rR C
@|:�p
�'�Bbem��Y��"�"�@U��I�'�0�2M <�bŀN�D���'��{�&\�G��)��b�1�P=�	�'sD���iJ�XsDkδ7t=�	�'S)r�@̂``t��8���'�͡�I�)T�q��(�)|����'�v��u��H}�CK�"mQPZ�'���فf�;A��@Jd�x��8�
�')J��ƌ,� 1:r�G�A��'�ZV ��1p�U�I��ի��ߐ�yRH@VN��A�P�6(Uy�+�y�ώ�RL���@�a��Ń����yR��<�~5�q��(8���e��y��
h��z��,p���oS��y�bX�Zd��O�y�t�qį�y"g2$/�B��#d�6�ȠH�2�yr�$q���1-Z�n�����9�yM&vc�ȅ� �c�!#u*��y"��c4��BR'�f?����y"(�rv��g��^�Lq�ϯ�y�^�o�@��d�D�J ,S����y��֍A_:`�bd�Wڸ�P�I�9�y��@�S����rg��x� \��G[��yr�B!^3J���ejC<�2����y�-@:p�4u�E̗OHj�����y��ΝH��8���ρD�����y2�A ���@O��@�
��y�j�n��"�&6�j�x&��y2i�'
`����#B-��*͌�y���RC�ǯ2b�`�ץ�v'�A��v�f0��Q&T��3j�.5n�ȓC��I�v�i����cF��ƅ�ȓk�J�i��Q�/� �ec	�"p*���|T��+��P&~�D��L.q�̆�S�? ���𡏥^�pI)�@��t�W"Or���J�P��q���%my�Y��"OSRoW�7���@�	`����"On����n�Kҍ9�.ċ�IY��y�"�$ ���h��#?"�1rဝ�y2S�qw0�U��*�r1`T3�y�Po �d��cĂ9�f�h��Z��yk� ~`Qӷj���(��7n�7�y��+I���(J� �`'-��y"B�����$�0y˰��6e��yR��}$
���ۭs��\Ж&�yR�K:<�BQ86��j��!�vm��y�I��}��a�WƓ':����y�G �|ds�H��
����k��y��:1���� T4�����yB�T)ʴd�%�wڠ�2l� �y#�/
" ����}��,q'c�/�y�Q`$�j �D s�$TZ��_-�y�OP:� ���Ԛ`�%��`ً�y�����E8�(]�8�s����y�"V�.>�cB�@�t�I����y��6VH��R!U�w@t];Q	ۋ�y"��r��L��k&w��-��j��y.}D�(i�\�ؖ�I!�y�ŌR{`��6�ИP>bqB���3�yR�C-PN�irsE*@���j��J��y�P�A�йZ3k9g(�f�V��y�C�yD�	����9z�� ۘ�y�̅� m���㒆m��Đ��U��yfV�Y�<��C]�|�7!�y��U���"E��U&��@�I&�yB	̪o$�r�ާ}���iֈ���yU���ܲ@�~�f��K�>�y�F@�:�<m�"N�JC�E?�yr	�a�|,H$�;Q�"k��y�'T�EX��(��D6T ����ԏ�yW�����5���q!C$�y�@�<��E�E2R��h��y��E�, �1�����@STDkVgD��yr*N�)��yG@�9�U�&aW=�y��#a�$iؔa��0t�4��[��y��=F0Q�D-H5P�0I&���y��Ӻ�X��t�+�\�"�� ��y"-Ў6QЙ� ��x�x�Μ��y�FnJ`��l
 v:����>�y��J	e� �AӅ�}�
pJ�!��y�,T��-[V�$�x	���yb,C ��iN4)kb���y��.]AM��KU%��mBWf;�y�D��W�������d�� �����y���;B
"3���0a;����'�yҬ�%� 0���@a������S
�y� ��	���y�� �pՖ����y��ƁGj���ϔ5�e�a��yb+C�Ƞ��d�?�x���J[��y��[-K*�T��Ύ	��Z��à�y"l��k`dJE�L���9�͊$�y2�͢oX4�u�Yofp�#a�#�y'�o�0e� �aN�x5����y"� ������D�T�����%ӈ�yr��I���'Gr^I�J���y��kƴ�r�ƅ5������y�k�5jI+u���4�4���HG�y�D .Y,����%���U	��y
� ����D8�C�E�d��0�G"ONP`���_e�\P�cS�#S@	zd"ON���]�H[Z�x��ܘqb�0ˇ"O����}12�4X�(�x��"O0�s��ϋ^J�ʵƛll�Y�w"O$b�{�E�SG��	X�@c"O��k �8p*��Y�f�	o�8��"O
��ɕ�k�Ÿ�R 5➑�"O�;�\�l�ZQw���uҰd��"O�L�х�'��]��G�6Z�b�+"O�ͱ"� =i86�"�U>z0`��"O��bv��<&8�h��Ӣ`-�a�f"O������U45k��3�I�T"O��&KۀH���!^�PWhL;�"O�tRW��) !@:%��-u\�]q�"Ofh; ɛ6]���q��� I&0�"Oʅ;dA�k2zl�É��Y)^��"O*��W�Y�N���0D�S���K�"O8�	fMS<˖��u� �L�<���"O4,c�,*]�b8H��(@L���"OF`4�P6_�v�{Î2/��Y�"OZ})"�U��( 
E�
T�� F"OP�2K�2Q�ܻG/P;�JD��"O���[�j�P�@1vH�ɰ��ô�yR�4A��xآ�R!g�@�3e��yb�)2n0]Ð�R:t�(�E�I��y����K���� Z�qO�pxeF���y�� ;+��Ȃ!N�aո��D
��y�h��'[��AV�$)���1芌�y�H��
r�D,�/+���@B��y�M�� ke�=��ؒQ&���y�ʓ�oz���	�p���eW��yR�GsCN��wG[ü��2�B'�y���?l�i	S���٤�����yN�
��a���Yު��7�y�-Q����G����Z���y�JY���̺�	��M[4採�y�E@�l�tiB��]%3�p2�(C��yRŇ�-��K�mD|9B�f��y�+�T�$���L�yϾ���aǎ�y�-���ba�u�ʄ#iİ�yf�� cA�u`B8$�r!�4�H��y�i\)Z@��ÀX��������y�
�~)�f����Y��X��y�ƠWITE{i�6�X$G2�y�ȓWDl�&��B���� ��y����#���`�D�O�p��Y��y�oܡ� �+�L��N"|��� ��yb�X@	���@G"?U��bJ�yB.-`I`�F�[�9�zHc�a�=�y"�Ɍhq�`�/-s���Go@�y���:L����'�Ш!������y"��I�}���V8Ghܿ�y�l�(j�0�l�� �P5o_��yBD��9��DB� Ӡ��!�̋�yR�ȄJkj�P0�
rI�j6C���y���;��t�ceX8\ר,�U�4�y�菽#G�EYA�� ��j�)M	�y2"T�$8('�CJ dx#B��yR�DRm6}���U�h��qiǈGH�<�d́3c����ϙ�\#�U6�LN�<��ǜ:����O"��C�J�N�<�р��E'~��i��W���k�J�<9&o�7\xs� '*4*HSK�<� XP�@N+1��	Dm��u,^�
"O6�ypƝ�+�z܂�nԋ(����"O�dX���	R���y/�F�"d�B"O�������$���^�f�
�E"O��94�ҷIҀ0��-�D�@ȳ"O���G�ë��%��-�k�L��"O�QŊQ�N�zij^��eOJ�a!��-r���Y/ *����6LP�E!�u~*D�D6m�%`�̛�R�!�D�5nΜ�s�L*LkZ���
$�!��4+�H`q�L�2^YR��!��u[!�D�9Gc~0f�1*�� �hA�t�!�D�>XNˏku.A����!�dΈ?��p$�C� ^�����Y�.!�dڟJ!K�"�-B[~}��%��!�UT6zF��adF�=XC���"O� �7���|_<,�Ţ�=>B�qZ�"Oґ�&�����Q��z�B�"O
����^U��<;e ),mz4�g"O�x���L�aH(��/L�\�-{r"O<8:�M�2�*�aů�]���j�"OIs�T�uk��k���I�a�C"O���'Q m~}0��O�!<9�c"O�00㯞&w�z�̏�s<@x�"OJ�kDN�$X��U#æؘj�A�a"Onl�iD�!�d��GI-F����"O�}K��A�I-*��6�Jik�]Q�"Ox�9��Ӏ���S".Ѥw�Lq�"O�yy�K#� B�>I��j�Ck!�����L�W��|��i�/�%W!��@P��9�
�>���b�g�G;!�D�}�Jy�a����A�y�!��7>�xI�%	�J�Ph��E:%�!�VmV�qR�רQ�pi�3e��~�!�D��o����l�!+���k�K7\�!�F8!�>� ��ΆT�a�("�!򄍵7����c��&1��#7�!�ă�
�`��ԻD⵺ԩ�;g�!�D�>�4�hT��=v���Aj���!�03ݚ4�s/�'�,@Sv�C� _!�$	#W����B��,�v �i�I�!��;0�P���
T��!���$n�!�O�=��D��j.��d@�3g�!�d��_H��� �y�q�� }�!�J9�]y��|w֘р�\Y�!��Z
L%p��//vT�I�B�9Y!�䇘]����自TB)�޵4�!�$��*\d8G$�&��� �p!���JF]�"1G� y��͝�!�$
k�詁���@Y��d���	�!��.��I�&�m�0�����!�d�#njd�Q�B9(�Ҁq쓒!�5ond᠈Ĺ/dй���j`!�$��z�^1H�MJ�3�z=�q�ՓT[!���C��ᕎ�
�Z��S��">!��F� ��ФP�*��4�&']W-!��z�6a��0W��B��ת%�!��Vl@h�_X ��ANF%�!�A+yǖ��`F� L@4*�L�'!�dИB���Ҍ�&�u��k��y�!�DU�)��5��Ĉ �P��Í�w�!�� =|�P)�C˙&��캧,Ζ\�!�dV��
a��K�,��{�k�-!�$��V��k�b�=�\�1!�� �`j��S*~���EL��#AL-à"O��YѤ�P��h)qd�F���T"O��� �;[��P
ѐ�� 8�"OTU�"F�Js���ɮ��"O��c���zVq�.ޭQl8H6"O4D���#M�0Aː;�L9r�"O�ճR�^&v�9!L��]�|�g"OX���!��/�⁺�ȑ0w~��"O�m(�� 0k�~x���N���"OF)�MR� ��1�f��Ӧ��*O�(���Àkʴ!�c�a�J)C�'V]pr�Ni����@�^%W�~\��'s��3@Ǜ�q�`���U[>��'��)�A�n�f�0���8/�h	�'�0�J�@ 
�ɻ�j�)��z�'�x�&��2�����R��8p��'6V5��aԊ�t%���S@�"�'6�ٰ��$�a!wi8=d���'n�Á���S���k���:	�E)�'wvl1���lc��P�.�:�@�'���iΟI��X)�ȅ�P���������g�
�
��E�ʌGN���ȓy`ɐ�Bٸz` D	�^�W#�L�ȓw֦��r�:
�0�0���	I�ȱ�ȓ?8�q� +��p�lŁq��t�ȓ�8}(3�����M� p�d`��=���M�,��s�nE8>n�d��(��q�C��g���E��`����ȓ4�j�� �ڸ�dnW�R��t=`�k5��7ư �'-��p��ND�ĉ���'g�����/����M��H�W
��a���͌+	�	��WȈ9����;)����'t~L��>���c�=V��+Q&�<=)�� ]�uS��(��Q��D^<�ȓ �qP(�#,�)��EN�;|l��6�[uB�h]�,p$�c/�u�ȓ��:�%P�M��"D8I �y��;�ኀ�g� ̡ �H�ܩ�ȓ)��e�נ)�(p���(Nr܄�g�P���@:2i���u~rՄȓP�C��ڤ$�P���V�vTɄȓ)�X�m��,��&C�=X:�ȓ-�����+Sr� i�%��R�L�ȓ^�ڭ�1�PnDxз)�:(	�(�ȓ�������_��ɳ�%��[�����G���9�c,�J�c�i����}�ȓ1��hP��Ky��Tb�WS��F'�)�&F��n���˱r���ȓ�y���Α7��(�V�M�4Jń�;�<Z���Εbы4L�ȓJ��@1�`�C�����ޅb-j��{��b��	E�
��%���l��ȓ2����@ǱL%� j��[=7�����6b08����}�ܱ��<B������d`��� oV!R'�ܸ�1�ȓ}0ST����@"�(7
�����#�Ȑ���U�U��m�-�3�����x���!"��>�6�G�vꄇȓ ����ᑧL�P�wNPfr⨇���Q�	Ւ_)&`kC�_�������D`��5�3b��ȓdY<kQc��85N���i����N���
M�"�I�3�G
&b@���S�? $i귦��V.��ԃ��:  �g"O��R�
\�9�U�J�I)��[�"O�2���R�ļ���ֹ8 D��"O(�i�?�q� -C�W1��S"Op<c�"�K��M�w���"����"O����m�"�A¤��2芁`"O@r%�#T��1��[D!Ru"O|�+RfL+o�e
�Ӭ%j��"O�S��
�qY�	B��.E6��G"OFh9CC��Q����s��,G��A�"O�b��^8Aa���C��w²HR"O�,����j��$�6���Ё"O~��ŉK'E-
���T
,`��"O�diDN���G�J �Ԃ�"O��Q��zpa�e&L�]�vX��"O����o�
)��Ӳ��/"��i"O�$3����[(��ZV$�"8pU3�"Ol�C��0F��]!�"C Nȴ�Q"O(x[�m8H�&c}�x�ča�<��Vq<�%��G
M�<�4a�<���^Z���TE�~j萁��S�<���̵-V5	7/�s�,a��M�<�a1�\)�2�u�9Vb�T�<a�o׌�,AZ�&�>�E㧈K�<�G'K4D�,AC���a��㖥�~�<Y���\;r����-8�z��{�<Y֤�#W�\����8���z�<�R`��Q'*<
�˚B��lZeL�t�<q�Ɍ�A�d����&8l"��Vq�<� ��2l̘ ��,It����j�<9R#^Q���%@��RX��eC[p�<i��"C�����U&
�Z�cv*Mi�<сe�$txܽ��m!t�¡���GM�<鑪�T�S��QUb����L�<a��N�"]��IW��E��I�d�<�c�I�E��Tٗr1~�Z�^�<��΀�[(�����WT�U�FG�a�<Qs䈧4k���Go�e.AR�N�]�<�5�NB�B�Z�@s�����Hs�<Av`�=`��h�>'R�C�D�<A�̕�[�dP���H
�z��E�<��`��hӤћ��aՐ���NEG�<1�"��
�<9�H�خ	[��YA�<1�ސW���[�I����v�^h�<��لjܜ��J�#���!t�b�<q��]�2�q Oڇ-�&a��`�<��$S�*B��yǡPO�ʱK��a�<����5��j�/\�˓�_�<��F�>(��8I4z���SDM�^�<����'��N�6Bd����A[�<1���l��1�D1"�R�k@o�W�<	���Ka$(�#��vB��PCQ]�<�V�l<�k0���I�HT�c`�^�<��o�-���&��*; \��i	A�<�`�U�|�6�X�
��w$p����T�<"�� �I6/]#{+����*DN�<��K�&��2�F��@�'p�<�!��?�X�Y�菗nym�-Kn�<��![.%�f��F��JFhD�q��r�<3�,V��
%�քZp����
H�<��b
#H�lzW&�M��C��C�<��"��uP�I���ړ7��4��aFg�<I 	�(o�X�3M��	�n��-D�IA�Y�3Ϥi�H�nJLuQI&D�� �Lb��gک�&9/t�!"O�X��wft	��h *z2!"O�4[qC�O�)y'-Y$A�$"O `�Lc>𳅆�2Y�}�D"O<�#�+_Dm�ǅ]��NI�F"O�D&�P8	<$��c�&_|�<8�"O�����?1T����@�<?m�B�"O��Q/�"��� �Q�y;�"Ov9��B(0<�֍S�S��`"Oh�AրK�N�2���0IB�I�"Ob�{B�U:���0��"M�2�u"O����QM.4���(����`"O~��,`�.�%�E>k(�b�"Ox���b
�90,��(Q_��c�"O�d	bI_+,�l���;_e
l�#"OT8��V�t�B�c�F�N�`���"O1i�h�54�$Բ��߉Yy��2"O�-��� *l�����. ^0l�&"O��a����x���W��3f"O8�� /D�5�1�R)hqnp0@"O��s�S%Ƒ8Ca�9ol8)"Of	��(��=�s7�CaH<�"O�����б.���/�+J4I�!"O����F�٘1S���Rc��{�"ONE�B��4�&��"�qK��! "O6E�`#@�tf$����Dv.���"O���1��F]��X�$�2K����"O,��s�ٳs���d@�#=��0"OR!a1��(��T�D�=���"O�!�
E�Z�0h;B�×(�&HiE"OB��h�� ��S�
�7�V9q"O􈔤��<~�=z���.0����d"OJ!���E4 ��$A�AF.>�^��&"Oڐ���fp<�E���&�B}��"O�H���>�Q;�e>�P4�"O�U����%0Xp 2/"��[�"O�ӂ6��i��Awg,�Z�"O^�!bΗ�4W���A�D�Uȵ"O�0#G�۫:�	;�	 튡�"OLHb�̚t�"��2N�#�*)z�"O, ѣ�t��H�vl��Z�"�q�"O���BO�=T��Q��]�<hQ"OSt@�T��0��'+�Zy!�"O�bS�h�JA�2�^�}����"O�d8&J�'B9<q�
ɇ4�:`"Ob��\�	ކz"�<E�|Q�S"O�ŉ3���\�x��һ��I1"O~�PC�8Ar�(&��+��eP"O�0xGf!H�(�O�%R��z�"O �'FQ����s��;��dK%"OXA��/9?߸Y:��<�P"O�2bӠ$1�Ѫٿ<�-�@"O��2�d��1���3�� "O*5	�V�IƔ ��%�2H�"O�h���]�x8���k��0r"O�#�l��^�|�zG�<a�f���"Odq�d#Eؼ��W�e)�t)�"Or8c���(����1���t8a�"O�rB�H�I��ȱG��J}44��"Op`�2���'<i+���:Y�Pᨶ"O��)w�x-����'��� "O���#d�<&h,-���E�b�AA"O�,�&$�-AL~�ɡ��2�
�q3"OH�� 2�(B�fՈL|j�`A"O� ��ÔE�.r�����%%L�x�q"O����7"��3feoEP�z��'k���R�D�9��/��0v�y�=D���j�(�<颁 (,�Z��h;D�2��[�5�&}��-B�}�:@K� :D�Lڷ�!%È4ȁ�\ t+x�@�<D��
�K��3��M��J\CE4C�;D����`��;���a�Xc2ȕAa$8D�0
r+�)50�,H�h�+h�൒�%7D�|����1���IES�*�ӱ�!�	l�'��	= �t P�Oϻu�4�@�*�O��B�Ɂwah�S�Mϥ���4$�*_�B�ɬ$�$M��k�3��a�2m�.5��B�	��D��.�1+�A��/
�_Y�B�ɤ�X���$�h]��7ȦB�I�EE.� �G�^c���E��h0�B�I"1�R�p!�m^r�����nB��,,�n�0u��4�P�H�#c6B�	��]I"M�R">�'�u��C�I�8*s.��w�p�����_e�C�Ƀ>zp)	��9k��QCŜ�\bhB䉤C��<���\��Ƨ� �B�I��D�@�lZ2L|e���=]�HB�ɑ%���v�˥! j�PGG:0CZB䉞Qu8�3�+@�R�:��4�#r�XB�I?uz�u�������ev�B䉘Vj]9� P a�9���_�D�B䉉��R�?\x��`�L?.C�ɦ��'
?Q�8��V&VB�I�$n���Rdˬ'���2�� 
����<I�'��p @ǂ�#�xI��@�B��X���x���3c�Q�`^�^(y�C_��y��ke�����*D�>1�tj�5�yB��N�eq`�Ȕ6��#̈�y�`��6�v����Z>H�L{��5�y�iӊReY�$��8�hB�����y"�V8c�ZPX�I��.E:h�$�yB&�PY,�H�@
	�H��c[�y��ҝM��hP���p�J�H�"��y2b��-H��+�-Ѱ~��ԑ��y��ʙ'j��b��طK�h\�@)��y���4k~ 	�A�4hz10��1�y�M��ua@�#��
0(�]���@4�y��&*0���ᩅ)!IƠ�9��=1(O��I�r���r���XK�N�?a�C�?� �y��^��U�*֋�����'�HՒ�N(5f��"�QC�1�':T|�fM)&Wt僴ĎY̌�A�'`�Hү͌uڀ1iC��eu8��'�V�A�I˚c�����D�S���	�'l|µCɅ.@qCf��4���	�'J&�rgÓx|(qgG*)��a[	�'H�պiR�y� ��Hҵ��@�'D�t��o�<�����̢���'>�-pg��}d�@�ˈ��m��'��9f,�tE��"�2$�z�'P�� ��S�Q*F��	��Y��'��m�2�N�g�H ¥��Tg���',���x��)�/!<��H���xR�ҁdpT�Ԡ?̠��[��y��������5�	b�.Ѻ�y�jR�wӌ��' �xoP`��� ��y�@�Oe���������y"ÛW��e���0��ò�'�y
� ��K"�L(���E<n��܊�'j�D�AX��LZ�`S�i�6!�$�!B�T,�ф�	1C>t��J2Y!�d�Rc���2Cʘ=�"DV�;!�$�(8|�$e��&�ޜ��ԛF�!�Č�w9��!��ڮ0�zH��ߟI|!�$@�D��ԑ���7�P�;���_w!�
�(���u��8*���Z��
@h!���shf�귈��)꼱����8!���
-0�Y,� \�bf��2�!�D߅ ;�dp�ctV\QSP��!���D���9$aD$rE�	ڳ�[��!� |�(�`6C�u���;�/ƙp�!�D�;f��x�K11�h@�-J�x�!�d����oG����z�lB(=!�ƜN��Xh`뙿Gx��r�
:�O����2?UZ9H	��Yې�$Zu!�DG�/�Xi�a�#چX��N�:Q!�dW�J<�5�E�].onB!��,l7!�؟-`�\cQ)J�mba�DGMB!�$yw�5��I��`�	����!򤟆N?�,� �.��U�P�N�!�R�?��U�A3�Ne9%`�4�!�A$B(�4��@ĭ��9�4h�!�$S���$+�͚�~�>i$�@�!�'�X+@�p-���ރ/�!�D�C �@
DLz�� ���*/k!��13�d��:>ܹ&o/}O!�D�H8%Z���2xg(�%�ʜ@!�D��/�h�&	�t`Fi��
I"s?!�Dǲ}�mh$��o�� 	;]&!��Y�Q����J�[WŠ���J !��F�24Z�p�`ڽ6vx��J^�q!�D޴�]��K7Ig��D@5!򄁡KP`���R�Z�P)�A��!�K���s�"H�g�P���
ԶM!�D"5�����Р">����¬v8!�D��!K� ����%s�հ�מt$!���vi�X����E�Zq!�dзo���� �Z@f<
��R�!�D�S�J���h�R�u�$>!��;�~�Є-S7��L�b[�\�!�䛩��C�̓fFkQ'�D�!�dīO��M��J���䆚�o�!�D��2����ٰ]x4�q%�%P�!��� ���)��']A���#$ӡN�!�D�9{~�3�D�qh\�'A�&s�!�ǇK�~$��@;o�8��D`���!򄋒8��$A�(Q�u(dU8�.з"�!�$��(lx<��M�.t��01\H�!�D���)(�	��=T�PK���$Hr!���&e��)��݃hOܹ�$��U!�d�/_qGY�sX���	�n�!��7U�*İ�n��A��Q:&�>�!�D�r>�@�!C��>��9�T&��p�!�$�!�l[� עT�Ig��B!�d[z�e��دP{���5蛫, !��Φ!�&�ӅAt�(�5B1;�!��ɾl�����$߱_���@���!��^Ŝ��Wa��{��]q�C�*�!��<H��}adO4Q2}�d��( �!�>)��I�'�S/+�>�0�Ƚs�!�$�:���P�ŏ�4C�$z��C�/�!�W6c�A	��J\&��C� ġcL!�� (b%G��� �.��j Ńe"Or]Af�@�i
h�`T�
�/��@B"O�9�bA�i�" iq�I�z��"On$A���->��H�֏�"����"O��e*�$p��0 NK�|�bd"O�y�c�&Qz���d��19�"O����O������)��G�
�:0"O��j�������L6G�25��"OX����'�셲E�E��lS$"O�	�T@/vn�W����4Bw"Op@p��k��C�aA�K2�1��"OP�e�;F�d���o:�R�!�DPu�N�B �:I���U���!�G�9�lD�s,�'k���V�Y*�!�ĕ/vH��eM B�"X2���:^!���8#���1�F�� $���jU!��oP@�F�[�kpd@���9d�!��*E��\�׀idh��q���;!�DE,u 0S�J�Ml���s*�(H3!��[
�
�[��N&=�5*]�!�$��j
�jN9a�by���4!�D�B�T��Bʰ)�FW��!�d���$��E�8����}!��84K$�q�*�	�&���Gc!��ݙ*�<�;ńʯCϤ�3-���!�́F9|�bB���'ɊqX�A�CF!�䜥�*�C��U��ukӀ�p�!��d?��E�Z�z��� @�"r!��S��P����5T���2 �"�!�$Y32gj0����MS@$��;�!�D��@��!��h���-پ$�!�B�����zs���;��C�	M��	����9\�
ŭ �4~C�	�e�X8�a�������� 4S�B��jh���'#ů����Ă�4tB�Ɍ'x(p��/p�x&���HB�I1�X��Q�Ωq9���g֗t,�C�I���Ă�����I�T�*�B�	;k��H��B*� C�6ϪC䉾���ق`�mæ��FHЭ.M4B�	��:ᑲH��JfڌrG���DC�	>f���^�bB�(��_GC�ɱ!�ư���W+;��A���r`�B䉺=V�XG��3���@�-Z�B�Ɋ~A��WB̿����A6d�nB�I�@��#e��P������t� C䉞 q:��V>)��3��@��B䉇,l��c#�&GlhU���J���B�I�a!��RG!H�-����$	� �*B�	)L�bSG
�r+�M��Ɛ�P��C䉢[��x�Ц�<,*�=Kׄ�_�B�ɠI�ʗ�ּ �zQk �߸n�|B�I�X���C�@�1�N������F�pB��_j�y��K��<�Yr��g�PB�I�b���k(����\�lB�	;9��ɕ�Y�H�ҡ
�T4JB�	�5�̡��]T��kV��T�B�	5~��<�'���{=d$���R7d��C�I���zh�-=\�� �5&�C�	�y�%`T�	Vo�%*��˝dn�C�	<f�ı�DH�lʉ;QDɿ#KB�9�tŊ��߬}��p���ZF�C�ɠ�V�A��H؝�B@�b�2B�I�8l�5��7p���b�nŐX@C�)� ̠8�c3+H�,�U��$Ҍ*c"O���bD�\�̝ĊO<��
�"O�����,D5�{e�?�*9��"OZ�b�I�k��(a��<tɦq�"OXи�F*\���l�{�v�y�"O 0�υ!ڈyà�!�$i�"O�	�t�[ W�(۷�0��mj"O�@s�L+]&�1kV�նm��i0�"OХ��-�	��lje�D)	���C"O�4	��p �'O�Z�D�v"O�A03�]'��L��v��E�w"O�}��l8�iE-t�98"O
�J�HF/��$�(k��t"O�U�(\�ܴA�-��$6xrE"OU"��O�w��A��mJ� 7��*b"O�h��N�m�P9��J�/3�H��"O�8�B�)a���It�RP 郡"Ol�I�#Af������$[�AU"O��� &D��D�q*/q:�+4"O�����X7�;�W���F"O�P�B@��u~��zǁO�cV|[�"OP8���ǓU2��f��'.�R�R1"O�h��
�jc!�?V��$�"O��B��M���bbT�u���#�"OThأV�e�DM��ҏ;��� "O������6�:ucZ9Q0��`"Ot`#�O-I�B0�d��?3j96"Or�p��kQFI1���W�*��"On���d	!�> ��1�"O��(�̌�t���G	�H]�E"O65i�Z�DE�K���6a�Ѵ"O��w�޴m&m`J��`E�"O��#��4�BHz$g��>�\4ч"O p���ѦJ����pf�&*��C"O>P�پ{�Ld�ԪG�f�2�"O.�R�ؠ/l���G�vI��"Od y2ˁ�rejV�ٷf�^���"O,���R%g�Q�t&�A��'��� g�O�fu�p���$�	�'��`j!
D� �Tii�LL	6 U��')�	��J�%;�x�'M��{t�!9�'�:���I)"��8���wM�X�'�`Q���0�H�ZR��u�,A��'4@��(��@���3v��2�'��H�bb�*kc|��W�=ET�8�'�`�>g+.�z6N�5[���
�'Yj%+EjͲu��D�0�Ս3��uJ�'Z�:G�C�}Kt����C��!�ȓ!�P�s��k��8@�%T��܇�X�̄�#ȓ	�h�g��� ���5K\]Re�<!,��ZҪ3.m��.�@���
���
����ȓ<�0}I�%h��X"p�Ӗ��(�ȓY>�p�nC3gBv�:FL�w����z���kQ���"�V��$F楄�.0vx* /ҏrZ�q���E ��ȓ}֠��3���x޶H�� LxP��sǤx�Ƭ�#:����Ш�.BA�<��):�� K�"`ެ��GB�<�A/	�P	p�S�=��Q�S~�<�4k�* (�t�B��]�!��|�<�2��9���caHN4)|LPf��N�<95��?!�.l�V/D����EI�<��jI.u�z��5g2sm�9+�HK^�<� J\�wo��~uaP�NԔD�2y"OV�hJ^4V�����
,��"Or9���ՈK�Tz��۴2o�	�"O��`fB#:��B�,L
!^z�S�"O�-���+5�`l9!J6B@��X"O^e��]3�%yb�Q�U��H�"O���0/�bl���֣�E"O�]YU劚Ò���<s$��w"O��3d%K7	��+�C��($"ђe"Ot5�3i9Y�4;��Ҍ8�i�#"OX��H�D�X)�5jC�}yХ�F"O%P��Bb�T AO��bm��3�"O�!�1E�y�ZI��'��Wc2"O�q�0��`�xР`H�1ax� �"O�� E	S��1��t����"OrP�t�ZVɊa����Tѣ%"O,j�CM* c�X������"S"O��"��=���q�A�~��MB"O5k� x>5�W��:�V존"O����f;�Z͈y3���"O���eo�:uhB΍3*'n� "O�T{�^>9�,4k�K�'"^e��"OVɺtLE>pCX�4)� �e"O�Ib_�R�n�a��#��E"O	�CdN�"��\��/n3��"Of8a�m� E�P�bh�!�\�"O$!8���$wT��'E�<i��W"Of���k��fJ
��E %ļy�"ON�q#GPn��i(�d����x"Ot	�w�ўM�
ِ�� �~p�jP"O�]�k�7G�rIQ#D�8W�Ų�"O&T[aB��I���;�i�%p8>�Bq"O��
�%��D�2JP��"O��+����~Od%3��M�> htA"O��ǆŚH=�-�� �5H�s�"O��b$Ym�:��Ca�+��!�"O�}�'�.^��0k4�$&��!"O��s5IX6s%�� �?ljH�3"OH��$V�M\�R2/D�
�&]�R"O(36	�?nKZ�qu+Z!:�ȓv�*��q Ya���@6D@��J���*���#� �*��� W����ȓ!0��#N��G�L5�$C��/D��p��](V�e�!'�A�pl#D���c��,j�SD�H��=��/4D�t[��"v/&������w��њ�4D��
&�H�Z��t������r��0D�dr�޽U���ivmsxac!g+D����.�&G�0�*WG�1/rT�i�i)D� p!"U:3c�h��a..��p�%D�4Qsn��d�(p��/ЙC霼���$D��Ga�Caޡ�J�Db�q�G/D���D� �"�p��˗ah}��M,D�h1BB�:sl�2�̖��@��)D��� f̄�"S�u+ڸƥ*D�X���'wx(���Ͽ �$a�3D��`/H5hB�l�7Ǆyɱ/D�������=�^�a�Lʋ�XɃ�7D���DyôX��`�=BBp�w�4D��hP#�5�zY!�0UX4⑆1D��K��H�_He:�@�>+BRb�/D��C�͝>\S!ED�B;�ip'2D�������E�Ӌ8X��u��%D��#$ͩo��jO�A*��Yd�%D�� J�;� �d�ƍC��A�
ي"O
1jB�ʶo��p� S9�R	�"O� � $��ɠ�ϑQ��,Pa"Oڸ넇�d����C��,�4���"O̽���)p��2�aS3S�p)�'"O�8��j¬v"2��OG�L��!r6"O�u�f�[���6�liy'"O8�g��>A�q0�kH�2��q�"O ��b��a/�|���3Vq8���"O� "�OD N�	'�A;gb��"O�(H���R��
��\	�Fё�"ODxP�	2X�ypF)`���R"O"��N�x� ��f�&�Z�X�"O��hӶ�4� �z�H��"O��`���M���� �A �`��"O�]�DN�G*cC-R�zț�"Ob�G��xv9��˙���R"OL��С�E��T�֩>~�2�"Oέ		@tjddI�Q��Xk�"O|x�%V@
T		����"OL���M!�j��ǘ;o�ճe"O:aaa��9!YDM�$�R�S���90"O"h8@EW:)�r-2�L�|HR�"O�Y��I%(�2�`�#�D�9�"Oh�ZV L4tb��\}���ju"O�<�fC�n����S�P��ꕑ"O�����D�"Ծ��C����!"Ot`�*S�~�J�c�#9����"O�i(���Q�gc������"Odx�d���ʩk��)���9V"O4���Y�T�y��Ưs�D��"O��࡞�190��#H^R��� "O�)2X0|����@��sB�=��"O�h	$�O���E��""[d��"O&hɒN��$�����[H2��"O��#�}�Vl�Q�֙34�`Z"O�U�
�/I%��D)��V򅂓"O��b+6S�^X���u���s"O2��cؘ��঩۽}��TAT"O��*��� n�pda@��y��A�e"O�a�oG�V��8�U<q�f ڤ"O���g�Kz�a⤎�aҺ5ۤ"O��8S▶1��Pk!m��S�T�g"O��C7lQ�ܸ�yցf�*-�V"OB�3",K�L�ņ�b�$�)�"O.|��߯E��DЅϲ�Y�
O�6��t`����2$�VAáa�=�!�� %�\�����f���+�'V`2Op0�e��@���E<\�X�"O,a�%��+h�8�,��uLBd�#"O��d��G��YSqM�<"O��:e�^�q)��3��������1Ӓ�A3DvCva��u����F�Z��%�[*U|d�2��+ ����*�4iσӒ�RR��>P�$)��}^lіƂ�a��]*��2m�:���u���E�+z֔�F2?Slņ�k� 1H��Q��)�C�Y��$����}��ԙ:0�i4%�)M��I��m}t��`Y� 	$TA��h�9�ȓWa�(��aئ�.�
��V?9Y�!�ȓ��������d�^�{�HFV�U�ȓ&iX}�L^�TƼ�+�K���ȓy���g�ۗW��t��|.T��S�? ������6*�����M�z���"Or	�,�0:�����׉^�Ԛ�"O��j�M%�iq���[��4��"O$P�6ćt"d�T�D#3*^%��"O@���3C´��E$�\�y�"Oİ �E��xxQ�/r��$"O,q'�W�ڨ���J
*a�"O��R��W��N��P H����"OB�c`�ζAXd{2B:�"��"O���P�gh8�*V4�̥P�"O`�z7�R6Rj���@�(k�X��"O���oñT�T��`�0 ����"O:�sE�5I\�3.ޔ'Ҫ�"*O��"�Z9%o�4A�L.cL$
�'�����),d��`�o�Z���#�')br�Ջ7��Q�]�F�����'o��b�� r@Y�-�E��
�'�:Is�� �JDr����A��0H�'�P���f�0���`�]�4ڶ��'�8��(=,� �IA`uVQj�'�P�#�C���=�AK�/�:�'�j-R�ʅ�X�|��`��x�j�2�'ʦDj��~)r�Pw�F�jNFݙ�'�,��L��+��kݢHt `�'�ĸxaa�j@�<*��UoL���'qL�Y�:`!�䊥��!uJ���'�u[g���*U>�J%آsbd�
�'r�	��U)�
ݚ4Ŝ.X錘�	�'�~��w��PG��bcM2x\r�z�'�,b`-0Lۦ�B �mX�X�'\�9��O�?B�e�N�1>�i
�'�~ԉ�hI<f��8�b*A�.��1k
�'u21a%cА>�����i�Q����
�'�K�yU��b��1z2��Q�<)7ϙ�R PBE�PWH���(�M�<�� ��_�<�5*�kF(�y�oDL�<Q�&U�z�J�³�N�4Sz\��*c�<�7bpw�JA���o��|�#�j�'�y��/������9Yh�$�� Ǧ�yB�A� Q$4��f$R����=�y�[h���R
Q���b�%���ybcJ�8��Hxc�ĜE�v�t���yb�F�¬D�a�$+����f���y«��lj*��^�V����q�.�y"BŮL����֯�0(������y"I�#.;��UO�%F#��r$��y�HS�Z
�j��X�EB �����y�!B*/��%ZƩM�EUT������yRKS��`��@>�:�ie�N�y"�ό ��h{@�ȗ$���ӭ�%�y��d��S� ��^�k �K�y"�	o���qᙝ�������y�d�;K��-Z���R���yb!�Ho���5�	H�I1�T��y��^��|�"/H>M�R �7Ɗ��y�D[@@Q��gO,e�	*'OE8�y�eG�WRơBQ
�|���)�I���y��/�H�f���g?�샶X��y�̑<�j* ��*�|صEY��OL��ȢJ��h���	A�b8PEb�!�DV9ef�$ȠD�H���P��_J�!�DL-�\iQHO*��8�%G�!�$\"�$qcUN��2�0�O��_
!�D.h2��I�4�L��eKO9s�!�� ���Q�;�H��f�-D��5��"O�Aې� 	A�dFo��^�H��"O�(�jF�g���-�>���8b"O�,+�M�)�^M�'�7>��L�G"O$�F���]��B�����"O �T�Z>MN`D��g]����A�"O�Y2%֥5�$�w�E�-K�k%"O���V�6SB Dh��FK4`��p"O,�0F��8��y0�(l(L "Of		��S�;:9���]<Gufc�"OJ�d]V!���jD��3F"O8D�%eQ�G��xr�E�CR.�"O���(ݨ��9��٢,��% �"O\	��"�&���C�G�)!��8�"Oܬ�wn�br�wmȽYZ�q3"O�mpC_P~l4� B�2�L��D"O D�eҋ+�L��A���,���5"O��|Z�C5�ʻ���pn�v�<YEւn`8�U��*P��}�<a��ۭ S��vBH&(r"£�C�<���Y--n0a�$'��i��-~�<����n��K'��) "b�h�t�<�D>
�R����G*��e1�#�m�<��̜�4Az$%ٴ0&5��A�b�<��(J?�Y!W�I�Y�^�	�N�W�<I��3B���֠Md瞱��!V�<�3����\�֣_$~~,�4f�Q�<ˉ158hXpMY�eQ��@&R�<�cvj*F��7������Y�<�7Œ2Bh۰ʯ)r��`�U�<&�F
/A��S"���(��a����M�<q���@@#��N%fV1@�h�N�<	�"%��P3�J�5�FmM�<1��[ ܼP5�L9�j�`�J�<��]�u
��cJ̑~����M^P�<�&nM��ܠ���)0="e�E�<�OSo��ǋV�;Z�A��A�<��iIE|��:A�]�1�wh�|�<��9�r��� �-
�%�`^O�<���Jt��Z�oR53JXy�G�<�%F _���S6$�es,�@�<�ʂ!>D�떃��"��H���V�<��˞(V�;w��5fIq���~�<���6.�9[ ����a�łIs�<q�σ�%�������e��݋2�Wq�<�I��4�D���a>�`��r��l�<�� \G(��E��1pXӦG�r�<�FU$3m&z�I˩	�-�`�o�<aC� &4i&o�%S���áb�<����i�� k���<��$	g�<)2�K�~�U�KΜo3�@I�+�b�<�3�� c�ȷ����$=!��TJ�<��� $��q��gA�+��iz"��H�<	c4`帍!�
β_����wD�7�}{�n�����+�X����*[�Cl����n��\t�����.D��0n�S�����ʃ> ��3�.D���Q�1�4*D�jS0ݡ�-/D�P��S� ��T �"@�"�}p��-D�p�Q̉P�Xᔨʗ�>@ˑ�9D�����³:(����#+A\�T�7D��@#kS�n	P�;�,�5��l�5�5D�t�Ԏ�$a����a�ƕ�h�yS�>D��(�AA�m"� �8Z��A��*D��@"��8�8��w@8�J1K�+D�� �Q�,Ԋ��e��%�T�����"O.��W��?=��=���;$��T9�"OеC�KTK&L+��V	`�8���"O�)8��S�L򁐌Q��9�6"O���*�ؙv�^�q8L�RV"O��eL�=()v�cl�_��$"O|��ƇtaÄQ-�� �aQ!N�!�dϖ9m���ڋd��� �o�>|�!�Ă���(�Ҭ��)�`MQ�.Nf!�Kgzt0����������-��cQ!�d\�-� �Z�I�ɚ�"��!��5�L����>Zȶ	��aW�i�!�Z�� 0EK3��ݪ
H6Q�!�$��_�ܠ���|�R�K6�]&�!�ȫU&�Da�H�N峇���,`!�Ą�H�v�Ht��5��0�2�Z�t!��QR'L�$���FI�K!�ąu�$��R�����K���!��\�H�$R�	�P%���äs�!�����
`Μ&x�����'�!�_JP�ub��x��xa��>Kp!�$�T�uBBO� %��['g��m!�5\�l9B nq�V�G�<o!�DLX]�@#5���1�I��43�!�
;B{ب��M� ��p4�� a!��>*�Q�E�ݰ�V�����Xc!���+|a�c&���|x�D(4!�dT�7!"{�Ȕ37ڄ�z�$ԅL!�$�`J��y���8I�p��!�U'R�!�$H"&��Ip'_�k4b +q»Rc!�D�3UN��*��5*D(@䎴�!��PO����j�=�:��!BG�(v!��C�ldN4�wƙ/���;�y��&]Bm�������.�N裢J	$6J�3�΂"�y�o�<���B�!b�a��Ϯژ'`�Y�On8��P��C�$$�%��F�5��Cc3��hb� ��1�īߝi\4d�R��|)�
O��t�^�mgL�� ��0�����'��@C���lܓ@Tq�T`�T��c��S5Z��ȓKo�#R ��c$ΠPb�&`&0�'�F���e�S�O�z�Y�ςMٸx	 ��&|�zٲ
�'�`%#7o]2[�Q�玔3v��K�y�.T�u����7^� �!�L�2E�A�B�8]{�Bቯn��tI��44��f�0z���B�WH<i�jҵYh�#�f�4S������ _�<�b�I8��$9� �'�Xxf�W�<)�@1|������6"��u8-�g�<!�*F-]�H�ҫ-��@6�b�<YAf͗(ZxY�,)sF����ʕA�<��L�6u
 ���epbh��͏f�<q���+h3�������J��s5l`�<�m�,h��������$'X�<���M$g�"��ǎN%z�R�P��[�<)&D�N� U	gJ�&_ST((��M�<1`�͉&��`� �L�z\��f�Q�<��N�'
���REnP�$�v́��L�<��1�R=�$�^F(���O�<�!bX 9�,}kS�T�a�h�H�<aP��?QRdIT�Տ���yE-J�<A¡N28��sl[dxl���y�<��G� ��U욍0)���(�v�<�g�[�bo����LI�+�考u h�<�㏗.���AG d����B��b�<ٖ-ɽMDd����G<H��P�<�  ]k�
�ui�`�2O��	�L��"O��f��v���5���$Ţ"O��23�P�p��%���K.%�L@"O��P���;�R�vbF(݈\�"O���ƫ�:R�h�PBH�5X\U:�"Oິ���3�΄��lƘZ�h�"O. �S����mXrL*y�&	X"O�LJ��+��;�L�43�~�� "O|@@�(J�d}�17JY7C�@X"OR���ϕj�~8X£
k�b	3�"ObhpC	@V��	DD>��b�"Oܴ�I��D��"�U��A�"O��S0�7�E
����@���ȓY ����M��/p@=�сE$:V�݅�u0!��h�L��7�ҢB6��ȓ=G� A� ���$��'_9��J� �1"� y$��C�+P'|�*�ȓX�eQ`�>pn���� �@��T�ȓ8��hpĒ7 }�y�D�F0@����/x�]0���<<��JƂÖT��d�ȓf�䬸b 	|��M�@�M�3$�͆ȓ:��`!�+R [�d�p�+�\.݆ȓ7\�a��+Z
mKډ��HN�sQ����;�&y�W�"�N��F�H,Zڶ����%�%�B�9[ �� �ϩgxTمȓ޼�[@���b����S��` �مȓlL�v�A�2���Ď�=���ȓpY�9����="��������Ԅ�|��� 8b�6����{�����P�a��J�[}����/)�b̈́�Z4V)9�̖k�e�qc�Ӥd�ȓ@=22�иK��e��/Fg��Y�ȓ�V�`I$(�:����<0�y�ȓM��,Cf�}rP`���I>v/����zI#��آ�i�e$s���<�u�r��b�״�h�\t��� �ȼ�����Ƙ��"O��p	W�LC��H�d�9a*�;eH� �v	�$K�?��R�BS���'��!��; G�!��.�����'�d0P�߭*8A��	 8]hU��&�͊��9�r�c�E�����H�����1$�<ul���*-O,8�VOǎ#�t�3��Wm�\y�/�C��B�OCB�����̟�]k B�I?]�\!�JU��a%� >�ʓU�ZR$UZ� ����׽"S��Bu� ���m�H��E��#�:���m �B�ɿ�tu�v��P��(���*F���3�׆i�P+�i�(�JI)�$���'.����ż42������M��X���*԰]��ҙ-��HD��`O��BÎT �څ�"N%B�Q9�$��6�@	2�=O�ě�͔�4����%�F�t
��	��D9bC�
�X�Z �I%��ܳ�ˇ� X���q���Ga�]�pȐO�}ۅ�U~�>t�0�ȑ(���6?O^}��k	��<�-n��Y�!�}�6x��(���5�v�#��ʷqd=�$aU� �!���.J����Iǟ g�ӣ�H*?����ʞI�f�!`���?������?��#`a|z5�'���a�IԿ�B�����P� %"	�n�����̪HH�_
@�����&A�n��3$��X� �<j�`p:��F���O�����^��\y'HM�r�3��I����R���.���`�[�u��9RaK�
z�0��H�l�<E2a�����ৌC����f�R�I����o�)T1��uKy�|��ؼr�6��CX�V����֎�M���3�Bi�S4U
$T�S���1�B���Oٛ`�tC�ɚ�p��W�#��xyf�Y�`���Q�ƻH1d)c���f���[�(F��,�B�/O�L""ҫ[y��a�K�+�έY�'�м"F�Ҩ��dꍤ-̎�Z0����$3�A��J��t�l�� �]#��M�rџ����֮%��d蕄D�����4�{��Ť���� �"N>]2��g,$�&���@��w�}���ٻS2�0p�����?�֠��
��Xs��R��j"$��<��A�6��hb)ϩ Oh��.��h#�J���a��ղ��Hw���to�"p�<���S�? H1�@�(0Fp���iz�f�
��R���J���k��S 
�2EM�CyB�Q̬�⥈�%�$D�B��0?)FAA�@�ޔ�$��>���!AFEڶС�+<L[<	0P#ɽp�ԍ��x�T�ˌ�$�#t���PE�zp��0f�7%���jTN����O�D�6�^(D0����T.QX��jO	}���� ��J�����=�����+��0���Ad�3:��rOI���!�d׃��!��!�?*��&?�`'J��N�@�nƷ-��K 	2D��`�IX�]�.X��m�p�b"DB��Ř�zwB���G�%E��O��@��O~R�.e���Kۇ�v�ڷh���p?Q���=*�vh��� "`d#%�A�]�E����60P↷QU\�a��,ܼ���X�2�8d��>e�}1�f¼m6�����A�RY�1��K�6�u�1�ElU��kVFKW��`C�"r���v�Hx(<9B�\&`p�#�X�6W<]s�qy�i�b��H�$�.m���U������~�`&V�
p3�gЦN4���bp�<�VcŨ������rup�z����Å)��#O�rwt�b�&r�'��r�B�(�-I|H��)I/h��U��d�۷���
|(%f�Z� e�d0|hr�H�@�Pa`d��-2LO,2h��_���;@E�)Y��X��'�PY�W�J�R�t�� � EA�3!f 5V��
oAx�H�+�!�d�;#%dR�!�+e㔉�c����1O���C��碵;Bb&ڧC��ä� =����c�]�>T��ڎ)����4:��D�C��8����B�3!8m'�9k�H&u�Ć�<@������ �`��7� ����ȓp�N��ҧCW��h�ЋT�=��d�������-l���vB�y)L	��9f����	.t���b[4$2E�ȓ>s����!�� �э.\��ȓ&�X�#�ۥN�>|�DK�����ȓi�=��(��+r���t��Җ��ȓG���/�0�U2 ���B��'a6����P:�L����X���!z�!�CM����$͢\�V�3�n�!�d�sz4��Rꌳf�0��&��	W�����'#��=��>I�B��;���⬌*_/�!�i=D��b��^�-��Da5�H�:�����9D�)V�0�v�qB�2:��� 9D�,D`��a��� 	�(C��r�. D�ز�\xW�J���:!� �!D��选� P(�'��al�d�?D��9��d�ڬ��ոr�h@�0D��z��tV6�l+L/x2�q�0D����] (vU�g#��K��z�;D�t*��=�څ�"�8L���/%D��s1�@&I�0�áEʰBh�\��?D�Lyfe�2x����I%+/p}���!D�j���=��Q�bA6(m
�-?D�����.8�R��׬S���צ>D��+A����P��2 �)D���r
����i"T�X�:���1w�'D���dI%)���$����5�cO%D�|;�A�>\�������e�A��!"D�P���L�2q��(]�x����V�"D� 8UhBY-X��F�d+T�#��%D�8�a8^ y�A�q><��@"T����hJ���2#��>���"OXy��\�1��
ŨQ������"O��1a�MJg��3�ǘ�c�x�4"O݀%�ۜ"M������c6���"O����E�1�"�I����A�@�1�"O�Ւ�d̻����w�WE�8="4"O�e��gߚAjr�`w��a�Ȥ"O�
�(T�
�I���+2J�0e"O�q0k�<my T��+-d�գ�"O� �۷&�	`1;��F�	��	e"O�%:q��T�|�5ዩ �X��"O��a�n��h4�ŏ�(S8t�j�"OX�#bT.�p��m��l-� @"O�1b���3�����mK�6B��`"OV8Z�I�04	���6\�X�Ԭ�1"O��A�jR�6�M@g�w� ��"O�̠��~UR��vl[�)�$z�"O��!a�A�/>1P+X��HI��"Ox�����(�к��V)�䡩v"Or���O�K�NaB0g�$<���j�"ODe�!��3l�,�ڃ��<\V��kt"Oz|��[#~A��P�X���"O̅�pj �z�0@T�L�*�"O�0�Ŕ��~�"
Z����٧"Oj<A�:8$m���M-.�t!�"OʴpD�
�o�.�� �4���"O|�%N���-",��%�❂"Of��C$[�c+>�pu��E��,�"O^� ��Ԭ\P���7
�9�Lц"O�Y۶G%�*yaG+�	pPP�h�"OT!ƁQ:)�I@dI'r0��h�"O�lx�g_�p��c��43:,3g"O4��
7L� ��f`�:�!!3"O�Dk��N*m��qrO�4`N�iڵ"O��U΂�r��U�#.%U*���"O8��d��)����C��a�"O�	Ht�׶|f����N�^VH��"O�g ��P�0Q
�NR�L3f���"O.8��O^>�ҴP4G�,7�q2"O�Hb��DP6�Ӷ�D6S�2��"O�� �-"��A[�&焅9e"O�8��A�6V,��0�5>�H]��"OZu��a?.�v�:�BO7�6�"O��RrI���x( �dьUc"O�%Pc��.
���"��F>;��	A"O� �R��� �m��VNmH�"OB��0G�"&�l	�*�2zGt$"O�B��S���+���i7"O^�p�D�HJy	�ʰI$���A"O����&�� ���J�dU.X/8U�2"O�h*��4m#=���-[�}��"OjŰ�
��	�#�	q�U�"O6�25�U?_�v��sV~����"O e���.��cB��7p0@ɐ"OHe
�� �5Ж��),Zm@"O|�s��a:��K�a8���"O�̰��E�K���p��.w�~ĩq"O�=�j�4��Yb�
����"O伂�B�7Rc�ĳu�U)Aj`|�u"O`qB��wM�:G�Z3�"O��#���Jx��Q:D8R�8�$�h�<��'��1b 0,��`�/WM�<q�_�EDr�Q�
�g�<a��D�<a�)W7}�Ա�F��0n��B*A�<Q���+iTu@f/S��Rl��D�x�<����*<��ۗ�ůDd�,��-w�<��%E>
�`o�%#�z�I���t�<Y���`k�\�l�qRz�WMY_�<���N��+��+Vi
�(P~�<�ҼB�*i�L�2"�	�q�<!2�H�jȑq�I\�S!��qNEP�<���8�QQX�J�93��P�<���ٛ92ZP�Ү�nm��AEh�H�<� �%;2Ń�+�ntb�
I�5T4�D"OЭ*0��}KXU��Q
)��"O&�FB�
�b�
Ʀ�T��`�"O.���R&�̐��@)Р��"O�|�pM�sI��q���4�؄��"Of�5�*�(��
��-�"Om���C�([��K#�^�>��F"O��$ۉ�\\�E ��\�R�"OP��F]4F��v�5/��E�"O踳ÀC��p�#��2 ���g"Oz ���l��:���P�jm9B"O��q�ɯ>����r@�ku8�8�"O�$�#��aj��#HA�p��"O�����~ʘ5���޷*�Μ��"O�e0�C���ã�
L� (��"O�5��'�=82Z�T�T"���"O�y��ɗ	��SD� +n���"O8A�$�0rFh�'�T���"O�"��ڑF@�i�@�(w�Z�ّ"O�(�d�<Z��L`!��t��;�"ORpAv�ö����M61��3�"O����&�Q7�\��ɀ �N�j�"O��(�1�R����qƶ�R!"OHr5�)G[b�0����n��r"O��[SAQ�}S����\>:[� "OH���L�Q�(0P� �o$:���"O^U ���3G1�ȡsn��b�.��S"O����T����$���*�"O>E	p$V�?�y��߶Tz\��d"Oh�Y1�ؘyP�IYC��8j��Q�"O�]{4�V�?@�l �ϕ�[��X�"O
�8f���+<��g��Kx�CD"O0"gnJ:(�tX�d�wߢq�A"O�,y��D$-�(b�F:r�%J"O�%B�*� �bls���Hj�"O�9R*W�!�^-+���e$Y�"O �ʀ�C>��4�5�ä<�Q˔"O5S���{�jR����R��"O��C썠i��( RC��a}�A��"O�Dz0T�s@���5"UB���"O�`���8'�H��!�Q�l��"O|�3���0���8vO�<f&�5��"O�:���'{�:�J�LR�a�95"O�ɩ@��:e�� �
�	'����"O
��qgˍs���i��ϨC2"OTx�%Й#�������q"O�r&FS3>�b���*W��`-�yr�f�:����S��]��lA �yrDʍ0Ϫ�3�c�x2|�UI�8�yR�Yt`a�ń0x�يm���y"d�$CdTm��cO+��A��CR��yb�E�`��%�:)�� 򔫍��yIِ�8�!ǸV��$⣀_�yr�5\anm��ė�bh�f���y���Q-��r����2X
�F�;�yR���p�]is	���܉j'��=�yٳ8'���K��(���+S��y��8/�L{DC�-=:.�6�yB��2� ���#�� �F�ڤbϋ�yB�K�b���3�jV��|����>�y��PT��!p# LO�^��#� �y��v���.LE�l9��A��yBɔ�RE�UoՔ*� �u�^��yR��4�E��/�@%q�S��y
� ��0͘�ls�$HW��$X��0��"O�D�����Kl�E9���;X~0� b"O�Se��a�r�`gI
=k�0q�"O�8���	ژ���gH�[m~@C�"O��z⌛,�PS�FR�rt�u��"O���	�d/�L�!BOֶ�"O<�V
�L��tk޾H����"O4��V Ë?��,����(W�B}s"O�M+ J}�(�Su!QU|e�"O���4���/�:1���H/X0��"O�Ȑ��7��t��	�o8~D� "O��z*�W[4Y�(6�p"O���¸er�,��>����"OlH:e]������\�*����"O�hS3 W�@# ��:�&"O�	��\�uNEP�C�2��5"O����FL&p��H��L�5�V1��"O���'�>�pt���F�Z��#"O�\r������*Ԧ8�v�7"Oz�ˑ�(���ϼ�MP"O�(G�ڜz�]*�O�R��12�"O�(*$��'s��5���+h�"O���*����A���x,�0"O���S��0�!��T�P��g"O�ڂD�P���5�1x����"O�����>������V��5+�"O�� ��/�*E	��͝X���
�"Ob�h#�קN�^usfo���}��"O�t����PО�ì��)�j��`"O(�X�d�6�iT���T�Cv"O�\���#�.�1�R�s����"O���B�2i�8K��!~v2��A"O���$KE�j�p�D�(+`�0"O4� «,a�b��qh0S"O�LX��ƐԶ)x�ػUwd9D"O��ya�S�vO&!ס�;Ħ��S"O��U#�:HӴ\���	j�"OJ��$�J�XI�����96�6[�"ON`��^�)0���GIA��0E�"O�ā��.��%sc�;q�8�4"O }�lL)O �`±cE �����"OƑ��K:_�zISl�5H�٠ "O�5"bt<y��	�)\{�A+�"O~�
�'5��Ъ���$.,9�"OJ-��X
�� *V��j�X{"OR��!ɰa�ujH�K����f"O��('Mܪu'�-���0�����"O�h j�*	��]��ΐI� ��"O�I���4�L�E���Q�j��E"O� �r���o��	���]!O
 �Y�"Oнh2bPKLJ���o��A��k�"O�A��mV�s%�@� btnd{p"O��� ('��}�.P�Zhhy�"On��6�^;5�8���CPF6��"O�Qk@G� A>���ĂRK~�#�"O����Q�*)�l;bl�t2��2&"O�
r���&r$!GMK572���W"O��PaU(Y�$5r���j��	�"O��S)9qm�DI�5'��L"O���aMЙ^�v�����
c�p�r"Oa#���#�p=rvBŔs��<�"O4�qqDڌI?|�� �Da��9�ҘH���#�P�h��I3�(��$�����ce$��Y[��2��-W�����Gx��TÜ
��S6�
�9"J��cJ���$�2�(O�>� ȱ��̃�e�a�p+��Q�jx���i�}Dy���W&n���
M�^h��r x�<)�O=<���Nļk�^l�u�Q���H��}B�e���'3��=����&}��S�Q�vVVy'�t�%�)��":r@�D��,�<���K<��J7d�<E��'�DhE��Ο�]�(���e�"�MS�(�S�OD�ms(��7E���@�a����S�	��0|����B�r����h�f�:�H	X�h�d�2��O��I	B[�q��
&���8�L�056�O���a�,akn�!QHK�.\%���	�_����-"�D�#@_�,Ȝ扏I��$jq��S��"�e�2St�y��+''�@��Iv
�.?NbYp��DP��}�'{���#Q��jlyj���a�T����	e>�Ѐ"Ȏ`��`�"Ň�)Ծ����0�I5o�Q�������7JRN8�e	�eǂ��6�xb �R���	����2���U�`ʇ�S�zr���U��>a�&3�S�OD���əd�HaydڈҎ��ٴq�<�<E�4g��	̲֔�� Ff�����rQ��b	�'��E�@-%̝��ဳ7��!�>1��-�S�S }z���d��)'�����7_f�OL�������d*x�h�@D�w��"fĴxd�	�#Q�"}�ダN[Z�Y#��m�:py���Ц��I+�S�O:	d�Mx:���B$�$���'G���3��_��Pб倊2�|�	�'i�q��ެkz� �f�ɟ*�5��'��Mr��1άx��
���fC䉩}'��#c��75p��ܔ6UB�I�9j��jB�TQ�Ʈ�%}�C�IJJ��" ,ޛj�����܎1M~C䉔M/��!��en�Q����7��B䉽.�f(�i�� f�1ϔ��\C��:%���,9U�l�0ā�1n? C�	�4�����OӒ&������4O�DC�I���]���FH|R�D;5�pB�I�5�J �P&^����F ;�C�
Y8�h����5���"��)V �B�I�!h�hy��]� ŀE��H�fݪB�ɦi�l�`"��hxE��ޠ�TB�z�5���0P�ȤG	��C�I�6������e2���ؤp�C�Ʌc 0��e�4z���Kw�՚ڠC�I5PJ@��mR�d����9JXC�	�o)�))�NN X�`@ �-�PC�	�8u��H�T?Z���Фn��C�ɞqT�<�V(͓r�^�xU*O2	R�C�I;F�<q�en�5 @h�#2��C䉗b���;I��VzPq��M�|C�əJZ�����|�T��d͆�fC�	=Z�!�q�_&.xj�hʀR0C�I#��Y�ecڰyXr�((2RB�I<�f!��X�.֍؁�V�BHB�	+S�nhQW�9�! ��'oFB�#L�-B�
5i��a�JS%cA���@�L�[3���H�ٺ���*j !�d��i��I��恪,��I�IA�!���I���B��S�!�%��<x!�_�
�Y�BnΈa�e;�eS�+m!��{���ArJʐ)R�f�a!�$�mn�k�%5���^9�!�dP�# ��tn��I���I�!�$��r��-�V��k]��"�֙�!��8.�楹��B�1Z�|�H�4-�!�DPzN��kA��%k���ǡ׽g!�$ձd��K@�Z6D:D��r`kZ!�Ą2�9��O\�3rȡ�fE!�� ��E�e$�a��^:��ҵ"O\U��F�Y~�PO�#�
U�"O�0j��A:���1O��}C%"O�����
 m�AME��"	�"O�iqSaũq�@U���)x,�3�"O��6�P�.ABQbդ��|P�+"O�(҆_�Ъ�c��I�V"OT��6�1oy��ȌL�(��P"O��J��\�2k�MySВY�J쒧"O���'{f���M�7��@1�"O��;�� 9��Y�>�8E"O�	�`%�
[o����Vr��h"O>���ΓA��P�b�Rp0"O`�d!E[��+�E� 	��"OtP���t	��JE�P!yޘ��`"O�Ҧ�ڀС`� �5��舑"O���D�A"pU�`*�_Z����"O��E�b.�܈O�7<��@P0"Ol}��&��I�2��у0��� "O��c^�E E��SRh{���y���P�رRǆH�
U0`���?�yX28-HlpA���*�#���yb��.0}&�^�J"d8�J>�y"�_�\ �% BU���
����y2!��L2��`�\�ZQ0ԅ�kW$T�QJWC/��8w��qҌa�ȓ5��+�*Ј]����b_�hԚ�ȓ6/R;dB�]�zH)�,384B�I�v���0�"�>jV����G�"B�I�a����/S~rħV�B~8B䉸(~�u����)c� �Oc6tC��.k���ф�+h�:�{�*C�ywJC�	�`D 4s�(V�	�L�b"O��J�f��Av��f�I*:��|��"O6}�!����ȱ����9!ft=@R"O���/�<g���Ui�+a�4�"O�(�5jǂ^w>�2��)5J&4C�"O��{w�B3.Ȣ7�Ša��	��"O���TIٸ���!�,��V��"O"*N��N�A�!N�m��C�"O�y ���_��y�`@�%xc�"O}��̌,� �鄀ۄ+�dE�V"O�X��0�L��.�9��1��"O��@ ��M.�1��n�S����"O@ �� 4�ƴ�� E�bP��"O�ah�@�$o��ԫ��1��ij"Oz�a1"δ���
�ʜ��U2�"O�;���(�αS$iФF�.H�e"O��i�]�h�!��*J�d��p�c"O\@9������HKZ P�Bp�"O�� ' �����S+o��`"O} ��	%��d V���0}n@�3"O��C�C;HA��N+w�VQ��"O"l"�.�a6���5�L���Ԁ�"Ol���o�L]Jx`
��E��ؚ�"OxS��<J�-���ձ�l�hv"O�Ą���[E�L�"OPir�%�_��e�Q�CaP	��"O^P#q�|�r(Z�ˇ#l	rX� "ODqc�x�6���Z��4[�"O���ϔz3r[EG�[�P"O�7iJ�no�fj���.��"Ot�D�Ja�1�ө��5_ A�"O,\�@'=�����׭PD��bC"O� |Y���	]j���F�)b���"O�<�W��T����"zQ��؇"O$<j�/��]x���A�I
s"O.���Z��4˵C�;�BE��"O��r(��|-�F�èe��$ �"O�P����8����O̹�B 0"O�}��BŠ}v��8d��tB���"Of�A咝0tr�P�ְQnD(v"O�5	�O�D'ݣ6A�La*(Y�"O�9��@ (%������&Z@��"O�d�1����gڤudʵ4"O�4{���<Kv99v�фaSV���"O��Cv��)mEJ;o"H�z\��"O��Xe:f8���;]^�IS��N�<A�=>,<�2��C^���UN�<�chѨ-⨡Jce\�N����fW~�<��K�\���n�?�����y�<�dh��5b��F�Z�[v��	�w�<��!J3M[ h*wcaD%>� ��d�@�	�3^w�L��˝;��H����|8�,;V��]� �� 0̕��X�����IA��(;�#R�z⨇�$F~�[U��!2�4y��ИMd�@��1sv��Q��0W�v�@6fļQY�Նȓf�R%P..�b�v$۸F\���ȓVx ���a9H�Y���\x�]�ȓd��P����~�P bТp.q��``�B-�]��r7(��s����ȓ8�0���ݵV�J,�2
>$�Y�'��~�
K<LY� ��W	�x���O��y�M� >M�%�w_0ղEe��y2�b\�f.F2N�E����m��C�	�b"�}��ឍp��$��ή.7B�ɴ/�Z,��Ȣ��0x���<HB�	�C�8�@=-.d����Z�qe6B�I7�@|��cW�nq`dc&�����B��/u�����$0�.N�lA���[�<i�☒w;�}@4 �z�>8�Qd�[�<��G� ��ܑ%�;&����eW�<٧�� h��CWEm�r��C�S�<ٓˉo�Ly�Vn� �5Ȇj�i�<1�>]% �PO
�u�2U��A�d�<)����&c
�2摀��k "�d�<!�c�?�� % =�:<�g�{�<�u�Vv��R�E�Zv�����Q�<I��K�c���J��٢Akz���*VL�<���үJ7�Q�c
�w$b�����F�<���Q��R3B��*g0`����l�<A�FI�~�")��f��I;��$�Hi�<	��)CbI��O��U��Y���d�<�b吧� @S��i9�};�Qi�<yW�dt����C�x��Ass
�g�<�c��M�L+�!_9�ys��c�<a-��IX�8���=&�qc�
�c�<�tj=k�ĕ�w�D�<��fC�b�<�&k L�0ԀS�ӽq60��vBMT�<i��N�h��hQ���K>Ś'M�v�<a���
4��z��\32[ Pd(FW�<�V�J��L`����s���U�O�<��D�`��	��pڲ` �Yc�<��
Wސ�Y%B�7[V�Г��y�<� FZ!	�goM�:�����\q�<р�^�'��h�)8��zЍd�<ٱ�D�R�X[F[,da庑��]�<� �SV#�"�*��փ4��b"O
�����|�dEj���H.�DpV"O�E+��D�FR��Qh��\/�xd"O�@���K�(��0IR%�+h|J�"O24#���(g��  �=�L�p"O�dh�(*�re�\>k��"O��&�)�(�B��I�"O�%zV ��4���B�*H����C"O��1s�G�x�<s��Š�$I�d"O&UivE�8����"��T檬�"O~�B�����jݺ�p'"OV��r�b��-�f*�=�p�"O�$ V�̩�r��cD�[�PMj�"O$������l�X�BQ�{��4�'"Ov}3��;i��x��{u���"Ob P��m0ܘ���C�8N�9�"O�V՟�^��5�1y�PͰ�"O􅠇A�������1��"1"O���1�9st���%��"O�	j֍S�Tr��,�2�Yy�"Od�ńG8_ȴ��	~�y+�"O�0��H�
P�V��V�]�P<�3"OH�K��U�K�����l� �H(�"O�P3d�51D������ I��Q"O~�sΐ�[�1��A�0=���"O��5�K"5&�:��5`���"Ot��Ĩ	4p�X����h�tU��"O����   �P   �  �  �"  �-  -8  B  �H  O  ]U  �[  �a  :h  ~n  �t  {  H�  ��  ˍ  ��   `� u�	����Zv)C�'ll\�0"Kz+�D:}"a�ئ�Q2�}����u��h�ӊvІ��狂?l�X�S�Zw7$Dqp.΍pL2̊ f��ʒ�96�ź��M��z�+��0fJ$7�I�d��]2��Y"%�w\��`3M����9���9/zL�:BA�q��S�I�&���ަ�2%��q�ڍ�Ф֏d��)؀@M�>�`��K�9�?�!@A=T�*��ޙ$���K�`B�'�r�'�� �0�D	��l���P
��X*�b�K�'�Bd�o8��?i�1��?����\kхI�=�:�Ȳ��
}�cZ�X����M#�����O��"3��� (�+��G/�4�Ԁ��~��U�I�E����6.v���	�,|�<�g��m���p,����9ⳍI�r��Tk�O�	K�	F?���-1��+q>�#6V�~�zD2S�Y���O\��O��$�O�d�O��$�|��wY|�RԀU��J��c��x�^t��U0���q�0�mZ���d˦y��L�9�MS��Ek���$Юs���r��Ko4���֩>D�I,B��u�۴�?�S�.s���U�;n��͡�̖�\w������e�ԡƕ,����!C(koXtAN>Ni	d�iS&6�Uۦ=�c�gIo�lQj�U	b�܌!���u�[S�]�9(���1����B�b����(��0�s ���M[U�i*7M#3�n�C���FkHM�'yQ�0��엺Ԥ��`����K�4E��vhj�\�0CeR�8�$�"���g/D��4K�� �Ks!�'
u�$(WdTN[�-�l�4� 7�]ۦ�
ݴ!�XI�'�
��rd��FZ�h�DqZ񈁑;Ђ`��+~��|��Y(���Z,T-�aZ	�`�����%����7�0�{����'�8���KU�#�������L:�4�?���-�VP�(��</���0I (Qc��?���2�?����?A�֧x�ְ�ԂA)}l(�R�iF����(��4Y�	J(��+�`vӺ�:���<V2	���0&�<��l���`&�0-�����! T�Գv`�M�5cTc�'7B5�,O���'�ZvŲ���1fg��E-U�D R�'��|��'��W�<��X�����	�[���c��)����� BB'Ǟ
��&�����MϧO�G�'Z^b�+�E��K�i�N^��?�-O���bF���Im���y硘�����"�rD.¥�K��?���s ��4R�����O��7!��iEj%8��,ڬyc��)1��H�'xf����&B��*�����
�1�
�k�F��l"�*X�i��ɋbٜ�������r>kE#̝<�� qIڣB,��j/�$�O:��O�"~B�Ú
t:0#
���( �"R^�'�^6��ڦE�|*�!��$�ɪ�Hy:|�P7�L6�M���?���2UL�5�	�?9���?����y'E�<���
�%%��E�����O�X���,LODq!r��3Sz�� #R�J\���HZ!��¢C��c�oGRc>c��a!�@??:5ƃ'>v�#5�NۦY�-O6�ip�'����?�OIg%+"\�E�uEB�{6>�9���OJ�=E���Y=>��AQ�O�e��D8���r~剁�M�q�i�ɧ���O.��+�> )F�@-8t�8I�,El��B( ����O����<�-�f瓅tt`�rQ���E�r�--������P1-5TH10o,��D��	�@�����B�4J1b6�E$�B���H�Y:v�����Ib">q��Y�#��1��	�$�1檙{����2�Mk���]��b;0I�0\�:�S�⁷u'������?���0>QGkˍd۶`apn�.�ݱ)�K��4�M3'�i��	�Z�:4;�4�?	��9/q���ЫD:T5��Λi�������?i����?����?�Qe]0%2�@���T�xa1bD^�-Za�k�#�6$zD-�?;�b���yj��Ն�+KFY	v�@"���	1���C���Q��F��㎅'JD;�HU%�,��J>)�H�ڟ��ڴL�v�'�6���c�>95"�[��U�}B�:�Q�$lZ
�?�H>�SJ�'[��ԫ@@�����A%�:��I�� �':7M�2� �EA�6o��r��5��o��(�޴SQ���"a� 4M�*O����Ʀ!��4���k�n5"s�T3�@�a�x������! ,z~�TQE4��LC��P+q�6M��K�<`qT��v��C�J Z%�"?a��ث�t-�O	{���d*��E�.ł��W	Pܚ���o��0�m�`{~��
�H6��'���0�5�F',�):�9��zQ�$R��dKϓr׸�O6�)�$�O|���<�� B�
26�0�I�Zlݪ��L^��xh��Mk��d~���')Pp1"��J�e�y�H���+e�V�d�O:���.������O����O
�tޅ��O���E��<.��I�]59ڮ`3h�������*��1�O�"㟔 ��|�����e_�sZ� y6A]�B�F�h�
M4.�+���Oc>͓��%?A�Ď�4�j�q�O�%\Ibm�D�M��Z��ZK�O�b>���O��B�>�41AWYLa 9���L�5F�Ol�=�}�b�R�JI8��t�
���5��`y�gl�ޙm�Y���?��SIy�C���葲#F��	.���q��7&Ԏ�*�~�����O���<q+���S�h+Iѓ�
c��à���!��=��ŘEbyY3$R�8F
Շ�Ʉ#'�-jS��&
M"��'%��k���e�V�&��՛��#n ���%��iF�#>����2<-��ӓeI/.<��0C�!a�"u�Ƀ�M����[�'R���Ή��D�jC��J~L1�����?���hOt0�L�^a�dC�I�P���5��O��n�؟D��4<'�6T>IP� ߐ�M���y"D_�xp�-m3��z��ɱ(LZ��	xyr�'�b<�D�x�F��v�z�F�`�J6>� �8���5�v��TkS�j�Q���'�z�ɵ)B�J���zծ߼��֫*f����e� ��y�N�)�0�������a��ė'���6�H�'�i7�-	��9M>ɏ��>扇�P+4�[�K�;B��C�\��$�¦E�'9 ��i@D��5����M-O�� ��զ�����O�P,Q��'5�y9�cç*�͚��ɀ2VzԒ�'^���D�)�cK%o<�8�N�.[@맫�)V�s��BU�O�����C_S��	T���E
�,�*{w,�8j܈L�ZB̊�^0�@��
�
TJj���P~i��?	��h���$�.o y7�է#*P�D��\�B�$׼ɀ'�1t�X��ۆA|�#<ѨOB4Gz��	Vb8HE`�
d�r�{1�I6ڞ6m�O>�|��D�'�?���?I/O(;�l��w��%)��ڲT��T�'�����ɖ˦U�����a�*��%�?ɶ(?��x$�Q�/��P��-X��q�FȐs\�QB�Si���|�S~��M�	:!%F8�H��$�J�(�6��<IwJ�$��B�L>�P�����hG���Q��+C�!�?Y������O|�?��'��:�s�T�!�55�d�(O�mZ7�MK�8ě�Z>���|�T,+��!����V���g!.�����C�1)R�'[��'�םƟ���|�E 9!1P�"5j��b܄�0̑��-#��0a��KK��3�����(ݯ_�<����I_l1�	Ծo#���ᒚ@5����
0��9��Hls�q �%M~1,�<�'��C㮑0w�(.���St��ƣş�!ߴu^���Gx�/ǭ�(J�)ϴq���
�b��y��#����c�o
���N����g��v�'���F��T�ܴ�?������D�/m�����ְ	�x���?ч���?���?�t)HEg�!��R�.~|�*ѦL�x�vmս6��1�'dMY�ѰÓJ� 5i���n��K�^<Ĝ"�.�6[�@�[�������ȅ:1�t��v�9ʓn����	��M�i��J�,�dз�Օ{���)�_� ��ݟd�?�O���)F��p�1'��f�r$�a*�0����즵��Fr��L�R� 0j@�dΜ�M�.ORq��#H$p����O�˧
����)
r�{Vk��,�<q��JP�U�����?Ib��?��u�2C�}�4��-��<�)��4���'RwМ9�.��.dI��P����Z/%�;W�d-�G�ā
�ձƃ�[�M&����[���+��ęT��u�'� u����?���	�OإZ�K�;��A珦n��%b��9D��a6*���w�ф!9���G?�M�/������QREra2�ÒT�~�h$*N��M����?9�����HC �?���?���y�G&pVH"tmT-r�5ۂ(STy�D�,k���t�6#�0-���$%U.���P�	;��-=;U��Ak�� 0��٭Ugn��%�(1�o�Y̧p,d�e���\�� 6(� `E�%A8@�3��G�u�*O&��'f�d�?�O
�TIۃ!^\Qk�?慳�%D�4hbK�z��l��f��vI�I�h�<�E�i>��	nyb��謜�DŇ2ִ{��U��`р#��O�2�'��'d��]������|��͂�0�ů�
/�̈��N,z���bňj�BI�Ɉ�M�<EÌ�B!-L`�рL0v|ҷ� I���KՀ����&N<m�и0	 ��-t�Z��ܶ���Щy��D�2������	ݟ��?	��iL7dؘ��	 �R�l���~�az�;�	��#�[2D]���NYu�'ͺ6��O���.UK�U?�	�h��ӑ�X�
��(�d�R���I���Z�/��D�	�|J�����⠂g�D�`�d4�U�)	�0H��dJ&��6N�\R%���Q����Qumװ!#����"s���"gٶN+T��ʎM0||I0&&�f�:����P�'*b!���Q�l��U��"c��IJ>!���0=����h�TO��~z�ܚ�,�H��p+�b}&�'dH�r6����%	�h�	GyFA�c�6m�O��ħ|bp�M�?A��c3��*���Iq$�%M��?9��Z-�p��O'o�T�P�@�zVZ(�!L�s�L�͟FDY�nϊEǰ�����#� ����� H��\Og��k��ݓKvy�/V����bV}����<hR�i%Hݲ8�؝;l\(���P�eP�Ax�x�F�t7��5���T�u>�$4 �����"O���7���A��y'E'v�h+V�	?�h�"]9�A�0���k�� }+��xpr�@���O8��->}J�����O���O��$��W��3g_n����ԭF�`R��V�j1 ���L0��!r��:)�c>�'���7��,�%WG�7j���6�6mg����9I��k�A[(k��c>1n�+d���I�8�h-A� �4�Z�X��/?�i�ߟ��I� �?��,�7v<��Q%E�W�Q�0�=�yb��P���	�V�[p����+�3d�����HO���O���0qI��=8�4����-@j �]��
����?a��?i�������OX�ӴEK��Ǜ*\��!��S9C��C#�9 3b1��oџI�)�'F��eh��+�oL^x� jɸ��O�?��]7�D/ejx� V��2X)Q`Ô<C k�,d�r剷.wna��GYt�|!�C�S�P��O�d�Oz�F�����P|G`Z�� �c��y���#�|���Ȏ�|� �I�F5�����'��	0	f-������	�q�be�C�];(�KQ"*C���I�px�%�������|�e��g3rdzR ݱsg.� ���;B2iB�0��p�gMP9L�
���[<�<aCC�0���dO�!u�3��6zzU{'�Ӡ�M��	EJ�x��D\(C-�<	�b��H�J>)$���|���:���|�;aTN�<Yb�b,p� &�љ*ee�Pc��ȡ��7*���@�A���5����+���%���� ��M���?�.���ؗ��O^5
�C�5>���ttf<��L�O���\�|���Sȋ[�4B4EȇJ
E�d�K�!d�'!�&  nE1�L���,
}�|��O�)�ԏ�j���@�+e -84g����H?�[��*(�Y)���9{"���1?�B�ğl��4��v�'�>E��W=��R�2�~���O(��?(O�3�%`������?4E����]�Mu����sӐ�o�c�	#��؂'� �u0���ֹ���8��쟀�I̟P� h�2l����	՟D�	�0Zw�B�R��G�w��=p'Ǭ[���ЇY+!o��1d�s���1���Uw"�'d��Orɹ�N� a��PDjD<=4:UJ ��)�r�E�P�2������71��P����b�D�R ��U�`�8�i0��O�ɔ'$�E�����?����?!���/�2|Ife��L���g�O�?�����D�O��?�'�0��-ÿ(�>�[Q&\&U��-O\Mnڢ�MH>��'��)O�1ȓ�
Q�mXT�D��ɚ�%"��0���Oz���O�D����O8�ӳ4|| jB�ղW�����^�7��#1F^8'*��zDK�1�6�{&%!
A��3'(L�k�mV0i3��y��(L��u����&�����'F�Q�r��lX����I�"��뢥]j8���.ԦZ-������O�8��Ix�I�E�^`�����= ڂB�	�2|U�����x �$≟p�N�O��o�S�I<qϐ=���8��RXᾙ`'	��f�!KE�-�����O(��"��ON�Db>�yn�%򢙹`�����V��S;�,"��6!`Ղ���O���E�픧;D�6�AU���E��-��҅RJ���i$lӽhlY����KM*���O2�|b4����x*� ���Z�X�]$�t��o��K B˕;�|�fE�H�jñ"�W����Ο��%#�%�6�ɴE_�YA�@0c��OT˓a�\(9���?A�������d�{�څ(��(o�1��Ț'�&��O�4�1`[�p�p��^�(���ǋ��5�:�T-��Bѩ��S�2�6Es�F~"g��Fe���("?�r�3e5P�����[}�	ܡAVp�yD`v�d�a'"�<��	7,��D�|�)§V���ZcL#4G���'ЁF����4H>8{6��%�>�����)=lt�G&�'�4q�uELe4j���"Z+n`h���՟<����d�aK�.�.]��ܟd�I���;]������{��I��e=v�]�fl�!����/�	_|�+T)~�';1�@b�ﵟt{M�2�HK�F@-@�,H�֮��H�%D��\
$���^�c>�{7K�$ik�DЊJ�Vx���K�m �)$J�hJ"�O�)D�'�1�1O�I�jN�C>���/�����"O��8 �\!����uN@Ԯ�8�^�I��4�̓O����ASέ
'�Z�_�J�adJ�R�V�@���O���O���Cۺ3���?�O����̓�oJx9��ڃb��uhU�C�>�ŧ Y�r��sf�2c��
�U�'�>��f	1WtQ�PmB���� F��-Qf��iC��4��$���Y�$X���A�'\`1CM�n��acI"+���:�V
�?)��iwh"=!�����)HJ̐`��;HC��S�Gާ�!�F� ��qo��H�<� @�>U�'�7��Oʓ:�ŪZ?��I6T������h�
�D�} L��	��d �����	�|JL�*hP5*GNQKl8j�n�0"���1���$1��M˶�*��@!-�'V �<�����������
��"���0���"���9Q]r=�ʖW�2$+Ћõ6wF�<QCg��\�4	��I�K���懌�|�n|ԏJ�w� �OH���&Պy�Q؋"n�(���˧f�����OFts!��5�\�X�+�[$��f�'E�:;
8q�	���d�d�n���ԕo<6\Y	�
+�J {�̏�W���'�x�A��"g��S։T\�6-�|r.��� ΀�R�`��q$�3Ҝ��'?���97p�@v�[\b,ɱ�<L���|R�L� �������-Y|���V~����?���i��7M�O�#|B1�jQ����1Y(�$�c�:޼�O��$+�;�R@����J�;L" �!F��V��Fr�pӸ�n�R�I�|� q��('ʽ��y3(�����P��ٟ����ޢo�-��ß<�I��1��%���SeF�����!m�I)s�F����yh��K.���ؤU�ԯ )�	�d�	Mh�˶/�-|��9mڗ�R�@��-�3�)� <�:t���5�7�G8I6h¤�c�rH�'9�I����ɟ�''V	��,��@�2�Q5/
 *�|=�b�I]�8�D`߭+%����)ް׼E�Ů<�Ѻi7�7-;�4���ɨ<���$M�l*b+�)Iʴ�y3�9��23 ���?Y���?�EL��Ov�$d>o���|�b�]Ƙ-��fL{�24H�*C�8T�Y+U	_����3�Q��H Σ4 (��Bg�<<\�E��ߺBF<$B�dO9&<ej�b�/>},ZgD� �x�?9G ���p񋄫J5�]"ЊY�r.���	�|D{��	�'��d
"eE�1aêK�B䉲[�l\�ҊE(+n,��(;�*�O��mϟ�'c������~��<	f5�l�#X (zaP�L|��3��?�v��!�?I�����ξZx��vgTvtPB�i��Jq'��4O�0���ر����E�L�:���N�9&|�� Թ[�4���gi���K� 8�)3��>N��@�茦C$�cIHA�Gw,����|�'O�0@�G ��ၤ��0 ����I>���Z�ڒ�Lf�V�%B4�t(��I-�?��F��l7ZX�bBP=r����\ΟH�'o"(s��n�p��OF˧N[�C�mL��÷-��cEdȆ
ƒY������?���P����V�:4T)R'�ák ��i�K	����;�1���W3$�fă��G?V����P!\i�\�n�,��%�L&|Jxi�B�O�M�O�.����
E(�J5�L���O�\*��'�
6m�j�O��ɕ�H����"�V�1�HA�NA!�� ��ݒfdC�,����rɗ�+Nџ�!���F�*�����I"W>`C��u��6-�O��D�O����(QXr���On���OZ�]1�&���p��	r'�/	B��1�N?E������
�!J�z�@3�Ӏ�\#�O0��┏t!�E�u��,I�1��O�JJ�)a4eR	f7~�zR�[$v�1��}{�?�~"�H=��k�c\��;�ٷ}1����<٢��ȟ��Sg�L>�$� /�2�pF�Z	�bq��3�y�$����g����Pō��`���t�'D�ɨ3�L��--��$��	:�� ʄ�bgj��Iğ��˟x�]w���'c�i�3%:R�`d+�.!0�����W3���T�aَi"P��z8�}����x1Rqa����`��YT�G�+Г�j��5��,��ӷ �S̔����3g���j��j�'�R���<1�B<�ЁS��S�-�?ɢ���h�HG�P��a�Z��89�"O4=��-Z�,m��{��;՝|�~���O�:C#l���'/ƴ@a��>�
����D!'�(R�'R�>9XR�'u�I��0�$�b#H)`�*q@A�(P�A�J!W��3e �hG�,����;�~���D��T��h2��J"N����զ!��T9��]���3D^�&�F=(��������$P�!2�,|���'�mZ"м��Ƞ1�5
��%SI>�	���Y�nŷv?��PT��"�d������?i��ޱ �6��B�4yq!�C�ȟH�'��x�H���O��'pW��q�e�`,j�.K�5\;@�%�dh����?ɳB��q��pQȊ���ݴ|&ꧥ��G�J� ��g�1ޖY{��&B��9�yµ@��4�"xӐm�^w�D�
H?- 5�K=��AB֌���4��L,?���Yܟ(2�44J�O4��Oy�I�!VWʠJ �"F=�u��P��'2�'����kV! ����M0n:��Q��d�O�9�'�1����#��,}�B�!ĭg�A���k�����O��Dć
���
���O����Od�D}�5�Ce����q�ٸO���E�
/ -*�N�Xq�h�yy�c>�&�,.p:i+�矺Z��1�V/P]�:���E^�EY^:m�]��E��H.��G��h��3PЍZqA� ���#?)�A���I��?��-�$Y�Î;hp�` ��^ i�C�w�j��&�Үx����qa�5'��5D���ԟx�'�B��� �$؊�E�.�(Q���}�xXb��':��'_��{����͟tϧVhsG�H��"��Α�K �\c���Ah��+C��"�\��'E�-��O�-��iZ"Y�Z��lc�Q�m�T_~��$iY ���1w��d���?�eN�$�qk2恞"	�A ӕC�t�	ş��Iq����8�(�)4��=z�D��l��"OR�i�DF=������Z�4��|�fӖ�D�<�Չ�}1��џ�aE&��h}p���K$�����Uݟ���/-��t�I�T�'A�E���<?�\�:C�Q�a�Ҧ?M��� -ZdK�����O�����R(`�x�1���+x�|Hש�}w�0�%H�h����m�m�b�?YTÔן�IE~BL�4����9J���0�
	���?	�2e���K֮x���c��5l(u�����?!�g4��3צ�<�r;7ߟd�'Nyz�|���d�O��'`����$ &�@����b(���]�����ޟ��I�=�"�(5j}�P��G>b?�"��v�'j��|P�c� ��[VB� O�,��'[��Pu*��v��	�0j��'��|G�I�;e�VA!�C�R���[�ŉ0����H�$�O�}J��ǀ \���E )d�L#'�Խp=vxQ"O�,���S3���R4����ɕ�h�����a��I�
M��f�[�aiӦ���O0��
�Z�D<��N�O���O���c�]�זM�^��7�г$��zb�� 3���WJIH0
�#��U/ �b>!&� SB�˵
ڈZ4��<w��[&�Hv��CA4q��d4�1b�b>�&�(����CM2m�Q^2]�z|Xr��f�3_�v��=�3�I"�-c��[�7x֝��eG(%(�C�I�{�~5�$�/�t�:��ʓ?A����N�	�8֎Łp��8�~�Д$��/8h���QXF��Iɟ��I��ԉXw%��'�)�4p�Iq�DE�Q�n�铇�>ot(bd]4lİ6ʋ�p=I%��G�L�E�C%a�:1I$��>rLq%
)y���[�J?\OR�&oÊIO�t�fnM;d|�È�7x7rjj�,�m�Y�h�p�b��i��&�O?P�.�+��'N�O�LqS-_6>T�)ߊ�����|�e� �D�<93�BY���?�R�mFC �����.%���L4O$�cR�	�8����A�!*��`:c��9X���$�$>����퉱jF�@: e�:!ʎ���;O�E3��'V1Ov�++�/q�rlJ��Hf��Q1"O �֍ڕf����pD�(b\�X�f�'���$p6��2J�-%^�=!��Zf��'�����'v>�	�O�ʧ���C�P�������N��E$	��?	�c�&���,�i"����E�W����Я��@ڃ�£w�ܢW)�_Q�	p����FM�^�h��f�P@�O�}�B�ԋ@�$*�o����OHIT�'����<'<ڸ�B�N�jtfBg�<q��?%"��!S?O�D�:WB�f�'��}�/ԂmG���b��&d�Y�r����#�+Sky�(�&-���O���'��ɂ�`�b@W�>G�A 4� �^�k�߲6X����h<�ɢ�Qg�g�X��Yh�lV>O�Uᖭ��f\@L����6��]��F��% o�g̓f،ԣW��9����Q@t�ID~G��?y��hOF��!�Ȟet|��BȘ"���2W�2D���5ƀ�R2�2 ��V+~�ڒ�<�G�):)O,��E�6js�i*a�l�(WL�^�`S1�ڦ�I�/ޓl�j(0aKC	-<.�Pٴ?m���#�iFצ�rc����߯	N����4dr��/^^�'Ob�@	H�TA�#ӧ e�M8�"X,^t� 7�^�4� �{-�x���0�έFX8I9��Y�9��8z��Q��tSc��|1��80�7>�̋w�OA�|XB#I�?��E ��$� ��'91��)p�׃[,��
 ��B(X���]����	�v��ځ,�_l4�p�	���hO�Ӂ���
l20C��Q�<���MǦz��Ɇ::X�4�?�����i��yڀ�D�O��%ؒj��4��U1,��y���O�mе���yq����l-%lj|�f#�]�`����5� �	�n6�|���W�Q�r�	g��}�+ڴ������*o�|x��]��|Q�K|2®ٜ@	���0�3���*VK
�<1���џ���w~J~��O��#Ɖ�i�0X�.�$�$�e"Of���N�,C����2͟6sx\,�hO�1E��NX: aH2D,f��� � G�'��j�8�'C2�'��l�A��b�j��[cY�H�A�F�T��5rEkX�V�PqȇEÃ��zv-z�dɆ�=Z]�O����fI�]W ��F@J�T �ʂPJ�{��WP�`����'�������A!���,wb��y&��U"�9pOQ$��ɬg����OP�=ѝ'��;�L���w���9\�ز�'&��3�2n����(b�����\���Sɟ4�'��d�ҐFS��VLޤ?���ذ� �\'r54�'�"�'�2�z�I��ៈ�'+���բS���R�|��ʧeD6��������F�$]�����9�yp�{կG;jPZ|df��䣢I\f.����tz�T��ĵ)D!Yp�OD	Q�'B@�Ѡ�?B<����'�	 A�Ȃ �'�ў�G|R�-Dځ�wo�!ڌ-ٰ�E��y!��RV��aw���v�	ᖎO���d榉�Icy�� ��'�?��O�j�!���lB�У�S+���L.�����?1��W��܉�ݣ]$��%�JN���i�v<h�s HQ�u� ��9mI4Q�We�`�'h�;���7�m"�G�1D,����8=-R1�'op�����Cm>���GĘ�y��O�%�'��7�A_�+&;x\�b��Q����ejƾ ���G�� 	gV :`�	� �F�(�/�O�i�' ^��en�8}v��@��C��ࠫ,O( ����I���O�D���'�žoNM4�Z=��ƈF9�y��{�pm�0��	O��$�6�I$%	��wɗ&)1���7m�j������0Z�,{�5O��	%��n���BƩhL0TʜZ�V�`!�I�S���ꃆ��9���K2�H%��D_�>IB������'��� �9ᕉ�D���6.I�C� X�"O���׬�D��E@׊^4��0т�ɕ�ȟ����ꎁ1�29�Vȅ�k��ZR��O$���O��v.��b�>���O��$�O���OJ���fƭB��k ���|0҄^8N�H{7GE4'8�A*�:].
�'Zb��9�E9}bDZ[��[�B���w�@6vw���U���G��uUC,B���bc1�ӌl��'�`�Q$��]�z0�ď��Z�[�^����@�O�`mX�L>��'�T%�d�#l���t�A 0�Tb�'-$��c]�R���ä�X*����Bّ���(�'����էݷ5DЌ�C�CG(���cܨ ZE1C�'��'/"�}���ǟ�ͧY��lk�
I�@`���F��!���K8u���L;7tPDC����	����BB>ʓK��4ψ��!��,EF��c���*�^�i3Y$��{�Bá46\!�*(ʓ��P�I�Is�|��h�2xАdKϨIN����4Jq��F|R"�(c���Y�h��bă��y�&�a�jŨ�+�c��Q�����D�Ѧ�	^y��M*��'�?!�OX\�2�f_�wb�ذ�h���)�1������?���Z�q[�f&Hc"�q��j�*=�v*ޢ�f��j����w읧O��T�t��Z�'�|ؕ/)]䂀��J:}�j����S�&�ISd��^�̙��Jđ�����4$�c���c��O��d1��ΰ��$�!��1Ҧ�9^q�ʓ�0?Y&�ȹT]Ȕ��I�$!��Z�RYx��(Ox�86+��T2��:���*jd�P���I՟���Oy�S>����<Y��=NsLmk����;��)�QY}B:O���<�7Y��>I �ώ>����!���;x�X���*�Iצ]&�,`���ˎ�"j�z'�̋1�ر�gI>M7�6��O��q��f���	�O���t�o���S�G��;V6Ma��9A�
aj0qmǟ�)^ܟx�*�đ�������5�J�3�A)3;БP��L<)l8)�+�?��R\ƀ��'����O��������03E�X�B� ��k��i��ߞQVr���O�I�A�O���ɹA���s��n�%�yB�"�5�AM�C��ǆ�Zgb�#�?��lv	�uV?��I���������n�l��sBJ��Xq`���?�֯Fןx�I&����Ƀ�?��"�in�,�d)�6K��l�T|�uG�%
"d�����M��'��dr��?�P+�
\�����d�O���6<?$�z0@�%3�b����Ɔv�|��b�hn��O�������yb�'�ļin����>+,�A�!nDjă�*НM��2O4$��'��HG���i�OV�d�猠hE HH����_�gyʵlZ��͓t؆�K�4Qx���OK��OL �C�wIܘ���Z��i�l@�G0��l�|u�%*�æ!���M3�Oћ����'��׉O�8<Bb`�Gְ�f.Ƅt1!�đ�*U��jC�*�P�p�J�-�V�'�r�'���'-b�'+2�'rZc�����FP�j"�ecu�(^�I�4�?����?)�����OR���O��dʼ�@BĊ�.�)"�-$'��oퟬ%��I���%�8��[]5BA&�
��PA��jK��o���	ޟH�I�����|�I�,pV'6���l�53 ��+�>�����D5ړ�~��&h�ebCB=uS^�s䅟����?����?����?�/O���E� ���7DB�x��,��fh��?������On˧���*�aq��1J)vP�SۗS�B�I�d\�{�ʮ.B|���,�M.C�	-'b�-���Elt G��F�C�I
|�@`�6Ɯo�P�'n \�TB�ɗJB���� �>kS���R�;J2B�	0�����
����2d�X�\f�㟄B���'Ј�D� B^���6�� �\ؒ@�ͯz��Ҳ�H`����w�#92��wY�#Ŭp9��	,i����N�4�{p�D��s5Y1��$l�ڝ#&H?#�zq")��i��O�@Z���3k�:��͛'�Hz��/����s�إ���� a�5(�4A4k A�ք*�	��`�CC�g�\��w=*�`thx�А��N�h�B�"���S�eQ6c���4gnǆ`�7��Dg2%A���D]�X&+��_]N�q��2V�`vb�V�`8��4?�"6��1! `Ȓ
����B��N���dܓ�蟜X�o�=J �����d��"O��#3-Q6F
n���oE4?�r���"O
��	%3�����L�('-��"O��QG��)Py����	�6}�Q�4"Oq���!`�����h]?>;�"O�${��l��R$��(U�ȠHS"O=��+�Z��D�c�Α8��`87"O�<a��)g� 1QV�\�,܁d"O0� 읠ǚd���=����""O$�8`�+eDvd�ϟ��8��"O�A�Q̗���9Y�M��%zD�#Q"O�t�sFR�%�}H��F�i��z"O� 2��d�،=�d����o� �e"O���Ɍ(���y�jL�yd+�"O�)�1,� e���?}�^"O�aS�jÒv}�)
wA[�,���j�"O�a�ˎ/7B$��-�3�А"O8M���ȅ,Ni�C�ZV���@�"OZ���dׇyQ@xB3+ݿQ�|�8�"O��
Ɓ7Za MsQ�W�xlՂ�"O��ƌ�E���v�O1�(�;"O(�� �U���`�v `'"O��k��Ȝ\�*����ߘN�$e"�"O��S��8�PmA��YU��t1"O�9�jФ(�>�A�!��5��8;U"O�h��M\�^ļ�����	UgFL�<)�-Gfe\����&G:���bJ�<��"�1����B�L�Q�������H�<�
*i> k�B)/]0�5f�B�<���׿2���5{ذ��|�<�sbު�d%����0�B�cEu�<)a�$�,1*���62�BI2�[�<!Ot��A��޳D���5�V�<٥��lH|�V�C�H�꜡��
H�<�voB6H��P����1��a��J�<�t�G�1�fuJUc��<n@a`a�A�<)#�B&fi�����	�o�6��3D�R�<�RϞ2P��\�Pf��c�H����K�<�Q���<�<�#�fŕ"FHx�7��}�<��KZ.?�lQ����|�s��w�<� ��iJ�xԋѽJ ĩ[W��l�<���r�ڴ���<�p��%b�<�s�ϽP����D��DK���b�<a �<7"X(!�Ԯ R���IF�<�"��E|�jB'�K�@�Z㣚[�<i�!M1���s�G�^��Ҳ��~�<Y���Zx$��e�T�8���c�z�<ybꃭ=�|4�4���3�\h:pK�y�<�5+^,^�e��H�'z��mQ�<A���Q����vS�貏�y2�F QP\�TE�s����7�yR���4=�B�K7iKt����yR)��������BА�$�yb��T+�������l����,�y�IH�#��z��3B9�Q��y�ˈ'5^*��SH̞~�S2#Q%�yB�(l�Z���
�v��B�K��y�oE�K$* sbbȀsU��*�(�yB% $��g�[�d��P"�\2�y2���#r�'��^J>���ʰ�y�*����;�&�X��MJAl�;�y����u�Y�.�^Úɀ�8�yR!�/;�L�ŇG%$i�EC�S��y2��y.�pU�P����	�yblJXN��%�K
}��E�V��0�y҇ɥ"�@M�W�#Q��AFn�y��@�L����V�cX��e�� �y��V�eH�� A�{,����C���y�AW�f������T/"O�*W�@4�y0+��P`�G޺N_�����۴�y�h"D��I�J%S3��V=�y­V#� �熑�w�`�֩N�y�E�#�Uk��S3{9Bs�.I9�yR	O�C�F�h�j�1d(��OT�yr�=P��I��V�p�:-���y�$ӳ@F�����J=k�((�`l�y
� PT�@�ķ+z��w��<m�Q�"O4-�%*�=C-�8� 9	����q"OPXC�I@".tӥ�&C8=�"O��B�hÍ,24�S#�_= ���"O\�{%� E��BU�{:�c�"O��9�F�!��@�ԫɜ&@`�P"O,u:@GmF��Q�� �R�W"Or�����y AC��q "O��X���ET�y3OO#a�<!�&"O���Ak��M��x�T"Oh��ƶK�t|��ns(�$"O]�բ��(8�8��~�B�C"O�rFZ�#m����#�?�J�'"Om"���#A�Ĝ��2���a"O����E��z��c��7�p�G"OtlX/B1�d��VD��N�ڠ"OxѨ��]�:��ac¤ڊCŢt�"O��%Å.W�ܳ�Z�>��AY�"O<�+fO	���p;�q����"O���P�h[��T�J�r"O��c��U�躳S��a"O%��F#TNl��RGQ.n���"O:���˘�l\,Q���T;�E�"O��0��$�+���(/:Xk"O0��͞+���#�c	�&��9�W"O�Apѕ2

|C�bأ܀y��"O�C �K��x����	��=�V"Op\��T]�N=�cN�;�d%�"OX}�'D""�����*9�D��F"O2U���~�t9�U�7:b}�"O��r��۫tg��*q7���"O���5I�6N�x�8rj��f3(I� "O�P��
��3b�[�b0�D W"O�t�[�K��WL��ah�"OQ�%E�h1��K�i>l@R"O���bCI�Yu"!L9��$`�"O�|S�霡cw��a� `�<�"O�A����%���׏iX�Xf"O ����WC1��0�xR.��f"O��xk��FHִ�.2-AVH�"O���*L�I�J,S�D�/ƖJ�"O։	�˛Fn�)�j�A�� K�"Opi!��J�0������;~L�*O�|z�H��>(��x�����'J�-3b$�"F����&>6�\��'�rP P.ޯy��q#ǁj����'�ЙS����J3�څ-�Bpz�'+��hEk�-B@m���S�#V\�S�'G	6�[tE���7eO�L�zu��'�t"2���c�Dx����`EB
�'�{T��(\�Z��G�,ʤ�	�'���x�X�P8{R��%t-)	�'X�
v(O�HȺ��E'a���'.�M�Bl�g�Ȁ�Vƍ�'���Y�'�8�ӶL��Q��\���2K����'�.���l���,��
� K����'�q%�֣=�:A;�l�8F����	�'v��ZpK��*��u
��7��uA	�'�Όp0*�+v��PQ��#8A�9�	�'dd)d	ʿ$�]�G̜6����'xXtCp!V�&Ar��A�C.����'���&b��);d�y1#A:9[N@��'�2� �$��yq`2,5��'��`A�hC�\\<��w|�[��� �()�g�k��!K���w2��+�"O�`�V&�XL�\:s���8��y"O�p��(�@0S�
9m̙�%"O��*`b�7� ��bBS�[�4|��"O�	"�/��<�qS@�]�8x�"O, q�H!\��tᆮ�7��,{�"O�s��1�*ś�M�$I��+�"OJQ8t��`�
�EـW��g"O�U�p��~��+��@ܪ0A"O�BAU�B�&���w�t�"7"O �£�B)U�Z�!�@�)9!���T"O���oS"Eԅ��B581TU��"O��`��|�j�IP��<G7�s�"OX��#ћ��ęү�]1t1j�"Ofe+%n�l���Ӗ�H�!�X�:�"O�e��J��))Gl��U}��"OBl
Aƀ� 9ǪK�CF�@"O���M�7@����=u	:���"O�xK�.!+�~az#�ƴ�J�T"OV8��.ȵ�& j5ID�X���"�"O̕���J�B'��A6(ۚ[T1��"O~�Z��P�vbVT��^�/P���"O�U)V�צc#�a��3ڮ8	�"Op�BG��j��p�J�Z.p�"O��aD��7}����	��7+��ӵ"OҀ��� �B�N�.d��(���m�!�$�O_P�7#��P=~=�caW�/�!�D� I� �0��T<��Câ�^�!��sfh�d?!ܥ��]4&�!�;<��m�HW3#fRT/�6�!�$*L����'�Z�x�.�"e�!��X�.�N�JrE��)�U.X�s�!�$y��P�Ö)hn� B��n�!��߿� ��L�O[��"�mU�7!�D�#Кm
�C�;_H��,��H6!�I�B�Ah`��%Er�rha!"O4d���!?ԡ��dT-O�f){"O,��C��$�Qm�=��iA�"O�dAf���E�k>��;4"O� ��(�?>C��E�^�F�^!"O�%��,D50�w$���Lf"O�b�k�`��(���D��eJ�"OlL���δ-��!ab��,�0!�W"OL	㐢�3rD���aVJg^T`g"O�M��A�>{G�ȶfA>S�5�T"O�\�nQ ![pXz��ő;ޔ\�a"O�U�Q߽J>5��`2\�
]rT"O�8b���/�\����/�" +f"O�@hda�9 �� ��3#�.|�e"O��Ãn	�t,��V�~�#"O�!!�G)>Ԩ"E��S����"O8� ��:m&�xaμE�X4SV"O��+bE�i�б6����Z2"O ��f��3PB�QBȚ�r��y��"Ov�bpT0��I��&ߑ7���(t"O~t*��1�u�d:E�A�t"Ody1��$B�`5���C�B~����C1�����$Ûq�����l\�'J(1�5�W�Tk��Y��ѐ$��)�'lV ��(}t�ZǈA"]�j�'�����B�K�:[6��cآls	�'{rm�'��'H��q��'Lz���'�F��[)k���I�@�X�<Xc�'�Y�qkI� ����1O8x��'��r��_/�a��(N�.4�	��� eQ�	�A�|-�3G�c`���"O<��6hD�Pc����DƘT�p1��"O���d�Q�*]�%[
�I��"O�yh�H�6*	4p��bʪK�Ds7"OT��A�7>$ ���0 C �c""O@%�3��Ig�Ke��!\	#"Oƥ�T":H_��I�nP^��L##"O
x���!0\ ���?3皐��"O�lZ�B@�J��9��P0@P"Ojk�M|�,	�G�A��R1�Q"O�(yƯفO� h�(ě"v�d"OHL�凥%C�	�p%D�nr@YR2"On���
�#i!rQ�c�.p�B-x�"O���vjQ�@	�Ƌ[�i�l<J�"O�����$D����JVQ�h�s"O�i��_�p%ޘi�tr�(�a"O4L��&�P%X��a�ѱ"O^�`��>�4�� ߎ�J��4"O��4E�67�̴��'�&y,�IP"O`�IPF͌VB-�B@�4t���"O�����W�1����f�Nf�cv"O>t��ϑ�^q&�V�J�\T�YA"O<E9�Dϴd�(5q�%Bt��"OT�ó,Q�n���	�*ƀ7��t�F"O�l@@�E�/Tt���o׏F�䙉B"O�$��
̆���cW.��I3T�"O,�Ku�1X��D'�ȋt�!6"O�*C"Q�z5S�#
j��xV"O|��3�غ/�YX'c�P�D�"O,T��oXn�B�O��.0����"O�ظ�j̜OiDz�앝8θ`X2"O@ �����d��T�7|h\ȹ�"O��oM�p�p�xG�K�~.͠�"O�L�h͟<�]�2��}@<�V"OD��d˽_�>M�4%ݛ0��!"Ob�"�G\\y24J�K3�M¥"O�`�oA�N������
�/�*b"OXd�	�((�̹�Ě� i�"O����(ĉ~���`��	�x8:�"O��y"i�W�P�Ad�f�(�"O�Z4��563�lJҬ�*r��Y"OԽW]�������A)-5�Q�`"O��1Т3��D��k�/z#�,V"O`o̜gܬ�r%�8b@
�'|\U{4�n���S/h��8R�=D���
  P2�!�NA��P�&D�вtiM�S���+����E�B!�K�ML��"F & �i���?:�!�DZ�n��!�K	O{ܼ�����
�!�D@�_�-A��>CN��� K�!��Z�pQp��� "_���]!�\��
�҆EӘhL�pH�#Ұ%0!�]9!6�S%�[�$��cN��!�DO-i��05*�6���L�j\!�Ĝh3�#��	T�֕��'b�!�J�&��A��i��uچQ+��&�!�<7Z�	���c��-��-Ҭs�!�F@�v�0�J�C��X��ʉ.�!�$��&\�}䏵`���Wԓe�!򤇴i����0kܓo�$X��C0C�!�dH�C94H��J	�4�$pR2��4�!�ǃw� ��OJP����#@�a�!�5]A� Kt�\5,u�c�\$ !��؀JB��IQd�pR�ܪ&B
V!�� �@���C�`��[��F>���"O*���cD;P�f���DL�8���Y�"O��*u�ص,��,R �^�}�B�J�"OR�!��¸s��j��̃4Θ�t"O����fx`��G�(��"O�a�c:P���2s���(a*2"O��s�&�5r��$H���*_����"O�t�5��O����C�&y���	�"O����دx�:�R���LߴY�a"OL�q��T�N���B��W��]��"Ob�s�I�r���Vk�#�P�;�"O�m{Gl����i�N)q��"O�m�p�Y�Sk��舯{��`s"O"�{�HA6x�Ȑp𨈶}be�"Oʴ�q�S-VU�p��h��G��u��"O�l��iʮf��Vo�i�ȨK�"OXz�Ɖ5##Z!��D�<��T��"O!�uh�E�z)C7��,&�� R "O&1��@�i{�Ir�ޕt�
�#�"O����@� �����/�j��G"O�a!����%m^X�~T�!���y"
�7U|�Z3���LG�@)���yrlTOC0��q��?B�#�l��y"i�� xQZ��x�Aࢍ\��yR��r0N ���ؖ�4ĺ�cS��yr���v��r/.��aa����y�HP9w��"p�ݺ�m����ybB2R��4�E�`IFa�֦���y�-
�5s|I�CH.��RGD^�y�g�����Z>�V���`U1�y���<��AZ�� 0����g�%�y�F�t��7c���]zG@��yBo_�3��L#�(	�d`����y¢�6jm@��#@h+m�?�y�q�`���d~��I 	���y�\}60�PTmؾR�0�X��W��yݓ �,��O�����I��y"n�pl��ץ���\��!��y"f��t� ]
P�[�����y��4$.R��p#I?R�@�e��.�y2����qc��-6Fz�a0�ͥ�y�$	�GmbX�`� r ��ƃ�yrB�%L| �3d�a�F	02A�6�y��7�6i�C$�.�~���dN�yb�#����(�Z廄��y�M.>��ܩ4��,}p�h��в�y,V���UV�ǉ|���v���y��]À�z�I��zh��!@_��y$�#%Br�B灕4}db�QT�S�yR�� )�Ջ]�tu0lqN۫�y"�D�EUN1�����l�r {�LC!�yb��8NT�ʐM�8
�j����y��E�-���0u�'��X�u���y�b�JV��:�]��M�a���y-���-�f@G�\��M�Pc���yC�.��x3DU f����q/��y�*�!L�y4CZ(BlX�"�y��34��=��eV-��hbk��y�a��
jȬ�E�%��5�1
��y�������3��-{�ES��Ī�y�N�p��,£Ѷ&:���N��y���<������/$�@@��E��y��H�4�,�D�3Y��۴�
�y�ÜSm��z��BQ*�d��ԏ�y
� NX+�@^b�EY��C�W��ag"OL	�!l��`�e�;e��"O�U�m�7y��A��U'���z'"O�����8n�d`��z�Jh�D"OV���%[(����<�~�A�"O��fM�d������ܓ:ႌb%"O�Q�&.ԊA�i�D�Ȍb|j��d"OZ,����llP�Q�O�l{�Lӑ"O��V�4�
i� ŗy`�Ч"O�E��(��'
L��F�Ľg^R�i7"O��`֕��
s�L$tA�E"Oj1�S�HƶI�B��'�楀7"O<D��o�_p,���$�R���"Oh�:��
7:����+��&�T��q"O�E�,ȉ3��!� ��gh�<Q ��SB�K�wq&�1-�U�<� ��!d� 9�dNU��ʣ!�z�<�g�V0T��I7�J'��H�O�^�<��C��B���BĹ��-@���u�<�DL� ~���q-�s�f�K��w�<�"MT�(��a��6_�h��!�s�<ƤG�v��01��ĝ2�b��v�RO�<��C�'�\(��lћy�&�Y�f�b�<ɥMI�K
�rc��yȍ���a�<�˒/�a��Ĝ�r`���`Ez�<)��
[1��ȷ��%AE��h�P�<����&=�0@��^7-G��)l�<�'n��P�c��M�����b+\d�<�gBI1$7��d�1�@~�<��
ʹt���@/�2V��9EF}�<�5�F�b ��J;Q~�}���_C�<٦l�5I�X�
s�^�;]RT���\�<��Q�Q,�:��6j+"UZPƀr�<�t���X��B�~x�9*q�p�<�p�_�l ����L�|�d����p�<���$H��4�x ���O�<�"
T&x�@�)˔g�H��1�AH�<���^1��T�O�	7��E�<3�T�y8�
��+J+|!��m�<Y���3�v$�󀔧W�tiugQq�<�k�=2Z��x��֦5. � �B�<��ҸY�_��ъ�-S!�R��p�[�(�6��d�!1�!�d߉n6u�(�1?��()FC�z!��+� ��+��1"���!�䄧-��m�P���d�VE[`݆�!�DC�3�L�p�$�$����RkM�v�!��Qj����|�R�
��`�!�DD-)���	�%�;l}�Q��˅�t�!�䐏@�:]:ħ�z�*�۴�i!�ݼ'k�0˥/�4\��	�^!�d�L�\�z��W>O��'h��iw!�$��`���!C���K�8��G!�b�N��c�N<$�r�����!��P.RNA���`�>9���Q"W�!�D*n��40�³B��(��K�1�!��	K��0���&��2��Y,!�D	��UBOO�=~�Ҷ��0aQ؆�`6�|R�gQ�`�i2��
�/�q�ȓx�����i3.�"���iʴc�t@�ȓ2�4�xB`ؚdB��r	��@5�T�=���U�:��ȥE�"�V$P�XD�	�ED����Ŏ�TFȘ�g�S$0 ,C�I�Z!���=�����k߆.�B�k����",#��U����)B��C�)� �↪�� �٨g�71[��T"O���S���Lzl��L� L�&���"Oh��uA 	�^��j�8��1A"OB�'΍�C[�0�HV�E|�,�`"ORPs#L԰j�Ux`%�/o$E±"O���S_	Z��r��/P(���"O��J��U*U�����@\�s�"O*ł�o��$4�՛`��8?`�$T"O�Q��cZ�;�n����=��["O Lٴ��z^��A*��a�"O��!�M��tj�pxS �-7)ˁ"O(ݢ�k�U�8�	�Ć�h����`"O t6`�YNPurACFP���Yb"Or)h���0/��z4l�-=�|ɣ"O��h%��(u�Q{6J� j2VU�"O$U;�l�+zر��	{OHqq"O�)����G�Tex'ۺH���
�"O�A2CL^:R�z`զ�|����"O2傦"�%,�����Ț�͹R"O�@�G�`3� �c�z��x9"O^퐡(��[>�<��a��$��E"Or��ߞMP�հs!�m{<(�&"O�\��gU�O��IPa]�q�"O�����@>`���EH;V�Q�"O��`�K�fFxa�ԭxi�"Oj1�tn��|>����Z,8�j��"O�eK�۾�|`cԁF�:\����"O�q
5��'�����J�S����"O���QI<*�K�.݄kEL�!"O$ek��H�5j,� X�!5fl�B"O Ac��>B��1D��2�T�A�"O����9;�$
43
�0
�"O� IEئBY^���I^�,��H��"O.�[��M��=ļpI�b���y�G�I
����
k��!2#R2�y�Í�~G�08QI��WuH�;t�[��yO�%~\x)P1�٘U���b޼�yA�$^
uj�'Z1!7z�c��X��yBi����@p�G�����݅�y�,7mЀ�w��.֬J�*Ş�yG�7<�4���%D�@��D����y2N�*ʝ�a��xX��p͚�yBc��b7J�0f�>h+*��DT��y��:&;���3g�"hg&��2���ybJ�	.�X���E�i�=�!Ő��ybfC7[�����c����TA���y�`�#���P[�XiDGř�y�lF&���֥$DN�� �y�Į%�X
bJ�1��K�m��yğ�@�B'��zO򄲠��y�L��C��C�*��X�jC��y"�D�}E�X$!3D١�M��y��F��$�#C{B�Qs�ݝ�yB���OB�t����d�&��rc��y"�Z�Y���K�_���0ׇ�6�y�n K��rSI1
�с ���y�R%,(}%\Y�NTH��y/.���%甃D�бi�dV:�yB�O\��A�.5�����y�a� T��<��׻�	���'�yR���q�V�'(B��`/��y�Ɓ
g�DA�� C��sS�� �yJ��r}�x�%hˉ$�!ө��yB�L�ix�b�A��i"F��G���y
� 2fbQjĶ����b���*�"O�Ӷ�
;��ؓ�i\�Ec��7"O��J@ω|3��Q���^Wv��Q"O���"ШQ�!'ULp�Rg"O���Q�Q"��|q���2�!8�"O,���UCF&=E��xG"O��;E��F�0;�'M^N�Ip"O�Ps�գ7��8�͜;:Rr���"O������+�:Q)�ˇ)8!�ɀ�"O>�b��"䬽���w�<H�"O�p��31\,��$-ܽ&����"O����R�,t|}Є��5<Kp`)p"OqHl�.�X-�lѯK`8QS"ODp �M�.\\��m��I���"O�4pV�_�e�h����6-��d��"O�U��%
?N�<��8,�,�b�"O����,�|�\Ű�eV�>d$��"O���v$�q�(���@�Qa>t2p"OP
3��#��Ғ�:@�.]��"O
����v6�9�(+Fd�5��"O�d�cm��v'� A0$E3�"Ov���X0P<`���FC(&�@�	�"O�R���O(D���Ъr��`x�"O∻�@;�,ܸ�$G�~���"O��+��ɸ�ƹ1�E�"��`"O�4�M���ʼ��ޖJ��)V"O�IHW�ݘ0�x�*$J�,��"Of rP�n�nCqK��
#"əL�!�$�7�<kת� ZC&qrc��W�!�T����rrÍ^��`��@��H!��H�L����^tҔ��4��Bf!�DR� �ȸ��k�3s�z�Y�C�
U!��Xꎘ FA�~��TÞ�{�!�dǔb áB� e��H+��-�!򄖄<��a�C�u��U5hJr�!�DE:??����;�̈Q� �C�!��(?�H"b��:GY� χ5k!�d�0ov!�/�RYz�9�M� 	 !��T7e�^�i��\M�#R�T�t�!��O_B��ҍ��E:�dz��[(
�!�D�9����~�V!����9�!��F�u=>z�J����uKΜur!����T��F	-��ۥ�th!򤅯\lVz6��;,��;�b�- dџLF�D��Ya8��ڽ.�8 :��	�y��߱F��8��N�'#��	�Y���=�S�O	�y�/��Z�</yB�(���U�<Q��Ԥ+�)�]�cN��(� �I�<I�͇%#ެz �?NG1Z��|�<�1��5~)�g�W:,;�\�£YT�<Y0�G;z�J�nȳ af}�EKUL�<��B�6� �G��q>�"�J�E�<����J�^� �ߑUͰ��.��<y!O�j[,q{�fӎ{�N�Ac��P�<�Ƨ�"%A��ym@�b�X����A�<9�,S6<Qp�S���ĸʢk?T��x$���F�j���_G�L�&�4D�`A���'�� Y%N�-����$D��eMO1#�z��5��VB���f?D�`�Dn�ʺ���^�2A��GL�y� ͮ_��s����)9�I fg���yR��]� [�
A�O^<�uN��y"�q6fmf���Ҙ`��X2�y�O�������Ǧmҙ� Y��y
� �l��G�
�B`z䯗w�a�c"OQc�Θ_��e�С��ps@��"O`����/`�h��\d� �#"O��u��!*�=;5"��,���"O��Su��v$jq�8t,	�$"OꐸS�M RJ�.I���G"O����꒔'�����O/�p�hp"O��#��Y�br��Q�	T`�Z`#"O�PI3Ϝ�+����*��H1"OxP�e�	{��ѡ��-�0 ��"OYb1I��i�b ��C
-���a"O�]�b��A�8��d�9H�H�P"O��+����ɡ��y���"O̩��	��ę�)ھI�P3"O,ܡ0�"J^V��d���8�	�ȓ~,9ru�]b��Y��� BD8��ȓ'DDɠ�]�r�	bbHK2�T}�ȓy2��J�"$,�e��aI=|>|`��0�|BFfܽq��I`��#j;���?|z4y�|&�Q��̡Gx<0��$b���nT�~ն���7",C�I.)�ڭx�Ȋ"�n�
w!���C�	�z����1x�QaejW�:�2B�	�(&�	z��3"��[��1h�B�I�sC�h@�#QkLl��,ι0لB�ɛ	���Y��E�6���L&c�rB�I�:��1!���b\t�`�^�`B�	/q��8�A�8HQB$]6nP4B�I�d��ԧ�=��D��*V�.mB�I0� y��Z�)�C�ӚdSB�,+J$ GX7@#(Y��DD� ƸC�I�֦=��\4� ��ӈW.�@B�	�Xi
���Y�L�H���
��C䉖f|��I1.K�$� �TS!S�C�	>Z�Њ�N� �p
 �/o�nC� L{��� �,�)b�l�B�>C�I((S��FjY���#���	C�	�;�~-�`���B�K/K�|xIUj0D�$���?t�(���U�b�2b"D��i4�)�H��Bն4���:�g>D�T��Ð"[�9�����教f�:D��z�J� �F5���02�S�J:D�4��@<���Sm?.����=D��P% F��Q
�C�@:�ݙ3O:D���P
��(�&��s_��JN8D�ˆ�H�eؖ�\��%W��q�!�d�?�^�򆅀%K���a��Qz!�$D�755��o:My֍�"��#_y!��B�����_�b�PI��Ѱfr!��V
� $Z�UY�[���R�!�d۫$<z����3NPt9�Iʩ9f!�$�HQz�p�KgC�d2cE�!��ZN���q��P��$�4b!�D�12�!b'b�"�T��`S�!�$�:M�6�A�_�5}.9p��ɷ�!����0�c�Ā�?f�@!�mWR!�d��:�4�@g�����*M!��;�8�S�1y�ZIE��@!��Z+v�^U�1b� ��	$K>L!��F*hh��C]�B�|�A)�:`@!�D�V�d3�M�*���(��L�6�!��Y�|q��P�$):�X�xǦ�q�!��D6!�>����u�B#^?n�!�dм&��=���� ���E��!�� ,p�0HϞ��Ib�
�M��"O2 Z%���T�h��i�- ��L*�"O  �稏 k�����/;qֱ�s"O�]y�ϕ�~��Y�TW%<���{q"O�� ˖4��ɠ�A6}���"O `un��9<�hH!@p�(��"O�� w���&����-4�@Q�"O��K#	�=��(X��9@��*"O�=�%KUIo�0(&,8�Z8��"O�Q0'�C��Y���=AF�26"O�Y#����b�1��	�Z���"O� �G�C�+M���`kW���"O�QHBK�5x.>�2�ֺ���+�'� h!��=̮�c@jQ�M��$
�'C6��2f�0V\��E�%r����
�'��e���0Ӕب�	n.lu��'R�·h�/`WС(���UVYB�'",���8aԤ�p�X�]���
�'[hJ���7v���W�J���	�'��sS�ٔa���
ފ!:l,�	�'j��Y0OĄuŚ�4%E"1jb(��'6�0Z��<T�UaM�*��j	�'���+עț"����0 �yѰ���'7�(Ԁ#Z��i����>�@]��'m�  ���;N/T;���1�.�!�'Z�=��sB�0��ǭ_t6���'����(۷�(!Aw���]���i	�'��]�4̞0c�|522j�'��	�'���]9TށHp�K51���'��H�'&'�r��ԠJ G��@��J8B�0��Ձg�hfG�&O���ȓ��yCt����8��Q�Ӽ/\���	���+�������`Zfч��%�մ����.O�5�("��.D�(����)�����ߪU���p�+D�Hcp�R� [�1R�ʟF�����(D�4�P��.C�U�D+HY�x�Y`�8D����I%(��fB1=p���&8D��9�0nh�
�C:'(N����:D��F�J��P.B�n�"WB�y2�2r|"V��y�ڕcq���y2�ȨV�p����k�.�C҉���y� ��#��^ذ���� 9�y��
�:�,��&J�Qb*\��A��yF.��prr�6.�������y����?'�x�#�'U��Q���y�-ɋZ��� �K�$m�������yB�\�
"0`�D�O��q���J��y��Ì'�(�ʳ��KF�W��y"���(*z%٠NB3����E����y�邀k��u�Dު�P��t/R�y��	+�8(ǈ�t�|�9C`�"�y⏌(�T�E"d&�5;#lJ3�yrDO�����%�L(�ڨ����yb���ک��G��h��k �y"��n�DHel)^�oΐ�yr^n�(�Cǅ�[���u ���y�nC�O䒙���D�W,4yR�i�
�y��ǌw�@2ȶfBa�$ ��y®1V�ic��ɒ,d����F1�y��'���;��A"4�&Đ=�yb�
��4�D��5Z�"D�#���y/��lA(M�F��*V&���$D'�y��5d��%X�ʊ�F�ܬ��y
� �qIb�D%"&A "��/J�}:�"O�$�a�o��@�c�L?�|H�"O ��C���`5뀟j� �"O޽{�Έ6��RG��*Z�sQ"OTt
�&�� �Q� I?:�X�H�"OTЂ��� ��G���83"O�� $"U�ѣ��
�����4*O����|q.	�6�'G�Ņʓ
����"�T��as j�|2����;~�u#F>W|]S�Jևy$����L����,H~D1�&E�n����ȓ��H���
P���QdJ5�@ �ȓt��jR�	M��§�* 6݆�-�^�r��++\����P�i4���%4�8���
"�v1���F����ȓ�űUf���� ��)_�j��ȓUR�= ���m�-���� 0H�%��
w���F�G�v�Rԙw�͢iv0�ȓ7{�x �Ė4LL�2@h�%)-�ȓD���V(؄n`�(� ��0$ǔ�ȓI�� "�B%!	
��V@J�ZX���ȓ[P�A @i��L):\ 5"ˠT*�(����U�Sd��u�2�A�['�C�	&���7D�%#�/ʺ"�B�I+nU7m�?[���v�2D� B�	�a,�)5N�^K�dB�o�2&��C䉒)ԘY��#=�H���C(\׌C�I�T��`�6��=03h����(B䉪l�]�׬R�in+��\fC䉒7�:0�g��#��|���-%�2C�ɔ�L\��#��v��p+b ףii4C�	�.����$1u�ՠ�9~�B�Ɏ{+��0���J AȢ��|	�B�ɱw�R0i'�N5/�� �t���>	2C�ɘwz��F�	�}��x4�S'�,C䉢��Q0�әP#���%
P�s�B�I'r�(��[� �8ٻ�C5��B��
�uR�-؉R�ūeN�8��B䉈t�
�Іl��	�!���J�=�C��Dڢ\��%JF�@�:<�B�ɵK��d)��L 7�``B�&�^�B�	?���"R���H�B�3���/��C�	�!p�h�X @E �
�V�<f�B�	�*<��Zs�	�1{#�"\�C�	�&��)�2͂�`��I�`$Ji�C�	:���s3�
���kt�G�E��C�	�[[�e+���M�n}�Ѐ�:�C䉂k^J��UbŝP�4� nO�	y�B�I>�������Zɘ(�x8(C�	1UgTY8�o�x.���iџ(C�I�[��e�	U@F�O�
ZBC�	d�f@�&��䔋�c�>�^B�I'��%����e]�D�w�7Z�:B�I�wX���#�Z�S�t���l��B�	:6-Ʊ�Q�؎N�����M�|��C�I�h��ԇ�$���j�˸+�0C�	>(:h��+Y�O�&-�Ǫۄ*�,C䉭z���_�y�N�ϗU��B��;F�����q,�3�	Y�
�B�I<e�L9[2��0]|:��wn�9W�xB��}�|��Ȗ 9vi(��Y?_ZB�	�pϺ3P�T% ���B�016.B�	�9�`|a��H�z�J���#�yB䉐 �<d��	�6����͘�[�LC�)� nQ��X�7Z"�Q����^L��k""Oj�b���4X�y�*U&Y�"Of]��,Vs�P�4�Z�7��h�"Ohd���l����C� ;�P�k�"O��;��ٖBw@}UH^�%~���"Ohw'܏A(T$��ʱ)�$�0"O|كFc�4,�����g��F�zc�"O 0q ,��)�B,���+3����"OD�K_)=�4�*L/�|}zp��k�<�G�_��>�`H۲�ІP�<���Ń�&��Q��+^F	�'�ZJ�<�#	 ;p��	"DǱE��uB��JD�<���D$b��c��\�C��E�<�"���&Ȉ���$�_I�<y�	�����H�h��Q���L�<�&&YC`@0�b��1����^�<1w�4=!��#N�E�>�2��Y�<��I�0{�.�a�� ;Oh��S,�S�<)�$��/��arÈ�#���OH�<��a�u��z�A�)s9d�CuɘA�<�chZ�"o8���O�bѪ��k�G�<Q�ԉg����y� %��Νi�<	5�R6~9��/��l^`41P��h�<aC���h���c�Cz�����Cd�<���ŘY�B�t�����+�!�]�<��υ�	N�`ai�
��lk��]�<y'��#F��Ur�O��T�A�a�]�<	���tX��rc� ��0�U�X�<	3��!szl��gD:z*�$��*HZ�<q'K�X�krmM�,<��`�RA�<q��W�s�����G���R��/�S�<a։Y�;�R4��K!{BL��EN�<)��JYa��l882^�r'��K�<�ǭ m)A	Y��X5���b�<A��7(��2Յ�3t�<,�&��I�<)�m�*8�Z�A�0p'jt��AWH�<!SFT�q�9ҰDF�:��#�k�<i�ǚ.M�����BD��ŏg�<��I:u`y�J�K�,�B�_c�<IT�KD ���'wo^���nK�<9d#�-�H0���, PI�KF�<q�r��T��c^�S����q��z�<��i播S�-\�x%R	t�z�<�p�Nk�B83�H��jM��&�y�<s͖�Rt`j����EJ��D,�a�<���$� 	볍ϐ�����a�<��T�l��4��ǔ� g�F�<!Cl��S�$p��GD	w��]p��Ww�<)�b�P|\h��,F w �#GNO�<a��̢o*(I�Vm��c�����lL�<T��<rt�����<e|��"�a�<YE��	[��C������:�"O��3�/� U܌<���%v�2�Pa"O��>'�8��K�c�����"O9�7�#v@�S�K�4G�V,��"O�#�d��2C��Ht�Dg�e��"OD��Rǈ/ >�HAB(�Nꎠ�"O�,k�� .�`|��gZ6�R��C"OzEJR�� h]�PӅƇ-:�H �""O�a�����5�,�^�<���"O��b7A�6�2Evሯ=u�2F"OpتE��*S5j�`��֗]l*u3�"O�k���#T�0�ΦR�,��"O�R�l�(�8<��F�8��r�"O�  �sf�]u��ńܲ@*�Đ�"O���Ӯ��$�����Q�,9� "Od50D��4>���	������4"O�((4�R:S�r�m�?wـ&"OT|a��p��i�1�W
���:��	ӟ�0rnV2=�&�'�d^?Y��
VE���m۴8����䏀r�0��?��@���A�\s��7��RtQ`�.��༂��M6��ɦ]2R��-8R���(Or��Q��-V�fS�b�-����
�Is`W6�8 ��oM�:U�LhӁڀ�� �{r-���?�C�iY�� 6�:'9 T��˜hAZU"g�7�����?��?�����w���)ɰ"�4 2A�Σ�^Tr�D���lw�7-m4p0�� A4	F�ID	M���eC�ilߟ4��L���eB�'��X�W3d�hU�
�m�:y����&`�	 vD�g%��U	��e��8`Aᗊ`3�x���|r�'�5���OFQ���`Lƨ��
��M3�.��Ra�A+ŐB��ȇ/�B�����A����mE�a��x)�$X*k}�$�C��ড�6��Oxo�3>�韚#|n2�>� �y�@�a�*_�u������\�?!���'"��:S�L�Z��A� �$�V�DygӘ o��$�ٴ�?Y���u�k������G�߅6�$��&b�4�d�O�q��
�+Lx���OH�D�O����?�޴V��	 ���%Dn0�n;b�� 6
��,�B� r�˳G�z1cdh֕V���X�#n�
O>i��4
v��҆!}�8P[C Э,DJA�0��	#�,3vOά%k�]�O���P�j�ɿt�PA��%S l]4��ud�&�n�/�P�	�M���	Y}��^�<��E���V�I�<k�)�&θ'V�	�ۨ��=��G>@-dsҹ ȆQ�I[!�M+Ǹi��LcӺ�4���)�|��A�HQ\���ާ��D�㮈�+.���F�?����?���nu������?q�g�(�U�B�V	8E��(�I"�i��JM-ҠY�%=\�\���'���r qGĀA�'��Y5�5d��H{@���A��A�h���IG-5�֝r��<�l�u��C*�O*UZ�'�H�#I�/|@ �6f��t81C�'"A�6-�O�˓�?��*��)(���	U ��б眳T|r�'+�EH<�uՉ�8�Z&�5k���A` �d?� Ѳ	=�FT��)�n���D�O��[=X���e��o)������q:��m�N��'\�2b����X/XKl�s�#X�4��UJ�
	\h-!�ƝD(T�r�ɂ�/�(Ov ��ښu) @ ��L(�.����\�-�P�PL�v@˃
��}�0��!˪:U��`QU��O��l�M�����_{���D)��;����Eۮ}��0��p��h��Ξ<R���IܕN )�WIC�p>y��i��6-~���r�H������ϘB��E�O6ыQ�צ��I��0�O}�(���'6��i�~�s�
43�ȽPQ`�=
łf�U�}�x��1�Ж'%�|�`��5h�^I��D���˧�z]c��
�͛"Yh%A�lG�/�8S�4y�dPPƆ�4<By��㏊^�N�PF�	 T�bI~��W�dAȖ��8��9��h�:�XoZ,	���DW���,O���s�2L��㕬]蠁@��H��*��O���2�Op<آ�� ~�,�!��$�� ��I��M���i��'\��������d-��y��>5�H���I�Ir؞谥   ����"O�Xud�tGz]+d`�X	��"OT9+�OW1u���#E'Y![��1�c"O���JF v�*Q��	��t"O��y��+.���T�F�fj��ڵ"O�Ͳ���
,�lkկ�( u�zv"O��˒É7�,l2�d�	Z��` "OL�b����%.����#��8"OJ��Ɏ7Q*�y�m�l��$�"O=�!�;|H�U0�6؂"OX;4�V����4��P�B�[�<���P�ŏѩ? VL���s�<�Dᗿj`i�%�%4�H���L�<�f��Q&���Î$)n��{7�J�<����,w���K���	z�{�,�K�<��D-<�$�Qk$a<����H�<�6�>�v�:u\���`�s��C�<�Vm9g���h�ńzZ���&n{�<Q1�R3E�=�Dm�6��I�R�P`�<���ÖQ7�����Ѭy���c�<Im�6#�\)Џ�?R�"��5�R�<�碄$pz
h�
����0���T}�<�%�;�$��P�ڂ4S�I8S�|�<���%}�b�P'���Rl�R���`�<!@�U�E�K:M1��W�<AKѕU7l�ZT�DKTlq��Q�<1���&ϰ��a=�(���V(�B�
re�4:�ޟF/ؔ�Ae[�ɒB�ɼm�<���%[I�^�mM�7D���̓�Q2HX��!�2g�$��9D�\��X�<�v,J6$9�lj�4D���Wg�Iq�P������Ra�0D���r��*Nx�)WnZ!8���3D����JF�40ǂ�=c��!�0D�袂���L�:Сp�ʍ����TG4D�� e�E)NXt�r֩�/�֭x�)/D�<W�2o�P�ƞ
R�ތ�q�-D���d��l"y�B!�	=���;�c-D�\��	�		Ð�[����<��HH1D�t�D -Bc�0Rcl��ǜ]㓌0D��9U-5GH`Bn	�d��A��N)D���#�˾FP�QV=.*�B�(D��)V O�}�а�7ȝ"��٩�@(D�`���:<i:����׸" ��R�"D��l������@T,\��"D�� 6ݨ��:H�^U�D�/�t��"Of��@N�	j�ف�ߓ@P!Y�"Oj�j�Ky9���bZ�'���w"O2�['��=h�N������P��"O�XA�96a�(Bi��F��d p"O =��iI��*Lc`��0e�#"O���3cO�)�&�ڵ��E�����"O0�)�����x@sNG6lԸ�C"O��D��+JA@"0΍S��"O�9!¬�2u�t�-)a>y"On�	��ʆ1�T���#p[X�"O^� v�K'�4Ѡ/ۛ(����"O,:�<R@�hC/#  ��"O0��A���}��h)���;i�*�'��0���xьaФ'[
3+��2�'�.��߃X��6��o��t�""O��B�������I�4����""Oj����Q� �ؕ'�L��\ð"O��KY%^�*�p�fޭ&ŚUZ7"On�����Ŧ�:�K �� F?D�Di���|� ����˲L���Я)D�T�o�.^Ru�p%
)���H�(D�Գ���/|�h
��h��m�$)D���@�ӵFrԨ�7�]�UF��0*)D��:� �� �/����CC,D�l�3�7��A+�Y4@���*D���g.�k��0d#j���h��)D��c4$C$f^$���,WM����-D���wb�>n }S�<~l�w�+D�����A�6�ܔzw��(��')D���!�i�^h{�ϹM9�H�M;D���'eX�mq��PgL-D ~Y��l'D���Al5��d�0!L#z�\�ja)D���6C���gU�S���" �:D��puBʡ
Ƞ��r�](9feY�	4D�D���/u߂�q���LI��`1D��(w��)��p"�1��Zh<9$%N�zL��c�c�*�qf�A�<� �Т5�d�7oD4C�̈H��<�S�*a��9�独
�B�"�B�<���*|��Q���d �CSx�<a��";Ŗd��㓒Y^
�h2�s�<��е_��� #ߐ�TL�N@U�<��["E~�̳gǁʆY�c�ϩ�y2&�>E���[c=�	�Ӣ]:�y⡈��u1c��%]|�1S/U3�y���  '�"��f�"�y��ߓZ���Q��4�d}r�CF��y�KЃ����T��r�!bd�yB�X |������΂\˝��ybE�Bh�������!�F<�y2����ը�%pZ���n��y���7�|���V�2��XӂZ,�y�a3TY��{��
=��K��y"�X�q��A�� P:&�ǣ�-�y��WƬ��ȷr;4�d=�yB�R�GҔ�T�R�\�8:�,�9�'T��2Ľnah��
v�z���'H���n.�f���ہtb0�
�'���#�K�n��5
s��;f[��9�'�pI�dG�-Ru���P��iX�'%^��&��M�'�(Nq��j�'m
]�aŭU���z�uT�Y�
�'�n(0����0y�c��m������ @�E�X7{��u�'��]�Z�k�"Oq�ǢI����Wʐ%a�Px"B"OtD!��
;I�����8��C�"O��@%�]�H���JA�9��#5"O��2'�6�z88eJ4|�z��P"O$�h_$s���{�	A
U-��B�"OZP��ϒW�hҁ�v��Q�"O$���KC���� 8g�H "O�����_�D
]���as("O��P�j�=�P�I�
�s��{�"O��K��a0A1���S
��"O�m���(V�HM+�`C ;d�0 �"O���1�900��5"��$d2�"O8-ENK_�����\�:��#T"O�	YF�*�da����\��!��"O�x[�&��u}\!p�a��$}�p"O��ǒ�/$�YU
�jZ��#"O�Iq��O�q�@99CJ�%W�8�"Ot����+VFEɌ8f,̘�"O��j6:���)��b��w"O��2em�8Kᰈ���A>o�H�Ba"O�����	n�$��g�����pb"O�`%[�T�T؄�TZ78�e"O�B`L\l�� �@�]aޤ�"O�"Pe
���T�!@שq�!V"O�1bN�#D�=!r�J��@�"O�i�0A�;7�У�T��q��"O��PՄ�D!l��+\�$��"O��7�7栴j�j\��"O�b���{���t�T5{(A�@"O|b�ڊ\�(��n��Y	 ��7"O�,XE'��*������ѳS�4��d"O�McQa� ��1yPFN��\��T"O,�C�K�+�rH��_�V�|��"O�T EE�^Uh�9R/��+߲y3�"O�a���~��t:EOc�C�"O~ �K�.j��s�mK�x�"Or|�`�"T0�Zg��I-Е�'"O���U�D�B�BH3�ɖ*tdYF"O�d�l��eD�ӵK݊.:p��"O 혁EMFg>(�"
�O��2�"O��j�ɕ�G7�B5HH*`NV��"O�)��׆�h貇��Ѽ9b3"O�1Vꑽhd�	0&��}� ��w"O8H)���/�*f��ht�Q�"Ox,	HH�d.`�YV�U�i��#"O���#�6HD��R2.VWҨze"OD(��/$=�bM:�/وKK���"OJ!H�gǱ�e�b�+6��Bw"OTQ��W%*YB�O!�еcb"O�y�m,UxE�R��z�P<r�"O:�j��g���i�� }ݔ�ۣ"O�z& ��F͌y���Yڒ��`"O�p{3�\<8�����V�� b"O��A-Ķ7��a�P�H�m�ԕ�"O�5j#b߁r}��b��o��d��*O����j0HV�@[��ЌZ߬4��'nE�$J;$3b��M��Q��m��'��1��ƺc(h���1�2@�'?L`����-)��� R"���'�vQ{�̑�/ƹc�9�`e�
�'�N�!��
�p�Ҡ��	��;	�'>��AٖpJ��'K���,��'o%�5E�5WN= g
������� ��Jp��B��M���=p��`��"O�q�K	-T[
!	�^�(mpE�	r�O�Xd��ݱmk<�@�	�&C���'�i[%�R�P
hБn6
��|�
�'��T���_6i/h��RE}��a
�'@:��tI 1���"{~�T	�'̾h���`%��A����\��'�`�!��LK+ԃ?��x���<!�bZ
ߜ���H�$��x��LXt�<���݃Y��� ԃہ~
��D�K�<1�.)rK�aa��V�YpzD ��m�<1�Ɂo��`d%ϺD�$�h���A�<�N	�T�<Y�p��:-�D����x�<��-[3ZJ��^@�0��BKl�<�d�Ĵ��՘c��Ds�hr�<1�JJ)|�t��%<RE��v�<Q�Ĕ�3�.���f+F��X�'v�<1w�:5d����
��m�6D�u�<��lWT�H��i�h��|"�X[�<�e
Ǘ2�V0`�::d��5or�<0��-Wk��`E@�#�xaw"Pk�<��,Tk��A��Q��F��Ch�f�<�2��#V�  #�+߮}�d@��M�<٥M�_�|��i�w<�2��H�<����{�xRR�Y�\����"!��X�E.�³%O4qע���/y�!���4��y�@�F��@RΙ�|�!�D�
F�$"w�T��sA��
�!�d��=zx��ʁ<`�8 ��T� �!��P	�E�B�,M�LA�f��9DF!�DW"d���%���դ��C[�PK
�'ֆ�!D��uu����L�*��@�	�'�<b�ĐSXd�9�.�4<��'��Ө��^M�m�����;����' ��Z�
�3�V���R$Fa����'�����S�r�ђ��7^T��'��8�
F�[|Й ��0���'\�q��m(4n�w*��"O��v-Ct����m���<��"O 4�"�Od��Y��U�E�R��4"O�`��1R��Tу ��` "Ol��U:�X`� !��q�T�0"Od|�a՜H뀘؂Ե[�̩C�"O6�H�ؔ*z�0�M�3;�ɪ�"O�:��,>r$���M*#0��T"O\=�n#a-�)��`ֶm6`���"O.YpC�=T��0/ئ��"OR����;&Ţx�G�A-,_x!	d"OZ08��N�W����M*^ȸ#"O�,Ƈ�C:(�Q,�&u{4��"O��"�GӣC���E��'](��"O�=�w�<5��iE%,B���"O5���Q:0�9�C�P׸�"O�=4�DF	 1S�Sn��"O��j�4aU�av�N9m����"Ol���I��c��Wϣr{�A�"OVU ��^_���� [�Gf�I�p"O���Ƭ��<�R�kv*˧oX�} �"Oz�"hU{�B�A2)�3#)2�{p"OL���K:'�� eM3��S"O��[EOK:; �i�ˤp�|�"O��)D�֒}���uָ����"OJ1����K���R09^�)6"O�5�K=U����+ߚ:<�`"O� �����1B���"e���-HD"O�+a�̧%����2cˀU�XP��"O@�+"  YDX]����z�,{"OLy��]��1���)s��<��"O�lh��R�s��4[v���S$��!%"O&QG�Ŕ9Q��hoB;�>���"O������,;�Ј:�,�!��L�q"O2�;$	Y�[5|���f����"O�cfJZ�T�>�q���	g���ҕ"O ��+Q2z�ܨs#ġd��$8�"ODq�Da8IK�Lӄ��!\w �2�"OLC��ۧ}����E�=|T�a�"O����4N漉D�]E8V"O�e:FkڍI���M�r����"O�L���%J>@�eΑ�L|�"O�<xe9#`��rvM�&O!� �"O��H�脔"m�tӢK7���5"O��9�j�V�iq�� g��<��"O�,"qE��j�2���L@A"O�=+ˌ5����蕈i��0:�"O����+�!,-va���;�@�p�"O��t�U?Lg2�{BD��,����"O�@�Q��WEN�'�6��U*Ot�:u��<-e@�x"�_9^��hq�'�8P$
�I��@e�$cޜ{
�'����Fk�/;��a�� E�Ճ�'�Vp�sOM>T�d���7�v��''�@��F��X�����(�&ˮ� �'������6XC��)R$��u�t��'�@ۗ ������rF���'��iC�֪��P�b �\�Ґ�
�'�dP���ՎY�Z���,�?�Ĭ��'�8m:֯������a3��@��'y<�0�J5H�˖�tlE��'h�[��^�x������e7���'VKWih�a���)z"٪��w�<����I��|����@�x"%M�u�<��diI�U����h�I��>рC�ɰ�@�E9U߬)k!��>^:B䉌<\Ԙ�r�gdx*�G�Y��C�IoW����f�2&h�#U��-/��C䉧��j�l.G@��j�mΦC�In�p��Q�^�>"4���φ�m�dB�ɯr��q�c˚0:Z�0��Șn�`B䉪R8�E$,x�,҃k��lB�t@��� C/t�v@�gَ�>B䉄*�r�$bXE�d,SW.ת]�LB�I)i�����Q�<���S6v� C�I�s��9!�J��M��ԩ�폷n�B�ɯ`(A2� 0�U&N���)�'R%AoبE�b#[�K��i0�'��Hfh?"�IR/�Sʀ	�'i�
VF�� n��p���+G�T ��'+&�ٗ��_�6� G�='X�'�$���M-V�)K��( �<x�
�'�����.�l���7m��Be��'�x�4hpdqWO9Ԟm�
�'2�Rp�ω@$��6��%US!�
�'+.l��1Iz�)���2T%���
�'�����	������⢜�St�9i�'�$�2f�&��B�e�D_X=��'6���G-�  �.�C�EѪ:���`�'{hq��ET�H���A�O�$3	@�k�'d �K��	g8|Y�"t-�	��� �y��U�M�*E12��.�0�14"Oع2+�v'��� ��Zw4��4"O��t%��sب�q'�= [�Q�A"OnM���9?܂1��ϊF��Hv"O~�)���Z�����+c���h"OhQ`cEF�!fUZ���!���"O�X�ӏ�m����	݋AX,q�"O$���+Xo�v$YFSK�ܳ�"O&��b(�I�
�C�	�@-��w"O�xze�G�f�&����N**����"OTL��W�9�>�s4ǐ�#ȳ�"O����NLRyq��T�E�`t8�"O1Y�
�� ��Y�WĜ�W�D��e"On����ʖ �LT`".Y7iTl�9�"Ol�a�H.QLZ�"M�?7h�@2"Od�6!�69 ��c �Z"*��"O01�w��*W�\ )��0d�"Oj��Q'W�6ܾ���	^�H����"Ob �@��TB�8+��G'j�,U�"OH�G섕K����Y59ӄ$��"Oh`��@�99�q��K��eX�"O
�/,���O�(%���D�N� !�&zz.�b�����G	I11�!�D=V |=Q��'̌i��2_�!�\�T��!+% ��)`���!�$�4�fݢ�eu�����Ԑt�!�dH�[~�"�
��2���K��^�!��
"p�L	Ԩ�4]� M�2$SGs!�PU��i"��0  ��26l!�d�/�8$��O*:�`(�#E�6N!�X�&Č�g���u ��Ce��!�d��c!(���4vv>�B�&��am!򤏅�����9L����� $O!�P_����U�A�5�����/c!�Ą�XQQ�E�n��V
�l�!�٥!���Q��S�,��P��Î}�!�-t�>������!������TQ!�DT�=g������k�
�r�bكkD!�ė�0;�x�ޢ!���p�⛙r%!�ė�[j5 �aL���`j�A�"!�P�D��cN�L�8P�C�ų~�!�d� #<q�aIɨ=i�T%/]3p�!�D�&0��A�	f<@�p$���!��e�� "���$*�P	"�i�!�
GX�	�� T�_�z}�$��\�!�D@v��D�U����A���!�d��IXP�Ke�˔�`S@���!�$χ6��y�`�(�����{�!��N"C=�1���w�H��#AK�!�dHD��1�p�Q,$m� �r�!�D�R����J�3g� �J�o�5G�Ii��H��܂�BR���qM��t��u"O0��#J#.w�|��H���)�C� |O���"A�w������$w%�U@��'o2��ט0�����J	�p�C� c+!�T.@��@����>0:���O܍*џ�G��N�<7��"P�D� ���W�Ԙ�y�E͠K�����$	%�qP����y��]�@�.i!&�F)��0&a�)�y��H�v�P5�#�{�bM����y��D�$`T�)���?t���*5���y`;h��6+J�oܖ��B<�yBk�18��E��fc��z�c^e�<Y�i@S��X�2�۬RZR��h�<� >%	�ƈn ��Y�ʉ	h���"O6@hTL��o�Y����.j�}p�"O�aG�Pg�d�"�][��3t"OZ�P�a��I~N5��(S3C�T��"O`�aM��ld�����T�K#�ܸ"O���R�G�_^��rq,I-%(x��"O&E�b�
 �D82�0�X���"O�T(7��7aǴ���D�2y���"O쨛�Ҁ[-�h�$��+��!"OtsV"�s�,xK1����`b"Opa�5l�{�ά���ȚW ��JB"Op(q�Ζ�~��њ��4��	�"O�g*�cU]	T44�S"O�T�dÙ!tT8�<z<�@t"Oz����D��p��J�:��1�"OL�k��ɒ$�ҠR�"�%g�@"O��"��.�	��B2`�T�#�"Ot�"�)Ëo�s��3�Z���"O^J��ĄR��]�R�]�	�̵��"O���Z�3@aä˳K�r���"O��ա�n!DI��Â"O���b#��n�:�##˖j�b1�5"Ol=؂bC�9�)�c��_p|ٰ�"OƩ��G$t��a����)e��٤"O\���[�$���Sl]�@cn����'{�D��-��u���	�i�ܬP��v!�$���9���� �&��3�ǁ^��x2鉀dU�uQu��14�h��B��C�	*����b�B��3� B��B�ɡ}�x!Z$@��O7���� �o��B�ɲ+����M�A��8RJQ�w�˓t�	;
�5[.�km��)!j��ū��/g�a��I���$�SZ|�9 �O�!�f�,!��_�P�fP�FNO"��$��X�v�� �j6�"�n�x�eI�2�^`b'=-s��ȓ�()�̋ [;\��7ϒTGx�M7���}"rC@���&G�LX�9�B�Op�<1���FN
a�&������l�<A��3<��*!��#5�8�J&�Ve؟0�[L&� �� 09
���Mа+�2Ԅȓ�0��`����)�2^͢��ȓt��= ��Ó9�H��:)5����#d�ҡʋ�/g�\���PJEʒf�<�'���d�E�F�@_J�B��^J�<yU�ќ[d�\8B'ؑa��( o�M�<1�Ř�x������6@�Lģ+0!�d�\Єk��n�[�Ć�=-!�$;�|�p��;k�,�b�.�/4!�Ù���Ӧ 6j�f$0 ��!�TQt�k�i�K
6U���Q�!�$ͼ1�`�3���.=�\+�n�9l�!�>�`��,��P�-��0�!�$޷IB~���R�U��ɖ�!�D�H� U�EGp���З�n�!�$�]'���Db�1�X�T�!��g����#���<�7CٌZ�!�Ć_ 5�b�όz���\>hD��w���{�lWN �K��@|���ȓx��T�1H,��H���óvA͆�TVz�!�(� 5��i�O߸P;f̆ȓ2]��r&K�2�q���+7�хȓK���w�T88�b�CL���!8��[��ޡu��Y��%�~�؝��k���xq��O&+��4�d���S�? 0aI�R�-�.U�G�	���lJ�"O��f]�r�d��C��\`�"O	�B�e�����§��`B�"O��{�D��~�~���-ǊMݾUE"Or���B�0�h��
F�=�
�u"O�x�?D��7HÇz�R홤"OL�8v�K�-f�k�ˍ(t�Řf"ORXQ�B�5���aE��Ch����"O���F�I�b�֬��䎲@W�Y�"OrD+�ͻag���dK�t�Ȉ�"OցH�Q�T��@58��-�"O�@�EO0��ѓÓ^�ܴk�"O�%��K�(da�T�$B�Mr�Ib�"O��u��mW<}KB#I*	r� ��"O���N�)�D�	��
S����"O��bS�'Q6�!�J�@����'"O�L���TO>�عtE)j��hw"O�x��		P���	PM��B"O�)��� WF�Y��#��t��1�"O�$hT���0��hӭS�"�rF"O|��׎؁#ɤQcօX�y`��"O�! u�֝�4DIF�Z5E�e��"OND`t�J���!H*aP~�""OZ� j�~%�������"O�z��8%1�Y�z�Ve��"OPUZq��*oH�չ��&���8""OH}��.��&F���@��	�x82"Oh�S�l��Lk��A�I
nX4"O�����==�ȊA G>0�X��'�����jJ��E�r h���'�ᨠ�Θ0Y�K8u�����'����0$A%k��}�̉D��Y��'�(@;4h�'!�RM�F �r@�'�t{p%j��#S��Q��'�z�����p�P`�fŪM�B���'v�$x��?��q��S�	��'#z��A4�t��'-@m�
�'& 9�A�O�\�xEć>2�9:
�'����g�Ǎh�|uj�Mngn�2�'d�SFQ���-� D�;  �	�'�F9����46T��IQ4��'H�r��F�GV�!�JC�};��Y�'�v�1/��g�P1��I�n="���'��m�4��Ipn�W36I[�'~�,�p"�	5�<�`X�I�����'c�BPnڰ--�a\3�?����?Y��ni���O�Fѝe�pj2'܇06��DJ0LL�I���)~�aЃ'	6xȴ���f��<��Q�
�'�`|��s��B �)I��MX��K�!�r�x�)�#�\7������z��K>Y3e��i�2/d<�$sd��g}���?q��if�O���ON�I�H`*ʅ`��L;��"�I}X���`I��P���ǪM\B�r  ��r���D{���Od���j˓=��I:�I)#�I��!j�X���J�A������?Y��?9�
)�?a��?���!h��r�G_3{�R�����I1�<��-*����ط*����D�c��Gyr�@�.`����*�")�P�qsD��Oz�|�W
�/�����!4���?G\~�Gy���?�?�ߴ(�IcQf� j��A�o5:R�X`�8��Or��5��|z�\����@�"�5���!O�G?y��)�';jF]J���ə�˳7�r-�i��zӚʓg��`��i%2�'��S�+�����߼[�4���>?lE&��?���?y���g���Rlr�b����G�G�	r��|��A@1g�:��I���5mL���d͘���q2剠*�$��щ����)�n�RN� Vh��qT��V2[xM�"ňָ'��`��<3�V�#�hӼ�ӆ�ܞ*ɶ�C��*6��=������?!��?q�����w^@�(�%�e�Q�O�Ibʙ��@��V q�@7-Ը�\00�B95$pD���	N]��Ҷ#_��mZ���Ik�������'����[�����iSV��4s��I 1�Ɇ�B���ei�IB��VL	Q�l��O�|r���5�`K0J��k'�EO��Cc �MC$�O�I��	��(Dn"PK��Y��HZ4�ZW��� �l97Yps����۱��(Cb�i� k��R�V�x}�������J���p�sET�9�iagV��~�'��Of�d<���M��ʧ��� ��F��>|��<��i��7m�OoZݟ���溋�*ide!Η�4�N ��b�'����O�=�B�'	��'
$�]���n�50$��z�eQC��(�l��sl��z0D�2l)��b�5�&���Ե�r�@܊1C8q$��&�G�HF(�*ԗ>�8i�����^�>���FΏk�܍��i��,���\��!�D��7޲(�֩�1m�����;R�	4O%|���Ϧ�����>�L��1�� �@����T���$ x�O��0�׋���)cCm
-D��`"��Ԧa�۴�?��iw�O��TQ>�����"����͋�j�ީ�$��:&�T,������	џ���9_>�i�OJ�D�vY&}c
[	T�X �P��#�ڱ���F��2���3�U9��А'�H��	�JPx3�(u�	oV��$)-s����gb�e�����@��y��r�ĸ��'�r���F�f��%`ֆg5<����[9W�F��T��/,���'�蟌�?Q��T	�q&��<�&�#֌�i�� S"O ���K��f�������%=���a�O&xo���MS�2�'��'W TQ� ��;����Ճ�O�Mn���M��-����)|�6��?�����X��	�R���4�� 3���BH��s�V�����?9�!��0�+K�J�(U�w�E�1�| R���&�"�"���.�VcW<8nQ0�)��FQ��A�b��o�✘�E�'�Q�E5r����C�f�>�+s��38��ԑ=�@���5�I�|�J������4�?ᬟ���CH�=�jѸ���\7("1o�(�?!���w��d��C�
D�
�◈��2�\p�y%�6�`��6�\�!���ǅ�)|!x$��VqO��;��*��j�� �   �?(�b�"OЩ8�O�.*�kӊͳi]�ة�"O8�v�³+>.9�4
�h]�I�C"OD����I�����AAاVBt�+V"Oh@�gYG*��c ��<P�p"OH�hF�h�
YQ�N�'���PU"O&=X��\-}b^Lҕm��O|�43%"O����gۯ=ʐ �0b��;j�9�7"O�u�"$DqH@(ӡ�VNZ�"OP,���v���*qF�v6h�"OT�eE71D��d�ڒ$Q�=S�"O��w�"|}h�C�	M\�8�"O����ϋ,\���۳#@�FG4ɠ4"O��%@%66����#��wc�d*�"O4�����JȠ��C�<3+���"OƩ ��[��u�d̙�"'�"�"OL�cj�.2�`�v���V9J�"Or�9T�A5�񘆊٢H�h�b"O@u
�@�l�ૢ��+\��`��"O0�k��*m�p��NV�&�<�`"O(�Ht��mS:X$-�3j��ycd*Ov҂��#Ɩc���a�+̣�y�̐v�����EԍZ���kǑ��yc�/h��kQ�ξ#�.��%R,�y�!6.��z@��%h]��v���OB���X�Hԫ�4�?q������n�e!�4�a"�i�@�X�Cug�ԟ��I��|�f� c�y(3��t��
3��r��}
�!"W��
#���?�8Y�(�oz^�<���9	84	� 
D$��(�HSV����c
�&��8�dJ3<�������dz�<�`�ʟ(Zڴv�O��&l�*Z%��Q�?A���cU�$���$ �)�}��̿�xI�*�/9���c��	��p>���i�6l� �	�EۺNMH)�3��8Sv ���O<�P���ߦ%��ӟԕO�4����'��i��q����g������(Z��Eϓ^T�pyFhƈ8�D�D�6^�>Q ��Pʸ�'���;���-%<1�Uc
 7;����i�>D��@<U���(�I�t��!`n��]'���}��~�4�J�h\h�hI�`��l��R	���OJD��*��i�$���"QZ��`s!�% �.UY�'�R�'׸��2�\���˝�GoT�P���u�t�<���i�7�>��Ϻ�%X�"�6��B.�7�29��ѾY,��'��y��$�/6��'���'�"ם��XlZ�4���r�,�d@@Pk�А\i���3�M�&�m�q{�4]=B���O���.#O�'��9;��ߍ'넩�ݗ?�N���R�*m��ո;9�)ٳ����I�A�a��lŅ�򄀈�$e���	I��k@	?|.��4M����@�aiJ<���?!�O�E��gQ�Ik��H�̵�����Fyr�'�������K�n�S�Ȑ�rW�D�v�O#w8H�k�4 �֕|��O��$Q�|���]O�L�sr-��O�~�+��ָ�셻rn����	���I�L�����8;���� /�.���E%)���E㆙�jl��f�%0=����ŠgZnH�3h+ʓ�h�K�d־ I@�r!J9i�V�吣v�-H���q��ů�hP��c$f^�'��L�R*�8*�L�zаi��?Nذ�`��+���'�b�'3�O��'WR.e�REa0�ӆ�3���Dy"�'�a1���?햙�QM�-�p�`��O��l)�M+�^�F�E) 0V6-�O�d�OW����I%ʉ�
�W ���H���O��d�Ob�3���v��AH�nǦ>c�ֳ0d�x�B�`�� #W��'��-EQ��ã� T�$��:#X	f�@�57HH�.�&1h�"�g����'@�S�
�<e�P�sش �q�� lP��L!�L�w�.hh^�؄�O8���C
��w���~�R���:]����'�
"?qU�i�l7-t�jA��D�"�L`*�A�3r���D����M��
C��՟��I�?�Q��������������S�>���,��'���F��eM��IЎP����鐕_~QF^���,���I�� �ƂC5]��[��6Viݴ*������b��Ӗ��!���C3��^��xL~��!D��A���f�~ݸ�[�&%nڨs7�����ٴ�?����iK0��DH�Y[R��`f(Ɇ��'jR��/ғ}ŐqB.�)&9���Nķ(Yt�Eyb*eӚlo�x���?��b�,1x�H8l�l P��3Y�4�(�|��'��`�� ���P������9���	���OF�d$LU�D����O����OV�d�W�D�i�n�x'�+w
vP�'�ҤG�Ш�i�G6�
�g�w8hc���*�l�ɇ�Gy��d�|r�H����G�Pـ �4�/D���b!E `�} ��āx�Is���(� � [&��'�����Ϛ�s�2Q���LB!�H�O��0W�O�nZ�6d��<������Ə$iٙS�WsX�)[嬞+}�铨�>�s�'Y�xt����(C6��7>�H7��˦�%�����?u�>Qu�� >  �!���X�|��$x�"O��8S�
�:���IY,!�����>9���)�NIJ���(�0/�u�vT�(�!�$��m3b���D7/��uh�4�!��F 1|yC�ψ�b�X�Wܰ��IQ����`7(H?t)�ьG[�8RP"O�= ��� �@ r��Y䲠q5�2}B�ɯ5�4�B��no����C�fKLB�	�o4��J����т$B�'��"=�"Ƅ��f��Y�`�`�l1"�KZY�<! d��L|��AM�G&�y�
�y���=q�?xA�	1)	R��-� ��w�<�g��3Sx��#J�.ٱj�<鴤�\f����Y0�A
��L�'�ay�e�3:�|��TǕ(Y�IuV��y
� Jy�d�'pH���XE�� %"OT��O�#�\����B�!G���"O�@k�%�;,��TB�xL$���d-lO�u��G۪R�����kF�E��"O(���l*0V^+~i�$���Hp�<y��Ӣx�� �`F.wL�����YS�LE{B��1q�� ��![�Dı癹�y�h��0j��I�NP���2�*�y��)�'~�leǤ؃}ƾͣ�I�x����	Y�0�26�R N
@�F˔�bE�'?�}��8G���	��yMR����hOq�� x���9+jM����-��Q�"O6R�A=�0sWy{��pQ퉡 �?	8d�ϯq/�A`�L�J4��#$��cزY?Zͣ�!��H1��'�z��Ӊd���2��ܻH�>]�w�"�y�J�7 �PC�(�+Z,�!�F����0>arN�c�� "hL�a�K�hVC�	�0z��R`M,|�qk�X8c�.C�	Y�<�S@�Pw��IsH� �'Lў�?�h���!cv&��
�_�TS'�!D�Dؗ�̳;Gv��p$��h1h"D��cB��Z��kU�ƷY�Ei��>D���$+��Vg�����@�1���(D�|`���x �K	�^z�|���$D�H� ���D=�Mb �ˍb"���n'D�@�7�W��m�f�I�F�<��G$D���A ��Ux�G�E8d��a$I!D�����VL�Z���L��C��>D� cF�R9,�U�ʐ=ȘУ ;D��ф���C�tu��D��I�4Ӏ�-D�,�!iʴOpR��%g[4a9��rR%+D���g_����ʙ�Ot���)(D��2���?t2j�1���-4�JB��� ��a��i�l(ᴊ�?FB�u��W���R��Q�%ǐ:B�I+T���r@����]3G�59�B��J��b'��?�z]�+j�C䉅��-��#�5f�d��a�9�C��,|j�8�f�A����A�2��C��0�4л��B�Jf��p%R�)z�C䉅fj������8ȷ��(v��C�ɛ@�T3V��-�N�zR�߼6�!���*H��Pp��=yj���	�>P�!�dH �$�� �h���W�ܢ�!�0�أ�g0X�l����i�!�DL�C2i���:H$���G��f0!�d�3ҕ7��/I��4s�h��dF��ȓ?���;!�O�2i:�BQ-V�Z\��ʓ$j����أ6
.M��'��+HC��6?��̋�-ފ"d,Q��d� <�rB�5N]�%{��5<��0��.�F�XB䉏?@��c͗i[�\��j�~�6B�	�L��}
s�?J�x�v"ȫ0> B��zZ��C��9��yc�AD�r�C䉟���c�ɰa�x-��K�Nm�C��W׎�I�/�l�
H���d��C䉥&j�h�G'�S�!��=$(^C�	�P�|�!()���rD��	#DC�ɉO�M�i�~!.�@�b[e�0C�	�Izjmʳ��x� \�ƍ�$>PC�ɀ1|Z�+�8K/B �c,ז�HC�ɭ(�v����H#��Út C�I�g�\��ԞH^�#v)W0y��B�)� ti�����5���j0�	~�H1"O�D0��҉h,ʬ��$�99f��g"OX(!E|�EPd���b-��"O�0i�&݂�)�4��93!�l�"OLT�,@(QXX�I�!H>E~L�s"O2�S�h�/���0&!F��p�"O,�s�Ɛs:Q��j�*�$�"O"U����Ko���*к# �p"OZ��5�њ(�"|�V��"Fq�"O�h�w/őx�8�[!(d�q�7"O�(⥃��'ϰ5h6��9��Xa�"O�`q�Ī#Y�lrU���u�jr�"OLY�Ǯ
�ؕ�tBS9`w�Ti�"Od%2/��)&���Ƈ�@n>�X"O���n�$ �Pǃ�yUx�	s"O�lavMD4fCpP����/)�f}��"Ot�36�
�:��� �a����q�"O,=E��:3�>��Tf��<���"O�e9҅�/#%��&�{W����"OX�W�����ecq�ɥ�� ��"O���%�ѭ ��a�v�?o.�K�"Ob:`A	�X8����ؘ]&�ib�"O\��p��,Z>4QJD��J�"OdpCE1c^M!�	܋�<��"O��F��A�	���+BN=�5"Op�1��Ҕx5�ǤC2h����"OFШ��	h=�H�L.4�FU��"O��ЦQ!r���S挚�b�t!��"O~1�5F�6'�.����+p�l��w"O`qk�넁3�����ؼ��2u"O��Ш��S�J]�b�B�j�Zi�"Os(�^2���q�P�_����"O�8K���y���fA�4�B�"O���H�M0�jA�.�E��"O����6ih���U��"O�,Zg����A��@��"Ol�t��!����Q�ÇJ$�1B�"O���m0w*E[A� �X����"O^=�wd
�x�R���!5�^,r�"OPM)�f�-h�*�蘌/?F\�v"OX5��b�4ĥ�`Y9L�挩"O"�s��nc,)�VP#;��q� "O��?ɱg�J	Lꦀ@���y�+�O�6��C��Aͮtc7�
�yB�Єn=�L�W��#����"�y��	VipM�C��!vA�y��>�BЁ+�T��d	�yR�6W�z�%Z���!{�@�y�σH*u(q��������B��y���K��%�U┐+k�Yi�!�<�y�hK=/@��B/�0הp�SAW�y�e%e@~��N�%YP�(c��yR�&~�>9�ᧇ(!I,D��.���yB�' �D��(Ф%�
a�'G%�y"�N32��۱g�0T9�R�y2�Ybɴ)[fo�|sr g�\�yR��<a��!�S�f.Lq9���y2�4[M
(�@�t	X����S�yR�W�����J�<1fa��2�y⏐4��e��F�� 8����y2'��m[Dc���" �H�� ��y� �|�R@Y��	#��M��ǵ�y�� b��	RE�p�@�� &�yrn�4#�B�b�1k�m���G/�y
� <ey��Q4Qj�[��s���(�"O\,� �ȟB�X�T��_�\��t"O.!KD!�e���a��Y��"O�9c�0T�(��� 
'�:-��"O�5�a��,�1{���4��� "O�적	F����-S+ӠI8'"O��f��#$-��þd��H��"O�t	�-bB���G���K�"O��a ������d]���p�"OБ"��1�ش�%W0},�Z�"OV��+��Tjܨwf]���I "Ozٷ!,�l�T坲!��<�"O=;���%5�H�#VcH�08���$"O\�f�٪��Y+���Hb��"O�
�͕:_YHDrWL-
l�؆"O���
��'����v	ܓc���y'"O� /�9q 0��ww��"O �HVGس~�Ft0���gZ�K$"O`����H�i���U�<rUI�'"O��H�|:����FзOTFds�"OP	s�G��٪0�u��>>T9!"O�!R�"�YJ��cVC�p��"O������
�jѠ�����9�"O����èc������`���S�"O���IKfX遮ӈ�2Y�3"O6КĨٝb����7��.�B�xw"O���NG 9PؑS5��%�0y�"O~}�N�#S���9wJ�+���"O���D���T�RD_�;�4�b"O�@��^�n�����D ,D��@2"O�eh`	�6���v�J�V�H�K"O�hHA�'0,��T	߆�\M�7���G{��鋝2�J�H��-L�|$j�'�*B�!�A.�l|��l��(`�p&Tk!��'pM��8Ή2o6]s�d�Ga!�䉟��As��K
�Hha��E�!�dR���;v�)bO�P��k��>���?�H~
�.\-F�X�"m�f��"��<5���a}����z�jD{�FA�<P-	�����=��ab��}�<yPN��CbL�րS�r����&WN�<���ĲDu@�{���1�V�L�<�##�<R�b|��@[=���S�"�]�<�-%y bI�==`�|;jMY�<���(L��@��:�H0k�+YS�<��/؀58���8LN��CAe�<6	h����VND�Bk�1���	^�<I��W>V��!a��g��I���\�<I�n�43�ٳ� :G�j\��GD<��f�jEiG�	��d[a�J0c�M�ȓ��5Ȕ$�&[P-Qf H�(��I� Q�qNX�T�d�`��Ck���ȓ�rX��t�*5X��ǎ�RM�� u�f�ݜL�08�4�M(���<~�=�U����sΉ�}���ȓ�	�SjA&d1��w���f��L���t�'��$Pd�q�0X�dǔS����{��'OLD	W��	9�HP�#	��`�F%��'�5rɟ�D�$k��,U��xJ�'}ޤ �a\;y��KR}�Px	�'��ӄ�Ԕf!p����z�4	�'E�p��M,uL��3BɆp�5S�'g0��ĈP�X����-eX���|�4�<Qq��`D�5���S^���� ��s�ҾI���K����"��h��$8�S���.3��! @�Y�Z%�D�>�!�D�,�aif�M�w
�e1��0���-S�'��>�ɰ&�P)��� o�%Q�h�+rC�I$k�J��΅�y���ڂ%�'?"�6-7�S��M��V8���n�,.��̒&�\Z�<�lԝY@p��é{Jd8�O�<y6J�k<f���@&Cz x�I�<9Č�. ���I����z�3�cE�<`N�;%�`T�B�գPP~��NUg�<	ve��\AVM����r��h��Sb�<9�� "�ktC��n��a��d�<Y1��Q�F�ʅ)F����C�e�<y0��o��lh�G�9�,�z#K�V�<��)�����J\?dd�	�baU�<1%/�D&6�;Ө�������S�<����w��2u2|����BL�<��h��Jhb�bW�-m~\����]�<I�g6cN`Ys�''�YK�,\�<�B�X��d��g݉G�,53⨘U�<q��Z3wG�@4'_�T�<c6�Zl�<Qe��P�V�	Gk҃|����Hk�<isnU�\��m�����$Kх�N�<q$+O(<00�q�[@Em#+�G�<�dkD4'ЮL��mFrUfP`e�X�<Ir%��r����`�]�$���e�Q�<��D>T�:���;yhH����Wx�<9�gڎ�Z�����xu��U��B�	�PT�	�`I�u�|��	�	?!�$�K�4y���`ޤ����ޙG+!��1�^ �JّŊ�r���82�!򤏗JURѫDj��� ���:UF!�M|��Y�Bەz?ڡ�.�'#\!��	W��h�e�$U3&�kA힒\�!��^��D�#�@�>&=�f�P�!�f���˔?S�\��F�*'�!�$B�o^��V���{4�\(7���!�$ܦ8���#�
��0���zDbZ�w�!��͏b:t�bfO,��q�aɆ�!�䁞��X����=�&�%�ޒl�!�W*+x��e)��E���Ȃ�;jy!�$�%����9�����8v!�ך$5����`6Z�ȩ��]�h!�d��O��0�!�ڦ	};A;(:!��~���H�=t������( !�[�Se��[g��n���EЯF�!��×#����Uh�"t6�,��*��+�!�$רp�ha��m��3v����,N�!�S�#pL��b�=BM{S��8c!�$�#h�*)�R'�%6 �!U��P�!�
,��A��T�MD�Jf�	Su!�dӗ�h���m%dd�ؑ�R`!��T���b$O�;T�=��M2!�$��j�<�`�~�e+��ϻ�!�} q���j��ьL:I!�D��:�b8S3lNN9��*f?!�dX�[� �2����M<v��D��l�!�D��cZA�d�ӯB�xmc@�T�b�!�Ds��a#�����`�%ɎE�!�R�Y����!�%�`5���>l�!�d �n<
@����-��ٮN�!�p
�� N��r�8#��	�!��8�N=��	En�P�25�L:Z�!�dڡHn�������Rd�;WA��{�!�� ��B#�%A���c�d-2��"O�P�uŃH�T��-H�-/"��b"ONԃ&B-f
䢦�W�z�,��"O�,�񤄸v�0Ec�	ױm]j�	C"O����q6�����N����"O��"�_�R��
dwpR"OZ���� C/�hS����Z�ac"O��Q��G��0Ս�::����"O�I�2 �|[4%)�&��f�nըc"O`1��Шq���(q@��I��=�%"O�M�dK�y��ӣ�8M�"��"OF���!8f{���'��*=���"O���A�N�03ѡ5{���)�"O]���7�z<iW��?2�֘ �"Ol9�c���ZP�� �&��"O��Ȑl��t��A��b��``�"O���r�ԟ2�]p�	+���("OL��i��-N6D�V��
�\u:�"O�tK����K��J�Ea��A�"O
�4�a����֧M+��X&"O
�q��(O��1�C&�8���p"O�ph�p�5тD(W Tm1"O ���G�}^�=�v%�p%�"O=�)S�~�X�ĥ�6c�~P�t"OB���#Q�^��D��&��YC�"O,P���Z 8 ��%�٩�"O�ݣQ�ў�zYQ�AL%��U"O<)�!#@f$C���2���"O$�!ve�0�z�y�DJ��`6"O�)�rl[�mT*���L�fA��"O|!p4��=(�!�ߜm��SD"O*����Y�	�PLS��3Nac�"O�' iO�]R!����٥"O IC�@���0��]%[��Lb�"O
��I�m%�T��c�0�vU�"OLD�����0+�Ȱw#��\�8�@�"O�M��k�2{�03�ς&|����"O~E3A�8S�~��6-"yH�h�"OHs!Ā�l�H�ҡƺxr��B"O�D!�)T�.�*ÆȍC��5ʲ"OP$)w!^(���R"��JT�Q*O�q#�P'-(i�π<(�XYs�'�R�ʄ%��'����NލIj~H+�' p0��ٹUy�Q�I9:��a��'dQ��ES�|BB�����
?x&@��'�p��c��.��ܺ��K;�
u�'�.��BBX�ƌ�: (5"� x�'�2������i�
�X�	��g����'#Z�8���O��(�&B�#R��	�'�BA+�˖�`��)ֳ,�9I�'�0٢�=c��j�H��
ۆ	�'\���Q�>�M)�Nܬ���'��)#ǲs���XsFȃM�6���'��, �۳|{��h���vM��(�'׀٣���bk��R��LD���ě%1�U�q�'R������q�!��]�X�r,T�u�B[�5�!�D�$��\q��=i�J�J`�]�~�!�dݛ0*�+<�����I�59��B�ɒ5��h�e	�q��(���%Q�B�ɟ_l�aQ�)��'j��qC��s�B�I�w�\h�s��Ħ�RU�&B�	�-���C�H>'�p�#(Q>1czB�	j!<�	v#�8x����aCM��B�(L�B���b���������+�B�)� ���bfըhd���Ɩ	�|A�&"O@�3EF�|D.���h�z.��"O�+��[�Q��=Je�A? �X�'�����N�5i�!��R(.��`�'<P��5-x��AIAV�$�%�'
�����3���!���+��0��'ɪ�p�W�r�ph!�����P�'"�DC�-�E�`�
�X��Q�'z���mOn|�ZǦ�j��l�
�'�=���y���F Ɩl�P}�
�'>�l��M���P7n��T�	�'��ͣ`�_�`��iA��]��]��'>v̰�DY2:0���"I��!�'�h��H�#�x�3��"8p"٠�'��\Iu�< ��mc�
�� �<d��'dDp{���v��q+��|H}1�'��(�!@�a�t��!e�~�V=��O��*ec�:=�azbC[|��<� "!a�延D�%��>�g-	Jjd�ώ�Ed��QD[84�e�KAX�茆ēY��<"'
%;`6�W��]��0Gy�ˏ3X��,g�ڥ:b4�>a�oŒ~�������>S����N*D�\ s��!���Pc�խZU``�-�3Ĩ�0i�7�PͲu%f�"~�_�v=�U��/� Z� �o��,���<�Xsɕ�YY�� �*
2d�8�4i(��e�K�'^�pL &џP`dg3�Zi��eV�X�a"%|OD�A�K�5(Bp �ݹ8�yئ��Rcn\���2�0��s��?�� �H&l8k�� �E�L8X�fM|�еqc�d4��aLU
():I?�Ѳ��Y&��""�#9����(D��b`����ze�3����Eƫ ���ʖ>��I( .(^b�|��f�(�oҹ�4�
�/C�bHC�i&D�ȡ�L������P%N�Np�	ĝ������te�ԯ���J̱�,�Z�'��٩�kQ6����a�4{��ϓ���(��@���`0?+p4�c�9(j�hwυ�9¦�� Ƣ5�3��6�On����\\6�i�'�0׶�2��|�gY0Ӽ�z܀�FE�ZW$�Y�1Բ��OP�m;$fU`��H2%�Y�Z� �'%zlXAn�P���"B��-%��%:2b�0�iE��)'=�r�h\� '~h$?�B��\#�y��q����P�KJd  LH���x���� ��At� T��߬J�|(_C�`)���(\����$�A�"��Y ��	�[g(a�w���l���p��f����Đ�P��1s�1q�$Y�Ƌ��8�|��ą�e<f�3��B�L�x�]IV(C�C6�O�9���
0��- O:=�@�xBCYE�h:D���4+�DAD�F~d� �ȒL�>��a�XX� ������$��f��C�	�F�r�##������X��m+D#q4�:���|��1@6G�z�_#��𑷁X ��ݥ?��(Ґ\PDąUNB�_� ��^/(�ug�0w�nQ�T�贰�E��sw�F�0(Z�A�O=mJ�p��1t�`(��U����K������i��)Yu;�(�F�=ғ2�Z�H����v�����L�8B�qK3����Er¥�G9�DJ��8�z��٦#T�D@�� �A��]����V��?�t/��]i�AC#t�@}k�+C�N����O�> j�6� ���N�(��m1aaB�w�LiK��L��JVL��4����#�I�e
�"�f�b��P�'��)H�lËǐ��ʐ��r�p�+؀!�,�0���5���IW�6��1x��ÊŐ��
P��x�@�w�H��R�P��-S���(c�
�e%@�0��P�L4aڇ�Ò;�x��ע�왐����$�á\�v^v=��_�]g����C8�5(ge֡����U殟��Q�ѱC��I��+{�[p�?�OJ�w˜���5:]�:Љ��3-��˵·B���L�7k�UaBh�%�k� g�N%c�FM�c]�8ʦL��:Q�hf�I���5(�I�'�(}�B�4�J�1�O��&��T�pΓO'8q����x2	�%
�&e�T�ӑ0�\�qA�_3r����C&��z�ѫ�o�6cgh	�<f�������ͪ.����`pv�-QQ�Q*���Y�.�bj�z������.ˬ� GB�6�~����V�R�B+#��@냠��q�lZ
�>r�!gn	�#�N ���Q�X��ق1l�6��0)w�D���(ڮ�ڴKcu%HP�q�P[����Al�2��i��y�F��i
�`lC�&p�Z#���'�d�Sb��8���Y�J ���̆0%�T�A��$YP.�`�3� ��P�W/KE�EeR�k�� �S9�l��dAQ%ZU����,��<H]���P	�=�&�����q��-Vh�P ��l������^:DE���R���L����ȃ/z�z�)��������D�k�2���'�O|�)��D;0D 
Qd�EϔT�ReW��@��ţK�tlh��آ�\�r+z� 4����e���� ���UJ^�Dr0�բQ!YC��Y��',�U�KAV����
Vs�6�0��^�zTyVm��r_v� �*Vb�9j�!�fׄ�"�%W�p�<�(�f^ p@Q�-s\���X�Q��& c��3��A&0_�0�DFK�S��-��
NF��YG*Y�Nd�� UKY�VEb�Ĵ_a��2n�-'�(ylZ�)C$���+M�\Mօ���W$'��>��(��W�H��dN��4�$�"Τz�4iS�l>M�q��Үm+�D��HS7V�ÑD�4�"�����&~�"Y{w
�RX`؁e�^
NR���V#t�
8�%&�OZ�R3�Ƹ4�p��ߙ!�(���ɕ�5�j�C����F_�"�$���)�.6�f�k� \l��!ڴq_0�<e��S���S�HQ R M�V����$�5R�
��&C�u���?�2"#@�-QP��b�=����S�0�}�2%�O�y��(��O���o�����P>>L.a�R�	��I��͏Wn�R���CI$cjd#�B@�}-���kN9�[9�K��Ypn�����͌����Ð�:�0��b��9��DX [8
��N���)�S+{q� Q��B� �	'2h�� ԏ~�<k�
O��E醵�:2��Q�e�:�j��xr�#�&q��[�l\��3�i�e�GG�1n�l2�j@�p�,5�� D����- d�Y�S�9?L�s�C%D����aL 4p�H�n^?���֡"�萦̈JR�DH�[��	��6���P���Q�OD�5Ӑ-p)�?� �G��;��D�~27����`��a@/�2��2�C?i��[]�0(�%ʲi����6l�tt�'Ȩ�B���r�S���x��ɇrIi��_:C��$õjT�yb��?���6�C"�d9����� �Xa�c6����2?Z��#�0��e��-��B�S�75jP��X�+��a�t�b���L�e�'����@ �v�}�C�	����#�W֑S�).�Ӹ|֊@�ÉT�c�~%8PGJ�P�|�	]؟��
?P�J� ɳt��T�t$#?!�������vT�W��=Z�x��#C�R�ևz�<��K�	Uj�)&a3
���V�q�<����d�q��JP�+�Pl�<Y�(��l`T���'$YB`t8B�s�<q�Ffo&��0,��<0&]��Ȅo�<y�m�TF��$k�V����Yf�<�2��?S�Y;¡ǙGOʄ�'�]�<9��	�ֹ*WK��w�(M� KQT�<�a�ؾ�,Mg$QS���Q�<Q�i�y�n�P�,�)4x�
�e�U�<�p�6��'vV�j�O�<yr�ܭk�Ɲ�',I(^2��h]�<�r/�2zk=�"����t��Q�<9'lS�J����C�S��	Yq@N�<�E�-DŶuJun�YA��x�FA�<� �S.V�JՍ� �A豇�P�<�&`Ϻv&1�lڟM���p�_O�<�B��Px���k�R����6.�H�<�e�\�eq2P�g�
?r����KI�<ib��(Q�J��P�0)�D�s��B�<ѣ��6S�hL��,����e���_w�<� �y�$	f&���������w�<I&�K��yuΊQXHᄫ�v�<���؁,%2���Ȋ&`���s�[_�<��Y*=���k��ԣ'�>a��Z�<��~�~h
�᚜|<QqqdS�<���\��� ���m������N�<	���@3:�+��zKX�	�I�<����1L� p�ԑWb���$FTI�<с���]�(��-
`q��Y�M�D�<�P+�(,hPd��k8c�<<@0K�@�<�7f�tᖱ9,�-��$���Z�<��f�����iMǴ�@��FR�<���ǹG��k��(B&��bKVI�<����%X�1��H����;.RG�<�s�%[󴭫����9}2q��a�J�<� �H�N@S�]���#bi�E3"O<�:�D8�E[D�<]�t�&"OT	��!�l�:��cJ�C��J�"O��l�za�+w#�j7�j�"O(=ۣ*Q��QJGb/I8)C�"O�ӨY]2�)B���*���K�<Y�Gy��釠M�	H ��	M�<�I�
' QwK���*ia�%O�<I�h�3�:��SX�F�r���Ha�<Pd٢7V< C�Ft�GoZ_�<	�[�}���Be/��h���@s�<y��'M
�BƆ�
TTr�`DC�r�<1$�]�m�1#�M�w/l�xf�s�<I�$� ���Sfُ[̄��Cl�<	��RX�e⇆9��`إ�k�<�M�-ʜ��v%r�X��Bd�<� ���-2�}1Â�!A.�sOi�<�X1zI �)�e��${�iƅ5�!�˷[� � �jή<��U�V@b!��F���{�L�l�`�;hU�ln!��C:���Mˈ��M�0�O�V\!򄆤)�B�y$��y��|Ӳ 5!�D�.D6�-�fH�2��$C3o�9-<!�7	p�T"q�S�J�q��K9G>!���A�P��Ą�p��낭�>�!��6*�� �s���)[��/g�!�d�x�(�@e��: tI�l]�`�!�Ă+cn����b?K��<Qg�Lt�!�d��,�h��1�Ƞ���@E�:}!�L@�u*��Y��
�ho!��F�Q)(r3���Y1�+�	��Fw!�d��	
j��Gg3��J�E�n�!�	!LV��Q�nڡ1�I�ק`G!�4(U}�5���9��+�,�*b7!�D�f����b�"s���S�ѤX;!򤄋�:My�A8C֘I��&p!�6G���I��U�4��3�� w!��;��4�K��`	PO�/$S!�ԉ/ ��#m��bxq���2>�!�D��I��Y���J��Ni��΅^�!��F�V��C��	��P
@��$M�!���>""�0cIV��B� �,�!�D1���6Ùk{j ���b!�@�b_+#D�$����nɂ���HKv��aT�/��݁�B�3d���^hn�1C�¾DI �4�2q�ȓ[B���1	���dDI�&��цȓQG0l���Ɔ)j�єm���ͅ�//�d�� �n�����T5V��%�ȓ[~�
B�� vȎ�I�D��n�C�	����f���]��&��#�(B�I�t��5��9����M� ,�C�	���0��5)AfLse���7��C��2o<=�Jr�~|�VOg�B�	e���������m{ ��*�B�ɭ2@�̲�� *a�w�^+��C䉦yCX@P��J,E�s��%Y_�C�� 1hN��Q�M:��]`��K�C�	�N�^er�$I�PEz�h�O� X��C�	)78̛r��Li��$�ܢ)��C�(%��i3�aU�/8!��O-	�C�I�u`h�q��1�,��*J�R��B�ɬ1������J
D��`;bGKn>�B�IF<@��d�t�|[����2��B�)� V��1K��RtX�Z�$��Ӈ"O�]����i���K�B��zĔ��"OZ��C�2 Cn\���	6��'"OX=�m��.y�L���^�iU�iJ�"O�d+tO�#9�J�{���cl�� 2"O,| EĄ���=���ԈwT��x!*OB��A,��Bp��J��. z� �'�hī�B�j�^���N�&^����'<D�b� K"3#b�&G�p��'&P}atƀ�p"ܱr�n�Y�
�'�\���B�xp��E!�t��D3
�'m4YD���8h[5jTV�p�'�4 ����!M8��W�M����'܈�:�JS�T��L�7��:=آ���'�$9@M��v��h��LP7l��s�'���ٹ��S��.S!.b
�'P<0B�E��n�b�9�	:V�f�y
�'�Zt�2쑴|�n$�`��:״X@	�'5�1
^7����W��(���'��	4$h��Bҧ�;~zA�'�X%C��I"L�@��K�l*�`(�'���e)��@�K�ǫZ�|L�'u�����=J��3 ����8�'��9�֤ݽF���C�z�d$��'\*�AwaDƌ�!���z�����'&v�#Y��ls�)�1-L�a��'��,�R���cO��0��ϻ
\0��'s�QѢ�1]��s2m�s!4y��'�Zl�!�@�Y��!NN�7�`A�'�P���\�R���l̚0�Ό|�<Q0�ִ`jde	4�EҬ5�6A�z�<1����T�ڤC��F�n�6���^�<�V�]�VUCh\�:����v��^�<b�R�.8Y�Ѕ /p�����J`�<y�f=>���Ŋ,.�,:��]�<A�o;.�ٹ��`�&0�afY�<��XtkC��$%�<��MW�<����	��y5'�4� �E��X�<���U�t��!�r��m���P�<i���Bđ���vT�M\O�<1A��8���Y�	�1X��I�C0D����k�m�M���\��E%D��S��ĕ%�R���"5
��b�%D��Q��G��XI�MF;���[�-D�a�*X�o�p,�RA��Z8�*D�����-�8@cH#���hS�6D� e$�&�H�bj�=@�H�V�+D�����[���ҀP"N:jT"�-D���h�7.���+�ϝE�&` �`$D�� �Ȑq��	�"��	�4l��#D����8$��e+F4k��غV.#D� c�Xt��dP�łd{��C D�h� ��2�P2�ǔ$�H�D�:D��X#�V��%��$-l` Fg,D�ٕk�D���*���uUF4R� (D�ȢgG�q	e�s�HH��'D�,�E3p� � � v� �ì8D���!�y�<�z��Փ:x�i��;D����)~Q`��(<p���=D�Lq"��w<lj�lS�)��\�V=D���SD�*U��x!cM�,=d���B&8D�d�E@Ӣ>�:5�-T��dH��6D� ��=N20i!�JK�)*���DC5D�t�f*Pvک��a�!T���դ5D�� 0e�҉عD�T@�I�#*XPJ""O�,ʢd�3g���Si�b �ӄ"O�\�v/���t�a&T��$+P"OI�R�3���/F{x�8E"O�q���"EԒ1��� Qj��"O�xz0�X�2�Mv��d(��"O��H��ČNc��Y�7Yx���"O����*0~B��ڄS�n���"O �C5�Ɵ3�|���L?s���"OΥ�Y�$Q�L��B�8{����"O�����D��(JU"�M�T��"O>�1e�+i���.z�D �"O0�Z���&i�����@Y�y9�-h"Opk���<q^k�-R�3�<��"O:�A��>� E37AL�j���B"O�,d'ǫ]������Yk���b"O��!3�;a}�]ۢ�=4^X�0S"O c�NY�gK��31�����V"O����?\t����]��"O���qm^�M@�����!Wt�hr"O��x�\�X4R|x�&V�q��#"O����R-o�İ�r*�5�t��"Oِ���ct\1��*	�PD�"O$@I�NC�n��g�0�`�2�"O��y����ap��cቆ�v(�I�@"O$���[MLD�UǄ*n5�"O̐KP�Z%��y���E,r<:2"O�	�@i�y1u�_!Zu�iF��y2	X�E(�,�ѣ֠ge�|ɕ�[��y��F�X3 J΋�E� Lr�ܯ�y�h@C�8�a[�;�Rb��y��@|�&���]�?����,��y���x�!�$�E:1C�qh��^��y�ML�$��d@,����ɪ�ybŔ�3?ġI�fܜ%'�ⴌ�yb����zѹ��7`T�8$���y�C��<��K�=���4�_��y�)�}��nN�-"q��L�+�y2K�:'=��i�)S�%�6D !��y���,�,}�ת�#��!jR��y�k�e��h�:o@*���%�y��ΓKJ
��!�ģ�M��.���y��F�mUh���a�;rK" �G����y�KF?���KP��k�r�"�����yb)�;Q��sbC��]h9x`�]��y�Z�0(�J"�JF����CY��yҨ3?�,i��֟ k&X��	�y��.e�"����]�_tӃ�� �yRo�#$�=#V��,��-S��y����(��ۢ?�H�����y��G?sƶ9ss�/.�h���b���yR�D�|�rM�U����P�.�;�y��n�P��C��RM8��J��y�&U�j5�W�UKf`:s�%�y��cn�EIdL��+������y��kk~lq�E��}3����y"�H�o� =H��C�VBA谎�>�yb�N�R�0�e˄�D�b��w#,�y��,yRbA1���;#ԍ�'���yr�հQ�	�0BX$"�fՁ�G���y��ݫZzxr4�ɞ��`&�Z��y�/L�/�$��g����� ���٧�y��V;jq�12�tf��
���y��ut0��3j����%m�7�y
� `�U�M5	�t��b�5���X�"O�Ơ�+L���r �1?�0���"O�tA�G_�8���u��7V�	5"O@qSK�<Gj�	���	�W!H:A"O��G��eo���#B&=�Ⱥ�"O֨�'-�-���`B��$���"O�������l�X����˚#݊���"O&��BD��"���p�&�P����"O�% 	ң{���q�e�>d�B	��"O�%q�ȉ�FLe�E�I�B�n�"O��e�+\�\E"�iK�Ju�p�V"O�LIE�?h�̃0�T �x�v"O���@F�w����Qh��!M �
�"Oʠ;$�D]�~���'Ѐh�`���"OP��+�7ͪel���c�[v�<���	�n��EYt���}qX���*[�<yC�[
^��4��蟊;�ސ���BY�<i 2"�r<C6¸I�p�J�d�V�<����'����P�l�x@�V��X�<�����R���ϋ=�V��_Q�<)Qc>)�ZdY��8{��J2z�<A�`I3����B�;gx,�"A&�L�<֢N�'�0�s�ǻ:4��aL�K�<�Q�^���� F7�hq�w�N�<����R8�Y��8��p���J�<9F�U-E�08��E����c�<)�A��6�2(�ϒA�V��q�<!���!O2��ٕ��<uZ�q�K�Z�<q���A�r@�p�^;%ͨ�YrR~�<���Ri优P���l�xH�Q��W�<y�ŗ�n���&�x����u��R�<�S%��d�j@�1��(���QD�P�<ɠ��)F6����h�y��E�<�m T��b����}� UT�<�P,ӺT�(�R��2Z��($��U�<q�c׃/�:�� ×v���'�ZN�<���Rq��Lх�O��`�H}�<�@Iıe��9��O��n��O�{�<���^
�&�6���˪x���Cn�<9��3l�J]C�).iJL$�f�<�&�`�JY�7�N�=�*���Z�<��.R7R�e�pI�g�ru�w��V�<yE`5S��z���)���{�<R��dI>ݡ�g@�ux.�QfIr�<�Q�ߘ4��R���f�(��k�<)��_9h��8��	��=�yA�Td�<�� ';���5��Mu\%*PH�<1!@�~�ڨ�AmC1 S�Ub���D�<)qN�!m�mA� z5z��'@�A�<Q6��FB�����<e&��Z5��<9DcE�d�����9*���k�q�<Y���k.d�x$�ԝ�r��h�<�aП�j���l̘Tʜ�8"�Ti�<	7@ְx,��AS��X<��q�n@g�<�ᕂ$��c����r�B_�<Y����Mz�DJFԀ9:8aӲ��%�����-ֹVl%PC)�A }�ȓqºd��@G�x�^����U�Ɖ��E�,�8�ɀ��:ՂWO��%I�@�ȓ{I�M˹=��%�p�"TL�ȓf4<	fVw�8�#p	E���ȓ
���2l��$^�f��"��f��rg�t�^�P�i�msL5E{�LN8	l�����wNİᥚ8���M��"|tʖ�PI,P��%G�O�hi8��@�nm��B�\p����OZ���3� P5A5��x^:僰���6	j�
�/�T������?a���. �a�D�R5d�0�4`č����� j�.QKV.�ޟ�0�)	�/���'0u$�)�@K�m ��s�˒$v��
Cg�O����H�7�.M�q[i>��f�4(>\�@�'�m*��}�ڈ���+b���D�!MĐ7-<�'vw�D��.wXP������b㙩lU
6�N�Jѐ7��$!��pv
;��(^�y�B�4�\]�B/���`���UG,�M+�/��m�!�O�0|ҧ��)/��lJra� ���5�A�}�
���j�&$TU�/1Y����S8K���+v�f�t�z�'W6Z�b����>b�|Th�m�-wzpa�e6���s$�QXh������(�x �Fh��1F8��ƛ,+(,�R�G�o�����E�y�:�����">�=�Z�Oi^����C�h�*(��n�3q���	-�d�($GP86�j]H��Dr��([k�Bs�k���>�V��e�b�s�Q>��W�۾{��B�F.9�H��ć�h��5���E��O�e����>Ppxұ�5)�Ʃ�p"O �����L e3@��1NLIS�"O*�9��G(1��������- 7"ON��	S:�b���[�/��h��"OH`SIA�� !+];Q�V���"Oh���a�Fz��`3��:c:�A�"O$���9`d�0�ɡbGL H�"O\4�l�	d&$�&�ɱe#1d"O�T�Ζ7i��|��
@�C��A�"OVu��/�
R@��pB�iX�v"O�y���� o,�MS�*  �L��"Ov(�qD߯r>eըW%vup%Y"OT���D�,�:�	&I��D����"O�XT)�w/�����S�4$<��"O\案�N��}���)u��p��"O���! ުV2T�.E 9�*��R"O\8�P���W�|@�T���@"OPI#
�t�ԅ;6�`��8X�"O"�f�͏~�<���N�q�0�!"O,��fOj�NT�mM�XΤ��c"OX���Q�%�H�bZ��CIەI-!�d����{!A�W�ب�H�O+!�V�Y|�9o�VV�x�ςm�!�d��(NT<�@_#HF�d�P4�!�� JٰL��f� �Ł�@�9^]!�$�( ɬ1� �3q̖��0�2
]!�D�,dyJ� @�~�49*��O3�!�$�p�@�#�<n��Aд�=?�!��
/�X�r�oP"D4��b��$�!��Z ��"�W�=R�KEM�t�!�D��9�xU`��</�%ȑ,� b�!��8�I�FH)J'|�s̍6i�!�
FG��s�$��>t�AI�k�'x!�$B��� �%�<ep�	Ó	��+!������+��;��A���D4�!�$L�h���Cc �(���"G��g�!�øE����֘"0����J�p�!�Bs������o.�{���t�!�ď#2��8c���<V��豧�.�!�φhr
�+@���������dH!��ņ(E��4�'6�@R�-D�@�!�&�2�p#���}��u15��L�!�S�T�d�ݘ �p�t8!�Dܐ`eZ�j� �?[��"AE D+!��N����B���ʜ���!�4Wݘ�'��F�e����J!�d=&q������*4�8��C O,�Py�a�61�h��$`��NH�	��ؤ�y�I��J� �JBF%D]��*b;�y��Y�i�lA�̅�$tK�*� �y2ς1LD:�!��	�����Qǘ�y�)�Q�@X��Z4���P�S�y
� �u����'�v1B �xp�"Or��A�9CG��#�,�/b8��
�"O��{!Z�*�����SKRD��"O�J�޴YBuq��GS���:�"OJY:��a��U���^�|$]��"O��2`�M�s�l��%�0 w:h*�"O�!�`A R�9I%�Ϫ @"O��	G��2x<�I1��f�yʤ"O>5k�f	�4z� CL�9���Q"On$���V�(I�-BՋ�)n�E��"O�4�Ǥ)�0�Dʊ�"m��[$"O��;�c�AڀʄH/�B�"O^�RY�<^
e*�I�r����B"O�@Уٲ��掙K�4H8@"OyR)���~]���)WMТO���C�Q����"Q	H&�c!�d��1����ț�_�0���
 (�!�+a�2��.E�%�9�'�X�>�!򤔥EJdi1U�9b�.��% �!�Ğ�b�t�K��.J�x<�'��!�!�$K4s�}���ǲ0��UC�+
�?�!�I�o<��`���{:�pKg+	�t�!�DV5 M�ȠЅ�U6,4��!�
�T�0�0��+�X�b]�!��0����'b߱&c�ؓ&B�G�!��G���T�H�5\���"�'�!��FXZ|qT�ٚ}7�@�U�?�!�\%f���c��?4^��4�V�y!�A�uu0�:�*K�{3�<y���}!���X|S�`[#o�E�3�PS!��ؚ{&�9hv��/m|H(���ת?!��ݷ��L:�C
 8��+!/A!�D�"V��Ti�q����UÄ�5!�(z$�u�q���=�&xAB��j!�DF{�X`��P�Q͊����	�"OX�	��;nrtr�ꃶk���"Ot���m�1�� �^����a"O8 ˴-��v.�Izbk_|���D"O`Q�j½3��X)�Ƀ�^�b=,�!���9TꙠ@eTG�Ri��	J�!��n����,N�R�8��(��Y�!��(h�i�dn��F�Mᇡ�#L�!�$ŭm�PX�wڙ-�u��&	�f!��+R*�P���a���r��:�!�d7$Ru$lE�Y�0�
�E��!��4*h���1�	:'F��ZufN�"R!��P #��Y�O��,�����-c8!�d�6���b!֔�+��'!���&3��R j�]d�ia!���?��s�Z_��h�O�J�!��3L	T�� LF�O�r�-ܴ<r!�D �e��p�-�M��̳fI�!�Ds��̹s��9Si��g!��ɾ<�fA�%�юz|A�2��!�!�d�X���Y.P�}h��� d��&<!�$!?Yڐ�_9�ȠA�Z/W!�ܘrb�e���sJ(r� 7:H!��E4�Y�R�].h��B�#ٞ^!�d�����3���[�<u�Q��,�!�ć.<ۺ�97�
R&p2Q��;!I!������(�<K�@�C��k*!�DٷG(��+�
�d�p��F!��324d=W.�(�(�CE!�M�Xm2�٧�Q�1��p����g!!�� z���+�c�\�ȶ�I1�Nqô"O��� &*�2����2�H!��"O����k�0 LD���A~�#�"O.�p�LÖDj]B�2v{`���"O�Z�,��NE2ŏZ<%]̄Z�"O�D�� ���53s	+�v���"O�YU��;4�1j����Z1�D"O� �	�܍i%f�~Ū1��"O9(���N�l�=K��9�"O�ذ#�]�1 ��:(-�9��"Oz� ���=)�ృi_
**�qY�"O�x�B����H�_�^�c�"O��z�$�)�L�3f[���"O�0�)M�)t�1�p�~� �"O4�R��?`�B%@��D����"O̱���:�e�v��6> H�"O��A��~���ǭ�;Z �y٧"O̽�똹z���w.�9�"�چ"O��Ѯ��,�,��S��.t)�|Q"O�\�f �k��J�L���A"O:�kc�U87��<{I� ��I�"O\�*��ڂ]�pX�aH͝}��ZB"O���F�e�k3b^X��t�"O��/�	J,
z#L�2�d��"O��!��;�ʠ��<#.Hha�"O��;c�Bv�]��Ad�F�B&"O�t���R#�Hv�9"�8Q��"Ov=zG�Ľw(������)0�"Od�)+SP��kF'
D���"OPe ġ ����/�+�1�'"O�`�l��hopL��� kE"5��"Oh�A���|e:u1�ǌ,Ӛ\I#"O�QC��'P���(RFȠ��4"O\H
�A\0Lix`�EƏ�4u�p"O��h���rj֜)���E��"O�EȂƬ$"����>3�¸�"O������B�� �� w��j3"O�iD�c*��熩Y��]�"O,�Qw�ԉI�T�Z%IW�,âq��"O�yP��.E�<h�p�K=8��(˕"O<Qz��H����I"�H-��ȓ"O��ɕ�b����k�;D	h"O^�c��d�T퀲��u�$�"Ov����J�L��ᏐV0~�� "O�i3uO���!sG`��dt���"OH�zƫN�b�r!p�E�#E�n%0&"O�a
S"�2������<}��u"O�a��'G!Lvh"qOOV�	"ORX�a�Vz�ޔ��ɧ_64l�"O�y��P:!���aP	Og�-["O�E/c��h:��8Mr5��"O �≪u�D)��(����"O�4�i�|��A�̚@���y�"O�!����;��I��Q���e�"O ���NJ.�hAJ������8F"O0���[�4Ar�6=�y�D"O��$�� +"Zѐ��|֔��"O�P��Pmn�#��V'&��B"O�ͣ�g8����N�8XI"O�Xx4eW'\$�����'h��"O8�J�E�e#��SCl��d�t�P�"O�]8��+yFI+��U�Z�PM�F"O<yI%�S�6\���Cv����f"OƹAV�
�US� �!�>���"O� J��-9)�.(�%�O�z�2�z�"O*isB��/���[šУ^�.e�4"O�t0�Y�s��9��ƛ�h���"Oz!���3Y�Э��[(p�"Oqe�R,a�X|C`�@<M���9Q"O&0AA�G
F�]8��L��p�+�"O<D[q��%OX�A�P��0�:�"O�U�B�Z�.#�	U(E�1$��	�'��M�	L���qDN��d*�z
�'�x�8��A�7������> ��a��'��\R ��.�fQ�F܊�&xp	�'�0�c*>6p�Zt�ש	K�!	�'Ҽ���A5����dE�P�`�'ܴ �e�7b��qsբBJ��$�'��Ł_�Bq��Ҵ)N�q����'���2b�B�0�v�Hd��%l_�8�
�'�ށ3�Λr�}�3@��i�R���'o�`0�O��c�̠BA��d��@�'C0jN�;q�yȐN�]k�8
�'}@���kM�~��$������	�'n �у�+�Mb��D����	�'��0���T }�$����ԐK�'�>��B�L,F����O[�dK�5��'%�Z玍� t����^ox��'����,�/|���dM]ؠ���'�~�W���=�P�0B=QQ���'�T�4G�D>&h�U'�h` r�Op�D�?m�� �4�?��'���b�t6���:p�D!���"�s#��?f
l�	̟l� �8#�@�@�i8(lD1v ���u�Ŕ��i]k\�"%����BBZ(sq�'}��*U��,f�(d��k7RX��Z�p2��"��n����b"J�6'�^(�K�x"LN��?	��i��7��O�b?![����XZB�cR&Db��Ġ����'��Z��g�8O2(��O����E�Ep��d`��n�n�ɉt�^l�'ɦs�n����t�5�f�i��'���U���d�'o�'���d-Z��TD�mH"c���`�+\?-v@I�2���ł+��)�O�t�� |l���/(d����S��5���@
�+� L�*��\A換�X����3�ٹ��O��9Q
q�qC�'����� �g`Ju@�J7`y�V��<)c����O�L<�CE�!���0�>C��c"�G Q8��'�����"|�'�Љ��BQ�O_h�wa�	gst�N�,�ߴ!1�f�|�O���Y�p�V�_6.h��*�V	~��33�|�t���?��?���&�n�O�$�OK��
�bw�Ԓ:k��@���T�걏�v@H�1�F�6���n�3b\��7��9Hbz0I��"J�YK�!��8�	F'��"�8�#�-5g�裭��W:�x��I'���3��2��A��P!8+`����O�������My��'�O���"�:&BI(�ꄼ/w�d��>�����	�Ş
44%���V�1��X`�|�oԚ1��6͡<�u�U�{���O�7� �52���-i8�-PTi��P���	� �D����I����v�M�LA��aW�i�Ќ��E21����7+;6+DL	���d�Z�jP.ږN܎�<i��E���eHP�<[S�U!>b4���	"3+b&�Vn���C0�3!B6�Hqܓ! B,�I�MKq�i�fŊ<��W� e�:y��ǝ��LY#)O��D�<9(O�c?!JB� !=�H����8��2$�\+ � ?�X��ImhBY�Ԃ��K�X�o�˟`�۴!��!P%X���쟬���u��nZ�z��}	S��-KHxs��҄A�����?Y��H+]m��ũ��Ơ��F�-JH(�L�>��S����2���.M�*�x��.;�O����׿j\6(%��!k�Y��//����.�^�G�٢6�p�@��F�/� �x����?!�i��7��Ovb?�8D�3{�Q��^�O�t٢��3��蟠��uT��dN�g�q���qrR�O0�=9��i?47�>�$�A~�q�+����)�0b��Xܴ�?I��?���H*k��C��?Q��?Yc��xH'���go�A��D̙h@�=8��dQ�P��M ��B�=��ʧ��[*�IhK� �����KDX,����BD�Y��8 r^'sm��2��Ⱥ��~j�	�n�;3 H��@Ǭ ��=	���(�L�	���
v�Zw���?����uצنp�J)�5hP�E��EBqO_�=m��OΣ=%?��2`��k*�:q�f9T802f#}�q�DtlZџ|�ش�?���������/D�y��蛓Xm�q:5�U\��5�O�Pjg�  ��   �  t  �  �  �&  �0  7  C=  �C  �I  P  WV  �\  �b  !i  eo  �u  �{  ,�  o�  ��  ��  8�  ��  �  E�  y�  L�  ��  ��  �  k�  ��  �  \�  �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6�F{��'O��V���&�;�+0:��x	�'%��"J�[�]�R�K2r��"
�'Oe#W烹�R}aC��z��
�'��;��7�������L	�'�:<*b&K"4����M����9	�'نx!c̓>�D �,ݻ2zX�R�'��@ �F�9<�m�7I�"+�a�'ր����>��Y�
�%&���'��0��3L�r5��M/� HJ�'U����J08fx����I$p:<����:�'�	�T���k����	�R� -�ȓ2�̻2e�� l���hޅ2�@t�ȓr�N {��V�%.�k�N�2�v!�ȓJ��kdF~Ѫ9�fA�0ul�'��"=E��	��ʙjs�=����-�6��?��'�X��55k ��`$@�0|(4�yR�'��UAԊ�Sƈ�{q���,��3���M�Oʨa�� �&�ʌ��^�|V�Y�')d�ʶ`N�@@峥/M�e"��	�'����D+Y3,�ɤFݛP0z��	�'=�X��HR8��
�H�_��0��'�v���/6.�����$���9�'��V����� �\>������IX��٣�LyV谁s��,`P�!�"��?��y�V�?]
�j�p��Ce@
� �P. D��#@�P�R��B	�i�\%��h?D�� X1pB"��j��)È�X��a��"O-ۧ�E929>TӣD���mx�"O��[���eB�YK�����"O�DЄ�Q�/�D)(�*�H�R8x�"O��vf�1��ʒ��9v���W"ON����8���C���0hVR�57O���$T�$Re:�h��N�����?8_!��9�Ap�j�b� A'i¬�!���";����Kd3���uh��]~�O��Jsn�{�d�1�� j�@��'y�'L)�F�Ȉj0z�:V���*`N�	��D O�533 GC�d<��+�A,�G"O84�ɏ4tSҘ��J�����v��_T؟��ī�Lf��1 ƈx�A!�o8|Odc�PDl�?p{ 92��w��Cl7D�RE�C���h��V�}<���2D����ΔQ�� U��i �\q��<�O��2��13.��2�^�*���Bd�ȓ�L�Ahԯ���#Ҳz�` �ȓJ���2�68ra�TeB�WԀ̆ȓX:��bc�?�r���߲��t��	h�	�V�@�����
�e{�־~��B�!-�5Y!_�rY\�W-ɦUh�B�əX���"�>z��� B�	��>��чM�-'H\1m��r6��=�%�)���L :��K�J	"N��ƓD��Hd� M�t�'�D�t�N��	�'� 5���O&3Z����y\��j�'�ў��8M�|8qk�Ah2��@E;Bؑ�ȓ7Mx@�ϧla�%@Ч������'��~b��v�i[*��x]2������y�DYi	F�ɀ)�wa�݀�#���'� t��I/{�XA�Q2@��u��)n��<��ҕ�×�����"E�_"�ظ�aB8�y���9��#o��n�Ʊ��J]��=ɍ{�n�	*<��b$Ͷq�:y��K9�y2��4wr�"��e���c-���y�P�!sdQX'��Wu�i�����y�h&L�d��	^澩 ��Y��yR�'���E��:t3@]�C���� 
�'Kl�*A�#�R��d�� 	0�S	�'kĨ뢏�%,!"��/ ܄9�'�H�0O�)f=��馃R�{aB���'b�K��%; mCEl	�j(����'�2�a��/<��ubw�\�e}�q��'�§Ɂ�/ZXa���ePd�Q�'�|��(ʘG��E�e��bQ�M�	�'nL8i�CL ����`��0)�'��C1-c�Aր��V����
�'��\�0`�M�ld����=�jB�	:�*�h���E_:�;&@�+d��C��7=�p3��T�;��-g��C�	?j%����
�p���ޮ/��C䉒Sq�\��e>}Ze�W�[�ٰB�ɶ`_

�%���@���͌t�C�� f��k�\�`}ɳ�̜Y0�C�I8��mZ�.9t~���I%~7dB�ə)	�0���ΫoȦ�(D@įYL�B�7F����j��R�P�;"��$QzB䉽Z����e�
R�*��cJ�7lpB�ɧ& R�@gɛ*0�B${���%WC�=>| aӪ�*Z��Y�q	��b��B�ɪ,�	�h�gW��u�Ŗ��C���4Itb��(�]9W��0B�)� L��a�ʟ)��%`CMӰ
"r�%"O����˅�e7n�(ci�(�DI�F"OR�XšB$-UZI@0	ڍS�Bqv"O̬@��<5��	@��8P�s"Or� 0H(;��5�#U��p��"O �Ҧ��gZ�t	Q�
X,��"OL(��jr6(���GR'"1D���mT�D�����;d�6 �BK-D��j�E�;��qɷB��5����.D�b��F�	D�8�Z
	�B�	�1��M�ES� �*���B�	5(�Z��߀r��)	$��k�|C�	9=��sQŀ�|�)��_RC䉂}�Mw�ʄEF��+���"C�I%Q
�
�U�&J��¤U*w�DC�I��xaCFb��p���n{"C�	�j��ђ��	p�H�Gя ��B䉍n.�C���~�����M�b(pC�vK��e�D�;�� f@�PRC�	'LIt	HSB�7Ƽ�奊!#�C�	
&��#T��<Rz̐���g�0B�ɝ.�<;���NdCṠ�j�(B�ɝ"4�qW�٣E��xw��_�B�	j0��K;$��"�B�{gB�I�`��U�`����K-ZC��a#d�i@�R8�����@@�g�TC�Iz���s7�ٙ���[u�-t�C�I�j��d�V픭E��F#Z��B䉸~jTq�O5L&d{D�Û%�B�&U�ld�e�"T��*�N��B�ɽz1�� � Ӏ����i�$0��B��3`���Dӌ(U�Pa���[�B�I�G���Gj��|!рѭI�B��&#�@��%F��=<����Y�+��B��
:ژ�A�j�&����l<�B�I8[^f(��Z���|*�J�v�&C�����
��\����(E�B��l!q�h�N���B��pB�	<fb��q�	|y6�8GC  [~C�ɍ@6r�� �4�\�.�16kZC䉡��,�q)ɵn�r���R0LC�I�����l��a��ү�-iC�	6v�X�;��ݲ>v�p�FZ�'��B�	�7��X!�96M�yɄ�K�%5�C�8�� ��]�':hK�GfB�Ɉ2v���8<eL�����C�	�!x�'�+@�P8��E�9`&B�	�~� 9�*C�t<q�6T�B�I�|,�y1a�\YdLF�Pf�B�I1ui��Z&&�0��Jr@��4~jB�I4J*�)?a����f�<Z��B䉚\~8�"�V�"��q��n��cvB�	?Y�ZEp'EV4��`�O�$+�C��	� �	��8g���P(�=`�C�IDo>=1PB]!d�E�`��%$�C�I3M�B�u��^p�h�"I�C�C�ɇ����CD�~*b���CG�|��B�	�T�ȱC/
��ZeXӎW�s��B�&$pr4H�� ��`:�cR~_�B�ɏR{RU�e�Ya�$�����>�B�	,��8 �;zi��32��v�B�ɽv�H���4�֑���μU)�B�ItB]V��z����O�'^�B��� S"�$QV��� R{V~��S�? D|P���3h���@��Of��d"O 1��/|l ��a*׹QJ�+@"O:�bT	Q��Llq!��=��)R�"Oа��� h�����%O����g"OhT@䚑
nL�x���
�$�1�'B��'��'G��'K��'���'Fz�쁖t��4*!kA�S���;��'�b�'�"�'���'���'���'�2L 7��L �HR��q�$L ��'���'���'"��':�'��'�x�!tI�3jԤ���W$RY(0�'���'��'d��'���'.��'������Y:	!��˶^�h<��'p"�'�b�'R�'y��'���'~"(ɂ�#���ۓ��3��"�'W��'""�'�"�'���'���'Y�eЪ#�\l�D��=BU@��p�'iR�'?�'0��'�"�'_��'g�52�E˽;���2&�K�D;�=3a�'G"�'I��'A"�'�B�'1��'I��Kƈىe��� A'D�(����'sb�'���'�b�'}"�'��'}-r��I�]Zv1�g�74@��'�r�'k�'y�'Lb�'>B�'۞M�eFՈh�%�D�J*,R�J��'Y�'��'x��';"�'&R�'W�A!�ř�s��gR%.<r�@�'E�'d��'��'��'6��'K)Sr����hC���6�xB�'h��'��'���'*��dӾ���OT��c�>�	8��!�ҹ
��E|y2�'��)�3?��i9�ѩ�n �v��E�5
�>�4Y[�`߂��Ćצ��IB�i>�Iҟ\a2��bJ��x�BVo��aH���şh�I&14�ioZr~b1���k��V�8
.̡�0A�)��(��=�1O ��<���)cq�0ԏU4^6�X��
8_��m����c���f��y�@�7/������9ό�(����pK��'��>�|r�Κ��M��'�"�ʒ�\�@��a!m\4=q0�'e�D[�@��i>}����IPZ*f�8�"C�>����dy�|Kd�21����.]mvM#E�p�`��n�4|k����O����O��}}B/��0�u �`�hA��I�����O�Ƨ�� 1�� � ���΁P3"�2�<�Ƚ���:��ʓ����O?�	��4������	q"+K3�牄�M�t��u~�dg�&��S�U���;��/*��%xro�&(3��I���	ǟ̐n�����'�i��?���)���:���]GF��+�h�M�� ��~�B�e���}&��D�-.��a�u,��T�a��*D� AfB1c�d�8����f�z�y�F1k> C�MԍH�<˖-D�	�Ht��g9r�,�gɼr�*49AA-SN ���?2L<eqWG_;�����`�,��C^A������/0�AA��)���BZ1 �F`Y#��X�� ,i�@� N�;��m����C+I	#
�p��Ն<R�7��Oj�d�O��I�{~�	`��B��MOL���CX����O��3H?�I�?����V���iT���e��/�p��%��M�@�_��&�'0��':�d�7�4��Lcf�Fζ�b!Y<��lz2GWަ�i"A�v����<y��R"R� �Lx�	�xI�ʷ�i��'���ϳD�O��O"��������u!�=�nZ���j~�l�����Iɟ(루���I�O\�d�O���ݬx��1��c�>qr�  1���2R�oZ�����Ϭ�ē�?������{��,EǪ�c�
\�+L��aI�����.���	��h�I۟P��s���'t
a�,�B(��ID�i:P�زeO.6�Or�D�OL�� �d�O�HBj�:{4je���<Kg:)�,�Q�1O��$�OJ���<��	1D���5
�z�ɗ�=ф�	�f�'��|��'���^!���G
���7�1>��������韤��ןt�'��4"N&�,|g��x�m[++=��8����j�n���,�I[���2n-�s��@L%Md���ȹM�rm�ºi�B�'C�ɮp�FN|������ɏ$U��S0K��h(��jQ-:}�'"�'>b��#�'��'��'`��Q�E��$CP��`�D��G��hm������-�܉�4%Z��۟���#���(@� "�gVD�l�0��(T�I�聃FE���&��Hd�I�2u�L#��>%�Ⱒעb�PDp��֦)�	����	�?Y�J<ͧzN��K�E�Ō��6��+f\��K��i��T���'���'(��O%�Ss���%���QA�֑:��\���_l6��O˓MM���(O��v�$V�?� �1��Ð�(�q�'�	ǪA��OV�D���`�.��I�P1)��8*Cb��V�a����1JRʓ?�S~��u	��qv�C�i�h� `��P-��"�i�Z�k�|��'��'��	L�fTѤ◴o4��Ê���G����?���?�.O��D�O�����B��\�⅔*���z�&��F�r�D�<Y��?�����9b��̧s<�,��M͛>��i���n����'n��'��]�����0�e����YvH� n8�b���,~(�B6aӰ���O>���O��3�� ���d��24��!��J)
<�x�g�?bm^6M�OR���<a���?�6� �?�*�2�;Wmi��5�J�5ٌݫ�aǦu��ɟP�'M� Sl'�I�O������g�mې$!'W�+�("4�i��IɟX��"]$,e��}��?�8� � haꄡt]h��!�<Ȃ��xB�L<KA���$/b �j��EO�İ�4ƞ? !�U�\J�iQO�n��p�`��3Z
L�Ed�W�TK�0 �h]�ZaBs�	�1_�իǄO�1��)#>~<�3ƊC�u��菬)�P��$@%Y��D�A�$z�Ƹz��
A���D�H�;-ܼBVꊦ=� p�C
+E8��� �a���֨Y��vE�~]�����*������O���O��dL�����?!�O�~Ƕ�҃�c��4��	
z���N״(d1I5�K&(^L �'~���TC��;U��Iir��'b1�s�B�6 9*kӍ6�b��%]� �Sz�'2�R�ە5Ǆ�Q�G'gJК�'ߪ�����?a��x�'�X�Lk6j ?)l��5��6B��t�0?��9@�����.F%���p���M��k4�i}$6m1�4���I�<�@d)7A���JzZL�L�LTʔr��ƈ��'�B�'��h!��'C�=�L�'��%b��e�
L:�\!� �<�p>�`�6?y�k��|�D�A��K�:9<m
qZU8���I�O@��Y���%�фch��Qgi^�DD��O��d�O1����^�ф��	lf,B���T���R"OX��Ģ�:V�܁Qd��K!�e 2O��'+ўb>%�Q�2�qA� *+c4ĉ�- D�$�f`	�9����1F��Xp&(K0a1D���� iVn9���7��A�<D�Pz#�]:1��ȡ��7tŃ�l7D�t8��ӈ$U�A���z�Z͓�*D�T薁�����dOH(|��%D�#���"�pe���욤 �.D���b�{"tlٶ놇U�\zt�'D�,P��_��0y��@�$(�C0D��+����p����ُ]�P��+D����)�9|+�q�0DT6$�d��SJ5D���r�ɵ+�vL�"iR(8%NLS��2D�8&��w�dQ!g%�@	>xB�.D�����3P���"`�=|P,�q�-D��ꧧI�o���co@�=�B��Ү,D��S"ϵq����o�,��r��%D���o1T�2A.@;B�4��(D���g	�
9"Q��]#b������&D����Ȁ�k��K�dƆz��Q��a#D���p/̭ox�2�%À<�L@��"D�<�����SV��Rj߀cH��a�=D���M5�`�(1c�#>Y�)k(D�|sT���Р�L�$�E�$'D�3%KE�]�F�+�L� f�[O1D�|[�k��VF
X��F5?�����<D���DѮ6x"�kS@�:���s#;D�p���S�"�����2���"%D�иrl�
?���B0l�l�F���&D� ��FQ�R��m)�Ĕ�IG�&'!D��b.�_�
�,Q3)�@D��=D��Ȑ$�#���:���U��5�n>D�qm�15[��P�����b��/D��`$�DI��(��!�D��0�j8D�4�Wa��;-4��$�¤i�����F7D��ZvF����H�_I��A�aB D�p�A�	d��8���,*�]24m8}"<�a{2ϑ+4�`�Q��ƅ>u�*�� ��0?�T�B�9\��w@#];��Qpb��=1Q&h�<Ar�R�CP<H�䬇,}I�E�eWf�'��Uiq�g�OJ�P��A�i{zI���8h�q��'�h�GgC�PtT�\�M�LJ�'�6��I�A�S�O���2hň5`��*#/�Ec 
�'mtX�A+J-lZ�-Y� 
an�4'o}rgْD	�	pwO�yAx���HO�A� MPH)�`�^�>AKB�'��1�FB��@�x���J2"�!JD�ͧg(D�x2)�sP�� �ʑ�9��}x�JD�g2X��	�`N8�1ɋZ5�i����MW��c4jM�0��-��C���&x'���5D*D��JR,	v����'O�B�	Cȡ c��JD4(��z4"�ȡe��*�qO�St���x0 f�� �@�u�,&��A�D�J�ܲDO�A�q��"nT�7��6�6�����	 W�ll!��/D�8[�jЭjQ� ���;�T����(^�f,6�4O0��D��D�H2c��)d��lZ@�T��f��#{���d�˷VA�D�GU�/f8=��@w\Ũ�mM�r ��S�Ί6��T�'e@���$��U�:t�䖛x0��=ͧ[}��K�a )
Z�PF�ԃ$�
h�ȓ`VbE�QL@� ��1v+E�wl��	b-F�x�E	��6�)2r#U�7���;W������I��,���rh����xg�΋
�¨�%�%��$���H~�C*��xK�ևQo��{U�Lx�'�8@�ER�e�l�����&��ÓlJ--apy���ɌF'v\��� f
9�����zz�(�g��Gä8f���H�i�C�'���cRE��O����b�?q�@(�O΄!���<?�⥃Td���*�S�{�O2�\"EN�r��l0E�@�CLz)�
�'�eB��X0T�a�|���ɦ	Lt��"�[U�S��i�<��˚w刄�u��6V&
P`�!H%+0,�#
�'e���a�W�PH����Iٵ���@��
���F�.
.�3c�h���`�G����Fy���7:4��K1g�4/��W��7�0<�%NO���Z5���@�[�M���ied�7V
i�E&Q��Ic���I^E �0�ގy���#e."�z�:��D�旟�)��w�d&2bAz��Yw$������2Q�}p�E˺���':ܒ�̄%�VljF'M4�M<�Є<��!hD�Q�R���L>�OB���a��h0� yT� ?�D@��H�m#!	T��[���wF��f���@��Յ��%�JazK>E��4[0��QLĮ>y�v�J9�4 F~��L�"�v|�bW�M�(��:XG���&%�\}��P�0���8��'�$|P򏃔"w8���ю4>4���O���iL<���WI���ᜧ��+�/M?�DI*r)JM�� ��B��p��KKu#B�I[ϒ15iT�;v	;D�N5t�7�I�c&&�ht�O�UA'�M#�~�'O;����|���d�rU ��V4y����>��H�Ҭ 98�����T�cc*�(
U9wM2���WiT�(�6��u��JaqO̠�S���E��h���$n&0�T�I�"�-qOS,T- q1�	�B��7m�Qb�1kG'߈:�6�Q����͘1w����gT����I�pt6i�S&׏x�&�k��p�r9~�!0�M�7�T�3��Uz4����~��O6z]i���3q�Ժ���5B�I.i���g�ښH��ѓc�[i4H���L�?Ʈ���']�����	�:�t	&��$�Ĥ&m"u�� å.)��`�|؟L�@��	��٧�U�Z:�8$�K݀��'.���p�,tK���q�뒶N�qO\�zKC`i���S"K^n�R�ɫ�IGM�R�2�tc��J.b6-�9"Z��Q�n�Z�쥀!O�^��!�e�=%l6���N*�p=١--YL~=�N@Y�)�"n�}y��A�d�٢�i���Ғ��f?��bMl�֝"z���t�ܕ>! h����'J�C�:����H��4��ɲt�%�6�Nx��R��ڟ�C�l]05�*�dX������(Qf�1�J'�\A�%H�>���h�f��C�N�1�	�4F��	��Dn��)"�#D��(�A'ș�`��O5XDJ݇R�9G�2)ʈ�6�'j>m����9x*�HSB��Y- ����E-�=�%L۰E�����цb���[�*ʃB�Y��'�4��@1�l��.��D��Oj��M�� P��� ��&��O��[�ߏW� Ar"'�vN=(�'<��FA�)$*�2�a�L
v�c��Q�,����D������I�.}���8�h%𷉜Iܾ���+G����x�Oh$��������@~5p�"=��E �h��U:���Ct�����?���(v��5��=eb
!ac��B��_�6�$��9������s�)#��Ĩcv����FվVP�		?�F���'�ڥ�"�n;DY���L3\}�1�I����My}"�M: �P�O8��af;��M��H��I!/0p�4��b"Oڱ���Ò�,$B#萒p� "�2O<-���R�����2���4h� j����"O���'��傷���V�UIe�>�g�+��=I3�^3�f�F�i� �B�́G�<�%��/= �3AD͟���a�(}�<�h�7�tR5eUc`�tz�<y�ѕ.}6|��^�J9F��Q��{�<Qa�H�"5���)�\�ǭ�c�<QWН|"�5(�j�*`
����IZ�<� JX��SL�v	�K�a%��#5"O��"�x즔�E��H��q��"O�=�wf`vE�C��,���"O��@Μ1�XX��,@�L�Q"Ot��։��<��A��D�j|,,z�"O������n�
!�_tQ�G"O4�c��ֱf�)�҃� c�+2"OҔQ�τ�$&����"]�l�"OT��/p�{�M���@(˥"O��L�0z�ڥLC���`�"O�B��f�2��g�`	��"O�K�
Ю$T<�ه:\k�d3"O`=S��h3�S�ʭDy���"O|i���IdD�/�D��+Ĩm�!�D����@�D5Z�x���kԖ�!��@ m��Q���:�(�6Im{!��n��Гw�ߡ�^5�ƈ4$c!�$Od���‛��F��8H!��6=�)C�H��iV���B��+�!�$B�-�ԍ���Տ;�j�;Jےya!�$�b澰� e�(sQ�	�EC!�CG,ʓ+?"�B;&C|*!�$h������өV�(� 6�
�]n!�����qd�&��ؘ�E�4[!�
�l�\Dkf� t���r)�A�!�D���P� AJ�Z�$\k��Q�x�!�A�e���-��p�@�� $/P!���&`���
Ę8*gt�h�e� 2!�*Y:��'� M���{��݄T!�$C�^�9Z�n�9��pږ�)m!�пy�d�Ѡh�l��N$W�!��<Y#,��'�$�B��6�־nX!��fV��Ö�V3W��K1Y�!�DB�Phx� �0U��x�%&<�!�D�7{�K'�ǁ[y�����4/�!������λ]���Y3��d!�Ãy�F���e�7\�8<�v��>b!�DV!,��}sG��"�i���P��!�D�*,�CK�q���%� "u�!����)�B'�?�l�7��/!���y��P��פK�ځ�%,�
7!�_]�ڵC��%�j ��=n#!�$���9��>�<(�B�!��,5�ƌ8�ձo�*��N�1!�䐆r�>�����+2 �і�

&!�$R�9�|�Q��P�eIH�w"��?!�*>Xy���4N�����%;!�D�+8\y�&T8[�����NrC!�$C�y� �1Vf����T(A�W.!�$�)� X����C�ԋ&2!��.���
�L]�~488��Z�!�d��)�<Pp���Hq��{�(_<B!��B1� ��]FQ��Z�T�!�"�x@q���xTE�TMN�!�d٥$]Z�GoܞY:FP3s����!��Ka��@k%	΄�x7k�gj!� K��`�OM=�앑�*��Oh!�ݲF	��S�� 4�>p��V'V!�DH�SR(yb�L�!,�i�u��Mn!�O�,b�J�oG�$"�	�"�+Uj!�ĭ:�8���L�3n�
��h!�$�Xn�D��j����BHFl!�$�{q�дj��~IrAj���8Qe!򄟴o����UG՘#�X ��U�a^!�� �L���܈,�X��1��*<�4��"O̸����
n�8"a��J��!�	�' ��y�,�O�b�	�nR�){	�'F.P˧NS�u�e��ޚ\����'�x�s4N���H�n��X��0�'��ݰ��̭'��§M�>$��8�'J٘���Ndؼ��	�"$�bT��'蠜��ç*f4� �L��Q��'�H�2���!|�L�b�D�:X���'$�A�Վ���A�F<���'��
3*K$��u;��A�*'�`�'�й��/E�{�H��uN�=*���K�'-��q�bK�~v�Yudũw�U�
�'�T�� �]U�UC��=dh`
�'�ʔC0� t�Na�5�%5��Q�'p*�@P�Q
[�R�pfi�,&�y
�'���r#��/<>FO��#���S�'�P1�h��e~���IT�����'A�Y�g�Xw�d�4��If��i	�'�2(�����d�s��V=A��t��'��I�a���|9�ii�m'd��R�'!���f��&�,aaAK/"*.�8�'�6�HZ�.P*���n[�P�+�'�^y�kD�Nt!	�+}�:��'���di�% ��i"I�p6��r�'o�(�ѕL2�	����o�q��'��B��\/{�ΔR!�h�����'���`��^%��!�i�aC
�'6Z�AѡJ�^hċ���kb�H�	�'&aTm	�y���%݆hYD�Z�'f %���,��#f��].�(�'��E Հ� 4U���N�)�,��'Y*�z�K]�x��y�O؟w��Q
�'�E3�l3v;�,�T�]�%!B�	�'��hM�A)X�fO�
_����'b.�� 	r�� #���M����'\*ũE��:�ȹ��L�nl �'��쑈3V����룥�	�y�kȱA[x�)�bR8!I��HC�� �y�Nڣ,�H�Dj>01�1K���y"��	(�E钫X�V�0$�K�y*QK�Hq�K�+zv���!���yR,�Bע�����u2�y���*�yRL�R�V�Ҁ���@���攎�yr�'H�(AaRȍ#i��`���y���M�c�Y�O�MR��O��y���B�k�B_*a�Y�PnB��y⍚{߈���+���qs�" ��yB�C�?���)��K�x �b���y"g��qFĀ:W��o�����4�yrZ�|S��h|(A��$���y�!Йt�,�s��L�f�`;�߁�y�$�-K��銑`ǫbj\��Լ�ybGґwrԉaeE��Zr�"cI@�y��;!DY[���'*���$�� �y�/����"G�Y'V<<Ak���y�	&vi��l�-]c���l���ybڝ)��P�UoI#gJ�۰���y�錇;��p:U�וp��qCЧ'�yF޹	]ra��WuZR��NG��y�oC�
�`��5jE�g��y�*Ex��F�^�CX����2�y�H�r� 9��c@�ʁ����.�yh2*�H���OH�� �<�y
� ��k�	arf�p3oҜZkD���"O�Cƃ9�@�c�gհ3l���"O�,�S/U�U�0��^�ok��`"OB�ɲN�-.y��Ҁc�(\*��!"O<њP��%A=��Ȇ��?{��17"O��{̦~�I���g���z�"O�$13+H�%���v.K�q�$��5"O���q��>�@@� ���c��\��"O�����V?P�R�J�LQ��Zr�D>�S��&���!���<HE��H��8C�I�+����%_
&������2�jC�I�L*:R�/W�l����i��xB�>
�Xr@��d*��
r��f>B��)~oRX��O�l���ԯ�<^�C�I3
V4�D�9Z&]h 4��C��;}>*���%G'q	�놌�/�C䉩t�QK��])\�(��� C�C��3oÎ��C���:��h2cX�C�'*�T�T'R/}��E�J�)�B�/X@E( ��/84��9�ˇ�B�B�I�u�`�b��7��m���.W��B�	�j���c��%/w¥(��A�aNB��#�0��㤑�y`�FfRwB䉞9���+$fY'_�4Y2�׽l�C�	'_WD��^'2�EW�7��C�I�U��$���5|��h$"�2/bC�Ɉ@�bXIV�=`���1'S�|(C�ɪ�"Ш�
_��xZЈ��C�?������bF�$r���	��C�	�Z�z5XB��=fV���F�4|�:C�>hI�4��IYtD�p�̸N�(C䉘r�nM�C�,"Ph���'��B䉞R`��a�- H=.@!�̈^��C�	3H�}v�Ül��J@��8��C�	�I���z�
[����Ĩ	S�h���$�	-S�X� ӡ�'#�l�+�ɉ�n�jB�ɧPr���&XV�+��Ƃ�.B�/�y5`S M"�<[$+�*B䉶�V-�7%\2+˨��f�&�C�I}03���u��\ 2
E�m�C��jΐ���	{����B� �C䉀A�\b��!(�h�IB��
L�C�	�\�C�F2E:�X`j\(�B�I7����kğr�EQ���aO�B�I�jq�Q�Qg�?���{�I�H��B�	�N�@���KƄ7�\��kI+�nB�	�ka�I��ؤm<���ـmRDB䉊/]`u��4��%��@��<B䉜Sנ�Z �E�S=��)&/��hB䉔S#�-�4�O�\��}�@�)�^B�,)��(��r�F��T9KIxC�ɛ���k��T>~��5��e�lC�I�Pq�8�C#	(F���"�O��dC�ɐXg�S���1\�t����C�HC�	�K�0��e�0hih��h��]�xB���1�m��b�*T�Ci�W�B�I�I�>Ea%ǚB5�5a�F^$J�B�	���7C
c֚h!�*ߧfV�C�I FC�����/r|1�͞2=�C��:x�!��u�Px�G��H��C�� Od���$R8*� h9PZ6C�I�@��5 jG�.A���V�:ADC��R�h�Q���7d��X���F�C�ɔT�Sb��P'�9�J)��B�)� �U����3M�n���̿.g�yY�"O�0��+����\�D]wMV�KB"O����힊h�-s��"G r�"O���1E=��	`h߀)�4��"O ��s�.s|4lb�#6�Ha�"O�(r`A�/^b��U�ͪ[�֭y�"O�8�bh�*]]�x�aD�1� �7"O�E�ul]#_0�0D�0n�w"Od�i�ߥ<~��(@� �B��"O�ʑ#��p!�(�ՋV�>��V"O���Ŋ��)�bu���$Z��ms�"O&aAr$�'[M8i�M2�Z<��"O �ň��Sf��9
�V@s"OxMysֹuX����

F>ͪ�"O��;G#�)�l)R��h�^Q�"O�S �%9=������Y� ��"O���5�K�K�����\��0��"O�!����2�lr��)	
0	�"OV�P-F�}��X{�	9$0My�"OF�Y�n*|�t�{� �Fxyqt"O�T���C����P�V�!n�2"O��"�� ��f�T�8�M��"Oz\��{��a�f"� �ځ�"OXp�P)�;�\�� �+G��)+p"O:��b�ȣn��y(� ��*ϴE�g"Od�SfJ j���`����"O��z�XXzp�%�.]���Ru"O>��V� 9l!�EËkz��P1"Ob��5��3�tд��=]\�#"OV�#g�d���@��ƥ|���[�"O Y�4���i@�����3K侹qS"O����� (z���#�P&<{��	!"O6K�b�=����N�"w��R"OF���#�j�-cW�%f���9s"O��	S��Or�X��A�u����"O  PD�"���9�E�BI*�;�"OD���P�!��C5�?iB�Q8�"O��,�6�N|�і4;����"O����(8�����-7V�+E"O����M	n������r%*�"Oum�1uNZ��f+�En��*�"Oԡ�R
�3 p���tI�-3���d"O�����R�y �H��*���A�"O��2���\In�	!ڻK��A�"O�P#b�*�TӁ5�"�B"O�d�ъ�*^�^I��*��H�� ��"O%���B�y�� LF��5��"O�	`��'V�����{���r�"O� y�f��AQ��r%O��t|iw"O��siA%;y-3���a��u`�"O�s��ϟX3��ZT�I�=:P��"O�*@gL!W�$����H�!���"Or��u(�I�X � �5>�v0�6"O��!d�X�&�q��g'T��"Op��bTgve�g%J��"O��*c)� 1�� �._j��"O���'�
w����K؎\Ι��"O�`�Q�]$W��]�T���f�|��&*OL46FE& S���U8"d���	�'�v8�©ӄ_�i`!g�6r:�a
�'@\��,߲:��1q�P����*�y/�t�HʃG�xX;נ
��yB�@ \� pU�ʶZ60�@
�yB��KQ����H�Q���[5,��y
� ���#�� dJ���� \�.ta"O�9���ׅZ��QR�ˏ.��dI "O�(���'}0[t�;}�*t��"O�}J�(9J�� 2��F�ۅ"O���
հ6����[6+�Vq�"O~�J2��+y�> �]2i�8
�"O~��BT����RB�X )����B"O���8ZC���'�\{��&"O�����˰��Y���c����"z�!�W'qq�]J���4_p1�e,�%(�!��b��T�_�M?���@�T�#[!�D&P�[S�@'BΤ���)/vI!�d�d�l}�'+�7u����*�!�͊?�����?i�����6%�!�F� 1��#��лU$аǩŷ]O��d+,�ՙ�B�#]���)�ND�<9V6�����-���r.�c�<� �Q�����b�&#�A�@\z�<�e�C�/>�)�Z�~bz���v�<����O�XPÂ���zrq���t�<�UЬ��,����>x����O�s�<�
�<@f~��A��8�J�#��I�<�����"�QuF��E*j=�� YG�<���1[���P+��T�h`u,M@�<�K�C����u�Χ�F�Ӷ�{�<��/evY�bC٥�ح���y�<i'�A06����	�r�`����^�<�p�A�d�I	���N}����@�<��Ç �	��n '@�0;p�b�<1ҁ�`���`�ᖹs6 +��V�<i	�7|��B��id��Q�\�<QD�յe�W!_�2���B�m�`�<yIY�Q<j0P7���!�J=�5�DZ�<Iu����$B#NUEXE[4�T�<��+B������&g��q#���U�<1�@Δ]D��	�n^$B!���"IF�<�� �L7��(��;���qC��<���T�fՆB�MP�Sn�� �YP�<�h%[�RT�0~l�a�!CI�<���Յ$:5��]-n�n` b�G�<��">c� �I�&6dƩ��n K�<ї�Ɍ��w!�8��� Տ�H�<��L�L�����ny`@@Z�<�gf 4f���ȇ�/D`�å·T�<!%L�g8R��
��H�6�K$��M�<��ԛBc�8Z�I	�r*�8'@AH�<1F�L�6�:�C����F|�u�,D�$�vf�O�dF�=F(21�+D���ѯ׬X�x�a��2�<3�f&D�RF�8Ih��BÍ3�g&D�p ��J�<9�Y��/���@;`
$D�$JS/�|��(P�/ޕIE����"D��	,�"M��S,�*E�HA�7/>D�8cC���+�P���-�l�c>D�D����K�¡k� Y����s��0D��b��u*�1b�Gy\� ��,D���������� �u�j��Af,D�90�׶q�~pI�F�"��51#�=D����˗.2�HdH�F�w��1	��.D��1�"�FN������M_z�xQ�-D���ԃ;7y�ij��Z�tp"� ,,D���UD�H;e�5��
I��e )D�D���_�+0R��!>���C�d#D�Tbu玝q���6�i���+�!#D�� ��4 ��>�D�#�kZ���"O\u��_�[Xbhp��C�;��X�"O�EiDmL�[o+"
�*!��m
�"Ox� 2�
\J�ׇ�XYt�`"Ol�1�@İG�3fgB�`"8�!V"O���M;4����9L}bI��"O�!����� �ADLx���"O���
ő'P�M�ҁU�/�0[�"O�H���28����*����"Oh�����'3�E���d�|D��"O��z�_"�^X�
3���w"O�HҠn<�`e�t� �CFZs�"O4u�EO^����v� �;�yB�"O���g�Xt��r��H&~2j�A"O�`��-�PA�
�:`�"ODA��e�	^j|��$���i"O���@�°I!�a�T���j"Oܰ�v�
2h)&�AA�7iψ���"O���JM.2������h�"O���`��.���B�' $�V��B"O��h0D_}�� fo��Q��"O4M"r��Đq�DV�'�v�`�"O:������� za�:U�
�i�"O��{�Ju�0���/�+��"W"Oni��
�4C�%�1�}�
$��"Oʁ�BÔ5,zy
4,Е�؝�'"Ob|�G"BW���R�S�:!��z�"OT����λS�|��À6M�!Ȓ"Oh(B��=Q�)!!��� ߾�A "O�<	�L��XH ����4=@�z�"O(�RǯԓY�l��%�.7�)��"O�4�S��|
��1P�͑x"zyf"O6\# ���]k�����^/ �T��"O�q��B'2�2L���'�H"O�:qEN)�F(9�ŋ�)'@rt"O��C�	��P���,2���"O���ֺ3 V,&c^�A�X���"O���@-98L�Ab�#�RMӀ"O���[�^��}�%�	~�Dh[�"O��Y%e�R���s�CZD�u{#"O��H��ZCh^	
1�ԏ?U�$+E"O@e�a��4��8�"�.l�Ƞw"O��
�KA"��
Gl�4\�&1e"O����R��8����,�<�@`"O�M9'Z�`>�c ID2l#� :"O�����~��������\��"Oܴ���ԒH\x��%Z?
-��"Ox�r�hZ*T(ش�Y%(~ibB"O�Q:���4�(�;�	_2�T��1"O�!�"��9I������9e	�q�"O���G�!d�q���.	^�[�"O��Џ5��A{B�B�F���"ODK��&�4�0QHMM茬��"OLqtLLH��r֧��%θ+�"O��3"mh�f���a��"O8�aH�@�.E����'
�*��!"O�5�����t$���K�6�&iHd"O� Z�� �zO�t��7�P�k4"O"t�q��'b{ĉy�N�/7�4�a"Ox��̌-z���dd�'|��A "OXQc�l�7��x�BҢU�b�h1"O�B����ph��"��{y0�["O��Y�(��K4�����?Ft~��"O�<��n��op��!3�R� ���W"O� ��5��5EU�XQ�LܥS��(B"OD�!m�	
j��DE�M� "OR�1U/�8k�*d��%� ?��["O�H"6&�3����ԣѨT�TY"OD �閥6U`@a%EX�a��� "O�!
��/���s�я�h�h�"O�Xآ�G-�BA���Y�48l*OU�G�G�@n$����ܛq��'`PTi��B�m{��*-�$Q�'n6Ib�V%�$���'s=��(�'�5{��V�}9X�8�@tX��'�\t;ԁ�[��9�gF�Z�>4��'D4��1���p_� b���V����'���b�E$>m,����MU���'��Tʖ���9xH*!&��I����'��T,�(q��Z��;�X��'�z��I9�"k��ߩ8:���
�'܆���ʀU6�8��哉d�$���'tUȠ�^,3���k#�����d!�'|"[�&V@q��P#?����'N�Ȱ�H�)k m(�JO*>N�1��'32�"#�,9ϼ�
S�ۯ	�����'z��FJ��^�V�q⡗���]��'�f�sc���M	�\�aͅ�Qf0��'��2���)' \ɡKܶ 9�%��' ��G�J��P!-�g�����'�P����p��0�G�I�����'�4 g̿J��7�"~��U��'ے1����h@����?o&:�(�'��	E�ė�R�2�a��9�'d��a�P�@�[G�vQj�'w�0�c��X�4aȞKH­��'$��`���HD�p��!pά��'UZ��U-ɴ@�0u˗iV.~��!�'�Y9�L,{s�8{W�F%w��K
�'!��fTm+bEy�,#@�R�'��j!d�9m��ѡ��{����'� ��j֨��1�QB�|Cfѓ�' �48�荱*s����@F�voj�[�'�x��C�RwPd���?l�*��'� ���GB�MԞ����H,��8K�'��X1�o�5-2)h d��]A8ɒ�'B���X�BN�DQ0�޷c���I	�'����@X}�tK���?P����'l6�����R�X�xGg�+H��|j�'0�y	�ǉ$Jz���k�6L2jE��'r�I0��J�&���RAŎpQ�p �'�xm��k��$ה��%B�c�e��'��7?!�Ż���z	�'䄣7)@'a���i���8�v��'LX�F�W9�X�A�	f��r�'ծ��S�FC����0`V�N�؀H�' ���!aʴx�����bZ5��M��'a^HkN�#��N?%�Uآ�͛�y�S�L0����	(��0�*_��y���E���bʔ�,Aj� ��8�y2�Q&��A��D��t8QbD��y�h�Qfv����f-�(5�	�yr%��DE��Æ�_[֩c�C	��yb�70[8կ�*!���fCߕ�yEU�m��#�\%w�|�p��B�yR@�9 e��� 6!f�=����y¬�
-ĜE 'ܦ@\�a2�ޗ�y���)c4Q(�-�
��Yb��y
� L�#��/���+��):�R"O��t��x�<�xp)�0YQ"Od���KݢA�.���HP�%�ȵkp"OZ���bB�����J�`���"O� ���|/���T��=�&�8 "Oȹ�T��(G��	cIR��<� "O*����Z0A��XA��N�4#%"OnLrp�ڮa�ޱ�U�F��Df"O(��1��[�br$/Sp7b��A"O��.�?-Nl���[�C�$C�"OJ�@%n�O-�PY�l��6RIC%"O:�(QB�e(��5Ŋ&N XP�"O4�-#*��h��%�h��\��"O��@2�ӇP��l!å��+����d"O�(�+ȯ���J!1��E"O�!B��5/���G�DAK��i"O�pp�
R�Z�0<ⲨWl=~���"O����i�(y�������-��i��"O4`+q�G3`WL��s��8d����"O���cH8S�JeRF��l�.�"O��S��˼g= ���N�&R���"OJAP�h�H�b1�O3p8�B"O�YR��&/�q�B,X�:)���"O&���l��/�h�,��&���D"O�<�v@�%*��Y�ī�6

d�8�"Ox̣�G��z�J0��>˄\��"OΩ:'L�"N`ڙYD邚D�hM�$"O��q!�<i8N�Jp�@"���H`"OT`�&��� c�e:F�J��"O:��d:@^����M���"OD Br͓2?M
����)S�X�"O�D	�"�P4����h�l��"O�T��OR8�Ʌ h�Dt�'"O<�����c���4d�P�:"O�|���^�(U*d/OJ��x�"O0��ū��UB�����o٪��a"O��0˛&Z�9�B��2]R,��"O�\��j�~ޤЫ�$����pq�"Oh8�N�Pӄ� r$V�v����"O��y�AH�s�����_:|��<� "O�9���"'s.�h���c�yaW"O����儊���HD`D�����`"O=�U
"<]��I��\���`�"O�9#R ڨQvV���H&!�	("O(U�&kM�t����(�..��	h1"O��K!(�pɦ��� !Q���S�"O~D�H2X����)Dn�qC"Oh�`��3�*�.K�t���"Ou	�$	~-�v͕�di>ɪ'"O�a�f��?q�"U�7��]tͫv"O�DCa��G���5�ϨF�t�i@"O�!����*���  "��[�L��2"O�T��E�$<j4Z�`_������"O���&��j�rT��
�Hp�"OhȈ�s� �!�&]�_q�0�"O 	��4u (BT��R��iu"Oey����M��A�('k�5 �"O��
��ȵ@��QB��	1`бIS"O �j&LD'uc��@��� AМ��"Oj�+�-�F�k7e�*>&E�"O0��Ehٚo�셺F�6z��ܚ4"O�U0sC�u�)�6�X��N�"O�0�eѨ'�K�m�=1cZ aU"O��1���B����C�zC �0S"O� ֔�mϫR�qz���8jg"OJ� F�L%h| �y��S�v��"O�(3d�.�,-���ɮ6<�,
A"O�H��)�7q>�9S��d!�Q�5"Ob�+�a�)>/�Qr�
ܾL�l=@�"O�<J��B<L���i�(�g�L(��"O�!|��`�E�]�P���"O����o�*��(�%�D�ȺU"O�$��K��^�]���ګ]ʡ"O]�q��$h# ���ޛb��1�"O:"�-Ԉ[���+�F�aQ�l)P"O�MR��Y5D�!6j�W����"O�$�vM;'�
�*��7t���X$"O��`UA�2w������)M�:%
S"O�y��	߄3C�S�S�t=��"O�9��Ȁ?J�p�� &�F�@��"O0�c@D��Q�RՒro�R7�2s"OLQ�w��LQ�(�"���!"O�eˑ�Z�\���J��� �"O2d���1�le��
 N{ Y��"On�5�>�J����ޗ^��,�"O�� ��׾l<@���U��љ"O ����I�/M�$�S�Ȼ�
QF"O����#߯,g�Y�́����"O�1i�	�2<c$M@�8D*�"O��i�	uN!Q�k�O�LD��"O�i��m��M��(ZC�G[<i+f"O�|d�I��z6��	ozq�f"Oڰ3�R}4%Y�h�Gk�$"O�ˠ�	y��J̷pKp��V"OdzV�x�.$���-"BЙ�"O�ū�J%�VQ�%� H	�"O��"�D|\]ত�?B;5�"O�Z�OP��Ѳ"�?,��""O̰�TeG�q8��
�A��O��!"O�i˰/��-h�$nH.Ȥ"OF�	� QgI�����X�l�U"O�����R�Q�b�@���y�"OL��4.Ӡq5�RC�$�|��"O|�s��
R#n��r#QBez8�"O*U	�jݤ7�
����֒AZуu"O���စ8���W��#5ޡӄ"O2U���ݴpf^���-ڂ-'ȝY�"O�(���_aO�d#�\K\��"O�@ۥ��.;
 ٨��;<6�!a"O>U��"��k2�=Z�#K�nNt���y򧒔h��\ɓ�N�An	�y"F�;��ӄ���
��q� h���yɛ:KN�Y1�Wo��$�rS��y�"��7�'$�Zp������yҪ�@��(�!�d�Ӵ�٦�y���I���f�DV�Hd�l��y"�^�d���iG�N�!k��Z%�С�y���8�̸ꔢ�B�����y���[����!�T6$������ޙ�y�ę�9,F����%I�����B8�y�'�pO��h�a �X~� C#���y��λU!���"� =}�f�"�U�y�O�?I��7��'"Q����5�yB��PY��""��=r,�눀�yb��uu*-��K�9DF)�`hY��y�T�qP�t��K\F>�zу��y����ulb�j#�֭ZĪ�� ��y�A.>HM�V�=+�K@Č��y
� l�0fi��Aum�EГ2��M`T"Ob!I R�!�H칤��Aќ
�"O�E3Q�5M!�	�V@H!G�v�XR"Od�y� �7�V�aR/��uJꍈ�"O�$����v`�߄v�Ԍ(B"Op��դ��Qn}����"B�ݲ�"Od��V�]�L�d8�pC+4Qz]�@"O�����s���vB@	5I<A�"O���D�_�o��`�2�6W0t�"O�Hy� 4<"���h.�U��"O���$*E�k��5��4SB"O�R4$�Ki0T���ֱF��թv"OzTٵ��=W#@;�+v��͒�"O�4��\ j��H�6�%x���q"Ojuc�8 t����V;GP�Q�"On,��Я?�.�;�hI4��1a"OnL�3��>F=X���*�ex6"Ot�� ߱F���:Wg�Qo@��"O��x aM�w�,���M�*mL�"O�Yu�]4jMb�9�ǯ-]�mb@"O�iK�BݍJ���i"F	-v�T�s&"Op�#=q~�\�"��8-�a"O^�R��#X12�@�-zo �D"O��
��L��\�.�2h��1f"O�������11��Iap�8""O��"QJ����l�숾}慘"O6<�q��o:���l��?�<	�"O� �rA�k yi EZ7a:P�1"O�@����%g,$�bI�d�ʥ:G"O����)�� �0�BENL�])���"O8P��
ChR����"�tM	�"O���S�_%q)AJ���-}ǜw"O:x� �.d�]��Γ�	�#"O^���.���..�����"O�h_�P�D팆cpDI�@"O�)@�mu`1!�e�?ČA1"OR��F	D%c"��DW�?��|�$"OD
�/��'��LK�D-4���"O��j7�C�w�|$���q1�-�T"O&P��%�?b*P���~x���"O(1�Q�8^L�qN�<oJ�YS�"O�0��Ⱦk���1��	�aV��CG"O�dX�i�$�p��H7f��"OܰӠ��09�8B��=Wx"OtPᤃ�?�|Kpd�A&	xG"Oz�$�X�ސ5;��Ӏ6d0�"OD����?���%��:jH4��"O�m0�&ܖ���Q7�7]�13�"O�Q�V.<y�a[3!��JH��B"O�]�&�22T�R��<?1��"O�$I���<x�uçK�W���Y�"Op�@mI��d0J���k�R(rB"O�4�f�8-�������z@깈""O��A6Y�8y�fN�l'V���"O�#�ɉ �NY0���-�%3g"OhU��"�xq��@�p�j5R�"O�`�  �'@�B�����	ΞI�T"O2�g&�c?X]$�׹+��y!�"OL�{ב7<���]�K v�i�"O�ə%�Ng=�]���������"OB�0�^9C)H<!���:Q��Q�"OA���{�Z�"E���g@0��"O@���%�l�1��C|�`"O��1`��9�!z�P�E�|��"O� l(�'��K��͒�!&}�٨U"O�	x�'N���Q!��ybR���"O�,���>��U;'�VLF��I�"O\�Fo�U�ڝ������>���"O\������
�\A��
zf<a#"O��A� �o�Z�0�,I:^a��h1"OX�c%��J�$Ԛ���1�E��"O^a� ��eQOڃD�lE�a"O>�3� ,�l`��%"�`��"O܁��X,ez6]��lȲ"�`��"O����j�*. �0_�Z��"O0�*p]6Q�F|� =<�2e�s"O
�x�҂H�M[�e�4+�*-��"O@Y8WoFpL�g���O�Ez"OxECb�1p
�d�	g^�i��"O�A�&�X�qv��d�. W����"O��;t��I��i��� �@�"OdA���h,y�־`����"Oz%;7�T5P�۴a��@4��;�y�H�[�P9ʂ�ЈWZ��P���y�nB�,а����R%JD�G�J��y�Mº{�1q�ԀJ_�Z��ZB䉠v9��X&mԝO������D�B�	�\�|\���
V�t@�@U(:h�B�I�'�,�P1a2uЈ�SW&ΠEiBC�I*^��)g��U�R�'NJ9t�C�	�ND�t�T ѫ,J|���r��C��%U��!��n��#S<8H�e?7�C�I�H��)áK@CD<C�!2P~C�	#)�I��+׃�$0�e~C�'tվ�@E�F~����a�_��|C�(0���XS,ѷT�tYg���21�C�I6*������d_.�{n�&�dC�?#\5�@��XXZ�a��#)8C��.ZtX��Bn�/5n.P3r�L�WzC�	�L���ိC�WGT��lL{� C�I.?|�����L�t��	v��B�IJ. m8���Ƀe��8Y��B�	�y�D���\�fR��B���E�:C�!<ВQf�Q�Y�^)��N	�*C䉥x�lɰ��6E�Z�Zf���C�B䉣}Rdi���9<Td=��'ťi�B�	,W��1�0�K%H�>�I����NB�	�W �
��~���r�F=nJB�I E�,�k�h˥=�xZ��B(b��C䉲/�+MB�t��Պ��	�
��T��'dԌ�cW�S?��AI��-3�Ȫ�'4��.�S����k�*'tN\i�'�J)Jed֖8��()v�4��'���
�J�Mb"�d�I�(|�z�' ���q����m�S����5K�'ޮ�y7�D�@oJ :�D�I�"���'B�'+��DY&5S�ǘ�<8���'�P���!��%�#��K�x$��'( t�u��_o��+��XPH���'J<�ʅ;��ے����m�
�'�.L��!��P��)�r5��'0�<����+�NL�!�ҟ	����'�J����]����L��T2ЉK�'���8udY�9�TA7j��\��9	�'��±D��h����[}@3	�'��̊�R��E��~N2��'�Z¿02�-̀`����w'�y �sj�hpF�T�C����ʨ�y
� 4�x��O�K�$a�`�ׁTG��C3"O|� ケi9$�g�ނMW�ۀ"O��yq��M3hmx'CU�Qh�e"OR�X#˷J�&����39(��"OL�WX{�u '�l=f�f*O�5�5��R.���뚨OJ��'�h��-�Q:���jA�GL�K�'�@����5U�*H2�A����S�'[����׮�R�u�����'ͤ�+ j�	N���U��!}L�;�'W�pі�Q�9��T1)�
�'�P��"�D�g0�p�ǳ$�8U�	�'�i
&h���IqB�e-�P1	�'����hs���LD�b��0�'?R}	�ɇ"��$30#�S��@�'���ǠW�t�t%����!J�e��'
Rc�]0��=��'P��Xx��'�|���U�%u`P�5�3|�>e0�'���R�!�H��+�*Dp�x	�'��u�Vʃ6)�@Y��'O�>7h	�'$PD���V%._�$��ʏ9'��!�'��e  �2�1��m@,~���'~��hd͊�3X
�h# ��81L�9�'�V��C��wY���nޫ*�XZ������5�(s6� s~��0�4D������2}Xdc��>�S3m6D�(��ͳrU�d����XS|!�?D�x����4�R�Fk�!	��n=D�L%�_p1#���tZR*8D�$���ǌR�Ψ(bgݢW��z$5D�p���}�t败�$j0D�/D�2	�H2e Xn�(���g0D�{�k��y�|0�IB�ZZY���1D�$�%ٖ9l��*�A�{�X��U	%D����gB $���d��!�,�Q�b.D�HA �O�g7�� �e�;)_"���1D�����1ة��#JL�e;D��S�Ԥ(`	G�7F�"�8D�t��'>hr�"�P�L�p7D���/!0M�l�-��oq�0�A"5D�X�F̀������!k���D.D�T����Pz����w`ʘ;�O-D�����t���m۹��A �*D��U�	on!sƏޞ/}0��Q�+D�\	S��+�L٫rn^�p�^�#f)D�lĀ9h�r�:5mۥ-Ð�6e4D��#g�+aڈ4�E�E]���)'�&D�`�W�J4Ot`;嬁�;�@�%D�0Ӈ���F���߾E�:��k!D���eą��@T�0�X��,�y��$D��#qN�N=� Ht�>\�Z��!D���d�G:b��8)��Ð{Č��$D�̂'���<�! ��@D"D���f+��u�x��&P�P��$D�̋w"�7��xY�fLe���"$D�{��ȗs�h�N�0"�8is�=D�x����G.�J1�H 9+����!&D� ���Mn�Td!��˱t�fܳ�)D�1�ა$�Ĕ�b��'_� L��&D�� f&VZq1���
@�\s#&D����e��P�ƽ$_J G�%D����S�/h���#-R�G",H�� #D�P�roKiR��ʐk L����l"T���A/�a���� N�(�n�{"O� ֔#��O��8X�D��:��%"O, h�+�+Xyި� ��^)6�ؖ"O�m��`E�"�x�Ba�'/��� "O�
�/l�!�j��L؀"O��1��Q*1k ��T�����"O����5�ޠ0�M��\�: �"O(a�!.��@hm,r�\a�"O2���19j��3 -ÕvӾp�"O�PQ��A�*,I9r(��q�"O��aCM%s��,i�.�@`�	�"OD��薼f�"mQ�h��Id�R"O��a!]�IH�Sp�/�t���"O؝yC��V��ձAf�|�u�a"OB�v��H�])G�4 �rL��"Of1��2���3�C��]��U�D"O�-�����i4�e0�a+G��$0&"O84:
[���T#�$dxR�k�"Ov1�b�,�L�S�ă�k��Q"Ov} e��^w͂��_)T@�8�"O*i�������	���Ydر"O
%'蒾���x�@�:C�f�#@"O�dS�����R\�،Xu�-	�"O՛c���uw8�K6�@�o\j�rf"O&�3�눻���b�W�"E�Ih�"O���v͘5�XY��
=
��8�"O�+�n�o�f��E[#D,0�"O��H�F)Kl���ҞE��1�"OzTA�\!M]��B�)�45�"O��p�$(d���u��P�ni�"O�a��O �4RC���~���@"O
Q�$I�E
8���LOl��`�"O�Q�`O�(y�`��ѩ���b��W"O6���,t%���E����)�@"O�8��@��v���RJ�^����"OxyyT��A0���qH
�9����"O���2o�*�ؚ�ܥgy$� 0"OJJ2jO<;$��J��oot�!�"O�Hz�&
4����ƛ;ozu�"O�бQ��D�9!�'d���"O�H
��]�(�@�P�r��ks"ON���a[�
��y�,O!z<P"O2AC��@p^�5�3,=�4"On\ 6Qgd!C���s�8d�"O^����ĜUh�8�IӃD�P;a"O��c`��

���%)ۃ\`��"O��B�B�p�T���
E�2I�q"Op����X��a�"�	�ə�"O���ˍ�V�����S*$��=�%"OHta��lzJ�Cto�l�Q"O��b���5�d8(�.
j�b��"O��i$.P�bY�5���T��i�"O$����ѥ/��1��+ ?0�[�"Oz�o��4WV]��ӈ��RS"Oބ
#�I�1�Y�.�K�"On᫆�<I�,H�գyo��:�"O��5�Tv��1%i��X��@G"O��@X�G�0���W�9M�pi�"O�쐠��5�*xH��X����PA"O$<�07*��u��#:�,��"OȌ��.]�:���Z�'��@!v"O@��
F�|[�q���*y�� p"O��bJH�c��5�s��r�j�"O��bHQ�~�2D�j%:�(p˗"O�-A�$���X��3�\<�HEÆ"O� DPb�X]?�43p�ũ?��Ax�"O�s�+�J��W�Y�"O�i�nG@;�35@��9"��P"O�H��!Q�hG��A�y'\�1`"O�E�5G�3FI0q��3A�0��"O�!YժU�:TN��+�&y+2\�"O��1�4,�95P�g�F=�Q"O.J���8�he���3:�Jm�"O~��"Ð �@Ae�fA b"OДJ�з+7�ɘ���/���"u"O��
G(��n]xߌ�z�"O( �����|;�/��q�>�pA"O�i�t̀h����ǻ�
�h�"O~��6�@�>L���_.)�*�# "Oh�[bNӰw���Q����x��{"O��K�.P�%4�2�ph`"ON1��/r�����kB9�2%�5"O�õ�;'{��їʎ�,�X�A�"O�4/G�r;hT�F�]�_���v"O�(�Z8dH����!�;u"OF�z�f�-a=���_q���-]d�<	�E��ATK��\�SƄ�a�<y'�1d���؀��?g
�SA�^�<a�cK�-���ϛ�"�lek�͞W�<��t[
ء'Y�:}j�±!SS�<!�D�6Wur�I���Zdb�L�<��a�;2��e�9U%�p�3	[E�<��o@�#_�h�g��*=��+Ү�A�<���ҍ!F ��E�1��<�CDB�<1S޾s����Md�蹃�F
j�<�Ѫ
�@Ռ��(@1}!��q��b�<�E$[�0R��¦�0}r�; d�<�R=m�B-���|��L�v
�F�<�v���)�t�[ă�6
�L;�Μ�<��Xi��Ȇ�	q�r�0D|�<q�J$H�UB��j��[��,ܙ2g
9#7n}�3�� �r���k�x�z@CH��d�����F�$ ��oI6D[�I��S�f {S���W�����z����ƌ�:T��/H�Jk������+�X^�8 h��DҠ�ȓ<1�Y��]�>��(��ĵw�^�ȓX���˴��-Z�f��0��4����ȓ!�� 7�K��Bt��gF-w�E��r�,q�3��hG�Ԛ�P+]h(݆�,I�A��+:?�T0�V��)����|���[� ��}"r� F�'"2���ȓ �r}W+)O������ąȓl��G�wsxqj���#�P����aB��3rx����4��<��(%�� q�D�X��Z~����ȓ`ђ�I�'��@�i�����~jT�Ƈ�/*vfu�G /�8�ȓӲuCQ�ݽx�c��1�|��;-��DA z�*4�E�M+�ȡ�ȓp��6���_�i���#}2�Յȓ�T,�q��S�.��1��8xL�ȓ@�J�gV%vv��゗�9�&h�ȓo�.��Q@H+b�:P�C��:����Ie���pd�8� 0���F�'[�Ԇ�X����$��s�$a6/����ȓY��QB��]>O�zfJ�y���ȓ+��<	@'�v�:I�1�Pp�	��~0J	胮_!��L��L_��h��S�? 8�h�+G�̓a�G<��m�d"O������7"H�gяWǴ�;3"O�=��$RJ ��
�"Q�,�h�"O���
\��r��#0�8S""O���T�.A��ؑ�M�/�(غW"Ozdg��MS��ρQ��D�5"O��z�+�ᓒbE+:�z�Bu"O�b�i	�4�V�*$��%�xD�D"OE	dˁq}V�ь�fhN0�"O.�qn����;�B0V�Z�"O�!��B���nL�1	1wM��x�"OH�g-P ���ބC�53C"OL���I	�LZI���H�nc℉�"O�-���Y6�Ԅ²L�d���Q"OD5��0ilR8q�
^�h\��2�"Ov�r��To-�Qi �S�*�S"O�<����\��a����,Ax���@"OJ���;v|��2PA�K�� %"O�����Fh���C�I���ҡ"O��B�پ-az�Kd��	x���"O|��-�+%�
2%��� ғ"OHɱCX:`�NU�G�+�����"Oh�[ �
��0Bb
<�XP�s"OD̲pg��~����7"P�s���;�"O*�a���%�Љ4�ܑi��\	�"O�5��o+,@TA1BֵoyD��"O0���F�/r� � �'P����"O�Y#��A�(y����0o�U�"O���?mrb�XdK(KnD|��"O�d��
 $1������I�0��%�"O�Xk1���!.J�A��J�,�2��"O��Y�+O��QZ�敔f��hT"O]i���
찠�g�+;�B�;E"Obtx��נ���t�H�wCX�J�"Op�>.h̣Ce�5I*8t"O�y�ٻcިE�A�T�T"�D�"O���P)RF�Q�PB10�v8cW"O�Y�bG¤0��P���ץ@:�:F"O���g^�t����W/0��"OV!B��Q�K�a�mϟ}HM�@"O|l�dj�B�P��쎎n��`"Oj=��n֫>O�`�,[����3"O��A��+<���+#�r�#�"OT�HS�ޖ5	������h��"O��&��	��xY�F�d#�e3�"O��H�4XD �cOǉ0��|xD"O���4�� ?V��%EԆ8|B���"OP"1k
(o^��CA�pk��xv"O�Qہ�Sx� #����EB�|I�"O�|(�Ђ%�T�{G�H7�:�"O�a��(}�<�S��6�袄"O���+�ZŸ��51�rm�P"O4����:~xJ�L���$��e"OJ����*U@%�T� �+�"O�\�p�m�� ж��<�F$��"O�t���1"f<��iL��rW"Oh�r"�� ���:
�\"t"O&�ۀ� 6�����]�#�X)hu"O��&ө�1�vL��|�2"O����k��T���fkݰ�*�5"O��˓�<y`
i��銧w: �1R"Oh��A�O���<3���!ծ<{�"O�i�V&�Rz� fF��X�S"OX0���3H�<�fO�3�rՓ�"O� 4}XG	ηy��ܚ��:3�}��"O4�إh�"��(�2.�$Tz(遃"O^�Q��٫ZX�T�D��Zx�y�G"O~}+���.8EL��+�)��1g"O|��g�R S��;��Q>s��ER	�'��y�3 	� �����������'I�1�0�_Z��HD�ѸC���)�'>m��n��5$�l�ca/�^��',R1ڕ�-[��y"�P�0�����'�� ꘗ���RJ�#"dm��'�5��g�u����MX>� S�'�ιkD�"�`�3���<�P��'��t�'E�E���gDZ?ی�
�'c�mʣ ˞:)��{��E2-n>��
�'��@ԊE/\�hG��H|
�'��h�b�XaD��R�I��Ej��ʓr�n�8��^�D�E�3;�L��:�3,͚��UR7�S�٘�ȓ\|� q2�I�#j��ɐ'�G���ȓV��հ%��5i2�a��@��qL����R�C�̊�%�BT颦L�d)�ȓq���J���-\�	�t���j��ȓ }8�ʶd� �Xk�$4l@�ȓ���˅�N)z��<���Y9�D�ȓ`����T$`5�A�R�R��ȓCU�`�.T�)#��z�ϟ8G2���ȓ�%HWg�.�V%�Ɖ1+uz��G�x*$H�h�`�����0C�IP2}�BH�� �*l��m^�`G�C�I�'�<x ̉�D�(��Mm�C�	�\�bTY	�%uP��eFH[�C�)f�}Rg�^/A�FRc� c��C�I�3]<�c�e�[���0��C�Y��C��+*��U r[�`�0%E�~w�C�Ik�YYU�� BR	1q�0l�^B�%-u�� f�q�TYBm�&}�HB䉟`p��!W G]L�a�HąQ�B�	8����� ��]�eIטF�hB�I ��U%�CV�Qx �V	@�2B�ɘU�тcׇ=I���t��:иC�I�S��A��)aY`�0��%��B�� �x�҄ �Y�iP8[�B�<hT�0��D���Qb��\��B�	9)�$9����*���yWA �w�B�	GYѓ�#λ{����$� �f�B�	(=����ӥH�q�H-Z���1(�B�I
N�Q Ӯ��[�N|���a*zB䉲NH�g��h-<Lѧ�aђC�	�26�9������{6-�2vOVC�r�F�*� [ ��AcP� �R�2C�I��$�㡒+Z�DC���?�6B�	8>��x{qL\s�( S5A�b>�B�	N���##O��2!w
K9 �B��)Y���`!� �k�j��ɣ<�C�7(0�LA���_J���i�5EǒB�	&�$]�u�,���H#�ļ&�\B�ɏB��$�����^��jB�Ɏ$����n�r٢0��E]9\>�B�IoU
T#5͒Pm*H���\71_4B�I>�Qۑ"�|�Pk �.4nC�I���p�f�E)=��3V�Y�R*B�	�`�r�j:j����5JU�R�(B�Ʌ��Yzt����~B䐻��%D��0c�ĸy��]�� ϼlZ�K$D�� �t[@(ٵ
p� �CiR�
1�H�"OL�� �D]�~��F��}�����"O�1ɗ�u]���èJ/o |-+�"Ob��#�ͻg2�z�'ĄN���B"O�Ab��^���q��؆_�`�p"O"}s7NI�Q���baZ3-�D��D"O�8��T��xX1f�H��-�"O��h���3>�s�h
��*�;�"OR��b�A~�$|K79&����"Ođ��$��_`<�i�7^��T"O����	 ���#􎄩�"O��ʗ
�'r��|p�-X�!A(A�"O�a�U�K�Qb�,��˂3<�m��"O��(@��`�n�`f� �O/$4˥"O�mQ�텗pa}0G�4k@SE"O*��5V�h���D� dD�q�"O�Ӓ�M�"A���"��:
9��P�"O�%�шZ��8�ц"R'��X'"OV�"$�Z6�1+�ݬrŜY �"O�M2a�F&$�0q#���Y�\e�"O����R�9�BT�v�>/k�(��"OfK�e5�2��j S��a�S"O<3s惾Fܰc�
�c�����"OZ$[Dc֠"?@*�ٯ%�j�[�"O���'Ϻ	���P6c_Dwt��V"O��U��;YBt�xv��}��1�"O��0���ΰ�
?Y�b��"Oع�b.L"$���\7�y�"O��lI;LM\ib��ÍmEڈ`�"O�	Cb��u9�m�nܨq�~� "O 0R�-D�h<)�4H^�ln��"O�}����#�""��',D;�yg̘,��7F��C�Bm��N��y�S�JpDZF��>�\��	��y��]`�YӬ�����;��],�yb��Z&�@G&�$m���ڷ�K5�yB*��Z�.9�b�k��x����y"/B�ye�M�G�mtN���?�y�m ����W/�h�^�`���y�̘ 
���r
ʂq�>I 1/��y�(��'֩n(���Q���y2jA�V����gp9�B�<�y�ʋ�q�h�p��vp�h#q�0�y��@��He����q]H,k����y�l+Uc���f��h��8�yO��l!�ѮǳYG����]��y��L�`H��d�%P���%	��y�IA%Zri��M��>�D��'��y2hN
62Ah6��$5��2���y�#�����D!`y,��ڌ�yRf�{���r����^�pi�t�� �y�Ŀ}�H0s!$,jV��T�4�y�K�Ze���ą�x`HA-�yR&́0�0,C��{v�He!���y�͐/D�����;��Ѵ�9�y�+�`$ЛBo�5C�S�A��y��ֶ7�4DdR:>����ڇ�y�Nݩx���r�3!�	�ԅ�y2j�|��)�Q9�\���]�yl��l�DR��\�0� �0Ba��y�1o0��@����+� ����$�y,��lV� b�-�����ޫ�y�@_a44`Vȅ(5�X����/�y�9lr\U��ȂZ6]�$"���y
� ��R��џQdX�&/
Yp"O�%�r�F��Hͪ!�ݮT :M`"O�-A���0�g�F�{d�"O�d�$��Es&U3� �9qdł�"O,����0@��[�i�?-��@��"O��@Q�h�]z����@�yA"O\qS���W;$Y�r��(*l`q��"O2�K��@!_�"�!FLZ�II�*�"O�]�N�`z9���\�(���rU"O��ɃJ�.*��s@Lf���6"O\���1�(�ң�8	�H|I�"O;��Ɋe��5�1�ܕH�8 �"Oց7�2[���Z��N�	]\
2"O�m9�O
O�>P���ܠ�$x��"O��G�*`���q��_�B�x	��"O���\�j>:T��O��k���k�"OD��1�\=�JLZ�/HGE��"O:���!GA�,jխč&d
���"O��@�a��;�f�H��J�.w6�3""O��b&��D��q�l�)|���"O:ё�&�,� ��鋋a��҂"Oް�%�'Y^��w�])��s��IE�O|8KC��*t�̝ ��D�K�T�
�'��ъ�>{| �ɖ�����'j�T1�>U��h��>
W��b�'��]��N�y�N!U�%}^��Z	�'_� �g�/��5z$^�,�R�a�ǘ'� }�@]�Dæ�֦������x���+4��i��{��]��R��y�FI"�ĉ��X�k"�@-�ybɴ/_N4��i�aV<�J�=�y"%ؖ7��0�����H����ybi?}�v�b��Y�o�)H��ܭ�yd�ZJ��q�) ڞu��b��y�LJ"YB����
�ۆ)A� ��y�F
�
��hp��ٕf�?!�d�Gu���v�	�@�0&ݓ>x!�Z8{��I֌H�s��h�wD�@E!�DԼ|��(����:50� 㦢H�!�d �r���ZG��#3�,à4�'�a|��æ\٨���70�fܒ��ڇ�yr��6:��C��.AH�Ze[��y��D�������o)�艒����y�ǖx�k�I�g?<P�§�y�ͧY��}�6��_��E��i<�yrȅ2~`�И�h\7^���[����x�'zԸólȋqt�����%r̋�O�=E��j /{>E�S)R4Wd4� �y�	���ЫB���6t;Х�y"Ȑ�RC�PV�qȅ�ɞ��y2���;g��Q�i=h��_�����'���e�Ҧ���D�u\��
�'�&U�f�Αd+��� F���-�	��&��7E	**��Y֋�>Vt���M�&��3b�Q��|��J:�~8�� )WK>c�����*�ɘ{��I�$��� ɔ�D/R�C��"n�x8w�Ak (1��	�c���'�N�O���l��T��<�+��Z�.�� �"OF�PQ�ۇ}�Dҗ,ۥ$A���	j���)��q�1(�Nu%�i��˗,b�!��B�rLQ$Q
.+��
��^�F�!�� v� �Ռ0&b���@�y�!�C�%��H���)&t�7
/n!�F�y�.�2��5_�c��N�!�� 29�`�f5NIp�`�
��"Of��pI�f�����d��Hr"OȄ3���	��\�4��l���;�"O2e���W(ăQҏ\ET���"O�RS։("�+$*F	A.Vx�&"OX�StD�M
\��Hסz7���"O\L�E*ˏ���p�핿E>v,V"O�͹'�]mB���EJ��Uȵ"O�i�1!_�,x[��䊕�J	ɐ"O`!�7��4 �D��Fq����"O��cCvu�@0-A�Zp1��"O�	3��6~v��%�Y�"�<�qb"O�� @���v� y��d�1���j"O���E�ӋD��� #��9�"Ov�W2=o܁%!(ɘi�C"O���Ǭ� /���a���$���"O9ʔ�X6-����v�S���L��"OT����S�U`��3h�{�"OZ���L�����������l�"O�M�'��4�l�ȥ/�=	�`�"O�|�CMY+q1p̓aTT ��j�"OȌ�℅0��b� Ts��-�p"OL���B��\�c��f�D]8�"O����ȨD��a9!eR:H�n���"O�a��"�p-@�C�s���%"O����ulj��C�7}�HH��"O"dH�"!5�9+싎P�� �"O`�B��9���v%�m���[U"O�q@�E8x#,lr���izv4��"O$�б᎛>*,�1�dɻHhN���"O�ɺӊ�$�(�QM� ~^b�p"O��P!�$uL|s�m�-A�}`�"O�@�ը�&-h�1�F\��P"O�9���p�Zu��("z�a"OĹ+�E7l3X��에R�~�'"OT�25���w�4!bI��7֎d@5"O $��g�J�ǧ�+X���v"Oz�w�@�o�X��s�,F�]�"O�Q�P���IQဉ""���"O�ٱ�j�3y:0�0�HB��8A�"OD��$A�0V�@
�NO�in�9�"O�8��i6B��-��|e�%�V"OP�+uB�S�ڨ��,8U��MQ"O&�!�FZ�,������t8�"Od
�C��:�
�K�$G�b2du "O�!a ���Xw��L(.�)5"O$��n��M�(cV�U&�	s�"O±K7E?��I�q͛�OX�AB"O�Ht��<�j��2L�4<2��g"O�q�h^�*S�`�wk�#�@B"O`Ā�D�UX�k0�:y���*#"O�ٰ5�M�}�B�Qԭ�4 �}��"Of�c�̊�}��x�CB�h���j�"Op9�C�����@s�$8�4xs"O�1�$̀��!`ǇVƺx"O���P��*L�4�-C-X�pQ�G"O�hJ�!6xu�i��G�u��"O�+TM��Ljt��0
�"8F���@"Ob=�WI�Oʉp�Jضv���ȑ"Ot	���U/��8�iR�f\��"O�)�g]n���Ъ+6�F�1"O��͊�E)C���L�`"O<P���%j`����X����"O� ��5hd��@�)	�1�,���"O� �����~�0$��L�A$�X�`"O��Jb�˴�|�����FԤ��"O���V�I2|��HV��qd�؃"O�,k�!̔8F@�	�	��m�5"Ox����B,fPl���r�ܫc"O���  �'���8aX:Tn�i�D"OBm�BƜ�D_�$�L�U`r�P�"O�	 Ʈ��ڬ�f���7U�y�r"O��#P (Z��c��Ћ:A�&"Oh��E�Z��`�X��ۈ(*���"O#A�b�����Vld�H &�n�<�a�5s�xܸ���]"ti�R"��<AT!Z(���UJ�^-B��A�<is�ƃY�H�]J(T���L�gj$���ƸjҬ�ql1D�|����{y�}A��^>H��\xM1D���#�
>��)�b��M�F�A"�0D���p�ǂ*���;�Q ~v�`�.D�xI���*&�Q��hͩ)u=��+D�P�##�P����1d��c�×�(D�t�r�ƵY�"�O�a? 	I�a*D�� ��:l^�0��J&(}	)�(D�����N'm窘8ր۾s���F�"D��h�c�>Zϒݺg�ؔ(S�X9g?D�Ԓ`�K|L���U�L,�`��M?D� ���ʲP��߫OP`�J�"D��h�f��
LeC��\�[g:غ�.D��a��}�ީf��9����+D�" "ZqZP��C�;q¥:1
,D�4�F![�Y0���C*���Q��+D�d����2�51��65t]ـ*D�J$	V���%��b�h�gl-D�X�4��u�ָ�C�@�Y� ��7D�T� k�Ve �z�b�r��� ��0D��A�$]!�yʥ�؁S���K�(:D�,0�.�
/DZ�rF�7e��2�C7D����Z�4���.�X�,�B�.�2X��`N;�(�!OS��C�I�~rM1E���(P�ΞR�~C�	���� ¥:1��)5��+RC�ɋ"�@��4t���#d/~�LC䉡S������.�jPnV�J��C�I�G�PK���Y)
L�D�
��C�ɪ!��tBCN��&���Q�EŐ��#>!�d�Ig�Ui$��>e��`�C��<葘�����(M��bY8�'ZH�<��Vx�s섵V�Xu�QF�<��J�(� ����F.���Z�<�K*[���R�ơ�li)�O�o�<�S��*.tEV�s����G�b�<Y��;�Nh23@��-T�p��g�<�梖8g���F�"�b,�T(�v�<�����A��hY��&.#,�V�Ml�<3L*%����UU� 6�E�<AB��%��d  O�f>1S�C�<	�O�F�q�W�$!h,@5

E�<� ��;F_84�֦���fx`~�<&h�Csz��ժ��C��$P���~�<���Z���ʠ�޴w!>�C7��y�<I�	Z����ˉ-�ܩӁ��p�<q��$CD�j���䅐�$�^��ȓ��<Rꘜ�vq��%�;M��ȓ}U�(�j��8ǡ2x��ąȓ6��D��ջp
t�©	�0ݤͅȓyS�P��ј �����W*Xx��S�? ��R4�T�k�by�g�D����U"O&��2
�q����G�*,r�%a"O�A��A�S�Rm�����"O�l���*xP�fO�Nw�ѸA"OV����C��2�ESTƄ��"O�8C���n�r��e�B�"O:�Z��(r[��s�@�:RY"OҐ�P�Y���0�4��x�"OHC��ŴV�J�([�]�(h�"Of��.�Y�p$��[��h��"OF�x0c�:i�NՊ��	.�"O�[uG!&a����,�Q���I�
�KUK�!$e�~��i	(Q��Õ-��IZ]ʇ�s�<�'�F�W}��U��M���2���6x�j�b�GʏPF�0���I�hG��'�F!�����t,W��Z�)��'�zLÇNZ����V�����4}�Y!�(��n��	x�IQ�J�џtB���49�E�3[�
唡xp`0\O����B8g,0��	# ���J7�K&>V�u�t]�j�bd��Ȯu�����X9-��i��E�c����l�0Jq1O��
��ԱHt���"j�Y_����.��S������ N*|�u���ZW�B�IL"}qC��7����a��:�^U���R4�RH�Ϗ�b��I5�S�"v<�Γg�x���'��I�5.�P�ē^���g��;�@��(M5V2	X�&�1~��q��딮H��H��Wl��'	:�Eҥ$�U"8��ݑ"�y��X��	�EsH��C˄$�4��"(B8w*���!�;i��dQ�>��`��N���&�'�,{�,�;#�QZ����|O�t��F�;R!���[ aF����g�6Im����C�d A�B�X�" ��/��PC�*��y2+zX���R#��0�!��j�P�F�S��x��	�w�<x�FO���s�(P�&o�A�L��L�&��X��(Q�0��a�S53�
q˶�/=��e�g�:U##P5h��܊��@�_<BPCfh40�QGz�l�d�����*k�@ZA���p<Qf��;9��q�)ē _�qd�>�^�`S��	n�j�O@�.�X����4�v��	�zU`���ɕ>O(��C��@����O���ir�7��%�u&N�,=�͚$*�#x|�qΞ \l�УcݗbE��!C�#�^0$�L��C�ɩ'�8I�'�Ģa TP+�o��x�22�7yLPb�BD�'�p�K���&�>E���"`#R\3��W��v�l��aj���, L�`�3�����H@�$ ���{G4�Y
+x�&���SK��HiVDSt*����I<v�"�l�eB8�-QYL���޻s��t�'��sk�6���J�	���}y���3.����9o�Υ��&LG $����u帠a��<)2��K � o(��@�Jr�Իb�[8Gj���欢?Y���Ș��b�<AX���!;u����NL([,
��sD�xV�;�Y�д�%b	?GR����:v��	a���P �d2w ��~�c ��<���*w4AIt�N6n�@0��	:'-�����@8�@��hD y�d�/)p$e�#�6n�X `��;$(���]�g{J̲Z��(�#]7O�1a�/5|O�y3����F��b.&����;���Ǚ> <�z�g����lI38��)a�闒<�Z����܈EŘ,�ClR}r�M=!���w�ՠo0D�����'�Dዦ��2w�X��?T��i��)U<o��9sgN4!	�I �d��eBT��En�DiC�@؅pOؘ�$D]�DY���T6%Q��F��=Y�-J�(A=+�<�q���b"<��5�Сb�����$��K�⓿]� r���)�,�!;f/8ma`*�%,F���(0�]`�g��8�I��'\P�A"�C5Dզt�b�וMU�MɠŅ&n hCtJ�-�nu��e�
VF�1����EՠX��M�H_�Q�]�%�IÕ˟�cJ�(��l�Hj�<�ۓ%\����	���4�6k�}��ҫ9u1�u;�S)&��yѷ�8/��׃��#�8�BR(ۖ~�����Kϸv6�irӨ�~���!>�<E���:��E �����'��
��M8�Ⱊ���w�R4�FA�-�İ[H�7ުݒ�.�
.�����`�I�-ڬ;�� ��@�8m�AA��A5�Q�<�\�M��i3h��J501+����a���6�2��4#A�(3�kܥN��}!s�H3a���0���Ht��,�R�����	0�΅����@�`ݪ��'�]{a�ɾR �DY��55��@��1��;�"�rwu3o�k�q3�㈽U �t)�ѷ1��X�^c�Z̹1��	=����OZ�o*���E:|O�i���M�IW����X=n΀$b�jO-$*�œ��Dj����LH#c���:B"�<x(f7�3yږQ��XL\�g�ŭ5��Ir։�0�ފ<þ����ժd��㟸J��Q�//�S�a׼|�qy1�G+T�]Ӳ"N����GK��To�p��ĸ� ��Z���<z��%�P���Ͱ���`WAK!=D����O��/�@9�e��w� �#dY����9��HS^d�pw�!<F���Xws �R%TZ$�M�*A�)w����*Č9'��� 	f��b�'n�5x1)�,��Pi�aZH� ��'���؂K4��99��T�j�!Pq�M/��HQC�'^N�0�w��� �q:J��"�Z.*s���
�k����&C�5F�z� �Sbj?fP��B 	Ŧ~��c��8%���CF��)�Vd2��O�-9���'7�U��`kb�yq�6A��h���Ii��015kX��O�\uy����f,ZP�
!|Bd�)Of0����f+��	�E����W�$h�f�&�R��G�Ҹ�4a#�)��(��CЯ��o���!�x��s��cr!�ă"	���&:� D#H�}e!�I�X���R�b^ !�()� H� &S!�DUQ�r�YgጰSȼ (��aN�'ά6�'���2�^�Z��Ȟ8*�	��P0@��劁ۀ���C��u�$��S�G�=��=���Ĕi����,ܘv�l��v�,+���Dc�Łf��Tq�C�G<�e�kW�x���!�>O6�����X�w̌1:מ�k�^��	=`m�����T?9%��ؔG�
%��:q���`-��s�<D�`[1^�(O�e��67�I�m7�,(gz#����<�F�~�P��� �lެ��H^j؟�c]m�,XȐ�Ί^X�1�AR ��� �FE�'џdɷD��3N�@)�D�6޴ 	��(�<E�4Q��I�w`����;[���D�_/M!�$6C|$��gJ�=��!�� �� 7!�Ĉ�7{b�hG�K�@��)1���?(!�E�,��1�uMK��mYԡ�23�!��V	#y pCQ��sB�T*� �=�!�ݦH�������N�%�#q�!�G��j6f 3}!�Cg�~�!���+s�ek2��]J0&���`�!��J�\X#��G�h�D����%i�!��	*x���H�2���b� �]�!��O��e:EhA4r�E�`�]�!�!�ē�"�� ̓�~p����S�!�ʣV�(��N7'|y�vF�)D�!���Finp8	�> ��k�&�Nb!�dX�A����CXh���C��!�䞙g���K�~� ]��Y<p�!��>H��6��ax.�cA��*d�!�ղ�>]VoB�jW��YWI��Y�!�$�)P�ұC�Dǯ1A�� h��!��O.cL��Xb�U�8P�4����!���%0I��U����W�
!�d_��)GK�5E1$���Ns!�R�gڰ�r&�"9v(�Tn�-F!�D�M�p����E�e�q�I�G!�V&1��h8v�/Y�*ex'O�c�!��N���e�A2y�E�ȂRlL�ȓoP,J�"A�8���@���DC|��ZS�I�����ܲu��<`���ȓ�(�
� �d��Uң�ׅH��a��t�j$�3�Á.����� dŇȓ=�����b�i��2��
��E���~Yad�� ��Qg�O�ؘp�ȓfI<��̈"�JTyeE�_@B�ȓ�^@I��]2b��i!�o��86<�ȓY����΃<D�� �ײ*�X��ȓp��h�DI�L'��/�).�̇ȓpW���Bd�*q"C�Q->�Z��� Ҩ����[ؙ��G�J��ȓa|�� �)��RmtJ�蔧-�td�ȓ ��`@15����E��0�&��VƢ�dk. `�ar)W�6%�ȓ@� #���B#�e�e#��w�����59�	�6 ��y�t�3p�M^ 0��K�  ��3�d���	����7� ����G��P\��ߏ>�$�ȓ�&8񗂁�`� 1�f��Ԥ��S�? >����ׅ:h���dØ[����"O����BÍ���?�X�JeC:D��x�"� �b�].�R7�;D��02���(��0�? \��ҧ+D�P+��R�%r�i���<X�#m+D��ʧnݱNC�����"R���Fm'D��õ��r�N��tA�>RЄz��6D��2�@K)�̀�S�s���i��5D��ABN$�:�jB(S�DI3D��B��ٷ$!���a%8��0��--D�P�G�ɋp��j!�¥-�����k6D���0آO���$$ �2����A`6D��Z�&/$x-���&�{"�1D�@�傠G�hCU& ,y��#�/2D��G�<F6����NU4���>D��ZeA�%��u���c,%���>D�X voNI���^�;B�ۀ.&D��@��u�Pt�!���e�&D�4��c�~K�q�R���L"�|�R!%D�4�0�	A�R�2a�Q�~U�<!��7D� sg`I�@��NP�X����D5D����h��S���� ��EN?D��P�#(L�H�MK�_;:1(D�ؚVGi���6/<�8��)D��3$͇�.�M3��%Id���e!D��2LΝm� �0K�- B�!D��k�h���l8hq�+I�Q:1�=D�T9�͏�{S0�aP#:F����@-D�x!�/�)5r$��b�R-t6��ҥ�+D�8�g�70��PY��!D����C�%D���թ��W���c+`,���`� D�P/�%UH��Ƀ�2��4�u�+D��� R�{nJ9!D�@�T�[��%T�TK��м,y��0DO���4��"O&��3�ʛ�|���}��[�"O�;����l���6k��%�Hb�"Ol��Ue�:.�楛��"&/��`"O��hRg�!�3�C�
P�:"O�L�6UM���"\��"ON�i7#�-� ����ߊ2����"Oy�X�)�v�-wŪuH���hV!�$FL�TaN�	�l�R�
�c'!�d^	���q�Q�u����P��k!�S9_���ũA�ܐBt����C�Ɉ~�����Nk�<�/��p!�C��j����`��g�l,���� 9�C䉍x��P�v.zAj@��C�I��dL��W�t�L ��F��E��D�<Qs�ݳ7� m$T�Ï�m!��ʄM��� @�3�v��΂?RF!��#TW\�ڒ�  Q�m����uO!��%�H�YUkӜ��<2GmY�!���.P��yp�'	��駬�q!��4�d��4K�p�pD��!�S�v�l�)�� (��a�
(�!�Ě���&)Ѯvx�)�*�#�!��zw�)�n�	Q@N0h��N�A�!�d���@��t�T�$����:�Py��^�wɾM�#�(��ئ�+�yb�Э��&���{�~��v�X��yr�NTpjr�� b�Ĩ�j߄�y2'GH��u� � w6��Δ��y2��.��1{�m\�Ubl�q�$���y2�ɦ�ư�Bϔ�K)�������y
� %��?� �!j��2�0��"O�E���V�7�L�h"f۝	���"O�=aT.-,R�{�Z7�%S�"O
�Q+X0=��m��~)R��"O�ّO������TlO�qH�P"O*#&F�=[�P1�J<l��p"OvJ$���@k���/J)(���k0"O$�P�,ڷL�X�IS��=��e�!"O&�*w%A}
���){�|j�"O�y��O/@����k��x�X��"Or\�NʖGr���̗FT@u�"O��1��܆rd����<(�Љ�"ONpk�LzmC	��
�<Id"O�}i�($20�h{F+LT��"O��6�Ď�qDF[��d�C�"OV�i�&]'rp��`&�&ӄ 
D"O�)��)ʥ)Ȕ�p�
�v�,��4"O��ǀ��z��*��E�N�����"Oޅ�)�W�h�D��y�တ"O���-'����IR T�f���"O�T�5&$$:�tz�b*�@��&"O������l&���0�۳j�y�&"O��ư1��m��Q�U;�13�+7D��9�΃Ow61��$�D�cw�2D���Ô)\���&N��!CA�7D�H ���F����WZ)��>D�lQ *@�"y�q	��HW ��%+D�� tA[�/� U�P��$��`d2D���lU�r
p��tj�1�j�B��/D�L
�A�=D�����F2#60m��M8D���ȉY?���DY-R���C9D��1E��5"b�U!D+7�B��;D�pC���>S ���q�D|��@9D������j<��(��9��|)P;D���'���2�z!�-��.��e�ǩ$D�$�#�x�@HTJS�lݘ02�#D�X����3$^,	� P�:�Z`j D�pzv��:F4��y6��4�H�Ӏ?D��
��/NKqэ��!�z$s�i7D��*�#V*fֈ��$V�(�$|�T�3D�0!�%΍���Hp*�-(	"��%"D��y�ȶk�Pu�ê��!��Ѹd` D�,0���$�偆��=A `�1�"D�����B,1����V)��A����O2D�t�����q��a�r�-���2D�uF̥}��a[�g�d�x��,D���ү�
�N �QD[`��Ma�l+D�d�5�8�Pm� ș/;;��K�+'D�<��K��c������=/� �f$D��YA��w��] Ňܨݺ��$D��� �P P�`�d�Vfҙ���7D�pS�)�8l����3b|A��'D��ʁ��7j�x���^Έ�r�/$D�� ��Ν!��@�cΝ]�.���F"D�T���Sazh��Ӎu�R<2�"D��9�M�7+ :B�"`��0�I-D���B�4�A��(\��h��H4D�[���Uf���PA��%|`z��>D���aC^�6����}W�(0��3D�$iD"�C"d:!&��"�h8 $D��'I'$쁵jL�ol�P��#D�`3��1:H�+a�L#of*(J��=D�ī`O΂42�x����L�Ԉrtf8D��B2d �9b`�G�O�n�@�9D�� xrEDN�V����WT���"Of��4I��L ��A�D�+i[p\	�"O����U�bUr��ccʉS�~ �U"Of�X�C�^��	���W��D�@"O� h��I���w��%S���a�"OL �	�����	$Ԗ\9 "O�ѫ7'V�!�� h�={*�U"O8��k�O�8d�r�^,U"Xyf"O��������tJc�G�-M�D�W"Oxz�8d��8 dQ*a�:���"OX�a��z5�̪���0��YQ�"Oj�[ˑ�p�0-Ya	ז:��xF"O��HN?F��1��4k4�8%"O�TcIP�@�!At�Uv4��"O��a���8R�6�A�Qo�B�"O�i4�M<K�#��\(L��"OB�فNɬJ��]��F�@�Y"O��b�ʙ�]/\V'��c�H��7"O.��
�6M*3'���G�>�"O��T$`����/ܟg�f�j�"O�� 5IR-��=	��s2��U"OX��n�
}�Xzp��-W'�[�"OD���Jټ^W@	���p,b�#�"O*tGK�;x��q�QAʒ��0"O$Xk1զw"�QyQ (n�` $"O��g
)|8�Ea��B��a��"Oz!9A��0(�e���R�n�x`��"O��&g���x���A�R�@]�p"O�,	�,X?QrV��e�#u�,�2"O^=#����e^:�'E��"O��)�H�h�Jѥ�@�p�p��"Oꘁ���\�n�xri�	��Y�D"O��(rv��,`���-�d���"O�(�.�D��q��xB�8��"O���5%ע_���Q�&@1GЈ�"O��A��S�,`ٔ�ӷ�8�Zt"O�4���ʤxj�E�c��T�g"O(�_O�d�QF␒CU�w"O�rϒ����j�L�R56�3B"OT1xS��=1I6�`��Р;DN�"O���k	T����nKC�x!a"O��S���{���l�����"Oq��=pl��Ie.;G&��"OE8t�þu��xBG�(f�H���"O\aP�Y��ԅ��� A�*h�"OD��#R:xi���w�)8��(jT"O�,Z�J�+NS���&o��l�☓1"O`)a'��QY����Gs���"O2̀P��1XƬ��\�(C~�ZQ"O0�����8[�<����ɑ�"O��K*Z�}�x���A3X�j��Q"O>��DƘ��=�`���P��"O�Q��/+!*�@W'�"o^�K�"O�P8VA�J�2)� k��L,[e"O��1G�˻a$^�rE�R��T��"Oȁ��ԪI��$	�DI#m||#�"O���M�?b%|��pIQ�C4��D"Or�st�?K�JiH�ꐇjS��;E"O���ЪaxL(E�O�c���Y"Ol�1`HU�V���+�/|{�T"O�I���-(2�0���?m����"O2���MJ9=�����!\//"&�3"OP��$�:�y��P'Z��r5"O��;C@F�ȄÆHՈ���[�"O� :���i�*Z��h��H'zΖ�k�*O�ᚵJ�n�T� ��N�e0XH��'j�b�VJn�tA�LY�@y�'B�²␑#��	�EQ��$�	�'�Z�s�E��_����4���d`	�'��]r����5��igƖ�hb����'�f�c�¯@l���)ɛ2�
ap�'�-z�c��씡�L}��uY�'b��A�cfbaCF��t��m��'u�U���C�z��dC�	إn����'��KdƝ�(�R2�W$1�8�
�'&��p�	�4zbHT0�$�y
�' JhC�,X|�����D,r
��-Pb`M9L�*�kRm�h����'$�a�We��c|�H��G�D]��'���u�S,8YZD[��4zݦ-��'o2�0 
@�
X����i=z���'�2{��̸7�� �#�k����'�r9�qN�`JR��l��%��'#z虳��xȄ��	)~ĠJ�'�x��
Z���A�"W*��5	�'-�Єm�='� ��IC���r�'!&�!���>l=N�BG�@�,n����'#��A��22Jl�SCO!*��	�'�D�S�E	t���� U< �Y8�'����G�!fI��\k-.h��'�M�1&[�F��PJ���'Q�	����?�ڤ�fF�:�'��[���B%B�;V�+P�J<c�'Ѡa[�j��Y�PL���	W��I@�'�^�
0*�#`|�a[���B��'����G�5V��(h�S�6~��k�'^���Qܗ5�ܸ�7@N�1B�H��'���CF,��E`��J�?6�d�
�'��1�JƍK4;Y�Y�3��+aN�C�I�	�6�Y�C>�ĥ9R���zM�C�I�6�`��\�ƽDF՛��C�I�n�:���S�ЍH"���C�	�}�(���W��N�h��Xi�`C��
'dN@�w�D�BR�`E�xLC�I�n���@6��z �g���B䉃YT����1�����ĭQh�C�I+v�� 7-ח*��J��ϔB��C䉗,��LrEoC1J�\ڄ�M�n��B�I���`p�ح6��="`
�h	rB�	�q��t��k��]���6i�15�xB�ɝ=P���Ɇ�u, ɀ5c��&�C�I+;v\�1�Y��cV�
�M�(B��2�`�N9.-�5����7�
B�	�kW��	��Ю1֤m��(�
n�
B��?I�.h2J� ��96Ɠ��C�I(K��)��#�f�:bT�S�C�J">q�Iܻ}`�x&��$E��A҇��<ѐϜ�� �≂77����"�Eʟ#aKr�S�O�|�q$Gֲm������|�
�J@엙��	�g�":�0���R���^�F���f	=U�4�����$z�`xa�ml��oC��H�(�W>�Ǧԭx��8ʥ�@�[�6)kaG��?�'k�#\�0�O�2wf��D38)�q��Q�u����5��9�J0���[�[�qSG�8\����)��k���;��M�@��ct��$y��D�V��>CZ�p$���F�b�t�O���2������ѧ~^C1lPj��"�M�,y���A���m�|n:�'Yu8��7�ϱ!M�|�bE���(�E��/zb��D��+V6�����rܧ�ħ�2P3f�6p�����`(:�bC�S`Tyi����<D	��Sk>A�4�Y�Ox4K����"��W4I���g�1_� 0;q_r��I�.z.�pR� E8'�`@���
�&��L�UR�{B,F�Iڌ��p�Q��C�/[�����-Di����_c=����*�9�@�l�<���Cr�π 8�b_�g32}A��٫F��)�ԫ�F���s�4/��=s�(�E�xc?1���݁|#���t��lv�!FMȔ��'���S��P�SܧJ�zH�FD�"�ȸB�������ȓK�"pSc="3�@��GF�
�.d�ȓ�Z�#��>�4mc�.,y��M�ȓw^�yP�Y�:�^����
./���ȓ?�usv�I�V^���U�; 8ćȓ=ΨɃd��lS��bH�j�� �ȓ\1`T1���H��1�X�~fU�ȓg�r-�,H¾� ��=qu^��ȓISn�x�b�6�"�"
\76���ȓ4�|�r?b�C҃��f.�)�ȓC����q�01���%o�����fF�e[bI�	|���qS�G���ȓ?��"RꊂSV
Yd% m&Y�ȓ|�He���L�y�t�aC�\�fr�E����A��9g]��2d��|�v��ȓ	�8�[��+2��_�ʆ��}�<���[�"�����E=@͢E��w�<� ^�L@u���7p��ۗni�<��I�Dy�dFF#F�q��`�<��Ǉ�K���݋���Gʑd�<�p(܃M����Q�^,''����`X�<9��Z�C�.���Ć(U
���e��W�<%-T\��5�` X=wO��SE�KH�<��ʉ0qP,Ðe�${ �C�<1@-^�9��� d%m�
�hpJ�{�<y��ʾ�R�"�HQ,>e��'��N�<9���
P3�P��[2xuhD��'�a�<d��m���J&��n&p��pF�]�<1$�

 ������0��ǭ�W�<�B�_6��-�4m֊g��i�I�m�<1#a�EQT�S2�"p�%�C �u�<��f�n�\=��'�;H0J1Bw�<a�,L�#'��9�O]-,���¡�r�<i���	�>ш�-۫aA,�)�u�<)GްV�����!8�Bp	v`II�<��O5$�p�;�AP&;���g C�<Ѡ蒿 *�z�-WC�ʵP�"D}�<yBgD�J}��q$
.37�@�Iz�<A@�� c[����L&`�:�X�RA�<a�儋q�4��siڤP�����|�<� .�?���;1J��s�*-ڡoo�<�Ʒg���镁}��92���l�<�B�?~t��3Ť;�f��S��n�<� ���HƦ1AHY�tKL��#,Iq�<iD��FK�Ɉ�e�4[�8���
n�<Ѵd/`���(L0U���4�~�<��O&g��B�h��@�X��a�<)��޺D� ])שV6���0� I�<�AI��2]���Y� v�U un�F�<Q3MYg:Dy�ͪj��礔D�<�L��`����N�B�;pf�D�<qel��'��q�@
�y�����i�<��� d�]9$Gbp�A���b�<)�@��X�ˁ��]*;�a�<� �]�M��Fd@�����HZ�<Y��K:qd�����r y2Q�C[�<���$�I�U*�����eM~�<�b��*L��	�Bީ9$�U�<]<�S$%���(� �Q[�lԄ�f���g�M�j�B�BP��ȓ���T�fI�x��<��l�ȓDV��[q�)b�j0A���H4����S�? ���y��lBVEC!JWl0�e"OP<�,�������[ܴ�{"OV�B� א��������q�"OF1ᵧ�"�Y����5�t�0"OZ��U��=��b��T�F�1��"O��)���/�l����]��X�ᑑ|�'���)Ro̝+U��(�ǱA��ً�'����%�b	0�iň 9E�yr�'<R��֩ܡEJ��#$�.��s�'(�pJ���e~��s� �}����'��9�CտL���9c�\2ga�й�'�6u:�Yl���:��?Pbj�'|T={&��:E��9y���[!.�B�'�vMӳ�S�jB(t�V�O�<���'9��XWŒ����J��M(�q
�'�e���(t\	+0���,)�yhX�m8����/	�X��$�y��!Z��x�d�-�0w���y�M])M��p(T���w���J#��yBIB�|���z¨U;]�����ŧ�yR��u�8��qI*V4���&*���y�L�j"ps!��U�(�Z%�&�y2E�
&z42�M�~�,uÔ(���Py"D��1�$��Ƈ� ؾ�A��]�<����O�jx�6<p(�A��~�<1$e��,��p`R/6SY�D�{�<Q' R '@�A�A�	<6t�kBn�<i�
B�__����q�R��3�n�<���7'q�q	�e�V ����T�<Y`'�~ 2������0��v�<�Jͺ��3M
�"�\q�<	O�;
I6}�,AgީI$!k�<��c�V����-Z�RiW�N`�<iT��lmHQ�@�]�)�T� EIZ�<	懟���j�h�)D$[Q�W�<�d��%,����%K����#�N�<�DN$d�4�aT]3r���O�I�<�uƖ!�@���1�><�q��j�<Yr�H
U���C��,\i#lUi�<�!M�u_��CS����z}����g�<�a���(\�'�K�]?ހ���Tf�<a�R�h�`I�Iܴ+;�X���C�	�@���C-\?��#T�W�XB䉓l�0iX����a��'�C�I����M���C��ƀx��B䉄%�,�Ar���b���a6�B�I���eIO�d��!f��2�pC�	�W�y0�/�4vɔ$G�
��B�IjBI��CD�8�x��a	�g�pB�	,.�6[C)F1q�R�P!�ІA`B�IF�(���3V�h�k6�ΎCJNB�I�v򉻧��$�>�#��ѫ[)�B��Bs�q�d�ņf��a�R�`�B�I 
n��W/?+�
�C �DC�	�4V�3�Q�b�`��F�e�~C��b�LLӗ�8}��T1T�׽qRlC�>]�ʤ��#S-�\�O�/7.C�ɯ-Ҥq村wӠJ���5%\�B�	�	�Q�h��gh�GfL��B�	��1H%L�,,8h���	�T9�C�vO�Hj!*�?'p�S��-n@C�	>W|,aPI	�Q/��H)��B䉴n�l�z n�깢c�����B�I4a���f�-65�11��^��JB�)� l�Ip�в3�T8 a���u����"O���c"L*P��h�ǰ{�R�r#"O�S�X�B����퉎	�vu��"O^D2#� T��e�#�,��"O\pk�
 )6�PA���<P�7"O
黢"��3��qd�N�����"O tx�F��G��R�Z�9b����"OnU�j��~̀m�-��"a��÷"O�	���`jZ�D�բN8���"OdЕ�Ɋ[^�����D�q�8�!"O�<�e.	�c�Th�7#�8�j�څ"O���f�**��1�O�`\kc"O��F-E��z�(M8H�N)4"O�)��"��	jYC�����R�"O��� 
jHUy4�ߪ
��1�"O ��ۉ9�b�駂�"?���c�"O �+���
�N�86��z9;�"O�A/��ll�Ryɢ�3�"O8�:����`��l�#�N̂�"O�8�����#{���IM� ���r`"O�����[ߤ@���ʥ}V���1"O��qg�� �� �͐+�p"O��M�}8L0�U�!Q�P`�"O�(��=_�����ޟV�*,;�"Oj�HQ�/lL�e�to�[�X�"OH��х߈h�� )�-�$8���۱"O���D�/���p듰u��\��"O���!�9o�\��$Љh���6"O��h3BA�Ko��1 i��XI����"OV����*Y]uS�B�2n��}�"O.�	V��"~���PEdEX�u"O�4��m�&56$X��A�m:���"OQ@G���Qx�����z���+�"O�8x�h��V�tZ��NP�X1a"O�Z�+�&*���l���Ѧ"O�x�AE�'	�r�0E��+#��UY�"OF�vC��u��Q1�J��j�;�"O^i���M�5��� 'ޕ%����"O�K�`�&�Ah$E�,Ằ�$"OD�Q�^^
�����%Ý��y�ʙ�G�4d�%IƉZt�E�U#���yb�İm�Ј��MI�P4�@�ّ�y���?1���K T�28�d�B�ybc��}e&\S�ĉ�D@�P�@��y҉�^@�!p���:_2Ԋ�B	�y"/�����9���6^���dR��y"��*��-(�ᘄ&̼J��U��yb��t��� 7�mZ���=�y��X�l���3�X�&@x��`�0�y��W6W|L��3%��	l	%����y�����,P`P��9st^�y�I��n�&=k�*�1{�nB���yr �:N�z�3���m�XQ�.�2�yBe�7.�Lq{W(�h�ȠXv�ތ�yR��`p} �L ^��ԑT���ycT+!z��-5~�s1L�-�y2���I��Y��ڜ"̜h�*���y�/A:7�x�C��]�.�h��D�ܺ�yR蔶G��x���Ř7�I� ��y�H �[�]`!�`�|�t(K��y���18��'f�QGdm��BI��y��1f�\�@VǍ�qO(y��`@��yB��nBLTʦ�P�W�P�� L*�y�K�hB�p�b��T�,�b�B���y
� ��)�b�h���2	2m�N�a"O8dq壐�aV��	�V�ꩋ�"Ou�0)���%񖫅%-����"O�%��Dͯy�l�3�J�
��<�y"��4`B�
��K0a(  po���y�GәOU�=K3�K�Wilʶ���ym��M�$akq�B-D14x�����y�"��1}��ar-�<x��:E���yK�Dx�u�R�^�;u8F���y��f.����Ƨ$�0�!��J��y�� B�@�$�D�"�b�$�ׇ�y�*�-N�Y�c	���Bڀ�y��Y���(PnSF&�*�&ځ�y�-�O߀I�0#��>s�X	`��y�k�2��l� ��:������y��]�ˎ ��S�4eʕ�E�P��y�D�q�0�4E:*ex�� ΁��y¨R+H P  ��   �  �  S  �  A+  �6  %A  �H  �T  ^  `d  �j  q  Mw  �}  Ӄ  �  X�  ��  ߜ  "�  f�  ��  �  .�  u�  �  ��  5�  ��  �  x�  ��  ��  � �
 7 { �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,��	⦽�'M��F+�~Q�HӘ8ި�I>��'lOJ5c�D��9=�L¤U@Q�l��"O6p:��˰1@�Q�Sc�W�4Qj�"Orr��̜+��Q�"�[���Q࢓|b�)�S�G��] 2LX o@��Ľ`C��b#�x+�m�:9��2G1P�.B�I!�f��Tl_�.պ��VA:Y�B�	7~���"�3'jes��]$	�|p�
�'�b52B�O�`��ub¬�4Z~�`�
�'� ģB �0��2���W�&|Q
�'?��q�O�p��)rF�ٴ`Dm"
�'������!��
���m�(]��'��a+�I��
$ǈ�M�p��{�)���`�`���	�u[xI�3i.(�!��/l�(I����Ed��#	���!�S jT��M*f]�<q��R�o�!�䟑k�v`���*M*����ïG�!�D�'o�{����n1�͹ыL,DZ!��,:�@��p�	@T��� R�!�ԏ?�q�G�9	� yQEō2.�!�d�. }6I醇S:k�*��Ev�!�$W'K�=��YڨY $�H
�!�7c��5z�@G� �>��s�Hln!��� jԡHaEI	�P!��A�$i!��:2_��`fQ�� �Z�-�5�a{��D�?-Ix��s�V���{��P!%�!�Č'`:*��)��t�
�bp-�\n!�5�M�"Ƅw՚�;d�OLn!�� ��J�DC*�0�&M�'^j��D"OP-��;)�
is��!�VqT"O<z�K�N�8��"��2���"OR8*%��,��m��E,v���c"O@XY�N��SH$��[Gx$u�"O��y5B�$Y�䭓��q�ir0"O��3�	<\
L�z��Chv�!"O^i���@�d��FW[��""On�CvF\��fiܸ5X����Id�OzT+ A���k�5n1��'����Rg�H����	x��D��葬�y�.̧F��A���,q{��J���y�"ԗ,������կ4���p +���y�#�n�Y�q�N�(�"�����ymP�^?�� dDJ%g���#�I�y��F��:U�eԯ쾱��d�0�y�ʞ�#��J	���ݻ�dY��yB
A /Ѷᢓ)��
��E��p?q�O4�׀I�c��X�bl�9Bj��"O���'#Ct���n�'�A�ט|��'�6�:�.�P���ޥ�J��'Y�œT��S�d��өލ	�^l��'d�A��MG�Ks$R�|ʈJ���a��0f&�"���fN�<�����?	��3S�̹�3'Ε'F���ҥ�e��LxR"3}���!c����%4��4kլ	��y"�F�P�$`CF1�eb�-���'�ў�Ow�C�T�=�x���Y�b�y��'v���P�آ&���۳LF���'�ў"~jP-ޅ B<���NfSzI𢄗Y�<I��dݪ�s��,���#�U�<i�'��|B(Z&8�̈8�HJ�>OV�(��Z�?��'6ў�?�y0iU�|y~�	Kh����G/D��6l��;R���%L5Ki�%@t� D��:�lZ/@T�$P�^�X��H�! ��}���S����˗��@i�M(�N%.@�C�I�+bn��Њ�l0�]S�/��W��C��Q���ūĐ=:���5�"�p듍p?I�F�'��횧�ӯ�򭢶k?i�O*�z��
������P�:�2��J�'��u�P�S�dR�a���?��|`
�'�qYuE[�A(3��'%�+���,�S�)��fP�S����thx���:F���>�3�ΟR�qQ�Ĉw�lsS��"9!qOr6̀b�g��HRm(T3v)4z�����R'd!���#IԀ�@V��9[b��DkK|�!��TPҀA��xP��*L-k�!�E�Ѳ�a�D?�$�H��X�!�$)k������b��1�R��=�!�^�\ ��Q�O�+��� ۮl���V?)�aP~�j��ì/@I�J��|��	`eb��z��1!`�H�N��I%FK�C�t��t"O�,zī�g���+��'P�>��Gj8�(Dx͑�6Z	����7i	"1����y���|O��� iĞx�Xu������y�E�y행(�V/K*=��D�(O��=�Ob5��D@ ;��EB���AU��
�'��T�t�3k�b���H�'L�P���!��qji*uY�"�f���ώ�	C��ȓ[�Lち�9K��j������[�Q�<F��e╢G�o����v@ 
s0��>��jY6(�%Wʔ̙�	"�y�����`�?�ɤFۤY�����
βp9����̇ȓ�<tsǭ�l��E�c�mA�,o�v(<� P��G�8\�a�T�)f3���4�I}�O�J�3�(�:U��� X��'� d�U�W-[)��pA�ä=g��Q��"�G?�����d��c6����X/KA2�T�'4�Ĕ�>n�r�ڏ/]�d� Ίm�^c�(�	�ei��ϯ}�8�H��K�0���?���-�)��](���ĹyI� bUg�&HC�	3G5rF�+t*b�17��7M<�ӺCR��'�ڡ��*��B$$W8aC�@�'���ď2@<�����`��]!�'n�s�m�$r$��Vˌ�F\A��'Ȳ(#��ߓYp:�
&f� <i�p��D/�F9\��v��z|u�^���=��{rᓨc��T T�I�>�B����#
bB�	 A���ѮG
)�^�Rv�Ϻ���~�i�y��I�v<V�ⓣF4bq���+A��C�	,L�m�GX��,y�Bb�5~�7�c�,�V�'�6k�KX#�2� �F�#��u��'�b�{��'�rq�4n��I�Oi��(�)O��r��ת3���zp6Odb��x0<O$�}�'�^�er��G�x�Z85C�_�<aU���8�$��b�LSW��[~r�x��?���K�B�(AV%Ɲ�49�g*D��ñJ�V휜��N�Y��'%D����Y��0��םL)�]�ы!D��AG�}�vh!�
בUt~����"D��cԅ\1G��=��Gm>��Qe"D�T�%d����J�l	h�V��E4D���Ci�%���dd�%d�$l��N0<O�#<&��!*�t!�D�J8	q<��)U^�<��-˼>^Ĩ��)p<�P�X�<i!_��\�Dc6mY�����H�<9F��=+�Z���@7@*��ɐG�<����u��ؒfOM�y����F 
A�<�-O.^��0�4r�4��&�[@�<�%IQ�a�]y#��M�$`Z���z�<�s�^	\�Q�/c� d�s�Jx�<�1�^�!�b����$�f!��+�v�<�W*7Ou��+�Mi"�P�hr�<�B�� tP�%ʦB��pE�ɻ�yB��_��K�H ��ur�g�9�y�mV5k@��N(	�hx�B��y"FV�wt �Eo��hБ	/�y��$�%w˟)
���Q�L#�y���&l�xQBݎ'��0��ֲ�yB*ݵh���ª�%x:X�:� ��y¥ŵ+o���u	�u��Ұ���y��O�B84SW�кs�&U�'B��y���;h�vP�B#_�ra�	�Vk^��yR��.3U���żk���eL���yR��-ZG���L��]!�P����y��R;oȈ��	�M���0JS��Py2ƿcG�s`��*�B���p�<9 ��9H�n��F��� E��"�i�<�3�3P��hk#�L$�,8c��CA�<�`M�<���I� \��1�c���<1���cÂmʢ�΁G� qA��Vp�<)���=	�Q��f�Ć�F�<ѣ�"���f��fXPP��\�<a��]�](��6J��XU�8���}�<Y��S�}) ���l�
R���kLw�<!�'R�Wf���f[�5���s�<�T�Ϭ0�~��	�+_��p��n�<��p�Ȩأ�
!?��|;��p�<� �׎'mR@k��U�,d)�"O ���+̇��P�"Y� 4A�"O@��@h�%�n/�y�V"O�=zt�ؔ7Uy�퓿Z����"O��à��:�A����u2��E�'r�'���'$�Q>��Iן8�I�{{�4���^��6`W�~�\������ޟt�Iݟ�	ߟ��Iҟ��	9���q뜴c!�A� II�{�	��՟��	ȟH��ޟ��������şP�I�=l�!r�	Q��	�k~;�L��ߟ����D��ϟ ��˟d��ǟ ��ux�=i7�']�,��ED� ���	۟��柬��ԟ��IɟX�	ǟH��KX(� ��F[�Vqɂ��P����ϟP�IП�IΟx��Ɵ���П\�ɍ.gN���i�<x��d��[>�%�Iß<��ȟ���ß �	���ޟ�� s�.��V�� $�KaXܥ��ܟ���ğ���˟�����|��ڟ��I1R�.�y)�gi&�C�M�8���,��ߟ���ҟ�������� �qaK8� �`V7Z5>��e��͟��	���	؟���ݟL����Iϟ�ÏV+�`쨐`�4P��"4�ϟH������I�����4�I�����͟p�4�K�<ȣ�0��\�D��͟��ğ<���������d����t�Iϟ0��5���	v��b'�Pџ��I�|�I��I؟x�ɦ�Mc��?1u�ƾ\�7/<3��I�>����Ȕ�����¦���[/R�j��1��xboZ~���6�4���b��i�a�!��i)
K�l�%"�Ʀ��	�{�N�m�`~R搶^����%HM�i�,�ڠ"ĆH08�<؁w�#91O>�$�<a�����2�ؽ���5���sH�!.�o�7��b���b��y�m�V�u���F�)!~��l���D��xӚ�IOyJ~"�ˁ��M��' 2����P@����7*�1x�'
�:�E s�f����i>��	�F�Ё*F
E����gI����IhyR�|ioӒP ���J��dT��/# �M��[�?̮�82)O���qӐ�	I}2��'���3d];^hX��;��˺�� �ċ�o�1�4��Ak�)�/w=�!G�
�����%�R�-�*O(��?E��'8�kbA� ��)udʤ(�B�ۘ'&h7-���ɖ�M;��O������@�Od�����i�Lr�'R�iO��囖��P�Æ'��@��(�8S������N��e��X�V�'����Ϙ'~t��ڦN�V�Y4������O�Unڐ�"��	ߟ���v�'C�z��VK�Z��b�:�h��F[�T��4�f�|��$!�i�HP�D�+���0�/)x���n��8�L�cMߺ�V�|Q��j�P�+���tğ��WK*�O��l!p[�����ztxr�k�(T��E�"o�PBd�	��MC�"ɩ>�`�i�@7�O0m�F�y���w䔧g\bSC�B1o7<7m2?	1L�x�Ő�!ش��'LeTaГ�H�=C5��p7�5ꡢ�3Ŷ��1��6B?Ș�6`��(�)��4��#�=H+��I��X�
����i@�T�� @Q$ļ4�M��Ē�d��I���'k&�
�� �4h�qӏV��X"c &R0\�"́3�hM	ȅ?>�c�ň4�D�C�ԁJ��,�a
2
�<)���+��a ��/�,M�B��.w�����M$LB�L�T|�	3���d����!�|�5@�/"�Y2F�>2Ƣ	�`W�
	LH�t�/r-���'��'��L�u\� �	ş���y?�F0x9b, "�n
���G�.���iI>����?����H9����Dn>)(roU�ܲ�@��iBR��>f�I˟�	ɟ%���3m�dE�׆g�mr�F� |������<����?q����dU�+����0�2&�J]��Q5u	���Qk�<��?I�����?A�~��e��#'�%P�'� Qꦄ��䓿?!��?�)O� ɻ?��쓀���kB�A&��ѷ�eӖ�$�O��>��O��$�0���u� b咖��A�S�z�`��?���?�-O�1���|���Uj}��΋�wy\U�ፍ�R>X�@B�i��|��'�b��j5qOD��$�>;�@���V5-X|�źiB�'s�	�;F�ДOw��'�ta��O���U�ʣ3��7'$� O�D�OK�0��~�Ck�(�$$[Wl�z���d���'_fDJ��'���'2�O��i��#�V�"�X��]-yB!���aӦ���O��ð�(�)�Ӫ4E�)��fķP4��1e�N>)�6-wpj���Od���O��ɢ<���?�3néi�ry�����+�ƽ���8n>�&�ӡx�O>��I�~������h�D�TH̋Iv��p�4�?q��?�DB��d�O�D�Oh�	}.�If��`uFӶ��äc��
�Np�Iџ��	���0@O�'Ѯ!�G /C0��[�h��M��R-��,ON���OJ��7���`�(DM�Q��P�Wȋ�8�+\��R� M��ĕ'���'�W��x�πL�	�a�)=d!y�J�:BE�'���'k�|��'j�d [�$)�`��Cx
�G�GU�PƟ|�'��'�	�&Y���V��e�٢GgD)��fƮ*An��$��ȟL$� ��ȟ��w��a?����A�qv�?8!h�
R(�b}��'R2�' �ɸ���O|*�� (�c�'{K���d�g�pp)��imB�'��	ɟ��O�R�~�`�E��bMReeK��v�{�KϦ��I�h�'2���S�8���O<�������?���x�
��I�'�i��ß4�������A�s��ث���+���W�i���VHd��?��W=�?����?���J(O�ӄV���kҮ#: �
D�!���'��	/��#<%>�[G�3Y:<�g�\9#����c�p�Se��O����OP�����S�T߃yN�ř��ɰW���o�&q�f��x(Gx��IN3~�Ykk_�QA���D�W�A���l���ӟ@r��yʟ��'4�`&�4xn	�5��O�mX��!�r��OC��'�"�M5Ԯ���
0z!�-��6��Oz4 C�b�i>��	�l�'ծu� �^-=�� ���M�H��41�+k�b˓�?y.O���O���?�"n�#�%a�jW�a2�:GfU<V�,j(O����Or⟔�	N?!6c�?璽��偀:	�����˦�;#?a��?����Dԇ;�ް�'?�`���f��k�֩��J_$A��'���'��W����j�$�'H���#TX��(V�ٺ!�#��>���?����Ƅ"��0'>�@�Ϧ[,^X�&�S�
�̠�S	 6�M���?�/O��d�|�����<k߾�+eŖ?=>����Js�L7��O���<�����\�O����5�M� 79D��Df��=W昨�뒓�M,O����O����O������$)���>5�Z�E߻HB��q0�i��	���9	�4&#��۟���)��D���d��M:`H|���c1���'�"�'��#�9O��禕����L��
ݱ�����c&�M;HK81�V�'"��'K��I&�4�d d�qz���Y%�NL� �����ğ���ɟ �'<�s�,�	v���+�jȞ[��y�#C%Md�Qߴ�?���?�5��U鉧���'�"�ԁ�J=��O�~��v$X}��7��O��į<��\?�O��O �QNOY"Ht�q�9	8��i?���,?�I����+��
p���1d��X��U"B�z	­�L<�D�{��?�,O��$�]/rU�@$P<mu��س-J�5������<I��?ь��'��dļ@(�!�ש�;f�xv��nH��������O���O�˓Q�R���4�. 13�����(a�U�	���]�x�	ٟD�IHy��'e�ß,���T����R�t��a@d���ē�?�����*M�Ҩ'>HՈH
�u��
�km�i��H��M����?	-O����|b����S*N~�e2fCϖa�Ip��7|=r6m�O���<��&K�OM���56ɗ��щ��F,c$�Q&�_��M{.O`���OV��O����Ƃ�Sb�
�*��� KQ�r�3R�P�I?R���	Ο@�'Q�TZ��]J�س@"��P$JUu���J6�OJ�h�DxJ|"�@Q4(�-���%\�,��P/ۦ�CDC�	�M���?����z��x��5��D4N�����1Hb!���M���?a���?)*O��<���t�`��PdEbź�����X�3Ѵi��'��[rޜ6M�Ol���O����O�NY>BĪhp�w��h����<N�f�'�剛t�t�)����?��B�J� â�*�4E�f ��ɠ��P�il��ҿJ-
6��O����Or��GA�4�OXՋTć*l��;$�I�A�,1�R�daBw���ٟ���ȟ���a��g��p������E��2��Z���)�Gm�"�d�O4���OШ�OL������a��e8\({Ԥ����$c�"�/}���?����?9����%���oZ�e�L j��0l�� �&�RH�ܴ�?I��?a���?Q,O��D�83�iQ3J�HT�&3�E(�o�#^�XmZɟ@��㟔�	�����"7|Hl�ҟ�	�j`y�a�#�8`0�2@)exڴ�?����?�)O|�d�X}���O6���.0⌚�Ǝ9�@$8D��g!���O��$�OR��G�42�n�ݟ��I���S�Qz��VF� �X��� S�&nfm��4�?�/O���ҖU��i�Op��|n�Z�L���N�5��9����=B�B6m�O~�$M�u�m�L��͟��S�?��I�;q��S��rl��W�ݧ�&�ШO\�$H�J�<�$�O���|�L?ɺw�O��vQz@)O�S7�%eKcӄ��������ϟ����?Y���$��퟼���?�Dad71?l�Q����M��ҫ�?����4�2��"����j.,\a�d��V��r���w��plZϟ���ӟ ¦(Y��M����?9���?��Ӻk���$���ƣO�R��F��0��<y���?!�6�ƽ�w�H ��Iܩ"9\@��i�B
ј[�$7��O<���O��d�d��O�s���,��c/j�#\��"�cc��'���'2�'b" ��ܹ0��?]���G�	��}Ӗ�D�O����O��O���۟�{W��0R E�E�;2w�D���[��ğ��	ڟ����L�I���B�d���M#@���q�g7!찁B��
����'�2�'���'4�ȟ��*g>ըJ� ����X9e���R�m�����Or�$�O����O	��A���I֟0 ���v�8ei��d��\�ÄE��M����?���D�O,�c:�T�'�X�"��XC�Q[� ��)͔ ��4�?1���?���j����r�iU��'���O�HI�@DX%w���T/H�p�z�h��dӊ���<���Ǻ�'�?�/O�i�*Z�f�0=���7E�+ٴ�?��?ƪ�j��i���'6��O��t�'{�� x4x�"_e�Ra��Aطjq�y�P�,���R�Q��䟸�Id�D�~��h��|��U������q" ����ĩ��M{��?I����'�?���?��ͤ`���*�/X�!�Fe84���0c2�|�Oc�OQR�{��@5���`��E��-OH7��O��$�O�ț�	����I�@�I��i���wB�ѫƊ�7Ah�MJ�s���O��Ct0O�S�l��ҟ�������ɹ�N�M*�HX2*��M�S*�b��xb�'�|Zc�I1D
*tO� �v�5E��ɩOz@�� �OLʓ�?���?9)O�mr2A�s�� ҋZ�D7��#�!�/$�'���	��&���I����o,tu*<J=T�EH��ԟ>��byB�',B�'��I)J_F]�O=�(Z �c��*ML,Z蘉��O���OB�O��$�O$�0Q=O-��#[#��S�+��eאՠt��^}��'E��'�剎A|�KK|���Z �Z�r@��!`���e��X���'�'���'�t2�'��R��ٙ gݦ"uR I��'\���o����	JyR�0^(��\�$����	u#��XM��hC�8��\"��Yx�͟�����l�~�~r��<
�r$��̀o��4��P�]�'���v�qӘ��O:2�OO�p��Aa� ��DvJ��u'�"�0m�����	0PO���G�)��=X��8-�#mؾ��p��,N|6-�&/�l៘��ğ��ӿ�ē�?�b�)X�9���\�F��:u�HT�vX��y��|��i�O `a1%Ȃ$�U���D�$CD1v�6��O��$�O�}	�NS��؟��z}b��8oP�� � xF�!�b��ͦ�&��r��Ƌ��'�?���?auEK ���W��W�����Ń?���'�N�Br�!��Ov��(����");Ȩȗ�R�5qZ�� S���1������'���'��O��2SIX4�r)B�FH��B��D31m�O����O��O����O���ul�%'���[Q�1�lQ�Ci��z����<����?�����D���&�'�-A1 DD��4����
�$�'#��'��'"��'(��'̖l�g�/]� ��@`�VG�@P�l�>���?�����$�+o�A&>U����3>���n9S H� 2�M[�����?Q�[>�A����	.�4��Q�B�"l�!���cܴ�?)����$�0X�d&>1�I�?�3�xb�ݟD,�d�� �-�c�8�'�b��P��e��rF4��� ��v�6��O.���Er�nȟ�	�p�S�?��	�9�:1J��^�Z���̙�X�f�ӭO��䛽aҞ���O��|zJ?M������X�+H�xH�NvӪ`
t�Gݦ���П��I�?�����I���b��Oz���)�=m�	����M둨�?�/O���O��O/r�^�9G2�@"�N�j\R{6��7��O4���O�9�bc��}�	��t���L�i��j� J0�)�W3�`���hi���D�<�G��<�OQ��'��ƚ(x̊��GrX&��BIֻ�"6m�O����U�Iϟ��	ǟ��������5�A���Z3k���b��Ugm$�[],���?y���?Q���?���?	���:"��u�A�a�䵩 J�7;��=`�i�b�'r�'������Or����Z�~�����(Jp���2���O\���O����Ox���O�y`3�_�1��̒!zlJ6�숣e��;�N0ܴ�?	��?����?a,O��d�U���˕PD���MSEN�<"�tP�\��ΟX�	�(�I�2��%��4�?���@E��K2L��Mϔ�r@d�9��B�i(��'�_���I�a����D�g���ht!�w�6��'F�
�8�o�� ��Ɵl�I2R��]�4�?����?)��w"*����Â~�JM��K�ج���i�"P�\���$��A�i>7-�4R�������O��buܬwHF�ZFN���3Do�6 ��I�I|�>1�
�|��eoĆCH�[�iM_�<qF+96(�ge���vx�!��b����c��xB��ꄐ0:(�F	��(bA+�g���&ة�"��~��8q�.�;5~	�,ۘ���IV�Y��l�e��՚��)
�j���1e+�-8m�iZ�.ޒ�� �ǯ��F�԰�"��:qm���FzZp�!s�/7O�P��}\J�P����?i���?Q�{[�n�O@�D9�9�ʓ��zd*U�ԁ,ɘ��I��9�LʿBm���ڟў��-��� ��CMG�q���YX$���/����K��BȈ1��
�?�=�!�]�O�����KXg��{c�j?it����	I�I��T�	OyrbX.Y�����΀���1!�8�y�@;�p ��Z�*�:��`,��e��#=�O��ɟ}��%�ش%��H��[��%�uFr�d3���?���?A�2�?����T�˞Q�d�Z#�>֡�RHRIܔ5��?�@a� �1�0=��La���0�ΖW�Z�ڕ��rh�� �;la�,�w��Dh ��Of=o�8 �,k�#��f�|ph�!H�H�4��'
"}Γ� 䱄�8��}�f*���!�ȓ	�4���V�sD0���;-�̓al�	ry"�R�D��6��O��ĩ|2qiG-�j�Ib��>f���sS��!�����?a�?F4���dD��*�X��$a�*�t�x�.[' �̥Y�v��l�P�	�>��X��>�yX�b�v�T�)S)��`4�Ы%T����\oIJ��	$d����[���4�?Q,���!G"B울�qc�>I��i�
�O.�"~�S�? �L{�����ztX��sQbQ83�'��O�,:���>��C� !36@�;O4�k�i1 ����O��'W\4Z���?A��Q��,�@Ck�1gG�� �j}�U�m�칎y*��Ab'�%J'�(y��Y$����BNR����������2��K�>z�ω`� -8��Q�A�ܘ�$�'�����I2���i���rv-U�A��a���(~���Or���]�1�@����	�$�;Lnp�t���?���,I��Pc1��+7��Yqėڟ��	Q����۟��I������u��'22�ҙq�Th�uN�0V2M���96m��DO-d�
�b���<[��,*��hO�HR��!t\�R���
���jf�C���iSe
>�ā�qK�P����6`���hR�N+��0�0��Z����wz���O��=�*OF˲�%2��}��ř�
4����"O0\��A�-k��%��C�^a6�z�����<1�#�F�gr���g߮i��u�[�6���';��'��m�O#�5�Hl�-���r�ɡsJ��a�(�r�x�A,�p>�sd�m�vd��y�&����8xuF���L@6i�:����3�R�'�H��#�;Y��x굄͊��@���'��Y�d��J�S��mC8��L�	�|�POݙ�y2*�H��T�g��"pP%J��yR$�>�+O�}K+���IП�O+�������lQ00��x�� Z�J2�'#r�B,Hh�]�G��6�*�P�&��O�j���1���b�tYL80�z�q��o�'��E#��A�V���TC��U|=��*د�D@A�[u��Ls'�=s��ek`��v�'�ms��?����?Y(��Q�X5���C�V=o������O��"~Γ&�싆#X	�v�#։�U�̬�����GEB��0"B*]���NI�Z�.�ϓ#]$!y�%�<�?�����)ѧO�����O��dK7b��E��M�4*����� Β-���6T��E�V��|Z���3��RT<}�x�G�]+`鴰2�E��p��w�S�O
�S��?�bD�vܹp��J�/���᲍Q�(G0����?	�O����O�A�C ���@=�CI_o� 3!;O��6�O~\"�(˥b�0�c�[�	fB�+F቗�HO�S�g���
) ��j�D�T�B�I� !S@$���ܟ�	ԟ�b_wI��'��xRa�AH��� Bk��1�PI;/�F)wo0�j�(�]����	6t�01��V��,9W! �`� :$FB�dDʈ!���@5�x%��?�n��V��b��1���^@$�y!��E/|�ѷ���4�D�̟���ٟ��<y+����E$ ���gٟ+<�@p'm�P�!�,��2�
�%���<W�h]8a*1��|�����D�Y��m��/YD���J��i���ۤ�2�6���� �	��8����X�	�|B��Z(G�l�ʑg( �؍���I�hc���e� 83a�S���<�Q�]�S�@�b�/܀�� F� a\��@b�t/�IS�Kַ��<�pbRܟ��	%\Xn� ����:�����+(���II��h����N^r�A��"A�jp�:\��dP�|6��1gҗ��@Au���y�̤>).Obồoͦ����@�O >�(�bj�4}A% CD�"\�E*"��'bBOȿjֺ��B��X���v�~����'Vf�ę��!jO,�: ���TFy�H;o�� C�8j%�a�&�0����;t�(�tj�5 ���oիa�ܢ<�ʍ�������Ij��LOf۔��������'nr��s�� 2��`�bE�#����!4�O��'�H�*�[��ZR��W�n4Q�bp��UH$����O�˧J������?���7U(tK O�q�ԈB�
"*�F��c��+3�(�i�I	��f����i��x�矶7
޺'u��xs"�2��a�G�A���]��}� �P�MHȢ~���t0��SaEM�^����V�S�p7����P��4��)���B���e#��� pd(yn�,c�z|��l�]H$�Q�>�T�X�]% �"�Gx�/� ��Ɋ*S�hK�ˏG%�xEm�*d����⟔�a$E)L�<��Iџ��I͟�p����dB�b�p���Ĉb7n8���8b�$_6'B���d�=xmf���+/$�L����S�D���o�����J�>�88dL��;�r����?9��D�C�t�$����t�'��Y�8z'{y-��%Չc�qz'� D�ġ���� Y���5Ɠ�PL�}��ß��HO��0�'��I�T 8ͩYwu���/F�z���Un1Y`f)�"�'�r�'�B�),~��'WB�n�bZ� M=����w���8��9k���J! ��@koz:��Ǔn��)�HǱKT1�2I
+�l�5�U5{��5B@��t��Jh��уg�O���B=,fh<�2o�,]�\B��p�J�o�͟|�'���4�d��
>Uv�D������`A�u�(�Dz��9O� T��b�y��:0�ӊ\P�*"=O��n�Mk���'��'�<���ߥtO�ݒ��BD=��'�f�:��^1�j�N8N��E��'R* rS�KHd�q�I�1B��Y1�'�4��B%I>d��b��4$�ES�'��I�W�Ҡ9�\I����+��*	�'S�l��I
�f�@+�h�������'�����%K*�t�0��6v [�'n�hv�&jw����S-2
y�'��j%C@��P|�T��'��AK�'�R c�x�i
4b����{�'�,Թ�c�%��I��I�F��'�.!�U�_(���b�2.�H�
�'�Tɒ��*���2��6�����'�v�!��v��a�[�%2��'9P�Kt́�J_Lţ�!�~���'�RК��Y=��sR�U:
�H	�'"�$N^��ݛ�E�����'�L����.�L��1�As��'o@���1(Y���Ȉ�8q	�'4���r�C�x�ȴA�h��,��'�b;���+k@L1�%g�z��9
�':�ȱcQ�se�-�%&��FN�	�'�b��ٽT�T�uh\&v��"
�'�
m�WmA�LR�k�Z|*	�'`p%��ɗ�:��{�6Tx(�(	�'?H�b�p�*������Q�X ��' MS��Pक़Q.;ߦ�X�'��iA5��2�LXmYb�ȩ�y�Zx�n�9p�	�zS�U3�-����	3lu�9�b�K�&�F��˝ ?�Ui�O<I/d-��ʄ�yR�ѻD�ڱ�f�V�NHk$�C�l��I�[?D�Ha��e�|�<�T�U�P�Bf�y|��{��Yk<�P�=s��t��OƉT:09`G��c��$�`pȞ2wGr$�e�I�.���:�B7�	S�m��D�-ЎXcg�];Q-��d�f�n��r�
smڈh���iV^� ?@(t�w�܅l�L`[�E.	�����R'=G�\�
ד)��%b�b�$D�HYf�6u�'Ȉ]���B,j$
0ŜLRM3���ǐr���(�,�;�Kr��\l!����D�býkCcK�Vxp&��E{D�`ǵkG�ԟ���Ee�''�󮃊-��;W�!*|����W�i!𤓪]�ta��*D�yD�V4=?��Ý|B�F}�����Q76�ѣF����'a���J 74��nh{�u�	Ó� ��E���4k�A��˯pVM���^�6����h޳�:�z���l�4hG��a	�<��#\O���"��PF0�mY�jd(2����bb)ʒNU��R` �}��4zG:�i����
(ҾĚV��6^����9D�DkfA��r�J)��.9�e�	F�&�䐹��O�t��$�Py*��I�y�+��'/6�DC�L����T��PxE�3
��ЭQ1�*e�.D��(|�$S���<�& P����d3�%�6��U��p��	AR�,D��0ʀ�X}���I��E���C���>�W��"l���̿l]D����K8tf�EL[�{�a}2���<wB��	�W~��kd���Lsl�:C�X3C�C�	0@eY3��kk@m�oڊ(�#=I��/O ��}��?3�`��Q�#������Vu�<a@g� vA��gnC1����)��M�&]rqO?7m"T l�j�pu8�	S��?�!�D<u�z�K��ęm�8�)��W�Q��I�L��m��'�������D��qR΋������C�,�����O�1#���2�������N�U��"O�( a�L�}�P��k	� ���:���)���b�S�D��塠�2H�z9�`0�C�>zu�Sf�(�p����,�67Q�.��-��{���i(`xȥΚ�g
�iv(P�G�@��'DT����Yc����!�?efp�O�Qr憨��=� ��#�PH��F�Z�Wo8���>��N�������ry5N�Έi��M�?�� h��?5����'��iFϱI,+�!4OX\��y	�t�X]��Ŏ!D��̂Qyr՟�k��@ Ibf�x��\o����O�i��ɭU�� �� �okI 1�J<pN�7��?$�AX�eI��ɍ�H�b@V$�,	�&�H"?�p-	��®�0<)`A������+I�%�0�d; qv�C�	e��[�S1��o�d�x�O�^a�!*�#Q+�d � j����DW�\֜�BL<��h���'�@,�*��d=6iX����/<�|����Sct�
�c���Px⋓���E!C�IS�l����H������~&r�'�|p�Q�Ζh�bJ�SW���O�p�8��T*��) ��!��r�'Wp�:g务bx����I�f��8JG��?�%��X,�k��C!t�Zc�A��S2��I�x��3�b@�b����@�\�d���D�V��IH������gQ2)YSF�-��9����+�s-��u����悉������'�H�[�� .]4�, �.Ҍ%�x� ��5��A�"pj"�Zv���MpHֽ<�{���d����	�q3�M�\�ܴ�4�Z��Px��Ó2�T�4��668<<�4�[}>=+�����è��i>�����O���;V�HI3�.��yr��(a�>��ɳ5F��a'$�����+G�9����A>�\H��H�����u�����?J֎)q����|�'O���@H(J���1�ѭ$���s��d�;��1"ѩ��((R!kă��0O䁈�Lt�Ti���m���R�O��?A�@�qJN����	�p<q7���>~8`(Cb#"0���7#z(���r��0p$
�o�|1��Ɍ.������&J)�lR���!=��#� Ƶi<�5��@�_K&-�B�R�b���ǲ	���wĶ�a θ}ࡁ3�M"7�NA��q��SrR"[d����tx�d�V�N���ط�D�'k8@��#X7ty�`�F�f���+O���i� F~|��P�
�`������	�V�2�)B�ØA�����5bA��pA�aPI��/w���t��+5. �l6@���vO�=G�P�
���O�C��R�{��Q�,�W� â��dͬ��E��xC�M�Oq��I�j�q�G���T�"��S���h�N\q8��Q%�"uj�Y�wV�85�H�-�j�P1�A�	^.1�`Ūs؀��5Ӟ�=ym��K��-��(	�l�+3ƀ�d��5h�d�m�db� [�M�Y#$�1��8CbҬ�U�4�7FZ;!�ệ`_0��H#�N,[$ݪ��䓄�B��sўt�.���N��6�x�2��Rc�vf���aC�!K!�c �k��ybcnKߟ��@F���To��̲%� �%��G���F뗎q���)�p���Y�(4~��	#5rYB���L���d�L	4�`��V���`��Kh�J�A
ުK�KXٟD��O�J�c͕"���i�x`��fS�0 +H�U�"�B�.g�&T��	�7����E�
�n�	�
�%�*6͕$C"��r�N4{B(Iр��5�\�C6,�>'nE�!��$mh����!��Qx�#�/�y�ݺ.w$��Z?�x��g1�Խ��eB���?~S�;���6n�2�;FK�_���3*^m�4-�C!4�������������z3C�o�8�I����Y௖�q�0�����E<�62w����OJ�p�j蚁�򅒗���G�,w>�P���	��x;u�]���s�%
(������%"�t<#���P��Hu@օ� ���b^�?y]:��E���"�m%�x�5��%" �5rt'�*=nR��Ԧ�5}sxX# T3G�r�D��]�Ұ`ӯT��;1��� $�ԡOc�'%���,ȩ�(Eb (цN���۴B������o�p�01
��)4��x�h�$�3� ͡CT@?yB��)p�a=j �/4��kU�˒!��Qǭ��,˓nˆ��L�&F�I
��xZ�O�Tp(� ��$|P����3En5�2�*s���F�Ѱj� ;�'�P���2�R�ɩb7�q�2JݺGC<�J�`�#>��97�#Ԭy0��T��	3��'�0}Q�FĈ#���I�l� C���;3�~R�!Lu��d��(�*!�T���� ��S]�^b��̖$����&
g
��u"�] f|��`A ��M�Z���w&�]�f}���9O�-K��\u�T(GNƀJ^��ū��Kx�4PSb0O�R�*�]�g��:i9t���,�d�|��.C�e���K��o��( C"�'^���X���>IM�<i� [�ARG��1j���띛��%�݋��'"�yU���#TD�	��O�#�ͻRTl�@�	�lc  �Dm�A8N�+�O3~Ğ��*�n	�'|�<Óe$D��)5���k�'Δ�E�ΦS�
�X���@eb8��D�0d�m8���k�4��O�ϧ^�8n��R�q �A�?�F������Ĥ'���ψq�z�����)[��)�A�9V�m���Ou�d�B��:,�<�c�H�v�s��Ӷ$g,�XA�a��}��Q#�lIv��Up�x�EJ;8���;G�m�׈n��`��ņ1iw��:(�����+��S�'����C�`�6��ܨ�C�*������SX�'8�C�h�v)�����)D��if��O�Q��n�5��I��>��'[\��El	��~2�J�7Cح��6���IcY�H�.A0�B�@}l�s�,!I�����Υ`�f�bG@	�O���G�z�BǄ[�Z�qa1j ����t�L	���O�P�݃��O`u[����B.��Y��L&2��)�rF�U�ꨆ��ռ� 
pؒ�ۘ��$)gW!%P���mټ�[�e�P��=�|E@�"\V���T���{����	�0�X��'��	���G$$�b%1VO�"m�@%
�g��v�I�s1��#�,6Q�ܓF��<).l� P ��ي��@"R����'y*�Ʀ<��/եT �X�
% ��������Q���"��T�f�x1�iL
#���T�M�W*��%�	1^��-ٹ�Hq�#9>,���	Y�,�t�	o�QA���7 r�,���R�~T"����5�0=ab�Jj��%Y��ӇL@�P�� 0t�W�(�PЕ���<1p�G�h��.[�D��U�H�G��Q.1�l�kK�0zpR����"�
6| �OΞ�2�'��H�"��R��)���[2��'�ȕ��Dɧ^g(ِ�( 1�}��{�OLdPӬ46�*$�)ӷ ����'MZ`!��S�Y2|	��'�LeRפvQ*�4����'Œݹ���{)t���(J�x�Ɲ�Q$ɽ+�(����O�t�O�B�+���ې��3�m�c"��?���\��l<��'��c�J|�S�t%�&>�
c5GZ^6(X��=U$�xB��L~�͟(1� 	�,�8rcխ3,6���R,���ʶ�C�S�$�֊�Xm(Dmׅ���[��� ˋ3�T�􋉈9�W��r�~MbL|��LT�\l ��pW/Dπ<����n ��0k�=�y�سK�<q�J��A3&�vG��ONX���V�Ps�M�yp�za5O�8!5.a�T���'�NY���1kQ w���p�x�'�@�ڣA�����8�rd#)mܨ<�������[�/la��ҁ4�d�D&�O�d���X^(*E�\&����T>}ۂ�ZN<�fN�q)�����r8�8:��ɫ6>�)	��L���၌0sX�h�k��PnqO�ӹ���1&�9!��ΓF�l��,�#%��@AF�6GA��O� ���T?iql�2l
q�[;)���7��,#�L)�Ř�<����8���0&hڴbތ(
u�Km�'h�ʙq����d�2���4�O�eB��S
'��d�'�SH��d��O�ɠG��M*Zݸ��#y�( ��ĉ,��O�q[�AU�[�8c��a���]~`+RA�^p���'k2�ڌ��F�b���/�8:F�c�����yw�T�h�U��2��`��#����ʸdG���[O��ħ(>l��.śS�h�S����m��Q���4>aB�{�^��9C%+�'A�rY��gG�1�5��2�x�P���\�x  �Juf���ۂ�����̏�s�D[GVM���چ �����c�>"!D�s%J�K����%��Xy2ǅ*%F<E�;��Yi��X(�M!̙��j牣J�4��'�(4����V�?�<����4�;��A�z���J;N��%
W#��R�a��,V���`CJ�0�Ұ��R6z����a���ZV,��]5X�#9�P"<!�j *OC@|#��HO;j�6�WNy�%Հ��`��Y2-���I�<!�Z<&C���Ee��K�L-�g�q���a6�K��~bb��~�@��yʟ�#�d�Q�]C�Xp-�3@�!�d��a�xk��+}0�85��9�-�9�M_��K%\b��j�4p(���6'B�l�s�(D��4��N�z�+�"��/U�I:��*D��򂪆8Y�<���A����ae'D��#1������!Pa��6�)D��3p��,~�L=�恵M˲��p�=D�@���#a(�Q�A3}g�!Q�L.D��"�ė@�H��-�u��Qt�6D�� 0���f{@p2qa^�mh��r�(6D����6�H�� 3�t���֥H!�$�0_} t�m�p��#M_ c*!�䃲��ӡk�?avjI����J�!��DZ�*��õ&p��Cw*�7�!�#K�P5[��W�k5���k9Y�!�U������j�s!j�'h*!��]4.k���N<
�&-��)�" !�D�e�\�T�A�i�L0:TIݏ�!����#��ǻ���@A�O�!򤝀2ָ�[�ˌ� S2��E��_�!�$�,��kPdO�lQ�^HV!�dY�S��*�� �`�0C��0D!�D�`�"�j֦�a=@�F�<A!��|�X4����6"ؠ�К\=!�d�&����邐t��	���W�n*!�$N�Aʈ��T�f^�ɐ���*!!��9tT8�#��ӠAYр�Z8�!�� F��VJ�Q�d()�&�)ox�!#g"O�	��ח)\|�BE�W�=bn�"OxX�,X+C:���/�,�c�"OtI��֏vW�i�ሂBA�h0"O�x)�C^�~����K2�n�h`"O4h2���LoP�&dĦc�bzp"O���A?H �\J&b'�^ɓ"Oj}(�!�R[��T�4k��I�4"O�Hf�}�@��%��&N��Œ�"O�h�TNJ;t���T7H�- "O`h �ő+t#�@c$gP�v���B�"O���q��#�Z�S�&÷^���2"O�@15Ό1c�@��QD��^L�B0"O��'%
2q�0�P����"O���/�y�p�����L�"OhL��
b����"E�Y��aj�"O╢�Р0b�tH�[7*�P���"O�ѠBٳ:��@{w�*�Z|�"O܌�!��4+�F�ʓ�B�A���E"O`�@�1k�1r�F? ��R�"O��S���1�Z�s"�=n��3'"O�q��N�0B@��Ir!�5;	��J�"Otq�/T�A@��W���(#%"O0�;��� ���P�'@��0"O ��GT7Hɱ�m�6Q���"O��p�*�iѰa�ԬQ4���s"O�Y� ��]n��L�!{�$�h�"O���'��s'�\�@L�0�LECT"O �B$�&�`��ίg��}��"O
�H�'�
!�V��vH"O�-��"O�X`�
ϙ!�\����V���v"O��	 ��-4H�d,�̴4�7"O�	��,����:q��d�r J�"O^@���[:G�ఒAtj�tC@"Om ���.��3&ti�5)u"O	:v*^>F�8d٥�ʳgP pF"O��'��6d����6��k%�"O�͘�
�$'b�bE������q"OjP�ף�:J���Č"]v���"OL9��bL�*�l�AD��bΠ�k�"O0�&��8�t�`51�r��"�'��'��x�aM�T�F�(�(ůcm����'�����O���TR��J���
�'X^�1���3�FM�"*оEiF�S�'�P2៦^�M��c�2~ !�'&�J�F�;��&�Z���l�����[�	��=i�Ş�0ĺ͙����!�d#����K B�n���l�!��2	��krG�*��̐�F�&Q!���1P�� {��I�1�J�5�!�D��2�J�7T�}R����q�!�U�)���BwiW.sCJ�	GA
�2�!�VU`�(s�˟:c.�S�I�w�!��LŔD@�K_�-��{����
�!�dЖ74r�����,@�H�5[z!�$�*���
:R�U�r�<5d!��SV�(WȎ:+�@���\�/!�D�>$5�=�p"�]T�ఠ+U�!�D���D��@G-]���2够%6�!�D�!;&!�t�20B4���!�d�]��͂`�d�`������!�$����9�[�	��٦	K��!�$88FMv�DФ5
F)\�5b!�J�24�ģ�)ʼc��m���:�!�� ��8%G�>VG�(#��E=ep�A�d"OxY��"�b�*��#â�"O 5/� +� ������H��"O���F�۸0ڐ�L��"��Dҵ"O2�	X,$�(��Eh�ua��'%�	�I'�,J���x
:�"d֩_?�B�I#}��h����~(>Q	�U1n�B䉟[�45H��+���0�I�B�	�*V���)�KϪ���@x!��@<�ReC�[�4�s��x�!�dO�FW`H;�d�3� ,9gA {!��*68�E��
1������7�!�Č#i��X��T7,��;�L:~!򤕊3}�I)BL+w"[%��$yv!�dA.Y_V$pѩ�[qj��"�E�!��D�Nِ!�2�@)�"��G1O��=�|��^#�ذ�hS�:%��@��u�<�'C�,W1���㙠[�p8�AAt�<��	d��b�L��l�S��r�<AţQ�"F��b�		uz��Rc��l�<���ό<��2�Bć$ANPuk�<��*��5���Jq`݈+`H\���Zd�<��m=~8�é� OŪ��c�<�g�Z�l�j��K�d"UI�f�<y�˃(�~=1U��:���� ��c�<AQJQ%A|�aq	Q���T�c�]�<��JFI��x�J<R�}����U�< $��0� �W	L��9k�Ny��)�'\�Z��%lU�q�6�J�W��9����|C�D0c�<�`٣|X}��&�d���̆�K�P�5#�%�zx�ȓ&:$� g�Ζ,K�����N�f$Jy�ȓ^���1��ý&��)3@�%U�Մ�	J�*C@ՓcČ4:�I�5$:��#�r�c�؇*���ЫZ�F�نȓָc'�.C�d
��P	d�^�ȓ2���G @)`S�4� ��7��|�ȓ�j����%�XHq$ş�0���Ia�$�����M�l��!�ĥS�}!�sD��o��
�a0��Rr!�Q�Rpb��"�ȍ�
1b�d�;G�!�$�j�I�ˤX��SiȊ!�D�5>�y��� �Ɣ�G��]!�D�+K� 
���&�}FhT�-;!��P�� Tǘ Y������p !�$@L9��C%-��1P���B�!�e�z<��Uf�ybe�I)R�'a|#��2�
 ���	�
�т���yr��Om�D�+2���a�P��y�f�H��H��F bb�� Z��y�&s#���6�ͱ%��<�1-���y�	̲E6,Q!��4�-z`���x�kѝ�x�� !�4}Kj!�`�޾�JB�I�,�J`a���!p0-8'Q�MiZ���*}r�˱X�*��_0+����΅.�y2��|� �c��.-�АX��ʡ�y[�CQR�+p*
=$>��:`� �y����z�H�.����}(0MQ4�y��D"�l-I�e�.%=-��ã�yb� �/h���KF>"���f��yRb\�t�q���M ~�B,9T�ֻ�yRƍ�D*�Z�AN�"A�hT����yB�ɮ��!�����d��y�*P�Q����ǝ>��l��L�y
� �A���ݤg��	"gY�q<Ujp�O���$�E�踁�͵>����P��
D!�VɄq����O�lpie�M:!�$ޠeJztB�Ė&�Jas�#ׯU�!��R3v��<@�cA<h� (��0�!��ۋ)�8�'b��H�d�At9MF�Ob�=��l�r�꜔/�:�Q��'E���#Oh��@цvl$���?~��i0�w�<a�K����)G�2@��X
�p�<��"�y�Ra��ժI�����$h�<��]V]�����8U
bl�a�<�1� 
a`�s!>{��̉���`�<aU��4|\x��Ń�v�:	�D�f�<If�@t���R�M--F
�*Í�a�<�1��\�aZu�^&p��G�S^�<AG�@�T��
�.O�Y&f���`�<��ƨQs���g|	L�� i�W�<��胙'A�Ɩ(�2)�Q�	Q8�lyQG�l����%
2%a�x&-$D��R([&�N��u㝃���b�`>D���GIɣg�ty�#V6k)����(D���C!F����`!���?A�tKN(D���`RL�X�4Z$�����هd��hO���F�_�<!%�El�r�"OQ�!�I��T�����N�tU�1"O6|�GA�T��\�j
#5,�U@"O*�#M�f,Ih���K+@�w"O���իm�Ԥ�ӈ_�r*��"OĈe������� ��BI�|1%"O�� ���s��dS�b�#;�D�C"O�F�����DG�$J��@w"O\AIRԷK��܉t�ЙK^~�J%"O�d)VB�?>�ls��'_]v�a�"O��f�"��{�E��p[����"O:i�G瓉-4��B�l�1g"ONT[tf�8)e �AΩ7��|D"O�9�ulZ�@�s���7��`!"O�!��ȸf��0�CQ�b�L��"Of�@W[�1����p��2,=蔁�"O���v��5|�x�hԃπj4��T"O�=�Rg��[dl���$��!�"Ov ��DЏ6�D50�d�4u��y��"O�L����&� ����ˀz��u�C"O21�F@	*��5z��P+��A9�"O��� �]1��]�P�ũ$����2"OF<X�)ˈ��v�ɸY����"O��:��c ���YAZB1"O�ؐ���Z5�D�0M�kSZaRb"O�؀��	�	d�i!�l�(FJ�I�R"OF����b�МH􋚄!�X��"O�uzߤ%0�O��7�����5D�dx 댥	�L|edlb��i0(5D��C����`|9�#fŪ/E,E��%D��l׾~�b�K��X6�����!D����Ƃ�}�|�
�V�	���ql=D��I0F>5�r�C��>���d�;D���A^ (3T�Pm=J�Z���H9D�`+�A��y	�3���^c\y���*D� /_�\����.Fs
8r�h%D���LZ�BZ< IA�R�0�l�d/D�t3�CD|�
��a�N�
���a0#'D�|�/ă~Q����5I��S��:D�x���a��{b	M�O�Ѻ2�,D�Ȩ�MW@���00fL!3cv<y�*O� ��9��J��aH�ˇ&�lh"O$q�$�2@ꄭʅm�)��m �'�V �ӣܣ�`�c�&� Ƥ��'��Q�	A��J��͒T���'�*����V�}lu���U�x����'bv�MM,vjfx*��̊��Z�'��쇭y&J@��
'�~���'�bP��>|�R�����
w=1�'E�$I�
��[S �i#ȕ+
̔�S�'�*�@C	A#S�
�����}���J	�'M�WR7�N���$�%x�ZP��'�N]�DD�{dz�ptA�r��ܸ�'�!�5G5$� uq�D��f٢M��''� �1�żOQV9��c��]X�'.����܏A�d9��MP�qQ���'�*JVbЛ0M����pL���'��D��	z@�,�p��/5Ϯ ��'*ք᧢�y��zO��C|�Q��'�� z���̦(b:8��̺
�'��A�@��)�J�[��(�~T��'�8��	�6�Ը�+�N�<A��'9z�۔ A;x��[�˱�H���'�������v������P�
��8�'�Z����C�%�*�ҕ͘).�h�'h$J�E�;Fӆɒ0�� t;�U��'��9AMH$N�S�
*s��A3�'X!C�J�Cc( h	S�j[Z��'��D	u�ыXR�E�d	3e��q�'H� E�R@�(���]
B,��'��$��&w�����Π�~P��'� x��_,3���
*=�1�'�:���~�=���ۉ69�9
�'�(��4
5Qˆ���)c��[�'.j!��m�;o�9����3X(*�Y
�'��У��2���%H>H���
�'�. �PPy �:��q��Ą�,��*�fT8-.��x B{%��"O��a�B�s+P$s�������"O�����R6V�FG�t�|���"O�yS�Eλa|���B4@�@��"O91��Za0�)b����U)"O�r�Γ']�؝jšs�D��"O�H�gX��@�G�#R�"�"O.���o��V�`"���5Fh�[P"O.�zGd��ar�Q*�9TP&Ċ"Ox	�&8N<H����C2����"O�A�-J)W��"m'D��"O�ձ7#F ���Ġ:��ȸ"O���#]�񞰂�dE%j�p}r�"O�)��E�+׶��cX�q>��A�"O:�Z���!]���sc�i$�Ij�"O\�S��~���⁐�>@�(�"O$��f���pwFޣH�苅"O@Z�� Z̳�
K�Gf�l��"OJx�a^�Bl�9��J�~U��z�"O�9S����6�Z�a��b�|@V"O @S"��@�0#t��59�|��&"O�Pr�S&l<xa�A8��"O��+���+"�fP*戎�}�Lj�"O.�@����Y�U*C�p�`U�""O$�	w�^wR������D���"O��$ξY��{�(��Z�ţ""OڑQ�O�B�B(K�T>]�"OZ(�AJ�6�f8�ԅպ��� "O� �hsUb_=�N%���)��m��"OR�Y6N3j��D���� ��lS�"O�y�v!p��$� �^���;�"O����BR&m�fA���h�؝�"Oa�q�^�D�L��60Ѣ ��"O^tQt�
$��l�����X�"O<���`�#aY��'�E�V���"O(uC.��֊J�>Dj"OE0d�H� j1J�M��	�D"O������5�Ш	�F�
>�FS"OJ�3�*$L�΁����?l�n�(f"O�x�*Š>��Hr쒈L�Nt8�"O��*q�Z�� �K�J����#"O�LZ&��5!Cra�B��� "Ob��	�K�6��m�4@J%���ȓt��P���t�%�f!T#<j0���Fz�%�u��4�������"l� P��U���[`��(B���p�/!o=���D@�[�Xb�&�8�H 54.4��jW� ���JVx�C��	SI⬅ȓFl=�����$����&S����6!��wj�?s?���H�E�D�ȓW"`�J��=q�H��0D�=](��ȓmX:�j�F$S�u�$c1R,����V���JW#�%i��yQ�)�� ��ȓ!�l%P�Aֈ/��]9����|���Z���Cn^:�:��� Qڌ���1TY���ܺ'g�!4�X]�V���X��)K�M��z���c�G�w��!��-j�Y{w�\�
m���Q��
_ĪՆȓ4���JWJ�-3�$����G-�|��k����W��%*�Q'Jnw�,��+��ܩ�˛�V��h�n��b�
���"��Bt�4a@f�����~�D�ȓ4K���ƈS(n%p�/Y9#괆�)j,4+�)E��D9!��7�z���80��!e�
G]z����7}^ń�1Nn�BM�1!r���RMԘH'�1�ȓ!N�y�� �.���->�ńȓ����#_�y�  `�N)���ȓ7�6Xum�<mQ�nТ>�d�����3CH�<}��� �,�J�]�ȓ<a�(��G*S=tB %��	�>�ȓ
H�8K描��\}�`dM���ȓ-��f%���!�fn@�J�bE�ȓJ70iڳ��/?�����߫H�p��X����Qb��xg���Y�b1�ȓy&��mZ~���Eݎ�6}�ȓH�T��G
hU�0x�'���$��`�:�E�M=�H|+�MV�]��܇ȓf�l2`��N�0ӵ�J�m:jH��_��m�t,��tke,�-Q��8��'��h��nI�W�_0��Sf$D���1�Z3�ȇ�")�ph[`5D��҂�Y�W܄�ن��.F�N��&!D���-ߋL���aR�۞A\:VI=D�<C�윗�V�21��9G�I�'D�lB'�����e���l=��!D�̱���+O��#[>b�F�"�>D�l`�C@KE�]9��d�^1���)D�ȒTm$v���àڿ9�Z-+#D��0���'7��Q��F��v�Jq��<D��Y1
ٸ�e�2L�4C��A��*(D��`REF�6Sȥ�7#�l$��	e8D�� bL��d֗kQ�i�e͕#/���J�"Oܓ�
س���h�nH1tE�T26"O|�����Z�E��--Z��h��"O���GK� �l|{ �F�:>��&"O.8(e�Ōo�tp�rd�W+�!��"O�@���,��"�	��P �"O��Y�-�-IR"�?M���"O���52�t��F6�t��'"O��3� ��r�ķ'�H,d"OM���ϟ����0���p���24"O���HD��d��e�;xh�'{��+��ܢr8�!
���ԔR�'El���� #M^���0�&
%���'���)��ۜp�`(�NW��	��'މb�&�H�"�#P��U��E��'�&I� ��J�{��T2OB�X
�'/@D��Րk����u�bb�	�'��%A�(ޟ&ju�W����栩	�'�8r0m����A��$*+�0�
�'Ȯ�z�ɔ�@N���a#Z�a
�'w�Tv�:;"+��O�=(���'��`3#D:����E/^��X��'�);#GX&�Υ� �'V�$��'�H9��X7��qi	�\uV��'n��QH��qP!� Ns�(�'���;�p��G�Be��'��p�NE>�	��AìYR�'���&�J�#�Ƶ�! �,<�x�p�'���#�.*��0A��h��(��'�t�p�C�{�ͣ�k��b�����'6nA`n&��U+A��E�����'�M3��WEh�@�%���x�'�n��4�+��Ǚ�p߰��'Br�����8H�"�3�DA�mGI��'����E�/��9�iQ\
����'{>Q��'�~f�h��!g|<�
�'�4�u�e�f-�QJ�K��q
�'tE����k�N\k�6��p�'�������QӆTid Q~%�E��'��`�ǩGY�^��CLޥu�v�"
�'e&P�@�<�B\�ä�v�μ��'$�m)gg��R�B��a�t�	�'?8� $صN} �$�`���'��JR���zM�u&_*WF93�'$1�"�"q�nH �T�ܐ��'��b7KF�X�Ω�Wl�`pE��'=�� _� �Bn�)z��bq���y�e�`�|R�����q�ڬ�yb/+ɘI��/٩Q���!�f�6�yB!T�L��s���C(�՘��
�y"I(h�d8�@��e��U�fk��y�	Ϯ0V�憗 Z~���Ã�yR�ŋ1�$��/�g����v#ߵ�yRjD_�y�mX8I#�e��ȋ!�y�D'���z4$�"��X�⤗�y�ć�K�EI�/J~֖����y"�ҐY7�Tȇ�_�q^�j�`�	�ybH��_\VUX���6JHL�eX��y�i��D��!�jKC¸A����y"�иy�q�Q��+7"0��C�;�y�g6A(��E�H�8`�@;&bۉ�y�V�W:}��΀(8� 0$�y⃅!R�$���D7K��'�Ů�y�ŝ�Z��r��$����C�y
� ���iR�]������V�K� �&"O���k� NN��%n��J��%�w"O4���n\4^

�@6,y����$"Of,h3M^"y!��J���k����"OH���!U> ���AB0Z���c"OZQ"��֝f[B�x䁒AD���"O�t(bO� %2�uj�7v1~��d"O^�9�LՎJa�!���N /)�Ҁ"Oy��3�}I�/7I!��f"O�]i(��S#�����G�����B"OZ��"%��d��9�@C�A�q��y��ۭ!��C�Jh��Y�L(�X�'�2ɚ�@�"s�j�!>>����'zlP��l�	v�Z��C�<.��`�'�F���.�������4Z����'��P�" "d�����G�)�d�'���Yj&�JsV�b�n���b�<q��G9T���{���2f>~(�6�\�<sc�<\M�,c��$&�\�t�JO�<9w/����*+��A�h�ȓ���1��P)l��4�{����9� �`-�R2\bF!�]���ȓQ��M����!J���/͘n����j����<pr�=����G��A��YPБ���K� Zd���h�g�ܽ�ȓ.%Z�KJ*i�u*�6�T��ȓ�q�&׊+�,d�d�|[n��ȓH���r��N�yR!���\8�|�ȓgd����H�.��E��������v0�=Rtg�wҢ��!�L Iy���ȓ%��Ig� ��DZ�%˹*��ȓ ������J�hˆ�7?~���ȓLb�����"�&���$����Ї�-;B��F]^Pi2�'=0���4ը,yp E�	��Rҍ�T<�<�ȓ!�
9;���^�J�j$?�Іȓ[<L	Am�[nz#g�/+pH�ȓ
K���2G@�pj�)C��ʕv�لȓYNZxvDO'$�4�z!h8����ȓ5����)����qA�0@&̆� �-�T�ܡG���M.d8���ȓT� 93��$^|�lK��`�<���B��� ��UN0"��	4�T�ȓ&,�9��-Z1�݂�煂T�`E��6����⌷X�T�Z�S��\��0���9$H�?wr\���?1�\��ȓXJ��DO]�XZ�(`Δc�z��ȓ`>.U�ϛv�l�@�::��؅ȓ 9��eF�oĲU�G����ȓHjʙ�ĊA{�xf��1y��ȓ3�x@`�d�3꘸S���)P�d��A�I�0�RRWN� �#ub���*BF�(���	G��@*Q�I@�(��F7�Tc� '���(a��L��r\y��$�X<�|)�.V�!�u��e~جCĥ����/�9��(�Ӡ7D�p��J̾G�T�� D�)�v �4D��Ï\P�-8��B�*��e0D�dk�.��I���"����j\�	E*-D�L����"7 �� ҅��+�B&D���`�i��IU'g��Yc2D�x!�T G`�a�uk�M��=q��;D��"aiG7D�x�sC�ԅ;2:��`%9D���`Kǲ[���o���(�5,5D�� $Q(���<|�e�"Q?Tt`v"O��"u�&}�����Cp�>-�"O��a�͵I���ɷ�E"�
@��"O�i��T7����Bž9��!*�"Op���T��"! ���*΂M�5"OڌA�Od�<a��b 4��U#r"O`" �v�N�sF)9�yB�"O�q�V�Ӕ{~��3E����W"OppX����HSk@cs:0	�"O��+�1y�=QcN�%4|�G"O��H��ǐ^��Ux���LpR�"O������ X�s#��j��h��"Ov�v_9�fx��k������"O�0Qv#Ʊf|Y�Ӏ�?+� ���"OJ�C�Nm#�A a@^�{���B�"OZ�9v���1,X�{fܷ=����"O���!
?K?0�9�nWv�|H�"O��%��K���a�ȡ�� x5"O�13F��0�&p$�4@�&�b#"O�p�o�( J%�Z���	Z�"O��&%��K�����_/���"On(�A�g���i�!���"O�x�M�5K�B�+��K��:Q"O� ���V	Y��� h�>�3"O��;1K�!k~dD�"!���� @"O���DI��K����a�9}�D#"O��d$�5%X�x ��21���"O���k�-n��Ũ�
��C�"Oz\A4D��6(�]zS��3^ΨQ "O4�ɒ
ȏ^���!�[n�,{d"O<8�'HB!ӆÆ'z���q�"O�m�E11���q�"&�T`P"OY�@�G�>�\1��D@�[$R�
�"OU�cAڊ+;�� ��V�LU�"O��H4�ޑ3�:eP���`��"Oލja#�>1�Ω*�n܏D
l3p"OMjPh!4^��%��%�E�y���/<ߌ����!l��Y#�.��y2�O?��T����m����KO��y�ŗ&p
]i���]�$c4N��y��ȥ$��P��_�S��e�]��yN�&���됆<���JEĕ�yB�;�$PEC=I}:5ZtG��y"�ٜH��%8�MػG�%x6T�y����F� ��)VDP�-
�y��M���`e��5U,u�`���y�mۅg���6Ё(4�����6�y�&��h�4�IՇ�0��dPp�[��y�'=�LAPĤ���Х �Bֽ�y���(wm�y���W��^Ԡ�����y��G�
�����(p�[a�\��y�!�2d�x@S+Q,P�jX[Af���ybbC��Yc&�0]x���O��y�!Kc4�2"hԮݢY3p�K��y�&��5�������GO�	�y��u@�� �lK�L�h	Ӷ.ͷ�yB+U)�XTX�n�A�d ��Ő�y"��g�z	!��ѩ<���[6I���y¢�zUd}���B�B-7�ޞ�yr���&3�x�iH�>�@�1S�X�yNݹ׼=ZNFE	B
)�y2�޷��p�Ư�4T��i2�Ԩ�y�D��qbG0J Ƽ�a���y�A-&��0�����:dzMKq��y
� dT�ul�Jo�1����W9rI�"O��@fۆ��P��o)O�h�YT"OPx�ژKV
�n�l Z]��"O�M�����v�����LT+����"O|!U�J2J�}j�¡�Hɠ�"O���B�P�=�r�#���'I���Cr"O�-i C�["�|���1�`��A"O��(%I��W��!�N7d���I5"O�=��j�%��D���4i*n���"OB�KU�hP�蒖N�*t�0��"O��(��)H��C�O�4=<�5�"O�}���R�L&d����_�^5h��"O�x����=�x��DNBG*�"O���`��){���b�MG).:�d"O<��R��o���4�[kb�	�"OҵjB,�#> ���e�1�ڔp�"O�<y �7a�f0�a�P�Q�6#"O�m��a�I<��C^�㎕Q�"OJ@��5>epG�f��I�"OVi�$'ۄ�.�a.��!T�dj2"O���I"�H\�c"ȹzZa	�"O8A�gIYb�C�����T"O�9����ȣ�
H�?� PD"ORа���7=�Y�����"O4��8���c'ޔA��͢P"O6XgӇ7����E�3,��p"O��Q��V�Rl�����&}L��"O�d�B��e7�4���W"�Q"O(4�W���Z���cJ�X��e��"O���'U# 7du�D
b�$1�"O�LS&ăt��7H����p�V"O����˟�8����т#�^���"O�!B���1W��׍�g��!S"O�p!/� �ģ��˥�>]�d"O���k�U��Q�3kꀅ��"O�Ba�o�i �H�9�P���"O&m�pǚ)m�tFhD!/�<�r"O�3n��6�^�	��ʆ@�$�b�"O��cH<�!�&��T�� q1"O\�"�A��L�`h�3��pcJ䒕"O~L	A��/M�\rDDF�eS���"O��S��яWW>���ߏ!F01P�"Oa$m �}��T��>eJ�"O��ie�2r��b�_"3��`"S"O�<[V��-)�h��A�T���P"O2a�HW�Y>�T/��G}J��"O�!c�� G5\���	Q|��"O�I�� VIhA3�g�cGȝ�"O�QXwe��FE��g_���"On�(�o߼<�đ)�&����"O\�cHS�h�M����|��Hb�"O6�"�f�Dr�G�:G���"O�XX���H�V���4�WU�<�"�C�w�@��B�������S�<Y�	B�lδ�!sj��%��5�$��N�<���X�p�"Nz!6,E�v,\�ȓ7�8z�,Ҽ7�<L�1gU����8��!�Q�G�(8�� Θ�gP���ȓF��l��D���¹;���@v� ��.!*m���=]^�O�$ ��ȓp465!D,�~�q�d��C���ȓHZ��Ekà>1L��'�Ʉ&�Y�ȓ,
�mzU]�: V)ɄF�8Y�ȓ:�~�%�J L*H�"�ջt\�8��S�? �q�(Ӯs�00�&B08��u"O:�b�˙�o�fP�o�y$@��"O�8Q�$� N�^r���t�p�"OV�:�#�De8y:2�� Ӧ0�"O�R��^���Z��P�3(~�@t"O�@��j�,C]$02%���v�Т"O����*�N>ȡ&��0
��*�"O@4��I�#�P=:w�0WX$q�"O氢Co߫]~�!w�Q�,k�<q`"O��0��ڲ�V-�gF��-p�AK�"O����"3Ӑ���J�C��*'"O*eS �հ}��!��k�_���"O���gGIb8^���Şl,�1�"O�4�;x9�S�	*DG�y�E"Op���Ĭ[�~4��H�I,����"O�P�AgnM�y���
 ޥ��"O����
d�R�y6���<e����"O���F�)�*�-��Ċ�"O�����3�� [�ˉ�.5�\��"O�S���NX�,H�08X�"Ofh�G���#S�7 ���p&"ObyB�'P?\�:�Ͼ=�d�õ"O(��$N� �R�KC��l��"Ox�2 ̃�U�B�1�R�!W*�0E"Oz\�5�өX��9z�%�0"�]"O���W�]�m-�d��
��֗K�<�THG�`Zt�x�b�)$�H��J�K�<!���3hr:Ek��Ȑ5Q��Z3!ES�<�����i�Φ7L|�[�D�Z�<A�a����`쟣���Oq�<Dj\>$�D�Z	.���p#
n�<��=J��8��.�Da�u�m�<YQe�D��h��:u3��׀�N�<��X�A��]���1@�V`��
K�<aVCćɀ��Tk�j��d�P�<Ic��0VHLp�@+RBX��I�<q"�S�M��8�h�`��0K�	W[�<��g÷x�Q�4��S<5�`M
s�<i$�p3jq� �M�ư�{�n�<!�DނB��G�
6ly��(@�Ql�<�pLA�fv I��P3[�H�Y!B`�<��$ D"��*FL�dƸ	���A�<	g��9�p��IŪe���DD_T�<�R� �:�rAZ���X�$	
�i�<y � *���� ��"���3��}�<�gnŐ1�Ҩ@ Ӄ`>�(�AmT{�<��\&7��̸p�R>g��e��j�u�<) 	�.z��Y�M7�"QJ�K�l�<)� �7���W��4Vm8d��$�c�<��L�x�h�C�D>8�T�qN�i�<�(ڻ0�=C"�l,����b�<�!IY��z܂!��*�X��kH�<	��A��lr�҆dv�)KS	�C�<F��\�rx��G�oL(�*R�W|�<�Ӭ�/z�͑2LY�4�b�H�m�<�L�7Inp�A�ҩa���T�Ij�<�q���;��adB/4�<�1�j�<IVA��=�����S�`�XP,�e�<a�E��	DQ�c��#kRP 3M^�<�U�,:�a�:���Db^�<�&]�M0 �(�aK�&�����X�<ip/�:�lt�%,�j�D��3FK�<s����,�跀V�P�����mC�<!�B�3V�J�!�aޗ�,(���<� �-QB�;y,:8	���P�Y�"OP	��J)W��+�D
b��ݓ�"O�<3f$M�o�R9��DY�!��u"�"O�l�!CH|�5I�A�.�ph#5"O��Z���%߾|Q��[����"O���M�u�!{�^�[(�j�"OXȕ Q:T�`��ćV'J�3�"Ob�4"�;D�����x����g"O���r��L��e��9KZ�B�"O�X
6I����Ǫ�2m$Ҡ�a"O�e��ɏKcv�!�_<� Bg"O�e�P$E�&|��B2c����r"O�
m�(�`�rw�+� *�"O�}z%Ȉ!h~|�s�-n�;�"O�\����Ri�T+�ZK ��c"O �9WMԏBH���߇VW��2"O��)we���8J��SO6� #"O� �*߈��}K�	��pԐ䡡"O�iȕi�
wBa��	��r!"O���S�y����� H�6Y��"O1��Kc�E��/)SThr"O��$J�bt���OB!*�V���"O ����0 w��#��߼0��0�f"O�����V�$�����X�#�"O�����8="�Ϟb͐<Ð"O���%f4xp�\����UQ"OH40���
+�8:1��W�<0�"ObTK$��7��'��)7���"O�`�b�4T0Ѻ%�	fcxE�"O�ܹ`LG��s	�@N8ܹ5"OX�2)�c� H� R6	��"O2���,�,(�TD���˃@|�B�"Ox�*�#�H�t��J� ޕ��"OLX�)U�J��;3#qH���"Od�9A�7H>�C����2���"Od���	ǬP��b�'�?Ђp)�"O�u����>.��D9d	�(���c"O��mS�wV�|�'I��a���	�"O8�	vM�F�Yj�g��m$��@ "O
 �'��^��$	�&rs�bu"O����F| �CeR$ k�y��"Ot�ۥK̓SFʩ�a&��je��"ObH�e�B1
Dy�Fקfh��a�"O.�FK�bw����ʑ7t i�"OP�����`��3�c�c��i��"O�{�C��1!��g�-��
�"O���O��4�#���T���"O��Ԁ܇(�*�AV%� ;��y�"O��aR���`�4%�G�~���"O2�1�蔓#X�48���<���u"O�Q��n�%.�	�ֳ9[���à-D����ܲ:|��+�5�X�cA�*D�� E�)F^d���_FtK%�(D�l�E)�4?>�ٓ표=�*T�e$D��tE�!s�ʐ{c���]���� D���䨜uP����4A��u��>D�v�H�dl�()�nb/�w�<)�h	K�5��h�M���ذk�q�<!�'�|�Y�i����%�&�m�<!p���"����l^�9�FMh�<Q��Z&�< R�kӖaMrp�z�<�I����a�bU��d��P�<i��� :ev z�#�2qA$i�S�<���.I�l�(�Ft������d�<� �\s��٤����H�<R��3"O���jP�'����$��=N*��"O���b�� B�hS��BN���"O�0�`ӠDf>I�� �

Mt�Qg"O��c�K�b��H0�@a:��0@"O���`,R	S	��@��"O��(��ŉOI�P��\�0<bE"O�� �U�}ؕ�rgD̸�"O�4	�"
�;k,�q�2o��"O�¢kE	Y��(*��ʃO�e�"O*�"΢2�HD���+4X� 4"OB��tOD;6< EkD��)pt��a"O|Z���++�K�l\q�^�� "Oh,�C�&$t����%!zޑ8�"O�|�ӢH(T�� y���vv��"OR)�g�R��B�����uqJ@�"O@@v�P�Mɾ� t ݆)bx ��"O�����!\
�H�SmK'yL��pe"OP�14�؄�~b�+CA�$JC"O&$ �#Kf;P�%NM"����"O��PM�??��RD\We.���"O8�C(O�J��P�"\ I<0"O�	˓ ءC�z!�%g\Ya��K�"O��$d
$�ڭ��.iK��[�"OY1l�0u�T<X�j��LTBA��"OFU2�Š��
�IX�0IV��&"O����T����	_���"O9�Eӂ�j4#���4$R�}��"O�%�qb�n����$�K�})�Q�r"Oj����C�jKΕp��("O�M`��?�����g`����"O��"��,3��X�Bf�.-m�@ 3"O>���]�M��LZ0e�ǲ�1"O��&'!e�m �mB��D!P"OPx�b�^�;���Rg.����u"O~T�N�:P�J���n�_��	��"OLH�o���`@��O��P�36"OP���2$���zT��%mP���"O�i�����oG��iWg��.M�1"Oظz���2c�Aڕ�4A"�q��"OhUy�jK:C3|@	�U�W2�X�"O~�y��Ǜm?\e�%�V"F��	sV"O
�� ��>Da�Ak�̚#ߜݺ�"O�c�/^4\I6x��f��`¶u�"Oh�i��[�*�:��N(G�R�3"O�:Ӌ@�N�t�C�M'g�l�8B"O�+�(ҋ~�&pj��E�g)�Ds�"O��ZEB(�9J%�V����'"O�׌G���5�-űl�����"O��y3�+H�ZGH�N�2<J�"O�[c�=q.��s��?�]y�"O8�*�e�h;��,ڎ�C"O�1�ȿ'ń�����L�`��"O��˅���=�3K�E�J�2�"O\�螳6@��X�J_���R"O��f�	-��qh�	�q� d"O�����a�)���E�yYV"O�)���'NJ�
c�� ����e"OJ��F��%`�|,ȓ�C4#����"O&lACH.&�ȼխ�-d0��E"Or�t��5�)9��	�4�"Op�I���|�f�풎G�)Pt"Ox	HW&�6� h��-�s�<D��"OpIr�AK�{�>���O6�H7"O� NyAW-�Hc`	��t��(1"Oh��4v��aC�	��VYH"O���3 �r`]�A�h�&�:C"O�R���&eҘ�A�W��p�1�"O���#j�;lՂ�h�h�,��"Od�R�ּv�P���0)�LZ3"Of=�/_�3@�I'h�{�T t"OVheMM��i��	X���I�"O�	���^��D�(�*��Ԣ "O�X��j�Y������ՍҀaV"O��A�aO/M���� ��Ed����"Oր��'Or����ȏ�B�~��"O$�a��B���N1g�$��"O���&��th�d03I�����"O�0�������XAH�-�^4r�"O��r�Bí�
��B�:���C�"O�:���I$ 4�g�� 5�1;�"Ot���@� +7�`���V��)�"O�j�^�H��ՠSHZ���y�"O���L��Z�
�f��"O�pӇ*��J�Ȳ�H%t�)�S"O�QWB	�>�'l[�kS"O"����ӥ=,�}	2�F�6�e��"O��@tN�Go��t�
����"O�2�7
p���C#P�`D+"OJ)sQ)�B֌�ҲI�G-F-;�"Oް0KՐ3w12B�$�I	�"OV@8�`Q-�а*""P�NR��"OաBeE�T��5G�#a�@#0"On12]�nuH`I��ʴ-ޠ8�"O.
ul����G����U�<!ၙHb*t�D�����rD�k�<y�r�c(
%��9�/�L�<�Q��=@^,�ą�x<�A�CF�<���_�guc�`׿s��)���Z�<7���=͌t��n\;U��=�#�Qm�<9&�TsX���gʹ>��!G�g�<As��'Fz9`���.|8���c�<��`�{C����]�B>���f�z�<y3̟�^<��w�؃�<e`�O�a�<�ǨU.<\�B�H`(�_�<C]S�
ي�,��[�B�x��Iu�<�2	9p�| �	�8(:�1(�E�[�<ɣk�8�� ه"4fJ@PץDA�<���S=2���늪&�\Y"A�<Q�(@. �i�åZ% J�`:��My�<9q��D��mџoA&��b�z�<g�Ϊ'c��c!��5�����}�<a�Ə�+�z�&��(��gx�<A'�_<]�̄�����h�� ��L�<��A8%[j�H�K�CJС� ��J�<�b�R�)��9p��./�b"D�<�S	ć~@��j&���,��E,�A�<�eI��^7/�4[EX�2�ѷ�y����]S�A��&Ԡ)�')a����ά�� �<y�$!�cO�k���ȓ,����T � ��F�V���G$�(�aH�d�zq�����ȓR:�y�c@�F�������U U�ȓ0_��(E�y^Pz�ȅ��Z�ȓh4f��!N��fۢ�ʠB��w����7�<]��@�wTj�ar�Y��L��ȓLn���ֆP�"ձ�a^7B�6̆ȓ!��9H aJ;�):��G�v���S�? �	�4y�@���-�`[�"OH��EMѫ"̞x���_�B.Q1�"O��h�G�#y��5Bq���M;0��"O�9�tD#�>A��K��t�n$٠"OZl��ѭe+��	T�*��|8�"O��H���/E�|�`��
�l�ҩ�"O��ʒ�xz��qМ;R��"O-ip)��7���d-�� ��(��"O�:�"ֶr�<�%.A61�"O�� .\0~�S�@�:����"O�(� ŀ�)Q�A�/r�~ɳ�"On���aS��#��	��"Ol�����6�����I�K�F�if"O�xI!l]�:3~y��$Z�j�y3g"O搋�h�Pd�A�4Dϻ?t��X2"O�$��ь��(C0Ă�	g�4 "O.�5��9 Y9�l%[�`˂"O�EqT@�)	���k>O>
]��"O���������!Ҝ<L�}1"O��&HѾ&:�R�(Ä~��I�"OTI�@EW��r�9���%U��,( "O�1R`	��tfm�u�1��}��"OpU#��'vv.h�V�P�{�
1��"Of������sd�5�7��-���1�"O���&e� $�&���)z�x�80"OP�B��(\�Ua��¢�<�)�"On�5����$��@��:T���"O.8#���9/�����~�P��&"OfH��M��[␠�"DY�<R�"O氛�T�v�RY�B� fE&�Zd"O��J�1c�m���1 �A�"O�p��T�~�,�Q���.l�8�"O������ ��W�8�6"O
��Q��+�`Q�An���{�"OFX�U��(ܒ�S�셿M���P"O�d1/^T�JA����'^��B�"OJ9�"߃l*̐K�8
y���"OҬ� ��ʭz��x~�S%"O�}���6:@N�[�dӰbp�աC"O�H �%�
p`1�2㎞XI��`"O ���jU�#,v�V�)>����&"O�P�F�5U.�H� U�Zڄ��"O��r�G	?���.�9A�*���"O��ѵ�U";���C��@-Ҕ`�"O�*KK;�Z�
�Չq$Z}�d"O�-��� t!�(���	���83"O
1"$B��k�ԴHoW� �dX(a"OVHҧB�!�b�J��5c�H�Ұ"O�Ds"�uk&���k�!�5q�"Ov�����	u#�+֪ w�.��D"O��5o]/@�V�
�ȑy�|�@�"O.=S� ?y�-;�MK�ú)!B"O�e3`��2{Ll�.јO!�<��"O�A��nhv�;R�!g�@ң"O�46c�+-�v�I�����4�2"O���k�,��er�kϾW�0��"O֥�c)\PhA��%��@"O<XG¡ *�A�.ؚo	V�#�"OȐ���}�"tb��=1��q�P"OD�[�)�8�}�$��K��a�R"O,��`9d#X�i��]|��"O`�r�	ˬd�D��@h��hWP��#"O��#Q��sy��i�Y?j@��rR"Oژ�M��i�$��S%P:w1�|��"O� �;�'ڡC�� G� U� @�U"O���)�����1�[8VP�"O� �"S'TQ�8p��[�S%,���"O~Q�F�P_@���y�5[�"O��2��g*al�+�z�#"O�%C��-m�����,+��"O���Ĵ
� E��L*<�(��"Ol�؅NIq��i�I� ��\"O����#�t2�����7gɆ5Y�*O4��`�.a{F����4Z���H�'�`�K�˛rJS,�J�hS�'��qD�ٖ&:7G�;�*3�'�tP ��4�0��W �)/����'\�=1�R�Fy����M��*�DB	�'��9w�-#�.`��K[�X$�=0	�'���ɗ�Q�%O(��Xy�'ج��A�åt�<�IS��p�8 �'�֜��X%p�L�r�j�(EҴ�p�'�t�i���~��u�a#��K�:�'I�H0L�7o���l0-q���' |@إ�&o���0���*[�qh�'|��ċZ�HzfI�+�'��y�'�촛c��'Qi Q5��/>�l��'�l�w�[+0�h{w����4�	�'4"�s�/Ǆ
�!��α����	�'�2�N�3rj�XQ�.��ce� K	�'jx�#��_!{�`��Ȃ.Yk��2	�'�&�IUa�:O���$'�2M�ޕ	�'��A��͇)�,ЈCD�B9�T��'Rn���%H��`���4,
�*�'� ��hΣ7mj	ғ rjp�'� �v�̨u��l����b�@��	�'�%IC�bS��U�̂l�J���'@Lt��_����${�p�EϚJ�<y�p�9��L���� �
�E�<a6�Ţ)������B;�Z�A�Z�<QeQ��a�'S����00,�}�<����?a"9�D�O�pgXQ�th�T�<�0���mB�g�����Oe�<�Dn˯U��i���;bS�5���J�<	��Kzư+A.�7R�����I�<��̅76FU��$G0U��Ȕm�F�<ٲ��<��`eY�B*�U7� l�<�.C!	�0*��U=nZ�k ��f�<i���>�N��u�B�<Kh+�h�n�<��B\�Z^0!
J8=��1���j�<���J6����Ұ8n���DNf�<�o�#5�`����0d]�@
�|�<i �5�Ai��J+6d��1���p�<��J
V4@�XVaD�H�\��q�<r�O;4��`�&X}�ы�%�W�<	4�A�kY�d���"4}�h�	RY�<��ȑ4/φ��%�_�n�,1��\@�<!���&	Ђi3@����Pi�d�w�<��I�/Y��Ks���|ml�G��C䉿ov����<R[8�R�fМ�B䉁_y���f�&n6D"�NΨw1C�I5.!9��7��k��Np�B�I�HR�90#E4j���"�ѧp@JC䉧
�.l��ɬh^03���h�:C䉀 `H�1�R�F���)ąL�[�C�5,p4�`��]�>��C�ꔵ �C�ɡ)�pU��jLF$����=ri(B�������h	:���BU�c��C�)� PT��P�#b��xu͕�!�y�Q"Ox��醔5���j�+�=;��� "O.U�j���H�D�S�!-�]��"O\���b��B{�E��i1$.�"O~XHw��6}�*�9�I�9/�n���"OD�i�"<1
�Z��\%x��J"O�P�FE7e�"�����"O4���GzH1#�l��r� �"O�H���Vt.��*��?�e�"Ox���čL�29�&ہ"�f ��"O��s!nL4ߤ���N������"O���dˁ�c�x]���U���0�"Ox%J��ư4��]���8�`��2"O�ћ �Z�H��4	�-*�d̒'"O@y�Щ�4���+��B�"O�tx �A�*`(�t��6F��|C"OZ����B�"d�:X�$��;�"O��Q�t��YS�G+>�J���"O���u���O�@ 󦗶����7"OЭ��KAC�L�3�4vptܺD"OB1��䏎.,�AtB�zaH���"O�D�E�ߵ8f�"���,[�h "O�u�c�'T�|��`ǝR�Hr�"Op��@�>W�JH�1J�Y!��I�"O���LѣD�%A���l��q"Od!��GZ�Gt�!�F��:1kw"O\tq���=~J.�$�0P�����')�����D�"2�.p�v��'����̠!�F��"]�0���'">�0���#f�KqF��
P�Pb�<�c��#�>���گ':�I2]�<q�kݼ�$�pb�3�P��h�_�<�Ei_�9�1	�ˑ%u��8��,Pe�<u��,v��vj�%l�B�h�dGb�<�$m�G��\���@���"KSa�<�g��>�k���'�� �u�3T����oR�4�����;EY�c�+D�<`�i[#�p<%�5~��}�C`+D�t�&E�)~�� [Ἃ�d�x�*
�'N�T�6�-��Yy�@J�35�e�
�'���P�[�2T��;� .jR,p	�'�(3�P�C�|�gV)$�Lu��'F���5��L��x�*I�"1b1R�'�ʤ�t-��^��x	��3�`�S�'���J���Ga:Dѣʞ|���'?^�Q׊
�e���	�{V���'ƴ��᝺
�Zq�T a%��'�ix�E\�^4��B$qڙ��'��l�Gʅ�JW��a"C���bH	�'�ҹ�� �2ɤ�C�J�9	=�H*�'��ə^3}����3k^�.ZЉ
�'^\��� /�2� #�]
���	�'�R��`j�}�Pi1e,�Nݒ�z	�'����"�"h!&��t�θA)�L�ʓ+�8�q·�H�����V��ȓW|���R�I�YE��@�%�Td `��@k�$r�j�&r�88��\�U����i���k��t���IQ.L�cD���O`��w��AJji*2d�0d����'�O�(�@��:���G>�l1��"Od����taB/�.$.KB�Ƀ�!�ē >��p'�l��	�g�+<�!��S$n�|mI�$�T2����?�ax"�	d����C�D�,Y����@�C�)� lB!�N2��a���=($���"O4LҔ�խR�4�Z��tRd�'���Ƃ�b�24��{߬L��� fp!��݉:QQ����`è���/ȲQ�~�[��Y�H�&�\\�Δ�&1���&D�$��@Їm�%Ӏ���&~��"%D���ۦ}CHу���1�p��F�0D���=M܊Hg@�:BY$�)D�0Q�b�:*���q$@X?`N���n"D��BCطrW^�
D�Ʉ���!D�8�ȃ�GfH	�T#g+$��B4D��3�d��\~)rv�D�# P{��1D���w'�45��q+�+�L�Rv�+D��(A]%2т�ⓌH�fg"�(D���dI���1ț� �\��ӭ&D�$��(
+�в�I�H[L���/D�,qӨ��7�� �gy�܁x&�.D�0Çf�5=�ZrGU�`G�E��+D���@��p,LI��Q:h�x�w�%D��ǉָD��3m��9�X�ڷ
"D�h���U.\2L�Zr&�(� �?D�L���<	��ʂ���_�P{c�*D��`�N�ࢥ`�2{��J��%D�����IcBt+1%�	WR�� !&D�����ɚ0Pt��`�%S�jxq�#�O��/_T��F�Z(��mۊ
P�t��3 �b�TN!x<�F|��S=*��2F.�"lr��	7쌥rstC䉻 �F��ѧ9��bA�#OlC�I�
�Ap �0\��j @�+*tB�I�}�H@��ȫ8"��o��'�B�I� ����K�<M�EJ0���Q�0��$b��؃iF�F�+��\A]F���C,D��)�Ie���z�@��`E�)���yb����xG)F�6͊x9�Ƌ�p4!�Dˬ)�Z����ԝ^ �+�RV(�'J�"=�}�0��a`�"#��a ��P��l�<Ys��([��p�҄@��C�q��0=92K���N��gǌ'8���q�kf�<ɤ��2����a� Bv��ĮR�L�!��!6�����#�����*L��z���ǲG� �p@��5��H���ިQ��}R�����M�@�Dp���OM`���C�4�q���"�"���/�6�UC�$�<�V8�ȓ+���Vh@<�r��섕dd�ȓ+��q5Kݑ{o>�z�Nh�.a��?1,O@�Sܧ��X(��K�AV�����b��H<!�$�zYy�ˌp�����:!�d���e;$���C�ED�"!�Ď]¹�U��/��eXR$�>�1OB��$��[���kqC�-W�1f��!��R�|@d[E���IYl�P���|���
O"li�I!)��!���M[���`��]����[1)���+�푝gä���$Y!򤆃e@N���F2[�&؂u��y2�	~��L���X�j1��seS�Z�L��Cc(�O��'��d�To�</K>�#���&u�)��'�!�)ڧ3�y�%Νtq�`��nf�&$��ROƝ�3c��Bh<��5<U����X�8�r�c��5=.�hnZf̓���s�@8j�CW�d��R�LC�y�@}A��'_�ɳ��5�r��}�Nd�P�W�	�����Nax"��W0�x(W�����hd�A��'�d̿���V�)FL�\�D�Cط�}	�"O� ȵ���l���skD�GjH����	L�D?��)E��cԒU��HM�](B�ɵcA���1q�X� ��L4#,c��뉮M��U��R2v�8�9�(˽!��B�	*ZS����k�&7E�㣌�4C�ɘg}h]iU���,A #�}�ڢ?����F� �E��L�3��ȡo�1a!��܃#G�aC#`�6�6\ÐB!��L {��y�D�F% �T ��%�,�D#�Ox���ݒ�EF�(^4-�B�'K�'p����z����K�6"��Q��'͞��TGHR�85gߋ	:�-(�'2�� D?G֜�j4��xA�D��'q~D"t�W�m��́��\�88�	b�,�#��P0�X˶��[�ĽhD�9D��c��C�Cm�}* %�d/b!�A9D�`a���|�(��ȗ�0�6D��b���ȪԭE5�U�'�'D��rCΉ�z���R�j�?.�!��&D���AŘ�b馩��O��؛g�$��ȟ�����^.r�h�@�K_��k�0O�=	���*�^3�ػ\�\ᥤɡ:�!�L�$��t���@���  �Z�!�$�:>��xh�l�L�0=z�B-h�!�d�f�vi:�"�%�~��7��%R�!��I� T�U�Ã�^��8��lѡ!!�D(nud��F!L&R�]+. /!�d��i��ݪ�"ӻU�ڨxǃ��H	��D�� ����W�R�b�G���j��1@3�	P���OF|��CW�3X�����\�<p��'����C��0x3��ѷxߔ���'���F9��m`F@�Z �'�>�H�NĿ@a$�0�	;` t��'��51��4j�����/0$J��D2��"��s�>ld@hX�&?U$�\���v�`��(����gGE���ȓDx@�(`ڜaR�L�2��S�v��ȓgZnU�dF�S��L{Q"�j&n���|>��1�"�lJ��T�(�مȓW2��F�pj��!��(N��ExR��(��'5x:q�r�C�{��UkRF1L�%����	ң��>�&Qsd?M�^�����k��ħ�pwΐ4��1���vJ.��'dqO���!�'�FD�-G��yY��
�q�	���p���$R�g��	�Qc�%yZ�/[����M<!���~��'B T��o�+	��[R���$�\<���x�M�#9�`�%�]�T;��+�'�#�y���8'[�)��5uv�}�4��/�y���K���ے�w/������(Of�=�Oz�I�*̸Y��9�"�) S��
�'(|�3(�u�v���"~��m ���ꦣ|�'�ԅ���{x��3�2�Y	�'atY�'^!S}���^v�����4I�<�����(҂��W$����Z9R�c� Dy�A����2�Z� ��W.*��_W�ި�ȓ$4jаԢE% �t��4
�,H2�0�'"�zx��C%b�5��T���J�C^����:�O���&g
����`��8��1��4Z�����>Iү�	16�#SdP '�m��MU�'cQ�,�O�� �����|�bhbL�
�'�܀i�L�5Y�d�`Ι�T��@�	�'��I˦��IA�����^�!�J!�'��P��Ń��4�!leI��d�<��Z8p�~4+��	`ה���Aj�<� 8!B�w<�K���l�`��"O&��u����� ��$[��t8"O��pC#�8MF0��  9�L���"Ó���&zU�`�j�V� � "O�9����qZ�����(IhF"O�T����z0Y��N�C�Ɣ�"O��c�Ñ`kLP��T�L�%"O���F(�2R�<Q�s�݄.����b"O��k�Ś�v%�x��C����"O>�`R�W�PfV��тU�w�l� �"OyQ�i�,_H"�೧��|X�cR"OZ9��oͼ[��Y��Q5`���"O-�ʞJ	� afA _D�lYE"O|ar�Q#�0�c@Ǘy%�l�B"O����/N��Ĝbu�!ʝ��"O������%Tp9��Ɠ�s� Ű�"O��"�l�{�
����Y�b���"O��e��3O�w��+A����g"O���%���BzA8�ů�pDh "O���ah�t-+��C�[���
"O� ��T�Hu���0H��:�"O�|�&��p����g�ť+�\��w"O\�0���q�@�h!��Б�5"O�q��(�'!^���`��Xc�e`�"O�9�.�5v촁�A�ݓrP��R"O�`�Kũ	J05�-�036�*�"Or$�1�Q�k�i��L�E!"O0��- 1rP~Ia*�	����"OP;���p�F�?d�f�8�I�m��l��N$Q.M�w��托2*���v�M=[J��tO��d�C�9rV��P�$�������5(�NB�I~�愳�bS��Na���<Y_�C�I�F&9`4�'�N��h�FQ^C�	��D��	�qbl�u�M�ZF C�I�x��3�aUq�䣡,�:Q%C�Ɏ*Jduss�_(e{��0�>k7ZC�	�o���ѥZ�[�v�� IC���B�Ito��;ǬH�)u�-�S��
a�B�	;=AL�[�;Q9�e�!��L/�B䉏k?�|N�z�b]8*�sV�B䉯�0@(�$\�+p�p	��	�nB�I.��<�@�ya��"[ᦨ�P�.D��k�
A(LH�0z��9]��,�a�/D���C~��y0�	V%2���;D���])At����g0���=D��"W�܅>�qx��#z4���u�.D�0"B���� �C�N�bp�K�.D����j�)D�"P(��
�68ح���-D���	4�D 9a�E�-���*D��c��Ab�a��Ó$��6=D�$� ��N:؅��_��,HB��8D�8����$��5*'\ s�
@b��6D���H+5%��ز��!�&4D� Ⓜ�M��]�U�עa��I��5D�t)�(�0`�|��Sn��W2�ɋ\~!�C=����',��P�C��vw!��ֆR��]�E�-HepZv
�j!�$N�NF���/V�����7?B!�̜���*�E�gZ�D{7lǃ2%!��U2%�衚2IHo�i�˕��!�U 7�$��S��>W9��0��@�p�!����X�2��߰8hX�Eo��g�!�$ �?���W�I �)6͈�^%!��	����&�:P�����ѻu!�� N8�UH�-<;�uj$��+�:�#"O�=F)��`�X�:�|��%"Oι�u��0U��u��'Z�vQq"O<�u�ި{��d��oF3V���AV"O|ipD�$M�X	#��P�Tԁ�"O�q����[5+3e�;}��)��"O�H�"��T�.���Ū��	+�"O���$C�8���0g�Q�����S"O<��`��#�)�c�۹��Uxs"O��cG�Q�SR��z�J��
�<б�"O�A%�J�e�bt�Eo��Ba"Op�S�E�T��M��[�F�h�"Oz 	�B�E
�л�l˓��{"O�)�p�8$�lpg�A|��(p�"O�H�.�# ���E�O2(u�@I"O��mN,��D��Z<Uy���W"O�)�G�ْ3l��3 G����"OR�b��_
5"l�Q�ŕ�G�LT{w"Oj	)����Ԩ�W�׼��ie"OԐ�a G�(�Y��F�e"��"O\�+4��"ٜ�b��dU�H7"O�8�� ��wR ;�bN)��Y�"O5Y3�W&3�P��@��#�D岤"O0ݲ�*�6?6�u1�5SF�xZ�"O�])���2�ѫ����%T!�G"O����B��̗�(�R"O���)�V4j�pK��k��! �"O|�)���6d����
���!�dFs�f�#�k��}���K4h�!�$֍^M9��j��[k�)I��@<�!��C({3��[�l��zV��%�Zz�!�P#D@Pb��xd4TB���'q!��$PW�%#��J�x���B�pl!��.D֊5�Q�V�Em�1����]%!����@
Rn���=�D��+2�!�$�I�� �
ȨvN+��LIJ!�D(<�� �����n	h���I��0!�d����a$�
P�+&[�'j�t��WXb%3C+^;����vLܼ4�D�ȓfm @�+)QL��˥K��/gZA��F|69� �9H��TB��m�J�Ey���G~21�1`�9I��t�z��M�.�J8�T�1o�~�;����y2�{�#@�N�`���Br^!����� ъ��d`�\�q9$�s���riKjM�Y�I"�j�(p!��`|��	6��*Q�����ur��:��]�c$Őb�J�h�XaW�O}��EzBm@�?�:���$M��d)�ê��=�)L�'�$���-A�<DTA�%�5HO�cqeWbk^%#�DP6|��d>�O�1b��� �v˵ I�%�b�����_h��d���6� �FA��ҭ�ƤY�	+)��(�%�@����"O\8�g+Z�`�X��#!�� ��zQkE��UY�hT�:�Y��J��V0����v���T��Ԝ���F�HN ��T�>D���F�z�LH�GhC-o�����^6cn!��k��y�.�FM�s���	��y�T"<�v���(�PR'G�	iL�DPu��,��ƕH�}�֮�"��]"À�.?����E䈸Y�2�	��\'7�Ų͍~��e,�<DLc4U�B�p�+�	�cBequ
��w*t�����7���x�A�|�0kC�Tӄ	i���-C�����TM�<Y�E07�p�9b�"'�
 1`g�E�V[3��!#�)z��zh-	tM�p��yWfG~��C�%ފ���6��y"� y�"�WH���2�.s��(�g( �6�nS;���o��O��s�*d;Z ����r�P�u�'6��a�h�(����$�e[ׂ����Ppޒ3�ЉP��Z�p'���k;�O��9�#�!�r����O#И�K����i�������L�ٴ#��x���ު��f��GG��@'��6
`�B�U�y2J̬Z�������2�\��
I$��Ԛ��;R��	���=o��\Jq
�l�$�X�=� �i�Q��W��9��6 �U��"O,��6��&U���b�5gSI ��l�vt��E+�bH[ve� 0.��v-g�'..tQ2"���v��ӎѤHo��a�v8f�Y�h�2��0a˓>d�Dq-� ����C�K쐰�s&.��Y�l��^n&Y0�����m,���<��-�@Ǣ-���Ҥ �jb>i�d�@%<��bH�[�Z�I� )D��Z�YJ�ܸ'b�R3:���D�{s���e$J*:T	�S�dB�?q�'|0˦%R�{������C͊���'�Ƚ�c��<�`a�t��Ve��`5�܊=�L��C���L{�u %�Wax��7(+�|��H��nӒ̹�����<����mۆ����~QlQ�2f�i�.���#��^�n�+���"f<��'�d@�P�8q�V���H�,Ұ�I>�$Ɯ���G��h�+���јOo
90톂W&Ф�tF�"�x%��'�P���B��(�n��0LZ�/D�y2�yT,��;�Δ:0Á���O�ɏj��p�A���D� @��@(B��Ir����]��q�ۗs����M���@a�c&�e!�:Is���=��G}>eȶ�L�?����L3Zr�bW�)LO��) f� )0p��b$��v`�=�70C&���:;`��Ý�{���D"����(��d�_���K�,;f�|TJ�Õ 1O~\R�c���uo\<&�D�k����X�4't�5m~H��P���?AS���BP@�Ƨ4lO�����;�����= ��B�j�# ��Xhu��:)`�O^fi�c@8-f��mZ�%].QKX�h�+�JDpS"O$ ���L��v�z��Z$f�Na9r
,L���χ,U>�Uz6��&�<���~�$P�,GLIH��ɖ'�D�rJ�.e��TR�^
�����]�,P
��,L����.ٛw���"`��
-�0�d�\鄅!�n��b$�0��!k��\�X�b����@V�����T�g.����/�>�����A�-2r7��6Q\��������!S�H��@ɪV�h�p�ѕ�?!Emt	b`$�*z�a{�,�]��I�
�9�I'k���M��; HV�ɸ#�tc�J��S�疌��]fk,�	�䄈��ӞFm�,�e��_!�z�����R�-H���!���1���剣/�6��r���)�O�:�ϻyvPQ���-�<@����
�\��4
�H4M�)&C1 >F�,=K#��
C�"���Aq~� ���Ux����_��m���ߞS*L�5�Z��z�GTV�b��榄�<!6�g����CM���G��Y?�7nP������tOF���kJ�l��H�u��oDqO �
�5'�дk���@�1���R`�-w�\ ��I�f�!��G�c���Bb!(�5¡���q�rh 6)L,U!�Y�2�|�'Jlb �#c��0�Q=9�v<"�'X�����J�V���p3n��x�.0��42}ZI���p>����2�r�T)A<��phF��Pу ���	�D9�e�ӊG�f�ca*�{��C��;+��Ps`�� /,��`CmM3��C䉉W�(YP/G9#�[ԩѕS`fC��(p�l �f��*t�%P&7�@C�I�"�,��%�Z�&��G*N5H4�B�I��L�1$D��&�k��O�)]�C�I�a<t����ؿ}��@��l��C�ɀM-:�
�D��0ZT����T�|�C�I;cz�;S���j��չ�kP�K\�C�ɚ7lL�Ѳ#�>:ŬUSgLQ2F�pC�I�h�
���^--���ӐD� F�Pe��xj��"~���E_�t��f��T�n�b`'�5�.C�I�$�8�$�f���Ga��ɳL�d�HA���㲮Q�d�w��6��s3G1|O.�iC��4u��ڴU�d����' 4��� ��ȓ@�.����)a+X��!�'l��?�ā;��}ȓk&ҧq�R(��%!D���kQ^��T�ȓF䔰�$��
j��	A�)ƣ)޴C4LN걈֚>y���O�\���C�:Ö�z1)QAJB�"O�Yz��(Z"1�"�� !2�����'���`��/�p���'�\��҉
	h�>99�H�)g�V������6��&�M���F/K� ؙ�\�?e@�;7��e�<1m�: ���c(��b�=�QJ�a��&3F�b�l�vD�#}ڂk܆-Z����X�)�x�(P	X�<� r�[�'5]W�K@@S-���e��f{�L�%%@z�*�g?Y'Cf�������M��-"���y�<�j�-+
��ZW��E"4��̑�<���.w f�S�|��� �]�X�u�Ĝ�p`f���IrdƉ��2O�% m��~Wƅ 0	�!1����"O�-�c�B/�����_�?/���q"O�tQӫ
)�R�
�&�2W��ض"O-w	�1�~$�6�Z&gr��"O�x�����TOL<bQ�K}�5��"O�}I/�0BP!�!)60�(���"O�-R�k�&������ybv�QQ"O\i;c��>�H���?N�m�0"O|�:����Yn�AzQH�318��s"O>X�hJ�`�6�rF�W5d��}�a"O��BC�!*��p
K�V ���"O������q��� `���J�%��"O"�#&D
�V��q��)�d"O�D�����6ى�iX8ǔ\˖"O�A�&k�%|A���$T@T��"O≺�	�InuJ�'�2>ﮁ��"O�A㎨Z����,�f���E"O&����G�
tu�̘#C��u"O��Tl=� a3#���#���z�"O*��f�Йn�0P5�U�6̰�"OJ5�B�.JFQ�d�!2�����"O���"fJ�<��dP��j�q�"O�3�K��,����d��`7@4�q"O@��tn�;������Wb4x�8"O\�nܴ+�A�`�?��0 "O�B"ԫq8݊��E��w"O�|K@ʞFH�JW�ɟq`�|�w"O��J�t�~Y��OU&s��Y�"O|y���ͻ]�$��1Ĝ�f�e�"Oz8��.�Q��m�`	��
�,�� "O��9�_K����Ɗ!k�R)�u"O�����(�-�w'�?6�܃�"O��zGN�0y�6�*a��T`ȓ"O�IiU�\�)��U���]�u���ȇ"O~5B �Y=2�I�2/S���a�"O�0�4��[&� "��-ɲq�	�'�:a��Ŝ�^�t����� I��)��'e�(x��)eג�i���>d[�'x|0�A�P�G� |;�A]0T<�!�',��HU`
R��TH��I�` Q3�'~�U"��FR+V�	F�Ib�����'� ss��qgx����9@�.�'!2��F�ɑA���yB	W�=1��'�*A�v��z�f4�Ɖ���i��'�V��djWj�DI�bІ��(�
�'~ТEM̷0�6
�}��,
�'���1��*�Y��t�f);
�'b��ɐL�-�V�:!L,z=��?D��S�˼�Pj���p,�y*��&D��@��:)���''�i���&D��J��zxeA�\2�
�r�F>D�L�bƑ7g%>��]2�I�@�>D�����L�a6��	��Р�3D�T"��X����5f[O�ބ��.D�,��;*8\i�C�n}9�/D��ۑD�?'i�L��T�d�vm��
,D��P�H�R�:	���X�Zme�,D���'Ƥv <�@'�o�&u���&D��X�iǵg[㫏��%�EV !��B1�p�p%��y[� )E�&�!�� �Q�A�:D�r(9�.`�}�"O:9(ĝ�@�HI:�")l�P�"O~Y�c�� � [2�DB�L�@"O�	���II~����=>d���"O�8��{�Z��an�7�U�0"O^dAeΝk> H�"b��;�����"O�y��t�!hc�U[���a�"O�*vl����U�?����"O�������u0`�H03�V�;�"O��9�D�ViF�pkjԻ�"O,H9��U�2�νjgb_{ar��"O=*W�ÈZ�H�ȇO]pؽA�"O�Y�Ё�q� C�dD�hܚ�D"O05�!��<:�z���[�8.��"O��{͍�"�%(R�dU�C"O��J���N��U��HW�b��m��"ON$*Ć&~�M8�\�C��{"O�mKsK�@ф���,�%o���%"O:�1$ˇ� a���@J|0@"O�t�vlT7M��AăV�#6�cQ"O����ڱZi~�A��p�"OԹ12�R�vJ�������0�5"OD���S�-9^iҢ M{�:��"O�DH`�.wԮ�e�����A"O��z��̑��X�5�7�*A�"O"�;#��2Zt(T�/\�z��tX'"Oc���35V�8��@7c�t�+T"O��a�!�ފ$��"����"OZ�Bh���LT���_���8�f"O�<9 ��;&��ar��B"O��҄�$iJ,�p*A9�N\�"O��R$k�Ԁzv��kl��s#"Oj�4�D�A!M��舰�"OV�z5�V3c"��5�RjN`(��"Od�����lq���*]�V���"OZԺ$�� ��J!H��V�*�+R"O$0H��F���	j�G��j�L�"Ofu{D�J.Y\��B�_�0
- A"O�U�s�� ��<�R�j��U�0"O�\�g$�>6Y`u+U��<w�z!�"O���Ļ���9 ��$u��r�"O�d�S4E���d��dz�ɲe"Or��a�؇KDE�ū��:R��F"O�����zI����_��ڒ"OH�D�qf��:E�F�9�L���	�HxƜX�Qpg��*e�ƙ8��S��<��HI�z�	i�x��C�	-L]������:m��T����3t�Ҕe��[oP��ƫ	�~Ղ�cpWm��y�mQ�QL��rb�?&V�q�-���y����dD�pf����S�^�C��)�Q��`h)�!�;7|�]�'�n"=�uI�8��A�SP䢹���\��L %.��*���I�`�>T���%}W:��埫AL��)��·=��I�W�'d�i�� � ��)1��Q��ݱ��`��>ZР��E@�D9օ��ʠa�O���h%�M��Uk�v ]�
�'>��P��2�2mr���*i�p�9�c
ayHӪR�T�����q;��D�T>�ll��	��OaI&)]� 1��"O�D��%�9�����gjI9[D�����]�A
��t��ą�������
Π]�+M��t��W�&|O��ɀ9z}|�A�c�'-�܈VF/n����:2�x�KRbH�mo���n/�Ov�rP�\;b>53U�
,;�t����,֜�@8u�v BJ^z:|�Rmi>%#i��Vb�ä��3i��}�Q�$D����E�&��1Bc �=����	H�Z�C2)_�6F�ӑ)f�����K%���DC�׮M���J��c� i�<)AmH�rD�)ԟz%*�ë΍؞tA�1(�F��w₱=�����9��#<A ��^��o� mjM`$�f�<� ���ʵd�څ;`�U8
"��'��RϺt�ܹta|��,X�	�@�$��:gb[��p=����-q����v�d�Pa�A݂^�Y0�4g��R�B>D� ��R ���
(	3;�d�12�?�I:Xd�X�Gl_H�O� �Q"���)y�X	�ND�Q�Ri��'�� ��K-<�S�j��;č��ψ�x���G��'M^�B�c�+T�������q����'5F���!l$<uy�ʋ�|���'��퉖L�ܘ)#�cʰr{���'�@�sց�6/�~�U��	`O���
�'���K�B�NIf��P'S,@T6t�
�'��e�C@Q�b���D�4����	�'�b��#O���(qr�X*$o��Y	�'�	�D]�h>�@�녠ll�{�'Cr�b��,\<�@p#T�g��\B�':�I�q�M�7�ʸ[0�߮[^���'&h��@�$g�L���yφi9�'��C��^^n�� X'b��}��'��Q��+�jv�I r�_�[|Q�'��M��bA� ��_Q�D��(O�8(�(^���<l��
8�H���cđ?��$�	�'j(S�O�1L�E�#.�MN ���熳7��,Ӕ|��9O�PڧaR���X��|�`d�&"Oʥ�p tp��K��֚6p�MR��'T5qw��gJj���� G_25�h��j*��ΌO!
��䆡a3�䨔b�!�M#唇,
�ոpS77���y���T�<Aa�B�> ����.w�T���>�8��>�vƇ�{.0�y(;����[�BE�)>��P��C=�['��z�<����j���t%^�#�z�C*{�y��;IW���u�MJ�Fe�Y��}b�6"��܉s��z��� l��p=�g�3h8�f�~���6��-�j�R�K_�
���
�O���)W/��1�	�8���i+Ѧoˀ=@�BA T��=q��/���D�<i�D��1J� �C�t�-�a*�@�xq�
۰6�`�)U�!D���qd�X��J�c�4�l�r#K��� �<��*Ms;nqS#6��͉�y'#V�PԠ��]�K��IK酤�y�`��s��Y0 �BJt�fM�^�+7�H��H0�O$�@�8�p;�ʄ�sxd�c�>d��z@O \Oq;"�X�0���'i&Y��o�5�~9ӑ���'�HI��'��ԋ�N���סʟvt.Ъ��
Q�x�k��,�	({:�*�f��W?�x���] �zTnL	:D\d8!�-D���ЎJ%�Ѕj�AȹpJ����:�L�p+=}KDV���䆇okf�`�ۚW���ȷD��!�d�$��4YW��L�z�
&��$ɛ�W$���'X ���X1.E�<�'�"D<1��Nyf):b�>���U4W]�0��m�\����k�<9�D2lĞQ����+M�� Q,\N�<b�U��n<(���|�*Q{7jq�<�f�!RA��Ꮨ$sm ,Ô�V�<qe��'��v��&PXJ����J�<�#�պd�.�3��A6�4A�m�<��-X�}�|�R�\Pђ�X�	d�<�3ET�l>L�1���W`�h`�c�{�<Q��/ySh�B�Ǒm�L!mx�<���_�U�����ד�� 1��\l�<�rj�� ����l*̘ݠ�)��,�r!�	�P�S��?A��^ ��RĐ+Q1d2d�}�<�T��~��#G�f�P�GK�<�@��D�5zߓ5�>y�rN\ܥ�O�8.��9��	�{�X��"�ݲ4֛fĀ�_{(�Q�_6,���s .�
�y"N/1�́�`G�"	� �����'l���8ZdB�G����.��4a�e�A����ж�y�A�]��2A�)�(9� � �5 �Ѽ-P�'B�>�ɧj�F�����
������]�"T:B�I�|[ ���$ɇInT�uo�M?&�D�iD�@�0�߰=� `x�ր�QF������q#�'>�a� �4wfjpn " P07��E6�}�UEH2d��C�ɛA�x���ԗD���p�t�����U�2���V�S9&T��e�͈j����T��;��C�ɬaL�uRW�
N���#l�|>H�2����v���L��F��'�ڨ�S��	PfJX:��X� �{
�'���Yt��&�b�r%�D�E��!�E�p�H�����=�C�٭�>�REЗP��X*�@`8��SC����ą|���RĿG���b��;�!�D�hpVɵ�҅B%�Qn�!�d@�6~Y1��Y�aǜ�B1�?"!�D��� �V�B�^����jG�2�!�$ޟO��Tk ���dUv8�R��0l�!�RE�P��R=<VH)rp#���!�I�&,���B0�cB��x�!��M�&��̫s�G�o-��b�* ��!�M�Z��E���\̢"NGt!��o��k!%�y ���c��y!�D'=U��0�i�1k��Q*580y!�d�28�lSt�F�*�%�)G!�
	A1���'^� ��H�V�ޫU!��-xH2�d��R8�6�ҒOm!򤑑\°#I��?�����%X!�d6p���weS�W�{��F��!��C�p-h5a d�М��̧7�!�D�`�H������D1��S�_)A�!���Z�J����L�a7쳶 �p�!��Z�Wm@�g'�Z\Jŋ��!q�!��O%��h5��&M�	��_!�$�)�|���=a��,����$U!�D&�Y���3l|
,`E��?zE!�$�	M���Q,\',} 88!#Ť6�!�DZ;}~	Z�nD�lXf"̆R�!�H�4j����- 0�����>*�!��Z1V �C(�6�`r���
�!� �d�l�-2@I�a-��k�!�Ѯ)tU��J5E-A��Tu��E�D--��d�VHD��`��caϠZN��oP^S8h�5 �'v4�
t�_�@�A�%�ÖX0xJqg)@&�����@L���.ؚ���E�]�,� Ԥ\,ꂩ�q �?Z��E�O������� q����1\��D04.�*9YZ	 g��~ھ����0|R���K�|U�K�&<�Z���EZ�)����Q���)%����(��F�ۄ|��1��k�H<��xBN�#��O����`C[ 1��!UF\�A\��P\����L��ԥJJ~�Od��$>���*%`�Ґ�qP*�$��&�(�U
6M9v�T-O>�Z���8��׳D��y2V��.G������ A�x=C�����z��Πk:Q?�d�� ���*�fS�8�Ţe�<eC��װ]��h"a!G8X��t�S�O�Ν�g	Ϛ���"�H�lñȜ)z��!�i^�*�IN>)R싘h�h
�l�D��k�$��aޑ��S���D��(�3d�Py�ϓ"���O��=�}R����Y�hhg�^�L��́�OPy��[�O��HĄә=�m���ŋI��!@�4����|J��a�Q)��ܜ�*��(��  �B8�*$��G���A�%>.��u�Ѳ3������O��O��!��S��q�E)T9���\�{��n��z�`�ӟ�����}�ġ�b>�A���
�i�i��)�\�#nӢ�IV�Ĝ��O�?����Εb��"B��%�T@k!"ғ�hO���H*��p��YQЍ��M��d�C�$!&	c5i@�<o�-�u�r�xC��+ېdR��X�R�r�*`E=a8�C�	�WoZ��v��+$�:ɺ�!�U�#<�N>y��Y66����T�zpâ[�3���%c�?jw��QB��v}�_3d��fg�%��iǇ3� �?牲nr�<3tIr���0\�)�6玳C���(���>��)��tȀ���XQ�[4����EB/HE!�dŰm�`���y� P�B�� F-!�� l��4!�Y��"��.|(.pb"Oj��,�]���w�_G�"3"O�ɦ�ÌX�xɥ��?�XyA"O*ɱ�#'E°t"��_5g��lyP"O��qAP)��Pt)�r�Fu��"O�1�ӡ�&Ew�I��ǧK�|��&"O~|B3�׳=B�#.�<�* �"O�@R��-)hq�ql�,ѐ���"O2���� 	N�l�ML,>��9av"O����_�T��FZ�`��l�"O�xA���e����1T�Hm9"Ot�[d,29�o�"KP8��"O����L�S��	���Ύia� "O� ��dHu�`
� ���]z�"O��u��4`�)�tO�4�4���"O,a�!��E�ذ�u�
�e{N�S�"O�I�0�L5���D��q�4 �"Oh��KįFN\�Z��/3!Ҥ["O���?cX��Yec�}�d $"O*E�"�LmEJ��S�b9�"O�Ha�O(��Je4��m�"O���*E�A��4 �0�BpT"O|ͫ�M�@��e{ӡ�Kz���5"Oĵ�DoV*m�bCB���-�"O�u���q����DB�(,o��G"O�A����H:� &��j�"OjC� ˂Xġ#�^=TivŨ"O0�s���X���ӌΉUS���"O�}�w�U���$8��Y�L���S"O,�rq���P��tW�_8hK\I9�"OؽHu��Y���G��\��"O\}	#P�V��4+1�O�����"O@�Rb��	�䔪S��!\�iX#"O�Ժ��^î�!�jԀc�J�	2"O�ICV�4�$J�:h�F�M<�y"(J�#~�3gE,@ʊ��u���y�'r/$�!%��1�AB%�܏�y��@�l�x� �/�\E�$ �c΢�y�	b���`&.VO�(	��y�F5/��[��MY��������yb��9���"W!��ƑI�!N��y"��@��dau+�e�z{�-R�y��@+x�A�����y�TO�q�!�DF�k�Ԩ�de�(T&���3d�!��C# 7�E�u#��/����K�!�d�L`v�Q�E9/�0�6F�!�Ğ&��41�6P�]pA��|Z!򄁇k���Җ@J.5��P�B1F!�$���fiȗ%Ǌs�`L�AB�!��--%R)���S��Н3ao��]���$H!mv�����L�t��O/�y�����\B��9r��BÃ��y��_"Rv���e�@1dz��"-��y��Z�L,Xc��%���{���3�y)���<Iib+��L����-��y���8)x'K��Hb�}�PMç�y�� t��&m9or����	��yBL��%Fqh��QU/V �e�1�y�$;�9z�G��m�U��y��Q�1�S(^�l6n�[5���yҧ�`R��qaՉmfF�pդJ��y�
�� ��iRa`|�*,�ǃA��y�� X��Ũr�C�o�@�Dԋ�y�@�N�A��f�!�$���y
� *�R!�{�tpstj�(
�\�	�"O����f����Ð�O��X��"O$:�.�L���Y�Ĉ�Ph3�"OHMr��#l��CC�.`���C"O�q#�+�6��H�eK�� P�"Op��Ƥ\�}�u�D�δM���36"O�,ʤ���Yl��C@ˈ�	6"OJ�`�g�0�b���e�P�"O����$<d��K��́�P��"O��bҠS��l`R釻�|BP"O2�vk�kn�芕�N�.Y��`"O���G��@S�\���ܗm��1"O ��j�12vM�T���W༓�"O$I� j��.Lt�;s%ȠI7��QQ"OR�����EY�-h�ͣ$h��"O�p''��g���q႙m�, "O,��@gC7s	1��D1PX��4"O�Q"��VG��`㎆�NJ�j�"OZ��O�!R"��A��)d�m#6"O�H�`���^"�W�R�Z@���"O���s(8�J�AD�
�N���T"O��2��R?�(x�����"N����"O`�3Gh&s,|�JF6r���3�"OPp�Q��jOf��	ă~�عz�"Ob|ٲ	ۘ�Ȉ���/b�0%�"O�%3�3H"h8W4~�˅"O���H�>``J�K$&S<8*���"O2J!��Z��+e/��,*vt�!"O>�1�S)P|��S�(�V�b��"ON�+�f��a�V�����	���d"O z�jQ4'u<��E�	-��j�"O�)�+��mƐ4Z�I�-~��yS"O��Bhu8�4� n�-ü�C�"Oܨy���sk����&r�<
�"OK��.��$qW��cv�#E�y�&��	H���j�\���o �yb��>����cE%P6�J����y©I6i�8�fÝVv�<�!�ѿ�yB�F+@&���QV�p2!앁�y� ��h��Q��F\��HX�e,�y��K��Xh4�O3O��ٚ��/�y�@@+}�V�ᄒ�s��@;�����y��_2.�\<:�2V�<0e
Β�yR�@�_B���Ā�~�A2UO���y�9��}��*!��t�IQ4�y��V�'��H#l�:s�q��W
�y"͉�t0���
� T�w��yo��bl� �К�h��BQ�y��V
P�Z(��KA�~ȩ�KY5�y�,�!�,�J!��f�<�Q�6�y2DF*]�A�!ϰ`=��0a.��y��E��ۑ��EW�Tqn���yR�B�O��z%�N�>��#PKX��y҅�8a�u@N��������y�,0n��3�Ó�ي���yR%�p����Ӫk}�p2�)�y��a��kq�'R���[�
ܧ�y`	�J�l��&@� P1�A`�;�yr@Ђ/"L�)#�ƾ%��Eڱ�ˋ�y��Z�uVh ā-+	���G�:�y�MF�B%��+��K�$�4"�ն�yr�,K�(��0EP�qVKھ�y�*ׯ?�8������O#�y"E�'� 	x�^3=������y
� ��A�]�Wʊ��3	:o�
 ��"O��%/T�X�8����˳Y~t`�'"O���sf�<ފ|ӑ!�R`��� "O
�`2����`���N��؀"O��2�$�1C��C��+Ѡ)�'"O�t:eg�9_���ٳ��������"O��:�hǶ�|�� IZ����"O���ҭLW�9é�X�.p
v"O谉�i�?@֕1��БC��ȁ"OʈA�l��Zr���U44]�葔"O�����>|A�h�AK�ES�=Q�"Of�W�G=1K&��a6Z96�ɗ"Ov��lǵm��� R#s�b��C"O���"����q�i bz�4�t"O��z��x$����0Z\�В�"O^EZ$HY�ZrNpj����VOtT�"O���E�
$Gx���rd�M=>2�"ON�!2_*o��B��!"1��ZA"OL��L4Y��1��%�����"OR�;�f��i����>5�J�S"O2�UL�F�B��e�\�L�X��f"OhQ̐�]�,|ڥD�8|�4�A "O衉g&ٰ/T�ශ׏G��Y��"Oe�����k�B��ES5v��P�"O�(���*W���7ᕄ.`Ez"O��:�aQ)t������F���� "O��C"��B֐E"6��rX�p�"O����-Ї2�f�� ���hT�}9�"O2MHfc<2���j�a���d"OB3��Y�.���a���'���2�"O40�uf�y8ٙ �0g�����"Ov��c@ {<̛����`ң"OXP�K2,�h㢠ѫaFj�b"OD� ��""��35N�
�,�g"O��cN��W�p��ǂ��Z���"O���,�3k�����JI���"O�ɀ�F�C����Iټ|(N��%"O���6�J�5�jZ"�W�_.�c�"O ��@˪a}�$ �F=H��%"Od��q���e&�$
$��� "O�� �J˺�$H����=d�3�"O�� Sꃌu�
�������"O�\{���W ��z�ƴ(��1s"OF@*`�#`Ŵ��%cj�t�"O�i�e�*`P�إDN*1M��ۗ"O��^6"?�a�V�>[ p`b�"O�����P9�̺$�t�� �"OV��A��k�R����!:�Nii�"O|�ړM�4|uB�P��x��"O\ �U=d^���T"f�KQ"O4�P$�B���F̊�A�6-K�"O�=��f۪_aG���Rՠr"O$([��SIȄiW��	,t���"OTXq��:&��=	Eo �=l��J�"O�ek0
�6Sܼ,�M�tH�"O�ȳ�ިP̕ХƄ#'S&J�"O*���+վ0j�o�
'H^ip�"O���!�}���q�	Gc
p��"O��ȣ/V�{9x��MY�+$��i6"O�۱�ת;FT��Fk^�u2�Y6"OM�ӄ�=��ء��G=�Yxf"O ��I��}#:P��i�m0
��"Oܡx�,M2�iqȕw :��v"O�Py��Z*-�6mz׌���QA�"O� ��#�m��Xn,���v�d�A"O2t��H��v�&x ���>�f�a"O���
 
  ��      <  L#  <.  �8  �C  ]O  e[  Sg  �s  �  ً  �  ţ  �  ��  k�  ��  ��  �  i�  ��  ��  2�  u�  ��   G	 � � : �" .) r/ �5 �< @C �I �O 	V z\ �b i do �u | �� � 6� z� �� �� q� �� �� B� ��  `� u�	����Zv)A�'ld\�0bKz+��D�/6�2Th���OĴ��5�?YV̒'�?��]O+� �*^
��e�E��~�`�*��=P��� ���F�w-�p��.�0�)35�����4|��f�Y0T+�
�*GhNdK�*�.C��)цG�+86:���Q�D��)�;8Z�r���?Yd�Z�BuLd[T�\
!$] �Ɓ�	�ڈ#��&������cWAR��<6m�E����?���?Y�oσ1��E��fJ� ��a���?��t,^��GKՍ��$�O�@r�����d�O���c K�h�+�[(G�@����O����O��d�O|�D�O�!���yBiV*D��B���:�b}D��`r���Ղ������ ��<Y�ȟ:R�Y8UhG�>D��!�!���O���k�i?����xWV �c�h>Y���� F�6��U�6¸p��Ov���O$�D�O����O��$�|�wԊ�86�L�{�
Y[� ���n1��'�v�u���l��M���6 ��k@6MִBͮ�s��p�a�&ˊD���B�VL^TGz��8��d�u�C"nx�Y��4VM�a���'f�� \A������@�R,4o�9��� �v,���Ek�O��nڈ�M3����D�O��n�NV(t �K�n��|�f��-��6�$Iz`��	n�BH�ȞU�LP�F�IU�l�mZ��Mâ�i��$P�C_[�=�U�#E(yc���3�F,�ŀ'I\7�[��3۴G"��"Q���Q��CeR�9��ܧlz<��F��z�<$�R�ţ��}��'�(QW6�"�i�(7����$+� ��؅J�M�SN��Cw�C�~�� �Z�?wVD��45�D��,\i��g��^�!i����'y��c�A�>k�<�3�A���H|�V�'��Ob�D�O��Φ����d�$l^r�FuZ���-(��m����I�zm�p��ҟx��Y˔U�&�@x⼘�M]��M�٤t�R����l�p�DɊ?�^7dpQ�Xh�!̑�FT@�/�)*!o9��l�q �o��I�@oU'r� l�۴wU�<EyE͓��TGyR'X�/4B�H3kׇ�P�x�U��?i���?�I>���?Q(O\��O[hP,�Oׂj�,���<k��D�O���V���40�O���ܦ�?�?!���x��%s��H�E�����L�矌�'��A��K~�$��%���+%'I�rM���kU�m�xP�@�������D؊�n�}~h4{F��k����)� @�i��%�?@ն�˒�11d �V�v��f��3Y
��Cֿ�h�p)(@R�\`$M�DZ�:���G��\�4�Orn��H����(+ށ��ѴҬ([� �:)tr�O��d�Od��<�'q��y��R�A����Gצ4�D"yӒ�l�'��ap)��P�t��Ǝ* ��͘ٴ�?���?!��f�Q��O&�d�O���e���?`yڅ������5�Ǹ<a��r ��IӓnՄ(Y�� &�(7F1p]8�h,(rS�i�PL����Ϙ'�&xa7/>>p%
�?��ٲ�i<t�B\�����?����v�ҕ3�k�Q&����2S:���hO?8�Jʴ%NQ�t��C�XF�uy��q��TlC�i>��Sdy2a]l,p�P�+D���HoR71��}P�>����?�.Op�'���J�`�}C#�U�Vl�w�.q���U�ҧR�xx�툼OP�yBd��0-�X���ȼ��爒�U��|���������O J�ĭ(��N�ЈO�4�� �A@-�6�@�]t�����Šb6"�t�R�Fz2��� xf$��N*m�f�Ps���" &���O���'�O(��GD�8@����<���p�|�g�ZEnZny��O|6��O0��صFN<8�c���Sr��ka���O����O��D�OLA�gV9z�x,C���Q"�*��D�u��p�eF�����䎭$9���$� @ ��V�W��Ȁ#N*H�IƢEl�pÓ�A�T4��C	�SKZ�����7��O^��u�'�6MH���I�E,�䅜.�x��Ђ@�yЂA�'���C�OH�O���I�w�^р�aXH�����S�0�y��'�剌�M#��7W��A��ʃ\��1XfE���&�'Y�7�]�r-�y2�Y�w!F��2g�i>�$�A2&�%��G� v���N�RH"�'k���� X��DKƂA)6;��0�WYܧ94�0�����2`�6 �� �O��Y��L�Zd�Z�H�=)����ؐCAC�$����^FP"��F�i��Z��i�'�<���$��e �	5���lA��L&m�$��2�Ăp%��O@��"���O
�d�<���S�2]��B�	�_�
��W�P�b&������M����&�'Y��
6+�9&����
 dՖ�� dz�v�D�O��dI
C@�|����O���O���kޥ�NI�Irɲ1�?)��ر�Z7�гRW��9�u�[+�zݖO�d� ���ƚWU�pX���	���a�*�	۲(�#Ieт�Qo�.�pb>��$?�Eo?^�]���	%�����M�]���&����'�b�'��B��V;|�z4"2�K)F�`�4�|R�)�SH҂�b�G�$��M��=������)e��O��i⟘�3H�P�L۱"�Й�F�:���II#͛F�'�B�'r�IR�T7�����P�l?R	��Ď*�Ҁ{���sPu���	>l�H���!<O�����C&%��pB�	����� о$A���0o�>t�lqx2�E�9L�yJ"�]�={TƁ|E����Y��^:�?1׳i�"=a��0��Ǝt��q���>F2�|��'B�	\>lx�BҧJ��I����;R����M���L�vij�`˧vFaZ�i�r2O�� s��Q�Z�k���'���
��'��I� �	�|��Y�V�BPK��M3��
�4� �ݻ!D�>~u���h�6v��I��'H&I����W�4а
�c�$�`1�O�P�}(3�ͱ,�`�8���7�6$���ă�iK|�>�' N@y�kG�b:�S�C�]ܒ<�J>����'�n
dZf��b�((�Gٮ�����ۦ�UN�2!vM�晃Q�6!cㆂ��M�*O.��u�Xۦ������O|Z8�p�'�h���Oն #R1H� �/9������'�2#ߘ`nE����|O�%���Y,:E��A�'4��S�`xB4`��O�.�����C��z2�J��A>\�L�+�
�4��) 6��7[��O�,���L�n2�w&�)u�p��Oj 2V�'�F7m�j�O��	�4��|��IT�av�Mڶ��;�!�d��!��pJ&^r �k�+~џ�c��)��C4n���Y.da:H��B�.` 7��O����O�\K����J���O��O��]�z]�Y�#���M�v=J£C3k�6�����@,�'oW� H��u�>��7�ē��])ẃ�@C��+�EIY)R�"��D�\l ��]S| ���LP̧j4|��v$��p�5�ۏnv���G�q�n����O��>��$�O��=�����"v�> ��ȋ��yR�)0x��"�
wm@YڇJ�,��DTg�����'��I�~&����pc��q�!�2F�u��L)kvZ��	͟�I㟄�Ywq��'��	�	� h��,p���vDL"@�G�ݛ&�<MJ��U�P.����/��_~���U7F���+r
�g��E��NP��RǺ��H�J *p��AD�!£YBn���o$d�
�ЀoY�r��Ȓ���?�����'�>I� ��eN���C�� J�����3D��[�F� �4%ŏe=V� ��-�d���IMy��W,f�b�'_r�����[��U�l4h�UDZ�]���'-ᡆ�'H��'�"4��j9�'�⨸��z{��Ӂ�30�B�'%ZZ0��~,�,(n�2���Ѡ��p�OD�68��#�J��
e x�B����O�q��'�x6��[y�쒤~�T����E�b���ƃ=�䓛�'���'*"?O6)�^�*��N�CH�@v�	����'�6mڰLF����ކM&$!�I*hT�n�֟P��4k�\䂂�i�\�t�O���2�$шBe�8X@�Ĕ-2�'���!%�iN �	�3cx�lZg�')I�]�� B�GYUG* �[�|��O4��1YFod��g�Ĥ{���)įŹ�1������</�����BS��JA꣙����o�O�n��H��<k�Pz#ɞt5hp JQ�,���Ox�D�O���<1���ͳX�����/)/ ��͗
��Op�o��M��y�=��9�#�Ɉ.�[��� )�xPa�t��$�O��Ċ�d!�g�O��D�O���tޱ�K��r�����/
#�ȣ�螒L�YK�Ǹ",�`�	�:�0c>��seG'���9B뢱��	ҔnW�9�������y���@�ߓPE�=9�iS`1v�H�'�,�(�.2�9���J,SlI�P�i��Ub����?����R :Q
���
g|�0�6I@	Ҷ��',�Q��Nח~����㑍���R/O(Dz�O^2T��p��&<���An�0f�4�1f�2y�lb�M�۟������Q�T�'�b�� �`���Ҫz������ VQ�����L�)�������ڴ"���"�(O�S�����F���͎%S
dz`$X�L�0)Z�:� ؊���!\�b��L7�(O�ps�q]l@���=cL�����=2�f��n�ӟ,�'����y�M�z29j���r�8�1�R�d�O���t����=7��:���1(n6�����M���W�B8�i哤o����Yw���'0�q����0x��Ӣ��W��Iz��'<eթ+��'Z�I+N4V%�SO�t�4�{�@��1ZT̒P�*H�h�)��ӫ*�8�a�I�9q���D*I�hU(QIߣ	��`5J�-h$*��E:h�f�`�ݾsr�}9�-�928���d� _���?�d([��Dc��]��`ұ&ə{!�$�#^�I"�E{�^�(��
f����OL�A��$W�����˃�v%�a�5�|�Ɛ\9���?Y-�������OY��Ǹd#�d�N$$F�*v�O���M�!����a$<P*ݣ�]W���Z�(��'�J��+{��PZ�O@vU�9�'��yh�L��`hr�]�X�*��p�"�����A)ҭQE���jP�)#���Y�I�O�����E�IP�Or��{#�5kD�� ���(6��N>������O��r��R�^��gj^ 8�^m��'/ў�Xݴ}�6�'5J7�z>����'ɬ��#��q��i3Nɦ���ǟ��	,\hj���ퟨ�I�����ۼ{�Lܱj���M�%
k�Μ�d�l�5o��ܕ��ުP���|�H>9q�R�H9�@y��<�6����� 7�0we	  �r�2�,�PnM�|RI>s�E3{<L���bΰv:,*wԟ�' �tP��?�����'ͼq��-��v)��&�Wg�y"O��ɤؐ$�ۡ��_�v���X��3��4�����<YCH�)�nE�![�<y>x82o�pr�d'�?!��?���'���O��Dn>E���Ļm������/�*�0���h����=�pl��ψ�7�dLD��� h�[&KI0e�5+J:.df� �[�u2b��T�_6J�r ʁ�:�n�֙�3,�6�y9�I4{zA&�ퟘ�4Q��'�r�'��OL<�`M^�'���E��U�l���1D�����JYQ��E��i�l.L2�O��oڟT�'%h��0�~���D�O|̢g@�F�M�0b['[��D��Ot�Ď-:.����O��d1q�"X�T/z�2Q��7Cr��1gs^pӵ/�*Z̸��ƍ sG4�Y��Ɉ|�Ԣ��"{�V��`�c�9�1fŀRG��Pt�	�)��q*��O���Q��	�e)Z���¦q��4�?�`G�|Ԙ���ҿ�����������Oʓ�0|��U2zJD���8�8Yh��t<ش4�F�Qe�0=��Î��D��i0�	5{��H#� X֟��IU��� fR��U7 mr��#[�[;�i6B�O��'� �*���RC`���'`��#\>��Oi0X�F�7�Ĉ�!eL�z���Q�O�Ax��a�!�� ��	  �kXn���#��tK�bX�зA��Tm��E%����\B�k���'>��|���\,W��{5��o" ΓU��ퟀ�Iן��'���?m�"�� c�`т�X;> <ᒕ�3���6�nӒc>��B�ɡ#�Jy*P�-k5�貵������,�I=ߜ�ж#џL�I����	伓p�RvUfhʕ�)6�K� :g��i�C=�?YQ�M�d{R��|�<oP&q�� �c*��}�@`;��ǈ"���;$�C�H�{��ǳC�>0�|⥊	o~bg���L"3��M��u+�F�_p�'��u��Ϙ'�97��9jAI4�ƦrҦ���'�8m�%��j�H�����m��.OT�Dz�OT�'9^�&ʕ�~���#aǵ]�`�;�,]w���'Q��'���u��IП�Χ\b4UCR��(��x�5C�tu�}����/'f4���n_Đh��P*V�-;��+ʓ;R����0]LЕ�ןuU�ex �J�R��&�k<�p�#�5�]���8�}�5:q�]	 �F����	%�Vty�˟��4|A���Gxr��%{�pt Ƣ̠[4\,�c	�y�.��;8�q��-��@��F��RU��'d��1L�p颪�����]���۴b��{��׀D���O�HZ"�OZ��d>�aW%@���=z�ۛ0d�T�����&��������-o�*t��윅�Q��,S�*�" �g��6Y����+�Gz�Y ��(Q������'�<) ��ן�Q��a!-�O\�n�����!$x�0,]�V���0yy�'a|⃔�s�.̑.y�<i����?	�']�q�F�٠3��� ����������C����D�O:�D�|�f*)�?yfm&,���&A���F 2�!ޟ�?���dB�����	(Ty�� q�I<+����OkZ1qw�?�)�1�Rc����FL\1`f(#?�4��^��S���I����4�ʳK�H��_�y8����Ȥ/�^�$��q��H_���O��}��'�>��ahє)orC�E]�M#LP�
�'�(��稙"
jRD��)=/������A\�O�8�:�ЃX��C���A،�3�if�'=�EZ���se�'�2�'O6�Ҙ�Tνc�6�BA�Y�6�鸁ⁱ`�4���N1.=��زBݎ<G1�<Y��e��~ri�0Z�-p�_	11�� R�5�E�&R�5�2Em@�%YƘ��>�)̂%-$��4�t��*h�0�i���'�P�I��'Q�	N<�d�Ov�=IA�PC Jp�6)�#��h;��+�y�U(nĢ�C#�&�N��sΚ�����r����'+��$�:P��i� �X�g�S<r,�#<�����˟|�Iş��؟����|"шJ�s9.Y�@e�3}��rRn��M#
�zw%[.;t������M[@�Ig���Fy��0h=&@�t+�:nz4�5@�'�t���cz�ҡ�� 
�od�v�zQ��S/:�I?p�YZ�@F�W�����X�s)L�tb�O ��;��O�;�Bֆ~���ҥ�M�c��+�"O���"�HM����7�_��|��|�(`����<�OX�A����'����2�7ȋ��\c��[�#���'o"Hb��'�B=��`� ?���S�*V�3�� iҏB6	�0�p�h��!UGH�c��ܚ�)^��(Ol�0��x���E�s�(t3��
*
H�2�d�+!��)�6�׼E�`��C�2�(O�9C��'ٌ�O2���f
+j�2�(D��A�q"O�p�e,�<`N��1�M[�K��,Z��'@Z��� 8��y���C�TԒ���ג$S�'JV��wӶ�$�O�ʧZ1\���N�2ȃ�'@����eL	:��81���?���O�i�!��(����x���i�S]�aӠÖ��r���6�����2���v���D�G��d��3��y��;�S�9L�a"ڐ[5�F&UH�E�}���M��d�)�E����"ϓ8�n�#�iA�9�'��|B�ɢ?Tzк�d�q;D=C�HK2Eʢ?���iB�6�4�䌲pC����Y�f���St�]�b
����O���O� j�	;BN����O@���OX��;Q��9*aCU�4�2:���E^>��N�z}���;Jv�����{��_#k2���R�mN�3A�N�"��u�U�)��7�3DA�\����� hP�D
Q�Ĉ�  o�6V��f�t��'~�������͟�'�թ��ό��h�T�3�0����	j�@�!�B0WZ�{1Cˀ7����R�<���i�$6�.�4���I�<�s.N�*6��6��1�����*"F���H�c�-�?���?���"v�n�O���k>��Y`���@E
�ڹ{���~�a *yF���!m������J�&���I$y\XЃ�/��t��9B�9:�F�(�f��H�<�Hf�6)�M��%i�m��R�N���"VkQzTL}t���U�(������d�I]�'g�Pۄ*�24P�y��J�M�!k�G#D��{�GR4C,����:��a��?��֦��	ky���*V(��'�?᦮_$
�+%��)�|��_��?���$t����?Y�OO�p!���8�T\hj������C��	�c��]���C�+G>|H��;�	���(O���*��M�:5�K�ʣ�4y�<u����X� ��+�&Wv���^�6�$����R�D�B�'���y�
��Qo�V|�\9G&2T4�O���Ċ<�m!t�W?Z���ͭ ���%�O���ĭP*��-��A9q�����$Y�0dymZ��x�	M�4k��Z���S�E:詋'c�$c�J�*�ǋ�8���'"<�{5���2p���\w(:yB$�G�S�[��?y�"L�3E|�P�Ԉ2y8Hq��:?�&��P�0���b�,S,N:���x���������́o6�׮ŎvV��/�I\��
9�����Q���	j>]�-*l��Ѓ%K4�����)D��!r�&K;9S�ʛwU��&�e�>Q!U/yY۔)�T-
9IW�Ŧ��������#!jq�I�0�Iʟ��	޼���A,"HD)P��a`����%P��KB��cxF1�S���|�l(r��I�|����'[�i���/��r��4jN�����k��=iq*�37ĸ���K���O�d�buB�q?�FR����K�c�<	
2nC��Mkt[� ����Oz�)!&���P����.P�uS ���Ed�<qd���Lo0e���.g��i�(�byb� ��|�����$!a4n�ȱAڗw�d[dƄ�gi
e�r�P0��$�O���Ot��;�?�������
/Ȅ,тL�?Ԕ��)A�E5�Y�jH&K��S0�@�s������=B�X�Ey�h�	R���%�=��Y�'��&��>8<����h��Sg�P��O�	�TFy�`H�:dld�G��mV>;��"�l���`|��kW���x�C@���8���A��ym�|��}qfD��(*��:����W՛f�|���5�*맥?aV��3��y���@yfd�@T)�?��sQ����?1�O����A&t�g�0:|f%:�-*_�l.t��S� �?����*ex`�Gy҃'gv"|+�&Ԉ��2�mP4eA���h�u��=���1�"�[�b���9Gyr�?�$�i�*���4�$5^������p�%�ԇ�	�zw���0���DHȚ~���ܟL@b�	i�<�W�ٵ-�� �Å�O4��?�2�i���'+哻	� ���\�<����S$V��ƈAT���I��d���IA��tI��T�e�ҽm�:��N� ȼ'p!�aI�P
�&!؆��D��/
�bjN��� Զi<�读=9�!�������͠��B�G�Z�§�� �A��O()n0��'�?1������lu@TQG暀!k �{¥M��䓸?��R�>%�V!�/C�Ġ'�2Ch�F{��'6L���O�u���H#؄��s�)�!�İi��'Db�C6/��y�V�'L2�'R9�v��UeF=r�҄` ��r͒I�v�K�w:�l"���<�V��$���y�1���O�V���ś@cV%S^���	3�����^(>F����[$&c�,�|�H>�2l����q�
�~����f���� �'��)����?����'H�C��c�����We�Uʔ"O�) ���tQ��7/���^5X�T�����4�����<ig�g&��O�p�^�2�+ r��Pd��?���?��Gf��On�Dz>��@%��0E�}��/Ӣ((���dL�_LpxkPS�Z�����@u�F�F��ͅ{�:��B�ߋkmr�#��'?|�\�-ΐB������5JS��� �I79C`�Vb��M��F��p�@�1�쟌�	��d�?����-5֠q�D&rk���R"� ~!��D�MEze�''-�p�H�0v	�'^�7-�O$ʓ�bq�b\?���r�α@CKޚU�@MZT�L9Zl^T�	ϟ�Y��矠�I�|�q���kWaơa�RtoR<#�t���,{n"�p��������Ԅ�4	�e�4,���2eO|*�'�!3��e�μ
T�1	�)?�C�\���ߟp�'�y�@�=+��|���B��$�O>)��0=9��HfL�ӂ	�̠s�w������!�,�0!)[�	w����C��17�	^y"#N�6M�O��ı|r2(K��?A�bɕ)WJ(C��8\r�rj���?��\�F � �
����`��ĝ18���VY?	�O2�EpTě�,u��[2]�'����OLxRD��N 8�i��H��T�҄##�Ӣw�>0EH	�j�8eXE,S_,�W��u�IԟE���'� >ȹ��E�7D�U�Ns��eR�"O��+Gʉ&,>�ԑ��ER�|�q��ɖ�h�*�i���A^�3Eܕ~����"�r�����O��dʲ~J�A9 d�O��d�O���|�e��'p��Ի�j�<}X�ZAX�O}v�KT�!/��e+I-Bw�c>�&�X�d`J�JR�`X$ʜ�SB�\µ%��{jlh�ǃe�f.2?.]��;��T91��Bc���'E\���̿=fh�OR��q�'�1�1O���qM�xq��r��6��ٗ"OH�� #�tm"DD[��d�`�Y�)��4���O���E�P��S0E�,-�� �/��
,q���On���O��$ֺ��?�O@�����3hP؃��D�6� �j�v%�'J��5��I*j&��+���D4�̻��<J��!3ē6u>�aWe����z�-�D� D$6�d|�T�+o(X@��4G��x�8�X+����ѥE�4�"D�'?j^ ����0=���e�41��e9t� �L*�A(5CV��3��F�'7創5D���4��	@b9J����NhP��W�,eJaxb/\��O���St���/�(_N����'��(����"~�hU��CY�FZ�=j�E��ax2+
��?��y�̔�x~� bc���8*��#� ��y�BP��cE�"<��B/^7��?Yr�';<l�eJS�7Pl��K����	M>i����?�B,y~bS>����6U;�n�pm� �Pb��\�Iퟸ�% F8>K����<7��m�S�O�D�eB �x B��O� Ll��O�M��P�|t���\�n�}�ǃU6Ѱ\��II��:�*�GDX~"%���?����h���I2 ���"�\�46�b�'�6�xB�Ɍoz8P)R �W�6��,��B�?��S�=�HM�w�(XL���!�\�f�4�d h~��8R�����?Y)OH�!3�#{�aP!dio����"�`�ӔG�ߟ��aG7L�c>c��p�j�5��9�n�	��"�JTG��5�e��h��̓:u��c>c�p�LR�hU:��ʱz1���I�O@�`�b��	�DF{"	ԣ\���N�(aAr�p[r�Q��'��q��GʎgB��,ʻ,ۺ��*O�aFzʟ��#UbD�p���.��`A\��Pu��r��YVnm��ՄF�2Q����C��i�*���߿"rH6�����eIL"�[g@M��P|"�O��O���OB�cR�wa�(Z�A�-� ��	6"Q���$E�_��	�Q%���g���y<Q�x�dɝh���0�#��Ӥ�J<={�1#,�3I�x$ێ:��@�S��:����O�c>��kCYҡ���H����a�<Y�i<��0!���2��%���©���	��$��X���F� P8���t
ōf(��|����I�k�d��	k��!WL��d�'�(A�9v�x���[�\x���'>j,�􇓐gtf���,~&�7m��hh#�2�X:⡇oXJ�˵e�2r�1j�t��GɠLL5J��Ԧ��S��l�>YC �ɼY��Q�O�ٌlۣ.f�����O���.?%?�'k��A�햄TyHP�7S
!�`D��'`�1� M/l&�t�KaR��hO�}F�t@�&&<��1�ͳe윳�*�+Z��%�'&�@��w���҂�O 2�'��O��D�4��UJ$(w2d�&��2��T  kq��E8���l�Z�9�B>��;���'�n��M����e�q���d���TkK"'���gڡ6(B��aJN����O� �>����bִػFH�)������Jl~퐐�?y��hO�ɾ �~��g�S;� !�k�nB�	�$�lC�)�bR���̩�$��I�����'1�\貀	��6%0�j��##���0��'�r�����矄�I��
Xw���'��I	�܄�t	�9i|ĕ�t��2i��8@(�9��vf�2U+M���%b���9fr�e�WF�cːH���3Fc۰ܰ�7L%-�Н �
�%c@d����֫/>��\�r.���jV�$U���Z 
��B�'�
L�7�2�&�ɐ�ݿ^���'LT�rV�ݧM�����B� Ǧ�c,OȐm�ǟL�'�\=CD�d��]��g�O��S�+>���� b/N��C�5�&���h����O$�dPJ��%�r}�Mbs��;��)��Cܡ"���� )b%�����=	ظSQ副"�>i�I�9]���%}
"RM��(n�䪥�m�V���̼p*�\���w�H= ��IӟL�|����3���$��$�Bh��!Vy��'P,�P��Q~	���	�j�cw�	+��L�ªްT9&���iDWt ˓Y>v��p�i�EY��'�ӹK("�����Pҁ˙N���2�ئw@�\ �̈́��i&
C����KƅG���"��y��{�L�f�''��YC�d�$B�e���F,�L&~�/��r�+ٹ9{\�X5�שKεk.� Q��Cm��zsm��Q|T�t�ЦXez�4����	矌����� D�AB	٘����.��D�<"�"O`Q*�+�0�ʅ�@_�r����퉷�ȟr}�bo�8��;A��\����BV	���O�Y�IY$'*�I�O �d�O��;�?Q��$�����P#�!���<�Tic�LV]G|i9���ZL��ȟP@Ӓ�I/��Ɏ���[�n�fA�DK"~N�D���@&5�$���6j���"B���r��>��J��	�l��&c�kÚ�q@��Y~r-Ƃ�?A���hO>扨lpƵH�A�Ufy`T^�.B�#}_�5pg���=d��U��^M���|���D�'剴+���å�Q�0���+		��F�Ї98���I����ݟ��Yw��'��i�x���h�H���ad��5�2�0�$^�X��}��d���^#> ]���S������W$b���͌�M�<5{���>޲q�d˷��y�*ި%�����7����$G��$�	�hI8��²V��x��'Rў E|�#U�r�`[<U_�����2�yB��*x�܄	��C��`Ǎ@ ����Ȧ�IoybH�2D6��O���{>U8T�F \�d��w��fL&<(D�O���/�O��d�OpIA��]=T��q��AC�P%:��i>���KAѪ=�)�&~�@�0�6=�9``/��t��e�����H��"%Y�d��X�&E�&"�t��Œy�@|F|�,���?�'�� &8b,�b*G0dB�(jvr9��'f��gN�
j� ���h�?&�de��YI剙^Z�jQ���*�<4�$��iZ���?���?�,O
�'��	B�)Yp�u��й�b͈����<q������m}����:"bmc7��1�����ߢ��'��F�x���A�Ӎ:׸���O�[fx�W�ղD�\�9ٴ�?�u�!�yȘ��?�������y2�7l��d�R��$(���@ĢNd�i!��iRᐳj5�9O&��tڟ�^w!>��Ƽ��j�@5-�)C�ܩ��h�bIj��'�ȝ�%��$`�E�I�����4��6Sd��d�v�
�� ڹ1cDyg֟���)h���I�<���Unzݕ�5Oz-c&��F���;�˝TԪ ��OD1x$�'����!]����?A��R�k��@���s���j�C�.7X���'�����?�p�ĭ�?at�'�����M��
�D��	B�H����@�b�ȾM/L�[��i���I���'Dv}Ӧ��O8��ǟd�I�?p���-|�r1�!�		�(yT�Ƃ$��<�����4�ɗ�u��'H�$B�'Kf�Ik�f�+�l�U���$�R�������:�dx������O��D��r��ş8��5�Z�-�f1t�A��]��<��4:Ӌ��<y �ݻ�MCĺi1���'g���4����R�''@d�2I��ɳ�
@!XT7M̃/���l5����?mZ0�/O�t���W�f-�7i��!�)��˾+��B�	��z�sfoh�1�Ȱhz6-�O����OX���O2�D�O����Ot�����I�&H׈�[`Å-,0�����i|��'	��'�������ߟ �ɖ.���1%��i-�i!�f�8�l�yش�?O>��?�O>I�O�*5)�l�j(UQiě*�&���4�?����?y�9���]��>)q�����1a'�l�^@�g�X@}"�'��u�'���{\�@����zX��cR�'&2�'��'d�P��'D�`1%R���X4��	0�t��'��'��I̟��O��'hB��tjC�[`杩wD�u�J����0ׯ�(�F����W�H�ȓv�L�)��l��SՓ��ȓdWZݙ���jo� ���
*��8V6�	�D֯O�P��n�ζQ��,:~��!K��m�f��V��E~��'��'��'�\�[T�س�`ʷ"�)^��+h�<���OX�d�O@�d�O�$�O����O��T��a�d�ju�R!�ɦ���˟P�	�����@�I��,���$���5��$���39V��{��^#�M���?Y���?����?���?����?1F#.}�:X���<p��؁��J���'z��'>��'�R�'R�'����%_����G��P4b���j<`��7�O��d�OT���O:���O\�$�O��D6]�d�3�Ҵd!*��F(�	��mZ�@��ğ��	؟��럼������ɠ<����@��֔�h�N�6�J�4�?����?i��?y���?����?���t�a�@BN'v�Z��DMG��f2"�i���'���'n��'����iZ�>[�w+�}Ϡ������7�Od��O>���O����O����O@���V���v(@0_�Lغ4�S�
h�	oZ���Iȟl���� ��Οp�	蟼��1t�&��E޳*�Vi���Ŷ51����4�?����?9��?q��?��?y��|w�hs�h��;�.o�NI:cA���M;���?����?����?����?���?����:\�(H�ː*jb^05��-O�������\y��S"`��$�9=�� WF���qnZ=Ҝb���
��i���R/O�����L[*a|D:ťW�g�.��~Ӱ�	OyJ~P�#w����*"��l�$���c�*G���ɋQ��p�ǐ>���F{�O����f��5Is�݅W3ıt	?N�_��$�$�ߴ3�
��<�� �H{#�ʈ	�P ���1u���At�D~yb�')��6O�˓c����5ڢb��j�g�~[ t�'���3CA�u��y�O���{�"���k��J�b;Xтł�T�L�� �0��<.O���&�g?i��	�	�x�⟠3ą���ɟ2�47^p��'��7�0�i>���+86,���#͍)?���e��<���M�Y�x ���Z~�cʻ"�x�f���юȜ*�X(��N.a|���Z�'j"W�4�|��Q�0�R�\�(�(A'Xy�iӊ%hg�� ���h�0�[��܇r������<Q��0�.O���c���Iv�O���ZU��:
  �B�Z	9K|@u�.lCpe[�O����J�^���R�&$���yb�n׾
�A!��
��������<�H>ᔽi���'vx�A�*��7�"���؈�*<���Q����4��D�O^7�}���V&ԃi�|�	��J�G�Z�v���hL.8�9O��I�H@)	Ph����������Pj��p$'
�p"�1"C47�ek��%�?����<E���Z�ta�d�/~z4�P����3k�6�����Ѧ��<q!�$`�����F�`l-p��G�<.O�7��Ӧ-���W~e��mi��ݚ�\H�Q���Q�֔8�L�bA��q!��T��q��'��i>�'���M�@H���!�@	#&��p|� iӀ����d&ʓ��q�0S�"4%�w��NyR��<���M��'n�O�Df�Op�	��*I�I�X9�HS�I���d�B�z�8a�'��LR\w�Mx��>�O>-Gy��Т�-�?=U
%��%�hyR�'���h�3?�Ծi�\!�h@�!r���Cϝ �5�V(I1�����9�?�g?A� @�ٸ�hݼ�$a{3n''$l	ش�?��ߥ0nƑ��?�q�;S=���V~2�ϯ7�[�B��w�r0�M�PbS�<�������ş8��{y�Ofe�k=\)`�3!��}���8P�i�b���'%b�'4�tW>�I�M�wX"l��.[�KFU�'Sv��XR�iq�7�ҟ��'
�D�O6�t�#V��I�'���X�D^,A�%Ұn	�ocD�`2�'c�E��(گ'�x���|�X�$�	џ��NΖg&)�C̓N�(�L���'k�'�I�M�ǐ�<���?�s�Dl�*�����
�V��
�#��'�T�<̛�K�(�	j�TJՖ4$X��')	�@�e��?���z��Y�-� \ҕ�,O��IB��`�V�~�h�!�-5������)��Q���OF�$�O�$�O��}"�'���!D%t������0��<���Ǜ
��W��'&7m#�	�?m��$2��f��}"��ɢ�V���ڴL��6F�R��B.͈6��d�O��36ǖ ⢙Pg�@=$M[��U�.%�dK���"ƌ�O�ʓ�?���?Q��?)��[�<�2��G����{����hZ�.O �o�l������IO��&��ņ�?a�x�dj ��@�fZ�xQ�4h�vB�ON�p��矜}�D��t,���Oʷn�\�s�U1y�>�#���<Ԣ<�p�ڠn�������%q�
��I�y����sdH�V�˓�?���?���D�ަY���蟄z6��7G	,eb���j|6bȍ��!ܴ�?�H>��X�L�ܴ`����O��3�Ӿo��t�G �7J�,"di�i�<���%�ɓ�C����|�/O,������i���)z��Ӑ����<
f�O��d�O����O����O�#|�dh���ؒ��Gڌ�[����� �	ɟ��ܴrJ���'��6-/�	5*a���C�X5b �1O(� \��I}���]�韜4�� �XJ����hP��D�>N\��T_5,QsckS�P��eSEEŸS�&�'�䵗'��'���'�}b�G��G��	ҵ!X9;m6����'[_�Pq�4Yښ!��?���ڟO	��ˢ�U	���� 4���/Or�'�7��Ϧ�����'�:�l�>�|)
��S>��:BB1��Tfcޯr�^@+O����b�µ�d` �ɨ<�Y����)���I�N=4��?i/O6����(�Ms�;�j9Iӌ˧^xȨ ��1����'6��OƒO��O��D9sX�����$�x�2�
�TS�6m�OF����� o'��O� ��-�&-@h���4�T匪,�D�asb��0�S�(�y�ܟ�'�?=�F��.[2�
a�8j��I���pϲb����w�S��M3�w=���B'7��9Bƞ�`S�i(��',��7O���?��ܟ�C@�� )����$t\��xq�[���3�_�H1�m�	��⤀�mW>�aG{�O��dU�︉��k�~5*X#�l&b��^��$�\K�4G����<y�(Ƚnnp-�"�U��q��dƆ�?�N>�"T���������T"[�XZ0�ܯ?���O0,R�'uν!�GY)F:�|��O��I�Q�|�a�e�ԁԧ�>�pa�E�D��$�3��<�*O���5�g?���@�R�6���i3�������\�ܴb�"��'\�6�*�i>Y��ꅵX�N���>$���C���<��4;��6�'��u5�
*�y��'��s���U�l�;Jn�ZT�/!����!C1��'��'���'���'���'��d��Aї�f	�3K/%rl|�X�2ݴqX�9��?�����<��$�(��5�#* (B�0��u �FG�	7�M#�i���(���@�	�+ J*�ȅ� b�Z,	�cȝ.dP)f�]�E���7w&�ggޜu%r]3H>�/O�����X�$�W-Ðl��-pS$�O��$�O����O����<�c�i�
��'�� �%���Ll8N�"��9l�����'M�6�O|�O̙�'~j7��!��R�"�#�l:@��=*pi��/H1,�	
C��I���d+]O?�;�u�k]��5*sEы>��+�@]�b�`{��O���O����O��d�O""|:��5T�AQu�i;��A*�J���L�	֟(C޴ �8B��?��i���|�"c\��I��Jߡo��t�.�����'��7-�զ9���qZ�)� )z�����o�:�z'HD�I~-�!cȬ<Q�� w��l��Ĺ��h�oy�'�"�'���|}J��e
��� �Ӏ�6?�b�'��I �M��AV?�?1��?������.C�?����^�S�K�A����d}�hmӺ�nZ�?�L|���.a�-:��� {��A�-N���F�0%�`�Q"����hMH������Ol���/�(�2�lФ1��l!��O����O����O�����p��F(��d&J@hQ
Z�K(t�c��9Ġ�hF�'��f���8��N}Rhs�Ȥ�$	��g�BI[�f��蠊栉Ȧ}Z�4u
R�PW/B�<��'+�)b�	x��y�'�T#p��j�n Zu!A�TT�@ju�'E�şh�Iݟ,�	��`��]�4��J+`�ZD�P��%"EK��g��VK�<T�b�'���t�'|7�~��Q�a<'�h��b.ѵ(�,�J�l�Φ���4mb]�����?a��8��q��jv�����7kC���q|I@֭_�ĳv*�,T�P�_y�'��	ޟ �I�����)g~�D1�`�cȆ��	ٟ �	ǟ��'].6�3^{<���O��dL�8ˀ�`"H��/����G�ܾ\���0��O �m���M+#�'��S2'�b�ؗo�=1+���*��Lk����O��3D`�7����@��<��''���6.�y2�S�WԜT���B�$���ЀjQ&�?Q��?a���?��){�l���E	c+б�ЮۙR�ܵ����O"�l6��}������޴��'��t!����8f�C+/�� �E��.��s�>\m��Mk�l0����?�W���1�z$�P�݂��� ˻[�Z�A���D3�-�N>)O����O$�$�OX���O��Bb��X����#GK!yr��<i��ii�0y��'�B�'��O�r�H�B��8a
�6b7�`Q�ǎ1l��sS�vGy����IS��?a�S�J�Ye��S��lrV	�)d�%*V�[W��H�'C� ��eާDYT�P��|�U��"$*����I�EIT5$���ʇܟ��I՟H��ҟ��	Dy��w������Oة��IR?:��*兹E(X���'?07-�O��O(I�'�26�Ʀ!{�m����C�̀W��y��f��Y�n�(b(,=�&�џD��#S}�V��c�MZy��O����$F<T;�!T7Dֵ���͡Y���'Y��'�2�'xr��q-r=p�J@�,�A��EX*5$F��O��\Ѧ�J�$?Iu�i�1O�9�@�/�) �D�;=(j���O��t���k`�\��O�g<��S�7O�ս�K��-e��U�ԃo��[��YE������ �hO��Ļ<Y�'ʎ(9է�6���fB��_,�����C9�KY5��'���!~̚0�1f��J�:�L�",���4E���n�<9J|��'<P��rAC?.?&��4KH8̄s��Vʸ4B��e~R�O��i���ǤK�1O!3�я+�Q*��i�\��R�\�Icy����O&|nZ�OsȉX��A!.w�0�$���my���<?9��i��O��O<�d�����
�M]0}md��΂w{�6��O�H�a���L��d�O�{c���c��,Pu��D*�K�0�q�Г(t(���WR�ӟ,�'�?}q�É"{�=J����a��8���Ҧ�QD�/�	�?=%?%#ش�y���3� H� �����2ɍBb�i��d�<���?-�I-	d��&i���6H�I���k%��:�8#��̙t��UԪ����CN����9O�\r���8�6h�S+����s2�'{�	m򉐕M3�A_�=�t�#q�"8i�Y�T.ވl�v%I�"Ǿ<���MC�'���5N�b)����%�n�)4m����O�]2��M�\�ܤ�"�����%��i�F��<q� EC�(�
c�܆P@�h�џ���h��ʟhD��5O�(f,�[�去c�� #��C:�e`��a�!�Ob�$Sզ}�?���/�e� dR�:�ab͜����b��(���|��\o�gCF�;G�|�X!ga̘k�;�
q2�إ�T1$�<C�H�|��щ�A�I(����O����Ob�$�OB��8Z �B��-!���3�U'0��r����G����'���iE'�f0����R �|�����'��6妙���ħ�����h3�h�-4N�x��ڃI���2��%(O $9�"T1�l$Z�,-�d�<ASf��I!�g��/�~%c�^��?y��?��?q���D����2`#˟,�A�Ng�I�4 F1'�pu�ƍʟ(#޴�?!N>	�\�*ش.����OL�1B�E2\p�`Mo�>%��g�#�� ��'�"�S+J�"�C�γEX���?�9�;O�� ��i���z�B7=S�x�I����I�����Ɵ$�Ic�O�d別�B)JA�p����WX�đ��?����vˏ����Ҧ�<�.ˀV�4,�QF�5D��E H��?y�O�qm��MS��?P<��УL�<a��:��q�ۡv{.0�a!�n�$}�uꈐ|�IK��#������O����O8���)���Xv#/��HP�A& B���O������y��'�B�O �	�`񂵩��]�N� �@2Y�剞��dצ10�4t�R����OÊ��HB%+hi@!(�]T���!JM�d�s/�+����?	R�
ļZ�&� ڇ�Ǩm������I�g�V�C�D蟘�	��IΟ(&?�'��7m0� �-� g�*~��T	J�-!+P��f]�r�'@6�%�I*������Ј]�c�Eiえ%��Ah3����MSc�i���D9�yB�'v��eH��@���W�lQL�� ��1�J�k�6䳖�R�p�'(b�'�2�'�r�'��S�z��Q��ԡ0X�7�[62���l�.
w*��'������'u�7Mh�t���֓Ka4��F W?$rn=+uǂզ�#�4��_�X��?����E��qV
a�ܲs"���0I%��$!��%3��,ر�J�O�X2�G�h��fy2�'���N�B�65IQ �+]�4Y��$3B�'B��'��I7�MS����?9���?�IX�S�3��ӥ:�P%��U���'��s�f�`����V�t��/�~H�3a?Zрi��HF=�?��7>L����j)�+O��IM]\,���b�$���(ɛ\��X0c�m[����O����O��"�'�y�k6����A��+w��He�U��?9 �i�j0[�O��nZ@���
�G�-I:z��Q��>����e���?���i�&6�
�AJ(ѯ>:����$!�KC�������׊��g	߃G�deiG1ip�%�`�'a��'G��'�b�'0�|�Bߊ;����-�A��-)�[�X�ܴ>
��?A�����<y�iE�+Z������g@��#h�����M{c�iKv��2�I��*���#g0i*�LvN8���N�`��H�'٧��˓-�����S�f�
�ZM>�,OT�CT`F����i�-'i�����O��$�O\���Or���<�0�iVƘ��'.�s �ͳ6Yt\[C�
ѐ	��'U�6m*������D֦��۴2mWԅ��A/]��`���Ź88E@�A��<��&i%�2�
��B+O��IS��a �⚲z��a��MG� �m����O��$�O��D�O��$�OT#|�C�>T�֪�ל5RB��]y��'�6��S"�I��MK�y��F�i���z�)��TZ�x�1b	�8��Z�$`�4_�V�O�`�OS��y��O,��P��MO����×*��j����%4��L��䓤��O���O��d���%@�ʅ
w�h�Y�jPf�$�O��{ț6 ܽZ�"�'G��O2�X:*Xv sEA32�I��Z<"�	?�����Uq�4-:����O�[��#u���9�8X� P��RD�}�ա[=|u�	�?E�Ve]�lr�y$�L�� 
�<VA�3��~�< f_ڟ��I��`��П0%?E�'u�7���A��)�-�"!x��d��4p*�	��OP��ŦE�?y�Q�T+�4"��ث3��
��X�g+O��b��A�iM�7M��gH4��c5O��D��S���1��,)�ʓ;��S��M3A��BH�04�A(���$�Oj�D�Ob���O �d,rыT�{|����սW,���`��M�a/���?���?iM~���K�V:OD� F�܄L~��v΄�:�>yӦ.m�(�n��?9�OT�i���	�.8x�V:O�r�a�/w<(��Z�]�.@�K�O<�҇��g�u���?�$�<���?���F�J�� �K<L�j�[4�	"�?���?�����Eæy�~��	�T�b�V+�`��A_+]0�0�!XZ��F���$�M��i�r�ı|��(�n�J��м>���!���?��_�^�"s�_N�tY�)O&�	Ud0BdAk�|q7NRmc�����)s�V`�EB�O��$�O����O�}ڙ'�$a��< J�1g_�E��q��)���=��$E���?��V��-��)g�W��P)��o�fneӀmZa�R�{���I�"�d�'$@)GF�z�i�C�9�W�܂�����W��Ry��'C�'`�'trbJ>3rZ�A�� D������Ld�I�M�]��?��?�K~
��llC"��!���:d�o�l��Q��ߴc=��M�O4�N�����a�U6�|�j�OH�F�R%)p	��BpXǏ�<!�$�f���*��������� z�X����;9$[0�Ӷy~���O����O����O(�כ�d[=r�ˣM�9+qdU�p�����A�"pӊ�dR�O��l��M���'����U�7�MBтP�=vX4��*R�.�P���?)`�8�jD���E����J��]�pf |뱌]0!�,���2}���$�O����O���OL��7§M� Y9���g`�����J�L���ԟ �I�M�Ui���?���uś��d��L!D!��G��rZ@�l�V���d�>b�i�p7����9ׄӀ3��d�O��Qg��9	o��rl+G��[���g�bEâcK��0�=�����v���C�ȭ�bY{�K�$t����O��O¦Ab�� ��X��IC�����ԉ/�^���J���dYy��'��69O��b����I���-Bv����Ȱ|�~1�'IV�)�(�Bӓ���ӹwULAZ���N�;`�Z�I;	�>�(C�v�pɗ'�RR��'?�ec���C� Ȥ�C�� KQ�Ӧ7�8|�OpmM��|���?!lV�z`�q��οR���Ѹ�MK��&i
�@� �<y���`ى� S�}�h��'0����\%���P!տNsxhy2�|�'r�k�O"jl"��N.�4#`� {�<yt�i԰��yr������Ԝ�s�[D�X`T@�:����MÛ'����)�O�m	 /����%�t�0tcL��]*��Z)kk��$D+0l�� ��$[j��=�'�y���4�$!)��\�wL���B��?A+OܓO��oZ�Wtb���`!Vn����@2jeRe �p�YJ�I�Po�<A*On1RRX/hq�Bf).[t%�u�'*B$��w�5 @뗮����x=ZP֮D�,�	��h�4�X�9��da��@1��D�O���O��S�O��� fs
@�y>@8QM�]��Ap�'�*6�i#��D�Oh�nZf�����g��i�����`\1b�+����?���i��6�^Ħ�xCJU?h����������N�j���hI>+7��;PB)|�Z��bg��3��|BR�h��ꟈ��۟��	���� X*O�t0GQ�^4�P��_yBb~����<	����'�? ��4\��+f��0�P����Љ=J�I��M�¼i���d)�)�����q��(*R�#^"�="1e��
:�UC��#aZ�6�U�1N�/:��h)O>�)O�u�Vǖ�D���e���a�Ox�D�O��d�O��d�<q�iCz��P?Ob�[bo\�Tб��$�&f���W�'U�7�*�����ā����ܴ�b����!�J�%�(U�p��W�M�Ʈ	�<)��1'����͆�q.O�����߹x��եR����s��Q��t/�O^���O����O��$�O"|:�!3qD�4LO�s��E�D�_ԟ8��ߟ��ߴ�l����?ᆸi�1O�U�U��{z`�/�?z��4ʂ��O��XJ��+f�>�I^�'�*-�@<O�䌿X�d�'E?M�Jd��M���z񯋽^gX���)�$�<y���?����?!j�)N�0dY��˚0m���ˁ��?������]馵�h����IڟP�O�ؽ��-B2�1r��ғf}��p/O��'M�6�������'�jc��+��,!AG_�YY��\Ƙ�cរ;\��9$˾<!��H�$�VG�,���T�Q
��h�����;b/\�
���?�+O�$%��<�p�i�H�c#�ֶg�<�Rr�Ӏ/����(���y�?��Y����4	�c hd�){v���a��z�i8"6��;�|�)S4O��	6#����l���I�E���W��f��<�p�۫q�x��Ily��'���'�2�'�r�?u4�$���K�J5N5K��¦��ay�����$�SN��'�7�x�U�0O	W��+�1Yj� �bA2�Ħm	������������	 �Xr��i5r�XA��$%�8!ׄ�y,����E�p���kM��O��?��.�*�Av�!4t�J�b\�p�
�+��?1���?y-Oz�l���F�I�$�	�M,���[�i@����� ��?y�P�(Rߴ�5�ԟ4�O�LuQ%�P��W���;wTY���?��!�#e���$S�����
�*w��U���J^� ��,7�Թ����,b�@���O���Op��%ڧ�y�	"k�����,r�؝�S���?A'�i%]�e�'yB�v���<�ӻB)\�L��xd�#��:�"��	��M���i�>7��-�$J5Ov���'o&	�GL\ W.��*7�G13�F���/=:ˊ��	9��<I��?I��?y���?��Î�,���%�P�^=�aU<����u�A�k���I՟�&?�<wXX���*O�H��(�H�%6���"�O��n���M{��'�O��$�O},Q�C��%} ���W���-�Fi�c�
"���*�V���o
�;��|�b�P@��vy *7�~���ɋ�B�PMq�ź(��I�����ʟ���yyb�w�f�(�5O�I���� �l�.����O�UlP�*��M�eOټ�M��狭$ǀ��r��alYB"�;l
��e��<���"�D��cĸ&�p��(O����ߑzA���1|��J�%R4��BA��O����O*�D�O\�$�Ob#|J�,Z=(�� W�\01��P������	̟Ȼ�4�X��'��7?�,^T�cɂ([ʤ|�aH�bR����U}"/}ӺymZ�?�c/^�Q�j��0���r`�1��4s��dSCA�):�p�8Ђ'��&���'�r�'��'�pmP@��Gf��lק|�b��'Z�P��"�4L��9���?I���i����X����:	|U*fh9H�I������mA�4Dl����O��|r&�T)���
D�7[��ڦHϞp���ҡ�n���?���A�0��$�c��Y�W���AG �[�V��a�nZ蟐��ǟ���e�STy�*wӚ���E�0��FO$!�z��1 ��I3�Ms�b�>1�i�D�G��`�<�VcD��V�z��r�D�n��l9`1�l���	�[T�%�!P�K>��'j uk��N����-
\`%���'��I��X�����I��l�	D�D*��V_&�U*^H���@Sj�]��V�K��y2�'d����'�^7mp�T�ˉ5[��c��>{����������4,��_�����?���WͶ��G�u�8�EH���l�e�M�P�V�П�;a�υO���B�O�Ey��'�k��/�m�#��ri�e���O�NN��'}R�'"�I%�M��G�<��?I�-Ҥtch<�� ڪ}��Rs�ʦ��'�Z�$U��g�d���k�4$C�b:%`���
B�rY[� ���?Q��7)n�!(�>j�Ty,O����C��-��y��Y¼Ma�

:yvX�U�V��?���?���?)���y��RFn&J���O�� �ĸ7��O��mZ71t��I�9�4��'��$�޴e3�m��їLbPp$�Y�2't� oZ�M�g��0,���Γ�?^�� ��ʲ��`#N"/.ih��DP�L>y)O&�D�O �$�O����OD�RFѥy�A!!�b�V�P�>�剬�M��ڶ�?9��?a�'����OB�b�g݊^��A4���|����m�m}��eӈnڼ�?�M|��'�����@��0+@;C��y�HA6K�T��Td ���D@"w�����RB�<�O�ʓ0҆O&@�$��6b�:��(��?q���?���?Q(OT�l�P���ɂVy��xwH�x������	+f��I��MK�"�>�1�ig�6���� +��S��&~)�5B��;i#��2�=O���]�S� ���P�*ʓ�*�w׊$�e�"MS*(rB��8v��k���?���?����?����� �� ІG\�g�=}R���\�d�	
�MS�F��?��]$���$�>P�x�ɟ�@Lm
q��\�0���>оiz6����A����?{|���O�e��h�fC`%��-� H��9;p��/t��0d�V#j��O�˓�?����?��}��3�+�E��9G��"ײي��?*O�oZ�W��)�'�R�O��I�?�U�!n@c�X���'c��I���$�ɦ!JߴB������O�}1�H�<
��P�X��p���оj�|Ys� V���?�JR�Ǆ �|�$����c�8xJ4��-\�c9l�� 
�����	���ߟP&?��'��6mU�r�LE��Q,�&ā2�Ψ��`8���O��ަ��?�W�H2�4N��NM'>,.�s���xQ��ԑ�M;��M�|L2�ϓ�(��2�Q+%Q��&Ó!�?	�'<w�\H�ȟ�r��	cB�� B3x3�4��IӟT�I՟h���p��u�d�E?A�IJA��V��K�Z�c#�&� K+��'a��I����ϓoX��G��o۴qAmʡy@j��ܴA�����OF����'�z��B�(ϓa�ȱ���i�T�q����82bq���mA9�\E�4x�H>)(O6��O�At���Βgp�AFN���?��?���$�ݦ��'���t�I�x����"lx�DU�Vbd	�#��m��tz�	1�M�B�i�X�d�|��e��	X`��ቶtx�c���D�I�|��耗�E;U�.�'p���ؐ<�\���:O|����	|{͓�Cݵ �R��5�'�b�''��'��>��|��A��w[h͐r�]'	������M��.l~f��㟨��J����)\2�tH���9j�H���M��i5T7�'g�]rE;O�$��]hT�k��Z$N���.M�~�P8���aِ!�9��<a���?A���?A��?IR�	��K�����ч���Ӧ���Jh�@�	͟�%?�ɤb��0��)Ŷb]H�.!+��=z�O��lڭ�M�T�'͉OX�4�O���Ґ@55K 	{Q�!;�0�hI�N���R�X�FJ�4ϐ9D��R�	Sy�$M!NY��8��J�.^]��U�b�'���'���'@�	�M{���<1��G#s�R��G�q"��:�@�3�?	�i�O��'C(6�Φ=Z��=#�-��\T����Bϯ1}��w�U�	>�I͟�ӭO�-0=���]yr�O���.�??- �q���i쭡P(#7���'Y2�'���'2��M�	�� ܢ|<]��Ê?� ��O��Ė�Y���6?Y�i�1OjI���K�� �bA5zp� �u��O��F=�Hm�n�)�QX�r�1O��dF-y��+2j��.c$M ���[Q�y2&H�9��{3&?�d�<����?���?��-c�"�/��l�v,��d��?9����dYצ%�B�a��I����O�f��C�IW��A�*jƬDP-O
��'t�7M��������'���	J�s���0�D��ި�͒ ��͉b���*Ț+O���U�*D8!#��5W<�A0ǊG{�5��эI����O����O<��,���<��ia����9�D-��π?�p�4e�5��Dæ}��T�I<��D^��9�PH^�8��D��"n&�� J���M��i���B0ț	�y��'�t��a����Qx7U��
,h� �n��P��2I��]�d���<I��?����?����?�ʟdmk��ϳL!P=Q!Æu
���t�V���9O@���O�I�|ΓP|�&0�Ȍ����|U�d{P���G~mqQDj�Bhl��?��O��������;8�,��5O�dEM�?<- ��	!<K��a��O���&CJ
\� R�d%�d�<Q���?I��.%�<i��Q/[8���k@�?A���?���$̦���-w�L�	Ο0w!-̑����>�����*C̟&�ȮOJ�l��M+��'�哪#�~����=����^4	Ǡ��O������-h�]�K�<��'��u�7M��y���7]�i�����ɗ'0�?����?A���?���Iw�(�I�� ���;4Z� �E�O� n�Q�Z �����8PB�R)Q������,ɦI�O��l��MS��i�f��*�y��'1]hͻg`
�C�MI���p��"��r��'�	���I�p�	ß���XaF�CP�Ҹ���;�f�C��ĕ'� 6mšWOX���O��d=���O�lX!�t�@#��]�E|2�i�LKD}R`s�ZInچ�?�H|2���BfdɧZrм��� *�Ts��R(b����B�4��d�79�$Ȫu#4�~�O&�_�5 Nԝ3pDq�ʛ�P 
��?���?1��?i+Op�n�1(���p��%��֊"?5���Oj4��+�Mk�R��>i��i�P7�����:��B�%� �ėFQ*��J�R�6lX�?O*�D�+^��q��*B�<��ʓ����w�R����S(��Bd-%)�P����?I��?����?�����!��Fnʹ��N\`-�,�r�'%"�'��7��,Q�I��M��y�I�5yp��*��͊|�F�K���� �"W�d�ߴRL��O�� �N��y��'u:���c_u֢Y��B��#ej��$'��p���%�)9G�'��џ,��͟|��%?�Zݫ��7R<�CB�T�i;@�I��8�'��7�a��D�O��$1��џY@�K�;D@R|y�d�>�c�i^�6�쟄$>U�S�=d��2�;$�B);VC�?H�b�ړ�C�0�,�s��hyr�O���O�.o��'��hc�m�)|���׉Z� ��	��'�"�'���'��O��	��McW���	&B-C!��^0��ҠƗ8��H�'t6-(�	,��$����b#��7��ڒ%�*�j� 1���M���i�칂���3�y��'F�� 5g�
z���uT��!�̛YRX�#"�
*����wH�����'��'���'���'�3� ��;�"Q!� �IwN��L) �4�i�2$�������j�'A��:O�:�ɞ'�p�P�:D~�Tp�-f�8�m��?a�O������	��ؤ�5Ox�R+D4pT(����B�r�� n�OD�[$t9vy��I*�$�<���?Ic's&�*0�mѰ	���?	��?������¦�QFm��	ퟔ2���Gvдb�Ȧ�T�V���t'�TC�O��nZ�M��'��S�,w�=sq$�M�2�3��� �~��O��AHV�C�Q�c��<��'?Ob=q%�!�y�i�ܲ�ϔ>�196�l��	��@��֟�	f�O��D��W8�ʴ"��H��i٠C�&a�� i����C�4��'O��ŭD��|���]���Ǩ��Bhӈ o$�M+�Jʀ_/n�ϓ�?A�̶ ��4y��P"M�\ BM	 ��IE�Y�7vf��K>A-O����O0���O��$�OJ���\:�nX�"R�ϊ�P�O�<q�i��tY�O���6��hJ�SBfզ<bx�ç��%b��ڮOv<m5�M��'ىO ��O�	����s4v���M!2����-ر�����U���VL߄q񤔺�!SM�DyB#�QK ��Ѕ�:�0uzc��b�'u��'���'剱�M3��<q @�;SX����K	x�����?	 �iu�OTa�'Pp7m�ʦ�f��0#]	��p�!�-�z�[�f��3,���4S�d�P��� �Sy�O�<�΍�0�����c@�q���+f��y�b�'"�'�B�'�B�5���J�S�;�g�f:&���O��������G�|�I��M�y��H�
,�l�V�Ҥ.��`��&8
�R�tXݴz�v�O]��Y���%�y��'_��#̍d����GN�g��W��4f���ċ�.q�'d��ğ�	��I�{��Ęv�
p�^��Wf�&`w���Iğ�'��R��=&���ON�d3�d!��Tk�9i��&|%bŀYyR�>Iv�i$�7��&>��ӦR�ƹK�B�7�ֵ`�ނp!x+5�Y�r��H��Qy��O�9@�>J,�'�.���m` ��E�O�LiW�'f��'W2�'��O~�	7�M����'��I��7��D`�$ߋ���)��?i�iO�Ǫ�'w�7�̍b�&\��i
�1̰Ģ���7���m��M�@!� ����?�a!G,B�Rd�Rk�&��$B#�t:�.�3��|ۄB����<���?)��?���?�ϟB���y�Z�$cջ�V��!�f�< �d��Of��O��?	ٴ�y�nЩu�mZ�b�D�^����
=���jp�R���a}"�O���OhX�6����y��ϰe�z�(�	�;	�����`Z�6%H��:����8��'J�	����	#J~ɫe�"D���U�E(�Q����\��؟��'�@7�CCX��d�O��$US�tZ�B��~���K���!�t��+��Qc}��zӔl��?a,����cȏa@������p�@l�e�'�G�[�TSV�7f����?)���S [�ΓqA,���'Z(3��yEmG�PR�����	����p�O����.���@/Q���0d�"y��Hrg���*�4�?!K>��'�\�Ѱ/U�g�Bp˴�#X
�U��]͛Fe|�(!oZ�Ckf���*c���I+dtD�QP>~��@S *��LM.��d�a��l�U�{�Ry��'Z��'{"�'�"BGk��`锁99hi��*F��I*�MK@�f~r�'�����8��1ZC�BX!di�G{�4�"��pӺ��	f�S�?A�S�B�c�@J�M1��ȑ�փw~��$�0>Z��'"�yU�-=�0h��|BV�4��揩<��5��
�
;Uv�x�b�П��	ן���ܟp�	oy�`l�t8�s2Or-�A�����c�
�$±
�O�nu�?��ɠ�M[��iQ��DJ�G��=�0�r��_�* "�|p¥�A~�(5�������=��O:��τi����z�p�̔0i���'���'�r�'w�SLHB%`c�āb$P$�6I�|ي���OR�D�!㶪;?q԰i1O�Ց�M g�ڶ�ڳ7+N`ѧ(�O��ᛶ(b�&�)���E����W�ˤ.�<xR��'K���&+F�3清��#ł%נ�$���'4��'>��'D@(
�kA�l�pMf�^~l�$�'�RY��4!�ϓ�?����IE�I[�-�oB'R�Es��V��	���ę�����4!�����%,�Iu��	%G���҆ȜN��#�c�r�vP��R�4�ӽ}b��a��Q�=W�I���PH&��B�!a"��Ißt�I��,��b�Ry2kwӤ�9��M�d{��G��7np�J���z��	$�M����>ᦴi����}��@�h� 2 j7�����B��Hpd\�4�E*� �D�ϟ̱���AHB�I;8oXt�P�'�	����I�x�	�����H�TCG�p1����vQz"�㍖) �&��:�y��'H���'�n6Mm���iU�9YbuC�I�A ^�(A�Ŧ-X�4T�BS��%?��4D̒%��I� L�ڳ(���B�Z<)��d��m�*X�!/O�8�~�O(��?���k.���"�
H�uOL��R�����?A���?�(O��o4aW��Iğ��ɞ)HV1r�o�#��	R�&����Ic��(�����۴8BBT>%A��5.<!�� ���a"�B�OV��"x�0�Q��'T����b��y�HP��'���;�	�V�q�Nؽ; �}k��?����?����h��	�j�X<�@܅4��q�;������	���!?�b�i�O����*~�1�/�,-����شm}���צ%*�4d@�&/�!�0P	�O�k��v(y0��G�6���Rã(ʼ��R�V���O���?���?����?����� �	�璬okgJZq���zV�H��4Ҟ�ϓ�?�����<���+I�\���)F(L3�A�*0�I�MC�i���D&�'DRa������lH0�̍��I!	ɇO��+O@��,?J>,��"���<��`L4b�!q�_?�<�4c��?����?���?����$	��Y��
t��Y�g�7�K�:{h�(u��5m����P٦)�?a�V�P�ش7�v�O�	V���hB^X�R��>1�,��S1f�<)s�O>=X�Ή7z��a�%�I���SgIJL�'�'>,dy��O��$�O����OT���O�"|��%��g$�T�7a� ��tէO����I���شN�^��'~�7�/�I'2�b,�c��1 Jp	�QqPx�IB}R`f�0�oZ�?�o�$Zc�������'9�0A%cU�{,�)3�M!�l-bi�'�|�'�"�'!��'jM�q�2p�`4�c,M8sD�����'��X���޴n���̓�?Q����i׭B�2���I��e����B��~_�	��dͦ�kܴR�"�IS�t�Dhj���d]���p�7u{45;���rI�uS�X��=,�L��W�I=J �)�Wx;ܐ�A�.	!d-����$�	ğ���M�Wy� p�d��*�4X��̢��������,ŸO�F�$�OAnv���I�M'e��*�
���"�����p���~�x0��i�?!���O����V��+��<��Se�����"F\�Ӱ�ӧ�?a)O���O��$�Ot���O��')�Щ�há0�z�cu��y��9�4y�|(,O��D+���O��oZ�<i�GH�?߶e8GÑ>1��j�/J�M�B�i��d�>�����'�����<�0G�Wf`�����+d��ۗ@��?Qq�ڭ!�,��&=�䓠�$�O��$�(wh��DEk��4J2�?~�P�$�O��D�OH���%`XR�' ���/B���tn��[:�Q84�P���O04�'�t6�̦�x���ɗ�ꂢ#Of�%������'-Z��U(	a�ܠS[� ��?2.�����<���me�٫��&נ(�b�� �I���I� F��<OHIk�?S$LiV�T��'�j6mu+�F���Od�nZa���*�"C�Z�`9���ĿU `��J��?�g�i�6mզ�����՟H�BL0��a��'n�D�W�J	Gn�1�C_�u��%�8�'C��'o2�'���'ۮ��Gװ6�Cr�P=WsP���]��pش/�n����?�����?��H��D 8Q��*�	X�\"
ߞ���5�M�2�i@F�0ҧ0�ɚ6E�{tN�P�'X�jw�,Zw!U���,O���E�G8e�DѲ�>���<�狼m9詉UD�0NQ�6��*�?����?��?i���$Gɦa�������Ô(�8%�¤I[F���a�U����Ц��?Y�T����4v��v.�O��wG]B �A�ڬ{���R5k5.`)�On�iR�������%�I[�ߍ��cJ�H}�G��Xܕ[�C�O����O����O$�d�O�#|��R�A��urr�Y�g�4�@��Zڟ��I���޴\	VI�'6�6�6�ɥ`�`̹�GI�` |��!��-��P�I\}�*m�2�m�?�C��K�'���"��gD݊
�UH0C �rQ eݬ$d��Y�`_����d�O��d�O���`�����,�8+nB��&f0���O�ʓYo�Ċ$�y"�';�?%�B"�*F<e�磆�M�Mk���<�1Q��)ߴ����O"�n�	ЫPl�×A�h4�@��Z�|�l���� P_x��<���g!,)�1(ڒ��f�d�U�<uX@+�%*@�������?����?9�������Ħi�TZ:�Z�41�񚗋FJ��m����A�4��'���ߛ�����
g�ռ}������*i�h7-I�=x"ǒ�z�����v�Y�M�\�'(�iy��E�"��@��E�DX0<��ʂ�i�"[�d�I��$������I��4�OnB����NZ��I�j-L�tH��i�v1���'-�'v�O,2�}���ɲESF� Ķ>���jC�?��ܴqi�V��O���R�'���jM�'}��̓Q�D�u��|�vk��ܑ��L�M��Qi�-�X�AK>y)O����O
9��_�&�<�1N��`0U$�O^�$�ON�d�<���iYpٻWR�$�	*@"�X���K�l���B�&�^i�?�qT�X�۴8e�F��O�ʧX���Y��/d<�G�(X^��	̟dC�m�^��x��
@yB�O����a
(k���rɩWf%E1n�A�!P�o�'3��'M���<�%��	-p=*�i=<���Љ�ɟ`x�4��|���?)�ir�|��O�Q��I۬S���.�9 $Dԩ��'�"7-BȦ���4n&�aq��<���a��W��l���܅2K��tKv7 D��J����$�O����O����O�����
	��B#S�"�(��˓���锝�y��'R���'�*�#Ta��TD�V���p���K��>���iŶ6��ҟt&>���?)�E�F�؀��/���<ѩf@�IZ�Y�o�By���)4.���摲	a�'5�	V!|�HdnXpC� pգ�6�����ԟX�Iџ4�	��ĕ'|v7�K�~[�2$�Xs��H�!����1#G�HY
�D���?	b]���ڴLS��!�O���U�
�Z;���;"�D�zƁԹrr�R�OR���"�TA2���Q��g�&�J�,��e���Y�b�O����O���Oj��O�#|*叁4�\�q�n��7ip�������L�Iڟ`�۴!8���'�7m;�Is��8�5�^�n |��'�9N���	c}��yӘIo�?��P ��	���m�d�%c�4���Ba��X�j�y%Ѻ|�B	ܑ�����O.���O��D-� ޥ���l J���Ί8�p�@��'HRV��j�4*�����?����i^�&$��"��; ����f�&��I����Y妹)޴O��@..�1����K��V��
�cE��v4�x��V�(��&tp�0�f
A��& ��%����>H���3b�
��(�	����Iҟ��	u�SFyҮj���%iP�^D��a���^$`�r��	�M3�rJ�>�!�i#BUI��	Z*]�+,���Za�r�$4nZ�P�Da�$?�ш��K����UL ���>Q��$�3꒧-��Ä�3^�R^�H��������I�Ob�	dEāM��Y+d�T�dB��7�i����'�R�'���y"iӘ�I6?�(5AB�<���aC?d�мo�3�M[ �'��	r�M
���,���مHEk�4-�7/ֻi��`��O����J�d�j��N=��<Y��?11-��?x�ۤ��@\,���R�?���?i����DMۦ�[�}������`���M���
&&�%!`��zR�@��E�I��Mp�i����|�"hE�	��ا�N=.� i��Oay�b�*-o��U��6��O���H��6����~ߊ88p��H���a�����'�r�'[B���<	g�l=�� �@#z2�����`i޴1��'e�7-+���?ey'�TĐ�1����Z��k���ܴc��a�� �FP;��	r��Ȏ�ul��c #�<�{�+�0tV�4�n�I@y��'>��'/B�'�"�C}݈���ƅ���� �9Y��I��M�E�_�<����?�I~�;P�(˖������
ۂf��0�U���4P��F��O�"}"�N=r�l-��-
N.��g�҈˦�8���䚑��+�g�>�e�|\�X�q��&;O/�-��O̟���� ���T�IYyoq�ԌZ�7O���g��k�h�)��	�"�h�i���O�nMx⟤[�O��l�M#��'��a�8| uё�P�D8�%�J�u�'�	�1�>'�����^��U׉y	l�d��+W�J%� �'t2�'u��'a��'Z>řNU�M��k���K9��Ru��OZ�$�O��mڹ[h��	�([�4��'6��KV�]�9B���c���E�xT�w�'�I��M[v�i����Q�L�$�O������&������3-9x`3�����8�K)8�8�O�ʓ�?����?y��0����d��;6$5��n�8:�tQ���?Q+O��o��}j�	۟���_��cU��0���M��l��d`B���du}f��4l��?�����5�������sn���-�@��H��+�=	ͨ�a,OX���[�,$3�<���}^P�3L�l'��yӎH%
����O��$�O���/�I�<1��i�aժ�����M�YCm�m���D�ئ�?��V���޴hDB�B�	O��Hr�Qi�f%�i�Z6��0D�^�Ad���k���RC��y�+n��C?�BU ��b���v�R��?�+O��d�O��d�O:�$�O��y�����Q�2��Q�p�0ߴySDA��?1�����<	��i��S�Q��2����,�~|���x@P7-���������<�IT�:�"��O�A�U�	�P�3��W�*:�D���'x�x���	�pM��|�]�@��̟���n�d����de�+�R��K���	�����Ly£{Ӱq"p����	�}l�j3�R�Mu(�q#+X�v���?1qR�<�ڴR��V��OJ�'u:X[�h�d�`**W�%C�h�'u�-qC�
c
��q ������I�q�=O��8����-�$
��� nB�'�b�'A���<yd�Z:}�tl�E%��Q̦�#'B�Ɵp{ߴA���'�
7:���?A���·Pv��@矬<�f�;�l����ܴF^��Jo�
,0�WD	��!=n:�8���=��TÅ@X�E�*|��H�H,$�B�r��My��'H�'~r�'��$9k^�\��Ɉ ^H��H&o%�I��M��<!��?�L~Γz} $*C↎`\jAX$��.��wW��Q۴��V��O�"}
d̛:�T���$F�Na*��"��y^��R����$�\�~�Y���:U���O|ʓk��A�#�-rZ���,·>��8i,O*���Od�D�O�ʓ2ݛ&���yrdK�s
 "h�(s2d})#ŝ6��Ja�� �O$n� �Ms��''�<�J�,Y����)�,���!�L����'��1F��-�Z��0������ޜc*�&lPH IhI�O�4��`�'���'���'	��'>�Q�E�n� )�苽/ȴ|�f�OT���OԌo�6���|J�f��B� ]$�E �D�4˜7��D�>�B�i��6���U2d�B�8�I�C�T=s��\b29�u�J�E���� �zh�%SI�IsyB�'��'�r��:��䫆�Q�V�cѪ��V���'��	%�M�� ��<���?a͟��y���]
���с3F�����[��"�Ob$m��M#B�'f��W�8����C�E��UPEiH�f1*aQ�d��>p�I�?����C�7p�l$����[;��3 �A�f���!ǟ@��� ��ܟH%?!�'k(6�J$�`T����3�|8�AR����4��'l�$������0�dd�@�cn���1X�D7�@ڦ� �O���|�i�ZWb�33�ɟԡ �F$���J��dc�	��'m�	؟��	Ο��I�����H���F�*-�D�fiR;"7\)��G�'H�֠�J��	͟�%?��%�M��'8�M�r�X:X�Īr�e61Z4�i86M�㟘�'��Oj����̦�~��Y0y0`�X�� �w�%P3cF��?��Z/���Z��A������O\��3� �`*�*�?	����͛Y��M��'���'��_�,��4[�^Uj.O&�$V)f[$ ʷ.ǈ8�xɩtP�^��J�O�,oZ�M�5�'�T�P5��@%I���B[�
ʓ��,��ㅜS6bzK~j��̉Q2l"�'w��J�i�-^o�dY��>JUP�����?����?����h����L�����G�{X�)�������$�ܦy�U�K�������M����Owz,�%Nd4!�q�"BN�{��'�b7�K��U�ٴ2��=	�cQs~���5� �ґ"YȎ�	v�٧`9�h9��޲�P�v�|�\���矰�I�,���H{G&S���RaF
s�=8���oy"�g�r|�=Ov�$�O@����3|����F�'�Bl�e�N�*H�'��7-P릉��H����c^�3���I`�>h�t��r���V�����̦<�P
^�`	6���������*�L���M�4 L]9���c���O����O�D�O�˓cB�f�]��y�oϬN�zX�ŏ�4�8�C�.L����f���T�O��n���MC��'��qt��.�^��7��q�l�`Pi`u��'ΊY0p������e���M��8��d'F� 	�0h��I$l䰫$�'w��'���'��'>�x�V7n���LބEg� @gģ<A�`���.����-�<!Cա/5�r�E/R,Ȝ�֬̀�?�O:Hnڑ�M��' �T��T~r�H$BJ&D�7L�"�L叐(I_�=�#!�9V�l�)2�|2Q��	�$�IџD��b�= ޸�����[�����K럀��]ybedӊU��:O���O��'Nt�(x�
	u`E3Í�tnƹ�'���rߛ�Hu�&0��x��Yz���M�!�4�sC�ѡ5v���휟6J^�)B�Lby"�O���ѓ&��2��'�Ƙ�"�����)4�M�,�f!h#�'dB�' ��'��O2�3�M�cF��.�j�蝣cpz���-Ӯ?;�'`�6�7��2���[æe�[�0�p��Íрe��V��	mZ �MS���H���',|8!�BB�: 	ĝ?��͏9�8��K�i���"�O�ʓ�?!��?���?+O��V�@ ȹ�#F�?O(�E�ɟ�F79~~�	ޟ���V�i��D���labR��[�{gB�7	঱+����D<�)�*hDD��O��:U,Ҧ:a�@:��Юf�i3��'�"��⊏)Y/ %j��|�Z���Iȟ(�D$�N\,y���ƀ1|��Y1�˟D�	ϟp�ISy�"q����'��O����O&�i��ǲZ۠=�u�GE�C%�ɋ����A"ܴ3�]>�0��<i|��'>fƹ�U��<���zG4��������'q����n�2�y�F/�Q�c�8g:ᣱ#�?q���?����?����b��R�FD?�N݊Vh� `WB #��O20mڥ[E�	ȟ8�ݴ��'%��! �-�!��a�^����_�~eb�xӸ�l��M{��@��'"\���Ta
����&Ff]�eʘ�f팑(��u��'�����`�I���	ꟴ�I�i��jǀD1�M�<x1�'':7m��A��ʓ�?�H~j��V��U�(6���f�?��Gv}!i�.�lZ�?���#&�	�'Z5nj�Eh�5p<feD��v�W�L0�FYM  9�N>!+O�	!'M�L�Z��o��ip���O����O ��O��<IU�i�4�Q�8O4бeʇzٔP�RMȯd2�8��'��6;�ɔ���R¦��޴?���R�n"V�Ӆ#���|��N���x@Xb�c~�睡
��u���x��Og��n�)���R`�48����I�x��'*��'��'����u�kjz�0�D�C\��B�'~��'�b6��{F,���O��nZj̓VW.QR���4@��A��5r��a����R���|�ߊR%p��'RZ��5dT���sB��1rZ��S�_�{*���J^'��'y���d�	��H�	9`�VM{ׂAi��`�%�A~-�	��Ȕ'QZ6m07���$�O���-ږn���~ر�ר&�,,����^yҍ�>Y��i: 7�ğ���󊛀La�+d�J$,/B�:�K�=K�횷�ΪA�T�'S��A� ,����bnW���89rW��)rY!pnM�FVB䉤D�Ad�U/xB�٢�י-Ŋ#>Ag�H; � ���	7&V�ĺ��5C��SB��()���ҪK�gt��:��!? b\���'��T��fɫI��A����>�rq�Q�F�S~l�W�?x������zu�Z�S"�3r��=V����E�I���Q�,�R��e�QT(��[Jaw�-r��Z'�?�tM�~�hY:S���
��L��I�z�<ab�3��]��d�D0hvlt�'��E��dV�n�㲣H�?(����MZ�cT^
�aS�ȍI�'�6:�&�{3nEQP
ޝ~aZ3�"4b���tdX	?�-T!�,9B��B��G[��Ê����#��4*7Lܢ��K�pH�`L�3��=C2Bƨa��`�/	%�.��`-T�_�t��ŕ�Fɞ$W�[#�@|Z,AL^�'�|�'�]�`g2�6h���%i l��g�0~iB�'���'���'%�*ƹk��6m66 �vp���qJ�H�!�SΝ�IM���	���(�	ğ��ɒX�Pzql����D�	x����I���I����ɠy�N�aI|"�����A\7]j�q��y$F��H�����?���e������?���?a�O�@Ie��]��y��
(V�`���?��gb�"Ӱi����'����-n��2�]A%(��r'D%���'�RI	3n2�'���'$�O��m{BC4r�@
�b�>�0���Z5 $&	����I6�,^������u��I�\d�PG'q�0材a�r!��$�O�����g��C���O|���O��O��d�O��d�O� N�[�/�~gL`b��G� �rG�i
��D�O��{�ؑ'?��	��9[��л
����GкR���'��D���p=1B��A�E�OC�KCI��l�t�<���	�p&̓����35e��K&��y�`�8Q퀱�p@K7]O�h$�M�a nY����;ܤs�g��W�t���Ǻy"���^n؜��KbՐ|:��#���K��0���̬UD��B ꙲JF�<A@�L~���j��8M[0Py�fO"���bܜ�Ne��xR���+o/B�'F"�'���ȟ�nZq4��g�L� ,`�q�K<J	�c�i��) �!� ����X�W�im�@pI>YA�,$�8�Q0���\��yx�I]�)1�k2�4i�'(ҟ��a�OכFn^���[,���t��8�};�,ԛ1}j<���'*��3�'Z2k�S�,O��d�O7��,�dDG�@*)�%#�fO�z���ē�f�C)�5m$L1���KBh:щi�<do�@�i>U�SVyҥU�8�d��؎b��ӫ7ZN}��R<N8b�'���'�U�4�'\b9���xdg��{(=Q��O+_
��0 %x�0��0K�G ��C|��Pn�8C��<���5Y������d�я	r�(�*��WFʐ���2x��E��46!�&�X��(O��X �'7�Y{1���Ak��K4d�(.I�=�0�_�<I�����4��p� jy�!p�M[8��Gz�g�- �8(�r�@�v�"I�∬�~2�f�
�OD���i^�b��i�/a��i7���®9\�Ԑ"c�$7�	O�'QH�D���ʻ"W<��bc&D}r䌇.���S�%²Y�>�XƆ���?�C��=O`<�v�U]?.�hԣ�|�<��!��d�D �RC���uH���<�/C�(���x����EL�<��kT1��Ó&ǐ+6MYw�<)$��-��=��G�0
����k�w�<)���=�$TI!f��U�T��pL�q�<Y4*�9=R4�P�U6.�����e�<i�	5jQ�����Yx칉��Ib�<�E*A�i�4Y�Q'�4.&�Ts��X�<��#B�|w��1�ȏ��0I���a�<Q��s��E��U�6B�HV"�u�<Q2f�vz(���R	F	��j��J�<���):6d(�i� [[�]�RFE�<�a�\�W���LSPF���,A|�<	sN�5R�(@�,��~(%@%$v�<1'G�[�\(+�P�)���C'm�e�<I'�ɣ'�4��!G�[����� f�<!e�H<	�1!�]'D�Bqc�g�<���YlK��Et���Wj�<���`��m��/V]����'i�x�<#�\"HJS�1f�{D��@�<I�e#lY��D,��f��|�<��ȧ"���S �4�XL�Uv�<��q5�&�?�dD�FA˰0�qO�I��%8�3}B�iJ���6�*�.�6�33ҡ�#$J�AQr%�*�by�f@γS����$ؔ$T���	�|{Ԩ!Ǆ[�6��@h�2d�Ь��I9'���Ʀ��B��%�'���͔5u���"����uK+D�d��Q�~d0lSA`U���ȒQa�<ɐ- W;��C�F b#/]\7��R�'�Q�d�H�<�w���{�,����9j��ocF�2B=�~��ΠS,d][����{�_!+��T!d�G�
~4�Aʝ��?y���>A^�ܱ7��b�$��W�[�&�֭2aM~)͂��p>y6��.k�pE�PN�^��M����G�'pM�?|�
���d���2j�X8H��ۥ��,"�눆6�!��E{��-�j�
�Z֪Y,Yp�	�юp��@�1P�v麳B}�OX��&I�k����JwN��'<�`�Oa=eK3�ü60<���B���,��65F0�;�� ��g�x5�X��p�c�A����I��d�A ŌZ�4�&fE�%f衲
�/qY֜����bgPl��	$�ZP�B�8}90 ӕ��TŚ#?�
 ;#җ�	�fE�'dq���L�x�tҳ(��u��{Vk�s�<��ɍS�����<H��H�I�>�"Ϗ�4��i&�G O�Z\���	:m*�ԩ��ҺQ����4��>9!���\���F!Ҭ
�V)���Z�-�5.P~?чʁ�s=�J~�=� �kqg�<}���l_#�h*r�'6�K!�W.]k���N�}�*�.I�=p���ƍ<3�u�'�\��������Q��!$#� �ե_j�|���Uk 51Q�X//���]<�		�2eϺ�i���'ɔ)3�%�s�t��D�u�$U�E�V?=X���@MZ&t��~x�xc��Z�M�d�[��L��B#�$��>I�YS���:i��yu"�y".��U�Lq��dz��Qa��M�O��	CH�Z��EH�Oʸ�夘�U`t+Ŭ�;L����"OP"�j����<�~�������'<�䒊���MJYlX8�,�>\R��#('D�<��
����a�h��X�.i�5 Q�N��$ca�'f�D{���jR�"���>p�l� 9SL<��#̰1�rYY��OaA�P�! GY�<����R��;5׷5� �¯W^�<���:�P�F�4��ɀ�-�F�<��	��Xb���])�PI���e�<�1b���(#�@�"��mᆃ�\�<)��le �JF=B�25��Z^�<��L���$-)ѥ��J��8`oPT�<���(j��d��V�e!�p���EV�<iPM M!T�+*֑=�8B�I�<Q�N�"�D0��,�f- IA��H�<q��93]�4�б.�^�����E�<����, &H�a�x&�5P�,X�<�ъòscP�n�P�� nT�<�S��/D�yY67-}YC�Q�<!F̟�9 �̘2;$t�X��H�<Q�`K<A1VT	�B$���s(\}�<�&�; 3���%G(b80�mR\�<AC�3M߀�c7F��yzG��d�<1�%J�M�3N5 ��p
t�Tf�<q��I_Zf52��F�`�\ Jr�o�<'��"��)���,q�
��4�i�<9��׍<@�y��(<�A���f�<��۔_?	��ǜT�戡��U\�<�$��Y��Ȣ'ǈ��@�梃X�<���J���2�d�9&�B���VW�<Y�NX��D6����*U�W��e�<��(	}�4�b+ڛ&`�q��g�<q��U$��IP͈;:�x��Da�<�4#RX�����;#N��S��J�<�0�U�v
�)�n����I���G�<���G2}�z@Ƅ�y6^��&��B�<a�m,��  ��/w��-���OF�<���ԃ1����7!�1.���H�<A@I�T:l��A�/\U�y(�`HR�<�`�)8Z��U�*0�� �S�<�����0�P�8���Z����na�<���(���w�ٝ%����GW�<Q�@/>�P [�PYJ��P�ȓ!xZ��Q�\�Ju^�
�%�c�݄�(�m����2���Wl�V,@��ȓu�r4���
Wh�
gg��[t��ȓ;W��J'jK���*��S����"O���G�v��31+�2�h��"O0`�t��Tt�!��;e���"O���ͧc�]I��Ȯc�]�"O��˥�� E"���A	Mڴ]S�"O*16d�1zk6�{6����$p�"Ol�c�-�w���F��:�≱�"Of�jV�Ì7 �� -���
��0"O�S��S<A-��( -�5*bBe"O�PF	/���K�LR�p	���"O` G`�"�lI)r�$#Br��d"O� �arǛ����Ѡ�?=�-��"O�m�6�H�-��h����^B�u� "O����HH(3P���؋q9��r"O���A��>�A��j�;)rҸ�"O`b�&��:�8����-}5J�"O:��I��3�+�	6�d"O����ɾq�4�c�؏N����"O�ڂ��W���ӏ�j&���"O�X�1#��#�R� �N�5W�͹�"O�5���М9������E��h�"O�|`�]�$2�y�n�><��`"O��Ђ?����B0\z,�A"O8���� l�P�k�#w��ъ0"O$�*���o�hɳ��z^��"O�M���28�b��d2>(v�f"O�X
��14��Q�#е�
0x�"OĀ�&��4#�x������NH�#"O�h��:o�(�Re��,��"O�3�V�"�(��c��� ��y"O����戊lx�"X(�b"O��iV';[�P�࡞�i� ��"O�T��*�-?����PrJ�
c"O���%��}��8ِ�N�b�ΤS�"OBZ��D�<���Ã��=Y`<�%"OT�5��34��m�Rt��"O����Nח��#�[O���w"O�)�$�Y$h�B�� %��RT>�H�"ObA��68�p�{"�ȯ}OZ�@"O^	s��/%�81�bۤ$�̙"O.�	���Q��T@��	
l,�]�W"O�QWҁB'b!���/"v��g"O=Ӈ �n���־f궜zC"O`-2㣀9{**=+#ʊ )�t,3"O��� ��h�h�sC��p��3�"OR�؄BN�0�r�)A��=f��#"OB�r3b��,����rB�NmB؋�"O�a����.LrH�!H��t���"O�;�`K�v V5�"�
يђ"OT�"���
L��5���!Z��M)�"O��gÈ�uZ�i�	Ʈ�1"O�T0e+���8K�!N�&�8�5"O�X�A:N��l�� B��$A�S"O�uxq�_! ͖xJ�o\ 5:�(4"O���@Ӟ[MА�OծmN �b"O��:BNZetB��4/�����"Or����$bYT��#��ǌ�a"O2���"�"�0EȀm��o��%��"O:	��M��3�H��C� �0-* "O4�:UG�<��Ο�t`Dq"�"O�)+q��*r5�ፕ=ob�!"O���KGr��)1��IU\IH%"O|<�p�؀&����^-	Y��"O���D(,M�a��-�a�*43"O�a�Z9:4$[0�´���%"O�E ��-Eo&��̄
E�U�"O�X��!�f}��6 ��D}�pP"O�)T��c��8��)�Gv&D8!"O@ Rj?T��5ұ�[)Wx��3"OPp���0Ry�pbV�Gb��(r"OJ�I��ē	~ݐ'a�w��Zr"O*ӂ�@*a�X�b�
'�*%	"O^XP���2]�i�Gў	74 ��"O����)��d�@���ݠ]sD��B�'#R`)��'g̡�b�S���<!�ҺJ,��;
��� >e���ь-U���ӆQ B�6%s�"O�L��t�z#b����4�d"Ol�Q���l6@H�9e�Ꝁ�"O��+f��;���T�O?cD�h��"O|x�a�O.4�z ��
?7���&"Oh��0� <쑃��0DL��"O�)adG6""P�є��*]3��R"O��A���+[-� ��	[z�"O������X�1mOF�9��"O$@; -�M�Z��,D$,��Ӏ"Oݒ��ʞ_��Q�(6����"O���瑹q��hfm�+	��"O�l�Kֆ.�|%yF\�S��"OD�{&nͨd�a�A��
32���b"ON�(D'H�b���j	�;1�h2"O̼h⬚<Z�F�2�֙K�@"O:Z!�4& �)�&�X! J��"O�����$P��RCAK)����"O��6|�C��/�^��"O\wk�
"���p�L>+ej�jT"O��h�X?g�rp��$GOV��"O:�K�KD�\4j���n�3"O�[r%X�8�#ƮJ9Fƕ��I9"X�9#q�N�e�蓄�*	7��L�% 4��C�W�8�6��!��;\���C4	Y��x��@�!��E�0�
a�y�^����9F!��:������֯F��DC�.(!��!sz��I	K�2�!��:�!�DC4��b7OVصS�+H,�!�D��X��������&�Z��C�{V!�dX�����ȕ<T\��d�L.!��:j$�{&Ȑ�5�� ����ru!�ղo�$�SOD�I.(B���>)!�΄wH�t(`���l�P3.���!򤘙>�� ^	���(�X
!�$йo�=����	���P�)0M!�D�3ʰ�7+߂+2|�P6!ŵ>>!�Ď�y۠@�O��B�A�#Y!��ߩP8(#�l�3��%����tr!�$�&S�x`�əf�l]SbA�D�!�D��m{di��D;4�L���5r�!��N� Ȍt��*��ժ�A��G!5!�Vz���3g�I(��P@(!�䛊<�pJa�	� A�!�u!򤃩!��qiEN/{͖ qsCJ7!��%_��Y����=|�"v�ҿU!�dܙ&�1�O�����L)�!�$F.tb����� �D(U��:A�!򄛍d$(�SiC;y�N�c�ۢJ�!��G��m��GD�o��y�PfJ	�!�D۫[V�Z�E��:v8��!�L� �!�AwX�%9(2o ����#oj!�ć6_Cڅ��fU�Of~�Z�;i!�ؚn�%p�U
T�A�[�Z�!�ҊI�0y˔j�,&����l�7uG!�d˘xf��SK�=d�� ���Q0!��*���k�&O�@���'C\�d!�D� F|"A�ǫ�K5�,ӱ��;A!��mtn�٢ �?"�`�(U���&E`���;����C�z7�m�	�N�`���*-��ZY �!5b�zE��"O���d��Zؔ��B�0�@�у�	�>�&I��EI1^l�@!���O<؉�J�[��D�8I�k%GQ�?�n��$�	�a���w�%���73s��$�.A@�;��_2�.}05�!��� �ΐs/�$��	 a�`p�gQt���sI�[;�"?		�^K�9�ţ_�+����'�p�� ���n�j��Q��Z��B�K<a ��
��5���s�
�~�f)p�l�R�f�'|zT���	�-,�(�sh�7?���ƣO�� %>X�e��.�y �Q$)�×*O�uzC$*�Doh�!��gF�w��� $9O���J �x�1�1OX4C�����{0L)7��k6O�5@�eE�zٓ��"��Ň.����硏90�*6�'�,Ɂ�	 A6$
rGͺ�TܑÓ(��	�'�H�[������<�����c�L�G�_R7 �Ed�~�<s�B$R�l58��j ���){y��W�( �b̗Ll�ݡ�BD���e��qc�yvjټ]y�C�
8��B�wb���ᇴpd���+�dz���ݾ�~I1L>���L,l~�E�=rϢ8��j�@��\P�Ν�%V>B���Q�̟X����p�� �b��'�K�\�a|r!؞K�q:tK"q�.yI�����O.�Q���	Ķ�-D�f�8.�|�R僢ɒ����ΦNNFB�(pE&m��|%�� ��r�,ʓ�d]�Ē"Hv�ҧ(���kf	IH�R�H2k[�BԦ�2"O1��`͂$w��`���C��kU' s���l�<0Ӣ>��$
�C��3�B>egl��N�B��'�Gæ�`��	�^��i��[�fPRPo�*ʚх���qØ�!��:g��ӶG��?a� kk�8�D+�IH>?��h�r��_P��R�,��,�!��9�8)�
W*Z� !�
N��/O^�HA�$B�L��|"P�N'C���(�k�53HU�$��j�<$F�/
�"��:g��ey��Q ��5N���[���gܓ0���{gM�m�]���F,٤,��ɒp��	T*��B�@��T([�&Q� �� %R�+��'�����5��}D�U!��D�0��U��i =��'��"�"�� X�y�	^3h�pT��%�T$��_#s�}iQ�ĊH��'̴q�U�S�
!�OQ>����� �B�{B�� �VM(D����G �@���G N����˙��	 N �����w�3�ɇ]4|0v*�Th�Y	fko���dȧ�|	hGB��ê��"��:� �9����6�4	��2S��j(�sX=�C`���Gң���@b�a��)1��W��]��ځkZ-2^rC�0y'���cF cc � 6�X>?�4˓Y���
ȼ#y�ӧ(�6�2�쌘+<$�	��֖^Œ�"�"O��A�j�����(F% �IK�Q��N}��Z 6���p�;��$�="b�XÀӶ�����U�o���$�b�b��a/�+�f�P�_<L�I��*�8\vR���Ƀlj01ʙ�F�0�!ů��?��D�'��Ĩ2�	ͶDʔ�Z� �"�6$pBC4PW!�dM�L���*��ʕ`_W��n+,9I�#G�=��S�Ox��׋P�!�B ����u1�M�	�'l��p��w��M@A��@#Э�..}��] F�Y%���{���g��$�-�Gm�Y(g���x���'�fH����!#�d�7+,�qe`֡4�����Z��%�K�(6uֽ;v�ǫ��Oh��̇m#��[K|�4!�;��RQa�f��v	�w�<�Q�K�Ga$���2G���kF
�sy2$^�H|�ӧ	I��ӳG�<�뒋�-ÔtP���,XC�ɾJ�����%up9k�kB1o�d�H��p��Ǥ"^h�&?� b`�ƶ\��A1���};�cm6�Of `d�� T7n��o̒m2!���L5!	d	@q�։��?YF[f�A� :,����d�'�l���G�`hX�&>%�#BD�Qn�r��\)V�|�֭-D�,c@�'E�(0��^*��'�<I���:\vy���6}��\$����D��8�.u��!��$L�ĉ�#�����MT:�O�p($��qO4�{�!�7d����環��x��'4�y���E�q85���|q���UJ�Jvz@[P�g؟б�o�*e�����ϟd��Q��2��!+t��V�2~������H�ZQ�y�KF�6|��""O� �1�ꅌ�N��f��_Nqq����H��
�C>2�$�"|"朁A�$�+�L
07x>H6�z�<��!�c�a���Q�+����L��i��N�aۧÉ��g����zg��r(����7������B���i�~�����6,\b��2�ު>���'���HPk�)���j�+xFp���$Q�9�^�:#����'f��D(uj�XŌ-qb��_�y��4��="s�D�]��O�6f'$9�'�{rE�Z���OQ>�iE� ��U��:v�Ĝ�s(D��B���.����3[��};�b���3'6���r��N�3�	�&5�Q�W@ N��u�@N�M"��$�f���!��&3�8��P��/Qr���=
�`0�nL���DW����r�J<:��GR'�3�r�8��J�ӵl��YB�a
6?�X�d4��C�I�$�dA`�!�$j	y���97��ʓ\�$b�I�_g�ӧ(�$p�dnؘ>󌭡V*��
�/N��y���x;�0ze\�;E(���3cX��'�	�T�ӕ'F�ϸ'�&�2�˒]�La�-4h���1c&�0�O܅l����3iB�sp�"��=z�\�r�.�O�iH5�^�2�j�"⍁>=�9P`��:���A��Fz�O�	S�l��zv՝C��1
�'��D{���)�~�P%_���؉.Ot!��S�<��	N��|�2�9X�� @���o��[��p�<񶫏'/�������"�ѡ �"/;�l�D��GI��g�zCB�x7F#�V���^<7ḃ��:�B��
!KiJe#�ƴ[o
5�w��q* ���'s����JO����5��'~ b��d�j�<��6ǐ��'!��!��BTx���n̍V����^�����+_�� E��0'{�ܖ'.�|��oC��OQ>y�%g�*�م�� fZ�S�#2D�<�4?nX���U2�nArQ�£��A�'.���q��J��ϸ'��m0pP6e�i8�<���r�_�l2�aJ26��d���٪ֈ��B��%a'HN�Q�6��Z1>tQ;�� ���aC�4hџh�A�D� �y�nЧM)ҡϧ(�J��'��0���I��H�&PBd��c��²�A�����l�p�̕'������1��,94�%*:?���$��N��t�/ʉ	�ha�J-D��(d��(=HQ*�Q]y�%�ůB�&A���O��-���\��qOb��怀R �p�%C�$�¡���'b���hR���9�CȌ8�, 'mݹF�&�{%`��̉���b؞ �g�\4��}2E	!a�p]yG('��2Q�A��D4e�h�q��\���+�

�,�HPo�ee\̀U���y�
R�'v!� �YS<����/��d |�dlt`�,+?��P�թHQ>-ie�.*"�)U�����,D��kѬO�6^��'eE$��qY2+��VM��j�-�*?�VE�B	�a;�qO��"��!t�D�Ti^(R=
<а�'+��&'	�:����w��6$T!H$� �'��Q��G��<��hAH��p=�5��~��1�+	9ݤq�`@n�'�����Ν�`��u��)�!8n�k4H75'F�Hw
K!�F�b��I0�!�+cv498�R:)����+�t��	i��Yd����@!�=��>�ȧ�\�(��&$��r��4�&7D�8�3ꚇ<OP���ؠ�D�y7��3}#�x���ߟXAĸ7��c>c�p���;$�.uQ��:|�2���i=���p��6@�ajE�m&|����g��m���Ġ��b�7|O�����n�)���*���u"O�AT`�jnI2U)��k>f@2R"O�4����_�hh���l<��"O�=��
�|�zt�d��T9��"O�Bg>��H{S�R�xكd"O�5��D�?d8 ��F%|ӈ�H�"O<=�gk��MZ��B���CZX<:�"O�	 �,
/E�`�b�B�|B	u"O��{�)T1��]:V��vA6`[g"O�[���zbt@�����	<���@"O� /ŋF�txG�6��9�"OD$:�& "s���jc W�� "O�y��d!�U+��?q4{�"O6�[�!��ӞeZ �a� h��"O��p�N�I�����X�1)�"O��5&޹F�.�J�.؜<����"O ��jO$]`pq�˩����"O��P��,�UOT3.d�BA�X�<Yvk�NH�e._.p
5 M�<��aV&��̡'�*&bؔu�J�<Q��x?�a`񮉪}Ё�!�G�<���@=M�0"���#Z���@e�^�<�a�ޛ2�z�ࢄ
�w�L	�F�]�<q`�֐�ne `*��F�r���\�<�"�7��2��_�N/2MZ��o�<I�gЪ#ތ���E�&�)ڕ�Ml�<dƝO?����7Ia�&Ml�<��+���*-����?3�p�jN`�<���r�x�P�&�:V��%k�]�<�Շ���8�xT�^��L��mZ�<a��;O��H�aDt_�+�PW�<9�dŗF���ȕ�8�M�@�P�<Y�FS�%g�P gFFz1��K�<�g�Q�ɻ%
�+�����F�<Y�c��0|B /��`�R@E�l�<����2:	r ��3FoTuk�/Vd�<�f�:|,:Ԍ֯yڀ� e�<�fgK�d�~S��0s�@�ɏW�<&A�:�X`�c�P0HUN��!�G�<��j_�_~�Dq4"�*���'��J�<�NI�!�&y�RE��1���!�G^�<Ɂ�'����Р�q���$�]�<A�]�bU��#�Ts�0���[�<a�e� ��}�FK�.��d�$_�<�Рy8=�Q	ώf�f���
�V�<1�D�X(�꓍�b��E��h�<1���"��ŋ'���-"�8�-�Z�<ٷ�!/H���J�**|�8"�X�<��S�T�$�s�ی3�d`�ϕW�<����������D�����AH�<�0��$0�P��U�^#�����D�<y���(!����5e��9�ϓF�<)1�;��}�C��3`��Ai�
�^�<�g[:�Ѱf߫#�A�XQ�<��c��Z!{�$8m����H�f�<ՇQ&"���3���{����ǧ@W�<	�J�$�d�sU-Q!��L�rIV�<s�
v��� JL�j�D��b̛P�<���>x4����^�mɮ �6�S�<9#�/Pe�����Y�oo�cD��L�<�VcM>gt��0��y_T���Ld�<A�l� )֨�0j��i��`��f�b�<�G�T�$p�R?>8����v�<�:}�X\�a������C�ɞT�`C��G�Z�rq�1�M �PC�I/�Dq���,q��Xh�+O#/�C�	>?A�YAUdT�"�L�2��>�C��"F��ԣ�D��LQh k�C�Ʌ0ǰE��.ڔ/dt2�+O j�&C�-
�m�d+G�����P.{a�C�I%|�� ��!Ӛ���S��t�C�I�%t^h��=z�T�6��qXTC䉚>!�	H�@� <ώ(3�e؂K?D�h�5*��[^ȺÇ[�V}�dHt�;D�� l8X&
�0H�TM�&��B�U8��+U^�flͣ��K#a v!"��#D�1��L�Zr�ئ�H�{c�@�D"D��c�G1|��5�h� 7���F5D��[D�":�5�P.6hf����)/D�$bS�������%�\(~H~�#��8D��SU�])re�t�q$�nP��bp�+D���Dm�0^���!�>>D���.D��R6A�H�!M�_ڸ���+D����B��'�R!:�+�;Z�~�[�!'D��f �;W�V}���H��h��($D��rF��Ut����3�H���,"D�,��KGe'ġ""n�;�&ٙ�@>D��ң��U1�y���>iG&�,)D�x���QF@�r��ԅ~n�0�0�&D���GMG5��2�W*��5�(D���,��s�f|!&`Թc�J��I3D��)ƫҼ����4H؈nIJlR�D3D����g�(b���!����Ѧ�y���Q���K �FNi���aΌ�yB�X�r��h�/P�/��a�B,I��y�ʀ���K��3`�ꧪ�=�yҮ$ �8�c,��*��h�g�_$�y��ف�<ؠ��<��8�v�X��yrAX�:F��DO�!������'�y�i�o�8� "C̑!xf\�"���y��F�^.�rF�]
-VNP����y�!Զ69�d���
�2M2F[��y2d¾?_��q�U.ɴ!�f���y2,��"��yFd�y3$42a
��y�	�
cb�u�կ��l��p�y�mڜT�-�@�By�Gɘy��ȓ)?0�B�M��0Ĥ������~\��tk2󯚄1(�=�Ň5܆ȓ}�ؼ��(���~�:�ڮ1ȓ~�Zh���)s�p�4�ŀ2Κh�ȓ#��Yz�ل<;�dJ4�B;2�6=��sF��{1��-A^4P�"%ΎV�pT���p���,�:Ǆ���6ODx�ȓjX��Y �n�x� ��\��KPq��U?v��\�R݆_~�	�ȓ>��j�e�#a��s�I?r츅�:X��i�N]�14��E��Z�D��ȓ%�A"8KBNx:S'[J�ȓI�]䐢d���i��[�!KR��,0�cӇ�23���D�j��5�ȓ�	R��'�ڜ��ψ#r^l�ȓw����%
�i�B�+�L��B�z%�ȓXȶl���_�J�	ဖ(90��ȓh�P4c��)D�^	�%��Kb��aq,�i�ʙ�%F@q;�,�:X���ȓ)y,�5L�9'���1a�":gL���(��YK6���`���F�2:ڨ��dI�U8�H"|�&�
��LB�	��Mj�D��GVvt"2/[1�@B�Iu���e��$W�fx�㖘7�C�I9S3D���� ������l�B��~v�ah�	Jr%*�j� )B�ɡ�H��D%/	pE�c�	|2�C�I�Bx4(�O[����SDD#��C�Ɋo7���R$F�3 	N�L�^�rD"OmC�
���p���'I��y@A"O��CS�Rd��G��D�0�6"O@����׺$�\�B�_�=�b킑"O� Ze���`�D���Z�p�|�k"Ol�Yt��h�a�$J�"ujƐj�"O�y�L)?n^=S���'SD�"O��3��åQ�MP��ͭ8�BA4"Ox��CMO;:a�pS���! -�y�?��5�Wߕ"�����yr��L���A�DZ���	��y"f�~�b���%:�>壧ă��y�ț�W�hyS$�[�+����W���yb,�-(L}���="�)[����yr5e?���]Q0-`�.�yR&��u3��C��0[",J�����y�
�#V�|���?�I�5(��yR�M\�*�����F�[b��
�'���p%ȒA��KU�����@ �'��	M�282�� !vYN|��'��죰B��y$*��&W#tP����'�z�X��ӯ`���Ҧ8����'���9���2ʄP0b#T�3V�P�'r31^��[� ί%�xP2�'#���䠎�H�ԩ� �֘L����'��=����{�\kPb��:���'�
�ҧ�^%Z8�=`�+0�`���'�<�(�@Z�k�0)�(:��y� #D��STHߒ#�d )!j��KtFt��(>D�ػeށ[�xxJ��B[4�q��;D�`;���G�`� 0��&x�na���9D��V���Z~:�rĢ�'ILx���k9D�p@�
�E&�z!E_���ID�)D���F���,<dQ˕/���jxS)&D��5K?8���ꇽH�<,���"D���b��J49���
H�89C�2D��2� ?l��Lp��_0��I��2D�rEO�Ec��_d�H
��&D�p	Ο�o���դ�F���'�$D��REꐉR[��M��h�4I��!D�������.�2T�� �F�,=s��-D�)���<�d�ɘCB\���'D�HyB�0x���$�)0Y\(�1�$D��JB)��xͨ1��z�\�c%!D�T��˝Su��z��$9EX���3D��['h�"����6Z�&�#�#D����O�-*���$�^qC=x��!D���#���U���po[��@���>D�I����W>LE�P�ď+E��a�8D���'ā7 � �� G�����F:D�Xp�N֫V^�1v�ʢ8�xHكK-D��#b�:Pʾ�2֤	4�ZX���-D�Hr�$��.wdHV˒����A�.D����a���Rv�L44AP!%:D��9�!�{1�H�h=~��:��9D�����U�K	J ]��AڰN9D������>����	 �L���N+D�T5dKn��Y��*B�9����Ĥ;D����)p�$0Ip%V0*�dy{N;D� `�`ѳAc�y@�ԓ�2���9D����eə2G�tQ��W+���1�1D�l!���7aCZ�@�-m!�]´�<D�HI��޼`޼��ī'x�)�9D�8�V�C9g���ĝh�4\��$D� R���W8���áHN^��7@&D�ТU�٪D�Т���NO�tBs/8D�8��*D?��sd�_*@�\��,3D�@�lР 5l g�GR$ �֊1D�� $�"�d#(TD� !: * "O$��N[?;[��x�(ы	�%0F"O8��梜s��x3j @� �؀"O��Gi�2J*Hx�
G��9��"OLl���	d¾aB�� ���"O@Y�ۤc|��gċ9*UV"Oбp1d�3��P{RF٠x�З��y�
G=.U�1���,,�M�����y� �Y� ���n�x����g��yr�X�m���1���w� !@&��y��ɱH���#�p��PB���y�@ <l���m�;q��Z���y�%I�-z8!�*A�b��<�ҮU��yk�BTܘ{ìL2b��!*̀��y��� �u	R��*`��򁋙��yR�A6��[�����ll@�b��y�B�pTzDҳ	���2C�2�yr�
d�12E$�a��"����y2`��\l���@Mj��ӭ���yr�Q$t��|"#��$��IYc-E��y�D���S�I7T�ܱq�d��y2�Ͼah^1�f��S]D0�M�.�y�� Wt]ZG F� �g��y2OB >��DhD�,f���7�y���,�^� ��
�NtKG��)�y҆��d���rdAqs&�F�y�)"`��x��
q����^�yb�X+x|��S�qr��(�ҍ�ȓ�^� �Y�Zu2��V̂$J�:H�ȓ~3�D��a�	: �AԎӢd����cH���(�?n ����_5L'8d�ȓf�D�6�C�9d�U�E�
�Te��X��iD2J>�U�r�M����ȓB���3�A΅!�F�7&�=�2̆�P`z0($P"6X�ɱ��Е�0m�ȓ\���hE

��YD#N<�ȓqH� �換8n�~�0熗%>�Յ�NK�)�� �9�(�x5o�J��=��C�"�jλ|�6�q��s�b�ȓ89-�S�].fɮJ��+�9�ȓln�!%�:�TT�W �>l�N��ȓE�,-+�)�f��h��c�"����j) 8��$<��`RR�	 ��pF��w+�<3�2�A�7?fRM�ȓ)ơ
�e�ʤ|qƇ˷�.��ȓ��jCKg��%!�+T3|��݇�B�10I׀;�>�@1G��b��ȓ_�HB�E6�`�,�3�Յ�F�)��톧�)7}��3�)O[�<�1G�t �@CQ�}�v!�wDS|�<AQ��`�4+ǋ�:�ta���M�<Ყ��&�J z�=lqt�k�fM�<Q S�C\�4M�ԌTk�e�n�<	�jKE&����V"���Ddg�<�E�0^(���'��	3���M�<i�CSAŨd��_\���r��K�<�bƎQ`P���Tx�x<*&MPn�<����+��膧F�+:��u��i�<��&٥FZ�<8�%��1ሼ2Lg�<ѣj�7�XIP�F�;f��$;'l�f�<� ��3`-p��#H4(3���4ːM�<9!��Q��M�aM;5��lk�!~�<I7M��#��<xa� 4Ȳ5aR{�<1���2{�D�e��0�0'Jn�<� �ma7`T*\�z�X�E�7>>̘��"O�%�eř�X�B5�D�Nt1�"O�!��:+>0K��m���f"O6�:��\6���*�(�G"O��k���8��$� ��8uv`%�E"OD�qE� 43h��{��	}.��"O�%�d�7�����<����܈6�ў"~Γw\ʹ(sJՠd�("�hN}��7�:P*�n��#)l�#W,SX��Єȓ�D��"�!4<�3�Gߏ#�$��K�Π�t�'�J��Y�-���ȓ`rF\�K�9(P0Kj�|�ȓT�^Y��)Z,Fj�
���YlM�����Y�>al��zsQ�2��ȓA�H���r�&d�R$�1J���ȓ,yb���F���!�`
q�ȓc(�LJp(�I�q�`�R��ȓJ��쁠K�,f�@��Əv^�P���DD)4��pc`��[��L��ȓ�A�����i��1�vI �>Q�ȓZҝ�� �Y�6�a�-9�\��;<���$�1M���� �W�ވ�ȓJ!jax�.����B%��|�`�ȓS���@!,l@ֵ�Bd ,���)�Rw�7%�����W�F�.M�ȓjCR=������i3,���,��0;�52�@ Zu���ƪ�l�F���Ko(��d�A�iqw��-=lP��ȓC�:A��J��ؘ��1��ц�y��H	�DD�3�B�Q��w����A��#�J�
��X	YBVX��=D��8"���}�3�ղ,w��K/D���TK�#{_6e�&��1��ᑇ-D��J��	�C��c�BP�g$�y;�0D���pH8�n%�Q�ʩ1ꐡ�.D���R50m�,��i��A��(�M:D��#$F$���+�e�2��;D����"ۍ\�n13O[3Zr�(k!��rAZ cX�h6,�p
A�8Z!�-gȰ�PEA&X3N� �izC!��ɞx������Q)!�ƌ�b]!��%D=MC�`]"xD��BH!���TC��-a�j1��+�d9!��D)̔1kħY�A�m��@�.�!��H�q�حZ��� M&q���[�T�!��L��X��aM(Z:�� shˣf�!�d̋�B���lˁ ��	�D)��!���!��e{��0Y�v��vh�(k!�d�`�� 1T��>y�b�i�埳G�!�m��9�I�<��ED�g�!���}
���)BA��#D>#�!�9lL��'ҵe�z�2ԠJjw!����aa�#�(�P`Ғp!�D�Ow�(��]��@S�P�X�!�D]��NabI!tՀ\�F,�4(�!�/!Wf!h �?�03�^(!�D_:���cT �X��a2jP�x!�$֔Ow���4-�nk��+7i�in!�d�YÜ�� �X�]�����:u^!�d�*�N�3�+X/rL8��gH�I!��G�x�b����УlD��&�F0x*!�aS��`��� Bp	e� :�!�d�u��[�D��f$M���-Z!��X�5k6��c��q��ڱRM�{�� ��	2, �|�2UAc�M�ZPV��"O���A��D5j��a��'hBSb"O�qJa� �Ro��[�N�'�f]jG"O�Q�@��;o
��M#�X"O��q`Ўeb䅛�,�l�"O�0ǣ��Q4�j`�m�ʕ5"O�-���C(1�D���i紴�"O�=1�/�$U,q�o�8N���@�"O����!1LP�����6��0v"O��#����J�IB�E���cU"OD��V�[�F�aU�)&�zX(�"O����WX<���Q�k�J��"O�����,X�� r�%�H�"O4uQ����ļ����$Wv�A"O�,����
8���E%3J Z3"O����H�uLM���۷���"O ��J�6��ȕ��v���"O�8���\�GH"�X ��:>x�x��"O�t�����ٜ�vC0"�$&"O�
��ST_��C�+p� �b7"Oj�Pt"ưIQ��:������(A"Or����ғ*��A���0��T� "O��1(�G�=A����6�.��"OxE�%�|��aIońy�J�"O��(�BԖl�@�-X�C
jL�"OX��Q�Ӟj�=��E'z	�XR"O$ �A��#)��ـ�OZ�$`�0W"O4&�2b��(&hV�]DE9�"OH㩙}^� �f�;y;^}��"O�`C҅{�&5�d�3F��"ON�ɰ$U�C�^Tʃ���Y8Nx�w"O���ɺ:w�8���|���S"Oh����ip@�"�|L��"O�!24�D�/T� DiDL<�W"Odp*f�W�5dф3` yr�"O�(sCؖk��y�'M\�,U���"O�����@R (
�ɋ?֨0 "O�d���~k����׬%L	(C"O��� ��=�D2��ldQٶ"O���`Q$~�	;g�B7{�ts"O^!҇�0|-���CO+N4x�"O�h�`M9�9�V y��!1"O�#3��7�,�h#V���V"O�Ie�(B[�Sզ�b��e""Ob,@�E�K��	KˈGd(�"O%�1�!�6��S��b� ��"O@@�7d�'E��U�"DG��Nl�%"O�B�΅5��1���Z�Ҙaa"O�AC���?s�@
TjZ��.��"O@����� E01VÑ��34"O�"dk�Y(zPS#���]w���"O�Q	�L�-rX1�W!� 5ml��"O�4(���y��2�OC5w���"O���A��t+ژ`����|p�`A�"O�aU KCN�A���QR���"O�r�B8I(�d��k� 
לJS"O�������xб͍���M F"O�M2�� mih581,�H�8s�"O҅��m����
��7��
g"O�M(���GE:,#��X�2_t��"O�lԇC/����h���"O�pj���
IIW�� ��5R"O6�1 �R�u�v��v'W�)��B"Ob�3� �!xc����l��?6�Xy�"O� �}u�@�4-�Ct���&6���"OjXd	�,cB܁eA�+Br�Q�"O<�82-I��)H3� 9r�<Mi"O� A�ET'�P����U��q!"Oz���įVk�}B.�:Ej����"O�u��f���er�U�S�p�f"O(ai'���q�(���N����"OX�����#PMlA+"뒲d�pD�"O��A�,����A��مY�JQ �"O:����g:Ъ)�6�^$P�"Oz��U'A�{P$+2I��	~��J�"OJ�"Q��&l�T���,iT���"O8�+���C�z��v!A3A�Hy5"O�X���>�na:2���}�>萇"O�I9�۾{��Cďݸr�u�"O�x
��βV��O�:k�RV"O����Ч(�����:V�$��"O"9j�/T�'��H�l,����1"O�8�Q
��cC���R!S 9�&Ŋ�"Od�J'd E�Ys�5����"O���3�߬	 6�zG��#�xr�"O�DcS(�
py�LA�I�q89@"O�:q�I/&Ќr@iZ;?hlkF"Or�R㛛;����5�^� 5���"O�L� �d�Q8��bQV��"O�S��0�1���Xe�0�Ap"O���a#~J���P�\�K� ���"O����eh~i@#�P$��d��"O�!���/ZY D G,��!�6�"O��pf ��@g��"쀀=�T�
�"Oڴ���R(T�^��UJ
?�\���"OP 2%�
>����G	�<	�>L�f"O� �b�+!�(D重�H�t%�S"O�!󒋝@"�%��N��z��r�"O֠��٧*|�Ca��=-fF0Q�"O�,�q&/a��m�� J�ikv�*�"OR��NT�"��0���	?rb"O� RX�$��u�g�ߌp%�L)V"O�$b����M
�N��W=�!$"O���kL6��� �ٵ6�NE�"O�x���Җ�e
�"��dsd"O�Yw�
j2T����,ƀi�"O�����>皰I�g_�H< �"O��ZLUd��;祘�9p�"O�Ԙ�d�O �9��-a2�X��"O,��K�}�d8�듋AR�{�"O�J�T�(��Fh�h�q"O2���i��h�h޷D���@P"OP;$�DV��� �xD�5� "OT���
Ӛ�\l� @�l8�"O��%�= ����%GXގ��b"O��S�Ț�~в�!�Ɉ�z�	�"OH-���T1��X�Lʰa':��E"O|� �KעHxAA�B�� ]��"O]���Tq���V� �����"Ob���Q �\QYs�C�+t\��"O�RӀ̆Pgnu��l�aV��9T"O�����"x�}
@,�K�>�r#"O�p��b� ��|"lI+�v��4"OX�R���!���v����p�s�"O� �F
.5(SPMFc�T�"O�]���ȏ>���EM_ ��)r�"O:�fgHv5bY���ъR��a��"OBAH��I��U�Ũ�	�.]c�"O� T�3�^��ȴ�fHY�
c��`"O���tN�+2�e��@�t�m�"O�x�a��'q�N�:��I�x`���"Oի�hB#|a�s��tBZ)X�"O$�� OX?(�����"s<���"Ov�g�P�\+��[
7�!��"O���/~r\�T![�d9��jT"O W������$q'�]k�"O����:^o|��GKD� V��"OT��#��6�X� �I��0Q��"O:9��e+�-�#kS�$���G"Ǫˆ�9lU��I�3F����"OJ�Iva�-j��U�ўw�hqQR"O�s���;�P;�gۛD6��X2"O�Y�Ι�H���s1��o7���W"Ox�I��C2^Hzŏ >!��"OnU(F��z`��� ����d"O�ڲ� B��܁��K�-��l:1"Oh\+Gb�"l0)����5w��s"O�m��f��%�
Qⷥ��
9���"O�=��IK%R��0�eU�ƕc"OleRQL�
���QAy:IaT"O^1��拦�p�j�J�w�l��w"OPq���.t���Q�5�V�8Q"O�@�#�/Fkx��"�@+`�p�R"OEY劖8c ��B�^	\����E"O���q�]�T{P��D�GGH"OlI���� �=0a��%�<8{""O~X��
lq�$j��ܳZ����"Op���.��pVH�Q(4��"O�%�E5u1�i�W�u@Ν�v"Of�����)��P,7bQ�S"O&��6�*"�T8��$O/x�T"O\t �D�&J�!���R��%�"OBQ��8��I��gRı�"O�)CRi�+2&�s2A�!Qqv��"O���3��F`�h�e���K,]�!�I
ME�`��kG�x{'ǁ�:�!��N�Bd����9�@(1�]�"�!�$j)X��n"|=Z�
J!u�����']�`e됣n`zt�����joF(��'�|	��@��XBT���+Ǌ�*1s�'38���N�t8L�an� ��A[�'�|QR�)C��\��A/+r���'Y������:b��R��{��}:�'u�,��mX�e�H|��.��x8l���'%�ei���}���QT�o�d��'yZ�`���%�n�9�D 3;���ʓ^GȤ��,��G�,�2�� !�b=��	�q(Sc
d{ �醌΁Q���ȓ`thJ�LW;q�������`ْȇ�j@$�@�Ыax���f_ v����3�̻3mٚlN,���z�B!�ȓg�|}�@I��t����:勎�]�!�$Y<DJt�m��SW�P� �!�F0-h�t�K�b�6Uz5(�3I�!��KJx.�7/ԶM�U2"ʋ{�!�޾
�ΔR�!�,~� h�AG�>$!����y�8���j��h���Ҷ7!�$['ZEvu�S�0c�-�U�\M!�86ɾ� ��\�w���Ӧ�/I!�Dö]>�x�pM6_d�=��oQ�<!��.\7R��&ˡ
c:D snR,)�!�d#,��K�:\�݂gC�;%!�� L��KG�>�Ȝ;�'ŵ1 �-�"O>��JݨD/rC��k�Q�"Of�C�)��{�J�As(L=&�`�(�"Odx���Z��g�8803"O����R�l�l��!� By� �""O,��2�P=:Ql�I���vv���U"O�kViF 鎽�'���zfz��g"O$!ѡ�9g����� Pq$�R�"OL��T�}*�i�n 6W��0"Ob��D�_(9��x0l�:(M��+"Ox�PFF!<q��	�(�P;J��	�'���F��O��UZSbK&O4h�'�0���(� 122��6ղ���'t*� �KI�2y�G.�s�	2�'�|����^�Y��鐼l��	�'m踠@&���	��d3�C�',53�[/0B�����%b :� �'�n�� �ܔ��A�X�^6�ĉ�'���q`˲Y��U�!$ǩR3\<�
�'�� *R�˴r���Se� "($�	�'L4]�AR�G�Hs�����ڼ	�']fxr�Ϟ+�4)�Ҁ�+l�%��'����H� .z��c2�8XF�+�'�2`�`��c0y�0`g�@���'����ւH�|���nZ��B�����ΫK�a�a��)j�b������y�^I�V���Ώ�X�fy�Gب�y�A#)�e���Z�tt�i�B>�yR�جT����t��>����y�ا4<8��4oV���xz�a.�y�nH�8[�=٦�E)𵺰�B�y��V`���;U��E�=�@.� �y"� �o�4]�"'S�Fp�����y2���^}�����:%a����yr&*�`�� {n|��␟�y�I�W�>ݒ�-r����dۘOX!��SR�u��&���0�#ńQ�!��D*N��QDB�0X�P��N��!�d#d�T�����u��q��Tm�!�dC�[<��0 KX=o\th�9�!��H^�x&��*Z���!�&�!�D�-(	f۲(G�Il8�c˚��!���l�@�`��P'qYt�T�\=$�!�B=�R�q7���7Yb%��F	�r�!�S!�r0hl��Q�P���"��Q�[�����	�;�������y��(�(e��KC#0x�1�<�y����E�*���j�Te1)�H�/�y�(g���k��'[ n�Y�,��y�D����Q�Y� #��#%i�#�yR� 8�xy���sE��G0�y���d��c�M�o�B���%G:�y�"Z^M��3��ձ;���C�-��y�F�=��,q�Z:�lA���
�yb��7B��Љ¶8`�4�� N��yB".iP���l��[�Ti9+��y���5 ��<b��]F�(��3�yr�Ч.�f��WcXDJ8XK���yB�)4�(!�Q�*ht�u��:�y��UO���P�&�Y$,��O���$��.qB���W9�p�4�6t�!� �=9��[�8U�H{BoU�y�!�\|$�%3'fZ�FD��d�p!���x���� >v=p��.6Q�I韌�?E�� �y8��=;�vqR�HY)ใ�"O&���"m:L�7�Z q	h�ɶ"O��PU� &2M�q[e�A�!�~��QO�O4��O ��$�/.�L�#�Bn�,[FƂ�!��I�Î��R�@	-V$tj�-��!򄌞7����M�xIrPk��F5�!�D��n�]c��Ǽ*_�hxU-J�y�!�/|.�|(�	�D�l���N#�!��L0|�h�afLs⎉R�NO']�!�ӷL�b��F̄a�� ����m�!���y�X���B���P3 �!��C;�pX���t1R�Y'���!�d�blܑ�7D_9`"�'�	=W�!�\l �=�/G(D���+7T!�D�l�m��Ն%$PS4+HBE!��Q�R��d��*`]!A�<cD!���]w��p��G�/��ׂ.#C!��V>d�z��B'��x�@��< #!�� �D8#��܄Wź�D�ՕU�!��L8
B(�*I�5O����0@�!򄜪�Ze3@jH����1��-V�!�گG��)�#�LcP����Ȥ!�!��&8oԝ��h��ra�af��a!�$G��"���+D@��f.��!��1�T�
�G,+��03�,�)�!�dJ���=��;7�fX��ݯI�!�d�;E�:�-F�ou�c*�0�!�h8�	$�%!Y��E��G�!�ˊrL����Y�I��ٖg��!����
�����#o��� )R�:�!��UF���F/,�������+*!򄃪 T9�͂mϸ0Y%͑�!�dR:Nl¹�Ռ02���U�",�!��ɖad��+�ާ�N����8q�!���EM��)e��d��t*�ǚ�8�r��(�O(4�c-�0Y>�8�2�AP"Orͻ'��|���J��.�ܩ���5��hO6�6lԱ%�4����̸N[rr�"O�ܐ&♲|��5�� �3OB�H�"O��Ï�x RQoۤY:�U�"O���ʙ$C�ME:6���0O���8&�||�g�םW�8 ���D���D�h�w`�+�!qF�Ҫ�H%��'��x�m�\8��A��O2��
�'�(�K�K�]���O�q�T���'ersIґi������ԫb{��
�'�ɑ�˜�b�xON
\hڙ��'�ڄ�'�ԩe��tp�(T,X�F̩	�'9ra�0Dˁ�.(� ��V�P�9
�'ɂ�wcW$.���R.�
VA2@s	�'D@�3@T�b�t�٧�X^�����i>UD{�O����-�
J��q�䍒��yrmѣK^�@��'=̆���k��y��ƽ-�=�sa�4���[��
-�y�k@�؂�HU�*-�I�r���yҮ�!�
��7I���"����y���m.����P	>̜�e��y2�
�njx�'D�/y�|`����y��K�L8䁤
ϣ7��E�%k��y��'3X����>h>Va[0&�S�PP�
�'��yu�ߝBa���Oٍ�<��	�'Ҳ�"���F����O.�hP�y2�'��O1�6� �b�y���ҫ]^�j9�7"Oh�14��<&���2� �?�^i�2"O� �ͱ2%KS�Q�ѯQT���"OJ����N]*��̓�S�@���\��I�J�$��"��D��rk��-��C�6夑�e�L�pD�Qɛ	~��C�I�	�d�*�a��ij�KVÛP�c����ş�E��EC����3�x�͕�yrF
�*˺�� @�0
����!�
��y�/�k|�����7~�*`�o:�y�dp�P���)y�⩲è֓��']�{���WDNٕoT9n�p����y2�έ[�i�Y1"\�����yBC�t�.8�	��Fg@qba�W��0=����� !zr9�A%�:��9j�Ą����O�x��U$N V��:�O֏Q]6y�-�s�<1PF�?�Jlbqh�0go�<I��4�h�t�c�97|xZ���rs�YQ';D�d�æN�F�$�+�Ɏ3����9D�ěA�T<i+�5K��J�/<�a�6D�h�a�]I2��:hIA2�a��A�'�ў�݊@�L�+T��JWNa�.�9!g����Y�Zy���M�!W�9X�+U�>:�]y��Լs�!�$K�L9(���Iߥ/0�q�¬��$D{ʟ y�)'3����H�ZJ�3�"O�y��gA2m�]���N:���"O���w&9���j����f�"OH�����c4�� � L�]� ����	�F� �	Z�@�(�<��d�ybÜ�>p �E�e�1�ׅ�*�yRo݉/c�!TL.i��d����yB._�W �����P"x���K�	���y�`'W*�`l;��ig�7�yR��6(�(|�য়�2���U`F)�y�oڙT_l�A�G�$��	�eF�<�yaD.
>z]�mR./��8�t 6�y�n[�Ra�UD:-�b�H��N��y�8l��mY�.+C�u$/�����O��=�|��)O/�(R#�U�8�y�v�<1"�!=��,� :�P�0�-�q�<��
�xV�a�K��ǜ�6�U�<1r�D���9t��3���Qc�L|��$�l �
3�!�R-�P��]�� �Eh<Is�*w�5g�q�S�Qk�<y�&�+~�8�����?�N���� �<9�����������/�@ �%^�R%D%�C�[�9v!�dH"_���"��&���@!��Q<+��iK�7Ṯ����!�D<��!Ut�H��G�.�!���q[��Yf��7��5A�%�5j�!��	��sb�2	���r�v�!� ���1ʁx��0b��
���d&�OH�hGeX/|\�9�v��26�k#"O8e�CW�9������F����"Ol�+��?'��<S�&��-l�, R"O�k�`۠f�$)��JkJ�Kr�'��O~1�D�qʸQp��;k����L��	�jv"U��L24�80G���8C䉿��zĊM2eR�h �Ɲ�� ���paS�%��l 1Ѣ�B�.`��>��B�-[*��,8N�pń��*��*ȶm��H�A�l�N�ȓ}�N�I��NԈ�C��9ފ`�ȓ���Ѭ�8v�>��b��7z���ȓON����G�p{�I��M��	�̈́ȓ�&�!��-"�tu#áG�i��@B
��� �m��ЫA���Ul�%��S�"Ot�o�s�x�#��R3D	�bT"O.�ɔ$�6Qk8�1IK�D�p*�"O��K��vR�I�S�!V񬌙�"O�-Zal�$h�F-;V��T2�a�"O��[�ʁ�W*��{��M�>Ř`"OB���3JH��Bꅾv@���	O�O�0��T�y�Fik�E7j�b	�'S��U�&Va�=� �}�>�3�'U�QրəV��mJ@�X�| �$
�'���c	�*�
�0�
��n�l�i�'�0����P�4���%_����'B��#'Ty����u�-&�Z4��'o�7Ӗ4�~�@��Y����r	�'A,��@�ʼi≥D�t1i�'NT�Y ���R�j@ ��ˣ8�Q�'e>��"�'-����FY�*��i�'0��W�I8y���F�I�B&����hOv�3�T�эs׾�5#�I;D�,@'D��!'��p%$����fB4D��q��گy��9S,@�,��R�`�]h<є�D�|�H4�`��:?
����`�<i�d<MNV�ن�Y���U��P�<9�씗=+4@�R�jX�Bd
[X�<9��/����w�ϴ}<>=��UQ��D{ң�$[�|�J �ul^��n��yB�5���!n��b#v�զ�$�y��S�1B���XҼ�; ���y�c��Z�����ȍ6Z̠���a���yBC،�8�kRG;m�=�g�ܛ�y�HV�s70(14"@>5��5��F+�yB$�>7"m[�ꅚ,:����@��0<����'�Ӷ�Ģ�Z���.����"O�dH�c�5G�-P�dŵk�<G���J}��a��	M؜���	�i�<a�f�(s��%��/W\� �Ji�<y�a�a2*�H�>���'u�p�ȓx,p���׵a��ɶeA�V��ȓ�A�1D
5Ap����D�4�$�ȓXZ.�#�y�L��pLņl��!���s����Ι�f����'g�� Gm;D��Z��8+����ϛ�9�ȉ:D�l`�ޓV��A���#]�tQq�=D��y�$B�e�T��Q���A�@�a<D�D)ALV:�ؙ�G�PP�l��5D���6hT*X\� �Un҇x��wf5D�tK`�B4
<	��θJ�Ji��O&D�آ��Ə=�R�p�f̀oAr��f�0D�P��7\�`�I�`��*�\�H�I$D��JdQ$nZʜCɊ#�XT�@�5D�x�7��y9�5C�~*���4D�`�`aښ;E>�g�T<<�l��0D�I�߅k����F�^S�i($f-��hO�SCV��à��*���GC䉓y���K2��8�.s�*x@�C�Ɏd��R1 ��p�&����=�&B�	"�� ���c�N���S�`�ZB�	;rH���P�1Z� o�
_4B�I�l�P�3��}��
Q��9&�B�I�T~���C�uE���- X�HC��.- �F�Y�kҬ%��_&DdC�I�:5�#��]1��qv�+07�B�="s��`� �MҤ��cJ�z��B��,f;���N�;V��K,C�)� ���+Lu;<!fI��+[���"O�p Q��4y�L5[�瓙08v�st"O�%�2$4SAx @D� F1�D�"O�L�Q�Y6^��(#PF�6�88�"O�:$J��z��lh�"� �"a��"Od}0D�H� }Ȓ��4�Խ�s"O��C"t�L��K�8�fE[�"O��\E��� �(�ov�K�"O(Q+wEҰPb��,E7	an���"Ol�"���x<���jW %H����"O���%�)|L�0���o+�T�W"Oj\��@H�fD0!�h�9F ��0"O����#S�<�L���FEq��Q"O���@J\���fL7	b��"O����c��yC|��k
40]��`�"O��92
M&Z� ���@����"O�$��D��YTe�6EБ<��LC�"O2ق�fф\y}�NA�:�F$�G"OJ�s��I;�(�6L��6�-�&"O,�K`"�:\j2�r�*[����u"O0Dy�g�'S-L���䀈w�ՋG"OB<����
i�-��G0D~0�d"O�$�b��7�B�`�"�l(j�"O�4bc�� �:͠VB���)�G"O��Sp(5;�f���g�
�<͸�"OBYJ0mc1(9�P�ݐI����"O��nP�0h�y��at���"OZ%ap	Ӻ�q�g��;
�"""O�؈��Y�hD��Ea��d ���R"O����B&Fg�S ��$J8��Q"O��s��gf<R�@�4FPQs�"O��*V% ;ap��fOL�p`D"O~-�f��98�N�I�Q�"Od�ҷLT/g�i�U�'Y�)�q"O�l9�E�&Jh�hQ7����E�"Ox!h�۬M���b#!o���S�"O�Ț�f�H��"p�B�{��S�"O�����C�t9��e"5��ZC"O�p��۲*+z ������#�"O�%��BH��0�hX2 �!��"O�,Ӽ@�Ҕ��Ʀ}X�U�4"OR�t��BdP�C�eE@����"Ot\��G��0{´��g�/�j�B�"O�I�.=(�4)&��?� s�"OF��4&�*D-�D'E���t"O���p?�w�K3�X-*U"O\1���ˏ
Z�=����m�^��b"OB5��L�"<]�BVK#C�LD#"O6)k� O�t��\B���O DR"Ohٕ���+��x��2?���Y�"O�x�G;uVX�c�h^�H�$lP�"Or��eѮMi�j�BWc�ё$"O��Y5aQ�f��R�W(wG��i�"Oΐ�`(��/��q��&o�VY��"Oʌ�F�q����@DQ$\�F���"O�D`F���U���\�Y����"O\�*�͌�V��i��)t��lR�"OapW- >��9�da_�x�bm�`"O�E"�O�H�p�%����1�"O�������CK�gn����"OD�
PZ<#��s�Z7#k��p�"O���� �!r{���1ǖ\SN%�r"O�d` �&O���QK
Q<-� "O���ǅC�f@ȹ���u%��"O� *��E�N�\7@$�p�C�*
Uʱ"OJhB@
�f>�&�����"O�Չ��L�N��h��ǈ�w5&���"ON����֤J�ܩ����e*P��g"OZh��ߪN�@ڲb��!�M�F"O4���ɝ�v�7[�:8�|x5"O"�Y9G����0��q����"O��3�"Nx�!��!7�8P��"O0᣶��UD|��T�_��0 "O��Fɀ�G�����	?ʵY"O>� �l���${5e�!W,@P$"O^,j�!/w���ƃ��&�0�"OP�[�+/H����}�8)�"O��1��[�-$6��7!]}�	�V"O2i���vO��#�e�b�)�"O�Y�k��Q��a�WĈ��|��"O�Y����N�}"��ϓ%w�hh"OB��'ˈCHŋ�%�BYp��`"O�=Â �G۞0hUbݠ[ڰd+F"Od���`�
�AI��Vhp<P�"O^����Zt�8t�RhMec"O�47Qx��V�	<0��"ORYp�ǘw��l��ڦQf0��6"O�Ha�H`�b����Im�8e�F"O�	TȒ�4?V����(�!"O���ĉ��z����f� ~��U�"O$��w ��T }�K�v�\L�C"O�8�v�C�'��Ё��ՌyJ�4J�"OE�N�f�L���)��*5V��$"O^@�.ޯG&x�ڳ�B�R��"OB,(��^%.R��#�Ћ@t�ب"Ov�3`ͣV�t1	7;�Z���F�O�<��v@�9Ub(	�փS�BE�q)
�'m�,� �@�dl80��ˁ+̴@
�'Z:Q�v!-
����A�'��Q�	�'��}b��R��

�% �ġ	�']�)����?v���ζȒ�'���q��<#Z�P3s��	u��X�'��zrbG`#�d��i��Uz
�'�*�z�*�a�p�e��\Y
�'5R@3�Ȯ6�mJ�M�eS
�'Δm�яE�#.q�Ě�0$�y
�'��Py�.� wn�/��H�g��,:!�DΔ@u<��GmW)w���� [��1O���OУ}Z��4Y
�1t�ۜU�>I�f:j?\��.O��D/5��5�w�N8����MT�m�!�$�+d'������S+�\9F�՘Q��D/�S�O^�h�I�rSPp��j�0S��	�'Zu�7��'^0��H ]4X,R�'-�����PF]�4��D�-;�'�H�ŵq�Z���ڡ3j��
���'�I��uӖ�06
@�)RiBB̅��yB�'
�C@��*�ȂU�P�"¼��'GPx�qppP#����!�	�'_t	��]�4���p��gv���'?�Ͱ���.a�~��qBO�o��j�'�6�#���	C�ЃvO������'�$�Rh�9�
yq�eL��z�'|"��3D�"�Y� )Ԋ�ޝ8
�'�y�.�TΎ�gǻ|��x{
�'&��������B��H�y�"�8
�'aΰSeN���~�iVC��?E�e �'�`�.*t�쌓�k�?8�X�'�|yG�Lt�$[t��7r��
��� ��X�HGC@�e��&S@��"O�!g�H[�H���<;��)�"O���h����!�L����3"O�0�E˛��8�$Eʗp4K�"O�񢉇�#rKҢ��q�~TÔ"O�-��Ru?��`� �64�s"O�ݘ�ǎ(��k5�^!�\(6"O�`��#�]����q�\�J�	��	]y����O���dí4��,�g<���xP=Of�ON��1��N���"��''�ya�G�$#M�ȓ-��C�e
E`.M��gШ+8-�<���<�1�P�����/�	ER�
S@Y�<a�Ht}a6f�����B�RS�<aS��U��QRD�-�03�P�<��E:.Gt�c�
�s� a3֥�d�<�e�!�D*�	� C<1� ��`�'^�?�h��F�H���9FFu�$Y� /D�L�%�1BZ!{ₐ[V�|�l���,�I}y�'��)�s�����%Q��8��͕��Ȁ�'&D��Q�1G�< ��b	�.�L�D�%D� h�P	&�����>H����#D�L1Сѳ,�l{Rg��@���E�?��hOp������X�!�"�&�s��@6�(C�	 )4v�!u���6MX��.[[�`C�.|�Z��e���=���	01����hO?Y���\E�e���<Lrj]��	3D���bm+cj8I2�v�I�"�1D�$�Bk��T�C���Y�'=D��Il��,UHX�DB�s]�q�#d:��j���Okl� �圩T��bs��/f������'�r\�D�)Fx�ߣXed���( �0Cj�	�jM��y2h�!d����F�'���UK���R�'�rT��'��O�M�C�@0�����_��̸���`���;@���O,�N1C��&B�	�m��,1�)Һ2W������N`C�	3>�ƥ�4�3��qz��ͣy4C�	!
|�x�m�@�2X��%�se*�I^���$�$70��K�`�9��=��D�+�1O(�=�|��ª��Y"�d�q��x�&%�[�<��&H
.��2F,���"uM�|�<�h�M�6T�����|� A���v�<Y!���F�8��ri�6#;p�IWb�X�<�á,�%IEN�7}��s�[�<�'/ǿK�z��'ʏ#v�)���<�)OܓO?-I�_
E����r��'f���D�>��y���O�(����e�T���U�4���87�'��'ur�'��ey_�d@Q<�4�B��U&8��Y�#;D����S�~�>b��+5{дRt�7D��ْ�P�V	�=C��ڗ}����:D���f�^�T�~���b,a&t�W7D��I�V�V��E�`�,�=��Mt����5��cwχ�pڲ 1T��9[*c��D{��DI�= @fM��nQ<��e`��y�ƫI�K� i�8�#��+s`<a�ȓsRb@����@��d�D
��:B�)��6��|aPOI''n>��eE�`�"|�ȓ] ��V;#t"1��-;tj$�<�����P"u�����T	\0��k6J�6VJ��bx��&L9X#"!Kf*��o�㖎'LO��<K��M�Q�m*i `B��Y	��D�O��d�O1����<qP�H�|�`ёXr�@����%��C�����Ѐ<F����G+2�{
�'O�5��I���r���<t��UB�'�<�ġ����U9ƌ�9ޚ<#��d;�g�? v�c�׹X���Q���(3��!i�i!4��0"�h?�Uy�-�]Z�qŤ%D�(�g�D'A��9�20a�Q(%��� �?�O��ٽG��4#�H]�	�`QĮ ��yb	0v9b�8�H�~��A�$���y��hb��"A�5GJ���E(�yb&P%+��y���;�h��LE$�y�$ٰ� ����+�HI�vD��y�-S�@�XE���()&��y2ˆ1N�B�X�Kˤud T;��3:��Z�������?).Oa�F�L/W6n�#Џ@�#������:4���3cB�PlӢdޘcN4�Ei+D�Tr����"���矆Q��*��3D�H�W��TzW@�,m��".��)��`�	�����o�I؟�ٰ-)o6n�Ѕ��/8��i���f�@F{��i��YVp��l�u&ȕ�PI�U!�Xm+T#�5
N$�qQ),��4�	Z���?!��~C��a��Ot���*n[4I�ȓj�� ����$�(ЯY�]�ڼ�ȓEV.1��+�`�
��	�#`C�4��~
��j��SS��U����7or�5D|�S�7}B�sa^�Ef.	г�x'�C�n� {%�Ǜ/�
�F݋��C�I"`�i8���2Ӷ�"	\�>�vB�	�Lp�`� �W���T	稝�q�|B�.!���c��ֿ3�v ����(0�C�	K�f�B.�a|��*P�"+*C�ɝ+5걳�N
>��@Ս��?�#<���蟤LR�I�Wj��rң�	]N�[D"O9�u�74���B@���4�Q"O���b�<	�!�2�վA�`IH�"O�M8�[8 %��C� P�r���"OftٖF�&T����ĕ|���u"OhtJP(�b�� �!n��,v�)	�'�*����%}q�pH��2x�5a�'e�U[�7sO�pK�a;3�� �'(h�e*��x7���U$9(�lk�'�������
L0�=�pJ�2$�x�{�'�8���#�?'!@�D���\��'�r�#G��u5>T��$����;�'���� �Z�2MAq'�#X��'Ŵ�0�V���l�䯉%S���)��|�\��]��<Q6�M#i	��rP�Y�o�V@�ѣ�y~��']��pv! )L�����1
�����'��`f�#�YaT�̖v)�P��)z�m�,���9�g�gZf�!�k�)�y����4�a�Ԑf�H�����y���`�TK�*Ln���,�yҪ Y:n@�Vo���B�yr y��iTϪ+�p0eG��y�C)vN��4���}�����y2eԪ����O�	��K��y��ּ� �oB+{Q`�A����y��&1B�+s��A�*���@ʩ�y�@��� �'PĜ,�AҌ�y2d�o:�`#�*��M�\�Q�/�yRD��c(�ȳKSKl�	� ���y�jW�MOm#�!ԊAh��0�gJ:�yr�J�\ȑ `�(@*����-�yG&b|JH��F���^Ic��y�ݣ�Nx�۪v6p-ٶ��=�yR�L�D	�`AK����]kZ<��'���`-� '�`A$��T��	�'% ����9P��F�ɳ ����� "�#�خ �� d���*je�"O����.���8�8`ˑp�<�D"O,e�.J�c`��@ί0_"��b"O*�[��މZ��d%ƸPkD�A�"O�A@G�ӏA���v�Ս��H�"Oҡ�h\�@�r��t���A�[�"OhM����T�~\��K�	�ʹ�e"O��ò�N�ze+wLJ�K?��x0"O`]���[?	T�1b�0 -�Ԣ�"O8-8D��/:���R@�]�y�7"O�l�%��&f�u����" �[U"O��hj@N?�d��:,�p��a"O�;�c[K��[2$O�n����3"Oa�FJ�=��Ҵ�&��h�"Of���.P���3�݄Rk|͹7"O��;a��F͊�ʓ"�T��ia3"O�
��Q�${�AK0�]rw���"O�H v/Q��f}z�D�%[��33"O�YلiU9.�=!aCM1yP�d1�"OL�C�e� ��R��X%$*�t�'��ɭ.�����+�g������!t/�C�	�P����aY/(UӯԘʬC�9qN���&ːc�6��M��r�.B�~��8���R�!:R��Ҋ�"B�I�u�<��)˿#6VHP�h�}� B䉯4*Q�c�I�$����ϻzh�B�I%����� �!����5��I��B�ɬfN�}���;6�BDL��"�hB�	0i��p����<d�b7�ׂi�C�	�/��qK) 8q�����G%DB�	4*>��G�@R 4٢��P�BB�I;8E -��k�b��Ƞ�/��C�>�j8��H2_k΀�I�c	�B�	S׎�����0rT��P"˞b���dD�as��S�Xjɞ��G&��D�!�dF�|�FL�c��&� �#��	Y!�D�W�n-���\��!B�e�b�!�d݇q'���vj��`�1$E2w�!�dW�gm��a��X�T$#�#ј�!�DH�}�L�b�@��e�
�a�ߙx5!��@1H�z�:c�t�d���)�!,!��P|"V���LM���1X!��^�v� �-،>5�Y���7s�!�D��c��]XFٖPX0�c��7�!�O*_�*qi���E��0g,�w�!�D_K�:)�r�� p�٨�a�?(�!�ǆ\�E�&/��]��|ZtO�!���0_�^�Q�1֨9�o�%�!����ހ���#Ղ|��B�/B!���.;���@�s��%�gB҇6.!�N?]Xv��$�:vC��p�Ô.)���d3�MN�%�Oǯ�yR�X�,h���"o͕y�Ȃ�Ϟ�yr.��&"t{fLT�q7���$��yB:1l
&��*8���*C�y�m·c	�`K��	1b��S�yҎ�5\?hA��E�q�,
�K��y�H�fO��Yc�(z`Č���ߛ�Py�n_�#T�@��K�s̚�Y�@d�<�!���l���6�3{���CD��w�<a2J[h��ո�C�M�ސ��nI�<A��פ2�.̂`نMw���AMB�<��fU�6T��NV�D�µ��F�s�<���+P��2�ML	,�{5H�<� ��"�hF�>A��2���y�4Ma"O|��Ň�=��)B��^|<ѻ""O��q�"�#Z�6bt�SDs�I��"O����^�
63p�]4ELX!a"OD���l�p�6�B�D�J;�iu"O�e�kX�4�"幁�[6+�ܡt"Ox��� ^T21���;�"O�A�DT�s�ļӒ��q��R�"OFp����6p�$�TB�\�h���"O��@D��~�x+�&IP��X��"OԹ
�J��3P2�Y��?a��D�"O���i�o̶�* ɺZ�D�R�"O4Q�����$Q�H��AE����"ODYP�&V�
K ����9-y��"O�������>d�Xz�!Ty �"d"O���c��-3t2�0��(9r�"O�$�U��<Z
��#���$�T���"OD9(6,ʹl�HL"͙Bf��Q"O(���$R��6,P�d B
�`p"OdLjV�5~Ԭ�R�60x�"Oti��&O(zh	�F	�zΪ��"Ot ��8�`��f7L�b�k�"O8Xyq$4GQ�ϑ#?쥠V"Op�0�#/�`%�q,E��C"O ���%�?3���3���!+��<��"O4I%����#�(^/h@��)"Ol�G�&3y�J�'��|\(��R"O�e�Ꚃ"��}�Dĉ�WH.�R�"O�15EӼI�(x�r�E�%<�%�c"O`!�%V
lF�q�*����"O��XT�W��N�I����"Or�2�W0J[j��J��<�X&"O�����+2��UjMS Rh��"O�LJ� �S���	ή(,"Od�F�)_4���r��wt����"OF�i�ìE�2�{P�"#�8�"O��cN�0Yㆬ͞��9f"O
i�*^h�c,�4G�,�ic"O���ͺ|�& � JE*7	��r"O�|� �!��E9��Ç_ �2�"O�5q��ӠMV��!�H�$��]��"Ox4� �S6GZP� �+P�`)��"O�9�Q+�k�j���ɜ ��@�"OJ$��L�] ��3��?]��U*a"O�٨�$�8	cTy'#��ZĨF"O��*P�F*
&i���6�z%�"O���c U�)�̙дoZ.r�z�c"O�-c$N�bt�4.T�yo�ЋG"O}��iW�՞�	����>:Lpp"O���o�-| I��OXƪ Y�"O~�;�NY�[��i7�R&��st"Ot�@EDF1�@�PVJ���A؁"O���7��Ĳ#��O$t�t"O\Uj��'n�8E��f01��"Ol�q�fX�%1$Ar�	(�"O��He��VI�ٸ��1`�"U2�"O�,��"J�w��9�6��>���"Oh�s�������f�x�VXb�"O��`��2(�x`�"I�J�����"O����&=��dA��9Bf�,s�"O�e��O��1�� �W �=~1 ɩ!"O>pC��=���x��˳*)��"O|��D2�̨��P	B ��"O�i�rm_�ULi��$"L����>D�� H �VHRÂX3A[]� 9c"OZM�!�j^�`�C@52<�8�b"O��SC��?U�|����5(�|�D"Od���'_�gH�H4.R0���"O���Tm��'z~��@�^�xp�x"O"A0��օI3����ˈ� д u"O�Xc�.�L�~p�3jݺm���"O.�IA���~��PɃ�U����"O4�`O۟C��婧���y�h��F"O(�;D�=P< �IdN� f=��re"O a�W�a���
P-,	!�=b�"O�!@ӋQ�.-��0c�ƂZ�Z"O&�6�K�5dt�"���G���K�"O~)��ˎ|����j�]m���R"OR�����}�6���>��8)�"O*h�f�V42X�G���̒�y�o;/�ҜX���m��h��yr���/���KR�v����N6�yB%�6�VE�G�R��,���"�y�Z#l�^���@M+N��b�%0�y�*L��>��p�^5\��D⴨���y�	�A]�`��*#˼tR��O,�yM�\["�1"�	���3��6�y�jP�.��q��ԭ��e2�F�+�yRDF88Rɺ��
(�N$�E-�yo�H�,A���[�
��1�0�yL���t� �r~VcA�٬�y�nVrx��eЂk�nsQ���y����]L�|yE͓V�:!��B׬�yr�
P �K�\���s�)ͪ�y���H���(g@׸)��䳧l�%�yRc�:^1,��ӈ�(;���C�(�y�@�6;(��2n�T��F-�)�Pyb
�E���Ʀ	)�<pR�bVM�<�Ҥ>IW�)�6o׊�Q�dK�<aaoĬ��ږ\;N��c�ˁa�<a��?�p-�cA�.BH��Ȅ�Lg�<!���%�6r� ��2�q LBe�<��R�(��lI�G`vh��%�b�<yg�ε)��`���&�h�ƌ�U�<7�--�8H�c�B<�b%�R�<9i�-z�&t�uNK�y1��掎S�<)�&Ň\��YW掾y�8y�0B�Q�<	�ᘍV9�]�2eJ�i��)3�U�<��"�1kLP9��:;^�Z�i�u�<��ٖ/�α
���.>�����o�<9�U�SMD�Q��̮%��0�Cl�<� �Jb6ҍ�ō�f5=�o�b�<�I[7�ũ�@܌J�Xj�U�<��Ɔ-˶P3#�X2[ё�&�U�<�Ǒ]�&�����f%��A�SU�<1�Z��h�$��*`ۮh��P�<)�*��,�N�[l�#r)�͋��I�<��eK�$��؉�j���N�gMF�<��hM1>O���k��8�䲇��}�<��A�]��m�_���j�^�<1�/ �~�-��E�hT�����\�<�'�.���
�MG�|��0�eUt�<ND������K�B@�5�9T�X�M�i����f���\��k)D�TQB
 �cz����0?����EN-D�x���9p��=�q�&s�n��u,D��9D�I�h؈h�`��',�N�Ӂ�*D���D�]P��ϑ bPL��6D�� ♒ Fգ+��Ι�N�`�u"O�C���Τ�g*L���2�"O6���B� �4�)�.y�,Xw"O
%���M]��s����gi(!�"OƑ���78�l��O��/\|��7"O�d�,��?��ɑ��\�-|�y�"O"���mߑ|D���H��R�"Ot�1ˉ���IW�S�u5d��"O��[0H7W +R�[F�%��"O�%▥+?�����
ˑKE� ��"O yfgΠ&�ll��)��p��1x�"OL�Ӗ���4�=���"O�-Z�&�'dI/C!�PR"ON�Zpm@5WF�8&g�  pX�Qg"O��qz�!�(9\��҇�̎ !���B`�� P$i>�h�4�R<.!�DO9r��d�2�H-z"vIȧ#!��-@��]�Ɏ�d�t��Ɂ-!�!��Kڮ����Ȫ�p+7.�`�!򤗸2�p�@�h]�z@��E�EO�!��\*B�� Qh��3����'��1��mh���ㆽm��X	�'��ՙ�$�^(P�{<�
�'�(�"!ˇ�o�H�eG O|�	�'ߺ�3v"��S>����ޱ���(�4��$8��s�X�Q�B�+㔩;a�n|�s�"Oܥ��F9]�^1��MU(�.u� �d�<	ÓgZ~ԉ�h��!����g��弌�ē.�H���5;ŨxɁK��L��diD�'!�dD9L@ �,��#�,}���*�!�$ܰ\� �	�IɎ4�$�U�!���0f�f|x�/W�a��m���ΦR�!�$�@�4�cd�lf��a@��!�_�v�ؘȤ��0�4IX2�I�Q���)�O��dۥ��!E�h-C4o�z}a|b�|2��C�v�k�OD+P2.Ld�X(�y�Z5۸�YV�����bα�O�=�O�A����a��IT��78���S�'��r�ĉ3p�`�cb� 0j� X�'+��BfAڎa5�0�U��Iу�'��2�	O�j��� �5~���'i6d[t�^��f��f�B-{)���'��m�蚎pS<5S��T<w�by��'_�8��ȡ/�X�f���n��UH>������*@��?�ܝ��j�7�!�ي�B5s�$�-)��\1���?�Q�t��ie�Ap, 3�X%+ܤ�d��'B�RcM(c�<pKDۼ$
�'��W[+�������m��4��/$D��@��! "�4����Ж�I�-6D�c`��"j��:��J2|���k8}R�)���8'���e�ڋF��Y��t��B��k�T�)�
[�V0H`+]�~B�I��\0h���n�Tİl�'��C� ������N�Eߊ��c#Bl"lC�	/�q�+W�NS�ŠEDJ�SP~B�	:oVn�Ia�bH��3b"RB�I�a��*$*ђ���i�׉'ў�?m��,0�Q�H�5�Zd�Pl6D�X�N�
������ ��Q37D�TT��'2�iY�	ǋi�΁atE5D���0 ��1�Q�/�9W��9s�wh<)F�D-/ChQ*ӦAp:d���iY}�<�w���P�Q
Z�캓B�m�<� �}p�8!]�-񱀅+1J"�h�x��)��'(Sbg�#=�`v�S>l�DC䉃C�X#��Jʼ�!�Ϲ_��C�I�L�5��EɊh��*,��C�I�$�乙%̏F1�y� )�b�C�	Jur8�DNԌ�pu�uiȫz�fB�	�	`��{q�� �R�pB�;
IJB�	36�"a��n2՛��$B,�C�	�'��5�d��L�=�R,E�u�C�I�(K��Z���(j����|C�ɽ_Ar٫�*K1=:�F
ZO��C�I��`EP�p�s@���O\�B�	�.��q��&D3P� �d�0O��B�I$DC�������@���T��B��7� ���K@�Hx8!�J��X�B�I�#�Ry��uA:�T>C�ɫ�H�9�g��K1�j��^<0�
5F{��9O�@�ЏZH�8z�K QD�u�"O�%Q�"Fgt���W�-��m: �'!��^%�U
3[�B�T=S��̙{Ba|��|�LC+R� @2��
��r%���yBNV�{(�� �N�]���iY��O|�=�OyDU�@�B���CTK�x�.��'Z� q�N$u d��Ģ{R4$����:O��� %	?rU��0ѯZ�T�:!�"O��S�h޳V�6A����z���Bq"O���4+D���xj�ě N{v8k�"O�� t�Ąv6|�)�#F_F���"O��8� �cs�j�!�8KXqBu"OX�xӥ��<�(�r"G%f�dPò"O9���/^�"q�1$"Ӿ,�c"O��cE	K�k�(iR�C,����"O�<9�A��n[���de�Q)�%�D"O����*L (�qj�Ö�:�z�"O,eJ�h�;@��1�śM���"Or��ϝ�i羝{s�R�P���"Ot�%�W=UC��+��B�[��4��"Oh���Z�0N�X����Y�(D��"OiU)�9�mX�����QbV"O<�ȣ�_
~,�Y��
���2v"O�pŏD���Uc���K���u"O~\H����¡�F4�$<X"O.�cH�Z�n �1�۱}��98�"O̋q/��9���B
Y�:�b���"O�}(ҩٙ=�@�B�) K���0"O
�ا"C����RC��X�!�"O,���F"� ����k��@3�"O�� C#�~���THɽk�<��g"O֥0�Ǖ\9�0*P&_�&rdP�"O^Hk���3YG��:�D� AޤP�"O^�����cZ&�0�M:�}b�"O�T�rOܲn�^�1�l��0���"O�X�vĔ�
Z���+���"O�i1��̖dtC��y���"�"O�����٢�x�㶊����r�"ONx�U���
U��Xf
��[�~Pw"O��r��t'�e�G�ف3�<ܘ�"O�����o�� �-�]uP8�'"O~99���4=�p0c��N�<u(7"O4�Qe�)$.�a���S7��cf"OI U�����vo�&�<�"O8aQ��U*���n�'&�ab"OpP�$��5'�� Dm��(w"O�0	�@�8����c���Y�"O� ܜs���,}MH�R�H"@�����"OT-IaO�}f��1��9K|�%�t"O(�����:�=ȳ.L O����"O���#� g��S�d�\��sT"O���%@պFt�8�¢A�f��"O���ʈ"Oi�h�ÐI� ��"OLၦ��D
 1y�.N�T�I��"OJ@8�/��i��̋���Q�r�!�d,[h�y��S���T��l��w�!��4�MT�0�X��Ć9L�B�I;-��Y��
KR|t��%B�	W�B�I0++�QV���+�p� u"��_�B�	�v�اG�$G�J���.�3F��B�ɏi�>%���y�D���A��@C�	Y(Ќ���<y�bP��(�=�C�,%��<�@��]2d#�ؗ3Q�C�	�@���#lނ/�N�h��Ӷ,�`B䉷[� �x�A�w�hy�%�ވh\B䉗$��i��e�N%R�푪%q
C�	-�d`�-!@�}[W_��C��+ЀZT$�'2�� ��N�z�\B�ɓ_r<\��<�)"�d�5BKxB�ɡ1��Љ�K"c���D�ڒq��C�� pG��`v��f��4{���!:�B�	�1
��'տ帑��h�d\B�I�)�䰫刕5)/��V�E�)�\B�	#�&��� ڍ>tΠ� ô'�<B�	&�&���_n����3l^�Qh B�;�@9x�]�pa��2���Tt�C��9���3e�6t�hq�Siײw��C�I�+	�`r G�-�����T�k4�C�	����E[&[q8��b� r�vC�	�nr,Dxpm��c縕
��9w(B䉮����\�ƅ�P��0"�C�I:A%H5��"�N�H�.R1!%�C�	�q2�Q�W�]TB�re ��@�^B�ɇ|�2���#��L��E�'HB�I�-�(9�F*٨@z�X?B��?��-jc�\����!�<j��C�ɼ6���X�oO���%HD��9��C�ɂ�Bɠ�A���I���9NPtC�I�
b*UZR.X* @���NDmaTC䉨g���i���$��4�/ �:C�I�td��S��03�t��3I�4*C��3e����]��kbk��H�4C�I�m���3cJ<��X��ݏh�^C�ɪBb4u
�� =�:�
P4\C�	e#T49���:h-|2�'{��C��&/V��D��;��8���f�ZC��B��S�J`?h�@օA .$C�I�b�ѰTNȫi�\�H�� �A�ZB�ɯl5.�b ��.=[�M�+,B�?~��j�F(zu,�XsI�(wQC��+��w�ž�J����[2MVB���h����m���r�bح.�.B�I3[Ċ`��A��9 �P�3�V5u�B䉇g �0@�D�$S�R��%*8>B�	�(�̅�͏���0sǎĜ=�B䉛2�\I�&�w���šDqq(B��4��B#C�#�zዄ/$�B䉨UHtk�C��|T`�I�h>�C�	�@O�]�`�5�4�ʅ��B�	nKP)��AԺ$zF��nDC��8Y	��Z��7bUА����XDDC�)� f٨F�ܞXf!��t"m#"O^��5�$���8�	�g���Q"O�8"捗-8	�X ���&aK��p"O��X�LrtY����"=��2D"OB����\.�=bV�Q�O^�y�"O&T�����,�*�eBf�$��P"Oܑ��@�$��C�Q+7��%[D"O���$�6�N�c��U�$�@ '"O8�ڷ��B`�	�8L�2 $D�Ha񥟇!�FMj�g�+���-7D�|j��ƃ�f48�$�M��i�P�5D��b��B�jn�M�F1	5�0D�4[DEڨTu��AC��4l�T҅l3D�@�v��Q�`t{��F�kn.QD�/D���0
�ZV����D��Z�Y��*D�@Ƀ&�-ߤ�'	C�F�B� 3D����=����%WB��D�2D��
�G�: �k� Es��M��n.D��"�M��1���;��Q�`�+D��$`�^�.��@ْ|��=��(*D�� �,B�wɂ��C@׷r1�5*��"D�p����:� �Ys
��9�|-a��;D��A��\4��@8 �^3
�fa�c�:D���5�Z�v0x[�A��6�6YH��8D�l���4e�"Ge�{�.Q��4D���TΉ_�4(:QED@3�X��2D����B���@95IA�L���s�3D��WEL�8<�إ�0�� ��m6D�P��J�4T���:q��}�t���4D��3%��v2�a���}����b,D�,c��Ů,&�	��U�H�����)D� B�	A=��hhF�?��{�)'D�� V��-�-�R�X��$n#D�|�� �'&P(QK�b&I����&�>D��3҉S�<���&i��q�����=D��3�+E q�x����G?��Y�dC:D�@C��Y�|^,y�`�Y�|����J8D�4(��6B_�L˥��>\c��1D�(�7�/~�0[QW�X�����-D��d�
�?na;���Xת�� l7D��R�
�?B9�P�jDk��8#�6D������	�PY���7y?�}��6D��	` m�2��d�� -@D�&D��q�EC�f�F��<j��j0�#D�Yb%�$v�Vܱ��߅U7yb�?D�P��Mףx�6QɃ`۷H�$y`�<D�� �咯"�dL#�[�1)��p�6D��[�:;��ÖM�K�t��i9D�� O������7�U�[��]�2�!D����
e��[`,խr2���$>D��˳W��p��a�@3|�qV�<D��U�Y���e�P&c*Z E|�4�=E�ܴ���S�����ѤH�&x��'8ў"|
��ЧyI7���kæ`B ^W�<I�� 2�9B��LxH���_i�<�mZ����R"ǋ��2C��d�<q�	]�"�!��r+�\* �d�<y3��&Z�T�T�B�Jt6m(�AK^�<A6O'?��JQb١X����TM�Q�<1w�܈~��{�Ϙ�G���Q��M�<ya�Ei�J|��OїU�x�1cC
_�<�N�3� Pu�Z���	���]�<I�ň�`1��n�q.}��T@�<9��ƤYr������' Y`�<� hPt�^�o֔�*�Cg|D��"O.09�� 7M�|P� ���G>�y�"Ob��E {�8T����Q��i�3"O���U��1����t,�7KA�mB�"OX�CR���dq��˂�QMRy8�"O��IrEܔs\.�cBjL�2/$A�g"O�av��,�7�K�4)���"O�a1�6<VŃ��
l`�"O&�0�S
���4!R��ay7"OR��".D�<��IU�M�ttčI�"O�h`��ۓj!���v-�*?{�� "O �X�f�w�p�h���'e���G"O�D Cf���Έ�E��:Y|���"O�u�.���Q��C��bEtV"O�$�CDT�9�!�OI*�H�G"O
����u%z��u ϖdٳ"O̵
D�T�d���1Ea�eg���s"O��*��P�_$T�t�N5@Wj�Y�"O����`�\n�8V�H�a����"O�ت��Dyڹ���
_�J��0"O��P��N)����P��H)��"O��!qc���%�ӧL�Iy��"O8��aB#7���㆜f<Lw"O�)�2������J�eT63���(W"OZ-�� �s�*[���@��"O�y�;]�T#�~�L��"O�s�*.8��S(��Gg�8"O~pb��]-#�D�� ط���`�"O�����&4,Z�CŠT�d%`"OB<����L#`/V�f�8�`"O�(3� �#����FM9-"��٤"O��Z� �$z6hq`&��C�0�۷"Of��K3b-�X�T��|�~��%"O��2�"$/��A�t�6T��"O�����Ϫ3:�P��WA���P�"Oz\��� Cy��Jf.�'�t|�R"O�`B�8�$ap��UZ01T"O
0a%�^�^�\�I!�A	A�ؼ5"O�<�����.��Ȥkr�����"O�M���ƪ1��P�H�2h�И��"O ��E�aC|�g�A �	�"O��2$/�n��{S+ѱꘁ@�"O�bqe�1rպ,���
&�\h��I�O�	YBM]8;Rl$:�L֯x�I�	�'�Axb�+k���Ż%�x��"O�@;�*S6��ɓ5 ��S�싒"O\����2*��@	��l!{C"O�r�AןL�� �Zx�b�u"Oh9���-����k�u��%�@"O�÷}����J��'��1��"O��(c��`������=|���"On�J�i[�s���WG	7E��m�'"Olay�Dȥ{ȰT�4)W!q�Tx�"O��ڢ��nX�1�0u:����"O�*p͖�8���Nʡ1��#"O�912�\�e�z{���2% P��"Oh5Ī[�]��]�Aϖ�%��b"O���Ŋ� ,���4c[Tu� "Oz���B�|��uB�� sCNmb"O`,��@N*�1��	<3��y�"Ox��
�f��Y��0��4�c"O�|����o�����f���*@"O�	����oG�q�q%�?5����"Oz�s`��t]��FԤ{��u���f�π E��ذd ��c�X���"Oȅ�e+�)I(����
��݂�"O���g�Ѩ>����a�5zzj@8�"OR"�a[6V��	��唆c�n�Z�"O�#GE%\ �פ�r(j��"Ovѡ�M�	�̐�F�� }\��T"O���v�A��A����{��k�"O��#"#�<�t!�������"O��#ϔ$���o٠��$��"O�d�
���5�4N�ɠQ�"O���p�¢�
�p��"�>�a"O��P&�=}��%����+C66eig"O:M@��߃&Ӥ�*��Q�Q$�ĉq"O�i��$�4�Z�R���(�0�"O��#g�N4b3��
��Q�YD"ON�a3���^x=��D�R#��sV"O�As�̡#��0�aI�)7�r�y#"O��fn�"���ꀅR<X "O�� e\�^h�$ѺzJZd˶"O��/_�l���s�!p(!G"O�q�dÝ���q:A�N1��E"Oh�c��,���쇼q�iS"O�M��*!Q(����ί1g��*O�����?sҸ ����	}Ѥ��'���"�΍�{��J7�Gzm���'�&d�Fn��W���1wfS
}�xdJ�'�0�[g*C�+��\�6���p�*t��'�6��WEͅ)A�e����r���J�'2N�ۡ��G8RٰRgI��D,��'h(��܀`�"�̔9PmJ�'�4���X�v�F�g٬`ڠz�'��<��h�;Q���S�̝{X�[�'�u�D�L6Et�x׈�2mQ\j�'�(�c�@�?HI[�D���1��'�ɱ�,�;4�	)z��}�'�V�p3��{��x6a�u�h���'*�M��(c�<=�U�lᮔI�'_�L�s�+;s69���6\7^,��'˪���T)�D�c��W/U_��'���K�A2p^���$�ǹN����'!��O�'T�T�T)�D�]!	�'C��w.Tr�H� $HV�H�����'X�S0��!qL:4z�B�A�=��'{lx��́�h���B!C=���
�'4X���Q�WC�5#��P�0���J
�'�,rդ�"D`�ӽ/¦�Y	�'-�Q#4�ޣ��틗�Z�]"�'��R��4f�L����|G��'e���!L40�<����2k��p�'�T�1�D-3�<i���u�����'��ڦE��{-�X�B�LWHxA��'�v�pF
��n��C��]�N #�'�ؙ# 	_B}*<��2	����'��("�O4�n]� J����E)�'f`1 �Ʀ2� Ѣ��D(/.�+�'�] ��I@Xxh�PWn�ִ2�'Nt���G��h��o�8lp"���'���j�Ǆ�d�g� _!v|`�'WR� �.زx��j��Bl����D�'��pav�P4�ޒgX�,��R$�Ix$� w��(�S�E��y���z딥��m��aE�<y����y�*�7c�䕻�O��1\�0w�K�y��S�s���C�I ^y���̀��y2��* P�d�N1���һ�y
� �0e�>]����jH����"O� �'aۜpn� 
�*M�r\8�"O�x9ID5>�z�yՋD�0��QV"O �Їf�
v=�jU�M~vH�"Oh��EO�m�Y� �9��3"O<��@8�q��/�'j��+R"O��9�-�&39z�%�,��� "O�p��+��D�"�#ƀ�A����e"O�d�wG��d�z��0ŀ�;~�,�S"O�� PC�  �z�hd��>j���3"O�ؒĠ��t�R����85��ȃ"O��SS��5�f�J�V�LB"O�ݑc�^�+rL��i��%��"O���6I�w�&���IX�C����"O+S�LE� ���R���
p"O� hU&�0TuD4 ƨc�.�["O�h�ţ_�_傕��F����-��"O�ZE��  2��N�� �6"O|�4J�/����J>��� ��Gn�^�h�Ј�L�@[����U��p�.���~��" >�(��N�)CO�DWS�Բ���@�G�2�*�d�$p4a~��Z1%�|-xesW�Mo�9��/6O��B�jF'U38|b#�<AHE=3�P�i�oG4 �8r�	�l�<�����젠�Z
���3B�Uy��B
hl$PH�g�	wTv�E��[�~��Ƀ�O�5K�5��L���y��&~6�!x�`���tp�Æ �y�Wc���X�C�>�$?��q$�܇0�9K6DƖ@ݮ$�B*�O@@���;W�(-Zǆ��	r�HA��:�@�8e�S qd�-��'�O�M`0HX+8��"`HS������I@�V�9��Y�Ip�Ҧ��L����K98��PK�#$6p;�DP�<Q�EL�/��Ub����	hS�NPj}��Rg��a��Y�p�\=����~�����<D����)�`T�C���p��(c�6��!���`�a �	U�Ӫ:DI�`n0����,_/�Uؤ �<����iC�gaҬ�0Z�Jt�F+D�4� ����R������l�X����(O�|�$B�Z#�p����-I;8���N;��O�21�RP�te�Q!M�us��� R]@% �ݿe�<SK�<"�dB�	*>#6�h$�1k࠘R3-6|�� ��M;���ls��ٳ�����d<8���<�2��*'���S"O��q��զ��0v��+,`n@1�JJdOXe��rfVy9�����gܓ^mJ��B�+��s1�ی!a�?�O0�r"�+2B�s��*y(ұ�@�:~��P�T�5�N��/O�ؕ�#�M1�ؙbD�v���y%�����ቼ ��k��*k֜�'z�y�E��k �ʫ	3�IBe db���	�
��ש��b�8�L>\�Z�'ĺ5h�k�}���'��U#@��P�iQ�ZX��T&?U��%��%>b!�"���f͔ C(��� �J<o,&�a�$~��?��D��|�2����CaG��a�L���#)D�Q&oZ.[*P<!/x!b�B R<i�DJ">���I�/��/�P�*���:9�p��ȓ!������GD�ը���UJX������ԝI��;��DE"��ەm��z"NQIA�'��Q�dȊ��f({ �7lV����'34�H��2��E�a�ÕI��"�'1�<�A��n��0�Ȳ�&��'��B��&U�l���םgG*�k�'�N��NۦW�Rua�VVJe
�'�Hp&��C�$��נ�T$"�'d� re��=U�^|Y�^�~����'l�q��d�$��]���h�U��'.T9���̱ ������$6�����'�2-#pKS�nª0 �GQ?F��'�����EX�jba;3�#V:,`��'�KGŋ�\\�5���_�GZ�T���� �m	t��2VmJ� w
��<�����"O�,h5��mN:�;j��ڠ "O� :`JY� ���:�`Z-�X���"Ot8R�-��BV|@s�e׻l~���7"O�����ތL!��X���Q"O^�� L
a�p��WCQ�	�N (�"OR�bG�G��Af�(N9T�P�"OFB�̷F~2����N�\H�"Oz���C�hp�f'Ks�]1�"O�H��P�$��,� Z�xe�p"O�Ҳć�Rdx%�w�E�'"O���v��&E5��q燬2ЎE�"O����Ȇ�bhQ�g��k�Jk�"O�)�(��)�"+ӒP�.<X"O\��p�٦Iv��4���zɶ�"O����	֍M
��� �%DR��s"O�S�̒��PL� N�,���t"OΘ���=Tc4�#���]�y�"O��ȡ�7f_��G�w~T��"O"h�U�@�x�gȫ^���ɓ"OB��׃L,;�$��tO��Fūb"O\|�Q�mz�lb��݂}�HMBq"O�Ͱ�J�\�"��2f�;�L�R"O�ɓ��R,� �AD�jk�[�"O���&�ݬ%�>�4��@��"O�)�!��P�u��Y,m��2�"O�#*� W�&I:�Ⱦ.dM�q"OJ�Ӏ�B�@�	�$�+�x�K#"O4�r�+L�[��������qd"O��f�Carˣn�Py�"O�t���l��	�߹��)"O�i�0��1��@ŭK\����E"O��6��kd9�֦��&���xU"O8��fKp�h�1�(�~!ܐ�"Obije���D4�dDM���"Oj�D
�{��ĕ�Q��9)a"O$hb��`�n�sӅO�k�v��"O����PY�Թ'�ז ��� `"O,��F�$`���GdMr�5#!"O.��g��7�� �2�
8��Й�"OY# �	������T�b˜3�*O�����@��D�x�a�Xz�y0�'t�y33���`#�"[ib�Z�'x���5-�"]^4xR(�U� 	�' "��9�X�+u+ u�c
�'op�%YZZ�Cu耩?� pK�'����G6К���͉7�ʜ��'�XĊ�d��)�2�����9$�z
�'�P�;p�&'"���6J��i�	�'�F��g���|��4�e�F�m��'3FX�sI��x��`�=<���'�rEs��/�`��Ṃ)6l�`�'F�8fc�f�� a�?Q���'�t���41�j)K��#~)�'qpɀŭV�G6=yd@��<3�'4�0��_	I��a��! S����'9xp�%Ę��q��%Р��'�=� ������e
d`���'�2�l�N��#�h�1�����'$�VHceJ(�W�T/�\��']0|�C�J�h�Z�`IM�H��[�'5��i3ɟ�_4��I\�TZH0�'*�]���!v�5�b`�e@d�K�'w��Ӈ,��z��Ȳ��!Q�M���� ~�k i;o� �zV��.��̫v"O��F� �j݃v��*���"O����q�XT�alP�]CA"O�8H���L�8��_ '�I��"O��[��E�IO* IW.��J-�th�"O4����݃H�"�P�?!v�$i�"O^1i%x���D
�.e{�`�"O�ɃGPcb��X���#"O��)��E��XK���`��D�c"O�+��H"�1+�&��Xe"OVX)��ـq��,	�%ѫV� ppq"OX)Z��[<� @�
��9�4"O<t�Ѫ�t�D��d

�,c\p�#"O�[W���Q��9�/X�Bj��;�"On�Q���VH^�x�fPA)�"O��S6��	6�h��-�84@�lc�"OR�{0���fઑ��.����"O��e(�E��������Ƚ��"OL��A�����RP욂RU��R�"Oh��J��>�-�L�>$�z$!�d˺G?L��)z��p�e�Ru"!�$�0^@DS��i�Y;�GދH-!��]N�,�%�̹?a�L"V�İ
&!���Z���ֈ��}L���NH�o9!���	���j'�ψa��5
Z9B!�$�%�2Y�&Eb��"���-J>!��P�H��� ��\��P�n�8/�!�DE 7$}JBO�t7|U��nɤ�!򄚹	漄Qu�^�&J� ��w!�drHpo_�v�^���⛸L�!�D[4H���@a��`P�B�j��?�!��.:$�z� �c���3�I�%�!�䁭k\i2��tԺ�+���dF!�DJ(3"��"�m�=�Jl��/4!��Ի���h5 
G�*M�Ê�Zp!�D�$;X\Ò�M�7��Lc�w!�ӅU�vh��V'3��Y�Bc-GQ!��y�p�b�ʃ@l�,H��^@!򤘟B̚�Ҡ�|5\�YqKu=a~���:�B��j�怣���/	�d(J6FM��yB�J�ʉ��ꆾ �*	ଋ��y��*	�)r�c
$24�e뤯��yr��LA�T
� �d�c�;�yb�G3y,I�`Ή��$��0�C�yB�W�i��(7A`��n�< �L����vzA�ůA	)�h����H�kMN5�ȓ%W�}��"ӌ jx���L[�0�����Y��b��>��!0���ɞ��dd�@CI���ya�0� p��s�R�p޵[h,p�Uh��B�h ��bt�qvj��|���"	��EǊ̄�.��)`�ڬy�(�Kc��9����ȓ0=4pr�ьLe,��$ޝ*��I��-^����5�0�%KŦp�ȓdj�3�n�6c�d� DC�VnЇȓr�]�� _�m.��P��2���ȓ+�his�ʹ��$��V'<��i�ȓp�&� �hG�d�BlR�	��PF(�ȓw���1��@g��2EN'�x���x��H���1M-�L����;U"O* �5I�i��G�l�bx��"O�e��%_  ��%�6i�"C�.l��"O���/�B�L4zA�,qX���"O.�3�^8����쀅 ye� "O� ���A��36��i�*�3l��"OB��u��5	�J�"�T&\$���"O�� �\���ST���!C�I�D"O�,`�e8~���C�4���"OD���.�1�r$aЪK$���"O���M�7�z��(��=-�LJ�"OT-�����XU;q�� ]�i��"O�Lz2B��zU��X$ǜ-_�a�f"O~���_b �˔�|6��Sb"O���&�LV�Ri2��b�"OD�3��%��I���&����"O�U
�Z�!���D=j,�a�"Oe�U���p�>I�f�Y�/��1"O��rRf>3X.� �!�C.<�J7"O��P�C�3l�k���ޜ	�"O�Y�"L�F�Й
5K��+�Z�p$"Ot��7���t���bR�X�d{Hh�r"OU���V�)�D!;�L\|�ۤ"O�1�ǘGx������).C��X4"OR���Bh�R ё>*�d"O������2��}�	F?@��$�"O�P�ϳ�����O@�A3\��6"O,e��Έi@�|ˣN�+%Jɓ�"O�!��dN�z����S�p"O�qi��i�|l;	Ȁ^R�"O�`�#��oN�ٗiJ0%�}�e"O� �4N���D'�2W4h���"O&y��E-�F��Ȉ�=߶(C$"Ohi��!6z���0�X�2���0�"O�m+LQ�v���8�&";����"O�)-ťL�E�Q�P�����"O�}����.P<T���l�jg"Od()�ɱu�0C��T�]��T�""O̼�cH��zS���$�i8�"O�q ���(�8��A`�HQ*�xT"O��R��*b4H��倳BXY{t"O4Z���5Q��5�Ć�4u0�]��"O�C�"ơw���0V/�.� �Ô"O^A��'�hd��k���t�D��"O�8Wb��6��,��d�;����"OL`��	�F�[���O���a"OnI�5�E�|�����ޑ�P"O
��G�Z�I涵R �&�z��"O�$�m���=s�"�����"O��JǮ^�:�>��sJ¯o�|�I�"O���c�[\>8"��S@0�� "O܁!ф��AuTqS�U=��5yU"Ol���Lߡ\Q⌊�l�"Ή`"O���OP�2�h�+אqS�t�"O����H�s̍2�,V5n!n|3r"O4�ɲ�N3fo����@��=+^���"O�E�Cj�(���b��S 
� �"O�D��&Q�U���w�Lyb"Ob��e͐n���A�-��J���"O$Z&��'l�}sr�Ps,X�_�!�d�2�p%+�ar����tɊ�0�!�d�--��9�uُ0�v<Дh3#h!�$ç;��!3㇧Q��l2��p
!��T�
Ip0��6e3�͒��!��fV.�bG��/����X�(�!�D�m�,i[�M44Z�S�iU�f�!�Ž ��ad<�`J�<�!򤈔C}l�T�
,���@�CdI!�d�j�Px�b� �V rB.�'"!�� ����Mv��t�D�>0	�"Op͈�����I�I��Eń�R�"O.U�P�N�܉Jsh�o�La�5"O�;�'"3b�ɔΜ� �d���"O=n឴{���:���`�kІ$n!��J� �su.�,"a��dŜm!�%"8K0�a����W)j_!�$�%}����LK�$}V���۶K�!�$õ؈`����'\����[Q�!�pǶ�����-@GH�p� ��
Z!�d3Y�<X���V�`HT��/ �!�d��lt6��^(.�`�кX�!��ŬI�L�[�.N�F��Y����(<q!��C5��2�U��M�G��UX!��'*.m�C�X�_��D�PI"2!�D�6H!��#�f�t�QȔD�!�Ē�5:���KƑg3t�PR�ª7#!�$�@/�d3"@�"b������u!�$GM�8i�R/A=4�\�c&��!�!�$V9S�\�	q��{��s�$I��!�d�5�Zh��_��h�7�a�����H�	AJ��&��C�W����y� �5@�:-JcIL�M�m�ȓ�\-��n�
�⢫��ɇȓ^Bf(ۃ�L�h����u�V�N@Pp��,�N����Q�;����t����ȓ<Q�����k�艑����ތ��}3r��Մ	+-p qYX�7Lʕ��Y�����`�-$^9w�H�V@��A��[�nF4&�2)����ʘ�ȓtϢ��%� ��(AWjE�-|*u��OH�I�@�)}�(�fONO��U��;���S'��~��ǀ�hh]��H[���a��/K��A0��u���ȓP��A�D�"N<ؽb�";kx���%Y���V�*E��#��׮<�fm�ȓKD�ԍ�0PjH���D)^��Ԅȓ_��4j�ɖ�� ���N�r��J�4}��G�.~�Br��?/�*هȓ{Qr�ł,�h��@W:	-F��8O(4�ꂔ?Kt�'���1C$L��M�t�y���1��9��_7��ȓ!2�����#!xB����	�h��f|����C�6$���}@��ȓ
Ȃ�z`��3+��X�9� ����\�Sq������C��\�ȓ<�Q��B�~��ia��J\}�ȓ	1n��#C��IB�Kә62�l��*>���Īf���#�ΐ~���ȓUt<]ʅ�Q'bz�j7,�7�u��gI�YC�
TL���1�hĄ�!i�l�T�H.1�b�J�U�jUf�ȓp]������)�ቊIt�ȓj�*��6f�c�,�C�� �	��Ks~m�b����r�%>d��a�ȓ)�t�3`ܾȾ�F��>����Wt	hS�O�_g:��F�-�����U~t���O�=�W��D@��)�;�c�k�R�pO*J8����MG��R�e�j�s`mӦ`,�ȓU�>�`�L7=�����B�I���in�����D�W)�9?�܅�ȓ[z&�)�.%q���r�7[�
��ȓ>��f�V� ��Q��'�&��S�? �`�KL��D�a�\\1��"O���wm��u��ؠ��\�P��"O�@ �&��L�d�V�N`���W"O6`�ph@i���B�6#@�@%"OD��4j�l�0xXE)��|;T�h"O�#
�=;���C	��j��"O��r���"�t��uI�".���"O�3�H�rbñ�H'/��[�"O��'˘�Q x4HO9C�a�R"O�(Z�	Oh�ؓ�h	��\P�"ON1��d��-�Z�Y���Ke4�*F"O��E���}��`�q��&b�p��S"O�<Re!�"
�P��S.	}^,B"Oz��Ȃ0�:9��D\p5��"O0����]��J����3"O\L*jߪz�l�sd/.r��H�"O�Y��%�t��ᤑ�!L�)&"ONd�H�?*��k�-b8iz!"O
��®��1��#��Z�I�Ԛ2"O:u�V�͘`%Dm�F�"�� {�"O-�tB�m���2E�q�� �b"O���@̅��j�9�`�<�"��"O��	v�A3q��:��Q�}�Jm�W"OH)��#��ܢ,J�>�f(�`"O���Dn�?!�2����Z�T�J�"OU�a
IO�xS�թ1�"y�4"O`D 5#�~�pHSM
7���"OZ}ca��e��I�6	�v�C"O0|��۳V;���#�=BJ\!�"O^-򡞺k��@�%Ÿ<(xX[E"O^ ���ȏg٦0 3�ڭ'����v"O��"�ʁm2��a)�
3����"O��@o�n�5:t����p"O� �$�ؠ4�lz/�1O�Ȉ	�"O��95��+'�8rϏ�\�L�)�"O �(�M�N��;6LP�W66�x�"OTPb_�=@�#O�jAp0pE5D�T�5ڟ/h $���7eX�T�9D��`�K�����@���l1D����T;x����Q1P0�Ҫ1D�@�#�����+4l)X�P�#�2D��c@�Z:h@"�x	:U���!򤄴g�n��'��\��`R�_�x�!�d�0�:����n�fЊwÝ�O�!�dJ�
���fY�m�ؔa�)�M�!�h�0�qV���^�\`��I�+�!�
��V,K�gD!Z<���T��gL!��Þlw&�"�W3k̬1:�'�8�!�D�9/8^]��hR�[�FYQ�Q
!�d 8&�bA�D�!�H�@W�!�$��W���PU)�%t��d*���!�!�dG8��Pq�*�Ԡx��� ?�!�J�y:��7�L�U��ɹA$Ɖ6�!�䆕H���$�-7������Ti!�d� b�찠iK%d��L�����VR!�d��Y���[���Ȱk¥	��!�dY�{]^�sb-Ͳ�^,(E]� �!��T���B�S 3��c�!f�!򄈻L�T��'��Q��a&�ؕD�!�d��rX$aH̘;��E���0�!�䔏�BLp�EА�"�
!��)�!�D%m)&ĕk�H%3&�L�,�!�d���*�
6+Zn�5"T(3C!��ǹƕ҆�ӴH4<ܨ��ڝ4:!�� ��
�'��Z���e��Sb�E�"O�-��#�.W*���(����"O��+ m*m�������`��I9�蝪� N*� M"1a�%vђ�D[�0��
䌀����㯍3fqOX����و3�ȁ��E�����3lݢ�	ٸ_��#�$K�;���\�H�����D_)�0|�ϒ)>�zy��kW�]۳��P}��[�X��\��͚EV����@�.� e�=n��-�H��i$^�#�F�XzɧȟVhXA�V7w�����
��"��C��jq{O>��O��QJg�  ;��:ui�hv�Y�}
�v�B���L�0�a[A�O.$����,ٗ5�'I${'`9�)�S>~��A�c� �iZ�'E,����XV��$w�X�4'��I��>`6�ΔK��@�>E�TH�-g��tI4P�5s�8�N�;��z�}�#��튖U kKb����:���F�d��LFu+çm�J@Ԅ� �"6O�V�:A�O�)ULބ����O�R-3Ч���<�diƻ`-�1��'�v�p���e�S�O5����F&x����#H.TC��)V�1(h`*�}���9"���q͜(M��H�����"���+R��Hm>��Cc�=���5E	�\���5�	:��<y�'@D��8���E�`�K��h�x�&���*��ا�O���se�<fR5y@.\�~� �٬O�5《�C�S�O@�0`fJkr��+9s��,�޴�H�q�T?��b6'�=j�eUX�����J��f"}�0N;�d�v>�&o���f���bK92��<a�O>`�Mu>E��f�5(�Z���_ХKĨ<�\�7�.�C��y>5�p�ۊBNĨK��>D �٨��>y2f
F��%
��x���$[=�e��=���Slǚ���J���jnY��٥D�
�8�W�h�<�W�Q2|D��K�d�LY	�Kh�<�w���`���n�x+0�b�<q���s=�ě7�J�|[���`�<C�
x�,�F�İ#/�I�EE�@�<��/Ƭ��t��۩O�S�)�@�<`����C�&��E�M#3��{�<i�c�o�jMi�d6�܄�wM�w�<�f�]�䠊�-d�ȓ6��.x�C�IJ-`�JM8K�<88���)K&B�I�8LJ�V��e%($c����0�B�ɇs;4�{b@R  \-�#�D�i��C�	�l�b���:<����3I��C�ɢ���Aآ7of��E�_"8(�C�ɭH��)�k�=^�4bs�J9��C�I�:�@�sa!�58���N�I��C�I
~>�x�s�nE9�wML1h$�C䉲W\�<˥��A2��t/�uЌC䉀h.HϜHrV.�*��dB!�m�<Qw�˷C�Fx d�j>���en�c�<!"��6����e���f�X�<YR=�P @0.G�l��Q!JCV�<�ʄ�6�&�@��H�2���'oHS�<Q��8t�Ќ�D�
��<lp�Y�<)a ��u��8��Y~�� ��Q�<��L
�\��D	0���kRJ�<v(Vb�z�Ђ��V����F~�<qrG]�#��8��ѩ }�I�3�S�<Y�4ij�ɓT��*Eܸ񔪆L�<��ϴX� ��B0G���A�]I�<��˦<�,p���G)+|�×(AI�<!�UP�6=���CA�x��M�<�D�� Z ��f,�
I#�&�S�<���2.��RѠ�V`9#�z�<�&L�T��ˠ�C%c��i@p��s�<Q���7R�����܋T�dp�&�[�<�J(;҈���0.�h��v�\P�<� l�{`lI�S� �d�'_+���g"O0�@Tm<
P�C#��:�E	�"O���-�bgơb���B-4�B"O`|�;}�F�PeG�;�K�'apt�#,D�,t6A��&�J��9�'"\=��"���ҕ B(Y�b��'꜡"��>A��*���L�R}��'��M�C�T�)�>ؓH��C�f=x�'�>u�����k� �*l�r$h�'��]iF J`(��K���i��%�'p��t�:Z<5�!�iP�qA�'�t���ѥ����!e�w���)
�'��14�%nO�16�A>p	��;�'�
���M�Z�$�%���`�
�'�l\eO.F��;��J�v���'��Y�Ы\4[��g��& :b؛
�'ZE!��P�>PY��C�|�iK�'��T	��Y+[��)�L>S8�0�'�ly���Ԡp��yK�LJ�9P��	�'y(A�T27+Բn>=�6%Nt�<���Z��Y�B4*�.X�5L�m�<�DAЩ���2n��u��.Ui�<#/��e��}�j�sUfpy�e�<�EIy�b��"���{���%�l�<Ae'Y �4+�'�&S�����o�j�<�dF�^dcLBS����i�<qT��o���AEJG�$t���o�<ar�%c�D���؊].���To�<��c ��5b�E̞O�pH�@�<��̕*���r���hݛ�	v�<��k׮E���Z�˒1gf�Kv��o�<ѳ��;�u�CN�e�h�<��^$#$}�7��Vwr��#j�f�<!$
�E� �x��H,8���a�<yԄ�0[�8��$_�)Ҟ�k���I�<y!�%r�m�աZ�MN�%�p�D�<���5^.Ѳ���iw(�
@JFE�<Quϙ9m������Kc��,���J�< �g�@MH�*V�m�z�����k�<��C��v�X� +(t�-�n�<�e�!��4J�<@3c��f�<�6`�&[�p�@-�Rv��v��g�<�Ǐ�T��Y2�O��8  G�c�<a�Nۈ(u��m[KLe�d�F�<�q��U�wC��=��`�l��<)�Jˑ����-�o%������<a�@�[׌h�O��6�E�W�<i�H>W�d�j�N������/�}�<I�U�b����$��(q��L�ш�c�<qCh-��d�� %D��I�� ^�<�@
O�Rl@(􅗣H�<Hc��D�<��"�Bq�3�C`��"�g~�<9p�_�E3�1JC��m�65wf�o�<�GDE��@Ig�@5he���i�<"lΘk�4��XsLT�2��P�<�5a٨Tn�1iŒ�.,2E�b�<�`�ڒj~�����		=������H�<Q����<h�!�-��i��gBC�<9�n�;�*H���*6:�$i�jAe�<�w�ۥF� �n�-���FE�<�HT7'�d��ǰ/(vစR\�<9�I�D6	:&k�G�8 �%�T�<	2�Gd�a�CA�*%s�L c(�T�<Q�gغt�f`{$(ݣW�< ��h�<� ��)Ƴe���p�:\�0�qQ"O�}�0��?���TAM�^�2�2�"O��&����N�D�+B�O�<�p�RR	�Q�V��F��g�K@�<�тQ(g����߳t�"�)� F�<Q�IC�C@}����� 20�8�AD�<� Q�tO<!j��$��@�G|�<I�Ó�{� �K`�?�(ȣ'u�<�E*!/T��"��������[f�<�Pↆ7[���saR�o�:�ВB�d�<A�nR#_�`yju��_	8���j�<�a����"�h� �z�H/�^�<1��M%�|��L�-�$%X5�^�<10�]k�BBj� �^hԏNY�<�p�N���Wo�=XM�qk��S�<�A9����`;z�����I�M�<I�%B�V��sD�]�#8�u�1E�H�<��㒢�3EC	�q��=`cF�@�<�'Ɖ��h*�GJ��#&��@�<'E��Ϯ�QׁQ�_B")�#�D�<1�`�W�� �
��-,=ѳe�L�<at�5G�&8�@�R�*y&�ۧ�H�<��F�v̆y�l�V~��*I}�<A!ȓ�P�8�[`�'v��=�R�Wu�<�t��+@�����:R���c�/�[�<qr�'U��ab 7�4��'��Z�<�lF�E�^�5;2��u�VY�<!�g�'�P0�0`P�A�q{vm�X�<��l ("B�Y�2j��=n�U��{�<a��s�lٰ��� ��Pjfn^�<�nZC�
y8c̟�}�9���c�<�$�����Lزc:`�&�I�<��(�
9gG/0��Ht��D�<ѓ���50�� %����7NA�<ҰP8C�1[�j� o�h˄���q@�(�φd�������Qev͆ȓ���D�F?W�0�2ٚ&����L�V}�"E§I#�5P!�;e�
؅�d��A���*_�����ݎ#U�B�I�gr��2�n��U��n �N*�B��)&�����!@�XŨCh��pB䉽V�~���nM5f�p���&�rC�I�l��Jb�]8_�j��ƂQ057tC�I�&��ո�@�h76Y�T��5]�B�I$Y�\��⑶;��qv����B�	�[KT����Dd1���2Y>B�0Cr��CэѼv��h!�܏Yt�C䉾 �lQK�
���\Ґ�LVA�C�I�T~y1		�<��AEN/k_B�I�X��P���q�v���H!Q?�C�I"T���w�P�>b��BnG�i�C�	�x�0�F�
�hqj��G��B�	�K�f�*t�Y�T
@�s7���H�B䉗88����-wg �� ��lڒB�	�b�̢�+�	��t�ի���>B�:a%��� S]A��P�Ȁ�wB�I-$D(�y��ݬk&����<8�B�I�fM8���Y�S�~8�0��8��"O��x1��& �^���Í�F���C�"O���K]����7U�)r�"O�q����B�Ē8���ѧ�#!�dߏCE�%KvI(�̹D�Q�j&!�$��z�D�����/8=��A�b !�4����p�M7z�Ê�X�!�� 4yY䬙
j',8���>�j�q�"O�J3�K�jTN��V��;B����"O9�g���U�
�@��k(��
E"O4<�LK8XJ	Xf�G5?@�2"On�Hu��,2����@١F\=��"O�`��*D7d��]c���..7Fm#"OQ���j`씈R�\�#%���"O~�P�����p�`��٫�"OF��$jR T����P*ޮ_�h�d"Ojm��B�%76�\�E$�<:�}�5"O2,��Ć�z|���N4D���"Ob�S�
�`[�W/�劔"OΜ�a�S�\jz���3!t���V"O�휏$N2�ѡ�"'vXQ�""O�@Ж-R,!�@X��-Y=I}Rh��"OT- ��E�&d�W�[3t~�y�"O�ٚ7,ɹ������\64f��� "O��@��S2/�ޘA��؞C3���"OjM�4L;`�Q���m��2"O�9��h �p���9�-CH��!:v"O\!��ˆ|B�]�A��<&���r"O੒�)U<Iܭ�!G*;�v�"OD)��в?$,D ��ɀ.����"OVdJ�(ׁ ���c
*4��郖"O�xY�BƮw�*<� m)o
x �"O&�8���K��]����\<�"�"O%��+%�l��jK�GR�$@�"OI�#U2igN��W*�4(M,���"OJ��D��XH��:3ʅu�b�cW"O:J1�?b��QG�O(x�����"O�'C�"�����[�1_HR1"O�t�3nվM��OSm�P���'�bl��� HoZΟtn�v��S��/t���+7�S�TE4����?��;�?��?�c�޴��8%�^�Q)�Y2�L�T��y����H������A>���пrp�yFy�׽~1&5�Ԡ@&pa���PGQ���ɗti*��a��Q^�9'bӥ_�@�Dy2HD��?Q��il�	Ax��ע�A�cr�����������IC�S��R�4Z��6`9c���r���Z7�,�P`�h(g��	0�R����+1L�>,���޴���#R��AmZ��$��K�d�;�6�a��!��Z�k�0�a�%3ocl�D�O��)e�F|^��bZW� ��\��l'�~r0J�7a~�Ӆ��<�X�9�bM�I��	c���* f�) �A6qÐʑ!]�I��;x�L�P ��U�h������6�DO��8��'��8�7�G�6�U�.����D
�7rqO ��/,O�R�/^
y�5�#�	}��`�����O��oڮ�MI<��I�/B|�����?P��XSF	�F��7m�O ��OZ0�ɍPR����O����O�D�vN��ab��z��(E���0D� ܴaD�|`FI�
�*y���p���O_���FR�?1`��!^$�;�A��k��=�00&p���"L$Ch�h#�7?rAc��:��S+Wy~@[�w�5�6ꉋB�.%�f*RXY4���D��,O��������?A��M�f��g>���]�P��2�"� Z��'���ȟD��'�+�@���#%��4!bĠL�أߴfқ�|��O,�W�*���\�P�k��R�c��H��ѠK70]XR�Y9�?���?9��S���O����O,��W�2!uz�T�Op����gC� #1�)s���5z10�tSNBF�A�֨UQ���r`��c�nX[�����w��)PYK�
ŭO�����)�3A	tP�&حs۶"<�U�M$\�ڵgٿj��4�WF�2&7NP�I<�Mk"�0}b�'���$�=���K �P�6l@ۇnI�:���	p��h�f�Jq�ƈ^��m �ƕ�Dɖ!0aVh�4�?���ig�6M�|�%�=����'�Vo��_"[�Z^g2d/�����$�O�Q���O����O T�/J����ƨ#��$��)֧]�,��jϙ&f<#rd^(�b�OL��Q�`��*��64�q��1 ��}�g�C=[) ���C�(Jq���Zr�H���@vQ���aG�O%n�!�~��� �0� �17��i��H��'�a{"�}�.�1��ݺ&��ŦI��	|y��,�?�����i��m	�ԶA�'�@� ����'o7-2!N���'��'��Ġ���G�+T�� w|ՠ�G\
x��d�O��x�`S�Is�2{^�'�@|�q�a�~��Ά/:�LS��غ��:0��~�I%NFΔ8��^Nоhx�B�Zp����B�Si&�����w�C�2h�/ڥ�m'�`��A�OTn��M���π \d
�c[=,$�H F�.X"��3!�D�O��&�D�R�T�j}��[&�i3�x��+OT�mڐ�M�N<)���>H���q��8|���NO?I�����O*,@4�  ��   1  �  �  4  +  .7  C  DO  j[  ag  is  o  �  ��  ��  �  N�  ��  Ա  �  g�  ��  ^�  ��  ��  l�  M�  ��  �  Q�  ��  � +  1 r! �' �- <4 <; B VH �N fP  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��	V~R�>�,�T��0`��,ap�0b*�W�<1A�Z%PV!р�TCM�-�#�XW�2��6r���=�O���2,Y�vg��B�@+W�d�
�'� 5iWڙ2���*g��Sf���M�˟�>E��B�Rƃ�/�V�	�D�}l� ��	P�YWly!�+�?M|�\�p.@�@=Pq��*!8ي�S�>W���cW.1zZ��ȓv�MP�""Hd�A�*\�D��ȓV���.�:���x'�Z&���'��#=E����'dAAU�	��E��*
�y�K�r*��R � (�YDL�;�䓱0>	J\3x^���A�!4�i�uX�4�<��'�Ę����:��u�Qi�6v�5��'v�:! �.\r��N�C*��
�'Z � ��(s��ღ%4�+�]�<��=H��Նx}�Y�2�c�<)���4[���̀0�dk�J�Y�<��a8S�YbF3�ȸ�bϙz�<	-�+Ld���g�d�^1da�u�@��jL�h�u�I2u�l�b�� �����6D��Y�O��0�>+�Hi�"3}�xB��G�b!BwAĘ&~��x��~��B��	$�p�H�I�hp��ĩ�K��B�2�� H�M��t��0�ٝAʪC��>x�1��;�*�X�X�0�4B�	N� �)�΃*I������	K,���(�� j1c��G��ؙ����'5Z"O���� O� ��mmϤh�ց��"O��C�k�+;���{s��>�4=Z�"OJh @�K-���ò��6u�l�"O0!��R;.�R}�vI�W�E0"O��I���*�M���\�pQ�p�F"Op�R��!UjzY��R�O�����'��'�*����5��ҡ.�A�� *�'�b���/Ţ~�*]Rak��;`� ��'_�f��<=�*�i$���l2�'��TR@�
%s�*[2!��X���hO?)��#l��t	e���=��fEr�<���?�@��*��qk�X1$�c�<���ǜ�LHFn`�ք�MI8��'��J�ʎ���m�4��bhe��7D����������&������!!6D���ë!%Lz�F>����2D���b���o@,{?�T���F�<��V ����ԈՠWzq��@�<����?���H���^�0�m�z�<a��
=k���sg�/Tָ#Umt�<���6٪�x�nI8D�� ���f�<�GA\C�|�'`سb;,��plOa�<�"_��$�$�/.Bvxa�gV^�<)1e
.��� �ş+�j�����B�<����@��!6������-�|�<�ℓ2-��Й�ŔYX�-9�o:D�$b���oF�����S>���;D�|�Wl�:�8��ŗgu�ȅ�<D�����M! 9��g3�&��`�=�Ո��=���g�����6O�ȡ�"ONm� �����#r��->�
芄]�D{���I.R�pm�/��oI��J�
N
4�!�X�*�� @�G;s���˵�:��'�a|BDT.mA )��T0Gr���NϽ��?��'b*�K�߷d��`�#l��4�p��	�'_Tↄ�f��Y��mV�[ƕ���4�']��P�H�j�eq��.
���|�Τ�'��0�B`�/Ʃw��܄�zV��c�IC�f��)� 2Ǹ��ȓu��H�h��P��Ո懟�=Q�t�ȓ�P�hE���8L~y��ǻV�P��ȓ��a2L����is# 8*���HSH��s�T�E��TC�$��IT����\�XX҂�?T�Q�� H7`��O	R,�e(�/V�Va�#�*�t��c��iy$�P�9���@�Z�Y�0�ȓ�b�PJŽ,}�qh��bzQ��kq�k�ړ?Ԇ�q�!��|�=��xT�uJbT|�~�5�� v�0��V��qC����>z�a�è�;�����T�����ߞ�����AP��/3��:��0�TLbd��2rP͆�y�XQQ&'�7��q$�W�3rXU��w�l�pC�M7��I1�0���z=zu��M:K�^�Y��WXXT�ȓ� �00�[6d��\�g�/rҁ�ȓ
�8m�5Í<^�u�V�����ȓD�J�[Q���6��Zwm�?'¸��\��� �R/Bh}�TEQBV��Hx�`� �?���C񤑆�����,
��M��m�昘CX��ȓ[�j��Fѯ!zD֤\�<ńȓ3p>䳁���C��L�5
N1���S�? &��u��W� Y�	\97pN��g"O�h��G��@j:T���2KF 1�"O��X�+)3�V�W�Z�k��-�#"OQ`��Q��� e�v��p�"O�Y�!��2J��D�I
Ұ}b"Of9��
�+�xc�N�@�D}#D"O�IA��
GN�!@2%H8)�Z��"O���숁�*,���9j���Z"O|��m�1�t�JF(��hs�u9%"OPuS�� �[�V�Qlʽb�6�[U"O��	a �<x�E۲-P"r,}*�"O���.\�2��0��ݕ@T�q��"O��� )FMA��82L8�T"Ox�g)l˦�EZ�{l���"Ov� `�Щ_G�4)��I�
^����"O� rph�t����W�O �"O�iCp��+���BrE�n~(`�"O<�Y�hݶ�:�`����T�D"O�(��(ȫq���94�L��lk�"ODt�A�����]I`��n�ȡ"O2Q[��1;V|�(��Ut��Q�"O��� ��dl� �ϖibP���"O�=�&^#rnݠ�ϕA^� �"O�JC���G���#�ʃ�R�@�zU"O�ЃV�B�#�Qs���v�x���"O��@fc�m���Rd�֥,�p��"O9+��ڂk�ysr��&���zW"O�g;Eh ��Z�]��m�"O�5�	9�B�:w�E�9Q�0��"O�Ezf� UX,A��� ?�ژb"O�������sC!�4��9�0"Of]��o�n�A ��'�@��"OJԠf�=#��&@ف@zYi�"O��P��6]��P��q]��c"Op�"�c��V*�t)V�RK&��"O�0A��)j�V K��R3*�␨�"O�D���u̜|J7���hcT�t"O�Ђ��2I2��1U)��u�B|�"O��Xe"Ia�1҂نl��ej�"O�lCp�בdm�`	�A�"�vx�u"OX���8m{���R�B�?t8��#"Ox��uF�
c��Y(�/�.�
�h�"O余toT�Q�|�ʗ���"|�� �"O�DA���f�^H�eA�,be�t��"OD��5�J�~�Jt�pX��X�"OJ�k��Q,9�b����ME&���"O:�0f��"+Ҁ���S:hXٰ"O���΀����Rf҅s�p!�"O���	+��U��u
�ēU"OLH����7��-���'o���"O����Wt��C�'>�8Yۖ"OV���]����b6��;`�2�W"O�!څ�ڝZ.aC�:�@yH�"O�@�!��' �XB6� �h�H�"O�hJsHZ>vE�u����$l��"O4���Ѕ^7.	���W�g�^Es�"O�(�CZ�m���e�;pޠ�""O��(��!i��3�؆8�*Q�S"OL��$!b``HC2.�/Z��1'"O�\����h�l�锫��4�K�"O\uj��O�$�8��d_�q��h &"O��a���1���P��Q�y�.P��"O8x˳�� A��(�$�[+u3�d#�"O6`��mX;6�Z��#s�T�8"O� ��!�@�YK^��A�@܋�"O\M^�����#J0 
Y�C"O�0��2�!K ���;J�R"O�Q1g`@)y��̣%.E�7�|87"O�@�� o�����ޯO$Z���'��'!b�'���'���'+��S8;:d���E���S.�ptR�'���'�2�' ��'S��'~�D�$)�k� I�5�����PGb�'5��'��'��'b�'M��G>\'t\HF��Uh���rd��'2�'�2�'="�'~B�'nb��+'uN9z�-ӥ- 2�s�HV��'���'�R�'��'vR�'B i�Th�b�Kn���s(F%3�r�'6"�'�"�'C��'x��'_�k�(}{Xq1����ED�0J��ɗv�B�'��'���'A��'r2�'���ϋ����ՌD�0dBWŅ�vU��'�2�'^r�'��'q��'X2M�29�8��M�#X�N����ڑO��' B�'z��'���'x��'ErM�>�rLk�)C�-	â��w���'�R�')��'���'xb�'�BL�;Ũ��c^�
CP�z���5�r�'���'�b�'$��'�R�'NR�_Ä���C}P���@�*�2�'���'"r�'�'��'e�MY�[0L����-a7n�s&�P�k�' ��'WB�'�2�'�l6M�O��D�4u�)�-�r��i!��^y�M�'	V�b>�r�fF[�,]<�Q�@Ţ4
��*KqV�M��O��oZh��|���Mۖ�+ ���֞h�P��ٯmț6�'�29�B�����`�@щ�����u
]@R*R7_o���PE�e�zc����_yb�%��鷪�+kڸ$b��
tf<1��4.�r<�<ً��|��=�ڱ��/=V�!�2>u���Iۦ��������3���ў'|�]�R�_�$�1#$�7U.Tpz�'��U���FʴS��i>��Ix�HB�b
���ZVl�J�D��dy�|RJvӐ�8��קZ�f��po��T5�%-ҩ1r�(Q-Ox�$q�~�	j}2*܁	��h;!��1H,�2V덳��$ù�Z�3π�~�1���VJ�g�D�$ʝ`�\��90��2�	Y�Šʓ��$�O?�ɾ�0$sЯ�1V���4N��P�?�M��X]~�f����g�8Aq�b��D-ѩ��$��� n��8�4"��g�f�B"�:p@�7-��q���X`�/> �����"�hO�<�K~�*;O���4o V9�$�a~�*}�8����3�S/�̄)�AU�|�&�l��X�*OV��k���IT��?A�Ɋ,Şt�A��r*�p �BB�U�V	SS�����������!������.}��5?q0�'=0d��@A�]8���E��?�+O@���G�����y�-��>�)�)�� �����yrEb�>�泟<��զ!�I
3���pr��<AJ�+�k�5(w*x���'���	02����rJ1��PB؟��)~�QJA��,H��I:��Q8V��G�Pt�S7O��D�<I)O?�Q,��-{��O���Rpa"扳�M���PD~AlӞ�O���`LңAf�S4���?��(Wiz�4�'o��g���$LwT�S�;O��hW�ۻc������ǚ;Q.5�U�*�@��!(B>x<v�!�2�0?ͧ���O�[$	(N
u���x�r� 8O��Oym��qy�b���OuR���#�O���
2E^�wd0p�O���'3��i+�D-�����p"bV+|�h�����*�Z�c"M_O%� kF�Q(�i�֝c�!*�C�u�I
E��q��(�3��2�T�I>!�I�h�'D���X�|��4~���3��п:��d ���"q}@�)Q��|~2�l����$��Z}Bhv�dA+tB��v ��A�:c�ia�����j�4-FZt����<��[m��`��Ab��AK/O��M�97�������xh�L�#8O&˓�?Q��?���?A����ǯT� �����|d�����D�#f�n�)��	՟���O�s��������B��&E��H���egv���%Ɠ��nn�`��IX}�O[���O�.�#�@K�y�WZ�\3c��rtA�I��yr��$�X£����'�����I+n��Pڵ��ڨ9��$u8b<�I�T��ӟԖ'�B7�Çgi��d�O���+Ob�!��=8Y��	p�B��P��O�lZ��M+��'~�I�yf�Y�(�U�	���t���	��8�+[�g�ba�qy2�O��e�q��}����3_0
Č�(k���/B�z#��'�"�'�B�sޑB�����1p�)ܠEL�b�� ��4������?�S�iL�O���>6�
\2#Gǭ9ӆ�#�	<j����I��4,�&ɍxf��Y�'z�F�+��yz$��:Bu2�Vk���F,��'A�ICj(�|�W�|�	�|��ן���Ο{��@�]o,)C��� >j:!q��xy�Ob�f�A�I�O����O��I0�i�>^$�	�O��&ᒰȘ>F ��'zF6m��������'�:�'��	0sA���h��D�1)�2��fʚQ��*O�X�"ٖ>NY��%��<iO�d6���&D�1g��u ��?y���?��?�'��NߦQ2�Ee��� k��\,��q�d��|%�%�u@e�ġ�4��'�r�/ϛ��q��`l��6kh�EX6P�"e*ʬ'a$���1&_���,�z�Ǿ$]�H�F��<���'` �X[� ~(���
-��R��kB���S0O��d�O���O0��<�|�G�h	P�0���4���@�\�<����?��iTJ���O�9o�ןT�'i�]ssL42���+T�<�A��O����fe�����'Uv�a:�1O����;@`ק��GV�Z��-k�d*3E�m(h�(ړ�?�/O��d � �v�@F�6Gn�� ��HF�D7��ڦ͠5I5�I�?	�Ӄ[�nC�ԕB���ِc��F��	ɟ�n��<QL|��'<`!���9v�&uy$ʔ)Dz��̳&�bA
�|~b�O^*T���$y��'n�XsP(�/ f`h�Ʋ@~B��V����Wy���O�hmZ�S�����\Ԧ�2��O�x��095�,?!��i�Ҕ|��~b�i�<m�ȃ#7A�E�"#^��v�s� ���9k���B�>O���/i(4�WB�]F��7�T��6BV�w�&��Da1AM�b���Iqy퓆p�������Ŝ�<jT2�����1衏:���?�$?��������U�ܸ�� S�,9 U�,;k2�i���<�S�?)�ɬ �l�!S�c����
:xM)��6��!��r�̡�n��A��9@#�\���D�'���`��˓Gkz�k��J�zl��'��R��;�M��#�k���%����n*���gQ�D&�*�B"�<Y���M�'K��(i�	����nL0�ꠣ�b�F�I�����郟D%h�
6�!?q�'�F�+U�?���
d��A���~�L�#$��?���?1��?��I�O:h#��ԫ5
�8S@��^|xzW*�O:�n�65�cכ�4�\)��,�0U�6�s���4W��9O��o��M��iɈ��ff��y��'��yɓ�:b�Rv��b�����E%������r��'��I�����џ���̟4�I!p�]�e�Ob8TK�@�])�m�'Z
7�E�eV����O>��쟨�'�?I� �$m���1�Հ+���TE�I���M�кi���D ���)T�_��H��kRD�;"F;8�� a�x���I1��Pi^�"�&�ye�xr�<a��ƈUQ��J���Z�e;�H�?1��?���?ͧ��Ц)c��럜iA�N4RSX�Z��l�5!��ٟHݴ�?�K>�FZ��۴/�F�eӰuő�11V\��e�8^h��"�!]���9O��dY�\�RW@�<r1����ƹƮ�e�S!)��; ��u궕�P:O:�$�O���O����O��?a{"�X�(�I�jB�5!ʭ�v�����Iݟ̋�4q�
��'�?1E�i�2^��p!DՋr��42�� Z�ĥi����?!�Oh�o��M#�'o:}1r"Y�<I��.LⱯFp����B�Es�5+����t��P 7J��������O����Ot�$O�z9�Y$͛�#�jI�De	�8�����O�˓>��͍���'���OY���#/����.�n�NHÄ�:��d_}��y���n$�?�K|J�'f��Z�oPX���V�W$X%��oZ�Ew.,x��6`��I�?�
D_�Q'��2��;g���!$	f��Ѐ��0��Ο����b>1�'�87M��))����)dv��t�Է~�����O`�]����?�^�Ȁ�4#�D���b�d@�s��oW~�� �i��7��JTf��s2O���IS&$�SDϘ}�j���w��)}�X��*�'`R��A<O.��?!���?���?i������D����1��M�2���߿<��o��.�	���	L���wbh���\SR`�vN��U�Fٹ#�o�9lZ�?�O�������ΒF�0���=O�!9c�}�Z����<�ޤ)Q7Ov�� 	ϑ4Ϧ�k� �D�<)���?�����2�L���y
b`R����?q��?���������
D��8����8�B@���- ;�F(3u�r����	��M�U�i���D�>��7q"���c �h},@!b��<��6:�]�b�֒GC@e�)O��I�
��ȉL_b��>N����խwE$`� H���'q�'72�S����)�9=�\5@7lE:փ��X۴"��S��?�Ӱi��O��CF�VP�P	�;��{�N�a�d�צ�۴�vM� �h0��'�d��P���c,9t 7Oʊmo:j׿G��tYJ>a.O����O��d�OL���OܑBd��(=���v�ͷ�����<���i\�E��Ov�d��ڒ�HUzՊZ�O�	3�Ϻq�pIa��f}B�nӼuoZ��?�L|2�'�ZW���]��!J���0|�x�bal�e���r��ډ��$��M��BN�"r'P�Oʓ|
�P*�Q6_�l��t�)fG<5����?����?9��|
/O�umڣ#̒��
�)0��^�
)J2��.|���I��M3�b��>Q�i�7M�Ŧ�Z@��/Ih���.u։�A4	��Y�ds�$�	)P@D�Y!f�-{h��'��d*a�e��T6�-�ش^�ꠉ��q�@��By�V�"~�u�O"�؀��(�,X59Y
�{̓C/��)�,�����&�`�E�>ʲ�z�)P��&-�A\�<�+O6̦͊��	S���q��e�,��0a���H��_2P���,7~ �sb�ʖ���[��)U�v�=ͧ���Od�0�e/�����p����?O�Oưn� Բb�P�Oerv��s��) &�ΉeoȀ��O�H�'eҸi��:�i柞()�ؼ_hf쐢!�8p�zA˦N��J	&<f��0��I�?ID��9Rj�'�@�+A�@�1�S�4<�PB��Ztyr�'��)�3?1G�i��xHQ�ɧ>(���/����e(���d���I��a�i>�	Цi8��
��� &�f�ƴ:`�i"�.@ƀ{�'RB�?=��x��4��� r�
S�ǣ-!Đ*p� �4�����O6��h�>mcn�k>ܔ�� ~�8p#U���C�'�g�'_��w���""�#b@U
����h��xѰ��O�6�j����j�'�?9u
2>|�����D� N��hC@�B�D�8Ǝp͓��t3TDA*�,$�K>!,O���O�@YC�-������$���E�O����O:��<�úi������'���'Y��"q ތV|*e9���Y���z��$�]}rDw�xxoZ��?��On��`�ԃ8�|p�n�:m��09O=��',��C�iT�0>��i�e��u>�Yv��9�r*�	9ʠ�U�g���������'o��'�b�s��9�᜗e�"��"[�,�JSޟ�9�4{V`�A���?Q��ih�O�
��HEi�b�.C�XJ�OZ�{�Ʀ*ش6��6@���r�8�'��R�j��q�.T��A�M�~,��k��ЬQ^�鷞|�^���I�����P����Pa�-H��$̓���(f�tp�d�DyRL}ӨD!E��O ���O����|���� �i5Q�[$� �O�Y�P��[��{�4 ��k�Ox����💥�C䎯^*���̍7(��8�T�C�T��Q��<��d�21>�}s��W!�䓱�d��y��j@.���T1���C�f���O8���O��4��˓1O�bP��y�I��BrT�����1E��[ &���yR�t����Q�O�Ym���M+�i/�ȹ��L��E�7O!9�=H7��@Wb-��'�b�ܫc����VL����?��Zcήdc',���%���Vj��r���<��?A��?Y���?����a�N䀍�vE�	x#V��/A:�yb�'[�!fӸ$؅��0:޴�?�*O�Q͑�J�d!Jd�G#��Q20hП��'��6�����#qV�I�(i�@�ɋ!��U� �W�:pv�ѷ�X� T���4��#dGD�	Vy�'"�'s2��
k�T��ITi�Hi�V�ª,���'���<�M3�*���?���?	.�<�X�J�:2&M��	�cǦ�R��� �O&�o��MC&�'��O,��T'V���Q��!?F��5��mH����� �VV� ��2��br(�C��)':yh��ǶQ>}A�_h���I֟����)�S`y�j����k͓{OؠS��Q�,��@��/=?�����O��nU�B��I��M۰*�[�b؁�M̝:^�i��CZ&:��F�v���&՗}��d�O0Ѫ��;"�hᣡ�<Y� 	F�8�+�Ǘ�" �2o��<q,O�d�O��d�O���ڛQ>�;��_'V�0#�`�X`�E
���M�6�R�?����?�O~��%̛�w�4Z�P�T�!��ppL��)j�k�i����>�'����6d�o��<!���>\����B��lC���<��K�r�� ہ�ж����D�O���	d�@Ј6A�
QEp,�����d���O$���O�ʓ.��b��y��'�+]�"��M� �S?�$8�̓-��O֠�':�7M��������i2�y�&D y��Y��&õ^��d�Oz��+G1<�I{��<���z��1f�W�?)e��M@*�-��	ӓ��?����?����?i����O	�E�;T�j�{��F	(c��O �oZ%~]��mO���4��H�K�r�8��C���:|��4O�MoZ$�Mնi���3"F��y��'��lz���h�ǌá��MJ'H��Ti�(:w����'h�i�lZ�8�Iݟl����w���X���q�!k�ٻ��My�`g� 	�Q?On�d�Of����=@�&E�V�

�f9�5.Ϡz��'<6m�������'�B��k&NBB���*��M	���5�Sp�ݭV��%�)OT�hE�X�l�R*��*��<iqCV����q����9��x�u��,�?���?���?�'��DL�;��v����JPt��F�ʑ6"�B@u��jݴ��'a@�s[�v.m�lXlS�F��[�F�ԡ$��o0��n� Qp��IU?yf��!pvʜ�m�<��'5�kl5_[&��`�_+|9�DF�7��D�O��d�O*���O��1�%S��4��nIF�Rl:���j�X�	ßT�ɫ�MK��^�d(p�Z��<Y�V�N`Q��� 7AC�TM�Y�@�ߴwX���O5���څ�y�'��P��͜�}��E�.~��);�㗦c������&-6�'���͟p��ܟ �	�Pz�зL09%�ݣ'�Ì.�e�IƟ$�'f6-Q�n�6���O��$�|�5"T2�ɱ6C�C��(Eɓd~���>)��i��6͌ß�$>���
_�a��$�O��̠d��R� m��k� �������*��� �ՓI>�РK�]��"�*FS���3F�?����?����?�|�-OF\l '/����H�;�8�C��C���z�nM���I��M�b��>G�i^�H�I��f"�����j~~���g�PmmZ�a�b���go�x���-��K�L���Q�'��)��`��Ȱ�-�|t#�'�����Iԟ��I�(��j��,@9wD��hb���p��c3-P)9�66�?0I��O��d9�9O0nz�j��@�1���]������K��M�v�i�x���>ͧ����!/�(%��<�3�F�0}(��u��"o��X��A��<a҇��9U�y�v	�����d�O����N��M����P�"��Cb�&aZ����Ov���O�˓uɛ6g�<�y��'�Rᙲ#��ڒ���+�H1�o�y�OJX�' r6-̦����䙙s�:Y)��A�J���Tn��I��O:T+EF�d�PmIa��<���-��b�e�9�?�'/4���Fڐ5	܁bDID��?9��?!���?y����Oj(B�T�l�0����G-~���Ҥ��O �m�Tt�����aش���y� �R�.�ab�	�=��3�d�y�{��l��MC3�_�r@)��?���@L|$KPdAi�? HB�jĖ$���&�ה�|K-���<Y��?)��?y��?Q��:tlu�AAص1r���ѩ��æ����HƟ`�Iߟ�$?e�ɾ8ͲRO 52��"�K1����O��lZ��M�0�'}�O����Os�Dz�`��$���[4���!��=K�Б	窅���$��نx��*U�p�O�ʓC�v�*�fX�7at�
%��M�~P ���?���?A��|2/O`!l�S� �	0:%$�цm� �B)�� Ŗ+E
�	��Mk��G�>Q�i86mXݦ�)p�#9I�@�⯑�:��*2��f�,����y�����"ג���-";���'��ԇ`���T��%�R䉐�&�9��{���Iay�X�"~B����@!�*�6I������w̓R��������覑&��Z����)
Y�q�,P���]�<�(O�7��̦��	Z�\� �l�P�ɮ�ƽ�t)��� [R�9&� R�.K�h@�qjOp����S����5d��	үִl�NPpc�.Ӫ�I\򉝣M;��C̓��)��hN�=)FCϮ>f1�5F5Z��I(���O�6Mz��&>U�ӛ.�ҽ��ʃd ��P@;^�J���ݜ��w�%?��'������g���������z�!�&E�Az.O�Ĺ<�|�'�D7m��m
 :�n�
ft�@ U�FKb���p�4�����'ÛvG�=:��D�2��!7�� P�M�[[F7-�O
�D@�?����O��	��@;��@����d
KR~D��˗0^�U���(���P�'d�>�$�פc?
���!���i��Mu��a̓��OY�7=�Vl��c٘]�6�CR�
)v\Kbl�Ɵ�m��<I)O�D�O�r�P#լ%I�'�P��W�H��4XIG%�f=y�'�p5�4��/�|�r`�|\����X��B�?p�@�gH�LJ�5��䟌��؟��	SyRi`�T$�u$�O���Oj��ů�r����I*(�� k��6�I����U٦�q�4&�B\���c�L���Z��E3'H8�R�q�|���u� �EfG�+�@��'��DA�7!�T Q�'h�e+�`�v�0��e�~wX'�'H2�'0��'.�>��	��7.Ȅ0�t���R�3X��I�M[&���?A��s?���4�j�6JS}/��6k��.x:�10O��lڤ�MK��i���`R_4�y"�'��亢L�+1�Y�N��TT�B' F�t��RI��C�'��	ş���̟�����`��4�X�Z6�q�숕\Q�Q�G��<	��i��R\�x�	}�Sߟh�g��&������e�̉�P0��$�¦��۴8�2����O �쟄�����-
F[��;])�H�@���|jt��'��KrL��H��ӱ�|R\��������eX��G�rXdD�'�۟��ן���՟��AyR������F�O�L�� W�x��%	䧘�i$0-�v��OְoZ{�X��I��M��i$6�[�L�� �)����88�Q�䎱xy
�'d�b
lM���!��I�?e\c�L�X�a��>U^�c'E��M��@��'2�'��'���'�\��6�\=�xY�/E-��	���O����O8Lm �N�����ڴ���(h��C�5,��R$˜�d�T��'����M;ûiQ$΄m�Z��'IR"\j��s� )$��L�	��q��j�TdC �|�Z��������I��X�T�L4tK@��5�S&�
�I#�ǟd�I|yRen�|I:'6O��$�O�ʧe��<��c>/� 
��?4��'�J�o���tӆ���i��?�iv��
��$��!{	zV�zӮ���	��zV��*O��i�/O�IIb�&�DK�3��	��(��X�EK��On���O,�d�O1���6���� Q<�8)�_�m�<x�H���1�Otl����'��c�O��lZ�!�t�bD�I���s����^N���4L���F��p�i��'5Т8f=2DO�^��	�(�$k#J)[�>523�17>�	ry��'z��'���'��W>I�Ǐ	`���D�,���ACɃ��M3���<���?AJ~ΓRe��wC��B��D��e� )�5#���3�{�|@l���?ٮO�	����6a�͛5=O,Ȩt�ʛA�D�)���	xj�ia7O��A��9����3��<���?1�L2B��6�T =������?��?�����A�Q��OyB�'e���5j0�B��ׄR�;���3%���u}2}�ܩmړ�?��O:Mӡ*^�W�Xe��Ɖy�p��4Ov�Z�Lf�H�n�;��˓��DN��g�r���5Q8��CAJ�Ĩ�[��r���?���?���h���dA�}�<+%�}�M��Tl+�$F��%c��"?���i9�O�ϠU�֭����>%��q�p犕<�dIǦ�c�4N_���D%��r�'�R�K�,��<1��P�p!^��'��qӼH"�c6E��|�S�,�	ҟd��ܟ<�I��H���=���S�b�)�v�0"�_wy�~��M�f3O����O֓��>"6�Z���H/���Sd:��ܗ'�&7�˜"6�|��?%�#p�fܪTٶ0Ot�U�<N�8E�qɍH�T�'�8e�ϺN(�9��|^��pg�ۺwG�"��ۧ����ݟ��I��L�	ß�iyRne�� �=Of%�$��J�����A��QE���52O>�m�q�"r���M���i�6-��{؜���D!"2@�c^'Eq $�� [����O<uR񅇬`�� ���<���y�k*a؎p��IA
.�C��

L���O���O4�D�O�� �S�|w���b	�� ��c��M�*���ퟐ����M��iO�|���;�F�|Ra�z	H���s#V� $�}����>�iS$6��B��`�?I��Op̣U� ���΅�E�򙂁�RV �Y�Y�Ta�H2���<����?a���?�aȋ�	wD�yV�T1y���z�^7�?�����$�ަa3�@c�������O���ڵl��!h�\�UL
�O`����Of��'��6���I��ħ����1����6��1�6���g�7d@��#r�B$�<�J(O��	Q��Pc1J,�dʌ_�����P|� ep��N��2���O����Op��)�<)��i}nt9�fي�J��؞X�|h#T�ƃ���E�I�?�G\�ش*͊��e	Zub�K���D�I(��i��6�^E���h�3O����!
�T9t�����˓��K�~�t��f�V�]�j	R����<�/Ot���O���O.�ľ<�'il2�{ph�	~f��B�Tk-p"g�ig�'Z��'���y� d��.�⢨��c-'f,&Ը	��mZ<�M�q�'��i>y�S�?-I�%�qF�	�g�D���B�V����'n��#�扆�xx�L�;{��E$��'��'d�����U�)p�O�qu�m���'�B�'��S�H:�4^j���?)��eLD����I�ʑ T��	=��2���>�a�i�l7�����'�e aժO��mؑ�Dbԁ�'_b��?
8�%��ݩF����?��6���u q�	�,�
��EF_�m�BT"���4���I�\����T��[�O&
�1^`�"=���F��A��(��� �!	?��'{�6��O�O�N�".$L�
�b�43elRʉ�5Q�������ܴG�&�Z�0�qY�';��)E��� `��6o�9T��@��a"��=���KE�|\��Iߟ��	�`�Iӟ��q ٵr�$�SGGN\v)H�KH~yr�l��p���O����O��?�,bY��	�7_&�uI`	���L��y�ߴ/H���Os���@S�͈�i�j�pi�n�0Y�04�`�-��	�e&:qq��h3|p&��'/S.��iN���v�T�2�0Q�'��'�����Z����4 �؉h�:��mā%jP�#f�J��h`���)�6�G}B�sӶ�o��M����.}$�I��K���Ƅ"V���G�<Y�ʦ����;y*�+Ov���3�&L)Ed@�K
>[$�ق���<Y��?����?A������x~���O�I|*�E�����?I�i�xm��OV2�b��D�<�A�D�2A�� R�?NIipF��5T����4-,���Oۜp�q���y��'hS��*4��W�#I��9���2���q�ٰq�'���ǟ��П��ɥl�v���[�H���1h��)�Iɟ��'�7M6>�N���O���|��+��wE^�rD�;Un	 ��x~R%�<Qòi308jG�'��O �'�:NTu0�`@~��P'��ra�i�5"؈X$J�{��'x��(����k���,t^�%��Y���37pаk���x���\1�?���?!��?�|�*O��mZ�,6�:�Ov:q �1S#<��Bo@������M3��ġ>�!�i�.%ȱ�
����y`�@�^�3��{�*Xm�z���"�s�8�	+$|X"B�(�n�'K]pӊݤX�ӷ�L#%YJ�'��Ο������	ğD��V���PD`��t�x�L�ۖ�Ϋ\�:7��Q��˓�?�N~R��#w޹� U�S}�L��f��U�):�F���MK��i���D�>�|Rg��i��4̓bxd\�t$F�y���j�^�j�>ΓYG��+Q떽D���M>!)O~��O���ኞ�V-���\�pp���%�O����O��D�<�F�iܔ5��''��'�,���b�/NR��v U�z�z#���L}�q���l��?��Ox�%��+h�����L�_z�b7O���Xm� ���<8��ʓ�bƁ	�d{�J,@��D� mI���#����@M�O`���O����Oh�}���W|��� �gy�-��e�\r����v!O���D�֦U�?ͻx��� fZ�<?�}r��E$)�t�XT�f)a�`(n���m�d��E�~}��Y�x��m�JO�hXg�R�@ $x�1Fj��]y��'&��'i��'����A�����M�Gʄ}�W�^#<��I��M�$������O��<����P˖�q��X>�S���[̜�'[��wӈy��Y�OU`�"DX�vȺ�!9�n�����(���[���Q$Mx��P���u�IKyR�D�!��*��F�[n �s	�/��'UR�'��O9�Ɍ�MC���<���˅ o�����*̔�P��<�&�i��O��'�@6����%��4o%��SPLʤ�R��Q`a즽�pkX+ Ǥ�̓�?1�nN�	��r̤��d�����1�n '�$3�N��QDݜ_����?����?���?����Of �,*2���˲f����']��'}�6��6��	3�M�K>�i�I���Є��!󨀈��[�m��[��+޴a-���O��x:I]��y�'�0�c�&f���Ç@�0r����KH�E���$�[7|��'����d����@�ɶ?�D��L�s}�X�Cd��I����ؖ'w�7M�co����O����|zv��e%U!�I�*r�R��{~��>QS�i��6ɟ��~r�d�'�R�����]�A�E���QM�wi��r)P͈.O�	D�\µx1C7�LJ��P���C"H���?YΘ���Op���O���I�<q%�i����dN�C#���'�9=@�X��-���Ŧ��	G�ɝ���W��A�P�}����?\���X�	^��l��M��)Η��]��?)t���4��$ .��dA�
�<����/NH\չ2eE1&Y��<y��?)��?��?)+�lPiuh�
�����	��e@�
�Ӧ�Ybd�,�	����h��'{6=��]��&�D�SVؠi��E��II��ٴ]�X��S�?}�ӦZ��Tf�� ���d&�W��HY��ԙl�����6O�0y���oD�Y� ���<	���?��Ίf��Lh&Ė+>B��ek؀�?���?����U��3�k����؟ Y�A�6��}k4�J>E����MS�N��I��M���i���>!�
��0[�*�N��L��KG�<A�x�"ypPNV�Y�Hs.O��)�1BHn��!��O��ւ�Z���ҷcT� 0�|�)�O��D�O�D�O£}:��V�5zኄ(�h�NZ�o]$,*��(
��@*~��'v6-+�i�5�r��1�VЀph�3u���!o��Cٴ/[�F�l�*��C��k���O֙���1*,h�b�R3r|�D��
	�8tܑ7��S��Ovʓ�?����?����?��� ;�	�`��K�K����H�2��Qy�x�L��f4O����O"���@9Y�J��pd�
���:��5:���'KT7M��!��ħ�j��BH"y"P�T`�!ac!}��pj&Hן�*y�+O��'+ (F**;�#��<W���3��#E@�8�����V�?���?���?ͧ��$MᦱHV.f�ĻBL�SKЈꄈT`�=��d��P�4��'�N�t���b`��Qn*0�v�!�@�*���K��|´I#���t���D ����C�Xy�O����%z� �L[/� ��.ɗIH��ȟL��˟���ן4�	~�'���P�B�Nϒl�A�U�q��P��?�� ��6�����1$�`�q�ܘ5��$�ͷE���aC^0�?I�O��nڨ�M���aw ���I��<A��z5N$�B�F�T�$��i��k"�����Kv�j�
T������O����Oh��Ӿ2�&�e	Y8��A4��Y���O"�c��vo���D�O�˧B�B�xU�%J��Sv�*5P�Y�'Oj�ef�V�v�l���m���?	Ѓ-1\oVy:���?�:��F�=xn��ꑣ� �'W���&m�J`�Ԟ|���mb��*�)'+�Fa�iU�L?b�'���'����^�8��4rG(H�w�J�`�AA���9X^E�vĈu~��f�B�۩O��m�0Z#L�����h�4�s-ۦk;�ܴ��6��3�\��'ceV�u;�А`O�l��+1V�Lr�01�P���Ζ<{��dy�'��'�R�'��W>Ⱘ�Izdl�u@S� �P�۵J
,�M2	��<����?����9O\�nz�])A�|?ЕH���G�5�eƽ�M#�i<T���>�'���'<�Lۢ#
�<Y�gX-��:B�ǊY�*�	��^�<9�"M�E����������d�OZ�D�6���a�m־^j&t�2lB�9Jx�$�O*���O`ʓu��M�;�yR�'02�R&'�~�x��O40���'n9 ��?9]�tHشI���O����+��9ԗdҊ����P�<Y�0 �i��^+PmhI{*On�)�`�H�1$��O���D$X���7g� �`��F+�O����O����O��}�;IU�9�ׂ,Gd������~0v����g7��8��$	֦9�?�;""��d� J�ɊU#��Gx�4͓j}�����lZ6�^p��e���I!9�	�����خ'�zy��aQ/{I�%�Oʟm��'H������͟4�I����	�b�f� �K(Y��k�f?�|�'�P7��w���O��4�9O�1yA-�D\������^��<Q��DP}Byӈ(m��?9J|r�'�@-�Wz�ܢ��0#��,�n�b�!IY|�`�,O�p��hP�? l�y��>�$�<ad�A?3%re�wϕX~4�*F���?Q��?���?�'���٦!����%!�2�
M��
uh�5�Lޟ|@�4��'�����H~���nچ[��ff�Rk�(�W��2t>�L�� ��kf��I��B��3@FZ �n�Ty��Ol�X�XL2�#�f_d��i/,�f�	����I�p�	矀�IM�'~}t-Q��W;e���և��!����?��tg��(2����'�7=�$hz��p��V<���ŀ� ɖ��Il}�AlӴ�n�|R�GG;�&�	埐�Cc�hiu��o5IZ���� C`=37�[6yV�&�4�'���'n��'�x�A�߼&�d)�㖥lQ��7�'$�^��AߴmB8�0���?������e)�R%f��ձ�+�"����$F�q��4X�����O'��L�j�Ȑ�g�V�����ݙ+^����oK�>�I�?-zSԾ/2��%����:7fU�U� c�Z�s���韌�I͟,���b>��'��6M���4�ҡ
v�Q�j;"9��6n�Ox��Kݦ��?9�W��(۴a@N����ͷ(����U���r/�����i!�6-�F]+�9O�䂖E�%PCW4q2�-�a�dG\&m�7k�k���̓���O��d�Oz�$�O����|��#J�(�H@/�W;n ��Z�r$�%�"K��'��O�S�l���K��q��a�#T�����ϔ�|(J�iT�6�H՟xק���OT��	G�7��(�'�������/aR��Y���h�c�'�liGh�_��u�a�|RX�\���t�t�]9	K��2��U
p�(A�֟����4��Yyra��X�:O����O��c�^+`$`#gG��xS��O�O^M�'U67����X�����6��SM�#k� �J��H���O�p9WK�8���5@�<��'J����/Ҁ�?���ɧB�)�w�Q�}CB1��>�?a���?����?���9�Hh@Q��,M�j�y ��#�|�ٵ�OĤn�9]�����'ɧy燇.�䁹�@��=����L��y��x�$1l���M���/><���?��� ₼у��qfn��@&ϼ�����%h�m@L>�-O���O��d�O���O(�z"=c��̸�jRֆAR� �<ْ�i�����'�R�'k��y���\��uR��Q�z���ֻ	��v!�aq����	x�O�~�Z� �|�D�T�c��8�HZ�d��Q�C�AV�˓����aGH�]<�+M>�)O>�8$eN'i���F*�*0�(��C�Ox���O����O�I�<��i�H� �'����B�>!x�Q����n;���'�n7m.��	���Φm�ڴ|�`Z#�$�eA=M\����]	c�H��һ��d�B���Յ��n���D�1)��Q� BX�/����)*P͓�?���?Y���?a���O]��*ツL^T�Bb�Y�r�P��'6"�'l�7�I*t��I��MK>�R�V�89��<������D�"f�S�`�޴YO��O��D����$N��d���,P$j��#
����ɏ�F���	�䓿���O��O��$F.=.�Y�6E�%�ʇ�Bv��$�O��[*��
�yR�'�RX>y( 
5-˜�P�Ο�az����,?�wR�x
�4_3��,�OJb?�`���5 ���/IDOt=XB � &z�Ecv�)k�̽�����]<H���3G�|��X.�	�OT��1��:"�'���'r��$Q��Q�4)����
G�(H�a�'b��)S7A�o~R�cӀ����O��l�!f^��1(� ?����l�0ؾ���49���� Dl,��O��qƉ�SVN��7I�<	��L��ͼH�~���F��<�(O ���O��D�O�D�O�ʧy�4��'�$oV�H�wn�*Q*��i*�����'�B�'��O�r q���	cg�(���B�[U$�P���8���m��M� �'#�)�&hg�y!�e��HU�\@����4v�$��)���d�<���1BK3^���O�˓�?)���4��tKźy�4��"n:Z����?����?�/Oĵn��CHf�I��h�	�Z�,�c_`rH����MP�?yBP�l:شH�����O�Kb����-Pq؝�ń@-fh�'��0I �Ѭ,�V�ӟ��U!�^̨c�'�L!kt_)�� s�!�>0�\���'2��'Z��'��>U�	"G/$H @Ƨv���E��9���9�M�рD\~2ep���杣w�j��L�Q}���hG�����3�M�R�i��6�M`w��󦙟t����T(ZǮƱ\�6|I��H�Č`�M��;\а&���'�r�'C��'R�'fPa��[L� �"��_"~��RR��y�4Uh��Γ�?Q����<i��҂�p�(��`�f�bG�Z;"����M�i�.�$�'@$ �X�k�`�4b�0Jlq��I�z8��-Ov(� k�.Z*�� ��:�D�<�����?�xyP6놡k} �jse��?���?����?ͧ���٦���c�����9M0��{b��VB��#b����4��'�4�O���-i�l�o�!c������*�@�F;�Mk�# p�@�`:^ASb�Q"u�=N~2D�ƈ�x6jӖQxD�f#��0{dh��?O4���O����O
���O��?�����s�	7�#bz�"æ�0������4d|��'�7M7�$ǔ:j��Sf��8<%dy��b	�L@@�I}"}��lz>Q��GI>px�
S��¡�&�X���D���2��M>v�x0 �����$�Oj���OH��7s�X�2���N�\Ÿ�퟇��$�Ofʓd���	Y�r�'��_>��^�*41*l�����<?��^�б�4�6��O����	W�nrœ�H��{�8]j�$߇y�ve���F�t ����<���̎R��u�L>��GJ�7��Ź0lB
��1g.���?)��?���?�|B)OL�m�=�v-p�I˴��T�7*ܒba�	ѳ�WH����MC���>�i2�ls��� �h9�I/��EB��`� Tl�4cЖ1s�kr�����
�|�A^9$:x�'����M��9cX��e�';�I̟���՟�I�0�	W�T�Qc���@�D��Y����@`64s.7MX�����O��(��7�Mϻ�pű'gIi�Ƥ���Ɔ��l��i�r6Z�,է���O��d ��x���'�������C�`UP�ML'r� H��'v�JU�З��h g�|rU������,
���V����e�[<���8����\�Iݟ���^y�v�Ѣ���O��d�Of�n�b�Ѣ��uKs�1�I
��d�¦�H�4F�]���a�u-�|xF��~tm��%l�|���g d���,8ޜ5�'3����=Y��dqf�'�N�y�'$C�f$��)T�Q�ftV�'0b�'���'��>��Ij,}��'�2O�v���Өj/��	��M����?�{ٛ��4�Za��(=J�@�"Y/c�U��4O`5mZ9�M[ƻi�&�� O����/dLf��!^�T `���'r0K�@�"f��"(��<���?����?a���?qS�ޥ)����(�	�Vu�d�����Mʕ&�����֟d$?��	&RU��cjΗ`�5��"uK@I�O>(nZ��MC��'��>�x#,@9;���9���%L��i�3Ώ{f�����Dyr�υ/�B�0��3+x�'���E���j��[�p�<�$�t�����T��� �i>�'�7Q:(���D.X,���F�r���I��^��$T����?�^�lK�4@@��Cw��K��/'1���LB;�(yA���a���r♟��蝲a��m��'�k��5V#þ/>�8��`"�q��FP��y��'F��'H��'��	q����CU�#��H0��L2I��OL��¦�*c�)?�þiA�'�8��[7B���e�	���	eO�O��~-��B|�L�I�Yo\��;O�DXwQ�P �kŌ3rT�p��E�b�VF�K�^ܨ"'(��<���?����?V���!���\%X(ܕ!F�ŝ�?�����D�צ}+gm�_y��'���R
L�YG���l���2%K�H���4��I&�M�ij���:�	�� �����,
���,A
V��gD�.B���'���*b�ʓ�r %�x���AH>Yv�Y�U�Y�����8��.��?����?1���?�|+O�5lZ�wVfiP���-E��P��Y�C]�DzG�Ɵ��	��M�rB�>�F�iN�E�g�:��u�^�D�u�p�j(m��\��keab�8��%޶��v�V�U�x5�'����#!ʃ_�(�`���UFFљ'����D�I���I����IV����d��<� ]-�)u�\0;*7���Fx�ʓ�?QH~b�����7(�R�*tb:A���0y#�x��4Λ&��O,��|��'���#{�F �1�ۣ��U*��p���Si&��+Z�4��A�5�hhN>�+O���O��j��w7��Z�㊥z*�7�Ob���O��<9`�i�V%�1�'���']�@`�
ƥFlX��L�o��
��'��'���t{�ƤoӞ���W}���� 궴C�a�(2��qd��y��'}��qp��:tZ$:4X�@�S�\@�I����L����P��g�C%.����eP��I֟��	���G�d�'7���r�d����As��'�6[�	|�	��M���w�p���
�&k���AD�0s�4 C�'�6m�����ߴb3��x�+�<	�h��.�=�����\#4�$�is�QՆ8���M�N[�O�ʓ�?����?9��?Q�]І`PE��<PCb<s"i��w
B��,O,em��IY<�I矘�Ii�s���h�J{nň+%^<@TڂO��$���P�4FX��SR�0eHӬk�Α�%W5D"p��P�jd�'�	��hH�!�|�X�����PA,�jt�_�P���u'����	�L�	Ɵ�SuyRjw���*Q>O,`aAc]a������RW7O�4��'���X��jq�lmZ%4�4s����|0KY5a�dIp�g�=	^�[���|��h
$��S��e�%�5��V�W\�5��R�VGȱ7���y��'�R�'���'{���י>j2�3�$�H��UAB���]c���O����ӦQ���,?`�i��'�\�EGˁ`p��1�e��nN���E��O��~u��m��)]	=�6`㓜���s��A���1���lq6���]�	�	K�!��%��'~R�'���'mxQA�W�w�YA�Ib�8T���'O2Z�3�4*�0��?A����:
 ����I5��Sh�x\�ɪ��d�Ц�޴! ��)�J�*Ibg�!z�@P` @��ȍ��H!�h�S��<ͧEwpЙ�eH���=�r4�3�5cg�q�C�CS�2I����?i��?!�S�'��	���Q���o�$C`��l�X���֛5�8�J՛���	v}�k��- &��`y���4%�.i�>��r�KϦQ��4O����KZC~���+�"�2��8Qu�yA �2vhɸ1W�h#�$d6�I�������ƟT�����IY�$�^�Q�H1J�7�pP�ȓ���7-Z�=-��O
�3�)�O�4�� j�(��-i�m*�ǉ'K�g���ٴ|��iP�O��t�O��#���~��n�I� �n8�x�c.��<9ᆙ#+D��#�����$�O��dH+cp����;���k
M�8�����O����O�ʓ��v�-z]��'iRlZ"wjiQ��W�m����
���O���'7�7�M�������$��mh�5h1�
��}�@��U��I*���!t��/], %?ْ�C�-_� ���0A�l����L A}|Q9�OB	\�����՟���ݟ,�Ix�O�B	�!�J���F��X.��Y�i���g���w0O����O��O�9�Ĥ�Tf�;�8 �l�;@�Hࡁ�O�nZ3�Mվi�H�"!b�&�y�'�ځ�WL��'fZ�*s��$L�5�n�u �H�.U#��'�I����I�����d��>(ƽ��iɸ�k~� ��HnyRmm�h�CG0Ot�d�O֓��d(b�Fq1 k���mM$Iȴ�	���>g�iN�6-Z���F�4Ww�TڃƓ.UEj�ʗ�Ʒ-z���VF�)j�	5�Ժ�eP?���%�ܖ'֖��b��R"�U���:0������'��'�����_�p;�4@zɡ�]�p�-��2�	Q΍O�>����X՛V�Dv}�uӼoZ��Mc�jY�i!�AS�q��Qy���?3rĉ4b�u~"��.�>�r��<�OMR��sҤm�p qS xrѤ�~�M���?A��?���?����O��������I��
�/E���Ӯ�$�O4�mZ�w�������g��7�*HC�d�_�&9�TlJ�_
�+��M�����$qӐ��4��:�3O��D��1;��7�>3Y��c�B�]RTċ�h	`F�,��'��	��I��ɷk�P��	�%�$�!	�u�
���l�'��7�ٵ^q�D�O��ĵ|��$M�_�8�!Q7_�dd�4n�U~��>���i�
6��ןx�~�u"�O�RYk�FX3T��P�%�K'���č4?l��.O�)<���&&5�d�*[�2�5Ò�w<1k��O+p>n���Od�D�O���	�<)�iYZ�C �XH¡�D�[*1ʑ�U+�y��'�2�|�O��I�M{��\d��8
2MI!G,�]���G�*\�Fl|ӈL[�o��l���o���y|�)B���G}�@��<��a�d�T�N�����t���<1���?���?���?a*��E�aE�*t���2�ʽ�2���(��	X�??����OB�7=�`H��?���H2�"=G�%����Hڴw<�X�b>e��M�%�L�I0��" i3JJ���:&�� 0� ���W�)h�&��'���'�4Yb�21�ӥ��x�d�'���'�^����4S�"�Γ�?��l���l��lP�l�T �ԡ�"��>���i��6m�<ԧ� ������6^��F�Ue��� ��hK�G��jԨ|X�	J�{�lx%��П8Je
�H�:L�%�#A��ira������(��͟ G���'W��E��!%��;vcD�n�	��'i�7��8U��	��Mc��wFF<@@O�iGfIۖ�hy��J�'T86�\��x�4��r��i~��7��,�$�D�J��bf�n�	���e���b��|V�d�Iʟ|��˟t�����ch(�r��b*�3o�2�s��Pxy��h��x��9O����O꒟��=p(q��E>H}j5cs�_�Xt���'��7��������H�\497�J��x�Sǁ4/x:M[e�,!ݺ$1e�<�5m��� �҄R������<*���"v�Ŵou"%���S U����O����O��4�hʓtS�&�T��A/ld�e $�!n]��Pp�\�<y��i��O���'|�6MU�	��4O9��1�2c�ѱ�G�;�L�@��@��Ȝ�'ZV�0%�8nYAƚ��ig�1h��CS69���;bzJ�9��b��������I͟�I[y����>(��E�2`Y�*Q�=�B���y��'b&�򩣐��`3޴��?��AIG�,	'I�g� ��8��'��	�M�d���b?nYJ ��O���D�I���-L���x8'� �m)5K� ��O�˓�?!���?��47j�S)ۧp�8��=P(�"���?I-O(mgj�	럴��L��E��P�4������_=|P�w�G,���XV}rfa��Qmڻ�?ي�䎐}~, ��ô�>��W>�Y�L�2�õ[���\� �0t�Is!g��>�p╩�@Y�����T�I����)�Sfyr@d��1�Ք � �0\`���Pj^�$�O<oA�l��I��M� -�2f��XH��M�n���0�/�)����sӬ��ҧ/���8O�r��aV�L�V��'�2E��"?ph�	G�2 �鳚'-�Iɟ��I���I̟��IX�E\MR�QF��o[��`�G5f�7M��P����?�J~���V1��w��d��ؘ8��ݙn��xҪ<�U�a�b8n8�?�O1�x�h �ӕG�J9xݾ��횲%XM�4�ݷ+��D�i����%��O ʓ�?���t�$��/ߜ~�ܴ�"螛v�$�����?���?I-OJ�oڧ}������\��-g�TqsG��?d��Q��އ`@��?!R�p*�44�&g�OB�"�޹ E$Ӱ>$��DwR�'P�I�ĤD��X���dFB6n��ZE�'XV�`�mE�<�]J�Yh�c�'�B�'/B�'M�>q�ɻ)�
�	��\�3���(bA�' ~���ɒ�M�f��y~B�kӀ��] e�v�x�%Y��
d����cZ�扡�M+�i�(7m�*g� �D������܈sl<p&jGu�q�jN�^��g���y)�h$��'B�'�'�2�'�:����9m2z�����D���S�Z�8ٴh',5Γ�?)�����<��E�O��{6���<�Ud��#VW�ɛ�M�6�i����*�'=(�1!p�E8�La@��9%�:���^�(A:��(O�4����aX�y�..���<)0Ʉ�a�6��d.�3e��CX�?��?9���?�'��$�ߦm�)g�,[��2��Y��
�>�T^f�C˦u�?9R�P�ٴ��&m�f0��A5�T%��+|�Z��S���PC��T�,�?V�1(�ep��5��ߗ�4�@���'�������y��'V��'���'�b�Iæ6'v8�G�W� MH���U��D�O���W¦A��/<?	�i��'�N�c�J�,j<ʥ,�'��eQ׌�O��5ߛA{��ɚ�0Mrp0d���;��7N"'��eTTi���H�9���c��X1s���$��'=��'W��'��$P5� ����nO����e�'r_�P��4kv��Γ�?����)�?W�Z��0Iܨ��  앑��I���ܦ%@�4Z���)[P
 -�'BT�/���er��@ǈ,V�}js��<�'z����ˍ��ά��P�M'g�⁘#�O'��B��?�/O���<	@�igp�  N� ����5��1�w����Mئ	�?��V��sܴDj��w���+b �/:���å\���r����R�N���5Jthhb�W�U����'����FB�_�h�bƊP�+�Xd)�'l(��ɅF���Y�xZ-K���c��C䉂M���'e]&j,� �_u��mHLR�zF 0�#�7��1��݋^�\K�gI�#��Xi����N׼ Q�iz5��������|�|j�C��]������84+��Ϊ,	��:������8#r�D��*RA��x��\�uf��6,8�N�%���zĬ,Z�P7��O����O ���j�poL��N^�Nd�s�Y�N��|a��i�DX@�'q��'��O�����IW���fɰX4J4�TA�A��	ܴ�?��?�ZH��O��$��ps&�ڄr:2���K	 /~h�6M�Oj�$�O�j��X���'�2�'J2�Db�I�./�
TH�C�XZ$��ٴ�?��a��v*�Oh��?����� E!:`p q�у{��Y2��iZR��4=��'�B�'e2�'�B�'T���c���W��$�I�l �$ [�;n�c����_�柈�ɳ4�A�`Ϛk�r�b  ˥.ʼs��Wҟ��	��Ԫ2e#���<���:r�\BvH������s�"Ol�Is��z�آOOy]���D��ɼ/E�]�k�־���tiJ�[�"W���IC[9h��C 1�i sm!B�u0c��D ,@���������FVj���GE/-����j;vuL�qЫ����3���N��,���?o��I�1 ��3�&MJd/�:��<b��#N\�0�ݻ{�*���ϺP�
� %AU:M�ƵZ�h32M�yE��O��D�?���"� ��W�֘x����}J^w�J-�_>��£	&Y�¡�+�N��B�.}2g��d%dS��z��H��t\�N�W���s?�<8���q��2�a�	� �'�|[��?ѐ�i�	��%6|A�4�²H���'5��D�<����?�|�<��I1O���r!/
E	��@���q�h��4R��ƚ|���G�ܩȅE��B'}R�7m�O��D�Oq��
ޠ	�����O��D�O�X�n��GؖA-|i���.��)K��X�l��=n�K�%q̧�M�F��<Yp��!X�n難n�A4�p�!����҉�6�֤����B$��p��4�iPL�'"�d b_L>�H�_7�D����-�d_6���L>Q��Rkcp`���֮Z6�d���{�<	� V�P^z5 E�.]bBL��E��<9��/+����n�ɚt�~%�B��+�<X� M+9i`��kۚ+I���ɟ��I��\Yw���'��i�[����tG��j��x'�T<���S�i�0�s�A�'�x��	���Q��J�jv�
�ko�4��G%h����Ug��z޲l���$j� �e!-S@<��!��^e��A��O�Ն�I�A@6�d�5vya�����B��
H��`z#)֊ڨ *f �Ehfb���ٴ�hO�S6��RD(ۨ������<k
C䉒y)�1A�Q�%p���ׁ�^��B�	anҰU�f�B��C�5<ÀC�I�M�\����D~�f\r��ƑG��B�"/f2d�v��X��o�"%��B�I��.���@�9�@����ô#+FC䉛TM�u21LV0+}&�pv�
4�jC�ɚ1�̠��4ML�����? lC�	����`1`���Bܳ%HLs'FC�ɂ2�}�B��<m� �J�FC�	#t�ѫ�	���������B䉫9nF��@X2��	Jf��"w�B�Ɇ)�*�h٠Q�.r�B�	#$.���-'uؖ�1��`�VC�ɝ�FQB��_�_���;��	6C�ɜ-S^�ːȔ)s~ A���Gj^B��$��3�,� d ����C#\�B�I&%D�<`CJ�)K�z��	U��|B䉼=�B� ���q��%�G�19�^B�IR�V|�E
Ñ��l�g�={�B�	�_���c�eE6��d�qS���C�I�|MH& �U*nH!�l.�xC�I�#�@Z�
҅U`� ����pRC�I�=n1"f���2`�uf\9:C�e����ˮ��0YVL��l�6C�I�*���ӧ��>O�D��Nܮ�VB�*F���0l�b��e�
�>B�	/I.� �T쌄ې2�EX�Pn8B�6'�Xa¤F�����Y%KB��C��}�Ty�e٭
�N���m-E-�C�ə.ڔ�B�D�Xmä��!`��C�ɺO4i1�N�>KC ��D��~��C�I8UG:�� ��CV>ЩSB�B䉖I��գ��-.�DΎ4�B�	�7�h�D�Ka�i�OB|�B�BN����M�6TF�t��4[�,�"�,��II��hGm= '8M��ˊ8"�2�' �p�b3�kcst�Y���'x�9����#�!�S��Ve����@����"�%ĸt�#n]�IH����5�� ��-@�/&���$H��%��f��i�nδ7�h'�ۘ�a{�ΐ�@m�}��K1M�l��Y����M�,Ff�d��n Y��)�y���dl���l�	�59����}�&N�5�P���D]+%7f���o���'�`�Y�bZ�x�֩@aKO35mݛ���Uh&��ݴj�
`;�ʈ ����K�[�����C+����ЎOa{R��Gn���ҫ��t��u�׸cu��s�ڿk=���A�.<���8T��('��}8��[����Fl����uNb%!@�TM�<�R�_i�pQ�
(l��S��/M�]���Y����z��ӏtr�*b/v�3�"X�Fᛚ#$�z�h� z@���;�!*��8���K��9#�f0XT�
?�� كL�di@�0�`�%U,a����}H�x
� �(#p�^=S=���ەlUx-F��!T�)!t�N>}�<���å��,@A�O*9r��e�*��g�^x5�m2����Pxb��%���D��3K���2a ��M���в�1xb!�?�e�D�H�+؎�S�s��۶��i�P�h��>5+ %��G-D�DC�!^7:Y�xX%L���*�Od�bt����W}b'G(��S�j�V��d���m{��-5���E��/jX]C�o�X\A�ߖ}k��YA��{!���!m\0d�*�󴎉�uD��N�
|�A��Y8�i�#"'B�"�REgf��C/�`�c@�T�$�A����<��
���T��&hԯj��ĉ�d��@+TA%�d8DH9�����.c 4�B���;Ѡ�x�t�-��v��!��:�':v��/�\�F�K�j��V׾l�ȓZ����&'F�h)`�
7��#�n�bp``@��B6�qsG�@Q�3�	�G���S�H<o���:c㛆r�B�	�r����ٛd���ʢI��?���6JI9./��J�`�l����I*��Q���,�z��Y�&��D�;۰�uB <�d�P�'�20Z��>ft����B \�{�'�`P�?j�����	F��b�}�L�1j'Xu��IP�O�����E�h��x�Sҧ5C��(�'��h�#�� #6=�B�<@i1rc�&o�r�6�>�f�>I����.���5�N���]�d�U�<�� � �BW�8W��S 'H����쓒h�`��'H��&�:2�`Ԑ��\wR���ۓZr����F��>4�d)����H	F�4d�0��-!��ؑ���h�cT�R�@(����h�O�|;C&��#�RU؎�)F4���'�ь4�w�ק�!��,RQiSŊ%e�>t�#�v���2�*�vլ�'l�"}�'�F��Oѯ����Nè��y�'��ܲQnL�]�����#_���۴�ʌK�ΞrQt��$�!�q ���=N<Q��)ʉlea{�ʙ*�0D;��\���q���?OZ���5Y�����(D���"I�	b�ӇCz�ƈ@�l3�I�q�(���d��>}��л50�*@�vZ���q�-D��k��.hn�(!M�H���$�ۙ6����n�i�D�W������&���T�A��z�hr��)a�!򄙭����F� !G/��R�ī&���+ǗRT�"��r��ԛ3��Usn���X5�|q�%4lO���	�N������*Rd�I�Qp�Z��AK�u���G����	�8|lA��W�4s�H�>��#ݼf�4�2ڧK�d	��ߧ��] ��	.*�T\�ȓ4�\L���/?�`�S�Io�DH��Մoюq�N�����Y� *Ėv`b�/E���z�(0D��27�� ����E��W�Dd�L�O�f�_$8����4]�N�K���%���c���
NVa{
7<yQ��՟�pd��^!"�,ћE�u��$D������2���iC5R��-xS�"��3���$/ B��>%YW㏈���Ո[�u�f�+D�h���?��ڀ	��r�-��M�J���C���M��T���D�(vX 4��J�0�z�+Ϲ
!���-4�H��sE<CZ���'��,>���.
)p����c@[\������G�oWf�sC!��^@,u�U�5lO(%����?�����Hw�@�V���a�ʦH�*P8Ʉȓ�꽱��׆ϴ�U�̔eg��>97m�9F�.����*ڧ+D�BC�Xe�5j�P�zc���4���؅@��[z���#E	)$�yC�C�����I�<��Y��2�^)S��i�'L�K�P8	Ǌ)D�� 4E�83����3�ٵb�z��fӦ�cn�t��9�
�{b�(����+1�NQYu���~w~���	j+NP����/v�a���Q���O#t���ԅ�y�d��`ܨ����.��L�4)���'&��٢OA?��a*A�w{J�AT��"������<D���T�t�~D�4 �:Y����eK:�Z�CS�Wd��v����E-;�$IBq�ؼuf�5��f���!���"���Yd,O�f�Eb�E�:DÛ��x�����A��D�B�	�:g�ME`Ǟ(tV/@�a{Bh׾h�VB �D�)� B|"$�Dl���7בHb`P�"O�8��
�l�(�r!A����p6��V~\�̘樗��h��p����e�i@�.	|���1g"O�4i�΅�n\�*�FJ�~�ˠ^�&l\���%}�I3�g}bƽ;�t��ȓ�}m�|H���ybK�^ְj�hZk�D�q�ۃ�M����:mL�f%"|O @�"ĵ2t|�{��+	[ R��'o��z!i�"*~@�ɷW6k�˶tCg�W0B�ISŬ	�Y�4���J�o"�����䋨m&���f���h� -;qa��(�"t[���K�X`"O�����=,�l����;�X����Z�ڌ�Q�j>}9�g}�eO=^,�i��N����1х�y���Vw\1{��V]8����#�M#��&�X��Ǣ;|O���*9<J�y����	�(�#�'OP�q7�!e�D���#��M�cB�05|k��wQ8B�I�]3>%H�J4	}2(R�,�K{.b�8���¾K!v����Y�ɐ�/�*�"AO;�C�o��9+D��(��`�wN��~��������1�O`�G��O�d�3�i��D0�c�n=n��W"O���R�
�
������28*�R��ug_�	�p�[Q�'�S&��%�p1A�ǲ�P� �n��Zr�

X���$J�) �1�L-��ȣGE��!�K�ɨ�R2 b���'�UO�O��K�I�3|�4-����+���e��Q��
�C�>O@!�ʳTI.ik6KZfpB�r�A�2��=I�삖&3�Db_�(Z��Y���o��9����O�U2�k5%#D�8��</t༊ H:����Ob�@y���q K�)�8��<�fe�7/�*$9$b�-5�.(��%�v؞���.�%%�e���(/��u��=�8$ہ�/V;�x��bOw(<��AL�7ifH�IY&{�x��1��Z�'bM��.�'qeޥ�%I���O��`��F�+F��O��J�ځ9�'�<��$[p@��C�U�AE�廖�ؓ_̲�T)~�Zt�I��H��I�:R���v t��Gǁ�|w]��"O�\��m|ɔ�ZU�ӥ"��@�ߥK_�`ÓDY�e>\(f%4AH�?iġ^n��CDC�K�-Q�D�b؞hjva�eʖ	QЀS=N���5/�v��@�#7F�h�ĝsR��䑛K��a*@j�'t6�E�N�"ḇOb������><股�u��"���۵T@,z�hN�&��sƨE4�y2��[�(�V4�(0H��l�(0����3+Q`D!U��t?P�Ȋ�Y�h��'P)h̚q6��(rƔ�$D�XA��ީCی�HH��Zc`�HS�5t��8�ř�$	�1Ʃt�~�=�?k�8Tn̝}�r0ړ�$V�v��I.�R�@�ʬ���s���k�Pň�� E�x	TcG7C��a��%�O��a��>K�8����X���$�$"��,��'��-�hR���']��1 �G����4X,z"|�ȓ:�Б��
!nߪ-�%LƩC ���d=9����ʂBd��Ij��~��S�D���@<�d40dg�9�y"A�(^g��Q�ެt��DZw- �yrN�Y���H# Y�5W b�~f�P��Ɖ�z.�T��� |���k�h��4�ք��1���g�xՅʓB|N]�-�&�^��ĺhpC�	�9���3*Ơ8F�Y��B�t�4C�	O]L�Ȱ�<x�B  3,C�I�*�0��%��L��]�#��B�?%)��BOH
vF	sjV�AJ�B�I�$z����?����� ÄC�I'F\`�GE�|%���d��o0LC�ɜ!y��S��З;�~��B�Q��B�I�5�~���ƪE�*��VA#&�B�<X���c�<y�d`�w��t �B�ɿ��Q���K>umJ@#nS&@�&B�	�},��w���O>��2A��0**C�i\�E�D(q�L�&G�g�
�ȓ+��``ΪKFn��+X�Fu���S�? �D�Z�]���m3���"O~���$L�'�a���;S ��'��<Q�ְ{�,�'�[�
� �A�'^4)��(AB�P�07l�����	�'��S�(��S�* �q"��T!	�'e��A���.YVHL�P�p�H	�'�5I��7w��o�l�h���'bj�[$����"��2��\m���'�䰇d�����jH�OG����'�7��M���d*�5�ت�'�:��n��
���,b֨�
�'��}0�^?S]fq#F�H�,X
�'��be&��f~�93���]���
�'$��rf�;[M�qC�S-[xZ�I
�'
���d9��M"`�Z��ty�	�'lԙCgA���U0W.F)}͛�'��|�-��"JJQa.w2��	�'��y��\�}��z�(�c�q�	�'�����-T�'�j]�P�V�V�V��	�'��j$�zפm�4�QU¾U�	�'p2�0�ቛ��"��P;�HP�'�Pu)G� ��ݓ��z�lx�'1���S�^.m�ı���Q =r�'�t�3�%t3�e;���z)%A�'�@��k���F����y���[
�'�� 
���q��@Q�f�d!�
�'�^Lr��<��D��l�]E�L1�'���b�"3�z��5�ǆ*��S�'i������;&y9��Fh�E�'���%
ִ��u���Ǉ]�"i;�'�b�ö�_&exR�J�%X.�;	�':�s�l�	�]�*�K����'���	Q0Q>9��gE2���#�'*	yƂH.��ܩ-�% ^�I	�'�Թ{��7y�-��g��V��'�VɹaܓJ�"��VF&�ܩ�'��m�K����0��O�b	�'��Ip��$ | �c��~�8dX�'���@ÒXL����t�n�9�'�x1�,Q�mx\$�dܲlu�9��'LPMRL��0�"�Â��h�0U
�'�z���L�Q�0�:�)�
͊��	�'�vu�G��/�>H��[
OTX�	�'������	8����g���(�	�'�^)�.ܧ�������/h��,�ʓS�f�z'䂔%�8x��J^���l�K���%s@�ek�f�Nb�)��H��)�E�סCm��*��I��jW�lk���yHm3W�L�8@�ȓ/�0=s�;r������^�������XZ�k�)8�"�"��k�bL���DQ��0�"5: �Vn#�|�ȓ	�!�Ủ�-�� ���8v<���5�1�c�*g(xT���Q\xTm�ȓd�v ����6YH $AcET���r���i��Q4�(��"oх:;��ȓ���2�(���4C�)>F<��;bt]����ʲe�Bfq�ȓ �ֵ�� ��k:xdrԮ�w{�8�ȓ� 8J!-�	G�h��Th	4/Ä��B��,ISnʇ/��`���Ym���'bў�|�T@V�P�-[�@T?]t0l�2�M`�<��DL#c�X��9=
�@ t�^�<�c��tn[���0І��HXo�<� �a�	PG%�5�Փy�\��"O�����I=0:�ׄșs68��"Ot��Q��� ,�!D��d�ui�"O���
�らr�$�?�6�;&"O�E��ִ 2A)���Z81"O#4dQ�r<���"G��"���G"O�1�#�ڌe����%XA�ȭi"O��R�+@�U J�I���<k���"O���R��T���!��R�d�����"O�X�P�V!7*��bK�Z��y�""O@u��LP���+K��1��Ө=B!�d�3���c	I�(���b��O�!�d
! pC���5X�̑҂CG�!�䖪LjJ��!��w���R�K�k�!�?������o� \.�y"f��6�B�=b�QI�&
&�yR�*:Pݻሀq�j@ 'E�(�x��'Z�]	�����	7���y{�'6X�w�M� ���#f.T�]vI�
�'->�q��D���@4釠\58��	�'yn�+��6$"�59�`Ѽ>���#	�'^<�����L�;@h��۸�y�aOOuZa
Q�H96*��lS	�y�	�ɴ劵�ƅB�T��B�؟�yrHS
?NTE�"��5��u����'E���3C�Y���"!M�r��'V�94���v8��kP�/y�*�'y \�ӧ*J��5XċYO����']"� ���<L��$�7�)B�':L��� q?X�@DL3v�uH�'��������Aq0�Q7t��R	�'�.��K�/�*��t�Hp_D�k�'q�Ab%G�E���E�d�05�ʓ[���G���;&���e�^9e�M��Hj]0�U�|<��E^�Y�B݇ȓ+R�����S���{�m�3H�@���n������6gH,�@�h�I�ȓ;��T��!�|�`}`��b0���#�����Cϕa9��;d�M� @bx�ȓC��a�%�1d��Əō�.y��Ah
M1�gK�| �sW��-���ȓ%;�1BP�9-aJ�Ӳ��<�<��2��0aL�h{��)DT�ȓ1�! 5@B�Yh���gG�������K&4�d�&Mr��Rc�ȽJ*��ȓ��d�ԧH	+���"�GP�G9T0��C���RD'Ai��*%B5:��Ȅ�*�eB%'L�)�|ɣ�����L�9�b� �TU�1iC�7v����o��@�-�� Z$�z�!��o�����!�]�Ջ�0:��q*�e�! 1���y�>�`�+�%#��sРT;�����Iv���ALԬC�-Y�C�V7���ȓ�~� CϚ/����qK�9+���I^?s�����)�5�<ecQ�B�<y��ʍ~��ɠ#Ā/F$�
3�B�<!��U�0����d�. :�mN~�<Q���h��X7��u�F����w�<�#"�NX�QΌP�s ]r�<�gk���u�Um�,͜d��k�<9�e��d��@��cH��p���M�{�<�t�@�',�Pjϊ2���%Ty�<a��:wР��Ls�h�JF�Wx�<�$�#P|%ypKŉ,����	x�<� |�(�d18��#�*o�@]�`"O��Jt팚j�$� �o�Hߨ��u"OdP[�D˛xq5��Q44����"O��"f�ʬ8�l�!%�	2N�ތhV"O�!i�#�"(]����B����"O҄��-4'����%8u�	�"O��@(� ���s#ģeS�IF"O���$/�z�$�1pb KK�J"O�q��mGd 4�a��
<Zp"O2����*�A7���O�8a"O�8eo�+��P��㕘$�8�b�"O�y��%��lPtBM"3���3"Ota�uµcQ0�:w���v��Y"O.)jסFDf��$�[>����"O�P���ْ2D���Tn��,���Ra"O�X��Z$�1�߁	�P�#A"O2a�J�C�Z�1#��**�~ɒp"OFȩ�ƜF����A�^3l��q��"O:�����c)d̂��&���"OL	�L͚e�Q���
#�@M�c"O�d;�$|�z �s��:Q�ř�"O��3)�{5�( A#�&�J�r�"ORliì�i�44��a���|��"On],]��T�dFZ�}EH��զ�yBgI1i�����B�h�{ħ�6�yB�G�53 ����%B6Z�BdO�+�y�
*,����a�(C�5$T�r�'2�� >|�Z�Bc(׌1���'yt��D��O2>@�.�"��
�'����Se�ln)�w�����yB`Q
����@T&sg���Ѓ�4�y��ՉA۾!i�^�6��`Si��y��T�Lجk"L�<+�����h�>�y2�	>��LB��%#4��V�6�y���8Er!X�C˴ZF�٠���y��W���,pG� ���;�U)�y�ŀ�	���%aߵl,`�	�yb� ��ݓ�	�<��A���@��yR��.:UJ�"t�B=$�Ip�@��yr�N�9hR1�2B�"t<	�g�A�y�߹Y
-�3C͂y���u$��y�I�=es�ar䔇�ά��.���yR����	��Nfְ�K�0�yb+��2�Dl�a�ݪ4N&�A��K��y�@�>2�P�R��V�����y��3�,pU ́�x�Y�(�+�y��M�*����ϒ�G�Z��$KF.�y�8���pG�S(K\����a[ �yR*�.�D-p�ǽC��H� K���y��>��!�E�98��Y�����yb�nR�����E�f �'l�2�y��6\�7-�i�(ٻ�D1�y��5�nQ��N��e�`�CŞ��y� ţN��"H�S�hlB��I�y��Р ���bG ܎@��	��W��y�K�(\Q-�D�p�X����?�y"E�+2�^A���c&���.��y�#�V��%
r��b[ƉX��ř�y�`��=���Ȣ���*�bpL!�y���C����έsB6��C7�yB��9��Y;r�J/j��g��%�y���TҰ &�cg*�#���y�F6�FTI�a�9\	�� _*�ybi�d�@�P��Ԛ0�zT�G�N&�y
� �!+V��+Dמ|
���!��!�"Ol��ǒD�������j�Xq+�"O�}a�ĝ'�����C�."#�e��"O,)g��<8*@1R(ڥ-j�"a"O�I2%���愒(b��v"O�ԃ��6��l{#ؓ����"O@)S�+�0<��)����#\�h�"O�	(6cݙv*���M�@��h�"O�deIJ
�,��#ܘ_����"O~���,���G̞�ɮ���"O2��dO�s���:�JX��Fdː"OB1�3�`�QQ�.	�H��U"O����H�tC aц")��q�F"O�X�E���a�(ŋ垳�K�yb ��}�}��Nߌ/�Yp��߂�yBH��:� ��c��'�����.N��y�c�d�w��! U��j��yb,R�M�ȀY��Ϻ�����F��y���w�4tx��V id�����yb���`�D%��fB	��DK4dR��yrc�K��Q���M�"���^�y�D��dК� �)DK����ă8�yr�ИB~ʐ�Lȗ*v@y� ��yrL�\ �,�={���#�y��*O{���l�4-��2&��ybe "^�"|��Ǟ A�8�!��!�y"TB4�I��C�E�6�y�	1�����NT�a�$[cg̀�y�Nw;�1q��-tF��sf7�y�G߶7 ���k��dF�Q�İ�yϻm�-����n��uH\�yRǕH~��[6c�+q������y��$��#-�2��q�&��9�yBɏ%Ai���C�*T��'^.�y򨈃M���p��].!�$�RlK �y�����Ԣ��
�|�P�b��y
��Z2$���]�w*��Q�%�y2��gq����P�4|�,��h�5�y��ʿ΢��Cǭ)���z�E��y2��+ ����"$���ε�y�LS�
��$�UL����y�� �K��l�����y��0
$Hm���<`�
艶���y���~�����k�]�H�&���y2ԃ%��<u�P�S��[5�yB�	s���3�&ڏ�B@������yB/5G�HX�k�k4@=S�(�yb�\��P �ƞ�L|h[Մ�
�y�� "N������w�3�,P��y��"} 6��%��# =�c�y�̷J
��ʮ����L�yE��,ZB1�TB��|Z�@��y��F#5:b]��H��|�8�Ơ��y��`�B� S��6IȆ�H7�R�y��S�a28h#��$I���#�N#�y�B��D:�`El�Ao�,�!	���y�胿+3���qj�>q�v��Ɖ��yҭȉ	�<�[�	�b����i�+�yK�q:����It|�n���y�!I�IQ�1����0yX�S�y�Hg�N���Ʋ#^  ���y�(�8$������=	fl�V���y�c��Wb,����#~H]CE��+�y2�ǩoS�5��m�^�lA3%�I,�y
� ��,*r16PÉ��}�W"O
�x�,�e��A�e'�Q����"O>��SEX�o^
t��eM�'_uA"Ox|�0���;��"�J�Y��aڥ"O\d��, �$�hܠ�)  �v��@"O�	�Ɵg�=)�"�8�@Q�"O�(��
 ��X�Jܗ0�6m)Q"O"ErE�݄������3�~V"OL���.
Dl8�X@)W�k���'"O~�u�͒$h�� �ٰ�lh
 "OJ��a���D!_�\I��2�y"�&K�����+R/,�Ҕj�"�/�yb�Iz�QCÈ-�d�sPb�:�y�	d�F��'�N7*.��%d��yRČ>HR�ũ6��/M':��Q�[��yB��mB��*ã�$;�
� Q͗��y�?Q�z�k�IA�94��C��ո�y�hL9
q У�� :�����0�yRB��@qb4K�C
�&��̲��V��yB�Z�n�`Z',9<�%8� ΅�ye�/�$9Y��J�[�vu�%�ߐ�y�L��_�\��@`*jHEU)�?�y��V}|P�r�9��c�� �yB#Τp���2{��lj󭆦�ybbM/��I S$W�a1�E�b�'�y�"N/��C"�2lX�� 2	�,�y�ɞ��5��!μidF:�y���Ő�A����#�.A��yBN�>�4��@�S�ЀC��y��<C�؍1�ȝ�].$2�E��y����.l ���W���#�%�yr�ڢg炀��I���c�&�yB�ķjJ<Z��[�	{n���_��y"�^�.�M���A��;.�#�yr��w� Y(�ؗz/B���M�y�e��%�8���)�	��M��M��y2�	�Cb "3� ��:�K�o�>�y2��(m(��Y��H䔥�<�yBg))�ɤb��A*�Q��.��ȓN���{� �#m��A �P���q�ȓ�谸�+��,d�,��1�DC則K���T�� G�(m���[�C�ɐ,��Y�J�-;{��
͕FtC�*�` ���i!��RB�K&JՎC��=]�,PzvDt��8xg�G�tJC䉪O��z�ʝ>=g�t������B��\b�x	7�Z�s`�P 5{C�yb����K-� ���L��B�	�E=h�*�c65h�C`'ޥ��B�	%_2�J�/f|dl�$)F��LB��0bh��٢d:�z��C���B䉘5%T@Pk 7Ϩ�H��C�Q'bB�	�uD�KG�ͺ��HD�#�"B䉴� ��6�E=��Px����B�	Ij��o�	Jc���L���zB��9eZ��Q%O�؜�G��^��C�I�8e�ya��g>�\��U�Z�dC�Ix�h ��(<��CᘃEb`C�I�,�"�Yv&\<]", R��^<C�	*a�2��q��
�@W�T"�4C�	�^����f��,A�̸ �9e-C�� x�©995��prM��+�$C�	�|�
�%!V<e��yy����
C�I
$.�@��˷v�vY#��.��B�)� �P�7�_�Z-�|��)��5�"O0 C��@{D��8󧙇LO�Q�"O�Q	��S,B�xMH�(^0$?��Sw"OJY
�I�#H���3K.j�k�"O�9鵁W-E��	�Å
�XZ�qH"O��3!G�8l���4��)E�"O�2�&;��i M�+�"O��$k�!=r����Ι�r��uA"O�-�!��iILI��j�4١"O������ >�ĺ2H�>
n"O^TR��-��q�ЏMm�"OH�X��0��(4(�V�T��"O�@��� z���hXrـ�y"O��)��^a��\;���Zb"O�+Qq�>��g��,9۞� "Ox���k׊q�.��1�F�p!q�"Oġ(U�͂Oа)���	;��I$"O���j	60Ҥ �C��u@�"O�xYTފ��a�Z�HTz����y�
���"¤ĉ1p)Ҁ&�0�yR_�o��lt ��	<ј@f��y�"K�]
jM80d�x�L���y"�U��	��k]�>��p��N��y�投.f�1�#�9z}�䄪�y"jA"&�p��4�]��jɡ�yr�
2���;��?�N�z����y���m�q�Am�3k�и��ϻ�y҉����HFj}BD�5�Q#�y�cS!&"L��GL�fͰ��H���y���Y�:���� 9X{(����yB�� dz�����"�j�K�����y��;�бi�uh�Q��F�y�d̒���Ȱt���ӤO��yɧ>�xċH�per���K5�yB
ܪQפ���h�� �l�3����y�m�j	�4j"�`Q��c���y��!Z�
	����OB��Ȗ��y��2���d�Y�-�^�L��y�D�"M��E��
X�(if x!�	��y�aW�)��)�B��6�����,�y�"\�T��(T�|�&��y�D�<��ѡ��ԛx@tᲁ��h�<�qG7g�:�X��]8&X�FȏS�<�ql�(6�\#gC�R,��ӳ��S�<��m�O`bH��.�/|1�ћQ�<�fB����z�ŏ/�jI@@��b�<��)T�q�8k󈙌v������t�<� �w�>,`dYu�Hũ�o�<�F�*;Fd�5'��f�T� B	k�<��9Z��ޖL�bT���@F{����"Ls��	"n��s�D�b���wlC�I2FF��2�C��]0�8R�� �U�>C�I9&j�zw�^0iP�aq���N�dC��`��˞��^D�0�D�h��B�I[3|�Ӳnł<�Z�@�Eί[��B��#q]$�;��{$<��<3c2B�	|����l� <e��o�S$Tʓ�?	���?��p+�q+��W4~����
>,���ȓ#��{�i_�sK�-(Ԃ��0����q |��A��vCT\Ja!�>ZԞ(�ȓR���{7�.��	�3�F�%8��ȓy6��Y��-�ġ5((\T��k��]����Xu�$�]/vM ���n`���K2 �ty�j)u�p��S�? X�@V/IRaY��K��.���"O��z�d�(~y,���JD1
@u�B"O�9[�M��EM��,� \���"O �yW�^�w�$}1�d'6� =(�"O6M:�C7<���aaK��l�r"OD��f��	)R�� �,��i`R"Oڸ@f�A�G�HUac���xي�"O��Ƀ��DE$8�@@��ą��"OV�:���?6(�*���.Rs���"O��Qf,?vx�A@�]B¡�"O�� ��Ÿ1;(�Y�h�/6.T��"O�麆Z� ��#�g��i�4�"O=#dc�_A��ȱ�|)�1"OvH ��cm��q��W�@r:1"O��*���='�R�p��$���Y�"OF��U��	kR����4��"O6���x9��
!}�Z��"O���˚�@It��2ֺu��t)"O�1or��m���ܚ7���"Ob`�Q�A7>���1L0:
:,��"O�b�遑; kA J�B�*u "O �ʓl�^�d�/S>TNF�K	�'���9��$%����c�A-���'r��hA�)���"흆"^jYS�'���&ʵc��4�r��i��%	�'��Bt�<~r,�rd��7�"��	�'�ư*���6 X��_275���+Ol�?y�yB������q ���0!��y2���[��|)RP�3��z�&��yB�'��!��%U-y�p���yb�:=wD!"����v۰�ؖj��y�"�z1�ܻw��>��c��A��?)�'�M������)!!��A1l�{�'�}K�E>_f`1�'3��'��i�2�@'5�v�)3A�&%�`�
�'_�+plؖ��I�lͺS�P�
�'Pb ���]p`�@
	"?�(���'ӒY���� �@�3�-� =�ڠ��'@\ E��4vX�|2�h��3��B�'�@Q�� R훶��/RF}a "O^��呇v�T�jbK/>N`ѡ]��F{�O�1OR�[��ί�e�E�G�3��)&"O6Iu�Ɯ@�qY�J�&a��"O�q�3q�B5��, ў���"O9�"��$��c�������"O�!Q�@�������l#���G��F��s���	H�,�R�^��9�/=D�x�4
M�N�f��DL�-^�A��9D�lR��G,&�I�Uڞ.��]"��*�d*�O���&iT�<����r��3G�|���"O�� .�7:����ߢ,�8�"O"+��@4���S�%Ͳ6�,X�7�	䟼G����E(�%��'�vTG����y2�I�E�"XW ��������yR��[��s�D��h!8�'��!�l�8\���p��T�9���)��'�l��d��e���� � �I�'`��hR
�>]�~e�6����XU��'K�Aj4[����(+"�����O�#~zdM�7� ���kY�*���i\�<����.C�X)اH/H�1���U�<Y�/�������)QfR�<�k�<36�K���LP�t�nk�'-ax���d\q@�B�*=ńH�a���y
� ��c6h\+ 7Є*	Z�0�ֵ+�"O�1˅.�Xy#�	7@���1`�'��ɼ&���Sc��.vT�G�B����PF{⑟���
N�9&J�p�CE
VA 0�2o1D�0���_?�1�C���h�*�$!��|R�O`-KW���;��j#`S ]A(��"O��aG�*���Z�/�%~8����"O�Z��ȑK�6�/Ѐ~/"O��&�˖y��䎂PI��Y��D{��6<t�d�C��M7$%L#{��ʓ�?qL>y/Oq�� d��G���F`A�m�b9	"O �j�����)�'!0���G��y�O9XE��/�1b����u*i��'�ň�-J=>ɸ��g�-�[�'��R�,�YQ�j(p} �'e�E�Q�:/�Li!����Z����O�#|���E:V��p�mS�c�	d�\�<)�`�<_��Y�X��%jԢ��. &C���%0"fǏyJ����M&jC�I6�*l(P`���0��s��\�B�I�-�jl�g�ͼ7�20�֭M�B�	�&���z���6�P��
Q��B�<] �ғ`R�X�����ȋ%��B䉀8	��rrn�w�W"�}�B�	:������	�(PX&A�y=fB�	<=��p�E�*��A)��L�6⟀�I@���TF5*�k�ታii^�� ���Py"�T����2ƪ�4�dx֏�E�<q��D��+(S���eȹO!�D	�6	 h�f�Gfɱ�A7+���?O��u�^��,g	��D�6,��S�`��I-MָSd���N�i�f��\��C䉳t
�S�i?��h@�J <���O��2�i>1�'�|ze����q���8w����'T>9��IB�d{�4Z�ˆp��C�'���	�:x�*�AZ%c$���'�X�끫��j�A �/��]��@��'��*u,u�Uks@[�Q ����'�PPr�-�>�CPjB�Ou��J�'�p` ���Gd�U:�[�5�.,�,O���4�OALH���"�		8c:-��"O	Hf]�\�jGHN���2"O���Q��7�Ȅ�)A+1� 	�"O��CO�`aV`�I�/?:��D�'4�	 j�te!�+M�hA$E  OE7nf.㟔��	$D-\�9u#d�d��!T3!��\,8��� 1�L"7%�(�!U�II���BR H3G��y�fC�tuX��h,D��0U�\5eR`�a��u���O)D���E�ܜ4�Lq1
��o����c1D�hP2n�4\�p�`f@]$#��f�1D��c,;�����1'XCv�1D��Z�̶�ƽk�mV�X/T��6�5D��ْ%���� #���6�Q�-�<��{f��a
[�H�����9����Z� Q�᩠�x2
��ȓEm���@�,^ڀ�@H�l���ȓrǊ@ fA;]��u�^~\u�ȓ|T��5g�ZG����I|����QJ�1jq�G0UE�p� ׋[a�ȓa�<�e��H��i�țx���K�'��8��*@���{#K�VI0�'LRpk4@��%� |��� *Zj� �
�'�2��F��%z H�@�F&<��x���� R��W�D���U��#N��Q�"O:�A�Ο�~�ڵ��+� E�QQA"O�E�C͞�S��D�*PdB���"Oh8 �L
�{>�k��IBB<,(R"Oi��m� 
Z��i��)�G"O�i�Т]-/� H�$�>y*�:#"O�ة��5A����(ϷLx�$H�"O~�:$��7��}��fʟ
�9���'1O��c [{O�b��W<�`�"OrQ�a �p�x�Y����F-�u"O�-�䐐l#pU�C�&|�ĩ�T���ɮj�&�#�xƸ�r�a[�wpB�D	0m3o7�A1���$a(C�ɞu6�ᨆM,���U��=�C�I�aT��V�6*@�R����d.�I�t�L��`ϙf����g�)3ƖC��<�pm�įR�UЌ��eH5I,B��M���J�	}��L�6ƶH��C�	�GF^ؠ!�Ƒ^ϖؐ�,��|C�	� T�pXe˘(,��z��y�rC�IJ:�ak��ڲW�n\�P��PC�ID� �h���(�%�6M�v��t�'Q�`Hǋ��u|�y*"��*��P(g�3D�`��YXS�	E�%� `�1�1D�@!���?���,,gH�����<D� �!@�nz�DZg�q�d��	8D�(��6Ufp�
O+ZP���9D��
g'��vʀ���9=}8h�'�6D�PV+��"�60��
J��h�/D�t��>;R�BW#Ɏ5\d�r�<����[�u���!@���ՅK�:��B䉯&Z����Ee�VƣE&lƂB�ɯ
uf�ꇃͿ2���#��# �C�I�hHPx
�E�!1,�=��eʋY��C�	�Zt V�Y
�v��
;P�pC�ɉ������)_�z��p�ې��B�I�*�|[�E2
�j$��bZ�T^���^�f@Q��:2|E�d��\!�Q�;�YՆ�(]5��ґKIG!�$�J9� I���� �y��J�+2�!�D��"�y��vb\���L�$~!�D��_��IQl��A�v��Zk!���̩5N��O�v-���E�WdџTE��53���iSdK�k��E�A�=�yrGɻX�ȵ�"��a�>��mV��yR"Lc���	�O����
��yr��>g�d�To�%K~6L2&��0�y�(ߛP�%��9M�Ps���$�yBDя�ʩ"�n� $�U
��y"0q>`)�e"��L�|�רK�y�K�#a�bB��vL��������y���U�����˂x�b$�3&�?�y�LP+6�*}R ��mL�A�
Z�yR��f?�Z�e]�l)�P�Em��y�,i6X�1�B�t�:=JU��"�ybo�}������i~��[�b۹�yB�A�`��t��8�&���6�y����U��yCČ�`���"C`:�y�G7�B%���w*�z1���y�# ��ٓ�����=aDN=�y�.� D��[�y�t��K�y�bDEO6��ů�!|z,x�#G܁�yr��[� �a��=u�|`�FL��yM]$z�����.6
��劄�E��y
� �%zec���/õD�&���"O�e�`�5N��h�-�G�j�[3"O�%K�AF&����!i�x�"O�x��»y���:VE��(�["O�AF�+�:���ɯ0I�4r5"O"m���{n��Ei��<���"O�L��D�J 8���c�����'r�݋��,p4��`�bFKpvdX�'��I@�+Yˠ!�b�S�.�@��')���P�Y�5Ͳ]��iɕS�%	�'���m<o$�r	�x	�'�R<���}ϔ�K���!.M�P[�'� ]���-D���2�l3�'R�(�%�N�5Y�Aا!�0}6D]`�'t�"�R�7ն�p@�5r�p��'vp��N�
��, *��k�楹�'�f�S��)�lp7˗�_��
�'m���djܶjW���f�J���)
�'�z\���L�<;�غ7��'<B�y[	�'�8c�/�/	��	3_P�0	�'9�X�ĝ/,�d��� "�  	�'�0�	f��([g�%(���$�(}��'8�i*����{6�Y����u�Q�	�'ː�9�eY7��i"�:��!	�'B���taM.#�0����:�0�'{���[���xRH�ER~��'��@9A`�
'U��	�$�:9� y��'�n��R]/ ��4+9,LPZ�'��܃��T2�<�Sc��%���'u�@��@�x�R���I[j�%��'�:��šV43�>a:�(�Z4>x{�' ��t��LMKA	�K2�Tr�'m�������4r�0&��<k|x��'�v�iw.ޖDG�Y���(:��P�	�'�qzV��[ߨ���4j����'*\�CG�� -���DT�<��0
�'�t�0��ğA�㓊]�2q��
�'�$A3��<�ܬ� i�)�pl�
�'`((�d%!��)�wc�U�x�
�'I�P����aL�e`7�ںM��	�'p��!���K�N-�FK�o���h	�'2���w�E?1~���H� �Z��'2�����^5�D�+�0b�'��=����N]�D��f��D���'�~A��$ʞ$�\��ױIjDP�'¼��|'����}�
�H�'�T���jI\��(�A)��e���k�'��D�q�ܗh����0�<n�����'i�٢G�5``	C�;p��a�'�F���1������$5qz�(�'��*i�7E��p,E���'✱�%���6��xC���!��'����+�\6��AЦ��)1
�'�܌bI�������F��	�'��ъqO�MqrԒ� n��9	�'�|y`���;fr�1p�U=n'A	�'��8�vJĬ�x�Itm~.����'�:��QF�vxF�H�ͫB|���'d��C��/|{h��Z�EH�](�'�n���a�8rx�]r'�K@��'�`���k�T���P�J�h�Q�'��Y��@@	8%���B�@�R���'Cv�!�MӺ=*x@�@�4�qj	�'Lp"t��ָ�10`E@����� ����H�![���r�(}����T"O��@EĂG�\X�T�<j���0"O��11��@�mрZ���p"O���E�E���q���/�d"O���▄&_��'�E0)d���"Ow�8<\B��I_B�iD"O��FH��.���ґH�-�1	�"O�m1�e�<D������#O!Z�pG"O��k�,V g�b\Xs@�"��z1"O�p����vz��"���^�P�S"O���p�U�+S�r��N�� QbE"O���e��C'*��0T;D"O �e2#��@	��#��xf"O�=
�
�d��,�
	�:�T��"O�*��A�����R�*�rt�4"O�Es�6BP��W���(�c"O�����"6t�H�N�[�N\��"O�\�S S2W�P�:��S�*�b""O�-
�׼VЁh`�2˰ap"OA"F�^��j��� ���i�"O�I��h���p�C�fo���"O��s��?b�2�awd�[W�'3��r+Ͱ'v�)�v��v�PY�o?D�H��I8�m�E׌j���ÆI>D�TA��*)l�+gO;Z"f�2a�:D� ��k3d|q�#��*Q��p�9D���@�:��4gϗa����9D���SǘlĘ��&���tF��	�7D�D����k$�*�蟼f��`�?D��qg�1�ND��@ 	WL�,���*D���6��2?�4Œ�m�)�|ĘU (D���գ�8W��$)_Qh��u�&D����k�^∰p���r���� �'D��x��*���]r�(��"ړ�?i�����8��ſ:����Go��iGH����'�RQ�����{�<IB^��4#�E�A�!�$��)�BYx6�ޤI�p@��E"`p�'ў�>�����u��!�a �:W��=���)D�$ѥm�(L�$uY
��S4��B�4D��A�#�;d/��1$l#g\!)�1D��!pڣ5��e����-���z�&-|O�b�t3Uf�}PF�j��G�ϜL�F�O�ʓ�0>Q�h�3n|�r- o���f�k�<��K^�~�)� &��vԌ��A�Cg�<q񠁵 P����Um�؉C }�<A�AE���Θ�r�ri����u�<Q�,��B���iM�U#jh��_q�<�q�ϿZ�1��.�<9J���Ey�<��M4��r4$5S�zQ �^i�<!rK�^�Ќ�է��^b^�J�i�<yd�W�h���6%ʪ_�&|�)�Z�<i#�C�!�d��u��:(��#V�<��'�1�x"ca��(>�^x�ȓ�d�W��)}�hW"U>�`��1����=�@�[��"2��utP�80M�6Y�^��u�D&Sz�ȓH�<L�U�!'J����A��K�ч�P��h�"G/}�<��Ш=q�8��^Fd���Sbx�bܤ7�I�ȓl�LR��Z� O���#�Y�8p�<�ȓ�"����Je�&(U�:���/�8e�#�=6>���0k���	o���)!��&�t���͝<2@ R�n:F���<AH>����V!�6�A�t�dp��:"�Pu�p"O� ~�2Û��������N����'��O�}�c����K	�^=iE�g����4�H;�c�>n4��꧂��9D�d�ȓ��V^�1�X�:�T��Ԙp"ON����%gB�{B�3'�"�Q�"O~�HBX `�g�!���30�'�$���V��x��
��"�:1���0D�����|�f-C��	�s�(Y�h�<y��?I-O �'��O�ʐ�0 �m����#آV��	�'��`�6�+g^���4��_c�E��K�Dڔ)A�]��H
� �(W]Մȓ?Bl�S��&IK0i3�	?5�Մ�l�'d��2�]Wܸ�����{N�|����?!��ܜa��
�����Bc�r<Ї�+�~P�G�E�|��E+C�N�W�U'�DE{��Ď�%5Jҽy�Z��P#h�	�y�D��vI��
�K�n袂�X/�y¤��y��@U�	?p�`�TO];�y2d���TXT!�lͲ�  ���hO�����e h�a�)���K܋=kr�'���'��)�3}�g�82�L�\�����L��yr-�>12�q����aS��ǁ����O ��O�� �g?���2�:�)D�Y@�0��F���0=)�l���D���B�ea��P�+�k�<�'��%�PQS��!�P��Fh�<�t����=H`Y�`qpgd�<��#����3�h�X؞q;���c��k�����x�B���1��.�<�LT�:ړ�0|�H�"8ހչ�C3^N�4�B�K�<Q���q���7��P>̘3s��G�<�a� P �qD#
�lH�@;�O�B�<�D��1y�T�H�o��V�qj�<��J�6`��I��΅|���r��Kb�<�WO{sJ���Fٺi�"t���\<�䓽�$�&����:&�J�#�j@������IA>-E��%�-�F"ܴI`�9A�K�<y��?���?Q(�D��<ib���U
�� NEd��eF�y�\=Yj�J�#D�f>���I��yRn�)v�,��#$\�;uȉ�L˨�yG�>�D�F�G�3n����ũ�y��ç^�HX�O�;"	������0>q�.ܗX�L���'�K�����O�'Da��Z%AR$���<���#��y"�u7����  �x)�`M,�y����;����=s�N!8�<�y2��)n�,�{v�C�mHP��@���yb�A�7Ȏ�4k[8��`�(�hOZ����l�d�����~���HgĒ���O���$Z�x��d�'Ak�f
E���}2���(FQTr� u�O�3�h�1� �<�/O���O��?�	����0@&� Vw��� �ц5Ԭ��0kh�A���^�~H!����ȄȓX&��%#�,lY�����nm�ȓ~�����T)��:�,U�����M�'�2� 3���X�E�gL*���
.O6��Dݣk�B BR�0x�|�t��mZ!�Wh�T%a�"�6�v�����.=5ў���_�O*r5��j�K� -���u$�PP���x�9��Xp )C y�	x�I��y�#�]�ɺ�I�E�t�5�C��y��� ~Z]bD�X9!�U�6���y�%X�?�,�XUlB� �tC���yKǴ!�HAy��U�D�����yR�Q*�����8yA�E&�P��	����@yr�'�3�	U�? Zd(����u�6�i�I� �V�a]� ��	�	n�Q�`�?0�RdE�>Y52C�I�1��j7�Y9)<����,C�ɗgn�-ѫK7w���S6+Y�lAJ�d>��|����?)�O��a�ą
�D�s���$1J��'N��l���OHp��O�<9dœ�ń"S\lH��'�px��H�X��ӎ�L��y���hOL��$�	�b٘ŭ� '� ���l��T�f0��[<����?K0�`P��Ku@�#��_�<Y�l�)d�qj&�>$��bwo�V�<q�L"��j�Ǉ	o\�rmMx��Dxr�	&4����Vo�\����P7�y2�ڄu�~���EE7<��1����y2χ�4JA��%��;ؖ0�ai�$�yrM#<�İr%�^;0���*D�2�yR��r����A��=$j4��mA�y�H�,�XSQ��73bU+�Jʍ�y�O#~(fR�L���R:��O��$=§�6mq��U�-Cuś��	�ȓ]��\*!' :KzXAI���;Ji^9�ȓ7)Պ��S;�)�ՠ6f��\�ȓDN���1	��1N�����J1~T@��X|�!{s臜H��� ��ބk32X�ȓז�ʅMDh��qb�<(4��DC�DɁ)��Tv�YC�%L�1�v]��sa-!�@L`:�m�V��)���\��D��T�`����g,�ȓ\e��uH+v��e*�H��۪���5+�S�#H7�m�r���%�ȓDI��r֨�L�N�#�aR>"`���ȓ�2�96�WM`@�fN�6
c�8�ȓLn�9&�	0�f�E5P�D�'��'��O�1�&M�A�C�S��A�s
׵i��D�d:LO����!Y���ᦚ=2W�-��"O�3".7+Str��I�eaR�G{ʟB�<�䩰����x��JD�Ő?�ȓC��J�M�GP�(��@�d�ⅇȓ$�X*��3H����l��Ԇ�T\8m�H��{��E4�l��ȓ,?`AĆ��%���` f�#26��ȓz-����V54�����-#g	�ȓ[%��f����h@ �U.#�`q�ȓ4X�3�\	����CkQ�`i쥇ȓ6w��W �!��	�w ��L��M����8�)�0�T�C#j��#�ͅ��Z}��#�:[3�m�s�
"9��H�ȓk��$إ q<�KS��pm&��ȓ`�X��ѢZ:A��)&g�	P�܄�)  �&�:(b*}��[�&� }�ȓ#
f)I��
�*�Ɉ��<~`2x�ȓ�\(�g��b�Dd@�g+�@��"���ٓ!ߢ���L�h�i�ȓ3P��KC�֏r[h�C��ݪń�?��� �<���xӅ9S�ܨ��<�(}P�V�3��yV���fͅȓ`���X�Ɨ�PL@�,T�a)0���c}���3گ)�ҁa�(ż��� �\�6�ǈ6���#I�1�̆��Z�Z��Q�Z���lI�>�͇ȓR�2!ہa�||��De�<c��m�ȓq�$� #/�&�v,�d$�	�D�ȓ~�B�2��rk4ᣴ�Z�D��ȓ�4Uiʐ�5��5���k�Y��`�:e�w�R.(���7��B�B���S�? ��#�1l����ɓ\7���"O&�Xa��-(d	b�]MN�R"O��A)Hy�b��D�Ҕ$@� �"O��P�jV
F��Kc̖�a�����"O�I�b�%��4y�_.4���"OpEA�T q#�d` a�)�J�S1"O&�����
TZ���&Z�It"O��@.��YlZ11g&<�"O�bJ�`֑8�-� ��"O��1��"h��*&�n��	�O����]G��*�  C.�`��3D�<�ud�11A2@	�#A
vʔ[��1D��y���}w�xx6�R��h=���2D��2g��$$ڮ��$K��.�`��E�$D��aD*�C�V��6+L i��`7�!D��͗:xC�xB3�J�[ �7�#D�ĸ��N�p��ܒgA8����!D�<��'�&V/bPiǪE�PA��` D��ó$�]24%٧�]�D�D����>D���d읊\�`y&��8H �Yh)D�HdXf~���g"U~�h�+D�t)"�>6<j$�3�3 4��@#(D�0Ƞ�3��A8��͚1���*�3D�xk1`��GzUAÌ�:Pz��0�2D�P`'*��8�r�a��+Z�:C�4D����/�13%�D
�AI�r�,�& 4D�p�§����< �J�6��hS� D���E�<�L�����+���3�*D�@V$�!���@�8;�rh��''D�h�@J0N��9�"��K��@`�%D���2�\]��zC��\�h��%D��cK�l֬<�/�<� �V6D���-T3�����? �=ҡ�3D���b\�g�2�������� ��m2D�4��G KeP%R�&�bNp��c,D�<K���]C�q�����Q��Y�*D�ĺ��ܛ[��1!GS4\�Z��-D�Xx&E�4J>�qB��і,l���-T��B�υ�u@b��	;2��"O,`i$� C�Ľ��ȟp����"O�	�2J
�<O���!*Ǽa{-i�"O$����}^�q 	-*{��E"O�ٺ7ƙ�q9n�ق����� 7"O*H���P� K(�<$�0Lգ]�!�T�pe�apA�U �,�@��'�-Ҷ	��A�ҳF:ufH(���Prso�/�u�*42�BU��y�$$.(�z�-�;`��ȓ'����(�
Pz\�	����#8N!��5�bX��F�\�ȩ1�O�-8x�ȓn8
�	�J�9"�xIE�&' ��ȓqѺyX��Q�j��xQw��u��t�ȓh����kO-)����(�8��>�,�rJX9["��5���#�t����2C�тae~Њ6-�#MV�������D�N`���vA6��ȓ@�s�Q>fPi�j�4�Z���l���4��>��ia��16�P��ȓp�\ه�T'*�\j�o<b��-�F! u �m�Z�0��(	1"�ȓWt���A�����H����
\�*���I�,��#�U�m��R� �"I|���&�3֦��o���S *1(���3b���"�˚HtB�Ƀ���݌Մ�S�? ��[e�t��y�`_�-�P�R"O.�95��hn��En�=u�`��"O��a��b�)83�קB.��a�"O(�J��D�S}�y�a��{�v�� "O�t�W�L�drRջ���>x���"O���$��=`��Y�VcX��B"Oʔ���.G�����T��b"O��[�)>j�ʘ t �����"ORQ:f�;3�$��jA���,�"O�飉ߪV���;�	n�(�xf"O�؂�C�k�Z$����U,^��"OX%H��1lO����C�(6�D�B"O� 0�b��H>M14D�2+2y��"O� ��ϔ�'*�pN�WT�kW"O(`xĊ�4��H#�,�#;QP�H�"OrW��_��
����i٦"O��#H��# %jG��GK=�f"O.P�,Z��,��iZ�s-�qR�"O�h%�Йq��`��	@ �["O���2+��6ÂIy�EH�LEl�2�"O\M "dEOM��E�M)RZ��b"O8�g�g:��7)Q� ���1"O T�� �=�Yx�g�N���:�"O�ʁ�) P�*���#��-��"O�`��`�$��/�-~j�"O�}�d � ��`�	'Q���3"O�	�wG�2VXDkMC�"BL���"O�	�K��2w���"U1�Y�Q"O"b5��@�e�Q���Zh��"O��+�(Js��P��["#���A�"O��;`�_5T��%@�2��mʓ"O�H���ގy:��0�O^����qa"O �`���#Y��!N��V�2C"OX}#pL���p�(�8���"O��U�0P�Е`��I+JW��J�"O��U�Po\v	@�DͿs&m�R"O,��c�C�{Tq����Lw��&"O�	�E��M�5��#��;g�E�d"O��J�ZE��%��+_TH�P�"O`�1�/�b��<#*�
T0���"O�Q����\�R(��.	�2W�a�"O�݈��Ķ�; �� r7(|�"OVq�� ��/qjsHN�j�u�@"O\1c���G^(H�����#�"OXQ��!D�O�����X$SX0��"O������\��)�tu?x��"Oܭ�a�Z/b��� l	�^<���"O$��S���IGB`:w�H;���F"O0��0\�9y\MQ d��>�x�"O���cl�B�`�蒓8�<�j�"O��i���I��¤Hܢ�����"O�8D`��yX�s��n�n<��"O��xD'W���u�Iai���ȓA����hY�w������jA��ȓj���s5���6�*a�E�֔���ȓ\�P���e���Q�ލBI�݇�@��th�(�=K$� ���r�Bɇ�I�P�y��]�q�5�C�(���+��̫�
E#wȮ�
f���L��B>��B� 0��Ɓ/m5j���';0��N��	 ��y����~�ȓC�x��bn�6o|i#Γ5�\�ȓq��db� g������ʀG��	��h���	�����b�>*�Fp��S�? �Ț6+oQ�% 6��2P��@:�"O�H0 %a��ʔ �.���"O��p�-^5N�\���
D�r���"O0�J7�W	{��a�c0�Z=�"O�X
!&�����C9��,��"OV��g/���qTiX
-��B"O>ɺAO(c|��G�QH�=:�"OB8�rN�-j�P\��DT?I���%"O\�R�Ύ�9d0�����54/ <�v"O����Q4Z���HU/�&xl�C"Oڴ��O*N����ԭN.[�L��"O*��Ҋ�%z�d����pp�z�"O��ˑl��4���b3́�@~��a"O�@���z@�`�B�Ȉn#�]��"O� ۔T~�FɠnR�d(�R"O��	t�N;wrl;�f�<?�u�"O������E�H\Z���� �<�a�"O�-)���f�Q|,��懇��y��Z@��q3�ѝG������y���+r�&��� v�~����� �yR	�PR:��C��WG�h��G��y�M�j�9�c���P�|�SI���y��Xl�u���J�L<t=SCʐ�yRaK:o@���g��y A�
Ҁ�y�\�~�zg��5|6�u�#H�y�)PYA5FO�ed�)cEÎ�yB�	�_ �ɩ��	�G����K
8�y����fҴ9�4ȔFJV3b��yR'��A]XjrED��Zp��yR B-h�*ck8V�1N���yBnI&F$Q�3���f�N��G]��y���1� axP$�ʺ�KwG�&�y�-Ê�����B���6�y"�bN��j�(Hl�q`d��y���X��<ó�\;2���bFǐ��y�*ԟ%r����R";]�U	É��yBM�"<}�įE.
�1r��y��tʐ����6G7���%G��y�.Ǥeh�T(f+Y�8^�1jf���y⌝�a�8��C�� UAVH�
�y2��� !��w$��q��^��yT�Z8�@[���96�|A��%�y��'M��q)SHC���oͬ�y��_g��8���p!�;0ʌ�yB���8d
�aO�8�@��yb�� �҅�hQ�Y�����F��yB��(@<Z+�\����(�y"��H�L���K
�$`� �9�y�/۸%�B�a�%Cn][���yCʺl�6Qb�ڞ%}�� #�y�"�̳ �V��x���_��ybA.6{D����P%$t��P�G�y",�C�Z-3DlH
�R�N��yBW/+Ιz%@�z�K�➆�y�T'M��%hǘ(`H��S�y�W����Y���GW��������yR��s�@VaC(tc�'��yRf5e���%�!f�ak'��,�yrH��=��KEA�*�:��5��y"��!@�,œ���t�ô���y2�\�5�@��is�芤�A��y�b�'��=� �,m�T��,�y��ܭAvZA�n"aZ|\C��F�yH�e�D���$ֶ��D=D/��S�? ��IӨ�54߮�4`\����c�"OP-�B6�* ��Խ&�<�;�"O�@�P�C/� H���E,��	t"O����*g���X�
�<	q���"OZ�k �X;M�\���+gȍ�%"O�31�5T�b��6+\{�Y
�"O6ESu��{P��2(L�1U� BC"OD���G����W�rI\���"O�,��%,=�!�l;@1q�"O�)b��4;���{�b�ʔQ�A"O�4Z��>k���AH�\I��"O��v�
1h�3�� z4e�"Ob�EP>�x�G��#м;a"O�M�E�I�R�<ڣ/�ִ
Q"Ot8	 �h8����I�6��"O,5��
�8��Y�C�/ ����"O`����G�]�B�	�@��QԴ���"O��1��M#��[%/�1Im*�X�"O�-��H6I�> s&͖�nd�H[�"O�Q���
b�,��޸h8���"O�M�@'άDoZy	bm�6*0=I�"O|T:2':6��Uã*׿_���iC"O�Q04 �OD�	uɛG��	�G"O�`�e��%?��Xم��"}��9�"O�qc�.U��D��z�J���"O�x��g�b^(�e��u�Դ@"O�����9m2�@� ��8��ѡ�"O��YU�F"��l�D�7[�����"O~�%@4��ěP$�/�.�"O�yp� ��}�T��a$X��&��E"OBd�@�J��!�b�ˈY�l�y�"O
�vB�{�ȫSb]�M����"O�镋��v�t�»7�xd �"O����-*2�Eh��� 1�|���"O�p�a¾W�`�IK\�tM�q"O��s�`�Pjx�������"O��0ABԿ�>d�QkY��\��"O�帕L��f����z
�p#�>y���)�/2�A���,IbM�G#K:�O�=��D�%!
b�hB�$��if8tq�"O҅��ū1R% .ܐ�S"O�á��N�0)[�D0""*y�"On8�a/�0A�Íh�q�@"O���m �+Z@��Č�#E�(��%"O�����	&��E􀎳��rt"O��2o�12���#�ݓi��c"O+͎>)��S��T�(�l�<�tH�F8�!Fb�s�`:�^�<1�Α�|���B�M(P�Y2�I�\�<Y��)����
�t,qbQ\�<��b�H�t�T�ŭ_�L��!N�@�<I����l��B-UP�ِ��Rs�<���SGz9�ЫW�N}�<��`F�<�cL-�fäjWS��Z��C�<��"θ)�$N�=�j��s��Z�<Q�ȘhB�AqF:+�R%��bEP�<��G�U�Ơh1�D=t�BrR�NV�<��)��<V�hxF�е_���aa�|�<�D/��R`
��d��"����U�	u�<QtIV�H)�+���(-Ht���	q�<����(�y�hpP��Îo�<q��I�Z�rT"$B!0Ab�z�hh�<IW��M�($�t"!I�|!raYn�<!�@հ3� � �CI�s��	j�*�O�<� R�c�,V��)#s�5�6EФ"O�\���� �e ���x�!4"Oh�F�#XD 0`G�6�n�Ȃ"O�|��%�3~j�T;�.ͭK��H��"OT�`��,�k7��5��0��"OV���6@��E!�%�;v$�q"O�!�l�-T6�0��$�Sl�@��"Of`�W��� �h�� �:h]"�"O\8�͏n���$B�{�!"OJ��!@M4 }�Dq�@�Ѝ�E"O���SC��.=4p���?ni��:t"Ox���$ƕ6Y4]����1\-�U�"OzaXSŕ�S_��q�G�7 )�I�"O<qxc�E��L�S��#�H�c"Ot�0'�68��37�ÕTF|�!"O�H�eD��S�D�<
Ɣr�"OdiR�S�y�$E�W�%F�98r"O�,�G�W�frDX��њ5���"O��!��Dp  )�m�:hfd�"O����z/�X�UOV�̕
"O�t��h�M�>��4l�8b�f��3"O����
�$���Q�i!�L��"O��Z88����3A�h�@#O�yb�I�rv&ت�ѱ�P�:����y2e���J�3�oM�	~��ɕ����yb!ӡM�B��w�Ѐ}v�!h�X�y��׽-䞙R�Ė�n������y�E#hu�̒���TXܐz�bO �yi�$QzT;V艆J���Ce$��0=ُҎ[#<��a'�v�\�� ��y������KTL�t��ZUj9�y�k̉��ij�`1��<�G���y��F�lY@�طi�~�k�I��y�L n�s�חj�bp���y��/us�䣳�T�f�8q�f�ζ�yB��:	*�RU+ �ޚQҕ�ҡ�y�h�~�8(��ν�$�����y��=:�<çG1~���U�̆�y��+Ne`��"�X$!��U��y2c�<���l��s�Dţ�y���Ns�;e�]RX��g]��yҌZ-;��j��G�����2�P�y���N;��P,�7r�:Y�&��3�y����X��TKD��^��cǕ��yr��xy�9�FQL��aA���y���gp���l�L��A�P�ȣ�y�$�9^�`�9w�^�8���d���y��ҳ5B����GFiRP!�ǝ��y����wE
�m� �V�Ǥ�y��_�K��4PԍT���iq��Y/�0=���2ׂ�g�:M��.2�y���^ɲ�+��� �){$Ȟ��y2�߶hxT1�e��<ڡre�P��ya�?CA���� ~A<���O��yB�Ѽ>:�h�c@kQhx���0�yBM�%B��P�Í�jV�љ�%�)�yB-�(*�Mip+_J^��I��y��o��tBe���__����F��yB_�A��HH��R<�2�l��yG�(�`�1WaԙE�lM�5��7�y�!�% "�,qD��B��P���y"�X'X ����Ħ4�x��W쏜�yR̫% q��
��"ϖ[w��&�y�2�F�	Qi�(P��� ��y
� x :*�-d�IV�܀ZǄ�z"O�-A�㙾e� )�$)��X����"O�,���5$�z,���^3��%��"O��/�<n��Q�(�"Y^r��"O�H&@9~�:�X��U/KE���D"O�}��Jh�Zƨ�2'ձ"O�$˕�(<|��0�'/W,&a�"Ohy{WOX�Q|��7!�`�<��"O�(k� �T����n���5""O�T�"��(�V�`��$7��E��"OJe�Fʞ)7� ;w�	7΢,�yB��pK�R���b���" �ȓEm��{��R�Ѻ��+%��ȓ7"v�1�Q<T�Va��_0T���l͢��QK@�<.�Q��Y�h��=�ȓN�,Iy���q9R��B�X�I�ȓR�)⦯��C_��-^�/����"�<�A�J!%����kճ5X�!�ȓh%�8:��������$5�A��M��УG���d�և�&�E��J�L���+�V���G4:Ʌ�:b�C��\	�h�Q�~I�ȓR�޸wD�p`АI�
t�����{�20F��LK6�#�������ȓ@[��`f*�Z��d��@>H�ч�7��I���ԶQ]b������m�ȓq��,�@�=�$(H7L�=g6H��H�p�q��	5i<��J[�3t��ȓE'b<hd�Z`��e� i�C�h$��~�h���*x���#�߿����qx�k���:E��k���\��X���R0��I�p�C�.�(%$����w�L�`��M^�q3��
��)�ȓfc� s6����^�X�c�}S�%�ȓOH8�6H�kޘ��@d:r.��b�( �pc�8��e��
��<��'���g�'%T������v"O���Jߒ��Z(��t��"O��"f%�YrѹR�
� �MI�"Otp�O
�4tT�dXZ�#�"O���F:]�L{6�J�W�9�"OHH�%�\�3�ph��OU>�å"O&�1%�2cu�������"O4��L��%�J!1� �[��p�R"O~��K�B��u�s�Z��
��'�$��&�ƮP p9��ޞ_~��kWK?�������cg��	�'c���S���I��X����s�`�	�'��=;fI�*Y�T�L�1^��@	�'�zub�A��V?�1�.A2Q6�(��'!<ݙ���($�H��hJ�'d8]x	�'�޼�@��O�Z�[%J	f���'�z�C�̇ @v��c A �Q�P���'���z�8k1��c�f�U����'Z�XUH��	�L��nh���3D��0��Y�D�ְ�dE�,�|07�*D���M�l(� [��B�q��8��&D��З ��!�Y��%��w��V-%D�4�J4m?�xժ�9  ̅��%"D�4�5�%�T`�3F_2P����,D�Ly�GJ���@�)eBa҇-D�T�@���9��9��؊Z��`U"-D� ;�-\�s�d|�j�${�LCTj,D� Ơ�,;�aKV/��G�n�@f(D�P��+W�s$����m	�#@88�n*D�� pqm�)!�C��O�{�P�"O�\��Y4f�~pA��9ak����"O������2��Ʌ X�W� �C��$W��S�!�9[h��}���/,�
���</�4Q��h�<�#!�?O ��ʂbB,o��p1MJ3>t��4`L�-)$���	Ѡ8�~&���J�R����w
.PtL�k�'7��a�F7[��}��@̉���R��8�h�T̶�S`f��K��!�r�rQ�@ײl��]�1�:c ��	3��i��nJC���9À�9D�,ega*P\ �Ԝ<L#�% Vh<���K%U�9� +W�D�N�I0�Vy�,,]yQ�Aw\���E�y�2��~�TgʵW���CK4Z��q��V�<af�ޱ	��RM܋N������We���`A�-�ι��J
+y�p%>�k���T�L%t�L�#���/Ω�Ѡ� v?�~2�]�1��m:�C��l� Q��V8$E�,��P:���f��"��Y��r�Y��$O��Њȃ�D{�M�]Ͳm�f�I���,��.�5�y�U,ڴm����շi�8Q@v���&R�6(�b��[��x��׼�iR�M~>��4n��yb�'A�<����H�Thh'Θа�A��	�O\(�4��-L$`"�KN	b���'(�i���Y=�	@���0vl9"b��!j��E�؁D�X)Sa������� �-�r��<�5oW���|�%�Z	�#�I��ę!f��z�<|ġ�(����A/�VW$)�b�5E��ӂ�� �X��P)\G- m�<y�����\o�ӑl
���O��"�M�L�l��&ḱx6�aq�/[��h�������ɐ��
d"2�-=�L��$�f⺄p�*]�6� �fA̠\���u���P3*Sn�8�E�Ɩc訤H���4�$������v��̙�(μ\��{�"O$kDˀ�*�b7K�b�YB��òA���Ƀ�wA��B���1���W�x��B�{y��U#(e0�B�N4&��H�R1�0?9�
ؕ.�ay��F�Q��h1q+؊"-��EV2cx�a��Ε���`R��Z�h�1�W��PY�򁄯�z�`�)%��]��ǟ��O:������$Ҵxe䙹l�Jɠs��\��r"�F�~�,���ۊI+$B�/%�n6��3rtK	�\�Dm`�Ѝ`�(i�#T�a�����8&o�u2Tuz��
Z�RE(�LP�c� e	_w��m���캛Уk5:D2̗/�D�F�Ch�<&�u����l[�d�a�U)�.vm��8��Q°}8`��X���:���v��o��Av�b��&��A� (-+�8��F灛{�F���M=v�",A�m	q�����@]�4زTn�f��TA7a*{ЀJB�H�|�yFjh� 0��%����'�Fh"7��1�<�K�o �h�ب��$Z�L���R���}�m�1?za#�)�44\C��֎:5��q�i[�b�0YcQ�����!G�8�a{RӀA>8���MJѣ⭑��y��Ñ.i�I���.����&҂E94ْf��L��͑);g��m�77�.��4(�B��YiR*�$�y� �?��<0J��1� �XR�G- ����RT�C�L0��C�T�i0�(�h�O���	
-;�h&R9��'�`� ����W?5�I�!ȓ�0QL�C�DG.@�v�[!�]��0�"SE�;EIv���,i��P��w ��5S��L�է�ej.؈ci�	����˖5Z�qVn�~��T#�٦��Z��_W(<ٳ��&I0��H	�dx<U�ӧLyb&t�Ҭ�&y�L���.O�h�)*1��9(
0�#1GZ-�9P "��B�	0Aj�����:��\`�e]N�;��Sk0�;PH�Z�,��(�E�	8;��		$�Y�mwؤP��
4h�VC��w�p9�R�HVV� y���(qMN��CW�.a�$@%e	f[����'��U�fG�.-1�	�a�v4e�
�][f�䣎�!;�d���>j�,��@%
:��Z#�M �8�"On<J�"��"֙81��3/�$���䙳/� ����F#D+0�}��~�ի�Z�F`|��&�^K�<)��ߧb7�iaQ"�-9@<@�SK�F�<a7L�83_v�)�cX.�� ��<	U�X�l������6 ��1�(�t�<Ѵ'�ڼ��Ն�d� !�䪚v�<i�#��l��H���B���.�ȓEޘ1e����Le�X�1��q� ��b�{x���r�U������a�j��!#�g�^u��i��hjCe��pd�w��(k���L*�5��#��@���I�jR�p�nф��l�tE�o��)���:}����S�?  $ѧ��,T���IǦ�+X�=A"O��BQgڸkݜY�T�T��kE"O�!j���IĬx�R���A"OPqK��ȅ��)W���"O�q[�LP����� g�<D�@}ڔ"O�!��۟^(L�C�g_�o� ���"O�4�H�x_�bVǟ��@�K�"O(�c���:��w&J�a����"Ot]��5��\��i}�y�r"O���b�*㮄Jf����"O��w��8&ĴRf�lo	ځ"O0��O)H�D����YP�|BF"O��[���':l��� �6aY.l�7"O�����Z�h�P����R)44.)؀"O�)���C"T��`M��v2"O�H
4E�!0���o��$D"O�ȱ F�/cm*��O��@��L��"Oh�{A�%��59���s�v��a"O<����aW��
#h�U�8���b�x
ucK���'�$'ɘ�ȓ :�Rc��?f��D���X�)�����FxQB�M��i%��3 ���^�\H���J�&��ӭ�B����-�ʅH7$@�GZ)��oJ�h����VAr�&��tD����Jȹk��E��.&:9���X��b�f(�}��q�ȓ�%��CһB� 3O�o%����,9�c '�T�R�H��.Cx���J@f]��e�-��\�W�
� UC�Z1\aq*D��(y�oX�o��B�	�`�J4;ㅓMXl}Z��=2%�B�I�{����åZ	T��D�)4�B䉲A��yIGE?�uZcA�	B{zB��- "�����6�T�8��s!B� %� б�W+n���$&�=�C�ɦ!�4�����.����!ձTmC�8c�t�$�������b��B�?d��ё����o�hy���ί
��B�	�4+8=�d���б��6i/�B�	�s��YSo0� �� QDC�	�b����ʖ2�Ry�3*�,��B�I�s�Nq@MS =)4�:� O`�B�	�u:�a8�m��&z=ᬗu��C䉴��]f��,J�T�!B��6�C�&���
��j�&�B�N;$��B䉓����҈L-�4���	1�B�I:&D���Ņ$grv`��gL:M�B�I
`�`S�0�P��A:9lB䉕/jK��d�x-k�N"�4L0#"On���J��Y�F�mqR���"O��J`k��E��`&E���L��W"O�X8�gR) ־z��3$�b"Ox)p�,�;$D)�dH:`���"O |Af�a�*U�֧Z��k$"O$qp$Y r�`}�`�ʠ/�P9�"O�������xaS�N\�MY�Y�S"Oh�a6b�?ld��!�["� ��"O|p��%>���ч�*�86"OB\���	G+�1��/>����"Ona��"Ǒ3m�����XX`��'"O�;�C�S5x=��@S$���"O��ӳ�)�*8�4n.K�:���"O�M�d��7V��#�lg�Ԡ��"O����5M�!�+L�Jz�e�A"O� vXR�iZ7ӊ����F�4��"O<��ǩ�:2�8���*@�U?D��$"O��S@�S�G��$(�+%����"O�PR���*L�l	�GgǬ��b""ON�C5.��n���87� 3ˈ=��"O�"`F�l)C ��j��A�G"OX�*�,`�����nD1"Oؐ�m�Xg�0HqO�*t��G"O�БBJ�꬙���Q�H�!�<��C�-� "�`�D�&!�A�z�f1�ddюB�����ʠ!�D���������9x����B'G�!򄊴 �8�+J%hz�R�˒.�!�$�(K�v|9�� nn��!ah0�!������9�HQ�i��Lsх��!�D�H�,%+!z�1uD�$n�!�d�7ksX�p�E>1j��ᄔV!�^�4�i95��H�d�@w%:d�!�S�z�:YsrC��yHS��נ�!�@�	���J����CV$	!�$�%��I�(_�/�:I�'���!���&Y�}y�̋�¬{P �n�!��I�~&��:%H��N�#$G|�!���/�"|�R��Val!r��f3!�$��q"��@6쓈Wo�B�ȉ6��d��)|�<��M�b�ܸ LL<haJ��>S!���$ �JT4�3�&��jM!��W���5�g�=N��j�!�D�.a	ѐ�ʶ�~�mR?�!�Ď:f��,ɟ4yJӰ�)v�!�䜄 y��c�	�Yo�2E�S!���{=,�Q�S�y\���"��0*!�D^<�ư�փL�e�v�A%�Ց\�!�$ʩ"�r}����3}�T�JcF�9*�!�d�
]��q4)�,���t��V�!����4���Cȶ��,��D�!��#�vL#U� U���tKރ)�!�Dؚ]6��r�����ThR�,�!�H�V��4	�"v��	� �!�ʃ���iT☮+uz��&����!�=��E�A
�<a*�2�q�!�԰o���S��C�IY�x�*�	�!��Ɋ0ʸ��$S��U���!�d��|҅`�c��[�& *�a'�!򄖄Шl+t�� +x��!���
|�!�d��U�- %�/&�h���L�.�!�$�b��C���bq2V �
=!��0)Bl%��Ǔ�Vj���ߐ8,!�� ��+�@�=��q{S�U�`!�$�<^�̱�]�x�r��q ٔ$�!�$!g��.��L��O��-Z�"O�I��@/m�X����/��4kW"Ot@ t��$z�]Y�E�x���K�"O���^�59�j���~oX��"O���թ���P`dֆ=Yb�8Q"O\5�f�қ#�0�$��f$�yQ%"ORY�BOsj��c8o&0
`"Om��k�	b����"�:��"O��jצl�1�� ��=�JU�"O�������@�,�&_k��b "O��*7�6R]���I�'Yx|s�"OJ����%Ei�L���=R�"O��H9Ժ��*�36m`嘢"O��� �qۂ�6���B%/!�� �y��֢1��D3�� ;s�`Y�"O<@R�*2^�Q���zP����"OJ�2%._�cI�(z��1dJ����"O���TN�,T<����	V�}M(8�$"O����M_�:�x�Ì4:С(F"Oh�cs�Sd��S�,4V(P"O6���I�"+&2�Rq�yKƦ5��"O	9&`ǄfM۴%D�.|���"O�*����ψy���߷#�}Y�"O�añ�4s��{���� 7���"OR�Bqř�(3t�K�<!Zy�"O^��lB�g����` �6�p �R"O�) 5 �6��xg�^�}��2�"O��vk��x�aᐮ%��a�"O���U�Y�t��@�6`�N�� "OsH�BrF��`D��:�,��"O�X@/��(S�DZ�&�Br"O���G�8(��ҷ�@�N���"O:Pi�-Y�����b���K?)�W"O�$�/����e(p�=D�� �Jo�B����9#�p
"�5D� ���$
����F��Cؒ� ��0D����Gp��q��d�c��,D�����FF�dy`X`z��2)-D�,��S;D�����EW<'�Z�*�A*D�<؃&�Y�,�@�F�X���,D��i$����R0aF�f�450��-D��x�׷E�p	� ��&?~�P�7D�`��J����
u��:� 9I3D�\��� ��	��OD0=���$D��K�@�Ed瘰S����"#D�8P�m_�1��i1���<n�x�c>D��#�N��%����
֒RptD��!=D�(㠊S�t��b&�j6%-D�����#8=z�ӬK�.�4H1D�� ��Hf~�9t���at�R�g D�D!d/�{�t�so75^�Ɂ��%D�(:��I�fH6p��N̼4�b�E	"D���6(�,o�vP �%p�#�"D��"�B^jt�����3�2!$#D��	&	�7w�D��A�w[�<I@ D�T�uO�=�&t���)g��h���!D��H��P��H�
��ec�k���
�'�.���P�%{օ[0�8��	�'OT�����iW�������'enU2 `��.�ҥ�X�a���P�')�u�1G5 �P{5@��o6L��'���'LC�l�|�Ri�[:"�R�'��iq 	7Y�$�#؏]78��'�\$�gM BkIq&K��G���'6L���x
pv͉�9�j	��'�p�1Ç]W��h�뒮5��K�'���*�+��	(�B+�'w�:5'�-Ϧ�jPN	�r
���'���A�	�`�P ;��D��h��'�ځ��ȩ=G�xV�H�#��l��'T����J!�����V��8�'޲�ҕ��7]Dr1J�@�-6h�c�'8-"#��4��F�!��+	�'�L�� �_�(����Q���'ڀ躃�	n>h�Ñ���`
�'�TxT���ilAÐ��li	�'�^��I����&�ΟwCި0�'Ć���T�4�l)��Re{��H��� ٠�M�`D�pP�@Z�u�&�T"O�	��"<3*����ن_�ȣS"O�(�v@�=0��Ӣ�؛;�&L��"O��	"<?��r��-צ�QT"Ot�� F�qG&$՜�a"O@i)���x t�Z�l�&��Չ�"O`���R�	����aC/4�DH�u"O�p��D�8.�GO�\��	�!"O�)�l�,	�mi��@��l�"O\$�b�V
�qb��5"� E"OP�AE߅sH`a�-��EP m��"O���Ȍ:@�ex�bЬ)�Yg"O.�	&�+">���kM�(6"O�Q��(JJ�S0`̭_$��:c"O��SV�C^�C� �tb�d3"O��3!��p�` �O^�^Fab"O6��Vi�+8�%��nM @�<��"O ��勔5BR����@�n"2&"O�T�v	ֆZ6Z\��,ؤH^��s"O����Mǖ__$�[ęV(l�1�"O
��L�	~h�pa#	��Sh<ʥ"O�1�
f2��7Fº�)�"O8qk��U$��tA7������;P"O���5.� \O@h3�EX,�l�;�"O4����	�H,B�EE�&�"O89����:h�����B6o��#�"O ��`�k2X�B�>��]ɑ"O$�Ica�'0�B��EBQ� l8�
t"Oy���T|J��'��#GB��"O��YA��$7"�@d��s��Ó"O&�S��M)'q��`&�� p�z"OH��F%V�#�F_ȰA;�"O�`�d�:�7�¡kH�A��"OU�)�.,� �V��I8��
�"O,<����w��Ĳa�Q���D"OBA�S�\�.U������cyf�q�"O����J�[�z�35:Ji��S"O�m3'ĝLTJ��ĵj�.�"3"O�)���ИT	��E�-G�-aE"O��5nL�Vvn2�*����"O`-}�ԋ%��1��L�GfF��yB��f��!���8��YyǇ	5�y2l�	)�2 v�"<p,�AF����yBAڷmi�ݢ�E+���x	���y��-o��]��䃽3�
%sUmE��y�-��H�gͽ֔ ��Ń�y�M�[ihc��b$�������yr��!̜A�)�Z�6(�#�0�y2��)A��9u�_(�d"O�P�.�&uP,{�5kG�#�"Ot@�Tc"�i��C�' [�"O$0�BΟ�v�Y�@��$��b�"O|��O�-����ͮQ�-br"Ojr�P:��[��ϣ�<|ɕ"O��8�ֳ�R��� ׽2��@a�"On�3�F7��8��ќ2�|`�"OZ��G�x��yj�H�$"��6"O�A	�k�=��gA%3��M�"O���c&[#u����&9l�r�P"O$�8�.A >������aG�e�"O���Ca�I�يFj=-�4Y�Q"OM��� 
N�ţEJZ�q��4�g"Oĵ�p�ڳ=��T���+C�Θ�S"O0K���9TxQc�o\?;�*�r0"O� T8��G8j&*�n��K�th�v"O�թr�K�v$���a�ܩ	Ӱ�+""O�ę(ԵQ��Ur����(֪��4"O>$��Ș�X�l��5�H28�XȰ�"O�ʳj	<5wv�@@e9�`�q"ORi�VJK'���P�e��`J��B�"OXI�7�	Q��5;D��f7��D"O���4d��2Ҫ��-�<�"OT��L�u�9l�HQ4!V:c�!�M?n `ǁ�/nz,xh��4(�!�^�b��d îҊ@B
���b��!�$�򈴣EۏEL�+!`�w�!�E�d�FQ�߷[��]�s��-�!���3gNl�A# ͔1i��0�@ō/�!�dN09s�J�^| �����!�P�6 4y(�
;
�(BG3_�!�d�(��7B)>1H|�sǓG�!�ݢle,(�G�גk���@W� ;]�!�ğ�Y���Y
քnw��PU$��k�!򄎩D���"�@{��˗�<�!��K�.����f*kjj%bP��24�!�dR%&.�q��`EZ��s'ʟ+/!�dN8G�9�񇆻]��i����!�dծ$������k�����mi!�D�?\���ưLuv��-��]n!�Ǩ~H�J%G]�)y��е@E!�$�	!��!��H
8���:v�P-m!�R�f�i����*A�Ug�?o>!��=h�����1\��ūQ�P�6/!򤗽T��2�O�?c��}��B ]�!򄖨��fkKn�̰��:�!�D�<vƍ���ѐ&U����w!�ę(X&�-#�Cۙl@J�C��3!��7	6�JsdWMdUPĎ!�� ~�ɓ�>ՠ�Q�Č�y!�ğ|��a��B-�p��c�a�!�$W�V�ԝv�O�O�`EB#�Ϙj!��L�0�B���bX	p��㖢��!�d�j>p���K��� B��P�!��
c�hyE苩2V�⢕&!��ۄl��(B�Rc\Tr����!���#rq��"`^�A��%	��P�!�J�`{pr$Ǒ� ������.4!�DI?��u�d��B��u
4FųD,!�L�`b�X��$�Ȝ�{�'!��܁r���foٞ���r� 0�!��l��Ɵ ��(�'���]�!�dG6[�|tS��F�L􁪂MդF�!�$loڠ�S�Y��P&��?�!�d��-�ΰc%l8)�ȡ*Ņp�!�$� ^�����o��:��I��^$F�!��T�<��;�L�	6 3oU�	�!��[��HL�s����	��ճT�azr
Ǝsp�87
��lЬ�`��"Ip��G,~ x�-�޸'�8�NO/5�M��O�Z1b��t�	�f~���gj�p�[�Ǌb�2\i��J{�$7�aʞ�PA,;��xQ���'N4r@K��rV�ix��ȗ%Ѻ7��	Fj�A�ʹΔ���}�Tdy�-ƀS��,��W=����
,��`ʓ:��裡���D�T���KE ml�,�6h��O�J�S`a�;T5���h���;���("X/*,B@��N
�}v0����b!�'w2���3o2��k5�Fw�:D�tͣ$��8��}�Ic>��6c��kQf��6�TE�jh�/�ɢg4�T�}J~J2�׮t�(��&E&jxi(QF�S��
L�(��>�ʵ���X*��stmQ)WX�I�K�F?Y�g�#k��O�>�	b�D��u@$+Q8e�L�)0� W��I�$/�g�? B�"��n0�ӷ���+����Q� ���'�Z��'>7��*��Ť .b �'��>���<�7�Z+>���b>]`D�Ct����$վ���1�6?)��	*}Vc��?�1�G��:��^�*Ȓ�@���&(�9�اh��x�@*�����&��A��d`�H�	�@-��}��� �I3�T:��	(����/�-s���}b��b>����.V��2&m��#�,]*��"A�,k�}J~J6�!w�6p���xȄ\� �E���F��>�OV�I`����v������ ��	���I4s���GGA�)ڧv.��G䚜_j0��bD�{b8�pǒ�{E���&#��R얡qУ��"Dͩ��	B`�)�NY�<�'�Ć�<�%��x�|Ҷ ��TDF��Кx�MA�m�����S	_8�YM� )�^�B�[}�ZO�x��7�ay�M�)AI�(��`8�E�Y�y���H�읚����Ơ)�T#�y�Z�V� "Ō;WvM�$F��y��+.]F9�ŋ܀E6&1`Aa�;�y�JS*$6ʔ��%ۻ:�x��p�O��y���q؁J��>��=Y`�L+�y����8F�|��L�ߴx��̓��yb*�joȩ���X��z�a0����y�C�L?d����`A�p/G��y"BѭP0i��n&T�\�RG"π�y"�ɻ@�sV�F�K�`0H����y��ˣ$��h����9sպ���Z��yꊣN:\�d�|��ڂ���yHJ�;��%:� �2 �*`b`ߋ�yb��uP��{�z�p�a�3�y�޷\ ����]+ f@ �y�c���^S���SǬ� �y�o�<!Шh����) ��C+���y�-�	z��@_$�5��H�0�y�A�1�Ƙȣ჊:��X�"�Ҝ�yD���*�S��Ȁ ��,�g�Q��y��#��e�ă� �"�������y���	2��;�ṁb��x:�K�y��1p����eH[�ȥ��y�jN�i�Kk��;��q��(���y��<�\HC��]�(�X�weU5�yBIŷ/�\��Ql�%���)6�6�y�'�)t6��4G3p�,<��'L�yrfNd!�1��#�0gpҡq�ˬ�yB��%�p|��/Ƚ1Qད�Ü��y�G�a��	
�*��wl��Ǐ�4�y�#��Z*�0`�Ѻn2� �G#4�yRa;]���r���a�̵
&���y"��`LPR/�<%���eL�y"���Qp%�%��+	-��(��Q�y���8y��Ms�斫=:�bd�/�yb�<]qb��o�2�>�"E3�yr���1<���
�:��ʥ�y�֑Yo,�l^�.6�dC�4�!�$t����lxP�Y�p�ǸH4!�dN�0�VVOJ��h��'!���0=�r�J�� @Խ����$!�Ą$M�ܲ��s�0��^�y!��5&[e���F�"��`uh:m�!� ���	JG!t�pA��'ڃE!�$H�^�}��
6�>ѩ�D/V�!�Y#:����;h��3 Y�O�!��-;����QE�<Yj|+��V2"��	R��t BϾI�$	��0�!�F`1D�p3�oH��d�:B�E�x!���GI;D��87�G=/��$@����B �7D�� ���F�FuzPcc!��Ȉò"Oh{V�1r�	�-��!�֙�"O�Eyaf\�-���I�f��|��!J"O6]AF�M�77T���Q��l(�"Ojȅ�U2Z~vyc4��q��"O��c��,���IᏄ'���"OΔ��H�3��{��P�v�����"O���s�A�č�!���R"O��X��Afb�B���`�̐ �"O�h�E��f��pBs�_<��8�A*O:��M�\y;dU��{�'��a����I@$Xw�t���"ODM�T���
�Ja��I�&��"O�i�w��#�4TQ�I8i\
�)E"O�� "�[,�R�s�� _Q�tX7"O��r�oN���`+u���2�0 �"OViqW,S�w,|Q�bɵW�@�"O��ҵ2�����$�����"O��e�tbT��ӭ��f�>���"OM��Bt����a,N l׾m��"O`YJ��M���	C��H����"O� �������Ӓiرg�
���"O�8����RvH`"�	�3��l�q"O���4�	DjN�b�T5G4%�B"OV�*���:>�x��v��5>�T�"O��I�P%������,�r�iR"Od=�膕Y�}IVm�pƦp@t"O�@�ҙX��U#ʳ��("O�,� �ˮ�ٚ��Ю/����"O� 0f[�@�y8����j�$��"O��$o�@uHy�����w�(��"O~���.9�ڰB�"��5"OP4���0l��t �A�;	�����"O�}�r �L��A1@��"��P�t"OL OLs:.��7�ǗSp��
�"O��Qc�r����e��hr�$�S"Od�H�zx��a�T�
t8Uj1"O�\QpEC�Q�~��fJ�l� b"O�ݻ���rHy7�ٖ]D͈�"O<u����#t�y�	]����"O�1S�V\�ƉQE�˃}F���"O���Ai_Yv��p�B�(J;��ѕ"O��(�f�2	2���c�L29�u��"O�ŒP�̮L�2�â*U�/��@"ON�5H4�,S�c.p��"O�<P$�M: >�`�:
;�x�"O�-�s�W1'�8�uCʰ-;~Ѓ�'�Ԅ�Ti��k��*���h�xa�'�6�9��G�T���@R���yZ�'O��K@f ]0b�\�2��Yb�'��y)�#B�Y��U�al�zT�̀�'f�pcR��~�ܝ�`)O0y�\���'�`ٛ$*�c� �ʱCԪleex�'�P�ۓ��s���@/ǥ<)ha*�'� �Ip�8���C�MR%F|����'�*��,G��p ���.F�C�'�j�9#�ֈ<0�]�To�p�����'���	IX!xi�d�
`��z�'����Vk�@]�aJ4�$fe���'쎤0V���2�z��0��?X?�
�'.VU��ڇ/~���&Y�%���	�'Z�A,Z�X�&��`��B0�k	�'�:�8���m'�P"���	�'�&���H�TL6Hyf�S:��Q���  �1e�1|L�@Q��W�H9*�3"O>���	�B�� D�9@X�0�"O��;�@���:ղcY�'�,���"O�Є"?ȼH�H�FRhq�"O��	RƏ7]�I��ޏa<$��"O�!�E�(m����cB"m��}��"O�d!&J�>�D�0B'�<�` ��"O�qVKԩ�)cg�	 ����"O��R�D&|������ۭu@�=jr"O<,s�H]*%j6�Y�Z�Z1�a��"O,1�r�W�s�� J��F��P"O�]�hR:�zhb2�͚#�:��5"O�=�B��#h����@3��3�"O(�@5�� ����	�0h,�Q"O� � C��9�G��EĔ�b"OVMhr&@��7����X�"O���u���z���Bw�"pT"O�	����Dr�ja�W�-7p��"O�M;��� �h+���n#��1�"OڔA��B�W�zu�E�Q
Df��"O#�'��{K�e�n�H���R�'�2!t%�.5B��KQ�'����'���Ag�LtL��QJ�<�D��'���B��NT�R'A�^t1�'�Έ��fՒW��8��O�2�(�'�XB�@�R1Й;Pǎ/pN�H�'� J�G�*����r�B2).�|��'���Js�L=o��@��4t�����'w$l2���R�h\���t&2�Z�'��H�%Wi�ܴ��J'X<�b	�'�X��(Y9^d"蕒+h�h��'bf@b��[h��b�U�%�N�8�'�6�x�
Y�~ʠ1q���F�.��ȓb��i�a�N>��A�Q&�e�ȓ3���2�)��(p*�/as
��ȓr ��{6�·V|��#F!jA���ȓ|l`d�3��=�����.�Z�ȓ�Q!Eo�?u����둀d[(9��v%�i����*���
7:�Ʉȓ<�����J�,t!uN�3
�݅�w��y���a���e%V�)Ӱl�ȓG��d 3�Ԛo0�u[��[�T*�t��*�@��!�/T�H�y��.�Іȓ=�mj"n�P7 �����\��@�8�`�Y�m��5Q��՝xG(؆�(�6,Q�T�����瓳�0��'��\�v��5�DLx��*c ���!�֕0A�3$
$�)��\��'?�QHₓ�?:b�{�r��M��'��[��!	h�A3AK�e ���'غ5�gQ�$f<}za`PVɼ i�'��P�e�#h� ha�݂LqNx�'N
l��/@!P%�r��x�9��C�<�RJʴS�d�{�&T�aܶ,a��}�<�w�L.-P���,���+Po�<i�E�%�X�͇ [����C�k�<!6"ߑAt|@R@͇�:Q8!�Kh�<)$#
$L{���Z?ek���F�z�<�So�H�h�U��;Y�Xm��&�Q�<���l�P(A+�='�F-��J�<���ӌ��y���U�x�[S�]�<9�j�>Y6Z�jVcڰ��P�<q����"t+b�̀$�B�)&n�I�<i��_ �X���˜�`�y��A�<� ���!�El+^X���Ky��B�"O�q@パf�yBL0U����"O��K2&^�rL,å��̹�3"O��qE�ڹ_�������W�N�"5"O�t�5 Y�D#�0Q��۵�ti�"On���kJ�!n���A��q���"O`��R�˂6i���"%�H�|ɉ�"O�1(aꗫ8��eܧ~��t��"O0ধ�A�"�BBo^2T�y�P"Ob�Ĥ�}�<x��X�`��,�1"Ot���\2���g��m�:��R"OL37k�!��T:�H�.,!P���"O�,�W�`�8!�E�H�j�ч"O��"&Q+R�Љ����a� �5"O��9�O�z��㜙f�r�"O�80C�ە�8at�$JMFx§"O�"ǋ��f��3jE؀�RT"O���V�,��HB6Dպ��V"O��JF   ��     �  Z  e   ++  h6  	A  �I  �U  �`  g  Xm  �s  �y  ;�  �    �  F�  ��  Υ  �  S�  ��  վ  �  ��  h�  ��  ��  1�  ��  ��  �  �  � � 8 �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�	#��$x�R3e 	F�
�Z�Bړjaӕ"O�1RV�GF��УD1�HАa��E�Oԉ�
�]�|5����n��u��'6���½`���!�Ϸ\�~Aۓθ'��I��ܩy>TD�QD��@�0L�
�'#p1��sR��i��̖"n��P�}��)��v���s�_)�y`7Dϛ !���d2��C�(v��S�	/�	r�Q�"|2�M��&U���Y��dy:AD\|�<	#�'�@d�AIڣ��w�<�kc~H"vm&#���硓v�'#Q?u�B.��Z���f��|�  gN:D���RM��C�Ze���H!Z�\h��N,D�li���Mn��!�G�o68�	�)D�@���u\���a�+4�^�˕���M;���>YW�O~�>7�5?�O�eʅʥ,��@��؋�)XP<���t(�X�6f�R��H��9V�N�P,O����+�H�s�&GOCХf˜�
+a}2�>����08B�iZr����F�<��4;�1�L�"\��^D�<IsaA�B�@,�b$�9ۨ��#�D�<�U�\dppR7� SPel�V?9���S	=��H3s�i���6m��<btB�)� ���e�+�h=��M�G��	�'"O \{��G�%��iP��X�7�|%��"O�X@�����i���e�8�"O,\psΛ�L�nE����84% 	��"O��h��A5� ����P��×"Op�qW'՞/�.%�r��V嬰��*lOV�C�̍*x=�a`d -<����;O�=E�t��N��P��hҧf+`e!����y2*�)*�e�fI�[	�T��e���y��,k�,�Q��D+�t�Rp���y�Ȑ(����O���"0���yªA�/����$O*(��`�F��y�!��@�X�r��Tr&�߭�y��Q�.u����! �ö'��yrA�[`͹s`�2d��� �j��yB�>fd$0e��K?X���(��O�#~:�!Q�?��"CO$//b�b\p�<ن���P��a�4��8��KӁUl�<Y&IWX��5�W�/��c� Dl8�lGz�+۟[~��S/��Le�&,ٞ��'���'�>4r��1K�dR���T�
�'}ܹh�k��l\d�eB�?EF�b�m�g�<i��1"VlՋ��Z�=ѐI�ң`�<�ue�9��A��+ Х�"ˌZ�<�V��)�U �K'}�fi�bˀmyr�)ʧh��A����ÂED3B����n��@��;h&��q䐦K���ȓ^��\{�o�%Y���3�I�Qh��ȓ7�.�z��A��^���j@Wz�1��.�����6MY�
��P`ԭ��|�9�-��N�|p��M�Ԃ���.�@���A44���SdgȢ����=PuhW��	]r�:�(��B\l���@��Y�ť�qVLEC�_�b���6�Piӑ�ͣ&�B��a2�0=��n 	Zw ς����Z�}�X���lQ�PRj�:��<��"� ^�zńȓwb�A��FX&hF��Ak��I����W�đ�b��Z���aa�%-tH�ȓk�T�kǨǟS�4xq�G�
_lB�����S��6-��gې���WjH¤ku��.3�!��΢?Ҕ���)�dhp�)��,lazb�$T'=�帀�ضr��(Ǯ��<h!�D�_�lqP��(_H.i���_�DC!�E�r��LtoJp/6�[0,R�+�!�$И�@-��" k��1r()�!���*�8��IN5Zw�́2H�, 6!��J��,�#��Q�G}ԑ���ӞK �1O��ג}2�P��J��`�K����<���$�gY`�S�F�f�����!G�i0!�@�vS�}1����F �̱�a�i�!�Ay�tĉ1Tx�X�r�Ǌ�;�!�D�9'傈@�LC v��ܰ0f	�7�!���>�H�25�=>HH�'��!�$6����WL��D8L�*�$��K�1O�	�����Y�hJ�"dMj�S��I��p�C4D���b&�XR��fc�t�3A>D��I�S`�phF���j���bv�<D�(�7f�,H�v�1`⚅<��@w�:D��:@�"!��� ��'otq�>q���өLz�
�)ߚn ��U�q�C�ɶ|	�pP���R*Q%̒�TR�'�ИDyZ��'d����^�mBf�	1�I�,�hٸ
��~2���2j�q慗�
��b��y
� ��;��B-A;r��7Be>�-�p�����'(�S&\A��a��)�^��D ��^��B�"����%7�����O2�=�gÃ�&�,Ӂшv(r-(�	��y�(�Y���(��g�mJ�ǁ�yb�84��ѳG��4�b�PԮ��0<��d�kH���Eh��U_N�b`E0o�1O���$�&(�v��2�ϧ�z4s��\='�!�$�-n/�y�6����(E�m�!���%���Q�,˦��l
�n�Rn�� ����Ƌ�h�� dZ�M<~����ǪE!�Рw��Ҧ�(>ܫ�V�4[�1�D�a}���OB4�@���x�������0H��8gO�P� (�1}|�lk�@`At��`�4�$/�O�a���[7r1���MAppp�'�F��O6WȤ	3�����S������'@�L1b����cw���:��0Ox5*��Z8p0o�#0H�ZE�'p�'�~��r� �ct��@`NNCrXPxak�<�����. FfЃ4�<����TG��n�$:�$�i���OW>ͨc>�������x"��!�!I�	:��=1@��;(�(�����.f-A,�y��<ə'rZU0H>�'9�M K��r!Ď�eA��x���&O����$LO�=�H��[�	��h^�z��W�U~���$=ꓤ�	O̧ZղhZ���Cf���H�,B���H�I��Mㅨ�$)/��:���~]X��-t�<Ap��5x�j�����"
��j�m�'$ўʧ<h�s'ca% U(�d��m�h�<��K�8Z��� ��T��|����d�<10�W�o(:bŚ�.�H����V�<�G�Е[n<�b���+4`b���LX�<��
g�(z욫����i�W�<)U	��T)�X�/�0�Ub3��P�<���@�5�l�RM�r��R���T�<q�����R�GQ�(}xt���Y�<Yd ̧J���/�\���[g�JW�<�$��SuV�� ��H:�A�hI�<�&K\ {�P�q'�LJ��!v#�D�<��G�V��� p�ٱ<���3�%z�<yV�A�1�J��VJF(=�f� ��^�<)��=,<yp�%����Z�<��^.H�T���9kŎ�#��3T�Hh��;�D`r�,Z�R&�E� C-D���p'*a&��kX�|���D(D��8d��8q(zD Q�6�H��H%D���u �|�Bt�	!&ڨ1U�!D�����)lm��H�C�	r|��Ȅ<D��j#X�J7��� R�.-D�h�GY�)� ��R�_w"J��'D��HD� 3"�+��[s����*D��bÂ��Nj �+r+=r��{�)D��s��� ���w�� �@"D��1�!@]5�w�0����;B�IIô�A���r�`P����F��C�	�0�Ń��\�x����ӏ8H�C䉢1k�$��)�<92ݰ$I f��B�	�� �"Q�Q�����ZIRB�	=@�V\A���2xI�9$� 2 B�	�K�5z���/�h�uSl:�B�I2_��qa��&�b�h�Dևs�B�I�a�N�R��I�6)+�,�,�C�"M^a �#�0S��lVmGs�B�I�!�F���-׿S����bH�(4�ZB�I�=Π��+�5��u�ƨ��zB�)� p�0(�gV�	�c��_<�;0"O:�6��yK5�N�j����"O�������Y��v�R��H�r"O��J����Ŷ�f��a"O �j��nS��#G�L�i��'��'>"�'�b�'|��'���'��Ż�+�{��!�`D5Jp�){s�'���'9B�'�r�'�"�'E�'��4K���K�*�a���|����'���'/��'g��'GB�'�r�'�R8:@��W0�a�bνkH�Is��'�"�'sR�'x�'L��'*��'�b={a����}�!�r/��"�'�r�'z2�'3R�'���'^��'목{W,Фw0�T+!,���B�'���',��'I��'/��'B��'��]�!)�mD�=���#C�){3�'���'��'��',��'K��'�>\H��m�]�d�X�����'��'}��'w��'{�'��'�Ρ�`�Ϫv��A�.y�@1�Q�'Y��'�R�'r��'���'���'W~i���t��ŭ�>3V$�q��'Q��'�2�'.B�'��'\2�'_�8���5rd�����sd&�i��'12�'��'�B�'(��'nR�'?���An5Vv����S.tV�S��'�R�'#��'���'��'"�'����P�u*�ZA�ͷ?er����'!r�'��'9B�'���m�J���OƽA��%B �)��³fQ�)ǝ[y��'��)�3?Q��i���eM	�w�8� �ŉ{��d�m�,��Ēצ�?�g?�޴HvZY	$¡  ����O�;(����t�i��(�	>9�i��O��
.��KK?a1�##flY�F���� �I(�I����'��>}Bi*y�D�+�i@�A�����d�.�M�$/H���O�7=�<�FƃT�$���� ��!�Sߟ8l��<�+O�Oh4E!ud��y"+VL� EIQmH�@P`�	si���y�R ����F��0�ў���������<M�f��H�p�B#g���'3�'�7m\�q�1O��a��6
xТè79�I2��9��'��d�Oj7o���'�\�8���iP��8e�˄v���[�O�@kj΢D������D�G��1�O�O�x��C/����.X�a���	�<�+O���s���!n�(v�A�n�cc���T�r��ش#�Ҥ�'��6�0�i>rRÕ0#�\�Q���"~��A뽟���%�ɪZ�@=yR�7?�VD�_2d�*\"\A��o�c��jQ{��4;Pi�	@�.���Oѻ!Hg�M��͠�iАL�Lm���Go���{�k�\�^5S�'?�ys��Br49en^�i8ѱW'6��t���P
.?� Ћ�DL�QQ�tӥ-^TrEB]�j�֜BՅδ6M�H�bG ]8�%J���,^q�����>�2�@X�~��|�T�%c���X���ux�u��'	|���u��@:�fZ�rTr��?W���F��YP���-D�A�֤Y���61^@���j ��+�b��Q��շA��6�'���'6���O��QG�����["D� ��G& ��?��F��?	I>�'��ӽ��4k�.ؙZT�@�a�14��7�^�U�oZןP�I����?q�������$>p��`JU�
;`��1g�t� �4M6* ������|�K~����;�J��}��E�6��"�iQ2�'���B�'��7�O
�$�O���O������,+/�4�B��<֛��'��	��8�)b��?y����웰q#�$ د6H��#�i
�Zh6��O��O��O@���Oj�+bĸv�
u���">���Z�@+ -���	�������Iޟd�I�vsh�PG䞬GV�Ő R�v}�I�#o״�M���?����?�^?�'�R�1xydѨҏ��ox�#цv��D
�O��D�O�d�O��'&�4�k�ixd}���IyV����@0����e}�|�d�Ov�$�O��$�<���4b1�'`��"O/�,�����8��I��i_2�'���'�'/v�Ũ�ip�'V�8R���id(�*�H'v�ά���jӨ���O"��<��?s��s� �i���sw O6��N7oܹmϟ$�	���ɬG��U��4�?���?���6��%���޵-�4��b)w;��A��i�BZ���	�V.�	�O���|nZ�j�f��E#�����BD V�|6��O�����lZ����ן`���?��	�Y����U�-�r��cy�F+�����O��1)�On�D�<ͧ��mrLm)SmM u��x�Ή�cސ6�N/mj�m��I������?���ğ|�IS�2�ԙ!�t%�g_&-`ܴJ���2��?��zs���'��'��qa���X9�]Ϝ�
��ǅ���'�"�'E\d��rӢ�$�Ov���O����Hl��� �ygk��qe��u�ic�Q���t���?A��?	��>�^X3@o�"�h\Z�A�8m�V�'Z����u����O~�d�OZ��O{��	���ّrM�W���R ��-#�	C������t��g��w.��%$�4XpZ9z�m�0X 8#��M���?Y���?��[?�'��咎'p�T�G�K#��1-S�G�}�'��'�r�'Ar�' B�@�7-N����a������!B��EVo�����IڟH����'h%����\c��ep�
��y{.xa�L0xx��4�?���?����S�v���z۴�?��f�!��2�h��$��k�$[�i��'��R��	:Fr��S˟�����+��H�T� А��!]�dnZџ���֟|��
<`T�Rߴ�?����?q�''�p�p�B�F��U����<���iO2W�X�����8���D�<��� � b���X$3���i�P	�A�i��'��� Br����Op������)�O���3`è#�آ@j��!��K�#n}��'x����'&ɧ���~¨F\Jp}�r㋪'0�q���\�5����M[��?!���:��$BM�j(�$�ݻ6�����$��=ڪm�;��#<E���'f�@!-͑%�:P)PC���y:�dbӌ�D�O`�$�t�A$���Iܟ��3	64����r��`��!WdM�>�U��]��?��?����k!T��z�Zf�ݖgћ��'��X�wN?���Ob��8���|AJ��C�6,P��x�p��[�D��a"�ß��	�ė'��M�"Ӛ�3`�γ.�D�n�N٦O��$�O�O�˓<���F� 7�:}�f��um$1Z�I_��?���?y+O�(7h�|��$�>|_�<H�D�!9�
{�C}}��'�R�|�W�x:$��>���V �~LЀ�MM0*=�u�v}��'\��'��ɨ,m��K|���GK�m�QE�'[~�	p���f����'�'��ɻw@�c��R��&�ȡ3��+�(,v�,���O0�=��2Ӓ���'f����E��i�����:�#�7�O˓f�z\Fx��D\���M0�:��:^��\�1�i2�I� �	ߴC�S��2��$A�E��$�+7^��$j�~ ��Q�0� �S�'�
yyի��5\i��/ۢ=��PlZ
�di��4�?���?	�')v�OBy��!T�G�V�r��!���!��¦ ��4�S�O��+Z1I�L	xe$0�Wj�2C�B:ߴ�?����?�Ƭ��$�O��$��� �S$4.��y�[�*���!R�8�I�K�db���I����O�`3�j&ps��
�Kx��aܴ�?���
͉'���'4ɧ5&�#Ξ��qeI���|Kt��	���:41O����O��Ļ<����1<�r��F�Пr�,�[D�!�%�xR�'��|BP����-�7<J���(T�����s�f��yr�'���'��I�ҥ��O�h�!�O�?L �B��,͒�ӯO��D�O�O�˓G�֠�'�� �'��3G�F��Q�ȹ1�O���O>��<�B�/��O��y�`ϸ�x w;(L�B��y���2��<)�"�o�M�4��&K�n[$@�Q�Hpހl�џ,��DyBM;k�����D4��F4#N�x�F��.�xɫ��H�IQyҎT>�O��K:%�%(��3�R��]#�6��<a��^!:�͠~2���Y�Hh×/H�0�i�#�
6,��B�}�b�I@�Ex��ĩ^�	V`T��(���"U��Mk��{����'�r�'���1�d�O�,��ɿ����Q�#h�r���u��4�S�O2��z�ٲ���t:&ə�n�h7m�O4���O��Y#-�m��?	�'V0`i%��Q_&i�0�G�t��X�}Bi+Ř'��'��U�3Q*�*  �r��m�G¨).6�O�=	�N�~��?J>�1��3fI�x3�5�e�욬�'�x+�y��'���'��I#,�bH�E�u� 1���%�
�4·��'G��|bY����F��x.DhH�%B1C�x��K�Fr2c�t�I���Fy��(q�Ӊ$�*8�ElS.~��lRf��@��O���(���<aTN�b}���/c"~�W�C9w���&����$�O,�D�OnʓTXA�����ر(�V�� ĕ�p]�����\�_ͪ6��O����<a.O($�3�?�D@l2 �6e�5iB��/΄ml۟���py�V�%�0����� lJ�`[�!`�9�E�g����A��i�'�I�j�g~��M����w�l1��߉lzt�Kc+�����'���s�}���O2�O���J��h ��q�R���9})vUo�\yr��!Sy�O�x�i��F��Ȉ1D��I�;�M˱)�|ݛ&�'}��'���;��O�и��-d}2��f܆��IB���l��|�<1��X(�M�p"(�Pܘ2Ó�*n%I�i7��'W�h�7#�8O��$�O��ƉD2���M�
[PP�-:b\��>�%*@�?i���?���?��0��ӄf99�Z)H/E�R�BMQR�i�� ���O6���OOk엑+/��0�A��w���#�LP��ɢ)�r�'� �I����	_y� p��t��,|,l:qI�'P�����]����?q��������2wa�#��2��!��L��-�����D�O����O �-d0P3���bb�,�t%Z�[�ڐ\�p��П\&�t�'��౬Oj�	  ި<L����.
B\�d�	����PyRbܸp�
�e�
�	��viōI�ౣĢ���Q�Iu�	{yr�����'���&�"
<V��W��8t�<D��4�?������x��h'>��	�?�ʖ��x�T��R"z21R�������N����x��l
����h�:X&�O#�괉ܴ�?Y��M�z�V�iD�V>�����$�8�:(�0�Ƃ���#GZ��6S�4���&�S�'}h�AF �f�@����m��>�Ԛ�4�?I��?���>��'�bAΥ!��=S��XҔ�9u��*n� 7�A�O~�"|j�z�� �Z�(MO�h�BlG.;�T�ַi���'Y�iW�;�O��D�O|�IlT�K�˅0<Uzi���K�w��b��d�1��ݟ��I��T)V˗�q���af֗c_|���*�M��50�D�x��'�r�|Zc$LP��%ڂX�Av�£2���P�O̕J����O��$�O�������7/ƅ��O�2pR]��e�*�'fR�'t�'g�IM]��4k	󘱢V/��.冥�&�Iӟ���ϟT�'�(b�j>�b�!��$UYF��L
�1%D�>���?QI>�,O��˵Z��k� �f5x�UG��bd�>���?�����D/1`��&>�.9��t)���!�n�§�ѧ�@Yl���%���'Ӷ�э}b/��kb��K�k��?���˴�V��M���?9(O��dLu�������k��c���a�����FQTyK<�)Ol@1��~��X��u��Y��#K
��'׆t�pӌ��O���O��EN���A9nnH�F�[.���n�Iy�fԘ�O��R53�AC�"(�{���Z@\�d�i�$ԑ��`�F���O<��蟮$�p�I�Ȍ�ì�7,B^�I4��Fziy�4kDPGx��)�Od��K�[�~\Hvœ�5v`���%�Ʀ��ϟ`�	�,��$�H<����?���BK��k��<C���'��90��M�gK1Ol���Ov��Q�NP	��IE 2]�XH�<���l�ꟸ�@J��ē�?y���?))Ok�	4�yN�n�|�a"�>�>#1O����O���<��Hع-Fu�eOG�9����Ơ99^���x��'2�'�����H�I?_�r����7ut�a׊�yW$=�f�!�	ϟ�������'ۜ��t{>h���*-�8j�4'I
�B��>����?�����D�O����(C,�ӷ	�	AV:mྈp�G�57�v든?A���?�.Oj��TW� Er`�c�N%���pǡ�1	�BA�4�?�K>�.O� ��d�� 7����'�����F4����'_RS�tIq K*�ħ�?I��(7���	�F|`���	U�V|�=���xb�'�"cҩ�O��3����Dp�� ��	)86M�<	тÄs�����~����� ��l�ЏZ?A�]�3�I��x�Db�����OQ1-�O��O��hp�@��|0�\@����f|�<�C�iD�Dxcf�����O���$���IrJ�,���W���p��!��C�&8�ߴ,_Z�B����S�O��+On��C��Q"���[�x,�6-�O`��O�)��R��?)�'2\$��N�1M�59��H�
VL�ܴ��^�
q�t����'���'���ׇc����	/З�r����'�@,kl=�	��@'��X:x
T)&,:	p�8"�۳H��:������OH��&��ũp�L@��� N�A ϱe:�Z�'D�ޟ��Ib��ޟ��I�|4p�"s��I��}�O��S��9��,����,������'�
�BP�t>q��;<d�����\�F�c��>���?�L>����?�QK�<���R�ɦ��EΝ
�Ӣo�/��	��	��|�'��p���#��D�S.�цGSR�c��b��n���d&�x�����K2��ܥO�8���DG��[��H�e��9�iA��'*剌F9�eJO|j��
���#�0����F[VQŤ��
̉'�2�'c6t�e�'Rɧ�ɑ�L*|Pt+��b?Ƥ�q�\�Ǜ�Y�<��;�Msq\?1���?Q��OZ�:ǣ��Rb#��o�
�"Q�i���'qP}���'!ɧ�O�Q��ͼE��l����{��]"�4ԉ���i�r�'��O�O,�$��� h���͑Y�ѓ��V��%�z����b��O�O>E�Imnl��	�0(���P����ش�?i���?IT�4~�'6��'��d�+M��J��L�G��$C��T|�6�|�� ������O��Jr�F1* �6,1��"6)[�^���mZ��������?����{'۰{�بY��D�H2��n}2�?�BX�x�	ߟ�Iay�`RrY���G�[84�f�y�n�YJ(�d�OZ�$6�D�OX��W�O�.5� �H�Q�MU�9K0�&��Ohʓ�?���?�)O��Q@���|r!�KD: }C��O�e�mӄL}r�'Ҟ|b�'���;�D�3>��r�a�&)�����ӽ�Iʟ��	�X�'��(���5�Iρ2&�ܠ�lP/^��� W�W���oΟL&���IΟ�f˟�O,|��K���i�Ö�0�pJTj;}���a��G�>C�	� �zӮ�}��z�\�۷B�1|�����Z!�,��t�����P��vx``�� +��1�b�ӑDC<kt�������$!�M�t�øPk0�H[?솑���՛H@b��5��P|~az�����m(G�H'e��m��`�1����ځ|(�$���|$��2���3�Ɉ� R5N^��!A�HS�ٚ��T,�H���"Gb|C���2'���ybb[�3!,�d�O����O����<JL�6@�%�
)�a(��Gm�t�P���Ym�a)a�iVd�#i͝)x1��7͜ =�$��}��!�uș>���١o�?�a�����k�@����*�����f�mj�1ODx�ǈN�q.��O�5qf�"��O��h�P�i>�E{2l.I�"}2�A�u����5�(�yR�N�'���a�(N�"��D,�����c���$�'��)� Ph�@��/|p��H�b�Dy2A��Re���G�O�$�O���3��?��OL�]�5%��B�<z�J��1��	Pd��=m?�8S7�ǵ}������|џ�q�+\4f⸙���@�y�f��9��%lA��tx�^7Pd��G�k�0B�>��P��(j(A���6�0*���f&m�r��I��T���
���[��1�	���B�I�@#�� Ѥ��8$��Q񂖒2�c�8��O�ʓ~L�TU���I!������hM���Sm�7p���ڟ@�b�۟P���|
MW�xG��Po]n��K�j��	���1� ~��4ba �@MR=����!�&""N��Di�� ��l)�S,�/��L�B唿hN�+EM;��H���ٟ�''�&eQ6QR}87�dG�	�y�'���U#Z�}R�PW؅Ua����'BF7M�,P�RQɦK��R�(ԫM ��$�<���9��V�'��\>1��'��0�-��*MV���Ӡd�9+D*F��h�	9e��K�&�q��Б�+'�I:g��=Ph.=�O�x{&���y�9@��ߥq'�PAN�,[C��|Ð`���Y�`�id��90ɚU�ט?9��@��V%�)��^�,HV�Rp�$}$��?���䧇�h�H	�����
�����p�҈y��'��yBb�2tܹ3�$�� ��RBO*�0<Y�	h��1�W�HF��H��m�$�>���4�?���?�1�Šn�$���?����?���Wrڴ����;E]cL�7+<��V��0$q��Iz`�@�G�k�g�I�B��c�˰%������%5M��w-ª2�r�I#3��yh���|��Ҳ~��!;��U7Y6@X��=xb�'x�%C�u��,O��$�.=mv�FA'Sb�3�N�[�^C�ɵk���Fb�����1� ����G葞��h�'� ����&2Lq�Ѡ�/y؁#2#����i��'1b�'#b'l���	ϟͧ,�ʈ�t�]9(xj8����|p�GăMH�Ё�GV���dZ�s�&�#b\�M:Ԥgi�? ���el! V��ge���p=�dHĳ��t�F�ci�4t�K�7�6a�I���%�t������?�Q�+s�f�Rl�YV�j�e�<���R��t�tk�i�6L�v�
d�c���'��IW����4�?y�����1b�څ8��rg�M)��"��?�P�*�?����dG��1�.�� @���ϓr����$n�(X�n�#���E6fq�㉬cÈ5�īD,v��}�;OX�2�.�Q����O�	D>Y��'1@Œ�7�v�>���q��r�ŹsT �(�<a��?����K;W���"O	�xt��ږ�ΒX!�D�ĦI#�MDp0x��Sa C7rU�P�����'5���5��>Q�����(���䅟7����%�9�$C�^�.�D���O"����Ϛ�
%���ȇ:^�,��|�/�ҭ���te(�Shpk�h�h��>���;!7�aQ�[2,7ȡ��	�
JA~�/�t����f��i �>d��ݟ�	���IO��@�l��#�������
�U�<����<a�_�&������y�B��2�@N��*���!�:��S�!h�K���a?�+��Rş�	������H4E��Ο�Iԟ�#\wX*U���.(�ؘ�wm]�AX� d5�\�!n�OXY���)Y1��'LF8�Q�H�D��F�X�JY����ɋ"Ј|��K�~�$d��O����)O��@���B(�1p��++��[��榵.OZQY&����?9���?��bèWx�kGL�=�E� ���Ɠh3 ��̅=,�x�k��F�(㤙�'��"=A�'�?�(O@�O����s�mWVlKѣW��RHI�I�O����OZ���̺���?��O�<�0H�[}���v����~U�� F?��p�F 5]��l	��'��@DA�b&�l�4�
y�Ը�ЧOrx�5`�x�Z��'y�5 R���?�REgR����gg	��?)��䓖?���'�.Iz�c7l��b��!����'�����C�xB��[���<ʕh�y�y�z�Ĳ<I�@ɛV�'�r�Ɂxd����У�U� �!~�B�'��S�'}�:��l���'���p���J�V6M��s�����)B8Cn-�F �.��xR
�?8��9�v�^�X�c+Ыw�2\�gV.;0� �g�;y�p��dO�\g�n� �'��`B�LS�	���C&�	s���2�'��'4�O>����Z�8��qmK/-lt�#S3�XZ�4W�F�Kp̀d8M�2��n�܌���G��1n�jyX>�c�����k�ΖL=�@֥�]�����h�	E(���P ~lb@���M�(��ʧ�.Њl�PT��#a��0h�n8�O��D��q�J]Бgٍa�Zunډi��������F��uI�ɉ�@ "b H���>�3�A�8�� ��'��
�6�q��( "�{�/���l�<1����<�c���\���FG�ea�c�0��3�4}\���|���'I�xkb�N'dp`��EV�6m�O���O�qI��C?C����O����O�� ���G��D��}���ʃ-�~J�' l�*�/���q	�)/�b>�OT!���M+�;c��� �!!
:�2�١����R�ޒ9q��'�t�B@B�dMv��F��f`�E���w��Uoӟ��r��ş�>˓�?	�EI�m��@"p)Oa�< ��O���x��՞=�Na��@�0��-���\���$^q�'#t`
��'�剝y��Yǂ@�$g���!'L����*E�EI��	���I՟�Q_w��'�B�Y3$��q��d�>7��[�
��*VT9u-ݤv"T|�o&1��6M���F�7�I2E�
��H��u+`��Oc�T��m@��X�hHS�6_0�7&<N�� "����'ɀ�և�����p*]���$٧�?��E��'�2�'��O����n�&���74J�x��9Oʣ=E���� �H�$oM�S�|Eib�/��'ɂ6��䦅�'�fi#�hӨ���O�Ep���)]w� �1��x���h�"�Ol�DZ�+���d�O2�S�jre�.L�\aC�^Ry��H�
I'pn(²J@�H���ės�xP��'q����Lğ$��H�f��A�z}�MT�&fr���
���kCl��9�����ɫ���\ͦ��O0IȁiN�� �ɴ"�m}N�J�$�OV����*m��ٗ=����R�!�$զ�A&
�a6@00)߭Vk5q���؟ �'Kzd�t�{�����O�ʧ\n��q������_�bK|�%�Чo3jl��?���I�i'����H��|+����j'��w�$�]O�E�C��]�j�A���	?b�rA����ʤ��EE-|��~�
��x�Q�hU*+D���"��Q�d��T��'A��'��V��J��?�uH�	Y,_�\M��$�Ot��$�,>��d�u�U**x��v��ax��4ғJ���C&N8|ݰ�i���V�p�:��?��!D�9�Q
�VF�9��F9�!�ȓ[�p�X�X�ɺG�ٻE��Յ������"�*�b����6>� Q��pT�d���P1=n��ps�.��ф�X}L���
C�q�^�k�k�s�8��
��h�¯L=��`[�Oй?��5���0$#�陸#	4U���0��!���ȉb��F|6{�d�#�'�4i��-I��U��̛)�p%�	�'���BL������F��.l� eP	�'���ʓb\�.9���,�"qة9	�'�FH3��I����*��P�r�'&�)��RS�$	�M�4,܈��'1< Qg摻!�~�Z���.Z�E��'�(x0�.*r����DАW��iA�'p4ɀ�D�k��Q+��^/~��{�'tL��ՠ==nސ9��x��Ih�'?:��A7^�<�'�ڀ#�Z��'�T�K�d8�X�%#������'V~+e-A��dq1��)!p�"�'���SIP����îB�A���
�'$�lS� �"0CF˗1���j
�',p�T$R%{Z����	�#���	�'�M��{��X� N�f���	�'7�d؀�X�����%�%��N�<�� �qg@p�ǨC�AG�	HW%I�<��F	��y��VyJ�'�[�<9�%�)V�6a ��I��g-�B�<)w�Є}@��s)�/@?P�:v��}�<C
�
�J=Ⳏ��0N$eZ#�A�<QCA2ONx��,�dk$`S��R�<a!�]~����
Q����Vb�t�I�q��Y�I N8�����~R�dîU����q�=Qܽ�������X�g�HX��yw%9��l�l����I����*,��r��<@��hD�0)�8��s�TcU����i��b�.^<��S�C$}u���7��"�	�� ^@����Y>��5�=[xi�d�WNex���a�F�o-��lZ9^��x��s�L�c��^��)�1��a/Z!��i̖�I��ܦ�8CnȫH��1���i=�`�$)O�4z���#L�;���;�6
��N�3v��hx��:�3�HtDRf��D��I��K�T��ԀBkYt̓3��G�T�E�.�2!�_��e�#f�V���3��S�M̠@ڑ��݂L����mw�u��j":uCQ˷)y�;��I7H*6�"���� �)wI�>wWl�&-���,�d��u�E£L�}{�\�Ű�x��y�'I^)���ō>��4@���0��`��'�n���ԟ!Kd�L�!�0XI�B��l����8x���r���1�<K�p������
	� G�£䘧�'&���4���8\����"��b�`ԦO�����UKE����,N�|Fq��D��`i���G\��bR/_�]������I�f{�#|��d�v�v��5,���1���_�hC��a�\�VE��^�l�����jG����� ��iL�D��+D�(u����e :ٓ�HR:�1O:ؑ�@"��TT9�_���2�B�	Eĺ����y�©�v �j����cs�
ٕ'Q4r���h�t�U
�!N�x@��H#��H�R���?�(R�����#����y5&^	nj�)Ycb��Q����i/��)�E�%����3&�]�=I�bT�<Q�'#����æ�{#"G.SsX�����r��(�t�c?���ȵ�&���L�C���+�I�'��:a�J6>[r�����^��T����w(e�!����oNY�.���hB�y� �
f:�{��_�3��pE$z��b��S�W<�x��4�4I���x}V��$P�z��J��b�R�d��} �5�%�Y�d��h 4,�X=����L�^c�Kх���C�$��z��|���	��D�Ppm�(
����K��9BJD}������9L�L��a��:CQ� ����?
��<�����
��p��^(�1��<�ˋ/���S"U�dIy��}~B�\bj0��t �1��x��i�����'���Û�R}|a��D�fij���H/y��+��6 NN�h���_$�C#0O���b�E�}:��Q� ڴi�(�xq��N���ۡ/�.�"�W^�T�֪�]���Pi�$TT¼y�'��@Pcåx���7��'~A���l���B4ٛD2��ka
N���B:騜mZ�]mlA�ش
*�O(/��	,O*��J ~!8�J"/@m�rT��Nn����\4���S<[�84	B��f�r���L��\^q��LҌy��{� �C��`0��X��͙�O�lvM�Ag��( e�<"t�<�g�x2��H�țT�A%:y��C����ē
�r5:֋P3�&��� 9���+V�C}��0�h�O�Y�:j�y�GϜ�@\TmRaf��lQ��񥮊8t��M%<O��ଜ �x�I@� 55�c��	�o�	��'8���i[��䤬<�;]5��b�=O�P0���� D̋ ~P`��@��b��'� ��� l�=��U�%��(�U�WE��"±��X����$1Y�N߻��'�=�獗,���I1M�%<�D�:��ʿ*�"=QU�[�2x䥚"��1���xG�<�EL�3e��]U�ۋ]}�<�j4Z$9R���u�	��qeD�/�v���$؊=Ph�D��y��`��NX�de
�'����/�M���S,M��H�L~"��1v{�X��yӔ7��/��1����p��4PgbF�]���-(�î�S���X��7_ў�(�-P]�.|[���tx�����йr��'�p�硇�S��6M�<A�O��,f���G���k����2�*D��`h�->�����ڰ3���;,���*FG��D6�}��o�_�lq��LL?���6\#��a�+�L���́:$�M��œ�^,����7W����$�=�`|�ࠑ7-|xB�ݵf���1	�= jfY[�K[�5�p���>b�|��b��%��b�� �j��e~�uYwB)i��!2�w�T�cjZ�%��K�+"h�xL�I�er�I�#(W8�LT�gbJ�E2HH�'	W`�P@��&�9Q����Wcq��ɿ*�2�!�	�8z�21X�@�>)��C� r�<3F�}8�ˍ�"^
�20g��Q�e� �/G��K<�~��)Ѩ@��d�c^/����@�k��g8\O�<3�>�4'/"Kj�Y��l��t�|([�Hk��b��Q��9��	
1�D�.DZ��$��J9�!��(�pрiE|X+8ޔ�sW!WdTDz.
�y�A��}إ�H�D����D�2�M#��D	'	$VmB�i��c���20QJ���d�͊G"�		��%i�ϵ;=�̌8��L�Xy�Ĳ<��&Y3H����'*� `��
�d�;#@D�E1�@�̭�O��fBU¨O��pC��!��!�l�5��W1O�@�R�XB �O�+���%��OM�m�N�EƎiY�I�f��̶֬`D��I�'����r�\�i5(�|R�i ��z̤<"C�վ2�O��'����,:L�$��M�|��*��5&z̊`a['*�Q���@�q�ɖԤ���56.~3 ��'�
h8������Cph|s�����y"g�v��'�*xC�O�A�PLc��Y�"�¸UvX q�(��H�d��k�T���.K���	����xVC��V���[���K��E)Hz=���MQr՘��9[NL�xc_=�V5�����pf
ճX{Z�밢Ɇh9jͥO�O���Ul�^1��h'<���'Ϥ��qj҅����'�!<�Ҍ��O)��'���O��S�<�Ls�t0Jܶ\��}�&i7c��x����g�0�C�m>K�	��D�$:&�@�7#�C���h!��@�T<huf�e����O�u�q�
vݺ!Ҷ����"�I��I�N��CŦKZV<�B�wi<�i������t�\���DZ��*8�XJP`	�F'�O^\���կE"�l��&���Z!1O^�X J���Bq��*I�.U�N>��b���E�څ� �j��M��!V�_����퉙I�>Ŭ1OG��#NN�U�D��h@/O�6X�tXR`�[I>������&�~��9�X���&�!Z�.�ka'����O��"$/���`��)� ����OǱo�����pq��3��'xt�"A��^��I�-��'�����i?���[;�4�� خ�:!�PC��<��I^����'��}i-Ov���ɧZV�I�����v�ԙ|� h���B 8YR��)��@��s�/�HN�	�L�y
�Y����mF�a���D�`Kd�Fx�>aM�@Ʉ0r�XI����$x�4QL�'�'^����w?|���O�(b�=�g��C0|�����hO1���O�/_2>	����~M\����47��m8�AԂ��ѧ�T�����#vҢ͓�6�:VO��<�&-ȴ�ըE͔'��'�J����HAv���(Î#�'R��J��@���"��ހ��'+d(��P+|�����	�R� O>��On��`�I�P���Š/P���'�f(�@'�HXx�
�
�n�ۉ�Ė=lJ����%���Ub�a�l���l����'zў��<\���iqF�Y�HL��]
c�������V���$ӛTF��ϻ� =�˖�:mVɡ��Ζ&�Jd��3�y�^�(�S�L���RH�g"�9flS$M�h,&a�
a�ƴP�����N�1�!��:� ��o�����	'�~�sb���LE` ��P�u��O6c��%�ߩ�JA94i�A�92G�'8�%[_y���@g�Ϟ /�lb�hӒ�-kL��Bc�߾@��m`�n}B'_���O�6��/�N�Z�֭[Z5YE�R4|���~0n��֢�
2��� �7�ў���
�!����"Ȕ1sr�A[���, ���'�����'/�d�|2K|��ƌ7*�T�R��20�q��-לX��y�fFU �p<A�eF���M-�T(�Đn�.A�$ɡG�R�O��� E���Q��Ti��.�2��e��A���0AJP�hўL�[�pji�d �h�L��'j�DTE�j<	�$Y�`7������D]����@̓ݤ���� nɒ�rkO�?����UA�"ȜdV��yGݲoh��$�,����%_����
�j^��ĺ�,�'y 	��F�2��`��� �J(�����l�4,q�!�8(����'��˄F-n���;E�8<g��Qf���4��bܞs���R����D�����u��=V@]�ᖍ�����Ơ|�1��"D���	 Stj��ߟ�F{ʟ����Cf���E�ԏ	 d�I҂x��)�c�ĹS�0��$��qrF	?+�Μ���פA��q�t&_�aa�pq��Z�ڄ�BP���'څ�F��
���Q/W�*�I�P	�đa8��Jw���[/^��4i"?��� /7^�a�$ja|�:6�wy�x�u$����톜"(Z�7��7����]n�+���:s�x����KJ�8a MJK�f���T�/I����l�s̓�hO�i�?~����Am���nԀmĆ���Oۭ?�ay2�͈A[���Fl�x1�ɥFϺ��@�:.�r��6�S�'nIr�h@��"�]zk�t���h6�Y�|B#=��(QA.���K��p5��P^}b��ZuĔ���'L���U?���Z�>�j�W��y����;�P��a�'�Ĉ�*׎)�Z���`�Yq���ߴX�T��5MJ+r~-x$#�2:{��'-�4��� ��l����Gi�(AE@�$��d/vll9H7L
J�2$�D07�ў��g�d�F���yaH@����4S��S��a���h�<E�1t�h4���K \��R�C$^�@0B�����jB	WJ�@�)�d�P�G��`��r��J
$�@�i�S�Ox�d��i_�t�$�#lN%7 �"�}RA�- 0�����==҄P�Ğ���r�����Z�\#��.��|=�����Oڮ�u	�)W����M��
ڸ꓌��a��9��`�:"c�	�����~Ix�B�����!�J~��j�2d0V��`K��G�x� �nFv�Ć g��8Eͬ,qZ�[��*U��O\�c�N�"j����%U#��a���^��s���i�[���1Q�Z�8Z�.P��`�h�=|��3U�J�G�Z#=�;�����a�-Zu+C1�����96��@�4�Ң72U����!l}2�����6[�3d� o����9X�e0UGW�-6�8b�"?I��խ^r��r�� _�,0Ø�<)�-�oW��ʧ���[d&�	I���q
ڴ^8R=CR�H�@,k#@��M��W�'�J�0�%��9$�$��1�QA�v����	+N���	�[��=b�A�^h�����'��g�'l~���T�2�����(&����.QjaHA!�j�l�vi������pXE�
�W@��-D��6�y��i+(Q���H8�4:����'��;����&�A�Yp��)ƆD�l��l�'��;.r�bY�s�2̀'�_��鞬M�L�@�!M{F�2���c�ўT�#�P�Re@þQ2��Oo����m�.�nɳSk��X����J^�Q����?ɅML��(�׊�vlPàC� wEf�z#D����OU.����8X.�t[�# D��Kwmέ'�^H�C�\3�D��>D��s���	e���f҆4r�\�F8D�lC��>[1�8!!��(2Pt4�D6D��� À+a�v���UIZh`�c'D� !ע�2H�\X#��1X����$D�� P��$^>�trɗ��l��"OȘ���X���
O�Ղ�RE"O�(r�`�B̉1"�.���r�"O�0���I?h��ж�L h� 䠶"O6��7l�Cn�i@Ժ ����"O"`��R�]� �jA���&x��"O��r��0�>��^��(��!"O� �'2�\�l�F���"Oơ��@B�A�	"�I8Xq
u"Od�P�ڤ���1tIW.	D�Zq"Ol��L�U�\іHY�} .<��"O,�w��;VXpT
D���`J"OQ�q	f�=�Is� �;$"O4ă�O�`�8�+� � pqT"O8�W-DPӸ| �悰+����d"Op���.pK�����\�(�� ��"OP�a��SL����'۴8߮1IT"O�U����3�|����� �h((P"Ol@[���P�d���˯Y�X��"OZ��J�H��Y�0!?c�l�B�"O�)b+(]��R�ɵ
q�݀"Odh���K:�Ja��D[~a�"OH�Zq$ �m13g�NH�;F"O����J0�����T�!9��""O��@�T�/$����@"?ª�q"O�ܱ��ܚ �n�+a J�5a�%�"O�P�ԯE��x�9q/�\�ڀ�`"O���4�6ppu����G��s�"Od����B�F�M��B�d�Ի�"O�<��HҸ&�)�(C7p]��"Oz����݇MF@��C$�P�$"O��V�:���R�X;��0;"O�\8�d�*'��Bp�b�q:�"O�2҄o���0�)T�\�8��%"Oh���,Jl!�`�ɠ�b�S�"Oԑ�nܿ{	.�H�H�$;��g"O��b���>g�>��%�ʇ'V(��"Oz�ȓ�V�w��xx ������"O�aW!��JX���h��e!�تe"O8��Պ�(!^	J����-|�"On����%1�&ܨ�Z�h���"O��V��x��Hz����f"O`Mj�'ĳuC&-���6��u"O$|uͅ4��ȱ��\o][�"O��K�Q�m�&U4
FY��"Oy� ��u׌	�P�D3���"O�ٙ��H�4�� w(D�q�"O�X�h��t�(�B��Њh���S�"O�p��
O�=R�q�A���z "Ot��K�4�*\�Uė�
La�"O��$X{n戀�K9,���p"O~�Kq��0�
��f�7�<�"O��9���>� ��F=k�tp"O�!`�ލZr�ӆ�NX� �"O�-sA���s谰{��>t4�6"O��r��Z�jA `+&��>fD�@�"O���$N�|��8�E�O3K����b"OZ!q���!v��L)����(kb<#�"O~y8�)�1D�H�ۣA?N8�-��"O���C�ͅ X9h�oށ%-�!s�"Oؔ�g�I�d�~LH��[ 3t�	a"O(�i�o�5B ���*z*F��"O��A"�;���b���:t"��D"O d6��	K�h$����3d��A�"O� ��1	����e��+�E���Ã"OBMR���kLɑ+V�8�̪ "O*��b鄭Zh�xU�O�F��%H%"O�� �G�;!������R<)�P"OʀB��@�=	A�Q]X��R"Oґ��.׎G���`�Q2q0�c"OPITK�9��#�)Gd�"O���Q(A�-/����C׭xTD��"OR���5oa4�%� D<e�U�z���'i|�(&� j����IV)n�0q�	�'�H�A��I8�� "1`�j��+Oأ=E���L8�%9����L}�H+�y�7=�x��R.!��(��:�y�S)R�24 �/z��* ����y�) ~L�a�R��J�$�d��y�#�4�
�:�.�����a��y҅��|4����l� |�&)��ɀ#�y�L?r�� ���%����J��yBn���f�H�|a������y�ƺ4U��)��zfu�5���y��P�wU2��B �(=z������y�(��'��2K�>^���x��٭�yԉs����nأc�l|j���'�y�Q}��Q����fWlm��S��y��A� ��-�
_�\kea���y��T:u�$|YV��(`}X��R��y"i�`�H��J�<(���y"$��0k���%�U�U��xa�J�#�y��
a�٫�S�����wGE!�y�>@m�a��CE$��ƥ;�y�	�^d�*��l�6�Լ�yb�҅;�U�h�^��Di�.�0�y�Z::�æ��c����N�3�y"�� }���Ip���L��h��E��y���.q��" �߫x.�8�mƕ�y�d��z���£��=U�<U8���yB�C��H#�+D�M���Æ��y����pq���Kb�M{�*���ybJ>W��(�Wc�I�Z�I��Υ�y��U1VF(�H����L�����y��9S��X���>_���!7���y��Ě(������S�R�ԕa�HK��yB�
iA��#w��O�yB%���y�DY-"��KF��N�z��T�y���>FR�X0�ܪK~M���K0�y2IՏ5_ؘ�jE)<�BՀR'Ȼ�yB���p5h�HO);�����eW?�y�:L2��XE����@��yr�7!;Z�Ah\:��\����=ыy⦁�:��	1$P�K��U��n���y��J}2�	�Ń��X阜�a ҿ�yr�]�Q�n�PV��K��t
���y��'S�@M��Z�@����viÃ�ya������C�<2��|,���x�	�6�ǉ��hA;�L!��2nB��U��7�x0�f�^=!�ĕ�è�1!슉b���� ��t0�
O�*C)��4�>�(�E�;7���r"O�C�A���E����xI�"O������2\��5�͓�2׶�"O��A�OT�d���"���e�r�r�"OX��J��|��dbӯ�����"O5��!�� ��9F�����"O�81-�b��zeI.n_�	S�"O� J���Ö_� ��e�@j!D�p�"O<�cM���JH���"v"O�kWNL�4�R<�Fx5f���"O����N�3��40q_�$SąkT"O���gޖ	���R�e�1e<0�r"O]��@�<��ҤU4~ph@"O �tG�$8���ݲ6u^�$"O.�t�]�)Z�u+Ο�jr���!"O�0r�g�z�(vJQ8=�Μ��"O���QÀi��衠��*yP�e�`�	���<1T���q���U$|�\��Fa�<�5"V�F�)��MT�Oqu���D��x�E׎u.�@��:*�p=#G��Q!�$��%��%h�lR1@�@��!�ãQ!�ĉ�QΠ�e�ؙO����R�*!�̈́9𦼘��ܻ��(�.�'#�ڌ�ē>0"�r��ۑs�L�re�3dY����~,����
����<;#��[�t���p��3g�	>��1��F�D��ȓm<tl���1|���+���5Y�zU��{ 8�:����)�C�
�*,�e��q���q����ȅ���
Tm���ȓ�|���
�M�c7)��b����oHi`���Z�С�؀�x��sQ>��^�%nV�h�@	�Cj��ȓP6�)Fz���Gc�$$��ȓ[lR �fB�%E�ej��Nn$����q���;�E���^'���AO3
��D�{����lH���"O4��������R;16�"O
}���ϩ812A��`�~!����"O:)��^ ��X:W/�?
(!�'jL��r焥L�&5!4�0�(�'���0i�+�r�Psnˍ{�r���'(����֬-Sl%�
pk�=	�'�����ߜ��� ���r>���'�d����~��Ka��=�ٺ
�'\�t�F��,�j���߼.�ĹO>Y���Iשp�L��*�=�`%���YS�!��j���2b�F|�lP�	�*Mx�T��(�̰*���\�*�Y�F�Z��E�"OR� �"\�`����w�Ա�j$��"O8�z#&F�}>4������nӺ��4"O�� 4��6^��P��X�j[
�"�"On�#fS�/�X��J�3-<N9����D�O���rRhY#���Ŧߪ���'8��Q��'>�x@�!@�(�"OF$�d�S�`��F��_(p��"O��ɓD�Fu�I�7��%}����"OF�)c�	xlق��ċa���f"O|)K��B���Td�D�\��wO��DQQ�]����9��2�m-!��_%��� ��q��|�!�dĵki~=��M�I�4���J#�!�d@,&�ʒ��k���fP)�!�2bm�[��B1}(�IXv�S�c*!�$��W��5�G\Lt��%V?x!�dN�LyN<�Eґ 9���E5(!�d���I�&�Q!VV�Ly���4<!�\�(�˔f0lנ�S@b��3 !�D�9!��Q��b���P���?c�!��,^� �⦁
�>"�B�j�!��?^�nي�o�-<�0���åJ�!�$J'1���@�%K#x�\X8A��/5�!�� L����:K@��k`�^ũ7"O�@��E��x�v
������"O҄+!,�N�Y%�W��L��"OPh�(��t�xE(��@��ఐ"O���J�5�i�Ӡ�y����1"O��qv�Ʋ[ ����� 8>(�Q"O���u��9KJt	r  �r6��"O�STdJ#rBL�0��p�|�"OPx�0��,9���n� 1�ܴ��"Ot�P�ѥt*~��A(ˉ$�VQ�"O�=A�nQ%@lx�+��L+2�j)�%"Ox\�B 
)u��r5�`����"O��XW�SR��a�"�>���"O�
�j=-ߜ�{T`�hR�W"O�t���[W&)��Ȕ�P,H��"O��*5��>~��� ��9��P"O���T��{yb�!q��&t�\�""Od�����v�Rm:�揕��v}!�$Y��}���
�D^� ��ڕ q!�D-Fr(Pj�>B��x��N�A�!�d��pE�Ɯ�N+�(@Q�G�?�!�Ğ�6{>X�5�O!`P���3�!�Z�VEX a�;�h$�B��!�!�d�6;j�j�Y1����#���\�!�O�'!>�1@��� $�t%V'RY!򤃤s��	�#��ax�+��M�VF!��Eж!�#K�;�e��
S�!�T�|��({��͋=8�Dc�*܇v|!�dNX� [����r��3�H�XH!�ă�c�u3*�7<kLYر�i�!�D ,Ƹa*-ŭxi"��S�	{�!�W���bR�R�iV,�(��
(x!��ƑB;�a sL���|񡊋�@!��T*��}80�J�x��K^�O!����%CC4���wKL[!򤝱cR�ڦ�;8�n���˃I!�M	���i�>|� ӕdȖ$!�B�lD��N������2!��Q�/:�!bP?�@\�����E!�$ο|���"��[�(^6�Ja\�!򤁶c���2%�֤�zE G��&<�!��%N R����I����f�!�d�e��[LT�4�CD)3�!��5p�rA�i�%id�q�#L !�D����V��- o�Qc]�/!�F�\ �P%�>7�!��� b�!���n�i4�F�[1�$At�R�M!�䎮K��'<��)B4�Ѹg�!��Md���Z$��gn> ��֖D�!�Ğ�d?x�c`� >T����d��Q�!� akZl��$VE�1��βK�!�Ĉ�}�܀A�Y%3�L�%�U7!�!���c��d��M�) 0��)�\�!�23(ԬaѤt.�4H�� �!�M��Ft�ԀĮY0����hВ�!�Dע`�ق���U& ehs��3�!�DK%�����?
�2����!��22�5z%� �]���B+Bj!���!:�2ѯ��'h��i�%nT!�dѢj��A��Ĳ%T����(�>!�$�0�)�M���" G��.)!�jV4�%ņ�H��6�3`�!��W�0�B�Lִ6�lUK�$Y.>�!�DD�aaFϦ1�\�2t"�*�!�� ���E��hB�a��.�rEz`"O�,&��Wd �1� ����"Ol-��^�t,��Љ�-r����"O.�2�
�?t������܋]���I�"O�!(�� �<�'�AT��ѕ"O���a,i�Q�T�W�����"O,��KYC�RՃp���4�&��7"O����$��8����=|"�5"O2�"���9�NtsQ�S�Eu��c"O2�s&��je�q�F�>�ri�!"O�++N�Q�� 0���;�~�h�"Ov��$-l�$�k�舿9,p�"O�!&�R�J�d�j����\��<`"O��rR)E���yD%�6��;�"O��)��B"J�=:�J�$I�% �"O@���J�7=7���N�@[~�	�"O
<R)L'6~�p�G�։W6�в"O�I��ǯ0��&�Y/?�QӢ"O��ѭZ0pfdA�G�U����0"O`\{pF\�k2�I!@�IY��s�"ODq�PD
�G V�q�'2���"O��#"꒨|�a`([0
���"O"!��#�61�W��-#���p"O��[�H�&D����́O���"Ojm��a��v��C�G]`0��"O��qE商��ഩ��^Z2"O&�KҌ�� �O��
U`�"O�4c���q��^���:����y� ��8aâ�^L*1�׉��y"ME��a�lC�O�6���Ղ�y⬓�l�ТO]�IT2�)a�y�	P���h�h?O���+u懠�y��
�~q��Ǟ�BJX�i��Ռ�y�+��s�:l!��P%lX�#'Q��y�'�.*�e�����qХ�#˅�y�/�H]���ꙖmAr9��7�y(�C�⭙�.®6$D��m�7�y"D�o"�,Ӧެ�,0sM�3�y�ꆝt���V�]P�9I�aE6�y�-��81�^-�(���i���y���&D�d�~��d���y��$!dXc�'h�Mi�?�y�$��a���f�M�	J.QF�$�y��"J�v(f@1���H���yj��_�������&�^@e���y"�ǱӀ�cgoݹ�%�'�N��ȓ.u�P &�ޗu,�����!cO��ȓm�^�G�}DD�G�Xw�(��p�Ȩ����?q��!q'��	� ��ȓ���H�����)��37X����A���L�P��"�R�k�:%�ȓ=*j���2;����U$��ȓ'�V���N��7������;1V���M���T���M/�`4�ȓ{��Rɋ�4����+D�(�ڰ�ȓ��7��,J�+M1j�*!��F���xנ�=H�ΨQN^�8�0�ȓM���*GJ��UFh�&�ȋ|0�ȓ;nY��Ü�|+� ��i�ȓH����Hy=�l˴��m�V��ȓ+7�zjY"UNӦk��l��(��j7�Q`.X�:��KfL�e����� ��3���`�R�¢�5þ�������h\ h���"i�0C���S�? ����䜆��ˢ�TR!��Sf"OP�#؈e���E�e����"O�1DH 	H���dV�K%����"OLe���&\������_5y8K�"OB��K�0&�$U�V��r�.���"Oap4C��.�"ё�a�)̐i�f"O� R�9��|3��� t���C"O��;��K,.���uG�(s��4�6"O8�����&�裳E�I���w"O�xȴ��$_?� �"�D�sB�5�"OdT�3���o��4����� `���s"OlU����C|��za	�OC�U��"O`y�e��.0��� �-TN �!���Pc���0�
q���e��!���kt@�s��^JD4b���]!�A;k�j	2�
KHl���#:�!�F�hz��`* $Ik�D�+-D!�ԇ5�f|kw��&4z�Q1�H+)!�D�|���#6!�?hb ����<1�!���2H�P��E^�u"�/ת�!��'P]��Q���o*8�U�ҳ
�!�Қ�j<�Z.7!n����5!��R1K^ʽc�%�,:�PYy"̚�(�!򄒦=U�����V#2�,��2� :W!�RVH�@i)�<p9�C)M�!���'l0���޲`:~�HA	��!�D�]��x���!p�Iw�!�DX%y���˂��/3�:^�!�܂BRp՘&'��Yj���	#8;!�$�&_yp�($��Q��	rw�ľs�!����`�4g�+��u�s�DRz!�*��)�l��+�D��L�%k!��(��aƦ�{�vpK7 �.lS!��5�$�aJ >u�U�P��lm!�d���zL�G��7fr�lN�Ng!�ĕ9LT���b�E_�irҌJFd!�d�0.Y.�cьI^u�WK��n�!�D��Y��ڥo[;>�<��*M1!�1W\���oH��s�iM�!�D��tt�=أ���H�V��[9!�ȡ"��d��@řQs�D�� );W!�䈞X�I{��DG�\r�tU!򄙔K�i���V	9|T0*L�%F!��z�,a�-�QM�eb.I7!��"k�UfD�G5�g_/{!�א]R����ꝼN$Y"te��!�L�`��Tně\r�Y�g�G�;�!�D�:s�=�JJ�fڡ8 d�$H�!�$J>q���P�5܉X �+i�!�Di�Pb0�ݠ%�b��F-:�!�C��(�Ar&H�\�V�#�  �!�
�/l�1gyD�ۥ��/{!��a��R�k�Up�T�v�!��R9�<���NS�[EϚ2�!��F-;�d��֯ü|D6Zd.�$L�!��۶��!��D�Z\0 ���'�!�_�`$��R���[�*X[瀔�Wz!�d'1-"����X�o�0���˄9C!�D����RH�1��Mȶ�K/*!��T�RD
"
��[$��ç��S!�$�*A� ��`U&I���FN�$!��V�e�J��ҧ�&c��)��l��@�!�D�_wH�{��5+��SF�.R�!�d�"|��ɖ�|�\����15�!�� ����>H� �e��(`���"OR	�J �N(t<����K�B\�w"O %y�g!f,p�7ji�"O�X�Ch� RY�X%�їIH$��"Oz)��mC�Ik�IZ�냰k8l�[v"O���"k3y6�2�kݡ&TT��S"O>�Ca�e�uT!�i=8�q4"O�R��4!��!p�L&Yzd!"Obu�P̒&u��kσ b4���"O��
@��^8BЖ�I�I"R�:'"OМ���B-mV٠�.R"/����"O:�P� �C[����^�Z��e�"Of��w�K$
wx�c�Ugz����"OPT�r�S�?�S� �7�앲�"Od�Bc${��|K�V6Gy�P"OJ:��-�����ЋI�h	0"O�*M�-P�F�'$O�>�tuv"OH	 
��i�ĸ ��"�� �"O�=�Ã-sn����o��a�6�"6"O�|�bΜ#`� ]3W���Vp�(�"OH��Mːk���4U鸁�ri�y���p��y��Zٚ@��A��yR� $\F��2��#r�i˅�F.�y��+L�n�ad�� v`�5���y��*t��)�E��,MCR4�k�y���;����E�?4a�3��.�yRŷyPܰ!PƝ�@,|M�"�ޛ�y�������N�6t]�eDS��y2�}�2�#���T@�d�Z�y�F��`���2�'�2[���	����y�D�0s����A�0T��Qs֏ ��y2�OGh���!�,I�
f�T%�y*^8c���:�d�2E�.m���ܗ�y��'^>V}Kg�=���GU��y��X�%�+4���8�:��@�y"(_#.f��W��}E���a��"�y��"p�L�;�%�'#yT�&�+�y�`Hw
��X�������yR�	�i�X�U��k�@�V"P��y��8֔��H�_�v�`�I]��y��2�6#��^��kg�U��y��B�J���qG�2E��1KT��y҇�(�� �L�?2��e���y��'��9b�ӑ6O4x�E���y��E�9�qr��.�D��3��y�M�Vw ����	�2-Q#���y"'�K��Q�	�/a��9��΅��yRH�1S���ӄ�V�M�6	�!�y��yPYA���H��s�@0�y� T?Tl8���*C�U�.��yb�Q�P �l�Ν�B�[!�y��0@�� 2Bȗ�X
����7�y�.�Uz�2���7h'�˔����y2ߧ}AL$)�a��r�F(��NG��y�
2�H��ɧif��d���y"-ʝ3'�q�$��2��Ѣt���y�$J� �4@� ��/��cF��yBG� ��	�@��z��Y�dD��yb흞/�
���Q�%������K��y��ME�*b�#W$�0i'���PyR˻D�r���e_'}���j�r�<Q�(NU��ӕ�*z
.�*U�u�<�P�_(�24`ͪA�����t�<�u��)<5P!/\�3����o�<� t�pg�E�z��c� }�f"Oh 3g��t����ǉ>-���h�"O�|ƎEW}�)C��}�P�7"O��� ���rK≈�a�$��yF"O�(�E�a�\�R4@��$�J�zu"O�1�L�s"�R�.Y�ܙ��"O\�`�
��ݬ�hu��6vHqAB"O����
6v^���o��u_L��"O6��Tk768&&�p.n!u"O4a�܊qf ���=>�ؑ$"O�
u�٩N�:�pq� ��"O�$]8b{��[���VQ�"O^�$�G&
R\��Ā�@zE1W"O�}�2��1v�����F[���"O��ǆ!�����)��y�Q��"O����Cu��PdO�. n`��"O�ؓ��D��3E�<Zd��3"O��� ͦR��z�m�:
#�99�"O�V+��Lp��(��R�rr6���"O����-��<���
fm`Q("OQ��mϛ����HS�aXV�: "O��G.�%��JS�xL �Y�"O0L �K
I �� �T� E�Y�"OVY��dՆL°�cI#<���"O���&��1;q����,N8��%"Oj�r��T�Q� ��[��������y"K�4B�H@@��[k��yP�;�ynטh匵��%Ő_�f������y��W8Y�X1���K��I�gOR��y��v���A�GG��M{����y��4&.R��P4Ab�5Q�'��y�(P��=B$��7>�y�oJ��yR���m�&��q-ޯz�$cA��y��:�j�ŤJ�R]3���y�"�^Lܭ�'jپO*�)�r���y�L������I1_"�i�J���y�`�"	 (�@`ɄT&3eR&�y2m֪̶��ujQ�c��Z#GK�y�R�.9��;Q+��U,=��fߏ�yrN��JT؊�D�Q�hpc�_�y�#���PR�
�Et�Eoɔ�y2�}�jE+׋8ȸq�R�ܢ�yr�+Cź�`tD�&19Ԑ����yb�C�L�T�ņ�/S����@�3�yRl�� ڤ�����~��Ȱ����y�����-�B���s_�T*W����y���)DTtɀ��V6�ApƉ
��yR��#��2N^3<;ܑ�b��"�y�+��ʆG��+������3�ybl�u����Śs�ٕ�1�y�c%V>6����ׄs��!ʕ+"�y2�Ŷ�05�g�#W5��S@�݂�y��NH1 ���G�@1�_��s�'9�p	��;R����K��"�'_*ġ"�ϛP��`�UH����'��Iy��K?;�N��������q�'�֘�pI	<Z���*�#N��l�'O���ߨ0���)v�UI�
�Q�'�V�Q� ���䏣<B��"O^`��A��B�z�Ӕ��iIK�"O�Y�/�,5�7�c�(�"OH��qc�7!Nn\)Beɤ;t䨋"O����X�8�<�AX�:wXӱ"OhDȵ&F<~��Ǐ)k��mK&"O� ft%�j��U"bH׹`~���p"O0ǂf��PJ�!g��`�"O��ҮX����(V,P"Of�Óĝ�� ��j	uU�l�"O(�S���4:n���o��K��K�"O,kR�W�]�����BxB��QG"Ov�U'Z�LP {T��\B҆"O��Fhզ�D�C��t���"O���]�N�h`�d��@�@��*O �{2�3NAX�!C��z$^��	�'���@$L�	!�hܠ$�̾n��9(�'2��r���`p�F@�#/��}�
�'Ô�cgm� k>���� *��}
�'|<2��P�TI�m��)Jh�j�'�Ni�HC��.�"����VHm"�'��04�|a�!F͗���Y��'I�q�!�}�f�۱Ft�*�'c�� �Z���HE.1�����'\���dϳ/ �Z4�'�v	��'��lz�M �e�J<0��Q����
�'� ��V� R����:@��(b�'����G�J�Y�(���ą'+F	��'�t�I�L(v�ݓ$�1>J5��'�(�
����r��T�ۡ{�M��'+"��cgh�b�Æ�N>���'�Z�������x�(��D���
�'��(
��Ñr`j��u'�?��

�'�"����QH����1� b�'ީ35Þ�c�x�xU������'"N;�N_.x0m��Ϛ�
1��'i���Ș%�ĥ	C�8 � j
�'���kR�*L��	�' /v�Ɣ��'���#7Un�q��EȎq��'u�xR����Q<.���/үK;��
�'��\@�� �x�{a�9o�ĭ�	�'U�\��iF2y��a��F�3_�l�	�'�>���ڭ!۾d��73x��B	�'y@�z�N^p8��A�}�Dlz�'v$Y�-ATCMA�/U�g�l��'�|�6A3YT5�Q/Y�S[�[��͹���P��%Ҏ	���#P"O���b&�"�dA	uN*&~��p"OnM0+��m��Ј��`�a�#"O.�x�CN�~����')�1b\�(C"O\r`�ޕu缈X#��.k��D"O�����u�f�p ��*E<��p"O��[�+��r�吣.DCfh��"O��!�l�/{5�[��&-����"O*�v!�ʂ�:E'�4�PP"O�9��Q�$�����Џ?>��"ON�شM͢U��\�2F�r-f�a�"O��R�K=<"�h��˨,wQ*1"ODA�&W�R,�y�!̞K"Ȱ""O�j��r��y�`��	V���"O�4���G�t�\��O��F> �!"ODtAD:6� 9[��	�" M 7"Obq� ɑ5�b���-�1� "O�e��ť?�=���$ A� "O��#�4Ϝ�)����,Biң"OέZC �	>x��E�
��"O<QR�װ2s�(���Q�7�.]��"Od��o[�4��h9��0�T��f"O\K���g\ݙ�6'��!"O����b��.��	�_7n�hW"O� ��[iɀ(���[�º4(~��D"OA�����,85�тn"��"Ode�WLM.x3���E��?y� ��"O������LӚ����ȆPm̜��"OB�+JHP>�xG��:�h|� "OX�)A�~@L��Ì$���AW"O��8SKL�hC`���B�0�!��"Ov��Iߩr^��r�B�2�>��"Ol�y�427�|'a�B��"O��G�\Xe��fYxJ8ejr"O�l�4�Sn�zH��@(8�9��"O�!� �ڹV> �Ę�"0d�@"Ox�1w�ٞ@����PNոb(0�"Oܼ �oY;uj�)�"ǋ���"OV4c��S�TRF����&]��Q�"Ol��wNP��ViP��#�.`B�"O(\�S��k��8`�EԊ|0"O
`X�I�?�r@i���Q����"O���qjT�=U�z�L�u��L16"O���Ō�v��E�Ek�$r�8���"O�p�vg�"�ԁ�	�/v,��"O��kլ� l��cGgϭ v��w"O�H@c�C 7��hh��P�VQ�#"O�ݒրʙWŀ�K5�W�L�Z���"O�%�)ؼ����f�9K3"O�8+� QN�7Dܯz`*A�2"O�kum��Pub鱖�Y8t!��"O.l��/��H�����S�g}�Da�"O���uE�9�F���L�3m�9H�"O��1�(�g�@��3��$�BU8q"Ov,��?�t;���j�zP"O`	K��۴c��DC���pN~���"O�AP��UI�!����]J��D"O|(��,M�,��@�۽D& ,�T"O�`BA��x�Tk�G�xZ���"OV3�J���BY��I�
>��"O�$;��ٿ�&!�1�P�^E"�J�"OvI��f�4�+Ʈ��'�1��"O����!��y�l(�,���l��"O�����W7Tr¬<5]$ ��"O�}���%��0LѕGEZ���"O�|�$�͕�+�+-^��"O��hׯgdru�A��62\��"OY9q��6H�4�#ч"���""O,)��a�%OE"�A
\<t�ɒ"O��Ç�c�n�%�11'�$1�"O�M�gE�9�Q����2B��6"O��Ȁ.EY�J}��S!�!�"OBL���'Ն4-ԤA���bv"O����9( �1�(u�TP�"O }yd a��=���B4��#�"O�L�UN�1���*�ɛ�}�&�#�"O��h� D�z2��NY�\���"O\��Z8�	6/���, �'Z�!�GJ�X���8(��H&X	�!�d�=.��q�� 
܀xBÖ�p�!�]�F�j�c��Лm��jqB��m!�DMy��y
b����u�RD!�$ڬ?���smFq$�y!��!�D�f�t��IY�o�f���V�!�d�05�P����9Y�P�`g�N�!��9�52.K���`�`�Zi�!�̎t�@dB٭@�>����|�!�D2���H��ڐ2�H��rk�:T�!�� �}kFkO�Q�ш�4R��
�"Oؠ[�L�,J��s〆�c �Y`"O �qL�����)�_�A���"OD���,L�Xi@��.}in\2�"OXt�4-�=�Ȩ
����7K�y�U"O�	QiE�o.��!b W�-4H��e"ON�����~.tȰN"3x�U"Op=��#Ү=JŋA�� o����"O��;d�ĨHE���KǑS�Yie"ORtC�_�B j9��뒭G��t�"O"����r
�`�«G&�"O�, a���Krd�OE#L�$
�"Or�x&h�)P�۴�~��R"O��j&&�8,JѩN��?¼� "O�9�U�G]�,�!LW���Mc�"OP�[��Xжu��K|H��p"O��i�.�ZL�]�WIǄe����G"O|@SH
�Pfi��iP9=�);"Oh@#c�/�r̠4
��?��Q"O�A)Ej�3Y�YZԮC3�t\�"O`�t���eR�9�f�I!=�,��#"OH}@Q {��A�B����hf"O��:F��M�f�q�Q8]���Z�"O�l"��?HX��C�A��8��@�"O�@�K�}�X�!Ђּ(�Tͩc"OF	�g�ɼ���a'-�d�"O^uq��! n��p��_�8�"O�����V2,�(�2ƐXm��s"O��2w'ޝR4�pJ���QkD�C�"OL��@ܪ&J�F�r��"O�͑A�H�J]L�z%A)M(��"O��IU8�U�b݁uv0��"Ot qb�yI��{Ђ�=5�!g"O��!��0�
�8�K@��R�"Ouk�G��$��KR6(Y�`��"Od���-�"ܠ�`ğ�%kN]�"O���@���TâEɺm�ޡZ�"O���ň]�2�0GEG;8���C"O�L0WE]`��ң�F��j"O�(B�%G\�P6�ˍn�^���"O�0��Grs�e�0�[��2��P"OZ�BՍA�24���s�:2Ӭ�{�"O��1�N�$N.��d/�4B�X\D"O�2�/׉c|����B
i��ܲG"Oz5 �J6"��ea�[��5��"O�А��5�-#�F
jLViY�"O�a�$F�E�Ƽ��DĢR�°"Oqk��W  S\m�v�Ё:© "O=��#QGK,HOj���"O���a�ȱun�<#�6���	B"O���pA�)f҄
���!mzy�"O ���*�;h����a�/���"O
��,N��LYaǂ�<�Ե(t"O�!A�I�Y+f1�w�Y�C�
B"Op�H�L�{u��Ðj[�:_�@��"O�X�DF,q�P{���6/B���D"O&=�4MGwƊ�0GP	̶8j$"O�)�����%t��L	�"O�i���n��]�E��5�N��"Oz}3QE��
L�X��jQ� }1E"Oh�N@�?�R�#U�P���"O薁��,a�ϳD���v"O(QY��B�OX��	{�"OΘx1�T.��i&�-h���7"O� ��s���B�R��M#|q��1f"O �AO!lHnj��'e�ł�"OV�@0��WfjACm�0ֈ8!"O�a4+0��AiD,[!F��e�<i&"�Y7��9Q	1O[0P��(�e�<�s���k/2}���6KT�9�Dn�d�<Q�K^�?�L��E���M+R��^�<a``��ZK���㈲g!t�A�#Pq�<�v���p�0�dY�e�f��U��q�<ٵ��*u�|0ʚ,Tv�{�c�<!`�'�� �l�JE�Oz�<�]zN�s�N�L��1�CD��	��C�I�"N����a�6�a�ŝ�W��C�I'��x@������C�!^<Y�C�ɠZ�n��ß;u�
�@�G&W�C�I7ʈ(c��1#��h���u xC�ɠ0Τ��IH3j�f( ��"V�C�	�1�ܤE�@2�j�	dFǉv��B�I��a��*�?
��+��F�j�C��.Q3y{�!R/M���iA���:B䉙dT$�q�UW����q��C��=F���C�B �N�v ic�R�Hf�C�ət�\��ᘢZNB�@C�i�*C�->9Xe�<d�.�H3琖H��B�I�9(&h�F,
�4$��	u��45*C�I�R�Ќ;�MT@��x�T�J�}*C� q0��a�W�1�lbR��A�B��<i5�pE�W�MB����!s�B��8�B):�YS��*��a_�B�	�b����%+��E��2��F�N�B�	+6�(Y3��ܮ�{�g�~5�B�ə�aI�	 �z��K�\B䉣G�X�{��&�d0�e!C�<2vB䉆_��0���I�N���A<�lB��{"��EF���Q��ޡP*JB�� R]�\1��^��ۥΞ�-FB�	��EiD��(DȜ�D&4B�	<�6`+X����W�C��?\]�#Ai~f����EY1��C�ɣ1H�dy`�!o::�;!�� C�	�i��WbT=y`ZH1�&֤^��B�I�>����anJ,2��c�3k��B�9�@��2@ (#�*����Q�w��B� j���J�M+ �>A�\�d�B�������/FA>��+""��C䉫�|�4�F|&�Z�`��NrC�I�E1�-;q�ؖQ̍��J�|��C�	�]�d�BA��U�3̊� J�B�	7zM�t��RW�$$r��J�C��B�I�1�Ah��!@��sh��� B�I6P$Z(���'I�C���6B�ɂ>�80��,v���c��!xo�C䉣u�*�x���+.Lpi�i%8�C�I�t ��J'.F(:QD�)�͓"I=C�ɩZY��9C  �g�&QIӬT0b��B�I6�⠁e� w����(�l��C�I����#j�#2 �����C�	(�YBq��"S[��P��WݶC䉲%�I�T��	��h�T�~C�I�u�h\�'i�.Y�(J��*�HC�	�{�=R�Ɣ.|C�X�@c�*�FC��rn�IK�ß�.j�@A��Ѫ��B��3ScD���!oQ�����;�B�	�*��q��L�	ab���c�1T��B�)� x����9(�iAt���=zG"Oΐ� ͈B�}�$ @��1P"O�;c��M�����g4*=ad"O<��QI�_qfAYD�e@�13a"OR��� U���q[T!���%"OB|C!<s��hF���B,�"Oށ:E�h) ��e�ʥ|L�5�"O���5(��M`�
�8C9'"O�E��b!B��q��KO�u;�8��"O�t�	V�}�Ha�A_*�|c�"O� �F���l ���ֵN�4�bF"O8�:���������p����"OP���!тc����@���!K��v"O� Z�l�#��0��K�_C��Z�"O��S!k�'@(��/�6;.�L+�"O*��ʏ�D�a����i(�`"O�9�N:��!��΋i����"Oh���93 ������$�tTc@"O���R����%��5�p=�"O2��A����N�Y�@ɱ=�����"O�!8��ގs^`m�G��+1~Z�I%"O�����R�N���cÉ`{�"0"O�8i�T�v�h�� A��vr܄�s"O|��7 ���S@-)�\e��"O�s�H6��MR�R6n�,��P"O$�A�
�T �q�B��^�� ��"O�̢D�'��U8�-T��Kf"O��q��'8����a�gq��"O����J�"�@��B�G2̀�"O��V�:0�.L��fU�8����"O@�ٔBe���S�#�M%T	�G"O���#���o`ic��<,q��Q"O��9��US(r�@����ȼ�Sc"Oda���_^�H�aa�~��	2�"Ox��rʲ����!�ƫ
��<a�"O:)�'DW-=�ZP����&;���P�"O.�
�@��e¹��)\�v���V"O��ц�N�0���w�Ǧ$ܼ� "OB��e�_5L3J��t�Wi���d"O|�{sF�y�lÇe���$��"O&@25.��2����W�Lr�T�!�D��>���طI�5r w�ÿ�!��d2V��Po8� sr�A�!���9���1�\�B�m��Ϝ�(�!�T�a��]U��.)��S!��	�!�ċ�s��jFÎT���g�P��!�Bt��H3�&�bhs���#~!�DU �}#0�]ui�Qhb��c�!���N�6�;�N�2]*8مD��i�!�Br 	yr�F�N�D�"e
Ƚ-�!�"��CB�S��$e�'r!�DƓ	�Ȝ�!�{w���uMvT!��_�{\9��d�g5;^���ȓk.P�dL:t��ưO]6�� ����ă$��%螪P�8�ȓ��a7hM�>�^$J䀍�e�f��ȓF�0Ѓ85��ՙ�nÛ+��I��J���1��X1]�#G��6}fx��P�����fҗN_tdkv �CjC�ɀ`�P(�o.򂑱�-��IzC�I0w|H1�ĺEz�%�!ffRC�ɦP�$!��C*tE�pe��bX�B�	�$9l(�uFНx܎tr�,��4��B䉾 ?�L��ğt#���"o��IvB�)� �Hg���, 8��D�/�.��"O@l��D�Y�� ���!K_Ҭq�"O0� ���Qx�Տ�?Q�x�i�"O��W�9#5T��rL�w{^ŀ"O�*������R�._���"O��{���#�0�٦Zu���"O�����E���4*H�iY����"O2�Br��7(�T��[
{G��)�"O*�1�铵 3�IA�Ƒ�Dұ��"O�+�hE�D%���EB��@"O�da�'� '�zX7jP�%I���"O���	�<7v��{��F3�cs"Of��
�4Q7����h��b:��"O����a�$��珫S|�ɲ*O�@�V� F`�ȏ�x���h�'�HaJ�ƂuF I D�VC�����'52�	��M$�K�(�JR��Y	�'ir�k	P�FhPrJ��0��'�����"%_��`Ѓ����[�'�6 15�ƿ(
f�# nC�B���y�@LK�&}�w�r!eQ�N�̠��'V�T��X%�<��ƍ�EDTP��'�b}�Bk
��1�гA���'j�8��	}z����aS
*����'���fM2�ڕ� i��p�l�X�'�\���Cop]`(�h� ܳ�'���H� q�)�����p�P1��'�T@W�60�W��p�81��'�����,�v)3E�o�X	�'j,���B�&1v�U�Հǫn�Fɳ�'�i ���%�Ϫ_��-��K^�<�䥚�mx��ф��>$����� B�<��J09�R ���X�Lt� 
�B�<qA�C�hF�y%��I;�034a_A�<yҬ;� �q�e�N`Pq{�jJ|�<9)�@�}��I�F�H���R�<I�
?s��1���@��*B|��ȓN(v��ƪ}�^��a���h�ȓj`�Xc�A��MElP�DnxE�ȓm��p�^���� y�v�ȓ ��4P�&A./����'c`��ȓ9��xF͌3��%���C>�&�ȓTp���g�\�p�h\��LTKT���ZЬ�B�g
t*�IET7u�T���h�❒%Nä.W�u��K^�Y��ćȓyЍq�4T_����E�g ���ȓBy��C�J�R��ԡ��Q襇ȓ.% %
$�V[R�Z,��ȓ\W��S�l�&�xH���(Rz��ȓQ�bt�t=�(��G' g✆ȓX�bĀE��>A��)��O!_�,|�ȓ"X,Z�`���A��
���M��i�������r粘2 �^�l%�ȓ}6r蛊|Bh���ah�j܅�1C`�mPi!��̋?Kl������������M*��#$�@��T����H�TY�cYO��Մ�b���-H�0K��+��ľ82@x�ȓ���b&�I�PY��ID��2���ȓZ��)��v+D4k�#q���ȓ;�,rE�]�g)�`#Jĉzn�ȓ7^��#X�@Ѩ�ɰ#.!	�"O��+ ��=������%�0�
 "Ob!T�va��ܦ!�F�Q���<}�!�� � ��Y�,�N���ďF�hX��"O��ō*Q	�h!��I��,��r"O���K]&U�PL�u��\��"O�3ҡF�u@tqa��Nh�$"O�����ӱ$�����K8(O�A�"O�I� �Y%�mi�� �ak���B"OL쁱/ݰf��d�N�ܸ��"O|��#C�X�c�B�0�ƭ2�"O*���"`���Ľc����I@��ybN�_�p��JX{`C���yR���"c@�C��)V��`�eR5�y���f@Q��f�wN +R��y� �!Q)>	+���%va&8ZVHG$�y�м.����/\
��M@�(Ʀ�yb��A��]�Э\����#W�"�y�L՝,&h)K"[d͛��y�j����%!5,U�3e��y���0"*z�u���R�Ӄ���yRWP�0)����Dz	�G�yRË�2%��a�GӖ2q��(0�yҤՠ�Zc�
%��8C�V��yb�& ���D,nI�Dqb7�y�ɔ5���tNu� u�@h�$�yrF��x�%�VQ�y3�A�y�Iɑ@"(�`�S4M���ؑ�ybBj�@4h�#�6pTzec��6�yR�l�D �oA,ktjM����yrg��^�xŐ�Z7\����22�y"DC�:��ʑdT� ��y,���yr�B�.	H�㠂2�^��K���yrdO$q���>@��������y�

�%��e��PJ��t�H��y��Lz���Ɖ�K��ണv�ȓ^��)���/���6�ޡ.1,4�ȓ&q!@Y6rV4a���+T��*�$`��ݙgx&���[lvńȓ�P�Ì,!��/>Nfj-�ȓ����/ zk���'�d��ą�<�%	�����-�֪ɝ1"��ȓf�TY�,� ]nI�щE$b��W��\ �㍌=�FP�&� >���ȓ	����B�s&8�ҕ����"O�Ր@V;��][`�8 ZM6"O�=�BmO+T���:�!��3QT��t"O�0cR�_�F���ɔKV��"O�	+7b@��|����O,0M�-��"O���pĀ�n�@Y��߂04�<��"O�e����8���	���eR���"O:݋2�75H�AW`��l沜�4"O
�Q��2�!��"N����"O�H0ď-gr,BǈM�y{4"O�]�q_
:���'P����"O��H�^$QB7EƊ�P�`"O���t+�4^Z�=� ONm�b�s"O.���A�l1�I�V�:(�z)�"O�-��/��1�����F�xq�"O4%�"l/�F!o�n8�"O��p��)�ؙ�5���U�"x�"O*��L6iԚ��Ō�l�����"OU��͝1�$0(p"�Y',m��"O����j� 3�40�ߟiZ$�"O����a�q����!1j<#r"O�QSB!I�U����W��f%��H�"O(�9�H��qC�oCt|I�$"O� ������(a����c�"L�"O,\�Bg^9��l���Q']��}KS"Ox�2��g]��ƀ؂t�4�z�"O���Ч� Q��arɃ�l4�#T"O�UӶ�Ĉ�N̠���oO�!
�"O�[P-�?tM�"Uǟ7+kL��"O��d�'_�� ���[�C	�(D"O�mh��҂0�(|C��I� ��"O�L 4���͜1�d��(�bšf"O��!�)�2�Z�H�^�r9�F"OZXÅA��U�rT@�ύ�i�"\`�"O� �!X
���0��W �l� "OrS��;$�	����%��`BB"O,)+0�@�;��13�N�H\��"O�p�b��5xD�j�o
�eq"O$Mz�(	k��fj�i�@ �"O� �Q�R�b.��˝�/|���"O��+��K4H���C�
ʦjzD�6"Otj�������&�\�`ۃ"O�`rh��:�*�A!L-��h�a"O�Ě�AH+wn���j^zrY��"OH����2uܔ���̋� c�U��"O�@0�52H�;A�Dv�ۑ"O&�S0C
%�R�+�b�&%�(��"O �2G��SNƙ:��#m���{!"O���G�-{2�V&�#�8��"OƬr�C�+� �C��W\�D�"O����#
�R�R%�'x� ��"O�!��'�]���He#A5r�\���"O��5s�h����f�E�T"O
tx���H���а!/As�,��"O�9����b�v0CE#�=���`&"O��{�	��
�!��5��|�`"OHТP�6U����!BP�/��d�q"O�A�oG �8PJs!�{w�܋�"O&L�Q��;�AP�m�6�
Qj"O���s������	��8Z���*V"OjR�[�I9XYA�N��c�H�iV"ORђĪ_�g\z�B3˞�Cv�4�"O ����ھ}I��!$�fC6"Ori��I��ĭ���.J_&r""O ,��D�?;\<@1cEJN� �B"Od�Q���.�d�5�*f.�a�q"O4� �L�¡�Я��~$9��"O��j6�� �~�� �.e�`Y3"O�y�sdŲp��@[!1��ɪ�"Ovp�f�E;>��30,
��阡"O�2caަt����/��E�D���"O�`fB��&Bh<H���|w��i�"O̩I�cD�|vV�x@ N?en� E"ORuy,'~1ֽ��o��Q�`@A"O:-AƄ�k����Y")�0"O���V#Lch��CK�.G
X5"O����HU�3����b�.�B�c�"O1��h+��1�A�7f��@q"Oވ�q�	�l1�x!�艚)VV�1�"O��M�&|��g(�<Pe�x�"O8ar$�X�P�h�s�b�Yr"O(i;ƪD4TC��re %#�X�St"O��G&�%��h��7Ǥ��R"OLH��!�'2| ��d�Ƙ��@�"O2`�$T�RH�2A�V�R�r"O���a)Q8�-ـ��0t�}�!"O���GC	+$en�����0G֭J�"O� rhA`,ę_����C΂BʔC�"OЙ�w��'a���!Aj�b�b"O
a�q)٬.|aۇ�ޔD7N$��"O����1�F��i�"�v���"O�-�U�uL��PE�A�$���Z�"Oh4��H�-J&��1��B�*�:"OJ�S
hwf0����V�Ь&"O�aI��(�X�땋��|*8��"O���g��1����)_� ��J�"OP@�n�%�sPiK��a�b"O����;G� �5�R�<�"�p3"O2�clܡK}F�v�Y�j@)�"O4l��\WV�9uE�"��%�"O&���1Y"��V
� o\�:t"O�,"7���I����JG� C����"O�=�!��-�`��T�I S���"O`�"L�Bb"�����J킅"Oz� !�O00r�Lp�%)y�Qѕ�'� ��F� �Z��1�׳31�p�فm��O2�=��(��IH<-Y:��0��D)���y�Gz��Ï<y���K��y��1��!�u�R�<��A��y2�ɿe�Q�8�Ӌ_�t=0�P��F��"D�T0B�C@�^\#�k�&Z2��w�+D��!��A��jj�I�+���F�*��hO�S"-܂PxLCPXdX��- 9I�pB�ɧ3W�����z�xP�c�� u�,��D&?����l�	o�]@&� �"ެ���6Sl���杺S?ؽ�'" � MGy��'����Q�|��RR��>�M��'e4Q3ǨY�x�`��XbvZ��'" I����I8ևXM�`2�'6V�# ?#�ĝ��#ŵV蠂�O�x��Eׅ:���a�V��9��"OL��U�3Z�"�7�(� 3"Ob�r�Aq�Pȳ����~Q<��"O����SF�hw�[�Gܮ��"O:���FـT�\ҰDA�Go$�S��yBȒ	�M�`\/{@�"��ء�x��'��c�����]2��_^l���C�� G{���َS�pDӇG����-�E�ܝ�y�k�0��Q��&X�%h��y2��7r{�A9Pưa���Q�T;�y��K.�ش��Jn�  ��
�y�*&vAB�K!j�#ELA8Q�yRC
/V�j��:N�5x�k��y	ɂU��JG�@�	����A'�8��'a{�ϟo����j��@ [�]��y�L�tP�E�7�=lX�!�f��y��˽K�1��OE� Z�D����2�O\���0Z�`�)��).m���P�p��	�� �P�N��#�TpA�N^ƠB��)g�zL���D�`� �PW�M�����j�r⟜y@BTD��k�O��D2@<?I�4�?��y�$ߔ }�T*B�	(z��Qe������E{��:�[AA(|H���s ��a"O6(�6�J�t��Ϙ&iJ*��f}�|�V�̉@��P�F be�˺;�t�sE�L�<�X*M�D��&���3ڬ��m�<��A�)ր)��t�� �N�<�ԊV=J	��Q�; ��B�Φ͇ �P��>v����A�NEy������]�IF=��պn�<�!�j�K'!���X�k�� ���0v�;(���<,O� �C��1E���K":���C"O4���/T0�1X%,�T@ȑ�"OV��U%�`K.9�Ԋ %�����7a'?�a���c�FY��Ñ/w�=��C Mh<�Q���!�z��En�Q�V]R�o�t}�9�S�O�J)�ʜuL(1��F'@I��'�y�iۥH�pű*��@_��"�y��)擌,:ֱ㕌�J�&h0���C�I+����Oי���y�k@��C�I��w�'-9�� t��/_҆C�	�![Ų��-����@�	:�B�(;�LЫB�T�GG|��];Ԇ���2B�l9Q@#�n����*�=4��ـ,Yd�߻>��ɖ��;{d��ȓW�t"�	���|�5j��<�ȓ_ ]�u�X)ʅ�V�0���ȓ[��3�$̀C�`T-ɬ8)�|��w �a2ɍ�&u:�wI8:]n�?��}�h�)b͒�X�,(˰�\�^���kar�CFL�0�� ��h��z��a��f t3w퀔X_����)V6%����h��}�����p�̙b�*S�8K���m�2�ч��*z�.D��$�5H�0�ȓJ�MYE.Z �x�΅�]����2����µ*�a֎We��QJ�4��$3�O����B
%�-�ЧύU�dTPQX�,D{��))$6����M�g���C��	p!�$�	|���PWD/��S�da|r�|�$�"'���h�&��̔��y-4�4��ޡ/� �6����y2JX#�^� �Ӈ 	�]k1��yRHб/6&�BK���v\�c���yr(0���ӡA~��@��'B��yR�	0:�S�悜`n<a;��Y��HO��$')2�+Ռ	DC��G7D�!�D̨J��pC&�-.��A��~!���"01~uk�	VdW(�7�W�`z!��I%sRP�4lB�%?N��N�!>�{R�ǒ:��9���Ru�4@�m�*R1On�=�|j�n�&��4Pe��/B�,3��i�'-ў�B��[�
<s�BH Ӄy[���q��wNYS�P��LS�u� i��R����7�_�g2�����C� eO"�PR	�"b.�K�(�-HN���"O�qs)��w�!0$a��� @kp"Ov���V�&i����� J�����aX��p�j�Y¹��jU�S
�6/(D�,���ϠNdp5�2e�Ըʢ�fӊB�'\Z~���'��J���3�i��/
�����+�~B1O ��2��PD�#�X%SE�E1bK�<����V� ە�!��[�'6��6A��)�DڏOM:�Z�"ĬK�!�D��2�a�Y�m��	elO�U��6��v���������#lLXI0�I�����'O���fnۅw��+!��"n�EI�_�<鰇P0_>ZS�Y�P��h�bΤ#ў"~�	�:FĠ�B�!d:���#%���C�Ib�b�X�J]�Ȯ��*R�C��#1F�[&jN�/�`�W�N	X*�B�IH�R�.9�<�Sj�<i|�hO>�[�Il�م�!.��`���:D���$FzaȄ2`�%'���	��%D��ak��
�|���Ŋ�(�U�F`"扟(drT�,�����Ot�1%�/e�2���!�m��"O� X� /��B�:Q�W�	BpP2�"O�0�R��5�8�Ү���|�e"O����"[<L>�J҈Օq�85�t"OT-A��4AɚY��CdĴ���"O�t:C��/oR�P�œՁ"O���Qƙ'E��($�7�ؚ���&���+W(!!/E�u��U��g�+b]���ȓ��X��l�_e�1�3��U�@QDy��{��#��b�_�q4f�Tf��(T�k����?a$I�H��Z�na�&e�i�<���D2N`5�bB�"��� 3J|}��)ҧ����D	xB�t���GM���ȓi:0jâ�5:�`�ksȂ����'%�I��8�A��%[�Ex�Z�[aB��g�І�ɏ7$�j6g˓N�UK$�O3EZ�B�I�h��V@�w�AҥC�eT�B�I?SG�鐄�݁�j����[�k�~C��%�<)B�TL�*aA6HM 8�C�I /
`9����;S��$M�"P�B�	"7QF@�C Y�]O���B6r��B�+!�૵�I'I����v��r�C�IdgP��j�K���	 �}��C䉒$�X]�p� �L�"�� _6kېB䉦-��h@��5G ��*[Kt�C�o9�9�ҪE�>�6�U�ן]7zB�	�X�JAQ�q{ZQ�b�(�B�ɢ//�U2@.W �&��w�� {�C�嘥� cJ!>������\�C�	�,u�0Ⓝ� QA:X@U��Mw!�$U�UQ��� g�_�X�[��ҲQ!�Dܵ:�\)�3�X�]DmG ��7s!�D#~��Q�f!O�1 ڹ�3e��S!�d]  +��d��-D[̩PKL��!��˵	k�"A�� NUШ�>12!��OmܚM`���
u�V9 %&ʸb�!�dB�X�r๥��=e�E�r!�Ğ'qnܵ��E۫}*R �ң�Aa!�$*�%( ��9@'*�seB^.+_!��{�T�v�l���a��W!�^:��=z���,�9`I�c�!�$�]g�I3T$�.l<�S$���T�!��߬
t�q��$Z�k�}�G��5o!�U�y����U�=�\YIɂ8l�!�$��E�=�Nة�m�!%Χ�!��)%Ǆ�CB��31���� (j!��/���rlQ���B⇩*c!�E![A��c��	,h�>�HOT�q�!�$n�И8!隝c�h�h4��\g!��#��h��dZ��A���ˈQ!�d�N�%bW�{�F����ʓ 2!��R�PЫ�°P�$5*šV�2�x���>m�60sU�� Uaz���I2��!a/��9q��b����y��ְn���{2��esp�������y"�I V.�h���Y�������yBEÛfhR���`?���4D%�y���U<�M��'���%L@�Q@��ȓ(�Z��E��;>9������ 	�ȓP~�%�aa�<z� �� �
>�J��Ś����1$���[�_����2�n�a6b*��h�Θ�*`�]�ȓ�:��d'a1D��0�JD.(��gDa�!\�,�88Is�k��3D���6��52�(�%\�)p���'b,D���bI�x�0���jI<:��q�%%(D�� 2��4$�>Y�.�Zf͘<%'��3"O�0�D�2+�`��-�ݙT"O\�Aj�*�̉ЂV�Jk* �"O6�I�	�'~f�q�'4QzIp"O��a�A���$#���)1؅"C"O����N�h�x�����'#���"O�ղ%�G�+��P� 4Y�z�S�"O{��R�@U���Ww�L�"O9��K�y?� E:9�~b"O��`�H��Ųe��Y���"O0�e��L��O�]���kQ"O[4m~Nt�)t�4>����"OtБ�����І��%����"O89�b�� �~dH��F�=�s"O2Ъ�7�d:�
M^��@�6"O�;W�P��(�iЉL?�Ρ2"O�t�� s��9�!G5z���8�"O����Y�4�"���B��,ٰ0��"O�@�7i��@c6Ha5�]�U�.���"O�����(�Н��#_2T�d��"O��BG*D7�L�)q�L"Rb}d"O2�sB!�v��5���	��u�"O֕�A��>�q�/To���"O�q��G�x\1CoA~�9�"OT �`�^��ve��$IT��"O��!��:���%��6}<b����� ^`�\؋�Y��7��9Y�fX;k�,V:�T��m9D�� �V5:Ot��wf��No����7?��o
�������D�= �XT��(\./N�-�#�'3����	ry��H8!���1"ƒ��d��aƧ���j��1G&,O,�y�M��T�|�С�5.x�q�5-~�i �R��$D�C@�0|R���䏛�T̽ㅦ��}�.��'$�A
VD
~�=(��F"� �q"_%baF��(O2��f៊�Y��C��'�� '��26>2Yri�ޒ�(��x��{��ejq��.1�<勁�	ohu�w͞'0b�bC��?��'�|�y�	?�Iޕ{h�@�Z`��G"�gay2f�	"�>���3}	���Ɉz�A5$24�z�C���2%��O~�{go٢��<	W�ЭE*�lXe�I '���j��Ly�a�&���b��P,i:��4+�J�qvђ�Ȟ>Ķ�����]*�������x�JZ��ʀ*4�$B�P���j\��������)@��@*�.�N�ց�H~�=yf*Q:�9���Ș*VbtJv �F��lxFJ�q���f�2�v�H�	�<I#�.��k`��q��!�a{b�$:�̰@�ٴGfD�d��#��O�@C c�c�&(��En���]w��������f4�����ŏ@�����'	��f-Q.1`�3BER�K�]h.Oƀ�l�MG8Q��؀q>�U[��)`��M�щ� �e��K^�tU!�Dϰr��@�� =.¤���ɣa3�<s'ML7���":~��R����{�@>T�=��ֽ�n������?i��>V�x���UL1�Ĝ�A*`��i׾e:X���ŁaI���U|nT� k��Yf�*i#�5��I Z;����*�*B+8r��'�~���ʚ|o�0�_�4_n��'�L`e�Ԭ7�d���h �Qp�)O<9��с~�$��3���-�N�}�/ِ.ԲaP�E8h9�y��%�v�<9��"t�K0A�Y����I;!8V��y��ƀ$���}�����I�k�#��4K�K$D�P�!��>A����q��퍬L�� C_ RٶiX	�C8�]C2��T���s�+��IܚɅ�I�s�v�[&Y�< �fT�h�<Y��%[�V� �a�,D�x�EcN�L�$���!v�H�[H+�I!w�N�C3(]5Q?*�	�
�t10/��P�H&�"D�<�U��L��N�Pm�(��ン\����=���>�ՅЗU�@0�	��Fh&4��Ig�<�`BT�%�D,*��V�W.�� F_�<�%%��6�+�� uH~i�@�[؟�ac+J�� �|3�!	�HJP�d��:x��C�ꉶQ�$�T����p>�iɀC&������S�:,x��g�'y�0E�F���Yb��n��t�!p�i����N�y�@Q�x�v�Q�W�ٞēEj��	�u!�1��T>'�a����79����ǘ
�����!�y��3r:|�2D�(}C�(�ק��r������iy�g��ű H��ą=�Ψ2'���!��6jl����A�t��$zH�B�!�D���z][e���;��)a��H��!���u��4��ᖂ��S�bp!�FUf�Q'��&+�Lۅ�C_!򤐟'�L����d0P�5�X8<!�] Dj�ʑ_������u !�B$2�����Q�,��2�N�<!��.�Y�!�;�:X፛�h�!�ĕ3X)4A��:7�4�y����!�f�\liE@O����1�C�!��}��2���D.��5�W�+!��J(�8���ȋA宩�E^�!�Dŕ	2vŪ�/�1�d�����2!�Dƒ=����,E,���JȽ:�!��>fR�8a�	L�ne�D�ªY�!���51�����W�;�FT��	ء
�!��P�hߤ�r�N0M�E`��T�!�OP2���'�}+ }:��E�!�[���ό^ $��
�h!�U^4>`�Bg�����JQ�b!�d�<Y�(@[֫T�`���JFI�#X!�W�p�f�'�ǂ�u��E�D !��>/i�m�E��5z�ɸWH7	.!���?�<Pc$��Y��H2M!�䊔Jʹ-�6���
����P)�!�DԹS3rY�qǑ)6p�x�Iƛ�!�]�N��C9Dͨa u�մ%�!��+k-U�U�Y����i!�DԄQ���+4aɔ5�"u�1�p"O�X0�]�ys����ۯ1c
�s�"O�	��͘�ъ�j��	$X���YG"O4���ĵ1L�lkӃ"�@�õ"O\��G��;7�U�!Y�R� "Oȍ�'�����/F�G��ˢ"O������pΈ�*I��"O|���'h���0샙
��ڧ"O�hv�M�4�hk�+�n��0��"Op,�a�TƠ��<:�h��"O�����$8�&���ʛ 0�j�8�"O���@P�{�Yr���7Kv�=yp"O�LhE�ũ%�hD�'��So���"O�Q��So�D$���S�yrR=�"OЄ`F��WAfp�lZ�xm\ܹg"O�hbBRE_b���őV��uy�"OF�䠉#�`����)Ѣo!�$�4b
��O>3jԲ@MI�0�!��O�N�04-B+e.� ks�T8kF!��1dzDCa'fBx0� 8K!�dS�6^x�Y�)��f0Y4[6p�!�Ğ!�����)m�iR`�
��!���^�]���Hm�����PyR+�#9  ����@w���y�d��&�4�ADn��6�K��yBa�?F3P%C�]5��"��y��An�^�
�,Aɬ��%���y£U�
�z|IS`I)#�a�4�A�y��Qj&Q10H�Z.��@�,�y
� �,���܅
}��3J�L�!"O��!�d�+5���(�����ܨr"O``8��_�zX���ky��
�"O��E�0B����u{�.�y�H
L��IS�R	%���õC�9�y��-����!7�jp"���0=��P��b�'�HTE�j�*Y�,X=x��r
�'8ڍ �F��NU�1(q/�9)��d �{2��jy�O�Ow��K3�O4nj�U/Vu��#�y�<��.S�R�
�� 
��\5��)��v�<�'j�8�M� *�,]j^�Y�^r�<�r�(�ʠR`��H��V&n�<��lˢ[�.h��^�L!}�i�<�� ���J�Q�Q���bSB�i�<GX'B�l��löi�\ BHk�<�b�?$7�9a�c6	>�	�Dx�<	G���=�Gǘ;Of2Ѷ\�<�0lQZ���0�f�9;@pP���p�<q��o����T���G
��l�d�<4�	�E2���36�V):�`W\�<�F(�*?gN�R��,��a��Y�<�͆��̨ʠ�U&H<� �C�c�<�&�P�]�:�ӣ�O�7ql�; `�V�<��
�U�iY�	DC�����FX�<�G�ϕG�đp0Ĕ�]n>+�AZ�<Y�e[�y��C�g�Z��<��(�[�<!D�Y�Ҙ�F"�'<|���O�<Y&��-px����E**�u�Uo�<I򭛊a�R��q��F�LJgc�<��D�2@0`�	��H��Y�U�p�<�tMR�j�N=� l'�<�aa��i�<	�P�4��X���"J�|3��H�<����&M�X�Ã�[X��1��Rx�<�4@P�O�x����[*8�갎
t�<�f�@%y��UX��ӛ~b�hNq�<r�%�&�!�O�^M~yѳ�l�<�te�>0L�#ă�.p��b�d�<q��S�A:5	�M�:بdC�a�<y�]`��� �e��,j&jA�<�%�	���h���N�X��4(�e�<!2��~�j�AT$�"!&�DTc�<�HZ8�>�Y7� �`|���P�<	P�N8* � ���F���K!�M�<!�(ԯ$��ժ�,052�Y�2A�f�<�kݫ{���s���fy��E_�y�X�ue�1���D5"�XuP��'�y¤ɾiO4�Yb.�W�|(Q��y����W)�%J��y�Aᘚ�y��t �۠��sNPѭZ��yR��d��l�)Z�&kV�A6����y�3�BXi���'vq���[6�y���E;��20��D����cL�y����j&�	�U�Z�z��&����y"�Z;�`�82l� U���C�'�yĉ6 ��ɚ�"����l�&����yB-�\��58�-����j����y)�I�!��m�$$I7ˀ��y� �^��P�����x7h�0�y"�J�%(r��ؿy~M��C�y�+I_�d�d��R�}T���y�_9�iՍ�U�V<aS	�yrn�&#@�ъP��'Hf(��E�y��ɗ���	S�I~h<y��2�yB�a-DDKs����`�[`���y
� �$Y0k��2�d�C[��|���"O�����:}\0:b!�>33@��"O6h��G�<*V�� ��;5�5�"O�m�W���	`�̻� A@�����"O������ZߢeF���*]l�"O������Aq��E��<_D*�"O �wiq�a�p�<sb` ��"O`a��k֣?Tt�{���zi@�2"O�R�IΤo���K���%���W"Ob������gDz�D3�Z�K$"O�y��F�g&���N6�zUJd"O,p�7��`��AZ'��*;����"O��{p��%Q�V��ё i��p"O��q��?d�^���� b=̼�6"Op�1�_{�@0qG�M�5���y��Xͩ-�� `����yr�
6�� pM�1\�*�kwl���y"�T�J�m�L��T}`bu���y�̍,m���'H�L@bl�4�_�ymEҦ�s�臺,7hQ���ѱ�yr��atn9(�	��^Ix��3Ć��y����c4����W;����O���y���.��`��ti�w/���y� �#6�����]G�F����
�yrJ�(��XGT�%	Xd�aL�y"ᓀ
,�p:4)R�n��4�Q#��y�$�89�H��J'`jR\�f�D�y��^Pu�N���4
�Y��yr�)b�Bh��HΣ�lh��j�?�y����]�%W3��S4P&�yR%V� UB(	E�z"��%��y�/\�"w����z.��P�I��yң�<�|!+R�[~C��i�R�y�#ԿZ�8d��ʁ�v��]%ƣ�y�)�X�(���?wTp����yd�3�e(6n�m���P�A��y����0]�P���_�쬑4K*�y��A�F��MAGBN�_�°h#͞*�y��<Q���
Μ#�B��b�	��y�'G�@�\�E85��I'ʜ�y��ڀV[�qC$ڊ(�8�2�CȨ�y2j4��dR0��sn^���Q�y��ԑ�r蘐OY$k\�"u����y��$�X��c�B>K/��A�(�=�y`����@��]�<��1CŢ�yrK�?�L�t0^��A��yr�Ğ{�@A��k��C8��A��y��+~0����Y�8Wl�I�=�yr�
&��5��)69v��� ��y2E�^��4pJօ,�ܻD��y�Ҝ2���n�� R���b��yB쎋!9��I���1!r�|�C�%�yң�^�J���H"�Й@����y���?�P�j�&f��%��ybn�(�Fh� �O/���i�<�ybn��((�3w�&?\a'��)�yD��(,�i�%B1e:�}HƇ��y��B�~π�H�#?h�f(J!�:�y�Cߏ>q:���?�� $�J��yd�@z�h'H��p�k4�Y��yr���\X��<���I4DY��yR�O�s�b:A+҉2�E�V���yRaÔQlL�We�(*�̡ʅ�݅�y⁗�=+�����E���z����y
� ��2jÿ^Y:�A�A�g�m�""O������uv����p�H���"O Qy�d��b��³�.�4	"O!ږ�D�͒�쏩>��%� "O� I0M�
q|��u�H\�hE"O!�b^"� D�5Ws9��K2"O��ҖX�1N~����]>3b���"O���4Q�V����8p t�r�"O�H7	�q�𼪆�Ԧ���S"O���W&ڠ	��!�0�e�҈�"Ox�"��[�dݒ���k^�K���
�"O����e�9dz�q(�KC "��a�0"O��!&"Ԧ}�tJD���"O�x`��kr �@�G�@��p"O�����w��P �ƷЊ���"O$�'��9QK�9#g��/s-�i�U"O6��%��+B��pc��[�f���(�"O8���8�U���B�j��h�t"OlX�DF��$>A���$\����"O��11��o���j�.�*�"OB�����X�DpgI�# �Ț�"OlG�2H
���Cf�(p�'"Op<q��EeV��Ėw*��"O��z''#Z��cd�]b���"O��C�G� ����B�)Ce.�""O&���LF����[�0X,��"O�7`Q�is��C� �*{�p�@"O�u�4�M� Bx���G�pjޡ�"O�#J�:'~�1H8�P1A"OJ4X7�X%�8L��{06-p"OL� ��@t�� ���d,F9;�"O�� �I��@Y�!�2t�H}�e"O�Pc��]�h�� +��`�,H��"O6}y�͡}���虙J*�(x�"O`}J� 6@�؂S�G9d
�x�"O��r���G�Zk��"6�^upa"OZ��U�9pw�̩�K�'h~֩q&"O*���K�e�F��U���a�JIÆ"O�2�ո4�fyc	Ir�z0c�"O1�?���a�R'_Y��@�.D��XU�S#�I`��S�e�fI	`6D��s��V3���g�O�U�Z9���2D��86��4͜���ȇ� �2�9��=D���k��Y���S@�'�ީ0��;D��yU�vz��b�l�k���f�*D�� �(K�|`�$HB�c�pI�W�-D�ĸ�/^�4�	���?Z0�$`�%?D�<c�*9X�"�NEߨ1��!D��٧K�b`��c]�G���;D�L��G&�YY�F�%��qz�E;D� ��,�~/
��#��L��e��)%D�,���:
�pE��n\	n��LӔd%D�01�c[�8�N��-]����'`,D�x�S`�:�,u�7 ֛a3�1D������K����IՒgT ���#.D��� ��9U$L��O�3�]��/D�`{Ё҈T��01b����MY`�&D�4q�G�� �U��a�c�n�B�&!D��j'��1+��k��O,rJq�r�>D��C!�%t�!�!�	�m��u�b�<D����]�g����� ��=V�(D�t
�jY[gΩ�c,+��՘7�)D��xl2?,��TE��a��*O輨q�������@~�ɣ"O� R�Cb��n��b���<l���۰"O����mV�#'�9�P�:;�~Ef"O����F[�t8
��[�g�zeZ�"O�2����q�f	���MW��"O� jU�Ԥm0�m�2EqaQ"O��ZCb�L��@J�k&PI��"Ot�g�zz�D�|I� "OtY�`Ό�5����m�۰��!"O��)GgE4T�LP*�끍x"$ S�"O����C�0����FM58�ebP"O�8)�Я]?lL#BL�x�՛P"O"��@������!e���I!"O|� �h�:r�2aA�:z��Q�"O��ԊK-kT �A�܁^��X��"O�Yu,I�Z��,�e��9�R�Y�"O��i�ʑ�k0Qk�
ǭ�.���"O6�Q��7Ѡ(PV�C<zA��;U"O�٨�	AQl��M�R7��P"O��&$�!Q�Lc�k�a/�$ذ"O�P#2e�?�� ��AɏC�^�ц"O\� ��U=*K��yQoQ%}�<p�"O���M�-V9�L�]�H�f"Oؐ#�@M.@Z�s���m	���3"O���4�S)
��鐀��Uq�"Ot` ��O)���fg��3�P��"O����6����І�zeԨp�"O��*5`�%8&�i���G�X�h���"OAJ
��w��| � (;B���"O���7�Y�8-�/ҦwM��HR"O|�z�j�,�R0���G�BByHs"O2i�DL���8��KL�QY"P"ON�ŌΏ<.hP���B�z��r�"O��gV�i_B�ᒧT	m��w"O�� v*W/F&0e�b&�FRBP"OPt��¼@��B֬�t�ps�"O�P�eX��Ҁ���3&0�"Ox�J�ҹf|lM���!r��ಢ"O�����C3ဘ2�AW� �:�"OVbN&m��i1 ޜ�T��"O�U��X}g���`ѷ��( 0"Of�d \>[ZTݣ�`]���y��"O*j�L�8
��'@��yO��@ "Oz�Z�$ЎEc�t�#N�7J8�"O��qVښl	n4��Nv�a0o�;�y��D�Q� Z�c�^.89�F ��yR"���p�AփU\~���!�y���e90�Z��J��.�����y"Ā�%����F*֭t讐cT�
��yRX�o� ]�Bo��v��1��H�y���BG�A0���T��ܲ�Á��y�QI�f����F�X��(�Ȁ��y��ԑ<�jD��^`��"���:�y�$O*}�����z.3�yR���'@d3�
2z"�h�3��*�y��?^`�"��E�pY� ҅���y�l�%N"^��j�Xb����i6�Py��`U�-1pI61z���c�K�<�`��,c��� �P�x�����K�D�<��n�w���q����8ˠa�J ���H�\Qp�M�ɩ�a�>���U}���@�G��|A��
14Ǻ��&�O��P��'Q��1�m=�$2��<�VP� ��*}p��+Ɵ5<��D���YSBb(I����8����6�'�����H)�(˿+��I0	kD�ѵ�4���"ڇ�.l��9��<v4k���C�:���G�T?=��S�? ��sb"6ƎI����\���wZ�\8fl�4-�c�"}�+�+G�a�L�	����U(��<�b��6��O�>9S��b�>�5ꄬ|�jE�%#���ڈ)���)�x�=x$��1h.��sM��$�U�}2	F>�E�W$����%"c0xQ���+�I�c1zU����i�+Z��(��x`]��	K(L�I�f� Ĳ4�3�)�Ӗr�@��/�F���H̘?!�H���hTAϹ �ƈ�I�r�D��yJ?)0�ʦ�h;@C������1�J��hBq�*�'��DmR�0�0�!PȆ�R���J�7W�$Q�=i5��k>!�Z�f�`��վ\u���2�>^q��}��$��wD8!� �=h�e��kݑ��I�,z� �?�J��*�������:3QZ�M�E?a�ԕ����D�$41ڕ14�]�N��Y��CqD� ��C��c��|2�"�S��$BH��PG#�	O����p�+�0���S?6�WT��baȵb�����ڍ{�nB��ħ_r\�񢪉�Ze�Ta6J	�H�\�&�P��?EŴ0R�LO�u�m���X!)L��z�l_p��$��"|dC&(
�H­����$�T`��'.��K~�ɢd^(��p�C�|{�PX�!��.D�������`�O<����LE�S&\�ȧ�*MX~�`(4�BB�	�y9��#e~���+9>ꐩ"O\�(��@�t�9b�)e7�(�d"O�`qG&Ԑ�p`�/$��s"O�="���n��iQ�\:
�-B�"O���C���|��`� )ƷP�ҥ�q"O��	uaG*���C�mԔE����"Oh�p�]S"��̑��B�aS"O�L�o�yd��@̗�Q�e9P*O���G��Q4��g�̛xk��[�'����#L�FbA�f�h�'��8��ͭ4���x��X���'NnX��Ƙ-O�`i"E7`��h1�'FɑŐ"_�����^@��'�]��Ò/�� ��+�NfJ���'��f$׭#g�-Y� %B�8��'�jl)q�Y�%�x�Ԅ�4`�XQ�'���%o&9��#�8����'p�u��H��-J���S+]�8W����'`ιR5�,
�r���K�ZT�\;�'q�9!�d�1�f�#D�&R�P���'�
��@L�%Q����K.B���[�'i�(#���:�r���A/;�r}�
�'��"�m�53����N�/eZ<��'Or�ڇ��	~p�Q�@/[[��	�'������1��x;�J�~�IR	�'pv����|�´���֡p�����'Ӑ����Ja>\Z�C�
hi`��	�'KP�Z�'"����QS�g�X�R	�'��u�r�@�5��4�A�žj>z$J�'B���"'��5���9`�n�p�'����.͞V~�SN0�T��'G6�$��EQ�b3�ʹ ���'�J,�t
5>X�
 �O,޵#�'{���c˄Z}��g����t��'ՠ�Sbd�s��(s�EԷ���K%j����F�(�I�k@�q�ȓ(K�ñ�Ӳ\��`�r'�<gI� �ȓu�r+gC
�B�	QeIMe��\�$����7W,�@���"u�͇�o���Ig��DKXܳ���}-�|�ȓ�
ё�Ğ<Y�}{P��-��lDK&��7z��q�WK�)/���ȓ3���+,���|`�G	K�^n��ȓ�2�B�e�_��d0�aB$A���S�? ¨ ��U-8�va	!�E�,�@�"O(�a��I\V�8�q.H���<�g"O����fɫx�@M�q/əV��V"O�4��e�&?]0t8��� ����"Od�v��J�^�0��|�A��"OT��a,óA�,t��$�Zgh��"O����M�>9�\���3[b9�'"O4LZ�#7Nlx��Q(J�͢5"Onx�fJ,�D��SH>D��R�"O�R��^�n��bG�;?'��0�"O֩z�V�k��h��.g��AT"O�����:w�`�W5 h,ق"O����jP?�򅋑��L�:Q"OرQ!���7K�XP�IĪ	KLY2"O�Y��#A��F��V�=
IJ,��"O�K�,�A�`���N,d��"O�Q(@ _�i�����/ fA�x�"O��Su�ݵX�p� �NV>O&N(	�"O:Yx���)O������j "O��S��Żs���C�%D���"O<5j�L{�W�]�3�Qju���T!���*K�l��!&,5x�b�����!�D(/�B)�E1İ`ƥ� 9!�d6?�d5��D̞+v�J�E$]>!򄈑L����0#X�ʛ \!�䓜+�� �DR�_�2P��$dY!��=͖�#���9�؍	���:a�!���� ����*ׇۜ̓�5!�$�1�a�'� E�.Y�&iy1!�$��G���Č��x�ZM�r��1!�Ė=��h��K�t�x��$�2Pw!�$I�
0(�z���.9��Њ6�OZ�!�䋹'4� 8�G`���#q�W�M�!�D*?��<aRa� L��3�N�:X�!�}����֦A��V�x�c .�!��ڕ6|%��ː�c���I$�]�0d!�$[�)�v[�B !��H��!�!�� � �9��]�gs� � W5�!��ў.=@i��Ν<�HH��_�$�!���~pR�k<]�L4�À��5n!�n�	s�+̯B~Xm��\�!��Z�Rp�`��_�D ���$ �3�!��N�H���].��)A�x�!�dx5d�3� �%LP��u�;C{!�ܽC ,$���%�h3Ξ �!�$�{~`�P��?����b`��!��M#>.��#d^H��1W��=S�!�$��W�,�)
���	DJ��B/!��:lH<�W�1R�TBUc�6w!򄞟a}R�'ǁ7����	36�!�8wu��L��I,싷��5Q!�d��8ϞY�&�6.2�xa�fO
B!�DV'd-����퉇$�l��08�!�d	"�͘��A�xEb� �!�܆=��Ai�	N6<	��CL�?�!�$��rp� �Rc���ZE+6�!��ZC��Plϱd�H,���ȿ[�!��G�|��@�ce�*0¨�ʳIP#<�!�d�Q�I��B�'،�i��RF�!�$N4S�:=�C<B��5Ӂ/�!��۵r8�tJߐ�~0���ċ�!�P<i䞔zq/I�Bw���a�V-hl!�D��?���ƨP�v[�9�4�͒V!�ć�I4DІJB?~��DJ=<!�� ��B�]1)�R!� (0 �pc"Od�#��&/��bfD�O���:�"O΁�#!�>\\�[���4{\�<@"O����#iB�u$)s�xi�"OaKe	�a5��X�c�4���(�"O�DX!��1�fؘP�֡)H�%��"O���W�҄�H����?#/��2"O�(� H	Xް����,��q�"O��r��ɿk��@aV�'΍��"O����Q2Z-$5Z�O���U��"O� Η;HC��r��h�3"OtiR�� QS��sw 	z�ڍ�"OtI����4L����A��n�B��a"O��r��R����N�<I����"O^`Љ\�>��]�G�O37[�"O΅�VD�"������0.���"Od�3&�0GI�B$�v"ju��"Of�B��E�(�R�>s��d"O����K�8��$ڦ���B�j}�3"OIs��Ɔ*Z�j���$�H�"O�x�gCY5jvu�b�ӝ`��DBQ"OTp ��#T�*��f��~�)#�"Oh�2�
E�u�v42�T>Pl��"O��ci�3V�B�W
r^�[%"O|��
�i$>�
��\#E�� "O
QQɃ�y�z(�-ǕnK�Q[5"O���ʎt3ڠ��n�����Ȣ"O�����Ϝ8�T(����1���"OZ����͖R�8�j0�R�l���0"ON$�!��C\�=��N:�05�0"O&��`̅�;P]�r-/�
�H"Ol
��I q�n���mܢ>��A�"O:��T
���b�{��U�<��a��"O�D�(Ç<^>@Q���)RgbxK�"ONQ5M_3���K�#9~K����"O 4�G�WC������-����"O`��N%|��MQ禄� ��@�e"O�ݣ7�ۧ}Y�����Y���@�"O���!.�2%7�5ꡩ��1�f"O��82�;E�]IC�&MJR��4"O&�5IS�"����!R>��"O`���A��C���0���i��V"OęYb`�8l���)��C"O�PT�H)8�>}�F*цs��4�#"O��9`�H�z���r�I�I��L�"O���C� %�����O?�nIJ�"O�iJ���wv���W�P���僅"Oʰ��W�5&D,���3~Ě�"O@��C��}02���֙*Qh�!G"O�I� U�S�R�k�%cH��CD"O�@�"gZ.Qga(�(�G^J�&"O�q�H�"M� ��J+,�X�U"O~l@f��eu*P�c��<�A#@"O�%oR�1,&�[�QM�4,�r"O4 (Q.	;��y�,וzu��P�"On��ËW�Y��3���-x�h�v"O����	Ԟ_�&��(�;.��РE"O�T��Lӟn0ZY9���80"Ov�Ȱd�0�Ҽ�`�Y|��"O�� �%U�FR(��R������"O�uIB�ϟ688�6/A��E��"O^�a�hN����4Nèv�����"O�Aێ_��T��n'�0e1�"O�ڱe�/�R��nZ�6�"�a"O� @��uf��u�`��Mכ|��ы�"O��P�ζ\;�7ď�,�|)b:D�����3�L��sℝNl!��_3��yB�!E ox0Ȓ�jǭ�!�D�SU�����Q�]��Ҫ�/\�!�D�.X�[х�$G@a�����!�ʯl/��0E�?�a�'��N!���b�����B�_#8��׾A=!�Đ%Z��L�s�����]0;!��\43���D'逐�$h� f!!�dV6
�s�
�$T(����Bt!��ޮT��l��e����Nڃ"Y!�ď�:���T`@ܪ�n
�J;!�$��l�h���݀>L��U�Bw$!�Ę7n���1FW.Y���p��ҁIC!��˵)m\�h5��@#FI�H�!� �mHP�I0n׭�8�p�� �c�!�䄙�.�Qt"WEz"E���=~�!���:-xjy*��N!@	p ㄋ��!����?+�E���c�T�ȗ�R
"�!��BPn���[3���e�Jys!�$�; U��#��y�*i�@�oc!��&VC��+��;s�\�7 � y�!��\.i����g��CV�])��$�!�DЅI� @  ��        �  e   �+  r6  {A  �K  U  m`  �h  �n  Ju  �{  ف  �  ^�  ��  �  #�  g�  ��  �  1�  t�  ��   �  ��  ��  ��  �  ��  
�  M�  	  H �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b��<�ߓ#d��t	H*"F��9S�U�ȓO�����0U���6�*hU��zЀ�L^4�z�׈�/Ae��?�-O,�=�Q�A�
�b��҆��Й�I���yR��)'��S��ı>v&�c �&�y��ܞߌ )0Ֆh�]�G	$�hOb��I!k��̹�0Q�A��
��u"Ovm�� ��q��&@?1�,B!�'�ў��s�\�=����M�2��l�$g1D�L��םC���@#
\��0�$G;��hO�Ӕ���N�\�jpT���{-�C�	�3Ľac�tX<1צ;f�c����I	)��p�C�w�l�:�ʄWg�B� /-��b]�c$���bD=_��ʓ�0?	�#])m̕H��S��20Q�X�<1a�D9�%���ѽipfH�Ѩ�<���9{���2���2r&�#��G2��''`"=��g�����P2�Q�eB�yrGäw7��b��"A��$��Φ�yB��$����F��h�t,�=g��!C�NP37$6Ʌ�M����;�|�3E�s�4$��W�<9@됻0� �S�%@�=>��g�Wx��FxR�
r���K�w�X}���m�J��\؟�k�U�W�� �$!��J$D�X5�f��x%�)�T�Jtf�4Lڴ����
�\>@�ȓ<,�dKNO*�$Kr�ֳUY(�'�<!���#X�j�K2��4W:�"P�Y�\7�C�7*M���]7���$��,m�B�I6�$QC��N�s�ڄ
�+G�r	tB�)� Nu���\.N��cHF�y��![�"OV��E�R6L��-�!�� �"O�HX����mZ%/�R4��P`"Oֽ
w��4B������~�x��D�>I���P&P��4SC�@�l��ɪf��*�~���OD�ԨKX	�U P��fV� g]j�<��&L�8Y�� G����f�f�<)@��C��г�+�����rN�j�' �y/�9&ߠ��e��2EE��pv�����e��(����Ej�;Z̹�g�N��-d"O� 9P�+V�d�B��P�6v�K%�'X�R��?�"(��gć[G�m�@C��S�!�O��кצ�c+�|XG�� ��
����Bu�ӺK�yBʗ)`ZD|�b��	�Ą����&��ޟ �?�B�Hի-�9�%K�:��/�)���O<,��I�:�n�[f��8J2��L'd�(M$� nZN*��O����V=Z�� 3ac��,�Ex�MN*	9����'��5@��j�D�FA���y�g˼<q��d�(61O"�P��7?c�3U%�,�:'"Oj�XW�0Z��*掃%ub�Xƞ|¼ii��>���lF�<Y��"]�9����:D���W��21��Z��s\�A{���O<�Iʦu�'�axfP�P����)D+3�>�16H�y2�	X�1r$ֳ&VJH:�/��y����h��,M���)�y�0������?�2��f���y�ߝRtn�I���8;�i�(��y��T=���C�*a�TrT��y�`������֏��5���rb�N1�O*U��IEh:��g��6:���J�,h�*C�	� g�()Ar�����EndjB�I�Bf|��� �&	�����ך@�
C�ɲq���M׮T~�l�!��L��B�	a�Ŋg�ɻ~��4�lQ�)��O��=�}
qD
�#LRHC��JL����HJ�<��-�C��@���jG�]ҁ�QH�<ٓ� ��P�{c��D��R�-�G�<�J!>�4�槛-l��	�!�K�<�tj����΃,y��Q1l�M����?wN��d~��4G_(����B�r�'�ўʧyN���@f��S��Qzw^Ѡ<��%�b�:3�K�m[�E��O�V	�ȓX�֨k3KFQ	z������K����?!�Z+ta�aJ��1hN؋m/�h��!x<5�D�Y�O���z�fճJ���ow؞�&�x����5^�J��&�_�0g|q�s�%D� �S	 �+D�	�E�H'�R9�R�!�~����a]�	ʢ	�%ސ�����5Y߉'(ўb?��6j_�>(N8�����lU@�H:D��(��� �|� �ʧ�pX�� 5D�����ҿ]�j�(�ɌQ����`4D����d��Z��Y��	A�>����0D�г���o�ȁBB��6� V�,�����'�B���U�X�X8�s'ʡ�m�ȓzp�L饆%WLJ� t�Z�a���Dy��#�S��G����E��E��I($�W��y�B���6�J`퐁"
���� �y���(I5�x�c֊/B��跥�"��It���O�ȫ�-O%O�nD�q���4t�O,���8d:,
�8Hwj�q��Ì4�!򤐘�6�BƁ=`��d�X��a|=O>�+n���ЁR�MI|�YR��A�*ғStax�jПm�UXM("��p�+ğ�'*�I�<��I\�1|dݑwo	�%,����+�!�� n@����� x����
&'N� �]��'�`��Id�N��U �u��i���O�~C��(��a#4 ��]��"J��	ey"�Il�ɋo7pI
Fc��mz�$A!#��B䉡[�h�rw��&�h�BŅ:��B䉋r4�3U��.���ǹłC�	!%5X�5�9�@���#w42C�	>?H�a��f�4�X��#p��=q�A[r�kS"�}��
�%�N�)�ȓ:�օ1T-X�ǀ �1���P&��'��}䘶ZN@������vqp�L2�O�#*QG
-� �Ɓƺ`/B�7�:T�<
 �� �H�X5O� ~\�Dh�0D��j��'^�f��(9=&�x�)b��G{��)�)��D�46Ba��E�qO6���y��i�,ɚv�pmq��{��Jx�$�vlZ� ȍ`��0Wl\A��/���E{���^�G�ڬK�dZ;��H�4&k ���S�t���aD�9F�t��׊ۀ0v�$�dE{����D�'d$\ui_�'"��-F�'�ўb>�C��<X��[��ٽ�`H��*�	az��E�f�牜�Qg�I���$�O�\�剾)��t0D�����H.O8���Φ1�6�� �x�#!��RA�E��-�HOh�G{�w>4�����9J
���!�X��
���yb;an���t�K�I�(� m��y�d�>X`�8C��^BB������y�J�E���5�ڟ��� �.^r�r��%�)��t1T�X�s�ڱ��� �;z�
�(;D�L�ЈJ;8d2�p�Y(�f��w&y���<�O�$�$�V;:�H�u�L�(�!���'��+�l�`hS+ �t��#*Иu	����	H≚(��av��<U����D�?VC�ɋ��q�	j"���<E�B��$%��P�1aJ5#�>ɀbퟴZE�B�� �p�C��
}�([?��B�ɴuKڠ��-�	g��P���%7@C䉔�V�?�a M�_W,DX�'�6ٙ��6�����Ȏe�0`3	�'/��0n�=?�Z�C��N(�vt��'��	�k�0s�X���W�QJX��'@d��i��[����a�ӰB�V��'���uG�9\t�L+B.�)Z�ŀ�'m�a�4� �<Yq�B�<&��M!
�'2L��Y$w Q ��I��&��'�v�$l��*�����':�i���x�� ����\�@8�
�'r���Ђ\>$����f��Q���
�''�H��	H�Q���a�� ;
�'ږ��m̀Uk��2�ǒYl(I	�'�8��*��0<����B:he����'т`�V��d>�e���([֘�'Kl��c���ZL�`c`@�9vG����'2
���K��L��!��8K�'X.�c,�pF�%�e� ���q�'&�#O&��lJ`�D�~0�AJ
�'��X���<8�FH��Y���
�':"$J1�O�}{$9�R
�+m,��'7D��bM�'�*b��[Y���'�D�J�a@�8x�؂�کNe�=@�'�n1�Ԇ� qx���F� Hr��A�'��q�/�*x�T�Z�Uz���'�����kf)q푴<�f,��'�4X���;�����\#7J��
��� ���n�?>�H	�J�as@Y(�"O�arA�\�,&yc��Xб�"O�I�h��+�pi�"�l~Z�H�"OԜCgi�9��pE��0~Ab�"O�3��^t�1葊�.p����'�b�'���'E��'VB�'/�'�:��Ga�0i3r0y��]<Y��C�'3��'���'A�'��'t��'f6YRV��+�)a�)N���k��'��'�r�'p"�'w2�'Z2�'�����G0F�8tLݨn� ��'$��'�2�'S�'r��'�B�'ZPK[i��dp#�P	REFTȟ���ߟ�����ޟ��	П8�I˟$H��Η�q�E�V� ��P��h�ȟ�����H�I���ß�����	ğ<�e�V�����`� �h��#��͟d��֟�������	�X�I�d�	ڟ���Y�d#v�Ic�ZY��Xş��I�t�IğL�	��Ɵ���ȟt��Xg"���� O�PL3#�ɟ��	����Iɟ�����������I��p�E�H�1�0�~EPq(���H��ٟ��	şp��������l�I��p3Dឿ/�<�k#�W�ke�u+fW�����h�	����	�0����\����<�'��J�:�RSX�Z��aC������I�(�I����џ����H�I�4I��8J�
�8*I���Y3f�Οp�	֟��	ݟ��I�l���M���?����g��=�g+�-8k6��$p��ퟨ�����Ĉ����@&��9�2�Z?1�B����f�eɛ��4���c��m�ቚ�)��ݸ�G­+p�5�$�֦��7Ĵt�uE%?��n�-I3ⰰ0�,�$a��H��� h[�5qp1R �6��'p2R�$E���ˠ!`�at��3.*V���׍a�.6ʾj�1O��?y�����șr�R]�T	H�\V�� � دy�½i��<%?y�������6+*�a���WI��싶+|uD��0�v��lǿj�2tD{�O���ѿ#d�1R����C ʖ��y�Q��&�L�ߴ:�:��<��	$�6\�/jFvER�lD���'�l��?�ߴ�yB[��X��*�2}��i�<z���2?!��	x=<�P�/CşR;0�q�OE3�?y�Ú�wg�Z7
�.XlD�b�2��D�<��S��y���9Ң�Q����K` ��́�y�	c�v�:S���Pݴ����4��T�P=9�iJJJĠ"!
��~��'R���'s�͢������<#��2/���BG+"Ќ���Ա�޼OS� By�*E��M�plμ>�e�A����:�J �޻��K�MT�8�DRtM��Eu�}�@��o��<��E;{�l���Ҍ;8�Q[V��%�xl�� !g1pu�Ba�?q���y��O�|�*V��A�M�F��TRq-L�z�x�1+� Y��y�D�J"����Z�0tM�R����.K�f�$���͏'A\`a�5DK3�d�I �41����=nW�$���E�
d��SȄ1m�C�FN'�4t	��
:-� ��O͒n�����Z.5dr�1�����&�0ծ`�ӂ�֩�M���?!��zC������W}�T� �Ԣ��}�Sd�2ʓ@(�(Ex�O��S$L����rX���I�$Ll(
f)Cڴ�?i���?a�'K�'�`J�j �x �O�>p$�W�̃g�7�ՙ���3�	̟�hïJ�'�x���1C�r��򏈒�M����?!��B[-����?�.������I�A��qE��#�� H0��&��'�h���9��O�D�O2��n¤�� a�a80��@��A�I�� yK<����?K>�1y4^�_8��㛁8��@mj}�����'���'��_����F�%0h��!n!^͸ToM��y�}R�'~�'2�ɭD���E�ٿlF����,G�kg!�I��X�Iޟ���џ�����������?Or��%		�J3p�*�Y��M����?)����?!��$9s� ���7�T�,@� U�	e���ν>���?������J�ҭ&>�*� ��9;Hp�.E0PWtQ0cě6�M�����$U2;%�O�*�R?2�4Ez4��5�Z��1�i!r�'���'$Z<Jt�'e��'i��O�u�@),�~��U<(�^�+��#��O.���"w��r�T?���iUfM��	X�W<e���}Ӟ˓��	�Թi(��'�?���)��� )��1ciߵ!RZ����'�6ͳ<�6�TL���O���v�' n���/�E��}{�4,�j����?+O��	�<1+O*`��GR�t�ȹ"5�$[��-��Ʀ�ʵֆ([�b�"|���TU�)�T�\1㘸�e�U��$�i�B�'��H�#�X6��O����O��D�O��G�<`HV@�7~��uN��4�v�'�2�]�_TDઘ�������$�O����+$X���ϛXx�-P7��O��!d�ۦ�������	�\b��:��%#bElTP�Ȑ�ba�
l�7��3\���?O>�D�O4���O4���O��ݪ bn�ӗ$�Bnb 9�G�+Or�1��Y�������	֟|k��pʓ�?�"mE"0e`l����#��=�d�g]�E��?A��?����?�/O���ÄW��H�NxY2���;Ϙ�� �k�
��?�.O��O6�$(Zj�$��#�R�H�'	�K��l��`|��3oi�V�d�O����O�˓���U?���
�*��Ai]!W	8��!��~��4!ߴ�?�,O���O���VtM���O��$D1,�*\:���v6�T	���-n�L;���O����<ɕ��~��џ�I�?�T��o7����ō�)rY#C�ʍ����O6���O4�*5;OX��6���π �IcNpD��#��m���7�i-�0Q��@�4�?)���?q�'}��i��Ab���MPv�8u*;Um:��$hsӎ�$�O�H��;O�OH�>=�"˔����k���Wfx�D�rӎ�H�	ݦ5��۟���?���O��E��0ck��c��yc.��H�x8Ac�iP�I��'lY�<����Rm��fN���Ж�d��ڥ�iJB�'�B�O�^C�7m�O��d�O
�d�O���0D`��%K�0�� K�#r���'�B����I����I���$�Oh��K�1��A!@F�0�0�6�Z֦��	D(�ٴ�?���?��m:��w?q���\ x������TSM7��T}�(�/�y�X���������x�I	ִ�h!*T�_� P��͌*v�8�(��4�M��?��?�R?u�'E�B��\��7��)ݓd��3�q�'e2�'�R�'�BV>ipR$ͻ�M��$AV��*�+t����G��;{�F�'���'��'+�	��{V�z>�𐩁/8J�1��<E>Lm*Q( �M����?���?	DY?Hba��M����?�g�/d��ٷ����q��K�R���'�B�'��	��i�bi>��Ii?9@��2y�^u�#퇜F���:�����}�������ן�f�5�Ms��?���r����7}>i:�Ǎ9y_�%�t�X̛��'8��矌w%u>���|y��M����H�еoD�E���9�����IɟX��n�M��?i��"���?�_
�"�.�y��L��O	⠴p�O��DU�AH�$%�4�H�O����ͅ7A�D����+��Aڴjhl���iw�'L��O��d�'�R�'�u ��$
�!Ќ@0;��2��d�`�`�O��$�<ͧ��'�?��W.b�"��J��#��8��.�#\��f�'B2�'�"y�?���O�����(��M�Qh!�/I38(xz�0�	�x�b�X�Iş���6JV�� ��zD���Ȝx��yq�4�?��hDU3�'��'�ɧ5V Fy�8�0�`��e���aϠ�����3�1O���O(��<I���HL!C^� ���n���][��x��'���|�Q�h����`N�� ��������:�c�L���(�	myr�>mj�����Z�-��%;uę%	���?a������3��'"�*��c!a�A% W�3լ��?��?�.O�e;�ly��J�5#��Y5]Q�F�W���ٴ�?�O>�+OHiҐ�Q��Y�*P�{^�� c� ����'�b_�`2��1��'�?!�'���c��
�v,C��R�ɶ��6�x�P�����(�S��%V�2q��z�HU�#��r���M�.O��`��N릩x��x�D�~��'�TU�2(S�2������X��Q�4��H��b?1�1DD;9f�4S@Ĳ z之��q�0iQ��ئ���ޟ �	�?�	K<i�2"��,�y����á�-6KHiQ��in>u����ß!أ�m�R�N�8{x,�����M���?��I�>���x2�'��O�Q!%��?!�:yc\H[�a����P�gN1O��D�O����A&ސ���i����ݯC�oZ۟�Bk����?����Ǝ�"F�)�Ч['b�,:R��o}G���'�R�'�"P� �W�:'��̋���'B�ި[�W�$�hJ<A��?H>I/O*�� ��?*V$֊ٝ(�L̓O�$!�1O���O��D�<Ѳ�?e��X�U`6@aD`�Yt��	��޺G��I���I@�	bycՓ��dE4o�<��'�I�Cĉcƻ6��'���'�U�(Ё���ħo��<k��قt��xR�ȆN�:����i��|B[��:��3�ɭ)/��%�V2<��0k���6��Ot�$�<af�c�O��O0�$ŗ�_Ix���ʋ�aY��� �)�d�<��Fi������E���5���Wj��:TlݳS>��X�� ��Mk�S?����?y*�O:��R�D�F����$<R���
v�iZ�	�R&#<�~�q��}�^܂�S��]�4�W��5��	�?�M��?�����q�x��'1ؘ� b�`�$�*Q��G���HA.x�H̚E�)�'�?�1�"qFhH��P/1l��v�2A��'H��'���+fO(���OH�ĺ��s˙:�ZrKB�Ԥ:�($�	l=��П����\�����r�L�I���`f��2�lL��8�MK��"�"�t�x��'�"�|ZcN��b�cT U?�]�RbC�O�-��O،���"���OZ���O��&J)�盼a3Q�B�[ (�u��F�v}�'�'��'�	+lߞ��%�-/�|�!lB�@�
�w,,�I����Iܟܖ'��S�~>��r�C�3IaB��P��X%�2��O�O.ʓuD��'�AK��H2`��U�s�I3`��O��d�O.��<)shؾ~v�Oђh���bj\j ��A�v��'�l�B�'�d�<Ѧ��S�D�Jѓp�F�F�V�hUG2W��o����jy�/��eM��r����
���!��7n�������3%�TD�	Ay"hS7�O�i�+
0\u��!ω6
���&�-#���o�֟��	,�����4�?�*�8���m~")6Z`0�w�V9p���T�V �M�.O�����)���H�d�Le�|���(S�'�>6M�_�:�mZ��4���X�S5���?���r��Y�5��&u��y��A�w�ƥV��O��$�O@� �BFa��Z���%d6�u�"�i���'�B.N+)�O���Ot��f���p�N?h�V���	�^|�>Y�Nh̓�?����?�#@���$����/�"�Z�#�V�'���Yr�3���O����O���k�/@�:�T��f쏧P�:�Bg%�y}BdI4��'B�'=�Q��Ҁ�'`ĠyĦYX1T�A���Q�H<1��?�K>9+O"0�S`\�j�b8���%�����rT1O����O���<�S*�{�Ɏ2H����+�+W�1�L�[�	�����I�I@y��؇��d@E`�]���5TY� B!LH�9Z�Iß�����ȕ'� �D+�)rb�
�(��5N�����'YB�mZ̟$&� �'���}��[XX�A�V)]5�d��:�M��?!-O��a3��A����S 8QYtG�Fnj��g�ŚX�$O�ʓ_���Fx��Н���=1�r�d�4Op��ҿi��	�hB��Aش6��S؟p�����B<�� �B�^��M!�aՂ(훖W��q!�S�'Ny�H@toGo���:( 6+�7�ޏ:���l�� ��ğd������?ɂg�q����
9T���iԮp��&�+�O>�	7� ���L�\e�bN�p��ܡݴ�?����?�a
P�_��'���'��d�4��j�5U%�u0��5v��O�c��d�OH���OB�[DF��N�D��"��!e,�bd!Tܦ���!9�Wp��?�H>�� �fxx��-����KŨj����'��$Z�y"�'���'+�ɯ>�����hFp���p��!H&���U/Z���'�R�|bX����N��\\�p�(%z8��֒*�@b�8��ޟ���ey2�+]���=/[�����߯}D����� �JO���-�D�<��@L}�ǽl��A-[2q�BE� �K4���O��$�O�˓r�nY��d/[�1���yFǘ����#���.�7��O��O�����>��Ƈ#��qz%.H� :Z�qa#��)�	�� �'Ryy׍#���O6���f�91���~e|�i��_�:�5%���'3 ����T?]BV-�4a|X`8��F6�~��R�iӨ˓T|�»i,��'�?���L���Fɞ��f��R���Y2�6�<A���u���O$Ræ
2��\�@�^{j��ߴ	hu�iV��'���Ok�O��d�I�\@hI�i��ً捑-t9��oZ$@#<E���'.W�F��L��������A�bp�����OT���;��&����ǟ�[�J�[�+C�R����@�-N���>9�o�Y̓�?	���?!��FG���e�	n䀔� �ԱX���'�p�JA�<���O`��&���"���F�)A��-b`��t����T�|"�<�	����Iğ��'w�X�A�S,�]�`ā���)�""�ROp���O�Or˓j3�`R�dL�'
L�(��oX��+s�{��?I���?�(O��0���|���N���%a��U&�����L}�'��|^��*�!�>A@��Y����N�gr,M�q��K}��'FR�'�ɀd�`|�I|� ��`�̕ ��F 5����	Q�l���'$�'��	�L�c�8Y��ǈ0� Q��"�^MZ�/u�d���O4ʓ+�R�ד�D�'[���Ƕx�r�M��Z�� K�G�O��@�V\Fx��p�@��	�j����9H��X�Q�i	�	�ֱH޴%����`�9��d��O�� ���G'�P���	H
��Y�Ը`�#�S�Ys:��ՅJrx��%�$n:R l��%9����4�?���?��'C�'(��#D�����]!���):!| 6M�Zk���3��ϟDK���W\Ո!D;�-!�(@��M���?���k�9(��xR�'fR�'V\�*�|��� ѱK"Dxa�>�	63�Lb��I��I�<R��d�<]D(O�%/�l-�ݴ�?�f�F�}��'�R�'�bY���#���R����qZ2�	eȅN�D�Xt�<���?!������t¹����7W��!p�F�-`�!�'Ck�I��D�I�'��'q`$[�#��T�|��4S�4�:|kA����'���'&B]�0�sKDQb�c��ZNQ�կDYq�D�"F�V}R�'E�|BZ�@�5��[?�䬎"P��  G	�HL���BO}�'��'�	)l�,%?�񠧚~a"��%�)N/D��$A��M�������d-WT�@����<1B�IU�%Z��"im�|���O��P�l���'�?���45�#��>r�\������ꕸt�x2�' "c¥mb�|��\�v"5��]ٱe��-��k��i�剂_��0�ߴ��ßx�����4A}�{ �۳;v�3��K��6�'�W�x�R�|B�� # Dٰ�S.~� ���%C�����%��7M�O��D�OJ�	�r�	ğ�H�~�x�����6"̝Z���M�s�]S�����DQ?qڠA�l �yQF*Ů͂Oirmm�џ�	ȟ�x��L���?����~�G�Yx�y��G�?���;0�F.�M�H>�T,]�<�O ��'��A�B�����R�ȸ���[X �7-�OX�1���Y��П4�IY�i�1�ǀ�OI�� �sؐM*f�>��؛�?�.O��O6��<AF� �]�׆�i  6I�-�����In�'Y�'�'X�'��<b�$�i��ظ3R�$*�:�M�.|I"^�T�I���xyr�M4T32�ӫ~��Y�hޭ6Q02p�������?������?���SW^���C�����]�-pL�Sȏ�yrH�uT�t�	ȟl�	my�	�q���x�Ȉ a`�e��q���ぉ��	h�Iퟘ��@�b�8�U���N�*L:r(J�x��Q�AwӮ���O�@P�j����'��T�S%-7�e�NI�Pll��CU6O��$�O���	U*E��Z^�tu��Q��}]n�Pyr�1aN�6��e�D�'C�d�/? F_�q�	��i\>]�@�Aȕ��������F)�ܟ�&�b?p6*�K�. !/u mq�yӀ�+�i
Ŧa�	ݟL�	�?��H<���R�� ;��S48�x�AZr���$�i|8a��'�ɧ�2�DN0M�Ra T��.[j2�1@Q�@mZ��4��ǟ"S������?)��~�!�����^K���g����'��x�Ғ|��'�B�'� ,Ir�;M
P�:�]�2���y4�x����Q/lH��'������ %���V]D*!|)�5�BoǦDj��E��yR����D�OP���O�˓\�H!N 1�R,xƠA��A!'ԃ8�'���'a�'���'�M��ҍ&a*���\� �f0c��RY2����U�2�^�{r��Zf�-�L~��
2��,
NO��"ք�P�<� ��@j�O�u�� �!�eܓdK����-R9$�8,��œ�u|�3���
u���"�8��A\�8�zE؀��9!U�!)caC�u,
�
ܡ5a���xdPs�	�<��$�U,�P>��aD?s�l��e�`��@:K7�TJZ�Kܜ�V�>z��� 4�Ù-0T'*�1W�2J��&}L����C�O�*��؈U����L <3@��G�ON�$��Z����0��i8N�K.Ѧ�qZw��]�R>]AF�.���:�N�4̠���i-}rK��D�s����E1��i�ם� �|�mi��"��,��U��mݨT�x��O��b�'�������FK�!-�ؽ���:�L��dA)D�$+v,Lذpa�j�?6 ���%O�Ez�͓b2쉄L�DU�d���=�>7�O����O2����%�*���Oj�$�O�nG�_���h��Փ{X��p��ɕ?|����l@�_�����45���1��N�g�I9rF��fތdvXQF�_*0y�)d����uI*=;n�#�h�
�q�2]`d\�\;C�f����,체�a�]�M��\�|y���O�I���[&�����b��6_q��AO;D����ҍJ� z�b_1�0:m7?��	"�M������'`���"�f3�du0�b�q��=����pb��d�O`��O���;�?�����&37��bq�C��}�BNU=I9�Xz�eU�!�� �M����y��X�@W���"O2c�4t��nŸ*���C���4	N�u��-��y��4d��Т�l[��!�g�7���C��?i���!�Ɍ% ��K�bֿO}��Q�[f�C��7a8��#k�&?fd�EM��b���O�ʓ0ر��S����L�Yu'�0�40���W)C�̀��՟����Bǟ��	�|ڇ��#n̙�$5t��Ċ*S&*��.E�y�h��֪�+(�xbmG' �:�f�8^bl��A�Ԑx:�D�C�G}5�܋r�X�"Z"��僼]�\Ey�%ʕ�?�����D�K� ��N�Z��ܪ�M�{�1O���$H���t�W�(f��,P��8E!�ė즥�W �J���)w�_Wti�C�b���'A��f �>9���Ɉ� H�[2N40(�u�6;l᳴��p
���OL-��$%}����DW�|Y�T>��O���Rd�(-��C�Ӛ.��QYH�(��둼}4Ѣ�d��&6��ҏI�(�#0�?�YQ$�2��Q5ˋ�Ybm�҈"}�
���?�d�i'^"}��'Y�*Q@"�����N�('� h8�'@ِ���5��9�'�/\b�i)Ó+j��@a!'ѯT�tK�b4c�p�@�M���?�L��#��!�?)��?A�(�n��1$��HJ��б��ſʔ틐QQyb[,���R��L>)M��f\���T�iQ&!hȱ4p�b\�t�W�:�q��'��M��U{�;u�N,w�B5���~�N�'vf�C�S�矐�I�8s���w du�D��eǴ�i"�N{h<��D�7]���E�a�����O~�:�S�dX��8�dPo�N�Ȁ�Ùp�ؠ��Ŋ����Oʟ��Iߟ��I��uG�',�1��x�Tf�15@t�pB�\� 5"��  ��X��H>'v@R�+:$�ax�@˟y��QjB+Ψ'�xT��]�͛��?�:{r��!ư���<ˈO�qⷠ�C$ �B�PC�$����ourir�vM&�����L�?���8`͘��1�M�7g����w�<ag"�[�(�i%��$[�\��H̓=���'���*W�U�ش�?���9�L5���7���P���i~�����?�Q���?������D�&k~\�����(�8���i$�[���0��)dP�z���Z�W��d�{9 �2�L��{쾍i�g�@s�TeA�S'"���k��o��D|B(�?I���� �!�� ��@��d V�D�!3O����O0�"|"Ån��if@V�"�D���NK<�4�i���䟖W#�3c��<gn�4[�'~�I�>t��)ڴ�?�����IHT���d�<���#҅��0V`�lC�h&����O���p��'���t�$׺d
�|�(��	�'[SB�P[t���а�>��!��9ȜA�pEK�1�F�"1̅I��%���Sf��LD��È&&��<�O��:R�'�\7M�O��$'���O�#�,R�9z�e�p��� J�e�O*���Ol�/<O���0��=jћ�-�5A��s�'2�#=� ��q1J5��lM8u�V<X�BS�Z���'�r�'��9i0�����'��'�֝�f�t�c�ɛf��b�㉶��ʥ&
�D����4sJ�33m�y�'EJF�z��`���@�	�rE$2��8z�2U��,��0q� �BM�t�x	�v�R�n��>�:T/�M��$Ԕ2�T��u��{�ƹ�ōL*ي)m����E.n������?!��7AE�׈T�k+�|��Gĳ�̼�	�'\�#%��<0R��d�"0��OڅGz��O�rZ�tJcb�6}/&5�dЪZ<T§-&!�pq*��П(�	�� �	��u��'��8�"�S�
ѐg�Nͳ�P�]\M��'��	4)ش8���{C�Y�� xB�܋�(On1��+X�4b��P�gB��A$'���:�� ��m�� ĦyʗBZ�TIQ��R���k�c��ZjB�d9��S�S$���]��ݑڴ��'a�b?I eR>M����h�15S ��@!D��"Q-��ݖ�⥇0D���/9��4�M����]�(o�y�'�"�4z���pfLc4�;�㝜m��'�hUY��'0B7�xe��ډ7N�pB#d�>Q4��e��]9���*dK �b�Kr8��2Db��W��a��,/�Ʊ�!C�U���{Ԍ��l�rH�Q5|��xB�Q��?��i`�7��O 1*�d:���eM��r���BC�<9�����.Z��/t��GַB��	J#O��m�cx	�5���`ƭ�W&$3�<�	NybM����6��O��$�|20`Є�?Q�� .���Zv�C�5���AA���?���mt��ڐlх.1��C��Q)�*�Rʧ8�sS��E�M�,�j5�O��5gV�
-6Uz�AO �8I�,�Qp�O܌!*�蕰]j^��(:�x��J��01��On�n!�Ms���OF`R��O�TR.<�BB/���+�y"�'��yoV�Y�d��V��&-J�`s'�U��0<1�鉶%F��8BK�hAX��x(�uS��Y̟(�I֟�R�ާ���������[Zwd|cԹ(���B\'ee�49��Ϳ�����D�kA��å D�Ce1�bO����u��H�˜%
�L�s�4P�hSD����S+��wq��O$D��GN?q&�D�� :q	BɻDT�	�/OޅK ���t�OO�OvX���� -���$U���t"O����Ȅp�|�i5�+t�N��t������?�'% ���@M�O��D8<�� �@�
<�`���?���?a�'�?I���?���G�:����K߉$Cf	�D1W��
�'w\u�AN�1a@���N53$�JŌ�8-Ī�Ba�M�hK���P���9b���3��G�NnX��'�<6-Ȧ9��^y��'��O:t�k��u(��m߼`�Ze
��!4��U ��2ҫ"��9�������OPtm
�Mc.O���Ū W}��'���ps-\�yB�Bg��I��%�C�'��E�r���'��I�H쐄+Fh o���r-F���P��恒P���%� ?"�`#b�"�.+�� �#X�o�f���L�?��T��	I	�a��b�:n�ڌ�GA.��O&!ж�'@��'��)�~.���C��
��d�'eʌ/��Iß��?E�d�UR�t�%��9B��!@��x�Cr����1��K�zl��eP	Z��1Ovʓ-��9V�i�"�'h�S
zF,��I?U0�agLB��;!�
���Iǟ��Ʉ�%�!H��'ڹaG� ��I�|����pmC@F� ��G*{����^��Y#f�^{�(+]o��}���^ 5G4}���|p4(�,�w�dO8Rzr�y�T@nڟ���tD]��v5��,�9l���"�r̓�?aI>Q��?�)O>Ɂq@�	QLqgl
��U�S�'��7M_ަA�ɩ�M���;$�u�V�~�@�aF�cTH���?��"A"�s�A�����Q�.b�%��H�`��fě��kq*"M����+��1Rd�]�Z�q�ꁛ@�هȓ$��@ ��G�$�:�Ӳ���R���{>d!F΅C���J�� f�X�ȓ�}�s�I�UBj�����o�Թ�ȓ��u�V�̒-�2U�s!#8$��E��l�d�DYs����*-A�Q�ȓ��31
�D����e��&$J���S�? ��:G&O�FHk(ʿI��TZ�"O��%"[�:6��6)[9��H��"Oj|���A#=Ѵ�H@'é/y�%��"O������t�`�&q��)4"OfXP��\@<$q�&��|Qh�8"O�l+�
�D�ª�  9�`w"O*�6i��&	��c�L�S�"O� 4�	�>���ؔ��=HZA7"O���Ҁ�Eガx�fE�iVD:�"O8|S�Lu��`����S�HI��"OD
 !^�W'h`q&I_�+휹#�"O��X��;_��(#����"O�U�g 8B�B�@��)bT����"Ot$��A����p�Ä�}���y!"O�GѲI�M�҉ޱ`�X��"O(z���RS�ܠ�O�=�B�u"O�L�2�(K_����-�6
��D"Oȅ�F�t�ddJ֋�LϚT9V"OR�1'T8���tm�.�>�X"O yL�5N�vMp�KVt��"O޸��d@�$!��*��u�	�w"O�DX�c��3�Pz��==�(���"Oh�zb� H���V�O,_c�5�ԏƉ��$�>iT�/r/���sӆ*R�Xf�Z)���R�Z�UiX�b%��bb���/��֝�r�L� P�bޝ�E�T�a�=�E8����)�L�����-_�&
U`"M���a�_�0��Or���&��#4|̙d D�4P֖xb�ȥ]�Pa�O�tyVD�.=�~�S'<
�O���|���
�#c�.옂BŠ|"���ҽ4-�:dǃi�T��/<OM �I׊ю��O�O��qʦ�� a2|��`�ܖu�H�d�ң��,� �OYT4�(<��6@�|x�%�4�j&�ܺl��m������(O�S$*�<AeoX�3�H���'qzD�v��3v��9�a�����8g�z睶[rF9������It �t�6�d$�S�O7�0��1qv`�s�h-p�k� �X�1�g�;z�����qPZ�O2��E�[2&���@1k@��J�\�Dx�%	3Bs|��1(�)�J�C�A�
��lKcC�9����@���Vl��'�t8���N�n}�5bՆj\�mIO>��O�E�Q�'"Hp
���\�x����'��z&��P�\q���=l��D
���O�O�U�Wl��{�h�D��%��'_���T�iChTyA�?yEp0�� ?
LT�2�V��HO�.��?r��b�;�F���îr��"��N;ĸ�@6
O@E�"e�yJ8<�e���
��hKR���'Z�U��ꏴ}��(��,��B&*��O<I` ��RxpB��7z����Ga�v8��I��=b_興F��-[B�.��n�����3mT@�A6��4��	�-]<�8�B�9$�X���I�Ԉe�7�X�'n�p+�	���'�ܩ�R�$M��4)��
�lz�����ģL����UƁ�)!�=1`�U�`hHC�Ipw�I�-H�x!�ǚ�h�sO�1\��U��p��"�ϊ�C�h�]&.({�lB�`�pH
3h�ZC�	3W�Z0[uV�m�Ĩ֩�;A0�`@��V3L�~�b��� ��)�U�C;7�Q��bǨJ'0�K$MSJ $�`�=�j׈
�0�I ]?�!���%/z=��ލ$V̵y�F�Y���<y�N�w�X��ǣ1?��Jf�L����'9498�.�'��,���f� 1@�K��sm�}`E޲-�\\��+N+��b�ݡ��"�\̹�JAk6����N�i����,��|RD�jU
�>F&��^5-��I�-J���IT~��O숑:�Z1hH>pAN��?��4�N��R�<9��>�lI`A'ՠp?�4ZB.WEF�q��ĉ������䨧��?��j��*�&y�Յ�Z�R���� m��I�� I���jy�a�']X`��'h�2MJ5�~�`�¥+H���P3�+�W L,�$�h���M��~rᚦC҄����L�(�Sh�-817*�>i�Lʓ}� ���h�H?ц��!E�
�<�萵?m�fNߟo�ވ"$D��MX��}��?]C�\� kv1S�iN�z�&��$��o���nE�#>�QϤ\λ��a�2l%�p���牙#m���	F��H�^8� �#��8r�+��9�d��&����O���G�ns�jG��bՕ�H�mE=���cN��N5~P�m�>	C�'���gFШ�~Q�e��QV��@kL7_��ayG��o�|E��a�O4�u�!D�7$���r�G�Y��)����{�	�<p�p#�*�Cި�SOP�$E�P`��8`�6���>.��O� MI���1\�d	�^�<ӗc����'zr-Fy���1��X�v�:�b�(B���D�	13K��k#��
r#=�;j����'�fމc!�սh2L���D�|-#���OZ�=E��JV�k� �Eh@ %����AK�]"�LEy"*ɴ+2 �A`P e�����I[�����
��պ����v�ޤ��#��:b0˓�Oj�J��S�&�R��ET=qV!��F&u�l;r"��3����6�G	�dіc�r(9W�+/n�r�H5^�'��Ɏgڦ��d^�A��|�2��U�>�d?6����޷is�Y�Ӯ'ZQ��լB�X8�x`pO`�
�1���M�TF{�O��q�H��� D"Ƅ�$��0+TB�9'�x�UP�HO��OȀ�cR0�,9���6jx�'�ԇ%�4��G�'�ў"}rpR?0����Ԯ_��Q��Ecc��jg�8}�Q�F��;~x��6���T��`��d�{�X���PM���e��`��&;X���@<�PxI��E)�V�J��M>l��MB���mQ\���aՈ$;������DI
��?%?�d �D����3,�	#Z~tC�5}�oH�Sƴ����S��@���'�Af��m�>����i�1� �	-�a���ԫfʂ�Q��1�؀
��:-�L�h�$=EIX���؁���y��� H&$w%�7[ۨ��m8.Y���l2�)��,Ox�*Pś�e|��g�׹�J��?9�IM�Zٞ��Q��K�U�UǚOy£���d%Jɪ=�f%������I�d̘��'�O��S�4#Q�x���Z��*,2<dH�hT�+w�[� ϛ��rZ�\�'�ΪD�qO�>���	hR�4�@HY$���K�h Hܓ X�$I0��x�V��ق�Á�o��u���_"*�� OԵ��^)(T��� �e�tP��S�9���`���_%0�B|�M�&[�P��ǀ�PV���d�1l|@I>�-��J���b�.� Tj�I��ǆT�'�U��C�'4��e���V�$���ٍvC
�$�Hڷ��[mqO�����E�>��HP(�-7���bQ��k�hU�aqO�>`A��-r@�k�K��b�Z�a��a�+-��ZA��x�I�������L��0r�	��\��'��<E9��k�'&���B�Y�a�	�'�5}��h`֣�md��8��@��u�G+z��Ӝw �a��AQ��	D��%���
6;��⟢Z'�x�j))��� x�6u�ag@�`�[h��b�������R��@%�`�K�S3$zB��?{&6�v�����%��s�S�A�S�f	9DK�����(ПGk���Ǡ.L�SDm�<`�{��1\�z����ا��O�������1�W;��3W�>1�kH�6�&b���39 aVhI_������1�/-oV\ t`�s�`�*E�	�%Q��R���R&oރR���Q#Ě�\#@4*b�%r�<�5}�ԣ<��0+"r��0�N����edItk�d��Ĺ��'*ў"}HEX2�(�MN�@H��H�H��"�
�H�PH�B��e2U���n��ɕ.!}��V�-"L@#�����e����,�Q���tn!v��0Q�$=42lkc��j���C�O�9��W/��<�bZT�����ѫ=ur<hg�j��K~���y�|PNJ�d�憝�?�s�اau`���CF��n٫��I�'��
 *Bx襣&��P�ڌ�A�'��O����b��?SD���u#u��<*-ȇͅ�q��(�5�K��@EzZw�xUX��+�y��N��[�E<[����,Ӓ�?�y�(ۂ{=���&DFm�'X�:LJ�!W�(B*���MH{��	� �1�Ƀ2B4�r0!��=�	��.�a��O\	$�̼�|:�k]0~l�m Ĝe�^�F�ص���?��Ӈ;���N�&R�\ �ӗ�A��ɏ%P4��L�yZ>|kE �A��ZMC LT �O�Os��3}7t	�#Oɥz��p�G]?~M��D�������	)
�t��ç�'zn�QK����'b�LRc��r]����Udx�#�:���'gp `Cmz�d��4Mf��t��/Н&�������c��^7~�kf(QJ������/Ma��	k-J�+��̻I��� ��",���$}D�aL�X`�L�Wm<b?YiUB[�L��Q��	ye0賤BG$"��OT�@슖TQ٧�3\r�a�c�>)��E�jQ���_�kQ�C%�&�V�'n!x�
��擂.5�PHǧ�B(У� [�nO��x&!�8#��\:o�T�I�'گ'�ҍ�4�O�x)�"]�|Q� c"���j~� V��jd�d	�<0v2��\�ڣ�O4/^��@�K�@?y��>���<i� *?HTUyr&Ц:�d`���ޟv^
��'�u���'�������
��n��P��Z�@i{�*P:C&UBԇP,�牖w,�7�I��Pe�O�]iq
˔/k����"�t�C�''��`	R���e�A��a���P�'2t��:ф2��(8�IP�[o�(`0�Ï�(O<�*ь�>� �ōw�1��'H8�˓k�R������	�e_�\��V���a���8J-�AZ��p���]�a�HH���K{}&ϝ<����r��;%@_c>~�������'�~���ɛ3y!:I"sG���$3����?
�z�1� �����V�n>����N*I~�CD,�p=�1a�'
��J!N�H=���3\�����>)����\�r�oz�� �0��1�h��Pg�g����rC�l�Z w�:O�����OHX�v�%Z���$j=�G��<u�.<�FL4�,��f��	%��3._���ъ��E��,��}�l�a�8��3�t�x��S�Z�$�h!���*��h�d��*)��I�!1O4	������:�/]��� �ШW�G>����T �Ɔ��5zx�C�!Z`�ӥC�/�����7r����IǒH�~�ś.3+�eZ�2' ��V�8�N�4V2��?��ƟHlbY	�P) $�Հ1�D�q�!�Dބ[[|4"��	�C���r�$G���L���Wr��A:p�8��?�p�,W�Z�ψqz���f�L�v{t1�e�}��d�}�~��K.��!��]�\����C�#�\�x�'Y�r�JA�'����	 XY��Ō!��Ȱ�����������'�9�L��eIU- �� #[�B�����uX�əuI�\���_n`�[�͈�ā�ō�+EAB�'���'l(J�f@� \3�*�=/�DX���C�3-����jZ�e�l)D}B�ڵw�䌨 /48�P�-�t�\Ex����DӢ�'H��k�dSJ���Q&E 
�X�p发V�6T�`�X{��u�D� b���*�w��)W)�0,�C�J�G@�p�����'}(�BF�{e�y���E.@0���
�]ɓ�D�!1��B�MW��Ä<��'j�� �A�W�,�� D�k��&�=�
4{��4��ɒ�O��I��� y���eT<h���cP!��/�x�i�N�8B�Fā�F�B��րW�fl�㟒�.%�cGH$4�P,S��
Xj�ᖗ>Y��T���"�%߅D��	���j��%�6#a�6,�X8"o��`��\[&�D���0|
����`}0��\g^%ca�P� `*H���'a�ɉ��O�^$ae�@��r�K�i�����W'�!I娃�!��������7/�F�bu@a
P�`��L㟠�'(��/��*��6B�
Š�<14�Q`��5A��֔�
�3�ؓvy��I3t[lL�'E�|:R��!_Ş��� �QNh'N�^�2(!�]�+0�'�LH� Q�1�s@�w+���'���m�<D�=I��:80ec�'2�Ix��fŶ���OV�*I2��'[�Ĺ�j�vtL�b�_�md0�`�'p��&�>�$M��Eþ_�H��'��xp�(��}�J�ʴΕ2]
�[�'jͫ0���c��k�ȉNT��	�'�*`��Y�O'�!IW�V�B����'�D"�"P(M���Ɩ'd����'��d���üx�{E���H~^�{�'D�RS<DҞ�W6�L �'~�x�G�U(&p���|$x
�'��M���H�U���Ѥe���8!�	�'/x���`�<a���N˔�@	�'o��Xw�ٴ2h���cn���h�'����Fa�2&��zծ�+�'ܲ`���m�&Y���D�v��t�
�'Ռ�w(ݷ+\M�` R
l|z}A
�'`�Kf��c+��@��ٽW�r���'��T@�@2Y溉X'�Z Y�89�'��yjeM>D �	���9XQ���'���ťQ$UF�1V%E�����'$} ��C r�I�#�v">��"�H����;5�[>���ȓ�L��a��O�}�&g��pw���ȓg�(��6���"���#JB5�ȓ�J=I��+\���	�KY>H�ȓ(ft�i^�?�� �$�,=�`�ȓwfvA9���3��|���VKX(��%m�E��&�]�bi����z��8��mF �I�͟9������%
Ʌȓm��1 [4}l���16.�\�ȓ���Y�B.���q֭�+,.����y�(ֵ&� ��C�ys�E��a���pV���yڣ�+�,�ȓ_�0l���Q�Ei<�)G���)ÒЇ�Yʢ��@(5��3GC<���ȓU֎��]t��������S�? (ͣF��<���8d�K�|��0��"O���%E����ܖj�Lr�"Ot]���3Ulҭ��BV4dI�"O�a)��5S���P��
�q��"O`�Kd���gmn(s2X9���ɗ"O���w�A%c����$T���8E"O�����.�y�#�>0���*�"O��[�.-������@�Xt��"O�Y��;y�!H`��,�0"O�pk��߉t�Qh b��	^q9U"O�i����@�"��P�Q��"O$�z%펞Z��x��\W10�C"O��0�O�>뼵�''@%Ӥ"O�Q����!	��P��Wb��A"O)�	;lX0}j�D/��=B!�J1d<�	z�Θ5?�YS�%Q�!�dńxg�1� �8Z7��R.µK3!��Z�wqрDZ9[%-�� W'!�$ũ	���K�nG�."��bR�2!�F�7`����W6r�8��ހ$!�J�P���uTz�0��	,ZT!��_r����B1<�Z��R#N�N�!�W<��b��߃-��D� `��z�!�$T�f����غa���R4o�T�!�$\	'?�[��)Ӑ�#FC�h3!�E4^� �	�Q.i�p�sFdJ+!�Q�,?�h'ˑ�	6hQP�&M'!�$!bF�� ��(y<Շ�{�!��
�$�l��G�P 6\r���\�!���+$�XZPo�JCj�С!S��!��τ'1����	S:H �mA��!���^��q��ǳ4v��ՎТL�!���*J��]`v�/h�H�kd��O�!��@ ��B#
-��Q!��ֶ�!�dǘ.YLș%iG�,�t<��� �!�d��\b���5�H��� �!�~�P���↱
�(��"e̓ RC�	��l��X�Q3�s`eK�u�*C�I��
UG�8ׂ�b����48C�'9�p�!A
Iv�wI�?��C�	�G��qk��u���׮�WZ�C��fb��W ��k�b(�
D�8L�C䉇s��1�v�E8<�,(�R*5��C��&<�"����?sh�M�.�FC䉰Ę�5� -QN�u"�/\�5��C�I�Vbm�e/G�c�ȅ�5/Y�Y���D,�8���Qp,Tl�Xl����C���ȓ/a�YA$�?6L ٣�̎	lx���>��k&�	%G8�lK��ɻ$��`�ȓB��u	�C��YI^����PA���`bB;Q����ǓK�ҁ��yP��j�L�.Zi�ݻ�N�7w*1��k��<Qr��d�:��4e�.���\�:͉Ŀ+��Ё�G�J�:���C�p��F�:k��ե��kO����|@���NP�w;t��!�$=��	_}�Gͻ0}Rx�!�.pQ���Q	�y�L�(�V�9�j�+l,0��
_��y��n1�:�`�;4�
��℘��ybAա1�>���&4b��$ ���y��ȡ6����G���S)Cq@���yR��	T}T-Q�З}�=���L���$&�S�Oߦ��b�$,�y���#rInU
�'��������f���$[#ԾA��� r	�t��B�ȄB � H^qA�"O��� ͨqX�Ջ�Ȕ�?��Y��"O���������$Ȟ�&���:"O� T�)0ȕ��a�<=-d�a�"O|�Rb(�;�����F�6`�u F"O�̐�J��H�@u0#[�
U6�K�O���fbL�ZY(���5P�L	H#�/���y"�5D҄�ac̴z��mQ���!�^� �𑡇�Y�*X��Z�h�^�!��R�v�����I�\qzU*#�
��!�[+!�@�s L&Y_ �¢��[��O���䚯D��HS�K�7�ȼږ&p}T�ȓ2G�-j��xR��ke�!|��u��':8�����n�4��W��G�����'���Z�"�,�nx����>�%K�'R-�X�=Ȕ�!kX�6!��I�'y(@�f��?��]pk�(��1:�'�r�`� q�P��^�.���'������̄mO�)2��J�'�)��'K`=k3�#;� ����U�^��
�'����ta��$�Р�!'ھ=sҬ"���'�,����|+�T�_�!��'Tֽ�D�� 2bGIrd�	�'%rM��ܲ���r���=���*	�'8x����20����̭=����'��4�Ľ �P�����1�Z��'q����'C�~�����&1z���'�X���o��4M��h��0H*-K�'VlYb -4C<ţ�-[m;�'h���AY*i7譓��$<(��'N������zk�yJ���2�xXj
�'M�dK�j�8�@��ӑ/:��K�'���Q��҄h�|����.^�ܲ�'r�%*�D˱+M���§A�8B���'U&i����#T{������jN�u�
�' ���E��D$�dz�F_
��'(,]`lG_���FN$]�&E�'�0�+Eo�7� %9N������y��^7�D����2߶= pb���y�G�r� �q�� �7��8C�'�(O��򤜣j�J�Y0lؕ?�H��fB� C!��B��I'J��nҰ0���%�!�D�ES�y����c��a��)V�!�_����C��/�^�ࠌ��t!�$�*i{�9�����궨�$�!��X��; ���� ��i�^�k�"O0���ՂG�(�Qʃ�*��R"O��8��ڛ0���K43v�*�"O:#%eK[*fQC��Ǆf�$I7�x��'՜���ם)��+ BK<���'�ҫ��U}|����c}�0Q��M��y�C�7)�h���
X�h��rH�y�
0�p��� ��Q@6�k����yR���p3T�[�C�X\��K �y��Q�eUܢT-�=���5E� �~2�'��]���3wqT}�ɼUv�B	�'�L�%!�	 ��ɠ'IIje����2BÆhI��2�	�"�i�1�?D����\�?Ɓ�Ȟ34I�e#��!��hO� ��D�TKҤz����vCZ�1B䉌L�pꗬ�� ����W��65��C�IM��TcX4X�M�&"V��C�I�p�$P@%QDu�����F�K�|C�I�kT�]��A.|BV��C��	(B�)� 
p+�K�u�� ��mV9�"O��)өX	�)�-Z�#��4��"O �)ӘZ�>yC������P"O� :�GN�l�KE%5u���
M��~��)�'�6���L��Zƀ��èz�d�ȓi(و���p� �Æ�A�"v���ȓP~����7�PE#��I�<���A�� B�*�2h�N��0��Ah���^A��W�܇	�d\KP
s�@Q��l�L�qE�&^��0�Ӿz^����[��1!��4'��Jd��0�Fa�ȓ$1`H�T�!3�(	�V�O�b^�ȓa�t�%+Ӟ�^�R�H��4�ȓ� ��TI^�_�)ꤋ�U8 %��!�\���ތab@ۏK5\�ȓCO���UbY�n~UI�ױ��$��G{���l��o�64h ���d*���yRE��4�}�E�H,� 7aԎ�yV�3J��`
�	lI3ƆX7�yRCYL{~%���*l��Rj	��y��#,OX��Q"Х,���A���y�ޝGF��1g|�R�l�0��m��u���b���`V �Aա;�D�ȓ�Z��P��0x���V'�؇�xQ��x4��Z�`��b�ΖA)欇�3� D���_�Q��y��芪 J͆ȓ!@ځ���R	M'T�6�@�+!\O�b�@�Q�]c���%gL hLy9��=D��۴
W i*Y!e�ߔv(#	;D�p;��DX��b�f܋{.u2#�<D�����
*4B֨W�}��)E�9D�8���N�dH�%h�0����$8D�� �ڊ	��Qa�/�&ٛ��#D��C�mU8_���8!P1d�s�'D��C��:/��B��P�<�;cF&D��@�����V\�;� s�g"D�$+�o�5in���Ԭkr�81��#D��Q,�/�
���'��I&򙱄"D�ܢ�H�5Dq��:]��EKUi D����?�����~��!B�F D�\qf�Z'TtDaZ�˔���1)r�?D�d�(��1Ŏ���bR1A�!�o?D���v  1r�����D��K�?D���wa���(أF�+3��N0D��ئ���V�BW	��E^�Ԋ�,D�$¢ըg��bQ̝W�$ZSH)D�4CPJ�[ ��b�W$�>��E�!D��B��ؾ�T9@�a��~ba�7?D��!�OD���X�O��T�!a<D�H��C��j�v���(?s��@� <D���%T���e��v�����n&D�Iq�ڹ%���B�a)��[UO%D�����9%�Pi��T�=˨3�%"D�T@pökA���KQ��d<D�P �O0f��|+C���WH:D��ʥ'�?���0�zO���+=D���I-x�JE*0
��q�S(9D�С`g�)�����х<E~!3��"D��@�AQ9�����`�w�,�3q�"D�(�D�09�� go��t
��:B�&�f�'�ҡ%R��R�R�|?.B�(>ҕ��S:RnaHC��,B�ɚz�jX�倕7s����.��4.B䉉Y������G	lC��B�"]�"B�)� �i��l���U�3�3"�ViH�"O%�&$�"?�&��㉟�d�`�z�"O�!�i2=1YZ�Oup����"O*M��c��&b�ã�-=\�!zD"O��Ɵ�)�2�s�͏6h��y�"O�<&�4},R�C��ZLY��r"O��P�@%X����U�X#Z7�t#"O<���ˑ�S��*bߴ^.B]�r"O�ɳ�J(}��g�^�t�b�d"OR0���Tw�,�C�	.Պ��"O9���WY$���9)�"���"O�\K�I������MVz����"O��@�66+:,2���� ց�"O�]+W��#C�ԫ�=d�� v"O(AY�
�j\P��
X�p;�!a"O$�q��OH�i���4���""O4��2�ڔ~��+Јߓ� -g"O���×)%J@�F�p��"O��1�"D[|����Ȫ�J}��"Oڔ�Y*)?���ƜtsrQ9&"O�@��o��bn��qe[A���j6"O*@�4N֒�,����hHrp��"Of���c�:b�>��ݫ,$���"O�d9�/ ~�P���B�$��x�"Oژ9�h��(:������4.���"O�	�㮌,f�+C���h�c"O&���F�e�Ĭ��j[�}��K�"O��j��@���b�gL�[fQ�D"O�=�lǓ	'��y���BD�}��"O8�;���\�M�=*<P`�"O�!ǎ�XL:�h��ßƠ`e"O��� �(1�,|���/�	r"O����\�dXՊ�-=����ȓ�V�i�
4C�+�-�%򐙅�z���ǂ�.�P݂�dƢftq���Dc��4Mv!�,�83�4���jU䌝>�	�Q��Kߠ`0�"OT�E�-D 	2lV��p,(c"O�1р@&��2��9¦� #"O��������i i�
u���'"O`���@�9���ݢB�tX�"O�	,]�&A����dZ�#�-W��yBK�96����b�t��t�Ȃ�y��:'DkBǒ�a���$f��y��R�	V�3���*G`@�c��ybd 97*D�JUb�""���f@���y��R)J/��3F/�#f-�e&ä�y�\9h�2��f.�? ��0BU��*�yr�:;��E0�Q�y�\�c	�*�yb��m>n��cޮ��b�ͫ�y�j�7��kgeX��ə��1�yr�PM�u��N�Ǡik��*�yF�pD�����}�X`��ۖ�yB�Ҙ�bL����|M��e+H��yr��"���c�s���%$[��y�'K�S�,���9o����Ɯ�y��a���Pi��d�j��®Q �yR�5N��G��Ҽ	ӌ��y�C<b�l�r�,���IWL�C��B�I+lq�W�E
 U��+�
�LB�ɪ~���ðh�S�Xa�a�0B�I;4��'W3ڈ��R؄{tB�	-j	"0CƎ�8� ���D��C�I;"x"���.z��Xp�o�/m��C�)� �ucg��4sذ����}Zv���"O�<sp�A�E�q`�.^�O.G"O�I�w�+P4=�nA6@M��"O8Q4*�/
d�{6o� �h{p"O�p�rg�) Y�H+Uc���"Oa� �J"Z�5�m���s�"O��
�m��,�Q�/\O���Y""Op���6It���q"�,g"OΌ)F	O����1L]�M��y�E"O��s��1\� z�떡(T� "O� �@ϵ8Fl��@ZMx0ES5"O
07��??��� i?`[�D�"ObX��P��l��d⍉Z� ��"O�8!gj(zG�e��ɤ1���j0"O�]�G]N���{�*T�VVe �"O�UH�'/b�&�Z�<o0K�"O�dk^r�@p�aA.\X��y�
Ѭ�yB�ǿ
���H�U��Y%�3�yB�[�[/d9��	�P�<9aT��y��(U��9qn �Wt����%�y�"�V4�]�vaC9損"-ʟ�y�'G6F����N& f�R�yB++wF���gG�@�p%��C��y2EՊ:Sґ@�=7豲��'�y�aC�|��
e��	F��q����y����e� ��b��8m��PN�y�H
#��W$�85r�dB� �yR�نh���uBU�-�����?�y��['��
�I��p�1�
��y��&D6� �б�p)�����y§Q
!R�`��Ǖ6h{p���y���P�(m`�ǔ=h�ؐ�\��y�
�>-̎����-P��)�	2�y�Z�$	��G�#��Z��4�y2Ó<�|]1tMh(��$ր�y�K=g}�D�w��"mX���.�y��
�C
�Af�;]�`r�h�6�y"���= .,��
"2�&��F��y��ؐMy��@7`�;w��2/W�y�i ��q'NL&�r�i�`�1�y�N��"�S	:
t0'�?�y���eU"d��	*�Z�'��$�y�_D�Pd��l9U��Th提��y2��q��)�� PP/J,y��ؙ�yBi�qj�혦3���%�<��d�ѡ,���i[0"帐�ȓz�@uH%I��� ��fV{�ʈ�ȓ?d�*�i��]| ����u[���ȓ:�NɁ� ��8{'�������=�"ܺ��Z��<#q
�&F��ņ�pG$A �M��LbN�j�h"�D���}�����B׹(Kp�@��E�X4���Jp2sM�8�1Hw�ǜ��Q�ȓ4��ɚ�l���ct��i�nE���p��G�3G%%��˪#p��ȓ�|īT��g��mh��0@f̆ȓ#����F;LD�Bo�(%�*؆�P\@�U�Cg��x�J� ډ��\�,�)��H�QXP�3����$����  �p� �QV�ȓ^�ex���2ZGx���Y�2��]�ȓg�65
̖�a��ZE�âv���-%)Yuj�ha�9���	0�R��ȓˆ�3i`�1E���Ї�S�? �p�/��EZ<I8&Y�t-�Ęd"O�-���6}J��V�D��R"ON���E	�܅���L�R<��"O@Z`I�u�N�S  μ7X��"O��i��9Worx�&.?�narw"O�<�'
/V���-��3�IQ%"O�y�ܼZN,��lJVa� �"O(L	4eM�EI�a�ҋ�>2��""O��r2/�."h��l�Z2X��"O��12Ę�F�\�Ӥ�;*JUJ�"O�E���؋@~*t1�,�R��&"Ot9�&��g		��듿s�� �"O8�Ŏ@����`�������"O.R1Ny��@(�HH&,:h�"OJ�����A��غG"�u�G"O�{�E�Y�$=9�i� �F ��"O��tcN'\�}X���4Kz8�"O�T�sF7e�$tx�C�O/2W�y"K�3o���&"ӅW��9��ǈ��y�ЄV�1����H�v�p ��y"� 	$(���#P���j`!�,�y��B�p�6��o�v+��1�����y�ꌂmd�)H�h�	�ŧ��y�	Xj����q�O�d����@Qx!�dZ:`�(H�,��	v�Jd�0%�!򄘲w8:lr�	>)�yٽe(!�6Y��b��{r��
o!�Đ�K_RA���S\�� �*�P!��%1���G�ƈL�DE3ժ���!�D�U�=��\�=at੃I��d�!�i1Z�sU�3ALƽy��-4�!�$̴%�ȐQ����"g�U�$і�!�����EC�T�|����Ӽy�!�D��@y����@�tcP�!�׏Z`�� c�!V�ȱ�!�_9�!���1��!�
�x�<�4ߒO !�×;�XP�F(�x���{GD�o!�D�'R:��P�����ĉ���%!�Y��@i(��r{����/�?^�!�Dһsuy���G$hl�)�Wo���!�A�1�V�ae��(uZ��(�Yw�!��W�Ri�0��4Ii�d��F h�!�ՆO��亱#�=NB��3�KS=�!�$܌.�Ԩy���:���Dm	$�!���O�V��E"�)
�|�c�L��?�!�D�:�p�ʡPy6]aWM �!���h�����ˏ�$I#b���!�$�]���B��-}�b��yw!�DʭG��$���</c��P4j!���L��(W

5��-�@��.g[!�D]�0��.%;X&�����>!�	B���I 7)��7`҉(\!���;K��@����!@��w�W�1�!�دQI��C��F�plˑ�ؙK�!�d 	�h)a��X,3�4x�b��3_�!��A�1��A��,�y����(y�!�ėo��A��!X���� ��p�!�D�>�p]�Sl	#0p��C'��X�!�9�t��U$F>A��,ɐ[�@G!�ą�7�X��p�Lks�,JN7A!�$�Pi�to�un
YW�Z&x�!�䖌"{�!k�M� MY81��̯o�!򤜜ֲy� ��/�H����x�!�$ݠn�8���X�^=K�j/3�!�� �E�ʖ��9R���d/���"O^�@n�
.<d��s�(F�)B"O���� �)lzػ���M荳�"O�D���G�(j��+���3"OP�g��L��	��`*B�R"O�E��Gn+@
~ڲ��7�;�y2��*IsjD�g���%[�k�zC�ɽIˊTx��Ϭv)H���"�?RC�	4U��H"�'�J�j�b�;HC�	gwd{C;��p3�"�qC�	�d�'�A>l��ʁ�.��B�ɺNX
�QO�O�X(��P��B�I�4ʰ���LX^� ��!{�B�	�TH�2�Ո;�T�HG�
:C䉻P����W�O����J�)K(C�Ɍ8jq��%M�����A	>T�B�ɱ	c<,�7�U�WAV!����}*B��?:q`�C�A< Hm���Mm�C�I3jY�ɡ�I[u
MYg�]B;ZB�I������4������+K�PB�	��T� ã�Qz�UA�lX�h
.B��!ZF4�����-(AB�Z�"B�	�!y,q�/�
������6F��C��,7!8����E��O��jC�	)Nx+���gBT��Pi[)
C�	�	�>(�G-U�tX��|��B�ɛ"��$"�(�����U��k�'X����L�i�bCPKE.a"�٢
�'j�;��
\�3�G�vX-��'j��q�@E@Z�E���	#��q�'�1p��(E�<P
c�v����'�(:rf�A�P�Q'Σh���'0��RoW1� ��f�G-b�!	�'�Ri(g��&5��*�Yt�	�'���*����/	�H�����'�vYj��C�!���+�X����
�'V�� �!ڍs�4�L��S�-�'@t%:�R�D,��EFԺy��y
�'~*�9�C� �rm*&��'�����'7l�����%D*�	#��N�b��'�bDٰ��4fD����|�2�R�'J���$30�p�$�IqԄ��'�
d�f�D�(~�T�s!�	i��@��'���� �/��p�c�"hNP��'��œ��R/֌ٸ�`�sm� ��']����W<:ŎM1eAi����	�'t�X�L ��cH�]S QY	�'��C�n[�J�9"����*
�'אl����}Bd�!��'2,�A�'h�r�ʧV��Ҧ��l��Z�'�҅�5��&!+X�6ƾ">��
�'�f���B�J5��s�	����@N�<�`K�6^.&\��ޮ-��B-TA�<��ʀ2)�Bq@'J��?�|p��}�<QX8mJUOнQ�6qJc��=Bч�-��L�B����5 (��d��B�I��&�FR���� k�����谢p��	zv��6�<J 0�ȓ�
E"%l�� ���5J|L����\�DR�+q���ʒ%v��ȓ$�|�t+@tԄ�c�[$w֐���5.�	r�؄TIhMZ�ˋ"o� �z�7��>4���N̤e��ȓsT����KKIBl�r!�.�0��S�? �sA1h�l͛�ϐ�sy�Txv"O.h����>�JMp��
�-x^��"O��CG.�8N7~4� Ōl���u"OZ QHݖj�]RV&P�R�PT"O|Mr��'<�P�A�3X>EIv"O�8"c�ߍ6J&m���_&*�)�P"ORŻ�&�6d:E��M6}4a�d"O�Pb�îzĊ,�֮"VD�`R"O��0ҎЂ[b&<����;=Ѵ��P"O.�q7`�S�J8(ፐT�*`��"OL5�π�`�m��	�;����A"O\�q�ؼ/6^m�	��!���S"O�1���T-ko�� çK_+:�w"O cώ".� m��9�!�"O���rm�e���0�W�k�2���"O���'�N�ATy���<q�4Q`t"O�1¢�6�7�Ϯg��q3�:D��� �4/���C�ϋQ���,D�0�t.	%o�1	�W�f	p"G&D�L��MR�6�mS��8)�I>D���W([oI��ʤA=+�x�C!D�L
��U6/,�4C�뛍`ܴÔ/-D��QDk[�;w�|����z���AK)D��s� _�f$���@��Rhu�#D�8"B������I �^�衮"D�����hT�e��	/�@���!D��jǁ��MȒ��f���X)�ͫ& 3D�T8
��T@��H&ۀ��(>D��ړ,�S�XQ�+�T�V�H� 7D����$^�|��$e�j�BТF*D�p9��<��]
�a�d� <�Fg:D�R�B�3��1�N�"�HA�@9D�Ă�l�8b��m�t�O��ph#3�)D���F�
�ϴ�H3%L�D�N,��A'D���m�7ɾ9Q��/���R @*D�H
��S�,��p3���R��Y�(D�L)LѦs�*P�tC�U���&D�(k��Q�z�#V;7�]�7!D����A�K��=2�]3tqxѨ�#D�,`G`W�m��������Viq4J"D�t2�cߵR�V9C���~|��1L$D�ԉg\�M���C'�B�v�q�).D��w������+v�:-9�(D�,
�烤&���5B��\�N-h7�&D��´hDS�`��`��F�&�@,%D���A�X9�,5RV(^�e^m���5D��;H�3~��
� �j���7`0D��A��S� 갍��蝖;��u�)D� B�MS0X����YaB��J'D� ��-�=);(h4�iԶh�d!D��J!!U;���A��"U�؉D%D���R+V�<$��c��gX�1-#D���$HD�y��])�'�$Z�v�	��#D���S�
	�r�`�� �����#D�xQ�fa@�`Td��@�h��B�	�B��a��"�`]L�yе.��B�I]0c��/�)Z��I�?"�B�	pTj���8&8�Cf!��&`BB��%?� M�����𠹣��B�	/�'�s`А�S�љsɢC�� u�Jੀ�1-��T@��?Z��C��<B_�U��k�>#���u/�tALC�I�mC�@��"V뮈�V���t�"C�	�wh{ѠD8(��8%d� �C�)� B���h��!2DE�`>\��"O`�D,Z�P�F}�&�
�H9F<i5"O@�����:��\+�	Z�A(�b"O�7��5<��+�Ȋ�U�\�S"O��;�J��j��Ģ҅��,^��Q"OR\��A�+�h�4�Q��,��%"O��	�JS�F$*�r$@�O��I"O�$�R��=��(�a�6.��Q"O"u���Q�N��Iȴ���.�Z�b�"O8�ː�W";�j=�G��^��2�"O*�r�	�=j�� �2}�i�4"O�H�D/�d�HO��w�c�"O��qG��6ҀY��� |%g"OP���M�w~D�M�3�d��"O���D׳?��"�këA�&�s�"O �� ��Tv�i�vJ��5�j�[�"O�䙒$Y?k�d#�� (�����"ODmБ� �'�z�a�Dߝp¦���"O�p��I�L�qQ��!�X�I�"O��yS#٬�0$���0 ��"Od՛'-��ځ�F+���h���"O�P
$��"[-z�{#+Q�a�${�"OP$���Ȗ~&�J�i��y�ZL��"ONX�_wq�I"T)�;1�8��"O��1�� �z��h�.,�B���'�h�" �'��0�$ȏK�"���'�9���!C�|]�"�\�X0R�@�'��R�&�ô|9BR#�z̠�'}�h���X�cq�=Ca%�&m�
�'�)#��I�:��3�Ekq�t�	�'*(YW��^�ZhJ��]>f���Q�'j���Cl�(}�h��p���B�'Fjt)W�ɜ�욂c��cF<��'�ҹBR�����R(O�E�,�@�'|Y�T��	Vt�-D s�:%��'���8f�>Y�l<�����:����'sTqcn�%HN[��N�>njQ�	�'���J�!
?͞�U,ҧ1��k	�'Ĥ�A���8�ni1$�9��	�'H䄊� �z��S�/-���'�nxn0Y���KC�sw�u�'T���DF^��c&���q}L�
�'�����CD<pnXkEG6l�@�r�'B�t�Ӫk�����5�)�'QMiC�C�#���Nd��Ub�'�.<xv�B4B�����U�`8 �;�'��`�
]
`�ƫ� V�Z ��'��ٱ�̊�Hi��CC�Q��y��'2�����*7�M`�.P'Ķ��ʓh>�A�'������\���D�ȓ(y~!9aO�#"=*q@!����g�J��q�S�Prs�k�L\��W:�m�K@7F/�ţ��Y�+�هȓ@ �i�H��9)`$�U���P��h�ȓ\�0�Ah��!4H]����ȓqNh3")�3ry,���T;(���U�1��]"ȉ�Sn�&F�L��]#D���E��=Xz�.ɹN�$��/wJ��S
F�&P��We�9_w�Շ�>�BXI5���Y��	�!N�4]�ćȓy�X�"d䟑2�0)4L����"O2HP�D��]���CHR.Q�2��"O�}�&��,�-I@��rQ�"O,e�&�ƾ���ӡ\A��3�"O� �IAO�]�a�f�D'3I*�"OFqcp$L"L	���ډ^1�8��"O��:4�H�5izux�d��O�A��"OPX��e�ah)�6"$QH�U�v"O���0%�W��`��#�<=�p�"O�X�"B��pt�H> <�z�"O���f��L���Q��0�"OBq�p+������1�J���"O��8�
�.(��d�T+F2�h�Jb"O�\��`�0��*�_��Z(��"O��Zm��+i&,{娀�(��<�"O )s��5y�@|��h;f@��r"Oz�9Di	<���p!iR�V�" �"O�K�A��-@���c����"O�I�C睛Hm�U�JNj�J��"OlD��ED�,N�	 
Ԓy~��""O��K��T	ؕ���_-uv�y#"Ol,
�AP�V�iID,�(y04"O�i�vg����B3��u#J���"O8�2D��F��)�W�o�����"O2[�P�d�s+�.N��A+B"O�ɨ`AZM��c�i@ r���"O9sQ�< ��dI�	�7�l��3"OJdad#�o{\h�I��ve`�"O��[W��V�,2�	Ÿ`φ5��"O��'P�^��P�苓Vͪ$"r"O4sp��� ��5aHʧC�~|s"O&����v]0-�%'�)6*��%"O�Ј��t�4a��=�R�3"O&�����+��x `���š�"O옻�O#Cwt��tIH�H�
l��"O���U�w�X�W��d���xf"OLx ��:J��0֠���Đ�"O������/: ��eBT�9�p!V"O��C�jN��t�����;�*���"O���#ȃ�a
j�xN�=iފ�"u"O��uΈ�rJ�@���mh*���"O�@˓È�M��$!F�ߚCW�|�"O�X���Z��Pl�`��	Vf���"OHmx�m-:�&� E'
S���e"OH�AG�LY%"W��E�9�3"O^]{�J�+M�X�ϛ AF� IB"Ol�%d�78�E;�HxC`�a�"OB���ı�pk�-O1:|�Z3"O"x�!l��/��Mj��T�#B"O(��W�ľy%�5��&W��
x:"O@I8��$z1��@�rB(�y�"O40:#�[�+�2�- �f�+"OT�p���D��(A݆$
�͡$"O(�Sk��g�.[�kT[�D�z!"Oĉ ��Y i�1D����"O��,ZPv��%N� ��"O��s���	��ǘr����"O��Z�$�F�Ω)V��U��P�"O:d�ebU�1[��߯svF<)P"O�0ا�A�?���x4��wrJ�)f"OF�c��K&}�4��̅�,b��"O�җ!�$)��IA�k�a�p
�"O�PŅoc�#
�X4Ԣ�"OT}�� O��hi�*�?M=T�ɦ"O�Hi�I�"�,����/V�z2"Of��C$$EL��  �a�H,��"O��1C
K���󉊃Z�,4k�"Of8��#�{^�4��;��H"O� �2�BՎ (�ؕ���n \pqU"O
� �,Q.|`р`["\p�"O^|�DݢT���.G(Y8\`"O&(j��ZF09�M֮V*�ty"O��*5
�16�(�WlL<��EZf"ON`� !B�,�fƚ5���Iw"O�"(�#=�:������wTL5�!"O0�@b�<�ؐ��H<oNv�"O�Q �o�k��M���FԘiC�"O���æ�98�^)��oD)�>5I "O�5���<g'peH1`ω]���!"O^]h7犼	D�9@.�va��jg"O�����-%� �R�BU6���"O�P"�K*U���җ�ߍk/AȆ"O��!�jD�s�h��, ?;2N�!!"Obh+4!�z�Tl����3��C "O�t١�Ccv��F�_F�2"O@��p#���$���'F�E	�"O��q�K��*�숣WgR�Viĭ��"O���aaQ�p�0,��P/`�\c�"O��B2:h��N4C��3"O�ِv 
k�h�
Q!����S"O�����t���2���3��I�"O�!���*~s�����2~Ƶ��"O��!�92Y�ț�m\1�P%��"O�M@�`��BBex�l�Zb,��3"O����V����3�\�r2
	��"O�*6��.Sz��W�U�A�"O~`��O�H�d=s�JI�4��"O��P� :9qL
BɁ�V�|�"O*S��$*I������>A��"OnH��FD�?4�ȧ �.,����a"Oܽ�dҥ'6���v�B�x�r���"O�`��.X�/TJlX�nD�]s``�"OPPJ��A�kg28�$�t�S�"Ozie
�%jb��1��mkh%H"O(���׃;��;�k]&Ne�}bE"O�+�J"0J�\ri̳.Zv��"O�M�P��88��"r���ñ"OV�y���gN�\X� K�o�,��"O�up�G�P/6�;��QO��b "O�\@���+Y;:�24�_ d��q�R"O�@���)ߚ��t�@L�JQIc"O���m���� (4$K��2�"O
EuN	�;�ޔ�㕧k��:�"O�P�f ��ږ6D�7W�A�&D����nW-J��㲤ܩG^:лƫ D��:A٫N��[�F�f t%82+=D�<�am*�ʅ����2F�%��=D��q�*�{�	VȂ�$u��'�0D���!n]�\;��"䇁�7��|��B0D�i���)�`�m�.&舒s�0D�<ӄ)�W��lh@!	9X��)�+D�x���N�`� ��B�R��Ҵ/D�`r�
��T|�,{G(�l�Ȩ㇬+D�4��H�,��m��2�8���>D��Z��@��XSꘪh3, �=D�|#� �{����V�8�"��Q�:D��3�e�*�*�C���e|�0�$D����)U/�~c�5CN�z6	!D��v��-��(�iI�y�X�s#)D�d�l��B�4�G�G�`�9��&D����Ӿw4��:m�!���Q�	 D���,���J�'���|@0m?D�� �,���n�4��5����,��"O"ip� 	;ˆ @���}�R�S"O����D9���� Ȉ4"���"O�Ԓ�GL&r��f�Y�)�P���"O �(�DP8X^����Ԋc�.0�"O0�	��VL��-�6�˝/k�x��"O�D���$ic��"tm]�-�*��"O*�AAKʝ��-L�v����3"O�I�⢟"s�ڙPuؐlI
�"O$L�Bo�.^Xأ�K�3Cm���"ODL2@�>��	����d���U"O �A�K��uU���'L�$oOp�j�"OX��ƅ);��!��u�L�1p"O����94�aY k��xs0-�"OR��WḺTY��!I�Or�r�"O��T˚7u�(qjDF�	wT�ȑ�"O֜1�D\����@営VB&D�R"Oi��_x�����X6/>.="O$��cK�`�6e2���I�X��"O���ׯS�w�����y��	�"OZd��!�6�=��+�1�~�5"O+�?�r}�񊁷�$d��"O���f嘆�th����E��Dag"O0L{&^�X;�H�Ed��C�e��"Ol����=�x1�5H� \Y"OZH�K_�{rP��c�0m����%"O�-۱!�0���0�L�6�Dy�"O� 1�fӳ@�`d2�I�)$s�%X�"OZ��.g�pyY@�!xp� ��"O�� iH�
���n"pg&]��"O��ʀZ��p��P���3�"O:Ƞ'`�rMZ��H�V��y�"O�Q�&�ʬ>�Je� NK~~����"OZ�����1B%�q�2j�"Pv4}�t"ON񨦄��V�>���k�Tx�aY�"O�=v���#��A0l�A�"O������[�&����?�@
"OX��I�G��q�2�&c5"O��(Q�E�UҨ�&�C/����"Op�l鍗 T!����vZ| 9�"O0l��ł�{ڌH4��e4��K�"O�j% �3sK����Ӻu$l�à"O��R��Y�s`$���3!��0�"O�Q0���%�0�kT�Իu�'"OP8��-�Q(��K�_�r�"O��I"Hs7���"�׸q��Y�"O��XU�h�x w�ltR�"O��ðɔ#P��%�k��h� "O� 0��̗{V��k�,���0��"O�M�TF̬ҊS��8�̡"O�#V7ܪ|��)��m�����"O4�hfOĐ))��p�� ]0�9�"O�K��<\5�UC�Mq�D{�"O��Ue^@�9��*X:L�^�#�"O ��"���k�z0�G"O�)aC ���k��
HX�"O\pѡ	�h�\-����2G�� A�"O�In҉vS��8�ʲ3�����"O�W���e6n�{#dBx��Z4"OPsAL�(t����]ɜ��G"O��`I���܁��NE�4|�"O$A��(�TX���uM�%{�'"O�0��ą>*+�XJ����f��"O:x���/l�p0NH;0�����"O� \�k3�wr$Xْ�*p+�D"O�m{��L,oz�m���"G`"O����֕F�2��C�^�( ��ɓ"O���׌E�A<���b�ް
����G"O@\�e�Agr�1�$	����c"O�(�� ]�X&t�d�*�,l1t"O�%#F�0�J�i�ME/��:5"O�����-����F�O.dM�T"O�У�oI+}$$���FX'L�z4"O��P1��j9�gŞ�:��"O�u24�V�)���̟i꘍��"O�����ަa��P3�ԡ�����"O�q�r�,}���Y���?9���� "Ot��ӢU6�}@�Hwڲ��"O�m�ׯN�Dr�i�6��	#H��u"O6���B�p���V�ĵ7>2\��"O��yU˧S�(��K�$�E7"Ox�[�S�(�%Y�9�\��"O���	�$]�(�!�($�4�a@"O�� ��/�~����)�¡��"O��U�ͰF'���!��R6"h�R"O�Ƀ䂟�z�X�@R�~;Ь0"O��*��S3)z�a�`[�)�	�!"O�	k/K�Bנ���R
B$2<a�"O y�%�'+X8�ZI0����Vh�<I�DV7z��#ʡdn<�!��Z�<��+O�er�*!IݜX�����o�Y�<��,ʊD�Ɔ�/v-���@@�<������ya&0�r�`��<Y�ƹ4'�ȶB®OS8M���Bt�<�iE�&���.6�A@��Yl�<y���EbP�;v��q'��;EO�m�<�Q٤H�aJ���,s}��+�P�<1�OF31Yꋁ; ���eYJ�<D�j��B���1�D%0cJ�I�<I�d͸ղ]�!�T�}C@@�v�{�<�p&Q�7���q�J�&((a��s�<���L�$MjP�.ެC72��UY�<ل I�u�8����Q�<�ܬ��'_W�<��
�ht��¢��@���SW��R�<!�9|�X䙤��(�f���%EP�<9�,oM� b�eƪR�.���B�<a#$P�c��,$�� a���V�O@�<Q�l��`KU!A�kVɸjN~�<��ٞk�2hQQ"�$���Bj�E�<��i�"5�^墵��U�>PH1��G�<��ՏU}��s�>>����0�E�<QT �� �xA��&��V4"�2gPD�<��	I�}���F*H1[�Y+�	�z�<�M���Lc�F�2%��|9��y�<��n
pnܱI ���*�)yT�@�<9��N�O�l��-@}��M��Ff�<i��P�� d�9]�8���`�a�<��,�2j�L���lx��FGE�<QV�&S��-�+�5p\4��'B[�<Ѧ��Sj��q�@�o���2�.]�<���D����Y,y'��%��r�<!��:<�l�`�U�S�x���K@C�<ɴ�̊v��B���r.����[X�<)�gF�:%v���Hݛ|�B�($Ǝz�<!*K.f�����j$40�I K�<!��J�[=x	%j��qF�&��E�<i��ԩ���`퉭y�&���	A�<�Q#�w���b�42�|�Qm�z�<� L�b ��>h]8uv��g�p�"O��7'm�Ry3���6I�dm��"O���uK�+�=��n$+�&��"OR5hQ~��ِ�n[g�R #�"Oސ��H��h��BM@� �~�c"OƤ�!j�+���4�;;�"O�$j%˗�W�� ��g�ƴd"O�q���I96��I3�K&����t"O��
2/�!��Q����2o)�]��"O�%B�Đ/����rDLuP1��"OR �D�У�������b�3A"O��[s�I�H{��P� ��"O�)���L�[�hҶ!��D&6�[�"O���3f%q�� �B�lj&0:"O�UY֊�].
�� �+��\T"O����P/U�J���� ����C"O`�ї�Η4d���L[�Cw9�F"O`�Q���:fb��J뗆=_Ʃ��"OB˱�[�aꨡ r�l(���"O:���i9d��ȃ�!XI�g"O�l1��K�}'f��W�"9X0k�"Or0Q刯Cd�)��5v���U"O�5��*S��h�'��t�Vx!�"O*��M�m��v%y�|!!�"O DN�9+�XI��L�'�̥�$"O��jE#�	���@qa�4p�C�'�ܡ��k�4$�����A"/�d���'Np󐬋��<��W���0��)h	�'O�MU̃"�ncv��:(����'2,�zֈ��<-X ���'OK�O�<ɰOL9f�	���'�h�0qk�M�<I'�� D�*��be��,���0�ZM�<�A�Ū`��uze`�>f�@x&��~�<�f�����ǆѶnR�t��n�e�<	g� ��]se�ܗhCf�b�<9uGU�)}��(�,[Nl䜸�l_�<I�F�M�bL�t�A��%����a�<a���%t���NJM+Va�#RW�<iӦ�7M�@Ȕ��Ι���y�<��)�s�*h�Ώ��Z��i�<��M�=\Ӧ�����r�J��d�<Q�K�-A4�,3!��1W�4U���h�<�&�/;=�ST�̫�<�R�eZ[�<�N�:F�	B�3$����#�X�<��.�*RY�C�5Oj8)8u-p�<���@�N�"��R��3ze9����Q�<)�n?��K�T.t�T�@+J�<Y�cܠ" R��"̈́�U,8R���`�<�u(��,dUa1�:<Rԁ���t�<1�ԘW&��N2�,�'L�m�<!4e2�*�Z���2x���ae�<�F�	�K���8nd�r�Ca�<A�s0:�K1#=Ҹ1#[�<��Ʌ+�{�dM$T�����[X�<9Ӧ��C��S2g�m�T�e��W�<���6&}x=I��M�Xph��J�<q��0h`����"9�.�s2�B�<9����^���.T%z��{6��<�'i��=�F�2@�p)���f�Z|�<��e�26���T�K#x$ib�s�<iB_�PY I*h�z(�W*Nl�<��.� bK��B����l��D�P�<��ѰA��¡�<7���P�I�<�ì�P)<ݱs�8X����ƫz�<� ���
a��)�D��#}�tA�"OFLz��T�@��q;0!ߨik���"O�I���G(h,Z=Y6�Dq���"O�M�3i3u�J��!�ӄ����"O�%�T��7j��l]8�^@� "O|����j�-����<6��D �"O�Py��RH�Sd)^����4"O�U��i�L�aB�ٴN��u�"O�`&B�ut�r&G>q�X�"O�X�i`~��%�}�>�sE"O��{�.�p�����d,�Py�1"O�hX� [&�Y�g��J�6�cd"O��9t��4� IR�?k�lr�"O��Aμ"ؠrCgE�hy�H"O��y��U�r�T`�b&ڂv��Ũ�"O������Q���Bv�2��B"O�Eq����n�D�*`�G�*�!�"O����R,L���cՆ�)\��!p�"O���%E���0e@��z1R�"O<��@-ĹxH��Ӷ�"b�����"O@II�ж\ٶ� �%�j`�"1"Ox�p��,dB��pO�}���s'"O��K��a�* ���C5�T�(�"O��5�J��ԁ��(� dە"O�$�d���RD�	�v�]�z���aT"O��D��x���0�+%��(q"O �R���10P[U)��8v�D,�y"i
��õ
^C�4t�C-���y����x2r�3l�n��@���y��8�2j�g�*�b�!�0�ybg�]U���G��*j�lA�i�	�ybM�8H�XI0��.��D��K�y��*E/�P���!��Õ)Ĺ�y��P�|�N0J����j�Y�6.��y�O	zS������D����y�БL09���Ӎo���3j�y���R�6%J�aU~X�E�+�y�aǏ����灙yc�=�!�"�yb�ٸS�h��A�;&�Tp3���yB#0"�Y�CL J��K���y2��=	V�*	!m����&X)�yBf1������r,�٩�.�=�yҨJKP�ya�Y�B�6�Z&�޵�y�O�g�d��D4|�`Kb��y��A�10��1���(�&yCƥΔ�y�j#2�R���
R�S�h��i�8�y��̞s��aS@mZ�F;���fR8�y2�_�kgri�bB�0�����i���yr�	*�΄z
�72Dư�5O5�yr��x�l�hSI�9�!qu$G�yb��-'���C�/I�;�B�t����yrI�ޘI�K&0�������y"o\9v-I���˥T�\9���
��y�휧�x(#d�N�Nu(53Q�yrf�[Ѻ�0�gL�LmJ���dՖ�y��^
��Y�Q@���� o�yb��|QLE
�'��`�b��y2EE4L(�y��s�H+a��
�y��Е��P�Hv9bl������y�f��
���C��,B���C�����y2�U�H�B��l�&�֐�7�F��y�$��"����<r���y�ʼq����h��b���g� �yB�Hm�<ra�+{mT��!¶�y
� ���6��X��	7/�T�0�"OT`�%Ɗ G�ܵ� Nܹr�dM��"O.	�a�gN���	����"O�%�I̛.���cP��nژ��f"Olxc�T39���z�F�+5�Ơ�F"O��B�`� ,Y�}�&�~�4 D"Oxy���ġR��x�Sz�8T�&"Oh�!#��D�QP�� a� �K"O�M��
���	����+F��0R"O�yp ���X�W/H�b��"O�Ș`�]�J+>�0��'<�k�"O�#���ݦi0��=A:�ݨ�"O����� 	e�����sV�]�"O��;1o^�EL�#j��IY�Ly`"O�(Z��A~s�Q�2���F�� "O�p�Q�5в-������֦!�$G�@phZB`B'�a�.Y�H!��M�$�hQ��ޢw�$z�B��!���!.$Qa.�R5�� ��L�8�!�$\9n�da���~����b��<�!�d�o����E/ ~�� 
��!�d��VN�1�(�{��c����!�_X�*	Ku�]9Z�jB�bt!�DD-%.ǅ��2���T��-v!��Z$���d[�u���&�L<[!�$T�	$��rl � ���%�*U!��Ќ:�)�5��70�l<��M@E!��t���#��~�ĐY�&۰T�!�D�qV�Ѓg��#S�̠c'#2!�_)o$��*��C�8J���`͑�E!�D�2��Aa��:1&�1W�=-�!�䚒3`�D���ʥp"��y'
 5�!�<C�-� �1;�՚��'IX!��%p��,
 �X%���Y�hE�d!�{���[�o]�f�Ą�(�4V!�D�gƤ��#9Y�p���=D!��%I8~1�Q���`�[Vn +.&!�ͅB��HK�Z�L�U!�ě�V���#�D\�Ku�N)�!�\��dc�&�:8��r���!��
����ӛsj8�!�$,!�D�Fd.i�H�U�^�1��10�!�d��
�ࢧ�ثx�R�OB!'�!��+� l����{���CĖX[!�32���Zd�� �L-!��30!�+m�:�`ä�!dҝ�G  7Q+!�Q�S���6�E��[��a{���6\h~A�E��R�H���J!�$�.�$�z�LU!U��Pj�(!�DC�.z,i�l�;:��ai��v��~�^���@9ѨP����9C���P��;ʓ��<	�k�-,�n�1�-��*R�a�u�<��D�r��8
���4e��aH�<�F)K�*;���゛LSn��e�C�	ןd��	 �1�䄟x�� �Ö;IC�I�(�!��������D��
b$#<)���?���,d��IC�j�����0D�4�$ćho6��&٠B��d$/D�$�rDʛG<}��g�:EcP��	+D�ċP/�?8W"�B�o�KRB9�4�<D���`<=P�qѰ��M$�C�{��C�	|?��{�m�j����b�1r#�͐��y�!_�Z�����h�j(�H{t�W���"�S��|��K$���Q1Ǟ4�<��E��y
� b4�1�9y�tj�
�!�Ԝ�""Oΰ���Q�fܔ�W���i9��	T�OO9�te޿�2ԩVhJ	~��)�:O�7�?�O� ����W�R�ĉڣ"O�ܩ#*͏Yu؁ !Žm񑅹i\�'�`�����E�P4Y!�9#�TH�'��B��r[F�2�f5r��H�'�\�P��7E\�"�)��- ����'��b�oS�%�ܑ׫ޟy���'@8�K�NL	X@�� p爵r4~�;�'���a� F��Q''ɨ�,}՚�8�'����Y��� �2;��
f�W��
G)2D��)CG�8}��ِ�}��/D�<a�W� ������؎����*.\O�b�� u�ύ@�RH:�Mđ,��qi�g'D�0��Q��M!�$��OQt���8��hO��¸�cL̂^�} �nU�,�hC�ɜ6<�;Agʹ2��� c�Fp��dE{J?i9E�׵|�t�u�	�!"�raG*D�{1nޝH�
���Ƅt1U���Gm�'@T�D�,O��YgŊe � �AF2jv�� ��"��?���:杒�@VM��3�Ǝ�D�~\��j�2}z��L6a}ܱC��M9\6�ԇ�8n��1��Qx\���(SX=���ȓ5���"�܀��ɒ� �#[�B0Gxb�>�M~Z�'���a��$5FNةT ��O��"-O^���*�h-�g�<'v�q1Fڀ:�	C�'��6�	MsPS�/G�+���@C�%:�6B�	�\�P�����5�����wr�	���?я��\� �"R��Ӗ x�K�p�!�@$@l�̛�"�h�\��eL�k�!���O�Ya%�T���ӡɛuO�'��@�<�a�=_@Є�N�PGAK�< �͂}*T '֧'/I8w$�I�< ���9���N����*D�'�ў�r�'���R7
E&d�JL�"cB	Q1�0K>����F�!��9�*L��`q��+N!�Z�3��O�i��O:8�!���[��B�䝧{��58a��k���=�O(�HT ?(�""��5��<�"OƘ�"-T5NA����=e�Hyq�"O�b@Œ�7��(C��2GD��ѳ"O\)�b�A�,�������)1�406�$,�S��*
fܫp��:U(8(��:��B�	�o����)BY&(���^�*�PC�	/x6N�fh܈.Rx�_�q�
C䉓aĊ�mۘs�>� ቉�o�B�	Kj�\�@M�u{b����"c�B�ɚ93�����X���i#�p�j��D&�_��1daK�F�y�Q�G�WF:$���|,�P "?����M+q�R�ȓJHa�f�V�y(���e��;�t��e]��k�!�(d��ي��$1>�Γ��?	��Z}���c-(!WD��1,�i}�'��2��O4[�h`�w.%�����'X�Azd���_�y{W���� `��'ӄ4q��n��[bK?s\JqO�̱`CZ#�XY��BX��<e��O�ذ"H]D�\YZv�I���q�!�Q|�<�d�\�F�tH�ȗ4ռ�V*ZO�'��x���}wd�B¢ب!�RU8�'�M�	�'�r��B�p��%�d�> �FUY��<,O&X �J�
$�e���+(�x�"O(pidu����'�~L!Ӓ"O� d�itM�:9��9k��Vf�Rl�4�	h̓��O�j9c�Z�u��} &��8t���Q�'�eCrH�;� k�4q|���ӓ��'��X���Y����n)`0y�'�P���Ǌ5${A�ؐa��`�'�l�(�
%Z�^i@���e��`S
�'���C'��^��3�	�Y�,�H>������!�V�K +!��;��i�!��77�������`�A��_�4�!�$�$Z�n��W��"C���9�ŉ+ps!��#`�0AG�(<�V�+Ez!�䈘N~Vi"�Z?�,X �4y!��v��' �9X���6��$w!�.�v hg�ĲqG$Dc�BH K�����,<O����-oX���C&)$Q��I�#�'1��/\�u�@С� �s�e�ȓ3=�(����&Hڠ�s�HKP$�Ez��ieў���X��L��0�r���ӹ|h!��C���a�-I�qs� P�nXP��=訉�Q='�I抑�#D؅뉓��M��_�&�%�")B�=0P�s4�HV��8�O���f�%,.�@��a��ޢ����d.�S��,��j��}��d��,r�m�I�#|BB�	�(�"ĒƊF!~`HkaLI�f�~B�ɼؔm��(��T��� ^�C�	���c��un:�
�a�
���D𑞢|��͐a����vh�JP2HաQ�!��C�(pnp�@՝j͠�
C�Y�x��'���6�S�ĨQ�3�L}"����	�@�y5�Š�y���kؔ@S�׆	W�X�7��1�Py2%.`�I(�G�Xyz ���܈5�6�FyZw���у�-���]Δ�p��ޚ�Py�i�)Kv��#�@�MO����D��y"��#,O*��d�E�$sDq���R(��8��'�@O���d����1À��V��X4��,LO�8S@m�+*)��爪1��3��_����۽i� �Qc�3+d(��uh�&a!�D�%D��MH���>7Hʁ ""�+lԠ���)�矀a�%�f!��7h�0�(��E���wh 9�#�%z�xL`d�7mn���	b�I�km4�i�n��aS�fږp�B��>���d%���V�%O�K�L�<�'�ayR����S� �R-��aP:Z�XP*�'bJ���2-��	�УQ���'���0`a����]�F��F��	���*�z�Ҕ��Ň"4iV�V�T�<��Vl~�2	�)�4�@ �S�r�ȓ^2��I`@��H��!8;6��ȓ9�����⎤1 z#�2F�X��x	�Tʲ��4a >d�π�2눨�ȓK,�� �O�'����rȄ�{5\`��F����K[�����.>d������~���#����i�ȓd�2}S��-2��!Ñg	�Z�ȇ�<t��)CD[;NCڀ����>y���<f�lx���:�칒g�8D��=�ȓ	��XQ���Nf}plW�E�����p���XfR0f�6�be;܄���]klɊ�"����l:��Q3
6��ȓe�=�E�"�2�o��d��!�ȓ�t��ZIx,��-u-�-��pٸ��"1@�"��~���ȓz��S�L�/4� ��,یY��ȓ`sd�	ĦG$�0B7c"~_�p��S�? Z$9���cY�e�P&�/iz℁�"O��8�ڕO�X�X��(c��-a�"O��1�ݱ>+%�׫ٱl��A8�"OT����9��I+u���C�@mU"OR	pG�MA ��"*Ȣ �*��"O>���dƗ �����c�5C�6��A"OJ�h�/F�V��H�� ��@kD�"O>0��-�+Et=a�J.A��L�t"OB�c3�E
�& �p�H�v4��"O<K Y/,�^��C��_I\���"O\(�����;�JT��&�:Q%�H�"O����U�#ĕ!��U6�s"O\��I�j��Z��B�?8�"O4�ab�_�g�tp
�>Z�l�"O�i �H�D!
!K�� (R8��G"O����+C .�N��1,��zʀ�"O�@+��lmq� H�o-�d"O����Dm!3�0����D8,!�E�r8z0�ul��,Kw�J�|NxQwCƠZ�x��1sXaz�^ܚ,��D�KΓ`
���y?Pa��h�u��Y�,{�ȓ)g��IUa�*yϢ8#��5a�r���ɾ堄�2v�jeg�6B�����c\��	��È�H���HY.%����K�"����ʘ����D��G ���i�fQ��\�#~-�S$��<�ȓVy��Jv#��x���㋌�P^T���. vh�g��>emHT����k��$�ȓD�b�-U�ȱ0r@�ņȓ!�����%��=�ԂȂ'����1��K�"1>�8��T�+{RT�ȓ%���B�X
�6aH?L쾙�ȓy���B�[4K��6nM���!��'�l��ҬG�+ʸq���b��Q�ȓ&'�� �zy" 	K��K����ȓUqPЭrglځ	�&���}cBX�WNS�(�
"�M 6�ȓK��	�a�	w���ꐣ�L`��ȓݠ������`�iƈ| z9�ȓzd�-����O����҂U¹��b��1�B!Bg�hY�N�#K&�B䉈hXƀ����.��i�F�.s�C�ɓ(��ep"ʇ<N���bF$"� B�	$-���DݯBU޴�'ř��C��1��I��"^�.��G,��"�C��--��=�W�����c�GDPB�	'���2tJ��$H �GbN!hC�I3ª�xbn��$	��N�'0C�	?z�((৒�bh~("���IC��*N����PnœO�H��U8
&�B�	,`��	&%�#�N�@��+ �C��#J���t �`�a�΂�cy&C�%d����"n�퐨�E�C�	)Qs*ƋOFj�;���U��B�	�5?΍"�J(� ��ma��B�3R���)p����b��"O��I,
�hݔ��!�3Y����"OF���ϊ�1^*��3F���%"O*a1q�aֆ���fQ!��TI�"O ����:.��b��8�V4�"Ox�
b�>Y�4����V H�"O~h��F�:Ɲ#���?Q���"O���FK��S��*r�ƎJ"����"O���ȏe
j�Wo�:ż��T;O��p��&�)�g�? `��6�G+ �Dxz���,c'���"O�CV�\(eѰ�F�� �`S^��	4�[�ka{�b�\�t�(VF��a$9`g-B��>A�C:.P7��1�ʰpCA#�L���CF�)]!�D$�l@����^�>��sA��C�ў�Cѩ��T�>���OM,P�# \�|����wE:D��i�iT>��Sf�?EQ��Z�)�ON�qPCO�丧��Fqp�#Yr�h����ź'�f=��f,D�x�w�D�y����C͂1 �Py�i�<�7.ϴÄ��� e��Xa��4|������#/9a~⊑�l���鸗dΙ}�$,-X�A��3��	R�"P�s�� �H�D�d���0T�ɱs�P 9όep�!��2�����e;C�ۈex�1�æ[�r��܆��J�k�˅#)ʨ�V5	���ȓ!N`�Šܠ~�ʈ� ��-W�2��ȓ2oJ��7��o����qIʗ,������X@DK����.�q�h�ȓ�|y���$������� J��̄���тKUW�2`�cϙp&�؄�y�0�����"a���"��=����	��[F*	Q� 3&v����W,��"�Y
p�l"0�,<�q����g@��@.p-��F�N;Du��l5� !?}����v��v-����M	���LCN,��)���J�H`q�DQP�)���,|\�u��z&P%!D��ZL��D��	ڊ�ȓF��ˆP���mӱą'���ȓ�"�����r� kq�5p���ȓ\�rLI�M�z��0���c�H͆ȓ,\t�B�ȑD�X2�БZ@2(��E9`h�R�?hĪTH�"�Y��l����ȹd�����Ə�y��M���ř+��\��P�(�d`<)�ȓ�8�I���*`F��� Ԇ0k*|��?0��2�`ܦdX�HRnۦ�z)�ȓk����g�:�\���/��#�����N-�����0!�0J�Gp�0�ȓ:eE!�$���`��,N>��ȓ/��=m��M#B\[dB��J�z-`�'i^�X��X�Z����Sf^�>R��'k�<�Q T!y�0��O�(F$��'����&(o�$�-ȹ'��-P�'�Ѕ�Тv��l93����4#�'R$D���0�� z� Bjd)�'�X�yq]�b!
X{�h�F����'��Y����R.@����J��١
�'.raB���w� aQ���q���9
�'�u��Nւ;�N1��űt�h��'=*�kP���s���;���u�<C	�'����7���b�Йx�F�`)����'xVa�D��9h�p�#ê��/���	�'5&hI��"hdy�Q�*r�<Bq#�u��(�Q��q�H%�g~RD�x��e�D�W���5b����x��<�����(�Bia�\ |�t ����<��A�ri��z2�Ǉ���:�I�'Hʽ
�MV��p<��ԧ,�|0	��6[������k�xlQ'M�9��V��� B䉶&�ȱ�P/Z%2U��k�*g���^�Nl��g�#W�F���A�8��	�]w�(����``�-<� �`�B�1}X`��'���h`P"N%΄!���/��+�u�=�4"�`Xd��R�H8#UH�p��t�x�	�z&�r"@8��P1�ƛd����$���&��2&�^���x����O�@X�_6Yb>�+��;ft�Ô����u��C~8�x㓏�s�a��#L�(	�BǢ2?��������>[�ƕ�I�3Ƭ80��݊I���� l"7E8�; ��?oxLsu�@&c!!�d�7)�*Qr�HTz�\!r,���;E�j�[�
Ȑg���85�Z^�$�kdJ�=��W?�k�Ì�D�4��n��#��O$D�d�P��y�>y �F�?W�d�yQ�4�~Y�G�l�C���-�d�@ޟ>�P�Hߪt��ʓP�
�3fW�x��$L��7k���퉸�y�&M��X��_�RU ��)Ñ)��H(��\��qx�E��.�&8�«@]�9�@�>�]^��2?^�8A2��4rb��?��'�� �w	Ŭgv�!2ׅl���!+���m��P�7db�Ka^�^�x�@�NQ����z���)���r�YfJ�]S�ڐ|�(���V�`���e	�!ѷ����v�QN?)�sJR��MAr��uB9!�+D���%o	�"]��+�$���<#���\���Kb��>WH4-�.!4(��y��pj���CjR��c�������9R�؂G+O[l���K�/33EM[O�X���~����V^1NDkB�P��h@���-<b��U�Ĵ'�Q����C�m�Je"�-�8L�#�r�v��-\+(iT��B%�O��Ix�����Eu�5y�$�(޸Eن��L�R��`g=�On� jJ����$'��G@(y�A>O��9��J�Hz �!�$�t���JK����g����� �FE0f�J�l�|���UޞC�ɹ0T��e�[smⰫ�!R&J�:��ㄹY�i�F;+4I��)"zR.uS�$O���ǶK}����2k:%HcgE�ta~�BW;9�A�#��\���=�xP��o1>I�� �NT>Ӓ���8����D�O�'�>��-��i�<���>j����$\�T>���E�Յ2P��s�8�]hŃ�J�b���Pt6�PP!.�� �Ƭ�p?��哟wU$ ��$�O"���#��<qw%]O�0��B�	;�Q��s](4��DO�O!��O�����Ç;f��9�i��3^Ĥ9�'�j}E�Ƭ [����� �b%����Ux�B �\�]�)�O���I˸#�
�s�_��~����^y�m2
_Q�. �1NA�p?Yp�F�?v��G��حPkU;Z�Zd�v�:#z��;��1�F���,E7m�J�#��ɓ.���3/(Ab\ݱs&Ef7�>��ɋ91�(�"T&�8`\�X�N,���@d��VJ�x u�,���JEB�9{��'7������3�B�㮙�6
=Q�'�X893N�8�1[S@�&1���	�F��g��'Zf��Q�F�?�.�����=Z����I�<���+�>���U&m̄�)���0Q�D����	y�R}��؞@O��#�I5{��$?�3�'��I�)�E��4;����g�1}m>���j<3TlD��B�:a�\(�A��8r$��d�-I(��pi����둡G�K�Ђ�2OT"?��S�m��h��&Ő!�@?] ��|f�}b�ƫY6X�p���2 ��Љ.X��(��ʪ-�� �p�S�k��C�	���*F印k�>���l*���Z�k*g_����	� �����*��z����O����᜛��$:�lLE�n�A�2��Kc�������`��6�R:D~%p�Q<H����@K�:or(˓G�"�F��O� �4֭h"fMX��4=�8����Z�n�|��e �f��0��j��DQ�X1`�n� ӵ��V�Z���&옋��<���W�a(@�'��R xe{A�V�*Vb� &�|rC�j�3�F��ƂF,T\��)YS�B�D�]'0ה�t���񤒑NkRe�
�6<�#��v*���դU����0��Y*@�Mn^IR-O�O���ä/�t�`=ȰaI�Ok���ۓ<0Q�ɍW}ҋSJ
�yr3d��)�z8jT�[��y2h�%����`ה9@���T��O����'0����y�ԉM�m� ۞H�Q��`���L:����7!VT�rń�+��В�ˉ$_V	B��4c+p ��^, ��C�ݐ4Bf�ղ]����K��];S�\.|����.���ȓw��8p�
B9��g�"X�\�ȓ x����=ƍ�-�4(N݄�p����NȰ_#�qI+�?7ތ�ȓ[N��ۤ)�4��@��J�nHhȇ�L��0�A�bT@&D0Cy�$��:wp�I���.K󾩳Se�
]Q���'�ք2W`T�aY�����0{���(t$lB�D���Y��G�\˞�ȓr�I�Ƈ�V�d������9��_�L��#� �n����eG� �ȓ*J,�&͈$��'�-b��ȓd���Ӕ��(@� P{�͟�w��0��S�? �ͳFbE�[��}v��dY���"O��[�LP1c؍�V�'��:a"On5�JV�"���7���N*,l0%"O|� �I��	L3�/��*z�%Xb"O>��#��!=�ƨ��R�va��"O��`4f��|B­�Vl�of���q"O6E#�ʐ�
= !���SM�	�"O��j��C�Z�����ׄn�l��"OX�Z�M�
!���3��9�lX�"O��6ʒx� @DK�1��iu"O�A���[F�09t+�-�I��"On��m�]["��D�L�\�pI��"O���
/Tv=IvfVúI�D"OX�B�ա4
�y���$dߔQ��"O�:pB&[x(0��|��Dғ"OV�{cJ�{�qY�kο<�"���"OU�f��P�TE[�-�
n�>�i�"O��+� ǀ[��8��-%��:�"O0�+�
�?Lze:AM�M���u"O\�6��^���-ېz��e��"Oh-���E:fy(%t��r���"OJ5+"m�Cnr���V�-�x�<	��6��\�2*��B���Zfj�]�<!TGȕH!x�$������Ӣ��_�<!��'H����w�
+z�it&s�<�d*G�$��\�S`��=�&}�!��b�<A�������ƽ0љ���a�<��������	4��QƧ�z�<�T��I�)p�(�^ABqYg�r�<a�*F&U!@�@� So���2�l�<q��˳b�L@(+(F����h�<���-x��5)�,E8����Ŝg�<A�� ��t)��D��s�NIc�<�J� 56�Wf�s���c�B�^�<��䔮g.�4�P�qOj�K�b�Z�<���9e�x�df�Y�ZQ���Q�<ɠ�d���8\�8<��iߩCa�B�I3X��DBќh%���UC�ۜB�ɫ#ƒ�:���g��u1���NB�Ira� HW�&:H��1�G�+� B�ɷ\��b��Q����6LQ�w!�B�[)Fq�b��m�1X�A�9S��B�I��I���:$��d
�,	�C䉱?j	�VI@�+�&=+�
¢C�Ɂu��DQ�E��J& -z�
\uNbB�	�LRl��J��L��I,fB�	/;B��G�O�'x��s�O���C�I�l��X#��U���;��ݳz�C�I�F�dh��LN��1^�ix�C�	�L�!ӲFJ�m�릂
0w�@B�I�n��UR���N3�-��B]�r�fB�I
�(j��چ(�z`!7똕b�~B�X�}끏�rĘ(�u�'N8�C�I�i[�pxrLVxKZ0�
N 8C��#At�i�@�̧=StY�b	�(�C䉛���h�F�C`�[p��:T�B�1xt�(0%���Y;�Lx�ż��C�	�	�j��G"0���q���9�hC�I�RS�ͻ���h�
�a�>t-&C�W�RթԎ+
o��hw��,t�lC�I�Wi"�ZD3o&�X�����&C�ɦ?Ұa�c`F�zz�X eZ�W�.C�$T�9QĖE-���g�n0C�ɦ�@T�'f�d���2A.@�6=NB�)� n����$�`��㐒7��`�"O|�9 ,�!k$��3��Q�:�&t�"O$	+2�Y�8B���n��e�'"O<I���uB$��색2����v"O�e#���P	f,�	N��9�"O����E�:"Ն���I_���zS"O� J�)�.�0�c����}���A�"Of�1I�Z��T�9J֎1h�"O�
g�I�p;���3M����t	�"OX8bv�U�=ȒL9���1/�Y�"O�L+���'.N�)�N�ZŊR"ORd�.B�/R(1���� ��,j�"O���O�r:�d�Dǰ���"O�d0�F�<G�b�f�j�4"O�Ixp �[�����Q��$"O ��(-$��·G$���C"O�h���0�Zpj��^��x�t"O8��A�hY�Y@�]6.�H�"O��c�CO���r�U�]ԙ�s"O�]ҒA��t0 `$�'4	�U��"O��1��]�#9�\r�dR�d�Bxa"O�tb1#
(֝H���<<�"O��`f�,3�m��%�.Ŝ��"O�5����.K��A`<��R�"O^k�$P����S��T���Z�"O�%���;�YA��[?LV���"O$	Z#3���ABL�i*:]��"O�ͺ�o��4^�b��&Ft4���"O�����y�JS@A  =�x�B"O
yd��!N�"�A��m.��c�"OԄ K�b�<]��@�C	H��E"O�!��)ea^RW�	�%��"O��w�=@����
�{�*Yb�"OJ�"V "y��kTK��C�l�0"O�huaU�9�A�VI/Ǫt@�"OV�Dϛ�.���A`��s��p�"O
I��K^
�&�R!E9e�!s�"O<�Cd�`,���R �ҡx�"Ob�+�Fƛ0BL�"΋ %pő�"O�!��J%F��pԇ$>�"w"O�	��Ȧ5ch�+�!�/2h� ��"O"��� E�ҊT�r=���d"O�U�8���y�nN� 0���"O�X�⎎)�H�b�L�J"�$+�"Ot�4+�H�p��˯t(��$"O��t��a-)10hraK�<�y��/(M���U5P��ٓ샟�y�B�<i=�͓GE�G��ɱ�#�-�yR�!@�2�a�0T٨f�^,�yR-����Mȡ 
#q`l]:#�ڦ�y� �T��P���*iI@�
�&��y�a1:;� �Qo-��k���yB"�r���0�!N@��H�>�y�ʎ�UC8��p�A���/�y�DSh�0	�$NY��YBƪ�-�yb����aA�/��)�uҮ���y�g�!2�9K�"�X�Ӓ�y��
�0�x ���)��������y'�*�n��;���3O�/tf!��Z�w,`�% �W�~h�`-�'G!��0��Q�ŗ*-�&�f��;J!�DA�
��L�$h�0p�e�w���O,!���09q�	�kضOc�pҀ��i!�����sNZ�I���:��^�&I!�� |����ȯgӢ���G�`���"O0I�#A�PB|aç�<r��Aj�"O�4+��ܲ, I곃�
w� ��"O2%C�m�J�^�����36� �a "Ofp3���^j��&�<%�y�3"O�Y2����b����>5QY�"Or�񐎘3]�<�5j��0� i`"Otщ�Âc��X�	z�208�"O���#ԓ?x�䯌!6�-1�"O"�Q��@O"��6�$����#"O}y���	������������"O(����X�kn�� �@����a"O8��5��f3�����O�o�,1��"O�萊�_�$s�jM*j���5"O�=S֮_(��}�q��(���5"O���`�rP�W�U�<�a"OD0���ڭ�l(�E���7�=f"O� '�F�Bv���4��O����"O6,{�kٞB\�M`c���_�A�"O�,�a�C>���k� U�7����"O�@1�I��U:�@Z0���"O�Ѫ1OR�a4��E�z��cF"O������.i��gCK37��J1"O��Sᖇ	�9
���|	���"O�Y�
�Jhp����%Yn�D
"O� h(�8't�-q��&HBe2P"O�%YF<\�8y���/@u�"O���Q��k����Fխt� �"O�Q�'�>F���hĦN\((w"O@ p���>vz��d�_�G t�f"Ob�e�Y�{m�[W��.��Q�"O�Pѭ�6<��ѵ�ďN���"O�qsw���� �"͕}�0��"OԜ��ʚ
<u w�]ߚX0$2O���c� �OJx�b��o`(5��K�#A���b�'x=KT���DM�
=��!�O�Q��Q3�`P<<�!��T4D��.��τ�����o�qO�ݹ��5P��#jr�ߐHc�x1�FB/)g�<"�.�e�<q�J�vH0�+v�J�#����J_�2�*�Qǔ|Ҫ�]���#e�鐀B['���W.dU!��xvD�B3n�{��L�AX��ק��1�X]��	
U"@#F�=
t�KÍI6j����@��l[��>�#6lFE��@�K&(!�a�y�<�Ä
�> �չ�@]��xy&�q�I|� �V���ȟ��Ҭ�*}��U{r)U	3�!�"O�x�aLS�}.@�r�)�(��IM��:E'�����<1��-j�z֎+|�$(
��g�<��E�5������ϓ[�t�9P�̞Z�Zc�/H�a}�(��F�p4�gE�'����s����=9��?px$��'�bl���+�`�	Am��4�jh�
�'�pfn��Ѻ ��(,�r���A�BM�d�(r���KROD	#�T]PqDW�<I%�)#�*�!\
\�~9��k�o�<1�ɳ*�R�Iu��?뾴�v�i�<0�Ųo���P�hA/up��P^�<�r�F�bb��a�	ux��ZV�c�<IpI�/�z�s�(�2L�8���N\�<i�"�9؊��d Y�<!,�ӳ�p�<�Ƭ�����"/t�N4�$�^T�<� �"~�LTwǇA;@9���W�<���]A8E�fLr^8���K�<)�(�<�>� ���`�
��)�s�<i��)�̙��hK�B� ��T��f�<��/�0R� �Ñ+s|F��"�f�<�  a��g[s��3C$@h(��"O��*��O�h��۳ɞ79�䅣�"O��ۆO5`L�u����x�|��e"O���DG�n��<cFI$D��eP�"Od]B�E�{"�= wj	�ƌ�"O�����J�R����L�Fr�cd"O�5(2�ϰ2����LQT�Q�"O:!$e�;:y�,*�B
-�
��f"O���H�s3܈�@��!o�x�Ѓ"Oz��B�q��$a��~�AK "O|5m��E@�G�F�z�C�"OvɗhZ�3��Q�aE؇F����"O�xAѡBkH03���/M(��"Ol��͐$���m�!]`k "O�`�d&�)aj����+Bz4�"O����C��h��!�7�ӕ<g`���"Or �T�J�oJe[�M5F���"O������ �C��7�`�"O�j��0b �%q�NX4$>D��"O��$��� ���k֍X�ʀ�"O�QLX�'�1zKءH�<� V"OX8AF��?����%
�/(��ؚP"OnB���}Ll�`h�3���Z#"O���o�	z`�����S �=P"Oz�k���P��R 5AV��bA"O���,˔	�V,�ĈG�4���"O��� ��pfPb�ܭt(�m���ݽ{w��&ae��2w�'`����� PT �����h�ߓ��'����V+E����ゎ	/A���+O�=E��CC�pw�M2c*�3>y�Ш�?�����+�|��-�E7��0�!M
<J �=�çA�X�wAR�|��DV��G�5�?���i�9��H��V9�}1��Z� )���'xPb�9�=O��	4Nɧ�������J"IK��ВD�*;<��e^�LR�D$ʓ�O��/�*TCn@H�� �ԑp�'�ў�~6,�!
T��*�^���m�'�a�d
������%L�,������'ў�O�����'��#��e��⅋��QɌy��'��T"��Tk�Hz�H q���9K$���@�b�{G"��?���Bz�SI?��J�6N�1�`],!L6��F�׹��O��>1���Q�BQ��"�tu�"��H�'"a�� ��X����$MMi�c����'�ў�Oe,Ͳ&��6J��4�C��@٠��M>�����B�+R�U���ҤW]���M�*��F�'(�|�Aiʤd�t	3eT8vmpyrA��O�H�����O����K�L1¥Y�d���`退Dz$$��T"2�2�+��Y>�p��+�S��I�+�}������a�SG�'�ў�>�����=�l8�'Ձsw��23ê<����Ӈ^~8!�%��%�,�[����v��3���f����!��<!�<�7�*�a��Ea�hL-�j�R聣x��D�1�����+p�Z�0 n!_Z!�d��L�Y��疴Zl-#/	1S!�dB�9�����]�P�D���W�P<!�4RqV��s` �kF 4�h�1[-!�䂗fh\��u�΁ -0���M�"+!�D@�#���򇚕&��cBl ��!�<n�Vi���̧j�X%� �(Jj!�$�Y"
X04ٌ}��W�,�!�N'֬Hrΐtw��K0,�\�!��x{,�yCjG� n�HH�¬�!�dѢ4�捫QA\�nW0���C˫!�d�) �=	b��^p2�Y�b�=rJ!�Dȏ���%OO+m�؆�5R!�� �󇇐�o�޽c��kª��"O�}b1���6�	R�U0�"Ozy���d�����K�5�ĳ�"O(��q	@<���{�Nǚf�@C"OjH�-C~]�1`��݅,�\ �"Ox���	"$�n��U��Q�\���"O���̜�;Bh�vؼy��"O��D�YW�d0Ŗ�"$�Ӵ"O��l�i�P2��`	��C�"Oz�'EI4������2�<x�R"O2��:�d)�r�����z�"O|̓"*R�'\4�z����d�"O��:�D�+T�(�c�5݈�@"OLP�a��9K	"�HPDHs����"O����mV�7=�dR7��bM��Xc"O�[�L�� ���o���!�"O��x�,�H���C�
�H��b"O���0g
�n-� ���%��U�v"ORTr҆��P a`Ӆ��E����"O��dK�'}��{��٦o����"OB����X+KU"�H�dMj]��"O��x�Y<I�~����3pAz �"O����k�E� �ɻ!���0"Of(x���9��X��^�A[�m� "Oެ�s����T C��o���a"O�
��*v��q&�N����S�"O$A���>\��W���r�@;6"OD(�Q͖�څ@�c�%U��\��"O�	@���J�N-��)��"dqS"O~��m|P�p/Uy�̡	1"OB��C06��4rOH�*��<`"O���hU�A���Kܤe��"Ob�p�ΔF2�`�o>��a�"O�]I&�S�XD	U�G�K�> У"O��b�Z���s&�Ñ��	ؠ"O�X� �@�Kv���4��Tz�P�"O^�s䫖�s�8Q��!+��9�"O�죗�Ä3@�i�S�].H�2"O ز�^�^򰈐�G�A���{�"O�ےg��`�����Vv�|�"O"��f�+�&�Q&\�!����g"O��i�n��S� )#�>�^���"Oj��&gW�i	5�m�޵�#"Ol���A�2`�������j���'��@9��+*x	� �I,�4���'��,�!�ўjKxd[u*�.&X(`�'ZR'��&��M�B�V�y�'����jW�A��B1V����'�M���Y#!,P���!R ��'O>��p@X�|�4S櫍�3�y��'{��{N�
T̀�u�V����'w2��2HG:f�H�s�FXl��'��q	�
CF�ч�ۈ?K��q	�'��ys�AR5C��$+G��3�L�b	�'u���V �4bX2-�SO�* 6m��'�����],X���/��pfI��'�:�:��'Z�<��b��2k���:�'4n �Eo�p����Z(����'�� yǩ07���A@�ƁC����'�v$���ͬ4� ��j^ �ЙR	�' ��%ܾ3��q'��I܀ Z�'��"v.U�OJ�����'Eg�y�'�b<�'źH���μ5�\�	�'��-�rk�A�Lc�'��
�	��� ��S5X:���	ցZ�~ L,B�"O�q��L�}���d���\�[v"O�PDK��O�v����o��(�"O���Q��wj�$)`L/$�p`:�"ON�[���g6��H�O���Nԫ�"ON�a֡H�7��=�A?����S"O���G��#bi�A�;^/����"Ox��6mS�d�|�atO�*d�<�"O>TK��ח��l���&א��T"Onl[�A�c0dk5��:l����"O�;�( ̸��5
����T"O���&L@ =(u��i/�4\��"Ox!��N��Q���k��ݾJ�X��"O��ƥ
=n�8���3椨�"O���C��$����1�֜5j�"O�ə�#D�N�R�)�hA""W�-x3"O騵H��2���t�]�Lu��"O}��h�1zU&���e+PԢ��"Oj�9�%��H�,\s���?d�x%"On Qu+���L8i��LC�"O�)񌙒]ZB�e
Ɨ_�!0�"ObP�����H�X�h�>M��$"O��"�bC������6�Ie"OnA���8��;�Y
�:�x5"O��`DiT.?�Kڼf�8���߰�yB��{����ÎJ&aiRQp&�ְ�y��W^�4��W��(��y�ɻ�ybh��'���P��H��x59��A��y2LL=:�Жm��ܒc��y� ��;��ܐ �8�nI�w�#�yҋÕp6es�d�������y�HU6J���z�����=E�:�y"��j3A@�)=� fK\�PʮB�I�:���N�$��S�r�XC�I�r(�P�P�-3����!�+o8C�T��H"B��\D��i%�1�'���B�@�C4T84%Ѭe����'���i�*�V���e^<cUL@��'�x��'799B���ӂ^�L`�
�'�.hp"/B�l`8���*z*��
�'!����IM�D8�8�n�.��M�
�'��\�^�RT�Fn�>`G���%��yƤX琈ؤ�v��U��y��=מC��B�k���rb^��y5?2���dD�p��`RW$��y2�]�cf�.I��4%���لȓc��H�H &wS.��흮������{���y��z�AW�R�������O!�$�C�f=���D!vD1b�F"!򤉾8�Us��Y�]{�I��+��f�!�mc���g(�h���X �C�	�0���k�<+� ���ٺbpC�ɖ{��+k�7���u��H�HC䉙'�$ ��� $����%*�$C�I*a����a.�"�lY�E`X�U�C�ɝC��� ��`G� ��`nB�	^v�7N	<w��*�e�qB�I[rU(tƋ����,�	s�HB䉰J>�x�D�U4+��Y#��Q�|sB�		�V,��+SX����ڹEcC䉉~�5@ �$e!~1z%,�2:��B�9%��arJ͚v�x�SQMػXC��W�� D�99ar��,�',��B䉫MV�p�F�W�E;P��#,��?X�B�)� ��Ѥ�J]�� !�!j<��"O���rə�m��x��Rl*�2"O�u �� ^�|!�����v�C�"O�p��t2)A��U�-r��2"O�b��E7"4(Q*_�iz^���*OԽ�b��X�E	��0���'������)Rܚ��7C	�;? �0�'K	H�7z�(�"�f�G>�l��'�����-�J��KȚ4�:5��'_��2�lϤQ�v�X�m��,�=y�'=�����(_<l('K
eUE��'^����>S�\ 2��!d�<��'aZ	Æd��.LTQ� *D�T�d���'a�P�\(j�YI` ն"�t`�'�������0!�̙#!�x`��'�n��T�<	-�ݑf�[�EҠA�''4�xW�Z�q'�	@%�<���'�������^w��!�L��/��! �'ޠi�B��p� :!ʍ� }�T�'�d�J�]�0>�c��΋SӴx��y�he��2H�)kt�=Y�Nx�ȓGvmV��;�0�8�+ŷWi*)��.Z�TR �D�}H"�P��
3H��h�ȓ?ذ�p��H�-���0��.4�$T������&^�uQZ-a�.X-Vd����+�v$�3�C���A�T�Y{g���ȓ�j|���ݎ�D�ŧM�H�v��TE�	BS�G1.%8�(�-|y��'��0���5���#f�V�T�� /@���+=�F�����aw�y�ȓ�x �����a��`�q/�pd�ȓ���S��!S���Ѱ"�'�	���ȱP��=Z�Rw�ͻ��8��Bg��:h�#��@�&�ҵ8����ȓ�B�`���)#"u��B(� ч����)��B�G�,bA��"c*���g?�9BdJT�SY�$��GU]"����a�Er�oZ�@��M�d�O>����L��d��K�|���>ṅֶȓr(���̸HA��ҥ7x���>�~ܹ'�ؔglx�8S�2;�Ḧ́ȓQ�|��	�*����(�̘u�� P.:�c�C�X!,}Ⅽ�G�<��i[=l�z�{1�Ǘ\�Z4��ml�<	���3nu*|؃��)Tn�a�#�M�<1���):���K�F����O�<�r�S' �&�����v����e�EJ�<d��;R}�]�Cb�E�X�R �CO�<9�!\d���ʏB�b�
�-�J�<鰪��K�p1��D���B�<����[u�1��B�g˺��2��g�<�M�1h�T)���#�lp�A�m�<IW�(^n�9k��z�#�c�N�<iD�R4PԪB��9Gz�cd�M�<�p^�D4�I9�a��Z5<��NVB�<0i��PtUz�����|�<���   �hB�z0�ȓ(ꮝ��@�_� M�L�n�A�ȓg�����*������%�br1��y n��Nڌڔ�
�-�W ��ȓP��k�d��_%�У5a��� ��ȓhT�AE@�(vT����P_�<�ȓ/����r�
:m �pt��}n�@��I�8�f�]C ��q&%aR��ȓ<�0��"̀�p�ƥ`w"PK���ȓN��
V'ӄX�&X�'��>����8VF��O�Px�Шe��?S����v	���EƢo��m��kK�Y����ȓS.���a�\(��K!f\��]3|�FI�3�H����N&8�ȓTd>� ��>ήA�᠀�
ܒ|�ȓ�TB2�ǎ=A��c�_�9��L��Le��D�Q��c""������ȓ!���⢇�'D��DS�A2��'^�ibFD
'`8�	���.B���ȓ)}
�"F��n�s�O��N�ȓS��ٵlʽG��BA� K��ȓJw�����>���IR�+f��ȓ#�
mZgb��|h XSn	�S�XC�ɲbE��Ku)�p��%��m]I�dC�	�K%D5j D*( r-*$�9F�2C��#i�0��mͲ�R�I"`F�'g�B�	7���2��"Z���-G�sV�B�ɻd�D��
�4,�U��C�C��j�4�� �F$;�1��C���B�I�vtf4�V`W� ��m{����c��B�	�zD�p���bn�#��"��B�IJ��4F�L�`�k��TC�	�dJ�c3�I,q�a"�GR2
��B�ɘ�%
�hS�Zr�4����sm�B�	�}�����d�,���"B�KV��B䉊]�C��Ņy�XYS� J���B�I*Ba+d΀	v�A���ƿ��B�)� j��b�ˍmn%���d���"O&	3.���u�A�=�"O60�oQc���*r��J l}ˁ"On�J�.��9���F�D(�"O�����3g�̲�N/���4"O( �'Ȟ�w� �!��.y�����"O~d""O��h�ά�ϫN�4aU"O��Iqh�	��h�'T#&��#T"OΝ������qI�A�)h6鳕"O�$�� �d����G-rcD��"O���𠋶B *Y��_3Ir��"O�5iW�?�zdz��Rn,�L��"O����ǃ>����"�	P&p0
$"ORpq"��5q��:�oG�B*x���"OLm���JB�5Z�nA/nP��B"O��@�P�l���HwmT?h��H""O�������~-~e�«\,J�>��E"OfM�"�H�2Q�]ȗ�v����"O
X�jԠ~\����$UU�*TR�"O$�Q��c�ʍ�C�R&6�.�k�"O�\b��^&�^���`�Vɳ�"O�	�ЅH�$Cj��aM�%9����"O�U�gN�ufJ$��f�0-ǮI�@"O�\*eʄ1�2\�&�3r�^,3�"OF��s��_���R�&�8G�<Q�"ODXh@i�;=��+�>�@�"O�ha�`I->740'H܃\>�Mr�"O�ܠsH�:"�\�PȀ�77��ڣ"O�I���8�-�� ����g!�d~�&��`hR$�0��$$)R!�DA�f�PSլ��l��B"�)
G!���ld&�� �Y�����@M+D!򄌂�@�a&)�im �B.U�x)!��jiru)a':v耱6�ͤ!�d�	!��lZ2
�d@l��*�!��&k8~M�G�-b&"m�W��6|!�D�:�6��I!X�9�[3Om!����M)pJ�'[L�$��ԇ?_!�DM�R"ܚ���V��ň��vi!�dޭGv�LJ��A+>�1Hn�0In!�$�c!�ܞ�F$;�̘m�!�$�( Db�+W*_��<.�2�!��hӚ�`5�H�ShRT�쒈?�!򄕫1���h����eH���kH3	f!��G�\��u�C&�s��i�v���cC!���/*�܈��L�J�-!��/�I�1�;H�Ȳ���2&!�̋E��� �	�h�ֽ�)��X!�D�z��U 5�R*x��qp%IڳA�!򄉂S�^ 
��yw<k1��XD!�䐴V��4A4I��1�uB�#7!��U�l�������v0���#�!���'~�|HRة�J�B",�!!���R�0���m�֑)a�4:�!��R�1�d�QfB�ׂ��u�#�!��6p�\�a��`Ħ$��Eɝ0�!�0#�Ty��#\�V�f��Wd��g�!��E�@�w�$I�yP��<#�!�$�5{fl�UhU�q� )E@W<�!�ݢ`��@·:��(�OXG�!�d_�<�@���$k��$3R�("�!�DFH^��:@o�(`�eq��/j{!��jƚ�;4N�/���R�D_�4!�P)� <Y��T�*�V��c��,�!��  =;�N�bQ�K�.��9b"O�����2wcͱ��Z�x�"�"Ot4��5w<y"��V_(E�&"Or��GE_�	3��xe$��QW�<�7"OL��	L2����]�\E6�:�"O���, |Ē�B2*�
T�JȳF"O@��M�0!i��� �Y�"OD�a���x"̰�'�+8z%�"O��[�s5���	Ħz�4E��"O�� ��0<��؁�V��ʈ�0"OࡧM��,�fi��ص
�R��3"Ox���/�=
����D֞.�l5��"Or@3B��D�Y#���\9�"O@��]"+�VE�U�RQ�ġ"OL�U�C01���W�S	{K�Er�"OJ9ՃѦ^P�&��b��""Oܨ�7kǖVv�V+&��U"O�X���\��xU�AJ��?�p���"OФRc�ݬ1���)��U�tш�"Ob4`W�+�2T�a���Y}�E"OR��ՆL�F"A�a��'YT��͸V.<��Kʻvy>-B�'�U��!_Ov��g�K'j�llC�'y 䐱�V��N���h[<b-��a�'k�aʣ$��=J�9W)ݹe	p���'6�I`EX��1��+�( ��'��@Bg�&iux��u��)�`Xc
�'�d�`@l��# �9��M���d٠	�'�I�VB�7K0���c�v;.y	��mi�u	q�ޡ*R#҇s� 
	�'���w�U�>�z  �m��q�L�'8X��E�W6�����~:�'\F�q����%e�H!Ɵ,t6`B�'�ؓ�bk��4�3��L���'ݎ�0W�ާi���&�C�S%
�'hJ9��⁧q��$��(�?����'&ܱ0K��H���%l߸=	�'�>�Su�ܟ@7�)yGM�`k~�	�'����H�U�����,l+�X��'���@��^��IA�@Z`����'Y\���cʥZ�$���c�H��'�P5�ի�<䡠䋔�%��'Ф�ua�A��`��O]�V\Ԩa�'���a��B����@J�|@ q��'rP�U�L 5�|�G���yW�5C�'R��s��P�Y|ZhB�aA�	e�aC�'�D�:��C; �ؠڥ�8 9��'N5��M�9z�H�	&K��m�ʓ'�ݻ��)L������ަ�ȓ�~䘑HF&��⦁]�A�>Y��zB��S�΁b��Y�)�*#�Q���>+x���f���c������ (�!�dڍ4������I��P2A@�S�!���D��2�>u�=q�.2�!�$\Ex��2N��%�>��e��E�!�D�7{�X�#��"Et��W�_�ў<��	�9E>X���oy��1H��?��'�ў�?)�ҡ]*Gl���4�^�U��1!h0D�@C�#V�"+N����]�=��b0D�Ъw �5pyɻ�hƿ��ݡt`0D�hI�� uI�xQ�"E�k�Ƀ�D2D�$�$&Һ<��1��6r�bȸF�1D�0�`O1� ��U�xx���M:D��L��Q�!k�l-a�8D�� ��P'c��B�R�s�V".�.�ZG"O�M�����W̐1�wd�<k�D��"O^�2�}�v���)皉��rG� 5��8@?>�0uŜ'D��`�ȓZ �zD�J�n�xt���B*$(�ȓx}�t�L-��$C%w�$��:�]�D,8l���\�x�d�ȓl���gD[�mN�4�Fv��ȓ`�x��%'8>N���f>�-�ȓq5b}[ /�"����K:a�ȓ-<�i��^�p���� 2gP<Նȓ3�8XSJN�+��#B͍�3M�������K��x����P ݇�u  \�4���8�������#bش�ȓ�Y��N�!wD��C��
�pX��4bP1��ц*�(�	���?U�ّ`�#Z�a�ŏ��w-�!��;�x��u��>Ԡ��tΝ� ,C�I�{��4��bC�[6�|r�,[8B<�B�I9ל|jQ`ۂ,ڦ�H�?��B�I�0�D�#�%���Ӭ�}lB�If�@���&��%b$Q(J!cD0B䉦k>��OP��ѭ˧ulBB�	�j=� p5d�4�*�6�n\@B�I�96�Pfȋ
�m0Q$��B�ɃU�8i%��&2�����o�PC�I/&@:��Z�++�!cp��b�C�ɬ�^�;��%1e��8�
ЉhϲC�I',dq@��"T^�� Q�6�C�I =db� ��ӃRL�ɪ���$�4C�ɳL��Ix�I,5���q	Ce��B�rG�YA덮D�$�Rd�)[;�B��)_ܢ3��T�X����q$�*Gd�"?��i%a�`�vI��r��2]�K?!�d��m^�[�e*3�I�p.!�D/�h���b�y��|vl_t!�d�na��5��;�,��WiL�1\!���[�[��1 �\P��C�gJ!�U�`���	��!���;3ǁ�
@!��6N%q�c�2g���C�oP+2!�dڢ1�5��G͕��=d�P�|!�d�4MƖ�"w-�N�8q�$BZ�&�!�,�\�"�[�?}�3 �;�!�DΞ$�攘���!yҘ��-֘6V!�+pH���f-�m��k�n��!�Q�l��l��m�
@^ƙ�Z�x��'�X�{��G�H�h�Y0�l	Y�'�$�
!�'o&̨���J�z��|)�'�M�ᘨ���(�*�gc���'� p���!X���E�H/`s$��	�'��(�נ=�)�PHN�+�tb�'��AWT����!g�`i�'?:�APi6cD�p��X�����'�|��s#��նQ*�
X�f�\*���+�M5�5�2%��J ��3ьաAPɅȓw�r�p�ȁv2�8c��\E��I��(�Ƚѳkx��
��~T�� d���B0m�`@YVM)G�H���Ɉc��.�b�q��)~]�D�ȓ1����2a�(@G���2l��U�2�ȓn3�Pť��1��YQ��T���������d�&2��p���8J��.��!@C�[0�hl��.Ƌc�*q��W��y��*Fg%Be�2H-(���S�? ��v���0�j[L��If*O��;f%��6�H�g�\�F.����'���`TBC2o�d���%�)'8Y��'֮(���"/6\�Xg$͑ Slly
�'�0���E���!�Q�..iF��	�'�@;&¯/��I��udz](	�'�lK���d�tt3a'�|��'��xH�m1v�*ѓ`��1H�ʼ�'E�8A�8{��łE���DQ�i��'�=yT��=doD%J
�-��'O����F�`��i�$+�G�U��'��RoK6+����2C�7b���'d�QhÆ&����2�.cB���'�d��	-HH��Bbj�[��x�',4Lȱ
��t�f�{a�S�e��'t:58�)!R<d
�d�� �Q�'� �1M�W0jԹu�����
�'��`�B �
\B�%Y3r����'Q|IKL�tE��y� �5�]�'��
dI��ia<pQdf��
�܃�'�Z�7l�xf�ۓL.K���k	�'tظ� f� ���q��Ҳ>�����'8�r�/�g�H��(��jN���	�'2(h����&2`5���f؆���'zV�s�IƋVo<��T�҅0H~Tq�'��T���'HќEQ��'�y��'K�y�@��_ d$sn�i�$h��'\�l0�G�Y~Rl�����u��'o�s�G�5�z@k%��@��'�2�[��[�H󄑀a':<e��
�'eD9R�	_�wm�
��/%� ��'�6h+�G�����H�Pіur�'�F1�!�ZH�E��A�H���'�\�Y�G�nS�<��̑997�k�'���C�,)�����F�0��`��'�X�`��9�1˔"�<�#�'��21��X�j���*�����']ĵ	�i=q�j�%�,&���J�'@v�)�I�1�h�ĉY� �ԑ{�'˪������8�l}8�N� �Y��'�2�sU�B�h?���)�?F|.Q+�'���D��
`Y�aȑ�Q7��*�'�6 kՋU�0��];rfQ�Oz4m��'g��@Ŏy d,xP�ˆC��	�'���8��y=:�D�<Hxh
�'�@Y@R�!���i'���1N�E�	�'��i"3���3E�qw��^KdL[
�'�HI���C�S1�A�fgG�S�X�'����'D�wJbt"F挱a�)��'&Хr��-d.�X�?�ڹx�'�
�Z�m	/H�ɊV�D�&�!�'��Qȥкt��;�'�?����'��!�#�؃jv�$�u�ʛe���S�'�.ĒuJ���,#�d�('�Z�1�'��u#r%!��!�Ⱥ Qz4x�'D )B�&:
�1��<��[��$B�#�\t[%���3�F��#�>u��$�<P��� #��~�<Q��CB�b�!��++�b��`!��d� �W<!@!�d� �h;��->i$��D�D�!��(ZY�r�EӢ'�Ҽ1��=R�!�xyjT[��ިc�zݨ�!�4|!��ŗ )��H��W4X��곦K
!�dB�~M�(Ӏn�R��#C� Vn!��� <��a�HP����"U�Kk!�� X��įҪugT�1Q+�;Ƒ��"Oj��3	4?��$3���0�8��d"O�u� j�~R �a�	8���"OF�!�̗�m�4��F��>�b�J"O���s�*
P����ă�A�\�"OxXF�ɷ��0��W�AȬ��"OX���RsY�!��ގ�H�3�"O�=�P�A6K�8���F^���4"OZ��D]
o�������|t!c"OP]pg("\��,���$�����"O<Q��&�_<�ǌ)H�z)�!"OL�`��i"�Ț_p�Ru"O|0I�̙���Q�ě5$@YR@"O|YE"� ��ѵ��+h��+�"O�̈��=xP
��ޛ-�N�"O޽s�G�
0����B97%z�C�"OČ�0� 6|\ڰ��	"0P"O|� 5���0�J|kd ��""O����`ʸ����tc�#O	>���"O8���!jO.U�l�Fែ1f��ȓzZ�a�-D� �d���H�b_(C�I�{�� j�3=h����N-�6C�I�<0� �+�A�p͸���)NxB�	�	���"�X[���g�M!�D�y�2)��ǘ4lmn��Ŧ�G!���F��HQ��_~���xk!�d֍��=�#_4��9�T�R!�$[�+]lhStA��#�"��ː(o�!�䒠\y��SQg�!0���S��d�!��̠>x2�HPN	@�<�˔/�Z�!��8�rh*��Ţ1˪q�S�B�4�!�dZ�:OP�p�9�U�fG�5z!�ė�o��0h��ĜR� Tha���BX!�d�-I���E%A"Vyt���~0!���I� �S4ė�aB��3,�	s�!�.6\��aػ@mZQ��Q�!�ҝWT@%b�Z�#KH䐱�7�a��O�I�-�?=��rcN�ŢdKw"Oh���oN�/jt;��8Y�~���It�OК9z�eZ�R��+�1@y�	�'ۤ	��0*{���W*K	(��5�O��=E�dl�7iv�IT�W�}��<����y��C!�������JtfH���p>��͏PM�A������)�b؟`��_�m#�;���1���T�l�ȓ��cF�	���	�ںʨMGx��O��=��8���z#i�g�eC挆0_��I��M�LX��!(��#U�`���'�4��7�GLq�(��D1n�z���'����!�52d|��Γx�Ҩ��'J��3!�6�x�;v-��y�)�S1IZ�̐uJ�\ȕD�*�B�ɰOR(��b�Bƒ�q�i��KN�"<Yϓpq�!%ӌMsbmJ6����U�ȓct�9C��6@��A5M��U1�'�$B���3�z�k�H&��9q
�'r����';��Ȳ,��&*�8I	�'����W���X��AOO�f�>8:�yR�)��V����Mל��>K��B��'���B��r��kC�M�WL�"<��{paZ!6_ȁ[���J׬1�ȓ7�P�*c��d�^9�w����@p�'���Y�8�v��5χ'W������'�XSg��^����U��q��A��� 
0IЍ��/�:\#���3�j����@���+SȘ��ˋC�3�	�9�����҇@�x����:zC>�����N2�@�Ɓ�_���CҍWCzmr i+4~��%;N;&���*L�6l�@B��X���r��9S��P��L@X�T��uX�=� ן�XYf��5 �����I��9"O���C.+mJȣ��=9� q��'�����&��>�&ɻ��EH���S�9yQ� ��nH-�1
�2�2���9J�(�P�Ѩ %���FS��[�;O�8�`��(!&����Ӱ��M�O�B�?��N6'���In	�0�FS�PR8��
EL�ALr���t�2�i!#��i�	�ጐ7Nax��7(s�F�@؞��VB�)6����ʊA�V�Rb%@N���3Tb��q�U����Za$��H(�� �8�Qw�ҏ
��)B5��J�<��GQ)w� � �E,7f8D�`� 
,�Rg�P�c^��2�B�!����Q�v��>�ݘ'7���ūf�N����<#�rC�>! ,�������^}pt���G2�S� B�k�X@��*�C�J�1D �.���Ŕ�Pc��I�/Ùq�ܹ�.�/��-�Wb1|O9��~"�o�+^��p���Y8���'�ܳ���B���ī�#O�|�����ֻЂ=B�E�*t���p#M�m�O�����,t�!+$�J�P�f-�qF[=.>��bW!?n�V�A׮�bE@m�!�]%X�B�I.P�Yid�[�m[Fٲ��G(@J~�"��E��=��.�f�R�F�S�IIT�;��g��*��!Ȉ؂������P#�D9D�TI�G�@��$(��3'B.�Q�aS�f���cf(#'��p�O:���恰2�1O�UA��z�P�M�2�,��S�'��4�.��:��y!"�C�E�굃р���񢅌�"EX&�(�*�9(�r!�[�az"SW/&4�w�i�
Q��D��'���뢤̧&�J`�/�Kބ9� �H�/K�p2�*W7��cʛ(i��zt
�0L!�F32E>Ѡ��*?�����Hމv n$3���Qrlu��?�V�8��	&W���D��3��t�-B�@1���żSB�fxTBP�]6'Z��N@5�9&�����ak� *Z��)���Xb ݷ$Rb���5�z�x��%�:H�⑓&�<|Oƥ�t���j*޹��c��a�dI��Gż}̸eQ'�0C�d�{��W6uF�w̚w!����\0B-^���B�4�"��2Θ=v��O���nr�0��ׁ��l� &˺`��E_,���r�5G��j�i1�~Q"O(�v�Y-N p}H�C�D������b2��ڄ��q[,|�/˸?i&�#&�-O!�Oa���@�!��ٰ8L�h�5ˌ�5y!�ĕ0����]�	2�,J똧vN�A���i��@���쒂���ϵ�U��yү��^u�|i� �:W }�$a<�0>�"�K$��'�H-lW�L9�ˏ�^*N�2�]�Ck�0��%˖'��`��b�� ������FPĭ��
f�R`��V�T!`�J���h���1� L ��H�A�<�h1DG�/ҘH�p�`B�d�8ə�^�&M�l wn�yÐIHv�S���QZ���s�*ةg��f�<�����;#�\�5LDk��cd�eH�\��eRX�B!EPc�� C#�,{v%�.Q�l·ebpp "����i���'�
M3�+�,:��	BS{F��a
�{D��yB)е1�ڝb��>,�4�)q���v��IQ��T �ےS�0>�������|	g�؊daV��E�'�r���R�-�{�AC,m�N��n�8��͔���� e��POP���I�<��S�Ty�pB�ƽ��M�`���*�x��M�ȟ��c$(�-���x��� R<���"O�r��&�
�8G��.&b}PF�ȱ &�I�ra�����y�3�I
2A+W,wX$E힗��B�ɭRߚ)Q��� ��Z�i!qI�B�I!7�|���(����<(�	åu�fC䉪`��lz�U+ !����0Fd>C��Yb����K_�?��k�I��C�h��Y��£J֮�����.#�B�IH(�Hz!d%s�Hp6P�R��B䉣sޔ�pΕi`!��.��6�dB�	���1�`��j.L�B%"Y<9O,B�i�BD
�B4xϒ�#T�RP0B�I8z`rr�\0�Bd+ hQ��|C�	%g��,�Ռ�|.@	Ri��U�LC�	�$E��]����4=��Pv�2D�lr"�ĔY�VYX�̢Uu�3�1D�� �%J�+.R_p�1�(D5� ���"O~�M`ْF �Ҭ��D"O$TY��
���Bf�4̾�9�"OU��H��\rQ��)�.p�"OhT����,<��ɗH����@�O��=E����	��EV� �jL��y�L]'sW�!9!lԆ��y���y'W8d,�[��J����# �y2l0%�����\@&���TM���yA�*7:���6.U�4>޹�$%[)�y�Nݧr:��e�/OZx���y�D�7#��p����LӺ�ۖi�,�ybg_�&��8v�'t���!�lH*�yB%��}�LXC�*6t�>e�⮚.�yH�N�ޕ�g���o� �
����y�ʎ�>�v��� ҿaUP�`?�y.҅����E��0H<N�Җ���y"E�^�#�I�7�ޑ�ҧ_�y2F��4!J�S�&�%k�D���xB�S6K�2�rrL �1�L����M�8a�ē<�@�U�1�^K�䖛k/̅ȓx
�@SU!�&��J�`�p-��5��ara L���V����L� ����:e��]�ƀ@	��X��<<%B�H[<x� �Y�$J�VWL�ȓY�������3������ [=�x��@Dp��<&4� y`�� Tc*���HDֵIF�Q�B]�g�?s��p�ȓw&��Z'Ȇ'o�y"%� �乄�ɍOߖ5��y�-Y.B���g�>3���iZ��y�F ���鈄Mِ0�ʀ��@��yr���?+r��UG�6z��d*ݙ�y��=x��q��g׆r_2���$��y��w��%pB햋lOb0�u�N��yr&��rrx����źc�$`@����ybI���@c��cx�Y��Fۭ�O.��җ�(���PVS(+6�!v��*�^HPG"O��p����t���(���Q����$"Oh��aBk
B�;�Փ6����"O	b,�y�Iا����9��"O*�J�$[��ȵ��$σ+݊$��"O8�;�K�-a�t��d ��Cf"O!B�K!H&�ӵŊ=��,�W"O6��ᙝa��m�1.�-j\d��"O�c0d�-3�| 6MJ7#K �QV"Oh��lAOrVAhe擢^<�隕"O����_�va ��3$�K ��A"O��j��W�=m� ��\�w4���w"O�t�%�J�EX���Հ��e<~9c"O��0��
i��e�5��63f� �"O a�) h��\▭�-Ӹ���"OR����;y5R�(�t�0�
�'~�Di�j�5Eh�
�Hτ;7�+�'��􈒥R�o�.i3�'2a�2��
�'���1KוF�4D4�M b��
�'�"��`LC�JN�� g�ęY; y�	�'a�Q�l�>�"9X2�O5Qܐx	�'j��Pp#V�J?\��!���d��604]����wx��R���g�I��d�t8�#Mɹ#n��h2)=1G��ȓ)rI3QO��!M��x4�J?��!��T�R-�SH�yr�Y����]�&(�ȓhK <Y�゜D+4�����fp��,(�<���
�2z�e���Ya���S�? �Q��n�.c:-s�iW��t9*�"Ot�I�!N��0Z�	{��3�"O �!�ݥC��H�&�L^!i�"O����@��(D�N�1(����"O���nR"e���z�Y�.L(�"O5���7 �z�*&(�<>�*5q&"O�
�z� `�S����
���"O��RE���E�;���2"OP�B#�^�.y�A���_�̸�$"O�@�U�Z&Q�Zq�%aۜ]�X@�"Od��el�#:��i؃AƩE�|�0�"O�h�b�>1eLl���W�s7؄��"O��P������
�8s(�Ik�"Oj؛�f^�r�|��ة\x,R�"O�EC"aϲ>#���&�ɘi��!"O�X1�F
 ���K��Y
�"OxLH!K�1c�ȶ��nU��"O���f�E���%�2Z�Fp��f"O��P�.G	!b��+P�� xPr)��"O�axà�~;���Ҥ�/lI�9x�"O�k���,&p��l�')3��Xu"O�l�u^=�����K�YZ��7"O����˹���hu�:H�}B!"O�����?:{P-�!�͔1@d�s"O(�OMT%+*�-2���(�M�r�<��&^+`� @��P�Pڲ����i�<	�	׍
��QQ'�>}1@���Xj�<	��C���� �9\
���`k�<I�	�T�����	g�q�/�f�<`�˄,�L�S���/R���Kv�<)A��/5)G��'/
�d��s�<9�o�4���:� ��
�, ��Tm�<a��w�j(��"�b���s��p�<9pC9��H�OH�'�jй6��n�<9юG{�>M5�B4��j��i�<�)�B����#�*����wWS�<��j!r+�s˘�"u���H�B�<I�hH����b�f�#���:4�g�<A�&k�X<#sʛ�OPU�Df�<q���'�Pm9Cn˜'M����x�<�ꏰ[���)A�C��ͱb�<��K�{V�f �J���i�Xx�<i���ʑ�M
;����+Ky�<��M̂p(� n�Rh�a�q�<�6�����1K��X܄��a	�K�<Q�[=_�}��G��O�`1�t C�<)�`Ȕ3|�Q��C�}^q�b�~�<I͋$c����E�z����x�<�1	Z���}�ek�YX����v�<q�AC�;��� �F.*r:���Oq�<1R����[f.�32D���l�W�<���ʓ��!!���{� ]*��t�<�_�^���.�b޴�A��\|�<�S���\�u��B�?Gjh����}�<)ÃC�	�x؆���
�\�A�Đa�<)�@'1�H����8cjM�ŗb�<�0��,`�]C�!�;gV�I�,�u�<AD�ˈo��9`��8h.���SEX�<A�-w��D�N�4?ĺ����_\�<)��Z.Y\V���7v���zb�@�<�V	5@�@D����8#�>�Q H�~�<1�/A�4��{%AB:%;��a�c�<�NT�ZȺ �`*��3��A�<I}bh�X�d 8���5O�4B�)� l\`�c
a|Z傍��ع!�"OR�3�f@8l�TIc�E=!/����"O�-�DI�� �"��<AZ���"Oz`��I%{q�k��(b�z�"O�tX�@#v&�s'��!��]��"OԘ
��.��c����A�"O���<����(U�fdh�%"O.h��F�<&�|��H�o\ё"OX�)��� !�R��ǧʆd��:�"O����4H�&m4�K���l�5"O���I�3WB�.�-3�4�C"O��j%�߄	\F`a��[���aC�"O�)�U��M��9�G-�
�ʤ"Ov�j���06�I�lÂ:�H��"O�-i���V��L�!L+�6px4"O����,a�ܴ�&�ώz�l�Y�"Ob���J�m�`MɷA���u"O \#4gY4�j��s��	��(H�"O��ЁkִQ�d�8���"�C�"O��s�$ұ5Qc���<����d"O꽩7�T�z�˷��6&~!Ѣ"OR�z3�Q���Z���81,��7"O���D���*B���	:�l�"O�b��*�Br��*&���r"O����ގ2��D[�:.�T|*�'8|`y�'A�jJy���GG��s�'���� ���d g Iܪ �'9������4�ZQ���-~2	3�'��1��"E��𫜫~=��K�'��U��n�!��P�G{nR�P�'A�L�d��2�nDauʞ�y�:���'�� O�$g0��d��)s�)��'�V�b�P�]�4'�"?�l��'މ���M=Ia,�x�l�&&4���'�ȑ�T.*�~u:�J	.a�'�4�yڜ^�����A�u!e"O�1��߄ ���*�HL�x��"Oh`R2/�g�T�rt�'l�*��d"O����	R�@D���-��&D1�"O��@��;@�@Y��̌k50��%"OyCB�,da��ٕ�].��"OP�����q�Ck\`�.E�v"Od�x�mH�A��a!
ʪ<��ГB"O�����e	TɚbJ��AL�As"O�R��W"� �yį]�1�Q��"O��RR��J|�T(��/2�=A�"O�a��+�z-�`��	����d"O�]���6@2�ai�E��||�"O~9����Aڄ�D�H�j��eK7"O�!����}n^$a�DK�G��W��y�c+=L���V�<�*�1�eф�y�ÍA�:�qB@��@��ͅ�y��P�7lЪ�gI���	P!EP��y�>Jh� �������M�"O^�`�%L�K�p�b�I8�((�"O��''����j�� p�iJ�"OP9 �|�d�B�H�(~�ƍ�5"O,pK��f?B�zU&� u���F"O��E�ޏ��De�f���i�"O�� vON\Sl�9;�*��3"O����E�+�Ç��+��V"O`�C @��ic@�O��6��"O����I瀠A!G&2���H1"OJ��C斡.��H�K�6mpR"O� P��4O�(��Z�E��6}n�b�"OH��@��X��= tMV�Q��`"Oǂ�$"�P��
��%��"O$�rDeƉ!��lC*�l��Q��"O��C�FR�����G\�wj�\�"OX͚�Bݖ]��Q���:XR@��"O�+BƖ�S
xIB'N;~f��KS"O�PA�V;�2@��I=.���x`"OL�yq�bB Rg���Z9)���M�<yc&M='�X`Ӭ�B�����J�<�t�V�l��\�c+u�8�б�In�<���Y%|&>�X&�I&x�2�n�<!TI��h�u,lʔ�T�*�HL��
��E90%��x�`�I~SDY�ȓHlDp˦i%����pm��IG���tӰ�s���	_BEc��ǆ}⬅�E?D�2^-R��A��+2��ȓf����ALor��s5Ό�^䘁�ȓ{�ƩBO�%�R`��c% �Ն�Q�
X�\6
��$�_P'|���XP$p��aL1m�t�eeƓoOL�ȓa{�щl�БU�Ȏ��ȓO�ra9��:s���F#������"�pF�  qF��E�yU�)�ȓ�P�p�E�0nd����"YŅȓjzP�@ˏyi� ��ɘ{��)��b����&A�+EF��1L$|��z��v
_,]�:dXg��n��9������'I�<[�ЀBU\�0<�ȓp�dR��M*Z�@������&x$Շ�6�h!Ċ�F�^PzƢP�%�y��3;�
���d� P҂��<c\�P��z��3R��ѹ���>���ȓNRH�⁫_\aa7�!iD���x �Y�b�1`"�ە�*]���ȓKmX�Q#n��@���+X��a��TtTJ���jp#S��o0�)��sJv�*RH�5Q�)��cֳ�̸���4�w�9$��Mj���=��C��1s9�U�3�J0���yS%W�.C��1vR�`�c��+PRP�h��!=!TB�-H��˵�l�m�%��EL B�ɭ *]��"b��]Ze���n�rB�4U�z|�i�����ũ�3Z�rB�	4�,ɈC;i�$(6�Ĕ��C�	�"�j����#e����eT�T�0C�ɧ0Z�U�v�ŰK�\��Se��B䉸}Zj\��oF:<~��;��ܞ!H�B�I�d�$�W'��kV������jώB�ɍ+QR��k�'׶����ܩkD"C�ɮ.�T)��Dj����!HC�	63-��DA�H�dተ��z��B�I)�v\`kH���;�
�0��B�R���K[#kP�a{�/؏\��B䉪g;�A� �#i�=�$hJ�	�'���+2rb<}[5�ۥ|��4�'7��z�)�">N�|�u̓�����
�'v�)��=2��ۧ�n!�M��yB��)c���q��r�:�y�	�:�y��
�XABl0�Z0���Q�� �y�gȝ;���["І5��L�$����y���+t񛑈���hW�G�DC�+ ���$.ȯa,�Dۅ�Cm�B�	FՐS�]���:� �6G
">ٓ �!}��;AK^(�-X$��<� fp3r$[�"�EZ���Q행�=O�#1��Ѧ#}ꄬ�7� ��@Kb��a�Y�x�H�P��.���]� �*�oڥ��5\��u��&�Mb@�/�0谞'�x�4�*�)ڧ_��Ejt�#� X�g�$
����	Z$FF�O�?�!�#2��T�1��?Wl��ٺ��'� 9G��<��D1BI��B���O2<R0��'㟒�ΐybO�P��5�`�)Rc!P��j��0�����.=wnu�Շ�5rG���G��2�~b��.>��O�>mh'މo�0�ɵ#��ĜY@E�v������i�]�ڠj��Kr�՚B�;N�?y��)���1����Q�@��P�h��$�t�L⟒���BG�>�^��RLB;�����>�Ӆ�����OdPL���9:�\d��ƨa��P�'L����퓄.BJ�'�5$ɀ�(V���H�2������N}Hdr��E�c�̘�baKdƔG��l�����C�^�V��$�5�BaZ����
9>`%�dR���Q�S�ӊ=9��:�$��ƴ1cJ�z��>A��E����'�?٤#� v��AA���'�ܘCFF?�S�N����h����D	�4t���@��S0衉�`�+O��M�?E��gU���8A�	|�<�a��� v}T㟐��O�&��OO;���rC���y��{��`��O�OF^e�DjW*6�|R$�5�@H�H�0����ا"J~"!o�D�~�kw����
�n�=�T\IL�(���{%qO��|��Tdt��`l<!!���}�I3`m>��ڦ��y򴢍�/�ZU�a�ʌ0�!�D�)B4n(k� щ-�N��A�8!�]#�z�*��ߌb�������c�!��H���g�\�@�R�f�!��ܜE�^��)� ������J�!�QK��P��� P�5G�e�!�d�'H�4�ܯ(����c�!�D���e���H�w ���OG6Z�!��E�Yzm+g���6fzɯ?_I�X�ȓK\��D#'��,)�_x3%��� 7	���r��-*�i�ȓ��I05�4S �y��'��ȓ,'��0CF�G{��+j3���ȓQ�.���jC	#�.���,m��� �UYa$��c��p�-�o]`��ȓPdԣ��U�kj�#�-	�9��Ї�z�j<�w�D�D��`�3k?o8�\�ȓ~8��� �A�.P4�{�`Ƀqf=��W�~Y�>>� �5TV��ȓg� tp���5ƶ�!���(���ȓA�`k��H�|����D�-SwB��S�ƥk� �*{^lH�C��x\�	���Dd��bȽ�бs�@ߡD�(%��bY���C)\�H#F�ەOj���c#���Ň���e(��B!x�<�S-�/C���;u��;u^�`�HAK�<��L��1]�̹�J�1۶e8��N�<��]�Rj0��BF�,�&dX��ZH�<��J�A���#&bH$#�� ���z�<�q �tm���g� }�Ы�/Ey�<a"�ΕL$�G��� �#Qw�<�wIT�N��������,�0Өw�<�F��]0�kF�+@�=� eu�<Q�
'��ac��Fl�p�aI�<ɵ a�Be�q�]����h��A�<y����F�2Պ1��l���6G�c�<�7(�c~h�$�̘x】�E]]�<�t�_X�B���`F��k@�D�<Aao�>8<	�pE�y�&���	�z�<Y�$*�eBG���9K��3�M�b�<� lx{ƫM�/:>�r��qp��"OPph�;^�I�ӑr[8 �s"O��!T-µ67�)�_�dO��"O�� N�ss}*��N2���"O��� **� ��e�P�b�"�"O@�ɗ��oh�];���8���r$"Oĝ�mgIjbT�wp��V"O2$��%����7��	6�!�"O�IRCne��Z�U�z��"O`9�ƫ�+Y���iǥ��!z}0�"OR-�"aC?C3Ԕ@e�!L]��bR"O���4� Y���%v>4�
�"O���&��U�*tw��_��9��"OԈ#��59`-��"١6'�a�c"OB��&��b�Jq�"��8�)�e"O2�s���;��h���,�d)A""O�T��M�(��l�QL^�;��=�S"O��zE��5�f���+��sעH�"O2��[���MѤ)3�d)ئ"O~����Y)o�F��2��;��Qrb*O�$�q̜�`�p�ZV���=ψ$�
�'�\h`�P�Ԑ�2�(i��	�'�R'� 1V.�b�@̚d0�AH�'�Ԥ��i�*��ucb.��^㲴��'���FA�!�̅	󋒗R�����'h�y�Ӿ#�B%k�AQ�Mx@
�'����R2<ΈR#ϓ2��13�'�j]�@&�8D{,)�V�-�A��'f�t;!l�6nB9��ǐ�M,@�'	 ,�#-ЪXt�'F������'3챔�Ї,rT���%87�p!
�'(I���+ u�t�
X�3����	�';6As%�@�� ��$'@_��
�'�msrm\<(*>�8���7>I���
�'�x�)���,�&H�t	,8��	�'H��ؑ�[����+D�
&��9�'�U��j��`�YXC&�&�b�P�'��h�d��$����@�ҨB�'�);���U�~x���S�k��'�|��h݄Rw�8��I���D1	�'�֭ $��2]������=-�}��'������$�����X;�X�
�'��ЖE��k'�=z���+����'���A��.I9$@Щ �X`9�'�2�(��*=�#
���qA
�'&��㨑 ��@�#a�ͨd�
�'
�i8dL�`�Q��@<Z�J�
�'��(�2��
�
�NCԴ�
�'m�л�*O�^��(��톌wt=�
�'XZ��	�	���r6��,j�Z�J	�'S������	~p�2vjF]k�|R	�'�d�cA�(F�"��Ul��Y�蜠�'?�]31��,�4A�T�I !����'�@��s�צ!0^���}���'�4P���}R��s`���d��'xZEF������5 {� 2�'fV��E-7���A�+	�v�
	�'���X���:���B�Y�W q	ד��'K>��⡖2Q��L:b���CX�U#	�'v|Ų�����֐�Q�V�:�xp 	�'dd��g�E%`���-ǀ5:��'��)P�++���3�D>}Ph�
�'P4��D5%�V���,�<�ȓsb"�p۱L���i��3"�����S�? B�����-5�S����y�ԡ0"O�� ��ǡeL���[B&֙	A"ON��WD��BIr��F?���R�"O����E^!����"�����"O��9�-��LOP�;�*�l����F"O05�h�pV�䇏�ɥ"O���
7h��P��+��}��"O��Z\+�QsÅ9�|a�"O�����}2�B���dA{"O��gԤ\��1�u�_�?�$��"O���E���rk�H�G��s)�@0�"O���BB�� �jWh�
Z��Q'"Oȉ�񯍧<��h�,<���9u"O�
�͠kQ:��q)�;C�ʡ�"O(8;�M݊�H�gŧ)�TS�"Ot�����E�|��-�iC"O���`��m�E䅞)%L�%�"O���sH�%-�f���6-/��"ON��@�ш=|�@���~lI�"O� �A-JόȘ�e��p��X��"O�t�'�8P�v��WE�7i���	�ȓG�<�3e�F�5Q�JR���}��S����V�~А�h[�X������I�W�|9���ł6�F���D��ً2@(}�ba!�]����xv����*� Y��a[0l d��t̶��J"����u�6	s��ȓp;^P�%�0!���.oX��ȓG��!�D�?z�EJ�J�+H(�ه�Q���!��Vih��!Q��&��]��
K�y�e��0�f�c҄.lf܆ȓR�\��b�:�ʥ��OÀo�"O�I	��02n!#����{%"O�H��ˬ3�8�14!i���"O<�	���X�F�C��6�a�"O^���_;ci �P�D'J���Q�"O a�I�J��<C񍀙�J��"O�<���@�>阜RCo�-R�b�1�"O,���((8t�P'
�&��"O`2VdZ�>���uϝ�ݞ�d"Oh���R�La�q�4@��@lf��"O�tk$��u0����ٍ+W�;3"O�����+L�	�#�zK�x��"O���W��c���[g�"of���"O�����8�:ȳ¢�2_�cW"O���`�}�PqW蔯!��Y�F"O�-��f��v)���O�S�fih"Oꔊ�EP/n�m�H� �֌@a"O���%ϋ*a�����oB�q"O��BW����K�@:#4�E��"O�`s�L�����$��%�P&"OT�*7�ï0�Z�2͎t��s�"O ��L�-��p�i A�>�"O0�r�#%]�2��F�.N�A"O4�%LY�MqJz����w"���"O� �#���4���&b4y"O��R��>Ur��6���xi�"OKG�tڦ0�r��`���&GW�y�e�<Ϥ�H����	�@��/���y���_�����'|���4$N!�y"�K�XgŦ%������y�‮Cl���dG�9��@�<�yչ%�z�� �c$�@�FM��y"�ܐ�5�j�7Xՠ�2���y
� Ҝ�%U	&��R��7���u"O|��G�ZDh�MR�J��"Oj�`����\�M_%.�RiX4"O�Q�v�	�hЦx ��x{,k�"O<������)\��z�"O2a�FOq��0FK!aI�P"O2���DޯT�.���E�nI�|�%"Op4z�Գo=�(��ܧy�\͹�"O���Vi׵`�z�Żg���u"O���5�G�Y����V�����c"O~�K���M�B�q���!A����"O�0u�ϕ1Y�M QL�4��"O���!�Q<�*paq�S�4�u"OT��3�ܥ��.�j!j���"O�}	6�	G���؍>XQ�"O��2�nS3J d0E慖m \�C�"O:)`D*э7��yAe�&duc"O�4l^�Z�RI�v�EFnYb6"O��q���?�xԑ�����1�"O\%��c=��u��-�4�X�A�"O�� �_0w+���Z��U�R"OL��e@�Z[�i�u�n���"OX�&�4H�)J�͕�c�B@�"O�d 5(ޤ�B���#Zr����"O�����*c$(���_!"]����"OZH87��zy��AFk�82��Z�"OL�Z�wÜp�0�Zds��z�"O� Hd��f�~�P�*�/`ڕ;�"O�Q�cM�dr�Ă��*J.��&"O\M�2 
  ��   �  �  �!  c,  �6  �@  �L  dX  �c  �n  y  �  \�  ~�  
�  *�  ܰ  �  d�  ��  ��  g�  ��  ��  @�  ��  ��  �  L�  � �  X � �! C( B/ 6 i< PC �I =P LY Da �g �o ^w  S� �� ڑ e�  `� u�	����ZvIC�'ln\�0�Jz+��D�/g�2T����OĴ��F���?YV̒'�?��]O+����I�2@Ȥ�ܛ*U`Y����X�Bc$=�[�&��u��1{��I�0`���)��0~�d�`��떩��L-ڜ�W�˨!�0�z3�J%�T(ѫ�(�I���0��'0�l=M�ڌ���˘1���Ї��L6�y��m[�>��D �2��D81"H�lZN�H���ǟD�Iğ�Ɉ��TB5"H3I�t�C+�u�\���+�|�s#�:�M����?!�'S�@���?��TTzX�5O�!l!@X6!��R�����?a&�i��'kV	K��'7��{_w؅"4'庻�͟�:�P��ۂ ��:���3[�-�'��^�=Ey�ݑ
���(�� �����nّw�R�s�R��̓���~��;R7�CBo��|�V��,b�B@"QC�)$��Y�J�����韴��֟������	b�T2����-U r]��y�
L�.G(3��'�@7���-z۴3�I��M��ƣ9K��-L&S��);�,�#m14�a��#8Xx1;0j����-X��F�|���̣�~�'�5��~�0j�.Apa��@�](��� K:&�}�B��:�������D�ش+]���O
�I����]�Lخ\�"�i�$��G"��K^�`lڽ,^��j��\ H���Ƌ�b���PJ�J(,��ݴL��c����U9b@����A�B�*g�Ӑ$�H ��(i�%lZ��M��i��z�-T5s�m�8{�8�F���1�N�6��C1i[6m��!�gŎc��Th��h�ho���Msr�2\w�ya�B�m�ji����?q֙2�+Kڠ5�2�_.m�Aq �i�z]�bI� �Fš%��."�Y��'��O\��PNT6`��0A"�V��L���OD�P��П@�Ư���Mɟ@�� �2�;!Q/Խ��'��I��8�	�|�#�M�;�ιy�I̚EC�}*۴XڄxZ�BI�L�(p�G\}t�{�78���Gc�/�R|q�8�?Qb��j��QZ`ϽH��!�Ĭ__�D3�o�O~�by2���hssV���v��95f��?����?)���'�2�'t�[�3����?3�]��B͈*\�2jxӞ9P��7;H�$&��7n���JCOǦ	�'?`1Iw���ľ<q)����-��|�*7aT^�+�'ܧ/���D�O�9Z�iӶ8��'��k\���۴��O���-�C��..ä�����py�`J5j:ƙ D鍢$��G���H�+�}���֎H�6���Hѭ������q�ZLE��4��!i���k�V�� nU
���2��|��'��'F?Ȇ��l�ԔQTMO	p�`�D&�����hi��b>a�3ђa���6��Z�BdnZ�D�'��*��O��'�Q�${@�#c�xv�AT����0�͐4�t8����M�o.�Mk�R>x�����R� ��ȥ%������2��M���jCD��a�ʽVe�@���$�F!��dŵ[4,��2R�nh	�ůI�P6�T`y"#K��?������|B�V.)�E�n�O�|�&��,�'��֟��B�O���,��FUYmMx/FLI�Z�<�ܴE���'ɦ6m�|��'��>�^$�%m��z�!�n?H�blb}��'{�Y�ؗO�IW�Y_����"QJ3����"V4;Q�H�a@��'�$���Ōrj�<"N��HQ"��C��>�s3��>0��(-&���b�]9p� �3��U	�+c~6���>#��^Φ�a��,�I>8
�"P��tH���c&T�Ygr(�	�H��k�X�afO+O�$;H�=�����-��֦i��4��d���dmƟ��~��#��H�j*��av$܉y�H��xy��'&27��\RNW�E
R���P;?�@�4���4L����؇
j�ű���DMaxB�2����h m$�!@;w���mL%6����!C�^N@�aӶ��GyB����?aӱi=`6��O����V٘��W�sA>M�4b�<!������)0?�
�Ly(��)Y���C �M�� ��4�"$"��ĕt�L�4�Ԓ6I*0P��i#�1
�Ԩ	҃��츖'��D'i�L��8W��<+1+Z�e�Xy��7��0!���?V�ԷdlR�; -pℵ����7TOX�>�TN�s�%K�a�) o:I�@Nw~b��gd��Ae�Z�99Z��
�gK�7�I�r�C,��V��"Z���đ����0S�q~�a�#�?AS�iF��Zc>)k�T�qA�ѥ�p-�#	+���O�O��D�O^˓F"*�h� ��u ����i�I�̝*�����?9�4�?y3�i����0)8h���:��XCT@�v��7-�OH�d�O6�P�� lJ���O��d�O0�]�cG����A �p�q$�_	f���u�Q(s|mZ�A*�)�a�\��'jh�4K�BԀ lºysT���&zҼ�(�)
6�"$�7E�;ΘO��$R�O\	�U��_j,���O��}���v�0�'~� ��Ƙ�?����?�ef���0F�K0N����A%���hOq�����^�a��遻&"�d��V��۴	I�v�|b�O��DV��k���l˳��6���~�B�4�?����?�+O��'��$�B�ay���ص5��A��	�-��6.�!'腺gB�!^�����:fd�k#�;_v�p3p�\8X$2P�v�+�-�!?:�!��DOm����5p�`I�	F�"T33!J�Yz�d�֦�#��D<�J!��!��ɭST�yc��g'����[�IƟ��	^�'|N�I�$��8q�( ǭ$�-��'�x6M�O��nZ�M#,��z2��즁���<I���a&��B�T�K�"����D�'�"�'��)ғ%��[�o����X��u�� P���@Ak�4lP�ǰC�<m�s�'X �z����b]b�&OF�tK6M�щ�~����
�iT�tj%�Ք7�Н0��D/q���j�꥔'��H��r�pe�޲N���9K>���7�ɼr�y��3tL���ӳ]t������0G�Vzu� U�@5`͈Ͳ.̬�Mc,O^|[�.����IEyB]>��	o��Y��Z���4�v��w� ��ǟ��3(��\��](s�'R�i'���F5�^���c�d *N=�U��jQ^~��E�c� ӗϑ��ưJ���>@�P؎��a�F�&y�4�����0�ӡו���N�9.B�'�>��I"*Lљ��-vNq�ul׍N��d�ȓ_��E�ff-���><EE��+ڧ�%��.AW�0�s7�� dw>]�	��'K�v�'�'��U�  FC�.9Q�k��/,�\Y�EQ�|��Ó ��tR���\̸�|z0$�"3�Iu-`�d�Z��-{�,W
p�PV�M�w#�,�5��?�H�'�#��&0��q��O\�q��]�v�÷N�g�|Iۖ�'��I�Ξ�d�OT�=I�"�/Z���8S��0m�Fe�e!֟�yB+B�}�Z��I͵]��{�(����dAY�����'�剷k>MI˒ PZ�C2,ġ_	@PXF��d_����$�	��\AYwJ��'��	ӍG8]؆�S�RR�*��	�2�kUJݞ}��agcE�h��� �>��\!�ף�.�*��"앆��3a���LQJU�˰���IfZ ��O<I)E��%��h⋹mS�8rH/G��'Qb��(§���� ��5��%��,G&�P4��:Ȯ�1h���R�R��`�D��F��M���򄜡��m%?�5fK�b�deb�%Ļ<gj4�V��O���?����?Ѣ�Ԭn�@��(ˌ-zh��r�؅�x�`�U�!�1�S�N�(-�y(��i`^;���:H�b7a
�>�4�QeB	u�`��
��1	�ʘDl{�d��ط�I|k���O�:ÜPP"��V���
l�v²$$����J����ԉ�����!��a��RGo �O��I�'�&P�F#�Xv5Ic�K=���<��`�E��&�'SB]>1�������`��,�H�a+�n)�qeAߟH�Ʉ,r����9,w�p�V�ʧ���-h%&�dk$>��u�A��t��ɸ���3���Ũ��鍆m�� ���C/ A`I�Q�������O|�}R�'���N��^A�@qb�r�JȂ
�'��	�U.�OBPY���T� q���F�O�JĢb@��	���I��� 9�h�iU�U�QiC�?�Iן$�IUyR�ڂ@�R��ߴl�ְy�	#u�`�h�F�2&�j��J�-]�4"��iǀ-)B�S�'*�a�hʘy|�@��¿o�����V�d�LT�$a�|(,6��֘O~�,��LB?	�&*w�n�HD��\
�b&h���@�'�����?э�O�r��ď�$� T;���J�C䉗U�<3A��&y� 3�l��x:�qd�����(�'�� i���0ճ�+ʗD��� %�|m��x��'���'B��O���'��)ղF T�d�èG��*��=#خ!���[	��U�R�Za:�-�k�'rS��;B��X���بD����PaE<�Z�o�6�J�"6,�{�1�&�s�'m�=c��J24����fV�nu{P�ڍ�?���hO`#<��e<�i�e��� ���˷��~�<��D�j��8h$��D���j��x���M����V(����O��IōnH���A+IRzf�Ȣ6o�M�	֟��� �ڟl���|���I�Y`�6���~Y b%U�N���&lX�3�q�ύ�i�������X�Z�<	',1�F�@��Ǵ\�i�jU�zǨ1�^�'Pf�P��>���Ӕ��2<�<a�ޟ�	k~�� ���y����2 ��!&J̺���0>����Y���j��Q�*��zAK�A���3�I"���c� |xFu�
1)ː��	jy�o�94E�6M�OD��|B%T1�?I'� =_�\˳H��6>A� ���?a��4��܂�%<:�qb2"M'8*�6�'|�mxR�I?�C��G�i����'.��Su��y�.M��)�:(�>A�a$˻J�JCpi��#	"�,"?�������H�O�>IEНx�fC�s�G��i!����yp�Ü(x�\�3�Ѽ�џ�Ȉ�I˒	���QJN�L�RA�#CU8312�'���'pZ�+�E���'��'3��+�^r�G^�d�Rq���2(1"˙�*UB�R7�b�[q�)�,а8*�'d��q��_�S9�l�F�B(Rzx�"�[�u/&�I�E��l�(T����O��Tkvg�_?qЭZ�D�L���,����Eo�ğ��'!f]K���?1���H�߲i�D%X��bQ҃M��]��C�ɭo@��À���`�o
1Y��˓|Y����,�'_�QLU6IO0��	}n cV�u�����'Cr�'��ON2�'G���O��i�&��MSn�B�E��MF�!x�-}=��fÊ�@3:���6GT� 8�Y@+�'��{��*'| ���l^�ێ��'�$3Рr�������bߑ]JI[�+�pQ`�[�H.dl��O��=Y���W�o �X�ϓ
(F�z2@�G�!�DN)����pQ+P�bɨ�H�y��'&�6�Oz�Z��Q+�T?���;*vt�2DJLa@nT+CU�e��럐AbU��I�|��T�#O�ql�s9p]�aǚ���@+�,�$EO�H��B�)am�Y��iY鲯\�.=v1�2lT @��ȚAʜ#K�p�r�.!�<!��Wax�ސ�?i����On�PC�kEl���A��%P��'�a|� �򤢢� �|9�Dn���?!��'�Hu+�Źu���ʏ5GE� �����H�d�oZ���	t����"�R�Ŏc��J��I�;���gQ4^�B�'�ـ��o�ţG��W
�� Ě;�j`���?�0րŞ���z�O\!fUzt,:?A,��`�ݼW�hQEF��$ ��4�'$�`p3��u�@�Э��8���'�N%���ɧ��������:w�� 6���"O�%�U����b֓6)��� ����h��̉�EJ$u%��	CHU(#B,��'[��'�rbL�8�a��'5B�'7�7��!��`Q�S�
Y[��bu@@K�k�jԅqK�5��m��ቯ�1�1OlXv"O�D�X"���D�m�%ʉAB0t Wˌ%Q޼}�w+\=H�1�1O���.�	aFB�$@��
�f���'��I�V8�D�Oң=Q7�?A�u,P-'��|�t�I9�y���d$<ї#�(�Иq ̣��q�����'��	��4q�%�Y� r��d�++�F��HT69݆u���4����t�]w���'��)8k���w��I�(� JJ�r4@7�"aD,��I�i؞�+g+̫*N����BL��I5�� @����F(i�~�(ۓc8�LHR&X�j�p��(�X*<�8C�[Ο�	J�'.�����$C���f�6m �pS4F$D�����!N8P.��5�@D��
/��Eڦ���Myr)؟s/�꧜?	%ݎT F���� ����jI6�?��[�l���?�OP���&��>?�R�	P�ǫ?=Vc�!B�Lñ�M���%��+'Z*"?�r�TR�	vo�E(���AG^;B�Z���h�O{�m#D��b�Z�Z���4E���d�O>�4r΀x5*C�$�8a�Ě�OA�y&�p��ɒ1�N�k�� ��} �i��9Q"�������2V�ʵ[��'s�T�A��O�˓}�d�H����'���Ol��Ê��X�AǄS�;��*G��OH��G�C8����H�b�Fq�PLڟ"|� g	�/@��X0��r�*<�<�-,�u��K*����A� �h���k�7'����U�(iiU���%_u��'7�>̓R�m��*Z;V����1�B@���ȓCNpZAW �m�"ny�����h��0+��,S�،���R8s�Ĺ;�'�R�'n�M��vdZ�B��'���'�6��h�ևk�.��Fҡ=�@�(Ab��Yڶ��F_�d
\�{ �Y�K1���Otx���_���y�a+4��Mp���/;�"�A�� ���m�`�1��7���>���	�/p6����G�
�$�BƙL\"��T���O���.�8���[Sl�%s�V���!��/D��PB�#-���kA���5оe�w�<��i>���qy��ɇVz�Y��_�66>A;uO
d� M��&O���'�R�'Tx����	�|:�k�e�4�  ��?�����.Fiv|��F��!y��
|X�/�d	���*`�]��D+z��+5��<8֩X�x�a�����@�h���̭~[ v�v��Dn�~�<Y�FϚe��pӆ%�3;^�!c���d�I��MKN>����F�'���/'�Ȇ�;1!j))�ضr�'4� z��'��'&��5��'C��iE-�-8���Z�E�9��,X��9g*�<K]ax��ԦU�dm��D�c��q�'=`�)BIsQc�(�w`a�T�~�D�\�}�2�CgvQSA	ԤsdƱ��Ӝf2�i'��G�HF3�~b] N�0`� ��l$�l�"�$��?���'G,q醯�)h
��#��&�<iJ��\�e͓
t�y��i��'��S�4�.��	�JX���_x	{���%���ҟXz��*$)i����'+��|*ɟ���#LWJ�V� �	XC>Pb�����`'�(%�X��Q.�ȟzQ��S�������*�pZ�����O0�d:ڧ�y�Aҵ�!��WŦ�
0F_��y�mB%s.!C �Y2�B4����O�1F���&_9��`�&
�&�bx��B��?����?Y��*��"�FC��?����?)��y�.�;,.�"Ta�J�002H8M�҉�1�ިdt*�A��� ����a#����`iKAX��sP\0=���2�M�V��L��9=h���i� =��꧀  Ȑe`���L �-�9��#0�'4���s`�$�O �=1 k��ta,��PA�c���)!�ͺ�y�oC/��`ȷ�^;Y2��
dO���� q���4�'��=\�
 ����U��UK�>A��P;0$��`�������	����\���|�¢�rl�yJ��٨<Z�T�C��4��qX$�Y�';	����z��0p�ɶ��m��F�ΐ���a#�-x4B΂
��/ ~����Ww#8�	��M��(O�Xk�m·I"��wک9��Y3[b�'Lў(Ex� P�V1Ѻ׮J�)nnh�ցM��y�hن~w��c2��T��h3�/��+[���'��	#bh�P��4�?q�k�Ш��D�r� 4H�.�S &�r��?��f �?i������	^h�)�(T�`i�`�LC��sc�#e1>��3))B�����I*/��)3�	`݊��O�H`'//�-���U1.1J��'>pyQ�$�'����C܃Q�h�D�ɨ�XA�',d(Y��m��$�H}0��9���o��|�p�cK"@�Ҡ��ԓ��#�"q⦻i�r�'@�4ū4��=J1N\)���7�5C��ޫ~����͟8۳�)Sr=3"��0{^���s��Z>�FmԦ=V��B�K�e�4H��o~�R#LL`�֯y�z=G��%̅v^��uL�9dk�8��*A�����s�R�u�jQ%>q�|*��M�0}��p%��j~�-P�e�fyB�'�|���-o�B��V��M�R��ghʡ<PJ"<1�ONao柬&��
 �@ e�X��&d��i���!�+�M��?�����C����?���?���ywkL�M�b�QR蚇
g������,ц�sg���l��E�$G�<鳉�t��$}��Q�*
4Y"&lҢA%聡�O�;?��Q����8T�f3GS5�����N�'��� o��x�RM"`D�˷żh{�l�O��l&���Iɟ�E{��ń&%�x��9�ۢIw!�H>?j^d��K�-8p�'�0j��HO�I�O`� �����d�HN���f�Br)�BO��l������?����?�ƴ� ���O$�ө�d1�Ι�I��R�`�B��P�$�{�B�U�M6S`����,J��A)f%L;��Ͳ�%��?0��RL�Tvl���41���ၴN��">١�΃ᅟ�&���F�Sh����ZΟ�����l�?���)Z�L�@�P���<�QFD!��[��;�92�D�Q��B���'f�6��O�R�4� �U?�ɁZ��IO��ȝ��
p�!�	���,�ڟ��	�|
���V������/���6l@�4k����Y�E�(����r4�+��\:_���S�88e�p�!JM�;vd!���+,��&��\����r�*��/��������'����tcɅ:=�p���1u��2I>����0=rlܗ;�Pyg��D{��A��H��hO�ӷ�?!ԉ�x�|Tc�bY�U��9�5m�ޟ��'���w���D�O��'Y-z9���6��I�U�7�"��6��/.�@h���?�/�&}�@lÑ���H���4Ta�맮�i�$p5�� ��L5��!0��VW�	�?�*L* ��#�(d��GiӔ�![wA^PK?C4���a;&�kɀ�Xxx����#?	�$�ҟ�@ڴ
��O��O󉉱N�����$+ޤ!�Ԣ���'���'%�	���S$p+����J7��]i����O��'�1��<��H5lԙǌ[�Zu<	�5�h�z���O��F�C��
G�O~���O@��nލa�@�a|\ 0��^���#�]�(��9������V�e�i9���������� 	��Iܡ��I���N�HV����F�F��+��I+��H�Y���Q���#X�
�"��H�wg�OP���O$⟨�+�r�|9Z���3:0iK����x���4�����3�;u�Pٖ'ܦ#=�'�?�-OZ��M�8�KÀ8P�����l����R�-�O����O��Dֺ���?!�O]�t+Dʞ�n��9��ʝO�����d�4���y�p\y�FO"{cџl�G���x���"Э\��)y��Z��9{����[t��FS�.��F���c�9��A�3w��P�ٔe̒8����?����'�>mx�gB�	�2���L�(��P.4D���M�XpD)��'�D� f%��\��	LyүW!a�@�'�?)r�L���B\�m��Z�B?�?Y��+�a���?��O�H%��J�\�HKd O7"X*dуbՍȚ1HFC[)e$X�aW�E"mDџlr��[�J	a�b�0 ���6��U�Ujs��?����Woۊ<�ȹE"�͕�?�������6h�H"v�	%�=�A+R=.��'02�'z�AĭP�-q��� 	S�N�	�g��dQ�R�d�(��V&�p��E���?�/O���a�VŦ�����H�O����7�'�b�jďS%�X���D?2�|�c��'�R�F�t��D"��7<`�ak�l�	$T���	�%��W�1�.�s��(+����'1��$ ʻf0re��
�|�����I�	|n]zW<{����ɻy����O��}����� �}+���
�VxQ�Ud��	�&"Ort�J�MV4[�N u�l��	�h��!�W��*%7�,sq�Ôgfՙr�y�����O��d!O�)���O����O��d~މ @��%�JX���$��ZTg��2H����H:>�}9���-r�c>�$��bb��5� �HC(�U���C�G��buP�� ��<!���2:b>�$�\��h]`H�17J�	ra\�bP-�q�IpaP�$!�3��sj> *򀍑[e�D؁fQ�Jb
�'�e�t/�Tvpkr&��?_s)O��Fz�OL�'(�9�"��-.�����Q�i���9zJ�2�'���'b�fݽ�I��pϧ~����pF˦tcn@k0.��w�$�+��ǮP��"��-\O���� D(� m�E��2!ź3�d B�+9��Q�ד�؁�d)y]��#�F
�n��@h���0��4 ����A�' x���?���dD&Q{ԙ���_�<�>��1b��yR����yn��&���޴�?�.O.a���W����O��*��C2�Ȃ�ߦ��
Ós��GxBi[����#�*�� N��0<iG�D�'t�l���N#_�4IA�]�9�:��Óus��	A̓J�D3�c)B���g
"dA�(�ȓd�v��É�+,*V�	b�YQ���I�?��BmX�k�N���`x�I_q�	�[� �� ������2<�6�	8v��a�����$
�OZ�dN�!����#[�
���o��"|:��:JҠ�DOMUL���t~�ȅ"�v�t&D=[��+�B�\��F���$�͊e�_��I )�D�O�}��'(��أ���[�d�ю�p���'����#��C#r�s`��9-^dy���q�O��;ć��G:Ŋ׌їZHnE`�<�V�x(O��Pq��O.���O"�D�<9�B�U�����J�%��̢��0*K��p&MN�r.��>g$�ۉ��y�ڡ/JPē��5-{��X�t*�=ӱ�&g"��/3sT�2���yB�Z�n�Tl[@���4�fA���?y�O���'i��I�)���y��ZHaie�%|��ȓZ1T�`�kֆ;Y���3�@�@W��C���?��'4�<�QE	eW�t��N%`� �ǅ7@��	22��L��O�zP�,��"��sR���D�j	�����D-̽���(�,��O��PP7d�؟��	ҟ�vG�C/�5��ꔇ������|"JY8%x�����Y�t�0F�h�'���r�$	'4��� m۴ �	��2I��E:r��
��9�S@���l��\�HFb�'D1�>�`�M�}p
����4 �٢_���	^��AR� 1c'�G�9]P5�7�>�O�Ȕ'�������)"� ����2_���2*O21���F����	՟ȔO48(3&�'GCT�#3�ёf����k8+ _'LĭhG)��u��0����O��~̧M��J�	�=�nl�e.�^w��-��a���i�r%㶁�
��D���n�u3T�"�Cϲ��!��1Oh5Q'�'B�����Dc��s*ߒYqH���HZ?�0��"D������ ���pCY X�D��*ړU��?5���0gĝ	��ʨ���\���ܟp�L�8j��I���	㟌��ԓ�燞-T���$$	"mbЩK��P0��ˤ #Z��!=5�*��O-�O�����;�2y� �\0h�4)(1G�}W^�sӮT2��󔌟�6��S�mK�
>}\&6�d)Q�^+���O���D�),���'Bў���Pb$ I	p�Z�P@�([E�1�ȓ#�)���%ʥ��á�r��I-�HO�I�O�˓u��$�R@���Ҁ{�A� :q�M�I��?)��?���������T��Iˬ[�
� ���(=�@𐃁�F|U�D
\$"Ӄ�J8X���ɯF���G�ѥ_Bdx�F�+�$��s'ɡ=V����ٶ������	z�� �I�`���0�Pb�z��4�D�D�k��7ړ݈Olĸ�-��J�N�
DŞH���"OxU��������C!)HxQV���۴�?�)O0�D�O\��LT�Հ��0�qS��=����)OJ���O4���$ẉQ�J	(-��0�κsG��BB�z��1n�:nt˵/�wPV<�T��z��L@�#~W���&��ޕ袦�9��ɤ��^��@��{�4�chED�'�PD���?щ�a�9�䥘qb��v7ة@�hE���&�Ox [3��F�X+�.�>s���	��'(�9�^��C�&\Tu���ŝ@����'ZLԋ��'v�S��Of��'�.<��8$��Y[L�������'�5�A��U�ȼ�B��2(C�<�af]!$�D�*��Ā�6QR9�v�]�*2RR���<��۩\鞩ɢ �^��� ]�6R���.0�S?+�,�Y%�_2�dJ��˄4�>�	T����O��S�W~
� >E`��Tg����̽0O���F"Ol�)�J�i)эԬJ?�����ɤ�ȟZ�k�WjƸ�ʴ(� P���OL�Z�p���?9��?)O�	{)�k��{h�����:h`���{��bK�	 �l�� �����I/]�Љ��Łh~$y@�*!J���A#�ğ\�`_�\����1Fx�%+$Hq2V(�f��+�f^"��D�*<�r�'#ў��Y�H�ѤK��bAdX�`�t��ɄȓSJ�5+��*�~#!��63uF����HO���O��TLh����@��O�V��j�g��?1���?i�����:�D��%K�h�	@��,"Nx��CR�:}����"�<Q��I	vpk@޴j���YWJA.��:�җA�ԪW�A�C��؄�	A����#(�1Т� +��-��D��%O$��$���O`�z�(đB�Ze��FqvR�v"O���5D<gf�X�biU25n���!Z�djܴ�?�+O<����u�	ן�ΧG���i6�.zU�1�I�\1���������។��+d�n�@@jH7Iu�̥hjXB���?��UB���(�T�̠iN���@�3�ג�#�S ��%���́c��Xw�
\Ҥ*���@�+�+��E��>�(O����'~>���eH�K#�XH�o�:w�)��.D��bΔ��n�7���"�0�OHu�'�V�0W.B-zE�`V�%����+O�D�O�O��R~"-D�2�h��B_<k�D!��D�0<���[��Y���UK��m�f!!N�O&6m9�D����'�dZF�G0|?�(�J�2ȅ9��i����B�DA�0R�'��t�'?��I�Lg�Q��a�=yZp@4�+B����,k�B�DJ���I�<�r!�xnzݱ�ȟk��?>\�`� �TJ�=��/L( �����?Q����yb�����O��	�O2���U$��u3�h$�� ��υ\���O�փ�O��'�z�s��N�i?ɑN��"u���	�B� E���?� �����IU���@�D�O����O��h��Ag�VlX�I��y�j]8QK��1Ƌ�O���܅Xr��a�x֩�?7��Ь;,�!($c
 �8�i�ւn��<�`�����0B>��'�?i���b��ˢ_�p�K	�y��کup��љ'���!��?���r��m� xԅ
�?�l�/~8�Ёϛ�<A���1\�.��㟸͓O"���	ԟ<� a+����?�6aT�7��Y��V�]T��� �HnY���ΓH�(�I���쟸ϓN��'X�R9�a`R��D:'J,I�dԉ۴n22�����?!lZ!�2/O��H�,:�,��
ȏ8��I����=��B�	2Nq�� �e�!iٺ1HF� �6�O��d�Or���O����<I��?��pR�ũ�HQ�*�KTB�>:H �'Yr�'�RQ���O��G
��A�)>�(��=�R��� �81��J�Nɦ)ۄ��9y��>���p<q��S�z�HyvZ0:�H-�.HD�<��$L"E�8�qR�	� �Hc ()T�p�f��uCl���k:�i��M=D�pp�N><�xu���I��Qu� D����T�P�0q�b*�9L*��i# D�4�A��9HBj)Y�O?F>!C��>D��P���- _�$X�&�g�FI�b�)D�����'1ąR��9v�p��%D��0�I��$´mӂ��RPPՁ'l!��?���?!��?�� ��I(X���D�Z��h!Lf���'���'R�'��'�B�'�bE��EZ�F�9X(��p��Ԧ#
6-�O����OJ���O|�d�O��D�O@�D�It@��"�
j���#b�Z�h���oZßh�I����I�p�IğD�	ȟ0��%�����c�NЮ]o�"�4�?���?A��?���?���?���o����f����d�e��F�n�u�i�b�'N2�'���'9��'���'�L��PA�V�h!a�7�0q�Q�yӌ��OL���ON���Or��OX�D�O&���B� q;&�(W&L��A㦥���\��ß\�	��t��ܟ��IʟDCR��	a�08�#��u�|= T
�M[��?����?����?)���?Y��?I �O��= �L�p�L��`h̻
o�F�'�b�']r�'P�'���'G��߬9#���g˃"sרq˱�Ή<v~6�Op�$�Oj���O����O�$�O���X�zQ*1xT��	���: f.C?8�l�矨�Iޟx����I����I��	!>vٲ��K4R4t�d��M-� �ݴ�?���?����?���?9��?���c��C@'��H'
<�A
����p�i��I��'u?IX��^�_c��Pd,R%uۈ���i�ɦK3�,��e�'=�f9O��pʏ8 y��&P5,Z����O�6�m����wv8T��4�~�&_#��HpEU4� ���,ʢ�?��V�+QX1`�kT��hO�	p�D"�҉ellã�����@�A�O(˓��P�f��'�� nhJb��5f�N�)�Ŗ'k&����IyR�'���4OL����)���� a���'��9f��'8�z3NS���T)�O���MRz�])�y"'k�.�9����(�S����Ġ<Y���h�����	`.�(�JF�a؂@؅m�BEd��Y)Ó���ٴ����T���'�p�قiP��9 �ȣ=���O�7��O���7�n��/�H8$�H�R�]:�q�f-ԃW�� �W�p] �=	����$)��*�L�I @"V,9A��+d˓>4��a���'I�aW¶���Â4�l蘴��[yB�'
�62O�"}� Hz^*8#D
PK4D���L����ńC~2�߳x�b�"��&�0�'����� �>2R�8fi͞t��蓓�'��6͝�GvZ���70�1�ߗ\�C�o��9�j�Dצ��?��V��޴	��v��OV���a;�tD1�"�3��QDǓ�:k4���'}�A�B�P��7����?��;$-���# �8!`�mB3IE�]�Ԇ�fѪ�D�E(�����ù$���I�[r �6�!R��� !њ���	1�LղA��aK�>J}���	���tQ�/N5�Tx�"֐Ц@I��IS�!Cd�(��UbM�c8��Bb�F	Cݐ�"1H�F	�4����':�D����&�|��aJ�w5���C R��Lr�
��E<����MN�"��Ra�-4�8�8�T?�����25!�"B��Y��5�HZ�r|3�d�;���y����$BR�-Ħ� U�l�bU�A�L��4ɶNV��� �DĊW&�e �]�B%�@��@O8� ]XU�U�ѢS�p� i5ƄK��`��X�9E¡ �l��Y'&�@!�(uL�F���:w�L�i�i�@ԂHӨ���)��i��HQ$�\l]h�I�R�t���E,7�!`�ط�d��f N
pKF�
�d���O~�rn�<����?�����-Da�V쒼0�0�1 �*�8c-O���B�<���O��d�OB�u�a���D�2�0g	��^���J���d�O���O��O���O����	*[�\tyv,]�S�qU���q����<I���?����	x*|�����sa���̴�r�|c���Oh���O\�Oj���O&]��b�O���@jY0Z5V�˄�H�j�,�!'�<����?������e׎�'�?q����m'JA(����ͨD!�3�?����䓅?��07B$�y��#]����c��x%eS1�?i���?1.O��7�|��?q�'M2h�2�ѲZ��h �l�Q|.��K>	��?)UJV�����(E$.a��cq��?Y���ȁ�?�*Ol�x���Oj�$�OR�D����.�jTf���%4�v������?1���?�BGQ����O) �:�ӞAR����Ϭmt,����a������?����?��'��D�O���� � <��B!B�(�.�3���$ޡ<)8��;�������V�^����R.��h9�ċ�M���?��w�d�8g]���'oB<O��STgJ_h|�	�ڬ`a���H-1O����O����1 72���I�%0бX3��<�����O|���c�<��?�����f<��aD˄Iۊ]@�ꑱ ���� \�O�D�O��<i`�_e�n�:�.>@BD�G��A~XYH/O��d�O�$9�D�O�D0ʈQ��ƃ_´����Cv�x����O���Ohʓa���ٟO�P��jܣO��H�AħnI4})���?���?�O>����?�j�yr�Ư��� QE�?*F%*��Ҩ���O����O��
� �+���@~�L���*$�	Uߞ���OؓO����O,(��OR�^T����K� s��c�L�=��M�	�����yr��g���������?A�ZQ���ȏ=
l�LA�)�k����H���g,��?�']���:6펌%�6��t����ly2HS�=��'�r�'7��Q��b��L*/x��E�_�,"��������	۟�	S��L�S�'Zt�T2P]^�<2��
((��,x��Q�ݴ�?I��?��'>����d	�&@#��b�
d��BJ;%��J�$���'(��'�_>���H#���!ZD�sw
6o�gK��M[��?���2�u���x�O$�'J��@��9e�2����Պ|�\�z�'��'h�@�Q��h�$������b@#�b֝F,r�@s.�"J���'P��R���O�O*��g�1$�	�ȗJ͔Yh��<�ᆝ�]����<)������O.�H�,�
%� h�P�]�Fx� m�0˓�?I����'(��'dH8bJ��"��e+�ǐ�\Z�`'U&Yэy��'i��ޟ��`gD�|j��/>̊�pD�D|ξ�ь�����	͟P�?����?I�)>R
E35���p6�
���t���1������?�+O���OF��˧�?�7H$�0X?������G�~$��+���p�Iz8�	�n*}��G���PqS:u�J�T����?I���?Y/OD�K��Lk��ϻ�,�c��Q�)�RD��dW����~y�'u��Y�b���7�I���
#S�t����Ky8��T�H�	�+�0!��ݟD�I՟��SRy��ɕY@H��'�0�2��31���'{r����@��y������N,=h���o�?�a�(.�&�'�'^�D+<�4�>T�/؏A�ҡ �C�;W�N�YQd�O@���O^���O$�d�����<��F_VȺ7�P_&���<�ԉ���i���'&��6��O�)�O���9� V4YG�
Iu�H�vόBb�Br�'yB�'���K+��]���'��dLp�Ҥ�ЬS6E�Yp�� -�b�'�J)*�^�`�O��Ox�ـ #GH�#d�"7~� ҝ��@���:��?����?1*OH�S�M�0S��]a�l$_w˒�Z�}֤'�$�	�@�Iy��'���4M�p���j�q!e�W'1���'��'���'��ɔ�F�!��U�6p�VE1�,dQ�B�?_���'���'��R� �IF�t�'1� ��jO�K���!5 �r�|�0R����ɟ4��ȟ��I�>V��ߴ�?Q�S܀T�D@0n<���
t���?��?�.O`�D��Q�i�O 牘5�p	Т�Ӗ
��)�D�ͱ-Gz���Ol���O��؝۠l矸�Iٟ���C�`]R ��e�����:xh����p�'-"a�>y��	xy�O�FeXQ���M|8a��3	92Q��'4��'�z�� Os�����O��������O��� ͥi/�H�X�.&2<Wo�<��D
 ������|�ȟ:t3R���}8H�2�͌6�d��'H"40 �c�p���OL��ퟐ�)�O����O�P/�2XT�����T�@�T�٦�O�`J���OH�O��+�)�O�EC���%SԽ	���;�������������	tB�����P�Iߟ�����ȳ����J��as뀘{��\�u'���D��Py2�܊��O[R�'�b%F:��mp���m�\H�V�ˍP���'�)��e���D�O���O´�O��|��bQ� z$�)���x���'T�y	�'���'��';2Y>�����z@�	7�Mg~��k���p�ߴ�?����?��j��Yy��'/�}��,���&A�����x���
�y��'N��'���'���'&��e�zӞ���C،G������M*a ��FC�On���O��Of��<y��d|Uͧe�""��C�
Hw��|� ���?����?����?9��0�tP@�i���'Od�v쌑t<�y� 0��T�'���'�b^����#[dt�S����kL6@��-�u�c�C�- l�	ş8�	矀�I�d(�޴�?����?	�' ��8���v==��n��@=$h��?�(O ��� ����4�� �C0Upt�ʐ,�t��$ �OF�$�ORX١)���������I�?���̟t9a��R�/��;�d�9vY�os���?Ie����?���4���z<�LA�G_C�r����e��I� �*ܴ�?���?I�'����?�4*�4!�D��mBG��9�4`�.W�py2Q��3?ͧ�?�P�޳���կ�g��=�7��v&�&�'�r�'��C�OB�'��'" �4���t5� ��*�	���'U��'���ў���'���'5 A�����7�L�d�<jb����'cR�I�M�(7m�O�D�O���e�T7O4����R�]�r��%R H�S���t/g�D�	Ο��矌�	T��O�^3�3`���U�I��C�::��l��,p�N���Of���O��O��I� �L�)�̙��Ÿ�� �2\����ޟ��	˟���ߟ�OQ��bw�����ƿL�RYi�HQ5}4|c5��O���O��D�O��ħ<Q�P���'�Ё�l�h�0]jfi[�J�-Z���?Y��?����^2a�JTnß���.5
<�+�LՖDrhi��	۠!����,��֟��'�2���䞟( �-O%O�����ꊠW�$�e��O��D�O����O�U�7-��5�Iן�I�?��q��B(%��&5�>}sRh	ǟd��]y��'J"���4��E��Ɩu�j�6d�,r�|��Oh���O*���.�M��ϟ��I�?���ğ(�hP�z�|q��e(�T�gSXy��'U�!`B�'c�T��U�T&t���2i�-n���0����?�G��"B����'-��'����O���'e2-�sE��q"쌻j՜�@p���;�����'F�i>'?�ɟ h��;6��zl�q�V)��ڴ�?����?!�kI:����?����?���h;v]�؃5�&�h�<�;���?I��?y�DA���'�?���?�$�F4y�����tm��'��?��y|����i���'�2�'Ӷ��y­\%��@�fo,n��m��o����dˋ���O��d�O���O����OL%�!I�^i����
_�%;�c�1a��n�럌�	�(�I�����<Y�"W
�{���>�Zy։�P��,�l�<����?!���?	����$���^֔Hʶ�a��'Ƈ�EDjʓ�?1����?9��s� p��d(8=���*��Y
�*D ho��'���'�RP� [�Ξ�ħD\JA�����d̻sF�-1�:M���?�H>����?aTK�<)�O�e�oX�m�*��Ag�%�
�?����?�+O�[)p����S8���ekI?#��8�1m�CǊl'�<��ߟ�RG��ޟ�'��S�A���§��GqI��(`�.�$�<�ĂܻL���R>����?�-O.%�7)X`� C"K�|��q���'���'�l�f�'ɧ�ORRy�S�»Oi���o]�r۠����1;��k��iB�'���O��O��ďNCm%�+p�uxE	Y?Y���,s~�"|��_�$}�wcݔ�l�g-̩UH���B�i���'�r�΍z�NO����Oj�I�K�=�E靶D�� �vM��3yV�d;��;gOT������O4�$�?;&8�A��76}�S�Ҭ�N���O�!�!G�~��?YK>�0C�BƠ)G&��=�b�I�a[5��dJR��ı<��?1����$��li�1 ������'Fѧ~�`xd��C��㟌�	M�㟈�Iv�? jJm�:AUF��Wg�*,��M�bU�(��П��Uy�@X�&�V�	��t�dZ,J��Ĺ�Ê�&S�	���	K�I������JD�ɡc���iBi�Y&xc�
���'"��'�S���������':�d`P�Ɗ<,qZ	9-��d)���?AJ>!��?a7���?)�Oޔ��˗2�����D���q��'�2�'��I�N�A�M|����B(��=�h��R�U��qc P
���?i��Tل �����SZ�Vr���1(E+K���Hb �� �'N���Oi�n˧�?Q�'I��U>9��#زc:6%��������O����+L',��8��I�.�r)���=/}�|x��֥#��G�x�6��O4���O���@�i>U�E�x]R]��ʟ�|��a2�$�s���4�I��F���'�h����M���v$Q���fӔ���O���ڀsmR�$��e~�)]s��|��Mi�����X��?	���?	�O��x�L~����?���s�̍H#"
X�� ��8D��X���?�Q�>{������ɹN�N�Z���n���q$��c�*���O���H�O(ʓ�?���?�(O�ໆi
�۬�X2�$%�°k�hB�v]$����h�'�  d��P���`�f��]������'���'Z��'r\>�ƍ���MS���_����`G.@_�;����?Q���?	���?1�����O��QE>�z����o���N�4�^X�gc�O��d�O����O��'Ok*���i."�'�@���/��\�,�Q�[#U�<��p�'�2�'�rQ�t�I�Pќ�s6�v�ԩ�+���\��Z�d$�p���O����O��d�OB�y+B����	��`�I�?�� k���#��i���(�m�ğ��IGy"�'N�:�O�V���q�Yq�O�6׼���k�3��(��՟8�	��h�+�4�?���?������Tt�)��*9Eôn�j�~��.O��ºd����Ob��|�ΟJ5 d�&`�be�ŃM>j�\��B�'��	{fCv�.���O���������O����O:Q�U�2H" ��Kͽ8XUJҢ�OFPS�O����<�'�䧓?�"K�"ƨ�3�#1��P�CЃ��6�'w��'�F`p�O2"�'c��'2Û 8���@r��*E��*�k6���'�ɪ���'?��쟔Γ�" �j��uG��xd���#���IП(���Jy^>��	N�I�T�Y��g�@�,�v�Y�i�8�' �� Bc��d�Ot���Ox�iy�sF��,t�����5*�"�n�2��'R�'&�'B�'aL��F F�`x��T�d���"ƤD��'�R�'S�W�%o)���-�;O��d���W,���B�Py��'G2�|��'F2'�~���$�V�br��&M\��ɛ��$�O����Ox�XK�(���$�>��X8���H �2�e��}9�'��'8�'�鑋{"��*U�i��H���4}���Z7�MK�
!��JB$
[�l��ẻ\��Aj�.�
5 �Oy�Խg�$3��Z5'h��B�aY��'��ɷn�z��I���	C��'�>Th�h��5�f$��b=��I"U���I�`�IT�	����ӟ�r�	W5+�lH��J�f>��H�G�Ц�޴���'!2�O��O�'��E��� D���p����p�6��X0�b�-Lɩ��]� �2姟��S�&k��ݒk�uA�gF$=� �mG�~�B�Ɇ!YB$h��@6�`4�C>a��t � \��,�7xp��ƬO ,Ex\���ľ�*�#��F4u���`�� V6衢0�K4�ZQO�B�2���54'T�b".'�\��Ī�b^8��@"0��Q�3�^�l('�ob��SIϋK�<�hϻ%h<`e���T�u�C�Pr��c"d� �?!��?��$��uӠ0㗋Ƕ}F�Ԙ�ط#�X�a��C+I�x��ddF&�`	�H���O#@����cy�H=iJD��BI� p0U��)��h���I@�� `ˊ�S�$�K|��Ɩ�9�
�$F~��UO�^p��8tˏ3~�0CB���q�O��(���9�����9�5a�#uI�B6D���u� U-��pC,�94+3C��T���4���D�<�0+G9s~��D =�K#�	~�WJ�?����?��r����O��$w>��Q�Ѿ(>���W�,�Sf4�z�a�ͷZ�
�pf {x���� �m�A����+���a�I�)�L㗍KRr6B_$lt@���K�'Ԃ���4Xj��BK\�BF(���&��X�
8���'�ўFz����c�>p3Wb�I<z�!q���yb�>B�R1��?<�bc`�T��	0�M�����$y ��O�b�i�����I�&�0EBT���"�-�O���)�O��d�O���*�&&���C] �T�9"��0�CO�:�B��^#G������D<Ot�cak���8C�0x����?!��u���X�~���ӎ	?�@b��d�$���'��O�H2��3@G����L�$���L� ��	WQ�h��i�S�t
3̀�dk���e?��R�}��au�H�'�>�˧��2���6r]����4�?����S
I����x����coA�P4qH�h�&��q(ބ�	s�����E�y@2gd�F�.�����0B��#7��;�P�MS7Q�h���m�V���:<�n�h���۽/�8���B��H��jN���� ~��D�̦�4�?��	�	~3���ϹM�d|Z7	ڍ���?�S�? ��;�Ҝ)�&�RuNȶ�zV�I �HO���f��/X
��PB��i�bt!w�%�~��'BR�_�cv�[�'��'�"�r�ulڛ>�@���-����A���|���ȉ�6M�(f��?2�<��O<��b�22�
�O���$	r�Ȫ:E��i�$�7Y�@���LV;$���'Ĝ�8 ��
KY�#ԧrh"��GL%?�w�џ���֟��?�]1���!�:� E��n��V�C��B1�)K��"��ޯf��I��HO��O:�D���Šݥ��l��	�5Җ����i"���?���?�հ����Od�S�T��AK��]���)I�-BeJ�:n�d�Z���&Β9p�h�G�U(kb|LZ�F�40��Uq2˗�.��엣%'~͢���	7򘝒�f 76���Gy�j�=�M�R"d�� H�G�����Q�*7�l��ş��	b��?庵IĶg�p�{�I0`kԑ�d�*D��{��0��� ���=D^���d%}��i�����<�@�ǞuΛ��'�B�iM Th4\�3�� .����	,M���P������OX�d�b���Q>�r$+�H�7�y�'���r`�2�I�-Z�= !	���O$ѷ��"nv�H��Ap8�S=g��		Eœ8F���#M�#Y"?�L���`�	$�M3��u�F#��uR� ̮)���;"H���~��'t�O1���8�B��Y�7�X�����AlM��ɾ�MC��%Fl�Ty���	�@����I:s�@PB(O@�bg�����I�̖O�Є ��'���c�9ur�8���պ�8�vkQ&>F�$�x:�9
���y�ĭ��!C��'��'j3�U�,
��Z0.C�f,.�'-J�)C��F
,*R�=2���E�����lLq���G.ԑ!����Dʫ7�b�'lB�'2�>�d�
=�F,���E�U,d{g@)}��'a{rꄢe+ʑh�bց������O��E�tES�M�|P[�E�1qF�,�pf��W>�D�OL�D�w?�����O��D�OD�����ܴ �xI��_�f،}s��.Q�Dy�O�RՎԸn��y��xf�Y�dZ(|��\�V�	<8V�¤�q��k�HXw،�H|�>QF	"��4��
"@�$	�/���ʓ(� 5�I����?A��?�۴$*28zINĬ)�	�e�� H"�)�矼z1�IL�R��0 ?
��b���sش s�6�|ʟ���l�F��I��� ƫȑ3��-�v�-�������?��?�V\?i���|*@�įP>��b�F |��I"$��i��Њ�5��ʤ���<�3�-$��2�,T$d�Pe�+��͋�NV�D�J�d����<��Nۦ�" �/���+U�D�|0�l���P [ �+p�B���<������*N(j2�`
£�c2��I2"u�<9gG�6EΌ[��.V���H���¦]�	|yb�2'���'��i��%�ӎj;f�����v�$�Q��O���e��O��D�O�ip��MY�!� IG�G����Y���c#WuK��z���0q�ƫE"��O^*��_�E�uOG>}D�ݡb��'�DP���Ͳ*Ơےc�5O��tG~�B��?A�i�f7��OPם��̨�w�&�&|�w.��a������?��?�S���'��^�|��鎏6�D��N�{��:��%�OƜm�Mwt�I��,Za$�1`�\&����B�~y옔O;�6��O���|�Po1�?)۴��}J���bk�����F&F�P����'i��[���[�n�c�.٢9�d�T>-'>��TJ���w鏴,e!��>1P�٧[=z�(��0���g1%�B-�~zb��e�Hy�i `��QKǧ{}�e��?���?����H�J���nҚrmT|�7DU�%�����>y���=9EM��o�xi����(7'�p����R�'+:"=i&߂SZF`��Se�%����,���?����ɑ�	���?���?�����] ��q�Ƣ��Q���[�]�H�nT=wJ`���쒙}U~��v�'����&��p��4� �Mؐq����F�;����)�	F�^�0���}���e��z1G�&>7xa����
P��`n��,���F�pI��,O��Db��E	f��_��9iU�� >R�9�"ON4����,rt\p���. @�*T�O>�Fz�\>�'y�)�VْK��M��iŶ`�֡��-��kﴑ�4�'��'�2,y�}�	�@Χ5p�JG�VX�)�H Y��a���V?��c�C�K�^���'R �R�%�94�@H�SB�c�2y��nϿ*c< BB�	-W(D0&<,O�t ��i�2|�*�a�T<y� �5!�;�,֦���4��'�6�|�rA�'l�.��1�Ĝ.���ѥ�d�<��e_�(J�-�vkp$����G�v�	Z}Q��в�Ғ�M��?��4G��\���N�&����S�o� as��'�Y�t�'�r�'�"�"t��8X��xd�ӮU�̅�;b���pvc#X���H��7�UG~��K*"XUY�hS�~�8�򫚭r6�x�TI�8 �8�W)��J��ؑ&˘:��OK��?���ħv]������h��C�@���j��'����b��H����8f?h��wń�5�D����A?� �2B����@��sL�� B\0�H�fy�*(:� 6��Ol�d�|rqc�?	�4CZ�`x��g���!!�*r���1��'�I�c Ʀ7d�at��ySD�y�Q>M$>��r�OX>�rVAUP	bAþ>Y��'R�<���m�*���� �ż��?幓�� 6\:�౧ƌ�H�J�>��!G����شf��6�'`�>� ܡo��y���ؿ��|��:}��'�d���ׯ�j
�i�O-~)�1c�ȑv�'�7M��M%�T�;4�V�T ܖ��ܪ@��L�xC��'N2�'��pI��ӫ2��'�2�'�z֝���'��*8YL��b%�(+�r���X)@�|e�`�j��\�&#]�s�v�&>y��y�[���:��ы~� dዙsNT�2R�F��MK����'�:����t�&�͕'?�E�u��[�P+ԉ]�W�x8`�dyr�P��?���1��'�R�'ޛ��N�iJHm����*�di%��1�y2g�NkP����ʫW��Z����~re(��|�����d�8��%s��_�B�B��NU3Cz���`n�/Pw��$�O����O�!���?�����ԏ̡L�܍���](޼0�6�ހ?ʤJe��(�P!c��ǘ_W�yRc\��A*��)'�y�����3Y��Q���S����	�Y��6Y�Z�|ɢ�gN Q�4���i�,NG����4�?!��?����?����?YI|B�\%+������ �o?l�E��M�<�f�ӟ���ď�)J@8�%�B��c}�\� �Å,�M���?��4\-YS��`�%���ZD����'���i��'�b�'-��J2��G��x�ˍ�m�XZւ.��̔�O��1+��^�l��)�f?�%�Z���ϑ*V�b�B���B�A����#ͫ�U�on>)�8Y�E~b��6�?1��?���u�I�bcLd�&k�"Xv�����*�~��'��O�>�f����2]��',�v��4�O
��'�D�EoP�
�5��������V�D4��9�M���?1.��MɆ��O�7MJ���CGH=UPExEkݭ���IXH�r!�m�]:r�D>(�8Tp�� �HQ���M�f<�P%���*�	UU�X���`�y/�8Ө�h�e�}�O��ur��˃)���D-��-+�OH��'��6-����U�O��EH�e�;[���t���uP��I����Q؞��H��,n�a�&=q�.�P�F0�~q��pp�f�Q~����,J@�:S��,iF=�I�4��2%��{s��П��	��l��]�t�C
DbS��+�4�������'���P���8n *l���O,82�>EJ���f���	閭ϩ�~xR�	�rX�b��~��Oa<b�|�WK��3��dѵ�,qa�ʘ$�M�T�iaRKS6e��:�Y���I�M�ҡ^(1��M�Aj5|m8}�u���hO?�$½uu��
�ěG����w���|���ͦ}[�4���r������]��c�o�(=H�Å�C<��;��������O����O���O���'vb-k��ɝ^a�@X$J&N�L��2Y"Z0���#8�l�fǴ&Q��?yNW�6_���"��1�.QadK�x�0I����!=�f�r3(_���M���$�"W��Fb.Y�0h�һS�Z�Su�@$v��4�M�����dV�3�Zw��H���J�
}(@�`$D�py|�i"O�1�Y��T���U��������޴������(��'b�i*"�+��I�\)
a���߫$C����"�O�4�F"�O��D�O"�2��D�]������3&t��ą;6�}���!m�B����PAag�-^gQ���Va :[��}��$�/��hD��m�J�A�Y��C� J�
_���h;SpQ��+g�O��o����90�%ɰ��'Q�2�Z��A9ly��'�B�'֔V���<�l��WjBx?����SN�$ו)�zU��̀]�v`J��N
Y�US���
���M���?(�8�3ċ�O�6��q��XGM*�@�2�C��kI|���l0SC
�1`��ub'P�4q��P���%��S&���1���P9�ٖP��+"(�o��ˠ� �3�0ջ��p�On\���iT�$��0�˒b� �O�)�e�'}�6mD �(�*��tӆ@	��3��mCTʛy���u"OT�
%�������$��2��*�h�<�!��02Iɂ��!��U�2o2W��J�W������ՔD���c����a�ȓZZ�z&�Ȑ�� a�wu���A�,`ݔ0��˓��=qBE�(i:W���3d�h��]�<�"�X<&I(�K�����5��E�<�a�ϋ7��x��$C0�pǯ�@�<��$FXL��+A�a�xL�Hx�<�f��T/R �������	�w'�x�<�\	_�`5
E�X�X��A|�<���%V�sE��	IZ����	P�<I n� U�P���R B�aЕ��R�<� .��+x:x�#[j*|��GQ�<� �|3FX����d����T��"O�i��Y�%#x�T�E
<��Т"O�5�����C�V ��R	k�Ԃ�"O��"��K�V�ƨ�f(6���`"O@�Iq����PQ
r*C4u��6"O��XlݺQ���Ԩ��:%K"O�E����&]���aM�D"O�aaI�)��`�DR�KJT�;"O $�Ui� 3���ZW@�>  �"O|��U�Ȍ?c����:Q%���"O��M��FЌq��V���"OYQf���ZA�u�%��>�m��"OX�`�ʍ9k���T&I�'����"O��#��{�D��u��5�����"O����R(��Qs������Q�"O����j@�n5��0�CL�
��`·"OV����:�8��ƞ)4�i �"O]�T�){�8��@B�'j=�y0Q"O��B�M�8}n�fҥCA��"O¤���I�3��T���^��SV"ODc��%*$P�ͤ<���)�"O,�a� /#�|��Ƀ)9�$ze"O�YG��/NF
��a�ϋGJ�c#"Op�Ij�͊��tYw�J"O`�Be��9aP��2���	�x"O����g�����f)l�^5�W"O� 9�ܥ0�c� �D��< 4"O�a��cL�*Xҁ{3�ېt���4�'�`Q�&:E�`��!Ch����{�xC�ɜz�$�J_"�>]�D�+q�>���B�c��#|RbO���b㈅	,d��D��<i��	]�&���(	1�!1 Kt?�GI��}7B㞢}b��_ k�t�"�ƥS*�"`��w�<���V����b}�R!�Ap���\� ӓb��ׄ3�x��"d�V�ҤJ��'���r�Ο����,	�wL��{%)V)Y�)�R"O0�p"�4<�5ABo�|J���	�%�]����#)h58A�L��4���1�rB�I���Q�Z?�1U�D�}�<�3�p�����L�_]�5��,���+���h!��L�M<$��ˣw��9HӡƏ>!򤖠r/ ѢQ�õ8ۨ�Q�b �
!�Y�%}�8�cB��Z�1A���Py��6VQB,¤璧9ٸt0�숤�y2�ұ)������6R9�C��yB�?���+�5"<*�3��y�,.=s������M�v���� �yr��-b���	g��)*�Sa���y ��@�ZQ��I��
`D�y�^�d��{��zvn�����yBhH:6�R�p�!��A�@����yR�:#r�9��TO���s�'՛�0?ɣj��?f�D�I�BY�uCU".0���Nz�<� �HR���cu�Q�y��)7×q�'�2�b&�f�OKD��#N�c�Ap M�6�p�'�ru���@> ��`���$d,P���
�Cpb?�)�'S����?��P��*�ht��'\�ux���nM�i�@(F ���,O�)�Vi ��=���ì"v��`ҁ)hz�䠢j�fx��
�kZ�����]�V-z�l
�M�j� �A�O�0��I���ȟ*���)�6 ����E
�_����d�8	3�i����P�n0���?h�ȁc��^�nOZ�(eO2z���6�x?q���O^�3@����-�R�n����!0O8D ��?�)�' +&�8L��	zť�tDԻ�i6��*���2B��܈�bN	xu�x
� ��)�� H�� 5�5ayh9��'����l��%a�ы�"�'�=��G�N�@5[�J_C�QzA
O0���MY3����J�)Tx�LӁH���	$V�J٘�cA+b�P��&C.U�P�	+>�B�w�hY�ZW��ȃg�^�37b$���vU ��E	�r�"k>���9ah,�X1I���@x@�K�Cm�f���z�
A누��Y�4H`��-"�F���?S�8�yK0�F�./�J�2��H�P�4�i۟x���|�]�f�3p1I �i��2B� �N[�y�Aï$�xҌ�1�mjs�?���� �yb�Q�2m����P :�| ��f�DF�E���A@�3j����I�C}�IÐȍ�c�����^Аx��ZY�^���+G�/�&O�x��e�UN)�x����%�&��X�^����+�>4Ir�Ҽ�y�!@N�z������a)���0?�D��9�XZ��ؙSr�1ʄ�܈�����Ӱ ���q���!O�Ι0�덝�<	@�Y�U}��ԭ�H��'� ��$gZ��e,�2�P����A�vX��Dlʵ�����Vc��	+�����&w����v�L�#�
�Z�oJ	��`zǊ�oQĨ�:����!I�7c�� 3|be0rMo�t��
%Z�'A�&���a	�w�'R8(ə���0t�j@ �x�����|
��A'�O�!s��^\q1�Ҟj'�q��Z�6/�|���՗QX.��ւ��1Q�I�TFMy%���4"�����j�*V���ú��d�cX�Af��VoƑPp��F8<	HG`�	rC�\%�� /JrcR�r�0O��8�h�g��	:��	�G�[� \| �i�2:#>1qg���\Q��`
�	�(��&�'��s̞�;���;W�&V��9�.Ȟ9���'�|�#��\���Ϙ'$p{DMkM��Á�v�r����h�X�D�:��	��F:Ü�h��Qu�'�Jq�ZH��i��ӖB�&`�R#W�-�x��$(�O&�qX"�&ɓ��Y3B\�HSCÃ�! Rҽ: �CdE�73(�)؃ �,��c�ذ��	&��0hÚ
#:�[�.K�% ���䔓z(]�  �Zu˷�[v�i�ĕ�u���Y���x,�eh@HX�'�`xG�0�i�*Mx�1���e���UDo���q�I 0J���"l��w������z>eR%���*�-��V�1�+v�)��5��x�D�S 
}�cI48� PA�1�y" PE5�ls��3 ��$�ӈ��h84NS����G�O��\@�"O*�#�/Ո!�ꄲU(��	
,2�d���T�ΨY�|U��`A#`O�3_�X13S�ݾ[���ハL�?��݄��8}3tEJ�lߑ44L��@�#��&B��'&�	ac�����I.,�$|e�\6: �[���1�<"?A�C�j争�A@
^5�ʧFb�;%�A�=�Rm!�@r=����Yb$���$ZT�`G�ޡ9gh5�O����Μ�Bq��b�'_�RyX�3GTV\
�f �E�T���n0�w�G�	,f} ]3d%�Ź���Y2���?�'��PaU�ڑSl��S��B���!�'��x�ELH5>��<"���=`���
�'�lY�$-�3x���P�*���
�'�4 $ J�S^IЕ��".�`�'�V	�D8J�6�+�B��n�3�'kD͠�!�+(�[Շ +}]�8�'�@}����TBt[���r�~�{�'Ν+"O :G�$�ڇ`��b�f�`�'�ܱ�@�ۍv�|�z'lEmvj�'�T�IQ��?7�4BA��YˢI
�'��s��Â>ʂD8`d[3CB�H
�'f����I�'j;� :'�ҰF� !�'#�EcN�ndyIf4n�$]+�'F`m!f��'e�� �ӣndn)I�'CF jm &!���뙚d �L��'���{4��L�rh��QǴ�S�'��<�⮋���J'���� 
�'"��G�V�,h&1�mH�,��H<1B�[�9(���d�)o�DQ@,��\�*����]��~��(�Z���B �e_�
w��.x�p(5&D�)!����٠�
����q%f<Tp���� ��8xM���42c�!8/�����ޏ�y�d*T�Ah�k7<�P��
;�ybŞ�b�2��CI��)��j��N�f� �#��O>C�r�I1��?w�9�19E��2{�����aw���̛Y��j�=���!��-�a~�JChi��
� ��Y`��:`�ꂊۦ+������J��PxR�[+G$�	�ϝ@��$���C!�OaSE(�3��ᩋ����<ȁ� S��R�ضn,�yҎK�	s~�{�DH{z�tr��Y�yg�cG�|��G�g��S�c�2�FG7b2��i 8H? C�	� 8����8HY9G,]�91��q��n�;q`��9;��̠P
����a�U�΢��~�(E�`���#��ޭN���Ї��;�Z��V�73!�DŽ@���	Ѣk�]i0�@�p��� � lܧI���UHba�)5Z�I'�'Q ��1�$D�6DD����IÿR�,P���Grr��2a�F<!�DP��=�`n �JU)%��&a��KX��$�>�h5�ݑ&�@�;���3f�bVP���!�^iH��Pu̠YP�R>2���ՇGK9`7�LZ�`V������\7#?� qSd(\O�)3W�I�;@�	�'�&p�#��&�h���bU�Ot��	�'��Kp'A*���Q��D�<�(�{�G��d�^$j���B�O$B����,v�R�-�:-�hM��'<.�3,Y}FPѫ~�cc�?�,t�M��s�<�5bˊj�b(b�A� ���r��]�<a���!���0�0�B�6�P-Hb��#4*i����xB���ۖ�I�g����$÷&`F�	���y2j�?<�D��n��ZS.B�y"矉7 ��u�ۻ?.�3n	(��'v�)��T:�H�E�4�C�Ap�0yw���1�ܪ��y����de"`�B
+bb� ��b�f��H���:\��@Q0c�>D�x	k�@=7/"B䉸���Y ��f�^�B�%J��Y�r	a�Ex@���l�#
&�(uG��|��;�`t��g��S���P��ͶwNpćȓJb��U��G�D�3�Q�PA�ȓy�0x�bb�!j�
�K�ꙵ YV��ȓh}���N�6���2 0D���\uȉ��LQ�V�c'�.f��ȓ2�.1�@�ݳdq�:���$5f��cۂ)��O�n�d	)�!JS����[�z'D��0\Q�CZ%_G���1TF��b�:a�T`^:)���6���� ʴ zD���c>��ȓP� ��O�]�I�b-��)+���C~�xr�I�@10u���ܟc/�}��R� ���Öjq=Xb§k^zi�ȓ$z<�넷.��<�6b�]�Jm�ȓ%~�R�g؀J�6���I>K�`=��QC�	K�H��>g&d��46w(�ȓ'�uc��Y��e�doI2��p�ȓj$B��G�
')�IR�g@,T[���ȓ'i� �T�M�@�*4e��~؇ȓ%L\�۰h̰��(JR�ߤc�̆�Jw\�q�J�8��c�/�9]����ȓ7mv���
�a������(Œ��ȓ���YF�Q8Gx���oH(ZJ��ȓ@3�Xy��^X�ʠ e�3-�����[l*�i$/	�~�P;`D/$���ȓ$�X�8�I.�$kr�=@iX ��E}�M!�� 7FΔ��'�L��ȓ�*��`��6r���B:#����K��3�kZ3m�4��@V�<s�B��+;�c�*��� &�2uJ
�,4�15�Z/�)����<�%b�E���X���3X-�B�ɔ{�m�K��hTL��2C��h�B䉣1@� R�I�d5l� ��B䉔o�~]R�`ٯg�8����Ϻ ��C�  �J!�"Hm*	[��
&X$�B�)� �iY!Ȏ ��Z�!L:t�xq"O�	��C�v1\��tƝ3�ZE��"O�j6�,jPv�JE��!vk�[�"O�R�ޑq�v�c�N�a����"O�	�s�6l�0��UΖ�P.0��"Ob}#1��s��i�-O��^Y�"O>�(J�\�����rT;T"O��Ǧ���~!s�_X��x�&"O<Yu��8s�:%����M�L��b"O��#���6n�là/��!+FU8"Onի6��g$����/%��"O��`�e΋)B��Uh�y�� @�"O�2M?N��CGɄTSр "O�p)�E��x�$tzSc<r3��{1"O�B���(:���Ò-v��"O���)��Zݎ|�oG�S# �pd"O��,
1�C�نl����"O"��$�IZ���  Q/$.�IPg"O�d�d�r�D`
pnI5$$�b"Oj5;��Q<?�8_�3�a�"O��"7�����>pږ�"O�zDmQ1?԰q�&l��oɾz"O~����%���2��[�H�+��'���*��Ϸ�ܸA
_�>?���GD4���D!Ǡ�n�{BlՌ|�T1B�D�:�rHu�F^��D(�aP0|W�E�W�ҹJM|dC&ϻ<�N�
g*4��/�
x�u�'�`�:!��7�
tC�^!����'3NaȂ @'@b��S���3�4�9�J�O��$��-D�ۢ���0eC`U�r�d�[(� ��oG�)��xB$�5�n�zƟ]u�UXѭ� lhD$�0\��#՘_���<��+ŸYߪ�ƎV�  ��YJ�0g�a�e 9��t��GP.=:� �Ot��k���t%�5%!���=Z)z�`pD@!u�z�)4	��A�С���(F�P3�W�az, xN�%�U�ܸ(jzS7B��F@b ��lI"�Ό���'�F4�u��|��y+�Gd�>���'����G��ф�>�bd�+@���jF�I?�2�Ñ�r ��%ĺe��sR
Ǟ��tsU�8O�����Y	\�B8��E�#��EUH�974�97'ϱhSr�G����'�r�Cȕ�+�qG
�3����yr��$ ���ī�5�@e��烂��I1�L��T'�'Eq�t� lB�cx�c`Ū[
���O��]���1��f�V���h��)Ԙ�1G0LO�8�@�(�����!(8��Юc��щ�i̿	.x��!sنV�V�\���"��ʡ����,r,�!4�ԣZۘ��`�@�
w<8�	ӓ-L\D2Q�O�{����g�q7��(�W���l�!z�T��	�0�\Pb�ԓI��PED�-r���F.�@B`�ѐYV��k�`�҅c�O�1i�P� ��� �?A@d��:K��Q�Ŵ,H,��FT27q�)ِY����$��aQo�9"�����x��^�4��H��`Y@%��i��e���V�N��Ô�%t�r(���+LO����J�\����ʎO�`�r�B�Y���ad���͸�G)c��'�|U'?E �,]�<8<�����  ����aj4��x�F�w�x�8Єi��30�#1�A:��'}bhV!Bj�'��� ��
P�H�7Y��`�o�Rg�!�B�-�����'�J�{��*6lM���Ãu��6�9;TY�䘦R��`�3H��`��(P�U��zx4�;?
t��#Jb����c��
إ�tEA�l�ع�U�9}bᚢ4Yz�q��P�Q�x�Q��,O6�0T�3.��hA���ql(q�TnC-Ul1��f�6t�@��'���q����v��Pr7)0��X�{���,	�ԧ��E�V�Q�������O�tbZ�St�ĸU��%�bEi6
O8��6���@@"��P��D�8,�i�P��b���8�z��O�U���Ʊ�t1��O�ۦDai_<	jY4A'����kqk˴h�,�Ʌ/q�$�a�Äq��yL��c`� I�
P�^f>M�����9��$+ ��>�{�䃈8vh܈׎�%z<�&YS)��'tx-8�I]�v&RA��[q�аȟ剸�J 1W�R�Y���I��\��#=�D�/����b!̌��K@�N}�/��Jx��GE�1}:L�Sa
ay�����<�4ѣ��!���������#�萪E�6�p���:�M�f�=5h`@Ԏ
�z@ �PCd�O���S��
?D���rC���~�j �a?!���S/]g���DR�Ech0��*V1H�
��qnϝ�hOB$�m�8Z̤��Q��y����N��"�	I��-ZR�
��D0W�:a�>�;�?Y��.Udv�� l	$@P��	b��E:�`D3��>�.��Z�l��b�! 	H�h�X���J��c�*Ĕ ���/C��Ȱe����'����k�F��CD2�p�0��L�v�b�d�$C�4T��Pw"�>�u 2Eָ��IAf!��utc��n\�!R��(s��*x$��n\�^�,6M2_��y[ǐp�Ќ��#���ў�N&q78����I�=�Ԕ��8m����2F7MEO���N�l�|ڀ�/鴑b3��?0�Y�!�M@��I:-$�� �,F��d�?�$q�!��*�"��W�����tL��~IŞN�x�g�@��ħ�?�7Ɣ�,$s�)�,d.�+��-$�ɳ� p��&�6Ij�o�`֤���"3����'�Ќ	���B0��J��N�etl+2&ދ�i)о4�n�K�p�V�=�X��3���-���y���>��m&��	���".�P�5BF{?1PD�/���	�Q����2##��� �!7������X�"@[��(Į�;hg(��'�|ӼqA `:]شp�%1s䘱"���r��n�=I�x��VJH58�L��/�(k�ؓƎ�I�T���\9@����9�4�#�ψ�5��A$a�(/�P�F�By�)E{�l� ?�H��ګ��ϻ~ ԑ��dπɖ�Y���nr�E�F):�v
�l�E�P�� KG�>�Ԑ��l��,pH���,�:||r��%\����fMt���8���ݺ(��D[���!��O�VE� Ҋ��l	�K+KF1�H�`������צ@}���d�A?	��W}yb��8C���T���	*M�y�UAͭG���Ks��@�N�����������tW:��9J� x�SM՝g�$�Jq�k>� �j�:F@��Qw+�4mp�C���)p)��a(O�T�Q���O�'H��"����;\9��#~�����&�jl~�P�ǝ#@<1�#@�(��''@�=a�'��d�s"C�fg��6�V�,���HVg�0�k�����%)e���X���`��Û�UF��9�*V�A>� B��Ԏ{z<�Zc(��S����2$��컡ˋ�Ƃ̗'H��rb��$A�ҘhQ���OX�%�O�0ӦJ�f�IVF\|$����>!XbD�����q�Q�o��x���/Q~�+��
@�%�dZ�����X��s����pޮ�3�Cd���'閯N��MZ�O\�\����4ɞ?n�蠠ȄU}Ĵ�'6|H�㧋�S���*�0*�M�e�O�詩v$U$$�r��#%F�h�'�R�cHRh׺=PUj��e訫���O��u�'Y`����
���Q�'�A����|��e�^u�%��&p"da��{p½9e�҅w�m #J6>~�Fx�Ow��yw��Ko�ͻT+��dm�ʅxwF���H���i�֍�!�T�W�Pq`V@^��>�/�*6���)Ԃ�[��� R��{����x��#vwr�Y�/�~ZQygC����d�
xi����	�2��q���#d� aԞ4��L�"+K�?�8Y9H<�4MF�~��p�vh�� �$�ؗNE����숿m+�:T��\m2�ޞO��ٲ����1ӕ��#Q����뚠9R�#}	�l1џ���rJ,@�q��6n�,�&P�`F��(@p�s'nAx`i��:�i�ڱ�ƣMQm�M�gĄ���2OZ�עմ\̈s�� 	`Zc>��O�r,P��#7�V4�g��i<ԸB �"U�,1p��ɪFx�=!7��:(�'3�YGjD0dDIs@D�$[ �q0gع5$F�D�&H��K�1��q� '�&`���dD��p~P2�7wG.}ɕ��]ܓc��Hs� cJ����J�Iؼ��O�8�,��9$
�i�g+�yrSl�4����E�X�P�F˓���4:f�+#����"��]�I��yI��iC�������sc^�e\�6�^0�xr��{���U�ѵ,C���5c8J�uoF�[���	|���#�i+\��`%���j����W�=F�F����,������+8��a��$��e�P��r<e���[���`ߒ(��0Z�N����'��s�,zCߟ��h�Ĥq��ڃ!�.	��"�s"x���B\:�<F{�`X��$�
���#���!�U��NLU�X�D��<ᄅ@��?�P͞�q�$�@���Ӛ$���� 4>�����A�*Z�d���!C,c���t��0P�-ȷ�'%*h����?�Bo@�t�Q'˄T��=!V�ˊp���	s( �I�A����qj`���ǖgD
u[-��Mh0��&0&�0+)�Kr4��,ߤF�m g��Br��`(�O�L�?i`e�?Q��ψ!k�.\�U,	06/���w��[}��R��5E�a�
گ?��ʧ�O��Z�B�\✕KEMG�O'|�Q���5��pFy�Ob��IAEW�������-��-4wy�(�,�(;�z��%��"[RAq��;�/�D �7��O��Q�N����������θ'q� W�^������SA�S�5:P�&F

N!R3"H��$9�I� :Q�W�N P7*X�N($�Sq�`����:t��R�9V���!�N�x�+"*|>��T/R�N<�c>Q��m��Uy���ۢu�̼Z��?}��k�{���_?Y�P����4`��	Ii��_�;`8a*��Z3A�l��́&k�d��F��d�� "�8���-c��%Ʌ,W�v_vh��On9S�i>%ˁ$�<Ѵᙸu�Q�6��Ym�P�L>M���IT��+������y�3dT�G�.�a�ϕ�R5{���/)�<���� �eȿ|B��߰>�@� BI��F� ��"����Gxr)��4���E��E� 
�M��?�W�Ii�%H�=�T
��qh�z�$����$tӤ1�G�f>���ϥ^�*�zp�~jq`َx�L�äl��h�� �ԆV����ĔJ��:�N�+"Llh��4��h�@��>%���է���l9%�L�8�U����!̶��g�c��q����3Pa:�ĺ *U1R�-O�As��P/Pk��@ʰ����J &h��8%!V�K#����i��`��Kj�')NH���(&: ��0�B�G�!%�����
�P1O������>���O�J�AƋW#) )�?!Ob�y���r�u�t�S����:"VB�?��'4h� 2��o�U��k�	�
��Ի.ҌUs����%��rq��mZ�:7�D��bޜ���S&~�*��O�HI;��^�f֩��gF�'���H������T{en�:y�f�y�'l}ҧ�)wc�郷��1:�p���=�άC
�b�ĝq���4�iٗ��Р�)bA�9oJ�)�?��CE ?�q��ƶ�hr�B�m�T�z>�-��@E�zL�%�O��5eѦC���'3)2+�9�jtzv
�	x5����S�#ړNON�2e��F�f%P�������mѴVV��r4��)z"��4�O?�����I�\�S)��,����V�6Qq�G��u���˔f]�O�nI:�]:IS��xe�D´~�^��&C�5�>��!�\�6i剘�V�%/U�!V�z��|X�L��e�zBt[�h��x� MڶJTF�lzX�`��C��dKj#t��go�Q��a��_�m�<l�6e]3xvƑa��I����B���J�'} m2P/�4N�i�2�����PMHN��U����5#rȠ��
ݔġܴ
6����nTn?��EY<
�"<ӯ]����1C
�r��P ��d����x�(I�D���O8'>i#�gJ
1c��g)r��C����'�'|+Q������Z�#CN�}�4���$�@���)Bۜ!�G�o�``�O�0�fP���	���M��i��kS�V��, �[��@ d�XܓmPD!6L�<R��al8�$��'4&��UĆ�Z�j��� ;�V|Z�R��|���G.%����`Շ��ף^9���&�O~T�s��u�6|@ReX3;"t��ې[����fe�'dՆ4��)RA������,)�oB�J
�P[�KR�~Ő",�ܘ"D'ڔ���.=�� P�@�jW����V�մ[��İ�A�%!7Șx��� fP}Q@�Y,����t�qM�"9|TD��Jj�f��ӂ?��H��jʞ�����V0#>-��i�Cbۼ0'�6�o	u�S�B�3��;4��C�Ш�`P5~U,�Z��h�{��8/�t�W�B�s���߅� �O�޽��Í�-������:�IY xI�	G��,�� ��'�޼�ˎ) c����L�
�T	���9:3��B��ں:qεyL��s�l��5�1Ol j��F�����5~6��Q��B��)�i�������j���goR	[5l�$\�#Uvd�O��#�������D��Qǘ���+0LO�8�"EO1L���Q��'|��v�'��5��*P��Z1Ư\0*�9�&E�OԊբ�1��i�����D���@���2醽R	�L���jf�	Q?�̓���P�

�7�͠4D�o�0�j��0u-�
u�'��������S�Y1Oz�J�ŷ$�hA�$�μJI�`ۂ�$=(� �p`�+A�OX�!�a"��o.	`B��-�"ə�(�7�80��� f^�!��I�\��6B? �*��Q�_r�p`☭><IapS�6�Թ���x�F��e�=��C@�L�Qʗ'�?�$"**��|�VOųYR����HC�<1 �L2]�䁱q]�|��5�d���<�1F��ň�DM�F�2�\Y�����L�8���O�x	[��E0*��+L�8�@���4��dB�BB<ZʖHI�C9�T҄-Mu��0��c"D�@�8S�� �E��@["�<D���fA9��A�G�����8D�$�S U�f��3��:1���-(D�l��i��A�����G0k����L D����i�/H93R)G	s�U� D��{�IT<�.��3�R�^�z⇅(D��"0G�'���ð�q ���Q�:D����
�CӰD��#�69a��j��6D�xѷ�L��M�5�� \&�˗h3D�X�N�|�M�F"�q��Ո�F$D��*T
=0�H���p��My��?D�<3�A�Y|��H��ʮyrA0$�<D�Di��݊s�����$�"P
"DCC�;D�8�g�zZ�U[4�ħH�I�g�;D� qh��� ��k>.� ��.D����AݛN%�Jr�M�9��"D�(qң�
]��<��o�\�����=D����@� (��I�dQ$�ι@V�0D���p�D6�`�C2�N8n1�e��d0D��7�P�ql�ِ�*��5��C䉦t��{BmR^�ċ�C^b[NB�	�}d�LHV]�]� Q�'_6PJB䉣<�"A �c.Xs�e ë[�YMB�	�O)����5�-�2[� )�C�	={�`( k\<~�4 h�2��,D��*G�Y�!s>�'��7D��}C7<D��[bڟ������<2�j��9D�|�͏z����>�LA��	2D����B�h���Z�a�ᘴ�$D�,�V�ߗ4�حI��/s�!{Ў%D�� ��č�CN�4�O �$�4"O���	��{mU=��"�"O�Qz�M]�UT �,ـ_�X��"O��EԿw�Ar���`�|�q"O�oNKz�ɰ͝�{��9 ""O"���PC�Ӣ�4k�P,�a"O��R�,W�p4�)t����AY"O��ʘ�Un|��	�o�rD��"O�Ţ�M���Ұ�W�^��lZ�"Oʁ�d�I�l��A�&�Cl��"O���,$[�R�b�4o5��XD"O��[g�הG��B"�l�6��w"O�,��	Ow������W�Nm"O΄{�kB�vt��#�ҹ@���K�"O�j���0
n p�n�n�=�0"O���N�9Be}�F�Ȩ�ҵ"O�����$J��ڂ#�9[�Ƶ�G"OI�׌�!w­p� @� �D��"O&4��@>6JY��oZZ�Q�a"O���a��"#*��t��<f[Ph��"OB�["))2���@bD�+=���U"O�
K�H�v "�l ٢�q�"Ov��fb�	Cܳ�m%1�0�#"O`;B��E��dʲ�_0y��A��"O����@<zP���jC�O�~�z�"O��qAʘ,>9ڹ*��3�|4�S"O�lF�44h+�N,+cp���i�<����i�3B��+w��X�eGe�<��$�a��择h�Q:"�c�<0�+0��U��@�v�ʅ��Y�<A##S��>�ȅ��!�4[V@SI�<q�LM�y�,`�J�Av����B�@�<ԏ�x��0�V��H��)`Ң�x�<���7L��y�o�1���u�<����=+�����NT/ڔ* L\s�<F��"M
 0a��t��9""�p�<��OИc.�Ź1�Ś��̱�)n�<)��˩!���*�N�)mea&i�P�<���/+]Y�_z��@��H�<ᤋP wV̹fA�:��d ��{�<�֯ε���J�NӀj8�!@a�z�<��%�(DHD�5\NH�ȇ��l�<A 
Z-i�z1a=��H
�(�'�T`�/K�Y�BPb��\���H
�'Pl�QFCT�~&Ha��V��hq�'b$#Q�ޛ*	z� ��!?�|���'��py����{>\R恆� ��L��'��\ �G׋ppv��Dōtz���'���B�&{��8[a�L�b�B�'�5+d�p�&-k�+đJ�~�
�'�r����wʖ}���HsE��`�'�\��G��A�<�2v*Եl����'�Ej��d*<��8i�K�'��(�s.މ`���DJ	T�I��'nq��"��'}�Ts�ȗ�Az�'&q�	\
H�8E밆� }���'��Y7l�/�d�j�P�x�Q0	�'x8���%*��iPJ��vk�@��'�~$��-�9Z�����'k|#�'{ ��'�ӈu�B9�S����*�{
�'
B��"˴�*fƁ�'_ l�	�'R��2&Vx��U�Z �8�'"��`LZ%	?�\P%D�3#����'k�������v�2�ƅ�0Q1��� f|��O�{t�S%Ɖt�2�"O�y��\�+����U����Bc"O�l·��+E�$@K�;c�X�"Of���MI�v$�PRUH�H���"O*�x��lE�	�%.I;r{�E "O�8�`���\�NP�׮ѓ;{(-��"O�ԓ$�J�SM6�G�9`h�Y�"O(L�W�׹~�ёB��Z:�0�%"O�����A#40�CB���= �"O��"�(\�7dԺ��(�.���"O6 4�ܤ3YJ<(6A5X�%�"O��3��%7�b�Kga :K0ޙS3"O���0���tR ,�捂:"0��"O����͚!LT�����-`S"O~9r���!����$���H%b�"O�)S�H�J#<���lI����rs"O*����S�=���xSk,q�H�"O���w� {�r`)�O0��q(�"Oz�CpVO,)�GL�&\���"O&5B����6�6��f@ȡ8���4"O,h�C�i���´��'E��"O�����H�Jm؅ ��6o+�$��'�j�C��(U��3��!�>X�	�'��xQ��1�=sB*�9�� :
�'A��C��np��Al؉<c$��	�'{�)8
�.�`��3j��h�'�0�s��Y68�rQ �b	6����4�PxRETa7�%���G�=�8�� M��=��{"bQ�j������IȖ��PI �y�
;|��@�B2�Ҵ�з�yR`|�����-pJ�  �yRbģv�!�$�Z&{�:�ᘕ�yR��q�J�;��pQ �����y��Óxo�x�d�ûjd�`���,�yrJСo�a��i�8��oA�y�i ;l| Ǣ�Y�v�PW,˻�y��So�Xs&��(�)h���y�&�Cw@�HTh\�z�H�Fp�<�����*aK�A�d�a��H�}�<���:��u
��Ð9%\�yc�Gx�<�Cǆ8b´2�,��O����v�<���,����d��U�j\u�<��b�O����IN�n�� ag�<Q�G�3��h
��*vl2��"�X�<!ף�Q5�yU�L98�0�G|�<��k�>Zz��6��$_"�����L�<���g;z8��]7zԩz�r�<a���(� ���5:|L�X"�Tl�<y�B��j5N���Ήq΢��!l�k�<�g"K=w��
7�.�6���A�n�<��s��[����x{�q1�T�<	s�ހ6�Ds�⋙R�2�a�O�<qO��6x�A�V�Wl��� ��K�<���H�(��B�e��RcIr�<��o^$t�`� b/V�%|��ƈ2T�,s�n�7+`p���4V���!�+D�HP��š�*����C>V,��Ǧ(D��s�n��ku��1�JA!F��<
�%D�Dv��8~<�M#�$(dؾ�8�I"D� ���t��e;���T�\@�h D��)S AZ\�{�G1k\ب��?D����#_m�pU�(ƕv>2�0TK=D�x1cgY��L��O26�ӷ�<D�$����)�>���eύ1� �Jv`&D�� ���h��$~8��uO�v�Tiӣ"Of���"!"R�'Y���� "O���i��;�4jEF�iB�!"0"O mhgN��#{��!$��r8ڜJ�"O���SN��u��\�0ʚr���"O�iSg8I��1��E
v
�R"OF�ۇ|�Y:Pg���!X"O(�aC;A��8W�'��\�B"O
8��	�@���uF�g�>�Z�"O�à%�>�>��QkQ�4�"O����|th���R�a��*s"ODy�G��}N1���'Kܝ��"O�4��g��9 d���˘�F�@i�"Ona`�m/#��T��
��~�r��"O��'ҙ{�zu�2J[�)��ܳ!"O�1Q�C�3�n�ij՞),4`�"O�Q�����8��q#�)�'�y"�"O�I��O�/�z=����~*���"O�����;�J��@���*"���"O�����x>ճ�"+�(9
�"O�y"�a��:��E�	�9S"O��2GP,Ra���*�x���"O,hi��L&@�xY���>Ԗu�"O<  3'Nx@��	�~��Y*B"O��C�Z;8��6m�����R"O�2���}犬���P��V59 *O$|��G�ucĹ���XzV�A�'�P�a'�N�o�:��S"F`��':�̣VB�GJ
��A�ڝvk��z	�'�e��*-"a
%b�H�nS� ��'k��D��\�0�PlɆ3װPQ
�'�0z`#Ӭ?�d Q�F܉P��	�'ӘY��,]&��L��>�x�
�'��qi�׏>\0�26jK�@���p
�'^ `��E1`�P�
٦7a��K
�'�A�aK�1K&2dA�	;�4]��'բ�h�8g8���b�6E�(��'`|�gA�Z8
�@Hڳj��m��'���q��2�P��fJ	 �	�'�֨�gFˠ:��	��I	9�����'�D@*C��"6��@����d��(�	�'X�T�E�H�t�U� �_{`Ej	�'��xp���Ci~�B�XJ1��'�Q�I�04Ć��1h�pM�E�'�T�)/-B�L��l�h�DlK�'�p��G�aV#��C�]eH	�'5�4a���?����mXd!��'�*�Rg���J���#T�N���J�'�*�@�Ӥ��]K� �NYx�!	�'���	�����8���px4ib�'%ؼ1��\T�[�l �m5����'��a�UI��M��Г@l�xD�'G��cG1+�H�,4��"� �y���*-[���*7C�Q�D�;�y��3%�"��D�-��LР ۴�y"�),�D����ݤ+�z����Y<�y2#��N��F��X�2-��y⎀5k�.U��].v��tТEȮ�y2����j�qfkް/��!wR��y�*P�4��IC	H�jJ�m�F'_8�y�U�kQ�D�	b�X�h�y2X�QN��f$O�I�<�K/��y�`C�A$�!�A�q�p�Y��K��yR��(v�CqO�p��x	�����y
� ʁ��ӵmeP����=>�ȥ"O�p��'I�~2�9ǀA#eZ����"O��+���$��LY��(w�@I�2"Oi�1l\=�֌���}�d5G"O�}�BnF 1���x��ܶĢ���"O@\�d䌢p��qcV쌠�F"O>k���3JϚ !�� �JS�� 7"Od��Dϖb�R4i6GӦ�n�:W"O��E��
j�e�)\.�@�"OP10�E�)�bQy��@�	�(�ѐ"O�4��	?�����ʻ�6$�E"O�xIaB�{���z�Ǐn˒i�"O(�2��|����ۻY�X�
s"O�P� ����4,���9�"O�P����3�+��:W ��Y2"O�}�ҭޡj���j�$hX���$"Oؽ�2��h��l�sjD�rPJy:�"O���v`ݐ$�t=j%)�!F7:��"O&�%�D�("|3���(	��"O
��������Ir�
��af��"O+��2R��tF�*j�+	�*!�$��K�*@+p�4V�ę���G�!�ěb� ��%�� ���x�e�	& !�$0;H�(G%;�x���cX�h�!�I�O�p3�,!14�� EF?�!��U�-|N!�3��$-�	�DL�L�!���y��مņ�C����wc�2Rr!�$!m��1�E���xIq �::k!�dV�~ȁ1pG^�~������(O!�$�#WЮ!�o�}&�P���'�!�$ԓuU��jAꕁDn �æOU�!�$ߺ~�U�D�:ht3!O�d�!�$�
��s��>�u
�D�Q�!�>v�4Apr�7#Tta�$ 5!򄕄;� �`�.i+��r���5!�	ĪD�P�d)0����sv!�d���t�V�J�9)�5KGL�>a!�]�/��0hb��ebx�t�@-/�!�ɝ�A�d�[е���!��Qa��*�%�F��s%>p��~�X�x�tnA�-�&�g.�IB�axդ0T��ڇ��y�:���+B�:�s"OR(;���%��#t�T�c��]�<��"��=�C�8%���k�j]X�Ib�,�ɔX�D���HJ.C��"�m4D���r� �_�����J%o��y�P�@F����e�'wr!�o@���?Q�'�R0�pDO�i�5�,
�5���'����@�I�v¸�3��-d�8���=���"�́�AdN ��&�X2��g"O��b�'�-H�Ҩ�T�T=N����i�"B�I3b\4� 6Cy�
��^�t6���$�H̓D?��!J�1F��gH�0%���ȓ�ʙ�q�S�i�5(̩H�q�ȓex0D0%��x.�9�!Z����ȓ�Y�C�/T^QZ�CY;e�����AbJ܋w��D"����W?�-�ȓ]�0��f#�Z��-]E����$hh�� ���#1^��Q�Q3�Y��M.rE�X;M�x@��09���ȓ.s�b�՚W�5qBҼ��ȓ	��e��E��K9n��u�6 ć��d5s5���i���*� L�)SJՄȓ �Hԋ�KA$T^2�b��K�s��8��S�? ��[��;dz v���-�(��"O83p�	?[�Ib�ǏJ����0"Oʕ����g���O�	��"O�8�#�~���e� $�XyF�']ў"~�A]#<P����
"l�ԛ�e�+�y�o�3&���eM"%l|�V���y��yI($�⅔��e�D��?��'��qaR��	�g�(D3�8�']�lYÁ�&;�E�F�Q�R*�)#�'��zt�~=N ��b�	N�$-��'��9�d�O2��|0�&R5L.��2�'�>��6A$@h�r��4�eI�'~`��-;IQç N <`�%�	�'O��b�#~x�V�H�.紅1	�'#��x�E�g�*�L�]���Q˓�(O%��?Z0u����i>tH#�"O��Y�
~v.�25P�z��BA"O��4��4D#L�2�f�Y�<lyp"O��q��+!�L�S$U�|�� "O���ޟ)h�誶�Շ�b���"O~0��E��G�6���ҬwV�"�"O���&2L��W�Y�?7~��%�d)LO��A˘}8���F�ק8,t=:"O�t�H67�b�!C�G�%*��[�����>C�
��c�%�b��T䇾cV��d>��={&��6Dؼ����F�|0C��48(��t ��EZMӓ�D�C�f��d;�I+Gn)�g��k�yr��ϗCD&B�	�;��l���S	���sg��(8�B�I%}����#�M4V͂� n2��C䉱Uh@�+�$Yl�nz Ϛ+N��C䉨A:H�B%C3���%�6��C� G��ē¨�}��,�9�vC䉕wl�P32��s5D����/*�B�	��zO�	g�q5�؏j0C�ɿQGd�i�O%pp8ECW���2ʓk�Qx�OU�]
^,h �>/�tȅ�P��X�1'O@�&���;21��O��=�4�рR�I3�U:��p�.�L�<a�ȁ�hL�DwK5�D�r�L}�<���ʚ6�����0Q�N�Z�j�w�<��
W?	2ФK!�ͷ[�)��Ys�<y�D�����K��t����MF{���ibX
�DH(����9n����'Q
9��g�^Kx!�'I	3�f�����1O(8���
@�}2��) 2v�"O�0����Ie^xx��݊X���"ON�r��J�w4R�8e�6C�H�z�"OdeKů��5���P)��H���ar"O �@����<t�S(զ5����"O"��ɀ3�A���)>�<{�"O<���d�[Q(XZ�kE����"O>-���V/R�0���)�D ,���O�0¢�8^�p��7ȇ!?L�9���r�<�u��Y�^�JG.Ѓ��(�V�Ft�<�@m�Y����3Ləm%t4�CH�<i扔s��9s,Îm�����B�<ɕ�ڃ^3x�r)�~:�R���<�DcۯI��#DĀ�]���Q�<b-�:P���Q!�45�$���X�<��AJd����4`��`�4��L�<����4>��u�Rd�!�0���K�G�<���A�I�sH�q�6"��VA�<I���uM:E!���B�\8u���<� ��×����kAX�I�c"O�H# %ҿ<?��1�Ƀ�8�8T"O�QŮ���|i���8a�̰ �"O�(z��ʴd��j�Hҽlsbe@%"O���D�&�6�h���Z�}��"O~�R5�p�D8��Α�*k�j�"O����		�zf����1:�	�"O��i�,�0S}�8b'L�/Z(�m�1"O�{��7l<.�j$�N�O��x��"OX�K1^�j�1��"���t�'�ў"~��l[^����G�g�r	�$��y��Y�b�Bmb\:��%��yrK#���J!i���,ж�۵�y����U���CCL/rԑ��nӬ�yR)͘9�6Ȁ�O�+s>�q�f��y"�=^m��c%,�<l�"�f��:�y.ȟv�6y�1䍋8%~��R��y���M
~�:�++�B0Q����y���X���؂%DS�Z�k�-\��y�¬K^D�C!��J�@���l
.�0?�-O����(H@��6�E� خd�B"O�`+���=�~AD�
r1�ac�"O	�R� n@� �Y>�S"Ol9{"ұ	^Z�T��4U���"O���A�_�Tv ,s#�?>b��R�"OL���T,<��3b��Ia����"O=���"{����@G6?���a"OiA�Mi̝A��.r�|hb"O���+?|��� ߀	ِ�{����0E��IE�S�4���(�.g4��A+K�yR)�S�8��!�{r�Yb+Y��yN<=��P�ؘJ|�P��з�y��-&�W�=�1�:��C�	�A~\$82  s��M�Q�^�I�B�ɻ$��Sh�i����ŋ\�A��C�I�ON�|
 ��	,q�� �(J�C�� ^[�ЪQ�M�\5r�+3��	�XB�I�	�E��L�E�� F.]3AjbB�J�T���A�v���?>��B�I8G�N�{�`��_$�zEG[�>��B�IX�,��$��t$P���!�:#$tB�ə{j4L��aî6c=�dFĐ/@B䉇�}�e�j��dY���{�(B�IF�Uu�ˍ%�0<r�$]\�>C�= I:�J/�l:�����F�C�3/P��pL,[5؁�0�ؐJC�	'l�d [�V�-F�����%*D$C�ɱ!A����I����2�ե_
�B�I12s�M��BK�<Mpp)C�6��C� \��7�#���L�%O�C�I�W���@­��E؄�#J�j�C�I0&!�REɱ^Ur��a=es�B䉆P�\�����M<��X ٴB�ɥzD�3ǯ�\�($��&�i�C�I�����a	R8P����WFW�drB�I,��0
d䕉 ��x	WCӳ �fB�IgT��m�x��:5Ɛ�PB�?��Y��؃Z�D��A��NB�#Nh�pqM]����2d�6:FB�	�S�R؂��*d�r��C�K��C�Ic�
��G�$a�b�;���=�C�I,e �Q��&g$�+��_4�C�x�^�R�C#;O ���${,C�	�8�@}شm��a�(����B�)� �B���5�J���R��d�"O��j�-�*#ߐ�t�S�X4�z"O�h.���i��"=8SF���"O*Q����F&]kւ��|H�i��"ON�h�1w�V����6_5�|��"OP��W���k�+M�1��R�"Ob��v���4�)$�N&_-`�"O*��` l�<<��*��$H1"O���pL+��;��9X�h�3"O�0vΜ�R�;�˓�y���(�"O8�8�dA���I֪G8)��E��"O���t��5�V��R�_�	,��6"ON<0ǧG�F��y��C=p���"OVI�0�Jn�ZA���DT��"O�r�(52�L�0D�(����"O~\Y��2W�,��CA2[���"OܸkS�K�#�e�&"/����f"O@���V��IaPG�
I8""O��d��P�,��3�M|b��c"O��PFnW�s�ȑz7e��٨���"O�(H���8J�`�a#�39-j��!"O�A!ʝB�@H�1�6��1�"OΘ�al��)bH�G �$���z�"O�i��쐲@&x������f��%"O,����o��c ��q�|(�"O
=ɑXb���С�1��9Ȱ"O�m ���|����'*$r�d(�"O�4{�)̨�p�
4c���°"O�D�U�
�/�����)�9�"O��z�"]�,����4��	Bw���&"O��t�U1t8iRO�kq�myp"O��%��8��}�Qn�kkh\�"O4t� �C.n�rXI�� �9_�9�"O�\p��G=L��u� 㜵fAx���"O�<y2�#`j��B��s��"O�lCq[�xES!�L'�L3"OH�A�D�15���A
۬ft�ك"O\(1eHv6<Se�=
Y���P"O�`8�W�5�(E!���wDr�j�"O8�g&ړ$��F<D����"On�[���*�� ��&�7v9�X�"OT�ڄJ�)�P1'c��8�I��"OT��e�	r���(F���%6�'"O�,k�!RZȣ1�ԴS�,\H�"O�Aac�1����ffV	E�xyc�"O@��sD\�nC��F	m�:(�"O��36�A��4�q���;e2|4�b"OP0���* ��O��*BѰ""Oh!`W�P2��1?"}!�"O:�ʾO����΋�aZb��"O ���2�,c��7��d؂"O�4��JT6̔�m��w�xii�"OF�1�M��?�������`��"O�k�l�s�f���Z.<��pX"O�̊��
u��뉒f��8"O>I�u�\,M������ń�(�"O�A;�m��J���b
	�:X� xR"Ol�S��
9l6Zp�\R�	�"O��R�ٞ���kuɝ%B7��$"O��Xt�Q1:Μ gL
�a��"O��!�N}��Q�f%R&~��"OD��4��^KJ���ʛXS\�ѐ"O���&��t�]����m<��"O&!pp��9{~dyԄ=m*��Ru"O� N��P$L0K�h�ڀD�t"X=��"O�3�K��	1����XiPMӠ"Ohex5
H+$D2����J��"OJ�[2�0�.h�EM�s8N4�E"O�p������6��3U�t, R"Oԁ��#�1�t�)�� ��"Ov�с� ;dQЦ��"I��T��"O(�S����cd:T�f�:[�֥20"O"调� �#b0q F,k�0�`t"ON� F�	�R�v�� o�c��Q8�"OV�7�%߅ɔO�Ґ� K�~m!�dI�ir�bc�)0f<R(��4]!�d�O/2ݸ��,L�q�G��8x!�$�ӎ�Y�׍m7P�h'VU!���=&h���i-J���иY@!�DXt�ȴ�q��q�lz�S9h�!򤎤���O])��J'#�+�!�D�[�:p0 _�M�p���ǴX�!�Ď�o�4�W�M"� {�"p!�d�/	r���Zz ��dIW!�ӻ=c&Map���Bn�rV#�pm!��"Ig��ií;�f�S�V
T!��Y�R�� y��߯a]6���݌lM!��B��� ��UQ6��f �!�dD�.��,��㈅'Y�5*�#S�9�!�$��1o��@S��,Tt&-� G0!�D�	��H%��8!gN��� ��u!�D��Hl�|�C�Ӻ1R��`/��!��*�"F˅$�Ѐ�րX�(!�dL�
�hu�G�H��8�����'S�!�ē�?�:%`��O�<�;E��2�!�$]c ��) ��HD �7H�!�d^�Lڨ��dS�2Ot��0/��Eu!�DZ�>]8�X��W:&�¬��m�%h!�d�7^&,l[�
2g����+K�R!���v�
�k�U��EQ�a:Q;!�"�貀I�$W��ejI�
!�$�'�ZX�I�5,ȭp6���!�ܘvn�#t�+g�B4b#ꝤU�!�\�jeJ��C�F�n͙a	�%�!��4T���W�U���ې�=c!򄕑h�(s4�<2�½9b�W��!�$�0 u"��I��aI�Fƌ�!��1�D�' 0~� 1��2�!�<t�h���K��%��mV�$!�D�=6ސp���3�T�"�!!��*1�\�r�C�����f�!�C}b��ы$s��X���z�!�d
� xXY���K_��Q+I��!� �h�n����*_1*�:��_�z�!���]�ɢ4IB�Y�b�i�i��!��W9/5� q�gR�/�ͱ4+H�(!�d9��T�w聄>�<xҠ�x!��\�9
ZZ�G�;�q"C�2s�!�d�.Dab,�&R�ʩs2b�K�!��$j)����$ 3N�A�q�t'!�$T�PX�KE(ݿ}Z:�z����'!�d��lJ��p�&T�]�3��!�$X��|����ϟ�$L�v��	�!�D�(�b����R�Y�a,�O�!�Ė.n�ؑ)��X�)s(�U�!�dQLд���i�.1�`QBh[��!�� H���q% ԉf�^����Ե3�!�$\*�jl;p�Ļ
ߚy	�D�*�!�� �s�O�.�#d�A�>"���W"O���i�1MZ���`y�-"OV�'K�/����T`�Щ+�"O.��eΒ�@�"E�$k�$b�j�"OfiS�i@�?HRq�?	;~���"O��CA�� �����H�*)�tu�"O��T`�<[�֐��m��U+�8p"O�U�oO�|�0�l=9�X�"O>�x/ղ�)��mF����0q"O.�H���?I �-XҍOB���"O�Z2Z^�~����2�����"O�,�݂[�6�
�i��1;7"O|,*�/M�)D4ҰiK�+��1�r"O MK��#)�����ӆ9���W"O���5���;�e�_9>X�"O�`@$�16����都#-@Is�"O��Ѥڠs�<<+H�%�|�r'"O�p�U'��~���KBg��%�&�s5"Oj�bp	��k�Dj��R���d"O�P�G[�k��)Ғ��"O���#A�9!������N�z�d̛�"O�yKs�ŷrE�ѪZ�{�Ł"O���	�:����2�"O8@`���)c��<�"���v��9�"O�LA�L��0����_�'�2�2"O�R��U���D�U�(��ŋp"O0�@s���%��z�h!�"OR��Cn�&t�Bʔ'gCȨr"OJ�� k[Q)X��c[@��)�"O�A�ԀI0R�e��L��R�"OT�PG��2M\�n	�dPl��&"O�aq'�A�u���Dl-=�yrf"O���꒤.�¼b`�!���20"O�Fḱm]^�X�ł�=��p��"O��r�Ó9RQ��7��?���v"O�DK��ȶ�&�b�%	(s����a"O
�r�� "�*-�CG�
v�T�"O���+޳%��q '��+K���"O~��㣊2o��Qae��Ѡd��"O$$4�X�-�6�㰄�*F_�%AA"O�DC�jԙ��h�!��9�"H��"O��G(@�N&B@�3��aЕ"OԚ���a�Mp��Ҏ8�^��"O���Y�j>�����V@P�h$"OR�P��rI�ł�9��\ �"O�HCFc�(���)ßR��a�""O�1� �M#�n�9'��2v���"OF��_�s�8mh"SoPl �"O�q6�[1t�J0kQ��Uܬ��"Oۥ*ûX����V��'lk�@G"O�92f��W�&y9U/�	 j��"OH�􍛁1��e�Z��z<�1"O(yaP�/���wd� 4���i�"O����R�1�tm!u	�  ���"O�Q��+�vTVc0�M��"Oj����+��EPPC�c�&"Od,{⇁qUD��1�ՈN�0y�"OX����8y
G��6��"O�@��S!0����kI�^42�7"OX���T��ӡ��),�!"Oڐ��BL���o_�/�R��"Oeaea��,B�\9Gԍ+��|i�"O0�� E�GpIx�,S9�4,8�"OR�٢��eᢴ�	��w�D�"O� �UKQ9��<{��S<���"O��A�Ɇ��R�l>^�
"O�9�끞*��嘁f r�3"OP��@��g'��@�T�G"O��!��Ţz�vj�	C�6D��"Od9zbA�	v�DR�:�0 �"O橛�F�PoB�a#ߠ"���A"O�8�i�E��	�@�P����"O��F��d��U�B?� m·"O`�[`�quB�jǲ�&萮7�!�K7	��(K 
P1ʭs3��~�!򄆣e��� $_�8�2$Rq$ܺ�!��V3渘�s��2���X|L!��ʿG,�K�/�5tH`���=!�$ bK�e�5�8 Zh5�qקhQ!�DhX���
Ȃ\����@�8qf!�ȺD�\|X��@�&;X��K�2~K!�$�$;p��m4����-~!�\�����d��7I~,p��(
!�d�iX�g�JU*0�,t�!��+�QQ�O�tR����˘��!�$CX�xh�V�W8Pεx�k�G�!�Ę�)f�+uȟ���qZ��2�"O,PE�Ϩ i�����M�r�"O��J�&	�c:	�S���2�)�"O��0��#bJP�S�ی�$A�c"O@l�䊚#���K
l�B��P"O�ٸ�Ă'c�ЅySCv*i{�"O$�9q &y:�cT7n^\y�"O��녩I,P�<�֏"��)�P"Ob��O�Z��Q�H�	r�zi�"O`�J�j�PϦ�j�޿&T��"O"}cS���3��<����Y��q "O��p��Ϫ�z|	�$B72�(0˄"O\��D�p�������[y�x)Q"O.u��%�$���IL*�KB��y���bZ��c��ݦ���
S�y�&B�h�XY��Ƌ�sۈ� ����yr����|]�� �h96$�K�yr�� {�(W��o�Tq� T5�y��_��|��َYA�l�׭�y뚃D	j��hƪ l�C"��;�y�+�c����i�$%@����ybd/W�l�kqBX�b�Ԃs�A#�y�-`� �Y�&�6X�\�`�0�y�,�<ad�)�IN
��Y3M��y�e�9>�\�PL��uj�0)sa��y�ȗ�y���
��A���L`����y2� +M]�y��J��
` �$J=�y�aн6��hXa���)�@���y��=����W��:���ϰ�yb�
[yl�1�#�1�(�G�F�y2��Y��h�B��=tf�(f�@��yb,H�Δ�@�"� �� F�0�y�JP��� S�NM�O������y�ĭJh��`�]�D �����y��&��lG�`!��M�l�A(�'�(��qH�/&W u*� \��F���'���J0Cւ ����0��'�����FOTI�f�~s�8
�'c�4³�����AJ!�^�tO��	�'I6|���R�`y���cۜ.�8A�'z�}k�%�x���qu�}�ޔ��'���֪�-=E�����Z�y��%:��� |�0l��U���@��#)�� "OJ$�"�<k~m���C!�V���"O�L!aN=ۛ��j��YAtM9D��Qs$�4��$��H�V�3�9D������UǺQ�f��>^�V�@I#D��I�	�
bxi��nY�gH���?D��Qu/�-U�B1 dـ�X����0D���2�)Z��9d�
�Ex4��V�-D�X�3����m�dN
u��ȥ�)D���#��g���s%��g��@�V�&D�\UΗ8�li��E
�h�#D���!�(0 ���E�3�0 �%D���oz�l	��J�����/D�� �M�+Ea\sqCч]�b��#�"D���	��dW�Li�L�j%a�,D��s�A$y�\H
^�X�t,���+D�ȠU�� �9�i� �nĩQ�(D��AbBJK����H(j'6��� D��(^�O�8�VC�5�"�!`�9D��vMM�"\�S-��&S��p�K+D�!�Z)4Sd|�u	B�C_|Y�3D��"Uo�8/'�!`�aS�v3B�94�0D�ؐ�&ƀ�ԛ0��>�R ��,*D�0a�gP;K� ,�B֢��@�f*D��@P _�3Ej�q���<�m�b�-D�T�NC�'���K��S�,�4a,D�ܓr��pf����҃9���Y!!�d٨
L��C�3Z��]Z#mWq!��S?���
A���w��!T$-Y!�D��T� 
ࣛ�Bĸ�J�JP!�Dx�B)�
�E	��"ɓ�bL!�d��.�h��2Mˈ7F`��Ay�!�Y�i1�TC��_�%��:6�U��!��Y'=�L0����5 Sn���!�G�K�Z�����@��M�o�R�x�'��EI@�J�z�ɣ�	�j�^�
�'��|+�j�dL1�ύ8��8�
�'*�L�Lٗk����<�:��'섔q����56@튋]l�a
�'̎��äC.]���g�_!fT
�'&�m��<_b
dD٧
�5*	�'��HXjZp�T�أȒ�L�ą��'���΀�!��dk�DϲB�&��'��ـ�(�%o�E*�\�6@"h{�'k>�����B�1�7/Yc&��0�'�~pT�<3(vLh�S�Jl:�'a r��E ,)��J�W��"�'<n\��l�l5�gчx�\��'7Z�{��N�)���D��Z��'ĸ�1���0np���	�8Q
�'�jx�1��|�6,�� "$�(��'f����M�"4�ވ��A�o��
�'eH�"��*M�`"'�Z/��Z	�'��$z'������M+�u��'zp0�e\�m^PYb�Z�S7��J�'��u6 � 7&}1rX6Q~�4��'�~�ʗD<:	��Ge�a��'݌�pWbKy!d,���D�@1��'X�5p#�[P6ph��Oڔ:dJ��'"�pū�̠1�*F)2Z�9��'��8�r�AW�1��M%�h� �'�ޝw%�p���A�T����'ń���A��@CBV� �����'�nݡ��'h�C��?~�&�k	��� ��"h�8�9ڂ��n�3d"O ��1�*��ǀ�!H�d�3"O.��q@�W4���QI�%j���qd"O��`��R*4�-�`M0t�ZT:"OH5�v���q����F�&i�d �"O����`��s�U	��ʾ/���G"O��$�O6Tx� ��I|�9�"OJ����7h���c���|�D���"O�@)P�/3�8�Ɗ1�}�0"O�3E�K27}|�9��Y24 ��"O��i�Rϐ���*UA@�"OJ��s!��=��y�4�ƣ,�Ԁ `"O���S�	��OI�d�G"O����44���� $J,�+�"O�@6�G%-EBuYe��^Nt۰"O ��dl�Kij��`Ɛ@I�Q�"O}q6�ñJ��X7m��40"O��H!��-��@ۥ�6ɚ8G"O|�B5O^'D�ʅ� c���\5ҧ"O�]�Q���5b(�0ugW/�LQ��"O�L�M�)3��$�V��7���J�"OX�� ��0`:pZ@�;!�� �"O���B�0idL��G4jIж"O8�k��Xy��4�J�bS8`��"O�����[�����M 8�p"OfI"��!`�h!*P4~A:,��"O<� �7��( ���6)��q�"O�)/|�E�i /`x�"O��c���l���'i'o��}:G"O�aP7�ۺ^:�0��H�1B(�"O�0��?qJ��� _	#�L���"O�]���ٕ7�b�*A@�:i8�E��"O�8�@C(DU�,�������u�"O�Y��'ӗ4� ����>4�:�a"Oxx0׃Ja��p��e[�cL���"O&EI��N>��l1�E�
��"O ��&
�|i���z-(XY�"Oj8*�d���F�	���@�6"Ol�:a1q��h���߳f�{�"Oҝ��B�)�@\���#�0���"O0�0�N	q{\��a]r5x�B�"OjmC�42d3��V�
�]�u"O��Q��
�$�J�P��"����"O���Ȇ�*F��e#���!"O�܋Aꚿ/K��CO�$[J���"O<�F,��!c��R ���(��"O6h�H�
�f���w��8p"O,	j���"8�|'���}��h7"O�`'��)[10���Z�iٲ!�"O��P��7�J!��Ӫ��p�"O|!k �R�ex��B&-������"OJhi��koV�I�,\�p񶘚�"O�LcGjK0D8�K����	�W"O�q��0kXLQ�lEq�*��"O��3e���e��lC�� �v����""O��QLV���A�I��	]*�
�"O�@�M
�qx����\!'�6h�"OV�p��&r�rE���<�f]�"O�Ah�	�0�����E�YĮ��f"O��IG �_����#R�}[@��"O��8u��q&q���һ��-3�"Oqa&��������+�Z�P0"O���G+oez�L?�8T��"O>�SC��đ˂.�Am~՘�"O� �a	AP�4>��B Y,+PNT��"O�j�0J��e��J�yN�PI�"O�����]�A�艐��ُn-$<d"O^�*�Y����vH]1YD�q""O�㒤��Iz6�ȡ�3"��F"Oh�BU�y�� ���ݼh�n���"O�)��EŜce����Kٔ��!��"O>l����K4���Ӫ�Ǥ�w"O�����>�0Y����+XHi�""Oz1��=f���#	�ʭ��!"O��E�i�ƜVW�s��b�"O�c!Q�r�@X��.˾q���r"Ov�S�K�I������'Q��5��"O���eڂf�������?���u"Oʵ����k�������h���6"O|�9n��q�� .���"O���5�¿JenYڢ��
��ᛐ"O"C1N;F,L�����?:����"O�D�Q�
,h%�1ʩ1��z#"O�p��
�~ ��d��X �Qb�"O���g�%x�ݡ��Tda��"O�d���)q8%�D�רE�4�"O�Yq!C7h�6���֊*��q)B"O^��9}��@U�*~d�+G"O 1�)�#٨-Y��D�ac�`pA"O��j�`�l~�P�5!��
?F"O���N�2[6��&�?(��Q"Oj���� �
��%�3�NeT�@Q"O��wL�DEJe-G�I��E�"O��+Ĥ
�������ֳ
�n1C�"O4�p���2y���u�,P�"OāQ��ò}ʂ��$Y��"O���p�Ze8|�ZQ�զr��@xu"O�UC���:0:S�ە7��}e"OX%�Q�(@^��T#Q5 ƺ00"O��17�^�fJ���s��U�(,��"O�܀�iǑ��[��T��vQ�"O��9'	Z�I���K�I	�C����"OP�#��^�-�ziP�)�.�\\�e"O.Ԃ�O��&�j�y"c�F�#�"O�<R��= ��Q�ĭ��u�@"O�|�� �BrT���ohLb�"O.��V�7�x�B��#�L� "OαX&�

[Zl\��1e�P4��"O=��Y�K��9���94B{"O*e8�I��bT��1�	�+�"O�4�`���'�p��R�i F��P"O��%UCD� �6��b�Lɡ"O��!eώ7��]��h�v���B"O>u�#���,����#	[��m�"O �	�I������ȁ�8ڶt[�"O�)�B�yG�]�@E��t�V"O��CL�5>�;%�,@f��P1"O:���
�"E�vA�EQW��1A"O<�:c�@�H��s�՞h�j}�e"O�]��˙�R�\:�A��?k(A4"O��p�04%>dˀ`�"	�0ړ"OpRj��%��L���a"O��2M�&���RG*�?���0�"O��±�	�z��<(A���Q��D"O*Ej�C��:�4�j�B�3e[T��V"Op��G��):^�0;vkD-���3Q"Oj�C�Q7u���I\Z�#�"O�� ��	�$�ʡH�9!�l�s"O� L�3�B�	g�<!��T�d1"O�c!+ ��m#�яc��\kc"O�$�CK�$���µL}j�ۡ"O@}`�L^& h�M��JfAnĘ�"O"}���\=j5f�K`mPp�Lmk0"O���jA�ڴ)�LX�	��\��"O�Q��N#AD�ƌ��b�"OPp��+
�{�a R��w�a�"Od�����*�J�C� J��b"O|�Y�g��z�~@�ע
�z3R��"O&A`��{"v���+^�*\|A�"O�� �_���	+�;n���B�"OH�za/��_Epm
%�G�P��!"O����Y�%��H���+k
TSV"O�rW�1i�<��ň�/�Z��F"O�\��)�(�xQ��I i�@(Rg"OR�R���)f�;E����xg"O�`�S	O�#)�  S�#��ew"O:4� ΂�2��!�$�=S�|�R�"Ol�կV./yL�xE�)"\@�35"O��p(H�f�������~��""O���a��)/��51����x�z)�"O�ū���?����D��)���Bu"O�)9��t������H3��
�"O)H�ʄQ����B�R�W05"O6p2c�.� ��$�
.�ӵ"O����bɺҴX��6��"O�ȹ�ü1��-t����� "O����&e
�L0� m��i�t"O����L�Rs�)�u�X(_���"OH-�b��%pon\K3!�gq(�:s"O�,�3+��X���OU5W�D��"Oj) ��Ԯ��,�P�]]	 ��"O�Q�ܱf�l���.!e�+�"O���D�!q���w�ũP���"O@�
�!�&m��B���"  R�2u"O(% �h�'��i��"�Υ�4"O���@.i<�4	�a��3�8)#"OR k2�C�(R�!"��C�s"O���A�95��kC����D�S�"O��R�ț�>�tK���2�>ș�"O6|!5鐴#gh�G���:��T"O�)�/����}shF�} - �"O�L"�KkL\�6H*��0��"O����Q'g�F�	Gff	��g"O�Y�V��*s,|qh���14g.Y��"O��It�L$Vh�<8��Dn8K�.�y¯�y� �k�DS�q��[�M�>�y��ީl`������N	�E����yr���NX��L�2E���+�
���yR̞6.\��nE�n���Tc܌�yB/<:ԭ:��7f���2d�ش�y�lF�h�^\cdӱ(T��&"�6�yroV�&��BG�#�) 7̭�y̋�p��<r�Jي!�4��Vɰ�y�%�${n�3EB�/f������y��߂l�8��I�(X��k�"̫�y��	޼`)1�ŋ���@g
��yR�F�$��Ic�b�hj@�c�*���y���*s	��ۖA�\�p0ѓ%Y��yR��q <�"��c$aR#��yBE��D�:6��1GD2��bE9�y�C)C�|�`��:7��GmM��y⥖�>��M�%K�6�`!�X��y
� ��#�l��f@0Ǌ�
<�p�S"OL��R Td�	���I�D��"Olx[��D�<�i�ѩJ�5��Ȅ"O����F�1���
�k,���"Ob1��HQ�G�(��,�0q|�*u"O��U�ƲŮ9����!Ȑ|K�"Or���
�-`�
�h7��h�� @"O����W6~��5�iC ? ���"O���II�s��P��Ȋ�z/H�RR"O个� ��(r�$Ip��t+��"O�!�� ��iKыNy|�Ĉ�"OB���(M)<=Ek��v�j�`�"O��RG˛{�P���䊬<\�2�"O$rSÓ�	��y��$�8W���s"O���)��n	�qyfCݳPrp+�"OF�S'M'y���Hw"�49Zjԓ�"OT�u��%��ɷ�ҍY�8K"O�4��LY]�$9���Ͼ(H�\�"OС"�N^�8�J�bL�m� "O`8a��5��4�R�e8�T��"O��!sN֑!�|��	od�	�"O@�L
��Z��bG��ͫT"O��*E';�M��["�d�0"O(i��߳,Nh�C���)�"O������!?����t wI�V��y�퉖D�v�jr�Y�(�����y��:�6��e����Z�&S%�y�
^=aC��� �4l@��W�1�yRb),��T8_�=	t�>o����'<(��_�]~�@h$k$8?���'EPA��M]l4�R�B�z�0�@�'4�q��똲�~�QG��$?�1P	�'+����T�a+$�i�o��p@
�'A�!��@�;0t0�R�&"	��z	�'��`uL
+��)UgL�z�T��	�'�5i�OH��E�_�*�Es
�'P��ja���8t�}��N�l M�
�'�N�	RZ�%{৕"~t"L��'$6��,������f�gD�y�'��U�v�ēu�*�ѡ�

#��:�'�ZMQw��VL�t�f������'G��pP����p&M�!�b�'���A'  ��)!KjI��'�X-:�,��p�ph���_�޹��'ZFX����)�B��Bp��'7@�A5_f�X�P'}����'t@S� ц9ND �d6L�v���&�
�Yg�37rj8y��@M�&��h*�s ����r��<Q22��u5)Cu+ CrT�-�-s�,�ȓ'ϼ�kF�)q�hs!ȝ'U�i�ȓq��YC�	�v�KA�Db��ȓ��\�����EϦq�fH�}�!��68��	`�϶>X.ӓɍbưa�ȓ��lsT#��Ւ�K!񺐇�od�0��E�a�� .*����MJ`�A5�R!��<BC�Ą$��"��F��/Z�����C�Q�Z8��0��d�b�"&e�8�w$��|�^��-}�ԩW�G=u�|�6�r��ȓ%�"`�0�N1�� ��A]D$��@.@hR���y� !�� ��id�<�ȓXz5�e�B0X/$�C�DK�̇�j����îX�e{���0�S��F��S�? >��A�,)訡#���!�`T:"O��ӆR�S��)�W1s�J2#"O�,��c�?�LH�f�K�i�b<��"OpTc@�%��]B$��Sg���"OQ��s5�0Z�ɚ�=���� "O4�kDJ۪g������3r��=(�"O�C� � ހ9IT����1&Ԫ�y�Ӆ_��`�֋��M�z�)Qʇ��y��.
��lI�bN-?���CbZ��y�Iݳ�h��a��
u~��L���y�	�4ok 5)u����xFOȶ�yB��,� ���^ �r�Z�&M��y�΄�+D�-��љu��᛺�y��8�))��q��x
�e]��y��	+��A�_�:�����G��yr�	f}���5Mϛ`-2��d���y\�S��2���"�p�D.�,�y��bd�=�EE�r�=Рf̶�yb�sQH|�e�Z.{����E\��yb�� x*-��p���2��y2�Y�:���u��2=��I��ؤ�y�FQ�6]n@�e��b�N@�H�'0��ZP��B�*p���n���R�'�.0 o�,�8qB� �|΍��'28x"�x~���B� )��r�'*�aB�Ŏ	A�*TA��Ƒ���'����ǫ��U��p0��p��'�& �͈N�X�ڄ��.��٫�'+(�EߞO�ҽR䃉<e>(�	�'%�y`iZf^�`P�	�d�ԀR	�'���@�A�/w�{S��H*(�	�'�4�a���$�V�����0:� �
�'U@��!G<S����b$�0,�p�
�'����"<������D$��'��`+��Z�P��9 �I�t<��'��LTE
��hHP%��Y<;�'�n��l�B %{Y~8��J���y�iJ"���F�r�1R���5�y����X1�#� w�����"���y�m�l0�F+]�<m�\.�
�yBe�9��P����?$�beeL��yb��P�H�G�E�"�#7�R�y��O*���/
�5/�@#��5�y"o͎]�N�z���m�����%�y�B��m}����E
+d��"�@��y�Þ�KH��q�_�U�9y�,F��y��K�^A
T��	<}��@�C��y��K�<��p	�&4�Lq�M�y2HD�j��#Kȹ1݀�6H�yre.+�vhA�V�0�|��E�S�y"F�%��9X�ʕ�6�|hB�*�y�^	H�`�#$^D:K����y2j�1T��@�5��\	="7c��y��ĮE��#�'>P�\\���y�/ĺT�^$ ' �#�LR%�C��yB��tC���0�F_��aS��B��y�`\F!tI��
;\lhӈ��y���P}䩕��Z�BY����y�� 4(K�ӼTˮs �G��y��ۚp	r�:Q^*P �D�go��y
� x��*qo3t�� �(�y�[@�>�H7��,�� 	��y�( ��Y��U�Ġ*����yr�,���23ۊQ�N�i�+�'�y
� lM���Ӯ
���D(��Eh@�1�"O�AQ�&�X��UXn��#gl)x�"OJM��.[�4��kG�"�b�jg"Ov\I�Mƃ�̄����t�~<��"OP$�i�q��D��^�Vq"O\PYªS&<c*!�6�Q:�PQF"O��yH�>P9L`R��L�)tV���"O�a1n���X1겠�B}B%�a"O&�*3�E
lFd�W
�[��d��"O�����!z��vKP�.�R1�"O�h�ݤ�֬ԃ8&XR��"Ov���Ϟ�Qp�yT���}�"O�P�a89�x `��ԡG�#"O��(�.L�07���'�2pmfi��"O�tiƪ�=�f���tE���kZa�<�G��#R��$ȏ�H�
�I�R�<i�E�K*"�h�J�)�9"��XO�<���+"����I�zs�h�'QO�<i�˙��,�M_�9a��#dIU�<��h\�wB� ���F7L^B����T�<yp(�8Yh�����Į/��	��Aw�<!�@�K��zŏG���;���u�<�'Q6X>�d#P(�6(!,��椎n�<	0��R^�9c��(A��Y[%�	O�<q�b�/9F4!#�I�V-�����L�<AS�Ǵp�b쐕BX
���jĦ�o�<�f6Yu����.z8��ca�U�<I��ˢ#P��Y�HH���yr4 @Q�<��
H��5�Pʟ�h����K�<ѶG˼U�x�&²�h@FG�<�&�
��Z��:}�,U��dB�<ID�	c�9"�nJ�j�X%��(�{�<4��R���7�߿| �i�D��t�<1!䔢c�$xb��,�]�g@q�<��q�f�*�ǫ9����w�<Y�L��1�f��F�//��*���]�<q��\�6Zʰx���V\n@:��X�<�6B��e�Z\Y2M�$��˅Q�<p*�Y	P�刋�9��`�3L�<ɢ	�'@��!R�=픡���K�<�K��6�(��(��um�A�<I"��Jp\����{�R��%z�<B� L�	��ϐW��ز��v�<�G��~hA��O
3v��q�k@h�<!ǧ�k^��íNt�na���e�<)���`�4�����7��%�|�<)+]9~D�� �hfw����EM�<9���/�,�3ƕ<���Q-Gd�<�0'&)%�% e��	Vpر@��`�<e!"^�h�(ԠO��f���Y�<q��J
i�uAAAP+%�b��A�}�<�5�t�P,�p��:�� ���z�<!uF�&[#db��a�����w�<)ֆ�L(<�3�`�AKlh�ȁz�<i�Q:��� ��[��� �Dz�<��#�$�`��D�T������y�<�1 \�l�
�scF��;%ʌy�<��ɇ�5'�la@�O�/`�Kq	OO�<�Ь �A����獛KD��t��@�<�r�^>ɣ���(ny��KN~�<�a\�Hk$]��ʻ4�q�f�D�<a�/�+G�|�wiW/���!��}�<#-���i�� ���W`v�<����9�x�;���R� 6�n�<� ~x�v�ŋn|9h��G�5,�{3"OR���S5Z�$�s#�N�K��"O�x����	�bP� ��0�g"O�3C�`1P��s�E�)���A "O��J�GK�o�@ȁ���f]ظ�"ON}q�(+/T�$�TiD�Vk
 sP"O�Q1q��@<J�؁"[!6��Xx�"O��.u�(�65`tlx�"O���A\"?����H�7B���$"O(��ET�����ش��"O�\��N�e�0pi����{���E"OV࢔'Q1�~���fD�9x �"Oڨ�'��Q���!
Y�.�3"O�$��BqHZ@쐘{�Ĝ;�"O�Tx&�M�Z�ΩY3�K�B��ia"O
�p�)ʝb\"����J�"MNHp�"O�Xhlh`�%/h!U"O�-��V�1^�`���	69��"Od��%iH��M�$:D����"OxB�@EL�и0'` �ƕ��(D���աZXP�1C_S�(M�h'D���V.��a�fE$_G�"��$D��
B�@�f	�ͺ%CM�J̨|�r"D��'APq���+I�.
,�d*U
3D��i�錒q�b�1T �	9�n��
&D����K�b`F-H�oR�,�R�9D�H�5M�(�,aA�E�'8,�I�d6D�������)"�ńV8"�c'D��9��tq����#°�&�q�(D� �d�H�!�!�N��ʐF%D�;���:�P��7�- �)��-9D�PK�Hֺq�R�@!͔E��8D�����R�:Ԕra`����8D�ș���
���xԤD n�0@�"�6D�`�%�E'�EA�%�PCQ`6D����a�!���$+��g�H��j3D���&$D���Q�h��L�hQ��+D�0JK��M@2̱�M��zv� �!?D�����vq$Ɛ�s��ڕ)D� 
LZ�� ���M	a�~}�3*OD�jfO:E�J�k�'�t�X�3�"O\UaF��G��L:�G̘0���cC"O(97a��r�*�pg���90�4�"O|�;1&^��U�5�7G�*�"O�Y:�F ����B�H�/{��MҀ"O8���`�/I۬���!o���Ҵ"O�I�h�l��P�)�a	�W"O u�����aHU�p�<	��"O��@Df�!BH��D��?R�<�e"OT�r`��. �a�
�U�8�q�"O�$�p߿3�M,��{PQ�""O�@�w
�h��H�
ۨn̒�"O UI� V�P��#�Ț 4
Ƒ��"O,{4!� 	��\�eǆ8Yڱ3�"O� ��c[-IG������#=rq�Q"Oȸr3����Y8E�@:�"O ܃4�ˈ;R8�KN/F6�AH�"O�X9�NI�$�ǉJ�K��Aa"O�=�mCu�������ބ�"O腊�-ն1��\:�@��y��	Q"O�)�'m�;F��Y� ����	R"O�P���*u� �:����3!b�0f"O~ $�%;�-���3D�`�C"O��x�)(f<Xeb���-۾I��"O� 8��C&&9�����*\�~��e�R"O�� ��L!{��$[$
B0G��$�w"O�l�2�/k��p���*��Q�"O�e� ��:Eb�F%�j��g"O���EK�R!���G��${�Rl�q"O I
0 �4<��!�v�Io�*�H"O\��#A�8����r��3B"Or���g~��cS,E
D�Z�"O0��@g��:f�x��#=
�b�#�"O�����5q���GYd�b�"OJ�$R"G���9�(6R܅Bf"Ov�sES�`�˲AL�w  �+�"OFl:`fW�:�( B�j�C	)Z�"O�)�`i�5&���Ӓ��C���A"O�q�Z1y(�d4*TѺ!"O����m\0A���K���Tit�8�"O����n�(91d�`P�1 �"O�I��.#h���BR:x<�UA�"OZ�@2�?�r��C��+5H���"O$0Csj/n��ݱ7��DR���"O��K�n*% ��S�R,$3"O��"��X�h!�8&.O����J@"O^x�Ć�C-Da�ԭ+-���1"OD 
�mY)5:Y�2<.��)�"O�m�{tM�K�/�,�:�"O��J0�1�9���	ɂ��"OK��g��XTl�4NtT$�l��y�"P]o�l�T�!J6Z)1�NV��y�j
�C��m�Q��H,��E�@��y�#Цep4�mJ(6r��j�!�yBdʪ���'W/Ó+����ybN�55<2��ǀ�;'T0��g��y"�ݷ2�������5%�R<�B���yB�@��4Q�I�3֦��Q`��ybÈ�*3n��Ae۞R8�\�*���y� ��L`��&�E�ZQ�� �yB����qp'��֊��$�D;�yB˄ o����3�Ѓ$Z��y"�� r���3(A��S����y��̮[�Dd�4,4!�D���^�C�o�b���;/�4$�#E��Z[�B�ɰB�=�@#B�j,���4#j�B�I#�{�g_�$4�w	��#�B�	4�L�qt�,A^d���A#GMzB�ɩBg��8�-g�*x{㇑9>!fB��-�����E"'T^@pq!
o0B�ɦBG@q��n�Մ$t�-y��C�ɴ_�$�"�L�~��qbǫ
��C�ɻ~)n�R��!#�E�V&D>�C�IVʎ�1& O�4L���O�$>�C�X$�x��K�O�@��h�0:C�	�K�8e�0l���ݨd*C�	3+�I2gi�'jtH��9�,C�	�!rFa!Ў�A����+�h��B�IT(Hױ0�C��%D�"l�A�,������:����T��%��\+�i��O"�Ñ�I+�A�2p4 �R�"D�ܘ1�O�:e:��+Τءf*,Ot�<	��*V%��el�<^3 m1�RR�<!���W��4�Gς5 �:�A�̞c�	��HOq���2SJ�9���B� ej��"O�ȋfB�1T����%�m^�X���^}b�^@�^�I)2��M�ue��eNPb���o�!�$ʷY�p�:���[1fY"�C_�Qۮ|��'XP�O?�)� ~ �r%�����7G,�X�"O�xaA="���cbXk�.�#E�| =|O�n�h����ܦ������'�f풁�O�]iFAO�����XP����"O���2�	ע	�T���$����I�<���d�,c���ǫ;d�&�Ϲe}�B�IL���4H	m,�A��R���"O�Ql�_.�SA��
������)T�(�卆!Zt")qce�%{B�!ap"Ol�ŋO$mк��f��s�Q��"O��s�5̄- �Z�,�t�[@"O���+���ږ��(����"O��
țl:�]��]R��!R4"OT˂���S�*(��2=궠�"O`,�� Y9Gj��D �d��WOX���B����p�DF�z����g�h�Bቮ|A�����e��� �_26�~��Fy��x2�UZf}��(��fZp�sdB̤�y"��mt�R�
1,�r�R�E��y"��+V$�p�ݵ80����&�0?Q/O�2���O�D̊ C�3�Ȅh�"O�P���;��-���;�@�
��IT�O�d!┦�|6�9pk�m'fy�۴�PxB+�Ur��X� Zp��I�4�yr�|:�y"�_�(�9#kN24v@��a^)�y���!Z��YV�O�v<*��7M����E-LF�|B��:S��ϔ=ݢ�;�����>�R�<	�C?F2���Ą5��[c-�uYaxb�i-�O(Py',�	B� �+�#Q@��'�#<YS���3&�S���H�PM��@t�<�C��s�D���D�a����e/i�'X�?)���Z )O�����^�1�<���<��O��M�B%ZX:7D�8k��l�bږB�a{�O��g8� ��@/?���S�_��ȓ"��e	5R� ��aH��E�|ElZh�'�ў�S�(V��9W!E�k4Fa�bH�r�*C�	�.�cg*׶rL̂��*Rܺ�O�=�}Z����u�T�$��.�B���LX�EyB��/|f��	�뛃�,y��B���'k�{j��f {D/*J�, �0F��<�'��#=�~zuI=Or� ��D�<h	�3ȎM�<qeď4M�X��	՟<��SiEyRY���	e~��/Eƞ��P�X�H����S���� B�	�q,4��D�:=�����ۢ]|!�'A�43��3ˬ9�O)a�A�O>1���I�c��1���]�R�:S�=g�!�$M�0��P1�	�j�x`�nH�*&!���A�(R�(\���(��Y'Lg!����A��8#$�EA�ʃ�&U�Oڣ=��DI�ҁ�1-n��[5��%C
O���P!��FӀ� ���9k�+��Z��OZ���U�5D�*��S�f�~�A�gA,X-���)�Ky�㌑c�T0��,��_���"b+�(�M���s�h���
�er��P�6��R鉕�ȟ���A�:�,7��%��,�Pmy�<�����T��Dj 88|��)E��`X��Ey�ԙ"v-i(���i��D��0=��$C����'D'''$D�geޖ��N�6-r�z�O�xqa�%U���G��/G0��"O��[c&�/�a�������(R0��
^���ð�[[�(	w#W�Hթ�%%���<�qO۱JdX��:H����'Sp(<��4`�&���Inq|��"[�(6T�?a���~bt!�/J;Q �.dhBEM�o�'i.(@&�3� �����QS��Xc�9���r2����'�ӧ��<���ؕxjظ�Ԧ$:h���.�I�[�Q��|r�c��hW0���Anv@5��e�<Q'��xZ �"��f���hLJ�Ic8�$�d%�=���i����RjE+vn�~�V��r��7b�fMh�`6���J!Ok鉙2�Q�aV�I�)�N�gY�C�?����&��If�`�e-�	w���O��=E����*"xH$��Î>�4+E!P���=�{2g��T�R�x煌1�
m��ʣ��kcF���M?I���8�Rb`@��`�L�r�!��O��:�0R�Y�dƇ6�!�Ֆ%�����?Bҙq4�B�!��9��X���7PM)%BA,b;!�$ ]~�Cr�4>��J	|1!�dH;l[���fM�.Nr�97DI.%1OX�=�|b�l�!`�X 9��V�"H��3�VA�'�ax'��%h���ʉiQ�ՃAi ?�O$�=�O��e
�EJ�0��"��v���'y�a�gET�Vv������l>�)��	W�' ����L�0�i3� R![�L�I�'� �yu�B�q��qK%�S�~�1޴��'�ў�'-�$
ҦJ%�L@�% ����	q�b��`�@�V�w��S�`�hL���x��= ��K�'ښi��!��S�Ląȓ /�H���#@��ȫc+.A�(���gyR/�@�@<y3�ײ����^�9��Ȅ�	,��J�YZT-c����S���d?��11�8��Jm��
70&��h��Ɇ!�D-b�(���I3?���	k�IRy����(sgl$sP˛+#���Ve�|���ȓ#Ɲ�1�F�~�ơ����y�"��'�qỌ=��1�&e(VbذB�R��A�!Is~݅�Iv?�d�A:��q&�'q���#X~b@H�MS�{�g�(��+q��3FFX�-��$����$X��Z5�Ve���
�	��PA�ȓ
,���O��&^��7+�#�f�lZ}�����vg̳X����*
�&H��c�i�"�ybE_�zN�Փ�@L=pBj��@)B7��$2�S�O|�1i���-���8%EG%V�̐�'�L3͓<C���cщ�D���O*���b��v/˓�^��hC'3<̲R�*�O��
k|x��iT,� ��Äj�t-��>i���BP)o'�=�@L��^��'�6�)�'&I��j``�r~���Ҩ��w����p�i+���%F�i`Ŷ&� �&����\NA'`�.RJ�����&?,���R��yR�B a��]B�e��X(l,�� �	�y"Hڜ"�E�$��A�,K�K���y��'��MIwG�7,� ӗ��*�yr���%\b�#Z�x:(D�#�Ь�yҥ:;$�;AA�5H�����'͜�y��L6����b�	B��M� I����k~��x���� EIV`Å��cňP!��yR�w���+M?Y�� W��1�O����L��x�C8$���y���*"!򄌐d,R�k��$��$qaL�p!򄗩l.d���I�ay�芛 !�ā1�$����֜x���c�P�S!�D�;;O����f�7xA��� O!�D@ [(ܵ9Wb�fd`�g��I�!�D��A�уEo�x	���tjٰU�!��Q"a���a�%�9Y&�ȹw�A�N�!��;K&����07FD�`j�8�!�� �(1�V?sO�x��O��:��$�"O���!�ٕ	�f�a�Lc��Z"O8���ǖ�8�i��h����e"O$�@$�E���x�f�XݪdJr"O����).f�8�����@8�"Oh���K�3TP9�/�`�@�c�"O����L�7�LI��׍i����"O؀�B�@�g`ix$�O���;#"O����U,B���bDE�Π�g"OL�[�i3�L�f�[�&�1k�"O�ibȉ�k�H���)�X��z�"O�iXslB-�r��3p�}@p"OX�I��uNF�
�ƽY�%�s"Onْ�Z2D�X�'P$s(��q�"O1��k���a�,/Dn�C#"Od�	%���s�RW,� 8k�(
%"On��f@<W�P�Pb`�O�[u"Ox�P#�S�s 0Q7 �\!8�
�"O8qX�&�䣢��&����"OT� �O��F����"=:�"Op�#Q�P7r�Q-ʟC��F"O̘�$Y
d����lF5��t"O�P07B��=Ȩ��J�?�P��"O����c�5��I��$B��D"ORE��N�?L�L�C<$�,4"O��KЊʱ[�R��bA�J�A""OĲ��Z��V89����q�r"O��!dH�?(jH:���@�n���"O��PD`��2�` ��J�3z����"O2L�t�&ؐh1w@ɥ\Z��4"O��31	K?��H���Vި+b"Oܐ �
Q���B	�%V*�k�"O��zI�-m>���	ѽq6L� W"O������܍�Th�S���H#"O�mZ�h��Le����P�1qX:�"O���׃�{`�Ad&>��!Y�"O\�!����+���Ε(r�,�""O�a��zT��_�Sib�2�"O��s^>;b��"%R2}@ T�C"O��,,DDh
�]+ĺ��:!�P�r��Saa[=��q(�!}!�d��&�>�8''�0 @�FM`!�d�p�XU c��?��t)v�!D�!��82R$8�˵L����g�Z��'\�5�D���x�BA�����	�'�����̆-��uač���:}�	�'����ǵ!gJ��BYi�-�	�'�ʵ�$␄4�*�+򌟄	�l��'Tnt�EݵzĤa�q�ä ����'�� {�D�^���B�Aj���c�'��u@!�(�(��LLe�칠�':�P;F��uT���IkyVI�'���q&L3�a �LƝeu�,��'�Ի6���:��\��f�W�F$��'?�X�#�&u~��h%��N���'x	�� �i��ʓ��[Fm�u@>D�hIRȡ���k�Q7hJ�X�e >D��R��\����e?��*'�/D��Km�>)�`Ԡ�`�0]<����+D��K3��:@���6&׫l4�);��(D� v��Y�D��l²���$�9D��c���z�}I��D��H8�1�3D��Ze�Ǝ�YP�*���h��D1D����%�5�P�L��es��	��hO?�� 0�WȂ��8���ۅ"O�c��4I ,���\_�ɋ`�OHI2J>)�U��|ڧ@#5:vE�12 �qEV�<i��}�>1�#�K�`��BF'��<y�������q�`��p����F���B��ٟ��GPbT����^�_�8�GE!?�������O�?<�\KjA 1�q��4�E2��9[�b���D�J�I��4 lAj[��NPP���,\FzB�'�6��R-N��|�Ў�%"�8��'j���ȋ0g�ʩ�f$i،S�}�'�Z�a�j��q��d0�� ���4�8U59UH��v� <�I�9�l��!r��`Љ9v��!�t�����hO�>��a��9\��J�,�V_��YWb"D�Tp%9����h	P�D��)"D�ĀPa�dD����E[<v���5D�p�$O��,;d��7&�qB�4�	o��<�@��R�@]j�b��bH$lµE/$�D��Ø�&���`ʙ
{�^�g���y��.$rU�.�1u/`���	�yb�Y<`�i��_�=�Zyb�֘�y��Wa�c��=�p%����xr�UEx|�p ǃ[��T+��͔C�I�w8�����WfF�ڠ��4?~˓�hOQ> 1ŏO��xA���b�@5OD�=��%�(�8�Ad^�T2�\h��Z�k֡��VC��C��9����A2D��Y''(�ЩvbɽC�I��:D���oI� �6�;��*L��K��9$��Yҋ�+(��2�C��Z�%.��y���$���d��瞐I�/�����'�Q�H�Eǂ
	�ܚ�H� i���`�7��hO����J�#�Ĵ{<(�&肿J��	@��H���`�G�2.�ݚt�]�-V	*�7O����d3�>
�8��g�78�pፖX�C䉕[8F �g�ХT�)��FֿY�˓_��	�Y��i���>`�M�N}J\��7o�ص�FC [�<�� j?�؉�LͨA8�Bq�*��'�Ey��d�PJ�zp�!f\?Ib4L��#Ŵ�y-P�V.�!�`[�A�.�	D	�?���S+O��yBRN��ԍ3`
��]�NԄ�3�<Rh�d8R���mA1ae����VȒ���J�~x�Y�j�Q+���y�:��g�B�!>�x豋�&���o�t(<a7�Ǔ&��l� 'G*s��D&_v�<���^�u���SE��I��{(<��4}圭����{(�Iش ��R�ı���d(lO^��QO�7��3G=W����!�I`X�Ȣv�ic��BpM����[��8D�؛V�?yf%H��6��KW��=�䓣hO�O'M��MR'iPDk� �pn%��'P4<xC.ҏP���Q���oŮ5����0\O�L;E$Hz�n��A�&,��Kq
O�#X�^i��A�@�|��%F����$��yR�ᓏs���k�K^�UʒDq�X�t����(O�˧��,Ky8�KS��R �y�<B䉃y6*���gۋ-g����Cɴ
�=�
ç?���!B)CE����ÅJ"q��>{���rb&� ��wM�6����`�'��P�烨K������=_�ީ"�9�hnZ�J� QR�EY-�NYk�*�`C��# �T	�MS�"P�xǏM�|�
C�=W�x��d��29(�i��4��B�)� ��xA"�^��ph��ҧHj�B��'���?%Ɲ1~�c���~��q�US�<�'O_*v�ʕ ���6��3�N�<1�lĕ@��I�aD3k?rY��̆G�<�V*җF2�l%�F�u&�D-�A�<�MD�hq�Y2"Ůf�FA���Q~�<yc��["\��K,i.~�k"��B�'@axҠؘO��l��'D�R��i!@�ʮ�y��ǹa*92&�	�V�����*N��y�����šRg�7T�Y�mQ��HO���DY�P��=±A��rq�L���M�!��,ww��Ro�Wj�钇@(%���swO���/K�	�@�2��0F���+b�'�qO2X�#T�&�b��J}�)��"O�)�̜�0M�H�� �/sB<��S"OT�r���.u2�u �4K,�
0"O9U
�u��u
g)�n:�a�"O���ҀڈA1$}x��k���Q"O~$���H%3C�``hV�>q
�$�������B��g΀"B�Fxr�	�?��'���ʠ�5I�%4��/N��'4$��c�:i��jN؊gQR�'����9OZ	5AP�F�Zt!��k3����"OdlH���}m��P�(+�pɔ�	]���I�`dp�`*I�E�$�@hфC䉕A��$c���+ho�E��.�|�p��$�Iv�����#n ��
��^2�((7�ǁ5�!򄆍L\��dʪQ2qذ�)�!��x�h�Vh�h_.l��O�>�!��Ry��|�b�SYD��3 e�)�!����YH��Xo^�c*����mV��!�DP����)���Vr ��f�ڿ�!��*,���"onp��e�!�d0{�t=�`��5R�D1�mG<�!�$�,�l*��W�3���W-�!�䛠|����E痱��`T-׆0��D}Ӕه(��J�`*��]N��ؙ�^���ɠwo*`��a�5U[�4���%)~B�I0?N����L��(3�d�@ C��!(�Z��DǕ��&<p�J��Ot�B�'E2*u��
0 ��Y����$��B�ɰ�(*5k6M ��էG�P\�B�ɇ�`�D�O�OOƉ¡��r��B䉭C������8g&��@ ��unC䉛rg���Bo��C��ț���"(���>	�#]�#�ؘb�1�#�
IU��l�'�@�,�<I��JE�sH�XҊy��'�jd0�+�@;*���I�*x>�I�O��G{J~B�_���j���4�����e��yۮ1�ȓ���'�FA)\�ag�9;D�A%� ��ɡC2�X�4�������e�����$-}b��Z�F-�@#ީ)�6��Ҫ��yr斋���q"�)#���3i�hO����e��a��.�V��7o�9�!�d'P|>`ǬH�}��B��"3+���)���� �&����f�	[!�#D���dAo����rk�=Eq� ��'D�����k�L{���E8c�7�O�'�!�T�2��тVh�;T~D`�'��{� ��>�
UγIM�|��'�8��NB� р�6BG�<�𐓘'��"&��:�0<b��[Y����һ�y�*MMz�]Ұ��2
�h��j��y"$�2f���f^�W2�� ���y
� ��D�
	F�xX�L�l��	�"O�IK;VL�V&�ܙ��"Or���T�����uc�)���x$"O��y��ǰ8����P<S�rt"O:��w�l3
�[�i�	��F"O�����T���E(��z����V"O��� �Al��)uf���>��"O��� �*s�F���gA�0�	0`"O�%�CgߟI�*}@w�@�b�h�"O�"A�x%V�Ѐ%˚(�^���"O�XA�ME�\�Tubճ� )��"O&ec��� YC�c�w��D�U"O$h�o�P ��ƚq�X5 �"OZ���+��,�D�
�g@3{����"O��!��,*�(����/٘|��"O��#b�<,Q��A+5j+r��q"O^��u�(3>n�D<(���i "O�a 'T�.ᴭ�ԡ��}sP"O������ZĘ�挳U�B�Z`"O��@�ڠP�ZW � ���b "O���q�\*\�xۡ�[6�,T2e"O>7oY�J#| X N�BFn#�"O6��U�C7'���4�L*��"OLx� �ǋ<����4+ @5q "O�pG�(�
��N����"OhHRR���U��d
���#��@a�"O�����/vBf�86΀)u����P"Or�A ӟPf����lόU\	�d"O����ȶ��U��նF�2�1�"O`���	,F��É�=`�j��"O܈���QY8��2�A'
��%X�/L�k���5`)���d�uT$e�"ٺ8��lP9#�!�Ă�C�z%)oO.p����B�V ze!�d����南f�n�t*�'o!򤀐0�*l��g���p%c�a�!�����0��D?ex����
�!��_JtV�I�F��)S�X8@�!�� ���2.�Q@ZP`'�B29l!�U�������O:Ӕ��E!�d�;j� )���+Lݺ�ʉ5J!�
�J�P��p-�?9����Q��:2W!�dW.W���T��
�8��D�đ��'�8��gC !s���4�����'�Da�Ճ�p�l�T�.���'VF��vj����!BD)H��A�<�P��Qz�Bcҥl�$�8�J�~�<�V����y�B^�A�ƙ@��@�<Iu��jD�i������I�U�<Ir+V"o�!rB.˭`�>@����L�<�g�� �VH& \�p8�#%�N�<aD!L8lNM�K�C�:<ز��Q�<�`�%#�C�Pr,��wUu�<�D�)g��1Kt��#�|�т�T[�<���<Y ���W��bȹ��]T�<كFL�p{�u
�9�1�6�W�<���*$��+��ŖI��*��M�<���ŝ-��4���)EC4�	�mVE�<�v��qn�B���.(�4�'�T�<A����Đc��6s5攲�B�V�<Y�aS>4���cJц�:c�n�<�R�OF'��Q� K���e�k�<yQ���_���BbE""���i���e�<��N��nuf4�o�
�mk��K�<a����k/�B��-Ī��s��O�<� ��ԯөW��$!�a\6� t3�"OP���dN�~=�N��p$��"Op9�B��$M�N�jԅ¼[�TA"O��t��Zn���ER}�����'�de;���hD���5�'e,�Y#ZW B�	Xk�����:hHe�RD��� �>��ُ��"|җ�A�$���@�.v����\�<ar#�a➁X�`�y+��P@"T?	�L4�➢}�NL�mԪ �e���dL�&��O�<��σv3�\&-�
�sǥ�p���8IUH	rӓ���rhͱ���El���v���	9^/ �zV��h���ywnƺZ4�ӑ&HLs!�d�,K��!�0�I;m�Q��lKQ����+�!>q ������Œ���Z�l����*D�D��P'Ƞ��I�RU��ʦ>qp�E���H�~���c��/���R�鉼G�XT��"O@�)���4�e���N�	#@i��"OHt��/�8?#�|�s&�M�p��q"OܽӧBB5�^Q�B�R�t=S"O��8D*H�r�~��Ҧ_�n���"O���@c�� W<�:�A�,%"�"O���#cG�`ю��)F�LI��"OLUx(��q�t�K\�J4 �`�"OԐ�Ec�=)�ց�Q��5Jj�V"O��	�fF�}�p��h�,U���"Op<�
��>���gJ�2
�:�"O�̓�J9�*52U�8)����"O�����JCdDXN�co"|
'�'8���'�`|����7h�:=�"�7q#6	��'��u�B'�=xv���H4i8^M0����*d��ę��i�$q��uib'�,39r��֋��!�ޠ'�(i��ێj���0�*xB"����=E�t"S�U�8��GJO�@yz�)WE��=e!�$T�XG���?}��Sd\%Oq�I��Q�����=��'P�J����5lч6�$���]x�(�%���}�lǲ�b��y�~H@�e��O�d3UEX娟flA�(�	8�`�Y$p�D��s�I9\�!bR�ӭCK6����&s��Ҕ��=������]�2Hx��+�~���x����8� MY�旈3e�b�G{���SlPT�S�O���K�	Ϳv5�)���)k�:�3�4x�:���N��'�����p<q4aO!Z���C@�_r�R`��[؞@��k�X �hPÈBG=TA! �q�Vy�2�BI��r��dH<��Q�܄��W�]= ��pjR K\����	!F'S�]�xʒ�W�k����cq<=�%:�P8�q	�m�����
�2���'� �j��Ƥ~Q�����>�4��S"G��dʇ��	���s �]6��'R������?��>�$J�a��EiO#^t�9�@H�'c�Py�Ì�x� �Y��@/2�L��uEl��I�2j�ybLvn��oZ � I�L�:M̜Q�nM\X��s`��z����	o\}ST7O������w���w�T5@}��c(�*�q^R��!ׯ��jH�z�	0C3�lq�GӖ.�Ѱ�O��(S(Y13$��)��G�-2�i��4��#Sb�q2b4����&%Έ sY�3&��F�+8�u� 2B�+��z�#�92��{��'m�!���!Y�d��pdɌW�n 0!f�04il%ʷ�G<N�� �i�g�c��V"|�vЫ��ȏR�d(8)���^�TS���)��%�xp8��O�I��ԃ�*��9<6�D���A���?��B��t�bQ�/;��!��/.�<%P1�-���3�<&��3�9[x(0!�� U� �9)�w"�d��) �I�6�4=+��H:^p 8���K�iP�
�3ў]�!G�f2�8$1�x5����l$`ia��3u�P|x�D�6�0ř��<Kg��S0Txӌr>a ���r�H|%�>���tj@��m� q�,��c�d����q��7z8��&�Yl�&� �S,D��<0���9h}�Ř�mCR�(�:ti�a���4y�M~"B�X����#2�ꩉ�J b�'EF���W���f�?1vPXT�OZ8�Qo١k�A�����m�l хS����1� ����ą)H����$B�\~����k��(HD6L�U�P�0��� �(K��?�%��\v�=�gCQf��ڕ�I�)�Α��']�~4�~��:="�)"�h 2��0�\0p����C�#3�lp�P(�5c�O#�=�( 4��O� j�y���A�a��\�lA��"1�'�d�ȕ�̸;�z Q���',҈�2Ŝ�$׈�H���PpH\j��͸*W�mhR�8��M�(R�O�R���ɐ�� ��Ӿ,� ��dV()���IHY�#�a ���$�\��+Įi��I��E�l㞠Y�bQ�����L��pQ[���
1k��U6��� C%���/�h`CZ<N��D�ư�@!S!��J�:E 1o��ybI�<��D[��-C"�� �E>$�8e�s�	�U�T���B8tR�sʟ� oV�S��4�N%3q�,�5�&�Ov��ѨS�[��KC�ap�D'T�-�А�O 95<X0&'�O6cE�U&j ��ҧĽv�����I+3�6]`nX�<!�+�P>�Z��P0�z5�r"˩i+J���y��Z,x0�Y�b޸�j�0�����<q5�݊A���Q�a�4�E�N���"��o���pe��y�G�s�F4!�C6P�����"}x�p�G�~�g��@]*�d�3	P�0��ݛe��;G7!�D�J#�т��:5��!�l�",
!�d 58�PR!ۙh�v����!�!��[������غ-62	��O\�/�!�d�v~�0�E� }^����7e�!�$�/*�|(8 #�G4<0wN2�!�U���*�|�j���.��O�!��_����B�R"���Hu��i�!�d�4w����<D7�����'<�!򤈵-���Zӌ�5^�g��,�!��1q?�����_�>�Y3�"�!��(ܴ]�B�����wN^�!��M�duy�剈khy9 -&G�!�'	=p��K�*:\(R��s�!�1M������
����M�6r�!�D�Bn怛��#�
����Z'r�!��C&鈩c��V�����W=�!��ӭx0\k�n�p|�L�@G.��'��0���Nx�X®۴����2	�(�8=�C�2�O��4�H�ld�H)�eW�{/�� �֬Gh�y+dF/$��ȕiV�5p,pk��w�
�Hэ1��8�r��$l`�>)a�陔9ܞ@��I�.L����I8D���B���W�Û���di{�0o
t(�yQ�>E�TbUV�� ��OA`��1�Q��y�N��C�I_�;	V��������D�?q}
��Q�ς�p<Ad��&H�X堖L6�$[EJ\q���
U��\�:H���R�(��]��Rl�bq���L5+Y��P�a}�l���2q�v�Y�`�3 ��C��+�mi�霖�6�*�EG/X�`H1���s�!��9;��Y���1(�Ȕ4�A�>�$���\9�"HL��)�'t��L���hl!q��WZ@��)Y�9{g�/h,�]�"�!�I�'�\D���LA-&P��I(Z�ģ�9==�4�
Ͼ-]���D�9�bUH���hv�����T��UO�d#`�W�#������V;)ziy��I2���e��	5`z��VJ2W
R�V`�9/��Od*�e���ȟ�%k .�*C8b<F�^4и"Oz �d����5x���A��%+ǁ K��I>�>��g�2}E�4wFG�Bs^u3��|�<)��O��<�CP*�GR�b��ނ"z� ��-�<�F��ɰ	.]
ge�-t��1�)>pA���D�upMZ�\�y�/��\����[�����ϒ��y"N��!~X�!�f\x̸l��=��'^<U	Ft]�E����
,�t{E��#�<���)[��yB��C�h�2$�/�J�:�N[N�[$o�-��	6$�Q>˓I�V�	�`)B]S�F��݅ȓ]9�E�[�'��4;��^+uص��^X�5)b+�s���LQ�?�f�(R���P!Ve) �2\O��biՊPQP��'�$y�R
��c�i�$E��@��'>~�AD�0w��)Z!�ͩ�C
z�����Q�]l#~� �Ç�[�����"]s���"O�ePt,�>R��띮y�8�Z��G�ژ�K>Q��>QajT���A&d��f��\�T�<�q�P�Z�����58v\�4/�����@ܙ�a}"���9t�%�S���S���r䚸�y�X�_� 	3

(d(�Y+�P:�yB��y#gQ�_�*����|�<q$�jo�e�ï6����n�<ɕ(�i
<���N[l	�`ɳ��d�<�&½3���-N!Y�D��͜X�<Q"X���@��h�i�` GP�<�����X�hT� ;\8�c�T�<9I�(R+�W��Lsѧ�Q�<YS@Ǧ�|�g�@�~� Y����H�<q"(�nb�q��W�7�P�Ұ�JK�<��h"��P���Ђ-Z��@�<�1'ªd��]�Ĭ��8�A�#�~�<�'��H�\9��O<N�����@�<ɂlS�d�9�΁YH�%�A�C�<A��M��1k`a݆!$�mH�@Sk�<9��&k����F G:t��8�dM�O�<�g��T��F�0u��C&�K�<!s+��_7jћ��۳�u��@�<�-yذ��b\*b�be���W�<�`B^V�|�.���SB�R�<9".O/3`��r� "[�H���I�<����'~�yc�dZDs��*B�<Q3��6�Z�isI�~�|3$�C�<����8]Z���f��{�li��N~�<� @��])q�
٦sԉ�eZv�<��-
5�Mq���Cx�P���s�<�˄�|)P��Ւl�����G�a�<1v�ɮ	J�#�O�n2zq��D�_�<�CƐ�ox`p�+_<I��bb��|�<��T�J:�i��i��<��{�+^y�<)�b׮b"��j@A˃P��Y�&(m�<ل˞($�����L�X*D�B�[A�<)B�C-f��JV!tDp�Dq�<Y� �6��m���|j97��n�<9b�zO���� �H�l�m�<�DIX-A\V��a�hA|��G�F�<	7��o�Ҽ۳C^�Q�u�#C�<�7Aפw����@�0h��Pzn�}�<y�.xظ��l� x�)2��y�<I�m�-0�3D&Ƅ��,b���l�<��̺/1���4�Â�J9 ��o�<�AEF9xtn��RGP�T�8�Q���q�<�F���v�h@c_��"5�0�St�<��M0M��G͏/l��͸t�i�<�)�-9�6츀�'A�Qpt�Z�<ys��z�ꒃ�9/�yp E@N�<�T��P+a�g�tRW��H�<�q/J&����+��Y���a�EX�<-|��"�V:�h�V��O~bP��Y�|��h�n�X)"��2�ZH���>9j�Z-���U.P�vxЄ��YP֠2V� ��)
�A���؆ȓ:�@�p,�G�P�ň���*9��m�ª�Dfdq��[�I�Z�ȓ  }��JҶf.g`Z���P�W�%&ez2MŋW��A�ȓ��Z�%$�`�2Eh�t����ȓU&�-҃�Ѥx<Z�ZR��È���!O>�F�@Y��!��w�4H��S�? �q�$O�8�2�2�gJ�yʍa�"O�`�7eC=AU(��,�1����t"O���,W�zX.Q��2�4a�'"OX" �4�z�k� T��,�"O��0��L�|�Z���I�I�@M3B"O�yѦ����9Ƈ���|�y�"O�*�l�q%��j6fȝ'�)��"O�A����i[$eީb>Z��0"OZ1Z��K;1���0e+�W��Y �"O:(���>Ÿ@��J��S��({g"O�y�cfX (�hY�G�{p�1Bc"Od�����=c�@,���^�vp;�"O�h6|l�2F��Dmu�w"OH��ȵ@��x��8_@�Z"O�0b�e{�Rp7)�Q;$"�*O�P`���3B >g��@�'
j�;�0|I�pG�(^��9a�'�~s��Q���'��R*�]q�'����AM�L�ļ�g?�䜨�'f�}J�E�dYX ���,����'�&��d :~���A����]P�'����)^�Y�X�ڱ��'��a0	�'Z��`o�=`�8��)�2�:��'���	�%єa�-R�(�Oj�H�'~Q��ۆh$���G0��m[�'z���EߑxR���@�n���'9X��4Ò'<p8��<G�$�'	~�C���}&��paL)lXe��'~H@#$ڞz��E�I�����'�(��7?\����+�
]���j�'�����E�5{@yz熖R����'�xi���P���ȃˉ)[��J�'}�9����	ي-[cƗ\��8 	�'���Z�p���o̬X{����'��5N[���kr K;H�be��'�Z��@.M��AR�KXh�'v�p���;'��1�@�1�ܥ
�'��R[7<'>(S`d#5��#�'���RឲCv|x���S�����'��:��7&��2���!IB�
����\��;��遱/�"}��&v������B.G�!���������tK�W*(f� ��@:qY�'g�>�����0��'5���BCDp{�C�1��d��8�p�I��}m�7m��[��p�wǕ���=�P����U�3枠K�0��&�x؞�3��#��|0�'/�\ ��F8=W\ȃ�D<�~�`
�'�
���=�0�Qt�׏��)/��Ak�D��u`a�<5�E[E-}�c�|f�7Z V��c�0u<L��΅>I����ϒv�bxf�O/�LJ7�F�S�n�����Vd�d�N$tcn�-���)�IK����J�b�K�� J��-{ ���$�_KR��Y_N��!<b�Ӫj��X���d�P��caR)H�x7M�6�8�s5�W��=�gg��U1٩5��
1�=�H
�<IUÑ�_��x�P�ޡ����''�|�#AB�|���*��HxؕA�_h}҃a��=`L�A�"O:��uE�mn�����a�!�R(��\]���Ѧ/�f�ӑ�߲/�4��Ueɍon��PN�k�5��8�b`�]�G4|5
 c�R��` ��'G:���+�m��d
�\wZ�q �ذS�z���a_&A�H�'�'�����;�q�@��YpP���~��)�̹H#�+r�&d�Ǧ�0͈O����Ŝ:cj(J�߇J��� �Ox �z7&1��Y�Ư��e��D��G�wb�s�H�%n��jFꏕ�����M��Hf)�=��< piL�8��d��g��h�sl��Ҝ��ș�(��Y� ͇]���3�nآ����I�>�T�u��<�p?a�δ#�\�とd�vq�Dݕ7�Tbꅱ8�rf��6IV�Eͧ"�R0�AÀ�d�|�'H$Ŋ�R	2�&���n�`c��4�O�%���J�B�A�e'vזX��e9��M�/^��0��#�kO�ܡB��ؠ�'Քb?-9L�1�ܝ�G��8A�6��ǋ4�%Ŋ��A:1��u�V���� ���3!܄N0���&B^%ao�=J0lK��	<H��TT 9�3�I$o9��C��@Z�KI��[�6扻3�X�{���6��S�O�����"�qP\�w�N�
�uj�͘$�)�q�Eu���"�!Iq��%�.]��qj>?����<[��-(g����w�Y<LP�͢��>97���8����!�}k���V��<s%%�:9<��SGڏTh��{�E��Cڂ�"����=w���/��V�TA�)���g��2�`Z���@�Ç6�(#>��ZjdS� 4�><�<��L�Y�����@��P���=A ��
)~���'RD[��Q����QV�7"p���'(�9�	�aCby�O?��p(ʊ���"�BI@B�ڄ�y��~n��)�VFruC������8�����j�(�p<GK�I�'e������p��pe��w(0t�>*��Ҡe�&s��9P��BH<���ˬy�^�3�	��t�)�*�i�']b�;�B�Y�'z �ْ�[4��9k�L���ȓ�p������0�0�׎��#}H��ȓu�xD��'3H��k��@�m���"Qv���]��30��)r=�̇�'�	��'�lJ�\�1n* |8�ȓ���Y�ȃ�z4^���&��x���ȓr�p�e�K����rGƨ'�FȇȓJ<X� Eԇ^q���@�ʂ3NE��X��m{��=��UҤQ>L�jX�ȓk|=j �]!Se�š%��9h��9�ȓ$F��ƭ	�}ȅW&��Xa�ȓ~�����oT�F�Q�(a�ȓ}��i�$�'��lK%�ǈ`��� �DĢMơu2��I��L����qׂ���^Y�P�P��lL�ȓ �f�K���y���U��"a�Յȓc�����+�v���:��V-��y�)�YܸQ��[j����"&�y�S6o�i�u�*"H���E���y2.�?F�ژ�Ff_�k&�k5 ޴�y�`T�`��U���N�g�^a8����y���/2����E�!S�iD(M%�ē&@�t#�0<O���� ;�T( �H�gJ�8��'8��82�L�bn�"�O=1W9�e�>�6=;�O�����&L��)t�	.B(���	�z��H��];d�q��Kf�6 6k�M�d&�呶"O��kҫ��{m����=Y4�[@1ONi�W��:�t��M�"~eh�0/5D<��gQ���D�ĭ�@�<Q�/B��iD��5�VM(�ǏA~�(�n.�� �_8�`��̓CVp�iSlJ?m^�Y�"5�Oиp1���Ae.�X�CZ�,�(i)�e��6t���	B��Px2 }h��������p���O���9;�$@��4A��I%䘛0Z/v�[��#�yb	;�tyV.:��زR�J��y���e/���#Om��
�^Q��g���ܘ ˙��C��k���Ȍ�M��H8En˃sb�s�(y� j\�:���ލ z�hu-��k>���W゛%��~�&� y2�FaӻT�vԣB�W�|V�x{�O�`!�$ߩ�
uq���
A�����j�pg��p�v�3u6����7Hїv�:(�A=���s����st���IM��X��Z�6�v}��h	!�BmhcU
 O������#� �h�������>�7��P���;U/���DJ8@����1�|��p�-X����4��7�/q`M�e�\��0>Q��Ė9���!$�ζrv��ST�@����ӭ+���0OtUZ��;rff8���[�+�6Y��"O��@�J^"[N4��!lȢQiu��P�g۰��LFՈ�:]#U��"  (	sFи<��H �"Ore;w$*J�2XX��Y [����bV5tKv��t�> E%�gyr��)Ж�q1뎨�V���R��y
� %0@&�\]�����+}���тc�x�%ހX)a|"KZm2~�@�a0�Xh�Cj��p=I���(�����g�t��GJz�*l�`E�;0 �#.?D��3�
x}����AJ���j#8rpH�)t,�qW?��gݫ1�-r��ȺD���g�8D�Q��S)�8�1D˚��X����7�6e�"�|�M �g}�l��w;%R��>'y�%qH��y"L]>I�8� n�]��bA�G��?���C-���$�-8c�=q2��4B�v�e@ήI!�D�&i��#KP�����Oߗ]�!�Y�sL�a�� !{m,|!�]�o{!�D��-�� ꗆ!X�ĮS�^f!���Ea�dف�Җhz��Y��U�	<!�R�
��e2�>H���B'�!���u�����u1���#jk�,C�I+b�P��D݁YӲ�w
S�C�	�7�HX�`��=7�Hs�3Z�B�I8"����7ǃ
��#`Iخ
B�!hb\-�$���SײQ��ؘi��C�ɊHB����HįJ�d�`��B�IW����D� h��蟧p= C�	�hy^���G�R��`.� J"�B�I�m�Zi
R̃�6F,9�Rn��'��C�������7~#���wʅ�OB�C�	�y�8�I��X��aᣟ�k��C�ɄKYř��@}��KC��*
ښC�IWP	��fA:H� �'	ە%RC�I�f��(��)[k��i	d UuW�B�	1K"���Y�H�������<��B�	�;�R(��L8M��#��+g�B�	,!:���ge 5k���V��s��C��Q䢅Y'�ƃ��C�Ӭ��C�I� ��%'[�2|�Q�GT#H�!�䛟ne��Ǥg�I��+�!�@�<H���Gpx�f�%�!��	*��Sg��H�$a��S� p!�ۺ0��0���BM: �!-Y.�!��,̢a'�+uM�Y���T*w!�$�%]#�(֡ˋ"����+�-p�n`�բ��e��(���>�d#S-^(� ���O�,���*G�<�y�V�]�@(�ա�o�ǣ��D�h��Ig32�k�����M�.a�&$x&�>I�ȕ8l�t�çH�*5hY�K	�k� [6E5� ��OPXB� ذ-��$1��	8�,�s�1S�o����0�'�Pe" g^�U���C��>E��$V;m]X����-(�0U�3K`�	:h�LԊ�Q����6.���ݶA���ʃZxI�O�/Pzet1O�8`����_���:��C����R�bEj��6-1�(O�?Q�W�N c:�����L�5m��#BCGu�'5v��)�ԥZ�ߺNb���fR�k3�O�݊�y���޻! @��Tk�pl�y#�Iæ0����kÜ>*���>5C�E�  ��^Z �}�P�<��)�'���
�Ǎ:����ލ)+����hO?����Q�]����k�v$�)Ҙ�HOa�I�U�A�瀍XT|@�6�U��A}"�5��)�5j��
0jߦ�N�����qO��	(ԸO��'
iR�'���8��o*b�d9�O��͓T���p����+��D�(�eI6;0ȑ��٭c�M���O�u�<�l�O�>�A�f']�J8�g∣w�씡퍜4i����S�O:@�Ӣ._>���̎8<I��'��'��)�'[����'K�0�M�XM(��'@"<�)ʧFZ�	�e��TT���fO �Ρ�	ޟ�B�}��i��U�"��3�̈́�y5�ąu��,�	]��W���A¢~�D��+5�[P�ǧ,�f-��@&�	9txx¢o�2k�b\��S�X��[c�уq�L��r�W�Z���D;�y2�.�~��eh,�F-����^��p��?��XC�"O� �,�)�	�b��	�^��"O��)"K�)�� �ˏ�p��l#"Onx��iY�7Vh�!d*�qd4�S�"OT-* �R�8��� ��ÖAV	2�"O�0�Go )�.�	�-�%צ��w"O�M*�BI��-e�-|֌�ZT"O�mޡ>�Ԝ�p��0a@"O�q�HR �XG�5v�Q��"O�Pc6ɉ=��2�BO���!�"O���ʇ�s���W���B�9� "OJAA#(�m�A��"Fd]:�"O����!h���I��S5C��S"O��8��Ǚl�*"�P�-ʾq#`"O|]�cb]H]h�qG��:�~�J�"O�i���]H8�E�W��L��"O� �$�-D\P����Q�EX��"O������n�����1t��*3"O����,��#���.�.� �"O���iY�p�I�A�	#�\@0�"O��"��Ԡ|�}i��׭n�^�z�"O �yTLј=�F� ��<M�:5�p"O�+����L���7{�0�ȅ"O%����0=e��0�Ut����"Ox  �OP�g��M�ԡο[����"O<8c��ۏ���ډR�x�9"O�Ġ���EHh��M#�"�"Of)j�iO0(,�4
� u}��{�"OZ�gY�bd�x#�����P�!�d��`��ɠB�[�Cb��a�\�v�!�D�(C�բ�O�$��h�M�%�!�D�1_�@�9��	B �0��Bx!�F�/`0U�re��Z�jA��
C!�K�,1bl��o%�^()�-WN�!��D>h�K$��.C����G�i�!򤕤�AŐ�T��,�A��\�!�d˛>�� �Ҧ�����@���!��G�	9��2���E�@$f	!�D��dے� �\pH�۶�N8Y�!�B&}݈̀�
�u~��a�$��!�DY���v	XWb M���ۆ5�!�%Q��`�& �VUj=�����!��	�qj l��%5�0E�D�}~!��Qwt<�����)�lEL`!��QbF�p�[���0!&*!򤐫_�Pjt 0W��9�D�'!�D�=o�
�Z��M	��PV*\!�M�̡%
�D���qOճEQ!��Ց0��<�F��p�bi��.�.]�!��N�< ����c��5hj�!���1!�d���\�Bt+�VZ��������PC� b �w�����H��y�
�O��ЃDΜ�b�:=2q����ybk090
�{��	x`@)ab� �yR��P`�Ia���~(FI�w@ �yjǨD~@��Ou���8FCӕ�yr#µi��ܡ��I�?���%d���y��Կ1��*�JL�8.
q�U��#�yRi� qF t�f	0$�\��7�y��8nPA�`�4tl8EG�+�y򧐖���jQ�8%�D��䮈��y/ �x$��c|a�k�8KN�)��',�t�p퐤ܮ�z��M51h:��'�h|�@�z]����t�ȫ�'S�Iy�LF#s�����+G,6�ލK��� FD�R G�7�$BPFO�Z}��	"Ov��G�\հ�H�"��@�c"O���wN�iB�Z O��;�L��"O���&�"dxh��C�҈��iH�"O
Q����@:8\�����}1�"OD�	�K�]��=���-u�5�"O|����J<H���k͐a����"O���4J�}Dz`��*�>x��k�"O0�h���C�P�$`͡2a����"O�$� �ݥ;I�Ub��D��J�[�"O8�H�
F*N�`��o~*8�IV"O��8�cZ,P��j�-\:~�`h�"O� �"D=`PlI��Qq�����"O>�iLZ�Z�ȩ ���S��9c"O�x	�
��Z��kc��<`n  9�"O���kߎ&����\6_���"O�9��T�x2��-UM,dj""O��J�.���A�2B�+ۘ���"O|-9ĬӚt�@�Ap��<Y�*�"O�Ys��:�c�V�.U���"Ox(���:a^F��%;"��t"ON"�ɖ�'�J0����-�u9�"Ov Ƞ�ޗG�p��M\�.�d�P�"O.��M�&/�zЧ��6���hW"O&E��䉠[��x�j�h����"O���nW�TQ2�/H�E�Ȉr�"O1��,>n:�"�+����"O85:e��3#glŹ����j����"O�<iS��$"m*��Ԏ��K�P��6"O����M9C��Dr�m_"qO�I�F"O�ȫV�OT��!R�~Bf1�R"O(HU.��ٓvJ�o>�&!�DC��q�'ڢp<�Pꒂ��!��S�t ➖n1`���bY#^!�1a)`�',շ*G*�;�&?�!��?�B�@��F�}[<� F;o�!�dQbU`��t�
"k>L�X��#C�!�D3r�^ �F�5 4%�dl� �!��[��.���I�@���h���_�!�H:6���e	Pd�"I�!�$��{�ڔ�0��� �p�C�v]!�DXk�,��ĠG:tu��ņ�#K!���F �$�4!PPl�  V{!�V�pi�t(���|��L�a���B�!�d�z����'.����.R.�!�D�0/Y�qC��q�F�����~!��'%�)g��g�p����ō%j!��y�.t�MT�G��,YUkC�5!�d�(<&8�RN�-@�����7+�!�d�
FH*��$�aA* 1GÌ�!�P~���  n� �)w�G -�!�	/$3�I��<#(B�!��'N!�d�)x��Y��yb(�k%A��!�Ձa@ hp�%?/�L���+c�!�օQ�pҐ**(f�C��ݹt}!�G.��wI��-���R�ɤ>�!��6��=)Ҡ��e��`'� !��D'q��}R��B"4�t	:�CI-1�!�䔛~�@�[UaX�Z��#h�)�!��~H>QI�Ǜ�/G��(� �*�!��Йd��=�@�C�)�lF%I�!��ȳ	�y�!��:^�;�˅-�!�ۋ9I��#WlD����+A�!�D���y�V��DVV�z��]�{n!�� �p��G	.g�}�e��.$�*�"O��R�a��]GlJ1E0a!�ջ�"O �#�M@���3Ab�=� !�"O�0JQ�3K��H� � <�XIhF"O�t�����h"yI��)~�1:�"O��(�+Ür���ښP61�"O`���h
�Vh2	���5N�e��"O>)�$�[���e��-�!6��EK�"O�M����K�(�H��c��m�"Oh;ED�<H��׮R�l��"O��A&/ԧM�0H[��[ :��E1e"O2���Ƃ&)QA�ڄ0>�|�`"O�� 6f�/*�6	3�5K���J"O}[W��`���f�f���x�"O��X��A3��\�p׏m`��"O����'��f�|�YË�S�^X��"O�R"�s�Z�iה���h�"O2���iE51�.�I�'U�	�N �"O�l:� h ���᎞5�ɣ5"O��s3�LY�lT���K��I��"O`��M "+VΝ0c��
=uHiI�"OL�X��/�0�Ӆ�]J���"O8h���_�v��(��썖x�H��"O�;�-Ƶ����.=G�2��C*O>��&��1k�%���0?��Ы
�'��x�$K�"�N�	�e�ܤ�	�'j^dE�
;}#@��qjfZ켪	�'n�a�!�W>9z�i¦¸a��U��'̺�G�Y
{�b�AN��Hٸ�
�'���	�n��Q�tX����A�'qΤ:�B�60�TD�Ɂ�bT��'��p!��ݗ�v�B�����+�'G|q�d`؂0����E�I�K�'���*�jǫXd�F��1�i��'��R�	�nT���2��-�����']�]�3�'G���c�^?*,���'�R���2��:E�&����'rfI*�/�D��@E�2�d�
�'�XIA�4d���wDW5Ҵ��'(�i3� ��5��U�k\4�
�'1д ŉǙ
�f��E�F�(m��'Uʰ˟�
!� �)�ܨ�s&�Z�<��/$�����C�%o��@`�IZ�<����l �{��Y�{�v���RW�<�-��q�|P���3T�t��!�\�<����}+00�S:,�ܔe�VX�<��B��f�T�ce
5�Z����
U�<�$O
{Ѩ@���V;���2aR�<a��k���scF���z ��U�<��|o����î}�%����S�<y��T�X���C��W�jy��ʁO�<a��O�������%&�|��B�T�<����u��S h��\�ZA�!��N�<��W/^yI���>	E��"FRK�<A�5IJVd�%��=P��d�p(�R�<�Fb \��Piؑ4����-�i�<�&��y�ZZ`�T
o��(�D�o�<�P�3 De9A�	 b-�H��d�<�Dͣ?����P!.�����NK�<����.6�d[��x�x�a�ȅE�<Y����Z��sB�H,T��vH�U�<ɴ鍱+c`p'G�w����e�X�<!a͐Yn���c�T5�m�gȒj�<Ɓ�
����S�^���P�(�i�<� .ՁסsȌ��&�.��QH�"O��3po�9v�n����Z0J�+�"O����JN6��ᤊ��b"Ot�� ˊ�R�ǌV V%�Sk��QcUXCCs�l듿?E��OD1�o��H���+`�>c�I3%��?;��7�D$9��ɑ  �.M�D�[S�9���i���k�ƔB#.>R"a��._/�����@!Gdx��\�~��a3Z}�F�b���_�kRLW:&��Z6 �pp�hՂ�&`�lӶPn�ş����>U�H�9RM�A(Z�6lx0Gd�P�B�'�ў�?u`�حV�r��f�:t& �d�*�ɢ�M�B�i�'W�Tt�O���o8/�$MhÈ$w
�]�D��~2��^47�;<O46m�-:�(��P�r�|qƀVD��|��A@�_ňdmFc��1�l�-r���'<�IXJ�[��K�9�� �w(�3t1�м|e�d(��E���0��k�!�iQ�O�!sG��"bK���A/ȈV��(I�Ý0v����M��iK�\����C�I�jy�<`�ꍁ��)�2��J"�<9�a�F�顂>uVLU9���V���Gf�Z�On�a&l��J˓R(u�ŷ�d7�1Am�Q2��-Iܨ������xR�'����ժ۳<E�8z
S�#�)T!= ��*�79�V��AA)��C'@:�(O� �t,^,
����e獱����/^h�8����=��$�3+"(�
�����x�'��	��<P��#"|����vBH�]�V٫H��O�$�O�⟒�f�zR)�p�[�ެn���z�>�Ao�C���Og����ܞ6霑��˒ �Z�jt�릅�۴���U�'"Ȑn�ȟ'?���c�@i"&�I#_X��x�H�:g�4�O��dLO�he�^�] �YK]6��BĄ�R�	 F0j��jÍT1��gUw)�OfM8���yo�Q����C��A�jR�u�4�8���nE..V1��'SSjV%���ԚUr�ʅlџ$>��k����823�5k�|��'�L:��d�<9�S���oH-8�g��"d�U	���msa{��iaR7��>���׃Vm�H`'��l ��b��rx�TdlӬ���<ͧ���}�!
�T0�,�3#ѧNN(���i�.,hhhJ4ƀ(_�}B�y���D c^�S�?�zw3�DH�0)�$/�(���ˆ_��P�dɽ9���Á�l�~���=yA���p�i�ɼ��K߁/;j�ru��8\���V�o>��f��ݔ'�^}������KAE�+c��A�#�&�0��aNP��R�'�~�1�!�I9X��D�P%:��Q�{�v�^m�n��?�����3�OX��V�XD�2hHָ�����HZ�K��M�ϓ�M�#D�w�l0���� 2�i��*��ӴOǅ��1k�C=X�z��3dR'M�����l��cut�aT!�KGL�J��ÔR�4qy6�JN5���5��tD��X^w;Tl~�'�k�f�"$���͋�8��qݴc.����;�M��V�	�t`-�PEG09���9����Q�ș��T>�j����C�0@j6'P_rx�oЮ=�Ƙ|�|Ә���<���?����� �  ��   1  R  �  [   r,  %8  �B  �M  �V  lc  �m  6t  �z  �  5�  w�  ��  ��  ?�  ��  Ƭ  	�  M�  ��  ��  �  _�  G�  ��  (�  %�  ��  O�  R ( �  O" �( �(  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!$��E{����K9��)x0+ӎ9zX�1�'���=��{"N�"QJҽ���U�G��L��ͯ�y��o, �i]�u	�Ÿw��3��'�ў����x��ˠ�`4P�2�N��"OR$���9jܹ͊vFD �.���	��0<Y��D#Zk���"�/�P�ăC�<����sM�g���^������N�J���� ��H��>�2�d,�Eǧt��Iz��7��C�Iw��ņ<g������ۓۂ���I&�0=Q�&�%%kЅеj��E��51��`H<qƋ��P#�Ҕ	����	��Ռ{m!�(3���9E��.-�̠ �n�7xmQ�1�'�L�O�0X����1��<b�h��v�>|h�')�T��'�M{�qp�@XF�py�'k��'�S��ha��j�v.���F+��	$L���:Z��(��Ar��-�4����*D� ���@$'z]"�j�\lš�*D���@*�_�^y�A��N��,#�-D��HVݭ�H���&x����'?D���Q@����%c�{���*��>D��b��Nc~����˜�[�X\ra>D�`jpG�cB~ī�hMx3���,6D�Hk�Əa�NU ���6���	�E5D�*�KHeVTy�SiˎH\�cj8lOl6m"񄀝!`��Pƍ�rHp��iF-s	!��ύ�*�z�ĢuAgI��v�	O������&K�g��T���D�L��Py2j�{�0�e�ۮr�2���R�<�d��OD���U%5D,���SP�'�?�sN�+�%�rȑ�W~��ҁ(D���cJ�+>,lhD�X ��Z��&?���ԟ�O� �y�#�tpJ�ɒ�XV.`͛R"O�Q6��d���3��Ց?���|�R��G{��&9��ŀ~���fA�1&xMH��'���)ش^WtUu��!dͮ	з���z�DP�ȓe�&% ���-u������C(!��)G~b'A(�y��1�	z�Rb&2F���BT��=@�c��m�|���O�6,;��� ^HA��g�W�v�
�{#)�S�ӿ"b]bBЂ@�H�BR*��Ll�B�ɽq
5S�Ȭ�0��GǑ�y+J��hO�O,��V�<� }�P��T6�aS�f�?M��OBɲ L�.���A��X�kZp�����}?9��	^(p����B�;T�09�s��`��|��xB�H�!U�EYc�(���*��)�S�O%��J�m\�U�b!C�"�2��
�'�4���#یZC�$3�.����p��#OL%��gK+E���i^�$��l@��d<�S�S?B|t�AMܦc/��"�� yb|!��N���eH0j`���e�~��8Dyi(O�(�l�1��X���E|��!"ORd�� ��g�L��)�@q�#p%��t�'�ў��O�MJG�M�)��E 	ƏX�\�r�'W�'�b�n->.�=05C�{���S�'��)w`Z�b�ˤE5p�N���d$O�`�3)�#��+'g�	�صI�"O���BGolВ��H��L���"OB<��mF�xR��6�[�Q�0��"Ob��b�T3&܀[�N�<�ӕ�iў"~n�$fi�,q��m�y�3Oe���d	o�j��u��̌.ip�����`��f<��m�pƆ\ss�3hUD�\R�D4��[�'Hj�Ņ4�	�v�TN�)s�>)�-��d	��*5���t��T��H�����E�gf>�#�b�.SX�ӳD+u�!�$I47�|��n�)a�jm
�/q�qO��=%?Y�QJD/p�f�B��B,S��I��2�I��HO�O �<�u$��fp�"�>�f��t�i��'�ZY+��`�E/Y�0�"�d�)�p�+�=D��s��-!�^4�b���.Ƥ��x�������cT�jQ qMX��?��'��蛶@�=���r+ ^��Dxӓ��'#x�24I�"�T�9GDXa�ę�ߴ�hO?76V�ղ�撬e��Ǡ��p�剣KQ���?E�d�ˬ\%��aJтW�"$��Y��y>}b�'�PR���PDRFh/uJ2���}�E�cx�lQF��(h,�4ό2fB�-I��*�<lZ8$�Ј���agX��!J�&�RC䉅���Ê �
���@��I ���6ړ4m$�����D/B�[����L$�XC���) 4@h5-��{�LU��U�a}R�>AR���m���Y��*"� ��W}쓗p=� ��H���i��,�s��|�'aў�x�����^\����Z؀�`�"OX�3��	'4��L3� �rƬ#c"O��D�@"Dz�eaG�]o�N@�"Oy���!��"�hO�_�0 "Oz9q��� �z�x��TG�9j5"OR��Y00��q�A� t�"O���A9$�L�*�jN8(��v� ���B |�V Н2� SǮ>)��|4y�w䋅TIq�\�6|���	f����<��JK�o�8,���
�Wฅ��"|O�b��M!X��I�p��ߌ�����<I�_A8�@c�4z� ��Ȇ�mp���	Z�I��bW��'��:W��:U����Q����� �E�U��CJ&4ٔ!��%���Z��Ir�����:)LIC���/�pIs
�$0C!�DиIkS���H�ڐ�E&]I!�%o���Ae��(q���ڦ�0+���'�q����E �8I�DM�0��!r�ᑘ'�!��#��3Df\%��C'=��O>�=��f�"�N�>�J���g��Y�p�24�\s	2^�t\RU,ڣ@�0X4��O����S���D�0X���A��Hv�� �1\�9���>O�ق�-�5�t�U-�,5�ʭA��>�����B��<Ӡ�)�Z�R,�T6�xB�%n6��i��?P�X�E�JC���c�$�I,��<�ĩ/ډ2r@��	!��2�~�<���Ęw��C�'I�`��AC@�<i���nǊ�S�R>�T�)�!�{�d4�O�h�'����pq��bOD)��"O,i�Q*�=�X�
�>9� � ��:lO$�[�D [��Y򣊕|G�y
u�'yB��Q�D�p�^> dm+.�� 6���p�h���+j�|h��˫+�h�E~�S"m�����)�3*9(BI(��B��y޸��D"R/tQ��ˀJQ�-β�hnZLx� ��b^�`��A����%F��1sA#�Poژ=a��S`Z�I�|���iTM��C�	�,j�x�o�7|@>�i6M�e���dS:�(O�T��^)��A���?9�h�"O��cR�XɎ]�U��2~��iB�"O�A�E,m<x��ǩ"k��� "O:�����^����%�ڍU-H�y"O���Dk�>i��qT�S=2��$"O�\��Т,�e�p��1&���D�O�OX�S�3?a��YX�!+�D�qDE��z�<QJ���Z�8 #�޼ň����x��l���D�V�Ԍ����=��u��P�j�c�Y5)Ǫ����pB�E�ȓ'�L��/D�B�`�C��U����Y�L�z&��)mtP� ���(�ȓH�DQ��֤gզ�@A�R�k1XH��@J�itg�CT�aH Ò( P��`6���� �4��E($`�"8F��ȓ,Td���%�l`�,Co�6��Fh4��)�=`����?n���ȓOXq�ޜf��	8�fS;zb5��2t��ˇeH�1!��7$|h�ȓ+�"���[!h.E���ïXRŅȓ7�z�c0J�y� ���ǠN!ԩ�ȓ$�99ФXot��rF��d)��� @c���ep����A�s;�`�ȓ!�r`2d8+j}Z��e���	�Y��"���,4l��"�H�q���H�,8�N˾a�Ρ��S��ԫ�ɉ?��}� �t�>��N���q�`�p�*�*
�e�ȓx�tu��F�9mXĻ�䏊u��-�ȓ[ B)W��t�(`Ն����ȓK��+��$0�ĭ36�I�l�~8�ȓ,�}�ѥ�;nX�k�#�n�9����9���	@�6DsV,N.4�*݆�uI�����	Dvq@S@�4yWL��(��J�ފ~�K���G����ȓ
��a��� x�|�dC]�J�X��M,�� �X�5D���r�-�ȓ��P�vM��-!2qإ���<�b��ȓg��dX$L��T��Axq�Ijhԇ�S�? ��Y#/�h@�ͪ>��`�@"O��+��I�m��yx���5^�	9�"O\]8�B'e�hr1�ر_w�p�5"O�c�hyj�OG agPB "O��s$E�S�P(��M Ov�9���'U��'b��'���'��'I��'tH0'`Q�Pd�P(��E�5�$ۦ�'�'�R�'�2�'j��'���'���!-D� 8Bd��G^�1y��'g��'F��'�B�'X��'�2�'ɾ�2�Z!-�"�$]<2m�����'��'\B�'���'�"�'�"�'6��)���=PRe2ć�
%�$(���'.B�'��'���'"��'�"�'%�5h(��|E�m��٤J���"�'R�'R�'���'t��'���'�t�PDC
P��C/F�$�=��'5�'L��'>r�'���'�r�'�h�BƸ��)�&�f���$�'cR�'���'��'���'$"�'Wh@�%�C�[+�T���'O1��r"�'���'C��':�'|2�'6�w�>���'w��"tU�7�!	t�'S��'c��'���'���'���''4��	�}��5s���o?�j�'�r�'���'&��'���'��'�&8Y�
�LHY1hɆ
����'u��'��'��'�R�'�"�'{*��1��4"�q��*]��xi��'|��' ��'���'iB,|�x���O|���� @���I��T�Y�DMpy�'E�)�3?�'�i����e�� E�t*a��{
��*�#�����-�?�g?�ߴ���jTK	�h�Q��&Ȃ?¤Aȁ�i����,p��������tłXR#�~,��c�FĚ�O�7W#��{C�_}̓�?q+O��}J��]��ҥ�U���W"���;�VCT���'�Dlz���� Q�O���f��`-,��Q����?��4�y"\���:�"�Mp�l�ɧh4���'	�N!�a��f�#��	�Z��d�t�Z_��D{�O�R���j��®Z�U Y1G�F?y,O�O|-l�j^c��.YdLi���ɮ"y�q��OH�A�n�ȩ*O��Dw����U}�w����JS�:|���%�R�����2r
q��L$�1��i˲�t݅��H溥yWƷ>�(���&}�"��,O�ʓ�?E��'�N��C�R�?{�|�uQ�s����'$P7mI�1��	��M+��O�b4hE��l�!��Y�*�)��'U�i�rJ�������z�q�X���� T������4����`f��	$�䕧�Ϙ'?��/R�=�I@r�-oi�|{�Oo�����'�B�	݁J���q�Q	rX؀��-J#x'���'mN6����MaL<ͧ�2�'	�v$�e�MU��PƧ�ld=k@#�`�J��.O�yPwl]q|5r�݈ Or9�E��C�PqUFT$9��Z�ف|c�i���C/)� ���ԸMhw'��f�2"O�tTf��
ԛHLCɺ�U���6%��\5/8�x��S�!�����$71A��tj[[{*%z l�Pl!�SH�F��� �a�;���yT�F��vu(��Ld0~hI��I�Dp�Z�!$��Ed��l	8��I�7����Q�APX�H�V�ֻAnu�fN=V�<%3�Ɇ�x�@�[WeU0p|΄ÕN)$�<����N#���t`'c��;b�'���[����}9AlB/w����NkӼ�$�O��$7��O���)l"���bo�0��´��A���]	8�DD�'%b�'�2R��X�$�w�t�'��(��V�w��0Ԏ6�,��fiӶ�$1���O���*�D'}¯L�8BJ�2"ԥH$|9�T���M���?�,OfXr�F�|����?9��4q (�0"��}�*�@��t4���җx��'�b�K��|�������\�uOJ��bF�u��6�i2�	b�=�	��������{yZc+��R�<Py8R�V�~,b��ش�?���=n6�����+F�R,���SaF#�v�
���M������?���?�����,OD�$�O �z�턣0t����Íro X{�`����3��Y�S�O���gd���C��<}`D{�ͼ�6-�O ��O�Qc�<)��?Q���~�[7�<:�J��4v���6��'C��鱝|b�'2�'�T���m�
����R2x5��BӾ�d�:��ʓ�?���?�K>��3:���GO�9\�� ��
�?_|,y�'��t��'[�����	˟h�'�"d�P/`�25G�
S��)Õ��6X
듺��O��O(�$�O"�
�A�M8l��F�/CYkb�3=�1Ox�d�OB���<���C���$m;}������+�A�a���MK��?���䓾?���{��tB�'
������SV�I���_�0ѩO@���O����<!��@���)�O��ے/C��&}B`���1�&\��nɦa��l��d�	.-�b�|3p�PX�P�������I�mx�6���O8ʓj{% ,�0���O���T�)�DU�el��.�����W���<'����h��[i�S���ҟm߀�	�G�u�>���&�?�M�+O�M�)�O��D�O��������a[.Hl�X-��=�<�����e�I��01D��ş�&�b?�:w���lRA�%�R�yB�Q�QOu���f-�O����O�����ʓ�?��[@`��Q�4��R1�I&;vЊ��iy�+���S��h�b�w.�P �I�H�@�U�ס�MC��?��r.�"-O*���O�����3dO��m"�<��\fdp��v�&��" �`Q%�|���8��=�� �)�� Bv=�0�3��ՉS�i�B��:`��O��O����<!+W� P�9�f��H1���E�?w��6�'8d$��'��	ПP���ؗ'e���W���/,0��m��`��:�H y]>O�D�O��ĥ<Q���?�7l�o6��f >���	
W�&\�����D�O��Ļ<��/���x�O@�M���S��lx��B�EY�|�޴�?Q����'��'d ѓ�/�M3�/�(~���V&�=g�T򳅖x�Iğh�'�bn!5 ��P��ES�)��$Y�)"@��pA���MÉ"�'9�a]a�Xu�J<� n- §�͒C�T��F�a�	Hy��'��R>��	쟈�s����%H0B����N�K���*�4��Oz�Ė�aJ���T?�X&i:Z!j�
�bt\����>��������?A���?Q����a���ld@��I�D�1 �iM��'AF�r�fH�����O�x
̧N΂ት��Dm,A�4�ཉ�iOR�'b�O�:O��
�y���$^�t��6�J&\{P00w�i�؈��'���'���O��Sn��OC����ld�h�����p:6��O��D�O8�&#�<�OC�h����_)
�v, �44�s���ݙH.�0$>����|��z�*E@�u��j�/�>)�|�Y�4�?��!Ԑ,N�����'[�_�*�,�$��dӣ�S�%��ubs�J#�Mk�]~6�:�����O����Ob�d�n4h25<��#S�4^�|��v�L25��'���'h�V���I�x�ճ9F�3%�-�¸��@�>kڅ�I{y��'!�Z���ɤ0���'%C�����St�(��r���m������~��?��0�4�#�����Qϔ ��mż=��=Iʪ>q���?A����d�(Zj�$>qy��2@�����ϣ#�\���D�MS���?q,O�d�|����)��=��,�sE�h�V�dT�inZ���By��ql�d����k�:/��ٰf��X.���n,��U����֟p�	ܟ�OX�i��9L[3.�&� tE�A�t��Idӂ�$�OT|"ШB���I�����?����Ц���\��&�E���L �����OhLB���O�D�<ͧ���"Rġ�r�X;f�,`�$N,��6M�=EV�o��I�8���?��	ǟ ��q�%)�`���uaNB�~$0ݴ	z�;(O���|���'j��𴉟#?fX�	F�RUn(��x�`���O"�$��3jLoZ��	�@����]5o/R!��CC��T���&�D6m%�d�E+�?���矼��� r٧I�%s��	�</��(�4�?�5/>hW�&�'�R�'��~b�'H\��� 9>f�q�H+S�<�'A^|��'����	�(��ӟ�;!�ó6o¤�a��n��Э�,'  �p�4�?	��?���n��Oy2�'#r�۰f���I� 2s,��1mȆ�y��'}��'��'���'7H��hӠ`�wD� +��aj�O@�~�b8xU�O�1�I����Iȟ���Ly"�'^��+��56��?\�t��ËՊ�=�b2�M���?���?Y�X?�Q�m�0�Ms���?��K�O_�93�戱,7©2�D�!����'���'�����4�3�r>E�IП����5�,��sG�3�E{�Aæ�M���?I��?)D��7h���'���'��DoM=�B(����Ľ�"*ě4�6-�O�ʓ�?Cb��|����4��Vl�<OU��P��۵h�dx����M����?QElZ�9���'���'����Ol����%R�Y�����ȅ�B@E�J��듭?Y��՚�?����4�
�O�>9H�,=ͪa	J �����4v���is��'�B�O��$�'�b�'5�x���̳C���P-D+H&FT��u�p4�J�<!)O��ɟx0�Ț�)�m�V�~���� Aʟ�M����?����t9$�i�R�'B�'�Zw�$x{aMZ''��+2/ثE:6uxݴ�?�,Oh��d>O�S��	ʟ|{ѧ�mg����U�G�M`7'U7�M���}Δ�j�i��'9��'���~�χ;;�D�e��<|�� rW�!��$�(<��I�\�I֟�I����1`}2ǆǐ%�h<*B��%hXui&@Й�M���?i��?�S^?�'=���4Bl��N�]�\$���łG,ys�'���'N��'?r�'�2CG@�*7��o����Y$(^F� ս�7m�O���Of�$�Oxʓ�?���P�|��&Q�j� �7LS�IK�]�E#H��F�'�"�'�2#�~�e��=H���';��\f�U+va�0t�U	6#�1Y�Z7�O���O�˓�?�jT�|"��?I`���\�S�j��u�c��5'B�v�'`R�'s2�
!(�6-�O��d�O.����H�4�@.P�1�fD ��lП��'+r�������'��i>7MN�,"��Z2�C�E}���C��4>���'JRI��[�6M�O��$�O��i���Ĕ�\òe�FP�R�D��	ľ,U��'�B˘�l!��|�O!�'��+��Ƞ�rh b�W=�o�v��]�4�?���?����z���?�����FV�9k��c M3S�����i�]�"�4�1O����C��=Q���! �e�.��6�>ql��x����hrؙ�M����?���?��Ӻ7Nl�y�ݏhU�e)��Ϧ��	myb�HQ?�O���'�N�|��E�E��V�	r�ƥ_~P6-�O(�@�ʦ��⟌�Iݟ�@����	&a�J /F��6�_	��h�����?���?Y��?�.���F�]I�~T�j͆<k  �����^�,�m�ϟt�IƟ4����I�<a��|-�1�kt��<��*��؃k	�<���?!��?����?���l <����i�~� 
ݑ��P�0�H�7~������i���'���'��Q���I��P�S�7�R�bA� �*!��A	쩐ߴ�?)��?����?��U��b�i�2�'�Xh�եY�@��aǆ�&Cii�x���O���<����Eͧ�?��'a��9��O�<��qA2 ,2�Rڴ�?��������,&>9���?�9�i�$#����ԧ�*�R����A2�ē�?�� "�Dx��@١�:9NP#�L���v� �i��I'{�j`SߴH���ܟ������#R��=�q�[�XmP$N�3��V�'<Rk�y�|��t�P�)�ґ��#T�@YTA(Y�M#�F�9ٛ��'��'x�dM;��O2LID*���Y?TF�IX�J7�7	'���O��O>9��Dq�qQ�g�������Տ=��+ڴ�?y���?R��F�'�"�'.�d"cvX쪆hU�?�0����+n4�v�|���"J�h�����O&��Pl��G(�4��
T~/.6m�O��3�]f�Iԟd�I�i�i:�f��'hl�1��mP0�Ĝw��ɕ.�n$$����؟���ByB�Rjd��#F�$:��d*�+�.�����I(��O��1���O�$��r���-� (|�r���-Z^�aB��O˓�?y��?Y,O��kP���|�$K��$:(�a��(|1$8+`]d��ϟ$�T��ϟ���D��T�1@����NĚL�)vi�<��D�O����O���l�����dC;�A*w�G)
�� P��IPN�6��O�O����Oֈ�df�O��'�zԈ���^�����b��ڴ�?����DF#F2��%>e���?���J�&�*)	��Kh����+�ē�?1�5�*Ȫ����S�$�Z�m�4�Y���1¸��@�V��MC+O�բ4��ƦY����埬`�'w�%J&:\`�3�D�1>��3�4�?I�+��!���S�Q.��q�/\"�zp��$��V�o��Qܴ�?���?��'^��'��$r����@Gu��(�M� $��7M(��2����W��Q�F����T�2��!��P3�M{���?�&��%���x�'-R�O�4�'eh�$���,n��!Q�i��'A2��Q�2�	�O����O�IT��`�8��H�H��զ��	)]��5J<ͧ�(O���tf�<./J�Z��N,O�*ȓ�i�֥N�R�'���'q��'�剳q/~]��IĊQ�"�Q2G˰?�F�z��/�ē�?I���O��#N�D[6�q��R�%f&-�"΃k����O(���O����Oz�cϜ���0��E2Ո��#È�/[BIr�Q�8�IQ�'DbdƟnq2�Q�F��M����5HH��A�H}�"��?9��?i-O�!�	�r��zI^��5�ְq�6U)ضf�Dbش�hO��$Ƀ)�$�O �S-r!��(A�jx���M�sG6��Ol���O��$ˆw�	oğ4�I��t�S�`��j��>b����,V�f�3ߴ�?�,O��d]+�i�O��$�|nZ�)n^85���Fb�1ft2�H5�n���D�O�8 5l�榩��ٟ��I�?-��ڟDz�(q�ڔpOT0��j��ݮ����O��8�.�Op��<ͧ��S0�h8Z1a�?�	���R�j��6M�
j$��l�Ο �I�X�S�?��I�\��=Y$���/L�~9�3��(C��l�ڴlEA����?-O�7�I�OTA�U(E����cFX&h����ۦ����(���3�� x۴�?����?���?��)j��Q.�`L��i�H��mZ� �'�;���i�On���Oh� �AW�x��1��'T����Μ���	�i��zش�?����?���T�{?��.G�N�� w��^�����Z}"C��y��'�2�'��']�SSƕ*'J�w;F�a̗l��a���]�M#��?���?ib^?��'x�E��S{PqA��C�0��`>"D�1
�'N�'��'"�	��@�i�Q��|���EA�qP#�"�ڦ�������	N�����ɚrب�	x����@H]��r���,R|�<`:�T�@�I�����Qy�E�u��:"FI�{I<���bZ� �
a�wcڦ���c�����I2v�Db��gL>S�6��@&ͨeR�!��`Ӿ���O�ʓ'�нs���D�'��dMM{��	�ҩ�of�ջa�	V��O����O(@ ��~:qR bNibja�p$�aʦE�'��I�Ly���O�b�O1��s��,!�/ӫeP����X�h��(l؟`���#<�~�r�I�<x��$BF'	6n�����T��AFZ���[8��� (N� ���X>Q�����aD	!�lYtƉ�y���;
Z�C�I\�l��ћp&��V��!�:z���k�m�KZ�˄c�/"
|&K[�p��1[�%��B$NP�D�"��P�M�XE��E�3{!���`#JKr�P^u��Sv�ʖ��U�J��(�@F�9o	�@���G<.'��9� ^4�x�i��B�L���)AU�'���'$���ß ���|� �J����=ݸ@:E
����6�Rj���$��H��a��V���Dy��Ҕ:�J�x�Dאt^YФ�+y �AS��.49@���2*J=�a�]��1Dy�	�*�v�) ���fU��k5/��<4`����?ɏ��?���]t	d�P�f�,�e � RVB�ɝc}*)Y�/�$��h;CH�6!�b���ܴ�?q+O`X�E�F���'��Z�KY5!R��s\�JÊ�K��'�R͡=f2�'��I�.5L�ۂ�Pl�VJBim�~�!㉨���J��((��̓��'����팾P�����)ҷhE� �ढWQ���ǥ�

�*��R�u*�#>q�ʟ���iy��K�*\�5cï�	��c^���'�{�K��v>phђ��(���,��x2�`ӨIp�f�E�j�q�4㜼�v��O��Pĸ�k���$�'��w��������&�D�5�Y�.�����(�p� �j����� � 1n�5�����	�|�D�y<��BR@��f��.���'UZ�`� �|����d)H�N[�8K����<��?�ˀ���(��I�Wˊ�8��I�e?}ϖ��?��h�����9{CT)s�!""�0���P�!��Լ	:.��b%�	Lx��*��*tax��9�_�l0C
%$�(r��A`�|�5�i���'�EX�)��t	��'^R�'O�w���Q��q�-h�/��=��,�.�a���ܦ�U!
h?xc>�O���E�Ⱦ�F��ӆB�"ČI��D�d죳k���M��BU(9�R�>�O��a�ȗY�j\�fC~{(�Z&�ަ���4�?��ߞ�?�}�'V��)E����&� �	�!/���$\�$>&  �.b�����XA�ɵ�HO
`j�'��	_��M�eP�6�-�)��E8]�n=i��?���?�������O�&��4y��V�'��I9�����
Q
�5!���6㍭B7R�hƠ",O��E�L���Ql�=,]��Qa�Y5l��u�ǔ;�,dbA��0axcU.��@�( �H t`[" ���i��?����'d�ԀS��BL�j4�VJ�9F~(��0"O*-��E-��I����q~ڝ�$����	sy���rG�7m�O��Ŷ	���vEB"���"6����*�$�OSѩ�OP��n>�{%B��'���%��M��h
�O@�BȘ��I�J��p���]����D��:_���{)ka�N�&z�R�CU�	<��ar��1����gj�NT��e�G�'^Rx8�o��v��>Y$FS
�,4���6�. ��,��<y���?����*X��}�D"�E�,a�T�ЍI~!�\զ�ci
%"��E����d�)��ܟ��'
�c�`���$�O�ʧr��������H�I�<`����4#O0�y���?�1B\1)���C��0�09"�i8��Q���l��) 5��L�����=��-��{#ܝI1ZP�J�m�O��ȋ���*9�h���/I���N��(@	�O��ۦ��I{�'j��53eŏ�S�:����S� ]�<A���4ړ1�ry6倱p�R,1T�vvv��I�M�2�i��'�2yA�NN!�v1���3�T�	`c����Ol��݁&���Q.�OV�D�O��4��v�!8x8<��!G�s��'x��٫�e��G� H!N�b>�O�R��v�V�Ie�cӀ! `
�'e�Px��E:�)�f@��So�PÉ�L>)����B�:QbI/O"8RA ˕�?	��?�����?�}�'�r��hIbe�v�O�El�A��iū��񤁽f��c������p�@;5E�	 �HO��py���"�,�JJ�`����e��+�\��0�I)+���'""�'��]�X��ПLbS�O��p@i��;i���bďI₈�#J)�Of\K�m�� KBu"�_;�x!���
�޸����>2X&qs�'nX��N�/nͮM�vD�2V�9�&�?�&A�'	��'\�O�U�D�<���F��������	X�Ae�u��i�B��E��%�@��4%��6R��脤�M[��?��fG�@����یu��$�E����?���/l�8��?��Ou���R�H���UԲ�W!2a2@k�j��jG���%�H��p<�"J�CR�8�(��9�޴<tf��v�E1hΩ9'nť��T��1���$����ܴ�?qS�
è̚"�	�t~t��a���O��"|�s"��O����EJ�(4��,���^<A��i��qh���sX�8c%�9�,��r�'��I9�֌�	����	U�T.�B3,��Hp�O�.��M���4���'v\���֬O�N�	��������c!�~�.�<��Δ,5��	��Zxt��I�>Ɂ��� � ��� H�c�X=��
�	Uq��Mע��M2����o�@�Y��>���8z۴/Û��'m�O���Ǘ�f��Q�	�����B�Œ(_2�'���'}��'+ў,����8{u�3q�D%R�V�A�-O�%l��M�L>�%-I�I�0�A���D�PуZܛ�'���'�h0�si�<�r�'d��'���2�|���	�?v��[Q�F�_6��r1͓�/�A���3�x�D�Pr�g�	3Q1�mz�Z+xC�= ą8+6�E%�='�`5�%��$Y�سӃ.�@
˓h��L+(A��<6`_��N�Z���?���b��X�S�gy�']�e���X�B�{6�(��O���#�R�I��<�C�29�E������$ɣ9F���<��.�0<~X�@F�op@9�c@T�`���"ʦ�?��?��=�n�O�f>�����!���F�̋%l�% Q`�y+~<����XD89Q@�i����qVIR��5\E:��@	{x��a�ؼc�T���O�~eꐀ��'��� *893OI�:�����-�G^,l9��O$\nZ��Mc����$�O^�dX�J��N֤r4G0%�V�C%D����Ŏ\��l3�`N�J�*Ģ(�5����<ywC|k�I̟�[_��H��'��<}�ґ鑯���� w����Iڟ ϧ0���q&���Y�1xrI�:��L���T��$aN�Gd�påM��p<A^�)2��A��4#��G[�����)�(������P��J�@Sbin���'��L��FȲ�۶!��ُyb�'��yGa�����DTs:,eؑK�x2lx�`}�`^���;���5�ܭ�19O:˓9f�k�i�"�'x�.T<��IeL��Q��:����ĭM�z�� ��֟|1��J��`ȴ�A	e"L̈±��	�|F�tvH�!@�V����r��s�dޮu�㎿]
P��i�0����Q���B�-pD��$�#r�h��o�!��F�����OX��Ɠ��pB�)X�F� ��L<t��S�D�O��� �E�hh�h���A6�� ax��?ғf4�2�)��`��P���Cq�iAb�'�B�
%s���I��'!��'t�w(�[Щ��}�v��0��AȠ���7�`x��!l�h� �Y)�Ϙ'�%IRl�-Zyx��W*,��Y�V���Tl��@��]2�r�(��ظO���'��<��+ ��%��]�1L��&m���n���qG�ß�>˓�?y
�)b����X#&A�C,ޝ��D.�S�O5~�Y0��#��tу�N�{*T`�O��m��M+H>	-��ʓh���I&TΆ1��JH!XN� ���#,FP���?��?-���O�dd>���ϟ.jy���	�&`��i	4Y���*,�����ϭ�MR��� 9��!�4k2��Ö�qyxdJ�|`�qHW���+��eZ���Ã�B�9�Q���s�ԍ=I(��dV!L�@� C��<#����7Ma����4��V���(�kr*	"�%Ɉ0����BԨ�8W�ߢOL��dF�N0}�<��i
�[�q����M���?��M�Pr2q���1{��vl��?���+f�q��?q�O!����g�[�D %*Q����
��*�24�X<-{�\[�o�/�p<1&�\P�jt(I�#K�F��4(�a2PJ��T�����i^�l���ɩuv�������	՟l�H��%� c���'�� k#Bޟt�	���I�L%?�'���$ Ӥ`T �Ul�)����(<�h۴8KM��-��} �ά\Vpϓ��d_�vamZݟ���J�TbI�h|D�G�d5�nՃ;�!Pn�gLb�'�̹�`��#�x\�"_�p�����XX"/�@<�DfZ�v��h���#��� ��>�n]�-fr}B�TR��RG�ޗZ�q�� p�Fن�(�e@�$��Ȫ��>A�Ο��I����R�'��a�&��a�tE�S,I�e�Lx�<�����<y��G#�d���_�f0QUd����şN�Lt�Q�D�q�L�T�ߎ��ߦ��I����//�mHf��ʟ���ş�����ձ���rZ�B�:ڨ��� #�P:U#�A=��RK!(����|�I<	4+��Gf���AS>�3A�z�Z�yEbT������`0PE�}�I<���X�k�Y#rOU�4����$�k���oӊ�d̯x���Y���	@1)���Q@�=�P� ($��)�Ɠl��ڳ"ܠgL��u�e���������$��~�T��{��� �Ꙋci�y�ֆ#!����d��ٟp��{�D�'��8z�>ñfQ���/�2������-.K��hV'0|OZ��aρ�t�(�6RAɋ�5j>�@cN�w�X�a'шt�d�D~���|�a�"��� �7+�]���lE�VFf�,���<1����'`F4)Qm��6X2��M����TJ�O����˫[HDZ�a��p���0�A�� ��O>�l�0�M+)Ofy���L}2�'��h�^[�H�$|��'��B��'��KV�"��q׉�?3x<jS����H�
R�3h�8	x�IL�~^�`��)��Z�b9�'>!�0���ϯۂؓ6(mCǃT�1���%��OZ`�4�' R�$e�(�Y�՘�i0�+�w�� \�,f �k�Ӻ3����
?j�6e�GiВ=���W���x�m�L���V�ﺴɔ 8v�̢��^ަ�'0h-ZrE�r?A����)�R���$�3���&�� ��B6ő�����O����1Rs��J�
֕�������+3��;��|*�JjJ�R*��5#|y�"aAt�ĞT�H�ΊKi@��1`&J���AI4����_��e�` ,�
�����#��[?F�I�M�P��?��u#�(WGص�s#���2G�Mh<�֣�|���3��]F��yS_n���d#_`r s�:'*�(��E�|{�AnΟ ��ҟ��#µ8���������ޟL�\wX�T�4y8Hᢏ��.�C�Ǎg������ɞ-]����o�%41�\O^d��kƷCN��є+��~3��r� ȏ��J�͋w˄��$�4q+q��O�L{tF&?�����I�2.%z�e�	��A�,O�})���d�OQ�O� :�I��<n�^�P��|���U"OH��d�_�j����ϤU
z�Y���(����F���IVy��ɚtp�����>2n�yXFa¶�y���̌�y�E�'$���0�L��yH�ᮄP� 	�|X	V����y��-Rp�I�ݱ0��FkQ:�yb��_(�5�G��	g�(P�s���yb��Y�x�r#�7Z�x��ր�yB��) BڜS����7+�@([%�y�C�_; �HC��	)���B�*�,�yrcC+,�BaC�(T�!�����P�yr&�9H�]���I2j�0�2t���y" �2"8B1��a/.��%�y�*-���:T#�ǀT �ߚ�y���9��Ux���.$�X,��N��y"�J�L4t�+��.TmD��쎯�y"FM�\z��R��
J'<�S���y
z���(�a�AJ\!��.�y�W8|z�����?���S� N?�y��{�X1"��֔W��sK��yb�S��8�r��3(���)V��y��Ț%���"_��z���B�y�f×(�q�"����	$�y� C�o���0̊e>
�B�J�y�W�"���D�C<3�����I��y���h��ջ`�b�� ˂d�	�y���5+p 4�Ѓ�Z�`���MԵ�y�n��<���#b�B�W<Э��ƌ��y�ּ*��e�t��,A�h�� ��y���bՙ֋�(��A"C��y�d��p:��TM�.v�1�)H���V�v�3�!X�o�&���	 U��=�G���=�Į�-��v���?�!��K�0a:�BG�sbB�H��C+�Z����3�t8#.�j��J��S[C�N�
H�X�'Z��� c@��&&�z��Wx@s��)�(!s�סoO|C�#�2m�z��A,�_��������_�� �W"%Z���O�lք�;3[�-bW�(i�
�˗�)~
�ɓ��!��1�-�6�1O�� �͏�_�=2&�M���X�I. [�y�q)�#�0��dή�p<y�M�o�����Zr�	fF��'\�1����y��t2$�p����T&)A�ZXp�e��h��R�
��D�-p�&� x>���E���{����X�;�G�+[���x���Dߤ��riS�H�݂f�'R\p���W�a����:Ȉ�J�E����2!��(�A�@��H��u�i�
E
�\qmR"1��f�(��޳T�L��\�SN,�<�\��9��Ԓ&*��Γ��M�<�1oP��D���lQ�3��%�G�0Ys�5CT�KM:WdO"
����_f#���'�]+7h�e��ȏ�7�tc2
�;?2޴p��H

az�ʏj�0�ђ�=8H����_>���S@�@���P;-�@�B��u���	d� XC�����A+`�<%nE
�l�YN�l���e���a���g�6a����؁�O:��j�hϕ?T��Q�����'j�Q �	ֿ4�!�����k��y�O��5�ƅ2����%���\���BE�0扡r��@A�@��n]*���]�8����?��9:Kl!: �M�2Cp���:>kԜ����C��%+7�/����'I��(U�
� �5��wG�Pіl�����
��N�s�A9��i���=}��[�daה-0���7BAY�d5Swn��%�vL�jUz�P�JI|1vd	��koT��֥V	Q&���OީjM~�$&�gWިhQ�Z�V\��i��M�`w�Y�$�i	�Ca����%��JW�B�,]� �'f�|��c �=I�¥*���8JQ"���˟ܑ� L��u�	��a��y���'�h1�l�go����܇8��9��y�̧xv�8�d�6CJ�`x��')�]��oy��	�t��B� $f�|����i�
�I���T���ܸO��q2�-O����WTs�	".�_iD a���
0~TC1O̰`b�D2f��$��#=2�H�w�ZU��ܵ:`�r*^3DB�	�*�v����F1|~��rBL��9�L���bG;^�j��
	gD�9����|��Sܧ3�������k����@�u��0��ɕdz H��Ӛ���ش�iZ� �<�*��R�" M���%���U�`P�g�ȟ( �,N}��O��4�;���1G� ]��"�&k%pM�<��*�+�pL�B��#�H�>�)� l�#p��%�ȹE�*w���zV�VB�� �UJ�|���M��0+܌8��?�!��i+��&	�>fBx�Z�Y".����ޡ)���g.Ԡw���3�)�D�T�B�pg�A-�htrdk[o?1�+ �j �C��[zp�V�XA�'ĕa�
� 9����o�1N�ژ�EAL9F/�-�{���'��h9E��"D�� +	6W"�5�1���Dj�*���Qr>�H�Ņ�2v��r��\S7��$m�ʽ�ЃBM�$c���ቆ��	�̝l��iYC�ڵUg)���̞q�1O(��ܾ1������u��\Yq�>���?�jD��ɚ�	���3΁yʠ�>�wh�O�y�M+�&����?	*��'Z�e���V���-��>���H�ڡi��ޡ_PR��O��S�.�	��H�0�B:�����&a�4�8��'3��"��[o1hD��#�+2�J��J�Bp&��a�pa��O\ha4�$��O�tjNS�U�i�^-�DӔEW�&`4$�T�I�;� �S��GQ4�L��HѩG�N;���v)O�s
R�O�ŀ�)Nh�Ӻ���3�R���� jO"��V��,3hnE��ܣ^�Rb�D	��̃ R��,¸)u��0��&}��X
� �`2@��,�x����n��}b�K�0�� Q���0덶�2C��OnA(�%�%�&��j�v8p;���bق]��gҀk,��jc���`��f�-d�#�,�&�� �I	@�*�'��<2������S�6r��F{���i�4QC6�D�t�Y��\��?�BFd�IH>�'�OT���N ��I�(�!�<�@E��Ev�;�.��)�h�EO�λSP���F�6t�����LA�'X����'�@;��)M��]�ĩĵX[v�0u�M�ּ(�<1q�]�YV�)���
J]��m���s��i'�ɍ^�q0�-R�aI28@W���6"�����'��I	����$��ME�C74�:��\�|�K�L�*|��xA��� ]Q�1�q�Gڟ��g�SR'��;]�����@D�� �����<��_oybΚ?Z���k��!j8��2�Ȁpƨ��@>Mǌ���n��b?i8b� #u��y�d��i���􋈳^5���5.�w�����d� ?�9�Q��c�.Ϳfo޼�`�C��5�Q�G'|t剝o�\�O�4y��&��<�����1u��׍�f��P��1O�R�7[x�Q3��1]x�i����'�0�
_�&�B`��D�Z�(�'����0Ab���Č�W*� U �4AF*��ҩʮ���c Y4��L�c�m��(T�F��D�5�|R�f�1O���!���r'hֶ}<|�c�V����[���a�U�6< a�e8ʓr�r=(�֖E�y"��ڟ0�H �O�!�F�ǥ!��O�܉կH�fd��bdg̀�j=9�'۽}�iB.��(O�doܠPzj<;�?�\Y��NTn(8yA˟�s���͝%;�	=_�NIZV�Ff�3}�-n��9FO��f�,��J�G�H�y�
Z�M��	J�Ā�#t��j�Â���$�#�h�%
'U��h�R��=$�\����&y� qS�%�5jPi�V��dZ\����9b �ʳ�
�8��Iფ�8x칺chÊ|۬���4~Ȫ���ώK?�d�W�,&$�BTI6\6���O��\� H�*O�����4�ՑI��S�#��{��@�'��k�HZ�!"�	�SWH08��H${l>Yː䟴0~�`8q���D��⛥,	~I
�C ��~��)�d����-N�[�Iŭľ�]Bb�K�1X�U���!�)"���3�r�	�d�Jz�d����962��͆�F����O�̰��'Hv��9��O��s6��8|܊ �3E�ջm�8J���O;C�p��	�I抡�s՟X�PD�V0F�c�[�i��P��\Y�b�O|Aᢧ�(2"�	�$F�!L|u)4�4n���20[�:K�5B�C�+�.옔NC�����M >延�Ү	i�S�Z�@��Z�Kk�훒Bi>��'�
9;"|�B��7 ⑒@��Or��3#õ,�}r*	Id��	�/�(}�2]�?�WF��VH��@N�\�3pJ͕>�YkA�<(��Y���+#�T\�QJ�E�dւ?���'+hH�k@��4U���ΐ�{�ֱр��F4IQ�雽Qkў�3 �΀5�4�:D,8E��h�/��a��>r�BƆ[I�F�p�o�1���u%��4V�x�e�K<tXq0Uk�����j2�Q=]�x�i gX�'��� g��%�����l�::X��'3u�aE٣'���#��UH�-�ꂗ}�<9� F,r�>�'��xt�� X1ȴ�$H�9�세�e�'G��Ȗ�{v�V���)��Dll�)��'�l�{t��2H�Ɏ aҒ�8��N�gG~(��H្ K⩕��d�yu��\�l���'Z�@Ƹ��ō�69=�!I.��O���t/IǚAC�'��A#z�Y�K���?�p�$$=�6�ϊu�4��rʒO��؀Q����)1W��rF�Q��a ��lҨ�wm�'���N:F���=�B&�*x�N�%F��Q���i�T�ց�36�4X3b�Q�?���Q��=`�C���9O8u����aC	��H��8'�f�#&�G�'I>������$
TF��3`��ԟ>�` L��Hl:��u�G3�5�t��<f )�ª�_}Ҡ��3��0�@I4V]�Ÿ���j�ɟ
e("�#���9��97AΛ8��*�bI�D �3�佋WƏ*��T ӬB`��&�>9*1�	�7��0a����S b�Æ��>���� &,�8��|�<���ґAV��se��k�H����Q�;�.`���\qBnL�-�:c��S�M��I5c�⑸RQ{�m�s)�3|f�T1�!�kE���F�~�z�j��j��Z�v����UF��M��y��M1&.vL��Ov<:v���"��G�JN��@�M��W1*��b��L3az"AҋX�M���F?�Eϩ �\��MK�s^��$L�m�t�	��U~�MY�h["�8��+�h�q�[z�� �� �}x�b��J'����'k0���g����pJ�1I]�s�|{�n(}"fMq+t����&|"���ԵzGl6m��v��ڀ�Q�_{���R瘍nb�Ϙ'gY9�	:r�*@�CۈO3�ku���s�#��4���2��,EyZ�ɚk\h 쎆d��P9u��8=\�;�΅�A@�iJ�#�ў2�#^/��o��Q���(�l.Z8\����!�O�9�)�O#���'����@�ܓ"�m2C.��m7l��и[lq�g�Y�V6�#Eݖ[6��*�h�[�+S�W)zj%��4m��Ȣ�V�%<2��?�.�24z��G�xIѢџP��l�-Al�a�厠Ί)@�i�����+�r,��p�IEH`	��O|�#!ퟂOF��KǦ����Z����g��	�`�u��릡@RC��T~��6��6".6R��DW�[W|����
����A��9gtd�q��l}�e�n|�y##ʏo�v�Ik�nQ2gK��|Jp	�$,�xw!��8��e����D��ɘK�D��	�,;���;	�l���A�H���r$�ͦ��D{��G�$��(���J�-�;��T�OĹ�0+ЕlgWi"z(������
M���������3T{��	so&0&��ၱ>V˕�`(>�C���OM�9aa� 5\���:p掝�Td�3V��@�˔�$�.�c��	Ŷ�	�&D9)Q
&�=�$�ƶh�x�B��R���b���Bjm���Z��8�'"(�1-�(Z�x�Pg�u�FA�����)�j�8i@��A�Hز Xe�b�t�����'HW�(!qO��Q#&5E��"0`L4P����,�?u��ɚl��T�� H�;b�D�N�ܫ*��	
�� q0ȰWI�2#i��\|�L��Tв�8��?�; .B��i�Q���%�� ɐ��?e���X=ة����F0�O��c�C.�'��-�2�X�䏙D!-��Cl��`j�E���0d����?s	BXp�;?� �F���`�Σ.�@��
��*��*�C�-R����ԩ!�	�'7H�w��~�I��R�@#k��ZJ{g��#F-�T�� �+t2f���7&�9`Ъ^���DZ&�\q1D�D���nZf� p-�=M����o]#��4cR�<�G��5|�Ӛ��ʎ��'lZXxv��d�j�����\�~(�Ů����$9z1����L	�^�D�4*@�B�r�µ̉X��1&�A�#u��%�����?�Ӻ3"�Q�ؿ+ ��V#
�Z��)V �K��֌�8L#���!`N�h�v�&?�� N�~��E1k8fITŒ77$�c̧/vj"=�׫�X;� ���*���\3H
ņ��9/(q�/&g��()�(��dȹ�sb�0CtAr6c�����!����>���`(:xp�!�#3u>���צ��T%KF&8�/?�� �:y��~�Ri�Ïڍ|���Ye`��|! H�y>V�0%Ƽf�er|� �i:O���A&vɩ爌�hQ��r5KO?�~ 
� �$�1̇˟`�^��.�>Ma�� G�\�i0=��O�W#N�#S��/��=y��Ev���`ǡE���Z�鐪W�~����rqj�R�D\�U�x�'  +��?�i��p%�>9��8*`19�C� OH����m�'�~<) e7@8���I|:� �FO���Nɗ���)c�V76 �a�l��/m�}k��_�r6hDsg0O�V`� E��H���
1�< B��i@MR$`�;k���O�n� 3�I���*qO<@��
 �p yE	Y�@c��a��U�" �6��Pxbh˪IH,�b�U)E��D�O����5g��hir��$V�*�0�m�d�\���f�L`AW?	��ܯ>+� �IN�x:��2�O*��F��K9ذh��2��9#�Ηy2Y5��R��(�a�b��}��/���ȑ(I~�L<���]X<�j Ň/J�ڈ����P�'(� 83��_�b?��Wȝ#�݈��وb
Dى��*D���u��*k9����ƌ�k^X)�h.D��Z�B�`�����>� �F#.D�쉴"��q����#a���8��Չ-D��L*i��h�#I�"���0D���4�[�07J�s��3�訐�-D�(���v,0�W��9��4��/.D��E��m5"}[V獱8Ȍ$�t�,D��K�lA���Ч�.Kl���`)D��3G�Nnr� �mE�T�|���$(D�����(�P�i�őQ���� <D� �������T℈A��pp �6D�Xە�[y@��a�%ǲ#��x�8D���&�TCX�g-W�
r���$D�t󔆞������,qW����'D��9��ٗO�Ѐ%om�hr")%D�0أ��v�y��Vۜ�*�.D��Y �ĳ��K��W�����2D�H�ac�N��-AP�-;��A�0D�HA"�K3����-^�f(P'�1D����.)��qr���9<��`2D���CJ��AX�j�VQP0e//D��X�e���u
�I�+w$�R$-D�� �� A�x�
�[q�˶.�60��"O�*Q�Yd�T��a� t2��"O0����*6b�+�O��D��"O��P���@�b�c" �w@z�"O�P�D^�X�޼ o�m�:�"ONtR��;Z���J?E�(d"O2ذ��9;��1�\R���V�9�yb�!�B���^02��Vn��yB`�(mK��@G�X��r�`�y�O��ण�[�P^�D�p�E�yRg@�;Θ��N͜����Q�yr���ry*�ʲ�^W ��r
C1�y�I�>4l��PB��Sgez�b�!�yRM0y�M�b	�B-��q�����y���p��H��i�*(�zH��@��y��Ϙr�@�`BH���d*����y�G�,�Ѝppd����wd<�y���C���$M�\p�`W�M(�y��
-mm*2MW�}(�T��y"%�ܞ�:�(��Kچ�*�E�y"lM)T��]��f�A$"��P�8�yR��+�x�[��Ա/
�9�ǌ��y"F_� n�,��fܟw�ڐrr�@��yr˹2��}��D$^��b����y��=�T���ɛR���$���yOW�R\4X��H�H��pAaJ��y�����(���;G�@��p)�>�yb���V���F���2�Y��y�%��Ni��ˈ@�P`#���)�yri�4$R�@B,;�n�����y�h�=�TQ�C�_�p���@�/�y��Q�=�����O���9�o�!�yB��97b�	F%P%p'�� �M[�y��ܸ��ؗ�ˡh݂��	���yR��19�DtB��Zc��B�C��Py���*M
V��!�,^��}A,DG�<�ƌ�Hg���.yl�`r'͚C�<�EK�M��R��Q���"�mk�<�@ڴ\�b`K<��d�։�d�<�S���m���t)D��$�x�G�]�<���9\�t�!�.&� ����_�<AS/����ʡ]�V�IY�<3���T�B��Bb?��*a�PS�<��i1Kh��fK�b_��"�k�N��G{��Q�w���b��Ip���y2�z��ؓ#@&	W(t	�F
�y��B�Fhd��N�,��8���?ؐx⩑�-�b��bʒ*)t��3��&�C��=V�T�1iQ7� �ˡ��3Hi�C�	*fY���*)n��iPoڜ�>C�I[�f�HuiP�p�d ��I�,��>�t��xaA-P?g=zip2�g�45��^���d��9{��xFa2z�:U�'�ў"}�`��!H��O�^���Ji8���H��8� �n�敠�	-OP����4D���C ��%L @1�F43�~0Z2C(ʓJ��ʧ�t}2&։ZJ5;�O�'��L��*B,2g�Yf�r�L�?jڈD��H6^�⇏�(*3�Z"�K�j�������QÎ9O��� �B�4"~�ɇȓo:�)��ˈ(��8�$�X�'0x�ȓR?��1D�۟9�H�1|_����E�.d0�V�4���4���vG�}����-�c�͆:���-�9U^ze��S�? ,p���U ��VM)[�Z�+C"O�RT˳R<TxW,~ײ�(�"O<՘�ᙏz�8��� #Ǝ��"O>�S���0*���Z0�[T��qE"OpL�baܧ,��U�3e]SZI��"OP���'_.k:`����H;Ix��"O��b�d	RVP�S�/��䀓"Oe�� N�$�����b҆.�9��xr�'M��`
5���Ap'��
imI�'v ��e���l#a �|��\Q
�'ib9�bΗkx�C��ɬI���Ǔ�HOd�iBb�<H(�I�(��e�ʵ�$"OZ��3�g*e��,E<Bm�E"O�8��+#<p"	(M�D���"O04[��+T��Mq���4�����"Ov��3uи�+#ã ��1B�"O�uJ�BD"`�H�����.=���"O��c	�yf��M6��(�"ON�[B-L�E���@IԶ0͋�D5�S�S"��Q
rOҐ)�$UY��^ sm�B�	�S�f�@6��G�lħ 	��B�h]�9�g]Q���Q�ʎgz�B䉶O�>i��Wy�.����D�Eu�B�	6D
ݫ�I�������U�S�TB�	!l��p�s]�� N�R�FB䉔zU�8Ջ�)6ح�1�%4E6-%��1�F�s~���ܛx���t=�O��	�lP�I�A��&0���c@�Y3�C��1nG��"���%OT�(V@^�QAZ�<I��T>��Hm�B�&#I�u�Z�8D�d�e*�8,���"�}��SF�5��hO�S��������fGN!+֒B�s&4�-L�> R����%ڎB�)O�y*˕ r��)�ᗶM�^B��|��a����/q��ıV��zLxB�	��}�����\�"�l�K�2D����a�O%Zy���D�t�6�0D�8�V��s�X�'���?!8��.D�Ȉpi��y���e.������)D� ��ٷ`�dbŏD��pj1b%�I~���'0��ҧ�0iH��i�$Z8����g̼���۬3���qG�4	
V�Ex�'6rX)���X0��3�悉J�p$�
�'�L\Q�D0T���y�NϚAQ��i
�'�j��v��p���QC�ț���
�'rX��?peP�L�B,P:
�'�P�qO��x8Д������J�����%f_4���/
��5�G��FG|B�	�w�Z�� l�=���Ѓ�ݕZ^d��p?���q�t�{s��"UH�YK�<��
2�����!}�N�ۅȁq�<9#-%-L�;7�
2���)�,s�<�v�&gU�(�cr��Q�g+Vp�<��F>b͋&�	E���gΟn�<a��7��iр!=^�d�`gm�<Rn�Tn���iM�Rvd��[n�<Q �LjPT��e��	:q��UP����>!!cdh�J��3�i����c�<�a !U���"�℁	=���3N�c�<i1MM�r���S`� "��Q��KE^�<y�	�-7�Z��V'M�yCX$h�!�t�<��SL����t�S�E:�8���p�<�#���}1Ո	�)N����k�<���/?,UZ�l�4+�dp����j�<� ��;����|m�l CK�9:�9C"Oh�Ѱ��0�܁��dV�.=���"O��0���v���Y �
�N���"Ovd��R�>ό�ԃ��i``��"O>�b�lX�[d)�U�]t�t�S�"O�QvEE���`�GYL�"O0m���\_b`p+N?E6�&"O��xw��hi�����N�j�x���"O�e�`�ύi* ���]��q"O����W#�R�" �iA�dYF"O��:A.�02wx�3+2<�Tc�"O���S9X{�[�'nЪr"O�h��*��'њ=ɑ�� >Q۳"O�����K�Xa87bV yV��x��'��ة7c�V\�+�ǔ4��
�'0��`�w!ԵA�n����(#
�'������xe��a'ݛ����
�'/|�!��6:d`�	'��
�'�(���;^������Z6C����'E�)����y��b�샲{4�Lx�'Qԭ�#��e� �;E�p�N- �'��p�D���8���
p��3=u����'���)2�� %  `n[�2�@���'"&�Q��&게;�k�&T�s��D(�'``��!
�����*W伇���5�EfE�N����(%�Z��ȓ���4�V.�����p�x��ȓ9D^�.9԰�1��&����Sf.D�8�`���.=�m��d^�}z[��*D�c�鄥L�┉&��nP�t���*D��+ �ѡ:��X�3�R�K>|�r�E4D�J�ưB�Ό��*�{J�Q��0D�`9��"~4��(���.`q����q�S�O:�=���Ԑ��!�Vc�.9�	�'��<�!�_ò@@�'� f�` �'��pp�� W��
G�>����'(噑"�2(�ĭ(��:/�$�'�Lq�L�K*KuG�%��Q�'3䉩"j�%4�(�c$��W���'�$x1/�}��0p�h S��h	�����Է^ B�s���3 T��j>D�@���ޞA���ڔa׽�,��#>D�lW�u0d�(Pk�d��"D�Tqq�|-
l:7i�f����}�<��̘ F噢��.cl�iP���N�<�2�٘v۸��a4ez`@��G�<��HX4*X���6�jP�T,�k�<��C��&7�|`%l(7�ҝ
0��d�<���E *��T!M%lH�#��l�<�ă0�ÑE��6�4)�Ch�<ɣ���(������Թ����e#�N�<I��V3H� )#f��I �`S�d�<����EJ�A ʈ O��)*��_�<�GJB�]�0y�u��L5���d�U�<9��C'j���!U�R����L�<A�M�*�|+��-��=�b*I�<�f��|�����*m�eBD�<i� GH�4��a�%cv@��w�<a�
՘/Y&��q�$l�h'oCx�<���?��(0�� #;�]��v�<��U��p˱n� >�A��l�t�<9��K���H���Nd��Jp�<���������Ot�tl�@�<�1��<"qH�M�*�~��aW~�<� &a�WJ�-9�,���J!lHR�"O<Q���3�rP��.MZH��"O�<���9B�p\���-`�X�"Op�S"�:pt\"1��;(�|5;�"O؄���>�D�+��ʋwGv� �"O 	"@��7�<�kx�0�3�"O
	C#λb#�Y�$@�g�ց8"O2�`�
.+��;S�.�*�"O P�W�ǣ,�܌�c,m���
"O�b/j-��ം[�@�D�
a"O(@�&�2� A����&tZ<l	"Oԁ�A��>ˀ,g@ڕ7K�$��"OXA@ԮKD �9w�/;V2Ёb"O��"Ŭ �2���ǃ}fj0��"OL9��!	 !�6�!�`ȴfg2��"O��	�oոō��5��4+��(�"O��AA�TP
�eS#.l�ܹ�P"O�$c2��3G~�	�
/H�͢�"Olt!�L]�y�ڐ����W^j"O(�E
 "tLfLz�@�/L�8��'"O��4�C>S�`M��4�rm�"O��)5��	֥�����jM:�"Or�g�4a�����Msxe��"O�q���O~ŃrBRBqR��"O��sǏ�}>��0+Yom�0#"O�4�	@�TF�xp*�7
O��"Oz(�A
EP`z�(I&	����"O~�XrA2HQ�C��43|T��#"O��Q$iI�[��q �)z�Ѥ"Om�a�=e�d�5f�M@��@�"O��!p��SS��.- t��"O2��T��0[&Ѱ"dV�g!����"O }�Z�}�t�S���}y
���"O�)�&�)�r�CĄ��d"O��e)O�S���q�bA.Zn�a�"O�i������B=:�T�+]2��r"Oz�r����%��&��+&RKҬ�yj�X�~�$�_�l�V}z���y�(�
��8Q��(d��H�#���y�D����C�IA�/�)k�cH��yR�E(l���`���!��h�P�K�y�6Qsm��/,fc�1X�Ʋ�yb�מ:��V	��i���#@	޳�yrė��=�1�\ a����Q��y�,�AeH���GU�@P6��(�y�܊2�T��t��L��q��o��y���
F��ڒ%W�(j��D��y�C��:D8Gb��	W��0VLX�yb�݉Eꈠ�A�4�ċ����y�/ǏR�T��bؾ5,Dyunȏ�y��&Q���*--�d�12a�<�y2g*5K���tc@�(d�J ���y� ��c+��)ѫ�%`��LV6�y�*��OT	��N5ʤ���l��y���5<3&���č_�8�B���yRc?x�M뤆���`���<�y�
�,�^�@@�־8T48�ƌ��y�Χc���`��rp����y���=�����ƣ��GPB��ȓM($���Րfb��[R)Xz��	��U��h��K#��L�"�DB��M�ȓh7���b���}ism�V���ȓ[�h��l[j
�z�Җ���ȓ	e5{��WZ��5iܷc{.T��S�? ���ШA�<��	�ãU�~�pm�"O�E���1R$z1��N,�By�"O���g�m����5���� ��"O��9����Yr�O.
�v���"O4�sD���xl�q �fN�dn:9!�"O�8�kE�bHAz�P%(˔��"OJ!��GX�H��	��J+a!�A�"O*2�'�!p?���FiBx�� i"O����Q�D����uJ���"O��b�Ϗ�^�(��f�ʽ"5>�(�"Ob��%��x���S+#���"OؐCa�̶$-��@�W�,�%"O�9P��ضJD�B3j�[��uk�"OƘ��l�N���Be陠4��g"O����� �e1'�Οz���	�"O2Qi'�C�
M�
���:V�`�ٴ"O�`2����*]��M��bt�"O⥛�c��b�l ��q�v"O�YÒ���I
���$�J,T��up�"O��w�@�@���D���,+�"O*=8Q�M�$ 2|cֈ	�s�eP�"O�$x��au4���Ǒ,U�"O�mq���#x�.,PrhˢeG¹с"O��p
�k�R�)
D.*ps"OBhq�ݳj��u��C�'qq�x�R"O2 ��%�3������mWި��"O��­�-Vw�9yr#\3'*��v"Of���;���R 	.]	rD�V"O����?>�]����; J�"OZ԰���"jD:�iT��0a��Y�"O\H��m�V+<i�CB�7ӀѢ&"O��b�w��yŎ��@*�|�"O,��`cZ�=t��7w���F"Oص���9�D�%j2�ig"O\��3.L�=��eQG�qB2%�B"O����Ҽ�H�����
&�����"OR� a
Ȉ���*��Ƒ� 9��"OZ�cP�[}rX[a)ĥPf��;�"ON�+7���'�����/u`��!�"O)�C�
:�b��%XNL�	�"O&`��&�S.4�Pj,+�j͉�"O�Pq��#*vvuB�E%��'"O��Ԁ�&��!*Q呆:$�*�"O���%�$pR����IB<X�"O��qgə'���g�B�u+��2�"O|�.5i�%�7MX%.�"��Y�y©�m���
3��-�2�%�:�yr��W� �B#��(I,�p�5�y�j�?!�����I�PL5����y�"� =��|���ɶE�`<�g���y�g�!'Q���3	/H�F|qUN��y�A�f�����'�v��+�E�)�y"��`2D�K����CENi������Py"�_�-�%�E�/��c#�<ن(Y.#���£'uv�0!�eEy�<�'��IլY�v�%f���停w�<��%�<Kop@d�h븴���B~�<a�B�4�E(#�E^��yԠU�<����a�fmk!��f� 5��N�<y`��g�@��F�P���� �q�<��ӿI���G�g�� j�<	 U�t*��x�
e�<�c��Q�T	����E��K5�_�<ɶ�A�q����9?2Qh�T�<� 4u���B,Y0��tl����)�"O����f҈Jm<p�-�5�ƴS�"Ob�L�3�b��0����"ON0av��,�2A:���w�Zx�r"O��*V��ܥ��d�2�z�y�"OT���#�����y��ؾ2�>�H�"O���ׇ��g����;Q���b�"O�9'dܑG��F�;oĈ)"OyS�fM������p����"O^���[�B�X}�v�<�(9�"O�Y����	\PQJơX�us��q"OD)��I"xR��N�.IT�x�V"O>9�wO��u,2�Y�ңq7�*�"OЫ3a�
hq��F��,'IY"O��	�f1��%Ӹ06D�"O�9��\t6J�Q%_�F$Z0�"O:�j��^�PdX��Y �F}�"O`|
eT�;�`t A�� P��q*�"O4���ʛ(C�-rK�"9vr�*P"OȰ�M�2\��j[�u
Ab�"O2(!R��$`�\��
%)cP��"O��fAL)]���w�^�sx��F"O*����"~�: iVh��z|��)�"O���ʋx�͒4H[V� Q:u"O��R�
B�,� ���L�Rc"Oͪƾ6�|ڷ��%y�l���"O���"S&�f4b��S�[~�!��"O�Ic NX3�h1�Kȉ3l���"O,���j�us���2T�D��"O��H�{�NC��˹"Vq�3"O�PQ�N_�r�D��!Ɖug���"O,�2����XbB�0Vʒ6J�iJ�"O �x҅�{��(i�FԱL#��[�"OD1���?Z�\��K\�`z�[�"OJahv��Nb\b�C1��x"O���� �x���(�dP*f�Us"OlxTiB�B�օa4AJ*P��!"O���A�#Vh3Df�X��"O`���fY����Ǖ*DL��"O���c��NK�LHTf�/^�F��s"O sW�ɂp߾1���79��¢"O�$: �~�`��c���y��"O<أpƜ�-E���ł�?M��\�"O�P��k��(�hO���"Ot��� _� ��@�N<���'"Of��K*>��4���H3\:x��1"OPh�ᔚo�̐��(ў/���+6"O�x@�ʴ�\��G�5�^���"O<�!�AȰ7{Z8�s$�v�E�"O
���@�}Ἱ*Xa�D��"�y����J�f`1� G!*Ʊ�VI��yb(�
�L�@�>���i��,�yb�,_�|x��Y58�m_�y��߭2��1��&�����5�y� ��(��ʰ���f�	a�B��y��8�>�V�������$X��y�E�! ��9Y�&��CG�tR�N�yBMT�ۅA�7-�E2�P��y�bY�b3�MA͆6��dH$EX��y��0���ۃb�z���h3eY��y�A�/!\zQ"�B�h���9�`�0�yBbұM����f�b� djc��y�i=9�RyॆU���d\��y2�\86�T���) N�BD���)�y
� V�k%��?+��M�"ݤZ����%"Or�	6D��%� ��B��"O��秂)`j��L�7� C"O������I����G�N߂ب�"O�$i��N�bL��`[�Q�"Y �"Ov@K�iǬd��h%���F��-b#"O�]ye	]:f�`��c��*I쌔Q2"O � C��w�t����~1f���"O���bG8�Xy��ņa&䝡g"Of�"��ʏw�xy	�I� ����"O�t�"�TH<.�:�)�$rf �@"Oz�YTl��mL�q�ƈ�69��"O�sF�
�Ϭ�`����dH�"O� b4��T�x��C�0:j��w"O����bY�lk�#��Y��"O�xh2%܌�\�cÙ2^���"O��q`ㅣ;&J�	�C
 �`�"O���E��4YDH=aaRo��"O�p��o��/�p�����F��S"O�x`DH�C��
!�ϔ��d�@"O�Y1�e/4��0b���u��츅"O`
�e��M"��tMO���!2$"O�؃f�F'���AZ���L{�"ODL tތZ!�qr2k��Y٘�P"Ort;��ٔ��H�I�,��'"O^p�hI(VnҐk���3����"Oҥp���|映���E��ȉb"O4�	�F�k�4`*�݅|iN�Y�"O:ys�j�� `�*Ԫ�!]n�5�6"O���'�fe�X��Z4"O�y���?$�ɀ�a�f�!�"Ovu����8@S�R�V�ؽ�"O&9���N7�D�3�N�o�9�"O<�#F7�aA��Z"k@Ȋb"O�d
���92���Cah��A�T)Q"Omz �I�Hi�zs-.���"O�pP��Ca���%K�?g��U"OƙY��l||�s"J_�T����"O������{�tA�Gf[:qs�"O�8�g��t�.�p��,xJI"�"O~�q�.T>�%����6�,;�"OH��2�ۥ�(r��6<��e��"O�1�b�K�QA��z���S�@��"OV$��EQ1��3uC׎-ͱ�"O�D���\�LZ���6̔ �"O��E�J�\S�h3"�b���[1"O�5�a�)h&����| MI�"O��ʆ��~L�r��]	n�Zt�7"Oސa�ʨSr~<a�]�O
 �t"OD!`Ec��|��5�M�_��y��"O��J#k�Vx�^ GXmە"O}�O��Xd"����[Yz1� "O�P�F��b2�21%��S.�"O�Y���=|/��8�C�R���p"O�80h�vP�pD�I5H�X��"OzbŋL�`�<��B��O�౩T"O�$ �
C/bbBH���7 ��H��"O*�:�&߽y4�P� ���l�0"OhP0�=dVڔ����?[76P#&"O���-Dyv�r@
+3Q��B�"OpI���	��^e�`�=Dݲt"O��:F(��&*��҉��H("��"Oμ�w�ׯBՠ��B�<;���3"O�	��(S;SjMs%��1�X�"O� ���BBT:����촡"OfxH��C�g����fM�~ ؃"O�{w�R�dQ(�g��U��X�7"O�ɳ�	6~7"dce�?Ƞ�)�"OXI�h�J50T �]�X=kV"O"�P��*�QSN܈J�0}��"O쨺���J���gd^7�����`�%�`h�,\����	M��C剼_C���7m�gY���ԃC�X�C�I�ZB��WN�s�n�k��B��C䉜Vn�uhSI����Б7 �RO
B�I�Q�x˲䀑J�Z�x���<��C�	�c��-{�h˳:�*qn�,�pC�(_��0W, :���P����jA�B�	�-�^ ����$^h�� (7�B�	�"0��J�1W�8���Hٵ-*�C�I6)X�xҌ�=!ܬ�a��$��C��6p l�d�B'� �0J�8xC�C�+`C��ɕ�q����u�:c�LB�	�~]̅a����[ܔ�AB�
�L%!�.PĜ��%#E1yb����g!�d�4M�Q��R&�
�펰L5!�$0?�0�
a\�gk$�1��� �!�Ѹ&V��rh�
U�f�� ��9�!򤍖[��8j�� z� ����X�a�!�d����0{'�A�yԈ���G�!��?e�Y`ʄ���)90��m�!��>-�:9��h�*+La�Ւy�!�-V��x�E�5C,ٴ���k�!�Ѐl�Ь��� .�ɩ�J�a/!�D]�I�}R���wtɈ+;�!�����A��qP<�Q��1+�!�d�Zeӕn�)�T?/?!�Dđ ��Q �)'�p�1ܻI7!�?P�"���_�BU�xP�Ɣ �!�d��|ї�0Z�K��E�!��i�^܉pLR,ur��T�K�!���N�Kɫh��1��]�y�e��'������g��H�g�C%g�t���';:y��.6ֲ��֏`~��R�'@��!ƞ
,�p �F��Y�X���'+J���7k0ZukQW�p�'�V�Q"I�2_��%�T�T�|"�'�(�(�rlnD����p�a1	�'�$y0��A�i�3�G�{��y�'s"�X��X"h��Tbf@Кm�
	`�'�*��R��4*u��&û\����'^j����D$��Cŗ`�H5r�'&\ݱ@��:U�41��Y��}��'���	�7~%�P
�-NTd���'��yB S�r ��āGӮ��'1��k��&��1�Pf�EIB�'?�AYC��9��w�^��-s�'P@q�3��*
� )@7jĤ�'��`��N*5%���@m��/�*�C�'�lp4�ے5!��
��E�-�mr�'��{W���fi65�P�� ���
�'�8�#�N��4�  \�Ij��
�'[tI�(�iֱ��IC�����'	���FG2�x�i��3c^�P �'���Z�
î���vMEH�:���'���K�L���թĔ>�&���'���dG>��]��c��5�F���'�Hr��5�f�'�W�"���� �9!��'C���9ga��54jac�"O���C��)-�J�"�o$��"O�`ˣ(ǽ(�@�B ?	b�`"O8y%�����q��P4����"OZm���2%u�J��ʻ�0�CE"OjX0�0�,0��L��(J`"O"Q�!+�V�8�b��r.UKW"O��!���,�.�S�"�?�prw"O�uH�	\�kO�����?2�bT�V"Ob<a栐�y��H����8WI�T�"O�5��!�H��x��ǛAn}�"O�8;PDD�A��ۀ�\�IO`�Y�"O�C�[�q}xU@��ͯ� "OL �E#E��3������"O�}���� H:��e��J���`$"O��:�,q��Yk�/zxB���"O�9�i�p�δ�A�Y���"O2Y�&��X݁��#{llx�"O�!Y��@.֥��G�*S����g"O�ܚP�ƒ$g��	��b��r "OV��v�Q2��X��M�&�P�"�"O�ecՄ�>[�(���D&@��U�"O��bRM�d�(ܣu)�Q��%�"O�:Q�fM����Re�0��"O �'䙿=nhB�
�&��C"O:�`��,xP�<��fP�:�L�cQ"O�e�g��W�.�3 ����9S"O�iq���:(���V �rͨs"Ozp���i�)��fJ�����"O(\�ԡ_�H]b%�fBY�%Z�"O��P#�I?v��[���4���'�J� &ϊ�s���Y"��Ldz�'���w�K$6	,�pQE�����'�z}K��*��MI�
O�l%�'L�p�į��MW񩒇 �I����'�.u���[}d\)��>��]Y�'�JŊq`
���8�/I,I�`�C�'�8��B� 
2(s�(:��@1�'Q�$��_i*�P���-��D��'	$T2@�ɻt{fX� �_sR�!�
�'�
P����
ʠ�-�<AV�
�'�(����!E*�R�G k"�M�	�'^�)���M6az��°bX�j�x�0	�'�:��$]~5���p��1f�"�)	�'��-��Ȏu����*��V(�y�'�0pjANT�[1T�! �ɂH{~,P	�'$�$�Q�MG�<X�"��@p�e�''���!�B}h����`)&��ɱ�'餵��g�oPq#Nj�0���'�M�&ʘG !�!��9Pg�%H
�'$�d`�?F��Yk�/��A�T��
�'�P᎐m�׎�"4�<ݰ�'R��#��F���p���-��
�'HF��,��^��`�C�m "��	�'!v43$Ɯ�(b�ܺ0ɗ	d��<��'P0�F���3P�B�(L h�
�'s���`mP %��b G�12%�{
�'M
���\Z����wbK�rXH@i
�'��� �%{ �Y[�l	�?}�\
�']B�JvBN$G��S��2�>���'���� ,^*�rKӯù]�d�	�'��@cU�_ ex���	�OA��C
�'��ݪ��Ɍ\��qS��*I�d��'�xI�ʓܪܑ���p�,�(	��� ��BtmU����y���2*�~A�p"O a�gR�m�(���T.�:��`"O�H�C��54]��(ԓ2�TYX"O���6�	)GJ����U�Tx̡�p"O�DXU�	Z���Y�p�ܠ�"O�c�:�*ʘ;Nh8�t"O��"@皫W�����A�`�h��"O �cKͱ]4��VN<9G��J�"O&y�Ԋ��P � �^/�`r�"O�}%��TP$Hт�QW0����"ORL(`ߗ>����X-ڽI�"O��+Qm��:��ڴC�> I�"O*(���e�\US%�ߝ3�Y0"O�Q��ȼ�����@��ޅ�"O���!@E�#v�a��;E�@m�"O�c���5dbR�]��AXU"O��5" �?<��f���Լ��"O0�i���h0�s�+� aPIC"OT���葴 [J$ieJ�]}��K�"O�csω�M��+[��� ��"O2m�����hz&�M9Uy` ��"O"�Y�E]�t�
�
s��Tn��W"O�p���̯ O��4M04��@"O^����,�^d�� $`�k�"O��X�=&}�Ջv��pT�W"O����GL`�Z��8B�R8�!�$V�(~�q�s/I:i����K�\T!�� L+�E1�I��a���'�'"B!�$�	�͓�H�;�d�C��70�!�d܃p9��Q$U�yͦ��JÒh�!��V85q�<{��mOn+�/�$�!�dE|����eI[F��Ķ!���6��T���$��`�*_;s�!�$M:3۠ŀ�상G{��pt�V68R!��5>�^�a����%]�y@��*;!�$#���S��M���Q	�=s!�$�`�rqJؔ#*b`	��̎P!�$N?	���B\d�\�� ��p�!��
On���G�B�^B��bt�Z#|!�����2��2V� 9����?!�dR&��t���3StPX�!򄚕9�-�7m/{)"q��AK�7�!���j�f ��� �1n��U�؂.�!�D��3�D\�1
��3���1Q�!�Jb^(�nX"3�.h�$ G<w�!���9ٔ�1e=
h���[�D !���"dʄ��l�Uv.=xGC�!��:t�԰�'�IsmK���C�!�$X<zIKD&0`,+�k��,S!���XG���GGL���I�cE!�d�rʀ�qbӶ�ވCD�B�i7!�D6A����ʒ*�����O&}�!�D�U���b���a�XmpхM�l�!�$�"j`��M,!}����[*�!�䇴P'L������ug�8	���!�E�8�z�1�II�O>d��%�$�!�$�!9<$L��-<j��5ӳ�!�dC�zg�Л�g�? 8-�O�*�!���E��˗=�p=µ��8{!���n��U`�?f�V�ZŬpg!�$XL�eZ�l��G�`,RK]`_!�Ğ�A��0ڳ� �jp�V�תV4!��Ф4���Z�O͍G�z�h��Ş]�!��Y�u����F���A�!���!�� \iH@�ƛj�����n�3c�(�"O
9�1H��$����m�Ȑ��E"Or�SA���K!ı���ܗ�H�i�"O�ɉ�K[X:����6u�� "O\�Ѓ!��o���2EO�Cp�̹T"OVH#�K�`�D�:#o`5��"O��BRJRb����� ~ä�Jp"O�½IC�T�T!����"O�1�k�2C1x�[���Y���[C"Oj�C��πt���aMA ���k�"O��qcf��r"N0�c)� A���H "O�Բ�񼔲��5��e�S"O��Kd�Bn~q&ξh.h�j"O�A�W�ڭJ��T�?cΖY��"O�=�����%v���h�0<��G"D�,A �^�zr�AjB��y� TH%I>D�,��cW�U ��JC�:ob��Q�
=D�,���2G�
U��瞏I�	�E/D���S�
�%*�ʜ�6<��+D��Yg�P�Pqp���[�8{r���.D��Q�M�g��L��"֊ &pY�%A>D�4�%�2��a_*Z��M;D��1� �}�� !7�1��5�9D� �Fd�3?f�ⓨ(!B�ɲ��*D��s��Y���"A��h���8��#D���ri͘A�T�a *\5&�� -"D�<���]+H�A���F����A-D������r�0�E�����&D�8C�L�O`� �'ֈX"�i��$D�P�aЎq��2p(�)@0ҭ!�- D�<{0�Y*c ȝ�P���Q��Ad D�l0Q��Nt��C�A�j)�D>D��:O�K;칃�1q�Z��'D�l蒈H:w����5S���&D���0#V�R�B��$���.\	�`%D�p0X 9#^5�"F݊�dSM%D�8H�N�[��:�]�5��j'g#D���FHF>9�����f:B�2 �?D��ۆcA�b��c$M�H����>D��;�n
)\ҭ�w �!X�`u��:D��A��L,}xd�\�
�\��9D�� �Ѡy��w$/1h�B�7D��!�DA�!L�`!��4 08�D7D����ߐF�T0rs��>�!K
+D�����}��<ŕ|
~�zP,>D�����0[ذ����>wjA��.D�(
�/Kx$*y0fL:�X� :D���P��S�4(�0B�.Nez�ih8D�8�6�E�n5F���X�V߮�#�"<D�H�hVDX2��4���L+���"9D��g+�<-P���Ş�:�ҩ�a7D�xPR(��^��EHSmR�r�`Œ�
6D�l�@�I8"b�*�63T� �4D��3oj�hp)�m����O�yR�U$^qb�ib	M�4 X�9�y�&	�{NP� �ݤ<�.1�Ή�y*67Ş��c��8f6v�R��3�y���	v����k�3��h�v���yr� -!���ਚ�/4�PZC/P �y���3�p�^({
4�׏N��yR�E?y%h�2LI<o��[���)�y�.��|����Rc�`Px�:4EU��yb.�#6�D�y�e��\z� %�M��y�!�3�L�h��O�8�H@�y
� �����v�y�	�>6\6"OH�G-�?aL4��Ȉ�5-~@s�"O��ã�͘IT!A-�:6q����"O���E��R�Ō�I�&@r4�Җ�y"�DAV��5��E{�(��U��y"!R��*� F��	A�L����y.υ@��уi�6��\��X��y�]�B9��29��ը����y�	�
B$X<����aTv��QG��y�`C�s:"����X���H`J�y�`�!R�}P�']`�d��`��yR���g��QB�j�2Q��}y4�Y��y�X~܉��1=���t�L��yU�>��[F�^ "�\��J��y�/ܵP�����#��h#$���y�fT$s�D�!��X �TQвoM��yDSXi轸��3mt�"��2�y�bԲ@�t��%��7w���� ���ybd�O�(�����"���yr�֞J��V�HyĈ�E����y(T =檈CC>~�あ�3�y���=4bЁ�D?KZJ5��M��y�g]�q�$I�g�3`:!K���y�Ei�"ՠ�+�W*�92a!]�y��"p�<��L#�� ����9�y�EU%�dSf@�<!F^�#���y��"tz�ش��"�	IW��y2GD��,*g�� k�2)�憄��y" �)�,��`�Z� ��M��yb`�x~@UkBKҫQ���������yRa :���1�Q3�x�������y�F#�\w&Y��!�P�ҭ�y�*@�5Jޮf��G���ybkP�,cb��g��k�<A�5�ͣ�yR��8$��zo��,#��B��^��yr�E�ii�$��c�o�<!2��'�yk�~^����V|X�W.�:�y����i*��Y�gD�{��(��<�ybC�*78�l(E�Ыw�I����yR�Θ�L��Vbΐx�D�B@n��y�c֫py"ik�APg��Q�PhA!�ybA�{��Ey6�
��\�� Ч�yr䋱@<$Y���Vb�@U���y��ƔQ�R���+U@=AD�]��y�mD|/�ɨq Z�q��3��ʹ�yb��t�Ԍ� �T�|匭��.՝�y� K?n��!%DӒrv S����y���q�t�Ħ�	d�%c Ɍ��y��=;(��,�$:B�P@)E��y2�	�j�fU{��Ώ ����7��,�y�ФRP�3��O�{$�I{����yҮ�)<
���6kO��V�L��y"���_�������
enq��H-�y""ǱG���k��b=2q�S�7�y"�N�0���bGH�P�"��R���y��T�*޾����N'�8���̪�yAh$Qs��X��#�%�>�y ���t��e��n�Jv���y��ĸ
k�X��+
r<@<aE��yRD\G�z�*Є
p�Z��d��<�y��;�.�X�k؊E��AV��y�FD�Ar��f�Q_�4�cnE�yb�	MS�	XM �3$���y"�0	�e�U�G*DY��2a��y
� �◬��4au�S�;6Ԫ2"O�y�R�z<ƘR"2&
͡�"O:i���Ԕ-w�b���.���"OjɆƝ�<~J8��g��I˶"O�K%�ģA�=�f�=߲�
�"O���#X�N�Ȩ����, �6"OJy{󇜢2�2<Zv d�r�u"O�ň�KЧKm�M`�/��e� "OΌ�Go��б�������"Ov�[%c�'wy�LW$ 8G����"O�=�"�@�o���e�?.�D��"O,y�uʵq鬰�С�b)����"O�huA�
Z��Q�@�;G�\�!"O´����9I�,IP�*����"OR��&-ѓ\�L�Pv#�R�౳�"O(L�B� ,xK�]��/S:>׌��V"O5�'+�4ȑQ�߽T�t$�g"O��ChS a�DY���4�c"O�"��)u
�!�:���Xp"O"A@R����#��P�V0U�"O��A����Tz��7�ӸH&�8�V"O������10���-y,X�s"O2d���ݮJP6 kT-4KN4;�"O� Xeϔ�y뾍A��dfmb "O����bS>.p �bUB���8�"O��  Пu�����F�)�L��"O��k�'<���O�3 �2 �"O<��g�7I��X���W�9�,�s�"O���(D�&�:�Rv�ދ<���Q�"O\d�+�E���(U�LS����"O�e��
N�AM~H)���=
�>Yє"Oh��w��+r�ôĿH�ƹ��"O�]�E�W�?3��{�`�u�nD�A"O�QpCeQ�XT6�i��J/ ���s"O,��UfX�b��Y�BCI�茈�"O2u�v��?R����n	&��A�"O:��4N�C粙�%���z�6�"Ot�e�C3m
>������ �B"O�M�w��ҨX��E_�K+���0"O~�&�v����ړ!^�Pa"O�Px�@2}9v	���P���z�"O�e�2�D0G�)�c#ڥ^��A�"O~<�E�j�6����B�.עT:�"O�AJs���B�v����@��h�"O�@�s�	�b���#�D�{�PxB"O�c!��	u�X��1�Z�i��0@"O�L���P��8cF��-��T"Oӷ�n:Ni�g�-7���'{��KI�~T���1;�0��	�'����l�.LVD�J�:@ �j	�'���q��uT\\��B x ��'��1P֢��@B���ħI5��(��'APtc�)ԡ{p�����E�A�����'�b!���;`��<����+mh���'����O�8�8]+�X4 Ts�'����d�����j։��y��uB�'��ā�!>`�:��AMuq.���'�n�ʒdP!-��شȋ:m.�p�'J��
1 Y
�tŚ�Kfy����'�d��S��t!�"�Lb����'QpUc@�v�^ �!L�G5�Y�
�'n�`r�H�a��Sǃ�>y6J
�'M�i�m�;y�P*'�حj4��'	�<�CH, ]���F*R�w��8+��� ��а�lJ荂�Ӟ#w��;�"O�p2���p$�����@J���D"O�m*樃�(@�g]O��|�"ObE��c�<|�d�Ƌ��x��"O�II��_�3o��(��y���#�"O���������|3gႽO�҅�"O3PJ�09��sA�b�X� �"O�y�u��3,/�HCA�/x�*�1"O24�Vc�8(�(�q��)L�B@"O��Jչ����QL��	H0��"O℣���K<53t�_=:�sw"O8��hG�EԌ��3�ϻ74,}Cq"O4Q'Ș��"�E����P�"O���0.�2 \�2�
�`�A�q"O :��A�n4i��$āT/�|�"O��% [6:�����J��"OrEiċRj� ��v�@�TIpŒ�"O.�9 &W0Z6`1��>!Xt s�"O�HZa���S$)"WCC885�1"O�툆O
�h�V��2����"O��R�JW-)���2V�ڤ"Op!��>8?������J��2"O2�ʑ!T=ie����g�Q&4�`"OT$��ɸ<�݂�耖0�H�`v"O��BB�9���
uʉ ���"O��↩	}�$�� I�����"O"e[ �"{q���6�
�d�.I��"O���Q�'�y�ƭ�'F�r�G"O���an_)*�z���چ�8xW"O�K���Q{2If�q	D��V"O��a��7=o:�Pe��
H�L�Aq"OxI�J�!nQ#�
FU���v"O,1�$@�A�69i
�4>�F�j�"OtXs�B�\��%�CՒ�ҹq"O2raE�B�J`���R�@���[�"O ��[�- �B��	۷"OB;��
>@U!��+���y@"O��l��.[���w�P��T]H�"O:<�Rn��{HB�˭\��e@U"O�AKsE��p��M̈́I�H<b�"OF��猕$28h��\�W���B�"O�,i`��@��%�f!g��pX!������5�gh��Q
e,H�W�!� "����I���p����!��V#[�Ēc%�y	J3�D�!�?�R٣`�3a�;�+�\�!�Zr�@|x�^�X
fK��!��@�mC~\�!m�����S��!���@�7�>E��� F�#c!�d2?��0��V����0�9�!�$~���J+W/X����>|!�d�?9�ĝqr'P�FN��΅�~�!��ݠ}xᙁ ?R�|`�
�Za!�D].YPp)j2&J�{�Q&g��/�!�I� �
��B]J'e͏U�!�č�JyոI�B�R�*�$ 	!��B� XD�!}0�$��z�!�dW��,y��l|���{b\��!���0�ri�b�Õ
-&�k�N�)�!���4���SaT	dB0��gcʊ&3!�d��[���ZaK�Rx)���A�!�$�`m@��S$H5x��b3�R�Z�!�ΪE�6�e
Ź~���c�]�V/!���9Ԯ����(�oU�!�� ��cF�<1tt�"�(�����"Or�3&
� ����Z�O��0"O�M��2��+D_-~��"OHc���2P�0���ffHР�"O~��$�۾tʆq�T�^�, ���"OHHQ`�_�C�v���ǖ?���""O��)��I-�5�D��2S"OtE��Ĕh����E�}"ORX�j�9,�,�h0J� gԲ�{f*O�5ɤ��D`rh�t+a�<�
�'��PRD%��RX(�#�!�8D��t	�'xt��bb��y�ް��#+����'�De���M�=$��xEG�!�.u��' ���ӭڛq0�� ���H�' �Dɂː�K+� 8�H΁"����'��ͪ����F�����mC�'.��k� TƜE�J�Ina��'��,�e�	B�XY���\���Y��'Ax���ϙ:#����EF� ���'�|���~��Im.���
�'�(p)ׁ@)!,4�����`��	+
�'�Y�#k�*EE0�(7�=O@(e#
�'�) &v:$I����?��
�'���0m�!A��9&�
6ȸ�i�'��I@�#_2��bE�
�%X���	�'��y��c+0���oG! #.	�'њ�����{��Ըw�7(����'wΝ��޿�\�z�EZ6�x�'�u0��v(��1�)�
����'s�ͺ3��,O��ZG�
[�9��'��yH@�D�AH`Ey��L�z;H���'z4ك�BE�H= {�Q�&12��'!���B�6�0�C�Q6��'��Lʓ�R�j��;��D��@��'��w��ka��Y���)}:� �
�'a$%Sa��K'��#K{W���
�'��y��m��/�=��nA�C3j�Y
�'[�0���<�E�%�8���j	�'m:	�S�X.w(B�90�˾7w�Ċ�'����[\���/-e@��
�'�.I!�N�w�D��YGT�	��'X�M���a"���q)�7Jt
���'i�"#E�&�j�횎XL��	�'����s���H.�!ᜢT?���'�d�c��Y�g�)bǀMUf�	�'SB5P���i���O\	L�ڼ	�'Z�ӅA;F�*`�EB�E8ʥ��'��-B�b>ic����
�f�r�"O� ��D�����1f��a�Q"O&���Л6ު�⪍�h��s"O��I�'�5e�P��7/�ZI�"Oإ+SJ�=j!(�J ��p�q""Otр%�(5�	�SG'-�Ȥ��"O:�'���S�3��!a"O� �!�1k@,�T�_��a�S"O,1�3�K=�ر���^��%��"O�
�-�5YM֨�2��N�V|jf"O<��ĐkO�q���Ѽ��4�"O0,H����Q���
�g�pʼ-�"O$�i%/�6 =)E�^"�@᪲"O|5��ɟ�6�&�D�!~���"q"O���QcL�q�ᒷ�F��b"Obt[�BX>l�*�:1�"�|�y4"O�����g�L�����r� ���"O� �=���*_�؂j� >q��B�"O<9�(�V�Pia����i�q�"OF�t�E� �`��rb�>pz��"O޸8s�ё3
�(�>=j|�"O���h�t��� J,cE��Z�"OB�%�P�}��iu��>�!D"Oĝ����{�`i��:5*�Y�"O�9����#ۺ}I$L?�,�
"O�0+�%48`asE9��X�"OR-���ݐD������TwX��"OR�m� ������6j���"O����-%����k:}�e"OvT�!�:n�����o��"�"Ox�D$�,1��P�ɇ'L
B�(�"O�5"b��J�N��)y�LM�"O�`�'"Pjt�{s�O2ۮ���"O���)3@�TQV /�xTi "O6�Senąh���p"��I�Lk�"Ox9�7 HH`U�K�>���1�"O�%�� �:E�S2���!�����"O�\�2�O��
`�""ȶD�����"O�l�R-�A*��(�R�Ȧ"Oތx��P�8t �O<#R�P�"O �s芘|xlq�B���4"O24#���Kߦ`A�ɇc-&E�"O�$Ct��7V[t��P(ɫT���"OB�ԨȪBw&tbA������01"O����&K8�����=���"OB��m�-I��+�Dդ3��Y�f"O^X"�	R�w� �U��z7�d(S"O���ֆC,H�����e�*8i��"OD�9�lYIR�0"����pJܸ5"O(�3�.�|\�В��Y��ɻ"OȤ�7 ��B���P��(�,�f"O�<��I��-���p��[��ʕ"O0Q��7�
T{�"ϥ0\��S"O24 ��(v�1�r�W�p%��¢"Or �c�0�\� �V�F$�(k"O>�0����+	�ŀw����2"O�@�cO�H��t�-��$8�"OB��åmV<�`�.�WҊ��"O�u0��óg��}�@M�� ޸l8"O�!�V����QRŌ���'�,<��	N &��ـd\� ��
�'�6�C�� �x���.UT%j���'�f��sKݬ0� A�@��tL���'h�EA��$�PX��(~���(�'\�#���ej���!�Bi��'a�\
�־	
k��!2 �'��=[��)3�}0Jہ��A��'G�,�E��;,<�41�@�/��I	�'���%�7y�ss❛��0"�'�䥓$ɹT|>��(
||�
�'؄�@i�P>0�b�
4}
�`��'iL�����DԌ1�R��I=������'<����	��<W p7K0�n-i�'�t9�� [�|����֮H=*�4���'i�aIA!LB�d|sV�d"�'NX��MI�n���.T�d�l���'��f�C9vB��/�)_]���'�X{ƨ�"�]�ҥZ9&.dD��'��`���<A�8*��!��Ո�'� �Y��Ï@kj�j�����Q�'8��"��kcD�y��ƳyN��C�O���� �Ȓb`L�G �3g�I�*����'a��(�<xIT$�4R��B��%{��5��x�)&�P[����K̝����V۳A2D�`�o@r��5�O>��3!3��<�ONMY@O'F.}��L]�_���"�'�'��DH1 ��rA@S�H��dH�ǔ;)i!�d�6[r(�0X;3��'�#P!��W�3�zȠ��8�z�ht
U >!򤞃 L����8!rX�9%�K9���8�O��楐�9>���c�,��xP�"O��Q�$-QaD�[z�샢F�MH<y#%����1�L�sPVIq�K~��)�' ��P���\y��R�s{�\��E���@%L�dM�$�7�;c;$I�<I�J��˔K��#6T�aI�9}<��2�0	�kC" ۺL���_0y�Zȅ���	i���|��M,+1�H��tF��Ҏ(7u�B�R)�A�O6�%��.O_
�	d�Rc|�Xp�'�Ox�qD��Qj����#c��Js"O�9�t��E�/ژc^+(4֨��d��Ҋ��B`��7"�c!���i(Xȵ��)jī�N�8E*`��	S�i�V����@�~΄I;p��X;@Є�S���'����#�ѼM���>)ד�����`�#B��� Ǒ�j�Q'��F{J~����.���b��L���N�g�!�?D� �� kj�����Z�!�QM������O�]B��"�ˉ5#N!��
a��L���|��A��H��z��+ZɫD��� �<0�ǅa��Dl������)%	��Wr�����$�S��d�0��Q&�hY���b����hOj#<�C�[��<��	�.�r@�t�Bz���=Q�)Ԗ{Pj����(J��	��g�����H��)�i;�	B�H����"��!"��D1UW�C�-g��+�n�w�P��v�F�2|���������hO��Y���HCa���������T���D8��0�HJVeK�8�\�se�I�4 �Eyb�h��n��"maa��]Ya!�F)D��
�F�?\gyH�!I�������%�-�O��� E�i6�;pC�J� �{�"O���A���q��@DY(�z�"O�}�E�0��QH��]�e>���0�'Ӊ'��
�/��C��1�u�����`�	�'������L�X�k��*x�3�'�(u��Dbt�֭"��(�����<�R�&g4���nɻu-��x�����x�T�C "���(�l�TH3�枙�y��'���"F&ɼ@���&g̛�Z��㓹�<v��{0C�"�z�N�-�d툉��s�A1꒏P������Q"�4����0lO`�Pk5X�	��n���0u�'m���x"��u�J��Cd8I��ֿ�0=��^���'�r�@�0�T��T�Ժ[����q��?�'�F�
���?�f�pT 0H`T��{��\?���4�?Ma��I2vtc�e�&|c�X��3D���E�U*��ha�	'8��Ȳ�l�>����;FH�(���٫Q>Ȍ�e�)eO���D1}B��/Ie�b�>af^|��ư���p>Q���z�-���-%��h��o����?y@'w#�i�`�ށX�"=@���j�<�f�M�K�2��g�� �n��%e�<����pBؤ��e��<�¹h�BL`�<� 2�
���25)d�����5Ty�`��	[�(�'t�ΰ���=2�pq���g��e�ȓpd�ࣉ�84��a@G�G-VA�ȓ
���y �3� ס�(���ȓotR�� \�Ѝ;�5)��Ȅ�PS�KGo�-3��

��|/�!�ȓ.����R�����e�:5�D��'��~���;t��cQ�<�K!
�zx���T��O�� �x٢�I�E���h8$�#�@t6�QQ��_7������?�fK�}@]�.F'Q,���RJ�@�b�>!��˾t���E��04Х��F�<A$�1��@�)Åg��p��L�C�'�ўʧ?R����(�@�`%x$�qWv��ȓy�<��ي�~����>#A�ȓ{����gOY�����	�0~Fp��>�����L9_�T@v���oYX��\�n���F��BG$Y�'�ԩ6&������?�B/ %2��I�dڗhT�Z���J�<�t뛊%�S���5r��"�����Fx��O|�>����Ŝt��e
����+�Z���b��<��#ГL��-�ə�K[D�ڣ'��<9�4�O2�=���D��@�g�Zۖ��E�M�<�P���0U��@�D~�ݩq��Q}"�d&��?��a �u.�EX�*�� H�T�a�*�Ov�'�j�"�H=��E��.�h�' ў�}��ԩGR�;�hה%��;b[w�<�RMJf8�)���q��e�v�<ѤG�0j� *U��%iH�����\�<ѤĜ�Wh$M���!&&�k��B\�<�#�Aꢡ��V"A~��HQ[�<IW`ۃMtz	قV��Hj�k�U�<9��$t(� �`.��`��T�<yPb\4q�v��J&ؽ:�g�Q�<yw�X�y�8�Z5�2�{Pc�Q�<3��+/u�uK�R��1�%DO��l�O��	=�ε��`Q;r��Q��&�"C�NB�/��`k$�͏���oQ�VSBB�	#0lZE*bq�Ĩ�R�Q4B�I*1�v j��wA�a��
_�C�I9r�J�ޅk*�A�*_y��B�	�m��� �pQ0w�J�2C�	������� u���j��Y�tQ�B�I�s����%Ē]���1�X&!����x��i���DFU:r�J�{��C!;D��cǓ�_ބ���5c�Z�!@�%���hO6��Ь߯3��`�EC�	�x�q �"D�H3C
H�x@�����
Ucni(�$"�ē�O�e8����.����dK�Q��A"
O�6M�"{˞L�!�أ=@�%�2Ü�R�!��/,��I��#��)�)�bQY�Q�$F���ƎNPt���ו$fT��p�ۣ�y2F�v�dY��	��!�����$4�S�Oˢ�2�"�޼�` ڴ+���'��U�P�ށE��Qj�B���;O���ɫi4�!�R�`t�Xr�l��C�-���C�u�:�YZaBa*6"O�}AW�� nM�q�Wȋ�;DN�����Z�O��Y��¥�^ă� K?H�4�i�'���+�8$�p	S�i��=V��
��������+K�W�SSgMC!���eZ	
F�-g���#���S�!��5~.a�v�Ig�(�rjQ6j(!��(kްtQ��F���p�ư !�� n��@ �XsAcC1�"��A"Ov�Y�G�=\�<��mݸ�X�"O��!�K[�8���"�~�`��S"O:$��Y.��K�f�V�\�B"O�u��O����� K)R�Y�"O���vd��Q��!Jķ�.��e"O�K�*K�^tH�ɘ�`"O�� @տ=�1�D�&g�dyP"O�s(�/"�Hȱ1��p݀ah�"O<�
P��? {��5x��9�"O@9�Γ�: ��B,y-��ap"O,$��WX��sG9J�)u"Ob��1B�H�v t���_B�8��"O~a�FŨ.��a����/S�q�Q"O2�K��N�nŒ%{��SS" 
�"On�P������	�N�?.��He"Op j��΋2s���N�t�H2#"O|�3���O������-3��y�B"O�}�7��2U�����(<�"O@rb��䇒kR؝b�W6b�!�$���^i�!Gԋ5@���'��*�!�ĝ�Vdu℡�)w"Hx��,)f!�R�p���y��r Ђ�I!�d��^g�i�V�
� s,@+�S�!�DS�eQ!f�v�p��gV�>�!���'�8��P��3a䑍%�!�4���rT#�h�^,�A��T�!��ӣ:��9F�0����2 �/	�!��ޜs#g䅎l��#�$��!��3�4��`R0�k�B�4�!�D[ o��\a�d�J^�`Db��@N!�䋯N}���Ũ�$TK栊ς�e<!�D�uL̈����#L V�P7�/<�!�Ϻ#��<�����_/�Z�2{�!�d�&��r��A*�m�(:!�dI,U�v�!w!D(}픭9CL� �!�dI'j��`�śy9j�Kǈ]�!��>��DB��s>A4c��"j!�^�� �QP�]�f?t��0���!�DE"!�j(�B윅b)�����U �!��[�B\���� u#&��(%�!�4.�t�S������=��L=�!�Ğ*$Ab�[ul����bR�o�!�d�4r���A#��B�z�@� 	=U�!�D��F4��N$rWvQ9��!�dƩu�DJ�i�5H@�Q⮎�^�!�'a@>){�ϏB=��k��̕	!�$ҶH�4yh�3_.x�RJI R!�D7Z*��Q��'5e�5�EƑ�"�!�V;r,@�-P%��L�c��x�!�ɠ��i"-��Y���+vd��c�!�DQ%U�i���+&��}Y `�)<�!��8,}\�i�NľI�:���2=�!�d�-c/&�`������i�[�T�!��B2*EĴڲAE�������!��ա��U렄��%:Fhõ���8!��(p ^�9�ϗ �9�aK֙,!���,
W�%�!a�$�2�
��'!�ă�bu@��F���j�G�X�!�dڒ-����"��*� ����GU�!��;2�|Ibe1!|LI�֩�!�Ć9�,a�n \���S�D�!�$ߒ*Ƌߏ'.�PRlP*�!�$�2R�Nx�ti��l�Q���
�!�� �<��f��\x��)b	(�"@��"Obx�eEK$T1:�[�#^�(/
�a�"O�U;#��=b���kr>Q���R�"O���"Jm6I����h�9`��'.����{"���A�0{b��.�t�!�d�P��Q�<͊0VM��V	���z�	I0�ᓥ����b��,\˓&Y1o�C�I�IgȠZW���#4,L�
QM�xc�@��jВN��x��B�²`��,A�D�x��j��x�"� h�Ei� �6)ں�J�����Q)4�_U(<�6b��,�U�LA�H�	��A�h�ϓ�^cqOb�+v#M�H�P�S��m6xГf"OA�c'�� VC%��r.�qc���"����f�qO>-"��oxm���:���`�6D���@�"������[';�����6�	sn`��:���Z h��^�C�@�w`B�(& q�!�܇c6��@�H1/C�	.o��p�bAO�3�e��gB#cZC�I��B�r DEMi�5�-R�2C䉅	�i崰��������/D��5a¿ GT��@�8
Y�\�0D���"��9T����M�K���A.D���ԥ����I"�s�v s�3D�D�቗%�|#�䋘"�2T`�*D��K���
�81��(F�N���Z�$)D��%h[	Z�Y�g�X�W�07�3D��{�'��\�s�΅&_��	�S�.D���	
"��81��T-��!RB&/�)C����i �7��X��eD�Y��(�PY!�d�L������R#�ZxR`ֲ >�I�������>>4�`�B!-��ek�G��B�ɔ����C��7����	Y�Oh\K�Bƣ��<�S--p���3�P3P�i���u؟`�vG��%ծ8y�K�c�x�HFg�����Oht�`��b9��! �	C��	�z=���#R�D�Н9��צ�2�^�+n�$�=E�$EJ�wR�j�K F��$"�̏�G@�ɋ^--�U��Ӏ9$��Fa��}]XE`7ƙ�<���
�$�Ò��;1���Ipd ��5W����Ma�:�@B��D&�"F��D�'EXD���6R蕑�� ��Y���G9'C̝������"�'�ެ� ��)X���X�O�#r�0q��
T�ʄ��d�(Y����/!�)Q�DX��@3)�1-
�4���'a����"-IĠ"JZ�{�
h(�-�D�����D�+A�����@s۴4�+�O��*jڿz�` O?�d�zx@�j�OX�s8 P`FW&�ax�U:|� �{�A��1� !��'�th XJ��L��(���{�)�O�����-��u��P���������%.X�::ɉE����ɸa��� T�V�o�JĚtg�B$�Z��{���v��v��&KƵ��H5c���j�o �i��ɷ_@�w�A�O�T�F��3�m[qEՒ|�t�ԠN�m��1pS�еUT%�7�A6N	�L�6��]-�� �`B(^ Ĉc�삏{�.����.��"�퐬?��hB%.,5����A�T�
���)�"\��rC���4BE�-<�� ��Q/���'�.���IKh>��*�!#Ă�����N�'4��$�)_��,k6ꞽ�u�B� ֕�' ��.�����V�q*� ra{xm��/�j�n52����@�$�1�h��#�hbU�˻<���
���ձi�,i\��4,�뒟]ܤ�y��/,��)�XC���Ԅ�c����^�Q{�Q��	c96���;02�lP����hz� #�����#��v�|��&�|�Ό�?̽��+�<���'~�x(�פJ	��XT/�O���cB�G�e���i��s�ùy?�QH$�ږ"�"���/:"��W#[���]s�O7�1ؒ�6�֌h1�^�1�� �4�Сi���!�j9�!&�)�?����dD���g��F��s�A�<�X@h�>������	q9L$D�,JRp3�o#.���/�"-p�->{��pZ�܎�h�Har�S�$j���m�g9�	�ؐ%�&�+�ќݰ>IBK�s_���+&A?$ h��&���9�'x4ʡ�D[(�'�x���h���m5���cA�J�hl��@ӖF���I�P<�����Q~"��G�"�08�%�B}հWB��j�!rh@�Z\�'M��� 8���(Y�Un�,���C�[�������*���
%f�!M�2����K��E�,��`��=k0�yꕢF_.��ґ|��#���	.bm�a���ެ1�*�=t�&�I6AK�XH@Mm�r�s���.clQ?5�fMɛ&��Q �8�r �C�iԐ�y��*�Od�u��S�8ce՟e �]٧B�0]�4� %a��1SZ���]�x#�3�\L���l� J(��q��	cT����`^��EN�m��hŏ�$_�����Lhb��f��R�6i`�%�^�l�F�=3
d\
cm˕t�ͻs�?ړ~XH�!�����h��E�|���O��0֨O >����QÑ�"��u��'�^	�@(҄� ��Hb��	,���a��������գ%�V���G��L��ҏM�)���l�-ٮB�	������ ��F��y�/�1�<|�qO-@�J�*��+��Ai3K�|
���x���FV]� ��p)�}�l�r.�i؇�\�V���s�0���6Q>нQ����TH)�'�D���@fA9$���e)�Q���9S$�\IGc�_\a1��nW~���6e:�B�9?ި;`��d@
C�I'n���˥��nJF1��+�$$~��$
>]�"�6$���m�G�o���}��AV�J�fg�N�(�B���9�y�\���çiU�OItJu�&��kX9|�P����"P��(ʟ��["!�'&�y��"X���G'�OFX��^�
�xQ��X���#��U�G�ҵ�'�#N �����p>A���f  �t! U�xHz���[�'_�KV�.BXa��%fi�S�9�QI4�*p���x�;D/�B�I�x�����F�����*��қ!d���'6A� d�(W��9��|�O+��Ы�(G���G �0��$�'Lp8��'��`�ʖ�7�N���d:|�d@W�¬i7"�d�3�I�rJ����m�3d2������k@C�	�sH�Ż#FߠvS�Ѫ3�%`_�����<:a�z'�'�ĺT�Һ,=�y
3͆�%D,��uXx��F:��}�fYW�P*�D�Ё��g�!�D��x�j�K�A�`LJ=Auېgϡ���<Hϐm�\�~��=� `�f~�Z�LY6�x��Y�NMq� G�PɊ�.F
�0<)W��=J�BN>)%\�t��)�Ƣ�e��\��&�c�<��#�mא���.F"9�lhQJQvy����ꌃ�	i��ӰIv$-i1��: ���6�GR^�C䉓X_��(�'\�g��z�hB;~�)�M�D�hP�s�'?㞄���׾�9�Q��&f�Rii�i4�OB��edVr�.��s�Z�KPe+׈1��A
�9��?a 
�GoP�B�L�0�R�����_�'t�1��0P�H'>�لO��Ur�)`�S5��5k�+)D�<����Bx#�&�{�L�<���I�`�B�5}��� ƺa��O
7�h��%�=p�!�$�%V���#��K�j-y��:
�JT�O�jr��p:��qO*�DA�0��0��
�"�����'�.�rD�
7T\���[)d�~1"#��K��@��x؟hѓGV�y��� �Q1*ۨ���=O`���G�%���O�H��� �B� Ш��zC�k�"O.��S�u�^�� ��!Jjd2��>1�̓B����?=�ƥ���&}���
wô�&�Ӻ��ւZ$����������ch8�! �,�X��!���yb�6G>B �FҔp��+�K���~B�6���[v�'��3�R5(���Q�Y5g�=
�z̠ �ّ`�|�iǨ�t�B���X�p�2,&��z�<��a^�Йa�I���1��JMr�'�R�	�OB�`
�G�ԏ���KD_
J�f�#��D�y�K��ul$P0AH2M��!� �W�>t7GG �,�O?�ɉk��]�Mh�:��e�F4I��C��&�6p�W�u�U)��:`�ɀU�h� ��0��zrcZI�(��΂�+A�i�`�5�0>����״тam��n�4��7�	 �J�CEM݋:pp��ȓ���(�<� |s�AD���Dx�h^9fe��t�O�*��p'7[�6�x�@�DH)a	�'�l�:��S	ܠ�Rf�H���@P���pX6���M�l��s�� UjW��U7̡KH69���:#"O4���R$�Z	a�
�P�H�@�O q���H�U2\���	�e�8�&�Ɨ������!c�a}m�7C��5�I V�uS֤��k���A��9�C䉊�l��b��(PJ��iU�B�ɴ�h@�eK� �
�7�K�V��C�	;�83��8T��aC����`ƸC�ɔ$����͚�~8�M=IlC�	�S:}�D��Jm�)�u�Fm��C�	�;X��nU�������>j��B�ɯ9��`��#s�-����=#��C�J	�I`��yq� ��A�SF�C�	��fR�\	!ø����R��C��9t�2��R�`q���� �G��B�I�)�f��� Y�� S@�'��B�	�YҊ�	�CCpqXC�@U�t(�C�ɪ�Dx�sn��}[R��p��KΌB�	S�mУ�&"�|5k���)4J�B䉊sL�Ȩp36F�PflY�C�	)k�r!�����U+����HU��LB�I�uҬ�0&T���C�&`k�"O�<"��V'D2L�A%cǣ`����"O�(�hC>8�����O^v�¤"Odh��R�~��jPJϋ#E���p"O"yP�-].�D�1�=�� �"O��AH�:>�F����@��M��"O���Ҡ]m
HۣAv��i��"OVт�I��rc�\!$��5>���"O�̋1@L%Jg�z2��~�pa"O2tirb
Q����cmJ�C�"OA˗�5;�zw�)��ؘ�"O<-��I:L��5oƶ�4�"&"O Qn_�0�Z�h.n�ҙh�"O��ծ�&?�*���X����*2"O����#(W�R�PZ9p�x��"O���< � i��	�8X��"O�Ke��B���D`Ɯ��lb�"OH����'N��ya/�N�b�"O�����Dv��2��5))���"O��Hg�62��H�d�4N8X�"O���0�+Vt;���$�l�1"Oh���e�}z�T���.y�6"OFH��tV~�:��5L�D�E"O@u�fC�S9�aZ���+-T�]P "O�e��oT�F[�ԋ�eqG$M��"O��	P�ӞI���K�F�%���0"O��aC��8V��ڤ��4j�5"O�}�w��n� �L�x��(h�"O�݉�c)@�(�2����c���"O2��!��fh5��#Ƣ2r"O�Y��0\�B0AU���4��"O�1y��C@�*��ы#�TT�"O��F�C�Gٺ��d�E����xG"Of�B�:9~��$�L�@� H�2"OnRL�#OD���m�3c�씁�"O�  ����$�ҌcRq����2"Onxc��C��0�@bB�;����U"O� b$J���$�ڰ^�	J`"Ob��6d�(7��)i�Tq"O<��A������VDdA"O���Rf	 ��)��/gbN���"Ox����*ݪ,ðiD�Z��"O��K�g�t�4��7�ͳI&��"O��@�G��4�`ԢӦ�$Q��@�"O� �cp'�bذs�݆����"O��p&O�N��(�A@n��Lٴ"O�5S� Z�����N�w��9G"O���SC�3vqvp�g-U�43] E"OL���%E�_�L����^8H\��)�"Oh$���b��=��+�>ۄ��$"O6���3h����L�`Ŷ��"O�IЕW$�@��/,���t"OZ�w	K+o�xDAt�՞&^LK�"O�XBB�"����*���!�"OJ��q�U�X��i����^z��u"OZ<�Q�	M&�s�Oڲx�"Ok�K���!r1�e��D��'kX<�BN�O�j�Yb��^�*��'iT�����a0dR�,U�_ �[	�'�֜��h^t��lS��R����'L�}Hr�
1v�p`��.s�jy
�'��(��� &���r�"`�l��'� �����0�Fi��B�u�>q�'p��Y�H�Y.x�[C�^bf��'�Nt�A��}��	�U����<r�'C�)�B��-�r��6��C�'0��s�&'I�b�	�.�
w8��'�N$�dƒL��*�,�in5��'�2D���52��R(D�sN����'�ݓU튴^�H<��Y�o�X���'���g�>K%Z�iffuj%�
�'F.쫕$��G�j��fB'Aƾ,��'Ă��gD	l ��ѶI�5Dp����'����FMR�hH.vn��'�n���F�6�|`���Z�u�i��'�^-���E65ɢHم�|�i
�'�.ACdH�To@�*� NHe�	�'�>1��گ9!�T�G({��hx	�'ܐx��Əj�ѡ�ԍkrrd9�'+���C�H�&��8Ү^t�
�'}�UC�?>��`����@�
�'�$!�@M�XGt@�ebZ�VG���'�~ɛ�Ӏ �����3`:���'~3���aJt�	Q0������@0�1�)�'S4 ��l�F��T�N�{�
P�'����e���"$�[r/���O6 �eT [ܠ���>&�qP�A*dMK�l\�f��|"m��rF�-R��	<X�����D�P8ʸ�E
�e�b���2OH4S�SBRU�qnYm���Ey��6E\0KT��Z�O�H(�r��&�����;J��}��'%x����_%<�$A�:����Eʛ�>K����R3M:ԥO�\���`� `��yҧ�*A�Dȓ����\z�`	��0<"�nшX�g��N�%��`-n���Ɏ� ��#���C��5�Ns,�w(�+]���dN! �y2c��*���y��Ppj�ɝ.�X�'I�BP̵�#�ȡG���%�eag&��"��<Y�n�9H �,\�Wkƅ3�"O�MI�L�%t��i֋ًvI����]�Ðp"g�f���(7�ы{�e1L	'v��OZ�ۘw#h�C%!I5� ��k�(j;z�x��&f$�����e7��O�?a�&eSvl�${���IF�P#-�6�#f�6d�A�W-f2)�r�S�b�"��0�2�^6cv����׸)x}��H ��z܂�pj˅\�\�m��	��]5&��pː�Y.6 ^5'��
Y�AKҪK����JS@U�p�ꭀ� �~Fz���ef�����F�Bg�5��
����2��av�_�)N��Z#����>IV��e��~��9c�4*26�����l��k�0�]�2�'n�T���(�����ȘqT��!�K/�z���8?i��I�E[3��i�a��Q2���$�9��|G,
hn�|�'Z'M��2j_�:�v����<N��̉"�M�!a�����*���Ӵ(�+�МH�F�r��On�I|��Ù(D�A�F�a��%�Z�@�`"��v1�%�K�.eҌ�	)L�6�a�Ɩ�m{B9���K�4ۮ�������In�m��OL�hv��8�c��>j.r��7S��CLѫ5������_R=��E�T� �8âOL�,D��ƩV�#�.Ѩ��N2)��$�2�mX���� X|2!y P�T/n�W�����N�rT��t���I]��z�K�}}�ǐ�J��`U�i��#WLǴ]d���^�@dt�8�9�f���'�8"
^4jC�H��0]��'��a�B�AN(�Oq�
X�c,�.� ��t��4'���$�	1r�X��n�yщO�2��s�?@<�CGÈ	~��	F���<v�'��!����J;C1ĵ��E]8%������<�Ǝs팜"��6}��	�K�8�# �}!p9:7cӨpň�
�?a~��7�`�;s�	x��M(A��n�'���j-�ϸ'���3��z@�T!l���`��'���'��"�#EZ�h���+��UP�n�i؟��j�-e~8�����x&Rtz��7Ol!ӓ	�e~̒O8�{5G���ށbR��}*�Y�"O����@"?&h�ť�{��R��>٦��;:����?��4 ]�8g|qӶ��%��!
 l,D�Xɕ��=D�Lm1��	}��)��(D��ه �"5�<��X61�h��''D����b^b� Cكhs,���"D��*�[�a7���7&ʮ:�2�a#D��3Ī���p�@�O=
R< ��)'D����N&r��eϊ+Un�l�'�"D�d@**TQZ1��"�M����1A#D�8#���Tb42���2xZf$�SC>D��i�[�
+���Qa�T ��o9D��jF�<g�f��!\�d�X�[3�4D���"C�3%��9�Z�t\��d3D�41 W�Y�JUC��y"$dv�2D��bDH3��tU�6��!1J-D���b[B�� �k4�f|�3�!D��	���o�q3���+t^���1D���a���`��`"l�s���!�,1D�`A���c7b���oJ���@ñ�3D��R�B�W��e��b��h3��3D�0�����l�A�5�z`�1s0D�l�s��T�V��w��WH��%.�ԩ��2L=���a�Ԇs۴ͪf �f�)��OE�F�M'�L%�Fk�	\� �'n.(Q4�I6[��'��p(�N�D�ĐQ���/V5�
�' ��f/1.rQ�b��	�A�(Oư�%��	"�,t N��|*s��<W����ƕ?m&t�NH�<��B�^D�%"&��|#p0UHÇ{,�i�J�X�ꑄ��g�k��Z�i}�xS���5E&E��ɔi��B�d��FY��ѥ�I/	�%��B2@��'El��p����Z��$�"d�}x���< 6
Qnӑ��'e���c��/D����vl�
E�M��U|ȃW� �4���J�F�*5�'�DD�0�_(8�OQ>��6�C&9r,�j�jOޤ��e=D����N�
|�4�6���_�a������/1!�����~�3�ɟ2଑#�'TM�"���g�R����_0��e��cR~�I �.tPI�bX/Z��U8�a��8��!��jM��1��$g�n]��,U�@C���H��
_\Ra/)R�°Ƨ8�.C�	A�%���(��ć�'���'Q�	���O�S��8�z�aG�K.�ՠP�zm�5���jr��sӌ�)����z�t�b�1�8�"O
�V	�S!Z�pe��
l��8��O^�*�B�*ynT���_�dn��j�m�<�S��	��a|�޳tH�q����L�9g��x��B�5^�<�:	�'���Pba�X>�RG��7T��}������t��!�(�T�K��*d ��AC����#�"OZ��/�N%<,A�Ԑ^������U�s�*���"���)��<9�Lݐi��]`GiͤW.����]�<1�铣Y��0`!A"-N%�� �<����
��4lOb��&@W�����ԏ�1r�]9�A�1�mK;[�LM� P�J�.��5V�C#G@Cby�d"O~�R�HT� �"pf�oHX�s��+p�n�(�� 6Q>Ų4�	fa(�ڥ��)�v�Z"e2D������<f:9Q�B�nP�B�PJR�[֣�T+�S��y��.F$��괠Ǯ������yZ.�@��
_3}���f��kn ��W���� �/��=)�̄�q�v�����V���"��tX�l�ed��hDR ��	���F��b���넨�yR��2IA|�6�\X`��A����y�I�A�h�S��U���q2�=�y"��� Y����a�AӢ=C�kD.�yb�_H���aW��C����'^��y�z�Պe��'>�`�&�
�y��͑J@HA¯K�5�&hb�����ybB�h\�kc���F�<I����y2��QY�"�`��*Yd+�/׉�y���
��`��-�I*���y��Y��DB�'M�aa�&�yRL.���?5b��Ή�y�K���օj�H� ��h�]��y��\�	ź(��f\����14�X7�y��3C�H��������M��yBF<:v%��̕P"�:�.�'�y�KZ8��$)�k7TYj}Q�"'�yB�I����&y��p�d���y͟:*R<�`�	8 H0��$�yr����R�.�T�8E�S���y��]�U��!�@PHxs���y���mj|z7KP�\��b,V �y��-O�0)��C�W���r�B(�y���%�dI�M.b K�HΉ�y��� �@
'c	!c�����y�`�$]�FD���G�@�!0*��y2�\
T�v���*�&&Z�
'@��yr�;*��h6�J�Ou�� �n�yB(�2��3lS;&!��B��y�a*"���rb�V�,���뷡���y�
�?���Kp��WFJ��C��y��#��숅�Ur��"�I^���D���#�P�O��ᓞK�!��NЅ��Q�QA� ��7M��d���࢜�j8(,էȟ��-+ҴX�e�y7�4�p��1pԺ2m�%*Q�I�0|�CK�>]6�K��;5�4�DE�&9�����E�x}�Y�*[4��)Y7������;$�T\"��̱A��q+�^�$)��R�Vg�	��'{{b��D�X�h����D�=�~e�'�@Y@SDO�<��;���(�7Uj,��(�Q�|���0e��ЊE�)��ەK$,K��Ág�$��Ga�4�� �<���.]�XФ`��G��qPE�]?�6%3�S�O������{����&HT�	aD��R����'`���=d����l�:��ȗ��#͜�'���O�=�|�I~���¥M`��@��KtBAʃ�i�P�ў�OC�P���V���M�BZ�BM>�����H�������0hb���gR�c��I��HOq�����Z]L9��C�_\���4�J)��� �Ī>E��ŝ�!R��σW0Ȁ�&�M\��I ��'��"���o`u QAP	H�qA�KΦ�ʫO�ɋ�M����p�}���[�?�����j��M�>���l���M��Dt�O��ت̈́�X��9^��u�n�����yr�Z~�)§l���&��$r���kA֗+�]���-��?��~�A�	��;� It9����m��'sR�<�
��uCC.V
!y"�<s�:Py��x��'��c�b?���G�2��Y�k�*GG�YIfB�>	�'��`�|0�}:���~y�B�	\c��k�I^��mP�̗�(Er��%F_�<a ʑ�U�a�t�[��,����3D`���t�_V�͹%�k�8K6O~���'6��p�� 528�� �0��@��S�? �� ���%{��j!���R~$ 9p"OV�@�
�i*�j_@��5"O)���S,TE���1ȃ�pF6e D"OH�ӥH4p~����&��x��"O���E�$��*Ĥ��dX"O�<Bd�Spf��e��V����"OHYq�.@X؎	s�ܐ&�l��!"Orp���̍Z�����[	w����&"O�h��ˎ=k�J�je EVHm�"O��z��oS؜�`��;
��B"O�%G�݉��h�P�5ft�I�"O ��B�X��M�5e��"On�� �H&�P�AF;pd���"O���h�~��C˞.�F�"O�x �䏤���RFiGV��H	 "O��qq�H�>D�j�-P����"O��(šD�J�&�d��_^4�5"O��@$,�:�
I�C-��\H���"O���c��:�\�R���14�xH�"Ozp	ׅ�!KݰlY��$�y�r"O�pp�GܙE���Y��J=��"O�A8�ƫA���S�nT�v��!�"Oʤ:5�
C�X`1������"O�Y��ӯ9+��xB�A'"�`� G"O"�:A� �b�PS/<���y�"O���։�H?��:�BL�*��8�F"O:�d��'0�A�a̎�*�06"O�q�g�B��5���k3���"O���&
�BJ��ʙ*6`A"O���䁅n���xfh��I�z!�o�<���L	ό��PJ~բ�@l�<�����"���M��\kn�B�aPh�<�Q)֑	pDR�M�U-�XB3��g�<g+�p֢�F��5�m�k�k�<�&���X@MNJ�`"�j�<1f��?rt���_[:$!p׉�h�<yӨ�&��Ě�ƖC  �v��h�< �V2��ŧ�-D���o�}�<�R�=$1�eТ�U*�H	s��|�<���M���� ��s�3g@�w�<�'&��;��w��5 ��D;���w�<o�;i�y*V�I�l����îp�<y4��p�Z 2��*:�\��s�<�w�
�T�q�<E���w�r�<��������ݏ5�\�+��Fj�<���ĉ~�~u	���x��!���f�<��cǔ#Y2�xp(�$f��SGgEJ�<��X3T��lp#-��m�щ�b
@�<!d��+�|��jB��g�Q�<�d�X�0�\Tz�L��z�6aQL�<�	ա@�b���a�=cήy6
H�<�R��Vް�)&MO:��f�WZ�<ѥ�]�]�I)�9kAN��TBCU�<k��"�^eZ�F��!3�@F�<	���L7�;4i��u���
�a�G�<�4LB�b�����_�D���
TG�<)!�� -�F @�ʇ�O��(���D�<1wbŹ#Zb��v.�-\�F��`D�<�D,�,���W�N�S�0��B��{�<����C�����ʄ��DCw�<�Š��9�ry�W�̃$fĽX׈�r�<y�'*`�Jբ�C�x�b�bE�<����,*�U)"�R(;%�V(C�<��#�;(
��vg�q�d�z�.�g�<� 0���Ƒ3��e׀�?4Đq "O����K*jf� 󳩕�|/���"O,�d�52Є�f�N�f��c"OTuƬ�5.�{�#�x�NlB�"O��Z��E))
L(��b��?� �;"O����+�d��U��d��y�6"O�Ȉ2k2t��h� �6LʹP�"O�<*ю�N���{/Ю8!����"OX���Q?�!w�@�1���f"O"�Qd���uǄ�+q�ڙȂ��"O�m��B��0�ɐEڤ+�u��"Ox8��2`�R`��A$M��)�d"O��2����Z0�!x��ݫ/v,�J�"O2E1 Ύ�Q�m�B.��Hr�!;""Oֵ����O��ht̜�>O<�"O�x�CA�?r��i���m�(�"O�� �R�{��B�H'�.�1r"O�av�4h��W@Ĝm����"O�0��#�9r����c�
\LLh�"O��cþG6$�Ӈ�k0���c"O�v@ڥ�v@(h6WLA�"Ol8��I����iQŦՃC�&��&"Op�k�K��'N
i������jTpR"O(�*��_��T�q�D�y�
�:�"O�$�檕5	��i �R�m��9�&"O���TAϯ?��ES1�D:1��l 2"O\��	�O|��Q��(ʀ���"Or9����SH�l��e������"OHIv�N�[Ƙ#�����0��"O.�@ �ČO��x��c 2ig�պ5"Ox���T΢����3x��22"O
|��c�_[�+���avV�3"OD�W�ǮA�X y2`> Y0�"O�QK1�N�BC tcT� �X<T��q"O����b��/���x@��)���"Ov-��gF*5��x"�G/a�Q��"O���� ��TpH�Q��<AZ:4"O8r���J��Q�GkD;;��p"O�q�o7I(�Iړꅀ(�T���"OP�C���(#_r�q � ]���	�"O�@˕�O����׬I' ԋ "O��W,�zL��&��gxP&"Ou�E��/T�,<�E� =��Q2"O$�kr��4#+�K��V%T^i�b"O�����Sl��k����ъ"O6�����;i\t1A�eF�m�f�c�"O0e�fN^��:�H�"�a���8�"O@eC����<iu#w{� *�"O�l��,�z�Pp�E��3y��B"O�mx�c���Q"b��%H��s"O�@%U�o���HЪ�3�� ��"O4���`��%6��y��M�/GT�q7"O�(R-�`}�&��@�c�"O|\r��.; ���
f�i�"ON�ㆌϤH� �zb^�.���"OԙS3��[����A�zF�c"O"��ц��l�(ba	0&�Q�"O����i>���7��[<�K"O>�����$��lsb� v�� @D"O�q��++Y���NyҔ��"Oj ӱN�$Ӻ��T�շtD�H�"O�u{�ߤQ�h` �c���B"O�����Q�-t q(��E����"O�[�@H�w�Y�R�]�5����p"O� |�YFL�_�nl�2��z}���"O���1��u�>��PE܈XR��CC"O���O=Z&�"��C�ߢ�s"O\;#.I0iJ�X� Ne��x�"Oh����c(���Nщ)���"O����փ5���$u����W"O�,�W -H�u��"B ��I�"OV���g_�#~.<B�`��>m�"OlAK�o��)�kB�ѱ&䀍i�"O|�P� �/Ҵ�K2���2,�|�"OLIz@)+~��E�S>�Y�"ObAH7�Tr�v "���[��4a$"ODaj�L�s���p�N�A�;"O�%��
}�8�ˤ�A=5��[�"O|3wǙ�n���οK8.�c!"O�A�R�Wkin�z1m�1XLa�&"O� ��	 a74A�7�^�s����"Or�g̪0[lU�{�ZV"O���f��!��I	�IQg����g"O*}Pf#CUv�!���S"���"O�����)$�49�d��F�z��"O�8�7���2l����IT�H�"O��eś�:3F���J'�*��r"OF٢"-яr!4<Z��͟V�r�"O ���`�_�x�{�� �z�CW"OX@�T-��f�\�j�Δ�0��A"Oh�92h�6,�̉��(��~: "O�D��e��!`҅��h��V� �`"O�H2�˗�W�2��Se �0XF"O��:�@��3*X�դL!D/d�K3"O&�I&�V\�a^X&��"0"O��a���Z��CC�фp���*b"O
 kw)�g�. 
Pj�=A�Ȼ"Oֱ�e&� 8N�i�`"�<#�)""O�"�$�^�^�!�˕:!�nM)�"OT20Cӧ�N���A�R�!`"O�8z��K+!���:w��=s��ʤ"O@0���NQɅ�jf��"O�]�tVBu�!&��Aj"O����1L�8�e�<w���R�"O
Q�*<���
h��D��"O��9@�4[�������,���U"OH�S��U袌�VD<C�V�;s"O��!jV(Bw:��S�d����"O����'�;��#�L�h���r�"OMp��"b<��� i��x�X�@"O�	f��4`���蟢l���aT"O�}0Y=Mi�$Ʌ
D�p 0Pp�"O4�cZ$c8�4Q��G�g( �j�"O`��O��.��|[�Dܿa&�H��"O$X�h
=s�(Q)C��0}�]�"O���&��i�4ye�	 -�5"O>�1v�	{\����V�}�'"Ob|�&�|t�m��b�5��L
�"O��yC�YH�P���Y݀�CV"O A%��1]L,Zq�N)/ي��"O�Ԉ��S6C�����Q/x����"O� ����9L���1Q�
�:�r�c "O ��dؐU+.d��U<eG&�%"O��3%ͧ%����#��r+:8��"O�`�Se�!��ՙ ��M��\K�"Ov!Z�e^�S�N}��U���%Ң"O������hl�)�'��5� �%"O5�Wč3�͓Eh��*["O� Y��n�p�(4HȎ�L�h�"Ou ���"�A(Y� �R�"Ox��2�Y��!i��:��b"O�Q�   ��     �  �  V  �*  �2  �;  9B  �H  �N  %U  h[  �a  �g  /n  rt  �z  ��  :�  }�  ��  �  E�  ��  ��  =�  ��  ��  �  T�  	�  ��  ��  ��  �  Q�  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p �'��I���S�O��ٰ5&q���R��|{ �	�����`P���Č(V���6nN8�ў"~�@�9T�,Sn�:㍉4�̠��	�<Y%�ҰJ�$:�N-JƲ��rk�П ���]hdI��?-4Y�FZ^�Db��7vTQ�Q���R`���eb�BB�ɐ�X��4�@-QV�Ț�BZ���	V��h���!�Q�K�ν�@�D�l���"OL�`S�#^���`���~J���"Obl)�/�Y!��9�H^D!�"O�A[B�^�A����R31hV��5�Q�PY��Y���U�����XAJM<2��P��7D��rA��6/l�\	���9��UIDd�O|B��7G�0lT4E�����o��N�B�I�l�R����ϲ%�8�����S�B�I�#?p��tK�K�"�#���3s�|B�ɍ*j�$� H�o;I�@V,b�$�>���)H~�����v�94%ے�,�=�ӓ[K4�˗�\�)JlUچh�� ,0��	���))�N�? @���J�O�$<9���D���"O:0�B�@;r���o̚I�h��3�xb� �O�U���7m�f�^HS��__��h�E����!�I�%�H-�r䎮\m��%M��wz��$���W��axBY�BDy�&L)as�)j��p=�}�jK6I�ܻ�ֳa�|SՉ6�yҢ�x@d1aI�_E�-��"\��?���T?��>��k��{����F@&�p�����w�<A�%��"F{�ézS�=��]���EFx���"�(yjĢ��8*�IQ�R��y���@E��q"�и7�B����yR���.� R�Q&*��t0 ���y�K^%B��h����d����$7�S�O�lۖ��K����ڑ�����<�'M��P��Ŕ')8|M� �R	$�h��(������Β&+T��5o^�I���hO�>	#i̶�ͳ���44`t�$�}�<Q��M����Ic��V�)���o�<2������,���`�g�i��p�'t�u�az+�����	�!��'\� ���8{������q��'�t�[g�̤W�d���ӥZj0h��'uT��
�n�0�5U�`��k�'���i!��U�Pй����	F�=�	�'��Yh d�M��(�ђ���Y
�'�6��S(O��9�AV  �6��	�'B�0��+�2M���b��L呂��'t@XR�Ԛ+R)s�/r�����'��h���	x<� y"�$:(2ْ�']\4�W�����gi�E'����'��qY ���=~��b��:<�.qB�'_�T�C_ά�!Q�N3���9
�'ٌ���M~�p��@�'�@�	�'PxЈ����KE���0J�%�6�1	�'� 銔&�.7�}�A�	"y���'���K�@��Ѻ��	d�Q��'����Ï�f��r��6 �x�'r:��'��-&ҤCjN64"
)�'������u�z$P��Q<=p���'yT�5���Z�Q�)�!7�X�)�'�Zp06!��8��})ч�/1��8	�'��������Z�OCV͠�'����3`ш-I 1��i��ɑ�',��nT�=�dqQ$O�C��i�'����ĨL�gIX]�CdX�qnl+�'7n z�^�*���J��i�RY�	�'EF�ӷi>,��a�j�f}�4�' pXk��&1}�5Bb�Zc�8-��'*4�v�"r�E�a�>#����'�F�'�7	�ȴk�R�`ٻ�' (���ӯD�Pհ���}D��
�'���+c���-:<�ᇮ�uX҄�	�'?tՊc�+e���F�	E��i	�'X(�q�-U�,���kS�@
L���'5B@+����Ȅ�`gC�D��tc�'$xW�E8aծ��&m�P?<�	�'hމpf�	z��6�`P<�x�'H4�J�J�=X�"f�D��bD8�'����jK7r��5�Fn�uy�'en�s����%:=з�"=��I�'�婴�7�fM g�#,�'l�q��iߞ
O$̲f�+,P�aJ
�'`����M�)��Fg�;bt�(
�'Qt�׏Pe�$P�j��|J	��� 4L�vM� �p\��.Z�����"O�Lx�A5�D�x!�R5�0و�"OLAЧ�@�O�}G��h��9��"O���L��2�^�P�"N-��"O0���X�`��KGb�c	�1""OBU` &M8Pll��F�s�$�@"O�����v*8ॠǔ2��Ui$"O�]pr�G�#��ժ͊2nǬA�t"O���s/C�V��)�6f��k�(�0�"Ot��	L�S��HӃ־6��E�F"Oj(�w��B��!`�����u�"O��
5�	�c�R�1�A�%�HY{b"Ob��3�͟B��I�� hT!�'"Oj� �/Y`B|Y$K�eO��jQ"O,��ڞL@E�v��E3$�+W"O*�e͜
�cU�9���bQ"O�y��oߪaʲu1S�Y>e���٢"O�tƃ��S$E+�ӥ.����"O��#Dg��	| � �芌�V�c�"On��q	ϸ�� �ĳӤ,��"O�4)a��d9
���jl�"O�x��oE.t�>��h��K �5�"O�y�P�uԼ���d�(
�"O�5�� �'t�d��D�v��5��"O9�bw��h
G.RI���"O*5	�f6�M�U�ė���Y�"O��JB�Y5{���i�KP�%�L��"O�5�흇H&���jI�ydLD�"O��'L��`4�������"O�A��yb���h��p�E�f�!�$�=[��IK��D&cb����,6�!���=Ǆ��DnM0+Mn�8��\�S�!�D��B͎h��M�`4�Tѱ�Y�z!��M�\A�Lp��M�2Bh���$�"b�!�ĉ�.l�s	S3@,L�	Ȃ�!����(�&�LW$�����˪U�!�$[���dUC�O-�=*���{�!�ז  ��$8Uz4��!�Ҁ6><��6J\�H�dU!�dJ3Xä@���e�YH�b�/4�!�DL#mN��:Ў��[��YsE���!�D��t�AW�ȁ:�%�Q��j�!�D��Kg�a�k�ܒda��y!�d�.�Hq�o�:B4��Ď�!^!�$[���)S���;h>�X�C�M�!�$U:r>�lk׭�LE�%ˇ��'�!��Ϛ#�t���NL�t���ɢ��,%a!���f�������8Y� ��1Y!�]�e4P�-�,O���AiP=�!�$Ѩx�H��TN��Y�H5�X�!�OH|�0�3
�-K����NX5N�!��v�b�r0f� O��+��!���ZJ(4ص�:\��$y��I)e�!�Vj>��W(�>�~仆��18�!�Q"M�(��UaOGz<�����Tj!�d�2>�`���MB(���H�K�<q�*F�� ��@"M7bm�q��J�<�!�@*�|�P�bzF9�4ȃG�<A�G^�gVT1���: ���5��l�<�Ƃ_9�,�ң��,���pTk�M�<daE-$hJR�+۰r3��H��I�<�N9sw옩��ݗp���`��C�<!���Cζٛ�C}�F)8���}�<i�G�@��\��.�2o���0e{�<� x� ���Z�Q��^�/V��2"OA$��S����L�t�@(�"O�IB��I�N�Hك�^4�0sQ"O�(���X;C��-(�%"�����"O�Y��O�_���сS)~�����'R�'Z��'<r�'<�'j��'����Pc�^�K�b�!9$�Y���'���'b�'_��'���'_��'��cdF�?2^ԍ*̲Hh��'w��'	��'�B�'{"�'}��'g����Z�j_��X�`]3X r�p��' �'��'���'Q��'Vr�'\@�D�L�c�����'��'��'r�' ��'4b�'�lH�!�'6Ĉ�+"J���3�'r�'���'4b�'�R�'��'2Epa�f?�!m��:(B�J�m�Or�D�O����O8���O�D�OV�$�On5��3$ڑs&�,?��02R��O���O����O����O��$�O����O̴)�L;6�����^)'��ԡ"��Oz�d�O��Od��O`�d�O����Of���D׶.��8�.�)~���PA�OJ�d�O$���OJ��O����O���OV�1��C�b(B�_�k�p%3­�OF��O����OD���Ov���Od���OZ��@��=V��r��^�l]��/�Of�$�O��d�O����O$�D�Ox�d�Ozm��5=4ׅ�?�˙P��'gr�'���'�B�'S*7m�O��D�8~������
�	ó,�T�W-�<1�����ر�4O٤TXҫ׎-�$1Bf�-�yr�mBD~�$`�Z�泟`o�ERhh�l�6���s(߁|u
�Yٴ�?RŘXz�'k��4�T�C�~������,�H�"��Z�Ɖ�wg�_��?�/O0�}z��2.��k�D�NQ��冄����Å$��'n�h�mz�E����;D�< (d"ך�F��!HK��?Iܴ�y2S���l��a�@A���X�4�D�
��eS�� -4P��H!(�h���^�L��=�'�?a3뙩`M$5��*�T�2����<.OP�O�mZ�W0@c����=\X���#����H}��]��I�xlZ�<�O���3�8
@:0��� �������t�ʆ[0�S,(擓X6$9c/HПt�`�3:R�x��Mw�S�wy�Q���)��<Yq�����酏A���8c��<���i��5��OXAnZn��|�S勬&��%Pխ�*D�V��`�]?���M���Z�@\	F�S~b(�}Md	�'
YŬ1��T
`OؘC�ݷKQ�y!T�r"�˓I�֩ �*�3�D���T���  A�@��?M!�BY��͚�(�,��*�*Rza:��um\/>� �����UAW'��V��E�������jA(WnYJ	�N�|�x�fA:6��0�
77�̱+��Szl�#�,_� ��N�H�ȍQ�D,$H=���=#żQ�%V���V���Re��b1�P�7��]q3ǕU�1p��/u��'o��'��$a>?��kѥ&ќ��ş�Jr�W�>}���'���6M|�OK�'Q�ĩX�ԈD(��T�C� �mZ�S����4�?!���?)�'@#�'BN����@�.֙1 �L��ƺ�
7A�v���$����h���Z�4�AR�K�7����%;�M{���?9�Y,r����xB�'�B�OV�ˆ�	V^@Z�&ͱ�a�T����H a!�ly"�'���'��d[��t� O�V��}S���!훦�'�2���Y� h�����?牿JZ�}����vC�H2�"L��ɱ�Oؽ�$�M.h6��ş���ܟ���ܟ�rG'dQ��x�W�X8�Y䤎hr\9��ɟd�IП\��G�	ПX�I2��M;dó!���c�B����$�<9��?����?q���?�gG����N	��T�B:M�$\�ã4�M���?A�����?I�>��{qg�ͦ�p�9�6�h���	/��w��r}"�'��'���''����_>��I	6�Yp$'�"S�Ri�І��%�j�"۴�?�L>!��?��ٻr�$�&� 0 ̈�}�d���w��h��jjӮ���O��)�$$@Q����'���H�?�ha��*$N�01��0ՠO>�D�Ox�q��~r�㒜}�ܘQ�D$!�A(�F��Y��П@C���t����	�?��	ǟ�7m�bM[у��E������§\�7��Ox�d[�_.�c��iӠ�䈨��g��j�͞<Lٛ�i��2�'���'B�d�'��\>����WT��`M�=G�K&�>�M���=��Q�<E�4�'hPp#˳8pluYu@R��XK4�n�6���O�D�$h�B�D�O�ʧ�?��'@����/5��`1��y߀X�A�;�	��iN|"���?9�W�BD�N�G{���E5��)U�i�2��1$̰O�D�O��Okl.pt��?1<�=��)[�V盶�'�E��V���	��d�IPy��'*�ի0ŝ]DI� ��:�6!��n>c��@y����9O�˓.2�3�l�6��F�B-8����,6(��'�Z�M�����$��Y�ϧq.)��!�!,���A�$C���'�2�'��P�����P�q�~�G��w  AX��,�����C�O}"�ͥ^�(�0f@A+��h��mƠ#��B���M�V� ����B�.���qCÒ��y�	�0t_ҥ�D�(u��A�n��~R] %V.X��p���D�>&��U�d�7[�ء7��]t�9ã�L�t�\p�K��]��@y�o�2����7�1�<�yv��I�~�� �C�Hw��M��i��8dj��R�� ���e,H]̡X�̑����ɦ��S@u{4�����	��Pq�4C��	�p5 �Z�O �$�O��2�!�[2<  �ʆ�M��$ѣɺRh<�&��<B�-I9&=Bp���q�������	�����,��(M�`둍��q�͖!y�-��F�(��Ÿeq��l�-iQ��
#d�[妩�T,J)3ʘђ�'�D7-�tyJ~�������R�t��0�	��f̋`>!��j��Q�� R��L���X�6Z��0���Ӧq��-T�zyHv�?*��ё䜯k�L���Οh��Ԙm'���	�����⟜�Yw��>��q�M��g�\������B�J��S��Ħ%��0#�h�P�W�i
��I��л� � k΢����P]9زƉ�E�x�%*�r��h��?�C��=��6I�X�����8��	�������^�Ė¦�r�4��'��a>�)à=w@E�����X����ȓ�eX@- �a�l �2),$D�I3��I�MS����ȱ*�(Po��逐(��;B|�z��X�sxv-����T��ꟴ8`����8�I�|�����5z,�у�2YK��ړ�N Xt<8�g�Q(`�����3�.�񄒆X_�����:7������D)���7]�d���3k�6�A� �t����c�nFFi�foь�V�EdKȟ�?���9O޸"�B��8��`
�K�&�K "O�X���Ͳs�bUA�t���a�?O"�l�ß�'�^h"��f��d�O��'N�~L`#�X�/NR�@��Hwj\�C"*��?���?�CK ���9 +�IAE�O��o�zP@�ő$:�(�f%ʥ?l�<1�䚋\Ƥ�A���=N���#���u��V�)}h�अ�b�ڰ��&C�)���$ڢ	�e���d�O��'g�F"��̶�Z$��!�I����?���?���|���D,��`��S�(8S�O�P�a|2n'�R�:.�2r�t�B�kS�J�^��D�C�P)l�ȟ���`���Рs-��'��	�b���OL�UX��d�o�V9(u�2�dg�(7d��uβ~�O~B��	H�$o��V�M�7�	�d��� �Z;y��k4�=iR�"E��=o���I8�Ͽ���N�7Y�����f���0n@�{M������?�r�i���OfI��B�$H����7�	����3Ot�d<��4ړ�?�e�N-5R��℺8����q�BN�'3�7M�禡���M�+�b���͔���&�."�������7����O�A���3ja����OT���O8��;�?��O��Y�wj��̨�Q'�A��q�N��I��:P�3*�%�G���|��N�9�0��<�wj��\��@B���}��&�N��i��(E Q���Æ�Sˤ?�K�ㅉ�1Ot$%�2��a�& �4z$A���O����'Ê7Mp�	�`��ty��ȗL�0E懬:E
J�����-�Op�%c�~9�)+��æF� ���Hʦ��ڴ���|R�����
�<��lڬt���4JI����C�<m���	������x�"��4������ň�����N �#
��	_2�H�A"��I����`@=�"����N^�=�dɛ��`�Ks8�S@b�8A!��"��*8&p��aN$E�:���^�sD2Dd�:4�To��>$R��M�?֌m+T��E�	Ly��'y�O��$�O�´(�2o���ŋ��}j�k ��O���d�\ۀ�Y"�e�@���ܴ!���_ߦaSش������'�B_>	zr�Ʌ��4[��O�*�>�1뜁<��l�	���	�8�����)��:W��	�ԝ��͐�Z�p"�S'8F��&ӥ	F<a�#+ ���q-?
{F�]��a�΍n`���7�W�.����#�-�N�Qg��rTQ�#G��O"�nZ��M#����,6��Zs&��T�d���n�k`���<a)O?牅1��}+�&¹F9|����
;~����&l�ǟ�`�C@�d @��|���v���� �)�I۟�O� ��'S��'ʂ���lT�\�@�VD˸�ɴMB�`L ��D�µ�M�����˧���<	A��*|��߄2i��Y�H֥w~m�V�\066ٹ� ~�]����'�D�iRHɮj�D��#-5��ڣ�T�&�2�'S��?F��s��T#c�xH\!��	���?!����P�I�D,)W�R�+�B�#<�t�i\6�:���?���'-p\T��m�^S�(x�m؟��I04"|{գ���x�����ɐ�u��'S"�O�1OE3�GO�JI�h�;*2�x`��5j^�Й��4��)��O�`�<!6��St1���7 ��HS�F�~-xƃ��p>�uk�����')��T�bh6�	-h��'CBFy�u�V#
�$��ə|3$ �I��MC����,O.�D�<���� ��	hsB��5�9a�ˈb�<)�"�L*%їiH.a�D���F
-ב�4�S���'�\���*e�*�
�#�.L�e��1k�I��?���?!�o�B��'�?��O�t��5=F����H
{�|���`��]�����M�|����'U`<�ϲz�<��Vl"<F��M�'bp`�&��$]�����'q`(��?iE�Q=t���p���^�\���ɞ�?a�����O���{����c�J��"Gn�>>��(�ȓW�����<>7>���&�4mH�j���'���Y�	�O���|� ���ր�,|H& ��/�{�~���#Y  ���O��䅯H�h��4�L7E,<���SΟ�'9�j$z����z�f�����yתyGyR�T�	�*h��΍z�������X�Dy�'_��< w��N,ty��hI^]*}Eyҗ�?QP�ir\6M�O`˧[��4b����yd�j5+I6e.�y�������U�R$���!�'{��!Z%�Mo�a|��.�^A���vc�@�H�SwCU>#|�$@|��mZȟ��	^���;`(��'=�BG�A���
�IJ�1�O<?���\,��}���@�>L��ʋ5�q����w,��9&O�%N��r�mI8���¢��J <c�R�w���`Q%,NX8W����Ͽ3��H�T���� ���-��S��^<C��$���v�}����1��\jv+]�W��j�a>)u x P�}���	`x��jCȜ:k��� ��? (E1:}��@�럼�R�/��x�dկl��A�cg�zh<iDK�����Sg+L��2��X�<�*J�+
��2���y��� ��_�<ע�!t�vd����v�^�R��r�<��/ fP�Pf���E&�	m�<I��0
r(
F,�7'(艣J*D������%x؉e�*�ƥ��A#D�$�W�ͫ�1cg�ɑA��ȉ �-D�BV��3�ļ���Ɛ�
!��*D��� h�LA����-@[)��� >D��I�:��H&a�;����"=D�`�$؟y����T�5&�p	s��&D��1�+){��P2��
"��|�Ҡ)D����H�O�����Mz)��%D���u)N�Z��ņ�+b� $�&D�87��	
(8�C�g�6|�A�K&D��ӠF�I�5�EDB��Z01T�%D�l�B���=�0a�-�G%�D��"D��\�'��3JK�[��Qda?D��{���1f�@*!��0��h�U =D�T��n��yD�Ix��[9r	z�u$=D��[ak�6I�"a��b�'\稉9��;D���щD��FK�3a
��@�=D�4Zt�2ddJ���IV)Lӌ	r�=D���AM$>�dA3�XJd� <D�08�f�{���hBGQ*�, 	f�9D����@��zR-�LjC�	"MU��� w���09�~B�	�G5�\�P/ ܠA�hH-B䉇ni���sB�s	�Q���lt�B䉮۰�w�̹g>�򇎓h�C�� 
t�UȚ�S�(�s�e= ��C�^SN\��ǟ
�*�p�����1����ħ/�~R��8 aW�\Jj@�楂L��p�D9D�����	�+X�yۆ,8�c'�b��0Cp/[�$��
W�4l�����
g݉����`�ȱ��A�Da{$	v� j� ��U�Αʒ�X�wj���ܺ1�)�T��l���D	8"�ph�<��i8�삭`!�O�<�d#H(�$��OЁ���>	��X�L��lXTC��^�бQ� D��He�	��|��Gy�`	�cΫF�*�(�',~ur��'��#}�'�����o�� �@�+�z	8�':E�B�&Xgz��c� b�@ش(cT)� �\/S���	Q��p<���Dkl1�t-�]|}�G.~؞�P����oz�Ã8MV�|��A�B�P��qI�z��g-�w(<�t(ښ7�x;W�1�Xt�/Lq�V]��	Wd(�F�J��L=��O���)��$�na3A(τW����'BR���)�\J ��+F��!,�82m�ŭDៀX�j�;��'n�O|[��˅U��1�G�h�t�R�'ʀ1��l��`v�:ѠF�Y��A��TPHbπ�S�ju(�M�P�(��E�'oF-���Z.] \
��J�7 �hy��dA�NVr���B d�ڼ�Lۣw#�F�LXdi#��� �f�@�菞{D�8��.xTUZ��3�Zl(D�ݐv�~��'���jS*l��)�7|**,p째O00�*�LT8K��xr��W�f��@��0�(� ��І�0V�-�W�H~9(��$�!��O��	� w:�K�ݮ&H�u.ׄQ�l�2��p�'lv4�DJ �39&�ak��~~�$��4z�|\!3#�6w�v�i��QT����k�fe����.M�<��J�J?����CX�H����!K𴂖Ög}�L¾(�4[���\6<�[vb��HOH�9�����dN�Aj�PF��	���wQ�h�:A�<�Sdl�{�Q�l�Q�G�)��A#(��Z���	�6[�z��V�?��O"�M<��.��Cr�%��f� F D,uO�n]8"%|O�)�ݥ��go^�*�ҍ����:�41G�O^�n�dh`��� @�V���kK�o�"���k]t��ii����|��D�k�PF[���v'�Eg>�K�,ɦ6�,bE�Μ��$T�?�a;B6f|�ȗ�s��$r�lC([�� Z���<R��tys��+�T�A�G���ɻ�Y��j,J����	 ƺ#=��i�8��p�7��,_����ެ����7��=3~��S��)�j���a7�=
���boWK���m��Q�J�ӧ(hvvd�0�'�B�R�j
<�9'ϑ���:�bʐ'������ˮ2�{"��JJ��PB��<�p{eD/-~P��P���@ǃ+'�<h��Q�Ab]X�ꑁ\�O�n��q(����O��P�`�|Xrk��!��i�����n�W��胇Η�Z�D��.O�m��*6�eG�ʂ&�����hz��a�Fd�DƑ=X�=B�o�0�1�4����	��&�p�Χ6�����!�;*ѣDï|���R�D;q�����
�0�ŏ�OEȵ�${�*�>� m�?	��M1#/\�<L�4�5!�OR���Ԁ�4sraz�7	�~ d`"��Q�Uh��T�Dj��!�6!1G�'k*fdC�� ѫd��$˨�h�ݩA�?F���j',���6'����� ��p'iD�k�@d�"��7*�%q����	��\�*�5A��S�'��
�fdߏs��y�E�ʂ9:,��w�$v��b����'��Ȑ�)�j��� KΙz���=)�Ȅ�5Bϋ�r����a��ɍQ�^͊��\g��S��B"=�ԋR��"�c3+��:� 4�'��ۦQ�I�4�f$zW/	�&s�p��E�';x�Wk�Z�,�"���\�^�R��Ǳ>5V`�Qh=�j��O2$�5��7_���+>*�HK�!S�Ӻy�	��y'BN=qM �� ��"@	�"��'�(�Y��2OT��WG�P�"1!@�*n:�3-��3<*���W%`!�D �Ϲ=�i���qth�	��>R/��y��6�`YC�Ƽ0����$:��qK��P"���pГ��K�h����00%��y��r��Lp�m��r�tAc�b�:��E�@�$�Pxr ݾ ���!LZ���;�lN����E.!R�ݚ���&�-:�fO ��ɐ�OU�Pː"��j�xd[aJ��!�D�M�֑�� �Er1 �Jp/�|Ӡb9�����-�Q��T,c≯6dP���C���e��� r�rB�ɘ!� aJ�`�[$���n$&P�B�;.�4U۴㑶�����$	p\B�	�=�P�� :.z��G��1�C䉣$����3X�B,b�D���C�	;>�(�Q��S�6⢍.O��C��%����E��*66$'o6QrxC�I.ؐ|sː!uVF�2�"�9�<C䉔&N�!9�#ޗ�f�ʁ#M1x3(C䉢=��3��JI��B�I:��B��"At	f�%r'(��h�GK�B�	�q��={�HM6=��w��hfB�	�r����"�)g�ĤR B�0Ss�x�T�ԤU�VX���ǳ '�C�	���(�QLڥQ+"�y��>P.�C�I�5�Т,�w�`s`NXCܖC䉮ǚTA��9��-*�l��P>�C�	��A:���.�n-0���b/�C�I�*[���&h[5�v�CŢ/	pC�ɷ^r��cB�n�2�b�)eƠC�I	N����$���q�bرy1LC�	2�����J%x�V��@w�zC�=DEvQb)˞9G<��ǡ�`!�B�I/���Ԏ@t�.��D���G|xB�;X^H�z�IF;B=,I�c���LB� o
0����FY.� ��B�4B�	�L�(H��HA�TI q�D�߄i&VB��*N0�㤉]lΐр �c�nC�)� �D�q� �"��1�/�5LV<ض"OD�uMјY�Q�F,��^A��X�"O�� BDۖn���r�j�-����"O� 5�H�J��i������N}�5"O�3��X>����t~Tۧ"Of��r�G4B�+�IL�ܠ�.�{�<�,��|�}��κ8v�=�B�t�<�i�[������m^!�+Ve�<!3�G~��Qx�-ʶr��W�w�<q���xx5[v.xh��p�<��U�6�,��A��:!�ug�i�<I�\\��S#˼V�*�[d�b�<a0cֻ"����W�E<6��)�'*_Z�<9D�:|e�U�!(��;�&�<���S�:��GaX�0Z½�D,�C�<ёK�5^��6/Y�S�d��`E�~�<�nU ��RT�زx��	!�A�v�<	u�֒I²5y���������N�t�<I��Xsw�ܳF�W�
A q�'�r�<�����h��H���Q~�m�c�Km�<i�2(3�)Acc��N�#�k�<)Պ�]���N� 5��@�o�<����;�(-:��P�E�(�f`�g�<ɵ$�r�Bzi�7P�؜�(\�<���ک+��9�"��nz�]�Z�<��B��N�V�@�Z*j��5'�M�<��FL�1�h�Z$�,)D�����G�<yCx��l���ٓ	ک�(�X�<��oάIS���D��G	dApq�|�<���W�zT�e
M�'��b�<A�[���a���hɈW��h�<I#���P�H�(P�R��*���.i�<���pe�y� �?#-����O�<q��n1.�i �[<F�DqdL�<��BAq��J;^8e��,�s�<Y��4@���n�+xC�q�tKn�<y��PT�L7�٪NL���t�N�<�ցJ)(��Kn�H�|m#VJ�u�<!%bX�H�
�
VK$�Qb�{�<�թ�c`���%׾t����%��u�<��ʃ{H�)S��ۓ
0$5ꣀt�<�&�6ZDA$ȧ)��5PB
�s�<���$1XP�y��8�`D/�Z�<y'G�">��qq�O����sw�P�<�1�߉Sd���t"Q-H��t� ��a�<�S���q�6�;F!&�:�ڧ$�`�<�f��'>-B5�*_�24cFD�<a�hا>,���%�SZ���peY�<��&�E��m�B����}p'�U`�<Մ�%�����N
]j�����[�<!AO�,Q*�Pg,O�6����p�XT�<A�.A'���K�FQ�"��H��%�D�<Yw��<�ʥ�s��:�D-2��E�<�SnLr�:��/]2�JW�[�<���&u��I,.�r�:#L�Z�<�3�M4"���= x*��3���<y���7f��[�,�3?dt�U��z�<	fAT��Ȉ�*).��1��t�<94��
n
�t�����H�V��ȓ;�FD�r�'42�؅L�OA���<:���!~\���+����~A.�[/�*O�᱀݆+��	�ȓ)��!���:r�iu��8\�2ͅ�dE�r�X1T���"��{u�t��S�? j�	u/�"xg�x�4�ǧ��4��"O �xP!�4o��z䏋Jˌ���"O���R&�bM���h�A� *�"O68�2���P~�wǘD���97"Ox�K����h���Ae_ �@,�P"O�H��A�bլ���CR.����F"Oʐ"�_�Q�q+W��?@�ZP�"O�X����YJ:p��Ŧ}�X�'"O83��V�6�r����5e��=��"O�H[发�f�nH!�˸U�8�[ "O�mRB�i%���hȺy�eC�"O.�CI�=�J�i��7w��q�"O��0☬[��Q皞 :L!2Q"O�u@��-��q��U$p|�"O�\�`�D.�����
��,��"O)��-�A|�s�[9O�|M�a"O��3P�]0fNxc!T�r��"O.m�� (N�ҩ���Ɓ�L"�"OT���l���Pe�����F"O����E:b@��Ӄ�� ��m �"OL�i���Q�f$��Ì�`�t%�A"O~ �6L9�,��m�=}|x$�"O�}b�JӎQ�F�3�L��_����"OŠ�Mȗ���Z�Dљe�x��"O��#�i�5X��E� !Ǝ8 H"O���D��jS<P�# �)A7t-aw"O�]��8x| ��݆]3f Zp"O|���F���L0R�v ��S"O�q jCK���F���r�m��yr�S�#�/Zg]�HW7r�6I��j�V �%	�.I�dmh��1qL�a�ȓk��tk< �j�p�	)R���Q̐ b'B�8:,XȲ�ߤ%&�U��N� `5D�'�tPáF:Qx���k� P�$��b��ƕ
3x���p	��YUA2|����$# #8V��ȓ#r.I;�iV�}#,s��F�/��`�ȓA;Td��iϛw��V��;VK0]�ȓ#T��s��6-P��`hQa�0���(4ZDbr��0��L*��G�~�rԆȓdڝZ7lν'�6���(a�ȓP�q@�(/�&<2E��A�>���SoR8hʣ�x�"�-O���ȓ1f|��	�3
�����'f� ��ȓCv�|AN�wV�H�-�! DP�ȓA��!H�*N���&�X���P^��s��Xr����"��)�r���D/�<Xwn� dq"	C")S3��E�ȓf-RT�
��W�Ji��ʵ)RR���1e��(��͋l`x����,��'U��Yg��|��j<�80L�"r�bmpe�$�O���k���5eS�Eȑ

	P@�t"%D��!'�ş τUc���
z8�9d�.D��(� ׇi�f4Y�b�$9pm2��.D����&�5sVq�F� &���1��-D� �b!�Bh����Z1��k�',D�,I ��(~��+��@X����(*D�����_�G��p�e�Z{�l3�"D�@`f
$ڨ(���]!	���#D�4k�'�$�Thz��ݽ)P�j�l$D��+��W�t�a@�^�6�d�<D�p��,�
7��{a�n����sC D��aa�Y���P*=B���s�>D�@ڵ��H&�$�(׮J]�Q ��<D�� ��В��0˨�{�ߚDX!��'��O~�p�!]�!��pr���
�"O�1���	{����x%	�"O~l�5��6i}���3�ϯ	��\{�"O��0N��sAL��`d6;v0Y�6"Ox�q��k��Y;�BCS[&��"O2$����� ��A��@���"OV���^!Lk�� �	�v�p�""O�����Ɣe�L�����	"OH�ɦ⒍5�5B&�
W@�q� "O6��u�Ԥfsf�H4'�*p�&"O�\jg�ѹ ��I��Ń�j��t�"O�#u�>~�����&�#>oH��"O����CK*�åŅ%hZ�;�D(|O����ڗz�P���ӝ ZT����'I������B�XT��1)ЄF{���'C�QYŉ�'�Q��L�(=Hh������O�#~z7�� G�D�z�fש[��rAUA�<�f�Ѣ�1Q���� �԰h�B�y�<�A&�%��P���=/S<�Q���O�<9uB_.ڎ���nO�2���!�O���=���J��� ��Z�؉fPT�<qã�)~L�Se�e���M�<)ǚ"ZG$@
JA�
�гF�J�<�2�D0���[1%��H����Z�<i��@��,W�ɖc�.��@�]8�(&�܃����>aj4�Pa��7ﺸ4�+D��xdݧn��c7/�:��{�*D��ـn�2o\�c���B8���#D����ީ#ҩ�.�@R|���3D��S��ڣP��d;dbD�"}"�z'B1D�6e�@�`PgE�3���@-%D���0�F�
QP�6$34�u�eM"D�,HbED\�j 	�k�7f���(��5D�Ȑ�<j��h��E� .l^�Xc�0D�hY'�X���9Q硇w��k��3D���cY<�*��wn�s@��L2D�dZw#HEm���'�l��CR�1D����G|5E`A#�2�ȡ��l;D��˒�% 8��
rbS�3>��jT�9D���b�
����j�o(F��ҏ3D�P`�cT�N��{���W�n�3
'D���WBV�0[f�0K�+3�BXF�$D�D��B��"@�Z��F���B��+4��X�聅n?6���K܏oTC�I�A&i$OM� �ʗ���[]�C�I�c�<(��G�l����m�.B�I�t�T8еo�*)K:�	�M��A��C䉙h�x��$��_r`�en *�C�	�.}t!$�F�/E�rlN
k'�C�I4|��@k �ȯ@��l����$H�C�I��}@$,�$��ݐR�G�`�TC�	6�c����l���%�#|OC�	
`���3tO��V���Ǐ25��B�I8���'(��H�,}@դZ+ ��C�	�-�&(�t,_����-�2o,XB�ɧTϢ1	�4���ÐN��B4�B�I�t���� 	o��LK�.ZDyՃ1D�:�FέV-��8pk��|��.D�;�-Y;��Rw�`��}�+D�l���k�@̐`�C�kX����j*D��Y����@8D�׽l�f,H�#<D��8��e:�DsVJ�o^�zd/D���2E��
��:a"�={���("D�� D��1h�	��9�q��GP�e"O�D�g�_i�\�p	Ǒ(�p�"O8T1#J��O����0(ͫ %�-��"O���4�Q�AC�L;���>]�E"OXIKF�B�'��@�ʚ#��x�g"Ob�K���G�	�$@�j���`�"OR��	1
٤9��ݲ��$��"O���*�y����g�4����%"O�9�1K��Q�Z�H4h04����%"O�}��횜)Ѡu[��G*�ZI*�"O��@�:?L<d�,��}.(T�"OZ}� =2�1R��ƨE=؈{b"O!*�.P4ra
�ʜ�d���"O~隒h� �j%c
�	'gZ�*t"O&�#�a��I(`茙 �ԑ9�"O$L
��M�9���ЦV&��@6"O���tl�p�V ���#L�"OH	+"�
�]`@��r�X�'�M�<у��A�x�A�`�;�r3&DI�<�p, ��L{$'�RFڜ�g�G�<����ު���+3V!�u
7!�n=9�� *�}�q��F!�ѻ)��B���-r �T����F�!�DJ�l2���闃s �	�O�h�!�E�:
���̟�?�R�-��Jd!��C3�)��!SPJ�AT,1�!��|t�����M�.��t*�J�!�d�3`�B�A��ҙq��0� �F!�^�o��E�D�g�(�#�)�!������V�ǁb�Fhw	E;H�!�d̓j���xG�$�t!��GʿQ6!�D�P\r)�T����]�	�>{!��J* p�犭-��L���,�!�D C� dP�[8H������#;}!��ՉVQ��@��	{����v�!wc!��%�]�X�-+�F�V�D���"Ox�Q��U�nؘ`+:�j��U"O���#�����A
@-ڟ5ӌ}�W"OV��w��
CT@�R,Sj/���S"O�y��oԡc���b��S�(|[�"OP����4�B���ɒ�G"r��"Oh	��J'#��S1�~*��z�"O�8��l�#O^�����8i@� sE"O�)�#l�6� 1�"�-R$�!"O�`���Y%p� ��_,"�	�"O� qp��C{&|� ��[p ��"O�t���\��@�9p�U�q$6(�r"O,Hѡl݁�����OS$��K�"O*�T ͅoT�yf%3 �j��"O��+��6.�T�Iţ���%��#�y��¢(Ψ��(O@L��Z��y��Й{�Bc ����-L�y��>b���F�Gl�A���y�/�2Z��
3
/G�y`���y��P�!�h��E`��7��)J�$�yR��y��бV(5d���J�k	�yb-�7'V4�H��_YY��-�y�O�;K��y0�.��X Z�`q�'�yg�=&����ר�MS�Ш#�?�y#�>b�����D�t�
�j���+�y��#aC���S��sP`�z�
�%�y�^,,�pI(�� r,������yB�5} Pq�[�2�Qr c	�y�d��:����-�xa`q���y
� �(�UL�'#�y fj�>1b<0�"O �̎����KUj�[/��"OXE	�㈿&,
U⢈C��5Q`"O ��F��;7�=!E*�;�eZ�"O�Ys� ��|�Q2�E���R�"O�5�gN@H�ȚUhɵ)����"O�yp���Y���5�_+j��r0"O>-���.��4���,h�`"O��¤�����#ǘ|�t�	�"O�(�!*����Q�>��i�"O�])CL�(S� |��O=4���"Op��ҡ˥q$���#OId�Q�"ODs��_�&�TMi�e�:D+��*f"O,l㵎L�1�^]��]�4"�B"O����[l$�)#n�wL]�"O�P�ф���K��\k+6��"O�Qq'(G""ota����'<�=#s"OF��\8^J��Y4mY$-���s"O"�"tE\�}��|I�%�t�3�"O�m�bh�3��L�cɞ.��Z"O| ʡ�K�u���㋊.;`pA"O@D�7kްqSN���͋�P���� "O�e��׼_��z�L�gĠ��"O� :���39XL(;Ra�`�>98'"O�����W�!)q�κy�P5��"O�HJ�냪_�
��)I��� ��"O9�0��p���Q�j�@�数"O�@�ҩŔ"����U�D5@�R�*$"O���A+0F08���0|�*	�"OT�P@&�.8|hՙ  �>���"O����΢Q5 Q�Qn�jR	"O;jY0s��u,�Ri,�d"O����ń]����V+A�:xZU0"O����fX����	�4T	����"O6�H�H��U�z� �'�6a\��:d"OR^c��A�= <I��D��K|!�$_�j�4��U�^�$�x����m!򄖋X|�Æ�u߸|�&�CN!�$�0eÂX�e�j�qFU�!�d>J.и�J>g\��
�$@*n�!�$94Ɓ�
�JW�`0�  �!�� ����LO�iVrxQ��W1
�!�dA".� (��#m7J�{���y!�d�C%��ܬ}���k3�FC�I�}�EhT-̓E
쬘��ӦVB䉵#��Z��%�pΐ�NhHB�<��`C��m�����\��B��T��Qg��`�yG=�&C�	<7�w��4O�0Ac7��A�C�I�E�H@�����%l/}�B�I�:[4��U5�΄B#�YXA�B�J�:H A�ƭ)���C��V�B�	�W3j�ç]�c���X�'�3�\C�/[	Fh�A��,mg��#u�R�*PC��<?*�9�ÀS  ��[�;XB䉕i�^݉�CK	/B�2�D���B�Ʉ+z�<h7�;��������"�8B�bi�7ƍ7��P���A>j]B�ɖ+"^� &��u<�4�&�>f�B�O�@� ���Bh˙КB�	C�Lm"P��c���$�-JC䉊��2��!�zA��	��&B��2H谕�i�%F	{ �b8B��	"b��"w$�����>C�)� X4����Qyzt)��X3<Uv��S"O�L���T�)��	u�� jK^ͩ0"O2�K��"}E��c��:}J�"O��pH��3�XYp0aI�
հR "O� �(<_�H���!Z0��"O��j�Z�0ܱ���εr|tKD"O�� ���6m���U���8 ��"O��i5N��q�"%�RkM�w��\�"O޹;�* $�r	 �0�y�"OZ2$Q�lm��;�6���`�"OD	�vLh��0k�H�]���"O�� �j������>EL�Q "O��H&�l� � 6�E�'��[e"O�����1{y�Ұ��tz���"O��:,6Z�����U!)ھA��'�xR�[�{�P��윍a�,�`	�'%p��FB%w3��C�G��[�:D�'L$L�eAа{�}���*f�h0�'P�Kbl�-;\��cTgR*d��'ò�A��m����x�h��'Lj9�K�1P�r�5l[v�*q�'F��+����
CU�q8LB�'���!oǞ%MfyB���6bd�	��'�H��<Cr�,�C/��US��I�'g�!R!�ɾ/�PDb
� R&��'X��3爙c��2��a� �'I�R��^JҡH!B��'�t�I�'�|�@��e6b�0�υ]�8�'����WV�y ���*$ 	�'��h��`�4��%H�J�ܕ��'�4\��O^1hH���u��9��'��zņO��Ԑ�g�X(��'����$Z�L��M��&�W�p���'E ��K�'#"��5!ɮP�'6.�Q�3e�0��P#�>Q�'�� !�	�+|��n��V���'��A1���E�ֵ��@K8d�~��'�6l�7D�2~f�:ց��XV���'��8�c��SZ�T�G�>N�p�	�'�����ʠZ�ʑh�&�V�p	�'6,-���֞M�)�棚PAD�b�'��H�瘛0tF	2��NR��Q�'��͸P#U5 T<���ƕ�9�����'8.	��5m�08����$�E2D�4y  �% �01�!L�'�ƹS �4D��[�L��@�pt �K'{"�-Y��=D����G=�	b��)o.�A*�9D��I��
��x!<P�;�h7D�xc�䟁5���!��$[LI��`7D�`zC�C�D��"�� @1B g6D�̪�	�:V@���t�ȯm��4��
5D���1#6e�x;r� v��DCH3D�H�����U,�p�iJ�P����0D�� �#~`hҮ�20�V���/D����눬/��oʉ^x���d�<�A�/7��Uq��� �)�!�l�<Q,��}�棃Bf���I�q�<�V�UN����ㅏ�b;ظ��Sq�<qDߋ%H�����	�d+ *�l�<�Y�XN�꓍ j�,p:g`�P�<�	ܒ9���i��ؖ�� Za�BJ�<mK�2� 	:&���C[͡W��C�<��^�W����TO`��}�"N��<�Tl�	ҬY��3�"A1�)Kz�<� -�#J�!�*���U�ࠈ�"OV *ƨ�
2
1ڐ��Ib�:�"Ol����ɕ��@ZNX�h[yq"O�r�])P���`�;S5a"O��0�d��ͪA�G[� �+�"O�B��U�Gp�CDǍ'�P�"O�`W\>!� ��h�T9�S"O�(��J߄f�2YVfM5vLaz4"O�a� �(�N���F��K>�l,d!�N�w��2K�$Y�@��!�#�!�D�kP�6f�qMt �G@W~�!��ͪ�R`5��@�����E�!�?$ј��@�]%K7�� 4�ӟs�!��  �2��Q�B,
]�0��1�!�d� �����n��@���:}�!�䟑P%B
/P�<�b����!�D�x��	���
��B�è�!�d pD0٦a����ڰ���{�!�D�>�\Pô(��J�xj�C�F�!�D��v-�4@�er*Ec�dR�~�!�ƞ-����- &m�T:3�H0z!�$�,wZ��%���@zp(�<kR!�$�Y�Ȱ��cU�i���҆ �!��1ኔ��� ,de0�k<[_!�$P*m4��q"#���"!��3"N!��G�_(Zbc(�
Kh��J�eL��!���_�
!jdoM�O�Y��Ň��!��Ѥb��w��0d�X10C�f�!�ѳ\�"e@�h�Ob ����-s!��I"[�]���C�:H,�8��R�dO!�I��̲� R@��Uá�L�/!�DԌv��8�a�=&�NɣE3:!�D�Q�d����7TuJr`�^��!�%҂���i�~j��*�,�.;!�� �~(�ڰ8V�����!����ui�Y2BՐ| 1�`땃/!��CPn,`�o^,�ԅ�FiO3!�S2ae�`�˯0�Z�k��!��X6_���id 7(����gօ$�!򄑥S#� �D�ý8ҽJ�e@$Y�!�d@�@a��QB��)����T�!�\<=8@����'T@��"�HZ�!���+&l�+��ɁvBʬs$ N0=!�L���h��wW����NٛB�!�dI��l���HO6L����QG��!�w�\A#E�4�V�j�C� �!��E{R��*�(��	$�!��'Q����d��Dxb�A/r�!�*��+'¥f�LbD!��!�U>n�H5a�N�c�l%�+�W%!�d�.Oix�H�"��,�J0A���&"!��#�
\y��9���"Ú	!�܈{
j�O *�tM�B�T)|�!�$зY��q�]o� =�n@L�!���tR`!�ʵ_sɸ�M��}x!��
�}�4l��o��R$�I�[!�\5����m�=hh�A@,Ӭ{y!�	-�*����X~��l�3�!��#C��������<����A�X�!��,��U�%!̶�a�ښ�!��>I)���c&�~� �Z�i@��!�;y>&��ܑ���GR�e�!�D��l{��1��A�\�(A�����	2!�\�xPN@ rŅ(�RD�$�Ɂ3�!�� |ț�N%�ୈW�^�s J�w"OL-�Ԇ���e�� ���2"O$5�R�G=�M��1\��3""O�� �ś�j^�J�a�}����t"O�a3)M:wYN| �L�hU�qR�"O\�R�e�lS��x�ZX3V"O:Y��mJ�H�\����4�
�X�"O��iDdOU�D.��i���x�"O���$�J:B�H|c�K/2xN9�"OL���Y�敚"-�na��;�"O����?R���DgU:�̄ȓz���g�2i6M�w��(3<4�ȓr�6I��E%[������Z�*P��ȓHX�ѲH�t�¸+C���Nd4��ȓ	�h����!n/���#��9�ȓn���򂂂|jl�"�!
�+���n�n�S�E}����|ҺA�ȓ��=b��d��T	vgÙu1��ȓ`g�� q��F4>���G^�T����/]c"$ޠ�&��(�2�l��Cʹ��큧&�fܻ��Ϙ5�u�ȓ;��6oH'�Թ;'�29�M�ȓ"��d��C��i
H��cK>Wr!��j��8J�h��iR$�
TL ��@�ȓ/��}�N��--Թ�D�A�Q��ȓ_~����y�m01�82i^܆�N��c�F�jbI��B6�e��A�X��#�����wLX'k� ��Bb����gG(Z���aj�;P��3�Vɰ�lQ�)�5d��`�D%��8M�)���B&?�li��d9r�Ԅȓuʔ���J�p�2��77�̽�ȓ;�l98d/��Y�����ռ�ņ�JvH#��\�ou~���d��D���F�!eB�0x�T��0lY�A�ȓ �Jp��/vĨ);�#I<g����~�	���3Pl�Dw����1I�'<f��Į��g��X�����I��'5~����P�*se���J�B)V���'��ձw��X���$��>4%dz�'$��eIGN2ZA�N��4X��
�'h��S�͒>.���:ˮ�	�'Q�h�w��k4��X�/H�a
�'��R2� �τX�"��WU(��'HX�*S�3w�T�x�I�Z��ȃ�'u䨂��G1K���&A�L��'�q@�n�:�ʸ(q�R� D��'��͐t�~�(-��FCI���'ܼ�s���\��"�Bj$e �'��݀����@�~X�AO�
dNxy`�'��x�r��K�"	 H<Vs �
�'�>L�(;}ȼZ��	�Q1�Hr�'�\�r3$�6.q2V��CӜQ��'*~���Ӵ	f
 ��N��QT�H
�'84���C�x,��8���H�0�	�'�N��t Y�ʍ�Ыr2 (��'���J���w��8��h�m�\ �'��БFG$_�Ÿ&a	 gv&�C�'M���TD��9� a����b�z���'"۱ʇ�A�@!2��'Q��I�'|�-�u#��D,����Q�\�q�'�4��N�.!�.Y�	��r���'�@8�fO�wʼ�CS�ȋBuB�'r�P��Wq�1r�+��0���� |�s���H����N�a(��"OT��$�X�Ι��MP�h蠈c�"OT����6��,[5�Z�G"O�ti���r42��2�AX�S�"O(qIz�Lq�äV�v*⸣4"O�$A���W�t� 5�ɛr,�Ta�"Of����9��tɡ�_�%���"O2%�5�Λ	�&����2Ko�9�"Ob�r"��i�J��NY�j�Q��"O�9��� �-���ý`��5S"Ot���臖|\$��1 )/�*h��"Oޥ�2�ڠk�����~��"OJ�AwI"+���YtH[�L���!�"O\A���P�dl�T�6�ևq�\���"O��+U�4ǂq��ȵJ�2ds�"OhqGdS!H|E(Fg�9�pb�"OJ�Zv�H �ĸɰ`�J0�t!�"O~�4%$[�@$Y���,�$"O�8P�Evt 
�f�^��l�1"OPZ��̥$oБ� %�
V��D#T"Ò���Úx@�PrĒ,����"O*	�`���1�j��)߂�vh�"O��"m�\���I��+�D�""OH��)\���	��90�uBT"OH�9��
s�4��Ʊr�6�t"OB!u懣w�F�7��4�~���"O���k��~������C�}����"On�3��X�
4� ���	m��j3"OT��	�T+��COO.����"O4DI��m�*�x�f��&( S@"O�Y��I�8rc�Ir�&�Fx"O�t:G��8nXm�*��r�(a�5"O�킠#��8Z�����L��"O̀q�[wV�8��
'K��'�-RD�)%���ѡ�6QK����'���iէ3F�,�%�Y�U"i��'�(-��� tw:�\�SV;�'ZIEJ�? �p�[e�N7��A��'�t	��a@�4�;eI�-��Y�'�(x�T�ɝ,�.�HD�նE��'.P�xb�ì^�b�C�%�~��EH�'�ԙ1�j�>Q���(�����Р	�';b��cN
g�F�Q��×1��B�'lDLs��.Q�@��˒�(�P���'�tT���E�j[����F�7�'_XLC�],�ѐ���Xx3	�'����(�88p��L����	�'�*x����	rV��PF�d����'�u`R%�J�����_2H%1�'� ����7R*l�w��.b����'�����|ZZ��G*S�y�R��'��q`��D=�-Jg��q���'��8��W+O�ʖ-Pz?����'ڤZ��SX���!Fb1m����'�F����R	-�����X2k��U��'�T��P#L�b,�H^d~�!�'��P#�+���S��BT���'�.��L͌w�2�Ì
�\�)�'4�h�m�ND\ɲ�d�*{�b5�
�'�\Q�"��SX)�+T7��e��'�#2��~�:��E�!�  �'^>P�(&uða��j��28��'���Z����	8�ZE�͡���'�Dx�G�7�rk�!Q�X�8��� �	*q�8s5nt�3K�3h>�d"O�93G"�( 30DL�"�"O�YYd����ʉ�A��O;��ȓ"O���k_�1�@�0$��+ȕ2�"O ��LD%eP�yk�P7x!da�"O�t��]��(m��Å�w�@P�"O��ic��b>d��A#S�|��u"O�m+"˟�鴍�G��*�y`0"O8�QCC]<�d��b �8 X:A�@"O༹�Z�a$��H�oH�H
H3"Ovp8�.�6��s@]�\��"Ole�R�t��������
�I""O�xd�ۆd�&�!�M�*�Ц"O�%�d30�����@N�6m��"Ot�1Oْ3+���
HM�$�@"O`Q�#(�9Q�A)��S"ON�I��A�m��a��/	����"OFpz��	]\�  W�r��%"O���р�2:t�A�ΓX>T�	
�'Xr'Ȇ|��mA�NRH�Z�'�ȸC�M��]�B'�ܒ	����'�x��&��i�s�(F�
'+�!D��c�ϽXCB��4�78�&�CT�?D�0���VM2��w �B���MG�C��R�����U:mv�@�gJ��8hC䉶9˲��,�}���g䒷m_�B�	@�& Eݗ솠02��"&�"B�,R�j|¶� �/h�q3�M�f�JB���)X#�[-�hLPnهG4(B���@��_�_.�p�����C�I?<��EF�45�(h��邃oߒC�$�",����-��p6�^�\C�I�-��`g@2&%��cdB/�6C�I�y��<{��_'+�~���#�7��C� C��l9Ʈ�c1>�����=�C�:N%֍��J؟�H�7J��GbC�'6t\!A�� {M�(�VF�2͊C�J�!EH�h�Ab�=DRC�	5'.�0x0J�}W��5a C�t����YV��Ƃ.wa�C�	8i�ةw��40VTX���!�B�ɑ[�.���j��4́�oΆpW�B�I��`,�s��6F�,x9E}]�B��3Q�lI0T� >�@$ӕ���)&�C�	(eՀE��a�6g�r��V� �B�ɻ-����D�_�n���E��K|B�Z_����	V � 	яi�B�	�	Z�
s��KH��p��S��B�I q*��%@C%�J b�j�����d֫&��2�LU�d�sh�!�#g���A���I���Z��$
!�� d��sse4>����Py�"2�!�S-l��0B���y�gۙA�Bu��J��e������*�yb#Ե�h��`��_�h���I��yb��he�BK�R��;am�y��.�i*$��!�IA"�,�y�珙}Sb�N�/�̡��fÚ�y�!͇Z�u�ÄͤT,i:g�լ�yN�n���!4 �(��,�6�ȯ�y2��C1�B�Y�?Z���j��y��N<ܬ�w	�/2����Ŭ�yR�Z�#"�iŸ#w�х� �y��H8F@�qeŅD$ �aH���y
� ޽���3C��!I�	�9jr"O�(�����A=Ͳ�
�r+l��g"O^d��A6�����O�F#�,�Q"O�((��4�	��BV4<�y؁"O�����W����J�e�#"O(�0a(U8^�F�д�Y6J��M�"O�;0��%U��U�
�z�R(��"Ov@b"G�� �Rdν;�h0z�"O&y��#�0���
�C�O�أ�"O��J��E̮�����=AZ��""O��Bb�2E�%�E-��C�*��"O��Av��kQj9���͖z���Т"OD!����MR�ū�_��{�"O��hCj�����S+�9��Y�"O\�H��M�y1�i㕈P	 �z�"O�yC�[�i0�9���("T�Q"O"��4,���R`�@�~&��"Ox���f3�V�
�ުY�A"O@��Nؘi!k۶$��"OJqK��4���b�l*0�ru�s"O��<�Ԡ6
�}�$ū "O&���Pr��Q�$;���"O��ʁ"�YZ
��'O;��h$"O�iT�Cmg��
&�F%D�j�"O�����i,x;��X3&�݁&"Ot��ra�R
.����&�I˧"O\��ه1�vk2��
"O䨂�)3X�´i�L�>�i�"Oz���&¢�J�F܌��]��"O�����q��0�'��}Z&d9t"OX`��F7o� ٚ�nK�h����"O�T2ca��0AR��B�U+�"OX�p�̋)*h9q�l�*6��܉T"O��[m������l�1b�,;1"O�ô'\(Q"�X�W�Z���@�f"O���p/�	]�A��*��T�
@� "O
<`���;��苁I��5|��!"O|��嗹%ق��ް~��x��"OD�[k�H~Bt���l����"O��`���b�n,�E�O�� �"Ol`!��C=�e٦A��X�μ�'"OzD���S�D�	����j�|}ö"O��g�9ObZd��ޔi�d���"Oܙ�V�Z*@B�(A�|@�pf"O�MkC��T(�܊�i��gVP��"O��D��2�
�X��ڄC\`p��"O�J���G�N,i3%ڋz��(��"O�-v�كp6��b�M=�u��"O �ɖ�Ү7H�K��ģ*�@�8e"O
�P5O^�xf�[���::h,��"O��U�'�6��Ev80�0"O \��N]�b��QF���nat�yA"O�� �	:��mB�� O��w"O���	�r{��B�L���"O)IS�L�e�����n��I6�=�r"O�A�ԫ��m!��QVA#7)�d� "O��3 '�I�Q4y'K��y��F9�y�T�'�	�%N��y#��:p^����݊1�2x��Q*�y��A�$<����ۇ)���`V�-�yR�Ԗ'�ܡ)�ˌ��Y� D׋�ye�$'4ēd�V#\Jm��j��y2��%o�ٲaL�����ƀ(�y�f�c���䏌.H���t�8�y
� X��V1"����Ǚ�P�Z$�t"O�ѡ6ɀ8���C ����(��"O9�#���X�{D`��M��AI�"O����W�ƴ�&�~�d��"O<�J]�re�j("~��"B"O�`h����()�m �ג%_��ʇ"O��r��Z�A3�50RGڠyY:�2v"O&�)0o G
�Ȋs+U6'RmC@"O�5�fNG����h�,';�U��"OR�je��8�9�e#u'��"O2%cd�5�Nt2��*/N�K#"O<�4?N�Ɉ�
�I"�"OЈ�ϱs!l�Z���Z�<��E"O^ra�Y;qDpb��]�
tH���"O�	C�Qd��%(���ynj���"O����A���Paǈ¥ngl%AE"O�Q�O؞�,q��� ��i
P"O���u"T8K�Ag�ϥw�0H"P"OR�bp�f���bf��x��0%"O0�kT'�'��X��ꝧ d��b"O�����܍Y�hp���M�/�j`�"O��[���a���QৗI�����y�.�`m&Y�5�hy�� �y� d�!:g+*�~D�c���yb�4
'X���ꆼ���S6j��y"�3?Ƃ(���Q� �j�R6�H��y��jmtcb@U'< m�@"݅�y�.��Nu���� �
�M�WK��yª@5)�ʉ����|��(���yR	S�z �P3F�2$�(腧Z(�yB^�`Z�BT
���4@ЅH:�yN�=��`�� �|i�u�+�y��I�tJt�rˌd��l݋�y�ކh*�*���x��Y��bD��y¢��Fq;���~����ď�yB*��q�$`X�O%y`��D��)�y�,�"�8�V�j �lI�Δ��yr��+�~4��lE[#�$�"c��yR�R�f�"wHT<K��e#�d��y�dĄ|Q�M�$ӼI��҂�yb N-nyx�:T���T#r��¦��y��
�� 2��	>�ܱ���y�o��e�>U���F�/h��J�y"�ŗm] �E��TF�k
���yr�3 ��D1S��R�����b#�y���p�z=a�-�	N~�%�F%�y�e�j2�\z��@�8U1���yKc=����0?�\8�*�y$Q�fe�!�L�&?�"Y+�hN��yb�R� ��3���A.�á%�%�y���/(�05�T'�1{	2fH��yR�P
�D$���uȄ��$�:�y�Ă��P��䊯q�Ҡ:dh���y�ƍ+Ll��h�A) *~;V�X'�y�L]�������@�h����Ҭ�y�O�'3E��bF�f��HdL�5�yRL�,�yɢ�ձJ8��1����y���8(���T����b�\��y�oB�X!̜��獴�0��)Q��y� �4{��)Rf��A�r䨔��ym@o1dQk���2k�hqׇB'�y��5D_tAcCLҞ'��9X2,�y�	@6i�*���-�JX� �-�y­��_��P�!QLx q!A�y
� ��C��\�=���A��&q`��"Op����/_!�}�GN�pR�"Ox����L�L �`G�1A2 a�"O���&�w��"�� �@��"Ot���`��z�u�`%�%$���a"OR�jJ�
V�	��T+r�q 7"O�ْ��G�&]B��O5_�:-�"O� �6)�+�����qz~�i�"O,�)���Qv��a��'[c���3"O�L�U���Cf2!&��OR�@"O$���t����H��L��"Ov�
`�%u\�C���P��I0B"O�h�E!~H4�@�d�t ӑ"O(XG�L�8L
W�S�i(��j"O�<)W�����`�Ɂ*�Lu"Oh@rwF	8t�~���G.K�,ȓ�"O��	��&[*��SOɛx��%H"O��2&ۯgG�9a��pG8d�!�O�VL��0@�'Wn|Jwg�A!�$�8p�֌��7C��񡈔(T!�䔄6,���J��l����"�\��!�$ݥ���2dţ_z�=�i%s�!���[nm��ID(6��y{�*�0�!��]�&��('m�:�e�$�^Vx!�D�?3��4	����g���A��
G!�V3ܜXL��/���A6Y�D!�̔�٢4�R'yp,�4�,~�!�Dۄ/��aT�
��J��!L�Q�!�޸Sf��# ��y��\�!�İwz���e�� d׈���m)Y0!򤂉��}���W�$�聂��-
�!��>̪I�T�W+q� �¥-ɩEA!򤂯�H	j�L�2T~���N#.E!��k�f���c�ݲݠ��=M�!�$��>^��EJ'L���,��v�!�$)
܈�# ��-�jZek��!���(�����n��ԸsgǼN!�G�}Dx���|��)���)�!�D�����a���e��|�q�a�!�����D	2А
0aE�HB4d)�'�neqak��)�"p��!�#�Lɂ�'�Z�C���< ��e�3����C�'9�H�ę �����׭b\� �
�'X���s���v. �pXz�� .�y�JC,gMp�ʰ��� �\��(�)�y��-V���c�ɜ�-�8��f#�7�y��+���w��3 ,�ঔ
�y���8 
$`4���ta�G��2�y��
Z����,[/
�Q*�枥�y��Țk�x�P��W� �afKߒ�yr�� 6�<!E݂P��h�,G�y����Y��f��Q{T�"`H��y"�
@ä1:�m��HԒ���&�y������Õ!�)�n��n��yR�F��8t��ߑ+�!��)F8�y��[%j��Q��0*�|���b�2�y�LѪr�v�0�,X:�z�����y"�X%���IG��+�ⰹ�B�7�y"
�1z	�bυ�*OH�CP�۰�yb��$��z�� �IB�
(�y��G
`3Jt�`
�#�N훲�F��y2�X�,QDLcgV��qaѬ��y2��C�m��b��~Ab`QQn�>�y� ԓ2T�c�%�C����͍<�y
� ��z`�9>���X�V��"O@X�cP0]�^ ��e�`�XT��"O�L��Ĭ0�"�PWbݮ`�.x+6"O�Y�6��2�� Tc�"f(r"O���A�������#2XTU��"O�	a�Ο�#�Pj�`
+Z,�qk�"O���cH��8X:Q�
�>:L�7"Ojx���[�wx���$�Ujp]��"O��s筀� u�|�T$�<_ZĂ"O�y��C"���6$L����T"O
U"팯��}��	��ru��"O,�`��)z|���AD�!�HY�"O�dq��;X�ܪF�޼K�ֽHw"Oji�"G��_
0�ŋ�0����6"O�T�g�1۞-ef��E�&�f"O�)�Vl�!w�p T'[���""Ojb
�Q��X01[=N\j�
�"O*]sw��- �vH��Z*J�]�!"O<�M�?k2
@���#R�D���"O�5�( F~|l���ڴ?����"O�Y�� hu�-BVER�U�*��6"ObՈ�� v���R�!Z�7z�
"Oʜ{�ʈ*si�W�M�T�j��w"O�݁�N���30%޿H�ͭ_�<1�L��M�����ѓ{1ء6�v�<��M��nɸ#�)*�ܠ�p�<�6 X�3A�����	U��P l�<ɲ1���\'�Ƅ��j�<�v$Ӻ �xX¥S'B��Ń�(�c�<�a4z,���f�C+x�`�/�T�<�2��*#�R}	RǪ�ʵX��L�<�d��9I$� fD���AI�D�<��dńw��ʣ�߽<3��RC��D�<��O�c�v5� dJ*��I��Z�<�c	Q �-��LM�T|)ᄅT�<��B��V$��+A�x�jv�]Q�<1�kZ���*��B�5L�Q��i�J�<AE'�C��sG/��=�I�3�H�<���y?p�Е�F�nfj<�^~�<�BI�4��!���=���rs�~�<y'��I�������"A���s�v�<��%T\�rÆ R�&z��Ո�p�<�F�'���C��&�H��iOk�<A󊏉U#d��ԯ��;
4��q�<��OP�fIL�q'ot��8ɵf�E�<!�۫	>i8�[,t2th���~�<�퉆8�J�¦� 1�<eXu�{�<1�H59tP�q#�A�QP���o�<����#�T�9�4:�4��AA�`�<Q᪑�um@�6�P�}���v	�]�<���+&8x���78XL���\�<���¼1!��+��4��4wD�Z�<�!��O �(�ueH/[�8�D�^Q�<Q���m���	�@���L�<A�g��,6��vO�w��sE �J�<IPk6q�D�� K7�
�w��G�<� �l�q�B�62�ha�#ΐX�<Y�*O�kX�,���7�����U�<��L� =R 9���kL�@�P�<i�W-�LDؠj�>Ӫ�CǎF�<��� �������<��o�~�<)g�T"��w#]8��d�СD�<�O�Y����LP1]#��qE@�<r�Ҿl���%�PV��!�[E�<� vE##���^�P�&GF,�s�"O8�� �Y�D�]���)+'j��E"O�i��A� a_~�*q�O�u	���"OP�*��=�� ��@�%+�Fe��"O���)U�(����nB�b�6]H�"O�tЈ?+v��$��P꜍�S"O�9 �f�FW���#��n~�f"O���
D��"qrw�HW����"O�y�5C̕$����EXu���"Oly���Y*�D��r�˧#��L36"O��QfE�6U��Z��	8N�.@Rc"O��u�����h�8z����s"O(;'G�5_j��Z�FT4)��4	�"O���D)'���ZX��Q�"O�(�T".0\����G B3��`�"ObH�6�D�\�zk !*{2.�ɡ"OhX�Ϛ�@�`	�ވ{^��2D�X�bnԻS��]�v��V�@a�2D�D%H��<�`�ȷ�[M�Q�,D��hQ�'`�`@���(�=�w (D�PY f�o�nI�ҧ��	;�d'D��9����yBc��G��ċe�9D��3��͋*`�T����~�I���$D����g�:��y@w�U��H�n8D���c\:na��� Ճuv���!D�|QG	,��}��T�9/��� :D�0ғ��6�t�!�c��*G,D�pHF�Cw���C�����s�=D����g��h8�8�r��` JhIv,:D��#��^�D�ȫ"_�
�ʡ�3D�� ��2*�^h����}���.D���f���0��a�!ȗ^J(�)�"+D�����?��#@�E#�[�*D�@Q�	H�9T��ejF>lf�D�c�,D�,�p���%�|�"'�B:B�ZT�&>D�c�N	qB��P��5���s0D���ο\��E�Vd^�5T���I9D��j�n�;ɒ��D��%YF���3D�0�D�9��4"Tl��*ĺC�0D���� :�`0�W%�+<,fN.D�Da�m٭&�ݱ���9P���I�-D�0�%�P���F�L��ثGg�R�B�I^^$�hQ����X"R�ߴm��C�	�
z�,�rf��C]�$9��th�C�<dQ! '( �o��� Fl�3o�C䉩���W�\Xc��K�F *d(B�m�H�{�D�GWD��1��o%fB�I$@��<H6��,F2hP�ǄːO� C�	�D�|�
AkN���ѹfH�;L�C�ɇ���c3E�p�p��C��C��2<~]���CD�^��âC?|�^B�	0�<���iZ4�d�:�䀺ecC�ɫ��튖��^R��b� �Q�C�I�T�Hv%��K�8��_'`h6B�	�@m��s���W�+�랇L �C��=XR b����&��xk�)�-��C䉬`FR�Aa�@�~�|�c�ʕh��C�Q��9����fD۶�%ta�C�ɼt� "�>��c&�A:rF�C�I�~'֨p�h,"!dtٔ�]-`r�C�z)���<t�Pm�GY�C�	#m����"0�S #2!fC�	v7�E�bV�\�ʅ�r��B�<C�I/x�-�0勋E���i�E�i86C�)� ΍1@e[4Z��Y#V��)�촊"OXx҂�U�	8�`�a��i)�k�"OęK���g������f,Z�A�"O�x�F� [��r7�"a N<�"O,UZ3)½r�0��M�>�4�"O(��:ޠ�c���$#���t"Ob����ʤ<�d���E-�0"O��y��ߴ�,��� 8>zi@�"O�Pk���=j���W����[�"O���*H��Q1Ц<��Ea"O���bN��0x
P,^�	���t"O�y�dȐ��@�`�ӂSPPt+1"O
�W��1PU��o�UM$1
�"O-�iT�;�����W$v?���"Oh1{Ӂ;uI� �T���Yj}�"O\ظ�dդ%|>��"97���6"O��2��-ŶԚƠP
�^�XV"O�8(H�%�������"O�eB��]�nyF��z���ȱ"O��U�PA��2"�X��� ��"O� ��<0��Ѥ�h�baX�"O�Тu`ʗ�1�4��o6�D"O�{f̘�">� ��I�iH�e �"O<{�EL���%�[�PB�1�a*O>M���Q�#x|
5.Ǖ�i�	�'���RѮ�6��y��F
g*�P	�'0�%[�%_,���#�lH����'�r�1�o�^B2�X�G4 eJ���'4��pVk�!om����l�1|���O�<�T��	(a��H.�Д��cu�<�dQ�%H��xr�H�	��0�Gs�<I�1:2X�(�^�)��c↑d�<)��I9�Xrοz��S��e�<Y���e�x�s֩�N�P%��x�<���9CJ��V�w.�����p�<�fd�_:y;��H��h�Rl�<с��+s��H��b�7|���1�!WN�<�P-�#X���	O���`i��`�<��"����d�.?�$��,�\�<Q��Ϋ>�h��#._*��|J�G�T�<9EA�Am L{'��M|}8Pk�O�<I��W�[)�T�b�G.FN�<�f�Ĩp�ɴ���wR�{Y7!���+H~�b�dҭ%�\��򎄥z6!�$�x[��#ӫ\�7���P:4�!�D��,¨K�B�z
�����'�!�d�#YX(J��4_�:�I)�0X!�d��{�F����i�TY�hM�OW!��M3$iӑ`�n+���F(ҐB�!�E8$ȾPk�B��Pa�=�!�$��bD������D\3
`!�MBo2�0���u��+V�Պ}�!���&j��(�S�d�ح0�ϕ�%�!�$ȑ���
�(]�e�l}�c�T��7�
�(t�@�\�(�.T�{����ȓv���e��V�����(�.#P����s���{7)����"G��7D4��ȓ"��X��UE��� �Z��ȓz��4�X90C�YV�
��4y���\9Ѣ��/��u+��fE��ȓ~��1C�I�2M�e�FC\/4ժ͇�w�f}��Y��)���\�G٦ć�?0���EI�|\�� M�'�Z���������7j��E�� Vk����S�? l���@ߢW�H�����,���"OZdwҭ"�R-`ĥ�4���ó"Oz- M4\������`F�3�"O�DA�ҶL\���@a�r�[�"Ov����� x�SAi��"Oi#$�	C��|��F�wc��	T"OD�ҡ��6 �N��S�z� ���"O��s"�H$)�5�V+� j"#"OzL�D`]A:�YҪSn/ҽ�B"O@�ݦg�ac��æ,6N�x""O�������v��Al��'��2�"O�(x���;������Q� 	x�"OfM ���v��*`�g���2W"O*�����>tojt"�BY(���"O���h��wV��P�� ��9 "O����3`983@�� ��Z�"O�}��^&[Yش��NF-'0B"O�p!��7��x� �&V�"OD�#$=u�@���0�H�T"O�=H�`czhp��Z!7+��q"Ol��R������ef��DJ���"O6�/M�5��5i�ş�_�>�qU"O$ �����V��r�b�"6�����"O�u�qcU�7��A�w��<�҄�"O��S��R��'�/l��x�D"O��Q'!M2������M�`�TeQ�"OpM)�§)|�1�g�T�SQ��P"O�d��l)�n���ո �"$�F"OŹ��$>��"� u�u�"O�̓�'E?U��|�A	�i��x��"O�����m%
�a�O�5��YU"OJu���S-g�h��O� �rP"O�9�U�C L!! ΙZ�8X��"Op�����)��Xu�Z.8���	2"O,�
��/}��񫢢��Mu�}@"O�9ae�Ĵ/�������{� Y�0"OB  ��]�� @.W�u��X��"O�my2O���4i�g��.X�"Ohi)��_*(%��F#�,�;�"O� H`��N�`a�u�Q�����"ODL�2N�/0f��%ᝯ*}\�iE"OX���d@�v��� ���9)r|��"OT�; bU/�k�F!%8�1�"O|u:�Ұ6���Ӎ!$20���"O.Պ�&+�^a"q�F>�N�%"O9AU)�s/�1"���uD��t"OPxB#�����H��+ɒy�"O�Hkd�ȸ	����7�žJ�j��*O �c`n	��@�pV
ޤ �n� 
�'�nL�S�0s��<!uFE?/�@TP	�'�^ف���ɩD�*�bؠ�'(4L����v$B|Zá���di��'��u�H�?�H%���'���'�Ƶy����b���ᕟP��$��'�i�u�O=qV��a#�S<Ar���
�'���#�mKA�>�;{�hk@T�<A��jꩊAK<lZ�Q��M�<�FN\w�1v�:_F�Y@2�q�<�G�L4.hX��cQ�ry���a�<�u�8<�~�y�%ܿ��%Ѱ�E�<���6�Vh���>bGB�HT/E�<�E L����Eҽ@�(e�G���<YF���j3p����<��v�q�<��E3�r����^%�z�S��o�<� ��f�L��Y� ^u�K�"O���ܞ��P���f�����"O0Ř4�Γt��;2��SP%�"O4�ц�U;)���JX�I�q0"O�X�D1����֩"'fN�i�"O�@YpD߳+�t�S��j�-�r"O���f^T����e�LTl��W�'��Iަm`��ѡ`���/K8�X@�e$D��k��		it�D�]�<ל$�\�y"���~Dq��F�zB�@�F-��y�M	�BTB#�övjJ��R��yr�Z��X�$�J�o��u�`�,�yr���*/�5�ak��q <�P ,�y�d%l]9��ȸ~��	X�iɩ�y��]09����iϒv��� qM���y"�s�z��!U�pN a ���y�_�0��
�*N�%2���.��y���%��	3�K2%"M�cY�y� Ij�|�)A�����'iH��y�$�|����%�� ��Q��M^'�y�X.�������fA�u���y.x�04aULV�xTF�1Rʎ��yb%D;v�`�V�r�0e3⫏2�y��VF�[�lȮ�p�����y�A	}��1��f\10����!�M�J<��O���zb�4�����蕬<�%G��D�~:�Dܨ/2��{�؅I@0�
�	�I�<yA�Ϻ'u���Q�ӄVd��Rp�<1W�X�Be!ׇ	H�^�F)Ao�<i�H�7�������� $���T�<Ac��n��U Ԉ;�"��kx�<��I7��"�B�J$��Ǝ�q�<9pCE�R����dB�@:��Rg�Pp�<�C*F�2Ʉ8�PNĉ,�"<��n�o쓵p=)Cϗcv�C�DX=a��l�<IM��r^�pĉ0&��J�_�<!6��	�Ġ��ʠ��=GT�O���$ٟa^j|�E�{� �ђ��^D!���ĵ{� ւ\�U��Q+�	o��H����2͕��f��`���ę�"O� �DH���҄3,�`�"O`�!��B�p����bB�n��ʧ"O�U��˘�U��I�b{�f�J�"OT�X0˕�0p���qk�={��\��'Q��+qa2�9A�Ė
Nu`�#)D�Њw'�n4����,�5>�i�-&D�̠�k�!����4��TL�`��?D� Y��/���I� ��0��� �<D��C!� v]�8"��S����;D�P�@�͌b ���u�Ěb��I��9D�T�KSY�%/ͣY�(b���@���'���x�VI	|KF�`� !�Taq��5D��R�J�&���X��%�HZg�jO|�S�3����(ni�')� �8���.!�$��.�6�q,�*�轙�dZ3y!�dĔP�|`����'�V7M�W�!�d�V>$�	�
��5���r�!�A*2�h�V��'2�t�lK�w!�$Z�;GژuEO8��{�Kܞws!�D��o� UxVnߢ}j4��6��~l!��7�`A���bb)96=[!�DĪmLi��D2eq9�*��>F!��2S�PQ+E�Qq>����_�J!��
�`��E��>�EaG�Xy�!�� �qІ�W�:T
��CC�<U$z��"O`<yff�4����D!ߤ]�UyG"O$E0�A�7-8��� ìO�!��"O9���L�x,2���!nv���"O*5��(O�$����N=Vzl#�"O�YxSDB��%M��dS,a��"O��� �5 �B�U�Щ(:*�R"O�I5!ǫfC��� ���=S4���"O0��IH(]^�S���(5��@�"O.,� /�r�.�zc��p(	�"O�4��cҵe⪥��e�$yqt�p�"O2��CLۮ=�L{T.ۂF_��"O*Ey�'��(b$آ��[0q��9rA"O:�0í
1
�<����3��ȹe"O���@eϩ&��z0��-g��PG"O�:4�Q�7��ͪ���-Oɔ���"O���u Z�|��03� �x�l"OҜ
Ņ�>eێI8 O�!�����"O�!��EY�{r����3;�.��"O�E�'��Gn��Ph�b7"O|��ো�;�你�)�`R��H�"Op���j�]���q)Z.6�]��"OF�b�C 	�(ͣ�ŉA��|ru"O���T�
�yA����F�9G��yb"O�L!���F6�a	�:r���r"OP�2�&A�H���dܐ 	tQ!�"O����#D�e�� B�nG-4K:�:""O�p�-�)'O���MƮsH�H{�"O��§�n䈃 b�<`���d�<����:'�x�D�?��5���Q�<a��QC8� -%����CT�-7�C�I-���:Rk��R��)���f@C䉿!��"k��Aj�Q�Q�/e�C�I�{�T9��@��{���v��42*C�I�����葛\�~���m*&�C��)4�(Ha&��)�|��fk ��C� vHi��Ƨ�<Őe�ڲy�B䉚<y�@�#,�pB�Z��@t C�IΒ�A�`p�;"a�v���R"O�rt���$N�Ab�����"O^0s,�)x�F@S�'OlH�g"O4��T�8��@�A�^�N܅*E"O�eZD��m08�r���>�z�q"O�8��;?��L�4@]�[~|qW"O����ȗ�$��Qj��F.%	���"Oq�'K� [v9:f������"OX�j6�� A��X��F TH��"O~��'�A�r��&i��/�lzF"O4�J1cA�*QBah	�A&�e"Op�!E��	;�x�s@k%Ji��"O0���S�Q��4��(�v/�U�"O�����Q<�*�(6/�4h!"O�x�!D�f� ��q�N�<��P0"O~ S�O�+
��%[2N���s�"O����ʲn���!f��!�V�Q�"Ob�(v�C�<?�MU.Q�h�X�G"OR;d�ˤd��(5̀�y�l@�%"O����p(��Ȧ녵6H���"O�; lÖ{�D���'X0(�""O��ǌX�Q�T	ה%-N��"Oh�s5�LHS�,j&(� .�7"O ��(οT"�@��A�8��� "O�uRʘ��r8�Gc_�=�R�B�"O���$�s�H��睚�x�P"O� �\C���<�����L�\���"O�	�MF~�V䲄�ޠ��=��"OR��eA�H��c�6$�
��B"O(��#;���hD(L�e��|�"OZ�[�i��3���ֆ�<w���A�"O�5�ǃ�6}�Tk��O�b��
�"Oz�P.Η"��I�fJ �rQ�`"OHHc������g�G~��,*�"O��A� <����5��TK�"O�5kĎ!1Ծ-�����q6��9�"O���0hS�!�����D)�ȫE"O`�g�9�X�K�h����"O��`�.�#\��K�g@�Q�\:�"O��i��@<��8b�~�a�"O"qz�!�|���%h
�i{"O�S �Ô]�X[gى����"Ol1y���I���$�{���ҥ*D� 0f	�/$^,|3��H���%Q 3D�ذ$��"RH$[��DE��I���0D��s�!=A�9�ufȬ[9���V-D�ġo�=�L��"� ��"��+D���6ivi:��rDC�l킈1��'D�4 ��׉,xm����=�x�!w8D�`���պ�:1(��H8g�~t ��1D� �� �r��I�#�������1D�x�ƂAyn�j�L]='w�q�u
/D��3���>���1#��=&ˈzc�,D��A�^�X�hsI�	��|p�%D��u�׶5.,MP�/m��* "D�(�t��g�ĹK`�M<t��A�,D��(����	�9S�#
��ə@�)D�� �e�e����(I74X�]�m'D�,1r��v�M�Uć�fa��2�@"D�`�A�;j�h�BG&	r����-D��W��,9UF�06eφ� ,D��)��G�LnH�e�
>v�AN*D��Qb� K��C� .p�{0�$D�X���2g򬠨���g�H��" D��S�'�N"�k�jbꄂq@=D�H�o�PeKI&a�A�[/�eh �(�O�å��=2�=K��+I��M��"O2`[���z�S��ɯPޒ�P�"O�a���A�0��Q CEӽ]�]B�"O��IG��]$���FG �����"O�a�e/5�|�2'�:� �ۣ"O)!�*��.e`!#�����E"O�a!��'��k�ァd��%�"O�=Q�BZ�L��f� S4()�"OT�{��)�xaJ�D��@i�"O��0!j�je�E0'
5b�� f"OPT""�=!�dy������X"O
� �@��lzv���I[/�h)�"O���q�Êv��0�W�B?jp��G"OҸ�P��%�y' őg�� r�"O�-i��_.��t��E�1�`�"O���E��i�x}�p�*9{�$�d"OnY�&b��4��=x5U#sb�c�"O�X(
I�K2d �<[>��3"ODh�G
�6	�y��u8&��"OJĢ`!ܿ;:$�y� �ʈ*?!�M;g�,I�ӹ`�#Xjj4"O~(�'�$:�hy��.�xq)"O)�@�A�������Z��Ó"O
����	v��3�o��'��]3�"O� ؙ��B�o�`u���Xd��C�"Ob���U�ڐ)Hq*şmW���"O�T)TD��!����(J�3���E"O�������Th1o�H�i&"O���sE�L��D�D, {�T1�"O��ʄ�hj��(�TX&h�"O�Q���D�qтH�@,tx"O`�؄� ���c��._9���"OPh�󬋪]�@K��&m-��ɢ"O �6�7H��c��X70
�l0�"O�HY�@E#'`�`��mA�g���"OFl�"%�G̠9�M�8V���B"Ol�+���0��<¤�ЉP슰b"O�	�0CE>Z�(��D�G�V��"O0�(�V"�0��Q<��X�G"O0�!e�]0�-�̉4�$k�"O��`@�I����΂2���"O�-�a���"��i�ʆ����"OBi �����lrG%t�19'"O��B���<p�VhHd�	�F�R�9����*1�Z����I�=�J��P(_�D�({@
�({
a~.=x��5�:�b�ɠ��Z�4�J0c�%'L��i��d�%�O� �OiQ��*�#�
:���q̒:HV�i�p;ړl��`���~�ʿo�pE�����F�I�[ 1FY�?�4�zr�^�n���)��I<ba|r�\BJ���P�|���H&�5�M���Ȩzdb���OF���ܱ����_w�Z��n�0&�1�;	ġ��
�����SG��u�\Іȓ.�ZE�'%�?fj��(p�D#k6��kU&yXR�cfF
�mN8q�R�+�PM������ڴ7"��; \t��ģ�#&w��'�D�@	"�o�~=x��P }����aQQH�P4�49!���ԢT&Z��e
A��m�qC�x�N7�
~
��0��;m5�6h�gy���8E�ƒ)���9�,9f��Ez%�L�<I[�ԟ�b�C��4_���)�'������i����$��`�<�`B���|𰉆��L��6;O����`�j����t� ��dB�\o� ����N��Y�Ue�,�K�!��Р�����E߇N���ir��$d�Ə�/Ktu�W��/4^r��)�M���F�q`��G��MK��I]�b��rc9��`�����UqB��}�pȊ�EY 59~)�Ѕ�%�-��LƮ
X�h�cגS7M��$����e��o~�J�Aʌ1�n�sU�ΕݬXY��ڲa��([`�kE�'�9+����պT|��#�z����+Cm�Z�c��i%��k�zra��i�\ձ�NųsGR�A�#o݁��w�.dS��C	$Y��Js �)u�2��䔼	ܞ5�p"���aΡX��Y�;��X�㤘�T��%v'ZyK�XM&�Q�(z���m�=כ^w�09�m��z���VF�j��D�5|�|d���XK���!'Þr���ǆN:�=�,O�!�SM����Oy�5³�2Q/��a׏ؘA*�Ѧ�O�>p�"n��3��Hd5��YR�х�Pȡ��	�[��$�I��"�V�Q�Ș�E
�D�p��NQ(��(E��Wl�`�ձw��Z����T�������V	[�I:�O6���7.����Lg.���O�Y�ּe���0c�Vh0�g@�Zv�#V�2�*1�����d�4��UB��K�ZC䉝i��p ˦L���7o�'ZP݁ơ^��\�di�D�%!�]�\��˗Ē,��[`{d����@.&
�Ӄm��z1�dF�=|�j*O���GX���O��ٰV�ٝMt0�q�˩>C.(3c�5#�T�4`G�T��ҳ�C�7>l��bL�H~8���D�-c�D���R�dU�����"�M 5=�(A�a�V$Q���p�a�t�S���lI2U	���RV��T�%J4�N8���b�a�E~�9�%�F ���]#p�AvD�����SB���\�p�قV�P-b@i\!�M{F"^)�!K�J�*F,�Kć�a$�:p��K���6U��V�f�H����z����2�ɗK���R�+f1�NʼJbl]��)
-@�̡�a�%m���*��X<���键\
��Q�&��$y���ai�ۦ�SR�I�5S5γ}>&]i�9O���AhLa�Mȕ!�8$n1�v�i?���,���8,�I�D�������.B���	��K�6qx���_+(�T���ܮ9�'��h"����h\2�(@�!z�f�fBߒ��OY�`�'m����V �]�p+cl�v~A�&�I�o
��˵�	�4�րq����n�����4{����0�4��LA"<�x���*>~q���Y�4ڃ�'<tmIc
�\�
��Ts��(���Q,�.)��� T� �l!x����i�(�)$b�(攑t�ԡZ?����ÿ[��ٲa7�p��,�*r�Ҵ��FT�'4�4�F,X�h����9to�� �#K�l̖iRp$�98��Da���W�P�BD��&Bn��3I�'�6`�K���~b�HA6����d�ѷ�X �+�0	8��عE����H�H�Q�+縸as����u�
"H�r��k��ӋK�,(҄L�*{�%��f�h�$>W�4SVeM6�0<Q�H�<Wj�P��˭#�]@@��=%���K!�
ڶ��@��D�c���?�@��'	�Y���%�����2N#,1(�lB.�AQ��P�a}�DM	,��mZ���Ph.\
>򘽊7K�L0�� ɉ�v�ƭ�����p��أ<� xM���\�f|�0OЊ>��@�"O^�q��DJ����o/Od԰0��'�H�����oX�4��+	�J���움=q�႓�-D���UtlA� �E "~L��!(D�؂pd�<K�k�_YR��'D�l��c�,J�9�g��x�Θ�G�6D�8�)�=^����5ꊀQ��&D��0l޺H�~@2UkE�5�j�d;D�lr���� ��t"�D 7{�lH�&�8D���0I$uƕ
 �́](Z��9D�l�a�YPB<jRˏ��$D���7D������k�\�E� �y�XU�3D� *ƌ�:
�@��2���XƁ,D��r�� ��fDi��A�Oe���+D���.�el>0��
��|�I#G(D��j'���-�i�rbܧ}V`Q���'D���N6.L4�a ���#DeX)&D��Z4�<*� ,��yc��xPd&D���E�e�<9�NFڕ��:D�� S�ؙE�̴��DMw�HI�*D��qv'�%p�j�����A�f)�D)D��9L�)@`BQ��1A%
����)D��i5��^��3�B9?�"1�a�&D��vl̚u`@��A@900�[�`%D�� �V;�*��� ��t@�<	d-D�LHr�J�W�)�'h�4D\��D�9D��� #�8�`/�LX�l�Q�*D� (a�Ե#�:�ӷ��&?,�a)D���u̘Mb 8��/�Q&�zE�)D����6.�ne�%&s��uC�H%D���)�,���(4I��b%D����£g�����]u8� r�#D� �W�S�.��Qč�]�D�b7e4D�4K��H�!%����V�'$aǇ!D��9�V38�h�AG���R�Xy�!D�T�DA�-2�e�W�I P�8��cL!D��[�"aK���C��V���uI#D���2(��ڶł��1�v!D�(�6gޡV�,\�r�υ�f����0D����[� `h|�@�ːnxX�b+,D� �B(3٢��f����)D�T��,�V~�4�D�ԸX����b2D�[v�	&T0���R�=����$M0D��RA*�
8&dA�qώ2z��p���%D���o�mk.����O~ ��J�C D�����[K�hb�CJK4(��?D�0h Ɉ+v��PjW��=a[�Y��%:D�p֍G�7�`=aa�K�*���Y��9D���b-Q�p]`D�a�D�J�6D�x�e��1����k-c���4D�\�ԅ�F ��I��*�e)��1D�����P7af��Ъ��g��qҳ�;D��e�[&J�f���N
��Й(9D��Q-�� �D	�F�Q7ZZ���l=D�4#ӯUO������;l��|��7D��YFF�"p��ծM��\��m9D�,�rƂ @.j���P������"D�X���I:�lpA�8D~؀�B�#D�`г��J�A;��O�\۸8#��*D�(8F˔_1�!0��}^��:�*)D������u�FA��8z$��3��-D�����CUBeL7;��S��6D�@0� � :�hB�=�dE�A 7D�$�7�
�fʽ	�Y972UA2D�� b�f͘%`"�h�7 ҕ�����"O԰Q��Ri`(��Rmз��t�B"O��T"K�0bThƌ9Y���;"OHx��/5|�F�Y�j��(�G"OP Z���w*<
'GI�FA>В"O|i��.�p�2l�G�ڇ_�X�°"O6���陱#�0��J�o6
"OV���勮0���4ɇ�b
�u"O�P#�BG�%^����[��K�"ODU��@_	��	�';A�(-�R"O&8��7.CH� &@<u<A�Q"O����F�825^��d�!zi��)"OL�*5ȃ�Q����4N��\^ر��"O���"Դ6�|I���'pE\��"O����l�D����$!?"O&���J�4.�s +H|&lu�$"OzR�C�:Bb̢R���z'�`�"O�X�ץY��ĺg�V�z����"O��a�U��p-S	d�Ƹ��"O4�d%�'�^[Pd���:�"OP����q.�����۲9a\�`"O���"����m*�"E�
��
�"O�e�-�"B1���	=��"OF4�a����\�P	�'+p1��"O!��a��g�0��hB8Z�#�"O����-,U�RG����Qs�"O��bD�T�'2��g�T�3�ҙ;w"OF��eeϔzf��fÊP��x�"Ol��ᎌ�b80c���6L�8���"O��rf!��'`��+#��^���7"O�=��ɐ��4� ռ	u"O��rU�%��Y�FB(}Ϻ�q�"O�!�.�]�`���۴vTu)�"O8�o6���0�$Ԇ7�P��W"O�3�e�
n�2�b�4%$t{�"OuXƏ�]��A�RB�>m����"O0�:FH
�lzś�$E�l�69��"O�� �k1m�0�(w޷J^��Ч"O
	1��{��,H�`R$e4��v"O`���L0�6��A$	= ���"OPAIADԞc0�A�%E�ddZ�"O��`�2M�@m�P�F/#'��"ON	��!��u~@�A�!� ,8�!D�V[�|���y�ja����y�x5��)�)�~������yRJ+4_���`�%h��y�!إ�yr.o\�q�%i���A�iN�y�9熽�FH�W�ν33�Ԓ�y���;�.��c�F�9��)_��yɓ3`���b[	kC�]�A���y��	-
����'[�w��ӱd��y�g9�P�E�%0<h����y2���\��hڋ,�R!;oG�y��\��	P�j��x�Ѧ�y��Df��%��#�9e��Q�T��yRƛ1��	��N1X䭨���yb�10��m�p%�%;��0�/ܲ�y�(��+�:q��[2��u`�O*�yJG� Y�!{���.A�h,�dΐ�y�K�_E<Ec�)>K�l��kу�yR!ɡx�B	�Eִ���*�y�/�},F!Q��K�n����L��yr�;���A��U7@D�{S'4�yr�B"Y�ry�$HP�=�2j��W��y
� ���IY�p��$;��6!?���"O��@ҝ!b����	�_� D"O(]�dJ]�th޽��B�-0��*OĄ�b�{��A^�lm�*	�'��hBLJ9L��1W�\+X�0���'HY�fº��EC0�.���"�'.ʔ���H����E��<0�'xl�"�y��t�I8sk*e��'��ܰD�G�B%��mE's�( ��'Y��$P2_%�1��*l�^Y:�'W�y$m�@�.�dc��j�A�
�'�h��b!\� -n�x#Hˑ}�	�'���۴@�@1�$��3 ,q�'ZLxPs)T�C�0��R�M6.�N���'����m��xF!ĝ+l����'M�j'!�JT��X���'Ů�����J��:T�E�c�fi*�'�a�'�C���B�"u��c�'qF�s�&��R�ޱ��'�*�
�' q!�&!Q^	P�!Pt�N�1
�'��k��@^h��/ľtҀ52	�'����C��8Il�P�dƴl�dI	�'֜I�I�=	&m�"�0[+f(�	�'L���UM����B�#�<Ug>�c���L�v��E���@�N�n�s�@Y6 �Ԩ;C+C-�0?��ᖃ^8uڀ&��
m�Š6�ܡT�žmH�؁�Q[.Ȩ�'.��'�(O��R'G�4`�3'(X�j��@�I1c���y�kMX?����4 �c]wZ,@�"��+mў�o�6C.̩�L�iQHMB��xwa|2��.�Åa@/1�t<J���&�M��A]w�>���O�9�Č��U@_wr���Аq�>!�;S��ƁжfX�Eae�K�9����b'J� u�E.>�y��[ql@u36b�	W}HԲ ��N0��P�U4g @��;� ���4�J��s�MӃD��hC )0Q��}Lع�N8�O����ɜ�op�s��<a��)���E����AO���S�� ���sT�i������O������<q��O��q&�Ѳ@�؈ZK] ���I*��k(��Jn�������"m3!�~�*�$�5Q�($�T�\��j���*qE�hs�mH!�Q�1�A8���^(U���K5�ȳ�e�F��6�)�0�IF�?!���zܜё�ay�Q�aF�)Q�(��ߵbyL�[ǴlĠ�;E@X ��P�1��l��'����JT�F�����A��P����\z�� ���:=��Itk�*������i��j��8(�b�9���'/F&<�2�(@d�!	fha{��'���(	�R���8EJN�I���)w�R�;w�Dr@Q��@n�=�}�&g�֦@A�O�"�;G�I�����O.	��ȶ,�����V��I3퉨J�ry�mK`?��J<2lNU^w���Ya�SA�RmZ �Ƅ^,ȳ�T8} �h�'�tp�A%�=�0<YC��#�pF�<`7^91���<YaKǐ`&�ʓ�Ҙ��h%��� �'"z����W�5��t:��a��<��O<�y�&�,#��3���������I�un���">a1�"�!�K	,
�1p��2b��T��"O�{g�.�V1�MRJ����7�Or��j��l��X�M��}rq�HS<\��ê10�d��I�d�<yBNf�2�q�˅�Y�5j��J��
d� �;T
��0<!�LGc+2��v(1�	�<9�nȺ#���&�4�q�8�*$����SF5�X�/��
�\ݸ��]�p�*�HtO��@0���d�,�p��Ƞ?����`I��b������	�䔈h@�-c�<�p��'���we{��iG(�*6�X�T�� �t�hY!0� !n��Q�ō�t��:$I�5sb��4*_�X��6��]���&n�4����6ivȑv�&{���'��T���=���a�F\7C�8���I{e>M!sO��?Ic$`�����R�H��|�7^�gJҵ	C!l>5��/�����,ٓvk���&E��Max)S�~��s��ݧ5ib�b���MA"ϵwB����f�O���C�S�+�`_w�6�	��\'��,��Ʉ	g�M�gM=PjY	�`K�p�R��!�t<1��D&�f9��HW(v�r]10J�r�FL�A�W�H�h�7iW��a�(�&�h9�4�v�"��B��yM�'��	z��&M�n�"+�>��>)\ZF���%l���0,���Q� g�1Dfɍl��9Jc A�L<�m�D���IV�Ek(8��b≶I������_	j�H��Ɉ�^ &"=p��&qj�]���O�����-�]R&[6v؊(�$CE�6ifEP�"�<�mK�퉁K>@�B��'��3Kݔ2l�:�&��z�:ߴyDh��"f�VE��D A� H��:�uG�U�2��[F`P��� �T�U���5���9�"ߚ�|u"T"O�Pc�FR)K����kP�J�� ��J5Wh.����;�A���
��Ds��O���I�K��w�4x��&�Q3r镩]�Z�7� �O��@��O���+�ϐ:_<n����?��%��:0�����j2z��,���7�R1D����B��@w^�Y�����FbˤB���6`��;q���
n&�D:d�'�B3�Z/1q��PeB�:L.��	�'~<�Q�Oޔ��3��p�ԑQ	�'!yڱI	�/נ�����p�����'�,�c�B.ߖ��T�� Z�*���'�������}n��ĽA�d�C�'tm�d*4��L�`���AO���'���VW{تՋ��W?FH��"�'�����-��ѻ�+�5�x���'�P��#f�.�L!�,_Z̖��	�'4=K4cN`^Du���Z���	�'Q���U�R�I󸝈d��c���'�h�Cf'W"v�ST@�e�T�1	�'I���p��:UK���@U�B����'4�	)�g�/R2(�R�|Q2)�'>P�7�U�!�TA��
I8Xpu��'θ��$��.FdX�:���A�'�X�k3i>c��� Q&D#O�����'[��Uϙ�q�l� �S����'&u{�5�t��./x1<Й�'��� �D�)�h�g+�.|f��(�'<��!Y�MK��Y�
tމY�'�<�W)X�� ��#$�1��H�'� ����sHH �#�'�`X��'ZJq8v�B8�X"ce�pdIq�'�e�u�W,4z���Ý&� ���'�F%j֏ϐ(����/�."��+�':�1���<�2ي�G��C �(�
�'��@���Y
H �#HR;0{�l��'���{Gߤ)�r�c�EԬ(A���'�� ��PKJ4�%C��-Ƹ���'�Y��&42��Q��e�$&�L��'�B$p�Q����ϛ4/0���'5[��P?8T��A
ߒmNy��'��mW�H�X�A�.�7��!�
�'�ƹJ�k�I���3�r��x��'�a��V�$t�[C.��&M��@�'��Y# �:md�c'�3y�H`�'-h%�5�I 
�([l�a��
�'���V�,q	#ϖ:��0�'16|H���$�"�cD��6�p�	
�'I ��4I�1aѼ�1�J$zt�	�'lN`j���4{we�����H�^@��'���`A�Z� ��P�[}>d�P�'�|�%I��\Hn��-�r�>��	�'%��`��� ��F��l��0�'�=�@��I~~�K�*0a�=��'q�Pq���:u�t�դ�j�\Y�	�'���
P#D�F�4��j(x0 	�'�=�P韲g���$i��5Z����'=��[Q��S��9Dh��Xx`P�
�'ޔ�P�K�\n5³%U�_J�D
�'x* 񥢕�79*����KE���	�'��5nC�P��  ��t��e��'�2��#iA��@	��
�bHXś�'`���`OY��Ĉf�����'9N �w�ީ�䙉&�Zޠ�Y	�'9�d�� l%<qrJ�L���'�� �m�v=�᱒-�7l����� ���%� -�U	��P�bݩ�"O�%�)\�\�D�5�H|Z�"O��2��,>�P�c�
GS��sV"O���*�N��Ub[<|�+�"Oر��J�.F^T��a�J�	P&"O��b�ʔwp:�p� !3"Pg"O��06bIbل�����m#,��s"O��#C�%�1"���aG�}A�"Ob%Q�jǇ]T4�bb\�K�|�"O�x��@�����"�(L�"���"Od=�RDJ��^�҃��98
4"Oܠ��m� h�y�7��<�YB"Ox<�5��3hc�5@�'{l�ic"OJEI��R�b���cj�9]Ir@�g"OJi*�$W��㣋�hM9:�"O������v�ȡؖ �Q*����"Od�M�3����֪A�<<b`"O���D&Bdɢ� �U�3\�	s"O�B��:Vh�q��i.u[V"O�R�k[���4����#=�����"O�Œ �ͼ]@���Qj�7�0��"O@��oĢ��%�B愒�<��5"O����̢	$ȭ�OJ�2�=�@"O"؁�)Yi)���&]a�q��"O���䚚��m��,\o��+5"OV�DÖ}��LK���/c���#"OV�
���>��9[�K�>ָ�	�'��cc��t62�B���<��E�	�'Ԋ��s����Ekb�>5��T+	�')'�H�^TjiI�oW-/H�<��'�<��#Z}Ӏ������Z=��'$4)rP�˃Pl�$3 	���|K�'���Q)F,D�܍@!� ���'�Y�7G�=��t ��=bZ
�'# =(�슈Q"V�3�	�7`<�
�'y��ق�Q�/�x����7��y��'OH� ����'���Ht�Z?P|`@��'�(бs�ɾWZ�9��c������'����'"��-��9K��U�+k��	�'���ÁE�kv�����=c�m�	�'z��u`E�a�<XN26����	�'[�Y�V�J�	�_�'��J	�'����	������n$+X���'�DxQ�ɴTԈ	�GF�4-)���'��jPF��*��ǁ�}�����'G��I�"� s\<��"��s�B��'ol�	���8��CgJG�d��b�'�`�����3>˲h"tf˞\��$����,?т��+�d�/Y�6�Geb����N�pƵ��,�)?��yD�.�ēS|�ᓣ%�򕫄/+d�9�!-�.}�<RJ<ytc(]�\�O������� ��B����G��ys�!C�@P�y�ȏ�lqV��'gX�4�S�禁)� �B�]��M���PB_4p�r���y�0������|0��J��p`����1oF��@�G�Z�v԰P��O�>�ۓG�� ���D�:d�d��2�8��'�f��
�'+���zO8C��l�1�'��q�<�!!S'��u��$p�X����dX�8#�d�:�r�>ɲlyV.�D�S�O�.a`��ݹF��qu�_��l�q�'�ܙCp���ט���r�9��]+r��ô7D����Cر�0��a}2j���0|���\s2��+ͬt2�;%�^/*(Nl�%�'&<��e���2Eȋ�q-6�*�'��q�Q'�J�\���� �(�3�'HL�Q�ꑨ8X�uӢ�ʧ#y2�

�'~���w�˻��ТL��6��
�'�t���&��(V
��2��%B&�5������ �%������5��MN$=X�l�D"O	!��9nt�Y�i�+xpHq"O���s��r&�,���.E^�I��"O�!qJޏ~�$+p�ɣ5h�"�"O����(U�7'ޕ��*L�f��P3"O��m�{��a�)G�?f�tIs"O�CS�5��Y�HmV� �$"Oh�TM�ht��p��]b�X�"O�������*���]QV)"P"Ohu�peJ+=o�� �^�8w"OV�hХ�
n�]���~�и	W"Ot�� �ӯ,Gv�!4�ŷ\:�QK�"O�(�tJ^*
�B�H � 7����"O�y�b ��H�� ��p0��`"O�j�F�CԂ�@ e�-V;"O��Ëu%�m�dN6D%����"OJ@�4��:����Ƿw4�T��"ONȘF����`��$��Z �q'"O8���֭ݢE@��E���s"OdXB��(EE��{��G.1?��"O@�p�G�7UB���Y�x� r"O�&�r�� �e��0�y�5"OΝy�+ܐ&���d�z	 �J�"O0�z1�۵u�^���B����x�"O�"��_�vc���j�d���"O����q�:P�DIQ�s�����"O,��O��N�S�.<Wz�]�"O����+�W���zwM�V`���""O��)���44�q���a$l���"OD���#�A�PɱE�Ni��Z�"OF�`��<"G��&N������y�*]�7�"TrPC\.�:d�f����y�&�aC<�U��(*;�`�ݭ�y2��!v,��c�� -
�P`����y"��$	����"��)v��c���y��������۲j���1/\�yB`��*��w�TE��$Y�"AT)�ȓ6���C���1s	
��@��:#$\�ȓ���gO��	���R�fL:�ޝ�ȓ^�nmR���&@��P�ᗳ����jYh�ס:2)
S�_ߌ��ȓ�J8�ሞ>�f�8B'�.H0`���z��pR6�I�n%f���g&����ȓ$��̑ĬƊp�$�yĤP�r��q���X(؁`߇5�@�ӂ� �Pd�ȓ@v�#񫌔Xf�y��˜{y�ȓ ����W�B?㶭k%F��)�6���h���:@�TEyv[���n�l̄�%�\��g�kԴ|b����цȓ*�D���E�Vx"S�TqYFa��s|M#��[�<��Ԩ�'׺'&��ȓs�B�U�	����i�Rq�p�ȓ/�!��G"�xh��لz.~��|��ZE����
��TXD��wGx��`Pg؝	t��Vz�L�ȓ`=�����N�4}�u��e\	n�(��2^�G�,!����OW��4�ȓtXu��+U�PN�*��8*�E��30��.�9U�(�f@�59�؇������:V����פ �E��T��R�a��{��̐TI�48�P�ȓD���p�݆Y���9���V�B0�ȓ{�b�"��Z�e#�� �I�=��	�b�P��_ 	K4٠<�tՆ�S�? �\��F�|Ԋ�ba�$�@�R"O����W0+Ёi�N�>ce�|j$"O�����G�QH� ���`'D�J$"OP�aS���co�ajá7%��0T"O�#4�X�~�����()έk�"O���%.O�?��{��4&��7"O����@N}^�r�eG�l��8�"O�8�@ޮ)Hjq('C��xt�c"OjQ��) � ?LE:��֥"*�x"O�UY��L'8�F���nE:Jd116"Ox@q�H̱1v���M�d�B�"Oəv�=.H��C��)w���c"O�h���^Lj8t@��M&�`�"OA����=�h�Iu�M�Q�]�"O���!ʃN`1���)v����#"O�8s���	a��9�.̫8��
�"O���&��[{6ɤK�S+X ��"O,�:RB��PDAf��>5�a�"O�D�$�7p����L�?T�%i�"O�4��bI�5)Y���DnH�"Or��:T���D�p���"O��Ȏ^��,s�Dǁn�4���"OTi��g�:��髡#��'�<A��"O�|�i�*N��׀�U��|(G"O��0������.��By�H˥"O<!0�g߻2�m�b� wZ�k�"O�ؗ��,:�ty��˚*mm�u��"OΙ�a�T62��D)�V8o}\k�"O�ip��Q*D����D_��u"O����=x�Kr�n_0�"O*hb2�-M��T@��5�b�A�"O|us�Ñ�u�L���# 2<�u�&"O��(�KV3WǬa��R��Ds�"O��#���8f��ԫ��3�����"O��dhE�l�z�z��>���t"O��P��T�	�бcԲ���v"O���I���=��;8�YrB"O�̪��!Y�����Q�	���0�"O0 �4_p��m��'+%J��P"O�}
�K�/g����5! ���"OnDQe܈5����f	�0	���3"OP���ͪs�{��I0~ڦ��R"O� �� �������,#�xyb�"O�(TIĽH�h�3�Ŕ&{�RM��"OZł�\�+�Ij�	B /��8�"O~�¯�GU��҈ֈW~�=3q"O� ib�J�X�~	[�._<mn���"O�Up��Y�G���4-Wj�t��"O����)T�F�d��q��b��%x�"OX��)�ZjqA �Q��hq6"O*1#�B�6A Ū���V���R"ON)�U�H�'2�I8d'�2cD ��#"O�{0 �M�z�@�Ծ )��[�"O�P��mE�c���u�;#z��t"O��j�I�\u���xP�Q3"Oz0��@!q_Hu�%+U+`'@�:�"O�P˅&@�#`(1��̬�����"O���$�(5"�0V�ڑ����"O���v!��4m�4V�(�ؽ�"O�DX��I�b�� ��G ��S�"O��(2n�*���ބ����"OԬ�P�	)�A{'(W�m�ވh�"O^����G)Q���arg]#%|�#�"OЁ��e���z��Q�b,�|hQ"O� �\���G-X�(8x3�Q �4 �"O���\$/a��(���D7L�0"OVX��+�&AT1��-a?���U"O��(�둗Jy{ Lו	���"O�1��0�-��
 {��mq "O��a��Q�ɨ6*U����ە"O���`#׼9��EB��U�d���"OTٳ��_��M
 ��X��r"OJ�a'yc$�RW�L|��1���)D��r7 @�ыu.�p1�A�a�<D�$�E� �Dg�,qF

25���9D� �RH��%���E+γ�0PG�9D�В�b�V��!�%L�c�J�j4D�LK-�2;5�$�H*^"�7#4D�$k��ll�=�;&(���k�!�Č��R�k�I�c#�d�ւ�)�!��ݴLԼ����1#�j�#��fF!�D@�3��Xx� ��=ha��'>�!�d�j^xQ��ƪa�vu�a�.e�!��[�*M��枒J�JP��e��r�!���2zIc�B�Q�ݡPǎ^�!�DP����p��0H���H� K�x�!򄓆MdЖ�ѕ'��`3�͍x�!�dR#|�����`f�IJ���?H�!��u�������� 7�ͥ�!�s,�A�؎�,��E�F?:�!���D�[�ƽk�`�#L�O<!��Ix"DipL��0R��:=!�V�3�]� *[�� a�M�;"�!��[�Y+k�SŮ��ʘ�r�!�(>�r���͓��m�'`�8�!��M�.$\	$+ߋa���3B8�!�\k'�yK'�W 1`�B�U�i!���7�<`e�>��z5NX1k�!��WWBQ���ځ?暸���[L�!��U�"��N���� k��U>H�!�D��=�,KDA�h��� �Y!��Y"�!I?KǄ!!���P!���'<ȂBso�
��M��j��E!�d�����ã�ȼ8�<l;�N�='!�Nl8ԭ�����NF=VHM"`o!�\�G_�(�/��DD����6�!��\�gKN�H�"@�Jh��M�0"�!�$��v� ��s��U+�€��Iء�dN�{}bpȔ�M,��T��y"K��\Ĭ�G�(6�Y��mP��y��@��@�A�()Ò�����%�yR��R�_-@�A�ק/u�@<��x������%1���h���6e�Ny�ȓZ����@�
]����B�<����YYV������^���C�4���ȓlO���'� r���cr��@D�ȓ3��b��#��:���0`���5JlD���Ss��t��d�~�4T�ȓkiF��,�)���ҍۄH!��ȓv�v�@'%�(c��u�#���1D���iyx=U�J�!�ݡ�f �����ȓw"t�ӟٞ�����4F������S`ENa-ۧ'	�'�B}��!�| c%�[rʩ92�lǄH��:>��鱏��w�@�Vb�Z*��� ��!�$J��K`�y;&k�&||�ȓ`�왱U�
2�F���>T
������LXC�^8vU�H��V�'e6���S�? l�P��S���i�6f�8�h"O���c�A*V�9��Q�J�q��"Oji��:�� c�`O9�h]�@"O&<�C]�P�\��aE�b�y�"OTy��ک?7\�q��[�<ٞ��%"O
���-1�vBfB�"m�ƕ2�"Oxd)B�q�R�!Kw��=9�"Oʠ+��Q�G��a�˭<����"O�}s�GM\�z�a&�=�*)+4"O�Q����W����c�*3`����"OZ�� G��FD.�� ��#��Q�"O�tU�G�+��L���8j���rt"Oz�!ߓd�V����%���H0"O�$   ��ɥ[~�8r��\�H�0�=�0�a�Ϛ'�b��e�DM�I5��
��c�65�I|��ҐY�4(��!�S�8I �O9&�5n#}Ҡ��-�lD2R��G�8���V'0ȋ�w ��
�C͔J��p�EV<J�3��a>�T�d���R������4�FQ�ذ��Y�o���	!�,)�P,�6D�@ɶ��h��l $E���6H@�.���qr-�� A�Uz����ͷ �^�	ᕐG�r����k��t�0VA�F$&����+�$�H�i���B�v� b�i��h3�iG52Ol����j.�B �={]d|sC� ��5'�F
��d�W� 6��W51O��$��$;�呰�5 *�E0ȹ@
C�%V=���؁���Id���48sr�2{��!8 
	ަU���ڡZXLI��I�+�%r2%%�O��T+�7F�����ER?R�O�h�%&V+[���^�F�¥�ǣ_gd�b�e����l���+Y�`�]w�xp���6Sb�rE�v�1b��)������r�^����w�ح	Be#qw�4Q�n*���~����' � WFK�Qj<�+P�E:��S���7��$IE�@_�9R��Ϻd�J�K�ˊ�Wa �uቓ6B^������L�-�fE�-q�i��$�G���!c�	�%j���a�O:~�(�KZ0Ę<s�H+c�D)B��� M�i01/��NV4��p� ����d?�tQ0A���9_�[��C(޵k�a�04�F�X�^3!�x�9at$#GN�9�Q���	����c޴iK��	Edĩ?�B@C�'��3A��Dz��5&D��J�B`)���3�"mlXs���?�<��#R�
�% ��+B����#):$@!@� $��ᄜ=�0�*O���V�G�yRJ0O8B�jH7�6�z�GC�M֩��[��y2fX�Y��d�q*�c�~�¥�P#k�a��
O��R�x6� r�	�ÍVEXy@��G�b�z�����;��yu�5�OHP����;C'�$��C�:��d)ĕkj�cĂ��*=�9��I��E�BL�F���D)��"�X�=��B9�z5al�}�&�ك�J�ex�ڄ�'���a5)�-/�A���\�1�\=8�ɺ4/�d���S|�1sN� "t��S�B�5	.i�W 0�V!x��H�1%�L�P�OD�[�+�j\�\Hv�M-O_H0�'�=@�ܱ����7+s>8��֦,,��K�
ܙ[��I�O�����V� ��aYpV�9��N�K�>I8�C�;��E}2�'�h�)0�j�)Z��?a�	�k
�A!f�W��ɳN�!�r�A���M{�j�Mv�HN��u�4��yDX���7'�D�4K�˰?I��	n|}�'c��h/"��6�C�u�ԌPAF֔|<p)�VBC�h�:�dMire�Gc�j),��f�ʼs�j�-�8��4����N[X��d�',(��r  ��p̀���3�8pBò%*l� 	�[�$�A��� [(c�7	�t����R�6�"<���<����8���耹� �K��>QT ܌N�<��.ث
W�t)��A@��Ȓ�[Ndm�u#�h����T+�5�>9��$�X561����N����$�1.�h�P�Y wP�����]Y�	g��I	��iɺ����Y@�dp�Sl�9,��D�����"�Ѧ2b�< tĬ��a��x|�h"�'0�dP4lە�툠_`��QC�GŸ})�aڌb��9�I@Ԩ�� :@`+*�d� �[*OwhT#	�'=d嘓��u�f����/;�@��#�9�l)A'�}������������4���Z��ڐx�F�xV%P"QPa}�슠F��ĺ�O�+f�*ҧ�n���PӮH�E��͘2���#|�~B����A��V.]R"�ֻ�hO،�VF�fS����F��ħ嶹����"�aH =3n��ȓ(W %�b��['�t�!Z����3��*q�p��ӧh���@�ZK���vB�/"�\��"Op�d���2p`�����g�P� �"OR4����!�F`��HFU�Q��"O�[V���!�U��Q"Ot]���4S��@*��=����"OFTrE�V�3�$��@�	���PAV"O��3��j)��9t J*W�x8C�"O�d*6���Y�2�b�ON�g�FU`"O��[��`�M	'����"O�y;�-�,O�a2.��!.��G"OH�C@�<���!�
f����#"O�������9!5^�x�\t97"O�� C"'o�IA	�Z���"O��i���=@֤��K�$�0�9S"O(�Rhʃ8k:�3�H�(I��3�"O����E-�D���Fx|ɣ"O��t,�~��P��� ��� "O�d����@��A��T�(�З"O\���KK;=�eh�.s��X��"O�eC�e[ 45�j6@ZI�FQ��"O�!�J�IRV��&�Ì�Ҙ��"O0��f����,|���M8b)� "OL��T��p���T�!MPu�Q"O<Z��E%�H��e��)�&"O��"'`1Y�)��HB%}�A"O��@ġԸ��ݱW�y:V"OXt���9LcjXY͓(>���"Ote�%�ǿ#��ar3,H
ܰ��"O����2*�b c6*� #�`P$"O&��Pn��[d0��p��1<����"Of���N�E�b��[/YL��Z1"O0Uj���8'� = ���'�ey�¾�NQS�)��`Dp9�'��MI��.LV�I�ѨBg��k�'R �d�ɵo����
[M����'Ħ0��KH�	Z�e���L���yR��i%\��D;J�80�r(���y�F�!i32�h"*|������\8�y"���U��{�I�!p�$=�%o	9�y�x���e ��U��B��y2
[7i�HI�F�*��ы��y
� *Mj���Z`ĨK���!T6	F"O�i��#3w�r���G(S��=`�"O�9�� �w�I��7j����"O2m�'��d�n :� �S^��@"O�	�c̍�2�~��VA
nZY��"O�I"�Ld�\�࢏͘c�A��'�^�����c�I�6OD�pJ�ex���
j
<�y"O(!��"�t2րԥw�T�S��A����J�������̛��5ҧD�H<�Q�5]�،B���Y��|�ȓp��V�ȸ�d� 0,z�3��@�]ORqp%ϊ[K�(��~�g�w���2�Eus�h!�صt膸���;v��*FS���e�D�]"�h��iÿ�lu͎YF����v���km�5>#
�#�,��n%�E��!;��<���Y�´���Ɋo��Lˣ�]��T��"������%�J�y�ˁ�8���
d��D�m�t�;��� 1c^<h�/Z&o��a�E`Eb�z:����P�d���`� r��-"T�ՙ�y��DV���(
7z�(ţ�ą�AZ��I$�
6z�&�� a��ħn�|I&�r&�(��d��k�oܰ�gD/�O��9�L��SfR���ԎWJtH�O��a���$�\ـ�ŕ3č��)�|8�غ4�D�3��������� !*�'`��%�Ƽ"���D�[|}� B`����HA+~���	b	�*hZ��'�d��Pȁ�P�T��W�h�f�X�O�y�Z\�h�E��\2L���£�4T�r	.�S\6(ZՌŔ}ֈ������6C�I?״��G��i~i�$�7h���-�+}`Ź'�V&O� ()S��?ֶ����~kx}ڤ(�2d�]�o�l�X��vX��>0���䙾'yj���-��F3T}�V�N;�Dr�MK+�1�c�h��0��''��ĉ�NB9@U��.��K0�O>��M�J��s�<_GhԳ��O�P�5��~B���L���[g��t��<�W����А�LK>�F�Pe#H?l�H�F,H:\I��ÑĊT2��k����oƀ�˵D����� 0$�]8LMt�G�BD�a�IQ�!����a�/r��	hԄ]��I Zwrh\��˜�u
	W�@`���J��ޔ����n6�,$@���<!#K�i�f`qrhŖfY��AV�or�*��H�r_ZpQ��3f��֡F�1��\C'Db^�/�HX�`�՘VB��ӂ"�,��D�bkW�)~<���-�YK���������\���+z:���m؏ZA����/�Ո�B[."�����R�R�
FA� ��Z��OL�2Y�ըc�ِ���!��$�D�S��Z�"6AӠ�P�� ��H��sg�?i�*e�D
J�t������;p��֭�6J���0W��;�J��S'?k�$E��
ˍv���0�}q̭֫\nU1 �0*&-��b����E�W����Rr�'m�.b� ,�3+�(#v X�KW6�\� !�?�H�b�g �v�z�AӨ���(����+"v4g�V�2�Z��%ަla�YɤG����;P)� j[�E��ٔNx��>A��A��v!�%&t\jp�&�S�9���EC�-�< �E'l�2E��N�\2��ѽ��£5r�:쨁'O,�`��������z-��q�B�14���u����O*98��@<�C�Dal�/t&!8$���(�y#��p�05��[Lʽ#≃2�"L!�@�VZJ��5������M�?���@E)(.p�rr�]��y��7y���Г��- �h��́�e��K�;������ͷ؛��=o�jM%>m{�DÇ{�扰񃈋"�0�2�'
�U�_���!�Ȉ'�&�j ⋥�e�g�È:��`�創�R�,�-	ތ��@E�o[:P��-Ō��Pm�@D���c>�
q�X�ќ�1Y�l�v�B4�F�r�JȉJ
nX
��!�\�ൌ�!����$ �$a|Q����Z�^�B��K�3��@&%��YG/C�e):!Q����@qb"w�8�c�F�s6���#)����>d(�)V����V�PDPq�ٷ��$�6��r.j%�� >�
�&?��s%���pq�ؼ ��ť�:;Q|0��=��s�"^�V\���c�?�G��>R���ͻ?Q�5�C� �
*zW.��2#��3]�?3��P���tᤐ�S�Od�Ti��Y)���R�����0�6�� �-F��)��)	������X+���Fz"���#�H:����<�@%�r�R��~~X���u���)��8lڣ"�\bPO�:�^!�b%�i�R��O�A���hb��6Hًѣ�|���!�l'������	��'��D܁����d�����_/"�Y���O�aVj�|� �EbC�GΩ�@CQ�b���G�A_-&�Q���yf*
-_O�(c$�[�d�퉢's+Gʭ^M�,'?�iFJ�;�(�0�H	���Y�n#\d��CO����A�Z�%�*	J%�:�.� ��t��f�9H�VD�fG�8�qO�-A���E ɶ����{[jZW�7�ɎzYfbW- K�	8��O2 D���&L�_�x���h^�˄��i�~��m�*��M��2Hp�����I�r2����-�4��m鰣W+SnV�P����E]�F�A���'8pX[���,lP.�ЅjT�Q@��0�`ۦ"��ä�c�HA�4�%B�qR�q���[�,�+/C.Q��9F�H9��>F�Z���R �j��#[0��{���)+K>1*1�9E�F��nޭ��)׬rS�԰0���Z�A��-�OаyU�S,eNd ������N�u���P�d���X A�ɪ0�BmwNߏaDLH@A����:S�&q���%m`���q�E�>yHY0�87� �'|�@,]}�\=oL|�S��g�k���ng�q�b�L�S�>��wL0."�m@�H@�)��$Ui�{Č�r"�&� PF"��c�:}2l�4B�0$��j�3`��I� ƨh{t��O�tqsf�"`�*]P�l��F�:0��J�3a�="� ����I>`��%R<.l2�S�A
�a}��͂�):5C�)�������'*Ҭlqc� T>���r
�mQ�L�͊�u9�,u�J)��������)ڸ\���#Q6��34�Ř%t��0S��	Q&�,�5�5�CZ�q"g[�0c��Ebm�"��h	!���x�E��qs^%���[i1��"�̏ R��0W��M��Y����$��� E>�q�Yhd]d����%(�(��)�Z��8S�̝.EhX��a�U@a���õ(B+��HG��H��p��I�9Rrx�s$3���$N��G��e�>Yv�&pc">���N�nt����  .*�v�Q2ҌY(���F[��ן$a<��U�ώhy��� `�/�t�)�f����p����R�������� �IQ�V&�N�25L�ay����Df��%��t��!4�a�j�cek���a0�hFN�Ti�G?S��Xh��p��)DL�b�h�{�+���y �gU6>A���%�.�8�9C�޷ψO���'	 v��0�ea�&<d�7�sӺ���)�{�U��t�Htqfj�l����O+�	7�E�a����ቇ�~�7M�� �조B�Օ9>:�8s��l9� ��Xr`X��A�M8��͓R
�EZ �FR���˙�?1�@�$]xtp�a��I2��A�oJ�C+> �pmJ��J�36l��1��C����(��d�DP�fM7�BTP�/��Ol��Ħ��WJ��!h�HȢ��Ho.��X*�6=¶K��+W|���3R䜁"pҢn�T� (�JAJc�Yq�� �����R��sQ����G�TN*!ځ�I�3-�eyscV���d���|���
V�p`i��KiD6|���lYq`'֐�������&�j��p
�wbq�4S�R<�ȃ\ T�X��"�|�F|r�VY]`"K�(,q�BT>]s%.K�p�@��'��$�4U�t竔t$f�{Ra
�D�>}KuN�ǟX��"��#t�r�}xǎ�1{d�(� ��P��4K�Ȳ��;3�Y.����dYD�q�DQj��� OΑ[w/�=缱;��5x�x!R�M�����n�:S���(p��6ձ�
�<丹+��DO82Μ��DΨr��+���U����1�OD��p�ߠ۪���`��yb'T9	E�␍��px�ͨ�Bɩ_$�$��"پu���#�R?r"������ K$��CW�'�̅ ��V�m��	�'�,Z���xV�ֺ?1j���c~݊Ս\�f�j��C#�?��HW/i�|{�k\7�yK���M�೗�� �29���7џ�k����:<�������.J�d��F��~\��re�@Ť��T*�k����w@D-)_0�XdL�/J�l��6�[�} T��REB��5�˒
Q����v�÷Q���	��,&�'��R�StܓS���	��$6� 蚩+
��وS���u�E>N���o[��x�.[^D��id��(�ۆ85I��	�{�f[�Ϟ,N��=�GOMɚ�f�><�,��@/ۍa,��#��;l�ԓ�愓_�����P*-V���"�(ZiD �u+��z�
��
�b�B ���l^lA����6���
�tw�1�!����(CMO�d�VYק[!mTxi�`�7��"Fj�U�$�p��ڠ/�Y)��ap��YO�(���s�5���ï!P�@�b��<���9׌�1 *�:be�/D�4�M�w�	�'��-"U�L�9�*��&�0"���� 1h��X��'64��m:�ɢ����ܘ?a�x"u)5D^��!BA�yȍ��H%W�Pl+�[#���g�;k�LZ���7@Y��)O�tY�b@n5�D���&�8C���I�^��!�	jl�QFB�W~��XAeؘRE�8qA���@3�g�5�j�z���:MDH{q�6Ft�1�d�B�-ͻLFJ#?i�j
[������S�dvVM�S�T���X�U	�]!6!b&�U�>�\�	Q*K_������"g|N}ȃ����PAe�\5&�Y��N�}�h�k�śP��uHC�'�E��Y�M�HUPK9L乸�!6uW�Y�T)�P���Ф߉�}k7�%L�La0�눸Jaa޴s�.��Z$��ڶA��:�<�k��F؞���_������S�+����׈G�~��s!,P/`:�d��.�}�t��w,������K�H���W�Fx��#��.b?�p���j� v���smȱ��TvD�>agD��S�d�1�Yg�a�!FsIH�IըG!.@=:��B9yO"չv �\��*Eh�"a� ��Wdӟn�1E	�V�L!���(C<�)1�$�L sQ��p�ā�ad��ڪu!��E2S�U[g�*J,�A� �\K!%ܶt�ع���3z^����ڣq߮5���T�X0q�GE��p?�wl$�2�����5�=�'��iz�IR��Q�A� y��� M.0Y"#�m02��$N��y�O�=�j�� ̊n�0p��������1)�aˈ{*�<��S�~s�����Ztçៗ-؞�;�,P42�2`�7}�I�r�8D�is#آ �JT�'�^�.ގ�k4����#���4$ZV��\�EJׂ7}����$�T����/`vT��0C�A�@z� ��J�R��`#�BطE/4��W�\�c¾ั�3'�Y���{o�Mq�K�	z�<C�%�8���@�s�$���Ev׮��%� �
���G� jBJ)��K]T �aA@{��d�pܺ�D ����h��O��DB�3��h�ւظk���{R,5D�@"� &a�%>%��l��`�E��l��1�t(�u�0���>q+@�`�(b�L8i�i��؍ ���@���AHǳ< n,����f����V�z����y��y��=��(��B�ab<]�g�R3�v4H��؄k�T�1�S�~�(]Xcoǂ&�E�6N�7�$q�׎7�|8@�`X�o�ʓ~}�a%�_�z�J赮˻&�Z����O��'J�Zᮔ#�*|z�9�E�=}�^�� �P�ʇ�P�o�����b�I
�"޺ {TA�F�ϋ)���`fiQ$a/��Ud�y�����9$�Ȑ�\%jO�!�d��)"8|@�1����A�f�ހI=ҭZRC�����(��iH�����&0rT��PΦ�gf^�j� Dį*K� D�W��O�g�M>W :���I	]V��O�.�uC�]��%�0<j�@�����S2���u,^�d���FJ�]�&�]wpr���Z�.��ҍw�}�� ?z�@�٢��w	,���f���7o�
;V
@;C.@8^p��~ZP�<��	@"E~�3�H���`UB1�݋�T  !�<f�P��,֥�Щ(��Cj�s�ቶ�d��p�ޚg��恋6͐}#q�ih�c�lޢm�(q��o :�EG�2���qF́e�=�f��L��� *�����ND5$�4 �(0�aA*��:� "j�� �%��N7[�r�P�ÏM]���Vb_�(��`�U)F�r�,Ԁd囊l#�	�bL�����K5�N��4#�t�a6�M�����Ai	�&�8Ez���a2�s��\�P�ě��C��v�8)# `��P*�xALY�+��koӲ P�r��S�Ȋ!(!B�9t�0%3(OD$;��Ĉ�y��-T�.������Q�$9�M���_�F�YD��4nD�1w%C�X��A���A�i��v^"��U*�� I<L�����
��0D+#�1J�dåx_���ԛT�y���8g��ԙ%��J�B�Q�[�="��s�hKZ���-�P�M�sb\;g�����E�N��.?;]����Xm��L�#�o�a}RM%o�XM����
P���"��,7��j�,CA��`�O�#^���'��*�*XXd�P�T��� be-{>��:al�D���B�6N�0+�;v��D!��Q[P��ܒ���Qȅ��:UN�bp �-�t��(U���ic�G�t���G�� �@��@�7rpHw�A|]~-!"H�_�'���@�/+���f�;�.����Z����K�hNna�s�Ҹ�����ά-����޴uNMߴ.#~/�&�k�S�b��-���M� �5�'蒾ǰ?1e�4H��]�Z!�|1!�7R%Z��W��7O�����$ ���
|:P�d�ݿX'�`B�P��3$�J�%�#�٢*F�
�Bl����3�֠k��"�Y��	�@�9O/&1��T�3�XȘ��'����0J�\����X��%Yb���I"<�'Xh�M�Q�2<�ǂY8U������N����oC�|-����2<NX�B(
�]���ʍM�!rB(��N-���A�$ު���mѢ&��@�Óp7JT��%��y��-J`���&��'s�ŋ�����vI��,>L�2O�|�9��������ƉXPtӕH�@v�j�/�y�r���%%$�����%f9�s���8$ʣ�C�\|�IJP`��>��`��kã>)8�~�Ʉ~�.5J���"Ov�a��Ž�>B�ɸ^�����oΚ�`�H��or:��*}�༡`�3�T�F�?�=Y fKk����S�z|�C�,�fX�z��O����N�Zuh�Â�� д��d_@�0�e�x����A)!����C�TW�̪�l2�I��Ha`*ȯE�>� G%5�&%̮����֜ �E
�a!�Z�r�� B<��i-W�@��'o��0��,OajդO�>����֣���
gJf�z��,0D�ܡc��esHIA&휱6�\�Y�I1D�`G%W�G_�{�HΨa��Z��,D��xW�Rd.ԣu������WM,D�,*�DC"!� �4���H-D�4�wD�!cl�]{�@�Of@��s�-D�P�'�͙��
Q"�0,��0�1D� ��̛)rNm�%cٸZLTu�3D�`T�A�@\�y�GQ��A#4D��ؔ$_�� hIu��6�(�@�O5D�D�VeI� ���ڧk� �HQ*�.D��e�[#m�8�
�b�8t9�"#D��ik��R�����	A	�k#D�< ��	;����*�;|��"�7D���$"Nz�H�#S�0���R'8D�XKbf�S��T�\8@bƔ�$O5D�А��˂4���Q�H؁f�LCW�$D������Z��3(
w����D D����`޻��L��a�_	"�j�#0D��; Ş�i``�$�|��]�W�0D��(�ke4��95<�{�d5D�l1w��:��2.Y2Ҷ�Ď1�*�pĘ��AqT����5z���xI��	��I�a�F���ϲ1=p����I��'<r���S�k�<;V�E��T�`���x&�@����3c�Z��!�i�4�R>i򔏃/0�ಁ�G)� E8q�ҦO�:�
Ӱi7���2] &�]��=]x���e���NH��,u��ە�i߲�'.����'X����r._�L ��S<{
���o:}�i�'x��'<����7K�ZIR���K�t�O±���[��1 J<�"��8pYI{R�����ѥ�|}"h�B������)�'&�LQ�!�;>�@�+�8w(m�)<`�f�G0�r�S�Od`XC�L�
U�!��ա��u�Q&ƵT�Fݩ@e??���Ou�|`Vk�5m�Pm�&��
u���@��f��`����O)P��&��$�(נQ�����R�4���-@��*$'\���D� Sߌū�M<�@����Db��<Z��ti��KD��	W�5���pʛ���P@f�д"68�:2�:��.M�d�I#b�,#��O�>��/�o��aZ�fL1W��BP�i��A���\�LJЈ%�"��.�Mr�����w��Є��^R�\s��d�V>� �b�뛯���@�.^�l	��dŗ#Z��8�kW�$=yK�+@<L����x�� �O����G��:�~]
��?��2��A<�?��ϗe�)���2�D<� ��)�1x��iS�Ū����77
��c��I|bX�f��~K|{�'�O�,��ӂ9�H�����8��1 ���)�b�4(��N&�ا�O�N��D�H j"�u*bK��9^��	�OF��D��R�S�Oyn�9��ק[�%9���+�\D�'�|y�5��>��<6�F�D)A�
X���*�\
�)a�Ƽ �6-��<ѐk��%#�Ԑ4����(��O.���pj�-���Ѥ�ާ<�4�*	�'h8���*oW�[��� 4˲�	�'YD�JLQ�j�g�S�>N܌��'����M�C��l;Kߘ�
�'�T(�s�+*��ƀX�?�U		�'�"��x ˵ �c�ݑ�'��	ӱ�ܠA�t1
�f�]�,p�'HRi��ّvT.K��/P�r���'��|�cm��*}�p�X�$���'=�\��F�]s�Ժ������$��'^����AI-i!���!\)ު)s�'m"�)��Ӎ8�@]j���4t[�'z��H&�Y }�ԁ����� hc�'� �4`��|��y�
�[����'tl!��k"me0L�p�\^���'iTh:�AD+(}@:J�}��'���!Dė&MX�A#��+�@���'R����3%�����F�0b�'I�{2܏Y�N�2'KH�!X�'h��"�ח��0k!$r=�'?
a������JA*h#t`#�'�X����Q�X�ҩ*�H2[7=��'DP�)ƳW,RiH�F��W#`���'ئta������C��Rv"=�'�d�ui�>pv@�e�K�8��'r>��ф*v;��p�	�p�m*�'�
 9�N��l�ĥ��˟;c�p�:
�'�u�Ҥ֛]�������]��q��'Ct�������gQ1h�S	�'�FS�o�g�M�r�<.��r�'�4]0ݨ2�TabB#ҲKZ~q�"O,0�e�˯pP:���"�#V9��"O�-���E�k���H`ᄑ)��X"O��fɇq���t�"��A1"O�,�`%C�?%��8V
�'�4Y �"O0)��57T>D��-��+�"O�u���6�
Pے���xc�	��"OQ�@�|됊I;4]41u"Of�Q�^�,�����X 6���"O ��L��� �s$�������"OV)�t
�' ��!���A�����w"O�4賄������o�D��"O���p���(�V��a;
F��P�"O@��c�*��ມ`Q��v�Z�"O*���	[�B��to�$#n9��"O\��u�ɱ��������|�"O����B(�����N���)�$"O��WLӪq��ۧj
VH9�F'D������4�2���BLѦ�$D�<�A��n����e�%0��#g&D�8xP&��{hƽ�Cb�OT�&D��hF$*)t4����%,��|���$D��:��#L�R�$>H��0��$ D�����Ye���$�|�q�҈u��C�ɝrV�I�*
+o���a���C�)� ���>@A~�0�O��l��"O(dm�0>�VL�d�	D	@�"OjMK����C:�{�CYx����"O͈��Ȋ�]��GWpI�"Oj�I�� q��R� F�A��y��*;H~M��<y���F���y�*��4�a�af�d,�M�p-@<�ybL�uO�$ZUdmwz�#P�:�yBd�b4v���e=]�)�r	H��y�%�o�hYk�m�1X[l�٦�I�y�NX�`@����	%T�@����!�y�Y�O� US�O�+M|��q� ��yreF�����[�t�`r�@6�y�iÍQ Sg��0u?��k�៷�y��U^�މ��U�f��<�W@
��yb
�?'�tmR3���Y����UIQ*�ydS�c�T%+�GT�A�~U�U��yrl��0��zDkѕ�P�c"ܘ�y��`�.M��� ���i�n��y2 �	��P�-�1~�)��'�y��b�݃��T�|�ia�$�yBnƄ"���b6#�UV�ڵ���y�ḽ}�v�W��/D|	8"��y���#T��C�b
2���ю���y�\�M�����N'����Ɉ�y"��1[��P���G��M�` ��yb��)�rCÌ�!D}\�b��G'�y�!@�$���s��>�1e���yrG�l�ht�bZ�7�*�#%�՞�yrBM�13�d�)4ɐh�t`_��yRM X����Д)�>!4�
��y2�02ؚ��dD^-�v}�S  ��y�@'T�sEC����$k�y�_��T	�"�_56ڀ� 
��y��
.�������,~|2�2�L�yR��/_[��c�"�u�(�P���yR��134���%M1tN�C��W5�yB�D�l����ch�U���R��y���;G����'�[%l�I�.6�y� ��k��l��T�?|e�G�ɂ�y�ā�b4���R���I
�y¢�gy���G���#W�@��yR��qZmiA��SA��fB[ �y�Uvr���͚Q�$�Y���y"'*��3'M3DcJ���ȇ�y"������w��04�<�1��В�y�/ǹ:l����e- b ���%�y�&Xk]>����6� 5�ъ�/�y�C&T5��bΖ1 � ����yBK6>pZ�@t�
�HZ)�II�y"��~�l����C��5� 1�y�B�	:h`�g��C��	a����y�)T�4�l2��x���Y��y�N+e��1�o�>^Dl9��P��yrK�����@/@7&V�4kg�6�y�"H_�t�@F� �8�SI�"�y�gV��X��a�1}�d��@˔�yҋ�	�J�N�P�낉�yfƵs��se�z����� W��y�n�,��m��&�&$���sa�#�y�X����&��2E@��,�y�
�:��(D�"YUq5hY+�yb��&w	J4��,!kc��E�y�B�'�08h$Ƈ�oox%�e�y
� ��@!̗H,��G �A�`��"O�x9$�V+b��а�fMe�R��"O���@�1g<v���fџ���"O"庳dȅ/0�"���V�$�"Ou�fiˆ�<�+C�Z*p���Ӑ"Ov\�v�B��m����_��ti$�%D���hL/f��q��~H8Vl$D�|�o�.ki���ט~n���/D�T����/'���H� =gH�S��/D�\�D�!�J�@7�Q�A����+D�P
˖Q��zF�ʊl��j@�5D��[%m�~Y��B��/n��5�S,4D�ԁemW������1t�j!7/D���3��f��,a�Ǔj� \��+D��x�`�]D���� F�BF�y�$*D�಴m�;{�J<�g�!���J�&D��Kf��8�n�x��N�8*i{cI$D�8�7Ȁ3 wr�{���$5h��.D�4 �.U�M���C�ٺm�J� �`+D���3!�t�f�"�#=��I�"�,D�Hx��h��)�G� ��T�&D������@�4�QFɟ2���2��%D���
G�Y�HW��v~||�ՇѺ�yRۄm���F�ގ7R@ �Da��yr*Q�DѼ���3+��$3�g���y�Th��9�2���l� ��"�y2c,wHj��QD�{F�R��yb�Q�n(�ǎc��R6�Ҝ�yRʍY��8�
�	Rx�z�k��y�e��xJf�sAW�|�@�R�ʆ��y�,GbJ����4q�z�3E���y"鑇:� ��`/ZSV*`s���8�y��� ny�t�T�����yR!ˋa�(�X%E9"eXY��A��y���6��a�� /NhDKր�:�y�$�����ʂ%�61ji;N��y�ș3����n�5 �VQ�O��y��k|�A7��C/���TA���y&�&��}@t�ׁ����Oh!�$�w�tU#���=b9�De��sf!�$͈�P�H�F�+j�JMigb���!��6dbQ���2LԸS!�.�!���a���(%�-cY�ӯ�!!��'����Q�T�Cר\�3�!��^ qE�eCf$@�_� 	��
�!�$�$�z�
�ؑ6����qd̹Y�!���_�n`Jq�E�d�ȥ�q�!�!�ŀTr�3�.A�kz֝��A�.�!��̘5KrX(�Kȏp@<ib�Z5'*!��j,�ó�F(}l�x����|:!�DX1X�6D� }2�X��D�8/!��ΐ<��僑��$t���ĈX  !�$ϏO��J�^������;!�D	5�Aj�/No����N2.!��1h�HI��P�\W�	Qƨ �6A!�D9e�Pr�$e�8�v(rA!��ů2ݴ`���M�Y�'�Ȋm!��ѣE8L��Z%v�E9r��ti!�$�\����uZ(A� 	P�!�Q1�� ���S
fy�e��('�!�D0����O��(EiL�!��7i�Dr���J=�f��S�!���f��jM1z�(��Ȉ_�!���6/�`tn�[���[ǄD�!�� ��šK�s	ZDKpj��=;�s�"O���Q&&�,j���U&�)y"O|QZ��8tu���S��<@�B"O�I撠HBH�tLI��ƨ�4"O��'�ߗs(���*9��_�<�f��D�dtI��ϼ(��T!M�S�<�S�ιp��5GѺ,A�x�TJ�<�6OӍp��q���͍-g���b�n�<qD�+����İS� <�Dϓl�<��D"z7N 30Â�\���P��B�<9V%�������,N�T=`�*�~�<�f��r���D+:DDXK刉u�<��	 Jp��l[)3� �`u.	s�<Ԭ;t�b�h�"�r�J��l�<Qub�( (  ��"O�tJ�N<���2��A3*f��7"Ov�2�@ǭ'�����Z�L�zD"Of��Ek]�gj�����F�� ��"O�X�oǀ>`z� ��>"׮��"O^Ń5��:j����r	�-t��"OJEa�
/�\D��@3`r�!�5"O�x����&�\����W�Yk#"O�4��o�EМE�@��+޾UI�"Or#S"R1¦@ZS@#F�,�k�"O�����G�<����T ���y�"O�(���-f�m��@�(�p�!"O" J2K]�}q�� �y�2P"O�\�u9�d���nE�;��`P�"Op 9��յO�1�P��/(��L�B"O�r��V�|�� 8��4*���"O,e��R�2�D�:�gN�m֠�R"O>�ANRx�JA�c�E� �����"Oh)����*O�X��.G����"O(0Hd����J�ɵe��|��H��"O���,�.0��|+�Cȓ%����"O��a񯟎,�虲��`lJ��D"O��:���6[��� M�&Bb���"O6� �L�"{��m�� :^&��"O*�kǗ=��u�%E�U��2"O�!I'n$�Jt\qM�ŲQ"Of|���YKgޥ���8�a�R"O�<��g�$K�-���TUy� �"O�mPp.�tb�Ւ�V3Nu��0�"O�9��	�/r�<����_f:�y1"O`�2�O�|q��@��ƨk�J@C�"O�Փ�EýU�h`�eg�23��\`W"O�t�v�T�Dp���@$|�B�("O����/F&4F�\b����%��I""O$}
��٪3X��ȑ׬��§"O��)sH�����c��&}��3"O��ٖ��8�	�id��s"O��TET#:� rcҍN���"O܈
����5��0����[�H}C�"OD��-�Z���lR&�5�W�*D�0�A��~z��� R.SR$�w	#D���
�
'�������b���?D���6���<'�VoH
7SUǌ=D�Li�ȗ'h 6���-)?3m�B�:D����k�=V�q+�¦NQ�E-D�Lc��pDP��"X	�B*,D����f�H��!f�:"䐞y�ȓh��P˞z]�̣0ț�0�0�� ܎��T%��3����3k4�ȓsh��y�$Tiݢ,�BM�p�Hd��d+����"P�7��Ak +C<��U��o��dr4Oބ�h�2���1_���ȓ)�Nl*V�$�a���ų&��ȓ&l� ���B�@����C�R����� � �ӱ��8�D'�e�|��u��ٓ���4k$���l l�T��:=����"� ����@�,I���y��m�9A<��1�Xh��ȓ�M�qAM� &��g�V(�Ʉ�S�? ����BU'�p�sG �_��0H�"O$4��L@�t�=g�����"O�|En�1�d��@��)p��MQ�"O��� 	I=W�1��'��9t"Od(wā� a���-,@�Ô"O��(7ĝ6l��с��-�@�"O<��C�/O�`�H��ܲ/"T��"O)j�	H�骧g��(�+7"O5�&H�ZGTPcu`̹Բ�;�"O��s�OB�G���`o��|�bu�"O�OC�O�����>dJA��"O.����۴c�x ��[�")(t"O�K��l.&yS I�h�hq0�"OJ�0��\VYB1*E�}�v�;�"O�� �F�t�<p�ɕ��|d�2"O0�sެ!:4�6�Y{��z�"O,%�u�\6`��@�� �%���Q"O������yq4R'��X(��'.����(��ʫj<ޭ��A��Pc�p�뉏k�.��FOҢihi^�-f\#>����O�-Y�C׋)I�˔�ŠJ�"���"O���f�e�~(�5H���Z8IA�� �IF�'LB����%�Ł�̋���a��j�@�q/�U���+��`;R��?qB�J~D�)@����gh�^v�I�����x2F8.28)G�']���i����!�#Ptؔ�t���!��ha�/��Em!��#!<�`RM�	'$ȱ+��֓H�!�<���Z�Č<��YB�;%!�D.�>-(���.�P����s�!��]n=q���#&�̰����'
ؑEy���L�Z�ڌ1� �/p1d�����yB'�Fh hQ��2�{D&�~1O��S�g�I�^��yIS-V,2?��4�T$m��C�I�t���X@/J�m<B�JC�NZ��VO��+O�g{, ����
u���H�"O�U 4M�e���� 
�u t"O������}��a�����%�H��ē�hO���S�F�9OIB�N�-o� ݱ�"O��h J �k�I��Ǌv�J���|2�#|OLT9�(�/�tS��V~�t��O
��f�TI�ga��hv����͠*�!��94ĸ�ٶ�ȕ�љR>"6џ����韉"^ldYW�(����m֢x�!�JaC��	�d��f
=�UM"q�!��\(�މ��%�))f�����H�!���>���z�d3*���;Q�Y�-�!�D"���АH?f��E�
��?�!��=�����G���6�Yq��,0�!�O���$a�"T""�zkQ
>�ў���6Q�qI��� |R\k�b�E�PB�I�\�4�c%��M���3둽U�@�=ÓV�L�:s��u�ܥi�@H�B��l��Ms�C\�� ��DN�=|G��!
HN?���S�Ċ3#FcR ��׆/��eDx��';��֗,���9�FD�6��K�'U���ƞN�@�*2dk�)��<����1u�p�&��,�T��dT{�<gV3@�f�`�h��Y�r��q$��<)�Y�&-��W�8�m��"\<��U��~�>&@����0"!
�<�B䉎O�JPq��\'��PB5�ق'�"<q���?m3���a�!���U�bՃqF#}b�'��a1H���
Lk#�pҥ#E�t#|=D}R) �g�? hc�I'�����'��{��Ȣ���C�O���@�/&�f�ж�X&\���ӟ'��RN=$�, ��T*06���sO��yb��{�@�U'R�5�
���c����2�S�OŨܳ�Lp9CcPH4|Q�'��iy"T<&z��%_�{3<d�K��!��'ipk׫��J��0�"AI�mh8e�
�L��\�~h�p2h

C,�l*«D!�AC��Rq���<Y(f�\;}N!��P5����
�;@�ҫI>'!�&{`H�3�^�x��:ut�Ii��H�p\ZfU�kp|�"���V6��f�<�H>E��'A2@3��'_|�x3�J"6�{+O��p�9�OrhKSB�z��s�k�$d`�2G6O�IC8��Ƅ��x�`�S���:�l��J8�xn�\P��(R�֑/@�`.m�B�	�`O"	PgP6�)h$F��8,8㟼�aQ��G����0iT1PG�ūqLd�P���yr��9xpeУ�c���f@��+�Q��?I+�%T� P��jr-:�0�(�-D��C-ʲOUh�"0�
$� Ԭ,�
�z�M�B����D�S�tYs��!�HO�ꓓ(�hL�n���Wѯwv�����ڣ�yb��4R�J�i1��?'�
h�E׍�?B�i>�Exb%�E�<i�b�R;0l6$�)T�y�M+�иh¤��_f�I�����yr�żP+������WjX񢁃��y�g�M����(�ND%!�m��	��'B�{�g"�:�1��[�zu�-� ,H��y�mݽqZFHa�x�l��P����y��$8]�#�	L�zF��(�C��y�)L�E�؝�ġ��r�%�&eÔ�y�C�;��	d$�g��y�BT��O��$��(O�)=mЀ��7�&P�6*��I !�$�#da�$Bd,�s� ��d��6�"�#�O?��"� L�}IC�آc��ոU/�o�<I�jЕs��|��TQ
�ض�q~��'��|�v%H,����eCk�Ě
�'.͓1	�n�0��Rƙ�i+����'�2�Q���G���k�Z ���'20�
iL,(�DI��m�1M�<�pO��#���2☊��*�"�K"�'��㟜�qhP�>��p�$���#D� ��N2W��-�Lh���h J3�IU���{��Y�5-K�`�N$@��S7> ��IB≠0h��cgE�y�Ac��ڝ�@���	h����ѩs���)UCHy�>��T��&S�Q����p�O�JQ3�EL�K�I�V�		YiL�Kܴ+�z��ē�?���.H�R���Q���Dt�=�|O>���]0W` �"%ͬ,�Pza �<��FR�p6�Ȧ���I��_�<�0hR�K�X����#y����V��E?�I<��O�>Qd�
XUAf�	T�x�C?D�0C��_�&U&$h�o�Tՠx:v�>D�H;!(�0R������?�,�;D�\�#�@��}�%2'�W�#�"X��`{�I�������,̞If�p��C䉏6�� �qfA.��]�G5w��C䉚w�^�	E�X1T�q�[�B�	�8���1�([�/�Z���ӿ4���hO�>]�U��^�2�$�ƳT��%,4D��{WL½o8���T���u�)1�O~�De�`j�`�$e���q���[�|AkÈ0D��Ae:?.�xæi��X�zq�0�8�R6�~� p�ф����`2fs}��)e"OZy�P���w�FCuD��KPJ=�F�'��'�jh��(4�a�)��tR��4 ����s��|bG�)�ⴳ�!ך.�����	g�����S�0��ش=s`��,
!򄇜oBa����b�� eF!c�O�6-9O2�ٓ�J6�$d�p%X)�*�[�
O}j���1�l�䓮��E'��y&<m�� ��	�\��(��֫�xR�'^"Y4��?mn¢@iFe����x�&�uoz��ΫE�&ps�����#�S�h}�A�T�Ը�4�L$r4�#�\��y"!�� �|MJa�#4(���b�Q�d���E�S��?�w�w<:��%�j?n�ᦂ�m�<9�	^�<�(�U!?sy���Ci�<��3�&L
��<���1w��M�<a*[$�d�Վ́}5DpaKp�<q��/� �Q���aT9 cDX�<��4�.1�f�������(�X�<i�@O�x���r���I�R�<������<8�,�"#��f�<9�R�{P �{�K��~�u��G�<ѕ*�}.�t2��Z4Hɢ�	~�<Ѡ@�r�,�ؕn�4�<[q��o�<Y��Va�X���R���� ��k�<ɵԝ5�"�Y#?��\���k�<	����-��P	�l��o��)��)�f�<��/�&�i3�G�00:�{B��e�<�#+ݸ��a��9eP�B�z�<����9�F�21�%�G)C|�<�6 �K� ���j�TT���x�<�*S�xr�c��0;���q�<I'��k��4�?^|�E� �s�<���D�<A�ļOT�uq��E�<IR�(���Hr��;��y
�f�<1�A�+����¿G+��i�l�<! 隶F|U�6���6���ǉ�A�<yA�Y�d�(xfJ>J`���$~�<���3!�V��cL�e��� Oy�<9��6v�
�+�Q5}��E� �Tr�<9���(@�X����̯+XA�V��k�<Iq @�=�T�Q��zh*M�S'�f�<��d�,�D<J�kE1=}�l1"B�y�<!⅂%@Ӏ��VkQ0f �c	[�<Ga��-���!�Q�sAL")�k�<c ����%Eԝ_�H���Wj�<!����&�t������f���f�<�G�)���
"��5$�UG�c�<1�Oɘ8]J8S�^1B���۲��v�<��c�Y�z��c�ׁLezd㷤�h�<	*�5�̐
WJ;.��a��@�a�<9�#R�Zj6ay�ɷid�b-�Q�<3�%Dld�֌Ӷx{�=QeM�M�<���M�m�����F6e��Y�RN
F�<Y�A?c,��R42L��.�F�<��cB�J�R���}���0LG{�<�0	�����ڸ0tb����s�<��A�4;�l��䃠BB��V��k�<a&M�>e����E*C�Q��\e�<i�ᛲԤ� �+<d�ڡ@�`�<I�	�b�|̲���?v�VXB�Pb�<���ʘ@F��C*@�&�����O`�<i'�V2�plЄ�V�
�ʙ�l�c�<av��1<��*Ԩ%>�=#�jJ\�<� �t���Yu���{��K(O��� "O����V�S�́�U�N+EQ���2"O���∇�Cv`Y���Q�om����"O�!�ĈOvd�c��-ư�pp"O�x��͔q��p0�F9�j��"O��� �!)�d���?6h i�"OjQ�T�/Ͳ��[	9/F�0�y�D�unU��L~�����HF�y��ޗpP���ڮo��x"�M�y�@GM��y�oB1hN+��ڇ�yRjAd�n�!��]���֥��yBm	�fh� �CYS�F@��y�/^��6	�
�k7*
5+r��L��E�]��]��-KX��!��g����<U��YFFǃ �!�dZ�)S�8��	���:/���!򤅡!:��8� N,��YcL��lt!�d�'e�<�f�AØ�;E�A=t!�$�'&T��gJ��r���Z�IP)S!�DۡH Vt�g��\~��X�-U=?�!�ā�i(�oC�	C�Ԑf*!�!�D���h�-X\LB��hس$��-��<��2�'$3~�k$W-�je)$OSo�<�eɘT�� ��Ύ!���#���h�<��A��D,��ӥ��\����%�\�<aG�F7f�`��P�M��#U�<!��]Y8.t�Cc�%#]~�IT@�S�<�`E�/g�0E�g���9���N�<�RfD�WZ\����Ǜd�N�5ɑM�<���	���2��%�J��oSG�<�F윤;�:ɂ������a �G����<�B �	B�(��x
E��AE�<�`ۑ*r	�!k�CH�����Y{�'	?I�fB>7�X�IaA�1��1D��p k�CC� X@FM�x!�ԭ�<)Q�)�'Wp@+J�u%��[�^6���=q�����(I�Sę� nL&�b�I�D��V��'����#~��6�ē`ը�RS䅹0,1O��:�yBQ?O�����@�D��vL�#�t���"O�r"k�xHk7��NƆ!zt�Imx�P �DFK���
8�j����"D����l��0��%�S
?@�I��E D�X�J@��}#�D�����e" �9�c�O��;E�	�@���5��,>H�؇�j�5{!&�g��\"C&�A�䐗'/ў�?)j��N�h��'�K�t�1�4��%�x�&�8�Qp�hC�Q���zV�]SV�?QE�+�'5e���L��>��M��lV< �ȇ�]�J��'M�o<�U9t��)�':b9Fy��i �
$�V�)��1h�b��!���/e�ҥ(C��{�P��CʳC[!�Ć�xz�&�4M�ؘ�Ţ��=W!�D7<6����)�� �7v!�d*6mN��Ќ�1�:WMj� �'�|�&̅*4����H�x=�
�'/��+�dX�,J��q�PB��3
�'LՀ�eH 2��G�#"�!�'ʛ���.�D�1������ɑ+�y���k(���  �΅z�*��0?�,O�S6��b��z��O�}�"O21�g�ϸ2��Q� �@�9q�%3�"O�Q�ՈX�^�1�i�?�F�j��'�ў���mZ�q�b��aCă׽p�8B�	�e��Y���ܮVU�]�0F�?i,xB�)� �|���)�x|��lѿH��1Z"O�B�Ⴟ	.\%���T۠�`�x��']��
bU�V� ��*u�@��4U����t?I�G�5����C�J�pbY~�<Y�NQ�5*�eW�DN��gA�s�<��_�(s��q :Q_j�iSS[�<A��Z\�H��I,xZ��u�
T�<�Ҍ	�"��@���
�L|	�&�YJ�<Qp��\w������T&Rܱ��j�<yAeYbܔ9@��l����Ԥ�����X���S��nнh�hYd�,��ȓr���p ƺT����P��E}��ȓ֪�8uI��iخP�aV��H-���'"�A��V�V�DQ�7�/hY�`����y҄Y+GoV�$�LH����"��y���%y(���d�O��3�n^��yR!	4j��r�O�Sd�ua��G���?1�'����Ao[�-���dI:8��)����xҊ�%#�(��P	
pYz���F��=��y�BI$4�(���Ek��y�F���y�.��1bVuip��e"	P��� �y�@`�Ne�ɐ�\A���!�̴�y���MP�W��&� <(���y�#�,s�a�$��4h�����I�y���
����pˆ?Y��hh�`�>�?��'q�iKr۟Km\}Y��T>|��	�'��]bm)���r1�H�~��'9� ÊU�4hҀ�_�9���'�f(��N܈a��=y���/��q�{B�'A��R��ݧ-�֜)��\Ej᪋� O71�L���ޱJ	p9�U%ʆ��z������B��)�h�=t|e遢�L����f<�EKSΠ�G�oq�19Wĉc��8�<���	^!<���aG0_V���^쓡y��O������&K)�����7�^C�'8�9���ނ�q�n�	s�E*�'�tJ�E��/$*<��㖉��PZ��DW�O���yVʗ;/�H}��%���(}#�'r�<��JP�B8�չ�̀% rش�hO?7�S�V+§U�_C���Ѵ0G!�D�����Q2%-p��G�Yk)�I�<Q�������'(z�T���^�f1zC�D��y"!U>�V��ƃ�~��mpcΝ��y2����l�v��u����'�R!�y�Q�r�v;2��E�mb�N�8�y��ôt>���@��>����C��y"\E^�adO��0؅+6f���yO�
{����Ov;R�	&�������>b) X������5>xLix��|��࡯OZ��%EN	L�~�c�l�)��r�"ON�XP�ڛ>��bv�5z��O��S���=���s�	�(O���*Ь��sC!��%�2����I	6.�Ș��B� �џ���NU�OGr���5h
�-@DF�]^\�`�'��b1A�\���S�R���,O��.�)ʧ,�p�5�Ej�����
�B����ȓ/�"�y)W�u$:Y�գ7*��ȓ|�(�z��*J�tZg%؊���m��<!�}B��&fߚ�92U�r��a`'������Oj� <4-JRϑ�0��L��]'ఇ�/�"1hР��F�޸���Yt���ȓD�vĐ ��J���
�R�u��o����Y�_�G�£�d\�@��5�!�I�~����i
6mF,��Ĭ�F6��~��(�� -;��5��@B�X6&��*�x��'iH}2�S�P/bMjQ���bx�O���<�4�])^���0����x�	���~�<9�ݱ<���p�Bnk��y�'�NaD��	��Q������X�#��]02l��y2�
$��i�h� �H1���y"�)����ybOB�\붊��'	����ۃ/⍲���5�O:��p�Lh" �8<جY���L4C�����)�O�������2?����/7yHZD�O����'�$*�>���c7��bRl�f\J�VIC��y��ϞU���更Y�J _���$3�O�Y��̎�r�d�â ۯS�V�	3"O( �F�1T����AR�@��"O�<��)�*�2/܁1����r�>э�4�,O���@��\�zțv��46�����"O��2C�ڿ5]ԣ�$�^�[1��b�����TS�@�%(U4i&��2G� ;ߡ�jӔؑ�h��l
ԃ���,e��R�E{��C/a����,�T�`EL�d!�d߲*v���N�t,SG)X�5T!�ڮE������F�.�	�'��$��2;O�s�Zo�$�����䀨�"OD��#
ʅ)"�c�֋Aľx�"O�s�C��Y4n����<����P"O�x�$Cֺ>���I�fJ: mH[�"O(����C���ű'j")S`"Op(��Kv����D0Ea�`Z"O(�����W���Ѡ�	�m1�"O�9��Òi.�)+��O�:���%"O^`�@�U�!�8�ٓ+! �@<��"Ot��b!.�`Cp`Qr~N|��"O��&m p�������g�RAxc"Oޕ�aHԫ	�D �E��,���;4"O��⇆�"�	�c�n3M��"O:<�i���iQ��9(���"O����OL76�ʥ�Q;iJe�"O��Q���L�ĭ��*�8t��9�	�'��$�n�:�@1�d�g�\�'�(=��� (��V;e��@�
�' BEh�m��|d� �]J^ :	�'0y�T$�~�a��/O<� ��'۰�2�/VcLh��+�
8XN(�'�R��P#��ߘ��Ay�����'@hu�rfE?]`�Yjd>k�J���'b2��p��I�l���ةe�J P�'�|��eJ;>��S
ϑ��x�'ʪD�ag;	�$p�+��@�4�'���ѭ�_I��dhAvt��C
�'��pxF%:N|tiNf' �
�'.��[�G ��1�V�\���C�'���A��Ju
faH�#���' �-QT�0N4d�EM�3��I�'�x�$ƅ1%w��fM1ެ�(�'��=�W(Ԩa8f��T�ɗru��'ż�B�h^^�����Za�Lh��4	ȑg��=�(���1g�U)'f��[�Y�J�R��B�I��0e���\�؉�(S�+ fB�	�?Ȑ���'��@�	���P��zB䉵1m��B/K�>b��q. 9wB䉂q����G�-	�y��b�jmB�I�p$|��̗ 8|�+@cȭv��C�	&U���i�`�1%'nԳ穆�k~�C�I7w����v�����"����C�)� �lID��t����
),Q+�"O�̪' ۫wVb��ucS�_d���,z��jGeƎ\64q����2�؛d�L���*�dv�9P���y�L�tk�ub��V¼mj�蓣�?I�&�Q$��q��w�:=�%���v��=a�$��	0��,��I�Eq4��ҔNas'"��L�2L2�D� G2����H7z!&ٔ�'K:T�L_e����L�G���{2GY�	�@{���g��hӥU%gs�O`h\�Ef�1(��9Hci�2� �R�'�J@UNúAP��釣ٝ�X9��*D5S�8�+d�
|=���ǎU���ܹb�'�҄��!�x�������}	L8��'Қ-8FƛBf�����S4�Tjӌ�ca��D�F,	%�4ɞ% �	�"�(r�m�;���C��S/v���[�v�AgLG�r�P�#�j�j% �Y���"�OC>3o8$���K���>ICDڀ-Vd+���%;�BE9P��z�I�Ju*��`��va�h[0��oB(�$���)����(�@8�|h���A�-b!���\��b)�{5�� �
΂#j\a��픘,� ��ף�B��,�F�W�SA��<�6�<Yb	ʔJ���q)C-��i$��JR�\��TO≓$��	�O1D 2\��I�>x�K�Ț��5�`B�;u����M3g��1��s�'y2����ۺC�B�sB�� f�4��'���G"ܒhi 5'��GB\�ieÔ��9r�c��W�t�G�E�k�uSR�P#5�^H�G }�a}2h��eNn�pl@�0�]c&k )��I���hf�Y/J� z�ᘐ]1H-C M@�fԞ��T j��[#���zRVk�(��N��]�wn(�O*�/������:�����ԍ�2��ªD�wczY�-�y|V�h�h�(�L$b�V9���XP�x��L��M�b��(F�R�r$��09IL�'P�'\�HC�^�R��d2�?Q�f�ҏn4l�0�PC��U��Z3dc,��v���xA@����F&Rm3|!EzҌ�6o~�R�헨D&8T����y�F/ �`�2��8��ɛ^�`�Uʑ�
��LB�ϰ4.ΰ�W!"W���nϙt�k�⎩y�"%M�а>с�Iꢽ�ե�IAx)ѡ��3�򄖖 a6-��G>$�lT	�B9nc~IQ &ӒZBj��<�洀wN�?S#H-*�^��H���'c��	�焾v[R�hV�H�%p�8`��ǆ�~\Z��a�� 0�G P$l@�%TRF�Hv�?��P�Z�H���n�5@j��U"��
񈑢�{�>#>Y���,R�Dx���ԡ��	͐X�8rb��P���ap%�	 ���Z��+��X��� Z�`p	�.v�2J�B?�QuBh��c��~����ю@�H	����Ć�t���O���ƞ�r��(��*��<-"<Y�+Јf|�', x �H��Y��@�g
�>IEf&S8 řTe8���Q�i��
�,v�%���M�V��Đ�jƢ=����r��:8�t�������ETe�e����F3��ȓH���X���aEP0��9S��ܹTMq�I�D�w���(̜I��O��+�HLܼ� �2�j���@թ�`��PC�']�Ⱥeg�C̓w^tD��`ꉄ�B�`dDA�CC����5��h��
ECd"D+�t��丧��$eP���FO�R����',"9�b�%1{qO�M��ǒ>jDZ��ݬ'>�� �$L���,��&�7(�x��T�^�@H�x9��/�Ol@�'A��YP��fխq'��8&�>�J�+Y�HT!�k�*�"V���޸�e.D����Ӛ~�(�񴩜
s`PH�b��B�=�O��I7��<>&�2� �6�Ĵ��e�q5��&#B�p��Z#�*_. g��l6*�"��D�La?1R�²�����"ʠ��=�U"^{�'�"0�(�/��|�㍟o;�\#v!��' �����5}1��ᆃ�4`�RR�ϱj<Q��	����bʃ�P��ts$�׬6����Q ����Z�S��S���P�n��ІՁ	ִP0���e'h��l�p"�[���X	�	�J�2n��E�ЂZ�d!$�z+G#��!�80BZ!Sb�Op0b �`>���C�s�X��*��<�~��c<�O@�(�G]�l���1g�R	�Mۆ�jUE�'pL
cFn�@߶˓%�£|�	�	�Љ�Ŋ�$s"𰖇�3m?l�>��)_�v�a"�&|2�!I6r	�36/�=rC��zޤȐ���TG�U���F�y��d�b-§��S�O70u�c�	<|A�	��B�TR�'��LZ�H�H���`�G�Qfh�K>�@�Ǘ	Sd���ZxT��J�[��p[4M�$�!���A�q��dű[����� � �!�:^ (��&�
Qn��W,HX�!�dZ>4�@`����#�L;��?�!�DN��՛'/ȫ`�(�Pu�'R�!�D�'N�� �@<h� �6Km�˓3^�8р�A�(���O��ɦ�ј)�8Q����IȽ��'̭3����m~F,��.Q� �n�����.��t�ń:���)� d���š5������&{��X��	�lmx�"��U@�B� �}��JUHPQFo��M��s��:�ȓk[�)��O�5��@1�­T�m1g��FB�"q���Y��ȟ��嘑
ep(%ʏ�ˤX�VcW��y$E8Bx���J	e��"�h�/GX,�	�{��� ��*W�N�b�����ъ�A����^V��A�,�O��3Re9T��
�k�j��W�ܾ]�ʐs`/�	��)�f�6�O�)ذ�X�z+���.4{�82�I;� \8�lH�f1�% ��ڟ�CA�t>Q��?�.�h�&�=:�1�O �0�υ7A���`�YS�kW�i������Txd��kˁu�6�i+��� 4�s���C.
8���"n�5��,D���1M��<��"cf��{uI�K�d�+�Cɩ2fd ��Ǒ7y��L@�	C�Y��ɍ5�b���g&T�t02��6aP��$4dZ�xé� ,_��0$��n�f�!���#�%ڏ�M�M�0Nl@`0� Oc�d�h󼱸FD��M2<uA��Ɂa���Q-7Ռ�	',Ϥ(h�H ?�T�1�O/>1�`;4$�Zt�x)�
O����ԎS����,�O($�4�ɠ2v䤢q"˗�q�J �������.Z��s �^�y��Z�l3�ł�	> ����w�1�y#�-���SR�����N��6nA�@��p�b��P$.B�I�C���dδ���IG*��h9�3l�W"0��D��f����RE�F&�5*���$jSa~B"R�*�)U�̓_����H) �f�׭�,* �8�� p�+WN5e���s�m� I0�E}g�0p�AC6�)�m%�� #'�0\��|�� b!�$@,^�p��bH��7�lY�6� h��IBЀ�iw�铄b�i��CA>mt�ъu)�%�FC� ���@�&)o���"��CfC��+T5�:�.� -��5�`f�7i����1�F��O(����D?�"��$����`l�<*��^g�<�$�[5<a8%�		@+!��u}b�+�&@l�6vH�d�B�)�$b����k��Տ�\,3���>�>A,�5x�B��KȺ� �X�D���r�K� �V��L[� [��'@n#}�'K�$jݸp�]�-�QSJ)B����+ �a2��)ՌN-2�k7�K=d��������)Ňp�\�b"l��P��-�N��Q`��5
���V�|Ӳ�UC�������:�
c��m�����^��)��l�-��TC��VL��B�	A�>����/Yl������7z���Q0p�J&=^[��;���Nn�I�5ex��"��ĈI���,:f�Ɋ掘+ ��}�!���s����@� 1�1�M�)���Xg�����ўA�ވ�����@/"8��%�S�c.�TSRaK�0�!��@.!0����c�!z�iCAi��]5ZqJ��4w ���
�2�ɠ 5�Q*cF�7��� �x��=�'c7�)(����k��D�1D���?��O��	�J��$+� ����Um�<���"E>�"�U<V��"GAǟ,B�@C�ahZ�	γ#w`�M��<	�F|�':���q�ͭἜ1k��܇�ɗr&j���Q�zu��B�� J�
m����r= �� ,A`?	�@/x3 ��|�<�g#G��	j�_�Ҩ�8 Pp�+9B$P����A�?ѓ�ɽu��%3�@N6$<Z���A�p�����	��tE�i�G*:YJ��&T��$r�$��hr~��K��a\w�2d��Õ)/Lz�W��ؿFƊ��S��Ϫ��$?��
�'6^<1��S%~񙆆N+3`��ڴ&��Xb#��,>���1�wyB)M�	��XSK~zuL�/���J@����Y� �N؞�`�8-o 8���'�| 
�g�����霕4k�y�_���"ɤv]Ƅ��%FxR�ŸP~��3����ذ���"��'n� �H·�J�%?5�h�6�T�0"��5N󼱺�w�Ă0`M� ��U��Ɏ��<�����cxtд'$q���( �*�]�O���A�bY ��������Ӽ� +m�nċƅV�_���OHN�<�u�	�h`Ȓ�I&&ŖKt 	ɟ��J��+�\:"�0F���e�iR�����̘OT��B!��U�,�
ˠd>�}��xZ-�λ����hP�'J�T�[�z�$��Bi�
Ah�Ĉ58K�M��(�)$��g�'�B��ebX![�"� &�ʅkq���
�9��`yF��. ��h3�e[��,=��B1<�"�82,�4FP��q�2�O^�q� �?SZ	<P'ļ+��ɛF	D�+���b��cբ����� Ԓ��ɠ���ۗd0��'�	�|�܂���,O��@5�� p^��Ə6��c��2�E�1��q����4� tC��y
ErR��v�bia L�C3�%�"~ΓM���#��R,�qAF� ovJe��n�N.�'�戚��H�B&7|#<�@a�fdG��O`x�W"=��(�D����Q��-�B��N���R�A}+l�*��9�$[$�ai=Z�86m��~'r�IwN�I�j�����n�az�%n�HX{��w?�ug
���j7�C�/�b�)�n�=�p��kO�'#}�D�۾����P�T���y3L�iܓp��1vO��ȟ.���F�֝�s�F�(�6L�H�;T�@�0��]Y�d0�g?I�O���H�;B
ƝR���Y4�ǜe�@�0�{�#.�g}��-ff|�P�+�&7�0���٩�?q6&��EJ�L#lO���'H6]�d���'ҔU|� :r�'~*UeǏ�'���l�U7&��%�.#�2��
�
�dOD$BE@����<��H���3
�[,횂�	�4�4���A��ݛ����@�
�������)��}���̹l�����ș�|�!���'1�\��Nk�X�SPb��p>�ZB���=�v�(�au?|\�O�NU��@�F�#8�X�a�����Frf����'�p}��KA��`4q�I#]L�ڟ'�Ԉ�G�S�L8�Ox-��Ü�'������P����k���\�%@Z>/���q&鐐u�!�$�hr�aU�ؗ�b\I$IE����1-< ��RS>
��d�;���O��,ӨQI�f]�[.X�P)IMP����%%"�Y���8P� ��gQ��1qg��'>��� 	:�AIVE*}"�sӮ�   �i�\���׎5ap����I5�4 ��Y��q�"Dh�"(�r��Ҧ Vj���vP������0)�zc�'�T9نф)�@K�.�wΘr�'JU�"���@�j�O�O8f�i�*L>PI�- �O��kt�0`(�*(b�h��JBh<�A�N�4z� �+U1St���s�S~��a��y!�ܫ$>�iR�5 ����͂7Rpqac��[,X�hӉ(�p?)%��	�@�����$���E!�V!� )ь�K(�T��h�?U
�O?7�R:�
`HF�M	�E$A�h,^-�����Y`�����EF!�U#J`v�9�O���$�,W��H)��<9GKߋz�>�c�-^)'�ձ���Bx�С�L�q���EbYZ�6�����>f�Tu�d @�<�b⟛)�>�R#�#�P�1�<�ZYH�c%7ʧ�P��s&�?<+r� ��^����"4v��
$MY6�xs�x�u���\��H7c�J����=n
Z	�ȓ'F������Q�a�`��[ʄ,�ȓb޵�7N[�8�\������V,E��)Ä�-J����*'�\5�ȓu&�H��P�,�1��РA�I�ȓVu��9���/.��h�b��2xr��ȓ-�����M]�@�wFJ>/P]�ȓ(�J�toJ�cy0� �:Ԗ��ȓ6l�ԣN��`r�F��ॄ�Q�F%3�cA9h�l��F_�Q&����p�U:���N3��y��ƅ}�P��'��y�S��M�H��aKV{���, e�%�S��My��V�m"T�ȓ
��$��^�����5@ۮiֹ�ȓ}�t�2�L�]�]sUB$=�e��RR��B%�*��P)p��`�<��,PB�U�A<XHr"c]�*�4��v.-��Àu�$���<Co� ��l���#�P�y�����'D�|`�e�":�8�8��HTȨ��G%D� 
V�qrU�l�2:���C/"D�����$��b�ɼf|,�O%D����X�?2�	PUh�*A�T��K'D�8�H�3R�����J�.�+U�$D���� �+?)H�wIF�|�ѳ� D�<� +�R �k���0�rm �4D�4rG$�s+�	5�XT�����4D�� �IPZ-K[�)0�%O�o���"O�9�wV?k�j��c(8�5"OR�{���R`h0C-L�<�e"O �t(�9�й��OAZ�Q�t"O���B��Y�h�ĢG-BF���"O<)��i!\:p�a�����C�k�<9S
��y�2��0��}x��]|�<�`/��h�S��a�p�cR-�<D����!���'�t�;СX^�<��f�C�QĪA��p����X�<Y��UB p��H�n���qd�X�<KBf�
vbA5#! ��R�<EIܣ0�9j��0A�%,�M�<y4�5B�.��/��](X�9�D�N�<��� �,�Pl�b+�`��@�H�<	��I�.�\8���)a��+�G�<yr 	�N�!1�,O�[���u�<�R�I�?�~:��R,n�����s�<�ŏ��g�*��f�Ӄ�xi��aS�<ف�0�4�S�O�0�����t�<���
`���)ܯ���3H\}�'��\SOHO�q���ЁOD�N X ��-L�|(E"O@��C�ե|n��i�1�Z�i&�O,�c ���M~4��O��}��Ğ�x� �r
!b7���F�VG�<��"C�Ⱃ"� j���
�Jۿ��d�j��R��o��3�,^ܡ6�����T)*\����	,��I�P���lL0ə�戠ak��2��ቶ�@D��$+�-;~���O��xd�\	�G=� �jMӥ��,\�=!K~*�o�#Ni�y�S�"��8qs�N�<i���&�z��"�Ȧא��A��<y�Lǽ-]�P���	���6� �� �**�NU�cF�`j�C�I�Lx4�Sy��kp��(͕'��d/��#xd�̟���k�*h~ �Ŏ 콐��?�OZ�zT�:Z��d�p�<*�%4�b!cn� ��D�0�-�O���cd΀:���Q�		[�n�����_~��! ��5=�8%?�
3�ů\Nu�.I
P���':D� �3��vniKG�^(D]ːC��<�3�)Z?��R1�>E�4b1~l�1���ۣj�p�g� �y2�J/h� �"G$��%X@��&�ē!I��V���p<AgI�7h�0ҕ���Uڅz�C䉊x� �@�%>N���wf�՞C�I�~@�t�i̳ -�CbHR9_�J�?q���0� b?qh"�4dD�0G��.)�z-�B�0D��z�,@�|���G3u@!i2)�>��'H=���K>E�T�ǜ~G21����J�zՂS2�y�A�'��e����<vC�p	�d\2���'x���b���eax�ˆT�����G/cl� ��](�p?aW�H,\D�H�L%a=�a���V�i�٣�GʠC���P���`�O+^$�v��)`"�>�� �鉲2�5D��%��"���\��n��5^C�I�G�Z��P����c�X<q,�I�'t��tLO���S�O�H�ՉA�zG�e�Ŧ�
��	�'pt���}׎D" ��w��i�H��4 U�=���r����J�@P���hI�`�4ȒCM�G��X3�!�.�f��R�^�,��0��o��r��'`��.�!�ش&9Z�HC�*M��9C��3C�Q�H{�c7������Tk�(Pm���`2*�.�!�DPТH�gLZ
@ ���F ���<b�X*�'u�)ҧ�:�	�₥DA��$��]�Y�ȓC��3���%�\$�5�	p�&� ���	ay�F���j]��d�r��(��A���PyBDΧ<'�1��H>N�B���
]�<��!������f��y�ΕY�<7.["����>N�b%��_�<� �|+�ȕY�r���@��\~��r"O0$�7@l�b��ќ9o��&*�<�5˅�Gq䴑�h�����U��
� :sN�kO���}���!Hu���Qa�4B��o��n�fEyq!�X؟���o]4).����A9:���H��3ғ�������O�M�@.�����I���1KN�~���χiFB�ɭ=XP�!�H<�3ԇO4(6M+_�6��Iq����B�E��MfL4s-RD9C-K"��a)��Z�<�R���D*z(Y�#Mr�zɩ�Ʌ,�����F3ʔAWN�\�D0��HOڑ��^55�
5�B��'*�h�.L8l%�A���YÂi�a�� Rw��s��W��4��'c�����,�p��Qȝ%h��S����32zMSk˔g4D����O�!C`V�	�<Y�
Őy��x{��,+>�y��'X�D��L��B���X��T-*cP��ٴIҘ��hٷ��.eX�n�ܦ=��"�0��5F��
04��I��؊��|�����yb��=](��D� �~h8�#��c<=���[BL�pi�� >������*I9>�'c�J�!\��N�P@�2s|�mI	�s~�yaa�]�L�XrA�L����qv��D�$��6-��bS
Xѱ �p<��(qS�'�TRb�+V"�H�'}�.ʠ��l���'�@8BgLU�p��&#��at0����X���!ѩGz(<�R��,��9�$��FU u9P��D�'R��T�;B�n��}z��'���n�	s�ة��!�E�<A �T�I�́
ԥI-w?4�����<�t*��FQ��J�#}��I�~
��� ���U�(�*��]�q�!��v�`���2j��<����>x�	�g�<y)T��xra�Z���k�Iŭ=l��k�]��0?����̚&e�\$sb�.��\�'��k��B�I�{B��EEK!��� @L�[T�>����RQ,�������c�U�"��CX�� 2 �y"	
/):�tR� X�G��9��hS���"��4Ҍ{��	C�@�Z5��obpc�8d!�]B9$1�שY2c��p�Y��!�D�?(.0G��vn�ѧfֶ>�a|bK>4�����Vr�{�c�(���M0�e�ȓ!�܈�R"K�1_��`���X%�?�1�#FF���IT��pjs$��a�(=ZݐS+�B�	�M����B߻{I����aߘ}���tm݌M-�O%E��Oh��gţmJ
Y�E�悉��"O��h��#��Da��p!����i����$٠9� ��It�{5%[�n�tA���>9�F��Dʶߦ�"�ܞ{x��P5�@B���l�H�����<<���ȓeuXM�B��v۔yf��s�`L�O�!�Vl̄&�v��t��*KB�>��_8c8��C*�%`:d�	0D�@ٖ��F�IB���{o��y��ݕh��;tI�t��Z4|�c>c�xa�ֳ_:�)�3s�`z�N;�pAs�ץUX���"{>��!-����u
%Ő�}fJ	�g�m��캇ɒ�B*X�ѩL+-� q����z�(:��4���AˌHoTq�ti�-_�t�����2���Ow�}ۂ(A�PC!򤂆Z*�	���8
X�i�gR�t��B�!HN>�� ��pv(�`7	��[*�91����B�7�8��O6�"�'��R��E 8�I{M�q���`�d�sw
�@_J���dQ���:hZ�4����y�F���D��g*�Jț�#E��'�n��}9`��bc/�
yI �"M!V�`qB*�Ț��0�S-�����Z����Z
k|��&-�]����ٞt��'0�֝-x��t�3�E�6�^p��5��=Q�`�4�O�+9D�	w����y2�muH��	�"�:�����MS�MZVArd&>Ē��'.taQ�	��'���/�1/'�u���=k����7,�[�`'LaR-IR�>���	٢$-Xр�B�o��ɧf���0�C��oD��g�'�֕0�m�W�Bt��,0%��x�}�̈%>��7B�v�	">�����p!XY��pm£@ޫX���0'
O�=I���~��eɤ��A���8BZGLP�gk9}bl�4$���poW0/���(���ݾ"wF\��Z�#�1�Bf�=JB�I6fs�u�GgI�?9���u&�L�J�D�6|z�,�#�=\cj���)Ķ�M��/� {v��|R��1jj��r!��4X�<c��|�Ē���#��� ��H��F3e�H�!UNV�0��x�� �if<[f�W�p�Y�*OJ�3�>�j#���|u�c����Ň�I�e����'a_VU�F�2x�ni�$�G�A�ڍ9�eԷkt1���'F��9�/�>o%Er�ɉ&E� ��D��A���f�%R��XD�@�g�B%z(㵢�.s�u[�Nf�'��l�GK�G�O�q�&C׻��Mj0J�\9�xC�y���Y5�H��w�Ol�
��� F��[$JY�].ݻ��Y R^�!r�|��9O�ԣנ�_�|�/84��R) ����w@D����%P�#|�'G`�3�Ds �hwBܠ�6���?aD�	w@Jt%�����h�k��$�����	�PH�Ի����� x��!�v[<q�JH�y��7���\��	֨^��|0j\�)�az+.b~01en�T?�5lP�!J@HE�C2+^,US�p��Ke�a��Y"+F�"}��C��ws�$�P�˚H��x��Xܓ$�F�*%��<�ȟ8@B��GVuy�Ѻ,��c�$ !(�!��W��)�g?a���|�l��O]�Z��=jfHW�Nuɏ{2�&�g}�#I���c�oU��X��.�?�P�@9 �.�iE�1lOr�)& ��0yDȈUgʼ;���B�'w���#*K%�z�mZ&!�l� �{h�+f�"c�O��wNL���<QP$�I���e����`��$�d��Lؐ���@ȕ5�������� 5h-8�h�(8K�AT�BB�dQ�f0$���� ]�I��vL�%w��k�jU�i����x��tXp"��6��i��f-Y:*����V��_޾�`��6?���&����$D:W�.d��\�w��4��L����^��%8W�K����,�t�Ю�!���v��Q{�b�r��1�)S�5�<<��O0D��w��=&���iO�G���6�0?-S�x�nPw�!2��J�gD��IPz��X�HH>8�U��*D<5h�z��<��F� [�N͡!�ŞED���@���8���T����
R҈�O �}n�8}%L��Ēj�+��,�$���$�?���)B��O�U���	���¥C�0��1��O|YXGg-P&��ϓ�́1���pt�iұK˜v�l�g�Y�g�$��ҧ�',v�]@i1Gv���օc��U��(��wzQ�%/4�����Α4l���N>JN�3 �4?Ѡ�M��4�G`�}�&�Yr����IP
� �c#�9�z�C�Gi�������826�3�O���Hh��C�$�@Q�$)C8�hYK�!��5<:ҧ���F�P���"�	`&����h���O�H�SE���OJ��b��Th��`fA�)D��K�O^�jc�ǲxhE)
�pP@�5��
u�.�U�e�@��	�d�T)WAE�r\R!�!b��ax-FJɖ<:����zA�!XR�H�M��J�-��kf&�E|Ro�4INE���S8z���8Cg���fb��yR+�1�n��ġ.z�{�.��y� N�F{L|��)C��e�GQ�y�!�0p���Q�#��	�ڔ����y��b��Tlх5C�|���Ų�y���.AgvD�%D�~���z�H�4�y��G�h���&ݹv ~�"�K��y���R�ޘK���&h"D�Ƀ 
��y"
�4(؉����j*��ǆ���y�h�r<$�F���e�Ryj�n[��y"o�#l�`���ڳntT� �H��yB`�'I�����kL�[b��0[0�ybm�2yG��З�9���������y/WUH�Rǩ6k̶�Eg�y��J�Vu��Z�h��`|��I�y�		l�@�S'H�P�8��n
-�yb�^�r��bF�\ך8�����yRD�6&`�<���'?�ŀa��y"��
�"M�PC�H����'��y�=hUk��'7V<�bF�y�C�u�g�[*r��R� ��y�o��@4Ʌj�G��p�a���y� F*V� 9�����>vD鉆�yB�	
5-~�{�
��^�d9x�@��y�oKI��Af�Y�e��8���ˤ�p=掘.9�P��I�<Z[2� ��y@gT�D��)z�
�F^Xp�K�uD�A���"w�`�i��E矢|�;�^�1�m�H9k�ɒ�:,t��2Ʌ�ٔu���3�.-��B�+)�a�$���HA�����F�8��!��;#ؼ��K,j��%cT���,D��'P6�����?,�!���W?z�	u�H�9)��+�'Q6���.�`��
G�Et�� ǅD� �ɚ��@�H�rdQT��p]J�r��,)o�	�O�������#���K���R��͟�0X�0@� q��5K���M��M���~)r��}H�����xQ�Pʷ<9s�>�~*ϟ0��`;wǞ��v���V�[V��3�L�7�~bNUX���*E1F:
g�.�?L��(�S�O]�H3���V�R�B%�:Y��
�'����Hm$�z�'����IǓ���	��#�Y	։�9M<��0d�X�~ARq" ��՟���#�H��S�?�Z�'�]h,���,ǅK
t0���Op)�O��p&�[>�pT-ߝ^\�h�E
}S�	�"*�I��Q
����	X>a��;�J-Qfʈ�W��)��b�>�EJ�>��>���4:��Mc�h
��䰀�U�[#Z������ǅ�?駨�@l� gQ/ ��5C���t�0#�6��ė�]�T�������O-0�`���q���'�Y$AH���'��X)�_�|IXd��6&�R�I�'xE+��AK�,��!,f@�		�'�f���MQ��h��t��9#�n�A�'��I%��S�O��)Ī����9��N�6��A�A�R��0|�dV<:*h���Q�v���q�
|�'5�"=�;+�< �o_��:�OE�M�4�'�%1�D�O�0�7�ϥ1ՉO
���~�§F�`���ӊ�P�Z� ��~2�<�A���l }���Ѐ�A5����	��M�HA3S�7�yb�>N�n�*@�Җt���B �yB��$/3��$IM
q*���6�ǯ�y�g�)B�p���U�l����yr��!z��s)�,K,:1C��yr�G�#:��*#B�
m��ʄ��y"�̄1�T�č� g���{�oX��y��� $"X�`��Y mc�@*Ub�3�y2"+7>9��H�v�xa���y��&T2�5јgp� �i��y�
�6e����m��`b���-��y2+�0BBHO�����B��yҬ�02�6#_N~
(S%ʋ��y��(&K*tk��%YhА)�Û�yB�Y�d����o�	X�d�	���y���f-�ux@/Œ@�ځ�Q
܇�y��_�I��񺠈��8/@���nL��y�LZS�ih�Hϼ0�T�#��=�yRcڵ��Hժ��%un1
�D��y�c.A�T� HU���h!�/ֲ�y�*�d���a�r�Ɨ��y���Q�d�S��S�*���⍟�y�,�5<�X��#MH�YgMC��y¬ܽ��X�p��>P��o� �yb��RL QR0I_�B1�*�/E�y" ��j.�}�T���P m�fʓ<�y��A�����Ѭ�SN�%��yB��-3�5�D���Mvt�����y�CW�Y\Z�CӺI
���	G��y��E�P:�n��Ur��7�y��20l��1���d�@�) J��yR�2%�^�x��;Zy�� >����ȓ3��%��eS�8k@HC�����ȓ4���"��)0��k�o���+,�O��I�8%�dϫd�	�p���L�FC�ID���֩�Ҙ�x��C��4���z���G-bm{�đ Ov(C䉜 <�x52 Z�)�$SR�C�ɗ���c�W{��)�b+0x,e��S�? �A��p��� fL�\5d��"O���U,���� /`QR�"O�i@d�3ZFXX�AC��\'J@��"O2�q��92�c6�ι'&Z�;�"O�9
pB�B7$�3�,+U"OX@)'�U?jj�2 *A#%�h�"O��@&g�p�j��S�j���"OY��P�'9P,��HW!P��"O�8c��7T*�
�FM�2��P"O8!S�E�v;�@Yd��?E�ԣ3"O�캅oGJ�NQ��$!��ى6"Oxs���b�`EkN(հĈ'"O0��a	M0Kq
AWMŧs�YC�"O��f��7A�9 A*F�W8t��"O.Y�w��(x� L���O4wSB��V"O���U#܇I���rb.��N]&8�"O�"'�\RI!/�9WQ�i�"O�šsj�v<N`�qKG5�(Q�"O���AJU�QW�qqJ^�u�)�"O�#f ;%sP�p�hN=|it���"O(\���������i�<d��0G"O���S(�w�����Yc���P"O͚�)��v"� ��I_���̐"O�ѻ�F�_���u	�J���"Oع�̌�}T`����ۻ�РY�"O�3`F��0�ف]:�r�"O�
Q)�09�(�b�K�'��IV"Or���'D�L�b�r��L�x�'"OxX�pj�V�������0�"O.�V������F�F����"Oּ#�.PB�� ���Rc�kS"O �˄c�*-"P�Dϕ�R�����"O
�(��U�E�`����^M�+u"O��ꣅ˺|�|�j�ǐ�.���s"O`���M�d���R­�4G���3"O�Y��54�̰�c�6Q���S"O8ݲ4�F���c�
{��E��"Ot]#���-�E��A�:q���"OĀ���#0?Z�cvF�l4�X2"O��0ޮZ1�DZ�g�<0E���"O����v��ypQ=}�����"O��Q����Mf�p��>Tа0"O����X�Y�i����>K^q�"Ol��G!�*y{��`� IU�=kU"O� 
U�.Z	�P�W�ݾV6~�AR"Odr Â�l���
D瞜{%�5)�"ON��W�2,�(	���I!Q{�"O��D�˸v��S&�Xw"O��Q��x�f�(�`��.�0�b"O�!���B���&���W��("O֩�Da�%c.��	��$�J�"O�	�b�<@7���gݷr��G"O(��@nH�	>�p�&qhHA�"O��B��0�F8	c�Ws� @J"O�dɃ(B� ��Ѵ�����Uӆ"O�}�s]�D<x���F�6z��H�"O��5(�)�I�G�ltbع�"O�X�S�K�M�d�X�L�S9�h��"O���U�1&� ��c%���"O�$;�ڢg�,LbD�*���s�"Om�p��	.mtE)��L�d�����"O~�ul�>&RP�@5��*J4�Ig"O|$34�B8�4�c5�I5�pH4"O�(He �D�bd���gH��"O� ���`d�*L2���2�ΆY`�XR�"O88#u	�~��c`�2R|%r�"O�Mx�e���Q���4"O�DoB0�@@t�۷sؖ`K"O�\Q�甦2HBԫ��͈C�<��"O��7��|z2�hX�Tl�i�"�y��TN��Jǈ �c�dq��T�y�C�_� D�B�oЪ]���Χ�y��H?�ʸ�q��3i�thP!�y�/ aZ\qpQ�1�*��B��yr�h'�p�(��A�`"��y�)Y� <T�Sf�7���81A�?�yB�Ӽp�0��a�߁2� @�A���y�?u���qH�0�d@�-ͩ�yjA�7 �P�(3����	�y"lD( ���c���NZ��hd`��yRLV~�H�����r����y���ڠ�7甕~�
�)�Œ�y��$�tC鏰u��0�Eԓ�y��@$a�ݙ�eҼn��9�f��yR���ő'.��\k�͙��	�y��Z�W��ca+Q�\��Xp �N��y�!�6Mdv����X>VD��뇭�yҏǶnʺ�S�f�I�چ�=�yBF�]�>5�pÁ����&����y�H	BɄeCL��+Vpp�E���yRb -2��H�����%���y"@_,�����b�pB`���b�y2K�a���V��� z1�4���yR�ֈihj<���ߦ�����)ܵ�ybM�/("�\j׬�3Yn���L��y2��-%C�!�§�(f�Qr���yr㘄J�(�A4�$3���(��yb� �N�Q�3�њ�F��@�(�y2!˙/&��d*[<��팖�yB)�7nm��6����'$�y�,���|�a��ܴ�&���y��̟8l*D8A�ޕj�d�v���y�ՙQL~|J����"�`����y��F�sQ��֪�7y(�=�Ů�!�y"�P���1sW���&E�1�$瓍�ynӤ(�J���MJ�
��e�Q[ �y�C��ʹ�p)�Uj�����4�y�eO XFn�b�3J��M����y�-��`�iECO�<���xpN�2�y�	�:S(��Sʗ�9�"(��HŤ�yR㚈%2�b"��1x�Mb+׊�y29�*��7/$7��D�p�_��y��*��hGe��:���1uf
�y�fXt)��H!�\>�8ѠweG�yB�_�~�Hұh¡.St�Z��ι�yB˒<G�۠$�- ��iع�y�hK)6]
 i��:\��B&�΄�y���9B'.̑EN�^����u	M�y2&�s�f4�`܉@�@�5%U��yB%U�1�B`�Wަ1RFE#���#�y"�7zkLU�/!*n�Ӥ�Y�y2�F?oxnI�$OH�m(�q��M��y� F�"~0�R�\�o�����Ό�ybc@)SZ�!cǩL�eL�eV.ݧ�yb)W	|X���P�*}r�Ш[��yb��V�@0W8%3�xK�� ��y�@�^@�p&��#n�Hu��y����N<��m۫l��I���y
� J�H-]�H�����(1c� �"O�e����)��Q�LC�Siv�0�"O�Ɋ�%�2�P��l[�P<A��"O����j2x��٪]l�i��"O|����͢0:�H�v�ߘIoi�%"Obds��
m3B��"H���"O�mHЃ
$!n�љ�ŕt+~�ar"O
A���.oL�H���c���"O�)r�N�?=L�S�Cwι�@"O�(fe��'�t�t��N�P���"O ╏��=�b��`D��aYڨB"O���QL^����;>v`�`"Ot�׮C���$8b�$|&��"O8e��*�:�����q�i��"OZ��"��Q�Cd �-����V"O$��Hh�0Tsw�$�DqAb"Oj|�p��;LW��ASEL4B|S�"O�q�A�,X�@����	�F1z�"O�hq�JP�4���L�	��9p�"O�����$1�\سbI�,�^�b5"OT8j�(Q�Q� 0)@���Ru(�"O��w�|���@����U�B�!�7Z)�ĲP�'�:�I�/��!�Đcv���5�Vw��)�f�$]�!�DK'[����R,<���c�At�!�DX�lnl�8㊌<�$%���.|u!�G�eJ�d#���TZT9�G��/h!�䟖69��z����?��z���"Ai!��͚:k�1�5a[l Д��#�qa|��'�ey�cN�5� �2WhyY� �PIH�"��X"j2<O��d��&M	YSO7c��ɓ��>�	j3��40oL �b�V!I��y��P�#��z�I>0v��a�8pIX�DG?zdR0zw-D��ta"f]�o%�L�`�:E��@�"�/�����o�8��c�#��s✽|Q���Q�H���IAy��'s�O���U�b@^[p�笛�A�,@��'g����	1��d��M\�c��5��'�b���ko���W�8�����z�=�L=2���`�_5t
6�0p�Ƃ@VqOf�DA�
$��}��*�N;Cĸ�A&p���(����'N?��)��B��(O�H1!��^&	�� ��4�d���!�OB|Pc�WݼIs!.��w�Q�g�H�'�F�9��ݛƏe�����~��(O�qg�(�G�,�4]�ǫ�+�R��4���j�Ҥ�ƴ\�D@[p�"@��|�BbӚDn�����G+�!1�6��`kB>L�Aa���XCҍ�_/�E��ky�Ol7-3����Є8��@-䅘����b擏*�4�e	�PUt�I�H�6 �YIS
MW������9�m�3;_d�[Co� N�6�P���BeeǕJ"�Ӓ"Ixu
1/�c��3�O�OD�+�'�"E�ק զe���O��mڃ���O>7MY�T�j�6�X�m��
�7���Oj��D�cD4�x2G��,�yi��͔�	˱�,�	��M3 �i=�'p�4���m��m�V4��"Ç3�����Fy"(
�=�6M',O<(1��N�s�@�9����b�@J�t^TR��	E�V< �4p�jxX�'~�=�0n[Q�I:�n��6h_"E��Q��͖D䔴 @LJ�Z��Yr�/�)���H��~"F�|�zc�4��I���I���NlRA�@X��?��ʊ�?��iH�����OL�;^ ��XT���Q0]\����O|�.)B-hǘg(�;��-�M�ܴJC�&�|��O���[�Թu@B�6Ԛ��w+@�"Gl=��÷ �e����nx�8���
���+�΃4I�	-�(�p��E��1D����J\�@��㒈I�nz��
W�'�Y�$��L��s��̋A ϣ7���'���Q��l� ��&*$0�S@�Y�A� �鉨]v>�$�������wT:0A�/H�+٠9�Fn�]�Iӟ��	c�S��F�0���KH
-{
m����y��� ~ȥ:��$�X�)Y �~r�q�j�l�xy��= 7-�OR��"0dD+z�`���!��{84�H����OP��j]��M���<o^-Ȕ�#Ъ�k���:;���Vl�'�x�kD���r�<ÍɀO�t�U�܁ӠY��L."Ԕ�ݗ*ٚ{#nY�=�⨛$�I�QJ�Fz2�T�?��i�T�>���ٚh�t��R�H�z�Q����,��ɵU�RAȥ���0z�	��i̩wO�'��"?�i��6t����^�j�8�1+ظDp����>���?�O>q�}
�s���   �   )     �  �   ,  �7  �C  �O  '[  f  �n  >{  ��  ύ  )�  ��  Ƞ  	�  [�  ͳ  �  d�  ��  %�  i�  ��  ��  ,�  o�  �  ��  a   � � ]$ �- V6 �= �C J �L  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�CJ�0S4���T:
b��'�V�)��/r�<��w$?��P� �d����d<?��A�7�ٸ& ģ#26�rԥ�]�Ij��P���	'&Ȏn"=�#+<O�㟘�SC�Z�\�ʐi�xc��p�"O��3�iJ
�	�ħ��\���+�x	/���OJ|ɂs��*)��ҋ8g�\B
�'T��T�J�^H�{�E@6v�����}��'4̀�)�_�r�)%�?s^u		�'t���Ql��N�1����� �:�k�'����O�Js&|0��Ʀy%����'X�,�&@�S��@)���p�"�A�'���XLK=�z	I"dS�sC�LK�2"<��k�� ��0��*��i�pfe��<��ne�q"N�\茔x7�x~�P��<E�� vhm1fj��y���ab�;�y��4f|�tN�m1r�S���'�����	)IA@����0J�ĥpd��xC�j�6)Ȳ��C r1�E+�3U XC�I�*86M�3�?L���� ���#ғ'<L�'"Ζ3�0؋�+C&,�1�ȓd/��A�8c����0
�%ܑ�'ˆ#=E����?>y"#�A�+i�l�߅�yrJүH��rTO�?C�|#U����0>�R����-���ՕQ%\�bǋ_؟���'�pQB�Ɵ�1j%��͛#p�ֵ��'��ha�Ȉ�4�Mh�iӭk�j|�
�'�"�4L�w����c�";�z-�'[N̻��"նeX��/0��-��'.�m��GҼ�� ��C�}!rAb��� 2l�e��CL�qF�-gT@ �R"O\,��N4)��E� c����`��'W�gDr���
��r	��`cN�M���ȓLVhw�%e��	��L .�T�>!����$Ox;"���"a������yҍ��TL�FΜ�[��+���<B��'�)�3�X_����4)���9z�Oڣ=�}tO7r��"��A����'�Cc�<�+�yg֡9$�F�ueV��~,�tD{J?��H��E�BL�%�Mۦ�1D�@I��^bZp���UT���4ړ�0<	n�9D>�1�Ao�
a'\M·$ \�<)�FO(	=\:W�B�3��ñ��O�B��@� ��BIE~,��c�Z`��%扶zW�@��@�s쉃)ϔwxV��l�����jBN	��4�CJأHئ$:��O����K}b��#���QdjD�;W`�#%	��p?Q�O����h�:��;e��4������IF����kI�;/M;��+�2=� D� ��ꁿ~\ �Z�I�7+)X��<��ȟ��hTd����!��%�!�#"O���s�>A)��c�S)x�P͢�;O,�#���SܾT8)�-ځx@��vO�y�c�)i��"�H"k.��(�%W<���qX���u���4��iR)U�/8|q���>D�xcЯU�y0���
�Bu 0�2D�4�F(S�C�&����"&����1��ȟ��p��P�fl��ꃫM���b����<��iSn^e��H+��1`��&th��Ë="�O?7m5R�-(���B�ݱ��[�'��!�V��~�C[�7�v�Y�� I���i 7�y�$�p3t����(��2sOP���'��{���d�b��WB��)�%2��=����>��'�9��5K���`�]`���'�=Pa��62��p�$%Uq���� ���<���;xHtD�!��Kk�%�UiUz�<y���[
����L�N�3�&�}y��Bj��(��M��O�����6,C�^���pr�'����@��M
I��p ևr�^�#�)��a��`	���:D�4�B��mU E�(ғC��?-���ɍv)�5RfԖ[&�鐔���yrA�=Z E0D�N�v�Ӄ���y��
p�4H��E�P�t�PJG �yB�ҋ`c�ȱ��wWyso�����<iH>���ɝB�R�0�BH`W�Eãܽs;�B�I�y@LR�G������.p�C�		7hu���G+(��ݰ���;z�FB�Ʉ'Z,\� ��,��I�/M:0�C��
	Ҏ�ۑ� �
)2��J�v�OF�=ͧ�Z�&w(�:��Pb��钠�;�*��ȓnZTPXw�B)5f��a/ȗMψ�Ezr��6�ȟ&Գ�6W��t���['hsj��"O�X��DN�p�W�alA� �'�ў"~z�%U��N$!��L8+b��7 W��y�`%5�(��#���,h��K�yD�!c�I��iM0~_�@�]�y���P�$��@S<jt�1��'{azBG�k�}�CٷD҂��SIЉːx"oJ�z�����r
� ����f&C�	�L��ݳd�W�\ǌ� ꃵy���� ��7����R�D�c�4�j���#��B䉍T=T�a��*OG4�:aoJ5?���	V~"ʞ�O�OC��� �-`r}�ț'~x��?�+O4�c���6��}�R�/\0��W�ɟp�ax
� ���/�P��G��x�(���+�S���Oy�LP�2�� ��Cl��O�u��b�"�t�s�ֶUU���"O�U��G=���5�J%���y��IK��]�'���R�B�*U(��?G����>(l,��dT���q��ݘ"5 ؆ȓL�@ac��Q�B����y���ȓ~��{f�Gz	��惼#"|�ȓ]ш��Q�]|�\�@-G�$���'kR��d�!x�H��49����8|!��ֶ@���j��*<�L��@�:!��޿k]��H��'��&m[�Q��E�D�U�/�tHH�4q[�ݓE��y��C�����`�:m��f���y�%[�P�쵣���85��E���^����O����J!+���R��*h�D�k�.^��}�aF}2�R�Э�Ħ��*��	��	��yr�ƒn�
�9�*E�$J���c�ݲ�y�m��|{ƭ���=J>��S��;�?ш{ni�>��'pm�"4��]L��h/rMh���s̓tt�Ӣ�� I�y����&����=,��`p���VD�Q�X
_��$��l�I���O��q���h�j��GK��y�\[	�'�ቅ,V�I�r���U�ZV��yR	I~��;��/�|t�� �c�:q��"D�\���?i���c+��%8t�$��>��$�Rp�WF�5$P�rS ím,��G~���1 3j1#D�\%0h��3��7����>I�
ϧ.2��ä�"+�����^h�'�$%�T�\!�$Ǧ��˃a�;OK��ȓ��V��JF���'~!ī�}�<��O�rJ��* J�e�D4JVS}�<���8���iѺ �"M%@�a�<���b�v�k!�C�Bښ���\�<���R1�Y8�HѬq�5��R�<���Ȳ PTI�+�%Y�J|�F�Mx�<�uf\n����)G�D\PhjTn�<�֣ߏ/S��+R#\41h����|�<y��J�I��Yy�H�T7��kc�<����5w]Ybm̵�s�F�\�<1vj�?�~ ����&(E�����Y�<�5�� }'F�"�cƘ]��ѫ �HJ�<���A4��l @&jтpCL�yBB�/�tI+q�)7jnȪf*˿�y��	AU�!�c�1���FbT��y�IG
Hyj�9�b�+ϲhɤ#���y��پh�e
!�0^":Ì��y�h��6�8��Ë�<=��*�Iߑ�y���I��r"^�0|ڡb�i��yBA�)�&�k��	"0��	A�yҪ	�n���؀MC�'%4���B�ybcA�ho��� 7��*�� ��yԈ1s���A���2��1Ӏ㓊�yB.Z\�eAp*%Q����G��y���jd}� OF�,���낆J��yBP"B�ʖ@�^]���yR��2U���1�Ç��lsҭ���y���,L<^���!�ĸ�tW��y�#�:;�Ya��_��<a�j�$�y��- ��Z�)M DD���F2�yb�	,���۵l�J3퉢�y���+%Z(��x��!X�yR��o�,��R4*=���yBO/|hz��@�U�|ٲ��C��y
� �� ��ț1Ը�N�$e��+V"O�Y7�EiF����J)t
��u"O�l�F��,��V�J9W��R�"OM�#�2M���d	ǃ^SR9 W"OV��r��}��3���a/pӆ�';�'{��'���'�b�'�"�'5���l?;��iFY)}0j����'�b�'OR�'m"�'-"�':�'�H�x�Dw�x��)�U8��'?r�'��'���'��'���'�xE�4�\ЅAi�v�a��'�R�'���'���'K��'���'�pm�%gM�yb������7z��<�b�'V��'Ib�'B�'��'br�'��� ��Q "f��p�S.%��P*�'�R�'cZ�M����?Q���?	���?1v�Y#8+�!k���/���A���?���?���?���?A��?���?i��FC��ոR3;�zr�Dى�?����?���?����?���?����?iU,E>|�Б�`#����˙ �?	���?����?����?���?���?�BΜ8�b��a�ڷ���Zf"N��?����?A���?I���?���?��?��cM5b�@����".��E����?��?)���?����?���?����?qD@ЃBP�A+��F�Wg�T@1�ڑ�?9���?���?Y��?y��?q��?�b��uWʌ�'�W�QK�	����?��?��?����?��rJ�v�'t"�8�fd@��Ӡ��asj��Gs�˓�?A,O1�����M���}��bG$�c�8��`*]�'Q�m�'
�7�"�i>�	Ԧ�´�A����ǟ�eD�;r�@��M�PӤ��H}~��G�e���Y���]�IB)!��X���-$]��1O&�$�<���)ͲYWz�� ��[͘k���30Ʀ`oZ=',b�������y�eޖD�t�jWh�:	����D ��,Y��dg� �	pyJ~26h� ��͓]R�,I�o`�\����n4���y��<�tN� 8|��4�t�d ������)P0O�d���%��D�<9J>�#�i����yrF̓a���Z����. [��	Vf�OBH�'�R�i���>1�J[=n�����G��T�VuAf$\~B�rg���am�0��O2��c#�H<%g��_���x���pm��J�%-��Oy�������*�j�;t�(#��}c�3�����q�';?�i�O�_���%qUe�&8bd��/���O�6M�O�-@����IG\�@��Z�&d�a�^�M��}P��D���s L�_����S�`%?c�h�<E�Hp�ĕ'7�\����!?Aѿi��8R�y2�I�
�V���+�pb�C�`��|�'�r�i	�#�����$��N�P `e�WB���%�B����l���He.�SG���:� `#�>ᷞ���ӂ��7�
�L�
b����Q̟̖'e�	L���Mc�<I��8!G�H9@aE�C���+b ��<q$�i�O��O���`�8�$�. +��Iƅ�%k�蠤�>i{�`f�̜df�Ħ��Cŗ?|����O��) �S���U���V�'w��ٺtK�<Q����Ĳ<E�D
5x~��f�*�*0*�DƂ��'�6폌M��*�M�O>iQ�Ȗ3��p R��< �q.�y�X�hl�M��X)x��B��<�'���
 'Ӽ{�Z��a��(�|#����t�ݛǨ�j���dS���I�[�����o� �T����x��	O�	:�M+u��Z̓��#�0I
v�0BF0��i�on�	���D�O7�q��'>��S	D�l�\"P�Ti�Ab�S|�6�B�I�%�T�d~��O��9�d)�3H��'k��H6$Q(x�h���*��(��'[��'�r���O��I��M�Ӥ��S���A�iP�l�H�b\
SM�� ��?� �i��O�ݗ'J�ֆO;U��q L�MΖ��Q��m�6-Væ�h�J�%��R�e��3eO���+O���!�s���3)�|���7On��?���?y��?A���AZ�{� ��m��\XWf��#]�UmZ�pT�Iҟ�Iz�s�s���#��>6�y�� $�pE���MbÛ�e�f�O�I�R�D�3ll:t{�4O�]J��LS^� �7&2�)�6O~���%*.Uxh+! �d�<�'�?q4��<EL]˲��<7(]�Ԉ��?9���?�����զ5�r��ܟ���(��ӣ�������J .�p��r��v��ɓ�M��il,O<����"=�=�M�)<�7'8?9�D6D�h��Ïݾ��'{�D�����>�?���?HS�L�� i��7ş=�?���?����?�����O���%!�ܜ@�d��'
¸����On��Ӟ�	؟�P�4���y�8!$�xVBX�#R|�*�ÿ�y(a�veoҟHC���O�H�I�(�'��� �ٴȃ���xc⫂9c;�Cة3O��%�����t�'�B�'�2�'�ڽ�Cd��pbR|��GAa>,�C�]�`��4
�)O��D-���O������ 8Sh�� �`Hg.�S}�z��Qm�<YJ|*�'�?9f�ى�^���D�36D5���*2�����X@~� �R��yӣګ \�'��	R�v�z�`J5 %���5��,f���'���'O�O��	8�M���ҟ�?)�G�� :G�@,KJ������<y��i��O9�'V�6M��5�ߴr���;
Y;(�Zh�/�����*@ L*��]ϓv����4\�zq5�Ԡv��O%0�%��� lU�'�]+#�(T���t��9O����a���������2R-�/ev�!���-�����(O��?���?� �i9-�cT� ��4��u��\2p��T�4`��`��zS����x"��O�6m��hܩ���"���O�7�
تp�g��^�8!��Ɵ�(�qq@ �|]��%�l�'{�'Y"�'8xa���V�l���dL��q6����'��Y��@ش[�T�;��?Q����)H>�A��d�g��t�y���#���O�����4|�����O�$d ��[ Nc��� �T4W�x(R�iN
� �0p+@ʓ���!"�V�K>��Q%�&��E}b�#d��?)���?1���?�|�-O�%m���@��,?�`L���ڋ(/L(�Q�ɟ��ɔ�M;��<�ٴU� �e��9=`� �4bB�[$�i��7���~�hA�>OV��w��%`��/C�q�'/hL8�H�g��8��@�c�X(��'���˟�	Ɵ��	ҟP��r�tb\�XV#O�sU�u����77�7�FR�l�D�O���$�9OHmnzޑҢ��"�\�)���%h*��'��M���ixLO�	런�陵-����g5OpéU�&�4�3C�i���?Ov7-�@b���i\e��^yB�'�"�O<k� %�Ï��U"��r�o�)>E��'���'�剥�M[R����?y���?���dѾ�s�J�@�:W銚��'+@�D؛�z��'����o�^~i�����5�LH;wFm��	��9C�C~�X@�+O����;��OŸn�9�T=Id#�=���"$�O(���O��$�Ov�}B�W��qBtb\�G�T0$�F�j��_4����-�r�'bB7M6�i����΀l��I7� �w� )'�a����4(��}Ӝ]p��M�7O��O�6MS�u��E����`r�����%yA-��$�8�''�'��'|�'�d���I��Qp c�ƞ�~�Y6_��X�4d�������?������<	v���@����
����Rk]���I��MkĽiPl��<�����[�O�+���dt��*��<�pxj���9w��˓�MC�DR�L+ƕE�|�T���A〹f�I�4MT%��!*C��Ty��'�����]�\*�4PdB��u�hç�	^�t9RuH�IU��͓QI����_}�Lq��am�8�M�s��X���(��N$��8�)���㔭�<���M��`�P����QR���S�ߍ0�iӼ<V�,�$!Ќ>4e�Cop�����,�	ȟl�����"��4�4QXb�U�|4�)��ݜ�?����?��i��q�CV�۴��yJ4
&�ʑdj�A�����ї�x�H{ӲHn��?�7�I�2����Ɵ�o�`,j�3$�h怼q�C�k�p`�"E-Et��L>�-O ���O���O��HD�ԐK�����F�Ud��J�O>�d�<AP�i2\�I��'T��';員I����(	���%� l�Y"����M3�it4O������p�j5�E����$Z��!e�ڬ���7
��5�'>���Q�� ��ǔ|����cD�@�$H��<B�����C42��'��'b���W�̰ش*���(�u-��G�>X$�x:Q�L;��GӦ��?��W� lT3
�YV�B+e�\:Ůǭ] �)ݴ%ț�+أ/�L�;�'\�i���eҨS=����q����:(��C��ـ@��͓��$�Oz���Oj���O�mZn����+lv� W�ȟyS�k�.��J@7��c����O��d/�9OJ�oz��Ӵ�B8.�ab"�[<�>4spH�M!�i�����>ͧ�b��0C������<�e���=_,�X�ɛ- ���$_�<i�4? 	GDSz��'8����ɟi�04�u�׾EkR'R�o�t�	ܟ��	��@�'JV7M̍�����O��dԧ����K�):th�C,F#N�@#�O:�o��M���x�G�W�ݨ�/^0��4���y��'ӛf+�F���[q&�<)��.r i���?	�Nעq ��@���'*ͮ�;Yf��������I۟@�	N�O�̚<�(���m��,���/4�R�`�lk���O>�����]�?�;D��`�T��b|i ���>p�P�.��FbӺ�oZ��ZUGd���צir�O F�|``�چ?����S	C`�h��`J������Oz�d�Or��O��dJ71����n��if���A�Nu�ʓ@śƍ�$A��'�"���'�̅�R�]�ov�PDҕ�]��b�>i"�i67m�y�i>��S�?�0rA#3_Yr��,�����,@ge�Ca�uy�i�˓%י/�.�O�ʓHU�Q����
>9kR�B ��@-OJ���Or�4���'��NМ�R#G�2�j0B�ƾX�D|��8�yR`���d��O��lZ��M롳i��1`D��V��@�UE_#�̤��)	�a!���'h�i6Zك���G� �����(�b�A%A�f����TM)�d̓�?����?��?�����O��H*�l[�T="���%O[�}���'��'g�7m��V��O�nY�	!:>d�c !��M������R� �0�K>�ڴ_���O���D�&�yR�'�����7�Y$Bݹ3�@�,.#�
h�	* � ��|rX����Ɵh�	��%F��2������+r�� �l�П��	oyB�b��Ă���O|�d�O~ʧ(��!�&�6|�X[�?;J�L�'4���?��4vhɧ��'�B� �+N��Ƞa N�e�r	A�4� ̙� �i`��?M����^d��$�$�F��H�4Q��̶s�����I͟��Iܟx�	�b>��'3�7�X�1�P�H�#��8j.��Ă�oX>T�4o�O6���Ӧ���G��&��ćצ���[�U�֠�	5b&<h��L��M���i��=�î�	�y2�'��f[C=�k�A�<� ƕ1��.���)0j��8Orʓ�?A��?!���?!���	Ց%F�M0�A�@����F�7�$Qm��	&=�IП���h�s��������ȝ�����R�a�Q�䯞,9��V�c�b�&���?U��
h���Wq�$�$�[l�0ʇĄ+X�Ti�Fa��m�՚�S�	e&�O�˓�?��5�4�"�Βj�Ш��oB������?I��?�-O�oZ*��	�t��-3�k�LU2p԰�3�A�!'���?Q�W��۴��֯$��G�
�R��'�$gR�U`bC%$�S,�L2��^�mE��J`c�O��o�M9Tj,�����(��Ic�S����P �Β��?���?���?A����O�̫���Ny�e��_�
�af��O�lڇ/������x2�4���y�i\�k��a���rr`�)4 B��y��nӨ4l�П$�4j@;q���	ܟ����ў
o�|:�ߪM�1�N��BژM[�OГ;���&�D�����'1��'PR�'�|��u��R	z��ީ@� �6]����4������?����'�?��KZ^9P��զPϺ���|3(�%ߛyӠ('�b>�@P,>f�I��[�=�j%���JgJ"��qb�Cy�%�/b�q!6㇙!B�'a��CJ��Hۅ.�"�1�hU	������<��ҟ��i>y�'q�7�ōaÈ�O�yN0�B��^u�0��f�)5�������?�t[��+ܴ����'ۆ�C2#W�uĬ��O�(�}	�$[�Dp���'�B��%����p����d䟲�1<�0`��%sܨH��
�t���̓�?����?���?����On�tC�-��#d	��H|-���D۟l��˟؊ߴ{<��'�?�t�i��'�(��Te�t�����חy�6i���"��C�9���|��YLF��'�(h�4/Y-2τ9ʱφ
� ,p�+��������س��'����D��䟀�I�l�H�d��Vk8�� O1J7>��	4�'�7��49�d�O�$�|B�/����z��E&/i��	'$�O~2�>	��i��7��c�i>���.W4@��.N&9�m�!I�	:$()��GlL����vy��O|
�sa�o��'W�y��  ���u���p)<qh�'}��'���O��I��MK�ؕ�t�{�m�)iE|9Ӏ,�t�XM�(O$�m�D�oE�I�MC�L�:�b�	D)TqQ �J�����'�� ����*�y��' �i���x���O�����ƞq����%a\����<Oh��?I���?Q��?�/O�I֏;v\��D�s���"��L3��lڂ6�$�I����	l���l������=._�\����:kU�e���4^Z���;���;X�ȐaQ4O�}�%Q�KP\��m�4���:59O:u���ZJ��\[B#�ĺ<����?��
�&z�I��L!���L��?I��?�����dZ��r�ϟ��I˟�k£_0oҾ%*�5P�n�æ�}�I��,i�OhoZ��M�6�x��X�ܴ+F���}�H]y�N��$@��n��Jě�:����Z���8���dZ�!�����3� $�4�
�����Ov��O6�d9�'�?�� CeNR�E�*=y�9{��'�?�e�i��`x��'�c�x�杋_��"��Z�%��i�h��E��I	�Mr�iI�AHV|��'aR�6X`�b�4$�i]	T<8"+S�,s~P�CM~��~y�O�B�'���'��MFL�D��L�A��Q��)q��ɼ�M��ω�?��?N~ΓA�Z�`&$�@�ְ�%��b�Y{�]����4!]�vl!��' d����Ņ�g�4�qeo� y�hh���,`��O�$�s�`��~�yI>a.O�-뵃�l1h����}�b�$�O>�$�Ol���O�)�<aжi|Q B�'����/��e!@�Ȧ�֥d��ز�'<h7M$�	���D�)��4QU�&L�D>���"(Y�_d�4fB^��D�5����d��@t���MG�vY������]
s�fL�P�Ǆ^�\���E�pl�D�O@���O(���OX��#��0[`(���F�]�,��C�� �	؟��	��McuHX�|J�� ��&�|��9h}��K�Kn���&H�/1O�m��M�'T�����y~���l�֑�&+S?���"F	ɘg�C��D�:���|�X��	⟄���h��*C�uq���ћ=t�=ig�������WyR�Ӕ�j�A�O��d�O��'e��0�	�lA`��+#���I�
�O��n(�M{��xʟ�i�D*nlh��#[e��҅�\�v�Zi���߷Z*��|�fm�}��	�N>1��=$+��-�	�"5�14�?����?����?�|z(Ox}mg�t��$�͞R��iAT��a�,�p���Ny��wӰ�XA�O� o"4yP�SrfV=ᚑ:��c�
 s۴~I����%D� Q�O�%9�+��{�@�	 ť<�r�&}�`@��42g`,ɔ���<�/O����O����OB��Or�'9��`Y�R5~�P���>��uCR�i{"ԋ��'��'p�O��z��.�9@� lbcR-�S��N�2o �M�x��� \�!~p��'cd�����>J�"9���636=y�'�i�Ԭ�z� �j�|�\���	ޟ�"%脰/?T�q�h�� ��	�Ȕ�d�Iݟ���[y2�i��=Hw��O����OV��4 	�=����mHfvxD�aJ%�	<����1sߴ Z���
�Gݬ���˘�D8����5?����3V�`1� #ȥ��'k�Le�@�%�?y��P$��(c ̕�k����mX[�<�@���o�����F75ZE�WK2�?g�iҨ�'��-v����0r*I�S%� J�0�b�C?4�"�$�M��i��6M�e����:O��Z3
��F�8�� �͓#!�,0���`� �+W��Re�0�d�<1��?Q��?Y���?���D¶ R ��)X��C�A����Ŧm�����I�%?�I�.�8Q@� `�}aF$C�M%�Tb�O�mڟ�M���x��4���8��a�#n��Di�A!4�:X;F#�*��2e�<� L�Ny�%�4�':�q%��9Rv���nđ~ܰL��'�B�'������]�4��4	X����hk*�Q�愨���,Y=|��q�]�V��Z}�x�p�n�4�MK&"ˢ$�i2��@�K4�|S!���!��Nh~�C�*�\<����&M��O�'*��C�tݛW�o�������y��'g��'�2�'�B�I��\�*�@��95,�Ѐ�P��2˓�?!E�i%*�O2oj�X�O&���M]�aĂ]�U�M>��ՒV#�Y�I��M�3�i���c�e�����'gb��i��{c�X�/়S)3pq������8r���Қ|�W����⟘��؟�y�-��>�̼�'k	�e<�%R1 �ݟ��	^y2+gӌ<�U��O���O˧^ք`�D��l��ܨ���3v�!�'R�Λ�ez��(%��2� h	�H�=u��8��D8c�Xi�ޔ`��ls�K��4�v�B�HE�%4��O���Q,
�i��ܠ�*p���O��l�[�6`8��
\N@(�A��������Ɵ�����M��b�>�%�i0�*S�:W���I�no��rKp�NoZΘ`��<?�EV��|�ؔI���D�i8� �؟d6��f�
n@�<���?����?����?�/�(�	7�"�/�7
X*�1��ئ��p��L�IƟp��6��y�숀E+BPC��B9om>)K���|ˀ��dӐT$�����HA�Q%*��D˘`�4ZD�A<Z����
�(���C�5����&��J2�O���?9�y��|���SM�@!�Ax�][��?����?�,O(�n�&�h��柜���="y"h�%%R�"'��
u~M�?�R�x:ڴ+N�V�<�Dȗ7�V�ԬǳL�tuq��'Z��	�gyy����L��9$?������N���I�<�� ��1;�$�(���,MЀ����l�I̟���P��yÑ�����	�E
�̃7&Y=��nӶ<��(�O����&���i��� ���<�t���5�tЉ�����	֦�C�4/,tш�A�K~2͔�,+���,
�6d����<}�����|2^����ܟH����L�Iퟜڃ(��D�LA��ҽ{���e@oy�f{Ӯ�� ��<1���'�?!$-��dL�b�B�$|�(pG	6$���˟dl���S�S�%� ���K��p���7�MI���	�[��I�'\$e��I�Zdf���|���0r��[�UB�H��e��E@���O����O����O�i�<�ҼiW �Y��';؁���A �L`'&M�#Ū �'ir6�:�I)��D�ۦ�ڴ��-�q����C�/qfx%���H�J�by�EDP���͑j�JUAqK�!R⒟���)�,Sen�q�R�E0�h�k[5�j�ҕgԕ3v�:���,�ε��+�&GM�i��U�Y=`P(i^!���BшO�p�9䤚ɮ\pࡆ�q�be0��QYz�ai�/,O���P�<'|� lc�U��8��A!�C�j���0�$[k�yӠ�(H��o	[��P&�2�!�1F�&r!��+pD "��?gH�Q��P$]������:��	�G�V���"��7H�@���5sI(5��h ��\!�*�8{8�=����zb�6��OP�D�O�=
�O�^�IΟ��Ib?�TUd�r���#��H���'e[Ԧ]��ϟL�	�C��d�J|2��?���T9V����N���gd�o����c�i��`���	��	�O�O���n	�"�č�E$P�,p�@[��_}2eB0~t�z�O8�$�On���O2��W��>�r'�%}�t�W*.��Qs��O����OH���O:�OJ���O@!
�n
8P�T��s�I�a-&uRc�4�X}���	ǟ����8��<;�T�I��ę��EҢ O"� ��Ͳ.���4��d�O��O�D�O|��f��!���F�X�yj��Q)�P����O��$�O8���O�D"l+,�'�?I�V��D�4MJ������;Q��f�'��'�r�'Rv�����ē�,�Xt�9Bē7D�MGn�l֟�	ȟ��	�a|�Q��ß���͟ ���&���G��D����&M�-���H<����?��k�E���<�O��C�Ǒ������:����4�?1��.2��"���?I/O����O����:}
�#T�az���ELm�\h��i�"�'>�,f ���<�~��ae��̺�A[�A(������j�&�MK���?���3�d� A��X��^`���.΅o<�4"<���t�'��`�͟J�$�:W� <m ɢ�&p�����O@�$
p{���?!��?i�'T��"(F$j��8���v^�Y۴��{B�{�����'2�',����@��(�QÄBZP���2��i��i����P���	ßt��J�i�%�I�=~O���@إP�8� ��>�$*����?���?�,OJI	�m��T�����R#hC�d(G[�Y��u�'���֟ '���֟�[�O`�0�hH5=-��	 ��Kj��	iy�'B�'��I�\b�%��.a�Ȳ� �0��a��Ѻ��UnZџ���៸&����៘i�/�}?a�`Ӡ(G$E��Y�H���E(^}"�'�b�'�剩k�8�D� v���@�w��8��WU��l؟�$���I؟�aD�P�,<F�!g��A��$��耹*��oZڟ��	Xy�쉂 �ٟ���?��'�(L��DY����kU.,�Ꮗ(�ē�?Q�r�1���� R`��%	��;��WY/VM��i��ɨ��L�	�@��ş\�lyZc��0#���f�i6��2�,�xݴ�?)��|��j���T)�J��Ȅ-ǝu���F���M#����?���?y��b(O��d�O"TR��іX#LH�Blћzf浒��N䦥bG��H�S�OG�j�)� !S�;;Ʉ�`/��n�6M�O����O��'�<���?���~��	sڸ)�`�� p�1�����'Ob�b�|b�'��''�)�{����A,�!1�VٸF�p�x�d��7�˓�?���?9N>��`,�b����KTV�v�$N�'(^�+��|r�'R�'g�,!^Ҝ��G��>|x���8hMI��̓�ē�?��������<+/P����ۣU�z}��ۛ)����O�˓�?���?�/O�e���|J����}ϲ,�%�'Y$��ѡN�H}��'yҝ|�U��"'ߟ$����j�l�� ��=L"(�#�����O����O��	�-ڕ��t��cS@���)�5�����K�(/�6M�O:���<q���?!�M���?,�"�����R���M�9�@Oզ9�IAyr�'^�Y�SX>��	����s���˥Qxtm��(k50�Aa,���Oh�dе<��B��T?�0Ӧ� *�*�p%�˟}0@Q1��>��;�P����?���?��'���>MB��Nr�t�F��,��E�s�i	��'�@19a�N����O��h��	-�ЙD�:}���4_�I��?����?��'��?m��-G�:V�Hԥ^+;�4t��ᇩ�M㤁ÚevD)�<E�D�'�����%�6�cU�&V;:ݫ!�w�����O����S:4�&��ǟ`�	�ϼeK��ի���V9!D�5A�4�?q���?��eG�1���k���']�dP0�v}��#�rJ��*�Be��6�'r��P^�@[��f�D���Ơ�z��%m�[����ao��ē)H^L�'���'R[�����
&�CR�$MX����K�{J<���?	������O��B|LX'.G�1N�zc��*�7-�O���?�������O��z���?�C7�-�FL�R�"�rE�p�u�2�$�OH�`�Iɟ��6(.6-�j:���<(�(���iM��'f"W�P�	�A��E�O'����x���@ G��PD�ū��Q=7�6M:��L��G��Z�@!� .��9�c�5\�t�c!b�n~���'��I˟�c&�AW�$�'4���5�*�_i��R�(�A��	���(�ē�?��v��]��RB�S�$N�5|�Up�M�R��DY�M3*O�!f��ЦIa��,���n�'�.1�#܅W�$�c�,��C8�m�ߴ�?��*�b@��O���Z>7�ΤD�j�DK�)�6%��ڛ���d�6��O��d�O���@R�i>)��' �mHf��i���	rb��M3��� �?����?	���(��D�Oj=!G��_Vq�*�%` �������	 ��9O<ͧ�?���c�*|Ha�(ա�oj"���i��'5j����g~�'���N�:2���W6O8R�)kN1Y��6-�O:9A	�j�i>q����Ė';2��rl�()���e�޺pp�*��lӌ�D˸Y�T�d$���O��D�<W!	���pT��~�� �cÇ"^�0<I��x��'���'��Iޟ��	�j$������Μ�J �iy�d���|�'U��'��Q����,��DP�olAA���3g����'������On�d�O���?���_��!�,/��� ��5fML)�q+�]8H`rQ�4��ǟ��'��_�"3�՟x����1*(����(L�[o��F��(�M;�2�'���_?#֐@bL<9��_�<V�-��
��@*)�������fyB�'�dA��_>����\�s�-H�'^L��L�� oR �Hc,>�d�O�����PT9u�T?�Sꅓx&�ԩ�-�48� a�H���O�!�^ߦ)�	럼�	�?!��ҟhy�Ř�+�0�0�ʺ
^,��C�S���d�OxD"���O*��<ͧ��S7�\ �aIN$`WbI�dlz�6��51��m�ş��ܟ@��?]�����I,Ƕh���� E8U�1�Ȝ,���� ��Iğ��H~z���,�y��B*����`R�(x��S�iN��'R���t��6��O����O����O�΁�LB��⩘ {����(J�3ě�'Qb�'`��!�����O���O0	�F��9$m8ӣ�<}�Rx1����5=dT��4�?���?���B��S[?�f�F<'�A!AK[9<"�l
�%�j}�*ә�yb�'8��'���'w��w�v��b�C�(.�Af��C�8`�t�V'�MC��?����?i�U?��'���@K���b��J�T�D��GS�<A��?����?q���?�vȀ�S�i	R��P�:��tMT6~����l����Ol���O����<����8��'(��1+�d����F$���� �i:r�'D��'��'J`AAigӒ���Of��G�K9Y|ɑB���t�fX�j����I�4�	sy��'�hH�O��a'TY#c`�c�&ױa�al���H�I̟��ɭ�P�޴�?���?��']�P��� 5e@�R�
�4��@]G�����<A�.�`�Χ���|nZz6ȣ�N�v���(?=c�6m�OV��)�Xo�П��	�,��?	�I�M���֌�]����0K�"�:�O����k��$5�4���Ok I*��^�	�� ���/1.^���4F����i+R�'���OZ���'@��'��Q"��F&�DdP��
Q��"�a��8 �e�O���<ͧ���?�s� X�y4�[�/9��v�������i�r�'�2c[�[�06��OB���O���O��ܽI���:���X� �ٗ�����&�'�	���)B���?��O�h�������b&I��Ŕ��޴�?9�㍓(���Lyb�'B��̟��쬋H�g&4�
q܈V��7��O�=�8O��$�O(���O~���O��$�/^L�[�.޴]^��&錰Y<|��k�����ݟ���ߟ8Y����?A���	��LQeV&q���ce���j�&���?���?���?y-��M�V�G�M ��]x��d��$�����M���?���?�����O&�xg6�����
q�P:S�����P����'����O����O<�d�O�ɹ0��ΦU��埬��a5y��X�uc[#\ E���M���?a����O�\�@9�X�'Ū,��+��i�킚MF�P��4�?����?Y�a>i��i��'`��O�v���Ǝ&[��^�(��n�����<9���]�'�?�,O�i�r9���MT�Q��(��{�v��ݴ�?���t��Y�G�i�r�'x��O�4�'1�H;�l�dzTh��@����>)�V��!���?i.O��#��ѠVrP�I���M�^��bV��M��	Z����'0��'����O	b�'@��U�Y�l���JP�Ow�@*'R�]��7M@�Q#^�d�Of��|zM~��^6�,b��3k�D*3��1g�L0�i���'m@�.�`7-�OP���O��d�O�N�|މs��ٷ@:�}�r�
����'L�	3:�l�)"���?I�O��"-��Un	 Ď��DjԘ3�4�?�P� .}��'�r�'�ɧ5^�ݐ�(H�/	R� ԁR�@u��@�O�e�O���?��?�.OV�Z$&��t� 90�-k����lmRE%�8�I��&�<�	���?r�~9��ƖA�&B؉y��ry�'=��'��Iwp�=��O3�m���)=_~�Җ��2v� ŋ�OB�d�O��O@�D�O���#�O��#�țnGB�:BE�zD^�j3�W}B�'�R�'q�I�K���K|�&��'0��r"�'j�Դ���ݨ6H���'^�'l��'���'v�ꖈ�#'�]��1�M��`�l�۟T�IPy�*��r�B�2������z��V���0�t�ʌ!�(�b��F��՟\��#� #<�O�ZY���j�5�fJ�)>$mش��;z��Emڐ��	�OP�)�T~���|�d��F�-v �#�A=�M���?Qt
��?�O>�~�6d�/Q�
��c7LZ�[�� ��@C�ڳ�M���?������xB�'�~�0���� �f"	�t�� iB(y�2�r�0OH�O>	�	3>3�!��/UX�q�$�	@�)�4�?���?v�K�^��'t2�'��d��Lp�KwiU3u'tY	�#g!P�i��'�n�#�6��O��D�O0�	��ғ<	����[	F���b��Y��'_4��0I<���?�I>�1��@j��@Ŧ��	��� �'�T�9�'R�	ݟ��I��L�'������#� �ω�Ű�SM��O���O�O��$�O����&Y�,#Ca$|�
L���H�D�<���?�����$\�4��ļ�483,K�Sne�5ʕ�n$z��'^b�'��'_r�'�rhۚ'�Z�
=,U��f�,`�&Y%F�>����?�����	1��$>�Ɇ-C~FPáȂ��nicClO��M�����O�r�c�O����?�K���<��.)��]��`Ӵ�$�OR�C^a����'�\c�p�s�B������K?X�9��}��'Q\��'X���ɟ��1��)Αd�"}9��)Hܛ��'�B�0(�"�'=�	�?-�����$J���S��.[�*�j�	Y�4��6m�O(��ցvU��Pc���&��CA�	q�����ʀ�~�f��z&6-�O��$�OD��D}BU>�0��"(��5�cHߺ��7���M�D�����'��Ĕ|��'����U��:{&h�ჵoVDXÐ.j�,���O:�DرC����i�O����a�|�t*��-AT��&P�
����y���I@���$�O��	*Pa�T�𣆪���!�߇H7��OV���A�<�@Z?)��~�	1�!��Būlj�٩���?_a��O�i��.��{��Iݟ��	��'��M�&Y��i�?@یؙ1O�m(O��D�Ov�O��d�OJ��)��֬Ȕ.U�H�G�V�1ON���O���?�bG�.�?�A��t@d	��7o\0	��Yn�&�'$��'Q�'%��'�Rd{�,҉�?I'h��n��UJ	�;}4�W��>����?y���
�+��$%>6�X�}n��.Lf��4E�8�2���4�?M>Y���?)��Xn�%>�2�i��7����媂JJ��oZƟd��Uyr@M��\�,�d�"������F��S��2	�$Ig x��ɟ ��:=Ȭ#<�O	���Aa7 ���E[* )�U�4����$ղmZ ����O�)P~b���c��[��Ӑ{�T�Z����f�O��dŇ0��b?�rd�,@eb�"��L�$�9�~���`����I�X���?� M<��M?����??��B�-J�Y��3r�i9h����ޟ�YT��h�UX��c~����M���?��|�>\���x��'�B�O��e��3q-�:���
fb�C4�$�9U�1OZ��P$ݥa��q�EIZ�Abu	����Y���B���L�yr�Y� ~���6���'���ϓZF��r�ѓh�xt�gbOpɅ뉴����dؑXx�q0� � ��	�v ��RM �N~����Q�(|��Î�0�l`�%�ɞV����5�b(�xk�H�b&p���e��`aҘ<8>��֎�Zfx�sR�F�7h�rᗡ|˂�Ȥ�/�`< �cג(d�9A,Tt8�ARa���>B ٗ�Z�(*,���s8:�c��O��DÝm��D�O@擯K�d�/LE8�9��G ����FFre�Ս	"p��`\V�'���Q���"f^���3/_�a
�	0�D?Jh$���̱z�}�C�9�џ$����O.l�/��$޹>�NY��I'w����		��d�O��D8�)§s�r<i���"��8�N�?	����u�V�Z*8r z���4;3��6l���rP�����_��M�'�?i(��I���O�\y�ITi�|4 #�UE�` ��O���E���y!��[ �B�p���؟ʧ��I�	�E��{�2��)�
o4����Y�i��&���b%�2��  �Z�S�iM�X#q�ׯ7-b�0���:r�'h\�b��?y��i�O��`�b�<m�F��GI_ln,`&"O�P""`1OB$ �_�A+�'�v"=!7��2�r�Q䅙�#n:u�c��5ps�V�'�2�'� {�hʧ'u2�''��y�IS5|
4���,F�]�����۔E��Ճ�f ���y��Mvcb�X��I ��2���J����FH�j�փ^��2�m��BUҰk��.Q�P%�E��zӸ���3O�H�5f��J��J""�\�$�m�O"�7�x��i>�D{��CE~܌X���x���EH	�y��ߜld�ݚgIF'Դ�;U�́��$Ms���T�'}�5B�qxLH�A�Й���w��5��p�	ݟ�����hp]w��'���أY�j�A��W�z�Ĺ���	��'<(�p#�ƺp��8�Ck7�9`Dp���>yź�Z���,p.��c�;�a3*�3p���S��L�M�C�
b�'s� ��N(m�L	�#���Sp-��?���H̒�Q&٘!T��Q����1?���ȓT�<�I��Y�NF�]����<{|��<Q�i��'7r`{!�~��"c��`R����F ����������?���I��?����d�(=GB����С:�H�)��D
�1[�K�4�@�J�g	�O�b���i�UC��$�--�1Id�Úp��Ar�@�Tjaqb�7QRe+��T&���'zӦ���IY���$^�Yb�OP��ˎ\D͋rHZ��I� ���O���dҤS~��J�S��VF��4�!��ۦ�#�.K#�/����g�iF��Ivy�C6U�l6��O&�D�|��K���?�a���u6Z�q��B�l��a"�]&�?Y�_]���%���ܵ�bB�7qP�7]>5�O+���W&�3#t�3%= ;\L���@F)j�,+b/K��"�aR�5 v���1R�K���[��I�SB��Q�>᧎��*޴��F�'Z��܁ӎ	'�[�>39��ұ���O���]�d!Іޡ-F=���:ax��>�x�����
�irA&���-P��i�b�'���N#^�<���'��'�"�wy�C��(a��+I8����@��c��98�O@ ��J�.x1��'�聛 )��r�!�3� �CM���l�ǐ�(FJ�ϦIq8E�q��'���lٽ&��@ʩg��)R'�'��ɔR�(���'�'�j���͗rh����McԜ��1Oh18�Ȏ�d<b���S:+�Z�Q�8ˍ��?m�'���P�	� �X�s�ύV�ո��O�Ur�cR�'��'
�)w�%��� �'G�90hH$$��S�)ԫe�~Lw�ދ;��#!�i��!��'0��UNxX���5d�5��}�͌�a�d�D�f�D��%E:<O*��S����p	�Ȇ�X�4|��&D��ci�:�$�\�Iş��?�L^�5�h���
�p��B�UY�<��ͺ'��9!����!C�ƊU̓u���'��	,7m�$�۴�?Q�(����҃%F\�p�eG�������?y�H�?1���t_�h�ݴ|CZ}z�glӞ�2�ǥ�05#�$Ą{�4�'ۼ�����+�lI�n�؊o�gNZ�R�ɋw�8U�Ѣ��>����&/8��'���'��(���mV`�c�\?__\��5[�h�I[�S�O��\���&J��pA�aRVZT���'Pj7Mżx��@Z�Q���?�t��60O��Ͷ�[�؀�?����锑TN�d�-4�0�ǁ�W���*��+�L�D�O<��N�6u�} �oH�b()1sA�|�-���;�'�b5�X!�h�W4\��>��L��4�����&Z�M�(��C,�H�����P�+C�5.��g�Ҍ3� �O^�!��'��7-����Y�'Fq\�Zi��gn���k�q̓�?�ϓ_�$�Х�&P���g҉b����I;�HOXL+r�I�K�(�*N,#���*����	ԟ��ɡw+�B�П��Iğ\���߭ "Y+�H=�4&�
,y�� �6@z��Z�Ƒ�n��j�E�@%�F�3?!t�q�@'�,��F�L 1��y� ��7 ����^4{r��PM=�&��	 F�P��!0�%C"$@ %���3شy �� ���'R�'��#��T�
4��A�3l�<���O� d��u��/j�-�ĭ�%+*)Z6��젋������<���j�*ό+&� t��r���h#�?����?���h���O���u>�ʵjɔ<IJ8za�C�k�H�#�+M�h�b���p���e� ����ф�(Q���b$��gs(�KB$L ���⑯��,���jǧ_�$`iS�H�.��h��͒4AQ�D$�Y���/�o���Z�(׎6�\�$�ᦵ�J<����?��r`B=�~!z"ME'l�rFE��yr���D��T�\6%[�,�@)ޘ'�&7��O�ʓ�����?���tl�Ȃ��З`Q$��牖�~�
�a��?)0�_�?���?��b7�2}�g-�N��i�<�ը��/T]�PME�^���.')v�qvc�,]��y4-�C5:����(q$�=��3},ap�'������?a�]����k�ֽ��Q>.
�Y�Jv���I韤�?ͧ��(.�;��D+4��MJ�u��l=����}5��bIB&�`�B�X�/�6-�<iѯ� 	Ǜ�'o2Z>A�7EJ�(8�"�	���j�� 1���)������W��9�+7�>�Y$�;�@Cd���N̖O�y�פ��4hk�"0��YJ�`[ä��E@6�"Ӡ�,�>�iP޿4L�	 �?�Q�#տv8xrѬA?��(��%}�Y��?�ҿi|�7��O�?]X�M`�����2D�4M:��"���4��	8|k�!{a_(sܜ5Ȗ����Ó0���s�ݪ0��	~x.ahW.�GbЅ��֟���=M�8[����	џ��	>�u7��1]� ��T%N�)Qʜ�7�;��c�ܲ{<
o��N���M,�3���!�dLb��ֳ/��A�A��-&��3�i˹F��2�����������Y	D�4L�@$Z!G��iTE�լ�$��IT��Oq��'/:(���xs�a���ƫ4>tKP"O�e��e�J<�|�ԊȬ%ġp������Ӯz�0��@*�"=P@a��(և+dlB��+
ߊ��t�ҁ2p49���դm�NB�I�]Ell��W�2xla*uӶZ�
C�+=�4���FOJm�Rm�"�-B��6C��1���L�Q�'��m�(C�ɐw��YC�@>B��񢃢{]�B�I%N�>8�ǀG�h�(Xd��)C䉗o�*90�� ~����K��B�56��x���f���;�![�1vB�I�
[���Te�!����&�ٱXh�C�	 ��,Q�,����h�Eg�C�ɝm�e��0#@�;�i@�%�!����ȅz��D�!6 �Qn��!��? !f�teЪy ���tM��`�!���3g�(sr�>�l�A,КE�!�$����P&T����)�Kہ�!���)B��u3  �#�����مz!�D��*�������H�ֱ��"Oʇ혼N�`�h�3<%�з"O>�;�c�$q�@�Z���'�P��"O���Dd$#nزR*ɴ76 �6"O�P�t�٘B�}�HS�'��A"O�xk��	M��4G�3?��I�"O�zal݂R����F��4�<"O��D�H���Q�CN�;����"O`��
*P�Ẕ
5��c�"O���.�;��q�8b�@PH5"O(�q�AL�*�D��i!Պ�"L!��^�$Y�Ag�|LX�x��1+����N�	h���hп3Q�e#��&h�&5��n�<A��H
�0=��oJ��
t.U��y��XX�@��L V*���N����Ϗw	Dx�e��5�݈�m�(��xb.F�B��%�_
%�~���U15fbu) B  x�SV燚iQ����:%����{4d(��	$dd��UHE��v�?�! N�"���(�(O�p�2%+#��V� �)&߁bHr	�([��xb3X�B���I�Y�B�|�ӡx?��V̊.P@����J���[3/�``A�{�'=� �����,c u9��74L�� F%n����'�6�|@ň��p�oO>~qp��ÓG���
fP�>E�zf�z��l%�$:��Rmz�㓝P����U�D�>P��'�ضy��8G1G�	ѓA��+	νSG�T�3T0q�xo�@`��D�<'Pm��L
2�J��$H��u�u͖k
$�#�\�����#�T�|�Pl��D.r.�)D=�� �1��d��hQ�ς
6D���	��v�'�-��O��zU�V�ș��2	����\�w�p �e���9��-���@��u�M\H~X*%k^�>�m�'? �B�ݸF�ε��ɀ��0c�-<ʭ+�]9}����I�c��e ńѿ`�$� d�]�c!`a1c͞2�ٹt��`��t8
6P���+�鍽'����$�h{~����~�.A���/w��I�k,����_����;y.��a�?I��p�#�(�v���Q�P��J�G�3+咭z�k�j�t�ӓv�F�5��Tm.8��R:s����L"h�@Q)RV�H3_8s	�  A�X�K�49���l��n:�t�k(��Q��.i߸���nA��hO.}{���o`�M�20���"�fY�KY/yMX�1cC��8)�f�	1���'�1��4ca�T��~BD�B�T��M&�z�Kf�/�?i� N'��D���x��� * 7�N�5����(�,_����'����Tkڻj
�����PN*��d�mn���!8cެණǚ<C�It��AmVMy"���M��9tn����6K�w���BW��h���+s댚).�pGJ4�(l��ɂ?ZR�i�d�7.�B�C�Ɍ=Ә�H��T���$�9;��0㕈ω:e�m��mO;����tƘ�y_I1J�*Ö5��J\7��O�]�$�F��L�>�`�A26���2��W%*����`�)��!a���,�xT��S��y2̂1'pPI��"��JH\ф*����>���T?)��E6�~B ��w��u�F�ݙL��Ć��A�b�O�eh�  v���'\:d!�������$�o�)��X�B��'�	�q	I�m����<9"�6?A��K�`��t	Pk��K���80ε�y�'5���p��m���d%V2cJZ���/y�\�EMR(��<q��U��X�OB�O�3?)�$DP<�Z
̤}P����o����O a�`jj�'x�i;��X1S���y��&v���$��{�}R����	$�J�酷"�R���k�/xubr��O^y)�#�9m1��$��S
w�r��_����,ë=�����.Z�M� 1 eN���G�JyR�t�	�6Qjl0 �d��!��8�O`1�d��� >���8J��<�B�5�1���<�Ӣ{��<�GO�Y��rƍ��7h�a2�0��+�nt��Dc��&�^܋�kܚ .�!!�0Y����ŝX;Ƭf�B8R�@%��O2˓]��q0���0J��DYc?=�� ��	7,v8�JFc����?i���Yp\�a1mK�Ci�#�πv�dʶ��C��!��k�I�0T�(@��69���6U�xa�d�`t��.� ���J��<Q�H�W&J)B[w�K�iG�YC��`�$�=+�$MXM>a�,�k0$LZ��A�vE�1Li�~�iV��<h��B(ݑ]޲�'��КDC��x�6�?8��T'?�	�&\�DGghV�AE#_,��ē�e�/�t�s�n�9��=��pq��X.1���
��:�l,B�S���GH�=_!�����P8d��	�P4@t:�i�?Uv����A+D�tFzb�CZ�:��0ϏJ�' T�}��Ȅc< �D ��0�T�D�|B��pnT��'���"��|��$�:��ң*{ֹʣ	I�J_��*�.��#�.<��o��|����m�Rm��T?M�q'Ն}��T�q����Y�Dh�'8�m*�'ުg�&���M{lܫ��.�#F�DC(�W��CD������^�q���'��'�,�n`S��٨I�$�cF��C<,bnaQ��Ɉ	O$��=�OL�x�e0�nd1`��xkf�pdi�'8��C�^����ˁş�F{ʟ,H�5�N�&c�Q�D�E�N���1�+�I�]��5��4C�j6N	�X�ԟ�d7X��u�0h\
H�>��̊�o7ўܖ'Ƥ���î0O���rc6��c@ �$3R�q��A�G���`�g�F��L0'-�	���r�$����2�JRu��!�h�;b> #�G�'��`��c"�>�3��x.�1����B�l�qO��$�ː4juZ�kU�9T�xb�dT�=\�:�؂	J�-���'<Vd�Gmѭg��iU`����iȅ|zP���@�U�V����+n�]�C������i��h+l�]�'����-ȠXz��2���D�8R̀,(U�-�!��O�r�GU�gM�&?�p�O����g�^��ިH�F�z�t�Eh/�I�:Fu�A`�8���[�㝪$�`c��AA���v$L�rj�/,��;�B�:P�=)���.3�؀��O�����r,��� �ƜP��-<����g�케D吖K�x�_Ob�0vΉ���.b�x�w
��>MRg���5GrА��B} ����ʯ
�V��O8x#�B>l�d��B\hI���O�#P��&*6U�2�(�:"��8�z��FmhI���'q� 񄆂�cr�!T�Ŧ<2X�5��� ����,g\m��+��S�X���<����i89����a���"\�U��PG�*:�F] �.��҄!	�OD��Cm�'D����*,ŏ��߅9bD;���9J9��e��r�
���a�ߒcƴ�Q��ܠ1x��<�"�?w���Rw�	�Y�����˪k�\�3׏I(q��@�-�ퟬ���3}��I�(Al|{�ݟ�ag#�Cr0�+d]�& �:�96�r�8 S�F�Dk�R�F��e)�"΋W���!�+������E8��uH�r&��X5S��ܱ� ��/Х����J#W�C�ON��ps�иug1O�PJ����1�0��@b��p���O�Ή��FϴO�V�f�͈qrF�%�<��M��fU� ލ�=�Oc�0�3�j@jr@��?H�����R�h���b���u��
Y�#čb�jA�~
u���k^�}�B�v�x����.s׶� ���3W���Dɇa���j�(�1O� D��6F���:���$18c�KUnk$i������hP�il~��
��z5��&5��O�j%�׊1��$c���	M'��q�F�?-(1��YV�n�҈y�H0u~�����T�z�� �:��%k��;���OQ��M3�J��(ص�_/<q��3�>I� E&*@BԀ��)��#7�D̓-k��a��U�0�BE��,U/�M5m�6d�'>����Ř7$D$�7FV�+XX�7$�x�^�{���)Q	茓���?V��șF&���4�[,a��:�$i��)�J�Kۨ�R6�'?`��ع��O���)5����I~ʜ$�(��{YD!�<� ��;�D Q P	A	�5��Y�s�đA�@��¶i����OKfv����6
6:M�!�-i���dG^y2e�47�Б���g�׏��v�v�/�|�! �3>� ��Ӈ��6qv�-�|�#�ӟ��g�S"�+�HPs'˒f}ιJ2�M̟��'M��q�l��X�R���1O  �O��<v�z1)���t9h��'t�G��?M�����=͓�\=ه��&`��u��
͞�{e�%,O2h��U��<!��gL:=a�iƞx"6ɚc�OXrZ�O���AƜX+�y����2f�����Y���qi��"�.�nD4@�@�6�R6�ɺ0�#:���?!��@�i��$�&	<�,�ai���0�J?��c��\��!���OD�4��[�6^L�p�-��J���.F�T���Λ)P��d{�KI��?�$�7����'8�Ŋ���������Ժ,ض$
�+O�8| )�\&�dò-Ah�g�?�� ��L̼є�3�$�'�Xd`⍘��?i!���,�`�O�!3��<�WN��Thr���A*��:e�Kq�V ] �?Y �L3l�g�� y���W�ȶR,ja[��'}8 ���9;%��	�u��p%�l)��&}Zc��qȣ)Պ|��%Ib)F�G�x�R��e�	N�4�X��-�ӝH�5x'/W�&�������r�܋H>��˵<�W�������O��L:_c�ꜫ��+oܚ���H�	�<`s��z�@Ty�K�5SH�I���Ӻ�ɤ���xr���r �愗.t=���v�*w��EsG^�Ԡb��+�(���\H�8�M/n>��<�d["V���y�bM"[3*2�G�Qܓ�?��X�`[�H%>�,Ox@b� Ϝ���EԸ(�X�C�#��G�����Y�o�T��F����uY�� ��w���R�B�Pِ�̜i�|��';}�)�y?�N>��M�ƣJ�O_�j���Y��p�IZ�Zb�yB�}R��8&P|+���~�d���ē"0�Ҕ'] o�4Y��S3SҬ*2�|��CSybJR�p	�t��l�L\J��� .�\����2���xk�8O�ʼ�j�8~>�*�K�0F����K�IJ����4!�aZ<]rA��9>P�#Z�d`��L&e��B5����m�R_$�E�<�PT;)�s��U�h�}ӢU+KU�'��'��E��*�?�`l�$�I�Eoو$TC���
%MȧH㜭��}�!�'��,��qމ3�ǦHmX� E�46]*̉��0}B&��U�'CP�)����:Gih��`���D�	��\�C�[S� ?����<ʓÓ��x��.P�2�OVP�F�
hp�J1e�^ܵ`�f��d�$"��7�Ę�qy�"5RM��'7�H�[E��8Q�)KC��.�ʹ��&D�8�ĉ-��tT�|�f���J�B�*�+?O8ܑ�ֹ��D�S��2��9�7�i�d�z���,��XG��'{�p��C�7��Ћ� ��/��@�Tg�b�\ 1A (Cɺ6�F5��̸B�(6a I����?�'�H�P	�-IXB8Z�O�JZp�����N��� -��e����C��-�� M�bq��ۆ,�0�p�!� �A�+'yI�l�'J�!��Ĥ��̻	��юĠ*�=��C�B]GxBkG�/�<1�g����D8Z3B\�d�P�=�>�RVGP�I�ޤi����z�J�Dy�U�9�.�PRO@�	_ޥk����:GJ�ڗ�ӌ�E[W�_'pN���� � �N	;�IM�1�T@c��\}rBȩJb��)Чg���{�E����ڰ~�ӮKLS� !YHժ-���ɲte��0-��A���P�ʐ>��	��ɹ#l d��d�#�F�"я[�rP�6��,���DӊX,�Q�Wڷ3Ǒ�`�@@��
�|���Ζ�0�`�HP���� ?�BX��0��4((
(�wޏ8^��SA�5.�D�@c* 4:g����w�0��+�_�8�(�N�/ J���I�?�FA��F�K687��E��*q��*L��� �ݑA�6��%�D�r�*�9��G#Pa�=Y�m��Y�Z�iw�|�e��*Z�ks�¹^|5 ��3�$!�	Qu��sD�bg�1E�2v �������U��!=��HFN�~jB�cc�ZM�=��kz�ؔ��ᆌ%��)�%�:-��=��>9V�[5�dpy  �2�0ݒ���Y�VI �c��V�.�C�F��!&�<b�;q���#��Cb�8[�j�!�0�S�W��Sbl�i�4�5U
��d���(70�:�N��c`XQ��	�H��v�'y�]�4�[TZ�<8���T��7L��%�<Qa�J>���y�
D��5��i�V׈�H^-i�x��	1ȩ!�,id�ə,��QABI���@b�>f�����\�4u�@A?���4t�DIO!N����g�wx�$��ώ�Q�&����I�\��*��=��KfϏ=u#db?�sv#�$*)-�K�]�d�䈉M~2�6N����P�3[NnE�@-��O^��%��<��h�IY0v�$[�Z���L�JqO�A�,B��Ty���Z���V��芤�����sc��a�� ����SE�E�\S�eR��G��]Q�l�!��	̾|�t=s(O��ѧaL���P�yi�hC�/�'�Py���!��8R�V c��hp���8�y
� �Ӱ��^�,�ʂ�Δ
ٞ��W"O�pk0�F�Ti��	��P����"Op�V蛌)]��j�ᇡFͦy�T"O��wE�,2��͆
�ݛ�"O�d"�$>�L��� ��[%����"Ov5����u�!�c�A/�	��"Obas�؏]��I�cҳ>)>�`�"O��õB�a�\���ɣ8>9��"O�0�S�)x�*�k��Z�!�"ON���#[��,Ж�Q���0��"O��h�%#�=�W*�*��T"O�,��+\$G����F ���htYT"O��yg��Z:�5A�}�\@"O���&%D�\�m���ԃqRUX#"O`YzG���a����	A4ll�B�"O"�Q�#ڞ1���pg�ܡPp��r"O��y4�6l<B�J݅E��x�"O(䌚X�pmp3��3>!�]�"OZQ�%��6{8��G�&�[Q"O8u(���lN����fؑEl�9�"OjaE�N�q���C�F���(�"O���"V�n�t����',)k7"O�D��7s�n!���G�<�R"O����CI�'5�#�'
�0�(��'"O!Ab!�#n=Q��A�t�N��r"O\���C�Y��,g��XP�"O��p4@1��H���,��x"O$x�*�(��+Vr��PS�"O֙���$0�b#W��|�T"O~!H�mP1��	w�3k���7"Ov�� �H�I����k�p�\<��"O�0cO$}�^�:�U�m1����"O0�S%
)JS�񁶣Fr\4bg"O��2Bǎ���i�@�0��`�"O���&@�`�:�[���)E��(�"O�hpfc���R���iO�D?dQ� "O�ɋ�(R�0g��Fj֠B-ҡ�W"OʽB���^�8J�)ծ=�$��"O��bЪ��>w�@ !��'���!R"O��U#Q)ʭ�O?/���Q�"OT8�g͛jT&�Xe�g".ibg"O`�iA�&�$D�A抱'���"O�! sKA�
L"}�'�M�=��L*�"Oz	��.$k����Wy&1��"Oj`�n@,}����b�o�H�'"O��ɇ�ԑ<�έ�V�G�J:���G"OB��B�R���w�>TT}��"O�]2SԿ|ۨ����!$�a"O~}�3�ԫ~2��0c�\�X� "ON���.OF�u�ǌ5fbT���"O�5M̒LaP����r_Ȱ! "OBQ�2U�@���-V��F"Ob���j�a!@�5O�5@�"O���$R6w�0*W'0oѸ�S"O<�k�ゴ���@d,˹�R%�S"O��I��m��.=�b"O�E��K��i6Ya�c�lP���"O�(SϕT�BLj�j5
�"Ot|)����~��T��8�Z�+v"OdX�@@ll�qI������"O��J�1�����6�Hٹ�"O
��0�߽Gz�R4�1s�6j�"OJ��qƎ�8^Ց�f�.u�H���"O��QG��$|�uG��z8�r"O� pxjU���'�M�Ʀ.ku�e�"O� �q�C���Gޑeez��E"O`-@'��T8��ې�
&p@�s"OVD��W�N
��A�<j�~d "O`AQ!�&��\Y Ɛ�w��Qc"OM����*�|�c�gK�8�*-�"O�x�wh�~rA[��W�L�x1�u"O֌g����<�X�ͅ>wbP��"Ot�0A�Ɂ0Ed0HafG�G��p��"O�[�Ɍ�.ۨ\�cW�ha� "O��qGʏ����y�΃:-y�,8�"O�)Cg�b_xER�C��Q�5�"O�� Q.ZK Ȼa���i �(u"ObqF��M� 3���$A���2"O)�,;2&����Ż;
` ��=�S��yb���/�䉙�'�X��hQ����y" w�>�p%_������:�y�B��>�0��t��o�!�p����y�o�Rc����� ���������yh�A� �'���Tli"˃�y� �4a2���x�y`��C��y�)܇$��@�d�ǜm_r]ӰOL��y��5}�� &�
�b��A�Q��y"n�<zaas��9O�j�V��y��P�lZ��J�g��8<��K�B���y"����A4	$}��'d�!
�'����nҬ.�ցX����d�	�'��U5`�*KD�X EѶ�qQ	�'[L!��L�b�\��*Ĵ�	�'��i������J�c3�&ְ�K�'kR)J��[ F�*��qO�wx�a��'�N0�Վ˷2R�qs@�Vr��{�'�d����5U��;pF�!e��˓�(OT��6�Q<־0�G¾CZeB7�	r����@7ܘ��W�z��x֊8D�̡��n|^H� ��:D��~i����J/��ya��u�niĀY'k�!�����-��+gkn�%�́�!���%b��JcQ�a��x�!�ā�;V��O�0H���r�9"!��N'{�f�hVM��5ZQ�1ā�!��A�%1�`TmQ�o!��:�@���!�K�)j��0_���c���!򤗮m����� =qFK=�!��ǌRmz���$Є*�`!��e�E�!�N�]A�)J��4E�� �`/�~S��)�.�]?	�b�po���2I(D��B��@	N(����M�(D�[��:D� �B��T�y9dMV0�����<G{���O89#���2G\K�1���o�!��_���ē�t����<�!�Ė�v\���eQ�l���b�$��v�!��ڸ 6Z�03��%��`�ǍT?�aR�O� 2UEE�	Z�5�f�]#O��Cw"OZ<��^�qg����Ӥ��4"O�t���ܺj���0���n1�"O�1@Gj�<�Ty2��6걊�"Or����05���u��:�@�t"Oܥr�*��/�ѣ 
�Y�,A2�>��"��(�֢z0�W�׭bVH��vD��ğ�;d���e�_�=�8��U��\	���h�@y��
Ф;��ȓ>��qS���B��ВQ����B�ȓq�̡ppFN),�rX�ʚ.Ҭ��S�? ЌA��uxv`ȃH�2t^��ö"O�Eز�� 'R@P9р�?\e"]Q"O�u렅H/&I�Q�c�ڶk=�șf"O��(���[ͦ��͙�} �"O�sŧT&�"MC�Ŋ�6�4[t"O�S2c�I�NEچ[�X��r�"O𺰃��j<�8��A~�@�p�"O��Q�l�������6�,X(6"O>d���qC�1+�Z�U��d�"OV�rBJ!P ���5fb�|�t"O8i8D�:�d��O��ɩt"O��Z2�ӌ]�S�O��p"Of��$�ɸ[R�=p��Ձ��*�"Oj\K1�:� L���?2j(�H"O��q«��g�PAq�d�.et@�#"O��P�cY.$`�Y�[IF�I�P"OT�U

���m�I/� � "O����@ԯ	b�-ң)��	@�"O&q ��Mkz9�C�H"k�����"O�����ei���%�8<�hɇ�|2�|2�'�B�Aa��N�f|�W�*q�p�{�'㌄f��C�L��FǑ����'$B�귢�9Z���)E0�x��Fb($�����P�	���1�8$��&D��X"�8���3��ڱpe(83�&D�4�#M�;U����(�Gn
kg�&D�<Zd,B�����i2�#|O�c�@j�U�7��ě3�YA�,}	Pe-D�sWb��s\и3�,��#"Qym)D��S�ܼT&��#Q6�5Ka�(D�Lc��_�.H#r�D�ݖ\j�)<D�Tjw�ZP��cU��*��UH�'D�hġQ�&v`� #�#N�X �D'D���0iE?w�) @���}���%D�D)��G�>N��eH�7�"���%D��pvC�7D܁��͂�;��<cr�#D�[��S%��@��2$�� 	c+4D����ިT&������:��83�2D�L���ŕ]���	D3	�Vڠ&<D��rW!��KY�-���׸���$�;D���W�:3H� �e�,'��A�
9D�x!��J��t�D�&mp�ذ�/<D��d�GS�`�xP$:mfbE�9D�d�@Aװerx�2�I"S�4Ec�9�O6�%0@�v�ӷ]�����j$p'���D���A��8sR-��O�"x�=D|r�?	M6M�`�Z	"�V��0�6�C䉶R��Bf̩K��#B"ͱ$yz��$?����ƽ1�D.�Ε�B�0;�fC�r��tm��>��r·�JaB�IcE��sO�~����j��Z��C�	 ��X���$^����uG�w�6B�$.�zyy��	@y�dP����pB�W��C���p�z�y�H�pB�ɲKBb3�)|XC�!Ѻ�B�?���i�J����"5��hB���&!w!��}�HйBƉ�IʺX٢�=�!�<V�	(�i�?���q׊6e!�$I�3Ҧظ��#��� ��s�!�P��T���� ��0��/E�!�ą�0�¡nn;Br�$�g"O ��ӨA�<cBD[&bN���r�"O��5K�M��qxV�M`t0�"O���˒�F)��ɖ��.S��UY�"O� ����N/4��v�!�4x "O��hІD�ov�x�g��=zʽ"Ol�q(G2�ũ�f,x��$�"OJLrd�C�b�M�B�ױ�����"O[��J�"FÄ$�_�F��2"O�����2�L���j���B�"O�1��"	��ej�D�:����!"O�	�g��R'�I��!NM����U"O*䣧�]�H��l2v*��e⮜1�"OfQ
�ɏK�t[v'@=��8S"OI�bH"B |�Ǭ�����"O����� l`���[�M��h!"OLaY���3:�
����D�TJ"OH�˗�W,mP��Av!ε���U"O
��q#]���PJ!ڂI��)�"O��"�"��I�X�Xφ�A��Ep3"OM �e�g��ۀ��+��C"OZYY"�P�6T2�X� *�$"OR��g�[R�P4 �PF��$"O�ŁCI�4�!���5w��81"OD�!�f%X�aѱ'C��{c��k�<4%جK�j��@C��n���q�<�Q����X�L�H0r���l�<�W
ֹ0PF � n�,��DB�eVf�<�Q#�
t2h����R���H&̇e�<ug!0�@�"�_����N�F�<a&'�'!�,� I�$T4�2#N�D�<�@l��j~\	 c�>2(��B�^|�<�"#��u�2�&�J�Uw�<�@��#�rQ�&��Ae��Jt�<!��Oz�X���v��4���Mh�<Yg�
k�p(�CΝ� 
�H�P�Ng�<	ԁ7˞za@G),���0&b�<���٤Pi� ���șZ�c`�<a��[}t��	K�;m2�%
�]�<QƁ^���|ґ�$��U��N�<Y�@_�ƪ|8���;ے��ҢYJ�<	$l�JYX1�%'�0^�n%����G�<����3N8\@�&�5b"����<!V*�"�HYr�#�_DhԳ��s�<����
5�9ڔ�� ;��r2�Rt�<� �7X'���hԔM
����-�r�<��N��q���D�Q�p�t�r�<y#�͉p��:#�J�;�|Q��J�<a���t���-Nf�e93j�F�<	�+V�n��% �LB)B蹛Gbg�<��"�l���q��M
��A�_�<y�̈�r�h��lH�v���i�t�<��Bيi�G�H�1U\�# �E�<�e����mW�v��vBB�<�7�+zY�$`�� ]xfpy'!MC�<�C���^����LV�W���p�g[�<	�d�='B�� �Z�C6P��f�M�<	w����i�,�,o�:�Ab%Wr�<�i0z�H,$���J�"�S�<��	ۻ��XM=��E2GX�<���ɜ���b��Z63�Z��FK�V�<���,�|�dhǈ �]����S�<��C«p�i���<x��)����P�<��eA)lLA��۴x�Ř�#_t�<��I�r�U��	'kB}��FW�<����/N��(J��*�$M� ��H�<�5�U�ubp��rg�'.��S�NZ�<���ʴw2ļ�Vl_ Ep�����V�<� �A�b�߉(7�L�~�P��"O�BK *zh�AB߹f��	A"OnU���3�U�����H�"O�����5��p!��9L� ��v"O�TA��5ouR��U� ��"O2E�����x�&`3'Nc)k3��y�R�Bn<(��C A8�!��j��y2/T<<�X�R�(�1�8��!���y���,'\p��ĠKf,� �y���7��p�!�>QNV�kF���y¢��pH* fE�NҺ�2�%�8�y���3Y�h��j�-M���13H��y�D�D���J�����(�y�g�d�柍�zP2���y� �-��ɑU��$	Bw��y�I�6kH��Q3J{���KC!��yb��Ͷ��V �pxI�I��y�$!-�h�X��N�N���"k.�yRON�A��UȘ3GLl!B���yR��-e���$ԻgΝi"/��y���T�rT��i�B3a��yB�I?s�t�I�N	����ŉ�yrL�n4C�!��J���0&���yIDE��A��F7w��su�5�y�I�*r;z,*�+q���q���y"%����"�NM"@��yYt,�yr�ӕ}�Y!��2=����T�Ɔ�yB*��e�Ժ�b�$64bIi4�X��y",Ʈx@����'`f00�g�;�y��ـo�
x�+nw��A��
4�y�e���-]�l ��G���y�g��3A�\��hQ�A��yaT%��i���k��hԩ[�yr.��5��uOܶ��qR7�X�y���86�4����<��X���'�yB�x�TYZ05eVP������y��	Wv�ŋ�^����S7�y��K�D� ���	�]�M�D\��y�TB{��:š�O4,m��i��y��ّ?�� �U���:Q��b&���y�-��M0�вV�Ί1�������y"��>۬)8C�,w�X���y�"Y:.�|��o)/��&�L��yRh	9I(̴�	°-B���U�J0�y�"�.Q���o;\�D,�K�y��U5SB��H�dt��2��y�5��p�sn�[u�p�ZI9�B�ɖ7��}�g�R�r�PA�sB�8��B��
��e���(p�z������{7~B��
G�`�ׇ��j@r#���-�BB�I�x{�tK�
�R�v� ��;&^4B��
{O�U�`��dx�I;[�؅ȓ1�\I���.9��E��- �ҍ���`�eS-O @�v�F�E��ȓ[��a�	A�o�CP#l_�4��r����s~������Mw$��17feS�mٕcx0X�O�!ИԆȓVC> ٓ�ۑBz�4{�
��'T��6\�q]�68&�E&�(:B�I*r)��x�O3�Z�@�ǖ�tfB�	v�(�Xg�K�7�w̒��NB䉎e���X��'����E͕�`_�B�ɤeCj����;Q��%����
B�	((mm#� ˃Y�`@�h@89�B�)� L4)��\Jz ����~[Lث�"O��['A�b8C�Yh���B"O~P��@�<U9����N*5eN���"O��Q�F\�n�l�)%圓(�����"OL��Ɯ�:�Hf#ŭc��h�"Ov��&g��rΎ�x#�=!w:98�"O4h�'�C�\B�Q��A�
nd� 0�"Ox:����\�:��ȍ'S�UV"OtI�/�	NKX���"�,^�x�"O���'G�	
���3 O�`xR"Oj\qA�H&'n� �$����&"O ���}D�J��S7���"O���,�YI����VM��P��"O�D�1�Y7SVhFQ5@���8&"O|Qɇ�*H۠8	Щ_E�"OfL�T]h�E���+;�I��"O���dE�Mx��a��Ͼ;6�(c"OJL�g(�rg����8u͠P	�"O�[�π0$���FA�Q�B�a"O�1Ce�+�U�J�A���q�<!6\�Z��4��̄�\d�"k�<�j�*B�)*����X�j�<I���g��9$G��G6�����j�<`�RU�|U���SvF�y��M�<A�"3c�^u���߈h⑱� ��<�@J�6dA4Ɍ"q�@)A �S�<���Ǵȩ�d�=p%iyul�X�<�ЏB9N��Y��P0��$�R�<�b���={p�;m�^�Q�.�u�<�5c�O�!h�$�4\l�3�g�o�<��ɱB��8�VJ�2~�xH��	VR�<iRri6���MGd�V�2b@KF�<���+u�j4S�lH��B�CJ�<1�-�y,UPS"�{����LDF�<�劓�e����A�0.O��r&�LV�<a���z�i�&n�)	�^4bf�NI�<�EMA�`0ZË��Fb$�����A�<AQ��bā"���ȜS�h�z�<ђI�}eޱ���ܿ����GGq�<��).F4�`� кT�� �o�o�<	'���nd(�A�����`�i�<���ˁ&�p�CVl��b?R�  ��a�<9a�ؤ '���`�T`�t�Wla�<��G�;kpR����1ol�k�jH�<��NF��ɀ���|������D�<9u�x���C#C�u�$�{����'H�D�mn�i�f��8��qJO�T�!�*
�����!k���Z�(�!�#tHP��-w��y��cE�>�!�dJ���%��3�T�PbЃ;�!���%��}�Ho�Zqɦ��k�!�d��b��I�!g��58�+�q�!�DĊt��ȩ�hT:kDZ8#t
Ļid�y�|"<O��!��
�d[���"N����"O��c� Z)N625��Q1o��f"O�0�K�s�\-��)-�N�YS"O��8#� ;dj�s�'R�b�Z�A�"Ox�XEjO�#*ASW� B}j��%"O�@3c�x1�Ti�ƕ�BF-A""O��xGQ6P2x�)�иC�4i���'���H��Y�^S
���+�9f��rn3D��I�,S9i ���I�J��{��#D�0J��\M�j�F��Ɣ`��!D�h���[�mx<}0b�['�z�w/ D�� :!��C�R�}{FX8G��y�"O��2���P��3BI���"O
YQvl�5��"vVp�m�d�|���!�'*Wܨ��!ҥ^ `_)^��A`V��G{��I�9 @by�R%N+;_t��dD�/e!�޷7]��Ap��![|Z�ŋ	F!�@�J�5����V/Ш����|0!�$�x��"��h�~t�b�G�l�!��W�ܠc�����P���'k�!���t
p��cԇ9(V�1gˋ10�џxG�T��?��EA�m�4S���W��7�?YK>!�����I;s-@8C�NȌqL�9ff@�JyXB�I�D�N�*�҆vu@E���PJ,B�ɴ���3g�N�3�.qB���� B�9W���/ A)-�f`�t&B䉛[r��X�J���2=-�B�I"��|s �̖yB�p���&���O��'?��%*N�X����-V�<:7�
H�<�/�' zp��ϫ5� �ф�E�<!0��
��S`�lH6��ĜE�<���?lM�͙��V�d%�V^Y�<�����?����֯�->�J��BnY�<p�;�6�@$D�Bz��iQ�S�<�sGN4"dr4z�NJ%;�R$�%aAP��p|r# ��0.�R���o�L�pM�O�<��$V�$t��̎���6m�N�<y�#�	-�-X�J�!T�j4�1#�I�<���X�#��O�����D�E�<	Ჰ�&�]�r�9�EiD:EҌU��EL8�X���(7φI� ��r�,��ȓ\�`�@�%r��)W�ǻ��QD��,p(��(����U�4�Z�$jVB�lj�$�'r��H���2sTB�!w �C���M��\96M�(XTB�I��I���)B)�|bv�6:��B�C媝ZD>ܴ�G�̞5&�B��X^QС��p�~0��ȆUU�B�X�l�I4�F)��ͪ�@G�\��B�IAfb���)���x�Vl
<c{"B��5Y��]3O�0n���3P*�DB䉴2��5�$��X<��DG�C�ɏL�Q 5�1W8(9S��� _bB�	�h	`����ۮl�R])2K�J�ZB�z���clH+��"��z��B�I�T����
L�����a���e�B�� ܌���)?� ��`�OE�B��/ �Z%��<I��#J°#̒B��>�:� �#�:���@!eŵ2�,B�I�>�,����5QL����P�&B�	���H{����9�(q)�/ ��C�ɭ!x����
6We�S���H�$C�I�2�&�����R�3wf�����O.�m����ɣu풉Iԃ�� �&0;a$,D� ���[�s R-�����d4
�RVl)D����H$���y���� 1�5,B!�$�/��i5��uk(��hO�!�$� `��U�UU:=@g�P�!�$G/,��ȹ틂wN�q)��7C!���J|����.��ya�ܬ%�{�Y�D�P�=�U�ԙp�|x��(p�hD��u��y��h\ya�\P�(F"R*�L�ȓ�ȴ�U�n)�o�K�؄ȓ�i�&ˉ0��2�+�$����^����N�		���k6���S�? XA"�r�e
�	4 3��B�"O���U.G/6]|$'��s���0�'�r�'��$FRt�ѷe�Uؕ��&L!�DQ�2#PH����t!�������%H!�d�4~蒐�V�ΌM��Y�Z!���9��� �!64�[��|9!򤂖^��d�Qhɑ-�r [��	�M-!�$۹(9�0 �g�30�0�#�r/!�d9%�ԉP�ɢ4ʆ� ⪂�*!�D��R��q��h�(� 	�=a�'_a|�#e��ɇ�x&T��hշ�y�� A�P�B%�x���`�c^=�yB��6�I#�Mߍn��T�g�F��yb��g�"d:��4g�-�l���yrA�pȴ����l���:�	�1�y���np(w(���7f��y�@���5����)�VZWkC��y��9
�Dm�F����j�*�y�ρ�y�m)�a�aj� lٌ�y�,�2W����� �vx��pa	҈�y"�M�gӪ�XQ�X n��dI ����y"#����'��"��y���ě�y�-�$y��@��I��:5���ɖ�y��М�d�PC��V���nK��y�(÷A��iX�&Ƿ �.�@Vn��yE��N9�*��H�A��e��(�y�n5z�&�ۭ1�A�����y�o�\XN�3H-	4�u��y򄆨�L@�wE6�D�۔ED��y��e��H��3r�!��
�yr�B�����&�N4�����y�.5fB]�0��"h�$x�Jƫ�y�L8dk*<���^�.E��E]�yrNݣ���pQ+��Wc�Lڼ�y2�
0,�F�{�*S��P(�����y�����}b7H�4z�R-�?�yBI�H��\�&N74İ���_�y��jdp	�F����BG�>�y��Gp� ���	�Z�dL��yR�o�@�� I2Vi�+ј�y�^N�Ų�#�;��0�"��y�m �!��Bd��
�x�;� S�y�J*(/�`h�(0U�Mk�'>�y�Ɗ�԰b3CM	LK|Y��ɒ�yH"v 9��%�J���R����y2��&\5(���Þ<A�9�ؔ�y������t�,D�P�I��y��7e(�B��4�(<Z0����yb��jR��b�g!z��Q�Fj��y��PH�{@iJ ����j
��yB���(�L�k ��d� h�&��y2G��/C��٣��W�h��0���y¨B�h�Tdҳ��J�$r�IV�y�l��)�d�4/�=�}�Di�7�y"�Z4� ����� /���3D�ޙ�yr�	�B�i�+\�][SL^�ybhz4T{�`�9��ZT��;�y2.ؓQ����i�>Ipt[V��y�!�{Ё�Ql��n�������y�.ҡn���r�.Ϯu��yu��)�y��<7�L��4@tF8�$���y�Ə07W���QHF-z��AQ�	Y0�y��a{d�-�p� ���"Ca���
�'48iӁ� v߸����=)��8x��� ΕQp��HZd�S-ͼ�:m'"O�1����R�f��Ɗ��J9"&�'��<��`�3z��P��J�8��ȡm.D�̐Ţ��{��؀��
IA�`�*D�<Q�&��4�z�����!2f���e�)D��V�;�8��D>X�	�`L*D���I���4I���Ëʽ�vB)D�di��քe���� 
�(j�Q��&D��y���5F���i��@ΐ�q��)D��%E{�!xeA@\7��QB�(D��i�a\,j �r�H.l�.9�3D�ģaΝ�wb�i��;����1D���1�PO�=B�oG���o#D�\H���?���k!ş%8�e�d&&D���K����o�9�i.	/h)!�Dգ����')C0�0H��D�?�!���-s�$�F�V�Ya�L�*(9!򄛑ERAb@KC�w�l�A%�A�(!��M�6�X!�#ǐ�����x�!�$�!0��LC��S��|A	S����!�q�j@�%<�dzs���=dT�"O4�d�DBj���M�L�6\z�"Oް(w*S7�]�עE�#�i@"Oĉ:F,^����a�Aj�Qr"O�|K��#ͤ�+4�ݧƄ�"O=ѡ+Ř�UC��+��Mb "O�ܒ��u��LQt�֬w��k�"O����-�N� �3Ԃ�>R�>�*p"O��a���KBI����.�Ԡ��"O� �d·8P�I��86�xH("Ol�1�� )�p IQ�B���N�%i!�Dtc<���� ��]B�H�!�$ hnQ�5"
�$�����I�"7J!�D_������.���d�
i!�ĕ#w��Y'�6j�L=�'�Z<eD!��]*y����
E�0y�S�#!�D)iP4J7�K���1��(!�ЀT�`�R���H�XE�`� #M!�d��p�i�u�Jkb��m��B�!�$Y8>�n��H.gS�3m�!��:��u�Wi7<1u��7�!�;"+�a����s�,٣l��8�!�Խ8��i`b��4YG��j!���OZ40���\& ZV�6xd!�Ěuu�m1���Q�s���.�!��,��%�Z9��MQ�DV.!�!�H"
�^���gD�8��"A�̑/�!��l����r+�9ӎ�qa��m�!�d�7XG�IQSI�\�l�PG*�!�Z�x,���G�C <Hj�O�?�!�N<:�q�,]V��UMԵw�!�D�;&��2��$O�6���*W�.-!��Q	6�����K�xJ��]:�!�$�-T�0�L<��t��!�^�!�$�N�� �q��x��`ė<�!��C�!y&��T˚h0���!�D��H�,L��i��+�H��W7/�!���o���IN�,Oƥ���V<!�Խ?���[p�D*}�^��	7�O��=��̄y�l�������.Z�b`�"Oz������h�0����6�>ᡳ"O��@BE��ڌ�2��*B���C"O ����n&��r�	��"�7"O �"cM.d0��&Ã��r�*�"O� �\�B-�;7�tY�+Y�M��Dit"Ox�
$>���x*B]B4���'��H���I�t1�!͵1��f�6D�J�X(Y�:٘B�=<��+gE2D�t�w����9�	���P"�3D�������w���+Se�Y��D�1D���6��4aڇ�W=v}��{�/D�T3ǈb����ٟv��XĊ)D��)���"��s/�-� B(D�� ֍������B�Hw��YQ(D�Ԛ� I*-�"t��+��%D��z�� �j����L6ao�@�"D�� ���5GJ���I0�z�ч�!D��q��I
�ʂ�ҁl��5�!D���f��(����'N�(?�rɣ�#>D�����K"`칀���=k:�95C<ړ�0|:�w�y��_Z�&��i�j�<1�f��T*�iP�Y�3N��90"�f�<AĤțR������tL �A�X�<�1�0��%	�E@�!Hx ��)�Z�<��"-V�� z
E������S�<��ȓ�F�6��d!˸?�D�yf��f�<ɱ�a䢝`��1"�IFNe�<!� �	�1!@�X(
�>m�`d�<1��Z5��` +�d��ؠ�yi��!�z(g�ьm��$R 钃�y2@I�b����"��g��ɸ ���y�\.=���
 �HHM��yf���yB%bg�ݣ��L!	?��a�Ί��y���7Ϛy����3�TK���y�E��h�@S-A�4���ŭ�y2�R�T` ����-;=ډ�1�\)�y��C.����E��$�}�@CQ��y�C
Y�֕�3@6�ԁC�lV(�y���|ި��Sm�d�4)z'���y��02����Xа��fhݻ�y��O�����H-`�W�$���?y��?)��?�����1,�I�	&b{���S�,^�!�	�_�HB�B�k@����R�^!�M�ll�!J�(�^�8MS3HZ�!�d΂:"��d��+"Ũ�b�'/�!�0Y1�@���ɾg���s�nәl�!�ċ�������BV0Qi#��:&�!�dȴA��`P��%cO�u�j��g��'Zb�'�r�'dR�'���>�����6Nz��� � ~�nC�ɮm��<BD��:��"���=$"B��$��0�厘�(�#���C�ɺ3�*��7E3��]6��o��C�"���C�dH-G�UR#m�S��C��;2Q@�k�����ix ,V	=���d�4��5�ScŦu��*JفJ��'���'���'��'��!}fT�
���-,����g��4'�C��".��@����6���9&b��\�C�,SĖ�r/�0�J<�RBZ�9�xB��8Bw�8��L�i.���t��X&RB��=tÌQӧ�N�w��L�)�06dC�Ɇ��:�m��Y�I��h�.I�0C�	)9t�Wfݶ���S�\ BdC��)y�H��+ڑ7�@�!j�Xl�B�3
�\D��N_,W�X��&\юC�ɯh�*�kA���,FÜ�S�"Oh"����P��(V)�{�:m��"OFq��+�W�4
�킫XȖ�"OF�k���P�T`�S//N���w"O� (|���F[~�����إ�R"OHQ9��E]"E�GE�v�hX*&"O.Q�s+�rU�U��Tv���""O^���d�=��� �J�k���s�"O�ڒ�Ѡl􊍘ΈB�L0�"O��)�?����H�����"Or	A5�EUc���_�K�&Q��"Od�R��TxZ�0�����ʠ���7�S�I�e�J��4�Z:h9�`��K^�'�!�cy�M�ĭ���J6/p!�ڬ7�����D�	���b�� +7!�dh�!p�Z"c����ӈ�!�ʐ
z�����E,�����K�!�D�/A����Ŕ�c%*�Ya�U�L�!��գ�8q���<<p;��	�g�!�d��Q��j0�ҳ������!��Z�M�N����_/Ja�b�ֽgr!�[�js.�)6������90hʀ�!�DWH��(�� ���@uf�|�!�ŌVh��R�)x�ġp�Ѽl�!�	*h��Q�r�÷|iP��7���!�%j���kqa�
q��J$E�!��A0T@ &d�H��Q��B2_�!��	ICl�"�`��"TڕXEM���!�$B�4�:�OL�AN��R.~�!��ۈVB��KU���];.��&؇�!���@���Sԏ��)���f&W�~!�DY3DӪ���g��!Z��`f��!�T���;�������6F�
�!�D��X&|��I%���B&���^U!�Ix~���2#ŌIrl�rk�8�!�X��	�a��d�<��é>E�!�>SD�){�e�?d��Z�Z�!�D�^[����k�)"S\�!g�L�U�!���6$ ���/c��l9^�PC䉌/
:��!��d�'/�r�B�	;J��5XG�Q�OD5�����B�	
(��!�$6����B�*
�B�DNa2���D�BA��[�{ʊC䉧v�aI�A�?�0����	S8�B�	x0j��blD���f�ׂ0�B�	"h���`�ݮ�:uMW"88B�I�@���2!�G9f��Dx�)��iZJC�a�L�+%��(�ZJ�/�*�$C�	�$}.R���P,t��7��=QL�B�ɢsH�XJ��S;n_x�kζB�6����瑿tq@y�%M��vB�I��JYb 6Gʈ��+�*�VB�I�.�~�b-H���xٵ�ԑc~C䉏v��Q�	G+n^�����PhC�	;.����B� ?����F��ZC�I8@j\��DL o�T���f�t�B�6P�D2Y��hH�vD�gHDC�	N�XLJŁY1(��%!HL�$C�� 5�rT,�Y�(UX@�G�JC�\��ܸ�-	�3t(`����p�:C�ɘ] �Y�؝��Ŭ��mPlC�ɗ�������4\��YK{JC��i��e�g�ǝO�R�H1��Z C�	��H�W�CRtJի��S�R��B�	�o�E"K[=43b�B/	��B�	-dfr�J�KР{*<q�Q��;B�B�	?<`���T�
�E �L��@X;v�B䉅og��I�k�a�Θsk��n��C�)� ��صĜ�5�J]�Q�� @�!�F"O5k�gK��xz",� ~�>e�E"O�QF����<{��2"��� ""O~0�r�Q#�И�Lݑ}�lU;G"O�p�-��)��i3�E7(h��"O�!$�\J��$c �w��J"OF%�d�6u��dct�Q�B�^���"O4l�@��E��dCF��(�
1�"O �4%̲'��S$L�/Ԇ`�a"Oԑ�6��(�	�A<�n�V"O�l`riBP��`ȓ*��c6x��"O\�A�F� T3	[�hYz�[1"O���f[�}�@�[�C�d�6��v"O�!���/$�HFݠp�<�"OhAsuL�q( ̪ eɨ1�r@"O�	�E�(I�&dk��	B��]�"OtT�G_"C�U`�D�h��"O��a%#��k�֩�gޙV�@%�G"O٪�g74<���E�?�:�i�"O�łG��iuC$�sS��b�"O���e]�.�\�h[S�T�E"O�d����9\���uJ�M �"O$�!FL�7:�x��`�:A����"O|��a�߁Ä��̊�p:JP�"O���'�#-��e�3]	1h}��"O��R�(�2BcХI� �R���:�"OԠ��*З_� �'�L�%���9�"O��Z��X56���(�?}xuI�"OD�󇡃�$R�eXvʏ~��D"O��h�	�R�2s��2lB�`"Oȱy�
�>�T��Y�2cDt� "O�ɹ��*�a�,�>IƼ�!"O�e�r���� ���UM[�s�"O�d��	6n)R9�V�]�aN(�A�"Ox,Y$N}T���n�d��sF"OҨ��A?�Fq�����$O
$�w"OPU+/HÉ��� 1C�dAQ�"O�``��/��zՌV� t�K"O∃∍�Z�Zt�-w���"O���E#D9��lk�o�zg��ò"OTѣ�K��p�Pe��ӭk}�ـ3"OH�*t��%c���kaO_�$rܭ+E"O�u``O�&:F�;a���;d�
�"OPm�f�߷p#�Ը% 2�=!�"OZ�"���RA(�w�T	z��]�u"O�8f��+�H��"�Y�l�E��"O��#���m��J1BƇq�"�+�"O(�b3��u�F�0VA�;"��"O ��%%�f�P�R@I4 o���"O`,a�d��:m�Q��^�~h� ��"OD��蛞c��3p%� s`jqc@"O�|Q�nQ-bJ8˳$�0P8�aR"O�q!���<L~l#Fcκ	~�*W"O�#6�EVT0���ʂH�F%[p"OƵ�U��	Kx��a'�p�N�Z�"OAr�� UjD��$/�@$j`"O�,����vRXLAgC]�xD�b"OƜU�/����3ɒ:S��07"O ����ձE/��
���u䪌�p"O��2Ƙ�iX�Q���7�&�J "O�5S�響�X�R� nf�$"OP�獾,\��h�CU�CV�̱�"O����;%�����'Νp���i�"O8���߃9��Q�B�Й<�����"O� �x��ϳ:gB	8!%,qA�"OJ%2'�שx�2����d���A"O\���>^L��B$�ls�,�!"O�d ؅#U�h����.mW��z�"O��(�F�	,�v�I�#�.�����'�	�wO�./��[B
"M����'�
̑�Y&3�Δ#�H��hR�'�p�feF�!��D�5����5I�'�fM[t
�B� ˃:���'��`�[�qr� 5�M�
T��'cF��@���!g��J�h�}�%��'G�(�P�X~��`�V�r-z�
�'4�p�bnQ9z�6r �W�p���j�'4�9�s�Z~%6�����i�v�C�'9��	5��U�29��K�a��d
�'qm��8�$m�!M�oєLa�'(d;�(֜����aЇa�
1�ʓo���l_�YGLm`��o�a��v�d��SH�Kwԅ��k�
�,1��8l���A�-~��:�!T�d"��ȓk4��-�c����ah��_����]rjѪ�땋=�q���ܾY�ȓ2�d覩�E��Ƭ$W2f$��K�l)��ȍ�t5�aȎ(�6���J.�]a$Ė[>@L��ʋ|��,����"�v*�+�ȕ�=�x��zV�3�,Ѫ�G�@��ڐ"O ���n��|qn=3b�._,��zU"O��2�5��U��F�2-��"O�\��@�,�r��صv�0$�q"O��嫙�G��,҂�H�f�0�5"O�Uӵo�����SkS�Y�wG\!�	�K�$�q $L~�nau��1�!�$��A��<A'�ջk~>pb	�7[�!�DI���ЀwL��,�vm��g�+n�!���C�ʱ�4M]��uK�(�? !�D�B&��a5�}��9����C!�S�8��hq���d��3V^!�����4A�i�v�!�c�	>!�ܚlD*&/�:r��Z e�H!�ج!nf����Wf0l2���Ku!�?.[t��s�РO�x	�0�
M^!��Ruli�4�[G����K��[�!��?��9EJ�9�^�STM���!��o�F�+ы� ��r%͞1�!���/�Tuk�Mf�@�	w��]w!�d7��D	-��g�E3��Vc!򄙙j�m��+�BA�iC�R5/�!�$lp�z�E�2a�I���!�B��"��٩iv���Ň�!�D�]����S$9����^�T�!�/tM� }k`��B���
�!�DL�*R�bc,�r�6%Z"B�N�!�d�6�`���Y��� 2+L�!�D�}��Qb�g�!���Ȃ"�!�$�1tr$� ��� N���w/��)�!�a��	;7+�5w	ళ��_�A�!��.�<��=3�`�*��N!�ă|3V��A��'�d�����lR���%kZԊ�a�3]F��Y��y�T2Eyp<�
�I9D��U�H��yB��2fx�(�f�Fn����]��y�eO�2)��ڨ��%�%%S$�yB�L����ƥ

`�Q�Mʘ�y
� L���#e8�=i��5V~<�x�"O����	]:_�&��4m����"O*��VBI*y올*�@�q��j�'l�L�D*��D|���3�0UQ�'���K6��%��XR̭'vt9
�'N@Z�/N�Ud�m3��(.a���
�'�A���N�p��K�1?z% �'��E��oZe,ܩ��#F|����'4 �!�(ZR��b#[ys8��'9I�N�qx��bfԤsc��8�'f���u�^�;J~T�@E�~p�q��'�*�p� ��XXc��W'r��x��'H,y�D�لeJtrI��q��m{
�'?��B��,rBQI&C�c�$q��'�Dt	ӆ�K��qE�ю^��xI�'����ŉ��5j��+���$�
z�'�= �D�bҍ�!%ْX �'k,�Yu,Q������@O�6 �;�'��@Q�F9]�L�Gf�(��C�'��ҡ��t�,�sǣ�7����'���Ô�[�jA
4J��$& H�'"��`��~�}��Lp�x�'1�i���h����ՇF$)�(�k�'
�Y��JG�9:m�4��+���'��-@gD�dJ�D��"*��ub�'�P��ϤʈT�@o�2h0�'��и����qZ�̫�'���'mX+�"�>�(��3D����@ċ-<h�B)��l�
��?D��S")�NY9䀗Z<��Y&* D���r��%)��!	�;'�a��(D�y�(J�@�ZH�d�2B��8E�3D��ק�u�$�Fh�.̦p�"�/D� 2·�F�MX�h}�|(�/D�`01��,6�ȁ�GFi�4*O@�;FS$����S?z��#"O �����<
�F��8��"O�}�҅���a6�1)H�qr"O��4��x�j���)e��#D"Oa��&Ҁ��d�p4L+V��"O�������М�F!�	p~�x�"Op���I�u��Aӏ�}�֠	U"O:Ū�!��F`T��^j�"O6��#�	�� �<'��s�"OZ�S��Ѣl4̋�(���V"Ol| �c[�U��H�lP=���5"Oz�Y%��<�h,2dkn��xZ$"O�q�ڕ4<�q[1��dM<���"OX�GN��7}��鑖dD��"OxQ02��5d&$Y5�߰8d$��u"O���Ӫ��СLL9IbBQS�"O�Cu�U3��*�K�<Td��@"Oȸ�BG=�z�Z�ə�d�8�"O�(�vKŜRW� ҡ�[���e"O�e�D��;�J�����g����T"O$���J?Ɍ���38:$S�"OhU+��-su`�+����'���"O�E�t.Ԥȼ�
��F
i���"O�5�"��3(E�y�g�� �x}�q"O@`�aDT�&z>聕#�<�p���"O,�A��$v�T+�<��+"O���kɢM���� d�SG֤�""OTq��aZ�]��!�E"1+�X�"Olx�'G�+�|H{Ѡ%G��U��"O� <�I�M
;b]K% �o�i��"OСSg&�b���@��	�kb6���"O�]�螦Oe��q�GѯQR9C4"O.�x�hˮ[�f��f&��a�*�4"O���U.�&���S�d�|�<��"O�xp���#J����ˬd�P��"Ozi`g�E��|�T^~$�8�"Oڝ!���5&��rh =>�4u"O�E�e�A����7͛`��H+�"O���rC��`���T�;���3�"O
�U%�%#�Q�Qc��f,<��"OP%i�㞱?q�IӣO'Jn�C�"OL�zFB�:esp�sV�-.��x�"O��b���!���$�X���"OF%
�B 
��YH�`�wr̊W"Od1B�^��m
g��=vdL��"O*@���!R����M�R���""O��ʗ�K�Dx�Y�զ�:w�r��"O^�A�
&zV �8��&x�ua�"Oe�Fk�'e�h��5-U�Z!�"O�5����t�6TX��=S�}��"OҸbD܁n��0��x\���"O���'&ĳt��x$ƚ� [r$��"O(l�u˗�QT0�eK�gU(i�"O�P���̣W��)2��%yS��8A"O^����ɏn�ֵ�L
k�<�8"Oޱy!$��0�X� ��p��ic�"O���٢pv��{/� ;�:��5"O1����]��L��oK�~���g"Ott1/�*:�ri��g�<��"OMRu��(6*AH�^i����"O�X*�N�"VW~�"MB>�-IP"O^�P��́tdh����.���X�"O`�H�.J�s�HY�S]��u�V"O���r��G��s`I^�_���� "O
��"NV��%r��οm�Ġ��"O�yz3�
g��(�B�}|��`"Ofݲb�]&+0	���53�Z�q#"O��Hw��/�X���C�"O�r-V.ݎ�b�DҨb���A�"O�-Q6
�0��TC�#yT�3�"O6Y3P��X�4��a�b��l��"O ��e��~��5���� ��8w"OL��a��E��xk�OK� v����"O�.����i�	D�R+5�!�DM�O�HB1ѪB�:M�Sk��R�!�d؍>@�@��k�STmb�G�5v!�?f%8�Pb뜌p��m��E��=^!�$F`���,ӈ9�H|�Լ&U!򄆕$:�SDJ�r"�Z���7t!�d�LA����EJ����,PO`!�d�PւXr���0-�,S�%��cn!��	;=0�{�g�e)��bU��H_!�$� ���� ��E�M*��@0!����´y7ꑅw���{V�[y!�$a5�M�E�ư^��m�E��5px!��U�������Ksh��h�B!�d�V]�)ɒ!ȚcnĨkDG��a"!��dD ���t@��j$'^	:!��Gb����G��8�P��+
 M�!�d�iCflZ��:���	����e-!�D��++(Ы��9��໐�66r!���0�L��%Ë+x�\�Qm�|n!�է;�`T���	�1t��#BK�3Vc!�� �٩��B�/z�q�q�ȷ ӊ��`"O��ej�:�A� �� qX�Ђ"O�E���
�}�*�B�\\�]�t"Ox��� �b֮�a򢕢v�<�r"O"�� .�2%_��ē/N��sV"O,m 1�18D(1�4�\�~��XP�"O��0���d�ֹ8���x�M1a"O�X𲤋*LrL��� �H�2\��"O�- WK��T����S49"��X%"O@d@�@A�X�R�k$*���C"Ob�0 :���2/�� "O<UE��37�	PwJ�18�	� "O�p���$< f4T�4#�.���"O�8�u��</j�uCC�$���G"O�)�g��i��:%�0^���sp"O@�#���.$-+�i���ڵ"OXk��2Z �8�ЎJ'���t"Oj$���;,����O�;Gq��g"O�M�Z�`�B�!{�
�P3��y2��R��9��f�$����^��y2+G�o��hdBR�eZb��'�y�i����YQPCµsс���y"����Hj'�0Kg��P�W��y��+Ò�q�O2k�6��n�!��0`�,S�AB;hk���4g�!�$�XU���5(�=qc�h�3ł�6�!��\�} hk�V�<`��E�P�r�!�$�T�p����;Uq�*����!�Ă�Y��9S%�;3	���H�D�!���H�Vd)3�ه�>���FD2q�!�ěl�ur��U��H1�& �%�!�J�A<��:���/+̊	�&M�j�!�5
�DT0���:�N�(�ą�3�!�� z}>��ơL�!�9@��۪j�!�$�B�I[h̔8�����a��Pd!�DS�f,9���B$4;fI�3G�q�!��� t�s��$Rl�V�G�T�!�d��p��;�f��l+w�]�G�!�˒�b�i���I�m��	C
=�!�K�J�����8NJ��	đt�!�d�= ˗lI B.2��� y!��/�FaFdU�o� ��B��!�D�.wj��`C[�{��@ŏ�%[�!�R	[���$��3@H-	"%?i�!���n�� ��n��K����C-Z�!��U�ZV��ę�%��q�7��>�!��3=���EF�o��q!7+�!��U���M�%n(N|�r�J0K�!�DϺ�֜j��!}�8�@��?Uy!����0��	����cK��5^!�dL�@TD�ELlݖ��	�� C!��ϓ}B�]���+`��A):$!�k�nd;���C �	qVx!��X$n���9���?\�yg���^_!��4���p�Q�*�3m�� U!��20�,5�!�߶?�@<0"�ZI!�I�hB��!Hk@d �r�oH!�DS�8V�D��!K�U���C�i�FH!�P1F� unL�$(N����8o�!��[�O�X�@� N`�M�H�!��T��@�1E�^z1���	#!�$�H'V�˂�V9@jL`�Cf�Bg!�DB-#�����Ə+x`�]�#ѱDT!�$�5��y�C��f�as��N1dS!�� ��� ��G7~!��c�+>��8 "O(�"�X-���7��!�P]�"O��F<Zm��p�
�:p
�Q�"O8}R��_�'\���Ë1``�,�"O��:5�L?4�]P��U��`<��"O�L�6�:-R�} ��H�� ���"OPغ�
C5S���B�;?�}�"O(-$HC�`��Ìς�x��"O��`�b�䁢Ǆ{A�ĺE"O,�����;dfX9a�Ě0)y�"O�wC�4p��%٣HO�s"
-X�"O�;Չ�8?(0�����s��s"Op`� ˉi���`R�ak6z�"O^;f�_��Ѳ� ^ Y����"OvX�	ځs-JMk���x�|�"O��3���d���@ �~��%i�"O��ȇO��gN��*`�����1"O@�Y �	n�VNN�K권� �'tBGy�"�Ce1WedI0�˖�y���q��A��H�\�NE���yB���[�*]� J¥`�f�;`&���yS�d> Ze�	31J �g�ƍ�y���+� iU�
�f0X@��b�,�y��+X�����a2���J�yb�V/밬��Ҏ$�̵����'�y�ϰ:�4yɔo�"�ppKwcP$�y�I���!��֛!F��Y�(�y�5^��u�@8Di����M��'rȍsE�	:���`a�6�h�C	��~bM��u�� !�F��X+tJʦ�y"j�|O"���)C(n��8b �� ��O��F�4�ʽB����P	I��[�G�y��`�?�S�J��Q(�a���i[v+�x?��Z�L%����
�V9Ej�+
l$����
1x�0�O�<)�����W�^�٠�V�v-����?w7�C䉧,^����N�&^���`b�_�1�P�OP�=�}2Ң�q
�1q�I��I�<�;@@�m�<3F@�D�n�A��.$���B�l�<���Kc�Ȃ�Y�!~r�h��Mg8���<	�'�)AboI OR����FTc,���'ݤ �@�ގq<�%"�MC%Ekv����6�l!Dy�D���N�H��Ԃ�f��=�ۓSj�-��
C�<t3��>w���=IÓl6���;+�L�Q ]�R�Ĭ���8!�7%xi���Ӑ�����ғ)%Q�`yC�w��G��`�vmA �&%�B�ɥ!�&��Pa��@�)	f�:@��B�	�@��4�[���Ljg��8\�B�;2Ŗi�c/�*8���P�^�BC�I�6�x�9֠�GG:Ac�/�4|�C䉚#���!�OCQ��(�S`�T"�B�I%s|�X N�OX�v�߫"3�B�	W���Ho4.y$YKw��F�hB�	�EW�Yip���"8堀x��b����I�-{0�K2mϢ
*
�S�i�.l��B�I(0 �8�'��'�i*J�iH�ʓ�0?i��%~�Lٺ� ,cRvt+s�P�<���:�
�D�ڣe��l$��K������`�D
x�f�(�2~�h��s���j�/U=ܰ�s����2F��d�İ�5�˲Fq�䝑Ќ���&�@%!q!Ét�()�c�%�t1���hO�>1!� U\Z�E;�(�&>d�qd=�ļ�L��ɄJ�t��kU
"��x3��4��'^a}
� �	�cT�D#��U<=s2��$"O��Zr,�;���`�
E����"O왒e��� R�����p�q�"O(�q6��/@��N�C(N���"O��1��%o�\-Ӳ�C�v,{�"O4i��S#G:�����b�@���"OB�KǢ�yݒ4�1I��\�H��x��'��!s��)��y�R�1.N���'H��x4�Zъ�P.ǘf��Л��0����]��dC�j�x�)1@J�4+FB�I4@_Rp�&f1��c���C^2O���D��N�@��⛐N�ЀG��g!��,Tx�L0��P�8�v!�F`E~�!�,[>�C��:ш��-/��'1�	t8��F�S��j��!F���@3D�ĚGIխmˆ�a���P��=y�Nq��C�F>><�U0��ɲ�NY
FC�7����M�h���0R����B�I"$^���gܔAR��3���R��C�I���̋b�;!��]��$S�i#BC�ɚz�x�����v���! nV�n�#=��Xߦ� �߅#\6!�W�ԏ[�:؅�딩Q�<22�<�R�A ���Vc��"C�QVt�P�''�m��Z����f��j!���
$F�'�ў"|@��j�%�u�@&D��X�g�Iv���O�*�q �G�69`a�����hˋy��'(p�˙�K'�@X$M��#�,��p����'��x�
I�/��g�̙/4h�/^�y����p�.�g�+;���N��M�˓�y�>	���7,Q�|�� 
e��Y�J�<�TlF��!�E� �z��W��B�<��˗�xg�p��	U�+)�pQD�GWX�� �Oz�f�԰U�* ۃ�%Z21q"O���j;6	j��$S7� ��D���)��Wr2�H#���2N<�X2�ƶv!��QGZ�jt��v6�P9�չVd�?��?15ň\& �0F
{h�[�Oy�<q�Ĵ�i�SJS3�v��p��P�<	�#V;XgͲ�_�^�A5�K�<	R!��pR�\�+#�(7K@�<qel�	q�仓#E�W�x���A_U�<)uf��@�w�Ĳ@�q��ΎS�<Y!�������C�R�nP�2mӦ-)�)��2���h�L᫖�J\R a:D�ʥl�<[�^�:�G���t�� ��<���'�Ā���װz�>�Z���U��Ԫ�'�"M
R̀�G�i��E�&HC��J>Q��9lO�X3��~}0M� �]x�e���'o�x��1&�D���(R<:4�A��NC�	}$ܤ�SH
+/ P�F��&�#?����(�<�	¨Š��4HX�~���+�"OԔ��荞�
�r��Ѝ�T�Y�"O�R�H7S8r�jT�8��́0�i��O`�)��)��	��ܠT	7f�N� 1D������1$ʌ���;�|t���pӈ��*�O68�a�#�^�!A��q.pA"O�%H#�ſ�,��jV$�tJv�'��'N��Q�/K�I�L@����A���h�'f��˝
(�29��"L�*gi����<�'f�R��T!_��H	2�	�em$���hO�>ZS��,n�	�wL�4��8ZqG�Oʢ=E�T`ٗ^��HT�W1Q)v=�g�Nu�	Y��̸qK� �d�[�@�!0"!B��!�OD�-O� D�5(^�dl�UR�ʲU���"OH�'�������T'VON@B�Ih>��@C_�B�l!�d�r/�}g�,D��c����Y�-���%o�vɳ#Bn��F{��	^(
��6ᑶE_���7�Ē@q�'�|�KT�-'�C|0H��4�ٕ��d��%��B�$񉤟�è�!��D�N�48��8��*D�t���,y��S��3nZ	Ä�]��hO?�D�,���h�ZG?��27j	a/!���@
$��AZM� 0��Ęn !�dc�Y���ߥI2(��IY�K�ax��	(W~���U>{jbP�1��C�J�I^���˔M�Qz�Xa�/��]��4	E!?�O��Oj�zdV�D)$E�&���cP*���"O 1����F�����[�[^�����0}2�i�ib�� K�Pxu�ɩJ~��C$6D��಍-Eҹ��+�=�=��2D�H�+ʷ���R�00�B���+D���@�[>.)�d�ǔ�|�ڱ��L)��$�O��G�$h��hqi�-'���9�"O<�z�ǎ�(��S�-H��%�g"O�D�ۄ��E��A��4F"OR%�wJ�l���4E#s�$T"E"OPx�B��T���áC�;.���T"OԤ
�`Y�,�0C�#�`���'��se/U,r[~�i���F�8	�'����.��@��L����!�'T�d�Q�#S8�H�gL��@�Y
�'�~�JS�Z���K�F$L�	�'���3�M S����%T��t`��'����AН<�$�֌�:}�)`�'�q�`Z�P�h���L��tt��'Þȣ`�ҪC��)QF��c��2	�'ol"��jLH&LBO�ta��'h$��Wۑ,�p��r%�$>.��I	�'�f����,m1��c�H,tt�X�'�V����PqbW*,�@���'��ٲ7ڰi��pŤ	axdJ�'�1Ad��a���& � )�	�'�x< V&�c}�%Í�#��	�'c�c"T,Q��q:6
[ �u1
�'i�R�i�-x�m�f�֧	G6�	�'����U�XU�xɒvEӤG��	�'�����W�R��(�8d�Y�'4��YR�E!s1,(B�S��R=��'�q00��*�l]���	W�X3	�''�r�O�9CD 1�R�@7{��;�'�@d��N�eKf�����\z�;�'S"dY7f�5aRu@hм
�j1��'O��R�G�EK��#���LP��:�'Tmq�J؟_���U��-#���'��	CA�\�hH2��ܘ�$,��'�����n҈|f�*D��2�
�
�'��}�2�R�mK�i��oY���	�'y������v*Ra '!�>�H�'R�iz+��c҄�$�
�E��j	�'�l�P����y���5C�'��L��K8(M�	s���#�$0
�'���s�+W����NM*(@$��'yR`'jK�G�W z�ذ�'��~�<a�(@0AH9C�R90&|�f"Xx�<���U�Y��m�V,�>D�<���#y�'z@3�+ϫ�DaӴ�鐼cP���3e)�����,z�!�"y� ���
bq�4!�'űJ�>)��h@�hy��16���?�$�>� ��*�G�7'L�R1藜BQ\��q"O`�X��Q�Vz|�3b��^n��J󾞒)jdɕ]���x��W#�ָ��	;G��=�ծ
 -H�-I�_���$����ք����)�e��:�ԋ ̕2H�U�F$����H�#*�Otч��j�Rd���˦\Ҹ,2S�|�K&]ְ8��~�dL��Eܸh&>)q�K��v��(.ۿ��I Sf:D������[�FhAwb_�LV�̉�N���	�%�w!���4���b?]9G�F?!W(X�<*�ⳏ�f�!R��Z(<!4�2�t��s�\��2�3g���JF��G�:��� �σ�pA�����D0�~">��Q�Gd�Q�e��I�X�q�/�H8���v�� ]f*�[���8*�Jd��'��@ a� ��ڨ��Գ.�e���a~څ�&M�E�i�x��TH�;?�E�/�^��X4H�$�4�>kU,�2o���'wӶ���\('?�Q1�@���~B��,��E$(�p�(��t�<S�h�C`�E��1Q7�éL͂�{%-��<�u4��t�ڍ|4�0�'�����A��7Z0�� 5Ŷ0r��D?s�4��F����p�Ng&]�N�17� �gM���g�Trc�a�4�١u��*FĎpD9&<ړP�]�2��j**��!�vm��(f1��BB(l��'��Q� 	�Rl�q�	�[�Zab��Ԙ>��)�Ο.����b"��d�^��S�^�p����Dɐ�.I�,�/c-0���aH%f�	�7�������!��Y0�D^�MO�#+YJl�EH2	��|�pL%Y'd!X��J,����V}o�pؤ���a�=Lh`K
1&BNY�G�:{��۷f��f��(�dU}/�����;x`t	ΟL,y7OY!u�����u>Dq���ڨN��D�S��7o�ў,A��V���F
}�t��7���D� Ը��8B��2t���|�TH�рLmv�г��@1��G�I1@�
,2喭%̞t�W-�0�䀣"Yv�:l�z��ʓ��\��ɲ#T�y����C�%z@ŮO�����X!Ĕ+�.ހ9m@��`��}�U,q��Hx�">�*���$����M
�z�� .ƒ>�p��]--Έ8p�(�t ���`>�R��C��z�D�F�P�2�<�OR�RN� ,Rt���fN�|#8��B���:p�ܭke������/N\����'Q�����F.�#Y�L����������חI� ��� ɼc�G|R�Բ4r��r	Xd�	34b��e@�[���X����B���&�A9cQ���	\�b�n��ng�#�ɄPk�ρo��\�iG =�P��'
t{��� N:�'��؆�M�f �3���X&diT� ]ϺX�� \�q�����NQ�MM��,KI	�}���R_@yBP5u��l��.�������k���2O]+||R��J*kJ&��.[�,��˧�ܘ�AH�w���Q�� ?-M�Y��	=
б!qn�5p#��0�;a�"����5��@C��N<�>�+F�B�k�D{`�	�i�Ls�'t>���T�\���`���ӊ��1#mrX`ՠ*�	�7����V�Pu�D�8#J9K��xSk�.h� �h���0����ρ	6���F|r��(1�t�Y��U����{�����yrW�fJP	yq^|����${�*H�s������xsH����.A�� 5`P��D0K�lɻ>x��,�Oz��с�!�H����1��$C���
5@7f3V�At&ڎY:6�Ԃ��Rpt{㕜Fb�I�ih`�&A�3���h��\�a~�搯of�}��Af��H��EX�r9�E�ӏn��@֊ɕ.\����pQ<��n�N�'��dׂT� �֫R�:p�=��Ժ���r����nIBp��Іd|��)ŉ%`��!͢iEiX��CU��qB�Q�$�F�'$���ӿd��@Qr�˲+��<�	߰ai� ��%9}���,��%�7x�8���D'�,d��c��Ř�g��=]��Xd�(��)�b���ǀ�.���K,?ɡI�PWp�dG�F�����$Н���g�=�RT!Tn� ��H P�J�0?!r��<t��9$� �G�ʕ�Fˁ�AI4��]%A@
Bቩ�� �'�ңG�q�Ɵ�m~V�>�@O3xW$5r��t �Wi$��b�M�^�D����ybDШH˨��3�ǶT�@�����$�`=����{��I^-�Y�@c��Q��X>�!�$�<r*�[�o+*����
��b�!�V��XR�Qm��15�� ov!�� t��ٻf�`�6<[FB�F]!����<����:3xzbfV3>!��&J�(��	D2�d�f��^}�ᙁ#�T�P�϶l��)���u�fQ�@�0�cQIW�~]K�'���2��G�H�ӓ-ͯ&����OR52�ܟnkv�1$G?��O��#B&�ޘ���6bL�0{��'ی%��6`愌����`��8� �P4),r�XG�-hU��'��!�� Fz0 ���\=V}���$�&K��C�@�"Cp��-�)U0�`�ݭ5�<���д�!�� j�Ktc�UqNlڳ�n�,5�`��9F0b!9է�87�=��i�ӟ"~�	3���s�et�ъ� �B䉾rr�WdZ4`�]*v�v���K�y@�mc��Z'am4���?�=��ɗ�l��1p*l� I8�ȁ��(hh�%eT-�Z=��C�0��E	ж<^��Uӟa�![�az��ȻE�@�sE"+�<ԛ4j־�(Ob�{�I�@�L�#�bo1�M�4V]��Kď��w�����&Y�t��E�r����.+�L`{�e�4"4@8 $�k�p���7$^j�qS�Å E��fK�/(�B|K�%�Y����p����|1^�pC�I�B,<�"O�E� _$�� �I�2�ȑ�����dߒI87-̨p�	�OI��D���)�tt��d@+|���Q��!~8����!<��B�'v�����N�C� ��L*ƴpq�M���A�
�+�ܸZA�'R �+�_�#՘��&Â"]����
�\����҅�:aV�Aw�[�vpa 5�:��
2� $�d� D�b���1!��pY�D��&�ܮ(h�'ٶ|kHb?AzU[	u�����,�2{��С�k'D�4bv�Ϋ?��6KA�d�lQ��O��#�m��[N�"~���Q�wZ�8�� �3{ǐ�r��>�y"��p�%�@5k�̵{b������ Ӣ��N	=��<����!��BЍ�3N��рh�L��DtǆwBZ�P"���� mTJ�%�Kh<��%�|g8}��d ��5F�A�'\�(�WƓw�O{L��v�? �[3f�045��
�'�l�;�k�#�@)B�ص!(E�
�'��l��EV# ��X��N�ę��d�RM2�~rW���a-� ��CL�m��E�竖��"��~<a}�	��:�y�u!J�XX�k�뚁�t��3 ܖݸ���YR�C��A?���ٳW�Rb���Da�xC�B�<Y'mY�G�x�a]�nv��G�Nr?!��B���u�3f�	p�����*}J~,��;�j<�A�E�q�t4�A#�r8���a��'���[>�ZKѠ��y�T�%��\U��C����a���|�'��"�2R���p�LM<����Z�T��:��	L-&�lӱFE('���@�-CFUxE"��aL�����)�0>���!�&�Bu��+G��17`�Pa)��Bk��?�vAU+Y�Rp�;nl��/#�BpyV���,u^m���H,#�^B�� A�(����)>U��ǩFZN��|EB�R� =M2���'A�w�Bdԟ��O	I�A�s65�S�Ƒ
t�T
�'�&�!�F�Ր�"��'zP�*gf� ��((.)�����g�R�л�a�F�TY�l;D�B�?i��ڈa.��|��
|�lYs�̢2*�p@��G�=����K�d��0�⍇�0>A�4�v�y�aȍ�$TaW�C/Fj��asN7����?�i#.p��p��t>扜D=����@�1A�p���P�*��ȓz��Ć�a�VŃԯEfD�갧͐HkV�	�m?N�N�A�z��1l��c>	H��@>2�NA4�&���
s�!\O�0� $��h�'���0Bn�h����'+ؘ��/(}B��9R&�iԟ��{R	�6<�0�oH�uW�У���'	�� ɒO����}zpd��J��pb�O�v�&�	���M���P�%c���`��}E�}��D-(�ܩ���7��|��dڄOJܦOT����6�:�����9T�i�Q	f���
�z��'����g8D�T�$�+��#È�U�`�* `LPM؍����94�H �k�<qgn)��$rI~r��/G�8�PI����Хʨ�p=Q����k9&T�r*h��p!��s������^>x��s�a�<#��|��)+`/���0<!�	�'RTjY�O@8�壦k�pܓ��I�E��0O�<���M���3H�(}9U�^9�t��������Q�n�Qw꽀m'�O��)�Tf���cBP\Q2��A��pE�YHM>�!�uK�}8�F:#q�5s���ݜVk/FxR��HQx��c�,D����[�@��m`�
�!Y�6<��k�O�qK�H��S���E���l��\W��5�S64PӢ�,t� TZb�^�m�:H�ȓ�xIH�ML/[	)�q��5��e�a��v�����@Q��FE[a,�d���P�#�@���f�1�t��/l�a~b��O��Q��U�G��(�O*:�8!�U<k^P-�.M��"?� ��1y���I?� i9�bH�F>�U�R�e����$E&���-���$E�2�l0����'}�Dyc��	"��ON��~g�#~�G�>-�y@��ZZ~vRF��g�ɕXyb12��I�~��?� ��Y%�L8f�Ft)s�סTՌap�eV%ĜK�N$}�+�g}"�Z�_�f�᷇E�dة�c�h�Uʵ/6}R�F72��\�xt��F�7C��ֶ�|yl��l����Wf	=:�a{��5U3@��W���k�,���MчL	XDcE�*{P^<D|R-Z�rب����˟���2|,�!�k���m	ţ(LO���"�Lߴʓ0&!k�m݂[ɐ��$E'�X)�>���6PE����9�'Q�t�j!%E�0��pS��Yi>U�=���
4�(���*3�ҕ���tZqs��3/ �Rï܋/n�'T"}�'����"R ?��l2���zC�D��'�Yx�n�9�^H87�r�5X�4
��IB�\	�b�LR�G�	
�1O��h��y^�Xz0`�`39xC�'�Qa�F!jl���[�8@�xK$ܳ��X	v�<�\�7eY1��<Q��׻7Ȋ��S��05~�ZtȂl��_�M���]/��'� �j�.�:+��p*D=~�����i�&e�(Ւ����F����W$\��t%?"�|$�ċR�:�~ ye�E/HU0c�(Q%�D-L]"�"���w3� �P㐄M�J�8�.�0h?���O&drB�(wS���䘲W�x�2T�%x����7mƥh�/�*FY�aҗ)
j���������%��U�{A�xG�}"$@0�M: 8��ȓT�$	k��΃z�1b�ͱM~ԗ'��b�����O�y�naBV�I���	_�T�X'r� �n�i�։0%�����>!u@�oٖ]�a�߫7��A(cɒZ��!G��c��B�h�T;�8�M��G���%� ��NM#o�T���G!���F{�kÈ:����H[o���jTC��k�B�
����1��%����u���
���DS&7�$��#�=y�x����
��>7,��gɗ~������'Z0���i�;[~�M�sD�#A��Ip���Єȓu����wLھZd��qLY��H=�'��̫AB��!8��J6�Խx�Y�O��'wBV��҉�4(s��ӎJAܔ��	6��I������������I�cF�u��e��*܎of�p�>E��RMx@��H�c�]�(�T��m�>�[ҫ�9m�r�a�<s	��'��y�ċ��z򍈛z�A�Ϛ
'BX�P��;��>Yǣ�;݊6m�$J�Xd��l�p��`M@*n�!�d�^��%2�
��Pʶ'��+�!���N{���V�eҌT�6�X>A�!�R�a�m��� �~LX��2 
!��O�gpƙᣦ�<Ҝ�XT��D�!�$4M�0�r ��1c���k�!��.]u6��a������O�%a!���0zh�w�/g#>u*Ue�$f�!�d�3;�Y0����,,9F�5!��ޓ,v����M�xx|�ve�C�!�$444�%�Ў=��t��e�j�!��ȧO�d;�JX#WLe�7�
.(�!�R�"�tad['����,v!�d��e0a�c	7�.�vDĥlt!��2{�|][��L� �P�����!�D�|ҕĬ�t�e'f�!����ðJ�)�V��E�H�L�!�������eѬqP�+(tM!�֜PL�js��T����K)�!�Ğ�3x�Yr�#G<z��E@'�6�!�a�J9�n�)7�-�V%� �!�d�1:�,�Bc̄�.�A%�+-�!�'ׄ}��հ^Ĭd���!�Y�Z�^â��f�`uY�O�m!�[�jI��
K�~�2�p���!�Ę(t(�'K_�ԛ�e�zw!�DY
��93u��,H�0B!	��=4!�r�@��	�/@���3Ug��jĄ���)|�����L�C$�%[�|�ȓzW�����2y�������ZC� ��%�)�uhΗU��x;�Ç���p��(�(L���H`#��]��l��V*
A��\n�jFE�	��0��S�? ԉ���M��SUJWzT`���"O����.Y���� ^1xI��!"O�&���AUn����%!%ɷ"OZ� (� ]B��?'��kD"O��Q��)#vdФ`J��H}�5"O� cc�ɵd�H ��o˳7��M
U"ON���F�����Q	�:�3�"O|��.A�4�S��DO[�msQ"OTx��%�r�N����E*#LdѲq"O~���I\�f�:,B��
��*@"O^�cB�ĳcv61���8K�|�a"OpX�g��� *U�5 ��L�"OT�j��~�8�r7�¤��=H�"O�P{D(��ZMș��P�"G"Oؙ� a҉*�f�j����\�8�8�"O<�hC(Tidg�� �
\R�"O���R�.Zmf�!`��7�jDc1�'�\(��˩$�����n�-,s��*�C$Y;��[�ObT���ÕE�ԅI�j
3_�d	�`�	�K~pi��H��1�q���IЃ��k��_�t��X%"O�q��M�
��P!.X������'ـ��͔A�q�Z�"~¦�X7C�6��%f˼uS��`����y����l�&�:�`V�lG��
�)��̃Zq�5!�D(S������I�x�/�Ί�3���<D��}�@=A�ݱQ$B#d���5@���s�oΒy�6(j�OB`��+n�|�ĭ�$4�����I&�1
j��#�6y�|
���C�t	�o�7p����!�b�<�m�9P�:0��~&�  �Fݟ�+���'|�a
���Ly���ܙ�Q�V#��G�	 3�Y�S��B�
�2�;��:n�D5�2�ѐ~T˓^��BuHJ�BK�AqÓ6��}�dm	;~X��ѩ��E�}��ɘD�aQ�i���9#��7���K��ݗ~�����X<��ʚ5�t3�րp9nA�D�V�'�Hq�f�/b�^��}�K@�M	�4g��бf]N�<�T�ɶ_���Z�jP��$1��'SO?	�T2V�ޭ8M>E���S���:�C\/1�|# �P��y�'J�,��U�&'��G�p�i��ԧ�y�r��I�i�� ���Wn���?	QA�&7�^�*"+Z�:jas!N��z�#��54� ��(�  ��qQ�*l��H�2�{�**ʚ���O��ě�l�n`�a��$��E��'qpA귄P6��QB��-,L��'JaPë%�<�O?	�f��%A�$�5����xz� D�( g�� ;9��`���3������!?с�0l
���g3OD�$��`��g \�z�(=���'��
�%,N���a �_5@8���3�1�vA�|(<����0W�4(��L�-���YGI�q�'��������}Z�g��t02ֱP�Ԓgb�l�<�7/�$Ű�vL."���r��<1�[�o�L���9}��	��3��E�>�٢�*�?BT!��
r�
� u����v��s��2VW��1���a�՘g��xR'F�A�a��C�+�ɕǋ/�0?��e96���e
��G���j� )u�u�Rꑔ]��B�ɠ_K�XdM�\,���G� \}@�>�$^G�,ш��T��
dh�c�*1�e�N�yBK 2\Pp���\��l91Ꜽ���ۇ�6�ȍ{��2�P�GN�U�h:q��+!��q�6PR���$���M5[!��s݈�J��V�B����?`�!�DD�
��6�t%liQ���$Y�!򤃥(�}z�%�f��f &�!��Z%&,�HS�(T�`lJy3f@Y.��4D�Fa��tq8(O?�(Q�V�4�@c�UL=c�]�<��T<x�$��@Ӗx�F̫� ښ�~2�о���w�<�҈E
� @���$M�=�Y�e��b�89d�'i���PSm 5��J�.,~���Yy��Y�+Є.�(5���'E�q[v�H�}wR�B�d�".d����F�kM�Y�EH�x}F�r�$:��a��eF�s���ct#�@�!�$�	G!���v��P��(�!"C�B�Xd��=h��Z�	�!4�)�)�矸�`�E���%�;t���7D��K�0qJ@"�˘>�$�D�T��?CG�&Dc��уj�1J�B�3ړ7"H�-v<�e�H� t<1��		!����������	�3\<��	&��,I$��<�
y��3;3^�p��'��#���1�z����*��h�����s@L�3�n���H{�7�9�`��(�W��1���?����@kBFh<1�BO�R'�� �Z4U��8"�E?s)�`BHQ�Yk���"�Z�#ׂ�Q ��0����I���҉��c�B[�]S�m��La�QG��>A�"I�0o�\����4K�d6�0N�y��C%��S�|��Q��!>��A�Pں݀D���N�Ru;Ħq��}��p����ĝh����L%.�$ �[1�4A;Qg�8;3�
;L�xy��'^\ �/(��x�m��"��,	�#��iEԃw����+(�E[&�ۻ&��%?$���J7�(�ar�K�V$���4ړR}h�r�°If�b?����9���!R��&U'RH�V�2D��q��H��2m�n0"d����c)��6D�&�>E�ؕ9�<��"�ع9�(��w�XY}!�R�!�:ْVj�"9g���E�ë#��	�X��)3W��ay쌍P�Q00,_�0�v�IQ�0?���öbbd�0R��t����B	�"�x�s����xBj�-?b��"��$yR2T�ϱ�O�H��cF?��D�C�gS�Ջ�)�?4��li�"O��r��&R�)i�m�@쎡("O����DSNC��� ��*of���"O.�0U	ƥ�H��ŋĂZU 0s��'�dT�0�TZX�𘡡ҷp#(}S�����(Ue1lO�(��W���� -�ܠ�B�A3u��� c��_�B�ɭv�@]�����q��%k�F�s�㞰Is� � �b�3�mS�EB�疓���Ud�D%�C�	--���ʄ0Ԑ�+�狏]�r�R�ϸ2��'��F�,O�q O rsR�C�"ݓ.ڄx�
O�0�W	[O�~��ę�� �֠�7I�����nF?I�D����4D��cQ�@=NTa�ٙp�L0��'���!BR
m�֬S5�q��QrAT�"�4�t�Ѐ�d�kǬ,D���`�� ����GR1����<�ꆞJ�phԨӼ(�<�+��I]�tq4�p�͑�NQ��G%N;!��EF"ݫp���i��,�@Y
�$S�%��J!��2���{"�	vC���ԁF5Er���հ��'�d�
�	�S�O� Q�%<'���`�кkYԠ7�ɤhda���� ����'�����B�A&D���,2���iK�L�(�'���'O�"�{��E�/ʊ�
S�<�4�]G�Q���.�����EC �yB�/M�Z���*����H��7^D���4L�:8���A�'�x�e䫟�yů�ŅH�z�წ�6��E��j}>��뉨8|��b�۞�������4���Nʲ02�BnD�O�u;�$Y�!В�qO*)Rp�¸/��q�E_�Dm�h���d#5^�h��у��OX���`0�(5�"
�``GX���p�ӋS"a�I��@�ʈ���Iv�3��Y��ek�M̩���366݋f��RޒI��<�;q�h}(B#Ԍ �X�h]��\��$^I���]�L��;�h�j} 0�`B�%!���4GN?1�b��'�v��k<��O���A�,�;�:� ���
	*�ə"�'.�mr�xt��͓���ys��f��9��As��ĕ'���:��ٸ�!���7P��E�T�C�N<��ߴ4���|��LI��Jǟ����HE��"g�R�K��z��HO۪��-U6+&U���ګia~ү��Ngj�yg =)�F�,S���ɇn�1�ƒO��g.�%0�ڐP	�k&Nt�4�y��Ƃg�`|�k�l����`��ybb;7ž���i��E��̈�?a�
�����"}ƔEB�7Ǻ���I;��%���r�V v:���爈G�Lm�ȓ;f�x�ICP��,p@cۼfE"�Hc��4)�K
�3��C6$�K���ė!p�̍���[���4���Ja~r'C$�
�k� L�I��׸1R(�a�@�
��nT�1�b��a��A�'�\BwHOh?p��N<��[�G�>A(
�A�n�{x��s���F$�i�^�����ĥL��� ulZ	�x+/;�In��q۱��I�O��%��Bt^���A33���N>�FF�15���)��=�'6ݾ���a�����bL,K�۾x�N��H��Y��1�N��i��L�ߖA�N��R��V�8��N�� ���a�g�$���d�g��!r�]��"U�9ƛ�d��0[B��r؞��s�-�89Xbj
�ua.5���>�,��!Oӂ$��DI�nͦ@�6 +��'��l��A�OIL���N�m�De�$� QI3'R����ȖN�\��WAL:Q���Bڳ<ܱO䠨V�δ%Q4�b��)T�L�y�PI�S��+&P�;�qO�� hM��0|�qD@8e��������%���M�3�̎��	��H����0J��ǃ�d��fŀEP�B�	�y�� ���>����锗U��6mG�Rqqrޣ�'�VyaRG�c̓�*5�dkҘ �~��,�;�:��c���� 8B���m�,?g��H�`K֥��$�0|��B�6<O��JWm�iA��ꝅL�aZ��^1Nnჵ�:�I�6���z펑$����BL����rc�iQ��m,� �=E�D�}��)������Ń#!e��������'g��g� y�8�$>�]���9���EJwD���P�B��%/"D�s�M��p=���F�x��H�P������Y�j�����w�YN4#��>%>�⧑*B�p����ϩ߬���aV�X�� k���!�$^'mФ�B%�I����7g��_��Zl0Erg;�vI�w	�0�P�O �'u�l�&��j�2�B���$��Є��'&���0׉�.Ee`a��
�U "Xr/� u��xT��z���u�e��,���Bc�ˁ"�p���>d;� �@` ړ �ܸ����>&&c?����6b����D19��|�����8#��<(�����'uʔq�
SYW�y!Эҽ$��t���7�:��� �(ӧħK�
I�1`ب��c���&ɛHۢ@d?D�b���uZE��ٳ+:��*�.?�0��2eR|Xau�ʜF�����b�T>ٛQ���b5��`�2���*�O I�B/�5s� ��c��v:B��P�E�HN��p�*П<6�Pǃ���)��HZ�[(��`A��"O�T}�K&D�����L�<$Ha��-G��9!�>!ǡ�q�f1:ד`��PlW-d�@m���N1����J9&�i��9m�-<v\+F*D�)O�(�'�v �@g� }[piV��8+�Zp��'�8���.�P~�0f�W�j��8h
�'��$�U*��X-u	Äm���
�'�Dp8��+���p���f��3�'葱k۸;Wd钓��1o����'dDj%ǐ1�����A�d���X�'�����[+�� 6��a�,�
�'�(`ҳ&��i��6�����'+@�P�βHA��P��M�sx����'j��t�D�;��!ɄkF�2Ŭк�' ��Rl�I���"��
3��%`�'����5�ږ֥ ��Y��:
�'t�����-)��ǏO�4���'��U`wN����S%��=�<b�'-����F��[�(�A�h���'��pC��Ǳs��x8bK�!>�r�	�'	,!9�f�֔d�!�I�.� ���'�e�E呃:�\L`����&z���'1�����	�E<N� �7�(E��'�,���փD�(�9 ��"� \��'��ę�&�?GYV��.4�ܱ��'�P��ŏ�At��Jd%A.�hQ�'v���0l>�Ⴤ�iv����'���{B��b�\[h� �ʓT��vM�1G�|��#����B�Kњ`�F{t-���?q!!Hk>��/�(wʲ��<�b���(a�b�z���-�^<Ƀ�,�N�	&�'�2�KWDI)�@H��@&O�4�*��;tD��(��I$|`��h�l�T�I��Jz�]0��� ӊ�c�hf�(�f��~r�4b�Z9�Yx��3� .�k�#1�ݫ�@! ���%�O��`��`���Y��������O�at���V-j!� ~k��(�鎛�M�"�*E,&y	�O��]#+���Z?�韬l�d�[�&m�}`��PR��\R�貟0a�il���RyZ��)*���}k��8B�
"Qgk�2��MاV�T (O��8ʧA7��c�&9p�dQ+���F~����O��q*�.B4:" �T� �P*���'�ș�5�(~Q���@��x�'�ʝ��E�"�Z�R��9)�,�B m�%�MKA$<�$�K����h�Oe�q���P�o��x�ɋ^iyM>q�˟lqM��k���K_+��� k�"xر6�K��~R'\�Yr����p��ӰB?P�s�%?�b0�#�g.V������~0�B>R�S�'m���"�4ZH��`q�_�*BxU�'i���IK?�E�O��mE�[�����0AKD�i
U���3(bӆ� Y���M�O�*ո���k����i	�F��A$��x�OR�j��l���R%$����柏�y2/I4Ҩsю�;6�u2n^$�y��L�TS�l����!�@X[��F1�O��G��v%9��ޏ;T|hc��V�eu#��� ��HO�4LS@��be.J��_�sI�8&� B���i�J�Yj�X�r{< �MM!l�剏b`�����t�)ʧEU�(���?ִ �U�Y�c��ZD��O�\�smK ^���S�S�	�⟨ � \ X�=�ia�)SI�<Kg!�$Q4n��Q�F�ŏD��t�T��,!�D��s ��Ӄ"�T�.��Ȁ�D*!�ǖH�����眩���s�!�ą#)y�L	p��}E����ہ/�!򄒚���s�b؞?I��Ȧ�5j!��!ޘ� �T�)��"�)X!��5�`d���/9�[D$ B,D���cE�0ow�S�@�R�$T2� +D�<0r+�;G�2�`D
%� ��#)D�����6p���`�W�o�m
W!)D��+�ٴk��W	ZbK�[� +D��(Vg�  �歨rm��������*D�hk�鋵tr,T�ԊGP-�)D���$̾xT�٠SGЏk��|�Vk)D��-�+|d~�w�̭?��أB*D�("���YVD}��ǋ/d6dD��*D��[�*�4;���xS+]�FLBK5D�T��ș�B�H `��*O�� T0";m� � o�bt�!"O��4��,�"-�����DlQ)�"O�a:ãO�mR��+�M^"~0<���"Oֹ�)��=P��Cqs6"O
E{A�}r0m�C3)�ި3�"O�E��ϩMDr�E�D��p�Q"O*�p�F?5����!A���E"O�����)&(̚U��e�+ �yr�I�4tQb�K=)-�c����y��Y
P�N����8 �N仴���y�$�$$�q���ۺ-e\��ղ�y�l0-O�SՁ0O�٦%���y��[�ضM&n�Ja|l��m¥�yRƇ[.�ڢ��'-�X �-�<�y��WX���hB��*F����0�y�fU#2���v&��Z<���!�ē�p>��EE'B:��AVA^�'�Xiq��x�<��� .�E�6��9Z������w�<�e'��5oL�2�ꆚJ�`d*Si�<���H"X�hXR���j�ó�q�<�C�Լ:{ȅD�b�<���n�<���ݠ,�&)��@Q#N��A� �n�<9G�_�y�1�AFG�gԵa�*_g�<IF�
<N=���D8S@��gTc�<� 0�󤍅.<��m�4B^�B�T���"O6���-���Q�2!��^
t���"O�A����=�V0��"ͻ����"O~+��_�G4v��4��j��8cR"On(5F�<J��P#�Q��[�"O�I ��"d�x$��

Z��1)�"O��V&�9x�
��A�B,�d�!�d;;���G�̢�� ZR� 
v�!��)�X%Pׅ�2N�����ź	�!��ߣ$ɘ���h�kΉ��OB!�d�F�N1ҥn�
a&�k�KE�r?!�d�)K�e)�gM$<�Ȝ9�̐g!!�Ċ4I�T�qp%۾,�$p9 nC+<!���<th�Ȇ�f��B�ӈ/i!���8t��ݪ���t62E�Ӭ�#�!��֛D�zL(�AH�.l��U�F-p�!�dQFx �c�!Y)�dBW����'����&$M2i䟶vw���'p�݂6oU�:�(Y��,�%b��
�'�X�����J\�!��ؽMvva��'�~}�4��$NHs o�9F�`0�'��i��ϕ_ʨA#���>zxr�'�4�I�I�GXT�4��-GL���'N�X#aޙL�3�1:A��3�'1JA�oK�
ORU�uaI�+\c�'B83��4�f��e��[ʨ0�
�'b�u���k��y�i��U���'�X�+���i"d��!�F�d���	�'(�� �^���Q�VQ�����'o=Ҁ�[� �N@�ѤI��Ȉ�'�>��J
N��#���/#��	�'�`Y��,L+_���p#φp.�(�'9�1I��Y�OG
@�)iT։��'q�}ѴOH2ERr�V�\1]�\��'�*ģR�hb���i͋Y�$���'3��2� �W����1G&{y��'����n�%OP���C�;����'6����'�):xTƖA��,��'B����L�y�`�8ti�?���2�'s`a�Ӥ[-lH��S�dI*��	�'N2qX1&M3)l����0E(���
�'�0���_*�􌋣�ߡD�=9�'�ʹ1��γAB��'���|\��'/`\��+S�TP��B�$�
�'�$�CI��yژz#ρ�v���'nL�VDǬ#�.�bnQpU����'���)��,QD�SbM UClp�'.F|S��B<\*L���#z�[
�'��1`lR�:}�Y� b�waLur
�'��d���̽p		Z���qT0�j�'f��2"�y�8�*!"_�h���'u�zBMA�6�5���\�M��!�'C�=�i���J��#�<��'P�i��Q2F����b�	�����'�D�ꅦeؾ�rsN�et�h�'�2@q���i�t�Cr&�2�]�'��[qm�]D=`q,�	+�\��	�'��|ӓCSp�&��PCԎ�͒�'\(�.7-�2�@�J�O�1+�'%��Ђ��$uҥ�C��MYR���'�� �E��̚GM�8Q�����'�P��w��@7��B�/y�F�9�'��Yr�B7�R�����uY&\��'���A6oٝ0D�3bcժm�jD���� F��F͑-|�t�Xv�E�l�EZ�"O�)�!R��f�HUlW�j�x���"O���֍�6+7���� 1�RH�"OLA��勈-tR�Eȏ���mz�"O�%k�EF�jM�(�D��,)����"OL�0T$/Q��A���:��Ea#"Oz��� Rhn`�*a��
�\8��"O0 f�ѧ�nM��c�pg�V0�y�㍖������A:x ����yR�$^]j8P�N�$E 0�"S��yR#PP1�|)�c,Tb��jW(���y�́<B�2�ˤ@Z�R�H��� ��y�%���%���Ţa"�96�R#�y� Q�5 �Thf�,	��E���y�M!R�T8{r�Z�͎�U�K��yRC�(L�{��ּ^=�Ё����y�E��H��)#��&���)����y�c�v
��(��F�$�n�s�a�y2M4R�@=:����-�+ �yҍOR����O��m��Y�y�gĜ;��A�r�֔�z�"���y��p�
($�ǜ����r���y"��*BS�ݒ�Õ� �ȱ� )L��yR*�
f@RT*ƆZ�j���+
��y2!�9f`��j8jC�5!oN��yb��-��ݹw��Ro<��R��y�	E���� �0yO,D"s��y��Q��D)Z%��qd$�r&�y�)��^���fM��q��$J�l��y��N�d#д0G�A��LĻ�G[��y��p��� fFI)��%(�"���y��G]*���!�$MĦD�E	H��yRe[YH@0��e�G�`z2����y� ց$�^�k��ʬ8��)��MO��yR��a���Ѡ#��} �O7�y"S������S�&�c&�Nv`��p������ǵ\8x[����U50e��[ޜA���61��04F��3���ȓ;�����0)$d��j��S����9�nPIGfn5��Q"�i�X���I0���$��ɨ6�%��9��|5�M1%G�?��mP��
�1���A�6m��*Xz�h�'H�#S�=��8��D{���6���� �(�0 ��[E���� F1^�{�b�s"�ȓK�`������Z�0�j���n�((��b�̳�@�!D|* ���9�ԅȓrE|�SS�Y����<�!�ȓ0���e@T�2M�� U��:Մ�]�	�2�L�r�Ba�P#�*5!�X�ȓ@���0Ƀ=\�����)S�Z���c/�Ar��/c��#��ȥ/6B���I�ֵ� W;m����M�2=��ȓGJ��jP�B�Pl8�˧��"F���ȓ ��MhWmV�?.��$��:������i����5tp��6I�iX�ȓ)�p��V����0�vC	
i.�u�ȓ"�(p�©\� ����V]Ҍ���F��!�L�v(d�����T����ML��Ҧ������,C'?V8��gaR�8�G�a>�����K��@�ȓdtqK�6xݮT�dN��ه�ê4�"@�dҌ����U���W�pt���)+��
-шs����S�? 6I:� S(q+N[�'�+s��i�"O4���HܓRF�u�O�3T:T[�"OPI'�2��蒇��,BL����"Oڄ���G5j��4�G�s2�Ts�"O�dY�+��(Ŕ`�(t��e0"Oά�d-�&
��a��
���m7"O��r���=��y��'�&ْ�[G"O���`�ű1�Z�	�,41l���*O�D�G
}�(D�L�6E����' v�A�<�`ؤ.�<�Q8�'$V(JɰBI�8aU���	}� +�'��ր�/�<�2�\�|�����'SBW�:ZR���Q�I�|��-���*D��P�S�Zۀh{��8=?�5(A*O����(I�1_49��������"O��Z�d�6
�ܲ�WH d�b"O�-�3�BG���F�]�o4��4"O������$���;Cm�{GF���"O�"�D+w�8i��M�P���"O�t��j�W�80p"[�
l��A"O���3#FV��W���@�B��"O���0兟Cg��G!��%�^�z3"O05�Ѐ�A갸x����r�ڀ"O��h%,X �L�үAK��$3"O2ͩQ�
dC��pP���/���s�"O�u�c   ��   G  n  �  s   �+  �7  �B  �M  �V  sc  �m   t  �z  �  $�  g�  ��  �  1�  t�  ��  ��  ?�  ��  ��  �  Q�  ��  ��  ��  ��  ��  � 
 � � �! ( _. �.  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�CJ�0S4���T:
b��'�V�)��/r�<��w$?��P� �d����d<?��A�7�ٸ& ģ#26�rԥ�]�Ij��P���	'&Ȏn"=�#+<O�㟘�SC�Z�\�ʐi�xc��p�"O��3�iJ
t�	�ħ��\���+T�@l$�HO��>ᢁ��r�P����:��5:�;D��У�E�[��"�#�P�ǯ5�	g��|PU*��M!d.
!P��@xf�6��
�Q��O���!��,�:�zuǂ$v-h�S�'Ԯ$�2�U�jn�B��I�^%��{��'Y@��͉	]"�Jp���\�zM����M��BK9v����H�1�L�CD��;��x�b�{�'�f��s���F�����̏� ���Q˓.n�	u��;�&\�$$C07�J|p)1?��O�b�"|:���1ԍRJ��2mh�b��(�S��+����Ӆ�o���څ��@.��=�� LOD���H\0C�� e^A�mHW�DS@��l��IB�f�
�͉�YJ�+�:�X�!���r��4m�5�,cS�>M�1O7�>}�	�A�]��N���&���tHtC�	"g�����Q]$lykSE<ߠ�<���"}�t��
7��h�m�R�\��1B]n�<��( !R(6�n�Sq�1a�k�	]�(pe�B��Pd�$5ȹ��>�O��Γi�&!�p	�4m��M7F{���ȓ3�xZ��3��e��A�z��|��Iu>5J2���W��cb����ȓ)�(�z�iҮ~�T�0�L0ngX��ȓg�<QhF��>�Ɉ����mh����S�? �U��7g<�E@ba��ToNH"O��0���5%{>D���I�{UЀ�1�'��(��k��S)E�jT�[7�����W`�9���F�'���ł�1b�D�=I��)�i`���0�Bȹ]2�`��K��yi!�DYv�2C�%24�y+��DP�O�S�g�m~xR�c�0�
]�3g��6M&��D{���&��j�,�2/S,OJʥ�j���y�A���Z�elA�DȊ��B�L��'zў�O��0�Elú^ZE�@�S�'g��
�'���`6%�T�D��#n��컋�D*O��qw �q�<e��мQ�p�H�"O��ۄ��C����s���l�V)*r�'�!�d@*C1���@�������:\}�{���'��"�6U��\q����$=�S�O۴��4��!6��'攫bp�Y�'�a{BM�>I@���_�����.k�Ɩ�����>Qv=u��#Y�c4�-h��Nh�'ax��C� ���6B�)�Nx"���.�yrE�$1D5{�!Z�p�9�`����O�"JA�I@�dA�N��*��q#{�<I��.ye~cs-�~�$�1���<�R&'�S�O`��;Q�@X�@��b0��:�'�|��	��l+Џ%m�$Z�O���I�_��D!o���U!Íj��C�.�b!��`��E*�%D�:��C䉳V���w�^%H���P�mЖ[u<�(�qO��=��r���Í��n>~��šM�e�㟸�'�?I�b��
���YTI��k\����y��\�b�*�)��њ&�Ѿ U`Hz��ɽ2��R�ट�=!���O�T�kO�#�^�R�ۭ7G�X'"O"�T]�[M�\u�-� 2��3|O�I ��N�'zL�6	+,����'4&}�'��P
"�e@�	�B,��A�Z�G��	��>��-�N �����1](,�#S�V��z`�>aS���,9�R�p�9
�
&qZ�k�4D����%آ}zdD�1U�)�%f�<��)5��Ot�}"�'��i�6T#�&�.XK���T8���'B��ܕxL��@Q#R A�Š���~���H$����51L@#�#����<)𭅓�H"=�!���h�ڒ& eƦȹ�OD�|�p,I�l��şB؞���Y�l�&�(`��"����>�O&u0��i(r�h�,�HPp��-a�j��'�0��Ô�2Ȇ�R�� (��J/O��a(.7�d�T�pґ?	�O�v1r@&"J�<$PA�S�Zd�@
�'m���o�$O���(�� �x��'�4SACi��AT�	L>�s�ɓ��y"�^9�y���{��yô�P�y���"?>�T�F��q��аTA@9�䓢hO����D�� CQ�n݃lQIH8Q�!�$��B�0��W|�x)�G�c�������'�@?f|YTCҀGS��y�d����@ �Q(�
F=@�mD�Y�4H�IR������I@�3n�`K�&�U#�11!�*D�P10-�%�p+Đ1���'D��! �d���˕�E*�A��.9D���^�DPf�zs	�W��HZW�9��{����v��5$d"�h����
e-$�H �IP��� ��o��=; �$�y��\�Kl�O�eЂԛ��M	�0=Q��	M�p5�� OV������y2'�)��᧡�T�t];�ś��y2����&�'�S�S�y�xi��$eِ�?t�\��D�O2�~��� �&'.H��� Ȏ]�t�Fy�Gr�� �=ϓ�:��9 D]�gU]q��$.�S��G�^,�LR@䆩�<Ɉ���J?�O�ț���'NHlȩI?r9�"O�9	�c��a6�A�}d2����	F��}̧!�>�
��$"���rDݗ�Z��ȓ`�����#��m��X���d����ȓ$�ّ�(�L!�XA�k�l���j�45 �(X�L#��#��B�5-���ȓ}�"834�S�Y%�(��
#(B�%�'���d�� zz\�o�-{�0J֧��}�!�$�l���AЧ��Z�<�g�üp!��ǉUO`��b���(q{ҥ�<fQ��F�4.��EA�؃�*��Rڠ�S!�yBK��8�L�SZ�9t���y�צ#�4�a%�ڬ`�@Y��	R����O ���
��=x�H��!��sG�F#a�}r��}��:_�\�c�MƳI���c����yr�A �h�h�)EdP�3��y�cZ1Ww&ɑ��6�|��Q��?i�{��nӮ��'c=|b+��s��x��a��mtq���n̓Q��a���I�9"c؝<���ȓZU~��U%
�Fx�y���~D1$��oG���O4$a�/�(�0ݳ�I7lw�#�'�ȗ��?y�\� ���2^����y�oL��p��� ���Ac�,�
J���խ!D�c!2T���3ȇ2E�\2l?�D�>)	�X��p�H���峓�B;�l�G~�S�!O�d�&!�3���0J��wX���>y��Éb����ߺ�bO�h�'���-�'D
���1Pn���Q�4�}���vС���L�VYãC�XԆ�c�FA�%)�JI��*U&iG~��p�6L�V!Ƈ��J �չM҆9�ȓ*��-�thQ1'N�s��!H�D�ȓ*Xl�({�r���@ӳV�Y�ȓp�r����I4�em��U�Μ��;:�aa!��Bv ��!��H��(0�*dĜ�i 0!��5Y&f\��B�(��A��$̀�d]-{G�P�ȓp�-�7DƱL�`(�RO��[F�D��,����	�Bzd��A�.��,��jOjT���Q/%h���jؔ	�$�ȓ�p @�GM����C�)֫�zt�ȓg�$��0+LE��c���O�t�ȓ�Ȼv�5��S-M
\z�Ԅ�f��8v�����ꀃc��ȓP� ��f�/�}����4�����bޜ@f�!h��d���$��o�\�Ö�̾9͜��A�C&6-�ȓ:Bz��'lF�j��g�> ���0�h�$�Y�v�"����X���$�ȓ��qǥ��@4�U�E��m�i��lxj�0=��b�� 0P�ȓ: *��g%I�C�̐ �OXc�@�ȓ?�I�fN���V��N?w~m��{�K�e���:&��[0`6D��a�懅*�[�@�.�^�0��(D�"��
E�(����+�d)�0E%D�����;")<Ik壀=uP5�$D�l!v�L�i�u��ꞔ\61Sg"D�hȕ��2�a�d�1���ӓ�3D�TTNE9���@b�$z�M`��%D�0��ę�DlJ����A?WT�Жi$D����S�r�
J֮Ѧ �L�­ D�� |آ�ݫnJ��� (�0%�d"O^�;��9rr��E�;�z� �"OBݛv�4�VQw��[�й��"O�;�k��F�
���>?�d��r"O��z�Ɲ�Hn�x��Q���2�'`��'B�'�R�'���'��'y�@a�Oҍ2��U9��ɏw�B��S�'���'���'9��'�r�'���'Ϫ����] �BDJ�E1nq:��"�'[��'G��'��'"�'���'H�=��)J�T�(c�J��=�諴�'���'�B�'���'��'0B�'��h�I^�P��ID��W^�:��'h��'f��'O��'�"�'���'���ÅM����t#��>pS�t��'���'���'���'b"�'9��'��A0��ɞhIl@c��� �6}�2�'b�'�B�'�R�',��'��'Ul�`�,Njs'�3��\���'���'\��'�B�'	2�'#��'*\�!g�������G;��`�'�R�'V��'�B�'k��'�"�'��b$c�8T�*�ô�'U�~���'<��'���'���'l"�'�"�';����o
heX�#9?����'F��'���'���'d��'UR�'ˮ����!j����甅�LH��'�r�'R�'>2�'u��'��'�E�4:��9V�]7�����eF9�?��?i��?����?y������'�%u�Jq�UC*��f/��ʓ�?I,O1����M�o��j��Q�q�߈k�`Y��(	�^8�'�x7�'�i>����M)Q�D�7ÄB�i��(����M��M��q�`EX��k~��̈́b�X|����?��S�gO o�-��Y�o	1O��Ĺ<����V���ơ�!�qx�M�w�ިm�R�0b�t����yg@)BZ&��� ��`ɜ�[d`�O@7mf����'�����,�<A��M@�!BO��H<���VE��<	� �������.�hO�)�O���!���t�˥@S�L����6O�˓��wԛ�H^!��'=hɣUI)-�Ɛ�'l)V0�����ty��'b�v=O��*&Z5I�
�i�h�����9�5�'Ȕ�{�Q�/@"鲊�D(�D*%�R�'�V�" �(`��Qc��	3*P��@2]�D�'Q��9O\Lc�m��yޞ��_�z�8��p=O��n�?;��/����4�#�IX�Q8���G{$8���O���`��DD� Ͳ�#g��d���%0��)w��S�H�I&�?�"�����K��E{�Os��o�SK�����O�����F4*
��h��F�O��'��V�a��/KǴ�p�@�.��ܻvG[Kyr�'��F5O^���I�O�`�7��c
�,�"ьx�Z�Sci�9�<�]��g��.H�Y�dɱhw�]��Ip�h��hɄ�����#_�p��vyX�t%��b�4nG�H�=�|h �I-�#`@ɐW�0)�>����4����O�7��O6p��-���(&lձNFL�)��08���5O*��1KN0B"�G����6x�1j���e.��_`] 欏(X����?�-Ob�S�O,Μ!t���uG��AP�b��\̓3���j	������%�����40��pj�ڶl�@e��.�<+O�7��Ǧ��Ic�
�b�a�d�e?ԥ�
ħE�\$�䌐�.5��y5��;r�Hl¥�%��|*,O|�K�X��7�@�Xj� ð�̦b_�5��J�!!�
;��Y�t��G^	��26�6��c������iyB�']��4OH����[*l/⤺��a���qł M^�� 8lq4J�A7?)��[��\I�&�.��;8w�E��bf��	o6�ɇ��";��m��t�QꎽLh-8�+�k��=�1�'����|�p��O��oڒ{{�kOԦj�lJt��gbJ,�ߴbΛ�ʣQ���O�9��j\6Zc52A@�<�S�ǿGS\�G��K��-J2�[�L"wD:w(Ԋާ2�Q��)l{P����W��͊��s���n�
� ��� HC�I8�4�@C�}�	ё���]��D�2��%,,�,i�d�$%�t��'��| 8R�ϗ\[�<�2ͅ�sV@Ѫ� �,?��)tf�.1�h[���`h�s�ʠi� �z��X6!1vI��<nU����ҩٶ���1S��q���ͶE�Pm:P�]<5�S��2rm����8?�:���,0���+��:��u�K�6�*6-�Or���O���E����d��>�Z��p��%h������M�P��?A��?�����O�2KŰ=�����5)�V�H��3p7-�Oh�2�,���?�-O
�$��ȱ�f��n��GC5|(j�%dK���'�
a�֋4�i�O����O��b����l���'�>L�E3���㦽�I#�z\�'[�'�?9N>a�KO��]�B�*;0��'�ٙ?��	���%rw� ?	���?	���?��q�T[h��F��X��m�!X~��ᅶ���O��$�OR�O���O��ڇN� �����%\�*J�����*�0�����ğt��ڟ��I�E
u�	�~�$�`2�=(��s��=�"��޴�?����?!N>���?�0I��O%R�o�C�<i��)D�G6l`������?���?9��?qC ��I�OTy�#,��@yVЋ�����ȨZ�������N�	џ��	 +`	�e�"�$I�`�h��`@��#I�!��Mכ��'Sb�' �J���П���?Eki@�?�u����=IsԴ[��G��ē�?a�F��q(�]�S�� ̐���_�47��@��Ɩe�8���i^�I?']�d�ܴ?��ڟ$�S�����bQ U���ў&oN�;1
.�F�'B�
��O��eK��S:Z h}sv�H 1LY`!�i*13��'�b�')��O���؟��	��h��gZ�#���rq-ՙ��yk�4�|����S�O�BF\�jr�5w�r�a��I'bN7��O����O��{V �<1��?y���~�NH�%�X}f���=��'��b�|��'���'=8��@Kct��@6tZ
�r��o���$� nʓ�?)��?�H>��X����X�j�y0ˈ�oD���'�3��'�������	��`�'�z]J&�Yg�Դ��-/Bx�ڤ�M1cq�������D%����dR4*«�����$;��)P$ޏ@}"�&��Iş(��Ny��<�	T���zi�okR@p�nG�2ś��'���'��'���'0I�D�O�@*�Άi=�D��*[�ߢ$�QR����矠�INyb��/��Sϟ k�U�(҄ {`O¥&>�a���4�M#����?)�$�푌{��*�@��4O
6s�֡����MS��?�.O�h�|����?!�'dU������y\@1�-8�zQ��xr�';�Ō j5�O���Yh֧����f� �J6m�<�uŷ�?����?����-OkL�AЊ<�0iL4�R����$r�6�'�	?5��O����0r�MIޘ�7���{eQ"�iB��:��'�2�'Ob�O����,�ɝc&��kɤE�j��Ύ/cD��޴p�4h������OZ�y"d١Mm\����	x!�c%A�I���,�	�+�:ė'���'E�O�y���7:���`�_�sE�+&�d�z���O&�d�O��Dȿ J��k֦L&�;$ƽ	���n��|�g���O<�'�?�����Y*�8qf� �P����:�<l�ܟ(�Sgɟ�'qr�'8�[�|J�N�l˴xA� 44YL�K�I�x_�t�N<!���?������O\���� �4p`�0X�

�Y���pFm���'g��'��_�(��l[���*�/�������:%������O����OV˓�?q��w��0�^ޠ
v���1��Er�L�#n&���^���	ɟ��'�R��&Oo��0�@fO�?X�{�f_A�:�Q�B��MÎ��'�f�e��xO<�T�F9�=�f��h���R馑�Izy�'$z�SPS>���ٟ@�s��)¥�5O�h1��bJ&�B���?�$�O���jF)J�T?�y≙yI�P��F�%��	 *�>A�V.*���?����?��������`�D9;���Ғb綀St�i�r�'7��cq�����O~0�g�ȽI P��O�[>�s�4q��-q��i���'���O�6O�遽%z|͸��1f,�!a�[� YlZ����Ο��I�����G�$_>��᎐!4hA��:+�ҤC��M���?!��EzH )O�\����3gF�A���Vh����D��w���FxA!���OJ�D�O̜0Œ�c�D�s�o�v�`&)Q��I��9{.P�*J<ͧ�?����(dx�H+�O#E��ؠ&�_x o�Xy��'��i>��	by��'Ԕ�JU��Y�!�aF�?v�bA�Z6S������IY���?!�k�<���e�=H��� �ߚ>I���j���%�<)����$�O�E��F�?�H�]�F���EQ4U����s.s�����O2��	Ɵ\z��3��6��t�B�׏ϫk{V4Òc7M��'�bQ���	�r@Y�O�Ҏޚ=��E+��*���PQOÆӶ7�3����|�Ɍd����:�$�)I��9˲KX.K_*L�Go�Uz���'rY��`���ħ�?Q����&f���kR�O�V�K�E�%�'���'���A�'��O/�\c���Zd��<R�	��J�u1���4��U�xf�oZ�����O �i�z~b���l[4종'�/���V���M���?�� ��?	��$�Ol�sӞ$Z1j��0D>t��I��iň��0�~Ӭ�$�O��$ퟖ�'���Q&@<�����i��`�r��޴v1�����?���?����򙟈��~v��!@@�x*@�C�H8�M����?q��7�-I��x�O.��'<�ep��G5���bDK��?��P�jr� ���Oj�䋧"8M���d�O��DE�.ܖ,b��5_?@�JS`X!K�ܨmҟd����|���?.O�,
䏑�l�X�I�/R�rp�'��٦5�I9)�0���Dy��'���'�	���zҍY�m����Ո| �"��ē�?��?�-OL�d�O���s@�>Ĩԩ3�Ƈd��dc��?2(�$�<i��?q.On�$[��r��<M�t�BA������7��O��2�I՟D��7.J��àlӞ<���?�ԭ"��bL�f�x��'D�	������TY��'�<0��Q�7\�#1��)�9�o�~�D���t��$+KXOġ�c��u�fYL�>|�n\ �iB��'���'y6:�~���D�O������󕯟�d����'�#�j��C�ۦ���LyB�'g���O7_��s��	ƭ" ��y#���#G����E�i��'�4� ep����O����P�I�O|pKƏ(@�h�ӳ��&y���)�@}R3O���F�'X✟��:��Nſ>�(P��W"*���̬�M� p���'���'����OH"�'�r,C�p�2� ��;X�� �N
�a^6� 92���O��$�K������'�2� �88Ǳ"j��*ѧ�*w}\��i!��'.�Ju�x7�Ov���O��$�O�n�y�$�WnӚfx��+�� �J�v�'�剛E��)���?���y�ޅ
��f��"1��x;��i��H�]ܠ6�O���O���T���O�@@��
#�%)��HB��cqQ�h#��g���˟��I��������	�Gl��&@E(M��ĺ��@&
�؉	S"6�M���?����?A�]?�'�k�h̄�x����L�"l@Un����t�'
B�'���'���'���6��H��hxqBA �X%+�}���l����	�D�	ޟ��'�b��,���G�X�`�k�NӻF��-'��O ���?���?	��?y��� ��6�'	B	��_̈1�S�9Q���Gڒ0ƾ7��O���O
˓�?Y�(Y�|
L��Q6�]�����g��95]P��*d����O����Oj�Ql����	ߟ\�I�?�`�%�d�h(��*� ��ZSf7M�O���?!�b��|
O>��-��� ���$yC�PK �u��D�O"��~��6-�O�$�O��	���D�s���ۓj���NВ� ��wN>U�'����"0���'k�i>%����#"O���bS/U9s^�8�Ѹinl�2IcӘ���Ob�d�����O0��O��פ>�@�0�=�|�2�QĦ�c������Vy�O�O����,8��bQ�Q�AFF�6M�O���Ox����WU}�\�t�Ik?9"dA5`� �ʝ4R�F8K7��˦�I��<�	�	���)���?!��`��W���zM���@m.�Ñ�i��7-�O��D�O`�D�u��O (��#�3p=��M
 ��FX��;u�l��	������IQ���E�Rv0�aFK��
��"���R��Q�hc�j���O����O<m�O���㟼؆�RM��і�˵y�� !�� lWDc���Iҟ���۟X�	�-d��޴\�Z�cઑ�cE�]�ք��y�b�:�i���'�2�'RP���	�>���s:c���`�x�~4
r*�d��듘?A��?	��?yA�Ϳ4<�f�'���ʍ�`q�����f%���)E�[�J7��O����O���?����|2���~�Q=tlB��@ݔ�q� ��'�M����?����?7�ۡ���'ZR�'��T�f���dh����H��������4�?i)O��$I���O&��|n�*���U��n	D �T���0&�6m�O(���q���l�ܟ��	ǟ@��?��I5,��d���0�jd3%&�6vbҵ�O��$K3��$�O0��|�N?]A"F|Qkթz��a��/oӲ��[��lZ����I����S�?��	ԟ��	�to��:b���*�KW+:ҬUЦln�Ls�M�O`��<�'���?au�Wx~41�1�]ٶ	R�_�e���'4��'��2r�,�D�O��亟Ԙ!�ڎ$&����p����}�,�O��"�'{�S͟X��؟L�V�\�,m�{�B��~G��`�hƒ�M���_��P�x��'���|Zc���`�Ɯ&,���kԒ_f�m+�Ot� �2O���?��?y*On���b��)$�u�V��8�$�B��E �&�T�Iԟ�'�P�	ԟÒ�d���d����SP��2w��4�	Yy��'�r�'e�<��h�ObxZ��.4����w,�5���ʫO~�$�O��O|��O�:&?O8�ЗJ��I���h���m-.m�c��u}R�'��'��	ju{O|ʡ��j45����|�����<{����'(�'���'C]��}R������ѳh@Byó,�M���?q.O:���C���t���DbEKG�\�f�p��K�A����L<���?yv��?aM>�O�$P{"!��J�N�����B$��yݴ����T��n������O��Ca~�*�5�����.=d	4�͠�M���?��<	L>�~�!��-�΅��ܐ5A�A3����I��@�M����?���B�x��'WD�)��(p��D=wd]�1�'. �w�'�ɧ�
�d�#o&��Ĉ�8���*RIG~
Ln����ٟ�;�-N?���?����~bė�4��P(��BʰHF O��M#K>���Ȗ7��O��'Gr&�mU����ـ_*���)��%��6��O8-XK�[�	՟���p�i����آ!��I9&�J'7ْP��>	��8�?�.OP�d�O����<�u HS�%hT��4kdA(0���,FP�1 �x"�'8b�|2�'9raq�R��LƂ-��$rD&�#i?~��'��Iԟ�����4�' � �v�g>Y��,[91Iz�ਓ�Qq`!F�>A���hO����$n���$^6*
~��A	�.&x���G�ZYl�ϟ��I�� �	ky����:�k�Q��%��wdLK�k�9��Iܟ�#$@�����\���/��MȇC�< �v9SM�צ1���������e�d�d�'�2�O�~y�պТ��ũ/�
�s���m��O����O���PL�1+1O��>Xq:��� ���:���O�7�O����g�pUn��������(��?��i��@�)D" n�ٷ�[�~�$�
s�9�䅾۠���p��Z�*�~]��$�(������䛆�;LB�'8��'<���'�S>uQFBٗqۢd#&h�	v��a��:�Mc�C�;���<E���'B�ᥡ�%8ݘD�J��@�����y����OR��_�1��� ���O���,��IS��K�j�8�q6��2ƒ0��yB�ʂ49l�h�$�O0��2���ǎ��t��5�!��Dn����󒆜��ē�?Y����S`"�T�D�s��Έ���(�U}�k��'���'s�	ޟ��� �P~�`� [�vq����������O����O�O����O����ʷys�e!'�ӧd���@�JJR�`�����	����{y�J`��@�x`#��e� Q��O)UJ��?	����?��7����'f"u��9f�p����0	:qx�O����O����<���:�O�ĉs�KԀ>���ju�[4+֠���bӾ�$6�d�O��d�7}�O���G�s�L�U��#?ST�s�iO2�'��I�I/��K|����:�ݚ)����c�6(P�ը<�'��'���T?á�4?u��k��iT\�S��f�V�p�t[ղi�n꧹?���).���e+��ІϷ$�����M&MV 6M�O��䓜2Z�b?=�K@;!�4�ed��hܸ��.}�����ۦM������I�?�xK<i�@T�Qw,�)@�hke*A�v`xm�i�v�ڊ����t;6���V0�Y�q➼L�"��!�L�M���?���kZz��4�x�O�"�O� J!�Q�礕�H@=t
)G�i"S�����2��9O����)�Y_\m*�I�4\ ч`~L���FE	6��2c(�(�a�e ��i�Eq&�Gc�
2*��s��@K䡆�J:�L���А}���D�	��L��+R>?�Y��M�Q�0A a�˛r�Z�@���.�LQ���ʂ�W)WgP9/L��X6&�V�y����|��0�r�/oI�P!��dxb��F�ɫ56,�W���j�&9v���h��Hq�`O�A� %�D_������Y�tf�gf�*��O���ܡ{j����O���&���^SD@�m	w���k��ހ��d�<�Ҍ{�c�3/=џtB� �j2 *0nG�F���iADX04�@��ؐ/�P�F����b�F2!؞�?q�i>���jyp�DĠ+'���,Q�V�4p��?	�����~m��k;^_�d��|o�p+�O��lZ�LPc����}$ ^(G����JyB��"i�6=�\�Ģ|��Ĕ��?��k]�/�H3�8<�,zW���?Y�{��P���̪@sz�1MQ�H*���'[�X|�c�66*����$�n����O�H����)"�$ّw�P��4�碈�R��O��}s�!E fʨ���`�#�thN�Lsw��OX��0ڧ�?)�o=Δ� e�^�A@�E�Lk�<�'/&=O�5���5UXD`�!O^����ě�	6,E��ܵzr&i�T�^�4w��o�埄�����x�,exv�������͟�]�E�&� -S�II����a֛ �(i�h[�����"fw�pS�K�'��e���F녉:�h���0�>�[2�̙\Ն<�����Z���i�'�M�(^�<���U�,��	l3�pR��.�?��Oh�������	1֖��FJ�).utݒ���?9�C�I/r�TMX�j��E�$-H�bˆ�W摞�ğd�'@fp@�j�ÃZ��N��)�/|w�]8��'��'��$f݁�	�� �'O�(�d@
�<?�c��4 ��p(Mih h���C��ܚ�߸��O��RmC3�L9��	���d��)7��4ӁL�
O�Jd;��u��7-�QTQ�p0E��/k�aZ���.Z�����LC���$#�Oj�9�㗀And�c#P�o�t�6"Of���4�,W��~� $�Ĉ���$���u������OF�2Gm�->xU�C@1q��\`�%�Of�W�	��D�O���L�e���(a�f�i�G�G���`ܐ��`k�jޤ��a�J��M��$�@�'���H�4~_�) �Q/?��2
�$p��	�{��Y�.�Ǜƣ͵�(O�P��'��6mGz}rΩ��*�O\?a�L����'t��'4���i�?��Ua��F�!��J�'�z6�||�P`�9 XDݪШ'�(��<�P/�>1�v���l�|���W	M��hE9�yx���$��mУ�72�B�'딠2jԎ#�}� n��ҝm�|�*�6-"!��ga�0��C�(^�c�>q0�� $q>  1FB:wJ�d��l���($?Ua��]�$�<��IQ3#��T#��0}���"�?�q�i�^6-�O6�?M�qȄV�}ѦH�,�.P�b���lx� �r��]�0aI'�O�v<x�srf9O�Ez2E�?��p ��ʞI���8%I��~iV6��O��D�O���_"rh�d�O����O���F}���0��\��]�e+ZɈT����"���	m�x���&�3��uF]��
>R��Yq�,�}z$, Q���#�$\�޴
�v1��'�3�d� v�2�t*q�5�*{*��$6?��k���>�D�O���K7[�$`�u�(jb��iE@�-~�B㉴nr�i����^	�� b札\n�~B���'�򄖮��9W ���4Y�7A���8��@�D����O����O��;�?�����+k�Yiw��?]��R)��[�1��!�D�Z6�G�n����˨=d(���[�*�\�@%�p�@q{wǈ�.�bQo�)�@��]0=�Q�Tѻ�ʆ	���9��O��mڄ���?�����'��	b��M�oȲu�D�F�be2e�
�'y���s�-u�D����0_���y2Kn�F���<y��Z�Ds��'`�O�*��)�����4�%*��\���'N p�a�'��<�>���,���O)�J5n:� � ��/6P�\�`�+j�de���'���pgJ�)�@�gǌ�s����"+b��0�F��L@��p<�aC�$����Ɂ	��P`��� ʘy�@@��'fR���'=�U2B�D��l	��(gBxC�	��M�%)ߵ�H��%�y���:���<y-Oa���ʎpDf��O��'m%������tA�e��8(7�د\V�m���?�6��N^V5�feԖ)�>T�
A���	�|:�LS�MD�ڥg[)�H��EO�U�$�-6+�-{&�"+b\�CF�i��~!3��]��S�N�tŋ݌��	�e����Φ�I�4�?��tD���DL��̍iuXp�B����'b�'O��u@B�a���+[ހ��|����Q���`���W9��@����M���?���/�0H"D���?Q���?y���Sn�l����雴
� �p!ʔ=�4h��k��yﾙ���E)<dJ�Y��d�x�'��Y��� ցY���'��> /JL9��H�sf����� I�~<����>}�Sj�<@P�#f}D��&ȓ.-�$7�Qy�E5�?�}��Ɵ �	/2����!h�e��������ƓL��ˢ#ױOx"0���0 4F4�'`#=��'�?	(O条���p��y����K��1�j6�x�Q��O��d�Of�Vɺ���?�O"
����6���1��7@=�x�eS�s�J- @�8)�����RX��LYY�'�F-P�Ú�a�4� �
��E�ˏ@���C/�*N�0@�#�uPh	D�N�ޣ<���2b�A���0�$
X�F���	�M4�x�'"��Vy�j�	5���qNl�3��ZX!�Dٚ|��RiQcR�2�h[�nK1O�im���З'�H�Q�'���'���#V�T qP\t���=sL��!�'�B��K���'�B��@� Y!'�^!���'�����ȍb��emݽ8:@HǓV���$P�F�
���̹T��\�u���Q{"i�r�F����:OD剔�'��ʹ>Y�K7U��)Վ�� 6�	�JV�<y���?���O	�'�ԵqV'_!l��P�T��*\
���'}�7��Ъ��#%*��{RK�).(.�mZdy�M�rL7��O��|�IF	�?����bݐyZ���
� PU���?)�����S
 f#iA1���{�D�k�+�0���-���`G��yo^@� �	)1���Ӑ>��!�!R"l��e��br�@Y�IC�Z�Px��+�G
[p�ɹS�B>s�Z���(�h��X�|���qӀ�oZ���╮��YDV`9P�q�bL�Cd_���'���'6���4��0Z�(	7
�Õ"',O8Ez�MӹV�6�Svl� ^:��iTGT	&�6�k��'���'���B�%�%P���'Z��'�4��+!�K���TZ؂���Ƹ8�F׫];��6�i��U�eט��v�¹ #m��Y�@U E�S3�~�h�kҐ���v)[f<<�POVܧ*��NaJ�q�͐t�f82��s,ʼ����l����?A��0�A��ӊw�&��fʆp�,���'��Y�u)�<c : �!gٲ���O��Gzʟ��2�X;2�y*I��^7xiDE�!B^�5�����?9���?y"��x���O��S�N��L�����b,�" C��@���M�G�0(��-"�a�A-I]4�7�ɯG���ЦE����ҍǛ��ABť�j���a.��(��P=c=BHC�	08�ݝO6Ȓ��9J�9R6i�O`�m��M�������O��p�G�O�.A��� �8)a��.D�������b=yW�h�6	�3B.扪�6�I~yK	�p�\�'�?AC���g�85)��͍r�!�F����?���p��H���?��O���pT���C�\-�U��)�ܐy��߆0��E���۵��r�R�Cm"�y�퉢Gc��u�
>c����T|�ӂ���>�'GÀY~2�X��"��@E{r�$�?��iwp�\-�}"@F��U�E� �K{&��<)����<1t��n�]⤭�oC����o<Ƀ�i�<�0�`��j�L��-��fņ��e�'n�I�>��	۴�?����)�0h����.G$�|v+I5R%�\"/A���O�tzb\�G���Ab�gV����t�T^>Uc��<:2f��*^��0��"}��g�Ω+"�Ҝ@���r)ʧ&���H�n�jF����D�"���O҄B��'�46�Q`�F��(k��B�,��e��FP���b�,�Ipx�(���M�*��dJ��Am(O�Ez��E&�IQ���yw��P�\��X6�O,���O�T�Ń��{��$�O.���O�٭+�TI��Ɏ� I!
�!=LE��O��8x9����m2'9�#�z�a�1OF��mR�{+���X���;b��,��%��@�7���5�
&#xq�x5"^
�y"L���ʡc��1~�\�*�������(U��Oq�2�'���R�;�>���q��4C��}ѡ��\7r-����Q,n͆M��gK���	�HO�I�O��fF.I	'��@��E�韙\�J����
5��Y��?!���?17�����O��QG���'ȼV�V-���t\��G��L;\je(ODܹ34G+OT��
� �Y�7h��`p��8Tŝ�m��e�An�5L���E���~0:���4O�i5i$4 ��U��d��j�BZ,x���'��'��'��O`ћ�"�8s� ���J�Z��@�"O���D��.]���KT6*��9��ɦ)��x�I��'1�*�QO\q��i� � D@T��ȓ�huA��
%�
����l2`̇ȓ8�j��,I��x9�.�9P@�ȓp.��;�c^`'L�x4J�qw��ȓX0��E�S�!@�l�f��lJ !��R,������/��{PBƮ$�����*
�e��B�H�.S��-G��I�ȓ;8�sEC!d�~�7�� �x����r|���ىK���jtH#�J=��[�`���c]�3TJy���~��d��K�D�#D�Dpl��a�$K0�����h�$&d<1�CK+T���U�p�v1k�X$��a��BĄ�ȓ���%��:��*]ͅ�h�<�ژqpF8(��T�`�����b�<�ahԅc�2q�q�U5'�h���Ib�<���@�p�lpx�N	�)Uv��V�Pe�<Y�J,VG�x�$EF|v��ee\a�<9�),��C�!Y+N��U��]�<qVk�#�a�U�ʊL/�1��@c�<�a�Ӣ&ƀ0cJ�D�9y ��t�<�7!Þyl���l��|Z���n�f�<4X�bSx�ꉶ#dE��G�g�<9 �I,��Y��R3�,���^b�<I� ��~�J�z�W����+XH�<i��" 
��EB+	�Ƚ����D�<���۸@͘D��V1@�Q ��J�<�sϗ�?�1���E8Ta:���I�<�q�W5>���ӥQJ��Y#�Fx���׭wy�	׉U,|�j��l؎ `0��,}VX�'"O��@BH�"�����-(7���x2��/�n�d��"VG9��>����e�"�������?�d� ���p Bj��d �T��, ^O8���4�ʓED��_}�$	�����)�P�m#N �+�%��^����'�2�aNS��|�����Dz�x�c��zz���,� �e�[������ڢ7i����'P��H��Mx��;��g>�Ax ��%�m�A�c��1v�	��hB=�~�ˉ/,����G����<4��E�RFJ!��;S����G�@X�P���E+����\���FBۚ��r0��<1V�
)-�bAB���(��S�S#A�Ì��x0`�bjח�y	5�ɀ��b+.\�����V���I�e� ��Յ��/��q�5G�w��x�?A�o�)���n,d}��C�y���-7|%K��]�>RT� ��6햍 !�IV�ҥ
J�PH �����O���[>E`�L3�P�b�J#"Ѩ�Q$6JD0�%�hv��0*�
>�?	�#��|���qD \M��壔�P�@�����OC��$�J<�(O��'����r�8Z��`fJ��-���ؿkH��Dɴv�tC��ΗC�%Z�@@�����g�� �{ЈN�E�T�'��y���o"���#�,jo�u���ܒS,�P��HO�Թ�D�sZ�q	Af�	J�@*��H�_AdP)��ʉJ��c���W.�1s�]���J�,����']J��N?�p�Ȟ�o��Y230iHC'%Q�2b��ѳ	�FnI���㠂G� Lp1x2�M�~�faД�^8
"��<��b)!�`�rC�@�Z��Xџ���k�d��E0xڀ��j(�rCF����-O��TH",ډ/3^y+3lDK�8�d�K� ʲ��6��|&���*�����śˮ�#�$~����K�>ݼX�ד"q���֧^�.��)E���H��h0��}[���F��ؘ$�����i϶���O=i�a�De*�\(�A��O�hQ��nKPh2�JH�@iႯ��)���(_7n�j�į߁I�.��I��t�R�V�~r�ƴ9ۉO|���Q����a�,F�(�@��\�%�l��H�>��! ko�-m$��X�4@r!����]/^n"L�wn��1����T��{��.�$=g�x�=��p��	/� �A� Wȭ��T0[��� %I� 2�r1��(Tp^%���i[�(`���|��I؃t<����yR��Yax���;��"E�L���!�Ǧa��tR�r~B@�C���=�g�I*~Xض���O�!pi�Z�|D~�*єy,4z�Ѡ;��X1�*�� ���	�q�&��u���M�T���D���~�R_>	7�Mx�d��� A|�PD`P�*���H%Kf��<q��l�"|c,��R
�SM�"��V��oK����+ad�9�a�C~�	!��'^�YW/\OܓZ���ǌT:]b� �̂P ���ɼ<LH�	"{q�H�	�L��=��((�H�ˡ	rx��"(O�?��	����jA�	���L4Tz��Ȥ���QkNơ%���B���jX�=a�LW�8T��u`�<�$"W���} ҩTp��:6lT&�HO28�#]�u>��'8��O~�X��*�bu!2���= 1�О>�FlX)�z`���<��|�Ԛe�t�Y�n�< ��`�˪Y��d�۴z����O�ׅ��d�7F'�ۊ@��L�vI�N�r� t(��FhɰaGqy�
 �$�=�\�ɉ{�	�� ���'͕�B��9f�0*ڴw�~�'�0bPb�'U��@$a�+Ḫ4�D�J�$�p"R��+�ƽ���Z�
��uE{�-�C��]�c ^��D�^s�)k`nC;:@�;�U�p?y!JYM2�PZ���v��yysM���HO<��$�Y�(,@�O�]ѮO�����^5�)Y������'�'��([����Za�#Lد@(&8`���Q�����g_JT�i�l�#���*TtU�O��O�<�fh@�*¤�Es�,(��R����$%�j`Y(OHHp$f�~���<s�
�{��DB ���R��$��@��Y�
F$%D		o%X��dz1Ol�z��:�L!��
 \t���Ɇ�W!������0r����{*���JQ/cޕ�Rጵ}�����xɂ��Cj�<9f����?	���?�c�f�W�4DcFٱ>�|��A̓~/}��!f�,rABS&4���?�	)c�<,�aB04wJ 3�+�84�=�+O&Aw�39�0�Gk	#w<�����.Yl��*��OU��k� :�����m r��PM�O��3��?��l�)vIT}��A��гG�O�T,�G�B<A&�4Y`�M2����=���V2l�$k�[]��!JW̓_U��a�J�=bH�!��Gٟ�I~���Wg��qBƐ���!�| ��{q.�<g�X�%�!�|"&R��y*�p���cf� K�ʽbu@-y�"pI'
�;bNp������"���O�����0�%�pm�� ���rѪ���0!��yҢ��F"0 ���O2JWF�
�"�ט'h
�᳎�5�V!C��p�:���?zc���b0 ��A�a`��3�|׋@ Mxb����)/uG`<p�	Y�9\l!��юRR�Ps�#g������q�1O���G��u�͘�%1�NȘ��	�� l)����������'�eж�~�L7�dM�}�'��r�"�9��'Mأ	,U �y�M١<u@�A/ ����>R�<x��B%@9�p ͤ&�:U袩r3��cH�6c��Mh��C�nZa#3�LQ�S��π�-F�ōV X)n n0��*A'<ɲ��Q
)A:�c�OU�$
�[- �PX.�S%8�����R��ID	�O�0�jP.G޸b�0 �b@^��+�Z�d���g;扃4�и�p�~6�����~=�
U��k:���/?ji��$��������O�PIG����d랮�=��Q�p�v��`S6���&�3
tsgW�Θ'B�TI�c^�j�>9y�珌E�*�K��-PF0z�-��6�|����$|�� QiC?A�c����>�
{d�
�. u2�O��
��<qK�9Ú��2C�
����Icy�ӵ��?�1EB�	��9���]dh��*�_�$U���J�CJ
��A�T>�(��E��3CcH�j�zd��*ΛV3|���P6|���N����I�\h�D0G�):g��+̑S�����,ܽ|��!9�)НJ�1O� ;�!��
&�;��lO�����Q�DL�i��ύ <"n��R1G��	B臔\�L(����2db�P�`~I�aÔX��,A�B��$�&7�X��擈f���듥�"ap7�e�AT�U���<IuE]�2XԊ�P5� �k�6v�.�'�����i#��Οla�'Ѭ��@�_;	�v��^>c���U��{���a/M�'�t�'�#�I�VhT���ʚ|��8��L�O�uz�_���� ,it�{& S�m�V+ՠ�����NW�'�2�=�`�UAJ4�e"TżSu'g
��8�
�y�E\q?�`0�������ɿ�TdRq�鴟d�vAY�)���Yu�C�	BZ�; 蝲Ș'�Z�9$�������vǝ�>U��yRG�*E�E	��D]&<[�O�n�(dJa�KT�[��}�I*{���Z��ϒn����2AZ���H�D�h [�E�XE()��ɽ,��B���UX��b>��. axu�T�\M8	Q ���+�m�����6=f�r�O�n�����Vy��ڹm��xg��j���Ƿt�Z��S6s�!�g�|ZR�1Jo�O��#9��$��<�dF%���ԯV�e���C3��4a�f�R�Q�'���dŗ=�F���wjNA�ԃ4XSVQ���ȅD���S)O`L[Ai�O�A�F��$ʓMϊ]�OV�a�@ޒ=E(�P�iߋ��c5���.5���b3Dr��+F!��{^��,���[?9mpݡED�`�@& �X�����<��
� �u�O�� ��.�MC��Ȥ�A��X�	Z�ϚS�Խi�H�3�	��X�O��O���$��.��g��Z�^�df� d�΍����{����I?�rf\>���|�<)�Ś'�rpH��ܐ_\�5*�N�x}��S2e�����4���fŜs�$H��Γ`*V�r�Õm��P��K�x��j*�\�2'=��n�vm��w(��ř�%�J]yҀ[6��[ ��9nۜ8XV�$}�H��?�ɵg�d�EǍ��~bi�;$D�aUn�UM��u��Dz�ǖ�mn�3\��?e���p���z��!����"T&��MZ��O"p1�h��D�U�Ku� *вd^/T��˱7��p1��iږ���!=C�a�O��O��[����M���:�
C���21���G����T�#�ę �=^h���z0
AYKqO�x#����~�jU#j�qk�X�l�¥w^��1ߴ���<���<5�]���^�~m)�P�}��)�WK�5OQꡨ!��T�'���w r��ڰ��<�	�n��|R0)ID��M�m�7�~j�IB�	_�ܴ6�&�"���1 a9��"u�����`ޗ��'}��#� %�v*	4jf��I�H���5���Gb�9������4��y<ʓG����b�] ��SVR�p8�hұ	(ȴ[#�����C���}&���\�uB���G��z�Z�O��O���y�� �=N���+�A������(�h2��&=��8;��Q>;�8A�D�#�I��D�6H��n�r����C�����M>�I>�2@!�'"��P�v)T8S%Α���J��h!�f�/B�1Q�+�ȼ�>9���r�(�9�=�6<)wj�q�\�l7z�`��>�X���4��?7-ڄ#�^�X��؅Zh�%�@i�@���.�I�eP|1��jͯ#�jDB�A�P�OZY�����t�h@k�5,>�顯����K�X7���VVr]!�@]������j�ia-Ƿ>g�D��F���@�N�C����w�Zo�lE;��^*$n48p�|��|��m�
 S��XU��1�䃚��$ioZdb= 
�0|QQ��-[�4B"���D* (a�y��8Ҳtx�Å����(��h����ɇ���Oz�!V�ի���xTK�v.0 9�?"�\��$̮=TQ+g�
.m\A��T:��Ib�(��<UV�+�'��l�$���f�h��O(	�E:�I�<��G�C�*] ��&+����1�:@�օ*6�ɚMu��K�	�(� ք(2��%2P�1w[(��0�cjM-/$�yir����'V���t�^�c��ĺ�H��V�]fc�Q�oE�W��U�᪏�l�:Q��yxF�:��M�[&��$@�胳*ԋ(e*�r�O^(@�'����7GϞ�y0�ԂN�h��=K�Q3���G�N��4��T��LN�8Dx�~���\ƢEP��ؽ]j�nz����Xβe�ٟT�j���	��%����9eҸ�� �*���T�J�U8���&,�7���2
:q�c뒄�r�;�
G�y�(�@EB	�~6.HJ�'u8��Jͼ3������i�ĸ��O�'�=��,Y5u��I�hSj�sa�^Ƃuw�E�Y����]./����#��0<ɦ�\5~hrxzE坤\�H-;�*�!*�$lXb
�g2�8!�ӈ5� ɢ�EӤ1���9�+ Ȧy��ԨHڴ�4>Od$ �J��U��`���z�Bxy +�=X����"L�ڜ �>��U�\��;,H(o�`�{��Z��#�tI(f,A
%:H��[!��H'�ȱ,:$q �,F�-Nr�Q��Y���'����V?��v.TI��)_J3��X�,g��B�l�1�PaG}r��3s���&�z��#�`N�^bz�b+r����J8v�t;,O�L{@�.�s��C�ֶ�Ȫ0jֽq�d�rm	)w�a{2&��lڮ,#�f�-�*��h�a��,т鋒qlY�Ǆݏ�Y���)��L>Y���0i�		φ<�����1�\���^��sU]p�� ̀=<6�O<1d�-�.Iqu'X��?�U�2���Х�i���M�?����%��_rPJ�D��C	���:�F�<����"�	�&q� U H�ɶ��q��-p�20i���ei�dk}�Y>�\wj� �П���G#(�ʼqa�	_%ޡ��N]]1~5����;W�a|g�s\���!F�-AJR��Ǫʎ����rӇE�]k��e�ۿ6��	����^,j�q2���)�t̃GȡX�4L��ɔ�j�》�<2���@������Y��F���!�-t�ܰ��]y��I^<3�<9��-��v�ڵ�O�^7lC�Ƀx� P�%û+G2x�C�ȸA�RC�I-7��AR%X�wL�1^,zB��%;�68BsnQbf
4��*��chB�I�k�*I!UA%�Q����( C�9S��\j��݀4	�����]9g�C�:'�eC6����E1�LW>sXC�	�Y�����P5�\�!$36C�I�>Ĩ��_9Uޠlp	��V�C�L�D=i2����Y�F`X�!C�ɹN���(DL�?P�)��kѐx;B�IV�<㤅@	d@�ђ*`(B�	��f���*Q�6�\h�I:3s,B�ɯZL8�)$Af��r&�5z,&B�	)X\@�щ�00-tA f�3_K2B�I�1]�!KEH�;%ty+fi�`DB�ɄOɶ�)S�ҖrpZ%���q�(B䉲g�n�ѕG֦�F��ro	:7��C�	��z���W�[�0��O�1&�C�1"%8m�elQ'<e�@����kW C�I�T����`�
����""EK�n�"C�I�
��t{'�I������D� ��C�)� dI��G�}$������c�a��"O��3EG�kj�����vSf�BB"O�is�ɍ`��ZWn�?�5�t"Op�3�çAd�"�/�<z+Ĵ�"O���D�D�[:>���o�-Q�Hq"OxHH��b\���N_�xL�ˁ"Of�KS�Q�a����`]�f��� �"O2�$!]�C���r�� ��"Of\���� ��Ѫ�
U� #�"O0H2'�J5~�\U!���+B�8��"O�0���M�L�aΟ�7!j�{�"O�-`�� ,��x��\C{�	Y�"O��!p�P�#�X�9@�>^{AP "O��i(U1U�ԛ��-s�4iE"OX%@�K�1>����~_(a�q"Ox�ja�	P����C�
"{8��s"O���Ԩ�"�t,ZѡC�fz�3�"O �;�`A�!^Plв"Or���,[�uw���tff�eA�t�<	�ȝ#$�����tu�L�`�p�<a ,�[�h
���c�:�ȇ�h�<9T���A���R�Z90 ǌ]i�<���������?8�Ƙ[��OJ�<�! ->gF)�ǦI�J;.M[��D�<)�BY"'Rt<+B�Fn���q�~�<�!�O�g�Ҹc��=�ֹҗI�U�<��-=m�qX-]�shdr�j�e�<�dW 'T�p�Dl�8s�� r�h�<��hÅMZ����x��Re�<�&P�M���13fK�|bDHHʓ^�<�䦏#߸�(@B�E"��"C��<�#OM+t{n���Ҿ]��P�WgQq�<�r+��HϪx�B�(��	���w�<���°%��0A�$(�f����p�<Q�B�t�1WO��-��<�#Lk�<�d_�r&�8R/�������q�<����9iM�[f��b+8j��e�<)��Ѻ&+������y(L�C�d�<���_��w(K�Z�ie�d�<���͹Q���X�Ώ>���!@G�<I�˺�И)��|����vȑ{�<��I�7g��ʄ��-���lPr�<����u���"�	O7v�M�R�<�
@�OXЛ`C	Y6h�@�Q�<�u��)L$��4B�O��
1/�Q�<A&��#?�X<��տ ��r'��U�<Ab*�$@@�Xa�]=;SL\c�J�g�<�Un�ofy12C�6t����g�_�<�2h��QȄYt��4!�${��]A�'�ў�'C�v|	��;^�i#$�G,m�*`��S*t"�Ȋ�t+��+X��ȓTWx�;�l�$/���)�͘�RN���b.������������z�ԅ�HlD)@Q� �@ `$�Q����ȓ��%��\<XQX���HS9���ȓesb�0��&@�}bk�"tFu'�DF{��4i]	����+@8b���N��y���L <a�ՀWU�4�� _�y�ȟ�L0����/ɇ}�~(���yB�[�Dюu�5$?L_���c.�y�ʅ~�NP���ԱY�����6�y�{n�����0;.ARQ�V��y2" W" D�l9�� ����yr��f��q��JW2d<Ր�#
�y
� 
���Q�ap��]&:!��w�O��=E�aX�j��	'.����	�y2��m�L��5��&8�#ゎ'�y����v0���I '�`᳁Ț�yr��b�� ����Y�M@�Ê��y�H�m+���.�q�D����yB�D ���
��1g܈D�1��y�CۥD`���Ո�fn�h� $P��y�i�O��l�DAȼY
�z����yb��%>��bu�i��vkݕ�y����*v����l�?-��{F�ƻ�y�M�vqJ�aF�f�C��yb�T�R��K'N]2|Z�6����ē�hO����A�R=�E��C�>��%�'s!��I)-��E�@4-��ȩHZ!�$]h(d$�� 5 ��Ҥ�$S�!�L5{i��I��b�!��ǂ)�!��DX��'A�`.����W^�!��ȮC��u�.A��j�Y�A�<�!��N�R߂���HD�������4�!�d�|��Q LH�:���	%oK�vh!�$:x���9rg	N�Vq��6m\!�$�m�詈�D4R�$eR%��HH!��L�ze�-�@X�k}���ƚ�dI!�Ҵ�j��QbE;uaH�3h�d2!��3Y�x떈ڝAx����E�5Q��F�t�ߓ����wC�=}-�=	�S%�y��M�W~,��!��Ka�ha�aC��y¡Ŏ��u�����6|�a�A�͂���dX�t�b���l�v�AU`K�+rJ����/D�*��[�g�������V�2d+&.D��ˀ"\1SK<,aA��
Cy�sFI,D���WD�k��&f��~�ı,�����	���M�b�P�L�Fm��P3"OyrA����]�NX&ٻ!"O�,#��P�^�N��FjI�W�F�[u"O*�(2�ťd�M2 �V�\�4}&"O�h��!�>,���Kܞa�-J��'��	1��r��Z't$�X1��P�DB�	��D�[D��i���&s�\B�!+�r����Ζfvx	sV��2�C�	6w�d ����R� [7��C�I�!�}ApΊ*���Y�Y�ZY��>щ�iH�E8�@�2NT���+��s�!�Ą�gX)�b�`��h�
K4y!�$a�H��1`��V��Q��>�!�'Q�K��4w�Be�g��&�!���p��� B��4��D9��0C�a2�O��ٖ�X ^ "E��#G*��+E"O�x�]�{�pg�G�h�"O� 6��|�����_=��7"O2���(R!{�f�`��k��A��"�S���0�� ԝ""}0 ���ȓ ����ʗ)(@�G�_b��=�l�rA�,<Pud˫L�����ҹ�K�?A- H��֦;h�E�ȓC"|�e�׆%�U�Q� >ۢi��L!�A�wʏ��9�%�3�N���i��� �^� ��ɗ�9������\I�Ќ�X�쭪UDP�|	|��l�b���,�!��	���C�@��p���X���,JH��25 ]��j9��T�@�Bg��9��tS�9����ȓ,L.L���.F�������?�OТ=�{�?  4�E���L�v�>x��z5"O�tP��2����TjF�����'�O\Iv�R35P�Y*���-0�IQ"O:��F�tR�H8Շba�9V"Oz�xqN^�w*��S��q���c"O�<`BFE��u�#%�7tI���"O.����F#`��y��B�e�(�'�d,�S�iV+z�P˕�X�"�	���E2~!���#{[�yH�k��sx�a1�jZ[�!��+�tس�c��uOhݑ�HC�Ul!�$D:�Y+󄅽!>�1!�\��!�y�[7ac+V�'�� �!�Ε�^0�V#�5�L�HCJ#-�!�3�������W��p��OQ��!���j@0���)���	tNV�8!��q������Q;al̩S�
�cv!�G�
[|DrҤL�6S�2�I3#P!�$Ω)QHeyaN�jR"���V�!�$@!��[��Ԭ
�����F7v!�d�'��� ,X���aFC�\^!��+L;�ز��4���$��v!�d�p��(qc/D�+�6�A��X�D�!��Q��8II�ꂛ^���eo��|�!�$�#o ��XecT)��.A�1�F{��O.��o����� �ʠ��'�6=Y�&W�>wbA*� �;��8��'ў"~:��~i�a��$�@%	&h�� �B�ɧ9�rI��K�42v�a7�˄#6��F{J~z��[}oX�Z�	�1��h�TI�\�<���|~	*   	"$�%
�U�<	i�;I���c�Z;��PلM}�<�e�&=WP�adDfjeȲ��B�<��Ǐ>ygD���%�aXi#lSd�<&$D	w��PJ��ɘ(�N(y�h�b�<Q��0�rH�FM$�����_y2�)�'}�,��Mה���@F͌P�攅ȓ9@���i��&���ƪƌA�����:6�`����mݤ`vK^�9���PΨZSG��V=���N�5��!��(08��K�Mr��;5�LDj��ȓqq��*qJ�R�P�VY2��ȓ`�d��ӓ�M�	Y��[	�'��py���ZTp�NX%3I~�s�' l�䁄� ���G�H�y�Vԛ�'� �P�W���l���1y���!�'�@y@o�;O	Z�1�)ʼ`��T��'�ę���M�~��̂��Z�d!�a��'u�d�D�lY^�AR$�c�HY�'�, �F�\�R�|I"B?mt0t�
�'�h���)�
P��D��#h <���'��	!׉�ڑ�t�Y�Z���'Z&l
� �h��YJhҴ��'o� ��*f�d��ǭ��P���'A"�c�4FQXjI>L�X1�
�'l��
1�'G+�Z��;O.�Pj
�'H�aZshD�>V���g֋Nc�@ 
�'^lӤ�j�?_*@��"�
�y�͐	��EHA�&C��-y����y�A!B�ZH��,ɏI���ˣA:�y�E�B��K'�͉I]��c�O�y"���Hh甬r$�#6or1��'�Dɖ���wZdX�FV:&�X�'nh��'�S�Pf\<+�f�/r��A�
�'�Lp*���2O@��æPh�x	��� la�m� �N`ؑ�P+\�RԘ�"O��b�
.��3�0�!rq"O�r�l͛YzvY�G�D�E�z0"O<�2W�_	O�L๓�ұl���3"OҴ6^~��R ώ?a�JX�*O��a���#E��dרM(C��d��'J�	Be�X��f�7D/Je��'d�[G��H	CS���Xgh@Q�<i*��C� �y�
+W�lqP� Q�<�JJ�+��)!����X��bh�<��a��P7d��fO��>��S�Nx�<1�ˍ��1[��B�h� ����q�<�%ɜA�䜚�ُ&X<�+��Qf�<U�")n�bb��	r-R-���E\�<1� �5�A3"^t����uj�c�<a"ҰS������$��PA\< C�I<Y~���(��"�FDYb�S��B�I�/�+��L52�`�mY�C�	�mPd�����}�̜��$՗.�C�ɕQΰ��A�f4��c�U���B�I.\��H�͘!2��XBbHR3"O䡂�l�
��a3D[:Q},ٙ�"Oԩ����/mR�Q@E�a �"Or�ae�P�cwR���Љ�P}Ӓ"O�H�K�+:%�H���3S����"O��	1�4���S4/4*,��q�"O�q8Q��;?(�Zc��5F�RH�"OhXat�U�v�����)�HI)1"Oi����,q`�z2�q���!�D66�Ai���/p	R!���;M!�D��|]b��T� D���ad/@4�!�f��ᒢE/��x��+��Q�!���1P���%�7B��;��= �!�D����\����)w�A@`֜U!�$Q�*M����!�-�4�Q��ޞ?C!�D��<GN$�0��.�҄�ݘN%!���@��
��'_�J��Eˉ�F�!�*��"�n��X�CL�<�!�D�����K�"�2-��O�hE!�$��(`���F%�����ϯ*!�D	�e�)1�˔h4X)��!�!�D�Ip�p(%I��EF�X�!�).��3���%Æ�!�S�f�|i�Wkݹ.���P��^�r�!�d]� rV��D�q���a��C�!�D�)	�i�e�4���)捇
Q�!��)u��y�͟�[��'�+L�!��$:,����!
>K��#��[o�!�dǒpJT1WO:>Vu���K��!�R:
�D��ӡ{�����0�!��J&j,�e�fРk��`eڥm!�Ć�F���C@��@��\�#k!�d�*�8���/E4�<𶂐-�!�D�*^? ի�"]7+7�ดD- �!�A�M3��ա��q3�Td�B!�DV�b2�����(|e��	٤E�!�$�u��X�bJ�0 ��a4��3�!�d��9����d.���x��F�:�!�d��F� 
�����*�	,e�!�$�]��T��^����i�:J�!��W�Xq`,;����h2	0.Ҩs�!�d�/�5�r�Q�P7�0p�B�!���6��� ��Z��8Q���:n�!��sZ(s@��(�X��٘v!�� 0���g�l���a/3H6���"O�1i$E�'�*����G�/1	��"O|-[aIfUI"e	Pb`�H�"O��C.���XVC�����*�"OdԱ�f��9�5�Ԣ]�a��p�"O�|j2��N�lQ���H�H��Q"O<��������FI��H.6�if"OƅZ&�O�jD3�gAP����"Oxu2$V�+<|����s�`�Y"O�b��çu�`5ZCˋF��`xG"O��#I,�^4u�A6f� y�G"OLT҄��4/b$T#6�J�w��
�"O�!���]�o�޴�
LX@���'� ����cH��Ё�ۮ��L��'&X����	�T�0*V�j�Y��',����W.D����� P�M�T�Q�'x��c��k�L�s�N�L֨Hb�'Ĵ��.�a���免�@�dc�'̈́\�@D�g��E��,F� =q�'i2�nF�$Ä����	@Iz��	�'��i�d_�q���!�NG�8:���	�'��h!��D{C��5j̹��'�:�R���E��,I�#5�$L�	�'o6ɩ��E�6�@0rmʻ0k4Y��'�A�E�0<]T9"���W�hlk�'�6mH�O�-C�O�Hx�|�'؜��n�� "���3/�b�C�'�i6�	02���-ڡ),U��'����ʞ>oւ)�Ā�'��$��'�̩��(�)w2�|	���2��0�'��s�M_�D�>�ꖦ8$|8�'�]+ Α�*[��[�G��l� �'��l�g!ōF7�scַ�Yj�'�P$�2��q���c�?~P����'S0��)L�c��1zRhǒ `� �'�����,�>�-Pa�Լ	;����'~\�9��8p���	�Ȯ4��'��z�N'6����u�ê/D�TZ�l��SԡS��6h�G�)D����o�xI�t0��`��Y$+)D��+��PP�S�V�&�!C'g&D�\��J��,�{r��!ht>h�$D���D,܎F#�m�q唣T<��A� D���Rf�v-�<qV�S�>7ءkd� D���#a]�o@R|@��V�0&�t
�<D�pJE�<]�&}w�X4<���Kv�9D��e�~����4O�4}�l����8D�������G��KP�[��'C!D����D��KH�X��B���ෂ:D�hCb)��vi8�H���]���&�"D�hr�h�P�a� �^�瞭��
!D��!�R,W:��@�ŉA��K�� D��tn
�!��|(s��5���J"a>D�D �ɗ:l�l�Q��	M�8S'� D�7�W�߲��ˡr8�e��B=D��JmHLV�c��� �Z��9D��ւ��_�r-��F�z~�q�B7D��!��.��L��Ɂ�6#����j5D������$���w�@�$Y��/4D���
G���4�e������`�6D�����w�:�I�a�1o��a��(D����BAR���Sl�=T^��� �'D��A�d�0MbV��#ǅ(3�	�R$D� �a E�_7�:�/D7x��&D�� Th%Ϝ3���CA�,�b�(�"O��*���\��%��(�"O��S ���x$��b�62^���"O�M94��3y�~�S�	B�hb�"O|��`&���\\�q�S"�"O��R�\f�
�@`f�H�FH��"O����̀1G`FM�E@�[�"O��Q�ʓUƤ=R�D4ҩ�f"O���b!Q9$��0tj�E�.px�"O���T %G& I�*f�(�� "O�u�d+��gd���*S,���"OB�8f�S2�РC�j�.)�����"OBx��h�j�Ҵ�=o����"Op�qw�X|t	2�%�$]��j�"O����WJ�`�%Α�}?�9!"O�,�e���[�22m߬��qj "O�i0��o,~�r�3q�8͂�"O�A��9������j��ze"O��8����l�4�yCZ>�V���"O����V�o�l�Do���骔"O����<x"�*g�&zڬ�"O|�`�9�)�
�� �ll2Q"O�L��[6K��&*H��d��6"Ozp	�m�9O �b�ߏ.���R�"O�$�R�]{݈p2nN�`l��"Oz�,p������̓a��	"�"OB���jP�!�|3"L�L��<k"O0z`��Q���K069T"O������[�����.ǻN1d`"O�4CT��g��]2c�W}"���C"O���
�(�@���b�xx8���"O�]�$B	#.�98ŋ�]vPPp"O5��[;JE��
V�y>��("OH��i�LwD�Xe��*
���"O��zr�^6:pT�a+�o� ��"O�I:5��
	Q0�:�jN& �TD��"O]�B	�
u��-lõ`nZ-s�"O�Prb�TTQ�*@E\(!!"O��Mğ1�y���"K9�"O���s�'�����H{=0Dӓ"O8qK�'�Z� ́R�R*�a�"OZ��,œ��<j���&
rb"O�E��]?$ۜ���Z�?x��Q�"Ol�2��ۍH��eᆃ@�0�Z�s�"OLtJ� �yC|��6@�=`&���"O�0`�BST��|�P,HEB��w"O���cm��n9����L\�G�La8s"ON\{�N�6O,azeK��hp
"O� ��C=��VD�v(��Cg"O��E�	�w��Hx
QU?���"O^q�0�� |�Դp�IE�};Ҙ��"Ot� �K��<�<9�7�.,����"O$q��Ɏ*���q�� Z�,T��"O�d���ռC����͐U����"O�-��=�(� U
�T���"O4a���gI2X÷)�?:@��"O�I%�0D`8�@Th��=p\��"O�1����0�:c��n���"OEavڦZ[x���C��i@"O�lȇ�ʹ6CH[��3'�<�k�"O�u�H�	�&��D�iNi��"Or��@���	l����RZg"� �"Od��c�R�!�&`��͉D}t%R�"O�q�'1!�
D���i� ��"O�  �IrE\p�x���ů_���� "Olܡ5-�4�X�Ŕ�E"OXX`𭟖K��	�e�#B�\�XS"ON��T�Ҕ $�g���"O|�{�k<P�IN��p��q�1"O0}��%;D��
�쏔S�l���"Oj���G2�����A ���ه"O"Y�E[*i��1f ��yU���"O��C�
�6D)�iG�Ҵ"O�ĺ%DMB�3t�^3ZDd���"Od��A���ca�$�J�Eɀi@�"O��1��0ƴ�R��A80�����"O�t���˲ �d=�6��&F��13"OP�CE�ۄV�� "W�V�\*6�2"O���l�/nM�D�0`�<����"O 5sq�L���\��d�'Q���6"O��	l\T	LArc[�.��!�"O`,��J ��� bO�>,���"O��GiТSj-	a�	p ^	��"Oҁ�T�A'0^(h�.�3lhn��@"O:Q����XM4䛔:NLՊP"O�$�S+�3!��8�H	8pD��A""O6L�цP�^�=:�,�aF�txu"OZ�s����%`�Kt�^14nI`�"O��#�b�`��i�K@N�"O �Y��)|CN��`F��^?���"O��&Nʬ�§&�3r,.5�"O�qpDJ+��\��ΛR���"O��s����h�c���a����"O
d�'ό+b��Y7$̞^�Ȁ�&"Or		�'�0s�����;$�Jav*ODd��#�_�p���M"1�^�x�'?*�J����LB���;��
�'V*�@#+ޠQaN�3���4�`�s�')�Y1�+��VEp(��dQ(:h9�'��i�QAQ��n��+/`P7"O"CG ټySdD�`�(S$�6"O�ɱ`!�2%�|=zs-�z�S�"O*xK�m�
 �h���5m�x�"O8m�eE vtKDK��R X��"O���� �j�5(��**\2�"O*}sE��.�V\�t ��mL��"O�9ٶ�O�\ޕ�G�޲&81µ"O�ɡ*U?�$ܣd�RX���"OjݻGd��|�2M\�
��4 �"OpuQ6��0L(�=@VlеU�z���"O��
K_�QЊe�'��B�ȬY"O�;#�ׄR$f�S��[f1�"O2툕��7"q�����D:�"O�	Sa�n/�(�E�!��%��"O4�Б��!e�pl�D$˅$;�!�"O���C!E�D�@ ��@�/X�@� �"O:M:���LH^{��U�CR�l�"O~|)�L&r���y��_BC�r$"O.�a"��zs����دB����"OL�B��Vٌ�z�!$T���i�"O�y�T��3( ����O��E�"OʑӠO�QH�����m��}h�"O����� Gƴ����.�N���"Oj��c�*m6@�Pu��wlH�X "Ox����<4�y��	�~��t!"O䔃����Y�yH�#��P��"O�۠L�hf JgdӑZ��u�"O�H:�ұ�� �t(����"O� VU��Y�vQjG�E�T)��"OLA���I�lb�mq�/^(-� BR"O-��a�7k���?:���"O&Q Q�ÏN\�PK�?�H0��"O<s2%�)�Z9���1vF�y��"Oj2�ܞ%TQRQ��s(����"O�m�p�W�FU(�!"��;
��83"O�u�aK�=Ϛ�����7	ne8�"O�p��(\f�U����](j��"O��Ɉ��Fa�3d�1!1Q"O �P��P:���&D��mƴ��"O��j5�я��e�.�8 ��+a"O^��&CM!|��(T��A�"��""Oxm�Pc�H�N�;�`�i���j�"OR��(� m ��	�^I�6"O��%�9�tMɐ%У{�X�3T"O�ku��#H�vi����g�F��w"O��q�h��T�
�)v�1S���1�"O�}qD��Y��@��ԔK��m��"On�R��20j�ʇdw��;�"O84*�O̟)��2�ޗdh<;�"O.�X&NR�1�nM�LL
P�|��"OF��0�B��4)LѰQJLq�f"O�)��� M2i� 	�-G1P,X�"Od%@+�l�C�.C:G��|� "O^t�J��x�� U,G���I�w"O�	��ٖd��a��%��3w����"O�cW�;f^�ł>^��""O|�"��3^Z���N�S��ĳF"O|Ij2�K�>�ac��2l�h5��"Oxm�ԁL�JKt	��ɇ�h��t"O~e��!tG��`�BC�zV�Z"O���+ 44T�&cK�]f��0�"OԌ�qi�(�*��BO�H�jT;C"OlDc�ɍ�1E�#7c\��d�a"O���
?]����&0���'"OZ}���?J��aPl�;��l��"Ott�ހa^�ȓ�*���fD	b"O���"J��0F��QJI.�8y�d"O�U9���D?b����1Q7F�"O�T �`�Q\��v��ε!�"Ovy F��Jǎ���'2��S�"O��(T�A%_<�Aļ~�(��A"O��*�O� `�捝*&(eC�"O�|@g�O	=�m��T�_{z�+a"O�P�k��*���)]*��"OZ����W0>�4�00�Z2ZvI�"Ol�8�&���h�P'�,L����"O($��䊬`\z08����J�1�$"O*�ZW(��q�9ڰ���w�.�K"Oj��K��<(�+��ҔR"O\�x&e?b5���3��%`r"O�<�� N�:|�!�Mnl�Q5"O�J�g��H�)ʧ��e�� "OZ��3�� 4sB�C��$����d"O���q+5j�<I٢ ϲR�0�"O@<)�IK�g ,x�/�:��J�"O�D�(��3�(u�4�"O�+����YI����E��B���"O"śg}̒��E���D؆"O�-[��+t,�AB��p٨"Otq`ӂl-Np��Hז"�����"O�Cg�n.����%�P��"O*�A6�J�=d�f�,9�~;�"O� �T��b-y%ځgN��&h!�"O:A��F�+A�>Ex�*�^}�4j�"O�t#���	WG�\9pꍨ1��$"O�����MXf����B
F�:\8"O�:V
L�6J��̔-����"O9��+B�5K�/��4t�S�"O�y�PFE?�4;!8S,�P"O��ȓ���BM�"S�-�g%ݤx�!�ą?&�$I�A ��wB�xL!��;Ol�=X�gίW���%bHv�!�dE�(�p�� �9��I�1�!�D�1&�|0+��S�M8���M�!��Ƃk��B�&/JBdDA�H�^�!�DT<�J�jSL��AB\b�'�o�!򤈫`��E@t��;������K�E�!�d^�_>a��*_8ׄ��6��(�!�$A�a�xAgȔ-.�,Q6���bN!򄙋S� 9�v��%}�T�"��;5!�$"�jlˁ�M���F�'!�ֿ0g�Eч��
}S�@�2FU<!����*W�ӏ(^�@�f>\�!���\T�=��g�9ZX��$���!�ض�੻�j2��`�Q��!�ɿs}�(��ݾa)6�i��U"*�!��D�#򍩐D�bDe�%��0�!�d��e�SM7s�@zp�V�~p!��ˁP�4�	�~y�3�6 !�_Cz�����
�΅{Q��%�!�DE�Z�|aB0D�?}V�R���!�B�$̈́��F�фf��U�G�!��!` }����3Hj�!A�#Es�!�Y�">\P:�Y4Z`�mY"����!���,��:��U%+O��wÃ��!�$i3�$V@̺^�H��` F?U^!�d�{%�i���Ӑ+�h2�ϐ�i!�D��Sah|�0,W�ZpBd`bl�3O!�d�12��Cڎe@=3��W�vK!�d��V�q��$s���b@�4:!�$���J�;�Q	!4Ԕs4��F!�dܠ|���$j�*�{P�P5!��d� �t	H�E~�9����T!��U`2Q�2�R�gv(�H�Y�!���!9��h!�´��][��\?,�!��4-���J@VHզ����v�!��Veb=��h%z*����J�v�!�Dٛjq�l3�n��8|�	�꙯ !�_W ��PD�z��,"4)4�!�=C�h�#-O�l(r�
��o�!�$E'2+��A�MK@�#�
^�C!�D_2�������v!cEꐿ7�!�$� /�(�`�p�q�e/�&�!��ܞ|�9�΍H�T][�-�B�!��`u�d����@<����f��;	!��.S�x1J�,�3-3�Yr���i�!�$L�/���S�+�o Ш��՝v�!�� �kZ�L�E�!L�!�+ZDx�SE�4~/4����	1�!�]��~Y��ǠC,�����6^~!�ɻ/��dX�kF��0:�+�!�dGL��50"���H)�z`c�"OI���o$ܙ)�����eP�"O�x*��ƇKڂARoίf�P�{�"O���U��6x�����$?�Pl�e"Oԭ���Y�Qy�5H��1Q�X�	4"O� :]!���G��eA�-Ӡ}���"O�i�6�
����l�H�<��"O�Ȩ��_�JQb�D٠]��"O
��T�F2=؃Æ�$�|���"O�C�i�m�z]B�	(t��-�"O��#w)C=A�z��Q��#T\��i�"OjHg
�o�<@r ��V�dx"O��.Y�s�4���N1\��aK!"O��Q�f����Qu�߯�d�` "O��0̕4�:P���gK���"ONY)`̇*: �h��T�%A�E� "O�u�=���4��&ؽ��"Of$K3��)3���%,KR<��h7"Oʉ�d�F<4�v�j��G�J���5"O��p�քV�Fay�*	7kN���"O-Z5떛Ŏ�AG S+N�l�V"O0��t���A��숁�5b���1"O�z,�6~��ih4�K�eH�l�D"O�hֈ�%4�� ��>��`P"O����崝xu���N��qP"Of����w5�l*G�I��B`�F"O��tK�10I
h�t��p7���"O��� �2Vj�
���C3J$)�"O ��C�34� �����`H�"O��ۇ��a���"s��%
�^�""O*y9r���,��')x�|�p�"O����0���K㆖=	�n�`�"O�ݢ��5<�E���
�V��U"Oh��Ŕ�n� E!Ȼ ֦���"O8�3#� 3�F=Q�B�v���#�"O�����3�n��a��{��
%"Oj�H�*1^�¨+�gV<��H&"O��R�[!B�&ɋfI��P�̋q"O�8�dÒ�/�6)����>N 2�"O��J�d�f}�bb6H�(Q`�"O�lY���C�Bu(D U�	�X4"O
�F��M��b4B8�V�"O��C�ꄜQ��qA����0r�"OUِl��k7� R��@�扩5"O��*�m�IP@m�WH��>�Tl&"O�Ps"�T�M�)*��R�.�@9xR"OT%�/�L��c��T)K��q�"O�C� }@��qC��*{.�#"O�m�7�Z���,Cf"O\�w�;��U�3/б^���t"O�i�n�B!�$@#�������"O$��#�Ր}����oш ��u(U"O�ɉ׎�1.Ƽ�Y�ʷ\�.�Z�"OT|����4I�)9��� z��1�"Ot�9W(��WjP@�n�v�H(��"O.X �H�x��!g��3v�Y�"O(�I�FY�?���7ޗ6ת���"Oh;6	�,O�����e�H:b"O��pS�V�v̂,��j�$R�h��"O�rk
[T�&�M�!DH�"O�Z��R��ˆAJ�M	,�p�"O� ����F�r$�	�Q�*d"O�Li�$�2;�F ��.Ԋ:HDa��"O�bS�L(Z\��ь�&	�t[�"O>XZ��
8�n����()����"O~qbX1lk��p��B)u%��"O�yzsE	~(�u���^�xL�B"O�S����uMf� @ �Z]s�"O�Ys$	7y�:U���^
/���*u"O� �yAa�7�����?o��tÁ"O�X�WJ�p/�`���A�4����"O�P���!����J��/!Ԡ9�"Oh�*�/�4_���Do�)Z@"OL�	�.�>&���m��-��q�"O��(Ge�D��`m�[�l��"O�qk�"r�!R�KL����"On���˩-e|��T�� ���"O��Â���M���9Ȗ?w�YB4"O~H��$�<���L�.�)jw"Ovи�`"K�h�̓?�ԐbG"Oh��$�_`x0Z�߫i|\�ڥ"OZ,��V�\1�bbI�'kc��zQ"O�!��m�$B� �bmNQQ�13"O�PRϚ�p*>��L]����"O� Oߗ2�,\�R�ئ^jL�"O�)8�L�$���P�ˏn_�0��"O>5{w�ݱ`��*Rf�*B��
 "O:Q[0��cp���\�A@ղP"O*1� Q$H ���3%��l��"O�D�4�O >P�hY�!� 1����"O�%X�޼8S�4˰�S�oh6�"O������O;n��4HY�Eu�0"O,�rA�g��i[��V�C�y�u"OJ��GΏ w�d+¤�9h���3"Of�4��73�a:�a�@`�˰"O�u{F����l��`��	/���U"O�[>~a������/�!G"O|9�K�Tz�=#�Km)�"ON P��0��)q�Z1֨�"O@qQ��t�\��� ��H $�ZU"O�ua���=,K,@�G 
' P"O��n� s� ��v��ų""O�!��:4)h��G�U	�lH�"O !;�c�2�����`S�kr"O4lAG��9=}���X.lbXY�"O����G�;ݼ���*��,Y|���"O�u�)�W��q�%	�l���"Ot�Sh�+-^����-�P��F"Ol��@�� �9�D� GN X`"O�Y�#�.~$��3�Ȉ>�҄��"ON��U5!ݞ|;1j�4ka�"OԀ�G&����A���&LY1'"OH�Ii I �P�xGfp@$"OrU�A�H&���ۺ&��"O��2dOT;T�*\u�<�T"O��Z�#¦������ИP[�K3"O�%x��0���G>=Z���"OX�s��'z�� �`����"O�Eq���:��Y���68�a"�"O�ٛE���Zd�t*Y���ѩT"Or�u�:U���8ekY>C�HR�"O-�WǳX�yZ�	Ϲ �`]�&"O*�{�`�;|����ν<�B�:G"O~,x�IӋ ���p�!ʠ/���G"O��)��}�a3�ƞ�y�v9@�"O���'I7l�.�#�2EqQ"O���C(Ni`#͉�e�$��"O��Q%�-���@kͱ ���{�"O����<Wf�	�l��'�:M�"O$T��̕�|\��e�xy���A"O�uPc-�9��,�௅�jd�1�*O��q�t�x���+���'�l�yr�^�Un���6G�B\4���� ����ɕ�K1L�P�LL]/���0"O�m�T�٢!�4-9a���V/l S6"O&�CN��m�dY괄Ы]PE�P"On0p�@V5[`��n� "@"O:tQ�B-R=h1H�A[,<��@�"OdA dOq�!�D�l;�"Ozu�'�_F5l�s5a2װ�A1"O�!i$�^j @�*���)`3"O�t�U(�񊜻I[�Np�2"O"����I	`��`�R�"@��"Op-�w��֒��ʖ�i�((��"O�$�S$ #j�����!s�	s"OԜ3�&B�"��l@r����l�"O�u��H����n�?��\#�"O6�86'��q���# C�+�i�"O28�D��6�i��^�S�2�+�"O�p (�),��!4�%���r�"O��@� �~����D�6¢��"OlE�L�d�P�ť͵c��t��"O��xGcգh��@`���`u�W"OX%C�9:�b���Ƚ<C�-�"O@��/։G��	�d^.uAت�"Oj��T�X�6��d�7�C�?4����"OL������4�IX3�42*D�c�"O�yHQ�>ي阴�
0"D0�d"O����̞x�E*@��5��͂�"O��蓥]"9�>=�'ʁ/%��!"O��k�M@&T<^y�e�١-�H���"O�ؑ1*	$��`���=�}�"O��A6�%"�B\@aY�5�-�"O���>V�*�"�/ؔ%�ٰg"O"A��5Gmi$�*5���G"O��y#jغx���Z�NFJx<hC"O����)D���W���(3�"O@c��~�lP��D	JR����"O�!��(T�U<4H`�: ��"Ol��r'Y.���eO�V5�$:�"O�t�F�q�j����Z�b'��!"O�dcQ+�*90�֭��=1��"O��3�H�DϠTQ���8v�ŋ�"O�}K��Y5C0�JĪG��|:V"OT1�!��"+���#��
%Ժ@�"O��+V�0��	I��q�6y"OFU�)�;cO������G �j�"O����3w[�p�u��6R��Y`"O�@3��X~?"���&M�}��yi"Oެ8�A�Af��HP��>]��-0"O��aa(P-wVԱĤ��R�&���"O~X�0쏚!>6�VCܟ]t���"O�p��n[:x�ܜ��`{��"O~l
�X'
�
V!�<zl���"O�$�K\>"��<�uO�Jg�՚�"O�H��#Z�zj-�rh�� o@Q6"O\�tk�]50��R'B kHEH0"O��W�� ]U����e�6b���"O�1�����:A\�A\��P&"O�}��΋8>�@�C �ܰ%힩z"O��j D�L�~��A�0S�x$S%"O.X�#��fA��87���(Q��"O��1u�Ѧer3f_q@��j�"OHђa��~�FXKA���}�xkb"O��:e��{�x����ݓO�tt	�"O�lCT'��[��8 �恙<��3�"O�[V��'h4#$�\�+{>Y�`"O� ����ǪBZ��vΔ�5Xpg"O�4Y�K'hi����'���d"O�q��50�`��л>�~�f"O���2�4(_P%���#@�ҥ��"O�Y�n��v����U
E}�Ad"O�A#)��:aifh��6J�A"OPh(0MW�?��{�F� I�Y)"O����hw�����B&S?�ZB"OBU����Gcp�pB���3V.�`�"O2�4�_�l�ek �R'B�\��"O~] ��_!be:9� @� +#Z��u"Op�[��L�G�:U��߳R"�uC"O�u`���uI�K�Hݾv��a�"Ox�Q#�PH0h�.P0 �� '"O��PhR#^`st�܅g����a"O,���.0�8�gM�-]��҃"O��N�V{fB�ʏ�:G� 3"Od�	 �Ѓ#<-pQ��=!.��� "O0��r�S�T<ԋ�!Ƒm1lq�"O܁ 1!#F�@�O� *�fH�q"O�	�����~ŉ�a��]S@԰�"O� r�@�U����`@�@��X#"OxiZUJ�o���ݏc(xc�"O���gҕi�((Yg����"O�I�����Zӭ� R�)5*O��zA.b	������q0
�'��4�v���GJ���ʯ"i�!I	�'L�h�d�FHf|��l.���'��L��ƌw���������'��x;Č�%�qP���.W�$���'�w�.tb�x�!���JA�8��'�ڽZ%IL{��Dpq�s6����' �ݪ�g^�h^~(��8�E �'�d�*�i���@��Ն%n��o�<a����� ��t%��!�m�N�n�<q�d�$ ��"f F�t���"b%�i�<��oZ"|�nm��פJE>h2E�Uo�<�D�	7��Q4kk�
��k�<��Y=4g�)�!^�Vݙg�Cg�<1%�@�?�1T�ד_ܦ9�wʔX�<��(���ʱ�'y��\bP��i�<I'��mO�=
���������Ye�<y���p����'S�|�bd�<��h��+��`p��o 24ɂ �`�<QRʁ�`|n@H7�Ř]��@��
�^�<Q��۽1��31�ѫu��}cªX�<�C�@7!�2M�v
�/ux� EW�<Q����/l�9�D�D,i�x�Jr`�Q�<Qf�u��j�k�9*���Q�<�S�3s30ܲ�m� L1�m��d�d�<i"���wP4Z���/�
r��W�<�c�$T�����O �7��!�KS�<�2-�(*�P����Ā���T�<Q���V\ ��(&�9��Qz�<q���1N�с�KY�{�l�˲G�s�<�Ve�4�k��֛c9�bO@q�<�'�,�H�H���{��a�j�<P"��`T��N�[�06*�g�<���َDh�j��ԑNA���fm�<Y�h�6�8	�l�,�<zEGj�<q�i���jɒ��O� �[ �
j�<�2Œ�c|}A$G�L�V4���Mq�<�3�ĿnS�D�`)ևAr������w�<��[��rY�`E��(�$x�<� nE���/ت(vN13��!c"O�i:s*��c�T%Q�.���D	@"O�$���f���awSe�����"O���'%��Er�-���F=@��5��"O�LئL^+�P����;u�4�b�"Oj��!�I��n��DǓ�|�z���"O:����ʛ?��Y��&�8Wx�<q�ޣ,���T��P�`�h�m�<Q� L3?�����-#�H�TD�<	��P}�,KbA�0 `�$�UB�<�QK�<�\��#w�<����T�<!��޷<3�4��\k��	ʡ�E�<q�j��2�<��٘KɊ���\f�<��$�1^b���v!�j��rJh�<��
7˚����Wq��Z��O�<����S-v��gMF>kSD�:#/G�<Y�AC�"�0�[�,PtV$�pSA�<!��]m�=�&��/pH��~�<���h� ��M�3��8tVz�<��Mƿ4�BwlH�!V�T����n�<����)���#�u�Ę!#��B�<)�,T�A�~��"��������z�<��F�#4�3%��+-Li+ ��r�<��oU�6��+@j̵>���BLBI�<��ޟ3^
	Kf+մ#�B�Z�[�<��׍q��D��cT�GeH=��V�<�#��2�l���H" ��;4��Q�<)�ϻPWx�)1g�k8���Rd�<1��ͪd�ЪAA��U�� �K�<7��+k%tj���0�ؔ���E�<1�b](m��EB��"�f4f��J�<q�`�H/�U�1i��Y�4�����D�<�EC���CIK�m��@�~�<�7?*��#B*ۨ�B�c�nV}�<c��W� ���&S��(�'�@�<Q�U�6đ0��#q�l���&�|�<��D�F�+`l��o!�$C&H�m�<Q �*6��R�H"`�tH p�ZU�<Y�PiW4y�	��M�, vo�O�<�5M�*L*�dY���,m� xvg�<��ZG�l��������ȱ�X�<�e�	<넑�s���bT��%�
R�<�P�J��:��GR>��1��AS�<���-��H��Y���b@ O�<���l���Ct�L]B"�����O�<�A��1f�4�7�I�~��9ʰ�^I�<yA��'%�V��.%cP��w�@L�<i�CN(p=�(�l)�D1 %YK�<�W��'yx�J@d�����k�m�< bZ1	G���ޢS��S-�f�<�&\��z�B�ǋ�(H4����c�<�6`���[�$�:hI"1��d�<�t�-t�6��e�\
E:�Q�֣�[�<A��9 t��R�@��RͱZO�!�!IOPjÛ-��u���.x!��":`��Y�y��ӣD�<!�Ѱ(����QJ/w�۴"ܸc!��#s:����ΈB9���"�:�!�D�K<�����}�E��nV�To!�$ۤ#5�A
��/}�,Q+&�J4e2!��,)UPu�a���srRD����y�!�� ք!�1�5(�x���Lr�!�ΫUi0D��삤4������|!�d�8�֌�aЛ;�j%X%R�o�!�� LXCb��DJLeiD��x=hMc�"O@�sD�]�f	y����P�5 E"Oh�3F%2����� ��S6X���"O�p٧�ʆY@$aTo�F��X�"O��i�G��^!��mA�t��:�"O�k���=��l;ux�{�"O0���L�/��ǫ5[7��*�"Ox���Ǆ"$Y
}@kł��m��"O�5��Ӷn+n���'(����R"O`�B�״T ��W⟐9���"O�H����;B�&(�����6� 1{#"O�9���+C(�(EJ��h|~�p�"O�9pD΍M<P`���х:�(ܲ�"O���$�U:6�İb��J�R$;5"O����ƧeO �*c+M5C�h���"O�@�"@��-�5�9��(��"ORms� 6��#ׇG}�ġ�0"OȔС�\�k\,�b��֓ �Rm�"O`�J�F�-d�p%��ԆČ�Ct"O�9@Fȗ6㞠��돺w�bL�7"O C�/K-Ů�x6 �[�ր��"OԱ:�	�tB@���[i�H�!"O �����x��!��H�0P�'"O�p"�� j$e*��ؕQ���zG"O~A�]�3!���&�āEd��;�"Om��jQ�|_���M��]K�-Z�"ON���GN�\ �GM΄8Z�)�D"Op��O�w芝�4�ERQ�	2�"O.�@��܌V�(IgL��1�T���"OB�a�`�i 0)��������"O�ܱT� 's���
�67���"O,��$5+P�{S(�P�8Lkr"O<)iB���d�4q��IҿQ���~�<���J�(��00�'�^��$#���x�<�T�9��L9.ݏ?�*a�l�<y��O4@���K�&I$�at��k�<i@ʒQ�Z�z�M�>X�8c�Q�<�@Q KN����ֆ!89x��J�<fF�/~̜��娑�MWrܻw�M�<I��T���A>{��3���`�<!�oR�0�0��BIͼo��Q3�K]G�<q�@Ηt����e��HɊN�<��OƘe���/��U[6��$a�H�<���4-xE��������rT	�L�<��ڂS\ Щf&�-8�T�:v�I�<��_�j�T(� �"2Ĝ�2�C�<q��:a��l	V�T�8l+�l�x�<�)�&,���rs���\ك�q�<!e0��ka͕=+1�u�a�r�<��'�oQ�x�r��e�80°��S�<�����D�e"�� �� 
 a�R�<�R挲`�|m��˼�maK��Q�<y���6-}��Qc���e=��gEQ�<ɐ���#�)K�/��8!�0JGec�<�LۼVEՃ�B-d�P��d�t�<I�Q?v�Hx  �&d���R�]h�<�� H�?C�4#�
>�����+�K�<q�!֪+N&P(*��&�ˆa�<���/�b�����YB�<)㘔k�^���IVna��d�<iUk�\��t(��U'B���K�<)f���ؘ�)�9Z��UJR�<����:�<u���8rM��{�`�M�<��ӑ-榭Z�BE� ਼�EF�<� ���A�9v���ħqgN��#"O�,��B�1�P���ob����"On(���*��4	U+�&�F�)�"O�;�l����!cڶw<��r�"O�$@��\�n�耒b���9N�`"O|䘑�\�Z�y�-B+\|��"Opp��N�(�2����͇�b���"OV��e@:Z��[Ձ��V�� ��"OL쨇��#,�4��2�ɶF�f4�c"O:$9"%�s��
7��0���"Ox�s��8w��ӄ�,s�pYb"O�ȃ/	B��-b��
`��! @"Oh�rs�U[�Bh�q�4�xK�"O
YBwLH9"��Ea��$l�9�"O�����S���8r�G�o4�Y"O�M�QN%4�88 �W�F�8�"O�裳G�D�{� [Έ`�"On)��Հ����RT�:d`�"O�tCS�
:p�"Ș$Iָ�"���"O0�(�;���8 ��W�d	8�"O�`�v띆/Z���tJ�x��"OP�:6��0BEF@��
R�5,���"O\�H a�Z�,\5�̢<jH�s"O�����Μa:�� cH����p"O�l���]�oV�{��ҥ�z��"Oi�	�~sM���ו��3�"O�%�4hY�Y)f%���3����"O��ᔀ�+e>p�BHI��ls�"O�bwdCr��b�_�2T�0YU"O�q�F�_7U���r�
 >���"O.Yj�(��b�P�	�G9R��"O m�a�Ӿ?�U�S#0(4�5"O�� �$Z3�h�xW��Q�0"O\�ibE���yH��
&�4Ea"O�@�S�1}&0yz�d
^H��"O��i�V?i�|#f�7@��F"O����K�>bB��c�ɡ�dj�"O���<�d��bl���Pg"O��I�H.�b�4�J�5Rđ�"OI��/X�:"��p#HT5P6-z�"O� b��,�TU�楊�en��A"O�-�cK\�P�z=��e�4��1"O^����i_�Y��M1s��(�"O�w��;5(d���S#�b	 �"O��`
�XC�\�FJʻk��)�"O"�㑀ک	�����?d���"O>�+b��t\r=� �
kH5��"O����ń?@���We4y�"On<k�,er `Ѯ%.&��"OH�Za�&i���am&9VM�"Ob�kWj�<��ଞ?e�
�{!"O�-PQC(\�q
��S�7�B@	"O��TW/Acl���k�L�@s"O|4��������TE�/#�(T"O����&W��+�$��U�-�'"O�,�2fJ�|9���kb�"O��B�
EDq1�;ui��x�"OHU	6K�q�pPA�U2��'"O ���� ʐܠ��\�"a�l��"Oƥ��G�
��C�^�XI�u"O���˺J�<0@v!A�y��ŋB"O�Mqf��*R�vP�� 89��i���hu�)�'N=r��S-����CM�k���4Ӑ��q/��6�Ȃ�(K7p�Ԇ�S�? b�yc/U@�iZ�*� �"O�%J�DL�xBPs�\ O1"O���ϊ�t����U�?Y���"O���ώ�X2�#O�&�p�"OZ���G�z\�j��T�f��qT"O�Ĩ��IH�1��hw�ț�"O^�3#�(��ȃ IP�>f��w�'RqOJC��\�S���x1甈�[�"O����G�B�
�d#�
,����	\�O� �C��|��ay k���t
�'�~����S�@9lq�-DI����Oj0Gz��I��I�̀"'|�V�(��1O��=%>i��C*ch\c�]!,�pza�>��ɩ�p>���K�;6ܨ�
�i��v)�m�i�1O��g�I@`�h�3��(J_�L���>4;tB�	:FcDTj����e.���V�_��$��Iy���6�X�|�z\B�a�~��C� 1�8$EӀ	<0չ�X�M�C�I|����I�����h
-T"��'1O*�~��k��A�va*Q'�A�j�C�!�X�<q��N�x$�Š��Tv��C��V}b�)�S����1�Ha��`�lJ�?�A�f�'�l�u��]��^j�֜�D�C|r"?yF�8ڧ|��M�pn�S�)pC�-Dtbh<y�UI:�ڡZ������AT?��!<�S�O� <;sI�J)(qGK�4�yy�'ߊ����L.b�� �]7��I�'# ��dO�(�`ب�OA>�L��'<����K�e� !ڷ��
�pl��'7 cglձuep� j������'K�mka)7���y��|ς=��'�"})� ��7�t�J�吰<�H�'�.D`B��$Q(�`#w��؀ �'�%ѓXHBx!�
�3���!�'�+�y�Ï:x��˳���)@T����H/��>1�O�Ic�`9e.PP�c�	���H6"O\ģ"��6<b�`�a��&���"O8����~ hY�5���}��D ��I^�OI�� ��C	W���ֽs0r��'-x,��]��"uRUԪg�}1�'J�L�$"Ї~������&
�8a�'!��@�ͤQڸd��+e(�H����IX?��犋e�l�Z�S�?��!l� �0?!�O^С�G��zV��4kU����	�"O&iȰ�I��rT�! ʦz�}�4"OLd��*�V4rC��%�T�@"O� )�(��-$d<��ž>����"O���$�2"=��*1��N�,��e"O
@r�hրuv���,"���Y�"O�5�B)3	�t	a�&kz����'�DS(6��)��WC��4(�Fv�!�$8�6� ǩ���ܫ���:p!��: ����*J���$'P�Fax��I��K�D��l}�bk�=^������ Ei�#=^|Qeh�Py�->D�P�qmYÊx!tk'e�*�8`*>D���T䛊�س퍢T�R���8�O���� �z�Ζ�pI�h���R[x7M2����G�uF���	
R����)7lO��,�	Z�A�x!��+eȥ�Vg6D�P�3�1c���U)O�xm�}��6D�0;��÷q��!����r�J��6D��z�K\?;c8�أ�Ȁi�5�'�8D�T)F���)ΩJ@Il���B2D�� @���%�,2ʔ|xc'�i��jѷi���$��t8!ą�92�b���A�<Te!�SePҥZP+�'sb)r��;�!���J�)���JL7\s� ~!�d :+��hЃ���3��{o�.a1O����̓T���1�� ��ҕ�N#M��O��D�O�t�N��;�.�gb�Ppu�'���T}�J,u>���Eh�����Nש�M	�'SF�ǀ������p�R(*�x$�ۓø'��\I��ߚ �hH�X�w��Y�{�:O6b������	��<��"�e������"O���#+�%v�ȴ��$I�P��|"�"O�Y���1�����ɂ�.|�l9V鉧�0|
+L��厛1��$�Ry�<I��_�Yԅ ��2���DS��ў"~�	�qh,�����ꝱ� � V�C��*/��jp�عM��5��ɞM�j��y��)擲X�*�{�iM�Yǚ��Ɂ6�RC�	xV�E�֢+�>=W$"C�=z4�)r �q�>q�t��W��B��WZm�+�~�t)ԆW�g�lC�I�o��݃`�_!'d!�4@��,C䉚{頹�����;��I!�S0Ly$C�ɋ��=(�=9d�KG	�]8�*}z����,�1¦��w+N�E蜄.k�}2m�<��ٜ)�t�8B�ʛ7� V)T�B��$gl��@��V�0; �Z3
������$�M��WϮ� �fE.7q���KS�<�%H�Kڀ�H%A����1Ke��g�',�\Ҷ�S�e�����H�25��EhgX7bM.C�Q����E�+�����Շs����?����I�-�@ǌo2�H�q�f]!�d��!"�١�+_(VI
���GL!�`b����бB)��!����[AX����'6����Bc۪vh�E���pt��A�'lO��� }2��Tb�! Q�$|I@\���yb�+9��}!g��l�D��U��>�y2��5W+�y ���\3�K��ʰ�O��=�OxI��H��TP�(�<O�\`	�'[���GT�{�I%gON���S�O�=E���*��m�
T.�rA�#o��IpX�`kC�V2�6uh�ɐ�;����<�����2�Ρ#���)�Ҝ��E�;H!�	���C$KC��0Y�C�C���Ȋ���m�R��U�K#,��I�@�J�d��C�ɩPfDr���j�8u��$E�,t�� �S�O3��ꂡ����iA3?��t "O$�g��A�=+��P����7�����I]?)��ˏ2�1P'�Y�@vt�KKx���'�Ip器k����q'�Y�Fm��O�YZ�'��$4�>�;B�P3���Ta$�pFBߪB�ņ�3�ld ,��|��H�)����ΰ?�cV��%i#P\ Y��e�<�b琯�*�u)�GƆ�4�X�<q-�M(�) @����!����N~��i>i&�<ꔇC�)�*�86m�#�Z�k�`%D���3nҮ^ĔY�2P����@?��hO���R��\7��qɁ��*�CO6�:[M��S��a|6���g�-V��	K��H�|p�7J�YCZ��W �[���"O*��u��D����DB]�~Y�"Oh���k�!'���sb��m
\*��'~�$:LkX�r&�Q�U���@�
&!�$/�98F"H!;��i��Η!�� ��aW�45FxĠ'�� ��"O*�����u.��V�OXϖe��"O! f������^�2��aH!"O��gm��Xގ!+Sg�.Zˀ�"Oމ�����PL� ��ÊfߚD��"O"��5m��0�tX"N!x�h�"O�X�0�Ϣk�,�9��9)D�H�"O�� ���+H�����DI#�$��"O8�f؆<i0bV�t
~8�"O����s�xub�*ۼ>X�2�"O ��c�}(�p ȿ?���"Oط 	�6g&����V<�s"OJY�Fý^���jA��	�:�"Oxh��-͛Psع�䧝<�`�"O��I"�z<���w��f5J�ѓ"O���B4	��|�P���9;�"O΀be#�#�5��kF#o�u9�"O��5���@t�uKL8� ���"O�أ�A��j�.�����>i_na�3"Ov��V�A�[L���4;��0�"O����A��m�d������rL��"O|tA��;a ±�h���<ye"Ol1�@��<��A��	?��TH�"Ǒ�r ܎�E�P��2�p,��"OJUk�.��-z�TKo�/*�����"O����4�<�����O9�=9� 9D�ث��N�E뀼а�VGt��#�2D��2�5�N9� `�6j��ȡA<D�<�aF�k(���t�k��e��7D���tǝ�T�"�Hvťn(�u�f�0D��x�6#�D�X��P����Ir�8D�����y�0qcD5:%��7LO��I�nۊ�h $�IA9@���L��Knт�gV1qi !y"O��{V���[#�T{���:*Z����"O�Y��d��Iz�9��Y�E�kA"O|)#��ÐJ{850F�\�,44�H�"O��3�ьaH|��oÙ���C�"O�t�2�ʖ/:����흽/�<p �"O��уf�7�H�p,ʏmk�p�"OB����6+vH9t*T"4Y�1��"O�B!�x�@��Ϛ� ��p�D"O<��B�F(�آ��<A���!�0I,,{���*^*�S��y���gLۑ'�0��U�����y��E�>1zV�3c��Q���M۱�U'G�l�{V �:hv}����!{��)d �o�-��xA
ד
����K�7Z��lYR"��£�T��-�U�HK�h\0�2�L�GA�4]�<L�re���~<���%D��(�7o/r1kvhZ+Tj�
*O�Y�@㋭h��A9��S���A3�It����@�?�~���\�d����)��V]!��M� ���� ��,�&��{���)����@�!��
� @Q|`��-D���WC����eM^U ���<�J���'Ƶ!���C��
,q4��ȓ1��q勜�����݄U�8���'��y��!
�S�z�s&�
I�꙱	�'�N����S���V�H2�ܠ���� ��)�j/��!��1:��M!c�%�2�E(�^B��|�>@�����T��P���ɰ@t
�P����H��S�O��B6-Q���ԋbW'K�<`��'��y*'�� �ر�BJ;��,O�K�"ʈ+J��dL2O���[L>M&�ۆ�.�
2�'�&�J���yEd,ȣ�H�o��LI�C^
7�� �IG�>�!�[�� �14��aᓌ%<vў����ÜfXP��`�g�? H�Qq 	3}�F�ڢW�B�A"O� �a	�~D�����C0(|����'��������*��W�"~�㑧J���E��.9��Ӄυ�yR$��]���b��	GEN������'$&%Y�΁�w9F��Ĉ'/&�R 9)��i!`�X��}���\��P"QBu�`�2O�b+<@����%��X�qO����˚9�l��g��,}u�����G(4`�N-X���|�1eX���Q�ڽY�v�B�~�<��� E�vQ���d�RA�W�K�<Y���YZ]kV5}���Ƶ�^DK�"�G5�1�bi�1!�dX�j[��B֠=#� �)�$�8xB0�-Ӟ��<��ϭ|pr��	w!�͡Ǡ���~�>�FIݬi��q@N7�H��Y���B��ՑS��S��A�`N`F~�d�*��x��bI5���z��A�Of�<1�昬�������[?9��E]��O>E��I�%�ح�T$4i=�������ybB� ��sAٞU/|,KA����2?�P�`����p<y�G�_і93$=vİ�"�Z��H1bAL�j2�(!�/�G�zTZ�+X�]�RD�p����֩�6�<@�(�6块-)��ؑ��93�����	��}L��&�,��q0*ָ|!�Ė�Ѐ�iɂ5"��B��E-o�DHE�4dC�Q/��)�{М���-hP�K� �<���� �af��~����RS&	�'�:<c%�X� ��D�㉑B-(0���
~�
Pi�+m2���Δ5��<:���.=5P��_�]x�c����"�����'^��"�c�X\���"n-j���K�\�z��a+��O����.�(w�� �MS>m7.dB
�'=�A�`�9�0�{U	>�|a��'ʹ��!ު{�ɧh���:7"_�|�~XK��/*����@"O��x���eĩCU�MG��}A�x�ꖛ��Շ�I&*�Ȋ�K�<�t�C�\�R݄B� Lʔ�T��o�|�5/Z�E%R��W�Yb�S��y(4i
E�8��)��@Z(^!B䉘Z������R�1ߤ"���(cu��$�09�>�A0}3���!@�T��es�\�ȓu����,D�_4�d�,zbs!��<�D`�u �3H��aFq���L>p�,�X���I�r��E(%LOT0� ��k�N�
ĢX-al`� V� ��6��!�P1
T`F�@b��DJ�y� ��p���S2ʝ�B�1O����\.C�����g�/�E8�K�~�"�ܡ %���=e0}�4�0v��C�	:;Ҿl���' �p�5��2�f��c-˄V�]"�`��\;�É6��A?�c��.<����@�p ���R�j�<Y㌒D�B�ɶk��Q��A9b�M$G1�8Q����i�H���%��XZ4�	L�rPxS`W�;�Z�P�B�D����&���ӷ~0tr�h��S�ޝ� Έ��
,�¥d������h�<-��h*,�t��zBQ�p�W��n�(1��j�m $�ɗ{@���τ�U~�Q鄎��+1��+�!�dԥ9��Y��텺=(�Q�U)FU�S��N��#"�m�FPo���7�6��Ͽ��	��gbT��e�< �
��RESE�<����<>��WI50l2��2�� ;lI�S`Þ|��Y#��ӊ+�$�' ���Tn���ē%�:f��iȞ�q"�S3u�<y2"VS2 ��],�l��DQ�cf�|�Q���j2N�C®��N�@�5f͖��v�F(sB��i�HX�|��!� ��!@���k�\���O�)�JZ�.���cǈ*�����=�Ra6單�J4���>�xt���ǒ��2�$�O�x��W=����b��]L������8�xœQ��>.Ÿ)��OX岇#�{V�eCH���
��w
�,~��0�T���0�?A�#)>�����h��`�˜OcRsm�*k$f1S�!�3P�(���4��҆◱&fӧ����vGT�d��8�G�8&�He�t�<1vcD�䔘�mSM����IVfn �`�ц3�RA���B/8��	E�t�Ҫ	�ay��ڸvOx�sb�Ի?yR4@�[\ƾ�[�G8&gH�룧Wg�5�M|��We�-��Z9t����4�W3tFr@##�D6L9�u���(�O>�rD&5�Y��

h`�8�S8)�x�SAؒ  ���І����d�cN�b"�4�� ��ഉ��n�3�+՘�@Dʥ�	O���#a�W��D��a��%^���Ndpv�ݢ���JG�_�o*:Y��ŀUe5�)�'{�ص��nO�@��B�KX�ip�wx�2����XΚ}�0��?j�RPq���J?�Vd*R��`���Z�V'r!�-��clW_�,���ʂ%Xx�`��.9�p��Un�>L�:h�e�~bӋ\$|�N}جO��4��lt���� D+>��r��'��q�cS.D3:qX��N�s�N$��鑜w�-�c҄R���x�KD�;��I���C=$�O�i/�Z������	P4�dL-8y�xi��ɏ{~0��0`D�hE���3gJD[P�ׇ�I�� �"��[+���i�8L��e�
�3+�q�TE��,O��[ŏ�Hobx:a��.o����OHZCӋ-`A#m�8Y�9�����26:c?��s뒅(V�zb�� 0�����?�"yز �$2.����4If I1b!��Z�K�S�F�(e����!\U�P��;w�(=1ޟ����C�L�Ή��	� �yb�]r� �����1Gy%N��?��LT���KwO��g8�(�#%��J�Py��� �q�`�9��L�9T����T$?��3�?O�<��	O�^u�O�̜H��2�h��N�e�f����ĪQ�ĈYƣ��lx,5Cu�Noa@�Z�k��WܥCD+�vU�s-B�Ike���d{���8�~�qě~�=ID��\�\	W@7_�Ґ2�oybE\ �p�s3*L �	���>T��x58�
9!��8C@�7	��ٰ��սn�v�Crk�1Q X�`*:�O�)֏@��J<�5��*�f��g`�ة��'�jP����}���/���R�Uo�(�`��'8����XR�p�m+&��\�O�� ��<	zH3N�;"�^5"���Rj��3� ǵ!�&�{�T w{d5�&I��yB����O] !���g=�5�o۝�J�x˓	�~�sT�78 ���6O`5�e�#}�=�WL�
d	�I�ӮփYT$9��cX+@���gܓ0���S�So����=|��1�<�	<x��J���'Ge��7�B�$�ҕ��{��9$���j�>�xro=�O~\�fņ���B�hyÇ��oZxD�Q�>���ُ
ѤԘ����$�T�*.O��k#���rΕ0X�,/jC�	�kgʐ���Pf��K���i"1�&F\��`6� :1��U�'nz�S�b-��O�h0�T�� ���'�X�ד&�E��G�3�:�	�h�LȰ�O��a�"�G�2�e2��&݉�
��=�E2�+2�p��'i*d�=) �ۑ1��m2�i�1��Y�m�6@E8b`͹-Þ� ��5O�lSS�1�@��M�)gr6�I�G�+����4!�����ZG#}�)�K��kU�>M� `EA�ПͻZ9P�d�7B�&uH�/F�
�6�ȓ4��e
B���TY���A  u���mںOB4P�
J�T1 ���;h���H�-�Zm����)��L�3��*�X���ɩ_�{��E0;���'㤴㵊�+CHs@ϋ��q(A�ʺ\�J�B�@6��p1����	8L��)�="<�"�' :V�F��d@�U�H��D ��P��8 �m	�� 	iW/�$n�:EgԚ�)	�(�(SSH�>7��9�����!�&�G|�`��dh�ʷƐ9A8��*fD�~�"1����Ŝ���� ���b�'�P�J&l�OI��	g$W�s�ܺ7 �&�(K>�g���>���=����)�&�F��*����� �\R��h&��D��'b�#��@c���"
������r:V�'G J3��>ٳ�P�P���bd����D�����D
�61\�8��'�R�A��њ>\d-C���%���X��@�����Vr�'ʘ�[�Ґ����^fX�p,S�Z}������s5S�%��MZJ�m���ĝ�#V�M:GF']|<�>���� ��acp�#ڧbV1Y��ܸ/ٌpR�`ߢCk&,�<Y���#An.$"��I�:Q�`̣U��$4qN��40Qs:�s��G�Y��'��"}�'�؜����0n~���"H�/Ȋ��M9ʸ'D� D�,OH�{Rk_�oɞP���̐{9.�p��iM`�2��ov��0aH�C�C
}�	s�FB�M�����9b&�`�2)�?ɵ��@R�A�`Ϙ)�|��'#]k�DA�0Qv� ӓ;\΅�.ſ$5N�QK5����>�e�)6��h7*(�i��7��d7�EW��C�(�K#�ȓ׭=�C�I�Bn�d!��Ϯ||�i��QbL�&0��� B3�˘Fzr�O`�]�7���� ���I!�#��g�t�XdT��(lO@a
�*�\, �(gȊ96\�J��'�͑E�v����OT!��˅ �����C,R��FղZ�(q�J�zZ���T&Q5XC�I=u�4��'ƌ%2��e�dQ��Z�2���V��F4\DC5�]�N��)K���O*fݰ���'/	����i[2�Q��3�y�W�W��@���(�,�x`j'�M%d	&�l���B�O���H��?Am�CD� U���"`~�EPv�'�]g�T$J�~� �	`��� IVp�F,�^��@��O \�"��3d#��rӓO6�����$|�'��D��H�x���F�Zs�S��*`(j�$�r�;}�="��ܺ	�M�&�)D�LQ�kަ?�r���d��>���0 F�<�1N�vE�����Y���	&���A�d+τ<��I0r�Q�g`�I�q���0?��kņY|.�9�L�E^�D��B�r�vBAm���,D��6+�$ܦO?��.x��Aچ�P�T�P; �_MQ��7ꚤl�>�A��ǖ"���҇@�s�M`�����χ=>�;`�'e|-8�!S����T$R�����KuX��w�חhax)8�GP�5��2���>�`�N�2�y"䘝WUTT�"
��k��ۍ�hO$)F�Օ�H��-[��88h�Ba�2XhzI�`"OR�M �F�q!r�^� [t=s@"Oz���;+���Pj��)���h�"O,���Ւ:��j�o�u���x'"O �x1��+1X�1xM�|��X��"Oe�eL�$���s�n�/g�$ʠ"O�%�7l���p�Ϊ7F�
"O�P�g	��l@�⛂L0�m[�"OJ1�,̗����gӍ3'���"Oڵ:b'ч ��y���,EȂT"O��s�@Ļ-�>�Z�f�}^ 帶"O��j���.
d���&�]j�	1"O�8�1�9��s��8f` a�"O���2�w���#��vCjl2�"O�@pu$�(\��z7�S9w3Jy��"On�2�i�;*8U�e��k� @�"O�ຒ�@?�2��2��cݞd4"OZt��66��$[��7���as"Ox�Y���Y�쭸&�ؼ^<�r�"Oļ��O�w�F��4��;:�9�"O>]���o�X$1�	��"O,!{UI��mZZՉ���;3��qC"Op�wʋ<֢�
����\l��2"O�swe�)�Q�$΢62x��"ORU����,���cI�_:25Q�"O(�d��on�qh��?6����"O��X���@��y	V)a� y�"O�ň١�֔�V���an�"O��ω[��#@شzTh���"OrS�!Y�]�Ԍ�� ^V�X�"O��Qᬜ�
A���Ո�"V0Y�"O�Py��Y4�d��4�N����"O�<�0mZ'r���TE]�t�*=0"OH�D�ݞ#�$\1����8�"O:�d�d������*�
�(�"O��"ɀ�~�TTSe�;M��!�v"O�Q2�GN�$V��C�M�p|pA"O�2gC��]��y��eZ<|��mK"O�I1j�<��)��d����,1�"OD�$�ˉ7����RaY�Jb
�"O�$"� �^5D�qƀ�o�t	�"OX�3��$�J]�v,�)y[����"O���d�
f�	ґ�۱,�b���"On� v�W���h��]&
ƚ�5"O�0j��V�A�U�d�=#����"Ohy(eg��G�@�q)Ԟ ��0��"O.�!�aD?c��q4ǒ:Y�@�"Or�r{䢘bch�<UCl U"O��Y��M�rΠ!�]��s"O��d/�=b������ ��(	2���O�6�3���k�J��!v�ǌ/��E�U
���
����زt&��=�|�K�G��j���ΓKe���m��v{vҧ������B�IV�,x6�@Φ���<D�� \�1��DDt�����
�Nc\�����7]x&�
�	p��焭���U#�z�V�P�#�OR�`��j{Z�AR��S��p�.�b=rg��'�\B�	�O��#I<�E�A@�����=�VS/z��x��/_���Oo�E;�Ȁ�=���)Dǀ�\~D��'�@Q�a
�6.5jqbc���N���s��D��#�$0�T��,O?�@Z"��� �W�Z�Ԥ��j�VC�I9q��ԋ  R�m�j#5O�/B,˓I8�U˱�?W��Ó��R��C*�T@���$<XZ@��I$>^JhʁȀ+u��)���T�S���"k���7�X^<��z�^��r�2ZNp�"�P�'B~q@0f�0����r�I@�3Yʡ���IQ05yƩI�6L!�d�?}"�A@Q���(U�	%�V�E8�ޡ��)�1>�s��~~4ܨe�<�^u��~D�MIdK��]���ʩH�(,�O����k��R�J��N6p�
qi4���ЙƤ�&e�!�$��K/^Dy@��4u�l`��"Ӏ�!�D�*V�X}��g̡���J�"Coؑ��j檋�?b�>���aW�'��$f�,4���"O^�c�I�)`i������`��OL	k�W<=�O�>[i����16, Bڙ	'0D��xf�ț)��� B����'0?���3�=Jo0O��ʧF�5� (k��Lz�e*��'�:�SG�<1��-P�	�*5bҤ �Yn]x|�!+ZB(<��$Țk��Pq\<V�~)���PJ�'�	���O%D��}�ҤLMe�����:��z��D�<�R
N�h�!S����	3���<�֠��6J�y�;}��)]k�>	��)ݞt�ڌ�QG�X!�׭q V�!�lI�jπq��R��IzҊ1���ʼ��xb��z�n���	�[
,#W���0?9��������/�7B��q��e��I3҈Z5�C�ɀ�h���ć,}`Ij ��l�#>�#�Ś�а�/�Sm�����o�Ljp%D�%uB�I��J�k�ȍyU�5{���p��	]Dd؃"�s�)�'QR�2������UUd�+�d�ȓAF̙ ����H�P�sq�F��&���Ǣ�+�ybl��V��V�ß@��}'$��y��vV���tsn,�)���y
�!΂�PO�b����R# ��yr�>w٨x�qI�� �;Q㒕�yE��pT��5��Y� ���y���h�B�"D�2]�8��
���d|�p���+-������42&Y�f��9��<xs�	�
a}⦈�.>@ ��9d��\B&Ɉ8��H2PaI�ڌk���e���9��V�ڴ�����[l~x�2�*ʓ,Ѧ��"�"ܺ��d
��'<�p<��  ��Ԁ������ȓ`ʀ<Z����
�(��׃8H�
��H�Q<��j�K`n%��𧈟�S�v�F��_,2�ZFn	��y��FC,ds��V�O�r}j��ȫ?�t���T�t��4�W�P������hO��R�^���@��������':l���_&�$�%��Ag�T3e���d2��u��^��0T�'��y�B�|~��!T(�0�~�S��G�&��Ict�
zr��h�O|�C�@��9�F��X����d%�7�X[	�'��L�g����<"1Q)1���)̕}����P��!��"�p�87�,8p*p�|�
A&-8�oȍi��k��M6d'B�6Xft�3��Ն|�40:���4j�`�ef�?!�Xi�'�A�FMp�ƫ?I���?j	&�P�va�)2�x��"\GD&����,�O�D����&8�7�Lw�$���Y6e��ŀЊ@�xF¼yߴA?����^���Va�[!�L�&�jǖvBў���՘�R�"s�@������] L���B����i-�6U�"��� z/!񤚶"J]BE��&��CVLL�ў@��퉑F�D�
e�	�(���2ƭ���mKj�g�!��O50�)b���g�2d�Fg�M��`]#s��y &��v��Ӄ��TK@՘+�~��F�[|rB�)� �A�ʜ7,�c�G?`E�d0%Q�P@S��l�����'��␩�C�e����t�f�
�t�l�2g���O<e��-.s^x��#�;c��t���3$�ʓ$�I�y��C��pq��C'�C{��+�I���Ov�QFLN�g��h0 �T���'��x�+T�az#'�E�F
�PC�'���kXy�S�O"X��#�������ۙc.L���'x鑶$M� d0!�e�M�RD����'���"�H��m��e��OE�g��US�{�P\hv��>i�nd<J�lۻQ���C
 s�<��퍈R�!�7��9��'�n�eA���_7�ȟRA��Ȝ,$�r�BH�k���	�'���3#ӊd*h��o��Au_�068�@N�(���<���!{�a�t��2ul�
׉C`�<)a�N�c$*@7�R{<�e���4�x���p�&M���>:b։���,�|9�h�(e����D�f*���ReQ�g��%�'J�ܢ� ��A�J���aM1�@8�'<qZ@h::#v����X`��S�OD�(#�����P�g�F�L	?�"'W*y����D��h�`#>C�I�`XKdn��RЮ�Z7A�;dw] ��7G�2��
(wZ�{�0��֜y<Z�G2r5fa���@�O��R�V�s:ՠs��3n�B�K ֜~�}2v��>�X�.ż&a|"�^�1����Y*O�H�ե����	��8�I�?��'�Qv�Febw���-�b@̻W
Q�v-V�t��`%�*k�Q��Y���RU��MI�PA@�V$R��xlZ�_�@@����,������6�͓
���}�7��v�dh�5l�wD\@�P��Y��K�ݐ�8 {d6O�Z��۪RBD� B�(���$^�$:���#�J������gܓ8��%��ݢw�h��[�<=�-�=��mV�؂�1�l!�S�:�(�@�&��
e�@7Y^rXzrH��w�tB1�'@������j�X�S&nB-Px�ءd�	`�ܻN��[�H#0҄�'�Ъw��I������<b�\�:���.K�6�S���F�<iIQ�l���;�&*=�Zԓv��f�	���
8lk�O���˓i���k���j̧J�y�cnD�̊��Ƴ"����뉑8�6�1쉸|���_�M�� ŋ`�������~�剔-u�ъ7#�)x@����I�7���J��$J�~�q�fP�I�㞰[S�E��Ҥq���HD&�Ԁ	6���z\���L�&
zLKAG��y����g��T<p�] M\�@C��L�B`$ħO���l��X��|�w.�
榁����y��U��QP�A��TP9��e��y�ʌLJ�=�-|���	�
�!�M��)ɲB�s2��2�TU�%r�69�(�eA1�6��d���GJ���&�&U.�m�A,<|O�`B��^���d��M� ������{Vd��(���L�?�8� ��>bO�e�Q^>�<��m�I�r�ѳ��s��MbѪ{x�DJ�J�:,؈l0rd�)��irn�BB�a�1"�!Af��a$�a}Ҭ�"��5�7�({�ዲ%�"��O�yBe�U�D���Q��3yV���Od�A�r��%m�(R���x�Z;��$ҫa��$�����e|EB���5\�Y�r)�$.8�'^�E��ɞ'+?$G��I�&K���s�|ui�.�	�lI�$��䓒h��$G]4��f`�f�)ԤZ�7 jԀ5�P��	4ceX�?�'�TJ���Q��'��)!ш���M�R��24M���ф6lOn|���+7s2\j7kR��9�p��2�"��ä��Ob]z��!�����@����t�$'���Q�l�J؄�$&���!iMm��ɑjH:q7Α�P<(("���%�b��X@(�)K�=�p퓬	s載ԯ  �P6�_�1M�b��@vF-3I��F�Č� EN�C �Ӏyp⭐�: �<=*$�_���u�>�rC�8؅ �$n}z�s@nO��}��Q���\�(���$sf�y���:���G'N�7-�9�,A5�����=���Q�r�bQ�+^�.���b5��N؞�˲��_�v����'4���`O�"���N߿PBR�N�@z���~�az�l�&d���I%G��,®P ��î��'Lu���ܳN���&?e���\3O��J-L'y<��IA�ok��q��ah<�e�� ��XЏ̟1�F����
 ]\�" ��H�.�z��D��ʼ���D�T��� A3 ��k%BEy2�P΄p��	)u�\Q��$��Ě0`��u���U�+G1qpIK���JQ�,2B��$R�=P�b�2!`�+����p藺q&�D���r�<� L=RG�Y�lT,ٲ��2!0@�Z�X���5Ɛ�(�nD)P��K�g�U�$�~
�M!T�f����2���2�Ax��BG�G���,$x7Z��X�*W�%����r��Y���%Ȃ]�O��}�	�����t~|�B@H����=	T��%b|��QG=��Pe6)�B/`���i\�lG�ɘ�l1kgHQ�O�az��+ybz%d@�U�F-aP���?�gfW�EK�kU-4}J|
�d�4w��
�?�(��M���-�2Ǔ�]}hB䉥�xyQRDT1h�ZT �o�*�PʓQǪ�R!a>C�*T{�i%XT� 	M�\�OK H�f)��X���捀@����i�ZmpR��4�l��%�/ےu�!�ʜ����7I�IZ�I�ҭ�G���O@Y+T��j�Z5����	$�D{�ɵC���6�5[h���b�5 Դ|�qe]�c�	����%ێ*�az� ��<bR�h�n�3'����6�>����o���'ƤU�$�*ਗ਼[)�Lc��֛Y�!�
Z��B�h@<l��!L٤i�ў0����5��>-���ʩ��w���"0IY&�:D��8�lL�%�$1�Z���6�;D��"c��i-(iJ߸sS��J*D�9����V�r����8=���%D�� 0�N*`�IcWA�����&D�b��$,6�I�DZ�2\�͊��(D��3G�g<�ӱ���q����5�3D�ZCm^�qF��c$D E�"����.D�AѧS�%�����D�R ��"�)D��TjO�
�ڌ2˅M��= d+D���3��L�q��.��a��$D�(�� U)�^���^�L���o%D�h���(4��R���i�{rA D�xrOec(�kI,E(j�DRT�<��ƯU��A��k�j�tB��J�<9@B�}�Xȫ�D�.0B���,�D�<�7��&���[U��*��Qp��C�<�3�Y�#&�:��+a(6}�4�r�<�6BZ(�0c�c����ª�s�<���J�(��g�hi̼��G�s�<�#C
���,�EhV���`ץ\E�<�O���;��_>�l�taSX�<�E�{���Bf(�n|�Xw��U�<sD�
�N�[��؁��IM�<駆B�.6���HS4����(�I��0+TI�Ff��d/��2\'.�&4���e@ˣk.�wb��p��lJ�(�O��S�O�L���C
~$����+���5�P�p�2L>�%QP�r�>7-1���P��R�R��M�Ef�6�1O�I�UF�v�ŞiB���"�^�!ZTE��e +]$��'B���+�)�'E�`��u"�%&�T����t���[&@XjRn�{��������ڂq�z��RNK�P�4��;O�)��'��Q�l��4=۴I
VfY�U*��������XeHT��S>%R��Hf��k��")�٫䢱�D&�ܣ,O����Z�9�̔R�i
>|���R#Rd�axr�Ɋ��eÖ�^�3��`�D�!�B�	U�f�#�Ŋ�j�~a���òl���d����
 dk�JM�6���K�[y���'khи���&M�S$ɜ`�\�K�QZ<�7�	y��ȟȍ��� Abzh`��0hM�d���I�0|�GH:),Py�*2��a2�Yo?i��>A��>����g�NQ��$�f�]Y4����@n����d��?q�ȟ��#u���s��8@��	8e��,��Jy� '�u�S�g~�O��-ӷ�X�a��4�$ :;͆Q��'6N���GӕZQ������/8���K�'v��Au��f$�@�(�#��d8�'~̻&�tE:MȀ���^MȚ'��I&��S�O�"�+�+!�VP�n��P��#�h�'Aa��!��.�Iԇ��	��@6�N��'�d#=��:�t����$l$,xNO��Pc���'9ܓO�Tk����9��'�P���� ��y��Il0�}*w�A�%�tIX��O�d�'J�횠J�O=�O�;�q��Сc���e*�t0�}rE"9D��Zs痃mQ�q�Re� TQ�eg5D�(x�� �=M�a7�?�$QC$/D�(;��^�eȾ�Z &�#�De`�.+D���ugF�[�H�jRf�v_�k��'D��b ��O���hQ�Ài���j'D�����+�r�s큷ZX`"�"D��y���B TSUa�zӴ�	vI D�����0�-�^H�F�r.=D��(�ȟc�ޕ1����Kn@e���6D��@�I�\��K�ᘢ9(M�6D�d��@5*n�)����o@�͡P�)D�0�l�
/7�|(���-UL�u*(D�<idA�z�4ٱS�O2~�DX0��$D��0Sg�$�Q� E
�\��.-D��@r�V�z�J�IAJH�>�v(KB�)D��x3��5�\)���(v ���<D��%5w.@P�j,vy��Ӧ:D����W'BMv�p	іs�� �-D�Ԁ� 
�oF�M����7V=��h�+D�0��A�	a��� ��K$%s����<D�t���ȩ&N)a��dy>����-D����Ǜ�-�z���+Xx}3'�/D����ߣ(b�=�CɊ$�Lax��"D����B�^����"��Q�95B�)7�=c�$�X��sHC��
dLй���"�N�f�ʯC�8]�4�`'�F����,���B�5���ǆF�]�H"i��B��n���G"ڨ3�U�����B�I
%Tv���'"Q����` .B�jIčЦ���-[�
!�B�I�tu�i�wB�+d=:�PpT�}<$C�I>������;�M L�(\B�I!MӤ���l��baJ��0B�	��q$�B�R��(��a�&nC�ɭ|:�����M6���5i*"bC�	*F��Q�c�F`�x -ܩR�B�I���@�ʀ.�X���*_6;B�I`i�5cEb�%,D�"C蜈|s�C�I0z����z8�ɣ�NU��C䉌`��� C�*a��9�����C�ɼy�!15���bЮ��q+�C�I�H�=�$�]0��׫��1FC�	��&8��"*��A�"?bP�B�	�}�M`�V|�d��"=�B�ɐA�R���̓�L�^P��E8 ��B�I33�r���(d��s�g߇��B�	�ywr��[4P $h*qnڀ@��B�ɂ,(t	�6�C�	o�i��� S&<C�	�C�l Ca���q�j�5f2C�Z�5(D�I"N��t�g'����B䉲]�� L[�*.4����C�	 ��1FW���!���c�~C�ɩF�~��2�җ �(�:�-ٛ�%"O� Q����H�Ѵ�G�x���"Oz��������J.t���rR"OZ�`!&O0@�����'�;uN��r"Oڽ�2#�-~&b٠��_�gd��`"OTM�2@P��Eآ0Q�T�f"O��R�F�&g��`b�g[�l�t��"O��p�J�z-
}�'͸Q��l�"O���F7f�1���fҍ��"O�  �'�I�:�� �FC�T-$"Ox)WGC�}AFʦ��-ɂ��"O��N�J
�����);�T41�"O��#A�U'?/:p�c�ڼ>��tx"O��-�
p�8g�ۻ � u��"Obq1�$� ��I!��@�w"O���II�c?�QJ�JݛR���Q"O08[E�Żh����#��X�P"O���#��4�艃0��,~��"O�4sa�B�!��wAӯuyh��a"O��cٛ ,R�	���?�A�4"O�)���R._�Z�����j&j�8�"O|x ���31.���-��0�c"OT��Z�-��};U��2�"O��P᧌�~�`�� D^	\�<Ex�"Od|i���%�6�BS�m��Yy�"O���'��0ez�Ȑ��P���6"O���a��4��M�_�R��w"OR��횮AN���fQ�0����""O���͌%��E{BL��e��!��"OZQ�w �*3��`�`ќ�4�P�"OĹ�D�c[���5���z�P�"O�3�B (~��zu.(�L��"O���ß���f��2���#�"Ov!���Ιw6�S�)4ϐ��"O���'�T֎͓���;r��]sP"O�a��D\% a��c�/y4�[�"O���+2����w���B�R�"O�8/y6z�p�d�7gL��YG(�Y�<��*�~��mh���L�$��aVH�<9�R�)J �I6�����˶,�B�<q0/�'��b�@ AL�b+�{�<I�$��~��YCц��W��-[�d�t�<��,��b��m�p�1kH�BIH�<a�ػOtE �J�'�PJE�m�<�@�V�Z.��m,N�BHk�<I�ɜ�8����2�� �Y��Bn�<��7-@��偎����� �Rk�<��j��s��Y�`eF�}��m��c�<�̇�P��r�ƛh��u��	x�<	4/�����@�R鞽 �b	u�<)�
�}.Xs֌�
^��`�&��W�<�oܷ ٦̪�DOn@��fgAW�<���wF(i���1)�P5V�<��J��m���i�������O�<Y3�ƫN��E��<34�Ӂ I�<���˿%�b��>KE��S���\�<1g�ߥz-�� ��8pB*�C��L�<��/����Z�"̪DҴA�F�<�F#�{��HA�!�.��e�w�<1��P@x�Q�8_��dƙx�<q�Þ5+�t9���ŷh�9��*�s�<�w�:6�aZ���=�|�P��s�<�Cή6q���DZ:<�(��M[�<�N8y��c��T M8N@2k�Z�<9#C��9���@��;�n�3���\�<��3ö�"��H�y
�X�_\�<i�� ׌�[�䊷YO���� A�<�'� _�����[���\���z�<Y\#hiH4�͕�kf����|�<AS*�;ž%�c�V�w�L�3� �w�<AW(E�7��٪p�E_n� `�w�<�g��mK��F!<����w�<�WŊ�g��`�#��[UZ�9��}�<� ��b7*N�H�	�le�i�"O��qM��7�M��fɐQ�qIA"O�,�����O�nz!��($M��y0"OȕP�B�H)�a����B�q!"O` ��O._ElYS����^x`"O��@p Ǒ6@<U��#�/�ܝ�!"O6�Aւ�BVa�TS���"O��DNU���ѳЀT�_�
ݢ"O�ub5��M[�,@S�(q2��"O,(���R4?1�\���!Ζ�K�"O�˖�^<O�4���nK�Q�q�v"O���pN�	��9�G�M1�E҆"OF�����43xE{҅H�2��᳅"O�X
U��<A�����c�&:��<�v"O�)ab̀F�R�h�@�;w���"O(}xt�2�P�`��[�KuT)�@"O�� �-cf*Ԡ⁜� V���B"ObВ��T���`B��EQ&E�F"O�H�"�~߂�Y�`�)O���w"O�I�2Ì�, �y���1�P9�"O��g˖�n���o_=Ǆ�k�"OLX*�4y=��($NޘK�tTXT"O�`i�! ؄}�_�&z�:1"Ofx#F:7�l�"�
B<R T$ە"O�@R���۰�{�
ۿ	�Er6"Ob�!��)3C	a#��x���"O�h�diƨD���bV�$d��2D"O�MQ�L�Sd�1��@"P:�0�"Op9�����},T�4m	�(\��С"O�(tiՍOhi
�!�
���B�"O�D���������]5�} "O`��'�5��\Q�C
d�0y{�"O4�)�P�qɶ��� ��/t~��"O.���ҝJ`��o_�_����"O�� rE� ~�i!�\0D�p �"OL����V9>�Ve�%*+6�jf"O
�0�!],T�1ȋS�,��"O�e�@ΊQ��q���ξ]��q�"O�i�W���?X�uC�HT'5����"O¤�ČƔ[|dM�VgP,��\X�"O�`�� V�8��/�	�J�JQE�^�<��EU,h/�"p��p�C
��M�"C�ɬhC����V�?�ĕ�G�&�>B䉒H�M(s�X�I��zw,��c:*B䉏W	�!"Ea�"�֘���!2TC�	�;N9(�$� y9�Ԓ䋌��B�I�����(f6Xlj�@�)z�B�	$R��T`͔(j@X`�K8J��B�	�����P�I�$HJ�2�KDr��B�2m�1p�e� P�tI��0"l:C�ɿ0�Ư' ����Fp9�H3D��!��Z65`(0Qn��9�R�,D��p�FX	[��A8"���� 2�7D����:$KJ�βxQ����r�!�Dݡu4؇LG�1�����*s�!���]+��3�+6$*�!�$��aT[$�[:m���۔�b�5�ȓs��Q��`N���	Yφ�ȓ%�
)�4�߾Xo�)��� ꒅ���R�;k� �@�o"���-D��Hbf�V�8�@�f�	p�.�e%+D�<3�훙t[̅)lԻ"J$�æ�$D�<薋ʁ
"4MӰM�e�8y�/D��rk�:8��Ua]���ɛK8D�� ���Q��=1��B�'^�Gb��C"O��+��I?OH%	GW�S�<�U"Oh`Yc�����f댦�,��"O&|(�B	��9Q�P׆=
�"O=鲡�15���s�Z �"O���   �