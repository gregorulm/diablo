MPQ    �-0    h�  h                                                                                 }�T=f�%�z���P4��B���}�t�շv�H� V�L"C ��FUcU�3��°�.�t�ϼ���I� $\*�A����t+���Tx�FП��3o�֤e�r��nj>� ����5�Y����,���F�a��8�Z*p��l������|7��ˍ����zŧV�Yiˢ��6�d��:.�v(q�=��S@�L��d�>F�Ɂ�8�(�x��&56�"7�Qd�ȳY�����q���4�ɷ�4�0Ծ�ILnO}2��[$5UǇJ}����:�|���yg���;B%�<|	��+��+xe�9��BP����rm�����jMO���+�C07t�̡7���T2�K�5�Ǆ��;k���@�������7=*�َ[�	��	mp����wX�lϐؼT�ٽ��w�B(��R�E�*��VZ@	���� �W�L��-���@��R\�7�Z��=J.�+S��Vs��"}���7ز�g|�с������>J]W���2�V��FΩ�[�@�Q��a��TVWΤӮ�;����]f0,;��g�y�
kI��e��XDL�9�D�
�����%��j�;��>�U���qICd���#m�b����#t��N�vzeu���2�uBm���wƃ�/:V:�Ƥc�t �H`pYm�'��p��N���'�J5���㐙�R%P}O{ΐ&�r���������~%�f�����@�V�v�(��%O]�n����9|��/�7+����ET�$����_s��Ɲ��y����+���G��U яh��^d\[5ӯ�űCq	�^�q��
*��q@Z�E�1��'�0��%�A����T���Ђ�2��2����C7j�9���L��z�uf�P����E�-���@�\Z<����6%���U�^�G���v��2���a]$���[鷧)O�X
�,S^D��KǗQϕ�e�m�b@i^�br4g���DM��ky�%�Kz����\��oa��Yfؔ{됩NB��
�¾9� |�Qމ�1 q�y����0�4o	�͎�[E��o��:T�Qv�Ry%κ�C,�){Y��B�������`�M[E�9��11v��S�I�&�����[�+��Qg���I����X��G�w����$�~v=>O�NZ�����#�So�O����q��ǐC3����z	��
+	����������`��K?]
!��Ǵ�V�0�Jq��}����<;4��N5�/*�&J�0�U(�[�+�*8��'��e.q�6���6�S���$��֋�i�#���\�K_�fO��v��}:�q���XT^U����F>o�΀�)�o�~�\�%o��t���G�e���xa,�t��7�"Z�J�����Fm'�	�j\#%����7]9慨�р?�d�8[��k��.��-��ӥ���GێZ�+s�ֻ����{k�G�d���3=��*PeZL,a��|�䙭* ��?�qƴ���"B�rmq� 4\��Z<j�ms+<
�n�nNC�%�;r`}@�
'Er5�� [�]�È{"�*����w�(qu�$�F;��%�qJ�7i=�c��CO^���Ip�g͟���b������ܡ����ΜU�q�@/JG F�ML5��Sc��T|�sy ��|�A$kH�;I�	<A}��c�|e6�!��6{%!�깿��w֊�Y_���1��h��[W੶���-��?�"a8|^�g��d,+�Bc���Š]�ؠH�ؑBC��y!�8>ť?;"
�QWDʏd��O�w��O��n1d���� �@'^?/�+�5R���ç�����6�D���Q�N;�}��ͧ�ċv�w'?4	�P���5�m�'�����[�����o���'r=Q	q��y�ʀcԢ�e�V�_ fأҬ��d|g��<���G>��u�[���τ}��)��f�l�a뿀����zY���O-�Gނ��K8���t)���t�&�٦�=�-��;=�Wl�a�ަh�Хt��h��*E��$Mӟ:`$�c\�*��?�����T��T+���Z��R��ˁ�v+��#�-޹�EL�8�'�/���xx(��q/˰'���EYDmĊ�������%�1�8`y�4�ȯ��ፁ���y4��}g�n`%*C��YoW�����i���7�$�9���l�����H!�e��2�pZZ `��.WE�"c���o����6���C��{k��YtX{Q�� s耲Fަ�ĥ�1g�
�S�	�i�[ �h� x�sg��!�=�Bߠ��2���nG�u��;;�s����M�h��Q�	4S�J1Q+,)��K[~��R(�L�)	�=H�)��_�GA)J��8�;Pp¥?AC��/��g�r�
���Fԟ��#��<�gKct���� �CF��1k+�u�	6��8$#��$�����ݎ��Zs�P��7.�f����(C�oƮu�?���s��"`�O~9ik`�S�R�f�8#�����fC��H���%i~��"���#5M�X�m�_9�v�Q��gWM�W���m���� �蘿�M�P��
�g3������%����Ù߇�v,�]g�pRl��`�"p\� t��|2����E�HbPT��[�/���� �����\��� '���f%շ��#?�;����Ϊ �}�>������v5aE�Ho� Duk����믉K��v<V~3��:�}Di�>���j�:���L�4ȹ���ş(�L��ru:�C�'j�e��W:�U�'s�����<��Q ��Yd9���n�i��a�Lȃ�KV)a�q��AZ��;�V�\�cy��X��?��h(wv�����M^=���B:�~�t-ch�Kb $�P������^�!�Z�Ic��eA&Ǥ9�x[�c�.'��)k�.�Y���o�U.Q�r���`ٷTO̻Э��q%�X�ǈm���V��u�e#�ȍ[�8���"��7�Y}";Z1W;�Ci�3_=�-���Z[�	���፭G���){�G�Ǟ8ܚ�'*����b����7�E���.�������n3��z��JE�n�ä`#1<�:�WK��;��:&Ú���/�g@�5�Z+�d����*���d])�����Xw��ʤ�/[u��)N�r�rxmmg�^5|oA��%x��|(�������t)�P-r�$ǡٽ�?�$2�3��l%Ml�����|���$�5Rp��=��O�٢>��/��j���7�7_kE��PX�8DT�o��i���7,�����n]�J].�y�{e�}d@���D�o��[�s7�����['tx z����mej��Pr���w��0B��,�E�y��qR��Z�`f��U">��Qɖ��٧��6�~l�7�7�����HH]ݹ��B�|R����F�=�-e[˖����a�����[rsޢQL�I*)�k-��>�H��&��)�����)2:a#��f�pb~|_wS��m�59����*<f�f�P�ru3N��k��͠,�҃��I�K��)`�!
�C�d��� G���2W��79�[�̞�-H�Q�7�ϕE�J�[��ze���>�d��ٳC����AHU�]YӴ1�5#/���HP���a��5��ґ���w!f^/��eU���ށZ ����m�"��ϋ��[ڷ�?�3ř}{�k�t��J}���!��pF�H���:��Ӵ�����{���d���O�)�g�@���|&���w�8OUE�ሽ|y�_�TH���'��
�9nĻ���[�U�wWh�sd���j���^�(��������;Zث�,�'W������TvAA�]�`��XP����r7��J�S����nu�q-��Yeˀ�J-T�!@�7+<S��������9�٬����vu�2+<�aX������b:^�s2�,ΉZ��梗�����"m|�%��Yb-�l����M� �kT�o�������]aI�ƕZa0�6Y�P{Ɓ�N}�b
DV�9�'�׬İ��q8��.�D�V�oB ]�)ԊE��ʿ�:�\v'�%IVC�{�A��?��$����[ �S9��X1�Q�S�;�&�C�d��ȓ�c�kg~I�:ܕ�bXny�G �j��[J�)п�O�,N8�����k�S�=r���3�l}|�"N3BR"/		m?+书�P�R�����Ї"4o?�!� �%a0��|��}#Qj�7���aB��c&e������+Ȏ�����`���\:��j馔S�(� �����������W�l_�ϕ�&����H�}�2L<����SU�LW��;{oc\��ͽ���n��i)�OI���#ehx\��t������3L�P,
�!bɮD��j����"�7�#�c�ћ,d������i��-=�ť��G6�ך�3���Ӿ�xW~�"����k=Q?WP`2L����7۪��폑� ȳL�A��NNB8Kq�����2��!�<�[��I�i�G�ֵ�};�Ce�6r�r��H]X�L{�6f�QpgB&�(l��$���eqe�i���:^X�6�! IkZ��mS�����} �9Y��~w-bL�vSbU����FDJ#��h��5@|wS����A�:c� ����f�kC`I
O�A��vc�t�6�����^!ט�T_{w��!Yz�����hgR3W���Wa-������"�B^���0�*+��c��i�;� ؛^�3U�Cu!�>�@o�;���k��* ��J͗C��O[EC1�%�L5�@l/Kэ�X���I�!	��=6s6!��'M����;#���D?���0Ȭ�k���W�kx���H}��1/C��8���R�o:W�'-��	�I��0�%8�!e����Z[ pr��g�(9�'RA۸B�y��uUP���&�yB��p�'�(����rq�{���z�ԩJ�;G9sE�4.�`nt�}�OU���=J��6�AWǫ���-�����/�c��{^��LhMn��`
3\(q����ީ�)<�G�����햕]uRe3�֨@o�谊��yZL\�~�)M�"R�BK���/&M#���a�`x�m?������<S�%�f"8[AD4ߏã������y�b�Xd�nS��*�%IYj�R�N�9�Ҧ���,?$����8+�8Yw��+�e���Z�8��IEW�Oc�	؛�������65{&�Y�#mQ�Ks�~CF`�_��1[��eg��ĭ�i���\Dx��gV��ż=��K��'A2_0;nb_�wT�;�=s �)��V���<<�d��SȲ�1l�)���K6}J�,o���K	������
_�]�AD��Գ�iPKl�?|�q��y;��r��
���F����H\oK�d��!�P�>1:�3|w+rL	Q%W)v#������(�x�>�U)���7�N+����+�(�z�̷u�;��׏��3�
*������g4�AK#$�b�B���k�
K�$�c�=dٞ�3�yΚU�,a�	�kW�Cl�/��݋�k�� ��g�߷BMw_#���gxTx�l�W� �L�J��t6���^9]���p���l����GL�2�^�./wӾ�֦��b�4�����/����S��{D\S���Ӽ�X<%pQ�O�?ޯ�֧���Ō}F�
����G��5���Hj�D�8���[S�/{H��:��Q?S~n2�:[��i�'P�����D�gBQ4C�N����cE�p�hu5����jH�x�r��U��Gs�Tȫ�LU�0 �H���i�i4Aiaf�˃왽Vd�E�AU ߖ��}iy��;MA��bw���y�VMYBh�<9�B�i~'��-�rK=z�����8��YXc����c;f[AA�Q9[�[�h,.b����V)t���5oA�$Q)�1�:�<`�g�Og����O%�����:D�6V��6Q #�#�[9�r��J���o̴�`;�_V����p3:C�h��C	���<	xGs��)����B D8�K�'eˍ�������'������/_.�L<ݕ����3�_	��	��iDe�������r�$�u'�����u�N:��茋g�Ն��䑔Rn��[����]�!�����wIެ�_�v�ʵ���Mb�Wmg���P�|ʓ���ɗ}��5���|���2r�l��{�?����;�هe�lj���/��83�5�Eĭ8]�O����W�JF�m�'N�rxME�2vX��T�B:�ҧg��M��_�j�����J��My�!�q<�8.���VD�����_�f�藅�E�'ϡ1z��:�'��e�G�+ѱ�@P&j0=�, �h���`y��q�@�5`f��5"ٲ�Q���皯��Q݉�.�
���t�,��V��]����K�RE�<���=e~P[���%c��sA��D'1�s�^Q6�:I���k�>������)����f���=a.����tNp=4_����543}�tE�*��f��q�3)0�k���;���I��U�Kس*){�
!���C�*3�SҲn��M���eWF�V9˟����Hp�7@��಩�h�S'���>�5�|���C�%w�܌ոX1\���#�y��bG�ln�n��pPͪ��n��#w|h%/��p� �Y* ���ֶ�m1=!�=��:�d�r���
�q�F?�ȁ�}�fc�@���fD�I��	�\f�	�ƶH�������O��"���y�|�����|��s#�E�=%�wH_)j�<q��d��B��D��:6U6>wh�4d��%�/�y���T�ˣ��&�Z�	��'I�'�Cߛ���шoT�5�8M���K���">7 -|�����>�u\'����˻��-�-@�2�<a���ObP��W�T�룞�vZ�2ƮaS���XFηkљ�zx,I�\�����ۧ�S -mwd�mb���,�M��k/DJ��#��G��F)�<I���UaK�Y\{8{���N���
�	�9�N��˗����qS���G��6o}W����E���%�X:�Lv.�%ĉ�C�m
{σ��x�\�{���4�[���9�b1l.S�Mj&���������?�g9�lI dx��YXI6�G;[�=�E�|7�4���*�NS�)��7C��3S��Iiv�g��}+#3��m=ϫ	�`+�����m*�(Bo��<�}<X?�%�!��X��?0���}����2�ŗK���G�&�_��KXh�_�+ٍ"u�[�캦G!c���P��ڧd��ΒYO��RC�_DY�uہ���6����'�8��h=UG.t��P4oj8�����
�*��)r�ec�xW�^tcz/���Nn�ˑ/��v��_�j�r���7.9�J�Ѷ9<dxy��˞ϤH]-����}�G�ٴ��%��˾��R}��\��VV=��{P[s�L���F����'��F\�'�^� B�C�q���R9��	�����< �˸$�@���;q=}6��s�r��ˮ6�A]�\\{آq��W���d(g��$i��T%q��Ri3��ZQ�^��T[�If�L��_o����������P��@]h_����U�S���}�J�E"�� b5�9�S�|��:��r� {�x��Ȋk���I%�pAs��c��m6)(��lPp!�f_����wL��Y��'M:hB{WV�µ�<�-�-��5��"ן�^ؽ8��5+�boc�����ؖ��Ԏ82C0S^!�d��X9;��ǟv�ŻA�E=^����O�1�����i�@��h/L�f�k���+�|B����65&����2;^�����氺���-�K�ު��_��
��#�%�l���&5U����o��'��	�ڜo����<JC�e$X1�U���,��"ϡ��ҽ��ۓ���^�u��h��Z��'��++��C<��bm�u���n�z�T��E��G��.��O9���ttP�*V�O��=�^Y�1��W"�+�T�}��/������'��_M	��`�>\��˵���k��M�б�����R �����7� �ףm���Lב1���Z�]���+���/�	��Bվ{�tm�����R��w �%*��8V)�4:w��Ggˁ���y*�;�3�/n���*y�Ye�����������A�$���� :�s_�~V�e���+;Zбu��#E��ic�|2��l��R���h���{�LY�gQ�=�s��dFT9���k1o����x���i*��^��x[�)g��K�WwH=����V�B2�tn} �8L;�]s[�7Ճ-�������S�ǘ1�c;).�K��"'�ڂ.�	���ߧ;_y��A_X��.m$P&6�?���8&��F����@
l�/F
�%���|�K�t����8�9<%����+-�%	l�g�9�#�����t��P�Y�#7{���*\���(��~��4u!�\���6�L�����L����I"���#_@؅��Y�� n�e6%���X3\����5�Ց���塀�W5Z���X������ �{����M��� ��gӕ��'Y��;�ۥ��4�O�X�차]Fz8p��lDn�ۘ?@�M�ѱ�Hә����>�bM92��k^/l���֡�-UV\��ض���X�F%w����?b����������}���Vӂ^c5��HHe69D+&W�Z� �J+ɉA�(�,b�~���:���i����<�����ݡ4����������s�Nwu0i��:�j����&jU	�s�͝� ��G ���d�$��iO��a�U�ǽ�V����SAPt��񩣗�ASy�'5�,����w�����/MTg_���B}�Z~B�-Y��K�,����P�9�THA�vac�@uA\�9���[j��.�C=�_��$/]�@��o� _QD̸�]�`�7�OB2��%&%�D�>�'���V��u�\#k�J[t�ؽ�k����>;��q��9�
3i���%� L���؝����G.�q)�b����8�n'���>Ww������Z����.�������d�3*Wl�*�p�d�b�����񍓚��^'��ް
������	�g���h�&�������-���]_�G���|w�%���/�i#�x�u�(߳�jm��'��c�|%��Ӗɲ������イ���=�r���Y?]?����	٢ųl��)�sa.5�;��3FOcx����d�eg��\����㭱�E$��X� �T<6RÍ~�߃șxY�E4�����J��Cy�`��$���r�'�.D���3U������O�'*�BzVYu�B�e`��P��{�����08d�,[�y��qH��0of
;*"t�hQ��e�B:��Eܧ��-0���X�g!���]�ox�� R �׎'��=��[�v��Q���=VF�&��&�s���QQ��I ��k�/�>85(�\�%)�������iPaII��\{�p
<_�U��2�v5/���ϐ"*��IfMwh�E3��k/+���<�����ܰ�K���)�S�!  �C���nL��M��ϯt�HU�WXY9��̔��HK��7{�\�{����Я��\lr�>	����Lw���C�w�w��S)���v�#�\1������� ��FQ��Rw׊,/k?���y��� �p���m�wm���V��֩�-���ŏ���!�)`�} �����&������7��p#�7��1G�G�$���OnP�ݷ��7_{|O���U=��E%���r7k_��K��
��
��/7J�����9�U�$�h�Ǩdm���ݺ��E���Q��~7Ǟ?0�ZP[��"��'>t�VY6��/{Tl6��'t�T��*��r�7{|͊�R�ыu���_C����-���@�M<�'"�
(L���Z����y3cv���2aAkaNv����P�ػ����9,�@K�f|������Jmr�zob�g�,�M�m}k
ʴ��d�K��¹8�<C�afV'Y�|L{|�UN�;�
z�A9��b�b�>�bwWqn�$����no��1�_1�E��Q�B:��vI/
%?!5C��b{
���S��v��q�@[v�;9�a>1��DS�]&Yy���(��&��g�#�I;N^܋�X$�Gv���:���Z���2oHYNnyy����x[�S $���S��bِ��(�3�L�X� 	��l+������u�×,�����d�?�Y(!7���!)0��D<�}Y���-W����<�`�&����ƱJ�:�*+>����J(�V��G9�k��v�������<[�����M��_��0�]��a��s����	#U�/	�хio���Zmf��;+���w�=�d7[e��;xR̊t�y��S�/�i���F�׫���/(j-J%����7nX��ٿ���f'd�I��|�	��#$-sK2�}�G�.�\�䦅nnh����ۑ<7=�z�PV�|L=����Ù��Ǒv����@bBn\�q���E��ǋ �����<{�<���ǧ�����}1�-JZrf�x�Q��]NY�{�.M��^-x�R(b[�$���L�q�y|i�F�5��^Ηf��0IaT,�#�@�Ej���^�>Ԑ�"S�|�ݬ��U��Q�Jx�Ɔ���56KS��7�6g�p�� v���RK�ky�uI@9�A��cp�i6d[w��Y!�T|�
��w5�Y�����h�2W�w�UB�-��Cϐh:"��\^��&@L+��]cKZV�qO�ؑF���;C��F!�6b�;�T~��`���@�+���&O�91����B�f@��5/��ύ�V}�i�כ���6P9��l/t��;�c��z�����߬�T�e���f��0�м��+��Q�Ѽ��o�'��z	�J���`[�q�Ðe��2�P1�&i���^��4�3��nB@��u��Y��Mi�/-���۴�^����T�P�k�U�z*��@ NGﳗ�|���֦St����Fߊ*�=�'ڵ,qYW}B����! ɕ%-ҳq}��L�M���`8�\�]D�p"��#�=��ë���,R�P���l���_�^J���ALR�Pȸ�X���XI5��8Z/���I�L���m5���|�ò��%�/S8Q1�4�~K�Z���E5y�]���nɈ**�rY`p��(H�H���w�$c��s蘏������e�SC�0Z���/�EMpc��� [���j~�� T'2{�\Y�iQ��sy�F�2���c1�������:˫iEޞ�ٯOx6�<g̝����=�߱�2�crn��m=[;��Ls���$���%���S>�1�/_)�}K���]A����	���:�l_4�BAzԩkP �?�(���즳�(0�
'>�F%&\�����K�
�W���4g̼�pP+�C	�@j~#gW��2ME����K��aJ�76��������(�u� 9&u�w��y���c[���40����� #��]��p�������A����s�|ٔ	G����G�(��D(W���@�F��/��a8{ �g��Uf�M������Wg.�ʺ����V�ҥ�x�*D��'#]�3
p��%l����SW8�h�̱$���t$����6b�]��#�/�F��Qy��HO\IA�ؑ��ǓH�%���5�?��ӒL���o,}<x��e+ӽ�W52��H`��D�3���R�e�1�������~�N':�Ni)�f�k�`����49�"�|p��we���u+M�T��j�qh���mU�js�f#�[���� ԆIu�q���ijC�a\
���V�>'B=AK��Lc���&!y���1,��oեw'�Eկ��MO�����B8)�~]s-���K�Ƀ�5��d�OX��k�c�;�Aw]�9fj[E�0.�# ���
y���#o���Q_	�0>�`j'�O}'��x�%{�]Ǚ���V��,��#F9Q[����T݃�Ӑ��j�];������l�3�XޕC»t���A��_�G��)�`ļ8�%8m�'��S���U���M�HA{�Cs�.���݋�b�� I3en���抨_ȼ�q�Lm���gx�k���/0��,���g�ަJgQ.)#R�AB-�H��x��@]]�����c�w�����5f�$���|�#V�m>�U���|��M�V���͇%�+��]쥶�8rU�?��W?��Q�d��ٽE�l`��׮�5#Q<�.� O�`��o��ހҜ�c+�nC+��
�E�	X�� T�I
�H�8���ҙ�rh� }��*�J.�qy���'c*Ϯ!��BOD�t��'��$%�TuzyK'�T4z]�e�G���$3Hg03Y,��u�By/�xq�ғ�y�fE�2"�Q�v����� ������uؘ�Mއ��匯�]���S �R���B��=[�[\���;b��X#�|c�;�sD��QltXI�[�k�zF>s����l=)���X\Z�!ad��ס�p���_(Y�͗5*��*�G*m�f/���i)3�Q�kj�$�q�;�������KNW�)���!{�qC�'���諸�1����W�D@9�����H&��7��������	��'��>$R��r��j9�CP���v��NAB�B��#`_���-�b0'|��� 9��@P��e=w2�s/&�'���O�� ahFL}�mgґ��x��CO���!K��
�+��d,>^�}��ؐȌ�w��yp��R+�R���f��,;j��è��H�O����U�Re�|����N���+�E�T�mF_߿��z�%~ʝ�K���lr�3Y�Ul+�hޡyd� �ӛ"*��!��J�6�Y���zZ,Z�̮�sm'h���)���T����� ��G�!�1���7��>��o��2�uR�˓:���1I�-%n@��<�Ϋ���r��J��T�;v���2��aI|Z��3��,��j�,?�%�Aw֗=h���amm��_b^c��G�YMD}k�o��7���8J�^fnS)���8a���YR��{W�N.��
��9}�|׽7����q�X�r2���wo�%Z���(E��t�۳�:@8�vdc�%��FC���{EhYݮ �q����L�[1�9���1b��Sb�`&�P�5�G��,�t�Gg��wIVX��lLX��G�إs�d��:��*�iN�n��yH�S�S[�ѵ^��]7��3F�3s�so}	z�e+uR���5�^�����3��?I�:!+
�vP0j� w��}��:�(KǗ\*��J&����A+Y�?+y{J�X��Qj[��׿�ԟ��$�p��/��w*���� �H7�_�˩���K���l�D��U}Q���o �������խq����e9\2xM�Rt���������~۲ Ю��j�A@���-7ɢg�U����dn:�W���?-���x�|GG���6Y�'w��?������B�="H�PQU+L�"��h~��o��3���]I�{"JB	��q�>��N�FWb���&<�oٸڑ���յ�@�},�|v@�r!X�l]�u`{�����N�(]=�$�ʘQq�]i)n��^	�lR.�I\��~�� B���-����e$Y޹b�G�CU�#���L�J3뎆�tc5��SqV#�@~���Q q<e���k4�fI[��Ai�cK�6��N�!�bu�eg�w­RY�"�T9h��ZW�b���g-�����`"M��^���o+\��c�ê��|،���D_�C�P�!����;���=hy�����;�4�T^O�2Z1�/Ľ25@���/�h��,Dx�2�n��6ku�+�OJ;��T��ߥ���X ]����� ��*d�⎾�\��ѷb^oKe�'^h{	�b�e${6���c�eZ���K̷�+Ҙ:`а^����I��*��u&�"�ܳT��R���y���X�(�+,����7z�/&�;1�GJ��7����y�t��������k=s�'mWؽv�ʁ#�<ފ���˳L.��QkM?.O`�	\9A�+�F�>Ţ���5ÆIh�F�FR6����Q���G�֋L͠�ȓ�F�Ә�^���J/7��2Ⱦ���m�T]�W�����%`�O8LY4𥿣�l���Py ���<n��*��Y[cy�_z/� Y�3��$�[��N�G��+�e�����ZF��.o�E�]bcj�7�[ij��@1�Z.���{W��Y�DsQ�:sT8WF�K0�s1����v���	)i`���T�x��g��ō�a=����Æ2�-4n���a�;�Js���չ:H�ۚ$�u�S�Pw1��)�K�9 �{�ڸ�	�Qʧ�0�_A����$�=P�)�?-nw�n���&���#
�nF@�:��|�ƥKO����J1�/�/�D+���	�����4#B�E�m�ѲI���F���7�pG�:����k(���[��uW6���Z�d��;�pշ��?�!����#�w�3	ј�8ǔm�U8����;���H��Kj\�������W��������ܴ< �s����MHKE��)g�xĺ��(�q	2�w@X����b�c]|Tp�Ūl�����4��P����O�Ȧ1Y�b��p���i/"3�<��cir\Ğ��l�����%A��
ذ?�E�1��u(}� �@�)����5��.H[��D�`�Ѕ葀낉7����~!:,�9izbYa]�&c5��s[4��W�t�A��A�u&Q��!]jy`֦Ò�U��s�Y��i�&H �U��2>����i���a�ޞ�}e�VV�AF�ߧ<q�H+�y@��KψJ�wbv��J�IMJ��M�}B�~x��-OR�K�Gv�<�y冮&�J���ƴ�clVA��I9�[ 7�.$7��Q��S�or,�Qzf�>�`E7 O�(�[��%v����jbu҄V5D���#!��[�� �ﺔ��!��~;F`��G/d3�^���V����p �M;�G���)�~���d�8H�'�D�t�l���:��G��D�.���1�{��3����`��Z�r��(�(K���[���-�~���&o�wp��cdg��z�9\!G��U S1�{d-]��c���wZ�ʐ����̵n�M��8�^�,m�%<���|�JJ��x��<��3Z�8T�<�9r��m��u?��v����l۩��ey��5���)��Oi(�*�
ޛ]T��ūI��#�lEZ�vX�H"T�|b�$��P�n���嘎Z��Jɜ�y�>���A�iK��]d�D��x��;��_�[��[�u�'��z̢��xbeV����w���H0.n,W���AlyJ-~q>0~���f�eO"�83Q�V����Q���4M#�Ș�bۇݿ,�'gN]ɥU��
�Rviڎ]�=�/�[7�ʓ��_�s{���8qRs���Q�l�IWkk��O>��!���L)�U��w��!wa���R�Gp�<_cأ�h��5%��ׅ�*(��fJ��^�83��k��^����n��fc�K	ٸ)̥]!��LCt�]���҃z9��M����WwQ9,�̊��H��7񕺕����O��d�T��>?���pE��C������Iy���Ņ#�#q���WU=�!	��|PU��h�w�/�/�z�������� <����mM���F��K�Tڣ�<�;Ņ���'�y|�}V���ӌ�/@�44+�mf�͍��A��gd!�}E����O$��S5��m��|L�~g��$`E[K�hu�_:�O�m��@��%� �r0��n�UR�hٛ�d#:q�V�}�����0��4�5����Z�^��8�'�������"�*Tb�[��:ȿʜ���ѕ�rH71{Њ?��MUIu�Y���l��-���@���<r|����//���n\�/�cvb�2�ƚaD���i�v�N����u,�w��r�xީ�$Yomhה0p�b��b�3M}:�k�5:�rG����/Ɏ	��p a�2�Y���{2��Ni44
��9x����͏غ�q�����wQo.�V͕�E�:��6E�:��rv��%5��Csb�{�
��I��l��'	�[�649�D1�S=Ct&ϳ���P��sίϕ&gj�3Iq�"܁�GX�,:G��d����5ֿE���N��q�� �.��S��D��O�X�Ď��3.��o�	��J+P��<xi������
i��?!�!F�n��!0E�L���}���#_�\����&с�ռē���+�_���7�LI���lx^�����Uok��ֲ�*s��C�_U�p����"�r�i�������U����OHo{���Ќ�J����˻�R�!�e��xH,�ttؓ���������<��ۍu2�00VjcY���c7$_�O{�!Vd�J��2���U:�-�0��s�G�9���v	�Bt/�d��]��i�=�5�PL��L�⋻#J�4: �l�a�����S�B��q�j��I������<qa�����3�B-}'��V~r�9����]D�T{i�t�=�C� 7(X?�$zM�q�ai��N��U�^Dg��AIW�_��D㟻9������@Fo=��iU����iJ�m{��N�5,2�SL#?�{�]�a� l�����k﹛Iv��A�kkc&�R6�!z�=��!ÐJ��T&w}F+Y����h��W�;���A-����Fyb"��^)/S�+7l�c�L�ŧ�v؇�ԟ��Ca�!#�,��;i&�x��ʖ���6�z��|UOGl?1렦�8�O@n�?/��<��st������)��6�ѕ�5*`;����Eʰ��>���m������{Ɉ���De���ѲR�o�T�'C�	�Q"���A�k�#�e�N^�F�b�-�S����P��O�$��e`~u�Ĉ�9�嗚�\��є��������~�ː(z`�1�6�PG�t���bs�mYt�\�,�� ̀=�$�"��W3Y������W�t�P�'����=Mڡ�`��\�����%��Y���3�6�aņ��z4R��°��t=��c&�)�lLH���n%�������/�����G��4:m+�e�2h��(�1%�x�8G�H4K�S�x���&:y��՛ė
n?�2*J�|YVv����V���n�NA�$t!�)G�$&�O�}e�j��;Z,��I�!EC�@cE�⛖�o�#6��8
�/{�Y���Q�qs/�(F��H�1�j
��tᇰhJi{*�ςx��rgB��(zB=���g��2K�n�#�c�];`�sDZ�Tq�֤��bkS�ż1�'�)�|�K��G���S��	�&!���_���A��Kԟ��P�S'?h���	�Z����N�
�3DF[�������mK�e[���A�*O���)+^�K	��I+�#7��#�����AA�\7���wY((��*�%eu���[>�]������Z�ͺ�3뭤5#�$���0���v���q�}5ي���ɊΆ��}�й�R�WF]	�_o�1ՄWQJ e���˔�M�� ��oVg���X_6��m���'�����g�]p��lUs!���4��k[�9�*�l:bt����/}����~�|\?��GǠ�	��%܅���*?s�����1��}2�d����3x=5h*fHV� D<���~⑛�����u����~Z�:�yciu����8��捡�n�4/R'�2��O*��4u!u�
źj4o��x�Uz��s^�>��]X��� �Dk+ˋU/i�şaR�҃X�VPYx�sAAB��6(�Piy0�'���%�w�����?�ME�-�
ZB�hp~��t-���K�!3�w���!k��E؃�!�c'��A�a�9��[���.ND��0�� �Q�o-�Q����&_�` g�O�S��}9%q���O�0#gVP�B"?}#�ή[%ý������)� O[;<��g{��"3���T�;��%����ۏ�6�G_e�)���.f�8#O�'Q<�r���d��m_�6".1`݁\K�V�@3�����CǨŪ�'z�ǩ��ol�a�4YG�a���� ���@�g��A�w �>8�.c ���]0������w���K;?����̻ӹ��&�mt�ڀ�\|6����O���!�o��޶wg�r�ys����?n�G��}��lVm��@;I�$�U5Yܔ�$�jOt�<��ȣ޶�Y(z�$�H�^�E�t�X�`TM�Zþ♡0�_�����n�R�Jd�uy���?�$�{�x�gDv�9�[od��c���M�p-8';��z�w}���#e�z���D�,y~J�0)��,l+�����ye�q�j���m�f�*�"E�|Q�V��S�J�v<��wa�`e�~��� ��>�]�p^�	5�R1�A�x�t=Q �[�`�ұ��eՈ���:s��xQ��I�r!ktp�>���-�T)�����8/ЬPa�����N�p�K_�ɂ��e5 #U��2s*㗮fe�x٬t3��k�Lͧg^��e ��9K�zp)�~	!q�sCOd��i��D�Y�`W2~�97��� �H�#�7,�W�LY���ۯ���9�>Z���h�� �C���H�ǸDј���#���4��Xː2�#�\1u���ӋGw��/�HS�6�E� �D���m��b��4���~��^\�W�� ��
����}�.�dی7?��و�1�HL����Ƣ�l�����0O�~����&|���Y���_�GE��ǽc��_��q�(���[�P���M�M���U��ghԵ/d~�����9�@�!��՞�[Z!��'k߇(P�=��Tݕ�Фt���W�	��"�7�*������hG$uH=���c˧)-[
�@�^E<�V�;9؉Ji�@�ģ
��vF�A22�va?�2�ě�	n�����,5C����~��t=���umc�f���bԺF�}8M�P�k�U���2�	��$ꉃm7�a�мYHA�{3N��j
K�9s*f�s$����q�J���M�RA�oit'�0��E����>:���v�+D%���CNI{�������g���4[���9,1X^�S՗&
�g�k�N�{�*�%g%�I�� ��f�X�i�G'�%��yd�.���h�aVN���o�5	�zS�m�����SS"���c3�����	p�++X�wf��X5��sŇ��?���!a�۴l00 �(�)}*����9�����o&�wF�7~�����+�c������GH��Xt�3��-��YIF7���(���i��>�x_��a�I�=f��6�6a��mU�������o�(�L�� í.˖��G�eo��xC��t�7��:���6���g~�h
Ůk`;j������U7���
��"��dd{��+ϐuq-D�)�n��G��ꚍ��]�υ߀��iH��B�O=XC�PG�|LN�
��5H�O�ؑ�&��it���B?f�q�6�V��Ǽ$��h<�r����|�nn ��}"=�,�0r�;����]��{D���x4Io-(Sa�$ծ��@�q�ji�����"^�U���IR���4Ѵ�vQ��,-|�����T�+�}�'U�s[�b�CJ����H5�o�S'���n'�A� g"B�c�}k��I��;A_��c,?6����z'!����bw8�gY�����h�`�WBL�&f-��bϡ�6"���^D��;�+Z�c���Ba�؂�i���C��!>=|�>>;D���L�1���19��
O��12{ĳ{�@I}/8���Y'n�L��gd��m�6�M��
��;Jb��KW��I����f����;�����>��X ��gѭbLodb'�=�	���[/��=16>e�6��Ab�7Vo�&/��tQ���	�Kzu\k=��߿�@�����ѯw�N���A����z��5�1��G ������'��t���rv�;�)=QA���W�B�@�Y�r����C��.��IGMu5�`��\�zˡ׵�tw������<au����Rl쿁����|׏�G�D^�L�/6�IK�I�A���/�:�z�˾��6m�y��Z��c�x%�M8B	4�T�3���A�yƶ��4	nz�*�#�YQ�?���y�ȑi�Y$��i�`��_iG��@�e��TaQZ��R�dO�E�Dc ��������K��=e��{͕�Y��Q���s
T�F@ީf��1��Z�,�D�k�i����J�+x�H�g}jD��e[=�w���2!n�d�
Q;;�sG�����H���6�+�SoZ�1�S;)�+�K}W_P��t 	���K9_e�bA��3���P��q?�X���_݆|�9�
X�=Fv���d�^�eK��Q�(Z
�%�*���v+�5	؆z~�#��6������<�Rr*/7g�Nˢ��4�(e���˲u����|������d�I�5�Q눚#KEf�i������#�˦O��+�����zj���Ɋ>���	W��Pq���L�[��� @��\�M~�����g?�W�L(���(�m/,û�;��9�]� Pp�?)l�_Hۄ^9����������b�����/�,1�!�ə�.\����"R�D�y%wu7� ~`?���},��L�x}��y���=�nk.5�uHQ.�D�X�F�@��+݉-����-�~��p:b?�ip4n⿜�j��54�л�	-��3��wP�u�Ge��j��~iU�f~s9�ԫr�\_� �SV�����i���a��R�3�)V�<0�.A<��]O�����yK���ꟈ b�wتՀ�DM@;�O6Bi8�~�hs-E��K� ���=�Gt�@H��|sc��EA��9u�i[�` .����8)[5��hjo���Q���䡟K`���O.�r��0P%l��Ǫ�듭Vk4W��"#��[`^��%֞�ģN�{?;�7G�ڷ%��3�@�Y����ӏR�G��)�����8��
'��C��eB��tɟY�q�tH}.0z��ȱ�1�t3tA����P���I�dl������|4ĺޜS�U����=gb�Ti�?��:P	�N��^
]�����[w�|������d�Ӕ#Ծ�mE1���.|��
k�V��DQ���
9r&�Q��g?������k��bl�P�����_Z�5�Q5��O��Т�����ۍ�V;���/��eE�U�X��T�C��y�@�K��dp�����J�Ly���8ް������`D�aF�6�	��2'%9��k��'�PIzBlH��MeLՃr��gSml�0$��,�
�s!3y�� q4�z�|Mf��"�1^Q�v	����1G;� ���Y�e�S��]6�]�[#�dR�t펓5�=���[�F�=�W�� ��>�;�su��Q��QI��kO�>$����uT)�7��-�X�X�a���H�*p��|_������:5o��;�x*��mf��T~�3p��k���BD��|��0�K<�)x�!���C*�:Z)gҹwC�w���W��M9RԀ̀gpH�zt7g���ҍ���eMX�>u_���V���MCD���@�?I.�S��#�'�O�������:�ya��χ���fwCT�/W6O�����Tz ���#m8���B>�L���^r�0�{)����}��M�=ߌ� ���c٣<P��*���.Q��L��Ʊ��mO���20�7�|5��4�	�(.E��|�^3T_�JT�㱲�v �I�(Z��v�U=�?h��d���̰б vp������2e�+��Z���",'y:�BX��X�TX�1��\�@���:ڕ��[7��S��?�ƃY�uÒw�˖���ɠ-��3@��~<(QU��~�e	�������2�v�� 2��*a:Ni����>��P,�.>��'���*E�Z4tm^5��Qb�e���Ms��kv! ��>����e��(�aҎ�Y��U{�ƇN߬U
�k9n�4���\�N~0q��x̀-�so�K���k�E�>���h:q�Vv��'%+�C)P&{��*�9��br����[b&=9G�k1��S��&En�Z6��毅�Dg�I�6��wCX�ƜGb��Dy�~�A���[�2N����Ѱ�TSq&�P>n�N�D^d3�/���	�!�+w��t-�/.�����DFg?zh�!|#Q��J0�;�(�!}����眗v��LA�&��ղW����+*�;�)9&�Bg�r�ѹ�H�}�
~o!���(X˒`�-�9��_�C��XR��_��n����KUNvͽ�o1}��F,��;�����q��P��e
¦x>Tt*���?�H����2m �C�����Tj��ᙍ7�A����=[�d��%��j���Ј-ߕ,�i��GXĨ�HX��x�X�ZN�DS��}@=�p�PB�L��	��A'�j ��b���nb�,{B���q��Y���w�W�*��<g���kTħ��3x�:}����rR]Ԯ�*W]:�!{�ܳ�����{(N��$00X��>Cq�4i�d����^� 8#[3IMȃ�}��1���[��[�����1.�~U�Kz��r=Jd���
c�5"�S��%�ܠA b�J����ke5�I���Aڜ.c��{6Ph��s�q!�L��v�<w��Y����"h��sW}=ѵ���-�
��	�"~R�^_��z +�g�c7� ��Q��}���U��C׼Q!Y"ȭ;x�����EL�,��e��O�?V1!��.Pi@$y�/s���r i���CA���r�6����	*���;�LW�戺�������Qm�����q~j����-�Ѩ��o\��'�XV	.�����Ǣ&q�e+>j�<]��������!h��	u�����V�u�ݎ�ͥ?���+��ހ��d&��W-��Q�A�fz�h1�,�CG[�=�h�.�B�t�$K�qئ�v�f=�ε!�W���j�������� i�8v�M�`�\J���\�������)��4��ȌR��t�b���J�L�_RfL>��$�����������k/H��5�S�ӻm!<��kÞB�%1B�8=�s4�ܣ�d]�\��y��C�z�7n�)*��gYL�<�p1f�4�f����$�~���5������e����>�Zw����E9��c����T��Y���?��-{���Y1��Q�Ms�|F{W�j51��χ�G�&�yi��#���wx��ig���^q�=��t�~�2�Jn�RY��;&,s�B�Պ>���J�U�S*�1��)y�-KXgI�ډV�	�0C���2_ ��A�+�ԕ��Pm�?��1�?e��f����h
�[F�����ɪ9��K �|���� S¼U�+�-d	�s�k #Ӗ��zo��U�7��_b7"��#�x�m0f(@a#�tu(��۽ڏ%��l�&�Ͱ.|�c��#�<��8�|��,��������ـ���U+4�������Y���rW��X,C��gT*�M�I W~�AC.MW����g����X�����V�Ö�L�,#]MZp�"llo�?�A��i
�����kK����bT0C��C�/3d��=D'ɴw�\5w����3���%�'���R?)L�8�z�gD�}(�Z���?ө~s5��\HL��D�����{扨O�s�s~��:�$�ik�hr&�WNˡ	Ů4%o\��v��\���*u��kVj�����UpP�s
�G��� ��}��$��©i��kaH�Q|V�{��BA7j߸�6�y�Ayf��j*���nw�-�CvM; y�^�B$(>~�O�-�Q)K_5݃�:��WD��;ؼ��Oc�fA��*9���[�%{.���f�H�A�#o�݀Q�=� �`�&
Oi
4�,?%g�Y���$XV��Sv�#���[�ԣ���п�o��OY;wSh�m����3\��ڄ�'W��D�^�YGՒ�)8��$��8�*'�4Q�Ey���j��D�/z�.K�"�wUd��x3Qɕ1!d�KP���|^Y!�� �WTZ����Ě��Z��Z�g�_o���~Ŕ4]J�&��,]f=���Cwkj�������߇��o/�w�m�@�ߢ|�!��Bh��9������KX���6r������?$2��Pо�)�lLT8�� :ך(_5��ͭ3�O*B�[�b�쾫�O������ԯ�E+VPX{$0T�+�4���fr���v��ಎ��J�Zy�{���Ϛ�V��G�DlF��7�"K�9�fa�'�9�z�������e�E��M����M���0m,"4��.��y���q�?˓W�f1"{��Q����	7Y��q��;[��ˢ�4a󇎐D��M`]�f����R�*ݎ��y=G�[��|�x�Q�D���I�+s0�Q�uI�	Rk*�>_�~�ccL)�ؽǈ�F$�a�X��{�p_u_��9:(5�iז�*Y%�f����op3KkVE���a�~�p�wF~K:,)�9!g�C���p��T���yF�\�W�7�9m�����uH��*7�,n��l�zV��u��	�>�N��^) � �C<u��~�Q�:�_��+S#L��j���N��[���ၪM?���1Bw�/D�r�;�� ͇�8��m�|���p^�\9���mB�K����U�h0�*��}'(e��5ߌ���e?Eپ�v�>)���������Nƪ���O5a���k龽a|�~n�r5�ռ�E,j�Y��_K���������̻<��tU؅ph�IVd4�Ӈuб�h�6o����fCZZWә�	G�'��k��� �sS�T��n�ZH?�{\��B����7B�E�p�ƞ��u>	������e-�y�@��t<�k���4��&[�6P����v�cS2h��a5�{�z��/��0˚,+:ɨ���)����jmYj�AafbJ�����M���kQG;�#��R�)z2� k��$�a�l>Y>dF{×�N��
��~9i�?�)�ď	�q��,�d���o�BE�fJwE���G�r:,�v�ss%���Cw/{1�X����]���8��[��9b=K1NC�S�X&�{�����\���g��?I������BXkC�G��C�ߘDy�V���SN����e����~SG�������I��ğ��3_xI�/	f��+��L����#i��r��Q?5<�!�nδbJq0ֹ�c��}`U��[�mi!��#&"Ď�-QL�"`+e̞���=������J�c�+�������c�������4�h_f1׷�s^W��5I�0��U��͸n�o��`�,T�V�Э����L�Q���e���x9��t�V��/)���ع��.��z�� �j4`ݙ�on75�����X(ydZ<s�����L�-zx�d�0G��ƚ�r֓<Ʌ��գ~۸��=���P=��L䈻Tm����a�ݍԳI�߆g��Bu�q��7��2r��Ed�<���Fջ��}K�Y�r�U�أ ]�'�{��ȳ�bl"(IE$��ܓ�\q".giL��|z�^���T�IH����IX�����:��r����k��DݳslU�C5�jWJ��%�G5�J S�I��,�V�wp� ]����k ��Iǲ�AUeBc��6�;��Г!������w��Y7�A�	�HhdF\W�ʵ\>�-�c��W�_"9�$^z����s+ȕxcr���xb��x�U԰,C��n!t���qI;�P�)y��g���'������Oxه1<��ĩDh@��g/��L�kdB��:H�Z�$6ץ��ih�E�;�V"���氜3��O�t��(j���(EҢ��#Ң��ѣ�o��'J��	I�S�Q���'L�$�e�e�7x��*�҄�<�׽���۵�u�nu�p��ȋ���'�/n��̽�Dñ��c�|ӳz1f%�'5�G��'�#�R�]t���L^g߱08=��ǵ� WD덪�\ �#���j��1S�s��M���`�Zr\�ݴ��5���r��8���2 �R�Iҁ�� ���z6�zfL�>A��8`��aLPEb��H�/���߾��m�ȋÝU�ٯC%�V3889s4\�ѣ���w�Oy}�UΖn�E*�YGo���N���H��`�$y}^��O%��O�� ��e�
<�Z2����IE��dc�̓�G�7��֭|�=��{C�gYL1�Q|��s���F���*�1�P����D�ǐ��@/�x}:�g�y���5=ו#�x�2|��nGn�3;�Y,s����%թ�ǂ�����S���1),)���K3�^���$X^	�e��d_�[7A����PH�6?����/�fd���j
Γ�F�0G��N��K;vۭ^������+���	�4t<#�vh�YUL��#��2�w(��7ݳ�>�6��K�(��Gx�u�,���#�n� �'\�A-�+���>�#�������w(˔�Z'A�����w��@��0�7��N%���WW� ��j�-A���; ���|J�M�ED��Ug��k������Y��c���qN�N>K]�,p�9�lf�����N�������ӻM��Vb������/����������\�T���EǺ��%��ϝ�� ?�Ύ��=΂��}������59�HG�DMV��()���׉#��NӁ~F�:�*�if������2��$ 04�-	��&� �����u�Fo�je[��/��U�Y�s�B���s��l ���<,򋆼i��=a�p7��4�V�ZI^�A20>�⍗4~�y����	!��_9wN_Jն�M6�X�7�B�7�~�V	-;<K:oʃ(�R��`"�6�C�2��cXA��p9k1�[�
.�d��( 1
�b��o^TQ�N䗀�`���O��I���%b��`�Ya�fV��8�A2#�[�j½[q�к���1�;2�!I��37�|���n�� ���G�Y\)S7a��*]8���'�������H������.flp��c���L3��$�̿6�F��8.S���/l���K�qr������C�ŗ�g<��#�����������g�7]����K�w�q��|��3F�Z�Jl{JO#mE���u�|GT����m�TQ����x�3�(��r\����-:?�	��u�D��l�w��ѓZ���5*�^��lO��y�$��ʃ��⫵8����E�vXvX�T^����z��h`�Zҧ�g��F�iJ5�y�z��z �U2j��(*D�JD���įK1C[3�a+�'LCz������eB�σ(�K��gO�0,}h��
y�I�q*ڧ�2�fl:�"��Q��d����]�V���C�������哅�]����t�Rb ��/(=�1[���#���E�
���4s�c�Q�I��k��>�����p<)�����y,�a�1�>B>p:��_O]��Բ-5g���d*��f�A�J�03&V�k�tO�x���y
���|�K�0)8ʽ!�j�C�rX��;������Q�j�Wc� 9����v��Hm��7ݞ�&euCD��]F� �>�]�����B�Cw�"����5�-�	��#M���l��#:�H��j֪�Κ�Ĵ�w���/�q-W���E; ��s�mnw���Z��F,ڏ&����q�n�Cs�e5t}t��NیHQ<� ���ْ�ѹG���T�SIǂ閧��|O���?�K��c;|��|��
�qE�>��Tq�_�GY�YEW�7�����Z�Z��Us,�h���d�_c�BZ��6Nɩ�n-ˠ�T���Z������'/��߸�����TN8�5�1��1S(C����7��W�+,ƹݥu��F�� ��Xj^-,a�@��&<ޥ�ljɉ�c���0ǣ��&v�N�2Qa0zj��kC�:@�K��,�e@��=D�d�����YmT�����b..���MiT2k,��^����uJk5�˃�K(ak�Y�%c{��ANU�G
s39d߆ׄw����q��q����oZ��IgE���\:�'�v�G'%!N�C߽({l�zݵ�N�X��:*[ؕV9}��1��LS�Jc&����<���So�;s�gV4�I�j��m��XF�G��z�HtA����њ�N���"�*�S��X��s��D�p����3�!���	�+�В�(���e9���nÇ���?�/T!��S���0�W�V�}��"�﷗�|/���&=oըj7�\k�+�0��_���8��iϠdş�~"� '�ײ֞ʒ��/�j_��M�L;����U��$�X�k TU��aͳc�o�=¼K��q�#�x���'��v�e@��x4lat����-��r�(�������#j�������7����;"��sd�̌����A�-{��_7DG�D����֮"�P�I���	��A}=),�P8�YL_$���q���2�X���$�톢X�B��qߚ�g�v��H��`�<]g�!vc�C��R)}�=��r� ���<�]0�{���)*b!(D�$�A�q�Xq=�i�Sr�Wq6^0��YnICB��E6*��X��U��Lh��i�o�N��U�[��s��Jڸ��@�d5��S����gǼ�`� Xk��t��k�0I���A�M"c���6�.q�*�!��8�,J�wi�vYR���[h?�W�7���-��^ϲ�"�y^�ےW�+���c�����N�s����CM�/!��;;�I�d���]��"�v�O3�}1W���$Y�@ڠ/�Į��_m��S��ܩ6�����Q��;���L����ɬ����b�C1J�g�� ̚�	Yɢc��ўRDoRX'�	dZ��̯}̡�d�ea�V�2�fHŶ�?wdW����ېA�Q�fu-#��ÑӄQ�<�H��� U=ɿN"�r�德)uz̃�"'Gv��ޑ��xy�t|�j�'��쑝="{ٵ9CW�$�q�y��t��A�����.�MF�W`��"\ $r�Ҭ�����3���!�m�5R=�߁���zz����� L4����������F��EB/�����o�8�]m!����=�%g�(834�J�d������y�Nb�0�%n+:�*��2YBl�&�u��o��U�$����d���� �e�q�eY�Z����|E/��c� ���L9w�7v�+{�0�Yg�Q��Ys��F��7/1�z��=�.��#9i�B�����xX� g.W"Ŕ��=�T�ӚR27�zn:��O��;̭�s�����������<�S�ػ1D��)o�K�F�~�ڿyA	��U�\��_�ۧA�ԋF�P#;�?T���u^�Ά·J�
��Fǒn�v�%�.nKvfn����	&�O�+J9�	)��,�#�vy��P}�P��-Y��*�7��HYݬc�T(����~Tu^�m�џg��E���S\'�ͦ��<"#���:䠘rt���%��������v����r�4���¹�� W�v�����&��Cz ю��q�MOT`��7�gP�źD�V��=(���Lm?��pg]�-�p��l��۵�_�
�ٱCQӖO�XK2b��r���/�2������6\+R�س����C%H0���j?�pA���DΝn�}K���Z4��5�T�HB�D�#��w���|���V�)��~F��:3P�ia_
(�߿�5�?��4°����;6�H��uE�v�rj ꙦJQ�Uf�}sʛ���n�-� �@��z�A�SiJXa>囃�8�V<Z���pA-jn�n[ŗ�"�y�,�Ƀ���w��Z�Q�AM1����B�g~�}�-�F�K�ǃcE�卝��1Xf�(c�A�^9�v[g�.:��ϯ̎����oIkQN�!�`�f�O�@��b�%]n�ǻ���V��-�#hz�[!U���rе֥̌�W;��6.���Ӗ3��@=�]���c�dPGK@�)n�����8�Ry'=���{ (��ib�jG)�='.��mέ��G�3ǙT�g~a�ATf���'���J 6�Mc0�x��M�Z�&����*gs8����\*��j:���l]�F���s�w!�z�7ƢN����-�%�o�G�m�ㅀ�h|���븃U�o���ξ�;�c�.r�c����m?������_�*lB�\�F��%95�r�%O�r����1�"�c�E�ǫ��E�J�2Ea�Xq�pT�]}ê��~[�ի�B�4��#�Jжy���Iy���A��)�Dbo5��~گ�`���\c'�l?zs
��{:e�o�Hٻ�<�J0�q,ؼ���`|y� �q���՜f�"���Q�����b'%�q�C����ꪞ�Y�.�]����u�R����ܞ==�_[~uٓ�~B�z� b�[�s��-Q%tI} 3k��>�`���$)�z��>z���a?]��(�pc_��ǽoKK5��L K*�2�fѯŲ3�<k����E�t���-��K�A�)S#�!]�C�~�_dҊc��ݸ��>^Wq`9�@���]�HH?h71U����pP_�+
��X�>ƌ�T.r��AC�����1<�0q��d�|#������D�u�U��H_��~8ٿW-wT�a/���H\ͤ1�M ����Bm	�&��,3�t�J�5����s��n��}]|��ӌ��;�����m��4�����Ǝc�����ۀ2O�G�����)=|yq���Ü�KEEb��O@�_�{�����ľ��f|����)U��h�]�d�8���^|�Qꑩ,�	�{�����)Z�`���G'����s���A�T����4��&�ðە�"�7�'���/���O!u4S0�\e�˓j�-�hr@���<9 �'����m�,1`�v�v2Z�2��Wa+@5�0�f��p�f;�,!���c����+m@mOl���b��؞�D�M��zk�a������p����̃Y�Da#�`Y4�{y��N��N
�& 9_
��}ԏ��q+������p�oU��͜g�E۴����&:���v<C%�ŏC�${���Pv-�SI����[�}�9�ۢ1D�8S�\�&������}�����bg��I�4���FX!�GJ2�8o���2��aN+͋�[{�u��S�:p�!>��?��U��3�i^P�	\��+��H�c_:� o}��W�U��?�C!�d�X�0�;�ς}�vf�
�o�#���}�h&X�w�#�N�7Ԭ+۴����1�3�F��-��~`�{����y�٥��1�s�*�_$uMT���M�д��q�����U�?ͮxqoB:�w�6���������Le�Gtx/L�t;��p�V�&����=��ԝ�Wa�jj���~�w7� ���w�ю"ydP}r�yJ��|��-��E�Z�3Gi#�y�X��c�ˮ���3i�.�=Ĺ�P3��L����$ݙ�i������ ���)�B���qڦ��-�Ǩ?�{��<��$��6��ZI�t}�E��zr�����+]���{���d|��w(?)J$At��,:qXVi{ɋ2�r^k�����I>���B��b�p�h������@ɮ��Uʓ�θ�J��7�[q*5��]S�����V�o� Sn���[rk�ޢI�\�AKV�cm�6BA�D�`!�VZ���.w$"DYmB��hYh�}W.8���-�u �ӈ"�=x^�w��>+~Q�c���Ů���nb��f��CI�!���$;�b#��dʝ��5\�v�lO�l71r��ğ�J@�d�/$�C4Z0�T����@6~r�zH�q;6˔��ݧ���x�s�����^<��}����D�Ԣ��aљ�yom�?'�hv	,��G�7X�'"��e�a�-�����|�r?Žz6R�k�"�8�u������焬���1u����:�~�M�׾�zg�����Gl�{���&�vt���ʘ�'�=�#�	��W�AZ�,�w���_��WC�n�730�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���șs	R�KF�Ǌ�pxC?�ކ�m�$�������D�29쩑�G]��f����qm�O�2ڡ�?|�>jGG�ZB�x���;�_�K��@T�V(uz�;G�7�L.���S���,\b!��IeT�������懎'��3��~�K7$�!2"�fyŻ���r���������������C
�P߯&��"k��������;i�M�'Wl��s��(��-�XD�2�����b�3VCU%�'��f��k����D��z�0�1
b��{�Ug�tjx�Zg�<�(ݶ�I��6��$i���-z�w��'�?!~�0�%�+ΒQ�Y��*	Zc�;�ע��D)�.@J�\lX�V�ۧe}+(���Z��?�)�3l�]x����-J��쾧��Ǭ���9�8�F��B�B^���?c�Y9(�F�UH%/��ON�ou-������S��Ҳ�][H�\6�]�H�X �N!?���hG��	��[Ո�?ԛ����l��5�v?�h͖�}�v���YP�`9T�Q��5�j�����r�U��8Z8���-69dû%B�=���̹7�~��c�ĝ��~�?0"�p^>yn��V.�P3Vm�B�܂v�m��0m��f���D4�j@��ɳ92h<3Q&���g3j$��w�uv"����h 4�2/W�!o5D�y���N�6.���Q�Y9��.R�x&^�ɘYV/�w���ΐ1������ �b�[��G���Y=%��)�+��֪�3�p�J��q-(���?Q���R6(X&uq��2�g���ϓI�%6E�R�'�ϵ�_��Yqھ�z�C{��I�K��,LI����Il���G o/���X��6���KvS��B=��-�\r�%�1f 2\X&�}�j�����IC�J���x��(�%췯�s��L�G�QE���M�.,��))�Fď��c����+-�����a���Q��K�h�>ٵN�S�~�Cz�������}��f[��Ǫ��lm�L�z
C*6.�66���f�3iK��x4UP�)������ar��װ-8�(�Ti'�:h��Ε�΂�h����小�R)����<+��p�����R�|	_?�^��\g����C>��c;,5�m�@��t�(�&�glb��|���AC���]tg)YC�(l�>g�VF /n1A������������� c�$z���?�%��ê�3
y(�vpɶ���_��ϱ�mJ,s*��6u��(5$AM�^��)��: �޴�c������]���+�G5�)��˺6�9���p I�3�ۅ�чgM�d�ل�X���jd���3֋
�$����d(^��7�N�`�E�W�S������U�5��dP�A-��Sn���`�E���W���p�Q�]׺�4��&'�-���{B�U���{�\7�ň����dG%����>�^k~���)x5L���hprcY�旘ޔ
��V3�k���5��R#�Q�S��An��:ϨҖ�۞�&[�(��	2�༻9&/�SJn��Su��{��Q�:���li��b�@��q�9k�HFH��5'�2FȦ�
�USZ<,��-�" �F�%� �Z�qg=mfPO�o�_����"���lv4,
� ��|V	L���o5)�t��p� �F�I�>�
�p�|��!õ�����J�6��H�7A�}I��a����
���6I#S-F$�4��>ƻ�z�� ��0H�"�0��#d�¨��u�]r4��3�F�>Uex0��U�ƹ�%ɸ!D�G�1kW���]�� Y\ϔ��Δ���ic�X�- ��UQ��ct�Y
�;�)䕎�5���������n)��h�����gr�wS�����ܢv$��U7�>@k�I�۱��|�o��ʱ���<��ժ�P�>{/�#�{�PKo6�$�?��9N��?:��z�'����he��B������墳�K�*築ʫ"�VKN� e+�M*��7\	H6I	�?�Xv���I�Ơ�W�{��U(�LEY�m���?0rD#���纈�?�u����E�Lo|��[g��5yԽWt٦�%��3�#=^����I~�j���տ��v|�n}*�F�r�s���Pz6 ��ۡi�a��x��E�5�be�M���� E^�%�Q�H'H����Z��;Hc��hC*��k��䒞mKe�\��(�'�Zr�ٿ�$l4�o(�d	��ݒ���ec��x��z��8@ ˁ�NB�{��vi�YP�F���%Q��+o����"��D��S9L���C[?��\P�����@� Qi�?�g�h~��	.f[ST�׭NZl�x�5��v\�hr1��X��( Y'��M�ң�>65�)��RT;դQ�~�5�"���8'I.M���sj�R�>~=ZzN�<I 1ia~{U���z��ۨ�߸��K���&q��#\�$mVv�7���I�vj�.W����:�,�؜�8@v��r[WC���ԯ��< ����qb�����H-+
�VԲI��H���>�G�3�l����b+������*�l�E�3|�b�_BoR{Tn�Yw!g���S*�A�M<�a��p�������F���4��7���O�#����#F��B�>R�ۨx?ܦ�6���?s�.�z�ѿ4���@��b����`0m-�9h�A嵼�c�5���ڣ�xz������B)�#⨒�?<z9!s��n�����g��<CB�!��¹JTsh�C�����ֽ�&��$p������G/� ���i)�*9
��wȠAn4�.�辣{� *�T3�z*c�H�b�h��Ֆ��E���)� s��R�۷��4d�DN��dc~�t*d����¦��ڙEΚ�n�/X�b�����6��l;y�e��j�;#�״t/�M���B��"5�\��}��O���I��	�*�H�Zؑ�ݹR����`Z�i|�Ve��5v��x�^[N�G>E�<d�c3X�-�k��l��2TY���0�"�O�I8x��z�k�`���x��Z|^dEi5�t@�x����
`��i�+[��ʖ�̅xE|��
�Cej�n��lѠ�i��?�7=���?�����,.%�M�'���t$�- q@̰�������'7,8���@WҾ�e���ņ�5Z�K��%�>�#����J���6\��R憇(�k{�Y�D�R�=��/7-�z���2�X��u%�����G���jM�'୕�m��riܙ��=K:�#�=����]�r2z���:~Җ�]����q:+Uٟ�W�L�pM�Yq���r�"�ч� :��or������a�.~""fL��9u.�&x#}�f��~iZO?��aB5ڦ�:3"����R;���<�d`�*u�Ӌw� b�TP\HGw���S;�����ʍ���L��^�ViF�H���mY=M���9����f������~��̸����������p5���\�^J��z��S7 ��\M��UM�ۈ#�\�AWS󀥒�ɐ����6%��)2��r=mA�aV�Jk��������H�����[�X��	J���V>�3;$�h��r�BB��\Q�棊��(���ŴG��}yЄ��<'�E:յE{B�"���Pd
J���m�^}D�`B�>pO@>N�|W�;��}
�
R�Qo�X���ջ)��d�����W���\C�©
�����l1����f��d^��	.��J�b�17�Ey���j1�Q�v���霂W���)�Ƕ2�����;N��������Ɨb�k�������]�} ��^!�&���d�=�aS�%��	A��r���S.0?��P�Q�^��\�J7����
eo�$���n�M��N�Y��.������i506��9Yզ�U��7N�|��'��'#0��:�s�ku�
�=4�"�V�z�Ha� ��ۦ�sX�93o�������·Ս~�v�:)���X�{�.�Jɻ2Ǹ:��G�2��m	�v?�_[1�M��_Χ/+�_��q< k��~�H_����[ԌO�b�ޘt��~�����bE���W
�*�{��I[�M��b��o�(�n��w)���:�6*��5��<�Zv�v����A� �owNK�| 7ɋ|�k�DQV��s��oe$)cp�$������惙?�]�Qf�I�3s#����t�+|0
,�Xނ������u ��8}��|0+�k����}�Z<%�GF넌8m�H]$T�^͞)�M'�sSx[����>���s &�T�[�*t�`iV����[��MǤ^$wC�����=�}Z��7!�6��1or6p��z�dR�z����� ��$~���]�sF�:����Ϲ� ��%��A�
ٺǓ5<���EF6�+��X��Cwt�,�>X�A�������D�j~��- �mL{��,�|9���}2���T`�!���CEm��2�ie?k��>9OhG�\H�M\�e_\e6D7ɫ+�eTܟ�uI�VG�xaL�爙�l�{�b!2��Xk�T�M��[\O�6�y�������9!a�f�j�����ru��^�� 2ˮY�\�����@�߾j���J�y`�������Mv�F�?�բZv�J���-�;����<�z�LbX�C����E#5��ѧ�/զ���}��0#�b���Ǥ�ut�3�.{׼+�݅IF�Z�:��y��ֆ@�{׉o�JCbH��!�a��|N���-X_��p�w����ki�Z9�[�<ځ�Cc��d�s��g���(N;�Gyy�p�νn�cIl��xR2���Bt��=�~�p�i�\$�Kֽat��x��t�=#���u���R���መ�x��@�/]���^�[{��H$�6E2� �+J��i��M�L�s� Ȳ���$m��։�	����tX~�/=�&���_�6��kß��B����(��.~�*c�v�ˁ���"�T�Jy�Q��:�P�ǖ��5���g��8��B�Jz��� Tj$\����2L~���D�p�j�]�w�4�v������ ��2�V��D�h��O��f��N��=�����\�F]��Y:ºhf����1X!���d���?ܿG��Y!\g�O=K+�y��3{y�4�1�c5}��>��Aj>M(@<��3�K��%�8ǆD�����[N6�@p�ee�\�m�1�EӚ�{e,^.0O��-ߨ��*����,�h�!��'���ס�9�K��t����۱��VdD�6L�9p��x��M�ǝア�_�����ݭ���/e�=�N;���:E��r��'�G��d�ٜڕNG�534.�`�HRl����I�Pm�m�B $��\��OUusն	3��Y>͑��:'l��t�;C���?�u[��:��G��F?ނOc̴Я�V��Xg&�mO�泗5\�Z�}�O�,T�[�������Ҁ)�Rq�L�\�PrZ��`�11���}�`��)|�gn�^���z8��`�a�Զ�����h�����>1[=/��E�p3���U?|��ء���l�	��5.�/�P6���Kjf��K~7���R���g����>x�t=V8�H&j��Ϟ�n|Ԯ�]��H=�IO�4�*=�q}�0Әz�)� g$F�`(6�z���)�+�Ƞ!�ȱ%A��������U6'n�0	r�7��T5��뢖�/�o�j,�:K���>�^��.�-,ͮI�跺u�8��j�?��$�#|�[бD���ɰ۷A}��	�+�H�u��xR\Rm���0C�iL;V5�a5F�H�.F���7�C c�����=k� �l]�`$����v0g7O���xX5J=Qk�]��vo(����|.�E9�6�D�x�"��Y^
0��i��\ҿų��nELkv
�1<5��>�<� ��� �,`7^���r�,��M�:I��$�4q񁰄�5�U�Ⱥ�%�,\A�:e���ҝ�ǜ��������I�>����X�J�E������N�W�YkK1���3�x����������X�e@%�D䶲��/���}Έ=��r9���̈́G:�D:߭���r�(��~����-���o:�E��eb�Lu��X>�]�ߵ��هbM@��VB��SSŤ3a�c~"�4S�OJ�9E�&H@+�	�N�O�ja:�a�)3�++��~;�x�<��C�����[� 2dDؾFH�����;Y�d��[�W�L�5�m�V9�cH}��m)p�ڲ�@9t�ɢ6�܃힀��ڜǶ��U�v��[pO,ǢV-�.5ִJcS�8�,/�(﫵H�,�WA'��uMk�`"��\���<���ʎyo�m3�Vz�J����ɷ�&������|+K����N��2V �;�~{h����mW��5QWF��Z��(����R-����}IUS�[[ư�=�ՅX]B��Ρ�W
o��=��}�B�-iO�UN��kW`x��M��
"�@of#I��3��\ dl"���NWe�S\)ȩ�q�蕁w1��=�6�d.'^	�i��N�ߧ���I�i�1�$vvM��"O�'K�S֨��˾�'w��vTмv��"N���;̎ҐP�]��{�!d�.��&�=�=RT����	xrm��S�
����ͪ!{�����o���Ķ@���r]����E��#\�����wd���j��i��lOP&Კ+,�Z����U q�k#^,W=�&!�&[�����5��X���P��^�P2IUhQ �Q��k8��S����P������0,Aox��&��&W�oED�yj�������m�~�Vmy���]�j�(Ǥ@�d��������s;�V!�;/�Bhr�\�%�c�x�Q*צ��3�(EL�Eq��jnV}�a��n�N�_CZ�X�BϽ¡L�
�o�w}��B�3!O^�N��=W�)��ป
L>o�+ C�˻ƺd߭�@�z��08B@	��
�M�kG6��,'u�؃E��[�{j �����ZL���4�6W=AE�H��g/`��W��1,t���p�?���{���\y�]*�L�X���:�Y"��_�����"�bc%]�F�"�~�/du4.P�87��-����
@�Ok���0������D�i�eP��7v`�<@̔��z��z��9�ӷ�Dg)6�R���D0�왮���W�t`.؍V�:A㹿.b\�|�#��p�f��q����z���������P'L�|��p��='�
�tx��O��+�{���G"̊��齖^R��3c����>�X�k�;�D�'��� I��R��}�SQ&d&��Y� ��L��,@��߼�ֵc���0KL)y��(:^�P�>�Q�r>]��kG�
[�g-&y��eѣKy$����S]��T��CNl��S���7t%`6����S���kb
�B�d�r--���nmr�`47S��z����Q��<��$��� -`�N�hS���l����H�gpg�q��ߗ̋�YkkA��5y������N�Y�P���@b�9x��Xܗ�޾�K�����Y�n��`�Uہ�(��&H������2%x&��˼�`Hn��S"Kv����>c6�M��i�w��/�@*�O�������Mx�h��3��WZ	�����"-N���M�ZZi�gʯ�f}}*oeSP��c"�2�t�04a>���|��#�5��o��o��
j�v�4�Zг��Ea��
�;Y��F3��eP��|e��@7��J�$�i�'�,S��M���u�$�u9q�X.��Io�j�.���,]����ľ�$��m5�hS��[���?�>4���(5Jw�Oӛ&���,=k��ؘ)������T�`��ۇ�\ͮX�Հ%��a�+����;	��ҧ02�=r���Z�:����0��޷nr�>N�~����[��0�:��]���L�ߴ�9�Ɣ�rq��%���Y،���ٸ� :�a���"�fc�����4~c�)y?0u/���TXi�E ���ee��K�;m�W�O /-)�(Jz�F�)~��h��h��Zr*���vE�ѥ�v^�GU�&�>9I�Ccu��BM���탄]s{�T�Xǌʷ�>5(=#���P@.�o�ʭ��F=9��\�;.������ҩe2I��a���ϰ��"�*���D)�x���)ee0�*��7(6C:�?�;�o"���W�4I画Ϭ~L�l*m�i�?R�D��ԑ�3�9d�o�t�YL)���UL��o�����D�R��V4�^��#j�Z��3�����(�@�=��b��ʌ| aL�c5v��Xhx�kE�|���͇(�d�r ���%�v��yY�:~�Z�k�;BC:͢"����j�Mz��g�p���Y(N��Z,|:��^�ln\������#��9����5�c���4�*8:����a�B/�X�03�YJ�F��%�xY��^o��<�K�ƾ�S��?��F�[yE\�Q���9��q ��h?U��h8�]	(�[B���숭�ll�w5M�0v�Kh��ٍ���-Y��E�=ԣ�:d5P�Y5���������s��G^�'C���3#s�g����=T=�^����a8�o�9���YO���X��Cg������Gv������鰳�.ц�R��:F�R.�čUv_~�[Q���طk�O�X��?q\�:���H$���Ԭ���#޸�w��~�����be��w�*����]�m�yb$^�oI�n ?5wIE��ZK$*�-ُ;E�<	�ۖHބ��}�@6wn$|@ޞɫ�@�6�Q'.��O[����)��D��,�����?���Q��%�S�#" V����+�8e,�ޢ@���u�����87�� !+5�ܰ�l}ｵ<EP�(#F��8�Y?]7�"�~F)��~���'ssL/�QD�^��ד�j�t�<�Jܫ`��/�ΊS��A��~�+C� �>��^��W���V1�1���pۨ�����)D���OY�Dx��z��
6)A�2v<�g��Fs=r+�H�X ��w��h��[WAR8K����)M����
m�i����A�9���pN:2�BJ��s�^�� ��mU�2P?(�>��aG��tȤ��V�Q_9a�����H[cT��u��JG�f�LZ���f��X�!���u��TK�����3�����*McO	!޲^f�k-��rҰ7�[���y���(�o����̻��8��z��) ���0�g�DM���o7�����t��4-�͚�s5��YbRmhC�t~��{x� Q����P���ٯzE�0�Q}b2�RǁB�t��K�����2��9��W�P���Ť@�R�����J`du��gMaݴ�N�v-�'t�L�w{D��K�w�[�=^��˛c�m�d��a*1��o�|(�G�G�xp��P�wcFo���L�.~�tkO=L~�+p����H�H�ua�#�ʵ���Q�=�����{g�����>{�1u��}��/:?0��L�{��=$�z�E�,C�5��DSi���)8����P5$*�
�q!_�v	�C�~�E�5�LS6�<��\�"B[�����̺h~-��c�9�H�H�����X�y/���7]P4��%��Üץz[��'������Pj!)ɴ2�2��������&�j�a�w���v�&e�)�  ��293Зb��D
t� k��Z���Y:ߦ��#{љ��:�Y��	�D�A�1v���F���,�|ԠG���Y�Wg�l�J+\�ex	N#�`n)m���d[HZ����Ԯ�?�ā
�:cЯu����b�����-^*m���D��b��o��)n��w�0��D;*�WϏ=��<K���3��o��B��w��|�9��m���z�Qi�kv��Q�q)�I���-���W��a?���Q�g}�ս"#�@��O�+�o�,��@�dP���'�� �<�8�=��Z�+w��_�x}�oR<G:j��F�318O�]9�����)@}���K3su�=�s�����UE��v��ߌyK`Ò��O���7��
�C;7���D0�=Aߙh����1Qp�8���zQz�0�쨷ڑ�	*~Wi1]�h�F��7���4�����I<�#��
��v��!�lWJF��+$��XG�w�h� �^A�;���.@P�Ll�O�am:q�O砠^H��5�
2J�&���|�A��e��m:�2���?M�>[<7G���ȩ
����'_~��C�Ͳ.T�2�uk�IG�K�L_'���9?؝B�!������ZTp���}MH�#�k�������|!��Ef*-�����r����� ��u��;�����|����`�N�����U[�)��>]p��֒��q�N�hO�[�ȅ�rJg.YW�!EV�+__�����{'�!w�N$�m��A	l�O��E��_�QdBz�g����9}�k���l�pX��^�M��s���*%'f'�9D��~�P.������?��}]�.�8�
nFػU���� w;��=}fI��ne�I$�Z$�ׅ.V+I 5�E�Բ�R=z��[L���𭙲�ǿ���������Hp�z�@��:���T+�3gԔ�#�Ħ�i��̥����X�̡J$b�����yy���f��E�)~.f��vS�����0�s�w��=AD{7��|	��.R���r@Y��_�K����)�-�{ ]� 3^���J�.}U;Ij��ͻ���`�H	x�X?ycD���~ì5fU^bX,]'��&�L�/�M�~%��mLG-7��1C֓�}<�^z]N��/3�4��h�~VB���	�w8�k�O<��s�Ȇ��@���"g��!�& ^	�MN}���C�ZJ�M������W����{�B"�f�0ǡ���W��W_��uh��&5j����8�0d*�*G𣣓%u �#@����Jq^,+}���;0�������QԎ�bԗ'�6��J������T\�+��H3���y�����l6W�a6鱧�(UrSq5�2Ʀ����\I](�6bZ?{��,�_��Nq��R�E��CX�����K��%L����)�~V�e�/���X����%+K�?�����U�S\o<%�Ȕf=86X�(}q�7����I ��Dcѓ�(%������)�L���^����u��t��V8�,>	c+ئ�X-�`���ٴ�QUv3�e�R��O���a-{����}���f�Rmǧ ٹRL�ϫWv*�k��S1��oZf\��K��Gxш�fwM�t��a�5,��j�8�&����7�H�k8ο@C�����-'�RF3��vp���t�m��F�sR��_��^s��g�d�I�
���,���}(tr^����g/5�l8|�hb�!X�%L�Y���NA�P���h�?�L��Q]�~�݀A����8:�y�©tc���L-�����j/��Qk��;ܯ�艁��#��K�7o���|:}#��f�L��}C$�O*�N�իm!V*�#���j�u�fr�DK�w�xg�c��7L��U�a�cܳ�S�8�!Ǆ���g�Z<�����P���<R�Q���a�����CRߍ��Rq��_�K^I�$g�A���E��+|3�,h�l���{t�K˕y=gſlu|�~�����Av�!��tZs$�;�����Q�i��ms/��A�wE�p��ݡL��V�n�U[�.��� ���x(�bg�	\\���em���,F���Fu�6{�((SM0U������Q%�cd,0�	0a�K��~7�]��QPno߂Q��焻�}RI3�v�ܗo��u���N%��+,�!��`����sh�j��B�Q�ȁ���n�C�M��65�<���ܩ���A{�����S��,�넟Rr6���/�H�P0gA7���E�1�W>���4Q����K���!]��2�jV��ך��R"��d�	�t�t���1T]��"�9�/���.�p7c�^��	;�\��O�޶��X��Y�D�,e�8�7H�~<R�P��"-�VG�=��VD��N��^��an��q��ؔ�78 �jV̴�sb�����艞lr�9���"�+2����q�ⶭ�N
�p/��=y������!�=)C�����#E�Xů��DR�3�fŴ�Q�PL�������h
��- [C�R�%��=\d� �kd�ȼ;%^��TN��G�Xk 0ݪ�y�,�:p!���ƌQ��>/Ѣ}�r\a�g���yŘ�H1w# �5<�3Sx�04e�N�$�Y�� ���__+�@}����u3�Z��"�����D���ԍ�N8�^@[�^eƋ/��*�1/]B�P)d{F��/0S������ދmc�BE�h�J�������g�:R#K�m��RG<:��m��޴��>��-���V�^�+�R�����Z���Y�"̵:3̙����ZB\�g�
�f|<YoD�V�="l���4�4��,�|�#�4�o�t`��I& �UeIV3�
��|\�!�zr/���v��֏�7m=�I-bȎ��g�3��g"#��E$�`�֣���!b�����7N0�T��\P^#�S���uh�^4�<����>�3Z0��U�G���!p�|����k�mk�	��L���@#H��_��~�X��|�7�;�+����%;�N�A��a��ך�����)p8;h�����r܉-�<
�*JvАUUE}>+��u�}�B6_��[>�v���xD�����|��>'i(#�-P�s�ob�U���9A+b��
���,��ԉ��C:e��X�R}��S��ܬ*+���7X�]5�CZ�e�@*Ǳ;7x6u�?W���!î�r��W����*���V�L�L�m�G,?ľ�DO�𑓤��k !���&��L\{�<���󌽃D��6����^��%��I�j]H�&*��Sw�?��r-����|� S�ߡ�I��b�xļ�E�{e�Ŋ������ �%����e����(Z�<;t2���ߒ�Wן?t�����
}( �&Z'��_l��5T�[����	�E�]|!�eI�&.<8l�7�.�B��"�iY|R�Fc��%2����Fo�.����pOfS�c����8[�y%\9�~��B� �̓?bsh*ɵ	ZKw[�-��BA
���l�c�5� �v�u�h������1�-�-YS�a���l��5����%%��.^*JE�N���9��'u���uFzs��8�B,=��gۆL�Za*uu�����ct�;,����T��PM�v���..��"k.�,��D�:B ���N��?�vQ��[�JшJ����N�q��q�Н�uY�H1������޼5��~��j�;��~��ܷ�b��C�)�4*�4�%%���@�bֹ�o�en2O~w�[�0�*Ũc�m�<{��H6���%Хr6�w�{�|�T�ɝH�!�Q����3��;�)���E����^��?���Q�$_�q��N�+�ܕhs=��'�OXF9a�7(�a��R����Z*#o��Ԥ�	�8�#-�ѿ�B����j�Y?�F�F�%����Wo�P�`r��sSH�Ҹ��[k�\�)�a؅�A9 ��'?
��h��v	7X[ב���)խ݈@l�x�5b��v��,hP������P�SY�dB��%e�W>5e����-JR��oQM�U��z�LK'�,���s��[=IV��D��a�����N�{�������C�w�!�Ӂ�v���q�^���[.��һ�a�:k8�����v4{[�>��=�������qQ.jØo�H��A��?�!D�����m��Bc���(Jb�bU���w*��@h?[����b�p�oa��n��[w�W����?*�9a��ˀ<h`�K@�p!�5�Ww�||u�ɀ�- b_Q<�!�,c��8�)x�s�'��a�*��	`?:�iQ�`ɖ��#wn����+1�\,9=��w[+�v'��<:o��8�����H+���g}��<�j�=�F�L*8�[�],5���)��%���s�' 4�_���g��i9A�ߌ>`�����T��㤓�CnVf�qJ�����C�Y�1d�PpP�ܹ�"Iz��u�;�[���~�]`��F��P�r�l��U2��nu��t�
�ߍ�� ��(F+p+��kX�4�wI����S�A
'_�ko��W�_,�rmRK�����ٙ�(u�2�@B��( �d���CPm6�2�T?�4>NC,GQӊ�\���]�_�[Py "� ��TQ��u^1GFԵL�h��"F�N�!g6`�-`oT݆�p�Z��N|�� |��@��"!�t�f]dL�e�r�������ug�NTt�';��uƤߓi�K����h��|��~�Mkh|;J�׷>�q}-��s�������xb
	hC9�q�z�͚��GS�����2��0k��b��.�9�t�Z�������ݚ ����j!{�@A�$����JuR�:��a��VN�l�-��Z���w3���\��/Q[���ږ"�c��id<n��~�'�L(���GN�pR�����c��R��ѥ��1&t#Cb=�̀~W�p`�*�q� $Hafx��m��	v�=X��c֭�.g�}�����5��/���ܓ>�{u��$`��EGcCIC�o	<i�]����d�Q
زr��$�VC�)�����>���~�-�߻?Q�P��6r�2��SB�>˶	��r��~�c�|F� 6ܯx����?�y�����P�d��(��{��2-/�i0ؿ������j�9�l��2A�J�ƥ�0�j]��wfav�u�EO� ؔ�2����D�K�W�]����c���<��E8��Qg�%�Yo
�=������1.��P�P��:��4��G��YV	�$��+���2�30��4<��X6��x^��S1��@�����v3Qpz�z���-�DDgUv�N��@��ez���"\1�S��h�{���c�����Ք�?M��v%h6�КE��E:�n"IK�D��. "�bj�8�싖!9e�xr/���C��w ��ޙ�ӫ�Qn�e��N0�ǯ3���<G$����@\ћJʜ/�N<��3��Q`K�U�|��I �v�"h| y����|ҚuMH˶ޮ<���ͦ��:��O��#�8Ú���u��:�p�GE��FT�kO�����0)g��G�b�l��\>�+}�_�O�ԾTBđ��r��b�)�V�!�r\xn�������͆����%-)�[�n�.��b0�z(�s\��Gն��������|����l���cCdQۈ��=U4^�%� �DA!�~��5C-Ǣ�r QHj[�(K�cD�-P���~��6�����)��8CJ0j�	e�3��|	���$Ľ[z�X0η����ha�	ܴ@H�$͑g�GR<�L���iۤ�V�fz5�=w(�=�b�����P�c���d�k<�Ql��S6���0VƅO�e�x<�k��ūǽ�J�|={bE(	��k���W������թ*$��T�A�
-&��t�����&p����bN����/��A*��u���2�*����k����z���]=�)?����(�8��N��A�1�g,gm��,����2P6�^(��fMu?�z��8�V�v�c)F��n�V�P-����Ƣ���6�P���v���Iʉ��9�3�J&�<�������37�԰zf!'���DQ���o;n%��4�j�+�#�k�YQ�b�R��	��n��H�*Ħ�Hc����I-Qґ�����b�QO������s��JJ��
�����m�B}��f�����3����Q�<*�I�͚R�fQ�fV��K&�xK�@� ���n��a)���n׿8H"�����q���/��y�}��/Z�g��R�yo�0���r;������!R�`K_ۡ}^���g�t���4��$�,L���7�)tlr4���g�/Zlف��b�n�$�AZλ��=t>>(c(o���-�έ
j/J��A��V���*�O�I����\}���9G�v�C� {�*
U(�u��m�c@p �F�mv��,��*#)6l�U(
>M����y�儂5��c�����ۺ�D�ٍ��;�5�nPҏL�5
��B�aHY3�(��{n��ٚI�2m�ԏp�!�B`��W�j/��5g�����n�/!MT �613�"����L�f;e{����w���Ǆ߿6�6�7e�Hv2Yg�U���0v1"�D�����{ձĶ�R/]�?��Θ���)�0�"����m�v�Xg'�X�]��"���/��r.FMA7GA�m�@�8Oa�H���,�jD���eF�W7,�<�Ζ���6�p�ů�ID�%
�H6G��%��b���$��j �7Vi�$��~bR����Tq��L��PcY�g*~���	Ϗ(���`�F���2Ip�9d=]���j�Y�&f�C3��.�=g��<u�3�R�=3YXAŘڗ������Ö:Й���� ��R�`�I�Xd��5�vd��v��"� ��LB�L<��<��0AH�y�v:ԧ��t<Q��>mr��5@��g#��y��B�۸�K�����$^S��T`��m�{a{7�"Q`l�K���STc��*ӥx��d�0J-�ufn�=`j���CI�E�7Qjީ��ѻ��l>-}7��|�?�������'��d.��w&����A$mkဇJ�M5o�o.I�����8�Z�rB��]E�w��	�S&IOƳ�^V2f��g�o�A	pn���S�*��:3�?d�n�i*�]���@@�hTo��̶��)� �Q�T�����Zja��c"���u�'�.�OZLAg��0f�$�o��?�v�D"n�5I_4B���2W|��v��oc�tԣ���D ��mI���
�.A|^~�!1������8�!֑�77��=I�� ���)iT+��#��X$�Gt֥�(�c7�6T�z��0�ĉў��#�KN��uj��4���@�>CM�0�l�UMb9�S�+!2���=pk�P�����Oj�BWz�;ח�sXuj�90��m�
��H#;�-�C�u���"ܺ!o)rhB���}r��;�4؉E"�vR��U�)>-�1���p�ħ��]�(�x��^�
�>U�>)th#TVoP4G o$���lU9�g�ϣx��������e&��7������;�*�Ĕ��.��,�Ӆ	�eY��*�9�7
��6���?كD��[��tO�W�6=$УC�JL�pm?�?F��D/���7�Э����#�諫L�L�� ��c@��E!�8p�0ԍJ�s^�W���owj[C����d�\��"���m�����>�� U�l��Q
���x��xE��Z@'�{-��9 ��!%V�W�v��gZ�W5;���͖�)�s�]�A@ٞ�w���0(�UZ "�.�]lb���Ҵ3�K�P�߲���k��(�8��􁰂[B�5Դ$a�Y��JF�`m%�Q���Oo�N�?�W�2�DS�՛�7g�[mt�\�^����� 9�?�=�h,�	�r[6���.��7l���5A�VvJ�8h�ӂ������PY8���`9�V�m5D�T��D��\pvR�jw�m�;6<'�Z�����sX���<�=�-��]
xNa,��z��-�R��Ʒ���"hW�֒
���v�*�p�.��5.E2�F�r:��<�F�����vSr�[���x���f�se�q�p����H�_��� ���v���,�� �zkbY���C3*��qg8��a��b���o �nt3�w=���,�*�=)��SI<��9�
�턡k|��<wbJ�|��&ɟ���x�Q��h���cd)�0�8v������k?9HhQzƜ���-#r��@�v+��,x&�ޖl1�u\W��	.�8+#��t��+)�Q��}㝨<�.2,NF8��]����r&)2_���%s�^�����m�ׇN9�����>��`�ۈ������¤r��C-���`�f�Kj��~�1�~pO#�x��zrz�����;ݪ~	��]���F���q����U���j>�U��
mǄ�I��^�wFJD�+�*xX��Cw�-�R��A�	��EX \Y�~K���!m1)-�A�ڠ��[ŧz�2������5�Z����m�
2}=S?�>�WG�wț�q�-��_�X����hT�Au�T�G�g�LQ����	��!Fa����T�;'���JѮ����׮�!u f:���r	�q�r@����w�m���&$��T���R�>�~�����Q��^��M�\':ն/wt�eiA-�f��
��b)��C8���Y�󚗴e��m�!����	<0���b	%��8#!t����?����nث�GC���@@����h�J����Oa`(N���-�|��@�w2�������� [$EJ��c��d{��|�&��(b4yG�p�\�Xrc]�����@$t""=��:~2�p�박���_fa���ʌh%���=7/a"s��3�)��0�(�V�T"_/��;�r.{{4�V$�E�:��
���?i�x���f"�0iE�1��$��M[V�d�BZ?9Tg�׏�飴�.$�����x=WS ��3�'-|�ZYC?}p���W ���Q�Y�ޢ��5*0;Oi��\Y�����+�(g��ZÎݴ�_J�(��rL���r��?�J��^W���Vr�m_���� �ܔ�wa�$�_���1�l�s�M�_�g�d4�H��%��K9r����=l4#Ŝ~��[݈����ߤ'�8I99Ǜ~c/�t�v8~�m�z���J�_nذ���1a ������9�	Ǆe���$v��].�o, j��E�Κ�5˺R�z���[�-���X������M}�Vݜ�i�H���zG`��9��ѳ�+i#��uY�拐���̺�up�XٸO�?�b������yyu�fK0E��.�u�c�2��Ȳ��Cs��R�%{���|nY.���& @N+�_|i��C�I)��{�� H>�ͣ-~����U0�Ɩ����*f��#/�fyxi��¾����US���u'@1�&�-�/K	J�����"�0G�zH�&��k�Q<^e]#~/��t4�K�3�S�	�F	}J�� ��<3N��q�ε���w��0�{m;	��N�s_��Z��E�Q�䐓��$1�����^m�jS?�|z�������]u�~u��g�"t7Ϋ3Lk��/�^��Ci�yp�+�~ڸnd Y(O�L��0�q8����,F��1����*�D ��ޅ�Jh�E?�6N���q�R$J�W˦tV�T_b@��7JƠ�w�I$V2À��lԃ��D[�_�:�d��D�ة�B�Z9�{��ET^lTT�4��,���2�x��m'��%9�	~��#���ZY��ZrϽ��4���+�����; �|��<l��j"��%he�3$5'	�4.�� T� E�9����n�z�t2[�h��O��P��°���{��s�H/K|z1(1�c�N�;�+�Գ"��֙�H �dU�Z(X桩.}b�`+����y�Ifn�E��.ʏ�~�XǍ�o?s�#��<qA{�E|��.�N��@��J_&?�-J�)��{��� �؏͍Q����U�?�Ǐň����GW��f,y"/����+k�U�G�k��'*P�&�)B/��]�=>�}*G�{r����� <��]MT/ 4[�����3NL	�:�ʪ�;<��ǁ���4��F��/����	~NNB{D��	�ZIQ㯪J�]�����{�Ȩ�]������4mz��p���	h�+B5	�M��[|�����i����l$���Ḽ�Jz(+�@���n���<�%����}�����JX?ϯd��\V�f������}���'�K�C�����P!�(�(q�@2�R��'�I\}Q6AOG���˫^_.�<q?���~�Cwu����K�7HLŋW��{t�I�C�K/�5X������Kr�о�ѝ���\��8%��,f|��X"�t}p����PI���=�<�%��F��J�H��͌���L���B���N�ċF�cj���-����)��\Q�	����ٱ�-��2��d�`�ܞҎ>}�=�fW$�&��9�7�}�v�*��ѳ2ݴk)�f��vKk�Hx0^,���-��3�?)��\&\B�x2Ȭ���u�#���N��Z͗�:������G㋕�u!��:SߥG�'FEǛO)���5�M	v8g,�?@��v\!}ݟ�O��Ts���9yt��ty)�5~��CM\I5!x;@���ͷ�=����f�O)B;vn� 6�38�z�������=ʛ�V
ȩ\�H����k����uo��IU��G�l�ݓ%��4�OJ554�֢>{Q�Xj��IK��ݾ2���积�k��A�:�88toVj�OϤ�B|��cPWKĎg��I�!������'�	-A&H4;d����R�#İ�i̋�V�+�5�v��u������xz֌��c� ��U�kM֕l��X��+a0笰O3<x�
���_k&����T�0|�4�E���d[xnt�@_Z
�mli�o�?!E���E��Q
XW��h�Sz��"�ҏ�]7�P䏈���n�,~siM&@�	��$0�Cq�}�����sߺwK�,�1�ѐ�)��'�D���|��f[�\?�>��3�B�jJK6ӆ���C_��׾�k������������u��^��GE�XEKW%L��6�W�N%-�,���#K� �r�>n�M�:CZ����Ih~r��C,Ń~"?r��I�Aܡ:{���L��w����䜵r�A����6���ci�Ej"a#�E"rZ	��`9�v\&�u�3V�Ώ�O��a�/���~m3r����;0.�<Q��z���۷I ��FX�H��j�b��;�ȥ�AW�ׇ�?U�7eEk�{*E�6������ɡ}Y�Pf��B�3%���Bu���c/�*?�v�_+�8G�fh��Kx�x�����4���?a{�G� �c8���3U��q�w�w�K�s�ފ�C"RR�0�������5��Rl�R�S�_��&^��zg&���(J���2m
,�9�	J[t~���/>�g;{Ll�?Թt["�q��A�-WM�tPob��� 凝�οt�/�i�A;E�����3�����I��O���K����i��:�7��Ħ(؊UɿB�#��}m���,����=6>R�(�M�F����j3�G�vc]�+��;���������1�P��ĂG3��:����Fm3���܍Y��+���d��aZ�!�̓`b@���r�j-��GD)�F*Jnr�UM&�~6+G(�t�9� /��8pT{����g(2��[M��,6�>R�o�H��gw<퐟�j1t�уH-����þi��k]r۞�1D������ө"5j��?�m�jS�˪�]J�"��W/�j.���7�M���e��R��O� �x]�����D'�e�eH7���<�䊉뛭����W̊���D�����|�S;ߵ4z<����$�v3�V;���\b��S�kܙ���ݞb�`��E�o�a;����֙����pee=o8N���ŗ��s`�썌�������cR�ճ3��6�*�@��Q��X7��C��Z�v ��ZRΌڷ��$dn{��T�����tV��'���~ �Nh�0�F9y4?8:��H��N�Q_|>�.��חR�hguۏy;����E�K�!6�P.pS�LT2P����Yݿ�7�a-`~��-�S��س�v���dE�"--�Qn�v�`|�F������Q<�Ⱥ��3G-�Y�s�*<���Lz㈯ [������8��&k��q\��5�Z�*8%�5Y"Ҵ�����k8��8N��@���Q�fK��T#ndK7�@�e)��&yX�ץ
���q����WF�����Rq,����QܔX��I�s~�!����"h�赒I�UF���8`�A-F3E�qpa��e�#�"���<��z��ٮ4B��?#PfF�m�>z'��r]P�)�я��*�mB��T�0�T��*�1����F,�y��R���w����� �iW��*'���%S�A�j.��r,�C���W�H�iN݈��;P����,gC��"D������۾(��f�'�P��`�`yC����b��xT�� ��^9P���uXK�����G���|_*��>�������c��!�F-%�,���g�Q�T��s�a� �o�3jܱo,V����}[͓f��3���8>��xc��2��%�"S\��}�HGO��[Tk�ϡ1�����)�9����!\A�p\A��3ͯ�
���@^�h):��n����+��z�g|T3�@���ә���ȡP(�@9�������>mBE���U}�i�9݋���.G�5,zȢ�I|�j�+�K��ݶ/��J
�����ȷ2˟8l��j��Ϝ��|���H2}Ć���A/6���'���	%�H,p|���R�v�Ĩʶi�|�V�;^5����c��87���Iք�zc{J��Mn�kE^�lՃ��u�#�10�p(O+a�xЬ£�k����S7�(��|��\E�,͆�{xf�
�8�T
��iod�7wȳ��EĔ
P�M����$�����u�҇��7��]䇴߃�L,v}�M�]$:$(wq�L���<����on�,���ш�<�����<�_�:'�^��T[>�"��:��J����~)=�;����lk�����G�����w�Z�V3��?�X=-%D���.eݭF1`���n��q�)�r����E1�:;�y�䱭A�rz�O$'~����	�9�f:sye��L��s��xb�վ��j����:��.���[�=?<aM�"jM��q�9��&�%�+�����O�3�a�4���3jKs��R;(Vz<x��r���|� �=4P�1H��@�Z&d;�h��ߙ���L'��L?�V��+H���m�n��*iJ9�b��揃e�/�c�����������6pǠ��0������S�"��W'@�#sn��45A��U����ԳF�~�H�a�U��$�m���V�����/�\,��	���)��A�p�Xi�V��;T�h7*]��Ex�WQ�C��-�(*E��ߴ��6}����+��dE��&�B-̡��
�J����}���B�[Oc�N3�2W�a��%�
�Uo�e~H�q�d��S��W�l\�e��R=���#1dq�A�d��	v ���U��W�Z����(�&1E�%v���ⶂ���S�*Ѿ	�!�D�V�4���4˄X�����D�����]6IhDE���&fIKD��=��ժmrZ	��r�K�Sv%��YK	��+�*�S��&?�*�@4�GrՇl׆�����w#Ԣ�̓#W���C�����%�vJP�� ����Z����=�kq���^�W�=� '&�Yᇠ��ʔ�� ��k�`���s�d�t5Z&�.�t�8�/�WO��u(/!�s%����m$�Ox���M��Ύh~����N�r7��q��ڨ�5��<�M�H��Cb��'�׀�.�ڀgU?�����n��{4�:�U��d'�$.,��y	�������³S?4EAU�����%�t�D�����r9�:�F���ӇR�n�-W�˙��`J�su�.��ӿ�l��L.މ�T��veb`Uq�-]�[�h�I��U\��j��R=�Dzp���-Bܦ�#G� �D?hzބh�	G?������3a�B��<�'��TxP~��3��B�Z�x���"����I��J Mi.S*������AS?6.P�c'���9W��i%*��˲;�lҺ4ޕC�'D҈)�3�۵�A͚?'�ȨP�	�� ��C80 �C���C�T�z���z^���P��Bu�
����A��@��W��b���� Te��}gx�F�'�H �V�};�[��B��%e��"b	��.I����ﾽ��K�x���i��'���x�u�)�^[��������X�*���H"�ثP`ƬHǚ^w'Cfs�p�Q�>��KZ�Y� '�i�20�v|�CqѼ)nu��Y���,�!���[d�J3������Y��F����J��W���V`6_���M�#W`w��c$�Ϝý��l� ���_��d�Aʱc���?�a9y�s��6�l�}�l���Ia����&P�'�v9@ex�-�8$+)�h�¾�[�A�)���N��8Hɤ�#hmk�B��K��J:8š�726��bV���H���Åm&�i2���?9�u>��G�6��qk��
_�Ğ��=�9odT�|�u�n�G��L�9J���W�	��!�Ǫ�fT\������kŇ)Z���u�-!�f�A� rǩ��͸�.�ڮ']b� _���i8��o��������ya����MD:n4W���c��>�ʓ�-j_�/�����b�C2}�Փ���JZ���i����d�0$[�b�6S�2l�t��<
���w������	^�5T#ꔴ��7��ZqZ;s�,��|ݟjoF�$1���{�(KW~Zɷt��lK�K1@�;{Ք?��H�g�`/U��A�8wP_���B���M�VYi'FN��%}��]�No�l'�(�@�;�HSP+Ҁ&[�F\�)��M�{ h��?ҏuhU��	��[��j��\���l�}>5*\�vS>xh���K��UY��k¤�����5-fb�ֈ��^��@��=L��g�'�����Csa��o=�ZRj���a�jn�癱������"���kDh�?�6��ԋvH���9�v鍲x.Na��o�9:ͳ�ïSrĊ&�v�n�[��;��Cw�̎�М�]q��`;H|��a1���ɝ_<��5%��
C��g�b�T��t��*Hu0< �J9Sb���o)��n��aw��v�W#Q*p��x�<�E��׀���q��5�w�l�|=c��H�@���Q�Hqo���{)@c����)�ޣe?w�Qc�}���/#?����+���,� �?�<�>D��r�C788T�ٽ�5+�8�ڧQ}��L<��[�F�18��|]���ۢ0)�Һ�[P�s��]�E@��]Aװ?3�1
ߧv`���k0@���>�[�C6�Q�9j[Z�ߴP�S��1,u�p�#�a�wz{a����ep~r<C](� Fo�
�:Uh��s���Ee�~$�
��Γ��u���6F�l=+_h�X��w�_�{K.A� �3�.�^Z �D�#P�J.���a�@Lv*.���!��3�6 �����zF���Ueڞ�$�N�lF�.�p	 �cE3���DT�#z�p[#h��㎲��c����؈(�+�H�lz�tj߻b����+kǕ��$�h��Ǡ=̼N��L�X[���ɣbF%�=��y��!fƪ$E��/.]� ��)��9u���s �t��{{n��| ��.I#+r�@>K_~�(���)8S{W�� JZ������U�a���Z�+歟z����yzg��}.ÃzUB��!'�@$&-%"/�<��h߃"��lb�W�#�������k�,S_}ѻ�!����/'�^�����gY!>j�D�w�J--��g�.xo�"��kv����륷�3��J�Ձ�_�����X0%�+��r�Y���q�R��"��ؚrD��8y�:��:8���TFr�� �^�~M��8��,&�:�be��
L Q�oE�2���}�m�^�!�)ٮ(�U�a.:`"��o���9�?m&Sd�ý�MLO:M�a�kӦL<93=�&�IHz;�w�<�����ӆ�� ��_���Hb�%�d�;dm9��v_�"{Lڳ_U&V$^�HșPm�/\ڽP�9�<(���<�B6�ڇ[�����!#f p���!�!Y�W�՞S�M��w2�Zޯ� �����A�M쀠����>�G�	�Q�o���f���m|:VE�����BG���$��F|��z�����KO�Vٯ�;[hJ/����=���Qm�e�I(nr�X��B0�}�^��F���7��0��B�f����
�4��h.}�rIB�#pO6�:NfWk*�ظ�
��o���v����d��_��dfWpl^\~W$��mu����1���!�Tdy	�|��%8��JL��`���81X�vati�&^��ؘ^��վ\Y����X�GG;��0��Q׬�����]�b��幱�&�E�x$=�׫� ��	|�r8+S)l��lhM����Z������\@'�r(�$�9)���v�#G%��f��"ޫ��S�ԩ��
JPQ8��h�Zl����zq-`�^7��=��(&���S9����Vޓ�*kk,C�>�sW|�t(d�&P`�X�Z8��yW��*�HbY!;�s��z�ɺ��d:�c[�M�?��F�f3�9i�ʶBqrd��һY�M����	k5o�?*V'^��-�Ә�?R��@L�4J4��fU/�J'3��,�+Ey\Ű�QE?���&+�4�!GSƸQ��7]B�g*d�;����WF6�J�Z�aR�����ܾ5D��d�s(X�����L���:"���q�	��`HP�-���J��Գ|�M��%l��M�z1N��%�B/�#�IN�W CzQh��ܘΆӈ���TV�B������T�t��[�
�L<+<��:P�u�B���CvP�*��X ��v2�/~�O}<D�M����Q���b���G!&�:�����'&*YDE����1����E�������OG�QY+���H+)1��*�3��(4�E��0˭(*��d5��W@�((�p�53���o����Dy��݋vNadP@�g�e/���w1؈���{/j
8'��<k��2������˘�h+Y��k���>l�CB�K_x�CiZ���`:����9�y�x�����h���߽��T��WDH���e�~kNŀ��Q����7T��ӓ��
nٛnVݜ$��N��3�H` ��ҝ�K.I� �w�, n���Y��_�u"|^�S]6��~-�[��:1�R��&�¼�Oy]ue8:�3GZmrF	�5Om�����M�Gg��>Y����\S��}�I1O��T7�<�}����`6)ϙ��0�\���<iU����{nU�0d�*G)��nNqO�w�z���Ȇ ���$�|��J��ȝ����B:�i��� ��t�U�6cZ�?�ו��m��N5��"�Z0>zj�8�K����C�a䰯񖓮�I|�~��88.XjXl��hT�|�`���� ��x����ʼ]j!	q�H�>&�<D�R�(U���%i���V�)55�=P.r����F�Pqc����πk��pl�G��H�lW0+1O�*�x���kj�N�#�t�$|r�2E�xa����x��1?
�w�i�J�̯҃�๱Em
l������  ���\���pQ7Q�w��;��,�$kM��M�$���qԹ�������;hc,����Tq�J�Z��.�W3��*�����o>�(cˆg�J�,�������r�z�k���ؒG�Q¯��2~�"�LӋcX	2�%��������������A���r�`9�U�:�Q+����rF��p�~欟��ok��:��F��WL9sD�ȮH�!�4�6�҇&-X��.V٧4�	��ag�H"6�a��9��&������_�OS��a�ߋ��7 3�RͲ�}�;t`s<���ӟ� ��!�H�j��&#;�h��?��_oL����V}�HA��mmw��v��9����˝�1�_{%���1}�W�����R��p�����rB���
SKm���<��7�o���p�KA�숀�^�$\~��=R��hš-�j�=�mU'�V>8{����{�i�=��U#fob���ւ�$�V� �; �h�§�V��b��Q�aУ(�����[�1}A���l���3��w�B`���W�
�w���2}�W�B믻O���N�hW$Bؑ�
�o�HmT�ܻ=��d0q���W)�u\W1,���x�٪�1R,��z�d��%	B����cV�#����^���91��v�ۍey�kzt��� �U@M���Ѐ�h� ��Z{�C��*q��َ]�204W���c&2?���5=��᪹$�	U�sr1��SBD<�C�e�v�ٶ�ˌ�eh�@ ґr!���R
�	{�#��M������R�?ĭ9*7Pj"���zZŰ�̉@�qƮ�^�S=b@?&�r��l,��1e��k��?��e�sGt�&I�Dq��8�W3W*���o!�hjsq�����:�]�U�|`{MH���4�x�߹���R+��[qKL��G��r�VM�VP �r�؜*'^T��}��̰#?k'��.;��ru�4�I�U���'�6,tq8yU��je�8^��-4��ٺ��qiC�l&�`��T��F�]���5.R��j�y��ܗҎ�7?sA�������������q���\`!��-�;��4���R�����|<m�z�Cٱ��B(�>#�����z��U4�l1,�8��-��B�%���?�T�d��ы��.ܽD]j��|ᔪx	�X�� �Kiz��*���n�A�L.c6�/נ�K�W���iqV׮���;3�Ж�e޴�"^�"��IEBr�|��y�z�`[��h���M�,�_����Hǰ�7H��<zN�� ����6�+�D�Pƶ�M��%���/�wRX�ug�T,b�1�Ԃ��y�M�fK0UEq."�h�JY������l��sea6�ybx{��Z|E3�.��Ѫ@3�_#j����j)���{ܡ� o:�ͪ���jX�U�����gӈp�k��"�v��y��2��V\���U�h!�'�t�&�g/�J:�����)�6Gi
��}K�1<�8)]��X/�Q�4�컁:����Ik	D��ʧ�<��N����ǭ��4�����b��	���N?ۄ2Z����������{׉Y�"�P��#����>����]�Fh�5&%��R�����f�u�_mZav���hu�5Y�J-�y+�ȶ��V����������� �9z*Ju8��!�D\�N������_P��6�F�(WI�>�l�m��(���q��2�l�a�+I���6w�K/���>�_�xeqp@��:COC�#K��YLBܟ�����G���|�/��XI�N�V�,KOT��;;-�ɚ\��i%R�wfy�{X�h}�݀긹bI<�/� ����O�%E�.��������
a�����'��0�9J�l��H�cg:����-S�l�ѽ/�Q����4j��-my^>�����}	o�ftv���K�uU�4aN���*�Dl�	˴�4f��K(�x��ꗢM��0(�a+�޳�g�8ʺ@m:�s\[�'����G��ie�i�
R,0����D�����1���RW�?_�}�^�eg����y`\!���,��˹r�t.��R�g�%kl[@ȹ$r��!��A�&Mt ^{����7N�o;�/L=A�F	�V�*��@�K�����B�����x���ꫛ����(��<�og����ȹ*m8H,���lй6�:�(��M�f���_|�+~���c��Z�/Q޺1Ԡ�Ā���m'�wL�PT8]���/��U��9�3|BM�=����K�t/��{!��I-��G@t���>�xPf}�b�"l`:J7���FY�|�����S����>8�
��d�gBזa���Y�`�F��'%(-�h��oLbu��"M�f��S����k��[!--\/.�4kl�.� 3,�?��9h��@	ЅZ[���8񥭰>*l,��5�4�v~0*hf���6�cN1YI��¯�ģ�1m5��>�v�\'�Ĉ`w�D�o��G�'�ԫ&�s��
V;=�o���]Ba�%<�R�6����`PW��V������FUvS$�פ[�X��.y?߻�T�:�ȭ��=�5"�v��[�=���#���g�'�5q��ë�H'�ld��Tƍ�*��`��Е�f�R�2b=J��*S=��Dd�Ob̎o��2n�9�w���*{���S�<��y�>�.�U�إ�6�w�|�J;�S�j3m:Q�9^��-�7[)+w�*!��\�ޮ�   �  v  �  �  �%  �.  K5  �;  �A  H  aN  �T  �Z  *a  ng  �m  �s  2z  t�  ��  ��  >�  ��  ğ  �  ͭ  �  ��  h�  ��  &�  ��  ��  @�  H�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ��|��B�,�r�Ռu3�h�C��'8!�D_��p-���K$��aU�/ �O@�	i�OOx�h��	:T�)�"��,n:�;�'�ś ֬y0<�Ɂ�މu\�	)�'C �8�:\[B��@�׵olV��
�'(��#t.\Q֕����c3��q�'�F|#�άt1�@+ 
�-W�Ɉ�'�|�Q��I�A��A�Q	5�d��'EXհ��IB�k�	K�PV�%I��hO�!�s+�'\�F���ز=����"O�Pr��� +�Q[2�[�_�� ��"Ov4�m�?Vd݆p:D�D"O�3��S�( ���1qZ��Q�>yG�'�j�AF�O��4���E�5�t��'Q��4hV�0i�tK��*��m:�'�K�N2��F!�9��hê�\����?�'%��)&Β�C´�;@�C%IK�a�ȓ`��s���8!m��Ks�%�t�Ў��s���Ū�1|_��z�%�"e:"���4D����Ƣ]!.�c׋X
[��Zu�����xbB�6����MT��
�� ؏�y2�*=2D�w���2��5�*��y�?@��2�r@@0�X6�y
� �E��U�x��\z��P+E<b�"O�0�䌆�n[�!�� �Tx��d&LO���h��Ԩx��E-�BG"O�D�������Mb��XL1�"O�	�F��;(�bhc�-��H \�"On%a��Y�l�{$���BS�"O�ఢ#̷F�0 �G+�VX�"O^���Æ�u�n���Ɉ: @�I�"Ot�!�'BR��F^�P:� ��"O�x�ь�(v(���{6���"OLH���Ti��a�dU*'�'�!���kP���^\��'� L�!��[5	�V����:GPƠ��e�Q�!��$
�
�"�Zi<`�G��.'�!�d)Bà4�cD����<!��� �!��1E)�)�ի�':昌�̘#o�!�dN�|4X�����W�M3��k�!�$��DX����-���VK��?�!���X���`# I���_#+�!�d�)%_�ʆ�f

*�P�2C!�$Yh�|\�`��� �Z����=!�ı�n�7F�0{�xu��M�<a:!��* �6Ҳ�]:�x4��!!k�!�DDL��y���Xl�Q��ͯYta}�>Q <hwR�X�%Ym|,[�NA�<��FT�(�� �J>v:Ț�LM~�<�"�N{\!J�#;5>&�$�Iw�<�GZ�F�Dzgჹ(�v!�t�p�<�Aj��e��,9��5}:�d��h�<y'l�]&
�1$�q�i9���c}
���hO��b��1^h@SV��>3��g�'�MP�0A2MB�Ni�����1KF���>��`���j���|6��s/�30�	��J�0H����+����glΕz�"̇ȓm�2\��L�x��\YwKő2OZ��<y���	 7��L���
u����a�k�!�$�g��e`	�9�i�� �n�➟����锅0�t�:c̊@����2���C3!�$�� �~��T+�6��uH7&��Q��/e���N��V�n5� ��)MZ�͇ȓ]�.��M�������@�IM�����z�E,f���9R��.9��s��)�}�Gԛ���$.3����C�y��	@lY��d%-V&Y����y"ݛVd&�������TPg���y���%mB�`��GS z%�uK@ȅ��y�葎�=��L��C#Ԣ�>�yB��l�|���i��?Ĺimޛ�ybo�o�d�Q���+:b|<�U���$�O��"}�E�VWB�ု�.��� ,@a�<�'jަF�7�ս}S֙j'.y���=��� d�ZP��n�9/�Vi*�SL�<1�鐡S�ʨ��E9��T2 ��|�<I�i^�%�>@ ��3o8��e(�w���?Y�W7U����)Ӳ!Z����z�<�G��U��j�L5NH��2T�,����N�����Z#�$[$�9D��s�ʑ8n�
-�Y-����/"�Iz���)�[x
@H���EA��d"D�x*螙HU���'^�Q�ƜR�o>D��[5H�q��iR��-��ibi/O"=Q6��\�y��bԺMw�հq�u�<		C\�z�WO�/��A�5��h��hO1�^0�"\>�T�'�
$��"O�  =�r��xN�1���>�1��IyX���q��<6�B}Cw�"tM��Q*:D�D"6�_m/t!�b�#��>D�����P
����uB7���O;\O<c��W�;t�ZMU���4��2�h9D��2��N*O��t��KԵhɶ	"��7�	]���'b�6y(6�mwJ����ߵ1�lX��*L=��ʂ�W�����k�1m ���6�\h�S���k�Q�%�)i�!�ȓ/����l�r����3��0cI���O',S����V/j���ɭ  �P�ȓG�H�FÙ�M�D�׀�2����>߰��,�TJ�I�w�[�v1D��<�����ӻ-����'�ۆ�>t��'Q�E�!���DfNd�W@�y��ђ�!�e_!�dR�^����;p� �@c�0P�!򄆗e(� 
Ãٱ>�TBGb�	]�!�;n� b.�6�I+u��G!�@<�Xce�1!�dU��	�R4!�DVD�R�#�B�E������~|!���9_�$}aFOڵL�pϋ�s\!��ܯRT4�&����$:���ML!��G�-,�e��j�і^=�t�s2!��$���Zv(M+6�*�l�Y�!�U�yF�X{�E�(:"��9Gl�|!��-r�<ate���(F�$�!�d�'J�L�W)J8l�*ؑ��I�!�d�G�X��M�L��I��)�8Bt!�	�z�;�^�
�� Wd�0s�'���%�=-+ΐ��-�w[���'�Nq�g��^|�EG�&q�"�
�'�����J(pUd��g؞d,���'4�ЃRD�#kĞ��t�U#V��<P�'�V�D�	<`����K��0��'WJ�`@LW��p ���s�;�G�<��+��@6ё�&�+�f����F�<ɰ�=N�"�B�	rH(E�UA�f�<!��6W\��f��6vz�Ѥcw�<Y)I/V�*�ȒH��^dPE��k�<����U��C1��ҤX��Ag�<A��?B�^�#�w���g�a�<q�Y�.�����1PO^(�R��[�<�Fd	xQR����O,�8%Hb
X�<�)G^��!�R�|�G`}�<)#�9�l�l��bi\H�v�^y�<q�K��s2$�0�j�5�@L�1�XQ�<Y]yG� '�ܶii��4h�j%!�D�
� ( ���6	�C�ªg�!�Ć#H�Y�2F�
�E0`�dJ!�DP�=���Z��8~���5P�!�D� �,��t�*�����m�!�+�|2��P��uصP��!�D�2��I�H<L�Z,pwL��p!�d�E|T��CL�J̓%�Ƣq1!�;4*�����[���`�G	�01!�d92�8��F�JH4�;��WW:!�3b���O_�73N�K�S�s�!�D̵i���ku�ǩS(n���8+!�d˽]Z�D[햻p��Q���T�!�$�i�<��mι �\a�-D�m�!򤆫	Ǆ�C�C�(��QE-�0Wi!�dªc�0�[�9�fh�t�=!�dK�]'�麀���}�J�*c��`X!�d�l�����b�⼻��@�2?!�� X,����� 	��+�h@��"O ���rZ`��G����	�"O�!��Nױ{��E+^9LC�0�"O�u%�SUE�{�ކ(/�� "O�4��j�WE�|3�ǅ�j<�]8��'�B�'l��'��'ZR�'�'�Zl��R'$�\P��'2U"h���'d��'pr�'B�'�B�'Cb�'u�d���ԾvR����E�tp4(#�'#��'-B�'���'j��'F��'/��2-��i�V�+���;[����'�R�'0��'���'���'Qb�'��LY���r��gW�"�ՐC�'��'���'��'t�'��'x!��JܒH�
�#���fl\ ��'���':2�'�'�r�'l2�'��u�W��>&adCϋ%D@=#��'�2�'�'~��'�'N2�'�ܰ��T� �x���6Qr�\���'���';r�'(b�'b�'xR�'��X�OɨZ��!��A8f��9�'�'�2�''B�'K��'l��'�dJq ` �9oQ/\��(��'��'���'��'vr�'VB�'u(�J�d�"�U�$����'���'���'(2�'Rb�'R�'�^H�F�#��sސ0�t�'B�'��'0��'��'��'q����,�ѲQ�T��7N1U�'���'�"�'Bb�'o��b�����O�hru�D�N2��R���!�� *�fy��'��)�3?!Կiڭ��M��FCp���`d�4�S��	��禹�	I�i>�	ٟ��)"H(,��E�N/kG2�J�ERџt�I0r��oZO~9�xU��Q�)ی\�~�S1+p�c Ù[}1Or��<��	�>0����U��-L,13f�=d|�n0Q��c����U��y��I I,DX��D�vp�$�[p,�?a���y2T�b>}�����͓^)
�iƢٻlR��U��"X�yϓ�y��O,���4�x�dT�� �#B�.�pA�d�[���$�<�M>y4�izv�яyB$u5n��W��!z��	���IE�O�@�'uR�'o�D�|�4!�?&w�Q�A�P�`�qW`/?���B������W̧B������?Q�b��-����� �DOv"�g�����<)�S��yb�^@�z�"�8N6�)�S 7�y"`~�<Dxe��l�ߴ�����j�?7��$)���@0MS�'�y��'o��'+ni��iJ�	�|���O��\��ׁ�hyZbY&~�Ԭ�aH/D�`�c���\�H s�l�t��);D���FnI�f�Xy��KAw�(sQd�o���&�<D�7��5Y��Y�o�w����IDc?ƈ3�f�s��d+��	ou6-��AH�`�R��@G_�\5�IQ�މnq�T�&��h��j�C-�MHWDM�t���EX�@�逤d�}�nX�!+еP��d�l�s=&�	Dlɪ �����	5x�iB� Vg��)ɞ"�C�I�:���� g�a�V���
�b�ɃK\-crePe��d풀� ���*��e�q�QK�`藭�X	H�*,�,)m+!d��Q�q�Z��ˉIx}f�H+�A *�,���*zj� i��yycT�
�`>����,3��%"�N�\�@�4&@US~�3�/Y�'K(� �/AןL���4�	4�u�'^2Ň"M~��30#��#u=S˞�C=�����O?:(��K���;C�"���O&�����Y̓�p�a1W$d���H���s�L'��BC�5��=���mB��֘~r`��>u��D�L�b���Gʮ'�� ��Uu����<SR�'(b�ħ|j��
�~b�� �,p��Yi��Vi�<!u�^,YX�:��'R�ʠ
�L�-����S֟|�'��t���l��``lD*�jɻg�0T�^����Or�d�Of�d�������O��e�h��C���<%�T���f�!�
C�dɢ�型|1]�"�'x�e��LH��	7��D>�mwĆy�2�0��D4�(0w�q(�8�t)��'�i�=��C�ӟx�	/�y[�Ƅ,d�T�cE�N�d1�Iw��h����(���X�+Y{n�EC��+V�!��#V���e'�j��x$"�a���W�����C�S�O2Xuz�\��ĀB��0j�p�'9&,��U��ճT�ø�JD��'/ 0��lW�#㐅�3��0pt��
�'�΄�T]!E�F�r[�S,�̃	�'_4��#Oǈ䶝��b��@X�	�'[�E���]=(�.�.ԄeQ#���y��ˎVA��aR#�=-�u���y�#F���c�M1#Դp#��;�yB)�Q�,��u���z�a�E�(�yb+V	��&�Ҝ^�t�Ō��y��@�ĥ���=P�\|���Τ�yb	_�ʥ���67Dh\B��.�y"g 7�� �ʞ+2}K����y���z�D&�83pڱa ���y
� 4�p)ߐ/��xR$��; rt(C"O`y��'7v����lɱB�j��2"O��A,O�x�K��7c�ذ�"O��F@@�X�a��$��ju�v"O�0�F4̞	��E�,��"O� b�/N�>�hbC�/,���f"Oh 9`�Ơ��ʒA�-,�j)ʓ"O�1RB,N?�h�2�!��%N\u�"O �I�'#�i����ي�"O>�i!F\�V@|�".�4P�"OV�F��8�l��/��G"O�tz�E�> �s�ēA%tDIV"O>!��HݹQ�����Ⱥ`ī�$"OHJRKRA�t`S&A�7u* <��"O�m�ċ�.�<�:�ʙ�t�%�"O�d�2h�+'����JN�0&�R�O��W�׋(��;6�V�V�
�K5�F�<�6��=%�1�E��4ӆ����NE�'���j�(�S-0��U�C��u����cX���B䉪C˞؈�۰+˜�������8\�\�>��<E�I޺Q����!\� ]�Ê�.�y�iT�H��h���َ���Fh��]F�p5O��j��^!-6��I?�4��)V�uۊ����˒=�`�Ӑ.!�O�hJ���1HP��# �tLX�p�#~/J)�`�%~��IÌ�jX��z�MV-2x32��!2@��`�(�o��H��U&/�F��5L(Y���
Z�"UA�a
Y��RB��"C\Lا�	`4�H3�F9�%1O&�QA�Z�a�����a��M�?qY�OQ4 'zyH�GK�P��0Sd3D��3jG�s��1���Y7��؇�s!v:3��J��t��=H8ʧ�OxD�"%�*���*Cc3w�c�'ni)��HҤh'oL(09.qQC*�e�@�� ��6rƅ ��7u$���d�2�A�Ƙ.	aКǩ� Cl��`�h9>�[gD��p�h��Pap���܃ _���bA@�LG�i@�a�iL!�$�s�� 	�G�A�B�9ǟ�`2"��p�DL &Խc���"+�1����)
���,���
�#X�S{� ��#D�09�M[�>h ȿ��%i�e�s��%��4m�����d�M��Or���gՠ<����_rb�LAd�'�!��kNl!2q�X���Tmޢ*��x"�Sǰ@�Q�.�O��(����nj<5B�ɒp8�U�A�	]E���E����![ט��	A���1�A@'��9�Q�H�!򄇚$FĠ�G����!	� %�dT,:>z�KaO�^�R&��z�O
,���u�-SȜ�5[0x�'��``S�V�n��(�D�@�̩�ƥ&vj6��S��i���US�3�8����L�S����/�����I�2�`t��\A��!�:f����1v:J����:�����I�s�$���jT��~�3�0XB�=	���	��&U���ORjiaaӞP.���E��	K��J�'#�����Աh���!���#q ޡ2޴{���8ň�y�4yy(O?7� �E��<�ڳd�h�3-ͺ-�!�E�2�8�۲��!>	�x�s� nA�ɶ5��K��#lO�B'��d.�U@զ��F	���'������<h���`9J�`���
P�`�'D�� N�wU
�1 %G1u0@�.3�7\���I��v2��0�ݤM7:u괏��	h!�$K�J$�H� �0)r%�;lb�V��<S�c�"~nZ�4V�B��7Lx�7eM�C�I��	ɂ�y����gްZ����8�A� 6|O����HZ>J^5Zb��,���;Q�'����s��M��l��2稉V�P6~�ҩ��VS�<�'!S���������l��Q�'Ȍ�!C)O�Q>�X fɒ:^��h���h���
*D��AH�tT8�zr/ϊkJ��Hq��Ot�IC�C�gw�O?�8ccN[_։ғH4W�l1�DZ(<�5/4W�d��I�?��0��ڮb��@�OX	d �U��� �@c��V8I�i��#W�JU�1���'7°J�F#?��,6����.�,p~�a�V>x�8��V"O�y�D��Df���!J�,7�)���CMS���$�s�0G�����Y�d��$��+>������yb�E�'���W��v�2�rg�����̟*U��i��k���~�<�r�rM ಶ��8Q|r��ōY<�v�<$`�u)�䈈P��	V`ĺAN
dA^�Lx .H�Qkaz�@!7vz���EI�j���bW`���0<�׫�=m����^�Tp�  0���	[1f�Y	W���y���
|%���qB8/���V�����(0���'��&��B�~ڕ�uU���Ɵ�(���6�H�<Y拖�*� ���ŋ�2����O}i�?�^}j�'n|c>7-)q��S(�"x��k�D�.40$g�;V7fB�IG`"�{��Rr����*HFu�V\�FH~Ӹ-�$吪A�R�Sa�|�?�A��2� q%�c0�!��EL�\�I����X�V�xс ��p,vd�'��Rx�$C�@�P	�jW�92|�#Q�'��t0�U�7�,ф��:;�H*(O�Yi�L��?�&�v��Eb[���g���d�I���3P�Jp@m8�	��yr�Ӫ`���9�ؖ&�F��<{W>�£��S_��9v�T?mkd�� ,��}޹���
�$i.T(�� ��w����dLW�US��� &S���Pc�}�P�J���Ц��'�jm��'
�)pt��{�1���-{JZ	3r�R��=����/��-E~�B��s����ɽ-�~p�bf��MAD�	^�{%�[?j�@C��P����(��r���)���r/B/��AJW�wNj�8�z��5Oz�qVK�4��	 \$t�i>鲑�Rsግ��m����Qk��$D�<9D�_������ѵJ�l0��oͳD���E�'o��q���~z��J��9��I��ɥg�*���� �x����'��Y���!�${�g7���:e�_�!���.��O�<�ቹ,ňA��V�xe���|�#?)BZ}��$S�NP���O��l*$��2���ȶFv���b�O�����'�y��ua���ӄn��|��OH�	'ȵo&u3��۵BC���4�`42d�ܲ";���g�X�v`�ia�"O��Ģ����>����ra����a�:��Ѥ�^�m��T?O�Β�O �ػЭ!��8(�MNu}a���=@�RӄYi��ڒ"�1ְ� Su͘扈��'��<���>��a��{1&���+�q����3dD�-;��݉5)�Y��1�X@�%f�	b�4уE+?���Oą��I�|�.�#3��_B:�8d�R8qM�ż����[i&(^^�O�����߶\�DP dfE����'�!`�H@�n�()%+Y��#"6
d�I1�MS�*����gܓ@Rܹe�%R��T+�	�ȓ2V�T2��;b}�=h+A�:�R�mڹ
�<�sC�P8��c�
%F\���@�_�4x�pb*(|O��J�G+g&�牆�
�B �����X%H��~B�	"�B�j���Xc@�}�l����'�-n�\�F�d�K��]��
�f���K�r3�'P��{a͙�k�5fN�[)���H�WV���J<!��>!pD@��||��X ��$h �OL�<�E ��ij,e��$��D8���KRȦa�7E��l��e	�J�Q�D^�"E�,�ĮW�a"`����"	lz�"
��<5�ːy�(�k ��<�0�,�O�<���k�Tu�#��Gs�ӑ�s�'p�H��d7���P��D2~4�⡯��j_,�ȓz!�0i�.�v����&��}�nZ5f�ބ2�}���i�v�ä��{��逽���3"O0-�I�.���tI��M"��I�]��r5���0>��ˁ�Pl�f�n]�ᯈ|X� ���G!�y��<z⼹��݁|����lY�yb��>*U2�K	n����!�HO���`>�h��RP�4�H��f�[P��$h�"O����da��V���=z �iþ�B����������O�e�څRF��.@����/��yc��r�t��/�Pв�X��Z���Ę�����'l�S�m�1�zaÁfWE���
�lJn|2���O� �x��aO\�<1�桒�+x� �B"O�e�1�[+x�ļp���Bo�2�鉁m	2���i�"m�\d��K�|��	�!K�N'!�S)�ƴSQA�	�����M��&	ͨ�*c�"~n�m�������=V����PHL�C䉉{�d�d�B�"�ġi��=���Sֺ���'��w�D����3!a@�@eU�� AJ5�7O�S$��-��PSĴk&eAS"O\9�G�"QP���&AT�Z��ɢnŠ���U�z��<���,b� ��U
(�!�d7PK$E6mD�Q3�\�_����O?HWIZ�^�x蓅�)ց�pR�<��G��8�ޠ���B�&��H�z�<	�!��8��I�̲li^��3J�a�<�4��1]&-À/�J��jK�_�<�ƠY�L��)���**��M��ÞY�<��b�2��!�M�|�Pi�-J�<��M�]�Ē�g�D�\���nB!��P�C"}ȀH�$	>�K�*��0!�d�I&x@��M���2!	I�!��Q�q��I�d�A�}�ܭBWH��]!���&=�W�]�� �h6�
��!���

A(@O	t�hu�R6!�!�ā�oa�~�PLӾ^K�9�"O`1�u�Y:^��4����|J��r4"O]K3-��RAL�Q4�2 ��(Ӥ"O>�9�펊_��l�F"\.8���J�"O"U ��]�	S�#v !K���K�"O<́�b�&D�`�"�ٽg� ��"O��Տ��z��h�BκR|N�#�"Ox,���D;(���с�� |��"O��0�X�S����� ¼f���q"OzH�����*G���oהR�:=�u"O�I�wCP�l�a�D�B�湑�"O�%����v)��;e�_�����R"O(��g$+u!|�֬ԔK^�;�"OD��ÃǿI,Th��쑳cYl��q"O �@"�d��t���Y�X"�"OHX�#dQ�E����3d��Q�,�$"O�i�W��K̔DbvB[���L��"O$�HǍ E^�{�!�P�����"O\����rg�B!J���-�t"O�ء2��01���o��[��p�"O$<2a�J�L�p0�o�2n��(�D"O8 s�LG������B�>�;C"O���V��G(ܙ;wK�H�T0�"O�(�0l�Z�Dк%c��n�xV"O\,�t��,$����b҄q�J�f"Oʈ�%�8:���c�����taxd"O���0�ǀ7��T��CҏQd�c"O ���9S'̹:a(�jl>���"O��ܬ]vd���=
,�`"O�����O.4}�ɱǅs�|��"O(,;1C���%pD�/gHqV"O��@w�Y�p���$6_��ra"O�����M(a��M�N0��q"O �0�Ôr�[X��,EN��"O8)���PY�)8D�U�P* � e"ON��� t��L����5�"O���ԋ�E���j�'�6,�`"O����R{X�0a�{g����"O04��e�::�� K�O��n_���"O�L�1C�f�a�&��;9m y1%"O�]F��\�X�а$<�Z"O� ��:tGј[c$lq���&c�� ��"O�c�/
�}�9��@�.V�0�"O�4��ݘ|:I�@�N�B1 "O
�p�G� DvU�0OPs�����"Oڍ�E��M���A̛Z'�P�"Oa{fE�*U��l�e��[�Xr�"O"2uc��4�K�.	A(�H�'"O�YK����:�3Ռ*472�A"O��j���!
�1j��c��Axp"O��ϗ�@�|}����_��ĳ�"O��aCV�P��PV�N�Jq���"O�Y�ϐ{��$YA���Rd�ʃ"O���W=0�ѺR��L� rG"O@�`'�Ɂ����bW�-����"O�dCD�7��m�7A��??ޤ�e"OTUSCL��'5�m� �K�lc�"O^����=F��F�-NB���E"O��� 3��t	�ڇL �`�"O�[��=�mr��ME����D"O�9
#���\�"�a���8��e�q"OP�[�L����G-�I�����"O�Wh��3:p@W��n{ yaB"O�ps'eы+	 ���/بK���	�"O.l�� �7|�jq/I8T��"OT��rM�h��1�M�_GT���"O�pHT��.
���Ro]�@G0�k"O�3��N(5Fp���^*/8�dB�"OxT��L&1�L��b/�AXi��"O2��"nY�s��"$@�*?��k"OĠcAB��b�
����:Z���
"O�{gG[���������hy2"O�� ��8%�,; 9��IX"O���엖+f�H�f��i]��"OH�[7��*E0���<%(J�+#"O��I�+�0f��=x�e�*\�0�"Ot���n�.I��١^��!� "Op�(��-:l�u	����Ѣ"O�5(���J$D��R�Y���qF"O��c�Nтr�ڲ`S��"h[F"O�8��(�|�2�U;(b^��"OEƩ.G��Q3.�t6EJ�"O<Q�I�=>/R`J���tZ���"O �ߎ��x|������!��R'~K�\a�R$B��t�LW�!�D�	]lp��_&���t(�!�,}��sF�LJ��Ti�([�!�DŬ8�l�]�&=0�yV臡Z�!�U)�\�R!bF4O����F�dD!��Ɵ~ˆ}H���j>ld됧J�r8!�
=;�~趡��Dݻ���;i8!�$D��m��%wP^�;eD94!�DU9m'��K3��;v9�����a2!�DJ�no�bUaD�t5���DmZ�,!򄊎&l���#ïv'��r�&"&!����bi"�.j����"IP�!�dP BM�%��ɫr��mY2X��!�D'g���p�����*f�D�Z�!�A;z�@U� �%'�e�4(Q�Q�!��,^Al@jʖ~re�A�_���)� ��9�&fjt=[c	��)��H�'$���A�<(h����@'�x��'kT�բP�6��AS�:;�8��'��|�g��m���rGMH�J�!�'�
�����]D�H
���/�2	K��� �4�eDYB�z�.uF�P�"O��`���.�t�6��Hf0�"O�@�3!N JE8����.(*`ta�"Of,�%��W$��!�n�bf��"OB���Y��qaA�*] � "O��H���>���3O"@�X��D"O؈�ك=q�HAc["Q�z=�"O��t��2Ŏ,���e��D�"O`	�%�1'��K�G=OY~��"O�i�d�ل=�4���KL�$�R"O�庲(B�����O�0d$X�"Oj�y5��z�3�G3'^h��"OfYI���z��1�/ÝÚ�"O���JD+v�R�#��P*�:,��"O�U���� �}��튏!�,T2�"O��toF�a�L�a&-ЉQ.ΥQ�"O ���ЇF�X����E$=u���W"O��d&��<�:"tW�`��"O��������U!���v��!J�"O�	���Y*�=Ib�<K5^�"O
�R��Pф����|��l(#�|r�)�Ә9pR ��:K��i�%؋^�B�ɥg�^(!�HZ?̚r���B�75BԬ��#\!��V�)�C�I!�p��u�"/�2��@�fB�I)"$�+`���}��٬xH0B�I
&U����.M�ča�܃{�C��[9R�T$ �'�!�a�tn�C�ɹu�F%y�(�?-Ƅ	�`�U;TB䉯��\j@!ֱ�B���6~ B��m�� ��Ö;s�a���MYB�I�u%�%��k#o��D��;N�PB��07�|�C��d�����X.b2B�ɴ�� Ba� Rit)����:)A2C�I���ภ�
}Î	�*�C)&C�I�{$Rd���J�b�!a��fC�Ɍq��!LM�p^�Y� R�öC�	/��YWě{ܺ��Z��C�ɽ+��Hb'�
�F� e)Y/*��C�I4u���-ѳ���HE-�C�C�	��4�!��ʼe$PYjC�N��*U#��nTrD�L�HC�	Aո�� ɕ.�`��	(��C䉘	�:��b��:_""tɁlݭl�rC��8r��ъ�6u{NLc !ܱX94C�	 l�y�5_3d ��iX�R��C䉆�b��g��T��Ÿs�ոQ��C䉢E�"�+f+Z�Gev�k���C�6B䉸?|.QI⯅�4Ɯ��6�@��C䉘7\�+2 �N��8�1*2��C�	�f8� Q�Q���*T<�(�5D�8#P`���l�����!k.D�|�������;�BJ�j� Q�-D�ă�l�?�`��v�U
��S��)D�����[;2r�r���Z��ljPH(D�,z�\�<�@��^�J����t,D��a��8a�!zB��(+x�)ʱ�+D��x����88dd#D`4�9�P�'D��C��)�=Q��;%'͌�z���'�
���lV+�����	
F ��'�*�*_�6N�
$��'R(�� �'�j��!��zTN�R�<8�$"�'�\�O7D� $��(3:2k�'~2�	�L�K0L����K'/������� �H2G;.Kf�����I��y2"O�yg�ƃ@!]*p��1RIj�"O���Ӣ�t��8�d]�RM�0��"O45	v�=J�i� �>B5d��"O0]��B�K���R@o֮;&�]�"O�x�Iۡ2���S-�A��]X"O�ܩD��s^��cËH8f�:(��"Or�h�U/FL��S�/T�"��Q"O`HQ����O#�M
��Ӵ!���j"O���)O�1��P�5���P��"O
����"����0��=!ָ���"O����	1�@�IF4�RM�"O��e�i��h{�G�4���Q"OD��f�L��9(@���a	b"O��J�-�/�T)�Q�W0\����7"OX�wB�=Th�HAW���;�L��"O$���_	oWZ�QB#��x���q"O`�3�̕�@���d�
j�Be�2"O����e�/p�18�l(xx��)4"O\p��:��H�E�� vY�"OL����2:�X�PܲA���"Oƈ�4��4[y	��
5�Ԭ	g"O6�@�ì2���֏x��� s"O	r�ꚴ<���f[(n�E�D"Op���䕘C9�����1���Rr"OV岳�W������)'����"O:Ј�BB/Bt���C�jp�1""O֭{D�i�>��7CW�O�l� "O��j���;a����]�?\!��"O��j�Jh�go�h�c"OJɛ��T��������273�m��"O���^f��q u�B�t.ZM�"O�shT2r0�f=(Υ��"O� ��V���[�Vv��0�"OzIC[4�i���2�����"OVEsKή!�$���Q�KG�(�"O���8u���Z��J�j�&�!q"O*iS�A3b�Y�'�W�x"""O�0;��WmÜm3e���5�ɑ"O�(Ѷ�.P�pX���E(r���"O4};u摪\���"D��ά�as"Od ��o_p�Ό�0o��k�ԍ
3"OF���eȎ v��;��I!x)hX�"O�����` ����]`d��"O�p��m�LE�A�҄Ўr��%ɷ"Or�A#ۉ�
2W�T	 �|1��"O�8�܎�G8�=�Ս�Q���J�"O�܂�C��i:���*���`"O>�2��v��|��ɘI��q��"O.5�Eϊ�h	v�i�J��D-x�"OB�Sq�z��J%ǵ��0��"O�1�% �=zbM�@�@4d�F��"O��B��Z�B���F� �Hh``"OT}���W��]�UI����5"O,�����K����EŘ�;�LY
7"O��±'^�<�!&Z�(bH�"O&xvLŇj���Cv�]U��X��"OƁ������H�ش���X8�p�"OH��L5�� �K��A$"OXHUgT�;MZ��A���q�(`:U"O�!����4��U��цQ��i2"O��z�Z:4���D
��%��hrT"O��*C�c�l�zsɔ�;�&eb�"O����%6d�$A16ꕨ/��ݒ"O� �	���F���1���A{B�)�"O`d�k�b�&P�b���Nc�ܢF"O.;1��!/谣���,D�8f"O6���)<Զ!����5"�:��v"O�IX���sJT����hpށ9�"O����ݸe��)AbW�Y���"O|���a@7"������*C(�H$"O"��D�	M�D�����L�a"O� p���_������ (8��c"O��S��ʇ^��0@2oǪJŤq�a"O��K�D����p�gP�e�@��4"ON�+�G��j@ ����W*�ZTY�"O�HZPA�/#��)��A�9�$	"O��#��$��P%T�l�R�B"O��qD�����I�d��X�3"O؅�$ ąUK��J�ͦC��Ř�"O(`:�[�!�A���`�)�0"O�d��
2iܠ����#^�=p�"O,��Bi4�l�n� AB�"OjX�dԤ|���x��%��\;�"O^�:�.,Tb�s�1_L��"O.e�d��-#h�ʡ���4Y�#"O��TlĭSJ�| �e�K��d�"O�+ǂ�740��C�r�\�S�"O<���y\aS���hX�"On1�QaɡY*��7��3ȅ�"OPL�$��)�)�|�Z{`"OԄk�m6b>~mk!��"����"OnQh�+�P��#`�7(iPLk�"O�u��(�-��=�R���K�j�7"O\q���'�y�%UDI,}�'"O�C"1�!aU���E��"OF��._8/�]��B�H�dXp�"O*D��,T	����P�n�6�� "O&��a�^)w�\��+���"O U`�
{Lq�*ByF�"O�%Se&�u�1ɂ�T�Dր�"O�=ã��:%׮O�	8�8�F"O6ٙ���"A��11W,3��{�"OT��k��@0�kLPt2�s"O��Ҫ
�_��]��d̕2���pp"O0�����B��=�@:��tZ�"O��!�մ/�AKE@��6� <��"O��p� -DZ�HJC�ӱ�ѹ"O"��(�5
���<�4�hq"O\4�f����QA��S�K�N���"O�p�0�E�<hh����/8���"O
0���W��'ԻK�QW"OB�{�b@�ZM�S�ӌ,�`�3"O��&�@�B��m
fW(P���:�"O�4Z��S�J�F���K��`�"O����>jm���_�i#Tm�&"OZ�'���	���DS��Y�"O�uZ�$��<>$p� ŕ ;�.��C"O����׾B����D��d�:�˵"Od��C
](�N���R��r�"O��"�	�@�ȧ�ƿ!���)c"O��p$�Ƥd{�܉4����:aJ�"O|c���nZ�)��-�2�I�"O,��B ˑ��QC���!N�J���"OP�Cg�o 	�O�7�C"OʱA'N��wmD�Q��\Y�xL�S"O! ����* x�ݠ]��ѐN9D��!,�H�m�Q;ܵ�6D�� ��b2��!XH%���_7�:eB!"O�s���I�*<j�)����P"OBE��I@�����"'��Р1"Ot"��9Q�$��m��v8d���"OF�s��P.�$����Ȏ (�p1"ONM�
-2��0���$a!���p"O��;���!�`�[3�N`���7"O�,
$�,/C��G��'�vE��"O����AF�/��E�,�T�XLQ"OVlX%�<l2\�B��/r��$"O�JՏ.�|�Aa�Շ��i*F"O:�(��H,h�I�V)�>"p�"O�� ��s�BdZ�H;���"ON���M��|��=<��M�#"O��y��1xP�9�6��Y�|�u"OH�5��W*�H�E�U�Y���"Ot��C�(�+��Of*Бa"O
I�D�)����%�2����"O�{ �Þ&���R��0RQ$�?Y�!�d�9:�q����f�aw�S(�!�˩ ���)ŠT1~�$����p!�D�;��eET���(U���Q!��<3��j�Y�z�2�����8l@!�d�Qv����m�V�q���61!�\�>-I2�ƖzR
��.
��!�$ÉK�l�b��FQ�y�`�ͺ�!���78���KZ6K��y�.Z R�!�d�10���9��ߚt0�P@.A�9�!�dەjg
 �tBǴId����N�!��$O� pa�	�<=��BŒ�'|�@(�7Gc�<8��"O�4i HU�i���R`�B�L�^�s�"Od ��,��#���J�&S��)"O�D�Z�9rHsu�{�J�2"O>���@� �8 D� Q���"Ol����A��L2,^V�Р�S"O|Y+�^�!lEzīB!�$��B"O��8�.(���B�K^,j�X��"OH�c�,Ӗ����E��p'I(5"O�0K�j��'��AB��č^� h;�"O�Lig��W���B��.~�J�"O.�bFCǬV̔��N�$J��"O^���"�&Y���O�9<hYd"Ofq!�ǅ=�X}��GT.���""O�TC�O�J�R��c��",~��"O��3 ��: �2���.C�uY"O���� ~%�${�E:z��A�"O�p��K�(s L4�#̳0��H�"O�d�@I�8���1�3U�"���"ON�� CB)!�������X�p�Q "ON��h� x���K6-]��"O4�YtB�27�y+Ń�� ��"Ob�1��J�R$|�#M<%��}�E"O��@oI>n�д���Ԫ¬}��"O�@�t$� H	����7!�@"OZ}8ЎO���@�5��q��"O�m����8�`
�C�`����"O��T�T�!g*@DV�LѠ��"O�lI�)B2;&�L�s���v-H��0"O��kS�&H��}��@�IZȢ"O��ZUFE8�h���M"<��G"O>�����259� ��$�z�x"O�j�C�5� �h�O�E�n̲ "OZXڎT���x��S���	2"O�  ay��ݧ���5�E�\�ZUp�"O<SW�ݸ
��#����@H9r"O�P����]Ք�1Ck�"3�t��"O~d�u�ٗsĮ=C�&`����"O�AkWdO�3-��i������"ON���G�*Q��ň�u��("�"O.�S���0pS� ��^�bt�l�d"O������U�L�b�̉0Q,�c�"O�IIV�M���5
_�_H�K�"O,%���S֌�P^aȰK$ܙ�y��Tu��� ��H�
�S�#�y� �=�@Us+S���\����y�J�-o���h�!�$8��T���yB��x=$z�+^t���)ٕ�y��d�(�Ł�5ePR9�)���y��[�)S(�4FIL�pAQ	���y�ú#y\[c�U�T� ��@M�?�y2oJ�z FmB�6�0%�����yRF�h�b�b���0���;��
�yb��3<�X���'\���a��yR��֞@U�M�%tؑ��y�>C�>�S�L�p&8��m6�y#ҥ} ����з;F�Hc�L#�y�GǌULP �(:נ[')���y� �)h�+#�N�Af��yVN��y�g�Q�V��G@�>�"�j����y�
��=�����͇:�N�D�9�y���>m����`�8�J�&�y�	D7n�|�s,PScT�ї��3�y�j(,� ����-txi8$��y���"zجKR,�l��Qs6I���ybA�?���%��kN���  ���y���KR�3Ңu5P��ɒ&�y�5!l�p�/�?��x�2G�+�y�G4(i�FkhP�b�K��y��؈UD�Rk^�+@�1R C+�y2��9�67fS=~	�(j�yң�v>)���`[�5[1��+�y�c�����^ۦ|�☌�y��@�G!�cO��V�"m�`BD��yBI�
 j��K���'G� P���ܟ�y�2�0��&� :*fݲgÄ&�yr�D(+xI��H"+���:��Ҟ�y��T�k:�3OH���lb����y���.0(PzPeS�b�F��q�8�y�!P"WW�az�	�6f�
D+���y�N�7a�����H�V]IT�Ͼ�yr����h!�:��:�!�>�yRF��,B�m�D��L�ai1���yb�͇r��AP�C�8H������y"D�
%�& �t�B"{�&��DB޳�y�]�(@��z���p%0����yBj�d{>̲�b�
g��-��_��yҫ��d��@�Y�r����A��yR��#=�2Be�ͪ=q���\��y�DF���¼a�,y�a
��yR��"��U;N�XY��b1��y�DS�{��U�g�ڲR�ܙ
v��D��L2X(KÌ5��a���L�8v�ȓo�*�IUdѕֈ4b"�� X3䔄�U�p-
�\�ׂI(7�Q�)��~�⤓'�P�Z�(�;�#� r0�X�ȓ'���g��e����v>�L��+@�A��%:k2�_��T@l�<� ���1�)ņH�j�p�5@"O��J�T�Q� ai%*E?W�A�"O��[W�� m��4٭2VN|�b"O�bc�-~/PH�ūCjتB"O@�jE�R�G+HPp(�9���f"O�)��!��&w�զ׺U+���W"OX�УG�H���C��(fN���"OHY������	�q.8v*<�5"O&��eS\J�y��A���S�"O����N<0&�ŉ�*y�v�"O|xRK2����K�0Q`�z"O�\�&��΁!�O]�R�|�!"O.d����"\s�}�w�@�CA����"O� 1�NMt���p�L�_��$��"O8)��ף/x��0*ٷR��hr"OViJ�J��`���:�I�/�Z���"Oⵁ�m�Iu|�FD/cШ�"Or�3uOQg/茑�e�L⼺@"Oz90v�X�T�ʄ)2�U���1��"O��C��\6I�X���e��L�U"OD]h�	@8+~=*�K�Pڜ��"O���%�֥?��)�`�/-`� "OL��s�ڟJ�Uʛ�|�� �"O. �g��$�H�FĊ�(�PhR3"OJ4�愍m�� �dE�<R��&"OD%z�E1+hδQpc�?rD�d�T"O�b�ѓ��ԀpK

��"O�ثMU-Ƽ��
[�A<�T�%"O^�/'{ ���k�<*:��)�"OX`1H���0A�b��A��H#"O�$�D�I�0��Ô�`]2�"O��A^�s؀��D52Q�X�&"O����G?8U0�(�lѫ=N*e�"O��+�Œ"��t�Q�T(F@�˗"OF�I��,1�8�a��N�gݪ�"O��;�K�O�D��U�� ! ����"O�1��A�2>,0��8I�@YA"OȕcR_G�Ω�ƙ3��u��"O��K�Q�Xn��ö̆�WDH��"O��j섰@ᆊ�@`
|c�"O2I���؏p���aV��5d(�	W"O�5"�X\�0xH�ؗg��:T"O!u98=��3�
@�t{���A"O���l_�),�Y���
VK�a�"OZm���A��A��x= H�"O��%n���)2��Z�0"DDQ�"OJ\����.��1�iF (���4"O`P��F(8���]�xa+&"O�A����10��`~͊\��"O��9�$,� ��F��2m�@��"O^�S��J��`�R���U�"O<I���*f��t� ��4�x�B"O����7=���Vc�a:b)y!"O�,��ɇ�i?��GA�2܉�B"O���!��h�ԁ&B��s4Q��"Or6y�B���F.^��NŪ-!�]��Z�QOP٫�&U�{ !�H/2ق�3��Y�a4��SGFG�!��F�(d��r� ��2Yd�%?�!�P���Fk�(�Q��!�$��@��Q��闄M�n�����9�!�DJ1[��1����7D�j���GF <�!�� !8�|��Fl�FF�&\�!��`��� �N���	�Mu�!��  ����]� x'��v=��H�"O�)��$��zd3v���r��%"O�����N�?b�x�.�>�xE��"O`阃�Մyy���r��1�.xR"O`��G3'5(��L�{����"O�u�Wꞹ?\�h"d*_�Qʆ �"O�xX�N��>V��IG��T�U�a"O~�kp+R��r�M[B>r�4"O*�È�j����e#��n8J	�B"O(�S�/�I�ʶ�##:8��"O�x���'�R��
P�4
f�""O$�ӒF�!X9�@1��L�^�<��"O4�I�+H���y�a����`�d"O��۔�1O � � �"��@�"Oxh�&��_r�SW/öp<�X�"O2� pj$�4<��M��al��"�"O|1Y� ֙x~�$[%�jW|�sG"O�Ps�V�g<�(�i�#aK�
V"O\
%��,_@H�D�W>g�`X �"O^}����=A��p�g+i�pbF"O�H(�/�5�@�2d8c����"O�M+�*�>��i��ͥ:�%H�"O���&�9hz�|bb�4b�&D�w"O���LLn�(�`��u�$�Q�"O�d˂��U¦ *"o�$<�~��"O$@;��f����������G"O\i{%A��5��0M_<WPza�"O���ҢY�p���cY����OL�<q"�6e�j8	7�"!F�P��J�<�OT%m�b7�@'U�l�0/L�<�e*n2.%�b��%����L�I�<1��*D" �q�D	`&�@S�i�J�<�2 ,�K��L�~�{�l^C�<�MUc8%a"hK��Ġ�GOX�<��"�a�So�p�={`�V�<ɂ�^6۲�FÝ�"��`1�Mv�<���23��8���O���EX�<�&��t 1����4�
#��Q�<q��m*�%�S!i��#�D�v�<��BN;n DQ�f�J4<:Ako�<�@"�;O5pY�ȃ�i��x@Q�<A�΄45<��@�.��s@�i��Jx�<��I�~��������	�}�<�3OC�k��}��-��Z"�K�nSs�<�������;7��i��кI�r�<�é�*�PԨu��H��$J�TU�<����*�YR.Ɣ8n�i �N�<i��0LX��S���h�0G!H�<1ǋ�?V՚q�/Ն  N���o�C�<1� �.qr�����?!Z҄Cg��B�<���K�Fu��S�7G��8$MZ�<iVH�<;3���r��5 P���JS�<�7.�%O��Aˑ�O�X}�f�	N�<��#.���S�)^<5g2=y�k�I�<y���� �8H˲f�0!�V	cA�<�E�N&�l��H�-?d.4I��@�<��	��"Ҭ96oΣ/��8'�~�<Yᤆ6.��ys�B�XfXhp&�S�<�6gS�Aº�h$�B�nի���N�<QE	C�?������	9�d�#cGV�<���6?�̨KCOQ�t�MFR�<�֫T�0��E#W�d�5�i�<�d�)ltAz���f��$���n�<�a��#F��R��&J��C�i�<� �ʂ��M �� ��c��E)v"O4akQ\�I�He�����w*O�d:R�� �x� �4u�L��'�`JG��]r��P��=�y!�'�Xݲ�˕M��@���F#~�v��'n$�+[�o����r'L�|䪭��'�y��Ɓ*A�"�̀n|u�
�'o���"=,��Y%����Ҵ��e��4(��^=!<�laD@��l��ȓ̼e����;v���	g�0�ȓv��sr�O5P�j8�6o	k P`��?��=��AT�Xp��A�w�@�ȓ<JpPs��� P*�@�����A<Ω�ȓd��s!�a�âCUڨ���Dמ�1��Dϔ,���D��P�ȓqW�P�?6���TH��.Q��n-�U��V�It�r`G�8]���j�����,�U�@� N!�s"O�H��[�1^��öeݵp�T-H�"O�4�l��&n8��e�,PҊ��"O��9���3'ر����,�'"OR偛a�إk�"W�qu2e`�"OJ�8e�T7�(��� N 	��+0"O
x1���3i��[�o�%2⮸ZR"Opx��/pv ���m�
@�Đ�"O��K�f�k�p{q�\�nL��"Ov��Z�J�K�+t�d]{"O��1�A�s��srk��F��A��"O���. ����:��	*!�Z�1`"O"�sq��!��¤
4Va(�"O��t��<3~F:���
{�jᚵ"Op`0�D0\�x0�Q�V5�m+1"O��� �N? dB��N�L&>�;�"O��o1T��sB7;x�M2"O�d�V��#�)Ò�5+ÎX"OD�"!�!�|��C����ٴ"O~Y S�_3F�ȑB^D��}y3"O�y��X�V���ۀ;�R���"O��H��C�9��R�Yw�P%1�"O"�{���+ ��Ѐ�U�/��"OZmC���!ف)O)�&}�"O�	Kt
E�$th��T�y�hL�4"O�\����G���PT�̱T�htS�"Olչ�;"�f໱C̎b�I�e"O���ʀ�N���C� S5[4B*�"O`-Q�f�\ؐ} %O[�2�"O�d��)CdQ8�*�c 5K�3�"O�u��]$#	z�����N�.8!"O�H�3n��9��ţflI6i ��3�"O�m���8C���B$k�\���"Odp�R�Ɯ*猑h��W%}�U��"O@�#s��/Q�ͱ�O `M��"O��f Pp��k̂-NA�9ca"O@��,�~V�زQ,�����"O6��s�I�,#��"f��Ȼ�"O�M�M�&z{������9T���P"O�D��o2(H9�ʟ�q�zG"O����*�D��O��QE"O"���㌄Tr�M���B�X׀6"O�`���2-�� ��j�&g�"}P1"O ��b�V=8x40� ��lr���%"O�<�P��f�*��O4<�2�C�"O����A�5Y���kU���=�*���"ORԪ��;����.i�*�"O�  ���Z�\y����jB�,���A�"O��J��.DL4:t#P"mvU; "O��� *ºM5رA���!"O�M�t��<���"�\�a"OB��gM�U9��I��{;�DA"c"O*��$	@4P�:sHJ& ��|��"Ol����N�`PH�XE�@N��I0"O�4��\�H5���=3���0"O���n�3'��yu(&�"O�t�I	�B�C�iT=��u"O(��#`�8~�I�w�[�hH` �u"OV���� s�$��p��H(`"O��x�Q���1R:���"O�$R��$]F9뇣��6x��"O�a�˃�
�Je����pE3F"Ob�qd��X�-�V�U���	#"O��k�(�#NV���A�*u�""OR��gW�O��9 *F�c�p[s"Oͺ��_�.H��J����`%��y*O�"%�N���JV�I��`�	�'�̴z�ږ
�v�+��]�w:�H��'�:Lx���+ �Н��b�0D�PK�'��!��:12�uQ1Č�9�h�Q�'��	�kq���p'��,�����'-�x��BN�z�.�[Sc#�\��'m@���H�[m��ɦ!gH`��'��N1
)��R�H/(!p�P	�'F�q84��s����!d7+^d��ȓ<���Bǉ)]��y�Ƿx�J��"D��x�ƅ
���!J�9���,D����&��q�Q�݊)TTr))D�`"v&�>q��ER�"@�,z��2��1D�p��/�M�xE�F�%ZT5�5E/D���"�~o�pc�{��M3�N/D�P�c�ߋ1��㇈�8n�ȡ[�!D�r� ��5�Eg2u�z�f$D�|Ȗ�[Pl��R`ғr���`B?D�t���&5�tUiu��D���'�=D���1�>�sv(�W���XE#;D�A�$&t���s ��8��c�4D���T!�0g�d� 2'ό�P\J�o-D�$��`��
��C�m�~W�3k6D�l�q�Y�2�"xkW�Ӡ+BbHf�4D����CW����\�4�J�ɲ�1D�d�Go@�p#8EY#�;Wj�j��1D�@��6Mr�(H4m	���y�P�"D�t��[�+��U��f+4]pa���<D���TCI�pc ҧ�B�!��<D�pQ�E\#`�;��ёl�؁0)=D�hP�OT�	����R�4��ѐ�D(D�p���O�@D �@i�3y�|�Y��*D�`��J*2����$���\�L���'D���P��(Htը O�.�2�H �1D����%7 Ac�� yYS�*D�d`�:-�c�e�z����`)D�T���ޮ/���[��Z�I��*��4D��SdJ�b Bl�b!רX�x͋�/D�t��"D�xKh=����C��u@8D���u�D"u0'L@�@�t`y'5D�D+��_c�c�AZ.'�@��Ǥ1T���!��4<L��R�I�eX�0"O\�K�
�6*��2�P�M�Xp�"O���۬sh�V�R2}���+D�L��uH��2�
a��QD�<D�� ,��L��[mx�,��:\6�x�"O��V�ׅ��0�ˏ?-9`@Q�"OR��P�M�6��(@�CRf�۴"O�	�%� i��3QOR� �[�"O ��qEĄN���@ծ�.���RV"O�u�
&�ܝ��-���AZV"O����
8J�PK��ߙp�,���"O���ӧ1#�``���Z�~����"OLUA��R��6p��P�g���5"O´�cD��}��<A�l�3Q�j�"O����J8c��pCta�&�Ԛ�"OҩGC>C�z`AYu8�B"O���+1W�Prq�F�c�"O��Ak�'�\�d�$TL�C�"ORB
����S�I_�;0 �V"O����'�o*d���T�B}@���"O&����J@��TÝs�j�i "OܤIg���yYxp��D�,�D��5"OΥ�d�υКd�wI�:�Ή˃"O\@���(tot�P`�?H��B"O�Q��@0Be��Yu��90�L+"O�l�"�øXv8iCG�r�z"OF��DD�^�b�Q�Ȯ#�a�q"OrU�B�4�@���o���� "Ot<�7+I���%��7u��h"O2��0㎙z�Z5AU&Z�v˺�h�"OԀ`u��_�Rg%2h��8��"O�(�d��#�2���T4zeZd"O6�k#�G�{݀Q���L� Lа"OXH�/�GIu"G�W#g,uK2"O���Q�;=H,S��IU)�l@�"O2��$YJ�Y�nĔd���"O`8s���9�a2gߜf_b9J�"O
�sF�^�?���;aE[��&	�"O ��E!u�-[�"T+e�\h�"O�y���1vB �G���t�j�{�"O��� L��a�J�İ?�FU""O.UB�P&|^*Q���%1����t"O�q��5L�UC�Z�gI6�2"OD�Q�D�!)��=ɥ�3w/�0�T"Oe7�QN�p;���?Zp�"Op(iL�6}K3�Ο� �"O0�q�G��\�t�+��E�f�Z1"O�����+fج2 �<�L���"O���2�ŽỲ�g�� n�`l��"OzĢ�n�y}:}挏|r^}P�"O&MC6dX)k���"�E�#D �(:�"O$e+Fl�7���&�n��W��yR��$����#�@�d��f�O�y��=5pxVK�L�6�)�����yBd����<U�ߓZ�b���]��yb տT.x�j���N���$(N��y�o���H�)�D�}�$���'E��y�i��=C�<F^f�E�����y2JŐ{\���B]: &J� �?�ym@�M�.I2EȚR���o�?�y�"�2*a)%�5�@��I���yB�"a����eʗ3�) 4'I��y2�]�x�H��2B��}�PG��y�h׿<�4���L�iQF4�7c߾�y�d�,esp1+�7Q�}[�o�6�y�5��Q`��7D��&���y� Y	b�T�٥��4�`́�+ ��y"C�jW x3ׄL�*�H��<�y
� v�#E`�/R�"�w���6�, D"O lp���e�1��L3� �)"O����
��a
#�`I�"OB!�7$χWJB�X1OHi���"O��`�$��v�<�j��X��P�"O(1�P���,;���`a���
�R�"O�`kG���f�H"�"h��ɩB"O��҄H�j�\���+ܣ�Xd�S"O�i2�.K^�� 	�*E�Tih���"O@U�U��R�����H�</U��"O�}
G���k�zaG�G�a�"O:u�EI�e��dߡ>��p"O�m���$9ݙ��Ř=�x��"O���e'9\���;�E@�b�����"O�5ړ��%,�HP�@�<����"O��4sHݩPƋ�4�1"O���@)L� �Eٲg� P�A�p"Od%�3A�55t	z�L��H�v�B�"O4�6�5��t�Ǎ1:8�)�"O�5�@-��4����FK�ZR(б"Of)�FHT7'�.Ezd��;4|�5"O��#�	)p$s3FR�Y�Z��"O����(Ӹ9��
��I�لb�!�L�>����m��JN���j@*�!��]�3��yS�f�44�H��
��-�!��ޒcg̥�U@�/3"���j5w�!��.h>��3�X�%�Läǁ;T�!�$�d!��`��9$>�P�Ʊj�!�$S��1A��W��L�q�ɢ%�!�dO�o�h��	Y�4ga�&܍B�!���w�,�"pL0��A��<8�!��Q�	:�����"|���s��!�ρL
�H)����F�DJ��[�!���"��3�$�>Xh���)�!��+�,ZQH
;N��VM��!�_�~$��C�-���'*�!�䛢F�x�)��!r���l��HB䉐��lp�ˁ`@18���8?:B�I-2�zUa�ȥHq=���
�zC��/i�`�儙8$m�1I	�9�BC�I-ޒJC(T�[�I+�ğr�B�	3 �8��r��=K��8 bgf�B�	$ZxB�����q�����l̸t C�ɭZ �%(�d�=/u412EE��!�JB�ɤ��1Jef�]�$��%z?LB�I4P��+EƉ�D�UY�_�E�BB䉚 H�S�'̘
�����N\;~�B�IM� �QW
ԉW�zɃ,>4B䉄):n-�f*�'�H�vI��v�RC�I#x�.�G)X�6��aEv3�B�I(1�jԃ���#�Ɯ�-ɩJHC䉣<�4�;䡄)qZtD�$�/?��B�	<7�@��T�ǿK=$�qa�fsJ���+�X� O��/��sW��S�A�ȓUf���G/s_G�	z����i��L:1��)[.�ă��Z+j����ȓg�d`Q �U�K�.ŐeP�=Ѐ�ȓm����T�b�,=)��$�F(�ȓ&���1�A=%n���s�A���*D�$�Ş�]Ϻ�1'D�!Z�+�g4D��%Z��zqY�I3(<0�N1D�Dkd&�6��;�(S�@�:��/D�X�w�R��Ɖ�2%�$b��+D��&KB�D��5�$����0���
=D�� p��ӭT4ra&4;�*\�A�N"O��
'� s�R`��#��u��"O�pZ�C����iW� s�J\Z�"O~����K4G��4J�b��
����"O��(@M݇1��$ca�Qo�mC�"O���B�'�艠�NӬP0�5�#"Or!X����&P�[w��"O^X�c�6+˴�Y��S^^Ih'"O����Λ�XBԁ�"Ϟ49Lp�R"O0��'��`u���$I�	:"O��{v��'j��P	࣍�L/M�s"O6���R�A��тޞF� x�"O
�'
^���Ѵ��՚�`"O��5*ߨT��4�rԓ5���q7"Ov,
���'ܘ�D��,�����"O�ҡEϙ)L8�K֚z�r�6"O`�!o(~���'&�|H3�"O�����B�AJl<Sc�/��q�"O��)q�ߕc���;�섅��pV"O��ApaIvwZ����Pe��,��"O�I6ϖK�2c�ԭj���`E"O\�1�<6�����
�����"OD���D- (�,�"�T�"O�i8�+�Y��u2�A�{����"O6����N8U�^�	E��^!U"O	s��)肴!�,��[�����"O��h�O��wh>Z�EQ*\�)t"O�,�`g$U��A��y��"OΡ9UZ�a�!"D��HLp(*�"OB��q�۬37�4Xd�Y�u�ӱ"O4�!��?N]Ѭ̤7�r���"O���B�6n��Y�,�%W�*�[�"O��6-á��y{gP�|�p:�"O�J�U�v�%���X
	o�Q"O��3�WX��h	��Z\�HQg"Oh5�R���q	 %�gS7o4@Ap"O���"E��@D�H�N�b	�x�"O�u��aB�EޚMӴdT�M
.8��"O����R������2x���T"Ot�cڄzT��GM�(�v�4"O$$�3h�\�&h#b����	�$"O��p&mE t'�D�di�^�Vq��"O�!r��j��4HY.M֜#�"Ov�����ER"Up!B+��3�"O��M�,t@ȱ����a�c?D�x��d�z��oB�a5X��>D�D�P�߆Ry�i��:u��`�<D�8�dA��"�c�3E��i$�:D�� $S�K�\�O� ���ᶥ2D��5�
67X�
&b��	C�*D�x�T�#R&�MRu��-Or�B��)D�@1 a��������Sm�`�$D��#h��T�4���D�1��˰�#D���B-42(@h�� %��@36�#D�L����+���@#�� -J�!4b5D�����V�L����$� bb��G2D�<�e���HTH�	W8Q�B0��3D����,S��T��F�� J�yP�6D�X �j�le�`c�L$�F�p#6D��p��$k6Z�;g/�'I�`��f3D���!�ID�U����t�W
0D�� �.M�qqv�As0�v:D�����N� К��cҕ5�*�
�/7D� �����Ar0ą*&L�(6D�� �i���Y�J�rU�ƍk@���"O�=u��>"e�O�
��`�"O�q��n�����O�Z�<��c"O�8�b��#,�p�+�M�?D�)��"O&X�#�%
nLP@Í��:��r�"O��d
#(�4}z�ʼP��}*�"Ol)�S	 ��[��OKŚC"OV�w������� a����@"OL�����O�d]ا�j��,�T"OBpPa͏�8���*�HvP��"O�* ���L�n �0郍]xIg"Oɢ@y��i  h�;#^a�1"O��c��A]ϖ�J��
	\�EY�"O.h��	h��	��4��<�s"O6�ag*ěuQ���	/2���5"O���6B�J�ˁ�O�h�Jp�W"OJj�F-Ҡ5��ú@0�0�"OD�[���vG�����=s�"O2$�ď7(�>1��c�:Q/��p"O�&�	��α@u�6TsV�x�"O ���@	�4���];4p"$��"O���C�/��\�6NM� QZ��""O�����һ{j4$X\ʨ�"Qn/�y��-��%s��B�^k�0q�� ��y��)I�����-T¸�@�Œ;�y�iO�1.�+'hL� �ڱ����yr鋥r@�٧�ń|!&��&�ˋ�y��Ջ|(T�b�	��D�0��m��yr��BZl-kS�
7��D	���y�M�#W6��Y��Z�8��ٔg�'�y2-W=l�xh2- >-240#	���y! �2�8��t.B�:R��`� <�yb��89�.���4g�dx�'���y���n4��Ѐ�ɹ+�ֈ���	�y�m�'1o�����*�=Qf�W�y��������AB���HƆ��yr`�T�TYh�MS�$�DM<�yRN��%�W�@�R� �5,P��y� @�jA�K6E1�����	��y�K�]�ᐡh]!@�4�	�e��y��B�a�F��a��6�z�3R��(�yBJ�a�.��4�Rk1f���yb�H��䰻U�S0^�Q�a»�y� \�{�����敢N3�f�ܵ��'�t�_q�Y��ҬR�\�k0�!D�`�鋮`Z�B��ԉ;�@#� !D�T��D�`F��+ ��/A��DZ4�1D��h�����nXbt��"�+a�$D���
A�(��ܳ�B����9s�#D��`���J]�)�$>��U9�A?D�xe(�TzθcAΤDh�9t*D��qQ+z1*�p�iW�sy�����$D�4 �
ߚH�TI��d�+�M#"%D���4�+o��jb%�,�f�iT�#D� �`�=`I����_�#0����.D��� D�j���hޠĬ���o-D�0�dU��<AW�F5ug�-�2k0D�����A`�ࡁ*�$\�B1��.D��q%l�k����"_ pD�kf+D�������$۰��W %Q���pb�;D���֧Ʊ*�J,���$6aP����7D�0+Ƥ%\W�)�H[�\�`a'�5D�b�I-8�d-�`!�*!~L9�5D����#(���Q
}x����3D�� L��L�s@Ȁ�!��B�\B4"O��#�I2���E�t	W"ON�0n�����d�&>P�P"O�q�S�^���ـ3��6 ܨb�"O�y��hA�P��	���M\`$��"O�q�2+D�.|���"O:Q�B�)��@��e�i�24��"O:�����P�V��&�%$��y�"O��1(M�rQ��t�#7&Q��"O\bg��f�����5�ذ�"O5���І-θ,��� �l�2�"OL�1�Ö�o�zi�7-����E҆"O:-˒��R�Di�bW�]]�|HE"O �ԁ@<b���;P+��tSpxS�"O�4%�S�V]Xث�)#"���CP"O$�2V��L��m %	�L��J�"O���ư%�]�2��5(�֨ �"OԵ��gl��"��B�|��M�!"O�}���6!n��[�e�3I0���s"OJ�h4�
�3|z	3��o.$h��"OrH��
B ��@�6 ����"O��8f�MxL sÀ�w|�6"O�� Į��
�`ďĳc��1F"O
�rd�G�S&`-ɤ�� J�Q"O���pe�TT,ԿnZ*5 �"O�TʗG�����Y]�4��b"O\Dj�ߣN���˞�z���x�"O���%-�9P#t`�dLb���&"O&q2����P�R��1%vL+�"O�1ʗM�<V,81Q����h��"OxD�B�� %��M�����"O 8#��-v9�2A�R"r�|�t"O�ja���,���ւUH��2"O�y{w�K���+��X��"O��kPJV�a�0Qƪ�	X�j97"O.h´f�!o�S`�ͼ!)�e"O�h�ݵ"�&p���Kn(S"OB@uE�� J��:3�¨r}��"O��+�=z��H� Y�ob�0�"O��I��K�v��A�!!�p��"O����
�@|v!h���d���k�"O��@�G�g�)k�;֖�	"O�����׀��p�4�_
Q��	��"O<���@sg��g#¡O��9F"O.�P�CA�#*^t
�!�g0�+1"Oeٓ7W �@��W����"Oyq&h��?��QP�� D���!w"O�H#� ϴ�(����|?�0��"O>��4���\�b�kS�0���r�"O��Ð�k֘��)o�H�m��y2,���B�0E��L��Ӡ߯�y��V:�P�%�@�}�"i �y"@ �Q�8�b �bo4H�5�@$�y2���z��)!d�
hd}�3�U��yr�?pz�^2,�rC���y�8A��HS��՘]a�\�#T��y�j�nЂha��ƥT�O�tWl�ȓ6|�`aG�I�����hܤ���c��RQ�׮.�9���F�2�t=�ȓ_T���S�$aC�Js�^a�ȓHb�f�
�vO:�P��ҍb�d݆ȓi��P�jj���J�4>h-�ȓUW4�s�#Ȋt�����M}7�8��6
#�ڶ	��t:!��@ ��S�? LQ8��H�#��A
2I!q\�c!"OBlct!�q�|a��.����%�"O��&J�7.X%
2�;>K0X0Q"Oz	Q�GU�p*l�1uf�7�v���"O���&$V�T�8U@P�J7bqP�"O�u��� QJ�Y�GͻjIzD:�"O��s���Nf^��F��t��%"O �FI�:�����ѳN����"O�$Y4HŦ;���ˣ��d��R&"O\K�O�89���耋A�j�LŹ�"O�-ش
\��	(��67L��"O�h��#ʜb����v�0TI�A�"On=Ia�))�|��A}=Z��"O$���I6�L @�q��@g"Oܤ�V�:@n�ԺGn��*����"O������D�CmلI��!g"OT���E�%-���[M� L�Ĵ(�"Ob��� �d��M�<�����"O&�#���4納a%��'R�`r"O�p��$+6Aps!Պv:]�Q"OZP����ܢ��v ����"O���DOQ�t�n;7 ��*��"O���"BLm(�$�2<�\q�"O��֐Q�N�aIڊO�H�"O��bvNE�R��E�ć��-�L���"Od�(��,i0f탂�U����R0"Opt󀭆�yZ��B'�����"O䜲���9)����P�D�b���"O��s.N�`U��ĉ�4yy+�"O��R��yf�L�GN	-<�8��"O[��!̅u�6�W�}�,�g"Ozl�A%y}64+@�S�L��D"O�ctf��}�%�VnI��<u��"O A2�L6=[��o��D߄��"O<d�%"5n
h�*ģ�72��E"O���� ��mر�_�`0^4� "O�h�"� Ah6��e'ӝ["��bc"O�	��k̸jJ(@��D�F0R"ON�x%*�0km,e2�T!E�&P+"O�˴��O�(��B?|�X�P�"O�X�-�!Q� ���<��r"O�<� HS=�t�@gEh/ج�"OP٫�G[U ��T��=��9�"O����N)
д\����7eG����"O���P-T�&��a�\?5b,�w"O>|�t�P�Gmf���GZ:G�3�"O� C�a��%ـ��Ȃ� ���7"O�	x$F�(</B�!��6?��})�"Oj$�£��B*�fpP�c�	5;�!�DS�z��M����ayRL �h�#[�!�'!B�B#.S9q��¡�E�&^!�d�(M��Ek�j-'͐�;�وQ�!�D��K=ĵ0����Xdo�>�!�dF1R̮heBV�a�Z% W�!}!�$ m2q�!��|H؍K�#T@r!�$P�,xT0��,��,LP��fCC�[�!�Y�D�P���&B5����0�!�D�	l��!��R�5��Ȱ�
$�!�D^�k�B�#Y�$R'j*H�!�dH\�ڼJ�	�D�=*	��"(!�N%z�L��"L7�|M˅(ҥ!�B�<{w�ԑK��)��a!�dšK}ZL�E���>��-÷�V�kf!���;]�\�f+U�?�|Z��qP!�� ��%WG��U�گk�&�i�"O2�B�G��i�lꒋ�<��P
�"O0�6jZ�3��仠OA<����"O�i�6ƊbP��ƭ��� Cv"ODm��˙�s:����,�+� �@�"O�@��Ff���s��.q����"O�
�����;T�#|�B�Ap�<A"*֜pb�pCW�H��`Q;0ɛi�<9��	/pP���@�X�u��y2�g�[�<ek�CT.��g_37��hQ�SV�<�U��2�Zp�UxT�QB�H�<1�d�7X�N\�C�(Dh�Hxa	�B�<�7��/Eb���O��
o"�� iI�<��Ɛn���y��\�U��e��#P�<�𠗳D�������jAb$��J�<��D�;8��
��եj]PG�q�<yP�@�,��pⱅ�r�z���END�<��Hؼ'y�`��+ѿ3~�(D��@�<���W�|q��ip���7T1�%{�<�$������I�P�X��t�<�aU�>@�5�Re̾"fV�H'��Z�<!f+	)p\hp��J^duh�S�<�t/6�P�T�YUmMht��e�<)7�K�o��B5f
S�Ԡp0�i�<�nH�(j~�����  �@PR��J�<���W,T��I<��ѓ���I�<9��Z&z �������|#�O�}�<YËI' 2���TN�[��۷��x�<� �ȧ)���")CJ��ѦMr�<v��k�$�Mrd	�$C�f�ȓ&к�X�*ǹnY�<���V$h
0��ȓ_&rmy�JO�~n��Z��TE�ȓX�6�сMF�f]�A*�@���V���YP`��?�`u��Ǘ��p��xM��l:$��U�%�@9��E�R�Z��v=�"��~�<��>,(�2'O**cy�T�f �ȓD��!�3~.P�v�F��dU�ȓlO�r3)G�q2ꡨ�-��z|���6�ۇ�؎mj���6iѝ:=���v�Q[�H�@�Xq� ˳7P5�ȓs$�P���@��dz'
*mh��ȓ/�2	[���#fu��l��<��ȓ}��d	[T(���͌b������Z�q�Z5� ��-�>�T�ȓnfj��b��Oٸ�[�������ȓ0\5)�
���� l�60V4�� h��A̚�@�<0�/A�D��؇�a�8���
}s
���W�%���ȓi�B����+V���m�!Y
���M�P�tE�+S��\B#�Ĳ
К���2l*�oN��RQ��,cZT�����<.To�pu��O�%G�����:����Co����P�U���#�PX��r��r�	�\�,�LX�v����ȓ\LX�i��ڢ\�.�z��
�hl�ȓ�:���q�Be���݅e����4/D���&�� �&o�>D��ȓV#�h�FLz�LU�n��yN蔇ȓA�����V�W�u$Ň�b|R�@�i�#k�b$C���	9�
��*�8����v�fA"#͊K��ȓ��Ȍ>N>��Si׿^����ȓXۨE�Q/'DnK^�&|:d�'D�� !�`�%X��0��s��Д"OJ=���ɖ|�����B���Mz`"O�| �%ͨ�NX[����pyX��3"O�˶	�����ɕ�G.$�B"O���#C�ӄX�U������ "O�MS�`�X%�Y��U�I���a"O���#B�t�h!����Qچ ��"O�XC�$W����Bg�	x�F���"O ҕ��,���6�W�T�����"O��C&�K��$��Q�-�(YJ�"O��x�o^��c�E(%`���"O$�(�S: 9jq��nQ�~W}�4"OB�w�N�SC�p1ůA;2P:� "O�`���k0h�vN�;n.`��"OddrebJ��(� KLR��p"OeX�$�9Ŷ�{d1@�1�"O��2����Nd6u��'̇ƺ�{�"OFDq!�:Rs"U��g��L����"O������"�䙭I��1�g"O
��j�orb�#�dO�K�tT��"OJD�6w*d	B�Ú4.�R%)�"O�7��72�̌�%⍕;x��0"O"��B�ՁzT����4Mc�zu"O�MA��_�T�C�Ըe�p�"O�y7NA�Lj�I�o� �YD"Oɳg���-���4�4��A�s"O��g�P�ol��3bZ�#��� "O�q�l	6l.A��X�es��0"OĘ���P	�ٱ�"��P�G"O8 �M��@ǺY:�I8y���)�"O�Ԡ��R62�A�`��|?,IѢ"O�	�Lݲ|�Jɑ ���]H5r�"O(E(Ƣʈ|�6�:2a�1nF��"O�H
aiү@�!�o0���!�"OdYYE�y	�= �űq��`"O\�3���d��Y�67�"O��)2⊍#�P��$�H1pހ��"Oz=I�(��k?��K"�O�R����"O��Ydo��L,�� ��%L��	:"O�����ĺ8��=)���I�T՚�"O�uj��2| (����!{uF�"O���Ḵ��"�͓1�hAP�"O��02)S
<�X�S��B���"O��aU���H	�P�P��(��(��"O�<Jt�Ji�t\�cBHcz����"O>9r���_"
����,��sd"OLaP�DJof\�z`a�RF�Ɂs"O (�S&ĭHJ�
��6W��J&"ObH0o�7fI2�P�NX=�"�9�"O�uB&�Z>TSx�)��e^���"OR�R`i&���$_D��xS�"OLMc��*kr�ģ�t���P�"O� 0��2S=��+ �I$.6�-q�"O����험XӞ���NB�65n�p�"O�£ W%"2�x!��?P��"O\̨�mC�@���XQ�F�W����"O(�˳$)�P٦�lu���"O�!����(Y�*�.mR@XBw"O%��/J��1�`̎�k3���e"Oa`�&��+P�U80��"O�9��M%!i����G�U)~�	F"O�d�V/,\��2���+��"O�TC�5�~a4 �+BB�`�"O�� b�bS|��D�_)k2��s"O� ���2K(. �5�i�(k(��4"O�)4�D1>Ƞ��ĜǸ��"OH�që܃���*��,I�>x�"OZ��ƥ�8�B����(:�t�+�"O^(J��F0k.�5Y�Mys���@*Onh�$.�@�!h��-0�\��'��p�	3P�l�E�W/S?��)�'1�|x#.;F�ݐ�i�%9����'T\�'�� rG�$�`J!I�l��
�'\���B���(�2�f��jRQa
�'�h�h�f�,�}6hF��:�a	�'�Du
QI����S5p��'}�<ɶe�#L0�IƉ�$5j�AB��u�<��K�X�9 "��������r�'R�M���J$Z�Ib�x��A9�'���q`�ǲ`����	>z�X$p�'"j���A�jEy�K?p?|�h�'��e�F��))�D8� �w�(5��'K@���e��J��0�GD�:�����'�LL�S#צ@
�$#A`�??�h��'0��B�7g|8kq�H�`N\�	�'��kUeϟo4�$� �E_$}��'cf�9�E_�h
�gτL��=��'R4���/=��墡�KT���',x�G�ݞ9�,�-�~b6���'r�Ԫ<0|�ͪ��W8��i��'�(�8�a	 &�zTÓ���>6�B�'�&�X�M�W����e������'����%_[��ٷ�ڋ�4�{�'W���TdR�ǦS���r
�'���Ä�4���_�bO��R	�'���Wr�5��d�8QK�'�4��w��.�]�D��R����'�$a	VA��L�!��8��,Q�'�ĨRc�*���#N�M��I�'��q2"���XR�;H^���'��0e���H�}A��w��t8�'�$pàBM�H�LA��� i�$K�'�(
�oP& �����/W�U�&(��K�a�a
�[�0���gK+K��방��O{┆�IW�>���-�����j)1-4�bՊq*\#�!��[!E�V٢%��p�t��	��B��,���se���uG���]j� �2��dߤɐ3���ykp%�C߳e� I9��*�5B4b���O�b�U d�1�1O�� ��׳�2HѠ�_6�4H�4�'2����۝2�,��5��6!HN���O�{>��aS�C[�`
�[�&��$�ρK��q�mV�Q�D"B�5<:�:w��]�tH��O��Sh��W����6X(X���'`�|���WT�h��=T3�����j.x=P���r��+��*lf�tF�D�F,t<��+�EK$��FK�!��΋��p�C�]�$����B�8������&;ܵjb�X�8"R��cX?�Ey�hF'x�' �*:�D `�ۉ�p>�#���m!�)�a�Qx�y �+�,h�� ��
.̂5yu�݄%�l���'�����͊#f�t��/]� ���K��d_~o.��G
IN�đ0e�8X�y��O�ۅ��� c��Z2B,��X(	�'��z�ј*��1��]���@*�*4h��1^�$��Uή��F�$0�� $ӽhn��h�"N�W�l�xS*Oи�DGV0)2���)P��@i̩Hqfӂ�ޮ{|�
�����t�q�'`P��f �I5�D�s`F�t�	�:j8xa��mJ��f��p1�5(�̧�(��� E��r|rǣQ��t��I��x�"P/K4�Ep�kU�F� b��B�hQ��|(�ej�>{o2�pǡ-V����6"\E1G�� "�|��pk�h-�ȓ�4� �6m:°Cs�XZr�|(�H��z�T�V�͸3h�9Ʌ��0c?�I�1�q�E˗�p�Ӓl�1"��F"OJ�@�ʆ{:�9��P�����&	U�F�\��di3�,[�k�J�ʄ�(O� L�Y��6!\YB�
 TL�R�'��`��(����(J�̰<<��An�9L�|��Θ��rѱc!�4���*�O�(bw��<vU�mC�0���w��W�{���ԥ�8l����ӓhl��7����-�&ѠdK����fL�9��Uo�<@'��~��LRT$ǯ���aP��}���)�CNd��p�	�]d9p ��B�Ƴ6m��.��qz�'�|!!�D���!t�I�儠S�,OX�ұJ�G��0����(5l��b�Į���y��d֑z�r��X�Aô1H�E�&8��z� ��nFIIiO3\M��S��J8Ǹ|�OԱnQ��q�����ȸL˶�a}2���z��mq�iC!e\��j�0Ӹ'C|3�h�+��K$�
L1�r$G0��ʲ'�5�fbY)A������
�!�$�'��	��Nj||�cA�N��`
K[{�͑�G9@��qP�S��y�o�)��  6�h)�f�A�_
|�ȓ}�: P���8cܚ���l
%D���爃�4�B��m��*��@b�
�?�>YС�,B�!�Ą7B>�q�fFAe��a�41"=��KP���Q��E;t�x��C�^B䉢ewd�rӉ@���(_=0��<	c. �du`�z��ө7�F`y"K��i���!_�o��C�ɷ]�ªmcX�Ct�C'b�t����<�f^���JL�IZt���.�s���`n��ϛMu���ȓ^��)Zf����0����)����ȓmQ�rȎ$I�x�N],p>���f�R܃Ņ�,%���M
�*s(��ȓJ�+1�<���t�#Ы'D�dj��L&֥�$(�,}bX�y5(7D�`s�D�A���db�����'7D���C�W<rJ
�a��$p2��V#2D�L��Ȃ[w[&��~
�țg�'D�$�`�Y�f�АT�~0"����#D���S.�"�x5��F�kM|Ib��2D��!��?L���a/�1ٌ�� @5D�P��ˆ#�Ht�t���3��#�B0D�L�����0Nl��ih�4�TO1D��j��C&�\����	�(��6�.D�
���%v �M�.����!D���G)M-��Qg�����c <D�H��k?��|A�G�V�Ľ�S!D�P���ԅt ��z��ďmL�y{@?D�di�Æ
#��e��A;�36s�̈́ȓR�bٱ�h���v�\RA<<��I��Y��kϣ_$
���%�s�Q�ȓ|��ZE-
1!>�K� 9Q�i��E�������&��Kц\�tҐ�ȓ	�p!���J+ve��S�ۏ%h@��q���H��Lh (�"*�!�`̇�a��i�c�Ψ4��!	Np�����:(�"��٤���gW��d�ȓ$� �;3��+Z��DHۍ8k����LC��gc߽&���f	��/�̄ȓQ���5M�������<KTe��@+�b�׹M�X����Bl��'��1��	X*4N$(tŞ�}H���LrJ�HC�p�HY�HK�%by�ȓ��3!��+?ӆ@��A��+>v=��h�Ą{2�C����e�M�:R��ȓm.�*��D��ȕ"��JX���S��e��J��
�z�C���!���������?h2His��%N����!02z��-_񎜩W%��4�ȓFWX|8�ͼC�yb ýpT��ȓt�x�p,C
|����ա��n@�؆ȓ�4az�΄�#�&x�f[�>e�u��hq�<H��!pՠ��Q�K]\���S�? >L��/���FA�$�P��"O��2.�\\\(r�@�76��咢"Of1��&��8p�/Ş>�(Q�r"O(-jc͔��D�����+5���Y�"O�@J2� 3 ��A�R9��9�1"O]c�H�/n֕���ɒ|�0ܰ�"O��
a송<���qTʒ=)�T�"O�iѩ�"1^ꑻ���.j�ٺG"O<��J��o�R+s���ZZ6�Г"O�����v�$%��b����2"O�=�c�rБ:U��<�$Q��[�<ɖ���H(���r����@N�<���R�j��(E� o��EH�I�<���O�f��Q� \.e!�/�@���5��"����#V��z#�'���#ǥ�R��C�	�g���kTi�?K��́��b/`�DB�1��4#�S���؈�@�	^�QPo�{�B䉡o�t��L�F�\�5!^%C�	�f�M�/��01�'�(:0��>YdG�'�4p��\�^��;qAzH<��cF�l?�%��O:��o�=?�`�����>���@�+�p=af��`��aMA�-* }b6�yX�Ġ�Cڃs]Z\¤�Zq�
�0c�Â�b&;#��Y��'��y���*g�\҇��=�1�$�ø��I,rS2I�u;�lPe��J�>=xV�ҍo�tI¦C2����"D�l����*���L�I��a�4O��Y�쭁�l�x,΄��*_�M�$�>�O�PF�ǰ_�",s��:X8>%)sO�HmG�c���Z���`��ٵ���rz8{6�-`*��zqX\	��d�@�2��R�Xp��7-ӱ.ax��  ��2c�o��QY�B!xT���`�%�Hm�)� )\��Ox��eIO	�<h;���GH@�ї��|�6��z���*C�,z�<��`!�G��Q5�LdoO����'��]����%��|�W 7zk����\$!��3�I|fP��_�^B�Q*"�r�'��WL����x�Ա�aX�d�X��TD�h��_�?��H�"�Q�F�T2ew��� ��"�� qb޵��<�FA����TS����D@Z2�i�@�D�j�*�x��TXA��J:q���eȎ`O��@�^�b: ���(��E�*R:���D`M�I���')$9��i�n����ŗ=kXIZ��i�"G6����t�~	[ĎJ�$x!�Dݵ+"����J�ABhH��_�5k�u�b�+(���4K<��`3��|r��>N��9C��<"���b� �PxR#ߧ<*؄`��U��٠���`�$��c`�I �9����h�鉶S#�A��J�QJsrψ}2���U�&�� �^$�t�FJ�8@x���cgZ�;������_��t��ȓx���N\,htp�DM�iN��&���0�#זp��#�3�ލG���E�D��Bj_�y�����I��yb��d����kP�~��Ŋ"E�D6=`�J^��	4+t)��O�7E�^L"�IG#J=�� a"O촛w(?�␊��,{nFU���x�V���K��y8a|"b��@���b��Z�[Re'��=y�<%T��F�
��0́0�X����u����ȓ+��@���?�Bq��E������ȓ'��(���!	cdD?!F.H����#H�`.�1�i�^x��ȓr�"q�G �@ u�n7���t���r���eCg�Q�`�ȓf��t3c#��W:��OH�FC�Ɇ"��@U-�A<�=�e@	G�C�	�o�"dw��}���*��]~s\C�ɴk!B�A2�]8���C�߾n)�B��+�Mb�/�`B�5_q�B�!o�	�KC��ZqB$W%�B�2c�X��CjK��T�X�C��XC�I#
[�06�yz4릧�9e�C��$� �B�V�(�Xa^~��B�)� f��Um�
�|��a�<\F� "O�I����Cf����
pTQ�U"O�ɒ�Մ4
 �6k	1/�1P"O�yxp�K:�\����T(@�"OL�R89̊@��*p��Dcu"Ozu ��P�ݺ��G&R����A"O��5A�l�����χ!�dS�"O�lpt�ȴR�8����<{�uAD"O����A�9����0�Oh���t"Oz�z��$�fE���${d�(�e"O�=�tbP�9D20�a�9Qrh�&"OJ�����_Z<T�kM�C\�1g"OV4�a��,x\NIӣ�YgL�\)"O��$H�,CE��P�j�v~�@�"O�i��1nl�(�éB�Yɂ�iT"O��j�� "Fȸ�*��&oH�!"O�P�CA�*��5q *ۻJ[�{�"O9	�`�S���0h�REI��"O�0�D*D�O��@')��Q���;U"O
{Qo��F��w�A06�hw"OH�nĿ6vL�`&�ad�:�)9D� ���кD��[Q�ɰx��0��6D�@�s�A���%�P-_��`��b#D�����)<˖�j� '�DSæ#D�8���P�]����UD��Ͷ0S��<D�Dx� Ŕ�9�1�L�'��,��C8D�̺�X�/0H�w
�'td�a9D��RS��ht=�w�ԟL�,T���4D�����Ք9�VX��:tTB�K'�3D����dƫ40\i�I�<�05�3D�0#��;ܸ=I��D�a���` .D�h��Y*����F�b.��2ea2D�$�D.T�f�dC���T���f.D���ceW�P�ve���0���q�!D����([�?�DɛCiǤbrA��C(D��'IL���)���Bz�03D���R���z
m�O�<|��Yr�1D�ā�N�'��p��̄b��!�u.*D�#��Tr̆�3�*C�PKԝQ�/D�Sq��7�V��n��	 ��y��(D�8y�)��L�NaJH�y�i�Ū*4�`�T�G�b��8��e˙R�PXˣb֌N�x|8V,/�O�s#:^"�(�U�@s�����'�B�qd+ 5��	��8ڕ�pd��r��&(���Kw�!:�G�?'TΩZ�F��!����O��s���xE��e�O� l6�W,`�$�e���
�C�'�
M8�ʋ����6��p~ 	pDHP�q���hܸ��s�@b�g̓P� u�T���]d�"��Q�����IQ�i�Q�H���� -V%�.$�TdǕ��b�+�`��d������5m[�0R<A���A�]-џ\�G'׶h�d��嚯�t���`	G���Q��`��S�B��<�}�Sc�O��Ð�~����<7�`j�Ċ3K<ɲ��\=	�?9S��ߚx�h\�N¸\!�9��y�<��h ��-ڮ��p-ݞL�4\�"H�)���m����ɑ��v��	�&&���n�4ڍ0f ��,�����X��`�gf�M7�#����s�M�'s��`�c
�u�Jh��~8��qT� #�8�r��:�Z��4�?U����H�-H�)��
s��#e�?9���@J5�&G>.y2 �)D��if� \i��d����+V�D�d��(�Ƌ~Hd�p��=g�B�IF�ɼ�b���F���z��K0i�R#ѥ�F�<	��@+Ij�v�Ûh�$u�M�&����mL*��f)�^����Ld�<��lܭp+P�T�ҚU����`YV���y1��}�Q�̝.'��i`�*��1U#��f�B�A ���M1�O��d�&6�tM	椝���5(��d�=n�@1��S���8���Yp�p���?� b�+�`�h�Bݸ���Wt<iل"O��rU��8j�.��aєW�nC��+S\̹�Vyq�OG2qk��b��$lۼ�5�O.`!b�R���+
^��s�g�C�<��KY�o������Q�>86�R`�^�:����<� �s�������+!l���<	���@���裂G��\ڇ�}�����"�,4���C�ϝ%I���F��_�0�pp@��v@�n�k� �����p>��@�y� �б��8/b
� ��C�0h���B��u��Ԡ�`�IIà�)l"�	�$z@�����B��m2eB�%�!��cԸ��@G���9A�L�U��h�mڣInx2��X�a��;�`،��O�^!�;4 �)��f@x�|Qy��T�5Z\��ȓ
Kpթ��=�~�S�#��0!F��dWk�: ��IV>c6�C�B��
Ix͑F�#�5�.���@]�+���X3��d�~؇�	0i5���I�:��t�E� ��LQ
\��j�)N�}it�[����I6�1Y���o�b�f�;9���4k�(]�K�(���� v�XH3�P25���G���!Gq����Ō&��C�	����(cl��5ڢ���HM wp��{
�1���bí��+��jg8�'9��Z�H�Y�m�<{X�,"�0}�!�U�U]B��p��F�ݳ����T�P�E�1�{d�<	�,E�`�ϨO�Ԉ6'���rJ�C޿lɰ�s�'��ik�E��iIlH�c�R>o�r�S�9��ɰ�y�a�S�lmqal�+e���"�@C��(O6Pk�!��R�niE��E�?l%��u%N�^-V�Xֈ��y��L�6�<$s�Ǫy���FF�yRm�d�~Y��ဟ,���ȁJX6�y�/�4h�6� 1# XKLP��y�g��l�.8�C�S�k
r�P�5�yB�K� 	YB��v�Fi���M�yr��O�hmi�%�k�v�W�<�y�.;�b�jt%��h�D$2'�\�y��D'�Q�#ʈo��4�ŉ	�y�+C(h-T�sB�)Z����5l�y2�0F
�Y'L�e��{U'�9�y��SN@��#T�T�)�N���yBOܸYպS�:Q���&ף�y­6��H:��<<*��;�[��y�h�=7���F�]�(pT(�`�A�yBY-��b��#���Z0b�(�y.�]�D�j���$�i���y��?)�F��`� 	�`l��+�y"�Ĉ�6����K�!�1.��y2�@�6��9��I�}��l�D���y�e4NR0��π?sB���/ώ�yR���@�ۢ⋕K�ʆ�^'�y���J����
��˕B�y��/���K7.�0�8��
_��yr�Ku�&�1E�ֶw�)�"��yB��-<���EIЎ@����U.�y�@	z�Ҝ˶EA7�$I�g��>�y⍎.5�a+t!$�y��\��y��śr�xK!l[��`�Y��y��׼;�f9U�7'Qz8�FA��y�C��[ L|!�$w@����V��y��T.i��qkD��
�e�H͝�yRDC9N�@ �l�xN���bܺ�y��^S�Ԃ�����|������y��E1�͙�l
5�J}��B��y��G	>���._�0�����݆�y�Z�F_�1���T.]�mqW�yB�ܞX*�$�`bJБV�ޣ�yR��m���4����i4�yBg
7)�MA�I	�6x�vU��y�܅rf �Ӳc���p�$���y��F�xBT�Á���j�xi�4a�3�yr�@�By"R�7uJ���,���y
� f�"�ĉ\��X���d��P"O`��׮P!)D2B�B����x�V"O )����g��ɒᄜTΆE @"O�JD-�3���GB�*+��$�"O���@�H,pҖ"֯�6��"O.�q�3C�b�2AaيZtr)��"O�T�rg��/r(=$FD:a}��Ɇ"O�H�1gF�V+:-S�&�`�j1�'"O��I6���;�0�6�Ͽ�t�zE"Oj��u�
2N������ʒD����yB�]3Q�J-�W�?��\�B��-�y��OtH�bZ4�J�e���y�0��4h�B<��ȳ͇��y��Y�s� ���!�|J�9Q��߉�y���o���q'OW�sw0��e�7�y�E�:+�jT���_�[��8�"�1�yIH#����bSx|��F՜�y�W� ���U4s��C��y�KX�KT�ö�"x������y"Cϔ>����5�ƀp�����Ո�y��ڷ1�h�s���!h��xc���y2��Rz^��4j�:�)
1N܋�y�/�f�2mZ����o����e��3�yR��3���#m<f�0B�폻�yr� �'պ-8�n��S	�)�P���yr�>�tek�ܖT|"�Y- �y��h�4�ycm�*�fԙ1���y���:��M��N��fZJ؎���S�t�B�ش@R�f�ˋ@:4��ȓsJ�����F�b��/��s�4 �ȓ&�=S�g�^Ѐ4�4L��ȓ	e@q���@�x0�0k�D��ȓ�l5S���2��Y�P�N�{����ȓ?�Z��4Ɖ ^*^=8g�/i}p���}p(r�C�9��`���Ϡ�"=�ȓPR���c�0da�X#��%6����^�P 
�M��r@f�:� �q2�y�ȓV��M��O����CG�N��`��դ	��hG
|B�LR%��T��z��#�G�,��@�ώ?~���#�z�ZD,@%��(���8'O�1��	�0�'cU	���!��1jP�ȓ0�ֽJ��W7��dY��\純�ȓH�l���}�8��U&P������`�Zv�X&��d��@P�rUD��ȓ0%�I؛�"T
��p��L�ȓUp��o�2e�n�)�)S��fهȓ�ɫ�B�b2]1�"��w����ȓk�}YWC,zD&�h�lԗ8���ȓ��ѥA����] ֮Fy��ȓ*� ��GI���,�c�F�q�*��ȓ�F��n�jO� Zg��,V��9��E��'F���n��NV�݅�5������¹XA��B
�a�ش��nb�y��Y�;	����A
{N���k���Q�Փ
s���O� I�ńȓ|�D�����K�f�;��a��I����-��]�B�˦ʔ@ L��ȓGff��ȍ#�����(k.$��_��(&�_{F�䇓+��P��}y2��D1?$ {��n.D�ȓ]C` �
�l%�a��+U+�M�ȓb�
�3%ʘ�)�I��X�4��n���CD5%X�Y0q��u�&h��S�? �-Bs�׭]�z�HdF�����Q"O(��#� y�Ɲ��îk��	��"O`�1#�5�|�*����i�:(�"O0M�3
�,51� e�%IH��b"ODR��א~�V鲒
�2�ܫd"O�|¥�E�)`xI
BOP��"O��x3Q�ͤ�ci��L'���"O~T�d�jQp�hJ��c"OL�B���c<��*q��!X�p �"O���@H�nLPB�Q�u6��"O�*�[ m�n�0��:#)���"ON �ȣ3������t����"O��BUjE�k㐔+������"O䁙�E�u��]PB�2>��m��"On@cto] ip�ѡ�M�7H�0-�f"O�ʠ�|<\k���-�����"O�P(��1~��O�i����"O^u�,��i;�Ͳ��[�W�� r"O&y���6{�,��8k�ļ��"O(��bE9�`9��'o8`�"O�YJ��W6�`2��ӡ|���V"O�e�D�ΨWN���!FZ�l��əs��7+��a*ȑW1�tsaMѳ>|0�ɰN�h�&o�:1��ę�n9T&�Dʆi��,���: ��H��
�<Ld@�V��?y.=���t��D�O^,���b?�+d�6M@�Xw�D>q�6A�$��9B�rih�O>i��i^s���S	����U4TX�P���^��q�H�����I�,�^�H<�}2QN2L��9JܔO[0�I$��ly�P�qR<iɀ1}r�!_�� �c]�b�\xR�
�7A�6M�:�x��D��S�0
� b�o3la!���;*����d�ںGx��ƱH6.H�b��1+vj�ozxT� ��۞�2O�3��|�'l�0��u��l٤�]61�@��'ݞ����}��O�>�@j�+
�h�c@�CR������ɸ�:ҧ�'8��O:8x�eʜ�4��)�VΛ'��H��i�N���ƕ�%���	;H>uϧ_x��aQ�_͎�Q�E<vԌ�q�E�.���̈��M�׮�\2���S aH�RザF4�B��=<�F F����M�ƨ��U������Ḩ��ߟ��ׂ\�N9�0�'�2�"�w@�কc�	Ǟ&Q� �'a��I[�TBb0�tc�8V�����LL���B5F#I6���g���d�?Q��C&�p�H2��&��z%�T��cHB�.$�|�i>�����Nx���Y��!���/`~��>���KX>5�v'P���Q�OM2g��M�@�6��3B�$`DxJ|��j��e;`�z��ٖ@�����g�	3-�"<�~�r��1\*�A,6GU�бz�	�:����<|W���Z2t��Ya��?�(6�ʴbu�"���i��a�b�GEx�`�猶:.Q�l�ᓸM��u�o�yV� �Ŭ��~C�I�X�"a���*�z�#G��HC�	9#.<XD�Y k2v��!��V�C�	G��@¬F�izF����A�g�C�	3�2��$��kfx}�b�+HB�ɠ`��	��׮�m'�	��hB�ɐ.1F�t*
�{)H0��G�u�XB�-Yfya�T,��u��!�d�;�>͉���q{2YA���WG!��W�b��<y�B	$Ӕe)ԯ�#0!�$G�M�ѳ��H�%��� ���4!�dT&I]:���P9�hI>Sq!����8�ṠӃp��]�(�/�Py"�O��&�sQ��3L�j�`����y m�p�"l�=qP��ҤE��y2���v۴�z���>�Ur��� �Py�J�+$Ɂ��O�cŦ��'J�M�<�g��[LV`x�"ْC)���J�`�<� �
�K�����J�O; �Ƞ@�Z�<�R��,
4�B��IZPr�UDV�<� U�v�.�r0[��_�D�)�%"O��Aƀ=s�m���ϒ3}�1��"O�t`��\:b�#�LZ+p��4"O�U��OX!4�z5@ኔ-L�)*E"O�,�u�5A��*�#�MI�"OB������A��i�>-��\
 "Od�ss,'!��h ��[�����"O�ta�ҙ��5�B)M�K��B"O�q	���/:'$�B�M"�pA�"Of�2pbS�4�6Sfm�/�t���"O:(�eO>u�����ڟoȴ� "O����@�*�0P�R�Z\�i�"O<��1�K;�N4y����HQ�LHb"O��Q�S+2��T�X'c�> 8�"Ohq�e��.\���+�s	:U�"O�p��L��R- �3t�A�<�4�K1"O�́�-�]n̸;���0Ǌ�H�"O��0Q�Wʶ|a�dW=c�v�9�"Oh����$!#�ʄ-n�z��q"Op�R�n�.
&��ɡW4:����`"O����btlظ���� ��	s�"O�� {t����ۛ2��i �"O�x��ҥ\
"�D�7<$	 "O2(W"V�,DQ���Kz��"O@�cvHM��	#��ħ\�N�Zf"O���t�;H�F��G�#j��$"O�U	L�z��@L���KP"Or�C�o	�*�`���6A�}hf"O|�{��:K9�t�G��*l!bPe"On�`�E�y$�|₌4[��Dڡ"OްB�.�L8��Al˪2R�U�"O�P�E��5��x�"VI����"Op�*$e�v�0��u�[�S=����"O���i��M�-���p,�q#�"O�A�&/]&J�p��3Hʕ|!y�"Ot؂ԂÅl���sA_��� r�"OHP��	�(Mh$AJ���P9p�I$"O,���'��T��҇J^3h8��;f"O�5�@�CV���;D*���"O�%�`b�67��@�bI��l�u�"O���V'�j"�x:���	�P��"Oh��F�#D?���f�-|@ɢ�"O4�bg�4DR��0�G
Q^���4"Od̑���v�)��ɘB�N��7"O)���`�0X�e䑤t���Xc"O�@	�艖LR453�(^�`��M#v"O�a���L]�j9"�,f��$k"O�X	!L̐Am]3r�U@�"OND뀥�j(�� +�9��z�"O@�ȓ�E@�(�s
N8nMD�0�"O��P��+J�,�/�;��؋"O�����/1^��`�L_����"O� �%���R��$����"O��3��\ ��,C�#�Z�:A"O�AS����{7�4������@&"O�l{T�3�`U�k� |`(���"O��4 I�w7���ˈb2�j""O�Hr����%pJ��q	�G�J1�P"O��k�$�vĘBh�Q7z��"O���VJ�8Ey�<
��F�*�\�"O��.��y����r�_�S�xJ�"OrHy"c��	x(dJ�����Е"OT0�tK� k�r &Y���[C"O �Z���rm��EK�|Y�"O� ��qr	̩��A�Ŭ�:d��q��"O Xq�f�t�YH�DC�fĠ@"O���#H�pG��v��7�:�Y�"O��X�c.�9��b��h�h�҂"O ,�Ҥ�+/̖-��]�S&L|{�"O�l �aЅt�D(f�a��3"OHY���E�LE<pA邪<���1"O���5b=&�nЁ%��^���G"O�!�7��/WoByA��	���"OR��"��}��i��J�+����`"O��x5��	I����#H�O�L��B"OX�;5�+'S@���dE�p�.���"O�u��Ńy5޼�!S03�d�"O`M �@G�=��qr�^�"O�A%���$q�O�{yʍ�s"O�5�!h8���҅�˩"�\���"O�@s��$�J��Ra�� �w"O@ف�fҝi��J����� q�"O��iքf����5�Ϸ.N�}��<D����� �P�q&Hѧ{�VI�Չ D�HaB��,\���"��]�1-#D���իJ5Ztb�8u�:��đD�"D�[��KF �g]6D���TL6D��{��U�_�@-�e�NUx)���!D�� �� $vI���Q�03~��A&!D��b����q,ˈd
0���3D�|���:�xE3Q�	���5�+D��KPN����� ���r��YX�)D�Ȣ�N�	�D@@fŌ>�d\�!�(D���a��|4��ђ�r͜���,D��;��V36l"�RvNJx�t����-D�+'a��lj��zc
J�Q�\8�ׄ)D��X�#]�_ANi�gƺ�H(2��(D��X�J�[�4XHႍO^�/X�C�I�f�!b�#�NٹQ@D;}gjC䉙e������9���c4)U�6DC�	�A.�$���(|����g�s(C�	G�"�@�] &F��2cݰZڶB䉟�x�2f�$ Xt�S��d��B�ɍ:��xFd��{�"l���b�xB�ɜa��qc ӣvT��`�J+4B�/[~�}� *V�q Rx�WL��l"B�	-K��2�&^�	Cl��W+�B�	OjL�3�	#��զ�F4�B�'xBE����,����6��;��B�I~F�1�B�J`&<���G�АB�0Z�)@%��,���C�F"D�VB�	�?�2��Âe~�EaE�?V2B�Ɂo�q2�N� ��C�KúgZPB�5J��ze.�������*A�dC��u-�͙�e�.OU��P��=ZC䉹okdh�ɬJ��dK�#	�p��B�)@L��G�S�V��: b�Y��B䉠[���� .���j@�~�JC��/����(�;`h�"�e
;!K�C��/`.{��:�8�g��E��C�	 w�T��ך^P줠�ƅ�>Q�B�	sڴ9gϙe��th���0I+NC�	�Nd�i�LǮl����W49LC�	�"V���nS�J�����9BDC䉾w����@)����y�DL�C�I�U!L�G��h�b]����l(�B��1u���X���69�"DfH�.3C�I�$�d����/O6���F�~H�C�)� 6`h��O!1��ňE=#"OI��o޾80h��T�϶I����"Ov�q�O��.� dA2̆ N�"O"��W!��#=����J^����"O)сȕl�H��
�,���"O�@����-��hعYvf)�q"O:y��(_�k��9yHėgBܢ5"O�]�� �,�XY �ُ-����"OڐC�@� Ek��a��<{U"O챉F_�-�����X�Z��"O0A&�W�Q�$4��Q�:�zj"O� Ζ-2�R��G�\���"OR���%��W��}I�-M�;ߘ�0t"O�S�A7��
w�^� ���'"O��Y�~2�t�O)��q"Oh�0ëO/�D�A���L�\h�"O ya(LV���)ܶ/�J�r�"O�E��oӜ�dܨ�-8�*�!"O�Ui�-��C*δ7R�a�D"O�����"��!��I�8G�ɱW"O �(�$�(Y-n�pT�P�
��e��"O\��u��!�2� �HO"C��=ؠ"O��)qf%^������](Yx�R"O�<���ÑM������gT��"Od�ٗlӂ(�R�QL��h=t|��"O�ܙ����@��d�I%'1��@"Oh���,�aӢ�>}��� "O�̓%�F�)ZD�c�M�D��0!�"O���R��"L�u��%қFY8"OD<��B��`�>�p�KK�=�"Ozl�Č�{8`���*6�� "O��pqꉮo�p3�kV�>��͊G"O~ 2i
� ��� %��,����'"O�M��5B|���3i��H���ȥ"O�9�L��Y��M��h.'��ڑ"O���ֹe�&u��AA9+7�a��"O��I��!R:�ȁIj�4��"O*1����]A�@��a�����"O�4�s��ku��B'U��\+p"OƁ��~f0M��H:B�ܰ�P"O�$9���lPL�c��ϓ+��A�"O�e{��?����#����"O�K�j���Ǧ�;���rf"OP0pt�j���4�҉L�8-A'"O&Hs�CO�O�|�	�h_x�p�@1"O䨢�.�P�X��pmM�a� p�"O�i:AoE�g��c�k۵Vt@@�"O�9B��҅� ��Dʄ ��"O��a��P0|�R�	 �?��Ƞ�"O��{�c^�PD�)"�IL�_�{�"O�q�T�Y`´�H��,Ԁ�"O�S  
  ��   a  ;  J#  �-  |8  �C  JO  7[  Ag  us  �  ��  ��  ��  J�  �  ��  f�  R�  H�  ��  ��  �  \�  ��  ��  9�  | � 8 � � % �+ _2 �8 
? NE �K MR �X �^ <e �k �q {x A� �� ΍ � �� �� O� �� E�  `� u�	����Zv)A�'ld\�0BFz+��D��X�2T8���
#Ĵ�g޵�?Y6�S��?� ��g+(9���!���3d�����"̓G�yC�m��:q��������H[��	�iqT��%q%���d/ڇ_I��H�*ԩ9�(�2doU�Q�� � �[t�5#�)T�[0��;k\ћ�'S̛V*!W"�I���V�d}�cK�j0� j�.>���8!�>�����<q_.�n�CR�t��������Ir����s�K1K�&9�4��/�R�� �V�A�D�Sc��6|����?y��K�<y�SޟL�	�"��@s��� D�UAt�.;v����T��ԟ��I����
�&PA����8v�0
Bˌ�	�����~�t;d��af!�/I�<�gP��1D�$D�Oָ�#���t�aHġS=����	����y��dġS��]�=�x�	W�ڈy�h�F��D	ջU�����ئe���h���D��ϟ��O��Z�yz�D<E�����^�-�R�t�yl���Ms�i��Ft��i#���9hf抬#�!psň�ː͓  g�$T#�]����Aß�p���O`��r�e���`�X��pm̔�ug����Fo13�nL�
�1(�� ��޺gdFTX�ㆠg!\�h���o�M���X�I>t��6͐�����,�.1�x�2�� O7�U����h%oP�����!�Mc�/X�DIڴy5���p�j���o�Aw���oM��s�c�?@L�!'��*�mZ
�M�ÿiƀts@�T��k��{��b�T�1�*q������d�fLÑ<3H3�R5{B�d˱�h�`l��M�v��>YGf�hed6?D�D�Ę]Y�|zqk\6�ܢ��1k�ԡ��i�n��Cφ=]�b�K4iM4<�����'��OV��6��52�Ȣ��x���^n0�(�#�O����O,�	�^�huFؼ�xA��OTl��HI,BA�,2(�QA� A"�O��$WT�����O�ɹp(��8��	 k$2<���ߵP���"8Ѡ�ɍ'��E�v�<O�9���M~n�층��6���V�q��s���>��Rs�H�d�axR���oy���!#�M+v]6 ��� �?���?�H>i��?y)On�d�5�� �!g^i�٣��ݺ)�(�$�O~k���uUԓO��Ɂæ�Ӻ�?�w�9|�8� ��\J�P�c���埬�'ٰE:�y�4��<��漃�l7f��YeL�!_^l���A�����|��#ɾְ�L���M{���˛T~��!� �=�ԄI,Q���I�c
)�䕻NRb��mï��1����^ӎ�i�,:P*��e	�'��d� xR�r�|F��:��}� h�E3PE@�F��F�hș��'��O|�D�ƫ6g0�B��*�������hO��	ܦ�H�4�?��i���SV8|�FdI��ca7���'��I&	���֟p�Iʟ �'W�YI�g���؋� ��[˲%��vݹ#�<�r��\6VY��+����?Qw�̒U{LL�gB� Ɏa��#�O_��FA�>ME����,�/ZU>��|��xR�4]6���Hv��1���7&��ɶ<�cd�ҟ�\�L>I�m�.�H	"!T�@�H��↋4�?������O��?�'R��"�Թ�Sf�2q� j���?�e�i�&6�?�4�����<)6��J�����&87���+�g�dptP���	ԟ|�'��S�|ڒ��8	VTUa��0���+�=F~�#BU�_�Yp����<���[t�{���,4d� 2#�/�*�z ۡtT��AAےEEˋ�$̀l�&jЄ(=��0WB�;u�>���'�P7M�H�'��O��'A#h�@���@�����b�O���O�=y�y2bΜ*�͋BíP���iBH޳��/���x� ˓�Pҹi�2�'M��1&`H�r��,�҇T#�r�ѓ�'��*q��'(2�@&B"XY��^�ڪ��pd���1�m	7��h�!Ft�L�&�' j xF$~JǂW,Q�U�� +�$S��ڒ(��=�fÅ+&�r�G}��J��?)�i�7��O�Tc1!U�4r���?v&�l˱�<���?����0|��N�����dHD-Ie�@h���?1��I�������Q�<^2ݢ�H�B ��AO���M���#����ܐP,l6M�Ovʓ���'�?�AGS9@�D�c���"Ą�u��+�?	��.��� AF��iΦ��4F�B7�+��+kH4zqʊ�6�����o3c���'"�=���2Q`��^��̎�Ѹ	�$�3bi����J�x�n��:[j`0�Qb��;?����8�4��O1�2�eBh���P��;V)�� ԗ|r�'�'�"�'>剶 �x��"�8H9q��U랈���Op����Y�	��M��6K�T ~�&��uHP��GCY��M���?��d��ڇm���?Y��?����y'ϔ
]�"}J��M��1XmY4?��)�7�<.��c�#0��m��Q>!H���V>�6y1��(�>��&J�)"X�e��mG�#V�m*�ӫU���*�E&7���+u�V	ҥ�d��(ި6;踃DLG�\��§�צ%k�V���Q��OBb>�$�O��dU+9S:9�$n�/?:h�� R).�����OR�D�O6��.�3}ҭ­(H���A ~�Z8�cČ�?��l�F�}�������a���?���N��G�R�z�C1�Z�h4*�B�?&|و�hU��r�'b�'��$�'�"6��e)W�ȽC��(j�-�3L �#�ȜPd:J��%�ʜ�gH�KPPD~��޴d}����o�P| ��
�D��cH:]���1��4M�I�h�$�`�i���O*�`�˓�^Tz��5� -W�qt�ަh�"�'�ўTFx@G�`��� h�6Q��uAf���=�yB�!̀P��㓗"HdP�a�I)��]����'���C�&��ݴ�?��27�!��8��P(��ΉA.:@���?���F��?q���?�6ˆ���dhFH����{�? �m�Aʊo/4��r�
`� ���'��B��Ҏ[=��ip�E�_�D��G"P)��Pc���qM2��G(ԆSW�c�)I���=���͟(p�4<��I&���ui3���ێx
ЃL���e�'M։cW�\[�Ll�D̌OFPm�>v�ƪ��(��"A�I�0�=R�SN�6�<���0N����'�[>1w�П�H���L�����\X�
6�[̟(�	=u�z�Fc��S#(Uaca�L��.�
�,/`�I�`V,#�D��BP�P`��'����G�(1ǀ��#1�����3}��k�B�%?��n[�1���aÞ�$�jP�X��$F=K��'��>����d�֙�p��dA<ȓ�FѺ{�ȵ��F2���Ɔ-lEXMA�;Au��F{R�'X"=�dO�Hℤ�֥Ӎ+�|i2�)ۺ�?����?��8����e�?����?���y�i	�fzD����	:R�`��*�1��X�e�Y�^j��~Þ�ˋ��" ��G$tb=1��#$�������,��b�����#ь��ʈ�P�I�5��'Q�AA��yG₞ZJ4,@�`NwX����O��?�O$�R��'kr�I-giz�B���*B���	Id��i�8YR��'i� ���tHpM�	䟄i��4��D�<Y��YO�\+� CJ.!�Š' i,�XFm���?���?���O��O
��~>�����6t*S��O�x�f!	�D�1V">�@E�)EY����_�g)�x��I���Pb��.��5�<3!��P�/8>C�y��h��x"�L���?�MS X/E�j���:;P�1!`����l�	E�'�̨Bő~�<U
�O� d�B�HP�"D��t�׫0���'�ݑ�RL��/.�D�IHy���,��'�?�A�}h�(v͔8�9����?Y��g�����?��O86�����3N�B!��x��iT��<8�Й�F�x�T�q��U=:�Ei��F�'��� �K:O���V*X5ur��C�2%E(<�V$��n��a�MYeT����bOH�'+�����B��F�<�㏛�\�&M�-
E����v�Ii�hт/W�T��)R�Yz���=��n���$�O���3�Z ^�$ɗ홢d�vݫu�'1����]��4�?�����)R�C���dN�0%Pщ��"ߎ�k�Ә[Ԙ���O��P��U�A��$)W�N�Y���ԙ?@�$t�{I�4I� +?��J��rգ�I�5D�Ѩ�(�T���б���ۋw������݀C���ד�Щ��O<�d5ڧ�y�*n$%���K7&�.Ecӧ��ybE͎`Pp1(B�Q1I�UC��+��O|�F�de�6</�%ҵ�B=�p0���́.W�V�'���&���ݟ���Ɵh�'y�H��IX^�Q��ȟ.<1Ч��<e���A�3��I��$�S�?i�`!M+L�ɓY�F��p��r����a��!Oc(�	��I%x�@���Mc�I�>�$E	,��d�Ee�����p�~�@S.�4)�jp�Ɇ&� �nڡ��$�5H:��O��3��W�RU0��f�5���U
��3 ��<����?���	����蒣��?F���%���2���OX�lZ��MK����vV>a�M��(��B���AŚ�+��yf	a���(��uӲ�D�O��d�<�|�4`K�0E��	Ɗ�}۴|���?	�
Љ7D�W�Ipt��?r>)"#kM�B*:dEy�GN�ctyc±\�C0#M�=�F�$�<� �H��O�_�����{l�
C��=>L"K>1s͟ }Xʗ���q�EY�N�Xaqk�O؜o#�HO>#<����WD�JS��,}f�q+`Bs����<y��&�l��HS��
�A&�h�+�MK�����x�`}o�؟��ɮx ���M�<��:1 [�ň��	��`i ��l���|��ϟ��<	ɉ�>��r"ǦF� !�'|��8�4��xqW�
AW~x��զzz ��I�xxZ���S�ɸT
���8d��-���̋lpB�	���H2��=5��IjuJ
? ���d��� pf�U�x��} �,�kQP���D1�DV,;H�mz>u��r�D��#���ra\P�W�HN��q�a�"��'e,�p7m
ww��a�+[Hh��o�|�ȟ��	�B?��=�����Jp��<b��?	���dZU��!ܴ��O�"I"��
�p�l0i0�͋Vb���On�`��'�b��՟�9�`W��*G+ҸZY\Dz�GM�<b�Z ��嚅(�{���ƂWG�'��>ғ@�x�z�l���(U��K��@æM���?	��?Ac�	8Q������?���?1�wlL�i���;�ǁ�8�r��@
\&���eM
xN�r����O �OU�ceA�7/"��w�G�9��w�\-#�Dyr�NK� $"�S�Ɲ[H?�q5J�"�=�&!���C�#R� �'��A5�����'����>�,�$�O�=q�`�a.E-����W�BZx *�'Te(�P�hV�2H>T}d`�-O\�Fz�O�R[����k�;�q��I��ݢP/�)<HX�ԇ^ğ�������ɘ�u��'.�9�V���`H;b)>��$DNM���uoD�V���Sd$�g"�|��A� e��6ߋ@�Q��g)%� DL1JJ�JV>|��F<i�`x�w��6̎��dC�z�2�k�8�7��N�r�%�$�7��_\���@OіT�8h"k'^�����O��� ��P�OW��#��T*p�dBGI�7mCDȚ
��'�x͊r��6)�䤉���>b�\M>q�i��[��áʋ�����O"$�`_�3�tx���
�R��b���O��Đ�����O�S���L��B��@���K�֊!E��J0 ܧM��I)�"M�Sς	a�剄!_`$;3�Q�]��H�`�f�n�A$�^U�1���ۑ~�QFJ#!�ș��Ih;���PѦ�"(OthIU �*�\���J�VŒm��|��'��bc�Γw�҅zD#4	Z�c��F�B�F�h"!(�DX����,�?�+On����Oj��O��'��*�;ȹ�E�Aټ��#/�p�XQ����?��(��Qx���SW9�Ec}�r�x��ɭl��hYE�	�,�|m�F�����|0�A��K�>�z���[ ���`d�۶t�*�B�Oc)X!0C6�Y��h�886)��ObԳ��'�B��<9���.L8�AsȈ�O=�QIS��Y�<A����^�.���hJ�pZx�T�^�'i��}���&p��P��
�G��c`/IП������̓o�*T`���	��IԼK�aT��$���^쎤��f��7<�� ",E Dn�m���|j7h ;V�	�,���V�A	_�*�P�ɏ�@��و�Ɔ^� �&���� �hЈ"MbT�Oaʠ��ݸ�yg�?�(�j �����X6�C-�?A�O^����'�퉟{�`��3��h "ăf�-g�2	�ȓW4z��ë�2��飫�+#�������ڌ�4���D�<�vH�o����� 'vO��I ���nC0u�3/��?A��?i�`��.�OD��f>��T�(�r'kN	�X���ɶ7f��bc4g�$����	8D�F����#�hBn	f͊�B��˳'"jL������x��3D�X���<#�mis��U�ᶬq��'���S�D� ިA(�HW���
��>5|���C�y���@+�g{Ft����t
}�hm4���,-\$���۴��\1t-2�W?���bEZ�KBnÌV�8ě@k�>
1������%.��@�	�|ʰ�j�b8�C�T�xJ�E"ȡg�@�T�Z,�pc�	#B�����0-���8�b��h^��p!N1oLZ|X�'ِ:�J2G"N"!�N) A�C��O��qg�'���9a��-���BRb��?�0%ZG4�$!�Ob�(���&-�����I/R�ܡ���'Ԝ���$#���p���PI���;B"Ҝ�����OF�$�O�ʧUy>%���I0�Sah�4a��4J4+���R����?��lG>p��9
s(A4\L�0N��]�f4��0��i_(@�z�����NU2A�`$B��	�R�x���M7X�]j��EZ`�i�)�� #W��?�1Áp'�Dyv-b<�d�$9?����Ɵd��W�O��dS�l�M����z���ʉ4K�!�DL�L�C�e��e�r��1IW�<ў�����HO��:S�̋lf�FDQ��Ś���O����O��$Q� �f�����O�D�O2��nޙ�0%�(<����D�O��4CqH�X<�p˓�~�.L��ʲ�
b>��i�(#��d	�&�:5��e@;k�F�jvE�	�Z�[ ,^�]�0�E�è\J�I��.��˧9�r���C����0ra&V�`�f���],<xb���
'��O��D&�zB��%bÝR��f���=8��y�'90��7z&h���"R).��x���?Y��i>��IPyb��+wmP���T"�� +�[�.�B���L"�'F��'}���'�b2��|IG��8.tGOը��$!E��N����q%NR��=�1	 
d9X�F~2 P����>
j���S*stn�:�`�
2X�=c@D�:^�{�
�zxfa���oܓ?���'�	(G��y��1f�l3D�����x�'���f�*Z�&e�c�U�woҽ8�1D�p�f
�D�%#��`6�	���0�dN즩��fyˍ�|cb��?	����w.~��N�u(�0�㞹�?����4����?ٜO~�,���N&JN�$e��i�z�0dd�[Q�4`�(�n��<d�	E(�#?	�#O�s7 �rt$	=}! k�h�7x�� H�\�E��g����:���y�iI�-6���=Ʉ�ޟ���{~2�S�vG��P���*��!�b�-���0>!�b)��`(���n�<@��Q������\A*'H�z�Qrq�P�Q6��Icy�KJYU��'�S>���Ο :@��?* �r���
x�|�@C������*O"�	�t�H�=(}Z��ߚK��ҟ<�4d�`��]14R�Q�6	���h�'8z��42j�xU ��$�Tbe�fݑ�Wi�A!Pi�<km40�O��,$�}�#���tUJ�\ZH|��ڟ�F�t2OXQQ�̞A��u�6�_�H��\`"Ob�r�E�X�fL2 �Us���g�	� ����V�t�X�� ����/C3g PalZ�t�Iǟ,.@~�{�	]����Οl���+�
�;� lQ�J�4�#�h��q D�p	Ƅw�,ը����5�F5�|ڃ�xb�
 ��h;���2-�JI˔f�?G����φ�G��ѭ�)xJ}���4K9�� V��$) �|0Y�Ě!�d���'�I�B����O �=�$���5*}�5/��#���ZQ#�>�y2���d=.`�+�\p��G�*��d�Q�����'m��?��CaJ�;v2]�@��j�FE�e	(֮Q��� �I����Sџ��	�|z��G#)�!9�Q�q5(�dh�z���i܉@0�q{�Ņ ->e���Ix��D��&�dO��[��H�A��Se��]+����J�c� g� ��M�7͉���0L>��I=z��r��^;
��'�Ԣ�����ʟ,F{��I�P�A3%��U��� _,���=��:<��YB�,^r�"1�N�M�@�O�tmݟ��'�H s��~���ujP�S�Y7q��}pf�?H������?�eD���?q����TnT�o)���`
�$tl�CaK�<\�L�B�V��80�B�.1������I��E�$��]HdƔ�dQ	�aܨ$@���͑qdH@�NZ�8�'�B��tsu�H>��E�s�	�3�v,�p,,�$)�O�x��@@^(�1�[�/ht� �'�f��Xk]|t�V�X?m�Z�00����P���"ɟ���ٟ�O��9P�'M&0q����^���1�-\�E���8��'�r(�Y�}YE�U�'��8TO��d�lm����	 �E�v����"�������P�I7rRLa�Fc�(Z{j�a%N���+g"_xP�-L1����IpP	���S¬��'����?����}�����$%�J0(7f5F�r���o'D�(�֬�n��[��ϔj�I�$�=;�>���Ē-��$�n�?T��ZWF\ئ���ڟ���b�$�Ѕ�ʟl��Ɵ|������\5I
]���R 6XeH�%z=�'G�ܑ!ʔ��Ϙ'�Y;$/��]�Z�(�ܙT�.�:�e�.uҌq�T�ؗ2����5mO�sh����!Z��iG��!;�#�+*��P���D��O��P��'�1�1O���� ]M��P�V-D�J���"O�l����
gc��0���/'�x�']�p��4�2�O6�ӥ+�2�4ԃ7#�x��@W��e�J}[�N�O$���OX�$�6�D�O��ӖR�@<��N�63j�  We�!K �z�B�}���2"�GF<��s�ߵ`Ex�D{��.J�:(�reխz���{Q�������oN(E�Y�w+Ʀ `�;�͔_���c�?H��'���)�}�<0;fM)/�����?I��hO�#<r˜?}v^a�1�/W��B�j�<9F�7_F8����%�bh����P��,�M�����D�%\b��Ox���!%�(OΓp�@t�v�@7kd��'�>�`��''B0�����fЌ��d$/kj@�/M<�F��7O
��l�)�!Mj����MI4�(O4�"������4A�� j����X5k�,�p&Q� ��:�&�42�+ݴ~��T�$ςs���'>�	�A�Yxe@��J�����>��OF��d�� @|C��q*�C�=(�����O~q4̓@���(&CK$k��T�Ll��Ms���?�.�n����O��R3��2o(�F-T7��`����O��$��Z���2r����430LS�"ʧ��	M�
�&#jdճ�!%�F`�Ott�-�:R%��B�@5��xˏ�D�J`��ŮR����ÍA>����~��'��>�̓&�4���:����F�s}�e�ȓ1���V�M�؜����3@~lD� $�'�.���#�~��ׯ��] ��	������c!�ʀq�4���ğ����̻���r)=��X�kP#�L����W���h�Á��A��	�f̧-�Ϡ�d�g�H�*�
� �&QM�`�t��o{L���l�R
�i�� IY�%?�lZ�t�n$�;E��BE�8�f@��3*�X(��Q~"�E��?���hO� ���"r�@]I-׃l0��B� -D�t{�`S/!��U+�xhb�a�F�<A��i>��	Jy�03�"�0F��j��<{Q�ƃ���(�ʙe��'xb�'� ם����	�|zD%	�x�"�be��=p��xz��B�Ub�E���4e�DXr�		<x�p Ơ^�x�b�<���-�p�Aq,î=���:�E]>.B��y��N�h���7 ^qzٴ&�a(��$= `�! jתK��4�Ou�PT���'|��D���U(r.I-�v�bHP?�!���*8CuavΑ�CC��g�2)�'��7�/�$A�f�X�'?�sF�<
z<	���65�B�O
ʓ�?��?� j�* �- ��I�Ah��s�'�(��gI�6}|؀�J��Np��cU� ��7g
X8ٵ�-g��T:"���Q?4 ��H��r�p�3�>�`��2)@�d�O$�E5��CM�M[P���l̯K"��&����I�FT��X�s�T<��fԌe�
㟬F{�Oz��$Ά i��Ս�1���[X��'q�9r�̖����|Z�4�ڰ ��	�.�`V!�x���?��߱5�2v�%+�Q����:�Z%��S��	��.Df�p`�d��j�ΐ�	�^y��mc�X	�Aퟭu�J|�Ԏ�#)���k�HǐQy���3�V]~�&���?����h���)� ��A�n?4)�D3���
�"O4��2	LG�X���Q�?�N9��	ğ����d0\ E���WFb$��i�!Q�,���S�(���O.�$�O�Ӻ�kٮy�4��T���<�	�$�=>�\i�ċ�ӟX��DW�xBc>c��		  U��UEAd�����C�P�Z�c�#E�\'ިp6�'��b>%9&����D߸D�����Q�b ̥Y�H�Pr���S���O���2ړJ�r��b�I�! �EI&pq�'���:����2Ğ�9�i4�԰����?Ѵ�)�+O@�U���z<p� ڌS�`�#w9&�8���O���O�ŞH�F���(��]NE�7(�
&	�	eb�C�Έ���P&K�	��'�X�U�#}}:���ȏ2:�hPGF�0�MsUiC/�����K4���IY@�'������G��q
�-����[�?����hO"<�U���h;��8!N9��@~���<ѥa�qĵr�G3z"^���ϝy򉌅�Ŀ<S��O����Ae�pq�g��L��Lh�����O0���Oh��g��1|�֔�~�Z�5�'�`q�7	�"o���-��I͘1�Óa/ִ �*\���c�T6e�\h��F>K��+B'�8�p���n�@��鉿?z��D�Ox�]���֮B�k�9H�
�#��$�4��	�]>c��X�A獼R�N⟜E{�O�6��"y*�qxB�β)��u���=�"S��8�F\yʟ�˧�?Y�!T�V��yk��xG��8iR�+���?�l�3C�2��� �-`}���������%�805����
�zR�ԡV��hڄ�ؽ(�z@��	�	I�x�'J�N�J|jS'b�8kÁߧ/�q!���~~����?q���h���9>r4a�KԿm��!aG	"��C䉼SN"a*У�9�J�8��,uU�=9�7g��D��A����Y���x���Ey"W� :gm��h��ܟ8�Idy���'7�D�l��K.b��&��>B8d�2�k��e�8�$��UkQ"u��D�M}�3��0&���� �p��aҠ����0�ȑ�?a0�s�Ј�'="a�'Q�1c���,X�x��������$��\���'Zўd��ʜz�p�hGd:�b%�M�<���՚ /��D�� �a�d�˟��I.�HO�@y"��"	Q"`s��vW!�GM�%/���O�����H,2i��J�	��'Tr�<q�'���#��B��Z�T/X�B@�
��?	F.�(�?���?��ƅT�>	��о'4 ��2iPL���gW7'h���iF��̻b�MW��Fyrdױy� ��o�6>~VL�0�A�cyf���-��.%,�+�K�o�Խ3�*ѝ;���bEܥ"�'������?I��k0C�[&䃡q�QvK����$9�O~ī1�7�>���/a)l ��|b�i>YK.O�8��L���@5)3�ŗ*&ri��W�؊���`3R"�ԟ<�Oo�����Ol��K>jj`��4k�!�8��ba�|��ܗr�h�3JO&	sd�T)G�Yz�y�'�O/����
H/0�J���iȓ�>(�'�^$K�oY'm�� 3lΈvH�i� �%ҧ:�� tj�X���u&�I��̓C����	�����ĜD����DV�1�&�2�!���^��T��%ƕ{�\Ȩ�$J(�ў	����]͞�ǢԎL�pJ�KW�R农!"C�O���љ"�,DZ��������O>�D��z��I����Į��N\�p��q�6_�8u㴨̅��xTh�.}+:�'<U�O��r����y9�A��D2�A���4�Θ�2�,�1���	~��O7�b�4��"qM�ahg���,��0?��Ύş���m�'����}��� Ɋg�Fi��Fߴ�!��� ���P�V��]v���v��7��|�����\S fi��n4Zw�Ȫ�gțGFr��u-������O��$�O�i�;�?�������(^50(#TL �S�B�6�L�8��͈]�D���ʜ_"�G2�}�Hc�DS+xk>ha�DݔLTt��EH*/喰����#=8ٸW�Y6lꑟd1�$�O�\�k
>3:F�#��^�-��Z7��Or�=Y��E,` �(�L�!�&t�U�ʋ %!�� 9xM{��ć$o��Ѳ#�*��	��Ms���P:NQ�e�O�>��a��m.xL�{&&�e��Y��'g^Ȉ2�'hR�'��(� �8�|��`�,`t�#��ͺ#B��T��ܳ�N^F��焚B�'V��`�L��Ba�R�b�^��Be�M�' �	8 ̅SBr䛲� �J�P����X�|M�4tAj��<E����we�uy"�'��q�@M@`B5!P�����|>剭P��$�45������{�ʓNn,r���?y���IȤ(����OL,�`��Q9ĩhbfK*��5��O��`�dQ�F�y�%&ǉo:P�
�fL�����	��� �kG(A�v r���v7�X�ب<��2j� ��"?���F�ćɰ��(�͂->}ޥ	�h;�y�!^��?q������$��� ~(���F�������
=�f"O��
Q�CJ�Z5Z򤟿��\Pv�	��ȟh��� ޮ
\��KA+=�,`҅�O����O�<K�G�P�D�O����O����O����تl\�(A�̈+��|�����V1˶�J��^�ӍA�K��'g�O���t�@3يB�G�>N��0���{y�	�M� >*U��O O�S���'yМ�@���M�0�Ǉnz>8��O
�-���'Aў�[ �����0���K�䖲g����J�&u:�O�;"�J|s"��[������HO���O��m���k4!���HZ�R6_�\Lh�� �,)���?����?�'�?�����f��|��ҁ�l��ƋV�Lu��vm��P{XH`u�L�N٪e��A�S���Gy�n"d����%
�D���ɓ�i���ǁ $����Y�[��i�s�;�� r�^�0��'����{
,-[+?x�����(�����hO�#>1&�%. Ę3���^쳇�Jux��Dx����c�@XC��N?LA����̦���qy��L�f6-�O�$~>Y���\+14&E;��/�`�E �O�dc��O���OpE��G61��:���48�0��&�^p�1��Or�:���18�C��S�-]Q�Ƞ#� o�\;f ��+�pJQ��]B�Z���9!�b�ǁR�=<��@MD5"HT�AlXb�4 @���b��=� �w�Q�S@>=ⴭH��$C剛,�
'�	��N��Np*�O^�=ͧc���/^�Ȉc�k�;lm��$R�X��ʓ�?���?!��?����?�̟$`8恎X��5���׫}z�4�4�Ɇ�h���P� �R�&(?2,����Cd��'א���F�d�96�9�Cd�7r���۔��$�6-�O��F�w��k�b�O����f��u��!��];z��"�0�p� ��/`��nџ��4&�ޟ�̓_�2��������&%���^�1���� E�O�퀔��?!��XP[�'����O���H��r�D�u�C):��q����?������_U��d�O�Xӓ��O�\��)9��s����yB*Ã9�(�4Ƃ�:"�$�b@�Bj���?���) �8$X?��ş������E�gޮ٠ϛ
{Tz�@���?If�Z��I �I�	'�?���[unZ�3U,aB�BT3S:� č�F���*pe���MK�'���J���?i�%��g,R���D�O��I��J�n�*[%8DQ���m ���4av�`����O��Ċ޺����yr��x�Դi�� �_mHŪ$런m� @0u� 2^�6O�=���'%�����O���N?>�Ф�δ-p���!�^
Lm�6����C�2, �4 ���O|���OV!�B@�T͂!Ye������&Vx�3er��MHTJ��1��O(��Sɦ�!�����O�&l�30� �ÑEW�	�0xQ�,D�T��S�L12��ӫ?"z�Z��i�����<����?���$�|��)NJi��әbi�8*�.^R�m쟼��͟t�I���	�ON�$�O�����?3�q	����쩐Q�l���'+B�'���']B�')B�˲b	b�A�nP
_�,۲#�Ki6�%�D�O��D%�"}����:�(��դ��n��P��k1�M������'�93ҡ`��F\��)�4c�,k��%l�wy�^�\'�̖'���"Z��)�SB3���IG$��ILyҕ|�Q���O\qۄ嘢d������9jQ"Od�r�(������m:ql$�s4"O�E�.�>'Daa�N�_�	I"OjA�To�/*��CnPÇ"O҅� �8�
��A�P�,A���v"O���\b��Q@f���z�;�	������؟�Z�+N��طĈ��}�棝�M���?i��?!��?)���?I��?��	
;�����e&h�3�rÛ&�'Y"�'��'�2�'�b�'U2��__�<Xr��S��=1K��bJ7��Od���Oh�$�O����OP���O���ɓkh䫶���*�)2���*:8�o�ϟD�������ٟ���(�	����I�|�b��p��8Z�t��[=�E�޴�?1��?���?)���?����?-�M�waU9"&<`��	x��ʀ�E!d���'I��'�2�'b�'0B�'��O�;|��U�w*\BEl@(Р('�6M�OD�D�O�D�O����O��d�O���;��k�=W��0�Y"���m�ܟX���t�Iޟd��ߟ��	������!_��0�*�:�� #P�'0{��2�4�?Y���?����?����?Y���?�f�lx��J��[ A�:¸i�R�'���'���'L��'2�'������v��ysB�h�)�%o���D�OP���OJ�$�O����O�D�OX�p���)�jT�ڔ����ڦ��I�������ş��	����˟@��Ŕ�VB5
�H��Tr���ר�M��OP�$�<A��ICp��0����)��H�C�J6M�951O��?�ߴ�yKŸa��eI�I��H�����K���6@pӸ��i}2����	��~}��'�Y�h�cv.I����.��������ŧ�
<�����4���	�7&(�腉E�N ��t�&)�`���<�H>�6�iK�G�ʀ ���7�6�
���I�0@}^�z���^G}2(n��nZ�<�(�\X��B��(#�0�l`_�L�cHM>%��`�d#?ͧ@@xe�e��yB��DP���%�/)�*)���N$��D�<��S��~�(�bdQE�3(]"P����?!"�i��Xi�O|�nZQ��|*�]s���pp)/��H# T=�?1�i�,7m�OB�2W-�#t��IWZDP����D��ٳä-ȴ�A'h6"��rh"p ў���pyr��N�o�6�k'��̽�a�TI�xp�'�l7��1Of�?Y�2D�>���nW���CF]?��ĝ��+�4�y��_��4�7I�'�� �����	��Y���� �<�����{�&�ˏ��6{~������2\,t,�������<�)O��O��nrp�ɴ<ת-8N³G��h#��.r��KΦM�IU�i>�I��MC�i��dI�;da��&�5.��eȎ\T���l�y���-C�l��mȨh%���]ں�%*��hL����H��t��"� �ʄi�'i�Y�̖����8�Ԩ��k���Q��#x�Dt���|�lj�L�%��ث�4�?9�O�\�QS+`�eYa �;#b>��3O4�c	�&�s�2�Du��5��?OD}"�# �=�̀���V2��"�瑱U�.%:��^=�T��'=}�9?�'���~�h���Y��Ai�/�@���O�O�l�5�c� �OI
�C�"2�����ܼ���.O�=�'ٰ7mҦ�͓��'��"��*Ო�עN�v�RU'fJ�z �II>*HH�0�8���" 4	d�Ei�'G ܀���	k�Ա*����y�`j�<Y���D3���TCش�L�i�oE�Tm�ܣU��WQ\���[~��v�^��s��aܴq~0b�ĵE��\YևV,(�I�iA��'=��9�'���!l��y�lO���
�G��r$̼9���c�n�|����<i��?A��?���ԟ�U�T�S*&�X�6&	�D���6�ӚtRa0O��d�O����|����>��%�fX�z|�H6e�9JےL�t�w�\(nZ�?	�On�I��I4� �b4Oܜ�F�A$6H8�*����R��O��G�f�n��)$�d�<��?y��T�:�TGM�+�|Z��H��?���?����������b� ����,
R��W�<���ǯ uv��Ee�~�	:�M+ҿi���ġ|�`�F��a�%�.D_}��I��IFXT��Z�~�6��'Y�tj�	T���9O�M����6�r���iH�yR*F�'4b�'��'��pYã}�<ӨN55�р��β��RO�Oz�o�4t�	֟8Y�4���|��'���Cu�V�H�&lC�a��o?XHb�4���'|ӊ`l��>�X�⤭f�D��[����K��M�	��@	4Rj���i�A;R��UJ�G�\y��'b��'0��']b����H��Ef�4'�۷C.剁�Ms��	�<Y��?J~ΓL��l��꟤q����ww��� .���(�M��i���D>�'5���q���n�j��6 �o�������S�L)-O�ՓP*Xm�2�;���OB�䛷km& )6 A���'nXB����O����O�dK���4����p��t$
�a���:uB5k,DX&BA*<s��'"�'r2[����4qn��O���`�
E�,���J�5P�	��J/���'O�"��4�4�c[m�Y�'�Dn��Ѡ�]�X���ac�*�~�Q�o�ϟp��џ���ҟX��ϟ0E�tl��o��<Ʌ@�/?�f�Qs�>���Orloږs��:��'Z�Ɉ/��M���Z�V(�є��8��IT}b�aӈ�lZ�?9�$$���I۟\�#�Z���m2c3�����k�( "��JL�F�&�$�'���'Z��'*���Jf -&Fڼ;j�k�%��ADT���ٴ����?q�����;"��ڦ��
�(D�U�����#��?��]����4rK��,q��h'>5�S�>��Ī��@�T��p���*�@��c�
r��Hpuo�^y"�O�Ly:Aթ1O��h�H�%R)�̧5�n|Y�L��~y���O��mZ�
�u�d�:l%p�k��,s�1��F??��i��O�9O�PlZ/q�z&��	h���(D&�Jt�ڴ�?��C,j]���?�LP�%,0���[H~�jǆu3� �2�\-}�4U�hY�gm�'��X��D��V.�� ��ȁkc�����Q��Ʌ���'h�Ԛ�dOq���ݿ?$�a���x:���n�dW�o���M�'����?����0���%3� 牢 �������^
u��K��(�Q��'MMР�@�ߦl�=E{�O��9Vl�� h؍`���x�cQ��V�4&����4YÒ�<asa��,���3M�/�0�bB�E�?�J>)fQ�`ܴ_қ�4O(�'q��M#b�V�xȔ�ᅕx�$����ĉGj�)���G�;?���X�1���7�y���_���h��{������<q��h��$��
q��٧�W�n$�$�`j�s)�~�V��������4�?QM>�'¸��ŏC'��i����	 ���`��>��&�y�F�$��|8��?O�dU'C(�4/Lk\w�Rm��,�>ռ����+^d}kO>���?a��?����?����?�S�'C0$���XE�d�b�<��C��	��lc�����D%?��I#%"i;��y5J���ǡ%��ܕ'xv7�GզyB��M�+�R�I���p5nn�	ԯ
�K�Dq��\�H�� ����<YŁ
��a�� D��䓊򄁆��[�Bي5����Ր1
����O<���O����O&�P��l8�~
� �M�4_�]�`�+�H�L�έ�!�'��7-=�����K¦�rݴ��U��h�RW� >������V@r�F[~� �J�>+u]��O��7r��`��6����ƢD�W@�'��'RR�'�2�� %��E�2��=��	b���/����e&�O��$W�����Y�� �����&����ۣh3d@BVJ�Hш�`Dk�?�޴�?�D�i��7��&��r!��R����OlT�4�N'��R7�
.J�Ez&O�d��S����'x�O�ʓ�?Y���?��-� 0e�8<�L+��eS|����?Y)O
�m4W,,�I˟���p�į� Q���#R������d�x}2@e�\an��?���Pnt��"ȫ�9�ԭשX[�XY!�]�.-��*O�i�?����%�$�0�Ȁ�@�\x�T��̇�>����O��d�O���.��<�ѿiTB��R-8$L��c�؊s����Q'�*���'q�7-7�	����VѦ](eC,:�*dk�l[o\n�ҳ�ݜ�M�U�i ��(u����Q0JF��2j	�|���'r1�<[d�I�Trq7��">��]�Isyr�'��'���'i?�ti��	�c�Ɋ]��L�B����������$�IٟL%?!�	��M��'�:$)�֌g��iJ̀01 ��w�ie�6���� �'<�O��Ij�  �~�.�=U��Z`[Pթ�Z��?�d+Y�y|dq�e%D������O�d-Vd��&H/[�VAI��h.���O(���OL�iG�F���t��'R��,
��}�T	�k��� g��3��O�E�'AV7�
ߦM:���J�"Q�*��"�	�I�0��ɥ4��0�V�=�n�'?��u���2w�p�\���d6h�R�̌(�l�AH�O&�d�O`���O��}"�'o�d�d�OY��b�A�YOA���oi�& ��#\"�'T�6�;�I�?uSp+�|�z��e�̕%#>�0uG�H�ܴ1ڛVEi��U3��[v�I%�kVN�3B��@&�l{R�r1�b�{Qo�Ry��'���'c��'���ɢ!���s��6j4��%�N��� �M�6���?�����<���ry�q�%S�3#$�)e��jn���M;��i����-�'k
��JD&�	a|L`)e� �c7�؁u
Qj`r��-O�� �"H9q5��Io8��<VbQ�l�ډ��Cf&t8['���?q��?1��?����$UƦ����`���#��440�)3� *�P����X��4��'��� �F����I��E+�"�8<�U2ㅒ(4z�*ԎܴB��	*Q|Ҡ���k�X�'?e��;)Z��`�FP��
�FN�c����Ο��IǟL�I؟D�	p�O\�QfgɌR�h�)���#��a0���?I�w�����yr�'�h7M=���& ���)�A<Z&�4`�N�R��`�I\}hӢ5l��?�: ՘y�����������s�EC"R�Yr4�ִr6�-��C�@Y�'erY��͓x��6�L�@Tb5:&��O(h��	P�I�Mc�� Y̓��O)��u�]�PUp���N��>%!.OP��'��7� ʦ�Γ��'�zTB�(X�ā$P41�4�F�ա~%䰊�h��AG��'���,P?��20�ė�;�
�q4�IY����a��E������'����DU�:���)�6H#�o�'w����ǐS���ܛV�'Bɧ��'�L7�>b"U����0_�b�vދt���oZ�(KC�1W� �񟸪�+1e���H�8?!Ԭ҅+�4ȁ҄���@��5��ӪmZRyb��M�f�R���x� �g�	��lnڠXTb�$��l��3�MC�w�����Uzi����F"��R@�i��6-|�L�'����O��c��B�,(�'=�)�� ��&2R](4/�����"��'%��dT�~��}8�i>�Γ>���w�O�~Y�	�43�H��Iy2�|��y��;���*j��碒�&+n�1���Ɲ�?�P\�\޴*��&2O��' ���8�M!D��(���������XBd��#�h�;��+?��'L�19�ybc��0K��[�������JC.�?���?q���?����a�XN�<)���!��/�I���Oj0oZ�]=.,�	�8"ٴ�?�I>9����u� ۫ml�<���B�\��Qj��aӔ�l�b
��Ny�l��3܄���̈́YE: ��Ȏa5�]��G��.0�!��#�A�	xyr�'��'�r�'.B@ �����F�,u�����ā�6�剋�M�7fZ&�?a���?!����'1���L�iwl,#��8!v��tR�L��4ě��OL���i�F!�1dP�v�dE��KE5'��a2"��O~�A��<Q� |8����䓁�D�2<i���I��6�W&X���$�O��$�O��d�O�/T�f%%J�2�[ e?�9���֞=��0WM6e���~���5��Fq}�Fg�*�n�5�?ٖ�_�­
���<�T�A G���U�f�x���� ����\ ��'���K���,�2$"#���7 5@�4  �'B�'02�'[�'`>1X��ހQ��r�#º��4����O����O�Po��&_��x����'��	�j��pR�O,�<|#�jU�$���J}��rӈ!l��?���S .X�����ܠW�"P��P2�<A$��G��` �cO?|� Q$�d�'��'|��'��	���R}�1�C	���!6�'��U�,	ߴU\��?��������t��d�y�ޡ1��C�?b剱��D�զ�8ܴIF2��d�O�ƍP4��.�$E�B!�� ��eܘks�tx`�R�:T�I�?�p��IQ�$�Rem��yઽ2������(�ٟ�������ݟ$%?��'*7M-� ���f�@B.	�$�T���΋j42�'��7�OO� �'!t6���V*��&�����b��yo��M� 	ޅ
�xp͓�?� չzK��ig+�"����&��,k��2�ƽx�l�h���d�<��?���?���?qϟ�!���6}�L��팷P��q��o|���Ǐ�O��D�Ob�	�|�����F;��T��(G�uZD4��ChMPbbӜtm��?i�O��������k��՚�9O1S6�͇m�lͺ��`�`�!��O�|�`�I��V�C�"���<����?� �Ǽ:"�C�)W.II8�2�"�?����?�����ɦ������@����T�a��"�1s�- �d`z�j�A�����,�M+$�i�����|�P��_ ��T��1t���K�����$�I�OM���4�оfl�d�'����^�~��%"?O�Q�5Ƅ�:�6��?zS, �u�'%2�'e��'��>u�U�v9��a�$I<�ƕ�#�r	����M{�DG~rsӂ�8�S�p{ؼ��툌b=h�c`Ћ&������M¸i��6M�;+�F�۳;O��d�#޾5X7�Թl��(����HԺ���2nD��L0��<��?��?!��?�S�B�_R�p�,9*6΄��*�R+O\-nZ�q���	ڟ��	z�s��p�MF�+��ZD$A-q\���$���[�4G�����O��4��3��@�YJ�8������3�"���bQf��� v�t�&`ɋF)��&���'���(uBK7�R���8@�a��'rb�'���'�S�p��4E�6��O��K�
 M��@5��dq�F̛���}2"`ӈ�n��?��M�4t��#��Y:AJ���L|���-��M���OT|a�+�X¨�[F&�<��'DR��T
402����W�� 	����?I���?)��?���?a��I�1F��Q� b�$�1-N�G)R�'�2�fӆ�qט��ٴ�'��!�ɕ�
��5�"A�u�! �'��I��M{7�i!�dH\�3�%Ӟ'�rb ����
7C�w���À�;Tm`���T�L5���|�_�<�I˟��	������Y�!�쌘g�OⱡC��� �	[y2bi�x�Z�L�O����O���}>�Q�JIgZ�X��DN��S��<!QQ�P�4�&��O(�`�i�PON�)�(��Q�T�Z��J.TʡK!O"��0P�<���@��#DcT���A�V���%L�EJ"����\r�X����?a��?�����'��D����fN��j�|$��q e�s
�n�	�\��4�?	K>�"^����4`���pdV:�ě3E�d@�йi;�6M���Dѳ6O��$��=:e���N�o�F˓
[����1%���*N�)�4	����d�O��$�ON���O���#��T4`��(#JM.=��xk�@՞�M ���?���?�'���O�|mͼ�3	#�~EB ƥ=��}����Mc��i���D�>����
��ghre����<aT�H2�IS$��)Ki��C)O�?a%cA�8��y��������D�O4�$\,�� zC�(�B) 3�Y�0� ���O��d�O˓��&gT,�y2�'2���&��C�S]�T���T�&��O�\�'��7�R��q�����C�-~<$�!fWs���C7�d�R�'v�5MO�]m��]����׆�C���<y��K�E�T�`���y�x��a`�ן���ܟ��I��"~�'D(I��ǈ�l{֠��۵o�L�+�hC��E:���ݦM�?I��i�L�s'��p���ppٸ�>�f!v�ʰo�]�y�x�D��v�l8�!�I�&89��Z/�r�J��E�FHd S`�a��SyR�'H��'b��'��B��Q~I�$Σ1;	�1DY�����M��̎����O������32+�y���*E|R4qcDH%����'�7-]ʦ����ħ�
��%��� ������Q!+��@�^"�|�,O�\���2Y�(���?�D�<�g͜�;�(@`u��U8�sQbS-�?����?����?����d���]+�kVȟ���#�$z,Å�T)?F�Vٜ<"�cӆ��4�d�K}BFc�n9o��?��%2@o�pr���#�R��������d�����?v�<��,�3C��9�'Z�t/���s���@E@y�SË ����q�'��'dr�'���'>��#	�<6L���+�`�$�O��D�Or,m�3l��������s�4��'76�OG(H����n؁6���e�'����M;��i���JT�pc�'����;�J�0�G)N��H`N�7=�\�2�	�=Uv ���󟀗'��ĕ)vy�}၈ѷk���BnC	DE��|��d�����<���ǵ"�p��ȭ2��p��Ly2��>��i��7Mx��%>��ӥ!Ĉi�Q�u	�[5�27Њ�2��7)�pyy�+?a��SX$Ò.��'�\��r�I)x���³[�R��.O��Ĳ<�N~�'��7-M�h�f���ђes�<S1)T�n��xe�����4�?YN>��<Y �is��S�NB7P	"�ݲ0{"��Il���$�9H-ؼ[f;Od����>-΀B���:Ma�ɿ/U ��'��,�VM�%|�pi&�H�Iey���en"��ը f�p ��F}?��mZ�S�c�����i��$Y ?�H�Q�W�X�.�(@H�.GP�7Dɦ�̓�������O��Q�g]Y�ܢm�⤀%��ѣ�d͖o;��$�!{A� rK��RKԢ=�'�yB�2j�eP�̸K'�����?!+O,�OVTm�J�c���V#�%-�Ф T��S�H�:�i��\&����O�lmZ��M˛'���p� ��W$��-�3�9D�D�O�ɰ/ ���ᜟ���i'��#���<��
�h��H2q��]���ӟ��������Dy���a�� �5`#ɒ >ގ�&&�=r��'�R7͟������OAoZw���FN�!M�0d����Xb�ܓ0Í��?т�i�6��ئ�if�?s�����8�	:,�Ĥw�m��ᨙ5TyX4��c�M��-&�<�'�R�'�r�'#"�'i��rD�_%Kp6�r�����Y�� ݴ�p� (O���.�)�O�014ԧ+����F��ӥ�F$r��� ��AvӰ���_�S�?���9=�RU��|�6���FxЕ(C��WU�l�'�����P���|�]�İS �� #8�c�ͻl�~�v�Jן`�	П����\�IWy��|�>i�7�b� 9�EŚcU�����m~za�w��OVem�z�k���M�ói��䂸2���e�Q�{C�d��(�+�,5[��.�y�'�!@����|��X���S>���$��gT�zTb�70�D0����|����l�	�<��ğ�G��%G�M��%y��^�w��P'	\)�?����?)ճij$��'�bdw�@c�TXrA8��U Ӡ�(Fw4- `nş��'u�7��ۦy�f� F{�h�I�
��ɋ���<�y��!/>{�ɀ�懁k�c`�[m�@yB�'�B�'F2��
\�(�L�Q�~H�����2�'��I��M�#Z��?1���?iȟ~��sb�#(���'��6�N��T���O��oZ �M+�'@�O�� ��m�dɃ+�ln���օ�*i����ݸ��|s�P���S�W�Ҵ�C��[�	�'s8�ɷBR�\�l0�bӆ_3���ϟ�']���P���۴$z.�� �F?�0���)�f�����y~RGtӠ����Od�l%�.��I�n�$p(⎟�2b��4pԛv��1
��[�'���Z�_�:R�a�/~B�I)BT��dÆ>"�Z=��	ٔR�t�	xy��'��'���'FR�?�&M��n^!{V��&?�v��2I�����k����͟���@��'��7�u��;v�ЎL� 3���1:�&,iю^���4�B\�����?��)��H�Bg��4CN��8��� h:4�Ԥ��4iP.H :+~�֥}�	@yR�'���%2<ٹ��߆`OZ�@�)�b�'R�'��I��M����<���?�a�0Jn� �6A#vw�����G=��'�2�j'��Ik�����F���DP�d �
O�7T �yCŤ�?i�?�p��g���8��-O��� F�X@Ax��i��*?�RAa��"(��L{�m�O`���ON���O�}J�'&���3�K,:h}����(����\�V`����'�(6m�O�Od�iG4YΔ�H1O�&Q1R�F�ff��T��
�4`U�FJN&3�6�q�'�Ҫ�#��U�P�C�,͞1�2H8Xoʤ��+ ��А|�X�0�I������ҟ,3�d%r��r���8�g�@Gy"/zӜpP���`�	n������V�5�YS��
1��.<�Ɋ�MS�i{��$6�����M�g,JM����c�:ݢ񯊍5|��pm�5p;�˓46ʠi"�Ϋ.�`�L>q*O.���m�\`����h�W@�<1��?���?))ODmڡ-��	'p|!9W�Y14T��`�G�&D�Q�I��M3���>�׀�l��{ִi،p	ìD7m�@%�B���%(�:�Ntk�'lO
!�v�ʠl�m��I�?�*�;E��t����8#��P퇏Q�l��	���������I��X��j�O��x8��YU_P$�#j��H�@�c��?1����ۨ��dDۦ��<i�g�	0�tc'�@�=�U��k�,�?�O�Am�M#��^#,�	�N��<��KMx��6#E#j%� �cۚ(���8!q��cT�\"������O���O�����M���u�2�+ԩZ�K��D�O�M
��a�Z��'b�?��F-ԣU ��Y��A.=�r��%�<��T���ڴT��6��O��B�	�E���t*I3�@�@#%�,m}�JV�����C�<���$��2ǌ���$�8�Ġ̀,�h@�UG�0��<Z���?���?Y������DP��5	6ꍙp:���Cb�M{�I�TOի` ��6�����f}�q�L��Ӄ<xaء�B�N3Ţ�@B�Ϧ��ߴs^"�K�L��<���<�`���f�8��K-O�� 
	T4� s���z�vI�2��Ob��?����?����?q������jo������,>{ ̢�
#S��6��4[����OJ��9O@Hm�<i`��n��I���Ҏ�ء�� �MsQ�is��ĥ>�'�j��P�n�#�C��<q3㗝`�D �x.0}(C�Ԍ�?���6	� ����䓉��O�䖵v�(����7� �f/�����O��D�O&ʓ��V�F;�y�'�B��#}0�e��gJek��g� �[��O���'ph7��Ʀə����ɓL�h�Ǆ[$.#���%�2�'iL�Y�=[��]�t[�T�� }���#v��<i�ǅy�n��vAݜYb��� �ԟt�������PE��1O�|3�DH$�Y9��q�:�3�'7>6��=9��$�O$�mZM�����Ӈ\E���*0A�1�W^�<�w�i��7m	Ц�X4��^���I�x�bb�ȅ�C&nv4ѫ%D�0�P����86���%��'y�'���'���'�N��'��X �Y�TO�+~�`R�P�<)ߴ:��K��?Q���䧇?Y�.��-�~HСa�C�`�0�<���>�M3��i��;�	��x��8D�q�"�-�@`JEɈ97��%��H��U�F�=�L!"0��=d�CJ>1(O���N�'P܆ى�_:���n�O0���O��$�O��D�<���i�f�z��'�F��B��cƨi���.�����'��7,�	��$�Ҧ�ܴ/"2�	[�<���B
?B��j�!��e����S�<��X�%Æ@�X�v�J,O�	��ߥ�fG�-���q'��E��Ot���M���?���?���� Z������~`�`���[#J ��P���	��M�S���?���tK�V�D�0n>�h�4�|���μ!�f�ĳ>Y��i� 6m��eyV��$��$�O�� ���"Y� �� \}��(ᒉ�b��|ޒO���?)��?9��<ب� �[�B�P�3�٬b������?I.OanZ+H�|�	�����?q�'.-��-��OW2#e�=`+I(y������N˦��4:�����Oj�˂B�?<%�"�.k$���^x�C;eA���0��W����(SI>�����# <�+��-r�)(�H
��?Q��?��?AH~R(O��l�@������lw ��.f������D�	 �M�����>	V�i��Q� .�E���A�8���F(r�`�nړ`L!`��4?a�Γ1�,҂ O���)�wM}1+6ąZ�u�����'O��ʟT�I��X�����	{�T`�`n�٣Ga�%��G#��T�M��f<�?���?��'��i�O�(m�Ƽ��I+	����a�OP[��rU$���Mcc�i�z�$�>��'���'r��IHĪ��<ae,B4i��0tU(<���G�	�?q7JX�>�td#��^�������Or�$�!9`́�'C�0���M5?n<���O���O��0L��*�+�y��'r�:BB�!KJ�,�|�@�n6��O���'d7��9������7Xp���_�PD ��b#΀S��I�!��C0c@�:S�X&?aP�eϭ9�ϓfc2�Q�ݗYJ8A@r��(^�lX�	ɟ��ן��I`�O����n(`8Jp(]���(eSR�a�n�����Xc۴��'_�tF�K��lJ'
�)q.�!�*\V�rLa��ElZ�M��iD<G�� �')(���%�j�Ѹ���.>�۷@V�E�q��	�8��'��	����	ҟ��I��$�I�E�ޝ��E	�k���k�h�>��0�'��7�Y#U����O���3���UjrU9���\:&��PT��\ɬO�qo���M[��'��>ݩ@������Ä�$�}�5%�1U6��
���Sy2�&3<���q�.%�'=�	��1�W�]�-P���(��	ޟ����x�I럀�'��6��K[���t�Ȩ��&����-*�B�LTl�$���?A�^�޴*���Ot��%�@]Jt��jΩ-$�Z	�$4�l��OhH�gc��IZ��Y �$�)���#�u3�Q�cR�F9��q�	�O��O��D�O����O#|�3���>�>�ɓ(�0f� �������X��ߟ(��4*��l����?���i�1O*��l�4":d�z��_�p��^�"\����4b\���O���cF.�y��'�*���S��b�c���O��)GM��R��=[B�40��'��	�$�	��	"u��уt� FV�qp�_&7�R����'֢6-��1��d�O��d3"BgӔ+}t�g�O>��0�_xy�d�>��i�6M	՟'>5�Ӟ<��D����{�(���ˁCX�E�C��&��U�Giby��O\#5��!��'
rT�B%��?�\|+@iL�펍�`�'B�'��']�O���Mc�Z�u��8��	�	���S�"���'�$7m2�����@⦭B���Q��$��ǰsB���Fh���M��i�Ю��yb�'�@	��C "��I�7P���$M�=Q�sT�\-zRUZ�+ȟ@�'���'m��'���'���>���%L	*D%�FeEp<oڨ W��	���	_�s�ȓڴ�y�cT&'N��S�B��?���LG�Dr���`����z}��Oa��O���p�E��y�D�c)\��B�[�fb�����l�R��e:��E�.:X�'d�I֟��	c��D@�E)�虑7��#��|�	ȟ���՟��'o�6-ǔ)��d�O&����nېxSdI-q�>�T��?b��êO\n���M3��'Z������"Q�ytU�@�S.UʓZ%搈�
B2p	�K~�NO�w�z�'�r��'� '�M˳O� kVP�s���?����?	����O����Z�y�)�H�ּ�&k�'g� �	U��?y�i>f�*�'��'��'���x	��3�/6,J�:�ӽF*����ܴ?���A�_���'1`׹ln�;���ǰ��ȑ?�)�C�G7Rl��1w�|RS���I��������	� ����3,}޽�'���nN�dɢ��ky*y��tkV6O\�d�O���|�#�ԝs����'�rh��N#'����Y�<`ߴ��v��O:�<����p+u�S6�BEB��H %��E&��u�@��'�<a�\ �!31���䓠�$7 s��h��J�vԻ@�'qB�'���'E�S�H+�4|;�T̓2�|���E�2R�a�g�ݶ&|�t���>�v�'��'�|�]��֠f���I�9�b�@V�Xe�� ��A3�pو JP	d����O�0Ò�N��n��T��<Y��BC��6G�
�y���5'��g��?y���?���?����?1��	��<��v-�9^�x'�C��'��b������xY�4��'���``�qH��mѬt6�s��'��(�MKҳiq��73*�Й'w�f�%���4G�	�>�J���Ah���w��"tuH��`�|bV����⟈��՟� Cڌ2W��i1�� 
2)�f����	Jy�@k��=O\���O�� �,!vO�:3N4a�dU�g�`��'c��6��vaӤ��U���?�I�`S�&^՛A�c��|h�d��TO[�����Ҁ�'N�D�5\�b�J��|R�C >�,T�mG�(� ;!ErqR�'�2�'���Q�8 �4/)�y�r�=
�ĩ����@�a9��G~�g��d`�O��mZ�xWVܺ�*�}� ��!�H�ej���ݴG���/� bn���'�"��::�t�C�b��"�剫�fTxCM˕[�!P�ոt=�	�	Eyr�'�2�'b�']"�?� �*$��������"��	���g��4a�?O\�$�O ������	�3�
 "L\�?�`�桅�D T�x�4 �Ƃ�O�듸B�'����~�@�� _���De�=f�r�ZalO�j,�C�VT����mڷ�VtaM>�)OZ��O�����%�6�!��˱R� � @�O
��O���<Q��i ܀�E�'J��'�B���"#g̦xVF*��ű���z}�i��nڙ�?Q/�*� ��d�As�MՇ}t�h�]�� �!�(֑h��Jm�1�&�X����<ɵς�+�`�mT�Z��!0�@S��	ɟd�Iʟ�F��:ON0(v�܏���1���M�����'ʶ7M�!����O Tlr���Bv��S���'N5k\<����?Av�id7�Sצ9�-L�2�@�	͟��beߙ���	��(P;�qr�+{t[��ڇڜ%��'f��'�r�'B�'���+"�J-N�����-z��1V� z�4C8Ȼ(OT��8�I�OVm#���>'hp�R�G��}z���0%Iz}��{�ĩoZ��?AO|��'�b����4���ّ5���2��S0gDMK������D�+��5���� Z$�O�˓IB�(��(H\�%�_8��8���?����?9��?�)O�5mڹ_]��	?� ae���K�x�f���@���I��MC�-�>)Ļi��7��ߟl���T�F&����3d2��`֣��	n:�k�=Oj�$�	b��@A�?�˓����wV%C%�L�* B`Y��i�,a����?����?���?����r�-#y#��ɜ1.A�@�Z!�?A��?!A�i����'��Jc�Xb�PZL=Ee�)�'[El��IU���'�6��������z��B��4?�Di�'\C�u�AAׯRezY����tv��bK9>�rN>�/O����Or���O�����$v�\���*T�xG�� 2��O��d�<餰iE|�s�'~��'���Aa	�	R'h�N���eY'8d���O�h�'��7�H�Y
��ħ�:Ve�K�Ե.U'�Dh�K#+��娲�D�J��=�rGSZyR�OȮY��$�	M�'�qi�g�46l�%5U����';��'�2�'�O��ɒ�M�f%�n��20劯1�H+�H�N7?1��io�O�(�'>6��-n��A�쀙)�؈��׆rc��o'�M�C;) x=��?ig�{&rxSC���$��{�a��C������.ӲF�j��<����?y��?���?̟�	Q�I�j2���i=;���#ggӺ8�p=O:�$�Oj���C���̓[��@�FN�D��!	&��ߴ ��Ƥ�Oz��*�'�bp-Ŀ]L�Γ �"|;�H�'7<=P�#óxY��M���V��F;�<�K>�.O��$�O�����P�H������)�T� ���O8���O�D�<�f�i�x�'���'�IC�hʆG�|Փ��ъ+g�}�v��}�LcӴ�oZ��?�/���,��p�.��{�$1C�U�0�D�&RȰ���OH�Ss�@!���O�< M7�J���M�,͠e0�Fǟ��	�����ӟD����3�yҊȻ,Y0�2AF6:�$��já�?�`�i��<��'��'�'��MX.U��nX3P:�(qua ,@�����E#ܴ
I�v�� N
�hz�'��&�;%���ׄ�2,����Q�	,���i$�-��ݰ��|2�'��IܟT��ş �Iǟ�	��4P�ː@��OP��0���Py��d�}���\�[����O��'���9�X!���/`T� 2(\0NRʓ^؛�j����I���O���O ^\��N>3�	�թ� ��bT��E8,eZ�U���fZ�n�����c�L��[y2�ˁt�ʶɒ�N��ր�yl"�'��'[��'F���M��
]��?)��;$����I�+����#�?�g�i��O���'��7m������N�$��F��nK��+�A~"��2h
�͟��L9�p<��L{y"�O�0֘"ST�R����zE��j\�>����������I����	��� F�C5w����	+�>U9��ǿg�ʱ��	!��a��ԟ���	�M30���<1��?)���?���i���"�T:��p1�ĮP/8�1�`��.ܰ�j�wG�vciӆ)l�>v����F����	.3
�*%E�;Z�6��[)��)�Ĥ�r��CNւM��'�^���I��t�	�x&�m�t��89�&X36��c9���	�4h���'q�7�@<��I�O�����	A+���xr��%����� �L����Ox�`$��"i����I��1�O��Ԣ�a �=r�b^7�4ERBn��	��TGN�Lh��	w[��S#�¹��-w�ɣ8�\���G��gh�[���W�M��ɟ��	�D��l�Spy��i�nuz1��2�)j�-�%���:`�Q�E���O0�n��<&�D��O��oZi��`�#V<u��qA!��)4���4�����P9XP��'(��<wq�E�p\�Z�X�zw镪06�����	&�B���ky"�'"�'���'Sb�?� �U�C���V��`�*x�DæH7�V���Iǟ�%?��	'�M��'��!��BR�L��01ˆ)��8PU�i]�6m����'j�$�O��DeͩbEv�ɞ'�ny#,ĕyZz���ֹ=�l����'�B|b%��-'kl	�ß|Z���Iߟ�������)Ȃ(��
�2%I����Iҟh�Iy�ca��`a��O��$�O��i�g,}¡S�-��'$�Q)9�I#��dҦ�`ܴ!_T>%b脤2�D�J�
�y�E�J�O2����P���5fQ�w����	ƆFh�ٝ'�f�sƜ5>r�E"�մ?@4�!��?����?���h���I#;�d!�eJ3-���ف,L�x�Dަ�i�g�џ��I��M�B�O���`���5t��(f;eV�y�c�'�06�G��)�޴@]�0x�E��<	�/�HTb���P_.��u	؋APB7�OsH���ˋ��'J���@��ӟd�	� �Iu�? �M���F�G�V����ɫX��l�3W���ܴFO�j��?���䧻?�� Y��Ш!��S�"L�s��,K�I=�M3c�ip��D)�'/Ǌ$���	1c���b��U^�YلJζ
h�M`-O,yѐ`�0p�&�i2�8�$�<1��=k���"d��zfv���OԳ�?��?���?�����DR֦a�g(��<� �@.��8eo]����Fc����ݴ��'3 �nO�6FwӪ��7fԒxQ��/.���_�1�ّ7L E����O��Xe�-/��`y�ǥ<)�'s�'4Z�BɳB醖.i�����?����?	���?)��?Q��-O&��jцP�t8`��эq�'eb$g�~9��`�O@����9�<IMǟ!��d��@ �FZ�lр��?�O��o�M��'
�Α���A�<���(�2�)��#v���ĉ'�Nظ�//d��S������$�O����O��$�7Mu\	w�Z�L)�T�S�*Y��d�O�˓w��V̛�9)��'b��?Mr���1|r��Ь��Y�8)����<��U�pq�4"��V��O��J��ڽ{ep�$��'�z<�k�=W����# 'n�m
��<���|�YP։���}K\1��h�&f v�8�_"l�fE���?���?y���䧝��ݦ��� �E\DbO[�x�H��ԉ�5l(��	�޴�?�N>i_�X��4Uɨ1�Xj�. ��Å�w{�i�׺i��7�W,wfh�p3O���7j\ *���E�
˓P{�A	�'Ν*堸�e��h��ѡ����d�O����O8���O��$9�b#��?!�.��Z0���@Z��M�c�"�?��?!����I�ON	m�����(�~[����^7A�$�3֌���M���i(.�d�>�������aԤɩE���<��b�)!��j�Ҷ]h,JD@�+�?��кJ!���fF!����d�O`����#����߳#��X���0�
��O��$�O�ʓS����٘b["�'��N� j�)�R'(Y(��d]6�O�e�'4�7 ��m������Z��*9�@Q	�1>��'�0�i
�	�Y�W� ��O"бC�;!�֮_�cj@q(\�wWj	J��å�y�Gż*��
T�	lE�3���0=�Ķ ��fȫ8'�i1�Iյ:o���ѩ@"��A�H/�<�K2��>*<tMj��; ��rY��u9��(��e�i�./�i	foQ�Iҝ�DI��}����&���9��ۆQ�<�qaKڜ<Fty���P]?��a&��z�Q�:�u@1��1.��Hb h�n��V"�?@���x�,�0t@�1���?�fM���𘥈��<���?9�4C.��2!�c���`��v�t<���?!���?�����Ofʧ�M�`#[1:��!��) �YB$���3
�I�x���x�ɗ��#vl�	\P�IѦU����3#���0��
~n�ZЏW�e�9q�Ǜ�B�f�̓�?1��?����?��t<��F.>dX��X1�^���K�ӟt�'�������'���� l( $X�݉^�8��t���	�Z���2�.`��gg,����ʣ�?!�'A'&�R�(Y���� j��A�ĕ�$�B����J����?	��e�����<ͧ�M����Y)�Y��!�;
��e��G���'("_�\��ٟ�%?lZ�&�Hrf'�"x�ș�w")?�:e��$V��?��fLm!�D�9����?y����0e臭��$~���d��K��*W��#
o��B���?�����4� ���O���>�р^"C����$�tuX4L�^?���?�����$�O�$�O���G,``P�<<�a	�����͋0J�� 0B7��O���*B�d@2P��N���OR�Dd�l���l�]l=b���J+��O���O����O�ʓ�?�/��6-D/]d��@�\�+Bz����_��B�'x��'&��'�����nG�^�����'���%��m�4���.ǒd�m+ ǏoX��5��FX��0Ol���O�����$�~���Q�xH��]���;&d\�8�RR�L������ʟ�'�2�i'���$ˉ0��4��̞q$�(pb�OP���Ò<��I�8~�z�$��Jx:Ň�6���w�v��Fe�����Fn�=]\��`��O���O�0ۆ��Ol�$�|��|��4D�l��u�D�TB^�Rp�&��C��'���'|��ҟ$��F�$��$���>ED�u��0:H���m!4�0�!'�n�a��!f��A&;���Aȅll@�c�	��p+��� t�-(��3B!@@��Dj�O$�~�#�`�7�8p�6�^�8vؤ�rnJ'dpp
��.+^�e��H�8X?�{���Nf���dX�x��X#��ۿI� �J%� 7f��*GK�2L��;�O�c� �͐x�>���1g�X8��kӊ�d�O&�� 5;C"y%�@�	ٟΓi �Sѝ��a`��=u� �I��T�Iܟ��� �F�d�'|2�';RnE4~NPp2� <����](���'�����!���O��'���/(k��BADJPX����T�h���O��E$�Od�d�O<�$�O��d�O���G�-���cfU�\)t��!�M|<ey�(@��?�L>���?	�`����]c0NZ�`#
-�ҥG3@�$���?��?���?���?V*I24���
V�s�2ՠU���@�g���䓠?�L>���?)����?�gN�D*^��c�^��2ca���?Y���M��BV�Wc4 ���O��N�x��9#:L}���A$Aָq��� Tݶ���ָ.@@��f�"�'��'�rE��yr�'��'���I�p]t�ㅤ�KҐ�!Où-^�|�'!�'@�'n�n[B��:���+Klmc&fN�,1HHړ�'v��'��3���yb�'C��'�.��Fm��Z��t��/��K/�Y�Iٟ̣UDu����ԟ����T��&4��r�HNO�0"`�Z5f�"�yc�?O�<%�	�����ʟ�IП�ؗaŅL�����4�	�p��B����$��h	��P�	��<�'����'���'A�s��� ����j<)Tz��bJ�&����,�Q<h�'0��'7�s���	ğ��I�F#��Ȳ��"�0��d��1��n�M��Jאsd¤Bq�'������'^�;�I3� .t��}{�#3:t�(�@��w���?A0���g��DE� mI�ʠ觢�|?�a�ȓ=l9�CMT�t�X(c�C�4��8ȡ�ױ8�\;'�Á;5�4�i��&TM+�L�e�V�@H� ���� �пS0|�#��L��3�ϻZ�L�jr��8��P�Jِo��%L��(;�ܓ��3���y��ʱN�	*��6(���J�/B�9D�praA�_MH��)ð�� ���c�p�P��l/ �$�O���O���;�M�B䈚a[6H�wϟ�H���Pm�+`�QU��Oz����=8���&>c���0I7`#��
��",��0n�;��F�'i��Ӥ܇5���O.��$,ܸ8�Z�B��H-$��'M��87�Op��A�O^��O|�'<b�i,v�QAdBuӢ)�Àen��'L�Q�aJx�jwGH�d�D���'��#=����<�'������_&XD
FX_�t`�D��+7��͐��'H�'��t݅�Iџ�I9��`�e�:� ��i�  *�`d�޴�J<9Q�ޤF�T�;	�3ɔ�`Rʗ�Y18!��+�(!����S��q�T���s2})	�R��%o��L6��$Ꙗ@*L�)�%�`�V����[��'���'H�O�����J�+�6�cD��p=Ɋ}�M�.e��0٣�B����@�
:��I:�M���ii�	0N&݋�4�?����M��e�>e��t	�i�U ,�!E��I���V���'��%I�R9BLh��5���X�� ��r�p�иR�X�@�	$=o�:���qܧ��9�6�̂V��¦�R).�2�F~��4�?��i�(7m�O �]42�keJ��3����c��<�P�I�T�?E���Ⱦ/�����#	t4x/���p?1�O�-�1�(QD4�xf/W1V��<Z���By���c)��'��Y>m��m���n��6Ty#��E.�\[%BԆ_86����*n
	�'�ƽuZ�m�FeóQ�FU>�&>]P2��/��E�4E	>~V��2t�>�D�F-,�=��ٸ*.��UH�(�̴إF��mج�*�B�PTUY�U�d�fm�O��nZ�M;���H�R��C�	�S &�@�!�II�e�W�>1���hO&O����A4C���!�d��e2U���$qܴj���|r��H��e�Y�$א�i`��2J�<�`�X���O���YZ걘�J�OZ�$�O �$J��yw�ϫy]4��wQ�E$�(�Ɏ�'hʓD��)�QB>n���'aP�fē!m�2�Ņ� ���)�_4��e,��\J�x����ħ�V0hK�x)�j����5 �l�)Nٰ��ա��z<�f�'j�i3��'j4�'>��?�ڴ#����%����M�2��9 V�9��'P���x�)�3����L�
�5f�1�.Q0���֦�rߴ��OA��SGyBL����@+U�$��E+fhʝv1���"�/T���'��'����������|j&:2�p���1}:�c�쁞Ojn�w![�`�ÅF=\O\�%�ħs�6�#v���E��H���+lԍ1��M�P�,��tb)oڌP�$`sr���W���Ы0}���H��i��6��O:��?���'.Z��*Ë
� `�$)��ՄȓX���֌	er �!I�ʙ�O���'P�	XR��[w���''��F.TQ�2�T�4���S	Zn��d��R���O`�D�:n0zYK��Y��,��P�D�E�@��l��陠E���f���O$���W�{�DIቍ�$$���'Za�D��ԇ/�`waF@�xTF~���?Aa�ir�'m�Ժ!ops��]�t@p�XGVH�Iȟ�����D�)��}@��m��iY�q��H�I��p?i��Ox��p��1��P�̈M�`�b��Lyb�5\Z7��O��$�|�mQ��?iݴSK��ӥ��('#����6o<:��'jt5q�ߑ�F� ]�C{z!r� �~�M|��Ӹ~�����Hk$�K��[}�M��"@�Y�
/ �`#/R�w�Q>ݻ�)pY���K!*���jG$�>��NG����L>E���B=|��Y�	��ܽ�࡞��y���;Ū�SBc+cp��c�̨�(O��dj������	H��D3��
|��idERy�O�K�8O����'&"�!2�9x SCu�܉a!.i�@����'�ў�����1o6�`�c�xH����+FP ����an~���I�Q��C!�F=�Fx�厞&$B�Iw������}
�a5�%v�C�I��D���SA�(9`"'"u�C�ɆH^�-9� 2dlv�Q�'GZT�C�I?O�4���<_� 9��-�*3v�C��Zx~�ˠ`s.�ŀпH�"C�ɪ~�eRtl�M��@jQoE'�(C���"���P����$!�B�	S� ��J �ٖD�I*u�~C�)� Lɸ�A�=@LhY���Z�+��v"O�A:@��$k�D(S��&v�$��"O�4y�!��*�(�{UvժV"Ob��`�C�
��j3xip�j"O���dmP�V2J� Ci�ZU���"O�K���#Eg�T+��ƽE7��2 "O�,�A#S ˖T���V)��t"O&�2��ŷ-��8�$
�p�IE"O�ʴ�Z�!����F<%0t%"O���'�G�,�� E�&	'6�""O�a�C�V�4�+�HKNz��1"O�5��#�N)~ܺ�.ϡJְ�C�"O���C��#%=rb�X<,Ŧ!��"On	���� ��2,�U'�Ԁ�"O`1rF90 @)P��?.�$�"O�9
@��(X%ƁR�풇$�Nժ "O��Am��6N\�Y0z�F�(�y�n�Wf���D�''x�W�Е�yroߒ,gM�bƃ�I��)#����yb���D�#\M5�vk^��y2�'?E���tF�v*TJ��͠�y�^��`��K�-b4�pr���yr���A.���2��&\�P�R���y��\**��5:!)U)|���KfI˷�y2�D#4�4�4&Ӡp^F� 4:�y�E�Hh���u��s��%�yR�Ѧw� ��i�3cΠa�F���y,ع;�@���	[��*�k��y򎐘; �҅x������y�J?zAf�Wd��y�@�Z6�M��y�@�+r�4/M�fZxtH�MI��y�"Xq ~@��n�
X��$����' �E�����@i	%jF ���'�6� w��/�ABu!N��I��'4�J7�@%#�x< �a0�`Mb�'Jra��g�-6�`�bq"\�<�!�'��X�͓q�j8iA���V����';�	��>-2�4Z 
)B݆\)�'>�����A,V�6@z@�C�u��
�'��Cڇ9���+�< P��K(�y"�NH~��YvK�z�,���AV��p<ъ�$��Z��������(��A? �!��[�� �d�
.ʠ3ׇ\8m�链hO�<H1&��\�E�9sB`)��"O,��E�R��Ii�%�7 ��A��)lO\%ғ 9#��CS-Y�P�5
O7��6���5"�5">���B$��a�!��'�����MM9:�ĸ�m�2_�!��T�t`��*���*)D �rA�'�!����t�@R�- N�A�!��Ma!�Adn굚�J̧򄔢�A�@e!�D��bl���Μ[�u{�@M�!��N�n�Lmx��>,ـ��shʎH�!�DL$B�<���*Ξ�#Ɗy!��׵AҘ�`V#>b�"��'iŵu!�D�Xs|]��%���"��T�r`!�,:�]���V+q�2�:`/U]!�d��,��s+>zD�{��Q9L0!�׆O_vp���J�f~���`�K�-7!���%-(�7��-r�Ĵ�#=!�7H�r��ca��"e&U���	�ȓD��uj�)#0�`��%H�y��K� {"&����U����n�*T�ȓ,�~�;/'�]�# V�v\i��S�? �ir`kɤ6�����Kÿ�~�r�"O
�[0�.6J�:�I �x��"O�YQ����X�!GN��4��"O�TQ�c�:�2��0S�"O�U��{K0�)�dH�"�`3"O�E@��Q8��M<����"Of��U�K�Q�t�A�MS�.&��b"O���[�e\��PU��?mD>�1#"O���&J��?{.5#�㏋H�Ĺ�F"O԰��I3�E�S�D�2�Z�h�"O�@8�� -#QM��ӻ�%'��y�N�#\༣fH�kڲ1ˡ"�,�y�őlZ� �R�o��f@���y��C<�F�;1�[�,��T	4i���y�b�s1�N&	/h��t�ּ�y�ċ�5D��D���w��(� ���yr�F�>��%�?��ai���'ĨO�i�ȃX�ORبѧ`՘K�}����8p|�#�'8�8�-Ȁ��Yx⤘�,���i�c܆ �1��&O�������u+�8��+��+"|-�Sd0D���mN&yb�`�pi�1n�<��f�>�fÇI���Qc�dX�<"�+�	W�ZP��4T�L���)�OR5[`%ڪ$���jH�*%\���f5)`��D-4,��Z
�'�ڑ�A�O��)8�.8WȉA���97�c��=*��{@��O�4�#3� )D	]�
^�2ġ�5t�KDO,������`I���ǉ!Q:��a�M���pK��n�PbSȟ�ô+X���y�7Pnl�s��.��Y#��'��<��T,��O���G�T;VڪH���ޜQ�
�yӪ�J��[�?.���A� ]H�8�'�On��Q��2Y�^ ���$�#��|�ƙ/��=YA����!�����,,��񊜑F�j�3��#�	11�A��˓��=�Q��5Ơ��e�<}���0E]	&qOZ|�r�"��Q���-���೅�,�^� Yw4����ݡC��iWB"50�Iq�'��<��Ǝj�<I�l��DF�<�O�r���r���p4�J3�� )�N�g?���C�{���f��t	:<�V�|��tJ��z�ɛ��T���[.�&`z��qO�	��΅|��Ѹ���D�:$���ODb��5�4^"@ъ����� �JTd=�Ou�f� '�Ƶ����9�l�7'�$�1�ɖ������
����,lOf�	4Ś"=CN��O�4l^J��+@l����K6Bv���G �?k��'h�|9� D�.IX�{�� *Vp�ȓ�N(S����~(ؕ����(aԘ�H3Wn��Wܛ~�
u�B�	�h��.G-|NΥc�g��.V��c��ݘM+!��;ml��!G�;�4ɑ�˔%q%69��Ɔ�h|���R�\�ZuB�2�n�=!G��?NV0A��"\�ȉz��z8�|w*�`�ܹiqFiL9�r.�:ti�����Lخ��f��)�����'���X�*ƍO\�d��
�4-�Q�L��OZ�$���0Dʇ�IV�x��J�|� �5���CA��+ϐɪ��Dm�<� ��t�+7�کC\`�C�����I�n֣f�iC�(
�}����G�s����
!^.!ڤ�ƫ)���a�"O�H��2(S6xjl�o��lbG��;y� �æE�$���Υs��3ғwh�2��7]U2�
����%��I��9p��(,U��Ӓ��!I���c�� pk���E
�._
�$� �2PJ)QѤ���߼g�r�D|��_!YXmp�
ۖx���\>��+*6x	�A�ؘ[���c� D��S�`�V^z��̚�u�v�%�d�|q�G
zø� �N�SgD�G��FH�k�P�p)Q=ZƑ�7O��y2JM�n���
E=it1���ۀ�ڌ���a�@�����,c�I{�?#<��`��pH>�i� ȓA���S�
{��,�$E���=)�S2j�F\�eD8�)�D�U].��D���>� �QT�B���	_��8q���I�'�)��j�*l��xq+%lV�'u�<�nܕS{J�pe*	���Մȓ9�R<C#��(=Pu�"_:�hΓ4�f�ZAC��*~�}�CJơ8��?EY�N��Y�V<"A��+�\����/D���с��X
���-n�M�#b�r�̓!9����O69(���'�F��L�(4��B�Oxz]��^T��"�@=� ����+F>9!��2Z����@��=,�l�#�!�O�}�iJuG�e�¥�/C�43��	 OW�2�-�t=ʟ�U�7�Įr���0��UmV	��"O�6\�@�)�#��4�l���V��:5��'P��%#F��0|�C)�-$�	� ��cv ؠ$�R�<E�@/�Ġ�l�/\�2�����PF
�_�6i�����gܓK"FM�əHYB�"���O2l��"�Á�*B����NR�o�< �Ƥ;:h�����0!zd"�^�1�HZ �<n���X�� �iHj�|8�l��Q�5��^�Ҝ�̚*n@@�Z����?N��ȓl� �a'��!s���z�ͽZ�Ȁ�ȓ 鮌!᫁���8vfM�ux����!w"��ώ>e�|�z'͐5u�T���HPqA�P�<�x4����?8�-��dQ�Q{��Z�lm
pɹ(Dm��)^J1��#E\�$bB�Y;T𰀆�b���:���54�$��bE�8XO����N��
e �;�p!wIݒzUhh��	׆�g�=2B !��HH�O����̚F��pB4���i��q����D��~�W��1+�Rc-ADo�6M�U	��:D��V,E$.(��u��!J�iiG�7��ȟH,�FU!ra&��Ȕ�'Mj���"O|���O��Hn\�@�呰C��<�"O�@@
�3+���Qd	:q�t�b�"O�� ��/4��q�cR�I���G"O��Ga�9\�:�!��4��e"O�Tr�(��v���JG.D��Q��"O�xӰ����5��W���\�c"O8ZD�"�a!5L�()�Ą�"O�q��f��"��̊H��;4�x
[��zBg�=\�����o���"	��9�!�N=m��a8��=@�5���!�d�.����E�/V�@�C
�;�!�$EuJ)C�iwp�
��8 p!���Y@����.�0����#6R!�DQ��F��B0�ZU���4B�!�$�(a��@9��n�je�����f�!�O6��\��A�� Aj�.��H�!���R7�E�4)��$c�83��Az�!���	 |��e�_,��E
ÆCb!�7zʠ9�(�8<��`�^�Vh!���2�0f�H�J`�H�O��*=!��E���w�I	,N��G>P&!�$ͥ$dA1��Ӝ���# �^�!��3:Cr�sr�M;}\�C�FQ!�D�<;���ɚ>*1�C*�2m�!�$.�X��V�Y �]9Q(�`�!򤓳1v��Z��J�[�0��g��!��eê��#� :`���半�=�!���艀`��?�f5r�lAK�!���X��iȻ_�������!!�$F&<>]��'�=T0Ԋ�/Zu !�_����7�Ӹ!L�����2g!�Đ6n���y�*�"��ó�%2"!�d����ف���?�8!8�K+/�!�dHf�~��.�jh�{�
�%�!�dN�(�V�)I��5`"ؐ@�͑����b��5���!��#|Od�!X�N<x1@�	p}d� 	�'y��Y���	b��HwN9���'���{s� �f߈0����-���'��E��ň>���R�R�,�H	��'l؁��82��}�a�?�d��� �l��k�>~ycV%yV��s"OTy��̑6]xA4/���0��R"O�|��&רn|�)�[�pA��#"O�rƋw��CS�Μ�8%�W"OLPcW�X'(���P�oٓgW`	�"O�!ӐJ��фRt��):��h"O���N��_���k��� 6��9�"O"��AF֯Z� ���)F����03"Oiu���<z`�3(X	]��<;�"O���F,��av+D8�B"OH�I�ێn-�r֫�(ao�0! "O($��bH�?��z�-����,"2"O��'�� >���b�L�;t��J�"O��!�L�n��01��7w9�x��"O8�%��0��j0랹~5*"O���M�*���#�N�d��"O���r��m�F,�dדw�EIb"O*|*!��ٮX��H� �*�25"O��S�+E=DVn�ꆪZ�s>�A`"O�+smٶ2��p�3(޴b&%Y1"O�|�B�L7&�1amE :@"O�B ���9�B���?j�"O>�c�2F��E��-E�}��"O΁/�f|����*w찉rT���!��Y�T�x�Sq.�7�d4*�U�B7!�D��G8��:�'Q��6��@͘� !�D[��1׎ɦ9�<-K�e�M	!�a�t<�v�ȴ���狊}!�d�(-u��Wl��t� F+W�!���#�.|�6;�*�sV�T8�!��
8-H�y��Z�H/^z@�'�!�[2�HܪƁ�:,� �a�]�3�!�×s�΀9# �>0T�p�w!�J#��𨔧�<IL�T/�p.�f��3^�5�#�	��!����OJ��P,���Mp�/B�bՔ�PĤ�NE����ˢ�Y��T��J���0}��-x���E�����K���y��+��8�PB��4{��|��'��)����c.x�����-���cJ�!(yx�q��'ғl�DYR��� ��3!� �|<�9�'�.�*����E���	qϓ ���q����l�Q�>�����A*���k�l`�� �nP,��L�<6�M�M̖B��=}�h�&���sV���3@W�*G�����;sPL�щq� ��V�!Q��qcF�	�:0 c��>�<��K��n��7�>6���!uD�3��?��,D�G��f#O3M��'�1jHB�z�b�O�e3�L� ���~&�#AA��+�$ϙ�j���x7$2�O@��)Jb�J#	9&FB��`j(]�	9`�DT���D�D:	��03"%@�]����*��a�%�Kn|�`N�L����V�L;$��f!ӭo�L�˔�eӪ�Pk��#`�L���\)�PB�AFŦ�s�i��@��#U4
H0ɪ�&�\
� ��`�&s@`���k M�t���E�6�C�5�(iТcUE�|X4�	�Z� �xg�6��pr� � ��᫁@���?��A��e��c�>lJ�GO�\�l���K�rs��C�����?}�r8��w��Hs� �9 OH4`�H#d ��'�Iq`�ٓG`�q�K��X��q�#��'��@��'����E�aks�E ���� Z�I�@ɂ{�&SQBۧpr��a�t��?7�K�� �DU)-���6���=���J��r�A�
�#a��(mZ��B��S��/�_Xt��bBH\Qp�OBM�eΓm����	�Q{$E�p(M��t��;��Ľ��iݕ�FЕԢ5�ebO�H]��'��/D \�D�'�6!;p	�Xb��@R$D�wNɘ���p�4dG ��$MR?g���'w�ӺoZ�|�w
��y�7"2^��J�pj t!ҊǞ��'�Z��We.�d���%�
a���>�7o�.dhF�y�a��:�(�.Vζ��OV���O�l�3g�$�F�{�i��z$(�,��DϬUB����J>i:��L�-����T-��)��%u铆��5ێ{�>�P��i e��Z(�*�h_0��6ЁC"�MsT� ��	����OXl���ıH����G���"�*�s��j��D����	�U�d�����%��0rH��iP�X�ZJ����G�
��08�� ;=���"g�عX����Q�xB�j�,�O�˧���U����� �y:�MR/y�R�cU�XE�2A8���IH���p���r$�@âؑ\
�fU�V�[id� #�@��P|kR����꟠��4�T�RH
�c@5RA��\}�D�(]砸��O� vH��E��o���q��{�f�,$(-�=�O���!(5�tK�[�^"�`1h��M���O�OO�R���@ᑟ�1�Lqф���[n�UHe��8#OџD�?�1Z���(S����X�kG��,��� �1�x2k�]�P倶<��Xz�Iȓ���)DCǡ��	rE�xR��|�� ��Yx��Z+�H)[���;:����"�A6��OD=�Ů��b�4�P�DY�7�8P)��>` E�,�������Y�D��b��<��.Ͼ	�
�D�O�1 dU�hj���МiD��fS��D�:$@�3�M's.�اmí�$��E
�p�u0��N�=ZqO*�1�'���$ER7nwLݳ�֙h��<kf�C?�M��垉;V��8�D����4��O�8����̩ ��U�rM�-qĎ����'��"��Oj9�}�s
������=<HJ��J� M���3���p<)eb�
I�4�ОwY� �ʅ9;ZܕzTi	�E��t�6���ă
��-p3�ːl��s�ʬ|&�t)�.�	A���8ǌ�Y��e�Ԃ$���lZ��V�M�Sz4�u�	\3��'�b �!�H��q�
4��ʜ'�q`�>��B,D30�!���0�P�nDX}�D�EU�9!��˅W#�q�][�-dA�!�ȩ�v�Ũ2b��D8��aª��'���V��!�8�B�r�X�r�l �^�=�'l�sÈ]���	/f0�d9C���&J
��݂*8�`
O@����	���Q��LS��y�m|����I�c�0L��߼�dL}ʞ����:r#(X��GZAX�P��韔B���+��;�����
�3�lh�����O�UZ���o�n<)��5
������h5�Km�8�2�Y3J���:s�7ʓs�~�j1�[>-8�6�I
���'���R��o�L4p�S7pl��	ϓ/L5r�CH�l�.�4 7�$J���! �5[.���ȓ`��q���3Id���c)F��P$���g!V8[9�Q
���_��n�Iㄍ ǅ���C�exd�#��3cE����6=n�xR�O��	,�ܕ��O�|��R�w+�\I[>�2 ��vh<y�ֵ!_���B* � |�pI�T�ʰo���o�'���[!
 W<P�w��$�R���D�<Q�s��dcR�iA��`W(��a0�b�F	�4m�ȓde8��% _�
\P):bl]��9�����$����cF�D�D`��$�8b�D�Fd��帘�����45����H��	�>�>Q���Ua�B+��2#�<����5q��YN۠a42c��XJӰAt�y+1��󦝡�.��yW�39��pw�[=~���ƭW���>�¥G�H1���F: a��W�<o��k���MK��
4l`��K���\�}�gF�4�.A� *A�����Ӭ�g}ĵ_na���\�>4�dz��D��hO� ueַ �0�-r^ 8U�O�eUL��U������Eg�sV�E�x[3�<k�xRr�F
W��dF~Ҁޖh}%����Q�5�e�:�?�үA"�L ��M3���҈�v≋F`0-QA��M ���"A+3[4��� �(-+��*���P�>%��/	�
��f�
�zB,��C�j}��'Ct�Y&��d�z$��Q1�\#5H_�C�X�*�x�� Z�^P9{���d���@Ao"5@R	�q��I	k�.D�c��)�j� �?���	�6��T9$���R+&	�u��=	�i�&T�#b��+�O��h�I^3P&`=��زe��Ш@�Rm4�i��g`rY�d�=Z�6��僖'��s��U�A�B.��5�CN��!"Ȯ��3��|"�g�,Y[P�.���% 8�~b�ʢ^p�DOA��x��*�� 
?K��ڕ�]�zVJY��D"����L؟d@^N肤f�Hh�i��K��x2!-�t@P7�$tx4���E+���4U�LAAY��!��M�\l��B�A�����Ia�f,��O� �F��D�^�yc��!FBy����,�?I&�]�wv�'�yJ ��b�49ϢDI��MF�X͘�*!��O�=�-՗w��`1k�4d�Z_wJDx�U�H2QJ]�gP7Q5�L4�d@В4��L>�'�K"*2] �-\���p�BGyr�Ė0͑s�I+q��H�V��j��h�e�\1t�܌i0��2���ꋦ6�A�~%���癡�@(ۡΙ����S*N ������]j���'�l��&��
L���e�>v�HwK/��ƀ�<B�"��E� g ���n�{ʾ�!�&��$���6S��%� ;��W�ӓ;��%j1O�=\R�s�*�Vv��d�y���:�E�m,�xv�i
R���R�oFY"�ȋA��ݠ�(%��ث>�ܢ��L>Y��PNfvu�C܃7�0�S��D�ɣwk0�Q�	��e8�`��'5~,�mD�=���ɂ�̬�U��6pѐ��D�'i��������ȣNR��s���1,�*!�'�t����$Ԟ��'�=PF/ΨJ��pI��)3�Rđ��� ���j@;zj�@23	�.$bV0HAʋ0|/����� ��1���	Xv��0:��`��dr��T���u
��'T���ϛ�vMcش=�~��b��<�xdhV�F�2J�ٷ�|R�V�r���}&����'x�]k�� �4��q��4��N����p���p~`�{҇�:{	h�
��>|���&�O�LA����^i\��pM@�\�� &�4D����Ez�?�ɧ+��OB�)�n�k,�DPd,�3�V�XS"O�����&�2<�D�D@��zP�O6���O � B�|��1S��O�(�ӰK��w�$������T�;�YqT�9a�r��A3��|� �� +I�����D�I�S&����|2�_�z&���e��`�D��h�9O&���H?ړW�֙�%䑡��l��)ҨP_^z1d�9�a�b֎@���Zt���6�0<�r��A�u�	�g��rk +�V�yRB�+28C�I�p�x-�t��$M��\�s�tOnH�`�����O�ʭQ�A�)`в8��g�a�&�R�'܄|��A�}=8��nG�� ���
S9Dax	�qwDtӥd	�E"&;�f��yڌVQ윉uG�!Q��j�GJ7�!�d�J�!�e�Q7$� 4 �|�!�$Y?Os2��P�R\I��F�G�!�����E��	�m��a��-|�!�$�jaF�JgJ�	e�����S��!��+4�<�
�Ξ�p���cӾN�!�d��Sшa AjG�$�F�
c��8u�!���3i�}I#FA"C� �L6q!�Y�;C��qb����ְ{�J1i!�$	;,wꔸȓ6�h��ꇲK!��	X��a(pG֊s���j��!�d�%���hãa@F�8C�	�/�!��F��7�D�I�h[����J�!�E!uZƅ� /R�[�JixĤ�8y�!�d	#q�Mz�/Xi�x���L�!�M�� �8��Kc^�����&W!�M�2����ұ@��Q�R�(M!��m4ҥxP�1=�^ț�)�-%>!�DE����r�[- �HPƨ3)�!�$�)h�
Y��苇q{�F��[!�$�X@��q��M����KҶm�!�J�8I�@�!D��s������(�!�Dۍv��}�).=q�`^�H�!��Eg�dѳ��L}�`x� �Y�!�DA&�`�h�5JQ��@�m�!��G(�D�У�ٻl&>\��fݡNK!�$�=%��1��(��	�"O�I��  v;�d� [$�ެ�#"O2��6Ɛ�$��#Rb�60�`�V"O��P���iP$Q�r��.�fC@"ObY;ҋ��t��/�i���a"OJ��P��w�V���c��A�8�i�"O.�xBL�)i4�}QRc�,;�t���"O��(��B����:��Ĳ0"O�1�C�0���ւ�M�By�"O�� �H��<`^���o\5i�����"Or��f�N!z�D�gϐ�=��%"O��5$�;f��nң'����"O!��I�!ϴ��.3rh�:D"Op�
��߼J��<K�͗�y�"�u"O�3R`6A�ڝ�������"O͋�%H� {�j��żd*Q�&"O�AAI�:}:Q"g�ӥ����"O�Ё��)�&q���^�k��p�p"O��"�məf�ԭ9uM��+D����ݲ'�`1�I�<J�^D�h,D�� n$�����:�И��M.4
(w"O>�(��!�H�IE�P=��P"O�Իc���f߸a�g�
�u"�(�"O.�j�'a���D��cjA�"O,�( �*+��Mxc҈a�x��"O�af�\Y����ҡ�J��"O���B� �VRZ�c�& �}Hs"O~�U�J�!��BBc�9���b�"O��!&�J �F���5ٺ�Jw"O��)��6��``�+��!�d"O�Q(MTg�A�T���f"O��dL̐S��X�m��n��ٳ"ODhI5��t�hTa�N�Lh���"O��B�E4#��F/�2��B"O.�+G"M1jP�
�늵b1����"Oj�@�m$52D��AS�/$�X�""O89ysߏ��y�D/�8|�R`�c"O����G�.��l��@�S��(�c"O��	%Z<8�ja��֨%����Q"O �YP�QH��dڱ���z�T*Q"O�)��e��I�i	b _�N���V"O�$KfE��,��%���D.^8�u"O}�@���-��V�:s�
1�ѣ�g�<�1���a*����E3�)�S��}�<�A���[���2Ѡ	���|#�d
w�<t	VY��`B�V�m��1�t�<ac��v����g�?ߞC�aOG�<!V#�9T4�	�7�@>i�x��D_F�<�""�%T�i��� j�
�C�<qT�^�.��S�OH����G�A�<A�a�}���yU��d�,ܪ�~�<)d#���7- M�Z�^h$��1ȈC�bA'Ce�H�f/3AvP��2ɎD�_Cb�a,U&A�԰��`5pDj��BkB	��'�q�"ɆȓYU6�h��K�P���l�?�ځ��ihm�_�
Ԓ�2`B\�%=����!;�!�s�R8SQ�a�ĽM�&M��q u"d�Fe�������%;�b���O�u�&�CR�<�t�����t�ȓYxP�	��N�	�����d�ḣ�1o�k�sR���K��;a��N�-�=j� ��GC.���,��'��]N�#5�֊@a���>pdm�`&%���*@�N������~,�#
{2����?(�6l��y�i�D�ˡ,F���PK2�m�ȓd7$�c� B�o�0z�J&td؅ȓz��M㵮
�Yz�%��|���ȓ0 i���(ej���(�
s���]y8��Fn;�8�#���~Bl��ȓB��sf[$Th��3CхQ�\�ȓ|�ԭ�U� "�M�e���l���K�FM����X�i[�	�p^��ȓy"��נ^Us"	�u�ۑ>�V|�ȓy�&��/Ѕm̆��îȋI恆ȓ����EL�p��l���q7����v�s�G5�� C,�=2�=�ȓ
L ��G�O�<��;f�х�UI��ې-\(V�&uC懶�bą��j�櫐7so�/	d~����7D�02U-� =�vDIGg�iLP��`�1D�ȩc�I�(��2��=-��xPb.+D�q��	z�(��-��9�=��,D�� �@��k��7zZ���ϱ�<�8�"O�(�@]S
plIv�#Y��4a�"O�1kv��lo�,��jX�3�ܴɑ"O`!����3,�0W�G]�1!�"OM�TDW9�Pu A��M1Pڡ"O��De�y*n*(���"O$�y@	�p�NI�nݘs6ĽC"Ox}���|�P)�C�=,�b"O��	�	�1:��0'�څ7���B"O@��ň�<K(�z+ȑ/�ֱ3�"O@��s��k�� ��U�s"OȑQ#�YQ���g�ʵ.��a��"O��pDgF���SqGL�+=1"O�����9j��<���k�"O<0swc��~��3D*��Ej�PF"O�))��F�%�|p�蚙kTx�W"O�@BG*6�0�3ȕ�eGֽ�"O�T{���)r�`'ŷHͤ� �"O�51C��f�6ԃ�,@�x D�R�"O��Ѓk�(�t��ᅿ:��X�"OH��T6���o�J����&"O� �©M!ns��ږ���JLj�"O~���ə?2!�#��6c8��c"O�h���REؤ��w�P:MP:�k�"O$����cc�q�Pf�-4��Y;0"O��Xw.Z�F�,��pJ��"���r"O�����L�QPc	��n���9�"O��s�R-	Ř(ӊ��Nl&�Sg"Oxbṕt�5Rb�Q.5U,��"O�P$S�.B����
KgM6%*&"O�������Z��K�A4*�q1"O�-�E,ZS�pZF�9>-�MҀ"O�dC�]+)��p��`׍rfq�"O�̻�O�*�Ĉ�CS�0�,
u"OH�s����,3b�.+.��"O(QSMF�i�fQC�`��F�r�"O@A�P�
�PQRQ���0~\��9a"O����ĮK"Pԫ��5:Ԉ�"O���������,�1o4*E��"O�8��Y� �L�a�Mz"F�X�"O�� Ƌ�7�9� �ц�<Ę�"O�i;�O�WN����F�{�!��"O���%
�O>��Es�J��p"Oz�@,��,Ihd�Uf��,*8�1"OL�1�N�i%�1!�Ͱz�Y�"O��[�[�/2��[�-�|�Y��'' �}
� �- ��9)��8�)+D������
*b]���P�`�,D�(�j�Jv��j�U93��*D��Ҡ���%����(@?�Xha.$D�t�S�F�Vh!0狊-�����$D���c�K�e�8�� (���*b�?D����Z�<EX���ӜQ�JIZg3D��q�[�Q��`9gE�v���t�/D�p�0��&)��q��U^i�c"D��	5�H�_���@���D�� +D�(��EQ�ɫ�*�1.Hh;2 ,D�d*��l"�ّg�g���ׂ(D�U�`��aZ�υ��.�E%D�L��^�e����h"A�&�#D��2U�^L�iB��ZT�Q��5D����������wq !��&D�$Rb%�Q����D�����*%D��c�"�i���"fѼ��(8� D�� �A`Ɉ�\^�C'
�9����"O!�!ӐΌ��`݃)BA�"OZU�S�M�z�V8QD`P�"F��c"O���Chʔ`Ѿ��t��U0��3U"O(�iE��&�a�A���G8���"Oڸ��K$
(~�a��+K�����"OȠ;�"ɫ7��)"��	@@ x�"O����bѧ\p2�S�D��{�r@��"OV�;�ڹG"�Y���_� ��"O�<A�e�`8`�B��/S�$�@�"O@��p���8h^��3�)e���iV"O]�ᄆMA&�@��=��qav"O�m��\.-6mb��(>Gp-Q7"OH�(�+*]O�U��*C�^3P10"OT�u�̉Y�,�{�(F5{��q	�"O�H�'�یU*�	�f�J-%{R̀"OFQE��T=� Krf�-���p�"O� ԋ��&7��9���"T��˱"O`)��E�l^R�A��~�l�5"OR��5��$4�<����X7h�4��s"OܵR���2X��!0m�>-����"O(�3��q�V\"Q�ܫ#�nPh�"OZ�AܾR*"v��;g"On�BU����u0"Rvxl!�d"O�	z�F�K�A둦�\vp%ku"OR�k@�ϳL����#�H,
v��y�"O��
&fN�S�Ĝ����>7��{�"O,ppR�v�Ѐ$�<1)��"OX� �H�d)�X*a��A!D4q�"O8�u��$*lN�2#��@uv���"O�݉���<U֮���2�-P"O�a ��՚Ԁ�+�8]�3"O �����<� ZbΕ�m���Q"OFI��fҴ?����R�O.N�4|��"OR�Y!MD�TYV�;$�\&�rA��"O�a���7��YX0/SR�(�"O�|� ��+�Dh�eMM1��͘�"O�<�!�Ō`��D	�k�'V���iV"OH���Vm�X�����_T��{�"O\�P�S�`6�����F}��"O� �D.{�*%����p�(�x#"Oѡa���\D��hp���4"O� ׋�R~�P$��3�l�)0"O����4�z�@%΄"Ly�@HU"O�Ի�Ҹ��0QF��pv�a"O`4& �9n�����P�y��h�"O��%�L =İUK���}����"O�%(�B��#�6�� �ˬ2�D"O20/Dc����Հ��u)�"O�{����1֠�;d&�ʰzG"O6���\� t���+�Ⱥq"O��05�܎%Ef�[��\%v"O�e��ŀ(�R�8�*�4%ܞȹ�"O�\�3���j`�V���[��5kr"OfHi� ��-���	ǁW�I�48'"O��z�g��.�贸�/Q6r�֩�6"O@5�#�-s�v؈3G�q���ZV"O&X
��"5!�w�6l��e:5"O��ڧ��9�d�{ ���&n
`X�"O����CL�8:*�ItB�&w��P�"O��@�E⬼�&�!/�B��a"O��ԉ��H�5�K�x><飕"OȰ�a�/|(�$ǅ-Z8��`�"O>-y%�����Fڮ_-��"O� F�Aj02�P1"���i�8��"O��#Iʶa� e[�c��p"O��@�j�-/J�!@��Y��Y�"O��{��ʒZ�b�qC%�>9�R\(�"O \��i=(�h<;עܽw��ѱ1"O�L(���"��#GQ��P"OT��v��))f�xF�D�]��"O�`�0D�)�V(�g/ �\�	��"O�,�5j�Cdʄ2�i[��"O�0Q��ޣ[�*ԙ⋛��fѪ�"Oθ�5i��$ΐ��+߇M�xPf"OL����,P���P�]�(����6"O�dx�G��l�viR����@�"O�����.R��6j���w"O����G�sr^L��I��yu�MÑ"O@5"$����X:t�I�Ysꗤ�y"aƼg�PJ�GE����K�y��*p
�2u����p*D�=�y2���6pJEYS�ڪ �Z%J���y"�Z�;��ۃ$�,~P����埄�yRŎ2e�	[���r50m*��
�y��;u���􈒪j�4@K��y�/ՅrKb��V�J�x{�&A��y"
���t,=r��D��J��y2���{ir\x���h���mЭ�ybNP�!�؄:a�6����a � �yB�d��Qao�s�F��.���y��I=*��� b(:;2����M�y�h�s"��q(N�5�0a P C��y����[��=Qc>�FQ��(P�y��Y(:.{*��5D@M�@��y�ğ3">>������ȹjuf��y#ӳr�Z�c&�	&���1EE8�yb�VV���+�d�: m�o���y�M�*a���S�G�K�Bx�����yB��aF����g߭I��zc�_��yrM�"�x=+T�ӑ1+|5�R)F��y��+�>,�5�T�`��bd@��ym��R���3�Ř8 H�`��5�y�$ɗ�Ug���f����J���B�I�匁���
P����D�C|7�C�I�	��ր�j�؜�j�*W�C�	,Qܬes�,ơJ�r(R�"ϲL��B�I.	�4+_�h�^��	s� !/��H؞x�2��8����%`��óF.D�<[��M����f�,I�0C��,D�X���F�>�B��~6�L�t�+D�P+��*v���*TួS ���rh<D�Л��\��� k�U��@0D��;�ҷ`vȱS�W*`3ҍ@2�0D���3��(>Ժ�
TT>n�����-D�(s$���k�FQc1�������)D�Zs&�"RbV)	���k<�@��:D���#�_2k&(,C������� d5D�XK�c�u8�F�8��0[%�3D��X�^("�Ҭ!B��!G��X;��-D�HÀ�z&��f�.-��"�*D�8�S��$(��tHD>o\TkR .D��ȧ�M%�&8	�%�r�:����?D��CD�XH��0�M�J\���"D�tS���b�P��,ЫY�(h8F D�����G���'a��MR��0c=D��a�K
�v9�#,��9���CE:D�	C�@�IDH�� �(�ڀYba8D�� 8��G+�:?�1�a��joB� c"OD����%S��y�@/��oF!�"O�:�⏘�\��%�Ź+[��"OZ�p5��'y�fy�ӆL)�M��"O�����0��\��Յ$:ԙ��_�x��	�TYP%3D�� Tσ�P�xC� pg��)P��\}^$zC��1T�@C�ɘT{n�X��_�m�Z��E��j�dB��w�P�i,-��Y��F'5�$B�ɗCwj<i��M*g�2Ahv�P8'C�B�ɴh��1��N�6�I�bɒe��C�I,Q}N��D��FȶDjD�T0�BB�ɣ�2i�∙-�|`h�ř2$�C䉙$�D��KX$FNHHy�d ���C�	�4�t1�,7- $R��Ȟs6C䉤΄S'�4o2�1�)��&#�C��1
W@�C��]j�)U��h�$B䉮F���`�_�,���!E�x�dC��X�JI��[�-��C4_GC䉻U��<��)�\�(d "Y\�"=	�c��<z!��
y�z���F%~�q�ȓGXP8p3.��� L]� ��ȓIe���@S81j�H� Kםv�v���a�8�hDll�$�scDK�,1Fh�ȓe��z1�x�<�
BA��}n!�d���p� rlL�8�J] 5Z�!�9.8��m�� �̍�]X!�&Ct�Z���A�� cPe�?MR!��M$�������� �m˾3P!��u�>+�U�t((Ҭ	�r0!��^2��S��M*�ic����Q(!�$��k��Mp�'�jI�Ի
�W��z�D������2��5�e��3�!�$��lb�҅�6���i���	�!��N2x
����/V~�D�uƙ�=6!�ğ�lkt��� �yr�C����!�$�=a���Bfı3i����
�p
!�$�"I8b��A�E�HI���j�y�!�d�3bF��3�(F��h��oa|�|c��9�>8��J�?5����͇�y�6/�8��G)�� �!�C+��'Iў�O;v��s��\�+P���`Q����'g* 0HN�qu�Aw�ǡmd��'�����"ÓWM�I�VJ̎��u�'��%��
��t2�H���m�J>��IJ����j?�]���F="2ԅ�*��$�7w\H�c���ީ��$ɮ i�� {&T,�V�[T�UV�<���0�	B	����⢝O�<�k��Tr���g�Q� ��&T�𲒄�)DB�0�(,���!en!D�h�$�N����CV�?� �E)3D��!D �K�����@����%D�P�*�&���B�ȃ�m��з�"D�Tˢ/P�h&���	�)8i��W�&D�X�C�6s�p3'�ރc�v=e�"D���/�>O��c)��`����� D�d���	!B6P�Sc�#R�8Ӂ�9D���)��1s�4�E� 蚨�&�5D��!�/��U�b�@LMx$�b &D�hx�	�%F�� C�{�hAQ�>D�\ DȒh��(r�L��� 8D�Ī�KɚD�8[�_#X�l`�O7D��!�hH�T8\9��M�b���#:D�� �8����e�Z4{�DK�c(J�K`"O)S��@%Q]Nh�BZ�3����"O��@��)�� R"��!���h�"O����"S�2삵b�*�Xy��"Oj$�%\� &��檄�h��q��"O��*7lI~H��K�', ��'"OD��A
B[S<�Ch�Oc�l��"O�jG�{J�H�5	�GD���`"O>՛���"(,�√�;<�a#@"O�E��J�nA��Q�A�
;�a0!"O��k�*)��1o��D$��s"�M8��c�ρ�#�~Ģ�Ț�'$,ȳ#�$D�T�I")��#� GV"0B�)!D�(�8/@x������ D�aR��4Z&�%�Q��<5g����(D�`�E 	{L�����ըpL�8��H2D�(HDmֿJ�l����,C�ěw 2D��ڶm-D������tQ�*D�$�4l�!)�sA&҈9���1))D��15�6}&�X�.��p�,��(D�4��·���4�G�9��%r�J%D���m�>p�<3��m���{��$D��H�i�>V���Kw�*�$\��c!D��*d���`���GO���h"BM$D���A-I�ބ��@�Jt����.D�� Aߐ"N��B'x�d�:��-D��g��=��JA!65D<q,-D�x!G�����bҪ݆%yPs&-D��X#N�)�0ir�*"06q��,D�$� �U��iy�/�	8<�P��=D�LYA�NwV��$�&�E�4E8D��"d�[�y����ɖ2[k0�%8D��@�W�}��S'� /ԅ{��7D��)�3?j�)���C�����M4D������
�X���I��H)�1D��CAG�X�r4�cD%)��P��O1D�4 ra�n��}x�g��b�(±�-D�����J$kH2�:E��@|�)7D�|�'n��]�M�q@�FZX�h3D���T���Zdx+(G�Ec0D��[�U�cR5�v�6�$d���:D�(��Ýfv4�(ш��k�2Q���-D��[0d�'r��Qɇ��<%�7D�8b��ķN%P<Ȧkҝ^  �:S�/D���f�
��F)ԊJw�h� �#D����1+����� U�4�d� D��tn�b�<�"뗋1��K�G*D�����äB�Q �,�"��6D(D�(BwK�6�d=��$�W�d�'�)D���,M/�vA��E[��t����4D��1 �4f�a(����O��9W-3D���7NJ�AfH�i���,�P5��%1D��JE��v_�dJ�`� B�	�3�$D�P�n�*�Ȁ���A�[�!D�t�[m��t�\0���xcЌ�y�b�>SO	HdE�/���yD��#�y��
?-��,�d��|d�
6�y"G-�DK�F��^<X k��yB�NCH��R��GQ�r�����y�Ã3EĬOJ�,�"���yb�[1ḿ!�&�2gv
0���W��yb����O��iJ�Y������m�	�',m�#�U}`�a#�(&�r|B	�'�	b@��6ov�:3�I5A?���	��� �!�R�߅W9v [CF҈<��I�4"O�\٣��
D<�� �ɗ6�T�HQ"O.�dfss�p�W�E�r<�K�"O@��TE�}�༺g��[p�X@�"O�2r�B�!|�ph��A�~V E"O�0�¶N;>U��"�j)P�h�"O��b�(�\�p�
���ۄ"O̤aǄY�:`�E��@���H�"O����)c(>�4n�~�x��a"OZ��X?6�h�H���#U���K�"O��q��	��0�t�	�
��BT"O�3���� �dS�Bn�x`"O{p�V�h�V$�����N����"O�]�4L��	V]) a��ON��x�"Ov!�Q���8��� �K����"O�4¢Y&���:���)z�6Ě�"O�1��ϔHZ�JP��*J��*�"O(��c%�&�!��)~L��"O�}#�cHO��S. �f�0�"O��Z��
��p��n<*^P80"OnE*ŝ{��p�T5W��9�"O�|����&�^(R���j���"Oʀ��I�.�I����"���*�"O�Ҥ�RW���gK�u��Uy$"Oӓo�%I����ǉҙd�<9�"O
�:a��q�i�]�h@�"O$	YGIV�t�<�	jU~��d��"O`�J�yZ.��Q���(�H�p"OJ<�q�@���*b�ΪVv�U��"O�p+Y]6��p�l�n��pB"O4li��I!0	v@�6�_d���"O0��I�9[7 �9����Рk�"O&����!_���%W�h�=80"OH)��d��>i�@j�?A�M�`*Oz��H�2���Q�!3ow�<��'��a���"�&A���;i����'bv�ГjQ���!tE�ZMf���'vp�D�EDl�i�#��Q�t���'�9v��'gvݻ��:6����'bȈgj���������c��u�'0`���ןjzJ�b瀊U�@Ġ�'��T����7Q6|�ȡ-��J2���'�軡$��G9�*1��3Yl�'�@w�U�+:y�j�ZV�!:�'���@�$)�� ĿSr���'�F����b����!6�9��'�N�	���{���w�
�e���'��,��W�F���`ӹX���a	�'�(���Q�x ��8V C�PͶ���'+B�#NL,K�ޠ"v×# c��'΄�� B<�DkUm��l�x�'��,8S
4l��$�r�A�'�h���jԀ~��QBg�L�q̬��'@AJ��F��.�`�OÕ-깱�'|VT�s'K��-z���)y�	��'��)p��n�AH�aFJ����'9�}��l�1i��i��G kipt��'�2���03���*6@ϝc��Z�'l��Bf��N%�MG;Z�\��'�Ha9�F@ ����7���e�����'�����E�a�Ru�G�e��Qr�'N\pA7��e�&�12�#Vxд��'�\\ۡ�]����vy�Z�'v����P۪�"ȊC�}[��� ��Sj�&� %�a��b�I"O`I�!h�p�j�@*L?b�Q�"OXyӣ�ό:�����S�5N��G"O���b\�6`t���h�0&3�ػE"O�|i	B! �dś�$��ܑ"O�����(ݘ��-d�#�"O���&ɏ>�p����b��� c"O�E[��(wG��S�ś*�:�a1"O���j�/8�6��f����U	U"O��LA��X���Lv�ݺf"O��	5��"s M��h�>����"O�ࡢh$- �̸�'�?�l�"Op�#陴e����Źa��Y"Ov����\�&s������*`4�f"O�dJ�Fq����hL!3�|�!"O�tt� "�;��A6�ł�"O����nM/H�f=۔�]����"O�}�/��Lޡ9�d��H�j� "O�1�!K�0�F`����5J ��3"O:����U.w�
�)���V<��"O���M����PG	Ƈ@�^�8�"OU�ϡ�@q0���	q�-Y�"O�I����G_�QKR�#_���"OP��d��,v!��F��L�"OJ �Ç�Z��Y�cڐ �04�"OĄ{"KJ�+��B �I��鸠"O00�'͘:`�>@p�a�%�@�"O6��uđ�n׸uB�ٵAn`"O�T��S�q4�!ǠJ`D(�"O*4��%�FP
�Y9lL�С"O8��ƥ.l0P`�Ѝ�G��`IB"O�!�F�"=J�-T��N�y"O �!-�#b2D%Lнpj��*OH�"�A�vy02� 
/�F�z�'�lEa��'�@���7Ӥ�	�'�~�j��L�w��0��ܓ&ZJ0J�'�K2.�<.1� �\�&!̵��'j��y���-�(m��l�.~�	�'�8�{�^+QB�Q`b��)F(	�'%�&�
IT�l{&H�#��5��'�Uu'�>5�� ������1�'U�D3��DU �f�)0�z�'b�y�#���C�T�6d��b�'u���K�?R2�5���'��hJ�'���#@�S�E�����̣i�f��'8�$q4���%J�y	\�gʤ|a�'MH�N8�N���o^�'��yB�'w�t�լ^=S�3����|	A�'�X-"������8��ϳ����'�鳵jD�>Y6%S�a��EBLA
�''`\{�Μ�j�Z��P�~]x�*
�'��X ����Z܂%�	�qVT��'���R#(/X�J�@�V�xE��'[|	���|$�{�m� ����'!�!0#��iR���o	�b�ؑ�'�j=��������jK����*�'^��@ E��F�.�-y�N|�
�'l4��M1'����I8n�4���'�)��.��̬y'c,�VPR�' -��NO�:�Bӡc|��'���0%j ���$��BP��$�yBe�=Yb�*a앾Bk^�R�EJ�y�E(�i�� �9�x!��ύ�y�	QP�`Ic�+�Z�"�w�ė�y
� XL�u(Q�{u�H�c���p�1�"O������-~U�����}s�"O�p�ǃ�_�8Kg��P�� �"O��UT+M���#E�J�f"O� Y��ٚqRl�5��6j��S"O$��"�,^AT]ZSOT |�P|�@"Ol�r�!-��<���
+ÀP�W"O*܊�O�8O$�*�n��Ą��"OJ)*���n���qw�ԑ.�8ܲ�"O��'�#Jق�R#���"O�T��앍CV��AV4�ȴ��"O�����
6!V�9�7�Y=���Z "O�<�Z�E.{B]��e�dzja����X���+{|@9��_��汇ȓ��U�e �+z2�;����&&jp��@���TKM���-Cg�P� ���ȓ>��۔�C���xc�'(��0���iI��$(��F�߬<4�ȓp�0���j�&e��� �߽�M�ȓTL���"	�Z���@�2|�}�ȓn{x帒L�jJ���F�[�4�"��ȓ>�^�(�L3yҽ�g�1\GZi�ȓS�|�D�3�t���K�ea�Ѕȓ"�����\�5�x�YnL����X���6��>"�Դ��EI�n����X�vF�IU(g�� /R�ȓy�M*�Ϋ5*)�&��9zZ�̈́�l����d��ZG´l�
0�ȓs70  ��8@,����J0^�@����
���j��Kr�+��5a?�5�ȓELEs��Y�~hd�__�ԨJt"O"�Y�SՂ=�n�?!��S�"O`�I�F�Di��DU&��(J�"O`��m��Z,0��E��56@�(z�"Ob"6�Z&J�: ��-_���p"O���'�O�uQ�P�wi��W�|�Zu"O���..�����w宵Z�"O�y�a�ϟk[&`��(�:˴EP�"O8T�M/7"��pȐ�
��Q�"Oڔ���ή,���@��4�����"O��q/_:PZ �r���o��U�"OZ؊��.�	"@�3?����8O��O�d�<ͧ��'Ԣ���$Ϭxum1F�"C�6�:	�'�v�����/~@��F�Ű#��p��'�ak�Ě�	 �d��Gl� �'��sw�_���ɶ��>�r���'7t`���p#(���l�.>����'��ثV��*z�0��<_��x�'@8(kA+Ƥ�q� 	O\qB4�|bW�b>c�t��N��El���,��N��9�7�$D�xYb�Nx��m��X�}tҭ9�'D�8KRn2F?���U��3C��!(��#D��ƥ�gF���AT~p�9��!D�<`,��`��r�(J�@��J#D�<i�-��>j��ʢ@Z�Gryq��"D�T2��H2���F@E��@���$D��i#�ϴcq��3��Id���y�ɉ�6.|³a;9�:�y#nҧ�y��9��0�E(͠7��<QcHP�y��y� #�^/�n��e�J��y��"<�<1v�5Vk��+�@�y2�Չ ����Y�R*%+� ֕�y�.*���E�5�6���k&�yR�)�' Bx����:,�c�
U#���S�? &�@'A�%a_�\���^
p�#�"O��)�M�w:�aSKV�@��"O�)���Z�Z�4��磙�$�"O���]9� ��ǬY���o�[�<٤ς.n�Sk	�`?��r%
U�<	W��(CdLh�Ĕ�Wh�ʗ��R��h�	w��v"���J�&|�E�v�R�BiBC�ɷ)h`A�Δ?j����)P�f��B�8csdDh��WU���?�B�I>o�)�w�&'T�8���ڞЀB�	h@���
C�[_p���ݬX�B�*(s�mA9�<��@f[/'�C�I�,}~i��
"%�Xdi؎s�����O���K�,� Eb�a�-P'(���z֠(D���Q��=��D��B�|�Y��%D������P/�l���/�]8V $D��Q��ʺ�.��`ۛq�����>D��BeV��$�@�Nԍ�p��x�<IBR7�zݨG�|��[V�j�<�AL3�RxQ�h(4�"f@d��	ן��	�'��0j��T~D�Mr���9k�>C�ɬ�b�{�L�C����JÞV�C��R�T4�V��%1`��"��6-�B�I�Wn���� ��T��� n��H}�B䉶8!xz�k��� %	�~��B������g���:a�ڝt�|�hF"O��:B�RE�4ۤ�^6|(��'��:Ig0��F�H���bQ R5tC�M��`a$A_
n|���DC�	U�*%�5�\!k|Nd�BFK�,�C�ɭd��Tɰ�ݯ6��R�"�<q�"B��&;�$��E��A�ƴ�3���B�	*�P��!!��3���%�	��C�� �"��AI�ʼ�u�����C�:n�2m�S�@�3��6�C� f�4�P9l��p���4:�B䉰#T0D�[,$h �R�Wo�C�	'+`�)Ц_O��9���46_�C�	�(Xx��U� ��(�5�H�I��C䉥o}�Qy�N5��ˆbFp�r���2��F�AE��ہ�\sM�H34�X%e�!�d�,
k��R/N/ND*	2�\-x�!�$²:-r@��& �lqD�L��!�_(BRn|�-)JR��P0{f!�$=jÂ �``�� ��اE��)d!�H�!ڰ�5˟/.�@R�c�,D!�$V,1.*<��ңo�<!uaܴR�!򄚴�Ƽ*JB��h[�`��n!�@�JcP� �ⅇY^ �S��U!�u�"��ߕLH�bUH��q0!�$^9V&�hQE�1e�L�AZ8/!�dΚ;S����	/[|]��)Ua!򄀜w�t�qEGVe�n�J�G{!��/�\���	�	�N��e/8h�!�$�=aU(�Ӭ��a ��D�!�D��. e�@���Ҥj�ܥ6�!�D>	�r�B59w|;�kZ%-�!��$����/�rd��1!�$X
�  	@p��X��܁#�!�ě�D���)�i��@����L�!��}�`M�I
�
q�=�4�ĝ@�!򄊛5'������eXͩ�d�� ���A���d�|�d���n-� ��*eD)�!�K�y�K&;G"8�U4P���5����y
� L����R�+�Q�$@��h�����"Ob��ܴ��,1a�ád>H��"OT@ѥ]��Dȇ�X�Fa8�Ç"O�]�r��2hN���.4`���#"O��YĠ1J����a�E�]E����"O�TQ��d[��'u�����"OB�B���Np�˧�Er�E�p"O�|��\��p"�▧f��5"O��ѡW�l���[�a��E"O��a�Ai��XW�E-M�� �"OH@�tL�-S�҉�H/t���#c"O�m1�F�=Q���^�p@:�@>�yb'�'� <��蕪4�l�����>�y��ѱ#�jl8uk��,Ip��S.�7�y�݇0[$]�����_��Qs�
�y�&�Άq
�`����Lx%�>�yr�nl4Ɂ��!p��U�匮�yRA_.nm�UygI�4�
�T���yR�V4-d���čQ3n~a�#+��Oz�=�O��Q7♽}�.��sB�%+��q{	�'L�|�"��{Є�PT��Lc����'�Ժ�Iw�����Y���(�',�� V�r�>�����%�b	�	�'�9� NW�k�npC O����Xz	�'��M�`�I{kz���fE�)B�y	�'VZ�QeGE?�9�G.͢t���	�'�0	�΀�0���`���"v��k	�'Zx3�a�2j{~���!@���	�'��yB��-����F�?%p���'�X<����>i�0ТqӇDU|A`�'�T�2B�[��Vє;N2��+=D��$�����<r�!��ga�Q���;D�8x�D�=O
	��(R.wd�%1��9D�<*A�!<I��I ��N����b;D��)F)Y�e�6�k`��	=h���(&D����G��d�rٱv�T�(]���&#D�p�ѣS4m{J<��eM'�й2ţ D��QG�Ar���k�.�$��!,D�h80�ޮ"�m�F��2ĺ�d+D�̱LV�xk�y(4�Ĝ� ��t�%?���ᓍc����Aj[�r 1b��@)jB�I	D��vL'<dʔ�a"��KDLB�I0��@�I�7n���p2m@ '�C�IsՀ i&n�a8��ݓ{n�C�	%G񤍹��-L��*�Z���C䉌Z��	 ˍ�e�p��`G_C��e���v�ޤ]�$eQ��ٮ}/�B��#�6�ST��!ZZ��u��B�ɣK��Q��X�T���Q
׬F��B䉣z��]PO�4C��8R(�j�@B�ɫgj�"���.a������X6OG�B�	m�n(C)ȫ{}x�ʣ�@�j��B�ɲ!w��@���sP��U�	#sTB䉺��)���)��A�L�?�FB�	8%����:�*��6M�C�*B�	?p��Ř�
�������B�	!b� I3v�ܸL���Nk��C�	�2�n�"��޺[E0@��l��_��C�ɿ.�!a�(5s����!]�\&B�	D��} �ȃh0��Ԃ�4)i�C�	�l+����D�
M�p�@��	o�NB��e9��xl��N�t�ӷl�!I�(B����%
U��68���I�.qB䉕DR ��V�\�	��!L�:*�C�)� �8z����&.�9���"�"O�!���X�0JVYy6��Qzxlq�"On�h���I��Ĳ��"Id)��"O�;��SYz��0������� "OtD;c(	�T��99珄�sq���"O�(*�E�R��XT$ߒgn�(S�"Ov\�16~l����D�k���hD"O�|;�̟�Z|d�Ա�:��'"O<L�5,�� C#�Ï��Mɣ"Ot<�B����}�&��*4�`a3�"O��C ��0��T�R#��A���"Oe�C��),�գRQΩrs"O�,36��"H��Ï/`�N���"O>����א0�t�Ht�S8s��aS"O.����
	�r0r��Jll����"O��b��Uf �sGm�*~g<�Q"O�<��k��B)�4I�Han<��"O^��Gc�8XAj\ ���
��'��Oĩ�N)nt-��f�.�r$��"O�3��(w��T��n�f���"O(Q��W�T2-aeeW#P�
xC�"Oh-X�䌛��y!'�Ə{���Bt"O*�{@ϝ�tRތx�K�-�䱢�"O�"smĹR�.�[��C�@�k�"O�5�$��)xl�H�7o�w��H��"O��*!ꗋg4�����T���G"O��)�-��qC�YҖ"�T��"O �LP	�-�х ��Ɂ�"O�!�D��i���1U՝?cn���"Op� �'N�Hu���V`=��"O��sÔn08���nя?G"Q�1"O �P憝��TpQ�_A!��0"O��1�+�=���bO��C��P�G"OV[�KZ�'O�ciT/Y��@'"O��QAOȅ/q��8`�]<����"Oʬ��E܄� @X�h��e�q"Oz��&J�j��x�F�d��	"O����ƁF`�EP'&J=QM�|�"O����0 ��Y���2>7� ��"O��i�Eǧ=:6-�eA �Qc0"OVm"��t�b�DH�ʑ;"O���P�G�QZ"�jӉդ@Y��X"O(�2�m�-b�D�D�:?r����"Ob�J���2G�Nq�g�7x?�!"O����;T֖\�"�
� 0޽k0"O���vl �0d�1���OD��"Oh9��������ꉇ^k�[�"O�X뷏�/+�i�� *.f��R"O�Cա_>?RBI�S�R�2��DYg"O��*6�G�n���u�28]�p"OX "T��'{R(SeOQ1q���x"Ot�x!�P7'kF�AD�F.�xly"OH$[��<-�R	"'U�H�z�9�"OT�㣊�h	��f��s�8�"�"O6xuH�#
�|��&^�X��"Ot�B2���b� `��]84H�a"O�@�ӨX�-L|�DC�.���E"Obm��!X�9[�a�$�?�P�R"O����nF�`�p��㏨Y����"O�XK�M�S  %��4�˔"O��{Bk�^g��R��a��H^4�!��3p1�oA�TqS�R�!��_tP0���ǟc�|�cJ�0�!�U�N3D��j��=@��T$%�!�� YQD�?-zDi��B'"O�yuA@���c�ҟwh���E"O���D|q4lp����[��Ô"O.=��*�.9�|$�T35>�}��"O�8��D�{"(Uɴ�V�3t��"O� ����o6]�1aۋS#��s�"O$����Se<(�h��P���)�"O������;G�XY2-_>lx("O�$p�hǈhen��֋̎7O,�R�"O�=:!�X.�3�LG*/J�}!D"O�U����6-ʘ "O�8۷aώ�J	���Q	6���"O����AԓwGr�C g�`�x	"O�=Q2g�3�&5�qo^�;��)�@"O&a��۹-�����5��&"O>�(�o�F��Ds�-_���h��"OL%k�/�E4�,�7K�5@��g"O&	�牞�l�v8x�j�!L���R�"O�`)��d��ič��a"O&�ʣ!C`t$ԁ��ہs����"O<�"e�L&3@����Ap�bX�"O*I��/рxa>9Y"��gw�q�"O.�!B�$F�Z�5�ޟh�5"O���F�ߙ*"Pp�c�]�Ūs"OBEKT�ga,ͫ�  D�lm*D� ��޹(��Cd,��E�l�Y4@6D��3�:/T�+r��ttN�Y5D�D �	Ǧp̓�� �"0�j2D��Pg"O�/�t�h5Ǟ�D�T�5l1D�����04E�U��Y58�c+D������6P$&��O�5X|�ȃ2�>D���`�#g��8 DӨU�|A`�;D�`�4oֿ~��o�wy��*M8D�p� ���AD�-ȇŘ�**v<ۧ�2D���3�N	2�Ը��=M��9gm1D��)�*�.Z�" ����V����+D�HJsN�
o��t�	5��x�a&D����)�3Ɩ\H���<|�l�9Q&$D���d����C�I�^�(!D�T�Ԋ�-�4�5�ʬ2�j3�B D�x)��G�x��1@F	��C,rYK�a+D�T�3��3n,ڐ��:!�@Q�.+D���h�7��!YC�bMaPD&D��:�*��@tȡ#�玼b��!y��#D��HZ�*�&!�OI8-:�U�S�"D�Xs��U��^5B"��=p�ΰ��?D�̑D���x����n'd�Xo<D����޳��M�M���	�#�цȓ�U��Հ#�VuBa�]5l�4���"O<D���LJ�n��3�~�s"OJ(b5���5 ����d�P�ڦ"OvĪJ71�D9Is+V� �(c�"O�,Cˈ7X}XI�*�&I#���"Oj� �C�	;B`�*ȘM�ȃ"O\ Y7*��E�r9y����0�"O� N�I�ix���+(FhB@"Op
�l�%/2R5
煗	���U"O�p���,�T�
�����"O�	CƆ@��0���.ҙrK�M�"O�(���!�6#t0�"T"O�����,�x���
*��"O���M��C��q��N:x*za��"O q�bȚ
	%����S����"O�����3!��݃5 ��bkx�G"O� ��Q*L[F�AQ�L�=U""O�	j Q#Y��ԋ�c�(%�c��5ړ��&��	�A%��4%5�ab��a8Ȭ�ȓ},^�r"T�l�x�aΊ��a�ȓ	�T�W.�j�� �˄2"��ȓh}r�����S`�34���=����5�Qi�48�T3Q���h�Ą�R���*C
��	��j�(8i�0X�ȓN]:Q�D�ZWrQ@n��tr���ȓxn0�3a3�����R5 t8]�ȓv⡒�#��']L��Q4U8����k�S�F[=�$��ǱL�u�ȓ_
���o,\�����MP� �ȓ����G�#VzX�I;򠥄�M�0IG�ˈ:�YqM����%�ȓC�<�;���49M�5���S�ЩFx��'ڌ=�gOZ:*���S���Xrl��'^�4#� �1u�|�9�L3�����'hJ�X���
N Z��V��'��Ƀ`�� +x��Α�L�	�'Vv��R��r|XxK񡍗�Z@�	�'㖨5䒃/X�M� �Șm��'c��r"oV JM	�'�+͢	
#�)��<I��P���5�gB�zYD�W*X�<�i�
\ܜ#$��."kL���m�V�<Q�#P$h��k��3d��h�$T�<yAɈ%�ૢ圢`��1���R�<ip��dF��e_:k�ΝqGXh�<At�؎>ފ��j�8;N��B�b�|�'��C�HKTnނ@��!�$b�(�y��|�'g�ʧE+���&�Y�*�L�ib�ж%�H	̓��?	�T�Q��D��#��`J�K��F�<pmE�H�F|��O�(ʒa�qJ��<�r��Q� ��m��Z%V�	0Av�<����'Z���.T/bqp4���Mn�<'h9^�E�%�;2�����h�<��'��`���H���k��[���g�<��a[�V�|�Z"���^��ըLg�<��̟~��Da�T�b��i�'�b���'��py⁞�'`]��NB812mZ�ń�h ��	8x��']б�"�5)�!�DO�&6he
��8�]�2kZ+=�!��H�R������5jײ�!���9#�b�9�iz"4`jY�n���=ͧ�hO)���^B���e� a�Ҹ Q"O<���6e���㟖 �RE��"O>hb�Um=��BE�yj*������D{��I��G�4�[b�9U'�� f�LJ�!��ӐE�2��K�~ �%��j��g�!��n�a���7u&��r�('$�az��D��	�T4S�
R�^BY�FҢL�1O�=1M>q��W0G*�g�Nr*2�e�<'b)Zh��k���rn	��(�d̓���<a.��ʧ'�MX�)�{��a��	 '��u��c".L�fZT��@pdˇK�r��ȓ<p����ɜO-�u�Ҋ	+���ȓ�݉w�;�(����ne�a�ȓ?\$�;�@��I�:xb#B@:A��0��T�H�7�AE�"
��ȓE	��H.#�<�8E���pd�]��/�������8<�RDs����<����	I����� G���D��-n^!�䒊k�F�02�:
 ���ŇU�!�d��H��ʨ���<8	!�� �F��"��x���/�~��v"O�� �흔P��Q�lE-H�Y��"O���w���l��U�U�n��͋��<�)O��'��i)��y���:G�����<_�x�O�=�|�sb���%gn��
����c�u�<��$�+~}ၠ�8u\��Ro�<ife�B����O���4��-ZV�<�QL�!,.����`���n�f�<� �o�]۶o�4]N���&��x��ɢhUt���7��<rr"�"/�B�I �B9�A.z`r�͑#M����y�D��S�O��$�R`�:��(G�N�6���'X(�c�H� dY�
�Z�Ƹ��')��$J0�R��F��S~��'ڊ]�@E*=yd a*��?���A�y���h��"�����k� ��#�hZ�~X�Y�?�S���Dǈ$�r�����6�(h�i�u{�ȕ'_�I\����ppr-��aƅ8�l\%ድg��	3t��"<��'�X�nӐ��3���s�<��*E���`�➹i�d�H�<B�Ǖ�����5x�s@�C�<�T��IZ<:���MF�E�t�X
�hO�i�O�� ����2r�r,�@
D�&k���e�\&�8������Y�>�R�� �2�H�FOE�c�!�Ĉ(@j�c�ƏԎt	G� P!�dȶ[rj�zAi&�brr��`Y!�$S!`����	��p1��@(4!�dE�.M���l@�r
���CG<F/!��sCn��DD&�F���ޤf�a||�˜�K;R��n��l�!@Q���yBJ	)k�v�{ފ܊���4ɘ'��Izy�Q>=�	���{UM��s��[�	 \)qa#o�'���>v*L��f��n�`�A,"M�B�I-Yj�Y��$��Qj���S��B�I�?B���p�\��Ö�(D^B�	��Zd�U�+��U��mqV5+"c���?�M~*I~� ��(k>� N ;t�M�7��<�	��X/�i�N��K��U#@lQ:XT�4���?Ap&ڽ~�8v�޸7��I���o�<q�ٲM($1dbV�T�B)��k�<��F��+ d��S$Ӄ"����%��m�<1��� �dL��=��8�o�f�l%�<hk&+<< O�qi�I�t�5D�@)p�>Y����<<n9�J3D�@QFM:?cU���E�Z��}�7%.D���)O�%c��@�b��9��-D�虣�( <H����a��$�f>D��Be�p]���qbÒ.���+F- D�2R��3}�c5E �R<��"�=D�L���U���L30A��*��H`Di=D�TB��i���q-�68'��]pC�Io0�x9'�a� KTC�(WL�C�t�dqiw�E�@�6a�Bシt�,#<)���?i�i.HJQ�g�
bqCk6D�D+Tj�r���"��� ��1	7f9D���@��=aP��X��ͤ[�ر �8D���r!y������<��)�K7D�DIѭ֍wL��B�-5=v�ۡ$4�O��/�`t ���~#(���F(�4i��4�x�H� "f��J�CCy<B�ɥ/sܬ�q 6Y5 ��4��y[`B�II��X��R%'��a@wC
+��B�	�H��]��n��@�)��B�3 �����<�c�D\����Sn���\��hOH�O� ��i��B�0r�FԐje�)�S��y�"E'(}ά���D����Z�y��07M�h�`G)@�<��S�8�yB�Ŵ�Nl81���r1��A���y�&Ƹ0�������{0P!�y"I�V��i�Ą_zX��R�ӣ�yr�X�p ���$��3`�ƹPA:�y�dK.���wmV7IH``qO��y���j$z�XOɵ=M&ȸC� 3�yR�M�KA�(����h���G](�y#�`��	�$c�4`��ڂE׭�y��RaG�ݚe�T<J=�b�G��y�CU>LuȠ��V+v����!ǘ�yb!Ƞ34�-9g:$��a�5kN��O���Ư4#hՁ2)O�|T�0�ȓ'4�!(s(�A1�:���+{���+��F�[�	Ď�!�GI'R����9���cè�>V�α�PJ� W�Xu�ȓ~s``ѥK�	t:��as.۝(��M�ȓ!� �K� 77�=ƅ�5$Ԇȓ%p�`+!Q @J�����{�|�<�	�W<,��Ĵ
�X��k_-�2p�'���'%&� `,[:lkR���F�\���'6D�3LKa�5	N�g�9�'���ѩyC�D�A��e.�0�	�'���ٔ��B!DY72ڴ�z
�'-"-���7��A��O;#8�[�'��1q���Qhcw�܂c~����'���3O<xH��"vkԒ[�\���yB�'d�i>��I�I�(+ ʔ2q>Q�0d.T�l20F��0��Y�5$Te��\Җ"O��k��R6(&~���c�4;%ҩ�"O%i�O	i�(��ԕW�Ɋ`"O��7+��rT�{ W�N�b��e�'��	:���0J�����7�ػ
��C�I�k�4����Uz|���Az���>yU�X�\��`��� y�� '��<ш��`ŌI)%�ۉL�����b����$8��	J����刘�&����G�U#c��C�	4��R�mD�9"��ԘV��C�ɣX��E)�aUK�2q2���$Q�C�	1����dU� �-��kǼN8B��5F�jL�B���C�I+l�Z,�% Z�C��Q
%cî!$�C䉰d�Q6)?V��m!�*C�5HtC�Id����K�'�tPF�_R@C�I8F ��Q��	�|�(B)_<w08C䉈[z���Hǎ���QrB_�d%�C�	�9�8$J�SG�m��݄vb�C剴G�䝳E	���
<8�N�<F!�L�~��I��O�Jx��E?KD!�Ⱦm\ l벌�3��!#�E&!�dU�1h%:v��m:*�q��~m!�d3+��|e�0�:����1t�!��	7r�� GK;(�+s� W�!��[w�4���P�)iç '�!�$�"��)��-�Cv�Ĺ�c�J�<A���^��E�ڏ`��8�3`�M�<��͚�|��S�C�8۔x��F�M�<���4AZ��C����n�e!1
u�<ID�_����nM�F�^8�%hB{�<���I�H�Y7@�#0n�J$CL�<�*̝)jJ5#��
#h\�u��)��<i�f�=G
(�̏m�`M��#�A�<� 2U��N���1��W!�6��"O¤�3�#�p��`�� :���"O�l�.=GRйJ��}+�4�G"OX�S��5h���s,�$&�0��"O�]��ڬո�sj/R�%P"O0�i6�+�y�H�
R��"O�]��'+_��g
�%Q4T�"O��1*M�3� ���ȳBh�#d"O4؊RlJ�4�h�q�ـ?Q6���"O���1.�46ld!*"ۢ%��"O�ѣ�ؓ'�����-���L��'"O ��+�}�|�aP�	l.|i:�"O�A�ֵ`b|h"�*�g"O�-�*B, ��4�ď��5"��"O�,�W�2<m9�GόE��C�"Ot�����(?��Ǎ�,|s7"O�H�`I��5]P�����@���
�"O�T:�)u���U���0n��4"OȤzӊӞ1��}��h����zS"OR��莇+H�Be�.8��X{w"O��4o��_2\�6FޏykT�4"O��� ����9���'o<`P��"O�X[���?	JD�e#0�|��"O� eDޮ#D�0*"a$W��rq"O��9��P����i�f��j�|�C"OT�h���� �0�+�ӹU�z`#�"O�h�Jש�����n��(�dYg"O�S�U����r���}�`<�!"O(�hT!
'�졨����QJ���"O��i�:=�bH�oW�+j$��"O4ps���(|������"P��#"Of�;$Z"^WV�T�-8�l�r"O��Cs�*B��t���G.Lwt�@"O���%���xY^��#lλuk*A�"Ox�;$ �*}����g`�V[L,
"OBi��n`���`�E��z��"O�hiv-΍2���w�C�"ϨX��"O����㇕GW�(�7O�*em*�Z"O~	����CV�!�cոE?��	r"O>�i�"ݽ|������ؼ#�͙�"O��@�Z�A���D�@�"O�0�� �9�`���'{�����"OJM0!�Ɖ��j!�@���� "O0���#�\�×/�t�hH�"O�a��)݆H�ؔ��N�?W�tq�U"OP��a�Z%#�Xd8wOϺf^Ơhq"OriGBA�*���A�G)M���w"O��A��'h#AńԷ:�^��p"O*��6�J�)��ճa�9j��r"O�Z�5Mp��ł[2q��9h�"O����-l*�}�w�#,��9a"O�"b�òv�ra�%�[3LH�g"O�̃���z��IK�cM�%�Ah�"O�p��*M-�\��0/ ��٢"O�uc�XC#ʬ��̔�r�~e��"O��"�4	�F�i卂�7�\��#"Ot�3ӣ�S-F�B͋��rt�"O�Z�mʫ���Ȓl_>^�v�q�"O6�����L�v�R��6{ߚ9��"O����C�q�v��(�$9�1q"OX=yP%��)�$�0#gӦ4����"O4`���Y��0��tHY*Wm�s"O`�PʋQ��h�$]gu^ ¤"OR�/X6-=X%��D�
s	��s�"O� (����Y�0E㡂��w��b"O~���b5&�`㢢�/l,�I�W"O�1A��I��@Q�a � �	�"O��)dBX5fЎ`�U+��&�+Q"O4���o y��B��e�&�"O�e��o^0yIz蚀�W��uR"O�����1"�`ȥ(�#�)��"O���@ʩ^K腰`��;I�a�"O8%` DG�P)��Ȑ�06��"O4ᣄ�� q�u�ӂB�|Br"O�!�&�H$��LB6x98"O���%�F�s�zh�D醗E3\,[�"O,��FG׻J�Lm�0H @{��
�"O����%�0G�Ҡ��ƲWe��"O�hB1ɗ$M#�����EDI�}r�"Op��	�,���0ݚ��"O.����9%��j#Ɉ/":��v"O~ə���F�܍�K޾&D�7"O 8@]8���6k�.oV��"OV�H�oֻq���J�o��"`�-:`"OꤺVH/��[q I�R�&�*!"O��P��`v��C�̓$�-Ђ"O��Z��6��Bפ��{���� "O���i��G����ucB0�L���"O�Ģ�d�1ժ�{��ʂp=���"O��*q�ŊdL ���[0c+8#�"O�-P�MD�D��[r�E�!T��"Or�(#� =}g%��R���{�"O�����9|a��1�HW�$�5A�"OP����(_��)��j=��,z�"O���L�.��� ���׾T�"O�Bq�s���v�ڧ���"O �a��S�?E��`�IƎ}�R�`U"O�\�At~�)B����ܤ`�"OT���[�K�|���.��->����"O �XR��"�� Foͽ?�L�j$"ODe�g�٢;Q�x�S�S����"O�q�g�_��y*7� fϞ��t"O �⊘F���._1��i�""O�{�G��D�vlS(u���"OZ��di ~�+K�'ޒ	��"OƠpw�~A"��Qk� <7�""Ot�x�	���j:;�0l�Q"Ol�HEƆt��ԥ>�<�"O�|�dJ��.�
����'Y
�8{E"O�9�L�k���b%�,0F�k�"Oy+�eJn.8	q��`�i�"Ov0� ��0r=C�$ر�6"O�-��M��Av��R�	k�"Ob�{#��U����3�_�X٦-��"O��I�8OK��D�^//Z�3e"O�
��|޾,����j��$X�"O�H��
N����L��0�0�"O&�0wD�%τ|Y�����x���"O�e�R�;c���uLЕGr��K$"O�XW�T$w�Y"a5n�>�@`"OF�2$睛p��aA ����*�"O��R�Z��k��'?�(��"O�񈴂W���AO�u�d{�"O�Ċ�
�E�9R�@�f_*�
"O��{T=��ɞ(�ƅc�dFam!��m�Z�#�ρ�|��]���D!�Kd�Yk�J^�{����� �!���S��%���U�+4c�"z�!�� ��I"�[3,�i�H՛�����"O�a��%J��pi�'��$殨
�"O�9�E��T��� GV*n�h�"O�u�X�H�ㆄ��*��b��$�y"ᓮr�$ʤ�z��8���	�y�m_	n��!J [�A!϶�yr� A0$ۢ"܆b�Ԁ��bI��yB�_  k�����I6a^��6�ؒ�y�B�8;d�a��((�V�U
�y"
na"��V
��s`��tdT��y���)(��ǂe�X��!�y2)��K����0+ЈRP*99����y�/ڽ��py�Ǜ(Nxj-�2��)�y2,�3��I�/�3Ƭ)�`��y�n��g�<�� n�2*�t4uA�y��D�M�D�A���.Kƈ�+kO4�yd�|x4�rP�=�2�!tɕ;�y��@�fA+"I�=f����-S��yb��Y�f����L #L��ye�"�}r���CA��I�Jb�C�4���JP�Ȁe������hB䉻k�R�H�HHX��`q���h\DB��>r;���ԍ��pp��"�B�	�R��}�CX�[5����)�6w�!���"za���gA��6�n ��
�z!�dƇ8�*ѻT�O!��A�L��P�!�$T�AX2� 
�D��xC,o�!���!_���`O6Wތ��ciRjT!򤔁A�d�R�V�БHюM�6K!�S�*�@d �+%�ĸ���g�!��аR��p��_�4ӸLi�oB�!��
#~�\���FȦ=�t@�",!�$�7]��#m� ҂��  �ch!�� 1�I�[�'�:��Q�%1!�R-T��� � �����4!��]8X�X�`2-��|�>�����#L&!���=D@,)��ݒv�<�A�ǉJ !���#��=BlӶ_}�4��^�!�5�����-�Ii2ap��L>'�!��?b�����k�c]��Af)�;�!�V�������
W�}�	8!�!��̀9_��1�A2}UjX�@Ǆ3�!���+E4v=���ږd,؈�1G-�!�d�>5��8I��ъ5��f �r!��ۼOQ���AE9|L�ʂoZ�RF!򤐂~�>Y	�LC6y*��2!�S��u��1B)���]��!�D��$6�h�[:`����&ݖ+�!�d߷3�N�7n��n��<[�f�.R!�d��b��Q�B4!Lj�z��y�!�]>{���F��s_��j��;w!�D�%8����PoY:J��˥�_ !��"sYV��B�:5ޱ &���O�!��-p�ق�#�� 0�� �V��!� �L{V��T ��|�.X0�$V�jt!��#iT�4	G�A�< C$��FC!��jy8%��"S4-��xJ ѓ3)!��T70ZMc�.M�~�`Z-�!�dZ�+?�Ó�7e�@�5O�>�!� �u]�����Q3x$���S3s!򤚨�2L��#Ћ"Ů�sA�V�e	!�S7q�r���ƀo`����ӥ\�!�dē:����G'�t-!�nO�q�!�@8WT��(��3)�^�8�.��!�� F����X�:�kնT�N4xrO.�B3��ho�,�"�O�7�<��4�XǦu��biS���YY������:j�⠄�Is�'q�51F&Q�s�D�$Z.l֚�)�'���pCV�;#��GlC/:5p���r�"�S�i �<��9@�K��)��ۚ�!���o���bo�d͂g�X�)*ў$�'��OH t��������J�0;xd�"O���f�;?�L�	��\�VLTY�'"O��νX�x���V��0R"O�йd�4=��лER O��|;�5�I[������8s���c�2�ޠ��-D�d� �V�KHF+���-`��8D�\�ц^+.���	��p�:D��`F�˶ �a�ы_���lR0d:D�ll�d	B���7R�[T�7D��҅��{[�[E�S����4D����:�����S	�,j�'D�P�4�Y�'�����U FV��$,#D������g7X�* oՐ@]V<�'H D�D[��C���vlԥ	(�;f�>D� ����X��@cS�D�[ꡊ�J!D����Z�Rh��_�A�Խ�U(>��p<)��aO@�f�D�c���1XO�<�"]�!^&� e��7vu�IdDI~r�'���H���S刐�U��g�������@�T:�e�#݋}�Р�b�S�!��rH����wzĪWk�n�Q�lG��N,_80[����6��j��T0�yb+J<�΅�ƣ�8<��<�7+I��yB���p8���l�Q:�/K�yB��zF�	Q2v��-�T�����p>��չiz ]�2ɸ=�*@¶-؟��#DL*fJ�dՀ#"�	x ,���A~�"5yN%;�ΝE�p�"ul�=��O"�Ɏ��O��(�#��<|d�t�Ԭ*<O�b�'N��`�H�ۻ?�d,���@��y�h�W��JN)6�Ґ�`�Q���y���<�vo �'_��yBc	1������h���?�&'��E��0
T�؝��H!tˍ�<A����;�\ms%jӐ��%&^�)IlC�I��&pI��W�d $�#�o���	g~�`�z8�08w��Jj�,���X�a��H1�O�O��c$eA	�F��1B�'�J4�E"O�Kڞ�6ވ�B�D$_ʨ���Y�����	�*!+����,�<o�T�'g�|�� *|@T�e��$r
��f�W*�y�ŀ-���lG�d����V����'VlBP�ёBl,�� 7N�xdҍ{r��?e��O�O7ZJ�%צ� ������A��ei�'DLM���f��q���<X|�R�'V�I�"�X�.��(h2�'y^�����'�����J���cԀX����'� �i��2J�Y�����U^�P�'��X��&l".�J��
,G:a�'�X]@S����K�
R(Fv��
�'���
G@T9/��1Rwi���B0C
�'���ځa�W�:���M+�5{	�'�(�(m=�.�HBE�*̊��':�����v)h�R�
C:IP�`(�'N��u�	=�X3�D�r�*�r�}��Q���'�L� c�Ւd��A�m�7 {��ȓ"b��t���U����� �(��'eN����y�% ��~�'_��@V�ƽ$K�t���	c1������ L�V�au���<#x���"O�Ē��<h)�N��k�L����'�R�x�� źچ�d���9 ��y� �����AL	��l��W���а?��':h SC
�11���ō�knz���'o�y�C���WIэ^�L�R���HOB�)/§7KL�ۆ���$�� �זbs2���'�u�c��P�,�аnN��~�8�,%?���i`�8��kZ����q# (M�!�$�OT�ض�Z$�:���N�U�`r�"O&�4g6wOƁ`&+U<9�Ҩ�F"O U0��� 9���b7���f�n��"OV\�w�	�j��@
�C� ����"O�xsl�n�m�gN��4���;�"O�@��l��,�t�3�PN�Y��"O�urs�֬U��꤬W gЌ�i"OhaB�Z�_
a��N�H}��"O�-Yw&�,+e��*�5 Fm��"O�NЇ7"x)B�J�	/(b�"O�����r��	�R��䲢"OĈ��
�|㮼����<\M�e"O��f�v�u(���@"b}�W"O�I3`�; ��+��٭a*u�s"O���S��O/�|˵� �p�=��"OD@�@f��)�t	��KS�^^(zR"O̥�W��t��h�Jd�"O@�IP�N�i�|)q�h4o7��B
�'Zx���
0?�2�HA�<�Fe�
�'Jڰ��+�S��q�U�\o����'{2l{�[��(;��V����	�'ㄴ{�.��Ѣ���&PJ���	�'S�ّ�
�~Q�if�\!F�yS�'0���^�#����� ��CH�0޴�Pxb!�J��&ƃ�%>�0��,�y�-S&� ˠFM1CuН�����y�ٌa��h��h�4dBh�fɛ�y2��7����DHƺY[�Q��kצ�y�'^1H��m�P�?�2�pp!���y��<���S�;8*�I �e�<�y2�҂{?x���A�,}��,��Oǌ�y�I�<#n���\
xVjuP� �y¦�-"y�ɫ4�Ӻk�V��6����y2��[�����^/��+FA��y��LWr�jF��"��(�ɋ,�yC�L��� �ɾG���j����yR*M�`u)��H&@96(�$-���y����{���3 �<4�0�dי�y2�L�~"I�`[�T�2h�#�Ծ�y�U7������M��{椉/�y�.:Y|t�6��L��i�ك�y�M�i��д
Y5L�4ى����y]%J��}��\Q�P���M/�yI�J!�؈٢K���� �A	�y2���"�@q�#eܘ<-B��냳�y�K�"��a��]�}�b��pJ�>�y�¸T��"q���(�
8� �Ŋ�ybG�:%̪h�2�;(������yký|5,����uSQcU �ybl��Mx� �����"�h�	�yR����Iꕈ��fΤQee�4�y�)V2��0�w��.z�|AEn̯�yG� m��]j$��2#�ĸC��K(�yK>ttPB5�YJ�̢6��y��U�y�(���J�d��!��_/�y
� bh�F
���H��
ɽ�d푢"O�Hp�(y�&y�!)�k�Rh{�"O�5�#-�<3�\�#�U��"Ov��S�Dɞ<�v��OS�L��"O� 
s�߼wӬq�S��<Q�	
�"O�l3`�u��e���C7~a�w"OZt��BW7V'�\3�gհJ�4�7"O��
��Vo>A���U2��}	"O��6�H~�\���팒l���"O�x��NNx�rK8y2J,2g"O|��S����d�VK�#����"O���.��z��L������A7"ODY�u�KpSv�S�ʚE(~�["O��C��(k��D��o�(����"O��B�
2S�H��U�˨"j�"O~�zU=V~��%Ծz�t)7"OB�Ke�ih�ZWE���2�C�"O��p B�:p}�k���a�6,�"OT����JXH�M��.�JB`"Oj1�T'������	֝X�v��""OJX�/8��`"�Z�ҥ!4"O�T3d-ȣ4�>��N�����"O�%K��=
R9�"$��IǄ��0"O�PH�/�NsI�b��Sb�Ԫ�"O!��͕p���j�M�Ĭ�G"OZ��N�?��s򉗔��L��"O�,��Q�X� i:��V<�$%#A"Ozu{qφ!_Q ���a�	�-�"Oڌ:�M�a�ʠK7�H		؈Ҳ"O�-�$�%@�h��GnŊ;�����"O�x��b@�>�� ��7�d�YR"O���擙*f��k�H����C"O��0i&-H�ز��mE& "O�<S6� �.�#3�M1j&H�Ie"O��9T�Q(fH��MƼ|����"O�C!��0Y���+QNQ�x�B�"Oy#��K4@@!���	�FB�b�"OB�(��3l��y�0l˪+,��K7"Ou���mrh��<AV��f"O���IÈ?��,a�+AY���1f"Od���ND�9Tr�3eU0W���i�"O(I���@x�p���)6r��[ "O��
"%�=9W�ɀP���
^68{�"O.�����C��� ��.0��(�"O�`���1�~jVo�/�:	S"Of��B�Qh��a��F��"O����JKl��}�%d*G� 8�"O��S�W�~E���G͓N�&a��"O��AB\�ʆ��6E4:�:�D"OR��r���ܸ��d�C��4�"ODl�DۍsH���R�L�R"O4���J�7��Ń��H�Y���"O��B -y�)�p��0O��T"O8MЦ�ŝsw�lx���q���i�"O���c�,�mS����~�:!�r"O�(ò
�1bWhQ����;p�"-��"O���4�_� �ne�0�T�:�1Q"O�ٰVk
f��L��hMp�p�"Of��DR<9����L2B����"O�uqdE@#?�lD��(�E�؈`'"O|!��E� ��3"k�"�"O���=/� 81�`]5y5�葠"O����,
��8����(*7��"O<�d�T�س�U�Px��k�<� ��Aw�5E�|}�-�35�T�#"O���J�'�UCl�2� �QF"OZ��Ŏ�ypP)F�}�(ȑ"Oʬz��
�K5L���I8�0�a�"O���i�D�;��'gp�:"O����O��lV����-[�T�V"O$t�2�ŗz!*d
5$O$4O��"O2�We��Ȁ���Ö�*0T���"OtT���d����bH�@4p刕"O��!��P?x�<E	�a�"0B��Ѵ"O��1��T�gB�R��y%�U[�"O����d|!*�,��j"O�!hCC�	���cg/�)>|H�"O�Y��*�q��I�%�6���"OB�.F>?N�ݣ�lK'h/�,�"O"���B�c\�Ԋ���+-����"O 	�%�Ҽ�^�t��/���P"O�2���w�r��	�"p�0��"Ovq�������+ ��% �$��"O찔)�
B5�5��]�|���"O�#�CQ�l�8���T/���E"Ox �T�H��qUg�^�ju�"O���E�Gq����f��B���k�"O�ؐj��hI��HѦ�%f�Йc"O�y���)16�@c�)<%B@�"OZ����� +S<�kV�,;���Kb�<qu��0>=
�G^7"myrώ�<���� ��`��
9R	����!�)?�b�dD{J|��C�	m>RE:�eΐ}�B���Ws�<t��-`���z!-�;�j<��h]y�<���r�����	(q`��GDJr�<�� �)��X�T�N~����p�<��Q�?w�ăkϚ(��"�l�<���+b��>Rzt��푴�!�M�iǨp�AE(L�a���!�A�#Ϝ9�`g��81H�/Z�!��V�	�pi@Q!�9F�-����!�!򤅈.�Ty�V!/hK�-��
�v�!�dC+q��!J%mO('-�����!�!�A3i�m	�H!��8r�[N;!�K������J��-�4����$v�!�؃<�-����:F�,8�@B83v!��9��u`�/M�^Ɯ��rfG.5`!�$�1hO�R�!�Q].I��^M!�F�O�2\z��՗ U>�У0O0!�DU�>��I�wL߲w'm0Ӣ8Y!�dC�V��Ajw���
�L8�Ԥ[!򤅛%N�F��5��E+����hX!�DK�Y�\ʤ�	>�Nɻ�/܄rN!�dB�R��6��j���#'�	V�!�DE�>j��2w��3�0(1e��*]�!�D�"a ]!�"7��bTM��p�!��PsL�-��>�{�E�To!��>MB�+�눪u��0�	�~W!�V�̄Ib/W�(žX���,hI!�DT0?�	ScW�ڙ)�ė`<!�$Q?W���˶o"x��0��B�k!�,t���І��Y`��i��U,$!�D6	UX�#EݼF�.�� ]!�"\����,߰:�N,��/D�L!��ڻe�r� `�~��%!L9*!��3T�I�s�Q1d��dC�bޫ2!�޴e2h��/�M(zl
�D
.!�$��]هH�f����G�"#!�� ���-�#fO�����% .�M�S"O� ��O*R��qk��Ø���:�"O�Ijó10���W��x��"Ox� �%��6Vؼ�A�m8A�D"O��Tc�5j���&��0����"OҤ�o;0��r�W-�*,JT"O��k��Ha�ȡ���$t��4t"Op��O��l����ŢƼ;��"OL1����7��m`��$����3"O�l����p��u��.;$hE�"On��S�ɒ+..��A���CUd�2��'P�T0S��L�,H)ؔd��HH%3D� P�[&���7Ȃ�sZ�`j#D� �b�R(��B[�F�4p�Q�?D���v ��� 	�Fٸ�Y��;D��1b �eF��BM�$�bU�$@=D��3��
�#6�P�,��b# D����k��9�ܨk�F��v��h�:D�\R
H�6C�p'�X�j
�X��,D�4�F%�(����әA���-5D�<��
�,��!���a�Ԙ@��4D�L�1��,�<9R�O�+lޥ���<D����L�E�����q�͔)�!�dA�5W^5�'l�%�l�&��q�!�d�N6�8�v�ʔ�!3-$'�!��Ka`�����=֤�Zˎ�[!�D��m���P��<S���!d��_!���$8���C/���E]!�$^��hȢaJ$��R�\�X!�D��y�����M�x��h3@���M�!�Ƕ%r�� ���tu�ECr,h�!�dτo8Hؖ �
lo�D�������yBቼQ���@��)G�d��d:�B�f3��A�m�� (�(���B�g�@ �d�' Т6�6G?�C䉈e �1�R̍?��1�H�9�RB�	��.�
��R�q�� 0���i�DB�Ɍ1az5FB?�z��a>�~B䉈f*��q�@
^vb�)�L�RB�	��B�FCőX$p��LN#�"B�	�L�h:��x��qT� l�B�	�n����F0u��-����+(�PB� 4 2Ȓ��ԧ��ő��V�b�HB�ɮL5T`'�*a5|����wlB�əq����KT	 t����>��C��=���P1���M�BiPF�%X��C�	)p�t�9% ,i�A��M	�g�`C�I�m%�X�ՆW�2��2��D��B�ɟOm�A�ON�Q ,}��.��<nC��%AwN�: +�
�ԡ0fҝ��C�Elq5ĉS����EAP(P��C�I9_~��1�JQ�qܴ=�bL��p �C�I.�&��P.��f�<�ZAU�'ޤC�I�o�������"G^ɑT�1`CjC�I16� ���\��x5�O9�*C�ɴ�~�`@��>hm��+-��B��!L2�ԃw�{6���uZ#"M�B�I�;����
�_�K=A���"Op���E\,�:e[�&׏w~��1"OD��O�>xGX�j�$��(��r�"O�HCG�1~��9s��@�Pa�@"O��a�J�DfA��8|�,-x�"OlQ���#IF�'��~��$��"O*���*C�0&���$J�r��kF"O� H�S$˜�m-с�Y&"Xq�'"On���FM� �P ���5+Dp�t"O���׮D�d8�⵼B�b#��yҮE�A݄�ش�Vb;��A�@7�y��N�`�eJ��6a�Dc aQ��y��;~�&���'V������+�y��N�h0�'G�VXh��Bĩ�y�(W<`�L�y2Ŗ��Ј����)�y�DS�L��%���J=bМ[�`½�y"�[!4j�ǎ%l�EAԂ��yr P�N\��C��U֨��"���y2�YG�Y@�FYZ�Vec7��y�.�j�2`V ��Q������y�5sƆx�R(G���X�䀊�y��.b�� ��� �V��y��iŮ��q���z�L}ʃ$K��yc�����m"��X�§Ω�y��&�Ti�Sbh�h����(�y2�܂p��1B�EI�Z-����8�y̂�Y�ĵ��"ߐ`ڎ7!^�a�!�Ğ�Jg���GԄ�v퉂��'�!�$2RppXC@��<E�0�E -i�!���B*4��&���s3@ Z5[�&�!�Y�*e
�5΄��h|a/�5_�!�r�AR��=v@ep'�;�!�䌄0�n���A�Wb�HHfkO��!�䜸�U2� ]���YΨF�\���?j>x�TmO !�z���e�D\ ��ȓrpj(k����bъ��G�����i}�(�JQ�+�J�
Q"ߜ����q�`\z���$�P]�sY��j��&@��,0�����=ar��"!k�MR������a�"]i�<�hKW��kc�"4�tcš�|�<�%oƂ�j�@ C���	�@Ic�<T�\Oٓ�j$HS��i�c�f�<	����,Ȇ�]�W�ZEQ�u�<���'¢m��H�!L)������D�<��*d�x�7��4=W �ŧ�Z�<)�J���`��D��~���h�U�<1'K�?eza1�R'E���a�^�<�F`��#�޼�Ϻl���a��g�<)���d\���ڷp���K���]�<�Gŉ�m��a� B.l����f�}�<�R&�vm2A{Bd�=l�"��u�\�<1��	S�@�q-^5,�8t[�Y�<qB��x"�������%��Lr�a�}�<��Tw��1�IIm�Z"���u�<�3+��b�>�yQ�{��)�@E�h�<��䗵Mk���材5 r1ڠ��N�<�j�l��( ���e�y"Hg�<9d�KmpAp���.�zIQ�%Va�<	�m�S����0	�$x�vLp�<1��H�Wj�l�bo�,`��|Q6lD�<�e7E��4��e�+DJ�Eb��C�<A�!��c�D���f�#R��H�-W}�<���T��jX��ћ����z�<7�@�0�Re�#���sF�h�<�d�*KŔ����D��V$3 �Li�<�ᖙ@�`�Q���*����d�<ѱ ��|�p�����%?���23A�h�<���4B�"H��@����)g�Gj�<�� C�v�	ٕiU�u dm�E�I�<�t[/g�$�f��!-֢D0�!�E�<tFʹK���r���s���i'�YA�<� � 1�£} ��(jp�%�"O��P�E�%F�@�Dg�9G�q;�"O���U�E+58x��f`o�)D"O�<�D��5��P0R��K�fD��"O<��p�88����i$S��\#p"O{G��S6
�j&H�$|�a
�"OXȚ�aȡn��#�G�k:���"O�a��ʺ?�V�4DN%TX���"OXUa��ڲz>���^!sCj�r�"Op���M#*��x�o��>�iq"O�P8b�T�iBD��ͅ�#r*!�C"O�+#ޙ^0��A�/�&�ր�f"O4�"�F�1/���K��S�U|$�#B"OQ��

� l��D�Ae|�+"Or����O'�8X�b�)cB��"!
Ob6�^�%��Iw!�$p�x�r���H�!��LpD�r%���}��t�7٤��xR�I=+�$AaV��}����z|�C䉦"�Q� ΂���+0kt5��'ў�?�� ��~�ִz�B�2Ԝ���3D��Za�I49�p����_���Y�0�o؞(D��	.�Ѐ0�.ɔh�C�"�nڀD�fT9tgT<:�(2%�	,C�B��+��� �B�8����$�Fb�C��,G��@��/�l���*;�ZB�	�Xo�ݒ��$6�Bxkq�խ:&lB�IP�����߬j�t����- B䉙�Ԭ�#�.$��Q�u�VB�0��3�B� ��dD��0�B�	�v�!��9̴�B�� hȂC�	+_0�E����2�ث#)�>0B�	�>��E��f>�x� �iC4B�	^c�5zІV�V��e��cG�C䉰p��4�IǕ���8�M����C䉢Ym
������a�2|j'�A�,	C�I�.�8\��⎞�l��B�	���i�N��	�m�N o��B�	� ��0`�
6^�P���H��C�7�<�c2l؟b:NExd_:*/�C�	2c�Ī���%�V�j��_b C�ɕ��[6A�>���!
O0t�B��!6���#!E(?1���`��K�B�	" L%���~Oh�O z �C�	�`IjC�>o�N�k�m�N�hB�ɰ��-Z&B�=lLB��0M\B�	�Aކ<aa!ܲ"##�Դ0B�	�4�b= e�Ù4�L��n�H�6B�	1r"��ⳡ֫JDIw�LB@JB�ɰ2�)�2GQ8l5T���iģ!�VB�	�YJ̩�	I��z)�w��B�əQLt:���\��]yB��.T4zC�)S�j�C���N�tQjcʞ�ZdC�	i`�y��J�Pt��ѡ3')XC��%H�dL�Pm��^41��m� ��C��,.-�ƚ�7�)��l�H��C�	3.+��a��bV�!1�W�7�C�I�>X��&	P�r�n�[5�ҧD�>�ENa�Q>�7�S�nTx�hQ�1r6�.6D�ĘԢS;����r��V�>"��O8}���ޟ.5�%�"~����;S�z��Vo8��H%�
;�yR`�t�";0� :5� �`�����X ؽG�ƳM,ay��^��(�Ε|�����P��p>�g`�@+1���D0�@��
�/i��ɢ@/��� ��*$�8ن	��
F&Ur�"l��9� S��7�B@��T�TDګ�?qC���� $����+�Љ T���-��O�j7 
[��hҡ+/���G��t����p�:�a�̟�RG�P����y��/ �(��V�$A+�aa�^���<�&MW&D,�O:��eF@�u)^U�q&�7q�4����c�� (���)/3ب���W�Y�8t�'_�O I�A�QX<�s����2e��|�dE��<u�=Q�BA�$���ɋ<�*���J�+!K��J+dđ��X�,nʓ��=��dDe��1C���1R ��fN�=OqOxlC�g@�#.4�u� w��� �66{�iZwwRTy������\S&+I�	H"D��'�P��D�p��Q�m�#X� LI���K�4�燛���n@�$�Z��4�Q�g?�S�E\��� 4��`ψ�`�WB������p�I�S����08hbp�D�(�+K-f�)�S �:(� T@���^�8�^�P�ў�=r�EW)Lm��	�-�� ��a���ř1X���PnJ�q��9p'JГkV�	�U����	s@���`H�I����Ҩ�Oi#<	ǉ",��x�� ���S���į��n��i���}��E�f��9�yΐ�n�t�[���qU,�L|�
]��n�3 �I��0rv����s�y�!ùv����ª��d���G�=D�t*#j^%,���W�MP�Q�0@��1���@��H�y���ر��	��O�'q�.E�P-���M�BP�P�G�q8�H1��	���e�0mD�$ƒ*
Y!r�͌Q�,8qf��L1d��$S�L�\�w���]��{f/Ӏ,*Q����&D�p��aǨ[��SVo�|BB �,aRP���O&���nF�<)�a�V����;�Q����Ħ�Z���e���gA�2/|���p�s����%��3X���]�(M�� "On(p�I̵B�@�a��Nɳ���5��\s�7�a�I��^��3�I���'9�@��$@ʸp�Xp����q�Tl��ϝ�$��Pw"�~�搰���;1��E2ڍv!:���z����ŧV��a@��۳B���F|b��r����C�"ZhcFX>U�	��f���I����r54�,2D�Ԣ�@��4_�-�ui
�hE ə��q��X�E_�����$�
��F�(�*Q��`"�*J�"l�q���2�yRo��r�@hVc�P`iT)U+W�ZPg�
���])�0�
E�?#<y�X�lBҹ��1Q�u���j���ʃ��3�"e�	��sƉ����xP�J�%)���"P�8�>�+�?�T�
��O�a�l����g�'�x��7�V�YO����"�R�:��k�Y�0��,0�h��(��Щ�) ����K�'@bl�C����(-�R�2r��)��?��葬`�tL�$k�*+�Q`�->D��c����!fJ4�&��O#���d�=u:� ϓAl���b�-J����''�ec��C��E���z��s@�'��A/Z1"��H�GC�C����F�Q����h�J�z1��9�UHf[��۬S�Ь�G����D~��;e�h����?@մ�$�D��%�6�j��7��~[���_��d��8"p��M."f���'V���A!K�l_z)��=��!{���,�}�cF3<� Y�q"O��*��5�vT���>5�ݢ��K,��$�|i�=�+7��� �lTS��1�11����9��𤁀c�,�Z�%��f��e�Qbƴ6�p���D[�§3����!	���원�0=���T%�\�H�^�b�
�9c�@G%!򄀉x���Rs	���eHr��;z!�dS`b��"ʔ}҂,#�*�Xg!�	��$p)�,K�J��!h�+~!�d���	��,)V$m�焓0G!�$�:*I���U�%\�;ǀ1�!�$�%A^q�N���Q��'�!�D�uhJ��p��U���Zdf��L�!���75l���`�-�8*E�8�!��Ά%�Ȅ8'��	ӱJ�~!��lL0������E)��	���>��M�Z�r�Lȶe����A�c��x�'���:'φ�p��PF�	���1��'��@�7���Pg�����=r�E����-�򒨨�k0m���C-̢.�x��S�? �8��pN<01�'n����"Oh�Bv��|�������-�n��"O2(��P�	� |hT�U� �A�"Od-n��eR�8�щ��H��"On!��쓽֢\��!No��h��"O*Hj�ߺZWZH;���?r���Q"Ob(�2jҳd���V#6C:�;g"O8���"���#��A�h�����xR"�T��zr͌v"�`�HP,� \������y�-џb���c"ǀ�9���!H�y2�yg�)2� U<k*�� ��y�/�8F�|��d�j�0� Я��y� 5�� ���T�kh\����>�yBEƦ:�Ā����Z�qp�ŝ�y̆J�f���N��b�U
c�%�yrFI�#����N
-S\�ÕW�ybR� )��P2� p�X����y2�$&R$��2˖�Ib)�����y��
�]��e�ra�Ը(�9	�'*����Zk��K2D�!$�B	�'I�@X�'��yp"X!�n0S
�'Ӗk"�J����Kq��	�dL��'�i@��oݦ��g�3(C	�'N�Y�EB�� 	D Y�O�	5��h
�'�I���0k�,�bd�<Z�[	�'�LrA��ꙡ1�ݨX�#�'|Ԡ��7E��sf��1%�����'�Fݸ��N N��Х( 3 $ ��'���'��!$d(�fS�1N��P�'q����h�+4�L7~m�Q�'"���g�Ls�(0��v^0��'Ih�`c�F`�h�A)eZ|�	�'I~�I�(	�7���z��ehaY	�'�А�! 3u y��IHg����'��PÎ��*aWKǊ&�ʭ��'�XP�'Zv�PE˧/Ʌ��� �'�$)uk���jD�JW3u��Z�'X$aƯJ�R��y«t���'����!�[��	� Me�P��'p�LȕiV����.��Z�0b	�'�����Y�� hă�7RW�eA�'��FNK�k�ƴKd��Pp�q�'�����Y~-s+�&��s�'��*����D̮m	�`
޲�;�'�\�WM�B��LcA��p��
�'=��2�.�t���Q�&�n���'QjH�4,R%r
:mq�#�HX��'&�	��*Z�4m�G�Ƃ%^�)x�'1b�۰BB�=�`����K��	�'�VI�0h�&A�qA�!	e�]��'�ƙ��C��S��͸�m��	��'ԸW�G0�:���)�\<��'���r�	�:8��)6k�3L���'�����+,����?7<I��'�����2U(d��P�$ZM0���'_�yQ2�� y=ؑK`c�^��`��'���V���?�F���
+N�\���'K<���]a'�h��kBh;ԝr�',����&��q&U��a��h��']̕��+�r�,m�⊍�6̞}*
�'�rīc�M�t��Qv�j=X
�'*ؚ"��K�����X(?Z���	�'�T)c_+Q��� ��4���'�4��7cZ>;&�� O_5��q���� &x�5m�;@:�E�Ԫ��(o.!�"O����A�+[��dS��PJA��Y%"O�a1�ǟP��P�tf �LHl��e"Olhs�V�8��q���ه@�����"Ol�I� �
Vixi�d�"�b	�1"O�ڔ�Ū2<��2�dąs����4"Op���$;<5�!}�|R�"O4趣��tZT H�/�+��͘s"O4|��Y��i���}��]J�"O���@D_�2�|ٰr��5z�"��'"O>a"��	�3.I�K��j�i0�"OΉ#����T"���(S�ĝ�"OX@�����¸2�����
�y���V�衰/�p#*��3�yb�1�ك�՜p�d�׭G��yB
Ӻ6���S� [@%:7O�,�y�g�~�LUɠNM�.��v���y�Ō�w�(j�gG!1�1�mV��y��ܓ�� � ܯ@]���fӀ�yB@B*l�H��@�D����֮�yrk��@N�X'b�*1^�T��CD��y2�� {L���Û75@�X�`֞�y�ș�F�e��.�7<�PFiϖ�yR/ɖH�L�H���,$��R����y�%��-�Xh&KJ3	�l�U���y��D���c@�H�p�4(X�yҏH.kp�+���8���c��yb�q��1	��rܶ���G$�yb�A�P�>p�b�҇rM��q0d��y���#X"��c-'o����d_)�yb�ט8^����� ]�0k��ʤ�yG'0Ġ�$�N6H9�����y��#΄�c,R�:�ƁB	L�yÈ�(㆕� 8 W<Б�1�y%�r�A�!��jQ���'�y"ȕ%cb�:'�Z�(��P��Q��y"B�2jy(�j�e�=aR�oF�y"�y�-: �+�t��'��y��~Kh��խ�7�Z|�"�Ѕ�y�)��BLz��ֈ�=Z@ѧ���yb��1���bmA�iz����в�yB�Oj^��g�?*�L��#T-�y��o�N�!�Y�'Ǥ�3P���y�JZ�V��D/� J�z9��9�yB_���ӧf��7��(�)��y���y{$|Qw�Ĝ/����
��y"��d�i�ʫ�:���#�y�`��N��,����z�CT��y�π m����,D�b���Ɛ�y���Z���e$��6T�S�P�y\�u�~L��_�s�20���2�y�
��0v�����tw��
'�9�yB Ѳ:P�G�?:�^ă���y�)Jz0pa�T�m�J��5	��yb��%E�(� F �-]_�h���Ó�y��-/�@�yS�RLaD�
�%���yb��-B�����%���4)�<�y�hH�0���Hq�X'���	4��B�	��B4pB���+*�DQ`�ܜg�B�#,�z�Y�IM� K| y�H�~�B�I�3	�S�^t
�It�W)]�`B�1k<�� �K578���C6ϞB䉼l�~��R�X?kx�2� 
-
�dB䉰r���h�V�^�܌e�F�l�BB�)� �<�F�Kc�*1r%*�'n54���"O�Ļ�D��U�bnڝ-l�#"O�hp���v�0Q����(P
�a�"O,�i��
���r�m�+6{���"O0`1���%�F���/�)}d�� "O*��&�'c.�kD�2 (�h�"O��6��L0��P�Ə�u��2�"O�=�p��'LÊ  ��Ć�� ��"O�uI��E�;� �c�K�3QΨ�"OnyC�jW�A�|(j��'s+Y �"O�eB� �I�.X�)�&]"Ov9���J�������C���"OPHȥ���;ن�D��B�& f"OJH�1�{j�Yu%s�y�"O�l��'Ž�����gDi��=`�"O"�����W�� QC%_��jrB1D��(��<g����N�>�a--D��b��ߵ5�!:��;r��f�-D�D�v��/<��Ae�Z�mٸ1V(D���P���uR�V$cb4���E)D�t���AJ!@�P��w�X�(D�P�a��_��aP/�%���B)D�d؆ݨ�ʬBF��2�=�1o'D��˘�:"�!�X� X�Ų�"D��C`���&�̐s��؎f|V��T�#D�<�� �,=��=�,.2&��`->D��#�i�	���*8�4�g�;D�H1�+�B�� ��-�>�\�r�-D�(!��Υ-��A�ы� S�����j-D�T�)@��@ ��G��3�t�R�>D���%��2yV�5�t���$�Ń<D��C��HD� �) ,J��g=D���$ͺ��Xi��$m�xUEk:D�@b�&ʅ&���h�ɞ�$y"u�8D�t�e��s�|��3�]�7hp=�"e+D�rb�D�
c��[�#W�a
4$#�%(D�TP�HA>��ʦ�/�>h�Ō:D��s�-վ%�y�g-�^�J�'D���̓��q@�7��(��&D�l���Բ Fj�p��BҎ|b �0D�p@�lG
BH����?Z㐸I�=D�,��o	�~�0��d�8rN�2�I'D�x�3�C͂+!o�PL��¶�'D����&W-�V�e��M�����
(D�l��퐐tD���<p��1J�)D�|�oK=O(��䞦,3��3â'D���w�ѹ
��8��FH�A5�%D�T��g_�\��	v����|<If� D�Lp�Ϳ(�D��'�mr$da�%D�ă���)y�0�����10ʷ�$D��c���=,>-k�Ö�O��}���,D�$�f!>��ذ�%ih�`d*O���Jqˈ����&�V)�"O��:U�U;38�;��A�~L�w"O&��R�ŭ?a`9�cgT|��p��"O�:VI�B>�%�5%�4.��P�"O �4�N8N�|�a6Ɖ�z>0�	�"O4����$d���(���kP��'�yR!��l:4��Ș�Y�u��!�y2l�^�"����`#���b�%�yR�ͮY�Yr��Ǧudz�;�*���y�숯6M@��r �h/��ӧ�&�y�枈e�
��U�?�\Հ��y2�ʥt����q(V1%20P�T��?�y
� ��sq	=l��@R�Q�"��#"O ��b�ybJ(�%G�L6"O쑰Մ��K=��e�VMt��"O�92�
Tↅ3�H��Nڅ��"O��g�S: ��s�gV�pF�QZ4"ODx)t�78�r$�G�FJ$��"O@	�G�7
x����/�����"O�%��KJp������a��4�"O�Qa`#E1A�������0���T"O�e��EԳ\P�u
��X��lAu"O(�K�H�,f��$s�iD�
9��"O����&�@���$H�gS�,��"O�� d�,n�60��b�$:G~l[�"O�<�����΅+р�wؾm�4"O�h WC� � �`S�.�p$bq"Od҇! `�t��V��I�T,I"O�����L�xa�P�E�N=<�v��u"O��m)h�4������"O�a�bϚ4`V(��F������"O�u���6G,���͘/��3�"Olp1��-�0�D���	�ZQ�"OD���ȏ\�p��*k�2�iQ"O�$ 3���
�:B��y���D"O
i9@�@�ez�!S��_���"O॒�g�Z"D�ԩ�6x��(�2"O�(S�`R:hz5H�L�m1�"O�4!À�+7��``ؚRQ�ы�"O�J���;��4�fY	gZ=��"O�|�Ə]\�a�gܒOzQ��"ONmK���b��&EI�,N��rB"O�1�+�X��{ �Q�jʚiB�"Oΰ�'�;ZN��JG
��A.�1�"O&}���[�raOV�\��<��"O�,�C� �'*�5j�TV8t�(v*O���Ċ^�@Af��և�M�J�	�'�]�Td�@�P�Zu%�C.�l3�'Ş�`A�5��ڰE+��'嶝��J�ĕ[T��4g�	��'s\x��J
�2Q\��F��+dX<��'D��S�%Ԩi�{B@O�<z���MUA�E�ŉ�.��O���׃�q9�0X$�Z�
�S�'k��S%Vrt��T/�O��c��ټ5��Uj5g*L���t�O�?=�e���i(�,��BhA�Ô싣_G�����~)�e�d^a��$l�T���&q��R���^�E��i/`�牫e�l5�I|Ҍ���_���5�,jW\,���	Y�I����M�U��e�~��Y��ɑ�A�ÀV� �,��$�/-�}D�i2�� ���ynT�[���25���#�2!�7��
sJ�"�7H��l���,[����J�$y�����';�Ⅎ���,�����AS� `�,�>ل@����'B�rih�@��4���,���%��a`�s�S�'q�¤Y�R+H�f���?$�N��'�XE"'�?�)�'=C�3�(,zv����hE�i��3�N�#�@��=��ɐ��;cd����#/��p�K�/+̈́p9V�H�i:��Z j��W��lHW�O��S�-,�	"GQ�nn�IX��uCJK�l��Y��{�@ƌg���i]')���@����Ҍؚ}�q�2��<ѱ(� ̊���Oz�)!Ĵ?/�YJ�O]ܰ]��ǐ؟H��B�%D����?�D�tb
��g.F$���I͍0���b��>x��@�O�� �O�b�+U�� >#d@��LB�@D� ��F<R�*�e�*�%�o>Q��9R���ٵw��(bƏU����'-ͬ�CddQ�~����0�����:"�6D�%IÔ&u�\Γ{�:�+��'�6HaBW��}����l����l��xjI -ʷ)
��f?Od�C(O����?���*��A8z�ӥ"�lߎ̊�Gjh<�V�ڪ1��$�V�5���P��k�<�U��Tw�h#�A	�έ0v��h�<�R�y��43A)�?�H@3"_M�<� �Bp�=a:.y8��T�%��`1"O��ɀ��6) ��A�q<P�"O\)�Ü�+���W��Y���"OD��vmΫF�Y�bO��@Ȥ"O�`v%��I��x3 Ɍ�h�r�"O��P*��XSnTQ���,�� �e"O�	�a�L����Wm�n��!X�"O`��1��x�h����q� uq�"O�tk3h�q���8J��/��I[t"O��������3�O��u�XV"OB�(�B׾Q���p�"O���A.Ȕ����&7�~�p�"O)b��؄=�܀2���3��x	&"O��S�i̚N�Z�ѠW�����"O޼#��4��P�"��*��-��"OL� -�eHԪ�ù~oP��A"OR@���U7+(\bǫ�v4�e �"O��	�XCpc��߬&(�|3�"OA�4��TA�a�U�:��W"O��mN�b��Ɉ��!2�Mzu"Ot���+�v�]��'���p��"O���%'�6,��#�eS;@�&%cV"OX�4�Z$����dF�l)
��Q"ONt�UW�B�: ��M�2W!8�1""O��� ^��H1f��sd-Y%"O�l�6k'@��ȇLێY���V"OD�����x��IR�`5c�"Od�#`��'L(&ă�NV!?K����"Oع��% @�pT��g��S�"O���󨋤��*ĭޣ		���"O<�*�M� AT��h����F"O|)�e�� P~`����W�<<�w"O��I%F�/�Q��`�	6�Fy	�"O��bao-ZJ��$�۴y�Z ��"OX�y�������Ʈ�W�*IYf"O`-K��46�|�Í�B�.�˂"OL�i-O+i
-ƫ����a"Oh���+�9,2,�*ܾhF���"O*!�A*lh���0"PY�"O���	W!{���O�/Xf@(�"O�Y�t�Z:	�R�0�..JM�S"O�$ E�֎c������OGĕ��"O:�J�e��?`��P .�&.��p�"OAa4+A���AC�^(ʱ�%"O��Ɖ��W�d)�$��}
��K�"O���+�9tt�sQ�i�
���"OZ�[q嗗m�(@P���;�6��"OE󁋈s����#^���Y��"OfT�k
�f�`��K�: �R�:"O� �p�J�N��\�+�q��Yz�"O�����࢙ST�C�nZ�D��"O�	X�I���<�(%�H4+R�4Kw"Odu�wE�.UL �"Ժ!�"O� ����I����������!"O�r`⟕9w�E���
!�ǘ)�l�T!�<I�h���g޴B�!�$��"Z�ps��c���u�@�PA!��.Q�i�.�j��)�֤Øu\!���?����I)��ī&&�>!��E�
T�(H�xY$��l!�Z-q�}�D�
�:�LhAO*N!�DƝ ���c+ΧF/l�`��9�!� 3�Ta��a��N��H�!��{�!���*��5I�8NL���0��8!�� "�[Gݨ?�T@�E�?x,j�	�"O�ʒ��w�0A��)1�24�"OpQ��Q�OD ݂�EB�:HPD"O�e�FW�&� 0P�.�VM"�"O�m�b��lY�J@�c4�e"O�q:#�G�Jm� ���F=iZ}h�"O���r��n| yp�) ����"O�Q���Q0X�T ��IТ8��T�4"O���'� ��j)z'�1,��0Y�"O
I�bkz���F ��@A"O�ݙrIŲ5�T�P"���O�ta�"O��k�I@��B�e�߂�J�"OTd0��D;y�Hؕʆ�d����"O�<��BZ4c�ޡ�A@W�^�r���"Oи�gA:MA|��7ϖ'5���h�"O:s��<d\t�͙�mx@�`"OV��[���=�LǍ70�IȢ"O6)S�gX26�>�ѨƁx�%Q�"OW� $K��Q��F��qG�F"O.hY�O�3i��sfT5A@,��"OL�qP��:A���$e��h.�ە"O���f/V�M!X\"�j��i��و�"OX}+3.��P��, Gʊ�\Rq�"OJ��'$ϽS2x� ��1���"O�	�OIB	˵�^�p�0`��"ON�I��^�5������V
؎�Z4"Od�*�)N�0��3�2��p$"OH�'g�"O�0�5kكs׸�8�"O����k��%?ĭp�C�F�p�8�"O�@sE�O�m2�*�!�8x���"Oƀ�p)�T7��C&�/eh��"O I�T��e��z1�
`a^e"O�9�QO��*�9���5N�Q[�"O�@H#�7��A�D�Jb�z�"Op�+��?6x! L�4��"O��*Fd�/�fɩ1`�:!�5�6"Op�����4J��a�z�|3�"O�A�@*U��n�2S�ļ��d)�"Ov	�O�I ޅ�%�G�@،��"O,����,n�e���ʄ:(�؉�'qO�	(ԠR�� X�f̂$/x��g"O��#w"',�\բQ���,�P����PG{��)N�)`�GI\�_�td9��&6{!��U/��Ųl[	hx�U;F��9*�!���V`bI����wu.yҤ�^(t���dw�t8����4~L�5� CHR!0p"O���N�q`���&$պn5v1�"O(`j�F��
}z�L�9 D�"O�ih4�"�h��Q��td�2"O��xF�
,��/W=n�iI�"O"����BXdP��`aH$�:�qD"O>�1�+��[�����P R����"O�4�f�CC�*���M/��k�"O��;w&քi�:��q��5z����"O`�2jD52�%�\I�( Zq/�X�<ie�I�>�MAŬd�h��@EL_̓�hO1��p��J](v����"*1�U v"Oj���LA5'_� c�_�#����"Oȡb" Xu
x8@1�) ���g"O���h^�n&�(��˥lf�"Ov�0��)bREz��ێ�^�Q�"Or컡�:,���aâ
����y"/���ʟ�kH4P�4��*��B�ɀD���[AꜽNp��#Un:xB�)� �q ��ԙ"?&4�RL�If-#�"O"�����8AR�XU��Qn!�"Od�S@&V1P����E�e��"On�"�I�\����b��p�|1a1�'�Ov�i�	�>n!x��7`N�x��+"OT@&e��$H��/Y�h�t���"OZ��(_�&����3��)0��1��"O�L�D��z�XB5$Y�+���2q"O�t���;��3$WM��)��"Oл�E0��Ⱥbd�1.h0��"OF|yR
 D]�(�$I�4Pz�Rg"OtPU�č0�(Y��`Nn4�2�"O ���aԕ<���y4/&*����"Or�`� �n���-ʣ4�hD�"O�����Ū`�m��́�qL$Z"O�81GO�'��%�t��q��i"b"O���bɁm�6�ìA��R5K#"O���a�ۤ(g(uJ�di��p��"OޘQ�!Ć�BA�c�Q4r���p"O��P�OJ�\�" �3�Ǌn��Y��"O��S,��P�޽����\��y�"O����ݑj���
%�	
FMr�sR"On�#Ь�*x�I���C�<"O�ݺ�
�f��y���;9��y�"O0
��
4��UJ�o�*/ۖ[C"Of|���� .�tHb�φ	=���"O�xH�&М`!���flټ5�ܹ��"O�5��'��'��"�,ՋJ*����"OA{r�Y=(�1�G�#�%"v"O�\�&"JT� S��3/�*�"O��BEc�;:�J�d�'�d�2"O ]Z�S,A6a�bK�
ݰl	�"O����a!?���㒊�X�:�6"O~T!�� �^	�d*���� "OR!�Qeʢ9��pw��"%`�p�"O��k��Z�-d�%�H�j�rA"O�1�0Iù��x��2.�93"ON��� �8jg�O&s4K�"O���BK	~M�Q��<�6�S�"O�1YrhH�rEc��hO h"O�I�BY$� ��A9�Q�"OV�7a�M�(�
vF��!�X�a"O��qĭp����F�*L�F99P"O�ZP�Նf�hդ��=N+�"O��(S��b��({�i��OG���u"OlXDS�.��B6�P#e�ڑe"O�Pu�A�|���Uaݤj����4"O
d@���j�)�֜ ���r�"OH��+I�D���UO�$��j5D���ǅ�bPdH�˚�X(<7!3D�(g�˰| A�B�؀'S��PA2D���3� oH����$U�
ص:�/T��K�a=�h����
$m��g"Ox4:ǋ\�y\,Ôh5x^�E�W"O�4����,7�*)Z'��v���"O��0��*EpL4s#�� sd�5�"O���p�ډQ��a�3St�e"O YS��",v�ۦa�5:�|���"O������y�ҬCܢ�"OBo�{wP�qT�Zv��p"O�%	S��[�H�:$cӖ3�:ݠ�"O�̨e愕v�l�q҂�:��"O�E��,��x�CV���)��"Oj�ٳ�*)괻���r��$ce"O� D��r�#ì)�AT���p�7"O��h�&DZ�q��#q�@�*�"O�@8֫Q���A2��Ӷb��4#"O�9����:8�Z�Շi��aI��[�A���۴�?9ٴt��O�{��'��'^���C>h��8�]>N��Af��~��\"����U��ݦ���؟��'s�A~�yY'�6{����Ω$+�MX'a_�F��뜹S�6$K�䛁uj�?�w�t<�D㒐�\x儗�8�1+K�OJ8m����X>��w��sa�U�=0�졗��;:��QO�O����ƄhKd�k4E��Y"w�)E�[�@����	2�M�'�i��'���O��aF� ��7�ʟg��%#��Ǐ	���:8^��H�O�d�O8�d�ݺs��?�ٴWi~ �����lh����/L����x�ϻ5jtʇ#G6�a{2�̴gI�u��M��R/�䲔dW �Ť�4'�\yv�é��2�-�غ��!W�`i���)�d�z�Huk��
�AQ+�/�� 6�?YтA�`Lh�'��eݕ&�\B�Pm�:=	%��.Q>mk �ҥ�hO?��P�(�l����*�~j�(�:j
]��4�?��i�"�b�h��|��.G~�f�i���)!Pv��St��,R>)Ǔ�?�gI?�x��o�>BJ��r��F��tj`��Y�����L����!g-C�</��GyҦG�6>mqQH@�/�8�+���0;:v���ϟ�8_.����	&`a��aJ��6��D�&B��i��#`bI1:0Z`G���m�T@�Ѷh&����<�����'f�'C�6� 3�ٛ��,z�����6,�B�I!;�PQ���aN����W�;|`R���h�vT�0�GL�%�u��'�rY>�
��ҮN(m��YW�C�a�P�0��O����Oh��+�3]�(�'�P>��=<�����3v�q��)-Sd��>ٱō
D�h1� �&k��Lp�bI�v�r��?�3�NL2=�p�j`B_&����%x�����E;ݴ�?�J|J��	�ܨ�H�
<8���h�ⅦD��'�Iٟ"|�'Ƥ��և+~����'Lٔg��t��N��lhӼ�|�d|���� ^��%C2a�����'�X�"G�6�OR���O��:o�H���O*��}��ŀۂLv��@n��U�1����oo�i�w��Ӧi�żi�8�'��i�j�7p�)���6?(�"��f	�'���6�J$�!�P�D���$E_��H��Ʉj���-�
0�d�r��p[Mh��Λ�+�<�2h�y��?���sJ�H�3�W-��)���E��(���'�ў�I1[��8heCR�$D�`PF��?�ĳi!v6�8�$��p�)p����$�;Tф@(V���l��C��H3sL��)�RI�	��|���8h^w^��'��fC��F=nd�D.�/�X}��/ÀF6�
�e\����	�cl
��w苒HQ�q�u6}�3ƄV�|���0T@�T`�ug��;�=/�řc;����~�`� ]�_"t	�EO�,����?��i+�O����O�O����`�0(��5A���
<E� �UjXVH<���Ȅg2, X�!����p��()�6-'��Ħ��S\����0?� �  ��x�H1	��u���'?��$�ZX0��Ti?�����s�%�w+�^E��œ�?,y�E?�I}{����j۹J��з/@yξ1�ǉ}�Y[T��;_��X�Tg
8N��b��mVqO�`��'M�7��g�b��h^�&_r� ��Y�q�7��e�p�Ob���O>˓e`2U{т�[��l�����,�Rt��I��MSf�i��I�\'aB#�L�N���B����t��ٟp��b�	U�'�N�I @ ��'%ʰ�B$�������?!)���]�'YH��` �7������8Tb�0��{�y� �7cBdr�O�;)�hX�G��8�����*K��a�A+�7st�P��u�88j4�I*�M��T\?]��)M2,���	��A#pH�xW�����?!�S��򄎈b���
���F���Y�JE�z�!z�|�l�s}�g �(�xr�Aޘ2�.(Yd��~�'�B�|2��/n���   �2�ߤE"�jUKPk}b����;4WN\�ǄM�y�ƽ�5A(6�&��	��M� �ih���� ���T��"F�����BW�(S��Oj�d;��㟀�Iҟ�'P�ҩ]�3,��Ҕύ�jp�d��Q�r���q4���t���a�/2�n,O�p3�˅f���d�O�˧S� �B��M{��
�nдa���z՚X�FR�'Y�� *.xE�F(ĭJ�f��̦��O��ֺKq&� $�@0�!d�	[+^i}%�Qx���i�7j�
�Y�L�T�OK�""MQ��дՠ���=��O����'-�6�E����V�'
�P��@�mbu" �S>p�u�O��4��M�U�� �Dĉo�h��G�!_V�Gy��'�*7��ئ]&�̯;J� t�EřQ���F�ʤCTV�T�'�'fay�HI�U $  ��C���081�f�rsa߿�Z#i�$Al����L<��	̔F�J�4��뀰0PK��_��6m�Ky2ą��?�}�I˟�oZ$~ju[5Q��8,��_�{�Db�| .]c$I	2��
kP��/@�Y���?��iH�6�7�d����I�>�R�׳- ��GHQ�ܘ��@��H?���/nY`  @�?�ZKJ)$��,�!�G�mO��%%���f�F�!����FL�?Icb����O\�l��ħ��	\�x��%BD4̱��h^	-����?��S��y2�i8��s!��舵�A��#;<��Q�'�ў�3�Mc�iJ��:`T>آ�L9'Xb�Un��Wl]�)� �(޴�?����?�'eS����?��M�A�"w@C3�T����Ä�;}>��'k?��&O ��G�L>�3�ҜD�.AbM�d|=��`<�lqx�m	�Ր� Z�/o��н��9�3c'�d'r�yP�N�jl\L���<[�2h��A��?IA�i��ʓ�<�E�����"-]�� �3#�is,���!�?	�M-,t#��пa����G�	6*"��H̓y�hk�֓O^���H7�Эq��,��[�qfޘ����/$
��	:����C�؟(������ɨ�u��'�b�i׶�j�Cƴg�$�qJ[�8��͛sM˾~S���sd
)˴��Ie8�� <+��Æg~���E|*=4����<`�&��<;���'�	vm�ɲ;wޣ<���E�Ez�ͅ
#ؒщQGڦ�Ӳh�Oڈl���ē�?a���ēy�6	��a�8��$�M2D���	\�z����\?�(%�E-�==	*5���415�Ż�4��|�F�O��ICȠ۴�Mr�6�3RB ���Xꔂ!���'5 #���'XBJ�+fre8Ql��0!`4FٛT��}xE˝�#�>�b�ƻrZ��+�ؐ�a쌡Ej�(����@���ES\�� �"Ҩ���E�Blz�����#�!y�nJ�$�+2�lɧa�,��	̟T�If��[�æm�� 	�?ۊ�BH8f�H�F}R��4G6�:sE�w��$/�z~H���i��6M�<5�=K��V�'�O���C�:P��,��dc�$�7Ǟi^��?A�jC&<���jU�ї]Ɯ!B�j��:��+��?�R�E�%�uӕ'?mM�p�>�Ƀr\��4�����s���-�~���]�J��֝,/.��f�F�Q�*L�vE�3�b��KB�Oul��M;��ħ,/�]��L-	��j��Y���˂���OF���O��?�UaL<A
?���7� �F�&��$P��lZf}2F�4��E 5�	�RVQ��F�/c<0���Ys��d�O��4�h<��o�Ol���Od6퍗���^�k|F,�F� p�<��`�r�0��i���m�,P�	�|�@�>aˋ!�p��ҡ-/4��Y= �d����x*��0�L�c��>1�§[�u�4�ޣP`���"���z�6�'��������se�'/8��*�u<L!���)W5��� ��?UC!cєbPP;unK'~��pB��?}�'��6��$���S�?�mZ�h�t��*I�W���C �>w8�'�a}2�ֽ   ����c�N��4fV�>ܤ0#3�E�1,,�Z.O���O���?㟌 d�R�Q�]�G���j���v���=}b�i��'��@k$�Ok剿i&hrc� b}i��<j��H�#����@��v��֟�	ܟ���%b]���D��++ߨ��'��p~�I5ű1ֵR`� H�r�sf_��IE�'�"m+�a¶*ń 8��@J�2����Yl��X�D	1�J���H�y8����c�OD*�� ?�Xp�2C�!�IJZm�x($�(���`�?�O,�H{^z� Cbʍ	=�|1�-q��䓁HO�-Ѷ� 

��%9IP�Yg�O��o�M�N>����?�L<9!�B4 .  ��
82C�'
����O`7mC�>�t1F
��Q�<s��q�6۴Lϛ֛|R�O\�_�I'�Ɉ:�5C�	�vy�MYU-��t�׊�$�Iܟ��I�0Ϣ�	��@�I�>��x"+R������$�B=@�+rr�8��5IQ��q	�
�9��=`8����E3n6�\�1�՝��)!��P�q������A�I6pd�Q��,���[Ӆew���e���ē�?i����ħ;6�U�ԏ�\��ʦ*U5D����~�'��@��#]r06'M�\l4���'��6��æq�'#*��f{���'b�OBz��� �WuT�e��R�2�{b�'L�9j���$/ٜ=�Qd��7�b��C""!Ip�q$��I�(1�ύ'��P�v���(Oeq��YoB�0�a���f��&���&Ν���WG�Qpb��j@�b6���;��<Yp�O6�o��Ms����)��z6h� a�#��8�]�)�"��IC��?���jl�Ky�;e��H '&�6dl�EHVB0E8fч��?	ܴ�M��Hϐ&�Ɛq!@ŪvV���ez?	wɎ�"ڵ{��?Q.��тn�O��}�<T�G.Z�Q�p��Gz�����\�JuR�
ӥm��\o�-$�V\>�O4��I�{��ɢ2��DdmA7 �.4�D7��$h5>���ʹ��RG`�5֨���B�"H�B�S`�C�]K�}�3��MC$)]Οp��4U��&#|n��~B�-�/Ķ
���b�#��Ɵ��?Y��DX!m��M	E�ş&�L���J�i�qO���
˦u��4�䓆"\w��1�D��6G�!+���/%ҊDK�)0��$lO���
�  �Wf�%mqy�B��(�0�'l\>��v����V��v@r��&`_*��8���O��?a��fE(u3�n�;#>4QݴQ�N6��|Ҫ� 	ɡĜ�nh�����=2!���x��P'����o�9��2�FCT�':�x`B�b��p�P��eњs(fT$�<����Oаl�ħ��'sx-b �MZ�b$�Gb��}��q�=���'q�'9h�KUFF #�����%��C6��|��i�*7�<�d#/:�4+D�A��T#�&� =���	��&�pG~�@e ,  ��K�V�B'?��l��Ɵ�INyr�'���b<�%I��ZUkpǞ�7Iv���I�,nZF≻R�-�M�V*$-cT(W�xx����2�?)��?��ƅ;g̠���?a��?Q!���|�Pј��F�^ "�����	X@	B�-�MC!�h�,(A�lO�a���'^ qO�5�����Ur��O�
�i"�Xy�)�m[���|��̄Ʊ��'v��*fE�1��x��j�_��pd����;+O�"��?���M��G��:��K� ��!۔��/��OТ=�O�Rx�jR%�NU��H�_���x�'��JuӰpo~���?��o}r��?ZAZ��.@:� ����
�~2�'�d�k�  ������'[����)��רOV�[7�'N�7�d?!�Z�bz�0��Ɏ�TmҴ.�O?I���?)���DHLq<�P@�̾��9h�σ���IUy��i>�X�IA�r�귣�q�R�ׇ�g0 [ش��D>A��oZ���I{�
��̛�g���=
2�ʞ��aI�y����O��03�R�$a��p�'�rT>=�Ob�bRBA=>�\1�ga���8K<	���9l\ �#� !r/���$!T3|�򔯻B4�T���?���"XOH��CwLN<X%�t����O�Yl�-��'��'d'IC@h
)5 ����P�zi�=���<A���&���)���SuȰ�& PY�d��pY1O��oڽ�M�K<�5'��O7�	R�+R�*)�
��YNB6��O���O4�0�֭3�v���O��D�O��X`�
�hcߐ'�|�!��04�e`䌍�F]�� Q�i6B�z�����Ѹ'k4���_O�8�A��1��]y�@��9�"QH��C�+T�s]��O�;t�Oҩ�1��)7��(��܌{��a(�,��M�dZ���Oq��'���韲P6@S���"�ِ.�m�|����)aB�k��MA���
l���Q���~B�'��6�����$���?��'^���i
:�&���ĉ�D�9�Ō�G˂��P��O ��O���Ⱥ����?	��3����aA>BȨ����za*4�vN	1� ����=tȝ�d�'sT���ɛ?%;�!R(�R�X4G��gR,8�f�)p>��"�' V`��)�!Z��"�N�S����?��i��O����O��O~6�@��T�ZTEͳ
��j����|�xR�ɲU�� �1\!�|��� /%��O��mځ�M�+O>xP�
ڦ���ڴ�����U>�@�4�W�4�	G�	��H�g���s��ѫBA�K���ȇg��̴��M�T��sh�� ����<I��<:�����0�L��'̰���� )ڝcn8�
�L�v�	c*��]���E�	z�B�D�æ���4�MӠFہ�D���/Uxh�h��b�	�|�?���?1��M/vf��A��+ zp�`e�2mw�B�ɾ6�(py�kb-�����U�ǦI�R�B��M�.O�$�6�����OHʧJ��d�ڴr�)x�AW�/;�u:�E��V4H+7�'|���4��jT�H�fhB����O5���T�}�Q �=�=X��W#�%�x�m\�墕�0�0��Q2�&�?Hga�,�������A���#%<�ğ:?B�i�bp&>�&>%�t�Y���q���
Nd
�9�	ܟ�?	J<��	!v��;���)~I�v�̹|�ў�)�M+%�i�'��u"'��{Mм3�.Z7}y*(�G�O���%�D0�W��` @�?���MS1�'�>�S���8x��,�A.�&i�@�D�)A��9��iQ��-�
]�ɻ�A9��<Y�K�(���s��^t,Q�F���?���?���?���DզIA������a��%K>LI���IR-:S��O�#��Cy�z��	o�#�?�kN*��mCw] ����r���.���rL1?�D�N>JB�-� �ҽ��'3 �J�G�*��D�sZ�M�����?q���?q��?����?��iܢz�����G�;�&@���*/k��'�"mf�����%�<	���'r]�l�dpV#�͐�P�Ƹ�2�'��	9�M��iV��o_�0���O��Q�D� ��`���ڨe�Ip��$H((��m�7
=z�O,��?���?��	�(�hS�#1&XJf$LO��hz��?)*OHn��˟�I�p�O]�]��� O>�!�5)T?MK�89)O �-/�v.g�`l��O��g]ĸK�Nɣ9ϖ�t�U��exV�G��� ���VKyR�O���	�$�3[F�'���J!����C�Iݖ!��I2�'[b�'���'A�O��ɞ�MS��ğ5��uI��X0pBUpR,�70�j�I+O���)�	zyjq�R��nٲC�t���ȯ4&�����֦%S޴f���#�+�V~ROٓU��$3-��&�Z=a���C�^ �p�Fj�T��<q���?����?���?i˟`�j���]E����X�2�dͨ�b�J8����OZ���O蓟�d�O���5l�,�c ���-\�q�`�n��M��'��	|�ӡ򆉸7.���3ܲ�sc[�G�,W����	�e�,��;|��m'�$�'���'�\����:l�Ja!`x�´ɥ�'���'��[��c�4��8���?�m\���U��n�@�`�7C�B�0��X��	ݴ��b�Oz˧�A�4e���e[ F�+
@��'"v4�&��़�r���@
�7�(��;O��[��@�SB�3�$F7���'��'�B�'��>�Γ?@8��S�+0�%Z�`�1C�	�	��M+qe����O|�(�'��$��'ק0I�%���*m�@�I�M�R�i�6�W�1*0�d��� o^�X�XC2c͈Sn��
�)ad��6�P�$��l'���'�2�'���'�r�'�ժ��pe�U�G���wyD9�R�|q�4b%����?9����<	�) '��銁'߀j��DK��)��$ǦU�ߴ���S^�Fi��h�>��(�ώ{lb�Rb�&j(\��'"�r�	R��5r��|�T�,�6K~�A��/Q�T��1H�� 䟘�IܟH�I˟<��qy�"q�:��g�q�<��GޚB��(ր=]�'a�O��$%��~y�lӎYlZ"�?!!� (fʈ)��n��T�FÎ'.�q�,7?I��_
=O@�1��1��'A%'jV�57�\(g`��[�Ъ���?Q��?I��?a���?9��i[�����/ 3Z`���E�XBr�'�"�e�.�2�<����'x)�Gg�Ppt�5kX:S�t���'u�ɘ�M3�i8�n��)i�O~B �j�푰e
2T�^��s�M�*�%;aEP:5]��A��'V$# ��?�S�1U�\�'`�P�(K�{�Z\��ٱJ\^�*F扴����'D�z0�U3�d��hx�8�A��t���F`]8Yt(j�䌾+@��Y�~P��V9���Z"��ur�n	�����m��/����!�X"m��0qQ]�h���� p0 �b�-;���3KP;�h��IiZ@��5�����)<OL�����\�����  e`�r�"O����,sf0{F)l^��0��b���gD�^r��b��O-p�h�`��=P.�Kd$#xv�4pC���"�҃�=A,��6e�(>&U�v��4DB�SCO�Y?�B��Q2b+�� �+*��9�`�"*%v�����:|f����6<jl�D��D {'혰G6*%�p$��a@���hr�����O�����@�'�����e��Q���-��z��?Y��nWXb���?����?Y�'���N�t��y ���>u�~$�D��$N��I\�>�oZƟ���П\��9��'������s36�Fg�	@� :��'>��e�'bR�'
��t�'7"�HA�`�p^�a07GG&L���д�h�����O��Y�m��>I��yR	�,H&���)�za�8��B��?9��?���Ol��1(���$�Oz���O"-#�͑\!��U,�6� SJ�O���$-˒e�>����Gh�)��̄,�� �O�2Վ����?a!�J�?������AW��G�nM޴)#�@�8�����b�Qs̚<�L#�F;���$?ْ!��ܟ<�I�@%����"ԫ�8�ÕmCP8��O�ԟ�	蟐��ş@%���Op��,x<���}��M"/�\���O��O��On��?擡O^xk�-�8���C��[�rB�	ȕr�*'o�b$�C ����ݠG�4�8rh�����f� <��޲7���gnJ�jU���SB�'o$��۰�'j��d�41l,R��դ;oX��hG�^=N�Y���FŠÉר"�\٢(�V����S$�]��Ğ;������eQ�>��$ ��2`�PCf
�2>7T4��ـ�Jq�g:�G؞H1��(n���)�ɓ�8�,�X�8\OTD���ϰ>H�z�%<���=~�wJ
r����'�X�q�Ǎ\�Reɧ��1p�����'$�ݸ�oQ1L�!g��r6���'����	F5w��E�!�w*���'�$�zE |ԂRW�{��P��'J=�ri@:,���R�}��M��';�u2�恜2�&���Ul^��{�'z��d���j�Ru���e����'����ᎾU[Z�12�Ԗ+��P �'w����ʙ(F�QWm��q��)
�'8D�sFN1ư�k�aӌ`O�ػ�'��Qu�L��z��5_��A��'{@,	aA	-X`��go�9]גM��'.
�8sd�t"��A薕��I�'9&E�fڊu�\��"V���Ĩ�'�6���dK�@Ք��W�.s�BP��'���;�!Ǖ=v�;�*Y�i7lEP�'�.�c�*j*~]s�ǵ[{`� �'}4*��^0�i�
<GK��'9�ixW&�q�f[�H�#��'��P��>xe�}@-�#��}r	�'r��AG@�!;(��@�4/�l�'��dd�{X�1�  %�����'l�K& SC;��Y"�ξ��u"�'������M�l�@1a�_�0	�'ͪ�[s`
�`'��W��%if��'�D�[pf�e��DӇ�
<�E��'������Ψ[��m��CKu*~M@�'{�P�Shۗ%m�����wBά�
�'�V�qWFY�����]�S16�
�'N�UB�Ț h�:Dhf�GMd�S�'�X���cF'FM�V�6N��R�'�$Ȓ�\�2��0�)��7�pt�
�'j�,���F���;�����A
�'���.9cJ1�IR�BV�A�'�v����L b����%źhh���'�t��F	N3��Ёc��<Ё��',���*4j^��#��.S"|�'��� i�)�,�q�ʔ5y��z�'0$�H��ӯ4�(�������
�'�(TؑGG<"�ڔ8�⁁y
�	H
�'��1���a]q��M;��	�'}�`���
�k��Zz�X	 ����MT4�J��� �$���Y'_�틑�� ^�lT"Oй�N̗Ew~1�'��<�����i<ԁႈ�g��|�O?7��I�X`* ��9_.YR碚�"U!�䀆,آ���H�%?��Q�W^�$ͤYA�8�a�������dK� �.�'�P)����;�a|��p����e�|�`���d8t�"�uFO7����J{(<�2��({i��Y��O�hڀ�d�,ʓA��ĳ���*a��y��/��]r �he�8;Lऻ$e�AӶC�	�2�.�r4h� x��8��Z�s�&	��C��h@ gو���D2�g?����" �2��6㶨:5"Ob�<ᰦH� ��M�� �7C�F�J�p���6HkI�s;� �ቒT,��f��>/�a����!g����dڦ~�^4*�l�Q&uZ�N��21�E�#i�V\2Q&� C��#Q2��$��
�R�C�k�6l΂���-YB8�X w	٥_��|z@Y"u7���ph(��KQ�<i!܀X�x��V�M�NC�E��h�5G�-��(�-k��T�d���PG��'߂�8g��O���󔄑�d��X�'��LҪ$�>�3�EJ'T�����.�
B�R<UQ�P���0<�2�ſ2�& yÁ�*ls��z��s����v�ܪS)�����|m��Z5��;�h� ��-]��T�FJn<����b]���r$Мdvp�"'�Rb�'�bEzt�aͪt�х�`�'�V�� �$QW�p���P$d�t�ȓ	A��_#M��D�]�W������3��I�ˎ@���)��<� E٠l��x��L=�~E
�H~�<�!�� ��-YE@V+*�ٰ��z?�'ɫ �P�xA�%�<Q� ��H��-*�a�!��`���uX�L��Aj��@tꇓFS$��L_�:z��A@��u�����85�*�㥭@	)o���c�Ci�����%|�Q>I�`�H�<����I,%����-D�؛�L��-_��q�ؘLި-Jq�+D�L�ӓ4�y6+u>���##D�|�RG@9{WV��vl)�d%)��%D��!FL��|(e�G��h�@=S� D��1�q��tɗ��z�R��!D����R*f�����$���Yk�
=D�L+!J�3V[�I��ԭi]�p���>D��K����nľ� ��[�$�C�>D�$��mX[\�}� �V�?r�<��<D� �5+��i���e��PΒ��5�9D��Y1�C%;�*��v�L�{����I7D�@X�FMOAv�!��
�9O�0R��1D���@�1#m
pb�;|D�X��j D�,s�^�l�4��&�ЭA��+&h*D�	�Tn�Q�!#� ���'D��Pt�N'0м�e.ͰQ�����O"D�,����8�>��ዱ?$�;r>D����Å�C|ƅI8V��ܚ�e>D�������J��l1�A8�D;�J6D��:�,�(���$%��-L�{5(D��!�'��ls�C8n�$��%(D�8��,��Di��IU��F]��"c5D�੢�3qz��3�؀U����0D�x�2��,�y�gΖ;A\�#��1D�d֬�=QHh��f`�M�<�C�C.D��J�oU2Q��F�V0�5���!D�t"�#�/l�8$���\Y�̳dd<D�PׅO%kv(I�Ҍ�ظr�=D�h�*)9L ����`��'D���<o�°3��R<&Rp��o>D��#���2�p��Z�ą���:D���s��|�����1҂�94&6D�$��Ə�dP�uqDW?R�a���7D��JРK��J�2�4�Fe3D�<P�
�{���JլS�L\8(K�e1D�� (`3G	�'
�	�(A�kX	!#"O2��1"D4r�p�f
lLy)#"O����c��S���h�Ǝ�V�:P�7"O���t-��5npI��\�(�
��B"O>Ua�lѽ�,���!U:0`�-�$"O��0CR�_�ȨI"�_�R�A�"Ozq���v��p��oR T����"O&�`N�;�����&C�8���"O&`q�܌3IؽB�.ҿC�4h�W"O.RC��S��i��h��H�D��h�<1�B������A�4AO2����a�<1bN^:�������!>�`��b�<A��:�j�*��ˉ ������A�<���~f���BT-1�n(
Q�C�<�Ķc��	� E*I�V���'Jw�<i�A�+u���&�Ҫ>1�1StJ]F�<a�Q�F�� 3�8c�F�:�G�<酁
S�,�ʄ�`yĒ5�}�<1�bEa�x�c�V�8`@2�,�~�<��\�2^�`�Ph�70�`��u�<9�l~^�U;s��)3���1�%�{�<!��Ǥ\�Tq��J >x��C�o�<�A��9��P#wn\�.�QY瀉f�<��� 6��$r@�_3�iI�`�<9Ĉn �@�=ZHy"����z!��X�S��m��C�0�@����[�!���4<e┫ť�#mg�����-!�!�$� {�i�ĈH!}~��R�V�!���}Fh�r��.~j��H��Ɗ!��H�o�褥Geb��[6㊭5�!��U(^>�V.	�Ao��Q"�W�!�d393������x�䁁:w!�Y�<Р�g�D�A(��d��|�!��.]�}��$.}/��
하9�!�d߂@�����ք"�J��U�!�$�l�m��E�(�ސ���-�!�D�"g0@��.�	e �R��U�g!�_7-̶��S�/B�=C悑-f�!���3+Rf5��n	�I/D6��!�÷Iq���bV�N�ĺ��t�!�ą1g<B(�@�*j���!���AP㟢}J!m2|���z�j�m~�Hd�Nj�<���[4H�5(w�j�ua��Xf~rNާ2��뉅~���7fx�D�I�|G���D��&�8�sfF*`*�&�G>�p� �]�6�!�dH�99���� +ݎ}��C�t?�1��ƱqQ>]���\+�!��(5���k�' D��B��"��a��*^$�b6kt� R�O�u,qO?�t�6(�e���^A` azu�)D�\x���J!ܔ ȝ�����*?9�P�(���$�F�P�pAe��\�:,hS��-X�~�%Q�����P}�4�&��0J04@�0n��y��PZ`�1bUb�>�D$𰋘+�y�&��aT���c�<KD�맨T��y�$�[���Y�Ks~�x"�F��y�MԹ+5|���Q�ޘQB-��y��_�l�)� By;�d�1�T"�yr�L�zކ�ac�֒;T"�"����y��0c��۱��+a�x�'A,�yC����PY0/��Otqw��y�b�/)���3�N6;�@���yr�l1~�d!���%[���:�y¦T�;e��ˀ+�6}E��ulF��y"�K�g���y`^*8k�����]�y
� ��[�Ȏ�I�|�x��Ӄ��ɺ�"O�؃f�7T@M��U�`� ��r"O������-bYE�,+p��:g"Of�"HH�7��͡�S�*���:�"O���G�c����3f���&���"O�]�NF�$�T� oB1Qh�*�"O�d@��t�T��( NU�@�6"O
�S�.P9;�x�0D�R�PAC�"Oh܂"Þ=\�����m �w�d�1"Obm��˰+�&����E$?B����"Ox��B���7~�H�"+�Vu�s"O@�h�a�%B�D5u��4�T
_�<A׈!e�`თ��12��h� �U�<�C��X�<Aq��H�\����n�<)���7�����Ӣp�� �Hi�<Y aQ�A"H1��H�5���H��y�+]"5��A�BbY�;�=Un/�ybA��g�����1�:�St
�'�y�dJ�C R��5���{qH9S'��y�ؑ
t���R�E6t���@Џ�y��$y0�!�Fv+BM���� �yb�-���r����i���!����y2)߰��A���Œ=�� C��y�d��� &u>А�L�8�y��I�;���Zъ�n��$��	דq,�Q:��S3�zX�O�Z�:d�sM��=�Ȉ�q���B�	��nq:@/V�1�̱� ���jIVB�I\>�M:�#�J"l���v�BB�ɨw���i��)�4�p��U�D.B��)N'�9�5���$�9��Ӟ�C�"7ƽ�c����n��1���!"O��{�O+3R�sH�0�����"O��z��I�dj�+ǴJy�Mp"O�H����C�~�G��f����"O���e���<kTIy�&�Q�<���"Oȩ�uD�/.鮹�hَ���c�"O��X\�Z0�,�$��!��%{�"O+���!d*�����a�A�4GL`�<ٗ�5r��Y�G�#Q8��)��\�<����	!��K"���E�Uo_�<'�ٱ~��$��,L6;����Y�<��	+]���9��X��lYa�XU�<A$�ڑ$�J㰁]��P�N�<��\K� &��,$��r�GO�<)�~��}��%�� �����Y@�<��&H��8�&OKn�L��e�{�<I��,t�xIs#MF>.�Q��x�<�PL߁Nh�����l�v��a�Is�<�AΞ�l�W��E8�90��l�<	���H~ɓ��ޘ�
�y�h�<A��%h������A&�|�Đc�<�3g�/y��(jw���Dm��g\�<�G�J�c^�=K7O��}�.a�­]�<�i �I˒�[�
h�4$g�S�<�� �-n.�P���.X����Rj�Z�<����$���
��*Q��X�mDU�<�C/�	D�H=Y��K�5��h�j�<F圛_�m��	U95�(*��Qg�<���`�d����0,�Q	�b
d�<ᦉǱ(k�͓d�ӂ���1��D�<���DH��}SU������`qn��<���!}󚁓1�PcI,���"r�<��.J��PK��(��9@�Tg�<�kB-+�<�P��I�P��)�v�e�<� 6@jV�h2������8�B"OxT�U@�,D��{�H���"OV1�N�ntܽa�"\���v"O�����WE��d��Q>f�%�I}L��G���5W$��)����h9�@��yrDO3 x�(�6΄�l.�r�i*�y�˕#���=E�t�81��h��#|dSs�ű�y2�B�F�R�� %ڻl_T�.�+���6H^d�Ԭ����<) Bj�$�@"�N6� I�u"v8�� "iϹ0�A��+�Ctd11J�qZd�Sf�!�ɇēcv�p��Xyc�ԫ��ٻ:��-Fy�Dǒ���s��@+���!���7J�����P�7ߠi��"O�}�v����q�6I���i{v#�'�*	��S�)֧����H�
�RT��M� zhF�u#C*!��׀880�zrL�L�~��CA�T���Ga�r��\�}��	�/�����Aմ9�8� �D��n:>���[: ��� ��O5��'�M�-^�X�����8�������x2��a>5�w䇴͎������'|B�gK>�}iV�0�S�	m��Qǃ��Ox�qk�
X5��C�	�Vy5z ��~�*��
7�N i�I�c�Zm��؟�~r��R�(P�jE� �ÂA|�m&A9D���s�ͦ8>�1�2�@�|: ;3	�OZm���Iۘȡ��Ӱ<y@�ZF��8��((�Y���k��C��?O6ؼ�N�t�|x�!=x�Ba���4-�neH	�'L�5(��njt	`
�3i�R�9��$ݯ3�4+����c?MP�n�^��d����/|;�@9��1D�$P7���x)W�Q�Cl�ȸF�O��ע����T:*O?�D{�AP��9[Ρ�s��!�!��v�.hr��U/v�F���	�3���;?n���2�G.��y�'$d�lM"�	�:py�����0?�S�B�_� �W
 kP֜z�%6�JY�[h�<i�ޑV\V��u�Q�J���"�P}�'/`j��S:C�Dh��8ɮ�(3�F�&�C�I�!��*�ID�}x� !��iu�C�	�
���Y�,RO\�:���yC�B�I�:vD��S���?�!iR��.(K�B䉛8��I�(~� Ă�$<�B�	3N���s&	7�&��ٙ2C�I�}$J9@�� ^����-�dC�	2���1E�T��2�W��B��4� �"�!\�;56�FV�=$B�Z,��3ꛬG�Ф�Wk!]��C�6m���S�	�)
Ĵ�Ɗ��G(B��@����xqd�rc	�7`yB�I�*"�����E��J��̭Q�C��]���Q�kԖq2�������C�Ƀg �#D�2{fN��W/=�C�I�[�l�{v �.o"`F٦ ��B�I�kx�s���#�D�2�w�B�I�9u�`r�H\W,��$���mĐB��&h���0 ��6�F�4A,$�tB�	�	굋�3b�*H�V��r7�B�	 �F�5k��$ޱH7�Z%U��B�IM~՛��~g����-$@�B䉚9�튠�S�i�9b0⛃КB�I���4AReN;K=]K �W��B�E�P�A'�p0Bh�T�҅"`B�	A=@ۀ͔9hR�!�+N3>4$B�	�8���4�ŧ�Ɗ�igZ���"O�`���82M���M1Z�$Q�"O�ْ�#�:=�v`(��Y2}7V�@A"Oj�z6�ʽ$R sA�[�E#��F"O�)�4@*k
�ٓ��X
���g"O`�1���-w�Ly��Θgg�1U"O� ^tyŮ��>a��ƀ�v��l6D���ש_�K2*��$�
:)"}��F#D�(�A�D����J�IJ�d�7�%D�(��[��ܢ @K0����c&D�${t��U"  �K�$p��`��7D��k�ܞ@r��SF�1QD�C�"D��������Ad���6`
pn"D����ĸ=f��9p�1C	n�R@<D��(ҥU)d�j0�7ic�]Z��8D���7L�| p�0E�2q8N,Q$:D�Kb��e�P1��Y:g�
+D�t��'5� l`�cV� �����.D��:W�����i��ı`�i+D��Y`�L�FY��Է\씅�Q�'D��d�S�*i ��JZ`;qB+D�:P�O��z�i�*�z͓Ӌ;D��I��*k��l�qjBXA�G�#D����&K�Њ�/�=/�J]�� D�����b5�<)�@0�N�#�K?D��x`bL�S3<<sə!IZL�caM>D�dq5A�1lV��'J
.���:D� @5ș�p��Es�<�Jly��6D� c��76L4��Ϙ"oC�y�7�8D�ؓ�dΆQ邙be�
?�����M)D�Tq��
�fqYf䒨+nQ��a%D�|�VƘ?G*�]��fF'v~Bq�g>D�x�vI�(A����c����a�?D����Z�%1�l
$f�\v�4qn<D���9�TSG5���Q(-D�@��i�<H�J���EZ�ʔ�!�+D��z� m���v���?|��@�%&D�4����?���S!L˥[OD��G D�x�4 �Fȋ  \4i�5�=D�4a����b��)3����L�25Y�N;D��Yb�� ��Ñ,��f���V�,D���G��?��QƏ;q^�|�o=D��AE�P� PR�]zq�0`S�.D�P#�"�H�<)J�B/m�ȌA��,D�D���_'�@XSBZAݼd�An+D��Hq(
�K�5� �ҋ�b�g�)D�hrC@VdgP�"���.U�4M�w�(D��"�^SO
��sJXdO6%P�-#D�����W��"o�1JE����3D�ԩ�d��"���"�Z?o��*��-D���O�,i�ԥ ��Lu�h��0�-D��E� [C
1h�	,ΜP��`!D��pF�I�a�8��5�Ȍ^,�2D���w�ӗ@�\u��P�+D��"1D��z��("w� �iӄ<`�� .D� �Æ�/�d�Y��ְ<y��'D�L�b @40ޤ ��Q�bn��iT�&D�pr�?3\L(�d�*��1��H"D��C� ��@�P�(���aB�Eq� D�t�bOP��af��!-�HY��#D���r�W�'-����V�(e�V%<D�0��;TAz�(mڱ[e�<�a8D�����
�hI3=[�yj�(6D��;�<[X����lŨw�t[v(4D�\p�c=X��a� 0o�k��0D���O[�5(���6q'��P�*0D�pA6#'z���kC��D'�}q��9D��Ҷ���Z&����X! �؂�2D���eO��"uP�� �NS0D�D�!��!U��Kׇ�e�v8�3�.D�� �,�4�دimT��dO�Z���R"O���ˌ6)ah@KbO^�7ȵ�"OP��N\�-V�9��Y�r�"O����3ެ�AJ^�:���"O~���(��}* m����>%���T"ON� ����\8d	��Ɩq0��"O���c��fcDiyq�kj8L��"O|�Ё�z:B�i���h;��"O�5ijF0|��n$+��j "ON�!`���"��y��#�!����"O.}Qu�@:��ʴ�;��Bs"O�%�&jN+��<��������"O�Z�G�N�P�:o��}�V"O|5�Ed|��i�K9n�*�"O,�H�(�*xF4��e���{eHp�"OL�W5?ͬ��B��W���"O|	��mO2%SPD8���0Wqd3'"O�����>x�@lpi�iXI�"O�A�gY�1,,�4��e �a"OX5s�<4����"�� J��I�"OD�	�M?8�� ��VW�^��"Oإ�$�C�M@�Y��� n�v��"O0�xq���b�&DKt) "eu �b�"OFT�����M�|`�`�7?k�*�"O\�!�N�.>Z �j �oOڙÆ"O����3*��Py�J��#�R��R"Oxѕ���(���p��Z>�,yѴ"O�ԣ5����0
���\kʄP�"O��+W���!�L%�7Ζ3@ZD@J�"O:Hk�FVh8RA�҃V/tK��h%"O�Iz',�5I�lh�B������"O����!Q<1~��� 1_z�*�"O��c�Q�a����	Topz�"O"�����2r�aGc]�VX�U�"O��@��FP1� @��	�"O��P���l�.����U"v��x�"OP�R���#jIn(sD��/\ۊ���"O�XБM�+>V�ٲD�)���e"OM���ή꾤����X*&"O��Z�-MdEn�3�@ժ2Ll�b"O����l�>I�~���4�}r�"OX�A7��>�q`�䈛z�����"OTԢ`뉆R��=��N)s2RJ�"Or���S�j\X��Q�$>�H$"O�xR��R_��b���D H@�"O *�Й&J	"��	�Xz"O$��1
������Dΐ2$H���"O��V�N?�ܘ�g�G	@�b��"Ox��G� X=
A(J^;B�rp��"O(T��'Фb��h0)���ꭰ�"O���2�
�~���D҉ޮ��U"O&t�2+I7R~R���N�j���b"OL�i��SiPάC���z��d@d"O⥣q%�0B�j�%�T��re"O��P���q	<y�x9p"O�A@ �U}D"��O�]4��"O�թ�C��5$��$��,� �"Ox<�0ǏA��,��*�p����"O�#�B	-ۆ!�1R�1"O��hxR*�ڒ��lb�B�"O��ɐ�R������ �6��U��"O2�@�&D�w�|��.�oѬ���"O"�hS��	@��AvG�0_�RE9'"Or!�W��ST�p���Q��k�"O� �fa^3���d����"O:���%����[�(ys�"O�(�s�_v�Ȋވ|4�53��=D��w �ZB@���9���k��'D����L
5�8�B�f"�v�{f�9D�x��h!W>(�{�iݧ�Tm��$2D�� V RZ&T��/W'#lB9S�./D��BE��?3h$��K��;�Z��U!0D�t(ԃ\0D<� ��@�.�0�"ť*D�� �4I`�Pȓ��0	(.��2�,D��1�DX�u�"���3�: ��>D����ծ.�����a#HXӪ<D���`Q*T/��cTi�Vǰ)G&D���4kSV��a�ܞ|%j�qE�#D��bb���P����ءo�,�I$D�PC�l\7l���+�"��%D�08!N�o��8�&DUf���A�.D��G�$v��A���-*Qx��*D��'�=z�$���B#6��9��)D��ئ���� GA�E�d�'D�$"��L6~��I�AB�3|�L�r��:D��{RG��0)`LPe*�6)I��9�������+�`l�����!��C�"O�����G�l�� 3�I>p4�"O���R���p��2 ���J�B�"O��X#Ê�,���)/R�F�N�ʇ"OĀzQc �� ��'p����"OR ��ϝ0�L5a����}�x�V"O�3�� �pm"x��������b"Od��%D
b|�����`E�"O�@҃��/*�H"5a� ]��ke"O�X*�I�#q E�!+O%���K�"O�󈁚49P���o�5rց �"O�<���	h#�Y��DR!"O���G���;�\	��a�(�:1�"OR=IT�.;Ol�2���q����"O���d�שl(�H@�� g>�r!"O-�C�]//�Vx���+Nx�"O�9h��F�}C�hxƨ5`i�5"O� PF/g���Wen�=��"OPؕ8F�D�q e+WP 
d"O6���l��A"�!g�
16ؼ�8�"O"��7�V�	j�(
�ܾpgV�A4"O��3�kD�":�ݲ "�8¸��"O�LCb@�SȔQa�%.&�`�"O`����8>�:{& ��M�\�G"Oz�z�	!f�ޭ8p�tr�"O�੗k�?	��k4�غ�i��"O6M@S':-l�i���xU�,�"O�t�Ĩ �JUH��U�[pI��m(D���獱J�p��������C�,D��Sm7g�t!�OBg p���&D�`
P���d HM���K�w&d��&8D�� �l](��y赋
�ܦ�i�n4D�8{�A�Bd�)�fH+3ܵ�u'4D������ &�	g�X�.�䙘5e3D����s���j�B��~% ��O3D��(�`�!#�:H#f��ct,�[W&0D�p�2aS8d��k$�R�'{�s�h.D�H���Q�d?�%I�#�J�e�3h,D����	|����Q�"eʍ�7�)D� �2n�?���/�z�EK�.:D�`���#?�~y�e��:<V��d(:D����I�	 ��{��9z�zY�E�<D�� &D�W���x1A��& �"O���E ̮H���P��R�"O��;���7Y֘ur����@*%"O�H�g6c��J3ꞽ:�D  "O8�W�M��,��`�TLv4hC"O�03A�O�JVr����\�|`f���"O�!a$¥[*�$Q� �7Ga2�"O<@A�ҁ��5��i�Q�-�T"OrMs����1��H��.�R$"O���R�fr�1����sBYS"O�e�e�@&��@���E�]�
�"O��@5!ێ��掑�i$h<;Q"O�u���=w�����h/TY��"O�%: �Q13y������p���'5N�����)}����K˷u����'�}�r�Ps���Y�L"}5�1�'����$Y��lsgd�phf ��'��E����s�J�EB�j&��1�'���Y0,S"X��_+VX��'e�+���!&Y����5V/2�K�'zL��$ݷg�$a��RL0��'��i0��Bl~��Ɍ�I��z�'���C!kC�<x�@�E;Do�l��'��wk�|w&�2�D�;��@�'Ġ��!�I������� u�'�r���./�ZuC�X�v��1	�'�|(C�`�g���h�.�o_P�B�'Cޥ��L�T�!y��2vSp-��'$�=[S�Vv��P�&]�d�@�'cTu��N	m����M�/#G�&;D��`�7?�̍Rd I�Y�,pi�H7D� 3�� �
����ȴc����"D�ț��X$5�
��q�t�!D�$��+��R� �t�O] ����;D��v�sH�����k��'D���Rj'͕�aW<�搫�f��yri�${@������v���0�) ��yr���f� X�F޹�uk�kX4�y�F�e���3)̼Z��x�B��y�B(�N˱�C/�~$����y�,>(@�aQD
�}��[7!ϫ�y�랠q&��'�Zud]��֫�y��T�*�y*��ȜX��ׁ�y�o�)F5(\B���(��Q�o�
ػ�'q�U���ߕQBeː)\�;qP|��'ɬ�%*ó.$�8�e�/	�E�'�ԉI�Ĭ�6�+��C�$L���'At-����X�Pغ�/Ct�@�;�'-����,="Y��'	6��ȓR�PQh�U��P	 "�-V�X��+�N�jEO��{(�gë�t��U��\��A�*�?QL"��ȓY(T]�7�ؕR�čku�߽+\�D��8��Ks�8��x{Ո�	<��ȓo��1��M�W���* ���B�L��BV��#��~�����gA8j��$�ȓ�5� ��
JW� �� �2~��ą�"�U�e�L�OH����
�v�B�ȓ�l�jb�Tn��P�����I�ȓ��|�M�Y�� �b	�(�^���1�����+�>K�f�upC �������C��X�`
�?CD��ȓD�|�Y�K��^��ς��h���IH�����@�!�08cr
Ԣ����S�? v�6��f�P�A����6��"O8��Ð0{������5ЬEJ�"O��#�#�3��ʔk�����"Oq��&Y#:���sȆ��\�� "O`�a�%v����-4�"O~x���̘B�)9�眆qn��Y�"O�Z4C�#�1�ڠn�
��$"O�4�`�&�ds���k��!�"O��z�OČgj(�	@����"O>�BCO&x�0c�ÉlBR�"O�Q��#4���5eL 3���"OH�S���Q����e���iw� *�"O�� !�6y1VA��C�_d�- �"OD�3bq[�#��B]�9��"O����@f�i(G��1:��rP"O�I��X|����1 �r�G"O�(ٓ#۳n7�;�P��h�"O�y*QaEK5�:�Z��"Oc%*��1Hj�0�/ĭ�|���"Ol sa�'�����Ӽ��Z�"Od���UX�TD���Q/�\yF"O�� �L�*�\@h��67��<�E"O�cJ�P��5Aҡ3:��i��"O���Ӂ�GP^���&+M8Z�"O����K�{jl�"W���f��<
w"O~D�%
J�lD��M�&S��<8�"O�����F�[��AV���H���u"O$�`iN<(j|YS��*�%AC"O��q����D�	睓&�(�P�"O腑
�5�4p@��&�x�""O�5�V��1$� ��m��X�BP��"O� їD�?Ø �eϚ�v-�l[�"O>Uɲ�Ǳ"�l���nS6{(J�y"O�er�e ����KƗ8����"OP�ȶ�Zx���rI�~?�x"Oذ(v���X"���߇w��"O6U�u��-0=��Z���<bl�ɳ�"O"�)�@�8��0�7n�>Q*@s"O�⦢ϕ(��ȱ��֩_3��v"OX��'��~��͸�iQQ"TT"O��b6��weh-뷇q<f��"O*`��s�F1�&�m<X؊"O��	b -7�~`�"FÙ6�9�"O 4�w�_�$���#H49;
��e"O�ᣒĒ>��!PugٽN�ģ7"O^]���0o������u�n�`Q"O $	��4��	�Ջ�#���W"O���$ �	X"����k(+�2rs"O~�2�O=l	�� ��;��8�"OV��"T�T4`)Eq��uA�"O�s���dϒ�B7) �\>I��"O����e�,&� ��(F�k��]2r"O����-8c�5��j�7�`�r�"Oxh+��#{"�8@��)>��t�<Q�Q)?�n܁C��h�D��Q�<�Ak\�"fJ�Xqa��3��[7�K�<1&*��,v�آB9C�f@"LK�<�j[Xo�%@���w�EA��J�<u��7n��A��:C�P�I�k�<1%�͛$=���e�B�_#�DI�e�<�Ҁ�g��$sg&[Rd�s��^�<����R*ㄅ�=���nV�<���I (Q�D�s�D�'h�y�<��T&tj��;  ���U�0n�s�<� N�zw#Ł�<���@<I�D��"ONexrbD!)��9��IS,���"O����!��~��I���v��Q�"O\��N�!�zBjF�}Od�"O�a`)S+5�L�"㋖+�`00"OJHr	�o�*8AD�	�vq�"Oy;Q�ˠ�$�˵���x�c"O�����\�1���O����q"O��z�D�uI�E`ÁE%$$ZW"Od}!T-��~9���� �:�Q�"OL4����!���X�&
x�3�"Ox$a�K,�y oPW����g"Ol�i�a$6lfY{� �P��@�"O���S��=��܂1b	�>�^�ڲ"O��j%f �h��`Y�A�&h�[�"O<��� ��{����� ��.e��2"O�IQ�nj��+3TR�Q"O�5�w-�-͆T�.	�7>�Q�"O�
��ȇr?�`����z-V��"Ol�Pd��<�Ĥ��J�����"O�t���-*X���Dj���j\�"O@U�#���6�E��˲@�<�C��#��ź`
N/C�<�QE-MS�<�4!�E��DH�$ѩ�U��OD�<y�*�D��C�Ҿn�Ph��n�C�<Y�g����pmM�S&��.{�<�,��/���`�*̼}��3"x�<��υ�B@�%1Ņ��$y�TRV�r�<QT��
n~��� aNy����w�<���*,H���)�&h�!��k�<�6Ǚ�C���B�鏣#���ҭj�<�5�\�K��(sEDT�u�͓�/�d�<3�S�\9�$�Y�1(h��J�k�<qC�(6�96�M�{��kg.	i�<���"�.���
sQ�$��b�<�fV-D{Vx
1d��n�t��SK@x�<����r�ڨ�3dԽ3)9�N�u�<Y� �3
tm��]:a��ᨶ�X]�<����x����m��I�`�<ٶ	��~4�r'o�[��вe_f�<����k����OC�ʴ)�id�<�Ō��n�B-I�`T,\��;fN�_�<1	גO���Њ���1LBq��g�@�h%E�9l�DQ��ș|���ȓ+Rbp�!�\Q�i��_��d��ȓg^�|K�N��\�T�����]�*<�ȓ `�U"��ľ|m�,3�a8oІȓxV�4Iw.�1w�Y�!ܮ$���ȓ���S<N,�R�.�'
$贅�U�^"ԣׅ��R�T�R����9P����?r0a���%BԆ1��<��0�@%�n[���	: �!�ȓn���-�"e�\�{ŏ��V_���ȓq�j�P�
CG
��A�� M��ȓ7l�H�Tm͌d]���������ȓs�J� �8%p����#ҿ(��T�ȓ*�N�8��N�VZ�@@�K�
�ȓnv8i�����ј2�C��I��*�@���u|����?m R ��n�jL#ՊΆ*�v��tc��~�ȓk�d�����AV�u0%��MDv�ȓa�����& zm<��� T*2�t��McPhX�぀ex�`A�Δ�;�t���sg�В`����hs	�#er%��S�? �q(�"Ծ ���F�	�Tp�m*�"OH5G��W?���@�ТE�1�d"O�A� �V\��Ԡ��]		Dj�r�"OT�[��	y�,�*!D�7�IJB"Ozػ��9!�fQ;t`]*��`��"O�p2B�E�X�ȆDF4�.�q"O���w%�����y�Í��0��S"O�1��B�v!�W�K��.�8�"O�Ċt�@D=�b�J�B� "O��adb���H4�TcڑԈ$D"Od���̂q�4�@�5`z(��"O��Z�M�h�*�L�,��Q�v"O��@C�-4�伳E��8�fpCC"O��1lͫ<���DA�\��aqR"O�L��L1v$�n@�Yd|"O�T����	*�2�B	�AKdq�G"O2��a	TIĨy3�`�"Hp�d"O��K�;Cf��W��IA��"Oݪs�>ф��%cy�4�sb"OB�9DM���I��A�_�(,�4"O����'J&*�>�X#!�+�D��E"O�K��(l�Ȉ��-�=��` p"OV��h�\*؈����mz�@V"OH@p����TɃ��_�Xt"O J�:P�[�'B��`�d"O �+�bJ'C��y'Oִ	�ܴ�a"O�SiO$��(*n�!tr�b"Oָk󡛇e�.�J��B�v4,��S"OFX�1�Ŕ�~�酯��{x2"O��i������H��t"}[�"O�����̴������4D^x�8�"O�]�",}��`2`�) �l��"O�L�g-ۉ/�ލ 4�B�x�v"O�걨�U��qh���!�N�S"O�Y���� 2�rTx5Ȝ�T�ج�q"O*D�t�Ѯp@�xw���JW�]��"ODL�#�6����*��ec1"O|�yՋdb�-��L�T��l:�"O�I�Rm�#W��5()_f�́"O��x��mt��X��{E"O���1ğ&8���JE�S�lP�-ʣ"O8!K1kF=�H��bҚJ��ڀ"O��j"�=?hd�&C��C4���f"O����A��b�E���"O6d��ϗ�s�F�B���%r@e "Oni�ŬE�6Egn׾[�`d"Oj- T�#~�ƍ��,��H�<�C"O�����T�[�P���X���EK�"Oꕒ�"�A��)�ɮ���"O��Je�� ��!��-� (皜�"O:�Q��M:0l��:#�	�g���"O�}�΁�:t4�b�+ɢ��h�"Ot؊�hF�츻vj
�h��0�"O+�C��@h7� m{� x)�t�<��^��d�jSb	��# �o�<Yp(�-�h���X�]���C��m�<I�$a�駃�'9�p����<'dC�I�g��U�ݶS���v��F�C�	�&��W������c�w&B�Is�	����m-�0��]�"�B�Ig��X�$"�.��|0%�h��C�u���8�O�b���tm���pC��w���k�DC�*>�G�t]8C䉗0�6��L��N�03���U/ C�)� ����S�6`�U)J�$��"O�8��V�9�����G8s|�"O�p�� �,�I`�9C�m�w"O��*��8��b�EM22\�Za"O� C`Y���ـ��Q�{,�0��"O
@�����6���烑ABt<"O���`�?U�(��ȵw�hH�"O,p�ƀ���~!"�&O$}�H-��"O���(�4(����80��u"O���։Ѓ&U̒��	R��sV"Oly�a��#}h��3�j��]���"O�q��D�_���oQ9�ZE��'bPЄR�FGZ��c㘭e��e�	�'�� 0*�LȄ�0�a��a
�'��{��M�x|��W�ҥ\f\͊
�'�l��'i�	P�mȱ�O�by���'>�@0��#���ɁJ�(��]�'A�0�͟�3d.���h�?2�b���'T4�p�^��@�B�-.�Z�'YhT���F�B�P�f�,�����')��
%&lX�'H�+N<MH�'͘L��m�9X�p��3[�JD��'N�X�[3�dSW��<z�'!���q�m�s�{k����'��!������6�Z���H��'�z�y'��բ���e	 {�����'�z�e��
Xeq�@�x��Xb�'����V���{�DQVe�(C�MR�'�ث7��
��%�%��Y,A�
�'l��
:]Rl�:P"n����'A&�PY>`�܌�d��ktԩ�'`���f̅;<y ��TL�
j�T�A�'FN8��L�Svf���d$����'A<�{U��Kh�t[�'k^����Ib�@�D+�<Q:p��
�'�(��m�#Z\K�I��]�Zqb�'}
������4u�D e��g����'���`�[�z�v<H�cV�]G`�X�'��<��)V�x:����U6G&5��'7��P�&�0<R��y�hlq�'�N�sw���f��H4u/�i�'N`�N	��� �m�W�x��'r�
Z�*"���`AIq
�'�t�s M^.~>�-T7��Y
�'��E����G����60f��Z	�'����C*JK|{D��U�d��'\~Qpg.� �Z��t!Z=BsL�	�'i��B�ߏ1*Y��U�/�̬	�'u��Hd�I�c(�R��[z��`�
�'�D#̯ �nI2�����'G�y��o5,��{1���m�J���'��:�K
;�1���X�m��'m ����+�&�@pό�i�,�'@h�	i�%E�:�ʷ�4[��
�'���a�=,ʌ����:���+
�'� ����[��t�A�H.�A	�'w��;��_#���&Aϻ+v�[	�'���T��O�
�:�,	* �-��'-f] ���8�X8+G�M�}ߪu:�'�����n�/X������|�� !�'0�<�wEE���1��� �l����'
V�pp���,*��h�#�c6��'�ZH�C��;Q/yX�h؈)rT]��'5��g�
j՘��V#&"0�0��� ^�1�A�i@h 2�_����`2"OP��D��+�l�f�����"O2�����!U���딙&��b"Oڴ�ƃ�5,�VdY��d�"O"�� �ޫknu#�ȉ"y�M��"O��+���[�pka5v����"O����%���! @�"eT�U�"O�M0B�[��2���5DT��"O\�B�g�13�� `��NU��"O��������T�_ߪ]�S"O����W7azz�@	Q�s�I2"O���IP�'���A�h
�Y���A"O��3��	V I���N�F��"O8-@����$����%\�9�a
p"O��Aԫ) ��HuC��~%H��"O`�Kٻ��A�p��B"O��J=_�@	�2A�%:��`�"O��qV�ڛyoF���ͣ;E�[�"Ov�٣GX���ad'��<W�ġ%"Ou��D�',�XK�$��r��{�"O�(0���,���B�ے�h3"O0���E,�꛹Ÿ́�G"OP�cR)�7��`�!	Ռ"���"�"O�Źp��=^^½B�_�,�*��1"O(p�+E!1�� ���{�,"�"O֑z�e:#��٧fF��8`�"O��iZ7n8k�%�rj��h�*ODЃ%,���R!�K�,_��;�',��$
�;̮��ᅜ�;�i�
�'�f��V�Y����Q��(phC
�'m*�b��!w+��hBI�#};v�[	�'�`"���z��՚�g��^P���'䎰BU���K�@�/��a����(�y�I[�pٶ��T����"b����y2$B�N�E堅-^��%>�y��H���!AbC<x-��!��J �yr��+��{VĜ3v͎\"7+��y2aޘN�Hh$�^v�x���/�y�
�(~.$QAC# �-s��.�y��
�qf�"�F#"���s�hH��yR�f��:��8kV$)JSiŴݖC�I2C��'I��P׾\�� �A�TC�	�#����Mڹe�J�� �Z:C�Ɇ\�ܙ�Ɵ,_.k�'t.<C�ɚ�^������26 `�B����C�	��8�󫚄r���W�C�3H�Z�+&��W2����
��B�	�B�DԚ�.ɊLV�!�ՅI;p�B�	@���;7J_@O~ՈV�)l�B�	g8�� ��=z���ȷm��C�I�s�5	��3�@ZVA��hC�	�|О4"V��D�@q��$��ZC䉅r.�y3G�!�>�8!B�;zC�	��(}�U!޶C_9(�ޯ%�:C�<=Dz�3��lD�R������=D��b�
* A���,.gf���0D�DS#1a�x�1/5eQB��f0D��qE�O�E�q� �9H0g�,D�����p���Ձ3`���h*D�dK5#�8����&-�8[�����o-D�xqb.� D(��9Do�ڈ�S��,D��'l�n� �V횢S�h����+D��I��[�])����kTn�A�5D����O7R`R�I$�I�:|�1D�� :1�s���_�>U��ܼe,��"O4��a��+i�n�.��3��!i`"OTu�fd�3;pd��F�-MJa"&"O��� �&���A���L/4�Z$"O8ȹc���r |522%G�3��� "O&̡�&����A�Y1p�d���"Or�SJ�x�pT"c��.~
${b"O`��Y#�XM�v`F.Km~H��"O�@�o*-d�*e`e]N��"O�M@&#ֈq�n�I�Ω<LJAG"OP�J���x�1�B>0I`�I�"O�8�@�x^���"\01Y�"O����S�V� "D�;�.`�"O`racH�`栤�j��l6�eS�"Oh�RD��)�l8v'��'�@p:�"O`����������f�=�.q��"O��˧L@#0>���D���H�+!"Oz)�_�wni�g��8&�Y�"OP��ˏ�/��m:���V���C"Od���IZ����H��-@�~�C�"O�q�I]�Hv�T����\� �a�"O4���,.4(�pK�=_�L��"O���lC(�	1u̯�1��"O&q�
�,Q���!��J���`"O&�Q��o�,��7�(u�}("O܌�yk�X�&Ä�7hB��6"O�	#���2+\u���Er]���g"Od�p�ԇ~b}�O�R�A2"O,S����ekh"��
%a���R"O�E٤�
 '��3�jX1�V�`D"O���mݪo��L�7���y�H+&"O�8��d��f��sv�2/���X"O�i��r�e��!�:Vq��a�"O�Ͱ�K�X�<��@N�=oX�Є"O^���/[��P��!;J�pv"Oh=�a�
=nș��ϔL'�E�p"Ov�����=Kd�� �:?,�C�"O%��F�4�~�ݸ^� �B4D�LDH���N-he�.J<R�:S"3D�(�&��&:z���l�����1#/D��R�h�6Ѵ]� �^�I��ɵj/D��1��k^����Ȩ[<��cK-D�ty��A�6°e�!�Ҋ3�����6D���EiF�A�>p�"cOH���*u�5D��1ת�'R�����@ �d�R�1`3D�l��`�]�F��*H�!-0D���k��w�&ܫ+�>�<��v�)D��: ��U�6}AdU�� �*'D��J�+�$g�dH�\�c"�|�j&D��S�O4�<��Re�RL�A�Ն"D�l@Y���A솆bf5�K#D���t�W�p	t�!L�A�N�0$K!D�T{giG4A >a(I����$`�� D��A���^*r�10�	4Uh�t	�,D��ʱFU�u�� �1�Z�f~�Ѫ�E'D��HF@�5N��U�E+O�~��Ǌ#D�hB�/�^�BCb���^e���3D��(�J��������h1�͠�,0D�)CcL�� 0V��D�~�9�.!D�	�v� caA���Dr��>D��Is�΢[�A#�D�-S.N��f�<D��٧��?QD��ɂl=r�4�Al;D�X!sX<2TCA�I8�4M&D��hT���|\����,7l��%D�� �L�R0bdZ!��((�|���"O�X9b�<� �j�!�!x�p��"O�TH�̈́7]9n���@6E�ʘѷ"O.��5�����@E�\�Y�P�X1"O���S��KR�,8d�ś(@t��"O ���C�e����ƥ 3P	'"O�4�6�&q��;`ɓk���"O������, �	���"d�N�4"O0I���yP>���L�=�"�RA�'�ɀB �#�@�# 60Q�>{E��]��t�GC�������_)20	�3J*D���	:�d�����S��h9�A>D��*�"�9pT��J�b�̨+��'D��	�EF��\p0B_�?�����)D�vd� ��ݰ3��*PD���	+D�`t�Mf����!���'��=�m3D�D���Ʈ.��FD�u}��P�1D����%q�e�oٙu��Mx�:D�0ӏ�-#���ą�������;D��9�ʁ�B�x�!� ��NLP�e.;D� (�5
$D�A�U#�*0q�/.D� �pÜ��8w��&2�"���+D��;�.�UF���wO��ؙ#-D�D˃mū)���aeɥ)�<�l%D�4���x�|� �]�3�H$D��q%D
z).XA��vF�$p��"D���A�Y�Z"��SK	M�x�bf"D�h��镳S$4�R�I�8-�K��!D�|C��5�\m��ƏH[
L#�l%D��'�Bz� H��<I����(D��i0'K bւ�#� �7:�Q�F�3D�,)AAC1k�W'�9��$Y��TC�.Wi�%��!k6��� �Նi�RC�	=`Ȍ��I!7��hC�BT@C�	(�l����	ASpT�C�1�!�DC��0�j��k�b����Q'R�!���}�*m(SaV�X�pAD�2�!�ۂ1X��Q�L%}�^10v�+e�!���+h�K��֬w�f�*��aa|��|�h�Yq�%h�VMy!׉�y�˞�G�\b����p���:�y�
���X�F�@ �J��QF��yB%��~���r,�!p��q˃��0>J>��#�7�H����Y�`2V1:�*�`�<q�MS)�v�J�6-N���PY�<v�>%ҤbE 4PX�d	�oX�<��.+-)>m�j
�z+:� @bS�<�J�+o��D�Ťұ@���`#��Q�<Ibmڏ���D) څ�RPJ�<	�H0v�ꖣ�$~U��[k���?��_�O�` ��7H@�+�h�g�<����
�6��e�!-�L�Kp'o�<1��V6"�)G��X8���h�<�����}��p9U�ܑqX֨;���a�<��m� �8�.ِ%�r����Ka�<�e/U�X��Iq�⑁-��t��df�<��AF3j.��)&N 'kq��铥X]�,�IY��X	�A�,ڊ"p����6J����8��CE�Egl�x��M�Q���ȓT��vG�1��Sφ�'``��	�c�(Q��j F�&W��Q��n�h	&O�s�"�Fh� _d�ȓE������b�$ ���ȓT��{s蘄s����̮/`�u��S�? ��"��\&=B�MC��O'^��y�&"O�dB�$ۉ<@H5XT��VH����"OZ�j���36�Nɛ�k�[<@)�e(7���hO�(f&V4͢� �IW,] �"�"OZ%$��lg��)wI�7[�.T26"O��11�S��`��G3/����W"On������zh� (��^ݤ9�v"O�EYR�V4�]�4-
8�,��"O��H���2qW��R1é<��S"O�����[¸��s�O�r���3"O�m��؂C�z��Vnفu*>��#"O"1�ać�X�HI�D��Bk&E �"O*��Cg6�pČ3
g~T
�"O�<����9`W��"Q�#�&as��'E�O*�2�H"1���f�HFh��"O�1�d Ր��(U,=�m�"O��+a��fZb�{���?X!v!�q�'�ў�#I�v�x�J¦G8|��A�s!=D�t�P�R�_�ڃ��e�b%s1@5D�@�	�6�2T���96�bX���.D�(�5`�&�P!YphO]����(�	@���O��10gت=�|)H�ǢVF��	�'y����t��U��"��N����'�nz��,C�.D	�oI)E� u��'�$0��+؏T7d�3��&`��'�Иi6�����&I��jTA�'3jxU*_u�~�Q�Ȏ�qk,x�
�'�^��B`O���"I��.���O2˓��d-ڧY�,�¦B�
��`��&M�fE�'H�}2a�A,"����7��������y�ȑf�u�1)JA �!�q�A��yRFoi�<C�J�aIuY�ϝ�y�b��-�9Qd� �i�X������y"㕜�(8�-�<  ��)W �y�FݽEk����G޸;��,���\��O�����\l��C�U!p*�p8g�i�<	�U�F�x��gM�)��Y�gKEb�<aG�5l�P���N�u+W�.D�����ڱ*.��b�BP��1�+D��ЇcˡL�f�C�B *c2�jv�7D�܃7M�0�E�s��JQ��� 4D��h6��~� �#�A�8!��s�<F{���P�~H����ܳ���c�U/ ��d.�S�OZ��/�6_�T�g���g���'��8���ʃl�b�杇eX�:�';ў�`��YXn��C�ױ6��K�!5-&L�ȓN�Qr�L+EJ�(pɝ�-B8q�ȓ+ڌ��@yZ��+�
2!��܅�S����`/=:�K�*K��!���s�$��K�?\��p�ݲh�LQiV�#��<A�ʞ
�ܥ��$�50�(-�5�H�<��DF2]Y��.d��� {�'�ў�'j�:���&��0��Wi�y��7��8J��\�PUJQ9�K�{�\��o��b�@��c	"%�''ع�pP�ȓ	z*��2˒�^H^a�ԍ�[�~(̓�hO?Q��>^B�X�N�O|�e2��>D�t�!eǜV�ڰ���Βuź��D)!D��x�o\#;�`��!�����1�!D�4�'��8���RfE,ށj�n?D���g��T�B	�#-yp�8��!D�x�j��iu�h��N޷ <���<D�,�!��S�܀��A�9V�$D���G�D*t`�-�o�a�q!D�� ������`l��PS������!"O$�'*9q��yI�+L��&#�d/�S�'a;p����F��G�)DV���ȓ"���j����\X�����ɣ0T�ȓ8B�SQ���d@e�^�����Y��TӴ���]�3
^"5�"��ȓIpp$���\;{q^P1+֢�eΓ����<)���Sv`{�%�"O>:��g����V�TPġ "�,���	Z}hϓ�hO��#��8	�1 sȑ`��&��'P�B�	�g5z��,ޗH����G�L�|B�I9��J�$ߴ{8֐��˱/�JB��68�%Q��]lꍋqd ;����?	�S���ĜW�epw�3�������G�!�D�5F�,ĀL�@������&�!�D�*Kƴ�R� g(� ҐM�!�DQT�pX��Z�_&4!��?�!�dσD��p�,� ����/z�!��K�/m��#�e�F���MC�-�!�D��G&��C]�3�ّRL�v��`��I��&�Q�����W��(Ę���OV�=E��- �MR�V+|��� p� �y����5:2�9B��)H~T��!̿�yrd�-fG�=(�EI;W2F�q�����y�e@�w�T#��!.���f�ۂ�y��A4�:y�N�^�J�Pi>�yb��0x{*��٩E�V�3�mX��yB�ձQ�6XStɴ&K�4�і�y�Z�p��,1�R8O�<���Љ�yR*[7stl�۰��tx 9�rn��y�GBJNH���F=erڙ)�O��y��2d�|�Z�ٴ\�����ڝ�y��6V �i�#ά��V	��yB���,F���7E�2�ru�%�Y&�y��G5[��U�N��'H���HS�yb$�0	�� qD�ӶG��1�	��ybȄM����/ׇz+��
�.X��O6��v��^�d�G� 6];4"���C�<APF>�� в�.O�*e;3���<)������z!!"TL"`�sMIx�<�1a�E��l�Qf�h�^0#��O�<Ir�Q.r���y&�@�+9R�DD�<�PjD� �RQi���>"᪖B[h�<�P��'4�x��Ε3<��T��b�<����>�00R��A�Ԩʕ��Z�<I��?�n�����8GB��BgL�@�<I�]<i��F�g"� �S�y�<9ć%Hl�u-B��^a��Eu�<q4�^�m��@��,ƲX�mi �n�<��!��oH|�I�+W�[�]��l�<ѵ�/�v���K%L�����O�(��x�mE?E鈠��D)AK6��C@�y���j`��Ё�7D uᥫ��yb�T��}��+��1��$�6l=�y���/�Ye�� a�ıFK�y�ݼm�pmQ�Jr��h�V�X��yb��>Ci�� �H�l֪�U�(�y�]�>bOԧf��iY�HK4�yb
��h��qb���M9e!�	�yR$K�zj� 7�z��=�4
�yr�L�,��ps��2q�ء#n]��y��aj�`�F�i6z	C��y�E�b�X[P��AAL���y�M��l�D����E�qP�M*�y
� Ȅ��#Q*hԴ���F�2%�� h"O�yP�X�iPl�z��͔|��iP"O�̪dDٽw6X���:g�� 3"O���myp<Q�c
1B���"D"O�qh��C�����C� d����W�3��<E��'YP�X��R&#:��*���r>����'(�҂L�x�Re� s�V�b�'���cV%5��HQ��P8c���ʓAx��1cE8��|Zt曄g+0���8�@���bC�gMj� �'�<��ȓY� *���NM��dJ$|����;sT١+�ez�i��`B��ϓ��)��\�@�gTeVĠsu���B�Id�ʇ-÷}����2dϭ>����?��0�@{CdИ�@���xhz��$���bq�͊X�`� C��%?�lQ�'$b�'�P��v+�0�X�᫟+A� ��'d�Y��+ڃ-�����(�Ơ��'Dpd�D/Vzq�%�9Tȁ��O֢=E�$HO�(4���H.t0�q ˗�y�G�>%�LsaS!�LPc�����)�O}���6V���r��� 4Tް�"O��I��2J�:�͚/�� ៟Д'W�y�J�sbX�X�'^bm�Uc��y"dJ=]���:�Nͬ\yd�r���)�y2]&A�E�7	NR�`�	UIȇ�yb�P^\�t����tf�u!D	
���O�����8hz-{��;P��xcD�J~R�'A�\����v��Pҫ�\�z���'�|�@r"�%7u�6�V�Z�4��yr�'İ�j׬	r�����W�a�'�F-h� ��kʚ�@Ư�7OMfr�']`-�6(�iPYȔ>Z*���'� A�CʱO�$��#Ն B��	�'�h}i��^�,��,+��Y<*ѐW`�<1FN8i��LrG�W�.�(�CU�X�<�W�L�2Inʣ��-p����y"NK4I�n��7EQ;J���L���y��(�4m����j��Ũ���*�yR#�� �(=�&�̥4������y�j���e�H��
<Ap4%� �yb��qt0�Zv�P+�6t�k��y�/��HpL,*�O� �b��R���y�́:Ps��q�&�~����`
ŝ�y��LM��		�*E{����o��y¤ =S T���Ӊ'Z`�R��+�y҇ҵu�&�r��2&�6l�%���y��V"��1��R��5��	�y��->Z�A/O�z`�aEOW��y���7X�𓠌

zP��Q�G"�y�E�?�P�0�N�k���� ͌�y�㑙O������v�R=��X?�y�7�p�U�P�>l^�+��"�y"L\i�D���O��'�H�y"��(�L��&0�DQh�Bݰ�y�eס��@��8S=&��sB0�yrk"E+�}�0 �G��*�� �yb�'}�O?10'@�	����jʳ܄��3D���D�DtDd�z�+H� Gxtqe@2D���4��>�*��آK�bA  =D���%,��k�(0!���/�@\c��%D�����$h��7�Q/w��"%D���J?M�J8�H��ʃ���ybOԀ1:THC���{qE����ў"~�S�? ;ס��$'��+�A1H��f"O^	Q�yU~�kCR�{{f-I�"O�	*�(�	jS�l���]rUs"O�QXM��#�,�KvM˽i
TA�"Or���bP�tl��A�Q�6���!!�'�O^e���ںc�ʙc'L��D���Cs"O0���W#y��)Zը���Luh�'�ў"~�R��<�湪$!J�8�^u��{�<iV��82YrU��A�pZ<m���L�<�p홾ul�A�fXs�XP��"�@�<ф,��V�L<�w	Q�p3F�Y��@}�'.�y"�ۿ[��q�H��~/�	���,�y�j��w2Tpa���}~�A���y���,P�,�K�	��n�>(p��U��y�(��2Zt؃b�ÆR�� �F��yr��8b�$��g(�2Dz������y2��:d�`9 ��
�;��y��͈�y�gI<y��1r��O%E߂}C�+�"�0=A��h��b,���b�/+��:d��y���T�'�n�
7���a$��뱧F�BwN�8�'�X���E?���B�E"�2�'z`6jʛi�1�A��%	S�R
�'"��(Pe�qTp=����#SO����'��,�T�
�b��I��?�fp��'��4�
6��b�$A����'g촢эC�0�@�S�S�tAv�I��$>�'¸���n�(�PTP@��Zb8��z+8���B�UhR%Hw�B� j�l�ȓ8�Z�����+T�0]��T-UZzH��v��ewM.A����k�/=�x-��=�։���4��2m̓2��U&)2+�&v�:�{�E�W��y��V�v[��P3E����c@��	^�'��Ț�EY�G~
j+�8
�&�[
�'�l,��ɐ%LqS�%_48Cb�
�'��#�IS,�����lŤ,���y	�'����d�kt���)xX��'�T5q�e�`!��6r���*�'�X+$M?%%J��+��aH�-���'�������+���	$́�W�������'E�I$�8L��zgI<Q�~a��'V
=ڳ D�]	+#��>Z.Ġ�'oF���LJ�`��[���5��ɑ	�'i�䈣-F�<��Q0իՠ5�����'-TъЬ 7g@~(hէZ'_Ր�p�'�$�4#x�б35�.) iɌyb�)B�+�@��!�	����'��:���<�-O��=ͧ%�Y	P"�{\�PA��(�6؅�g�^�Z�X�&�pЌ�~?�D�ȓ;�l�c��7�L*��#g���ȓR��Se)�&�5K��p�y��͂<��b0zQ�7*7s2&P��v���3��8B2�iA��bþՆȓV =�c�d)|(��g^i$�F|����b6�Q-n��HJ˽3�4C�I�L��M�QeR�BR@���8R8E�	ڟ��'��Z�b>�	�*�
\���ЉT*P���BS�B�ɘ~w����_�z����Cd�]��B�I�)����AB�r,��	qNG.�B�I�Jߴ�r�e��\�}��i��)�j��<��<����c�p�s	��NI�Q��]�'�i>�Q�	�Sby����4��:#e-D�<�fiC�cW T�b��v0H�6�,D�iT�"�f���ږo���!)D�� ��s��)7$�1q,�9�fhE"O�K4�¡!-�T#�
Z�4ꊑ�0"Oxy#���#Cb���4I&u�6�'|�O�J��Zr�ȴm@�9���0>O��=E��I�omD1��Ψ^Ͳ�FM�y�/�x�|I[�h�f����0���'��]���'��O�Q�&R1*�(��p�T"OPi���S)m��V���p8'"O\ܰ�i�3�5�E �@ז1* "O�aж��y���q�/�$�ZE[A�'��O0�sd*:7��jsIԩK^�͚�'#�'2��[��v����e�% |μ;�'�ŋg��!մ�SEE���P�
�'uEJ��l&|\zѫ�*`iVp�O����>qƈ���+�*�#HرuH!�$T+%�����˸O�`�I�GO(0!�FDú���Y�,]C� (!��',��y[�R�L�K` P�`�a~"P�H�m�%\�J�����&k$P�v1O�=���Q.^�9��,��i��E�?���?���?�*Ol˓���Ԧv!pHr�F�@��k0�ߊy4�d2�O�q�	�,x`(N���#C"O������ m�	��?�2��"O"A�FD-rú���^k x��"Ox��"�:2U�d�gŪ?s.yc�'���|r���]H�� Da�2;�^��yB-LJ�pE��,B�U��R��Ӏ�y'�2z �DQUI7J�*���%?ܡ�d�L̹�B
�1D�f�U១]�!�$J�f����F�<g�M����!S!�7`i0�4ƭ�X��!S�Raz��'��S��H��F$<8X!��#ccr���f��E{�O��OP��F�CJ��![ac�N'n1C�"O��bmM�J����睜J�Y��c�<A���?��Ş��9O��P�I�(�b�%�sR���"O�`6h�!{"Z)��:�A�?�!�䝀h�yp�$ыF�vT���"�!�d�-nz�d{�%��(a@ �"Ea~��'UD�c��ls��2w���S�f��O����Q2"@��"�.'�.����W�D 1OB�=�|ztYq~횱��3ST�����<��F�	��(Lr���&�PL4��� +�⌁,/i�=q����}�J`��~k��rD�0X��h�Rn��i�ޱ�ȓK��	NZ1��d���`$�����?Aeӫ@�n����!8�4E����l�<��.K �2y�C�]�48�=#0�e�<�`����l�釬:�M�' ʞ�?���?���?��2_�x�t�J!)F2���)\�Tp�I)D�����Ԯw���R�m�}�^ �,(D�h`T�q���d��	b�E#�&D����֮i�`����YQ���%��C���)�O8U�#O0_��BE�E`� p���<A��4�����J9Am⨐5+�,\BP��'�t�R��!���huC�Eژ�C�'���''�X`�F,e¥(V�0�Y��'��E��,Y�m� }��y�"2�'���X���H~�aC ���E���
�'"DXIe�ϫnEb�аG�)9�R`!�'3�ͩ�Cf @drs&;[r�p��'�2ݢk[����
���L,1��'O�eB7��!J�Ō�T����"O������i00H0�̕	`(��"O@�y��8I|��4	���8�"O� ڠ�M� (���qHܮCl����"O�t�U@��|��@�h=IMH��""Oz ��kV�3Ǌ�1��S-O42U�D"O<l��	�x�93�i���"O~���P�1c��9G޻x��Z�"O<�
���290^�QDE��-Bܡ�r��O����� gkP�aV����t٨�I�+!�$+�p�Մڿ5~�L#��ˏl�!���n�����L��T�E����!�d�|i�	yto��Y����S��j�1O`�=�|�2nJ�2���$�!F�t��Q��f�<�%� �n$�� d�c�Zc�<yw�G��S��xn��#4�I~"�'w�{Rko�h��wM4p�Ä�yb��1�>�Q�s�8�ާ�y�"�Q��E�"��S� ��q����0=9��'N F�D���g�Q�u�1O���y��)�'G�X�5.�.<��4�`B^	��Dx��)"I> 7�y���6��H��NJ�<yp�!W��dbץ�"�2�q΋l�<I��������� C�BL	����<�Ë�#�~�kV��8IoF=A�I~�<�U+�> �Dt*eN�-�<�s(U�<	�c#��-J$��'sd�!��kF�<��攰T� �$��_��d��%x̓�hO1�H�㰉��_�Љ���B���أ�'W��6ӈ�B��^��Z�Hd�_,{�<���>���(14���� $j7����`�<9MA�z��4Y ΃�E���S� �B�<� Q���t ��Or��3n��<� � ���	�FNL�& ^}�<a�jK3'�1������>�z��Cs~��'\�O>��sv��x��T�H9ȥ����>���Ox��TM��|ߊ%� "DN<ZU�!D�z��
�b��rҭՠd_Tl3D�P:����	i��"���K��&D��B%�S�Xp/ˤd���y&,1D��@��ڧ�.�+�ϻ8l��2�*0D��b�@ǡ=���Ή �����9?�H>)��	ƊG�9��(^<ƈ�WF_,���.�O��Q�֟3�%"�!Y�r^nz�"ON�RR�(R2$��a�1`M�t��"O�)�F�ϰ�����)v3vy2�"OD�h�lE:�ԉ(�N__u�P!R"O80���
*�L��Ȓ6kg�%s�"O������w�nq�7�� ,DA84�I��LE�D ����1K��iE^a�@�A �y�@ظrk�4bC�Z*t���­�y�G'bn�p"��Aw��̏.�yR���,Ь���.5rye��3�y���/1�r)�� e���4&O�yb�«W�����W����ӏQ��y� ��j�����K=<�0��Ymz�O����<1L~λ<�d�E
V��h�{�)Gs�hUI>�.O?�)C������ɵE��d���;23�C�	D��	��I��;#"�I��эL�HC�I4�<�R%]�m�$$������B�	�N|�xW��,6�����[T�B�ɀ7��q��g/MEҭ�4e�	��B��-�|��A?Fqv�cA�16��4���4�'���ɒ�v�;҉Q$[E"����
�{U�C�9_"����!��I��C�k�hB�	�]�z��jͳhi��/B�	$~��Z�iJC � R�;k�C�)� `i��k(VK���W������f"O�}�����,���w��"O�H�VbV�'�8ܩ��S1jk�0�"O 홷�S�fx��q3�J0MZ\Б�"ON���m�V%�qH4KҳfR��"O�q�-!U�$�"�HȪw��	�"O�����w��Ϫ���
"O��2g�S�rR���S ��!�r"Or�	����TX���w$_��f�{B��O`��6��<E�C��& �-C0!H�E[$���ybɚ*^pњt�L��%X�C
��y"��}-4�8�m���{��5�y"�E	 E¤�J� e��/��y��	�����hő�bW�y�(Ҡa�8�*��ڷ
ʊ��#���y�	O����#�N4G��#��?����<�(O��O���L���r���x(�Ï�!!�C��ϟ���$ď/d��{�-�FQƼ��&ah<9珒��b�a3���+ �\��oEK�<q�Β}qH��Y;/d�7�PE�<��D;j�; �"�Ġ�~�<�+ҿI�>ȨA7%>�u�Q��|�<i#㊊8�8j��\+g���ST
R̓��$'�'u���v�1�p`2t"Z�Nȴ����ʟH�ɡ^� й�@��r|E����5]5���s�,���c�82  <{':��H��Bw���<TFlC�P4v��l�ȓ}L��C��c�r �W5�ZE�ȓ)0x@�c��	�(��I�
x��ȓE�l�h'��P`�6��]"���ȓF��4K�A�!.�i���J./c.}�ȓV&��YBhP�(mj��C?p�p��H�iZ��C�J��T��YHȆȓ'M��uM�|,8I3e�ܧ.����,����GG�~�x���-��%�ȓmg�("e�!������~��U�ȓd�v��I��{�<�P��]����-l$h�ËANyE�Qb�Q���~Mi6OӠTT~��1ȃT�$,��L�ά��JJ+B4���2��|�ȓ7�dIa%� 1l���UHMND�ȓ���⃒:A��� �-S��ȓo`.]5�Ģ_����6��Q'D��SB��ւ�h�ۀm���h�����]QbJU).�+�]<zp��ȓ�J�����(u����#+ p����ȓe�($r���ty���V:�f�ȓG*dhQ,\iS��b�V�`2,��ȓ��`��&Fo�AB�_8M����ȓ�P�v@��wa0MS ܰS{�A��\�x��G�.���SS0/qU��#�&����'
Q��� � , �D\�ȓ��dsԏ�5*(b�
o�X��ȓz*���ҮA6M�6@�`�rS�І�sd���c�)d(�a�ׅ!w����n�c�.�9!�y���=:7�ȓ~���W�5��%�ǭݐ&`���)҄�Y�>�򈺄��W�u�ȓ+���K�"�����H��{gD��ȓM��q��~�(] �,��u�p4��U���@ ,�����W�U~ ���Y0TM�C��/{T�&��&��ȓM�-�WH�p�Ő!�b��\�ȓ<�@|W#�-���D��Q�n��S�? ������7�HHBH��P7����"O.E��ښt4D���m�l��D"O���l@����p��=|�9p"O��{Ë1>M� �D8S>^�C�"O>1�"�NQ�z�+��1\qHB"OT���nAGf�m�5@�&7�)��"O~��6%�ac���Ο7+��@+�"O�e�,N�jH������R,��9 "O�a�A�_��F䚧d��/,	c�"OJ|K�/��7J(Q���bp�hS"O� �a̍�5��$�k3�T��4D�1b�X#eOH	bM�>A���D�&D���� �N8���'�iR��J0D��!��b�.(��o�;)�D�
!D�(�g�	k��}��b���j>D�"�C� m�DX(q!�(�t��d;D��س�V�o"�(p*�'i���K%D� �e�P�f�8�;�+Λy%y3�1D��S��J4K�Д@PC��<"�!0D�x�����iꢋ�$"�lӵ%;D�$�@h^���AƦ�\���e&D��I5�ݨOE��*�̜rbz�8R�$D��0��nK�5;r�\�J�|\��-D����k�$^�<�K@�_MJ�9��+D�ę¯,a����t�7v���u(D��r���9]t8�'��(�ܠ�)1D�8�$��>����A���0o����/D���V�� ��L��G��o��-���9D��[g�� 3cԴ�-�	c,ČR�6D��I�(�"U�����Xh�(�.6D��d�:����@!@.��C#3D��͌>a�>�cfNQA���1D��ed��q)��s�Yv`��y�<D�����R`-�aX�*~�٧E,D���@JD+U��UҪA�Uba�2�*D��H4jY	�M(���5U��CpI#D�,0e`�6H�pc�1D�`,D�LP�E �R&'���b�4'Ҫ%X!����ugN,"�\�n戴sFΥD!��ٯ�t�B�-��i؊�#�c��d*!�D�4�@�0e���u)!��H!��֧�h�*�`�B�;ϕX
!�dΉg���)�OK
f��ń�)!�V�%�l�?JZ�����!�$ 9T���ҤCLa�$)���!�7IFr%��d`Tb�H��^$�!�$O�w��LqS� ���鱠�,c!�D� Q����uMB��������z!򤙧l�FB��,�b��tKW)4!���1�g�0a}��#���`'!�Ğ/=	�P�Ɋ-^��(��&!���*6 :�B�`��E��}!�d��b.�Dy��)>��7��-�!�$Ρ�"A)��٘H�r�)w&�D�!�D��z'
с�ɦX����O�!�d��l��Ơ QdĚS�Rf!� *<������"92����Z4!�d��zϼtc��/p��8��9r*!�ЭWZ4�ʡZ�s�2h)��^�!�D߀6FJ�jэӍ �a�I�6?�!�?nx�c���E�� �%��FW!��\�� ���E�/�N S���!�ă�9R%ۑ`2#�0!���R%g�!���4S�Hm;���h����SJH#\�!�� 8Y �\�!�X�k�Ƨ��\�#"O� �Ū��z��Pr���T���"O^=�Uᝓ|b�	��O��<��e"Oٙ�OW�"��T����1qq���"Oj�"3%O86MR�S�&q�2"O�A��%E9@��QNEO���p"O|�Ҷ� fM:1�1��d6��8$"O��0�d���j\QtlC���"O���PH*` ���$����vX;1"O*�;R.[_��	[�OͳE"OL�cק#t����X&N9��s"OFLI��ɨ;�T͊b�������"O���%NɼCITq����&w�N�s"O�P���
�����%Ɇ����"O~h�1-�5l�1���Nt	&l�\�<A"��,���1Ɏ(;=>�8���r�<A��ȪX��A{g�ܣzff����Fy�<���_3	x	�V�¹7'���Ew�<)�'�4��a2J:I�("��z�<��I�,w�D�q�9G���2���Q�<��O�0LLP�
���-�)�A��K�<9T+�,�*���/g����.E�<�G��)'�=!0D"�� ר�C�<� n�tH�a��e�\:�H�{�<����$&#�HX�~��H���t�<13e�9_@P9�D^�q_���	h�<Qb�;L�Ј�W��>~�`�#�Nn�<a��G�mS��v��70���S� �l�<é��
:T3 g7
�䫓�O�<����n�H�,�-������M�<I5JRMv6��]X�8lA�SF�<ɔo��,N�ʂ	ȏ��X� B^Y�<	�蜼]�"���-��P�X�Yv�KX�<��R5D���� �!�j0�5A�S�<AV��0���Y m��G�­#���u�<qiߙ4�X�$!�^|��`
]�<��C'I;���� ١>�BW��V�<IS���W�x: G�G�5� F�T�<��aN 1^d� Gב{o$q���F�<�&&�&b�D���
�l��"���x�<q�.޽粕��
Ϯt���)CƔr�<Pg�<;���"Y%ft�A�Mo�<�&O;(vn$��hءU�D\�֥i�<1卌7]c�!�TN��c->�j2`Yj�<ɦA�zd���T�x�fDjC�K�<��A�53�b"h�5gP��Wo�<�D�Ż:e`|8�S'q�0�`��B�<!��;'�E�%�<��8w�\B�<��a�O���B�_�D��R�	�<�0$�kGʅhT	�"�䄹�O�A�<���6Y��dkF@��tF��0f~�<A�JF�����I�e��z�/�r�<���K
c�хG��"�@chf�<A��ք! �q0�K~&�م�I^�<��lJLܾ)h�FB (�2�x�m�]�<���*'�Z1��a�83,���R�<ӃH%4�$�BK�U?�䳦mPK�<�V'M-f��<Qcl�-@r����H�<�6�F1\BQٖl�<�.���K�N�<��X6��i���ܑc�R���Bf�<qA��N����L�Tp��
Fl�<�P�����y6�
/�Yۃ#	j�<�B�ed���4cٽNU��`�d�<�v.��M�����7{L�1��%�e�<� ����`w�H�s�8m��P"OF��ª"*��Zgl���.h8�"ON�z���c�T� EH�{�T��"Oj!0H�"UHb�2��Ч�<`B�"O� ���C���t�E74u��"Or$�����`p���^�̶�
�"O���DF�]��딷/Մ(B"O<���D98$`���>�"�R�"O���hM�E���:�(_�'�(�S"Oi��ʁ<n}zʉ���1"O�])�X�o�25زG��W��Ɋ�"O���GN��.&z]a�@2`���� "O5��f��yˑ��+Z��yeLq�<��K7 �pc�Ӑ�yR	�E�J�H�ȷpY��:a����y�ǞDx�a��m���P�yB�� E���e�o�ZQ��)���y鑋tD�h����kKΡ+w�4�y��L'D��03��c܀E@V�ɸ�y��u-���%VX����e"�%�yb�M�7�l�&�M{����̎�y�C/|�l�A '�Fzvȱ��	�y�
Љi��%ヲ(	n9�L�!�yr��&)�y �E�������y� ȴA�hO�8m���'�7�y"�э-��|���ң7�y��痡�y�i�l����w���,ޯ�y��ۙ�,spXD-��JC��yBjG�& H��5OޚD�nxGU	�y��2R�(�1@M=��T��/�y�)�$A�5�a���X�稏�y��#=�&t����<�7��yRf�&Q����	؀Buf ��yR�X2���W��-9�eõjW�y� ރ4��G��3��=q6h�;�y��:����j͕{��pF� �yZe^�}��*^�n��1�рڔN<B�wH�)�.!`m��A��1��B䉊D~�� �ܘIl����NS)lB�	
*%��*�)�_�����T�"S�B���Aq#JKԀ)�����ԖB�I�,�����R�R��G�ԉJB�ɝ��=��Ǟ}��d��B� nU�`&��z����gLV��C�8&D�NT�X@>L;�ᔝZ��C�	�}�����,ULk�GX�E��C�		x-h�����%P"��B�C�P-�����S�d���� �2e�C�I�z� Z�r��e�ߐo�@B䉂J��
��$'
H���h^4yW�C�I=/8��W��'�@p]^'�C�ɩ,Tx��椔<<����eF+S��C��#&���0��څt|���M�?{}lC�ɦiB<�I[�N# �Br�Ѥx�C�I�n�&���B����y�g�=P0FB�I�D���1��=�ݰ�!�,x<B䉴S��qV@Θd�h����&$PC�	: �Ը���V��^!��M*EyDC�Il� \3W� 0i�DaIC0�C�ɩ��|��L^te�CT���>�B�ɏ'��80�U�(C�.o�C�	�>!�OI��Z�8�$	oPB�9�0z!�(gA  x��!�$B�2Jll�P�:Q�^xA0h��ViB�)� �����(m=��[ /@<��r"O"�9�%�Hkht�!��(9�T3""O�\�'ܕPE�9�ˤ	9Jq��"O���s��%yjx�`�H8�!"OZ iGGS ޜ W�]-F��2A"O^4DQ�\(:��9}0&�A"O�Mi�)G.I}�M����')čZ�"O� )4��Dr�2fe.N��I��"Ob=I�)�1Zx���c�l��|�3"O !m�֓^���1��%o�20�"O�D�c@D�z��(��g� ^��K�"OBe��3P>��T�``p�B"O����Ą�R�= �)��b]�iYb"O��s��]�"��0�A�`���w"O�<Z�H\�=\��0' 8��L3�"On ��F��X�R��"G��(�;�"O�đa��C�*5 R�)��@�"O \2a�˅a����74����"OV� '���QO���5�4v��""O���4#,"ܺ��R�?o�DCG"O��W�י1��R1�4P�"v"Om���9��`��FQV�4Ѹ�"O`�UF��k����R�^)	�"OTIRF�I�>rv4[0)Ml�c�"O���GetN�{�`�%�jd�"Oh���F�#�9�A�Ҳ.�����"O�%QdKE/_�
��.�7>�6l"�"Ox��t�]�L���4�Ȧ��dc"O!���v�<Y6�O� �ve��"O ��犹r֎�3�`ϱsX�4�b"O�	�W ��9����NB>Q���qV"Ox��ѯ @2wv��9�A"OT<s1��@g�e8�o�(�LQ��"O�(a��?p`�aUɐ��a�""O��L?hY �[��&k���"O8� a-8OB(���A�x*w"O��CA6�t�[dJӗy�̩V"OP@�(�~3�����B���2"O0 �4K��`&Z)�"tH X�A"On�AP��@	���O��Z�"Oڜ�.���B(��6B�T:�"OF�Bj�WO\}Xp�
3P��Mh3"O8��ĀrsRI�u����8��"O�k�%�|����$T3��ä"O@Q��K$���bF���p�"O꬚c)L�[�e �_E��Tc�"OHh�-�C�r����	%]����"OT	 ��<s<б��
 �����"O0���V�V Huo�\@TT�"O��)����p:��t��~7�}��"O�4���	�� ��[8����"ODı�'ٝ"F�l���	�!7H"D�D�҉Ra�􊶅��#|���e#D�B���x&vER����C��qhׂ D���ׯ��#����K�B��(h�C�	D���b�V�@��)V��A��C�Ikd̩Z�����m[d-UT8�C�I�P�zU	�:A5�Y���G�x�C�26z�k�e�����Ź&(�B��sl��F)1�A�G�VB�2�Q:�H[�L��gB��S$B�	7Bg6<ِBTKe��R�HB�3%�R#H:Bp۲�ڞB��.	Zh�1*qv��i��9uB�)� !�E�	$G��@���R)m�l�"O�4B�h`u�	��&�01��#�"O�kQ��焍*!H�p��8�"O>a�w��SŁ�L<(�r"O�9!R�X:|��(Ձ	��#�"Oޝa�F�.Kܜ�B�F��e�l 9�"O����b�  K���jTo�|A"O2�)��ʙ`�&�i�[�`0�"O¨� l�v!	&*R*8�8x�"O��P���-�(�W��`.С�'"O� ���;�9�F�I,(!�"O:T˶�V	�n���ە.��"O���*��mY$��Cڌ~���v"O���CM�%s��8��ũQ�"�"O�A��Ϗ�AU���̞<jl�Z4"O���AgG	g{��ec��b�rػ�"Oڄ3��T��$��N�`"OH��1&�?Y�(�����6��[�"Orp����~��ir�`�E|jٲ�"O�Lxp�U���q�s G$l����"OR`�D���t
��!��`R�DBa"O.q��:p9����B�_-*��"O�} KҤM^p�R �<�y�"O��I���|Aڗ�g� �'˻�y�X�S�ɹ��ƣp\0��$���y����A��Q{q��d'~ܸ6�́�ybo�X���	X��`�&[��yb��&�,�q�D���	�C��yd��T�"h���и  �<�1KG�yr��23�6�!TFړ�r�p��=�yr�
,b�l"�,M2^�A���W��ybm�0I��M�椋r�摈`�
.�y�lE�p�x�AŁҪ|���#�yb��&o��p7R	�� Cc��ybF�$Lj��"%����B΅��y
P8n�� 'ɒY�#�\��yDʬS*��s� �/�	�����yr�4B̊��Gf�{2���B$�y�"��\b� +ʈA1�e�"L�y�K d���3F�A�6I�_/�y2�U< bT���ߪ1�yP�?�y2 ��-���P^�<��5��d֠�y���D���˦#�9~��/1}��ȓ{��1�O��P�Dm�B��+0�h�ȓ7�!K�$V$z(y�ר�4��ȓ0��̙ͺ"\iA���g���ȓ6��]� �LGs��8�/��'�t����XP�%@�~����EW"d$��1���cGnQ�Y@g!&��Ȅȓt��H�j3�=�KR���e��.[���2i�	k\�GA�+(vX��>���qň/v��8s��Z��P�����,Wn��jZ�{R�Ct����8&�0�$YF�PMG̍U����_�X����+qd$p��`�����zl��f�B6j�,��&	r:n!��~��xs���E��U[7��y�]�ȓ=��E
v��WD+�e�����ȓ,�>�X�ƍ+oA2aPp*�Dy��R~ ��B�QR���A�A�M���ȓ7�I
��Yt�� ��׽����ȓ;�F�������Ql��xg@�ȓ>Y���$Tl�T�I ��U�ȓY+bpz��	M �[G菝9��<��S�? ,j�e�;��PQ���2u��uRQ"O�u�R
�<C.!��@0Q�bp)"O�E����]W��0LO��~�q"O�,�+�xD~m� BA����"s"O\�7m]G
i�#jL }���A"O���+�5Pʉ(�)����ti�"O�P����'�]��ٝO����"O�S�L���AT�O���"O�}@#����{�&;3�$��"O���/�<o�=�S"[�x#�"O
p��ߣ&��1��T����v"O��3�B�̀���q�u��"O�AF!
H�ր��6m>�q"O��
��iٺXBN;%V<��"O��r��E1A?�`p�MV�Y@"OFd3Lۦ;tf���L@Q<h�4"O���$d�����ta:ͺa81"Ox0��k�[h��)���b̕�a"O�	Lժ|�`-����n�TA "O��q'mA6S�4�RS
� +X�9�"O����C�b�C��,X
��"O�׊/*��rצ�.@D����"O����B%-�E���%R41"O�(dDˉBt��b&�N�E�"O�(����F���;դ.�`� �"O�u�4�ơp*�li���'*���"O$kqd��1�Q��"��V|�5Kp"OιS���.)�,�Sf̨r"O��� ��q��TҀ\�+\ƴ�"Oh(3q̘27~!�V���8s��6"O�cC�£����T�i,D�U"O���2O���h%���)�Ne�b"O��0�
�eyT��B�vp�("O�y����i��dH�b	�SSQ�S"O8�ʒ�V�o�
b�!�r1�%{�"O@]��"�Y��2%O��/��!Q$"O"���B�$݋��-���s�"Ov�QC�^-
�����(߼C�d��f"O4����L�Je�8���T37z�k�"O��b��I�x��� ၧz��5�b"O�Yy6	ͩZm"U��)�,*�Vcv"O�M)�N5NTD����w��AC�"O�Uء��j�h��e���q��"O���3�U#`Kt�'bZ�4@Y�a"O�]�mȷ~�F�E��zp\aS"O<-����!�$����R�4x5�A"OT��[���	{�lY�n}�"Oju1��B$����1,Λ��d۴"O��M�u��q!����e\1�"Or`�`�ݼ60QeA]�"H:p"�"O<Q0%��\�,���/�y�T]�"OnEh��T=D�S��8��$��"O�P`�ͯ�~�d��=�`&"OZY�U��6oB�8�Aś"�EQu"O��r��*�� ��ɟ$0`�x"O�њ%�ܝQf���(!+'Ęd"O�I��J��9;'@�$VI�"O,��W,��^�U�`@?@"��"O���2��|pȭ+`ԉ��́"ON<i���8c��3��
v
xBc"Oh1�.� ���k�KLwrb)@����D{��	V�]@l��2K�Z"5���4{����G{����q�I��	��U��]�t��B"O���e��n└��C;mV�,;�"O� AࢌZ+32����^%a�p�"O��ۓ���W&h���fITЄ�q"O@���.Q�bͮR����1���"O�ip��%b%j ;ѫC�Bꀘ��"O6�2�ǐ83��hyc-P�>Bt,��"O&\R�j+����r�D�<9$���"OB�9��F!WI�(��6(�r��"O���a���:&n�30ЮQ:�"Oz} �K[���!@�MLM��`A"O���C��T��F�. 
�"O�t���<
����,I���"OFLz�i�#M�� ��aK8���q"OhtC�D�	�d����I��;�"O�|0��#��\r��پ5�C"Ol��b�߆@�(5s��Ap�z�"O&�����)͎��(��djd�"�"O�{R�C�T�����ǉ� z����"O
�y��FM�sԯ��E�ƑH�"OȽ+�)R/k�Ak���L,�cF"O6�(s'�:-��I�I�.�|� "O��r��[�����ΏM�v@$"OzS珋=��xj��k�d%"O���N<��xi��ў�\ �"O������<5D�UiœN��px�"O�0��" 
pr��R
"�LD�&"O889��GmY��ãH_�$I>�K�"OV9
�O%i��@��m5^�h�"O���Ԍ0jfQ���|�YC"O��oA�duf�R׃�}�iig"OR����j��I�
=UxV�9�"O֠�1!�g�8U�,�5²t�"Of����="<�%��e�����"OP,�`N
�
(����ß������"O����PȀ!��L�f�h�#2"OT�C��`vb=p��À[�M)B"OTY���(-��2g'�nZ�!�"O����A�@v��1�M!�x�0"O�h;7�>jT��g
:�:}���'�1O�a��i¨V.���H��}z�x"O���N4h�]��<2e.��""Oh8P�U/T&����m.nر�"OH�J$Fܤ�����}'�%�d"O�����\�Q��H��2���"O��7�?�� �Q5]AJ��U"O,x����(h˵�	�)#�0; "O6 1��U-"d���A�0zfBY3�"O��s#L��qV�� �
�m�v5�"O2�KT�N�r����䁉�" Vرb"O��y�(2���s砃8�<�Ѱ"OD8f!�$>�hp���4|���"OԕP�NV/��RaNN#cwܵ�&"O��0��6/|�s��jqn�*�"Oʐ���&l���Ql�gXI{�"O�5Qp�_;
�*�L�fZ�1+S"O6\zan<��q��&zTR-Z�"O���Si�l�f���B�M)��)v"O�� ��K�e�X�ΰ{�.�:�"O�P+ �3Z���@�Ⱦ��%G"O�%d@�pp����)�"�Ct�'�1O��S�ck0U+�$ŵ3?جh�"O\t�U�G��0D2���=.��G"O��
�%ֹfu�D��8l��z2"O��ZХ\�9+z ��91�ԓ�"O��ʇ������^�i�b��0"O� `�[g�I/������^U�r"OV阃�Y�j��U��*������"O$��MY*;ʡ��'F	�0;E"OxIu��z\�Ӫo��JA"O�Њ'*�L���dhc�u��"O��9�umFɻ��^��n�X�"O���E�v�n�ӳg�A�����"O����b�J����-q����"O�@��k�$���a�Z� n�"O��:��]����
�I޺] a(u"Op�jӨ�#>V��^���'�\�!�Me�	�$E��]��j"d
<j!�d�*'��!��>{���S�L�!���,�6]��^"uT�Q�R�ɐI!�$�[� ����+ Z�`{7B�-�!�f�i�+Ϸno�ls�A�V�!�D�b�y�T� b�qR��þ4�!�$�f�f�cU�C�W��S�*_�x�!�d��+�F��NR�?�j,�ǟ�s�!�$ca��C�}8��c��`�Y{�"Of��m�@l��[��Y��~��1"O�ٱ�X%��t��+��� �"ODQ����#e?^+��s!�G_��!�Y�?)B)BF��N6����!c�!��$1�D4E��$A��yv�V��!�Ď}L&����:$,�9�`FDj!��U?1 �ة��ռ/�]hcE�(`!��,���c��s^��%J\�_�!�D݊�f=0r�	�?<�lЯZ7!F!���IZ��*u�R$!��!c �:�!�²$���!�BC�~ؔq��V�!�Ď�h�J	E�jg�P�p��	v!�T>)�`H5��`�ո�-ߩ^!��E��r�G�'eQ�9��n�#7!�D\$y��apgV?CW$��@�*K�!�E���lI�`r2}�uN��!�V������4mWh ���'5s!�$��tU�C懤V^��3g�?nk!��]����1��<,ON9JR�@�VZ!�d\)a�������`I� �9R!�$H,fǸMs�[
z�0#�ND�RC!�DHA�hq��S��"�#[�(!�A�t<��4hRW l��%��B	!��U-�"� s�C�Y�P�S��� s�!�Ŏ3�\1�0C\�9�l�
A�X�!�!�$Ь'*���/ݴ;ܠze���a�!�%1�b����T�5��������!�BX ���o��q� AXN!���]
$�t������JN�P!�d^ =5\��%`�`0�� ��1z�!��Ėa��E�-� ���!h#}�!���v%A��O�5e��y���S�!�|�l��&ݏ?n���uY�'�!��/ N��:vJ��{_��ؕ
M$Jf!�d��j��9+�_�JK.YR��fD!�$ɨ7��}�4d�(Y��S��+L<!��_�1sգ��Uz�;��
�(!��%[.����Ck@�� G�!!�D�V^��p6kԾgJ��Hf".!��ٞ]��=@clެM�Z�!C���!�d����]��-�>��"<��z2��=��� S�:Z�l���ηM9��4$�;Ƹt�P�YS�<�N=(���K@�,UK���P�<!�&���:Ggέ'w&����K�<� �ỤgF�F�^dX+ʻy��D� "O�]�@�U& IBT�ɉ�l�;F"Oĸsw�
�o	Xe"����� ��"O(�2�O��Od�[�"�R�.�Q"O^�ZvO]t��X��<E�y�"OV!�"@��4�d����ˮJ( ��"O:��T#	��p��%�JVpv	�"Oq��a^S�$����s��*�"Ou�wL�;���T�T5o�hS�"O�;���#M0������x�"O�1��C�	yj�[S"޹h�(��"O�l{7�E%%W�}��!�3{Ҁ�"OX���Ȟnzxc��֤QW�<`!"O`�,-(@.���Sgb�3�y�$U�w9"l���8K�����y�n֧S�q`VHэ8В�y#���yN�MqdEӵ&�5N�8ꂤ�1�y��M-iT�w��+U�4�h��y�M�6�X�C�	,|Ra��ߪ�y� Y9@^��!�ݞ$Q^��c��y�S�OePx)��J�T9���D�y�'�O`V���/� �������y2ǆ�9�b � �T�.�����	�y"懳U(�,�J&n~6p�w���y7z D�7ꗥY�xt�0��yℒ�F�xȷ.T�RM���_��yҭK^�v]AQ�W/J��0
��� �y",W��A7	�5r�X�Ƭ��y�m:.R�97'�kt�����ybn�T�n�#�'_�V;,��%k�0�y2�N_��T)˗Iu�4��ʎ:�yRT�)��2�ܓ@x���χ��yb�؃��T��" ��X��B���y".�3YP�@�'�C�7���+cч�y���h0�D�Td�!)7$ [�J��y&D�Z����V�UC6����y��  ���O�$���"-�*�y��X�e�Ձ�'�pi�ѮX��y�)�*	Z&�S��f�t�a��y2���J���6� P�|Q0�^��ODqbp���(�L4@3���y7�hz�*��0�Nm��"OV�8tᕭ-�vV�CSdM�����Ъ�d8\�s�>E�ܴz��4�HE�X��.3QH܆ȓS~�D#O5bT�4��ށ��d��y���BQ����˓$���`J��+��ёogP4��Ɏ}��l�B�	�h�R2�ЭDz��Qaʋ
 ����7L�*$¡���'��$�bX �(�.�B����(�n���S� �N� �)J�$�2X[#��d��+Fe����VZq1�n܆v� q��|�ڬp���g��E8�ѦK�z<��J��~��Y2m�đdGεB�P�T�yҫ�%s�H(���C��AA��?9w+��@�Z�$OB�Ը�W#�	;@�_^#n�(��.q��%���S���B'��Q(�)�&O
�*`y�n]�YB|!n�i��h��3��$+�K�!=�E����e�?Q��B�lLu1�"G}\������F���o��|E���^��y�*K�7��yp���G�hm{��-��h9�ބq缵1d.��?����O�\hg�*<��8����ڝ�p"Or�P!��?~b��*[~�н�7�'��a��T����gϝ
~2ax$W�țC��&M�ܝ1V.���=��M��`� Y��	�T��y�"	�[�T���[*[I&	����xߡ'�h�Zu�;9v<�d���OȘ��a�GGV���j���O���ҵB�Kv�|���TK H� �'�T�H�eU�%ۀh�׬Mˠ]b��&XZ�a��ȗ}����S��yb�_�W��q�ۯqa.H�	��y
� �Dx���=#�|��O';3
l��O2�1E��%y0Ɂq@+,O�}ے��LA�YAGH܊}!�a��'�F�S�I?nY�	%$A�aw�9r��*7e*��P�Zh<A �_.����@êVA��&�u�'!
���ET�O7պ�ǘg.� #�M�3��Q��'a�;�@V-	]�0�2�##)py��'��)�oC�_�$��AJ��4/N0�'��pӄ�]�Z�rF��>� ��'���bK�4C���q�MZ�1����'A�x �G�V�FE*��e� ���'�j=��n�#9Av��w#�*]��$�
�'���g��o���u�T�<�0��	�'J�hI���'b{��yE�O�>���	�'Sn� �F�5i�4J�c�(2��Q9�',�P�b�!��&�!����'��)�Pτr�d�@�n��+��'܈�v�6p�i�c�7�@9��'<�� �_�& ��N'�Q��'!L9i�#�\�t���aT`�-��'��P�F^.D Z���H�cz���'G�H����in4yQ�G�X�"��
�'� Pei]9m�Y���ޞ+�64�	�'���━՞4�pC�q5("	�'y�(ZS�هe؄	��e��X��'��� 'h��:<�-pG�D�Y�>��'�n��p�يVa��xp�GU���
�'��T�UNR>MF����??[z�!
�'�xl0&
R�r���1I��d����'�x8�[�e=r����(����'�`���f�=�fl�Vi��}q\��'���ia��r��$�%�A���q�'�vȣ�$O�t�%�T	 ȅ�'^����-�7�UC�
�8V��H��'�<�!�=?9�\PӬ�V���'}P��%f�`|:�OэG^4��'`�;?=eJ����S�$td��
�'��H� &�6�$i'��Hn�
�'Ineq�a�p�I6��?\M��r
�'Lѡ�K��aZ��R�I�0�	�'����Z�4'���$G�(��t2�'^�\�!�	!�%
D�#,� E��'�p������p�'�j�J���'�>y��@�:i$�iH�ˎ�`�$i�'�<����L�_���Z��=*E4T�'����!�3_rЁ �&����'���Ja�	�0����צ_��'�2 �CLl����_�C�HK�'�&����9u��Q�'��E,�;8�d�(#<q0�x�'v� 0P���E�l�3Ś�zm*���'$������|�vl�K���'�4�
�_y��8KƁ�6s��	�'zx1H��6�����CH
��'�HEӑ.���6� �F�$-1�'�J����KH��'�H�<����
�'-�yʒ��0R̚)�R�D�|)	�'Uz�Hp��b���!��D�Ԍ��'J؅��d��X�L5���<�X���'�� ���{Ӯ�	IV�{OP@�
�'�@�*��++|�hpd�/i&L�	�'zH�;ׁ���2�*[�k����	�'��1�7H��4��;Fǉ�ȭB�'�`i�e�	�ʸ��
���F�y�h�N72�Q��/"��� 1@�9�y
� ����J˺\^���@T-L	�ru"O�\уlV�h:@i��$N�j�$Y"O�,�f�d|B$�u	.` %"O�d�E␑g��c��/��DZ�"O� A��D��4Y���G��XS"O�9�cĿwԨ�U��W��*@"O�-"Wd@^��V�7i���0"O��1�._� r�}����.P0�"�"O
�(�ɖ"CH�a36� 4h��"O�x�%JD�V����J6P9~II"O����@^o��Qa���(%k�"O�81��V�c=��h�h�uH�p)v"O��%���%�:}B7�]�	P��ٕ"Oθ�TNL)c�R%8���i9,��"O�= e�'\".LJvO�A �H�"O�ћT��U*�i�O	w��Q$"O�9�d���P`ΐ�t���[��O�,�%�&�)�'G��-q'�K�\t�HS��]82Ƅ	��?�-�͉F��9��[�tw���'�lB�Cw���2H(��#K�3d6��;v�*�O�kť�@�]r�YP<hueJ9{0B�"O�EY�2�H��TC��+�&��I?+��|�3Q�E�3EE�6�4���^{�B��������-�ZV��>>���
�JD�r��ӘW�8i����0:,��w�B'_�C䉜5���zB)-1�I��CA�p�S_l��v�%\O�����҈kKؙ��W�D.80
��'�����i���9��X9�ԉi�
�(ł��'�v��u�ʡQ4�c�'G	x�\��	�'W���Â�%JB�hH�c�Cظ���'%|�rFX�J�Y�IZE=T��'��@��ҷN�t��B��r�l���WMf]C�G�|`A�D\'u���q*������^w4��ę��
�ȓ.#B����jn�U+`�q��1��V�$9å&+YL�(5��.ܢ��ȓ�"�`ᆎA�тR�I��p��@Ѥ Q.
G��E�1�<���p�<����Lw�<lҵ)ϭ�t<�ȓ	��`✙??�2�ʈ�*��I�ȓ��(0Q�� FS6�e�S�]`B���_��}�-<hx��@EӺ'-�$�ȓ
���*&��<�Bt�b�	1_E��ȓ.8=�ȋ1vt�]PBl4����1�1@w �Wy�����7������6�R5;�C0"��<�����
�z��)�S�:��Q�EU�$�ȓS���SF\�xv9�� <�:%�ȓ)��x�V���?�Ȩv�� -�%�ȓ]��0gd�I�G���V�J�ȓ1ޔ��"�[��0,1��	��-D��B�ӝQ��D�I��,�Ǣ+D��Beb<2ЀcK�1��kQ�%D�,���@q@�Ժ#�R:Tሁ�p�#D���ݩC6�8%&�3�|���-D���P'@Eh]ʷM�~�8�b�7D��e��m\�*G�<J_J\2�E2D�xS�
`n-�G�ہ6��[0D�`�9&��|�%%ն�����/D�T@���M��)c� 2�p!Bc�*D�H��/Ȍa�v�IW-P��*
r�<D�8@�\�R��hU;t��sB?D���!⏴-2t}`WQ���� �g9D��R��	,�rT�K�1L̴ѩ�B6D�� ���\�%P��C���
�(�a3"Oڼ0G��	�����B��@`"O�9�0y�����YZj�h��"O2`� �A!;��y��O��(J�HS�"O��V�4gԄ�tN�8%
5Hc"O,����{p�X� ��=v�e�D"OJ£ �0��+u.�)hk�m��"O@S2#�)YG�<��E�!�-�e"OT)���9Pr��'Ľ�IqC"O�����QDj����rI��ɒ�+D��p���%�@���1eg)D�g ��qf\h!G\�<�.��3D��A��Dm,��:��\�Vަ���'D�p���[�]64��4]8o[��p�a$D��em�K�) 2��!�D�$D�h��mR��B�˒,$V	�K@4D��{ ���I2 ��4T�90e0D�@k�FF�z��mY�X�؉��=D� Q�����q�e�80��� ��,D����eΫDF&�9rbƈV� ��<D�l���$Hxqq�N:j\�`� D�������T�L�c�C<N4�S�%D�|���X�&a�s�/�"-�q!9D����ꘕZV� F�ܐ<��a1!6D�p`���.�嘗�=���S�5D���DI�;
�nū&��3`��D��7D�L�E�&!�|�W�X#мM{6d3D����`�d���C!�W�4���t*O�I�B	�v5DઃP�M�\p7"O����M��PZ ���Pq(ɔ"O�q���,H�8X��XiR��'�>�86e��٣F$�2)��-�	�'�\�RI��k�	RC:/lV��'̹2�/C�vԚ""�'�v��'�
h��$�0I^��"�(`Fl�`�'@H��&-\R�r�E�=YR��
�'�Hq*a)M�~yT,���F�E&P5C�'��aHe�h���_�,�ș��'�(A�V@�kQ�yz�n]�'�L1�'7:$�㏐�bA��j2GȌo_��i�'� S�*.����'+O�M��'�%y4˒�o�c� �K�e��'*��G�R�!�����5ll���'r�qa1B�/�̵[!�H�]7�,�
�'ࢁa'�W�j�R'L�U��(+�'
(�5���Vy+�T$s��ġ�'X�M�E��p	������{�
���'��`80���+&�L� ��t*0�'�� ��I
$�F�rpf�%m8(��'�=���IHx�'�D�r[���'�^��p�C�F<)g���|����'����C	HR�a�*�k<����'�x�*7�	�|\,5���aW��h
�'�)hr�H�q������A��'>��ͭ(��M1A(_>y{V�
	�'��r����^D�����&r�&}��'�&@�L�
a�`pf�v�,��'��]��Z�W�QX 犪9t(�b�'N�g�Q#$~� [7�6Є�S�'*2�B�a���Ł	%{�&Qh�'m��k���'�z�;�G�� {6��'�`�R%��n�2�1��G�ypN�x�'� ���@�e�:���ڋ{*���'O5��\PG~����1q
h9��� .�C�d�	{����I��{� �1"O��I��^�R��,X�F�9Ed���S"O�U��Q6D��Ik���Yd��"O�t`枹�
�ȃ�N���A�"O.� ��/�F=`��<��MA"O��AkY;������ j��v"O�Y1�=�V�$$�Q�q2�"Oh4[�k�8]��e��̓�E���;e"O��a�`�"9�9��g�H��"O,ic��!��㱋�<5B��
"Op�p���%^�m�djڴC� 9��"O(Ⱡ�1��|�@�9uʮ�c�"O��p�M���|c�@51��)�"O��rP,D$j��m#� �+h����"O���`�%�HA1�k���u"O���R�Ik���3�C�;�\D�"O��8�j M@X��wI_�)�`	2B"O�$%k�K"l�����,рA�"OH��_zzܔ��	>Or��R"O��8q!2T���8��7(�h;�"O<(�K��x�p10�@�­��0"Ov�q���W���C�� S��B"O��h��0q�@8������PA"OY�B�]��-`�,J�,���H4D�,��dH�i�s0�2"��d�(D�����Ѐ_\�ೕ��<�:|���$D�Tb��5eY�ye�P�_1(���d1D����d\_0x�d�5
 � J.D�����A�z�Rpl4�3� D�Ts�d���v pcG)V!JA��2D�����V8@\[�I��hy3D��R�� P��UAH,($Hɸb?D��തD�`��!��eaH3D���(�;R|�9 ���,��|fD7D����G�ĩ@��k�:��'�b}�tJ��7a��)6��e�pe��'��0����
֔���i��t��'��@!.B�a�uaʌ�X����'��S�đ9Ϥ��`ȩC"��h�'���G��3E�
��-�	�!�	�'�xe�E��rw�
ƤY���'͸�c�n��Q�z,Z�$R,\hz���'�"5තC�o��ps�E�I �Iz�'vР%.X�n����d�׫@~<a��'8:�*M%c^� c�΃�@*"1q�'��
v�G�"�*4k0�Ԯ8�.��'G���J�	��diu�	7` ��'�l��$��7BV�хhV,)���'�j��"O'�4���Ā�'�	�	�'�Kf�[�2A�q��"ax��H�'C��VB| fѻ��[�y	�'Kp`p҅�1U���S���e*�	�'�9 0/L#H IU��(
p�	�'z�-��Ǝ[��TQ�)�,����'�a��/E�\F���Ćڇ��$c�'�HK�nW�=��s�膨-:@�'@|�1C�^n|���V�Q�X9��'�ʸӶ%]"0���BBBe���p�'���3��N�Go|�	�Ӫ@shI��'�Z��҉β*@-��!H^��'�n��t	]�5P�����s\0�
�'+���@N�qX�Q���&e ��
�'��5���,Eyt �o��ZMC	�'�P���W�hb#i�	"���� �y:U�Z�F�>��V�+%'�y�"O����MS�+��-�m�8�j���"O�Ȫǣ�+i��j$�z�ı�"O�-+�
8�c���s��(�"O��ɐj�\��m3� �,E���2D"O�\rE��랈ր�"�����"O�lp5��1u$�����.,q"O(!�*�26��³�ŵQ��y��"O�d�^6�xDуKدz��q"OB�
#�ř`' �3'J��
.}1`"O�,H�D�/��YS�E7--���"OX�
ThV�H�R��H��履"OfS6�G����`ǫ3@v0)%"Od-����<]�A��+a~�"O�5�P���6��S
'l*���"O���wcR&(����C*,.Y�1�V"Oh-KU���|�1�,�/Иy�"O,ţ��I�.�t1��d Bx��"O�e9��R`�K�Lכ"��c�"O�����M#B���"@��X�XT��"O��pvI�=0��2cOU.F���I`"OR� �Y�d�h��P�F�c "O��2nD'z�(iH�� �3u��8u"O6��AQ �$���nڃ���""O���PP3v,��֌E�����"O�H�L=r�h�J��`�{�"O�A�Q�Z�^'�Ub���F�.qS5"O�ERp
�������m��.�h�f"OH��R�1ݰx1�`���D"OJ����:0�X�  �P�V�>��`"O�TsvH�."tl<��h�Q�q[�"O
����҈�zYcG��=_��1�"O�����(�6��% xu�ݣb"O�D�B-�<��YN��\��\h�"O�(���e�`�����Hu��"O(�RB���x�t�ӭʁRvx�R"O��2���V�*U� ���w\8��'��8q��	1�z�iC!$�ܬ��'lf|�%Y�m�l}*��=���'
�xA�� ���J���r0��j�"O�83(j��u��T�S*&Y��"Op(ӅL�oG��8��ϕ~2��"O��!クVp�h��NRZ�:��"O����Ԕ|n���fE�N)pԑ�"O@�YD�ƑHI�`��(T*N�c"OB�24*P}�.-
�G��ix ��"O�z�i=|��s��A�{�J�ʥ"O��rH�' ��A�օ_U|��Cf"Om��'��9���T��)�BL��"O�<s����E�G�A��Ӷ"OT�;`S=�"�s�e�_~8��R"O
���	/	^��G�@e��X�"O��h��G�G�85��Im�Ti�v"O����F^�1`�&�]�|��"O�ڄLU g���ѧ)F%^��"O4-�,��2 T!C�j�(��"O�h[ ̑�a�xѨ#�QO�1HV"O��$��Z�I�P��,�1�"O�L��F5]��C&ɖa�\�q"O�L�$�j�l��b�\/3�Ԁ�1"O�ep�l]�^�Z�	䀊�*�,�Y�"O2��c�7/�,����$i2�"O� z��2m�d��чF�X��E8v"OFu� ��		�<l�U�s$�Eq"O� Ƞ��a��5�R�`�$�f2Q;�"OdT��ў*�<U�g#K9>g�#"O.��s�G�c�.��%LЉ
g����"O��e� �6������{!|SR"O����N�o8L�#�	�O0I���'���2R�K��Ԃ�GҷĬ�0�	�+��H��j�k$�ȓ6O�=���D�_u�l0�X~Ņȓ<��x��M$�N�����\��Ex����0|� C�֑:P�		e
�u��O_�I�e�q���)H��C��ϊd&R51�&�`��u}T ;���a�S�O�
���lE�@ T0�m�����42��� (@B�S�O��(���vc�h1��\�	�f��hPRѪ�|��S
#wd@�0e�6	$���Fj�^��Dx�k�\��� �0P��@'.�96tP�y��@9}3!�]�dE*t���QF��,�"埓�Py�/K����2n��b�pɑ�^��y�#G�P�
9��#�pW�г`��yb��b`5`!-��d��cҸ�yr���'8��� �~&���$M'��'��zB*܋Ť���b]�&�J"�-�yB@.rI� W�%����bR1�yR	�I�9{�#?�^d��G
�yr�M�T�la�CH��D�׎���y2�ۆ�t5���[�X��$w�J��y2�^@��x�&��#H]㵧^��y��J�J,��r�����H��B����y�'],��P#����a:%.)Y[�ȓ� 2D�U3��j�e��,�ṗȓ3L
,�QBQ%s�\���emV��ȓ�02�ž`h������cG��ȓV[Q9S�� ���*��)�BQ��OJ��Ză)u�:t:&)�� {����6:�R�ǖ.y\
�$�{�HԆȓ{�(�M9�=x#�g�ze��Rv�Hq,�b�\�S?+�l�ȓ3����ӕ<4|����/=��ȓy�p�R�a�# ?Lh��2k�"���wT�%[�(�.~�3�E�9&��ȓ<n����Ŗj��i[T@(KI���'��<��ޮ6�آ��ms�h�ȓ65�IH4�ʴE�� SoX+�~5��J��At��|�X�`�.�]\ڥ��7�>�� b��|���xЦ4�ȓX�|��kٗMVD�cΏ�n�xD�ȓ/�$9�3�G�i��y��L�H���ȓ'�6��T�xE���b���Ĕ(��P��Xaꝳ�|<i�l��,l���ȓ!X݋e�)`�\I�f� ^~�$� 9�t,�<�����&Co\��͜@P j=��u(Ѩ"'�T\��K�p�b@�V�uF���� L�P�ʼ�ȓL���#��yP^p#��E3
!�$�1�^��$BZ���X�L�S�!�D˚vK���%�L�8���[gG'!�d�S�T��ʘ'�މ�"$j*!�č.F;��%`1$��!��#�?E�!�\6Ѷ�bb��4n� ��(�Y�!�d�$5��a�AT�?WR;���=�!�b��m��G�T�R�����ms!�߿�
5�� �1���ޏ a!��02b ��DͶ[t����^J!�d
dN,��#K��	X����,SJ!��0N�p�W��AAС�G�H�bc!�$�:F�>M��G@�	Q��ѹ/a!�� D���[�M���VD�	�m`�"O���`I�ukB��b��M� z�"Ox��"b_0�Δ��@U�&����"O�uC�&�_<"�h7����"O�U����z>��0ӊe�~�k�"OVX��L�8H�X��-�2p4��v"OA(ƄWp�d�H�
E_��:�"O*PhfBZ�]6���_$H��prS"OtH�s�U�P��MaӌE�J|C&"O�Z�{%~bs�ג	�@	�"O��J�Ĉ�u��{c��q��1��"Oj`3g!�$W�-a+�+A�>Lz�"O&��A�ƙ.�R�����&^ir8{�"O�#"ī[�Xv�Dki`��"O>ـ�Đ~p��S���N����u"O���Yzp���0��;�^�{U"O�m�1C�5�$�fR+V��z'"O��'Xyt�񰤯���)��"O����mн�Rh��N	�~���#�"O���b��Ol�Q-E�U���K�"Ozy�R
C�M{*�p����Y!�"O���V�B�K�>P(�L[m~H��"O�<��)�� �v����y����"O�p�#i/a��(p
�=�`Y�g"O�[�+D�5QrܣRDH�a�B�х"OtI��gJ�W������D�z���"O�lh��N�,��$rq���d9�"O���	 	�,\��c�3qu4��"O̋2,�'2�QB�Did�5�c"O���R�.c
�g2[\�zW"O�C�/^;4�A�r���*G�u4"O0��ݫU�6��'P�8"^dI@"O�-B��́s�Ьs�b�	c�q�"O2�!�щKtv�R#��ߪ\��"O�db6�ކ+i����V'2Һ�I�*OD]qTF¢k--&���N�%3�'3ʔ���=P��;ĥԷE����	�'Z��褯Djz��Y�őrj%k
�'�͛�/�<�"���ă[w����'Ӹ�Cő'�u*���-~/�Y�'/�X��S�ɒ�#�O%?S�X�
�' �Q&M	�D����: ״1��'w�%���Q,	�LiP0DJ%v����'2�+u$��&���/Ե=�v�Z"O$����.R��r0�L�d��"O�����Cu�u�Ӎ�-��2"O�Y�f��9�PRoD�y���$"O���ֆ�	( ������by2`JB"O0��O�/4�֩��`��q�t��"O��G�ԥ,��I��E}pB��"O~���k�>|��@{&��f�R�C"O~!�B�ȃA���ČNo8`Q��"O���L�~Nm��K�$'4�;�"O�� A"�dƲ�+F�ܙ&
$��B"OƼ�0a �m��Ki�87�j��p"OxM�1�O�
V��	W'�K�%��"O9 �nN�5.bͱ3���&U�"OP������䵊p�V�Dű"OrE�6�<���cǈA���x4"O��bd��
r�^QX�čG���e"Ot�	eB׆&������L����"O �����
&���֭ P64�H�"OLpDO@�$)Q���}�)[�"OI����ZB$�!�;XiKD"O� �X���M!Y�0)���m �ң"O����AM4�ID���F#,3�"O���)E< �q��SA�,���"O���$իA�θ�0EF3@��"O���i�$y|�� %Z��I6"O�����V�2A�b�bS����"O>�!�ba�V�� '���G"O4�RҮ@+2�����OD>M[n|
@"O8�DhާVV�P�ߛeW� �E"O С��^�(�����G��r�F�J�"Ox�x���H\Q��E[)8~���E"Oй��D�	�,�C��*s4�"O��� bA�P��(Q�bNV�x+�"OV��šܟ>��(����0ވ��"OƸp���vL�xB�홃Pf�i*�"O���`F�0\�nq�ĭ���@M��"OFYZ��X=]I���̉?"�i*'"O��p �WX-0�K�lj���f"OJ����<,	
c���ZfX)�"OxUړI��y`"�c�A0�V"Od͡�AG0Y�8���ˋi+��3"O���+��:�TٸD!�q'�a�7"Ojd@��j��`�g��+)C�l!"O�q�@� �d�@(0Ӥ<��"Oj U�2p��pR��lꐩK�"O^V��j�9�Ř5*����F�<�pC��;�� ����d߾yX�fB�<!��ۼ[D;��0c���Y��Jh�<q�B�p�p�����|Tȍ�C�J�<��b|�1�aj٨]�Bya��~�<��G+W�*��@(\�Q��ݠ�M\{�<V[�.��H@K��S��8�6w�<!�J;N��mP�"�a�y���w�<���N�!R�ՠ&� i����Y�<���ڰ2hz�!�kϽCa��p�YS�<���i��a�EB�T�|�A�a�i�<鴢ݵ
��T��`H|;ZdI�d�<�eR�'��bFOJ�Il�����E`�<�b�N�Dxr�i��(���3q�Z�<A4���D��dևݾU��e�Y�<3)[<i߼L�Ь?V6��7#�N�<�����ah�k>5�-Bb�r�<AV�G9<DkW���B`��_v�<�S�� "�:���L��I�G�t�<��lU&^V���b�)eG4���@Z�<��g{^0Q� ��"D@�Z�<y��D�q1FMZ�&�8*�<��� Q�<��I�
��)ZwJ��q��س@a�L�<�aD�;����F�|^N�%c�S�<�e���s����PD�p!aP%N�<���+K�z٪�eU*H6�D���S�<Aլ�9!�&�ۄ�$b%\Ȓ�mg�<���C2zcV�#�G�.TB�%�X�<Q��3��jR���p#�Y�<a�pI�Ƃ�NOV�@Wn��o2ꔅ�|�Z���GS��DW/I$�Ȕ��/�!P��2!{bT𤀎��*���6��A��8%8b� ��Y2�.ć�-�ҥ
�CZl"-�bߩZ�܆ȓ%��rw͡��Y��
�t;�8�ȓ+.��
S!Ŋ�h��F.���ȓ��1z��L�cu\�g�^	?��@��2�a��e@������D�HX<�ȓ6����+n���p&"]�c�fE��S�? �xj�.��Y� ��c?u�zl�s"O�yQ%jG�4T1!H�A�2�ZS"O�K4,C?v�#���($���E"O��RD�9U�>���8��4(�"OĄr����r�j|Е�ѯ7�0l�D"O�E�'�ʢJ?(Qb3잯���i"O�@c�8R~<� vh�/4�2ݑ�"O����$� ,���G��@�ތ��"O��I�	5\{��&�v��ұ"O(Y��z 0�HQ
}܌r�"O�("r�[wb2�)�T;�\�#�"O>8��F�hI��m#yTxX%"O*kUn�	%>P���j��/-��e"O�8�v��>{E�HBg)�
L����"O�`Z��׎M�H QU�:���1%"O<,�#,�5x��(��-�5"Or��æ���Ƙ�P�(l����"ONy3'��&Y���$	O�4���ʒ"O�܂�߇T&�@Qq�ݴQ|�(c"O����O�h�؉�]�)o൱�"O4D��Dڱ4h\ !ߋ!ix�p"ODx�2��22 ~8�R�VU�[�"O���Ф��7���`��I��l��"O��"S�3.|=���-52���"O�<5kR�XtL��ua	�~4p3�"O,{���)���sG�H��Ԉ�"O�� ¬*X�s�eӻ5+����"O`�0���X8P0Їg�x N��"O҈�tB�8>� �C'����p�D"O&�JRJ�/p�ܻ�5�4�A6"O4�e拘%��PBէ0��ɋf"OR����hl���fd�x���"O��!���F�=�&�����zV"OZ��F�h�@���-I$�+��'O���i�4�S1�Z$}��)UD��3��¥O>��d�O��D�O6ز0��O����O�8�F��� RN��L^@�Hs��Z�)��H(/����Ɏ}���p4A��K@BL����b�Zn�:"��'#/*Hl5�l(���P���8���06�.�p�Tʎ�Q�������M�������O���'J��᳅�ь��(�w,Ԕ]�����?�
�*�4�H�K��)�� �pc�N?�2�L�?[�FS�$��Ř�u��'�V?��AL�l����*�g�X�áC�l�&�B���?y��0O�8[�o�?Tl �hP�l�Ό��g�V�� *�ED{��H4�r�����g�{�'?�d*�I�}@aυ�I�z%��'c���h���0OJh n�0`l�`eS�'�R0Q�8�f.x�~�d�~��
	)����ЛR��l�E��0+�B�4�r"=Q#!ϿJ[�x�%�M��^�iQ�B8�X�ٴZ"�V�i�rQy2M��4�I5�S/`�TL[�'��0�ɦ�BZ���;�M�L<���/�u /I>6���d+�p`�ǓO�`*�i�����(4"�q����I���Ͽ�t�NM�Y[6%��YZZ=��G�Φ��Se� ]��К��F#py��Bǁ
JHDʕkʥ���s�����h��������0��1�M+�ڟ2ߴi���&"|n��-j�+��ߦ������߬$>��X��?!(O��d+�IR}S�H��,�@�ښ_�ɹ��7�(O�o�6�M�Ke���'f�Թ�04��"[T``� �H>�4�Cǟ��	(S�N��F��֟�������	�u��'2��!�0l�2�L@�����/��=w�@H�!� �x�������n��b�Ν#�'�r����d���ڬNR�<"�	��|0x���Z;�l�;4%{��G�P��8�5�]���L;0��"��1�U�n�T��p����k��$��Iݟp�'����)G<�<��t犦U��ێ{2�'�$�����r����fH#Rj.0�5����ܴ���|b�'��D�a����L^�R�N��H�P2V�u��]�����O(�d�O�P��,�O���OT�e�	��*ueQ�'MXa� �8|@�sV�̉�����Sz~��J�P�Q� ���"18Q��	��QQ8�%���	^����-�@ ��h���3g�NgQ� �tF�O�M F�Î2ў��˪!��0�$<l�� �'*��T>��`p�:,��`�
W�I�, D�
S�л6T��B4�U�@�	P�ߠ�?նi)�6��<y���&Fe�F�'�rT?�+ j2.��q�v�7(WT�災\������?��#�`�����O�g�? �t�R�P�	3(��E"��O��9��� -��P��M-zc?�J'Ú*h�ɁV�B����j(0�B�h��	��M�&��\�"(�ر7��~u䅫ݿ9���-|O��j�� �/�qN��� �~�0��� �M���i��v��;V u�u��6�����J�2��Iן���^��[�I��� � @�?2ӧH�>X�H��dѷ�RJ��c�'��5o�,��"<�{�_�zA��A�M�(�ÁM�|��ć�N| ��#���x�R�C6�4���ZMrhS��\=�̊t�ߚs������IU���$���_HW��ȓaF�� 
�-[ށ���B��M�ȓ�(BabV9Y��+�&�A%�؆ȓw����_�&�¼C�L׷Q���z u�C��dW����X�F������zD�h��і�� j-F�b<��"` ڕ)�'`�nћ�ύ)+��Ն�)���V��@��H��ӌ�r��]��R��&o�L�(����	�ȓR!�Y!�o�6<�2�Q@l:;�x��ȓ�1��D�f��lѣ��S���ȓ8E�Y����m��a3f��\�ȓn?����@�:[JQ"��޺݇�yz���`
L�zp����-�9�0݇�OOF���tɘ�@��M�%�tч�%b��D��"����/�jD�a�ȓ~�XUg	4]���D�~�)��/��xKDꒅ)Ɩ�1���-W٨��ȓf�±##i�*�2nݑV��T������W͎=tA�]�ṗȓv�8�RG@�:�H�AW-K8�.ՅȓlE8Z���V�z��M�]�&��ȓL�4��Z�
�=���J?~a�ȓ(�pA�b�>Hp����8��I�ȓ���Q0.ؽ"nx���LY'�΄�ȓs@^�Q�'&:�5���ß7p���9:<p�f�2I�i��R�GG>���	�8���-r	�a�''Zd�ȓO44 �Ӛ;�V\{`)D:3�5�ȓ12�����	���2$��6y�І�]Ap<���Ȣ邬�ٲ熝��a�ݒa�#6x\��oޱ%S� �ȓ[�4��FH�+Q����Ƶ#WЇ�ba�{� R�!�@�9��H/�҉��t6 -���)N�!I/�m�b��ȓp�ک@P�>xhh9�D47Ύ���y������1��x���Ԕc ZX��T��ia�X�x�QH=�B9��=ynE��G<.��=b����i�n���_�Ψ���DS�E�0��2ƌ�ȓW��A�X�T�A�I"8,�Ʉȓ0>�]A��1����v�]f��Єȓ4|��cՀG�h�ӑ�T�[�~��ȓp&AS�oņ�&�1�Y�9訄ȓ3-x4��ųy�z08Te!����S�? ,%�$A�]������
|6&�CE"O,h!)�5 ��R��@�M"l�""O�Ń@�6F�bRV���dw��C"O���AE×P�|I�UL�r�  ��"OX|�Ѝ���a���2�ҭ!"O�蘁e\�p(w��;����G"O�����=�����
���p��"Oj5j���=� 9!�JԬa ꁀv"O�MX�M��A�hs�jԹdDb�"O��Ò#�*W��� �j���d�"O��$g	�{-l��a�s�>hu"O�SPi=NY!tɖ�p٦��A"O�X�@@�42�����ݘ]�҈ٕ"O���l�'6<� ��;5��\0!"O�L�q�
�T��JW?	0�@4"Of�!GY)x��ʇ�H?����""O�dC#jG������^�%���1"O������c�������^�Z��"O&��`�H={L��b�N@�P��'�<`��&��x���8d��'� \:Y�y�M������# c�<�v����FY+A�]:X	����ʔy�<)`.G
lRl�"+��Chqc!'�~�<� �@�^Q�z�=/��ы���@�<9S�R-#������ٺDUj��f�<1�P."�������H) I�q�PZ�<AE{�Ț`L[41Wh�)d�KU�<��J��k�E����y�\Tq��w�<y$m]���8��kϙv�R|�U�^�<IT��J��"ܽ%�vD�ef�R�<��*�Vb袰�I�� iQ��V�<!hۆF9��c�ƒ��@Ia�U�<)𢅺g�z̨#��
>���3��{�<��*��-#Q)0���f�v�<	���z̺ԩ� L(& t�G�YL��hO�O�d����2����x�����'�t�ɠ��p���xĦ@�Fu&5
��6O��≁&�urC�̓q` �K"Oҭkd`��6L,���F]��p�Z�'�Fk(�	JX����A*z�Q��ό�?�`�{s#.<O�١�F=���S�x���M����&�V��*=���,D�T� �,~o<�p�.�Z3�$h4�,�	%���S�\?4��l��A1 Pi��K=^��B��wή\ dl��*���	�)�nb|�s�i�'d�𙟌�sR�D��eZ�B�v<H�b%D�,s�&#
F���Re$<���o��[���9ް>���n��T�W%V"[V$ ���X���B-�-��$\|�E§��sR���흀i�!��T�/�� ��S�Ai��25�|mS2�?�)��7}� (�\*|Qb�C$D���5�O�)�e�p�<A� Xz��ןtb���s�X��� F��	ڗ���t�e�`�7D�p fF/�5 HBziړ	j���z���䞾J1��s&�f�`Q��F�a|B�O��	�C����A	v�VA`gƷ]�TC䉪2�x�I 1K����k���b"<��Ov"~��_�$��4PӋ�6h��lc	F�<���� *!XXq��(N�J0jJE�<���L�&�c��)y�`����I�<�$iS�e��	�fڢ-d�\	"�p�<��))W����$�ĴP��cż��ȓw�x��aD[h2���H�ntb��ȓeP�s��'
�J�P��Y�����ȓ+y*%�Zz�	K7Ή�	C�	��S�? ���](|�p��lƬGj��"O��D-��)p��@1k<A�8 p"OL$�eS�a}&UJ$�O2r��"O^����8{�L��Sʊ�D-�5�"O��3�'S�>���$X��Th%"Ob����&���ޡweę�"OT�  �5;;��zB�E2!]*|;�"O6�K�\���ʖFE�p'\��"O"!���>I�.��V�6K<��"OL�&�ƎMC|�3@I=#j��sV"O�$
P�.B�6�8�@�5g\�"OH�wk��w��y�"ϋ:tI��P�"OV\���1 �T����[�<�Jt"O�Ј�n��Y���o�?�Fd�"O�Q�9dN)Sf�[3D^�uw�h���0D��  G�DC�A!zb*��ȓ2W�Kc�S�`���Ǥ֝E�X9��E��xSW�=��R��W�8|��O���3�ķ6� ��m��;S�ԆȓA�A˰&�KP�Qab�b�`��v�&����C�i1X�5�H��ȓz8qۂ�+�hд�2���l���U�F�p���sk�|1����!�D1ע5Ҥ\���q�� ��c�Ġw�C�G�~�[T��
��ȓQ�}��ӏ�V�f�Ӕ)ۺx�ȓjLm3BU^�-P�
�~|����,\p�*	�>�& �7��C�@I��5���'�׍X�Tu���ҳޠ��m��=�Jͨ��<yTe;գ8D���@M˘%7dܐ�  � exG�#D�(#I]�_Bʱ@fd�ـ?D�$�(ƫB���h"-U�|1�t�ҭ9D��249n��hy�E(Z}�6C6D��i�¸'.>�E�����t�3D��"�pz�ؚ��"K:l�C�1D���H �l�8g��m0��s�/D�,jՊB�/��ty�i[�Y��@&&0D�4�&�&'o�t�$m؜UU��3D��@��_�r���-ѹ��a���1D����
ڋ}k�h��c2��	�� 4D��s��F���k$m��"�P�"g�=D�x��eR�/D4$�q���Ac�!Eh<D�P��K���t���Ԛgk��a�L;D�x���Ѻ2�0O��MR2%9D�X�V��?Z�=Rl֬,�\Q��5D��xơ�H�4 `k_(nF8�#��3D��!C��$��=�uě�i��bA�>D�`zG'�0��Ha`����'$1D���éN��A� ��p*U(.D�|ї-��X��Al�@ql��1D���&�td*vM�aN�H����'�~�Y��D�Q��lD�*��2�'�\`$�T,s��eC$�="�'����
���0Y�d,�tz�'��(J�O*3�uB��R�l����'�����
6\ܸ�T�+$���'��T�(�xҘ:���yQ�y;	�'��Q�'�3j���s�ߩl4�p��'�x R���,!�Y���Ѱa}>�+�'e@峗�3N��eB�֫\�̜�
�'�&P�I�6U;�$���3"_�ɓ
�'0p��FJ�:�a1�&F�I�	�'Bh���
�U�C�@3Ij��	��� ��#����4�3�EN��>�`A"Oh����ZW�͑pO�!}�LQ�"O椁�%�G�}�w.K�Hj��zT"OHq4�Ǣk?
��al�?y`d��`"O*Q`�D@<=�B^�NX"��"O�yJ'I�[���6߿wKPi�"O�1�d^=#Kn��d�C#F4�w"O�MJ���-(�����y΁ �"O�e��V�z���n��Q}�t�"OdB2���.��0�r��	Ry�H��"O:QV��"($h�*���__��P�"Oέ!R�]'%�$�Sn�$9}]T"O�̓���
`RjQY@� l�	�"OJ��CLY�*��@�e�nd��jC"ONYXBH��1��� g�	ba��r�"O��AB@-l�2p��T�U�lQr"OL���05r��"�_�?\���"OB=#�8����B��!W4�Z�"O�A#w㞉u�L���d\ �Bx�"O��#�̒�<k�!��C^�3�&�"O8bP���Ѭ�7��?I}��A"OH����E��A@	{M��"O�����T�@��t��a�"vn�(6"ONL ��8q��b !ڄ5YJ ��"O�q)��ȇ+��H%n�r:��""O+�ŖX�VU�䬐�_;�e3bD�p�<���\�|X΀����<Gt�:�"@u�<��˔_@t�*�)E�2�z��� �Z�<I��1Q�BaPc@�bJt I2hO�<q"��bZ����,�CۈȐ��
N�<ل�J'��u�ri9�� g@`�<�q�,   ��n��8ыR�^�De�)ODDzʟH�7?p��tc��:,r%͕&��aC�6�&�'���'3�)�ӈ2�r�H�0�Nl�J��1w��8�iD|�1 l�5ǔ�cP`ǔ��OV9Bu�Y%i��(�ӄ&�`3-Q� &@�sa�\Ę��O�rh�`�U��)}.D���M�4@��(�Z�M �����ON�D�O��|F��h���ty��ܿb���#�� �y-������R6�h�j@��-���by2���:K������H�,�����J�wFheb�'��Iڟ�	ԟ���S��픈j�
��g8b��1Ee�(@�n��A��n��%A���ގ7��U��	oxaBt�Y�F��Jsl'#�]��B�5sJ,��3$7�N�����ǟ��'&̀V�؈`_\M�c�H4���sN>��P1�H���,.'X5*��Pb��t�����?���ќ@~�h�ׯ�a��HQ�h՟��'KJ��!T����O�@s�% "鎀SE��t�Q�d�O���
�bк�9$��,(	l�c��9"�l0�����r��() �ԃ��T� �M~R�43d�ѕGƧ)��i#(��i�ZE��n�>K�.�o�C���)���@r!
�O*�d%�'�y
� ����7\v�E3m���&"O����W�b)��aL�6 �T�	��h�n�c�@Q�$�Y9�!�/��ya�'��X�u�4�Q��H!k	-rƲ�;�OB�~k&���(D���Γ$an$ �a'�~��صl*D�4�d"G/7ÞtYr�ݼLE�D�'D�h��퇕r4�0�@%Q�5�+�3!�6@r��V�ڲ�ܕ���GBA!���.C�>��q&!(h�jsJA�`9�	&'{���DX9 񸨓�3�*0�&J'+!���5�TeB���5�*{!��ٛ찕�KK��d"���(u�!�d±B���f��v88�s��*\�!�A#"�=;&lW9ip(F6.��}�Ǚ��~��F2�i�!�$�P �N�Y��4�ȓ;q)���.RDF�T #�8���I��!_0:00 QCV���ȓx�^��i��N^Ы���Qt���j^���g�(�<���@�>��ȓ8k�@#�Y�����"�>28E{�����4�Җj[J����D�9��=�"O.5�pk�:B�p��O�>=�Z�j�"O$���L���`Cb��T^��"O���"oO�9`�����+��咧"OL�I�NC�7�.���A�#�(�s�"O�͓ -ėm;4Гł!�L�1�'/��"���4#�(�م`;e8њ��=#�N���)��7鑣-�5R%��;e
�ȓuv���T ��n��pK]7.��ȓ~���'ٰe͌,ipƗAl���ȓy�(����� c��x��	�1A�ه�{Pj��D��S�&;�b� ]%���V�3:j4�cg"Rl��:+\x����٫#?¸���$II����;;�H,��̶ 4�5�G�a.�)���X����?�����@Bm�=;Ft��IJ�xK�(BJ��*�l�2�bi3EEݏU��`�0gEM�'#�Q��!�"q���Ї|�N�jc��K޴U�'��Y��iqE6Z�
��p��~�'�l���u��V�>�)�ʲe)c��#E��@6�A�@]�Ie��P��D:����BG�lxb(�O���'���1ƌ�e��dYV.ѩ���*,O$tKdb��a���@�O_��S��'�b*+SD��@��2,����"^�p�BE�^)D��3o�b^:%���i".}IE�T)�1��Uqg��}Iw"��%!ܨ��=O�<�BN\�dH��h@E���@��d��!���8t���?\_��@���Q�Dؐ����hD��	?���Dͦ]�,O�O�ӌ��Ak��/�V�b %�j�\C䉓�jБ��	����x��EvL�=���K�j�(5�˜E�*m�or[��E��ԟl���$'v�Y��Y�����ğX�ɀ�u�'k6�h�f�T�L:�	N}����H_8�d�)�>�Ж�J��3Z�A�	�@ޜ��h�n����'��?��b��m���)��Vu�����-��������em�Į��T��'	@,k���?���ds�ؒ�AS�ܕ	�]����i�G2D�Cs��U�yK�oД��0��O0,Dz�O��Y��XVI̽t���@M�������- ��lA`Z-s+���I������u��'xR6��p���~�VQɂ�*��	�6�Ʊ� ����M�x��I��S%��B,��(Ot�0�"�"c���X���Y'V�ne�W�A�mT����mI=eV�k�ɛJ5ܜA�{��%�?1��{IN� 銱Tn��͕��?����'��>G�RW4�
V�O*p+ B���<A�706�X��բx��YZ��@yr�n��$�<y5b�au�F�����1�.a�5+�"7�H��WF�{�6Abb�'���C�'u�'���2��!���]3S�!�ħ|��_z��x��4Nd���m3����Ώ%oȚ�-�D=,�ȣ@�$+��h��W�L�0p�7�ԥ_KLT`��\�'u�a���?����N�`�X̀T�$D��ɠ��
��D2�O<	���E/d�,(5F̀ s:���'��ʓ}P���3v,�ՠ�"��ݖ'U�i���'t��_�4�O����'�t8k��R0�6�J"+�|d\�P�'Ύ��3��t;�!J/{t4��*��|��>�!���7K舡�U5;�6-��f�|	��M�/ڄͲB��	Kp�(g�Y��H��X��LT 0)�q�������4OJ��1�'������S�? �tz��G&T\����2#N&ȹ�"O�TY���
.�h��r	��BP\t��I��ȟԥHP��n�h���a)0�L�8�c�5{�b�$�O1��K�}5L�i�O��D�O\���O�����h&� Ka�	�L^$����N�Y VP�F�B?#rJ�租�~v$�'��'V���J�3\IBc��::��ɡp����l�@"�2��`�����)H0s�XN��H��A�\�~9���+k(���e�/?I$A�����S�'L�d�� ̊�a�
r:�Tc�_>/!�ē���\����:7�(�RΊ�?G4��|R�����o1<��j��}�@�QB�G7�b ��MD�[� b�O��$�O���O�a>a���Z����+)�e/~}Q� ŏ��Uf��0/2�z��Z���Oޠ�fI+C�ȐCK���v�@«����)�g͍�lYk����EF~�-Q��?�B	�Wb�rV���b\"�ça���?ٌ�$3����9���o���i͞z-��Q�'�@�`Ɓ�J����D5��=�,OԠo��ܕ'q�d�#.�~����d�ү�6q+�@ؒ_�d�1GB��?)��X4�?���?ydm�2SR���F� >>Z��A��D&�4U�I���"w��!��D1��OhX�@G%y�Y��B�J�˧x�j�
�B�O�l���Y����E|bT-�?���O{���gl�{�d6����@W�ԇ���	=�u�T���a��f_-!�����RyB�\�L]�o�#\і��E&��d�On�d�O���OZ�'�?!�O�x��M�6$��'�mr p9+O��!g�ĕL�'�V���DI���
�`��!�����E��'�F��	w��f��ɈE���pN=TS�y���g��Ը���I�/�b�D�O����O���)D��9���z�g��&%�M;�/J֦�	:ବ�	�<�B��rnz�=��OX�Nڐeq��H�H�Js�0��%Ѫ�	��?�4gH��yұ���d�O����O6�Brx�� {P�+ď^(W,ih0��O`�$0@����r�H� �?7��P���'J�Z��F�N�H�tH��7�����'lfX����?I#��*���T��Ox�)�Ҡ��@�Z����<y���V�[矘�UJ�O��$U)m8�������?7�[�<䔝�V�&'�L����*�*���Φ�Γ{���	�ّ�<���?���YY�y��i���6��H �ŲMG�q��'�&����?qv����p�tK' ��?�mZ<A�|4��	lU��S-��q`$MzB�G��M#��'b�Ő��?yv���Sܟ����A��ѣF�K</��a*�p�����4y�tݚ�'B�}�b�i]�6�����D�Пd�g�O�QcEmԿDv�{ ` �Y�8LC")�Φ��g(���'V8��y����By��Q���h�=L{��I��\51���"OxA@T�W�zB�0MH �1Z�i�"�'1�'<맯?Q���ih���jF�`����cѼ ��<sܴ�?A��?I���?)���?����?	�O���ħ�'a�)���B�r��Iݴ�?�*OB��O���O���|Z�#\�H<�4�A
�1��n��,���[�l��͟`ь�L<��$�GB���&�P({( �C��i}��'��� V��Y��p4�B.m1�H1H<�	���c�*އb��*�Nݰy�D~����?1r�"�#h��<��
�59P�(0�>D���q�ć2�x��@�0�Qb�?D�2��n�|}�rH[�wnF�ڗ�<D�����2f��PJFm�&5�@b�:D���&OU�`I�ۅ�Uv ���8D�T���SzNB�p�g�9���"�:�?a���?���?y�I�'P����ъ������`d�3=���'��'"2�'�Z��'�'� ��1D�0iW���V�Itt�s�v�����O��D�O����O����O����O�hK�A7�r$�ʝܨv�X�y�I韸�	ğ���͟<��џ����"F�o�.$ R�K#����pb���Mc��?���?)��?���?���?���A�[@h�"�C��:i� �^�.{�F�'{�'`��'�r�'kb�'M�H%��]!dA�#7Q4��UD�<;[�6�O ��O���O4�d�O��d�O��X���A�� �4�9RG�R�fm�<���h�������՟���П��"(��3!I��V,Id�!]
� �4�?���?���?���?���?!�&B��E$��4�ؐK�NH��$�i���'��'��'5�'���'���[fEJ/���;F��M��]ZRIbӺ�d�O��$�O\��O���O��d�O�Hk�X��@�q�%nL�X���æA��ߟD��ݟl�Iß��	ß����(��n�~b���o�>0D�qc�.�M����?���?	��?���?��?Y!������Eߪhz����= _�v�����Zy��ӵbD0@Ҧ)�Q�5L*/�8o�H������I�?e��~��iD�n�$7*���	=�,@;d�]�6M֦����d���i�O�1zP�����DŃSД��iY��\q�#���f@b�DH)�f��a�����=�'�y␄@A�Q�5J	GZ���"�?,O�Obam��q=Nb�� �)�@
ٕ� � �G��{*�0�dq}B&y�Dn�<1.��T0 ]�[e�u�R�k�Hh�RV�<i�� 2�}�$#?�'3
p��vBC�y��1�2����\(ʜ�F��,��D�<����h��D�N�15!^���8'$U�Gy�F��7����ߴ�����GĒ	D���6�˜�$�	�B�Bhzӆqm�����R.\��o+?I%a��\HP��^���(`X�3�>��X9q'��Z��=1���d,�:w��)�4&�%s��೤�T�j-.�L����>̘'��l��+��B��5Ό����b��z}�h�L]m�<Q��)E �X${����,E�m�7&�9Ef�ք3/���s*H(S	ͬQy$�1��C.�M#�	�%Ib���k�'1�X���_!X�L �BO� "���5���L}���[!�gj��>/6��F!9�c�h��F�;�)����z�i`�A�kyFtZ����U"������7dC4�]���2�H�pj�{W�RbGט�AȀǀ�1��дcL*/b\���ԁ_B�s/
0t���b�3��,��o�6��<#��!E�]#A��3���Zs��{���E�0��X��.�#���6��,qg��B�jAkЭcD��f����7'J/2�ΔU��'x2�����6MzD�CmN_i "Ǡ�J�H��X9Uj�p��a�:9�D��:��0$���8A��2J�xP��,Z:Qf�*0i�j�y	�)��Mcv+�OԶ$�ĎޟX���)�N�3h���Q�I�}�0-(fn�L���"�-�s�F�xG�хl�ph4H�%D�*%P�/&/Qh��hQ�c$ ��\��1R�ˇ-,�E86f�ZM"�y����ؼ����Ħ��	� 24lŨ&��%a�jI�2�\͋��˟��V��˟���BHf�$�OŔ�1ƨ�&8
�f���01�'�b�'���'H�\H��'=B�'�B�O�r�2&�/�ص�#�`���p�|2�'�RG��b����y�O�ĕ���^X���Rd�Û�Y����?���P����?�(Oz�	�O�/\
N��u�.<���gS�}cN���O�$�1Y��"�����?�����&�j{��X�%��'�B�'�2�'<�t_���O]ʍ�u`��T{�8�D�.R϶���'�h�DhW<�������C�A������E���VB���O����O�1	�e�O����|����yRŒ�`��0�f�҃2�`X�aLN�h��D�<��W��'�?���?f��
1��9Y�#��19�	�1��\��O.*'�Op�D�|�����1j`ջ�K'>9�$̃:�*O,���/O��	؟��	ן��IП,�P.G�~�.�k'�9t��0��O\(V�l<�'���'��|��'��hϋ#����C�G�h�B\)U�#3�6ѻ�%�����O �$�O�ʓ`�Х��O�r�"�)|�p��F�Z)|��-O���O��d�<����?t��q� ��Sy����̡7�y˦fBKy2�'���',�	�$�Ҽ�H|bTnQ]@ �%3f:Ԩҕ�%�?���?i.O��D�O�D8���W�0�e!��4X��p���'8�Y�������ħ�?��w��U �,��:�q�ߠZ��I�����$�Oh��݀kJ1�l��z޹�p�˅>p�Ⴅ�˂MƜ��'��O�ʓ!��%�ÿi����������D�&%L�h%��o��[VB�rB�'���b$�)��g��Z<Ԃ��д�p �w�d~�,��(�7��O,�D�O~��Ba�i>����9G�<0)�lD��DE�7�ݟi�cASy�'wB�Ϙ']��.f����(�&�]�� @Oˬ�M��?i��%� U�b�x�O
��'#N�Kg�԰v92��T��i�Rx��S���	��3E"%���@�I\�q�'c��%)�#ţ0���#7��t�I�FXL�K<�'�?)�����ӊ �$�s�hЃl̪Ġt�O�<XD��O�I9���O��$�O��S�����.�#�l��Ĉ��H��@��@.)�'�2�'PrT�L�������Ӕ3f��Tf,p�l�2���T��c� ��ҟ���_y��ݷ(�T��]?gzBF��-*�<�2c��L������	�D�'���'��S�O2�tk�/�\�� ��%����<����?q��� %p��E$>%k�`��j�؃bj�� ����N۟|�	��|�'m��'�X����N��8�S���El�,I%����?q��?Q,O��0�_`�Ꞔ̻:K�\c�O�r"���&�{ &���uy��'��k ����5,��Q����uZ�k��]^��D�<�W�խ4��]>��I�?�(OƨcF�Q��h'{op���'gB�'P�E��V��'��O ��Q����J�a�]I(��B�'j��(@e|Ӱ��O`���x�'��ӗ)G:�C��R�&4Aw&�Y����YԔѕ'cb�'���y��'���{��U2����-e*���hӂ���O��$B�R�(%��ԟX�	0,��-��C�xH�h�F_2�6̕'V��'M�4q�y�'2�'
�m#���83 ��`��2?\=R�'�r#��O���Ox�ħ<qũ�m�����^"
��Aq$��?���>�.��<����?(O����8Li	�F��B\IP�9KL���g�<A���?9���'r 9h�R���2,d���J�:��]�M��On���O���?�S��&����3��z�D�6��4��E��I����IG�����N
a��ݹ��O#V[Q"	g��P�<!���?�/On���6'*0ʧ�?��M e�&eH�BH43̽Q&/R9�?Y����'��I<f �'��Y���ǷP,Jq@�IS8[�F�����?�-On�$G�@Yd˧�?����� �Mz��O�v\9ŀ͒�,���ı<�\X�'� t���c��(�B٦7gz�ڥ\����~����	�����韘��Xy��� x�u��/�6U�A��!J��	ԟ�
d��*y�b��>	M�a��,�D�������O�|��O����OX��꟢��|"��LP��d��wU(a�
�����b�nL���_m�S�O�b(Z�#��p�Š[&����!)uX��'B�'Y+�T�����I�<��نQy�P� P�kR�k	 �nb������{��럠�I�<ѱ�݈�Vix��zdT��ggB������l��ŕ'�"�'?�$J1x.i�Q��NS�H
E�м]�	��Z��+?	��?�-O:�D��&m ����U� T�S0,�?Oz68A!&�<��?�����'{R�AD�����,�:
]S��%O_�x�fA�����O���<���E�O�p��a�6YDA��.˝?�RY���?���?y�R�'��i���ʽ{~$QC遲6��{��%S[HQq�]����ȟ�'�ң�&0�S��\JP�ɝ)L���?"�V9�F��X�I{���?Yĭ9 ��P�Oڍ�$��/;��Y��O^D�l���'�]��I�m� M�O��'��$���%
`B��h�׃�&]�Ox��_�U�(���ԟV�C�
9H<(�OƔC�&h[�$�	.6Y�	埜�IП���ay����H�p��-n�6%�g��a�џ\�r�Z�t��c��>}��KM;^����)����G�O�\�C�O����Ox������|���"�b RЍ�
�d0K]m<��<"�X'�y�S�O���E��������թ :/���'���'�f4��Z�����	�<��$�J�De`���) �����e�|b����JDe����I�<�Q(��$o�[�Rmv�[qN�������'�2�'�2�$��.���w��vZ�JG	��!��Ɋ%�퓖�"?��?�.O�D23"��dLh��y`3��	@K.��b�<����?�����'w��Ë?~)1 �3o}0K&�ĻtWd��H�����O��$�<�����O��yzEŘ.zv�b�l̜^�U���?����?ى��'���x�H�0�.��L�G��tCD6-�(Q�_���̟�'�l�Ce�S�� �ɷo1<); �PP�Ψ@�������v���?9�C_;O_�`�O��5(F;y!^$�+�3�8���'��P����%h	�O�B�'��4	��y2Ƥ�DK��v �dP�O���Oq���ԟ�I��	�(=��	vؗ��P���Ɂ;\���˟P�IΟ,��Jy҉��A��A��-�y�b=��n4�I��|:B`ʛ%�Db�b?���NelMҔ�&�Dac��'È��D�'���'.��OE�i>���+Ɋ�!�F�r�贛��T)fd���@4�Pf1�)§�?�҈X8W[$]��
r�r�z�kO��?���?1��a�<��-O��OD�Du��CW�[�v�����S��[á��j1O��	gC8���O��D~�tR�#��fPp+A�_z���&F�O��䎸2�0ʓ�?��?A�y"�J?rk�r#�Ło�@�����#���<@x�束(�Iԟ@�''�O
g]�+��Y��a팵;�0	�T��I����	W��?���
�=���D�� ��](V�D+���#�_~��'b[� �I�V@4\ͧ�*ܨ��U����#`P�!����ϟ �	�t�?��� 2T)[���:E�kg+g���5�м.�8���?	���?y����D�=np���O��.H��)�7�mFZmsCE9��$�Op�`���&��H!�	9}+�47��|��BP�_�Z��F��?�����d�Ox�"��|����?��'?�T@`a�X��5S���&I�ѻ���'
�)�3-ݹ�����3F�t�;
\��r��4��Q�����|�
��	ʟ������Ny¸Ĭ�uAZ�"f�����T�#�СY(O���C�0�p5�p�����/�ֽ�7�Z�6O>I�$��L�B���y.R�'H��'���S������+%dO�3?>���l�0O��C����y ���`�y����O���N�kG@yv��;S�*�)q&�O �$�O`�$S� h���|���?��'o۵@�<���+�ʏ.��Z�N��^L�M~B��?y�'z�8p��2F:إh�M�,v}����?��	���O �$�OX��*�oԬ:�\��_T��� �X��p�!������?a�����O�P���<-X�@I7���>�[*бw��<���?�����'uB =�\����E
:*Vd0(L<���@"�����O���<Y��wyX��O�n����Λ:t�jTb�<6����?���?I���'0��0��L� 8�-� V@�06H�EM�8Y������$�'���d���h����Z�nTg�4�ZIw�����Ia��?��	R���H�O�u`��T6��=�V땣P.p���'�BY����yF%�O���'���IW̀���E?jX��(�#~��O����tQf��t�ԟ ����K ����6�C�%nDa^�x��q|������I�x�S_y��S�5���
��]�ؔ�òf )W��I⟄�t�%~[�b��>A�f�Q�X/�U�be�^�j���O�����OJ��O �D����|*��р �x�!J���6cՌ&|�q@C�'�4��6dԮ����V��0K�Q�G�5HJPY��ǣB�:���O�d�Ob\7��<�'�?���y�`E>w)�U�p'�E�q�G`8(���<���V���'�?9���y�A
<{�� `��y-���֣�?���-/OH�$�O��D>�I)�I���;�,�൤�#<�n�� Jmm~��'��[�|��
�%³N�F{�Q��E�6�8�c��fy��'��'��O �Dʀ�8tH��Am~a �GƢE����k�8kq��ǟL��ly��'�ּ��6�v� ��	�m`!��O�ELQ��'�'�r���O�A���n�䑡�T�}��▄�'1����<����?�*OL���\F:�'�?��"��dnDa@ ����
�?!���'%�8'w<}�I��K���86�44�����^%���O$��<q��fZ��*�����O��	(},�	��IޥRO��?����ɔ-�����'0�?���L�L}� �ӵ�%��<f�I۟X
ǎ�ԟ���۟����?	�'f^��c�=D��љ�)^�=���U���,��{Ԉ;�)�C<�+�aT�.�f��E�t���䃀 x�D�O��D�O����<�'�?�%aIF��̀�K�_�hM�'��?�ã��GFJ��<E���'�.������s��]:uJ��YY@���'���'�R	�(-:�i>��	���̓/*�
RN��U*'$ÆS�%�O-�Ʉ5��%?��	ɟx�I,x-Be���CNC��P��<=�xL�Iğ�ˤB	 �M����?���?�dQ?i͓d	�@
%IR􄰐�D��n�8L��/m���kb����ԟ��ן��z�D��vE��D�:z��'��9,����'���'���~�(O����m�ЌrM�z��쪠,ƣ%������O��D�O��$�Oj)�j�Ѧ�A%�-�����K�4�����X�	���ʟ��IzyB�'{��O�d��!-� d.6��D�#(�Ae�'�����1ob�'��S�:�ذ�ߴ�?���l�Θ*�mJ���Ei�,ơy�1[��?���?a(O��dٌ5��O��D�F<�����ב?0�I�TG5�3L�OB�$�O���2�P�m��D�I��H����DC*~�d h��:d�V��	��\�'�]�����'R�����ܴM��y��g�Q&d���/X
�B�'~��V�<�7��Ox���O�������DI�}�43�H�t�`V��Y�˓�?��������L�X��@�B�|,"'���2��L�O�
��������	�?������������kH� 'ϻ`����C������ʟ�'���J�S���/h��5`һ ���H�D��M���?9�klN�����?��?���?��
ÿa߈<ȴ�ށq�&*^�?!�����P/P������On�DؿU,�����.s�5�­ߧ"�"���OD����Ӧ���ٟ����p��0�&��x(a+����,�mhʓc�:����$�O����O����O�m2�$M�a�7CC��v`�L�Ln�ן8�	���	���)�<���h��T`&�	�Lĸ8+DKH2n�4h����<���?)���?����	ˢ9�`lZ�2S� ��A�&�~-�&�	!^di��͟���ڟ�����$�'k"oƓ����U &�B�C�Td�,�ѶDY4�����	����������؛�MS��?�'a��tc~))����8Z �ReM���?A���?�����$�O�%zG>���$�O��Aㅚ"�HYy�B��NT���MP�d��d�O����O�QcE�Xڦ��	֟P�	�?�tO�0L-x�Y~��j�]Ο�	}y��'W�xP�O�B�'R�A��O�t�cϋ(@��117���l���'�b�'�DH�Ѥf���O��D�j�	�O�h�V��-R'���A�<I��d�$���?�(O�I0:�կU%蝹�- 6��Y�mH՟��d_/�Mc���?����*���?1��?!�! v������19�qc���?��������yB�'�8�� ��رð���,���sӴ���O��D�/���i�O��D�O���O�`��m&H�@�0�)5E.ڔ��Of�$�Orl��kD�u�:����)�OJ�D��KY~R��B��)�����*���O��h��A��������ȟpH��8��	[�2�3 ��KS�ɱ��-� ��܅|-.�au5O��$�OF���Op�ļ|��`��Z���`7)�j�m�1M�L�;бir�'*��':�'��D�p�Ү�%P2P��r ��Z\T@5Lʍz��<���?���?�� �1�E�i>��$�	b�%{s����1����?����?1���?�������O�JG8���'	=eL0e�@��|r!�'�O��$�O���O��D�O8p�IѦ��	����C��9n����G�k=8D���ğ���Ꟑ��ky"�'^J(�O��I7A�F��3��#t����s�Өq�M�3��ןD��ޟ���<J�a�۴�?���?Q�'0�&p@w]���q�Q��`V�����?A/O���	-p�˓��4��)[�.
L�L��F�H�A���O����O� r��Ԧ��	ܟ����?�Sڟ��]M��8	�˅=(/,
d�jy��'�
l�X�����O
�� �4��iA��2s������O��c�O֦=��������?���\��ݟ����#����Vy  ���G䟘�*�럀��ry�O��O��M�W�>���7+G.���^>3�6m�O����Oj��3g����d�O����O��d��s���׫�ahnH8�22����O^˓2�P�pO~r���?���$�2 �A��r���!$��y���?A� #k���'��'�b�~2��� ,�0K��`d���ꏯ���CW�@2��p�4�Iܟ(�I��\�	c�t�ȊA0J��@,��&�����T<u�a��tӊ��O$���O���O��I۟Pk��Q�4u��F/YFҶ�ƗzK�	֟����d��ݟd����&a�-�Ms��ˋ04�� ��i�\�*�#�?)��?���?����D�O���;�dxæĜ,Rj�$k�I�Ƙ1���矜�	"�����ҟx�'���c��4�)ܨs����������	B��s�d���OΒOf���Oni��;O����%6�b�j��F�l��<�	Ο��Ilyb)K-B�B���D���Z4n[�P�裗ԓq�̅�&�<�$�O���ߊ=���d+�ԟ�eȧ`��L�F��f#�6Bdr5�'�ɛ[��xش��)�O���L@y����ظrG�g�NA�'R��?9���?�D蝜�?yM>�}�Q�ێ~��7H�J\I���Nꟈ�R���M���?A���E���,G�0ҋ��~Э9N:y���٩���=� ����$!3Eͷ����_
v��mʀ�M[���?A�vq�G�$�O��I,,�AZç\ ��ШQ��-9 �d:���!T����d�OT�ӮO�H���O��RDj��^�~<����O���)�d�I韌�Ip�	�?�)��%P�2兌 4s聕'�6 �'���ܟ��h�
1�8���)��"'�ۃ$�9 i�����?y���䓅?q�&|�$)U [�2u1u(�.bS�i^�?�-O��$�O��d�<	�D3q��D�S#�Ua��_�LrN���W9����O���)���O����f�D��0�����޿pt�a�2��` ��?A��?�(O��*���v�6Qh�)����p|���C�2o��������&������p��
}�$�'�r����h�ԝ2�M%ao�����?9�����_�n,e%>���?Ɂ3��K��h�̈�CdN$�6�AO��ϟ �	�	�	M�?�!�]l>ȋd�;U�ص�)�OX�C��:�i'�ǟ�ӷ���>��i��GM*q$��ˁV�'}RI	�m�ɧ��Q>%�^mچg�/~@�Lu���ٖT�IA�t�ߴ�?��?���r��'��锢d�佃4*��)�&�1j���N�yr�|��I�O��Y�n.
.Ƥ�'(J�31$(����ݦa��؟@��;0��}��']�"��H5���+��X��rP@���O�t7��$?E���I�6��!��)��[Z��kQ�B�>ŸP���誡bY�ē�?�����D�4]�Wa�-]�r�����).��/O`�����O�ʓ�?����?�*O�y��G.N,*=���&b�xh�a��o���>���䓪?���%kR�0t+��
� �䖀2"�	�l��?�(O��D�O6�����@��?	 Cn��gp���M�����1ϲ<!���hO\��� N���G�?��|�"�:z�p��Q^�����O����OD�$�<��@P�O\���2���N��"6��4X^d#R�'"ў����"����ڟ̧%A��E@* +��@�
�A��9�	L�I[y򡙌.�����dw�9�F��_�8��D)K�\7pH��*�IΟTB��埘��W�'p���񎆇�R��sad� ��y"
J��7��|����\���� $S��4P������<���
nz���?1�����,��U/��"m��"��>�R�_�B�'��I�?��'��	2
��PF	�7�H�Qr��-[����?F.̂�e+�)�'�?A�$X�x!�D�˼-7nekDI�|H���'���')&qX`)�4���$�OP5����ꊕY�cͽ�F�	��2�	�#��c����ޟ<�I�]XY�[�rѤ���H3F�}�I՟D�R�ݟ4��v��'d�'W8I�ӥŒ!c�P+Wj�A�NQ�`Z� v�j���?Y���?I.O��x�Ңt�t�W�
�?vH� c�\#S�� &������%����៰8��^�h�ؑ�J:��9�B���%:c�8�I̟P�ILy"a]��|���.%��M`"�H#X%.=Ya)��3�	���a�I��I= �R���kKU(7+[�er����Y��˓�?���?y/O�@�&�K�S $v��P`
�u%1!l�.Hh�I��%� �	��Q3I9���n�B�'�mvl�A�ԄA�����O���<��l�/��O��O�� �S��&8�jŖh9FQ���-�D�OD��\�qO��SN��a�N�^Քst��9	[����<�4��(䛶U>����?�:/O����?(2B��"�����Aj��'2�'E��K����R�oIE���,�ب+ 3O;Ri�<e7��O`��O����a�Ο ��I1]o6�"�@ `�&ᒑ�Z��P)%�S�O��M]�Oކ}�"�ܝ
�hH!'���7�"�'���'^4h��'�2_>����<���V�YC@(���B�5~�-z�c��b�iC'Mw�ןl�	���`����dI3�$�.��h�#D؟����p(|��J<�'�?����$�94dN�g ^_�Ti·.�p}�I5[,jc�����\������	g,@�E��P�F%�?~F}�5 ����Isy��'��'��'��P�͂`4*կP�`؀��4MY�eQ��O�I4MX�ED�^���	�iǊuDX<k$ޓL�DP#��ltᅡK�"���"	F8�P�Q���?����?�K>y���?Q� �$�@*ӥr�ʨ;��"O/Ե���'���'j�'��S�?}���?iu�E,W�YQ�I�,;�%���K&�?�����?9Fɟ�H���sфU7\��!H7b��+���xB�ӆ �&��#2@H����2�'X3����g."?)S��Ym8aa��3���Z���E�'�\�r���}h���DMU�~ܱ�H��x��q�޲*��M��oj�^(j�I�۰���n�!%�nA�n��l�Hd��դ�N�Ai^��ȫ5
�&7 ��3���Gק-�U�B#M</���� ޴BlL	qNS B�l���-�3|�bF�>;������@�Q4��X�X%��P�LZ,(�������?1��?b+B�}�X�I�oT>!���jV��2�$0%�9���&*V�4�ŗ�9�"=�����DA�+~m�q��oj�.ʪH�����L+�т�Aǩ@K�����mm(�O�����'�1O���x(���^JabY�`׈&�zC��1W!����=X\�rVo֣Ma��'rў�S��I1AfH�B@�@�&���H��&5ը *ڴ�?a����f�"���O�7��3��]���|��X�,s#|cs˒�+��H�4���F�y�S���i�"ዱ�:v�����8@ {�4T^^�Y��ʸ!�d�r���So�?7���%�J8jD���ikW�Fu��ƤQ��?������ĝx���(Tz�gN(9�5�"���yb���u��D�Al��+i,E�Q�&�(O@�Ez�O�F�=�����Ȗ5�8�	
"I���D�O�a��'��o���$�O4�d�O�8���?Iڴ-�\K�A��%Ӕ�Ǒi�JL��I�O�����)]ֲ��d��_���DR6V��Cף\��$`4ĕ�to��Z�\R"1@�I�=sc�@4P?#=!4�T>��;�+L�n� �Rt#y}b�~y�	�D{RP� ���,����A<=.�� D�T���#|�B��1y7����I�Q����Sȟ��'����	@Z�X����l�~�R�.� ���h��'x��'��L�@P"�'���@6�4 �#�->�Tآ�.ZO�^�&�[�X��q��5*�l���m�XD��N�=K$����O9uX8�����2��%�6�ߡKv4��䜦2����!h�t|���.FOЄP��%%�(���#����6������w�0��-�B�<1U#��l&��`����B�L0pk
���l����|�'�I�^7M�O����~*T+�`2b�{�$�+?��'W�B��i��'B��'��	K׎�vW�I4��3?�<�T?�ʑ+߉!a����	�p*eA��.�L�u�u� �����ԙ��S(wQ%��S��`Ȣ����j#=��(�������(t}�y���5�쵂D��n�!�Ċ�1\���-Dr�JaP��O<�|r�:}R.��	� 6��Z��`��1q��E's���n��t�	`��#���'ћV�ܜx��,���	)a
�u{r�/z���$�eӮ� �� Ro�������)�s�@]($
^�
H̳�J��d:x�Ѿiq
�@K���J�J��U�c�8���RB�
F��] ��W_H�H`D@��5r��O�9$�"~nZ	�n�0K�
��E�fţ�`C�	,'���񣌮�J��c�E�K&�<�F�i>�lZ i���Ј�0\u�&�^�X���?i���+&��|X��?����?���� ��wD��!����bPгE�>��,c��M��dR
~��EG^�|`�3�tL��c��� �2�Y�G0W�Q�G��͉�FU�� �����	�~�ź�(;G�����֔[t�F]�)�I\؞��3�D����/�2Ȇ�Z�!%D�8�J�6[ȴ��1�Ė�HvO�U����m�	y�4[%��\˲�C�
�=W0E56��-C䟰���D���/�(h����ϧfZ��"��o���R��Tɠ�1 ���%2
�H�ƙ�4 �F��OtI%w��PX��A:A~Tcu��ОBŲ�#��&0�U��+�
 B
��WL�< �����O̅A�܎6���s�
��1�Bo�&�y"+A,ö�������Er�ǂ�y�w",��qE��$��C١�~��h��O<)+�"_Ѧ���ҟ8�O�-��"��/���.щ��� �n�3V ��d�O��$�U�>9��?�����
M��0��Qc��*"5�h�M��F�~@Ez��G�>�(Ie(쬑�� �j[��߷=O��P�`����`�/?�����o�O�D��OW�kC�Z�bK����q к�y�����Is��,�fHI��p>a֚>a�m�g.P�(��r<
��#��e?	��An)�f�'�Y>�kG�͟ �I��#��V�T�]h�Y�-Dh$)0�>Z��iƮ�_�|�� b
�F2\�vk�?1�|�1#�橫Qa��86�¥Q1_01m�BY�,s�͆ev2���B?65"I�d��/iz�avÅ�\c��� U�)/�h#լ&I��@"�4A9��	���S��MC�Ə�Z��@�H�P]3�GU�<	�f�Ow�1Kf����!��Oi��?� �i>�mڳ^Zm�A)R�}�^��D�6|�p=#���?�Rk)Q�0U���?����?qT������� 
(��]�Gw�9�'�V�,��}8��y0"U��C��1�8��r�'g��2�FЀe�6�H!�\�W4��qD@0JơȅM��>Qz��N���(�	 v�y�C�}� L�3픨g�6��OL@賯�O.�nڴ��Y� �	f}be�(,��a��З
vQ�/E�y"�S1�M�dfN> ���%�pF5������dz�Q����4ξA����6y2U�X9<��$�O�d�O� �A�O��$|>eK���;tD])�oK90J���J����Yt�$��|��܆%�`$��h�6��d$bU#Sd}�S+�y�,��i-uE��㉬BV����5' �3���X木����<5pi#�'��u�e*ƕf�J	�B_3�`���'�n5B��7z��� ��1]Lu��':@6M)�d��^=T��'��^?B�a�;���� 	�c�v�a��!6(nt����?9�n�J�[ФH7-� S2V��'fJ����� |��ؒ%�|z�iDzrhϪ�����Θ-q��Ȳ�*2J�������,<��9�鉙~���O�D�O��'r��ǥ�<Nޢp�׌�IZ~1!��'L�O?�$ҙ8̼x��2c|Q��]/#=��hO�W]��A
]�0Esq�X�pQPxk��Y*7��Ċ)�B�o��t�IY�ԀD����'I�"�9z�,Lj��@#q�)*�cǱ ��KΤԠ%��'���M�(�.^�C� �_|��2������CQ�f���A�kh<ѢT-�5/Z"|�1-��aP�
5q�����-���o=b�D(�)��U�@�I�� �8w�5���c	-D�#�)#3���)�a�6l��/*����S�A�D�'�f�
W���t�⑬��?)�^]Ɓ� k��?���?a��u���O�.�� �"A�
>a]6qY6��4�R<��&$�d�W�S��a(���-ExR�ǖNH�M����Q����ԇ>J>�����9��y���Fb�aۯ�(�)���u����(O��3�K�|1�����Y8M�й��]���q��O�m��I.5�`���T8L9�MY��C�ɛ69�E��Z#��s�	5B��d�i>�$��;v�C슽ړ	�H1p!s%��=�`����,�I��p�I
^�����џ�'����������Gu����*M�����H��Ę��Ne�(Aw�͌p�p��!�_�}}>27�W�u���z�jE:�)��a�?K ��Ad�u�'��R�/�0U��O�%zD)��7#=^-R��IC^���d�W��?�EC� �fA���T�݆�22#�t�<����oV:T�f^*}^��C�g?IuY�D�'���k|Ӻ���O��PC$u)q.�+&,fy���(����J �b�'n�*I�f��A �ۣV���%� ����wbD�A�,Ɉ�X ��F7T"=�SD�"1Θ`�F�gO��Jc�̔I� * j�Shz,�1OI8���M#��t:1��OT"}��#�4����σ�G�x��ÅY�<�Z0H�5��^:I�2�@�%�_8�1K�����.MR����OVl��e���ذN[��M����?Q(�Tч�O�dgӬ��o��')| 'S	(��H(pǊ
M��8y��ߺ:�E���0�sӲ����y< ��pz9y��i0 0�5��6D�p�C6'f|����iT|)1ϑ=d��b�
� Җ�2�4,!�)�	��S��M��o��W_.���ª'�t��%Zx�<���M�Vy�ᐣ͆�1M��Ӗk�z��?1B�i>�l�
Y�����E?}�n����k歘��?��N�ҕ���?���?Q��"��w�>�
@9`LIT��<.(��+��ȟ�HR�ʔl�xʁ�'���w�\�b���9+�����LW��q�Y'r�p�3��^��dTx˰~R�e���'�^���-N�X��A���Yl�˪O��j��'�,��D�'X�|�� .&Z��G)O;!��T1�ȉ�)՜C<=�����W�N���4��O����Z���X�X1t6H�1jM� �8�"��O����O������$�Ol�ֈ����%���馪ִ�@��Þo�<�K���]�j��)ن��Ox�j����&�v�+�؜Z�OߟI�@Q����J��I=w�i�4��9q��.�����I�l	�@��k�)���QE-B�z�i�%"O2�����!��YrkH�5v4\���'���<14CU2L��)��!ӕ*ft�J븟���4��I�a��i���'���� <h� F4i��� A�wa�	h`I���?���?�'Bԛ>�R����$6-X5fO&O�����"+A�|�51g�
uᒩ�3}<�Gy�#".�af��P�
�a`�Ί<�B%~��)��-���E$2�� tG?ʓAv�����MC��i�b\?=SLY�k�܉�F!�C���90��3�?я���'�"�HÆX9�=�+��]�	�C��ͤ�Ha���1�ܠ#��d���b���!�?������*N���$�OZ7�>+��P�C�58����+!����/ >�8�����08��m��d!���:�s�� x�������Q��'���Ӥ�i1��8A�JM6-�!{��i#C��1���h˅��s�ҡ!�:+�r�1�ɗ�dgPY[��`�:�['�'o8�O?7��k�iv ��C�XM	�V�]�!�$�9d֜����B�b���I�;qO��dx���$�i�&İ"��'/"�Ѩ��CT:����O��$B P�Pۖ��O2���O��Fĺ������+�?;2�a�H.6�6xXҌFߐ�� !RD:��K�ώ���'>���H��OھE�Ɗ��Q��-��c��4��8��7c߀��׫���N�z�bd� n��˓9��puL�_)<Y+� ˲hv@d�'���j��Y�z�-�+e�����K)g�
<�ɕ�yBi Qp�1��´�b��dC{�(�Gz�O9�'b(8�/�(?��݃�@ۋ�$y��,�'J@��3�'7��'��:?���'��I��p��x򳭑&}��DgM$��YS��$`JH�wNL�X<���TB�'���P6D�t)���"? �����u�� �Z�l���s�(0�S9:�$����\6��i��ˁn�$E�ڼ9gn�87���1J�O�d�<y������Z�jaR'�Q�e9����'B*lO!�ۍf��dN�5%4�<�FC:����ۦ]�	Ry�_0��6��O��D�~2eH�r�Y*5�D3G�b��&C�6S�LH�'	r�'"��R��@�dn�B�&	k}���e ��ܯD! �مi3SE�<������g��w�\���i���0���?�����6��ZǄŷ�J0�&�+ғb[�I�ɍ�(��L�aO�r�ڤ!T���C/���%"Ohh0���yx�d��D�D�'���'��@)'vH����_!ukiP�'2�Щp������O�ʧ}8�q����?�4 ��}�˕VF��`�Ҽ?d`� ���V�\� r�^�3�l��`�H6��(d�r ���\cA!���*���'�!��	ٴG�llz�*�Jx�!�� @Z8j�n�";�!:�($�\cǜ{Tb�A�(!A2��h�4�شa�J��ə��S��M�!i#6Ģ�z4���5�h�2B�v�<� �S<q�� !�U��bPR$�m�'}�#=ͧ�M��G
�8Y�p.�Dnn0��͏ ���'��$d4/��'���'~l�����R�\/ mh�#
=[
=�A�d�l�愝r7z���޻an�h��Y?)����Я���UB�K?�@
C��p����(B<J/H��!� ���dX?�SbMo�D�r/�<��*�>B���J"�tJFuc��	^}rgW�?�&�'���iD@�4v|���ݤh���'��iЗ���AM�l��J$oj�<��By���ԓ|��ÕO�6��j�#�Rʢ�C���DA���'�2�'(n���'��8� 8s�䖂�Z�!�%Q��|�A��=7bX�i2c
�t����+��'�AF~��B�+S\$sv��8����f���m��m�N��H���ź_5zѰQh��<K�/Gh�T����n/�	�t �"X0�("���`P "O�\jT̖�<�����EJ�N��"O>��QI>O�d�E�!G��8��O��>�6oA�`���'�S?i��	�pR���"O_�^UC�6p�&4P��?��ư�"�nFG>f�z��K����j>U�WLZ�:�
�;�PF#Vu0�n/ғUrA*�^�8����+����![�>a�$h,B�LŀJ�hE��V�{�@���O.F�Dl�,ld��sٵED���m	��y�iխ(v�����q�
�&���p>�Ǜ>��#]��T��#�R�iC��0��z?!�oRQ����'��P>9�R�ҟ���֦q��2 ���UO�
M6���In�"��Lo!$��&K��y*�~c>7P�j?|l��[�x�(��95��&	��_5bxb���(%�,������6i�!r�9�HٗO�:�ڂZ��Mn����J>E�ܴ[j���A^�[$^@*�ᆺv�V-�������c
	3��r�D7a�D�Ey"�+�S��*T;W��(�HM�ơ�H�d��O�jsѥB��D�O����OhI���?��'�t��dhǕk���E���608@m�|�f�u�k2�y!3�~
F�	
1�J��ݫQ|\ q����n8P���t��@�}g�좓
�~B6h�1>Bb820�<���4�a�]^r\M ��	S}B��?���'5B�.Fôrp�Y�L0�(��VQ�<��bǠX3�	�lz�1�.Ѽ_�@щ�4��Oz�@���cy��J�CߗN��lQ
vɜ�E��O����O��D^<y����O��ӈA�,��xӶ �FT�|ό���,
(n�B�z��'�r5ۮO�@A�ɗ[�͓���K�f�B��'��͈��#!(<9��ܫN���N��a�8D����6����ʚ�p �}��"0D��JtJޚmDP����G���ꯟ���}�ՙ;4�7M�O.�ĺ~��i��j�uᐃ��;�F����7j�|x�v�'3R�'���5�'1O�S�D�H�"Ɣ ��5Q�6=�#=�c)M{�π ���vb�/G�R h֭�&������fVJ�$c�O�l�JA�D�#ˈm�u���GndAs�'���C���?�ƽHR�,F8A�iO�!��#��M?Jʨ�ؓm ,C��^A�V�i���'�哽Hk�L�IҟpoQl�T��*$��T���ᑵ�F�� LPb䏿p�(K���mx��K��#���&>���[Se΁a���6%��)�A�C���*?c��Q&��w�P�!dc`��5f/�-#P��m��O�B)�u�M��e�[K>E��4�2ѥ�>f���s�'[�S����ȓrJ|2b!�^=��g�J�<~Fy28��|�۴/���Wc�0k�=+T̉k)е���'R�~�H�ц�'�R�'�R*lݍ�i��H��U�G�V��cL�m�$3�U� �wĊsQT�:��5,O��O#m��I�.�0[�h�U�t���@d�T}��(,O��(U��@ �)�%ӁF0�p�]�"!��Or���I�sɬ�H-��#��ەf�,:�C䉁oP0�$�-t*4�U�G�Af,���"|B3DC�nP��e�7Y�>����(�HpK&�3�?����?	��z�d���?i�O���tNR�6<���j�Yͬ��e�S&o���ղiE�}���-n�0�G~�h�h-�e(�H_�.�d��v�˟l�As��^}0��YN�PCC>u�bqCsτ�㞼�g��O� �2�D�K�$�� s�����_��y"�H�~�Y�+_�:����y�T�K������8K�d��𣘾�~bA`��Oz������9�I���O44��l�>&\�U@�6zt @�"� ���O����5h� ��
�'|�S��HԞ3���]�|�yS����HOAgl�N�Ƹ*��H'i�R�y W?�)c���2P��O�6
|�#(=ғB�Ԅ����(��쩥X�v3ڙFJI�����"O�{'Ǒ�t(�k�Ȟ���q�'� �'k�0�f�X7~HdB.�br���'�]�B{Ӕ�$�O��'<�[��?yشV�QA��?2D����a��th��R
JE"�b�Z���*�`h~������5v�}[��ɒ�Y� tٻ���M�"�ҡ#7���У�6LV�ѫ��37�0E��E.
o���5�b��B�4��/L=9�l�P�E��MkC�ٟt�O>E��4T$RIұG�2k�Č+4�T<-�y�����I�bA3#H�" NH�|�0 Gy2�<��|Jݴ�*l+ N϶ry�m��R+F�nXZ��'��$JHa����'�"�'X��r�����qP�!ݺ%F,T�w�_�^a���V�<p4��DO,}���QGoX?]����OF�B�큐�9r6�¬t��=H"�I�}���Ѫ�^| ���k����V��9�3gR/g��I
Mٺ�Ȃdې��	�e�	\��'߆�̓�p=��+,܎i��)ɚ�a���t�<Q�N� ����7��;l��3�J
u�"=ͧ��Ne��ڷȈ�n��<��:`��Y�b��mL�����?����?	�J���?Y�������"�*��mLƸ�3��[�6�¥鈷#�$�GK�$s�|D��#?�BV�^p��e= &ra`��TB<Ƅ���Y^x���z���e�Ԧ	���Ƴ5�"�%���*�O�6�٠~.��@�@�[���5+KN!�$C�n�!-Cı*˗N�b ���HO,�-�c���i�s�>4���Op�o�P�I<i����4�?A���I���HE#Eh�4�8̂�A)z����)���d����#;�4�W�נ{�8Q�gZ%p`�i�O������lئM�D�2m�0��H"jc��I�[�朳��I�� ��	?�,C ��#X���U莇1Y��3����=���N>	��������	��xW��
㎍,�9�$*^�!򄑒]~�h��3�N̙�蘿J��hO�C��)�d�;���C��`��'G�wC��FC�n�����\�$DA�(���'$��f�x~��kD,I��pZT̄!ijVQ�Ǜ`��P�tn��E�܌�e@���$���m�E�7YUPh����r�=���i���e�NqZ0�&[V�qJ�-�
�u���o���eɧ e�pEEԩ.[L�1e$��%��Ox�nڬ�Ms������\=?v���Z G�&��2�U�~�'�a}R�E-v��\�0C���3� N��(O�Ez"�O/���1i�1[T/ο%{�̺��՗Cn�8�����hO�Sj��*��O�o?V�0q%�#�B�	'�� �0��vnAm�v�b�����4��I�Ub&ՒWK"1	Tz��X�/DrB� _�p�q��M���)�#Y��C�I�N�0��`
�t ��+_�I C�(f��k nV2���k�/oC�Ɏ=hRY����-m����*?\B��#	�`8����UIt�� M�g9bB�)� *͘��X�r�S6��@}f�0�"O���#��8��%Td���C"O�u�N?��8!����C2�A	A"Oz��n��~�=@�"�,���"O��p�ζ
7�u�#ϳw��!2"O
`@��X�D�]D� ���"O8�v�99{��2&B?�t�"Orp�M�ZT�1����jiu"O�����C"��Yf��3/����"O> jHϫ9����R��	N=c"O�D���ܥX^J��w����,+"OT��0���,���#X�Mv�1;�"O�C�@�\�Zh #�W�Yh�qyr"OB��@� �.�����*��~�^�B"O<�� �}N�@4H��	��<0'����(��L�
�)�#�$<�Ӏ�$N�=��a�!*�Ɲ�aꙔy�0g�_���x@=�T�!��R1+�R�:���.| �č�_��]�*��D�t���^	@�؜�U��p�FCd�������|�&�!�˙�9CD<ba[{��\��nC'r�Q�Ǭ)�H�S���h
 l�R' �#pܲ,T�6>ؘ�栂�.v�:a���?�C�M)j���p��l����c�6hѴ���6#>�4�/=�܉l؇,��5�@�٧K��͹C'X����+2�#��\�8B�a��EH�}� �ӡ��0��M����C�k��`0�ƕ<��x��_�W�B��iR�qg�4��)ke���i��@ppƔ�y��@�^�S�,D�֩�1�vP�C���	M U�aN�&@�& #�*'��ܘL��I���(J�0(�B�4*��Q�ԀB�R�r���0*�}ۂ����V�B�L�21�7$�E�b���Z)h��U(H�H:�³a8m2u�u/�y���	��S*=ay��^#�@�ɣ�H�oG���P@G�V�J1R�G���B��v�(bT"U�#Tp�y�+��jN���P�ǦV�P"U�������g;�ђ�e����5{1F�~�Q����*U�c2���$�F���!cm>}�L�f�6<$c�OX5^G*@��k����:�#C0c��m��ă6H�� ��n?��[,&�]��� �N�v7M�d(6�1,�S���r�|��e-:�@�LU�����eX�}��y"���Ph5)�+[�m���H�b$�(h��>)���(�N�/iII1dgH6 "�ډ�R�愑G~�PC�R~�'�(�y�P1{TR!�&W�gX��9�,B�V�ۗEգl~	Q&e�b�2�!U��2|YRj!�V`Q��Q�,B�SI�e#1�؉$l���I�gG�]���4j��`��I_�'�(�í&���� �C�?s@����[�1t��b��5�<|��Ջ^0��[��"q�L6� H�gU^7��s��*f�p����f�l*��ǯ5FU"�CC'V� {戀&��'�4Cf�A�df�
�D��p90pr,��c�@ꆆB�$/ة3 ����,Zq	�-hd0� "�]:�Ԩ����#��ܒ&ƃ�&*́{�(̘���	�ka8��先� q����� ��\�\_��x�"��j��xq�`�̵��
( Q�A���xv)�(ZR������Y$X�㒢�
��`O�"xn���b�=*&Z�8��
�~�G�X\#RݳR"�	������<��	ԩ^�Lu
��K���Hè� j�B���t�H�#o:dAcĭ�+T�,���`��?������5E�*�je�]�$����2�65�q�t�?�ȝ1")K�)VzIpc�[�LЎ���
"��I7-��=K#��7N������z+�U�E+�"kr��G��8u���W��X�4xRRf��_z3Gظ"�}���'$hr���'�?w�Ы�P�x��p��^�.Q��Jե
�~!��7a9?��
�z�T(2�C0�:���O��\��O�����P�
4�@dauEȾ;�8�ٰ*�6��H#��VW����I�	�K�?�W�(,M���t�Vo���9���[�a�� ((x0M�8�����:b�2����)�9�!�%!:PZ�oL�=�D�r6�B�.*\$KPF�{v=p�#�gm:t��4cиإ@h�r�,��Z^�p�@L�[�:�:`$F��M3a�
�~��8S�h�	6��K% ��rȲf�TU�0C�<T�%{����{��0S�`����?S�1 J,]�U1q 6|��0�
�C^X�!ە �m�� H�K�|S4%�,^�I!P�$᢭іU�bY��T�3.���S��.s̎�[ck� a�Dah�=?��
�LX�7��	 f
�2(�� ίqɄ�[�^f�PuPsy��) �Z8�6+Ҵ�Z��� ����'�D`R��(}��G�,L�S~��Q5�B	
�й�㭓�0��egh�U�&��P��<CJt��5)�l	�ޭ�#'0����Q�$���)����}��Mx�薧| 0a(C�2Kb�w(�A�z]�g���?ͧ|��Q8$��$z&Ih3��0Md�Vg/����@�G��@��F� j~���!�Y.>��X�O$\o���'�$������C��`���΁�M��kr�4(q���z�rD����1����5����J�${�6$� �Gp�:$c�^�y�|L��1�b�yu���^Й C��
M%���̰V	 4ѵ@�S4�`D�Y��(+�@\
�	�C�$���@� b�yeǕ�i4����k�`�B��T|Rݳ6ᓊe����vǮVo�uHՇT�o �Xf/ȸh�d�J�F�W%��!T�H_T����@  Xp�b\F�T�e�>�h�9:����k�3VV�A*��y4�0
��! �J�&ިe��Aݻ*�8(��l���D1B%mȅ�B�b�)CP' >,V�x��	Z�pⰜ�p����!@+i�fuk��ǔ!M��B#d�O ����6�r\�$�>90����y��
%�v�)2�D)	bMX���UJ���B]R�|[c�����u1u�T�(�Mu,�51ov}0qIPX��@\�T�L�6O��x�T�uY�Y���/T�Е�O���R�ȣB0i�B$�/&�R�
��^8(˔����/I�
򬄨2��5A�đc4���
Ev�2�ɑLX� IJ)fÉ�|�B\17�̌H>9m��Ɇ	)��X�Tb~��åV Y��A�GA�y?�kE��=8Wv%��${p��cX1PkjԳs��"_��mJ0��4~0�!#��هDJ�{�J��V7h�.tƕr���@L�sO<!�@H�	���.��:�l��D�P�4���^�t��2�z�����ϝ� ��9@w�ʁ)&��'h�*��=H2���s� ز��z���a�܂%�� ��6�p8aE�Qw΄�� �ӛ��$��� ���Sنp�@�$i��8b�ߊ!���9�� "�	!&:� ��{qē-h+N-�S#8BGh,a�I�M*�V"�;<֐3td�T���;�Ē�k-F!�3�:FOxYe:OF\��M�=$�kWB�Z�kEÄ�{ݐV[��܅(B��ğ� �%�#�Z$�N܊'p01nUQ�a�v�� e�`�6#@�W˲�;�%C6i��Jf��6o6�*��85S&D�n�a�$�sl�h���Fy�]�T�˗d��5���Ec�Qʆ��Lʢ@1��� {?��xDfۧjt�I�d��d��1�Gc�Co�yږ�N�1 �AH :��r��4C\h�u�Y6��K��Ȱ�g$(y�[ T�Q�戊��s�+v�1��(f��}�s�X0N21��G�j��*�M��9|�Qc-t�-A&�(f��A���yӈL*҅�}�$4���^oB�Y��i7W� ˧�2T�Q��$'+��@u`K�~�4�A�_�jH�y�b)�5Q�$�Oäa�$8ӋD�aRM�fd�����d�@3�D$eFmÖ�~����6�Xl2���5jC|��l����οG~�	0�őDB8Q.�k���ST��!�q�&�0���WHO��6͑Z�����";sz��%Z C7>٢������k�gӸ6�M���suNC�4�J��Q�?}�}a��c��[i�$���*6��٣ 	���
���fH�M�6���
�Ұan (]m�4���6��������������D��D�	#�(�B����a(EJ��T)��>Ic��>����$��Q"�ԠA���19���)�SVeR�M�~�&��$
2ذ 'g߆|�W-R�M�X�p� �8]N�I�k��a:��ƛa�)�JHi>N��d#�q��#�d2X� ��#�I<t-H� �AMH]ӥH l2T����t� �Kd�7R��f��/&�*�4�Й_�Zh�wD�=R���:����N���ȅxK��%�Y�yH�i٣6���p�ɖ��$J"<�L���LL�ps�
��<��,T*$����'5��� h� 9�\�:�a�ML�`c�����LC	?E�Qb2��>Z�4h���aW&��$�妱�w���*<��ql
�y�'(:��l�q�`j�$��0~j@��ߧjVB��f$�H��
gG$g��M�Ve��lHvTJ���-3t~p&*ޥm_T݀��&F�IVn��-3����ߦ_,l� Teťc����"�8�J
J��ٹ奆0;�jыd�D�����l]�4�c��X�Q�;'Θ7PXؙ'O�e3u�:t�}@���&�#v��5T頁W�� ^D�1N¿s�8�E�����h@�[F8��X��i�)���l9E��p���Ŏߕ���(�ȗ]L,/Ia���"&�@	 �eT�
F���-i��zЄRZ�ɰč�b	����(L9xa�N��3���<4��ɀ��)���E��FՌ	)ɟ�kʄB��?_y��Y�6��Ő�!L����a�Eӌ�ߎå�ޞ>&3�B\�L��a��!�$���#���1/­��7Y\<r� = *�n�0�P��A�_���:�)\]��-����%6�L�u�	,7�ҡ�e읃K�`AC�#�\����i|�Cg�ӹ]ݐ��#��%�.���}�y ޼CZ���H�H��\��aZ�����'�έ�D��=�揟�(��hjGD��sl(���E^�pd��f-�VϺ��$U�V��xG�.h��5Su�ʓDJ騱垌pxho넝2VE%�f��OM�Zr>aq!��`Ԃ!��3W�2����� �Mǯ�,;�,�M��b�+�ɸ%cG�$'I|��D%�M�\1�4K�Hһn�� �7+	4P����Ճ�B�0���/���dC��LY;�{��9j��0ؗ�Wx��b��;&XR����M�4D;% G�*flY��T�`�N���]>��uA�
P��}kYw�0|S�²	≂�"�)��lH�'>8���*&`x� �8ʖ,�B°���QB�>A����Qp@�Ҿ:��aq��������%��qI<�룬�4�4�I/^f@PQ�R�
0oK�t�@dL��7-��s����z�����R@^e�2˗E�i�g*�	�f�juD����[�Q6`dh��%�$I��e"
��i\�f���w��tZ����C�^��C �-~q∙G�,4$��E�]�n�����y@��Rカ\������)Z�u��.T�cX�!����8|I�e&=�V�QV%� Ld�㧄�n�OZ�2A��l$�ХJl��3��/���VrӼdy�z�8�s%B�z�:\
�K#��]��`��$d�G냠>;vH��t��tN�**�ܻ�ap�t`���2I�֥)�E�|��e�.�Sc�K�-�lm��E�z*
��$�T��ɤ���oaR�WB��:J���O*���� �O�p� �E71*�ʒ�$;�`a��5�f��P�((!��a��*�X�PRFd��d.�>���Y.<�=0EE�Jt�]谊�m"1�`�A�Q�Md�Y%˪[�0)�'-��pú�F������u2�'D.�r�k͡`@�����W�.$���J�U��}X ��;@~�!T�H=�2�H��_��ԭ�#��jv�	,d6����և�y"��d2ԍ�2�S�NMjy�
çw��db���}0�[�ʧE�ƄAw�M$����g��:t�lbN�v��b>yJD��ټ�̉%h�-�Т��q�p�-�p��	�;��Q�A�ԶRs�iI{I6��K>yr��s=�\�S���:�%�P�D?.x��c�7:_� ��.��H����	q:�x�<��q��H J�<���R�f�Ys����Y5�%��4S�b�Q+Odt��d5h�X���̾H�r4��L���4G\;�� !�	��]!���䡟9Jr��;g	8vqO�bt�
+Iyx���)2c����a?��C<S�L�q�h�
�bЅT%>:�iT3��\ɘw�  2��Zk���W$�78źt�b_<��g�P &����W�]'V�(�A�	�#8��
�x��E25L¾r����%����w���*���x�J�=��P�3 �@P�fP8��OPe��� 6��Y怄�?��r*8�T��'ZnX�P �&zi�S孃�L�,�rE��H��F�zX���d	Ws0`�:C
��8��|r�i�OrMW�V/7��AÃ��&E�4��D��p8r�j�*޴=ˮPD)�K�zѹ��;5�x#g �9t�� ��ːx�CH��� ��-Q�q*����L��C<���q�̐_��	�b��e(�*�����џu#���ф�y7G �v3�!ѕ`K	h�X�Y� ���>I�ڞ4y gJP����J�htv$㦦3^�� ���=��)�gưkg���*�����ꝃjs�'�Bar�F�;�\l�a��c��L<Ѱ�� �"7��'R��4��)dĚf�%s$ iJ%�I�y�@)��3|��V
�	M��7���&.�An�d��˓D\��#�V+��cOѩՐ8Z`��<5�:B�>0����I� LL��c�!P&��;��Q�Ӝ bd�M&����	�]�^��m��FqY�D"�O�$`b�]�r�h(
�i� .t��r!L 1^�9G!T��$����-� �C�r�l$*��N!-p�=�¡�8N��-F�:�Z�Gi�QT�U"GE�+�J#?��"��H="��B�8(M�&*^'���ݙ��,�Ʀں k��c�C�=�ءAȃma��KR�9#1���M����f�[8%g�)� �Qp�/�4Ǡvf�����:�Q��!F�ر7>=(t���.(�gL�gؒ�IC�N��0��0{��H�gE!Cj�$���+8n)��imEshP�8@|�1S
Y�|mFRB�du��c�L�94�qzff��y-��hv'�!:c���cS��C�/F�?g�Y����"#�JH��l +/Ӡ)����P8��ʑ����8�
�-�WI1�p1�7�9�f�i�(#L�$�(&d�c�ǘQ�xY��2�~7ͅ�t<�`�
-!N�Z↓�q�dYa��Z��Ah���09����<aЄQ08��7Mt�b��O�\��m8@$��8���	7�i]����?�F(�ץ�e=�����7���sJD|\p(F�\�(Z��H#���A�"�<*?�)Of��5Ë�6$К�NX&C��\�SV�^1�`01���YR�*8�`Ѯ���'^�����V
�za�e�1���C��˧Y(x㐪�Y�8���2��T��!B7��OP��p�<�4��2��m�aNM�a�6�c!�C�,@�c��a�B�(H��!����� (��S�<.Y���_�f�4%�#����\D�D�48
ў,�g,�*N��T� ��&���M0aZ�ό?��,Z��H�*� �~e��Յ+UJ<]	d���?�8����PY�b%�RE��#� 1c6� ��BJ�wb\`��U�~��	3�Ȥ�f��
��,Ɩ#z@`ySn��o�X����b�d��Aʛ�r��ȿ)��%he���Qqo�1/И̃�i\T��9aK��`-����>+��1�'�� ��I�>PgJ\!�R�op$�h��	2l���C���&f8����	R��)ߨ1#�'F�M��R�q
t+8�V�k���@?&�{��2F��)��OD>j֙���|�U�7H��{�%h��,ﰽ�W)�/�|�W!܀3�<��a����	� e�ml�6�>U��C J�(P�Fb3��e0�B_�_D��`B4l&ў���,+e��'�x��Ƞ-�a�1���(S��E�F�
2G"pN<��-̔"o�x��L\� ���#%�P2�jb�H���K`����]���èq��sWH����dJ��v왧/"?{�1����iݲ4� 
Ɯ~��s�>� c&F%f��͠�f��`h�s'�R�4ltDZ�ݍkj�L�A&�=s�:�SF�%g���3}c�c_\�"����Y��|u�xb&�Q���۠�Er�Y�o<�)	�&��'x
xp(6:���5�H�,`�%���@��BA�s�>[����"F?�y �(f�UyU� ZD=iEa�+����ѦQx�ȵ!U�R,�R�O�8����+!�(@H�B�1U;R����M(G�F�`!o�2q��Yt���7�QZe��(��y���.�&���,��2�O���̰e��l5nĦO�E�!k��N�`̐�#�'w>���F���Wf[�'0r!�'�� �ʹGr�D�G:�@Z����O�~�b���Rm����ߩ��#�W�w��:Ŗ>Q�>9���H�bMY�s���8wF`�,���U�.ޚMoXqa*��|2'/8}��A�)
v�S(٥E���QJ�y�@�<��Y��ɃyP���,Գ.PV��0���j9��f��]�H%�r��T`SP���p<�qȚ�ZФ��SG��x���ҡJTX�L���nc�Mb0�
(Tx�����H	�u
N�es���z�E�ēS�� ��=p�.�h��y�8�<a��x�>#u	��:�����b��o�8���ڱz���C®�y��ݓc��<�S�UY�S3m����5)��J3[:��O?�?ҸdФ˖>1Yc��6��C䉨:T���iÙ'�>�zP�N�|�C��?4�T}q��N�<�,5�r�Y, vC�

���]$�����Q�B�I�-� �qHΛ4��(�0�U	t�C�I�s��e�G)�~��8F"� �C䉒.(��f�+�zX{6M�0 G,C䉓<H|� ��C ��X�iÝ46�C䉄UZ�i�"C2^v��� کwB�C�	?`�A3�
�l��y���ZhC�ɟ5�꘩b雖c�ܡ@T�ٲEfC�	�9�(��*1�؉� �U�YVC�:�i��F\uL@d-!|(���"O�qr-ѧ!�
0c�D��Cv���"O����V�U����	�W3�Ay�"O�̀�����m��&�P8=��"ONC�@Z-V�ŲFD� j�(�"O�����I'oJ�`h�a��a��<�D"O�XÂ),r`�e���Ap"O )�+��HX�c3�j�T�9t"OB]zG�L�B:�y稗=]�Ը��"OP��J$M-)��"J����"O�Y�`ߢ^�Π��g�,-m����"OJ7F^�a�y��H@�;o�E��"Oh���ODP1�A��"KL�0�"O�xc�"F�P�T�2'��v�����K�!'|rE�$�O.8K1��gԨ1	1ɗ�>	�!9�"O~�V��G�n8�!AќEx�"O� �B��T �E�W�["�0|�W"Ot%	CnR1RN14

��|�5"Ol��'M�7��H��)ɭ6�����"O�ъ"52ʂ<C�H��s�=��"O^�m�"U���PT�	 b+~@��"O�%��K�nFn�����vfA�b"Opq��Z�*�+%�0x��� �"O���'ҾKW�p����+�Lu�q"O��Wꊅ9��᦯<�*DR3"O���a�F�MN����ׁ&�r��"O�u��E��ԁ�M�{�8���"O��ǍN3��SUj�V�<}9"O ��QA���x�Y��	-���@"O>г���+2�Y�������YR"O�UA!�S&��ӕ�՛`B�"O���e�/	��m����g�He��"O,�ȗ/Y:Oڔ�����8�I��"O�(��P�,��m �
ȷ5~Jh��"O��j�F#�"3i�nr�Ѳ�"O�TR� jH ����ƾ_[�9X�"O��)F"Ͳ���R"I����"O�� 1BT;���D�}4� �""O����U�1 !�G�8�l!"O���#H���Z���#b2R���"O Lp#��{PI:.�+����"O8��E� u`�����F�*�,��"O�$���M��A�R��=��[�"O�-P0�ֹ9�t2b(D�!��]��"O�YI���ՈY�GҀS:��v"O*U+�[F�J��q%ޡDRe�w"OrP"g+S�A4�0vcLR��"O&h�#JߞY�12��X�`�#"Oj�i��W����#���!�x2�\��4��K^u����<C�|�w�E#���Q�I�9�pY�@̾s0l���?Kи�ؗK�E����3Ӧ?���� �',�q����E�v-[��#G�
�Ja	X�gǒ�H1p`��@�dp����%8�,X���n�J�P`�E㐴gab����ʍ,n����ߕ�퍟^y� I�+ȉ	Q8�iF�E�1�^��c�D����K�f��b>���S�&dڕ��ݾ) �q3E��Bt�@$��B�����6�
<�1$�XB
X�g(1:��H�a��0jp�jBDרk�N��^�T\V�ߺ��̪�`�K�m��P��iDHϘ�����e0�� �@G�R^���`�����H���X�FP��U��
�Lқ4^�́n�����R+ ���) ���&V���%È>^����FH�8(���+�2��䘒l��A ��MF!��gƣt��"dѡY�(�`L H?��倢��G��-�� �OQ���S��ko�H�w/��W��p�ID�x����w��TX5�?1�,u��Α p�H��FOC�q�����Z���	�9���?�q  rd0���iD6rZ�C�>�́����>����~x|�q�"�n{DM@����9 Ec"�	mJiC�C2��R$�P���H�tѶ8&,��{��D`$�7ОIe[����B�����Δo^, �.z��[^�Y /�t�T��h���ژ����5$����C�D�Hϖy��L��Xi���ܰ\�6Q�w��;d���.��z�,��a8� ��D�;`#Rm���v�ڽ��E]:�4�2*Ŧ1i`)k��͛IT��J� ��l���)Z�OHF���)5,9��]'	p���C�9�����weL���)�T�ڠ��K�\��V�\(�bAH��:��A��Je\��b)V�! �'2��P(g"�#�\�Mȍi<��
F"G`�tz4�8�(�nM�E/H�8 w����QuY�]R�(T�b�P���6�?A�h��pa����|޸l �O�)�HK��X9!<Q��O�@���K3e��PZa	 �C�z����>��� ��PS	:vvyk�d��<As�A��bc_	28!����vZ�I2/K�N�p�'�
/�##M��$����P7�D��d{���W;�q�����>}R�M�"�W({��p��#>��"g!�'j�I��$ԟ,"���蘾qQ�LB�S,����&*(��C8l8ڣ>�]6c��uy�C�<���f���d12�M�GO0%�'i���B�(��e�8��]� &� E�L�Q�+R���	dj0� ����:"$yTn��k��&TY��QS��h�hQ��@)�큇T�2�b���*pAH?���s
�0����69sd	��G��*x�'���&G� ��a�u��E[� �2 ��}�@�Q�ή(d����0h�b�#�:qv�̊B�����z�7#:?���l}��Y�	��!��'�JO8��"o�$b��RĎ�o�|Cd+M�/а�E��8e����5�E��|� �u�ax
� �`���x�l8te�"�`�;��>�t��{�4��sf�"Z�`0L����x��_(
r8Y�N�#d�Z��E.�'Y��B�I��U�}���X�Q2MR2����l9E���T���iHė�~�A��D�r�> ��$�DQ� 1�� e��'	�mCf &J��cQf�' ИE�|��:Q�Q�*M�;ㄹA4�[�B�¬�	?+�Ż7�O��|"��A_�I�l�|�c��4�N�@
�"����B�P��XJ7�1	$`�(� �?ӧ�@� Yy3-�7t�,l@�cC,N�T p �dS	T�>�2jI��G��5��� �2!��̑9a�D`r�Obd�|jP�A���A��<�����c[�0#F�I*^�V����#�I�L!9��"����aau���e˲X`�	34��Qs�\��MtӰm[!��s%b^�k��� ߟ�ԟ�I��@���$s*��Z�'?�'fTuK1�3�n��k�S��}�`��W�KU��9�	~Ֆq��ˁ�B'�v��?~G8�!��O�(p�|Re	<�I-^��;C��}��y�sAU4y�4� dM\�w<���A�8�TD��@2�'}�$�`�M��,>蹫��g����#H <Fİy��.�DD��>�]7gH+�J�m�i�����2�ƀ�F�4X��J�T?���Y�D�4z��p2\�y���$��ч	u���SrG�Ȁpk��W��q`%�==����E����2�����[Ц@K��� �i�U��	��<���eC�� ��a����>IІ�o��(c��_��yPo���I!>�w��0�QawE�[��S�z���A��r_��Y�M��@⊆�U`]�a�_�u��5+�d.h�Z��e�d���O���`� �X-	���5��f�*H��CV�ŲɰHX"N�d����d�3`��OqR%ͻ!��Ia�M���J�^���>��A���M~&�`�3�	GJ�q�Rd���գ-LJ�h��ʐz�4�橍4���%���~r���,!($���r��2�Ƈ?7@�k��D�e�v�I�і��t���!m�������C�}��5�Il�ɞ)�l�3lM,)N�����~�h�j�(" yJ��	Ԏ�.�4Bv�X�>k�������AL�#`Ϝū3f;x����c���XW�
*��Il�	5#��I0�H�]��:#ϊ��X�`������:f5��ǡ��Zd��CR��z�ʌ!R�Q<�y�f�9 M�������'	\x��^(�Ҵ��Au�<]`�4o2t���N�v�z9j�憇KL�F{�;�����i윴e��HHц��C?�Eˇ�eh�ᑃ0S���c��44|I�T�IZ�x�"��"/����35����Vg�ڂ�j�F�2�[��DPf?�J>a $ӝ%\���R�K�Y8� +��H�1+x#��VY�f�V� BX�u,�}0�4$v�?q�}LԹ��,[1A6���5�عGyZ���{cI35��1�RD��~>tL�'�@pP�N�T��c���h\��d'U���[E�Vh.���)�	�{Ҩ�E.X�{�(��,��1�fGX0�i�h_<e����2���hOkL�;W;:qX'�ԍ0��x��I�B9
�ExR WA�S9��+�|s������S҅i4�|ȴ��GKў,��'!t��pi
m}�~ƀD3h��>�^�qE�z�� �cX �g�U8W��Ѻs�h���u�]���]SzL�r0�N�!�@5��VO� �b��w,!H���OL�3%��)z9�h"kȍ(w��#�(@"��I3�ne�ׯ��\����\�D�?7-I�bR!!�]A�y8G��	zQ�쒤/Y�"�R #���10�!򡒇�f=P�ŀ��=�M��x�ě#w�¼%?�LA�,F.%�}�E%�@[�]�e�jӜ�ʡlR�o9��OQ>Y���I�;�H�!�`Ȩ'|������iu�W��92�a�$/�ȑi��_�b��9���Έ��OT� C���:i�\�J|Z��L�8�&��$/T�;�i�<�#�a\|܀q߬I�P�bêW]yr�%<3&@��K���TY���&J� �@����'B�C�I`��T0���z
8��
*T��uJ�:t��5(hx%?�LYVd(X����������<�L[Rl`���Rj:�I�թ��A\M#0�| ����/pbI9&ᅵj�8�@d��G�џ��!툤WV���|��
Dr�B�H��ٹ?�^51a�C�'p\�
E�I[)019�OËf�l�p�'�LAs���y�*�S���6q��A
��d����F2s�T*�
�-b�I�|A�H�B�ޝx>6qCw�K�~�����k��܋�k4W���gO�<�Q�,���ʹj�(Y��A�P�9���x�M�҃��*��a���.l����͕/�*8��Ղ%�4�h`�ڤs��]��Oڭ:6E2vt�`����-�d�ѣ͊�0=y���61�2����i��)PU͞�op<𡣪�1a�1��~�T49"�2r4Q���$t��4`��&���� л�Ox��	h��k�$R+vʹ�3��>Q��T��p���A�p��QDi��tUUB�b)�n'�L&�d��e�
�z�3k�0`er���]K�vѨ��Wx3�R.�1,i�x2���H�b�B��9`fܹ���23��)�p$Fd�:0�nֽ[�j��D	�?��Л���X9N����86Ԕ���O� pt�ɕ>U ,�9����R�>�1�7lOT�RbͧwF���4 C��T��� ���q/�"4�B�	=G8��A��A�И�4LY�>z��(i�O_:6q�7
�&s��>5�#� A���2#��1�~ł�+%D�8f�Ўi�l�a��9ȲA�篍�#V욲�F<�`���$�Oڣ}��z�"�Y�$к
/� a�^y�$��� ׈���%\�O�Q�U�2�� t�8��(Ok��,r��kԉ&��8s�N��R�����i�y*��V�M�U�ؙTFȭ��/\�W`�X��d=,O��YCIO�b/���ٚI0JI��2oNfY�!JNq�4��7H�T��4}����%^�ͰK��fb�h�O�Z��ܴ,|H�nO5.H8I�$�x�̾*ܐq��A�+����-�/��'�f���1Or8B�ܒ&?���f+ �Q�,�d��,k��@K8�`�tCsS���������6�� 33mQ�p���s+\���nӁVK��z��R$�| 2��5�O\Щ,�V�\B�O[GupTzv��DrPW�'7�$�0"*�B�*E�Tj��[�蒤t��'ER�{fg͂
�3�'��J3еD����r)rE3��V�"���s����'�NtaӅ1eR�b�S�J�|�sP��s.rY�9p�4�0�GG�>!:�"��aа��9��d�oX����k�\K4��9f��m�:�� �Y����8>�Ԑ:��Ɉ�:���ڿu�H��7F�˘�*������=�C!X<UH`��%�#�$ȝ��Q�F��8��iX~��@��r�Y�?�U�B�W�jZ:u�g����=���Cm��	�p�I�\��Ѻ�Q�;�0�beR%�j�'y�$��n��u�c�:G<�I��WI"&2��Yw]>A`f�աD���э�<����3D��H�g�*5êp[�%�+O�uc�'ƭ4���P7����˓�h��D6zJa  �&
��֋F�:�!�W�J��9�Ȫ
3��mޒ
�D[�cO���4���p=�'��',A���,�D��G�<c�4�*�
g�۠.?��� �Z~�<�!.~J��ȳ��M�aQ#��r�<��A��!J�X�k�y�����NS�<�B�S�?NHu�� ?�Dh��R�<�Ӂ߳gEL�Ą�v;�%����P�<s���0��Bb�W3"�lD`���L�<q 5H-�s,��f���L�<��BЧY��J���f0dyc��I�<9�A�1���R��H�\�;���H�<YfC�"&�\�����>V#Xi���y�<ق�C$
>`�"�D�&[7��s�<9������x���A&	KV�Lh�<��@�5��h�E�.�jeR�o�<��.M�NwP\x��V . ����_�<)R4^�Cj��2#�hGF�e�<13"T/|(�q�������N^�<	�)�,�֔��AU���@c#�Q�<a��M# ��Q��_�|w�8���h�<��aQ�@����t�R=}Vغ�N]�<f�U�
b����d����hj�]V�<I!Ɵ:o�a���5'ĸ|�fWT�<q�@ѓۂ�'�, l.��`�e�<��HC'9���7*��H��<���}�<q�֪Le���Q�^3$���b�]y�<1'뜛w!���%A2.���օ�P�<�ʞ �t4J0IC3֬�04��L�<��`��^cT�QF���1�u0TǔG�<��O�a��*����QD�_�<�G��M�������W�(����R�<I7$75�V )���L@��	�CCL�<��O�;F�b�"	O���]�<q�)�@܊�(��E&����RIR~�<ǮC=�p!�"	;�l#�mRr�<���o�yhwcպ?��aP��k�<�6��W��0���Q�t��%HR�<� R�wg�(�✙�a@"O8�"�'��X.h��9B"OR�G
x.pa�� A�&Y5"O:�z���70X�"R� �ġ�"O���Rb��a��J2��F8�""Ov�5�T�[�<�e�	�U,f�	!"O�ZD�߁/����E�@0!\�q"O��W�W0Z��v��9$��
�"O�b���)Q��Z7&׎	�yxf"O�MQ����l��bF4uM�0$"O*-�#��$r� lz�/c��X "O���!Tn�K�aމV:@X`�"O��0�n
�#W ��á�6�Y	�"OV(���ޒ@�z��E����ZI��"OHْ�kF��3c��d�@yC�"O��(�#L�ya5��� 9���2"O ���Es���:���[8�9H�"O�d���J+�nص	�}xd�O�<Ѧ�~�x�GL��Bvf-P�DI�<PC��T[�L�&�/5�^��.F�<�u�Ǉ|d�,
6"M+���k�<q���
��(��G�Z���'��e�<���%= B�k�H��"K)�"�AK�<��:f�a��4��؛��J�<�S �)pB��uXx��I�<aE� ��`c&)I�H,� ���D�<I�� OQ��.ۊz��[��}�<�N�EqZ����uh�Ȳvh�a�<YP�X3t�8�w��;$2l�����I�<Y2m��f�tX�6@��S@>M2 o�`�<a��؋�x�w��i��L*�JXt�<i%�A�)�\�dB~a*�F�<Av�	4a�*��<]���N�E�<Qw ҙeըX��L44:����v�<y�U��ĊWT&~| iQpF�o�<����5�6o��xQ4��j�<1��ڕ]���Cv}����C�P�<)WeЬ5��q`��ϔ@F"��Ug\u�<��)5�^���-ֵ�a(�'N{�<�f)�ek~C��ׯ6����Bc�<I����+�v`��ȗ*g�L��B#�a�<�O��s*R#i��^��QdWa�<q�j\2q ���W�S�!Y�Q���F�<��e�"W�H�AZ>]�xaY� D[�<�PB�*e����ц<�F��U�<�硒.:��ݹ7" 5mo���G�'jv#~�0b��;�l<�æB�hD5�a�k�<A�$Q;}�ܳ�G�7K ��
�Kg�<9-ˊyo!i� 4F������~�<�M_4ܰ�e�Xn����a�<!c��%V�Vy@QmA*m:�t��^�<i�d��u�BUb�';,��1L�W�<����v���yӀ$!A'TN�<i�I^Z�v��a��#g�� �M�<��ǽ5Nh<2$���L'��(W�M�<a0�L�%,^�+ ����pX��b�<��������"ˊA��hS\�<�E/"4�LC��q�nmu�QZ�<d��EbN-��\	a�Z �@EU�<Aom�$Q@҄�mAM�2B�I�<�c�*}PH6�Ԙr�l!�'��]�<��5y�P���Ү�J`���<�A�?N�誰`I�&�4٢4�f�<���W���0�1jA�Fx�bPe�<� ���)KX8�؅	�6E��C�"O���PBK���Y�G\�X0�D[�"O8�	6C]Wb�ѳ�S0"�4�e"OV�SKֶҸiR��J�I���"O윙aΘ**M+� Y�w��d`"O*��� ����Â�ǻc�Yp4"OH�c��.�x`.%I�Q��"Oa��*U���J��Z���
"O�d����Vbx��j-z�i�"O�\�`a�8FO�A���H2�B`T"O�!���D�N&��jńR�L&"OD[�$Yk���PV�L�w�|�2"O���򥓛m�n���蘸e���)"O�tȃ��W	��6HU�u��Dx2"O
��/�K�����E#��\s0"O�|Hv��	����բ�?�R-p�"O �� �P���˶�Aۊ,�c"O�eqr�_f � j��k�ʁ��"Ov��AJ�.w�F{�"����j�"OȨsq�Y4<_.Ԣb`���ʆ"O܉*��HI&v�y��րb�T�"O@dɁ�B
μEa�]�4���x2"Ovd��CW<frl��2T��b8��"O2���+��1X~�ye@�8K�X s�"O���(U����F���OA��"O�-h�o�/8XdK��{Pr0�b"O�-���M��@���H�0�"O�-�d���fz��ʄS���pU"O0����Bb^@��g�
@���f"OP��g"�<��%z�F�� �"O��(4�����M��D��U�pa�!"Ox�b��L�?�YS��#(�)"r"O*AI`ۭ;��(0�A(7�EZ"Oa��,*���Bde�z�����"O�³�/lz���#ӉRxD��W"O��n��8=���]�4��l؁"O:���e���:����ݱ\��#D�(�b�tX� i�V)�a�S� D�8� �!~�RЧُ5��2�!D���N�*a/傀nY�.��lHp�>D�Tceȱ/`2u���x���#*?D�@{�f��?TmX�
�)\��Ăc>D�TG
ߺEdp0��mh,��0D�H5%JB�L�S�6<�*� d*/D���4x�"Į�Kt�#f2D�L�7C���)�'��LF ��/D�0!D�·r70D�N���¹ʷ�/D�L��ńjWf�ҦjG%M���M/D�T�d$U�D�:fą�YT���u�,D����-D�!���PJBL����*D�T�C�05�p�� /G��9$3D�X�$��t��s�N�S�РYg)3D���G�#QL�㭞5�̳B�0D�L���~���ģ�uW@꤉.D���6�y�hP�'�� �@cR�(D�l�f/Y��{�$�/}t�A)(:D����bZ��S������ щ+D��jF�ߏiC����R�d��-5D�xQeB�r6�����'PL�c�2D�$X�%]`�=�R$�6�"�I��0D��x��?9U���P���8�j�9D�l��fX�d���CĎ 2�K	�!�_5ͨM��B�.vN%�N�0)�!�DG�a�ܐu��8Lb��;0g!�� "daV-N�#�.�cBL�K���â"Oz����B/�:�A�
:��p�"O&������@���e��|�B"O�a�ܥG?e�n�8����"O:��dOoJ�M���0r~�5�a"O6tCgj���6� &ɈfRLH�W"O�P��Ar;��C3V	x?�K2"O޸P`���K�!8��p{�"O\�sG�D�@�UJ[�m)D�X�"O>9���+���ɑ隟u!NY�"O�#�$L=/Z��#)� �&�"OZ9�!&�8#d:8a�HE���%�S"O��CU�
37��c�&#�6U""O����e�8�����Z�~�
�"O�)�� �>�hЂ�P�a�*$yq"O M�C��$E&��s�E�
Ҥ���"Oz<��	S���F%ˣ%)B���"O�$��&*ƀ��r��B@z�QS"O���v�16�(Ɋ��H����&"O� ,�%[���1�����"O�i �B�]M�����3&���"O���=~�(�d�X�^�8��`*Oz ��"I�0NhH�vm��L��'�^Z6d�0x�4�w�QR����'����,�0fб���Q�58�P	�'�z0rfL�=[��#V 1xlM	�'�A��'X�:��*F�&RѨ��	�'��T
wI^'*,�` ݋4Ү��'�d���	���
�Р�=+�'7(�iG�ؒN�eP�-Ī	����'���vʗ�nH� _H��'�J囐,��$�% �zP�<�
�'4����m���ēm�0P�
�'��9�a���AR�$�?Te��'a�u�N��W�q��<w��D�'AF��ddM�n��3a��p"����'-�i��#5p!������<I\pB�'p��+��K�?i������#n����'��!{�����ܑ����.I����'�08�� 0a��2΢�J�'t���gD�Z�N���4o��k�'7�8 �M�M��j�,(Xv4�'�����0��Hѻ"��x��'�T�J<2$�=��a���2�'`�a`�M�Ud����D&T:u��'�4� D�*xԫ8qp���'���1&	�F�	��؇g��"
�'���g	�fC����CgHA�	�'(b(�G����"Uj�[��A��'G��@#n�w˦9;��~�8��'J�P��η5hZ�2#g�6y�D-a�'d2���A��OtV��,Q. �
]��'����cؐc���:`KC|��'�Р�0Bxm���w�A3v�(x�'9ԑE�H#}nȰ��D�@�'��:�� :>Y&�*�īmY~�y�")���vAG A�\�_�V��ȓ\��&IA�Eh�gC�2bu�ȓ8�=��)a�yDOؚ9�\фȓ:��� ծ�q2���ʁ0oV�ȓa>�z��Rr��7 Rq�P��T��u��r%`TQt�
.=��	�ȓr?|u�!J��j&��x�`�&ELش�ȓ.��Ms���B��CG]"+gLl��S�? �]H�+�?\�m"�n��]��""O�P���ŵU+��fnY���"OV`�OV�c(�@D��RA�"OLL:/`�H���M.^��I�"Oj��&n�}�&��$�V O�|p�f"O4A��6�T��l
Ve��pv"OZ C�K@�3�"A�ԏTZ�M��"O ��P�װ�.�[FD�	�4ٰB"O�)0�k�B�V����_v� �"O|���1U�sGC �^r��"O �{bmU�1�fd��+�tL�('"O:Y�E�O")�v�q�hY ����g"O^̨b�:
�4M�e�<W�6�Ju"Ov0U7b*�k֖�,��"O&�9�/,"��U�c���~sx�8"O P��$;�H)�iB�]���"O��V%ɨ:ǘ�Zv�'e�x��Q"OB��B�\ 
������ /�t�RF"O&\[P��h� x�,=��9��"O�P+i,np����<���"O�4I�iÓ��2��\��"O�pX�m�c��l�B�U�_��4B�"O�`t�f��hЄ�/M��	�"O���F��^�
gN dz���"O������e-��OL����"OY�LШ�R1�凘�h,� �"O�0*���(��3G!��"(��"O�dwc� \G1!�m�		�5�G"OƘY��K�P�*����c	6�À"Ony3	��jR������=�dy1"O�-�FUV8�H�)�b�3�"OD��cdJ�~�����Җf��e�E"O.�i�!�3	����7��8� ��"ORyD΄47�4�g$��Q��y�#Y8g�JA�� ���dX��y'K;o��٘����P"S�N��y���+�D� e���x��2@��y���2��S��]��:���F�2�y��^b��ĢU�7"���Q�V��yb��DQ�!��R  5&�P���y�@�?a�tQb�`:q���Ê�yb&� ]�*�	�E� ,P���Py�&�:L��xC�!3�@��g"V|�<q�V�Xp}7k̔\:D�YBM�y�<�4B ~��Q��g�4-1Ga
r�<b�]�[�T��֠D<���G�p�<��f]r��f�
�cHh�Z�b�k��U8������p�Q�ۥ;SB�$6D���vi��z�z@��@�R�@�5D��9�Lvd-��KF�8{�@z�*'O�"=)�\�X+�u�Gc�B���ه�L�<�5�/D�q9� �FV �C�F�<�w�:)R��@-�-i�@�!$
�l�<a���'A���'��p�"��G!�h�<��b�?zV͙��W�w�dd���y�<AQ��F�Lj e� [�b��n�n�<�(�[�^ �aY��Je
�o�<�$nߌ���P�0��Ð"w�<���� Nk�hZv
�T,����|�<�PkՔO�!3"�ս{�x��WC�{�<�W�F5X���'*��T�w}��'[����.?Sg�}�ř�X�0c�'C��B��IL�:��Ҥ�=� `�'T�˥�:�f\cHƜI����� t0iwE�7}�ŀ��*�����"O��CƒJ֐3u��3~h2��5"O���*��n��C���Q5��"O2@�cA��=f�$�����_�1�"O����ƒ6$RV��cՇd1�y�"O8���A�����VYs"O�e1��G�R�R��W�rsR)�"O�5C��;�8���c�2\�C�"O�5�j�A*� ;W��#c�H��"O����L�A�����B\\�[�"O��r@��3���H��X��"O:ibt���� �"�F͉4� a�"O�y��]�1��91����X��`"OąJ��U �>I:R��L��= �*O�q�*O �5��ʞ�Nh�'0f���R��Q'W8?yX�'ѱ�n�8|f�6M�>i'�t�
�'Z`��l����X�LPc5�͓�'�D�K�%�=�|� ���T\r�9�'Ȁ�3fE�I�,�Z��=}2���O@��D�%W��p+���@��(D��}r �<Au�Ԫ=/�D��ƛ�\�����a�<atlL�x�$�Ո�:da6,�\�'a����n�4�P�%(��@,A��y���8tiP3��t)�=`Ԉ �*y�=�O��P�<ٴ�_:N<�+��^+G�<��HQ�<9	��O�&��ӍЮ#��)���L�<!Q��"h�,U@R��>_�a���I�<���M]�V��ÇR�OL�B&iV�'#axR,�l+~42��_ۨ�Q'�$��'����S)����iU�s�Bh G�W�cn��	�G��J����iWb��CS%,D��ڴpt!�d��`<����%� U	�
ԚM�yҦPp�����f����9��K|�pm�ȓ�lHK��׳	�l芄+̑)��-$��хW�ا�O�d)��G��?7��B�Q�BQ	�'t�(��bH��"`NN�i�h�3�IF��~�X� �#_
sh�AvA��p=�}bdȐXv�)`�����E�5�K��y����(�ߝ{&�Q�s���y2jY�a�č�P-¶s�h�Ƀo���ē�p>���W�FCxy�&+�6H�>����T�<q�ߖ3��!��R�nf��p�HI�<�f$��}S��A6
X;c�ȁH�CC�<���{����T�Ү^�P��3lF�<q�璅^FV��2�.$�s`�A�<���)�
����(|���e
FX<1��~��Q�c���3��d�@ ~�Ɓ��Wp�X��=5т�9�`�yX�!�ȓ-ǘx��M�\�֝��C�50�I�����X��7l�z�Q��׫?�|��z�2yH�#kz��QG
%4�<�ȓu�����]j��i�L"B趁�ȓf�[�)�{�N�v��+���ȓ_�z���:�he�L_���d��F!4� �l\�#��%�`��J�ȇȓL�������!D����NB�V�Gz�'NΜ;UIHF�f5ʶ$��c��%��'`�}�S�ͷT���C�ON' ��'��HP5eƒ#��1kv匱Ff6�
��M��{�Kۃr���G#ZdYE!�b/�y�γ3��Y� �5�~	#ӆ�(�'�h#=%?)y �9K� �6nL�^��"�5D��
�Oʬ�f<	�ϔ�f� Ћ��/D�� ֡�t�ʷ_ �3�*���V��D"Oj!� ��*`LST@�7sɨ�E"O4�`��L��ԙjZ ��"O.$y�gȑ eB�qN�6QD�k�"O04)�}�V-1F�����Od���]�� eʓ·�G�:T����:L��l}����m�6�����I�n�iQ��Py�jF�`)�+SM�Fe8���|�<	7�߆�Re�eoF�mPD��"F�Dx�l�'�dzA�R�_r�e8��ۦjF��*�'��:�뀠EGhc���%h_�ݨ��(�S�ԭƱ���eNխ+��*�d���y�G߬5v�$�Vm�+w0y���п�~��)ڧ. I�s�@�N��h���W?0p�؇ȓE��4���\ z.0�vh�`� P��!/�hH�B"wJ�L��Xr|iʇ"ORrL����s��бO�zp`q"O��S`��.�8d�Q��%� ٚ"O�1����\s�ܳ"�O�e�ZY�U"OJ`k&'�ޕ3�냶?Y�!1�'*ў,���4������V)u�	[��ih<	�!�p����]n�iS���W�<ɵ �x�ZB��62@����I�<Y�Ԑ<����h�0	���jQ`�O�<�b��v�B x��B��az�
�K�<�uQ�P}�I1��pdR�(�I�P�<٤���7IFU{0�Q�	����Gk�`�<�5eX>����bԑ9KƷ!!�B��:[�d�=+R��eI�aw�B�I<#o(��SBZ-������C䉷&�6Y+���)R�`�) �Q�jB�I�/��su�/Ϟ9��A��*B��(P�!�$��3�0�$��2��B��K�J��.S�x�j h�Z2v%�C�v ����.\�*���n�g��B��6wp���m]�m�
���DO��B�I�z戜�f)�(�
�U�RB�	�Q�5�d�љ'9��aa�6AB�I�y��Q�5[���QhM�C�I'�z�H�j ^v�sCB;W�.C�I.	{�L0WąN����"@Q./C�3@��%0�"�:W~t5�H�"��C�I�q:�Q�S�W"*`���#X+�~C�I�s���J<(����#W.4�B�I�:p�P��҈�D�ì�'L�hB���
�*�C� �����Ϩ>�&B�Ɉ(������(J�D��DG| B�I�S����)�ZF�<	���T]�C�	�8l�(�4����N���# �d��B䉌z@\ȸ��QT�*��g�4I:�C�	;<Z*mQ��W8r���%3OJB��&=l.���\&lB�a�ϕ8]�C䉖{���b�P�\�� ��,�:9��B��7X\��%��:��x@��N$\�B䉛G�����S�Wo��JP�R��"O4���5H6����%Ƞ"O�L��޼q(��c��N�54� "O��p#���!��@O�y���je"O��:�����X�[���4)��rw"OJ�fÌ#�eH�Ļc"-��"O8�p�̙3�U���e9�@3"O���T#��j�Д�*�)�M��"O�	��&�7G�H\���?�DA�"Oȑ�w,А�4�eg"r���I7"O� �IStD�r����L%R9�8�"OD�pl�
`�w�9]��F"O2a3a-1���`2����9�1"O��㥥�#�MF
'Y��Ï���yT7l�p2�����S)Ђ�y�L�,ذAG����z9k�/���y£T�h8�l9vG X�&���y򧀲�x��v��R��9�����y�Θ�q߾]���ݸM6N'����y��K�v����d#�]�V)ƀK��y®V7S�,��PA�Z���4^-�y��ЯC� ���&K�p�*S�yl�R�ZTq ��F��݂�����y���4���DG{�QS��yR� 0cj�J����YJ"��!�y� oU�Ɂ` �RV*�{�bB��yb�Q%Έy٢�[4R��H�K��y�nL]TP�´���3�&�z�M�y2FZs�a"Q@�:@�=ˇ���y�鐊��=*R�H6n�0�&/X�y"#��{��H�a�� fP�1f�R#�y2�KNQ�FH*{�0��(�-�y¦�%2�~�h�hR�T���#%ċ��yRg ��8�8�+ F�p)�̓ �yb�Y�V�l�#�h��Dl� aC?�yrdعq��٨�^5A���� ڔ�y2G�4�Ą@d�B,9
�`T���y��B�J:-S'A. .Y�c� �yRn]�"�1��H/Q����y2jǭ���ItB;,!z ��yr�˟�ژ0 aH��^�u���yrA�1	4T���*���A5��=�yB�G�5[�}�䥁�.5yT�R��y��^1��P"bL�;��((!���yޢ!L ���/�R_�trPGG��y�oN'veL[����gĝ"�y�hR
�yi�� �u�I��=�y� �����%F�3Ex�Z@��yr�U>J�Ҝ�#�CU�A`��y��7VXy�6 ߥi]
 �pM˂�y�b��|��3���
�(�y���j��a�*_�.�`)�ؠ�ybb�z�(��$F!8�2h�AɃ�y�	l=	dȐ�<�i��A�$�yҧ�>��%K��<;O�q��ܛ�y���?����&�)5�p%��jщ�y"Fg�嚢ݻ~��#?�yRbѮ�<��ka����c��yb%3 �=(��5�Ф�����yrG���D�-	�*�C凫�y �W����g�4/�Y#v�X�y�ɏ�N��J�=�D�VF�/�yR�K����#O�9�.��B,�	�y`+r#­���7��Xb���y���;
��[��
)���˱�y�ƈ�itȠ�6kզ��{@ē�yi�1\�Fԑ�F�'Ȅ��F���y"e�>Qc�,��'�L� �p&X1�y�֚g� ��f�yNhP5����y"��S�h̸�mP	)����&X/�y��μQ��}��l��/�*H��?�y�"�9|�r	zA�Ya�(���T��ybO�2>� �1@�Ț̅)���!�'�`�8q��r<@�3hԓ|Lu���� i�������'�%T�ਜ਼""O*]�4�XmXЋ(�(#��( 1"O�=rgQ�B��`R��V�t��"OT�	HY(!���x�&��}P:�
�"O�ݨ6/��b4���e�!Md��7"O:m��[�B��Y��$�:	ZZu�0"ORX �j]�;k -3s�
3C����"OF���R%H�� ��5Q�����"O��Z6@D;*c��sCٓw�Vي�"O(���C�4D��[�߷ĺ��5"O,�b�Ę�d�z�cĮs�ް��"O�9��?)&h�o�B�r)
e"O�a��#�dJA	�C��Q��"O4���I�l;R4p��@�)g41Kv"OР˗��� PR�q)J5rx��6"O T#!j��@��	�M%�Q"O�$�F��iN�-���W�DΌ��"O��@቞�bL� �uJ�0 ���"Ov�X <Q�<�S���a��"O��c%ϖ<TSj��e�J�]o"��"On(��$�r��	��f�PP�p��"O���իG**@�Pʤ�ڠ7Lq��"OX��H����Â8-$<Ҷ"O�ɰ��@-1q�t�؃1ʉ��"OL0SNU�O�9��K�P���"Od�S`�g�r�C�9㤽�W"O �	Oo~<�eD��6��%"O|��2��'��m;3�e�IQ�"O�KWd�m+��c�"3,�P�6"O:݋d��
�2��$=h���"Of����_Ϯu���Lg�>(X4"O�� K�T�P�j�я�x�hE"O� ;q�#�<��#.�$A��"O������5r��X�⊃)� ݩ7"O�(�S*X�6���[q�Xv"O��H"ci֩�gΊ��x�"OD౰O�:|�X=�F�HGӨ�r�"O�9�T�,��C�I�c�L�1"O��ɖ\�$�h��7���cF"O�����c�t Y���4L��዁"O�1qp��H��i�jug���"OVTrC��E}�rRdΡ1�L`�"Oh��Hȶ#C:I��{p@��YN�<��J�3|��5�rg�/KB�t�DK�<�Q�N�7�LlQ�ˀ'�L�8��J�<�dӊ]	�K��ͽj�дQ�@�p�<��+�0:D��cFc�21�&��6FC�<�΂1R,x,��5P2|D�QfTi�<!2nG "�]Xu��<�.�褣�b�<�5o�T=^P��g�rb ���^F�<�2b�F�d�sEV�9��B��\�<��ÃI�]� ,�Et��1�
R�<�A�Ԍ�3D�';���!�!\S�<�!fQ,P(;�e�,z��}�⌒O�<�tAF����g,g�XY��F�J�<i��S�9dhuI�+ ��Õ�K�<e�
]���k"%�0s��c��B�<Ya��9P�-`�J҆cEҁ3&Y�<��!�)��Z�gV�h��%SWJ�U�<a	�]5Zɢ�L�5�����Q�<�u�A m0���2���bU��G�<A��	mUM��O9M�|]��$C^�<�3����|�rg�3���@A�]�<iNN8iU�bs��2��Y���V�<� .�7�7Q�D$��̈��(ܱ�"O>��4�~t>���.a�5"O�������Ъ�L]4���"O<J������(���F�i@�"OX���"K:ƀi¦��,;.t��s"O�q���ˮ^c���S���zhk�"O�hS�+XW/��ZR  E�n�p"O��Y�A�hڦqKsn'sF�Z�"Od�p"��7Ѽ!g���>m�\��"O��1D��(VV�X Ð�FM$t�"O��CRbV�K�Z`��U5rD4�	#"OxL��m�<Pk��{B��Q:�p�"O`u��i�E�F���P�m4��YU"OV���&Q�Xa��H"H�X	"���"O´Q�	��!��i�,��#`��"O���H�I��5[��R�>�`�!"Ol{�,&AH�0��-�^��"O2c�	@���z�lӖUk4��"O�XR�.�Ut�I��E�mT���0"O�-q5!�,Pêِ��?H�K�"O��rv��=+~���q+�3d���
�"O��R�C�k|xsI^���"On�я�5wy��dU#K���"O�E�d҈X��k�m��'��r"OTpj��F=��Ss#�	��l�b*O��Rg`�;����l>��'a�0�����i��S�����X�'y��x�����J3Ú1%3�'���`B�S"%�Vd��ߖ��K
�'���T-p>�U�Dˌ0^�P�	�'����nF1F}��q��cp�	�'S(�$I�rp��f�D���	�'�V`Щ��S<>H�f�GZ��8	�'���d��JP��+sO[>j{�[�'۰4
%P�<�#C�[/�4��'������]/�(��H�
DX��'X�H��̽�$2�H�9B2�:	�'cbP#&fV3C��d�D�`�����'M�}R�G\.���G(k��X�'~h	�e䘤��a�%Mrn��'���K�)"qx4��퇴}�0��'�VibC��aW��ŧЯ ��A(�'
~��B�25謍���<
���
�'�hPh����j$���J��
�'n̸���؜)
�=0���U��@

�'��¦�H�5ZvpVa�/Q��-�
�'R����-��\�FҮ\��e�
�'��(�0�Xu���Cp��	KHĹ�'�.���!��@>j5ے��a��	�'S���䂈*#����!jѧt�nX	�'Έj�ǃ�J$|}ဍ��j�"�P	�'�R��F, ��b��a*��Q�'`X(� �]/|�~�����n5|��'�]Q���s� ��
�_A��*
�'3�!���*cn��p�E�!���	�'�P�C��_f��p���D8�b	�'A "��RI��4����:m�i�'�� ի�
 A8�v��8Vl`�'z�HJ�'��n�˕���:O�I�'�< 0���,�����1:��
�'X�T�$�ʇ\V�i��Y�1oj��
�'���3���̒iqK�l�9�
�' ���N�(r��b��,1
�'k���J�A�:m8���"O� b����@=tD��� �R�� "OfDy!fۍ �%Z4�Y_X�<*"O8�i
F1b�`u��<��T"O8| ,E�"���OY�j�~Ѣ&"O0�Q�[��zcѯ�� :�"O��(Ej�?���viֳj���t"Oҙs�A�#$��\����4I�Vyv"O��)�i<-.T�R���+0�T�)�"OV�B/�-Mhd��b�N�I����"O�`��J�(O�~���B��7�҄�P"Ofx�w���%�b��2�8R�"O2����M c>�(���5���za"O"���e�4Rd
���`-f%i'"O�mC�ᙳ626�Qa��;f|:g"Ohݘ'#��-�5S6n_SX���"Ox쯚<Zr�`C3$�*���H�u�<a'����H+�KR�\0CTo�G�<�' ��$��`�mG�+��j�HZ@�<q��ϐN�	!M�F�r)�D��}�<���=Lf0�@�eC�6@r@X0��|�<	�O���(a%`�h��v�}�<�'�ͿD��a���W�?\Z)�u� A�<���Hy��i����6=iR�4N�d�<�a��Fi�bk��j�����d�<�L1QRh��C��k�J�d��G�<a���G#~�؃A۞r��S1ːC�<�a�=>���!�������@�<���d��$�J\z�� %�8D��2�#Œ-��O���yS�9D��nF�Y'<hS'G�I��1#��5D��Ca	�Q���RnF�QY�҉5D�HV�ތJ ����X*��3�1D�dۑ���"װ�rqʖ��D���2D��jV��_\�[aɓ E��4b�I,D���6�݄y�n���g�.
����U,D�8H���2�F���.Jf,q&�(D� 1CY�<q�x�5n]
�N�( $"D�H0��H�c�\z2O�+�H�#U�5D���E�h��sց�-d &@
%m4D����C�;z�9I�N!+2���aK5D�<��V<��Q�=+�H�K&D�(�.^�.9*�� ,д	n�${Qf%D��T�F:�vy��g��=�,T�7J$D������f�B��[!�a�*7D��e�H$e.��b�lZ�+��9rO5D����F@m�@!cӤ���D�/D��j���i�Ph�W�ծo���0k3D�8 a��-BޡZ���P��4D3D��I��"t��,�.ؿ'�>��r�;D�$z��Bu�,){��"��\ZC�-D����I�8>6ب��\�@�Ĝ�*D����쌟5��:�l����LxK&D��91%
�x_�h��×�;�`,��(D� !DbE�s.��.ˉ�n��',D�����Y��;qN��5�X�(�h)D��+�I�0�2\�!Y�7�z��%D�l��*�X h�D��#�jͲ��$D�J�Hg�Բe�*~���F#D��Ӗ">e���JS�؈��$ D���ᆒ8�zBD��u��꣍<D��(&�[�R��(�u�W95A�����9D�h���pn����W]4��L3D�Ђ�ԑ�Έ`� T胶�<D�lGI��2/B���D�;0h�`/D�� ������l��5�$��8 2��31"OL�a�hԹ+Z����M�:�Zf"Op��ѥ�=GԀ�MT2Qa\(�"Ot��pg�R���@�[�VD;�"OT�"��&��pJ�Hy6ܑ��"O6e`��q��� ���"�"O��t��0X�ؔӃf�"M��Х"O�a��#F�y~����ӊ0\U��"O�e21�G�\��!X�L��Kf��1"Ö���ֵV�~y�f��& 	�"O\E ��&䊭��)^�J�T�"OR��/�Y�vkS�:��"O��`n�!�D��F�K�v:c"OZ9�M�_v��u&2���*W"O��aVܔ%*����,����"O |�ЊN�≉E��t�
��"O��`�F���丂��&O���	c"O.��vH����Y�d�h�R�"O@�M߉z" \��:u�:�j�"O0a�i	�|4�S%��o��d��"Ot�"�%��y碸�N.h�8f"O���B%��$\��pd\�Dw�x�"O�u�UK3�H�2�ʤZ7j�C�"OI*%�tg8�@$�X>�*��W"O� ��� 3n�%3lZI��a'"Ox��w��r��e[��K��1t"O^:�

M�+e,�1=��8D"O��V��
����q����̒�"OBi�Ջը�޹��i�1y21"O�Xp5k�& �� vi�l�a��"O���!��3h��[�b!jF�k�"O^��_
����T�0i`���"O��#ȝ�AϪ�����>e��"OD��C�)nc@qPP�x@����"O�|H��J� �6�ibCY8a7\I�"Ove�ď�+\�v��GJ�&�܀ "OlM�r+�0�R܁!J��#	���"O0����8^��O߷Y� 5"Oz��R�����1�( %�%+�"O\;bc�{�|���˚�n��� "O��Y�.![��uj"y��Tc�"O��B�(]���s�H�5�!s"OܕS�"�Ƙ,�6#<X�αʑ"O�l�5kR�%��!j���I��p�"Ov�[���d���iwa^0���r�"OY�C��>}��3���c���)�"O��r杨/�@���9�T
�*OX�2�Z94�hHa�1fdj}:
�'�X�bi]Eu�0;@�q��h�	�',����W0!:�̿mq�c
�'b���� e���@��O��Ī�'F�H�wQ0Iȭx�lϩ�<���'��X:U�Y YX �8��	bF{�'�p��'T����4%D�k�<��Gґ��� h���	'萷Zl�Ņ�r�活!�E�J�y1�T?M�2<�� ���j��E�i	�㗀tx:��ȓ5}��B&&Ʒ.84����>��Y�ȓ�L飑g�,!z��-�E�^��B0��cF�o�������(ȇȓ~X��Eɱ
"�e�#A�&��-��),f�G��;	��0y�FS����ȓC�H�a)͉a�l( �� ����R�XU(�H�0Y�n�(�O >R��ل�S�? �q�`�V�%Ɗ�A��@��f"O4Q2�:L����&�9	�.�"Ox�
q'F:
MFH��EH��9V"O�%Ic��o�pD���C�0�"O��B��������2��%�:Ls"O�����ڲ��x�b��I]v2�"O��`%�M�����0z&UIU"O\�A��%'<� !��X��b"O�)�K�~D1�q������"O���"m!Bj>�Kƈ�B���"O������8��t�'�]�	��"O��@�&��q�Vf�,`��d��"Ov���g@�9]����Ō96�d��"O�Yk���]N��V/t��)R�"O\���B5��HشBE<U�ĭ�"O�U���B#,��(C�P7S���t"Oz�9�ɞ"h�I1`�W��F��"O��ȒŐ]jNQ[6O�  C"O�ѻr�B;�2Q'��j��Y��"O���B��q�Xa�>E֢�C"O0-���"A�Z�H�
�;6|D`�"O� �"P/����Be��Q�"Ov<a�K�*��̐���)|M�`��"O�L�����p� G?��c!"O�����,��]1���O����"OtȐ���D�n ��I��n��b"O��=?�,D�#���0�"O�196@^�H��8�'�f�,�C"O.��%�K�M�,�!������P"O�e�"��.�t[����`k"��&"O 9���0�<����2ck��� "Otq�w�ݝQ��
P哷ky����"O�Up�ڴL�9B�Q�+rpT�"O��0���os�Q�WH��t
�"O���e�Y,@���L�	&w�qC$"O�(Cwh;�D@���!��X��"O\M��K�T��F� �\tˢ"O��j�{ÐL���)v��ٓ"O��C�**�EA�`٬z��a"OT0��h�9&t"�R�d9��5"ObH��j�h�å)ˈ ҕA�"O�hk�JX�֠0@�U)JY#E"OxPS��Z9:�N1;aO*�����y��Sj8X��.!\��Y
�!�y2��,T½!@DȺ\�Asf%���yC�M�����O�P���Q?�y�J�!�4���$�w�X�1U^��y��7���/�8L�w���y��Ư@*��1Æ�t,8�7��%�yRK��`!�&�B�m��3�Ҋ�y2�ݝQ\�<(्�oz�r���yE�'`\��eI�/��1��j&�y���U�h����#.:�x@"���y��)��Q�
P=,_�I�i�<�y2�M�SKt=��C
!��maf�^��y�l����2����
ϰ��"�ͩ�y����<��Pp�*��rh0���!�y�(��j ��fY��A�"k ��y��
! �ȴ��{���r��yaõV!��!��Ü^����'E��y��%"���N�;Q�f��a@���y��4�l�Z�)ƯY�h0��)��y��A'p�D	�O��3P���yR�� ��p���B�JoF�`w��-�y
� >В �D1^8��vꈍDۊ��"O�L��F�GC
��6'��A�0-�$"O��B�-eЖI��k��2͜D�w"O<�ʒa�%x��Yj5��_+0��"O���#.}@���p��c��V"O�h���ƣp%x-a�C s�ZI�"OZ9S�O�vLM���C�� "OT	ID���}����P.W�Q�Q"O`̋E��$b��U���-:���0�"O��w��<���69TFuB�"O��!�lIͪ�sD��Q���"O�m(A�ݥ|��Rf�;L�����"O|��Ǌ$���!B��lz2���"O�s�^!k�ũQ���H*M�"O\����*s�a� σ�Zk��W"O�1kC��)Zx��,cw���E"Oj|d[�|��0�uh]�
Zr��"O�hҋB�*%�PӝxITA��"O� �͜�c
;��0>�J��E"O^b�k�/��ԍˣ;8 �: "OF��P��3q�V̚6+P��"OZ�QU:�V�:6n	%]�|�a""O�P���rʌ�6�J�:��"O\	L�RQ�Hs���d]�u"O����F��9(v���kD�N��B�"O�ip&|@2��C�����@�"OQ��I-F���'lSA�PJ�"O��u��1]�݊����k$�u�"O����#
�-�&D8�@)6 �b�"OD��F䓴�B���M�D�z�3
�'��1pцLsBp+# X�o�4��'�X8��]�:�`�hbh1w�5a�'��@�b_�Xq��O&D6��+�'�����n�l���b��'¢���'��1	�^gEd�C$���;�'�H� �%[B��
Q����P��'!����a���! ��6�Ju��'��s�nJ��0�)S�0���'lN8	Bj�-3@R�9ֈ�=~4�1��'9��JŌv}��H�5`�v�[�'��	��˒F�8��C��S^e2�'Vxr��@�8<�"\&Tɜ}��'���3��h�x�p�˙�E"\i��'肵Bc�۟k����
��	�'}��C.ay��7Iդ�bp��'^���F��:��fI�-����'m��Ha�¿:qV;&`
5�8���'A�q�V�ݕKH4�+�/t�mb�'?4e ��۞?���b��_;z���'n0�0d) s-�����X&�Ѫ	�'�H�(�
[��9�dˌIA��'�t;�"�VKp���C\(�0�'j�E�!�*����WE��&@1c
�'SF�U#J,~X8`�Q�A+i�T��'�n-C�ҟ(A���i��'������5�dLs����t�R�' �t{���x_0أ�������'�N$[��@-ir�A@ׯ�}Ů�*�'� E�т� �s�/�4oܢD��'�&�ۑF������LKt���c
�'��QO�+>�ր�!���]6f�i�'��H���V�lJ�p��,*���'�4mЁ�݉V�����=)**��
�'����%A?$T��eL!%>l��� P���,�|��B�&$8�S"O�X[#BI6>�����NJ��"OE���L��у� 1:�2��7"O���6N�v7�$IT�xp�"O	�@F*!�L"�&��I�XY3�"OFȩGNF���Z��=jk�P�"OƁ�햒H(��Y�k`���q"O�DY�d35]��bJ��~��"O4�9PMwpA��&�*.���2"O��!�ډj��ukpY0�:���"O���!?L��%�R1!`zM��"O��p��� BPm��ǢDk�d��"O.TQGeGL�������x1!j�"Ob�y��2���3�F3?��@�"O�$bMF~O��ڣ�����I��"O�Щ��Q>��=[4
L E��ɱ"Oq�3B�q'�L�|��,�v"O��v��5 ��|�r�����"O~��g����e#��7켝�4"O������$r�tk6lL�J�@T"O���F�T��̩K�5�� "O޼
WB�.^]��KۖwH�X�"O8��rD�1h���B#��Jlj@"O�Y8c&Έ;��"@��ЩC"OL�"��G2��`\
n9|��"O�篂'A~�:
��h��r"O��aFM$b��B�H�>���(�"O̔��f�9oZ4�-B� �4��"O�|��ՀW����h� #c"O�a`���$oP��4��M���"O�񋧌�A�p�caG_��d1#"O`) ���%��0V @8
��J�"O6d�.-&A7o��@	aU"O�%�����42�M��kE,z�Н��"O�a�`��`X�;#��0جM�"Oj��e��]�Z�@���(� "OY���._��@�3�īz6�J�"O�){w
�_c�X��/F3t�4�"O��H&�:*d���&B��g"O�,�k3��`r�?`�F�g"O�i"� �X�Yw���T���"OP�ѧB�}��ٳ�,�"EL~�Y�"O񈢀E9J'f�<Q�C=0 !�\�#$^�A3L#T��� �B[� !�y���t�Ȭx���U#S��Py������Hud̓-)$Y��:�y�P7\Z	zWoׅu�D�J�&��y��Y�iR�ɤ�gNL��ʂ��yA��_b�e�E�A���bg� �y�Ri��|3�K�
����ūL�y���t2��%8-jT}X���+�yb�7n?N�1�m�$�P�`�O(�y�ɔE����E*�RQ��*�y�%�+�8�Kt!(F����e���y��G&��b`�>{�����Ȇ�y�0nI���oA7qT��j�)��y2�G�M��Ӱ�ܱ`��y#è�yb@P=P��irGC_��Z������y���:Z(�휘T�(�R �y�@�8pĠ�[2��I0���6(��y��VW̮MB��Hyn��c�֐�y�ß�J�t(�RȖ�J�����"
4�yr�ƳcV��V��y_\��6��yr����HcZ�j%P��M���y
� ����.��&]bt�@��\ic"O,���3���%H� �`!"O@}��F��"�ޱZ �Y'���D"OJ����4U`(��IS�&�� 95"O|40E��Y����)�/Fh<�R�"Or�å%C�l�L���`1�<��"On�`@(ފ��s�N ��T�D"O����Z�S�ā���M~�S"O����.�?�)�פD�tR���""O��e� �%B��s�b��#"O�飄A<�2HU#p)�T1�"O�ĪR�,� ����X��� !"O��C�%�V�� ʋ�v�a"O ɲO�~�kCXttJ��"O���C�_�±X�DA�|e���"O:}�d�:�:�s���S�|x�"O�X�6�W�^�`�)%�~%15"O�<c��Ę X�(�Bd3���j�"O���Ã��	b���㛆x�$��`"O��ڠA�/bXd�+'�E���:5"O$I��l)����>8�� @��y��E x$�IӶh�DqO��y�S4a�ex�&�g��Y�����y�*����S�Z!��p��yb���a5��amL1�,S��^��y2h����$ E�@&Z	�rD��y�LT�SB~�#��0��J�yҬ�	Be��a��J�f��Q�)��y,Ѿu2.�s�$��X���N��yR*�;	��m�d�^;	��(;p����y�cI�H����C�μd:/^9�y��מݶ5�#�-
�%3�釪�yRNE�6+~M� ��(rڌ9��y���5k4��� i�8\�� M�5�yR��Np����D<��{1� 3�yMx�T�Å���k�<�ࣚ��y��@��E�`ލx���q�/(�yB%S�_������0x^uZǏ�<�y�`<� RlQ%�v���Ȑ��y"��2�,!���f&�Y��?�yb�P8��p��._���a��yb�чKQ�Q�`A����Ȣ�y�$::����`�V���)�j̷�y"$ֈr�;#�B�����2�y�)�<l�|ٔ'ç��x�!j���y�@�����I�C^� �o�"�y�	4#��0&Z4=*̹�ԁ�yrG_�It,,(gM�+Fİ�M[��y�d\Iz #Q#��Z��yqi��y�G�b���Hݥ$�^-�&
��y�	?I��IS��w��`%��y�
=z��1&H������O��y2ғ�49o��0,0'���y��^;P�H�o	��9��Ш�y"
ߣ!�2��oQ�T9�(����y�@W0e����J��@=�1@��6�y�B]�/hHM�vK��(ɎdX6h��y�A`���Ӥ��"��|�EkI�y2�� Ғ�7Ϗ'2e�̡��٣�y�o
�
Q`u�)a5v$���!�yO��1���\�&X���v�+�y�(h|��P(*@��Kv*��ybFJ�XPv1�	���<�ŦT��y��M�`������tY��$��y
� �X��c|�M˥MK<@l`��F"O8�U��]���$nK�O4l�y1"O��C#ΨO�8!�d̉K��(H�"O��(�ʍT��ȏ%�4q��"O�}�A�k��00��U�Nq�@"O�@"K�1��H�$=q�-��*O\	z"/J�_rdy�=S��0�
�'>����#B	��a�͋Ehy�
�'���R�]i��K��.�q�
�'�m��b�K��h�̚�q�ʱ*
�'��A:��H;"lt�"��T��t��'��E%e�9b��1kG�;�Jt��'GFl�T֕���������'����5��G��c�M!���s�'rP82'D�ބ�"Ý�#�
I8�'�>1��A�eX��q̏+���'%��*��P�
7t�i4��Medx��'��ҕ�?*n���d�-sz���	�'<0X���<x�ܤ2�ˤY��(:	�'`�dK�H0+�X]�A"LW����'�H���oY�a'2})!��R�MC�'(�IY�DI�Q���ra��2p��	�'�D��v
ٰk��idK�
)#�d��'�~��W�)
�����w9RXI�'�l�(��ĩZ`�Q&+W_K��r�'�ٲ�"�*}�BI^O��� �'��\�@G�<P����"�E�����')�%1��:ҍsQ�L�Fʚ���' ��ဪ�4:��ؕ�S45� I�'��yj�ՙxȆ|+� O)O¨ �'�x�:��?I.E�������H"�']�Lg�J�(��Pأ+ڮ�,u��'u��7!�!ĚL���
�=�5;�'�\aÁ
H��K��S)wx)�	�'S2�*�N�:��yA��$=2b ��'��ujp/<���(�aD�kyx���'Ú���#G<i�R(� ��������':P�F��1x*h�����'(O�9��'�n���-����M�&+�U��	�'�b�bd� \�2�x��������'�2(#�⟷i�j�I���^��A��'�V�9To=z0+f+ج""�k�'� zf���Y�j�9e���ཡ�'��ق��hA���%��l:>5��'O��!���w�L\y��5�0;�'��[UŅ�4Q�0Jamƽ4ܸI��'+�HIeE�+�^�ڡJ��+p�d�
�'ްi$B=�I[Q�
*P��

�'|�������V��FށB���	�'�<i�2�͕ߨ�@u�$=��`	�'��\��C�P&0eOS4]�
�q�'}H��!a6%�p���d�W���R�'ߴ�H1�P0����7��Ulz���'��]#��� �>=3�#R��-��'^F��L[�xB�hR-LYh���'_x�h�/g4�b3�D�o"@���'�aR1�. Vd�3���li�5#�'`��e�Lt��s@�D�a��'iq:��_I�ԁ	��@!U�����' &$*� ^B�a���Aa�Yp�'����2��v��x����Dyx ��'̓�@�-�Z���N59�N�c�'�|�蛰R��j��C�6R~Y�
�'�Xс��ƪ<`�3�lڌ#:�I9	��� ���5ϝ�[���� W7
P�x��"Od����\�F|�u���
EJc�"O2���Q�}� �Ps�J7"5"��C"OV	`����l�8�B�!�lQ����"O��@E��T�^-3A�		i.�b�"O��PdjљYHȨ�Ȇx"���"OX��lS�ƹˑ�D�x�Xc�"O�y#�F5q���s�S,K���"O��4��:}XUb'E�?]~�1�"OdDC��3���i!D�!�z��&"O�Q�/�c	�ɰ�`��*Ŷ)bb"Oj�H*�Wl�|bƏ�~�a�"OHTP�@�%]	�t�`�ZUv���"O|jdO�},R� �5��  "Ol�A�&ˌd%�!��P�r��9r"O>0���J$&#�g��X���t"O�((���	0�!���21&��¶"O`U�Iƴ50$9��R�P ��"Op�U�U�!;HX�p��7�
��A"O�pf�E�@��9 3dXC�8e��"O0�@�	�ܩg��7y�Xځ"O�#+@V��*��9���"O�8�7��aLb�(;A L8�"OB�k��;��9��3V��(�"O��au�˓j	z��e'B�-��"O�q�f�Ɇ=�q�S�'>3� i�"O����c�Mp�[�&®U&�@`"OF�J�/X?-�ܤ`u��; u�yA"O���#Ä~o����Iy�)��"O~�@��:e�K�ƳYw����"O��ÍI����8%A\�s�4Yi�"OH�9V)�4T�:�i��\�U���R�"O�li��q[bL�cm���Z@XA"OL	�F1�p-:�L'4��2u"O�I6��!IR@pG ƥ&��t�"O�e��ßD�N9zd �b�>�Y�"O\Z�AɷE:�P��-Hx�%7"O�d�&���(�#�Y�xT"Oxȉ�ȋ�,;�"B9V�p"O�tőK��Y���+O2�e+�"O>d�C�1*[���@��c+��1�"Oԙ���ҧ0�,X�o�Jn���"OV��=/�h��m�v;<D$"O�lx���8�<��L��b/d}	"O܄yp"p�(�,!H�"O��1�ՠf����_D�$"Ol!���r��;6��'���"O|��SJ]Q��l!C��5)� �e"OV#Ċ�3��q��"�
]� �SG"O�ls�:�������'[JU[�"Oj����:Wh���ӍS1��Ö"O|8W�O�ԑ�́,Z"���"O�d� hj�xWk�u��`"OT�ؤ�^#%NB�A���ge���4"OʴP�Y7F	qU��V��K�"O0q��A�6�@�pu� �>��"OT��%T� jp=�UO��{%:�)�"OH͑�%
=c�Z�ك�^G� p�"Oy�sM�#eK�ۭ.M`H4"O�eco�)�P�A �mI$ 9�"O��!�)F=y<� �۲9E�Ց�"O]�ş�[��ek�.�vΐ5��"O@�6�X�rـ�MT���S"O��A�.��alb��� P���#"O� ̡pa��+!l2=� �b�"O� �1đ4����W�|�f�:�"O��ʦD�&a<���Giڲ�.8��"O*Q�O��U�'ۘa�
���"O�d����7w��D��&rN��"O2��S�[��E�N�taj]�D"O�y���ٞ'E��񕦛;}P�S"O�1!4Ϙ1,����$V�T�^L�6"O|1�4�őK���pv��9��"O� ��K\}Ը���8PfJ��4"OQ{�N�Q�t�@
��dg�հ"O��1�C`�����<t}^5�"Oҥ�C�5>�0�`��N &h���"OH$A���f0�� �zO�,�"O����׽</~$�V揗_����"O\u�5LF�F��}�`%Y5Ρk�"O�-�%k�Od�ҧ��R6����"OF��*C�5.�eQ�N�%4'v�)�"O�9WM�f���	@��.��X�0"O`��C� 8m�Z�X�-�#a�r�8&"OBɘ���XQ��)�m�c����"O�4'w��A�F
=#�R {"O��q���}�v0��?F^��T"Ob�J���P�mJ��U6$:�H1�"O���f�>�N=� M�f3�x	 "O�Ӥό�xH�#��|&�9x�"OZ�E̘,P*��#��l\�"O~=���D>Du�siTiI"Op��@ӷ	�4���	� N��"O
���Y�$(:�@�]��"O�3�Z�!�Ēc狏n��8��"O�C⣜$s(�)�:~X��"Oh�8�g��<e�Ȁ>B|���"O��4��<ڸ��%*	�5H5"O����7]���#V�L�R�b�J�"O~��p*΁g�������:7u���%*O����V�*eP���4��{�'lp�pah��C�^t�B�+M��'j���ޢ's>�x�aҦ�f�K�'9N����"|x�`�놩Q���'K���Ō�?�T��ː�pW(�:�'z݀`���o�������4�[	�'�>���9y��y	ĥ��w��5 �'`9*�-F5
������\��
�'���P�Cݚo�$-�"m��m�P�p
�'&����㛊{}��%d�	P�h��	�'�Fʂ�M2��<+����:�
y
�'~�tѦФ
Ő�*ٗ3�j�h	�'�(LL�3�U�H�&��y��'�z��e�DO�B�s1	�"^�b�'ʹS����d��7)D�0#�'��`ڗjA,rĂ��̴AB,#�'�$�k�'X�j���!(��9���C�'J�A0� �nS6\ ���g�:�'�a��
C�4np�Ɗ�Z^ha��'�V���A%�N`�Ux�ѡI��Py��	z�"��Ki\�vd�u�<)�'�yBX�%��"V�i���p�<��+@:N��FS�jX�����i�<�'�Ҩ5�,�ҕ\�Z��$��g�<�T`C�_�i��e�8��gQM�<AtK��0�hIY�&Q�K��	uRF�<���ԭ�R,y��/Wfy�e�B�<ɰKT%^�N ��	)i�P�`�}�<� 4�*)� h�$�"
ćs.9#�"O�	qbH6 ��̣�(�H�.xS�"Oj̻�J�=w����f�nu�tJ4"Oj�3�$U1M������Ouab"O��UbF�w���2h�8�R�Q"On���1/ra�l-c|���"Ox�r(
D8l�LV�Fp4�"O�(�2�N�{�P=+g	M$p>���"O��SS^�B*"� dkɵL���s"O��1�.�L䊨L�~�jdY�"OL��Ơ,u����T,�qT��"O�e��dKT�p	���N�`Y�9C"O0���^z��+�b�d�E"O��P��1Q����kھݞ�)�"O|ɸ�&ѝ+�$�v�=X�B�ٓ"O�a��A�$�� V��^m�e"Oh9��X (�8)�pOށ]RnP0�"OΘ���4`~��Z4H�G*�k@"O~�HQ�Co�$���f�7)5t�"O!yEeQ�u��9X���"d#.%��"OH-0���J�$}1B�͟���"O��#��aN\�y��5t�l�"O����M$$���C���$)Bd��"O��J%�ɉ�L�@���^��%"O�5�U �,�)�(د) ��z6"Op@NH�(�d���hB�QCd��Q"O|ha�ן*��͂��x*��;�"O�4�͘^�6��'L����"O&��Kٰ0+F��l ��w"ON-`��j�B�*!'W,A�>��"O����/n�*x�GeB�#��e"�"O�A)�OY�(�K���AP"O�%�CB�]�P�v�L=c�����"O æ�[C�H0�`�[���b"OF��sǏ?Q��Œ ��t9����"O���])���A�\�R���J0"O�m��iJ�=V�LK����q��ّ�"Oz��r���nH(�/y2�=�"O�(U�X%iHV}[en�?�	w"O�$`�d8Tx��#&n�T�8�"O�@��I�7�*p�ɺIݼ �D"OҽꖃU**������>_^t!�"O����[$F���2�j=S�ذ4"O�p��H#`{�)JP�q���h�<Y�ڙe�@�R���$G0(����L�<�qM�@��`���	&m��Z���I�<ac@ɼkc(h�� AX���g�]�<!���
�2��B i���P��Tr�<��V�̺��2O�}�hȇmFV�<)c��p�j�H�,`�X�R�<I����:��l�Ģ�J���s�D�<�@*�<�4��LE�[�5 �QA�<���3oP�2@�L��!�y�<A c�o�HȤʊ�32����x�<i�.J
����ޅQ��i�e�y�<�g�A�B�hy� ��@����T�Q�<� ��21ND��h߃b�� *W�<iCo��N��(aDD�z�\"0n�T�<)�i&I�ɺ�ϋJe�u��I�O�<i��D�h���R��Ll>�jSK�d�<�r�T����ԉ�u��'�K�<�&�q4�aԈB���h�GH�<�mL';r�}�o�Q����t	�J�<�TJ�CNxPka�u��U��N�<� �`A�Ȅz��IT��' ����'�.�<aP/8
A��R�̀��E�z�<93�D�FQh�0�-
9S	\!Q��y�<����V��c�8f���0�I^�<��,Z ������� �J�0U,�U�<Q$��:`@�a� NJ9(�D�ҧTX��Ey�&ך6u���$�i^N��n4�y�*�j��� ���d���ᷯ����O�~@��u$�+TdX�P�I"T�I�<9���v��\�󣍩Sj�8��C@�<UJè"�p�sRMإN+L%�1D�|�<yp/�?\����)ԤC�0�`�y�<I�b	T���k����0��4@�~�<�GI��V����1r����bL|�<y��F7�2Y @�T?K�n�2���m�<��G�T5��"�{]#�P�<$�5���hֆ�8��3��H�<�w��CQ$�rv�)n���+�M�<�A�K�v+�T'��J�����KM�<)��ɑ.�Z���I�+d��OYE�<�c!G��8���*��xq�A�<t@0N��������63�l�d�E�<���5�֝i��X�����j�A�<��b»7��� J,@:�icL
w�<�2����@AR�*O�(�v�q�<�"��,VC�X����</l=�qA�o�<y��ęVh~� �P�Aw�m�<A��O�i���ѣ���8dYDM@�<!�,�=B¹�`�ܖ5@��U*�C�<�����Z��x�6.��~l�T�"DV�<�f`�WL�d"��$)�d��l�<��jq�$iq 
8n> �FcSs�<�!���a�^���e��Jp|x���u쓾hO�OS�Т+Ƃg�fY(��V&e�J�'Uў�}Z&bO�2�K��H��!r�,t�<9��W:a_xe����6R~6tز�Oo�<Y�֠E�x`����(3�����i�<����	��0�����#��e�<���V0h����B��e~ȉ����w�<I�lF)>�mU�� Z�<ۆ�s�<��)krZ�r�G�3c[xA0EMDX��T�([�ޟ#pYZ�* �NT�4D���޿\�� ��Ü�,�T�s�4ړ�0|��Mf����V��]�ܥ����e�<��Wk��y;5Z�'��x�p��m�Oҧ�g̓2z��`��بj��Q�Ө]w���I�bkSg�� %��q�*!��Oɳ�y�f�3V��a���l�:,Rg��0<���D�'P�(��c��F�.H�F��&U!�$�Vr>5YK�8��,k0c��w`�O\��D�Aa�l��D�.x�du��	�<!�$D�z70lBC�N�cX�ۂ��(b�<��ȓ[A��آ�y��H�Dr�D��Ʉ_�4��<!�����Z@��T26����䔪��'�az��B�J��q���]���d���X���M���imc�\��ŀ�|��Ū���!��-T�����.���aC��v����Ó�ŋӛK�NC�G��8�I�d
,T�4{ L�V�DZ5NI�PNv4
�'�!�d��<��T��B�E�ĭ�!hqOdO�}�v�S�Hd��5���*� �5�A�<Q�$�3��1ө'F���@�f�}�<a��\�C�ٲ���!Ɛ�ЦFn�<1�,ylqr�� �L ��am�<� i��˜q@>i:��b�zm�c"O�T�$E��+A��٤�Խ5��U�q��o�OtN�4�K�@tt #p]�z iQ
�'�4�8jӟ{���*¢��
�'��١ ���,&n�D�%�r`+
�'"��d��pJ��f��,"u�a)
�'Mu�U'�2c��q���!���
�'l�x�G�8R�D�J�*��+[ X�	�'�v������H;�Ș�Nm�����'���F��8��q��j�`��'y�ʳ���h9��  ə5[�X�	�'�1s!!�X@ &�%\i �)	�'�ش�Rԉ,�f��*ԴE��{�'�Q��bWijȼ��-�::3mY�'f�P% ȸ@�͸�L�;'��9�r "$�hAd��0&4�r�f�i��R �=LO���>���3P�8ԓ��.q�~� f�Gu�<�_�(q��F^�\zlp�K�X��C䉰^B�B�&$p)�!�+F�BC��,�1�Ҡ���B|W���'�a}BJ�p���&B*n2�K����$0�S�)�>W.�/,Z [b̝==9(�C2��u�<1�
�c��٣ H�"#�<0��OG���0=Q�+E.� �r%$\7���C�<I,��z/$�kp��0IWd`GbJ�<�aaM��ҴA�kQ)p���#X��hG{��)�1H�]9�舛`x����ۺ@��C� W�u���]�@
�Ҵ�X ����0?([���Rp�Һ�PTS� �e���(���$�)�@��ڸ��|5L�!�d��)M���S	4�����@�G�!򄌞 ��A��4L�^pyd`_�7h!�V��.5��L�	��)����:��$�D��h��9x!g~��slD��""Oj�#�%�'Y�=:rh�6��x��"O�����.�I�(�9v`�u"Ol��F�NJ
eBE<8n>��"Ox4x�$֢t_t��S��3��kB�'�˓��ɓC������!M����%w�7--�S��MK���!H,D�t��7�4�	�V�	L���OB��"�h�]A(`��x[@��
�'�z�#���#|�`�Cb�C��,�	�'�PYB�,n�Թ��� J���J�'��ۅ'L�A��P�b�8F ��{r�0�S�x7�9�0��_^�t`S�<chC�I�?�5���E�}�F�Qj��d�<�˓TvY�*Ɖ$9x���)$����zv��Q�k_��2�R�"���Lp�ȓ-�r8���2,=�q�?>Pd���`���c��?��� ͳ����jwf���)E�% 6gG�ö`�ȓz�%�@�wjH��Z�h5�!D����׮���%ih��r+D��X-I&��ؑ�$K�R�H6(4D��I�ȧw�(]R��/OX ���1D�(��$O%<j�Jv�i��)Q�0D�4 ��Zr��B&��l��c�2D��i�nE,^HZ�Ϙ�/wPLHf�5D�X@�
 �z��B�q�� �M'D��@Sf�e��`�1.Ѳ2��Ţ`�%D�L�F �fA0���0	���l)D���w��
0�zͱ1n�$w�q�o4D�d��V�;�dɹ7�˟-_����/D� +&�ż7԰��$I�G�����8D�� J�J�Z�A���eHa��mї"O�Q�E+�b y����*J �0"O�9�s*��x+~hg��+
��"O�e(���/��d)q�"=�԰a"O�r�ŏ�`^��C��ܸB�X��"O�d{v�s��A&��A���F�^�<��eкlB���F�/F!iA�p�<��@J'd�t�%�N�7֞49$�i�<��K� ,'�P��G$ZUh���l�<��E�#
��I��%��9����B�< +�!"���A&ٟ|?�E�Ǭ�x�<	t
�2Ia�h+��Ȟb�R��Vx�<d�vBj��a 1�ܩ� x�<��*̘Pv�2��S��a@�
�q�<	&eʍe�^\�f%H�[ @yx1O@l�<�W��?\-!��E����!�R�<�d�?�j�d��k~8pPG�TR�<�X��b�1�tH2$ï
�rB������:bE�e	s�]�;�hB��<�,�!Q!5!����㚠K�C����!��� yb&s�"չyZ�C��;8���xL�$e�@ꗈu��B��;X�� ��0=�u�B��Bx�B�I�L����ץ�����J}�B�I�Z���ALM+ ��+�@����B�ɔc�6Ye���D4X88�� e��C�I��XŻ&lo%�)"F"_�VjC�	�,2�k6�ֆ�z���,؝f�6C䉠(BV��	S��R�`�gֈ	�ZB�I�Xd�C��,uBm���T�@B䉸(�̐B��)�2�Qů�1\�VC�	���3��5pa
�r�C�5q�=�S#�$3���T�*�C��7@%��y/֐>���9p��iTC�	�RzB�Rg��,C��U��e�lB�>S�~�# �[?1�V�*�mݼy�B�I-'�Ԁ;���+y�� h�k3�B�	�Ck��C�k�-+���%p�B�ɫ �AҰUf���ۑn=*�C��>pn�@u늺3 �9̗I �B�ɫ,b����GG���͋1j�76vxB�I2��5�hZ	J���@�D�mhC�I,F��50�둤W��¯��9X�B�ɨ!�J4�2��?ו���oDmr
�'_�a;���:n�`2	l�"l:	�'�@�w��4���шP3a3��r�'E A	BOH�>��3�%C����ʓO�0($�=~�l�� �B4ن�(�m�2�U�6h<�!�'�	}`�t��{�uP�dD�]�j�T�\k�����>4�1iH�NZ��Q�a[9b1\�ȓf ��c�c��5%3I���'0D�(
���/�u�Gf�9��D`��9D����ȍy���%={���$�,D�@���
&1�[� �~��9�!I(D�����Ae<<:���=H{��j$D9D�X��"U0��1��2jl\���5D�� �J/�T�B�U�@>��è3D��X ʄ�K ��:����?OErj3D�P�wMV� �p1�!�X$��L��C1D��E/ׄ3 LK�m
*#���93D$D�tx2O�L�f�b���{�L��6�-D�,Y���Q�����"O�
.f��7?D����,"�M)�I2�nٳ֍=D�� X��A�G�1��IAB�i�����|��D0��'��"����qj��:�<i����y��5i/�0TB�l쉊�nŕ�y"�˓F�6�+"�Թ*�x�#	�Px��iz�h��%>e�1Y�@0~V^���'��`@w�B'\��0��CPn��q	�'�0�Yʆ�-�L�m��k�B|�O>I	�5��ؘ��՝Y���6k�O::ه�M���;+*����a%X���Au�'k�x��<-¬�vF_6k�@Y	� ��HO�OeS�O�}��w�x�ȱg�t�\9Ȉ�SM��j���GgK65�H� ɕ�z{�5�<I#�"����O���㔀G�V̩%Ģ@t�e�'����+�J���I�:����G�i���<1�S���"��`�����IpZ�iO��E{����B�0��M3��W71Rb���̯�yRH�*��4���0�������'�(#=�'�yB�C_���a3�	?(H��	%�Px�iS�<�עT�>$is�9xD2,г����Y��~ң)����/c:BP� eF�sF*�	r�I;feJ���c�4�S�9_U�h��=<(��mZ�Q��6�S�O��<���(�b�h@�κrz���'L��т$���* !�;�p���'+����ʀU���`�X-Ғ\*�q+�7�T;`�1�-�U4I�q�5G�!��A9�x�&�(��Ѳã,�Q��D{���� e�ڮƄ(�"ťR�
1:��5D��z�d@�.4z��4Q���p�2}��)�SK�����	 ���m֮o��B�L����fQ�e�����D0�$/LO��Pk��
����d+ʹ(t���f"ON�(��ˁwL:H�� Q/E2]zp"O֝���T߼8�o["Tc��1t�>��+ҧ<<|���ͤ>��)ЀM�mzx�ȓ+���0�	T,轛�!`��ȓY�,0���#0ˬ�b* p>(���M�w��v.ECA�n\x1�GA��ē�hOq�Xa㒧�L�������O3bѫ��'$qO<���ةA@R��R�\�;��z�"Oq���̅���v,NF7*���s�'7���9ot�����r���L���B��#E�@U�$ ���\��'�ց=�0�':ў�?����x�����k�
4[Sj=}R�)�>����M���U[�^��ؒO2U[����ކ=��Ȁ�o�_Kl=" ��=G^�<Q��>I"�� ��A�/@Ў��$�Q(<)ݴ �&@IC(�<j�8�$�2~xy����	��MK����u��i"R٣�޾,�L���hR�M؀3#�;$�ܙ򯒝~�6��+�X�<�xSD*D�x��k� p�B\9�<sX�ã=Of��ēu؞�ۄ���m�D��H@�.���>������"[
l��l;G��҆�	��yO��>�R���Һ4�P�Q�(���yR��",� S"�ޡ2x� Ý2�?i��$�8��'�k�� 84Tyl�2�V��%?5�!�DA�H�mAVH�3.��y�&�-t!�Ĉ H�LD1�([�@K�u�%����z��'��_=��3�A�������\�0�Z�"Ol�c
��e�&�e��"+�Ⱥ�"O.�(B�~� ��1"4PQ"O�A�G6�N�j�.H'B���S�'�Q�,�'ʱ��]XB�Y�K�6|0fM̂Y�R"O�P�K�;�Vt"� �xA�Ѐ�x��'��*G�&�쐒E�O�Ү��
���y
� ��x�ʛ��1� ��nDA�S��ϓRў��*`e�˥K�8h�@�@S��u���	���'?b�pt`��g��Y�Z
/��h*#"=D�!�d(�@	{7LVھ���
H�m��|r�Ov�I�"�\yȁ�����A[�K 9�n�T�'L�l:��±_�B���6:N��/4ړ�0|J�"ƞc�`��pU5 �0�Wfa�<A�e�Fb��A��U�x9��q n�Y�<���c)RD�fN5~��H�6�NT�<9G!S�hڰ	�.U���0�aGS�<�1BȽ\��3�Hǂ<�JYzV�Y�<�k� ���DIA�L����X�<�!nLd�Ɠ'	����V��M�<�1�J[����𦉣vuBt�Ȑa�<�cגk�EJc(S0doUZ�<��ɼ <�"'H4u� ��o�<�3�3�0�����B�R���'h�<	ϗA���I"`ULw��#�k_�<!�h�:`�ļ�2�:9���^r�!�D�!9�Pb��PK~<:�ńm!�$�$x}�g#6[,F͚CŜM`!��Xa/Z�w�ݖBD�Q��D��<b�y��O��Io](|B�/��FMd,�ȋI�C��z(�]c�f��a�8����?��C�	�4�+#�2֐*@���&
�؏�d<��]8u�
R����'��}���"O������ U��-d��q�҅Aw!����P��e�A	}� ��! �Y!�$����ٰ�c�� o�>z�!��S�*wf�Z'q���)pD�@ϓ�O��"�Qr�nX�� �j��xH<ɒ�ǉi��E�u��0یô*�ty��=�h�s�gJ�f� `�7�Ӥ+zC�	#<���u�?D��Jb��fC�^H�`��7a� 5����B�I怸�q@�17RX��V5P �B䉑N���/�?c�DM�2.�NC�I�o� 0��-g���*E(U-��C䉹;�b�7��.j�Hd,R1戣>��'�>M�wV�- J�P�cW*+pRAs��7D��K6���)��0��5���z���OlL��JBx�93���aOT��^��* �3�>�l���/伲!��<Z%�B���I[���Mk��d>�	�7k��2�o:8 
�O���E{b�xaD/A�@���r@B6�U9�y� �6i�8�f�F8~�AS�����<I�'k��ҟlH��(6$�|9$IʀEuٛ6�-D�����]et�8��II):�Pw�?T�l���ŜV;��Ť�+��`S�"O���C��4��I�U��A��	M8� �Ç�;y}9x�Ӱq���1sE9D� +O]�T�E$8Li���2 �<�󓁅AiF���#$3����@Ui�<	3�D�+l�Q� ��l#��r���K�<��&�#_o
9����KX��f��E�<�f�L�bP��1P�v��I_�1��x�?y���~*��ڊz!� ��.h:	�v�u�<I�B�1Ui�5�U+�Ԗ%�"i����IL�S�O����/f8��e�{c��""O0gɳ{���KE�Ur�/�y�	�%u�]R���p�"�ɇ�S�y��0zT��(�1k���'���y���fƈB���f�|y�W ��yM��U�$-1��[�sVZ�� ��y
�  b���| ��!�M/���j�"O��FV�7���8��M<'H��"O0Y��3�t�@�Ա?&��"O�MI��
%����n��,�(��"O� Si�#��EBt�R�+6"O�@���b��xx��C
�F�� "OBa(�osXd`t��*�HJ7�0D�(��F/�dU�0��{�z��6e0D������~��܉�h��:R,�Ԭ;D������<�JZ�t�2��s)Ot�<�.;F��)����y�%���Gn�<��Jj9\��4a[G�������D�<�5�L�B�d��A��]���谂�f�<Y�ቦH�4	U"��e�<th ��k�<�  M$�ub"��\��@��B�<������A��L�L�S6,|�<�t+ғI@@�����k����t�y�<ٱ�OGM��kؙW(����s�<�5� �?�*5h�c��s6Vqa�/Ro�<97�P�fXz #;&怀� g�<��MC6e�X�D ǔv͔�@�`�<a�'>ڦ%� ��w�ܽ��,�g�<�G])}v���T17,��e��`�<م��E���0��F	B�| G�^�<i�#آ9�P
Die�4C� \�<��(&+<a�#����}B��V�<  ��:���e�8jIZ���Y�<��@ϴA�x��T���7F�,rBq�<yt�Č�c�H���9�X�<	fn<�2�K2̞=�2d�C�W�<�等�#w�E�AX'P��`fȑH�<���\�)@�����kՐX���G�<���Z\� �@�tԾ�Z&*�j�<)cc͇`��tX�e��{�����.D)59�@p6Ύ��>a�/9� iJ�e�
�d�H�<� �C�Щ)��=��d
���H�<��.�q���e�5R��9�I�B�<���C��|�@�^�BU	fFOk�<ɱ��>^�����a	F��qV"X�<�#]|����AC�YTp��T�<��	��]7��� �����y����P�<A�/̔���� 
�QWR�<A1�Ÿ�r� �'JEd��'DF!�y�
��j�@}���C��w����y"	=`O4EX�֎(���	�y���=p��g���"Pa7C��y�Í�F�&ܹ��8xZD�;�yዀp 4t���Qr����p!@-�y��7_l�pR��M&h*�-�f�yrK�w�|{�e>�컆���yb��(T=��I��?_(h.*�yª�8U.]�sF�:��� n��y���?{^iiv�h�� ��y�Մ/M���ǔ� ;Ȁ�M�;�y"&N%F�ޅ���2SR�M�'�#����d����H�tr7��w��$a�.����s�+UP��'JׇO��P�D~����	������A	N%y�'��v$��'v� RP
�+=0��дQXzt��E�����#�L9�]w��U�' W�d	�蚭Xt�����>y֝b�͗�e�T!�h�I������G*�p�h�U� ��<�$_n�t���m�
d�V�I�2H�����O�Ab��IL��˔ !ς9��5Io܄RQ�@�W�j�4�0F��H���M�I0�hB%F0~�s���yO�L�T��$Qn�A!>��M���d�'���2�#9�P��oV�4`B ��+��)��	��^�vxCFD 朁B�!=�@�����0hR,`��/�j����%qLVIs���%#����KF�:��'GHi�L�'E�e�sA[�}�)Y� �I�ʼ�d۶8��\C���dh͛nO�M���x�)At L�؜�V��6��8tN�?�aN�C�d�T�ƫ�;wM�<�cO�C�d�T�ƫ�;wM�<�cO�C�d�W����2}F��݁��i��"X�SGG����߁��`��/Z�QNO����׈��n��!U�]IM����׈��=o$��hA�(DLPB?�%���=o$��hA�(DLPB?�$���:g.��eL�"LKUA=� ���6b܃!��k��-$*��P�Ҋ+��c��#-$�u�S�Ӊ+��c�� )!�r�W�ш+�n��jt�,"$3E? 9�]2n��l|�&)(<H3>�^0m��`x�#/(;B74�P>c����ZM#I�R*���a��ד�#��[M#I�P(���e��ߛ�+��]N!I�P(���e��ߛ�+��]�_��g�t����_B�������Z��d�p��YB�������R��j�z��QL������Z���'�Gn���f܉��Yʹ���-�Mg���bވ��Yʹ���-�Mg���bވ��[ɼ���"�A����8�z��w�蝧[������1�p��u�ꐮS����:�r��t�랭U�����Uk"R1�T�����޵Wi#S1�T�����ݰPc(^;�S���۲_c)T�{����!��ȶ��������Y�w����"��̰�����[�q����+��ǹ����ɂ��^�s��N=ӱ	٘+О�`k�%	�h��O>ַВ ܕ�ic�#�j��M9նѐ#ؙ�el�/�e��B6�s�X6���m�$�g��yf�r�T9���e�-�n��wk�x�S<���g�(�k��ti�x�S/3P�y�fF$PпfLp&,3Q�y�gI*]ܰ kL}($ <^�w�nE"QвdGz. 9�z$��aj84�O�_�O7���t+��im=7�L�Z�H0����w)�im=7�L�Y�N8���|#w@As�m���Z���K��#�yOO|�`���W���Dq��!�tDHz�`���P���F|��$�zN@~�L-w}es���_����K+s~gs���_���	�F&~um{���_��� ��N��^Q��!����^�����N�\R�� ����_�����K��QQ�� ����Q�����I��/E��C��b���'^�<�ܾ-F��K��m��� [�>�ܾ/E��B��e���-W�6�׵%Lژ3��~���U�g�>�$�>��v���	σ^�j�>�)�8��u��� ňR�`�6�,�9�����s��>k�m�X�� ���s��;l�d�S��s ���y��<k�b�R��}���vP*CD����M�U��ϚmJ\%CF����O�R��ė`GV-DC����O�R����hM	["IO�������"��-���Q"�������*��(���Q  �������'��(
���Z,�����Bf��61m�������Ol��32o��������E a��88g�������L7g�j��۔������y�T:e�o��Ԛ������|�\2k�o��ܑ������|�]0o���\J�:�o���J �	�]��Y
B�0�c���L��]��\H�?�g���G��X��Z�o\�3k��i�z�8)��ڥV?�dW�;b��i�w�4-��ۥW<�fU�8g��`�|�?!��ҭQ9�gU��Q(t����;�6��(��P(t����>��5��#��Y.q����6��1��'��X"~�f�Z�;�k���9LN-J!�h�Y�>�i��	�2AC&@(�o�]�?�i��	�2C@ G �g�U�/���rV�ߒ��<J~~�#�u��wS�ٚ��4Bv{�!�t��yZ�֚��:L|q	�%�siED��Q�[ٛ[��u����U�dIN��W�Xۛ[��u����T�gMK��P�^ޟX��u����U�fKM�z�޶�N��p�E��~P�24s�ݴ�A��}�N��~]�<;}�޴�K��}�K��t[�?9~�֣�����{�<p�%z\�h������~�9t�'{\�h������~�:w�"|Y�o���^kփ]�5X��ԶO@*��eSb؎T�7X��հKG!��lTgیQ�?Q��
޺BO'��mTgی���x�õZ덽�W�c«���z�Ʋ^�Q�dƮ���r�ȼU僵�]�fģ�/�'�1m)
��$dQ�
n�'�/�4n
+��,m[�f�"�-�4n
+��,mZ� b�'�(E����y�7~@3��{x�|��G󹘱q�=uN;��v{���F񼕾s�;uH9��ys�w��H���82�T "0u0��?���v*�
38�R!1u0��?���v*�0<�U&7p4��>���w(�40Ｅ�	D�S'��C�-�3E�Ӄ���K�R%��C�*�6I�ދ���D�Z/��C�'�=L�ډ��� L���wy.+4�
�gW�n������t})#<��`Q�l������qq$ 8� �oQ�i������{~7�.uzK��HC���U���p<�#utE��AI���Z���t?�&r|O��ND���]���t?�&�2�a^}*�F�7S�M!8�#�0�f]p'�B�0R�M!8�!�9�nQr%�H�;\�F$>�# �52*9Dn׵gO.��>�44ٽ2)?GlַdH&��3�9?ӵ5,<GlַdH&��0�?7ڿ> 7���c��k����ޱ��������l��d����ܵ��������g��k����ս��������h�⾠�c�醡{A_�ɭ���跨�f�膡{A_�ɭ���ལ�k�㌫qKU�����
�⼥sK0K4���J�|?I�����tO3F9���C�u5@�����}C<I6���M�|>D�����~F;A���m�wx�/¥|�H�ۜ���h�{u�#ȩp�D�ћ���e�|t�&ʭu�C�Ж���e���H���w2)�����G���: 	�����B���r7,�����f��j|���L�~��'g��i��my�����M�~��'a��k��av�����K�x��*m��a�l�'���oM�d���b#�'�϶�&���oO�a���i.�*�ž�#���oO�a���k-�-�ϲ�,����F��\�+7J��ʱ([�6���G��W�+9H��˳*Z�4���B��S�%:C��ƽ$S�4���|��Eb���9H4����T�w��Md���9H4����W�p��Fi���	3B>���^�z��@���ג�o�F-� &��u���ӕ�h�A/�*��y���ӕ�h�C!�/�
�x���͙�m����y�~1c�{�Μ�g����p�y6d�~x�Ǖ�a����t�r:o�qv�ˑ|>��\�>��-����_{v5��U�0��.����[~u4��W�6��&����Y~u4��={�o��M�؛&�D��	*D:}�j��E�Ҟ$�D�� H7q�f��J�֙%�G�� N0v�d80eoE8�/@�/<��w9Z1:cjF:�/A�*:��q<^28bjF:�/A�*:��w;V:0jb4Q}@�'o��I��*(i�30RA�)n��E��)*h�10TzE�-c��F��##a�:9\pptl��q�dhM�#z1!��Yuqh��p�dhM�#z1!��[vum��w�mbG�*r6$��P{b�n��k�8*^�"ueӔT�L�n��k�?.[�/yaҒQ�H�k��c�1 U�'reՓS�K�i���[�۬��l�Fu����L�[�ٯ��i�@����D�]�Ӥ��k�A}����I�X�y4`7�#��^�:g����v=x4`7�(��T��4o����u<~3d2�+��U��6l����p8}1e28L����g~ LH`*`��3F����a{%IIa(m��
<O����d!JKm'g��2F���7���Y,G�Q��`M�F��4���^)B�P��dH�A�� 1���_)B�P��eJ�E��9 8��E)� #���S�|j��TbB9]��U@���/�0���ǆN,6��uɘ�u�+�H(�űAf�
�x}�H�zH|�(�,S�Xr��>R�t1�!��B�$��'��R��<���,K0�� ߩE��3�a�)) �D;�皝@v�Iɣ�=6��� N����c��>,q�(��"�PR����N7>����K y$<@���0-~qɥ�R�h����$������i�1O>�� n������W\�,���ƈ��	�&g�����(<6�H���?QZ�D�oދ+���#s��aB�����d����rh�>0�\�Q�A>US�hzV/_09ꈑ: J��A�N�R�2jr�,�#nX���50d�U.@�$󆧬|���U��ې���$��.532��o�
n_/bm@���ۘl%��n�5+�V�
�ŭq�������{�B�4+d1ȓ�L�S�#D-�xn$҂`��2��5�e�8F܂�&�033�5V��#���ym29�R��04��P�Ş�E�DZR(��mƎ-f��b���<N���eBj��	�jxJ�!2Č+Np�V���Bà?��6��251���%!]oV�9�R(��!������ܐ�<@�!T 
�"a.�ߵI�L�M���qR�-E��-�� �O����N�"p�
d��*��A��I�kB��$��;[�8�O��0Ynha�U�yCx�lZak�q� F-'܌*�/	�r�<Q&��i����T�r0�7ٞ6+���U�E>_j�{J�3�M���ś������
����Od�9aO��_�V�ځ,�W2��SG�M)4��3$���l5q5�ؼr�μ��Û�:F,�r`����f/"���%]��r�*F>
��Bc�-xN����(݌��!�A//6O��� ^^h"��ϋ'~�� ��Z0{=$p�J=Y9
��f�ƈK���A�7d�����A�i�j��'�V�׻��mS$��$tz�'����	�8�� C�E7m� '��Q��I�m��!A&� ^2m�◟g��-����d�Z܆�x�ωX�HˆK՜�y�-�5����5Hİn�P�)ç(�:��ؤV֘a�f̉�<��McP���w#�mR٦o(�s�[4*b>=�#[��;��^�/D���
�?E�-�ЏԱB��	+u�� ��@>P���K%Eh�ZO>�G-P5R^�,)j
�h���
3oh I�%͐w��H��+2����6aP�PY��<�!p�iQ���7u��� `��	��p��d|�t[G��p���ˁ���D��j>�aN���&l�<�~�Cg%	��������s|�0"5���tT��ҁቒQ8�!
���߃RGX��h�e��Y+�e��o�Q?y3t�����5B��bb�߱E�� k�o -��mK�w�])B"�/t(Ji�u�G�
,�j�`�S��8�"�����QLhy�!n[�#9����+�8,��IEDV��} �#�;�(��"���jq�a�xRC�X���8(ˎk`�YʈOnD����O^�)g���?ys)85�C0b��2�x��������3(�3 +ҤC�/��'�N���X�,���-Ea0��B���y�d�O��rD�S�*PI�nЛ%J�$���ڬFi"���bU���2$�0O\���P��64����A�m=��֋���xrC�j���^�uRL�fL
�N1����ʆ�L:�IK��oĢ,�����d���޶q[ `��K��yǉH�`�d�0��UG��T8S�����>)c@�O��`a�@r�6��L�.
O�)끯_V	y!��R�xʲ풠�0���85 �v�<����ۯH�'�*�g��+c^:4l,`��3�ĉ�uj�P�4N� �����4��M ��ô������&W�L��Wg��|b���!Fָ@�pX��U8|r��w��`f��d�:z0�#���HQ2���J[2�ۀ���4cP���l�ҐHP&�� �!J0MXю�'�$���ӻ~Z0���2�Lӡ΂0
��{�Å��0?���ѹ.�-����*L H�9�&�	�8���!N�ꍂ�E�rn>-�@�A �!���+N'D�qWf�����JE�r2�l��ԓ��C�m/��`���0��x��F5~TekEǊ&�^���\�8��3B��m� D��i~�LÕ�C><'�|��	÷Z��Ж��5_�*ă�"6i�6t�',�j��ι0��LҶI�v�䉋�Oʉ����	@��cGϜ<�\-���]�{o�d�9s���3��0�<�R���#4fRe�)�=#�z�S�B�ϲ(z�Դ;�P�+W���OzuHC�A�%o��3G,�H�С���6 A�&��q���o�$�AA �0��C�/J�F����� pJvW��:ƥ�W�x�� �a|R�ۉc��-�Ǆȓ8����$M��!��B�IXƟ8��
O��QbI��d��Q�Ҧ��ÉZ?5E:��,Ҳ	��<)�E?#�P�ʈ7$!40Zw�ɘߘ' 68JW��ئ��7� /IF-�6d��E��<���ʦ�b���z(�*�G���YI`�,A�6�G@�-rWx@s�*ؗ?j�"�S,|>�J�����u�'�UH�jA�r�P����d��B@)х5�qQǈ�	�p96!K,���j̓-�|�a6K��l �O*3��Jr��##.A���'r�b[r|�QiC��#>����2\�l�)ჭ�Rd��
^�8aR�u��q8��y�l�t(�B�h��\�⩱�0X�r�)঄-&b��b!T(]o�z���m�'����7�@	� b�`�*\d�a��M+*8��(ixh(��iP����)NU�3ぴI�6(۳�U�T1R��T4=5hӴ�18aLјu�ߔ�6=P��@�kT�\0w#�q~��ǀgи���9`�"����$�h4 �mʓ	�l��R�+������?X���hDOЉ�Asª�Y;L�n�@��蠎�5#����e���\���@����8!t��
�U��h�_�i�dE�%d�ʐ
�Q��@�g�Q@D���Q34�&�!�ßz��iW��?s6e��j��z$���GJ�5wJ����'҄?���g�?ғ�5V�4!�)�ä@�/ �!hr�ߦz�qcb��<F찲�^  ���'x�4�1��?ODՋ�OРh@�m� &��U��I�����|����(Mdt0G{���{�\�򎞆~;&�g���Z�H�� V��2�.��Fj����%��]�2��C���
|"�
ÓX���)­9?�������c�x�96j�:ݦ!X6! (hz|˓t�h�&����ݙ5�Y�Xw��� �7h
�I�����H-R�Nͳc��1A�̠���Q��&�z5=9���;*L��(s��*�n>�'6.�i���~�^q�'	�B@öc���̘�j��[u�@y�@@��ħ��8���0�ǐ
!|0B��R"d�6�z�ƛ�bdr��!p�"5Z�.�*��O�� &&Ɨ;�Ԑ��8%m URq�E�1��Y���̋)Mµ��=H83�k9?a7dL�N't�HF׳*��� B=�w��i9�F�$�d��E���@�YtD�#=E���ejU��=H H۞I��%�ȶU8|�zpBդ���Or�X�@�+K
u��=�'U���(d僭}�`�"��*?��'��ѐ5*�Pv��cj�4��\����ژO�eۡ�F0t, �5Ku�EJW �6�nSג>���>�2=@m(y��K�F��)R��4++<�CT��%�:	B�.� #pQ�|b�n1}2͗1A���U�H+0�HQ�R�\��y��ͱY������/b���JqU�dR�O�#m���P�J+"�)� ͧ�ڈ��[	�p<�g��'�`�jDk�|y�KzX�������
� ��׉v�f �k�
$kp��#A���a���u�tB≢T>4ABWM��R_V��R�1
bc���rƏ�|d%R�#Ӥu�����3H<|<4&BT+8�e����m�<Y6m+��0��_3k���Y�l�*e�¸� ���ӧ���$�1.
R��4C�)t��M��4�!���s��L O����k�FK0!�!��Q�;7Vڐ䋬����E~v!�]3,T�۰���"Px!)��|!�d�/d�0i4  :tb�e�/��,V!�d���Ƥ[�L%?Z
����Ƀg!��4G�(�(���oB,��.[6yU!�X�D��5`���1 �7��4�!�d $�DEjC�X;c!t�1��j�!�Z�L��� '�j�r��iѳ�!�]/)B�X��� �M�n�AGe�1�!�P#��y��l�:P��6�!���X!�%����9�3*!��$w
Ȩ���0 |N����Ԉk!�S� �݀u�ێ
h����#!�׎g��@+1oq
�dm��!�Qtpp�I�=~l:�#�A�!�$�F:�ՂH,Am i��#6H�!�Y5)��X�wc
 5Km�׭
1�!�$,����ɡe�6�{4)�u&!���bX�eߔvJ2ѸSI�B.!�dD0F2�m�b̀UC�7hѴ�!��K�mQqW�)L"$̋s	]3h!���"j_�:�Lh9W��Q��$P
�'�����*USF����C1čS�'��ٲ�F
b[�uxtb !:X���'#|�;�B˞ �l�ȴN_!
��	��'���! Ěvt� ��7a<da�'-j��
G6=���0�ʠUj.��
�'e�Dqp�G�Ե��@�qF �	�'����iC,�<�	`HE"a�\9��'��H3�.M�F�la؎	P{�1c�'B�}�c�.0�=��
ÜL����'�*�A1� �Mw�T wH�Gp��`
�'��|��E�&b�q	B���`����'+T���N�(EK�щ�NE�N�(�P�'�Z�0#F�Uj��RDb��',L�c��P�cK��Ѣ�	�|^�s�'�*5j��y�z�+Ɠ3/2�P��']���&�ħ~	�`�aC^��`ȃ�'�8M���)8��Qzw<i�'.&�CwD�QNxT� ��,~2j�	�'���fO
w�6!"�*ޜm�����'�d���Y $N��V�^YL�z�'�85[�*�
~rz�Bc.HP\���'\č�PKP� A�V]�4��'�
�*�eXh�8�U4_d����O��QB+��*^�i��O�~����֣ ��@�V��/8�
�Q����$D9�a�Cth<y�œ14HCJ@{b�X�a=�~R���S Ȕ�CD���1�ҩ؆�1%��	<2@ ��~�y	.�&Np����,6�@�YSF&�OԜ���92�"8�V��?L�	G�ƮQ�9ip킳i���ГA�s`�:�l��((�v���`�/���wEp�I�IX�+� q���7��2�.H/;�2�%Eބ!�� Ц�.!�����p`RҎq�Jg���̶���seTՉv�M`���ϴ���seTՉv�M`���ϴ�����>e��`�P�|�Qf��]����>d��d�W�t�Yn��Y����:c��h�X�{�U`��U����6m����y��A�����( 1�O�����y��A�����(!0�M�����y��A�����(!0�M�����ŞD�F@��rΜ��h5"V����E�BD������j8p,V��ϔM�LK��qΟ��b?u+^��ĜF���@�#~Xw,�t�����B�#~Xw,�t�����B�#~Xw/�rƢ� ���J���p�>���2�?VF�� ��H���{�7���0�6^M����B���u�>���<�1\L����B�183���6Ɠ���"f5/=�183���6Ɠ���"f4-9�60:����=̛��� e0(5�:5>����!�Wu����$��9����)�]z����(��:����)�\x ����/��>��� 6���4V�b�/��v�� 0���?Z�m�#��s��<���9Z�j�'��y��/��G(xh���4\�� (.ێ:-��F(xh���6^��&/&ӆ2%��B+zh���6^��&/&ӆ2%��B����i�{�U��LP/�͍ߑ����j��X��JP)�ǎߒ󧊓d�u�X��B^ �ăМ������sU���{��E���	~��T��y_���~��D���	~��T��y_���~��D��}�y��X��tS�m�F��4��n��r��W�m�O��=��l��z��Z� c�D��:��m��|��_�e����G�!���2{�U�B�ӑ���F�!���2{�U�B�Д���M�,���:|�Q�C	�֖���L%��|����:�j�}��?��\�(��}����:�h�|��;��S�*��{����3�c�u��6��[�/��{�}�L�1 ��*��^�G��S��|�I�9)��!��V�A��Q��~�J�9(��-��X�O��[��u�D�=���S���E�)*���?���[���L�&w$�͈7���Y���I�#s'�̈7���;�ū�q.���.��0m齆�:�Ĩ�q.���#��=o鿂�<�­� ���/��2f㵊�1��:�^�('�����<c��|/D�3�Q�"/�����8f��{(B�7�S�"/�����9e��s!H�;�Y�2}���$�a�٨2����6�=|���!�d
�ѣ<����7�6w���.�k�Ѧ>����3�<|��|RaX��t�Z��o
�NW�6�tZi_��w�Z��o
�NU�3�|PbR��|�]��m
�NW�4�wYjmY�܋V��a�1�ǲ���fY�މT��m�;�ʳǨ�m\�ӋW��o�:�Ž̡�i^s����d �@�B�(uܸ	s����h-�M�H�/pߺ	s����`%�H�H�"|Կq���\L#�������������]B+�������������[F(��������	�����[F��:����)"��A'�`���:���� +��D#�a�����9����&-��K-�o������О�o'F\���g1���0{�ɡߞ�j B_���b6�=v�«י�i"B_���b6�:~�Φؔ�objw�I�|cO[�v���hgd~�N�~`K_�y���bllp�L�y	fJ]�s���bbcfT�N��S 
k+R�/�M�k[�B��P
k+R�/�N�lS�I�� Z
n(P�/�M�kY�G�CB��"jj�B4x�
t؆��CG��*ed�@0|�
r݌��LI�� %mo�L=r�rݎ��IN�tw�e�s!e��$�n��ͳ�t�ut�c�z+n��.�f��β�t�tw�e�p$b��/�c��ǻ�q�ws�q�xΨ�x�24Aa� %�kr�sơ�x�?>Me�%�hu�qŤ�q�42Fi�-�mv�qA�f�����~�!�����"C�f�����x�-�����,H�`�����p�#�����!I�lɲ�&\G�OW=Dd�Nf#���!YE�LR5Oi�Cl*���#XE�LR5Ok�Gk"����C��Wp�(�+a���0��M��Pu�-�"j��8��@��]{�#�-e���2��J�/m�@s��b�w�Q�^�Q?F"a�Gu��`�w�Q�^�Q?G!e�@r��e�t�P�^�Q?F c�/��A�bN8����=��}��&��A�bC5����0��s��( ��B�gD5����9��v��+��;����+��c%��+�����;����/��f ��(�����;����.��f ��,�����3��3/�c�#Wb����̼��:!�n�#Un����ŵ��?"�h�*_e��������?"�v�;`z��߬��	QN�m���v�;`{��ګ��UK�j���q�2jp��ԥ��YG�h���}�6z ��X�<��O݅j��(���r/��_�?��K؂b��"���w+��_�?��K؂b��#���r.���Q[��cM^Qx�5uʝ0��VZ��kDT_v�8vΞ2��T_��iFRYt�7~Ö=
��XR�s�Z�Z3��(U �˾<z��x�S�_0��(U �˾<z��{�V�X7��,W!�˾=x���Z���r�{P�?~/��=CW~ɜ��}�zQ�>~.��1LZv����r�uY�<~,��4I^tÖ��z<hQA~��\��ۤ/��)�<jUGyȇT��ݠ,��+�=mYHt˃W��ݡ*��#�1e�u<���w9W�(��垩��~6���y7^�"��ꓭ��}4���q=S�/��햮��}4����C�D��8���&,"H\����A�F��5���'/"H\����H�H��7���)!)MZ����DQ�n��p%���D�=C���Q�h��r$��	�N�0N���V�k��r$��	�N�3K���]�`�9��|KE�p��ל���)��8��sDJ���ڝ���.���4��xHG�p��Ӗ���%���9��w�s���ox�Fǁ�M.�Etv�y���nx�Fǁ�M.�Gws�q���er�L͋�E(�Aqq�s�7761
WZ۴N{�����B�g035<TQѽGr����	�K�o9?:3[_߳O{����	�K�m::=;��>�b�{xs�q*�E��5C��;�j�vw~�{&�I��?D��6�k�wsy�y"�O��>I��63n�X���v�sW`H���O:d�W���~�{^oE���L:d�R���s�vReM���N:d��f��tc��@��5��4k���j��qf��M��5��5k���k��~i��M�
�5��7f�	��a������*/�i;[Ň0H�������+/�j>\͍;E�������+/�j>\͍9F�������3R�@5h~8M*��R�w�4R�C2d~6O+��S�u�7V�D7ip5D#��Z�u�4R�x�9��A�6U)��u��@�r�1��B�6U)��u��E�z�:��O�<_#��}���K��<H�q���6j�x�%1�	�zOH�p����1m�z�*3��wCG�����1n�t�)4��wBE�z�~@$�ϙQ�����'^���J~A'�ɑX���
��/Y��OyH.�\�����(S���@wH"�R~3���T�$࿥����y�Xu8���
Z�'伡����}�[t8���\�/촩�����[t8�k}Tj��6�!���{1ӳ ���l{Qo��>�)���{1ӱ���aw^c��1�,���{2Ѳ���fpYa;D4��T q���؉�5��2N2��V p���ݏ�2��1L3��V p���ݏ�1��9D;���"&���Lx���kI�^Ҩ��!$���Bu���hK�^ܪ��'!���	Lv���bB�W١��/+ve�!�1��NWф:r�/襕s`�"�3��NWф:r�/褗pd�$�4��F^ێ0{�*ﭜyj�+ަ'y���^�5Ś�U�RѦ'y���T�:ɞ�S�Vԣ.r����Z�3�R�U֡/p P,r�V�Na�yRq�=�-�&�'?d9�D�&�����Q�n�\4JdW�Ji�aj�	9� 5�v�"F=z��Vi�<I�R�b�I�i�0%
��O���$hԪ�0�6�!�t�����M�D�:) "l�":@,G�o�R��#�;H\i��ƍ���v�T�8z^Đ��;j�l��Zk�X��G�;JZm���ͅy���l�8{|%�c�\�ȭ;A�ŇU�\HR�+V�?%�5x*���^xH�H�%f�l9�B����ɊJ�r�B���>��dN O�lY��=.N4��aO�H��dj�i��ݻdR2?��D��:�ڵ�d��<�tl�=Ì�V' W �e�3e���S,�?e�@Q:A���0}�t�ݓ-����0wA��1&�_23�н����h$jD��(�6����ܹW����b�%>�B�1cL��ƵSg�AX�\��4��1k���SƘ:v�����$h������!��-��k��Y
 ��z��p� :��l�HҴ��o�Cj�k�L`�O��GAe�v�֥%�ݐl4l�����j�lm*�H�(�Bx�fO��BJI���W$'������6iB��`e9ov�������لd�/S>����95P���a�K���p�Q�M41dp�;LJ��2�M?�œ�%T�t��	pAe�75K
%Ӥ�Y�~WVqGm߁\P;c�0H2���WU����`�&��u���ӂ2��X����90<򥹶`U�w(h��Ix��d��iXu����5��T����63�� Tr"h��[�=(��`v���`%ʴ�Ѝ��R����S��b���O`��D���`$c��`�\�i*����+>�{��4V�.yY�%#s��9UU^][u�SSSzBw���BDS�S[N}%��QYj5:��T�h�@�I Q�9k�Eϗg��ɏU�
PAE��0W�\A6��U�Q?���)ܩX����&�2Pޞ�dJ��Y�ح���H��MKƊ�1$�J�J ��R�*1���P�g��1���,��3�f/gq�1��d	�_ 4�X��k��b�i3�8�w+�H�j�P>�		:H�p���`��Ո@�ֿ2ZtI�	6,/t�ѷΝ�h�S3aĕQ�KV����G�F�꽹ª>���޹q8>�� �9�2 '�L�&���C������c����!3�9S�R�l��T��t��\ZR��1pF$*��� S���5i	� � L�u���f3�IB�>Y��ɉF�j(�;.n�պ���@�	�06��p�d��M�&'Y6
t�'@=�0���h��Q�&�L�������"
��4�f�n>u@��bG^�.��Abg
z�D�1"+p���G�&r@�Ƞ�O�N���7I��M�e,�'c8��U�U �Q�ԫ�%\��m��;Z�J��|:�CP:�y�Ҭ �t\Hd��T�d1JV�ʜg�.�rVT}���(w�瓸(w�|"�x�
�'A.,4N�����gVޘ�'�=uH̒��U�{$`1jV�Mz��[�yB��ٺ��ءE��(��Hŉ8��8�e #,
�JĎ�J�R��koY�I;3H*%z"�.1E�MypHʀg�	8wɟ4�0�0̀�7鴜�@BH s���P� kFppA8�I�MUJl��AGFs)U<32���';�8 ���I���q�%,."}��C�#����
A��.�����)(�|{Η�-�a~��{L�(�K��yƺ�QfJ�����n��m�P"o�l��ېk鈴���ģ{ž����O�5�!�J�WX�i��a��v���c��>'<�MIt
J9i�>\I��'{J�[�C�d�p1�t&�G�B`�PAX�F�1Ij�DT  - ���$��R�Y)V����3N'e�I-d�ڥ�"�>�� �4B&��zf�\#B����ȰK+M��"I�;����.�&H��db���ҵ��O�a��J��i��PP��$i�ƕ�ToZ�:�R��f�M�2�|U�6-��L��I�3JT.k��@`c�V�l�н��?�EQ�$ME�R;}���y��'���A@��3�n}8�@^�6KF�T��17� ��R��c$�:@��<#�j@�tQh��4NL�#)*��$$Ȉ�أ�G�����g��OM�'�ó�ݦ=�v�	0g>�ԓ�B#�����l��Ӈ�I8>c���N���)�!���{G�����	-/���Q��ayrY�MZ���DP�b-����eGe��Ȕ��ON�C"I�jX|T��X�I]�����9g&������b���$�U<M��yb��'��DS6�caZ���ɱ1��}
������C��L� 4�	��X5A�"��0�	�a�Ҝ�AC�q��a��

��{�-;$"�Q�Y7B�2�8G����5�V�2$H40H2.�x�'��1Pn�6A��5a����s$�=���24��0�兾G��JO��C�f%3�mL�YZ�[d!��C�Th4HW�0��,B�D�A����!?"(P�c�T<X�Ĉ�J������XR}����'At���ަ%	Th�i"��'��E�LH�D�����4@,�q���>���F.�?]3�b��;���nFB�'C`躢f+|`�"�?@Z,��Ư)h����V�S��6'?nms%T�8�x��r+L!.�q{��@�xb	�8���@Cύk�@�Bd�� �0>Q6��#�D��M�:~�F�Pq��M]�����O&���E�t�$e_Gt�H��b�L������̳�(M��a�a&�%b��
��0L�o�~b��o��6S�ih��Y��аD
�}�ҍ_{���S�%�`�X���
A\�3����9$1;��F�f�,l� d���=I��2 �z� FlÅHH�SqY���P��-8\�K�/�0S`h,~6�l8��B����W�Y*6$�#�ƺ��y�=މ!�ǆ��]�U�BM`�e�c�H�jp�QOڷ^/>��6ߦ؉�DJ�'
n|H�)P��,9����ѱ���C�ň�.">1O� .
&4&Q��H��h�4	��ZJ��#m��a�@�Pm���uT:�hO�@���D�A8��盧9-v}H5��U�`����U�c���b&IS��I&D�����Ɣ5F��W���S��T"dj���bT�����R��� _�@�ɰ��H�ΐ9�`���$�+�ƽa���	�xM+��ى9"|����0c(�5 ��%1@'�d���QW"R�I"����\�p<HhZ�r):	�D��R��9q�g��a���y�K'��6�v!��E�-_T0!�,��33h�Qdq�r�#�иr��3����ʗ��D��!�&�W(&�ҕzG*R�z��C��nj����q�6��1gνV�z-Dz»��K���΀{��
�`�Z��W�.'�d�z����r��@@v
�^�$�t�,m�*8�R4�5dV�V��$�H�4m�Ty��狭��lP@K��hO �EM�Ppء��A&%��2@C N��@G#@�_�~�R	&��`
O=E�b�b4�P�	�`4��B�?��O�C�%��͆�/
(��g�� *�2��a�ay�ބ8��`��Ά"�>A�1CJ ��M�Ȋ%��3� @*��[�v����	;5x�dF��v#��0�/�{z���C�׈CaH:��
w������ɶb3{��['Nr��bP#Q�y��YK�Ð�aנA��'�-1	�g(?�i�Y` �'��q
�N���h�'3=�r��6��ѻ,�e�=�S'�i��yz��;��}	�c��,)h��BN[,n�.�ѣj�F4���B⇨(����Ojh�%D�RV�e��M[�0{x��%�Qq���UDU�-�y��� FAz؉��P;r��C���[�x)�aC]�D�y:���pj��8P
Ǐ3���O��1 T:l����!ҧq�� ��8c���ct�� s���'��ٷ�S;�pɑ.��.+7lP��O\�r�Nȣ� �תݺ�|�2����&�4�Q�>!E�>�7�"p�]bӂʃN�`�Ɍ9xK�	����'2%�$�$I �N��|�	 }2$Wd���"���B@� ��y�� 9*P8Ć�	���I�g#��T�4p���Slr��4�%x3�Pp����BJ0x�F?�p<ar��*&ڹ�v/���f�[NX��c����?"�m�6IdEH�e
&wP���#�& �� �Њ �\�B�I�_HB���F**w��h��ϥV�2b��`�O墤A�%"�U�a5�S�o IS�G�Che���@�B�M���z���{G�i8�+�
x���Tʈ+W����g�>E��'u���'d�!�@���=�:�	�'G&�����b$|XW��=`�l���'�V��B�T`N�!�F#n���	�'d�ʲa�2��1�g�V�f��y	�'VD�i�'�H�P�� Siz�	�'��"f�ưYC��p��V�C�'�k�E�qǮh ��	C��hP�'f� 05��S�\x�D҅GI�r�'�)r��Q"����ߧK�\p�
�'$ ����Z�����4��8�'[�9[0��VS��a�(�
�2�{�'��y�j�*`�kGOI�X����'����~���w�!Q\H[�'�fI!�C\!>�I�v���r����'ݘ���05�p;��b�"ڤ�y�D�G�\s&7ZG�k!G	��y͓�>$ )H���J�ǈ��M��C�6�F���N�)-*��T�^-pD�C�I�d:���,�3A0��6 �1KvC�	!JY�P�B��'W�+a�P�L�xC�	�B_J���i�Ĉ��k�$)�XC��	d>~m����|�jHr�ƽh�<C�ɝNPk�Cͮ� ��1�%��C�u��YS�k��{yU�����jC�	�(�4�M0=���@b�HC��pՊA���z����U&,��x�M�7�b�E}"�
�^�i��^wۖ=H�K�t�L���ܣT�\x���t�ֹHO����+o>h�!�/�L#V��g�Pl��jV ��;9���⁕l>���!�1Xf��e��,N(���<�1�ם@K�l0��#}��	7P h��h�2w0$��O�����yb'b��?M"�L�G�Y��Z��S��^�M#�dC��}��y�B���ģq��8��ag&_"|�"p81I|ܓ�0|&S/������p��fE��~f���O��x��ʎ����	�4qTN])kz[�(h*�;i�	,i�8[��U( ��S�ONH�nxLH�B_�I��y��4��I���)�M}����L�/#4aⲈ��U�<i�,O��Dz���ҋ=|���d�|�V�A�3Y��GY����>Dy����`���+	5����T��0|�ԫ"w�hӣc�z 6<�dBx�'~�"=�O%j,ҢG� v�hI��L�p��+F���-{��ue����g�	7E�X�É7Aa�I�7/[X��xCd�-1��b?ac���?�c\%X>�qC�I�9�P���l�<��c_����h�(*�䝶[4��4���\Q\�:b�� bO�m�>)	çj}@���M�CƠq��O�$3.��{��@����Y�x�\��[��� 9��R�'���72�Ib��e�)§ �he�!��-��B��%Ֆ�ΓX؊ ����S�O)Bq�`�F���� �|��x�T�h@S�(��|5��WB� fB�H�j!�v&~�v���<%?� �)ґ���P\p6Z����:"ߢ�X���e�0�����m�\���ڴ(��]�3�9p��ȓ&�H���W�܍��-��yb��0�
�QE�De��<��Sc�e�ȓ]�� �(8�^M�$D��%�,Ԅ�O��d%� G��Dc�ߢi���ȓ��i���ʣy���T
�c>~��ȓ@��A�@l��Ҵ=�X�ȓ>�Ա�T?o�����Av�Lm�ȓO�\��Ԑf�N�I0ㄜ6��J��pϘ'�k�����ȓf~���N�t~���W�!�P��ȓ%�tIS5#�XlZTÌh�ȓIVXx*�nYI���` �E�fԇȓ�@�Q£:����G��l��K��� 5��%-b��IU�|bVQ�ȓ&%�H87�ز�4��6�ؠB�Y��/�]X��T�P*r�k���:��фȓ.m�<0 ����5x@'Z����U�,�7�W�`��`+B�tW5�ȓ��I0WE#�.�#��NQ�l�ȓF6nA�#��
��h��`G8hA�ȓ+ܐ`��C	4�Z���ԑSʈ%��2��	�PlT�q^��*��/���ȓ4�,1��=`�(8� cJ2E6 ��St���޳$.b8����~��ȓ]�I��-M�O� ����ӿ��H�ȓw���kq�I�^��4��)Y2:&"X��N5 �"ŗ�Bb�uz%g�36�ȓ:/��iǪ��M8.���7=w�\�ȓJ����B��,��`�G�0;�����(t��gV�S�H	�AIĔ�$݆ȓ$�`��ch�5K��R�)����ȓ}$v���F�
���'��k��a�ȓ[g�hpc/JU\�
�E|j,4���@�f[�I �(�J�:��d�ȓj:H���!�R�����nӾ8�ȓR;¡:��>�,k`o_�>�ȓVҔA��@�~�����t����ȓ&Q�|��Œ�J��F�Q]�=�ȓP9l1$�Zx�����V�$���&���Z��\�qц�Bp�2-��>4nĹ�m�[���Q1��X�����w
PZ�J� #B�=�܅ȓ/�<Rw�O�h��P�{¤�ȓ"��a��C�V���� \�����WPbT:�������1��V�ȓb�5�Enž=g5�pJ�07bꌅȓp[40�G)&>�d9�����]��4S�����  D
�r��ԲJa��� ��Q�D�nXi�Eh�nj-�ȓ;���
�d�=A�`�:����E�ֹ��+W�E[���V�ȉ$@G!9��ɄȓA0��*gҪR�0i�dP�B��}2�ȳ���D:āU%N �\��p[��"p�_�$�:�9��:V���ȓv|$���ث�|l��^=V_���ȓ,v�P���Ue)��^9w��A��W���*׼D�y�cn@b����ȓ,f�I��߲0*�ӣ��1N� ���	G��q��4H�d+Q�۩o��8�ȓy����ї�� ����#K�>���A�v� �a٦����۟R�ͅ�\|��6UD��iB�@�<�����S�? �8��ȵ����椘�vQx�"O����H�t�VH����5�w"O"Q���8<@�� �Ud���"O�Uy�C�&�:�s�d ���P)�"O�AQ���6�VE�vj�.D��$��"O�-p��ݓem6I�.����%"O�}�s�ΰT���ʊJ�&���"OtE�q�F50	0đ�lA%�XL�"O��0�iQk�ȜZB��|� 0b�"Oj�&�~�\P��'ߟ0�ޔ�"ORm�C�޶X{֐ZVD\��>��"O���V7w��S��6�Dy	�'3�����8 M�@���}I���	�'�rD0�mJ
9���c�� r��A�'`�������!��9v�� ��'�R8I���?�ʙ��;qL���'��""S'6 q#��y7�3�'��4zS���Bt\ �Q G7i�.	2�'¼0��@�q1"�@ѫ��`�����'�.���[�\Y� ��� T�8lh�'oT�j��3~���_�t�:̠	�'��laf�����s-�4o>�l	�'�`"C,B���z�@yG�Dj�'���q�Vm{�HKF˹H~�b�'^~! �T/��D�V���B�C�'�5�$ Y��l�9C�� �.���'dA��+W]`i���@�s����'�|M)����;b1�b�F4[�Z��	�'���tJ�5d�;��+[.�`Q	�'N��A0F��z1���a�X�N���	�'X�	pU� =���I��K?>����	�'�x���SE���̚-)�`	�'#J]��ڵZ׊����7u�U��'��t���⬈bo�Zj�!�
�'':�s%T
Y�� roO 8 9�'��yW"�+@�9�c�`�$}�
�'�R�B���t_ވZ�#�8���'�:�hUMн'����� �4�I	�'s��څ��h�tl�0��gIs�'bF(�H���ɉ�ǘ�yk%y�'�
j3gN�lO�A���udY8�'��!Ys�ΨOTP��)V6l��*�'�J�[�F8�fu9��U�/ԡ��'C�MQ'��.I E�s��QI�'@���K�&�����M��q�b�
�'�Ib5�߃tt��@�e�i�-�
�'�"�C��(+ۀ��&�ڥa߰i�	�'��m��.�k�@|�Dˇ�TGv���'�bIÀ�V<!	�LM�K�j�2�'����D�R L=�VN]	p�D����QQ+՚X?.�!�K��8)��\���p/��b�(P���A�Z����Y�٘d���kМ*��d��;81��({Yh<����H`��
Y�])���U�&i�& ��5%�H�ȓvr>���m"�p�nϭ ��ȓn�Z�����2l>�4h���B�< ��B�Yhp��A��qV	�r�D�ȓ7�Y� .I6�5���64���ȓ1�����E����W�4�~���I"�� UMM�f�v�VF�x~I�ȓ]tX�s`��2C�Ր�Ģ�.y��:��ģ��U*Q��8Q�[3p��	��F�D�3L�Aߠ H��B�7� ��S�? �L(Ջ(���r���((=@�0"O1������yQ�D> ��0�"O�t�ңVr�r��5��i���""O���#)�M\�q"u)F�~�:E�*O��C�g�y1�T#�ُ`�@�
�'�>�2�G!u�������=�[�'l��4�� Q0�,@R�<M��i�'*��)��(X&����@>�y�IA�	�����h���=�yB# ���HU� /�p7aX�y�K[5(�|�QA�?:�Dq6.��y�H�IpfЖ�V����F�$�y��H�'�&���D˚/�.�C��H��yrD��pVj�����	c�̠	�'��ؒW�T eѮa�s� 5	��m�	�'�Fl�B��0h�2г� �R����	�'����K��t,1�`��53�����'m�u������q'#��#����'���8q�OG&�@�� �L��'���2Ą�-:~�a@�̺"g�1�'��x�g�ŗ�8�[�B��+����'H���CD�n�tc޼+<ZP�v"O��YVk�-@�� �V o-��"OJU�&LK�
�|1R�C�r~d=��"OZI:d��	Q�T�[�)�a_�ȉ"O�4�T��9 k$)Q��]�f�,%9"Od��`�Bäእ�G�`�"OlQad�Ôbf��d�	`�x�p"O�<�i�N
T|�ea���1"O�4�gC��G5&���-P��)�"OP�e鄆���jgf��5�BpkQ"O���Ů9�<� &ڟP���g"O 1��1"Z�X7���͋4"Ou�F�M(��ROS�l��"O^��6� �30l��$�(d�W"O��[�"N����$c��`��y;$"Ot�ّ$�Xܸ,)e m�����y��[�	@� Z�`ƕ]@p���y�aĝcjlp!��Z�L�aS����y�ҁF4b�
�f�n���Ï�yR���$�"	#�
S��@��ᅳ�y��[�#��;`H7\#�͡!Q��yB&�(0l�X&c��e�Y��lU!�y�]l�p5U2M��a2 I]�y���an����/^!B�2A�Aڢ�y�+�v��0p�E�t�ZW��;�y���HuYUaE	A��!�v�'�y©�>*)�܁���;�N�C�JW�y��A�hX	:pf�$9H�)���y�S�n�x��ɍx���d�E:�y���8�y��Ƃi����#!��y�N <HA�q�H��\چ8 n���y��3.�x��kL�X-4�g冮�y��6U���C`�Z�`0����y2�A�n���a��]W�(�F��1�yBO)��=k���V����ybX2r��P,̅G�4IS�M��yr�"gd�Av�H;iFB�YS��yb@'�4�) k��+#|1�;�yr��!s��yh�%l�nE���:�y�@_hf���+߃/��tIp���yB�.����!U�U�N���yb�� +�T����(b�	�w�Ԧ�y�ǔ��.)zt�C�_y��R��C�)� � DF�U����_8����d"O��
7�	��N0q(��b|�0"O��",�/s�4,@�@��:��0ȥ"O�ɫ3�D'�@H�5	Z#4��b�"O��v�ύX�jAx���0���:�"O4�X�!\�D|��2�h�i�Ѐ�"O`��a.u���S0I��l���B��M+�O�ĉ�?1�1OV�)&(�#g�Hx�j}��H����=H٣2�Ă}Щ��mF	6T�(ʟ&�	�%l�q�w����b�Vb����3Qs6��I-��jT��	M&p��Q�$	���~�t-��&S��W��x�v��0>tdqKY
N~e��48�l�v����)��O��$d���(!IP%-	�Y��O�#�썐�#�[�I���?qL<y��ԉe�4I0p�ȾC2H�:s�b��զ�3�4�?閺i�b�O3�4P?��W��H�aפ�o�)�O��\����i��y��'�H����ݍR��a �A���4���-�'�D@��Q�͛v� �Ѩ��(ORYe�03B�����.�AH�'�uXT�BEQ���铱��p��t�X� 1șB�{��Z��e�]���ˌ4h���%��vO4���'5�p�2LF�j���A̟���qT�>	&�i�nc��?��3�0�����D<5�b�?�?�iP�$~�,�nx�4�1oU�7��OW �]Tk$�	�2��3���O��d�%w�DD��&�MK����2TeF�a�4]ra�������`!�Xj�ȝ� Q������7�򝐒$�plv��@��~��Q��Ú2ŶM�үѽW&����R,Un�8 �D�*�rbk����up�Z�ϗ�}�Dq�SA������?�������O���3C�2d�в���,w�ݓM�x���9}@��c��>f�z����u�X�W	�M�-O0���e����	~�S�?%l�Dp�%�â� K	�5ځi�>2��Iܟ\Bbߕ~��5�N��@xX���?3�=�G��|�d��rTD��5�I7[���o�_�Y�����Ǘ�3H��H��m�n��U��A5<u��OF"���U�~�`A��842)#H<�4��⟤p޴C>�>-���l[�U�t�P�X�%�k�T��=��-��F�� �#��9B�0���G���x��z��`m�㟔�ٴ�MWaD�r���j�3˰`(CƙfV6��On����\�'	J�z爒�V��pC�79�0+�Y�A�(�
�.*��Hs�N�g���?�rr�J fv��+W�
� dK J���*1.�#m���1;VK�`��	+0��=�<����g�݊"�� �c�kw���R�$4��h�i9�ʓj�J�i>��ēh�f�r ���U�q����3%x�Ey��',���2=��� ��dӎM[��>���i�06-;�4�L�I�>�撇��3��_\z��i�� ���nӶ��D�O��@cj�3	N��A3+��ub�ْV㘐5�,%�Ҧ�ǂ)ʎCTE��U��ā�1�ɼ)�j����@!Y�����Q:,��J�<8sH�����!:n$PօM�KڶQ���i�qO.u �H7{ ��e��]@�	��A�$ �"�x��'�D�I�� '��n����p�d�#|N��`���:$���	%=�\q��H���j�+ғR�Q��i����'�D7m��%?������Nѓc �  ��      �    �  +  �6  �B  �M  �W  �b  �l  �u  ��  f�  ��  :�  ��  �  &�  h�  ��  �  1�  o�  ��  ��  5�  w�  ��  ��  �  ��  { { L" /* : I WR �X /_ oe �f  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���Ex�%*�S��F�N�~e14l&#��0ɠ萑�y�O�:\q�8P�� E*U�æ�y��X���}�'Gӑomr�c5�y�O\)𐥀��̩7�.���-�y)�*{r��ܱ'F6��E?Q��E{*�,������ ��z���_�a"O� I2�ú�]�s��J����6�S�ӡ*�ɒ�wF
�ؐaF�S�B䉵�:TQ�(���*Ċ8:`�C�I6�~���j ;A]��G��+%B�I�FA�ٓ����+��ʷb��C��>@�B9��ϒGA���&a��'��C��;,��#߁y���J��Ǚ= RC�^``±��9:����T���5�B�.5!x=�@�rɔ����X�9��B��N��yr��+H|)�$'�I�B��j�P/bX� �O�4P�B�	���Q%�>���A8�B�_C�yV��<h^|S�瀉,�B�^���XsjL:l>ђ���I�B�	-�X}��i�2۾@B��{K|B�ɩ$�浃���1_�D �d�[�u�6B�	�c6�X���d;���m�3fjB��"p�V$� Z���� 8���� �q0#���U�>�@Ò�&rlQ"O���d�NR�X�aM�+*$y�f"O4EV�m��T�UW	)�`"Ohq�7ߴe�Љ�✚	C�(��"O)��%1�BI��l�_B�q�$"OPp���U�mV̢���ђwJ���yBoƛzt^DAR���	������yb� mǚ�B��O��ҁ&_��~��)�'a�(E�s�'-�p���ϋ@D��FxR�' B\B�g�		,��s(D����	�'N��yV��y�8����aĺhp	�'kZ�)��[�h�`#�� YSʬx�'�Vy2�@K4"��=3e�דd��t��'Φ��tk�`�
�ZC@�=Y�X�	�'| ��'�l�F0{2.|�,0��'a�J!]f��{�k�<KLyǓu~�"<i���b��;"M	.��ء���m�<�v-]k��y��?�����g�IO���O�t��M��rYC��1�ؐ��'-��ڶ�	�d���c)�I�h����~؞LATJ 6��r�H�}7��0\OT��y�N
�lc�,��)V!If��]�y���#L\:�〧|�����J%��'qў�O��,�A$�BP��*�xk"U�'�,�� -������nJ�Qc�'\a�!P�j������*fC5�E��p>iI<�W!��Ջ�L�:2���j�J�<	�_����m��{Mnh:�/F�'�l6�:����>Z�8�Xc ��s������]���:�OVQ3���6q�԰⍗,�^D���iś�/0�)��PU�.4�Y��N3qzw�#D�0��gƃ���F�B�Hp��_k���|��� ��E�����FB0Ec'ۈ��?�'XЌ+�����Ĉ��9�f(j	�'@|�9��W�\'0�"#��G��ʝ'�'��)�;�&�P#bPK�Vm�����H��G2V�h`��C�X���C�.��ȓL�Μ�s���XQ�\Jg&��H	��Z4��QWH1,�Ũ�o�&W�t%�ȓl�9�G��{�	�TeLv]��?��}aҏP�-=�U����]ޭ'��E{��(ش����LF�E�	��y�n�4x� �$B�I�Y��a��y��mc��"EOo��-�6d���y2�Yr��1 ��%\�h��uKQ#�y�CF=c�!�%��YĀ��7����yBV�rpfO1dRe�0�T��yb��OS:�Y1I�.q=,��F���ybe�A}���O�vh�H6���yR���4�ly�C�M�m�f�fO֕�y���$�D�1�۫i��<��ۖ�yRKKDF0@��:N��[sM�y��n�+â�XԽJPg]�0?�.O�Bg+�[I�)&�Ur���x�"O��	�B_�hWz��0���o *�C���7���pKR�I0.yi�^�Y^���"O��Ғ���=���~��Tr�"OU2�oͫI���Qp�Ԥ)n
���"Ob�r�'ǉR�qau�ȍ_h� ඣ:4�R��O����zR�R�d@X��2&$���/��� �n�P4��0�0��sק��B��>e6 �2�#��R������8Q_���p?��N	f�>��vě�us
��tOK�<�e��[S�}�~\�e��`�<� 0��#اV���"�)6 �����d0\O&u A�2�����G��<��誀OB(�� &�����_˾0���D�<�Q�Y1dp��Q%D�3C��f��'L#F�%���,G��ÎYa�y[BE�^��C�ɵN�����B�T�\��mސO�pB��.5��[2��e��2ca3%ZB䉰[�J�Zg-Q5H$F
�c_�#<!1�'7L\b��\k׊�C��SH�z�'g��Bw���
ƚ�c�����A�'֠��Bi��.�4�K�"4P��'4y�%(M���1+��9w�Y��'":���c
KΆ��ң]"Il�����Afyr铆]EdQ��F�TE�s��,j� �L��I�s��! ���U�0��D���|o2����O�� ��
o&���D� "�k�"O��s$��t�Kv��7O$�uA"OҕC� �\m�M�6�Ֆ[�l�"Oth(RkC�&�\a�s�1V��%2O�Fz��I�, �h2�잁o;��c�I
!��]QX��r�
�u��I�a��V��Itx���C�L>1Yr����4�s�%D�ț3ɖ�^�ؙz�΍;3̺t�1�)D��Ac��6���*H9�����G:D��1�ݟfB.�ps��:�r`7D����hY8��H��P�Ls��X�!(D���n�5��0��'f��aZ�(D�0G��W�F]P�N�y��0{E�%D�h𲈆��bł������@*"D��`͞�I`��`� L2�m�!�$D��J0�.��' ��3 4��a!D��a���f`"#��ʵ�P���>D�h��
�;Q��J���j���� D�@{Wj��Y���*��(R����A D�D�B�Va��IW,�y�ǥ0D��ip����\|I��b>-��d��y��ɱ6��{������`��yrh_0�<�W�Y�	3�����yB�-�z�XB�)��(􂛈�yrn���,����)j:y*c�M(�yB�#jڰP5f��q<҉�B���y���mTMs�Bl�̼�����y2�[:H�ȩ�bR�hҞH�Ѐ��yBK�*jpl!�A�)�0��l��y! �K�Ng�iQE∃c��ȓMFz�HF �5��)Q�.	�(^B�ȓ����A
�j�識��R<{i��ȓm;9[c�����Y�!�M�M��Ʉ�:��݂p��2��!�&�c�6���Tn��aHH�%3�ղ�(��rL,�ȓYY��§���0�`Q�"�U)G7�<��:��$S�`F��A�w��y B��ȓ"����4��;B`@�T�F~���\��mS0��c�P{U��_:T�ȓN�b�YS���WiLQ�#	%xn���P�Q*3�Y+x4���N�,!�洆��nx�fn��L�����	?%GZy�ȓ*�nT�f׼#����s�W�]���:�	*e�M�C8��Q�ʛ*QP4�ȓ�<m�W  (e.�ID�){2��ȓ��Q���88���1�/أr����ȓA.ʙ3�"�7XL����B"D��L�ȓ{�N���]�L$��"`�R�#K�p�ȓ	)ʈ9�c�I�T��@F�Rߺ���S�? �1R$e�3�d�� U���"Oa�$bE�>;��Y�z1�HX�"OBy��F��!�(�!a['J�z4�$"Oj�ʡ�m9�6�^�>f�M�v
0D�d�"�ι-D���#6=j�� ���O����O����O��d�O���O�$�OF��6	�+�mC�Eځ1�"��'�Ov�d�O��d�O����O����O>�$�Odq���^s�j�Q��Z#B�A��O����O��d�Or��O@�$�OD�D�O���æ�Np�����x4V�3��O>���O���O���O6�$�O���O��YQ/[!V!���C��Â5���Ol��O��d�O���O����OR���OF��T�ߝ
/�0���U1!�"Q�#!�O����OR�$�O~���OR���O���O`}i��8'�x�s��bN�d�F�OZ�$�O����O��d�O
���O����O(�	b˧B� �sށX� |���O���OR���O��D�O��$�O����Or�A����?�����[V�
e����O��$�OH��O���Ot�$�O���O��i��_C�Zi1�n��`��O���O���O����Ov���O���O����'K�  �*�:�2-���?Y���?���?��?1���?����?)���)��h���d!��"h���?���?����?���?	��?����?��Ɖ�rr�t���2)���0�\�?����?I���?����?a��v��'���Wf>4)a�ß� 隵х�Y�x˓�?a.O1��˓SN����.1������9��G4e8����O��nZʟ�$��
�O�Qo�=4pa�P�S� �R���g��L��4�?q����S)\\��?��ߣ\�0����C~�*�/IN�E$n��$a�A���'��Q� E��ʝ�i�0�y�M��x����ү��7��1OX�?u ���K6��=�"�rK�0�m�d��қ��yӚ�L}���I�|���' �;0�ٍ%,��XD�K���Z�')�]"B���y��ĸ4�i>�I�C��Hɧ���i������K0���Ty�|�D|�dL+�󤇔`f��vN<<a�ոA��-tAx�T)�O�o���M��'��I�N�h�ת�1�n�6�����
b� Q��z0~9�|���y6�9��zdҀ,�+� Y:�H]9���)O�ʓ�?E��'q�d�C��-ޤ�6��o�x�K�'x6͝�
��	,�Ms��O�̱z��O���Z'�P/8s�`��'��7�������/gi�|*��2?�F�ßq$�y���cQ  ��lm�\�$��t	����Ԋ$��	���A-E�����mK�^f��9n�.t��
��%�T�S��9G��e �ڷD����AQ�I�7lW$��-��-qM4��Ч�/k��߽P�X��F�8� ��>V�>�2���V����Ŋ�
p�p�Å�Ѻ"gPY�%ꋜR��`��R7F�v}˳���B��ID��l�ZP�!��:M"��y�,�'.
�! x��䌻4L�pw`ͅw���x���,az�h�G�m3���*�=�&`��Q�%HZ���芣Nϰ�ũ�j��I�Qc�V�|�ܴ�?���r�4�:ՙ�\�\o�aJ%����kC�!�M����?	p���<�cX?}���?�����j�f_}�*���H�#? ��i��}R��'e"�'���O�B�'F�Ӿ4�1�V���dtT�7�N��T�	�4g=,oSq�S�O.�˚'5v��˱���ʙr��ԂWgH6��O\�$�O�ax��<Q)�h����8C�?��1�E�y�$$)_���'���(�� ���O����O ���m�x���[�ny��O覩�	(��<����	�����+�$*^�V%pQ*גv���貋^5�XY�'5H<�k�(����O���O����O���Gڢ��A�t X<���2F�"m���?����?�N>���?qU.з6�b�%�vf-�j�p{������Q~B�'���'���' |{4ޟ����皕V-��&&q�~�(ûi���'w"�|��'vBϜ*����ܴ�n}Y1H �I�<لcg4�Q�T�Iڟ��I�����K�@��Ο�I�/�v���h��X����I�Y���4�?1J>����?�vm�!�H�&��X3膭�}�2�5\�U��y�v���O$���YC����'j�\c�,R�.��x��fz�����4���O��Ċdy>��sӪA" ��B ��R)x�Lр�iA�	:l�Tqi�4���ʟp�-��dR,v�2Mc4(�cb<҆.������'�����m��)*�g≢[�{@�i��hZ�m �7�ȲD���nZ��|���������|�3`K�1�'�u^�E�B�U�Xs��#ս��	ԟ����?c�h���Œ"�O�Đb��4��th۴�?����?a*�zn�����'��I
�o\@9cgGR�.a���eEI�,�듻?��D]�<Q��?��.��e`P���A�
X�M:F-&)��iroAC�O���O����<iP�W�#��ӡ��>_�Hl�r�>u�f�'��p�y��'���'Y�Ʉu:f��e�4 ��@���X�BÞ����3�ē�?����?�.O����O�����ϳ�Լ*7��wU�5��%�3Q�1O��$�O��d�<�WlW���	Ű�f�$�	"N?� �`�2m��I�t��̟l�'���'e������P�ISc��1[l�Ң[�\��ٟ\��Vy�S�n�f���KU(	�+4��Pd�W�n�*(	����!�	���'��'������4i�`�&4����е1�����M����?�(Oȴ�G�p�۟@�s�u�@.D���q� �t�`�r�p˓�?��"D��|���n:� \�Qa�Ȩz�Z��Q���P��Ǹi+剋����ڴ`��S��h����Đ>M8�Ï%��$)�CI�}�v�'�� �/$�)J�g�I>.��sÊ=63&\C�ߤ.��6�@�Ma��m� ������$���|�Q����MH�+I�\n& ���?�&&é;��Iǟ����?c��	�[�\����D�F� 貅�]�s�4,R�4�?����?)�bW�1)���D�'a2��.@<@�(Ͼ[Ӏ(�)Ń=�0��?���"���<����?Q�����$^L*��� �� B�pAq#�i�N(�"O��O����<��G�-6����>�`�b�I �ʛ��'*B� �yb�'4"�'-�I�rvApd�*�d�8�?1��Dk&�����?���?�)O��$�O���D;z~��1M44��"łY�:�1OH���O��ķ<�5����{/���d��<ȹ�B; ����D�I���'��')��ˮ��Hr^�i��)k)M�@v�u@0S�����T�'H�k��b��S��(9t��1�v��O���=�beC��M3���'���\���xH<�����|�#`N�O��ɱ�O��I\y��'�hu�cZ>��I�4��-Z������@<����8�8�}T�D�G�'�Ӻ���1'�$A���>[��qq�HZ}2�'Oa��'R��'�2�Op�i�k���̡���Q�_�P2�c�>�(O �Z��)�)�<8���w����ؚ"��/���ą?���'Z�I�?A�����'p0X&���A��+$�ƈe0$t���>i1��^���O�b���Pе#���F!.����Ճ�x7��O�D�OXhR#C�<�'�?i��~2��BU���Q�()Y3֤q�2b�4�-�ħ�?!��~��M�U��)D�s8i"#����$�|.pʓ�?I��?A�{���\�$�Ъ� K7�\	��4����B���AV��h��ҟ��'��Q�3�N���^������	�N��@�_�$�	ʟ��Iz���?)E�:,�8m����mc�������0:�by~��''�[�h�ɱ]}���'Q4����J	)�źfJ�A�0oZ��,�	���?)��M���5����zG�.@�t	�V�X�f���"�>����?�+O����sӈ�'�?�#�ʏ�0�'��[���6�S6!����'��O���ߏ"M�$�'�xB�iߺ��0`ܔN�j�� �Mc������O�9�%&�|���?)�'8�H�Jqd��T��)W#�� ;E���O>�$�.j�1O��>@�P�DN]b"��1�� "wd��?A��@�?	���?	���(O�Ņ�X����\�rl�`[+|���̟x��,�$�b�b?q�rK�0����L�DO�Q3I~�zq����O����O,�$�����|��L�Ȉ��h�VP��(�Y�MAc�i���2%ݵØ����D��H�#g �	�̥w�܈?8��o�ן��I���ۡ�Fuy�O���'��D�~X�0����2�ݩ�: �<�f# m�O'�'��D�����c锥"(�b�O5���'=@	�DU��Ip�	Q�`�������0Uu&�;�,6��'�D<�®���D�OP���<y�0�H�갃΀%�<#��
X��.�-��d�O �$�O8�`�I>N��`�"����Aj��Υ�x���9�<��?����$�Of�5c�?���
u҈�s+u�P���)zӪ�d�O��d?����\{c�Vǔ6��&��`��:5@k �?�����4�	Vy��'��A!�V>���]�f�a�aT.*Tt���Î/~���Rݴ�?I��'S���M����@������U��@b$6b]��n����'��LR9{���ܟL���?Q�!B��Yk��	�jP:]&�)W/��'Rd?�P��y��n9�DN='�N��Rʘ�̓<���ӟx�4��Ɵ��Iby��O�iݽxso���aS)O�x����g�>��dB�e�h�{�S�[����vM,Z�D�ႋ^�2*��l	����	ß��I����[y�O��L5���M���Tӑ�F ?�46-IWrD������H�LI�&^�T� e�tn!p^���ڴ�?����?!P㘖��4�~���O���[���d�%JHu(托h&4J�y�JF=a������O���8%7����K
|k��s�.��������,%��'ab�'����މq$�I�L�%�𔠱�B9��Ɍd�n�jrH;?a���?�,O����r�Lۂi[HP�׋��s<B���<i���?���'A2g#
���t�V��
vf�n�x5jS�S���$�O����<)��!��L��OI���/cCl(��h��`�%�ݴ�?����?1���'U��+d뉭�M˅�˟+5�`�Ā|��D�Z���	�� �'�b�'���Ɵ`�իD�h`X�2�� �
��TL!�Mc���'�ҮG;����K<I�O˚&9)왇W�~��]ʦa�Ihy��'�b0��U>�Iϟ����5���A5l�Dܩa!��'PU
���}��'#��
������|Q�Ő���*j,Ӡ�&��7��<���E�?����?�����*O�NތJ��#���F4�Sڧ��I�X��!\#/�b�b?-x��*u,n$��狧��5`�|Ӵ�jV��O��d�O.����L��|���[�e{�� `��uC #A�P��2D�i"!p�� ����R��Mc�? x�#ǆ(@��%��(μF��)4�iD��'q�Q�%��i>��	����/b
ݑ���wʮ\+c�A�*�&\��dЗH�ء%>����X�F��Jp�@E�l;�C�e\�Hm���N�iy��'�"�'�qOf��Ҿ)�≛��׆M6��C�]��`���Z@��?i���$�O�Ҧj-Rq��K�* h�ۃ�F������S�$��ߟL�	K��?q����Q &x��H:����B�&���]X~2�'(rV����$g���'W}�Q"�
�(P��a�B��DQn���L����?���`����&��Պe�K�I����-�}άC��>���?1*O��d(0���'�?	¥� beP��l�)U�$�3��S��V�'P�OH�$�<K��d�x��,R¬R�%��rӴb	���M�����D�OJ�!�G�|:���?I��QȀ�q�J�_MxdӴ��7#.�����OVQ����U�1O�S)��!�eH3x��g�A8��듮?�CS��?���?����)O�N�6 &btk4�ќs�A؆�d��	�t�q��+��c�b?�xq]�d��e#!D�C��e�lp�l H`l�O�D�O��D�����|
��M�h�Xc��\�\��P���*9	��i��if�D�������dD,#��`5�\i�U*!&Ɔ�n1lZΟ��������Ŝiy�O���'����c�c,ǀ.w��#�	أ>��<�,V6A�Or��'���&prl�����lͨM���B��f�'2j�ف\�0�I��L�	vܓ`����0l8��&e��F�0��'�բÏK����O\�D�<���j��K�jø%�Ո@力5�����8���O��$�OP�����X�4i��^�H��2o�.K��d�Wj[9>��?Q������O��1�?�"E��R ��P�I�at�5ڴ�vӶ��O���,�Iџt���$;V7��_�{�7l7:�(�K��.�������	uy��'c�D��]>Q�	�/	h�0G�b\,u�FN-oV�ڴ�?ɋ��'�~`�%�ņ�ē�@iJ�B�T�p1c�͕g�qo矌�'ob�GQ��S쟜���?��d��(_���x�%X0b�p,�v��>��'�2�Ā7\��A�y��`!̈H-L�d�՞g�����[�@�ɴV��t��㟤�	�|�cyZwm�	0g��'Te!�AEE:A�EI�O>��V�k$,������Ŷ[��X`�R=z%���-�_j�f#M���'���?I�����'��Ƣ_�8�5i��c�vI)��l�Dh27dY�1O>����~,�ZF@Эd�H����]H���4�?����?�ШE=��4����O@�	&'>ٻ l��Q ��a0�
j`Ƭ��y���[�8��$�O��I51h.�3PB�z88�wJY$&�D��K)OZ�$�O��$'��u��"��.+�	�U��R+�en^�V��P~��'��X���I�YW^$����T� �S���#	*��6FyB�'���'�O�@�G+�!ap)]7	$ �1c��C�K�íyh�Iן��I͟��Iğ���U��M�pKC��J���R$!�Ҍ"A,T ��V�'�2�'4R�'
�ȟ�Uj>	�B���a��߂LD�m3EL��M;�Ă���?��X?�
��8�M���?q�c�4	; ໦��Q�<rS�6�'�B�'��ܟH��EAܓ!:��SBQ�L 0���g�VMmZ̟��I�D��+*j��ٴ�?����?���5���Ǔ4S��5�6��%
�<)�u�i��U�T�I9x�8�Sԟd���<a��s��q�d�Ѭ���ӄ�3RL(ٓ�i�B�'/�e v�i�Z���O~�d�>���O���b�G�D`̚��9t���8oQ}r�''b����'r��'���
�OH�':�K���:I
�E,�&m�@n�t@�Y�4�?I���?��'�����?���_�֍8�o '?dn�Z���?#���R�i�4����'�r�'��P��O�Of��_�9�i�̊'���C M��6��O����O�uHPɁަY�	͟T�I��x�iݍA�E�"� �6Ɔ8B�Ѩ`�'�	(��b�d�I�,�	
������E7,����C�$es��ٴ�?����8{��'Ar�'�"a�~��'��J��M�Jn�h��a��ѩO��0r1O�˓�?1��?!���?q�N^�b����ɓ4j���h��j�6�遺i�"�'DR�'-P����O����X$:��� �Q29����A�C�0*�d�O�$�Oj�D�O��'.'��'�i�"y�j�&*������)-x@
rӮ��Op���OJ��<����>�ͧV��$�SHY�c�b��M0x8a�^����ٟ,�I˟��ɐu6��ݴ�?)��8�jm�$2t�����Ƕp�����i���';�Q���I����Ɵh��<NRI���4ua ���@0Z�n�����I�$�	�\��޴�?����?���\���C�G�f�N9�"ǌ_� ��i"S���Ip,�M�i>7�RP�����G��9�1�b,��X��'�RbФa��7��OT���OR������'(_�]�#�/>a��s���mX��'6r.\!k�R�'��,� ��ԙ~j�n�B�,�׎�.Y8���a����{�4�M����?A���B���?��?�� ���r�.s�����S��f�۪LY��'u�eɜ�������O2�i��\�'E��!wC�+YH�C&Mv�$���O~��W�G�T�n�����͟p��Ο�� Y����e�[ƋBN� 7��O6��^P�S�T�'>��' ���h
�E�*a&�<O�����i���p-<	l�ӟh�	�$��#�����Q0�&:(���R�:x��B�>� +v̓�?Q��?����?�s�  ��E� s����D2���
Э�-S��'KB�'`c�~�-O����#ys@x�
��������[ K�`$1O ���O4�K���O0�$�|:� �^ۛ��?��͘��K��ճpK-gЮ7��O���ON�$�Ov��?)C��|��-��4��A2�nG�H�=���!;뛆�',�e�'�rg�~�r(T�gK��'|"�Fc�e�E�G�x���$�,2��7M�O����Od˓�yBI��|�M���pA����1+ɓh����c�����Od��O�m�p��¦����`���?C���U�n�X�V�r�$���mˠ�Mk������OpXc?���d�<��Iy�H�4d� I�D��C�e
R�`��d�O�������)���L�I�?������W��P��4;��ĭz�zH*�d	����O���W`�OXʓ�Lhϧ��S�0���R4M�����46�J�fx��l�ʟL�	ϟ����?��Iɟ��	4L���y�o!ӄ��bc�;Uة�4'�b=),O���|����'*� HP
A	})Pd+d��<���"!h�:�$�O<��͝W�	m�\��ş4�����	`�L�u2k^��d�r�J���!T��i>E��џ$��9�
=�"��%ؐ�ow�-��4�?�
O�x��'���'{�~
�'x�IĪ[t�	��6��5��O6	ؕ2O����O���O��'�?1ǨA��>m!���e+��9QȈ9��i#"�'L"�'맖�d�O���l �+B8T��*4b���S0O���D�O���O��D�O6�D�O���ONЦ	�&�ߒ	KHU+s"��d2й٦k��M���?���?	���D�Oн��=��L�Q��B�j@Y��,2��L3��CǦ��	ß ��ןx訟bU3��증��ş�#$�=�V`k�ՌK��4���:�M���?������O�U�#8�����|�M@Jd4QqHP/t�`���aӴ�d�O�d�Ox(�s��ۦ-����	�?1`3�h .�s� ?�Z�x�H�M�����O��2p5��$�O��r�;���oV'?�B� ��՝6�č:��Ң�M�,O\���n���꩟N�D�֝�'v�Qs��1etnKਝ�Xd���4�?9��	~����S�'S"����,R���g�R�n2@��`�ݴ�?1���?��'P��'�R�X(k��"� # ��rOD�:�6m5:�$$��S����s��.�qCC-�IM��Y����M���?���#�97�x�'&r�O�ATR	1ؑ3�  S���B�i��'��J�:�i�OD�$�OUa��6���f�
�~K�,����I??�R@�}��'�ɧ5��|�jx��$�*64+�'����Z��J�d�<���?����d�/]d��/U�3N��b�*Ib5�"E�~��?�N>����?�TEׁKۢ@��葈#�Б;�.�9cg������D�O��7�i*m�\��'8X�l(w����l��?��'���'�'���'�\ȝ'w6k��� ���+ƍ^#6m�E��>)��?����򄗕l���$>��O��Dp�n�Y�^y��,��M+��䓮?!�
��|����ɪ��p�ŭ�0@��1�gg^7m�O��<���4F�Ou��O��x��.�v���Њ��R�+7�$�O �d�V���$:�T?�'�5�<Lz� R��L�u�t�f˓T�J� �i1H��?i�'lc�I�@���١ɔ�m�!iM�#o�6��O6�D�6�-��)��b� ��
Ў[��q۰��\�fo�coZ7�O4���Od��k���Ls�8=�xɑF,/L<;`�N��M{����?�M>E���'��x9�d�� n�!�;*̜ܳ�gӦ�$�O����In��>I��~�Ҽ5���qӠ-��	��إ�ē�?Y�ύ:�?�/O��O���38���2#_�;�r�u�	�7��O��g�N���X��D�i���h�'�LTq�@�&U���e�>�2��<�/O�d�O&��<�E���@0��C�@l�J���<fjt��'���OܓO����O�=��� 4<n��Q揋-R>eZ��O�x^���<����?����d���(iͧ-,]��ïw:�L �� ;�,��'��'��'��'J�iV�'���+M] <�G�^���4h�>����?	���$���X�'>�
$���6� �^)v����-�.�M;����?1��:���2����	e�
!a�1A%�1"c��!s�7��O���<	5eÎF��O�R��5Gذ}�@@B#��t�-� �0��'�i��k���'�q��z�kݼ'A0�Sg̜�k����i��	 ����شN*�Sӟp�� �����i�,EscK 4G�d�.L�J��̣۟�i�͟���t�O"�e�Q3*=����HX�m``%��4'*Js�i���'���O��O��Y�X��Q����}����e��Am I����������;�H����5��q�OX�z,
���z@0mZ���ϟD�v�����|�L�|i��Mw6T�b,��[�t�jrNfӘ���O����B=��$>��ן �ɢgT��ӄ�6#}�-趢�-V ��i�O��� -�On���<9����p��R�Y/h�zd��)��5\���d�<0���?����?�*O��r�.]2p�#iW"F#�Yz@�8�%%�l��ԟ`�	F��!rvTi ΜYװ�+T'K<_�4�K��S̓�?Q��?���?������F�%4��г��2pJ��nû�M+��?��䓓?��%ڹ�`K��ɲ�H�
o�12TCI�a`��p���>y��?����d^�r��%%>!0
� t�I��Q�F��i�!�^�@O���i�ҙ|"�'��L����'���JDC�g݌�aI�%4�JM��4�?)�����:p�(&>Q���?�JdA�%<舋g���+6�2�������?���<,�Ex���qP�:]���{E@��Ec�ui��i�ɜX�� �4yz�S�<������,��2E��o��L)�ӧOg���'��m�<�O�������ő1�����ˇ�N��21�i@�A��r� ���OJ����bT&���I�&�(��$kHBR���
�$R��zش`"�Ex��)�O�ezS��-.��:!	��OP�G�6��O��d�O�ܠ(�C�I֟��I^?F��"1��9� Dr����z�c3���<)��?���[��m*Čķ8y���#�[4V6�Qӻi�҈��?�bO���O&�Ok,ɣu��$�bI#u���S�����|c�����I՟���%X7h��g���po��|p���@uyb�'���'��'���'��궩[>qb�b�Ɓ� .D(��WdD��O>��O���<!�"i��)�1t�N [�%	%
���	�E��I��h�	�(�?��-�g���4d�x5(�Ӎ)/��
�Fб����OX���O��$�O��P4��|�i��u" ŏy"lj��H�L��ie2�|��'db��n����O<���gY�[R@)*V|�s�F4#�ʸ��U-q�Y#RDK�
kl�r��V<�ZA���4v������[���B����
a� �2e��N�<!�"�l�����h�h�c(��c�ך.sTTȁ��o~�A�;V�I��@�
L��P'dǞ �h�`鉈d���A1�՗Z��XS%�=�vX�U�t�wjۊ`��h9 ���1�N(	I ��P���*}ᙢl��80\L�p�I	Bh`��ڦ#dq��K2cZ��-dV����<��)���?���? ��l1�"�&��f%��ȡ�C�[�M��sgR�^:0�8��*�nc>MK�Xz�o�s�B䣂.��d)l�v��?3�~�9�j
��d,�BۈTO���H���ɑѦu;A>�"}�r�\�W� �����D�����-�I�F�����|"gC1<x#�d�8��@��\�yr���bJ�%���b��EQc���y"�'`�#=ͧ��z��9�s���t�T�*BM�i�D�b�-��8&�����?q��?�s������O��"k��� P���C���6&]��5�Vp�]��䄦d����I�0�����g�FP�e�I�u5�T�W���(z�N�>o�Bx��Ɇ����LCw��1 M����$��O0��/���'�<$@!ɓ(U��phd-�ڱs�'�I��0$:��VE�$�̬8�y��e�>�Ŀ<��M6Q������*�����Y25��:�L�K������>o���	���ϧ1� MJ`܆	��eBW%C"�M�
`RN$bb�
�=	�\j"ˀU8�@үD��(����45?�oZ�t~Aٷ䍿:UK���u�r���7�r�'��u�(�jFP�|�"ɚKhb�p��	�2"�)3gD� #�c�k��˔B���M�$�qML�q���z ��BL@��?�/Ot��ԂI�e�	�O`xa��'[�H)wA�jc��p�ur�9b�''2G�<�`@P�ᕫ00t�(���O��\���X3H$��*�/�48G(����4`��sl�J�ȸ��P�O�`eY���wt�P9�/ԗ�RN���r��O��%��?���D�{�P1ѩ��e6�`C�*D���I�@6�#p��1m(�f�.O��Ez�Z��1�G��)F\X�T���7��O��d�O�����8�8���Ox�d�O�NbrL�E_�j���A�Tn�ya�K�`[(y��Z|}1�d2�3��˸5z����$� �s��,G`j��X`���k ����|b�ϤF;f��� �d�� `�섆 ���O�`������4>�BN>6� ��F�
$�Ʉ��&@��M7���b�o���<��'��"=ͧ��xR$ �	�>lȲK\�M����V	(D����?a��?�ļ���d�O�'ljD��LԈn�.�
Z�*_��1�h�^P��>B��
�'�<����<%@򯌩J�A'(M{��S�k^���P���\<x"?�CM�	���8�F�` �y��O�|��	%Ӱ?!�7b�}2�dO�D��y��)�P�<�L�	!n��� I���~@���Cf�w��|���,"�6��Ov��ѕ`�X��@L�r?��L��j�X���O,��%C�OP��y>���JN:nV�����j�Z�h�I�\��8��EA�$&A1u%�D�x��71� ���QH�H��*\��� M�}Q�ud.	C����I6=���-��I�)��@U�L���TΜ�5!�$�/D\��"��!j�4��-�3+!�����)�G"�0�px�7(�lan쒕E�b��l��ݴ�?������Н �D��Y"6@�f+���L�rc��B���d�O����N�
�*%.i"P��5��g��^>C��y��m�厱0Q��!gC9}2��Qa~�� ��!�5x��S���X�%!
����Χ*]p<䎃�Zd4��Pꄼi�2��O�x���'���O�� *41�O�V�rL�vB�'w�@f"Oa[��W&H�����M)��Li��'@�"=��J��c�\xr�54ހ��n�-S���'��'l�ҥ���W R�'Z��yGGʞ;��M��.W�Ph T W4Fhl��+�/��u F`�.gdp�bU��(񄖪c��pY�¨#��ERQ��,�1;gOD�33�;R*��"ɤ�����:�$�Z f���,�]�P%�"��xU�<$�8�"�Oq��'�=��d�-z:�ZA�φ>�tA 
�'|��4}T\�kϐ8,4��O�UGz�O��'~��@$ΒG�zU��Ch/�11	Jb�h]D�'c��'�"*nݽ�Iڟ�ͧrPE�iٰ-ƹ�c.Yu.C�P�T��eؚ�X%HCA�*'����3dL�9d�⠲G%8���s��'}�L�hĶX���O 7Jv�����9^��*�O|�	8\��܁�FST�J�L�A�����O�q��ɻ�����ET2a_�V�S� r����)�$Ť �����Q�?�*J�Ɩ�%A1O��m�m�I�WC����4�?��X�P�@����[�d������0��)"��u����ϧi�*��VѾV�)M~�4[$h _�*�N��Q{�<)����O��-Z�-��B�*���p�*t\Z��s��}�c 䞊.V��?yыҟ��4B����'�l��Ɍ�?ݠe9�%�}g�\B�Q���E�S�O�"�"H����"�֌q5�l��'K�7�$Jj��	e ҼTI6�""�Y�g����<1��P�GL���'��]>�B4ɀޟԢ򆗨�@�Jbk
cQ�������(�~�1& �28ӧ��|B� oS8J�,C�-�F�7o�_���?<���=/,$is���^\�K~#���4��~$a�7!}"銋�?�4�|���@�82W��
���E;�y�-��MpܕP�ǌ;�2m�6����0<y�	�}�N��5K�~��X� ӯO����O��Q��K�m�r�D�O��$�O�n��WTj@2��x��5�N�E�
y�,��C�8��L>�։2s�`
�X0_0��(�|� ��V��9d�T�?q��'�R�h3�3,���*�^(a�����I˟��2�Eޟ�>��y�����<#����%��I��M��Z*6���7]�p�(� #��͓�?)�i>��I\y��[���!�F�� ����jD���'���'����,�I�|R�J��u�����8%��B��l�Y�E���>au�0IF���2K��T�#�J����\���U��$i�]�k۔y�i�'��z�D�'�������S��CѡF��?)��@�p@tC 
�iqC��?Ĉ��ȓJɪ� ��-��w&߮t8q�<��i��'��K$!s���d�O��h�Ζm�����Yt^T����OL����Iɟ�Χ:��5�%��� @����?/
٫�̒C��d�2@֜}�(�b��ާב� 󷣟�7˦̺�/3y�~��@�K��mQDH@��H���ʮu����I
E�����䅣{r�
?�ÒAa�p��C/=S@�2t͎X�!���7���Df�"Mܸ���<�!��C���+��)���	�K�;D_��� ��	=������|����)0���Ds��"r���$1��^y,��d�O�]���L	U�4����B��	�A,�|�/��Q��ݰ(��� �oQ>���p��>�3��,f��FK�=���ަ�(��J|Zs s�5"���vF�� 
D��j,�t�v�E���O���9���2d��*���@r�����(r*jQ�&��v	:Mpŏ���ax�d%ғ6 d���^@�r�bFJx��i�2�'��e�� Qjq���'���'K�����g�B�W�vm�4��	)%>����X�q6Nغu6� �䃥�1��'oH�bb�_�B@�)	���/Ov��@���&� �"�y?��JQ�7��O�Y�S�`����V|j��t*IJYTL��/]~̓I]T\�)�3����A���G�Q?d�F�8l�!�d�,:�~1�� �&)>�ÖkȞG����HO��#�ĉ�>��PG�޸0�8���&
�R���=[	��$�O��$�O4Ĭ��?�����4J7B`�e
g�)/$"T�\+h�}�6F�&�1	��hA�W��<0�j5��k8���D
-ze�|��Z�|ҮA��gGC��Cd�,0g��R���f4�lz`�U���dQ[؟��
_�L
�x�e�k> ҡE5�O*�O�-��Ν�q�������m�d}0!�d@��&��QR���M���?$aģ��c��!h�°�����?���/3)���?��O�:0�1#��]�0����\u��EB�|d����R�8��q9%B^3�p<�e �H�<H�GC�O��l��"���؁�E[Q��pǓ�\�j�B2�� �hO�x�V�'�O����ګW��){BNX�|�����"O� ����b�t���][dtYO~@lZ2,o�!!#���:, i;'dݐw� '�lI����M���?�-���[ad�O�%3��	��(�	��mӶ`�O��d܉�z��/m+,�
��9�98�O��� >�RbG3N��
D��?uز�'۠�8Ȓ)N�j� T;R�hٕ�y��c�[&V8,ɭ;+�p����3_97g@2*芙�O�2�'�ғO����`�2#�舠���0����3"O|X�nϖ4�*h���,C�Hh��J"��|"D鉓S�x�rb���Q?���B�_�PҺy1�4�?9��?ٶ-35(�B���?����?ͻ������ yQ����B��L.9����N�:!:� J��+��OV���3G��<�1B�2 R=��@��=m�j��5$F��Xp%�+w`�	� �ѣTIL�}r��]7lz�I_�p��O&+�9�eA�/iW��@�4"ݛ��'�n]P����$�O.e���2s#�[���X0����D74�8�]��y���9n�y�s̙+Y��ɒ�HOZy���O�ʓ�4\���
r���Q-q\Z�P�H�,U���?a��?!��h���O��S���8�ءREakp�X�Y�|ar��c+n����-67.���L�H�'sP�m@~S)K�Ę�9��4�V� �e��IW$R�D%N� A* �]A�ȅ�N�N$�)�=�'ƴ'��r'�^�8W:�`��_p]�ɫ��?9�$�xg\1����S�¤a��f��&��#��,�(s�ٟq2�xAc�,�	 �M�J>�bE.H�V�'^ҍ��y�a!C�D_2D��T�B!<�2�'�����'"?���@�\�}]�I��'O:,��}��]�{���$�<	�ZГd'ڐV�F~�i<u8��W&���XıcO��Sj,i2mT�eB^�т#R�u$)8&���FY�5��CܓS����ə�ē&M6����c��bf�)c�͇�v	�\����7cr�J�&ؾI�X���	��f��6%M���M���P7��1dG�'��!�7�fӄ�$�O�ʧG%V[��n�+e�6|�P�#�H�:V��B��Ov�/�@����b�J0dίL�D�O�SZ׀�X�nmp�b��3���H��e��?GxE�F&J�{��(�"A�n2h5"Bᔅ�~�I�>ⴜ��͜�@Ĳ������99��$�O��d�ON�?=�I���t�P	f5�*�	ʟd��I;T�`���JT9`T���2����c�'l|R'�����`��;_�,���fӰ�$�Ob�$�4�F�v.�O4���O��4�5[��J+}*�h�`��Āታ	֪E�j۬O�AE
χ]�1��'y��i��F8%�(�ʀA%�\�d� �� nZ<Ji�ڗ ��)�q���s�O�l��BS�)�X�:��^�b�$�� ��f�`�,���|��lً"��G��� �U~�E��5�dL�u�J��$` �$�^��'k�"=ͧ��~���R��_�E<�q����h��p$�<cxD�R���?���?�׻����O4� �|��KL�k�x�-�7-s&q�⃭+�����N�3�&���aR>A�|Á�	�+�D��'�+FrdX7��+j���fD��u2X"�J�]��]�a�ݕ[''�6d�#&�	1.ح�g`�)�����*e\��(�O0�������&
-rq	���9gS�C�	�hz�$�@B]1lF�ku�.@Ьc�$�ڴ��;���0�i�R�'������n������{�l}�V�'�"�B����'��	ٜ'6(Ph��M��}��iD7��@�#m�7B���(W	܎ ���@��M�'`�s�o��y����7��.K�X��n��:y��H��W/E�>�s⟦���bش'ݖ4s�{�ʓ�?���x���AV�h+�ba�6�*V��
�ye"i`\,�ea�SӠ�r�����x�`�p���ц���PTIнXt��3'7����H:�l�쟸�	r����
?�"i��@%;�ے;��if��7�"�'�6���/��vx�=��T������OK�(�Z�ӣ+�mLDAAA;����>	p�!vt:���k3Kt1H1뇈(�@����=L��!=�Z�;�-�W>Ra���Ӻqv��'�t����F�ɧ�Oq�xZ���@@@�N�P�'�RQ8�N��xZj)"OAY�lĀ���D:��!}Ġ�:Q�Gs'B�4iS �M{���?Y�yZ�j%� �?����?�Ӽ��N;7�~LIB����"�S'и%0��`iʜ ����2*�&G�@�����?}bE��%�(�Z�aÞ$�1A�M�rv<8Q���f9�L`ޕbʒ@y'b��Ӡ�p��9�� ���!B�@J2�E$m�tɠ2�Kp�%o�|���|��U� y�.�)u��ɴgK��y��Ȗp˘��֨�qh��m
/��D�b�����|�+��$Л����b�.9���Ρ�P\��*_�',b�'�&֝ğ��	�|z��J2M�4�CH7 ��4�eg�qx����K\����~��tsf�iD���١r��g#����Лg �6$�Z�*�>LO��30��n�^MpA��f�\1�H��I�r�5�Op���Ӂ8p��@\>O�b�"O� P1PG��jk�X{�ޘ:���g�T!�i�йi�"�'fV��HH03�@�7���P�1�'���3y��'S�+"kl���F�������	�x�.YPD�:.P�Ţ�!�+��:�,�H�'m
����[+Y�)�eYw�����k����/GmM�Cb�;:"h�*��5g]�<�=�6���bK<)�
�� n�	��G�,��$�)J_�<9"iS�|bV��b-��k��
f<�նiM�q��G�qr,���j<\����|�êB,^6��O��d�|��?�D�y�xh��D(jФ�H���?��9�4��Ș����lÚO69�a��/'��"�"}R'���O��b�0#^ &(Ë.��X6�>yPLPǟ�I>�ʖ��, �,җ.��PX�E���E�<��T.t�T��,��4U�t�z�\�����pܩyu�գ~p�,�W�[JDmZ����֟ 
1�H�J�&����4�	���ҷ�K�&6�Ab� \�1|�[�c/�
+]���Ę�M��z�� �A�X�!qO��jB�'I|<��a� 3�P1�IN�Ț���'��N����L>bGH%_�BX
B/Y=@ԕ�eIr�<)5���,�ڡ eC�6`�q�'M�o~�%9�S�O�� ��v�)#F��	*
��-�<+.�A��'@��'�"���;��?�O�8�WI�5\��2Jƚ���1BO�K��}ꆭ\�ϼ,YcLԀ��#?�Vh^ M�x�Ҥ�Q�g�L( p
EU��\H��V�Y� �{g�
:Ϛ�6I@M����o<�I�^��DPg��s�Җ��?L�4ڧO�O�$���/>�Ukʪp=��;0�G��C�	�[�.q�%үXC���T#�Kіc�\۴�� C��:"�iOR�'�"5[b�P\��H�u�_�f�8�	��'�b/��_�"�'��I�j�r�`W��P��	�R�t4�wkن>)ԁ�M'{����S�$��!�.��I2D6�X��@�i���¥ɓ-@���[)=2�+�ė:\n�أ��6`���rN�"!�_�~�<�rÅ	+\���MX�q!�d�ͦ	����8	$��8��;r�՚��-�	YO���ܴ�?I����)��;`�DM�1����	�.H�P��FS�R�����OP���٬���A�B�#� �3/H����Y>-{��.���'�R�-Kw9}��B�/|LZJ)S�@%�De�/��K�GJ�_�
��'?o������0�p�Q1"���O�����'A֓O����� sJ�u��f[�Rjz�C&"O�@yWG�9 ���F^_4�)Q�'��#=y �H�u�,�#&%�vۖ������1��'���'k�Q3�R���'����yG���;X��Cg[� H�lµY�� ��H���G�2e�c>�O @�� ���F�R����3��L:`���@\��㌀�Jbq��'�,+��o<F4Ғ��Gl$x��!�D�Gh��L>�!����3Wm��
�(��@*�x�<)Ԁ��Ȁ�ơB�KYt��gCGq~�b<�S�OKbM�f.W?@C�=����N�(A����H���j$�'�b�';bw�%�	��XΧT����t�< x.��~����D2o�:�x�oJ� ���$N��:E~�	[<b�����ηf�0���DA$L�0,�����cIN�cU)O9_/�D�Պ�P�@����d�e ���煬W���7�� +AM�v�
ȟ8���`�d��!<E@�@HB�|G*���v.�0�h�5�@���\]����<9R�i��'< =r�h�b�D�O��7g�9����$�Ig�q�2��O����a��d�O����`�h��L�U�����/�M ��0 ��15��A@�<�)��g����O1�R.�1:~D�b+�
�z �-C�����BA�4�{��'j��:�(F-Y�鉏{b#���y��xG��f�(�xf�C u���3Ț�y2��X?lY G�
ju~y�n�9�x�,r�`��TO֟j��R�KQ�tI����&6���?��l��h��L���1��hԮ1i�Y��.	�[�:p����/���'���&�ì.N1�.Z5	����\r(��Ij�4?�E��,K_��2�>��J�X�r@y� �,����u!/�뎘?P�IpB�f��
,Vh$�%+U��l��é8}��V��?��y���D��;mIW$G	@,�0�eI��y��׀(r�`3	_"Ph��ɋ*�ў�S#�HO:�id�F�L��k��$��h�@�Aߦ��Iџ�ɍ%���m�ϟ���՟��i�a�t��Q�|�)���p�"p$EI/^�(�8Vm�0_�UA֮�A=Ld�|2��>A&��6By�7"�
����S�H�P ��\X��jQ�@�m;�A�1�>�M{�`d�A� a�,$0�A8u)�&TT��5j����WP��)�3�[�|u��q	�!b�1��(h�'ޘ$����
n��piwH-����'��`2��|2L>� @�������M��oZ]�'�ۓ��2�On�D�O���Һ���?ќO��;��� s@�Dj�CD8 {�����S^�T"?QHDC�A�xQ�#?����lM��{�
V
2�q�2.V�ց����U�Xm9�GV�-��){�)S����wܓ_ly�c]�Q�����|u�YcS�t�.�n؟$�'&R��/~����MN����TV>]G!�^�/��E�KH�{p0JIS&1O��mZҟԕ'��`�pMnӆ�d�O$�B��1B��5B%Ƌ�-a�y&+�O8��zo����O2��u�F!�&�1a�E%)
�(�X�`��N�,���,M�
�,C�g���O���'��uf����2v2��2G ر���^�iu*��v�U�+��!{'�;Q/,� �{�	���?	B�x�ȓ�3Ⱦ]�qI�>���Y����y��g�NX����;d����x�h�z\��:{�<@JS��/L�vYq��'�S��y"�YdT�ڤ
��O��;Geբ�y"C� J�H,�Dk
%L���ab@�yR�0J�RQBu��9�r�0f�O#�y��-4���eO�e�� z����y�FUbf��1da�
e�ح0�J��y�OE"��{&��V�2�sa޷�y��_1k�:9	3#®�VY�b�-�y�o��Q�N����>|k�a�e���y��H�?��q�6GΦt�ڔc��y�-#3�2yR4#Оx�.��`
�y�T�a�P�@��B"5؄b�Bʑ�y#%/)����)޵b�j��y�׵etR5������Œ��y�d7~]B	2��6��D���Pyr��9z�,�!V�I�uA��;OM{�<�� x��kT�\�-UY��\@�<Q��ӟ�2�X�(�B������y�<�t@�C9(��T"޶��0�`�Y|�<��
�QRȖ�s��}�ufNo�<I���{G�y�GU�`�z�*B�<��^�a�\�1�Bߓ0��q:
R�<y��˹�z�A�e�[}�QJt�RS�<a���f4ya��3m@���@��e�<i�b#�5J�>e�  �e�<i�a����]Z��D5iV�swd�<q�Fs����7B�QF�����E�<)�O�.	\��� +ۂG�4̉ӣQ[�<P��z��:l?Q碜i���_�<�$��;T���5k�<φ��ELX�<�E [�Q�H�å��7&zHk��V�<i����,���2~؞|pB�I�<�'��KR�`�)Hrl�v:$B�X�ؤ�Ѓ�%�Z�{��}�TB�I�<���#牗a�"����
rk�C�ɨx�J��e�_u�`Av��k���=+.�#4"Δr����)|�B�{��ȺSX�:t�	+�1�S"Ğ7l��9�Չ׺7�%>ʨ0��J	2Yj�öfȫ!��z3�Z�|�Sg��r���p�eݰ���I,�|yð�T#8�vi�u�\c�ʓ�ء��3�P���^0�GyR�P��n��PhS1� 9B�e�1{������F)J�pw��F�S�@��~����+�'�f5����ff�k���F~es�dF3_?<<3dn�[8�;u�ACƬt���4�Љp��ʑW�1f�B��H���Wj,�=��w�|��`ʒ�y�8��A��U�N���l*���s
N>��`�*�/_�}FמSd�:��P�"��'9���B����!��P�t�5MV�S:�&�V3:�2�F��	~��[���	)��Fx"Ɋ-5d�U����<;�|��⟋S�,�S�bV����#@F����bÀ��\�r�) ,�a%;F�D��+\#4�H�$+-ʓ�t,P��M�t߶Hc�f jJ���D�2qε	�a�V����웹^ t-R��]�4_�Ia�n ���U�IH�#��2k��@�E�g~L�[�EO� �
�I�X���F
	ȴ����#B����E;(��ђ�E�-�ހ9  �;��DJ-�����y�gR,4ٸ%L�?M�P�[��ł�0>	�Ɗp�}�5�&?�;��O3��Z�ɱ~���!D����d"#����2���aV<� 8;�8y��I�n�)��ؠ�$�\�Њ��OڐǀČ7Ϊ�G>)�z����QL��9aHL�,��0[��E)3�4���f�/7�D�W�J����E5vk0]�%.C�>ؘ�Fy
� j�vD@?
�H�G���&�n�Q�N 	�����L+��Ijt�<U/j�rLPJH�Cɔ�fg�I�v����U�z�4*N)u'~L�����e`r���q1O��ˉ�D�|���80�	B! �
�A�`Y�-�����##��!�� _��
��� q�,�~�9�ZuQ��#�vف�-L�C�L�)&[�Ӱ�T�'���c�U9m:����ָ()���k٬ƐA���ɺ=�ꍦO�Ä�Q?����?Q=��Xe�?��RgD4 	�@�2�),H�,"�/G���Gx��1��E�i�2���}�"��t#m����9Җ%࣍kZ:B3�����$=)l�x�ҙ~�'����H,�yp��'xD^����E-��R̚�g'�}�A蝪9����,�J��9`���BffY�P�1OX�`u�CF($��'��AB�I?}�>��MX�@��;��:��	,�bF�Cm<a���O�a�$�U2w�=h��|�'Ԁ�u0+�2l��Q�'��;��I��`E~�OQ�<��ɨ+̠� ��-��7�}*q��^��h�)\��9u�̇V�P�#��cL~�íG��u�ƪ�R0]7][J�H���,3IJ�"O�a��Q�i�¤H?IV��Z&$!��ƈ�j̊��`�L�i�`����A��.�[�L}sfh����:��[3a|r��%��٘�癍m��$͐6cP�`���ٔb��+ю���v3�$� )��<Y���ef��SFf�[z,�CE�'�H���hShK̍����"_���Z�S�ֲ�N��d3��y[��Vx}rMe+��0�e�a����M�b�p�@ ���e��y�ΞO���'K.����C�}�i_��g?Y�F�5�(�{S��0�N)H!TL�R͑��J�y�P��6�ƜP�(R�V�ʧ4j�b'��%d�l`K	I�;�b�E��͟X@���d�u�G�On��Ɨ|ch��0RC��y����[y��� �/c�4��3A��~��$R�/[ �b��|��u��<{�P�"�YvNĔa��7���7O�'����'�I<uj=����
V����h\��ŁT�Ƴ9���ba��<, ��k�%��b?%̻_I�{wϔ�s�F����U�XK���'&�)1�Ɍl,��f��Bh�=qU���A_ bR1�bJI�b�Qӭ��<$.3m&���$��?u]��瓞����4΀+YD��3���Lݢ%����Ox���g�#���:�o�DIƋ�|jŪA���(b"j�$q�(88�ϑ,�)U!����C���~J?�~��nZ�fJ�5I&O�j�-B� SM��h�,I� z�`Y$��  �0���hj>5K"G
�A��,@��O�t&�k�<2�X�/N���&�8���MQ�Dʹp��,���8�bJ�I��ңm�� c*V�`�L#�̍4[8 <���2r�r�I�υr?�Ӵ<퐐A�#]>����5��.��K���a4L�Op6��]��s���hO�0�d�c���;@N�4^�X��TJԸG�&1��cܹHti�E�O�<`1�Q�\c�DB�C:,@m(!b�O��O؁��AI�xS�Ɂ�9��
2�Ƀ����t&m�"��#/�l<�#{p]C�BD�M�	(V��dz�����D���L��"�<�H�/Ϯ�3}�ϐp���3�)����3�5�Cס���8wC� e໴kM�dp��'�(����O��4��O
��VS��ٵI܇w����d���#�c��Oo6̓����b�'�<9��)�I6b�A5��:�.x�Că��y�#P���C��0<���J)�^�A!0>�,��.��Yi��@5�E8d�H ���/dK"�	�fG�.���+"�B�>7�e�W%2Z���˾&z�xR�|���>z�PUm֊"aa�T�$}�Fx����|0�{$�ˎQ��-��� "�yB��C��a`�$f
 ��ښ{��Uȉ{b�|2bEsfe�t*�`� /*.m�N����RR��{;x(����1��9���ee^�����r���J	�m�~�;ե�:���kP�$}r�[�5�.�kӠ�)�\(��e���'WI��nrS�@f	��V4���Zi8a}RCm���E�B]r�I��]�+-T�p�/@1�Zu(�-ǽ$:�tF{��Z+U���	T�w���\)2, ��&.��S�i9�A/��(O��Sd�07�r�+"��2��2W��O���ئ!�H�SL+�<8a����$�/M�,�ũ� 6��l1�ݔ\��I=�(O����I�8����fZ�1!~(j��K="���%پ�Iw/AE��A��4�eY��Ks'Q:1��g���/N���<L���6���	�����gʐW�����MԠ%�:��?�薏,�̺��Iތ1G���<�v �L��Е#�����79�dʋ&c��'����J�F>�݉�ʤ!�Hej�	L0M|��)`K˿X��T�0�
���Z�/��S$&\�5��,�e�C;5^���va\��To�=�tj�λ?��:�uW�[�rb��'\n���Ju��T3pCm��'�n�6j"5���	�u�:�`��$#�A"V�	Oy�����������S�S�-#����2<g��r #Ѻ&����d�.|K�k��1��M\�Lɷ�]!.�TP�0p�z�@m޶8���'`�"}�'�:$�!.Z�3:��2��,-�xH�'\r!ʱ)�? Mk��%9�\e��4�6D�so�-�x��DV!�l����*p6DYP&О�a{Rަh����ʅ̟rtGL�!�s�f�̽˕�2D���Kәsڄp��K/��a=�I�w�DC#����>��alLJ�|� G	�C���Gl D�� ���rڙb���I��	��%R .k���%�|�`yr�ӆ=J-�CfP�	��,��i%D�a���?׬��u�K�'#L��c�u�����늵1:N����*qR�mD=#ĖAa%j��]����D�
T�4�a&Q�v*��"���=\JlI��6,OT!A��;88�ږ"���% E�� ]҈u�ѡ�+wde�ҍWH�'tH!��V�"/ݓ��Z�@��2 �~���1'�K�nQ�GAG�剤nI^��A�%q��@a�ώ}�̢<��(��,d��8I^ȝc��M}�oQ {��H�F��n� a
��HO��𦟈>�2����ɀ��Գ�+ɱL����&�iX����S�|W0���	#fc� �
�.90��sMS�����w���1�/V�p.���W 7���*�?<
��� �H�D�R�JI�<Ð�v���S�#?A!J���z��dߔs4�Ԛ�]ĦZ%FK3	�\]�5j+v)�(�V�2��5����5#ư`����)�.�ɷ�|��健i\=s֦V�K��ʓG.�s��I�-.�q��0mGyD�?v����I�c���ܸ�ybq��3�	�!N�̌IL���O�pIg΂�a,��b�J�<$
 �QV�����
r�)�@NIM�3���X��`�p�N�vQ�wK��4���&}1�����(20����4`�~]Q�gۂA�� w	C �a}G
3�l����<]R��	2����O��2cK\.o���-_�y�0�ӋN�
��Я�s�xh3ec�L�C�I�Nꤨ�fH�+*�j�s�	E�eW���^P�Pˌ��2,���W5��tEz�5*!A�2$� }��;�I�\�P���m���S���c���	�s�>�1��Ģh�4� �gȐ&��@3c�S<	J-���'���ċP(qZ�P�E�U�v)�q@?<�|�hwޙ����"O�d5b�F6o�D���E)�O��5�_7e�hh*��'{�L�x����;d�A+ܻ��O>ؙaJכT�#'a�Ĉ�i�(
�	��d�rxW ة�^ݑ����=y7(���$ry
Sȉ?m�I�n4Ҝ���ؐP���1u�J�iW��wF��xp͜�#�
L��%WZ���Ez�a����i�2C0!���0V
mٰ�X��4j	�a�X��HN�mFR��:B�RXvHTc:DѲ�Ʈ�l��'���AÆ�Z;>�"P-يPA�C��P��$��ܖJU��
�'�*����� 4�W�D� �X�/̠yQ&A[�`( �剞p�D�(�|�J��h�S�Z�����+��p���)7
#?� �@�-�]���-��ӡSK�A�ffք$9�|�a�G:��ށˤ@�bnƤd��}�e�W�<�g}���}{�|)@�պ�F����ݗ���[!2,��j3
�,|l�e��ӯw��\I5��!�@���Z�>V6��۵�� 5_>�t�gm#ON�[��_9G%^�``&^
^:,B�┞�򄑹8�ty� �j�3��"z긕�%�T!'�1��B�(����ȼt�pac$..�(�a��<Rj��FvƂ��6�"�O�Թ��/\�	k0._�U�(l�S�ɝWMx �&FH�1y:����"�1-¬���L���=BD"O�����2 (9�q�#.l�Z\�X��֩O��a�>E��m���&��$U�CDU��yB��L������r@��y�AT4��U�N �V�`h=�yR*��d�!�nA�q��q$��yҊ {M����E$�� ��y�OÁ8�FЉw�];�,8�'�3�y���`Z������8Sb	�yR�W����Q׍Z� �v%�\��y��w�\�"A�����(!���ybiG�q��I�Ɲ!Dw(ysNH��y�@�P�T�b�ߘB�������y��D�W���j�lN<2���qm��y��8"�n�ת��K�T�sfÌ �y����'2�� ��[(r��McFB8�y"��X�P����>^���ᥤ.�y�?(��Q!�0V f���J�yBN�} � ���S�����dj7�y2fѰW'TIP�_�D�d9tG�y�k�a�nUZ����9��]�C��3�y�J��"�\)
jK�.	��ز癑�y�읭rv��1�DE�W��1P���y�n�G(�g�Ô_����y
� ��1�@�\� ]:KI%f|q��"O�ՀgI)#�9�K�%{�\@A�"O\���%^����r��H�X�{'"O�q�UM�4T��:�v��|��"O\9󷏈�%+��s.�v�Vt��"O6P���=t�Q	5Kޚ\��-��"O���䙼i�EC+�Y�x���"O��;ä�D�8ա��׹)�@}[@"O�����,.%Ȕ��II�{| t�E"OXZ�o�u@̬�sCט=c��`"O�9�b��;gM�Ar&d�B�����"O�P�sK�'|����)b�X	��"O��aSEO-/��|2��^�Z��"O"��a�+�4��񏇤km�q�G"O�u"���9h�!s����Ilh��"O�4J�C/9sx�;!
#)HS�"O�@;�ڰT�qk��i���"O��Q ���M҂�F_�n��D"Oj� 2�Ӫ7)&��W �Pw$���y2햗K�"!J�KK�|9xVB�y���&<��9 e¾I� P���y�l��}zd�:�%�<;�
�q���.�y�NN����섃[Dtڢ��"�y��E�0�f�ƞ^Q�)I��2�yR`O7\�mi���k�%��f^�yr�Qxp@7��h��!9�ܒ�y�̂3|��ڇF	�^ 
���+��yr*��'Pi�J0P�8���#ݾ�y2�Ҏ�F��@-@P@D �Ê�yB
�+T&����4Ai�(��`��y�Mĥ]2�A�l�Q�<(Q靧�y�F҉s�,@jل@��-;Ga�>�y,�Xi¥�G�:
�1	�#P��yR�
�dY���B܎$$��C��&�y��ɚ^�=	A䞬",�YY�/:�yb˞���ٹB���D��i���y�Z!�Ti ���,���$�yB!%m;H qe�+��5�	��y�⏪s\��A��3 u�H@c�'�yr�ΒpԖ�0@�N��iۧA��yBC��N}����MրDh�Q��ڀ�y�Y{T���U�5.] ��L�yRÄl����/�"��'�_=�y¡�=S.6AѳfC
^��0EN��yR��q�t�
W`S�Q.��pFț�ybe��{q̅��K^�Pպe�*�ybEXT�����.V�"!s�A\��y[�{��(�&��Lۼ��(��y"m 0�@y�!иJ'���CKP6�y�.6��t(�&˱?&:t�3&�,�y�!�*T`�8g�2<��2��S��y�,Ԙ8�T9����A�썣����y"-_�sϜ��Te��80�����y�/�:�MQ@6T�a`��yr��Kra`��5-JMѷ�]$�y�G�S�ك�.
1.��4F��yB�Y�̸uwO�&��\@�E�7�'~ў����I��D2e92Y�$eʖv�4�"O>�� ��gJ2���RJ�~��0"Op��A�$r�ԃbCW/�T��@"O��*����q��I�a�+4��۷8O6��DU�!b�؀bNW�8-L�A�·B}ayR�ɨq�L|#!V����R�{��B�p�0���gޫQ��a��mӼS��C�)� ~��5L��[ft`�$M� ,}�hB�"O&�Q`,�7/<��\_L���"O��	�D��uݒI Eb
�"��y�"O��%�:O��7���G���"O̬�Ïɠ2��i����*r�@��*O�(��fMR�θBpN\�.b���
�'?����m��P*���@��*@bРI��E{���mM 4�`�J�X��V����y��]�8(�\p�b��a$N�(�y�JC�#��e�vo��D$�*p�O�ybFR��qt	�j ʧ����y2,���@�gc3r���6����y"�W�d��8�KQ�?r$��J���y�g�TKE��ΟD�ĩ���yrn��5�^�YA�><Fm���Ɖ�y�M"6Dz�Jc.	4q�$���y�M�6IHJ-�Ã[0XݸA���O��y"�F�����X0'�&(P!�[��y�Ύ/^�襋���G��eV��y�*�2e,��J�j��/�TH%�Q�y��]�w�T�R'P�*}eC��yBjY�c�p��G�
��m����8�yr茍E'��Ƀ��W�����yBj�=v�)��B?{b)�R�y�)�,zL$d) C�D'ʩ1�CW�y�AV�r�����	A�)r������yR-H�Z���D�6�8��u/��yE��e�x���@?����bն�yi�"#"(�iҖ8���cd���y��X V\j�
�@X�&�n`�t�V���k���Ow���$��[���dL\=2�u��'��̉!�"hj��jՊ5����}"�-LO*�FZ�Iz���E^Y���fO������+���Sf�\1��XcC	h�<q�R�2Gb����ح���Xb�<D{b�ˏ^�4�ZD:��sP-V�����p>y���Q�@����f������i�<ٱC�{��Mhы��;~
M2p�TL�<�jY�3�TY�ˎ�{�&Y��M[p�'�Q?�إ	��#��;��d�U�4ғw�a�4��-Yn !�H +�$	���[0�y��S?{�ؔ*��\�!H��"�,I����~�S��y��K�*��6	վʊiJ5���y�`��4z��pFO�xw�	u@�4�����> b�cNT��6.f�*C�UT8�� `� �~ҩK�c�����_/!��J�0�y,79l����HS_t=�F���O@�D�$�ӆ\ {)���ZݺQn
��y��Q�= :���NЫE�1�I���1�O�Y[��)O��9�a�
Af�(�"O�H#��F:M$�}��X'	�c��d>�S��1S�hd�C�l�4�S�Ӛ(rC䉸@jD��-\"Sh�=�$�+��B䉱p&�DbU�ڢ'���˧���B�	� rf�C��j�tYQ�(���B�I�p��EϜ�?FM`v㉪)0C�	2j�J�*Ĉb9<]z����$C�ɪ�Y"�)�x�*=J��ܨ�=YÓZ��yA "8�2��0 ��ȓI%ȼ�R�S�oX�#Y�(�����&.M��Z�X�   H�e�ȓ'j���, �m��C .
F�2ɇ�8���TVe�peR�ra�E�ȓ	��p��3(|Xq�揀 -��S�? Ta�%� u$�AV,�P0Tk"O�Q�eV�&)�2,�)�9pb"O�T��̎�9� %� {�V AR��[�OX��$��/ _v��&a�k X8{�'��8���JW@���F�:)�	�
�'Rx�kBj��S�ԙ�=-&< 
�'G|d�!A�sB� ��/��"ؒ �O�6m �O�U i߬.��{��A.J(RQ���'���;��0��M�R������>/r����eg�Lxׄ���2�Y"�(���x��I�i�*�jP�SP�$
�!��`ZPa�s�Δ!,"�(s
@�VTp<�ȓBϲ���]������̀&�(��GT��W�
�A�f��ʊnL��ȓ�`Y����,�S�J ����''ў"|����$��x�Ǭgp\�"IOd��lZU�'K�P�匟k�*�AE']?����'�|�!�Y�v��e��՝�@��	�'E�A	a��Xrk �P4:�'�~R0(P)���H0L����}�'BQh�)R�m��%j`�ՋjdT��'��Fˁ�r{�X� ���4.��e��y���(be/_(�(Gd���0=���Bd�p�����z��"�yB�4<ܾa	�
�D؛d�»�yr���L��B��B7�E�§�:�y+�d�օ�0�P!>uB��Ҏ��y�e��)���2U�=^?n�����y��9~鸧�I�QJB����G4�y"*80FyR3��[��a�S �(�y�b���$#�	ќN���2�H �?����*�j]��ጘe.hr�Fh�H ��1Vµpc���"G@�"m�����ȓs0�2疬I&hz��Iz�Hd���f�x�A�;`��!U.b*h�ȓ5>XdR*�$dJk/ן�����Pu��O�7ܼ:r+ڑjlن�G\a��O�<X���!�Y>���ȓ-�v�j��%�Qӡ%�3��Մȓy��E��O�r|��rNR��*)�ȓx�<4q�-M&xp�lAG����l��ʓH^�e@ABT�&�~�)w��3t��C�I[�\��f�0�`��Ȯ�yRKN�s�lK���|�d�[��/�y�G!v�2���Ŏ_c�je*ϑ�yr
�g��E)2��[;���t��yRd<sq����Ym�(+e[�y� !�hZ􋖀X:(2Dh���y��ݵ3���R'��H�RyP�B��y��۔d/�ŋӁҨ<X������1�y��u��0�*��@ļ1�AJ�yR�Ķ7��$V�O��x�0�G��y�&��<���e�ݱ8�EPp��y�a��"�k���"H��bI&�yr�1F�B\ɠ!4��hb�gN��y���a�h�A��Yc���u��y�T-v�ѓU��V���"tgڒ�y��K���X
�2R<(�1ӯ ��y��/ra��Zc�� Gn|HV�D7�y��U�S ����A�3�es��G,�y�/��C)���#��?3z!S�.B��yrmIt�L��9�ȩZ7�6�y��?� ᣷�4;��  � �y���Uwȝ�� �kt&�9�n"�y
� ��[�h��L���;�n͑? I(�"O�ٹ���h>\D*�>o�
�ّ"O�����.y� �i1��	��UY"O8 �@��d>�xB�Uw�	@"OB�����?5a���a
QsJbQ"O��Y��()�8�@� qk�AF"O�A���	�s@� A�$޼yr��J�"OE��J[f�nW9S\��"O,HC2JK��$�cƆ�L�d@e"O����b�}�$��
,$�t"O>y�M�7u8���&�PvH�#"O��V�ߖl�,"�ő=r6T��"O�T���E�p2}QeOT>2E���"O�@�a�H'n[\�N�{;|��U"OT�p���f�ڐ�҆�	.�)[�"O���*D�u*��V�0%B,�)�"O4A��X'O�	r�n�
\<���"O����C�3���A�����"Ov}�E�R(oH��V��`�~,�"O
)iT�"�����بB�� ��"O�"�(йo��X�,�#q�51s"O��xk�I��H`EQZ$ep�"O�5���yh��BK֑Un��s�"O~��
�b(hHѷ��3j��[�"O�U �*<w��6��$T�t�"O�yH�+[hՈG�M>U�)q�"OBi�DH[�o�i�2A PQ ��v"O0$X�EI�U��x����v��r"O&�z��Q�"���C��<�"O����kT�{7m�cު���"O�����>.9lU:%� 0M��x��"O�ɛ�V�q�B;B�\]kV"O��A��ӞK�x��J��E���C"OLͻqJD�:��$��QM��2"O���GY=M@�7I�9,�"O�]鶩�
SXĄ�R0m��< P"O�0b0mS	8��ّ���5]��"O��9S�ԝj��<��-��b2ޝ�&"OʸXdI!x�B;��VDƒ "O@�*2��yT舙r�\�����"O�ja�[3V�В�FD�}X-�"OjH�!j�=��9����(l�ј "O�2��gv:�R��6�M,y�!�D8<��`�*]U���@u+C~�!��P.Q� �0m!1C%I��K�!��,v����b_5\�0d��+!�n�sNN�3�U�!!
��y�"O�I8�����81�T�2�>ې"Oj-�Ė3>�0�٦��3޸Q�"OH�4��j�>4J d
,�4Yb�"O�ٱ��*>D����4}z;�"O���� 3�$���,L�/a�͸u"O�R&�	�nٞ��%Qt`<�J"O���n݅p��% *�Hs�H{�"O���"�T�E���H�
ƀ��"O"�p�ϱY�h��扐�6�zȓ"OBDPB%�;��8�)��"ՔZ�"O���QꚲUf������.f˶�RR"O�0�CK "X�"(�&'�q��"O���&�ӻb�:ax�ΉA�L��"OЁRĆ[o��
�֧� ��"Op��T�R��8ZfOˆT�Xx�4"O6]z'�B�x.]WE�5p�v�b�"O�|!���%!N���!���� "O� Ԥ�h;d�	 V��b���X""O���⃙�7�4˔#ĝM����"O��x���]��� A�> �.�Z4"O�lK�E�?]��$+a
�*м�(C"O8@[âʑE���0тQ�i���C"O����[@�q�P��x�Ԝ��"O�C�i�
���֞�ځk�"Otq�戆�8-D9��B�<ޭ�P"O��YUh��Ύ8�e!ݝ<���R"O�e��DMj(p���>*�H*"O��Q�@RBx���o�l�Ҽ#q"O����K-y�5�S���/��4��"O�pr&N�X�0xԯ70��|��"Or� -�D i�������"O�ر�ѷ^�����8C��p�"O�G���]b9`�OU>0P��"Ot��ƃ߫R�Z r$�ƭkݶ��f"O�pY�� sځZ�)]�!n�=c4"ON-+��8Xd�lA�H؏z�h�"O���f+Ģ���)�y�ػd"O*];`��]�"�X�I@�i��=c�"O�1f�]�6��K�b�]�U"O�Z�5'묨�Ce�S��xQ�"O4���U?�Je�A�D�?b\��"Ovd�e ��tr��4`�3 5�8S�"O�a�g�TS�l��.K "r�	V"OfA����I�h(�+I)'����"Oj�Z$�Ү`�ɲ�
�M
``a4"O&�3GD�4i��)%��e�.ᚣ"Oz�#5_�>�͓���	��t��"O�,��*ܰG�$�4
�(�.!��"O �W"���P�	�	�@89j"Oh]`!�}����R�[/e+���"ObX���J�bb��DcO�sH��"O&$�������(^ ��2b"O>5CR)�Zn���UO�? ��hc"O\��@�R�0�MRPNTV��L�"OxݸVf��R���s�N�0q���ZC"O68Bh�>c����$�A	�@1��"OAu�}KY
��KÇAb�: "O�8���Gf�����Ǔ$�p��%"O"��w�,�~A�Q�͂\�T"OrM��	8w�}I�f���`t"Ot���u��i�%�tɖ��"O����
�0����CD�w$h�"Ot3���Ip���9e~�I"O�L�F۰~Uڍc�5-a����"O�m����Rf���&��?KgT�҇"O|��!�0CD��RB��+8@���""O��i�q�h}{C�%L0�0�"O^ñJ��c{( At L�P�]"�"OLqj�'�6,�n�Ccj0|����"O\��w�T-�2��f�?o��#"O����뎘L�^|���I��2&"O��Pg&E��)�c�-є4 "O�p9Ph؍W���-+���2"O^���)�2/S~���&�""O@58���[�$a0�ӱ\�uY�"O
e:��f�����'h͐t�T"O�Y�P�U\�}�B��N����1"O��AqEځer�ScJK�lƔMSp"O6�b&�`*���Ӧ?X�@A3"Ox���؏ �()T*�%W^���"O$U:�� k��	0�@2��՛�"O� �БŠ�?u�*����!k>���"Ov��'%E8$�A�&M�n���"O�a*�mZ#?9�lS-Ƹ[ʒ\S"Od� �H�E�룉��_�5c "O�]; ��F��@VIP����"O8)�A��4�ܒ����	��1�"O��C��"2J��(Q63��Ḕ"O���-�.{tB�X����,���"O��Ѓ�lh(����8I�\�"O�yaN�8|�����S�x˸hT"O�S����lܘ�8udЗ3+��D"O�DG�)!B��2a�0Z"�4�f"O(���	ދZ�l0aV����)�"O��Y�60�"��&9�\Ԉ�"O��a�cрm֪|��f(��@AF"OT18�.�*v�H#�((^4	+�"OF����m��|!P�@�K�`x��"O�3����2�,�h��L���R�"Oji�n��� <�N�;s|h�"O�u����l J �۬r\��C"O�ݢ�A��qsa�z�"�B"O8�C�lpN�A-� N�@��"O�s�/��8BԳEa��dk^�j�"Ob *@8VP �rc:�� "O"$�wc0����J%�f��"OX�r˖ j�xY �L aRb"O~	�C!S�����nZ)[�x��"Oƙ2�	@�KE�v�Ҁ30(�y��c��/eF�Q˴�P��y��ֵ[3^�@�+�\%��AW����y"�ƶ{�m���ļY:prv�Ò�y� T��$��J�'���aN��y�O�6�.�2�H�"d�DI���y��ܗ\%xeC��N�Q*��9T��
�y"-̨QM�u[�x�Z�`sO;�yr퓢*(��3�ں#F|�A�+��y�'%+�0ɪ⧅� ��	Ǌ�yr(G64 �I���B%�5
"���y���n����
D�J�@��р�y"���*��V'���g�#�yR���kH:A�IH�K�����M!�y ]1(@�͠Ӣ�3�|L�6E�#�y�B��%>/X�h#�\�y�/�Y50e��δ$@:|�N��y"�T�V���sڼPLhF���y�R�y!&�%\؝p�K��y�ُ:�f,��-�Q9@�7�y��N�]��%�k\�v�U0a�.�y��V�N �	�u����0J.�yrcD�g�*�zX+D� �2��ȓ0�ݒP"ޙ/̾���cL_"��ȓq��1�GU3x�Vႄ����$I��4l�	�hPzH�T�$W"r��I�(e��-��\��^�J��ȓ06�a�ȅUJ�sၐ"~��ȓ8X�	J1���t�T ��� %��OE����dpiB�N2t��ȓ +�lY�J�Y69��kH��x�ȓxf.��� �U��ixu�_�	�V��ȓW���R+A�4�b`(@��0���ȓ���
�~�8M �L�v�&��ȓ�@ܱ0�.(
L���ȜU��q�ȓ�$�ZI_�	���A�v�V�ȓ,�B�æ׳h��ĨdWtR0��S�? �H&/�<56�ذ��5���a"O�,҅G��y���V�e`c"O��R���	���	�mƨ9��Tz�"O%������D�b� x�1"O̼���ղc�t��m�6 �$}H�"Oތ*�#ߔp���4*��*��]9�"Ov� F�1=�@,P�N���c�"O^z��
q,�������d�r"O�����1��]S�R�*��xs1"O:��R��J���P�	Jl+0"O:iɔd̐��`��K�v�rQz"O����@�"y�U�v�@~��h��"O`�H�Q�{W�5��Bå=�fU��"O�*�FA7��(��KӮl�"O~��r*�7_.�PrBA�_��	d"O�`�D��=*��y�@��b���U"O�\@��<���h��15"OL�4(��\�B �t��I�hr"O��+�'	W��I��M�#��(�Q"O���Β�m����R�^u��8��"O(q�pf�G�R�	&L���t��"O��y���41�T�%^�*�|tQ"O*#!F4h �҂��9��0�'"OB�STg@����`�͎�"O�mk삎
q�5B�kC)��H"!"O��C�Hm,��q3j�BӨy��"O������9��L� ��@!t"OXY���77���h�i8��E��"O�=[p���z���rƉŗ7���("O��Z�.�e.�Pe�%V�ɘ7"O�1�!�շ>����I���%�"Ob�8���n!`���-��y��zE"O01���4
ۦ���솖���"O8�sN̺Mn$1�PAJ�X|��34"Ohs m�#�8j��;],��A"O`p��C'�h�Wl� W�d��"OJ����n ��U�մ9�b�� "O���Ќ<6hv��,]��s"O�U���+q+� ��ߎQ3Ƶ)"O*�p!
��ue �����B$�$�5"O���U3.d�����o�<�"OFicB�]�`��f��E^�H�"O]���&��q�@[�v���%"O���G��b��D��MϐoY T!�"O�	��O���6�3qBz(��"OR`�ϑ�\�`1p���=�`�C2"OR��RKѐ@��'M�VY,��"O"X2����X-+��E���E#`"O"T�����v�hU�X�����w"O�$ cJ��vQ�T���S:>� Dp"O�ظ��H?L�X��N����Xf"O �P��#�(E��㘁#1��7"O��T��:8�#��,�T�a��(D����ML�	�x�&̃7P�r"k:D������$�T�r	�7�}3ƈ6D����.m7<�#��}���Յ"D���eƆ"+|u�	W\��z6?D� C�KX8��9��/T(�F�
�*>D�\���Եp�TDzb���)��<D�8i���6Q�$ap��uj 8�e�:D��*��rp^�Q���(���7D��8 �2iX8 �&�e\�1�):D�$�s�U�) ҍ�j�)���i<D��	��[�v���Y�����:D�� VRBJ<NqIe��/[�x9��"O�� �U��[�n�0>�`F%D�dr�'�]�P���g�)S��Ć"D����J�X�p���>dv�kB�?D� "@ʔ:���AX,���a=D�l�$���9R�,B>����!D�@��F�JqY+u�,R!��QD� D�P
��A�~>20�R.�5�����?D��TmŪ)N�Q����g�|@���=D��!W�(}r`�K
:Ոh���0D��c�����FA��n	����k2D���妇�r(����E,�����/D��)樚��F|1*4kӀi2�e-D���6��@>j���։q�>�a'�?D�l��ѩV&fЋ��R�/��|H��<D�����J�ek�q��Ț4ČY�>D������f[6<�3�ֈ�g�'D���2�ʵ�S 5Q����;D���EI=i��(���<�ڜ���:D�\xV�(;H� ���7[�L9t�"D�(����,H֑��E�n��%.D�,�ԭ���U��Q+aZ���,D��J �^_���bN��vyrsA=D�̋�$�?��`�� �|\����;D��8�/W�&9�m�+�K1�@�&:D�8���,����F�,d�lP��8D��Y�Ȏ06��9�!�/q�R�7D��1ĥՑ��ģ���/yn�$ D�P��M@�Q��j1 VT�`�>D�������J��h��H'�n9�@7D��� G� &��:G%��e2T:�6D�DIq+؁ ��[Ƈ'L�8���  D��� f֤�aP��D�;}2]�D;D�(��J�����P��ji5i5;D��"�Ñ1��\��_� 
J����&D���4aM-�*̣���Av����8D��R󤙍^A��3fL_�a�Z����*D�HJ1A�,tKj�#��o�P�b� 'D���S�d�2p���p�rCO$D�L��U?E{�@3POT"=��`&E"D��8���k�!T'e� ��#D��`�H�? �8�8�͑%|k��Z��.D���T.Q�{�q�0��?�}Z��!D�$x� Β@������Wt�M���;D�гR��c5F��ʊ|��$;D�����1l�4 rn	2vA['#;D��8�*��G��t�`
�[aq"��8D��"���e"~�`b"D$~F
M�C�4D��I�gF�H��x��EP�� ��i1D�h��/O�rK2��K�*�p8)�.D�$�E��.)����F|�p�ȶ�2D���V��i��.�n��0D���i��@��LI���P�+g�)D��JF��?� �
�P-C��&D�x:q��h�Nt���R�.�Z��9D���`��
jĉ���2.f�g�%D��S�#dا�T�&���CP�%D� � �U.i��"�g��=v����F0D���öi��X3���+K�x�D9D��i�#Z�N�θȷMَ"���O2D��;p�� }~�"b��� ���Ņ1D���3�^3��)VoR3����R�/D�@����	hڀ�a��}X�<�uG*D�`!�Բt�����m�2T0n܀�H&D�� ���8?.	bd��9=U"OR4��k ap�Ɽ��`����7"O���G��UE���$Z9i��Y�"O���F��f�)���t����"O20��ęG4���b)�?�y��#)`h�Ң��B��b�j���yb$Z%2��b��@��>�t���y�?l9��$�	@ԥ���Υ�y�@"Hv�)J�j���a5bՔ�yb!۾N��q����S6t1�I
�yH!B�ԡQ�M������I��yr�0�����@[L%#j
�'����L֥+���Aa�Y�t�p��	�'	
P��#ʪ5'*E��,��9�0���':||9��@�¼�G�]]�|�#�'���P$�q%v=;�D��O�X��'J���F��5:�I�s��p1�i��'y�s�J����E�PVQ�'^^�H'�3T����G��^G��0�'8�!��<&'��� \��k�'r0�+�g\�S@���F�C �8�S�'lJ����CQ��C@T�\��'z�Xy��F^SL��է\=s��uk�'b�� �=B��0���
o�J$Q�'��"��I&6\�+0���d��a�'�*�`2̞[-���v�ϗ����'F�*c+׻��$�&&�oy��(�'�d{����:�3<~�ؑCD��y2�ַr��]�D�	4t�Z��ئ�y�I�Q��@�䜘}V�l83i��yB"!3~��ӕ�߹_���:�D^�yR�1e��� KY$VY:Ug�W��y�I_1'%)K �K e�������y	�\�eiSa�6�����(�yb��a��(�!G��@���ǩ�y2��:�zMj��S{Q��R򪍜�y2�ׇ5���祈�x���2�X �y�a\�5����hG�s������ńȓtЬ=#Dܳ!��)��a��wjȨ���A;$�ϭo�8���ʡQe�� #�$�#K��2"�@�L{�q"O����.� U
��!���8�}��"O�ظӣkw
�iȧ�r���"O��Q�ϊ�C�	q5E�9t.N���"O�բm 
=�zhp������:�"O���N��5U��zP�H�4�j���"O�M�u�+�vKa�\-�|���"O4jG&ƊbX����K�}�I��"O�ܹ��;2O^�� g�5/�8@�"O:y7��	I��):��#pd`�"O|8���FM��a��-�q�g"O,�@��ܒ��|�6A��@�(�"O6$���$3!th�a���0	ܔb"O��3"M+4[�9i�g 3 �Ւ�"O�3���W�$�a�f�P�d9�c"O��d�=E^����%O�c��$�"O����H�7!!)���A��X�2�"O����E��7�K8X��"OF�Q�C���:�B#"O�IW/�%� 	���3`̬AP"OZ`+�Zk"��&l߅T�`�"Ofh��@ZP�*@ޑoS��J0"O�C�a�&��s���-Pĩr"O>��֨�7m��k��NCX�B"O� l��C�nk�,�)k����"O� k�i�OO�ȲQ�(�x5��'YFx
���	@��+T�^�_�D�p�'�dC4 �E�j\�B��n�P���'��k�OԴU��w,�cv�#�'E��פ�OSh��ɀ�[	�'j���C�D&J�n�+�޵��'z^�S1��-&(}��ȁFLt��'Ѣ��� V�&�z4cĽ�ʡ��^�<$DE�R!r�0g�L,$���k�@�<)�l� q������#W�Ux�<�b��"�$(0��0N>i�bXp�<�Ų�� �G�)L%8��ƚx߀C�ɅD��%��Nљk�8ᡐJE�je�B�3�����#^U�4ҧ&^�B��B��5 �j4#����� �p��B�I-;��Y�WA�e��ha��يe��B��-a� �4�ۨik�:/���1�*D�T��ʁ.;���J��,g
N��E=D�Dh�On	�ِ&G��v��A"':D����#r�v����M8��I�p�6D��H��V�h<�g��72�(UH7D�@��m�䠕m{������;E*B�=X�Aq�R�D�"��Q��P�HB䉌1����D�$��̺��NM�,B�	+�R��E#�9XAٖ,P0*nB�I�!���@����L6u��C�	"w����r#�'Zdȕ�eE���C䉿5րm�4D�!.V��7-R��C�I�-GTu)���y�q��]U	�B�ɔO��cR�(|�8�V[�x�RB�ɣ*"���W�Z�-��]3N�|B�I�+9.t��jT�Q��u@���&}�xB�I*&�hS�GV�I@�j�4�"C�IJ��͐���g܄���
�-`C䉄l���´oɀK����2`C�	'd����gݔlz0��[%-��B�	�qȶ��p�yp� X��W���B�	7Cs�Pڂƈ��(9���+8C�Ir0:d0�ʜ�+��D�����W��B䉊A��Ā�"=���a]�Mh"C�I�ror{0R�"� ���%�B�I�T��:�
��5��ei�G&B��B��k�������5x���%�3ԲB䉒y���I1"�� � ���E�--��C�ɛ#�!��-͵^y��y'$_;�C��:J<��A�G�=y��PBN�g�:C�I��< � �8t��]�錐H� C�I�b$���Ãͻ�z-�עM{;�B�	%u�� :�i j%4!2��k}�B�	?J.����j��P��9w��B�ɔ!.* ��
1= �E��*�t(�B�Ʉ_�Z P�f�&b޸	�W�u>B䉢t���av!�>[��9�R��6T4B��4o��S�	�^?��U�A�B��2rF`��m�(�d	��R#Jw&B�	�?
u�u�gŚ�ud���*O왪ei�L����"׃w�z<	�"O�!�%�c�T�Fa�40��4�"Oj�і)	̔,7!�6&��jw"O��t�`9ʀ��	�9��4"O��2��((x�
e�^�'$��*!"O��̈e}!�d㉷+B�Z�"O^詁	J!hx�!F�Tz�C�"O� (%�d��Hy�/�!p�[�"O�m� ��a����� aR"O���V=����F<�2�XG"O�@��ݘ>]��cW�E}L��"O�ub�F"D��X�gf�2Pn�X�"OZ�yWl	(g'�)h�RC{
��1"Of|{�@P9Y���s5	��P�"O�E�&-��&=4����ht:�"OXMj��Y�|������E�b(��"O� ��/� <��0UǮM���c"O��A2� �C�-bϙά(:R"O��aJ'R����0�u�X��W"O ]x"��pۢA��I�A]\�!�"O�T	uAP)r�rt���"���B"O���3j�2�ȭ�3#E�L01��"O>\i�df�x��Z�`j�10"O�ѱ6��<�|*�d2���J�"OT�3�MW|0r��đnȰ�{�"O6)��!Z��;�`R ��踶"O42F��
-J�3�@DMXla�"O�� ���W$B�B�~}�"OHD*K�+!������1x���Ѷ"O0� ��!�y��Ҽ�|-��"O�XᗃH�b0�m` EY~�(�"OdQ�`�DV��2%$$*�n0ٱ"O�M���D=`��%��m�{h����"O��̲҄"�+N�3�r|yb%GX�<1҅�a��"��-;I^��f��z@�X./N�82 �Y�z�8Єȓs��}� ◽�n�z�@�ae�|��1��	�˒7H-`���A	3h+����M_L�+�Q�:�Zp&�R_�х�P�0�$�߼+p��y�g�^����&�§�Q`ׂ5��ύ-�r���(�����lI�t�(SP��(z��ȓNg��+d'W49�h5�V�ۢO+t�ȓ(0iQ�*TIB�*���2?Ɣ�ȓyU6U�r	7�H��#i�d@A��wPl�H�,V�4�a/ج[9���dT�g�ʘXst�ō�U`|8��U�0	��A\�*B�c�	#��̆�rj��S�h\1����:S�p��ȓ*).m���ӆL��zb�ĝT;J���3���FAth��cb��1U.>a�ȓ�ii���.\��Bn�^�\��9u��g
�/?��5b��5�PȆȓ6A�D��O�1B��L*
h���D������	Ua\
�Cќ�lu��5�&��!ک�qӍ�1(`��l#l�:3�³p-~ ��+�m�ȓl�R�`g��JKH��t�Ĕ#�]�ȓ�B��Ce��)(�Y�"S�k쩇�/�1-؂*�8 ���/[�m��N�2��:��HR#�Q�F���4�J�S���/;���&F sf̆�]n�ő5b�����c�dr���ȓETEj�#L	�P�0*�(T����)+�5y��6~�Va��\�`�*���� m�U��$+�����ߥ&��Ԅȓ*��@8w�ژW��$���L�`�ȓ;N2@cb �	P�<��/�$H�ȓ'��0(�L�,����B�r��܆ȓ��)�P���Hm��I��Q�@P���ȓ�jAȇ�5L��qgG�o�\8��S�? �-�t):Q��Cu��qE:�{�"O�*�<���P�!&#�@sD"O��KΘv9fqx�焍:���"O���w���`��}i��Ux:a��"O�j6�ҙ��1X�&[�B[��9�"O!"�
� m��G��!KT�P�"O\!�ѧV�A��m@F�KD�ݳW"O��wHUQ�)���F(G�>BD"O��X1�-.zd�ء�8+����"O�M��jW�"���ޏ
?H@E"O��"�b_	ve A��H��Ԛ���"O~�:�m�*f�1D����5`&"O��(w��o��I� 
e�"���"O�kC┃)m����ЛSz�0aA"Ov�B��H�]g���1I�-����T"O8�R�OΚ�zЍ߿d�n�+T"O�\KrJD�63\ ��ȳ����"O�hp���$�eK��ǀ1Ԁ驅"O�|�	И
l|�HE�Ik�8���"OB�S$��?'����(��A�"O�}{Vj���6�0��"{����7"O^�h���T,�P���ҝr�t�8�"O1���A�59v�������x�6"O|�Pa�����z�J�>�8�h�"O�5[0�
E�Bw��%O�,���"O�0���!T����ѨH�(��pK2"O��8�o@ p;����%Q�Ҝ�
�'�
��󯑠h6�E $B�}f�:�'#R�a�D��{wU8��mR��P�'�j��TA��f��{A�ֵ0��Y �'�x�1��l��b���$0=��[�'I4i�#^0BV�@iD�,�:�A�'���8eJ$
R�4D�x�<q��'v�AP��X�Y�$��s��g�xq@	�'�Xͳc�\0�v	�HަPY�'^V(��a��u�2�+�ϕ$/}����'��X��Rw8�A����ٻ�'�)T�X�y�����!:��:�'����]kN�z�D��J�ј�'�"�ᓨĂLxe����`��'�2y`V�9w˚��%�(J	�'�x���+"wTL����$nO�)�'m���B�߷YK��bbC����{�'$r��p�]6S��I��J��Ď`��'z������-9��Pxr���,u�' �X1DM7Q�� ��)ՙ�n��'���(v��}W�����L�����'��4�����=>1Y!�$0��݃	�'4@�:CDOK}�Cd��S":���'H����V��Y���-LG�(
�'�<�H�'��;ˌ��cb
.�8�	�'��Y�_+^	�TK�@HB��4	�'�dU�FaP�n����3�Q>���p�'hZ�@��dA��s�#e���'�p G�!v�X�#P3]�nhb�'=��[��Ԁy����Ĵ><�'ҩx�ɜ��0a{��G�� 	�'f��h�N�8#���`E��'FUj�'F�I���<l���z��(-�5��'��IZw�!wV�ě�,
&���'�F�&�N�T_����t{�̱
�'�`Q�Î�.r$4q�`OƘp>��
�'���U��v�`���
2�2E*�'�n�ib�I���Y2��e����� ���,�%r��7v�u�%"O(��hV�M��݋��O!�(���*O�x@��#��(�i�]YD���'���!��,j��"0J�S� }��'�`��Rh���H₥\D��)�
�'��(�ãV%I�&�R��A�(�q
�'�"x[r�L{�0�Rr(߮e�x�X
�'0�A"�[
ڈ�ڠ��VV੄�z�n	��Ɵ$SV��� �s����n��8��F�3`�{ ܪ%`��v�>�iׂ��uG���`��2���ȓ{�}Z��G�a��X�B-ϲd����ȓ\�����d�)j�T �!ՇU�l��ȓ4����J�7㰑c��ٺk����g�z�SGK����+sDG�l��ȓE�J�e�	4@���q�D��+K�̅ȓx`��(sNAaW0��Fʝ�xv�<��Ϧ`aP%T!G�P��ǣ�d����<���@�<wF�!��
	<����ȓ����M5���؎� �昆ȓfN�����.wE !��W�Q�Ƅ��W:Q ���,��Mz#�	5x���(R��S'/��Q�dP�@H��Ɇȓz����'_զtx+��C|n���@��qIX�ze��X�"�1����>B|H��n�� �|�fR&;H�ȓ=I(l���6i<��!@�),��@����k�3���E#XSk\��ȓrz}��� ��,���ENQ���l"��Ə��wz��t�X�&����ȓ8�M"�X%F�ҭe�	"\܆ȓ5�D���� t�B��qmI�\��D�ȓ_Ɗ@+�[�<���؛w}���ȓW&�B��P#N`*��6�� �J���YW@t �@L,}`NH�N��-MTM��?z>QZ���(׸P�t����H�ȓȸ���(���ٔ�;N�l��d� a�'X%,�	b��e�̇ȓj��0���)�煟9�z$��Pª��`�?#*�af4ZP��<�eQ��&���xt��t�����Joܼi�)Og��� Hũ_~z���F��(�$�M�Бw���5)��Q�r�h�F�<6�^�Ԭ�(S� �ȓrs�h��E�(e�è̏Es�y��|���9vb��`.�qB�x��T�ȓ-x�h�=�-�1��[fx!�ȓf�vx8�]<�L"�k��+ ,��ȓp��0H��L�P���A��k&4]�ȓJY쓔��,e�D+��w����5�r����o���䤐�:��u��gVܡ�߀fw��HC��i�ȓ	z�4:�lC�'�"0v�A�c����{���q��w_*�C #�N����/lԴCFj\3�09����%�r�ȓ}��2�#H�`|2���o�^ʼ�ȓZ�@�mi�h#Wk�-�r�ȓ46�2��	3�H����9��P�ȓ~�(�C�!�;k%<-��������_��x�V F�	z�ЩP/��K�؅�0��e�d&J�l�^�)�DF$�%�ȓJ�p� �]ys��H�w����ȓl[ֽ���)c� q�"������3T(��̍�;�B��݃;�����S�? ����Ŗ3R6ya�b�Ԕ�"O��S��g�n%�����	ZQ"On����VbSnE"%�I*$��ق`"O|��`�1}��XQ'�D�{�(�Y5"Oֱ�2�O�0x`�ŴD�*�:�"OV��g _ d5����b[8A�bD{�"O��ÁbFFt6����q�J��"O�!��e��:%�^�M~
��d"Ov���C- �����c�-$"OJ��&o^=I���O�B���"OD=a �V�Vl�LA��WmNI�`"O�%�W	��┫տ�"�"Od�!�(Štkv�%�/�My�"O��͗�o
y��#�"JW��zG"O܅!W/�F�4�d��%<Nh��"OP�8� �C�,����;���"O2! 9�XU�a� $m����v"O�����2@�4�ҡm�~ xB"O6m:N��}"�)�w�_2FqZ!�s"O��!Sl��DY��
�F��B"Of�	�@�_�|����:`V�a�"O�=�6�a�*�B3�I�.�6$�1"O�H*���*ɰl[a��>�e5"O�ܚ���2.�(
".�3k`dy"O
�����.�0lS��b��2"O����*Պk�)W�H�Φ�@"O��	QJ�e���&+�B�^A��"OZ]B��\xElb�	�.0��h�'"O�iƣS/4�����h/^|Z�"O��xE�p�Z�*��ۦ(Q�YX�"OZ���N��t��mU'nFTx��"OpA����Fl��D.N����W"O����o۬)��!3g��4���"O�E0&ٰw��t����6�8q��"O��:�MF�	u��ؔ���:L���&"O�P{�T�q�@Z#��]��"O�컃Wt/44+7BP3Ƙ��"O�`s ��b�����XE��'~��vm�2'7�\R`��^{�]j
�'����/�y��Ȗᕩ]��hH�'�|ƫ�a3lxQ&�UI�
�' y���g��9���'S�D�j	�'YHq��k6kp�`�斈|���0�'��!ؓJ���b%/Aμ�C�'�`�R�^�Z@�l�$n��;IҌ�'/x��@�Ҡ@�Zy*ӊJ�4�¥!�'���Zw#%l۴�b�M�2+l8{�'�"(��%X&}Ef�sg��5�@!�'��L��$]�g،	+r��v+b���'U`��V,��_;���Ƌ�j��mR�'¼�)S�ۘL9f�s�D�e��
�'�z�Ba��#]��A�i=4��<��'�� �W�C:I(`@!̒-�H�Z�'��U��"����9q�݇(��(�
�'@u��J"+��y�65�8@�'���rg�ľT�6�x����#�l��'c��z��$@���p�H+fx��'�)tF�R� �1Ь� ^��ʓp4�@b�C�,��d�q�� ���ȓ06�M1�ܼXjQ�Ű�4�ȓ	s�c��nt�fө;p<�ȓ_d$�j���.P�i��νc�PT��L�@�y0���Rz\<:�P��ê#D���IΞk!���P/\��0r�?D�� \8&	�\DI�W�@t̀ڀ"O�!��̖�"a$�Bl�R<�1	�"O�g��0�R1�v �6'z%i�"O@��+�-��,����i�!�"O��(W矟*�85�U� *^:��k�"O.��Ã?W�1؀K��W�F��%"O�yɄ�Q�:J�IU,��.��"O8�)e� l%8y6��q��ܪ"O^dWhҋ4ܚEk��M�8�N��"O 0S�^�*NbQ2%�1yp�&"O\����� e��`���ZrV�(1"O�wo� ~[�yOFG�R���"O�}��K8���!�#��9��"O؃�#�_	����BN0�l�i�"O�}k�% �0��qڴ�O A�Z��"Ol�C6�9qz0�`���7+@�5Pf"O<�#��١I)�lje$rN~��#"O�)��� r�d��X8��"O��÷ з<�T�gJ�X4�ɳ�"O%�pJ^3�1"��վtA|���"Op��E�nX]9g�	�1aftY�"O�x@?=�T�i"�ɵ]N�,��"O��j�(ߠ�d��SkT?8�!��"O�<#a��iU�i�@�_� ��)"O���$O�=f,T�S@�DD��"Oj}3�?SR�٧�DZ0r9)C"O�`ӓN6��F,�"��"O\!#�-�2O��%�b*�9 8`xY�"Oځ��Mغ*�&T`��ѤV.��:�"Op$K�E�%(��,��X�N��}�D"O�4��曲
8��΁�-D��"O����I#�֥���N<;;�Y��"Op��AE��N���#5�ϊ8�tU�A"O�͸0/�'P���yP�M�{��١�"O.�Coޤ1��	�be�Z��"O�(G߀U
Q1���l��)�"OԬ"4�Մ->�R�H�)�:� �"O��*���'C��0x�(�s�ș�"OtݠG&�Y�4P`���-G�x��"O���)\���b4eק2,0r�"O��9ЄI�g�>��=$�"OP�!kЙww|�����K#r��E"OP�k�)�ƐI�1��p
	i�"O�}��%D�l�v�x ���,
�bd"OL�))�Q}q�p]d뤽�'"O�%�4FM%.|i%.�
\vh1�"O4鋶)�r
&H� � �!�L`�"OL��3f����O�p4�|#�"O�X5O܄dZ8�Cݮ(>j�!�"O��6��<��$c�:$^�k�"Oz�R��%�Flr&H�[�X�#"Ot
�iޢ[|x5�7�Ny�4��"O�I�vLQ;v[jIs�ژB����r"Or�,Ul��%�ϋ$� ���y��SK��D2#�TLj0ё��+�yb/ڐc�r��5�ʲ&Ѯ�A�[��y"� �$�� �%���E�Ո�yB,���zy"5�7����Ë�y�èxP%�G��(��1��o��yR	��_��Kcgۇ$`l���
�y���u�J�
�!#/�4��4����yrC�SmpHӕL��"ܒ�33�,�ybFXr��0N�61��p�U��y��H�6VL�����6�B�3�����y
� "��fkʰf���[1�»4����d"OJk1�Զg�X��U�K�<	�E"O�=�fdJ06�|r�E%9�Bh#F"Ov0���K8&Ŧ��eV)4l�v"O�����PA�$@·�	f��}�"O��ڄ�W.@F�� b�#]�	
F"O���1���bѓc�tBla: "O�I!1�@�vެ$`s�N#9?H`*�"OT�* *Pn��I񀒊G��9p"O`4�d�,!�m#��I�e(3"O*l�1��z��=���8	��D(q"Ot1I�AP�B��ѫD@��$Z�"O�Y�AU9'�4Y���[����"O�9�Ѐ9=b>x�"�aT3�"Oؽ� 4\�łA��$}�"OЀ�U
P��H��.��p�4���"O��k����N.�L��͓�qy<� ""O
Y�,� 6�1b�ADk�L�"O(U�E�������g�f����"O�����H�]=.%z��P-gPP��d"O�(Q��G�r�m� ��4�(Փ�"O����ρ/\rE�iG��]�0"O�e �!3�&��	o��is�"O��Y��.Ka �@2�C..�z|��"O�}�`��G� �(A�{}�"O����6۾H��M�^��ݩ�"O�������G�X,M�a��#D���ԎV�j���H5�Q1�B���*?D��q5��lS ��a��Q$)�V�:D�TZdR�@�y���+258�H:D��bD�*��  � Ԑ2�]"Sm7D�p�P�a�����lP�E(�c��'D� H'����UO2;�޼�a&2D�D���\E j�*#E��2��l��/D���Ɗ�'3��DH]�"О��/D�p*7�M>V`�9���=��yU)D���Ήe�Z`���otԲqA)D��'eK�̑���8q4�
(D�j4.O�o2��4�]Q�Ph3�j$D� ���ȋU�Z�PFc!l�fp��"D�x��:6hP��dCG?N�y�Ɓ"D���B.Xnd(�@Z���#D� :s� l�Q��6n-�])ק/D� �6���-�J����_��i�j,D��1�K	�
8�=+$ޯ}7.��)D�\i�F]W(�*��T:� ��&+D�(Q�8�b� �O��̊d?D���Uo�	�>m���J�prAN(D��FB�moҰI�&�eh�9f�%D�)$n���j@"G�9u�Mٶ�"D�����K����,��H	��bp� D���fBM$;�ʼ�ec���8� D��Öו4����#�NDv�	�#D��ك�Ù$��!f�ح�F!Swg#D���F/$<���b&T�$˱L"D��pA�
*���C�>��2+ D�T@Giܪ<-��P�MR�hqz�?D�IK� <ظ
�U�~��)>D�t�q�����B!	K�jdV��S�8D��i�&�1[kJ��'�۟y�`��aD2D��8s���(�vQ���=r���r$.D��S�l��3���b�#�,D�8�Wly�؛k�u��A�Ca(D�h`f��^Jy�"��
Z��:�"(D�� �����d�,t���K C�tZ�"O�m�A)�2V�B��B����s"O*��"�֕p3���w�� �,���"O|��f䈢V��p���n���"OB�����E�¥C����7"O��J�#�.z�bŠ'.�BA��"Oh� �i@�}���9P��5|ޜQ�'��;�8��j�r�$(EjH	]�h��'���?���d�5P�<�v��
?Z�P �g:J!��M�:�z��FO�V�E���wh!�$�+�<��֡_
���:&f���=E��'��i���
S�RxѶ��%s$�X
�'t��JVA$�[֡J)
�r��}"�)��P�G��	��f�|KU����B�!��	�� w�x3������� �=q���$9�*�#��pK a�%��@��
O(6m�Mz�`��
��9vO��I��:pDaxR
�10x
�O&��hx�+���>��5�yr��)ac��{��7h,�%I�E��yGE�x�@�)7�CZ$4���$�hO"�dq���o�'6�p����'d�0��FF+ú��D�	/��m�%�;f�@y:P(��B�)�$8C��Q	+R0CtB��dP?�Ѥ�9�,{�Dʚ$�B���Ŗz�'��x¢ёm�%�jao6XCC��;pO1OX�',v���H�缃�ˋ�#\�5��-�4t���HA��<�����+!�xh�YDљ�D:%��	Ϧ���T?��<�m�������Պ|~�u��Cw�<�2�C/��S�YA�٣F	�q�<���7?nhc����P���	k�<��\�q�=���JR��R���(O��G��O�s�$;3L�ۤńpd�O��J��Mi�$͝.J� HS�ԘY��V�)��U�s�B�dzT@��mȱ^��*��)�O��Oܼ���\�UH�#N,H��"O�  �оl�J!�bBV�oJ)��W�&����'_���ږ��-XV�0C�TΉ�ȓ�n` 5D�k��P�����2���''�t��Ι�8}����B!a|���d�<�!!�
~��)cf@K�>�r|sV���<!�J`h��dF�FR4�G4�l��y�(�;e
Ԟ��1��l_+^۪��`vh c �I�V�L��K�)'||�ܴ�O���'��zdc\��4��a޺B�
�'c�1��J7l��R��y���K�І�I%fo���(\Gu� ��A�`�=Q���?�i ^)Z��Ż1���쵋�/0D���E˺L�KL`��鑤�G�J	a|�|r���ðH�=%<x'Eȼ�0>�K>Y���%�,-J!掛l]�д�Q{X�\��[�\�vJY6w�*0:�+^%D4�GD=�i��#~z`�	\��' P6&�����L�s�<9DJB�j���I6�ٳuq��c# S�HO��'��I��M+��T��Y��	HH�^qHv >`���7�)��<�vfݚɦ��GB�.W�n���ZJ�<��N�$P�+�+�(;���҅�C�<i�@J�F��]��C�.�h��3���<�.O���>�cA�u���X�m�(ׄ��$x�<Q1��y�^\��KJ6������p�<	A!��B)�X��/ao$�#r�nX��Gy�gފ:Ab1C$	߉^z,"FIS���/���j\ғF�/���r�G�78�D��� �r�U��FHî-},�ȓSk0����Oy��hU,;��oZZ?a����	Fԧ� ��PRh"Gܼ�a7N�8�D�h&"OV�;���Ĭ����xr��r"Ox�`�°2�����!A��×[�0E{��)J�&���;�	S�6�PeC��7/�>���>�E�%E�� ��.��n��Iwܓ�hO�O��8�&�m	20�%OW�*8�'�� �!,��_/�`��$}�zقN<��'ߛ֙|���˓�F�$��<���r!DڤK�
݆�z �8H�Fѯ-���TkٛJ�~��.�IL�TE}BDQ&B��� ��,`� 
/M�yb�#%\����ؚ��ɺ�D��n� ���$'�O���J���W��{���);��'��}b��>$��l��Uf�j�SW�	j��C�	��� 2��cT�Y$��S�C�x��Pi��ݚ���f� �&�VB�	?��p-����XH@ @�-N2B䉊#c����9Zv�����l�PB�I�L;�\����C6�)����|v4B�	� KH�)�� ���a��-usB�'x|i��%��j |qt�=Z"B�	�K v�+E�;���b偪1O6B�	iT�u��H�Sk�9S�^0m|B�?�P�p2;�U�@臼R'VC��'O�y06��7Y��y�7���B�FC�I�@�bE�m��oQx����ȩOv"�	��������A��X1̑Bs#K�5�d��"O�Ȫ'�A+d�\�
?1����"O�����L+@��2C��(z.z��Q�x��$Y��O�r4�fȍ����IU�_��Y�'B��)��H?+X���φ�H�<��'CfY��
ֳK�B)�k�?"�i�'�e�ԋ�6<�1�+V�ɥ4D��F��5\���f!W	O͆��% /D� j�7�PyK���.[Z0r�A!D�lW�9�ްSEm�(]Q�Q�=D����A,��4$'�2D�� ;D�h���Mz�0�O��IIƌ�W�n���$�	H�'b���Ц9�B��p�̳'���I<����i�68%�R@(n�|����I7!���,Q�B�i�JE�)��M���)!�D�A�02un�/����&D��P!�P}>.��fIG !"H�Pb�O;!�.':�'l�;,bJ]��.�/]�!�䇂$ŀ�jq!Q,�䤋� h�!���3!n82EI�f���ǳ�!��!e�����&l�S�s�z����p?�S�+�����W
<K�Fo}r��_�,c�"}�U��?0��2�o��Q 	; ��l�<1�-g�c���3������Qe��y|RR>�I�\$8%-� ɖ0��ՋL������<��N��1Z͓RHO	M�¹��%GR̓��=Q@f^-QM����(��@0�r�EL�<��MߔcV�5+O�^��"�DXR}B;O�˓�0<�gJ��]���ѱ�/]�Б� E}�<Y«@�jO�ؙrˈ2[$̩a�.{�<�0Bƿ�zx�d�>��y6z�'?�?a�#A(>j�H���5�\�"��<D�c2K@<vl�ra��g�N!sf.�$=�S�G�ЃNP�0�c@�˟~t��ȓ4}&�1$O(f���*�5m���ȓTc�QA�h�!:�	����B?�|��$B�B�K	?<��APJ��I�����I[?����#aVt��CD�@��B�N]�<9�̻~��}��C�I:^eÐ�IOX����I�S�? t9���.x�z1�ʁf"�[�"O���� �\���='����"O�q�K�
XZ�j�/M�|s%"O���!�n�i���J�q�X�F"OT�r�J��[Д��F
�lq�@�&"O���V)�[��ʋ�����"O��@��I�+*�i�V5^�6c�"O�q�$��#a	��Sŗ,��U�C"OL�i��L�}�Y#.��1���T"O��D#�,��T�_�#Āx��"O��I�*؅*�~�9�. F�VŊU"O�	�G:
�p��焹^��<r"O�A��D�;���3����`�"O��� k��zA�] �i��"OL�kGo�3=4��"n�*lh"O`�R��z� eq�l�=n�� "O��*A�_�m:MA��*�Ѹ�"Ob��b�I�*@T�U@�%W�d�Rg"O�����!6b�������(�{2"O�B���/a���4�K&��}�!"O������0m�ʑ`lR.0��A"O����<:p�	]���;@"Of����^������5E�p�#d"O��;��Ժ1��=�I�*E6Y�u"Op��#�([�:�@�5Y��|p�"O�����K�
�>e0�G� ~��R"O�tcCG7 �0�H/k�Q�"O���@˺2��p�]��*(0�"OF8���[H�i[V"� -�R�y$"OJY���6z��P���r���p4"O��� +@,�0�i��̓�"OVŲΓ�',�/��16�nw!�B�8	FIB�,,��Aל#�!���i�u�� ^����"��5E�!�$żL����ǡ��QɄ��O�!���
|p�\���g����!�@����
��5'�hk"�0x!�D	� �1� ��5r ��r�%�!�D_�G�\� ��Q��!����w!�dǽC�@X��C�/I5{-�02g1O	��I�5hh�C��E6}1�:`��	���F%�q�䤻 ş�)i!�$ڶ ��#
D#@8 D%��S�!�D��7�0Ex$m�|�n9��oU:�!�dKq�\x�������s�nͧF !�U�:%��9q Z����ف�̛!� �Y��8�n_+l�ƽRЌW^!򤜀E��h�V�GA�N�%�OK!�䁥B�9%�â��D�
�R�!�DT9��'G�T��������`z!��^15�r]�N��f�¥Y��Q�k!��'R<T,1�-i�<�yD�ڀn�!�&#e�pP�ͱn?�p/G�!�6|��y�P8�E�f�ٷp!�M<(T� �B+	�>�I3��!���#Xs�$ç{�NEH����
z!�dE	s��5Q�d�*�e��ji!�
8�M��ԉ��۳j@�k!�DD�H�b��GjՐ��1+T(�1CO!�D]0���pG�ߢVRT�JqFA Q!�����Pb�\ @��y��۷ .!�X�5j�)�D˓4F����I	��{r��<:��D�'��ZG$�	��ԛ��Y�= m��.ۭuEv�0`��O��ȓ@�&�R����J�n�� j�>Ihe��h�$zZqO��Y$ҽ,�"XJ�'� U��e�" ��m��Ҳ-�<�ѧ�Q�&���2T�s�|Y�����|�mzB֧�y��l�L�҄�/�ڂr�=���|��i�H�Ѕ�/�ۀq�9���|��n�H�ׁ�*�߇w�?���y��l�2z�>�Ηb*����2��.]ӆ2z�>�Ηb*����2��.]ӆ2z�>�Ηb*����2��.]ӆ2z�Dh���l��yDڦ�NAw�@l���n��{Dޣ�HDs�Bh���k��A٤�OCt�Fk��0w�
w�X�׷�;��f�0w�
w�X�׷�;��f�0w�u�\�߿�3��`�2-���1p\:��;iC���&͖�=zT=�
�<aK���,ǜ�9xT=�
�<aK���.Ş���Z�x;c��_�]��*`Y���Z�x;c��\�X��#jS���_�y9g��W�W��#h\���P��Rl�<�pwG��!��"^��[e�7�wrE��!��"^��Xf�4�usE��!��"^��X���:[��$T�dy�Q��K���2]��&W�`r�]��I�
��0P��._�mp�_��A����o�7�%˾6ޒ��6s�M��n�4� λ3ڑ��6s�M��n�4� λ3ڑ��6s�M��k��ò.-2�����e��#�;��ǵ.(8�����m��)�;��ϻ' ?�����c��#�7��ɺ�,}cY�Ot�r|:�g����#�,}cY�Ot�r|:�g����#�,}bZ�I|�xw6�h����$�(~ԝ"�� ��T�i�f�rz�DNޗ&��*��Z�`�l�|q�OKْ"��+��Z�a�n�u�HCњ*�}��1���[�}�|{�}��1���Y�u�qv�v��6���^
�v�ws�u��<m��A2��(n����ы�;�e�E5��+n����ӏ�>�`�L?��"f����ӏ�>�`�Lm�_az��#�_�h��wu-�b�Sjp��+�X�o��yw,�g�Wgr��(�T�f��yu!�o�ZgM1u-0Z����w v�2� J7s(8Q𸂋~&s�3� J6r*9P𸂋~&s�3� H5w-�P�ʯ��/Z��Ȋuf�ᬵP�ͫ��!Y��ʄyi�כּ]�����,Z��ȇxn�믶R��wD��E��y�m�{h�h)�3�tF��G��z�n�yj�h)�3�tF��F��|�g�rf�a#�8�~O��Q_{��q��F[���53d_Ru�|�s��GU���71`ZUp�}�|��A]���8>hTX|�98M1t����֖<�c��Y98M1t����Ԓ9�i��S24A=����Ӓ9�e��\<=K6�K�b!b�����<���sk�F�n+h�����9���yc�K�`"f���
��;���d�L�e2c����]�"3t�����=9i����P�)9r�����27e����X�'6p�����<5d���%Π�>���X���ϫo�熏!ʤ�?��P���ʨm�〈)¬�7���R���ʨm�る,���.K9�W�I�t�1&���'@3�T�@�}�3)���,M3�T�M�v�>(���	'��Mم�s)&����ߏ����I܂�y#,����	ޏ����I܀�~+&����҂����Cԕۙ�^�Z>� ��������Ց�[�T3�,	��������ג�Z�\;�,	��������ڙ��"6}�z�����D$ň�~E���"6}�z�����L.΅�sN���.:v�s�����E'���wO���(?$����7Xs�E��=Guz&Nɞ)����5Xr�D��8Cvx+Aǖ!����5Zw�@��:@s#K̛,���߅�C�����X�Jv�rЈ�I��˴�\�O|�x׏�N��ʶ�X�Ix�w׍�< 	K��Ah��]
W�����2.B��Hg��]Q�����:$
O��Dm��XS�����8'HjF��FɌ"�d���1R���q`O��C΋%�c���>P���veD��AΎ �k���>R���p`N��&���]���<N����"���W�
��4I����"���T���8B��	��*��Ԫ��R�ցQ�gNu,�c�}.ӭ��X�څP�cK~!�c�p%خ��S�Ҍ]�cIs+�g�r$د�#�<:ۓ�bHrQ����Z���"�<:ۓ�bJvT����P���%�;=ݕ�fKsQ����R���.�63���rV�6�������U���[�;���ʅ����P���qV�<���ς����]���j%bv�'�U�WܕcW��K�?b-jq�"�P�SߖcU��N�2m-k|�-�]�Rِg\��G�:e(n|,�Je_����~�,�Q&����(�MaY����u�)�S%���$�BlU����v�)�S%���$�@o�+jc�2�A�*b��Oϣv�-o`�2�M�&a��J	ɪ~�#ai�8�M�&l��AĪs�-ng�ʥ_@q��M�if�����ͭUK
|��G�nc�����ͭUK
}��C�kf��
���ϯT�<6����v��x�!�EI�x�5<������v�/�OC�}�7<����v��v�+�IG�v�>5�P+x�b�n�T1��pэ��P+x�b�n�T0��sҎ��Q*y�c�o�W5��w֊��U.}�%8CE� +'q�,�e��"9CD�$(~�,�h� �*6KM�&,{�$�b�	�/U0+�5}��q���� P5.{�7|��q���� -]8,y�6x�{���)_9#x�L�W*�'	�� Ω׽_w�A�U*�#��ͨԸY��J�^ �+��ͨԸY��K�]?��>�>x�;���~&V�|R3��3�0v�:���v,]�s\2��3�1y�;���w,\�wP	?��:u��k��PL�C��T५A-�p��a��]A�I��Q㧫A-�p��a��^E�N��Y믬E.�r��`w���
�����#�䃄Z�{���	�����&�烄X�|��������)�Z�q��_�,� �عk�9}L��_�,� ~�ܼl�0wF�
�Z�)�"|�߱a�4pA�
�Z�+��?N���=xJ��[�ú���5F���;}N��R�ͳ���5@���:M��X����
��2�Uէ���r�G<��2 ����^߮���u�E>��<����Y߯���z�L1��= ����Rӣ��~�X��`��!�Y�ʕV|��q�T��`��#�Y�ϓ^u��z�]��e��#�Y�ϓ^u��}��򺉓�,�����ھ�̒������!���Ա�̑�󽍖�"�����ݹ�Ř���&�e�9��E(�C۾�SnT#�m�2��H#�Fؼ�SnT#�m�0��O+�Iհ�_bX/�j�C�L���a4
�� ~�ռ:M�M���f5	���,p�۳7F�D�ʗn:��$x�Ծ4@�D� �@ ��	��-�?�sG�/� �@ ��	��(�7�xJ�%�/�O,����$�5�~L�%�*�M�c8s�����t��%��w`�x�i5|�����y��(��zj�r�d;~�����y��/��qg��n3yA�Uw ��-!gH��wTS�[N�Y}��!-mO��xPU�YL�_|�� .jD��zPT�[M�]p;g쇺��P�������T~�I9d脸��Q�������Qx�@3o䏲��W�������Qx�@1l��h���r`� 0w��)S���O�o���t`�'7v��,^���H�o���uc�#0w��+\���@�b��&�q)��54٭8x1�,�H��"�v!��?>Х?}5�-�H��"�v!��:8ج5v9�'�O��%�s&���F]�04z#��9���1����C[�75y'��?���1����HP�><t)��<���=����G�X��!���p�����vG�X��!���u�����~@�_��$
���}�����{J�S�G��%�"�MK/��Q�B`�@��*�)�G@$��^�Hj�K�� �*�GA&��[�Om�M������t$o�:�SF�{2!1�;�����|,g�2�U@�p;.;�9�����x/e�2�[A�}7"?�;���� ��!M�3�$���cG�ea�TR'^�4ƐCS;>r�RF̥t6�cC��5�4��K<I��"I8pp%Ϝ�m=���`+СR��Pbd�P��e���	�r�`I�#H8�	n:�����"U
���$�A�I�7$��Z-�pΈ�4(�0$[y@T5"��e䈤O��r��&��A�S �|CdJ�0�IQ*C������͆F������6Hz ���
��X0t�@ޟ�aj&��	�Xw�2��V�=��� ��2c��p���jѥO�P�aa�H��cgԔ���#�L�$��� ��9}V0��
����$V�����C��"ɼ���Y/Bf�I`L�>;l�2p,Z
	����Q�V������  ���#�S<U�*|��#�j >**�;�a 2\� ���GI:a���sB�W�Π~B��Q�Ĺ婃�0�+'/�L34H�.��_�$6�p����1��-�ೋR?�y@�N_����mG��i�m[)Mz
@�$�ӌ/z���d��֠��Dg�O),�Вg�m@�ם7l�8�p��H1��GZ�`hD��O�-sS �@U�m�EOU�~��G�@�@$E!�'^���8+9,>CPy�F	�?P���s�3J��� XϬ|��`ѷe\0�T��y�)�e��ke���1M����[ȢX�& �4`N�e(�2�:e1����4��d�I,\����'��  !^�nAt�J�gk��Z��)&$�V�X�H	0a� Jf��B��uj�l�
0��<C�K d���[jߤ"�L�S�ɱf� ��=F��n��R�>����!_�9����B� lC]h����Ս"[��)�,]�F���2�ѧ�ZErR #2� (���5�� A��!�B���Y�Rs�L�ĵ0� �"1�*4�Eiē2��<�'��("�
���RS�!��)�!��}( ѲmXu��?�(�1��FIA' %;���<U�h�𠣕��\���^�H���jƉ=Jq(���6/��I�d �>�a*� xn�M�/�'���j���,K�ii���C��YBU�EH�z�	�<K$�%nR�p,�T�U�� ܮ �3�ã�Ms��ĜM�lу2$����'��=+��u�0ޏ��C�Z�\a�l�e�h� U�UZћ��	C�d�9A��a`6��7��1�4,�a�V.��y�f}�R�� �p�y1���``2������E�(4�r��Ab��i�46J����ߒ#�vy�� �N][s�Y���b�]�<�o<�B��oj�1c�@=�e�f-0sB�����3=P�]g.��O~4�pӽEp��I�
_4b=�f���>��'�G��I3���؏@�AgDB�K��3c�C�M"<�b�N�h:�0�n�1B8(��.Q�0��J~"@	&Y��Y����ةm�����G��F&9R�$),��#=��m�x�jq�#�M��9x"	T|�jI��Z�?�rY�FHA�d�4�4L�l¬�&�l��N,܎Mc�gn�O(X]�@�o�Z� �ڶ45��р��%!ҍ�F�D
ER�I#�H*^Q�`���X��kLC> ��{��$G�a;�	I-T.XX�3�J�f~b�'�X����ɶ�ا%�V�x�'�|���?����8!��P0װ,�H�� �8o;8���B�������>	��=yぐ�V�Q�v�	w���3ҍ���\aeA��jf���xC�E��Fá*��$�v�����72i�aȗ-QK��#��(o�4ekrχ3�j�Rń����>A"E��}}�q)'Aפ뢨�'U�D��g7�bZ�-�n�yRE
�
pI����%EЮ�(�ۼ�0iJ�5���W�Ĩ-�|���h<��^�/����F�%�NI�a圦h��͂��lw4�bU�^�q��K�.,�����璛'�J��\�j���D�L��F��ţ G����<)�-͏S72-��!���ܕ@���4ev�R�LM9KH|�A�`�D�X\+1�G�A�����R��d�D4`x�=	��FFX d��O�X�����|�;$� �2���|+` i��
�*�kb�)2��ۇb��0�uz����+*"!A��I	-X�I`���c� X���'A�<�F��Z89����*@$܂���n���	�ӒY�|����kL��Ə�R(�M&*E*�ҞwBf��s�A��3 -~�K3$@�9��|2M�+�o�?�����'�1��`��� �o	�{~�- �LϥL���a��r�����7��@����8�'ɼ�8�� :v$	�v��)P���"b�*��u1Qn�u�8TRXح)�B����ei��"i�(��@֙P�Xh��8Ī�A��O�k~�QE�� z5��&n� Fz2�E``�J��S v�h i6I�f]yT��|z<(U���@U۔˗Fgp�Q��W)b�0�	ԴL�b]qT���R�2M��GF�JGЭsѦS#3f�u�j`���I���Xj�A�'��XBa)�z��7��&@�A"q�щ!�@��z��Tj�aݧ�� �)�j���O$)<��*��ØKu�Ts�*(�X�����2�R�J�������#�i�A����S	�Sr���-:8��� �
*?���� ��x�:�ӃiB����㩏�Xf�g�p=��j0�H��#M�R�Db��Q���V�P�PG�/�4�����6��j>,z*Me�ã
#dNuj�b#5��P���Ѥ;;� ���%  ��N�J���l���x�����IK�d�gă=Z�<3!�F/��4���K7��d^UFU9��ȕi�|؇��|�|��a��>�X2��X�l�`��h�=-(�/��PFBہ;��9n�0��a��oz��bEB
0c�~$'���jd��� 6�BR?����9Y�Vd)&,�e::|�2a)�ڹ�a�O�f&����O�'9��ީ�ޱ�Q
��b>��Rc/�r�ײ=���h�n��L��� ��҇r�j������[�i���X���/dy��Q�ܿQ�i���kLYN��tؤ�"�H��͘�	�vp�4�O�
� 2�Oh߂y� ��HˤT��kP�?A%��(b@,��y� ��"-�$�3G�� �JA�Ǭ�b�̀:~��h�.��#<AfIN�n���H�l`�4�oF`��L��JN����VF
)��'����&�ʓ*�|����}�4\h#(�;��t�6��y�����0����w�W�']��1�Da%�1�С��G�`�z��B4`��d�O�d�`D�x"	<�2h�S���a�3�X졡������r, �!�l����$$<�	Z��-�I�x�x9+K�u����4���اh@4��ph��Y�h���+�>~	���2L�6/�0Ԁ�*:~���׀�=(��A�"�Y�l�����<z���R�6�yE�����Ң�Q�vm,8q'i^U�(�g/ج( m9G�r���q�}�����O���dO��T[�!^�He�P��L�����2E/B6p��TFH��š�H�+V�2DC��IgQ�� ���7`�=/zN��l���b��;}vћB煚>�p}��N<'����W�x2C��{GHQa�oA�s���Ci�=���c(�Fj<��'ٸ9��}���/%�8Z "�~�!vB>���h�k����`E�M,ՁC*	�d��z�P(���U��jX#^�����8���k҈@�� ��a�M�,��}"�Ҧ�At��@	\�����mP�@"'��|"%��kx3 �7K&L� #�ݟP ��@5
rU�4"��3��ʟ��F������^R>�۱D[�Z�����#N{�Dڥł;G���E+�n6�̰$�M$_P���ͻ1��q�
�-Wj�",����i	�!m��B%,q�<eI�\V���D
,q.m@��\-O���	��.���R�Rg�������F1.<���̙��9}b�ɔ
wZp�!	�!�\QB�ᅬ0=#���Z����'fJ6'�:	���~�|�K��-��KS�L9 ٬x���9Gt�CI<�TO�r�,䂧�%����`Vf�#��<�$L�\⟌����
-'�q�A��tO@�9R���
��N�q�#߭��`��'�;�0�|�>\
��*�)�'+&D!�����;��(4&�"��!�B"�)"�sAʉAd�L���*'�>�][U�Y��QN�N���nT��C�I�b!L�pu׻%_�I�K�;cvP	&�ԈW%t�C�%�F�n�f��?�=�$�ٜ	�
4�喝+n�Г&��Mx�ԛ�IJ�����*Z-uz9�����Tp/_���JG��c��X���A!)�赻b�C�!� ����;�����Ǯ
�T��z$qEC�|R�Y�p	#"�"�"OX���d-[/L��C�&D:-� "O8%��"��
�yAĎ*v0��
�"O&a:�$I0]8�cC 
%*m�C"Oq�-��%�$�>8)2"O,��Q'�.c���6��
{�l��"Oʈ�u�.i��}��@7H��t�"O"M���vFQ�u�Y�?��y	R"O��p��R���S&�%�V%��"Ot�d.τ�&�xs�۟K�����"OH����u�\u�Sc�<�Rd"O�`���Z�ܘc� 	p�"O�ٙD��EF Aㆇ�_�dݺ"O  �aC�T/��v%U,��z�"O��pkɫT��yDA#"i�Ԃ4"O�|��i�/pL�L�4R�_JI �"O�4���Og�v�+�y�h[T"O@Й���7�,Pх��.nH-�f"ON��@(��$��D�f�ؓ9S�XS#"OxؐŎ�ZJ�AP��5gX|��c"Ox��a��MZy�u�P�U��hr"O:�ғ(�L󬑰�N�8Q��Aك"Ob��2D�#T`ځ�Cb_?{>{w"O&=hf+?���T�&4x�"O*<r�K�
J �u����G@�r!"O�E�ްޜ���À�Ľp�"O��+c�W����1Q.�@ĐD!v"O4��#t�I�N�=;J�;%"OR|��׷-*�eC�kǤ����"O4�����i��jB�^�b�.�yR���a��I,5�ؚƆĴ�y�B���BfY�̰����"�yb��<&�i�FԐ
�ސK5KE6�y�(=b��&�E4?�yEE
��yҋM6]߰��J0[��,�4�1�yr`D�cj�����Rh�����yB�^�LP��)ن,reR�e�7�y��^V����̊~���s*��yr�P�t������)�F�떌8�y"�q��$����V�� &���y���N��H"��>F'ެ��IU�y��TR�m:BH�<:lTi��)��ybʶ��1��)�����y�Jʳ+.�c�o/����N��y�&&*�����	TM�0!�4�yR��m7@p*'�9q���j0Mؿ�y
�  ��2i
�b=dY�r/�3\�j���'��0�ō�p}"z��Eŷv��#fA�w�tաg!N�|PV���?`�j����Oj$IЁT�`�������-4
����Ė�txfc��~2��"O��0P�C�Kx(�b�?3��L�`���<��+#+��+éO� a}�!�.�h���J/34��M�9L��
�֙:�R��.s�Z�˔�.�`����C�11�2�M9�y�"�;xxf��fa4��ex�
���xT�Q����CJ�0y^�e�-ִ,�H��k�>��	���2�h]���T�R����3��1{]�a�m�.�D�;���B�葊��0"��2R˘�s�aykcBH�s䤗���=�C��2ax���po�
rR�r��id sf�O��b��@�����a�2b|���o&�ăd��੕DN�P�%��E�o�]�D|�$sۤ1�D��}����0CJ�eY:�hg�[�NԄ��'+Ȟ	�tY��ʙQ�1x���O��9�WHV�\h��A5(Q�v��	!X�t���fU�EqO@�p�#�;>4�l��mG�W�dᚅNUq7���##
�|�"���[�T�0�#�9;?�@�P�/S�x��%.���św`H�W����AD>������'�XZ%@	�kL��@�'�����28L��sd��7~��u�Ā�� <��DZ8B�u����L�LKñ<E��Ԡݵ|��i��ϗ�2óN�:�,P���_�i���6g�u�џt�ڀz��=��$۟doڽ�g�ΑuW�ܨ�e7�m!f�h��5	7ʌUjIA \f���ن��rW���A�'�Mq�i٘n��	a�E��Db�J3Q�v����2��@c.�W�N��5K�|��hj6h�[j�-B�N�\T����h$g��8!�B8l��4A�Ⱥ��iB��(�;��۟�m�71'B*�q`�BC3�(�A�!9�;&�V
���,U�R��Hؚ:���+���b�Z�0~�����HQ9"�F9ZP.P�N4�wH�>��K�U�~���Di�57����AG�5sV�)��O�`m+㋘qBU��}������$U����YCM�Y��� W
߫^w���BF	5c� �]0�p��ީZ�ȐB�H�3n��U+���M+e��V�$1s�M�x2�iJWFZ�4t�$r��L4V]���'���-�PsGɢ�ēL��\31�O�C�
�ɶj���9C]0��ј=�r�WQcĊ¨^��Y��(J�lt�44G� �ҵ+ޕ�����ˇ�KZe
�[��1��Fħl"�Ҷ��V��T�7� ?!��ÊW�|�POÃ%�܄�M�Cٛ�J,&�Y�d��(�h>��=�	��.�P�n�1)�����h�	��3a���"�	;���0�ܰ�0�(6.
�,�q��
��x�M�g�Q*�����%[��]#�7O�� i�L�i�5}�@� E�.p��b�-F�j����Ę]��Qz&(Sr�Q�:4BX1P,�6a1��B2$D���#�͌qc �0?i'��0&x�seJ)�^��4��*I�P�Q�F�R���rHL�ڡ��-�1+x�C��(�@���͜(L�@�	�BF>V]�aYPWE�f��7C��h	Bq��]�bM TM׿6��.O��E�7[�����EX��:Y��e0���p颤�Q'�j�f�Å	���diW�	z���F�8]��uP
OצMQ�Î6U۪�bw�"��P�2
=`8!"$�.���'�:H�a�I2�4
K��!V�ӓ#G���X-'���`���4��7�/A5j��Ǐ�
7vi��`��~`�2d�ֹ}�h�83�V<��G@ƮB3`���/�5z)�^lZ��6,G5:���Y�8&xyؕƅ؟\+�P�<��	�b׆XgN��fLG�<%�i� :"K�cny�w�%��i9��_����Bv���{H�Yr��X���%��.bjm�'Z����#����_P�a�J^0Hh��*�5�v���e˩���٥�ŴI�(T#�W�yV��:�ʛY2Jp��B4 �~Ͳ��(y�6�f�Y�t#\�p$
�R6 Բ��S�eL�q!��	C��;-O�=	��݉W,�:$�������|9f	y��BII p�đ;��	��#p�$И��P��H �3
_�=dY�iC�H
Q`�<���C�3P4t�����X#����Ͻ
�˓�j�`d�O5:�8Lb��T���IQ9���� �P1U
�Y�rD�t��!B8Ԕl�1ǝ�,N>���@%-2�C-Iv�i��$��
\�R��=ބp����)D��xb�ЈIe�yR��W��0�z���#Q��t�Ov�x��Ԙ>�T��(��6�6=P��S�^�����.k�`gʚ�c�tm�'���Aڼ�1�&� t��)Z��{�̡�-�fc�0(Ǫ� f�fM�O��q`N`9n���D��!pl<�T  ]��X(��F�F<�Kb�Kb����e3z��Aē�${z�f��Y��X փ�#pp �+U��*`R\9���!B�g�9T���r��2A�'��a�EL�(`�p���OXdؕgϸvt�� #�;Q��Xp�;�GP>l�0�:�@H��Go!&g
>h� N��Rl��G*!�$�ie%Z1�yZt��>v��'�qBD�_��5�Z�@;�@>L���㗎яVG8��q��5T�̄#D� 1�a��FXC�n�;Ek�h�@�����nE6P�بK�F�
4 ��э�\8��)�Bd1�lA4��10�Aʒx�:�9��O���g�:_����!���	�[=x�
����H?I�"�+3/�<f�"�53t�ĭ ǭC�0�b�C�C2_�=KG�\t�.�k�o>`�6(�M<y�&9 m��G���h�@��!��2l|�cfX�~��=�� )�U`#fF��MSįt�]C� ���"�qÃ܁4�"�� �J'̍�C��*�1�f�B�*�@�a�]=�B�aI<�$C�:7r���C��3$�HXX�a�;'�ʙJ䧐� �!�#E�V�3�ܩE}�cR�Z31=��C
rLT�c�"|L�i��ƈf;��I��U�y���f�޵w�.,+r��d��'��Mp&�S9 8�rC/��>�dݫ�n�aO8�;��T��ՙ,��Q�aȃa�B!���*\�B��2�؆l�(8fi��f�Љ�5��)��u���b�H9��ܫ^�L�� �/O`09aC�4U����"F�W�պ��S�<�YsE��o-h([ŀ_-Kg>Q�!�1X�����3V	���T��>Kt&���-����Kl��Ad�a�F0�B�l���d�>N`*vDc����~5܌�SO�&�ca/D�{��P;V���M�Ѥϻa/�6 �/#ےU{3��<6��a���?
��z2M73)��s����ih���x5ʈb� ԰E��y����c7 E�g�,}�#�8�z0�o�T`�zv�-�&$�!�ŭ��P�Vd*SYx�8��C2Z����H%jH��BE�u�, ����/�T��[+PYz�HG�°ynx�UOI���|Q��~�.�k�O���҆�4(�:iBw�)����a+`�L��4N���Q��/�4U�$�ԴC�%
<�r�2����2]µo�CR����,,�pm�w	s��7�P-�p���
�Y�A��R'�u��$ۈ�B}�A"�+9U4]� aZ�E��ر��4"0��C��%�A� �Z��XI�1B��8R<iZ&��!�@)�
�J�"v�dq2�1"�	�6�l�Y�"`�5LO%7,Rq �f�$XHi\tD��7H����H+k��l�j��M��扡Q�xA��K!^��	�\l�ΧW�����ԩ'��d9"��u�(2���UxI���La&2�	�,� '-T\A��>�#�فEGN��2jN Mw���Bl�g�? ٫�@���je���d�,�����H��*����o��'�p��"P�K�4D3�̐�V�z�)�Kw��"�L�W��}:P����������Q�* F�	θ]���iQ�_=I
�$T>-���gF���yQ`�U;&�l�Ȅa�sa�bQ� �L�;OGJRYc��^+�YشsE���!���h���s5�K�C��aQs ˝}x}��G�e+�t �1��yP�%Xv�yQ���F��I� �{ti�%����th��0
f8���H״mL5���lqh(���	X�x]��������F'Ƴi"��5��u�	�f�Ir�A׈H����C��A,��h��]�@t���aΨ^=���B�P��Az�1O�ʅ�܏G#��U��EXu��H��_������4��!��K��t-���5��'�:=��k&bL[�#�J��B��C�Uw:0�ŋ�"['�(�u���$ 1��� Z�8�5� Y���J a�O<$�e�� ^-� �;j�D� �×i:u��z��@��
�wp>�'� ՙ���f��H�"C̥*�dq0�+[jA���,:�hx���X����"?� JJτ"c�AK�%�K�j�a#ȣ��|X��4^���dF�'2�4�
N&k� �C��0&���>�E	�@�<���x��Ct�dY���p�0�K��2 �	�_?�C@G�\�Ω��GJ1�0�r��W��4��.��<s�6CߥX@�к��Ӑd�ة3󇎖f;�}�e�ʭ�����C�v�y��E* ��;�-Cr�8��W�B�L�b�@I?V��*��#@��2�rO�?���s(�8Zud�N����)���s�.!X�'��^�|hHAi�' ��o���d�
Hv�IPΟ:}�����ڮ!9��K� \�&�,I��:g��0�?%�y*�Ӷ'�l�3&kP	'3��;B@�$"� U;bN��c��h#�n0$��b��[���ؠO�Bw>0�V#By}B�~p�<�3�@��qq/�,@Dq��d�h��k�¥p �06J�ً��y�V��&��	Zkc�[��H���U�n�ιH`�Ĳ2@���7>��9A��G�F�`�&�a�сDDJ9*X9Tn�Ukĩ; F�LN��g��/s^𠖯֢������/m��h�&꞉l�t�@o]�>f蒆*H�h��������ـS!��j��\�'��:VE	P����VlٌG:Du�JB.`]0�h���n͘�P�#��?	�eT���ٶ,Y�D;L]AC��fR*ɂ׌;,�	"SN�"@���ݒ)�~ِ�b�7�nY؀:}�����׫�����S��ɕa�t50�e�:t�` �(�)l��86c����7�@�FLFu#�`���0�r�\�z� x�4o�
�`�ցGP�ɒˍ�z7��6䄖*o��(�#ڭh���6 "�t1�FF*�|e����=���9@m��dv�(5� ~�>����\���V'�T9���+;�)i�-��`x|�85À��8���1�и��(�GJ��;�#��\���(a+9�p\I�DN<�?����
����ɛ<��)3�$î~�P��@�T���hS�ܲAN<Ĳg���RQ�p(H	5 �!;�$C.�\�������DI�g�P�����	x�����IX&��\rh1i�Y��hO�1��;{�)�"��44C@ C�R�O�=j N��~*TPksd� 0�$��dA����}�'aEr�	B�Fʕ���ʦ�!���;&�*��e��5�V ;��� A��M�5�%H��s��X��O������
,5����-�W@^����O�	0{���:�m�0�UE��oD"?Ȋ�F���H�k�(�D ��LolʙI1���L����">ʈ��=�����P� ��I�: ��߭b���P�IϏtu�D�#}��^���~����#Y��yB�E�J��t�B�ǺU�c�#C�P  �ԟNp" ���Z�::�z���N��$BRܓ	`�I�=7�D�phɝx>�m�I�|� �{�i
!�CoG</�X��O
L�0ȉz9�E�@�)+�DuX3:+��U�uᆂF��l��/Յ1tZ��
�z,.P	!�ʮD9.��#f�D�^���7��Z��'cx���+y+>xi�C�-C46��SƁ�D�V��;YcȀQ�Ix�N�RR*�6M�u��p����O��L��T�6a�4��`W��?��O��LCF��2K
x��"�N��B��d�� 8���'����؟q�ƕ�$+L�Z<���?႙#iךe�j0JGg�<�l"���<KQr�0�g��(���
B�ȧb�$���e�t0��JX�%}�d�h2�O���+�܏Y�,�֤_	;8�%�\PclI= `@hCI�6~`$���ф7ˈ�sa ��7�a��`DBV�R�*�>|�j�Ŕ+ R�aŐ)4��}�*��z�� �6�I� �4�x�I�)$�}(��C�F��pc�����:R#�>�A����y7m�$=I�,�s� )!|�r�
�&�p>�Ջ]*U�n6-R8��@d�M.��m�O�?�����E�����oٖ0����#�,:��4 �-��q1CK�;8�Ī�\=t��ު2������A��� �?�1�ޚa�|����<T`:A��@ ��9�KG�j�� .ox���a�Jjf�h��dc�1�hP�����$Ԓ�bfQ.r��t9�L�#����	�z�x@�ga̞�R���P��d�竆6y��]q�ٜ'���KeH��np�׏_�&9K��Q9d�ܤ��ݷm��M��*?V.�{�mM�_�����(!��P"1��r掙�-Y�}�H�R
L�#��K�ێ���T�$��P2!�ؾu떵�YD���Q@Vʅ������ӧ�Z�D�hu��9\O�%���Q3^հQy��& 9a��Eb���ČA�T:�!�!S#MXԉ�F	�H�`sE!C�d )Qb�Dj���D̀4R �q��%�ȱ�֡�-#��riI3}�t1�y)I��d5a��])k��"�/̠E��(�O@M���ϑ3W�9p��* �a;���-<�i� QU�-�R"4g �q�bcN�5Z�DxD�P�ԍ���,��aÁnߤ?yR�S�/\
�-آ��6���0�+ ^�j5����N	y����#Q�����g؈]��i��	0�j��|$џx3P�M&5�a�	<��șP���uB���'<<�$nV!=0DQ�'\?����2I�|-�AC��`(��4�������V�I�l'	�� �)��8��V�����"��:И,I9N��bgB+�����bcX�x$�UڦEHs��8���kC�͈�v�r��O�0H�өν3���X!X^DѰS�3������j�Ҭ��%�9����͍>q����VO��^SR��#)��O>1F�.�B�c�O�o��Li��Эa�d���N�<"��)�F�L�C��r�W/�R�Gxҭ�6M8��
�b�*HEG�_�HA�d��F"�) �
� V�|�O�%0���U�v0�u͔5H�P$#��خ<9���@�b �Go�4�Ŋ�Q��hO>�٥��@��#1�#C�V(�A�� ��X��N4�(,*%��$m�Exd��	#9��H�m�b�QҦ\E�J�� �q�1�M, �&�I�$��q���	��D\�df��g�F
2����P&�H��]*�&�*|�|��p�K,tL`�����S�r�������j�d�<>�>}Eh�)i6�E�0�,tNf䃳��W�b������c2k_9OØ}t�L�4&~���[�$�汣��EMޜâƣòUXB�8M��y��=�p��Od5�Ј )=��d*lpP @�������#�%B���f�l9���� �(Op�[��T�P�
 ����HǨl `AF� �Hc5���=Vx\����v�c��x�����Mƹ�N����S�R0H8@�
S������j~4�sae�hO�2�U.?zdH�"ۜt����W�U�z���)H��4��ܞy]J��I��y`��89����V�0�!+%��?�Ya�<]A�J��G���*�'�[�1���IQ�Q�l1qè �R J3ܞn�i�T}��i0 ��Ԅ�p3� �~�G_��l��4V
\��G?����o�ʧ>��I@/
�x���Y񮖆'J�9� �� Ӈ��p]���şA�
���C8�b��핈ܢ��!L�?MܩFa��y�mZ
zΘ���c�3ʓd���3S�C�;U�t8��G%�,Fk�3�4���%̅�dx�qk ����O���ɏZ 0�e�_[�T�֤�8	����R��6����	 uX�țue��i�h��V���;�O������"��5 �)��:�:��0�.��u-�y��!���O�RƠ�=l u"'K!2K
|��R&��MR �Ռ@vs� ��NŗA`��O��J�<8�����ؑd��*O�娆��6⸧(��鹓�^�N�Pɉ�kE,���i��:��T�Uk�Z��bk͞t���E��wָ����+b�Шb�$�\	�'��LX���OQ�̓�������M�T�l��$%<Z܆��O����љQN|T�qቜsPxS��!�}B盁#��$��EF�ir���<�<��%H	7
T@T�&VPa~R�\;��)E�Ҳi�Z1�B����Oī�T)Jɢ�bM|2��/�B,33	��8Q�an�b�<Qg&�/N�,���+SFT$��/�G�<��o,�5Z�/��M��õZ~�<A����$(b��ʞGJ0�;�'x�<��eW�+���iR�RJ� 3f��o�<�FD�W�:)�V�W2��9���l�<�ǈ��"��p�R�)�HcaeWm�<�'�V�H/*�(n�� �Dk�n�<Y�GC?m��L��oS�;��Ʀ�]�<�ЃH��|(� ͖o�P���Bm�<QT�0��
�F'��l�a��p�<	עݤNJ�B@"��)���e%i�<� G,D��\�7�Q<�ʴR��Od�<��ō�6ǜ���Z�%�z��G͂]�<��LQ��D�X6;z4y��ܹ~�!򤞕t�n��@E�a\�=JB�R
^!�$�5o���i�[*�Џ�0O!�DQ75��0'FQ""�8r���1,!�d��i��y0hǫ@��VDћ!��ޜ8gvŻ0��PD�@��e
!�D��`X~<�4�N�P�4��%1-!�U�9J6��b'�Z0���1@�!�D4ް�a��Vڔ�ِ&J�v!���[��wIV�1�D���&y�!�D�(v�1:v� �`��\p�j�"O:�at*K����j׭�>_��H��DH�X��tcGB�A���AOZ,q�1OpP�WB.t�V�q��M��x�a� G%D"�J�M5}�.!��<����2.*	�eOI�H��a��#*��'3(��>��EH�ܡ�ٸa�D6a0��O9}b�^	m�dpw'>�Z��o�.�a��k��� [�t!�(,t��X{'�>��<%>��`�v�53��_?6����&Eu�h�"3O���O�"��@����C�C�r��q@������3p�qO�?��� �����F�>����AEZ/Y����Ox!9��t>��Ǭ�<_X��k��F��t�hFB�[���<=(�Ѭ�J>��R۾yȀ��yѬQ����>����<�v�"}Z��~
B)q-B8+��P�ȰҁĦE -O���O?7�ϐ �.$I�^s66a�B�7'����HOQ>���̙�4u�U��{����O�MDz��iެ)�.��N��r�����$��|H�#=I
�'r<Ոe�ǵ�T��d��8���k,�	�?)��ؘOX��>��U�3�īq8�2�#�4����6��a'\����M��D� Da�J
���GFN7F��Im�(- R�ԟ1O� d1��Q�]|��#�K<S:��"�i_�=B��/�)�2��5�&&�3
�r5�p�S�sM�!"��C�&����\�d�arD�+[&�P�MvqO�P �O;��-��O�dX������7^�~����yy��p��֋����S�O���Z�b��@�ǝ&h�U� ���0&����S�O���Z f�f ��f$ ,�p�d��O�����?y��QZ��xR(nxZSBf�I�e_'���I`y��iH�.3%x�/C5�8ċ��
 �!��Ș2ڀݠQ���5�Փ$!���1@���p5��h�t�ۥ�Һ�!�۷=G�ebGi�F�5R�.V�I�!���_����S��9ᤍD u|!�$Ԣ�� ��d��L�W���W�!��jA =yŅBU��	s�~M!�S�K�bM;���$����Û$;!�W�yG�t�"N�-f�!�¤N�-!�T�B�^�BO�0mYX���Ü��!�!7f���5��@D0����7U!��m������.b��#� pR!�8|��X�V׎:D�����u5!�D	�=F���Üc$�	�T��g/!�$���Ι*�G��r�}Q ���!��J4Q���G圈1
�`�$Q'�!�dߓ	}����*f���s�֨!w!�D& erl�r�� ���s^!��+-��e� \�j����g+!�$ٖE6p�I� ������B�o!�$X��`�rA�2|�h8Ȁa�8!��:^X�8� �r�D�#���u !��6V�����̂p����lY�O�!��&j��;���B��Q)3�F��!�d�q���7ۜ}�*!��iA?�!��/-���&����&�B01X!򤃖gʎ�3R�C��L�ND!�d�;wJ���lD7m��R�<!�$ 
5k�@y1�=$����ME(1�!�d��s^�p�M��7A�-9�/C�v�!�D��~�����3i:(	��ci!�d(d�Ƚ��$ؐ�\�i��*T!�$�:|��-�&(�@���x���!�L&BOܠ�5�0;��]��:���Y�q>\�:6=Um$!	BB�y�]�uy Xf*��Lp�al�y��Z�%�l�j�n�;f���#��y������Ak�*TnrR|�0̎��y���	�� �UgJ-l�����^%�y�&g�������U��q��I�yRj�?�@[�FOb%�!��y���S��8D-R�oP�mk��j!�'��X��
��pQ� a�O�}Zj��'�t�"Pz��G0P�����!D���F@R
��,h���lJ$q�J!D�ti�埗al��wFS�`�Ӡ!*D���RK?��8C n�(l���I_<!�Ũr�r�(�ۉB�,�@&ʚ="3!��"D���c��\�/_\��SF�}B!�$B=~^����E�5Z&P�W���r:!�d�=�B;�(W$DGv��Rʊ9*W!�$��61U��,*(I��KR�!�d7I�\���@P�s�0 �^�!��>JQ�1�l�k89X%�9 �!�ĹcW�"UIN�=���"���8r8!�d�i*\an�#=7�!ǂ�	(!�D�O�j�U	O�q�ν3����|�!�� �1臋B�H��	-�@�E"O��(��Os,\��!P�]�"O�飄�Z���T�6�B?l#VѢ3"O��!���4h �Ö���o�yJ�"O^8{�	�Y�t�Y��P\����"O�@KN9 z� �7I�<&-\峀"O¬�GdG<_����N &�l�"O\H��*H>��孜g����"O���agY$Ed�a��L����`"O�+��V[���!�X.��k�"O���q	N�U�Ɲ�5	ކ]� D��"O�<�ł'8�LأEX����""O��B�D�^�F��e\
I"Y:W"OnY�bM��S䮴�DS2>ܑ�"Oލ	�a^2io���5vy�v"O`��B$TWl(J�P�i	��x5"O ��b����[e��4�t��@"O�`)W���,��.�#9�-��"O��T�S���z�,6���s"O��0���{�~m�P�M�P�x���"O�q��Q}-��Ҡ��W�D%YW"OX)j�Kv ���D�����"O�m�+.	����`Ǯw��uke"O�홲�� ���� M�n^ͻW"O]p&�ٔP2�$*B��0p ��"O�ř�!�4)�@�Κm_����"O��bދNצu�v��b/�e��"Ot�@�#�	`l��OY8;��\!T"O�,��)ӺD��raGR�����"O��е"�$L~(�A�_�^�����"O\IH�G�L?��*"*�E�@�a"O体��3c�e�%F��'|��A�"O�{U����E���� +1"O�i��	L���҂�.F� ��V"O�|pe������*QD�l�"O:�R�.�
�1��%
���'ʀ����`}�EW�_���	�'�0٘C�Fb�1F�M�l\��'w� @BbY�y�|�s���#	M�',��F�� rfaa�
4 �潩	�'D�P C�,|0��˖�͑%�\C�'n��g��1qeDxL���Բ�'/�9�_�s"��zf���� ��'����Ad�����Ǟ//{N��'$fI���Z�f��A"��V7QX��h	�'���!�ǐ��ܱr�邐G"4�P	�'��A@&j�1A;���+;3�	�'�6��d���"���
�8%��'���R3i��io�m��� ��5{�'aN��u �M��6N�
�jdP�'M�x�D����Y�l�x`�h�'¤���7���btD<uB�$��'�ڀB���
sn��D�O!��b�'�ؘAv��'����m��I���3�'� yaC���0F ���ʸI��'�Byk�H�2c#|1��`�&
Az�	�'8��`�� �|S�t"!ֽ	��'ZLz��(WF5��ѴxR�k�'�IR�0C�q��	��r�
�'N�i��^�jWp�₧�0u%��Q
�'�(��� O�v��Ūl��	��'�1���$H&|�6�N�l���x�'�.�见Ȩ98�����a���'�d��ᎾK�H�(%L��W������� jP�S��>Iq�K�	�	���D"O\`�'8�M��� �z��"OpX�i(F];g���-�"9"O�M�D�(���3��gc���"O�	P�@N[]#V��7
\�"O~0(Ê��	��;�f
;o@a�"Op5�ᭉ�l��}	��,Vݲe�B"O�mI��N0l�8ebT�"!�%Z�"OH\���I�>�`y@FD���T"O(ظe��&t���h�j���q"O���FG� ���"0j��`@)�"O0�1��f8x�1���O���"O]Y��š��,	�8Ͼ���"O�y�m�#<9�u�A�8}�Z�9�"O&$!�*��\d�	P��"w �Dp�"O�4��_�6z����²*����"O�tC�@W�0F������0k�"O$�Za#��bu͹�홛_7F���"O� �w�P~~I���H&$��G"O�j�kG4n=��#��%!^q� "OH�V�,X��tH�˘}�t��"O�Sq,�>�P�)�'K=,�;�'���"V�{��f��h�` "OD- aƜ�9��1�E^0u�����"O���)kt������Ma�"O���G��.B�Y�3>�*HS"O:��$�Wf�B�:v'
-""O�`��Ӣ~ȅ�`'�	6�JT	f"O
�*U@+SD<zG�Z�p@a�"O���cӎ0kjD &�IiP&%P�"OP� U��&mΉƤV�N�$u�"O�pi��ʚI��Q�D[�B� w"O0uPƦN�v� ���⊺�(m�q"O8p!L5�|A�n��r�����"OZ����Øxo���p�;i���"O�LzBdƓ!:Pg]=YȰ`�"ON��r� ��x�&R2 ʐ"O����H%2=�XX�eJ�b � s"O�=�w�Ъ'�B|9&�EkF&�(�"OL遆��r��ucA��Zq;"On�	 !΁[m�6L�Lv6�'�ɤ�� Z`je�R�7s�=1�'�H�`eĈ	!#�@X�&�?]0��)�'�6$j$���e.�����9Q�@J�'c�q2g ��Q�$�{BPw�B�
�'�Dӱ��x,xQrM΢h5��'F2`R���wb iz�)pi"��'6Q��M�:A��*�-�����
�'4T!K0!>%��s�D!m�bd��'I�eS0�7t�.��%�Da��P��'i����A�[�:P!u�U�$�A��'�Fd������闗o�$}��'4]1��G�}9�Xc�A�$R��Ы�'Y��'"Ssz�K�.ѮDyBU��
f~ճ��M�~�H H���c��ͅȓ?�\��ޘ)�5��T9npp���_�T)��Fk���	�&�\@��8H�����MuN���S�}����p�氓a�_5�r�O�(T���E�v��V#45p����܅=�����n���X���f�G*h�u��D֨��񈋥��QićK\h���ȓY>�ЈA�ŜR���qF�>2�4��ȓo7�����,3��5�1���[�Z���S�? B0pn�>)p���ǀX`@��"O�Tʶ�!m����ҍnf��(�"O���$6sRH� F\`n�RT"Olp�	4��E��bJ\���"O6�a�%F�iS�Hy��حD[�ܙP"Op��"ܟPR@ ��f��jzR��"OƷp+
�8@x�Ӭ\A��@"OHe��F��!��iQ ]4w#����"O�$Kh��Yi$P��n���%�&"O���th �(�$�9�,�6`480�"O�ْ�/Ǝ]Y�-3'��N"O����^.I�R��
Ӥ~�$;�"O$80�g�5xbQ��1��m�v"O��B�   ��   �  i    �  �+  n6  A  �K  U  !^  �i  r  {x  �~  m�  ��  �  7�  y�  ��   �  F�  ��  ̽  �  S�  ��  ��  ~�  ��  >�  ��  8 ! C $ �+ 2 b8 >  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��gëF�ڙ��n��R�p����?�  ��[Q�q�oY1]N�$�u �P�<�0�	���)���eL����N�<��*�%[�J�z�D�(lf�䀅t�<i�*I3ъa�n�!q���H��@p�<�/ӷ,X�C�ni����\n�<aS)Y%֌[�eʱ�Xp�Lj�<	�gA m�&���nݤ,Y�%`�Rd}�'�D���B���A�փ+˪Z���I�W�\4�u/��z,���bC�Ƀ�j]*b.�y�8Fh���B�	*���2�W�X���)dc#��B�	BY�pRVz�D`���Y)���>9�c"�'}�2H1!!Y�~O\@�R�4�&���w������
%`d��I�2=�<��'א#=E���S:&`��#J&�ja�K:X-�ȓlX��0��CC�}�B6YXl��ȓVp�� jЅ (�A2nF�W����L��A+Y����y�*�!v$���� �maѨ[�.8 �mIa�(<�ȓ/L��8s�A-~(X��R3�愄�����	�8�Z K&�ߛNBa��"����wi�=[;�8[�]����S�? � �fZ(�D PA+ֽP���"O�H[&Ҥ_��I%ˑ�Y�"�;�"OfPYDaB-6l�my��τ{���""OЌ)�������r�(W��9�"O�|����*^|��/�iq�B"O�E@�B�*;z����I@�]Rg]�TG{��)Ș����P�؆���J�>�!�$4,��(�����l�����s�!�d��	r@)�,ʓ>����$�62!�d11�Nd[R����H����!�޵2��9r��A�Zvh��)�"[[!�$S� ��qHӽ}P�����C�dv!�DZK�2�a�-
�p�e򑏒�9s!�Ď�*�~���fW��`�44^!�$�T@n�%��5Nl�D�Ɓ5P!�D�!F�m!�*W�M5`	� +�V`��Y����G�]9y��s�D�>N%J��6�O�T��s�κ6�@qa�U'	�ܵ�ȓ(ߤi���GB�	%kס2���Gz2�~�gjg'� H	y�Lh
'Xy�<�-�" m��5bE�g-V��0j�r�<yB��$��h3W���]<���mTl�<	F�I<y�$��aD�	X�i%���<�����"d=97��
{V�)v�Ɩh��B�ɹ+<|��FEį,xX(�+D�_.Ԣ<��T>Qc�kЈep��2҅��7L (zf�)D�(�5�٭oJ�����2�&�BW�-D���e�P�4@mRg)��-{�p��(+D�,8fN�7c�X��eZ#�X|@Тm�p �]5f�۠�?�Q��gÈ|�qE}r�S 
�Hٷ/Ѷh�b��o�u$�B�I�b��(bD�1
�M�P(ܖ
��C�	�"r�U�@Y�p�F�;5!6r�C�	�`�Z�ŭ�6z=$����|��B�ɟv^�9��	�G/!b�핳f�B䉦o�Ձ�i�l �\�w�1J��B�I�C銹1�� U��gH�Fi�B�I-G�L�Ӏ�
g:h�r@�P-<k�B�3J�C''ȳg� ��g:+N`B�	�l/��3`��q@�Uy��\�6B�I�����A?Y��@�[�v�LC�I�D�08��,Zz ai�jx~
C�	G���d�ѿYڽ���	�B�	�q ��A�/\�{��aX�Y���C�ɶ9Ll�ba���=�h���I\�?�B��z0pbS$��V���.[�L B䉠|T؁3d5���jX�4)�B�y�� ��ꄘ+ܘ����r�~B�	�)�RX�"��
�H];��xZ��=!	çyS8���FP�Z���n��'��=�ȓ�l]
⬛5~͆��Q�4����ȓN��ģ���M�ne8�c̑P"���S$p��Ъ>+�m㣏z3�t"�'3 �D˦\P�i%�Ca���C�'I���%> Lt���*��LK�'����p�ծS�*z�ϵ��}��}R�)��Ӳ%P�E�g ͆A�� x�B͓	�!��4� �2���_��8�W!��a{��9�IK�@��d@@3���pЩӼ ;FC�Ʌs�rlk�	�nDS���
��?�S�T�8�DIp,=ی�`�gL=�yB��?I�L���J5rψ�qa�ʍ�y�jZ(���$�!:��7����y��T�c��i�Ύ�f�*��7��y
� �-)���}��Ɂ:"�0�p�'�1Oʬ����KvbX�i��m�j�#�"O��3�x��T�K��<%)b��[o�����-���)� X~H�6�ڡ"
B䉻(�N�
dŔ�7�0[���6�8C䉜^~�L�A�.NV�lsŬY�t�*C�ɇ^��GƇ Q,��Q���Y�C�	�S��� ��3�x������h��B�I+N��<񵭝�[�B��R#�%.�B�I�j0���@�	"*�U����C�I;`+x�w�S�W����5-�1לC��&+;�x�S�/̜��!�/bNN�	S��h�]@��S�'��&Y<%K�&���yr	�0���@ͅX����&�ē�p>g�UXe[6�K�!�T�h �W�<	�H�g*�\RUDҥ6r:*Ml�<�'�á=�	�@kTP���(ͧ{`��XG��w�� +���/b�(+E	Ӆ`��4�˓�(O�,[&(�Q>����R7 �����"Oj��R,�!���fCWh��D����l��OR�X��hq�fF8?��H����;1�А�O�y��	+yC.0$ �\Nڡ��
�0����O���>�O�L�l�¦��?����'T��!x�!R5ז�
B �]؟��I���)��n����ѬX���N<i�4��$1�0*�؈��^�N,�8��U�3DT,��I]�'��DFK�r����AC� �Xsݴ٘'c�)�3}"oQ�s�b�C��_�!�c�6Аx2����t-J'���Z��P�O}��Ҧ���I9}�c�l��B㎁X�t0�j4D�|�a)��b���!�v� ��2D����㓾��`��E�
ت�g�:��hO�1���U���s4RX��� o1hC�	 ƠLRШ��f
����u3PC�	�i���	�Q�As�X3d���LL~C��-Z���*e.�t��`s@nE�2MBC����c�m�8'�����K��w��B�I�7J���FLP�H����u#C��bB��^���(��O�K$r���՝c�0B�I�$J���T�sET�&h�!FS�B�	� d�<��m� p�D�(wVfC��;. %��^�_�`�s�_�3�dC����|��7
��1V� t�C�7l\j\��	9	�PhS-]��BC�I�i��A�b�W�2K�+ ��L�C�	�-��(Q��I%z%�whD��C��4C�����l��@#jq�aGA��B�(%Al���7�vرE�_��<C��]r����ݦ�����Q�E�ȓgm8�
��D�tSh���N�n}��B��);�MD���yE/�����XL��r��'*Hn������IKRЄȓ���g��F�$a�K�)oر��m�n��E��3`Ml���Hj%$9�"Od@ѣ���JZi+e�[�f�su"OSŁ��B��Cbf��Q�q@�"Od��
P%���d�T4����"O�bRe�3*4y0�A�3�Dx�"O\s�� I!NaA@�,-:@�"O@p����=Gu�\Kϐ�b�rT�"O�i���E7 ����rN̖y�(I2�"O��&��ʈ�w�djx1��"O�ix�#� w�(�ـ��5x����"Od,;@�O
WI����&t�l�r"Of,��NM�:��<���.�\e�S"O� ��ž*�Δ��'�ppQ�"Oj #��`(����l�k�:%Z�"O�Y�@�@��x��/ �zēB"O�1�R`�����G$S�*)XF"O|1a��>7�����B҂J{$aB�'*��'B�'T��'�b�'q��'��x1hD$�ZP�@G�}"�t�u�'���'y"����'��'T2�'�pdk�H�j��L�S��/'O8DJ��'���'|b���4�'�r�'��'����q("��x�@�Mq2����'�r�'��'���'���'��'�@�+��A�wC
��R��5^� (��'�"�'�"�'���'x�'L"�'�:��2k��~*���o�S/l�2�'���'���'��'72�'e��'� �C��!Rd%�)�4x��H��'�'���'zB�'*��'rr�'��b3��;���3���i�h �R�'�b�'(R�'b��'-R�'���'��Dj�F��(��q�6�ǁZ�5Yb�'Z��'���'��'���'S�iL&	,��ࢀ�!ɎI���E!>[��'3"�'���'��'��'Q2��O� !��Ls$�����4�'�r�'���'u��':b�'��
+M�-�gѾ
ۀu���� "�'b�'�r�'W��'��'
��$<���V�. �D,FT�2�'���'�b�'Fr�'�6��O��$Я>w�`r�ä<��\(��ߨv�h��'�bQ�b>�FZ��*�
�H�:sIłl3h������t��O�(nZҟh&��s�hA�4�FTS��8K���~�����i�r��Nț:O���2?<aa��.�ɯQOV���M4m����yюb����My���c�L����T4aȐQp%k�&	�4K���<����}��G�p��f��/{�Z<SP�E;K0
�m>�M�'��)�S�E��<n��<����	B�vD��N��e�	C�H�<q5h�7F��8jF웰�hO�)�O�AY�(��O�ڌ��p��)�9O ʓ��y��e���'���Qv,A�
u�Q��K׎Id$���M}r a�j�oZ�<��O\�PǛ�[�	��U�1R}�������M:) 0�$.�S?#�(�;8/���,'�ڍk���/�t��bLB�6I�IZyr������"G�v4a4��Y@4 w��Z���ڦ1���+?�P�i	�O���X����4]֑!n���dЦ��4�?��$��M��O���n��R�	�-�w��Б�gt���k� 8�ГO���|����?����?���z�:P�0n��*��@[Ə)u�^k.O��o�0*D��I�l�	�?���y2��8��q�d���L�{@I�Y�\�ٴ�0O$�����O�D{Î4��0��k5�.9%��*�Z�(`�<)1�F"�x�B�
��0Cc�H)%-�tIbc�"f]���ː�7��.�*L:$��h����T�����G��2h��m4�-hۑ����H�tl�'�����Z?���[�d�{g���<� ��{!����y:bm�A_(�MR��y��� kك
ب �@�#[��a:�)�
8�N�	�
Ts����E�� �l֙>�x��C'�!�p0�O���#��������$�X@�$Έ�6p�S��*N���H
s�zx���4��\l��s�LI N�3A\���dN�k��X�O��D�O��d�<i���?q��|��N"ro����C�<�$���L�&����O���O4�`�M���i��"r�h���a)Y��`q��Kx�j޴�?1����D�O���\�w1��Mt��S>PiZ���B:����Ǧ]�I�ؕ'�x�Sw�1���ON��ƸX��Z�Y��8h��%�����i@�	˟,�ɝFc�c>%�I�?7-
-�h� �ɨ,�.逌��S㛶Q��(�oI��M�4^?u���?eA�O�t��(B�j�f���'�(�NL��iTB�'1$lITR���&���$G^	Z@�_"i���y��Q��m��Ɵ����?uyM<�']��(P��h����ѐO�F��¼i��)[]�x�	ן��3�ş�E%\$\�b2�:%#P���l#�M����?a�)�H �x�Ob�'�p��A���/�M��&ܕ9fm�>���?	n̓�?����?)Cf��{�0��SU}\��S�ÉZ�f�'\���#ů>a)Oz�$�<i��Wk 8c�!�V��`�F�k�U}�#� �yR�'���'	B�'$�ɵFg>���ȱ�)���P�a�&ԙ@%��D�<�����d�O ���OM
$d�6��9���U��n͂mN�$�<���?��?q���J���i����ֆܽ�$����1Xz����`�6���O���O����<q�S�N���[�L%i��q����4X�@`�L���	�q��0��Ɵ��Iٟts�I#�M���?iS�ęJ��	��}ʪ�k�ݫ��F�'��'�I��X����~y��O&�3�̕�^��IrwK�LUp;��i�r�'���'
�ѹ�$y�x���O ����l)�@ʝ7_y�$q@*��C��Hy!Pᦽ��oy��'��A��O�2[��s���(!mȂW��,�"!7J��׼i$��'����*iӎ���OL�$������O�Is�,�86�$m�F=Y4f�8���g}2�'����!�'$�Z��L��R-(�5�Ň����#�^��֫�#`f�6-�O*���O��� �d�Ox���`i#!B.~�T��B�n�^�<L�	^�i>M'?a�I mS]�PJ\�\E^�����4O
l���4�?I��rڴ3���P��i��'-b�'ZZw�Lqi�H��Tr�|Zj܂`��bݴ�?�04�p0r,��<�O��D�'�ҥ=� � 2v�Q��ҝ��(k
��Ǻi�rJ�#uj�7��O���O��D�p���O��	��R�*�`4�$�O�`
,\��_�ȺQ-?����?	��?��?�5g�U<��hv䁱<z�x���
D��i���'qR�'C~꧹��OX�!4��,'�~� c�?wL��'!�a���OX��n���OlʧF5ʀ7�i�fՉ����,���CS�p�x��gi�>���O��$�O���<���/f���ˢ�08r�WL�^2���"T��'{ĝ)#�'"��'�b� 4G7��OF��6=v���"��H6�qC���Ky�Dl������Ɵ�'���.���X���0&>v�(5�Q�X0�j��X&����ȟP��ȟ�	�o��Mc��?Q��B�����t���qA�Q��'nV���'�����C�No>-�	xy��M���B%P�J����z�T��NզU�	��k$�[4�M����?a��J���?YWi'N���6�P�k�dh�"�U���	���!�	�ԟ���矜`�Gv>M��Ќ�F��B�xqh�KP.J���%�i���z �y�F���Oj�$�T�I�O����O�	���:����m��	\� ��M릍�T���_y�O��OVl�%
�B�r3J9��J��Q�e47��O6�D�O��aL]�5�I��L�Iڟ��i�a���T>k�f�iV蛉?�&��t�|�T�ĺ<��"A�<�O���':�ꔩ����LK�n(p��?m�7��O��Sr�ͦE�	某��ğP�����	�M�z�K���NWNL���YH��i�$����O8�D�|���"�:pJш�$�z�TL�<�R��tKO�h��v�'l�'�̱~�,O���'9������KIT2Vh���2���:O���?9���?Y���?�u
�8��֍F�jrR�KS-�
�X<H��C"�6��O����O��$�O���?���V�|ғjqO�)��hӛ wN]r�/�4��'f�'3��'���?1��6��O �$��~ [�&��J���?�$t	r�i^��'{X�|�	�h���� �	�H =pw�Í�B�@,��d.��t�Mş8�	˟L���v�Ĝk�4�?!���?����j�+�i�2X�8��5V�Z�°���i��T���I��<�Sӟ薧��4&x2�`KޖW����B�W��J9o���ɡ?)��4�?����?��'���3~�e��̳W�r혁f	!V<z1\���	� ��'V�i>�ӺK��ҁ{�Nx��oG+4x�P.���Q���M��?����b�'�?!��?qu��o�����20�6���>2S��R�-�b�|�O��O]R,݈y帍��αHrp�` �I!�6��O��D�Oj�y�)Ҧ}�	����	��$�i�ѨA�R�"w᝴=a�I 6rF�v�'9�	�F��)��?���"� ���,:�(1�t���T����i��޼`h6��Ol�D�OB�A���O��'Η�_b����;O�!3�i:� U>�y��'�b�O�r�'��$����憔�X��-	E<m�y�H���M���?����?��]?�'>��W,)��XVF�:��1� � ��XA�'b��'(r�'�2�'��ùd�6��4}��+_�u��d��k�&�^ym���IʟL��러�'("�������.�,���+d°���2��6��OP��O����O����e�TloZ����	?K��U�M)d4bE�5��Vx�)@�4�?���?�)O��D?;���O����)p�-�xM���c�6�O���O��d��x:2n�ޟ`�	ڟ\�S�@�$�سb�9lz�RUa�+;s@`
�4�?�(O\��ֵ+V�i�OT��|n�/A��B%84�*��G�$Ң6��OR��߽e���l���I�$�S�?-�	�f��=�Fj�=m��+D�Ȟ!1"�Ob��ׄTc����O���|�K?	
"l��z�xp�)\�@���jS�s����������	����?�#H<!��C�& yp�_V괥cL�#ZI��i P���'�剾�H���dǉN�XcE��8��Ux�� ���mZğ�I��rF'�ē�?��~��:D��]a�E�}�֔r�(<�MkO>�ł�x�O��'���.Q4h1q(��5�SĘT�(7��O�rA�v�	ԟ���~�i�]ò�������u�إ)yJ�����>	gh����'���'�W�<9�3V*!��91k6 ��6:�#K<9���?�O>1��?i�-ͅH�(�# ��aV�-2�
�?-��͓��D�O��d�O����͓�0�zp����6W>8
�iJ��Ǚx�'��Iԟ��IПl�bOr�LY��ەs�X]귀o0(����	���d�O�$�O*�9��dƝ��\*ji;v�غHH�(#� ��V6�O��O�$�O���,)�I�z�h82kQ��,��!�J�:6M�O��$�<���>7�Ob�O�h�S��(u�Tb�G�u�Rh���6��O*��Z L��6�T?a;���,6*^U��v�,	���S����܃�MkZ?��	�?�c�O�౮�0|�F����M*wW�;�i=��'S:a���'��'wq���+�䑍�~X��^�FQB\Kֹiת����}�T���O��d���'� ���&|i��a���HD���&��M#�4W\Ba8����S�O�� ̠=������sâ�ȖA^�Iӌ6��O���O�3�iEQ����N?9�̆�~��co��#!@p��eJΦ�%�H떎g��'�?���?	��ѧ�����ѨUH�z`O�2$8�F�'��sU�*���O���<�����h0A���j`aA��5L����Q��	��O˟h�'
r�'7�Y�d2�W�Xp%{�؇-*�0�.L��j��M<���?�K>����?�s�ڽO|H�:��6��!�˗��u�L>����?Y���$U�l/���g�? � ���Y
w���Ӏ�s���Y����ޟ�'����ޟ\���������9(�W!��f�itFȚ���O����O�ʓi�䐀ǒ��@Ζ7tN�1q�]+#����	L�H:�6��O��Ov���O�d�G��O:�'FV��g	�y��@딍B5R�H�2�
C�ny)Dm��q���R���//��$�ԑI�z<F��#|�� �w� ���-�~�Z���UR|pz	�'"LÑ��|Y�Ae		.J<��5^���'%�S���B�̆5((!D[�sF��QT�M'$���� �?C�aB�F�5&s�=:��W�@���;N��� վiԢK��!D; �34@�/]����>���t�1Z'h0�ᑈ>h4���D4�$�X@j�]YpEܓC����0��D��j��'"�'���h݉�c�RG��bfF��V�� �sm���u)����?�@�	���|&��b�HĿ�r����Rp0�ࣧ�55��h����?h� �aQ�	��>�����H�c`ƓS���C_
��r��7OO���/?�S�@��S�'AT�@�%\�k���Oy<��'֨۶m�?U,ͫ%:}�Ⱥ�O��Ez�OP_�HG��3h�(qr%�q�M�Ч�:d\�ؑ��ҟ��	����2�u�'!B<�͐�I��;а�ʇ�ߥ1�<�y6��E�!�[�%>H`0�:�|Y8bn8a�0�O0X`�H�8"�鈶 I4J���%?�rf:�O ��Ȓ�5٬u�Ǉ*q���q�"O��[���Gў<*t�?�:	����a�_2
�`f�i���'�Hl��H�"DY��(J��]#��'���ڇ(�B�'��i��2�"�|(O�9/^Ix���&JTQ4\��p<A�g{�<1D���S�Im��h�-�|��܅�	/N�.���v��_NJ���b1W��U����1_2�B�I�Sr������p�6,�b��	��B���M�� �0܆m�"��Ibx�$P|�d��84�i�r�'���c	���I3A��Q�OA�RȈ�I ��8�����ş�w
� �TZ*я-J�i�S�$^>��G�?O#��pB/ Y�#l1}�`S@�l�h�;w�𙒔��O�$i96 ��o�>�@�JP�p���'�.}8���ɧ�O��В�aS6�|�[��DgЊ�X�'�.,[֥�=�xZ�/B&em܍��Q�He��7.�0�"E$���g��
���Ot���O�H�d�M�w�����O����O��=IR.|��N�aRP��`�<�A�Uϼ\���O~�Ѵ�1��'ofS��^)��Z��n�@1a�
�fV4��!��O�]��Ƹ��"��xt/�/�HC��W(	�>]J��|�aW(�?�}&���q�ʳ(�ahceV� &58��2D�\2�"L�4��|8$-V�b�ƽ�#?��i>�%��z�b�.VSZ�ڕ�N�b2��	eG���IȦ�����ӟ$����u��'��2���Ԫ�%f����b�>�(=z�@�bɊ�"��4y_�p�+��1g8�F~" :	�b�r�jU�`<>��e�'A�n�!���-]�xYc�^Jb���o;��s6�Yiܓ^Y��i�ƌ�hN��$nT���T۟��2p���Q�C:|P=�u �W0B�ȓ{������� P�@��߱A숰�<��i��'��}X3.p��$�O*��F`+>��9����i�A@��O��Ċ�.��O��Ӻ	�d���D7_���!���Xh$4��I�m�x A ��\�`4�dϨ��O�ъ�ȡ7x@Ast��[����&��<�����T�@���CQIH)J�	àH�?'E����{Ri���?��xZ�x��&��U�&�GΙ0L�X��BEX(��.�Rp�E9҄��XՄ��=��&�,�bUK��J�����EBj#�'���Q�db�@���O`�'y.pe{��t���!��:Ot�i!p@�7bܗ����ɣ�~6D�e�4���:�A�?��O���k�
�	cpyH�[E+�e�O��3��٬����E(N�r��4a�25(8�*��˭U����>�'%<D�M�"� &P�Ky�4�Ɇ�M���i�R�i^..��S��8d� ��v!	18 1O:�$�<Y�����y�����o�pMk2���d�axs�$mo�<HhC5lB'�Hi� �\�(}���۴�?����?	4&�0H��R���?����?a�;2�pd�UM,�&|����RI��*�y�"���<S����l��9M2�uܓB Љ��	R'VHI���*�y���D�1M>���ϟ�>�OhL��nЛ��h�q�c�~@"�"O썩��ġu�h�镍&'��C���L*��ᓄR��z�҄E�� �A�%��9D`��:I�������ݟ�r[w��'��	ؚ�)�I�K�~���h0?&-��^�B��y�l�K���@�k�'���ǫ��5�8`[�C�8"�X�XV�D8u�b����ɷ[�(
ANەRvJ ��+�%�x��=�U˒#QRm��cC)	��r�%f?I��<��?BDX�:��5ۡ��'I�$e���GU�<� ��𗏍P���`T)A�u)Ԝ�%�Ğ榭%�L	4����M���?YbKX�M�^`�s��`��*�Ш�?Y��`sLxY���?)�O��(5��u� ��S��:$Ÿ+-r}�D���k�0�gF%O ��G$M��:1� �N����ʄ"�*�K I
t��.S	�@�.�	���Ɂ�ēH��B4����,�д�ȓvP���rB�����MYT���	����V�9�d̲��ұ$Ұ����'X<X��}Ӕ���Ov�'��(�n��%	�~�-�cLM]���X���?ign9��`F�ɑ7n�X�:B����n�T�P#�X���,l�B��-K=��%`��Q&�zQ�ă�*!i�����B=���E���{S��J��H�.��6-<DA���I�Da�Jo��mZ矴��卝K.���#굸R��^��?)ϓ&]28	vG�@�P�k��٢J9���HO~��5�>o��S�mH���L�$�즉�I� ��<2*�*f���h��ȟ��I��ݳ��L�|qW'�=��l+���$]�`r��CJi����r��>�S��	�s��Q;�A	;L?��慃	�2�x�hQ�qX0cw��uE"�(�hC�(�O�b�b�����OtN\���ւ4n��e�I;]��'3f�������BKd &��%
�v܃�/V� ͚1��5x��b�Xiw'ʠN��)R��#?)��i>	&��C��4�=pЭ�&N�� L��{��Pꐀ�ßT�IٟL�	��uW�'�R0�`����F7 �y�Ə¸E�L�S���&h}j�!�J��<�((<O�pcBU&;lC2kr����!� ���M�q�H�)���Kx�����n��Yc�F/{�5�U	W��t�$#�O�,�W�+m|��� 1!g@��0"O<��A�]�d���5$T"@r��DʦA$��cP����M���?r�?���� �0|����I�5�?a�P�n4���?!�O�t%!f�B�K�@��Gϖ=&lA �Ъ�d��w�1(��9
4�Ԩ4��#?�ץæc2T�I5
��iȊ%Ѵ�ٲ�0`���E s���3�m� SB�C(�
$���;4�"�ɓ}]����Q�	U�^�"Tŗ.\��¬R,~fB�	�-h�90�����2��&ZB���M+�F�kH��td �['�]�����z�,lh�i.R�'��S�}������)+.}�戝�C����N�E�� ����8�쐥,�T|0��L�Gn݂�йt��I�|2���v��Uz"�����H����K���4Cm
��C�%F�drPڪJo�$[���i�Q�Og�<:��L�,�������6t^�cI�(`���O��&��?��#"�x�p���&y���vG#D�d�Ѡßx\F�؅۰8@�� ..O 9Dz�� 1�]j���`V f$^5qͲ6m�Ov���OP1�"��Lt���Ol��O�.M�E��b8b����mل[���ӄS/f*U,�*X�^M1�����1;�|�zݙtj�Qel
;QL��pH�0U� 	@��O���6�ά՚�O�R�@$j������ɳ{�HKd���#���h% M�Ř'���H�S�g�	�d��H8�MB�o
BE�a,	qrC�ɪV|��3�Z�V�1�ĖNp �ZK���X�	�L��tB2哈dx8�ǰP�0�X�C��$��	ԟ��Iȟ$JZw(��'��	�8�3��,)x�M0@΀�A�x��RMQ,AZ���4|O�ys'�!dV�t���͜�bU0ah=*&�{W��v�:\�P)��(�RAF~���;{�ڕ�	���LtP���k�ɒ�6�a2"Z�7\� m���	�y�H%F�[PCِ,�j�9b�ʘ'{�6�*��R<7�,�O��`�A����v �; ��%�'_D8��'[��ir�'}�5�BPJEc�6�p��#��rX�z�$8|��|R��BU�p�L-5$F~��"x�(r��_�S� ��*��Uc��/
Y�T�� E 2&U1�U��2E����c�'�4E���Yg��B�>����=�
�q�R�P@{��V̓�?�
ϓ
wT�`B�7��Q�dT�e����u���/0�$�a�Z�R�t��t�\�#��U��:��Ҭ�M���?)�6�§$�O�h�$�V�2u�I�,�Uڰ��OR�$�6I��r�]8?��!1"՝f�����O��S�:�(���
�
9b�a+3.�'C�S��Ɂ"�ܒ3a�$��Rf�=Gx�8�R∽7�S&s2Q9$D/cv�֣@�i�]��$��2��S��+�\�1��=*�0E�	e�,�ȓ.�i�������)�M�1�T̈́��HO���A�.�LT²E�3��-)4*����	Οx��u�E�����������i�ͻ'烙jH�2��*SP0��N�&O��v���4೅*<���|���>i����}�6���[j�9UK* z���n(���(&�ޗ[��k��J��S�C/���8��
�9�<��%�-X.8�TM5�I,Z.0���|2�A.x���)e�V�Y6H�@Eٞ�y������ĭ^>"hX`3��2��d�B�����|
� ���%H��+I��i1�;D������tI�F��O��D�O��Ă����?��Oz��;t���682<�lK�� B��Q��	�W1R�ca)_�wj�TF~b�ǛM��D�̟+7���3a#J�X����ˣjC��P"��v&���������_pD%�d��΄�2�(�'�+_-`-�2�*M�l�D��=i�4�?�,OB��-��/ΐ Rg��4�6�P��]8>B�	"\�D�@��^��(��ۑK�b���4�?�/Od�r�'���1��矐��Q�T1B7C�	W��Ze�^ԟ4��N��������'w^�h���;wmSNR�-J�a� !Սs�����kػUL��!��@:u����7�6N�-��� h�0�j�;~ �cV&�� ��"��T���򀁜�T�Pj�J�T�I�V��d�T�I,J��yi���in ԰�
�	WB䉌�Q�5`B/&![&%��_�""<q��4��Yoڗ*�t��JȐ��S��?�b�D�����M���?�(��)�A��O lq��_*8�=!@�Ɂ _�p@�O:��5�Tsa\��M�!`G5fG�
1֟˧M]��Kr�� #*]Z&ږK�@�O����J�	�X��"/FJ(��2�C	�|�nAC1.�����J�+q~�
��^ >���cB���I����O�l'��?Q�QEO���ڄi ����w�"D��9ƭ�PJ�3"D�����) O�}EzC��-���g��qk��c�R�Q%�6-�O����O��R���AVp���O��O�
����0�*I����L�.Q�-.��,{�����V�\( ��/�?���fNO�P�qOZ�R��'%��;����g� ��7@0@�|H��>�� 0D��L>��h��M&�
'lRbhT� �DX�<Y7
Q�J��ʙ������Qj~�(*��|�H>����v%��S-��*EjH&fiY4@��?���?���w���O��Ds>�f�XBM4�*��&B��(C�V�h�Du	�CW�u�#4���������D��),|���?��E+EC�����i��_���1��kMt��êB�OH���ߙGOqOr}i��C"M6eQGgԫb�N�rdE�F�r@3�O����{� ��uˎ�t���z�"O����+�-<zf�r��ɳ{�E C�D̦'��J���Mk��?��闈A�޸�F�Z�[u��O��?��6��p���?y�O� @ /iP���@�P�~]�v��Jކd��T|�h��ʴRB�	w��M�'��l1�4J�����e%�q�Kݕq�y�r�:mA�7�ٲ
����l�' ����l�'a�|8C��"��Ĩ�_�:��Y�'�f��&��;P6��4'Kh0��'J�7��[LВ���9A[�� �#dH8�Oɨ�eG�m��ʟl�Oۚ	)�'R�A�FBH(E
@�Q�)(hNh���'D�aLm�rY�c ��<:����D(ss�L����I �^$�3aޔpǼ�H���1S/��n�q C�P�Μ� 'TW�h����b��4'p��!_��@���K�XYZ���P���'�n����?iL~�L~r�B�� �6�3c��)X��mqC��k̓�?ϓ[�Y3��2mVabaʛS	p,k��4�2�EzR�Ώ5�xh�ᛌFM�es��90��6ʹ<���Н�����?����?��Ӽ;��3r�[J��k�̌C�y�2�hQ bS �ʔC�5hdV��1-�Y̧Z
�m���p����C1~������ٓD΀�MJ��"�&��<H��
�>I���>U)��>K&��1T<�R�B@-/�  A���n$*�l������	J�O��3�$� W�`Un�h$���f���!���=G 	FD�[�d��&,��A�I�HO�i�O���>` �J� N�;@���8��eKA���8���?y���?�ĺ�,��O���uW�]s#�ͪv���ʎ�0��E+���:�~cԈU+:�0�	C��Eq ]� �	�:ވ\YQ叝Jk�x�P�������2k&\�@� 	�a�bɗ8P@\YP�	��Ѣ��Ѽm|\x�\jt8t�ޗ��,>�O^����9�xa!�,�K� iÂ"O����
u�h,@�Z�e�Q+��$�Ϧ&��[4�Y��M{���?��)N�j���kVCI-'����?)��8A��*���?A�O�$����֕��#���d��M��e��Lۑ��R��|�4�6�D���f�?>f�F<j���9V�#xy#B�e��ҰkIZ%"�;����ֺ� a���O$�(�K��	P�kц\�yrF�⧍%D�����X�C�F�1c!�2Y#t�7�!�8(ܴqT.��cX~0(b�N�+zZ�YO>i`�8p[���'�P>!q1gS��$(�H��z� �� p�������	63���H�긙!Bn'I��"�);-�H$�O����i�w�5��HnH��ZL��!�ߑ5�Nܲ4,S!Ok�1"��̧�عP#�?�!�G�{kxh��Oў_[^��!�.}�G���?�7�|���l��9A�ҐnfD �a�9�yb��Y�|e���˛S��s��;�0<��	0pmF)��<}�2��T�A0� A�4�?����?	��Z$>�ȹ
��?Y���?�{�? Xx�S��$B&��
�3�f���%������P�H	�5���΂b�4���>8rqO���F�'_��@4��
=<���L�:�:-�"d9���:���L>� "ϵE6�9�N��k��l�Ga�T�<ad��6+H�8E�۸%������R~�e7�S�O��U���25�	�G��gܰ����3-U�9��'d2�'��t�U��۟�'E�l���I�a�n�Ђ��3�A*�Z�,����i̒��BPFW���O<H�cW� ��0yB���OO�Ł��Uv=ѨF�7C���ğ�O��?�,=:�ԭ��L /������"�����?����o�`�g+D�y5L��m�J�<��D�6��TB�0�fj�́H̓OP�OxE��QԦ��Iܟ8�F��
+H��q�H�0�,��̟P��w��џHͧ+J�x��3�����޿B�|��S6]<��ʱ�вUI�x�Ҹu��a1C�	�{��	RR���V5���\!e[���;�`��I(�M���iZ�Ő1�l��`m�+Ɩe�5D0P�I���?E���H;\��L�15.n��E�[��x�@xӚL��?m��� �EW�N�MX$>ON˓|6�`'�iJ��'}��F��	��]
�@]pZ¡"c��o)�u�������1Vީq����>�ޝr����i�|
dh��2@��ôhR#P�o�_ ��<��8N��]�U.J��c?���n
�hň���{x	���4}ReQ��?��f�O|�O�8%rm�)�e{Q�̷r:>�B�y"�'.�y2Gy�
����9��f�@#`"?��ij6�#��J���M{�В"���2�Ճ9{�m��������Ԣκ�&9���H�I���ݘNqԙ��'"�tx@a�S�t8���<y�e^Tx����ág��t�'-~���S�'�I�����d�2��b��k���kч$�l%������Oq��'�Ȕ�s�
?h (;�L�Z���'B��� c�VMCV`�Or��)�O�PEz��		�n����i��,mq�‚���G����$�O��d�O�����?�������L^�!򮈌$�b��J+ �k
�'�X��6C���";'��%�
+�x���6��uX���U+F�{�h�!���B�W?a��.@v������V��q����yr���8�
L۰O���#�BT��'c�\p�M^�M3��?A�
`Ht�"!ƠcX��A�����?��qfp9b��?ɛO��2����=yHY�&�6K�0Ҁ�]_�hل�I�L�����	"pp칢�N�@P�h:p�$O��1��'� O2+�(Դ*~
�I�]�RS6���"O$��"�G� �1�%R�ICO�yo�1̼��2}�j\"�Lë7=b�d@��.����O�˧ynX��Ш͒'N�:M�*2��X�\��i���?Q4�^�$VPո��X21�tY��T�|��n�cҁ���K$���m8(@	�����ɍl������1Ŋ�K��F�B�~
�#</�Y*��@2�����Ze���d/R-�B�D�t�O8,���^sr����f���O���,G-I^F���.�"L�w�'Ɣ"=��U���<sC������9	� �i�B�'�r"�	�*��a�'�2�'7B%l��Z�nxqbb͇t���
٪2~:�󀗌�?q���� /��|&�ԩ5$X4pJ�5k�$���RŊ��ic�r���(�?y�͔2U���>�O�{�H�("�T�6�BB��{�ɗJ���|'�2Tz5��$t Y�wjǆ�y�r�d��,jtf��i�����W���T�|R�(p��Ӣm�d�����K�=���mМ+�"�'2�'d��������|0!
�*�^�xQkؕ>n1Kң�g���	���  �������7J8�ck�D<�@ ��L9��Q�2�;�Af����	>��?�V�ԌpX8�� �ƣR
ă�+�H�<��札��a�E�{���`ǥA�ea{L��i *5z!�W���q�f��y""��vR�S�cڜa�~`�P�X:�yB�	���AL$W'��; $�5�yr"��;�2xaѢ�+G��됆޵�y��9�T8 @�D$��.��yA$X���f[��8�{%@�$�y��?T����&�^�<��Y�$��y
� `�qN՗0��F!�[����"OH��fO�yd����A!�"O��#mW$g����'2/yZt"Ob��$$L+4�X���N�:|q"O�ڤn�]��@ׄ^>L�Ve��"Oh�%O7qE�y�t�t��5�"O`��[�Jc��At�H �H��"O&��Ӊ׻j���-�<�ui�"O�8ꂅP��:I�)·+��I�"Op���.D��St�"H�<�T"O��P�Pi��':�����"O0����t���V7�v�x�"O�L�A�D� �~�c/�m�H�"O�ZB��=����`������P"O��b�o&Vm�<:�R$r��t��"O��r CU�	r���!LK��Ӆ"O�pG�?p�xa9A�?]�"O�47�Q<X���	-0>��D"O����B_źt�Q�.e5۳"O�������D.l��e�5cT"O�$����m�WaO�����"O��ÑTU�!�?����"O�����0	mr��"��4�l��4"O*�2Qɞ0g[.As'�j����"O8�P��=PJ�Y6G��j�6!@�"O�)�����+�\�iNR�Թ��"O�H#��ɔ��gΩ&|x�s"O�A`�'�%?�%�D=ae�8w"O �Qf�м	�9����D�*��' �Sb��QhR飂��~#|mq�X�Gn|��'�������l�fŹ�G�3Q<����ĕ �e�0#�}�'_�K��2�t�ϑ�y+ʜ��I6O��ֹiL�YU��2|�,Tȹ�ˁ�<`�B�߾��3��|B�o����_ y���	�O���ݞT��I-O�pj�۝,_>13#�ۉ�
�{پ}`bN��S�����S6��xExb@�6,�sb�(}`Z��P��M���ң�Nma�� �P��I2����Ð+�z��5i	�5�Z$�U��9p�x���7���'~�q჋U ^�����BNh`��(�Ok�?ku��caRc�h�b�V D��>����a��Fk��|V�U�(��)��8�A	�)P��I��3�0<��Α.
pN�8SF�OD�@��ʴ1��`k��/�d���k=/%�?���u���a��Ŋ<Ta��BN���	"C��|�wF_0@�L�S� 
�<�' F�:R��!|x@`�B�Or��	�O(�F� \�B+�	)4�y���T�\h0�i�h�1%�VBv!��+�0<)E��6��D+֯F��!��'%h��'1~6ͨ<���ċ�Ylm1�+��S��*lŧ��9�!�''�QȪ�p�4 r��O"�zź�étɈ��$�-@�N�IB�'@�\�2!:	�d,���`}Z!��H��  s�Ô0 h$U��l�.K��'瀤�P�֨GD�{U�"x�,	�J<I�2O�X���4����X�U�� .?qD��	��P*R���Ua��@1$���E�Z�A%"��e�I5(��	�W�t́�C�(��u ��I�9x�{aA�<h��q��`O'�y��'<ʵ�aW�Z�Mig��'w�����L[�'�ў�];H�=Ңß�V<ݻb�C�K�L�ۓ;�lt*�kٵI>�x�-�ykf&c���(�h5X r��Ř�Ƹ'��^w^����țs�J5�E��5���h��"��T�|ñ��/��Op-z 뛌c�d��e�~��u�ˁU$ȻB�f�.�b�ŀ��~"E�:��1Ys!m��|r���
G�d\Fx�I�q�b�@��#.~�Ə�
x�S#�AT���i�����g��ɱi"B0���N�;J�	�.Y�-f��"*�
���'�4�O����%`{z���^}��%	x}��4�?��LHQ�@ɊO~��H@�5&'%Q�]Sq�F�<#��R�Y�-p����^�a���^3
"Y10�,)}t�J��UDh�FEO9g�z���C��?A��V�.\�24�i�t�H��E�|��M^˼c�V�n�Y�K�	���׮J�'m��b�F"FQn�ϓIa�����A˼8e�O Д��T?Z�4q�ȃ16~5�	]	~H��QA'<9Fx��gs�D2ADۓ0ؤ2��Ҝp�{2�[SĴ<�'�-֧u�Dڡo�X�1��ʬeL����VDY¬چq�xѫ@�v�й+�cU����i,�O&���ո8�Ѐؔ��~@�ԑ�mB	��IX�� BTK�ie�DbO?���4,�k,:� ��b "� >�8��� 7��wN�p=�d�-eG���y1 �3m0��c�W(.����%c��1��jy¨�"��k̟Bp;��A'����Oxxi���VI`�Kfǋ{�x�d��=z�����O`�Ib��HS�-$$XA�+L�vP�@q.��M��`
;���Q��D�;.I� ���8�"��&��XJ&-�em����R�E6�T�m��$R��Y�nM[�(�I5oQ���?Q��^�J�"��i�,J� ��g���Cc藴l!�T��Bт$�z�!�t~H��'�`y�en[�A`rtj��En�
a0��'Yf�I�WŸE(���8�db>7��?�xv�0o�3B�FNP	D�[�'�a{�@�)jhy�Zc��X�D�H>����6T�9 ����(�d(��#?qD�O�����E��u��y���ý)��-�(Z���c9�t�v-9 `��;��0�'-��?h����c�Y�]R�$�P�f|���'���'��1���0���4;�1K©>}�i͜ix�C��
������8P��[��׍q�<��O���uߴ=�Z�I�T��(�!��>��P�5���?bА0$"ݫB����GS�Y�')������deZ��%��Bz��2��}S���'w�7�0sCM'��3?a��(n\�ܨ�.O�ht10��C%v�X���IA:������D��g�0x�B���*V���QANE
=��1
O<���,��
V��Iu�-k%�41(�ɗ�H�[��	)Y��-i!�R�*��i�@�'�{��F�p�H�cɤ �����ِ��$�O�`�5��݊i�\�r-������95��Mdk�) ��#m�, �.�QGb�46&� ���~R�Ȕ��L>�P��3{G�,z��Â/(�c��$�(9�s�؂g�<-�����	�7hV�Rċ�{����%�?p���{�n����$ϖoi�i���.�s�1bǍV��ij�X<l�ȔZ�"�O��+�%l�p��GGq�[�4�Q)���@�/O�M���WŦ5z��~�gT��`�O�$Qz�$��7���5Aד`r��0bc�'#�<C�C�;)������Yy�v��O2]�A)���PVk+U"��@�'�5Y�0�U�iJj�$�����'28��e)�<��,��nϔ
6�������w'ݲ<o�M�d+P�:�8��S���yg-X�ns(i ���<�
��J1�?�2��A�����'��zg-X�	xr�ڋ4M��1垈7Vb���SV^�k�m��<�5=��y�BV�tx6x
�3`���%;��>)�[6�R�H��Y7D���p�ʃ�@����ʣl-�tAp0O<�`Á�Zk�=��ڟp�a)O��/g����CB�l�*|����A+ΥDy��L�o箴��KR�l*}�����?���+�R��'�%1��l2��ک� �!ŜO�]l����d`�$N!��+����!� ��Q�Ġ�T4Y��FI-=������	�:�BAHc��l:�짿�P�Ĳy+�,�p��	H5�[�,���ۂL�8�ߓ\(x�BvoL�!w��!�L��o&0%ˁ�I�ĉ1_LaH�'w�5vߟ��s��.rj�� îR��� E�C@1a|��	r�����0��C! �ۦjN�=�^���B�c�<p�'���B�O86��\r@g�J}�'�R��"�gƊ��SC�&��9`Ң�O MX0U,FO�)7��6��w�'C�ѳ-��y��t� U 2f^�Y3��-Eo�``p��Jě�`�,O�榡�gy�-�/���4
�_:-@%�N�"l�"&�#�����"t�¡갵i��)��w�@A��B���-���nh�C�z�@k4F͢	��X⢉F�0<	V�N�T%�Sb�%�*��4`�� ,��PC�<� �àA�SR�O�����(3JxJ%͊#~; � ���;��=q�g�\�G�ĿK��QR��f��1VaX�kBL�ٴ��>e� )k�Y�\f���瞑JCJ�'Xd��߸
A|Z�X,n���DzM�l�lp��`�>�pS$�����6��¤@؂1ܭ2�J$�6�5	Y4(��f ��E��+����	=+��R�M�d��S �5X���o�ʼK�4Y��
cd��)�s�9�c蓥�bi�G�L>6~0耱ɟ{>X�'�=$��a��.X����H�8ta��Q0� ���V'`�G�q}b�/E6: y���%k���'E�& �Fb��1o l�"%��jMQ�gB؞�3JS��yw'�Hq�����ܼh��		)�b1��O �M��X�H�|��M�8�H��.���f��& 	���cըg�R#=ɓb���h1�h�D^����b�S}��� �&1���-m��-��FK%�?��c��M��5O�i��	����?� �ЕÖfE:��(`�R3���n�2XҭJcRY�lT�g���S�s�x)�- �(�W�5}�
]ઇ�2�P� �R ;U���@.�x�I(X������#��EF3Xn�Uℊ%}����&0�|��������W8�����	N&4,�5"?�OLiZcT�2�����A23��: �@�x�&���.E/x%�5�L�'�d�gɄ[~Ф������ݩ[����oL�z��qFz�� KR���Ħm��|�3�E�����l�Iz@b�2 �`��˻N�%�8� Bշ71z��	C��|)��6h��3��0�OR B��6MZ;t���Xo��#!�� D%���<���؈� 'n�*p`$d�o�ȉꅅ-2b�F�@���@�^l���Ǉ�,;ʴ`b䘹c�E��.^�'9d�{?�)O��'����l��%��8���H�&��3u�'9R�rӷ���� ����0�k$�g$���ǛK�
A��c�Hr�O�&��6�$��y1�IE�q�Bj�)ّ7�3�+�y�"�=�Tm�PlHr��-hE����I�G?-!)c�xÖ��3�$Ő��0P��5h��}2'O�<IG@�:hV��[wr�'t`� E���.�� �X49���ߴT H�p�m��$�&�H"T}��&�<ɢ�I`}"���s�T�V�].:����V4��$H�6���
#+�rx��*���D���;C��)Y-�x1(K�B.\�KH>9�(J����9
�N�hM?��w��s���&��T��dxO�=�a|�.ӓP�wOҽP?d�a��7u��" JH1O��&(Z{�'��I���Z�h�D�=�ֽ�T�"F�*#>�Dc�1M�æΚ��C� D�<9��Čl��%� X��r�&����'n�$�YY
�I2Hh06ū�OʀH5f�A��}�C�P�W$�ѳv5OVa���4�yAj+�ʁJ1�'y���c��E~.���a�J�y��'�XuC�>�&��0i(O�رEBO����``.awluP 	�=������D/����"]jj\RÀ?[�E��I�
`�w�v�c�GD�,�he��ؗ	8VH�%F�MµJ��;���g��:�,��_�C>ʔ�W��S�'�ͱ�A=A�Qه��_�J���Ol�a4aV�W�e
(£j�XD�	! H��`Ҍ./<=�,@�Ud�-y�q[�l_�Xd�3�ϼV-�lZ.˞��c��8�F�oZ+e����=��R�BĈX&s���v���h0�<�WMM �d`5��..g�ً�۳?U���D�a��y��R5oZ`v�].Љ'^��nP��2ƍg�g}�n��@���W�<iв�"�U�khy
�2NP�o��L8�Ȑ+
h�I��Ȗ
�N0!0nʤ�M�fM�{零�җ��D�Ayb<��3�wm�����,�T����f	�u�
�'�I#���$v���xu3VȏR�XQ��C�1 �l7M�.F�����'3 +@$�)_�r%�[C���	�'���x"�6ZK��ct�	�J���qU���M�Bc����qF�o�\��Z~J��F��)T@���o*!���=��Y�R�y4�xk�ُ{'!��?WH�H�*"`h�L]�t!��+\��c�-ux)W�Q�3!�$4?0�,aP$UDk�eOq;�!�	�!_�����0`�d�N�6�!��
s���JD��{Y�drFF�4m�!�R�Qb
D��a�8�2�E�*b�!��3�`�3*�>��]P#��k�!�d�:F��-Rs^D���%FF�.�!�Dm�081d����JB�	��!�Đ�p�"�cX�:Rm`T���}C!���5>t%Z�g�1�<e03'L�J)!��e&�A��R�P�سfA #!�D	�a�)Sc��$=l|�Cr�R"V�!���6�����J�B2]K#�Z{!�d�2<���[��W�J/�=8�ϐ�ud!�ď �
��,�0p�Ƨ�dj!�$Fg��g�"x
%'Y72`!��TJ���#k@�Q�Jh"��Xv!�d4#��0"��бY��[C���!�d
�0�z���M:6�\e��R�"%!�	�ISttk2kE���5����?!�$\XfI��kG�JqQaß�g(!�$I�k{���!�)=�$�۵;G!�%Pd�'�	@ݮD`Abu�C"O��S��7L�&|z��]�Ol���"OT��®M�Wa���d�F�f�Z�ar"O�i����k��#��7=߰�"Olm!��ư\�Z̹�G2��}��"OR@n�Eb~L`G��r��u*�"O>���A���PUX�%�5fU���"O1�*�	m�8(�#%�/N�����"O�����Jؠ��D�C�pYc�"O�y����3z�Q�#��8M�"OdT���Ů3�0��B�0?���C�"O* �G��}ҕ F�0�t�c"O�H˲A��h�N1���	)J���T"O� �ɢ���T�b�	��hThT"O�D!�$W#
m�$Ifd�B�H�Q"O9�&�ݠB�٘�)�8X��"O�� 7k	(���u�_2E��w"O�D2���j��T8ug$&�y��"OX���	
�~��s)ǬfV�Ñ"O��C�.�}����
�$��"O<�#�!�U��i)�D ��Xa�"Ozy���.%��fE���*(h�"O���D��(���
�c�E�|�{4"O2�Q-�;O�z�y$�?p�l]q�"O1!&�1U�ȹ��ɛ�
�N!�"O��j⭚\b �	�Q�w��bS"OJ�Kcf�	
���q��ɸ�!6"O,m�G#ٹ=��jVE�z^"H@d"O���E� `�"�s`jөb��S"O�BB��1�����ߵ�P{�"O4���B=\�=@0ȅ�C���"O��i�o^VN=:��ܹ���"OL82��Z�M��$�4�ƨ)�@�"O��#�(B�P:td�p���j�"O~p��l�N�Z�jAB"O�P%�.,���ZQ��1*���@�"O�h�cI�\v��a�*ڼ}�sE"OT��W�c���4�8x�)h�"Od����|40���V>r��(A�"O��HF�]�A P��s��(<�`9[T"O�� ��mʵB�6�0��"Otȫ�lK6�"��+��$i�d�"O��pî�
�.�;��LR���"O�@h#�H�p��\X&���t�h�{p"O�%���(֔hⰁ�D�h��"O������S~�Ԑ3 �/�ց��"O�|��G�S5�<C��F�<�F�z�"O�(���E�w܀cQ�4
� T�3"O��䇌�B�Zٙ���`���	d"O"�s��b�d,zR�	%�l}:!"OX�{!E�gE��H߉Y�xm�$"O�]�!�.9�x`[D֝�j:s"OƬS�T3
�<��f�_�P�D��"O��Zի���F��&n<`�Cӻ�y�R�	l~�{F�ӈ:~Ԛ M���yo
�PmV�+Pd�
5��S�eX&�y���0%#�-�qO*yX&�{��Z�yҎA�b���s� �[�L��y�d
X�����g�Jy�E�Ϻ�y�ђrL.p"$fN4�f�1읦��>��O�ٚ" d�$��Bf�5�r"O�mؑ� D(!��Oê,���i_�tE�ܴ5�2���i�)N�M��.Z�N�����?I�F�-�8aqsNW�P.�����M}�<$�����b��h���S���4�չ�B䉾9��T�w��(6Y�"���2H�`l���ƨ>in4�(U7^D�EI4B�!���O8@ P�ǬF���ϙy���6"Ov\�Q��� a��h�K?]H)E"O�����5�رq���>%��@a"O�}�� �Jm��gM�+�d�ab"O�;�P���=�� "{�
��"O�iR�#�$z�R���J?p�9R`"O�S��f�6����X��i2"O���4��
!��q���	H�1"OV1R���{�9�q��6�m.�yR��j�Ĺ�ҠA�BT���[>�y
� ���b�_�m�7ȇ*K��U3�"O�9�`��^N����ǜ9d	8]�"O�� GȌ�s���
Ѡ��~$�P0"Od��!�P>I��O���:���'���U��P��Ģ�$��D��N� z!�dB�D%�(J��ņk٘鸴��#[!�ӋiҮ|w�� 62hQb�òM!�d�/M�޴#��Q�Jx���#P)F�!�dԷJH�hvoX�Q˘�T�T{�!��T�|�j��⌺ZP���?�!�d�v�a��@�9:M��y�-�=�Py�_�)���T�G�R�HIQ�)�>aI����X�Eߢ՛���q�l���3D�(�,��`=��cp@�AH��)s�2D�x�@)���ʲ�x��(1D��p�M	%��B�F�27�hp�B�+D�\h焂� B���m�!a`��T�'D���2�ɔD�*=�Ǳx�>���f'lO2➰�7�вF�YAÐ�"5ʝy�!D��˶HX><�J�U�S+D��I��L"�t���Rτ�*�m�W���w!W39\���	x�0��>�­ك-Z��8iGzB�'��M�T`w_:x��V���i�'� �F�-�HBr��
�Q��'ia���K��� ߕSW��Z�&U��yG�;3jt)ֱ3��|i  \�y��ю$����B��%�f�@0[��y��#u���p�D�RDN.�y����)J�,w��	�+<0�=E��g�`-#��,\[BU@��Q�u5Z��O�=�ң��6� C���_ �'��A�<�,�a��2��=|h��Bx�<1��hJ���0BX��l*Q�CN�<��M�>wr�t[p&D!�h���i�G�<�Њ�P�\B�\�܁��N����'F��K`oR%z[�qj�
9z 0
�'x�qأ ��x�r3Dc3���	�'0r195Lɡ+<�)t*��D��'
�S�كc�����FҼ=����
�'�\1�H��!JqE�ܫ2�0��
�'m�e
�i��ѩ�=T�q)
�'�0A�@a�W`��
��	
&	�D��'�̌R�拙H��T! 	&-2N�3�'����an,4KHX#��(��,���5�S�To25K�-���P�H���
�yrm��n�n�i�!���R���mƱ�y���C��uFW1�>L��jĽ�yr�αV~kG�]
��� �O�O�=�O�<��"����)4�	*���+�'&�;6�>8<%�c/ω$ժiv�)��<�'��n` �M�L�tY;���r�<Q�B6E�ћ@͎�(U� õ�q�<��#]�~�2%����\�0�C�C�<��DA� ��p�P�#�5@�b�I�<it�@�8U�Zr;�mD�G��hO�O�N�+Rd!���`��*�� �'��)��J�NW��3�
�7�`0��/�H��	�Jy<���_�r�d�f�:e��B�IvQ	RA�8:,����`��5��B��>u�]��ʶv�\9��d�9�B�	�&c �Ѐ�&j�DT.܂L(�B�I�����CԅQ;D��G�;c�B�/t�>T{�̳26L�Q4@�q��C�	�!�`@�6  }��b͗&x�C�)� "P � �'( ���E��Xg"OZ��3F�
o�`%��d˽q��9P�O���dP� ��aa�Y�}ꑻed. !���9=�-�g��p.���aČ.Tw!�Q�D���fTU�BIN�!��张P��G�Z$��j�ι
�!�dI5#6�P�$���
�-f��#�S�Ojz��CIB&w�p�p�F����
����*k����Bg�����k��	�yb���L�b�!#
���)�����y(<oY8������@��6�6�y� 08��X�{�yf�����O
"~�˟8h�a��ʛ:gf���%%DF�<1!�ƮU�ݱ�*�:$��ia1K�A�<A6�A��!	��?jJ�Hw([G��@�	T~"�C�r{�蒑�į{���p�Q:�yҪQ)����'�.(~]aA�B/��';�z�旑x�:��5��U\�쐥����>��OZY�uB_ 9;�A���'1��\z�x��*�'֚�����!�8:�� ـ؇��V}��>!E��(������"^A�x�.�z쓛M�˓#�`-I�G]�P?��A�-��ϓp��"~b��_�:"�����_�8u���syB�'a|R�C5��]j� �~`�!«ű�0>�H>A��	�'�x��!*����A̜k�<�FV�Qƌ��)��z�N�(�m�g�<1�%D����$&��Wx	H��Vg�<��Q	���b��?ɋ1O�e�<aI� q�X(����kSr�FcBe�<S��[z�(A��G@���Ō�d�<�bI�In�D ��wcW�Bj�<i�*W2���3�ѭ@�P�0�f�<qd�Z�d��0� @Y�2�B�ʶ��b�<�$��3��1K��k���JQ�X�<i��I�%�ʍ3L;jVx:g,�{�<���!=]��Qs�R% ��g�u�<YwȒ���t	^c�h���p�<i�-C}��A� D�(Z�����g�<	1%q�~x�7�E�'�l]�Ɓ�n�<i� �!jK�E04H��0�6 �e�<�4�e3�ɴ�N���C��J�<Q%�N.���ψ��Uy7�QE�<)�F37R�1A���G��=ɲ�Z�<��[�R~Xa��iI:o�@�0��V�<��팜*��9w \�NF�`f	�T�<q%Y�4�膉��9c��#iHI�<��E�=G@ qã_7H�h��7�	I�<I�JG:b��:�.Μ= ��bBC�<�d���Ax�LITUQf��PH
A�<9Q�8?D�i�g�=89��Dd�<a���w)p���.qk\�W��\�<i�M�P)Y@K��:���Wo�<�ġȈ)�d b�AQ&�	cD�j�<�S�`�j5�ᧂ;P�*�1�Rf�<���G���q@�ڮO��F�d�<q��iε�`���y�4�K�z�<��#۽h�0Q�A��o}f� ��[u�<Q��ǷWe.@�,�Mp���o�<I��j�R��c���U���j�<i�.�8.4�}�b�#-���#A�P�<��k؀G��Q�6�L�gJ�<�q���Њ�Ϙ\�"%2�E�<�P��J�hi��O�m�왷�g�<�g�
�D�l��(��P��Y��AK�<� �|
U)$�0�)�X)V�yH�"Om�A+��UT�A��;J�e��"OVxp�M�ݾs�v$"�T�y�X���Z�b��@�� �ܡ$������q۪�����:���酅�4:܅ȓ,UX �4 ��(6�!ˆ���I���Y�%pd�����Y�B�ȓc�-��U�6��y��D�g�6͇ȓ�, &f@~�����e��T��&$B���:&��z5��yI�E��+�� �"�.Pahy����*/`��ȓ 2u)�OK<*Ҭy"dO�cbB�ɗK�,����H@�Er)� oC�I'�ȑ9Q�M�:rܔ˖F�<;��B䉼{-ʄ���WxC��S�gA1$�B�	�;Z��EQ& o~uiB�߸&�B�ɑ��H��5J>�@;B�ޜp�B�		Ip�����V�E;PݱղB�	�vԑs��_'��i�E@��B�	 4.�0Wʊ$:نq�n�8˔B�	�e�6��UB^3��eխQ��B�ɱ|B�ŁU�J�dh�W�T[�B�	:n �zE̗4J(�XFkH��B�I�O�֕�#M(n��{�d�_%�B�Il^�� ��b� �2eFʠB��jHH�c V9dʼ�� f &B�I�E�~$�w. p^�d�����0B䉲l}R-��&A3|���@�G�-� B�� 8���a�މ4�v�CG�C�.��C�	�6��5�DY:���F ��C��0_ �H�aT�'�&Lq%�W��B�	�r�= ��]�A��\"5#(<�C�	SY;1h�����	�rB�I=_	tHzDF��6eb]kc��#�C�ɶhw�(� �T�T��!E9��C�	7Q�-P��28t6!��I�2��C�	�I&v%� GB�+�$�xr�7�B�I�H��i�h�QbY��i��5jLB�I�+�A�%҄{��:��D�h��C�ɥj�I��KW��H����ƽe��C䉴,�8�x���Jv�a1cY�no�C�	El}b�M]�D�]�Vb�Mk�C�+R*|����M�@���R�jTBjDC�.3M���6	��A!���07�BC�I��rQ��D[�=�e�|�C�	<��dl�q}�i[f¹[�8C䉀e�в��Mд5��K��pC��2�v��*RD@��A���C�I@�l �) 7Q��c�͍�2��B�I��� ��ϙr���%,L�C��C�� "�$�����>*��=Q�.<^"C�I����K �Q�|�I��F�iT�B�	�'Ve��k�9%�UXFo� O��B�	�2`j��8ߴ��C�Z$8C�	�!B���h[�+hƘ�w��:,��C�	/v(���U�P)�ިR���>��B�ɵ���hE�H�,�� �$+�8>�B�ɫ1�9Z�"�5�� ��݇e�B�ɫf�Tmۅ.8����f�>�C�F�h�ըE�L��@��^�0C��4R�^�1�-�cz��˘�Mg�C�=<LB��T�"a6�b#��(�C�IV��l95��p�f��v��y�C�I�pHd)@lY*S����	p��C�)� ,<�G���eT��xJ�"OB�@ѡ(���g� �R�bq"Oh��g֪uN�x��E9W~����"O|�5�ɞX
H�GK*b�0�d"O��C#�˽\��E�K��?w��AD"O(|8F��E(&̉k�X�T��"O�Œ7@ǚGJ���oP.	�@rd"O���Z;Q\�X�ԣ�) ��"O�,C�zG|����=�z)��"O61K0�ڶ4Mش�.��&�"OJ�ao
�-F4�yF��,��"O6e��ꏟK����#�o�����"ON5���дa˕w��"O��uAZ\����jud��"O����&��q�D�pWc�"OV`c�HC�F���$
��N��q�"OVͫΝ�a2�Br���@<���"O6زcfD|�V\�u'�WW��ۗ"Od�C�Y�>��Mأe�:X݄���"O��{�+Õx��$rDA.6¼�)�"O�	A1��~m ��� T�T�1"O���u+_	m:-�1��{O�|
g"OBT��-2Y����k�UR��`�"O�Q@�ė�6uX��Z�2�9s2"ObD�a�F?_��##H+)H���g"Or� f� �[�Ȑ��lX�CF�Z�"O��YKd�Pԑ6��a/�6"Oи��M_6?�I& )]7vEC�"O�Q*dD��_4�-��/I���B"OV�Aǐ�N�<2���$ �"O.���C��y�-"���`:"OV�X�K�#��4� 01�BD��"O2Q[��܊jR\��A��D�9�"O�\� �C� $��0`�-���"O�5��o�?o�mQ @BAl��"Oڈ6��h�&�"N Afp�"O�ݹg�<+�de���Տڈ1�"O��	D�Y=+���6Gòo�ά�"Oj�Ƈ�3)o�;�kJ'���W"OB4r��crjQ���@,b�sS"O��P2a�o_<�÷�_r>��"O��#��՟z���B��ՓX�P`20"ONA!ף�D��A�&E~�Y��"OZQ�c/K�?��l���1z\�,�3"Oxh�U�`!�v�ڹ!��Y�"O 98uE[����IP@��b���@"O6-�fa�.t�Z�����BV"O����CS7U��@h�.!0��tS"O���	*xG<�����;���z6"OxP
1��x�x
d�N��܊�"O2m�Qj �yI.�k�͝�6:`R3"OaaAhC�B���'E|"M�"O
h�/��>��y�IɆT��"Od;��
�1#�T�0�J�?d8YF"O� 숵F��af�9OD@��"O�� 뚸�x�H�āp/��	T"O����1j�2 {��#A6�"Op|Q��%j�h��Q7Hy9@"O^dW�(`$`�B�0�@(`"O���%)�Y_�er�i��I� ���"O^��1�e������#]��k"O��,K�;�N���ץH��X""Ozqq͟�#	�މ,�nxk�"Oz-P�#�Dx6�]a"pX��"O� �k��T����K�B�?vl�"O|*�_��Nx1� эd��3"O�y)֨4"��x�/zS2��&"OZ��&�.8w8cp�RXb�{�"OЩ��c�#`Fm(���,5����"O]h#���^1J��W�Z� a�"O0���d�85��)a���00�	9�"Oxu�wŇP>1��h�D���f"O0�XAn��Bc�!��u0��"O���A>H_�иtc��pd0%��"O:p؇cM6%�V�Zu��O��yr+Kv��"�$φā$�K��yR�?ZQ˃�������&/�-�y�E*e�n!���p��5�Ul��y��� ��MǥV'E��E�y(ŭ� MK��Y�CD��4�6�yb�(�!��ɜ5:/����J�yb�4�@CF-C�	I`HJPa��y�ꉩR$yy���y��٤�T-�y�E��)ڜh�� ��D�	!���y���S�1TNO�s¤:pe�y��fI~m����f^du���)�y"�R%��e���6���Ǣ
�y�N΂&� Q��.&�|��N���y��אE��:ҥ]�HLneq���y'Q!�����
Q�����'Q�y���&i�@����F�D9@F�#�y%�/��9s$�8qT%�I�1�yb)
3�議�$�FjԹ���߶�y��;q] ��w�э7_����y�C��(T��r��� �zpQ��[��yRD�p X��I�e(����\��yRϕ�D�R=k��^j�5���y���l �P��aZ+��.ޖ�y���>X�TӠNCZ����y�*�f�fY���E ���>�y��-+�XR1ô6��x���_��y��"{<�B��]�e�NQ�GG���yr鞽]a��@��2c܄!f��y��F��x@P�E?/=~�B�&G)�yRLC�K�P�[5�ݑ.HT�;G�9�y�$�N}�[��΀8���8wIH��yR#�M�D��G�31�p�g�3�yR_;32������ iH��a�ި�y��I2z䀢,�r���QD��yH��3H�9��Z�m�n��0�2�yr��3(R%Ak҅vf�) ��y2M��d ��v���l��0Bp�P��y�cH�
�e��%vc����9�yb��G�.��B!J�<a6��C����y�d PU~1Z%F	�-�85�"��y�i1�MH���-�5qR(>�yBFN�.Htcr�J��`�y��"�r�&g��}��d����yB��&6]V4@�'	nC�i���y�7"�v�hᭅ�tӀA���#�y�g�4{�)�HD(l�-*3ˁ;�yBH�Y/�a��C�o�^5�⁀��y��Cbf]b�dF*k\
#rC��y"*�E���r���;P��?�yb��C��+���|�l̡�`Ղ�yR��&���EzкE9���y�X�R��P�3�N,K�g��y"O�3���A�f.�"���7�y
� 4�SL�''�����%E��ة&"Op�1�kA5��mI��E�֡CP"O�� �@�T�2���C̗;��=�T"O�@它!	,��{��G�0v��"O� [(�b
4��F	)�Q:6"O�*Do٣8�@�+��7r��p�"O�x	e���w�P��䃿^�0��$"O�TBԅF���yz��ѥJ�t�"O�� w�V<s������W��*�5"O���+�LO��y� ��n,]P�"O�XKT�,�����(Kv�,�6"O��3�Nͯ'D��XTk�|V��"O�`�OP�(�H �*�6@OP� "O���1g)BG�E�`�C���T"O8���� !�h��g�>��&"O�����y�b��á"Od|S���&N����$K/CR���"O>,R��)�&Q#�Ѹ�aj�"O���	�0��K�k�2���R"O��UhAR&H����Վ.ǐ I"O�4�(��`��8���Y��, 0"O���&��$3~�p�*	�{��:�"O�u8bgD�ᠨ�e�|^�	"O��)�h��!xhp!���`a"O�M0��y1dM#�E� -�Գ�"O�<�W�	G(v������0z��24"Oj��#/�e|%1��M4��T��"O�x�gM8i���I�o)Rjh݈�"O@p��! �M����ѱR`��a"O��9��\����eh�G�e� "OZAcZ4}O�� hכ>P�X�"O.iJ�l NM\�������aT"O�d���5|� 0s�)GA�USR"O�ss��F���G��pH�w"OzyЬ˾ { �aB';.�f�8�"O��Y�O��bn�Z�
����4"O`�(OX8x���O,/��u��"O��2U�˽��C��|z!�Q"O�UӤ�:1�r�R�BE�Z
ذQ"O���� �GdL!�!��
�G>�yr��a#��)�!������ ���y�I��;V�!��D��5�U��
��y�I�����	�VX�c	��yr�[���J"ϵ�B�jc�ρ�y�o'+�F�y����5C䤎?�yb��h~���"�!����t�N �y��חV����bI߮k�����͏�yb̏'g���פ��_��%��\2�Py��]�9�&A+0	r&Y�N�h�<!���e��U�z��k�EJ�<���;!����l�*O�u�E��E�<�`�-*vy"���r���B�Wf�<7�RF�x��J	�bذR/�F�<y�
�Mz��v/��J%��P�OQX�<q����:���2Ⴠ-��]>�B�#3�&��� �*��y�ъƛ �rB�ɪz�\Z$��.dO�Q�0c��a�jB�I.5�4��1
�\��y�
ޠ�&B�+2���7(G�@2�T[<7WB�;Y�΍xQ�5H�LB��N�C�ɓ5��LQ6b��?06���`�� ^�B��5�.�R-�3]�@}I"��y۞B�	�?�n���A��u��l@�
�2m2�B䉐�H=��a��&�t���,{QDB�)� �z���@�6x���/O/Z�9�"O�\(�.H�G,`-��T���"Oj�[�h_"/����W��$���˵"O�(El͒b��t����a8��p"Or�Є\�y\25r�����ţ�"O6��#H̘��uj'y��'"O��㰭�y�0\�%�.O2X��"Oz��-�Y����(+>��s"O��U�\��FQ���Բ7o����"O�P�c�U=&"��p�BU9����"O����]�gZ�'-�Q��3�"O$` C[zø���+?� ���"O���a�>p��Q��9=�n|""O$`@���A��{�IfAxd"O�H00��/�2�!UOP�@ �V"Oz�K�D�e�ā��+�X��"O��aЉϭcˤ�X��O5~�!�"Oִ ��P!V��(�����Tz7"O�P�OŒ&OЀP�O�::8�'"O:�P�+�.`W�Qq�ˁ񖅫�"OP+�*��:k��)�0'�ر
V"O ��$��dCF#�*w��MɱkԖ�y�A�AQ(X��=i����*�y���!R�����&P��p"���y¯�6�|4�c �<9�5+@&3�yB�[	u����dk&0��\��]��y��J�=������',���` �=�y�!�. 0#��\1�j4k����yrh,7�@�Qn�?.�h�@G���y"�׊_L�i�@H�o�BD{p
J��y�I�-��Y�0�$4bVL�Hؤ�y�a�Y��q!���$g�1!g,���y��N�k |@��^�R3h�ض�E=�y�nM�h�ׅN3Myz�x����y"(V�n�N�8vMQL�Q���y�Γ=~S�"7�C��Z���;�y(N�
�l2�# �.��,p��	��y�N�_��􋳪�0��ၣ���yr$�+/w�z�Aӏ* $��1�y'�%E)z���d��U��P�aB>�y�ыB,�5p%��N(���̟��y�iΉz� �x�n�8L���3�5�yBiʂI��Cao1*P �0@(���y�ݘ�Ա�(E�+�@h(��¾�y-I�)���b�'V�"=�]�f���y�e�x��}�����sܴ�����y��F2E��$�ȴ�J}*���yRg� �X�s�΂u�@ �h��y�#ҋQ�ށ�^�Ba�kތ�y"���*]#-׏\)*���^�yB'�P�����e�dYi4F��y�(ӽk���j�6	D�����y"��*iZ�����U���{@�3�y2�[�-��@C���O��D���y��ߛ��)K�+I�@���0GL��y��V�! �d�8�"�I*���y�#P8}���ڟ2Hr�Ӕiߧ�y���St�B�"z���:���y�n] � 
��W�v�ٱ#�H��yRG	�N�2��j��i:s"
 �yR
]�si^�X1툜0�,���<�y�j�((�9��*S��*��Ē4�y����*�(�ʄA�E��IkQ틅�yRe�+{�p�T���CO��$��?�y
� .8"b5��D��G.X����0"O�8��bV�]���Pf��$-���jW"O�E�х99�Y��L��j�"O�$��q!pI�e�3�TT"O
䀓Æ�:��z`K�&o�Uc�"Oh|	Ռ�?�D�PԫX�`��:V"O�`��퐃R�b-3�>�$��g"O��B$ăo��k��{�p�"O*)�u��'�$鷥Z�-�ڀs�"O��(��>��H�����3¶��"O(��O:��4j'�Ϋ	 ���"O��K4���^�d�	҆��Q���"O�Q
p�F'�e���PQ����"OaA�]�2 +���UH��c�"Oth�
�42F CbB�(7��7"O�5'�ݝ8��9��\�q͖�
�"O�ebw��;;r��R�
�\���"O�}B��!*%�2�L�|�@"O^\3E�A�G�S�V�) ���E"O�
���+=:�P!h�� lӢ"Oj8��U�bX�p��L:b����"O����r�<9q.Ëy�>��1"O�1���+/��b&Ga�(9p�"OFx��-�+Z��,�	Ԯ\�t!Q#"O��82H1d���1*�*b�Li�"O���[y/��&IS9|�>y�W�q�<��$ZQ�z��$^�),��+p�<q��X	P�yنoܫX?�LR�k�<���3GL\`C�&����c� _�<q��ku2�N�
^�ju�W�<�ԄN�t���j�MևsHƙ:��<T��['D�P�v�js���%�D�b��;D�40��>;<�RE ?>}&����7D�DxE&�@��C��\3�"y�$�4D�l*"��x�<�d���#ҫ0D�P�댁�&�kcةz�N���i+D��!S U�7�zu�ҌS�C��ĈT%D�(�5"^�r�KV��#=}�4s�a$D��*J�X��83��T�^�Л5�/D�(��� oh����h�v�~�R��-D���d��FNм����D7�q�6D���Ɓ�T��4K`�4Z]�-�i D�DaS�S�'����ں-0�i��&?D�\����+CJm���O��Q K;D����mL�l�ɐ�oI+K� ܀m7D��@7��$��l`���.\��%�#6D�`���K?�i��Č~��)�bi5D��B�K�0��#�@���ap�3D��qF��8!p���eZ%| �$pb�=D��#%O�32�l��bW�y��405m8D�h�㖟$���1'�'���ʗ�2D��G�S+;���1���2}�f�k��1D����i��5��5Q�K�HM�f';D���dM�iؐ<�ԣ�A��9D��"�X�v�z���!q��}z��:D�p�矏5�̩��B�ɳ %D�H@0�ՓSϲ���(f8�@��&D��󵏓�H�,)�
��:/&��'(D��� sJe#�f�eY��q�%D��ks�Ӱ�^q���
@.�L� �$D��P	�a����ɗ61����!D�,z�h�`�|��TE +��%:D�H3��׍(b4�6�@:0W|Hk4D�@��ѯq~��`�]�UL���2D�� ��i�(H�N�0��թ\<4A"OhB���:b?&i�"�8m�(""O>�;�
lJ1G��&��"O��P�I�m�\���"��{�"O�\y�Mڬ.R\�葳3x�R "O4x�C�F����I�,D&a�@"O�\�שކd�y���S�4UnD�T"O� ��N�	T�^Ij�枬UHi�c"O^�a���	p���*��$��"O��c�)ۗE�h�)�揊[w^�{�"O�HѲ�!��Pg�]"&^F��$"O8X!vt���0IV?-|XL2�"O( �b��6t������	/wv�ȧ"O`%1�C�B�>1��� v����"O�����S�θ�M�Xn8��"O` �ao��_�M�3+�>qG�=8�"OR���+4o��$��<u���Q"OT��g'�4:]��*�1lv>D��"O^cc�^*xДItj��7�����"OF� Dg��a���i�b�q��"Oȵ�S�ޓ��� �!�Z݋D"O��c%M�l![��L���c"O0} Q��g�d�����dZ��Zc"O�,���W�+��t�SN[�JT�["O��3�V@�	-K���ф"O��'�̧Knb�ƍ�z��|��"O�|�P���B7��:@���rậ��"O���b�5#�ސ��=>��-�q"O��!��[�Xwڐ�%)Z�O�B�`�"OD|� ��	��I�t(P�8�d v"O`�Gi�-H���hO�l�q�"O�% @JO���]q%H�qr�B�"O� +7!��E�"��fX�k5�ȗ"OPE���B ;�.[+R��h�T"O�����8E��T:v���n��Hs�"Ohݰ�)�)!Nl!@a/�MxP2"OƉ(�� QM����.^�Th���"O`�@�t�4z4	$1U�T��"Oi�s�ܻmc��pK�8��@j�"OR8��͊=R���;]h��"O�`����/4�	�)"x�1��	O�O<B�P1��Eh �B�'�� n���'��<���6��m�sB҃�~5p�'.�\�1+D�Zւ���N�6 f���'�ht � �M6���1��"�H$��'��d�Sn��ȂV2�ʉ�a��g�<�'�/ �тTfC)fPDq���Vc�<�����6X>d!���D��}H�-�^�<y`g��`����׌<\����-t�<��(1��}�Gˀ$C���!
n�<y�Y�;��`���|�^(`țe�<�d+@q(�A`@�9vUpS�I�<Y��H ���"��e4�ܻ�j�C�<9��C���I
򎞸_G� ��$�A�<A��X�>��`�"/��=����}�<��ˍ}2�4�1�ԟ��S � p�<��.�Y�������J���.�g�<�`M[5TZu�ʀ�"q+com�<y���"&�*7��� E�h�<)�jA�d��"V-]�v���+A&�J�<��.*i���ԩRI�?36B䉠F�|pN�:��Xv쒉z� B��=9���!���m7�8{�m0=?�C�I(:ͨ�f�V��3ya�B�)� ~\P7�V;B�$�r�;V��L��"O>��w�	�{�ڤr#�F2R�Z19�"On�(v�ǅ`K$������A"OV(RFB����<� ���q��"O����ܵ?��2��F�4N6{�"O��ÂnΝ	d�9�F,��:�"O��b�/�Q�Z�cr#J�l��x�2"O����a�g��볡�$m��� "O2�P��L�CS�ER5 Q�@׼�x"OB��v�.4��˕I��=�:\��"O�aC@הPX������)��yV"O����.�'xfl2f��@����"O�14� �5ȠpP��0H�@��R"O�a��@�C�AH���r���"O�L"���9�\U���܈w��3�"O�qB3�49����Q�{>�Y2 "Oh(Ja(�~���s�W�T֡Z"O�y{�*ڎ/�
trd
��dY���"Obl�����I�6aB���/��x�R"O���I�vm�$	e� u��qP�"O2(�RH����:>�$���"O�2Wj��JO�����4��`1"O�$pD��#����lK������"O�U�fI8�,'ˈ�k��Q��"O�]�3NR�z�xa棈�|�,a �"OHu�4I]T�ԠJ�?���"OΨ�j��K��8(�J\d��r�"Oy�'�P�s4eJBϋ�H̀�4"O��9!,�+�U���Bi�C"O���m�fx�<r�n�M�%�u"O�<t�!��a��v�  !"O�p�׆Q�1���4��5)U�"�!�dH�Ul����� W�5qBd�213!�da�i���W�"��(��Z"s!!�$�7��=��)I5��� QoD-H
!�F3`�����2y6Fd�5.C/L�!�DL-gꥰ&�G�M3���&�S,>!��H�9W�`ؠՂ(��pj��!�dR30��Ъ3�ѩWS���HКd!�dx孑�g���y���ɟ8�)��gB��;"�WZ*�v���7�\<�ȓIҶ�I�e�9��q��>`� �ȓo�U�0�O9B�������V����C����!/�8��- ��3����C�J+��>�`t�S�I�]�Ʌȓ
�r(k奒�\k&��w��9�&���9�B1{ӯ�3����w��3IR��ȓv�4���GL/!�D�i��,��Q��7��E�U�A��(���p��@���2�F;���BPFԇȓrl���I��:a8h(�#�DjH��h�����@,�����#����l($9�'n���D�s���΀��7�Z�hנ�3Lb8;�GO��ņȓ���*���T��mZ/��@�z���W��:gT,"*�ABf�ő�m��<v�1����Y���)֧RZ�ZH��/����/(5�4+P̒�����e�FM��G(TM��NӯC�B1���h�ɧ��+T�&t2�A)�&P�ȓS�*!��N�kW�����X��4$I#��RpY[�/STS����af�H�$��,2�vcw
�E��h��F@�![�M��,d:V�u5�y��S�?  u+�E���A�Ǎ�(b��q��"OHE1�o���(l4�ɓ[�<�I�"O�QP���t�8x8�ϱ;涅"Ofh1�D_�i0D���L6DɊ�	�"O��0`��X�������l�����"O��Zr&ľ煝�'�v8�!AB�en!�d��K���q�T0q�N��eI�6Sk!�Ć>^D�Ö�Έ>�,�r�(�� -!򤁺2��F�|��4�7�]0!�D��N��S�&�3u�F�" �ֳh�!�D\K�D	bHS=u�h����֮ �!��[���Q������UZ0	�|U!�d��s�������}�$�'I� ^U!�$җS�,�"��h�Q!�$Xh�ht�Gn��TZ�'V7!�DC6j|-:"�7��H���)!򄄷u�Ըs/&JΖ��e��(T�!��'8k�#�J��z�֩G?!����̹r�X���p�4�N�"!��;t!Y�ATb��D���'<!��C�j��@8�튓f�JM��i G�!�P�I4ـ�&�3, �ȧ�!���-<
�H�/�P�i�FG��g�!���M�Hk�H�/6�x�$��,b!��ʰCnf����H�	��H+d=.R!�L�NN^�a4�RU�"�i�54!�ȑj�R�T>x��h�5�U)_$!��7W(,I����J�^����Og!�.ۚ�Kf�.c�`5ys�M�&_!�U�)�L��I��=8���,f!�׭S�����I�n��I��]K!�d\�?��`�lX�I�:��߮nc!��W,1:�9� *�8��E�,jH!��ϻG���P����,��m�.!򄎺u�<8�f��]�Dmi"��!�D*A�8�+6"�]��`��Z�]!�D����@sVb_�V�<�#��:|�!�d�:;hT�ckէgC�+׍Л�!�D�&;�l��ʽuY�2�� ,
�!�dη%\��2ᦂ�t�x�p3d�[�!��F8E��uB����"���"��[�!�ܿ��yx����Km���u�H�'�!��1+Ϻ@��� }�Uap��W�!�҃[�=��₠_n9yTg�U!����"$R.ܴSup����T�!�$�s�8�;4+Pz9ȹY�Þ�A<!�0/N�㓨Z�V+���O�O�!�$����!��ہhX�c��2�!���%?�\#��k�P�LY [�!�D�O2v@2���'��"f�*�!�d�3A��(��	��2]�$�7�!�Dõ=�!C���.E����IE��!��H;'=�t�[��̿�!���82����(�+i�
��密�:�!��0���Hev�|JFO
�\�x`��ox\A�.]�n�}���+�"���N�|,K�D�y�U�I*}E�,��/�R�Rf �\x�$�D̈���ن��)���l�����H�,�ȓ{(tiu&@���H�0��#;T-��<.��)".l|���
�AX��E���c�^�7�!���i�&P�ȓ7���6��.V`=@�G�XL歄�lH���Y�G�*X@ǩ u�L��S�? ��3o�'@ް�Tn�S���A"O}˴�v���MH�C�X*�"O�� ٠hm!m����"O�]ٗ&K'Ȕt���ҋI��y�"Oz�Sba"MD:�P�AC%>�2�"O4������D����ӡ#�F0��"O�5S��&�X��-�V����"O�Ęfd͛h��awj�r���C1"O���ۿ�����bz��SA"O�#���MDA��Lz��H�"O�m�G��4eq�FE�0s"��5"O��C��C�d�r���!��"O����� E�2����]5EE�u�3"Op(�߼%��Mx�cW=E;b"O��b��G #J
� ܻa1 ]��"Oj�7�A3L�@-0U��Kn�@w"On}9G�4��b�K�=��PX�"Oz��C��B,:WM
�t��*�"O��ǭ��=��EǢe ���"O��CF�-��$ �	ٛuQ"���"O(h��X7�@��7UB���"O�T�'M�$&�(�`��'W=����"Ob�8#�J�
(��tሼ;ٺ�"O4YǩL��&YCcƸt�����"O�X!��U�2&F���.\����"O0���i^����G-+�Xh�Q"O �p��F�b��m��O�-���#"O��R�$T;Du�D�
*6�(��$"OZ9hs�]�z�0-	��4R�X� t"O61�D��$S����'m�6i��$��"O�M ΍�����8F��Ce D���pC̸m�F����Nr]�ť*D���橅�,N\{�,G�fv~pS �+D�܃" .P�� 3j��|��a)D�0���ş:Sv�pELBN�&��C�%D��`�Twp�$��
U�4B���yBF�M�l�	���x������y�ͰVS>f�͊����y2 �28`h��\:b\�c�*�y�]l���Y�f�}�V�h��� �y���#Y���8BR!t)ҭ�")���y�aɫ`� =fh�Cߞ������y2a�"�$���:"y�Y��y�CW�4
�d��I��(���y"f�7����V�m(�pA�V�y�8_D��v��d��y��߿�yl���~�CmM�uQ�@��l��yr�ܪw����m�(}��8���y��ܴ����W�o�>�8��	�y,�FD̻a�Ƥb�"A�`�	$�y�-�����5(E0fQ����j��y2D�h
j±�^�cW����m5�y��
o�֤�5ꓵE�|]0'�-�y��'e��(i��ԭ����e��yRʘ2H$$4̎;A"9c�N��y� R#qzp�"u�F����C����yr���00T�{��T�)�+�yES�@���ٴO�3�����FJ��y��1�Ĵ�ȓ~L��'#݆�y����0�45sf`���Ҋ�yb S+�٩p���rs$@�v)5�y�@?�)�
� �0ia�n��y�,U�05Q���z1�������y"�@!dt�tFZ&k=>�
��^��y
� ZTZ3ѤY8�k���$����"O�E�u�f�	�@L�Tʊ�`�"On����X	y�&psա����C"O�q�uK��XR��S� ��:$�p�"O�2G��&�^�ہ$J��
B"O������A�DA�ըG�x0�g"OT�ڵ/S dQ���@�d��$"O4%�7��&ff@�u��6yŹ�"O�
�Ǝ-U.�����,B20�v"O�cHL� fN�㕤�7B%�m�S"Op
�l��5�*��1d��O*@A��"OD�-,�|CU� �
�T���A�i#!��-9��h"�)�2S�Jເj�!�D�,D\r�OY�9�H]�0�\1 !�D��x=a��=����g�>U�!��+��)2�h@n�4	�ց��!�d�"eA�Qs�͢�x���玭_k!�$L��� X*ӴDy�D5_!�d�w�e
�M
k�����K�\!�^?(��p��^�&L��H�]�!�$יS澩
�l�2L�j��$�@�G�!򄇵"�� ��j�' ܜ�"C��),�!�d�=g.���MQb5dtځ�Ѓ�!�DW�	H��a��k+B�3��X�!����������iڸ=�!�%!
�h�EX�~Ԥ�S�I��J�!򤐩�)
�a4�����Y�!��R7��\���F�8�P�e����!��1g�����(Th�y��Ձt!�Y�N��0���dbnKuOY,+n!��t�h�`��)+b�D�0A�!�ә}Ͱ�9�"ݯlV�x�B�O44|!�d� K����Ε�f��(�4�!��;�� ��ʏo8�-��E��@!��X�[��4����p%E?O	!�DՏ*���
ń/i��%	ao��=!�d��b���ò�<>�p��@�	!�DΡC�* j!gU5A>�85M)D!���605xA#���>������+�!�D�9yl���D�Z�T<eJy!��6x���M',�`��h!�C���Y�� �[�y�
T�u!�$ٵT�1j��J���9���#�!��g
t ���\9CK�Z�!�����'e�{�Lē�IЏi�!�$
>\�B ��C+�HQ{��@�!�DN�8v�,(R�1%��A�h`�!�ć�o�B��&'�I��9U�_�/�!�d�:%�r@v�˳P���vbP*�!�d>PP��S�*Y���p���!�d�1afQ(��^�Z.ي��V@�!���H��P�ǂCFdd�QȔ|e!��x�t�*�"��c ���7F�
t!�=@�l�n_�KE*ai�GP!�D@�|Z������J���SDK�XL!���)]|0%��FT��z)㶃;�!򤘍5���i~��|)u�D�J�!�D�{�4�Q�"@�Lܡ��<_!�S���q�Z�EIx��(�&!�!�$R:[���"�i�f9^]g�Ƽ�!�D��X
a�.z��zc\6O<!�$C��>��CeXL�r��B�|6!����1�Њ��j;�1���(:%!�D	Y��h��+%��p�Н+!�� u�CA�/A6��r7�#:�p�"O���u-�<,�x� �0���@�"OnȚ�k�?<;�����6:�t!��"O*�x *�d]���H�8�HB"O�pH�m�|?�@ �*׿v{ta�"O�93'�D��rY�腈<r�Hc�"Od�" �#z<$��ř\`��2G"O���$Z�����!H�u���4"O�ԣ7��x�n�����P�*�o�<��o�I^ ���
2�F���*�e�<���� omaGd�S��S��b�<7J��L_F��T�ê%���R�F�]�<��Ҏ`�6l�� l^
����R�<���'Y����a΀C>�aY5kKM�<Y!��D�(�CT΅3]���
¤�`�<��+L�o��@��үY��e�E��t�<2�5�D-l*i��ʏ�7�ՆȓK��c��;=���퉽�Lq��m9�8����<"�a� �:�~��"��.[�l�R$�@?��-�ȓ@鲘!�C4"����}+A��B�@m�#�	#��p"R"�a�`�ȓpA�t�Vl�.|2,��f� u�����
�`�;�Y�Y.�C� �x
�(��p�h�csȝ�MԘ!��#ԏm�b!�ȓ"��8��d�50�@�6�[Ι�ȓc�6�JB�*o�sɀ x���$�،�w"ȭcNf�2��;o�^��ȓ	�t���8ri����KV }�y�ȓ3����r�]}D �f�]F4Ņȓ:�#�[
TM{���=e��!�ȓ]<۰�bX�3�n��O����T<����e��@G�0����j�hEȃ�_
e�a�!�2D0`��DJ��;��=}"q9%+�qsF�����fl	^���3"#C-s���]4DuD�æ@2	��n	&Rdʡ��!�6�� H.*��h��	R�1��d�8���E�"�.����@���ȓ ��@WN�#T ,U`��h��� \d9{��W�.�@St���� �ȓE�% F�	�$X�IJD28ՀЇȓ�����/���ePe%4p�,��.���BO�fҤ��g΍&XI��3ny�$�A�{՜�	

�9��=�ȓI)z�x� ��C�rL���R�fх�6�>d���Q�|e�	�A�{3p�ȓB$Ρ���Ì�ᑠަ��ȓc[�Txq�Z�M����`-��i�ȓ(��0�5&�Au�U�oP�pr��F����;Ţ=4�71e���ȓl?1Q���	wl��sKH2�̅�]�q�3�ͣn��D���H�S-���ȓM}ش�֦Ǜ;����W� ����ȓi��]����b�1t��_�h��
2��R���9�r<��e��A�N�ȓ;�H���P���K�0�0���Z �D�4������( ߘ(�ȓ4���6���0�^ �[&p�d`��4���'<l� "�$}�H��� D��@��'�N�ڢ��)5�Ԁ��$�&�� $ʵ8;��`��(8�vم��luC�%�%tt���H�#^��E��=���+C��k��D�!rP�8��S�? �¥��+#��#�*Ј[��0s"Ofĸ���=4��a('Ro�N�[V"O�l�hY=]�AP�I.�>�2"Ol��Ac��"B|�ۄ#�V����"Oz��FͲX����M9m����"O2�)��*~�@��!
������"O(	�a�-0��Y��˘򠱇"OdU!� _��P��v��k�"O\DX�l�9FH��qM�He�3"O��0wJ�qQސ0��UG4%�Q"O�DJ�LS:Y���3���{3n� A"Of���i�; +���vM��;N�{�"O��[WI�(*�>͢C&ޡ��P"O-Ire�	8q*�����t��"Ov\`�A�hWLٔ$�-r`(�"O^i��J�d��4&�ib�#"O� ��\1�Lʖ�5+[J�+�"O� ٗ+��t���Ё=D?��Q"O���G�F2���`k�\RVp;�"O�\�R�	+)N�2�ѡ�4�s�"O���C�`?p=���W�q�z��6"O��u�C$q؎!��ɤ[���7"O���v��z�N��K�6�x�#"O\q+�ܯ"�v�@uJ�8<ŦI�W"O��E@��F���	��dE��"O\�x$@#O� �ʴ�ͪ/�$,�A"OL��Q�
 ���E��%�
mu"O�YGX�_���#��&��AB"O�X�Ԉ��g8�"B�̬��hJ�"O��p�
;UzbTۢ@:K|����"O� �J�
8n Q���� �"Of���P9���8r-c�[u"O���s�#Y��	��lT5{��e"OKW��+r(0%�(i�� �a"O�M��M�m̚ы��>����"O옉��L֖DZahJ
U�(��"O�2ŏ��l���F^�Wz��"O�xqE��d5�ĳ�e�9[l��"OfQ���\�xe��6EDڬ�5"OP髁럯I?b\"R��*H���"O,<��-�;�iH��V��2�"Oz�u�9~���y��Y�BPqc"Oֽ�E��&k�Dwk�/oN!zc"O�]��bE,KƉ^3\��8"O� �@\#}}R`;`�?Ra8��"OVE�p���jM��ŋ1a����"O�1�!��sR!o#"�"�"O�91_"U4*�B�J�%iX5��"O�x�SNQ F��2��
g�Bx�"O�T8��\!��D)������`�$"OF-�D�@m3�I�!����Q�"O��)Y�?��֊̼5� ��w"O<bsNaV�)$ci���G�f�<Y׷}������ V�+�	�d�<�b�� E��J�+���[��F�<�Gk��nꁊq�ԇ*=���l�V�<� �C�R�n��FX�i��P	�/CL�<1$�W�4�I8d�#f�|r̘]�<��h �VDP�/���&�W�R�.]�ȓ�dx�@�;d���G�<w�����.�yr��qA�b�
3'*���Ź�y�oJ�[�,ag�Lg��Af��4��OE���R/=E�(x4��#�Ho%���ȓ^�����8�z�胊Gz�a�O ��<��� E@W�ɝm:q��*�-���"O�ꕂT��hS��K�|��#�"OX�$k� i�i_0pi@0)��D�d���'~� �S��_�N�R���?[�q�ȓ:I��`��G/����	ؑ%�n��O��(?O��p��Y�<�rO��?��y��^2sꀰ��)$��hO��ɏ�p��s��s�z	�s�3p�Zb�0���x��h)ã�)p~l 1&W�,B��>�AV$U�A=�Ց��0@��C�ɋDg����=��ak0�Uz�C�I����[B+�b��9��KG?�C�I"u����W�E5 �V Z�*�	x�C�3y6�t��h^��8�+5(P=j!�C䉭vJ8�7����^�q��̰w%(C䉍1sX  NM&^X����]��C�I�[��#b�^},�z����~C䉯_45(���7� P�@��T,�C�EWĝ�V�Z�_����M݅L��C�	-dI�W#W�W�ԕC�ܖl��C�	�(�a�����f!�b.���B��8���B5�	�N	�=ٕFȱ%M~B��T.�YãLBD��Ԭ]|B�	����%� \X�5qFhR?,%B�3W���hǲ$s�y��CF�J��C����!�g�$�$ ��C�Rx ����<���X�5�5�Rᙺ{��̋��E�<��fF�)8������o&�q�W�<a���A���OвM̈́�3o�|�<�!��p������s�|��
�A�<�RdǓE!�=�"d��M��e@�<郡��u�|���N��:�m~�<1LTIM ��O�n;�U���^X�l�O�@�4(I�R���k��
�xQ�"O����oB/xFxrƋ�#.�n��b"O� Yq"��W���鰤P�@�������=\O�0qC��$b��p��[�n| �
OF��A��n@c& ��^���f�y�/�"s pw�[�.x�҆�ݰ<���,6�+ǧV���)���T�0�!�d�DaTUH��f����t�Ӎh��IN?������$��9��Q+Cǒe��>C�	�J9�A��T[�8����x�d��'r�q��A����`��;:l�`�'� E���V�[?�8`,�V~��Q�'{�C�U?a�RxF*K,#�.��'�vHr���c��Ÿ���!*BJ��~�C
n��Ƭ�l5�j0M��O<�=�Op���0K�U`N����q.L���hO�\C��9):������D�$!�&"O�`�n��v}~)"a����R�"O����j�?.��8IZ�"���KU"O�-�d�R���N�-zZ���;!���,אpv�AaL)�ňƛ%�a��蟀RҨ�!�P�W)։ �u�0}��'�x[GF�Yb	���6������7�	���$U������^�ND�<3�B�ē�p>!u���p�X�r����y��Z�'sQ?�� D;+�P��$��NCF����,D�t�4BD�*�B$�����h��,D��fl�?4~ȕ�a��:$��ux�,0D��0�m��pL�3 �AS�qhR+D��C�(4�.){��_�B"6@�֊'D�R%��\�:9�4�!L(&��%$D��zSl�2~��l[N�!�G��>��d5�g�? VjS�7�	��B�%��"OX��d���n�8� ��1X4e�V"O���&Hԝ^z(ܘp��J[��h�"O��*�6��x���F�L�fx�����(O�|9�IrDG	<ie��I�>O�p��l =�Q� 1Qn��� ;QP��=������$D���1!�G�@���z�$�6�y�h��Od��K�,5'D���'�yrkF�	T0�5Y0��j���yrBU�^�\��3�D>#��P����yB�7wr5��.��+���Η0�y���Q��m���o�~�Q����y���H��t
Q^ItX��A��y� ޭYE��@��EQK��Ж���y��eXī��<G���6�[��y�+�5$����nŕl��	H�M��y�H��P\�QH2��Op��ȳo���yBd0�R%��%�@6�]��+��yrO�H�z��"G]����1�yB^7�����D�*�k���y���*쒽��݇�%;$*���y�'�l-\�#��"L��y�IH�N��࢈0���:B�Ҕ�y2*�?u��-R�/Ԯ,AR��V�y�&�cb���B�jt�4�э͞�y��@�<uŅ�s�d�B�HF��y"/.Hm�Q"rKq~.pˀeV��ybћ<��qc�
f{�{�,<�y"#�7mXL!���d:��p���y2GT�N�*�0@�R$	�`��G'�yB��&ZF�A �w��T�FM��y"Ej�r��F���i$c�ϵ�Py�NK�����V4fc5rbD�NX��Fy��׌�2@u&��e7b�� ���y`��-�n��f��mFr�����5�yҌ&4��D��̜m�������y"��++*�{� 3$���jD��O�=�O��(��`�.HxR*Y�v���'l����9�!�Y)f�f�$D������u0(�xA��*b3f��w(���0-�t��x����.�������O.�=E�T)��<�Xzȗ�$Ǵ� E�$��>aJ����Ê�2&�U�� �0ON4�d�/D��JGo���MHP��'PXT�Aց8ʓ�hO�ӭ \�-1ai
�W@�9���frC�I�~�B��)x��y��̏c�Nc�,F{������x�xq��g�7j��4S�� �yBń�B�
h���^�L\!���y�m�y�tA��TO]���ø�ybɐ�Q��CulŭH�,}��,��y� ��r����aE�9�J�\�y�צ��[GAUf�*�Q�E��ybČUTʜ�%��]άKU	��y�̈́�a���2��O�l%R�lɯ�y��Z$m��X����P��+A���yB���RT�)���r�,�rw)���yR) ���Af�z���&l��yb����%��ʍvh �
�P��y�J��H@�$aQXx��RkQ�yB�A�?�`�6��FpJ��ϵ�y�OL�|��J&-�$�d�$-]��y��ނj|ʝ3�Ȕ��20ɗHF0�y�
{�ک;0�OY9�9��#޴�y� )J�~b�JF�M�2��%I���y
� ���� ��m�ƥ�sXb�h"O�����_9Mր��R��� %"OK'�:�h��aP��-��"O-c`��w�0��;��Y��"O�$A��^�B����[�x��]��"O��c�iF fj�<#��w:�� "O�k��aM(}B�4v�AW"O�`�c&V�R��3#��K��D��"OT��l��}�´�`)�7H�"O, H�oț���EF�x�T"O��#����j�t1{4be�vi� "O� ���V���ن
�V�H��"Ojʕ���Z��dK�f���+�"O�{GB��z�h���F����9"O�r��̂qP8i����5ۘ�J"O@91�DfEh��r�*z�>�@�"O̀D���L1L�c��1YU"O����mժ��8�w�s�h�k�"O\����\�p8	�)S�:xC�"O�TX 6Y�>���H! a���"O"�J�F�	i�h02(W�Y24�d�'G*$ad˛+�]��)�0�a"�E.�$�ٴ�C%C� ��'6��u�.I���0��&e��P9�'�2���F �L��d#�H.��[�'���Q�_5�V��&ᛇAt�J�'h�����/ɴx��`�
�'c>�Paǿx�H1H��G+�)�'\z(�@%��.$���b��y����'�2��f䏁7�i�e�Ӷo���	�'�L���Ӎ�vmz� \�e�Ľ��'{���#�2��U�4,܆P�����'�t,���D�G�b!1�K
?e��|*�'2.��b��'A���CG��2X�@�r�'�P����";�ށ��j�]_�=��'�Ta��L֌d�`q���U�XeC�'5N��~��� /QG�괘�'�ePW��x�Zw'�B�Pś�'c$ԙGJ 	4J���ѭJ]��H�'�L�@ř}!�p�V�,t��:�'8��2�f�fU���e�3^���'0!)6"?�D	Jb��p�ƥ�
�'Ś��7�\!p��}�f`1�
�'�8�����|�0�Ⱥ:B����'�)��	S�*��)��m[�3���'�г��Y�bPz�3�&�8�0���gO�I�a���g�z���>��c! 	�wJ!�D��0 `�#6A;,�8�镈Z��3Ҹ�!����S�Odȭ� !�t�p�$R�1����
�'~��AC�&+0`%8W��<1�p���R0�2zd�%��~�?c�|� ���lɯ�zU� �{��HA))$����Lڸ	=fݨEkeֆ�'MYLϬ�����aǁE�,bB�(��B�d�F{b*ýEe�U(A�S$��N?9���̋�"4���D�1�ȸU?D���&c�+vr�O�'F<��a�`@k��ŬF�,$�d
��C��Mӂ�M{�|[�'L�8�0L���C�<1�\dM���iI���������7�ɖ#�01a ��5]�����hO�L�2�XL6$���aubDؒ"�'i��#S"V�ei<`���`$���fԨ2�<A��Q3����`�BH���x6��!a�\P�������/�	2#�L�iaL�9F�&5в��R�O�t�t,�[�iZ�B�6R��
�':6�:���r�RH���ܐ"���x��S�gDXr'�D�O��)n�h���V�$��] ��_/|�fIPTE)��|2a�	� X�uk	7n��(�MʥJ:�y�����X� تx�d��4~�^��mO)l��>y�	J2>p�!� Q�{�x$ar/�j�'N��s���fx� �A�n�� rD��R�,}1� ��K���~�qKxA>����;P,		��>��`�k�����*/V@�%�SH��M�ʁ+�!���Pu�� ;��\�T�]:��Rom>-λ�Г$A3Zְ�� �{����9&\Q��D<��1��	/�H<�����^� ��V��b)�cu��!�:�R�'��,#�H�'���;� �8���BY 㤨#ד ��{����-�Q�#ω\=�L�G���p� �)n�x��e�&zo�d��V�U�L��&jכX4Q���0�O��p2Y
Pd0q*9�I( 7��X%l�v��h��D�D�B�cHW��Q� GW�K��"��˒-�>���ؙH�l��T�K �p?�4iϨ4�aH�V�TR��-L��R��^2lJ���H�SSF��ĉ+?�M��)T�PZ����2C�`�b#b�(m�bSK�E(<�AY�
$�RBʁg��4���n. �+P <)#�X�JȂ[�-��?(����`���U��i!�䓟|�^x"�(4��!�'�@џs�锸�dȠC�]kM)���Q"�a���.?Y�@�m��|�{��صi�؊c�ͦNچt�@=V-��Hc����_�f�:E�
�j�{!B�>A#�*\L�6#��纍���,S<Z��R�D�i8xn9o�%�)� O��ҖF�h��K�m���� =#�s#�9I�&����K~%��bA�0���M:��D�փ;(�Cc�9H�.��� H�.�I��pۣʖ�^Q��R�Ŏ�
��~��B�:(��.�yM(��fl�M���@i�"�ة��D*l�4d�dJ��S���Y.�}D>����C�J���'`ze!�Ȉ1ي%i2���h$��� ��� �ِ#���1,�)odYY"
ҧM�2{��C��<³a�>
�>A�t̒2� ���/!>�yb��c����䖣O��C�֣�y2�ZoG`�tM�5.z��*�2d�����W H��8k�b� x�V	��a�PIz�ڌB^ݠG��Z���D�	`����WC��p�6�2�A`�N�� �$[���b���r��Q�ˉUF��R�n �0��n�0^���u�}5�E�׫;ca~Bk�����*̊���D~�r�B�BF(@H,�i��X!�DH��k֮A%z�zt$S!��!��Ňz�h�:t�|2�X1%���)L �@�i�f�0�O����1*�q� �
2��xc��2eE�vѨGn��`oҜ8�ē��g��4����4ѹ��.<O���eD(�~��gˍ*Y@�q�=OD��G�Mq���B��B� �����bC��:Tph��J� i�M�2���+��9#ċ^�F�(���oQ�񤛜_6X�I�l�Ec�8RZ�aʬ���DR�ʘ	��K"&D�)�LZY=J�y�MGf��d[�g���a�ܝ��_��B(z��A#>�a~���K�,�ũ��>���3%�-{'�l� ��3s���ۣJ<S���b%
�dKg�L?;���k���|(�'�%Z`�Z7?�]�VgQ�y��]bH���0�N�#��	#E&M�F���B��6L�2D�I�}>�"T�ђe�x��o�"I�������u�@��<��<I .ҍmh��N43%*�{���V=k�dsӢ�?P���0��kr�k074->��(��*� �9}�	��9�Hݳ�ʧҰ?�d� qi��cq'G�$�D��I)y\%�"�8|j0B."@�����/h��sQ���u7h�'��]iD$˛>�R�KT��D�Z��}�U�%�:�.�8GH�lL���i���{$�!��X�Ƭ�D$,�ŧ&k���9r�'l���K���!Zu�D���Ο'��d�6L_:IqO 4+�kۍn;P�XNW_E�\�v�Ojx��jĠt���j�%�5B���[m2F� ����XJ�p��h�����I�* �$�΄�m%3 2-�@
g�zRiL�r�pY��ɖ;�F��Y�%?D|7E�7?q�L�3	T-Q���p£�$rT`�s'�>�T�BuY'=Dxj�E��;x�h�]�zY�+$ �`�f�mP���DՆoV�5�'E�4S�|� ��ڱ'�(hK6n�
��T��׉VQ�[�+B7d�>��)��U�j�8�%�0&�*dcFn����0n��2��-z�<BA&QW[��=l@+��S�k�:�^�q4@ ���¡�1L�ᚱ�ĥ.�8��KD%:�PS�_,rX@�,S�/�@\A�CM�'1�}Zd*I*P�1��."���q��D���JU�P�7���z�k�c6�mBDJI+S�-)�ܯ!���QVc�Di�����O�^�Hs �)A����'~�pѹ�Ը�o��2��PTg	"X���ɍ�?��-`�K�Cx��h"%���ؤ٣�^5��)�wy���bg��v�ą��%�>-g�	�,c�X!,.�d��ƝJ"J�G$5ꡲ�,G�|�1�Ҡ&�Yb#+Y�z�`q���O@�S��9p��(  $ׁ25޵���$�����$94�� �sj2UYw��|�v���)��V)Obm�GN�o�!
�p>��	N�K^��ghءP8����̘͟��z��!ru�+�J��N��H�b, �	R94]'�P3t7�m�D)D�����'39�\�s�Z4[�ޙ�2��=e
Y
�cJ4<`�iӵO�*)�@ʧ+��O�����IL��V썓ؠe���'٦q�A˼jK``ѳmџGjPDɠ+�x����oǔ8��&���6M��-�,�E!��ꐥ���S�}פlF{�)%�Pu �@ĸa����$K4*��L� /�R���ti�8&��C���,f�!򄍃/ jMY!��)r*��ʖ&Y<U�0�"��4T�ׂ�,id����L�,&fYy�5�jޥ��ʒ�V(��b5���;���9�*+D��gC�3GN����=�teK ��|9�k�� [2������7 [���,�eE(�|��O�Rdjƶ[��q��]G��JE�'^F�K7�@>�^��g�h�? RȊ�5s�-�7�ӓ&Pz�H���.}��m[g��0|�(Qb%�	�p<��GX�=�<�b�h'n�*V�l�o�"!&j�-Hz�Y�M��u� E�F�d����tG��N\A�uh�%}�L=����u��e���0�4i�ˇv��iu@̆P�V�qg@PR�n���'��U�p@�鄛r%k����IU0�T�Q�p��5i�ST����-�9Z`ԁ#f,4��0�g�w���R�o���m��^�3Ϻc�L��Ӑ|��5�^9<�C���w4釭0?��.^.=�m��B!
 �����n��"�P�,�}jw�W�2~$ۢ�]�0��C��J��|bsA�1*U���U�N�=2�D���g�'[x@��k�$�=/,kg�ВY0�O([�_?�P��͒-R�PJ@B�2p���4+7�]�s��
��  �_9^�8Ad̢9�4� �O�mcԌF�%��h34�^ f�������A�v81r)M7@&�%0fo	>�QoZ&G��������yW���B.�98�]y�ܢuL��xr(>4n�akV-X�v�����#��g��ɜv?�����'�z���ˁ"���y�O`�`�*�@F�$*��_�?}��e�'G�0D��:p��j�$�<=��7�8tAq�S4��8�tÓ��9#o���$�(�(�!J14%ȉ�D�6Im����+G�>� 4�&=7�'�8�D�N�8:�P�d�;��J��EL�\��3O�����.�$��L��!B_�Y��J��'��2f�W
�̓�m	7Dc��p*٢e�6�!5�=Zۚl��ȈC��=J�Q�諕�	�Ec��@�w�@8�0�#*� �8��ɑFY
���'�����0?��CaԼGǜ|xUk��yp1۴zl,������zQ+@�έAl`��7fC�}��!�`ʗ��!�D��1B+��P�,K�.�H�w�/\O4���B	)]�)�C�R�TĘ����V�r��A�O<O"Bd��L��-��u�V����B4\��"JQM�'SZ���Y#�4�聪�L��k�{r΁�O��"	�[Ši�id�@W�҄$�D牃�����!�!_N@p���$o�b@�j�iL:��'o����ᄖ6�1�0�%*�J(��]/xPT���^bM�bME�+`���'�H���Ӕm#aͻV[�``e-�e��ԛ�L�/
$.�`�O����^LT:I?���"���j=��A���M�fAЎ+�bH��V��M�3,�00�ᅜ�N,���)���M�#^��8CC*Z.V*b��b;�
S�1�8�����	Sj6<ؑ�ŨKF�,��꘺u�d�D�O�c+�m�w�?9��+��N��H@F"{h~U�CC�t�H���g!�]��'6��c�,�q���>p���򯞳>)qOJu�7/Y�6d��G�H"J��S,Ux���1a.c�r�@���,a>��ƕ��	� ��R&��b�c��fRey�Ȟ�b�v��\�rp+b��ܴg�́Q���({^�q��@�a�[�)\�P�$�ڧ��#� ����2`�ҽ)E�i��03��gʠ!�w7ֽ�sKN���x`F
U��C�ݺ?��8�K��"iօ��
8�����]{ʔ �$ �2QCb��%�?_����w,HL oڬ]�l,��KT���/�,p�^�z���w���7,<n�v�ywh&"/l��`��$uT�&i�u��#?i!�]�'+^�s��<��$V�6�L�1���5#r���N)]Lv�#�.��gt5)���=�Ƹ��vݍ#��ĚXDĨ�!&ϸ2�b��B%_��P���A�T�.�ش����'��bC�M�(���� q�&arA��"7�d�4kT�*����Gi��I���q�b�79$\��bL̬~���d	��!&�d��,���7������ 0�i*Ui�1�U���=�� P���:e�Y�X��!0:H�کRd���ѡ�)��@bޙ��&X�$6�,��-MMn�dY��śhl�-["�-��h���"RH�3ړD|�0�E�_c�]�D��I�� ��0^?���5�ٔMO����N�F�8�%cϜZn�a�D$كM��04�N�S�b� d�6y�۠��r͜x@��Da�p�����ࢸ$b����k�+�*-AcDW�s��t��L�y�v��2��1Mb)bWo�%K�8�W���(�"=a#�סs��@�t�z�x��J�i�N���mI�c�fM`C˅��'n�x�@i��fޤ��So��H�R��P�O�RmH�M�Wp��CI[;��X�e�5Q
q�q%G�;����,�6fP� aS吇Q|��s	;��O�
�ÁN(2Y:WꋲxC �j %)C�$0�4BR'v��ӗ�V��)C�> ��ⓤq��$���~�.]�@����p"���b� p!��*��<�	̥gK4q�m�UF{�,Z�`�0
5h�;Jjp)��Y�ʮm�Q�#P����d��C����'c�(2�HϹNzXAqd)İQ��^1۰9��#�?��٣�E��Q�͛�o?џP�W�OFx�7�͆,(�����Ñ���4p��b�\��I(a

0Ȝ�.�uw��yD��b��M�OLE2���b0,�YC�R]5�H���H�v@]�@��a6 �q��\7� Xg�Ԥsoj�
�BS�q�h�M<N�|K�i�\x�W�!Z����)���y��)P�[��`��Dʩh�F��/5�X6-^�M�XU��	c����0O?7�x��2��++`�{��L�:�f��'�XU�@k�
ga�!͟�X�F�5&���ۗ�ü;���0���E}��^�e��!TL�L5,"<)���lc �Y� �.D8�2�Lڡ��ekP�ؚ4
2���	/X?�;�*�`l��B%nJ� ��B�	�l��R�$�*y����1��IBdB�ɗ%��kv�P6�zIB�+�}rB�I��|�93�U"*"~���62�NB�ɀE�i����F<��M[�.
B�ɹz�|�1#n�R��v�W+�$C�	�,��yC�+
��Y���Ֆ8�B�I �\ԘӤ�3>�e�P�O���B�)� `��2��1q�'�%dR��"OЭ�ԉP�aPRL�:'S���"O��k�	̃ dt�i"N� ��"O D� >����� E#�Ȼ"O����+��,���(�_.�@J%"OL��`o��5�B (%]�;
Ys"O��'��s�*�qD��:q�8�"O,=�G��U^�@��\�>y�)�"O���OB=G�4L����TW�ESb"O� #� �2Nތ�A�J�i+x�;�"O� ��I-�h�E�^
�sW"O�	3%�>d}�XC�d�o�(�"O�Xڷ�JE��c��B|}{�"O,��raW U�uIC�NR����"O�ia�l��C):�����)c�Z�"O�����E� ��9%a����0��"O�QoԻt�ȨRaJC>3�B�bG"Orp�4jK��$���ǢD�^�8w"OJ۳��(s2�� �̴S�Xe 3"O�p�EV|��]���k�䴈@"O�����Xu�p���ٺG�%9�"OZd�����-P/I�m�L$S"O�z�%��h��g�V.j\X�g"OXͨ�	�c(2��ժP���\ۃ"OT�pp�� ;t�0�՞{��:""Ol��Ɵ�{A>m��� ANH�q�"O��a�'k�����4'?����"OԤk1`��Px>CQ"�Z(Z��f"O��CV�2h��7�K�>  �X"O�QB"	#`��XP!�O?|���"O��`��_����"��/(�T��"O��j4��4m� ��
2sRx�"O�1"�Oܳ4���'��\	h)�"O�}��DA@�
�Q��Fe*�"OR��'C#j����X�7��+�"OU:����y����U�	���V"O*X�ָ4��1�T����$�6"O,������`�+ �P�L�h��"O���Fĭ,bd�Nʵ��8�C"O��ɐ��
z��0���<�p#u"O^-c���!��4����>(�8}�!�D
�a^~M�� 4 Ҷ)KX�!�>�$T�dD�-�"��"G��!��Z�c ���Ϗ�iC<��X�f�!���Yx��	�*��㐈�U�!�$̇G��u��#6�i�(���!��-I�r	b����d:�=�"'ɩq�!�dK�.��[Ѧ�?�y�G��%n�!���I�R����2D��G���џ�Cq'y��>yJPcC�A~f(�5oP�,�n( 3k6D��� .J�HS�L���	E�l�S�>�"Ҏb�F$�G�x��)�6Fl�1aDysڱU�H�d�!�ȔzS
xQ0�قp
���ݒ&G��,� ��:'I����'����kZ\���T�0{
�+F�%�t�V�v^iH�{��YN;=(^�`'�%Ra����8�)xj�)&��)�F����hO��̎x��JI6~��gب�A���s��U"�B��L�����Lp2'��$5�9jq�E5=���o��O�x30ć�B&ڐ��G�5�ȟ�)#Ԩ��i@0�vt�a)̥�y��+a�$3%��7	���D'
�"���n�e�L*qF@7��hi"ԟў�
��J��H9B"_�$PEC)�O�� ���AH1y��� ��P(bm��uJQ�bH؏g�v�@���p?q0� Ӝ�������k��Lp�bΚ�1f@��0+�{�#ԯ�Q��x�@a��v��	b�`�(H�\t��"O� ���a�=/��,U	,�޼�'l�r�n��k�H��R*�
}��>�ɕH��-2���h�X�"���26�����S���kVeүe�p%(����OC*���R�Tz�ɫP�W�#�fu��$C	M-4�1u��>	�t-D}��؀��=�_��9�����O4��Ͱ6I[���&,0AK�C��>� c`�ļyRP�g�M�liDB�mT��W%��p?q��29����f�O��͸Fh��h�9��n�k���d�Y�h�v�+&߱>����aFڹL������0m�H=���oS6 l�!A��q�<QG	5�,�7e��O��SQ��}��(C�ˠx[�ب�@�6��;$7ܤ���"90-c ����~���p@Z 
�mX-x���T���p=f�^(g(�+$�S(����!�#JD%C�߂{BR�wB��f�$�+b�D�#����q�\���,"�e	���1�эoM�-X��
r
��=y���8� ,��xP3 B�N�+@��1��qu��4V ���_�v��DK�ON�R�`)hC�'����lͿ���y ��:BBE��a\�n��ȃ���l���7?���f=���Ap��պUmn�Y�0NS�A=�S����L���,D���Lֹ������Pl �a@.�r�k�M�?"�ԑ2E&� �м�R�8��{Rk\+Wc���O0t� ��+D��!��N�>�B�K��'�"�+Ǝ7W��� ç�B\� b�1 ��D�N�(%<�� ��	+@,{)��;�d�j�C�	ґ�(��"��j��)5璷&9<�3:�ɓ��=9��P�~�h[ �*>���1i_�P��Kq��:0�
�RC an� �R\Ɇ�#s� �O ɑ�K�.}t�@tNR�]j ��P�Оl�:Ԫw�V�C�:��U�ѹ��kC/~|�XTޟ�E��w��e2燐rt��Fk
 e����'��ddI;��/:�,��l	�|N-RB��A1�ݚGC�ÈLC0G��'*��Qdcެx5��'�~� 1���%	��05�5!��Vn��L��LaF��e+�IA ���[���&tO�U�
8* [8,PmpO�&3�������*1�R'ʇ߸�Ӂ�0�qOT�� �
R�t,X�i�=^ �6��똵0�� p7���t�D��]�6�0���QO��e�@�}OP����
�f��W��[ ���[�>�� �G�y�,��灲~KT�O�,杆J��m����/�X}����kD>B��b�Xvn�	t�E���ѬB�t���a��*�>V �Rt*a�ՓQ�85-ʡ*�|r�H�2�����6L~�HDAR��<���6N{� �ᓇI8v��TJ%<=�	a��(BBzl£�/qJ�h�#�ٓ0`�z�DG'>��y 	�WOr�� CN�9��vj]��ēp
�)�;3��"
�vz���'�P�c�,�+�")�҂ՠ<�\i��G�4z��i)�l24����&�-�r̘@g����!�v�+~f����{DR�I�h�|��'F߯�z�̧��5�(v��T�GR���o,��d� C7��G"$؉�5[ AҤ�[u�����q�"]ZD�@�-=R(�D��ޜ!#ȡɅd��Gݺ�'�d��A���q��!Xy�XK`�<}��T�B��4��O*��q�ʏ�l0�E'�6��Ycem x�D�@�_�(0hЪŎ]��xrg��DX����\��I�P���p��8/E( Ҁ�B�.݀8�'��m��x<P��D��RU�8P ��$I���hK�r��Q�$\�J����:�3U��:"K��$	�L�x�f�]�zX��'d��t�d�BjJ�i_�9�pg	|I䥠�L)��|�v��{\�)��s�H���oP�!���ɭ���2��K�ޜʲM"�Ofu�.VN[�X��'��Q$�"//d"�'H�$ؖi�4"5 f8�bb�v�\0R�X$L* u��@��( z9Z0�	��'��v�	�Rv�{!<���Q�'M�|��K��}����N�M�6.�	Yl��R;���	@g�jI�����.�D)���*�Z�	��9k�@�bM8:���@�I�f�@��
\`eN�<a4��T	�V�X	P@�R��#6c�<M�t�" � 
^Ta�nʾe?���"�.����&�XI�#L��}2,�Xhxb.�=	O�`�D!�����u�����H5VNR�0@Ϡ9��A���>D�|#��� ����p���'|r�����%h��7���Y�ў�韂p���i��^���e�1����A74$&5sE��0-cB��h2x4T�B�S\6�b�� ��(�ga#���/��`]���SK���<�I�[���P��=�.����1��%�	cZ���#����,�0P>�eL��1���t��u��$Y��7D�xd�$�b`�P��9���.m��%j�NS�R0�t֏jixQY�	�!1� 5��a�b���F��f��.�+�*e�N K�Fa�D��"m�}b	�dX�Jۤtޒ��瀁�K�" Ce^7J��awجz
ԋdk2ES�e��'rӈ��Wትpۼ5�0	ʃ� }��h�,`�2�=�$��k�2p����O�4��X�N���
q\�T�DS*[8	��B+� ���*C0����'����)�39��Yjt�+	�8�/�.%۳
]&A(ƌ��/Z	6������. ���ϞS�ЈĆF�\���2 	 �E�[{,HR���ze���Ѓ�5T܈�'¦�4�Ç��J�4c6�ɁO����!�W�ӥ���%4�D-�4�
9�dD����W'�n�T�
Q zLP�.�qt�z��͉D�
mce�.1b�ܒ��O��hO�a[�<F�J=I�M*����3k�76$u�w� c���0m��"�:D�� H�Ѧ�ͶJ��3CD�uw,��ǫ�l��`�D�ڹ0C���'=y�Z���)��H��z�%i�
����4Ϟi@/�W��C�	5F� YP2�V��p��AɺR�|m��$�ni����r��c�lv�ݛT��9X�f���<�dR�X��0t� T���k�b@���z"hU1>�ִ(0���K1j%x�GH��@���L�g(v��a.�2$Gn ��M�\��p0�����dL96&��+شK.���O�1O*��b��
L�Ȉ[�ΰ��i��8)+����;2!�12K�.PG�4���J�,��U�Н�PxBc���A"w+E�#��$�E5K<�ȉ�Z&v�^򌍰F�Lx�Í�
��e���|4.Ŵ�y�KG�b�4�!"�ӊ&�$�3DC�3��xB��x"V\{�aB^� ���&k�$�W�Ŵ*�,�����P�
f���"70��яn�IV������2j�	[fHʷ2����D��1m�%;��44�� � �� ua�9ZtO�HsV� $�C���X B����ćT<I"p ԎHA�'���q��9s��pբZ�\hX��N>a�b�!XcB��/��"V@����Q �1�uft���CC�F�<]v��B��9-y�l���Zw�~8��E7�O~F�رea( �7#�����Ff�!S�чQ\cR��^�`,m2e�ºs�'�-�yw��Vd"ͨ2�.%D3C+_���x�_Q�<� �E^ F���#E2 ��pL�Y�ɑfH
�[P�Y�-��sRr�y�Or�����^r�h� 蜫94�����'s�|�])<9���C�.>�v�"s�D�/�V@���-�PR�l/1�^���ķx����a���~���$K�z�
5CAW�q���⑷(G�'p��1���5-J�����2�x=p�M�g$ E�4O��:)�$�!'��5wX\Jd��NFz���' ̅���%#N�B�݆OP<)�q��
fvmj��U+G��q��R�ҹ`��%X�zdK�NP:9��w�|��aM�D(��;����I{	�';e��E<��DXFW1X���C��XV�p�۴	���"f@�6_�p4��+˞)u$�� J�f�p��o�㦕A̘����.�C�!\O8�;2%�;m�N�)�"E�3���x��o��\�`,�]F�׭N`�L�f���<���E�u���0�T^�'�"Ap�dQ�BKEy��I $̞q��{Ҥ��e�.����C�!��	j�Ȋ;Bl��<Q�b_�0�$=2pDŀY�5Ѣ�ٷc'�P�H�DV���?�hK���[��.tFÆ�O,:����)�  P9���-8���.Js�pQ�7�yGdSi/z�0���)D[���g�WE�I�S��8IKNs��g�u��"F,�G�YR��:�r	g��"f�jp`4�iIb(���$�>�!4��Φ6��~�i�c��Of �hb �8�ژqW+�n�@!�G�ŋ$��#���-6q�Q[5��"�,�H�<LȀțg ���p5�Y��>�T,�?~	�a9��J�Pl�i���KŖ��� ���,��(ԋDlA|/npCd�T�Xe��6��'�
�0bZ�g����ڣ�t((p(�+�]YF�i�dP�٫z���1q�\�3z`�r��sՊ���Y��ƙÇ�+�MsP.�0S�n-SK~n%|��r�^<�<�;2oO5@Pa��F)��јs�>'�d|���ŗ"bā�4w�E��D)�j�̻k*�%�c��d��d�2J\�92b��Ƣ�28��xƊ$+��!г�hF{��y���:��N;N�T���^��%�Gݯp.�6-AH��\� �7����.Dq�<�i
��u7��>(����W&@xu���� �����Щo�ti
���S�n)���[�HV�f�y�ٓ9��:f���hU;O�`���o#d���A��5�uW�Y#eL��c��ٮ(Cd��X�Xft-C.�:��*� �j�n�`5m��B%M-Ck��z���Sj�<8�m	���w�6ͤ02It0p2���v�u8�Z�'������#d�x�A�0ƶ r	+��'p*���FJ V\��GC�SN�()Ag9	d�xy�e�/x*A�J4�� ��%]J䲷BPK�,9�w��=� ğd����L5Y2m"��]�B�)p�Kw�҈(cŒ������I0}S�}��ڏ<��x`�M$0[�0��5~e���s�e7�XRe��}Q�e����;��L8���%3[�8��4�. Ђ�Ä|F 7di^F-(c��.�8"?Qp*�8%�p�Zcj��B�G/N��I�`�!��KG/0%dԪ �!�-C�뉂C�v�r�bG.L��i�`��'�� (t���3#l��Bf�3}��d�p���'�< �'����t;�*Ή6q\�p� ���ޜ�D��Qک�Q�с]����P�͉O8.UA��)8 1����
�҄��S����?	 gY�M���E���3E&D���w���aZ�ZO^tb�æ8(B�1P��9J�����1F L�SݼCe���[S8H��O_+bx�����P1���%��H���z6�;�Q�g�'Ui����~6��u�A&-��'E7�JLY�R�Y�X8bϼ���mD�v$ͱ��� "��ǥѴ�|���3�R�#bJ�4�ttB�V�{LrQ(�	(�Xꡍ�(X��A���K�Q!���w.�b���K��ӵ	��:U"��hJ�U�:M�Xw�@��w9E���t��E��h�
�Xc�#�8�0R+��(Ov+ԅ�k��h	��!�>� rk��AZ������^|LI���Hv��6�J?�����+/����I�}�Y�����z-�扦LLhA �Ǯ�jMɖKe��0��		�"�����-(���s�ؤC��\%#�J���c
 *Yzu��z}r��� @ I�*���I+h}R��)��='�	`p��/3�*��'�&�)a���z��G�52�ˍ�?+F�@��G�Z�`C�)�&���)�	E������T�-s@� �LaCg�;w!�D�}�R��A�ęt��D�F��]4!�DV%rP-�檌�M��J"/^l?!����%�DӰ���oR-.!�� ~ z��C.M��K!
�6B�]�"O�x2�̊�rƌ�� �[1cJ��"ON����G%���PЍ1�\̱�"OȈ3R���&@�ł:�N��"O��C��ϳK� ��e��7-�`as�"O�=jЎ	4`��9���'�l�[C"O�A�3��4�:�S 
1f��PA�"O\ �g��n��$I�C�3�(|��"O<�p҂ޱ!�<�����4����"O���@�m��}w�E�F�&H��"O��[7��>���BR��@1s"OftB���Y�Z\�s�%A�|��"O��sp�U�}�
��&#C9#N� "O����k��h�Q���=C���"O�����(�1�/od���3D�Da��B�X�����:Ae�h:�.D�d� ��F;b�C�o� Y螸Y�,D��Yv.�x���"�CI�`���@,D�H�n��"c�9��5��F*D���`�PL�����_%� u���<D���nϣU���+�DW�S� q�#.D�T��mڙd���8E앢B�h���*D�(У&��/,X9��cօd��@��&D�<9G���2��Y��ˁd�ʄ��$D��S!�\�X�$�1����̀��%D�|�� C_�������`��1J!D�h��M���B��̷� D�o0D�ЃV�'?n��Cm�U����%D�LQ�D:CL�CSE9��YSg�!LOҝ�ҁD�K!�K) ��xx��J�Z�Pa�[Cp(�'4��S��$%V�d�	�ύ� �P��&)�+ASb�O̥��mx�O�Z����C�,qE��ŉ�n����5}B�˓/�dy��5�Y?�'��y���}L&�E���=z�E�'���k"a/�)�'*�0�Y��>(�����]���lZ2
��O>		�'&�F,���w�V˵%ܠfe��h�M�ryBw�1#��'�x�	�*Dd���D8C�t���\�x���Ӻ:tk�ꦕ��:�N��8~��p�^'F��� >e�B�a��xr�0.k��S��R>�y���fK
������EZ�~����'S��gǟ��D^z�O��C�k(1vё!eU�N3�S����T�S�Ȱ�������>
0�M1_�D�A��e�JxpQ�  ���<yA�O,��h��E9vbUؠ� �.!����	v����M�.mZ��H�������<�M�y�
p����~ʓi�Y#�'�.��	�',9������=^��d�`"�`H"��	>?ٺ���M�(O��7�S�&����q͝>?�Α���>&��cROJ*�?���<���!�Ƞ�f��#3�r�(Ӧ�@="�������	w�S����N��0�	�^�����iU3!9�L<���"���G�V�1CT��L$P��5�V�����O�`*��'���՟�;��� �,|~��2$��ELn{6j��~��ԡ�7�&�T?)jJ~�s L����`���<��� ME�=�`2�(�vݛ�'�<��|�>��4gܐ5@�y�/�,4D R%_�Lr�	Q۴>��	���x����3j�8��%�'a�-�2��a�,�:�O��P�ըN��"��I�#�ziI�'�Dq�f�9LM�1�kKz�O��1@�6nҴ���'�����BH�cۆm�6m�Y���rƴ�?�'m��U*Zp�d��1
?�b�'�΄���
se��O�
.�p$�
�'��샵y��$D�w�BXH�L:�y�%ê6	(L3ce���`C7�G��y2�ΟV���ueA�)��)�	8�y"��Q�v�@�	*MK�A�G'6�y�̓)g0�8���ޤ/�]�6H���y�V B�Ό�S�	$lȩ0�K9�y�a�w���
��L�dM�Ա��@��ybB��&p;�"��'Q���Ι �y�)��w_d5
���,�����!C��y
� ���+�~N��B]�,�ȗ"O���v`W0 Z�āV�,H3�"O �
W#�<nDD�#�K�8팥s�"O=b���M�4u�T��|����"O*�`��P:sl�Y�'I�"T.\�w"Op=��j�2K�I����#.�:�v"O�,��F:P�uf�	C�t�J�"O�i�
�EQ�`��#���q"O�5q�١d�I�3� l�By�"Ov�Y` Z����é)/���{b"O���2�т2�Vpj��\�x��6"O�)���O�~�q�)	!s���"O�1���TrY:��Ǚp* s�"Ov��Q*�d@���n`���B"O����/FFS���R�!H�i)�"O��tǌg��rF�%eX)G"O<Z�+�_.2�����aF8�H2"O̱�f���pjR�y6�7TRHx1C"OTӬC���r.�G�\i1�"Oą���C����/X�$o��"O� R%�����.�:x<����'; ���M�HER�`��I���R�'���4eQ%hyj��I�B�x��
�'p�I�r����I��J�A�h��'�J8�H�}\���3藘;kx	�'�h�$�1#�i��<���^�@��T�8[
9�`,��A�Ꙇ��6��эN*H�����C�ˍ0�'\����+^70�����L��'L����X+w�!s�/Ǿ	a��'�8D�E�V/��}1To�;Q�(q�'�h�{F���@�Z��B*'`L�
�'x��).U�>-��a�%|�M��'��H�J�7�X-+A����q@�'�h�@'�21�֡;���*$��(�'�T4�}ï�'��zy��1�'$r�qR�k�؝۶��|�E�\�<�oD6|�yذ�D�X��<�� �T�<I���&^�����C+|	Nݚ#`�L�<1��S� ^�=�f��>��"6/YK�<��?]�&�s΋�;B(�  \�<�s�]9'6����Z.J�4�
a�<AS�!佚D��>�"U�6ȕZ�<�&��9y\l�ET"!c�kV�<��Lߢ#�t<+��(h��U�O�<�eء����ǟ�	 Sd�L�<Yҁ��ZH�=>
�
;1rv܆���A��`R�IWNp�b��72^��ȓL1�jB⋻8k�0 կ�,^�D��|�p�ڡ���g� ��� � A2i��bD�s�!�/#$ӣ���60P��n*1"௘�T�S� ��U�ȓ<h�F����8Qj$<_^��ȓn�qQ�a��:��#��O6P1:��8�����S�t��6�X-�ȓ�a#���?>\�!��j��|s�Յ�K�Y96��ur�]9$�_�4����+S�c�͑*�� �v#�5SR���ȓT|$=�-D����C'S�= H�ȓ2�6����|
� �A��]3����F�Zܻ��S����� f���ȓoj@i	��ղt-Xtj1KD>)j����I�d�c��/X}�u�F	Z8P�0,�ȓ)��R��7r�����M�=/h&���S�? ��Z4� �9�8dh�� �>G����"Ov� aۮtK�X�S���2�Pu��"O`	e(��C�$PǦA��bY!P"O��;l��$�B{�Q�"Op��҆S1����V�d��,�"Od��M�5�� �ʊ��L��"O�����+2h�Q�I���D�{�"O��j'�@�_gve�P��\㨵��"O��XrH�,Q�t9AF� ���"O"��!ܕx6Y:E��[@���"O�d�e��]l�p����2X��c"O"�2q��>@�r���#C�P�@�R"O��#���|�V�����H�p�"O�,�G�<(k^���!дF� 1��"Ot9�%m��2V�R�/�6Y��˴"O�0�u �-{r6�E%A�`�ĭ0�"O``(ǁ�=�PȑW#̣n'
`;�"OJ�zq�0\w����j��2�"O�M�眭t����%�R:�`Ը�"O��{�IĉA���� �b�,���"O�0!NJ��Ι!��:m�ry
u"O�C�C�H����*�^��,��"OE(����k�� �Q
|��@��"O�P)��R���(@k�44�N	�"OE���A$6<�|c�<x��q�"On�H_G�x#���"��Hc�"O����צ+Ԓ�+�̄9 �F �4"O�)�D�E�uJ����&�I e0D����F�*�N���I�}�
�)B�9D�t� k"6�!�L�(u��8S�,D� ��I)gqDC�&_�<�ҼQtE)D�xpE�ڊ0'v�ǎB�`Z���(D�4�pڒ(Mx�3���6^�����H9D� ;#���h�Ze�ǘA��y�8D��GY���Q1�k�|5x0#D��x�BE># Z���N�]�"X�'"D�(���7�Z-�W�'7����!D�������|$Q��;�$���?D�䫥��"1�¤A��^��Eh)D��˕��#�2t���H�,؈t �!#D���j�/+����a vL�,D�����V<�-z���-V�D�;u*D����H�	�hA���"�J`�A)D�ػ��D��B̪U�.|�1�(D�t5`T�k�^�;�IբC[��F"D���t�G2)�0UB��S�t~�A�ש4D�L�i���l�* �Q�/�A	�*4D�8D	�F�͒'�N�hH�ј��=D����T�h� ��̖P�e�6D���@���|�xE9�ω[���s&/4D�(KP�ΧZ���se�̫;^FY�1D��k2�'F���Db#N�r�4D���,�$����E

�gA�:c�0D�Hp�Ŗ!q��3�-H��� ��/D� DO�[�U �#		qf����8D�d:�!P�y�9`hǛM�2u�� 7D� ����o�x�h�Ǌ��@�i5D�`"��X*��ct��.�¼���&D��z#(�|xQ��ퟕ���eJ7D������7R��)b�]7x��芇�(D��q�JU�!꜋�P%z����&D�Ȩ���Kݘ[W��dLH�is�%D��:���rZdXI���\~ �*7�"D�\����D���iMY,Gk���'h4D�� zRbH��[�ЌQ���	=�h�J0"OEʕe�LY)��	3���A"O��"��7Hc +6�r���"O���F1y��+Q�N<]R\ "O�e�� Y�\G��cf#A�x��A"O�ٸ%L3?�q�"]�@���Z�"O�]ڢ)֢q�E�������5"O^u�2b�
!*�`s4�iwDQ g"O��0P'�8���Å+%��`"O�dk�aE#2�>I*�!�/�詀1"Ov�2D%WL���XF�=n�xr "O<�qp�W�m`'K�0l0=��"O�+����d�N���:�O�*3�!��4|���L�v���$�!�!�D�h��L��V��8%�0�!��:K�ԡPeV�%�f�	���!��5px���]���t-��Z�!�$����D�F$<�D=���w�!򄒦i
����_#��Smҷ_�!�[sz�Eb��]�h>�A��I7R2!���9	��,QS�+�|��Mh�!���0��t�vQ� �@�[Ȝ)v�!�Q)L�>�ҴݺQ���W�	;�!��#)�L��HA-jf�*6�]
tb!�F�W>� �!��tƊ���!���4r i��S�,J�� "}�!��L$>��6��2m����-m�!�$N57�5�e@Q�'�"��DhW�p�!�΀�F1�����P���W�Z�!�K�BI�� l�0)�^9�!�M�)�.���ʤAb"��ċ�4H !�)��S��&&I�5ȁ*\�s�!��&�b �2DP4	���3#�!�F�w�&lAp��T�F�c���V�!��^%t�D�� �Xb6<˓MM�r�!�$������Stl��L�h�!��ę>�q�)I1*��Tl{4!�d� �z��sI�zi�Q�bk��{!�$
9a��Bԩ\�=[l������=�!��K�(�� �F�)N���r#Q�_�!�EΚ<�*��)�k!�QxW!�P)Y�`f��kRY�pǀ�-2!��#�u`ch�q�����X/0+!�D[����P�Ƌ���`C%��1!���/E%P=����e�l���d�?�!򄕒V���r҃�
S�ܤX��=~�!��@*ĀR@H�,�8	�v����!�/��4ʶό R�:}�FI��9�!�$�	W�Z��C"A)'hx��V�B}!�$��(Uʭ�ah .|h���f�V
!�ɧB��� Gd��`eeh�!��}P��kј&�hq�F�R��!�d-t�|Q� B��\�~H3%�G#�!�$L�{R�h;�	��[��x2����}�!��I'I� ���\�{����$�^�!�D�<�2�z���u�LeH�d���!�D��} Z���EP~����E�YP�!�䎺'�`
`e�[��-S �A�_7!�dL�<G �  ��     	  �"  &-  w7  	B  �M  =Y  jd  �o  �z  K�  ʋ  �  ��  ��  U�  ��  ۿ  #�  {�  ��  .�  p�  ��  ��  :�  ~�  ��   E � �  O$ �* F1 8 Q> &E �K dR 9[ e �k t /} l� �� <� |� ��  `� u�	����ZvIC�'ln\�0BJz+<�D��g�2T����OĴq�g (�?Y6�S��?� ��g+D�[��L Ln�2�IV�2(���l��US�@H�"�`qIfk�'�� qPf�	�jz�	�*E2q�c�L-,h|�Js
�=)�\��v�ں'}���7J�.[z8p*3oӲw���0��Tk��#����T72+4J��C�#DL� f��-%��a0EO�O����Q��$�#��Фy��n� c�v����������ɥt����Q��l�q�)׊gڸh,Y�ȩx%�R̦q�Iߟ����?���aw������X�)dƘ\S@R*+�U������A����	�N��6�T�'�<K>`=|I��菗4-�4��
������4�yb��d�A�G�i��Ov �5�Z�\��I�cF��R�z&��U>8��y��d���dSUA�a[�牃B{|5�׈�!h|yѲH޽�H�$Ӧ�I�� ��ɟ�S�h�O��n�/q����[-#Dĩ�BT��bu�xnZ��M{վi���wӴe��Ѧ�z��/c�H)�e�0H��$��M�"a:*M�7���M��|@�(&���?1%+��|�����O��VÄ`'d )fR4�׻xI�Q�����$$Ϯ3�����414��d��i��|JTJM��M��%OU,Uyv$��	���+��ʙ�M��jU�rπQ�0�Q8QD~Xy_�6mUF՜��$Kb�tm��MK�����g�� �Pc���x9��P+G<='�Q���i��7-�Φ	�E,�(@��?o� ��놖;��m�T�ty�6�ߔ,�԰Sݨ^�J���@���M۴�iM�6�/���+T��|��e� ��[��]����%��!\�j�bbϽ0��6-;�tqP�L�������ҕu�n�$%�Ɉ�冕�'>��5H�aLj��X�7���4c�O����OD��韸yzBϞA��e�OX��c`
:SZ	Q1� )��=zU�>��?��ڏq6�	��,�IT�
�
I8���x��y�gH�axbm��I\� �����
cl�9f-�G��"�,[2m��a���:�D�ó�9���r��J�]�t1���M�Z��x����&KxM#�hZ1�<�%/�O���OޓO���O����O4��57і&�QiJՓ'aɆU ��d�զ�h���;`64[

JW��a� G#�M�����fۅ3S�7�OD�����?A	nd윫T�ݒj�E�!�ʖ�?��BW�ࢦ�	�F���Si�V��W�,) ��p`��4'��������j��XR��\1�騑bK=F{��w����#i���p�a:��%@�.�����l���6Mv�O���Gdjd�өj2��s©�!j�"�$8��
n4�;$��QA�<�`
ծ]��%0��x�TmZ��M���|��v<O�B�¯tV��+S�	�HQ��'l�\�\�#�韴���l��ay���mIb���O��Bt�"h �,��6-׎u� A(`D�|:��d�'x��H��֘#��`
�aǗ~��ݫm��6ì8��ͧG{6�ؔ�)@|�	w�:�;�a�В�`]�tWHT�Vim���'������"ȟ�'�T�Fb�zj��V�W�>Ap�%�'6�W�L�	\�g�$Z9uvV��R��>��mP�#==]�'�Z6�ᦝ$����?��'@
���w���;0銞y$����P����?����D�|O-6TK6�K��T��ԙpϖ��Q��0sv�0�U�Y}J9x��'7^��歓�dQ��
��.v���8Q(�7|�ҹ0uc��dܠLK�oF�$�џ�R�b�pdL=!!��j�����i�#�����Ҧ�R���6�	J��hR�=(4u��BM�}i.���ɟ���t�'�1O�Y&�ZD���ݒ.����|b�~� l�[y� �$����y W�}�y��52`\��/2�?�)O��d�On�S��ʀe<M

�ڦ������$e)Eo��nŔ%�5Oi�ة�0CD������K"�q���_0�iq	
�r����@<t�.�E2��%�?���ihV7��O$R�nT�t�,����T��8c��<���?)��0|�ta �������R����r��hO���ئ����9.`jPۖ����L�7M���M,O�8��d��f�|�$�<���f��f�'��aA�/�h(l��!�$/��T�$�'�2 -u{&�j�jx֛����	�Ҥ�9Y��m��dI�O����e�Ah�D@
I�LU�2�֗d�^�$��]OJ���*�l�qf��n�!D�%͹�C�	$��p��s��O�lZ��ħ��O��|�T�S	fH�Sa[�Yu��hK>����䓛?����$�=ܵ�h��A �5 �Y�<�a��ڟ�����M;��B����'I��	D��$T'�YCŌ�=��� y��d�O���M%`~,����O����O��Dk�Y���T1�H�b�-���S����f�ʦ�����5J&ٗO����#T��0Q��7� !��9갶��+�.
��@\��gF�i���#<b���')7@r]8��;q��9I��m_���[3 Ӕ���4;���
캝�Is��h���P`֣B
Z�0�ɧY�4�&�^ʟ��	럠��џ���Oɛ�ǐ	�th��ǚ�T0�����'8b,d�`EnZ͟�Jݴ�?�����+��Y��ޓ0��1�U�D�2B�I"k��.�<zpM�O\��O6���Ӻ��?�O׀h�K�*#�r��u��*4b�BR�y�(Jq-�n	*�q`�
�#?9���m���Z#K�w
�<��,�M�f ��폳�^9 �&ț0��A���,m���Vl��^ �4ࢨ֎^|\P؅��OR�,��O�A)V�Ҹ9��Z��[�jXI��"O<C�-Cv1z�C���+��|�t�.�$�<�ኌo����?�ࢦ�@�m��H�y�P�"�OX��?������t�=9�f�;;8�䤇�� �q"��HM������W㊡�1��>�^�A���$X��"�'c�D!�R��";�lq: d
vZY�%��Dr(!౨Z=:+8m�7qVF(%�d(�@�O�%m�����.v�<����g~����`W.Zm�'gџp�'�k�FH*�R����05�z���'I�\��G{�O5�6-Q�^(<��-	5z��5[DeZ�0��Un���$�޴~^����?��?���k�0���� �&�֞O�6�����M�U���?y��΃[�V�����i�@6�7���Ѡ
�
X��s�Ӳh�%J0�*Cn��t�؅��O�܁�`Q#��1cW��惡�2N\;�"4�� �9L�� �S�g���k5��qQ��*`СX���2ᢰ�I� G��?O�%�5�G�8���E�R
o��)Q7"Ov�E��u�Tʢ*��c����	�ы����HrE�ζ��;��7]p�QoZݟ��'���p�Ox��'�2X��^'���a^�,<�@��"r�l1!��$-{�a�C��|��|J0eǚ#���I��7'Y�f�
$e�<}�၏�GS6����#@G���3#�4�p�O�ܙPp�B��yGE�D�\���
z8d(�%.U�BV�M�<�C��t��f�L>Id�WC@�|xQ��.�!��J��y���[)��e �?���xN�7�?��.����ߟt�'j	��KM�7uHS�gW7��1���AR��S�'s"�'��cm����؟��' ��]�]���·e��`*�����X��9;�,ѵL7$!1��C'+x���S��ԇl5���K�qW�1r�O=g�x@	��P���y��:� Ez���!Lέ�`l@�� L�!B!̀#_���c�K�c)/�r���O��=�����=bR�X&�T7t~��g�	4.�{b�dR�t�u��:vt�A���5=��'�p6-�Ot˓R���C��i���'�DQ�S�-�2��#�C�S�bu{�'�-�?^R�'��)�6;��7	��T�`A�e�Y1j ���C�ρig��@�'^�D�� �bH���O��Z���.����T!݌w�^T T�Л�(�� �Ç͒�FĲ$d�D~2�?���|r'L�i���BX���:�N��y�-ڥ_�0AP�A�OSE�
��'�ў�Ӌ�y�$7h����0쟡n�(��ĭ]s�ɀ&�����4�?)������X���$�	|rY*�U�_�0��R �
_����Ox���N%1���J���|ϟ��c��Ő}�6(2�"�4jL	%�� IGoH+H
 1��'A%�)E��S<H��$MZ�xdx1�B�����Z�8���'��>����O��s��%1�H|�2I��
|>���r���(���~ K�JE"�yG{��'�t#=iq+F�����&�b��Pzw����&�'���'� ]3�
Z?R�'��'7��Ʀ�b�FM 9���id���L��ӱ��5Q�Yش���V��n�g̓lhD���H%5�j$�%�Ϋ=�����d.�b�c��i�� v�W���Ϙ'�vI�Q$x1�Xl��"������<-��'�2�d��E�l%�!�x�f<�bS�hENB�	�:G
M3-F�J�b�SF��p��d�O��Gz�O0bP�Hc�+-!AJ�(�GY�@w�	�CߥC�R82�EΟ\��ҟ����u'�'�2��%*bmD1��
�`*f`Ղӆڸ�F���y�c��5tF~B��w��Q�	>&k��1����h �p�_�fx8|[BG}���b�m��]��n_9�O�M���R�o�45;�K��̤�1�P�I`*3�O�ub�	S$�ᢡ5E1bT���'1Ol�14����i($o��}��k��|Ҁa�d�O����lAC���'I�q���RTy~��j.=�����'�R��3|�R�'H󉚚c>��ĨM4��M�F��OPt�ڎ`��Jvj�%d�m�s�'�����"٫C5�y	@�A�]D��-2?�|���3���hA�I?�0<����͟\ܴ.��ɀXЩ��Hp�)'��(R�|�O��D$LO�E	�m£PB!0�Ϟ�f�,��'ў���?v�[�3�ҹ	�}R7�^П��'Kl����>1����i^<�����8%�d��@����!�PÐ�jƖ�D�O ��bN�)9����� �x%��$2��t�?��B�Uc$0��lU r2����'?��0w�$�{�ܖb?Z	�a��4t�
e�ʸm�1��'#���P�aA	1����,��,���'e�]���?����d�trc���_$yc���> (4�Aj$D��WHEL���S
��P�#ړ�?��鉊�D%�$:�|�G�%�b02�4�?���?���������?����?y�w�P�� �.zI�"��]�@ݱE�wx9��)t�V�ٕ�Oq�'��AAQ��ZQ~�zg���k����wj�#��a)��0Gi,��e͘O�'��%a$��u�H4�q�����'��	�JlL�d�On��=������6�ׯ ���U	�W���'#(��ܡk�u�!凞9����˟�A��4���$�<ipÁ�� Ԁ1-�m��B��7�@k0��?9��?�����.�O���m>YCC
�q:5�c���z6�Ѡ�:��p�Eޚ/{ܴ��4��<a���f�? }��.�8$Cj1��V�t�h���R����"�C��u�4�Z�gA���4葰"��O���D�ےt��\JW�D|.DQZq+�3,)2�'ўDxR割}��1F陋����d���=)�y�ŏ�/�Y2O�~9�12���#��ƛv�'E�(4�6:�� �D�sL�%y$/W#<O�A�f��1g����Oz�� �OF�$`>i`HZ�<b,ٙ'�٨G�䠄���ɀ㔨P3�%ȕ�S�e��D�B�dΚM��&S�yVJ�k�FO�rl�37��h.��@���L�(��7�	9O|���O��cn�]� ����� Ц[cX@$���	g���J��Y����C!厈9-!�G�;�Ib�����O��6��;\� ��K�npUq��'��	"rI��[ܴ�?I��������S%"�ZX�B`�r�fYhv��>�p���O�X�횅PG(뒯=�FĠGL��Ԗ?!�W#�+��!��'��h���EJ#?y2�B')S��Ф�ݟT���xp��3��.i�lU,�t�p@�ſ
�$�e���j� �OY$�"|2��P�'�����1\�d*/G�<�]#$����DKK�a�>��`��@�'"�6ғF�Erqb.]<�BP���@��i/2�'+���[V����'���'0��BL�� �d��.���!�)L���p�I�V'j�K��W2�1��D&�����A���Q��L��m��cʱ*�<�ҋ�.��]�t��nxb>]�O<q��ԾKtdᐇ�!>�h�@�+ٟ$�'{��J��?��d7X������E#0������!i`B�I-D҂HY@�O��hT�%�֬D�n�A~���S͟��'������<��I�@�
���7c�������'<��'#��tݕ��͟��'*5�p�5��*?���#�і2��L@#�O	o��� �W�^���΃���D���3�x��R�d��n��Е����|���	�AK��y&�B�m����cO��M㠎Ġ8��Oځt��)Kva��ͤ��5���P[ 25�O�"�"������S$z�f"O�IP�Fk��$�� B��e�|�%��O�7�~���'pe�0�BG�Vԣ0�3��*�'��n�/�'�~�N�����"�+�ܺ0���&���jn�	pt$���0��[5N �n@Ohm(�N�t�H�����)��SW�9|�y�����O�C �'��`�J�sw�����đy��(�$�5�d�O���$������J� !�+�%�'1��O��=�'n"M�a�|m�dK�1޲$��o_��?�.O������������ԖOQvT���'�p;�)ʁ/"�<� ��~ؑ��'�"#1���&��)��:q���[�����	�-}z�TY�5���!޼.�	��B�!p.MS�ĝ5]�e��k�E\��A4��"�����o?"x�'B4���?a��	c�0��G*X�A����W�h%�"M#D�(�e5�ޕ�GN�NL6a�O+�n��>9h$I9E�"�RB��^O��b�K�æ!�'�2.:d垍h��'��'�>�6%`"D�	@~���KZ(���_� #H�E۴9�,�7�i$1��%�H�N��u�9@�+,#��ת-1��2Sg-3����r�L�b>��I<���Ӎ��EӰ�
�9�x��[?�R������O��$&ړ΄�i���P[:]rӯ�8�J���'�V�c�(~�
�K��C�z���-O Dz�Oh�^�h(6�öLpЕI���iE�2m�p�ӡڟ��	�p�	�uG�'eB?��@�q��E���'��T@|��A.(I0�D%T�@A��Ix��?YR�UY�m0���{� `�GB�8q�e�Fp[�d�O�Q�`��$�1Tuxi&��N�r=Qp#��8d����'*��'0�O�"|��@�o��Rd�0j1��qb��v���<i��{ʞdjp��jTc�j�ɴ�M���򤝃��ho�����ɓ @��Y��=�>��E��ϒ��	ܟ̳VM�����|b�H�%k�dh/��H�4
D?3@z%�0�*O��R2������↦�;���d֮��7n�����Y/4A�*ش`CzMY#a���A�%!҄G��z����	^�*��8SL���_/Uz5:5-÷�!�£WLh ��&�V|Wm�u��O��=ͧ3��"�(
6hh�"��s���Z�`ł��qP4�B�i���'>�ӳgE����NĽ�%�D|�j���K��]V<5��ß4AU-�	�ԡ�fg�9/�	���HS�t�?ڷ�Ľ~ؒ�Re��L��1�#h4?AW���0��)R��0t����4)7ʧY�&�y�LP�5T����� )��L�'l�����?	���r����H�3	����㮊��4�v�0D�X��M�F��z�+nRlhH �-����>� �۔J<���-f-.��t#�m}�W��H��?M��ޟ���Iy�M�/�M*D��p��$4[��q�1�ݤR�tI�!��x4@���]>�S�[��'Ŝ[ Nڶ
�\ �O��1U�-2�lm��I��� ��%G�l��'�|Z!�i������� A���SY�!8��MEƍ�e�p��al� i�Dϟx�|�'bb`�-ʾ��W�Q�Z6tͨ򢇋;[r�'Wa~�\�q�T�z���?=��+���1�?	��%D��#s�>�O��i��˓C{�T8�"��	�؂��(=�,��W��|�\����?9���?!��2���O��}'@I���.=X��䘓X�R��+F�~2`\�@�(��V`7Ԉ�oŦ�nI;���ҢQa5D�c�����H!#�(`U锞4�P��s��^86x�"�'�h���Ğ]$��#�fP5u���PbF�!�D�?;�X�J*RU���!C�a'�'�6�#��H�~���mƟ��ɻ9������)b&|AQ�^ wr�	��̂���ԟ0��ȟ�Պ6~j�H%�Ћ�Fڮ.w�y��K���Q��FF�8��iO�xd|A�	L9RZ��شyJ� g��bT��7���y��-��	8�Z���Olܗ'�ԩS%��kȈ����I�{�H�����?�����'�>-����(wTԒ�A�:h+���J?�O
`l��11���S鋵7z�5��,��_���۴��$�<J?P�n����Ia�tA9%��K_1/%���A�C �`B蜸)�R�'��`qs@�^�iҪEv�q��K7�DQ�?M�ӡ��ΈX�ƪ%�@]34�>?)C��U$��4N�&���s���uD	c�F�'DWz\kA�)Ѐ`�bP�0���'U����}rɧ�X�Q �1?:��7=�Z�Z"O^,��<GY`qag�D�Z|P����h�|(A�m�;~݈i����B����gӤ�D�O��$/1���:Qn�O���Or�doޭP�%ד[��ݫ%!T:%0ܱ���+�Ԯ^����'�F���@k>LP���gh��JȈ�	� �8��nӔQa�
�lI1�1O��c�Ґ
IY�B%q�@@q,{�Ba�',�#���ɟ�'9���2�M�jLhŧ�1爁�'v|��'�D}�����<��A�3JP�e��8S*Oo��$'���ܟH�'��R�ߤ)�x�C�@�<IB]7cңF�x0��'K�'#�/݁�IП��'j��mJXʌ�V�5Yl`H�P<t%��({H~��'�5��Ǌ�H�q{����^xrm��x�Ĺ��X�P�(\���'�$ع�B�b]�&HC�y,�hu���?���'�h�q�n�?�v!�%��T撚�	�'�����4G�d!d>V@J�ZL>�ֻi��'j��I�~���0p��R��O����(C�bDI���?����?�����Tc)�A�	@�{ �u/ꔺ���@�����]#V����)j��$q��/����AΜ��M� �D���`ԫ�(C���C@[�Đ�D�O��$1?q"�D7R(�Ir����]hQ�TV�S����
^�mix�1�+��bB
�ր)�Of�ɹy��A���W����Kݽa���<AP	N�t��V�'�bX>Q��j@՟Ļ3d�C��9�#A��n�<[�@������7}�|��,D�v,(���bX<s�py�O��$��<8�獣k�$-;�LK?���o���#�N]�^̡�A7	:�|�#�4J��C��q��A�g~b粟��	B�O��R.;�0�[G����x�2gD��!���3����@�v��@�3�ҥc�џ�Ë�I�D`i`�ĝ�18PE���ūz{��'/�'�t���gY�B	��'X��'y�N��(��²IH@ r9!wK�29�i �d�2,�J�����H�((�Q�)]H�����'ɠ�Bq�\W��]Y'��7k��0�
N�$	� VLG�T�Z�)� F��O����v��nN!�R�I��B�;�NT�g���FL����/�O��=�w�,d�!
�&;p��JE�S�?�ɢ
�'��Mk�Ł�:4 0��nB!;��0j+O-Gz�O��V����I��u��+�9<���4�S�?e�Lxa�����	ß����u��'��6�p((���3ͬ��� �MGDHr��w�=3"
V16��ٔ��$-@��yW�(�(OD=#b�j��	�0U2Ժ�&�3=��ФM���O-H
�7-�%5����?��޷"��#�C�]�~�rL�D��I���?q�%
���$̞=2��._�<��&�+�$�!$�;n|�U��f��<�M�N>y#!�q��O����6)y��r��8s�jd�����O��D�O@-�j��T�y�JP�,0�5�	�f��DZ��Զ �B`CR���%WD��$�h���������dK3k6��0�M�M��q�2N8����Z��Dz�퀦�?	����y�	 6��XJM��X��'[a|�ќv���M�&N�sq�I<��'&ў�Ӆ�?�2`�Vv4J�,A�)�T�(��� �'ڍ�QP��'����O2a���4�!B.+�Ȓb��O���H�m�X�+59���pr���"|2���uϲ�KgnhmR�� Gl~�+х�$h3Ej�*���٪J�A�)�i-gl>\�k�U�lJ�(^8k��	�M���d�O>�}r��� $L�R_�p|���h�D��q"O�E��`��(YD���O/o]`�r#���c�����:��K�mΝA,���!C��ʓ���	�:���d�O����O�ʓE0�U��fR�h��,-aLҬc%Z�(	���3�'� [5�����Ϙ'#>��%�N&D�=zg��jCb�T��j32�33�^?Eu=�I���O�����>���.t�Z�R$-��l}�5�fj�ß$�'���k���?���d�BFVq�/�'j:�*6��wnB�I�4\���[�/�J�����Z�6���O@8Dzʟ�ʓq��3g�2&XH��$ ˟/���1�G�'�?���?������� �N��ʖ��JLZH'�]3���c�"]�[	�h�E ɬG����I%l}`�*"��Ԙ�.\:A�n-9��c��Aᡕ*�=r$�4N��!���0�`�7!C�a���H��1����O�d&��Oz����<�|i��:+��|¦�'y1O�����j��Tp4�A�wހ	�|�O�>�+O|�&��|�:��12*�i��rce� h;�D�<��?Q�a�^\���-Fʜx�5����
�$Ϥ�s�Q1p�L�
�ʝ�0<�ԫҩg��=*e��<<4`�	�v?����'��5��Ys��#�N�sdEU�K��@����O���&?Aq��DZ��R�U.�N,�W'�O�n��a򇜝`�ޜ`D!�=a�2���'&�Id����l�O�����u�{��P�(� �1��'Y��9J�$�����|J� ���r��I���p�[&G�����?��\=hd�
��Y,M�is�����
����P���g���X�����?]H0��gȬ\Q�g��>)J|r7��$krD)�"17�`�J��{~Zi����O��}b�'q�XZ�Ǘj��u 8Y4���' ��Q�i��~�1͕4U�԰���O*�Ez�n�OV��L��!�"+ ��I^y��F#���'x��'���xF�����I�\�m̤��y�dѰ0�Ҡ�Y�.�C�-X\�g�'.ԡ����?V��������b8@�@T�{�^EZ6*E�EIt���[�'t �<��P���5 I�s;V�`�=s�^!��@�O��x�Z=�	؟(E{�d^>���CI!�
�� ��=4�!�D���V�,�9
�8pŃ���R�'4,#=�O$�	3n�`(4��2A�b��s�Զ6J^�=�[�!�
-PÇ��I3��O��<�Z��b$*ʐ�,�2r}���'ڠ=�2�'���'��()1�W�<}Z���/��4�\i@\�>����-�RdTY��Z��4z�e�G�h�2�L[���QL���Ү�2[1a�`���ɺ%;���Oc>Y�`E�}����S'V�P���Ϊ<��2�Ҡʑ���
����ϣGJ���	����D;��g� >.��M�EMF則 ��P�I��'��S� ��{�)�`!G�\WΘ��fpdF���$y�����H�M�4`�`��I��͹�SD̨dQ5�8Ut�g/��r�I�b�1"R�J�k��p"*�t�z�h6���O��yc���I6	;1��4:���r�'������?�O�Ov�I&��Ѳr!�>v�	V&�0^b�B�I:�f=z!�1��h�	 ��� �	.�HO�I֘8 \\ꢌ�N)� ;�F
 �d�<Q�@��?��?a����ԟx��)�p�p�[E͋XN��ڰ�yب�i��оo�b@��S�.�:��'�nAӠ�ۻ.�j�A�ݎ*#n��si<)�x�ѫ�ßl�Q�Ҟ��i�6��&�P��!\��Xx���>g�N�P��3?ɶ����	B�'
�
:Ւ\�#�9]�jr�����5l͸��`��f蝪�	��dDa���D�'��	v6^1�%�u:���mҀi�PL��,�۟��蟌��`y��$�Ԩ:�1+����\�|�g��5���K%���Q]���7��<hδ�0���e�'��]�Q�2X�"��#$T4�5mХ �����<p�ZA@�j���s �%�HO ����'.ظ_�kv�H���2_5�5c��'�ў�G|�,
	āY�I2C���K1����<��D4��4�s���8=�g � �	��M#����D�14QP�~RE��:\jH�6�V�>E��J�h����O��$�OP��)Z�-�T��/A��B��vf�
�u����BB�+:�)
�-R���O4a�ІA'��I�Q9UIx�+ ��5mT ���V�q�ֆEF(�q��I�'BJT���?ُ���J�#�!���P�,�vi
�8��d2�O 2��38H�`�Bٵ�Ń�����hO�vy"�ۈ7�L����	��8D����ĝ�x���Otʓ����Ov�d��H�(�S�L$;���P&e�uv ��������Fu,l1d�1x�����)�jO
� d*��F"����F�?W�Zzϼj�d�mK�d���
\&�5�S�'����E@W "3JpR�ӇL ��\t����$�䧎�� �t�FB�oS �2a?�j��"OQ�B]<9Z :g��G�̤����O�Ez�O/,� Bc�]�\��d�#{~�8'�')�I=S� ]������	矐���4��9-ɚ�"�/�#E��txc%H��4���E�V�����C 0�L�ʟ^Y�>���%ZeJ���:�������:}���K�`��%����O���ئ�?�d�3V���Y��C���eÆ�&S�	�,�x��O��=)�'��̨�L�*b�xx0��S$�u��'}��K�hHd���	��D�����'tx#=ͧ�?!(O��C�cs��QR�Ov8���\�%v��@���?����?�*O1�����$xi��$,v�x	�hO�xA����.�>@RuG��0�<@��R�'/8��ǟ"?n�z�eʍךQK񎝛#U<aЖ�>]0~\�%�. ��q�>ғ�0��	�
�d9�3`WS�r����2B�I��V�'X�,I�	H�n�#@�D*��$��+#<O~"<��i��:9�Sf@�A5p̩�My�q���ĭ<y���Y����'d7��E���jiƉ�&���dn�k��'=�&�'���'O*���%�lC`U����tFN�
d��ݺ��aΙ�`�g�U�Y	�D�6�Xz�'7�|��l�Lec���z�T3$�o�Mۦ�V��r��C4g��T� �۩Y������E|�	�[����=�i>qRF�8�c%�YO�l��$D��SBP	_F��㶯�F�ؐ�%��!��|��\�0c�L�Cl6����	h�@@b��<���?����?Q����)$�C�.#@�Yum�tӠ�ht�w�E{�o�d�z� V�(P���W���'��RN<���Û����x��C
�)�
(ʚ6m�O�y@A�b�$
���Ot����,�u�$r�?Mr��2�� f�쫦/����l��$��ޟ ������ם5����
Xc$�Dȹ�*0hP���,��?��~����'��.�O��d�����b�$Y��ɡ<�v�q�#��-f<d�qOg�d�D�O)���O&�I�?���s���r?1��<S*4�(�aS�T�H9��P6�?�bS㟘�I�#������O��i�O��R$� �54�ɘg�Č� bB�TER�4�?��"6 S��yb�����������4�9�#Xo�ي[	�h�BBAԦϓ2�n]����$��'B��?��'bN�p ��Hq�F�xЋ��j���Ċ��y��
�?��bK���O��/\���ߦc���6C.x��#Q�U �T	�ʱ���<�A�ӟH�ɫ4N`�'�?Y�LmZaP��T~𛶉ؓS����ıi�m�W3O:)sR�'�b�O6"=O��9����R��_􅁣o [z�*�GuӤ�Y���O����T�i��I�<�S�8��,��O j��΁.V�fpH�'�5�J�G���.N���Mݴ�?),O"�d�O�d�<Q-�kL�r
S�g�*[�h���]��IƟt�I��`�'&�Q>u���TE��)xW��B���`��>!����d)�W$�;A� [�H�cF���'���'w0�� R&EAF�c ,ݻa��m�'���j�e{$f��f�O�*�ڰr
�'���Ş�C��UWꈒ"�М��'^���ㅅ H��y5E����hy�'Z��heM��1\���a���,���h�'|� �%��7���@�� �@���'B��JĀS�c�4��D��4]�I�	�'-���r�
�88
yg����Vԙ	�'��qM����EqF�
9�l�@����Op�D�O����O�г�^�j}V);�(0]��M`æ�����H�I���ğ�I������0�"�F�:F-ش�a�,��7�g	mڟ��	ҟ���W��?y���?����?����t��a�N�ǈ�9Gg�-ݛ6�'���'���'�R�'���'�����#r���F�<%R=���6\�@7��O����OT��O��d�OL���O�$@�9��l�7`��Y�}��,���mZ؟H�	��0��۟��I�������ɤ���zC*E s�:(C��M�0�J�4�?q��?����?���?y��?�#op0z��0C1�A�GoԀK�FY�ĸir�'�"�'���'�"�'���'S�	�S�A� ����$v��:��oӶ���O ���Ob���O,���OT���O�9���Smfq;S��� �'!ޱmZܟd���T�I̟���՟��I��x��5��(��yFt��f�<%W���ڴ�?���?���?����?!���?	�h��b�;m�b��;����S�i�2�'�"�'b��'lB�'ir�'�z�r$/Qm~I� 2x� ���s����O���Of���O.�d�O���O��nB�c�@��H���9��mu~"�'G�	N�O%��IA�_��,p�܈$�|����i�"�K�y��I���͓n`��� Imҵ��VL��޴Aޛv1Op���'"���*�h?1�$�?@HB�2ԧ�yI.d�bE��P�Ε5Fw�9���v���d:ON�he�,ƨ��H��B�|Y�!�''��b��M�0�Hl��� ��BI�`ׂ�Q�Ğ��B��$�^}Beh�. mZ�<�+���K� 	kx"<�B2�����W�H��&V^�z��.+?ͧ6�<��V�y�@+h�����a�tZՀ,��$�<Q���h��d��T��AWn_�Ӥ�h���&�lwӪ�����iش��������N޹�t��f��3Gk��U���}ӎ�n��,fk76���Lw��c���4xkםv��ŋ��A
M|�8��G�i��=a����'�S9�P�K 5��%��@��e\˓4N��/���'Y��x�
��z�b�!!cֽY}��W�h}�l���o�<��)��M�f�b�B�4H��tJ��" L�D�L�.,��%"�Z�� ���[��`�b���L��t�#�ј.t��C�?D��(QlJ-Xf�9鄉\(bd��?扝(`b�:uo�ϰ��&�F��e(B���]�������M� d ���r�}j`��( *��pd�@.���a&߼0J�]����y���A�憴+
*����2BD1��7R�\��p�\3E@U	BXgc*-�UN�[��z�V�+p�Avf�2[�x����]2EDEY�FYns}��B?�����e��M1��]��R��K�9[T0�9�J�Y�6Z�Z��M҆���Y��p5MT.>���(��ڀ=A�����v��!�Go�	mΔ�+��cFO%ӈ{`�I5@$�.t�����"ǠU�eL>+��)��ڈW��(�Ӥ�U��R�n˛8����ʂ)9�!����?�^l��Ֆk�ȒP��a�$��`k��"���Ǥ.\�E�վA��˲�L=tX����H0ie�}�
�r88�T�ֹX���	� �ɢ=uN�����")W6�����_>��I˟�&��	˟<��Z̓F��$�wǝ�DX�#QCM�y����	��X�	y2�!J�������?�ɠě�[��<����7NgE��"t���@�		~���?�'JltpaU��3��S`���y6v��IWy�.X�9�2�'Y"�'[��_�p��E�H�2�P�Q�M� �H�#^ПD�	��4k MTJ�Sܧ8���s�!�X�Li�� C3�����2®����$�	џH��Gy��'@2�HJ�����mM4Rkpd�TO� Q�2��5��O>��	#~��A��)ѷqEƜ��:��m����l��؟`��^y��'f��'X� �����h�d��� �[8(B�O���0 (���O��$�On���.�So���Sg]0�\E�&+�O���X�QS���?���?AO>�RJ�%A���l��+�'ҟ��W7c��Od���O����<��Q�K|�t�U�h�|@�j*��L�-O����O~��2���O|�ĕ��세7��oآ�9��I�(�>�jR�.���O���O��<J��O"�ݐ1D��K� ��Ga��a����?�Ʀ}��x��x�	�[*�ϓ$B>8ҧ֐Y�=�s�T6b����'sR�'�b^��!'hc�$�'���r��9P�p��ȏ�F�h���'I��|��'Hb�B�j�1O\z6C�d�������<�"h1��'_��'m�	�2[��OiB�'x�4��hvLx�a�4P��E����!��'���'�Ԍ
�'�ɧ�4ΐ��|��!�YY
��0�,�?�(OlI�r�O��D�O��D���ʓ�<4�뗟:J:�#B�!{p�����?������8����20 <��A��9t�は���?!��ذ�?���?���")Oz�D�O��;�&� l ��eǙ2 �����O�)1F�+�)§�?���.�D���s�E+$��� �J�O���OP��̻M�"��?a��?��'�H�$�(U��(�8��͓��'2"�'���	DA4��u�۳(y"�QFȔ]��'�,P�K�>�,O��D2�$)0}�4��
H��ٓBJ�)��@J:L>Y���?�����S	r�j�f��鐐A�� 8���Z�՟��ן��'W�'�L��4$ʟ2�8,� �ڥ8 �WdZ�ym��|��'v�\�4�g-Z+�P%ݏ40X| g��U��roQty��'�r�'��Iן����<����	|��HT+�5Y�<�CЮ�e���'�b�'s�Z����-$>�P�Iּj�X��w%��
���F�"�'��X�$���,�`L����O�/�0�U���<9�����Ol�$�<)��@ ��	(���$�Oz杖^S�-["�K���Ac�q}ƒO��D�O�����
�1O�	¦	�����.[�I��#my�Iʟ��"��\�	������?u�'�~,�������U��
۵I%(��2�'\2�'I��*�mM%Ә��O��8:���̠�%�)<DjYP��]� %(��?���?9�'��?��	I�oz�d��
Uع	�M�p�G� >iTb�"~jPC�
<��(81�@>8�rY��KР�?Q���?���+Ĕ"-O�Z~2�^� �d������Ɔi�`킿>��<aa@"��'�?����?b I�lFd�� �7����Y��?��rᲈ94�x�O�R�'0�	6?�Z�F��?��X��b",��	��*�E�ޟ����4�':�ڟH��͈5	'�h�bM`RlK�R=�\�'q�	Y���?)�' (֣B!N�&��2얹}�^@Z�����'��'x�Y�<���֨��s%�>�0�R�с �fEP��xy��'F2�'��I��O��A�#'"d�y�J���-�0�
�3��'���'��_M�!O|
�G	�k=Hȁ����N�<�@Fe��?���?�,O���|�����I�k��@I�'	$�´ڷ��_WB�'2��r� �c���'r1�� ��Rgn��z�\M�t&�*����|b�'+�I"�"<1�-sh # l/� �0 �����OD w�O*���O(��㟒�s�� q���`6j�;���(�0�����?	.O^�9'�)��Ñ!�,	�[+N҆�(���?�u]�?����?����
/O��C�Hs��L?l�(Ke��IgR��'�Mz��ᓺ5VrR�!�,($48Y���	����	�p1���zyʟ:�;�`�s 	�@�jD��(R�+eH��9���'�?����?�7�44:�)�g�rSVU�Fa��?Y��8���i �x�O0��'��IN�5�`C���vs�AG�3z��	Sy��'���ӟ����l�'��u6�1g�v47혌d���T�Fr��O���O���<���?I����JT(�x�
U��g��S��d�����?1����d��"�$���`Q2���A�b �W�[�8��e�R�\�	͟��Jyb�'5R�!G�-P�n��'�b)��aflC7��I������,��⟐X9��7��O��d�9RuF�8҉A;�L�����> v��D�O8���O ˓�?Y-��|��O����(�.2����Ў>��-� �'���'+r�'��VFx�8�d�O>�d�:)r��n����D��b,6)�O���<���_k>\�'�?�(O�阖`����`
�buP��G!�/Y��$�O����2��n������֟����?}�ɇ|F�q�#�'#~0�m��}k ��'9�-�,�2�'��i>��OޤP�0�
(=v���E�ăd�N����qWh"V�i�"�'���O<���'7��'.�UX!��>�F� �`O�
�p1���'����'�Z��l�S͟��a��3r�,�q F�ooq3����MS��?��2��0���?a���?���?Q%�@�Z��	����N��?Y����$8B��,�D�O�����Y��F�$<��cvC������O�幤!���m�I4����r����	==Bl����`p�:KD��:Ǿ�̓����O����O��$�O$�(��[Q� �����[�E�}J�lZ۟��	П,�I��)�<Q��)�j����+��5kG����38d���?y���?����?���?�d�G;�6FC7vT L��#� V��riP5q?"�'3�'���']�	��Ty��r>u11��oخ�h0jD?K~,�Sm˟���ǟ��I�����ҧ@��MS���?%K%?a��"�(�1���� _��?���?������O�Q��1�8�Dv���&�^- �v��f�\7�s��O����O����O�!@ă������8�I�?�;A�7:0Uk�K[�	g�(K�F���Jy��'�PQ��O(ɧ�D���F�j��I�4�p(K!	�%#2�'�R��)�7m�Ov���Ob�)�����	�oTvMaE \�)<� ���)͐��?	�Q.�?I���4�x�'�T9HD+��W�j��#�+%=���ɤnj��aݴ�?1��?����R��?I�6hPH�$�rR0=jp畋UU,��i���(�����|*O~*��N(���A	�$�g�22��!I��i)��'�7q���'}�'��')~�6�_�=Q�dk����E�H0��'��'G��1���'��'���Y�.L[�����C�	� ����'��a�>%:6-�O���O���FG�4;O.-Q���wĺ�p���(s��L��'mR �"�yb�'�2�'%��'�哓�jk�f�b}��	&��q����d�M+���?��?a�\?�'�bGsw�m�V�T�b y���Äie��)�'#2�'�B�'T"R>]��^��M��L�	q�*@�� �6��6*Ƒ�?���?	���?�����O��Ra6��1���=?�@b��ɷw�H�����O��$�O���Oj���O��������I�|� ��@�qRe+[0���E,[�\�	��I@yb�'7j\��O���J���H�h1#ْ���Hٌe����OP��O�����%�N�l�� ���@�ӗ*��@��H-'�n�j"G�a� ��IΟ(�'�B�?	8��ky�O8J�
օÚm^$a��g۠P�j9�#�'\�	\u��4��	�O0��Tmy��/3��q��98�MC%���?Y���?� jv���O@�<	�&�$tv"�gԉa����&k���m�֟���ٟ���'e<EK��U�Q�.pĮ����m)��'�����'��'���ėK�0Qը���0ٳ@Q/c8N�m��0�Iџ�c����ē�?9���y�`����'�6 =������?1N>a����䧗?i���?FJʷj��������E`�K7�?���]Xf�
��D�O��O��bY6����E�J���CǒdC�ɉ]T�M��my��'2b�'�剕�܀aJ�C;b����ũ��!�	����?I����?A��}$/Ī�p����8rN�T0Od��?Y���Iv�x�O�*0�eA�k�>C�,ֻ=P|�a)O��$�O֒O���O2H����Onu���ȡ6���y��i��D^�ޟ��I֟L�'s��f +�I�|W`��(�np�4��5dB
���O6�O���On�3��O��4>�ݳ����8���ۡ�[�q$�������	~y�.S�j��\�����yP�/Z�싇(٢V����c?��O�����uK���Ӯ,�|��Ԭӷ���@a�4gh*��<��<aӛ6X>y�I�?�.Ofi��2L�&��F�G�+FNşl�I�� �-|�Sܧ99dM��LI�#�`�a��Ի�h�IP�x"�4�?q���?��'3G�'B� �h0�$̪D���3,Ϝ!��'�����'<ɧ�4�d�J� ���>۰]@'��6�$�mZ˟�����T+ݚ:�ē�?���y�L%b���ÀDu��$c 㕻�?9N>9u�>��'�?����?)��J	Æ�R�
ܻp�����2�?Y�wyh${6�x��'��|�66��R"kՋ"��`#V!�.t�I��u��'����	o�P=l; ��2ZV����a/�Ś����ē�?������?��h�`��Ø�VqfEc$�Z�����d)\��?q-O���OX��<�֌U�:�����):x��n# |�1"�%����O��$���O����B���1Oi� �m���x��&07$��?���?�(O���G�Wg�Ә_h0t��J�}�S�O/8��!�	��t%�$�I��lyvl|�&X3�)Z?_XH�2�U0�	�d��ty�Mò>����dퟌ��
�C���9�����I9��<���O��$H	�&���(Z�M!���2�
)�*\$-2��D�<y�d#��F^>u���?ً,O���^�Mj��ك�<=�R^���	�t�I>I��썾.�@uM�x<��+�M�O�[����M��ޟ���?�H<ͧ-�>m�C� T�2�S
-�N���2�,({���?���h�x���)'��iQ���g��P�Mڵd���D�O����O|��`��<�+����k� �I�� c�}�f�y7B��H�Dn1O�����3���O����O�x� ���v�:��TJذI�z=�M�O��$A�!�t '��Sڟ��	o~R�ʙZ��Ҧ �>||�l
��X=���L� �1O���O���OB�$�$L��$.$>@�Ѩ��ג<'ԙ&��<���?Y����?Q����\+0�X�K�$���ĝ)k,dU G@?}�r��'���'�bY�(10d���e�d2F�:!��j�l�)Ly��'vB�|��'wB�R��~"D��w�\����@�)r��:��d�O6���O�ʓWўI3��Į��`y�ƅ�g^�=`�ႀr�'L�'s�'��t��{B��,K�T(�oI��hM"!I��?i��?�)O�y�&)R��ɟ��SmE\*'���%��k��_<�­&��	ş�g�,�SJ��[Hx�S���$��Q��x�'N�`1 d�˧�?���}#�I&�ҝ��HޓJ����O7D���O��d��r���>9:���85-V��8'L��V�˯3��/٦�^6m�O��D�O�iK�	⟜��b�4yA���!s�bI��Q؟|��&�S�O!�L�E=�c�,�,<[�0�%�i��7-�O���O|5IG�r�֟|���<�d뜈2�&\-B��X�j͌�8���'0���H�I���`s�58b8����ʘ9������\�� .y�l�K<���?YL>��E<],*U� @<�`�(���dH�A�1Op���O:�d�<!W�ǰV���Z, ��0���a�	ߘ��r�x�'sR�|�'rb�F�n(��+�A	����Ѵm�2�y��'	r�'��I0Q"����'B� �(ցV�$f���`�>$�ݗ'���'h�'���'����'a@�I )��ۂ�1[ܐ�/O$�$�O��$�<q�M��YˉO
�D
PnP����1%(H�6iy�'�2�|�'�BdƝ��'���i��N%k�ڐ�B5
|���?i)Oz�d�TV���O �$�O���C�2$�@"�r��([��D�5̼�O����Oz)�ʹ[M1O��g���r�ȟ4Z�U&Z^^�[�ȳ�BR3�M+*����jD�'U񡔌A�q��.���?���?Q@�[���O����iΚOI�0��Â��l���n�L5���i��'��O͒b��Y!Z�F�<;`�,O�~�k��Rן`��b'�S�O`B`�N𤉫"k�44�2\�g%�<n��7-�Of���OTM���z��,�I�<9T�%�2E+�_$j��Ȼ��w��W�i�<a��?	��$Y�rX&
�$`��⊣���i��?An��%(�'U��'[�'T>����N�I��M��T���S�H���8����	��t��ϟ���!G9O
z����B�	��HRm؇�?Q���?����?!O>���?)B.�+����*v�|�B���>���<	���?��?i��z ٙO�~Q�F���i��D�/�w��������O��O����O̙�u΀	 ����TB�AcZ����Z��I��e�<����?9���$ܛ|	�d�O02��b�Π���!����w�K�X,B�'���$3y6c��ڠ��1gh���N��|u)�O����O
���O8x2�ȩ|��?��'.�d�r���L�Ҷ I>/YZH>����?�ŊӳxE�\�<�'���Фm��9h��� ��R����IH�IА�@qcǜb��A�����8D���?ͬ;Q�H�&6�!(VnG�D�\h��G��n�r!h��'�	��'Nr�'b^>�����ɭ��?�B<˂f��3�ƍZu�ΟP����4%�T�I�d�	����2Y�(ش0���%�&Bt����d�Iئ-�ɮ���Ob�D>?����0n �%��X\�^4@K�.m�*��đ"�x��l���>1���?�ˊ�ӯG0Э(s�܆9Ul0�KF��yb��+4"����[�Dv�Ȼ��Ԯ@���Ï"G��թ����!N`]jE�yM(�%+׽ ��DQ�F�A�@��� (ԹBoҀt��Pal�rn��L�����'/ڮ��a�n��x�jٖ`�H�
n7�C�J	���ӱN�	{0 P��,K��Ҳ�(#�(YQ`��n����蟰��џ(X��\��q�4��I�%l\�ʡ�ރJ=��a��#D� ��5a�4.����e��$��|�'��� EB�:��eh2�̭}
*\� ֆbFnx��o��$HۖǏ��u'�iXR�q4�O���5����D�P	%+ܤq�>膁QӨJ��'��'��	��$�8 ��	Sޒ��ҋ%-�z!�<D�|S�/ؕx��;�"��	���@#�;�C���'��	'@Z�D��4�M���6b��e>�`ؒ�R�0���'LB�J+��'�W&*T<PؑOޫ0�u ��ܑF�np3��^��p؞�(��9P�d��Ҥ�V8��ʟy�P0�wV��������<ip�^��4
p�A���<���P�l.*����?�(O���%�)���[?
�Z�&^}rj{�.F�7z!�Dǥ/�.-����A�����> �t �4�?�)O`X�6gH�$�'���0���W)�$t�����`[`�@ݟ|�	��X��k@,2Hl�T��-Et�ڳ�Џ"���Aݺ�Uh��xUД2���R��$sU�b�����a.��jFx�0@�i>B�����8���13r���Im�}  1�}r�D��?����H���HvJ�#SH��b�W�sj����ILH<�dM͙c�qi���+oD�4$�F����{�-^d(����IU�8��!XߺQ+������IȟP�i>�!��Fڟ��I��ml���[����EvV5�$$�.6*v1��C�q-R�[���
K%�8+��XA1I1�S�y���#�6�2��[0J�9�w�ˋ}��\� HN6u
���'���MPp\��H���6 '?���w��h���%cּ���Ϗ��
c��ON�m�>��D�c�>��w����V��=����b��(d���7��O��d��� MN ���P��@�qO��Gzr�O:�iQ4D�tNM�jH
��م������Oو���6Ј���O��D�OD �;�?�����G6?�@�X�NX�&����7�`��d��7�B�!�H\�\�Dnݍ�kC7'�Ov)C�c����g��o`�E�7�۫$R��B�Iu�����?HS�Ng�j�X'��g�_U�٘2�	 Jn�$'X�i��5mZ1�U���?�I>���?	I<Q㨁�����*Jv�iBЭHO�<�60]�N�XR
��4�(� �_�'�>7M�O�� � ��iś�!�'P:$��EГ8gp�J��i����O$��Ę�l���O������̚�]>�
נ�0!�t�Kt�^������+`���jڥs A c�	� �~���6T�1���D�
���{�����U�V*IӅ�ÇO -�F��㟨���O(Qn��e�Q������qE��=#��Л>����?A�J~�
�3P6�q��	��\�	�j�<I��]9Q$H 8d<`_H�	�.��$6��Oʓ��95Q���IY��"72����ҭ
�ڵC"A�����'��'r��#�ı!PF(�p��6>��T>��;?��@IgII4��Q���[�n�ְ�>a��-���'Լ1\+���j4u�pPЫ�b���6`(��'b�����?���?IH|�+� l�1�j�$�p���� ��O���<�ѣ�1� ��@�
jhJ����X���k�{��ܶR�iS��p����!*��!֤���Y�����i>�aw*������ɟ�o�$ndL-���-"T( �5'ð�����l@�Hr1�O$C �rR(�?��|�'<D�A�G!�x�@FĐ'.��� %&$�$apu懜<Dވ���H��	.I6Y���Κ}^|�do(^������?	���?�()�g}�\��ֱ2bm�=|}�=pa�\p,���?�O�z$���:�ȥR��2�Z
���s�'��S���ÐK͓s�|�Y&e۟L�4X(p$K��?��oP�Nulɉ��?����?I6��:���O�,A�M�yS�@K�#O�DC�Y!x���\�1d�1BG4HD��_w����J�W��( L�q�+�*��udX�������$�X�kp	Qk#��H����#�4iE�����Q�����+�@���rۆw*�� ��?�0�in�O����O�O�Rv�Mg�qP�'Lk a��'L�@�b�z�l�
�n2&�>�C���Ŧ��	By�o�%f�,�s���2eL�FI���� q&����	ޟ��w�͟��I�|�t K��i1r��6ZO(�ӱ�,T��)��ßh�<���))"4xc��Ē6z�ߛ<�x1wCȅP��9���\�6������cdT�!F�rZ$�A��x�ܓO*�A��']�7��?�*у�Aּ,4���.�_���[�3�Iڟ"|�'���ytF���f����a���@���,�'+�b���Xp�P������ H���o��$�<��|���'MrT>1X�M�X��:�Lk<x<�mCe�������ɧa���)%�@j�%���YV��+gKO�Q~��;Y��z���0�h�H���3Y���>��[&t��y��,�?��Y��ur'��* �n�r��2vB�L�i�3���I>�i�ҟ|��4mě�'��O��j�.ǌ*������AZN��4 /�I�"|�'+�H�1.ܖ�*ĢB:"��l��'ў������ d�S8FV�Y7�L�PЦ�"L�s���kD�Ot���O󉏮,�����O��Dv�2�� ��T����0m�6���R����%a�7*�dD"uKl�p��O}��6��*X~�-�2��Mņ��Qi��:������)�7�֠*�������aB��}21�\e"ı{b�r�#42���u�U�d�4@Z���'?zD��O�����Y�prv��ɸ"&Bu@ �Z�����	�Q4��3N-)(Z��ߐ���޴�?)H>1���?��4k�ً1M��X}0����¿8�ಆ�'���k�9T��'s��'{2�֟��調���@�y#`��h[%h��p�e�ڡt\ʴ�ǦQ��nŃ6� �l�ΐ�2�>�B��e��Ԑ��)Ch�$]�|�i�/��pw`tkGL�8/5��4�d@Y��9�=U
�0?�r�� V`-c�b�%	�'�Ob��!���OF��"���]z��Rƥ@+9O�$�TaB/!��K�9�>a����4]��SU�3l�Q��8�O �<��U�a�ij�V�|��Jӣ�Q<�]��C�GE��$�O���[F�(��O���\�fQ^9��+�Wnm! ݿb'𙊴��H �|��T4B"Bi"�$2��O2��rF�h�r��l�2W�Q���VB��a�k�
�$R���L~,i7j1ړD���I*�M�Q
?4���'�F�l٥͂2"W��[�����O���P}�d�/�*�h��'zo��@�˙�y�e�U��}���ۦ~��-��ߚXJ�4��ƦE�'��#�u���񟴗O8��f�'b^��qQ�=Z�(,St�Ҽh�2�'%��*|��}�Gk/J;\Y8�䍽j������Q ��oKb��4;2�Μz�w����Y ������Vd^�c�
������ ~�ݛׇC ���y3�d��a|��'ȑ>�A�iH�N��|Zb*�j�̚q�S��?���h�^�5�ŃqV��)՚5	���I���'�`<�q�×<_����F�.�����βO�2m���I��ӌ*��I֟��	Ȧ %*����
=S.�Y��	�,䂈�k�HD2��M��?�џ�b>�*�\U�穇�S�l��'��f�ȑ�K��<����:L���$�J���D�*f$�bb$N�D1��@�]������MC�X���H?��R��mL@B����Z�H4�T�.y���� 0��D�e?xbu	(�铗?	3鉧��$r�L\��"��NJY᱃��#����˄ן(����Ed"��	Ɵ���Ɵ@�Yw`R��U��,]�0��Z�L��^Ըi��O�*"D����D�X�ayBM�9U:5i��9%vV���l��}��Dk%��a�
=za�ؑ-����\w����%b���'&<1.��]���C�ʌ�4���b"S��\�F��q��4�?�,O~�$&�D�/=KdmJ�A�z pK0DlP���<9�Ox9;6a�S�0%ią	��2����M[M>�2G ��2)O�Xը�ܺS޴c �t
��"�N��תօu��8f�'���'1N鑗�'�'��P94�il�F���Q)7�m*��s:JQ�� �����'��L�Rh״��!��U�I���C�˲1Þ0�R���:������R
�p6�։TvL�[v@<�Ė�T42�'��]ŌA��JQ���޹J�!��E:P�Z���	S�S�aU����:��%�"��a�d�>)��xӈD�BJ�d��PHb�4��w����Mˡ�i�剕"�F�#۴�?Y����I�}�$�"s�����I��ZX1�H�)�O���O�I��eB��p�������@@B�Վ������a��6u&�ĸ�b p�D��na ��I�R�@۔c\(��ԯ;:?$���3r����M´�h���>z@2@�H>Q��������ϙ �|u���w��%�fR�D�!��R%H�8�ʀh;`��3��.��$4��|����,B�t�G�F51�B����-�^4��I��M����?���|
R%M��?����?ݴt�*�2t@Y�LqR#�L� �3���*SiX��&�<%_� �΀j2H~�'.6k�C�G�Ɫ��!��D�6���#B�:$C�jA'P��H����i��EQ�a�=Q
d8����,
�83��?ѵP�lx�:���NA%`ʀ���Ԭs��1d�\p��ix���Q#��֕h6ǟ!e5���X�Llb��kݴ�?ɉ���'�v�)!zʐ�`�B8t-c$��;tw&���;C�.��R��O���O��dS�����C4CD;c��˷̍Ш���l�5rZ>�;!�6U��p�!{��ܮ�8��<�O>�,3&IZJ��L��Ǫ%��p@�A�H��!1��x�֝��M�CS�~�RP�M�$yPf�N�r�
B	���C�n\�d�q����?Q��?y(Of�D.��$��<S��T~��3�/
���~bX��� @ xNT�ر䍫!1��	p�=�v8�&�'���M�ӟ\�K���2(�0�Ԃ�8���"O�<�! ߤ �,h��I���9H#�'�<̺�L7- z4�1�Z&IqZ\@�Ya­
Q�X�<���L�/�JɹG�ӳ��:F�|�<��.	�y������''�pU!Q���<9��0aJT
˞g\,H3bG�x�<� �З�
>O$�d�ր�P�\P��"OH��oF�vψ���EW��ِ"OL�h�V�f#�Xj"C��Y
�0G"O�]�0��<1���׫4_|�c5"O�u{q,�
`��`�kM0.���"O�M���أW�b�Zt��'HyB(q�"O�	�VO�-�x�_y���r��YX�p��3� A�������iwLU�N���)�$�5E��Ԇ��`�(��g�D�兆:U�|�Ex���2���cg��t��Y����T���%FV1��$����@���y2�J�$aB���%H &I��;�y�ǅ�� �Z��zxlk	_4�y�)�;9d�u۶��@���f
�yBI){7F��5��xj��5��y�M̵
�@Q�C"�HD���y�F�}V��T��U�Qb�NE��y2�]�a��b�/|��s&���y��ER��+��ݨi��͉�hX8�yNԷyՂ@ȗX�^��qx�&߱�y�JQ�Ţ���J�\�]�䙈�y��B1hjx�ڬe2�hhGJ
��yR�G�w�fy	���3Zj��&,ط�yE8�b�r�j.&��|:���y����*�r�3*� \c����yR�O�M~�Hp��N�3���3�yB�T�`צu�Ff�@L8Y�Re��yRe������
�/<{�x�5g͗�y�V!_RI�%ϫ%~�ڧDO��y�*Z�.؛�c���x��Qʝ!�yrd�~|hy�T�R�2?ܝZdAC!�y2��>Rf(d���B*ɈcB7�y��#8� hF�,��,У'�,��$��1�`I�F!\O.Pk�&���B@B&����'\�$0 �	�^�a�C,[:x��PMc@��h�k�<�"��6ȑ�`+�� x�i��(\b�'��{����"j"�3A�	��	�Mj�Nν7�R�"6L_�is�@�@��d��h���&z��h�jV�(��$ˑ�asXqr!G݊�2�Q�ʢ<E��'���%�T'X%�� ��Y{\�9�4���9�j�+�p>i��\"^��`v�_2<�dL��<�u-�`{��e��2͘'z���!C3N���������ݣG:.�E'^)DmB��8�^ӊ�Uv�l:RoM�/�nP�m�.}8}0G�Nf�y4]`��O� ��"~�Aޏ(��$D�]
,�(��ǡZ�'�2��,��]��a��Ъ

����aW�z�����Č8i��` K�9�>uܢ|�'�l|S�c��%�,Q{�d��6QڢLF61��ʓ�uO�)��<)E��5�p.�;u�5�WʖR� �p�cQ"�H)��	#(�-C �-Tb0Is��L���2�l�zU�S5d����<i�7b�����Jm� ���F�1�0�c���d|@�!�OV��a4���5W:�@2%�Q&�2 ��M
G��t��!W�����>4(l�5�#;8P�p关g �"=	E�͒�򉙱5C��ӣѽ�@�Ġ[�^K�cC��
?<�p���|�'�����6r�~�v�-x�����'�p� �� 1��� �cHLI�=Sߴbl�3p��p>!��W�&�t��Ϡ Y֝��L_}���%]		���?d���U-R�`~^� "D��C����)���թQ��2Ռ��3d�C�ɅK�V,iC�\
s�J6�t��C�IY�ra�2��R)�H�d0<��C�	(R�:��8|��4�WK�ES�C�	z$dL#'
%S�0{�^�F��C�I�p�~�Ce!ÚSd*4�U�_�nB�ɶ4ʤ�gC�&O����ۻ��B��]y��h�̟(w���	V�(C��5�(�H��׮��L]�C�:;�z���Q��I0�f�;p�C�)� ��IG�>!�	a�l���0�U"O�h���u�B�Sdk�!3�,) "O�8���Ӹ.x8Ѡ+@�C�"OP�� Ԡa3��:����虑�"Oڸca��4dtZ����qp<��1ODSf'P ������st4��'�Н����z���b�jX�7��(A�'��0�vX�E
ҩ�Q�3����/O!h��TE�Θ�ҋ�((��O��D����ł-5���#��MtX ��	.��8���"g��L��PX9Q`؄$�R�)5F��L�@Q�>�s�����I~�'žU)2�:A����f�
�� ��$�a׾<IR̝!K n�J��E�����L�\��ȓ+S͢Y�@,C�M��	���YB%�9|OzH����3M xZ#�H#J�
`�iq��#�&Jl���(V���	�A	�T����Uv���$d	?l�l���g�A�ȓ<��%ɧ�X��$qr!'Z9�E��+[�}z�����$x�%9�C�:��1%�Xc ���yW��)F��X5G�Vs�y{�$ְ>�DɆ���	��B(D����~�������z3��ܳ!a $FXpҥ�$�f��}��펒8��0�qM�68����qd�1O�.p��H�L@�吆Q>��(��n@,As�yy��"T�d��@VM	'mf�-BߓQ�^q�� �9	�zб���6��n�+O�xW��?:qqf_X��'vf4�RBͽ)�D�96�pV#��8�N�"E�_�*!�
����ST��I���YP�� kܾ�X��y�H(1c	V���bJ�oӠ�x�9��C�ڬ��=�tL��H�/6Qb��@�&^����.��㍉�~�� �	s�"�`��V+h�Ġx�MG�`�Oƨh��
�(O0���,��`��	�'��P*��'kh� G�Kޘ4��O���'��{�B���A��V����"O���d�[�T5�j��^E{���4z��::���>E��M'��QY��.Y��! N��yR�ۈ_�����^�V�����/]w��O�ÔlP.߸��B�b��7͝�w�T帖%;|Bm�����I�莥>���k5L7��#�L���T�sN/�O%Ò-T&�=��ӌH?�b�'�4Ѱ�� i}"�%l�I����?a<�y�� �y�(I8]1u� �ϖ,{�8jA����'.�9;Հ�R�Oߴ	��g. h���;S�ʉ	�'����o^A�iA�V��d��ʘ�H���DG��'L>� �EW�0ǆ�0fE8V��1��'@b��Ø,EQP��!O�HȀU�%d� (<��de5?��ORz�=�q��4?����㋈I��R�@��������"��	7W�L`�)�=*��G-�.a�q{�LD�B�
��	� ���A	۟f���@�� o`�Dx2��C�	�Y��YЃ�6��I�r����&�]�$i�UN��k)!��J1Hxʼ	&kϯ �����X�p�1O���a�ٙu�����ɕ�w���Rp�$\R���iY�%�!�#*�,0H���{���x�'ّ^�R	�b,B����2!�(#|�'�0�[���#<�|��%�^�+���'[�Uj��_�E��ē� R�3A����%�����d��|8�X���X�c�t}��R��)a��-LO:@���\U���q�':�����B��̨�%�
a��Ԃ	�'[2�[�M�K��.���z�O�O�H���*��.�~B"RV8M@�ꊿ_qv�+�MJ�<�4�
s�6#��6��� �HI�0�F��O.z$>�9p�ei�+	��xc&@"��d�ȓ^���ᇈ
*Q`B��X9b5�U� {����'"�*d�ݹ"�F�u퇀D�nlI�OR� ֫Z����uw�' ���e�ȟ���Vb�\*��ȔK�?D����'��DȀ����	"8&���F�z���؄(Y��Mc��Έ,2����C���O����Oͮ<�!�uY&�X4)��k6���,h ��"5h`C�-��E(��0c��)�Lޚb�Z`�@N�^��X(:}�e��w�M� ���'񈼀��K�/�R�A�W!�ޕAK<4È/%F���Fޑ��PSE_�C6��bbd�{�TE6}T0YX��J���m8b&�'�yb��b���ZF����h�8���5fЦK��4���B��|��`�N�To]�t	Ijj,�И~�4���h�w�юv�pah�dJ!�<�#B�%ӊ���|�8�*�I+@(� ��e:HX�u��(E����@ү
��fc�\�ܔz�H+��m� �I萒��u�fʂf���+�O pG⡅��61P [T�\+ku�B��J�"� ���&�I�=9����6|����Y�'V�\��ӝ	�	�=)�	3��Xea��]�as�Z[~��£I1���F��72�L��bǳ�<0�C�8i�vX��z����4�ӽKut\�f,W2B���L�4����'m�v����$6,����ܣ�ܸ�WE�!�d:ci�!��hͪzY�9RH�%��IQ����$HmXи"��F�p�
���b��+�O�ܘro B��J��%?beɵX�L}�8d��� ���r#הY�By�4@�*�+��'��|AЈU�w�6��BMڑҘH�@��S��5EBo�k@j`;⩂P�XAna����`'*G3G�2��)��`��1��c� t�x [d�ß��t�|(KD�#���r��T;�+M:5�� T#]`�4ht�T�� V�L���ݡ/�P�����Lr4 ��~BU�2[�db�F+g�=*ף�j�<	�'_*tz9bb V�_\ �ŉ�"&v��! 
x)����1^��J|�K�b�,�9�w�1�����ZC�Q�r��'"g����9�%���ՠ;܈���ˢ.��s�i�9uN%���Db��83�N���I-+M��a�͕?5�ȩf)�/z�?�(�,5P��@��[�9ޮ��#+��?�qZ5`7x0����j�*@z,��SoZg(<i��O7qnȵ�!��PK�E�gL~R#����ۄ��!b��vnM�t4�l����nM �����nx@����#�y�<j��R#\�u�r� �\>��aF��g3ƍs���W\u!���)� U�/8����6�ܱ�Ă�7�C�I��n��u�C�\3XS5�DY�LP+���Y]&T��T�V&L���ŷW�f�?�rH��M�Z��u����өD8�xza"�8s�[�M�=�2�I9fcX���&�>L�y�MZ8��;F5�O:h�rF�n�J���Y�}�؈p�x�ǟ3O��5�a�T�����+vt�='?��bG>U�𔻕�ܵi��(J�K%D� �]���R�X�!�:P��E�4���߾,��7m�@ �)���_�O��I����#�ׯ����$
�/c��B�		��T��C]�$p��j�24�7��K1�h���{�ĉ�Fx��xǊ����m:N�x���
8D��pb ۜ_�ax���(b���� �8D�LYV�=��r჎�Ge��[s�=D�ȣ�eO��Z�$*�k4�Lp��9D�p�"h�������`��82"$4D���sF���> a&�±Fl9���5D����mK^���Q�g^�  ����=D�L�f��?d���mߩK�2p�59D��Al��WN�h�`�_�y�!Ra
8D����&6�U�mV(ݢ|h��7D��rЉW�"BIsfg����1�0D�8�Uj 3��ǆK�0r�	��:D��i��Π.��]aWG�@2A�;D�D����1L�L�+Ғl���:D�l35N�!�)��R�=
��j-D�4Q7d��s��q��랰SV��-*D���K��#V�hX��_>�zչ��*D��چ��+CĲ��\69�|���-D�xh6��A dHSf�
$�~�i��+D���P� �9'J��G�H�>�>���c'D�dK�NJ�*�V���+!$�q��.D���PhI�M�����Z�e�wm/D�p����?�^(��̏I=��8ׄ*D��iE
�'
e�\�gMj�P�)D�h�p�˔&�>�[�$H�v�Z��&D����fהu N��b��:��)Am%D����#)��g���[}�("�#D� ��%��TZ��yK14�ɻ�l%D��Ы��^X�I����?��1�*O���⩝0B� �$R�D1`��"O>D�f��^ͬY��̤P�.p�g"Ob��(��J}��ؐn�}�ļ�"O��8炚+\T�	v팪l`:��"O���H�-�ࡈ��T^?ޝY�"OB���J2^��œu�T��5"O=*�X�3�MUw0�ٔ"O������!� K5L� 2��'>@p(�99�"�� ��(eg]�[�l(��9f̖�E"O (�u��F~���F8�<��"O��E����t�_誒"O�]�%��!�.l�cN�MO �q"O�Q���U�3�0���n��p@���"O�pS7�I�pz]`��ĵ76
E�s"O8� �k���x��n�@I���"O�<8��K�f�Ҳ��d#�,��"O�1�G�@$>�B|��]�j34uZE"O*�{b�8;fH��Q(2����"O�}�qbQ�(���q-ɱ H��0w"O$t8��� �얕R7�|��"O�c�.dI�T���j�\��"O���F��(Fu�4+V�p(����"O�hA�GQ�iU
L8��9G�`,��"O��vƜ'&���wAI
;��I1B"O ��0�_���0��Y
Hs�"O��0%�:/Oh	��[T��S�"O��:%�Y�d��! ��	Ur`"O�M��!�R!�׏�9C	.�s�"O�D��M�`�����װS�8 
�"ObP۰��o�V�(P�ԟ:���+%"O����eZk�4�[�E��Mn�#�"O�y5Y�ER��G�J�J���"O
��%`R��m(�#Xq@��"O�ï�9�
�P�@�>Cl�U""O�yՄZ0s:�ɇ��93OV���"O�}�JE'D.�3lݨjM�p��"O�;��@ 7:�P�vC��Jq"On]�G�,DD����b�2hR&"OL�aQĒ;{8L���"�4*�v"O,a�
�4X������9X���"��0��1I�b
9������UR�?4�M�T�H.h�DJ��T�'9<���O�(��i*��$�p�-O:ub�cW�HX�@�����g�Sv�v�����-ڰ(���9V:���OBAcP)�
> N��v��#��dㄳi�*$Y�Щ5^�1"ulϽ,p����dB�tPf��,ӲpI���'.װg &�Km&��Q��S�Ҳ�O;f��@:D	8X[��t�i��_[x�����	g�.�~+6,��'�$*��zu͗�wU�d��(O�O/��0�Z}Vi�
�9�f��d7@KЌ8ʓDM�h��yif�	�l1O�@�'H�����˔B�<X�o�9O����O4x�J<�"R"o�
�	�]g<4�3$��+�珀w�L���ōNE��+K�B��	ju/߄�\�Z$�D$=���?���|Q"kQ�S�����Vv���0���>�R��e5j��疱MM�)�� �I�'��Z�o"=/�*�JG�q�$�ȎE}&�<Y��d�."z���ꓱբM�E��1r�`� ��M I,>ǓO��5���r}�)p��ϟT"�
��<�ܬUǞbyR�ON�����<��u#��Q�H�`�u
�I��S>��]H ����#]��`zR!	�^���ǰ} �&KH�!�R���y&pxkCM�H2�P{T�*͸؏yZwH��./���AV2*:�mڃg��tC�D�!����(P���D\P3P�X6E
h,� ��ݣ�M�j�ö(��<�!.	w�	12HK}:1��8'�Ĝg��a�T�i�q�,P&R��Q�l�l�u`L<	���$"B�`Œ(���!Ħ� ��0K&*ԡ^<�R+Fd�˓�T?��'v�X�TO$]⑒�C��|�� �e���u��B�-	Y�t��s 9ʓ|�� �᧋�J�&ѫѧZ�!1���$DD��z5`_yb�G�P����d���ѯJ~��ѵ/��ٲ�������+��١��K�,��,Eyr�ذWW�ɛw��	�أ��[X�$���h��=9W�Z�z&�� �KS'����r�̑7e�$��O���[�dJ�,r<4tp�w�.��h�q�`�E�zl�UR�� [S(�>�T����I;.�}��C�u�����-ǘwվ�Wj6�	Xy�'��
Tm͉*�.a�5�M�oA��O2}Ӑ@��)B@�s��H�<e{�/�M��mZ*�~�����h���?�R`�۴��Y�r�_�?�2e�ٙm�%Rw��'"
�p�����{�N5W9r&��N��<����	��h�R�#��[���)8��@�r'�4/�(-:�F����dڽlR�5��؟vy;�>��W�-�v��h�_K~��!��+Sz��f�Ɏs��P�cُ?����e�O���L�9u �!B���L�*����Z18J$��U��#VKS#�b}�@U� �)��; %� +�+��s*��ϫg�p�'��8�dD�|/�Ty�P�nH?ɢ�'	�XM�������a冱I"B�z����'�.�(����7\�R8�4��P~B�U��D�`�#6d	SĥO5!�tR!�]��?aG.���O�{�t�\�M� na+�F�"�5AT��@������b�4=#��A3�q
PN���OZ�ݣ*�z]h��N��#Q�	
�TH�|R �)J�TJ�O��������������	�t`ʸ�� ��h��ԅZ{��W΍4D�$��D+��nT��bЌQx�D�(Q%tsraB��ѷ7�h'�`@��!�$A4�r�ɗw<i���[w	�=Y��6
%0B�H/L7K�<�B�ЂD���v��&Q�g˒�Gy Q,Ҽ*��mx�doN���N[,�#�' !��S��>�>Wʚ>\����Vj��]�yR�g�-1%����#�.%v���۳VzN��v�ˋ)]��#U�IIV�.׼����M^8�X�򤅞5K�	sSk�?e
�dA��Dw����E��'g�Lc`��

�� ��e�m��H'���QRTd0Lh-A�`���0n�'F��91��Ӏ@��ʃPrc�@��|2��SS���ڣ�rx``$,Y-Е
���4%K��S�,��I�v��([�Č�XU�a� ��VhJ�=�l�3��s���<p�� ��[≵Y��I��w<��pd΍=��b��4��Z����"/íDh$�ᮖ	��Щa��nx���g��9e̴f�N�A4F�	Aa��>6��1U�\�!��5@kԼP�����Ҽ;�.�~(�p
�j�u�4���QK�5��5���cl¸��O��c 
�V
L��աA���Äb��(O��M�
M���Ł[����O������k�0ĩ��#A���7�'P ����?E��X����z��$SZ���$W�1�숙@N�S���	e9z��bO�$2� ��Y�i���ˮm/�����o@2���cO%G��	v_�e�ɾ
n`۱��9=<�S�h��Ɍ_q�K�
\J� ����Y�b��q	1­i��*c?!�嬍	<�0$8��q�����"Fʹ��R�7��S#Č,0��=!����2�*I�4!G"Д�E�#�m��4i&�jE��R���#p#�	�V���c��I�u�6��Ǹə�NԦ&rT�c�C�{(�ȳu��1.����٩��tiV���T����K�=}��b���K�?y���Z�+L��~�hD2�����(��`i�.?eT)!���N=2+O��cT��$���u�'�B�9��� w�(�ш؟? �7�Ζ{K��f/2[���u�z����?I��j@�߬_ ��Co۝e��IS�x�U�&D�lB6��4Ͳ�O�m��&�j�(��8(�4#.��I���Ix��:��M�F$Vy^�՘E��3־��P��*�b��,�r�f�B��(su9��!h��� ���MAkށn'x�0 E��?�Db��p�E��{T�3/������41�A��\��"���>>����ݻ_�b�3��Ƀ�b�lQ�A���Jf�1p�ʍ<c�04ʜ=B�,�i2���~2�����1��AN�F�]s�nZ0��5'!^�9��T��'S���a��IqZ̧O�Y�D�V���?W\�p`)��D���v��-�z���e�-Cb���^�e����i�|9���E�}�9Ѷ��ɮ@���ՁA�4zT���(X�/q<������l�
�HOq��,AI�j��L@V�2O����"(�0 t����`H����iQ��)�`�j@@�(�6$�E�7h�1o�"Y�"8O�H��^�y�F=�v)"��V��!��l
za �h38H�� �"^˔px��̡z�F1���韪	��K�Q:�݃>fV�DېNS��J!��1JP�I�FY.d�b��	pFH4j�-��Mɯ�~�]�wJ�q#'mX�i�x�Z�@ԑJꨕ0aN����(�'"�UPC��)3�h�� �V�1�R���Y���_E��
��с�ԙ�Ч8�>�Y7��Z.<Z�I^��\��'���0��РH��M�V�C<	�ƭ��Ol�{Ӄ�G��`£J]�	u�|K���s���9Ѐ$8���[x��"��A���<��4H-+bB��+<���ț}��`�u�Őf�t)�F+�0{�xGy�'=w�ac�!ga��% n!�d��V�&��]��qBr��H��l!�y*�X�� ��f�@�@)
�tR���ǃ�80��a�KQ��)�[�R���ϒ�;� ���
�� ��䆝Yʸ)�W�� 4R��7�:|O�B'(E�?� ��L\o+�Y�T
v2�0�PMS�_��Ē  R��E���*���r�����<(��Z�h�È�r^V�	�V�HRnMR�(R��d��'?��.A>�?�D#D�|����A�M"q�9?A��W4��8E�;I�օZ�m@�I+6�	 4|D�!^����,{��'k6d�A-�e(DE�צM��q0�nS�ZTr�Y�JD/�zl�P�'�0<�&���6ЙI�
	,<�\�̖�,8i���T.���'(�%�?�g��|J�lԉ7Pt��%@��J�*=gN�DNF��>�G2��A�qf� ŸO�h]#v�P��( ZG+��<\�:Ղ�5"'
���2�)ZC#Ѹ|�\�8YcW��`#�'5i��x$-��	&�hX@
v��qP���Rҙ�d
��b>�D�*@�P���"Gd��gK�e	^M�sd�}z�d��=6�0�O��[��<���⮎!a+�����N�~&xBOM�an�$�������!��>�|{bGX�	# -��'��i'�e0��'����4
�k�b9F{�`�)-�̵P�噝?�����	d9�V��#i�I��r,�I~��'��\�,ɤ�k�i�La���F�T�[@,A	�蹡��;zMc���=HT�YD$Q!I�-@���出
�й�ðq>��d�~���OM%)h�l���tc<}�i�_�i�g��q+ ǐ�!J��	��X9�s���B������W(���0O�'v��h��̩<Fp9�&X�h�`]x�'
��[M�����VEmխ�>��Zx�m�sbD�+�H�ӧT� �H�I>�ѧ\�9H h��OF4���~��ʄ/w�py׍Ĵ��� ��M�vO�7]HM���DA�eA��� ��0���u���KGE�G�n�#�Q�*#X�%�>?y�G���H���4n�(i�,�0����
�~y� ��A�Q�x�f�),�2����J7~x��<A��Z?���r�,7 $�͟>t��U�Q+�1�.�3aT��]_=r���S� %�ŏ4.�t���� 	���z	�df�0i�hb�cW{����ҭ� ��O:���Ԯ�B���4AѢё�'�=@�p���
1l�|�' �"���5"X4��" Jz������0W(���G�:D8�)4Ŕ=p$��>}2��-P�)���-ݘO�>	�u�hќ�:@_�.�-(�l���Y�S��H��'t��:R-А	� -�0���tP�FW�C����R~��Ǫ6�-�	p��M^�>���K��\�< �O�W߱Q[� fcF������5���a��O�:�H��M�A[��9?)q.�Y�<��
��lt@��<���b�_	:�F�!E���1t6�F}�C�V^����c�(2�h�Ek|yT����NV�@��gIɶF�(�1���M~�ǂ�-xP2g�ǅ[�ݫĢ(�OT���K�E�"�ud�@��}x��O*-���cc^�2��3e��Q�����ḑW�T���K%�X��J_�l�.�*����RFG�</����'�L�QA�4c�D�H��DD�:��.u�aB5�B�yB@\�#jL�SE�6t��s��]0�DI��	\����aOќOR���Y� �Ĉ�Q��w�.)���(#�ɫ�O�95j�{��2nyn�3�|��.�n�1É�*p���W��
o�Ś%`�H����Â�.��L�㉠1x"�a��>yg'��M�p�	w��(�Ȁ�}�
O��;UD�!{�J�i��5#����!4�L5�U��ENl����	���.��f5������-�ԝ�')�����IVk�s���K��8B�>Z�a���G�*m��&��a�a{b)���9�'O�4N?��RjD����~r�'�%���5�^��!�p�^�;�C�E���p>qVI6mb�Dr��/s�(��G�7�U�ȡx�R� vtA)���=��Z�����#�o��՚%/V�r���A�G%Sl�|�4'"��"՘!'F�2~��C�O�]ð/C�d�WD��DL�SA�,.=ɡ`.�9x�8]x�KѼx�i����)1��Ox4+r�2&���Ճ�L��3�G�b� AeJؙ�H("T��|khi��r�	2����ӱvs�0�P�
y�(�ہ�
q�xi3�#He��]����en�zD��(BU�Ca2��폽n���dX�b�P�:�O��0��.�.ØlQ���|yx���(^bMѕmU�A����$ˊB�ء�'�!%؀)����;m�I��M�h��AP�Sٳ`� ��0��eX�(����<	���D��} șiW _�\��lP��]��|2	A+dR�:[xP���=$ޘ��A,9�fģ�m�'_��aDꝙKŐg`V�?�>i����7J��%I�U�����0>I����x]�h���/!O�U�&-�n�����Y�r����LL���?Yq�B�M���%�`�p���fE_�<���&�l]��K�T#���DC[�<�S�z���g�5J<�u��AA�<�� 
�2g��96@�0Й�C�U�<�0�Z�\���Е2�(�QJ�F�<��*�#J��PP��-V
���V��B�<a �ǋ`��e��F������d�I�<�Q�°\T��f`�NoF�a�H�H�<iUKH��
���(�o ̐q���<����t_��"�^�T�)V�D�<���͗Bw�@�����J�P1���<��(K�)�B���%P��E9�Q�<a�'A'n��F���J�~		g�r�<��#�9��P�ď�}�,���m�<�EM�C��;��7mv���e�<��=��	�0�+�T `+Ո%�!���U�Nu�"� ���TJ�&b�!�ܥZ�Y@l^7
�q��Lj�!��xd�	���b:�P�H<!���FD:��bZZJ�(�"O�@s!�D�5MS��j��^��Q�sA��KV!�d�1'������/��eb
 >h�!�ڂ(_�kG痐d�^��!	��!��b&ŋQ��:X�ĕIӇ@�=�!�������r������-P-dQ!�d�0���aS�I,gα�e�W>�!�$�GL`<�WD�<�B�膷{�!�DI�M��� ���w*@����$=�!��**>}�A��7R����h�!�� �̣s�"�haeN¬<��p�"O����=��e�A.�06iB$"O&1�F�#����e-�N�l��"O蔛࡝�I[r��1OԾN���(�"O�A���٦�T��lާ%�6P��"O~TS��Z"9�~ّ���$B��QCf"O��jgoK�{�"'��z�� �"ON�rw
2`5�-+�k��gv�#"O``%�-�D@�j�''`0� "O��jWˍ[c���^wW�U��"OtX+ֈԾyQ�1����,gKH�� "OhAh2��.�L	 3D�a1���"Ov���fJ�b_�#äȇ .jc$"Ot�R����u�����T�
'��H0"Ox	��#V(H,E�5����a"O�$8Q�.`+����nrf00�"O���wl��.��A��_8�=c�"O�\�@�	0	�.�%�ڮp!��;S"Ol�yul��č;R!�,!���"O*	r^:_dJuӤ�W�a���'"O���!�֒=Ŋ��ӄ�5�RןU�<a��KY!\�C���)`r�9�NQT�<I�G]*b��U�0�)Pn6(���k�<�1MD*;�rA� )��	�L9r
�B�<1��ߴ�T�"Q%�	%9��ShB�<1Qʍ�:��Xf�D,M�}@pHRW�<񠤒=+�ժ�gW/�b�*��U�<�b��<6���)o�b��7��G�<9#�	�W4��4��+anN�;�N}�<���ж*���b��� z�Lv�<9�\*o|b%���D;�}p�Bt�<�ϐ�aƆM�@�K�,�� H��C�	�>�\% v��%���5&�!EdC��6�4����$q����M�S\BC�ɵ;`�<�S+ϔJ8��ر�"n��C�	�	���*���&`?�Ūf(θ4�C�ɍ.��څ��4�4mL�	�C䉏 ����T+�wnT�K8:B��1Dڄ��p�7g0��Q�KX�\�TB�ɂO6<�,U,Ss�h��$+t�bC䉷\�H�eù(Ȫ�ZvF�UTC�ɽ�N	�"(�+.����E��Dp�C��-*_:]��ɜ�/CT<3��
;��C�	6���(X�0�>�0 ����dB�	<t�����D7��� ��GDA4B䉟;�D@+����xz�<	�ʆa:C䉣l3��eH�]�tz�I�(�(C�Ip)|�a�eZ8U(��R�ˣY�B�I=&��Ir0�K�W��u� 쉭?v�B䉲"��e+u�J�)|��@���K	�C�	�`BNC��]1V!���̙F��C�	=G�t�ꒀ��`��i����SB�I�n��Wț�G��%3�e��s$�B��4*N��B�.ǰ�pU���@"ELC�I1fd��ȏ@0p�����rC�0C�Th����'d���"UL��C�C��%x|��نDuKn����DB�	t&Ũ�"�]��(J�Ö<Q��B�ɻ&y�h#P����DH!���{z�B�I{��,��Ӝ[u��2�kCr�C�	Y^l�#�W�&lm2u�ߐf��C��;���FB܊@aTDB�p��C䉓ST�����A)v�(I�� *$ B�	�~���1��9Aⱊ��X"��C�)� 0 �sʞ6Nt�%�X,�B`E"O���g	�$ +r�8��
��t�"Ox��ƛ�#���#���(���	�"O(j�J�)c5��+P*��=�U"O��a�̖�����J !�*M�G"O i�􄆻3C�i�cKU	k}� �"Ojy�e�I-1���Z��*q��"O�B�C�[De0���?,����"O�� TD��C��h��G/G��Ma�"Op vc�s���w�Ȼ6�l��"O܍�"�X���Ѧ��5KԴ���"O.L�V��  �Di���3���)�"O��J�;>�@#.��+F��{U"O��ۀB�r��,�Af f&Դ�"Oީ(���)����ЦV�"m�e��"Ol���M��C��a��[�Cc��0"O�xР �6|��A��W��I�"O�
���*�ۆLG��8%*�"O�p�c܆g"R���K	�-�2�K3"O��
�
P����Eʀ*cyY�s"O��ңBhܰXE�K�jk*��T"O��/_�
��AP���54�Ã"O�p�F.V��Ic�P>� 4��"O��:�˗Z)v���ʠ}Ӫx�"OP`a�)� �%R�ZĪ<��"O�1�nG�n��x��(0��%h�"O$"�b��S@"��ǎ�w�P�+G"O�	C(C'?=�b�>��u:T"OE��
�A�P4Sk�7��h(p"O<Uzł�JRB(9�	/v$P��"O����gIQ�D(�E \Gc��"O��'#+d�@�
S:X@�"O<�s��Ұ ����$��	4����P"O�$)$AP��r��C��2�nyd"ONl
�h[�.��mq��	b�UI�"O�z�@�K�fL��NU q�4U��"O���A�"��ؔ-�� ��!;�"O\�
`G{0���Q�\hw0 2�"O�����k��$"�+��ap$Ʉ"O�I��
nM$��eT9D|)��"O���U�HxK���b�49�ah4"O�2��!6�`�K�"I�O�12�"O�T���VX���@���p6́�"Oژ#��C?x\*2�V S<8� �"O��
 ���_�L�Λ�B7XL0�"O:p�n)]�Ʉ�_�J�"OdrnɖRHY��>�XS"Oj`1�NW?nl�&�Y��l�V"O~��GC�.�r��!�
u���"O���Ɏ�F����&T/!Xj�[""O���ґ99��z��Q�6=���e"O&��B�L��	[rH��j:��%"O:��fB�L�Lћ���?�0���"O"��SFY%���q&מj�j��"O!��뜈S(������d��y5"OJ�`�♙p���E����e�"O�Dr4I��[�*A�Ц�|(q��"OʡyԩC���E2k��c�	+�"O�@{��@:-��ܫ&!�[趼�"Ox�rM۽wl�i#�[�Xӄ`A"O�G'�$L}��j��%Qo$�"O��9��;+F��a�AP�]+�"O�q0G��L�8i�5m�g��`P"O��iUL�D.�9�N�>0�e��"O� rD�6k��")
T���Xv+rP""O�mIQ��#�
�Q������"O����S]t���燣q����f"O*m��%�f�Pm�@�u�6"O�:�!�!���Ib2iyc"OQ���i0(r��}1���""O@�`1��J�-#��2(�.C�"O�<1 掩2P�9�1@zȰ�"O��H�	̓Bu��@�z���"O���dh�9D�^y��Đry
���"Od�R�N�*zQru$� ��-"O�e�P�ձ~h�� �: @n)��"O<{0��6]�x��OՐD/��)""Oց���UC��-z��@- ���"O��f$M�*$D��L��r>ͱ�'�(%r5���3(�H=b4o��a����ȓ.�2Ay��M3�Q�jm���Ey��|j5�BS�̠�Т��A�p�C/�\�<Q�̚X� y�C�:�g�[X�<q�=?>l�{U�u�-;5D�z�<a��ң�4�t�%fѴis%�Ot�<A���� ��9�"u=hH;�\y�<����J�Ȇ'��j4��`�Wv�<!7�Hl5N�A�!�9��6���yBh�L��x{�ʐdaHA�'a��y��$+I<��sM/3"�HxdI	 �yZx��'
�*0���r/�A2��'����Eș�ϔ�#�R5V��x�'���)B�ɚv�mQ���US�'=������s�8c��:�T��'G�A2@{�^YsQ�Jr���
�'�>`�f+_�L4ԡ�p-��l���	�'ͦ�(ueO;}��x���w���8
�'H�m��I0 6<�A��_�v8�4�	�'�ę&�H�M���L�(�,�s�'��Y�w�W�_}����O �l(	�'[��Ҁ�%=,���ϊ1jly�'�VB��ͺlpZ%���	�vĢ�'px��VH�3v��Y�#� J�}p�')�}����<:�@yc�֝y����'��鸵��2@N�x�ReF
"�؜X�'� �9R�(nd4K�c� �R4+�'��	RP�ǏX4�;�G�&P9`�'�Xp��L�o�&�ZQG�&�)�'VMk��%��Q���H{�i��S@T��(�|���� �ȓJ\��L��v��0�� � ɇ�r��a�b�B�UDih�U�x-�ȓ�� �@ܫv0.�p"�ތ7�=��^�jh�E�Z1Z�E�T:C�&+�8|C!��JDi��KP�9qBC��*�B��AD�<`��t0#�	�B^C�Ib+�5��hPP���e�;��B�I�wy�����g�T<2T
	'g_�B�I�/r��Zƍ�z���P0oS�*!bB��fռ�BJəS�;玏:PB�$ȼ�y�q��c�*RC�	 e90�(��/,���1xC�	�~�茊��<�Bp�&���]K\C��#3 -:gj�
w�$pc�d IC��!V�jԁ���	��1�f�6e�B��' ܾ�4��?9���Y殞�/ָB�I�p�Uôbʄa'�t�Ѓ�.KzB�	�=��1�c�'� t��l� �bB�)� ^H���D�*<�x�J/$����"O��V.V!^Er��l�&2���:2"O�I��Iʴ�Z�L 3d��!"ON=�!'
�s����>X``"O����I�2J�zF�$��t
�"O0is"&H#N�у�X:?��1�"O޼PhH(=�$������8E��"O6lٱ�9:���kC N�l����V"OB���ϛ8��XCBQ7!��xW"Or!*�Z`EJq��;m���"O�u��H�@��$~�`�"O,�9� �1[���4/Ϧ}z&l;!"O*�I��>vm�mZ��.b^�9"O�-R�f��A��t�GLB)}J�ux"ON��E���tTZ�KU!]Mnt�V"O����̄!iP�I��=c: i�"O:� %	�7d�Y$�Ӂ�J-��"O m ƌ�X�B�R09�^Tc�"O֠�&�[���T��g�(��� "OR%�Gθl.��G ��+��[b"O��{��;�n�\ش�7"O�0�`�K�	����P͙� ��mq�"OV���.�3-q<Y+�̀�y}j]��"O��R��!ϖ�����Dm�"O��!4�Y:���3��Щ�(,�b"O�,(�EH�J���� Ĥ(�����"O@��!P�}[��)$&֛ey=�U"O��R��C���꙽s_l<�"O6�A��z'�`;���&lC���"O�D+�MȄ �ڨA2�C'?-�4�D"OYI��S�!�Ȫ�/Z�|/(�c"O��ۡ���& �\�N�Y[C"O M���B*G}vU@�`���$�G"O0���S"]��� �J
���"S"O�U
�K�oct� W�1]��Iy�"O���ć2v����AI�r�u�$"O��'��8X���X#k��ecJ1J "OTh�S�WD�"I�ӊ@ ,Thu��"OԨr�	HA�Dp���̑RQ@��"OV	HRM̜i�z�`��Мw&hؘ�"O�T`2+?8� -xP��1�(��"O������l���@'Lz,Y��"Op��T/�>j���Q��V&]4�Y "O�`7Hлw�4�c��ٵQ��Q���7|O��{R,� �n`ҭ���n�*�"O�\��ɅW������N�2�q�'���[��ɇ ���oB'm���'4��y�.�2FH�d��;�
���'�D|;$�
렡b��Ai(�1�'�<��P ��di��I���Y����'��pB�߰��$�v��R��'EB���톕�huٵB)~}�`s�'��ɢ���C^���M�}��᠋�d�0|����H�t	��:~K2����\�<)�M[�F��A`��2.��!7H�Z�<��B0h�@�`'�Ʊz�����HMp�<�t�1W����6&�84��4p�mAT�<���LDJE*�ĕ�;��l�Ԃ�M؞D�=���4KJ*�߸(M���R�Np�<� C���T��a7!0��,Ep�l���O���'K��	�b$@��
Q��'�f�W�L!T���������q��'hʑ�SL�--��aL���.	�y��)�S�r>8��$aN��#3n��C�)� V��C`~�&����4��"O>�؅.̘SQ.}1���=�5�b"O��@�O�3�� c�9!�ٹD"O���C� ��۶�%rs�P�"O`	�I��?[� J�O�$s�-�y���	,�K���zx|�������yB����v8�b̬k�@d�䣘"�y" P�A��Q��;��y4D�5�yB�!ݶ5���
) �N�a )J��y2��J���"��F����F%�y�G�;r�)	&�G�;�h�w� ��y���p�c��CJ�&awΌ��y"���l ����H�@`��m��ykL`�.�zp�SG2Ƞ��F�yra E��RbH�5=���F� �y��
;R�`�o�3��=@����y�'�'q@5��O�;�8B��P��y�ƙ�I��a��ۧ8O��d���x��'�2)1�K�S�eP�#�+s���'�
d���� �"��f����	�'"���|�)HrgM�X��3�'���̔�Ld@�@Bȡ_:-�'��?�y2,
�^�����-�#[�y�K4b�,�[�lN�ʲ��0&��y�nү~p�d���ދ9߰���V�0=��l��%���k��7���qB �yB��
jNV��F"с%�B�P�,Ϯ�yRM�?r7�8g�9	����>�yb�N��P1c��z�H8"�k*�yB�Νd�h���m�1��䝠�yjK4D|	�#��]�`q ��*�y2gB&�e(3�EY���䎳�y"Ƒ�7!�d�� ��`��2B�yb�ܻ3T��1l�Y/��B�c�7�y�į,�l,cU�S�W[�@[Wj1�y"!Z6��};A W*UNXe�a��yBL�SRҐ��g	�#�����̿�yRCҨ��T"�'Ђ��DP�2�y�j��ao�ݩD��_t<�W�V"�y��CD����	��*bgF�'�y���|�����/δu�$�O��y2�č)LB}��(��t� �����y�T-X���(�i��d8ņ��x��'�r�C�l�.�����Q! ���'�F����ƼEiv!r��ܦ�H��'��@q�2t��������z�'��0�E��F6A��+��E�D��4�hO?7� n�6��M±H�T�ې@�~�!�@;.�vĀ���*��7@�<{�!��^P~ܡ[�ʯ84��d�
�qm!�dNp$u����:����O�Ar!�d΁8��IA���4x�ԛ���p`�y��d�R]�,�	Yw�UsVjW$=��B�	�)_���!JA1i���zlS*l��B�7#���Pu'\���fеuC�##IX�:Ƣ%vZ$��gD٨�C�	�Tމr�~�ԭZ��Ľ3&�C�/��EqdǙ�G˦}zqE�@��B�I�N��`P���=m͞�ef�
��B��8*�fM��Å�q3�ó��R�B��$#��):7�vo�����]�lɼB�	7s�X������z�k񨉯!L�C�1W<l  �݅6�y�WF	�,�vB�I�l��Kӊ\< @�a��)��`�,C�)� <�A�MK>t�����S�\��Ott�wCҹ#��z4�ضT�*t8FCG_�<�d�O��<�*a��/�F,���[�<!S��('`ăf� +y�48�	T�<Q#�L-x�����M�(lʬl�	O̓Y���b>2�-�".-P����P$0�2�R��%D�t���V�Z�:� @L�1z�ָ��g9ʓ��<�G��4d:�ò�J:\�Q�(�n�<�)Ï:f.́�ʝWW���Νk���0=!��P/Vg��Ц�-%�����AA�<�b� :cJ�I#ɐ�)�m�RaKz�<��	�ERd,z!�AI"��㑠�v�<)���5od�����d��� &K�<�0�/�$��B�W�_\	�a�D�<��"�����:ag\m�ݒ���\�<	��E�"��Q3RJ�'c��2cV�<���l�6I��3-V�U�
U�<�rɁ"6��谆\F�%PS��M�<��-$����R�q�J�<��"�f��͡�E��G��,�K�<y@���:���XP�@a'�P�/�G����&�:���+ʽ4a�2F$G%�P�ȓk�*�*���s?�D(�휋5b(�ȓ��XuES�!n,pa�]K���[�V(A5 �{At�����A��F�Y��E ~=e��a<�Ņ�?�\Y���;d�Xb� ��I�H��ȓn��*��B:��T*h�>0�̱��W(>����;4�����EJ���ȓ8e��#w���/�X������ ����Qybd�%dM؄^(i�n$�J$�y��\&E�N�:�_�szi�CQ���d:�S�O5� ����$�2(P�l�<�XC��3x��I"'�K
%�ʕ��E$C�I=k��)PK�2�����ߖ3C�I��Ze3���%j�2��#��"�C�ɾ���cX1^LN�j�FH?p�>���I��t|�
����s�򰨵�˶/!�d�
��P��R�^��sa
k9!��P�V��-K�M2{l���Mb|!�D������7T��P'�^Kb!�Dń@0��6�N�V4�%�6+IGS!��\�N�*�Ať�f��1JM�&!�$�4b!1��^��ɻ�iØ�!��ݚp�x�#'��}����"Z!��-�>Y3�$�9��}ze�O!���1%x8�@D@� �V]�) cM!�d2XXP2l�/|.ţBG��^2!�ޒE�l���,X�HPR4��'k�$X%�
e�ڸ�� �Mkj��'��X�	�$��Ѧ�PU�0��'Ϡy*ҍ�vĔ�cQ��s�(H��'x,��7�%�.p0���r��:
�'�=
����:D���Pm!a6��;�'�d�����DHsFń�0`2��A�<��G�e;��"Չ٫4X5V�Q{�<9���SҌE�sE٥��uzss�<��K�s"�����Z93Dz�QFUg�<aw̚�|K|I#dT�' �a�PN�<Q쒩(�������o,��l�H�<a�&��WX�궠�#ǈY�E�\�<I&�Ӓbh��F�!$��j� Z\�<Y ��b��]0�"f����`A�<��H�$2y�7鄴5OL�f���y
� ���s%�'���r2#_j�	Q@"O(t���Q�&��L�aʆR��q "O�\�	����`�lVL�0"O�r���*[�X�r�� a ��"O�Gd݇`����MDdUR$"OB�3"c�$0�UC��nf5i`"OA� ��U�(AV�ۯ\�PuH�"O�!��G�b��귢��%ӎ�B�'�0��1U�"�x0õZ� H)
�'�������^x8�k�%��Qj<�	�'���v-��3�6�q��	s
hę�'��ᨖ�ұz�����V6g�*Q��'���#$�E)%xh���C�\���:�'P�� ��#9e��{�O��JfB�Z�'�� Z�7Qj@����DHBy��'��Q��!'��D�G�H�,8A�'����r(�L����)H�@�`M�
�'9J��a��0bO����jh�dY	�'8�A���D�o=��2�@�cy��R
�'��J�Sl.
qA�a��� �'��u�����tj@� *j@Vps�'sh�Q�ǍK��{�Y�dc�;�'�I�P��a5(4b����)�'�"8ys�+E2l�`�+��'��mR�k��G����éP�X�1�'jV�j�.�5@� �����4Q�����'�1!5&۸f��0�B$Cn����'�B@�"*����bU�)E�)��'��
b�-&X�`���+�`{�'R�K��J�g �i�1�E��~�i
�'���+�#1C��Y
�.� 
�'�Z���ǥg7�����82Ĩ��'�4QR�@��بg�k�x�'gNpy����|�� �VjL�/��b	�'��kg%Qy�8��j�/Bh	�'?H�$	R�g��@���\����'���*�)ET����	6z�'��1GT���cD�V�
��'�±�ef��z�n`��ΒH�ֱ�'nr0��LJq�y9p�с<�b$�
�'F����F.]\���rcԅ-�l��
�'���KtꞆ�\�3��\?� R
�'��أ�	6[�b	"cY�T{	�'���H�M�#��<��I�������'�E��˱kP  �F�%/h9*�'��!ء�U���U:5�%7���'�pE3�x��eF"R���sv�j�<�U㆛1OF�gB���%���i�<��(Փ.�B�S5'�N��aI��c�<���\�P�bM:$rRY��/D�0;��M�Y�hI
!
����� D�Xy �r����5����gD!D�do�Zc�t煣9���*��,D�h8��$D>|�#�0f�� Ԍ>D�H���8C��(�f��Q8D�P�q'�-J�|��0��0|i�D�l4D���a�
�{��}��Fэ$G�L� D��K甋@<�p�a�O5!������3D����G�&��ihT�>_\�9H��0D��chQ!NP���營r��Y��L-D��ѥ�S.8ܜ�V
S7>��1!�,+D�d�0
�X����9u�y�*D�����O���}C��R�}�y��#(D� ���D:y)�d��폠>�,0�գ'D�� �ݓ�I��O�
mӧ(+nu�ȓA5&1QG�@�dKR���Rl��ȓP��hrE 7��2�A�����G֔
����8�R��B CD���B/<�Q��56�x�٤�*n݄�!mZ����`t�	�L64�����h�!��Q�snN���3ZL���ȓ4�Գ�
�tnHL��b�-sմՇȓ��A�3	FQA�l����M�T ��I�tP�E�;}=t�&¤hUص��	�����O�B) �"#�(9���eH��Pu�r	�'��Z�ڕ��<B(Yr�#��`��H�G��$�hm��,c���� �p��(KE��8�ȓ�B�����o�9X��M�Z�,\��,�jm�5���?����ʊ<1��l��Mm(���đM��[�
�t�0��s�|�� �/i;����y�ȓW�J%I #EH6j ����5��A(![z��3���`%4=��.�k��@,�[��Ȩ7	�لȓe1+����b��ާ_�~��H���F���ZJ�y ����ȓn�DC��H�Rz0%��v�:��ȓFE�y�Ec�s�ެ��Kd����42�L12J�0<2J��a�]���}��!�xtq)��Ъ�˱�� &��$�ȓ=���Q1"E+w��I��3�֙���n9�%�o���{�.�'�]�ȓcL�{��%�=c�A��;�|M�ȓ�H�ƈ�"���:���%������ʃ�T�=�l
�IΉ|H���=�^Y�	²j*��k♄�}��@�@��N�f r!L�=@R �ȓ$�-�ҩ�-g�f�Gn�0�|��+��X9�웂L�����gqX-�ȓ�� �E� Wt�����&�F��ȓ&�xD�Ju���A��8Y.���<.8�z6`�a�������p�ڕ�ȓ;jd�e�U��yr���3%�H��q͊ܚ�v\
��Φ+����ȓ|'��pR��jj�Y:�jȮ"����ȓ)U��!��@\b�xvE�h��؄ȓ=�^Њ��ӽHQ�HЄnQ.4B��ȓX*���(@�Ql�1`�!�(#{2���;뤥2��$>U���_b�<���^�`I����'d�۠��\��M��3@���ǣ)z��T�mS=�H ���XpX���� �V��Cȅ�tp.���pez�h�a�V����Q�X�ȓ!rʼ;����Q��t����n��ȓ7@��a�4y2�˄�أj�88��(f�3�ls E�U�R��'���J��V*�dX�# �:Uz�'��8�!��W��daNR�`�,%��'��A�Sđ��d���K�qd�'���I�"*��3숎
����'��9�.��R�SR��9\�+�'���!���(�~X!'���=��'��3�o�yzj�R׉R��P�y�'�
��2L'rVd�,����'�rc�F*U$|Ph�� 
@r
�'� �07��N_tH�ʗ�Qr�M�	�'�������S1①�@Y���� �p*S&ZY �y�/Z�-��A#t"O������+D�j99�)B)a|�T"Ov9�1A#,P�A��&�~�#"O"I�v!� sC��`�2<@�"O^��aL��K�$�pcФ9�=��"O��auD��a"t��1�D�7�5��"Ol|V)���8E���D�E��,x�"O�$�F�h�*�q���~�I"O"�0ŀܚ@��ѡ�$̳'x����"O�8���7�&��I"LҬ�G"OPy��C��`)a��
<+�j�s"Oܸrd*ҷ(��Xr�!P���*�"O�����K}z��$� ^�<�"Oy��aS����N�aVr�'ąg�<Ae�.|���5GD�d\y�"A�a�<���)eS�q6 :Bu�H��T^�<9����V| r��:c�JPB���d�<����=�8m�"�7}�J�.Dc�<a??2-���$��@��k�a�<ه�6_�1���M8g_����It�<���<K�<aʑ��l@R�"�Vn�<A��ؤ�����'q#�x%�_�<Q���(1�I�+U�~H#�+]�<�M�QÂ�cW'S�
)२�,�X�<�7�>�t����t]pt�W�<Y�D�""�� ���0hz"�!�
P�<�!�Ҽ}��R��+7���5�H�<A 	��læ�*�'M*s���AK�<9����Y�3a�_a��:��l�<�ekܭBz���H�+f�5��E�h�<	q��H�([-i�1�F�e�<�n���A+[�BeA�͍|�<A%�d(s�AߧR�`�Sac�v�<�G�ѕCƸ(G,�*G�
�j�Gr�<9���8�v塤�ώw�r	�q�<9��+��U9���Q�r�	�	l�<q$�=y�T��5����dNk�<���7a����a
1�$���d�<9�쇚O�݀WjE9���P`�<)� �qp	��
G��|�W%T�<iC�ʻG��`守>Bu�G��S�<��ƕ {NA�n	0gl����g�<!d�R	cQ� �P�"�E�s�Gb�< �	 ��U� ̩z�ap�o�S�<Q�<�B�bca�<?��5XG�H�<Yg�]�(�\ɚ��y����%MH�<�R�uB\�0�/ⲝ���DA�<ib�Ox}�X�F��u���a�B�<��*��*�,����=nP�1Ò��V�<)�る��9���#s���S��m�<��Q�z�м0t�@Q�����Wm�<AA�R�=�Z��E{�.AU%f�<�W)�.��MHs�@�3�B�b��F�<IFRG�ni�nڢiz�t����v�<ITL�H0�����a��P��_o�<A3�L�ԸM`�ɚ�� �Ū��<A�kZ�&M�a�T�I	k��Ab�Sc�<Qp!^
�]Xv��sR�����[�<i�HX�(��7�9x8J�Q�<)wb݋��ձ#����ȇA�<qP�ιP�z��͙=(~��� @�<����/{���#A�2N<*���}�<i�Ɣ�(���C;��Ң�r�<�'��B8�9g�ܵvH(�)X�<� b51��S8�, t�U*`�*�"OH�9e\1y��Sl�&#^t��@"OJ)�q�N,;����R%-$�ѣS"Of�{H�v�^ek��L�vPP��"O�hf�B�f�\����P�2�ٚv"O����	�8m0 ���DF� � ��v"Od�R�\��9�T��vܰ#"OT ��aվ5`<�D"S�f��0R�"Op)��)AnJ�ٷ�ׁjtF�1�"O��R�.�a#�a����2Y>�"O�5P��
�_#�����&p`ąH�"O"���۞5��88��\D����"O>qA��'H�D�E�M���"OT0i��۾y~�u���Z��y٣"O��+V3{	$p�
��Q�@}�5"O\홗��g~��h�`a(�Ȓ"Op�'56)V��7FǬD7@��F"O�u���9�����_ 
���"O�ES-�!<�ba���=Y�e�D"O�݈�MA�X�xR�&�$��"O`PBJ@r��J՘ �"���"O��
 ��\�yQ6��I�Tq��"Ob}�&ы����G�Ч�f�"OZ$��L��Tf���Ȁ5�Nu_�B�ɮjWy�ѯ"a���P�FԡY��B䉯�q����6z���2���PAzB�	�#��=���JkJ�)�R�8�BB�	�!�Y�Ï��r4�,QA&B�I�9M��aݜ��a�%-�@B�I�~�܂���;Jr�%U�Q�4w�C�	/)7bXK�� �n�;()�C䉵{k@8!A#��@	vY���>!�C�	
TNL��5.�[�Xh��W�T��C䉚N�4��fbB'E�r��� �?��C�I�s۶9�H�)
\��JS��0�B�ɒ��	#���" �Y96`B�EhR��S��8|\��%�8B�j7Z�*Eq�^}iUȜ5xB�I�*આi˘	�.!�& 4gCNC�I�NȦ-P�b<��C�%
B䉟X� 4f2oW0�p��<��B�I�D@`�'"�!Ѿe`��;-XB�	-_%��q�8)�-�J�7l7�C�Ɋ3�P �S��R&�	b7����C�	=W���O�Q=��"�f?b�C�I�k��`-��y2s�A�#&�bB䉷08%�bI��Rq>�:���8u>B�I3AȪ�.���qˌe>F5(�C D�<+�ϱ3d��	� �0�!�<D��33d�
jdlc���(�*E�do9D�X0�ׁ<���[W+	�6F�]� )-D�8ڧlG"N���4F[�u��D+D��K�B�(3�r`�A�+3�x��?D�0�⁉Z���Ý�*D-AFJ>D�@�)�!,y5X��	_%JuC'D���&F�M�v����:N
Q0�� D�xp��˕4]� �J�w��ds��>D�P!$O������.H�x�X��>D�<SV�3m��C4�D�^(n�xtJ)D� ���;C/j��Ň�D�P���'D���PZ�雧	H��&�2�3D�2P�ظj6���Ơ��p��!s�-2D��Z�N��_���dA38��2V�/D�[姂^}"��3�
.����� D�� t���k�)�J���I#!Ԥ�6"OV�:Q���#���6"y��"O�iXg�]�x�ua��Z�O�P�("O���c>`��ˢ��opv��2"O��Pb��q
��/IUJI��"OF�B�ɏO-� �`m��"O4����7'9�T��&��p#���"O�H%��j�DQ3� �X���[�"O\�1p� 0I������J 'ަM��"O<T�aO�{��h��L�e/҅S�"O�3�) W���#�)~$�=��"Obaz �>4jX1!N�P��h&"O,H�R��
?��n%���)�"O��q�iȾ1+���N�
�6=�v"OFu��MG�	8Z$�4���Z�(���"O�� ���#E�DQ�$
�~�h�)�"O�����;����SNT*�X@I�"O�����ռb���!P�F7Gs\4��"O=RUG�M�P�B��� ���["O��@w�n�Љ�Ūόߪa�5"O�W�T�T��	r�^�G$��:d"OB�NA3 V�����̔t�ze"O�h������.�Re�N�!��\�"ODq{)X"Y4��K@d�Y��L�"O�E"4�]Ͼ��A�ڄ�@"OT�$��D�*.m�|���"O@e�6㐦H�����ŧ,�zX�5"O�l��*B #�\"��O�&�f�٠"O�P���,������̭:�p�۱"O-�nѡb: y�@
n�fh��"O�H���	:ڴ�:f�6�>�r"O�Q�����(7���@�<3>���@"O���0]Q���GR��a�"O��kd�O8�^M�:H��	P"Od9j�� *�iF��&&6�9�#"O��2��6���@7kE�&6�x�"O�<�T#�;�t-S7C :1#����"O��q5ّ�Ւ`8H��"Op��a)I6_��cI�[İ�c"Oa��`�T�ӭ+���S"O�1 �˓�V)P��0b�tm��"O���a�ۏ/�YA���(��$!"O�i,��J��0t��1��Y"O�=Q�@�p�T��S+?]��A$"O=�f�P�NtY+������X�"O4U(�ЛM8���@ �e�-{"O���6dM�~�Z5+D}�� b"O��&�(]�dT�rT�@����"OL�a0��
a �"b�&`�H,�$"O"Q cc(B��\�`�ݼT���Y%"O�,���ڒ_�XJfN�3(�ڱ�"O���S��d�
1��m
�y�w"OX�X�O�q;.=�[<A��!"O� ��n���@a�Ս)+����"O:��&�ǅ?d)RA�D?C
4�b"O�Ј�Bz�F)®"��i!"O8I�֏	-EL<Ц%��w�L�2d"O,���U �x	���5lt����"O�}	��\��i{�
"l`
)[a"O*0r�$��$$���Okf-�V"O��k%aJ�ڨP�+�4��"On5{�I
�qR �:d�3qL(�U"OM!�K̬d���f�@ ��|��"Ob�R3��,&�e��k^<Xnx��"O� ~I�դ�	+Į���
�*��"O�̊0łj�2,��*�T&3�"Oa��Ѳr%N����E!%@�"O��À%?U������ C�z��"O����ˌ@�f��d�@��p"O`e*%֠���Rub\�h�bu1�"O̥���ΣD(��2 G89���v"Ob� �P�/M$�3�D��wsR��"O w���]��Lh#�wV��з"O�5��HҼlC4�yfcZ�+A c0"OzѢ"�H'B�,��+M#?/<��S"O������q!^<�3뇣p+tY��"O�|{2���L�b�X&*�<��E"O�5k5��0��Ԉ�Z�2Ћ"O�T��D��u(G�#SFL['"O�h!N��\]�u�X�Z:b�j"O��3��sGT1�f /@�j�I�"Ob�C�F'��JpF��9%p�q"O�Y�,\�\8�EW 0{����"O:ś�hɽ-�ބ�QD�-)d:�{"O´������0����mT�p��"O.]�įΤ"�F1V�U &P��S�"O��:H�0s��;���y"R�S*O�9b���W$FL�����}2	�'At) %P;?�,P#UEǷj��	�'\tdQ'��/� ի��D޸��	�'�L � ōu�TܐQ�u��s	�'�T�I�f��cm��0��928`	�'���"+��D8]��
V��<�	�'�E���H?*R1֏�C��q	�'� ���K�<�Kv�&�
�[�'�Ƞh�a�|�P����H�����'�fIf��.RI<`�$�m5h�X�'��H�3��1�ujf!B7d�3�'Q�E�J��+�(t��ʓ�-��(��'z��e��-k��c�O�:8&|M�'�x�[2��la�U�B�J�,⨤b�'$�qSs���p	������nSܸ�
�'}*|q�*�8~������?O>~d�
�'��Yk�.��bn2��&�>8,��'��UIr�M�|)���3F
67�B��'H�ܺ1.�u�%R��x�� �'�̐�c�w����]&~G����'_���F�d���QB�� ��'(|}�q�I�K�z��`��nY�'Y�ĸjBg.��"�	z8�̰�'�[#�ׅ{)N�s��BB�as�'Q���X0f���(B���6��t�'�@��m�%@H� )��@�'�����O�4_�$�-tcN��'�l�	`IY[��ENŲr�����'hV��Bʃ@�L]8�$�VINDC�'1,� �C�"���k.H�h�c
�'�V�`Pd�����rh�1*��'3(HX��}�*9�AC��v2�3�'^,����<�:	����b\�9)�'�F�:e�)P����[8Hm ��'��`(C���Ї��+	�'��p����u	��AJ�!%ִy�'�*�1B"ʶFp�	�bY��"a[�'e��cul��T�ڡp��7ym��a�'���v�@5#d�Q�	�D�ȉ 
�'gz����]�G0�1�S*C��@�	�'� ��		r�2Tӱ�9O#�@���� �;�oB���Sc��-�&	�"O�BT��L�����!챒�'����Dh��1�R�`l� 
���'K���0�G
`�>�:t���m���'P����6��!�&N1jt�̓�'���;
��x�D,:�n���'�-!VBQ�[ծ�*dƐ]�(�i�'1@a�7/ׄx^Ɂӡ^,R��2�'���nK�8���#��UU0k�'c��)�Y-���j"˞�O�@���'�"���	�!�����'3�U��'N^��^�L��0	�#jt�9�b�P�<�kO7U�@��A��x�. I�<Q�͒5/�qi����<x�p���]j�<���i�d�)A���kR��y�g�b�<��IQ/(���0!Uv���D�E�<ц����:�v���꺩��s"O�����
R�4����1�|�3"O�3Ѕ��#m3WIrL�0�s"O�p�Bh�8��s���yA��a�"O8Y���Q�AU�_�Y9d	�Q"O�� �I|��Xc��'t$����"O.@��m�"5@���%���Y�+-D�<8L�y�^�8$�I!._\�e,7D�dY�@ũK�����ȳl���`&:D��Ѧ��R_P�1���F �u�8D�l(
�L���c�BH���1�!�d�*����	�<@4y�Q�Ƒ8�!�$�(��a����*
+��2��:�!�D�|�~x�D� *�q6&A�)�!��F �h���g��@�T�S�Y�5�!����w T.n u�u��i�!�Đ�[�fm{����L�bK�I�!���$:�h���B$6��UR��]SU!�$ҎHތ4��hN�H�"P
4��D!�()�p(w��3 �A	��!�D�e�`i#0gF���\( ��*!�O���qj�8H�����ۤs�!򄘦3�	�����#\��sKL#l�!��01; ��gaP8=$�t�9+f!�$��s��8�2�۹E�q ���$y�!�DN1F�q�!-��8���\<�!�\��(a��O�!r؞�H�/��<�!�D�I<6j�F9\vĝ�N7�!�$�[��u�&ꓪ&X���)�!�D�&�Zy[�gO�:�N�#����Q�!򤜭"j�GJ�bCl�0��5�!�^,XF������!�Ft��%ΘI�!� ����Vd�$0�=���'2!�ʷv/����+@%!厞4&!�D�&t��J��ܬ�qABd�R�!�D�D5<����*XbEq$n�K�!�dZ��e(�Ȣ1*��2L�*�!�̙e�@���"j����e[q�!�䞠R��P#��u��Ax`���iv!�$�v�F�����HO�#"}j!���_�m8uF%5L��!Cd�[i!�D�,��q���.D=!��	T!�$ӧmQ�9�.^7*l0�vCKJ�!�$͞`�d�'F�<h�	� ڭ|e!�Dπ?����bg[�i����)`O!�� rl�C$��&- !c%Ԅ^o!��+�.QA0�Ӎ9/�!�8J�!��,G�����I�>��H��M��!�� v� A�����%�0t�h�qw"O�ĉ�&�%h���^�!��J�"O�أ�#	d����k�_윻�"O�!���&Y@����$k^z�!A"OhY(r�Ο5�T�ر��gkZh2"O�ez���l�p���+�YQ��3"Oh���@��˷럙wC��#"O� �2"�Mxh�u$�;~$����"O����d\�R�t���!TD�z�"O1�oز=�`%�ga� �D�J"O����(OURa��	�,�z�kt"O*�J�F�8�M��D?.�:q� "Oș�֯T�q���R%e��f��иu"O�q�a��5%*�z���K�h]8�"O�0�B�T��i�@#
�d�� k�"O:%���;�ʕ�w�ˤj�pD�"O�!᷃�")<���C2�⽁�"O��Ϙ>[��a��\7�Z��U"Ol��Dn\�]��[�ϲI�NT�%"OlYQu�ޥF��c���2n���""OX�$J�( �+=td&�"O��=V}K�I�v\��E"Od��� B2�ԥ;!�,x�n<Г"O"}i�'U����K�-���ab�"OP8p$FD���;5��k�|I0"O���2~]��R�<��y�"O �f�+��!��$��l��X��"O2���а<Q#���;p͖`�"OP�9��%�rxGÀc��"O>X��lI8�8��ܑ]�A�"O�q��O�b�h^=C�܀0"O�Y�j��/[*�aQ 
Tθ|	�"O�# ?��Z������"O�����<�pCN�>��#�"OfiAO�Xu>���ʷb0���"O:1���>M/T԰SH�Vvt��"O�!z#!T9�,d���MG�*7"O��! �<sznl�  G�VQrB"OԴ��ˈO�.���������j�"O�q�F�*t�4���JX/$"��z�"OT)�j�_�i�
�h�v "O2�j��8o5�d��G����"O�X��ўW��0�E�[�V�X��"O�x��O�!g��ݻ�N�|�$��`"OZ�j�lE 1@Y9�D�) �D��"Oā�sFD)���*��T� $�%"On}� Gl�i����&�|��w"O�����l8��CUhҚ�0� �"O�� �ہR��3�����j�H�"O�x���P�y�I�Wn;R��2#"OV`�t�ϣ5v�`��#Q�-U����"OЩ�jW>.O� ��BN/�袵"OrLЧ&�8l@�yY�က
��k�"O8�Bg�g����W��77�̺c"O%��H�U����5A�&:�2��"O�A�*A�n�H@�ºL+����"O��f���=v1k���%�$H�"OθТC��)���S�'Zm`�"Oy��!���#��}��jc"O����	N0<� �g@�5��U�"OȄ�t�rĲ���	G������"OZ�sЁ&<�R�*�ǔ:MG��bS"O:� ���8�J�ᐤU&6�a#"O�a�����=�$�#�;(C��"O� .�B�CJ6����P$���"OI�����8���5x^��v"O��D���WpI��̵\�,�"OP����"2M�JðDdl@�*OV�`̊K� ]���=F��h�'� �SQ"�-/�~�R�m�	 �JEI�'�-�S�x�FT�#-	=q�� 8�'�x���e�/f)��0��Qk�|8�	�']�$iL�D�t)ϴ8,޼	�'�0m�#m�, ��`�l� (h�P��'�n�x��Ƌ�*Ex��ǯ%�rx��'��9���];wj��T++�l��'�:(�1�ё{����$㕢3�l�8�'V~� �R:��q�C$L,S��X�'�>�x���3���!A�e�љ
�'j8�@�c�.�n��UN�^w<��
�'��Xk�g��6�� �'�n�j�	�'©	�OK�26t����Q�`^�:	�'���*v����鋅��Y�8��'�`��E�c���*��� ����'��M��_ZJ�����&���q�'l�4�Ц�?J$�<�c
��%j
�'8 �T-�1`�X ��aى-5��	�'d�Br�Q{�\<:��:*Рm��'uX�`�&�ġb#Œ#�����'���m֮�8=��Z#Ey>P0�'-n�GA�/K�4��fJ�BehEi�'���)^%��B��#q�b�'�@P*���g��Z��]�IAx)��'�&Qj�Ԅ�<�X��\<����'�젉�.ȃx�
4����-�� 	�'dEa��D�~~�+��p`ɱ�'�&%�d�Z1bŮ�֧ݥ=�@��
�'�-��)C�=]������y�,�
�'G�)3�Eh�4q�+���
�'�``Uj�[�wo�Փ�'�H)X���Tv��d��>_V�Q��'����/^`�#�Yg ��'�
�*a�LcRF ���7hr���' ��Bqj�Ep�k�W�g;줠�'H|MP���;�ļ�v�ۍS����'����3���V@��.��
�'�!3�*G&v@~0��i���4�	�'줕P�e��P���n{�`z�'[ZQ��*]����lϻj���'��<{�Fƺw��óM�"\�ޡ��'�.\:�I���d��Aۧa$��':*����92��8!h��[�r9(�'�:�x!��2c(��×�H�P4���'��yڤϙX�ԩ�"h8HJT9�'C�J��ņ����� ��K�'�,E�ׄ^�))���N�'` �;�',�����@
.��g�>�����'

�RQ�����x!0!	d���'Z����i��`Pq�Q�|?��'�,��0₩q�a� Ŵx�B��	�'slR"�̗4Q�X�kX�~!��'��J򃁵"� �i)��q�����'�4�*� 	�lZ4i��'~�ȴ�	�'���s�d�H��t�S�-c�<��'�Di�$�Y�0�C�%�2P�H	�'�x���(�(,�4 �ׄ��	��9�'��D�V+%%{�@����V����'���-�9+���)�^�R��� Z����O��5!�iƕ
P���%"O�q9c�@%T�iC`	�r `���"OV�rsɋ ���@t(�� ���"O%Ze��/�I��)�pU v"O&,��oW��>=�W易B�����"O2� �b��2��e˔jΧ
����"OTAxM�Eׄ�q	Tb�Ƒc"O>yc�˝�w���y�N�"��=�"O��&�pl#� L���t"O��s�K2#��p���x|xJ�"O���$f��L��Pq�\"�"O��`���a����X`�P����yR.��E`D����@���yb,��K�z�S3�?P�Q����yF�=\=�qc���_��HCfF��yb @u�0���F�#ЌE�4+V'�y҇�x�����#G��@��Z/�y�-ԤK�����͆L��4��$�#�ybǉ�%�A�m��D�J����yr�B�rȡ	{kJ�sw�=�y`�)c��XY�l
�$('���y2���!Y
\���?�p�8v�Ŝ�y��C�>�����#Th<h�/ւ�Py�	��0�<�YV�h��d�b�<!�>:=z����1���_�<0lӔE� �fHѻXq��%�ES�<Qb�T�ziH��$o_���C��G�<���B.3��	(��K�5A����oi�<��&yz"l{�)�\{T���CN�<a祕�j���KD�߁9���AKH�<I��؏f�t��!�H6	��PJ'��@�<AQf�w'��Ǒ/r]�qʥ&AC�<)��R)
��E�6�I!v��57��h�<���++:1�0�Й!� ���g�<A�NQ<4U`�a]�[C�L�s�_c�<�׃̜[έJ�Z#	O��`d�H�<aM	�j���8d&�/vrx0�A�<���U�aR����IQn�����<�aI�Jh��1��PF��6��F�<�e�PvT	�-*>$�S#�F�<Y5.ũ������	k�)�q�GD�<�U��T.P"�)K���A�C�<%��o�4�`K�$fw�9�5hi�<���Ӱٔ ĎN�K�z��{�<A���-�pA������Bg��P�<1q@p	�Y���d�x�
a�J�<Y�.
/7pҘ�`b�=��S K�<I��ʛi�(0���8P�f0�ΌN�<��aU)|!0cE�::�n�u`�n�<󈏥|�9��!�3�ҨI�C�n�<!vmY/SĚ�
L�t����@�l�<!��2B��{#���\�&@�m�B�<AB�7]��в�]�~�K��RI�<���D������e3n�1AF[�<��;���2D�z��5J]�<IV�
a�"̓b^����CSQ�<�ŭ��X+�iD�M�RW+ f�<��C�X`�gnוo��$��*�g�<a�&G�j�ֈsc@���iѩ�z�<�G �8�.x1�W�#��	��Iw�<����H��z�Y�w�l-�0'Lt�<�7憐M���)g��y��0�R�q�<��gJ�j����n�2)��k@f�<!ᦊ3�EI�"f��@W� `�<� ���я�B���A�5(҈)7"O�	3����V��y��cF<hz;"OT�Suf�Qj��ʧQ��|H"O�����
�gn���Ԩ �f�*Q"O$��un[4B�+ .��W+P���"O0�K$�u��ZL������"Oڱ�`�!^������}�P "O(����,NET�� �Ip"9�E"O���.(BC�DБ��4i@4YrE"Ois$f��c_L�*3
ԧp�� K�"O�1ƉRy�ls��|��ٛ4"Ox	K���<`q�CɁ�zh5�"O�y��o7[���+�T�"��Ւ�"O؁����Fp
���A�Y�n(��"OTUKBcT�Y-����F���|[W"Ov�ѣ�ˡ��|�f�E�Ѽ�+"O��q5k=!	����C�����Qp"O� �"�>{���1"�4 �Vp2"O�y�ի�	'
D����0�j�� "O��)V��([@�n���qd"OD�[#�\`�)��'���u"O��O���F�ʶ*+,���21"O6���ᓖ	/��;�)͈ ��H��"O�i��H�2 ����ҥ�/���4"O�)�rM�L����~l�g"Ovq���Y�5F��kũ��!��"O؍('��;Y�2�А�\�K��� "O�!�3f\1 �h�	�0l�V`2�'m`��o,(����[6��|��'	Ĥ�U"шC(P�*�)Q�4Hذb�'"P1� FP-ީ@#��3"�D��'� <�bNW�gɪ �B�'r�}8	�'�y+��Q�BFN��W�Q~g:��'9r�ң
љ2�\i*�n\?`��\��'��)�B!��j�@M
 �S	o��|s�'�`$B�-%z���i�7�  )�'��@�ª�+P�IZǊ�[����'�j=��#*P��!�5��N�����')�tI�Έ�`�t5)$��#Ak�)J
�'���t �!"��{�؉@�vd(
�'DX��2+Ƣ ��]�����1���1�'��K`j%.�P*Gb�6#�~�'��\���7R�Y�GB^��5 �'��UgG�T9p�㈸1���@�'�ni��ԥs��:�/�]ʮ��'��!�$]�#
`��@+P$*X
�'V֝!�M�h�;��^�H��u	�'�8(�3�έbd�C�B�	`���'%�8���þ
<:�h@O��,Jh-�	�'�
�`���?H�P+��И(��H�'��dW�
�
���L-W-`
�'l:|h��;$|�rL�^���	�'��ȉ�Ʈ5�IAA��Ky0\�	�'}:I�����A6��h�g�E]0	�'���3��O$7l�倷j܀��0��'� �sI	��\8`GJ��JQ�|3�'VD@�F%�dЈ�&#�-D���'S�����V���(�E]C�4���'�ʱ�� .G�R`���M-��5��'��8�A�-�j	CDH������'1B�����9�J<+�-Q�'M��k��(y�@j^́�	�'�T�Q�'��"��!x�R]"
�'D]��g|�4[&�8r���
��� �9	���y�b��A��

�\�"O�mJ��D&-t�\�BE/vLtX
�"O�9 E(R4��4k��ǀ_�di��"O��`d��.9���h/=�b8�A"O�9y։O)f3�QHqiL�Y��ȱ'"O�SG��	5�X����#Bl�
"O����d����&G%9U�=�"OL�Ȁ�߆:�>8��$�
jF:��w"O��Š8d���j�M�|7>4�V"OF]�Ņ߂! �5C���僴"O>�����):�f䘀뚓^�t�""OȑY�m$SqX-h0+! �
���"O��'��,S��)��lK6���"O�� ˇ�s�xi͒>U I�5"O�ث�i�봹�P���M?��9�"O�Yы�5	v�
���<8��"O��2b��y8V�kR�Y�H<�r"OH8���>�,TƇU�w|h(�"OF��nƲm�xI�@��{���S"Ov�e*4�ހ� ^ �X�"O,�г�K/
� ��Q�8�*�"O��s�'�>Ɣq"�[�X�.A%"Ob����P�N~$j���h�,�0rl!�D�R/<����-X��y����*i!��
�BTIƈ{�>(S�`#IR!�$ϼO�vhp���Gy�����!���HYi�hZ�y�t(�(��P3!��e,R����э#t��@��1.!��S��JŃ��^e�������!��/	���f�Ɋ2()��:�!�]�HX�%���% %�=K1����!�ĭ3�fE!�b��0xY�s�C3\�!�JeP$0��r�z��C�Ƣ:�!�*Z����&H�PS��߇<}!��2�A@�37��`��[6hm!�dک`6���'84V$���'c!�d��7�L�K1���A�9Hw�ڨ�!���Q��H�$�1�L������h�!�d�]p�ɱ�eƬJ��TI2�̔�!�GAN@|Yc*��R�:�I�_�!�d��*{�Ո�ׁX����hE!�$ �;s�A��׊)ܰ����@:!�&g��k��!K��ܻ�@	�j!�͋|���%�iL�p�1!�D�STָ��	X�xX��UV���Ĕ�;��X���;~�����@.�y�,� ~͋�U)z\@ݐ1���y�)�x�v@�A�K���p�)��y��A�:L@���֢ >%J�\6�yc�$5��1��nL�|�Q�8�yRg�/����B$��{�k���Pyr/��@����sHʑIZy�'^N�<!�L��|���x�!Y�J�,�*ei�P�<�%�*$f���I�`��O�<1!)Ӥ}U��p���x�IujVG�<��K�u�h����\#&�Z�<Q�I:GJh�QQd��fH[��P{�<��c �Q� �2W�H�p����G~�<	�G�-GW
͸�V�X�R�� t�<�1c�/���qgFߚp��M�4 Dg�<��N7Y�	���8��ad��e�<�3hP�;\h���֓�ёbN`�<qN_�0��q�H¥z�LX85�[�<�.�/W&8AP�Kɇ 
Xv��K�<� ��c�Ҝ1�:�"cE2~��l �"O��9`H�0\zp}��L��I2�"O4����C!�8�K�5u�%��"OX�ED
�h�̣c��y��Z�"O�C��:'���÷��/�\I�"ON|�"�2i1Ұ��@�9�P��"O�Q�e�1�ƕ�� �Al�� "O���e�z��10RF�<-#Zu�&"O��xq�R2�*�3�%V�8�ZE��"O��d�1*����;z�f�A"OXY��l͏ �2�N�d���2"O��	F"L�>����ʳg�MC�"O�p�Rb� @�6L7v�*��Q"O��r@C��)^jUI�o��2���"O�uC�U _��˧��~�h%�"O^\�����\�3/ʰF����"O���p�i�tG�,@\I"O�u���eY�pĥ�/ 20��"OnH:f�G/u��˳�ۡT��06"O�dY���-k����L��:.��e"O�,A$Mש@G}��`�]����"OXW�8�P��%��[vPʅm�}�<�n�C/T-���_4C7.�"��c�<QΐsJM���4j���^�<)ӂ�C��\��/E�N	ɢ�H]�<a�@�m����@�?��P���X�<���͐0��c��Z8Hs@)���~�<q�gZ�;E b��Z61�A�P��z�<�6N�P�<���%�3���h���s�<A׀[?\E̜�DEI��QdGn�<��K@8J0��:g���2�!��U�<����+]��Ȃ� ���'�O�<��旳\��y(�MO ��ĉD�<)����F���s"�>U)���DB�<����.�d5C��^:rrK~�<��O�n-l���J)\$��I�J	z�<9v)O$���gO�A��ѡ�^a�<Q��<"���jʎQT�eQ��D�<1Ѥ�=Y�{bˀ�6�~-��*�@�<���R0�4���ő�P��u�z�<Y��L�?��(��g�.G�Ƹ�y"���HF�@6Q{��Z��y-٬8Dm����H�7$L-�yR���	�>� Wi)L1B�����y�).0��r���.Ԋ 	����y��I�
�!���U�B�X#C��-�y���V�:�F��	 *��SMV��y�'��	�����٠Bj�$�yreF�{�N�)煛~,��AL�<�ybm�~5*������l~�ѻ��H�y"o\n��d��N.^�z���5�y�*�~� 0%ہR��Y�푹�y�
T�*Z��Po�G��%���є�y���|G�ia�`�D6���@χ�y�*�1�p� ��QT� @eiM<�yB�8N���d��+G%�%�&���yD�
2�D%�Q�ڡռy�ca���y�i��*68p�E׻S��X[�kݚ�y�LՀ���-
"|�4·w.��Q	�'k6<�����kjܑK䩛oY�Y��'тq��$�3	�m��k�`.:�H�'��0beD�Y@�]��X�$�'�l�B�Ć�q��}�f�C=�DI��'�td!#���V�f��eB�5 �]�'�h�Dy��� T�SP�����9��Ù?$0�b"O����
��;��Y�Im�((��'�Q����#[���fB��a;��z�D&�O�wxȝ����	�v�y��M�4rP�DyR�'��u	$��82���0mӚ.�z��	�'%��S��"2����+�L��'	Py�h�&*��`�g˞9�� 	�'Nb��Ag�%?<��� �h�̼�	�'T��/E%l9�A�d?J��q6GU=�yhd8����J,�)��Y�0<��$�M���/�*�!q�h#a�n�=E��'R�A@�oq�x*P���:�Vk�'�:����z��"���B�p�y��i�!�dKa��ȥ$Лf�0��e�_�A�!�J3D���~	H��4'��@!���U�x�W`��BhFxX�%�"�!�DO�}�)�c�L6K�Hr%đy�!��#xx4�\)T`pgՍc�!�Ą2��҄�u���s�M�$�!�divd��qo���(�%��m!�d�� 0�Q�ؕ?�� �f�V�2�!�I6��LѺ&��䒳�οPu!�DW1#al!�-�+�LA+���na�D%|O�S��P��*̾[�K\ JhɡI>�O�$��3�����ۭljz,Q�!�HOa�T�23�^4(�E�=h��PAjA��O%Ezʟ��ʐ��a��Q{�3"�]��'��D*�)�T�L���+�2 Ux�RE"6�:	���!N�Z��� ix@a��\."�!򄈶Uڐ)Q��b�||cӎPo�������)��:�նf{ $	#.�O!�^�<���͆1c��R�$E��$�S�O��eg�(X��C3J_���5
�'��l�7AP�/�¡�C�Z,�l\@	�'7�e�S�M++>��b��*�m��'����f�!F�d�rB܌r����'�Bq�㭉�IW�!J%V�h��	�/O ���H��BA�M���pMT-(�!�d�7��7��g�T����$���=ɍ��T�f��y���Qe:5��F�/1O>�'. "~�C,�/�����:w|Z�3��D��m�d�[�����@�@�xb�e�a��5X�B>D�Lq�LbUЩ�e��' bX���N'4��9(�. a�1��-G(�L��7Z͟�F{J?Y��>)e*�5sK��SF��wo�i"7cFA�<QZ�xV�)��QTRT	�~y��'%1���[� �B��=0�(���{�)��@�l�<ݢ�埖cY�LKK�:!��E�- ��ã[�=M�8p�,D�b!�]mF�]y�Fx:����] k�!�D��6UKf�G��
(p���!��.AKL$X�)�0^���Xu
�
y�!�$-�uZ-ݫ"Uc��;.j!�ĝ	I�^�!���$|�1�)M,`�!���o|eʑ�2���b�D�!��#n���$R�KU�����)M�!�$^�}Б���m�F���F#�!�d	5$�`�;��ĴL0�UG�l+!�����j��\&1�ҍ�p%ȗ !�I@-�a�ş�0��؊CI�>Y!�$ȫA��*B�0a��s�O9H'���߶څ�<O���[ĕ�7��(�y2�'�f��R'L�� �4.8���	�� ��MC��̪U�\4���5��2���t�<� 0�8TN8�B]@�	۴< �Y!ቸH�	�*�>�*�y�������(��Żrb�q��$�x(�="�:-���O ���T�C���N�)��hR���CfR�1�$7j]J�M?�	�k�Q��d�2�E�|N �k@g�,��`�x��i����>i�{Rǟ v��`p�bR9���5�N�nu��=�;t�f"<1��5_�]�0� U Qa�K���_�&=��rS	��r���b	X�n�"B�ۉ�ϸ'b����a4�]��>��1 	�'��$pGA�5���"g&ߛ
�R%h�'�D�P�I��h�Њ΋3�*���'C$A�0��Dpd���F,/#� �'�
���#��4�48���+Wh�	�'"�iá��b�:�t��82�R	�'�0I����pY�@f�<4脌x�'���"Cb��Q�z�*���}: ;�'p68���
�S@�ܺ�o]�y����
�'S��A`�ݢ:����`�`�Z	�'����[�t���H�T���	�';�������1@�+ �P�J�	�'�������<6����Ai�
�'��i�F���^"�}
���h{��K�<�T�(4����5|h���FULX�ЧO:$�'$ޥ��ĀMw���D��P8�'J�т��9$"t�A��FUێy"W��bb�'O}��`��k��b����9��C�	$h�q0��� hy��8�^�t�#<��5O�S����'�r�[�a@G��퀱"OdeY�C�	
�"< ��|��Qz"O�-��h�NU$��ąɃvXY�4
O��QE�ŤS �!)���x=
��DȢPDA�B �?0J�]Jv��Vazb���PCR\�o�
*H� D��>]���~��H����Cǌ@N�Y�c���U"O֔�g�I�'���Z�E�'l&�h�e����I�J��g��� ��k�"��ШB�	M	�	k� �	>���ȃd^�36C䉀�Q���
eԎ�rC ǝY,\C�I�p�������]�x���]�TC�	5p�� ȴ�_�R+�X�    "O8A���Q:B��ŲA��B횭�"Oҍ�q�ߧt���p��ʁ��@"O�Y#�T�n ��0�[0_��1��*O�j��+;�.��ӊ,Պ��	�'_��2�V0����wb&;\8�
�'1Xh�SA�j�X��"�<�M�	�'Φ��$��*J�ȃGl�(t�<�
�'��N��"t�К�n��&yd�I<������BG8aj���! ?� �C��]~�z��$�� �` =Ң�;��ݐ��+��U�'��ɾKT�q*�&׬&tZja(Z�Zh�B�	�MS�+��@z�r�
$)Mh�+6���<!�}��MV�Op
�#��J.>�V�;th�11����r��'�HhQlT|�����1K����OL���b�<����,n/$p���=��~"W�,Yf��i�T-)��B$��0ɤl.D�а6��5k�R���^�9�����*D�X��J��V�:I2��%;��R�k(D��ѢF��:tKq�ґ/Rvt1	(D�,�VhQ�v��
�Y|*��m+D�H���[2��5��8�L�Se.D��á(S�Kj��k��$M8���(D�,��9�����2@�d��:�\B�I���W/=(�j�ά�B�)� ���#��aOV)ƨ�g"O����О��IãN?G�����"O��� 
��|��O-�+
Lt�<�&�E�<�zTa%�0$�}����m�<I���&VX)`W� ������j�<q��WM(�!�g��&���4fM^�<Qu)@ 5Iyh0�Zz�n��v��Z�<����$ބ[3jňf#�	1�RZ�<Q��K�R��Yҍ�l����A�V�<�ԅ��=DU�"J�-�x�T�<�p�%f([tN�(BF0�p�He�<QO�t�z�A�#S�JݢW(�Y�<����9MWʽ��\%~��$�6AR{�<1���&���&h�|	�(�p�<1���X@]��[�8_�!G�l�<�+ĴS4��2 ���5� ވ�y�7:�����b���y1	�y���RJΕ:hL�U(V���@X
�yRe���U��B�
K��Y��yR,�	{�̅Pb�B6I,�E�-Y/�yR��9(N���%��s���0
��yBfأl�թ��\�sA��X����y�|eX���n�U@ė��y�6@�d;Sȅ�e
�x�%�>�yrLF-�Ɂ䬅$o�Ѕb�-�(�yB�о�:��#�|�H��G	��yR���b�|g��&n�P���hD,�y�̫D�>8�u��:Pz>�j6���yr�_6���ҭGUdIcK_��y2b�9C�NU�Q���k�ZIH ����y� ɗvs�i��I�a�Z�w�-�y"��4?�@1�1�$VT\��O��y�Gئ=��IHJ:A��0���A��yBO��}�%�^�;.�a�lO6�y2���'�Tk!.�8`�=2�AT#�y!\�1	���,:0�4J��Y��y���;o���G*ߟ'�� �(V��yb��W�4]�MJ ݔ��mB�y2CWh��n[��Z�X����y�B��sg~]���H����
DǍ�y�A�D��$�7C��+��h���y�'�:6��m�� �n��yB"EK*&��ᥕ�	�P������yR@T� �@H���#{'H���y�ϝ�(�&q��ğ.+��r%n���y2l	$�Up�̸A��(��Y%�ybѪ*@pr�N� $���!�yb��2Jc���0@R�R@F�B����y�T-q�Ns�N�MmƑ ��4�y�)U�o0������L�fՁ�ʲ�yBA�P�A��K���Q�=�yB���\�'"�U�̔���F
�yR�SfP����2P�Ќ����y�a�0{�@4Y�e&1��U87���yRB]%y��i��H�(qP��ɦ�y�D��%�E��3��hV�-�yb�D(���3�\�.��ņ
�y��K���8�kB
D�1+A�y"�
����L>7�ex�U�ZӔC�	�5�����'�pՑ��� �:B�	?=r
m��ǲ
�0u�u��4B��_���3k�]��/)ZB�	�ar�C�)����o�*YB�	HLqd�4P��A�uÕ<g�F��D4�S�? ,�)�;YeH���7CK��"O�)aw�ي=f��ui� �Ոv"O�P� �;0L4�����M�m�"O�H1�@*(������L[R�ˆ�Oܣ=��a�5L��q�#=�ƈ��j܊a�E��I�0��D�#�t4���Z�yg>�k���D!�I*D�v�ӔA��'kV�Qk�= V��D�$P	U
��@�xQ��4��2�M(O4ʓF��>���Ʌ̖��B�"hM�u��a��/K��#6�Vi��Q�$MTP��ȓj�8����0tFE�� ��m$��<
�qF�pIe������MU?tT�<��	�!u���*�4p�#�(�V����^�G4���F{����zU�Ʌ�8��`�� q"6���'.B0Gx2@�(<U�*��݋e��lBP#��y�lӻ9�t�2�KáXi��As���~�D��h� �A�搹D�H��<�D� ��'!���'?X	�g�8E�!@F8H�:@��{Ri��\9��P?3��1��Q"U �1�O��ѝ'z8�)�j�6[�4�+�H�l���L>1�O�c��>u��-�[z����>V�ܥ���1Oh��d�~d ݃�X>m���a͊�(�!���=�x��N�#�t2BZ=Lv!��!#j�!��`�=Y��Y�N]!��p�PT�Aא)M��!��_<?�!��vIHw���&�*��ݴh�Qv�.$�@#��U/<
]*�*�c����@G"�8m�u`��Iu$�(J�}2%��(C�	*~
���t�;:�d���/CjB��D=�8uNiy6��9�x|9��39Fx�b@u���	��N�.Lbq,U @X��1 � vw!�$�@�2\�T �+x,h���N���yb�O���Ϣ��iP�\�V�B���4D{�\����^�S���d��3YƁ��`n�t+vNK%7�de0ւ��~h���J��,�lоpB"�S��<��I~����@�n��J3�&%_\(�ȓEy���l�6K$P& �#,|��ȓ+@���f��>�����%{��H���PQ��M\4 PWϑ#C����'��~���$^|pİ �+������޿���hO��>��A�-��Cm܏��`�/N^�<��L[��|���X�*D�⡀W���0=!@�õzF���6�M3���� P�<!�����z&�ڙu�����.*rOR�y�Nπ:m�pu�� R�"O���aN0Yj��K�9ᨤ2&"O.�`��X�r^��1a`.t�x�* "O��K�oк�E`��
D�x���'l��i����3k ^��Pv��@h>�Onʓ�hO�	(t  �e�h,�����*U�a~�Q�x
�*E̤9;�G�8*V 㐆3D�����4E�6l��E�]DXC� 2|O�c�0�V3.�<б�囏9ZXۅ�<D��h�NK��p2��<G�b�L9D�[�lU�
#H��'	(ȉր;D�hx�jͥ)��W�ܱG�����<���<��M�=E�ʜ�ň2o��S%�r�<�'� �j�4S5 �|��Rj�y��hO1��|Ɓ��F+f0r�$'����"O�9b�$�+���qL+Lݾ-�1"O��r�M�2�����5��XB�Ir����+�E�h�X'�~ �y�H5D���� �'Ԗ�+UJXcV��+���O�B�)� �Ұ*��"�"��t��/G۲�Q"O�y��!��6�+afQ'q6aI�"OR$P$S�+_Ԝ#���l#�@��"O��Qv�Q�_p~���8*sx���"O�:���5@�
�y�*�sxq�"O���Y%v# \�pk�'I�O��� ��*{9N�aF"�@|ab�"O��,ۙ1�$q�ɁH��
 �N��M[�}J~z��
EJyG'Ũr�p�r+Xa�<�d���8cB�M%n.��0�b�<	�JH�}h�!�,xa$Ow�')�y2L�.i�`�C�6�~�1��W9{�ў"~����K�nJ�W��va(D���ȓ~ߘ�ZDH��,?d�TNN�S����-\�AΟ<*���0 �� ��	�]�I�R~t"S�ɖ5ixTs�M	=sMFB�	'v�.�HW�>H�L���#u�^�>Ɍ�	ٛD7b�+���{�1Yq� $��2�O����+�]#c�<�9�"O|��ŢK��,��a��G�(ĺ�"O�0s�"�\ȚM�`�0�����Jx�r�W�f@�5&]� U:��)-D���P�PO�U��nPnFL�Q��*D����m�o~�g�\@���G)�Ig����%J�.jV��t�t8m��;$��#R)$ �m3wN�.!���ۣk�/nj�d3�S�O����D�Y�"� �Z�Dj�=���HO̸@�cI�}	j�#K�`Bs�"O�׃J�yf���d��jŊ��>y���)���Y�qNij��ˍv��)�S�OXF�w��=o$�{����S�N$��'�����
q8օ�p=V����O�����-l�\-!k�$��hD$R�&6M:�O��3��Ԁ��K={�@Ɔ�p�,����c��B�$�c�L|����hH�.�4�?Q�'�#=�)q=ڦ̎$v�����)�C�I*p�(�Qjɪ~Ê�XQ"ԄH���	��4�~&�|qC�$�̰���ĻzB�0q�7�O��_b��Nǿm�Z���`�t;Jm�W"O�0�B.��-�|����@�C�"O|�q �ۤ >�-{ U�(�)"Ol�8�
�^�9�ԣކ �ԉ�C"O�3���L(�0�1�Ԏ^�\��O�Y��lΦLV��+�(�E�:�"D���  ��$�"Ϣ�q6��>|��P��I�v����W�*̙Ћ�*�*@CUN/D�H�'�O�y"tF�|��1um"}��>�Ó$��k�AP,�҄��
45l �ȓD�0p"¥^�V)D]�&�T4�YY�'J��p.A�@��z�JIY^}*	�'�<�ŬЀ}���Qhָz�9	�'���D��2p�t:%��G"�`	�'�5�7
�!#��ҡOV�F7.]�	�'�$|�a���<���PA֧=y�l��hǽ�(O�>�A��t��SG���|@��+̙�ȓ/a�8p���b%�v���������	zy%.�' �0�!�� N�	h&�g�v���X�?:E i�&�	���Wꡕ'�0��O,��d+U]��,�$w�&��'�a��}b��t#���V&.�%v��BqN?D��ҡ�����p�dW�%>:5�,>D����g^�>�Y4�V�5��e�A�7D��Ƣ	*n��@U�16�a*�E5D�¢/ߴ�T����T	Rd��&D�� �ۣ����h!�t�%�V"O��5+�^2�B���<m�h(�"O�� �Kf[d`�Vo2\L�u"O��K#?\3�E��# ��q�"O���fB��j�&DȰ�a:x�8"O�[� �7v��xP�Y�;�008"Of0:�ɞ.a�U*t�ԇ@��r"O,p[#�4A8d1��O1�5��"O��kĢQ�(�1+�yf��ۢ"O��:�fF,eV�"K]VwQ0�"O �h$M�<7�E*�ˍeC����"O��{�ڽy8���%�V� 4��"O<� ���/�bx&d^�1<�1"OF�z�b�l�ʍs�(XdX)7"O��XV"�X4�]���%*g��`0"O"4h�n���	sǅ��U�.���"O�,�q(U1G����T�4��8�"O�����' O�����4��s"O�lP@�
cŴ����0�J��"O�-�#ɺ{��UIC�
6q����"OȤB�"_�i�c"�0"���"O�TɅJ�f�`�k��ߚ]�X��"O�ջ�b�Z�Q� �[y��A��"OEa䊎0��TO:��P�c"O4(p��VQ
�C�!B�Pc
�'!��.Ra�X�ٱ(U:e�d���'��a�ΈV~���� /fr��'txQ5��^	Јc��1.�j��',	����^�0�[6$�^�����'φ�p�7���&/�^�@���'(9ڴ��!ڬ ;p��\~64j
�'̘�fC^#d��U��R^�
	�'����;��HZ7 � a2&	�'�TP����6��J��X�Z���c�'Au�ɖ>����G�Tn�P�'gڄpFFS5��g�>I�z�0�B�:��%#1�P�"Ծ(y~�	�
Z�in�܀=D���C<ULt��b��%aĸ�9��:D�Ș���lS2����"L��	��;D�`��hЀx@��g�#s�E"&�/D���C�I<H�����`�8���7D�|��@0V�ҹɑ��Y��d���7D�,�K�	�>9!�n4%r�q�!�(D�0`DG� 93^��0�S:X���	 I'D��ڵ�ҫ1!�*cL�[����� .D�X�q� 'Y�dA��KT8t_��p%�:D���dߡq��Q҆ճ'_�D�S�:�O�T�"�R�6[���V"�*��L�@��O�d��6��m$C�	WF�:���'&�Ȑ���;0��#<q��8)��zEh�1NNt�)I~���[����'I�T%*Јw�v�<!�Ñ"JX^Y���	uh�O]r�<�� P����ۖD_�p���P�<	rkZ�|�>�jV������N�<��o�5!��I.v!��GR�<���3��=h�N��_M�L���O�<��MO�0�z��XWӌ�ҥ@[q�<�G��3b��y3��5u'̵��Ĝh�<	�C�X��0
���t�vI]i�<i���$�4�ˢ�̈́X��=J� �i�<QaƙMmp�x�eUP�9�a�<i�h/`����Ǩ����ЀeHg�<I (�$YZ�9�#V5)�LM�fa_�<��n�*Kr�Q�I¶��!�cȒa�<i��\�r���L��	�0k�[�<� �X�W�ݒ���Í�5b1"O4���ߧW�Py��㎋cӪ["O
]�s�ǣW���AA�p�6]�4"O��.O�/FHq@Ц|��e"Ol�ꐬкP0��k�Oߦ���#"O��٤&A6)>�pcD!F��HS3"O:Թ`�ֳM�H�`���;y�i��"OV]���ߑ2�TP��*Q:%2t�SAW������W��-��ɾkc�ԛA-*s�ǎ�����L�>���oZ�D��$�#E٣GtH��RA�A��p	�'�X] B�HQp�˖&H����$X�@���D��v���?/ ���F��X�j���P�� /����{��rS�U�.�PY��F/z���B�)5sH��A����b������Dְ�*c+V��)C�4���[�j<Sr�'��- �虶Q����R�B)�V	��'��uKŉ˚.�>��b�K,�0�����y�*�4�`Xs�n�'Z�=h�EL��0>����+m�P5��}��
�d����`���]�^�ȏy�
A�Y�J�G��h�O`@�C��P.�J�,!!R�S��dr ذ@G�L�5��?��Շگ{y�cǩ��\�h��B
C�Zq�Ղ�'=}�%�G���$�7�6�
M�hZ��8@�Ê/�mA�(�e��$��E�<E��'ǚ�Z��ǟI�^Xzb���8�t�)�f��d
Ť�0>�5�ӗ��=�P.P��$�0���<���Z�	��  ���'��p�nÈ���ϓ5��$��		�9zb�.��q��ɹb�* ��ō�9�Pp�EO-��2v��)2Jh�����-�M!ʀ"���a�S�7,/��RD�D!=�f��0j�4���[V�Oɸ�h��Am�t�un�9��2�l�
���N��5�<	TFU�RI\�$"?��\��j�r�<���-]�jp��$��D�ӂR�U����,zd���	���H����*1�ZB�Q�  ���Ѯ$�ݳ�O��2�a�Pl��b��.G��T"OH�ҷ�04��S�*S�1���"O�Q9u��5]��p�hH�.���`�"O^�bf�ݧZ�V���ɋP��"O�H��ʔ�^��`̽�7"Od�Lޗ+3Z}��]"@ΡS"O"��
I!K#�`R��#5RD��d"O���6vH����pъ�x�"O� Q�Q�9'���b/ݛZ݂D�"Of`6n�-u,z�S0�ȋ��bR"O�x��*�w
.89�,Y�C����"O�heͩW�T�aRj�7l�Y�A"O��ԮQ)p�$�(�j �M���I�"O,t�G��5��1���T31���"O��
�C5I���g��!��i��"OA;`@V�}�|PKtf�,놹�:Of}˧��5ĸ��I���s7���P#~@Nux$��uQ(��¸�!�Dd�h�ۇ�=7�j����B�v��I�f����Q�ӗ
����0ez�W�TdÌZ���*�,;.,(�R,��°>Y�ة.��t��!R�P�Iա���|��iԉZ~*�!e`�V��'��@�3* !7�����N�I��q�%ST��e�	�+���T!�J&	~� Ҳ)K�(�x�ΟT�p�t�����S�����Ǧi�*���i�Q�'7�͹C _;���`fܼi�>)ش8r�# �F�rƔ�G�U�!l�O�(�I���JA ��I4�Xk�	͞�� LB�8B�	Pi��P����,������'H�J�@�&�ru�Bn�u�<x�DUn�OrmȄ	�˼�� C�o�T$��D�:���VXX�|ü�6Txx��A;,F �u��g�\}����HO\$�f��)Ъ�n�$8�hl��D_.n#��(Õ�HO�h9���q<:�#�ִ�v��)���!q���{˸h	��B�&w��j��i&�,2�/�)�U��	�G����¾
�!2cB�${��6��=�@�7��9BjT��OW����w���hF	.+aB�*I�V�Ȑ5��%�D�;�yb��!nK��s�H�&s\!����>� �i����Ϊ2@��cBBݖOf� v�g�}:�H�d���i�P�t�As#'�O𨩱�� [N��L��p�!�G�,@!��\4h!웜r��O�=x��(OƴZ�d��R�BaR`�à;�+t�'���J /���O� ]D�ˑ�zÑo�@�(0"Ok���*^?��JD��m�@S��	��H�6�4:��>E��9y��9"�]3��`z�n�/�yҎ��rI����O�'^��wj�N�ʒO\��'��̸��l�&Q�G��%��Is��/�\���I���yp4�V��8v*���r��.O�JT��A'�O���W�Ǘ'R�����I��	v�'��͠��_}b��9m��1QE�I�"8
�B���y� C�!��1�@J�.2�y�FIV���'�&�r1 �F�O[�ht�S�a0|Hb����J����'�(�Ó��M�\���J9G�,y0���9�➈G��'�d�hv#,i�ޔ��M$?�H}H�'D�Cݲ/;<��Ɠۖ�Ȥ!��;���£#?��Ouƣ=��d�4X���bi��H����Ka���� .��ɾ{�v���L�;�M9��Z�;��g�yɼ�+	�<�^� ��Ea���Ŕ>Six�DxBJ.z�ɢ1��d��ߨ5���[�q=T=�į��fEE�H"�Py�)�	t2�!$G�ޞ�Q4-0ۘ'ܖ��m�2_���D��-"%Ɣ PK�$?$8t� !�y��\�L�E�a!��.]	6Cǻ�ԅ��n�D�$�t7>�(D4;��ΈU ��Ej�-}�v	�ȓ#@|)�a��XPeʤ
�q8xT*r�D����A5�OxU����uUL{Se�c�:�ɶ�'���rK��T��l�]�H���"�)ڰY����Qs�Ʌ�P�����O�2/�E�`�[yfa�<� '[|rA0E�/�fHp��G�\�[֮CS�[�Ld��ք��P��"���z��ňDn�l���*
'��'����� �gټD�z���'I&c��P�<D��p(�hjD�i���[¦!�G_�
�������>1Ed�>w$�b���p��m���Lv~�,���=���?����>2�N�dЬ������¿A��5��$�9�!��ܠHՀ-�c�۶wԪYY C��nn��Z0s.toZ�kR�8��ۚq�*A��|����|�f=8��9�iȶh�j��ѣ�I�����4}�\�����7x'�� ����4�.iish)z�|tA�D�0*`b�i��7��b^� ��S����<��BX�����HJ6�0�1��a��l>�A���A8^ � ��V;Q�cD>��'[N�d3�M�U����]����R�(,�m�2Z����$7G@:���.�~�n��'	�,n�e[T�I�ɉ7k�=~��5,D�y{L?���o�9Q���� �TP3�g�<ZdI���Ј?/`B�I�s.��Y���!V�u�q�R�c�)K3b�s��JE@&}K�Z�4!��	�Ha�4`nV���N�u�.X�`��1�<���j�)�h���B��e��$R�B����v��Qd*H� x1e�ȿ����q�X�'_ʴRr�'Y���=���?J`2��^9�EA0iLw;�I6Y9��@S��d�p�.�$4��D˥��3/2���ޟT��ք��6�ْ�,���>�2O��YS�/�.��דz������,Cnr3��A*%��(��ؙ[�$�
��G�a-�
���y���'a�R�	��R=k3�B.H��u��� �LZD������?�/K ���k�#.6q{T�Q�E���'`] z��phBB�Co����x�9�ˉG��=:��[į�=21k�Nv�
w���џX���?>.�qÈݺk\��M-�` S'FKC�:�v�ֻ4���뒋�wg���#����ve���«�"�V�0!%��7�@�v㉹���D�BKдS�Y ��:��29XT!�d�R?��p��ҩ9���h�*���(�|��w"Op��5�M�S����&%�S	����ּZ���z�ٌiY�	��<56r��(�3�Ayhh��ul��!KX�S�3�C9�����ʽwi�����X�(�����	��
�2U�fcK�H�����N�X��Q��.�l4�x�Oυ���w)?cm��e�Ї��OxTR7��8���!��/G���a�	%J咂�'e�H���*�{��@�
O��'�X�cZ���pG� ��1�R����qAB4��%�#�.� �K��b>�����v|����,�!�Vmh�,!D��0��Ѱ#��}�w�#V��MZ�� �4� =k��~uT J�m�v�b>=r�͞ey2�Q�C,�x@��66�	�aQ�Px¸�'2tSjU�iZ�i��ǎy��e��@47�N��%QwJh�ȇO;���­�#�"4���@� ��t���m[��h@j�,/躒ၹr,z���ͯ:�&)N�n,j���������dχ4Cp�kэ-<\�f��<O�'Zz�hg´z�4���&�n�|�eGK�8�j�Yr��G�*ĢuA^0{�C�)� |)�r,�UtIJ��ԙERThuo׃/�x�JE�iօ�����#|B)O�(��	-��(#�R�{:�3u"O����@}������_��}R�i�x��|��Y�M)���A�
��b�D�4k
쩲�Ni�!��^�C�|u*�@
�`��2�T�`�!�$fb\�R��\%+�^q�$i� p�!�&hl��GG�.�L*�(	8[!�D�zwf �aڵW�"�Z�fJ�w;!��c���U���g�Q���=% !�DZ�,��!����|z�]����}�!�$�5}: �����6�V�H��y!�DW�L	l����C�y���*	�	�!�Ċ('�F����1Ԭ�xb��#:,!�ĄN�:���T_ł�A�D�7!h!�@�����J�|�k&"��!�!�D��zv̝P�3�Xt`ǃ�,:�!��a�D�! �.��L�a�!�D��+?Pm��+~N��#���.Q!�䏹F�!�U@J�K_b��Ӏ��#\!���~�R���&2����Ƭ{�!��#Ʌ�6$n
�c�^� ��(�"O�x�u�J��:�e��w�L�"O0H3qR�@&�9b�DX�D� V"O¡�d��P����t�>
����4"O�q�dO�>���;��ës2�:�"O��k���#h��A�!�V$v{VE�$"O�9����[�0��P;Tl6`�F"Oj�+GA�^�V��&��bDv���"O~��u �2pUZ9��e�#}�ȸ�"O�D�&!����$��x��"O@������8P��H8w���"O�yAf���3`
I{��?z:�P�"O�uJfc	�]>�i,�~���@"O��K3�A`�����R��"O���DB�	M������B�A|B{�"O~�B�6Ӽ81�G���"O�T�4dX)9R�0�늼R�����"Oj\��A�,AP��@)[�p6j��"Ot����1oR�8��Ⱦ8@�03"O8Y+��K-2��B �D� H��"OTР�H�2�D� 3�J/N�DJ0"O�,�A��#(�!�AM�+4��0�T"O~p�'*EčR��V�@@"OHeQQO],)�@9���* *��F"O@5(EO��U�Fh�!OR<�"O��Y���S�ع0@b�44O6`"OZ��S�N��J	H5�I�j�D(B"O��zq��(�5x�gڵ�z�s"O@V�Y�ppS/��0�r�Co�<I�A"��;r+�((���!�Hr�<�$�?_v�[�C�-h��d��r�<)t�ݎB�}{�'X7���J��h�<�S �T�N��#��Q� �B�d�<���@�h�Ѕ��oR熴����a�<�
:e(�BT��"%��!1�_�<i���'CKl:��ĉ_U@�QCE\[�<A�!A�~���ȨY2B�BRL�N�<�
G�B����u揧BH�8��O�P�<��L�-+� 8G$4L��	��*BR�<��eP&/��1ȣCI�CT>��W��N�<�'�2����c�T?�����[F�<� �(�����%\uЌgj�J�<a��	ʥ��L�|H[��L^�<��D��p�`Pg
�99@-[PH�M�<� R�ۗ'lf�B��>`����"O�M��⎝o
�{#"K�&� "O�4�p.
3p���/�"`!�"O d�S��d���qa	�(��"O���`M[��	Ū��z�H��"OD��(�X}���X�n�8Ts'"O�@�E�&�Ą� �	�K�L���"O���5d�<3V\%KcLG)v�֜�4"O``0�H�_%��X�� F�~��"O@P9f��F�� 6��/ �$��"OJ!`�L���08��Ԛ��4��"O�"��Dق
I 	#.��`\���dJUJM��ɋP[�}���<_9�M*�C�j�n����4@�ᒥ�Tm8 ��GH/QP�T��C��}P0�a�' ���G�+I-��6� ���a&N��QU�X�?�z6
��		�8�#�Y#:�2!�G�f�d0��{����u��"
���H�'�a�>t�'�Ϙ\aZ � ˍ�P~Z%������\�R�CU�=b6�
āD�li�f 
#u� ��7�'rN������a�Z�k�u`d�'��$y�f����ey��D
#��yA��Ʀ�y2 A�i@H�e-�L�E �$J��0>q�͂3#^z0��5Y~T���ĥU��j�
k���y��o�%�I�O��mzG�6�\����X�?�!���U�g�tI�4��7i��?�c�v�`U�WꙔp%�5$<@�	Y�O6}"ˈa���dX���0�V��T/>ݣ�W�Q��eۑ���jOt�z���<E��'>q�PiL��UYpF��K�u���Q��xp�	��0>i7��*$�)gbΗY�R��2���<I��q!�`�%�U���'#�|��T�-�̓<P�\h�iH�]�"�٨9�8\)��'���� />T�X�ECؿm���E�vq��]�\�4tZd�-��#~�"��I�@��Gp,�����s�'d���J�z�Q>���Ũm|�U�dX�M�|��'��
8fT���'9}��n���d'$���nO���c H�D�!�U�^���Ģի$��ܫ��I?`��ƫ^�R�j��'�H�y�/V'P�� �˕/�X�s�a�X���>�DH�+�`���(P\x(y'��h�<i�]�
ftp����'��� ��Pe�<���K�&LC!C̪I�)�$	O\�<iGK�w�h2�ԡE�ƴW�Fu�<�@�u϶�2�Pe����̀u�<A�\�h�h1xT�X�/�8�+q�QI�<	���cϢ�hQ,FG�L����R�<��ρ#Lı�pcU~�ɲ	GJ�<Ip�E�i;���c�haʉ��NF�<p�E}��#��jL~��ংE�<���?M��C����d�Q��E�<)4�V�;k����s���Bz�<9��_.eM�yQf�M� E#]�<a�c�T�\�jQ.3����]�<����Y�΅���H�"f(�T�<y�!
I�Tؔ�(j�
`�\�<��DͅL[���'(h�@㼟�r�Ҧv���n�
H6��u�>D�0"��jҨX7e	=���sE��<A��!�,�cNU� ���!L>�˟��{���6.cֹ�w�*<ı �'y88����}
6X�7E�$w�<����,9�t�S��~V~XR��s��������Ď1�Y��hd��=j�P R���v�Q��'ғ}9vb�6,��oE����F%*���,��������z�7�D�u_̨�eQ���=Y�J��x�����Ӷh�Rt30υԦ;�OΖ�Ld�Fm�mꭀ��~���ڧ��Kq%�Ol�jŪDl"�(�3�ծ�z���"O<�2�e�^����N^2u�^��0��,@^�a��)��/��{���)�$�
��x��_�VR�$C+`i���D?ڬmI���r[��d�N��Ĉ�-O߶PQI�o�2���Ͼ�n�DzR�E�jW����w��`���!��7B���i�aв;���Fz¬�1P���À�#O�愃@�Y]�dj�*,��V���,=n���͈�MC�%�0������'|O M���'p�⅓��Q�h&y��i���ts5fJ���'*�X	��f�@4�JX��
�D'f���R�T�B��(��P�p\��S�? �`�q�۫,&B-Q�\D9�dx'��ú7�Ĩ''`�C�H�	�Z��P��w��6ơ̻#~:�Ҕ� 3U�D,��`KhƆ���I4bAP٣)��'�:�I��
�Vbp���+z0�
2�B�6o��%���7nQ��`��{lx�Q'��.)H��t.2O�SC#8tVzYQ2��4��JRu�pغ`C�����0D��`���e�%�O�>L�bU8?A���>r���"}���:>@6����ۥ[euX��9�!�V2h�&�u��
Y|�,I�#Y�L�d!'�(Y��N�q��'D���n۞K����k�Z�;�'�`�1�i�$]��l
�drd��E��L����r�ޅ�"�U�I���kp��0�(B�	�0�:��C ��UT��ra�ʩhB䉿Y�v�JgӔ�(�M
��.B�I�n'b-�*�R��AsT�ȯ4�DC�??N�Б��z.��[���^�$C�I����E�F_�����U�A��B�	�P�f!���W��N�[$o�
���,VR�đ>�%a~���$��dr��`"�\�x�ȓq	�r` ���x����'(�y3A=QP��#�O�xT�QAШs���Zc���@�'i�-�뀬2ZLx�r�0��S��Fz��Z�阿x��ȓl\��g
� X3�Z6T�2��<!�hZ4Q�&����8�'_�����R9e1x(�r2@�b)�ȓU����<K�
�Z���l�(9�K����'� ��� �H
�"vn���@�0r�)D���-J]w^���٘SE�����P�R޶D������|�!Ck���@��8%��L�@��0=���T{>\$Ģ��	'��	&,���b�2
�ZUn=D�x�CM7k�F\ٕB"��͒��,��"����0��=Q?M[�gG ;�:�)�)+��Q�1�*D���֢�<3<���`�eY���eתj*��#�>�eKo����4Zȝ����;;�1�R�A�"�!�DV�+�@���A�i���	W�d�b	As������X�"g��{���Tg
*!��E��9+��.�i���ɝ(n���3�'ӈh# ���H�@36�N>.�ְ�'0 �ś^1�8;f���B�
6��c$�h��
�L5
�5�;�$����$i&��:0��2t���B�.�?�E�R�O�Q�R� #Yix�Wf<�XQ;��*�$��G����9	QnpkMO�0���-YV�)���O��)�����~yx��N�*˂i��l�~b����4���ܑ-��������<ALK�yf�=�BJ?\O~� �۲_]@i#S">v����P���r
�u��Wo�-:�����[w�,^p� ��)���Z�5�h���	s�!򤚒|�a��%^�ҩS欕�n��'�7�?�`�8c�Fu�.[�z�u'��¦m}�u�f�A�>uI���>[|zy@��!�Or)А��3�½��B�-(섡F�G<(x�Sp�	A�J�	���tqO�pU�Kܤ�E�?�2L�'�I�P�v���L�_^���@̃%���$߯ $�H�T�Q��1��W��y"��pX[�QY��D����m�d��c�YUdM@A�f�TȆ���K>85�%�hxX��~Z
-
/������)#B%b"�"FL�y��4�����jlx�ʆ��:�P(z�U�z���f�Ưol����Ʌ�B��y�
ň�&Ǭmi�O��w��=�ҡL��H��	\YȖ��e��lX�o��ތ�¤%	�����$G�t���lͩ)IpA���+�DM�(KtI���&Ÿk����,T�@�{�$����'�5م���M���K2�cu%�-j�[?��0�B�4�t��e�^�w�(#�(D�q�+��se�Z�R�	�퀑%,:�B��>8[�U�5lEa�E������4-@y��(��
/��y���x�<)왠n�H��]�WA��{r��5r�&AH	��(�D�$C>��ę�>�ƹ�1��.8h�-ɤ9�azBJ��Y�6dSm����������1�`�u�n��Յ�e(��2�
�~��̫!"��4��<�q�G�,�2&�M�!�J����I/?��(����+`�bNp�!�d�*3��`lW/ 2����L��R3a��r�B �OȠ���3?y�"�9G��GG
@U�k�F�g�<��V,7@�;�(G��t���ݴ��K�V����b"|O� rmQ�׿Qr.y��̈|��zG�'�$��&�;^J���'�Ml�?>:�0��Y�*g���	�'�Z%�D�o��PKU���4����yB�Ţ7��:ai�0��>5p�M_�X�6=i���#b@�\���1D��hK7J�r ye��c��!��@T��e�D
'}R��@���D�;Q�H�b'ۍ������!�!�Dقp�H@H��$X�qI��#\��.�		�6Ȃ�'~n��_�R��`hviY��bd��'�Z,����0be�P����y�'����pb��1��>.�8	�'tp��$ DK�4������-��'�V�5�K�2a��3��ݎ#�`�*�'߲\x7�<95c0'C	&0!�'@ձu��rn�lcVɈ%
��D��'l&q��B�u;����J_�x��da�'�҈`��/C�� �*�ljX��'��]96��B�p#���3�H!��'l�J�4�)�����B�'���N��d=�-rto�5,�9��':F|�E��=N���&��4K�,�'t�yMR� HH�0�E�)����'t��"����f�0��/���i�'��(:�ɋ���vK:�t]��'�=C���4_��0vj�x�\Y�'�r����)4��-�%��
����'�m��i�;J�)�
(|��)9�'>��u���>LA�ɜ:\p��'�ڢ&99�:E��B7*���'��lh��*+S@8CEX<+r��	�'����A+�hz:���B[�i�L�z	�'.�y����7�!�A�a����'��<!��3gL�k�%k,|��'媼��DL�(��=��c�=�`��'�Q�Ɩm���
��MZ�D���'ԩ�̜�I�@�e�����'`LX�eߣ1-���dd�T��	�' �j�� U|@�ٳ��Ii����'�� ���<�^�¤�O�F	�'����/F+��p�aW�I�Tx@�'	r�)��4ְ�9�kP�N�EI�'Vaä�5q� H!�
�DV�

�'*,`˙Z���t��E��  
�'D(��w#��� ���0= }(	�'�8�v�+pm�]�r��3�"�B�)��,�@��-���5胼nCt�ৎE,��E�b�y��M�.���ȟS�G���9E�-�v��f��z����Ĭ|3�kI�2���)$�ՇE~(⟸��/��<ͧ9�bٳf�6䐒S�X�D,Fx��)B��8� �cf�H�_ :Hz�U�<9Q(�x����6�tiזi
��1�5{rR�iC�A�ti�֡�����?�)�S�UH��"#��K�2-��e\�	��HO�>A9G菳Qq�:@㓤O�j1AT�O$���Ӟk6����k�!!.a"��!��<���T>5A@hʓ,�^(x#����P���`�'"ɧh���Ů�L��aEʊ&C$ ys*�Yyb���LH��|�OT� � �N�@s2Y�R�^� 'ġA�'v��=
@L�K��9O��'~Hw��0o����ێ
����ǐ|�N?E���JEej)�@ܧ���� ��(OҢ=�OM��sB�0t��B������{��'��=9r���}����G�
o2��(�1#&qOҢ=���w�ʮs��F�$�(\���|R�M���D���h��c �Jtܡ�B^�@���I!!�Ca��KN?&��y3�� �r1�U����'���"�O�#}:b�̪{��R݈:JN��L�#��I�v"�,1�kL�Ma�� ���Ο K��踕GD!JHD9eV�\�g�-<#UJJ<E�� ������τ5�|�`Ъ���M��a�T������x��)�G ��G�pQ�1:��R�C_P�Xa�A�;�'����)۶"����O��x12O>M�i#�X���ԫ�)x���4�
�	��u�ԟ(X[��N�%��1t�@�9ܸT�Ţ�5e?�Ѕ�	�z��H�mKO���$��
a�bB��,��U���_d�!'i�7UǜB�I7��ٖ#�,R@�X�+c>C�� 7K�ĘA�I�|� ��EN:BC䉥+(ĥSbM�*-h���V#˻Hx4C�	��{w.k׆��d&ʿ%&C��26}�s�a�[v0�`ǃO9C�	/7�D��l�!�#��t�C�I
�,�	�:=���yg��=x��C�I�@�6Z0B�x~�����$�C䉛IV�	�&�  49@��VnC�	��ƍ� ٴp�#�u+fC�<e
!�ǚ�1��{�b��w2NC�	�c�5����x��)D)� C�IB�x@ZP��i�I��̗J�C�	;o�U�j�].)�`J'P�B�Ƀ5�tI�7�=0����ƮZDC�I�N߄�x��*<�LI�e�X.C�g���yUCԽ>M����B�I8*��F@�TU"��#!��B�I�~)�A*��Gt9;e��L��B�I1jxX����@��st���DK�B�	Z�x�Jf+�:)��Cc�0�xB��6uJ�����QM��4'h?K�>B�	�5���'�F>{��d)򏌲W)"B��.��(� �dʦi\�tQu"O�e�W�Q�u�b#��A?���"O������wIx*G�� k(Y��"Od���+ ~�5�"A��z�"O�e���>=R�]S�m���"Oh�H��X�e踉�GP�S1eX "OD��@	Z^4Y��ņi
A@"OT�+������ !�*��"O��أ��������Tn�D���"O��AZ�E#�e�&�Вt��Ie"O�=�/G6����bɾ_��P"Of-8waQ�t������V¬Z�"O�H`�C�l�N�bw�%�>�_�ƓLs���� �l���U"�--ڰ�� Dʔ���T�aB�),�]�ȓ E�q��MJ�Fu�Й��ѡ�,��y���S���@��D�;B��ȓ���($�Fn^�����-*�8�ȓC\���Ad'e���;�ꈔc7�ՅȓlLZy��͚1X�xq+Əzd~��ȓMf��ɕ�M�g�F�Gd�ȓ7�2�YfnӫE�"���D�S��ȓ }X�z���y� \��aA�mw(A�ȓ	w@�al��8xr�: C 8����Ej���GڪD*����앥<a���s���dkG#)�l��7 �g�Z�ȓJ�N�`���
u�.�1Ei��
�'��m�FB	R�z�YT!B�6��ܳ�'��L2�&��>Yqsט,���8�'4�`�H�I[�ě�랃#B�|��'�&��խ��l7d���CY� :�'��I�T�M�X�N�;"�G�F��q�'4�b��$+�U@"*�����'���$�ΰ�x�!K��*�Z5J
��� ��C5N�[�����!JOJnA�"OR�A p	�"�bB
���"O`"�#L�G�
a �!H<�Ip"O��	�MƩv�jA��O��2*,¦"O @��$@�%��,��	ġf"O���-Aډ(���04��@"O�I��]��������"O6 �C�Ƣ�e`fG�5�*�P""O���r�-Y�"�y�E�	S�-�a"O�pℨҡ3r
M�U���]��@�"O.�3CԹ`:�TC�ʀ�����"O�A�0�A-_<���0)	
}*p�"O1�7�֝!�j)��V	-����"O�1�4��$r/�E��O�+��A�"O"a@�Ӥ- ���B?G�8ݪ�"O��agl�4"��C3A�<T~�icU"O<�:��-%h!h"��F���;F"OĤJ��L�Vq�k�`$"Ob�ySI=_���CLWq�X�#"Od1�� �`���!D͞��f�a�"Or�qGj
d8D����o����%"O��Ӏ�@&o��u�g�΁G:��JD"O�Y[s�.'�Mp5)Nv6 |:E"O�9�C��p>�a��.f���ɕ"O�{G�:9Z ��6G��e��"O���qf��OhY��� q�&-�!"O�Aq� =�\@2�/R�ZP;"O�E�3��k�<��c��D��"O��cE��&���b�$���b"O*����/��S֡O4y�F3"Oj� ��?$��̠5ؤ5��"Od!Aה-s�$!��+Ǹ�%"Oر���2�8���`��M�Ή��"O�dв�T
_?�"���A���	E"Opc�)g4"��(	�%�a��"O�]a#a�U��٢�h�1doz	��"OX�����,�����h�m��
�"OȈK$*U1h�,A���Q�^4*�"O�(���-|���֢,#���q"OZ)�����+<
A���ohY"O���� ��q��P.%d<$y "O�����"���	V��}H���"O�ݻ�(+=i X��k�g;�)[`"O�І�P���A�,��<:$��q"O������ňl+U���Dä"Ov1`U�̑����֏7T� ��"O�MIC@��D�y�JW h�@0"O�K���>a!�Y"Q�R
�ʴ	"O��{�(�6s�  �\�DF�+�"OT� ##G	b����e�U�Q����W"O��Jq��V9�a�K�K�
�k"O��:�&&L�&9[4@��]!QK"O0����В!!��66rd`�"O�&A�r
�)�֨K��Z"O4���M�c�4,r�q[P�<D���j�E���{�W�h�r�J=D���ff�0�4����&8�z��9D�Lc酋��t����,],$��'*D�D�d�\�f��C�f�0ZH�i$�(D�X
� ��Q�`�%)[9a��%&D�����|t�*d��Tf��`u� D�����6l��x!��nJ��{�f4D�ӄ�O���$�1z5����0D�, ���D����Q�,TNi�,D�� HY��-��va�Gج.��0b�"Ou��</�m���6ȶ4pG"O~�A��C`m�Q�έ?��G"OAa�S�i6nX��LT�����"O��	7k�<$F�+3�U�sg���2"O�y�oJO��h -ǟ<��;�"O�*�H�fDf4	TB|�%
W"O^q�F�U\B(k�@�e��ˁ"O\Q�d�E_rAI�/��U�й��"O��B�<Q&�*u��L\ �I4"O6�*t�ފC�L�""CU!V���#"O֍��*�?�0d�#B]*E�$Mp"Ov�0�h�l�͹R�8�h@��"Or+"�O��l���6B�D�Q"O �R���bV%2�l�hDԱ6"Ob(k@*�&R�r��됄d:�#�"OXW� �Xp�֍��9�6���M�<�#�P�:?
0HՈ�!o�e�T�<ɡk΂e�,���
z@T�:G��`�<Qc�!�r|i��P!]8T�Ug�W�<����.q���VG�
E�Lʤ�K�<	cΉ3&l���[�^-BL�I�<Q�I�r?z���	ņg�L}*�B�<�%��(C6�������p ���B�<tB�NR^1؁�u��F$�A�<��I�*zY���!}W^	1����<�w��~�
����G, ���EM@�<a��ؘ�(��b�p���:F�Mb�<Q���>�Ha��^�n �:0%�C�<1R'��'�fhaEc��87* C�<Q#���u��a�sNC�w5���F@;T����U*`�L��l\+F Di�$ D�����":>���[�3��M�V  D����#5��s�EG.�d��"	=D�$�w�;��]J�<.�>�jƍ-D�d@�h%O!�r�S0���?D���O#�PI��S&�.EJu�*D��+�׻ �ƀY](�7�(D�`F* ���)�Y� C�5�'D����Ř.t(�|��W�z^�MTc$D��Ç苼~hd���kV�m��}�ţ&D��8��	T�iz�ǟl�^�3ģ%D���"E�g}�س���lhbu�$D��rA-�0S0�u�@N��N�.��"D��ˆ�7#�͙�c�1kޤK��=D�P�ҡ�Y����@��M'��[�!�A�(�qd�F�`�� �M<[F!򄘝`P����ħp E)b��(C	�'�,�����_��0`�D��B�J���'��l��N66;�KP��E��
�'D�@Z .T6�ر*h��r���p
�'��ڤ�*�>	0���gx��#�'R�"Κ*&��H��	ճ|�%i
�'` �t�-n��I�ə����'��U�"�-w���0d�qg����'���Z�c��h�0����y��(d(�)�=+��x@$���y��l&�w��vT��*J�y�$Z&{���I�lA�e.��C��yRi�6��x�%�./}0��m��y�&O�sr�ա�͇�<"P|���W��y��P��� �:2�$�ׂ��y҇������t��+qO��Gw!��*N���J���ly$�v̟��!�� ���K�{ ����(H��"O�귯D'T/d�#B����b�"O�@҇W�j��q�@�}z ��"O։�E(ӂCI �,Ltp@��"OA�%��:W|��I�\b�"O�С5��+V#P��[SX���2"Oj�"�$ot���M9 H� "O��A1���A����I\�.p`��"Ot��k�  "p(��[ƨ���'e�a�5��]�C	��o�I+��݂|Q����J��H�d�O��$�O�}�O���'`~8JviM[^P ��9U�(0���ͻoN��+�∮n�֘�i.<O~U�Ĵ�4�P1A�;�Vl���4����fh�@j b�jt���ቷCs�7-���Zl0d��v�bɫ�$��ul"��4S���'���P�'��O]Z��"@��m{"�[��Bד��'�X��w+�M����r'��i�HE$�l(޴i��v]���rC���M������S$8�Y.�nC��q�bI�v�Q�p�	�g�y"(�X"zUp@D�,E�Ա8aF�����C1K�H�pA�S?D��b�4��!+�fO90'(��sA�e^�\��d�`3S�àX�����D�5�TK�*�+��hk���O̅m�8,�S'3�\���)J��xwj�'2΢u
���?�I>A��)D�,i�Y��,Y�KJ�2��
0��~��s�lI�Eֵ@�����1 �q�
4g[��n�T����i������O��	�f$���&�\�h�e�bf�P`��8)���Fc�o�dHHt@ �fC�4� �
�f}h��Ͽ3��څ8��ly��Q'�d�2�U}��F-₸!��$�p����un�xrNzF�'^�l P��ؒp'D�4p�'|�x�˛V��Q��3�S�!#@��t��Tj<x�'Y�n�'�r�$;�	>��PJ1�:.Zz1q �:i-�>9��i��6�+��j�ݱ�HS�.�f�3E(�چ�b6o��?��?QT� /�����?1��?��oq�}H��2;X��PC�w.4�BL�f@n���iH�!6h��|.���;XQ����Y���h��>-���Yq�C�RV�Y����<�2���F�"��� �I4c:}���� )+�Y� �`�QrM* �}�'c����i��ƒ?�O%U�Xh��ϝ��B!hqɉ�����l��[�i>�&>a�Ƚ/����vЌ�r-��?�r�i6*7�O��o�{�t�Ov�90��A:��؝?�d�S�C�i&. ���G4���	��<��ğ8z\w~R�'."�p����t���f%��ᖐU/��jj&nQ�1�[2.s���$Z[_.���80v:���SȄ���Mށ �����vF��$^�r���B?i��(�e�$٠Py@cZ�39��oځ�ē�?������§�ӗ?4�r���q�v�
M���'=�O�`�����pC��c�
ӫ��I�Mc�i��	)y�&0A�4�?�OR-�r���\S<DБa�+
��U;��	��(q�e�fs��A�#A�1�����Y�)CME
eF�Yd���g��Xp1(	���<qBmF�Rg$7�'U�$�/I�� �E�5�"�&�\C��d��g�K9��ExB	9�?I��i-B6��O�֝�;�,�G�ʓ|{�qq1CO�Q���	�8�?����?����d¤Ej�)w�Ԥ�S�c��~��On��c�.Vt���^F���.�Z��'nF����'*�'\�'���	 @ ���     �  ^  �  �+  �6  $B  _M  �V  c  mm  �s  z  x�  ��  ��  @�  ��  ş  �  L�  ��  Ҹ  �  X�  ��  ��  ��  ��  �  ��  ��  V�  �  W � % \+ J,  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�?�Њ-�S��Q $��9�3탡^�]���`i!��@mA�!JCψ�@�t-K�g��KY�~RT�����ԯ��-y�/Uf,�:D�+D�ĉ$��e� !�7�8ϰ8�f	k���[���xSd�L�p����TH��zu�蚔"Oj1����`�c�瀔j�
,�2"Oz��̊^�H�3t�- �ܱKw"O�1w��]�� E#Z�|- �"O�h��[�L�R"�D��ȹ���0����e�~��@�Q��0��e`��.Q����4?q���\�z *����S�hUz�	U���O$�T#�G��E* �Xw��s���H�'/ $�"d]	+
"=K!b�166)N>Y޴�p=��Cڻ6u"8-y�h�
t����hC�Ʉ D�A2Ƃ��91��g�	\�C�z(2���Ȟ62F��G��F{�B��|K��ݤ	3D�$c
x��B�I�O�D��oS�|���b��GM��B䉩{���RL�1`��Yi�a�+�B�I�F�r B1'�����"מ~�\B�	
�t�Ir-�4F�89��!B��B�	�!0H�ek��A9P�z��=9lB�I+������<x<ҥMɝ:5Q�T��I?7��w��!k2x�aWi������v؟ ����lь�u�I+/�Р�rK��0=���D^�n�T�Xb��1B��%��%d��yB�.��R��`�A�!UPp��ac�Jc�������`��#{TDT9c�x�h�
"O� �"n]�i���J=_�����'�!�T�%K��0�N�0/�y[�\��{�8�$��Җpp�P".���١JӅx�!�D��|��;Ƨ�A���D)���pD{ʟ������(i�@_+x�
e"O�)�AK�h� X���ã n`y�"O2xZ�"Hd�� $@b�&"O�A8��[���`"]��M�%"O8�J�h�V��j� Y��"��a8�t�bJF�5���Â߇`�����9D����-P�I��v�F�*.t�Q��8��6���'��E�D�Ww��!M������2}� 5�t��� �3�Վz��ݫr���'��8��'��盨r�������W2D����:������A#�"�7)(D���� ָ2Ȉ9A�H��X�:�	�i%��O~�=��l�� �p���q��	-L,%�3�6��x��Զb�R�25� �3�(%:uK��HO0��U]h�1R�Ԋ=d�<�0+è"�ax2�=#+h=q�L��`a��:cK�a�B䉄������gcd��W��-n��B�}!"� B��Z5�t�3vB�ɒU��L*ӥE0w���{rO��>�ZB�I%O$L�Jw�S�)U�aX�Ê�\2B�ɦq~����?g�=�b�	U
&B�I(��@�ɘ"�*�a*�C�	�)o�m���ɿa�0��$��&xC�e{�; @�Ȧ���B4lDB�&%\�JӪ��*��x2Q����C䉱`<����G�_�읲��x��C䉣7��A���*E���C��@UrC��/�f���kk�M:�ʑ�#C�I�[�&$�G�6ޔ5�NE-��B�I�j��ytJ��r�ңL�	z3���,�S�O�)�\z}�Xx%J�<�⡓wO�r��J�q/���Q�X}ΝqQOV����0�Ov�
Q��	Ԡ��N�Y��(��'�R,�'-4��H�*�S�ŝ8��r���z�#`h<�@Z$�.ubvhA�=��Xt%J���'����ȟ�1�r� >|��%(�(�5g� ,+��'�4�GxGڒ,�#SHȃWv�Ku����y�� h��ȟ@Xr�Ar"jH�A [A� G�;�Ӻ�]��D�2QDM`@bײ{/�)X4Ã!��7u�|��(~�x�G�*�@��B����M)O�QcF���4��v*�,WX4�*�U�XP{�eB��y�����)[�$�1P��Y� ��y�NL�|p�!1bN0K�֭xDϖ�ynW�gX���.&���Mڃ�y�̅�(�6|�d��'t���3���y���	%1�p�æ��!��H�S㑁�yr�tT̂�Y%'6�#ӑ�yb��!&7��r��(n�ZQ�/;�y���wj������9l�T� 4O���yB
.
� ��MO�̘i4�_��y�̇]�촚���*B䐐I�y�	�Y��,S���M!.A�0+��yRe�1`���;	�2z&
��'��yB�J�h:=Y�~a�J̛�����p>��"[$����R�;� �F�s�� �'Z�a��흻�����΍,PJ>��K��Bmb��A�,�s�o��X&�Fb^�\p���$ P
{6�p��ve2�S"s�<�!K�`�*9@ċ5�t����oy��U~��(��觏[�j�1P3�\�DQ��ad"O� ��@��#!kB�ȗ�/\����"O�u����$i�̂��ټ0��"OB�@�� ^�Зd5!|(����(1��!�OFu��j��zZ�E��鑰''Tp*U�'��O65�h�3��ڡ�����!�n�Q��D{*���d&���dy���V���$"Ol4C�W"JI�U�M+i�=�2�	l�����,��0 S LGr��Ҵ�/D����jĤ=/���P���}����C-D����h��h]��G4�X	:�7D���� =QN�r$h_a ��T�5D� �2�w�ɚw���u=
3m>D��P'�ʟA�֨)�.I�'�F���;D��5�k��Hr�nG)mz9K� .D��{��&rD��QD�]uxA��e!D�49�&.���d�,(�nM�'� D�8Z " �I��ID�ƖJW���P�;D��r!K=I�.�Z�'ţz�|�kw%%D��EG �]���はz ��(D��r�*
4W�)��%�A@\�A
)꓆ȟ"e ���-=��l)0�B6!�����D8�\��	���Ѕ#�Z���b��dG{���ܨL[������]Ot(�������
O�u��� ����B�&���Z��+�Opb�Hh ��4�%o"��ؔ�V��A2�����xr�J4��L\�.T$�,L̽����o�hib�C�C%�?Mz��A�� D�8&�V�=�����ϝ�U!"��S�{�����=OHb٫G�ܔQ�dU�B��t�bC�-~Al���ܿ�(���,
w~C��/p�*�ze��-N��)��Bȸ_�tC䉜e��=0Bb�$t�U˒��)XC�vS�Cs���R�d��u�%V��B䉖l���%BФewJ��&�F�>�C�I�a�r��0N�p�Աy�+Eew2C�	��t�B�җBk�i�@�Bgr C�ILB�Q���#(��u��7^�TB�	
h+��0����~
�E�.&�B�,d��@�7L�j��He�ğ&�hB�ɭy��+GA��@���_J>RB�	�h��E̕(�,�ZVl�8P`.B�/h���DA����bg�ޜG��B��g��E ÏG���$�92�C�	5L��qׂA�hX����.�C�I���X�g#E;V�6�׊��A�@C䉤#1  ���L��Am�:C�ɫ
���yG�I;���(c
Ж	jC�IL/&�`6���%�p��i��jj>B�I/���ȍ2��cp�.j�B�I)G��5�ȕ-O��(���J��C�H�:�P���jh�0�o�k�C�-L0u�����3 !L�y�`B�kbr$*��Ѫ tT�I�9(B�	�L��YR��/�j��ʽY!�B�}t��#��SJ�QQ��@�B�I1=&���W�� ���!'� z$tB�I��Zp�%��)J� 9�-[%B!�B�I95����M�@���[�G�SC�B䉕J�Y�%Jt(P5�ڝ�jB䉁l��sAj�1AvDc�bZ�v8\B�	�rGtd0�(Y'0�d 2��+�ZB�	#3f!T+�8a%z���K�N6B�I0\�Δ{"<x-dBM)+=�B�I�Q�9@�(	y4�SU��C��B�)� �Swk�1*�FP:CB@�H�^�x�"O���n-�5�w ����ui�"O�$(���\ev��o�|�x�"O��c�Q6:{t-��m�n5(��V"O����B�FC�`h�(��M+V�z��'�R�'�"�'�B�' "�'��'�8�(%H�T+B)\�,�f����'��'�b�'���'��'0��'Fl��-ƮZyL}�)�.W~|`�'�"�''�' 2�'o��'���'s���!I��6C��	խz��5��'���'�b�'2�'�"�'*��'�)3�D�aJ���{zE���'���'�"�'v"�'gb�'�'�@������l��`-ǼE(� �2�'<��'�2�'1�'���'���'��T��ˇ �*`���N�j~���'��'!2�'���'�B�'F�'����_h��3`�2�T3���+[M�'\R�'�'$��'d2�'H���G	����B,h��5@Q#{�2�'���'b�'!��'~��'�r^�0�H���K�2!2���
S��'`��'��'���'#��'b"���KY�uq���֒���N�kB�'��'���'�r�'��'a�+ՠ[pL`s��8sh�bh��_��'���'�2�'
�'e��'���$V΅�0_6pe&�����Ut��'n��'J2�',��'�$7��Oj�d]8�����3z�Ĩ���P!�<q�'��V�b>�:�&.�#��l1�Y�! ,{Z�jQ~r�f����s�H �48�$�ڇG�2A�(����WH�l���i��"ɼD���O��GL߶�&=
K?�5�-���b�C�9�VhI��9����l�'��>�Cv$��Z���e�&�4�Vh�0�M�B�k���O��7=�]C-�Ep�ʁ���9[�Z7̦����	(9W��98O�°��X]�Ap���:��=��9O>�� �2��(�J=��|��h�촣��ۖ���`'D��;��͓��=��Ȧ���#%�	5N,x�KG��7a/&hh�cT��VT�?��P��@ߴÛ�0O�K�LYjw쓄%Rl�$���B�ʥ�'a�XH�)�u��Ѣ��4nI����`�'�(XXt	���qA�Г,��u8']���'���9O�y�r oŴY!��C=VLE�5>O�9l�:+i��,��F�4�^�sQ�8�H	�L*I ���=O\�o��M��b��#p�j~R!#x�m8�ܟJ$h��w�۞q���&o��{Ϭ)�2E��G�X)���L�_�θ,��Y+rĊ�M� ���jJ�E��H�vΟ�8k�Ȼ�%��>>�);�lO�6=��R3"�����)�.D���цW,�SPaܶyt=�(�97J�8���>a�	��A����kğ(Y�C���r��ypd�L�8�`8)� ��7����'�Qʒt)��<2X����n�����Z(n��4����Pܭ��t�PbU-�LY��}��d���$\�a�P�̙o<�06�N�`� ��N'� x���!�U��ޣ,�VX{� Gz(Гƅz`���Ox�$�O�i�<���ޏB�:��d-�'��(J陬z[�F�'��bW�H��O��T	G&�$hv�����KSpHsP�i�^	���'�2�'2�O���<��42QK�(]6D��	G38}�!FϦ�8�ɉG�S�O �I'���6-�1ER,���Z�{>D6��O����O�u���<����?����~R����bٔ3жT��$����'�N��ĝ|2�'�B�'p�[F和&Q�� e�ϯMx�x$E|Ӣ����~�jʓ�?���?�H>����U��dtl��ys���-�
x�'8|��|b�'��'u�4��a@Վί����`>L�	�A��Ny��'�2�'�'�"�'W�*���"�T�w��T6xsG�;9�'d��'ir[���V �MRV��R�䭓��Ȕ&$2�kq����a�����IN�����I5 ,���a>
�(�կ[��c/U�g.�i�'�B�'��\�d���Y���' |�2��N�ps��KŪFwn~I��eӼ�d*��O��$M)F�^�,)���"�M��B�5�ԩr�iӄ��OPʓQ� �*�X�$�O.�)o�l�[f�S�HnB�(3���&�89M<���?!�c׮����	>E.:�DG�
Q��bO4J'��X�DФ������I�?���5f�[1�,H��ݭ1�H�@���M����?I�,������O�(h���ܖxj\!�� �l��4/�#��?���?Q������O��dMXߨ�X%�9=�x����:p���lhX��IN�)�'�?ap��
�P1��:(���U/8���'.�'e���4U���Iݟ���\?�@��;;4�`6N�		�:@i���V�$���
O>����?	��z/���+��z�
�Z�b��|R�@Ҿi7d��H(�Iӟ��	� $��X�9���$E'�<0�Dˀf�L��L>I��?!��򤁊M�ܑপ/u:�A&Ê����<���?!�����?)��0�T`�ˍ��0P��
6d7*���$�	���?���?�(O��s��Z�|z��Z�J�h� �.eĬl(2����I�'�R�|��'�b�4���ز�&|rvc��N\����n��	������t�':��Ⲭ)�)��}���gP�(��������9o�ϟ��Tyr�'>���9|��~*reO2� �C�� cr%	��٦��ܟ�'U�3I9�I�Ol��Ʈ�aWG� I:ţa��.9Vђ�i��I͟|�ɕ/F �In���'��\� >�"o��	�J5i� Ӛ#���2ĵiZ�	rH�DzܴV\�ğ��S��d�U>�B��W�WL��
��R���'�����A*��n��CAA�]V �l�^rI�%j��YA�)�O���O������S�TAX�34��i���Xv��Ɛx�R7��4J�,͛f��:�l�cQ��UE��c�G�I��e	޴�?!���?at�2��?5�O�٠ "� ov�49EA3@`[�Br̓B��8��i�O��I80P��x��Ơ>J�@+��%=��7��ON��e�<Id_?��?��,��	|��%�\�:���WI� ��	�?��)BШ9�	����'@�?^�8bgT��깑�fP�U�P��P�H�	ٟ��?)���?���8 ��a!�,��e U�
60�y��d~�'rB�'-�	O�z�O���
tf�79o��vM�,8�1��O����Ob���<����?���X&�?�h�$D��4�&#���� �.0��	ȟX��Ty��'܈��uT>��I�m�|�(�tX��i�cB�6��QB޴��'��V��R�=��ڲwsx��-)�HՐd�Σ��F�'�2U�t+r����'�?I���ʖ/�"`�Ë� r��, �F�ݖ'�'4��'<��yZc`dlQ0��<�Y(��[�"�2T��4��d���m����O��i\Q~�;n h@G^��l|7�Ѧ�Mk���?��?�U���'^�sӄ���%D>���H�b�`!�0�i�(��5�'���'��O��)�\�yr�� aԊh�D�dރcW���w\�#<E�t�BM.�)���	J�4�gnՊa	F6M�O����O��XV�<�O�LD�����ߘg:J-����a��;��	���OV��O����K/��|�Wm�29��H���i�"��|��	
��i4��0%���{��&E��yQ-U�\]�5	K<�M�U��?q/O��d¦'g6�TMA��h�*���(l�{D�<q���?)�b�'D�.n��4�-�.[�d�"A ��5��6B�#����O��D�O��h�pT?�����-go�5*# �%���Q�4�	џ$�IVy��'E�ݟ@x'�B �����=�4A������d�Ov���O�ʓ:������TDE�VȀx�E�+g)�� ���9"�|6-�Ol��<���?1�ٳ�?�J?U�K�-i�B�C��5V��\�Q�r� �d�O��X}�������'�\c,(4�-�'9��H�0����4���O"����8z����|������qǆy1F�,E򜭛⊜����m���ɔ_�m)�4�?Q��?������^r��shA=J��0힠\��� �V�T�Iw�����a�i>ᦟ��ڤo�7�����c�rq�w�i\u�-r�����O��D��P���Op�$�OF�c,�NذQg�'	}������}�f�F۟��	wy�Om�O�򄇃sL�)�ѕ*�X�K�mL7m�O0�$�O�8�ңR�i����@��ǟ�iݩ���y�tm�!Ǐ
�rh�Js�l�$�<���<�OHR�'��;��ĳ7!1,�Õ*K�H7�O~u1!��ݦ��I�(���������	3V�j5;���e��L�ź-���P
N]Γ�?����?����?!.���CB@%�]b�a��NENҡ�*{�Yn�។��˟���:��I�<���5��9��Ȓ|��C1.��Ւ�*��<���?����?���?Y�A�L�ĺi� `��WEl�;@�ۧY�&�W�i�N���O��D�OH��<��1J̠�'m��b�O�WAl�*$LA���˔U�X�����	�p�ɂ
h,�	޴�?��*6(!`%Ĉ��S�]\�Q�i���'KP�0�I�b�x�S���iOꍨ���S��8���O��H��4�?I���?���g�"M[f�i���'S��O3*M�#�	[�q��O%e�k��rӦ���<!�?8�8�*O���|nZ?)V�ə�.B9z�@���w��7��O���g�Mm��|������S�?)�I*~8��dL�g�ZM��I�&����O��d�|b4�D�O���|�L?�"v�ι ��[q)�	���p�4��qb	��E�I�����?����<�����[v�� �a1`r4�E�+^�>dmZ�oD����N�i>�$?��	*����cEa��ջ��G"�sߴ�?����?��*Ӎ훆�'�B�'�r�u�-�8A��F�!��gB3̊�o����'�D9������O���?}��֓lL`1���R��1`�n��C ��n��T���$�	���I��P{�'w>2W�߸u� )�O�>)���<	/Or�$�O���O����V���IB�>����.BF�9��*Fڦm��Ɵ`�����H���˓�?!&@>;@Q!��R5?s�@H��EG��ϓ���O����OL���O�䊷�����!'�8.Y�!� 5o2h�G*��M����?	��?������O��p=�k�F�pN]��F�
>U�YȵnN+Yꛆ�'&��'�2K�~�ŃTJV���'�N)	?��GkՔ"~xԨ���1U%�7��OH���O*ʓ�?q�f��|���~�@�z�d������Mp5�8�M;��?9��?���3W1���'���'��dEY�h�ȟA���U�77m�O�ʓ�?��h��|����4��M�4�DMI�i�Hݖb��S�M���?�Ql@%���'���'��$�O=��)-X8������ ���ئh�2��듬?�Q�?)L>ͧ���?8��x�6*L
� P��Πf4�7�@	 ���oʟT�	ϟ��?���������8����e��=&F�9c�������4Lh�Y.O.��|��$�'O�� �m���Ϣq~���J���0�Q��i"�'X��ñ-r�O����O��	�.f&t�b�N�!�Ly�plb"�b��b�9����	ß��0
QW�He�z��ܡ��@��MC��6X��t���O
�Ok�-g���קQ�E�*N߾�R�OX�(�e�OX˓�?���?i-O��F��.'D��ĭU�J�0 Z�h� ���&�h�����'�l����,I ⒢G#������u{H�d.B�1���Iy�'4��'&�	�99nt�O!؍sto�S�<|h�m&6`�J<����䓗?��A���)��p�>� Ǣ/&ѼT�GeX&Da򀐢V�$����t��TyD�y��̱`�� �(��O<w$����ᦥ��G�I՟����;H
��@��+i\ �[`#B�g�����zy���'+�\��C����ħ�?��'a\�|�C�N(N̖����zO\�p��x��'���~��|����b��$/���L^�N:���5�im�I�-����4DS�֟d��5���f�V�h�H!�J�R�R�g=���'�B�R#rV��|���-�#g��2l�?l��x� b'�M;�י<C���'���'��(��O9��+9m��`R�X�4S|80�XǦ=�U^�S�O�B�\�#n����6E���)�o؈5�$6�O"�D�O�@��CD�	����	B?Q#��%`����Z57)(�d�}�j���K>����?1��r�b�H���L��y5�Z�"���ƾij�C�.W`O����O��Ok�8L:!U���pJ��/J�SA�ɝ����	Ly��'X��'1�	�e�N�I@f�!}=ZX+�I�@@r�#�&�ē�?������?��-�%12�և2�p}���͸e�N�X�Ax���Yy��'��'g��s ۘOj�	�b��n��ly��=gFN�@�Op�D�OȓOr�d�ON��$��O��T֤R�b0����;Y>�hu$~}r�'o��'X�I�o��8cO|�5�.n�2�k�!�m�5S�Z<7}���'��'o��'^
��')�E�r���/��F8qe�� J~��4�?������/���$>�I�?�Z�.F�H����w��K�F}�7DȎ�ē�?���&%�X����S�d/A�zɎ��v�Å2I��� fA>�Mc(O�?e ,6�X���'p���"?�tc��yIA K����f��ܦi�	�|�E�[T�S�'c(�Qr��2n;�pAO#od`mڨ-���A�4�?����?��'Gˉ'3bgȚ��*u�v<��oN� eD6K�J���"|���t�ء9��طf��ZSC �
�V�`��iu��'i�HY7	�pO�	9}Bb�E^��C�6N�xi&@��MC/O����02��'>��	���I�E+�̨R��K�v�KuF�fE��4�?��C'����剨�tcaF�'R��DOé.r6-�O 4�Ѕ�OJ�d�O����O����|�u�M3|��q�7芿f���C�)�f�S/O��D�Of�D?�d�Od���(���$�9�UZg�q��������|��'��'�2W�X�������z�>�ZAl=3Rt�DJ�'����O(���O<��1R%�~j�łP[F��p��(�,��b}"�'{��'y��'/$�V>��ɋJ��i�d� >�����q��x��4�?�L>����?�4O���e%���V<iÜ��&,��e�lebu+i� �$�O�˓5cd�S��$�'���Ȗ:���P��zKXt`S앏y��O����O��3Q�~*�OU
?�D�#7fE�e\�\R"�̦��'�����r���O���OX.�x�>쪖��7�f�kI��/T$)m�ǟT�	�;Z#<�~�L�'�ε��)5~���D�Mئ9��K��M���?q��ךx��'S,�`�Q�MS4(9@�ڪ3H����h�葲�)§�?��(��PM�a@�倎a���D��2/����'��'e\�agj4�D�O�Ķ�DGƋ�Y�����̘�x�0
�>�	ab� �	ǟ��I/�����%)�y�
~�*53ߴ�?Yc[(N��'/��'�ɧ5f��,#�����<�y� ����d�Z�1O��$�OH��<q��Bn
ղ�X�q�<�������έ0Жx2�'bb�|"�'c�kY_���ҨdcDՋ���Zظ��y��'�"�'��E_&���O�е@���$0!c��X�Ge�	�O �$�O:�O"��O���!\�+�.Q MB���%V��¯�>��?Y�����x���&>�K�L$,ML!wCF�_��Q��+���M�����?���8J��>�V�F�F�<��0�%d�Y�S�Y����	���'���� �)�O���D[]�Ր�7X�ؑ�RO��EH�]'�����4HG�,�S�4��..�& �HR�^f�����/�M�-OZ\�Dg�צ������$��ft�'%�,1DD
�a+���T��#q�N���4�?	��G��`Ex�������M���Ov$DcA�K�Zw�VnA"/���''��'��T�'�O�����.�'H��Сκ2���Q��i�����V �1O>Y�	����e��R�b���X;w%�@ ߴ�?9��?I�t�O�����p�`�#[�Є�q��8< R1J-��hLb�,�Iҟ��	�E����␖\~�` ��=g����4�?�tnUp��O��>�����`rƓ[��H`��'�\��[���d$�Iܟ��Iş<�'К� ��Ks �X�&%��F�e�r�S���H�'�2�'��'�"�'ܮEjt�+C�1zg�?�v)�([�Ę'���'�RQ�$�tk@��d�/�����[�/q^���^-����Op�d2���Or�$ڡS��I�(���mҙ`w��ҧ��H<x��?����?����?��O׹�?���?�� Z��	 %
M5p�HT䊘.=�V�'�'\B�'����}B�ըk��D�5�ʾuhQ)��Ӝ�M���?����?�!Q����<���Yא4Cb$׈%:��������s�
�ē�?���}���w�S��L��$)+'��;����Vۍ�M�/O>���������,���?���Ok�Ī�b	Zq.�`�x�rcm\��'��u��d����'��Q֡�A��
gL޿al��ߴ"��Mx���?���?I����Ŀ|B���&nPd�8X�D(��+�[���S� ��y���X��T �&D�vx˅��,i�)��.Q5^�Xx2�O�k*e�HTh���Q&�"E�������
f�V}0��4�Oެ2E��k��M���.he e��n�_�v�Ȥ�ޱ`*X◄T�6�N�4��Vkg � t]pŊCl�K�Ɛ	&�էL�"�"��-1�^+#��#ck�9�1���!��lr�oӼ(60��w�ݎ5�R�y�O�*��c҂�)wL"���ۃ~��C1*����X!0A�*:X�u�"�'�"�'����'��)�2���!�#c�8C�	1��&J8�}�a��#�pQ�EFi�'��Q2��?m�̀�Æ%~x:C��gL\�0��;[z�a��G;fH��̐��{RFH��?������ȴ╫P�f���W�J�X�I��?I-O��4�)�!�X�u��ك�w��-\�X�t��
��]�)F�c�-Ѥ�D�~�`%�[o�f�'���&j�Ԅr۴�?���I[Qr^yz�dKI>�҂JҞvI��x�g�OL���O�`���W����䘟��T>E�GHA�fdȘ���S�	�8ɛ�M+�b�PĨU�9T�(;G듏3��P�P��JwJ6���f
�T4̐FyR���$���Bڴ�?-��8�!,GR�b����{Q�����O�"~ΓRN�� �j�N(�c�[
�L���ɢ�ēW���@�Bi(Ь��
-yY�h�0ȇ�i��'�哿t�4��ٟ<�ɟ�n qí�/5�4���+r���Y�mH� �:��Q��+�`�:�n�80k�A���Mq
�8�~ɱ@L<v�N#�
�48��d�0��/+^@D�i$�}�5��`��HS���h�_<c� yK�E�!�4�[��J8���D�O��S�Y�l�T��ML��ա�/���B��6�м����|h�][�쎙A��#<���i>i��y����C#��Oh���N�"Xp,U��ϟ��o�l�>	��ҟ(��̟��_w�b�'��ĳ1��(�l<S�����@<!�4(q��<VR���#+B����fL�Y8	�<��H}���$O�5A�\�h�8A�Lx�$L\C�\D[7NX�6Y����M�'-ȯu��'?Z!�qϳ^�� �c\%+��Z�'y�����T⛶k:���Ox�d�<��J~� 8�V�)7 �8�
U�<IT�G�BL�gf�%7ł|�M�;*������'P�8�z��ђDC�a~�|hЀ0���O����O&�Dӛ-����O*�S6~���Ҡ�4Y|P�;�!:M�<*@�y]��i��٢uN=b�#�l�4�ɅyQ��AT�=�}�L�B��h ��aW��PI�v��|hQ"TЦ[�*G��'h\� ���?E� t���cTK��U����������?�������iŸ.��RV�3.�
%�CD&7^!��E�9;�ӣ�?��H׀� F��Φ���^yB�C��t6��O���|BGÍ�|�,�{U��-%��<ː��:����?Q��Aڄ�p뉗J��4�V�^�#� <cF� ��T���)Y�F(!ǝ�J��@�ZM�'�j��m԰i����"�7%n����� !CZ� �&n��= �@��; � y�RG��?1��i�����$ٸ-�t4�%|�M2Ħžn7��D"�)��<a�mE	eJ(���U�#q~�yU�n��rL<�0�5e�0up4.�!8�����<��F��Iϟ��O
�[��'q�'j�h�V��(�J�I���P�3�G]���mX�@o*�I���O�m��(`ÁB=�DI	D��'1�k�C��}�� NP�s�yy�E$�?E��ބ���%��G��j0���ݲ�m��?)���?)�������(�8䢎�L��<PFKN�y�'�}�Ʉ�xc0��瀷J��������O�`Ez�Y>!���r��q���y�5���(�	Ol=aA!^�����ğp��2����O|աңW�F��y@�(3ϾYk�k\z�cwK� Sn��2�H��p���S�4� �>Lj(L�%!q-^=8FB�-��d�7`O�Ay��s�?�=	�*��|E����բ@���yPҸ�?�G$���?����?�gy"�'��I�EŲ؋	w��XR��K�=CvB�I��T��U/f��xc3�Ӣ1p�я�d�|r.O20�����u�e�97@}���Ƙ=�ZTY�"B��������I�@8d�	ʟ�Χ�����	�E?^xËV�\��$�aFR4rè��1к]��v bpS��(�F`���ʞ�b-braV7GI�ԉb�Q%2�f�4r��`�\�� Ad��5`�m�{�κ�I��M� f�:goP�=��At�@�����e!m�Iğ���T�S�D�V|�@ ���ޘ1�x��$�y�'�^�0� ��
�#	X}!��ɡ�y��lӒ�D�<a�/X8 f�Sҟ��OYr��	�aR��౥�6d�4���%����';"+I'R2j���ϑG>2tဦˬV���m���%��0���H�R*;�n�Eyr��%`x�F���*�4mЅ�3�nX(���68�A���N{���D1?v@1��F	]K�'p@9�O���/�����;|A ֝>ٺ��Z��ןP��	�O�_�\U�F>a�m�Т#?���4��$�x�S	-$%L ��N�v?�5�G`b��>�@l�֟D��@�D�T�GT�'~�J�p�t��W�(�̬2�!Y��L`t�J-�՛�*�OH8��@㦤����wX�Rͱ'��@�򆓩Zt@4ȅ�5�2���	 ����f.T�# ��T����|�ݫ
/2��D�Y�;���7ԭ,rv���"����k�4_��F�'�?�d!uv��u,�cB�p����s���O���d���`�ص�C1\K�Ԩ�, �1O����w�'�@�	�5Oxܪ��y:ʩ�2��k��@���'���a�9�V�'���'�R��~����<p�ŏ�Fp��V�ؒr�i�`-��Ǻ[L��Ò�N�l>�#?A@N�q`���Aƙ"�H�"ֳ2��EQ�ŋ�	����BdI����.\��#!扞Foܴ
��R!\{�1�� �!	Df���)�.�����M���,O����<���y��\������u�W�g�<1�A�)RB$�$`8e�2Q�2�Ӟ|<���'��'>�9U�'��ɋ̒ �Xw�0�r#aޣA�$l��GQ0+�8���' ��'ib�K�H���'��)�d�F.2�"DS��RZ~�hꢥW5(�VE	�*¯V��-�u �..�����е/�őv��`��{b� �~Ad��î�2 ���BC�*�M�F8O01+�"D��f�\�����+�,X�m�ވ1��_�:0�DJk�̟x�Im�S�t,,�D�PS��5M_��C�m��y���U�l��Æ0I�p��!3�y"�>	(O�B��_����۟ДO���Ӄ�>5݄�QElѪIK:��2�	�;$�'�����DL���6�j�Q�Ν�2�<�'�TqI�T�0��C+%>܉Fy�'P5�Dԣ��0b�쌲� M�-�3��\�DO�9¸��w������I*)n��D�����ߴ�?!*��aX��DE�])��B]�pA�%�O��SH�'m�����N�H7f,�D���=z�١
�%ț��~����F�P����W��%~�X�'���a��$Gy�}���O6�D�|������?i���?A�L��Pό �U�	�{��Dش�@%l��Qq6J�jS�P���z���.�tc>�$M��Xx�$+dQp%��,y'�3N��Qo\)C �py�\�g��O(6�u)%� _��id�L��(��aC�O���%?%?��	[y.�����.�%�V���A��y2�[	A:А�N�7C�t1��	��O�|Ez�)w��dȾC'��K�MR�q?"�!׎�Eh��O��[Rg�E�����OX���O.����?��U�$B��v^e�笎�
_�<9��'����cؿn�8���ǅKF{��F�,�<�3W	4Myx��g)ݼ$Ĵ����D>���E�D�B��hOR�A��ܯ ;�����1gzVx���Op	ف�'Ǧ7mH¦��?ْP?m��K޴ms�A�\I��%K&�t�	)h|a�A�N(@��	Ȑ+
(KJmy���Z}�\���g����M3c�:��I�ғ[H���
�?���?9�Hԕ ��?�[� �C�JŧU�ߜ�2�iI`�(:s�f\�)�
ӓT$�A7�.��0�2�١���>/(@*��J8�Tڡ�L�k�th��G}�'1����>��_�p��$�Ф'2�Q-/[�@2�"~�
��<��������'�,3$(î�ܘ�@MR74Ԍ`��hO>Qk� �d)�!J�@�E�TqQ>O�UٗB㦽�'��e
ҏjݝ��ޟ �O���{���Eߚ,weA�0�8��A��!]"�'7R�K�"F��1̡f�B� �����8�'?�$9��0�t53�"ޕ�Dy����ļ8�P�	���
��2u�֝�2,8q�j[�G��uH�K�&B�� dDˋ+�d!a��'�26m�O��'������6�l2b
��XM�p��������$D��Y��ٶ*��T�1ǉw��s�'��u�LUl�ȟD�(�cb�Q�#+�0�b��S���M3��?�(��<zS��Op�$�O��R��]@$��R�g�!m0֋�5��HTG �:]�&BH(j�0��?��|��)h��(P&?U�+!.J"MK �c[�|�L��b` �+���Ӆ�܊'M�9r����ɪ|���mdY����2v��xs�I�xl3��C��?�D�|���'�D	P�م{P�Q����/#`0�'�8)�a���	��- �K�y2�'J#=ͧ�?�C����w��R;�xK���?i�� �2H��)�4�?����?��P:���O�L�dr�%��C ��}L佺��6Q�spB'&����6��<����}~�CqN���dx�&ܳxD��u��!��Q0��A�3ړ{�\�9�&Q�hK�@)�+�B	N���4���I�pBH<!��?q,O� *�9QA\�*��u��|B1���'j�A�y�`М%xP��kڭ+�Xp0m�&�:7�Of�O�)�O˓`�ĹA �i�A�O�X1dܘsh��~� ����'�B�'�r�ԁ��$�'t�	�Iu��PC(���Z�ʛ@��[)"�i���C�^�ݨ��&uʑ��PEN�I��H-}e��# @�ND�$��K��Uh��TƧ2�Ҽ�ߴ^��)J�팑��^��)��ϟ4
��PZLȁ1rO����9bX��<��Yy��'��O��
f����&��j�<D�q@V�8't���7ړw
��BΆ��L���$`
!�^���'��'�6"}B&-BK��+�ctB͉f�	Q�<Ivˈ�7��X�4�U�$�Dh�e�<�&^�By�6&�8��E
&`G�<�U(P�+h��{�M8k�t��@C�<�����j��P��`����9��Xx�<ac�]�J�� ���<B�	���DJ�<���W�v�9��9
3�\�*I�<����0�b��rE��E��!¢�FE�<q扂�(���f�]
uK�K�<�%j���p�r�+T��!A�BD�<I �=[>@��&ܻiŬ�!'��V�<���� ��S��7`;~�!!�R�<�d�_�5��ȱ m9J�l4��&Q�<�უ+��-{�%���)���v�<�L��9��H�M��wy�X��l�<���T&-�J�Г�p�-�Ԉi�<9ujÌJu~Y��҂!��,Hd�$T�y�	�� �ɖ#A�U����0D�(��b��B��Gd�&.tb(��(+D��
���|���Vkؑe�.�;$�;D�p�mZ�n(J׭Ը�
DX�.%D�\A�(V�C=VA���P;WxS!I=D��AwHF?*@2�*I�ӧ�:D�
Ai�Hc.��iK�]O E��2D� Q �6x�z�a�I�z��E��0D�@���O�nt��Dȕ,
��bdA0D��a�Z}����6-�6{v�����,D��{�	���k��ސ"<B�B�8D�l�6+��� �
g,��2�5D�Hxpb[�(�Kc���G����Ee9D��#�'"�Z4�u]�mdx���f7D�8 �������ګv��������j��wV^��!hM'W,ӃF:�?���%��n�t d�Ue�����<��['�^TcU�Z�/����-�v�'?f�XÊ˸o� �4 �a	�mk�k�u,�����g�'��	�U�L�z��a� k>9r��0��5i��7<O>8p:3Be16𒀁F*�!���1Y��I�)�i��	P���,��G��qa��ַ`�i�gN�׈O��Q��
n,t��	��c��ͫ�2O,iK���[����/ �b�n He�|�'Vy�%��n�n� vJ���l��(�1�?�e��8y��p����5WO��Scd��<�c7��Xq�u�VI�a��X��?7�K���*H g?X��1 1)��I� N~���kP"Қ`�d���\"<Q1��l� ��<���b�	0Us��"�&�v��?�<��+��af�H�2Ҳi3�\�>�b�4 \p!�%�'ej�λM�`  �dp�8G�ָ*8�t&��F{J~
P�z��c���6�л�)!�G���sB-5K�x��Ý�*6m<+���$ϑ�3�b@Jpd��=��K��z��<�q���X� �S�p�� ��W[�^�Z��_=�}c ����d��v٨�
!��������M[��,��|a��>ɰKI�G��vS��,�F%�\y�@�\�Ҳ�
�L�2�PV�A��6����� գ���I�"��5��z���e@j	�x�شt���#Aη��ʓ�~��� �C�f��邭��@)�,�'��+Tиc#�nXj�	��͒;Bhp�F�	�/\��!f��3&�E8Cb��A(N)Y�%N2V�#B�<9�<OH�ӛ�����F�1HC��M��I�/\��$P�	�9X1q�\6Ey�K�'L�]i��'�D{V2q�߸Ae¡�EP?��m0o�W�P.,}�`ߪ��):p�d�w�lN����<��됫 �(��Olݪ��L�B�D�9Ѷ��<O�2
s=��G�]| $�gI]]�	�rY@�AI�e-tt6����p+�=DA��]k}��BD*a� K�Z�T�p�B�8TB���N0��@�)C�HS͟``+�k��N(���J��q��L�H΅��ץz������'��u���L8Qz\�sG[;Y��p���D9
;n� t�;�E��5@���L�*kv���G֝7ք�X,�_I$���hW��ɸ�Ί0[k����\��'�ڸ�e�
��l4��L�*�P� ����f��Fy���|���M�j^P�"��'�0�/J�&��,	a��#O<�'p��kF�ٲ�9���h��1�-OB��~��B_�<'P����1�*����^L�	�q$*����N,)����w�S�I�p���a�*F�*�1�Ƅj8b5��)K��˓�?�ɟV0HP�P�i7&U��'Nlk�FO8t��A�-R��1�2�ԖF��A��ʟ� ������M�OM��V�Q1|�S�jQ�B�ܡ�Q�'�hd��E-�(�*Z�Lɏ����(�UI�@l�e�IN�J ��ɞ��O@-��t���-}" b��hâL?1�`P�gO<1��#dR�v�����d,*���+���M�]���<��A��0�3�
M(�0x:E��k�%�	(����O������Ǽ{�H� m4�d@C�\���j�i
C�I�>� 0;�l�4F�����L�c�tچ&�a�͙�C�%N���`�[���'��b�'�� �����Y$�<��`�/TN1҅�4%��%�4#�\���0E��`��IQ�Yc>�ڀ��#F�Ji���Qf��1��O88`����	�Ǔ)��+�bD�|�
�t��BC͋t��{r�h�		
��9�M��R<*�k�bL�f����	}�J���Q�qŚ �C��8J�ѱV*��Gi&�caH�lv�%����V��$�,��$��Q�g�6_��V�^�z��ܢe�Ed�u�̻A��O
�����W���?9���p0�yۂȞ�z��T䘰CK�'a	�P��O����m�X�K>����Z��cB2?q��rcgI	H��A�e�E}�� ���(;�N��4nUnT���'�Z��G�'c&AR�NUX�N�G��S)���tfHZx�U����Iɤ���'�Xx�#E�+h���b�Qq\PA����~��#=�;P�����C�Bb�����w��^}��Ѧ�~&!��j�!gM����'������?��d�I��F�ͫ#M��HZ�W�� Ҭ�v~���$/L�3�I-X�{q��b�<I�eK7>8Jq�(�rɳ�V�=F�'Vrȱ �'�Rl�օ�K�`��b��|�g�ŝEh���`����%X�§9FZ�[�O��YR�@,�IU�d9��(�'�#O�Ȼ�#^�@Նѐ��'�<�`��[��TPe-y{�)����w�~�؅F�0�L��1�Y�#ZY��}R+Ԩ��c��"�+ժ����ac֝+rM���?a�@X��*&.���&)�4>Jў({�GH��'�����F��l��-�`	^e�8��Aϫژ'm��AΩ^atY�����8*�́Լ�� K9� ={1k��?)pmrBj�Q��S�R��������Ĩcqa�������9�O�EZ��l ETNp:�
��w�$ d���(���«`��	�G-�i�	��H1C	�#/�|�(�I �G~���q��t�s��T�����A��矬"zڅ9ঀ((���f��O@��s�\�f�� �-掬 �i�={�K�U�8�����$+��h�빟�P¡�&o(�$[��U�O1O��D�Yǎ�!-H�nF�	�DHQ�������^�ݒ��b̍0�hO$P����Z���Q����`�$�*�l�1y�"�L��[�|ј`�O��R�l{޵Pnr2"}Pc���fዒ�3}�(�8�l���|�g}��C@e&��P�H�D@QS�$.��XP(@����	`a`�`��'�re�c�MG �(C��DJ-*�'>�A�
�w��#]._J\�x���p�$V�>�	"༑� �|������H��tY�&��LM���+z$���@�Af��PlI�W�<ͻ9N@��RnZ�5?\Iw坋k�Ez�=�	�/�Lew��>c���a�30��=�D� �VeZw�NZ�=��韚<�@�5`FD���IXPq���h��M)�ݸ����-L�yb���L�\)R��P<h���%w<�EjeJ��.��� �`ͷV	~`F	1����'-�84Ȝ<R��\YW�]���R"Ѝ��d\7 Nd�9��UT[�ȱ� ��%� ��h�QNd1��>O����'[ȝ��"�m��YJOǲ �B�'�R�S'�=��bB�T4;�
`�5$հ��͓T�b,Xe�/O�Ջ�OS/~4����ɰB �7%j(����Ʒ:Sl� r#�ObY&�ӝo3|\��W*d�rȲF�i�A�eB��T�J=/ZIB(óD(�I�cY^I!�9D,��<�O���r�@ҁ/_<]	�b�yM ��@ʙ�8.4<���õ�(O��j�"9� ����|�k�ʕ�TC́.��r%g� @I`�� K�S�DAp���0���q�O H�G$"�a�fX��� c�@
(���y��'?�*�T� ��� -h3�-���A0$�� �'���7d&�$a7Ah(}h��}�ўx��	��L�:
�Z�áL�����J�
P8Raf3
��SA��<���H! �!nv�T�<��*�"TT��-���]#uh�I�N�A~P�ŭ0� �$^�d>�%��\�0�B5葞�.I���z�\�NXB��		���p$J̻v�"?pLI���3h��2�.�O�!� N���I��AK�&\���02�r���'�m�����|�p�h��3��0�����?��8w��;��)}Zw~����)�T�̻([H�"��p��e��n%U�r��9��Q�%˅4c(�(O��O��#.�&2��:�a �.1*�	m� +������C_�I8(��[�����6�A�X���'����8x|<U�`II�_?�0z�ڌA�����'�r��U��Wf��H��R��������݋_�.e ��ڛtZ)�3�دP���$Vޥ�6@��9G~�=���W?�\�+W�=R�[A�ϑF���RB�H��刱CJPk��8�l]v
H�"�g��IJf!����5� �LQ�,�!x��	7��(4H+:ړ(Ӕ$�q N`��L��"�'B����^sb��.8Q�fuBQ�C�]X���7#Ǝqi��cNt5�U؃�]�F<}B��y�v0�mU4d
��C���0�`1�{�DAҨ��|���g=@�2�e%� 03�aM�N�����cY�	s���kT��U�Rj�=~��۴Xy��Ī{��-k�a���������	"hO�@�������B�8~�!$��F�(^\!��1JH*T&܃��+ѡRռ}#��*m���Z}���HxBTat�'P@[W�S�V�B�#T�dh5
4"\��	�b�9`Â_�d�� �7��R�c��!'��|ر�CD����3�L3hpڙE|�ǸO��q� 4��k^�y��A#m^�MA��7?q����F��4�dE�PY
|rr��o<Qi��&��V胳{D�|q�Z7�hAp���Lq�8��ͥG���:�c��<��ݠ#��]x��ʌC�Vx@t��a�ɜc��X���3PCJ���n؄=R�-��T|�bT 7��(�M��� ULD�S%V%0�ʈ��b��yڐ��EG�Ta&��� ��@��eT��O>�+���$>aRm#W%I.zo$�Oڎ��Ѝ�	E^Rq
��U\w@AB�꘻H]��R�-�yX4É�2�y�N�0#�5X֦Ǹ阼�7�M��M�b̤fJ�[1,�w����U?5ZҮט�ħZ��`E%�57�^p �-��d7(ۖO��bA��v���Ʌ��(cR� ����a��|�^�3d$�2��8A�_?���b�c�̑��2?�v�yS�N?o>}  ��U�`@Ȅ@\��0<y��!6.�� Zd"�t�V+�/M��$5�L4�͹�*܁.�$iӆk@qS`�ɼ;,��@�-8%3����Hґ�B,���0Zة)Qj;`?��W�<u�J�`�")��X��� w��QPU>O~!��+���0����0.$�k�b_�#��%�e�:Q	j��HB�V����$@�C�t!I�#E/%OZ{u�Ş>
9bF�4���Q����w���̓&t ��:Q���t��QP�pA��X��$����ITB�	���m�̔�n��-Z�&S�|�&i{���<q�lM�l�r����	����Œu����f��g�l��D�EZi[�RT�����)���dY�-JP���>{d�)`RK�&�����O�m�U��]"0/�f��O글�CT"&��
6	�\����"�<���F� C�U�2c��1O�T�6k�6��I�p�����{q�
	��h�*5i�Ji9�GڪL���"�y �Q�������y�A�54$����hj��ԭΐ/��\A�HJ��������ڏ���I�	0V����mê����-C��z�a�e����C���m�'�W�m�剡��J6�\ܓNwr$��G��[Bl����H�.�Ȳ�X_*	�P��Ap�	�
.�ʶ�H6�*��K�t�>�� �$u�ୃE=/�:�&D
x8��@&�\� ��g�h��x;�I7�$�vx8I��ӄ8���y�F҈j�$�8L�`߾w�$���(�!2�(hR�|b(�#6���YBO�Mnи;®/0F����ϻet����cl�� g�=<OB��L?J�~$Qƞy?l�[�/Ċ
Ht���FqI`O���C!"��	�b�˃�ʽB�I8&lԮTD����.j��Mz�M� &Ni&/5?��p[�+ʿ5d��
�'��a��ڰ[���#'-E S'4����=���U?7mQ2)1�t)D��U��M�E/$�Q�$��^�t��[�ʹ��� a@-9�	���>Q����gX�7߂�#.��w��DX*��־!��}	�S?#=�#�~��3��	�鬡��HI�'k`$y �N���
�1����+�!cL�E�5�*B}l�� � )�P 1��K�㫉 �O�Q���'p�*��fi�*u�F�X��ɮ?T�h��L�J��XX�B�D��lņT�XM��2N�<�B�#�y�Nt�N�"�;_.`�j��я�y@�*%���P�j�x�BO�.�y�A҃����)M�>�,�c�@*�y�ۗ'� ��G�"d(c�i� �y!N8��Т�C�,�h��Z�yB(�.C���au��"��R�-��y2�ǛW��!+�D�,�\�y�� ��yBG�;;j���g�&Pt�:v��+�y��ݘ��͒�� ���e,�<�y�*�		��P�⋻@�v�c&dU��y���6V�.�;E(�eId�x��^��y暛4�t� ��+
��J����y���{����\�	�^��$��y2���	����́	�8��C���yrO�H��s'�R�, 3 L��y�nW7x�lhH$�������8�y҄S�=Te;��]�
�,�Hv`�1�y�Ə�VJ�{foK���e��yRO��r6d:b�. 쨄�4Y�y�$	��:բ�E:�!c�I��y2E��b���$�G1g⨐s��y
�  m���9��iP��'wc���"OB��*ň�.�(���N��Xj�"O4�p@�¼D��	z�o"w��y"O�qb��_�a�,p�᧐�XY*�"O|�q"��4���8W'�;��t�"O�yp��i4���E�K)Z��"O"�S���6Q��ͰR��|$��)"O����/��;d/ó4?�X;S"OJ�S�YyP�0PO��=04y{4"Oj�®�l���Q"�K�Z"̥q�"OAkUт]��2�F#t$!*"O
���;ݜ��T��2p���"O�8��AQ�'�pp�P�>��p�"O�9yg��&l ��&�	j��	0"O<u��߈���E�WCN-�6"O� �'�2O�~\�b�$M����"OV8�@�ߴ���+�/]�^�Z\��"O(I��*&�P���6o̫'"OT�R����y�OX�8\8�"OvM
�ɞ=�@�ծ�t����"O�("�O	�dS��2��T�m��TPF"O��*2��
���kԇ��̚��T"O�l�1!I��� �F�R$�\�1"OjPX��*������A �"Oj����F��� р4�*�bv"O�}{�L�4�;�dȪ��8 F"O�T��C� ������ݻ0��	C"O�<s���PD�q�gMG4�@�"O��c��oV&,�gX���"O̤�g���zRؓ�셃���c"O�8��Q/&��`��� �$h�U"O�i��G��b�,�
%	�:6�(�0"O��2�'A�0���WȜ���x�"O��B���y����©�5s��̉C"O���� ���cH����$ $"O�����g������e�j�"O��I�@� >�����F"X����"O�,�$�?����'ϭ1y�Lj�"O0ň���7c ��`�H��ZU0��"O����I�E���ƃB]�ɛ�"ON=��ġ&��h'��m�9��"O2A��ɽ^:�a��H[�"Op��B��&�RpQ�Gf��|�"O�s�:j<����Ƈ6HM
�"O��S��LH`qa֊��!&a�"O֕je�ؒ}�	+"��9���'"O�%�qg݀&?�X��Zƽj�O�E̔�XS0��$`�6����$9D�tPU$�.\D)`Sa�1\@�9�.!D����O"A��1ٵÎRYx�d�"D�<�$v�$%��̇12Myf�!D�pK�N�(Plx儇���� D���Ƨ�%F>=��bC*D��3��<D�l��M'|4A(��L�����l7D�� A�]%t�I0�l�_Y"���4T�d˂��?qa�pQ�.ݠy��	�"O�t�b&��p&��,���J�0O�)H���$LI{�-F� ����`JX \B��6X�ʩЀ+W�=qU�6��B�I�[�.m"i��Q" ��P�B�I�?@`�����!)/�� u�<;�B䉷W5�U1�@<k�n}��"�� �B�<��T>Q;��Ǝ��Y�@�Fz�r��/D�Jf��P!�:&:����.ʓа<� �m����Quش� � ~�D��"O�� �.�z�\�1�Hςa��"O
ذ#�^>�Q�,�o���a�If���%G3F�p��S�Gp��n/D�X0B�߃t���s��3PEZT,D���բZ%ʶ��F�Hj��"?D�D��'B�w�:4��T�V-����;D�0��oSV�x-�
T)j�����5D�d�"�w7�����" ����Ӥ!D���5n	3G/��k��$�0��n2D�h�![Y�p3F!��Q�]0�2D���iX'-~Uل��.y���0D���AtpȢ�R�?èXi�,0D�̺�Q�W��\�%У3�����#D��ѢO]��r$sDB�-Ԛ91�,D�D�U'��x���c�f��i��4)D�(�! �'F<���G.�x��)&%D����aC���M¤�A/[����!D�D�$�S6Ou�A��Ę:7�<D�p2)ޝj�F�b��B�*j���P�;D��5D��TJ<Ѐ� 
J�`B�4D�({����Z�J�,]�"r<��1d3<O�#<���ơU�Y�8c����!`�<��I
�t�0DD:T`b�
Zx���'���(v&7
�i�&�!|<�X(�'_BD��b��(x�uB��V1w�\�!�'RR��TD�?�mP�ʎ0J�$Q�'z���g��hm.�1C�6�H�'l�3�7p{
�hp
˪WU �����)����qg`|J`�3zK`���-�yrN��h�"��QhE�q	� ��Հ�yB�Z�}�)іFƙk�\���Iץ�y2&
!ߦ�[��nO4��"���Py�['��
B��b��S���E�<qV��"T8DQ�%W ˔��AD�<��h��ݚ��0a�3�\hZ@ D�<I��K=T��!�ǉ�9z�����V�<!A�]+MkE�T�W��6�k�A�S�<��ͼ8�E1q�O���h#��P�<A�"͌y��T�a���fVZ���
�N�<1&`_�3[��Ut3 $ ���G�<IE��5X��8�b�a�\�0��K�<��A�:������_;�,�pk�\�<�:�p� dŃ�h���p���9�!�A��0��DU�So��͒�:�!�$T$V�8r�0t�tk�sj!�D�1}���b,�I`8&
˜4��y2�	'���b?�UQ�Ȓ}�PC�I�@8F`��e@�r�ЊQ��B��?IS�p(���%,P�s��ʏQX4B�ɂ'ĭi�DJ�20�2���$j?0�'Ta}��w��C�X08�e�+MoD$��'�yq�ß���	�s��Jd]9�'ɐ� �:%�Z��g�ؒz ���'M�tB@��_�X���Eݥ%Q�I!�'�>�����?��%��>�r��}"�)���4>�� ��	O�i��y�2��?x�!��U����E�Īn�v�h � �Q�!���tM"����1o|Pb랾di!��"L��0ĨY#~|-h*��.[!�$ާq��e��U�p��ඃ�#)�!�D���~�+����{[�����i�!�Ez��r�"ǧR&Y	C<M�!���9T�l1=٦-��;��C�)�  �3d@�!�zAX�	�	VL ]a�"O:�E��	f~��Fƍ^_��D"O�`Ӂ�09�T�@&�۶6;\9��"O�Z3�A�DDp��@�-~=j0�"O>�C�ժT�(�#�C��tG|��a�'��OD���?/���e߄QG8љ�"O��aP��	k# :&���b:p`j&"O��d ս�Ѥ�C90� ��"O���b�D�?�TaQ��#^�l\���2ғ�h����S�dJ2*^%p[����
�!�T5S�RX��*rV�mYa#C,k���(�ORɩ���#S1��#�
i��!U"Or�@��Q3`P�"'�*i
���i)���K������HE�|�T���ň�u!�d��P3�)�jϡp�A�ED�(k�!�DPF�0q��/� ��!��	� �!�d�I�L:w�Z�j��@:����GI!�$MK������t���:��� 9!�DMnŴ��B��#�I8 a:!�d��z�*�B�f��&���
�!���Hv�X�����WX�pb��vL!�ӻ�.����hG� q��ȧJ!�����Ӵ	P�w0F@P��w'!�>*�)�oF�t-܌��dՇ!�ē�?�������A����Û�ay��i)��l��
��S&�5\�{"O6T:�?\��v�\� < ��"O�@�Ҍ�S�H�!�ϩL'�U��"Oȅ���< rȡ �/Q�0�e"O����#��Q�l�T��2N��U2#"OF0Z6$H�5�2��P=��%ZP"O�d�e��q�����aH"W��h��"O0<��M�!e�%����5~�X��"OVP� C$#���B�t�^dCC��^�OBtB��	46����a�0��}��'��Bv. :����ۃ,��lQ�{�'�X�fC}/P�0���5�A��'�"��� ¢E�i�A�>0=f`��'<�Ea1�)%���Ô����'lY�Đ�pFl��a!��Vh3�'B4(X����"u)�.J0xn�`��O:�=E��N�a�ã�@7t�th��I��y�,S���d�A� l��=	Ǧ	�y���i:�X�e�%l�Y�k���yr�Y
jx�k�aΤfz@�u��"�y��V�iõ�AN��R�͐5�y2h��%�|x�E�=�:�h�`;�y"F��J9ZI `�A�*.����y�h>SH|]�eCޝ�!��K]��y�/I$x��H� ��0:2��e�	��y�źY����ĽKp�X����y��p��b�K�t 򫇼�yECB^�u���#HD b"h�+�yl�8V��ӧl<� 9Q@��y��E�hϔ|����;0�����y"DϨ.��X�˒�Dn49P���y��I"_a@e�f��@f���G��*�y�g;|$(�Э�	9�~����yb��!7Fp��L�6�%�@�.�y��0Kyd5�W�!	�R��R&�y�eSp�ip�?�T��b@��y2☊<�8"��LkN9) L�;�yR�I) �d���h�:>�9ِG"�y��� 9V�*D��"B�����y
� �`��ӈm?����oד�HB "OF�� ��RX ���O�D��"Oн��Q'j�i�aM�`��5P�"O���A�K Vh-0R���8|��P""O���P���(Ԝ��ҬB�ceX���"OD5A���t�"!X6���#9�y��"O$�yã�8t����cBH8X�"<�2"Ob!�TA�;4Z�]X�b�7�L���"O h�D^o������7��,S�"Op�a�3���K$݀�1�d"O�]	�	�2`���	
b4�XG"O�+0�� ���%	L#��h�"Ol��cz�����,�A"O����k^tU��f��,n���b�"OШbtH�-&��[��0`�`"O5xS��3��D9�r���"OB�"a.�2L�Pݑ���9 �H���"O��&m��[r���Ǐ:��̱6"O�0���!X*m�F�	\��L��"O`\�(v�I[�f_}(U��"O�Ic� Y�H�ʔrQ�H�Uf�A��"O�K��ܩc(q�R�M�=Uxyi�"O��
'A��ܣ偆MU����"Oj哐A�*S��,*RaV./LxQ�""O��;�%� X��7���lH���"O�*�%�L)B�6Yc "O���ȋ=��i
�?H��"O�Y�ثW^�X��^�a$��"O ��菖#���# Ǘ�iE,�"O �A�%Ƽ>�d�q�	�a3��{"O�LAw�6T`�E	&�@�"O�%#��'s:��"���
^	�C"O\Q��!
�g���ؖD�/�v͘�"Ǫ��SS��1	�A��;hԐ�"O�D2�e��!��͔w�niʧ"OD1�ve͖�H��1k߽86��B"O~��B� �P����u5[�"OT��� 		F�Pʔ�+n�i��"O.��䆘�|�2¦ʣZa����"OD�RP�ګA7$Pj�#VOg�U��"O^\ ��� E���2b�.N�X��"O���R���#�^�Z����i1b"O^ARa@וg3�Tg�%�H9ɳ"Oԡ�P	P�k��PCa��~�� P�"O�Yy������j���P�"�:"O�qꅃȵ�|kc��.!�XS3*O���� �P�(�����'�0��/����:�ѥFrt��'褜R퀉
r\��'k���q�'xTl��u�(0��kH����'FZ��A$G�`S0.�ft��C�'� عЃ
�yM"(K`E�b�X��'�ȅ"5��Pc��'Ī@	�'����6@��5#V��2*	�<���'�tȒDޟ1.$MPa�M�}���"�''�`�%��:Y����Ɇ�D�{�'�X��#�ΗgB���舽h����'T�4yW��iYD	�WdG")����'q���U��%���۟v�lX`��4D���� �r�x�(�h�64[��)VL.D�laU�3mX-k��?4�2����+D��kӇ�	5�8�*ĵ���f�2m�!�D��d{B����9������ЍT�!�DT?І� �_�lI���X0�!�� ��Y�+� Drlh�.P3e�d`�"O�%zDe�2"����ΜK��(��"O��#�<~T�P��S3[YZ��"OH䆨8�D�0�16�pИ4"Ol
�b�;��	9Rh�R���""O�����'�5 ��-l�,r�"OnUBU�Ť##���B�Q�� � "O詢 �Yr���
��
�>�2�IQ"O�L��C�-K�ڌ�����g���j�"O~��g>O��Г �.l�
��g"O�	�
K�cG��a�M;�P�a"O�����"7� xa!.��`�4u+�"O�)�&ݙW���u�<2T��"O0��$�d#Pq"�O6'/8��"O�y#�0N�fP��K�S���IV"O>И��P/;�`6�}�D��j-D�H�С�4٦]7Ȑ�j��tZ�,*D����][�%9�cP�>J���$D���1G"F���hA@C�j�[Fc%D�(�f�X����b�'NF���=D���Bd���a��²e�� ʦD:D���5�4[@�����{���j' .D���I��%^dp3aN�����˵�+D����7"Ąc��*)R驲.*D��3@19�y"w�\����ن�'D�� C(.���tnZG��Kǉ?D�����"�teٵBס WX��'�<D���/��wA��;��U�L������8D���ƃN��!�ӠN-x���W�,D��N�bB<�d.��%ݼ�"�,0D����H��Qe6P����&�tXF�*D�{���&.u��ö���F|T�k26D����'_~�A1�b���n�r�J)D����WV��@ -ߡe.Q*��;D��Z��KE�M+ł�,T �1�e4D��4oV�'TD)�4�Z )��Q�SE4D�`q��F�w���+�/y��5��a<D��F�TI�I���z�ᒭ$�E�ȓ3��DV��~��d���Gw4m��5��u��x\j�Y�Y� ���p1�W�����T�C�pS�I�ȓ#>lB6���H��	!"�4��	C�݃��˄$�@3K
���ȓB���ee�5{E���
:>|!��s(�<[��M-@�(M@0���+q��ȓ�4 �&ӷ=נ!���6P�D�ȓ� ڄ��A��k�,��E�>��	��ӆEH1�T8k�0g&m�ȓ;K�r�csIJ�5n+N\�̆�)�]�o�,?� ���A#D���ȓ
��$-�=D��aD���M�Na��c���0)�1y���	 ,ϐp���ȓ@����5	�b�hY3|�B���� �gL�8�TMA�-�:5h�ȓ9�ZQkᆃ&�dQ�
�94�<��ȓ-7D�R��Y�dU&-�̬2	�	��}&LeᰥA
�d)FHݪX�����,9Z���)d$X�&j5�ȓe�<x�����S�8Y��-�^֢��ȓk�ܨ�i�76,�P'h֗<@T�ȓ!�V��`�*v��Li�hR�nF,�ȓS49���I���G�5@�X��K$���H��Y��p�oN5T�����Jq��	���'d&�-B@��9t�ć�S�? ���Pa�"k�5���۪ o��ʥ"O
��L��u�Ӈ+	9��j`"O��S)��;<��&�H�J�PP��"O�4�c��	j�A�D$�AV\��7"O�d3b,��z�0hAE�0v<p��2"O�1��Y�؜@���ҭ��� "O�!�i�[����9�Z��s"O��$T�/���g�$_�&��"O��*��W���+�ΐ�U��a��"O9+s��%�e��̒z���"O��2�@^<�HY3��D�k���0"OH��b��M��"Pn��`ꁳ�"O�L�$���n��e�%��s���"O~P��#�"x� R�n��`�"O 5;�ǧb�zy���u��Y�"O�X�Ҩ�u�����.P�Dy�0Qv"OJ�8t��/�	XbL���5"O��w%��\�{ ��
 ����"OxIר�&c���ǋSx�T��"O���!�_�����CČ����"O�I�dM�P��u��bRpqލh7"O"%�V�*T�e��X�Fi:�"O\�@#��D���-mPDA�t"O�-�p
��9��mҲ@W�5N����"O
����)u�(�SfFBNhCt"O��`�g@2L��l��n���!2p"O����J�c� �+ƃQ�0����"O�E�B%�t���1�tͮK�"O���֫ƺA���ȣ��
�вv"OJXKD�,s����EB�8��P��"O�%��&��^*�T#�Z`$��T"OJ4�2J4�1��bP�)Ap"O@��,^	a�%b���=>F�Ё"O҉A�&�M�2�!C'^-J4 "O٠t �^L�H���"#@�A "O2@��"U ��xg���4"Or�3$�R�<N*)���o�]�G"O��pD� (X�F� `�_�{�0T�"O(��!����W[�5ˤ9��"OLYZ�C~�q"'��%��T�"O�hk�V�:�&E+3�W�g�f\��"Om��A�0��� ��%�(A
�"O�(��� �bɠǄE���yb$�E��L! �WU5����ڦ�yR%ڄG�%�!>�<�񋅚�yr�.
�H�� aPՌ%�b���y�$�"q���s.�9yЭ�4F'�yR! !.,X���C��#�e��
��y�/�`�}�r�ۊ{3������y��@,j�pa��Ɇl��<A���y�"�tu)����)q�Ʌ>�y��9�,�KD�S�$?(0"aQ��y�'D 2�H;W��h&�Q �I�y��
@�4�g��2��G�ŷ�yB�&Y͚	2�ϴ9��	:�����yrM��]��`R�à4�4�����0�y2��U��p �AX/Z�;A�Y�y�aޙw���څ�@L���1���y�!J�@WĹ���u�l`� ���ybP+R���:�kHg��  D*�y�h�orl)&�>[- yr���9�yB`��R@��!��AMXE�J�y�H�"���j�1J2(�2)��y�ػq�kUo_<
����6���y
� P�铉���6�I�߮	�J�!@"O�-x��%���'ܵh�v��a"OT��5��F�hm[�c_�>ܼL��"O�iw��"U�Y:���lپ%i�"O�=��V87�|��' $L0A"O� ��ή=��|���6N .I	#"O��*tO��KA�E�e�bߖ���"O,1�c�N�1�� �td��n�A"O���B���\O���b;�����'��h��- `6p�gα\Y��*�'ʒ�J�� D0e��n�j�XH��'��������Ń'Đ�.�tt�
�'T���MȜW��q�G�&]v*S
�'� IȂ�X�E���d�ғTLl�	�'��%����S��C��$<�Z��	�'/Э1B'�O� �
��?$���`	�'О�"O2)������P��'���B�A�6���k���
�ƙ�	�'dYI�� 6����aM ��lT	�'���s���|�B)r!"�2p����'��3I��"�2`R"ꇮ�HY{	�'�~rd��Qo�`�Y�T�0#	�'Sr!��$OM�t��BV+���'� W䐆#qġa'�̟:�~���'����u#�B��9�O��2�nT!
�'Pv����`�����Q�%c:��'u�� 1'�"��Us�@�<���'�4�F!��tT;�(�'�t�r�'+Lh��d<�{fg �.P��'V�T�b�"<¶�AWJ��j	�;�'�.��G��8����fgO2+�'8���K�GQB���툸e̠Y�'��j��=iZB� fO"d��={�'��!t`oBdJ*f��A�'�Y��!-w`!`CEĔr�(���'/d�K�:ݨ��z��Չ�'i��E��|�Rm�f����'b�X0�U��b�I��^GM�A��'ΤP2�k��Vr4�� 	=C��@Y
�'G�APAoL5P.HI˰(@�=C��	�'3�4���;l`>&[��'Њe@!h�!#�9�g�Є (�Q��'(j��S���c�>��
�JReh�'���6(�AϺ�x%)B��z�{�'΂H��ʜ�����(��c���'FR��E [�y_�THŇʙ
�F�a�'��A���

B�Ѡ�b�wF0pz�'�����"��1������7<���'lԈV��xOdy��F�@�Z���'��QPѤ޺+hx���F)'�Ԡk�'�z���E�%
�I�0�O<N>�+�'4@�P'�K�䭱�
 0�&���'���	 ����A۷���%����'��h�a׮��7��%�|��'Vؼ��#ǵ"eT��l��<��y�'����P�ֳM�ұ��.�#lR�
�'y�H��-Y
J*ҡ�p�)n�mJ
�'�L���LN�(�0x�W@U$#� ��	�'�>eD�� I����T��'�4�5fW>.��li%F�)����'���2`U?S�VY��
L�zRR�b�'�z̒�,�x����KC�AV�z�'_�,�t��j�Cƕ6�2=i�'�f���g��<�`QvH	�-H
�"��� ��
�Vi�q0�ŉ�	{�|P�"O�!{b
w;��j!nGfl�Pr�"O�������9����eZ2"O(��j�= �)��<I��<��"O8k3#өc��@�
ʑW��ty�"O�t�6�nb������Ll�R"OD��2��^l�H�EGR8�z5k"O\4c5�нP�LL��Eګ`��c"OP�զ[��tCE��B��"O:=�E蜍8���1D�8V@a)�"Ob�E�#Nz���!�L�	G"O�<9�@<�f�*�Bb��c"O m)���6?�0��-� Z���"O\��@*Uf��e��*�X`d"OTD)���9�v9��iR# �6 ��"O8����d�1�Bi�2��!p"OHI��ML;i��)P���f�t)�"Ol��ԇS�Yy���JnLA "O:���d̄|�h��p�צ,l0$�`"O�=x�m�o��xiP�ƌ*�ȸ8�"O��)0F��z�1�4"�b�|ڑ"O a�D��n��������� "O����R�.��}84%٣l �1Q�"O�px)K:L�[��K�F��*O0���/£ �� ����7

F8�'��������e��M�H���'E��aCO�OHM����Ҁ[�'
X*DE!'t!�EDܪ7D���')�h�AX�A� � E-1Z�~xC
�'0�s��͆k�f��G%��M��'ČS�*��x�l5��
� g�T�'�&Ecv-.qCR���n�����
�'��݃�
�3p��juj�3`l��
�'�8���̈,� )��ٵ.�J
�'w��(VD�7+~r0��ߨr-r
�'QL9�u��6��y��,�>�B�
�'jX#Q�K�}���:�+�� X���	�'��8P�0a�zK��XD9x	��'���Q�� ��d{6��<$Ѱ	�'xu���Ǯ�H��HZ��� 	�'���@�</Q����V)��%*�'�����L�'��5�#�{+*���'��豣Ꝝr�ȑ�C�W]w}(�'�J3�Y�vQ�隣�ՈMl�dP�'�Z]S����e<^�r�bפ7Ж��'_b|bd��v�~�#а\�vL�
�'I��_�n�`���J���8
�'�L�ҥ�Q�T\`��'Nv!��'��������>��H�+��b�'K�5Ao���Ml���`�'�"I�ˋ�J��e�krx\�
�'\�P� dkd���0b��(!
�'�"@���N_� �
�^�j��'%ȋdЪw�q{��G�� ;�'bq��=��h�9���c
�'Q:�s��k8��iB�SH	�'bny2�4}O�:p柍{"�0��'�"p��f� ����W��x'��
�'�q� ?j:������=�����'�:��R�D�d��	g=N���'����"E4��	;A0��S�2D�\��_�E�,X am^�4n�{��#D�|��(��4Ⴍj��}a d�d- D��q3��5g���@�X�6a�ш=D�� ��I�R�<�y�%D1 9X�"O�P�7I�S�t�0�����"O��J1�ګ��iYt��bO�ŋ�"O�����A�L�1����{>Ą��"O��S�&�C����!K�*����"O,���T�z^�-qB��kkJ�Qw"O����&#^�X �G�(bXIy�"O
�i��b�|�	Γa��J"O4y�+^�boJ a�BH�.Bt�D"O��! ���U��	x��IB�<�1KՎeY�Y����un�D�G�<qrN�%:)\��d�D!u�GM�<yrH��.�����ǔ!N4urD�D�<�☔ ��4"�f���ӡ�CC�<1$lʺp�h�����o_<ɻF��V�<��J��	P+��>��e��Mъ=!��X�����T�lxP�0���2!�Ѹzl��B%�=a�2���˙�.4!�䆩�$90��3y���03�X�i�!�� Ԩ�;%�v$��D��p!��B�#H\�&��`����D�!�!�$�u��X�A��K��a
fD�0	!�DǎR���oD�e�������9�!�͸x������Bin܉W��&�!�d�91�2�A���֕����2�!�DX�RH���,��}������ٸf�!�Jr}ѳR �Tf8e/1�!�DE��Q�+7�]��)'D!�$x���;M�D+�i�h�<�!�D$*��ț�f��[�z�I����x�!�$�@��#Ǫɱ4��9�� �i�!�$�#A���V%��h$���!�Kx��� �G;R��V�:%�!��8�U�]����M�&�!��N�<�&8A�#�7t��L�ЬM'1�!�����+����s�̽3�膔u�!�D�*_쌊
ל � d���#�!�$��)����wV%S�B��T'ϟqw!�d3@{
�E _��TZ �F15Q!򤏮6��TD	�g������#<�!�Y�:x����}~(�d�N3!�	�C�$<녋�Mvx	&(c�!�d�3����5$T"i�q��*\9nD!�D>˪X	@�Jt��c򊃅6!���'V�	&x���r���k�!��{o�H`��utԘ�t���c"!�D��8f��hQ�E�z���W�^
!�d�(��!KX�[��!�aa�1�!�d	�n�X���gL�;�Ȅ���Q�L�!�d�6%T<(��/�捳��2W�!�
�p3�]�bLնu���"#P+�!�$�	[�"48�%W���lr���c�!�d��Nj<uZզ�1}���3��9X�!�d��e!��jBN�;k�dq֯��i�!����g$�v�B�)h�(v���P!���x=\z����v�9C�l�7!�$]��D�:� ܘV����c��Y!�J2kI|0�f��v!��z�����!��

s��@�C��0�tMhU �1JD!�)8EXq��(I�z�|x��K�!�h�Tr�L�<�@��G���&�!��z� 1��d��)趥[�w!�D�/q%�z7�T�`�:�34CT�?!��3(�� �2ꏔPw�혥���T!�� l9fAN�c|xq�%@.@ %H�"O<%����9��(!�&Y�H""O�9Yl�c�8���cFzc"<`"O<��d��K~�	X�b�)FE�0a"O~�#fh]6%�n��'� g>�=�`"O���w�/si�'/c9�"O�#�M��Dd�K��ڭ"{t\��"OLA���'U��Q ���.���"OXX�CJA0vK�؃��Sp\`�7"O���橒.Cz�Q�#��FD��"O6����21Be1`��u�$"O�m"P�@��
��G7z턘�w"O�qJ�	��-�NH��5OAz��"O����m�^�䐰J(H/�$�"O` �bo���:uN�8��"O�M���^�ua� �x6��"O��H�.ЌC��T15	��/Zyx�"O@ ��*�L�%�߻8��T��"O-��;Ob���Nd!�"O��r��tq����(�nx��"O�D���M/+�̌� �O��ɺ�"O�0!�-�$.�Uj&�޹��yp"Ol��ܯ%�n���휸h��)�`"O�`�@Y�m>F��w�T�Y�2U�q"O ��5M�0xp�Q���ʺL�|˷"ObD�ƩK�|��U�Q�G�f�J-	�"O" ��dX '�4Ӑ���	4�h"O�e�p�U1*��e�[%v��"O^�[r'*��p ���$ 5 E"O�5�7�ȶb����#ʪ���C"O��&�׳'� y;F�����hc"O^�p�K<5
���B ���4ae"O��b��sP@��q!k}�HS�"O� �"B�%d�z�qj��}@)Z�"O@-3��I��P�ID�|$��p�"O\�I�9Y�r@#���'t�ı "OL��M7;D:�H����1b"OXҗ�EaN�pGLW0@�&��"O���4�{�q#�^?P|�i;�"O�dCf/U�@� ��7ς2l�b��@"OȲ�b�6!��w틔k�<�G"O�hڳ�����9s�Sd(���"O�-$��9g���*��˺6X�xr"O�K7��7R�R��$��V���b""O(���EP�W8U9qJ-���	�"ODX� ��~ � ��+�T�Y`�"O^�#�	�/Mc�ݣe����l��V"O��7AWA��h��!.$�X�1"O��ɦ�ʲ'b�M
�jۀ	��zB"O�X���^Tu4$����(m��L�"O.�b`�ߡ|;t�ʄ�� mJ���"O~	*@��0^x2�� +G:j��I'"OF��aT�8TK_�5��"OH�I3c-��b!���,��]��"O�L)&��#nx՚`��Zk�S$"O�H*CDH769̓��N�9t<�"O�Y��E�Y�6l�'�R,V���"O\yj��_�K��]9iK�e%��av"O�s�M	�ZMb�"�*Jz��U%"O� ��k�l���
�r�L��5"O`i8�(��S�|]�Q��"R�J�"O� `�o�q���`ޜW�+��y�fJt4P���jY�h<�B�n%�y2�ϡA����EE!f
��CE^��y
� �a��˕/����K��8o4(I�"O���3�%|��U�G�Y!{2�\Y�"O�U
$]�<R���k�ˠ��"O��:f\�h�*D�a`2b���1�"O�e�S�R"<v�`�	y�Bpbw"Ol [���}� h�92Ǽ�"e"O�$iC*���0+D�P�}D��"Or�����F��Hr��$	z�ä"OX��+�b�Zh�d$��e�r���"O��)�� y��h'�0���$"Ot邬Q(�4�G
Y;�U��"O��C�`��c�Ċ�HS ���[�<�a�ߛ{�Jx�aO��7l�a�u'J~�<���7�U���0J=�X#1A�E�<A�h�q�@��b���u�lSBK�|�<��L�6��%�`�Mf=r���w�<a��S�RM(�)׭W�z���XAh�\�<���$����jNs��2�AO�<!ª9dA�Tʕc 3��uXgI@O�<)En��G �2Ѡ��z �l]J�<i�l[je�]8��U�ڲ��W�Qk�<ɤ�Ff���Ѧޙ0	&��K\�<��f����ŁW0v�xF�n�<9p��&�mhA��`��Y`W	�k�<�!.H8(]~���I�$� (�e�e�<1�EؕIv-r��)x
�%I7d]�<I��ξDtt}� �
�eE�)��iS^�<� ��.J��C�G�9YhP�F[�<)$E�|P<@@��]����C�DR�<ᄂԩ�� 
�Ȇ o��@!�D�H�<)�M֦�ʑ��!kj�<���\�<!�bL7|V1�G�,�,0i�+�S�<���=Q�p��nD�/�0���)�Q�<	�iE�w��1�� �,�~Q`Fe�<!0c�0�8�c iΧ@�ԣv�RJ�<!��@"#�@p��ɚ%)ƀ�1��@�<yg�.q6p"�M�$��I��jJ�<��CҤh���"��eu�=3g�z�<�&DV�<8�e�D �J*A2�+�y�<ё��Z:x��C�&�>�I���u�<��I&HP:�@ _Q�P�0�S|�<Q��@�J�V!Af�12X�PQ�]v�<��cҾ�`�X�F��R���G�<�v�G�	ں�J����0$=� N�<�t�ӵ~�:�'?~(���O�<�"#,���Uh]�{��	RL�<I4��.�Kζ[����KIE�<q�H��i�J��P�t�!��#]e�<���
=qs��` ĮK�ИA��_�<��+�&h<	�mǫ0�T��
e�<񦇗!!�`��.�|�F�� k�f�<�+e@�"�ɇ�8$c���y�<�lԡ	��A�F�p.�T�rE^q�<A�aT�v)�hS��Z�B� <(e�Ck�<�"i$v����٘����g�<Y(W"���s�],ZP�y���\�<iFw��h���ׂ{�:�Bs�<Ѷ���h��SH�5~g<��b
T�<�O�[��5�)�ˇ�&�bB�I�4�,���w��i�Ą	Z�2B�3kF����]�[a��wN_	��C�ɷJ���#��cUx�S5��C�I�3)�0zV�FD�[ģ�pILB�ɠ]�֤��g�"F���GJC�fB�)� 2�+�"mL"1�O%���0�"O.p�׈ܘ]�p�* ͂k�����"O�m8T�X*j��a���ZJR"Or�y�^$q�<���G�Ue��Ф"O�{��%Z�<��`�5OF%�0"O���W-)Y) P�Ǯ�-]�	��"ORU!'߅�qʂ�J�~ �l�t"O
�+p�N +���˵A�J��!��"O����^��a!#��(���I'"O�� #��E���¡)�1	� �b "O��#p�I"c|@�CȂ"0��e��"O1�R�O�D��͉��	�WX	4"Op�fKM���`�V�x��	s"O
�KB�s{��{�h��$ɉ�"O��ڗ�K� ���&��6���[�"O�����ˮ;%P�c�	�<D� "OZ(����d��i7�
]�(��f"O�� �)mk �2D��X�j���"OP@s���)bH��������"Ov	HBߵn*HE �e��L(IR"O�T��K1��-)!� 7�
Apg"Ob0��"<��%ḽ�A0�"OL�8�&FzOJP�1j�,�2�{6"ONL�b�Ё���JBƚ53�8�"O.Yj7A�!HJ�Ѕ�&lv� "O��j�[M�R�	/4��"OXL�uʚ�s=�M:a)����1f"O	I�C�f�|��W=6�HL�"Od��Mڃ)~���-�,鈌�"On9cLܘ\�\Q��4� 4
F"O����eF�s<1��̕=5�BEA`"O���Yz0��M��0�P�
3"O�ej��8H�#�KC����T"O̝� �7T��e��`�	f��:v"O��� ���o�LxB0�	-�8�p"O��y�ϳ
�Ȱ��F��nȠC"O�A��E����5�\T;p"O��ɂ��6"9�	��B�?�5ks"O�Qp�P�aք�c'�I57o�D�"O�<�%�]b $P �)g�\j�"O�d��?u�� �oK X�,A!V"O��Jr�Y�K��]��M��W�P��"OV��p�E�S�U��*�4��F"OPԋi�F1@qb�.2�Ȓ�"O�:%Jܬ"*~��A�G,U	�|�"Otpb�kWew�0�!Z&�A "O�e��㜈;�ӀO�-ݴ�5"O\�r!�9�@�cb��_�����"OㅺP�#@�2$��y���ֱm�!�DX����Ëm'����DHӺ�ȓ[㞌z�B�v�nd���V� ��ȓ�����HφW��j�Xb�r���r�p��"4�	XQ2V4,�ȓnI,�A�-
�""�Hbc#)|� ��K�Z5YbjY�q����ʶ ���5j����׿Mp0{p��o����Z*p��!>a,iKWJJ-,'�}�ȓu��0��D�.���@	,M�ļ�ȓF�q�"n_9$�Lrr)�'�0�ȓ}�h��� �96ȹ��#"w��i��9���Cգ{Aꌉ���,�����1��MW%8䙵��W�� �ȓs=.��p�Ժ-�\�7ػ_	��ȓ/$�Dxtj�5{�!b���1W��(��S�? P��r��,��iGF1x�ΡrT"O�]JQ���,��#� }�&HQ�"O��D�l�P�9Q�$��`"O���7��"N���&'�s�X��"O��3�S��4=xed[��]b"O��{��W�g�*����
C��Xip"O�<ӆ�u<`��"�Q�>I�"O��6�*y�1�B^�_�bx��"On$��rYrR�RT���+�"O؄(���,��5S��B*��`�B"O��'���#��yS#�{�u� "O~���o�Jfhq��B��E@n#D� ����?���5`�	h���;s!D�8B���A�P�CDgC�Q2J"D������;6�Bp��DU�m�tE$D��XA�RMH�}"!�u�j]�A�/D� qu�#6�²�*�|ъ��(D���hA�1�`�2�JוD"��QЏ&D�xS穛�]�P���X_�l�֨(D��q4"���DU3EZ���Xp�)1D�� W���O9�9�"��8����E/D�ԣ�Y���F&D�qB�,@�9D����̐��097� �|�dK1A"D�$����1��@�s/D 6|���o D����&W�'E����D�;4� �0��>D���iB.p��J0�B j)*ȉ';D����D\�� �(dz-�{a7D�<s`�/)\b�Y�ӮW�ms",6D���#\�=W��W8lJ��.D�$:@��������@�R�H���+D�\�o��''�Dr4��>%Z@�ZC�-D�x:Sȥ2�uڔ(1s6Is�,D�,��C�-/��K�͛N��Qv+%D��p���~��V�� ��)��!D�x�����Q�`ë|�6�b��*D��r"�,���8�)��e�<��"�&D������T��p��� 8 HX�@2D��cff�;E���0qZM �5D�,Z��7�x �Ox�&U�cF4D�h)�a�$:��A�K�RN m�@#2D�����O86��8b�H=�RaZ��1D���p*�!f�\��g��8֌��6�-D�`K�Q{BG"ѹl˒����?D�d[���6%I�Aê�|M���  D� ��͓	Lv>E�B�D�jL��#D��& �� '�8���R�i�,�R�!D�������T������!�D��.?D��z�X�z�[`�AN�$)�;D� E�O"H "T��Q�"�l��&9D��hrIձ<��)#�K;,l�',;D�xb�'/>���S�� \X�qo=D�Tf)�-�@��c��3p]�!B�)D��b��
1ᴉZ� B-#�4��%D�$�aK�Nx��%KT1~�A�#'D� ��Z4l1KUH��v�`�9co#D��
�m�*(�Dг�
�����k/D�P���ѓ&�tۗ�ǉH^�Iڔ)-D�D#�!��a��M����_Ҭ�[ �6D���'�A�� �U��pTe�df7D�tքԠv�pl�#��v]:&B)D�Lh#��E�p��A+� N�
(
�'$������x((0���@�>Hh�'�ށA��(`m|`PthG�7�
�*�'���b����;�27�\�s��� \��ć�Wy\Q�擸 ^�u�Q"O,���.r�&�QE9��9k#"OV��4֋Nl�,�uE�k3�90�"O��I�8��,�d�E�vyr�At"O�<J��� ��A��eY�V��b"O�u�t-^5FM~5�B��$37z�r"Ol�Q� �)��g�Uv�LQ�"O��X��*��	M����g"Od�Uf�~Y��(I�fb��#s"O��;�ٞ
E\iIU�N
FZm{�"O�u��ꄔE����A�9��,�"O�x��ؚ-0,�q� �zN>���"O�����~��� �"&���"O,YjtB���Wǉ%\}�]�"O4�X5db��9sv�L�pl�A��"O��1fK��9�����dҐm<�b"O6�B��
4Rm�T&���w >��$"O���]��H��F~RT��S"O�S�I~���#� |��r"O��з�]4�&x�T3
.q�T"O�2 N�3o�	�ĀP$u��`��"O����,W��)� �(b���"Oh��g�j6>��7`@s�HL��"OR�qd�:-Aΐ��K?ՠ�"O IK¦O?|�b|�c�/p���Y"O�I�*ϹG���PaIn�� �'"O������\V��R����"Ob���I�.����ӳ!�J�XS"O��A���J��)�g%(�6��"OV���S=c��亇��V�"�i�"OXIX�E=l��+7@�*���"O�$�c��t�ZqpDMHf�x"O@�����r�Z0j�.$]��e�"O� �I���5䟤}\��z "O��)��k��XpsLJ,Qbt $"O��0�\�ж�F,.[��!"Oluq��W���<�q+�/
�b���"O�Z!�^������8]D�� "On��n�"��s���/VQ�#"O a9�U]|,���'�$�\Qà"O��f޾n�X�w��E;�U��"O�8uAT,|v���?!��Ԩ#"O �Z�	?_`��k2
$�P`3D"O�u ���3*��h�EjD�g6��b"OBd�q�_�$��Q�v��3h"��U"O��æψ�'��SG�T��Q;t"OXs�-/�0����(�8KR"O��KaE�9lr�e���E�4��%P�"O:��&+\��� FUw$y��"OmX��_���
ĢA�o_�%�"O�[�.(�
�{s+���y�V"O����I�I��a���,$���A"Oxl;��g\t}�qI�e��0I�"O�34-	I�@���G�M����"O`�V+���8�@���v�kt"Oꡓ"+� ��G�J�蹙�"O�؁k�_�v���-Sx
!`�"O+A"z�rl�g�E�Iq֠��
K�<a�Y�_Ċ8�͌=Wl��	�^�<1��(�@�Z@@��R��ٚ�N^�<�e�ZB�a��7'0��!�X�<�TP���V�>������ _�<1Q&�+���Ӑ�#��dk��u�<D$�
f@ �r�ԪeH����t�<� $	��S���5�g(R3{�X��`"O���� rtz�9a�%lV!؀"Ob1A@�5H$���g�2>㊀�"Ov�:&IR�J(��C�DȌ��"O��c���'��
�葯�l���"Ob�#@�ӭHV�|� ���g�@D�F"OXšf��68w��0AE�B���A@"O�l��&&/���	��h���	�"ONA q&�|I���Vm�S�ei�"O�<s�늶S�	!�B�Yb��2�"O�I���$�&�sED9WW�yq�"O����ޗ}X�� �يPBJq"O\4�q)K.�*4�A�*2��4"OZ���J29;`�
�R'��"O� 6�LD���gG�w��=�"Ol����Чo�֥:+�N��9BA"Oz}�eD(t^ �KG�<�blY%"O(�SJ��o���b�P 8�l��"Oh��ę5��12��0��I�"O0lZ%#������K0	�8����#D�$�v(Q?8��}y���0j:F��k-D��@�e��2�$YrjG�j�֔�@H?D��q��&��P�W%y����Ei=D��J�h�X�,z �d�C�I�#BLX����ZNbİ��M�C�I'gx��P�ⅸk.p�ӯP<q�JB�	:ac佉 �)D��IrV�B�	�1��HI��	OQ��*bcG*tz,C䉑#\�Кvd�0#"4��@>E�C�ɛo=T�q (/�TM͉�0�C䉘n��;Cj�k4��"D�92�C�;z���fB(+� Yv�ǪU�C�ɽ?t�1

H�8��@,Q�|C��<^t���4�<U��QZ�EJ;<xC䉔(�<�1��mۘicɆ�&xPC�	}IBhB�fJ��t���o��&\C�I�d׮(��)jr��s��]��B�I�c�t��
�.r TX�AS�[�B�ɏU�Ҙ�	I�1����^7/H�B�	 �LQ�@Z���a���7�C�	��{�mP,Y�����[���C��4L6��W 6���;�囆h^C�ɩb3(AdLq:�`�e٪�DC�	�(A�H
��H�6p�g�#M(*C�I[?h�A5NT� ��`��S�.C�ɯZ	6��g!��a��	ǯUlC�I�4��x*��S�V]l�0O��VBPC�	S��I���]������K��B�	��z��p	1l��er��^1��B�I�1@ָA�GF���y4f�d-B�IP-"���ٌ �r��`��BS8B�	��������	B#|,P��E�^wB�I~@&��dJ�n�lH"`��G�C�	�>��QQ�.O3{WN(��b[;��C�ɦUl�a��5!��y�bAZ�WkXC�I�bq�}�6�V; ��"���j�ZC�I5YOt,�ǁP�bO~5aC��{��C��/I�֔Y�
�1��DStEM���C�����xS�^�m���k�KS�B�I	��1������˴��k�<C��1���c�=8��B�]A}�B�	�Q�V�13*�	�u�q��.�B�I�b{�UH𠎯yq�ѣTDעq;�B�ɿ\���!�%�0�Q����m�`C�)� �=�p!��y/�A�w���T���� "O�Ը��߅�(�;.ݶ�$��C"O���B\�	T���w�sy>\��"O���4#�!lL�c�G���4q3"O�Y1�Tw�F����8�:]U"O8tB��Z��E�R�W�xajT"O�Ac𨕲 �z�I��3>��(:s"O6 ��ņ�A�&}�Ĉ�+�*i�%"OڀK�#L_��2�]�*<~M t"O����~�񐒡�xp!�5"O҈�TO_5���!t�2���d"O�����!I%@bgτu*��c"O&X�慁5ew�Ʌ��!�6�0Q"Ot|�"
��X��$������"O����A	'`�T9���	 C.�є"O$9� CE48�`Q���x�,���"O�y�U/I,��!��Dr�1�"ON� 5!�.p�x%!R>>���f"O�x���(+��Pa�ЧA{�]��"O4E�mN����Ô`�?P_�Xr�"O��jaI�N`ҧ�V�i{���f"O� c ,ƚ8Xx���>B��c"O�V�#,�Z\��4.<���*OtD�����%��lGJU�
�'��$�tOP�sv♨��T����{
�'`Z��q �g583��ѼQ��'c��9#
�]�` 2"��T����'ڴe[p'ƪg: ��+ý`NZp��'\����J޵�X`�`F9]!�
�'Ğ��"㊶yw&��w��ap,4	�')F50��-d���i��#�(E�'	�e;�xX�趣ϪbHy
�'�Ƭ�D����堣M�L�8p�'jj102G�)&�`���-�(��'��Rw�~(h�c%�醝P�'�qIc�S&?���8ck��	�.�'ׂ9�D��;>Y@���*�le�l(�'?l�b�e�7R��p�Pg��^Bغ�'���K)٠H�lۇ'F�Ex�
�'�V��0*o�����E=-9Tq[�'[�J�-�5+Bt�i\&�ج�
�'�AƬ��tJ~���G���
�'�jX�G�m�e��B>e�T0
�'mP�*� Q�S�q0�jյ/�l�R	�'�Lx����"-,��
5?r8���',$�J�#Z�@r�`(3�62��<��'J<͑�+�7\�P�" K�;�|�	�'SXM���\��h�C�H�i�'_�胹w<���	µ�$��'/���Um= ��cBl�$F����'�:�h�%��;2M��Ѻ ��'Q���"nҦ@/���d�E��
�'u��'�<	2�R$�R������':!�q��!h�ͫ�R�
�T4��'�R<�⯑�]n �h
�!�'���YS&�EK|�,�.rxpx
�'G�������Ijt��E�UdD�X�'��8�&#^9?�~`A�̏�P��a�'���ۧA^�o��e��O�2��m�'�,�'�U�Tɴ�#�&�l5��'N�
��� 3�&=�R�^�Ƭ�z	�'�RY�IJ$%���dd�*`��'Z�4��!�-Z�u��,��Z�X�'�D��t��	O+X4�R� ӨE�K>���� ���q��E������wSR�"Oz���>M��Y�DmM�gjn�S�"OX3`��/\�iV"�SH�+�"O�0,R32���a з\4��: ��x���=����`��p�.4�׏_9M4������W:�>-�Q'\�3�pp���+,,H��j=D���`@C����_�<X@F�<����))�nD��G�!W�
�?��	ɟ �'pay��Xh��A�w��>=�n4���y"��'~�@���aF9U�A���,��x�H=�i�"M� ���v��>E�!�䛖68&]3F��c��訕L�ax��'����I�aw.(3gW�@��'�ў�}ũJUҦ�;YH�K�� V̓EHr�<�|�����.�<����� k��afQL�<��_�ISqj! M+�^��<�!�#ړ6�@�'~	�r�C�)��¥
˗�~�h�'#0��K*��4���>�`Ca(<i�A �3�����i�J4D�2�F@|�P9��I�X�D����nKza����*����l�~�>�l@P�3��p<��`#��g먼�<!a#8�Ş.�ؽ	���hc�e3�ę���h�ȓS�(�8�D��P�d�*��Q�P��t�p�B�G�/�+TA�ya�0�ȓ;�]"�É�:��4x@��
5/����Q�ɖ^��Ur %�!T4��Q&Q�<�&B�I�)�xɹY�0��������d?�	i0`+E�ƕu&@�+�	�B�I�8V�p�@�$���F-�r+@c�,G{���k�1($�鐣�"��LI����?�@b+�S�OP�-x�)7rH4Q)5]��"O�]87����6�#�H)�L��i��$	lX��P���BnaA���6R�(@9D�X ffѳX-2bP��z��-��6D�ġ��F�,X"��g,ל\y�yB�F7D�`��c�,w,�$���9P���Ѧi?D��1�F:(�P�A�ŋn��y�en>D��k����:�"�an�b<D�\I�ʌ�|p�j%�37�M�Dd%�O.�ѾP#���B|ʑ��*�U�ȓuY��(0��i2��u휫��!Dz�i#ў��ǂc� |�FhE�g:pY�t�]4_#!��e:�cү!T����-�6
O��b���&hxl�6��Jb�À�'��Ds��Q"�-��HD��9��A��l�Ĵ��A� d�z5��	��D}��ȓj�X�[B�TY�H�����8R����{n[�f}��b���G����oN`��G<&��1��&~+��	m�'_T�	�e�Y����L�lIL�1�>���铸{����f������z���?A���ޗ؂��-�<ySjT�7��W!�dȗ%8(�R�e��s9����=d���F{�����a�='�^�C��ۻ4Q,�r�"O�T8t(�:2�|;�O��
�`b�"O��"3�ڮ`܉���&C
����"O	[��]f~e���-MUF�9�0O��dY�n �JPB�'�!�Ǆ��v�!�I�&��`�ͱ2�	:���6ў<��	��R�)���"x:����E�׆C������� �Ajb�5C�B�-�R:BG�..Q�Q�F
T�+��p?A�YAD�b��m�`z�oEfX��O����D�j��,�.�7�.Y��"O� ����8���	���
~,���"O�$�7�E�%w^�xsB$ut�8y1"O�͈�/�5KcF�2BH�6a`���"O���ĆF,|�y�� L+w+섓D"O.�cU�Pc��I2oH H���a"O$��'kA�S���(�-�2T("���h���)���\|i@��#��@+�!�M!�D�wL�i��%�"�q��T���	�4�ا���І5��|P��G�$���P���Xm!򤊲l�NQ���Ƥ/�����I�!�J,$V�A�)�G�"��4ØO2OVP
Gć�%���tG݁AF��+wR����|f� ��<�$�����*B�I!MGZ�ң,H��\��g�Z��B�I�A���Cd�bP��d(C�Z+�"?i�d/ڧcw���%�::"n����� �6e��C�H �ԕG[tt
���>um!�'�ў�'���߇w,"\�҇�$c(���/�I�!�d�(`�����C4(�c���\�!��P�V.G�#v�x �5*��T�ȓ���#�(H�D,~1�eA�9D_����g<����9G�&�c�H��N�Dc�k�g�<y��U�|%fLq��	Rd���M�<�ǔ	!��Hksa׋^�F�w@RŦ��`�h�/�4lɶ8��Q{����	� ]1Ob��ɰ%�����	�+������9lO�<p�f� 0�=yu�$�Cq�,�S�'K|hE���Id���xBOǺ�,�ȓ{ʎAю�5��8��A���4�Fx��'t�h:��S"Wz�s��M�E���JN>i
�uʸ찆[o]^\[�G��l�^C���<�TMY�I�ڐ�]3
��Li�om��(m�G����%̲�ِL�'ĩ��jA�џhF����<�VAB�(��i+��Ż��'�ў�O0���"�G! P$��&Y;�Dx��4�~b�/�S�O�B�kf���6�\����Ӱ5c\��	�'S�:e#  F=̔�#�@�P�*0�.�l؞�(�h)�}H�iL
p4�$��H=����:��>z�\ɉ@� �;��D��GM�	��C��i8�Ax�┻��B2��0��B�	�5<����Dו����"S0,��B�t*����Jo
̺栆�}G�B�{Sd��Eg�VI�F�D��l���9��&[F~i��C��2X�6��l�0B������3��$�p�f�/s��b�|qR�)�Ӧq �JQ.��h��,<\bC��������U����!��%b�ⴘ���>��� �H����?��@K��Y<F��l̓<������J=(!�l�D�K�?�a���691��ΑO�$�����4e莴��.�n죗#N-9�Ĩ,�9u=X	��a��]�A�/A6�x��� j���ȓz�~�I�ɜ8p�1)!�O k �P�ȓh~���bΚ�n��Őf	���P�'�0E�?Y��� l�[(y� �öZa�XX��"D��3��h�ndK"BM�`Mư�5�a��>5Tҧ�g�P�`����;����2�Q�0a�UFzr퉖J+"HLS❳���Q��q�R���$3�O.Y!р�+`����<@]�A���	T�OO�XuV
!�.P��7�i"Oz`˧�Щj��I�A�%αq"O��(2H���^u�G%�O����"O6mh5�&�. *bC�l�|�I"O�`���ߣD>����F�f���"O� ���ģȒ2�^u�  E�X���U"O��ôA�?z��G�6w���4"OP���D����:�o���-A�"O��@ v�&0��>U��:F"O
��W�U�΀[����+}�U�1"O�X�J�C���͐92	���"O� AW�ޜX����AO�M�
Dط"O~xj�G�/fX�	����,\��� "OY!� �.L��UH�n�+`ub!�"O��%�P�%��Bn�Y�1 �"O��! @�k�5z���R?��C�"O��"�	
B��׃-3x)z�"O� cw�׆d"����A��m"�Y�%"O�Aq���[ǰ�Q���,�.��q"O����^�Ζ� ��d�$�T"OzĠU��,�*�*5ذN�2�0�"O�(�%��W�~�[Ă�&f���!�"O����'�R��a73����"OH���ۙ(��,�ᛚ��+"O�Y�iˊz��)*�!Cp8up�"O�z�W�;�^��	~2�`B"O��Z����X^(bqb�??�P��Q"O:d8@���Q��M�>a�q"O8\0�$���q��H�}�q"�"OZ�Z�n�)���4M��D�n �"O������,���F�D�w��9J�"O�q���_e�"z�z�h��ݗ"r!򄅚p�+��Y�
ǦL�U�Ǳb�!��H�g�������&a��!D#��$y!��R�S���P��2b(R�yG!̵YQ!��Ko��P ����w��+!��U�HҲ���*�I�"<s4`�
!��)~00xb�C*I��d�v�Q�@!�«�lZ`��d��h�'�G@�!�[�D'�E�k�,�����f�!�Qi$����� .V�R#�,wl���mVj�x�"	rLt8�nl�h���+n\h�4E0|^$@IPN7D������5'
�q3���>6̩`�5D��p'�7-D����B(?0Cd�3D�4iL�r*�Yw$�=x���3E,D�Ȓ!N��!O�`���&��ћ0.D���′%#,,i�H��4�h���N,D�x�ҫ�n�Ta��� ��B�+FG0D�l9"�)ww�����<Q&	ҥn.D�0��
�N�<E��DA�+c�-D��0�E��M�@	$�]�-�$]��-D������t|F�a�ʚ�\b�A/�k/��P�'�w����M|�@`���c��@-jDԩEb�[�<y�Ux�*!�U��1-&�bBV̟`�w뒢X~���!$f�D���Y){��P��q���z��	-!�=�� �#
;�Zh���+f!��0=������$�8��d!U&$r!�$��k���G�A��xuja�!�$1x�f Ge_#]n�:��S x�!�d'o()6�Z�g$�QA�j�!�DU�+��ĺ��E@��Ѐ�>Y0!��Z�`�����Q�/<(�1u F�}�!�Ę�q`j��ϋ^"n�C-�=!�䈵;�UY��"&�s��]!�d��D����I�8�l��T���!�dYȠI��J��T�2�uiR��!��"68м�%L�ajPT���'�!��C!ycP�*�hHYR���ċ�(�!�D� YǴHxpJ��?�0+7	G~�!�� 
5�FG)�L���_�:`8�"Oج(BfD�Y2fp�� ��@D\�"O�����V���R�jZ2^���"Oά�VM?K�"X#�N��D�"O�mqp!��<�9é̝��@"�"OL��
VS{�in��E�"O��8�(��|�����X�d���'���w��7Ƅ�(E�� ��rt�ޝ�^�jsO�pY��C#p�ж�ޚvw�4�4�	/�d 3�΃�q����+�%~�쑁hW�c��s�"O(��E��� �ǜ�U �sp�'^�\
0�kv�KEP�"~�r��'^�b�b5��&-+�4�7�6��D�� n2aQ	ߓh�"Xy��SC�uZ0�O�x��'35�_Z���r�϶��'X�l��[�i��+��^��(�a)�H��X���>���ج���E ��V��!2��ݤ�^�C�@
<�x�y� Q	2�H�]b�Or�@�EJ�1Y��7	�-�����ם4�~����k��c>�b��
��� �sp�# �-�j����@�S�S��y�͘;SƬp �P��v1
#���?!5,�$-��p�W����)	���h���%?����%�	ђ�͓7� u�3O�Z���[��*����̷l�䨚�*�=m�I�1٢��*ߨ0X���<�S�_�6W����'x�~pa2ǥ#���@��n
��I�o���wǖA���BS	[#=�x��	*�U+4I�n�+�}K��J�7���|�Q�CӬl�s�*�@�V�w�'<n��0��oy���}ʗ�+,�^�9��J�BY�3J��}͌����� �dҧ���\�}H��0��0ܐ�R��rr�d�yڈ�d7��S�5񴵈gd�`�T`�����	�yCz}1f�E�l��zB��>�8�!g�˗g�0����\��p>ɔƒp�*�4C�T8������<K��آG��ȓ�Da!�ľb����3��ˠ�GzM\�o ��D���}�<���B�C�����E�y���!LH��D _-0f��j"��yr�Z+���)g�L,2�0��aː�y��_-@,Ƚ��(Z�G�P͓5���y��=1��xPA��!4q��K�
�y�g�*W�8'eYD���;�"��y�(M�u����dm�0@h��dC�y�c��%ؼ�����a��5f�5�y�ڷf�����;|��T!�B�/�ybG�p��\xU���k: �2tg�$�y��8P�@@�J�~��4��MR)�yB��s.�P���
A�z���D@�y��K�a/�8RU/ڒA�+��]��yrKژ.\2G�,2�����y"iK q�H��� �ݴ�mȶG!��K�1�h�ЧhT�I6ɃpI��9�'2��P	͕8�,�ʆN�S�!�V"G�<�A �bd�*��S؟iR��,F��Q�qH��:R�WɉD��i����̀�`Uq�IU��MSֈC!���5�L�Z�p�y���f�'�< �i �_��0��L��V�ӝc:m*&M��pT�"�����	1h�<���cR�hazr��r"��A1*�;�&������~2���U��qpT�Dmz�4�R�'�)��:���%�sip�S�|,PA���&��1��'u���G�?Q�H�'�+f4hZ6�X�zbR��Aϥ|8���惦d����fE>��I�O��k�� ��C�V�(�%ڊ}�~Z�&���M��}�@�3u)����O�(����*�=P�9�x�o��~�:"��V�{��٠Uh��M��q��9���D}�\_��i��X�;����o��|�#��4�nEjϑ�D9�ĺS�O?%�ҡ~�,�qf6LOr�J�I� y�E+�;��kG�O�ڟ~�^�(�ď�b���1��L�I�Uǜ��CV��4@�q E,Sgx%��ΆD��y�
�'��	E�C�KV�`လ�?��+RJP�Vn2���Dŉ�U�3)�<&��1%f�)��	�xI��A�0h2�/?;	��kf&��9�a"���J�B�OI�1f�K�=\����'��w�����[� O�1�cG.�j㞜J�g۫3l}{gM�n�H�vd,�m����2ɢ��[��D�]�02���e2*(��������N�Tʬ�
��v��OZ�$��r`$"Z �&���`�&'P�1M7�g�? ��5�U�I6�Q���&`��0�"O:4;#���V8DX����|�0�#F��0���O>�IT�,�3}��V�Rr�*G嘞{�6��R��y"_���1����h<d�Aㆿuc��`@��yi�}�j˷�F��ҏ�n�P�1����p=i��[:c��Wmy�(r�Ƃ��r�۵�ێ=���u�*D�Pr!��+���b�
�T���S�))ғLL&�(�%&�'AJ��T�۰&n8U�j��~o���ȓ%aܽ� �\�4��(G���lZ;Tֹ�b��s�h�O�p4%b7�Z,Q�@ܪ"O����|��g 3o@�	�^��S�͔� �{�^&䲙)TȄ#�-;�m��>A& %7�$�����C�V3���U��+��D[�������pR +A��BW�Ea��Ez��̀\�z0�'���35��e�&��3h�$=����΂<�y2��l�e�A�.3ϊ�扙��?i�&�6��d�d�Q��E��(�s�<6�P�u�ˉT?pA�:D� 1VKYchh(i ��z��H`���aF����	N��~�bΌ#\\[���$��X� �y�у�v1aB����	��N��?�q��@-���I=lO����EIt�mR1��-u൸�_����O�
qO�)��mQ�����M�� 7~rpI�#@��U�r���<Q(�op��Tc�(���$Hu~��F�!R�ACg�P<l.�� }�n���$�B�.Z1��AL�S�b!	�B��>I�E�w��EHu�p���k��>q�4MS�+�!;�^�QWR{&�O��*#�][�g?����	�����vc\�Aǉn�'u���%���������wb�O�
 c5��+=C��q
�L<��S��V�B��CM�5�����ғJ��4�'�h�tQ�
�x�(9����.w����
:���)�	�;�ĨG��Of�X��z�!�͘$+4k�"O���B���R�|)i���du	S�H�+dH�1Eoul�kѡ�3����bƄ�j�O��	�w,��4B���!kpg^�K�ͺ�:��I�m�'��a* 'Kf��j�������f,�z�e�-��b�"�DF�(��<B#�S��dhv�ڑ E��Ă 	���9ݨ/�"����4!*��mo>�� �El2K&a�Cc�k�O�<�@���'�!,O�	���Ț_Z�ŒyJ�熘�%����DL�(۲�0�3yf��y2�=F�O����2}ą��' � 4��b�6L����@��HH<1sD��KsδHF���2(X86@� ��̋a�V`��Q�+����L{д ƛ>i��'��ѐ�m׸6[Ԡ[P ^�f�I�����F^&]�����X� Q	�/����Cq,Q�6�����QS�x«�%.�-��@]s�=d��${���)X�#������x#э&�a[�m��'=^anκ�CF�?=v���-[�d�8�`�e�yy⃋�ii����#QVX�|�G^�`�`�Ao�A�јE�7]~�%BƎ
���J��ZΰA������!��y�Fk�y��� �N>Z���1- &��GO�X�(ʻ@m��D�LQ���MH�����A@T4yZX����\
܌h���:JI�O��nQ�U�������<sl��Ɔ�r����� 63 �;�G�Fm���v 8T�B�֝@!��Q.μj:�!�T(R5f�%�p0g� (R�n�&����D��Pp��@Ho��jկ;�^��es�!�:9�Ђ��@�<ӥj����D��P$�_�D"�a�҅z�	�Lp�(LO8��p�]�"j�q�f#�A�CB���3�¦�l:l� `d�<&2���>�N�=5X^ ��*: �qs4i��P�!�D�=��T��D�"*����Ξ�(���c1NN�O~<�b��*��Iڂ8��\-0� �� H�����:�f@�%h1|O̩a�ƥ]��!@�~�����L�Gh���'�Abo���g����?�ÊY�+�<!�F5&լ	R�n�@Ό��uǔ�I_�%@f��hN���e�ӯN*:Sq�Qb�#���"O���C��My�8
Ӄ�"e� (K:�X��TI"28b8�aF͂SC�>�	�`M`aA���ZK086�P9\_�B䉣ipL40#ҘH�*��Ρ7�$�V��;:��q�(a��� #�H">�M֤Nt��v�T8R4���JS����PB�~��Q��V�-��((à��Q�P�K�խ\ϐ�� 7���	&�j��6��,�!��I��~�`2�`R-F��
#�!4/V�;k�g����+�
��儻_U��s����yR�G`�����NL�D�`@�R/��B7r�8�鈈h��<B$i�5,��9���p�\�A.�<��$`���|���.D�� ,iJB
��y�> �$D�ByƸ�!+R'&�"a��I�MJ� �4<j�3�8�n�S��
�|�lȨ��EЎ����
]DI+2jN��Ɇaט`a�!�CD68r�@��t�4�:#l,�O�0���O�,0��ئ�*�pa��"O��+HF�� ��T��� ����"Oh�Cԣ٣O3�����p�(��5"Oΰ'�G�p�B�b�-;.ƾ���"Oj-a��A�>x��/��f�,q�W"O�,Gf%o��-qtndB,Z"O�p�S`W1 OD=�r�v5$�cC"O�PH��η�ѡ��n2b"O�!B��21Ud���W	~��b"OZ��S����A�Nf\�@w"O�����H��\�ьǫu� U"O���UD�#z6i�0P
65�V"O�1ar@ؙE�l=+$	8 �" q�"O����0q5����P6i�
�x�"O�h�g^?$��F�U�pT�"O�e�W/P+e��Q�.�� <p�PC"O��[bK$vt~`["�Ԫe��P�"O6a�A�[��2��0�],axnqX�"O��Y�<7�f��"ݮry"�t"OXY�ek�!A��-���0td�:�"Of�b� ���P6ƞ7�ε��"OB�2A^�n���֥�gv���"O���&�	�L��%�ń��Cj��"O��R$�@�];"m���'^I6�jt"O~�Z���4f͠�3�#A�*9���4"O:�1EPt�����Պ*�	��"O����(�?B3^p�"[=7�𙚕"O x��� ��q��X�f5A�"Ot<[�I�of���+�Z��hҴ"O�T��ᎋy%2��f�?�lʧ"O><�a:H �`�D̎9.�!�"O����I>X)��P��_	����"Oj��# /Rt��a#��(P���"O��Y��@j]H@��sRtt��"Oh�v�� � �W�d��;"O��9@Ǐ�r��ZՂV��&��"O����꓇V+��5 �<p�DZ "ORp�W`A&�Θ80`r�5z"O�Yð�� `i��
�*U"O�= C�G3~��`s�.��l�@Q"O�H�#�0���=Y���"O��Pn�t��P�C�;W��L��"O�4!�R����B)��F�H9�"O���c �:�v�Ȗ� �\�腑�"OVܫ �V�V�9sbg^�Nȶ"OL)���Xz��a'B�v��7"O��HS�(2�eS��?/���"O�8d�U��0�H��*�
�"O5sv	"WT���a�Z��g"Om3��0�0�fHƔ5�~�(�"O$Fb� Tr���8N�j5�"O��Q�JY�2{�<����;�4���"O���`� ��,	��'�1A*��I�"Oڌ �k	�V*�T��H�-s
���"Oj�K%a\TC���N��|�f"O
�Ѱd�XS�h�M�-+�F���"OT��Ba�)�@�Ӕ�X�]~e�b"O:%	�/��6���;�)�)1ΐ�C"O*���߿U<ԥ!ե�FB(���"ORP�Pa�~�yc1�ɩ`.���"O�-a!��.ڊ�� _�1�9V"O� ���D��
W���*Z�⤪�"O�i��`�U�<�) C0�lUrP"O����(N�E���D���*1"O m�oD�jn��7�Բn�6"Or��%�9|�v�r���Ja.�&"O�X��[�Z��d�D��o2� `"O%q��#oހ�Æ"�;��A"O!��͈Y� ��ЇA�1�4"OD(���B�iHlI���U�h=$\�p"OI"3�E�
�Da{qCOP�p"Oh�Q1/�2K��t`7��?�:i���'[(��E�"�����N�~ �x�`�; 6`�:�O �ᢉ.>�����P>��{��I�P&V �cǖ�q�ȸI�.މ�ҕ� %��[�d,B�"O�-�u ��/]8E�vJ@�*׎�1��'��Ȣe��k���b]�"~:�˙�*d���Opب��F?����/42�p�ߓB"�0�B�w�,���$��y��'_����M~����$H&:���s�a�2��b��b6|(�H]$(n�<�D�'l� ����i&4�	�`P�P�|���)Ȗb�21OΙ3��1]��	L�6� ˍ,F�V4�u
�8o1ў�(#DE"
5:�"S+ç[W\q�u"S�D(�� Z�j�P��5�Z���
$}��9O����d�ȹ�(�{���ȵ�'�"-���_����wX�"~��m��	N���(�<
$�Y�y"A�Tc�!�rn�`����C�?�F���	4E��E*���<	�!� 	��i���'�
�V��~A.��NU,�`a�sѐ�V�C��W���>I��?@�Z���W<�k ��4x1	��N׾*Zzɋy���/Vb=��GP~�O<`��4bS3mШ}��YI@\��������LxB���5��O0,�a�-Ԗ`���.��B(E	!CBB�VEI��Op��s��� �,{�<��#ȯ;�T�q�����;�!xa:�%��}�5+G
�@T$��T�:�jGB�<y�@ށGB|Aa��#\Or���-�a1��(a�bLx �'����aA��]y�6)M�Du��'��%[�� �yb@�-X��s���5�}����%�HO.y! ����h�b��������6 T�2<xpS�"O�1�t�A�+�
Q��6U)�8R�"O�L0���P����$�
�)썐�"O�M�)�&����F�
)�zI"O�I޵-bl���N�^���"O\  6GW��X��
p�>y�1"O.�s�E&b���Q��Q�8���""O�ћ�B��ͮ��M��xS"OD����vΖ�H��
�e�@	J�"O�5X�B̷VP"x�#��*fz@"O:Ժ5bZ��ބ2"D���sd"O�(["��tY8땡ըf�ҥ�r"O�i��#��pZ����_�t��G"O��+œ;����uX��C�4�!�䒿hl4d��G׮?D-E��uk!�dv*�p&)�T.���&�H(T�'/����(U�q�b�I�S���:��ġ�����po�I؟H*!�'�Dl[32��H���*AsIż�c#�I�	T��M�f�i�r�^.r�eh2�Wn�'��d�Vȁ tU��R �ن'��S)v�^Ժ���)I,���Ĉ��*����@UZa�M&G�az�lX����ڰcc2�	6�ˡ�~��:ڒ5[�A̰sY�I�(�i��c�4�S�X �x�H��#7pViy��Y1��x�'�jL@aGX�B�y�0"�*E��M�p�M!�ئ)�h���r| �����>'��Q;"�^��fX�i,`�jv�e�~c��Bᖸ*�B�D),m@�Y� �|�eҔW*�xP�bR7 U�OP�� h�h
�$��y��Q� ȭwe��.�4"R��OA3R�9v]���rʂ#$��t1�O�ʕ-�2F�.há�_�TZb���'۞-���(�P���	+Z�V$�qG]3{jH��)_"C=��	�9����CK�H�)����,A)�j��btc)Y�RL��d~ݣ�j�3<¢q[ )7D��PC��	/��C�D1b���	�J�=9|ࡠ��4�J�\�S�v�; �-��'�L��;x�"�������4���	�.b�!���;��QB� 2`yFl�R�L�U��mڲ�)@��b��TP��5]��'Őс� �j�qO�X�i�$`k̂b�#��8�����\���Q@K�*`�x8�d��|ZS�Dj�5��)�Z\�f��{y�@�*�T��	�JBNI�3ꌊ�2:C,J+\�O6
�l�.T���4�S;9�`XÅZ�!����B�,��B�I�]Q�Mj���e�� &C���u�]$��I�;'�!��Oh�t��T�v����*ڽ!7"Oؽ�N#*�1ɱ��^�(#�]y�%��.;�O�	���R�Rٮ�Cu�_;D��q�'�T����A~r�շ,�����fѦ��a�bID��y�c�0f2Y���֙�.�A����yR��F �O�|�N���K��y�Ks��XwDL|b4��P��yk�,O���i4��y�4�t���yRd�	}
rQ+�Q iў:����yr�Ht�� Q�85��`j���y#�
I�t(�CQZLn�ʗ���~��+��Ԇ�ɪqnnkWo�*l�(�ĝ��\���ĉ'��x �J�O^\�%���;l=����	-V��5"O�H��{D��A��
W-�6�d� g������7�H�X��MY�t�4 � d(1��V"Ol���@�bV<V��;t�eI�E��HP��@�Es�+�g?Q���0HΘH���_����țI�<����a���k�ʅ��ҟ�`���0�(����'�-9D�A1x\�Ь��y�
�ȄX��A�*�7m��eh>Q�4BT8�zeX�O��(�!��,Ah�\�o��;�蔄ʥ%��O�D�dU�_��d���i֛fŖ�H��$q�C��D=�!�ď9m��G�U�h�Li�W��E}�I��uBP�O��}�.��9� �H�,�p�!��ȓ*p���=Ij`y9E�S�����>H�ͫ��֖RUa{B,�-LؔI����4��H�����0>��ǒ�6��e)�w�ZU�S��qP�E1W犋L�a�ȓskh�x�=Yvĺ�(܋5��+���E�?Ic�D+2��'���;t�) RFΏ0���4�ǅ/����ēu����7S#�T��	AP��e��=~*|e"$z��O(t;���l����P�4��URT�S���x�W%A�܄�	�Oc���xQ�Q�/!��@��(��
�$��'���3si�g�.T��	�i��Q��U�Iid�a�0��M����ȋg�*y��+��_ê��e�0���l���q˟�.s@�i�+͵a��ٳ����x�!Uj�X�G��%y�A�":�	j��
4S�z�DTRP#�#Sf�p#E�'}�0�L�RI�u���R��@)l���V
OP�T���D����lޗ(Pl#�[�o�{�����u���x��I{9���J�I�"H< c͗¦�C�@mÖ���̄7U^8�F� `�%c+e�69Z0׊��Rp-;�<A[��S���T�(P��'�TE`��R�(�0�P5��t*�:�OPi��jѻ�D$��(��k\T��Թ@4�1P�,b�ז���9�+(�aʅ��#��x2�� �@��@
ҨA`.�����$e�$@1���$�$FB+���p&M��N��`*2}�4��d�$A�4�Q�BЕ[�$0b��'/���$)-�$�"�DNx: SA�84v����B'MT���p≅J��B�OF�uD E���Xٮ��B ڿ@�z�?�D�ʆP7xM�"� k���AH}�Y��ת:���Ӗ	�� "Yj@g"}�m�C@��ɨc�r����܈T���q솸k���2�nט~�Ιp��a�`�����)a�v�E��;A���2t�¡z{�eAa��2y@��G���Z��>���H�	J�T�Q���ŁAM�;�������|�	\�'�1Zs��)J��P��ǭQ[��(sr�"ŅѤC�

��ω;�8)�/Y�H��t
7�2mA輈3�3�O��adgx�t(#dJʉ� d�6��/�r)ac��83�(�h&h��'L�P��_�s����Z���ȓe>Z$i]�h3�p3TS�p�
pr��D� 0�%�FO�AP8m�4�h��$�. ��19�⚮T�t�!���?gR!�'�N�Q�ُq�Z1X
�WBM0R��`��¤��`�'L xP�`F�8	 ]I�@�F�$|OD�K&��j(T9��]�މ�"!ڎA\u�G�A<~ B�)� �0G/T�H~t��u��B�S���݃a" �1��_�?��"|���Ƃ�"F�.I�&,âKx�<���1�`ՠ����t�6��"�?,ՠ �0�Y8��'��>�I�.�����O+����#]*
C�	6��=���Ŏ0��!�'���牓xmV� ��#xS�zB�����b���hp�X:�BQ��p>yC�X�j�f�z���I�h���^�V�ӔO�|���"OD����
�hF@٨��(1"O�A '��)`?V����*F���"O:Y	�hA'}XV
��4DؠZ�"Oڕ���A�:d���D+
��`S3"OF�"�)�
U�n�0��0}ǄI�"O|H�3π�[��Y���)�Xd��"O�8��k�!���� �
BVzY[B"O��)kG�R��ѢQoݬak��2�*O��"CĔ�/��%�7���I�'ۚ� ��?h�Cf`�R�U��y���Y��I����2?c ����y�6�X0�fD?7ϲ-с�	�y��<lz��V��/+�`	�$�y�	6yc�łI�1� �QO��y�Ѱe8�$׫	�Ra����yB��!+&u`�Nx���������y2�#�n��(V#w>2�dIҾ�y2��+0�:D�_=c@}{U@_�y2�؝s�y��Xu��]�uG/�yb�17�R�X!�]`�LK��&�y��M�d��Hr�A�Y���!�"���y�H,@�5&H���q�g���y�dߎ|*�����NbF��c�+�y��]^�[��;D���	����y���
{����JW9x\��.���y�Q���`��:<,(�E*Q��yBM[�/��Hd@�%"�N��1+���y���t��|�ѨO�](		��yr :M�Uђ
��<�FH��y����N	���}���i�$��y�N���;��&��EG�ʉ�y򢄦;���2��-����
���ybB�1V$��8qH��[��y�
���5J��.֬Rv��yB�Ѣ`� �B8�H	�fN�y"E��m+|���?�d�c�y�N�J#x�cD
O35�h��RB���Ȏ�����x�T�FF��qUVАV>Oh���k�j^~ zbd	XlRY��>	�䈒����?I���A�|�,�3��['xV��5i�<����(�v9 �h\4B��2�C�#1�"mcv�'��A+��)ʧY0�x�͐&�1�E2U8���g����<�x�㑧K�,Q[֋G�n$8@�S�%��n%Q���C48��d����{R�T�k�`4�$C�;��)n��d�{�)�'QNM�թ]�<�%����l12�<��)�S���D"v�;Dmqn��Cj��I1k��#<E�Ԭ%w�����չ7�-���y�)�'2�vp[��E	qHr�1q�UH�+K>9)Oa�$	Q�4����)<-d��7��&�?A�
�8M���~��,O�|��ف^�He��eɽC��|��k�7 (���'J�'��>���N�/?W����@�z��T@���7��O�tiiŏ�2��8��S�D,0�'�ў"~���O�̀�@�2=t\r%F
��<��`����?^�s�C'e�([Æ�<{`>�l�k��ȟ�<��oQ������*�k	إ(A�sy�gk}B�&�g}RA%s����mҽTn��A指��~"O�T��h�<�r�"L�^�P�&�@����a��wA�	Zy
�'%B��h5�A�m  �*�2��EZ2d�V� �)O���π ���$�2t<]�UP	�"�B���9
Az�F1��рr SB�in�7\jU�q�>� ��n�Т��x���G��hI��BƎN�g,�����>�~�V�vup9k!7��S%�
X � �����@�S�aY�`��Ir�1?� �M�"}j��'[��XB٬Y�����yB���칩7C�P
�A�7b���y"��:,�`�0�ځ=T��+�C��y��ØB�Xt��d�~�C�Q��y�	X�q��(�@)F.q�%�b����yriՇhc�1��O�/VHV�`�ᐽ�y¦@�U�Mk����Nm�u�
�y����S�&$�t��D(�]Z`A��ybH��x��o�4�T@"���0�yRk�~s�3c�2�ɹ5 ���yb)�K��R�Ј��pᇤ�y���*�4E�'aV�U��BgNE9�y2%�e�F���,:����%�yҬ�9:�q�ŧ���8!�=�y���� ��	9C��u�U��\�y��� u�����A��p��w���y��<x-��(����S��K��yb�gl��"JV�p\d�:ZQ��C�	�<���Z�fX(pA
�:nD�B�I�as*�r�؋������# �B�I :5��G��of�Ӣ��C��B�	�~عb�J��M��F)txB�I74�J�_�� 3C�	z�pB�	�(�j��g�!*I��2p�X:y�|B�aS��̫V�Va���T�)�C�	!x�	{#��+=툴i���)l�LC䉤#���b��#x8p��T�E�8%dC�	�D�<��j�x�p���΢�@C�	�R.~m�mu��0�1kZ1�C�I�2%������-��HR��=y�C�	�jB�x8�$�&I<1{w�3~�C�I�%�|h�6�=ESR<с��#@�B�>��ȡĘ<P�N\�� �7|�B�I(5��1�A��TUpɂ
tlB�ɦG
��Qk��x�uA�!Dk,B�Ƀd8��A[8�*ЁV� �xw$B�(Y��('Ã�rb8�:���c3�C�I�:HP���3���.�:c�C��&/�z��&ɏRJ�-R@��x2|B�)u��գr
��D���`����7rB�I�:�бQ4Ufv2p�}{B�	�~�U9WD�g�VI����c�B�	,h�(HR�NՍFq"Ah#G!~�*B�	v
�D��]�t��ؠnCRn$B�I�=sRD��&ɪnƠ<�hZ�bC�{ζ��N��d������^C䉛{缈0��KT�+4�]>:�NC�I�9,<��� uH�ס�V�C�	��lB4HDJ�)
!�נ>` C��fЖ��d`͋/ƒa{��$(�C�	���!N�%|���!S)t��C�$\��4�t䟷o���r�O�(VC�I�r��1j�i�$V�B�Xv�΀s�B�	2Z�p�� 7���i�;[B�	=(��[@�T9t�:�5&U� B䉢}�C�L�8� �(s��w��C�I�_,|�Ϝ=��D��	B;�C�ɒ`�����C�����7͕0J4B�ɬ1
D�e��w��к?B�	�B�p���J�_`����� ">m�C�)� b8���r=̔`���p�Jp"OZ����oD�چ\|��X�"O��P��FB�@h��Q.vIzU r"O\9[B��}���+���>t[6"O@����:DL��5�,J � �"OX�8�(ް5��Z�'<��ؑ�"O��k4��qʄ�a�	B8T�3"O(\I�C�x$R=H�d�,!~P�@"OzU:ACM^l�Mx���L(1�a"O��YQ4<�rO�ubP�˃m\�<ig(��<�(1�b�)���0��Y�<��*Dui��Op����US�<a `K�z������\~�٪���i�<���
*%�HqF
>���y��	N�<y�.	%|t�J���6��4[5@�J�<9`m��N�h�cܭ������H�<	���w�xi�N�+J��U��N�<y��X�o`t<������я�K�<9��(�����n]�*78���V}�<q`�V�)RfA=]��-�&�T}�<�aF��"r(��G��	o
t�Js�<��ۅ$��\�هp5�DJWGn�<���8��q�O�(mq�A��h�<	%nV@@"�Q2��8;���	�k�d�<��#$0L|��ą7!��f�d�<'��w�ȐHaۊ8������v�<���T!u�.��a^� M��s/]r�<����3Q�n��"@GG�<�"��PT�<��#Ɔoڮ)�-_ Ӛ5��[D�<�f[�5�&�s��;:���D��~�<Qbk�N��|
��-k��NDR�<����=X����,�#[��(��Dx�<��'��eTa{EM��X�
�����}�<	d�ħ8�� �T���]��z�k�x�<Y � 4�½��!�>`x�cM�z�<�D�ئu���
 ��9J���ڲ���<YD�Y!Q��)�eh�]����D�<	'�]���s���=C+�А����XXtY���S���e��'��ȓQ�T�����{�i+s�GC�")�ȓ21���ɜF���nV�#�"Ʌȓ,:���O�jՂ���̈́ȓ@��`"gT4n}t�c�`N�M��ȓKr�0����%C͂�땢��G��ȓXYXSc�y馨���Dcݺ-��W�8qX�%ߟ`n���A�_�l�ȓg��VJѼ2�i�wN�N���ȓ�0	�� ���X��g[�Y�ȓ*|���W���^*���aj m��n��E�0G���QG	\:i����3����y����@�
:��Մ�RJQ���6~R�TP�Y;^æ$�ȓY>F�	�!נH"@�T$E�i9z)�ȓ��@�2 M9@��;4J4�,��J�,��x��`ߥcG��ȓmװ���D�b��a��#N���\��k'����I�'Ub䪗F\�hЅ�K(�@�%Ú��d�q&�:'ڙ��uO*��3��'�xت��S9�0ц�M^��B4̘�$	��S��r�.��m#P�E�6�`��9���ȓ$OY���"����#�>�f�ȓJ�~�#�)�4`�;����2ĄC�<1�l˃52�R��2?B�`2�	k�<� LA�!LO�>l��p��Y-�H"O:�$�S�z��ҷ�ʫ
+ء�"O$�9�	��Q�&�XHl�a�"OB��#+=�8H[A�߅ ę�3"OL�˕�±6�,Iu���?<�"O� B�w��sV�CWЬ:`"O"�H����(G/l@�"O<Ī�b�|s:U{"�q��	"Od�`Ce�1���#G���$eF0S�"O(MЀW���Uo��.rbA4�3D���C�̇SA U("��w�:��`?D�z� ;Y8r�H��H|h���9D�(a�Y�?TTD�M*T�`�#V�,D��pP�W*@���Ą�y�y�F+D��Y0a}p�[�@���y��+D��)0A�=5٦"��߶q��ի�d=D�@b^gl�C fݖ`��8id�<D���A�{�t͙�Eۅ$�p=�$>D��P#i
L���P*�8^�0�6D��K��]�}�u����xi�����6D���t�/���+�
�.C�B�	$*��*WLȐX�1!Z�/3�B�`Ǹ�zÄT@]�xZ���+5�B䉼W�>��ߤa�0Ks��jB��h(FTP5���#d���/\[_�C�I<b�v)��뇤e��a��Jr�B�*ZF�x`���֥��F)�C��6_��D�%�/��5��
D�v(�B�I�V��@t�W1�)ydE�;�C䉭P�"A$���q g��j�fC䉣Z`�	��+
�H��5���Q�I�bC�Ie�i0 ���܆�g�
�)�hC�	�U�@X�QAV5� -r%L'2�\C�I$)f �!��)�:t�%;lB�	�i��`���5~^��cB\j��C�I�`���cm��KvA�a�M�Q&^C䉊'�h�f�\�"�vU�֣ȉ"h�C��h���C��xZhyR�)�!91(C�	�v�C�*G�,�3�]�2C�	5�Z�Ѩā.뎄�*ݽ
��B�I�/2�����׵L;p�E���n�TB�I'yzD��c��ڔh�%5�rB�	]E��J���D���(Q��CHB�	�v�X�6�QI��r��Mev�C�ɇd�a� _ �|2��ɴ`{�C�$1bF�+^�Ԣ��cZjC��83���pei1�$�j��̭+{^C䉑���3H$Ha��%V�BC�	)&4�I���^�aYXq���9C{�C�ɋsxD����T�V�a���"��C�	6B�"�j�-� \D��|e{e"ON �E��do��"� :q�\hY�"O��p�撅�aa��)�^�!"O��q�:|O��G��e}���"OR��¢��k�풵���VW4��"O��1K'Q
�6o�B���)�"OX4I @^>0a @|�`Tc"O2�	r5 *��aF��!]���"O�X,����d�f�Cy��"O��@jߒt�ri!��H�c�cA"O��B�[�x��7�9Hލ@W"O�=�#�O��� fja�Ä'O�!�D��*�����m�K���M�	�!��C}B����% &>ȡ�0��E&!�� ��LǱF猕c%�B74����"O�<�m]�cݶpS���&����"O0���=�4��uV�|p���"Ony
�d��/>}�jK�]l\|��"O8�2�>k�����f~�E1T"O��r�,'9RFl[3�.*v�5��"OVB�h�?S�lz�bյ{��QX4"O|@���l����T*�`�bF"O���"K��u�h+�EϪhwD��"O�� �
 
  ��   F  �  �  �  m+  7  �B  TN  �X  �b  0o  "x  r~  ҄  #�  f�  ��  �  .�  p�  ��  ��  9�  {�  ��   �  C�  ��  ��  F�  R�  ��  � | � ' �&  - B3 �8  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h�=��K"�S�S)?\��Ǳy� �@u�A�B�A`���d�K~����,�R�ʢ<3a<O. �ӋQZ�im�8"j����'~ў|97G�|�X�P���
�F���:D����D��o�X�Q��/�4�q��<Q��)�'i
� �'���`-Б�X.F|�ȓ!{�jvf *�Й�"
���D�ɔfah�p_��1��>�,��4���=�ԟ|r�Z�� 0T�  n�$�'���y�U�M�(��pNX2x�ʭ�&$^4��>��O�􋢢�u���k��I8a��INx�;t
��]�p�H�6
�4d�S�D0�hO�	%�Y�rU*���2rHl�I��=А9�It<As��g��l����7
�^�I����<AC�O�"=���Ď�p�ؠ�ʏJ�
�ȳGW�!����� `��(@�������
m���#�O�Q�L�=f��ij��K2Q�W(�y��}n H��
+�Y2O����$N8�(O�>�Ӵ�'>8
�e�9� =���?OL#=ї��%["�S�o�b� ���lB���=�dQuMą�#�H\%��!�/�{�<p���0Ll�bE��m"PP��@}�<�w = ����Q�	�n-1t��v�<���H�S#D�HC��rc*���Fr�<�6jöaU�m"�������n�<����w�X4 ����/������E�<��+,�:� \ ��p�ŌH�<�feQd�	��C�W���
o�N�'�Q?��'�R�U:B�i��]���芰�#D��I��[�U�2���ZG�4�� b��qK���sӆH�����4������H��'-��� &�
6 M�n�l�3NA����uO�	_x�li�oN�6,�4�I�\(�y��(�Ob6M�<� �Q�� ^T*��;c�P����"OV���&*�z{U���V9q�"O> :dj6:��2P�X7iF< "O�q���j�H`B��T2���'4�')2d�dMF?^��Y�F)۾1R�/?�83d)�u���(�'�T��t�Q�>D�@��M��B�86	]LddI�;D�Ċ�%P�iQ4��f�&�` �b6D� b(B?BI�a�Ê5Y6�4D���@�E�d�|@w��M���%6D���"�@�?Y���AO�0J:�ղ���hO?�D0:g����EQ8m8��N!�D�	6�Z!�X�\�f5aD�Sn�!��=���EG�%�Fv	?l�{�k�q��S+��	U�^8]�p���[" B�	u�T@���Ñ��G�/d��˓��k��)*K�q��"(D$�ظ�j�nP�B�I2u	Fݨ�+��M���L	"<�%+K���O�ϸ'$�¦V3 ��B�-ʔ�L�"ߓ��'��$��(
�|�^L� ^�%zTa�O���dӒN�^d��K�<#�H��@H86!��E�
��_(1ʔ�� >����"O`DH`*�yԌ��&G�H�8R�O�=E�t�==5Zd��������G�y�B��mrhR�Żf�܈f����O^�҄E�=�e/].Po�e��˒E�'0�?a2㍖�`�r�%�YG����3D�T��%O<s�r�6nX���)0��1D�H�GG�b�����Ĭ jyP%O����� ��ĳ(�N�Pu@�;<H8B䉲7d�p8g晢n�8'�>@�(B�	�x���+L@� �Ѵgd$�>I���� c�$Q��E
��5z��ST�!�䚟ck���&D�.%{x�b(E�I�!���j<䠈��P�@h��r�fI�(�ў���I(!�l(�4�k߾tyţQ��<	˓BJ��COZ�<b�Ű�,}7�T��Im?��Ï%<��	�"hV���kMŞ����i>\�b\��Z�H��J5& �ȓ��Ħ<���ԏ�4"�ư�r'��m~�!�Cк�y���5u[�C�%w�$�W���y��E����`�/!=�9�3n�2�yIC
{�^Q����o[@q�w�A�����6Oʈ�!'�������Ad��j�"OB�9qR�Y����E/�^�FŃ�"O܌���A�B����?�b%h0"O�j3i[07BҁZ#쇦
�!x�"O��BdF�if��mڭ�P�B�"O��YӋ҆'�f���,
��p�W�'�f��'�x�C��ͻ
BH��5JU�S�a[	�'��sdي_'l��4��SC�5Ј�Bi���ɉ�P|�Xgc�T| ��C��6!�Z'|������&e�ͩ�o���F{���'_�4��AڍL�<yo��z�����'�|� $��ޤ	�*ҴP��'���D#<�d5��kH�H�0���'�h�U�A+	6]EbP�Pya�'Ж!3��\�'U�ȳ�Υ_��t��'����G�o�.�cI�A@�E*�'�
�W��1��!�=�.�(�'oR1�N��tn��g�^�8�:ES���4�',k�%��)O�m�USv��!�L���B>�$Ȓ�K;��(�3M�].|�����<�����hE�8���W1��=�5��e�<� �mC'o�� ���A!k�QҨ�u�d�U}�@�v�<��/���A����<|�r�\�K"@�	�'�v�3�oڌdq��j�FtF �
�7q�c� f��)ZN�:��K�p�)�B4D�p�W� 38�E+�v>��#�0D�lQqHC�nh	�6!�
ztP�h;<O�"<1iJ�;ͺ�i��y�`�f@t�w�<�Ԏ��S�0`��=B��ж-�O��	���)��L3z��+&�U4(�B�*�,�����!k��b��Q�A�>G{��9Ox��D��>tB�p�B�o[�5���	���?ud���Le�x;0�_=��vKܭ�M����hOQ>�XoX�$/VYQ�烀U���,3,O�<��4�X��j��lr�ds!�x�<��ʌQ�	�RG��5i��`GuX��q�]�s��R!,~�+��6]���`-D��I2���P���C�EՄH�)��0|����<Yr��@0� l�J�<��׎g:*���f-$@�x�G-�B�<1a΅px�e�D�%p�����U~�<��D�ؖ����_3�i0 �v�<IF�ƲDK��j���/NM0ir�'<Q?�І*͡?�B��!�������8D��S�f��$�&�NP#%<�§7ړ�0|�b*�1B�8��D���st�mx�<�'B��r�`Z��za9#ͼh�]2���䒤��S����P"}8�c٤3�
�jsIQ��0?ѣ�ǡX�&�"\&��**����Ň�yBG�o*eC5�ދ��!�B����O����#ҧpj�YR�-W�URtdOE:M�H���=��\h��]�`{�8�`�@�b��e�ȓ%ꐹ	��?S��Q���la�ȓ��P�u ވE����Є
Ga��
�B����×D�>�!^�輄ȓb��0��	Ƌp>�<�p��g�<�ȓb�ta3D[xJ�q`	�!&Ʌ�W�����-��+�eG+R��ȓN�(��b�K*P�����*ʥ[bȅȓ6�x��hӱa���B�
%S~�1��z^�l'�R!p�r��G:�x��ȓ��x��O��|����'L�~gx�ȓ\j��ь
 !�P0F�?�2��ȓc~�x���D�k� ���)��H��d�U.�=/��ၖ�mcxe�ȓS)*hu�ȅ���;��ӫ3��E�ȓ&���QV%��lh���'�5�4T��@�ABD�RFϚ����R�A��ȓ�8��j|T܈���3�ȓo���v�U`$-���7�Z�ȓT�Hext�:/t @���-����U/��qR�ƚU,��BV�[��X��`��)�b�
�if���&�	�4��L�u	��/U��kv�R�vl��B���`d�T)/YV�BF'O�-!�ȓ#V�C"M<%��izA�-UҢ݄� ( 	+KF."�Q�3H�+Z^���hK�H"����QFPb��$6H��ȓS%��Ґ ޽Q�Y�u�C\�ȓ0J�m�)�>�3�(Z�n��ȓg ���4(ü�v�å��shم�VB��v���
��u{���$^5��ȓPP�0G��Zx����#�d�ȓ/(J� ���(���=��ȓTLЅa�D��2IuB��Ko���S�? 8�ArdB�@���)#Jb왐"O,���
�U+f,�H �kw�X�R"O���
\�:�.�*���{s�ԁ�"O���ӀXx������BhA�"O�8�f�G�:$M�6�O4x2��4�'i"�'���'���'���'�R�'ٸ}K���|׈$�%	�'D�Q�'~��'^b�'"��'���'��'ntAx�*m\�Ѓ���3�6I��'���'�b�'���'���'Er�'�r�XA�Ǫ#Y�d�E�/n�q�L�O>�$�O(��OD���Of���O"���O��S�MvFEdm(���D��O��D�O����O�d�O����O��d�O�l�u&�$��!�&X�z醵���O���O��d�O����OX�d�O����O��9š�45�`A!t�۵I(��6��O4���O���O����O��$�O����O"8�%�;x��劃�ހv�:,����O����O(�D�O���Ov���O����O�4�C�7�:�`,�J\�Xvo�O���O��$�Ov���O(���O����O(P�'Y�?�<ES�DJ�XJ&��Q��O��D�OV�d�O���O��O���OH�9�����|�aee��#��i�V��O��$�O&���O���O��4�?����?���P1+�jXs���Bߜ��f���?���?���?��?	���?i��?�����Y�-@2!d�aZ���?a��?9��?���?y�e���'���S4 Y�����\�n�t+���<˓�?�+O1��	��M��/�5�U9(Tj����(T�xT�'Z6-/�i>�	�M��+'5(�ƛ��H��������',v�:�����dF�P���q�Ť����8�^�jި`�Aav�ί���<i����5�'������i�;�k� 2v�� �i$p@Éy��	^ݦ��PGT4"g�I��:hV��X0ݴ&E�8O��S�'7Oʙ:�#��<�L���@AN��n�Z�*��<1k�,���I��\*�hO��O�ݑ��;�^��
�����0OR˓��M2������'و���* ����-@������	K}�bӦ8n�<q�O�\*�z�
tS*�p �����LU,��y�-�S	)�I��џhX�eF��hQs�Mŗ���d��FyR]��)��<�@�� +�����=�^���W�<�ѷi�ba��OJ�n�L��|
#��;�bh�7|�H���BD�<�v�i �6��OV}���¤:\��1ZP�!���J$ޭS�a�@FLJR
Y�ZzT�V��z���4R��%?E��I9\����6 �]Չ9?�V�i�ڴ�y��O��O�V�i���-�u��
Q��`!��������ݴ�y����O@��N�LI��(�K<m���3���������D�l-��h��ndX�M���O�d9�T�eB�ͫ�ŕ4j�tQ��OB˓��,���)r@t��0��rF��q4��-�%��t�����IC�i>�I3�MK��i"A�<`�DDb6)my���4��:�L�k#"�͓�As��"5"��:E�?���x�I@Ycp�`T�Q�J��a�j�>~<LS�'��T������hM�Rc����C��=!_4�ȑ��J覭@Ae=?���iW�R���$���)a⦑8-�j!��F�<��ODlm���Ms���P���č�<A��d$`�0X���24K�}#�,�� T.*���%+E��hO�I�<���X}��J��L�u$P�z=����ck�faQ���'��t�Of.�K���Ļ��#F��O��'�D6͔Ŧ���ħ�
�"�!C|�1pQ��)49���n)R%z#gI(bxU�'��DO�Vȴ�0�|��O�Jޭ��#|-�u)�4��K�4N��:L�B��H(ۍWP�XbUmU��?)��?Ǜ&��`}�fz��ɢU'�HQ��`(F�Ч�)ش��D�� �f~�@�!��丷A%��A�$�OD�r:�s��4Wǆ�ByR�'c�|��g0U[긢DCE�U���q�`Ӛ�"���Oj�d�O��?}�����ᚹm"�� �^�j�����I�6Q���d��'�b>����ضOj�扮��M�4�	`��ԙ���1p�V�I�I#�$�V�ǜj�9&�(�'�剦da�Ժ�Y�E�\�pBG�'"���P�%[��͟6�i�BG�x��!�I B���aƀyy�Oz��'�6BѦ=�J<i ��_`���D�x�����W~���;�b��BF��wE�OFu
!�͍w�� L�}�J�<��`���*�y����vQ\�����7��8
��@!$��^����OR��ڦ��?�;�
ك�g�
!����G�Q��,�z�&�b�x0n�g��I�T�(?���߃����a	�=���z��2#�!aP��I�<��K>y(O��?����,o�ms F�4nFF��Uas~��f��9�G�O����O�?��`�4#��X KˣM��s�꒳��d���=�ܴy/���O�l�����B=2������`��S�h}b��QW�4'ϗ�y:�h"���7�Z	�U���F���8�"�(��ꡈ�K#I2s�9*��!gi��� t��#=����B D�n�+#��K��s��'��T��n��<������'�4PQ$�@�#K�8�`.�"-pE���H�<��ʓ��8�r��-��\[X�`���@�0�������3	�"E�w�.�j�Pu$)6�`�3p�P�w�2aA�/�	c+: � ��%=��������(��#7̰)r� ����
�ĥ�	�q�u�4�2�Hq a�_�o���Ƨ�vSZ��,�+�="�Ƅ5bb�T� �ie�U�5�J/b,��!�<m԰�Q�k�>y��?9N>q���?aT��?�R�1m)Jir�e�RN��[>����4�?����?���?��0g<51��?y��o)�Xk@��8�.���@+>:ic��il�|��'mB	�Y��J<i7�T�<ٖa
��Jjs耨 ����I��X�Iݟ�C��i�4�'wr�O��T���ӏi��HW셸�L�0�7��O��d�
Z'H���T?
c���"��D�p X�K̩cg�sӎ���O������OL�D�<����?9�����}�L �^(@��[�V�%�Iן$�vV>t�b�b?��p%�.��J�(N�wΈ݁v�j�s�B�O~�d�O(��@���O�˧ �:Q8b�S<����V�Pݖ�!Ծi����㘧����#P������~Q	�E8Zo�Ɵ�I�閆WyX>��	S?�r���5+�q��	KPq �[U�1Oޡ{�D�n����Iğ0�������$Z�!�2	�R�D�+�MK��rw������?Y�\?�	r�ɪ��(Y�(G0@�9e�a؅��OΜ㲋�l����|����ԕ'+k�r��`;A�]�L��u�;�j�3O<����?�O>���?��D�9ʹ���D`:\�y�jʃI!x!�<���?i����d�D) ��>].��9��>h_``(�.Rt�6m�OJ���O��OH���O��R-���3W��FhlY�C��&��aA'�>����?�����D�?@�~ʧ�?��e�.��x5�X$s���+�A����'��'/��'� Ls�d�g��
%�]*S�nm �		�K���'�rZ�� �Gs�4�'Ar�O�"���,�t�pc�U���镠+���O�����](h��Z�*�s�	sP�M��ԏ��QmEy"ӓ��'��'F�t[��X�,+�Hp\3d3��2�ɇ:�06M�Ol��
�
m0�b?���b��
���ũ��.��i5 �T`H0#�O���O���˓�?��Ӟ��6�B����!-���R3�i��2���֟����Ρ��d��^7�
yZ ��M����?a���;*O0��OV�䬟T��(u7� �pȻ..* )�+>�Ic=�&�\��ݟX�	� ��ԡ_�,o��Y��e�����4�?I$�֑��D�Ot��O��Ok��	?�-0�$��W*��Xaa�*"��ɡ5�x�&������p��Jyr�� ��(�P�,CS'ΈbR�T�0R�`�IܟL��@�	ܟH����=����?��gԊ#�B��7�VS��Ɵ0��ߟ�'19tҟ��Ф�j�6�s�.G
�R�$�i��'OB�|�'Nτ�L��D�S*�k�	)l86���ӪT��I����'���]>���(Mj�����mr\s"��&.�ݫش�?�H>���?��!S��'���#�B*b�����;��Q�4�?�����L�/z��'�?Q���FjK)9���%$5�(�b��'I�'�D�Y��T?�S�^�d���F� ��djwӈ�;z��0�i�v�'�?�'~�I6[+��U@�[0ШKЪ�4Pn(6M�O��K1�dE�d�'2��Z>7M�8��[��2XZ�!pD�cq���^oa7��O
���Ob�)�b�i>�X�*�bS�TS\�:�K2ĸ6��,4���O~���O���|Γ�?Y2&_�Q��i�s C�%��f�nE���'t��'H���V�(�4����OrI�$�R�Z�j|JT�N8���pŋЦ��	͟��Ɇ��������X�I�bh�<CP���@w"�;}�0�sٴ�?���f뉧��'��^�8�ѨN`d���6}��C����M-O���<	��?!�����S��� v-��jr��SZ
.��f#�H�	��X��Ο��'�rݟ@%Q�hV(L7�I!ˀ8t	���i�R[�h�IΟ �'"��R~�IC%��Y
V+�:���z9�U���?Q���d��r��fÐ�*�άp�o�.���aŋ�ē�?(O���9mt˧�?	W%�^� ��U,���������O��*��m'�8� �^B�V�Ȃ]��8۰Kw�d�D�<9��'P&�+�����O����8`��X�>8�Br�Y�[iz0�a�x��'��I!g9�"<�;O@�٣��1Wq`Hr¯��(�t��'B�$m���'��	�?���uG��<oI$K@ƛAԾ��wȞ�M������D���2y BL �+��$ȕ45�fmŻiz�M3��z�J�d�OH�����X'���b*����O�8�D���n�s�F��4�?����?����d�|Γ�?iG\<a�t���&�SC�y"#����'�"�'3X ��5�4����O��k�͋=Y�,	�LQ7"(�E�Պ���ӟ �'�P�g~��'���Ew����UT8F,�-S2���k%$7��O�����u�i>!����'��H��$
+5����\I�r-�ף�&�Mc��a�y����4��$�<���\�$a��
��f�z=���O9��h]���+O����O����I��H�R�B6b=�$9C�äo4Z%���*X��!�3?Y���?����(:�X�'E�u0$�� �R@�H̘X�ڜ�'(��'`�V���IڟT�b��П��p��z��LW�KP�P�Ǚ�����Oh��Ov�]"6p
F��t��C
PK">T`�7P�G��6M�O����<	���?����?�K?� �	a`/�/.
�Z�j�9(x,�C��i\BQ�D�	�"�4�O�2�'H�\c%��c�T��r�I�lJc&��0N<q��?)
��|�<�O�T]a!��{���+��d�3�Ot���&6'����O����O�I�<��T�xU+�!�+��#��4j_jXnZ���	2N���c�4�)��'y7ze1�_�Hz�0#ŦY��b7M�(D�h�o�͟�����������|�1I���hs#�z���kd$ͬ̎mZ���I����Iџ��d��'F�Gphͺt�>s�5kÍ(6-�O����O@�C�\B�i>��	����%���/w� `Dlp���r�я�M����?���&�0E��Y?�O�OT�ѷ���l]s�Cʘy��lQ�i�b̚x�	����>�ɾMo�,���L�)?,�VďG��8��OF�!ŗ]����$�I��l�'���H?hFTY�B�}V6��w�QZ�O����O4��<����?Q�.�&�ڹ$͘�1l,��	��x-
���$�O ���OR˓#�Rhxv8�F� H�/p`�%��l�����P�8�	şl��]y��'�dH*_Y�P:��faف~�t�00`۪��꓊?����?�,OVT��MON⓽!�F��5�
1�]����9�v�a�4�?����d�On�I�"����|�ŋ�
���-�+!��1c���K���'�I��P��M���'���5�B�?��%P�U"9�� ��&���?����r��HMO�S������� b�ɵ(b�)cuK�;�MK��?QR��?3����'���'����O�rc��H�
�i&�Ȼf�*�۔�F$$�Zꓹ?i!P(�?���4�p�O�	P�#2�<���Y�2�i�۴O�
X:ѳi��'���O����'���':����$O��P�d*[<Hxn��&im����&��ON�O�<�i�O���&U8� �nĤ��&b�զ����4���Y̨�4�?i��?����?��! �d��'6�N�;��ے>���l�ٟ�'Jj�#�����O�d�O�d	���$�yr�h��A� ��!͇Ǧ1��e0\�Jش�?A���?q��U	��M?�4��=�N�����n������TX}B<�y�]����˟L��wy2o�Og��зJ;>4����\�.�� ��	�>�)O����<����?���s>�i���T�EKL8�򅘍?6 *bE��<��?1��?�����dO�b�ZU�'c�2�Bf��)2`����k�NhnZDy�'o�	ğ��	ԟ�yvm{�\��IΈ`06X�͞����0&O������O$�d�Od�D�O�X�MȦ��IΟ�F��3*�lq��ҀaB�l	��:�M����?�����O����8�@�d��КWǞ0��}���V��:2�lc���d�OZ���O�<QS�S����I韐���?��G�]1\T��Щ��S���d邳�M#������Od�Ju;�:�d�<��e�/��6l�B��\��c������OR@0�i\ߦ��I��<�I�?m��̟<Hu��'/�*�C���!�*��͒���$�Opc  �O|���O�ʧ���Wɒ�i��I�jt��A˯"��6�J�[��lZ�T�I�@�S�?����p�I�$�T<�3���ТƩ)a�=�޴F$N�������|�H~��+\��'��;�v5��(K
"Da�i���'���;�x7�O�D�O����O��
�xѨ|C�ſA�p�{W+�Y��v�'���2mR��)2���?y�x�*��H4m�4h��+�nE#B�i�b�K1>�zO,���O<�Ok��$B��V��Ֆ�2e�
Jk���O��IUy��'a"�'T�I�Yu�xy�D��3�t��@%�3L�a��)�ē�?Y����?Q�m��[!a�|9��M�`%N�B�[3�?�(O����Od�ģ<iFߢUG�	�Ԡ���w/5���K&��ߟ8�IH��ߟ<��k��� j�x�X�/�1]���ʘ�4:~�2�O����O8�D�<A'IV��O.�m�#��[�4]�Mҿ �x�CQs���8���O�D�.v�$>}b& $12��e�L6��mܷc����'��]�8�����ħ�?�'@b$�JnH�G�N����B4+�鱠�xr�'i�� X(��|����H��K(l�؁�&�� x( Źi��ɴ!�4�4{�������S���;iZ$�F�:S�F,a@V=Ar�6�'��bK��y2�|����ۻ?���U �_R|�Ғ��s�@���MS��?����C�x��'���Q��뾴Y�B�u���m}Ӷ��5C�O\�O>]�I�cTZH��΃-j���	��؀�ݴ�?����?A��,��'���'H�Dؕ|c:�kp��,\��	�E,�;Y���|�*�N�8�|�d�O
��V �#�S�R�����b��6�' ,����0�$�O���)����ʷ�P��ʴ�F�k�e�C]�����m�@�'�2�'P]��@���&]�0�LN f�z@��at� ��M<����?�K>���?A���N@���%��e+����P;>������On�D�OjʓKݠ,�T=�`�hH;h�(H��)�(u��^�x�	ڟX$�|�Iڟ�Rbn����
4H�m�5���C}
"���D�OH���O�˓`2������do��	pa�gRsiTE�C�Dh�7��OВO����O\�c��Oj�'X��ʒ'���tc/F�@�y�4�?�����C��U'>��I�?Y��]�ق�L�Nb�@k�a���ē�?��2:μ�����S���ʏ.("�P�A�C��«�M�)O�,a�bEئ�
��R�$ퟦ��'��:��R�8I6���\�5��L��4�?���$m6�����S�g�? ���&BT����ǎ�qS��3�i4^P�t�{��D�O����~x'��S:�>����<)���"�=$�B۴������?���Wh�>m�I:@�VQp���[h(-r�'�� ڴ�?���?�C
>tC���4�>1��ـv���q�fV�\� ��&���}�'�����$�O���ـy��0���<���+�N,Q_2�o����HZ#���|R��$� 	�f�*"͋
��k0����6�'J��"��'^��ԟ��ɟ|�	ϟx���ώT�B�8���1�"Q��.��p����ʟ���şL�IN�şH�I>v,�a�K
AV����((�<�J��]�i@���?���?�)Ö��k��|�wm 	1D��av
ej%dG�n}��'0R�'��On ��W?��G��zN��M��^�h�ȹ>���?a���?��;�T����?a��<�¼"9?[Ƚr���ȡ�žib�|��'c�k�!b����H<�$��V����d&������I����'���1�:�	�O��)�5{%$�Q�!�c;�XrF�<j
*l'���Iß|E(�S��B��ѓ�̥n�����M�*O�ܫ��K�����������LY�'U�){���0i�,�Z� ��N���ݴ�?�c"��Dx��DH�-2���.�2�@�PA�M��eD��?���?����*(O\�'_d-3ST�D�+����-9��i�&��fg�����8��N�u� U`���3h�pڰ L�:a��m�����ߟT�������|����?QT�%v���#&� �%�������}z�O���rk=�D�O����Oڥ�t'΍*Ӱ�3VHԡx��#+�ۦ��	eF��'��ꧪ?M>�s��ry�E�!
$Zhpu{P-�32���6-�tD$?)��?A��?��tE4e�d���x���Hy�`�����OV���O �OT���O���猎�=�dD��J�TQ�M�k*�U"��X��ğ���Ly�"+N�V��6^����L�T��,�]裬O8�$�OF�d?�� j7��'eJJ����:���Y�Ê����'Q��'u��'��*_yr�'�b��  ����f��6l�Ыc��6M�O��Op�d�Oj�`���'�5���:t�"I���R�AX޴�?y���Y��Jx%>!�	�?u��	ہ~ri
�%e�0\C���ē�?���I���Fx����Ag�Z�:I�y����bX:u�i��	q�|��ߴA'��ݟ����DC�Ams�L
3s�ma�[�!�&�'��k��O���E�D��aUzmB���D�q�K�����L�M����?I���
���?����?E��F�� ���o�����˴1�����%b�'�-�~*I~��M�`�#�A':��Z7�T&E��%�нiR��'�b"G��7m�O�D�O���O�_4�V� h�/xf��Ibתכ��|"*��yʟ��$�O��3)��k��Z�/���"�	X�nZ��LHHֿ�M3��?���?y�S?��7q�PPT�g�ɨ,>)MJ<o����gy�@��ɟ��I���I䟘�	�r��K���=o���/�pwz��&�O�M���?���?i�X?=�' R�3JK���ւ��<��8dc�)N�q�'$��'���'sRR>99UD=�MSrD��G��2L�s�M�v��ƛ��'Hb�'���'�����iBa>"�C�	O��U9�D
' �����$����O���O$���O2�sE������I柴�į�	|p��C�I>Tp(�1�M;���?a������O���4��˓y0D c��V�R ���Ǿ9:|P��i�B�'�"�'��3G`o����O��D���ya�Ǳj8�w&U9*+浸��ʦ���ry"�'�4
�S�����ܴ�P
A�#Z���B�	
D�mZԟ8�� �����ƟP�'S�D�'Zc &t" A1:���[F�	���4�?!��DX\x��}�S�'[U�1�Ù�^��$�1bT�:��IoZ�L�6�۴�?��?���ab����cB7H(K�R$M�DxcE�_�pɀ7M�x����3�	⟤ �jѹb)6���$V����aA���M����?�J���+ONʧ�?a�'�(�#�&gO��Q��)<z�c��>�	�E
M�N|���?���Eu�9�UKF�V<x�7�P1}��+�i��?|�7m�O��$�O���t���O� ���R��ÇK�<r�����ia2�-�y�^��������	�����vo̝*U�[n�0r,��a9�h����M����?a���?ybZ?��'z��Ŭ[J��ڄɔn�	���K~�:�'���'&2�'�S۟@�#.�%�M[��m5� [��v
��C����'Nr�'�b�'����4Т�b>]�Bϸj������2A�0�e�^��M��?����?�V?Mi$���M#��?YW-�~Q��:�ɓ�s�􉨡(�$l���'�b�'��	矰�pok>!�O���"��>&�U��hҜ)sLl�׿iNR�'�"�'	r0��+j���D�O������HI���4o5�0'N:C�|��� �����	Cy��'��Z��4����D�]"���)Y��J���M����?�!�+$ݛ��'0�'���O�blWs��|B �0b�N�T*��m,H��?���!����L<!eaL 0�h	B��	.|Ds�SȦU*&Hڽ�M����?����z�'�?���?�`��;���� �/��者O�!�&�W�F���'�i>e'?)�Ɍ{����
�7L�9bS�Ɛ=/��B�4�?����?yqD:���|r��~����Z�����%={QaQ˝�&�2"<�'����'��'?j� �u��C$0�H��S7j*}�ǻi�Bjɹ!��s��ɟ�Iu�dϮdxʑ�Y3�U�C�zD�'<�'
��'k��'����"8N=Ҧ�	3d��K�iE�P�\�Q�������I@�����Ń�-%8��E�)_mX�m6FN�JK�D���̾W��T��o��J�h후�?�	 ����źI��K�B����0D�ܩ��2H�AB bN)�>��-�j����N7#��q%��al� ���#r�$�2��L��a[�iQ�9��l;#��t�"�iT���.�:�nȭN |�Ԯ�x��Ro\��^����� @�� (�n])jD�p��A�P�H!���!{F��8��VIS$���
�5��D�V��1Y�Jn��!� �	9w9r��?;��y�u�I��c�E�2�J���O��Y#l�;l�*�%�x�6�GӺ��jČ��I�^ubL���(h�<E3�j�	y��p��Ջ���,7��0"MB~�X5q^w�p%36I�~��۳���:��8A��2gFj�߮q��n���E���O�p����-�m��.A�$@�͹O �j�Ð^yL��T�LH��'y�#=QĤ�3P��Y"�˾1)�U R��#Gl�	ϟt�	�c�g���������"�uJ-V�6#/-s���r�J5�lT"�H���xQ���$:�  �iNt�Q�'��x ���7:=p�����7~ "���f>H��0�K	%�$�X�"G %�"�)�¶|�D�(�H�]	%�P��
K���`bTe�RN<��i~����i>]F{�.B��ͱ�c�%�p�v���y2iS�]@Q���Ԙ���`�B��y��'��"=ͧ�?q(O��9W���{D�Y�"�F��4I��J+�N�A���OT��O��d�ɺ����?��O|��� �I���,�Q<�a@��a���'�v�yP�E��2d#?���'�ҡ�ЦF�F�x�B���e�Ή�r+X� u��c�74[����i ��J&'@C��'#��
4 � ,ɪ���}�`��X7�?���i7�O��d�O �<�s�C@_�H��^�;H`���5�O��O��zҦ��t��)ѭE�]*����������YybJE���'�?Q �K,XX�MH�r)�+ ��.�?9��s|:@����?!�O]�q4a<MO�9��4����V$E�E�Q L�M�<\�),�������_�'|�-آ�Az�||"#Y3ҴI��H�	�� �
e�d�l�\\��4>��|[��$]�ob�'�ə�Qʁ�� �س��qZ��>|O�$�P��UP�a ��>��Y�wO�nZ�Jn2D(�k[����feʐ�IBy2�I�T 7��<�+�D����O
�IW��ulU@�G�>(8�����ON��T�c6Q�C��@@TIɐ4u��1�ǐ�v:�'l��1C UT�ZT!"��f7��O�		Ѣ6@��\��+�1�l+�O0es�l�~�wB��m.	;��8L����Pw�׬q�2�'��>��I�|9Dd�e�C�uk�޸/@�B�I!g5�ثK�(����
�
����$�b�'�pu�(�#�T1��"�?:A� ,w����O6�d�5U����$�O����O6�4�f��pFU:�~	
�O�O���&e۳=T�r�W�`�*����wTdc>��	�?@:�d�]-Hi��l���~���.�39R�m���Ԝ��y�sL�|�НrBe�B�SȦqrBgށҤ�,�������e��!a�Lڟ���ПP/�ܟ�>˓�?QPN2��-�T���>���D��xR �?G�B�D�HA�b�*ҭ����d�n�'T�$�'^�8.H0�����4-�hx��X��|Ð끖6P��џ����8�XwX��'�iI37\415��)2."�J���U�z}J���fH� ��2 W�-6�'����$j��54��M֟@P��wgV?x�V��R��
��YxWcW�0<1���>kV�{c�Џ�@h	�l�p� ��)�MK���?���?����?����8m���32f�\ ���-Lv"!�� ��)�mK^�����(p1O�`�'���1�����4�?���l? 	��o������l�*,���?��˃�?����t�8��tp�l� ?K�ma���a��`
7烜tC(x)C��Q�x����8��C�T�كR�Y&"�Ċ�����B�"�'ن=!��8��I�:Q,�D�O���O��ؐ�>t!��*ua�2�|�u��<i�����.eP!Bױ�x;���:��`b�OИo�*4E�l�"lE,awM� !�t�d���Eyb.�W�Н�!�'�^>�8������iU�����R��!��m���	�y*�
��S9+�\<#S��^'NT�^w��A�X>}�MN�� ·6x~i2Q(3}"%�?���w$�/	1B��Ǵx��L��4I�O��9	∑ F�*,c��]w^0BK�XH�"�O��lZ��'��'"��)� �+���2��3@��<�����<� Xo 0���Eb���
�u�����Q���KРm+��I�@��T���l�ݟ���ܟ�8�)X-#������	ȟ��ݷm9A�L����ez�cR�\�Pj�hߴ!��6�3��g�Pߔp�0� �T*Ld+Q�D3�>m3�K�� �x�Ą�&dĨ�I�rܧ3Bb��Nw� 0�d]�MCp
$�"Uh$Ġ����M��i�BU	\�O��<����i��J�"��c�? IDu�H>����� L��lH�5��U	�H�[�q+��|S�4��f�|2�OE�U���ƫ�?������*U\V�Ѳ��-��0@���@�	ҟ��	�?��I矠�I8����ƕ�vuI��.�x�� �0=M���0��n,T��' OP��ucH��z���$Y�xrB��&o=Z8B�M_(>@��G�5�&��%�ɋg@I��&�6���+bLTQ\h��*�O��n��M����?q���?���?)���"Q���bvXT@�0T�h,��������Ss�D�-�9k<��e�},��$����4Z��FZ�����ԋ�M����?��&,f*p� �FP�dk� �?�� F\
��?��O8��B�ȭi8b�b�&@q�N�l��K�ٞ2g�l�G���u�$"?!�Q�K���x��W&u� 2'����	��lU?��𸐆ؾZL�Ԁڴv�Xe��&�B�c����	��M;�[��B�"���l�_�c�h�3�	���I��?E�į@��<`1 �j�`ݙ6ψ��x2@�4@1u�G��H�K ,��>]�ro�O��
��m;f�i��'	��:5�]��N<�]���#�RRm"S��X��͟`�%�45����I^}Ji���QHD�)�|�5G]9h�^��E�M�{@��7!X����L�a��L�ʦ��ԋU75ڴ(�;9H�m�$�2�u�Ō\��U8��$���5�T���I!I��$�MjI|RL~J�B��u��U)u�(���]D��?Q	�;A�0��^/v}�ࡍ�UǺ���4��XDz��Փ���J� %/68��c�Z7�OT�d�O����T.���O����O���bhj��K 6 �pd��"h�H!�>!d�p ~�^1+��&�3�� ���m ܳP@0�L��GT���͒Ii����p��IzU��|�EÈoV-2�J|@rϕ%|�26�ꦡ�ɀ���)�<���|���@�[1��#�Ԗ2.l�n94�8ƫ*J�ę�Ń�\'b�R�9?q����?]��myb��>�sg�·>�N����f���e��'�2�'�bk�Q�I��'��c�g۬|I��R�DC/H�d���%6<tkT�P%$'����'A-��O@L����Gň�I�%X~���㖖d�dx�1aQ�*�v�;F��S�iѵˈ--3�u��)��hm����чR�t��D�HI�����J���3ݴe����'x������?�@%�r�hEd�2z��7��i��$�l n�-A�L"AR�xhd��%0�	Td�	ey���e֝џ��	�.�nQ�k��QD/L�0,����4	���˟����|��|um+�%J1�ޅ�SLG�2
��ar�m+�JK�gU�9 xD5FU@�'-T]�l�Κ�x�$Ҳ͛I�*����� C&�p���D� ��r
��p���Kz�'��X�gx�v����$ʈa�x�I�`�J����"C�3"c���?Ɏ��IKQy�ř!B�N����C�S��E{�O�|7-�F+�xZPHZ�0� p�c�$kG@�$�<�cH\����ԟp�O6JMR��'���BS�4ƚ��MH!I(T��)�O����V��4�g�I�-���#��s�ʧ����F)`���k��.�Rmr�.ƹ��E*j��bPAk@QA1nզQ���TB9+�`��)��Z�h]�S�Ϊ��ɴ}�t���ܦ��ش�?I���NA��T���bV�>�LA����'�r�'MfAH���'��	����+����i>͂��M�V���p��v��#an˴JgN`�'���'���"0LI"�'c��'-�ю���h�,v�n�p�պA>p�CkE�t�c�HQnO��Q��]�Hf(��Y>��tk¹! =�%�	!�H9v��J�2,z��I��b|�	�#�jye�
\��ch�8R%L0b�4~��	�B���4����+�I����_N��d)�8]�C䉄v�\h�è@��1�v䉮%X��y���4�ڴ�?�.O��;�NT�v!����+J0G:�p�6��.�B1�"�O����O,��뺫��?)�O+|��DU'G��гs9*9�Ę�|K�%	l0҅:V���':P}���ɟR;��[QLR N�0��y� � ��ͽ#�2��$��w�pa�d��@:R�?KD�i�����f�H�ˌXؐ����Ɵ�z޴n+���d�J�'0��-�aܱ6�59�-��!
����IX�	 ���[����9�rg�p)c��:ܴ�?)�yB���F�0w��,�AH��B��2��I>�y�m�2N��Q�Ǉ��>��dE��y�KI�_)���7`B#�����!�y�bQ�)r���	�S(hg��y�"�3)����,9v+>0҆�F�y�k�P� w,Z�jM&�G��yb�B�-�Ҡ����&2{����$�y�f�:S$p�#gO.O��
���
�y���f�u+&�ܱ+*����ֶ�yr���9��L��)!F0�q����y鞤n���+�ɯ��Es���y
� �����[7LJ���~Gv5;�"O�$���9��Ъ�;k>��"O�Ba��3:��BTo��0|2e"O��C-H�v��<�eNE�e�pۀ"O�y��&��%��L�3��Mbe"O����c$O�|�q�k�3@�lI�"Oj(2�-Y�B�8�c�B�l�t�0�"O�}j�n�z��8Y�gI�d���"O�xiƯ��m�� ���6-*��"O��DGN?kL�@�v�ީZ |XyG"O�@�F�\��6B�T<Q�����"O��q
0�`T(�bֿ/@|�� "O�1�.˨O
P83�
��P]�`S�"O4�Je&�IN6�xӨ��91ּ��"O �����O}>ဓ@"���W"O���S؂�&�ɤd)L�"Ot��%܅rr��1��?���$"O�1#�dC�\�Hu1b'|��ay��>�f�x����f�&$�m
����O��ݛ��+	p�@��h�
kq�� �'��Ĩ�b�G:���5-����`'Z�*�\rP�>�?���H�͘O!�X�O$ɀࠕ��<=�qM�!&��(��� �)�s%A$G-ԝ���Ѭ+
�����;��$���I
b�ݨ�#Q�J$,�	�R���V-]	Ulڻ{)�%Ez����P�����M�Z�B�x�o�Q���	�捏}��E�Q!���$4ړ� d 3�*���F˕C��qGP&2�pd([O8�\yեݰ+r}��eELDST˫<ɉ�4�V�o�^tk ��d��嬈�w�����0=qRLݛ<��\�s�G�@�.���a�4�d��KX�7��
��f�'MBP��H�G֪>�4{d� ����y<�	�N�c�e�b,֣U���$ƃg�C��it�3b�AhF1OP���"q��3��|HIA�x�o��cx�% ���"
� Y &���'�X��$Yب|��hV`l�3#�իNɒ�#��ڗh
fT
ӓST1k�^$�n9s� �z4:��5M��C&�3�����0�+���6N�	�T���Sz��dK.6���m�f�:�;�,�0,iD�"�<lO��P-����D]?�z�z���+e"��S�O�Qџ����(/����G�|	ESӇV"D(ʖ��9�8����?� �>�-ҭr@�1�'�.�spW?h�~�CB�%�uPUM�;�@P�\9]`
I)Od0B�Ś20et�+d,��TT�FPԼc�88��N>6x8����'zN��Wd��'���!�O�=�w*֞"Iv/;L�L�w�7�`Hb�/]� y��2	�*y!�֠d���q&�c	az"I�8���{��R?XY�T��s ʣ�ξ�>�m@��O�iP (^
7��D�P(ܥTP�ʧ��'�����q��rT��@�Hq"�0���ע��豎&��')ԩ@�̂��Đ#��Z�<9v��4�(�y�\)O��%k�b�&��'I
��!��/;t�!� �ݻ2%<\铤Q�l��	3��H�� [�q�P�N��T
b�h9�uxGHE�R(��ʜ�w�d<�kL��'a$��r�B����30���@��[5����T闋z�a��%���tk�I�'�d�&"V"Sӄ���Ő	Ԑ��C (�b$01E���J-��=�f ���S~0b�m xm���b��x 
	ۓ~�P� �M��?ޭ��Á	>�;V'M��0>��.ٳz�}�������j�C�@�3��@XT�%���ImyR���J�|� �� �C�aS��)% L��ӞJ�8}�B���w�����	�)S�`�WA�o��Tp�&G�R9��M�?�B�pgL�?h�QʀF���I���[j�ۦm��Q���'���f��rM�%�M����'�pJ� �4�@��Ѕ̀O���F|��2Y�(�{W*�{ �ɡ7b�[�n	�ՌR�7%���`�>>���1����OPhH x��ܙ��ɻi0Fհq� ! �l�~�'pH���s?�u� #���f�<n�F�Ӄ�E�W�g���7�A<T ��d}�9:�m�
FO�A*e�[7n�N�D�j?yvB	\��� B�P�2M�c0�pA�
�F/P�V�ŊV�Š����E�ABF~b F�r����o\~ҴiԼ8H4��g|� *�+M2b�P�O��A�hV�$l��D��7G	f����< v�FN�2
|�Dfa�._:E7V��% :�Ԡ�6W�(����9 �#��>�{��y���QW�H'W����5�Å5h��1��eU�u2AbH+S>]Z�Nި_���YZw\">y��ER�q�E�(t,-�S���W���U,U?g�4=�?E�m#!�� E��3!�� ��|Q�0�\l��0ʛw�R�h�+�/N�<P���$~�xK>���$�������w>R�j���5�l�3
�XG����@���O��Bdm����8fğ?G*l�I��
	e�"@J��'�v�J��1%z]�?9�lqӔ8�!��^�����#���q=O� �8�49�����ϻQ^��Q\���� �]�ތ�F/��"��k����'�*�� �?\�DI�V�gŐ}CG��ܟ��aA��,U^�sR�4�뮓��hObm�#��q���[gK_#k�f�i�,Ɔ�~���:��'>�c�ŬY�����E8c�8@2���.q�Z͘q�P�'\�1�s:.�]�2����ƙ�mَy��Ĝj���O�x��4�i>7�
�}qʵ�2�M##p�2ck�+$�.t"��B���'Hi�T��w��Kc���.����O뎖�R���9�`إX$e+S�M�3�'�:h�֦\��?qS�t�����,��t.͟L뇌F�..89�cQ=6���CΔ>Hh%�抃�{��a'�������'4�'O�#9䄅�&/ʘ�~5)�+I��<�GFH�/r��k��F�F<���hO>��s��!3\yӈ�8\�(�� �3}�!�	$�1��<b�ON8&��e\�-J����	42���kBn�'����MY��>��B.K�I�A���-���[B 
 Lr�I>YF ��S����O�r퉕,1�U���G�a�^�����6J�)��y���
��(���@x�|e態��8Sސ��bUμp:q�K:s��sO<���͕pf7�ʹwd����O�oN��������7
��	P���s�vؑ�D�3(���{���@��;�e�=Y�4=%���?q�#3����DZu�H8z��/�?1w�ߡʤ�RӀ��g�0� �C�'��y�/	r�iW`��(p�eqL>i�B�2B�j�G�ͭ$�Tq_�h@0	'�@�����F�Fު���!Ds��c���K]H��h�ǭU< ��'U��ԟZ���#�H��`_�\P��8#���k�.Q	������BCB�(E{�����9�ӺC���Bn��GoD0z!�����K{���?i� C#k��݀A�Ψ tBmٗ��w?QQB�,�T!���[!5�. C �,Q��q��D[��P�d�B�RUJ�|�?��.oN����ZfءJ��?��,[�N��mF�]*�9��N�'1M�`D��(��D�@�"C����K�4N����\4��'���?�qsbƇX����璸L���Ib�?w�f}���DxC�_2P��y�����牪L	��1P\�CTVI!A��9S����R�R�?�;0)Q[!������_�#{��۴dO	U`�0�1�	�^NLȣ���~��u�3�O�2�a>����/ڤZ�Oܥ��4;�n#�I�&��m
f��+�4�K�����V�	��td�l�0 ��W��,�f�\�tI� �F�"�lDB�O�� �|d5��2)6�t	lH,3E���QMpS�̂���yy��0W�
�\��%3-��|����x�G}2���oa�g�C0������~h�K���R���p��i��ϗ�u�� 21O, Q���%��xAH��=��r��0ex@9Y�9f
����Aϼkt!üf'ܰ"����^�$�v	
�F�2�ir�2���DRQ�}=�H*��4
>��2-��Q�� {!���>��#<��K��Z�������O�v5�f)̕-�V��!��h�2m2��J�M��h��B�k�F�(�S8���'�J�K"M\9/� -3EA� o;j<�椔�dRĔ�v���)�q����럒�#P��H�i�:S��:Cܐx!�8 '��46��7�ލsT��]h�'mZ� c�$m�e��AI	,�A�'��H��nO��D�v�B���O��>!$-V6rH� �mS%7���"U�'Rbd!��?O�!��D�n�.O�IJ�u��%\y�Z2h�3@��,L� \���e�O�+�lМ' ��k7A��'�|9��:;��ZW�
�zH�"<�RY=i�<��v�;4�`�>��Ud<fN<�`�ʎ�p�,9�h �ɳe�����8L�y���=���ɡ�4�f�֚f�v�S����󎌉��A/�j�kBdGe;(�)5�O��<96.�����n��ƽ�rII�D�#���%?o6:d�+m��H�ȐrMn]�_wQ�P!��+TXrH9�kN0��x`�p��@�-��c?�� �H����<�O ���ޭ@;�= gĤ1�tI�b�*bq�����cX���ՄD��]�TeP�&S�:�@ƹ���DE&e�P�j6�O��p%ӭC��ɝ'�'&�IpE�F�f��`۵�Y���H@��dD=I�L���ĭ
M���~��b$Y,8��L\!�M�vĀ*��@����ny2I�1���&br	+D�~z�.�1?�]j�- ~ݛ�^�'o"��H�7)��@.O���kl ���δp���=lNZ�IVa��QD� B��L�����>�H�:y�$�|�<��BO�m����¨D�XpPq�^�<��/�M��'&�Љ0�����4�	"YUr�i4N�*E{�T**ؠ��!�Q-�c�xR�� 6��HW�XFxwf�"}���l�X��H�$��1�,��A;��Oba3�+���5��R�� ���(O,�yt]#�O��i ��,R��J��OHd�1 GHր��pgԔ�\P�.-ғ6����+@Tx�7bZ�'�.)�'��9	���?�R���\�fh������p�p��*����|�ɿ) I�P�Y�K4`Tͧ;�LT�DU�*����*v�˃�ɝ
�*x@��K�B���x������>��m���V��*$�jhy	�&�Z��b@˦�R�'G2!B�Y�tS !�[���-��ƁV|��nɣ?$��!R��+8`��dك���#V2��p$�52���OG�T�x�� ��O2xc#�Ds��	*�O{t4J!��I���t�\�m�z'ؘGC�$���քB��ԘT`��@[�0C�^�q��Kt+�O6�IC�$h��K�D���h�Γ8��qLÃb��D�Ύr�<Y�ǂH0@4=*�Z� $��*ƣ<��׸>#�ܘ�/E?�i���!z��7
ح	xR�ae�6������<� 'TBXHS����% j�� �@�f��2F��1�V��+E�4��c�,V�(a�#.��P�B��f��?�6  ���8 m�B�\(�E,*�� �'������\\aA�Y��J��Ту	��ԓ��B9p&ų��J���R;y�&ı�9���M]8eS�!�f�dF
]��ۓ.�ĥ�e k.�чT�q��$1��S
1T�U�R,y�Ru��K�D_X�"e�8�O�] ��rt��4�Z	��jA��,��iСA#b�P��ò"�T��j�=[�&�A�,� !�� %j�Be��%���`�ҀL�2�b��!���5F��A%��b5�*�"p��	
a]�����<y'ʑ(X`U�Š�:@��ח#u�9bsƊdAL�2t��n`||;V��v�C�L��Dڇ�"$Υь�s�*\���\�=��V�\l����	WYf ����yr�̔��ߩt�(E���@�X�Tt	v��6D	l���[�{� H�'��5�SIH�yd��1ufn_:4V����B��yr�J���i9%�L�Ê˥jE� ��H_i�v��k�3�T��
�0H�<��D%��U�CU�����̟|�B�P ��vm��#�e�I�5Y��Y�YH��	yt-C4�aX�[�u����a+�I'o6��!���h������	N��<�d�J+6��%���z�ـ��m�,T�`hR�\YP��%��%\����~w��ˑ�:~}�E��h����reI�b<[v`	0ʼ�I,�n߆E�$Ǔ%��C%���@	���iP4x@r�d+tB���$��5ϕ�D	i1���j���`�C�>�y��H�K���cBF�fn`�j0j�$�u��i�-$���'��&'����C���[���h�h�,-��X�c;��AE��|�aǕ�R��|r��?�Z=�o�8R$.h�`H��q播�}�H��F�ݒ}��i��P�>J�����/��[TOX�c)`a�f��,���Ʈ�|�ҍEznͳ� l 7M]�(Jy!ST�r��I(��,�Dтy$�1��P�-�v��d�2 ��j3���:������� �H����1N��]�����M��E�G�]>>T�I:9����زY|뮜�4�Bx��k��&�Da�l�'=�!�CJ�*�A�
U"nࢴq�c�$I\8u�P�=.P$��'2fm�D�R%-:��O�ڹӵc��y7\�W`�c��!i�8%��̂�Px��&0+�0�$�
�q����<F��@3��J��[c��.NZ���g��/p��1� ��1�O�����\V�����/E��Pbd"O�(��N�Ew ���C�;x���7;O����.H4���	s���9EĤl�D�h��ދ9fHC�ɣv"`:D��5�T͛B�[g2C�-du�z����-4���>�C�ɲi��A�H��[(n{��:xC�	.>$��:�+��(��	0�ƠK��B�	4k�@z���,|v�s&zC�	�Nƌ!�L�c��MN0C䉖
��r`V
��)�2ȶCv(C䉑&�(阖LL�V�y��G!U�C�IR��%�&�P�^��3��C9B�	L��tc�0���/U�C��.}$����c,U�v�$6�B䉺h	�|)���|�}Ӏ��;tS�C�I0K�FT;"�T�S�MB�\�#+�C�I>o�P�ST9Ss�τ+s�C�	,2���z�@���j7���B�ɷ&��y�`KE�7#za���RB�M�	����P�6�Eĭ[�`B�	�{$8���C�Fh�	n��C��:7��(�ݎv�ij�F_#�B�)f�-�B�E�=2B"C�~sFB�I�~���a�
��Rw�M���3>`C��C�F��ߟu�ح&�ʾW�zC�ɱHL�w���:��!XC	��R��C�	6`hḥ��,5f`Z��GK�BB�I-t�g�'�d��n��<#vB�I)��[�aQ3DIJ�JB�-�C�I�k��
S%�	RB�\sj@�i��B�	�?�j�9�	,u#&�z�^��B�(p�D,�!�[�A|R!xP�Z�x=�B�/8��8�f܌&��+���~�B�\�\(ٰ`�]��Ń3��C��1qp�x��!+>S��u�7mb�C䉈�|�a(T�P��=�B��9LRC�I$r��8�i�1����F�|��B�)� �	�q�؀NyTe��dK�k*���'"O�]��fL�X��` �P�(�D�"OV��J��w
DMZv(E9	�)�"O~��vŇ6F��剏�T^\���"O^�x���2�|��晛NtMӒ"O����%I�x�`9����<,=��C "O��i%f�1��j�!�5&x�@"O�lX��x�0)�22ϊx��"O��AmR?I�N�� ɀT�
���"O�dٴ �3q��TaWm�!��-Щ�HДB��T�fL���!�ƵU�X�z����H�s�
�>w�!�ђ=o�� ���Y�^@G)�%�!�ˑxX��"�ʟ-��	��X%?�!����i����
��l�E_!��f�p�I�"3�
�;q��S^!�䏅-�Ac�{�fH��:\!�DH�}��yڣ �! �Ah�=7x!�D�=/���QJd�lؑ��]ea!�$<D�A��i�&���f wN!��p��r4�� ��P��HW!�J3$��QcT�Y�y����N!��GB����)�y���gD[!��.K���Q(S�IqJ�{Ѧ��k6�=E��'� A��@���ѳ蝂*2ڰ�'Zq�U�J'Te Q��&�N.���'T���)=I����A�LF<�Y�'�FUr�'�(�*yx�ǫB��)�'܉p�?���b��Ý:�"l�'A��2/6k�șB��+E!�9a�'��Ċ�HYY�pB�D�9���	�'�:�B�
ׄ3G88�R&ِ*"�h�	�'] 쨒�&t�("�\�!�T �	�'"(��1�:��4ʟ�N!�][�'{.��qB�yB��Ĵ;<�{�'�i�F
E����F�4����'��E��C��A!��&ƠK�'r$�C��8��룍��|���'� �Y��BO~��g���XIS�'��XA���|����",��(��'�:�����+ 킍)��##��%pǓ�HO� ��,]�F�P�������"O��82f��@�d}:1o�<Չ�"O� ,�9 â�e��?P�x�Cc"O� ��ȝ��  F ;B�6�� "O�(�D�����8#h�@}���6B�B!h�h���9�N�c���p��@�nF�]  ��ؠl�!��7#��%b(?p�-���I Մ�0%.akaj��VF��5�k��ȓ%GnёP�OU�(j�MĔ^���ȓ?x{a'��<K�&�}V\�ȓK!�5�2H�.�~H!��O�� ��~n���Df�z�IQq�ĳT�l%�O ����H�����4&L<<h�c�!��;C�>�*���i��!I��\�f�!�'Z�L�1�Hԇ\M�c$�V�ў���. ��2�!?f�٪Ą	-�B�I-:5�hޫ~+&��M"��B䉪"������#!��H@�vC� N��IX`��_��D@G+�'��B��:_▕�`
�.���	B�B��B�Il�]P`[���5��% Q=B�I�L�U�v�F/�ޝh�n�M�B�)� 2�I�M��N��	Vn�Y����"O Y����l`��ɚJʬ��a"O�H#�#l)�H�%�,���"O��"f�*~����� +��|*B"O�rwE��#���"QkI�N�Ʃ��"OBXz&��������L]��@�"O`�wB̅o,� p�*N�RG6�
�"O�A����W���:�j�9���A�"O�)��ּGF�1����qF�F��HO?��>_]Ҍq%��f{.T��`�LX��$c�$���&�T)�Wlұ�yC�r�\@ƭ_yDZ=9� �yLB�BJ�5۲,X#m,������y�،Z�v��WIL6^�� a�_��y��C�CVi0�	Bs0t�!k9�y���`����I<�$���j���y�I=n�<d��-h$�K��@�y�?k�t�a2f��>�j�JΌ�yZ"q�qy�L��[�p�����yb���(�b҉�,S��MJg�yc�?c�(��-�QS����=�y�T��T��ۨJZ~��u�١�~R�'n�p�ZFȑ1j5T،��'.�dg 
����9uXI��'���S�l�;(N�3r�U-6b�'~*ɉ��_�]WYئk���]��'�@��$(�9YT0VB�~<��Y
�'���l���]`����u8���	�'
I�a��h��2��,#��H(<Yߴ�*�E��;l �v����v���I\�i�8�/�3��*�+�.G�� �ȓ>��ѳܾ\՞�A��T�f�:d�ȓ"����`���N����%e�,FuT���A���P�JF1&�n١�@�>N�Ez��'�:���فb��;Coʾu����'~h�R��ՌE��5����6sj� �'��-kf��&k���#�f�f�J��'�P<�#ˑ*h92�T���G �$����*�'VD�HQB\�*_��������ȓ7�`i�� 1Y�.����
�Z���J≀lmJID���z�|}yv�.F�C��/������� !+ ��0��n\�C�ɢH�&\i��{����
X)C��Q���V$�Flȑs����1� C�+���a(�D��}�@h�_�B�	�q�\5���S�[�|�4#J� H��p?���ۼ1?� AG��h�`0)��	e�<�����0��fS{�IY5�`�<Q�+КMC�"Q���7��2�_�<��h"��)bgCW:���3�
Y�<!�OK��Ȁ���X�R�!֤	`�<�7
�:-���C�U�d�FmQ�ΟZ�<9R��@3�h[GW1a�ޥJ2�U�<��!B�la�Iͫn:|E�eNGg�<�A S�TV�2E��cR���a�f�<��N�}{T�[�l=r8ʷ�^b�<�4�	OTeU��w�4��hb�<�L�j�
�b�>@��JhEv�<q��H�e��H�^�{SK��,lZB�ɰ*[(����}������&��C�	5Nc� �G��%LA|�Y�l�z���	}����
ɛ�$(����F���т�"Oj:e1��`�V5��\��"Ot�qt◩^J�X«�!��4��"O� ��)rL٠K�iGkB���i��"OH���|�R㞛^�V"O@ $�2E�N�P-��Q̊@�2ޒ�hO?�	��"��M$�hB�O��gRd��D%�	!R��Q�'��dy����5P�BB��+�J݋��0i����������d�>6�߮:��[�ǵM �Ij��_{�<�`�h��(��+�~'�5�p�z�<Y�j�� �q*Ao�����`eFL�<��n/~ ��b!4]D��E�<)co�~�"����R=���1	�D�<Q7g	�"Jд�d�� ����.�C�<1&ց��H�TB�X��HbD�}�<i'K��D�P<���:���M�<�®ǣf$:�Ǎ8Y��[q�Jt�<�&H��BI����� Q����E�<���5�0(�� �H�0X�!H�<��hPw���u���U�����@�<�ң��3[��0��\1b�:QViFF�<icG��(p��(���|@Ö�K~�'@?��mƍa6|�#��%�ju*s;D��S������ �a3�|���:D��ifbٳD��A
��L[l|	t�8D���h�H̰ u��XImjr,2D�lyA�B��s��Z�^�@-���0D�� 2�(yt<z�#��O-�%	�,D���7��.6,\��`�5~^�A�6%5D�@��!K~�Ց����5�#�2T����c!C'Ε ��Ӎ4h�!�dMV�����,�A
2ى�lĭ�!��-��ys���!]�(�I&�C	J�!��~���N�j���JK�!�Q?5�٪5�X JPd��� %E!�$յ.v��J�	a8t��E��%9!�dګd��]�`���<A�5�H�9{!� ��bD���EZv��R$�?uo!�DZ/z暸�f ˺l�1f]�:Y!�P�	7X�y�a�y�n���T�Am!�ľ:����`�&�p�*�f9d!�N�C��Ч��]xY ��	!�d ���t�ѤV�yO��ծ�4#!�Ē�^��;�o� `9��ٖ.!���}�<�Y0DO�J+�u�S�"I�!�DC��{�L��ᘳ7�!�
6^*<lrIɥ*���8�AL��!�d��f_�y�lQ>nǒ�ʠ�8	Q!�$�$u
��3�J(s�� �a��x^!����RvJݠ)�z�BC�N�Aa
�'��t;��W�:nRH��Ŋ"n�|���'馩j��^6���%F�4`����'ζ��u�k\��+r�&+2�@
�'G 	fC�dpi�an\Ɏ���'����g�"_̼� jW�n�	�'��G��Y�JT"��L�
���'�J���O�0����Q�	9�+�'��K�a6(�<sp̲O���
�'ن�bsa���<Ba��z�x{
�'���:e�R�aw`��@�m����'S*1�gC��p��@�7 ��Q�'��T�A/\sx�)����8@/�T`�' �R��/Y���#�-	,i��y
�'�^��$�_�F�� �#^�
��2
�'@�ڔf��kl��� G�&�a�'��u#��ӟd��'�|�*���� 0�+�Q�#B�ѧFY�>��	�"O<�� �U=K�ƭX���O����E"O�AD��$���0'�qjY��"O� i"��Dzl�F͕���D"O&�C�ɸy�2�2��Opߢpa�"OL�k�R;�F��e��(�ʝpC"ONH:��?\�g�(Ӗ�)5"Op�
����GJj�����%���Q#"O��3'i
�6�
%�ݲf����a"O,H��A�a!����2D��"O�Y�0�^�L(�����D�B`!�$�z�0̺FA�(j��P����t'!򤅌A�Zy҃"�/��K���1K�!��ЭV�$���*;wnM�eۡ �!�$΅0�`��ϔ0��*�
p{�!���L=Xrr,E�TL9��"�!�$E�4�Y���
u��A�L��!� V�,Ӳ��1Ь����x�!򄈱P!��7⛵>�"� 4��T!� @�Lt�d�-�N9yeA�h!�d �d�*As��N���p8RK��!�a_�c�l��wK�800*�'c�!�dӞh�(-�`JܕWK:\q7��1p�!�o�T�fB���T-־qC!�$O�SP��M�.d`��w!��S,/�T:�S�w_(�R�-ʇ_�!���48Gǒ8>� ���\�!�5c�.U�0�%! acJ�@�!�d@�+��}tKH�/$Hx�RL�2!�dK�d�Rm#K���֌��$!�d�O������#�H0K��p�!���t����4艧�J{3���r�!�N.D�����70��IY��2�!��<i���g �7�$�PQa�v�!��J�R�9G#���d ��ˋw�!��n(�#Jĺ#U6m���R�r�!��̬%��g(؄-NT���u�!�䀮l�T�:�$U�c3H풦�A!�$�DD}��hɱO0~���I�Z!�$6P���iէ���DR��!%�!�D�{����̈́ �r��aB+x!�dO���:b�ԁ	�عʰB.Co!�.G�]���D<���y�"�F!�M5)�b	IpoŊ4v�h����}7!�%e���C�׊	 ����I�$�!�Ā�A�!U�+��l��dQ!�$�z�x$�l���J�1Q�M6A8!�d�;ɐ�b����C�,aCBK�35�!��B*���K��t��� :b�!�$A�lޜ����{��Ui2�A�h�!�d�X�r80t矵dv�(��n�+n�!�*3HfD��#[�\k�����ۦ?f!�D�Q��h�'�@-_0�%$ʜ~e!�D�jԊ�a��V$¹[��T%c!��?���*B�_(Q|\��B�%%8!򤘮v� �Q�*J�J�L}q���r!��#";�(9����CQ܄ T%0(�!���&_�|�BG�x�ܤ��m�#b�!�d�O�4��uIۂYŘ���!��=9іFC9V���K!9�!�$h#l�s�a@�"�$��ąG!��-):8<���X��p2�$L�F�!�dF��p�f�{��)��N�(�!�D�.)���{���V� �bOH8�!�� .�)!�ŏ8*����ACgR(X��"O4�ȵ��p��J�`��oF. �U"O��"GK&�Q6A�.!'�d�S"O�Q�����I"��w$4��R"O~ )0�@�0:��e�au�e�"O6��E&��@P0�3U}E��"O��Y�� ^�2�� ��y�`�q�"O:��`T46L�"!�
3�D`!"O�az�<e��`�?��9P"O�ȡ�\.D�XC�N�{s�A9�"O��&+� Y����7�=c�)00"OnyQ�'��C�;O+��2�"O(�r����3�V�����&jM:b"O|f�RD1�H�>�P��G"OY�uj�=)�R��Ƌ�1z�Jw"O"��F��V|ct*�"%_P1��"O���#��?��YyB���YY�)(�"O��贪\�ot��[�	AKN���"OAZCgP�B��x6I�=SJ%`"Oxy{�.H3|���fG̹i(PXP�"O$�B4�\	����#�](V̹d"O����"�0�B���#Y��"ONp'JK8{.<�
��F*#��Qq�"O93��w��L�e�ұyބ�"Ol��Ɏ���
D�C�,<"���"O�]p�E�R������χ%�š�"O6�A�v��d	��M��d�%"O�51!ϟ�@�[�$�2p�HM;C"Od�`���'th{&��[��Y�"O�����P�{��I�(�"l]x�"O,!8�Leź����@�c	2�37"O��k�r�F0�7eB8!$���"O�F��(?Ȉ��D�n(7"O(��!�F.���C]�2e<eCC"O�Xʡ��$�~��!e+j��s�"O�!x��Z;����DX�bH����"Oa�R!k�%�g
N��h��"O�T'�!zP��&�U�[� E��"O>p)W?
�e�ɾa�f�a"O}��O1)zJe�/ͅ.�($B�"ORIp��;��Ju�H�s��Yc"O�x���8]4�X�mƽ4i@$�t"O����E�9ƪlK7��(_n��"O`)	b�N4t�ap%�1fMba�T"Oʩ)��;y.�����=�A�"OR��l��N|m�����/.VI�"O��O�iinqI�
��j(B�H�"OF�P ��#B9
 �Z	1 t�""O��{5��l�R�0D.(w�D䑧"O$E�'��&����V�R��aP"O�Ԉ�L7�� a1�ܬP��X�"OJS��P��qwJ��pm�6"Of�z���}��Á"t�ȔI1"O���ƆG�r1$�Qqh��G�	r�"O�{�o }�nO)��
�"O �s�-]�YuV�Af�ɽ��G"O�زdix,]a�.
�x�|��"O� z2���_�NIs.�7S�bݪ�"O�5�/|k���M$`��D�"O�8K!���<q�8�F�P^��e�"O��`R�Y�s��YW�������"O�mB��ܚJ�x5x���R�^0�"O:��o��/I�Re&Xђ��"O�|@ b�L*5�e�WY~$yR"O� bqcЅM&W���	�"�FS�D�'"O�@���9� �L��t)�t"O��v�p2�в`��_� ��"O$H��֪2���$�)E��"OT�B�J�*
�� ��A>i*~<��"O�]s"	�F�<0Z�c��S*�IQ"O`��M�%+xv�"!Fؾ-�"Ob1�ąďR�6�y�(-=�\�#"O(ܱ���'S2AcgyT4�"O&Pjeֲ�^`)��P h���#"O���Ge�1��{#�A�g��5�"O�����W�4�9��L�dC*�t"O�a�dʄ�0�����0$qAA"O�Q)C�	�2��Ts���\���"O��� D�m��,��L�mT�0!"O��C�,U�Z2�P�pk��2;�@ "OR�;W새r+�����!"��b5"O�i:�H�[f&�Q4��+4؁u"O���1h�.(5T�3�ߦNz(:"O�ًħN�X ���b!�IV�B�"O�y�׮;JX�"ᆲ<� 4��"O� �D�R5)`>@C�Y�{��=h�"O,���*ޝ{�*�G�Yٴ��"Oz��
Z"^�HSȚ�,�j�"O�љ���]�hhS⊧iT�T"O�ʢ��*������5��8z%"OLRuG��!��$fج(�"OR �5f�8~hx��O �{�V5�"O�ŉ&Ϟ*n�UѠ��#��)�"OxM�P��b-���c���H�"Of����df��أG�s6(1!�"O��G �Tn���$X $���"O�ds���A-"%b����x�@"O�	��/GV-�)�W(�?Ҙ��"On��6��#&��E����Y�v�#�"Ol��D�ƴY��!xf�N�o���xf"O� �WM���ti�&��
b�&�"O�m�IJ0%hSQeRMP< %"O�	��LW:Jg��2p�Q��:B"Ov��Áq�h���P�]���p"O��rh�!0�-�a�6Ur��F"O T3��3~����$y|p�"O��K��T��A+DR�SW"O�PDFQH�C
��]�t�B�"O8��Qm[46lJ��).&��A1"O����?t���T(v�@�"O��B �4f��<�� Ѥ8:��"O��t��?k$���n�m- P�2"O��a�聀Gp��0 ��n�k"Oک�
���Vd؃�F:Z: x�"O�T���8 '��R�E�;22 �"O&L� ,\J�R�����}h%"O�u�QmЀ,i4Ax'/��j	V�`A"Od��pCU�@q8"o�^_���"O2�XTGA%j^t��fM��mF~p3"O<!#C�tU���0*X6D��5"O�����65�tY�%�@�H����"O��`��p#D��E��x��	 "OX���O�|�Bl����!�*�P�"Oz�����_��1�K)ǌR�"Oj�QvH�}x��Td��1��-��"OmK�d��Rĉ�I^6e�U"O�A��I�S{|Ȼ�םW�}q@"O��1�Y�pJl�H�KM:K�b�"O� R��&ZP���,`CL���"O-�ug!X�� �R;O?����"O��� �6��BG�}�x̊%"O��@F!߯E�u�����w�h b"OF�
�N&68�b�	0n��"O��åG�Kt,i��	N4 :�S'"O���t�w��X�g:K�`<R�"O�i��jʋ]�����K-a����ȓ�f������Rʱ��̞�mE���ȓ[WF��P��A�0�[�E38���ȓX=�[��F��F�B2e�d�ȓu�0GO�Z�[b��]ʌ��t8:�7�\�}W�lj��˪D�ȓ��Q��/��T��U��/n�t�ȓqc�L�hL26�r�awa�gsA��p}�iC ��]�X�a��xx��x�x�CN�a�iqA/�]&�����Z�L�����5�@�d��ȓ:�1���_�&�&����[�����m�Դ����.YҦ<i$��+�*q�ȓ	�Fd��(�-e).Q�XՔ%�ȓF �[��(q$���OA6L��>���[2N�u��D_�Z+���Q�Dy����*��QǕ	1#̄���Ա+RFT:�$UC�G���ȓj���'iL�)`�C#-��m~ćȓ/"t䮟�+W���4%ܳʒ��*� ��H��=�Q��1"ؚH�ȓ~|vL����;��a��j_,V�\ɆȓW[�2RV�w�����$5�m��jG`���.�u�L �o�#.��/]ʍ��T�Ml!6C�0�����b_^M:��]O>Y�@IX �`���H�Ej��@Y�A@�G���������z�G΅4�~4�V >n�)�ȓv�9���Y�	=t�C�/�<w�<!��2�j�Zĥ�fd�Q"LŲ*X4��E7x4�Ț::[A@���h!6��ȓ���^0)�A�����w&�p���̝��/S.G dj7� �I�1�ȓ,��XRF�Cl,ڵ�՚L��ȓ7]D����K*&��'f�c����5��U!ڄ2��e��K�u6��ȓ�Q�s.I&X���ۑ)�,X��R�$�I�)ʪi�<((��\_���ȓ-H�+ �� 6�>8��݇�D�@D��'���%�G8CT6)��<��d����g�,0���1P,�(��?�e��	�+Wp( ��I�^u,L�ȓ3�؁��M3Nj��b2K^EBi�ȓwU�Z#+E�#Ô�*5�"�D݅ȓ@G����ȑ�L�N�* 
����ȓ^��(+�-^�/��sAP��B���8����ē�[���So�Oٲ���h�h�$��o���F�`�D�ȓ��})g�ٕp�� D.د�����	~l�r͗X�^���S�]\䈆ȓ�����8��ATTنȓq�ެ҅g�,%� IxU�QV��(�ʓz��u1��"?�V�dE��	g�B�I�iV4��%�s���Jp�^�W{��䃼D��$�d]���8���A!�\�r�e�E�Y>k�"$�,؝�!���-��0GB�l��ɫ��4|�!�� ��S�Q;8�����a08҂��D*O������	�����הS�mi�' |;�Έ�2��0ϋ�{y2�K�'�<�#v�A�>��
�oQn�x�@�'�
���Iۥ
�\q�Fȷkv2���'�� c����0�N���0k]��	�'�q�u	D�{r�a�b*Y���'R���/��Q���Ӫ���nDK�'��"�^Oq2Pi�+���Z
�'�td���rd����
�]��'��0F�G�s����#�/q�^d��'2ी��ks`4S�)��g`����'�LT�҂J�>�CA�iq�� 
�'�BěԂ�#<
���]\6��'�l����16Xl���[,���'m��P���N��E�Sϋ�d�L�z�'w���$i��c &z����&H���'�����	�X�ة�P���Q�~��	�'��%��Z:!�B�6MH(K�\��'�zts0O�[����Q$w����'��s�b�XX�5��;r_8���'�.	�R���b!j�L��d?����'F:�)#��yT�M�f��P/�X�'��@��� ~�ʐ����"|p�'�,�T��hw�N�C�e�CF�y��L�{�L�c���T�ܒ�"Z��y�B/�T���wZ1@n��yR�S�.:��!�{f�<�m��y���gB0�� ^�^dQ2S��y��P>Mܔp�1U�8��"a*�y�e�1lr���#oĀz��0���y�-ې~==��'��[��1��&�y��v�TH�G	�Q�fd��з�yr�̼E��y )�=NU(Eر	@�y�"�[(�ʇ�\B��0f���yb"�=by4�� �Y<b[�qb]/�C�I/_�$՛���.R%��k��a4�C��!C���BE�CW�ԠUm��B�7�|�cPL�r�ʠ�ʽd��B�I14,j�	�F �'m؝"'gG(�C䉄m2��Y�٥'.�E�&�ʀ0ϸC䉇q(������v������D���C�14�&����֔��ek@MU�4h�B�I���ʔ���>{B��bD��2��B�	�2x�,1&��A#.�JR�@a��C�	�|�^բ3g����LSɟY �C�I-��Ђg��2S��R�ܑnA�C�	$����r�?/�t`�S ؘo�C�	u�������Dj,���YŞC�	˔��@� g\Px���Cf�B��|���;ŤN���c�bYTJB�	 WP�8��l�� �֏5�0B䉦8�@�zį��<=��ǔ,^B䉟G��a˕�ςr���$�$v�C�	�39�ŉ��)�F`���	8�LC��7^|�K�鞷H�P8�%�SC�	��t���$�0�Y�dc�#xC�I�A0��w�))�� (��\�C̤B䉧Lc4�1�ˈ�N��h��/\L��B�ɳc T�f�`�|���O#ȦB�	kQ�ؔ�T�<Dm��n��B�ɟrgX��E�F�0e(����A}PC䉉5�X�"�Q�w���[�N�/tpC��!�@٢j�IWp	4��� �~C�)� �XۀE�U�&Ikc�	I��"O�T� ��wִ�qRϜ�1� "O4�J������)S���O�F��"Oy�B��I>FE�B�h�z8@Q"O2(�`�Åa�b�CG���7�-P�"O�<Zw�A�Yy�1�p��
Z���SU"O�!�0$����E�С3���"O*��vl]&* �xDl_��P�Y"Opܩ�Ć!`�jYXk��&H�Q"O�!�C"�J�TJrkܹo��5"O��d�U�QU�%�J�0h���"O�+�@���8���\�PG"OԜ9ţ]?q|:[�ǅ�r��²"O4���,9�(�'�
�D��m
�"O68��g�8��eZ#e� ;�����"O���c _�f7Æ0�"MI4"O��X�FX0'�;�$�>��E"O@8��9(�� 0ᗇ5	�"O����'&����ӀŁuf��A"O|x��È�o3�r�O��pakg"O1dd�G�.BE�ݙ8���{�"O����E[�a��aӿw^U��"O��!�Ά5g�x�;�M�(;d�Q��"OH��g�0"���{`
0OW�0G"O5��k̈́���+49��Z�"O8|S%�ۦr�B�	E�UQRh��"O� �bj+���Ѩ�8I�a�"O2y���:YZ�{F�Z!%1����"O����k�)H8V����Q *��v"O�����S�r�ن ٰ18)��"O��7��)�1�S
���� "O�z�H�4; �1錂\��`�"OP�$)�0@q���W����B���*O��:DƂ�./Ƅ��皍m�ؐ�'t�1���G��y�7d߉6��z
�'�t
�̎�L"��Cˀ/�x�!
�'v	�@�<W�
������x�6�	�'b�M �MݻKZ����ߔa|� �'�Ҹb2�ɉ\��FD�&b��'7����M/?��<F�Pv��5i�'ڔp�&��~�ޥ{e�Ď�@�
�'*�dY3��(��	x�.Z$�j��
�'�̙���?\��b X�y-�i�
�'�^Pɡ��+Ģ�ba���2)J
�'�$���8��
�<_G�lk
�'�܀����{������f��
�'ܼ��֧-k��D �g�w��	�'`�B@�:Wq&�b��ˁj}r� 	�'IN�QtH��|��K]%W ��'��QK�,M�4Ab��
K��\�	�'JĤ*�#ιYϚik�%ݢ,��X�'��15�]�Hz��U�#��8�'����ԫ�1oA�a�ҏQps�'�V�y1	�-r3
����;�m:�'�lh���#@h��f/&�N�{�'�
����8sD���� q�zp��'�x]Y��A�9�hta�Әo�$|)�'M�I�רPܨ@+��f>zxI�'W���.#耠���g��`��'a؜�s�� 	t����/[�&�x�'gF���o�+D�D{�-��	!@H��'Oq���g@ʩ��BB. �n�c�'����D@�$n�4ˤ�R�i9�]s�'�P� 6�ރr���G��iz� ���� ��5`���b�n��e��8�b"O
�sT��1,�\)4��j}�a
�"O(S��'��O��LbEP!"Oz ��"�P���p�W3w���q"O�l+aJ$}�0ŒV�4t�F�B�"Ova�s��@�|�UkFR��2""O�P1�=v����U#Q�0��C"O�Q��[:	�D���˙{���4"OD��0l
>i�f�Kr m���"O�]���֕E��A3!��Ju"O"ḁ�S�rV�z�5\ϰ�s0"O���a�8vǌ�Au!L�8�|���"OV )��(}��T���X>����"O:��d�
�'�H�R��%Q��p�"OD�R&@;@"RIf�Q�he�ȋ�"O���I]�9F�'\1j�rH"O��pAo��_���*��5���1"O���$�\�&16d�cI�?�H���"O����
�:�"�%��r��ȡ"O��4�R���UfD�V���g"O��CW�����y���ʧq��h�"O�!P���`�b��d�:|�b�i�"O�����^=��#���Yfp��"O
�)@a��8����E����"OR=@7��@KldⶡK�ؐ�"O� cĥ��H����Y�z�νc�"O��0p"*���!:o��tf"O�I;4� D<T�r oĿy��R�"Oҩ����
�|3���?��P�"OR�O�=.����lK	VQ�h P"O>�hU�=,zȬ�
�$~@��6"O�l�嘽AnL�7�y2ؔ@s"OB�ZԦ�?�ڴ���Q�P�pp"O^�҅�0�x�aC透<�=Z�"O��sw ��i����U���r�(B"Ob����"q
�#����>0|�2"OZ0FA��q�
A�6�ЕEG���"O�!b�oOKR@PK�2*�)+�"O��W	Q�ݨ!C$jKi$���`"O:��ULU�XT�����
#>^�%"O@-����/T��ac2��?l��\�5"O4Ż�F�$��m�6�' �L��"O��òe�������J��;����"O*��D��e�-�ǈG�(��|Ra"O8��DaX<^K��/���e"O&+%�7���Em� ��=�w"O�ؓ�
��q�F�X��9�Q"O�=bd��>(�VpH��M�m�\tSG"O�0��N�$���Pq`��}[C"O�	m�Mn����O�^W�%�"O�� 2

�?g��iv�Z�U�@i�"O:�sdI�K�,�xq#J		:��R�"O���E�6b�vYHva�@����4"O(�"I�6.��jå�����"Ov�ӵ�U*B�<�S�C|vR���"OV��'�)@S8)Y��TB�%��"Ox�q"HJ�$A��iCKn�J�"OleRU$;l�0������Z�f���"O��1a���5�PḟID��at"O��b��D0-�E���W'���"O��"d�ȫ9�*("�cڎ' U�u"O��;�I@*<�<J��Ġ	.��Y4"OH�9f@S(���S�a�~�A"OЩ�U&��+Ӡ�p���20�� ��"O� �,j� ��2v4��6e��qI�	 �"O��Z�M)o�|��C�0T1̴�P"OH�Q�П%��i��噰(�z�B�"OT��-ĵL���d����8�"O�䣡jH�`��E,�h�L��"O��-M>I�8Q�'�^(;Z0Q��"O�}*�g����c%ݖZ��E"O��#͉tJF�CE�� <�4"O�ś�ʙ2c����5l���{1"O2p�7���PA�Z'h�Ř�"O
!`����:g�ڬ\�rlK�"O�}�B��R�bAQ�nD�n�L��c"O�`�4�� ���яȠ;Ҁ��"O�Tȑ��<8�dM
��D�4�܊�"O8zs%
P^�Sl+_�}��"Ob�)1��%+�)����t�e)e"O���@6(0���+_$�V���"OfE���N
!<�B�0P~���"O� ��J^0	(��Zn�7M\���U"O� +䅍�Ĝ;�m� NS�|�4"O" i�ղ4���ٔL�۞D�"O~������"0���,��oڞ8��"O(����Q�6T�J\�˘|��"O<�l�4S�j4���)2�� 4"O��1&J*�5)�'�5ab��"OfI����O8fH*S�oR���"OZ��"�]�tJ���u@��23"��"O�������~�J�R6 $�4��"Oj,�/Z�+ � �M-O{vXȲ"O���t� 0㦂�EIڨ��"O�Tⅉ�Z��q���A;qC2"OZl��� �}���gK�$���*�"O��"f/��`ʐ�"���%"O�PS$'Nt&�Ӵ�I1�~Dj%"O�Da�I2�����/D"T�ȍ��"Oh�3�� �s��Y��X�U�z�k�"O���@i�r��d�T"'i�� �"O�APtbD�O+����t��A{g"O��KS@ۿ`�,���L*�b`�@"Oh0�CD�1�ys�!�Gs��I"O:��
�4�
���/^�.f���"O�U"V<L�|�҆��2?O��Ӡ"O�Q�)�:ڢ����J8eF��Z�"Opi�D�B��s�_+VA�鰵"O�8S% 94���ЂO@�=.�$�"OR��^��ʔ��-� )48��"O��I��\�-��}�˗�_��j�"O~���Ł:��qG�/]<�X1"O����>�U�/τFR6X�2"O<���о6���ð$5X��W"O��Å�ϼV)��x�� 3^�^�A'"OXl[&�3 �r�N�C�F�YP"O�cg�F\��-P�̟"oo��PQ"O�ҰM�XY1�-{� ��"OȀ�6m *��!o��Ƭ� "O�=�7N�����2͘�6b��1"O�MʗKT�V�`r����p��mJ�'󠽪!�>EZ\�5Fњ#�z��'醙��T��uH��:A�đƉ;D�,rD��B�5q�H��{��M��:D�(�j��v]�a��kU>��I5,:D��hׯ�e�N8�"���P:��(&F8D�����i����dP�AA<L��7D�hZ�$ۜe�Q��O"�`�+6D�� ���Z/+́S�2�壴"OfX���:^<P��D��jxj�"ONAB��m���s��"b5ժ�"O��5��t���S9�=2�"O����j�*r�-�W��5���"D�@�F%�D���J�&fnI�B�>D���gHV�̀����v���A��(D���b�C��:����]�ɩq 9D������Ke�	�4 Nh[� *D����W�>�@���ܦ8t���(D�0�sB ITh��t�cD���;D�bcLΝaƄ��&'L<T(����*9D�h+���Gj��kr��B+�!yf�$D���&V�+wp�������a�H D�ZrD�Br ���YeFp�$2D���Ə�i
�� /skR�#�;D���2�^o0)��hZ6��7�4D���&�^7b��a���Cf��St�2D�L���YD���1��ӆ���f�-D�l���M%GN���"��)_=�� �''D�x�F+�
�����S��0�"5!%D�([W�ȲX��M��[�\�+ �!D��"�����"�O@2�[�h:D��ER8_+(���C  Kj�q�I6D��bnȩ6�H��e�]�^A�g�'D��,E*g�y����KZLC�F1D����+R,f�t���?Y���XWD1D�@2�ʛM��yq6N���x�J-D�(���
*�Z͉�l)E�(�B�).D��H��P$U�̍�
�0�� 1(+D�ĂqCj� ,�eI�TF���f�(D� ��ܼB�L!�e�:h�~�
Q�$D�p;ր��8j����Dx����$D�pB�T>f��)�G^�"��Ge.D��Eŷ,(8p�P�r�����i-D�ȓ�aM� u�F�V7�z)fL(D��SELpT�R���&+�}8&�L�<q׋L�(�" Ӓm�!LH�P�B��n�<��BI�^F�� %��C؆LxՎ[f�<9"��#gu���N�C{����e�<�1 �'c��j�F�& fļs�o�{�<ɠ%�_}L�a� ���<�bJQ�<yqA��+�e�%
ǐ&�t�gIh�<�'�U/�%R��U�v��L��k�<�DĊ)tPB�^0/�����e�<9�,ر*��p��*F�6}Ga�<9`NR/bθ�U�ݨc4�5{3�q�<AR�K9�>�qA�P&��L�f�d�<)�'L$p��7�W�����4��_�<Q�޶Eq�{`h� q��BQbZv�<1�nɾL�ha��niLv�<��#^S�P,�K�.L_�%�B��p�<��蘷x��)��U��dlyB��T�<� n5,Ĉ�@�%H��kv�Q�<�l�P���!-��Dn�h�1gK�<��*�Y��	� ��Y��k���J�<i�gN8�,�Z�Y)��8���F�<a�J��[7��yYBQ����@�<�撝�N`2�Mդ2��2-@�<y���4aKڼ��� +�`\a�͎x�<���Z+K�
���i���Sk�q�<A'� X2�	���Zc$̐CKi�<��@+,�L��lƘz�\�ڧ�a�<��^�Ce�Co[�-G[�S*�Y�<� �Ģ� ��s�pQR�痺x��a$"O�ܹ�ET�y�B��T��p�"OX��p��)��h[��^d��iZ"O�@�bi�9l���1�F	��d4�0"Op�  [шa���Y�HF��"O�P��H��2�΅P�V���"Oʝ����5B8ٴ+T�u��Q	�"O��KV�ٴ�(,'}��"OR�A�k�%~f.آ���*F4H�"Od���գj�$-�Qf­{�^��"O��X�1��ӃI*���)�8"�!�D�.Ůdjv�G�#TWg<f�!�$^���Yc��%	�[ gß�!�$6'k�X˃(��ɛ撼zs!�
*F�@��ʝ�"�ƭz2#_�|�!�d�9|x�w&�h���jR"ω%�!�Dʁ2e��i��T��M"�`X:�!�dZ2n��B@E,:����ƨ�>|�!�D@�[I,�,Ip()A��6!�D�6KTD���R�-����N-A�!�$�/	�ȡk��͇Y�r���)]�)�!�����R�_� �@�cf�J!�@�g�<�Ig��3'��I�c�R;h�!���8#J�IBÁ����0�m&t�!�V�*\D�w�@�A� u�^�:[!�d޵>�p�]a��sL]� !�duӾ�&GT�V����@`֡"{�B�I�.T�m)��X,����Ѩ:�B�(7*ıɁ<;�1c�L�T8�B�I#!sm�$.�`���4鎻Q�nB�I6��G�H0vGδ�1bG��>B䉠�$\����:?��9[���i��C�	�33�!"��8�q3���>C�I�,T&��"�P1S��@q�&�@��B�	;Y�L��陔t/����J��,�$B�I�!nh�T%[�9L蹀v��uZB�	���L1��[eO�=@!e ��B䉝&�a!VZ�X=�r +x�"C�7w�lUceM	�n�$�p���'�C�	�)?�bV�B�E��J�Q�C�+�h0:�lZ/��A�^�Ly�B�I��t�KD&����3l	v
�B�ZB�|X�N�9���A�KnC��$|xx�(�%��4�ِ�e�&?B�9	?�����f�iB��2��C��"~���%A�X�܀���3�C�	`֚h1ₙ7A�ʰ��I��8B䉫{r���"v˰I7�G�k4hC�	�OB�0�Ќ
??z��ŅP*gO�C�IX��m�g�Q!}�h��k\1"C�	�0F�p�.��62bx�f�?6BC�I�d�M��h�b.Y�C$�C�	u5Bǥ��f>"չ"�'��C�2��<��K!
��$,�H̴C��\��T��4�!z��VB�I�T�^�0��Ő(ى��>:B�	9
F`��ܬ*�8�j��2 sB䉎\����V���k�	S�H7v6B�	'*˲���C7O�,�&�npB��0��i��(�8Z����e�5�:B䉌P�HH�d61.����ϳjS�B�cB���c�D�"�x7(B�`�!���c(	q�Q�T��I��#6�!�D�${6�c!�O1I��aQ聍k�!�� �Mx�슂��9��-�'`����"O0]��,~��)qM�6:��u�"O����9%F�XY��G�7!��I�"O$"4�O,>�a#��.�xq[d"O�D�BN�>���`�Y�\�"Ov�rh��A�n(#��,^�
�"O"�g"X=#�H�	 F� ��-�u"O�*�!Sk
��!B�;=�"�2�"O��J��KK���KAF�v��4�"O�<�r/�0PZ X� #Zk�%:�"O�1��e��Mh�KS/�2g2 e��"O��`��%��Q�VZ�"O�|{���?_�6�.Qqa���q9!�d�l��NL-���&�7!�䖱l���F�.�Pdx��T!�d�U�L3! ����EiI(t4!�=j9�E�s�V�bi�-*D)!��-�D����&�P,�g�D']�!�$V&ȜșEʂ�w��1���>�!�D̘>�Ę�Ӆ�e����؃�!�L��D�m�m�P�`�T�!򄊎7���z3�s���	�LX?�!�$cX���Vn� w!l�L��!��<%�x@R@G@�$>�XeK�*a�!�$�v�N�S��)\���2�?U�!��(5WH䢀��*K�œ��ʢM�!�d�?��a���2s��Ͱ�'�Z!�N�@ �Ȋ��ʿJb�)6'�0'X!� *�ޭa�Ϧ�:�֠�G@!�̆dՈ�ڤ%P�f� @��Y=!�$֧����a��/W�� c��l!��f��d���l)A5���8�y�'��q�&
�q��4ۧ�?n�����'�<�u��KbP$i��"�D�1�'��8 �J'$Ӏ��nK&(J�S�'����6m��p Pn�u9�3	�'��%;q�S
��Es�F�~��B�'��"�� S�e�'��&|\Pp�'0\ĩ�� 7�ZE�7�${�^�	�'P�
��uV���.Q�FD�I��'�6�J4�G	��\�֥��qp<C�'��ӵlӞ/t����J{���p
�'Ǝ�؄.���t@gK&rL���
�'�@��Rm�" �b�R��&:�t�
�'����.����X�g
/����'������C~�U��O�M��'�^4��H�<���9C�ăLLZ��'��1��τwU�b"`�-2��'�n� f�e��q��	)�@8�'uI3�"9}�@����#5O4j�'h�T#s�ʵB�t�Z�)��b
���'fL5)A8�r툓�F�V�v�'4*�sFK,n��Q�W�%UO ���'.�awO;r��,ۦD�0!`���'�n�r@M��������0���P�'J E��l�1q�b�R-|.�`	�'0jp@P�S�:�u�a���bz�(�'PX25� Y��ikҥ�0Woƙ��'�b���&�/%���A��X�T�d���'������D"i��Rᤓ�J��%��'�$d��ߏ	�JA� +�A>Τ�
�'�33�w�ƥ�〡&�R�*�'�<U�倽�<�jw2��q�'|20�t�܇���)B��
�R�3��� PpFG�6� �
q���K�X\�e"O��Ae,e� ��O� ��U�"O�%�s�^�@�h�H MB$&	�g"O"%�7�TO���j��V�l �a0�"O�`#5��.Z898Ջ���I�0"O��K�<�4��̂�t�ਹR"ODبW'�"jX��a�LU�d�|Ղ�"O��ٗlڠmR*�����<�TŃt"OP�(U�ŗX��I��V�!�y��"Od��bb�2Pgb�a��F&�x*E"O�T����@�L�P���P�N`"�"OХ���QMtl����)rH0�{7"Oj���IW��8�@߲J2�P��"OZ��M�`ܠ�S`]�����"O~@��,�D�sG 2rv�A�"Op�ʴ�5�:��@�(q����"Oz�Cw�P�3�P��͌9f��"O�	�W��8F�da�,�O�$��"O�YI#��5t�v��+����'"O�cC��
�d���W9
����"OJY���G�%�~�a�
�ȶո�"O�)`2j�)T�F���k �p�jq6"O��:��\�E,b���I�[[ʰi�"O=�e��:*���/O�/L��P"O&��,ֽ���SnQ�nA�M��"O��s�U����o��:
D�z�"OL��QL �a��4����5P�;F"O�5`��Y�eiH���Y�qa�"O�y�V�qMDa�b���d�z�J3"O\�ʤ���r��}+�@˧	���
!"O�1# ��r�@�ȒJ˚A!�0"OޡR��� ��N����[6"O21�G�.R*�b��T35��%(�"ON��-�#=:�B�g�p��X $"O84��c�^����Fw���"O�qkpÎ�jq�B�&�=W�,�""O�`ѠlJ�KY��Bwe�zjؐc�"Of	�FY<$��CDQ�f^d���"O��b�U6�~���CPl�JQ�"OB��;Gd6􌌅!�Z 9a"O��3�C�dxE,��.���u"OF�2�������2bŋw���"O��3``��Og�iʒAA�v����v"O� ��`Ƕ��1� �΀UT!�"O��Ҍ��$�AK�F�D����"O�<B�eٓ<o�Q��V�b�x}c�"O��"�Gܺ��3��ߐ2�$I� "O������o`��B����g<v�r�"O��h��9آ��$Q9+Q"O��Fσ.+�Py��ʅ��0�b"O�,�g��=3x���?Kl1��"O�aҵԲTZPk+H8!���C"O�%�B�+A�ys�*Z0M�hu�b"O�yh���j옄�S%�Ր"O�t�`�C�R�\�[$��?O"D ��<qp�X'�r�siC�,��! %I
R�<1�³�B�u��o���H�W�<D���u dD(��6. �sC̐i�<	��
#UҔ�%��h��a�0h�c�<�2��89�(��K٭@,6�b0j�z�<�d-Edhvh!��ݯ`e~�J�AI@�<�q@P��h�"�E�H�BFOD�<�w�L�Ȅ PDO��Hyã�~�<�2#�/�p1�2���f�HA�P-w�<� T\R�Ѿ2�tAJq�ȯZ� x�"OJ��3�\8Ef:�hr��I�j��"O~�C��;� )�S͒>j�X�Y�"O����;C�ba�2��.���p�"O~ U�9��������}�04C4"OP��cɾ- ��� xe���"OT��ď޷`��������X��4�"O�M�	G�p��\�4n�?9�h��"Ov( ���0�7͜%.�4�R"O����h\�`�-�1LӞ;�0|�T"O�,����f�9A�;?��t
�"Ov���
�#P0JsGH<Z`h��"Ox��dk��(C�yB훑@q6p3s"O0P[WM=g���3�͌[���"ORM�TY����f��9D��X�"OV|z��˚bf����H>h#e"Of��b#�*���D��|��C"O`����"W�I�vȖ� P��3"O�iy�� �T-h��G;��٩�"O(�*�+�;J�mz��X�6��I�"O8t:��ϞMmHكF�"`��9� "O�\��C�-R�!#�_�V� "O��J�o?D����0��D��"OH�ځGʦ.c��k,E}��T�"O��Ѳ���1��}�٬t/n��7B>D��c�	�P��+T�o���C2D���=C1e�7V��iq�-D���Ҧ� ri�y��D�H�90*?D�8Kǫ;�.�CAD!�~����=D�D0���(�0lI�#<^��n:D�t��ȏc�XQ"���#�|���:D�(����P�ڑ�d�"S���6�<D�\{F9r�̩XTi)H����k;D����!Z�i� �Y"H@�EuFT�"�8D�@�u߃t�b�X��75�,�
�H5D��K�ğ'��$X�G�D��ݱP('D��� &3C.|
�$��K���uB&D���N��H;��p���H��@d�1D��s�GJ�'2�P�V�
w�<x���;D��q�ŉr�~�3�D�L�(8s��;D�|J�-#a(�M�UNА3���"�$D�,�2*֛I8ҵK�(M%#���㔫5D�,c��.\䴣i��B�t%[rm3D�Dr���e�܀`��R�����1T��@P
anV`*U�T-��bOz����RKX�iq���i�92�7D��a%̱)w�B^_Y�+k�*�yB*�8s����F��fp�ɓ-O�y��ԸL9�B��E�b��k# �'�y�#��\Z���ƈ*$0ث5�À�yb���&��d��N54re� �%�ydQe��(�kI�s�j�HhP6�y�,*�� ��Y7zf�$ P͆+�y���kjl�s�3r��۷�H1�y2*�?w��36bc`k7G%�yB��+i�A��ӗ^���VЖ�~��d"ړ-d�٤c�J��a��3��"�_!�S�n}|YA�g�]�tc'�y��O 󓢈��U)��͸n((�"�싀 �8`�'�S��	,�Q�AJ0u�c�n
+v��K��(���ۀ��G��$�Ee] D8���S�	���E��'�h��I8>�Tx��C��L�O<��D���
�)A���P͏%�|��	S�٨OT�dDK�6�Z#;���	1�@�!�� �]�dΟ5���V��,%<�`�i�Oz���X#+�t�"� 9� ���+�!�$�erD����_u�`@0��K�<��'�ў"|�7A>�ʝQ	M���s��	u�<��/P r����fA��3��X�<	��	�6�V( D"���2+m�'��?�:�k�� `"��\wB�K�6D�h˦+ޘO����)�A���nh�4D{����e�<���IH�UCB�J�O�i%!�'y�0�ըތ[R��HX�!�d�?`si���\Bl�X2Ν&�a~�T���3��>�j��s��#��aO?%\���d�RbD����'5$��H99�qOF��D��n�����
��e(�'��O\Rqϓ��?!��/e�2���Rs��Ys�<yp���M0"�
����:H9T��U�<���� �gG#H��Y�'�ўʧٞ�f��-nl9���!P)�ȓF�L��s�X=V"j����f�d��ȓ
��*ulZ�k�QHbnR1:)4h���2	��.ɻ\���#%��/8��=��x���K2PF4%�a��#^@Ň�eM��p3L����5��%V����^��@��8t��q�Bi�FsP)�ȓ%�E���1U}�D񆅑?�Ό�ȓ �:��5�&$���Q*
C���<̌�bÆA
m�$Ya*G�����Iԟ��a�N�*�nQ�D�L=�N�mC�xmZp(<�D��)D�R 虲'�v]�W*Sj�'�x:A����ǅ5_e�=)����y���O%�qc&M,k�H�r�P��Mӟ'�ў�|E�Ռt��Y	4].h�� �F�_�<��O�c�"~�r�[�L�B���	��N���B �]�<a�ȉf�z����@�x�GX�<���J?F.��8ՆK�E���4 �V<q�E�N2еP�B]64�a����At��I�<��.��0�6)A�|�L(S�C!YE�E"�����p�#ї�x���@�d>`UyB�?�hO����@��N!{`��
mr�aݶ{��ߟ��?E�$�DT�(���
<-�,�аhk=���)��l�'X�t�G \� ⧕7UC㓖~�O�!��oʫI�XUA���v�N R�;OD����r`&��?9�R��qJ25�!�D��rĎ�A��:�|�BǇ� 9�ў���(ư(jԦ��i�½:�"�+7�t7�0�S��Mc�*!�xq�5�<dtL��ϙ؟��?q��Ĝ�D��֮6Zt���\=O�Z�'�5D��+� �n�։;v��D,J����O�l�7�D:�S������� �|lΙ� �'|��z�Ż<閍�gښ}���*BaYiI�8�<��y�ҕە̌	IZ$! �q|؅ȓ��(K� �-�&� `%�0���ȓQ�jزv�4S���@��D�c9
���R~��!:@(;dC�5G���b�.�yr@�:����fH�<�%�����'���?�@á_��A� Ac^���'h�(����		���'�L(*�,�G)Y1`�HB�	2v�� �p��yD�W.{$B�I/xXH�+A������L�=$:��|����b�:�����iw�N9�qJB"O���P���e
��eȗ�j�����|r=O���Z9!�a(�B ��TҴ�ΆM81O���m�#�$R�!�b�ۗMŨ9O��G��m��`���Z��h��P��(9'rC�)� P4� �f�e���о{]L�@5"O�x�3�߄��!�ՠ�	6n�Ja"Of�[%�Y;b}K���cX�"O�i�C	�}�P8
C��S�$0[f"O�(��=m�L�r�M(%HN�h�"O�%
�k¹A7����4=<ܽ���ZzH<�R�Y�r;��F�6�P܈e/�c�<AEү`����h�0_\����{8��Gz�Lޫey���EϜp�TY0&��MC�'�R	9b�L�dch�B&J q�Q��O��=E��⅞�*�`��ٚ��w����yR��6H�RU+1�y��E�W�?��'��9ӓ3�a��hޜ�*�V	ӱo�����>ٖ�c�v��a)���hȓG	1h���e"Ob(z$���4nD�і������"O��a�$ s�9�4�\`�T�5�jӌ�=E��d�(R�1KA�L�x������C�!�$M2dD�|���d0�x��M�5��	c��຃@��T[����K��zi���0D��:s�ڱZ\�XZQm�_lN�S�i+D�����L:[$&������Ji�� *Oj�=��O�b�HE�q��"y!+�BV�B��&P�n�sA!ׯ{u���2.N<z"�B��-F��:�DST���t�M�c���Ħ<�H>�*�'��q�l��^���"(/`\�	�'4����W�4h���lIYFC���S�y2�	�-��$h�h�)�KˈY�|����O����'�+���J+��i�Z�4�4D��y���t��E�Q�:Y�P�X��=$��;�,V�s`�|P%Ʌ�6�:1J�#@��M���sӬ�&�S0{��I���j�4d���=}��%K�թ��3kܪ0x1�5)ƦC�	�@�0�mA�a%r�H ��&i�vC�I! ��Z!�M�nV�ªL�J�dC��	1ʤ�$��
K�uPdlH$)�B��92��W�)q�6,�Y`l���.?���$Nڎ�z �� z��AjD՟G{��	0I�v�Y�,�,F�b�gD#z��B�	4/1��k@�2��9�����牿-�~"*�� ��#��jn��ѳ� �yre�*:���
� 8�8t�K��y2���}/�9����3|T�B����y�\2�-�RHY�2�������y"�SS�	p��12nM3�+@��yR�)�'CR2� ?u��CCXh-n ��~ٌ�:��@r-H��B9dH��ȓaN͙3 4<���2�� �ȓh�H�Q�� `UL'Jp0�ȓ6��;�EF575.��A��p��ȓhI�|��&�>@4,TKs)�)@�b���W����#H=4�ԩqC�"g���ȓ?��Y���+)x���p	"0��s����F<Bb�X��i��P�na�Ӯ�8h�@��Co��<X��Eb�\����L�>���ƪ�%�ȓ���ф �<l�0qQ�����R��ȓ*��t���5&?Uu��dЈ�������O�,施�S��+XT�L���,���{t8�ܨ�ʉ�ȓ1����hQf�j���-T".����B�����)*�:�ȣ�ȕ@, �ȓQ����	f+	�3i[�'�6��ȓU�x��cE:R}Z0H��tW����RQR(�cC�'8`f &/�/ƅ��S�? ��!� W��R��!.�}/�-�"Oj���L;A&�C��A+B��5)�"O��b����]"W��"�h�0"O�a��'8;^J����W2H�� &"O^�r�S'�R�k����邓"O��p�	�|i�U�ș�D�p3"O.���p���8s.Ȑ�zԉ�"O���i�n]�!�%KZ�"O P��"H���w�CG��"O�Ly�J&1�
T+a��3.��%�'"OɈ�n�61鼬���0�Z ��"O�\͋�o�x�$ ����;%"O��Qd��Bs��/�w�>̋r"O�mQХ�
��P�d`�1~?�A�"O�ѫ$nJ],1��HY<��"O$�ᕂ�{����Fה&I��f"O��E	�)n8���e�}.~u���'�X`��A��$���Y�MM$}hEE΀?���B�a����#D�Ģr`�*'�>�RfT�*zE��O D�l�������a
��S�5�z�"��!D� � I7�NL��͞*�v2��>D�|Z�зBƔ��	h���pV<D��#�DJp�>܁��98��[��/D�<�Se���4�T�
r��c��0D�� ÈƠzA�(���S4AĈ,�/3D��C挢6(�,��P�a��4�"E'D�@��˗�M4t���i��|-���Gj"D� ��g�&k�$AR�N'5&�|B��/D�`�s���|�[��ӂaIv�as�0D��i��S � ��vJ�6b�\�a��%D�0��G^��Ԡ��o�^LQ��%D�x�� Fp�Y5'��V��D��'D�����Eib4���J�I�Ҧ)D��p��d�$X���٣F��}*��*D���$�
�D �q1�K��MO�E`��(D�0Q�ʈetA@��T�Qj`i��$D��y��O�U8�`2��6Fj�h D�tX���RQco�.QPm2��>D�x�v��'=�DqGkR*�0Un0D�@£`�1�&��Ӵ�<@ۑ$;D�xX���R�!RQ�͗v��y�q�*D��b�`�ɉr��A'D�\�'	�)^�X-xD%��b�)#D�$xF,�J<.����,�p!)�,#D�Ի��Qr�b��D��%�N90 �!D��;�`�(NKp��!��x��Y�%�9D���DA�>���;��Q�	k�)��	5D��X��Ӷ=���� �'2���t�!D�@;s/b'~�Q�iِQ��
&;D���OҰw�ȥX T�Jx��:�O?D�p��E�W >H
��ԵqB�ȩ&)=D��j��<e��-z���t�v��P�&?Q���*�n����q�|�iʻ#I�\�fᓈ3,�}r��	1)�x ��ڇb­)�FG���%{����az�cF�v�9�O��{�^~UFᣀ��?m@@�e�.R��PsoL�+���l��{�cX�:t���eD��;ʓO���5�ա9���i�VZ(!�C �'v���)`�L�M��ʋ$ x����t��s��`��֘�J�C��Bp�#厌�]b�'"���7*=�3�/m�Q2B��$b�C"#�=)��	�P�z@�+ߓ��x��]4��X�퟊5)`j�.ŘU �� � ��A�����:dB102CMr�v��C̃�&<ȱ�uo\��i��'`��p�־ z�'`a�U�ԟx��85�� �"8��􄑎���J�
=��O��(���Z�L�tGX�!�HN<W�tL�	�?�'f��X`XO��ՂO� ��nژi<���H0?��S��M� F��d�K�D3����#k,��" �՞N���'�Rl+��5�3�=ޢ�c�i��Je`�Z�B�����N�HeJ�C��x�cۘ"�,���	$���(�}�>�y�(�8�8��ɢ5���戣y�qQ�C5)�����D�`	�ተ�'׮\sG�B�z�-�'�*�zQ����1�׊ڷ �������_�xl��,֎��O{n�b�AZ�'u�0��k�,�H<q`O�(S<(V!/�'|�%D�M�k��X���,Lm�	�A��P�viY9�Ƞ��O?%��K�P-�D+v�H(]��@s"�([�~	M�0)�&������P��(ps!��#���t�J9.� �ȫ�Y����2R�e16� �?Y���0�hhs�A=����1A L�Q���=�Bi��g�> �!�7AAt%n�S�&�1y����$�0E�" �I�ĊN�3�������i4�i�Ь-�4������k���Ο�	@Gɉ&ic�Ism�$p���d"OV� �����²KB�`��S��+�K�--<�b�L>�U�8e��c�hՖ�R�;5+&D�SF�6jF������0v*��fq��Ce@X(�B���gܓ��,[�Ƙ�;HP9�$�"2��������Ć�x��h�7���i�@�	Mt��w�F��ȓ�B7	:l�4�C2)ʘH0��*���(x��R�
��8sʟ~�$-�V��ͫӁ�:4Nt��"On�zS��)9a�I��*˸@-N%i�S��Iw%+/����MN>���z���a�1"q2ؘ3�'D�8�dA��L�4�����R6����Lf��Daʓؐ9u��I�*��	# ��mv��2I����7� � u8���Q�,@E NDB8륃?	H���_T��&�\?���4�OΜA��4�^<Hs`V�H�t��X�&��������� ���Hʟ�*$��p�֜���A3bNF��"O$1b��N#��Q�UnƊp9�51QJ�!c���Q(��Z�v�X7�]�Q>=1:OR�Q@�7f��ab��r�k�q��  ff�n~�j�D%�i&���ׄ��TgT�j5�F/�4	��H|Gp���P���p����-�z�0��3*؄y���2��OZ�;VAL����Y�oH����̃Z�Vx�e@�|��#���a�v]�E��W��g��8�0?9s�G]45!nV c��
��J�6�jx��O���VAm6ͨ ��'E(��ꠀL��uW�q޽i'�*K;�3� ҫ����e�/�@�^U���<�*�aZ�(˭�F9��KV8� �a�&7���*����-�p����o�m�7�L!/����}�d��yQ`�JC��-.����
��-����`m���6�ԟ�X��I����N�/h��4�0�V��O����@�?rh��y��S�h�6l����.	�܉��D���p�f;G��91��>�-��s�*�sB����	D�I��� s�d"�틎O���8�AM�
6�B��87ܴ���JM��̋��̴(0"�0�J�zB�\���C�j}�ez���rˤ�O�mj���
sϮ���K�<ܢ�OzZ�C��""=�Uj�1C �=�p��(El�$�����b�T�
&�)��� Q`֥��u�T�#)\�=�2[	�cW� {��>E��n��5Ҥ+>,�R,h@P�B�d��O�4ݛRLsӧ��FQh�o]�uB��"^����O^�+�/�l���ӓVxQB���8O�TPGf�9_�d�'��� nLv���>	�a�/t*�"��R�`03"'��E��EzѥԼf\���$�-p�{�A;Y�%q�Í�|�a�R"�xdʤ��}��ޘ7�x9��dO�O�\�ʡ"M�=dp�K�X8<<f}���d��U�|�p#���^�c>-!Q���{
�J ��(^NX�Q�V���ѯ$ҧ����"���K��״|G�)��"��?9�	�#le�������S,�Rp� ߳"���k��K��p�������Oߺ}]�����H�$hb���M�L��D�"���i#"�R�K�Z\�>��G"����4�ݩgF�Z��z��9��bK�*��}��/�ƭ�Ċ7;cn`Z��.2��!@�O�z�d��$�<^��S#3�'/(���FhČh�;G$Z�&�4�E{fˋ}��!z�c��1�&m�s�d��9{�fZ#�jY��@R�>���`�;��s���ŧ	pϠ�x�J�6\9l�*�O��1wL���L�Ճ�<E��M+:ڠ�Xn��*O(lY��8|��MڎF�xd��ĂV؞��e�oF��U%�4]>�e˵�<YĊ��z����W��
�vŰV�VX�p7�U	l��ԋ4Ɣ�(�8���kMta~�f;	�@tS6��*yҒ��n��5X�E@\�4e�<I���Z�,M#@�2�'1��i��B�"6����:8Ӷ\F}"
� �(\:r���.r�<	c��9vT4��͙����r�I��b�Ԙ�O0��R'c�\����s3��Y@!�:���#��G�Y���D�{c4�+O� ��[�H	�y_n 8��e��S`�'����7e�v9�9�퉞6e�p�T�X��t�U��"O��c�X �ҭjy�'I���� �Z���l�,pU�q��+�a1� 3`(� a�C�I�g�~u���/9rt8$��9�� �	Wv�	�2w> ��쒮o41�2<�;
Ҵ@Q��<7_�����(@�z��ȓ�\1��%J�^Шs,���8b��A�T FH�L>�;PX�8�2��>t�(e���"�C��j_X��D��X�|�a)On�B�AW�.B,�"���T�HЅ��-Ut��b`D2)s��X��� \:��I7"6Y�a�7N��D�f��6vt�x�N�O܌�����&�T8EOF0"��x�K�?{�F`CZ0) U�'�ja��*��} ��N�*�i��O+6Z
��'V�9�B��n`ac��b)��b�L͛*�6��'��5)�+��M@z���	~蘸�/O2m8���z/�3b�޴�ȟ��T�вD���q��M�[��"O��B�(�AI`t�0�}[�(!&��-�(���
����3��gܓ1�,���ꈦ'���5χ�_Ԙ��	)3�8���	W���X�Ź_;�$y#�_�kL��	���wLa}rD��A�a��;x[��[���O��3���M�p@����)I$ʰ"�%�|R�c��d=!�B�2��(ҵ�uk �ɇ?NL�I
^JƅQ@
�$�()���)Qs�E�u ƍ)5��hf
P<>9nB�I3Fp�)#��&����G](f�L([d���~�G<i�L-����{��S�o�<���?I�`�3cf���'�b�;sF[^�S�ԣS;m'�xz`��:�z��*ѡ �&3� ���'����@�D��mإJg�H�O�80���<b����?ر����i�q�L#�~Ǌ��[,� ��HD'M��m��/͆�xҪZ���`&N�wK����� Č�g*J<f�<a�đky��(*�����	�2׸����ڼO��L`��?3أ?��'i�4}�b!2}�J�h�O���)��F�AC��%2F�Fk b8"T���0>�Άh:��!)�lP���c.�[y"N��nz�Y�B��jn��1֟ u�M�z�uh�O�8�����D�0s"ĳ%ծL
�'��`��+�2i���g���P�q+ɇi�j|;�f�|� ࡠ4��t���"�� Q���;!`��k�
ׁ�B�0�I�w4`P����kF�TkAL�p�V�`�'F��VPJ�m��3�Ρ*�$
�d\̓uވaX�m�(Q,"<)���:W�쮶[N����3�Q�8;� N�(�B��Uď�k�)[��d�i��lC�ezd�E��?.���PF`�~�.�'�O�ثt�P>��rrgЪ(�~
P�O��4�?�@u�6��U�AS��CtH!��(�j78�O��`b�.,L��SR韅h��IK	�'��-���Ƽ8�*��ʸ�!���lGdث�B��6̓����{ݟ(��Q�ʺ�h�wA���D�ޥx��A����nLP!��W �6k�{����"��
�4�(���F:��w�X8+lXu����b���Y�Σ}������g��1;��"�U��eA��?:}E}��/(EJ�	��ߕ"L���!�0:��
RI�f���" !!�u	"��г��[�&t�'��1IT��:u�vA#�c:5����'ҹ��[��șY5�ԤWƖ4��@:i�����i���D�y�=�%�7vJٚ��<BpM4�$D�H����+4࣊F�V�&=��bC6_�ʜ��!�>�j ie-�-,8x�uM�����U�6�bb���q
&����Ӫ~�腫?�Ot��#�#>�*P�d�D�M�P����_�K~d����O#J��t���M�Si�t�}� ��U��c�pZ��2��kt�ԕ"w�x�K(�~I�UO\�g��4�d�^@:�ɇ&sO�r�dO�O��6�GYŲ��$NI�A���iW�Ӛ��=!KRI�A۲"!y�Vt)��DPyˋ��ub�E��D�Њ�ПT�0d�ӈ+��8Fvݽ����^��Q�қC'B�Y%G'D�@V�Xg����̍D�tH@� jg��e��LE�~T@����gs�]���y��B=[�N��\\�B!�YC�%[�D �`9!�dY���Y!���9���{�D�CIl��#�n��P�?��	8) Z���q�b�V9`�.K��|U8A�S
?m�U��	���@�ާ�I ����d�Έ]!n���kbB�	'RvB�a�'�����a�%dȴ���L=P Pa�y�lO�PRe�=�|R�(@�d�(��|@�)@�6b�C�ɹT�(RBbF$wKx�����U��C��2.�~�:CEQ'o�4������jC�IkI��0݌+�����Ȍ#xLC������s�Z�4}�f/O��B�	�#��8�5�����WÎTDPB�)� �Ѳ��H:
�����Z�{��'"O�E8�i�`-���a�Y�t��'"O渰��	x�Аz��E�<���"O`�J��'No*��Q�o2��V"O��u���`�8UK��ȠA�:HA�"O>$�艖`.��2 $���`]21"OP=�n��rD��݅H��3�"O�!1���Ft�\�P参\;2�Y�"O���4���)V��+)+�% &"O.#Ȑ(�z��b��X6�숳"O�$W�\yh�s��0g"B�Yw"O�ܺ�xt���W�q�8�m�P�<���{;��������QHpA�W�<�J�'�:4��� 8U�.`X��u�<ip�B�`�$�k�?�&I�ǡ�w�<yu�N#ed��ˡ�2"Ӡ�Ҷ��G�<!���^��g)�.X� Eru��V�<A@F̄`@�B dV��^)��Q�<���:#�(y����ZI��t	�R�<�dW�,����զH�sL�5�]B�<y�	)RԞ���~���p�<A,*[h��T�
�k���JD�<�� �&;S&����#j�� Z&��~�<y�ϓ�]�dq��B�%��ĩ��l�<��FH�ƒ���	�)Z`SM�V�<�b�M{}��.ĴP
�#�"�W�<!䢋�:6����&��^��B��QG�<Y�)JvV����I��@(9�G�x�<��@����t*���	T��eje(�x�<��[�.���a� \�|n���y��۾!P��-�}��s���y��9�^1  �$n0��G��yr�ܙB�T�q��!"4E`�!�$�)�&euOװOI�L��eL�V!�D�6]����U)vJ9�L0(�!�$�pctH2�˻t4vLz�-�7�!����歹(]#��R*G�P�!�ĉ�x���� cD(:�� `#�?<D!�$�\� I�씞|�xT�9�!�dA���tff�%�VT�� �W�!�8y�
;� �<)A*DP�Y�2�!�ă�fY�� 0\qDD¹q&!�*H>����+4mk (]/!�D̀6'ڡ(^�h)P(�%*��{�'�0�� ��	(h���g��YC
�'���R ��K�|HCr̅�����'�0�����2[�A��&�J��X��'���'ېب&��/Oa����'�@-#��i �F�7F��'���K�!�s	Dt8�89k� S�'&�yy5	إb<�4�%ߒVT9��'ݜ�A��E���b�c����'nd��̏<O2���L��zH��'��؋BH�2�᠅Fev�{�'8��'�һ3x��6M�*;N�;�'\��"�ji�t�s��P�L��O�t���p=�s)�!_8��w��EF�Ԃ`-�lx�В ��-9���S���D1ƠBdh0bw \j��spa�25	�x�]P悝�" �0���OG�NpFzb��� 4C��Q�'��`�f�I�H���5�9qv]'���u�K;urY��Y|����Ӈ=!�Gl/h�7�ϟxȊP��c�"��)���QaR ���VD��1}N5t�1"�O��B@D�g�I	-?lҴ�N�q ӤF�=���q������5���, 8�:2��}�9����+�8���Ҩ&�f���B��+D��H�� v9˓���p0�� �B�pB���F,7O��P��W�	*O� #�a���h��w�OVS�<9U�I)(b�����y6�l�۲�{s
����e24 �x���'?�z 80b	m�Oj2�Ic(W([�d*��L�f�iz�41l�j��.@`�ҧ����O�K�݂U�H8i���ah������D�>	Q#P�3���'�z`���
-r<�a��.�n���OR|�C	���`��mZ⸋����]��x� E�[�4��N6���>O&|!�Q>�6�s��GL�yY�)4GF$�@�p<9��ɥ�84!��<a��"U�rT�f�E0H�T4A��BW�'�$�u�Q�R<.q��R 4��%��%G�ZN�Ր��M�ɎT��0���,]�?��뀌�@����ԝ4@����O�����
]�H�Y3@�/�~���@�9��A�7�'��M��K?�髃�[t��W�,�p�~&�$�vNo�$�r蚘jP<�5�f�O�e)T�7-rHj�?㟬
�կj!�ƍ�i ��I��aP�B��VB�����U���P�^�bH[f�?����QO�	&z�aD|r��hɈ�O�� E��((�F-8�(����#���E���O�h��M�(Hd`ѣ�=s��y
�'[�3���cg��j��A�U�Vr*O��yB+ 4 -Nb5�)��f��*F��8y���:*����G"OJ5z$�C�4E�VI�!iz�a��"%B�ɵ&
���g\�3�I)[�x�3qK�PM`M���z�����
�X�`�S�'����`AC�C��� �v�S�	|ga~�D�1cfL��!)�'V��eQ�����O��F�Y�Lղ�5�A�����U�(��R�D�<х����U�$�Ih�a���@yB���wu*�����?_a�T��/"Fd�vB�� ���À�y)L�A���(�'Φ3\� �V�Ơ���sy�d*���2��B�g�'��	��T�>H�����C�4-�hzۓ?:�a��&��O�@Yf�U��4���_�.?|dF6YSC@(�<�
��m�,5�HMu�@�KN���=1d F�$]̍Pc�Q)#Ehp`HX)Ah�J���2�W�}bP�"��W�	���<`U*Wg�R���#� ,k�4Q�3Aקv��j5i�>���Od�O�<IΓ�(�pnZ���ʓ p�ȓN4�	5�X(9�����"�}j�D��U����`upA;����&`�,�O���S�X1F�5�C+�	l����	b���r�BZfb*���n^����E�;C�܍x���U�E�q�K]a~"�L�*�e�ǚ9�9KS��Ѹ'�����j�+di�ey��×u4��9eh�Z�d-Kk�,YF�с2k�u�D���O�T��	2��O����H�0k�Q; �[�4I�3W�
� �X3�� *��^1�(���'}b�r��B8D���Q�.��E��'Wt�(��B=�ɧh�������=+���U��%�L���aN�L���̌/[B\MI"(9��ۄ�I2 ���l�	�������z��C 1Q���a(�O9q�!^�c-��k&@_�.���E>-���- .~6��%O�:�^���K�H�j��NO"8\ ���dL=ShBI��@�O��8��y� ��N��$��� �;L��#�f�d��4��0ĝ�C����SΝ0Q\">9s�G̔��H0�S��,����f
0Y)��rNtK`+z��X�@3}���'�|Z�	���84�ǐY�:�'�n����D�r�O?9B��&4d�(h'��&}g�h��O���	�@8�"��'��}�d
 U�=2�jŐo�n��O��+��$�0�:�}��4I��٢4Mۧ	ܙ�'Gۄ`��ql��4�8H��ɚK*`�.\Fp�ϻ:�,�������p��#q0,xa�T"���PG^
>؊��h��h	��	��
ȩ�bϷ!�<�|
�n�8f)�P��_AK*}q$i��� GlD��p��K�"~�I������A�os��K�/J�d�b�$���
��G�����S�O��5[⥄NF0qRc� Rg`���Ox�iK��2�C7���rMM�i�֥0�(����'��
WB��lT��c������T#̬�@�I'ɌP�lr�ӃW�h��IP�XA��o��1�� �6�f���vO�C�]h�Y���(�H���(4��:��4�F�ݷ[�P91b�	�:&���-'6ʸ�|�e�=N(Ѫ�o���j��.<S>�{��-��S��y��J�+T���/ �^�x�r�K?�?9��>K�غN�(���S�K�LLJ�B�Tqb-ԋ8D����:,� P�U&g�a{rG���bH�����C(���Ӧ����út� ��s��d��O����Na����4V���qG�;"$|� ��K�_�p�����~�v��w,-� �U��֍5퀔bb��#d�� ��إ��'f��P"٦(Ij�D��Y UΌ�АM� P���ا�;��O�@Ō��b?�ّ��'w�Uz����kT�\#r@�Ч����y��~�ś�԰���!N��9���П�ybNO$l�KT�]"D����$ݺ�?�"��B��zt.lO�x�T��~���r$T���K%�'�H���P��pmZ�<���$`
}��0�ø\�BC��:{n(҅�c��%Y���dr�v�$�@���:���1�n��7����M3��B�I�V�p$��F�@�j|�ԖU�a{���2=j�'�"~��pe�g�����@CGF�����ȓ_����$�H����(}H�U�ХQ�M�X��ԉKȁ§d�UF{��϶L>������������x���7z��{HЛ$Rt��K�2z7v��g�=e��Yb�'GT�����?[�<Q�wŃ�t�z����dR#8�b��$	����⩟B0H��>^\�U t-D�kخ]��"Ot-8׎'�x@�����Lz�T���a��3t�:��_	�?�(7��?���#�GOG4���2�'D�8Xe���9�L��BN�Ԍ�)���ST���'p@i�lL�E��ϸ' L-�f�h�����]��k��GBc�+�L0*�CCd�-�J)r�@�9��)��#Ӽ7A���$��ġ#������	@ $�џ�;���	[�CƈϦ�tl4�q�m\�#�r{a�:~C䉿�� �W�n�$Q��`O:$�*˓^5�9��)ˁ8�X���$�'o���	`�C��w�џF�����zeh���GXR�d�����
�v=�'F�(o}�D�\��Hh�9���<��}��-Q�ڝ��|�!�Ė<��Y3�E�l+>)����p�0����4�ZP��3�O��9C�ŞP�@��6�ިq$Չ���;�PDC�=�����-нP	��'�Qرӎ1b�ՌT�nM�݅�1�6��/�;�L���$��3��S0z���O�G��O�1�dM�|"X2WK�F%
Yb"O��`#\,+ cB�{)J��dΏw4�I��1'Ea|�թ*�eӆ�?�:H��p=9�ƷFD3��|���e��>=�5'~��1�>D�`�d8�cR%�#<�J�I�3�y�Ɣ�EIڥ1B?)�����$q�'�>z�r�a��<D�HCC���IԅT
����62[�����9}�#�h���d�t
|��`�\�@,i"ƃ�!򤖵l��X��ؤi�鋲 
�T�hQ�`L�sU�Q���'7��CBM)p��rd��z9 i�ϓ z���$
�1,yɜ'���q`
 �x�r풇TX0:�'=r89&�8yG�q�� =p"((bL>a�( ?u(< 2T㇒�����r@�	-U�4#�Ȇ���]�"Ojx�b��B�j$Z�U��)��%�,B�t��>ٴ�Ig���ɘc&���o��9�������wy�B�ɵ*���x�U�w�!��9_\E��H �B�K G]�la{r镉#lvH���_�$�HT��2��<��߾"�Pd���0
�Z7킛d�F� 4��"����I_	] !�N z�br�FY%�� 1�K�/d�''��`��ʶ*h�4��a�Ob��y�.U�:�v鰀A���
�'�&��Զ��ge�+���'E�"!�(��$F��~S��>(��O�L�IE�_�*�aп5�0H��"O���0kU�7����D-U�`2DC���\�x�HEB܆�ɘ�x)�f݄)��C�brp��D�)�J�@CÙg6��Bq�Y�	���X� ƭS&!�$ �C�f��M�#EbD�۠A�O�u3T���G������i^4}��sAT�M ���AP�u�!�D^ -xH ��43t��RZ�V�@�"��^�O?�ɴQ�<��۷a�P�jb�چB��C�ɘ|���Ѝ�����AS9�Ɇo�8�`��'��U�Q��"Zr�D�FI�b�	�'�X)���F�g  ܩ6	Ve���{�'%�!iA@��Tգ2��!v���
��� "�
5�H�R_���Є15�<Is�"O�i�pA� h��c�c��9�z�y�"OF�7C��Kf����+T�e�d`g"OL]S��g��Q��A��U�F! R"OP��0F� 6�ޅxdET#"�z��"O��ۗ�O�-x����cE;i�n��"O�t�I�u�d�k���;b@�{�"O�E�n��vZ����Q2�xp"O�*w�4�Hy*��=Ep�W"O��(�� 	l&xe����!x���"O>-Q� U	>�`���8S�	�v"O�Rw�u�xDXk֪PB��e"O��gf�r�|	zR�4<C.��"O��5��4�2�)a�!BI�p"O��I��V���="��Ũx��8"O��0�FO��P���ӍP`Z�#G"Oм���>#�v�@�S�<Y["OZ(�-�@�Vx����|UC"OvUS�L95轑�JӵS�����"O�9{@'�s�1�r�5�͒�"O�L;�dI��:1�M�X!0@x7"OB��e(�t��٠�LF8&j`jq"O(Ȑ���&�J��mŌ"
��v"O�`:��F�;b���%Ԕ`�"O:qxƦ[4A �i�+�/� 0�'�����[��8�0IB01u6��+�CIL�z�O�/	���GGS��_&0i�OP��İ��H�eV2��*�FC{̓2��"�f{>����T+&N��w�BEe�Rפ<?Q�R ��$�<�}���<��@�S+��L�<�� -��$Z�>`�T����|��ʂ>W�V@3J���0k��-��b����	���ػp�p߮]Wk�~�$���=���0|���2)�jD���C�J\���Aϋ>߬���eퟒ#~��.�m����A�V��'�X̓A�T��7�ZX��?�v�����D&r �J�J�G7�,�OD���ɂ((5�V$��x� ᜠG��A4�(O�>`d/&��]
Q��z+��i�@G�vA$�<E�D�O��ի�d��4I0)��_�v�LUZ���)J
a�TcD%  ��	O!� ey惃%��'�aq����۹?bpZ�W2�V�;RL��o����'���餒���F'�(�����I˹�0�"R)�1-KХ^�U�6m1�ARF��}>B��M�""R,/�b�Y�DY�r��	J��m���2,��Շ�3�j��%A�.*��A�Y
3x�5�O P�ѣ�3g��}�)�Ư��*��	�����Hg�Ak�P?�Dn�͟@2,s~��	X
z����7��r��P��K�5<��	�x�L��?E����H��Ia�%�M�؜�Ŭ���?�Tݔ6Z�OQ?u21��gLތK��(>�~q�$��bj]�>!�'e��:�녩s� :���*x�%X�'.�� #��䩇�O��`i�?k��@��ͩK�4%#��M�&���ۍ4�ܘ�ti���)$�'wE���T�M?�>�Y��(4-y�4w�H���Ǚ�0Jt	���&%�0o:ڧ4��m�2��y���
 !S>#x��H#)��("�h��i�- 0�;��N��?����R�p%�Kj�� �T�K�<Q�Z��J=A���(� ���)�]�<�m��qB���ʙ8nt!k2kW�<�@ن�X�G ��\�R���V�<�W�đ2�l�����YjXA�,g�<Ip���W2t��tR+�<qH_�<��H�E|b�k7 \("�8QbT@P]�<Y�,O�D	�	�]؜b� +��0�ȓ�0�`�[1?l����ϋc�FL��?����N�l�vQ��fٛe�8�ȓ*�!q�AГW���f��r�ҍ���$c�e�3U��D����
+���ȓ&U^� �J�ވ�sJ�;'�ȓC�&`(�N�6	l�s��̶Z�|p��S�? ޠi �Vx0Ѥ�0	�J Q�"O���/ � �2mā�ذ�2"O��b�A��������|�g"O,� �m�'��L;��B�I��aQ$"O~�cjS%	�,��"��%U���˕"OHȰ%
ڪAژM���QVqV��3"OT(i��J<+;��N_��R���"O�:fJX�r��0薭
U�� *�"Ox\�I 	���YABͿzܢ��"O��d�e�� ���(����"O��k�!*�qp#h�l2qX�"O�d�E(�R��%q ��G�d��"O�`1��C���<�t���%K�-��"O%��%c�ds ��\;،R�"O6��� 0��ظ �S�D181�E"O���Bc�8o0���w-ɜ""�Y�"O8�(���
R�$�����
�p'"Ob��CI[�d!��S��8b5��"Ovd��	��JI
h��#\-wl�`�$"Oxr���*����U�TS�HX&"OX�b�`�� L꓋�PJ�#�"O&,��C��EyS�G�+ۨl�"O��!�kC�m�����4��Ay�"O�Pqsa�Yt��	�
�����s"OQ���Mn�6O��4)vo,D�h+lګ�>XA�ݧ_��H�(D�� �+�[,U �HQ/�}�f�&D�����WU��᫆�Y|�J$D��{��L�{d�L#!'G�8�XݰŤ&D��s5��50B�'J�5?�<����&D�lS���-c9�h���:Z��X��"8D�12�\N�$��D��?8�����:D��9`̑�B'�R��E 4h,�*Oj�z�F��&0iE�G�>�8�XA"O�S�,��[t�Q	
�� ��"O�DB��X�d��LЂN��gیu��"OX�0���	
^Qѧk�W� }��"O@�2"��vuJ��F-֘YՒ�"O��c刕b{Z��pe�wԘ\B�"O �R3j_�@�����d�,S�"O*��ehL�9Q�uzcD�t<>���"O���vL �"�b��& ̊p,2�v"O�a{GfO1O,��ʷO�v	Z,y�"O�ò,�G(QQ�.��B�܉��"O����M�"�����E��Di�"O���� N-D�B$��zh��f"O� �7v
�	ݲH�< ��"O�	K��{��τs�:�QC"O2���-��C���q���R$x(jg"O1���L���e�!�"O���T�5s���[��Z=|(���#"O��+V��V�1y�L��<I��"Ob1�`"S�h
�%3.�T"O"�#MD�b��� E݈���"O�̱�g�
��\a#Ɛ�N�"O8'*ϒu&p�a4�QR���@"O(�	�� 9��H��K_��ђ5"O*����0)�,�$)J��!X�"Ozc������ �N�?Vx6`s"Ob�{�G
�8�T0�.M	%\J��t"O�I	��^�	,4a��-�$iCD J5"O����>���"Sl�	nm��"O6�he�ƈ_�0�lR�53@�"Oz�x!�3\��)�쎫&2tq�"O� J�Ru�Pi:@�"�	QF�bT"O0lZ4 B�r�rH(so\*�"�"O�m���:t*ޖ ,���"OT1�X7dL���TL�<����"O��5)ĎT'
!�â+�H���"O�s�����y�T;0��m�w"O�+&����,�'/�67�48
�"O8p�g�5@� c$mɗ
���z�"O�<;�B3w���b�l�#=�t` E"O�q2@�D� I��!�K��j݊"O��*�P��0�I���nR���"O$h��ә�(y�&�jP�x�"OV���W�F�)��)6@9�f"O�ؙʐ�<��mF2Z�"O�XI�L?d�M+tRHb��"O�a�UÏH�
]+��}[�LsW"Of8�)Σ,�|�y���6U���"O(e8V�}�0�c�[�F�Y���K�<�S+U�I����b둋}d�z$IF�<�!�b�j����?zB� 1�Y�<q�iN�Xnpz,R�A�M�#YY�<Y��ʰ|�A��nˠ�& QdCZ_�<����60�$U�M�>��P�g	g�<i$.�6'F����!2���	�d�<Y��a����U:m�A��ċw�<�e�6M�����b�q�<Q��	%��P�tBڌbb<�� B�<�P�F�1?�)pKW:�ȭ"Q��{�<1�'�+/��=p��܆!�d�Hs��K�<�Γ(	�@`q��N��j�q�<I�b%���#e	{֩y� p�<��E��.ڢ�����B�R7
Rj�<�dKU;{�2��P.�!J ��B�Uf�<9@̀j��F �N������x�<Ɂ�!b�RAK����2A*$ 6hp�<Q"Ē2n����=����r�<��֢eu�!3qN*D��@x���m�<�L�{PZE��F){�1�b@�<!T� ���[�.�~�>�b"�Ex�<���V?L��Z6@]#,��aF�PJ�<�'/
!r|PcV�C�s�ҹЦlDO�<Qċ�+�&p	��P�\ʠ�[5��s�<��*��������%Js�<����60���V��S�� +��G�<��7�TT�Q�Z�V(���PE�<����l���Ů�!��1�HL�<�m� x��1(Fub}��E�<���Жu��s��D�hvI	q��H�<���BR�u`!��"$��#$�~�<qs
��2*ax��	\�T!��DO�<�FM63���D�W:���Ȑ�L�<7�� r��԰�f;H��xqAG�<	�ނzf�(�u+wL5 0�G@�<y�-C[�u���¡�F@�!Ûv�<9a�ՠF1z��C�OJuh�X�<�`�?DЈ���}vа�Y(]�ȓZ�EQ����6�����
�'�сgf�N�Ǩ��ș�	�'���CG� �ڃ��	-[h�i�'F�儀�
���b��Z0U�Tp�
�'p��i��:O�p981`/S��m��'0ֹ93��iH�	f��z�DL�'H�M��� n���0(Ҧ\t�5q�'���4%�w�`�AQǒUIE!���  �c�01�^$#4�*�  @"O�h��E��Θ�w�Ii�]cC"O�x`hl��I���d�r�"O�xsC-@�����"n:pf�@m"OR��	T:�H2mUJ�k�"O��:����Vm�}��L��_i���v"Oh4��
����i�j�Up�p�"OX���N�r[�i+�*�����"O��@�i
!$Ϫ�@(��/��L�"O��*�������` �����"O�(H�
�d ���T��SV���"O؝��L�B �	��%V6C��$h�"Oz4j�
Y������Y�p�"&"O������p�S`�<O�(���"O�	s�LG5
�p�H��F�,����"O�颂�Ȯ����2*F<#' c�"O2���ͪ,=����..A�E"O2Dȡ�W����:�ȍ����"O�L��n�0r\�;&Kp��|�"O��ՠ�67����rdܽ��"Oj�m�9�R5Q��X!]]�c"O�����+(�jIY�L�8J�	cP"O��S /H�~*ҩOA��q�"ONՒP�N1�T����**�J�"O��CHǊ��3%��Jz��a"Ob< ���S�4=���O�0hz��p"O@,z�cY#q���;T�}ZĝH�"O�,K���apz �A�	-���"Oԁ:���݌40�_�G6 �e"Ob�G��PQ��
�~��"O�a�0��&)r|x�ńw|̨�G"O�Z�H�LR��k@/�[M�59""O�]���6Z.�
5/Q�̃�"O򄘅圯,��EG�5o���5"Od��⍈O6�G�77�b�"O���5�ٴ]1'V�~�.�y�"OL�32�
�h j�Ƙ�J���R"Ob�x�䂮>/�8z�eF����"O�}�e׺Eq��`T
P�5�xIq�"O�<)Ӯ���z��8����"O�26n�;0�z��P��
=�q�"O�̈�a��#>̈��V�$��U�"OzY9��u����T�v�R"O,�3�@,lz�ha�f̶Zf��c"Ov��'��FsK�D?���"O�,3#�'
�٪�*P0>�"O���%j��#��)Ђ%�ƅXF"O��2��Y(;t<L:R�����p�"OJ(�jąGV\�3*��#P긂a"OJ@��P�y��y(�ǖ�@(��E"O�T���zOt]#���q%ruA#"OR�R'��d��pp�P"Љ9�"O �q��3����4嗚xĐ�c"O�q"��� aQ�x�p�Ć7:�h�"O܌k�
   ��   D  V  �"  "-  �7  |B  �N   Z  Pc  /n  �x  6  ��  �  T�  ��  ݨ  !�  g�  ��  	�  K�  ��  ��  �  T�  ��  ��  $�  e�  �  � , o � y  �& /- �3 �: -G �O V |b Ik ^s �y � � ��  `� u�	����Zv	B�'lj\�0�Hz+��D��f�2T(���OĴ��'L��?Y6�S��?� ��g+�4�tˌ :<��k�!Onٺ#"]�g��9�ud͵<�M�b�%��'p���ϸ�F����
fk5�\� 6��J������ƖH؄���A9}�Ɂa��p�2�;pj �B��Jp��e��5J�Ia�!88�$Q7/
�Y�d�s��'4���䕭
�}`b㈂x�fun�Ŏ���០�	䟴�ɯ#\j��1�M�w��'��<"���*`�&}�I8�MK-O����;F��'"ė9�Pd�beP
5sX��I���b�'B7��O8�D�O��$k���!R=c�2��F)��ӷ"�+c�)k�P�q=�ph��j���'�n��@�U�Eba�b+A�(<:Ce�I�or	(�#X���x��x�}��P�\`�p+3	*7��N3f�{f�(Q,�Ez$݃g&�Av��d�O����O���O�ʧ�y��%#�x�{SCX2X<�$IC��2�?�&�'i�&�d�R�o�ןT+ߴ��#`�i��`���<n&t�0��3�p{�F!U��r�!�>��v������e�A�Y�|��O����.�<0����"�}#S�U���2�,�x��a��7	80hl���M�i��T�{>9J�E�ئ���X�w~t�Y���4���"!�٦�i�k��4y�� �]�7�$�0c�i��с&K���mӲ�mZ�p���?�ls��D<~5���خg��y�s�ʀ�M;��iu$6m�3B���`e�z�>%��O�p�����I�T��J$�F�i	��ے`��/IjH��+ߨJR��oz�M���i���@Ԙ/	� �lߵ�tMK�gS�}{f0�c@�*В��BI,�47��{{�Ɉ�@�=}�)Y�צ5����6�ɿ��L����5}B�9��G:>���p��8>"6��I�d�	�?���FJuxh�/>����$e[���޺T���{��-E�)F{��'�M���ۣI��M$>	1`��m:�a#��{����"O��R3��e�ITƌ�6�)13F�-Hu�vf=;qK3O@&I\�=�Q�ZSd�{2틩�?Y��i����:Ȃ��<C�&<�##�4-�6}	�'���'�'���'92�'Z�iЁK�.�Yd� �!R�2�_|H��s�l��S%�^DhQ�*��[>Μ2�o�Φ���0�M��ː%����'����?U����Tqk�xv	�v/�:};$���QƟt��4A�5�WEưn��y�m%'���)��IT��'n���f@�K�:���m�#L�\�0�O����&w���s���f�Lȳ!o����\w�����O�����f	
B�D�BwM� @b AQ�O��JE�'h�6M�X�O3�ωCݐ���hàS�<��U.�ў��'���'V��S��`�B77�n<x��??ق�=I�.ϛv-i�f����9�'#Q�(렋��&KnZT��90�����'���)��'���'��[�,�@l�%Sv��0�ȟL�ȝ ��P%��Sf'���M󳌚" `ȉ(�p�?QB�7�6H�&��!|�5��3*M��#��ώ]��+6 �
ptL��|RՖxB*�%'@`��*�l��1q�Fw���k�<IT��ʟ��U�L>q�%��
�>����0��y0W��?9�����O��?�'P&�g�pljU8�ƌ�`�����?�p�igl6-%�4�L�	�<�f ��;H¤ss�F9H�M	���e�b�b�T�D�I��h�'c��|r�E�t��q��Ȟn�+�o���b���XODx�B�K!��<iF-�~��� �D�h2�|�UN��Q´Mc����%!�n��)���6mi�0�eO�����2GA7.�rMhB�'F�6�\V�'��O��IM�2#� 8%�LmqV��%A�O��D�OҢ=y�yr.�8+�@���&A/\����"����#؛��h�T���Lʒ]���Ɂra�t`�M�2Z4i���vn��IßX�DП��ҟp #�Mq������7v������-yq(ԮM��0��E�8'y`���sҞ���ǔ��� C�s����D݊0� �5-U>=P,H1.g�'*�<���{��F$j�6�D�/x�<�v�׿kk�2��@�m�$��?)���?	�'x�[	r��&%n��� 8�<0�?!��4�<lڬ���:����P�B�w�ܻè���4��D�;��]�F-�O\�����i��
�1G�n P4a���U�u��(,���'@H�Q�p�x�A�i�Am�@�']����'���.�4B�WnA��O�գq�ȌL�`�÷I(.�:i�ք��3����
������ ����ù~��%
�iתnE�	�r�r��SJ|r���`Ʌ]#&-c��%AwR\�5��'���?1L>I���?-Ov�F�.1��E��R�{;�hIpE�{�'�2��O�6��O6!m��P�V�V�|�VD�mZ&��
��� �MK��?�* ,�P���?����?!���y���`s���� @?c�L�q�)A�Bc$D5i�v,�4"tE�0^>�p�2Q�H����O\�\�f ��(�<R7����)��/���h��F�v�b�+��q��/#bڥ���xޥ�qKY�=��q2���L�:�����R�<����Orc>�$�O���O�3b�T��U��\�����O����O$��/�3}Rh��G>�� ���+��˘y���Iɟ���4�f�'�^7M�O��)��Jʧ��c��Ts�>����8�|�3��:T�AY��?���?�����$�O���
W�^���
̣Y�Y����RY�u;E� ��� �Xy|���(���BęH�� ����3{ ���l�L-� ��:g2���E�O���D �{���H>�'D@\5܉#0C۟)�L<BE��Qi���8��b�����q��� ��8A(E�&7�HpC�'�1O�@ra˛&�d�P�S�g�u��|�Il�4�d�<��%�Ib����xiĢ�7b	�,��	U�A�<@�g��8�ɫ(�J��	���'Jf�!���r����aD*u,�� d�BׯA Z:1�6i��j���؁��D�ȸp��F-3䉓ǯ�L�~-�a3~�"	#�J�d!�ȳ5.Q�9�h�ZC��2*r�;"��k���O|�;e�'����`�c��>V��q��ИK���7mr�'�a|�&۬;�n��1jY�7��x�oN��'�ў�S&�?�bП˜p����!���T�Fӟ��'�����rӀ���ʧ�?�s��
>��
P��1OxR�@V��:�?��g�ʇ�t&�8���9����C�>x����	�C
2a(sEY0d�������q�)S�E��@rV����)�N�v���OZ; {��z��?T���5w ��$˦ ��it>���� ?!� ��]��噑�O��E�dD,K�HV*�6iV��#!�aAў͓�M���i_�xӀ�4�D��B�0_��p��)94Mo�؟��	ş0`��#h������	ǟ@�;'�����
%�P)BE(�8��t�S%[��xxq�8z`�BO�`̧
{��������q��]�IT+Ťj�f�p3,���hL�M"��b��),�42S��4L�1-E �3�wp���A`�$0��}���ǒ�8 �ic�#4�����?��������c+��@c�0�O�/E���	�'�=I�&׵bn��!'�=����+OtDFz�O�BT�ܘ�|��S�����;u@3F���������	�t���O͸1r��D�Qp�ˣ��2;�B!H��P2����׹����X��ҹF~���=;��=��˚H4*�J�e΍X�) ߴ7��iAK>O�tH؂V9���Fz���xǄиg�_:'\6H���j�� ���?ю�;�P�,p�"�ƌO<aIqJ�,�����	T�`���#���/�)q��+=`'�Ԋ�4�?�.O�QjįW\���'����oٖC�#5j�2)��T��'�rk��T���'��i�1�X@K��:
����F2s�f<k �R�8Q�k@�#>�P��J(6���X��$�_�ʀP �L� K�aQ�oƲ�xLn�e�.8�ՊQ�dH4�`�"K��$�+���R�R�q� `�'�4���U�y�v<ن�ݰ ��-�I>A�}���TA(!��y��	�!.�M�?1��4�X�I1 ��ju�D�p����ƹ`m���<�v�I��V�'�rP>���	��<��fݧI�Zur�g�t>�y�g�����I�.��)���$\Z����7bᶡ�Ow��S\K4`�O(�@�=&���$���1�$EHl��Bņ�K���E������zd��eENU:�2�/����
��,xӠ�G���O&�����Q�5Hr���G���B�"OB1(чD�4"\�xLU0�D�����h�X�Z���*ռTk,)o��qavӖ���O���>JD�<�g��Ot��O��DG�ߵB�!3���k�#�'B�8@��1�2�C@J�&�M{�F;#k�m�|�<���	e��|����a�a	5�:�� yE�K�6�����@Y���|�֡$����P*L�-�$�?i�Ol1Z4�'���'Y�O�|��-������O�c�VH{�I#D�{�S�'�8,�GK�9����O0�dM���4�'T�	�$��t�@��EԈyKF�ܽ\���3�B��M{���?������~`Hm�S��)G�RLh@/��/�<iJ�*U�=k"se�˟0��\��ݿCκѢP�	�=q�UR�� u,�q��0��tC�פe�bT��0V�,Q������L�~1�)Ss	6��ߩ~�Lpt*E=jp��u��/t�n�S��'�V6mu�'(�x�Gj�6<_�}��l͌c�~�H2n.|O�b�D��ƀ��,-)��Z!�ӝj��'Wl7m�O0˓����r�i��'=腃� �-�X	#Ɏp��}�'26N"�'Q��w �a�ņY� ��EC Rfh-�F�.=�ЗD�]�&��g[�j�"Q�����.<��4�f��t��xT��P��q,��6��,����M�8��FL���� (%�ɹ���x�.� ��
"����E�ʉ~��B�ɿBd���t��d$�D���E�U�p⟠D{�O� ����%��p%�1?�X�EV3�'���`�!|�t���O��'L�ʄ����J@PF$@2LǞ`���	ud-s��?ID�T�r�%���۲-̒�L�p�P�g �
�����u r�)F��7Q���F�b�I�XpL�t%ɇ��)�D
�B�� J�BA
��Sʍ�?9��
�&hf��b���A�f"?)�-ן��4�䧒�O^���2���qq�O������/O����Z��5X`�BEI��I�@����Pw�ɤe��@�ҪO�'��G{B�'/�7m��]�'��pㇶp��d�@�������1(������?1���?ٔo�p����?����?��w7�I9��(;dL �4�/��"%�Q��)�0�'#���֡��Ϙ'	�bAh� tԘ����;eJ ��Z�$��14�'�p�`	���Ϙ'm�= �cK��@` -�i^M�����(+��'�ў����
8)$Jې6�fţ�N�<Q��AaC(���M*2*(���ß��ɧ�HO�)�O�ʓz�؁�
y���4 >�UP�KK�@�)��?���?鑾���Od擿9�X�˫L����>� x�J��/qn$˕N�7h�Ѕ�I4�� j��ׯޕIItI��N�8}�ܩ���o�&���b�C"��D�o�d�4�ȃl��c&dWLoyht�'����d�4nL  �خr.r���e��rB�{R��s�D(!�րU?��Y�dL-I%�'�*7�)���#��U�O3�dǙ=2��Ac��H2�#��Ek"�'��A��'"�0��3�'�7���1�̠Ee��q@�\?l�(��F,_G��ԦEp�M��C��(O�(H��7O(()��`p��Mbv!F�A}�t#&&D AF��!fܳ˨� �,Ub��G�1��G,UEb�'P�	
#Pj@M=1G6��T%�D�|�O:���՝ �p|8�B4�|h�%n��O��=ͧ0PR6G�h�q �|}���I��?�,O^UJ�ɂ���ퟀ�O���@@�'�.\����;�~Й`��%J0ܠ���'���͆3����a��0�h�#(��h����	�7�LY0�\x �֬u��	,��t N�
���Y���;r�<���oW2����i˔8���8��d�)*2�'��>��0�v$�2�V֠2FKT5
��C�I�"�`���ц1�8Z�M��;� �=��zg��,�ïR*8���䄬~^�p�6���M��?��A~�}� &�?���?���y'�F<m8^T3�V�S˾LS7dؘ'�`�r�%ڴ�wHțv�j\��F�i���<�G�v�������3h$NI�3�2�^�Q�iBL�	3�R�d3�3�	�j��k�L��
�m ���=��B�	7Fm�M�#o
z$���3���V����_�{l��Qb��-9f��7�\�[�.|�Qo^�6(�Iٟ��ӟ�YZw��'g�i��O��2r�Mx�!8!��E] ��Or)S1�ޭp���3�D�5���֩��0�!�ެpHz꒏	�h�a���T�C�')���o�6�(��G/ �"�:#�^�_f!�D�9��$�#�l�@���%c��'|7#�F�F�4�n�ğ���:g�<�F	M|�ųCo	4�V���ǟdr"���h���|*1�K����<�E�U$Dr��jc�Z�y����VJ_l�<� ::3ڑ ��=q�̛��L�'�ܕ��C%��dh���i�b,U��M�kN��B�	��ɡ+�-�Lң� 9����$�ڟ��'
Ќ,r���r��`e�(��3=��lZӟh�I_��*C�]K҅B� ��l膌Iھ�h�/� j4��'�����ۑ6�>�0���\�Ik� I�l��?q�qmZ�;�@REIN"��uP�#?�V��8*�1ڣd[DB�z��Ɉ�(����8��)�/J��mX�n��dZ $C��O�=��	ɾ���^�)§f�����z����d�.}�a�ȓL�$$��D]�A����Ɇ�K|�<G{��'vT"=I�'\�HZ4���$H��" V-A}���'�2�'1<�K5/|���'h�'��N�'����Rd��c��C����(��P� *�����9B]�x���iI"B) ���'Ul�Z�N
�Ā��k�6dN��7Â>g�.y�rk ^����6ǔ)O0�O�h�b�!2�y'%�fB�C��I�d�XA�'N�d+���Ϙ'�vH��ͬ@�X�p�H�}�����'I����Y��|�a��^dDS���?i2�i>�$��HbҰ|=Z$!�I�.M�s$�BͶ�!�ӟ��I����3�u7�'w�?�����
��
P�CX�B*�%z�I�*2���#\�CUPq�����F�+���(On�˲�>>�����$�Z*�`D
(�x��7����aj��Hg���C.Qb�|�åJ4L 6�� n�<l�DqZF�T�EvR���_���f�-:^L����'�L{�A#|O�c�8�fL)AS��Q�,]��,k�k?�D�Ӧ�%���������O`��cb�&z�T)����}~�M���O��Ď'w4�d�O��DɵM�"��%����~�?�޵I�ሦI��]���A�T$���'�����Ԕ5z����ǖU�ڰ¡EQ�(/f��T,�:�]��eX�v)�1�e7u�v}�=�"������4QH���')�İR�Q�q�~�1�U�rגՈ5^���IJy�O�.���!�*R,�:$�S�ؔ���y2�)�ڴ[(F[ƨ;� 1�� ��e���i��I�D/dpp ,S� ��I�T''J���Х�	�2\k�1��eR,XB�'������'^�I� ���	����㢃�7��I'@ފ;��V��"b��4,���/�h���2��J�o���+g���a�����WN�OHoZ ���]��O�Ry���F�sV>u��%[�'-��U�P�r�R-��mфfH쳍�$�>1�iE�7�.�$�+<��	!�e��Y&Y�w�:�����O��D�O��!I�
�����O��D�OL���ء�D�~��ȉRG�P����c�O�� �Do-T!p�3�I����	�O�@Ғ�\�O߰��a�ݫGp��s����΅Ig�F,_���s���;a�۱��|�5ό.E2��{�? $h: ��/f}Ѣ��4{�9Bi`��ї'�T������?���?��Y9V�8�ԇ�MHк�C߶��3�S�O��!`d�H�n�fk�`
"N��`���?�i63�$����<��=Z���I��eK����K2�ƨZ����?����?���[��n�O��$p>Yc`l���� W=y����2�ǈA�LH��d��\��,g\J3@�r��P+	?]E~�
EǑ;���(#��1��<�U��X8ir�Ӵf��Lr�I_��d��4��?��Ǝ�j�`�Ɲ(obQ��
�w�<ِ)Z�>Zb̂UO۬P� Z��k�	�M3L>�B�2_�&�'�RL99%��`1K�9�(4�1�R�'wPH�P�'N"�'$ Ayȍ34�'%���1���Bت袀Ҧ;p�Y��'W>����#�v ��C�f�7M̓��h�5*�:9����RPu5ax�,�?)��h��ɹU�28��M�*g��qCC���b���O���?��q�O�P��F�սV�����D��<6�����C��#Y�x���!���yi��Y�9D�7��<3���=Λ��'KW>Q`��ӟ�9B��%d�z�� 
.�&%��PΟ���%gzp�׮:mJ�Uq�a��W����`&
�K��!�O�%�f�}\�#�� �)z�l[�Ot��csd�u�:Wܬx���a��������I�Iʢ[c�t%b�R�C�\1��&�F��KP�)§Hz�-8��Z�BuV�*��$C�@��&|ب��V-�
'��O��GR� �'TW:�p#�7h"Z��vhA�#%%J�4�?Y��?9��߹@ t@:���?����?i�wx�@�֌e>6m�� ~��"L>�6"�3~Xm�㉒N�ٷF
(:�� Q�)����f�IkjP��46M���c�[�g̓6� �q�	���q��B�h�|r�4x��	�������g�	@}q��O�Z��g�D�anL,������	f�@��p�/Q�4��r&P�{���D��&�'�ɧ���'�I�_�����	��(@��Ɛ	j�L3�m�y��d�������🀲Yw��'�)��g�bhKC X�t���e��+mHբ1*�$kN�"��Qx؞��V��.?���C��>Yw]	sd�� �J�P- !9nT�v�܈��<�E��)lC�Q�fH2�xT�&��4)����I���?�qQ�h��mY��3u`6�z���g�<��	F4J�"G	Z� �EB	�e�-�M�L>QՅ ��S�`�bW�bU��x���{��:F�ğ���	G�&�����ͧJ:t<	�lƷH�R�KP���eF?22��	��o	:��-OPD0� $X��%���)5
:Uo�!&����
7x�@�#���8{6���E�r"�'V�I�c���0��<�&i�e�6ؓO*��d/K6T�KG �-J|�=�O��҂�Or�s�*I�V� y���O#�n9�C�'���$4���ݴ�?y�����'0u����|Q�<�A��DĘ�"F��$�O�x�cA�Y
^X`u$�Jq���G�|ʟ�8J���@j �S�;M�j\����@q���A��M�w%q��@��RV�@%\�X�b,၀��r�����D�O�}�' �iE���8��p��?:~�\@�'�`Y��j,Zi`��[�"� }X����p�O�T�[��SVu�]",�<	�dS��?A���?1�F�>.�����?!��?A�w���'��%�H��+�^ H����M�� q���^��� e��"��O�<��DYy?)TDT!!�RWkU1J���Q�P�qeޑ3$�F����nN��9�O~"޴fV�r�w�̄������� ʜ�p�ѡ����T9-�b�'zў�aQ�E�
i"�,X?H�8�֥�w�<Q�eF��]�'N&�
<�r�py�. ��|����dУZ+��@%]�.Y��:&NC�BC><j��.Y���O����O�宻�?�����LCyF|q�E�_:�m�r#�<Hw&�jAD� ;��FE�P�ʇ�O�y��Ey�CĄ2ߺ\�d�� f}��k�5J|ryb�K&�<i5AU�A�Ċ��i4�͸�2�	����1#ǿf	㱇66�ڡ�Ń�O*���# `N�@��a�, �'�*ӄC䉥s�z�I�WDb~��U��w�F�O�do�q�{�@�N~�$S��J��3�`0�ӎ@�`�'���'���M-<���L4<h6j3l�O��q���;(M��2W��4
��M�'�� ��1mX�qɤ�"/���{�IT�=�(xأi��W_��h��Ű��9��N/ғvy<l�I�|�'Gr�#��V�48������#���cJ>��L�e+��Ӊ)�:�
�I�-2,M�?��4�X)�I��ŁP?�.�1R�+��d�<!�M����?Y�O_"�_�6��|h�B�Ҧ�����]h���?yu���Y�����$�Jx6��vh��%������LӚ5�@����DPR�T�K�`���;j�r��&RJ|C���-Y��o҅�!��A�K~2iߤ�?���h�Z�)� �l;��.;L�Ԯ��,�T��"O�8aɎ(V��͓2.U�a�yѷ��П�I����}�"�OèL��ų%��-0(���
�c!�$�O���O�ʓH6�a���.�ʠ�㠃�l0`�a�x$L�4�'^�؁uƞ���Ϙ'.���1
N���adA<}��< ���`D�@��i`�'/�b>Y ShҺ��$\*1��I�eOې�"��� 4c✟<kE��O���?�~�� ��ջ(�p���NF����'�L�5b��@v� �I+j�j���?���)Z,O\(��#'�
��\����ƞ@e���O��d�O��Ş{n�E 7B� {�ai�l�U�J#��<LȍȔ��.�!��']�F��=�H���IߪP����<�M�B��?��Y���eR]�[�'	�l�A)(YK&�s�A�PΤA�I�)�?���hO8#<Q���,dTLU��,ȿ2��13A�m����<I5-L%?4H�����W�օz$dg��>����<�7��uP�O{��C�E��H��h*�H�C�n�������O��O1(f�<�4���dܯ-�,p���|uQ�LN�%P�%��Mq������q3�l���@*��F�j��D�D�,[x��N�/m� ʐ�
"t퐼Ez�M��?������
G����C��6�vAR����O��'�a|�.X/\H2�EF_�f�P&���'�ў�Ӓ�?aPl��t����#��풆�����'l��i�Z����	�Ob����{A(9���1S�H��Pe�O@����\�Z�Bvl�ld� ���"|Z#�X���dA�Z85���k~��)0Y��'A	e
��zC������)�X�P��uaG)*�L9Rf�#W|�	ST��d�O��}��'�����_�̙#��-Z�,z�'�z)���9G���O�=6~x푋�D�OGz�G�v4Q��nKz=�a�gH�9y�I}y���i�'���'I�I�n��y)�Kʁw��Qb��N!.e�����R�v�A�~`����V�g̓1��p��ɘ�T���2���p�(�G=�^�qƁ�3����P̧�4��[��P�ߢl ZW�̄{Cr���O��
�d�	���G{�OH�OTv,زP�tJ�l�cj�0~�!��Q7�b���Ȅ��,:E��!B���'s�#=�O�)� ��`��8�R�c!���400x���!zϓ�P�ã��&C �1���*��J�]�KL�q�Wa�72x�mZ�ܩX�$�W����O�$�z>�9�#."0V�;��9"擢Mܹ�Q�2-�d1s �M�K
">Ɇ/N !W�i�ߵVb��B�?A�T�6=aJ����={�$3��*�+��E���t�|�׌��)�q ��9� I�%"�Qy��'�a|Z��Qpo�K�lLp���x��	�t��I���`J��t5���oR�xf����?������Xdl���O(tA A�[����@�ׄs�2�c��Otpæn��;��9������|����eB�M��Q+_��D0$DS:�y��9ZR�5�v��s,������;g9�5��pT]�ǫ�a��I�\���O��S��^~���o���A0-B����˳�=�y"��Y8}�򂗷�����hO�4F�4�V� ^z�AuG3֥��W�l�2�'�r#.��!�&�'Wr�''B��ywd�1$��q`Qk�8Br�z�b� X�$�
A��$�L4����G�����?io#�	�4�����w�X�TĈ���+�.�0��A�NRȂh8����\�ʤ`��<'��j���:�Ɋ�>����	v~��?����hO��	=@a9����<^�i��x>�C�I����ެ0�$����(��#���0��4�N�d�<qs
��Q{�5S��R.L���F�P�y~�d`��?����?/O1��ЦM�
���E2F���0�
U!\�p�#\���w��cǂ�����TĹQ��$Y��0+3#�d�z�Í5i&�͢���"{8 l8=���Fz�$���?�B�_�a��z�f�"Ta(LC�����U�'U��k!�9���+�fRF����0<O�#<	A#0����AoO��\\"dMQyb�y���D�<y���o�������' �f��qKS�3�([2�S�V����I�r�.e�����I
(��p��[7�"J�z��Ô���.�R,���T
-�Н�d�[�	B�[�Ir  );�����F�J����a+�pQg�ђj����r�ǫvxi�g&�^����
ɥ	�b����
�O���1擔=,��f��0]�I� ,�+e_,˓�0?��kD*w7�\[6��2xT5���F_�	[���$+�<���F�N<6ё�$�=B,X�`!Xy���o�r�'Q�Y>	�'�Ο��I8:9jY���hFp����@��y������i���*��	9��1����\)��|B����z�`�0�j^�$1ئ���<)��ŦY+B�X]�z�{�.��H��5yA�3��3G�����(D�2t���T$��		��d�O��S�{~
� z�ذ*�)y�Y��V<D�>�*�"O$���Ԍw�`uc���W�<X�q�$�O�Gz�O9tE�" �b~�A!��4g���!��'["�'�P(qg��T�r�'�'����'�0��gX�t��M�/B`TB8-(0��;a\�3�e@��:wJb���e�]+tլ��P��2��,�k�)CW/��#�Sq�>t���[v�X�$�=K�q��Bc8�9�����Q<�+�_T~���?���hO��I�l��@8�hV�mo��0��)q�B㉐Zl<�� �V(���J*X�	�HO�)�O�˓��wER�>��k�Ņ5\l�6�Y}�r�'l��'��)��N
���/�I����,R�1f��Z!���w@m��XT!��`i�-�&G�6������@�b8+��e�O_ކ1`�Ҕ@T�����HOVQ���'U���coǂuN��XD����� ��'bў�E|b�����r�Z�d!���ĭ��<1���M�2����s�V�.5Db�d�P��	��M������J�Tt�!m�ϟ����|B�jQ�W�(�a��l�xKJ�y"�'�"�I�sդ��&�2Gn�A��T�B{���`���z��
@���ŦZ�\G|b�#h�<;7g��(�hd�T�g��rb��:,��N�FuI�,8�ASN������O�.t:�FZ���Y $��#E����'U@l���Z��B�dG�6(�IM>��4�$]�'�f8  @L r$�e��� �a*O��O����Oj��|�ɟFԳ�b�;#hy���?\%�q�v�	
�h��I��M@/R�J�(��D$���$�:#N�'Ԗ!�II��
��F�=�-p@���L=c,6��O��jcJn���gl�Ov�d���dh�H��(�4���(A*ݎ?�<t C�O<F��8l�����ѧƟ��jF���������<E����"� �Cq@���TX��@��?i�l-{�'��O��d�R�${�\J�n��5�$�&��3eP�qV�?�H���O�����O*�	�6���s����y��<Pz(;�P�D���q�f��)�BEG��?��dj�X��]?��I��t��՟���]�dQ���-�P����!��9�?y�%�������2���*�?�-yn�9c��r���4a�|+���?T%��d�^��M�'O�y���?��!�iB���$�OL��?��	�����w�64�p�ԝdئE�s��#���O"��Pĺ����y��R/�d�i��� f-�����C�ϻl]p��e�^�`�b8O�˶�'3r��.��	�O�DP_j�0�aB&Y ���� s�5nZG0�E̓_L���4]؛�O"��Op�c��'ePn��*�C�xD�1]X6���o.@�Ģ<i��O{�f��V��?������*�����څQ�L$x�NW��y"okצq��Ix� 9O�MC������O���Oj˓���F���k��dR$�@�O�V;2���i��'G�'���?����?!��&��ZƧ�9����eN�&'���i�V�X�����ӟ�Iڟ��	8>,t<@���&��M1��!��2�4���?e��1}R�Re��3̈́* %�������:�O�-:ƅ�GMP���$�F�8�;�"O@�!$χ���(�!J�>F�pla�"O��B�nT��jc	�3d�����"Of���*��i�1�B�;���Ӳ"O���`
�@���*�?>���˒"O@��6bV�"�=���Z(]�\!�"O�������m�X�b�	ٯ^�,�y�"O<T�3� R�Xi�HQ��n����ܟ��۟��I��,�'Ӆ	Z�U��
�7C��"Ԛ�4�?���?	���?����?���?!�>fIQDOO�R1�[R�ډ
�>��d�i���'*r�'��'���'#�'��-���Q�h	1v���N�sW�aӼ�D�O|�$�Of�d�O,�d�Of�D�Oj�Pv��?Δ�[0�&FO�t�6G�Ӧ��I��d��ПL�I֟��	��h�	Ɵ�Qb"Χ���ye��@f��YA�&�M���?��?���?����?	��?Qwb�3p��t��J�!x����C�U����'�r�'}�'���'�b�'��Rz�	ț]\d��dՑn�H7-�O��d�O&��O��d�O���O��dM6^B�M8��U	B0#$�ݎ6X(�l������ɟ�������I՟l��ğ��I�	p���Ǯ�tȰt�� {<$�4�?����?)��?���?A��?��Y��|��A׮SK(���(�%u-25����M���?y��?���?��?I��2� 
�� ����gEz�<�V�i*R�'t�'�r�'��'���'0@�2��?N�詳d��@r�#��c�t�d�O����O ���O��D�O���O�t	rP�۔=/)��Q���>6!46�(?Q���� �C�	�c��?�x��&�8~�x�4Yy���<Y��Die���/rf���H��|�L���Țm���nZ)�M;�'��	f�S�:��U�����({3��$z�x���亃�eT7�?�%�
$b�(HpAi���hO��c�v��M�V��JD
	��!H���O.ʓ��c���U�՘'� �����٤zo��8�F�?
ec��m}��y�^AoZ�<�-��ؑD,��r�Z���ߜr�1AvX�lj���)Y$�1�a:?ͧ+X��c��4�yB��FZ���+͊*@��F���d�<���h��d��5��踃@��"S�X�@D�|"Ok�p�h��,ܴ����4/ݵ� "f�LRJ<��Uh�2;k��`ӌ�m�ן���J�;t�@�:��7��6���(N����%;�� �d!]���=����+�S�C�l�%-PXR�q�[{��Ri��!M<��'��>lJc��/0�3/��/�~�Y�!�j}��`Ӣ-m��<A���#�֤R��2M�
1�7Η�;��ABd��	N�	%!���$��
C�p'���'��9��.?�}9C�ЖP�ڠ2��'��'�R�'|"U��zݴnl�	��*&Xݱ%������4��OeD	��d���ėH}��mӾ�m�<`��1PfMҔ��!@� ��k�U鎤9 u�t�f3�9@D*��˓�"�w>�]�V."v!���J3c�"mJ���?����?����?9���ҩ:RbC)/��)r0��x�'#r�'G 6�U�'��D�O��o�P̓���i҅����93o��[�l�����ߦ�{�4�?9����(�U��?qwA�o2�8aC��I��HڂG�P2�S��$;r>a��y��	�d��!�L749^8aa�T���B�	�QаS#ޏ^�,T`�lV	U�!1���4?�̀e*C�~�@)daRa�>+�}नF�d�(����G!����:��r`��5�b�a1��`j�Q"�sN(;�7V@�f� 8�x��e����Q!���tB��`�J��4���Y5#B�E,X���e�xs/�^' $'A�0``����!۪0I4�Fn.|�:e���^��dc�*���f�g/M+L&h��%/D�X�bA�B(��̋�&Mf�XQ/��+�	�υ�ܚ˒儍�J)�������.��2e6�-��7$�͒�,W�_�>X�)љDD@7`�3��uZ�o�(������zm� *Z�sԎ8!#,ړPl�( �b�=���X �;v��T+�(Y�6��uH��wY�4nB*L���ҳ
�Ǧ9���D�i>��(Oȸ�ªO�fR�i�k�m=�����'�2�'����4�p�	P��ɶL �4lK�(�V:���]�&��ߴ�?I���?��+����4��G�``p+ˁ1�.�Y�@�6���֬��d�<aH~��?�0��/r	�űY���H�=��i�r�'}"d�6Op�O�I�O��x���"�'l�Dq��͖2��ʓ���R3�1Ob���O��$	�Z���; ~k3E��MU���O�=� ��p�i>��I՟��'����u�U=k�Fq���G�zw�D�a�'��e�:��'��'bW������r�򭒇M	k��٩S�	2g��1O<���?�K>�+Ox�z���2Dn�SS,ϖCgH�s��oZ1O��$�O��Ħ<�G�H���O�Z�R����㸍������$�O����O,��?A��]���'h	ޅ�U�� ) ���NW-~�'���'z�_�t���Y��'1���8biƐ'
D�1��F��5;��?i������O��N='eq�̨2P-��YUz�zsə�Kuh8��'��'��	��.��N|���y'IX,!��I��E���:�'O�?*O���O$=���l�46�\���	d��Q���L�'qVQx�(y�,�'�?i��1��hꄍ9��I 4f�9�$�Ss �d�O���<v��S�����	:X��(+_� �������Q��@�lԟ���۟H�2���|�t�{����'ϗS����?٧I���O�����1O*��X$L���'���2eJ���w�zInƟ4�I�H)`�Q����|����?�@�����0�+B7sa��]�����O��� 2?1O����O��D�WH��UM��R|�D��H�����O1�Ц1�I蟔����X����	w$I1�I<nf���lS��ʓRxY��?��?	��?�,�L����/`$���FED��E@'+�v���n�ğ|����������	�<����`�B����yE��2��a�p��<q(O��)p��O����O\�d�	���lZ�#��d���BTsS��ord���˟���韬��ȟ@�'���=��$���x]�����&a��Ղ(,���� ��D�	ןԣ hZ��M���?�2�B?�~舰�	�@ql:�"�?����?���D�O�ؤ8���D�OJe����7.����dŤ�A��N�d�O��d�O���A�����I��l���?Ї.GYĈ��,ʷ�:0q��O՟�IGy��'jXD)�O�]��,����V��a��ĞN����������9�b��ܴ�?)���?�'�2�N0��ΜT��2�#Rg�4�-O���JD��D�OF��|zΟh�`�/>:\���� ���a��'�p�+3�u�����O�����v���O���O�I� ��N�Z0c7��G<hQP�b�OƱ&��O2���O�K�:�X�������Vv� :���?�� C�)�&Υl̟�I؟�{a���?��	ܟ��	�<�	�3 �� ��~>.�B�7C�M�	ϟȕ'��05��4�'��4�0���қ2����GM�9�����'wRD�E��6��O����OH��RZ�d2O�%�� �:P^aXF�00h��c��'��T��-�!�yV��������I؟��ɏh��*V�!��l��=�(s��$�M����?!��?V?	�'�� ?0��KZ�@V�@#3<�:I��'���'��'q��'�FǶ4r<7��\������!8,�৊�
)}j�D�O����O����O���?�U��|�� ��8Q���~�i�(U_a��0W�'��'���'��S#{��Q�4�?a���}���571��*���<SC�@���?���?�*O$��5{���+?Yq[:�l�� �3����e�ӟ<��ߟ��	��� ,Y��M����?�����QcТd��SD!(���� �?�������O� �a8�z�$�O��;�<�~(z6��n���1��T�bp`X���O>��O��B��}�������?���矄A�i�Ulx�	�¢W&��V�SYy��'^X8���'m�!_���{�"�2�z�H4$X´���犤�?�K��@�V�'�2�'<��Ot2�'j��AF\�Mz���	I�Q�T"��2��*i��	Iy���4���B�;Il����7.���A�D�1%XmП8�Iџ`E��?�	�0�Iޟ�	l&���NG���)Ţx����p�c���&?]�IΟ���1�R��P>z��,��٘e����	���	ˌ�M���?���?�Y?�̓=]�K�сp^lhTdn���'H&���'N��'�B�'V�T��R lA��Mʦ)��d��F*�� �4�Z�Oʓ�?�-O��OD�n����E��@4x����8XF!;On��O���O<�Ħ<3�L�%��䫓3l��0��%SE@���Y,�?q+O���<y���?1��X_ȁΓ3z&���d��8��
�qȐ����?	G`��?y����28F��&>�H �|����)Y.c��Y0�����	y�I����I$i>��	\~"�H	v�Ȕ�T��IN��!J��?���?�,O���B� {��៬�?	iJT i�dE ��$j��&�`��ԟ�h2�e�D%���=G���V`X)XZXS��< �D�<!��j��Z>�	�?��/O��Hr#�C�|2t���&%�����'6��'�θ�A�'��'�1�|�B�H��#��(��?�,�V�'�ڄ�ҀnӬ���OF������%����# ��jS��8OB{G�6X���	�Q� �p�)§�?q���?eyƤA@H��`J&yAc) $T9�&�'	R�'�HE'��O��$h�l�"�k��@!��=n `��A�OܓO���A3�	�OT���O�1)@�M�F�Ȝc#L�.T�l�	�O���?�T�&���Iڟ�$���W�5YF��hs��X�$�дh�\y�&��yRS�L��˟$?iӴ��l4�( d�L�>��wM�*z�kI<����?qO>���?���^��c�cD|H�t1�hŽ;+p�̓��d�Of���O��Ap����O��I����
���:����>�h+O$���OB�O&���O����O|��bԂjo�a
J߉.:�j��<i��?y����I�$�$>�z��݂�[�")��I�~���IşD%���	ş|�4�s���'ߦ
�Ɠ+_k��3���_��i����?�����'�ҭ%>��I�?EXD��"U��<v@L�.��ԄFc�	П����8L$�	b�?)��S	ʌA�ƒ%�&��Q��O>�BQN�b��i��������9ԩ�f�E��,���B&��'o�� �B�|��t�S���WC�SC�( B-��?�@iK�*6�f�'E��'h�Ԫ&��Ox��
B!����V,���XȪb��O��ʷn�O��O"�?��Ɂ/�N�(0*N5Wc�� "sv\���4�?����?as�͏*_�'���'D�dɗM}�j�'^zǬ8y (� ��|b�B�ر���` 7'Y8�A��J�;zB���R�~-�GMW NކPѳA��,�z8���$w�Bu�KܟH�I�����ş(�DOt�:禖�o�0�+	���
��V��n�Ɵ����?��?��O����I���5����*&��q�'�b'G��p�eF�$ax2D�$j� 8h�����x3#ۦm�!�d��y�@8�%G�u���٣e!�z�`� pKZt��+J�7N.AҰ.B�k8���v'B�a��"f/�
�[FB�2�6X����f��;��D#*��}@��@��޶I�dd�3J�݆8�A��r����ej�,2������2��P�slg`l�H�.�<(I�|ˠk��
�ES�c�͟,��柈�I��u��'���i����[+f��8RL�Fn��4f���j��]!+@)�'.#<O�`���+��#!'Da�����i�� 
v�]�ZP<�HZdx���ʙ�;d�Ys��ջ�xYۥ��~��Y�S(�6�w�t�ľ<����ē�Y�'f�-mb	�&O*.����ȓ�q���եY�`�R�� �!FybO m?�)O���q����ش+z!S���3X������P���b�'C��'�v��P�'[22�jx@c�Z�U$���j�؝�肁�((�҆����%m1<O��x�\�JXu�uK�+���AY�o����c)��Q�$���2<O���3�'6�6͔�PA�T���֌{��(�CT"#^-�$�O\˓�?��J~B�)�"Z�v��Wŗ� ]"Ѱ /�h�'��?9Ha�	V�0�RFK0(V�i��i��7��O��(��L��V?e�	\���T�0Ȁ�+���	l0�1�iѫ,&��a��'��'��k�$T&�L]k䭟�X>��ݫA����l�c�)
,\h�q��x��DL���46����#���p�ȘUG% �e�?Z����@BXp�t�r �H7n���f�$�7n%B�'�>=!&	�0byP��4���b^����Ǔ�x"��[F0��'d�"
��:�����hO��D����Ba��
$�L�w5�X��%�7M�O���O�	գ0,v�D�O���r�� ����
Ç Ĭ0`F�("�te����x�<1�ߟў(���]���[��K�ESh97J���OȵG��O�՘¢]�	K|1�7+֚��QC��^̟,�H>y��>��HO�"��5��H�(X��(��\�<��N�4P�R����R�Tܓq������iH�z��d�7�	�E������	̟,h % ?}�@�	�l��ƟP�_w\����k��P7�R8'l 7(-a4���Y��3�F�b�@
�%�:���Iz��[���*)��Q�0+�n�ⓦ|�4�D��+7� ��x�ME}�-�8/��P8���p�T����� �Mǥ�ʟ���4)��'�'�'x� p���h&>�ʶ��>Ϙ�K���d�;cڵ��I�+E�@lC`�R*GQ��[ݴ�?q-OYU��ʦ!l�!�2́���iB���K?#$����?��E�S���?��:�qG�4H`����.
4�a�$@1X�RD��F��ņHq1�MC8�L*B���2]n�RQ#H7:���͉O*>��^�A�G��uQ�E��S�����0RX#3/�����U�#dTT�@�P/v��9��}y��'��O�O0:�ã��XA}���vJ�h��1$���D���,���p�)fs��B.]�8}���z�.˓��s�W�d�I|��c@)pF�����-"��H��`��88����'��'0�8r�?�87^���(�ƥ~�[wT֐�Ǐ'1s��!��:	��}�+����! �
�X�"L	.��'a	\{5`4+�l���$Z@��=�>�� ���� ش@Q>����}C|�X&��L�f쓗N��v���'�4)����*j�ӣ��w�vt�דG;qOd�)��/jh9qw" ��!WM����4�?����?�'\�n���2�4�?��4*��Y)c�^4���ҵ[��@3�-�*JH����i	�����u:��"v�LaD͉�RV�rS�I
^�s�ֺ�8�x�l�V�H@�ޱ&>��2n�
X�n�N?�S�wD��j���o��q	KL�$,:E$�O��m-�M;���L#}�'��1�^�rTL��nY�))⨒��O���$\�,e������9 l��E%R0$�qO�Ez��O��i|!���^�k�L��D	+$�Bɨ�a�O�`�$	��E����O����OH���?���߹��CŮLB�L��/�J�Z��~}�P�g�A�x���H�b�x�]�H+ �݌iS�����G3�Oab��#*�[s`<)�
K;�u��$Z��i�ㆢ:���
X�^���1�.����ڴ#����'a���M�K<���U&uB�$;E�+H�(Z�C�I�.:�T�2@ē6 2쒵ajE�p�iQ�'^��'�����b���\�$�8թ.�, ��\76D�u�'���'E4
#�'��<������޻ |���G��6J���֣O�(�#Ƭ�do���GY�sΪ��w��&�(O\��6*i@L+X1�j΃w�zY�󋆇XO<M��/5Y�8<�T�˺����ݙ���O�����'�R�i^�����c�Ԕ9l�$mq1f`7�	�"|�'�Q��$��`�L:ua�-���:���0�'��C�ؚ""��s@F�Ay�푱c|�
�į<��Mό��>7-�D�	x�$
�OƘ�GG�RB�?A�?���SD]���Јs��, �J~�'����s"@TZa�gNt��x(O��*���% 10�#R��<����"O��2˚�%�B�����*��1��"OV�2l>JP�,g�_�9�^\�6"OŲ�K�$j0}�a���O���KB"O��9�%� G�ƘZ�φ7�(
�"O�@���1 ����W�c\�Q6"O�A���x�r�0ӭ
3tZ��9"O��$'N5]H����RM$x��"O�������˟�i&*7%D�|��(W+�^,p1U�?0"@��&D��2�վe� P#Kш!�!Q�"D�`j�ۓ�)hP�Z�f��}�t�!D�xP����t�ta��&m�	A��>D�H+1
��%e��PE�j��`#��#D���Ky.�i��R{�d�A�*D��P		/8� Ѳ	��x�	1�(D�<�cCN�	��5c1H@2i ��D(%D�H1F�ZJ�\H�(��R(xa�H"D��Y�A_`:-�g�Y�6��C�!D��/e z���bC��JţU���!���[6$��j �o�XH��
*�!��G�|��5�9D��3d #H!�� j���b��BT)�׭΢J@X�i�"O���нU �U�2�	4V�a@"O\�;u�O���z��F	.���"Or0���#
X�`��)�#:,�X "O�x�"�7f�"%X6y��o�
�!�ŧTND���4@'��Y�I�/�!�H=,e��H�/F Ra3��R3=�!�DP?ܔ��@H� �<X�$�9�!�DC�@	��p��Oq�~��G�ֽ/�!�$�_f�b7D����K�l�5`!��<p�ʧk_;{S���rȐ�kp!�D2@�9ab�?AXm�BM��g!��K�N��x�h�'	<ąr&lP�~�!�D�! cV)��8y'4�wl�r!��=�Ԭ��LK7	�\#'�Ii~!�� ,1SPv�Շ+
�1���f�$�d5Zu���'ضPY�D>��]P�$]\B��
�$L�1��Ľ,����[�y#VA�)����)A�C�I-f�a{��Dʚ��S�@Qq�c��*���n�����%ҧW��6���C.��O����c��r�<�2��:P� �&(F42�l��4A��,��;���b�f�|�|�'���LS�l�~�uk�2w.h5����� ^~�a��M_@�1�&�Њ߮>>Z�*��ԙ}�de��!���͢s���V�@����'J�*�l\:(� ]Xw���T�����3����ЄwrR%]�擔u�"��p#��m}�A� �v�Ν�#�Q>�hԌS�K���� ���#�Dj�*��H %D �����?S�Hl��K�a�h:��^����u.֦M�c�I�L��w�N\�a����H�РNٟA�����d|5j��Z&P|,��܁?p"؊ �̋q8�AC'�!8�1��C�	�δ�C��7|F1�s!܀=t*Ȫ�,�I�)︥�ag��;n�bd�}P#<q1!�+q[�U㏼W~
�8�H��2��8M� ����^�i�	}Ų躣�ʢI�  ���لRזȅ�I�>��%�
��$u*�hC�}�j��[��Ƭ�+�%�&��K�1=��5�P���2ARa��;{�x۳H�_��p�@#�i�
]��X�dC�	�Ss"�R�,Q3p�%�ה�q���C�	k� �TFtM� ��Ux0�B��Q1u
�x�$����qc�P��ҜVG�`�∔��.��DD��1Ȇ!C;6�x� d	G;��x�e��1���3'�	B�x����΄n\�91C*��w	f�X�i��>��TȆ�_��ɢ!��`�
�$[�5T: @,"<YG�HAH1I0.ԽN�Hq��C+rL�|�đ?)
����I&B��Tsl)z�\���ѨU�XZ���d�z��ǬK���)G'8��I��O?"�j���9�|P�3I�R��X��+A"�ѣI��=��u�N�2���6p,�0�CU�)d1Cր�'
�b�H�� 8\)�
��U  +`�_?���]!p\6m0����(�؅��CF��%sӰ,րE"�dt��H�8E�P��w���ے� �x�j�k���J�d1��<�Hʧ��Ze�Y�2�1���A%oׄ+��bQ�W.� ��OV�~]�r��#Kd����7���9Տ,��,�T�H�k�K,8�
ƌ*mg[�J>ʓ��Q�b��N'.�Rv�ިhj!#Q�_�.�]#3ɞ�W�t!�7K+j�&�`��4��u 5�ց~���������a[���M�l��0J��]�>���5�U�J�����Dڨ�CG�U�4�����4�ƥ	D��8?r�9jU��(I�l�Qcm�2Y�t��5+r,(FA�
j� ۵�ް?ua<:�dK�O�����U` 8�� �gA������<E���a��Ƃ6m�1����W�џ�y��F�*��$zD��#/�\a�%�,�0?�DJV>2^M�q�
%��" �N̀�� B֋޸tڀ.�-��6͙�RZ��#�I�YÕ�[!�5��>����X���s�À.1����,�}�'mf9z�OM����
���0B�~����!	~�)(ť��I���
`dR�g�)�'ZUS���IN-K0�C&-b�'e|�E��3N��E�w.)�t��O1�ү�P6�)�^�P��Ǎ�H��y���Ū�H㧦$_&|��r�LQy	Ҏ/�ZQ��▎*����D��$ֶ��u�*MId�k5&�~
��
�-Z,Z}H��$��?Ql���X-#٨ъ��D�NOlȯ;dL�=̻c��\����7:&�|I1�0_*�ȓ /���4���t��0!�fH��{ ��O*:U� '͏�x�)V�? -���TB�&
}��p�k�`G�I�4g"0��DޠV�NLc�F�_^���8����!W�Ĭᠭ>&��B$�a�&e*A�K�{� ِ��P�.K�]a�͓$>�8�wMҍ��O�<2&��:��0��N{����|)%�j���y�e�<x�� `I�wY5��Ѓ�����*J"	�й��s!�q�.��}�:#z����E1
��b���m�J��`W) N ��\����+Ź	,`���D�	��B �Ѭ�y�'T����gE�yT�!G��"�y��� )�T���I�P��M}��1ಁ�Ma>}��!̴_�����_�)�\��f�J�d��k������F>K�Z�S�B۞{�Ќ�@O��p>I#F�=4���A/3� �R����=6� @��ԞY.��GL�Ws�t���I�R�P��A��}��:EN&:9�4�2��!i�J�����-Ġ���. �'Z*Iz�͘�v�h�`%�=��9��&c\܄:#n����H֌
IW�H��*6��Q���H��v�1���ˑ�B)H�b$��l�c�;�4��t���.����������A*N�9(���	�¥��(b�2��`cK(�lB�I.;p>��1�K�~���dlG�l�N���G�^�X"Q��Mě���_p�ţM)�DcQiW�|�̻M�n[�JA,j�9k#)P�ck�e��I�7�<H����� b�O�\�JÆ�?s��Qz�o�&.d�D�T/1aV�K�&�0P� �C�R݁%��K���Sf_K΄ G{"���Wpre�	�#|������ӱ%��+��!]ʤ\p�e�Xa��3A#v�r%�U���"Uɨ5�'���C`'ز�򀳷��)���y��νr�5àNN�|�ְ��h����{�g0
��I�@��0�;���(E'��~̂��%�G�<�0A�ʓ(u���sa�~'�I��\�s�X���M�?RD���;?UEN�yy&�����M�ཱི��Y�RS쬉1ݿ)PIE3y���22LY~�����/�D�PY6��}`5�Сe;JM(��	o�<]�l�<u!i �	��M1rBaa�ُ�O@��+��T/|	5S�c$��zq�|lS�`#��B�;�4 "�U�>�f�]��N	Г�M�IZ�� ֱ^Ϣ ��g S�8�T%��7Xn���'WZ�ub!��뵊��{��#�T-].0!��kJ2Y��a�'��'SV���BS����'N�N�%�캢CG*�f����ĳF*!�D	!5(\�@amU*0wּ�ƊP�t{�@�B��P�nZ�5�P�'2Ft%j3`��Zd̜$޼0��n�0Հ7�^1���Ԍ�;�ay"/�t�c�	Xq-��'m(oJ֤BFO�M�T�a�d�'��>C81
�'K�D��jZ1�ܔ���ξo�8�����8 *�ف��FO����(Ř��	z�<MZ���wKHP󃅎-ڔ��	�M���VE@��Z`S�D�Zf��� �L.h^�hp�%�O���@;��ݦ"ta  ��'Z]���7t��A��"���r�T�IM�%-nEHش8F�וU:�a꤈ ?P��d�]�e&!�$�� !VtY�ܢ&"��3�ĺ+S|��D0��5jB{Ӏ�x7�JZ@@��r�:C@^T#��Yq^���uĄ+f�e�G(4yq��#׌gY�\�˓h���a�O�,Ĥ���M�)�
TR�'N���K.�*�q&A�c��A�@�E�ʠ���̓lHj��X����#�\U(����j�]�r��Q!*�$,=�����yq��1
��6@�K��=3<h�w�Q:��U�B��E�vl��`�<���x���-Mz�j�V����\
��@
�"A.�L;����)�ѠɈ��0*t�
77l��!!���X0�M�B)�P�agޥ;sEC8cb��*�S|�s�%%D��q�%��"��K�q�T�H�䚳IЈ��K�)e��SW�T�UJ�=����-�
��˼r�X�`�$Z2Mʴm���|�Q"��zTp�Xp��w�R���ޕ]9�Bi]��Bӡ�X�l�L�c-S�W)���1eN�	(�=��+ō=�,� eB�X�8��b3i�ў��$&ȒpXa-��a�@Xx�� �	��-2���!Iz(���7QK�i{�A��&�i�DX'gG�M�%jC�CW���@H?iD�iB6D���0?��b�):�Y���0s�Mh���u�I�c�"|� �ܒl�F@��%��nYP�3V�"�)�Q4%xfL^M͠]h�Aϒ6!�$X�9��+�l�������A��`a��:g)l���ɰh�����i��ɳNM�g��:@T9Q�j�TC��R��t��^�S���D$đ0Q�C�,L�>���S�k"KCL 1ce��U�џ�I�������Pq8�8��D2,Ol!�S�M#8�f�)��&?�4����p��R��
��z��}�
����
�\`�"��\�p�� ��ؽ'����Y��ʙ���+ft]�eK7��/=� ,{���0V�<�y�-µqnFC�	9,~�S��B�7����G"�-�������6"dc3O���Mː%�C���$�>mؘ9����-z�u�H�!�O)-�8�@Cr����+����B�!xX(qDW_؞(�1�I)F?n���oD=0&:�B�I6lO���7FD�_�0�B�O����U.����&���>c�1�ȓt�4�e�B�'�t��(a�(�P��I%���+'�)�']�P�z��/>�)�%!�$�х��x�[����Q������Ks!�U�ȓg��\���[�q�f�#G�0�j؇ȓAuh��@�B��p% ;�и��]"��Θ�o.>�j2�nMh`��2	<U���@"xy�80	��DC䉖d&0��S.ח/���	ˇgvC�I�-��p�$�Z�v�bԐwbIm�<B�	!��Y�C�Q�xz�ďW?�C�HA��X7D�	N&���c	*R+�C��%_a�$P' Ƥk!�5����!sfB�)� �@��DG"`�X=QS�
';.໔"O>�1e%	*Jgؽk��	�f�T��"O>QKL����*K�i�̤""O�	���\vt�Axti��?A����"O�	��L&�����B�J`0r�"Ody*�'�Q|�̱��HN��2"OU�!"ܙet��W-W�e��\K�"O���#�M�\��0���� c"Od�U��=m�L����FV͓#"ODq�E ݎL���T�/;��""O�{&L�4y��:��ʹ,ֈ��"O^���l���@0H�	&x*�K"O4��F��.Z]����1�Q5"O"4�
A=;8�X�G�R���4"Oе馮�'Ne�N	r�Pي�"O�I��M�:Q�l=�`��,_��r"O�	H5��(^\Ȥݛ#��(��"O�=��JR43H
թ�D�����"Ov���/�9 }25؇�v�z�"Ozms��Ȁbr���BU pS���!"Ot$�¯��D��E�G*�vL`�"OXY7(��$�l���A�0�*]�"O�d�*�9%��x%ڛPo�QrV"O�	��҉[��}k'Э16|}R�"O���h�<�f�����;28&�f"OVx
�b�"-֤ͪ@�G�a�p�7"O,m��*�"D���R ���`�����"O`mR�F�sfv<���'x����4"OJՈ5�#d
���G�p�P��"O�M�`���M�S(
t �a��"O���
.��qy���;_��*�"OZ��0JT6�nD�Q� ����"Od%
�HX:�#&M�`˰,��"Ox���$y����M��T��X"O
�x�kA5dp�"!	�$�T"OX��6m�("Q���wo;"PU)e"O� F�Xd�ܙ����2}vd1"Ob�*6M���Ġ���R���"O�]�""�(�^�ЗBQ T���2"O*�� ͒��-z���}���Y"O>KG�X�Nl��ۥA��l{L0�"O~U1t+�$��ȋA�wg�-�&"O�|�W�84Θ\���9"O�*��E�挡4l��j}&�:`OXi�<��gL�WA��*p膈VC:Db���S�<���_0@��p+�Y�ά*�U�'~�`�v��G �����^�АR)Oֱy*ٝm?�0Q�%B��4*Op���T��最c͹Nn��'�t4� �Xp̜+FF���л�'�%`�
D�f"�"�g�S�
�'�li��o�3Z�8#��t��"�'��Y��ްx�v��O8����'Z=��K�z�䭚���J���'y���ʇ�Ac���6���M�"O��U-ɫ��Af͞+&��"OЬp� �	�B���� '|  "O�4�P��= �N,�#kB�S_t�!F"O�@�&ҼD��.QV���;�y��$Y+�P���ڡJb��[R�\��y"$æ��5C���B|f�`�A��y���2U{�MjĊ�(:��p�h���y�=C�F�د0���{EY6�y�A�	W����ִ$��4@�ϋ�y2*��t'��b�D�(&���%�2�y
� x��*�4Lp5�T���D��"O��!
�;�2��#,�����q"O�U���k��0LԐoj!��"O�2u��h����FKJ"���"O�L�5�MP�ʕV�by�A"O�\���N���lN��}#!"O�K����ţ�>�:�rW"O^����?Z���� ����)"O�k�A� ���(#��ဃ"O2�h�A�	I�|�ǈ4�*�
'O�M��W-.DJ�X�Y�m��摕=�jCቄ#�ѩ6��(2�r�B���9���d	lz�h!�Aĸzܔ�W�X2�����>D�DpB�M2q��@ ˬuZ�pd)<�$�����<�*���'f�.p؄�S%Aw,�� �L�
��+���"G�3R�и�!�U���N>�1)�,� �}ڔH�Hy�ӎe��u��,���Gܓ�x�ì!�ݨ�g�h�L׽D�$�!s)Яj����:@t6m��|�>D~"���e�񑪞{��]Qvi���p<9��W�:��as�i�d��Ahʒq���+�0]R� 
pL.i\Z����1B��d�iI�U���VS8�H%�آIy�\��qҕB��X&%��j?����k��O�r'IcST�keJ$P�;�'�L��"�ƚrp���(kJ��w�i�h�+�H�>	B�I_�'z�֕��'�l p�c��pvH���H78Hp��'������Y,!��(��	X�A�Ic`�O����J��,�p�v�����"
�(islU�>F)�e�H2Q0�x��ݑ9>��H�!bID������-�Hy)��ܙR�ui���"6�Mئ����ar�M*���� )!�.zK�0"O�"!���c@�Z�`�(U:'!���.|)
�z �PJD��yF
	Y��iEB��VP=��>��	����X�I	���U���Ȉ:ɐ�U⏯�q��OF���'m\mi�g��~吥�I�G�Fl�	�'.��xu *zm;A�[
'D�[�]h}�c�)�MsN<1TMr�|I��";� �	���!C4���O f]V�s$	C�}W:)k�|�t[eƁLU�\려�10慢@��=��8�+��7�5�`�<	���@ޭ!Ҵi�BP�g�ƾ�(Orș@�N!�yV ލ;Fs��L��P�[w�2$�n�&���C�=����w'��i�(���6���怪:G:�*T���P��a�;�a|�ʆ�~NF���	4^)���2���'k�I��lԍ.�A�/O��%�o��t��*n���#$��;<XQVcY�z�J����'O��! (�Lx����M�l�TQ�*Z8A������!���@u��\�4�A��W�Jj�D	#�Cp�*��(�"���3�)S . ��vv���� jƶ��@��`b
�8"ܪW�tI�;��%�F��"@R@�)���ȓh�" H���GA \�?Ab�X�^nL�9�%�*�j�ҭ�y��� `�	�WP�2>�!Ю�+s�Np���Ze�u)��	"�ɡA$V�(	�,�3�N="Ǌ�s.�<Z�b�h�2|����
c�M��[=��"vcO�z �s7��$<���P?B7v��(W��L��K?����OW��2Xt�,�w��>����A%�xR���B��P+�8��(I&)K)yp��u(/(� �!	��D�2����Q�<�����\�X7-h��
��J��!�"(�~�f���$�j��a�D��H�x<���[a����k"I�CB��Ӷ��wl��H|�0�<�sd���?!�l�ddx`�5e�Hy��ߢB}��؆#\)�J���'[p��%��|��):�O�%Ez���_�x����c�t�YP@��tE |�Wm�;~̠u�	_%`�����ov��pÇ	�.u"� d�"��OJ�X��.8d�y�I9<k���Ĩ���`i�O��7!�±������,q/q����'��Q˖���Έ>
��#a�ߨ;��	��y���+N����Q�N�_ȚU٢m>���N�!jTa��%���lҰ�\pP�܆q�CDMP$$y
��kA����`*" �W��(�	:�bZ�>k�kR�،=����ƄY�:
e�'�ɂ�V�*Ҭ�Y�X����t��ɍi0r�9׍W	>0��$Ճn*�R�|aRAX�G]T�I3o��(��??Itk
�\c��z���������k����?y��
�bl�Lxp �K�ֈqBd�>y$�чt	~D�\��(ٱ �pr<��0O�L*֯.��S�D��m,�1�>�����0"�,h�KY��l8�a�O/� '�'�N��H�<3��ō�S�[�:���V�2Ab� MG�'��$��@��RȊ)Ҕ��6(ܮ�#�U�����I�BZ�q��G���H牽f$D�D��xX7d��"��&��\�'T���]��<�6A��9fd�O�=1�ٜAR,l�+�uɖqr�^�H����d��$Y���>�7�d͞g�1�AcS�4�u�GMŊJ��P����^�6�HWE@Ǧ�ZU!0
����� ���Vj	E���2��_/)��rW�
��D�a̓�X)2���p�'\�@������R�jCS_�����t��|��M@�={�CX�>�"��P�4ޒ�'�`p�4�(?F��֝6��yI�ocӞ��OU�L>����&VΉ��;Od��v�0���O.�Q񁊐jj���a��e���r�z}R�7?�v�U��	;��i}<���d���ɹxZh `C��
삐[U)F�Nu,�O��YQ!F���	;R�Vb�'�b�Lm�t��t+����(%J�9�Ҝ�QF׹7���|�D�1�*I�3��xb��=Q>�h!ao���*�(�u6x˓!�f	`v�x�Ʃm���i#eW�,��M��aR�h��A�f�υ.��prF���&B�	�t��E��
���C�t��aJ�&I�l�H���Qxyʟ�$�=�����6O��K7��#J�:w��2vA8d��
O֤��1�̔	e] N���u
W��~b�\hk�Γ8j<aV�����ęQ0�I�tG�}���3K�P����V<bd��P&N,�@1���q|��-ͱ#������8�l̰'�_<c�d�r�	*q8I����,�y"E6,Of�3�(�^����3'�8z����>��o^�1tR6͂�Yf!r����dΟ�I�!�T�����jm��� h]'nT��'���e�>:�P9S��/.�d���o�`�z,P8Q��D�P>��y���)j�ʖ*;�U0�.�%w�a;@B>�O�(h�*DJ�LHT�/k�4���ѽql��8�7��8�m����V�h*1�1}�aZ�9�*�K��	�D`�7��HO`��4�ռҤ���)���PT�P:�R�-�P�c7�P��)� �3� ٦6�AD��"��xr-J�>c�Hس苝A,�Q���A�Qע�7}���������d�?`2���*�x�" ��}�����	�=k�,=�H@@�m�3��yk0�3ۖal)ȈO��I/� �gn�L�"��V˞d #��/���%l �	��#>Y�bɳL���a�a�h�o���y�A��B���Ѯ��1M��z��N�⟼[�f�6Nb� �LP�6��k��%}B����ŊW#]��9dI4<���I�qj�IZ5��/�:-�u
H�[U��*��.U��@H%4XnU�U�\�r[���V�� ��U@��F5��x���AF=��) Q�>�H�$�	j�x0*l�#x�'T��?��"��2��#4�Z�*�� ��=�a~R�g��SG�C�X4  ��:߮k�%S�?1��'��}�B��ń��ː�kD!��-�&��@�)�~�?���'&4�	2ԤI��k�:P�x��q�N��c�@�t7"M���V�i����t�[b��Hs�ء��I�t��(s�+����qd��-��ʓp�!���Q1N���ā17T!��'���Ӧ��G,�HrbԬ�ܻ�b�-ZL��û�d�F�(�"�]8��K�;q���� ��8\lb$�>���������<iR #��>�OP>]肩%�\\(1��(5� �� �'�D@2[c.�B�
�-IΔ�wC �k5r�37�.t/pِ�DY ;�ADy��+�r�13�����E�N�b:0�z��]�uR^���.�x�r���n�矸�r돚ʔ�0��m�����&��=C�0�r��?u��()�i�=[T�'�X�$�<c��x�axb(����@�1�E���M�gSl?�{yb`�(뵀��E���$�,}8>0ۢ�3��:Ul@�[�"�Ѓ��m�XQ2�B@��0<I�h�_WB�F�:%��R��6�zӲ��=1��ZH�\?Ƀ���S��@oܶ%�I�o�8D�p��w�'|�L�0�tX��æ(��iu��!�UR �D8ғMB驠��N박���_�x� �v���+ړn%|q�S,NG�HA�D��$����q�~���!��j`�i��!ݧ1֠���蟘l�~b
/1~���)��*��4��<�y:7�3+����mܹAP L���3C*0�v� 8(XƜ �H��ҧ�Y�<��Ǖj���5C�>94�5U-�IZ��Z����%E�<Zˋ��VOџ�p �4?s���
�xx&�9�nW/GrL@�7�xr$͎�O�y�\��g�R6��!�0 ��3�5lO��	���K¿.n}��R�^�����&�484�Ex������G=�j����O�`ͣ�*˾6�ቐA؈G6N$j��� �9�Td�sǗx�"	��֩�󤉌k���_�@��Z��E����P`~��V}Z�i&�ʆ��� ���a1� � s���r�=����'���D䍷7p�ɛ�'^�pQ�'g���>1#��3=�"�C�c�9�����3s"�=ѧ$4�]���o�n��ҮI?�18��YJ�0�d
��0��k�m��W�����g� K``���O��m�C�
���B�*_�V 0�p�(�O�Ab��Iިe�V#�:)�)[d�P�قvV�D��+�<9P<O�X�m[O���p���n�?͡uj��T0.M�!��Vڀd�UN)�'�(H��^�� j�X&e��Ӧ
0�(���H��|ѵտ]��7�6e�ܠ0�'[P��BɆ��)�v�tO�8Kr��ܑ����8sq�O�-�螄4%��@ȉ�+��$���=��V���,���N�p�4�� O>$�%ڒ	�(�� h7�ʌ��Ih/pI�F�V '�d)�c��o}BD��
�($r�'�1Oh��� ��c�`բ��*��i���Ǩ1�O�0h��)i�"�h�͇4eh�8��I\ؕ�<9��9�I9Z��76e���@ˀ�&�paa�dW�et�y�K
^nQ��j�6V�v��UN׼';�q���p�-ѣH���:�Hc�W�W|^��	{̓�^��}
���å��t�x$�<�e��#f���cW�q7��6IX?5㗟^;��$_�y��ɰb�X�Gy�Ȱbrb�"e�T>|���b���yq�)"/�H��	�[�6�2�lZ=-����W.�iy���qg�#I���=���)���Î� .�P���0|� ��S��n����˞dH�T��U!���� ��Eo~x�=A���B?qW�[�4a�+`>���		�����/`��p��oډ: F'O~ q�H�#$�F���C�t�I�QD��u�U��>tbqo�
T.��'.�ܢ��;�V�p��9Hw�$�|:�5+�K	�6�v%�ń۳Rۘ}��I̸<)���'<��4a��\�9�bB$����C�-!g0�Y��A5���p>�`�@F_�f���f��z��V�'�@�FɎ�r�)
�X3k��	��S�f����ݛ�$Ʒ �0!��T�<��Bӯ,R��B�׳nŔ����S?��b4
>�t)�Dſ$l�Dc��S�5ۺuc%��fs"iZꑷ��B�	HVb��"���c2�h;֎��?s���ش��DV���!ܴyÉ��'�1���3`g%[ 9��M��'{�px#��5h���&c��+֥
�'�]�&�I	T�'ㅺ"�L\K�'��%�A%A�h*���^:��(	�'!|��k�-�1 �˔46���'*��Ca]~���-5fȴ��'�F��6�]��Y"�� !9p\��'f� :�L̍HC�U"�a|�)�'�x#�S�Y�&!�sK�j���*�'�������+�8����[TL�c�'	��
6@�Ϡ��Rk�*Q�zDx�'zDL¥�Qb�\�Rg1H����'��-��.�=���1���1U��4#�'*��+�ㆾWzI��E����'_��"�Oo9p��� �6fHP�'� �1ehZ�N� 4Ѱb���R�'����4�×��4�W�[��ݛ	�'� �8�M�~����1Vm��'ܘ��rN� &�,�*�hZ��L�C�'�����
]�Lxб�-��!c��y�'d`y ��A'�l��2���(�'MLM�"㌠8s�
EE�B��=��'���+��,EHC0�mz�'���׬�b�z��CY����'t��bXqxx@Q�]9k�n���':$`i��=D-*��!�bٌl#�'iJ3�Eە䴩����JW؍��'��(�g"�1"LvȂ7!�S�����'�:$�xFT4��!�c*���'���jSD�6�vA����a��z�'w�h�����a��dD&���'[`q1e�I�{pZ C��;T>X�@�'��@�µ%�)رϑE�VH��'R(���D0A� ]�I�;�
aX�'� ���ղV�7���|�z�!�'����fB�\������~��]��'v�=
e��o^��f*߉3&I��'�)�PS��E9�O�H��#�'Җ��v��`4�����\l��x�'�b��s��(e�<�tm2e����'Y��[Ł����bEV^zZ�h�'�.��oW�J�L��E�=X!���'y8]�Rd�k,XU��B��s�'�}�R�Y4��ŭ�?�Z(y�'K&����G�b4BQb=Ⱥ��'��zWb_�>�� ��!������� ��9��]V4ta�`c�x8��"O~a��"��M�Rh[C�Y+z{��y�"O�e��C�,yތ���֔Q�N8Z�"O8Y��?7/�(��#E:�� �"O�H+���,%:h@q"حMc�,�"O�p��-]�wt51c! �B��"O@\bW���zm�EJ+�4n�Jۣ"O41�僛0Y=�0pI�:��[w"O�!00�S�l�y��ҪO���"O�����g/� �{ʢ]��"O��q��[8 ��A)�w�x��@"Oj)Zg��)9ɐ��f� 7�Z��0"O��I�׹?���Q !-=����"O��
*��X���82��I�"O^Q���oFl���/$G��P�"O<�(�oX�j0&�P��۩"�:5��"OJ�x����f��a�,@�6���;�"Oz��AN#X�`���^�A�ĒG"O`͊��	�|nĘ�$�X�.�U��"OBͨ$F[-r���y�c�L�v���"O�Q��l��-�@�&2��"OԔ���C�Y��0!�7�nD[U"O�DQ�������-͑9����1"O 䱰`EM^֝z�l� ����A"O�����f��(2�kX-_�,1�3"Oh-��nņ;R�aq@�beԴaf"Oz�CI��|2���b!)md�9p�"O>��U��f.�%*3�]�5L����"O��)I��<�b�2�%dkX�s"O�q�ǁܐ�J�r1f�+G�L�[�"O�xkF��[���A5Ń��@r�"O�aA#�~���d���0
!"O^a	edU=F�
х�H�Z"����"O\��
+*Qڕ앗�L5��"O�t��������Y�'�ځ�a"O��Eh
;�|�G�P��4�"O�1���G2W. hi�GJ�-��-+�"OT ��J�/^1�Kk��["O��Q�
o��˦��"�`��B"O������5I
�c��Z�z<D"O"ȊQc�O `Й`�Ԏj
Ty��"OZ��Ui �P�\I&�*\�9s"O�x�@BIF8 �ԵU$(97"O�pS�$��u�f<�À�&���7D���S���\Ѥ"�WC,[c�3D���`�_�lw��i�BG�jL���0�<D���B�˺@��1�!�"��e�s�<)t�$6Wd5Ke 1'Bd;���u�<� ��;$�=��N�>'�,�ڄ r�<��� D̎H2$W�U�j�<��y"��`w��t��ԙ�k�i�<酂c ,�U�X0�*��&Sf�<�Q JH}ڠ���	T��Z�<)�M� #���	�zJ^Mƍ�Z�<��N�|��m�GN�v��O�Y?Q���S�P�n�a���8n蘒�JM��jB�I�w&D��
IA�3) #�ZO���dɁ	��!"�ӥ0�JD�׬>!�ĉ�/��Ŋc'^ �)��+�I!�$���8�[�fR<(�`�g)�F!�D��>��bԁ ./��̛ 
��e�!�Đ�d �r%R�i���+cIK�JE!�dN�^/.��JU)RL1�-v�!��|s�@I&�J�P����a��a��B�)� ���R��ID�@�a����Q��"O`,�fJYO_D�cj���}H�"O�AP��͑ �F	J�8��iIA"O�j��Ap�n}(����^��@z�"O��z��	�^��;�`��:���f"O�@����7i�>d���=v�Љp"O�p�\7N
��
!�ՁnH	C�"O����'X#F��U)B+B�A��͠�"O�4z׭�@��x��)�%s����"Oi��nE@���!���Q�>��U"O��@��
w��PE`�E鄬j "O���Poy��!�dNS�6��XCw"OB�ۃnw:<P�0n�[�D���"O�T�LC
PA����M.WL�D"O�a'ǔ�d�4%�G�Qd�5 �"O��K�o
�}@�6�+4����3D���)�4.�b� �/�(|�����4D�p�କ�>|H��E�]����4j/D��� ̒=$��e�(7���B��+D���f�AJL)��Fڈ!�F��k(D��idb"4x�a[pمH��ˀ�;D�p�q�ģMȾ=�a�W}�()��6D�Q󡉷n���H���RTn��!��&:�P�J���-&��(�K�vG!��%�r�(���l�0h�dI62!��D
G�Ĉ0�g�/���q�Y<n!��ƨ=?9Ѱ�<�Ȥ5���O!�ΰ]�"�����<�Ra�!oܰP�!���W�>Ī��Js�X�E�7�!��8x��z��t�"H�g��0�!�đ��Rqq�/��X
�$ӡ0!�
w^�AqG"	}E&�0B�f!��>J(�pȖ��-E�U�5�2 !�[
:���IۜE:Nأ0�B�c�!�$�d��}�,�D+2�S7@��!�d��m�m�g�c��9a�U�#�!�,\�LJ4ÒA$8)gU�I�!�dL�]����u�쐳����'&B�C��YL��1��|u��B�'3b�@B@�aE�l���\7J��-Z�'�����
8�J2VHO�u�����',�((�B�#iS� �Z�H�Z
�'��Z%�g���c�$�t1�'�JW,�'gஉC�.k�T��'~��ueU	IN���n�w�>��'���(���K��l�W!�%w�Ѝ�'�!��kRs�� �7NӔp���R�'|�tx ���||�$dS�`���
�'?�ZC&_(~Q�1T*׳S�5i
�'�D�@"CZ��Η2SW �	�'���hE%��\��0S"��+F��P	�''���B��Ur�������j�>|��'��`��쎂Xz4@��An�Ta��'-���f�ȍJE�	�w��x��-��'���	s��9d��q��K�0����'�|��F��	B(���n��h>���'�*��D�ڶFq�|`�o�Q.����'��jp��:��A
�G(��:�'Y�����&+���'B�H��q��U*������|ɀ="q#޹i�(�ȓl�Ĥr�k�LL�Q	7�M9~:���E�|a��E6��|*�
�7B�����D�dp&�!t���G>�䍆ȓ&(^�1M���h��F[�e���S�? �����}#^I(��NO����"OրX�Oװx��C�M�N�|h �"Op,�aL���D�T.]� [�"O����n��b�� ���LI��Q�"Ot���/���u�W1|ɢ"O���AaW¼@�) 	w�SP"O��L��%�Lك��N�p|X�"O���O��zX�!f�29�r�`E"OxQ&�[��-�"H�NÈl!w"Oz�����/��7��K�.�t"O�Dx )�6O���3F��2��v"O�p�HE7�8���X�H�2J�"Ox:�������̜;E����"O��;Ҥ��4p:���l�R�䲡"O���% ޓr�\D���
'�z��"O�����" K��7kB�ك"O���p��+v� s��#SyvaC6"O� 	4��Ml(��j�� Y����"O,\��A�>`���x ӚtF����"O�x��V����I��+t`��"OZ8ۡ���+�2����R�}��"O�	Y���dḇ�Ό8�L�W"O
�Aq面'N�p���}�J4��"O~��E��9szЀU ��`wah�"ONq���-k
���`K=(�ޡ�&"O"�bV����M��NU�i�l��B"O^p��*@��(�*9Q���"O�K�e�(p�vm�,��Mٔ"O`Ԑ4A�=��jt
B2^�p�1"OԐu�20e〯��D��"OH`:ԩC��ȰS�+@�W��av"OԑA3&���*��Š�jR��9t"Oj0��
�����J�>����"OV�BUFߓi}6���蓁K�X�0�"O�� f���~TL��G*e~H�G"O,����ßx, i��ס?Z���7"OpP���Z퀁zQ�A�K7�pp�"O��	D��!EZ1�̉�!+6	��"O �Ic�J�bLM�����U"OL(��KͽH߬T��싯/�*+�"ODT�A�\V�"䈄%��f����"O-��j��qt����z�b1"O�R� 'R���뱣ܯde`|�g"O�����B1�~ѻ`CҀeH�� E"Op�b��X�+qTm�����X���b"OJ�:4$�m|����ݥo���Sf"O�<��η-�T��e	ìR�fE��"Ov`S˟4L;�@����5sx��"O���D].Awr|Y�I��9�&(+�"O��P�4*�t�� )Q-Dئ�:E"O�����W4>��#p��0M��q�A"O�-ҧl�/	�x\uZ�P-J�"Ofɩ�z]��t�+�Ҕa�"O�Թ���.�ֹ*�`�iF�lB�"O��6�7KI��(��D�e�}0u"O<ha C� ������=V��+�"O,��2/�<5+��"kđ�6u�!"O H3u� W���Cj�-V�(��"OB8��@V\���B�� ��}��"Oz�+�,�5���c��<\���*4"O�\C��a��A�w��Hi4-yd"O I2��BP��r�`F�Zb���"O�!�gj���8��l�
>8`:�"O�zb��$�6}��+�H*�Mp"O� F�;Qm�!+�I��	��H;�"O%h1bQ
B�:I��dY�G"O
8Y��
� Y���~�<���"Ot���q�*x��+�� ����"O(H��5i�����w��h�"OhP��(G�3Ӳ�q�蟤8�:9B"O&�"��C/B�nܛ������Ñ"OR�B��h���(�ھ���g"O��` [8��=�U�D�P�Ӷ"O���Ab����Cf��m�r�"O�e��ՔN���*��*[��k&"O�Q*�!^~ϲ�b��=uPND3G"OZ5�H �]�ځ� ��/<�@٣"Oر8H��2�E�Ʀ�+ ����0"O211���v��1��'�6����w"O��!R	����E�M��i�"O��	�GŔ?�2���K Ȯm�"O�rD@Y�D!����.\�t�"Oj�IE�Y���pȄ��� �z�a�"O���a��Q>&Dz��p�B!�R"OF5����15�lqT�B:)�P͙�"O&M�#
$w��Ÿ!#��8 �@"Ob�Ѳ��}_�ЀL��{z���"Oڵ��h��X��;���q��H�"OL	�&)
H�0MJG��8B����"O89���#�شi2�0'��Tp�'���Y�?+�乓�3S@��!�'����${#D(K���Q�9r�'��"��K�)��5�$�A�)i�'��큢I��GE>�Wg 	Ok`5��'�����@�*@;�V0MR��"	�'�*x��٢^���T�� B��\��'��!QF�F H����k�2j~Y!�'zYkeݗ@[�ۆl�z7����'9��wǊ/z$x�����r�]z�'���M_��	ydl�<���0�yB���@h*��Q���3����yrM��=VM�m�7�:�l��y2Ń�l�Г@艥7�h�k�ô�yr���B�x�Q�jU4�$�{EG�6�y��ҖoY�Li�Z�+��1S	I-�y��0Q�]��U���cO֩�y�H��
��!�/5s�	Bsg��y��¥T�PdY�آ/�6��WW�yB*��*������	sǢ(iPm_��y�T�8	�l'i�D���ƈ�yr���j=:F`�_��`hthɶ49��.x!'��"F��Ô�;8@!�D��������  芘LO!�
VD�Z$��u����F-�V�!��V�GL a����!L��!��K&L��� DY�@z��FK��
�!��J_�#5�F�}Z��S��$g�!�$�d=P�����qE��"�&Yv��I`��H�����X@@��Ė'V����"O�{%�F�;�� �t�NAdʀ"Oڈ*@���._f@{s��Z1�Űf*O`]�ŔY�Z���M����TZ�'��5���c7B��6��Py���'�8�W�ن^��&�� � 
�'�j%�j��+!���C�Ԥ+	�'��)��@�D�y��X09L�S�'�������4xЬM��o�(�Ƭ��'w�ay�e�7�� !�!��'N 5X��� �Y���p�6�����m߂-r`"O$�Մ��`�z8׍*H�h�v"O�� qIX7+�iK1혲Be�A"O4\���P�,x�t��>6��@�"O�@BER$j&�i�J��a�Ĕ)�"O�5�3�.]���($IM?+�VA�D"O�|i��Ⱥw��Ia���N�@��A"O�<*���s]�pБF�t��0s"O:| L�5�~R�"���*�"O����)>Q���@�f�6��6"Ox�x�/�t�I�F
�3�Έa"O���"��2C����ك��T�u"O>�ȧ
��$�*A�p�v�Yه"O��I�m7v�.��a#^Z<�w"OZ�Z��#8�ȼpF�B�mS"O"$���ˀb�bH9`L�$zPb7"O��Bq�Yw ��@�9}�>�p�"O�i��'T�@��a��C%�u�d"O�0���"���ؑ����<QT"OLQ�\4�����Ć`�H�*�"O��΋t��Q�ƋT�W��!�"O���sBAdtк����[�(�2"O��#%읐QT�@�J�]���S"O�y8oK�s�0����R�9��a�"O���mD6|��uNַj�8�"OΉ��mŗ��4�&��y.�S`"O|ˆ5S��M��NI-tk�=kd"O�x�uOO4�b-��>95���"ODݠȇ9"}Dd�U#��*�0j "OFL�5̉$|��kWc�Z��d�SOD,i�#͢k�5�'��
^� �8 �?D� *�"��{[v@�-9���A�=D�8�0)N�Q����!�@�v��Mգ?D���3�M?G��3��=A1�Ay7A>}�`c���O�)����܆< W�D�`-����'BZ���b>=��	�c�9p�'4�UIl��L�����U�]�N���''��"TK�z�٩�Gܾ�K�'�F����	Is��SQ�ܹsk��R�'H����-#^X,��@IW�x�&|(�'Ơ�aUʒW�=�֮�l^:L�
�'�\l�s햤c�2�g$���yB�Rmq�lx���b��A �
;�y"hĻz`*�RpFEL�b��y���r^"�
��Ԝܪ,�5#���yr덋Y�y���C�"G��P!��y���I�~���ۣ
0jp*V�ܶ�y�LA�$��|��)� ��,�,���yb�5(����A�|���9�$V��y�n�9I��W���_YlQ�g�yB�ƴo�p��&�Y8)� ����y�aF,V|�;�j]�N�ɉ��	�y2�ɤbdp%2��\��#AF��y�/˂��51խB����j�y�&Z�YX��;��4��Т͈��y2��5b����Þ�#�P�1E �y"��:f#�: W+	z��ѭ��yb&,�dL���}N��M�'Qў���L��`ֺ'VTC�ä4Qj��q"O�]�&nw��{w ;aZ���"OdA��-æn� �[�/��])���"O��fD�%�<�[�� Z���"OJ|rT��1>M@��x�h�g��S���)-p=$������L����Gb O�!�� 2Ȋ�G@u�����:T�!�f"Ot����1'ڔс!�E��<p�"O�y0a��8�ba�i� �J\�S"O�!�ic��ճ��\�~���q"Oȁ��l�D������4I	��IHX�艑��;�6�"�a��K�40�� D���Oȼ.���2�eV�P�5҂*3D�K��ވC�艣`C���by�$*3D�P�u�O��ہ\	|6�Bs&D�rS�A4E�1ِd[�C��``Sm#}B�)�S<�zA�3��g��њ��Q�<C��	B^�Cf4Z�zu�U��dG0#<ϓVQz�bq}f\��LH��d�%�ae�<P��O�Vr̅ȓ:b�a�� P]6}���׎n˦�ȓe�n���$�D�b�bG\�<�A�ȓ5$^�K �r~*���"��fD�a��-��%kf�v�b\��#U�q�ʥ��@z&Lq�`�A�R�Y��>M��ȓk�4�#��MP���7\	���ȓ_5>U�4%8y4:\�N�$n��ȓo�<)���B�1�#k2����"uSA��%C��i�AnG�b��`���>��,��R��?#ͨ� � D�XJT��J70Jы�h��:p�<D��ّ
גo8�� Ga���f<D�\$
�|Qn	�Q�TSj�Y��-D��i��O�.��9��(}�H-k�>D��qq$��l'�a
S�͆\q
))�K2D��BAo�"S�%)ƪAM���ǎ1D���F�mq�y�rK�(b^n����.D��JH��d'�ت�"ސ�"q���.D�x� �ǉ7�� �1ɜ�T����/D���*^�R���3ֈ�-;�,2��.D���╽+�lų���&U�f�3��?D�BW%Z�-y~YqB疒F�6��ш:D����H�<fW��z7lQ)k�&���7D��U�Ц@��-�,8��f�m�<����
'4���)Z�,m�,K4�Xh�<��iѴ7��h!���i���sʄg�<���)Q�9Eg�<MY��g��w�<A��X�=��w��5�(�yƇ�t�<�p`�vZ"�
KU0bq
���h�<�6��xP�"g/���y��g�<A�Ñ����2M	)u����cf�<�q�Q�Ȁi�mI!� �� �	H�<���C�>�,JpgM0�H����X�<�W C�qh�Yad�n%Z1K&�X�<q�L��]���5_%T#�AQ�<�u�\A��%W�M�.���N�<	f$rEx�8�&�!`�C��I�<��G�n�
]+$�Ǜ7�4�K�N^F�<Q�*�{(r��Cn#�A��(��<13b�="O�uqh�9 ϕ3Rq
�ȓt>�-��k[)8|	���HM��ȓb��m�2C��<����ͯc�,��`�41 F�C ���r�U^��ȓ!gF=�c
;;	-z��V�K4�Y�ȓ�V2��^����B�֩�F�ȓ���2�j�]�\��'�0�P@�[�<�HPO��(F/�.!D��o|�<�rBM���+�ロXD�M�B�<Q�.�B va	%*�,m���hѨ�}�<�	\�W(�}���E�;��p �os�<� iq�Iþ|��
��Vg�Z9��h1��#�Yx����9�: �ȓs�@�RP$��lݬ��V�<d4�ȓLĂX��DA�^@���RV~U�ȓ%�&e�+^�~�ؕ���)cq����`�̊��@�4���H�.*�N)��7�n���C yH�@"C�'9�l��Mm�)��`�7���`���s��ȓ<,����*�,\�1�����@f��ȓ9CreGF �>THҍ'�FЅȓ}b��Q�Nԋ?h�Z���)Vх�%Ob��D�L,T�hPu��:�	�Ǎ�3F�0�
�f_���؄�!�z=�1��8��M�&�9�J��ȓme	�r�v�~�c��';Bj��ȓ�Di��&��Yo"��B��N�LY�ȓ=��9�
^�F�9�f���6}�ȓm� p�g")$����K�-[p��ȓ8�J]��AQy��w��,l�ȓQ%R�i6�͇~��2Ƥ
02����j:�@�R��A�z�@	ũ>��5�� ���Z�,[�2̹9�jX�Qy���D�phvg��t;0�0s-�"g���ȓG�<��2�t���(�M�n�.}�������$�Ό�Ŋ��H �ȓ}4鸂��)h�p��@�*m4$��Z��R��ԾL�P`�jA�Bp4I��V��V�(KJ�p��U4#�9 �"O��I���f�܉aT/`FW �y�L��ȱdc5��eΌ��yr���h���&M4�Dy�c��y"��S���*�둻G����s
Q��y��U%7.�iw�@?0�s����y�f�!`�^�Cd���:G��B����y��X�9ޭؓh	�C�8���J�	�yR!�w��@r�i�h'Zu�F�
�yr�Ul��(��ǜU���;��/�yB��X�P!���U�:!�Q��7�y�a��V��y�P�	�I�v	1��y�-�|���
�&ל=L���j��yb��4��9+��K,^je��)�,�y�oϷA��I�ET�(���+�yR ��b~��3
$3�����+K:�yҮ��h�:43�`C+(b���D��yb`�
�>�@ǆȬ�
�`�����y�eX�EcP��=$x1`�����yriL�5�Ѐ�1
�(Ȭ!R ���yr�z��0��L#���+��y��φB�.Y�&��A���!ب�y��Ω�H3E���5�K\��y�/Ɓ�S-*	�0[&����y�ꔠ>t�S)�#Qw,˄����yR���H�\����Y;:ߨ|�j�2�y�O�R�@�JŢ-'��c3�۬�yR+�)m\M�0��T&�=
��O��y�$ =(n(�H�@@�#��y���&=�ij3��u�iz��H1�y�!�]A�U��J�?P>���-ѫ�y�7��б��ˎ~������y��7g�l�"�"\����ZE�I�y�D�]к�p2����ES��š�yB,��,�,�#Ԫҗ}.D�t#Ι�y���)Z*����@�BF��$��4�yh�Dn�up &�:4f�	�#�
��y
� �8�Ş�#���ZQ�%,r�5"OH|;���%-����EF]�1�"O��i7Õ�z� ���d׏Tg�<Ó"O��R�*��_�"i���EUR���"OD����ѽzE�L���C�pW�D��"O�����;s&�tB�!Br͉P"Od I��_Pjp0qk�'`�mjG"Of傶g[M�Έ��L�)A��"OQ�$ЕzS(��F!}_l�s�"OY��E+F��� %�"=Ըk�"OD��#�^;1�Q���K�!f �"O ��ƥV�Ƥ�"�43P!�"O�u�-Mc<�e�̭$hXу�"O�5�� _"��i*djN	R�*�R�"OB�q�%�B4Z!R�[�$�"x�3"Opd!@�aq����[8-�.��!"O��X��Z�h@C��ę8��th4"O�Tq%�U�?'�]���ky0r�"Ox�KֹY�X!�7���Va�k�"OV,��,L!�R��!!�'t���"O`�+�q�Ti@1��+���U"O �q��8{C�I��Ԙ1��xP"O���&��6Jj. cs	��|��"ODY����$X=
�GU3krx`�`"O�y�������ȼm4���"O:��S�17��сp��,/}�銴"Oz�q��G3@gz={�	�c�"O�������H�ay'�ÝZR�5	�*O��I%�M�*��YAn^��|ѳ	�'U�azwE͈v HЊ�I�-#�rA 
�'Q��t�Ǿ,s`��DDN�#g2�k�'�	j�!մA7�q`�O\�"��)�'g�5bF�&D���DIfԝ`�'K>a�ӭ��E�dI���$��p�'���z�)���X�F���g��'=���!U5�TQ�6�G3HLv���'�`����~�>�F��?C�L4��'�Rě����u�)5a_,>���'��H����TU���(Ӥ!V��b�'6�d���V�"��i5�]?oиJ�''�hUہ��T�۽'ή�B�'��4#s�M�o\!B�!����'Lt} 6,�i�����@ETpAS�'#�y��`�%qI����9��k�'���R�J	w~����kїal�m�
�'�(��"_�;��Y�`���*����'5d]�7#U�O~IP㗂M5�`�'(H�qC�� S�`X2v�a*�'��%8󨍫dsN8��MF�d�:a��'<ځ3cT&V� ��14)�4"�'c>q���	��PY۱�9&�p�Y�'�р�E�7�h\��ק5�f]��'B��#��&`��@��
B����'���6�1dc� �b��J� 	�'K�l04��>p����ЌC��A`�'���T�[�\l�t���� '.@ �'Daڤ�![T��Y���%%P�)�'a��b�(�l�!ʄ#܀q��
�'i�Ԫ�E��X%X��K\.���P	�'Hne��F5a��-�C�C�	���Z�'�ɂP���բTQ 12,3	�'�Fq���6G�����9i�J��'��͈���9Y��+g)&Pct�
�'-~�Ya�ބx��%H��@�@p������ <թ��R�S>,|:S���uI�a8�"O����9C�`��ْa��ʶ"O��S1$ xQA�it�	�"O8�!焛>`�0q��.kV��`$"O���U�������*/#>��3"O��I�K��[X4!2�X�� U"�"O�5ͨ@��H�.C4Jo�Х"O�T֡�!9�LbsRz�3"O���DʝY�� R`ì^cꜣ�"O�ؓ�=G��3�/k�1R�"O<�sG�%��EZ���~6n��"O�"��?N{d��.E<("O�QXЦg �\���H"!�W"O6�!'��Cp�!D��d�$�"O� B2� N�\�CE5!�����"O�qp3! �[<�}�Ta�|�� rR"OZ��r�®B.�sN�;tA��"O��ÂZ�*cË��$�Ò@�Y�<��fͬ��X��� N\xs ]�<�g�7X.l�EC�2Ecq��Y�<!��4Y֬qd��%1�j�ˊW�<1�&B�s=��wR3W�b͙&�U�<���"C��Y�`��8a:�iq�*T�ĸৄ�)%����P;(�P!�*O�Yt��n����ӵiE�mXd"O�	vK��"Z0��G' ];���"O�, ����\��8:��݈Z1:�2"O�i����<{!�T�5ą=uJd�z`"O6Y�!�0Ķ��!EH�N4��B"Oj�2� &Bȁ��nK/)�b,0"O�Zb-_�-��;��	#]�PT�"O�@�A�o�t���+��v��ò"O����� ���24KG��̓&"OF	�Ǟ�:=X�� �x����3"O¬�&i+�5ksi�R���1"OT�Sԫ~�΀q��R=U%@T�<��ᖊEc��aBV�xa!���j�<i�cV�֦ȫe�J �rJ^d�<	���3bF![BE&xF� 2�`�ȓKp��jA8i�b� �fυ]��ȓ6w��t�VG�V#҄Is����C�ZM�ʀ) $�]�1��B$JH���Lx��X#�d$(3!�1[�T����Фڶ�[Z��$��M,Q��E�ȓ
�����;���B<d,�� �����̿7�-:�`�=�2 ��UaL������f'�U*`��^8��ȓ:^���C��UU&�� E�s�DQ��2-N��a*V�J?�$�2�	.lX��z��U��k��5B��g��9�ȓ��y���P<Z�af_��Մ�Z�ͻ@i>gj�P�e�={�B��ȓ��|��o�H�jq;��K�~D��@E���$��q/�Xk���;�6���0	�q���pp�P[,W�n͆����f�T'v�:��9Ać���yBgS�vH�i���)ȮXV��yZ(��.T&�&]#3���f�)��'������,5�왢��?[��C
�'V|�t��O��պ�EJ�RV��r	�'_<-� ��)���H�P�t���'�0��+�$�(�
�@���	�'b��*�$_��H,H�#,3ɨ��
�'A����W>�,9�"��u�� ���� ҄���:n S֩լ	�a(�"O>�Ӳ�?=�90c)۪B�X�Yq"O���5�E�
 �t���c�"O"y� �ǤJT�Ec�?a�J)��"O,@i��a��EJ��p�����"O2�lX:Y���*V�ez4c"O����&R �P�(H��	�P"OF���KO{��S6��$/�p�pC"O�YX�lH`�2]0�#�(
�����"O�>;����Sm��18�'�EE!�$ё*蚔���ȥI�%ù4�!�d&Lҹ�2�Q�=Y`���.�!�� �|�]���
+2S,Yc#��o|!��4%��Q�K�Pp��5�Ƀ]!��O�&Ϯs�#�~��A�T�$<!�ZX*FmA&�;Ler�⃤��-!�Q�Z�d�S��&FK��X�T�q%!����"e�^eY�eQQ���!��O �=��B=	<�ee���!�շ:Ö$���a&񱇤X�%H!�$�&�ơ�­I#k �\���ڿe)!�M�oh�[��	}Fȡ�Ǽ;!���Q�HL�R����Qiڂl!��|_�,c�͋{�|i5��	!��I�b��-r@l��m7¬C�o��)�!��Q�a��ui`��+-|�QŬɯ2�!�d�>l���2da���U��
�7!��Y�
?�1&�V������=!�d���\	�E��z���2g^�E�!��dU�@�6��$f���ͅ 	x!�$��7�L�`A��/�
�	���'d!�$�LW�� gM��$��QBM�4K!�,rGj�$�Y�zT��鑡�%h!�ˆZJ�zp�@�Hq�lI��,2T!�Ă�qX����A�|�i6f�<,!�]�a.��@D>Q��ܳ�j|!�ĉ.Z�B��G��6z���vOC�,!��X
b���E��_[�Q��,(�!�ҋUd�!�d�,Q�����m�!�d��2�4`��ǀ?4K��r�o�$K!���J� �"W�3�
X��k .,!��,Sy����˓#l�lUqaIHY!�$�0#�!�k��?�QR���-}�!�Ĉ�� A�9l�0ѢчS�rL!�<V�� 0i]�Hu���i	j!���RJЩ*�':t�0q��+^E!�R�:x���)`;��`��V>�!�L���yb���- �C.!��$���y4O��T���O�O!��4Ю4��C��]�,m�P�c!�D��<t��N+�V�3� U�!�d��$�0`� �:d���E91!�DԔB�Ը��L�}\�7fP�uJ!�d�3k^���D��&qr~�sg��08!�d9w�"'O*&Z��+�Ȣ/!��O���qQ�J�C�aJ�)�%BG!�$�o{��T�0��E��h�Q5!��ϓ���AG�^*�P���%�=>�!�$B�:�,m��k����G!�č�d����`Y)TV8�*���%.!�+$k⩃�� !!]:��l�3!�dO 9�u�ե\JU8a #�� &!��u�,A�됶q7։��k\�b!��Z)E��Y!!{�a0K�@�!�� )⩞(����
�@��c�"O���3��"/Җm�s�Z��q�"OƵ@��V���
�
�>���E"O���M�xb�����,�D:�"O�K�g�JJB���K�L�G"O������V�|�rEB ���e�"O�E��d�'2��PUb��AWZdX�"O��
���\Vh�S��Io4T��"O�h�w�U6a=����.�p��M2"O���6ρQ�B$�#c��C�ʵ��"O6d�"������{��-���e"O +� ͘T�rI"�/O�v\��"O�Y����@���#	.M*$"O�y���}�ژc'�1m�`4"O��D�_A�(�ÍY;��B�"OD�8�*^�\�XM��f� A�"O���c,�&G�
�c",Pcw����"OVT�\a�h8Yu+�y�N��"O�r�LÔpMB��R�N�}�iU"O���'B��j��ѓ�+V��Zp�@"O��!4%�(Cᆘ�7*?���s"O��@%��< fQ��H, ��a��"O|����� ���f�4Z�>q��"O�����')2�Ĺ�O.M���0u"O�}Hn؜aJD�!%	38����"O�	���¢1���|���*�"OD����pO�t#�bH�c����g"Oh8��KKIޱ;%������Zc�<�A��&��ؑ4l�:0B�}��b�g�<��HP U�V��7��>{I��M]�<��.S<��E�� �����c�q�<1A΅.H��90�ǂ�l&��*�k�<q�;)���T(G�rQ�`��e�<�4�N����&jc��rU��^�<A�L@.�bMB!�%�Bx��eT�<	����n��e�U���@z��iM�<��i�X +��T�x4��	���L�<ɐ��g��Rfz0`(C��C�<�W��4��2�O�J� Q����F�<Q2���1�ĥX���z1�#D�<��_ ���ZRiC�	�z���$Vj�<q��ؑD���j����.HNi�eMj�<Fb� n���d�]
t���)�FKK�<��l\�7Ҏ<qv�ͬ�~Q	�,�<)g�'y�t� mҦhFx,ɥo}�<�����E0zp�震[�X-D��<�珬]]0<�a�[*}$�ce�Jy�<�g�� ȢE��'fFJ�#�&�_�<�G�X�|����ĆNtQj�&�\�<��b�$	�����L	H��#�n�<!S��xq��%�[}�҈�Ag�m�<	�M�#�(��F�	�"!8w%El�<� dPQ`�*�:>p�,�l�<9���ZŸ�{!�:��#a$a�<���tX`A��%�6i��a�w!ZB�<��͑6d���ϰ-9��S���R�<�u�4��uX��N� �F�c��N�<�E��7~ & ��q����I�A�<�"Hߔ\��8P�"^��䡃���<93G�M(��N�I$� �ϊy�<�F�*,nD�Q(Λu�������l�<qD��*D���P�s�QH�Mi�<ɤ�3�����_�Zly�Tc�<1 -Н]�%"��*]m.	�̓\�<� �=�� �1a�lq+�#�Mz��"O0��T���	�B�<#;x}j�"O%�B/HxQ��C��TT8��"O�\�.X�~���@E+�.�H��"O���f�!	6H���J�	�0��"O�a`��C*�� L�F�LZ�"O�p����I�t+P�9����"O���"�j��ۧ��/�>T8!"O@b W�h����,�^@P�"O�p����0���=^�����"O��% T�[q��Y�m�z�vU��"O���D�7&��\zu��)%�,�+�"O���(J���1�^$i#���R"OP�����Rh�Ƅ?�#�"O�-��� �U�4Z&=��M�"O��Ш
]��i�F�þ].R)��"O6p�!H�D$�ؓ/]F�l	�"O���~E�T35N�3��s�"O0̊UE�u�hy���ď*�@;�"O����뛾j(��Q���B����D"Oh4kC�8f�p �d��k�"O8�87jL(�ҁX %�m��1�"O��RrN�?RK�lr�D9`��h�`"O�DXP��V~Z�P�c/wz� �"O  �@Trj�c�T�$d-��"O �����!\�|o��'�|�0)+D�$;3��8F����3��.!���(D��XE��bш���`v�йv(D�ts�m�r^�U�B54ۄ�# �$D�p����9�B����AB����?D���Պ@%�xs��{���Q��?D��3T�\ov>����$&�4S��>D� [�m5!`6� @���G�?D��{����$wNK��g?�����!D��{�I;<�Ys��\m����ƀ?D�${3l�Z6z��-��|�`�C9D�Ȳ��Z 9!x:��̺Y��!D��`��_���H®ƷTƖ!��1D�t����1 b�*S��~l�ŉ�c-D�  Ȋ�4��
'��v�|�a�f*D����;%�\�H�i�gP=y�:D�� !KO�1��H��̧kG*�c��7D���a�l
F����ɄS�@!�`1D�買���.L���L�(��"�c3D� rbŅ
f	xD1�D��I��/D�DC��?I�`�jQF�T��}q� D�(�*T�bg�,�eiԇS\�`�`?D��3�ɑuÄ���@ؼz ��#�<D���E�ГIͲE�� C����Z�!?D� �tǇ�hi2��T�.�N)!$C>D� �ԈT�{z�EZ�*SE\Bv=D����+��u�V�Y1bS��"�;D�0H����A���X�ѻ�%G��!���{q,@��D!Y������!�$�s�=2�nM�~��}�#�4r�!򤑢j�b��,Q"�-(E�(=�!�D_�<*�%/��/܃3�\�!�ߠ&b����3�"��s·	^�!�$�+G�8� f@��Jd���qx!���8G#b��V�܃f2�hB�ۊi�!�d�)�	:�%�M����ŚX�!��F�`�a���l�0D�f$�!�$��" -+WP�{��VN��!�'Y��b�
5ah\c!ψ
�!�� 򰊶O��7o�E��o*��aIf"Oy���B��\���ޤX�jQ��"OD�+��Ĕ�~}r�ܨ8�����"OB4�aiݢ=���-M�c�̡jd>O�=E�d&ϭ��8;g#� SI�l	U����y򢂽a �Q�W�P{��:э��y�fRs"0I�5N��?��5B�f��y�bf6 �:�n�i�¬�����y�/�	��9	����8���0&�y�a��H8�E;Gf-D����yҦ\� �`Cd䍽'W���J��y�	�.=v�=&)�p�p!��y��@�b�d(��Ɲm�&�b��	�y�K�}�j1r�'�0.����� �y�oF	l��p�����$PChL9�y"�R�v���̘}�>U#%��y�fY�:�d��椘�F:(�a� �y��W.@I��\iMF��c�9�y�é;�NI�BdƁe_�PP�J��y��X�4Bƙ�e��FHl� 䙕�y�e����͠"gΖn?l0�G�y�i���T���֘b�������y���t<x5��!a,@�y2@��y��J>M�R�c�G�$�@e���y©}Ɉ�#ȫF���h�#�U�Ƅ�ȓ%ݤp���G�f�����+H	��o�Ł�%aZ���� H�r��l��bφ����\��pm�A�C�A��}��*���TgU	}3T�� h�-&�
����%�U�R�7��m��o@�kHb؄ȓ���� �F:2�4��d�O�S�d=�ȓt����bHG�$gD�I�r5
 �ȓKFvʠN�)�u��Y�����ȓyF<AɅ��}����$�f{�Y�ȓ$���IR���EM��F��u��2���w Pz�tI�僔2�M��!b�P��Ɵ}&�I��G��M�ȓU�f�׌�8N��W��u���heq'��y��0�CO�Gy��ȓ_�;�&]��L C��8�����|RxK�i�>N���@"�!�f)�ȓ�V��fB�>sY M�2%�u�졄�oT�C&�Βd���-��@U�ȓj4��'S8J4`+v⋑g�
���n��{T�2,�����^f`Ʌ�[���'a��~P�h���1U@��J�t�*��6_��Kg�8T��ȓS�H�5B8v��d���.�Ψ��k���3�s��$�F�����E���T+F8HE�y��5oD��ȓ3+< �R���-�~�'GC0:�n��2�Ԩ��(v���i�o9�؆�XG�da�ܠ�U���e��"O�I���M=D�fЛ#�#� �#w"OʍJq(߼I��j�EB0p$vMz7"Oa��+Ǻ#Ͷ%�Ag��R ���"O)��`
>^������,Q,�XU"On�b2$ݖpl�,A%Ҥ4)�"O����D��bQ@x����ZƼB "O*�b3��'�p{�L��9p"ON5�C�	38�q�d�@�oڕ��"O�u��uB(���� J[��q"O8)j��^�pzB/�]��%��"OFE{���n_v�� G˓x��݀�"O� ��if�D$^�:�ab��.rR Ö"O|Xs��W��� V�Ð.ND�O$��H�>X��5��(@�����U�n�!�D�8<���x�*�j�|5��`Ğ�!��4& -��hT�h^F1��ݾ !�DG����kg^�A'�H)� �;n�!�d�*ZhT��撥b6T�'iQ�!���4$_�0T�۹#�
��蜀;�!�d[.�`H���5��83r���!�Ć!`X}���׳	;��A���[!�>I�Z���"�a:�E�j^�D[!��H"r9Hc̈]3(D�*A!h�!�:=T�r�*�,~��v+� CC!�RQq��&KKoB���-Ց);!��V<e_�`�O�b�Jѱ�T?�!�$�|ܴ<��W�[�8��Q��0_v!�(.J��
?fX��B�N@�!�˪#��3&m=(���w!�d��Hm��)RD�7I��Q�n2k!��l��@��C�; p4� ��!��8)V�U�
�(
NM�h�(�!�D�% �
�2���6-�4%M��!��O�Dr����E�j�X4$���%�!��3|x���e'=MŸ`(�l�7I!��0.�^���+O�0m�ǀ,?!�Z��N���EӣA�2���)ߪ:!�� O�����;�ea���"r9!�$Բw�`гCB�C�bЃBe#$2!�G�Y&6�,SC�=�eJ*�R��'���� �L�.0@��*.��'�B}�я��B|~��j�>fǘ��'5r�y2�C��i&�2sB���'E$Q�s"��C�/"ؠLs�'�u:��߷$]���4D��H3�'hu�T&0s%���>#<���'��}� �I�KH�i�.� �8�'�.Tq���%�v\Ze���:���'�����: 9 ��+#�#�'��y ��,8H4
�Y�)Q�a��'����q&ǚb+�[p M"TA0��''��#S$Зi���;G1��0�'^t11�0L���� +�'Ӑ�x1�Ӣ:��27��8j��P�'z�q�&�y��.�:݁ơ�/�yR@f�@Y)$������Eӯ�y�BH+���8C�'��C�,��y")V:B'-�w&L�p\TH��'D�yb�F�ؖ�r��ޅڽ
�AA��y2!A�+�� A0NӪ:��� ��yr� ��& h�U4.�8}�eH��y�b��wrd�%N��n��y�����y&B��(�Cd*ƈ�DGF��y�a��OpPT�s��>E�Љ)D�_=�y�a&x����#��(o�CF��ybE	"�&�X����Ԏ��$B��yҭ�I��,!�ؓy���G%� �y��Q�0h�dm;!
4튓�y2)���� q�[(=h�1āE�y���5{�J�S�iI�SZ��{V�V��y��K�r��B��Q����V�K3�yb@ӯ]�4��d�L1C���з.�y"�Y.T��j��_�C��|��¸�yBM��Y`�E��iBd�ae� �y2I
�b�� #����J��y�II��y
� \(��p���H#���"OV���Z��e���×M�4 ��"OT�p���M�"u��B�d�X�pw"O^�)��OB�}ѓ���2iز"O�s� ЅC�^u"1GS�<4\a۱"O�p��� ���Q�}���R�"Oj��+B�>_@]SqN<���G"O�pH� ړj�J�˥F� \{ތX�"Ot �b�2�	�g�Ξ ^HD"O��x'��`�!k�H
L`���'�J�SݪxvH��#�<P�����';��k!�B�e�yX&��_�L*�'�̰��M�oH\$��,',��'��T�����,=(5́:ꐽ��'�x8J#L;T�����	Z0v��)�
�')X����W�.60�����t��I!
�'� �������
6�Z�sH�a�	�'���h&�0��bn֕nP8���'F&8�O��4�R7lƎU@�l;�'�`���@�w�L�(�'��P�� ��'��x* ���=��	$�L���'���d��}�q�+�u����'�.�HԣȪ7�c#E]��*$��'�Z���o�*'4�s�˙oi���'�Ha��U�Xx*@#H�?Z�>%��'��p[�)�N>*LJBʜ�c�$��'��P"�ܑzTz�`&�
Vg��a�'�ZTDCM�F�P��Ռ�:���@�'nn	$k�1���÷3�r�q�'�a2�Ir˄�@#�zrb���'�f ��AvR�5,�qܒ(!	�'E�|X#�T�#e�RB�g^<��'@��oS<C2hI��2Wp<��'���RU��,r8��� R��V`��'��=�5�H]}F�jB쏠x���'�$��'NL�)ʱ���ġ�'?��+ьk���
(@`e��y�bat#׻t��Ɂ�V�����'�ڠR��I(��lk!f��Ʃ��']�t�5K]�>�B��`��1/Uj���'8�� �Y��@�I�*UzMR�"O���c�!(�EJ�OB8�)!�"O�`� ��4[�(T�7F\ S�<bf"O.��=qE�p��A�:���Y�"O�I��l]�F;�q���Dv�3c"O�`d�0*T�F�޺?y�܀�"O�1�J
Ewv���:[8Pkq"O�82�/g���³f\�NLP�"O�p5bޤ|�0��D��WCD� "O�+"/·!3����暻���X"O����"vJF$�D�Y��A�"O��SS�Ġ!, �3eI]�Ay�Q�2"O�=@b�#l����- �T�Ƅ�"O��!�0�l؆,PC�$�p"O�� w��)	(�:� �s� \��"O��
a��m��������"O���AA?|}���S�A04�Q�C"On�[�`�q�R�@C� ""O 8�e���g5j��FБia��"O�e  �"�rCf	�}���+�"Oź�]�1
�h�B㒅3V,9ڐ"O���������N�x�5"Op���{Kx
a��}�8UJ�"O,��G�V�rV0d��ϛ�S�<���"O� ���g��
SG�y��'�Wh��1"OA	�!Z�P5H��P+Q��6"OPE2�V�>J<����1l�y"O
��viE� V<��Ϥq&*X�D"O�)��	�OW�с�'��sS"On[�a��M�.�i���s���1�"O����Z=�� �(�2��"Oސ�@N�#�!�`�اq�ʜh�"O�2G$�������,I4<���p�"Ojh1PgD&,5xhb`f&��,�"O<�;��C_n @"�*��%)���y�)г`�@�La؂`��y�BJ�8���)�nN��q���y�F\z��3Ȇ�Qs�A8��к�yb&�h��DJ��:�*鑖B�'�yr,	f@��$���.2V�t/ǉ�y��5)�	aJ��.9�<a�[��y�f�'����e]:2Np*`�E �y��_,q�pDY
~5~��g�U��yb��ICv�j!�O&+!�F���y��G:����S.k����A��y�o�� i�nL���aeE^��yҫ�77�D91֊�4E:Bgޙ�yҦ�:&㢅p�Ț{4��qHH��y��5~!�h镋�)�m[QO���y��n{/��3��".?��`'Ȟ�y҄��Y_$�*@��>�|P(����yr�P�T�:�mM�`$P	�f�_�y�φ�K����m=Y���v���y��7���g�<U���CF��y��<\�����]eRH��ĄM7�y�ؿ2��!�	�[�-�FO��y��_2��h�r A��U5�y��7_`�Ԙ�$��:�8���;�yr&�	8tLp��/4M�A�����yr-̅�*5 0��{��)¤�׬�y� &;ETQەo0H����#��y�g�0(����U�8d��*�,�yB�!~�}C%���`�t��+��y�Ǐ!4*��`-@�a��-�2�9�yd�/F���� ًB�8|p�� �y��
g��9& [�QhvT)��S��y�G�����Hk̻@ˀ(�y*èpM�A c�x��
ω�y�cH� �fF��z&���7�D��y��F;�F�eS�ٴ=g,���yBg��	̬th����{&tI��HF�yr��@���G-^#o��X�S㔲�PyNM�7d�<�g	��Hײ���Y�<9� \Np��0CN���A^�<yB��(hI  ��#Ѫ	����!�\S�<�	�[r�q�C+53��*&ƝK�<��[�Lܤ�AF̦(���35Ko�<)�aҷ
\m����Xڞ�C�	Ec�<��LN�hp揕�lǔE���\�<)�͝�%HR�FQr�^͚5��O�<QT�ڵ$ur�� kr	�V�VM�<1�LN+t�
=H�%��Z��l�K�<�F���q�.4y4�$	2�I ��F�<!��B�*��-�q� T��ՋDC�<��$��մ��2���I ʁ�%-C�<�dl�F\�J�)�����@�<��
E.X���M� ���󠊅t�<鰥�����P��H�TM�`�l�<� ~���B��9"�`Y�������jV"O���$
߄]�tȐ�#���""O��:oN��EG��l"�mq&"O2��N߫H�ld�!G����"O�PJ�(X2�Q��@�6� x@$"O�S��-!At���U���"Ot!��<�.��A�x�|�C"O�q�W��m�c/S�:%`	KA"O���s�^�2%R%�G���"O�50˒+~²��Qo��X@t"Ozu ��X�]ބ��e-F&lc\��"O����hť	�xY+ ��cf��81"O��zFl[�@~��� \R0a�"O��@�iQ7N�X����/��"O�8Q��L\��C��YKn@k"O9I�C	�C�� 0��=�Dà"O���L�60P �BLș�f��s"O4�Pgk$V������R�q�hDz�"Ol@��O�Dq��+���V��)��"O~�fCН�T�0�Ҳ-|�� "O�i�@�ǈ/��h�����(���"O�	��؆t\H�B0i�-q���	�"O���IW�Re�sƢ[��x�"O�	�'�/n��0���<L���[t"O(j�E�:Q��)�*�T����"O�4�+Ϭ�$+�/�5B���r�"O���ģ��&F�bQ�N''���C"O6L�e@	i�$LYū͏i���r6"O4����@�h�ZVj�d}DԛV"O@q�'�?K(�$�W�`���@"O
��$�Ӱ~�H��Ѥ���n\)"O��'�^�2�.`"���"O"�"�,�zrlS`!�.JD�0�"O=Ӡ�{���Z��ٌ?��G"O�(�DC�W��Ơ�
��"O�P�F���3�<M9�̑~����C*Oz��`�?6��t��)�SGpK�'Bj��v);���+Tox��
�'VL���ǈ�v���&Κ�Bޢ=`	�'�Q��IF�̄�1fF�B�t���'�r�7K��a�4���<�,��'˪H���Ԅ�̭Q�E�:����'�>I���ov�]�R#/�xT��'W��؁�K�`E���H�{�����'z8��#

�%( ,D  @<Mc�'��u�uE��~�i6��;kb�*	�'���9�*�'kh��p]3zt0r�'иqǀN.�|J'č�-Ҙ���'I�<&,�"B	�&咇Z:�q
�'o���a ��G*���`�P;M�q�	�'b�E��d��r�P��g$�/���k�'�z�*�+F��pA�EA�#��0�'���gL	����2J�@���'ZN��w�іE4��j�dF
=sH��'o�0���=k���0eK"8,� ��'�.1[ �F�d�b|�R 6���	�'#��+�Xo�t�q���4�>���'���(�ʞ�43�"�Ŕ�*YL���'�L�D�
i���j�G�(���I�'��S�b�:�|UJ	*5^���'��m�!cW�X��M B�U@���'�J�(��%[�5�v�27d�|��'0y�!�3`1�8� ��5N��

�'v����Ξ�*�) ��V���*��� ~0	�BP�vtԡDo3~���
�"O��u!tb#u蔙C�Ld�U"OT�K�卋x��x�c�Z�r�F��"Op��M�,�pJ�+�J\�g"O����>��������""O�<� ډB�xd{��Rzk8��"O���)��BCx�a��"S4�J�"OP\P�Ɉ��8��J-@D�; "O���Tg�
6�����W�����"Ov��'+��w��R'�F- yH�"O�{a�=?,��'zfv�1�"O2Q����9p���R$�:dB�i�"O���whÝ�t��$S�'2)*�"O�����k�
����%L1�"O�)y� �5�P��cD�@~���"O�u��%	2��H³JΑO2���"O:���O�f��1������B"O��0��P%~x��R ��+%�L�"O�ѲA��t�>t9��6+y0��"OZ�(V�J�C�@���EGo��+�"O�l��T!
u���e��n��š�"Of��A	p�R�y7�Y 䖇�y��<�%ŋ�QǨ�sFǬb�E�ȓVA�	�s�͖E8�h��,�$f�|��I������*���b�,\�����6>�x�S��"\{�iCGIT0�L��ȓB�� ��CUj6(�ȋJ�R�ȓZ3�I���[OvIh�ʙ�d>����="����FXS�d+�Z6���ȓe�D=�$ğ+4�2���k[�8�����f�%�b�H�d]Z�0�G�}���@OP�  	�:���i��gsj���5�2�c2���g�И�r"^~YZ���Y�h���Vn��,��L̃k� �ȓ%e���ԪG�V��2��6����9�|t��$\�����s��	�ȓ^zL�jC.O�(`@�;����ȓf_�q�1�H��4�{�"O�|�����e�D$)��
�K�z"�"O��B�?��A�R@�2|��IH�"OJ-p�ѷc� 0U%]�A����"O½�w��|)Ru�Ԟ76���"O:�Y�j����}�s��V�T���"O��P6H��3D�m�"L�T��U�"O���f�D�4��xГ�w2p܈�"O|�b���ڴ��$�B'"OPHbu�B,0����2f��%���b"O����#ښ�f�%F]�6P�X9�"OĒǄ�:��%1�%%o;�i��"OF䉢�J�l��IR�=s �48�"O>Qh����8��CN1��-�g"O��Q֨
32�0���ؽp�8�ѵ"O��SF�! *��"�/zV- �"O�d��e�3S,,@*5J=j\�͢�"O"ɡ1#^4'�2���V	�f�9�"O �˂
+�T1ʑ�A8dǰu2W"O>a�c6Ay�9�0G�3:��	�"Oƀ4�[�,���ܖNаZ "O�!�N�<h�0�e�ӆNjh�*A"O�q���%���td2d!B��yҋ� ��܊����@8
T�ְ�yr�
�Z��$��C�G$�yBj3�4���A9�h�[��7�y�"�	X:�� �lV�r�Z��y
� �X����1R��C�K3.:\�[�"OZ0*pĖ�^����F�Y�t��"O�Ыv�Є[�����,Z8OF��XP"O$8PB��':������l@vhb�"O��g�{�B����|8�L��"OJAGѭ,hp��G�0ϔX!$"O�p8����6�#a�8Q���#"O�u���K���u���-�"OH���G��N}rvH5y͆��u"O�0��m�9"v��a���� ��"O.�W��*��r�Eڇ�r�9�"O�����0�t�y���J���"O�d�G
���څ`&A�@fV��3"O�԰4�Y^�}�0���Z��P��"Oh���C
D	2��aC�1;?�!`"O�8"�b�68�y�,Β$^�;`"O�`VBO��+�i@�ir���D"O6�g!�#8l:�+C�QUz}Y�"ON�C� ]nM"��(�8a"O���!*�5k�����W�3� @��"O�EK��,:���k�d�%.��9�"Op��F�b����@]�R�"O���`	-��X��BT0y�D�K�"O������x!��ּ;��Љ "Olг6B>� ��cL }��}��"O��8�I=0Ź%���*���!"O��ʡ�8vi |���V/ ���"O"(��`ߓYg��:0�١	3�ĉ"O(|�QB"((�q�Ä_-ё�"O�
#�ŽK_� �D�i���"O���vG�3.��#$ĉ� HqZ�"O4�;e��Ĝе]	lr�Ö"O��u�� �T8�ځ2�*u��"Oܸ��b�m��\(N�E;B"O>����+^%�E1i����"O�@BB�֬&m�]���:�̌�"O����#rh��
Tz�Xc`"O&��dE?Ax`)�ܸci�D>D�2RJ?S��� �Q�I��U 2L;D� Q�i� 1����~%l����:D��2/��]ل살M\8g� ��f;D�O�;H-Ö'�m�&Qŭ9D��B��
<��3r۸O� tc�B"D����L�6�|l�EY=;�I*�?D�DjA1ef^���٪���#�>D�J��݀2h�Zu�5����g:D�lcā-m&��a�T
>L�h��6D��R�Лo�d�8�,�� 6���'E!D����4m��iB$пj"�i�EL;D�4�f	�F�8<��"r����h.D��R��C�&���J�a�2��D,D�bTM�*G����9*���rh?D�D�a�?~�Mx¦��j��1��=D��v+¹3��0x�,�xp.Qh�=D�`�,G�z�4�&�U���u";D��C�J��e�l'�ã 7���b4D����ߕE�r�@U�·9���j��1D��Z�n�?/����M^/V4��l.D�P� d\7|���uI���tRF-D��y"���L�) R���h"G�0D��x�˖N��L�s�@i~�PB�,!D�|j (תSq�����56و,hC)!D�D�u	�qz~�{���?��T�?D���b'	>+`0�S��tG�{�k?D�� �@H6�%A�����U>H���s"O�I&A�Kn�� G^3&�$���"O}��m� �!恹7�,#�x�)�|>�E���*&���+A�P	%irB䉟X�J�ʈ2�8�W��C|�A-OL�O�3��vР���a�OBqe-�6����d��<���s�����a0d*u�U
A")ϡ�D�4`�B!T�P$
c,<iD���O�#bd^P�(9b�%�Z|)o�<��.�&\@p�d�:=��`���m�<C��#&:�+Ӡ��;���j"�	f�<��V&o �T˵��Q�����	O[�<1��?opP�95���
�"iYW�<�B�ů)��U�0)`
�h�S�<q�K�Qt�8�n�J
X�o�I(<�ߴq�P��ajS@�9#�(�@̇�Zz�H D E�7�� T�Ի4������h�'�ڸ�sh�(2 (�c�i���'X$ʡE��{���&-�#K��)�O̢=E�&�o�	���4�|H��E�y�G�%.� RG�/��ɉ� د�yB&ȦU
ĝA1B3� e�r����?��'�0��s���P�YN^I��A��'����gV�k�E0��Ö��)�'���Y�' $i�Ir��f��'�ni�sl��A �똖��d��'���s��w��zD"V{���'Y|��#��)d
��t*6j��H
�'R���Ťa޶(YC/�4K�'��T�c��%
�(v囒X��R�'���"���o�ڰ��CYJ튥��'��p˰)V; -��`.���ȓ`��+F��+`,:<1�����ȓ���� �{{�(9P]�	�81�ȓ�aX��z�~ ���ݹv��X�ȓw2$ѳ��N"0� �u��4D���ȓ\��Q1�"�
$�|�SD�2$�Ň��0}�ǫC3��2DbTo0�h��2�����O�#dH(�AV@-8�ȓ1)�@@%`��5Э3�'Y�.�����F~&x��.�
���s�! >5�t��}*4��kC.�r�ʤ-��؄�e�WI��@�`���,�D�����V+�Y�G�(��Al��s����bIB�G��~Jt���$�b�(�ȓ~�-bq`�Q�����/r4ن�s��$y�A��M��'oPf�����a�t#;����ޘD@�����Q�H?�|���O�0�ޡ���l Y!i�;[(���jD�L(Tфȓp�ȹ0�l�*'S$x�� /�,��ȓCl:h)�'�<oy����g�r=�=iK>�$2h�����-�!���Ȱ&Z`� �ȓ�JT�/��/�\�pr�ÿ|6���*k`�[����W��7iDt0w�'C�O�6�۽	_���ŢJG�d1A�Z.d�!�DP/�Z�z�K�m��d�@���!�$�.g��iB�D���&�:�K�K�!���j��]ZRo��a�t ��#���hO�$p���m��oŝdZ��c"O d�g�D#F^B�Sp[�!b�h��"O����o�P!7TcN	�G"O\������12%�oIl�@T"OB�����]n@��O!}���1"O� 24z�$�
0m`,��,��Fؘ)��"O���=�HA",�5���1R"O�+�n�/tQ������A����"O��Hr�ԡC�ƀi��"EU𝡳"Of�KwHTĖ�#��
�K�6"O2%����2ZZ��!0j>͆�2�"O���P��s�IL�S���2"O`,���ͰZ +*	��rQ$؇ɰ?�'28Qy���!2;h<y �R�����{��)�)��>j|8G�������i�"�!�$Zc��1��
��@a�Ї\O��hO����8E���'R5�T��"O�����9����QA�@A�"Oys*ʻ��rdnP�$̨a��-ʓp��O�Z!����Hkv����/�B4��'�"��C�c�0�*�N�x�Ï��b��t��O� W�
*H=Pc�"T����O�Q#�{�8�)��z*�]K�f�#��xR'�<��;�%X���ϔ#�y�J)a���"�ʏs��({E����ybH��OG��Z �۴nF�x��ؚ�yB S�G�L��DG/n�89*���yr�Sm�aҠ�	�Pg��Zr/ٜ�Oȣso�"
:i�q
@�j�"��� ]e�<9�J��c���8���h8yDG��<!�^�<$��g̓G�e��gU�B�D���߅#\��D{b�!�'$����_�t!�S� {]�uX�/�t벁L�'����ӯD�9��v�#LO��2X�Ib�F�0'ϐ;���@a[('W0B�I�gL<9(���"+�"�(c�׈\	�C�,x� �8!\! L+���)�����W/"��	�W>����
��qS�J�tC$b����ɠ)HQQ��g
Ju��6q��C�IȦ0���칲7E��?'�$��i�{y��'�x�{��LfMR�K2Ȕ��'RN$�4�v���qӊX�:ٲ,
�'i�!�H)A��J&e��;=�Pa��ĒS>��%C��2�耑���	O�t��k;D��r� � �&�Z�*��78�h�L;D��a��A��t�p���y �\�fj:D�,!�	�@T��J��W�/k�B����a!�KD�ny�a�\hC��/k�0��`�CrU���c�hB��%������"N���#_�gC�� x�����S�m�D�+��ܱ%_2B�	1Ѱ�[(r"�ء���B�I�3�)��'G	�\q��\2�B��:�$��g�&A�Ԙ�K �z�B�	��$l���
c����l_
�lB䉜�j�ʑ��.8)��qB�J�YRB�I��� �UF�)ܒ` '�ʺ8ZB䉕Y�d����M��I[��C�+o$���"�pj@�g��Q��C�I*{<��B@SH��6GE�c��C䉨IB"��%�%j�*��Dm�!{��C�	!e��a�XL#�)xtC��BHC�I"J�Zeˡ��
�ı0��	C(C�I�
�س�#�T��(���S�kvC�	=Ju�!s򉒩~`�IR$��B���J�9��P�^@�aOҳ�B�ɍM�nȐ��A�C=@��%Q&^��B�ɏR_�r�"EL4f���Q</7�B䉴tw�����T[��R�;ΆB�I"L��qb�-�3� X�fpM�C�)� $�����J)��?f�<{"O$Ȣ��;]HVQ��ʎ^ �P2"OTP�爃8� q�hL\�>Yr"O�űR
��]o��P�ɉ�.ЄH�5"O�D�3�,Sv���q"�+Z�[�"O`�K��F�X�� E_�H��"Oĩ��/�s,����!v���t"OR=���3,Ґ񒅎�$-����"Oܐ�$�tj��U�Ϗw���g"Or-��ȫd���G�9{��e�R"Ol�.(bT��k��\�8� ��"O�5׎�.uZt*cD�=-�����"O���C���eL�|��Cۨa��F"O� R��ty�����ɖR�T� �"Of�s$��(�(���, v�!�"O�L��K��T8�)�	F��y)#"O�ثbM�B�Nx���DLhb"O�\�R��#K�27H2I����g"O\���F�Oe����R���aS"O<ia"�i�����u��غ"O̻�D�蒈S�[�^�i�"O�d����%~"� ś�3{��) "O �xS7Gڰ����H[����"O��:!)Q�L3����-��`��]� "O`�&�Be������7p>d%S"O�,�5�Pa6(S��'$/dXX�"O���(�d�d�!2�-a+�<��"Oth��)1^ ��+62����u"O�d��Z>J�p$R�)�j���;�"O��S�p�P��u���\e�]��"O4i��I�*�@1�	ڨEG�As�"OR�h���(�+>uM���1"O���F� w�� 0���-a39b�"Oj��]�;N�q�&O�eI:U��"Oi��l�-�n��끐n��<��"Ox��aq�p��,H���
0"OR �$�"*z���� h(�:1"On���I�	:� $J�9B$pG"O���,)K��Ŋ3��-�5"O*�� Ñ�Z�`��0j�8/�.(&"O�0z��/����	\:�fL�W"O
0�F���Qp�]:��
�F�R�"O~��mG,!N�1i�a	:� ��"O��S�Y�DX�RL�w���qV"O�z��|��[�F�R�H���"O�H��Õ�}J�y�n�?
�Q�"O�Q�D�63��,�p@��3��U�D"O�mz��U��^�����$z�Xq�b"O2LB�I&]^"���-O�?��l""O������]t@(�� ?(�;�"Oh ��$@>�)�֚]�Fi�r"O�t���9X\3dlԦ�J�"O�x6Ί%u��<�Bm\$a "O,�A��V�m�`�9,O�q�g"On�9�HF�`��9e8PDTA���*�S��y�͍�$-&qi@I_M{F�I�K�y	�(_��C�f�� \��eɉ�yb��p���C�U����A3�y�M��jXH՛1C�=���(�_��yr ۑ���1���:_����4׈O䨪���(4D�nJ&�����<�!��FQ��L�&��R���5�с���<�S�O8��KQĀ�e�pĂ��Q&L�lm8�',p���;s�	��?�$�P���yӦ�� �Ŋ®� kJ�+�mR;XF�t��"O6��  -��m�7��2$+�hB�"O8�x#JK�*���!�� �Niqe"OX�2K*+����R�%K&"O����T���3�B��B����q"Oj���o���Ij��B�%���"OΡ�&/ү-onP��c�f=8�#"O1�DJ#:P���K� 2fd��"O���(9�:a[E�ϊ`*8�xt]��D{��I�>5Bt���3Ρ;��&�!��b6*��W�N�=�T��"�e&!��ޤ*M+)Q�i��d	7�)�ȓql�����P�p%������!FC�I�'�N10�Ɋ%vpiy��!E��C䉩�~�PpCA-w����ᣛ�]�C�I�Y2�H��P<����V�D�C�ɠq!.��1Ǎ;���Ok�B�ɮ҄�xS��-{@b\c�N�B�,q5l5r�"(u�1��J�B�#F�z����yo�E��R^�B䉻<$Hsď�\� �a�3=|�B�	!L�4T� D����1�	�5 ��B�5HU��K���'��%�����B�	��:PG�"_A��l�/��B�ɶ���р�S�91ބr���c�hB�I�K�T�D���$h�裂̚�#��B��>cz��i�j��8ɖ�Q��Yf/�C�ɕi&��s�Iߑ?�ĤQ�k!l�b�,D{��t,�;a���Ќ�5 �H��p<���Q�tG��� I ��s��=w!�$\?YBX�����Y(��ܿp !��J)�Ao��,��ܸ�o�&�!�͛O��ak�"U&������.an��d9b�8�&���-m�別aL2;�C���\�UmC	C����i��>�dC䉽\h�]YC�#B����҆�5k�.C�I�nK�0a�'�=%#�y��B*C[RB�	� �4Qtl�2�h�ҳeڱ9�FB�	"_��)�H�*fGR��)xB�	�f���`D���u-�E3�#�T�C�ɴ$�(�R��{�M�d�
��C�-���r�Ȑm���QIƴn26C�	��(�ك�1���UA�i��C�	�c�!A L���.-;��� ̨C�ɊzwF�{U.\ o����C�{�4C���R�ۧ�`]�R�@�+hrC�b(�Y�C�&�yhî�?�<C䉉F&v}+t�_�j;P "��+r^��$o�S��ƴeH(�F��#^���d�%D���VEϳ|�B��D�@��4
!�Ʃl��$řHibx����!���8�tiYb��dQ�y���$A!��P%&ޜ���E�����:%!�$����$�G\�2Bh9K��%MqOd��D�FEtU�E�ŃRJ�"D�56!�.Q���g�&I���0��F/ay�剰_R�1�c�
�:y�㫄� B�
s:x|qU�*z���C��zb"C�ɪ\���h��.�lSt��[��C�I7?�P`�B�6v��2M�#5]jB䉽: �j�,�'+�`d00#Ӌ6[N�O�ꓝhO��y���1� ��J�J�S�	U,B��-̱8�!�.OO~a!�"O��sSh�>�tQ��	�a�"O� ><�D͖�_r, ��J<�z�)�"OHu���V����Ѣ�&Q���"OR�9P�P�
yN!R�C�]q(��D"O��k-��)��sTc�0�(��y�l�?�x��dL�$ I�i���yr"�JN�x�B޳{zi��蕆��<9��D9�!�kN8���H/�!���5����㛱oIf��#��i�<����EN�u�E��H`|�pՅEf�<�CH X4��U��:$Ɍ���^�<����),�=��蒼|���S�A�pX�@�O�L�$�[�^l�8�m��2�∛��'��)�T�QN�3v�%(GO�IO�O��C� ��Ro�"��� �T��u"O���H��G���"$`(����2"O4)t(�rJ0�oi�� Y�"Ot��k�3n�|��X�<>�A�O,�O����2L��F�)N�$�p� /m+!��� 5G�3h(�Y���t(!�$C6h��4
 ���1j�9H$<!�Z�ڐB�e|FM��I)	a~bS�@��Ɣ6Ҁ�8�*R j�*�I�HO1��)��!_W����"��<V;�0�C�IH�O�$@�SșqS��Ѧ�Sj���b�'��E�2+�$V������ȴ]^��ّ�"|Z�'PX�[�h�	�Q:ebCHߪ���'V2�w�Q�C��:����@M~�[�O�"=Y��¨C�%��nP��j`�5'R,S�!�d�,���Ct��<��3���*���hO�đ�$.��vC!#^�\Z�m��"O����|��ܔx�(m� Ĝe�Đ�'a}�HS+��C���i�`���0<Y�����*�n��Ǐ</�h �g��x�!�$#e������vlP%+�!��3���!��ۇ���薟E!�D����S犃s���Q��)[!�$F��9������d�I�|�a}�.'?� OC�JS����oY�@j��H&��d�<ir��&;f�$ND�*�,hx��KE�'{x�����{��YP NV�pĶ�c����<iǍ"i�$P�1��	IW ܫ�"M�<E?O���g���@2G�g��E�� ?��=�ȓt��q�	�K�~Ի��V�r����ȓKY�T[R�K�q���w�λ>N
��ʓR���D�r��U��j���'ª,i�⅑gfV�u���]�:i)	�'�<�0�D;��2�
�W��*�'�<�C�5}1
9�D�ԈOM� ��'E&���O��Z�� z���D���'��z�ޛ8d.�YD�?��I�'{h`��M�)Bж�#ի������'��Yz5JX�/���DF�`}:�'���������IP�6y�Z�j�'W�t!�ȇ<>��4��>y��0�'�ԉHbb 45��{��ϕ��|�	�'i���d@�$�R���|E1�'a2�y�f��
t��Y��(�S
�'f�لo��O� 	A��_�yjK�N�<�c/#��!b�&Q7H��`{0�I�<Yeh�Lk�$���3�<s��I�<q�OWy� īw(��0���B�<��g��T��	�\�b���<��B$�q+އs5�$b3�]|�<��j�Cx�������<ʑqᄀn�<� <|31�sP����U)rc���"O⸓��J(@�`�	��Y%�X��"OT�S����U�`�Æ�=��S�"O^����E�&�������R9�X�G"O,iq�V]4�5� #�?6l��"OB�%��% F, b�%I��٪�"O���P����KS Y�P#�9 "O"��b�5b���:f�5<��ӧ"Oj�X�1R:���L����"O01�2�-4Od� lפ&ڍp"OP���(�f�r��Ǽevx�"O���JNc��IwIܨ!Xv� S"O(Ӄ�R�l��4�v/T�څ�"ONA��˪8�
C��&Y�l��"OP�A�?D4���T��-r�"���"OhH��"��A�TYф��x�&Q�&"OP�se>z��fD�>��@�"O�$#e$�
/��U�Ą�$ /J��T�ɯM��[��J�(��i�4d� T�_��(*p$��`Eو��)�h��ȓ7C�M�F�(mN����N̪Շ�g��9W
ժ�$��ĖJ㰴���`�w�G�x�a��Ój1v��u�]s�_�6�0��2F��$B���c �M����!�,U��O� @*�ȓS����0'��Y�j�0��%��;뢭�hH�Fu�����X�;����q���Á4ge��� ��2X]��{~�wC�$"DT���+qG�ȓ�f�� 5̺�1Rˡw�����oѲ���[�n������9�Щ�ȓ����7GT4V��G�0瞍�ȓG��6#S� fVTr��4jBv̄�!�<e��ُfC�����5�6���J��tyNHp���q�-7�X)��Qm����<�I��Ҫf�|ɅȓE��ճ��N�Q$UYgL��YO ��ȓY��)Ȳ�@�Z�F�*�hL�c�4�ȓ+Kҕ���N�6���զ�%#L�I��Y���Rҏ9th!
QDV�t0f�����x�""pG)j���?S/>���j"L$�4g$ 0}�c��a����!��14e͌r\A5�δ쌄�uI�4�DgS%}�H�@`Đ�����4e��ʷII%K���ʶ �ȓ� qba��p��\9� '"O�hrc<p~x5z�!���ĉ��"OTQ�b��rs��*ť�9�x���"O��{c#�+"��8*U�D3/E*}�!"O*�����/E��	{vܓ,n����"O���p@ؤr��Y���^$�R,�"OnA8�� W�Xj�`�g�z��3"OTq�w(3AEI���� :w:�x�"O��y����PU��MGy��`�"O<PC��;#^�2Fl��%}n�Ʌ"O�eC�(�-I�dx�lŷs����"O�8X��L'���z��Q�XZu;d=O�p�AL�.w�a|���a�n(	�A�F�������3��=q�-�.N0;��'��!!��E$E����,��>%>��	�'��U�u�O 7�nD��'4�JEɈ}�d�>PW>�I��H�Α�G�Fv���fMID�"O���g�b'���DT#1&a��I]�?w�$���D��(��ɟ|&8�]�WRh�Y��5ar#>��O$�0���jJM̧Y�AK�ɮS�^��G��/�)y�%�5gĂ�r�ꄉy�����_p��	�jd�;���]�h�DN1�!������ק��艈5�5�W�,D<H�� D��'l֮,r0s���s�.\�2"Od��n\�8pD�9��>O��d`"��k�­�#ǔ \H��$�%/~ �f�ܻ;q��(�t9�d@d��q$��0X���¾�teCpL1�Onh����FuU�F�%�н�p�\�<&ꔰ��Q:4"r��-(���C��N��B��&�ح�0���'T> t�ϳr����&�D��ʍ�D�V��\R�ȃc�!Z�M�3�c��J� �P;C�oZpS�a8,��bR��47�R�@D�0ؘ���'�J}����"���l`S�˔�Y��"�J�#M��X��!Ʒ�Da�We��,1�Լ�pP�1m��Q��U(�b�+(H��LG��D���l+D�#4䗯lm��X�F��y; ��LĲFJlբ6_cbB���c2J�H4K��֮mo��F��?6 �le޵��۵%d�s����t,(L�ta"�OȵS1AK&D�� � >$)`p/�$=a �4�x)���*�:��ђ�^U;��I528�O­!!YH�`�m�}��`I%ۖe���+�k#~Azq��+"��B�O5+Ɔ鑗��hҰ���O��8�~a� C58��N�8�5��ֵ	$�i� �%�ቹC����~fmh��K����;QD�>}��1�Ad��Q^:H�1ࣇ�up] d�i b�G��6@�1�[���5x���R�L�;�m���?!p�.W����qȐ7=j�|�Nܿ�6����� a��O7P��7MקX�V%��CѢhr�ԁ�*\;�yW��-2��9��ʨ`$�u�#����0>)�,Ü*��a�aW�Z�.�WkڍI��E�d�%U�,�E���p��͸-\�L�>6�Z&��i���7����6)�L���d}�캓�ʊ_�n�b�a�6�P8Ey�h��gz���3�Z�x�:E��1�N1&�-����I�<CܤpB/�*�h;�o�x���Ka�!��)�l����t *��,c.y21c��<@dP/Q��J�.e"er�C�*8Ivt�P)4����S�<������j�4��݀5#͢r�V�;�lB0cf�#�L�\4�<:��)��1	!�Ԇ-J>H E�Vd���B��VQ�"��`BD+�(.��q�HuӀp2���o�Ɯ{�wԘ�h"�j��=Z3���UP�0�O4h�FZ2KX�ˣ�ƶ'hDE���P,�P�D?8sftS���M3q�c�����iEȼ�ĥQ�0,� �Oh��Z
q]��+��!U\��3��j*�ei��,�@!�#ηHt<a��B9b��{���P��Q���Y�#�0h��Ɲ?0&��x�k[k6�}�I�*3���$��6-4D��D�1۰�m^`�bO	6j�I��05��	��@D/���!ӆ�cZx;U���X�ʞ��\�`�/V�B����',4Q���'4R �ף�i�䫤��NU���0y0��Aq���O#*m�@�2Y<���yݡ��r�)���R�D"��k��a ����d.D�d���ͪ�Rݘ��_�\��ȕūb�U�
�����'b�`��'�������p�JgEC}��"<8�j �PrbEc���;�p=!4�\Z�V�I�nG
��+�DK�O�.T��a�h�H� ���=B�ؐ4��-������2�S0�*�Hl�z�	-��)/N��ѣ4e#��m��A���RX��Pj�k�*m���&o�&.>��޺s��94�hO
!�Pk�mݼ~����w���>Y�h@�c~$lSӈ�(\�&%��D��T�t���1�"��E���F#%��ds2HC�)_�,5��d��WI]�m� �f�K��§e�A�<��G�(t+��ǳO�=⦝��n|
aôe�d�ġ2%d���L$,x3�/2K�k2���A�TO��a���ɏ+DքYxc�G8�\F��,A,�;�oA<Z�L����Ѡm}���ve�ԋ��U�~�9�gL�o��&� �\�V��ቀ��S�EF�J�Δ�P��#Z�#>0�g!��P�霚0�+��ʼ��t-��j=JUHpk �cp����L�t�f�U� ��I.uz���-s�H�*ݐFR�	�CO�z��NI��!!�Ą�zd�bdd��~�|�$
�BV�ӎwz���c/��:c�HQ�Ɍ87�C�	�i����v�P 8ڐ$󯋀N�\����9j�9��32���)X�M�HaϧAt�=�F����1̻7r���&׉:9���#eؗQn(��I(5���@�G�@yܰfۮK�I�M�'J��g�mI���L�QҺ@����Gv���d:�f3b��mϺ}wb-���ɕt��HE{���"�M�r���:�a�/����RG/G�^,�&U�I@J�d˫<�(|�J��HoH�����0>yq�/H#
` ��M8e������U��db��t�Ƹ+�ߙUҩ@�.L)LX�O�pآ�e�ɹb�ŦH[ 5ѱN۳1��lq�G!D��Xƫ�V�R�"PE)�||
�@�g��5quj�kL��vQ[�*T�Wļ �QH,L9�엵l�t��#LT�m�����p<�鉪
�<�z� t1�@+t덈k�b�'�&R�m���L�RʓS�X�ցڹUF&m3�B�� ���)��$W�?�`����,<ئ�! /@753�'ڠ�Pπ�64b]��kG������ �dcC×&<����ʰ�
�1���0j�����].xǾ8�PO :a|�o��4¬Q��g
����e��c�D<���Np�T!Oe^Vda��E�0˾u�D+}�<�0���#C�}�pS�:�D���OzI��fҘzx���
>��:�퍁Ko>��a�WڦY�G��C~��F�[c��r�PL#� R�Mi����ϫ ��= �/�X��;��'C:�C��^�H=⧪�YZ&�ِ�S�>0L����Gw��0�E��<a�0-��:�Wr,�$m�O�����$W��ĘB,+$Xᑆ�x؝UA�8����>zU ��4jV�X��QńK�?�����06��)�hL+[��a�uıy�Tx��4�Ԩ��+9�O� �T�VŐ�CJ�%���D�L#�lY'��kZECTdh�X����r��H��eq��8H.�fnu��B��*c�a�BI;q���!��5$���N,Yt0�"�%m\�*���r������@`+�Qn�+Pax)�Z^� ����M7��j�&��;�����	?6�Kѫ .��<Y��k�JsX����&;�ԓg��cE�٤��
�>$jâY�	F�D:G��-H�V��k 2%�����'u\���ԃ�, "��D_+�pkR��D� b�	 Nt�'��!0��Z�D���#5CØjE�@��݁EG�Yt��=Q5<��pD�GW�A	J���I���ҙNV9�%���f��D�:p!z�sp*�g�6P��c��;gB����C��äN5����ᐹv,`��JI9d�8L���ފ
���Q�h �6@��/�	����b!��Ԭ^ZH�Q��6b̈��\gP�����A��Lkv,"9��q&���\_D�a��
7aʄ�S/��cJ�nZ�e0@@+� �،jF��|����G�7��Aa$i y1�� ��0 >�h􆖸 )�)t��(C�A`v��!@�4*�r�kM�ў(# ��@��pH↉^��|(`&�I�+���̀(7�����ə##f������؈4���QDK4dI^��E�D�$���x�o�:�0?�"���p�x�Z33f$L�_�O�%f�~,x1��.u �(sD�2g�OTy3jV�G�гE���
	�'�Z�:�bP=x�$��!����,D&�;p��2IZt�q*ؽ��O�|��O2��F�M��t��GS�D��OĬ���:����%�r�Xs���,���Á�;Q����A�D���ъ�$�18�`�	-]Ƞ�uMD��ayb���]��S�[
%z�i���e�T��ɤ���1���J�q��.�P�&8Q�R�@�eG92�D�0d+0�$�90�J�p�уAf�3��E�%Yq�V ��.۳CG�D��O����ݑf"O�;�Bɉ;&`�Q�
�'��H�5�10+�����6�E/gӂD�e�3?I�k���X��c�qڱI��z�<��G��flx��B�)�ީ3�̓�i|��K�FǸ)'n	���'� !��Ծrچ�S�ѿw+� Q	ۓH�=ڷ�E�!)����:i�"8���SpQ�xBwK�!�H=g����d�uG~�:儉O��4��)��%{�"~҃#�>,Ӱ1��
�f7Ԉ�B�f�<1QnSܪA��è$]Q`�œT!�DQ1�\@��OD�C)@Y#��
�!�>e;����CTn��3�թp�!�dVv�rt;�+�l �]�T&�#!��>!����fc
U���9��#B$!�ͫE<d%���A�JUS���
]9!�$^�Q�b VԈ1d>��ˤ0�!���Rg�Ϛ)� �Be
)��p�'�����Z��<M����'�"=;BN��8̙f@��°A�'���y�1i�n=A�A��r$	�'9�bDnL1)�֙I���M�0z�'��uW R\�h���=�D@��'�zP)J�0܈��	�B^ ���'˞�`�(ʞ��<ãDњ��'5��xp	��Q{���VB::5�� �'w0ђ#�d9VL�n�*�'��6f�D>�t3����ZJ�c�'�܁���ZD�qS2	�88�NE1
�'�b��`�{jD�Y�ϒ=�Zk
�'�llsa��|�(��F	T�5_���	�'g$�K0$؞+�"Q ��9*�Lm��'����T�&�t��h��t����'�� j���s<`ur�
Îa�iZ�'h���t����Xu�[�tc�2�'�0������s��:>[ƍh�'U@�k�AQs3��(TN���'U\t�UnI�	z��ɣ��+R;�d�'�L`{��Ik�T��bIݠSf�eQ�',�ũ�d[p4��e�JB`�
�'�ƌ0Ad_=nn:���iSL���B
�':�s��"�B�2���)
İ5�	�'K�!��Ou��Q��>5�� ��'D���R#�Pc4���%�P�<� f�s�D�:~�] 0F�%O�<s�"O�|Q��c��-ZrP�#zh�"O�`dC�5pab�K�6x��b"O�az��� c�\�YW�B'u�.���"O��:`�]Ot@�+\yM|
"O���E�m��4������ "O���c�#` 	R�rk��`�"OlDK�m�e��(�"ߋ`V䐳�"Or03V�N����!�RMP��"OV�el��!A�)@ ݖ:)�"O֤s���}��jn�%\"�s"O���7AȾ#��YR�`�w�F��""O�ah��ڎ]2T� '-Ӱْ�"O\�OәINh����<��%H�"O��В͓�w�ֽ(B	�T!�"O�a��i#!��'LI ),j�1�"OJDUH�gWy�s�ܯT �U��"O�! �W�3c���gb� �T�'"O�)�����AP�GM?h(4ؖ"O�D��_�T{��T�^�n����"Of�{w�R�gxzc��RF��"O
)�㓿o䥡��@W�\`"O��#�ۭsB<�셟A�}��"O6�j�͈�� �eM&Y��I��"O�a�M,Z��p�Fl]��B �"O�%����/At$�1'�0�\Qa"Ot��`iI�40� �Ѭ��uͼ�a�"O.MK�$ƃD|��`��5C��:�"OBD��C�?~�r7(ѧ7�p�"O���F�݉F:�X�g�QL�I�"O� �e��k"ܛ�(��u��g"O�E���G~b��U�Z o��;�"O�����pp�cZH�L�60�!�dl(��F��a���B��C�Z�!�䈚z} �c����!򥆂�5p!�F�qѸ��ǉ�N�8�z�M�q!��M���;�e?(d�Q����!��܋Q-������ *����)uA!��(;�:E��l Y�Y��捏K2!��ؓ7.@/	{:�(%Õ�<�v��	�'b�а@H"jC�l���5����ʓ5�<���O�/`D����-&abE��6�l��Ҥm� 2�m�@1d��T(�Hz�H�Qd�f�>v���9�����i�i5�I�6��L�ȓG�"���^�LC�L�d/F�L����ȱ"VE_�-^賄����������h��܁֞l�EZ7W�nU�ȓb7z��C�_���l�L �ȓX㶡���9]>�a��F�U�m�� �� I��-	VI�Q��#G�Q�ȓs�n왦��%H�����"�"܅ȓX�@\*ѥ�#���S
��
n����N�"��Q)D�>��@�`�`�4�ȓ�F���1p���p��V 4ЅȓB�P�kօ4g��	�VC�?`���ȓ=D���ޡt�m[g�~l\B�I?�^]R�`��]'`��D����C�	�����"<�r�Z��j�B䉃Spњ̈́�w�L�2�&�4���I-i�H k'�4�O ����ar|!!	ĳp��탦�'�F0+��߿iI�d�Y�dQR�>���rBZ�Zm!�BC�"��e��	j�m�A A�B<�Ozh�g�c��0铧-V�k��G�E�FM*�ߠC�6B�)� *��& V�}
�@USdp�f�)g�X�m���dC��(���x��P�*Q��<!�r">Q�@O�(��S�J[�'k0��3��R8 Xq����,纄����8���`C�^<��	?Q9q�C����9r2O�2(6��З>��A�-�"%�%ק�T�o���X���Q�ئA|�0����N���,Y:!!�
Q�@�q��N�br��Ԭœ�� eJD�v��@vG� H�D�q*�T�N�A��i��8)piي$<T� �6�[D-�6��p�Q�C5^�h������v��qhD)N���XV,Q�<��������Àa� )�C����QҀ�{����,X� }&Ls��Z�Bݖ5�ue�6	�.�{��#���!ԴX��	#Fˋ�iEZ�f] CD]�u(ۀ8� ��M�RI�h(��V� 0��Z|�C%dO��n��� P�� P�*KZl}��k�(ss<(�
X��L������
GS�S�� iūOQvA�q���vz0 �*�}.��⢈J�L]^��VC�!�D�

6�t�F�ͩ�:-��f��r�&���#�j�ƨ
1�R�ih�篂�?�|��L�� �6ƀ=w��.
�4E�a)7*��@���BE�!5�a|RE�)#�I�e�%&��B#��0J�9"�$�'2��D�L.5��cD TJ
-HR�"J)���CZ5A�b��PB�D��f�{wh�?�R�صc�la��X�~�(��8DT��D��-N(HC����a�Z�Bf��$ad8�v�@������ĩa�0��G�m� L�� ;�0<��k��;��(�2m0S"�wI�M����Jρ)�,<K�B�v�
��H)>�����2U/ 7MS 7�t1I�ΐ@�Iyb��d�^Y[�BT4|� 	�'��L�����
�[�GU�X�
�8r�y*MP�FyX%�  ��	�p��6M�!�G�("�I@>�@�����*=lI����v��b�'&�H��kE�)����SK�2��&AA����P�G>vL<M��.S�m�a1���	Yb�7$�M�(ɀ֡ؔF������>�1�ʽ �d\)���!��\�a��a�'t��AC
�$�rpq@����`ؑ�<�����=P>�(�`��\� �p��6)��{cK�ft�, �Pu����_��� � jQ�-��^�sߔ7m��Qg8"��9��C�nڱ?�tS���!Fۼ�#�>g���A7vDJ1�#b�-�DC���7���:�D��8 aB.Շ ސ81#��l�ve��(K�Q�FQPPmH�7ڮ��fhV$���[��юI��ʻm�|y��ȋ<�y7�U�V��B�M�[�Q���;�0?���]�K�6��e"NOY���慓Pݬ�Y�nY/����%ްLkR(��[0�����ΛLQ�1�D��Tֶ�!3^��x��J�zF�Y���B��SL;�*�D�91�]/zEh2���n7��ʒ��<;gZDY�'ێ[Ű�p�'Y��˃F�w������,�m�e (�	������ս6��tjE!�U)��'l�������X�F!�5W���I�6�Qʄ�d }#����`�{s��G�Azd��e����@M6�O.EK�Q�T�d����1$h�y�ҍ���ua�LǽY�P ;r�\$)�0y3a�S�r��u/Dq��w���)&O��Q��l$�X�.���2�'�`��$���g��9RT�+��h�����L��fꙡ@掁�҈H��4��f��-j��ٙ.���odj�����I� H�NIs�}��	�;�\{�����8�BEl��z�iػ����JH�/Y
�� _-q���;�I	��">�h@�|�����2�0�:u�T�'�
Oєs{�a*6AڥT��=�r��d	�a����u�ݯM.�mZQ���c.a���'��A9W$�)_�iH�)�)<x0�ҟ'Gʅʅ��c�<��s�R�z��}A���[�Ip���(>{4�'^�q�Юȟ\n��үH��8%�ȓl�J�!�a�,�+Cani�6J_�|iv�̱9�<�Q�W�n�N��o���E�L3����L�S��q9DY�������
uxJX���<�P�c�O��'v �Z�D	)s�`��lD9 �:=���(CF��j�(���J�R�	W��]C�e10'��+�$�*W4�">1�J�5oî�X�y��)j����y+��h49��b�!FG�u������HtN��I�.�p����{[T��E�8��I�#��x�g��I_�݁Q�
)�n�abk�}VN���eڞ<���0��+VG*_v`XB"ƴB�ɌN+�Th��"��W!�&���tBP\"�Ñ�|�������E�|W�D��089 D����Pv�ҕ�J�9��yz���l�����B�QM*���&O�820���˼��|cQ�J�'B�l�c��z�����ڲ(�Ď??&ՁW�7C�� a(=K�
BGK�l���=i�MP�j^�z�ꎑA�����=#�}���
#��1��c0�`U!Agƿ	�: ��8
�UP5X�D8b��H��a�f$j�@Ű1ov�0�L^�.�"@q����R0��u��Ie"`��;UaX<e��`�����Ą
�y�ȓT��y�	(Mo����Ee�@L
%`[�V8����[Z~�j@�0�|0!�	�50����P�
M�
tS.J*�8�QDE��5���pgd�,�0=��@��S_V��@� vZHp ��G��'"[�%@À����'��|I���� �t(h��L�60�	I�ቛ)�lҖ�Շ.�$P(ECݸ9wp�O \%�9:p~�� ��hT@A��lÄQ0Ё��W.� h���
O�8x1��%P��A��V S�@��@$J�(��D��V�(��i6bDڵM[Y���I������XѲ�����D�`@!�`��{�0�)U�%���╩�1x����1N%$�dR�BO�IB�y���>h]�<��ǎ ,����X�M�G-���dS�`U��aS)�6�ٓ"��>2� @q)��!��@�L�7tJ����'A�)(�=i���Eܫ)�L�i���fcL�k��)m���Z���:u1F���m\�,���$�̜egD#<��	g�(TӔOڦ4腰��Ym�	�Oo�S�Ŗ0]5�9Pl��e����P|�u�'`�h�P��� ]|ɚ$��&��y��M5��C����0>)���(|���"&FL�B�|-�rI��v��'Ȭeo��pD��/�ډЬW��yҦ�E�nl�;�yǉ�4s�p�ň*�t�,��x�ͦLL��Vሇ0@f�Ԋ�g�i� DUn�x#�i�V���L8M��R���	l��p �T�L"ޠ�d�H+\�yE$°� 1��,H\R��	`8:�Q�j��\����3��6k�*�s�e�.J �M�ڽ~>\��)�?7Wn��`��j��W���D�$�3E���O�MS���0��<�Mɛ��d�S�xbg����d9܎i�́�4�� ��-��H��m�b�0���f���QS�W%-��1�3e�E���!o��4�a|��?]9"��х��{�����;-yD����B�Z�E�Ǩ�=Ө��2��[4<��a�Zx�Y��M���y�+Ȍfk\� �f��XisD*�y�LϻW�4:��,HGN�R��s����!G��ڤE)��=I�l�:Q�3�lY
B��Sꔴk��i������2��*E�{DZ�דvƬjb�TtHE�'�O�
�:]��̧T�����`�%:M���69A�@2�lJ <Tba�	�,iG{��r�4�����'#���8p�[���'"����0qα�P�N;����h01k7!�KU��P�m��kY2H0B�`�4��$�Z����}���m'ue�0�'H
hA��K<�!�ۘ�K��ܒC�a���"c� %>Y��g��4�`f��	���9D�����jPZi�5�K�Fz�%�A�?�f����\j��1!�W�R�
b?�%��>�������GJ8yu�M��+�xH<i��ӎ)!�1R͌�ą��}���[D�-+�=Q�m�AH���i��wC0�?�E�JX�jU�W���Ĉh
)�kX�в�o�s>�=��dӲS�d@y�� ����DX[��2U�_�Ej��	�'qƠ�'��Eܤ�yU"�$��	rL>ie����-:�G|jix�-Z^�'%��5)��=P\��(E͌�OD�ą�]!��s�B�Aֆ�CD�Xrz9�e�H�T(P1T-��1E�&+N����	A��s��S�D ��U���,��B�I�ZLt��t�
H�P`��� ,�,E��$G9O񴹰�ņ��=a�cݍQ�:`���
�Z(7B�b؞Xq�!T*�NDK��'i��ELB*�P@ؠ���J���3�'�ri��@�(#��y��;���j���To���b�!G� �o��k��;u��B��:l栌��@20�(!���$oN$C䉔�hժ���UP(]�AJ��v7�B�	+k}�;���$n(SPf�Gq�B�	.~�,�Ѐ���X���.u2�C�IS벸I�*�m�M�si�/M�B�	�d����2��<#l0A�&� j�B�	�G5� r��� b�iCCCܢyѺC�	A�Z 
O\�ڑCqj�A�C�I�-�H2Bk�&?n��*5ŉ8V2�B䉱zX�I����~���(F=��B�	�|�@�w�	`��t+Da��C�	;֜�s핐q�=2�$��{B�C�ɖ�6��p)�yk�$*��@w�B�Ɋ?��QG*�5;�bXh���!�dB䉁'�hE1W@��~�|@�!�� p�2B�	�D����@���͋�e�8�<B䉼|�`��؛����f��A`XB��j��塳C�7N�&|�����4��B��(9$��O�0����d&K��y���;n���D8&�л�h��yR�ЭLֺ4#G�Ȗ&7S���y2��.��ip�oZo����y�*�!ڌA���G�pо�Q��!�y��!9T�
�cA8��1�j(�yB+Mp���Ѧ�,- (���)�y��E:(F��K���f)�E�"�y�g�+(a�	9�C��x��Gfͳ�yR��?,\Fh�*�<~�}3g��y"�m�<H�i�t�r�QB���y��=0�m0鞟a���ٱ�Y�y
� 4�!�jD�a��&E, &8�#"OdC����s�X� �U�S��er"O\��K[�+A2d�U��4$�DA��"Obu萩�%:�PQ�(�~�}�T"O�	y� �;�A�ZWxȁ�"O�����V1D	2E`�=!�^Ղ"OZh#+Ȉ��p�EnJ����p�'�^]���Ւ�"ЃZ�A�bR
�'(�q��-J�LP@n!;���	�'	��[Q4P"jpJ�L��^8��'G�i����=@Ӓ� Ǡ��G,tr�'F���B"o����,S��lX	�'��U�P��z���z�DX�E(b%��'�T �c�������*��{�'��\�b��nl�ܲ��Z"RE���'��2�^�R���	v�݃R���	�'M�񳏁-��9@f����9	�'t<�x���.�]�0�_�%� ��'�b�c�d�1Jf�;g���;fD��'@`��ÎV&'T�+A%Z�0'J�(	�';@���ʅ�~�0�CT�6�F<Z�'�.\�ԁL	p*��ej\1dX��'������F��=p"�@'3Ȉz
�'?D҆,��6S�����]9((H���'������Ug�s�A�/px�$X�'�@��wH��X�h�җB��tC�Tˉ��6�\����^_�v��g�[sLR�E�|A�O�LQ�,�4f�n��a �T(4�TX�l���7�'�u����a�bI�V�,;�e��YR-)!�>apG�	-��Ȇ�� ��8Qsƃg��ԢÁ�	:�'f>6m�#0�Xp0� c�O�Ҕ��gԐ.䤬�$�ڸ{x۳�	n~�D��	�ĩ�#��=ma�國eݪ��E�!ޕ#2�͝�~BE] .�Jy �\Yl�̅�x�}��[$%!"hz@IǖBכ��#0�p���M*ӧ��vu�RYJ4���9�V���a*2%��d����S�O]�N؉7	�� ����ʐK(#��p���	��#��0��OyR�����*i����ƂYD�%��թ��D��ŘUD�蟬��1�J�;�j	���,���'��O�6��azx��U�]0;�F\F�d�;#��l»9�x��j	xf�v��>u�Ip''U�B6Ti+�,ҧxg"���~��:�XH������(1-�4���+C�����ˊ�~�ÂNS�Oc���O��)� *U
x�)���&q�ҽ�a,ޢ	�P��g��y��+���4�?�}�P��U]�|bG#L�E��|#dߋ��E��x+D�K�Ot����ڢJO��iƄ��򒯍��8�fM�l//��|��O(�}���K����K��8U:D�&�F�@A���$�m���4�?����O��GP$����[.S.X������a	a(;:��&�"~���Q�P��sO�5q���#b�{/���.՞��'.��E�Ծ��a���e����WK$�*R�]F�	�K%�7�,�Z� 7����iQ�BY�+$2�┟<۲�Ų VJ`K<E�T	��@-p-�^��Ȱ	��~�K�8��:`�>��	_�pp\8qfeӻYzG�ϓq/��œgW4���O\�#���ǉx�`@N�a�
�,�:���ã� ��@aF�<�����Mʟ@0�����Ӷ%��e�V!�yWt����4HjhS�&h��Oh����:yҴ��ᄱl�ҡ�VnN�n1!���%l��a�΁�P�l���Y�p!�Ĝ�bt��٥�7x�TL�чݰ�!�dG8'����+_��P�� F�9B!���$�B�k�ŇZ�*3S����!�dӧ.Ev��5��X��u��9�!��%0��}��S�AL�F-Љ^a!�dKAzh[3�Ϣ��X�#���*.!򤈒�{���.1��=�w�R�_ !�W�/kJ�z�K^9~�v����I!��8��Y֬�29���ӑ�؁'!�䄳P+V�!�M8^�8ҍ
�X!��M��s��G�9��Q�tS!�D0V]+���d�t�wL�'!�� �� R�S�dJH� �+&�(h�E"OVa��-H�qZ�(5���L�` "O�����}R<p��/ƴX6�aG"O ��ԬӘJ�䝘��^@8P�"O�};��4��2Um?@��AJ�"O��r�h
�i2���l���*��"O&i�$��R��e�	�f���[q"O�����T<��X�^�y�|P(@"O������39�HP��B�:��}�"O�i�ت1`�dC�Cϓc�bI�s"O.8��D�\��0��{J�}��"OL�%�{�T�[�KC`"���"O��@dƪDFP  �.
"J+�"Ozh�E�>�Y��S�\�Dݢ�"O��b�7,|9�c��{��K�"O�8��)�2THH �28�f�I'"OTy�'MA�H�ҧ)�4��"O�!베�F�2���̹^� 8"�"O�mh�h��b(�8:R���~���Ч"OJ��ƀ�}-�u�t%֞f��I��"O�(5m@>֘���Q>�B$0�"Ora��%�Jh��2��}�8�"O�`�E`2M�q㵡�:mh]��"O�E$I�)&�ZuK�5#�J}Xu"Oİ	Z��0r�䌹_Ŵ(�"O��R�Lخ'�,yq����R!2"O���(_�)A�$ǌ�2�2"O:�1 �)$�a0�c��n�h�2"O�� ���20R�c�4-��E��"O4hq�"ɪN�$l��_&���
 "O��y��騠
D�\+R2�4JF"O�Y��n?,�z8(D�1d��!�1"O�<Hǂ�പ�B���T"O���3KrL0g�Z��H2$"O�k�i�e,�(��N&2��"O�
VC�;Q��ɱ��ԙ�*١�"O�ذkҢ�9�Q.�A�0�c'"ODu�d�^�5�l�0���:�X:V"O D�S`�{��`�����m�5"O�-Cg��-!���
[�
H�%�u"O�T0�F2_�nc�(�&K�Pt"OP��c��)������Y�+�%�2"O��鑧H<4�08СĚ��i"O�P�+�5���q���ʰr*O�A&N
���@+bJ��d��ݙ�'l%9�mE!6(D�I�o�(s�>Y��'�Lh�fY(
ҰL� �m��#
�'�T���kH�E����(6#Ĺi�'@X�1�^.�Ҽ�K�0xʈ�'o`
�_�*HѶ� / �0���'m��r�	�q�~02w�X�)w����'�8��i�\5��览���yH�'9ॡ�I�
QUl$�4oV+eX���''&�X或K�BE�	T�vX��'�VQGε����E���'&5��'|�<���K�/�2�+���_�=8�'�DCt(��
�����O"�k
�'�d�&'"P�K�������	�'�T��KA�b��t��v�ҩ��'�Y@Jĺv�4���8���'Б:aI�v���A��z� ��'eh�Hp 1������|�F�[�'2��HbaАA&<� pa�{`P��'�D`)s�)}$P�ʋ3rj�lI��� �:e!��n��"Έ4(�~ *�"Oh9�����d�ޕ�L�b"O��dO��D��C#q�>�"O� 93�K:����B�Ԝq��y�"O����&V�Y-P�R�"�yv"Op0��bM8U�=�1)ۼM����"Oz���K�/;��4y���T�Jl�"O�(�� '����Ǚ�ʢ�"OH���݃�R+Ff��"��c"O(,�"!�.	je+5�;=�`:V"O 4Ib�̚�RI�	��"O���F'Ms�J1Q�,l�N�""O��8�˅5r���d�r�mȠ"O�\�C1G�T�`���Xg��#"O�̊�ӵ�`䘲˛�:B~a`"O~ )���`$r�p�:O�.�1B"O�@���'"��gH�-����"OB�Ѧ�K��,K�AK�IoE�"OV��LW�P*����ϫ=X���"O��Eo�	x�u��F�Vx��#"O����S�S���[df�=g�\�
q"O�A�G�gq�b�+Z;&�X f"O"0�5S5���#j�0% ���"O�ܙ�B:2�Z��'O	߮��p"Oz�R�%���,�*Bg��7Ŧ��"OJLYeޛ*Y�rFV�v���@v"Of��P�\�}���XW%ɠK��5��"O)��%��D�E`W��%b��͚"ODh���� ��i֫�@�"h�5"O8䚂�@��@l� ��
����"O�]֤��V�l�GIQ#~z���"Oj�Y0M.�qhW�F!`z��B�"O�l�tǘ\���m_}nd�A"O��a3kƾ�J�k��ۅhҌ�"O��9���'�0���L�*x�PYط"O$ɰ�jW9\璌*^Qaĝ��!��J�`���
	����'�Z
o�!�$��Lf��>��bw�Z�&t!��8�f��SSm��eE��7�!�$M70˒ah���ag�<P��0t!�Dİ��P�T�8l[��ñ�2t!�$V 
����3�J�xF"P�F֓6!�$N�F0�d� ���N4Ry.9@�(C�'hJ�P%�7�2@���j�ݺ�'��EGҷ@92��B �[��T��'=p1��>{
}j�`� T}a�'�r|#�cJ(n�Q��̓F�H���'���
s�ԝ.��x�ʩ���a�'3@q�Td؇?S�K���:���'�\�Jv��]+D��c�l����'KV$P��SZ���K�	R]4��'�����m�D�~(a✂B/�\��'<HC�
�+��Q5��@T�#�'�0@�@���ul��t�N�v`�	�'@�Q$��7+$�
7D[��'�ʔ�3L�1���s鉳l���'�(F��Sf�]B�Қ8)�t��'�B��'#г+KX�8s�Ļ.쪩p�'���#@�S�X$�ʂ��4��E�
�'�&���&YD[
@*�K�~��#
�'��3v	ɒ��,��IU6E� !h�'�l��)��Q��A�lL8?;�z�'Ą󫞀_J$�0#"V�;V��*
�'?�x�&E�1$�6a��k�+6�d�	��� �Z`�ڇ
�^4[�;_YSU"O ���dG!"qJ�{�C�JN1@1"O�P7��"<&�+@h
%$�N��"ONͫ@���?�&�7%B�n�@u�b*O:5+&�[))��;#IF�f�Bl��'�*�q�J
��`ě2�5:�	�'4)�4�ǘ,`�!AQ",*���'J�=�D��=t6���(۵*5,$�'��P�&D �T�H�"Q�D�LqN�j�'r��!L�1?��u�p���<��q�'�8��F�&wKJ��Eϔ�0e�-��'&0�	��8���U+�&��̑	�'*P���Ɯ^<���edR(.�ꡫ�'qT��#�]F��8��1�0`�'����2�S0w����$������K�'�R9`oO:s� �2�˘X�,� 
�',zQF�;�����ɇ�O~��
�'�be9u*��FK��c�E�Ew>(i	�'���ꢣ���n%R�]7iK�pz�'S���~w��i�$�4@�t��'aF�� `��O���Y���� ��y¤	�8���o��
�(��D���y��΄Tr 1�S��9F�e��+P��y2`X	:&X@�e�.Rh���#�y" �"�Jc'@��l��n���y��6\��E	�@�� ���Χ�y�lAe����e/p��Q���,�yR�ή �D�@-=$ty�b��yrBͫ,���â��0	��[�,��y���L?$�qRN��y@��
B��y�e�$b�"�@S�t|<�W����y�� ?e�^�i�Je+X����	�y"�Bf�D��`��\�6 ����y�#ۂ���T?X9��eɀ$�y������4O�%CM����.Օ�yB�+#
2�aQ��%.��i�J��yB,�DʸX���+���B��,�y�K*)���2$ɡ-�&��Bg���y�.ه��l���ϸ&p^�r�`��yb������#��(�ty��+���yB,�%�)X�.LX(����yc���UȑE2BP�G�5�y+N'	�� ����i�t���ybN�z�z9Ѡ�0}fdY*�Ò
�y���D*�rs��_���'���y,͖Si���nΝK��� ��!�yb\9��u�Q6/0�-B*��y�¸`�ވ!1�E>,�H���yRMY��ؙs���Ot���P���y���Z`���ߣB�x@�Q���y�H)Dtj0�b�	8}�HQ�L=�y����FA#�.H�M�0�3'B��y�/ 	��L�'H���H d3�yAN�v�k5a�<�@�d���yrg)zb�`�Á3�~;�E)��O���H��!�4�?����M�ࠔ�`S�	���R�J8�K���Y�b�'��@R�=	G�`��8J ��� ӹd�R<�@א{sYbG����OT�"�̘n�Ɛ"��"z�B�ӿ�X ��H8Gk�p�An	������	�?D����̦�9�4�?�Zw���D�/l���** I!�'6"U�x��h���J�f���2�	/T�D����D7�S�4nڐ1�����YR��ܱ2>��jl	����/%�`�lZџ$&?��S}�"�D��#��iW�1���$$-���Y)	�zU�ug�J:L"A�ŴD�L5� +T^9���L	Ga@:ClZӆ�H�#�����\��$V�V z]��C�es4�s��l�:���L��̿r��	Z��MV�4���Km��	�|n��$ЦI�~��� �����h��m	Uċ�I��dXf�O����O�OP#=y*I�t���R��1nd��$��N�'�l7�Nަ�&���� �|��CU�n����҇�ia\���?A�����ۄ��?���?���?&�I^�	��l���(z������iZ,�����M5K�-�Z����?i����>�΁�h��4JZ�a�2	Rp�S�5\�����C�!"&������}���[_���C�n�>�hem�pR���{ח�,O�h�:��Ө�!	�GK�W�:��$�On�=E��I�"�4jP���
��D������'�(7���&�<�S�?Q�'M6�b�Ǚ�]�-u �&X��=Yn��-��'2�'�R�x�E��ϟD�	81ݸ$%�Ô0W*�J�3/6�cE��,�>̑1ΘG�6��
���h����f@rR��#O~��[ FF/>C
���K9@⼊���%1�L{��$�o�&-�#����� A�:�#D�j�)n���HO�Hnڦ&P���wq���&('��mBH>����?�O�OzH�aA=X"h`e���&`H&����M����6Gj��4����Bk�ݦ��	ɟ@m	Z������&���m_*5M$� ��?3Ĕ���?Y��Z�Vd���B��R� k02*$�];� p�!�)�f���R&�"?q2 � Vx��d���B�I��]04��Aȗ���L��X�A��ͲcoN��hO��e�'!.7��R�Ɍ; s�x�+��n�R�����}��8��ן,�?E��T%�(daS�X"QT|�f�5r����Œ�����")o(J���DA?���AhT�� �s�Jy"mތC�F6-�OԒ�j�I�>)�����n@z�!¡D��y
�ɍ���> nʜ�vJ��Q�2�bs̅#���{�����wrn��A�C'�8q���"Ut�جO��%��=��	�>� =�$�;!p,0C��J/-�a@�A�-bp05
������DC2wBqӘl՟�G���N.G��@�т�\��MJ��ݒ�����H�I���'���t@�?{�8�R)��yQ�H���O��	�$������G9~����ê~��Y1`U�j\z-��L��fX��fk 	  ��   �  X  �  s  �+  �5  �>  dJ  �R  �X  E_  �e  �k  r  Ux  �~  ل  �  c�  ��  �  1�  t�  ��  �  j�  ��  ��  )�  ��  &�  ~�  s�  � �	  �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���	N}�iÄz[�}�e�	D��Z��L�<ɖ*���H�a�I�n$����}�'t�'���	h�X3(��a#�ϼ)�4�"OFȐ�`YQ`ei���ls����.@��-�O��~������}��A�V�� �2�y2�
^�����0f ���y��';��ڗ@�C�<D��&�6(YX����� � y�S2Cy����ϒEEF0
b"OP�BG"ښw�i�cBU�@ ؔ"O��=Fy��_vH�"O����O/�8��#��B��"Oj�A���8 (X��Z�>8�R"O�@�%��51c"�-�%&�Q�?O��=E�d�J"��woF�aM�A�0���y�CL�j'����aR��1ZQ�����>�O�ᚱ �8|�r@�wGު<D���'�ɀz����� �,CV��
��C�	}�`����@����:��<r�NC�	�3%���<��/GVhJM��R(�mЇ(	�@9�g*���n n�\�������E9;��%�D��Y3���q�F��y�gB�h�*����J�XkaI�,�y�M���$X��>GP`i�l���yrG�2�B�@X 8%J9r�_=�y��Z�b��.�|pc�.��y�f^wX�ؐOې8��8�#���y�M�:Z��ڒ�0!&�L������y�E:i#Z�i���9a� �jr����yr�\<'�
��Da��}�D5�Z�y"F>�&苕�
�0�Q$���y"%�1*�2�(�H��C���cAN�y�蜍�%�, ��݋��9\B��3*�j}Q�ʘ� 4R��$ӱJ��B�	_�d�4k -c����c�ѱL@�C�ɕ4<�Q��%{��'�C��$9ހ�yRe�p�����BBB�ɩ!���N�B�Tճq/��B�I"#�d���b����/	:�a`"OF��'�P��>�{"i�E .A�"O�\3���������̩�Ppˤ"O�1��(�V��(IAKS��%(F"Oh�&Ya�Ё�0g�n� U"O�E������n=�Q��(&}R݇ȓ<�vh��KP5K14Uk@�H�p��ȓd`MM3�RA���9V�ȓlzh �f�4a�h������l�&U�ȓ�&]����m|�8PPe@$?��D�ȓ���*��&sZvͣ�ޙ1�&��ȓo�d0�M�������s���E|B��P�$Sf��!8JT)Q����2Ŷ��Ě8`:88 $����}{�hC�$U!�V�9&�!.�tބ$�f�$;N!�m5�P2��Il���G	))1���O��0D{���;�t���@�,���jc-O��y�`��r�88C�VnUdt���yb(	,�t�����iy4P�a����0?�-OpTc�G�U�X�[����;�d �'"O�paA!er
��n$(j�t`T"O:%�-xQ�uO�`p��"O�@0'V���
Z�cVv5{A"O^ c��$�Fa��NE���G"O��)$l�K�h ���R�X�"O�\k�`TC� ��p���H� ��"O����'Ѯ}����s���}+Dҷ"ON����: *�\����e��ɘa"O\$A�%�+mrF� j�	�e�V�y��חYT4�9eI;>�|$ce(F"�y"��6A�`q�F��3TTH�ᯄ<�yB%Ѳ��uX�+�0��YH�Þ,��9�S�O�~�st��P��)�B_��9��4�hO�>��IOJ`J�J
;���R��}�i�"O� $@�A��|�
�s��K1h��D��'��Io���d@a�ZhYpb־&��B�ɀ#Q`��3�nR��1� �/IhB�	�5W�d��@�Uˈ�*s��+M"C�I¦U�aHW�5e�5hP�@fh�!Ғ
2�I���<1�/�iEp��7�R?D�x�R���c�'��ي�/��5����b�����yj����D�����e+^�u���+<���I�<E�$M�-2�F�� ^Y�0��J��y"�T��UR᠛������ ��y�ĞH$N��P:U��[�,�,�y2h��`Gr��FȌ %Զ[���y�#�M�d�SÅ�n�vH��y��S#,��q�kӃ ��EM�2�?��'A<A�r��(N�Y�A�I*WJ2Ÿ���2���y�S�2H� x�A.Mol����T�1��C�	4,4�PCF�)8(^�ƌ��x��6���L9%�)�'�� {��*^[ޅ��E��t���B6��w&ǥ\.�و�A *��:H<�-O.��qOlp�a�#<Q��{B��?fS�k�"OrLy��(e�P�+ʄ>[H�9b%"O���΄�O�,�3�	��c8$M�A,1����O� ia�"P��bDj$f�X
�'-N������b�"��˖�й����M�+Or�S�O�NH�Z�8���=5�ٰ�"Oz�"���?]F��d�V�LuaA"O��`"Ήi��-$��<��U�"O<qjf�H66�(4r`�_�06j���͓��Px"��x�~x�"!B�q�X}�`F��y�cI"À��u��=@�������ybNK)?td��ݭ@|�di$����C���OFNLX���#��l{�	�<�X��'�6�Kq��5I���rH^�h�p�{�'�����%H���%uJt4�
�'z�1���2L����$�;7+YR�<�u��-�LR�n�7ki��$��J�<q`�!l�%)�4�3���I�<!��5�(�
��>�@eZI�<�� ���YǄ�(�����J�E�<Y5��'����@W(���&�ED�<��� H�H� �'T���~�<�ծ�����&	Ԧ3��ba�{�<aE\�+�jD	4��}��r�v�<�g�ʭp	�XF��4/d����k�<aĊOJ�VA����EB��Lk�<A���g��h��`��SIDj�<)e�n�y�Q�"w%�G�V[�<�v���.�Ye�tI�W�^a�<aց0E�t,��_>|$:׆�C�<�iՌ$�F�hƥ�z�%тbZW�<1��[k�h���Β`H@:F�Q�<9�#%��@0��^� .lA���c�<�	Q�$˞�B�F��G�hH����`�<��a�u��+qA�;m���l@D�<��س\��tC�Κ�6��\����B�<	���0<�Y:�B��Z_0��BmXC�<�ci2-�A��ıx ���CB�<qR ڝ]�p %A�l�L*dNG@�<��00��P�i��~մ�Z�E�P�<�.K�p��Yj�'L!-�IB5'^L�<�b����،��E!y�a��o�<� ��l��\�LCr 3���a�<A�,�!^U��b�;[���FKS�<!"�K7��a��']z�P��O�<� vM��A7X`�I�?ɈC�"On�06kG��� "�6�`���"O X1����� W�N�V!f��"O��ac\���=��E��}{zmR�"OF�B�@Zwm�=�u���^ŠȠ�'BV�\�I����Iȟ��������FQLm�Of��U��S�%�	П���ş��	�<��ş$�IП��I�.��p�ݤS�^��7ˏxT
!��ݟ���ş����������ӟ����v�,��5*çM.�XF��$�������H��ǟ,����|�I��@������I7}:ɱwB$n����������ߟ���˟����8�I� ��֟���]n��d��SV^�X�Ǒ�i�ށ����8��֟����\��Ɵ4�	ʟ��	�7�i�&! �P�sfק*�2��I�����۟h����쟈�I���ɺ'�+�ym`�he�w�B��OJ���O<�d�O���OL�d�O���OV��≍�]�8�j����xT�	�1 �O&�$�On���On���O��D�O��D�O:��֢�4��2VH�� �RY�U.�Ot�$�OB���OL���O����OF�d�Oh�dL���:��/G�Q�>���G�Oz��O�D�OZ��OV���O*��Ofr��#.fqb$.D 1��˴B�O^���O[oZ����ʟp��͟�	̟��b�ˠ�2]b��Ew$���G�ğ���������P�I�������M���?��$T舅b�A�I6�Yz�e
�[N�	Ɵܔ����������͠@x�4�1�џ<< F%dN-?���i~�O�9On�5�~mX3��'��te��6R�[�4�?s�O��]�'$����H�Hݦ���O�=k"~i8'$_(l�ѣ2��O˓�h�� I��7����a�<J��1@��ڦ9!C<�IS�'\��w��C�E��z�*`�[��L�$,j�2�l��<�O1���	��L�I��$G����@R>���AC�I�B���
�͓ѯ_����=�'�?�W��9`�Qg�$|��i�2C��<�+O�O��l�����yBb�%:�P��*^�=�6�8C�%�O��'��6����ϓ���Q�p:�ؚ����Xo���^�J��	?U�<����5��c>��"�V6��5�	�Rl�ً{#z�AE��.o��Ŕ'.���"~Γ}� �B7AM[a��2��(C6�ϓ`8�f(��������?�'4'�qاL5�:�#���D�6AΓ˛��u�"��G>e�ܙ�v���z�gM�k�й	񈃥=Z�d��D�]�|i�K��(\&�x�����'���'�2�'�A`���:h"��sHȹ,ľ���Y� �ٴgCu1���?����'�?I@IU�l���PE� R-ACmC%g��	��M�7�ia��4�埆����r�X)�A
�J���M1?�}jS�@#_��#��Xi�#v|�J>I+Obd
���@��wF��(�20��O`��OL���O��<q��i�@�97�'�P��Cc�Ђ�
�P)'�'��6�,�I��D�!�ٴ�?a���c�-#�I�>$ȹX��߲`��X�$��<Y��P)V=($.�{�̸<Q�'��f$S��}���rb����7oZJ���j޲K�px�`��7�&ݮ`D�5��
ٸ2B�p�b(	8�~�#V

j�A�š�(a�k����?��c�
��1��Ł BS�h:��C�<�J��t�� N4XB�G��i�Rt+(C0U��j!Ɔ.^k��z�F�(�T3���,��X
TOο[8�4���\�/�n��1K��J�̬�DaN2z�%�k�&�����LɱG ���c�Y�;�>D2�A�d�t��v��0�_�7W��ٴ�?����?	' H'g<�' �'�����8����UI��,��y� �%�OV$3�O$��O6�8Q�|��'e ��R�Θ�g�!ly������|z���_7��P5�b���S�F��,�Q�_��p�l<�	�����ٟ��'�`����E4�H�Q�O#'����g]�b�^O���O`�O�˓%�T�1a�P�j�l�Z�e�,H�슥m	U��?����?�.O�*K�|j�d��3Ŭ����+#�2��3�G}R�'���'��	��|�I	- ,�Y�$ i��̸&�2p�*º/p�5�'-�'*b_��T%^�ħ	H.%CIӒb�����S�rq�apV�i"b�|�\�$2cC4�S);� �JM1D����B)=�7M�O8���<�ҩי�O8���5ƍ�,@��Y��Q�j�����C·�M�-O0�$�ObL�6�i�O���i'���$fV~�^}Se���y�(pR�4��$Q27h�o�(����O����|~ҭ��a�~��6�G�MnAQTL���M����?�EF���?=�3�D@'����A�ڏv~�\4?���W>t��6-�O���O��)U�i>��b��I��@ 2�\�ޥ��4u&5�-OR��O���D�O�M���[!�떊��y�vh���Ʀ�����`�ə���H<�'�?���;`F)[r4�p	U�!��8��dS����O��$X	�1OD��O��D̏B򘉓H7N�Ȁ��OI��lZߟp�Eh����|���?)O�!0芰&ppa@&	�l�*%
����Y�ɭmvb�p���|�	ey�$Ԡ|D^�j�D=g�Dp�'�J	�mBǊ%��O����O�˓�?I��do<���V�(Ų�#@�G���[��G��?A��?����?ѕO�qߛ��� �T����D�]���5DX9Uz�6M�O���O��d�O�˓�?�Ec��|B�jǽhR�AQ �Y�%���8�����m�����۟p��>���� j�FIn�����6�� ���ph�9Ȭ�3��G��@�iu�''�]���I5xW��Sty��t�~�h�C,|�E����][� ���'u��'���7cx7��O��$�O�iӯ\��P�Jȳ|����:Om����'�r�؏����|��MC�`5b��a��B ��@��ɦ)�I��0�Q�T��M{���?1����'�?�C-�
!�@�B�
�4r��0�N2R�	՟�� ���	̟�ڐ�>����ؑ���%��{�e�<"h���i^��iq�2�$�Ot�D���	�O�d�Od��m�4�Z5k��F�~�z�S��˦�������Oy�O��O
���9��|��l�?@Y�	7E4rB6m�O��D�O�IVϟȦ��I̟`��ٟ��i���Tj�d>�R�H�3a�4{'Lc�F�ġ<����<�O�'�Bj	.��y�r�ۭ
����Ɍq�p7��Opr�a�����	П���؟�3��~�IZ<�@�1�ˬ�r��R9�P7m���$q�7O ���O
���O��$�|�fƽvt` ��,�T��|q�(�w�H��p�i2��'���'��'����O4mH�g��gC7�,([@��l�rupS;O4���O*���O���6�+�Ǧ� R*־.�flZ���Y)��TD���Ms���?9���?������Of9��5��u)�Ƃ�{�o��V�@)K���}��,H��'.R�'����0(g�B���O|,p�"R��ܰH�.��x��"R�F�����ߟ���cyZƛ6��>����'4�DS�l���CaK�SFN�zD̜z����'fr�'�)Q#h1b7-�O^���OZ�)��wcД���G�� ��Үz�D�mZڟ(�'���L�����']�i>7MD�I�6�bf��!��y�H_��&�'��G�70$7��O4���O����������I��e:�<F�:i��\;��)�'����'�R�|�O��'Y"ԳԤƞrxU�͝���l�����4�?1���?A������?Q��� ���"�D�P���
U�4l��+e�i}�I��'\��'Z����O��O��t�E�?@4D ���| +���
2�7�Od���OLT�Q��E�	����џ��iݱq����(�('G`�Lq� ʓ�q�4�
�<�O����'���ϋ&$z�`?8�0�1�oB"W��6��O��Z��Ʀ��	֟���٨�N���Uȝ4�?ssT��%:^[��^���'Z"�'���'Q�ӑw�<��Fkj�$1iD@i�~X:�����M���?a���?��]?�'��݇@� `�P�h�J���c6��y�Ȗ'	��'T2�'��k�6��FH�@!��A�.e�U�ҹv�<�o����������矴�'��l^-�����	�d�� N;m�6���W�L4�7-�O����O���<�e߲(��Sϟ��AOO'���D�Q�L��`:��8�M�����$�O����O�Y�:O8������_,%Zx;�
��n����c����O^˓.��1�_?��	������~��yd�5*�����#�7��8�O����O���,+X�Ļ|1/ʭ����(B�:͖ 	֬�����M-O�<Ҡ���1魟D�dៀ��'D��X1(Ls��i �_�s��9��4�?���En�����䓷�O��d��$Y9���`� B� �%��4(�`�P�i>B�'J��O�lO�����ݛC��.@�`{�옺=1�l�Ty�I@�)�'�?�u/B�;v���a�<s�N�YŇW�?���'U"�'�f�p"���OL�Ĳ�$�w�Q�p�RE]�h�1R+lӬ�O�8�҃VX�ԟ���|rq�9OFŘ�.�O�h\ *K릡��3 ��O<y��?	I>��t����0*�4g�\�3)�*Ʈ	�'�:tx�'���՟���ٟ�'^���BG6�
�YQ�Ũ"�&��G�f�rO����O��O����OH�z�*��#�.�텊j�8�cD�$��$�<����?1�����3z+���'@�bp���o��%h�O׺vv��'�'��'�'��);�'08����\?[|B�+�	J���5w�>���?q����;s��L%>�+��H�>��e)�A�:ֲ��W��9�M������?���y5>�Γ��
���Y4�L]� ����A��46M�OB���<QU�/܉O.b�O���)v	H  ��	]���3� �$�O��£�,��$�T?���Y��Ia����@�>s��j���C��@ñi����?Q��M���	��abf+�mz�)3w �=�f7��On���V��;��)]o݄��A�+(�2���V9<���L×3�06M�O��d�Op�I�F�Iޟd�&�y� ��"ꉚ]0���l��M����2�?iK>E��'s�	T�җ]v��d�/<#�q�jqӌ���O`��0�� &����͟�L���L�!Cc�8����8�m�X�I�!�tjK|���?��0�4����n�i�P.(4�UB0�i�����e��O&��O��OkK:4�p�VBX��lP�ϼ@���&	��	[y��'�"�'m�	�(޸� ��Q�\A���DضHbd�Y��ē�?�����?���p��Iy���8������>N�c�]�?�+O|�R)��L��� �'{m6@�c폮8t��f�0�.��ȓ@B��������-W�؂XZ�I�=1v,�,/بR�,*�X��/��P�:�B�&/�@PS##�,4�����"h�y&�>?&*]!��4�-A�[�]��0�%�
\V�! ��	l�u8��$N���D�i�Q��+7�A��K�A�T��Ս�V�x�� S�L�V��W��[��]�FH�1:Z���g�ȟ(��"��D�n0P�fעJ�pɑ
��X�	s ��k��D�&Ū��7ĭ�ʧ��ĸ~6��� ӄ	�]�ҋU��/|V��$�-ǄE$!�g�? E�ߒ�@w
�IY�!y��>����DX�43���'��� ����4��KB#W,ޢ�`�$�O����ʪ`�(s�e ;
�kblс]ax��&ړb�]p�LE
=h�[�K�(�#��Qş�������kH�|�i����Iٟ�+^w�6��s�橊p�ʏQ8R0�2a�:�yt��O*xiR81��'>�"R U�*��H*��
.w*H��F8"`���1O�On-A1 �����_ 0� �#y5 L"�͎�e��9�M°i���C����,OP����X��f{�@З�H��C�ɡRY2C'�åf=��!��I�{6���񟠑���������<A��`�Xu�e�ɎIj����3|���)�$��?���?A��d��O�>�[4�/k�=(�`�$^Gx��Xm��L��"V�BGlɃ�B�(���6�#�Aײ@��Տ"W��U�{o%�!�Z�r�Ai�8I<�}��F��&�J�ad��w��<YT�${�Ա��HS���A.р?-@���ן@D{2��\36=��o���A �a�=�a|�|�һ-$N��+V�I�J��1b����'<�7M�O��c��`���i(��'�6���Zc Y�0J�rhz��':�ܒ
���'��)þl���|�/L�h�%Q�F��~�6��a��*�p<�d��B�s`�D��*	�5"%��2:�̭��������L�k$�x1PR�`v �rW!+qx~C�I��*R"	S �I�/�F�jC����M�Tm��ea�p����^��#$ �k̓F´J4�i�r�'��GD]��wp�����D3#C��'/X��0��	�t��"�H�E���ApR���S�_>���b�\�"�m@n�1A;}r��,�<!��6L��9amW�\䱟6Ճw	X��7�Q�#�� ם>i�o����8ٴ1�O��O����2FO�z����B�Z�c�yR�'��y��W31EH�R` �?����d�C&Nў擮�HO�-�#oC�>��8Ч�F�����%��y��ȟ��ɕ3�|ا��ş��I՟����y[��6,���K�B�v������dl��G! X�pc ��Y�|'?c�H��� �~I���#�e"Ꭼr�����	���{G�>2"�>�O�@p�_�p�Na�qJ�)R���㲁�O��l韰8Uj���>˓�?�J�w��q㬏&j˾�1wҩ���/�S�O� =*��K{DȺ�o	bռ4+�O�lZ��M�N>I+��ʓ^Ă̙��$��|��c�56����_q�(���?���?�ſ��D�O��O_���3e�-F�bL��J�?��Z�ēsEcU�?�d�XP��x�'�x"aF+޸���T+���ؔ��2~�Dȁ��/5�!� �Bt�џ���ɓQ(1�Ɣ%��ݸ��N��DU����4��'�b?�i�$X�e���`4i�y�|�K�J(D�@��V�E�>��P�l�@B7H'扭���<Rꃾ]'�F�'?£�/��ǀ�:>zi��E2��'�()�#�'P�6�H)����

^���P�)%�|�#�T*aVdjB��
$�p�v��K�9G~Rf�zΔ�����5	��7V�\�����5vR��`,�i~	P$,I&��0a˩?���t����O�hl��M�2i�E �IA�;�-C��,NydAj+O2�$*�)§���f�#O�&j儂"�����bn�����<�C!c^�u)#�?�-OZ�Y�ʓ�e�I��O?V�	d�'��I�fe�;��Y�B��07�� �c�'6��U6�{����|�؆�q�z�'��V$M����B9kY���7埮Q:�R�xp�$i�"i�4\���#�����!�כ�~�)���P�<�!UN�d9R��bc�plm�ǟ��O8�S�,�ԛv�\l�xa�FƄ�Tilb���	fx�d�)�BR.=8\�RR:'��!�ቾ�M�Q�iI�'�`�{s�P�h�.�j�.p �`1,�>����?bINX�����?���?q�;\N̫��1�J,:��Y-G_�=p�〮M�В����H����\���O\7���<Yc��r�lu����הY`I�  X�Xmڻo!>�i�X�K�R1YSO�K���Td��3&2��r%��@P�� K;<�ZR �O4�ux��i>���g���3�dR
$�b����_[r8�v*��E/��/��;b~=Γ�?���"�M����d�=�&}+r/�>xl��'�=T!���/g,��$��W.T�t� ��!���n�u��$fZTQ#hCG�!� ;�2��pn�@;�0"�FW�$!�$�9M<,�Y��ە�y�C��-c�!�$ƅS�.Ȳ0
�T> ��)^"�!�Y�*��rӯćSݚ`!k��!�$ӪO&6@���)�`%� J�p�!��̀8�T��	��5�A)Q�9�!�� քi���8�����O	.`i�ҥ"O�y9�-�"[L2A���f2�"O���L��f���c����	�"OtuK7G=t*�$9�ƈ�t����"O�3���b��䒍a�6qj`"O0�h���+T�3�ɇ6LȾ�xg"O ����	�!(Vyj�iC��*��!"O$�:b�υw�x�*�9��u"O�Są�%���q�PG�z���"O.�@PI3+b�,#S�r�*��"O�,ҡ�� ��(s�+� ����"O��d�N |�KD��#?9ژZ"Oʐ� "�1?~���C� _�T��"O�����C�֐�.ŸH|<[�"O2
��=Aw�ܹ�O@9P�yr"O ��$-��0Yu-[2`'� �"O*��޶u��Uc��H�A.��P"Ot*���� �z�� H�
���"ON<��F�'��|�.����q�d"O(i���C����A�敆Jج��&�O�\(�e-�)�'Z+@ H!f�?i���:& �Y�-�ȓ&��QC�� �H�I'��T3�a�Oޱ�N?lO��1�b��(���Tn�r�b�'.�d`Vϐ*��{u���1��DigX$�Rd�ER����� -Y-�Q��Ċ�<�b�)��3�^�Eࡣ�U�%YD��A_��pu	7��h��+�mS{�<��	غ7ǴX��
}q<p!k����y�D��J$ ӛ'2V\�ٴ1���i�19��F�O�/#v�F��#�C䉐F���p�!+ݚ��#ʊ>a�^	k��� H��9�R�x�DX�#���ɀ�.MZ�'�XЇFҦ}X��q�C��8ã�>�O��SWǒt��­^��Ǉ�$��tSP.Lh�@�J�!�l9f [WX���a%�r�+_���`��d�Q���4��2 9ܔ�VE���hJ��O��ã�1c�.���8&���8�NQH<)R�^�W1��t�M2Cze�C�T?�E���{�#�>g�+c��K?�~*�������9'(����1s��w�<�g�T�Q��Y�d�qfN�[Ei�>�N��!�u?1w�

��Q�6�K>Q�I�2�nD኷BÞ��`GT���Z�+��J���H#~@��N��f��H1ᎅ�4�T�'��ȰQ��,��ëre�=�bA"c.n��SH.��tzQ��'�,iA`��-�
��k�耦h�~'�= Ŷ�F9�>�ɖ\\F;��.��O�\���y��`J��t��5O�pS�o�0���ص)_�(��]���>��m͓V=,��FŮ4C��s0�H+)���h���@�a��Y�Wޖ��/X")�@�"�I�Yɚ$z�eɈ�䓙yZ���)���̻{�L}
�j�.��DS��<eh|��	%�|�c�ćy�TQ�/�(�$�㴊����I5�yR�'+����.O:�jHZ�ak��p�d�pS2m�1MB|��
 �0M�eGz�$�8�(���f���x]���Đ�;�B�6��$t��+�rE�$Ա,#XI@#��!a>r�+S̀�{I��Jc%�WM��81�8��"�tӬ:�Y2Q��T�'��u�d�8��	�;��$�0OI�L=���ecѬ]���XOs�����^;�MD�-	|��4��-�|�+1�����d
n�nW75��z��
!QhD���8oba}ҩ�1^���宖@�d����%uO���S&d�~#>��Q�,5V0���Y�a��xȀ���<9��ݖEjzq��_~����M�'�v�ٶ@]c΢�;���7CY���uj��msҐ�U�]�8���2	{d5�'%��Bԁ�/р(��OF�`�ґЉ���F�r]���@9/H� ��"�H�B$�KM��l�j����Ѓ�;D�\����1~W�tۣ*ƭLY��y��T�y��m��.�T�nZ6$����,Y��a9�ň7>���Ę9(��Q��3x"�g)�i�y!��I��?)&h�C���Ĉ� .3�a}�IL&�T�R�/�w���Zb��&9�p�*R�;i�P�O�+P�
k�y8�)T�)+P�s3BI�66𽻓�!����K�+S(#=�F�];[x��KB��4t�qЭ۵ITZ���� �~�5��\�kB���L�3%�`�<�D�e��a�	O�+�D;�.�k�.~'^Ւ£����ǆ5L��6�ԋ�x�J@ {�ٲ�!B5|ν�#�_!�1O�.'HB��R��'a�U��D3/P�Pr�,D�lp�y�M%.��1��Ih�X�x7�Q�Q�ĕ�S.I��Ń��T���WNT����'@X�z3���O� �	�b�x����K�Qk��y8��@����j&e'�x����H%{T�Gm���2����#�
�D�*�!�|"��O*�#���5��Z�P�!� ł4��P��蟀�HOAM��i�:O�m rCYT�d�V�p"ĝ�qH5y�l�Ef�1A���Ol�An���	#J̙\TQ�C�x�˓U�YDi'"v<D�w���M{�b� k (��@̞�<9�	G�Ck����?��瞯G`t������&��v
Y#���b����T�L�-�M"d��bp(�����F�O�v�q��M�`yt�x����g�NT��(�On$�
}1���2�0B�E�
0\���"�����	��!B��Da��:�䘃p�$�0͕�,LR�8ڴǚq�i��Lr'!�����V0J�m�I����X��5��Q��}���Q<4�d�m�HO0ijpG�2c����P�@مM[��ļ"H^�.�~��u�X�nн;������V�ܡys�UŦ�S���svb�X�5��Ԭ�E�M|�|qb�fx�4���5޶�1�Q�X�1��a�T��~�>���'*bP%�a�8|��kՎpY(3%��F՛&�O�t��ۓqF���7:7vĒ#A�[�f �p��x�qgO<�~2�c��ԟ�I�u�G�<6����7�,�#����?�D��&#�$�%�0 Ľ���	�D~�L���i7�@�p�<@��O�����ļ����$��%���5K����@�1� �	VE*��OR�m�%���@����
�v�Q	����Q90C�� �0�c+Of0B��,E��	�{�nU����'Ȭ1s�z���(g�H������u�.�"GB�Rel�-1�D
X�dZ�E5G�P���\8{��у�O蠐��'˖��������0�مx��a �'�i�5h�-sj�\�C�	&rK����O�s��h�>I��`��m�2\%R���X�<�e�W�Ejd�;�ḻPv�@iÏvxuY�N�[���?7�Og��;2�.?�(lΓn�R53�
ͦ?���j�G=�>��;��Mᐢ��i�x(sv!��p���*��77B�U��'����R�>yq'LK�i x)���0~�O� �Q�v�Q�k��zz��ZR�I�E��b��]��X㧎�y=��	U�~pz�d�4q�>`����E�FS���GΖI#����=Y�nM�nZ���ɤY���'�S���˓�]+6�!�0#�0Az�}H��ͺ�HOk̘����I�2����  {�!����� �MȽ\>��gfA+T2�듭HO�lv'�/:���[��,4Jy(�-�#W(^���,2F)(��L�k�'^���O�4ɀ�A*
��-��N8�B�,�Xb���$�N���D�K�)�A��l�D�T��H��aC<�Ia�$Q�h"!��۴f�;0q��fP2%�`����F�O,}B,4N|���*Ơ��R�9��8�T��qX���FhJ���W�#�� �R�̲/O](�P 8%�'����r��
ЩF�pYx�:�CRp�Շ������w�ٟTAG	Oަ�hЃ�7z���2�O+,O�LQը�/t蜉a���
��)#�şrN��ٵC�1;��L��l�X�'P�LG$�ad�7m�.F�Q�7���0OI�pih��P�ӟA�tA �:}©؇��H#��(�&���'�0�!aJ�JZ�y� ߫Uz�����]��E� �e��y�BR�0���'�^b���W�MA��Q���Z�cu�,=U���L:5�*Ɇ�IWp$����N�z3l��&b�#uW����ݐ9�xZcKD�XV��U:���4IB�s����vg�I�?O�9@�HR.*��)b��T8DZaO�#d��P�@MX1SŶ���)�*�y�"պ���N��L�P�`F���HO�Z�b�a��+&d����tؒ�@3bu�HE4/��ťO��� �6(�zP����N��jB�$�+%_�T����'�ؠ�c��\Qr�P��Y<��'��	<5�@�C���>9���;�xB��]q� "�GP�	��`�熑$�����<|O�Ab���$����6f�Rc��j�il��)�v,#1Nϊf��@�Ϙ�uG�Cb��P`��'�0"����=��L��B�DQ �4 Vł&��R,V�	0 �u�8��F�X,(R|<"�j%ړU�JBlMc��9�w���� 2'W<U��H*a
�I�}��Q�B�R�7���pH�]�ش�M�{y�+�rj�{�J�Q!�Tc4�8u�bOBI��`
�1jv�B�H^�>Q�0�DܽX�l�dAC�`�p��n�܉��ցVU3�V*���}��j5��0<L`��!�N� ���������Yr�P� �]�� ���6b�3����+ɂ�� ���d�O�6��c�)��k�v����0,��� &ֈ1���DS5W���5�,Wv�h@`���%o�f����a�ܸ��''|13�?�3D�	P�S 4�8����"U�t��K*o��T	���bՂx�tl�oT����n)�'��I��
�H7\L��D��7����"������:_�N=�`]ᖫi�1O�i�����M�����L��a�!&�6L�HH�� ��~"��e�f~�`>c��Kw�(�#�/�E�n�IC"_�4(����\By"mR�&LO��7�I<1��"��U�s��i�w����ɔ-�l �O��R��m�O�,E���]vPi&eR)
d�'�J� �3�`]� �q�"�0>��j24!V
� F�<�/O
�^?���G�Q���O\�I#��̡RG�t�V�S�'C*qF�C~���G��i��O*�1d���ne�I��-J�e�����1���R>O��[��;��Oc$��}�N�@q�Q2�ӭvL]{G'�).�
	'� �(��ĕ7���]�y*��i>"�ٳ��С�#ͰgŪ��0�C b�<YT�=z��y
ۓ*J@P+�6v��CR�1N %�桚2P�J�!�4zi��θ<�����Tk�Q?�ݪm�t�R,�s���X<MO��$��/F�hx�`E�v��Z�	�}�4Р1B�x5�d˃_��q�����O���Q�뮖�,�� �b�"�~�b'�\�U��cV�!.��<����b~�`#�L�?�a��?)�4�h,0���0<_��ے�R:f<��'��iy�-�4Lxe9��EFr4��D��z��q���בvf&!�r'I�lg4���"�xzkcnk�����4�(O�i�S�#V�E�Я/��]�4F��SA�DZ4j�
�
���G-�O4����Y�e�DI0`܁H�*:�K�<,Ϝ�Fz���3�Z�u�M�r�ٸs���*3�Q��'�U���"m- �&�F	�
M��(�D�p@p�k�7��$A\~�E��Z� 5(0�z�K$9��R���C��-���t�@�%
0Dy�����A�	�R���p�P�?��R�D���B�-Q�Tʑ��5���!@��>��]�-[�\��Xa�C�}�'fL��M̤ !���7�Z���4<a���(� 7=r���F�~?��9�uGȖ?&�0�V�E2O��h���T�Zl�a��'o���hI�zw�b�`O?Qz<��.��<�s_����O|$X�U>���^�x�]�%p��`1i��,����F�3�FB�$Vf�1J!ل2�� ��S�iJxH`a��D��L*���y��7�%��?��HԁZ�+���1�iLRp���Ɠ_�� N�)y��V�G�9�� �شZD��;�(�<\*��2�J8d�:UG~����tࢂŝ�0�`�*G�ݓ�0>��EBo�%��hH#7���h䩙� ���6I�4r�r�q ��a�EQ�D����6,�#�A'�Ȼ�(O��m���M#���Ц�M~rpbA�[7rD�B]�y��Ͱq`�C�<�e	@����f<o�E"W�<!�Ű1���aƭ	�0�e��Q�<ْn�[���a�@�@��xf�]I�<��"�0P ��ˮ]�<}��OE�<A 0d��2c@�1����u��l�<�ԍ�Z����;87j��Y}�<��JY��Y[F蛺	�X�cƉ�~�<�MȀ3��1�c��]B6�'L�U�<i�*7#?�Qْ�]0clp�����O�<1gE��|��d�hF�w!�Q[��C�<a�\,��4�B��R.���2�K{�<!&��U����UN<$�@�@�<I�@��#%����OH�������r�<�`�M�xT؉���hlT8s��m�<iSL��zR�Y���e]��:�!�17��a���D�Y��=@�d\=�!���Rp�T�FӔ�b�a
N�!�ā�M�t#V�� R��oB�%%�B�	�!�~$�qA��^��!D�,C�4"4� B��"=Xiq��Bz8
C�	�GCva��Ν;,�y�L�N`�B�ɠ,q@���l�XI����pC�I<H{�ٛ�QC<JIQ񦟟m�NC��1X�b���P�V�P�ȱH�F�C�	������JI�EjB�XS��2|�C��vtY�$�ſ	�T,�TOY�5�hC䉫L�h�&��3�p��P��:u2�B����e8�C��tH\E��[%(C�IJ�4�F�oz襈�����B��;c����p���t� 5��j[RB�4x,{�:��������T�0B�I���]#T�*�ؘQ��4`�bB��no����B8�d,{�`�7aHB�I�h�ܹa%�%.���5eV�6!pC䉘X�A�����9@LSUC�I�'>tA��J�5Vx���C�)� X�8a�%��SA�-I�F�R�"OxM�W�ެ�\\@䅏%]368r"O��5"� '�Q��&:S�=X�"O"-��j�XM0a��ąc4�i2"OR)Z�-���(�#Q�R-�!{"O8�3�e�N2���h��;����"O�x��l�I�����9h��\"O��ҍ�SV�Z��	���@�"OH4µ�K�U�؉�����9�C"O�` I$�Hs��/`�*X�"O��u��^eB<� �����d"Ol@�b	{<����Q�@�"O��2���ũ�&ʬq��-ځ"O�����H�m��HB�T@@Hf"Oڭˀ��2�P��ŀ=I&��X�"O"�*�X?m{�c�唋'�>���"O��q��Ƴ$�L]"CO�q"DҐ"O,pr ^����gKÇSW$ԩ"OQ�q�K&�U�C��Q��!v"Or��O�=ӞMA�
ܟI�5Y�"O���H�{�b���KW�
Hq"Od�B�P�M�x-��	��֐�"OT���F�?v�	��IGb��"O$z��щ iB������P��"O��S�@X/*鼌j�H�?F�XD�"O�qRP�_�΁ �ϛB�*�PB"O�!�oکAt��Ơ��,����U"OR�#e*Q�̝(�F���li �"O���/ŽW��<A�T"���"O~y�J/Bz2��l�"o�Z4I�"O���_Ǌ��F���"U�\��"O�ٖl[?AX�:�
�?LR�C"O���BE�e�pd\'l�����"OZe���Ƀ,B���U�փ�e"O�9Ea^�,F6P�%.�1�^��"O�-�2���� Z�L�2<RA "Oz\Y���?V�`��F�-,��Ғ"O~�@Oдur�p���� ��a�"Op9Q.dg|qѕ���(�*���"OzY��a�� �>$�r�#ue�""O��UjE�S+J�4 �p]x!��"O��:��ٜ^��0���0N�!�Q"OdX � �E�R�{P�C�*�	j�"ORX�@��=�I��-ZD�T��"O�]�CNڭ!J-���S
:�+�"O��@�̩,T w���X(�"O��3�E-9�U�*ԏja��P"OR1+�X5[��yzk��E��P"O��{4�&^��x�C�_�^a)D"OF�شf�;g.,�v�&Q8�\`P"OH����H:J�!:��6B�+r"O�����ʱi�%:5GK�t�PR��E{���!��̔�u>�h�b�Pn!�$_ePtq�ƭ,B�Xy9o�O�!�d�6MT��[�j�[�������A�!�D?'�t���\�gw��jm��i�!�]Kp ��VB�UcZ�a �i�!�[�"m cr�J8F�t��I�~(!��"0��Ye²�*��R*U�~2�|x" �,P
`l���ӱ^B�i�!�D+�yG����u�\W��a���y�'M�B/N�@� G(J]6�d���yRȀ�X����dJ�/���'D%�yR�I1C��1��(Ym�(!��L�y
� ���(B,)x�C�%�P
�"OĤ��Q0��ı�H��w��)�"OpB-	�2D�2-��pi��"O�@���(`����k�8�"O�Hq!�˸Gʐ�k���34��e"O�p�ANQ!8�F��@�
��"OD�)!�J<��:�Aܸ���!"O��*�I��!
�@Uc�r�a7"O�MCP�N�Z_n�òoD�5�r�P"O>�3,�R�X&Ν�r��AS�"Oƀ��g�9M�C
�,'~����"O�;G��z�*�����3C p��"O�����Ԙ-r<��Ϟ�_�!Re"O<����5Ӡ\�u�:t����""O��1#c�X&����e� �V"O��y�"�f�t�2#�;��ݣ�"O 9[�ț_⥠# ��9~�mX�"O.����@1F�:�+*̛kBF"OJ ��nߣV��00��'m�0�8$"Odp;�g�^E���!�	��0�"Oʰ���C�"��hq�¤	MX��"O�pS*ǀo��\" �cᆱ��"Op�{�o�-�j�!�AO+q^1p"O�0�FHm���ꇡ\$>�z���"Of�x6��6D�������K�H� "O��"���uq~թ���>��-Z�"O� :UB�{
�9���%-��}*"O�h��hV*��$����R��]"ORUz����Z?j��Q��3���E"O��I��ܮmΤ��e^��zm�'"O�I�*
�x%�U$ͻ����"O@�g��"M|��r�9r���2�"Oz����&8�<�A�U
��ɳ"O���#�G�u�T����(mB�S "O�P�'�,mXM��d	'[yx�Y4"O��C# �)�2�=c�؄Q3Z�E{��=5��D(5
�+m9p��O�o�!�X�XN�p�E�	0���g/��!�d� [L��W�ȅ/#�l�p'�
�a~b�H[?14 �18`(S�	j�R��M}�<y�C@:V����+P�k�ޕ9�/
N�<Y�Ě!9o� j���0���C�d�<��C�$�d�cF�4`xd$@Z�<I�
���zaI�R��P+X�<Q��b"�qf�Oc
��� �J�<	P�	r��U��'0��!��D�<���CQ�����m����8�vL�{�<QӍ�#Sf��x��9P�0�#_A�<a��C#V� m����%�~��e��b�<���5Hx.y��2rT�эJ[�<a�IP$"��tb�kD�9�zAr��Y�<9���)G;n@
C�X�$]<���V�<�wdM� ��=HS![�g��	���O�<��`E�H�Dc�ÂwY���_�!��I�}����7ϗ"'V� �-7:!�D�$�"�.��| ���jG�9�!��ͻ{J�E3䆄=D8��0��u�!��x�0뎤Q14ऍ�{�!��,��\zT˽<,0��B�8{!�D� B�f��H�JA�-M;�!�,�`�*�ǖ�>�`�b�l�!�Ľ#�I��IC1���N��!�Ğے�cgg�u�N�{p��K�!��O�hG@� �>���1&t:�"O� |ȉ4���U�J�bd�A !t�x"O�)	�FIlgVy� +��+��$�@"O�����ۻs���xd�KuB��t"O��J�q�z0��Ɍ�h^����OTh{eȵ�� 󄯎(bV��Q
;D��*���N���
��$˒t�g�<D�ؒ L�"��@3�/\�%C�Ha��$D�T9�	l���;�$�gP�� ��5D��Y�V36��YA�Ӝy�EK�?D���g��B��-�@��_�婴c<O
�=�u��1=+�Q� �c����s�Jq�<a䎓�&�������Me;�cVp�<�O:(�p؂�ՋP��d��(�o�<�Bؗ7R(x���Ucb�ţ$I�k�<�R�^� ��m
j�.Zz0B�f�j��\�'���Q�H/b�V���ˀ�lR�e��?	�(� �ރg��˂��4H;ʤDb�ӝJ4 �+�d۹�R���g��B�	3s"�XV��*$`�
��?t��B� o&h�$�'������ژOm2C��H���E9k�8KuI�:��B�Ijt`��D�&KG�Tb�I�B�I�^T�ó�M
<�)P$Z�{2�B�3Yd����*�\p>Msg�n�bB�I&��%㈻!�H�P���?�6B�ɱ���5��hU���&l@
T�B�ɼ��Hū_�	���n��!@zB�I�/O&�[5aL�h��]r�""{^B�I�pb�Q����8I����Σd0B�ɃTd�my�,I�?H԰��@ѽ&�B�Ʉu�)�ń<9�d��t@O�W�C�	�^	\ �Q	}�m�!H�4l�C�IX7�l�k#x%hGg�\��C�ɎO�Pij��[�e��I�C�f��C�X"xe�6.�)Q�ň���Q��C䉓W<*Y��<-A&}r��\�Z�C�I-&A��G8z�U�&�ne�C䉘�h�sUᕽu�<Y���nrC䉏"�\\bƀY��������5�����%#(8���p+��u�R�!�D�- ���"#�"H� �'۪x�!�H�f� �+c��8U \#�բ4�!��ɜ8����B�Iؔ���&S�!��]��)*gV,d�0Qs�r�<"O�F���#0И*S��y�a�nVh( ��)#�*��5���yb�0b+�X�ac�8���h��ԅ�!�>hʣh��R1V��VG� p��P��9(���&J�vY4��3�!n���"�|p* z��kA*����'���7
��Z�i`h�9 �iy�'kd�)�2Ԧ���nC!/�
�'�2�����0-��|W� �p �
�'�"�a��.vf�$�v�J�'B�	�'$}!CֱZ��m;�Èߢ�P�'2l�����;q�I�!v��'����oߪ.H��1'P�n/H��'���(�
5�u� ��`�0��'9�����퀒ofN�pUJ�8�y�*�:�*@2�N7a�
�Rf.��yB.�-��"���S���C����y���x�h��L�&7�B�a�N��y��G":�ܓ��U�Yl���J��yB'g��4��C�QU>�BWDK��y
� Θ"��_g8�.D���-8�"O,9{� � D��M&���pD"O�Pb˨D�(�"����e	e"O* �fL ^j���MO�0���"O��d�,l�\�ӂ)Ō�&"OtT&b�!8T\��Ó#Ţ�"O�놢D�/r�%��'̏x�Pث�"O��H�20f����&�9z�IE"OΤJ婋��B�(%枋H��9�R"O����BCakP�a�EHM��LB�"OH�t�)w�,����w���"O��{�?_�����l %Di8��""Oz���[�b1���{HC�"Oz�I�T�|�$��E��m^	b#"O��Y�+ع[|�4�EXc�Ti�"O\D�e�@�\���F�7�̫E"O�	i�a�]��-9�E���B3"O�a��kԨG�j�PQ�T;t
��*�"O^i�d[�4���ь�?T,���"O�)3�@�,�V��A�0��"O�t����#d�H,�1B�6p�+@"O$q�E��,�a2�ǅ����"O��rc���0OǻrBr�W"OB�$'�zƵ ���)^�\��"O<�r�	�0����\��@��"Ov��V�!O">u����Y�"O��� �#y�f]A �B�)�n��"O@��E� f� �UNQ�Ww��8�"O���t��6-Z~v|Ը�"O���N�7>D�QA�A!pjȑ��"O��j�D �	M*�����e��%"O�aAC�EP��)7C�#Q�z�(�"O���BW�� `��a���+"OD�ۂO�	�xqQ�J?�}8�"OZ�rB�A�, j�A���k�2i��"Oĕ���F��<��0d�H���"O�A0���h�D��C=l����V"O�K�����Rc�~�D�;�"O�a� ��/_=pЫ���0M�քu"O,�(�)��BIaK��W�x�l1"O�ɔV��� 2BͱE�&h��"O�L����Y��b��_�t�$���"OHP���Ȗ@�P!�"�	�ԭ��"OHu�ԝt�H1���V�E�~��"Ol�3g��Z�0�Y7��-e��h�"O�J��4$���@i8K�~YrT"O�Z���{O��Q�bN�Z����"O���r'_�>�Q��AE�T�b4��"O~�S�j�%��u���B��%�5"O\5���
u�� SD�@��� D"O XA��:�聧`K�m_8� �"O%Z�/Df� ��OGM��"Ol�J!�4q�*���Ǎ.����"O�E0�"Z�t���6-��|,����"O�xst� �K�~�un�40�jh8�"OЕ@�k]6Cu�,���r�ޥZc"O�L�QǑD\�bg�W�|4Zb"O�=�A�ϑ_C�H �X;2���u"O��Y"G<2O�\ ��"y�n��"O*DJ�(�z͘��H���q"O���H�"7Jm�CiϭO��[V"Ot\d�]�=��HSG�!O�)��"O0�g�$n];q��E�T�F"O"UB��\�yȞ�ө�1��Z�"O� p5�3�µN�pё�]�["O�pZ�a�-�F���m`�"O���&�W>8�PD{��מs1���ȓZ|�h"S��'�.i�(t<�y�ȓ9&�P�e턨Ai��u� j��I�ȓڒ\X��J	K�P������<م��I��.m�|}��/U���H��El	ɷ�Q{�IC�ý"��\��i��VHnF慘CÑ8[������� �G�0N��A'_�y�h��>t�#���M5�
���aZa��;� A�JI�q�#TD��a�ȓ{�Dܳ�	4_��Jd���H���ȓu��X:a(֡*Ԛm����ȓ3/v�
@�ٵ9�q���uQh�ȓ1/d%��E͍m���r�&Uo(�؆��+�?`�JDrVkɫp98t"O6��6��
�~e�F�\���2�"O,CR��Ald-�C�]��ԁ�"O�][�C���q����(�v���"O<ᨣ�[�R�1V�#v�b!��"O�����,����|̚�n��y��Z#HtY4g(3�A�sB-�y��ɉ�@0����:�r�9�CQ/�y�e[���,�$'�gF@���>�yb/�
Z|�E�:,@ ���D��y�˚�{Ԥa��*�#�N���y�U]$HE�/ 92�b�ϋ��yBl���\�$L���MR�N��y�@��n�`)x��L=˚��W����yb ��'�R�hC���-�(Y��c��y�����ԉ �hȠ���3{M舅ȓR�pʑ��!�0b��J��`��*�X��ϒ�9�a��G@�vl��ȓ>K¨�4�ER\�m�v�ؼ}2&P��U�f�3�!OS�Eb�� <M�V,����� #ǮM����۝��H�ȓ�Npa�Ȅ�xP̄"^�3A
1�ȓ��U��.�3&䛂��Y
F�ȓE2X���B�H4<�e��?�@��ȓUX�
v�θFL E�[�bć�_J�1�Q�pN(2e6�ȓ�m@�����N�P��,`\�5��q�(($�6SxDY���D�&��L�ȓh�rĢD�S�(���f�O$")�i�ȓ}ɠ�����5h�l�r��PI����/����	��:�Q�J؀shq��~�-�w�/Ll4��A�@%u؈��}����#��-�V`��J&K��5�ȓA	�PȤ�Z�rNAP+7a�݅�yU(A`��H�,M�<Z�+Y5͠A�ȓq����~�̉�MS36��ȓt�P@��J�+�� iQ�{\��ȓ ���)�93��	��,?0XA��k���gLχ_�Bm��f��c��h��o�Nq0���2��&V0peX�ȓG�x�*3d�mK(���$��4|@�0!��M��!cQ�̹?��Ɇ�.e$QB���6cἩ�c�A�u���%�"�
4�C�UY�}
�(�|�f�ȓ9}9�s�Ը2�r���1İ��!z�P�/=�jq��L���b̈́�OFv0��%�/%�fU2�kIG��a�ȓ/�s	��HEǕ4 ����S�? �A�&��Ҙ]ygG2V��i �"O�5�ю�!7�
Y�Q�ğ��!�"OI�E�iAnH����/9�ٓP"O�X��Q<d��l�Q�h"L��	�'' e��ID�	�'$~x*
�'�NT����V��aSE��tޢ�0
�'�����E<%�.P�ת�4s�Xd��'�A�tĜ�8���wi�BV
�H�'8��[&�s�iQWDՇB��,��'�>D�� @�/Jp����';H�dY�'���P��4����DC�3��"�'�t0dc��*C� *����(��u��'B�4+���>���	�-T6WH��
�'�>]H���P!"����S�R��'��r����� W�I���'�I(�e]&Z���5a��j�X���'�8�y�d�'\�h�#��Z�I+	�'
�!j�kG�#���B�T�1�Fh[�'����sb�Ո��҉@I��z�'V�C�
*~��!�O
>e�)��'�:��&��/�VdI!kZ��`��'��U !W��d����z�z�'w~4� I�4���E��)r��X�'4:��"��
{�ۅnݨf�3�'6��u%ȃm��Ԑ%NK�k���'��K`�_z
@�F�z9T��
�'AY�s��̸웣G�/}\�p�
�'?d���B�-�`%�����,J�'�Nq�>�h�c3b��Ν��'>�2mܩC���B�1vlr!��'�zI!`H�0
��8�nĢl
<
�';��P��S(ұ ��A�QF��

�'j�l�?F��1�M�N �Dj	�'���p#)�#q�A���K��l��'h��1 ����rH�4��'�,�Kqj�:{��`�O�|:�c�'� �2���,���S�oۘ#g�؃
�'�|��Ml�!�DmN�eR�,�	�'�]
��3�z�3me����'1��b�5%7,�P�%�	Pʭ9�'w�Q�@�;�����ܾx͜��
�'ڐd��N�U�� RR�E�a�Y�'3� �)��r��YA��"\l��'����*~����g�S�J��'tDbg�_�N٨�(��/F�[�'_�=�6��%{�}@gV�.�zH�'�Xp��m'$MN�Z90Vr$��'���dkF�f����a�Q�Z�'` IR��&L�R�A<y�t�x�'}@4���e�y�F�;c�8��'H��G�xsnHHv܋*�^��	�'� q ���`i�TjI4��b�'�:�Qn��:Li$A<'���'L�RM^.6�jI�ӿhǔ���'�Q�7o�>j�d9���w�ܛ	�'ǎH�����ch�a#(�%w#	�'�`Hʄ�C�Y��Ѩ`�_��	�'��՛pd�$1���;[��y��'}���Y XWک1��"QS�0�	�'<���R�9�F\Q�9TA�Q	�'�h�:g#��zV�D��OH
Y�H���'JHe 6��?��lx�ė")�\q�'��)��<T蒉�r$���Q��'k(q����-o�Œ�g(qB�a��� b) �mBL���ܜX<"�yc"O�\	&�͵i�^Qi��!B��"O��j�b�V� r�"ʸX't�r"O�m��A��3� �*��*�"O>�p�Ğm���*4·�n���+A"O�$���$�p�%�ߦ/	�IQ""O��Ci-g�8Q��F�0���+"O�HҢ��(a�!W��q�"O^x�;^��Aǈ�{�x��"OLaip�ڃ2L ��hчS���"OV]!��X�Jk�]�c�F>�R�3�"Oؔ@�J�;�&XPiLH�RQ�#"O:qY��ىL���QGŬ\��4{g"O�\��I f����c@ė@m>��"Ol��4F�	&RH �«\R���"O�!$�Ĩ �����`S9z@x��"O> ��ԠAH ��F�ЗIBt�B6"O�)
N7)�e��0{8 �["O�1�,��s�,s� �B���"O:���PC�Qb1i�c7�H��"O|�b�cO��>�Y�I���r��d"O���`9.� F�Shɰ5��"O:���$G�`��	Eև8��� �"OL���`�XP�j�d��y ���`"O��B��Q��6A�D��i�1"O^d�c��$���cP!	���xg"O�w��T4�c��-�*�3"O6��QDP�d6#󬐟eaV,��"Of1���dv�=��a�1Rb0�"OR�N�=lAB�AOX���"Ov8+�#^��\y�3s��|��"Or��q�W'y*���7�%/0�F"O�B�ń�U���A� ���PA"Ot%�Rd��IȱCW K�*�͓�"O��S�⋘]� �7a��
��"O
���W�J;��Q�b(n�L�2"Od-s�'1IyB �"K�O�� �"O�,�����tPb��/4�.(5"O�l��O\�G�u�F�]�HM:�"OZP����5#�H|0@��0pqP"O8�y��Œǔ�Ud�+���zE"O`��q�>}"���߈!�bA��"O6����+{ݒ���!S�r�<��"O� 0 �6S>R�x�FΒ1¸�8r"Oh�w��Z�T�%��c���
�'[�}i�
ΨY��'1��x�'�)�v��`���A�(�	����'���u�U.}uN�kQN��{_���'{Tt�F�ڭŚM�P�9b4���'�����+���8X�h�	�'�+0�G������%B2A	�'�"}�f)�L�� 3箑|(@��'�L����C;�T8S��A1�5��'��� �.`�X��UCH��Vp�'~���	̈\0�"P���~lj���'���1�fƭ zH@�
��ar89X�'��(��σ�.� �P�c�mnfݠ�'c�`�榆:oD�Qr�^e�J�'$����MB~�k!�ބI��}0	�'�^j�N/M~Z�{�͞�D�^��'��xxuO[��"e��	�+�.P�'m��m�+j���[p.׈&㢠��'��-������l['f�i8�4��'�戊���)�:m��E�h�P	Y��� ^uK�J�8������^bD�"O~DqC(�LYbhB��"2"T�"O�����/��ȫg�5�p5�"OB �+�eFvĹ�M����DAW"O�r��Z�AJ]�ql�-��Y@"O�m�g �n��2�ں:�t"O�i�� Dv���R�H�W��i�<!�!Հb;��D�b���c"e�<-e���q1��/m���b\�@�VB�	�{����㗮j�,݃7��g?JB�I�,[`�@ Y,WT�C��	O��C�?F��x���}$6䪂��)Y1�B�	�kzXqCq�V!g j,��y��B�ɖ�(����2�=P�-�3R�B�	�h^ɡҌ҆1?����Ѵ��B�)q���S�I���Ԑ�J�t?PC䉳&���"�H�^Q��2��=]J�'��[�%�-m�2����w�l��'پE��8C]�)�Q揎7�dC�'��إjǦ �q:4ß�w��1�
�'ht�!� ���$�q f�9$V�k
�'K8�&I�x��
������A�'�<����9.H]
A�zA6H��'��()�M�+7�$� lQ6>à�h�'�ز3�Yྐ�� ��C���'�t
f�
;��8���?]�'eL��!�Y\w �Q�ʐ�6p|��'_u�����U�(Y��E`��'
MzWL��L�P(�w��+ s�l��'�2U��^'
\��(6��9��<[�'_��
�-�(;�������%��
�':�IH�f� �t�B"�P.A��'u�	���F�0b�t��h�	�'�0%���O�Đ����2>��	��'`\��H�e�Б��-	-=���h�')vT�F���ʃh� :uV��'�)�S��V*�l�T�
5���{�'PyJ� �&�쩴cϩ2+jq�
�'z�X��#�`��9)��s��u�	�'ClH��5��4��(�q
�Ia	�'?�e;4LI#�V9S�j漳�'��)��ې�t]��a�%h�"���'�`,(�%[�@�p�u �,dl��'N�+��1z7�3�iZ:e:$1��'� �Y�/U�3�p)!!A�V��ȹ�'JtJu�
	m�aB'��0�����'(䠋�hǸ�t�&��<����':���̚(�]�.VI�VP�'�&!�AC8�tʠ��$4*��h�'�yp��5j���� (�V���'���)p�_��DxTe��ie��A�'�\L�U���I�(`*bְu�h���'���fA�X�޹� ��y��D��'��qR.àV_��kPi�� �p���'��(Sc�X�K��� `�X�OFu��',8Ze˒8�"`�PjNh��`�ȓTi�m�1%B+Rj"�r�$�"��ȓ9B�[ ��<j�����V"12����Z�&�	�)ٿM��AJ�[=�ȓ$�H ��q	�Q�;��,��-�|ӬU�s�I��Ң��\��R�f��ԩ��1���P��0��@戅S (�=jf0q�	�c��5��H�,���5T|I� ������S�? �dA��,{��@��.�T!��c�"O2��GH����p�^"�)�"OT@r藪�v�:�e�g���p�"OVp��h�~� �2uc]�o���0�"O�u�0���d�Dd�� P�@k�B�"O����H�X��} �O�"1|d�"O�� ��o?@��D���irYB�"O����J�V�p;B	]--k�i:S"O���0�Lv�f!�2Q_d��Q"Ob��Ro�}���[d�JYT�]X0"Ol@p�g* R�#˦E�0"O0M�, �i����B�&ġj�"O^5���]�[{v�uB�=)4�s4"O\�7�D�H���y
s�\�"O����A���8�ա����)�"O���t�	@0d%�"���z��"O�	�M/5!,����ZxN �"O"UQ�՟L7^4�sʗ�RP"O:<5��:9%REPE���/��	"O�ّ�A!o����ج5��0jF"O`,��̍-
��$��/��B$4��"OĬ{$DP)*���i�nϢc���"O������Vv�eN�nj2��@"O�	�(^$2����X�U��5"O��;w ׊���"3��(I���F"O4ppï�- �	��ꚦ�h@�g"O��)wk�Wa��Z���`6H}br"O<tc����.`��s��G/(�pV"OX=�7*Z��JA@UȘ"O�X�c _6#��Pj��X8`����s"O�� �P����9�K�+rP\�"O���@i�<��0$+Q� �TM0�"O�����0h�i��U�o�0e"O�cc�M+�J�P��M�]NV�� "O�$J& �QJ��KV��D��"O@�f_D���U��C>�G"O�U�v�
(6�0ő�=Ą8��"O��94�h��Mڳ&��W����A"O
�Y��G�HN�js�T�_c����"O�a��\���rpߕ���3"OPtPѯݳFvJ��A*l�D�1�"O�lY!FY?!���U�ƃ4��4 c"O��i��\^�R��6�������5"Oؐ��OY
j]j��Q�ЊH� �g"O.	`i�������es����"O`(��a�3����B^��U"OJ�x��-QVb�� J�*��xv"Oh��3,M����J���u"ON-�cH�SZ���	.-3��S�"O&"7X�L�`zv�@�8�@yȣ"O�XP�p��Y����;�B�+5"OT,��8(��XWDF�v�^`!�"O,e���73tj��i�2)��R4"Ob=xr靄�Q��޻B��E"O�Q�Ƅ�<�"*�
*��-��"O<y)�b[��ڝ2�+)�XJS"Oj�↣Y�m��x(�>.�v�2�"OvTXpdXk�X�R�ެWT�P�4"O��Z���;@b�Ys��,ݴ��"O� ZR�]=$H�)�P��Z�dHb"OPPӒ�C�u��e�Ձ���V"O�%�0��4��1hׅ�
v�^��7"O�U2�h�<IL�� �]3�̐�"On�I��"OXD1�J��H�"O� �2WiΗJ��=�D�W*Y�pu�P"O��[�B=�vm!���)���"O��Ze���i��HA�I[8���"OD��G�ԏf���gh[��D�&"ON�x��O"ВV�ÈI��	B"O�Ecdm�A�xh�f�-n���YF"Odq	N "t��1P��7mF4`B"O��K��G?n�0{7!Z1��m(�"O2P8�%̍!XD�*!@�-f�.T��'1O���b�94� ����dMaW"O"�C��94�4�
^%p�5�"Ox-�foX�^�#�ӸM0��u"OT�ۇ�8Zi�1�c��%*(8�"O��5�3릑+�HƃHT	Z�"O
i�7k]�Av�dHfh�1�L���"O�HӃ�\0؜�zd�I�N5\{d"O>8���	_�9p���b���"O��K4m��t�������0�@�"O�h&��*2�N���l�a�^Xv"O�܁���&5�؝1�ɋ6���"OLH@��Զp��Y���acB�Kc"Oh�9w?Q��
�.f3���"O�����&^�1IsO	���˖"O�`�(��Cx�(եW'\ٖ"O`�)�C"6_�A�b%̕s��%"O�Y2�	�D�ˤ��\���"O(E��A�||�y��EMw��"O��y��@�BJ��%�(@�5�f"OP8�B]�D<����U,{�ri�W"Ox�k�O	��94b�)��=6"O�T!��57� ��	>�Hq�"OT�0�j
4[�-!�耻.�-�D"O�U�%��s���h��U��Y��"O�`@p��4�(�����~�!#T*Oz��p�K+s���� 
�e�L�
�'�@�jT�z��4���\s�n,�	�'�hY�fԅNP@EI�j&���	�'��� j�'R�@�T�Ԕ0��=	�'y��9�#ܹ7�ad'L;5�,�*�'q6�R�	�¸B�nB�uRr��'8y�IN.��مgZ���':j��� ~��JT �>^d� �'�`rЇלT���,�,^�`Xy�'W>8y�6 �b�>S���'��p��.*J��*�EKL4�:
�'ʬ%� ��J�H�ƙ���'�K�<��CU\|0���
W���&Ol�<�vbB�u�\$�N�?��%+c��b�<�ӈ��S�����:"{&���Ta�<9b`�a=���X6v����Ff�<�3D>&^�
�'�
��kSV�<���,t��kB��~s(1`ԈS�<�A ���J�TρX�<�w��ve8���P�:�&xItY�<�e�%tĊ	v��Q�ˇT�<��(����S�MW�)p�M�Q$L�<�i�	�*= �,׺ёN}�<Y�#Ԓd(P�'WaQ�|�<ٰ	��cx�=��o,*(�t�bK�D�<"+��M� ����ɨH�\�2��Z�<1�C$6�su��9<ZH]r�
�R�<�5��]:
!��jC7n{���s�HM�<)%���;RȢ���	aXy!�r�<�gT�rtf+�g�.;lZ呄I�o�<� ������sY�d����>T��Y"O2%acIM��)B�
�(;&"Oj���A.Ul�B���!�����"Ozȸ��W7MU�q0s��~'`�Z�"O
�	��Y�����:yX��"O4)!Q��&�Ġː�	dl�p�"O$�"hO�I(`)`�ӷxg��!�"O�!�F�.�p�����cf����'Dў"~B��#{&��Uו0Ŷ=q� ���ybOC�_�����*A�+UpTc��Έ�y���*|^��(&�W�+j@�@`&ќ�yR"3,Z�u���O�\1%[��y	��\��Q�0k,4(A�pFZ��y��L� g��G�������N��yb��		�i0]�i��TKY��y2�E23c�xkf�'(�8��N&�y��dBL�S�ƣENP��R@!�yBɹ=����s���?�2<�Q�y��) ���O�;�udɊ�yr�F9:x����&��I٢�Q%�y��E�y�DS���\�	��y���#�l�2�"G
yɺa��'�y���D(̑�C0x���㋯�y�KK1EEƅ��u���2 �y�N
Hb>@ 5��_C\u#���y�9OF��2�a��	,��8���y�_�H��㎎TH���ά�y��.^]nP����R�F��y�k qg��� e<|�@lpG.��y"��|?���댕vTm�A�A��y2h[�i�EGX�r�^l�AAU"�y&�t��y�V�Ғ>=z5�q�ʙ�y�#�+}�0	�'��0��u�5h�(�y"�L�|Y�!�m�51��`30���y���{�@9��&X''*ؐ�P._��yRG�J N�F�'#nt	Ї��y2��Kq��Yt��#/A�<�' ���yr
X��2���ҼXN��
��y���c�a�1��49�J�v]�y�/$#L�8�	�,-��-:�Lg�C�	�n�B�R��yK��!�5%�BB�I�c0�s&o�(#ǒ+�%o��B�	�?X|�Y�/�
)]`�*��G;j	�B�'�I�AAƒMt	RdHD��C�:�@Yqw�M7C����!��_��C�<|�<K�@GN����$�=Vl�C�	9�<���߷Yܘm��MA�d
�C�ɴw�9V�X�����o�*Q�nC�b6� �/i�F�(F���#�>C��T@jȥ�M�V �0�7�Ų/>|B�	�Q�)�/�8)��|�Vk��.B�	�j����݈V�$�#+.iW�C�ɰv�e�-��v҂t BhW�p1�C�I/VY�T[�M۽?C�����Y��B�IM�z��C'ȤK4�!&N�5��C�	8H�z�c!�S}�v�K�4"B�ɲ�H{�A�h���V	<��C�	)��SG�mt�[�p�B�J�$8��4}��q��'�L%�B�ɺ}�@�����P&
2`B䉢#�8!rr)C�O��a'��b�FB�	Dz9Z����T [�OȸMM B�	�Ub��e��vn���OG+1�B��7M�]3�E��N�<�D�EZjJB�)� ���#����x���.|$�p��"Ox|� $M[�ț�E�I��x�0"O$���6�<-��#ȱk� ��"Oz�"qi��a9�Q�^
#��8��"O2���72m�+�.�.a�p� "O&0b�L�V\�q�gc�E?,1�"O`���9�����.R��"OV�����bL���l��>A�+U"O ���(�sM�0���.0f|��"OQ���¦5bB��PQ��M��"O�0�@��t�|�b	J�
v����"O�C
��~]c����Mh�x�&"O�4 �㛵v��:I �}Rl3�"O�A ��:;0����й61* ��"Ob����^K�W�<9��x��"O��8�dTɑ+� �`'"O��t�a��E0 nсb�@���"O�%A G�.� ���k���A�"O
��ǚ!b��9� yu����"Op�C��A�*5`��aQt2e"O��0rA�T�b<  \Z��q"O�-�c,�Vx	!��Zt���1"O�d{��>"��Y��\db���"O��"P���d�P��$⍔AS@���"O,[,��6��T+� �dF�`b"Oʨ�'`;K~5���ۻ0B.=��"O<|����T<��h��Q"O�X��(�.Ċ�͙0�z1�7"O��$�k�v�@"���?�fp��"O�˔��9/@�0���N݁W"OX%���TU��}�T�ݚvͲ�ȶ"O�	�aLS�8L�crGӂ/��)Yr"O^�ك��]�f�j�EDQ�ꡋ5"O��ҥ��k�@�
�YNv	��"Op0b�� �l�x2Þ([�] �"O04��d�%��PBrB�Yj �"O�	J�H�"qS����A�^�4� "O��F��	������w�4�A"O��q�hPNYЌ:`�)��]�'"O��!%E��:�>��6Okz�]��"O��K����Jh�a)bF�� ���"O`9[2NVa6�u��X�d�R8�B"O"��KE�)�l*rAS�Q	�q5"O�AG�?-����R����cp"OĒ���+>r�d�K�6f�fI*�"O��0�灓�n�
��IKs���4"OF�"Ph٬Ow�3�$�Pˈ��"O�� *�#9���d�AEi@А""O��!�"I�:�j��(Uy<�S�"O-B��B���$!��2k��s"O���s�~�4�� ;as�"Ot�W�ޯ3`]�qc¸T*��'"OB�s�B�3Ut�2%��<%4��"Ox��m�+�8�Y�`ݴ,�T�"O���e�:��"��)u�����"O�(�%��\�"D�@,7m��T"O,�rt�ܨQDl���N*"O@U�d 2d$��  �8MZx"O0�{�m�u9pxq�$AYL<���"O,P4��*H5����?@E8d"On(��܆C�XYJ#؁}+^��*OL$B���p}Ha����Q
�'�A�)ę?��sPK�!��h	�'>�x��)��"H��d�	}�	��� �\�͒�d�v��u�r+"OH�*4&D�R$�K�ʑ4Q
L�p"Ob��0�;$��0D
�K&��"O$T�2�	'��(Ci��V4�)�"O���\ �E���1?0��"!"O~E CÉ��T`"����S�OVO�<�
lA$��t�WP� Ik��r�<YCI��j3`�(������T��r�<	�k��TnL;�GR�E2j��w�W�<�cL�� ���2懠R��4��@Q�<y��B�,{*ٰH]u8$�	�K�G�<1gf��Km.x �T������E�<����;J�)�%']�YB1@qjE�<� ��3j�4��8&T�kdw�<�aI�>����8�{`�q�<9��?]�i�IY�;�t5�XQ�<��A_�_�ب�Q"-0<�"wi�G�<�'O�f��r���ړA�J�<��Δ�B�X a'�ۯR�c�XC�<)q'*Z4��QR�۫w/���l�A�<��'�ay�E�r!�tSୠ�+�{�<I3��1"#��%�K�Vs�a@�${�<Q��it(����P�b��7�LM�<�S��ohN�r��ɲ�>��[t�<���ԑCm��+'�2Wp0�k�a�K�<�!m�z��b�!2&N�;C� J�<iB�?Ȏdի,|0y�gD�<��m��I&9� H�j��*A�<a�O.a���J�g�?N��N�<�$Ո<V�����4
Y��!�F�<�'雒Q�|�ғi�
o� !_�ІȓK�HI��=�bp�%�n�|A��R�Q�Ǣ�V�Va 4��jb�l�ȓ��,)��_u� e�֐?	���XT\�z��_*�� x�E�%��a���lD�IW��mAm��:��ȓS�d��Bo�{rn|8�J�P��5��*�|�D��̰����-��ȓ,�~ܑ`e'?Ԥ�3 �f����ȓ-��9��g� "+��c���3������-I�S���"bG�B�,̈́ȓ2��;�ʇ9.dP���Z	����8�)2�+�#=�%�@�.-jFфȓW@(�2�J�Do4,�UM $����q��Q�b�\MB�b⢈�����Q�\�s�CN�^��#[�u�Յ�X���R��-&eJ��7Ն��ȓ&�R�"B���_��@�U�ze��ȓYw��14-�1$�5"�!d�p!�	�'�j�	&�&@}|�C��$���'��d���c��9y���� ����'p�� �F�'޸i�4P	(�
���'e�99���0r��{�d�*w�d���'e��a!��k -��k3(�b�'�*`��*?���cF�qiM2�'���ժʅ5��h�	Noljк�'7ʌ���Z�T &��*�@�Y�'�N�(�m2!*@��D�)���'��!{����5�Z�QcJ�8P��i��'P$Uz-�3<V$��A�K��h�' 8	)Q��;#f�1����Ʊ��'�f$9��1j���[�T|=��'G�ԃ�@�(oa�A���#R�R�i�'?�Wa�6���@�Cݐ�a��� ��ʉj`ѓ`G��0d�c"O:�8��K8A1�{���QѴ��'��ْLF�9 j���	�P(�'�6�B�� �b�7�X�}����'�����I�-}2Bi�SgS?(�\�'�ʼ���
8��p �(S�6�����'���X� ��$��]M]4+��d��'�&���
�7>ʼH��
;.��'��c1hؕs�J�(e�!��Z�'L"�BF
(�j p���j X
�'���Q��J��$�Ǐ�:1���	�'�����Wbւ��W Y�j���J	�'b�R��S x��I9��6+�;	�'X
�Z�	@{h00�^&#�
���'����%Vx$pF޻W(h�'�F��!n4}�(tZB�nX�2��U�hQ�0P�#�
���$7D�H��f�
��� 0J��h��CD/D���ŝ~�b��i�7J��	�%C,D��¦H	S^a�����m�>D��7C��$��0pvO?!A�;D��` ݙou�����?s�!�P.$D�@�F�ģ.S��!\��5D�|�qӠh��R� ´F�!T�.D�d !�Q&}����AS9;���'!D��Y"ǈYkV<ڶÐ�4���C !D�P�tC <�B��Bˌ�E����)D�P*��E�.�`��G��{vb���)D��hԁ qX�ԓ�*J�<�6�qrn(D�T:�F�O�N���Ģ}W���m(D�p��@�)��R��2&J�L#h'D�d�g������aL��h�p0g'D���"��}g��2K?r���G�%D��1P����h��s6��a�#D�<As�l�
)�A�T��L��4D��!�<b�������lЌ$8b�6D�D����1>����b7+���&�5D��{4i�%|\d�&H����AQN!D�`��^�H�!q��5  x�#D���mE�ݠ�q�(H���3SE!D����K�'D��`ӪF�w�:0�� D��C"��Q����C�P_�J@�!D�tP�0�>�e-Λ8�Ka>D�8����6�`�"̼�<��r+&D�d�윯���KW2��\;�+.D�\��_�S�
 ,Wz��H��*D�!af]X���a�;�P��)D��j[�����LPx�{q�(D���J����6'�#�����'D���F�?�
Ѻ��N�F�4Ib�%%D���G�*M�vI�&lǬdg2c�F6D�tFhʼ��@�b��N�,59�o4D���ß�U��R"j��b�AY�'6D��!�&�!"ʸ�#�i["b��8 �!D�Lz����*%||��� i_�S�C D���#��)�(�)&g�ų�0D�(��� Z�)��,B���Q�#D��s�i��k"e�p���n8��!D��y�LP�?��|0b.*ZܤY�� D���Lޭj��MX`-d/��Vh:D��br-L ���7�
V��+�4D���0�ŋ~��͂va�?e���3��6D�DS��Z�U��(`��'2���$2D�Xj�AE�F<� 2E=yv�[dg=D�� �5Y$��s&Ĩ����N9����"O�`p��L܄ /��Y���"O�����\�b��,{��"ObUc�W�g��p�f�0eF�X�"O�̉$�vع�F �T�@q"O���ܽ<"ȥ�HS'���#�"O��D�,��7`���V�r�!�Ҙ%��eՅR�$"o�%Z�!�D�	u1�Z�ǩ.�������2�!�L`��)�≶	�cQ�L9c�!�D>g�tI2`�N��f�Z�%�!��BR{d%�$��>՚  ��^�!�dݠ)�� �&K�g+l�YU"U=�!�8�4+��W.}Z�g�Y�y!�D*ye,$���+Hm�-�p�\�^!�$�
6Vx���C�Nt9Q�ɀh�!�D����C�Si>��_''��ȓA.�4`G R'+�HHi5$ ) @�ȓ]
���BL��\�L����
��݄ȓkk���"p�J�����u
��ȓ7{ �����@����� 
�ڵ�ȓ.`̳�y(�,Za�W�x����T���$�C�y�|���l�/�Ɇȓ{Jz�C�FFX�p!Ϯ<�H)�����b��H�}z����֎�ԡ�ȓo�q�6���+�����,,���ȓ<�ŏ��Fւ
���B��A�<u
�{yֵ���
�2G,,�Q��E�<Q3�8\2�����l���&�@�<WI	�
�[��ņg1T�qNS@�<)5b*:H��1�+��O�\YG^~�<Y���c�0�CR�Ϳ&e�]Y#K�<��<���!�J�20�P d�S�<��Z������tj�[%/�N�<�%&��@LBg��KР����H�<�g�qZf��X&l�USB��B�<�q �
!x���� �zԢ����Q@�<�%*�)uϔ�C�l�u>̝g�Zy�<����=I��Y��Mq�.b7�RN�<IA�D-(������:	��A!��^�<�jO<����ÿw: 9�GX�<9��7L�8�ذ�߸<3�1GK�<��R)C�:�hX�1)�h	�e�R�<���	�co�T���O#���� lBs�<�@ˡp3�)p�A�?ۮ{�Dx�<�!Ãxq� K�XYȐ�N�<	�ŗ'm�)���'�n�9���J�<Q�C·^.�ɀ�*[�UPL�b�[�<�Ո� f��6�V�R����%��_�<�@ת\zU�Y
+JP]�l^�<1��(i ���(�!6n�BJY�<�V2%`��Jӛ-�lEZÄ@p�<!Un�9�(y�A�c2��U��r�<Y�J��B��
5n�����e��Z�<�!':��V�v6�;q��j!�C>j�)Ҿ����Q��<N�!�Dѷ[��e[���xF�F�w�!�
�b�Ȫ0���K���I�DU�p�!�N�7�x�V��m�(<YF�1G!���;����O��� �4�!���L��{���+#�
�A�I�	�!�Dф'��-SwD#Y�$u��K	u�!�D4f���DڻM�@��� n!�dֺ7) d��]�,�pl�`��Y!�� ��F��	���+[;
Y(�¤"O�,��D��4#��C�lҏ3Q`��C"O4JE�u� ���S��Ε�!"O�H(A�[W�@��gе��ct"O"��vi�o�d@2��i����P"OxD��p�����@,3��Q"O�u)qdE�K:���֢+����6"Or�ce�]�v������F�w�<xe"O��k���z�8�̈́Z�\�"Of��C�&/�U�­T�>�0�k6"OP�c�o	�SS���L��]���P�"O�$�d$���H +W�*����"O���!G@�]t֩�V
��GD���!"O(�#Յ�a����I�&b'�0�"O��`NH :�z���'Õ(�}�'"O:(�R%�`h0e �+j3h�"O�XZd�T��
arTE��0�>���"O��#�%Bm��C�ʳ��#"O�D;Qm "n(	�,o�X]�4"OnH��)iG>�
-Ǐu#x��"O�Ip3�ʚ~bV���ܝM&�2$"O\�-Y��3�^�'<5������y�y��y�ĢŤK7LxRd�E�ybD٫4l���G�z��r�����y"Ȇ?�ư���e��9��(�yg��3CPT�D+
$aI@�@Q��y4�M��^V�b�h��y��PR���]���at�B��y,���З�k!����?�@���'�j)Ct�ݽ-�m�+�2MV���'���j��-P�"�J"^Ut��'d���V�ʒ��$�7�Y�G<��8�'��A��a�/���Ǎ�9�(���'�d����T@]�ǉ0�j���'O��(&��k�Dl���@�&}I
�'��Qq䎚�rhD!�'	�Xl�	�'&���땪SC�ȋ��\�󰭢	�' L�r�܊F|�����ԛv(� ��'����f��P��FN:^��*�'�n�{��$N�H���������'h���=�H8���ۮH�B��'e �]�>*�ۤ��OK�=��'�R��m�tږ(Ӕ
4O�H���'�����LF�M���%�Y�������HBD�Z�t ����6!򤎁%����E!�|���!�D�*(�#��\�S`�R�F3(!�ģ2����q�6+A���ţI$m!�V� 2h����x3�z#܄7S!�d�M��;&a��sN�0wdϔ7�!��q%�e����N��(T$�'�!�v�I�F��M:X��a��W�!�d�v��c�t�%�ǀM��!��Rͦ%���p�|� �@��!�$�4I]B4	@���}�Ǎf�!�D�.S�n%A�F0PU��
@��H��y��>����V��>�^��G�v��B�I�9.L�+c_DX���(A֠B�	Ak��ШI�VVtٱ��/O�B䉩I��q�F�0sG�+�l��8B�	��8��͆�E�!��EL?� B�;I�vp+c&C�+Z��jT��7�.��ɫ��?�ӂ���\��@�1P>��rʍg�%�xbP"X�l����ռ^���B�%3D�� ��� ,�l�\�P��J�V�p�"O��p梛�`b ;�%G�7��(`�qӢB���s��/0W�P��Q ^]�C䉀g�(�.�4vU*�Ƈ9#�C�I�u�q'�$�\ݣ���FC��Q���҃	1���ZXC�I�
�
��P�,^��J���a�PC�ɥUܸ1e�C�j���� �P5{y
C�ɼ]aZ�*����m��p�͟/*�C�	���p�ђ?�����X�k���� ��īc��S'hV�:p�xQ�d�"�!�
mؚlec��cP���Ą�!�!�$��A�4c�&L�09%�
�q�!�$@�����-,^t�`���!��
��t�0�	&H����9I�!�$�0���4���'�~iJ�n\=�!��6���ʃ:/μ:��٤�!�[�4�.�� @A	�pDk#��%J"!��?O6Q�
m� �����	!��D�/�.D�r@!H��!��ޔ�Z|Kv���g�b���Ҽ9(!��Q-@3������	r4�*�FԳi!�L>9��M!H����+!�D̈�p���AT� pRP&H�!�$4eP~�2AA�*><�ؖb�!�D^��f �F�%\��%ʁm�!�E��Y匙08���� w�!�B�M�d�I�Ɛ8y���P*��il!��*n�N��EE%e֚��]���<ON�r�
�g�l)y�ės��lړ"O>��r`�~=�lA�Ć�r'��������	3C-2�3�G�K'�Z'M�>;3B�I-B/P��C� =_`�t�ۯmF
B�	"r T�F*Ǡ�����#�DC�	�+�V�C�΃�O�=���'xy��hO�>��ե
�IS e����G����,0D��p[�+ʥ����$���C��-D��z�@3o�&t8Q+�f���;"j0D�l�P"��1C��cvI��"�5���!D��'�Z�*���[`�J�	ָpc�m D��{u�����s��v��p�l>D����^�m��)�bj܀3�`f�=D�����Eȴ3�X$">��1D��9h�k1�@��+�U���"c�2D��� 1O*���R��03a�5D��x����,L\% 0�O��R9�Պ)D��a�"1��IT�sMx�Ӱ.&D�x�d�ƷuBtmQ�.cٖx�6�/D��*�ζ%!�В�ߘw�����9D�����R��Us"�ȘP-�tb�b�:�=E�ܴ&��-�H$b��0�ą�3�d��2��Q�RM���2�/L�t�D��'��|1,�F�i���֧0�ŅȓH������&/���̌ Ǥ���K�(����߷d� PĪٙ8O"�E|���9)L[ F2n��QjF-��B��/�|9�Z�b��x�S�<��B�	�8��uz�X�mc�L�V����'�a}r�(jD��޾�`A蚐�y¥ �M݈iY�1~~��6��2�yBǈN�\�r���=z��}��W��yBk�-p�*�x�i\)C�^�Ce�ï�HO��=�O�,��1E� ԡs�ș<Y�����>$������<�Le1�2�hlr�.9D�� lZB׳?,`�qPԼ{�,���"Oh<2���U�����D/z�T��"O�X��&�#Q���"J�pk����"Or3'(�$]X}�a�[�DTH�3d"O�KWG;>�����<k�ba`�"O�qA��C/M��U����*C{D���"OLI�ԫn�X���ʀ�&�QHT"Oj0�BO�uuF�
����Yn2u��>!�0��(
�9Rx�x���!X�U��D�Hh&��J�T�Y��s��)��zB�'�H�")I���/7�Շȓ`|��:2+��&y������*�d�ȓC�D@yc�
y*�e��o� 6Gy��'3�5�6퉞�j�:�nDh��L�6C6?�O<E���yM���S�G�7Ұ���#�/tCf�ȓK���U�n�ެ��%بn<1�ȓP�\! �ǚ��s���g7�,�ȓxI���30��p�lC>���<�O>я�i�{y<�k!�$'�49dLO�1:!�$�k��e[��pD!�p	֖&(!��(pv*�(ݟHr �ș,p!�d�S�(�ز� �ߤ���g�?�!���A��9[�=Y8z(i���ўdF{�o�O@�1'-W�.zf�QR@U�2Tn�t"O�y Ƒ�(�0�6�ϫP��Q1Oʣ<1����!���2\Sވۥ��[�����'� c�p����D;t���_#T߮M��n`��=E�ܴ�6���a�`At�B&�3���=�����4�ɚ�֥pV�[51h@�P#����D<�O���u$<G6R���N�l~�� ��'2�	��Q2���+���)&K��C��2��-J�j_�@����t,=P������5���q���g*��R\5��BԱe��C�I�ht�<����(�N�
�D9U��ʓ�0?gȄu�4�����8�μ*��C�<y�'��C�*�8��=q��hR�a�C�<Y0�c���
3��9$�`�W@�<��F��m�LQ2������3�@�<iLՄc?69a`�P?d���
�s�'�~��ď�[�<�Y�n��70��:�N�6u�!��S1l�QD�$>B��Ю�7
e��(� 	SWn=2����lv�]:��)�Ҹ'�
��N�q	�..8�h5`NRl,��"O�`A!g�-3��) �� x-���"Od�Iܣm��H�5E�!�x�P"O0���@�j6$D���"F�
��w"Ob��!���0�rq{t����a�"OH��#�,	n���@7�>�w"OƁs���1�^��ƫH�F4�"O�E��9J}��*�R�"O��Ѣ*P�Xl4Az#�F��e`�"O��t��&w퀍�`��/v,x��"O�8s�K:6��L��ݓ4��	b"O"	i��A�D|d���׆=��"O�����",�Ą��(bE��"O�}��3j�)��c_�B�r�"OTDH�'и��D D��EJ""O��CA�,��ׄ,j�jHѥ"O0�R�ɧl��r'&� w6�#w"O�U"D��i��ē�+؎$L ���"OB�Q��u�(�mU�Y0�!c�"O@e���bMȴ�'�2��6"O�P+�C�Y	DL��ס}�E#�"O|5{��C�^�pI�#��$Y�"O� T��31�[��1+"O9!5��7� �17i�<|T` [e"O��teр��=R���}]4�"O8��G���H���ꋧ	L����"O�-�2g>��(;�H
ZB<�a�"O6И���aHN4��_|-5k1"O�`��-s r}�����"O>l�R����:��M�h�.8!�(D�xCdfAyX�B�H��F0���C%D�\�G9$��LIr�G[t�y{ �6D���f�"�^�P��š[����06D����o�7:��ׄ&�P�2ƅ5D��2�DA(0z�t!�jW�s�XP���4D��;p'%UnzH�V�Z|����7D�Ұ*Y*r��Ek�f�?d�Yy��4D��3���5�b��t���ٷE1D��C��+��#@��]�ʔ:�!-D�TP���>p�N8KK>`A#�*D�<�R-A�.�ё@@ޘ
���� O5D�<ZKV=TVȀA�Hݡ�% �!�S)U�>���!L�c�>h2p�r�!���K��TߠT#H˵�a�!�D�M�T�2�U�(���"�ST�!�d�3*i����N�;\�p�����*#!��Wpg%�g���aT��%QD!�U�u�d4 �I1�%c��̋Z�!�\<䁐fd�D�T�:}�!�"T��f��9��`��/U,l!򤊤N`�{P�M����#2#�=x�!�dQ�^XX��MV"xf̛��_�!��҆^�D�Qf@ByB@��Q�h�!�$�6TM&=CbԿ �Љ;VG��k�!���Nl��0�6)��`��S/e�!�<IJ��C	7�&$Xv�K#x�!�D��C�Tkю[��4AaC�)�!��ߵ!MR<��ak�i��o�6`�"Ol)g %5��PG�S�l��"OP4�G�
=/3�1�C˳f���6"O8�rO�!1m�(��B�)y�"y"O��zǥ]&a�~}�`�Կz�P��"O�[ G�i�:Y6/�Z�"OX���Fm-<=7�Ýb���"O�\�V'T}N�R�N��3�J�
�"O��)�c[43�H0 r9uאּ˃"O�{�%�&H�� s��?w��c�"O ɑ�͗ n����-�/e[`���"O@y0 %M!(�M:��*=i��Iw"O(�ʆ~\��PEb�2}���2"O<t�V@�_#�L1�?)����t"O�1����y�U��bF5g�̱�t"O��AI��Ð ��#ݘpQ�"O0i�㆚����ǅ/`��H�"O�H�#B��=�V��Cؒ�Hu��"O (�W�A���2�e� �~�b "O�=y������{��%{͌)D"O<؃���4xE��#�Þ�d��L�@"O�Ę VuB,l+4���T��]�`�|"�	�U��Y��y��DN	;7��A�Ǐ<T�a:&����y2�O�PO�mJ@�?�)�'ل2��XM<A�O�a���'[d�����$����UsT���'0B�B�(�*j��eME�Q���ĜF��a��Ƚ��>��)�j��S)B���%mZ,zaxr����D�cL�-k�f�T+���s�d��dEȉ`hХ�&&)D��2�M�D�(�u�;J�� ��O�@[T���Zc$��kO	&��";O,�U��J��g�? q��н*�҈�%ʀey Un"lO�L�r�YJ��Es�͚���1P�-P�>B,�M��}���"��݂� �dO�jy��	�l�3���@�t�a!@�mB<:��Wg�Z㞔R��2r��
�#M
k�e0��)�u�,\*j����ׯý0=�D�q��=��|X��F
z� �kcC��s8��Ě9uWT�JH�6Ạ���)c��k���M��hXS.�h�ԑ�q�ڹtRZ4�$*	1���(e��ݞ?:���>4�zD�����Yo��d�1GFD����3����3a�u��{D�?)�F);�k_�=�e��a�����R�fnn�#a�B3A��!�H�De���ÂM�CJ��+���3\�����	BO��{�^�Y������93Ұ���O�1��=��k�1�&xa��
?��$9�jZ�/��	iÎC�0վ���N/�?]�;�Lo�b=���ݚ48%�4��i�1�Ł�5Ö��V��}�ֵyC��<T��F�=V:��U��BL�	6�i�~ȲӅ��]A,(ߓC��5 3 �� F�9���`���7�3�a �eOn��c�@��)8�@�1��A�'5j�����5v��K�biq��;CMڙ���<��xR�F�suR%�0I�V�aJfř�t~PHWgU#�(��A��eT�!j��FsyL����Y�U"�e� rf| �g��l��xCH#JW^����g��y"ȏ�I^H���N`�ش��J�I�
���3$S")PfLѦ:�Щ�$�//C2�ES�`�Y��\�N���B�ӱ!X1O2���+?y��w���Q�Q��|b��Y�}PG��cg�{8����eXw(���[�m�� ��f�*?D�vF�&Af�!�&ΰ>adE�r��.hdv��DO?B�Z��`i:(<�ly�eƊC��k��D���G�E������%u�-�&B݇L��}�Q
�+;H�p"G_ k���I@�-�P�؇lü� h"�O�5Z3�]��e"��2]+H݈c�Y 0ʪA�U�]'`�X=��Bԍ9$��l�]��Izfm�X ^����7�,�z�m�Tz,qc��@:n�a��'�^u�N[k����ܵE�2\JE �3V ���`bʂ7<�ytnC�UB$C�bL?	)� �!@�(h"����P-��H>���� �FQ�3�;5��t�G_l�#� ��wk��m�#�e����zb	�z����Pf5cZ�����ԯC~��Q�( v��mKV:|fV�RT_F����!���`ń�n�P�ȫ)�B0	R,XUJ$���F�|���riŐ&Ζ�5d�a�a�'	(/�R$!R�̭v}|E�� YT���'ݍ,��B��6�>��$��"u{#h�)|��ICkR�I�a�@�52����K��(��d-P�*e[c�X���睹a��D��l��8P�!J5����
4���V+�.s�(���,MZ���E
2e���z�oB�9atт��D�-P�+6�/p�88��&V�K@�%��i#F͑9P����7j0E�A�-,O���G	�,e�X��0bڔ�v+\?v��Y%K�JZ,B�KU�n�ܙ��ǈR�n���d�#��<P��	�����i�:z3j�I���Q≠t�lȺ3N�(%PS@��}(1*���.8�Ȍb�@��v�\)�I�]�~����M��ƀ�@O
щA��]�v��Ea��E0
%rr��b	�E��]��+��Ѡ#���V�_�r���'E31B�1�$L�E�d�b7�{:�	�Q&ե��xr�ħ����F���W��u�B%�*��M��h�	h�\()%m��)X���'}������DQ��I���(?)%oߤ5L�1�s'���X�ԉKvx�8�3��1��p�i�5U��q�"��� ȩ��1>нb�EG1)�$d��A28�c�]*U_|�����y@�>��P�(;��'��\�C��:�x4��Єbd��S�M�:�*�k񋇒�q�F	�pJ8`�#�*N�x�!J�dm�؆�	�5�
Ы���	9/�m��t���)]j�a;�oş��Ġ���{�� �� �^�A��K���ا9�Q��%�(tѾ�k�h��4�,�"Oʽ�$��?l���ϵU��0`l�O-�ƭ~z�Hse���ȵ��6z��6S��H�'��d��(�s}0�#S*X��4�XדL�̄:f��+��C�ҞAix��&��Pb�H��iC�r���QDfn�vtx�F�7?�,�q�GfQ�,�FS>N��-I1���Xd�/�����L%{��q�d��Ya(�"m� av%���b7&�bg�!F� �9r��b��;v�<w��B�C�%�h|r!L�`0��g�@�S�.����$�8S�ݿ�M�5*׆9O���ؼ�@"�� R�M���C6e����aTZ�<�A�R�E����ǺKsv�ä��}>}���>�yRǗ�K�٬;K��Qt/��4��/҄�~�j�;[b4m�g��agBdj�I�$�p<٤EzH��9��/����G�W�[�X�F�6BIc�e0|$����J�n�8�9S@U�@Wx5���[	XQ�4��.�C��� f�#Z��� ,?i�!�!C���#����H����I6�X��Ƈp�]�QeQ�f�p8C �oc�~B�Zc�� (M��)�3�ۿ&���y�!��
�Ĥ����";���c2�Z�I#9���S�wt�Y�C,�� 
to��ao&U���k����IѡaU�ՀČ�e�zmYSY����^>B�'�"�E��=K��"�	1�j�'��՛sF@�x�F�qc��+b�!��$��;a
d��LU�<N}�򆑜E���#��[5�yi�gЬ����䩗��MK1k9+$�(҅��\�&�zŊ@���O$!�w�R�'�R������
�(�C?!�d�+SR���q���A� t:��&wFR�R�E_��VH�LśV�<o���2�NӸm�`�0��{X���_j��L��٫><��'g��,�4�g䜷J�����!��z���ϱz@�7MV1Qp�	=��-Q�w�f�n��5OL���B�+k>����N���Ӂ�:� ����!%P�@��,#G���Α.3*�DE%~�I�t�f�91�%|�#c� r^���Hh�&ՂG�8����P^�G}�� �m�F �mBnb�`U�O9Bt��U�@���8��T�Q�V��d��A�V�2��PYa卄�H�
�!�(5�n��3�EH�<��1�@�
����,F��Ȅ|�ld�#o4s@�=�RD�w�d�7���M����d�0�� �5�� u��SR)F(R<D��Ď���	z�i/@1��X�O��$����3���Z��	�a��T.O3�MKDf�[�f��l�2s�����������`Ǌd�x��$Y8� ���C����#TjZ�J��D*F@+<�I�+K=C��=��+'dD�� ����k�j��I��lr� �Z?q���)n�� [Ǣq|�YiצN�'dHa�E��s?�ۃ-�:5�|��f�K�P9 �'^Ҕ9RO]��,��ĠL/�D��A ��	@K��O�TS��4a�,�+G�C�4q��B�Z������G����ͪ&М0J�-٫�ԭ��Č�;�ʘ"�	�[�=Zt��]��,(��X�%D1�Ŏ���?	�	Za�ʐ5��X�б���r���0f+��Rʮ��%����qG���e�ƀ0�[Y���.�ܼ��)W�WȾ��������ɫ�g�V(<��кD���q�%W�Z���3LYk�ސ3T)]� U`)�U.ɾ<Ɏ�ɶL�E���a�eא[��Ã�>�FE�t" �h�Z:s��¦+�b���*׈�zi��o@�.��L���*7����HV5/�H���{:�Z�)8<O�!��#"B�W���u�ВiQ�(���Z�'N�DU�L,Z	��9��ʷf�dS!A�@��OT��B�	�R h���i��s�%r�XK�`�	�O�ҼH��s��t2w㑨�d�����>w�vб kQ=���ԩ0K6B��7����VW�d�&fW�<��QC@.��y�d�a��ʇkjd�#�:��*=�I'1�$B�jx�LQ'I�/P!J��d��Ld�%K	W���%P3Z9�����U�����%�.#Z
9���'|r�d�̶*�~�p�ʔ9���dR�1ަ �a"��+U�t@ �O�?�K6��8 .�lKg�D0ӄ�;�-6D�����$���d־��5B�5?qu�-#v	[FH��蟰 �BL�/�v���-�*oL�"O����܄a����<���V��m�� z���e,.�3�˃k�2L�E� �p%K����ZI���B���U9|�مl )-��4�Ί/��~�
V�hLW���"�� L �y�� m�4E"S�VƬ<��A��y�jV�?��4Ҧ,��W��͉�-�yݯ�h|0�e�:@�Rtg\*�y2��QG&%�u @u))�V�Ʃ�y�f7�P��Ly1kП \�ȓ^j�d&���r)#����h�LP�ȓjKl����$B�ʔ@����9�ȓ����A"@��j�.�5�ȓ/�a17�6��Ա��Ą8��x�ȓ)̕ɧn^) ����J�~���t�M�ʃ�*��J&!<c�5�ȓ1���P��ںP25�R͟Ff(�ȓ-�eY&ʑ<J^�� �,�[
Xԅ�>�8}:�J��9ߢ4��K͌=r�|�ȓ�2,�ԣL��V�R@nY�r��ȓ"SƘp��q��s�Í.`��*�r��"U� f�	�u�:e�ȓD^�ݰb#��rh:�4΋=L���&0֝� F�S^`���"܆ȓ���a��V�.��4�`��kW�t��wP�LJ)D�{XPp�I� O�Q�ȓS��1)��Ӻg� h�J�I��Q�ȓ,�^����ËS�lأ1fܫ4ҖY���B8�7
��d|́w��%B�D�ȓ�z�R�)~�h� �X�v���.P5�Qc^ah`*�
�>K�X ��X%DIѦ钲'w ����4=�Ćȓ ��� PF��}���y�~���?U�u:" J�/z}a�dF*W���	��9����q�q�1i�:��I�ȓC����S'Efb
�W���m�����q�u�mQ�v�xHs���.5~Y��S�? ��+�_�'���K�:Lza��"Oj h�O�)�<�y���<�z*D"Ofh�J�$�Գ��R���a�"O����YD2K��]&����C"O����✴+��i
��Q}��D"Orpk��!N��pV��iDµ�@"O��(�嘿[(E!4͏�$l�{�"Op��HC�tm�AiB3wh��+s"O��x� :jAj)�1,�cE6Y{�"OpI�G"k\��j���
{0��[p"O��&i��H�e��K>(�IP�"O�	H�F�b�.�pì�1 �R�c�"O�	C&/� �W҄I���3@/@@�<��œ�Q���҂�����
_|�<i�ûM�L{g��=I����Wq�<9cаH�m�4�4q�=���I�<iCK� 3B�@�Q?8�`!
�.�J�<	V��"2��w*R�y��7�y�<�f		�+��
�É l�F��0�B�<��D��k�~-����'h��c�%x�<Q&d�2�����b #؄�d�^�<9r
<P��ԋ`FZ!^椸���B�<0Kԫ��	rD�k���H�|�<a��X;H�U��-�p:�*�v�<���K�@M^u��Ĕ�*	�vbZq�<%�_�N�X�֩U4�h��C�n�<y6d4��捊)���!��h�<9�� V��*Sʐ�{�$�	`�<a3�ȃ!��0�(�,8E�]J�<iT�9r�l�h���!q�J�(�|�<Q0���;��ò@$zZ�Qv�U�<� '�IJuX���%U�jh��y�<����UY�M�9�
]�Eɍ\�<��n߀5a��b��AO�����T�<IQ�I(Ll��f&L��$�W�<�����@b�#Ӫ\��,�L�S�<qvhAT���nÃ<svđ�KP�<y���f�L��kF�0����c_G�<�qGWR�5����y�L9�!^z�<iĪ߆`�D� A�w��ڣ�q�<�����
�13#c���m��Uq�<�����H�#�Z�Sw(K�<�g/)綱�a�̼{���兏i�<F�N�}�5��r ��h���]�<A��ׄ��a��O[8{�@#�X�<�%o@�&�F"�i�e��xQ�U�<Q���9�ʔ�&o&j���(���V�<Y���+-�MiT��80�ZvC�P�<�7c�"w�
؛��T0qP 5%_j�<9 �} ��ԅC52jl��"#�M�<JQ}����A2r�ӐCS�<����`��N�]��5��Ra�<�C�x
l�enQyr�h�X�<���h���P!��':A}��B]�<����3�jA�Ǩ��5oh���b�<I6Δ�X��Ka蟂��	� ��W�<	��B�z�.������ȩ��nCN�<�t��
asD��G�&9�>�u"QD�<Y�BF K؊����W �V����[�<�V�V�1�x�P�NH���o�W�<q�������/�1a�2��(�p�O��i�$(�1Oq���+��43��c�^�h6�<�4"O~��� �,b�%����I"^�w`W�
�'�B��o �3��up��Q��2$:!������$A:�� N cjՁ29hx* ���\��H�F�3�Z	��&�O���h'C[�5QsF̊�-��'�>	�BMI0eXd8U(�>���D�E^f�� �խ:]�J5�s�<!b��DR(pP	#@�&�)1���A�B��8$Rn{"�R�{�`pI�#A�$�OD6����͝�tL�#@��2��`�ۓHt��f[��`�R'_ENUB��5��m��e��^�<]�%D���?A��X�^V������}��6^o�5ڇ��F�d �����'4QOC�]���J�->U�@8�� c����o.i���qw�ʐ6Hd4�0�]� 8�W���q�� !�F�p>���;3�:����M�Қt�w+l/��JÙ��y`-Iz�<����Ѻ0�.��a �وh��μKa��A�V}��2O�M��Lh<yQ@��	(Q�0]�TaCS�Дb ��0!��N�5��0�q!@> �-`��ղY�D}s3IP�a����.h��rDG�
�lEp����<	B�gA����2���CpN��k��Y'��b����P@�5z��B���u��@	�k�;F-0S����aWH�T�'�H���,Z�
k\X� �^�9�X�L>�`K�2�l�-թ´q� ��'
��)�#�K�Z�����?nM������q�8K����3F�6(nXQ��'��MRQh��4�`��B��.�
�'����0k�-O��ڱ,ѳ��Qj!HX2�~����ɬ�ۧKx���UE�a����E�W�a�&F34��8EK]Dj������%|��ak��W���Q�&�o�Q��h��F���)Ek]�Cd���afY�z��UԯٜQ���ǭ�q�N���"S�s]q��y��%�Z9#�nT�6��M��m䪜!�脄E�(���)� �����Tt$�O l��J���2j배yP�E@ 1Ox��p�t�;���޸
Q�|��X6�ʔR���iU`}y��V9D�E��L�(b<�veR�CN��g�2#A�,��<Q@�AE�tuD{r��&�`��u�Uc�BB%��T{���n�ʅy��\�0&>�9R�
6�����Oܙz�iC���"��x#1��
h�ʽ`�L�!"��)�:H&�H�J����B�I4g��Dy �T��H�Q��P'c�q�*J��@��P�gLmB��7`��|y0kU�^�	6���l�Mkvʋ�`ډ�Q�]G^�`z �U
�r���Q?�P@��8X�D�!��R��ЬkC
�18�����C0(�(�) Lͺ5�T4CS��*8�"8�Rh�ʘ���267�'f�!e���$�'����}�	�bìq�%�Dv�V�#�hU}7��b��^zZ��� �R� ����@�7u��+�ś��RU<g�B3��yx�|� ^z�"�$h��S*
�m����Q����J�|���"4�vQ��퟇}�<��Ԉ\41r#-���={������I�h��%{� !�Vsh<1l�?~�  QV= ܴ�Fۣ@�X��3�
^v�[p-�
i�J��T�;y�<(�V<ؼ�`�⼳�h�7T���j�m��R�j����gx����'J��l��՝zDѥ	
�g9��" 莊KCN�Q1��\��$f�ڭ����U�|`�e�K��J��#@R��H*�(BW�X��	$-칱�F(T����`��V^F��vf��f�����^�h����(nhȴ`�W�I�0T�U�'�AQ�d[�[������2Tz�H{N>�ĩW2Uy�T;�ٖ#A�I��
ʒH�`;u��7b�Yq���>} �e�䮎,8x<
T�-	���W�w�!*�Gf��Kd�}x�@W! 2�,��Y?SOxݣ���r�jÃ���`މ����y��$��m�"+��9�fI2D�,�@aR,D���˜$Wy�����<�*t�D��eU�_6���)R-G��sT+]�Pv��t����yt��'ڶa��؇}t�ICf�L>s������ۀ|��=*q�
��|1���3Hb�1�Ǌ |��w�N@Hf1���Dk�����I�%��]�q]�v�P㟨k��P�(��UC�'LH��PCC�R���b�3N�&����hC�$�'ٜU�A#�=`�a���z��TH��E�m�T���kR|�w�S�BT�&@�6�ĕ�'FD|��p ���n	�Pϧ�yw�D�nӺ����'K0H��Pa�&�yb&ܤc=��BŇ;���c���"ki�qRfC(WWpȐ����s����b9��
�eF�<���Wa_a?�W���`@W��D��!J�w���i�i����DۧƗq� E��"V-n� <Y���51lq��'o$|���37pm�� t��>醎�*F]��̐�Ν!Zt�⟔B�k�F�$�3]��8�!H��$N9�v�i^�˱��,L�$X�i� A�0I�r�I�p?q�␈gI<ݳG��J�J���%/ � F$�|t����U:
�l�(BQ`F��;�H��'�y�/dN��T�߃29���&��yR+�1��q���L�x�#�'u���ᣙul��&k?(Q_w5r���\e1")ZH���A��R,��c� ĪgML�0��x�j��%p�Y�pK޷4d�Pk7��7ʀA���P$Lz�0�	T6m*���ص/� r�Ƌf�^Y��3͎�>�kD8t�<M��oڄ׮�� �U~R����Ms��/�z�pW�ҥM��U��/Z�0h ��PB|�!Pº�v��
V�	j��`��V�$��䜽K�.zs∌Sl� a���u0�����"0(��ae���\�B\<���T�jw3�d� �ґ*�8�$��]���'m���Tu��\�p&�m�ic.�p�b]�=�8�YH>i���0>�6���Ï,�p��Vf�J?�"��)x�	X᪇�-���Rj�B�'!�����h��[�+��ȳ ���؈��
DR^�hd#�)j5�ilZ�ށh���vX@���b�E}
� :���(H�4a
�X�c��,I��OBM��	Ң�41�tǈ�L���iU&Y�8	*1,S�V������ 5U�ڥ��/V�l814$]�^֠ps�'�>���D�(�tL�w�Q��)8wM&�Th��h��xfy�� �M3�J~��p��=Pg,h0��`:Q愿l��� �R�ِ�N�jM;���S�Rl�Љ��bq�d �':�@)e�OH��GB�z�����狪U"�D�δ��P�өR޽a�W9�i��<�d�<���E��b�`���wصO��耆�S�`�6Ⴙt����+�oz@)���o0�3ǉ@k��	D}�!՘a{Nl�U�_�t��d�����-_�0�Cp�֫&� �R��² 8咅O8�n�nZRn�郳��4E�uڝc�(�R�蛽=RUs$�'�����(O�HCv�Ӵ|�d���Xm����T�A6b	<A�7+@�o��mZT��l�
P�&Oi��n�?=�BŢ��@��C/ �M'�~Rӈ^���f��tP20)\�Rjh��5��mT� �`��%��Y[�&�Y�<q���Iftz���7Qb|���鳟I���v�Vp��Z
D��a��?�-�����b��TLRfς-�� �B�S)38>��D�ݙ��)���q$�ZSC�=Hyơ�1�^3j͐Q'j�'�$��d#�8?��Y#� ǻ|K�V�<�C�4a~���D��*�.���9��e[V�8{D�4�2�I�|�hU�0 �bgDvS`�J���&�����99�% ��Q�RS ��q�H�[^����Y[
	C������U%��<�= �呲SQ��1iH��y'�c.x�j@�8F��	A����Px�)��y���2ta 6��ͫ'B����~��j$!��4����עE�j�D���,)B�YË;}b*�#-+���iƂ\�܉���8�p?�r�H( ���J^�p-N�`Y$�q*�)3��Rg�U�sK4L��Zgx�@���P.x���!�r@��/3�_l�@%aÄW� hH2	F�H�"p�e*9�h��እ/P�)�Z�&c�O,#3��-+�Z90����u�5�OlU��� �2����`Κ-
��!4cV���0|�&�C�GTQ`5ē;Pv� �"Oh(�2�Ƿp��ԙ��Όu2��A$� +drd;W��YN���c�AY�':�qO -�Ӫfan�[�/V�`�� �'�j�G�:Q���#�ک_�t�Xi��b�D�[��Y�8����U,��԰=���	N2����B�x���0�I�'$j(��[.���"S�Ь.'��I%W
>� ��Ԕ)���t�2!���(�3�d�]I�C�É�~��I���@�����D�T"�*"�y��� �:�k���7�y��$HQ�T�F�ٵ��D�WJK�jH�L�L���Rϔ�X�q��'�@5��a^�$m,j��ʎK�V8#�'��\c7鎜f���_.Qs�u
��N5w���a�n�z�L|ɶ���-�t_R��ȓ3(�X��,��H�:��d֕7t�q��`Ϥ$�ь�2_"H�GK[�d�^�ȓ-� ]��KX�=V0IY��e�j������0b�>-�j��' �b
�U���R��GG�E�݀�%9`����ȓ:���M@)̘�t��5�l(��B�"f"�[�)�֌��4j6��⁑4c�Ҙ��拍�`�ȓ2�t� F�j0�g֧zY+$D�P��v2�:LW�M%N-�te/D�pC�I��)��)���GqX�JqL*D�$���%Y��aad�,L�
�[E.&D��a�@Ñ7g�E{V����HIR�:D�|��
,�ꑀ�)å"H�홠!,D�DbV�+I��Cj�1'Qƭ��j6D�$�cR*Z��pbs ;Fz,�bB5D��!RO��lx�H:m��h�I0D��i���1�`:v��?�qXEf-D�DشNU',�\�"i��b��j�(D��SF �;f��&�Y@�H`�$D��#%.�=T��ԙ%dL�B�����#D���D�%=3L]��F�������5D�,�u��l�	S�YV#�A�q2D�Ls��ǯy�B�bCA��TYČE�,D�P���A����AGC�@xԜ��n+D����HO�)�������x��
u�(D�܊�-
�J8CS38��P8D��@�Z�8�N�jI��y�=D�� 
yC�B�jnj�ᔂ��CR�a(b"O�<�H�(≮X �k20q�"O
]X�i�S��i�REˠ"���"OB��W�V���ܥM'*��5"O^��7���r\�Z��3.�D��"O�����}�\�r��:�R��"O�1v�Y#t��yG6'���"O� sMZ�S�d�`'e�\���Q�"O��j�<	t��ӳĚ�.��T�e"O<�!ר�%b����Mϲt�=p"O�!3F��X!��ˑ�<ʲ�Xb"O~M�6�ؿS2� �lYϤ���"O�8ʴ��-'ͮTc5�� A� y{�"O�[թͲ|�i[�おq�@���"O�T��oC!{{��Po۹fɢ(�"O<tSPF�e�$�'.�C�Ԭї"Op̀c��%~D]��-M�z�!C!"OM9��,��y��)��I�"ON���G.h�T�AJߏ\j����"O�50򢑤^�r$`���
(=sD"OxtQ�� )�N�Q'ISF�H�E"O<�s�HP�o@�Gik:�*"O>8��"K6-@z8樌%*ԡ"OU�!��(FP�P��Ajdps�"Ot�(&��"Tz���&V]Z^��"O�)ȅΒ/cn\Mb"kł)4�y4"O����)��2���x��U�)��#"O}�kH -�X���*}�5��Or	��i>�c+l-���OG��$Д�nŚjD8u�� hbD�QJ I1�,��	S>)�2�&U���vF-'���"�t!$�A�U����'��x�t�i�ɦ˧������  ��ղ�$R@n�/�Mx@a�(�b�Bܧ@�"��Ā�ⱻ0m�-eD1���,����i�n-�0�9��=擿v�h��ՄE����Їc>���O$� RlV8l�<�1�O��@��aׄxz��Dnշ=�T�Z-O��R�R9U���ZM<E���ʗH2���$�(D�L�@cgE�~b�O�$�F%t�|����#"�,���Bh��x�oO(jq�=*�B,N�.8�'���%>�}:�FJ�bl⢭D&i��;oSiVu��[��	�4x���H�:��I��'iqc�(A!i��%�wn�G^��r�OM���<s�t<��'4��>Ŋ�@
n��0V�K{���VJ,(
f���L3a4�p�'J�h���݂�:��)�$]f�y'(�uK�dX�j_C�PI�uFw��S��%���9�������%-�m���AsEH�-�
Y0S�\Ӑ��ƽii�5O���S��Ϙo���9C�U�Q�w��>Z����>���!�0|�"�� Z��P���<5�&ݱ@	�9,s���O�I$�΅J��7��O�P����12H�'�ɰE�����24��įps�S4Ϛ>\�)�%b�i�&��?S��-��$_Q'nE�h���;�h�B�S�OF�����h�s��ͱe'�vdO/n/�ŉ�yʟ2�?}�2,X�w�QgI�2���pӄ�N>"dU�oVq����,0X�
X�Nl�̉h�^��I<�4-ؓ1�D�8K~ҜO���)}���&ڶ��s��3B���0д�0@N�=Q�ӧ���$̤I8��Qs"�� HE��!w-�H��N�5&�#�l@�y�ҟ�"}
�@=��s�@�3c? ��.H˟Tأ���9;� ?E�D�� hbu��D�^l�A��T-b�� ,�l���'��VDI�v�����%�%�*�g�<�/t�zx�,�9%�Eە`�e�<�$��ii6���I�O�<�`�x�<��i�/����(; ��pP)�o�<���h��`��Y�$uPL�v�<��ԨyтY6f�0_5�0�k
v�<ٔ�J>��E�%.uU�cF�s�<�!A�F�t�@�$Z���%J�<!�FM4%���Ӌ]�V=��jH�<�vh̽Q���
�U2� u����X�<�̒�TH�%D�@��%C��X�<1���,hv�����y�ꥲ�gW�<� �+��4"ҬHf�	�0X:�"Op��2���Aw�4���ԕ9��p�!"Op,�F̍LQ�-�q�I�iLz]��"O�E`��Q�)���rd�L��"&"O
0K��A�nɎL�`�]�j�-��'ڼ<@a�H�J��H!�@��;	�'d����cV�=^H�b@eTN�*
�'z���%���:�j�u���(
�'�
����Օ3���9�ƓgQ3
�'n0f�@�o}������2�4X�	�'t���0����:$($X�'x���B�F�1�B�5K�H�'2��q�߲����G3�@IY�'��x�c�W�f|�3����D�h�'|Tuy�Ѹ9yp���kJ�d���'�H�BJ�5V�x�p�ݮZ���'��0⩊F(�c�U:w����'���d�<>W�x�'&�g�C
�'���S.T<:P�����2�*,��'=h���� ������'.2 +6��t��`PR� 4��'+�a��,B�y�x+q� 6`!
�'a����&N!n��@��Ce�5#�'�@)W#_�2��	�'�ڌ;*T<��'�P�2�_�Mx��+�fW��B�'{j|�L˃]
z(�h5^7lI�'%�@@���
�F!��K%S0Dɢ�'8�ʄ��8�P��n�-R:=�'���A�H�$�f1���O�4�.M��'4�$r��H���Ȣ�X�9�!�'i�$��۠�,:gj�0`g���'m�(���:6%@݂�Ώ�*���'T=I2��	�E�ň 9Òq
�'�(�r�B�G²@����*di�'���B2�#p ���'ր	L����'���䉈� ZbD��u��,�	�'J����A��(h	��i�F�q	�'��ňWA�[���t���^)T	�'����o\�[Ċ��l 
Th�
�'�Aw���{龀�@��JZX9�'P����&u 
�`��?l��9�'`���0�/i$i�R��1n���'�6���
�&}��Ɂ�u�0г�'jِ�.�%i�:d��)J���a1�'5��Q�Ŝ���hת�Ϩ��'�p1A��0����.�9K
0�'�b�� �H���8J6�P���	�'|����^�H�-jEG�J�����'� ĩ�#�hN$	�%@+v\Y�'�XP�#h׀_�P˵�1��)��'�"�� ɉ@�i������	��'�T�灉
.]yjӯ�$���'8����Y�:��zh���hػ�'$"�0��+B�L�i�i >����'�1 �FG'd\�r��H���'� ܁glY�P�f�Kf��q~���'�8��-�_��r"�!ZM�+�'˰I����y��L�Pjp��	�'��3u�@�t	 ��C�Mw���'K2mɆ�Q'q�����ϱH벱�'�B�Y���}��sC	������'C�\��+�
��!&���m��'�*=�a���՞�����H)���
�'���h�J��y�M+��:Ap��
��� "M�v�aB�#P��*dvBh��"O�I�"�V���2��2Z4���"O< 3`��J?���ӎx:��j�"O�$��*�o��ջR�
� s�"OLRA
�V����l��(��q��"O����d�U�t��M�;y��"O�@P����v;9c��?`��Qr"O8��F� ��!j�K�U��10v"O 0�RO��
�T��	
!U�Œ�"O�!"mE3}&�,�6'��U�F�  "O���3�6�n��RhY�L���p�"O��I'�ŉE�r|*��X�-�$��V"O5Җ+96��H'�S���;�"O��
&������$e��w���K�"O��q�u�p�	�P��$�2"Ol�Bv�?G�JPȒOۀFt��9�"O�9"U��#f#6�3 @��B�\	X�"O��3�JF��l�dNSc~�y"O�(x ��:)q�CtM�;`r<��"O�!(gn�6�u`B�=*);�"O�B�N.3lTY{�/A�V9�aJ�"OD<�q�����c�P4-�I�B"OЁ��M��Qv�8��9;�4*b"O>�5IO�(��)�s�A9J�D�W"O��+v)W<X�uE'J7�:�:e"O���Ԇ��x�C%��)�L�r�"O��YbN��p5K bHF0�yT"Ov-�v��' �PV�̲8�, �"O`��%��X�&@0Sc��	D"O,���7r�aC,�&,���W"OJ�!qiJe�Ҥ��k����g"O.t�юL�Iv��.,��4P"OT`�@�Ҙ&�b �!� �"����"O�U#��Y�0���e�8�>���"O|P;��a��
wD�8���'"O���a�1:�ɓl��	�i{B"O�-�eZ�{H�y ��8^㤌��"O�i��w��)h@IH�!�>��"O`8p@�80�f鰅H�-mతg"O�nKI�|*�h�P��8�"O���X;?���6GA�Y��)cg"Os�)ԟb���&�H%Wr�p��"O����E�QCb�u���hdD�y�"O��	���:݄ #�ʇ�O���"Oh�d�9�p�h��ҼI1(Y�"OFY�`J�/�
42��ڎ<"\!!"O��D�A-#y�D��	^� Bd���"Oj(�@�޻S�a˒9R�a[�"O�Ő�)�D���1a^�P�yW"O�E��⋴JJ��0�ឌj�rhb5"OJt�5��R4t ʚ@M��@6"O���� !�*\��Ƌ�5Z�̊"ODTH��Ѕ{��"��N53D�$��"O��keEE���	�"X^�hhh�"O�%*�
�N>��P��d��Rp"O`C�K�%G
6<�`���a�"Ov����X(xTT3R�S<�,���"O �� h]#%��c�A ay��*�"O$�fn�)lJ�)B�"Eƚ��P"O����^d���{(E�U��"O�X	��(M��I@�,3.j}��"OB)]X:���5��ԩC	��Q!�E+.�L���A�6����qί?�!�K%k;`Y�b�ށ|��)�A�+*�!�� Fl1��=4+$�	U��:~����"Od5��Z�&S�My0���B0 "Oy9C'C�S!**Q#�5~w>��"O�e�3e`.��"�"(J�MÔ"O�Q�)GJ�j�Kÿ�H�@��s�!�d �Ft1p�ת���Ѣ���z�!��1�%�D�.C�`�d�Z�)�!��Z:��ٓ��?p8� �E�<+�!��e]�`��L2AV�1���!�ϚE1��t�� S�� UA	K�!��Tf@��`��VS��t�3��B"O�-��K�l��+�'��v��c"O�<J�/b8��h�F��[����1"O��x�܈Y�L���/���҇"O����A�:�IЅ��p�Z,q2"O|4�@F���a��'����q"O8���ϭ��I�PB��4t��ۧ"O����;T~pF�P=t ��R"O�,RvΒr�����.tI����)�yR�Oy���z�،\T�����]��y����RZ6P��	�"@�@�&	ʱ�y"��&;�����F�m�>�B�j���yٻ2��hp6�٪d"�$�Tg��y�AT�Yy[q��1B���O��y���pD�C�vC�H��'���y�&KL޲x2'���g|��r����yB(G�P�Z�PT�;/f��b�yr��>�R�jS����n��yR�d�8 ��������Tjy!�'�<��p��� �Z	Q!��-���	�'�֭��Eߙ^������%���	�'�f)�%�e�%��*�105"�'!����dӚ���"חf��q��'2*�b�ۍl���Q�-,DD��*�F���
.t� k��F�9��	���S�"��q�fc"30	�ȓIzP���b{����A\��@;�M8D�Z,I�K����CAS������3D�x����{�h�e� 
4� H7�0D��ka������! O�v�B51��.D��3b���6�i�4�M9z4�@�.D�X���6Q�����LI�<	�5z`F.D��3��!Fp!94�Ӎi�$9�e%1D� '�[�Z�"���DN
*��l�o3D��cҽg(�}�%��5mʌDB1D��9/��*$��^�Z�����;D��q���v>ބqgd�2��'�3D�L�)D3����tEZ�9d����/D��0�?Q�n����~�ԩpj,D�Nt;`��iS�K@"��F����ȓ+  ;DE&`���nìK<���0���	�ˀ(�p�� ���]H�t�ȓ!EV@���� _d52RB��A�"}��3�����9�Fx�s@��0�݆ȓjv�c�^!U���fm��?3H��ȓ&�`pG�*Yw\|�`�V>k��%�ȓMD4 ��X   �  �  y"  $-  �7  �B  N  �X  �^  e  gk  ,r  
{  N�  ��  �  )�  h�  ݠ   �  [�   `� u�	����Zv)C�'ll\�0"Kz+�D��`���b��$Ò�y2�S��y"��g+�Qے�Ǵ^�ֈ�2;de���L}��S�(��k�fY�+���\���
 (ϲ�	�J���pl[�=�@�� -k������@���H���3�Xy7�΅chP��;n��ؘ���?�#(A�}���8�&�6>B4�����=/@ ­L~B0@����> 6ퟛ����O����O����<�J���bX�E�UR��ףP����OE�����'���3$�*��?��u`|�K�*@�V�^���D���?a��?Q���?a��?1`ş�тB���@c��0 ��� ,v�Qv�S����`c�L*O8<"Gă��'t���ґx�#��ٚA�<������<����٘A�ƨ:�H��1����w��)�E�Ͷ#��z4��K�kxӜ���O��$�O~�)�O��'�yA��]�P��Ћm�@	k�]��?�7�i�6m���;�4�?��iR�A*���ڬ-͖0]�)��D,&��tQfg[
*
�x0��A�'g|�tVay�,��I��R8�]w����q���e�	{�juZP���Հ�p��Z�b�ۧ�mZ6��Ц��4��D;��( �;N����� �̭֘�Q�(��(����zV�V$k���6�@�4e���i� �
u��jߛVIa���o��*^�+��_6qX��D���{)��BHHr��j�*Ԯ�MQ�iݮ6�N9\�h��j�^��؃Ш�^BZ���ό�*Ian��'��I"phT�[�<����P��o��M�6�i2��
`�u-䕒7FR�CBH�geN�]g��S'�$d�"hpc�W!G'�6-7>�D��P�B�Jcl�R0�����D8��8j�.�Zd�^�&��2�K7���vB�E��U��ڟ �I�?1�Ӵ&��+���KÊ���x��Mͦ3~�뒅��eوq�	؟��E�����Iߟ�Q�k��A2�Is�"��S�ZI���h����O0Q�p��*\
J썅�	�gZ	2�Mؼo��PQ�����ݼ$m��Y$��؀��A%O�-iSX�P�.O����
�$:�v);��C+`�y;��'�r�'�'�B�'4��ɟ �gL�:^��g�%O~��Y�g���I��FQ8�T]���?Q0��|�7�'�V�2`Ms�Ȃ�]�!d������W���m�۟�z�w�Иx�) k�l�ᢚ �r���?y�@�-.t1 �����<	�i.���� l�D	�b�� i
��If�'?)�C_�Q�ƴb�.M�	����޲6;��hѓnH	~b�x�C�I� ��=�P����O\�oZ��H����h�2�r��I�?�Z�×l��Uo\��!��o�O����艏m��p���x�nh:��I�<�ڴ�%A�ǟ@��4�yBb?PLi(�h[mf���@�)�?9���$�	����Oz���O�˓��ڑ��o\�0����ZU4��"��6/%P쀵�i��|R'�J�)z�7��'�L���˟b{l�s��	Wx�R�̉�x�"i��Z�	*� Ifc�4��OE
O�l���V�� ���	(g�!;�o��t�'IF9��*̟�'�� bU��*5���C67�^���'�RP���j�g�ē�m��}`��u���$D���'��7�[ߦE%���?a�'������3g2FT�"ȹ8]bwH׊.r���?�����|�O�����iҮ>�V�P��Q�'��*틡d����훓7V�
Q�'�9�aˁ/Y: ��.���Q��?r������4z�����.fџTˣ�C�(�)�3�նf�^�C4���!\�D��ˋ�?�	GJ��j`�P��ȁ'�"(�	X��F�'1O*��3�C=|��9W�ֻ�&P�|��u� \mZdy����JL7��Od�$X��A:qΨ~>�sե�0{���O(� ��n�� �I6kK��
�Y�p�qe�������&��ӁL_��22�	|��C�B7DH���*�1cpN\&Mk�9��
�j�BY�c���kJ������#]������1��4�?�I�?y�ޝ�g�s�*�9t	L����O���O����Ң	�~u#0N��8�z����r��ON�d=ڧw���oZ��(+��XK�  ��i��\�7m�O\4o��k�ft�4�?Y-Ox�i���Dգ?pyEdӁT@�@��L 2����OM1vcD:���p�2 �ݴ��O�x�e�h��-#e%H]��5���Ju��~�f`��LE�uլܣ � W����g��k�^h�ӛ��0�DTyr�"M�̜@��I~��5�?���i���2c>I�Gkܕȕe`\"�@�`1 ����?�H>����?�)O��fl�v�D\�#�Ȼnv �Bj�o�'��&�O�6m�Oءm��|��^�s{����QK'tm�g��M���?���}�|@ԍɾ�?���?Y��y��]/.��墡��Ar̳D��+ku�@�S����� �O��@aS>�P�B��K<���
�pd1E�(�P�@��u+��C��o�>��p)W�:8�S�&;�Ѻ�!f�A2g��7��LA�$čU���!�DE�U��V��H�*�O�b>���O(��އ*&\���Զ%�L��Wf��$�OZ�$�O^��-�3}��#]��� `C�`��B6�K��?����vӚ��	Ŧ=���?��c�4��	 ��=k�M/��ʳ!N���x1P(`��';�'���'��5� ]�b�0zڽ�0����Ԑg/K.K>� Raѓ)fq��FC�l\G~�,|$��GP�=᰸�F�Þ>�PYC���mdȥ�A(�0_z��I��0֜��	2�`hC���$��S0@�Q���`���O��,��OR�v,�*^��Y��	�,B G"O�(�ӁO�8X4����+
�-ٓ�|Rb��$�<��N�!�f�'���Ļ]�-�`�B�U:�D�s/T��B�'�b83e�'�r�'��S/�.SRN���y� fL"��B��9�$�� �,I���'�欋%E�5	������vA�	�CJ��'K�!l����L$[�F���È�K���=�Q��柬z۴�剧b:p!��(V�Q�P��CU�G�^�'#`ń�a�xz�ʞ%����S]Q>��LԦ��r�-S��H3�,jn���/�%�M#)O�����Y����O�Ёb��'�T�
g�V28�H4å�͋br��b�'�b�+eu)�צ�5��o�˧���CKِ5z�%Ɵ/:��u�թ}n��y��P	ǲC��!�+zoPdѰ�<Ӯ4�FI �?�����^)��[v��6�0�*T�,?��Zß���@�Os�%6$*�1�c�	1�pS�&�U!���\�s&O��(�)9ў��I��HOLap�I���\�'"��(t ��!�O��D�O��d[*� )�O��$�O��$eޝa1 �:hܸ����2��ͪ�O Kz,�@"lz�!Î�}�.b>PH<р�7�t�b�ۖh�z1����>���l
�fpmqG*Y)hw�@�|
��x����c2�lC��A�%I�$:0�ډ�?��O�`It�'!B�ɱ|(�A����<:"H��G�3�B��"��V��*BL��+1/<�'T�"=ͧ�?!-O�ъ�-�3;���Ea�B�$3�1T��	A`��O���O��T����?��O��AJ�J$R��a�gJ��
x\�V���ut�Z�	�'G���ÒXI8�x�RL���%;E�V�`�
4i0���1�ѫC���i�
	�1B�xr�l��xX	ֱM�˲��8�b�#�'2�	a�'Vr4Q`�<��-
�'�[P����'�ၢ��2�Dݡb٦c��L>Y��i�]����.����)�OB�*�jH�w��U*�
4�J��S"�O��dC	���O�S @��(��CU$���P`��j��rc@��$�𲫑H&�XP'��V�0���	���1��IX`9Seŉ(#p�3'UIb1C6K��-�&��iN����7��s �Dʦ-�)Of+U�@7~��I�Y(	�B�|��'���3 *�΍Z��F�~a���i>�*��{Oz��N�M��T���G�N���I\y@@9e��'X>%KWm�̟����\�8�����&��)fg�ԟ��I�gT�|qM�QV��6㜐o����W՟��d�!��f��FA��!�Ʃ�'H�3�K��4%$�z��̶ZD�bs�<��m;RH��(Ux]�St��S�p��ʟ�E�5O���i�9���Z�kȰ]
�$S�"O,��Ӯ/��D�s
��R#f%r�ɀ�h�����$j����O���Ⱥ��q�B�D�<a'D�2����?������u���(& <Qg0�)�ȗ�4pJ�Z�LG�T" U� �5�Z]C�C�|B��L6���� T?�p`��A)d���O:�%+���	U�"���Q�P���iκ�@�f�>L���0�@�����c���l:���dY�
a Mj�S��Mcr^�@��Oz��-&��	��@�^�"Y v�_�^n�z+�ȟt�'2�'�?5ـ͖�`�,����2�L\�+Eǟ��	0�M#�iS��b��ʧ�r.�$)а#R�k�|!�"��P��e�[�nZ՟`�	ҟ����O��,y��A�~�`V�ߴr&%��ݕu���`�)[E@&���ި�Pd*��(O���&��F���sr�^�W���t�ΫN�2�V�4P��P`�v"����V�61C B3��^�V���A7哕C"��+f�ӊ|��;�':7-Mv�'z�Đ���7.��E ԁL	%��5Q�)|O�b������p�@��b���,6��(��#�dF�1��Sy2)č{#�맔?�"��eA*ܱ�녭C�X�.R��?��eɂ�b���?��O�e��&q~�bd��?8|����N�F.�Ӄb 4s���^-�,ˈ��Ϩ[�����[4�xY7o�6���bc,՜u����T��'HI�-kR��t�'������?��O�|D�C�+���q�Ā'_�z��|R�'���EB֑^1� ���43q��H�g�l���Ybg�	fu0��f�1�?I,O~�[��ڦ��	����O.4Y��'���*�K
C�TD�'�ϛd�ԩ���'�2+��B�"H��2*2�6�F¦˧��	%, F�@2�y��*1X���UZ:���+�r��5��"I1�M���D͏�Z�R�3&�)%�0�`�Oͣ���^%RK��'��>��	�2w@yT"	9f�ఐ��-p[�8�ȓz��T l��P�P@ΒF�<�D{��'��#=��d�B�<a��0�D��e��V�'��'�����G�)���' ��'%�nW	12�1��e	������6|��qEQ1:J$�C,؍;"��r1��UV�I->f(ҁ�2$�c�nGxM�B#λ'.ʕJ!FC�FH��uf:擮�ēp8�A��&E��U��ML6��	z~r$��?���hO +��T�#��z0�I�O��D ,1D�L1�Z�Lή8h2l�e��R��<A�i>��INy�B��NF�x�r+@�v��ZF�L�M �Qg)B+���')��'��֝���I�|�S)K���J�&��� �����.їb���xmFVz�`۴l��Gy��\%�� ��Фh-̈́�T���CvLjQ�j�L y�*_���j"�jӢy���\D�$�dࢋb5c�&�F�(����2r��d�Oh�d2�IH�O�\���lZ�`���b�~�KIn��(�<�q#�0k^����&�	c֍Vl�I��M���@x���O�"HDN����$$	~D@8뗊,���'�z؈��'��?�<QCwI
�h!���e<��|I�L˸U�����XL2���,~4R�N��(O�+fC�H#�9�V��7-����i�4�������K�d��C֋{k�IB`hÇ�(O8p���'�6Mly�A�.[P)�2�,B}��bR�L���0>f"ڄ{G�;�&�;A=R)���o�� ��7/j��H�
P=h�a�-(��	uy���!(3��'��V>}r�'�0��LԒ]�H���#n�N�@0Q䟬�I�t���E��7����6jY>]Ɣ0Pן@�BcJ%�5M��$�d:5#ԅ"�4�'쨀��K <SL@G��Sצ5Pa�.��8��x���� ;�`�L
Z�Nv��	���F�t8O����o�.��ҁ6n%�`w"OM��n�3C�uq!Sc6�E#��	�h�bi�-��.����`��&�n����'�2�'N��ɚY!��yU�'<��'8�9��`���X�h�ψD���&�^lty�Rj�u��AӢ�|}1�,$���A��*cq�DR'\|���僵,P(S�!�=!�Iɇ�Ġ'}�b>��L<�o�t�>������$��-ן�'.�I��?����� a$�q�͂q����]�]a�B�	���F�N�%��3a� i^�Dޑ��S����'Le
�/�p�0 �gϪ~�=�1I9]h)b7�'0��'x����ΟhΧ��"�#ӓ.Ǆ��ď�<(�%��)F<'�ފg��	� J$"�~Ds����ۆ���d��QR@��%ܰ��_�r��$�@�Ɵ�!��Q2s� �� �܍�l�&u쁄�$�8�/P�yBf�`��l�
�'�8�ڴ���|�6U?=�	�<b�I:�Z�*Š�����6�&�����R�[�l���|��A��M��.� �f	�0�Ծ.|�ю]���]���DcD�i[���:,��<A��?��ᒡU(�Ir�a��
��arV��1�8UR���8K ��C*�Sz����߹��Py1�Iܟ0�'�t!���ݣ7W�hiE�Ա\�V�iK>y�c<��S�B�_7���1�Ql�* �?	��4����I#r��̷���Zw+.KR��$*?��m]ԟ���ݟ��O\����'\rUr��M
r� �;c;�t��'��!5:��2WeE9���sp�I�{s�p@�� T:��.3ђ�_�tm{��f��������!�%)����5���$�5^oxD�2��?b�f!�z��<�r��W�l�4#T�ZN.�,7����͟F�T1Ode�g�V.Nw(�ӧB��H��(@"Od	���9	�Rɲ�녻*^(8����ПL����G�"(�G
��b��C�xw(��O���O�d���� ���O��d�O�ݞ3���9�ba�eE�H�Nt82+�1:��ՙ���z/l|�)�I/�����Op���#��m�)�(	R6M����NXX10�.y�^�2󤓔^d���e�|
���z=��ͻm8]�gF�H��Xܴ��'A�	������O��=�6`�Z��hKRoD�Ns��z���-�y�E ,
|P\Rx}�l#G���?���^z���S���'�|D���$U�4��a@S�g��4�Ph�3{R�;��'/��'���O���'��i(+VL��J�<ra�2� ����$���ǝj��,
Sc��f���dHC�՛)5zy�¹4�,F�0HD5ZuaN3��$HEb�����h���Ue �� ��'|T�7�p������L���)�&��?����hOJ"<�p��:мh[v+J��T��D��O�<�6m�Qqli�"N�DI�Ȓ I�;�M������	Y���O�O֪nv`F:z��Uc�!pb�'%xaʷ�'�1�b=��d��l�f�21��1X�)���K�t�|!�V�\�����=`�F~֕E��e���K�MЦhR�ؔm�aSk�3���p�	N0k��L	0��r��1�	�W�`���	Ο �'���p�_�\Cd���_�BO>Q�����s*�-[��-���J`�	j��\���~0�=
む�&*�! ���;�����dy��q r�'��Z>Q	K��|z�&��G*@�(�΃\	�@�T#Y��I�J_��vf�?{� �uK� Yu՟"�ZI��z��̒HX�ԃ���U�F|�'�n���I̗s�̕Q���9
P%��g�"�6YB��%d�����P;+~!ą�0n���uU�������E�4?O�����07� �k����/�|aQF"OhT�U��!Y�<2f�X�>�IA�՟(�����4��m����YP�jG��[G��m�����۟0�v'>B����� �	�`ϻrp��p`
C1��,xtf83�4�%1�p$8�-��Xo�%J@H�w̧o�'L<����B<��C�ˆ71��u���!,��k����0�|�ZLW���O�O� �{b��^�e��H̥qm��Xf�'@�IJ���O��=���<]H�ܢ���<D}�!�S��y��^^����ő(N��)
���u����'K剢	)�ݨAň�:ܙ��_�T�� ��٘$�(��ן��	Ɵ���Ɵ8�I�|R���g�4M
`�*i��x&ˁ	�v��H�3��t�5�Uh���	�s�*�� �L�ܑV���}�b�#��(-N~jFM_��\д���M�&c�y�j��H>�c�jRDp�F� 15v� �GˑNR���ҟXF{B�	�EUrI���� b�8<�&`�=����D#�	)&k(]x�F^gD�p��OPn����'Ɉ�ˑ��~
��iyި�Ӥ�:GR���7��x<����?�V���?	����A��Y��qTJz�)��!�?��]��KdT�2��E=eK�aa�`2��C�P'f�:�
O0u�l�9�a��y���b�({ �S�|x�'�r����Ň �*@�����XI(����&�D%�O����ȥQo@ P�Q�45k�'�<�d�1� �`t�D�!VVp+��@�t��_���%L��H��䟜�OT�l!'�'����w��QeTp�jA�C�FUAs�'�RG�<#�Ȍ9խX�N|��i�k���'��i@�8,X�����=W?|�c�If���LڬD��@/,���i�AȲW��D��*J6z@��s�^�8'�5hj}�N�6n���'������?)���~�x�� ̱�x<��"ա}�v-j�?D��	��˙�4�!��LMSU�;��P��>����
B6�h���!<��@��Zڦ���ޟ|�I;-Ė�����ȟ,�	�������<U����E\M� ʶ�\�'�'�DT`�mU+��Ϙ'�����$�W2V��`/��Y\�e�nD�Hm�uqddأ�ԭ)�B�$+�hh��byRp��$p"���uvz�8W!Z9�z����l���Ot���'1�1O�詆j�p�r@�0�ʰ3@c"O��87��]\H'�T�z�d|�Q�����4���O�4ö�S���9��� �xj�hT-�h+#*�O��$�O������d�OR��cY�y���Y��p\Ѧ˛��^�+3n��,�BM���[�`�˱�H����E{��3d�R�F-_�3�� ��@�~�� �F�H0i�n��P��h���J@�[㎘�%+[#<R�'䈘��Kߛ���MG��E��-L��?����hOX"<� R�~
�)#��'��l��\e�<1U.��EN �f�Ĩ]�y� G�	�M�����"���O'R���!�@	(q�@t�%a�=^xR�'/ND{�'�1��Q�bɯg����7��%^vn݁�"ѩ��_	�z$�6.�#���`߆�(OP�ydH�ն��$��#����3�L�uɄ�*�`�2��y�
�81*6�תl|�?a�mA˟��Ig~���r��i��JpCz�*�/����0>y1c�/[���R֍²��=���x��p��{`Lh3U�*,�lk�
6�LY��py���Jm�6��O4�D�|�D$ڪ�?Qƌ#�4�,�#H0U��$J�?a��%��Asq�^�-��(�@����Y*���'9��xZ0iU�#�9��k��/3`\�'�`:AK�
9&����ij�)G��ʙ!E���ɶc�>>�=��#�=���R?I��h�&�.HY�y�E��?I����(P!�`B�	*V��%)�!yo��s񋏐 F��?�a�>mf��	Gmò¶T*bN�8Cz���O��D�O��!�E�Zk��d�Ov���O睒.�@Q�&������TD�F�0��*��Yr����n� K1%h��.�;|1��'�O���S�X� Z����QF�t	�$��DP�@#<9ZI�W�װo]~���7-\5V����N�T�q��*Q��#^�����-?a�e������V�'\��&D�':ь�j���&�4�8c"Orx� �9��YbMNl�p�SR����4�����<)g��1K"��2V�ʗA/8��4Kӳ��Ze���?I��?���K#��O���w>EҐn��~�+D� b���`�J�"S��j`�dc0�V)����K	62,Lڍ�$
�k@PA�<+�L�CT3M��4��)	 2��@�P
Y D{1��e�ցx�`N��k8r枚
��u+E�Y�;V콛��Ο��,Dl��ݟ��x�5�X��Ԅ�ȓg/ �E��$s��|G��%ָI$���ش��>��������N�3<@����G�s�i��?�?�(O����O��d �'Ȳ���
�8	R%�P�R��˳�ʺ\V�$U'��`���'�>OvY��Գ*� ��R��u�:�I0#^|f�s���c��C3+�<�$�X���g�'�89���?	�ON,�	V�rb����9F����W�|��'���a��]���A���/T�|r��i>Ey��V?��)�nئ`����*$���	]y�K��U��)j-�l���	"���2e'� &N"a$@�j��O"L��v"
������E�)�'6���ф�eve�b���.��'��<�qɩO[x}{�`����������l�4��:|4��@�����j�t���Of��7�'�y
�  �#�ԌI�h!�P��4���B�"Ot`��O�>y��2� ���@!��I����ğ/.��0d+��1o% eAF�˓�򤛋c��d�O`�d�O�˓���c`I�.P�8����E�00�w+K�4�,Lsv�'0��+˘Ϙ'����c��Mf���f�M�������,_�Ȫ 
�=YZ��	�ʘO:�A�7l�>�'�C�GA�����*
�dțg��֟�'�ɐ���?������uFl���U5?�bL2�h��B�	' ���S�A�65&�ȀН��d�O�YFzʟ0��mC"@�u���[��G�Bw�x�/  �?���?)����J(7�b�Kď�&md�l�?[|���7��sܦ�#P��z��a��	1D�t$[�\U�X�S�Ox૶�kӰ<�!��#Gd�S�I��M��0U�I(SX^=�T��r�),�*j<��C��O��1ړ�Oap'�=G�*���nI�[Mt�'�1O@��RF��KRͩ��!*�=���|�>�(O:i;��y�w��Q�b�S�F;@��(��{�*�$�<���?���l�l��g܆o����m�M�d�y��yS���@v�3�!���0<IdH�0@&�� ,�<ml�2�ȟ�1fz`�ì2t�����F����I<���tU�Of�&?��F�yd��B�;jb�st Vh�I{����ș��uStiޚg�-��7�	w���4$�OlX�"݅?*z���M8�h���'4�ɀh�¨���	�|���Ƥ����p��p�6c��VE�8(��?��+
[\h6��0� Ö����M1��-��lQ�F����ß�P��&�1��a8�#S����$禵�)�i�;9�V���l�
7��A��@�@S�	n2�d�O¢}��'%�A V��<�u�H�s�)
�'5��9��4(�dmB���/"N
M9����O�Fzr�	^CVLAc^<.��$���]V:�	Ky2$0U*2�'-��'R��m+2�ya�=�����"6�� �g|���g>X�H�da�g�B��y���X?B`>uKQ�UE�Mw�Ԯ]\M�.CT��_̧<*��ȳR��P��'%� ���ƠB�r��f��O��B�e���G{.�<�(�kV�ؐS+T�� ن~�!�dɼ�jE1�K@"\��.��=2�'AZ"=�O�剶!T|C$�K�ޞ!��gȳ1���x�%w�-D�X� s�D�&P3E�����X��u�������y��<�:ZV��?r�8+ĭF�?!�j"�?����?���V�:�r5�Շ|�Z���c��ݵ�b_L��p�0���"�j�c��!)�Qځ˞>Q���b�4z�"�*Yw
z����@�4��bl�39�aY�����X2�'a1���a���_Qh�zaÝ���P�H��I����F�g�0�R�/_5|����ĀJy"闘O�d����ß�T\:w�2��d�i&���O���|�Չ�&�?1���V�X�S�� ��IO�F��R��-�5���ͦI��2s�5r�V�R¾?��|�!G�=u&}��^x�:2���<Q��-'|Mچ��8�*u�"���
�>�yq��"D���FN��r���&n�0ZD/�O���(?%?��'���&')8��&�S0��h�'�nԸp��+�4  �(O���ҍ��HY�Oraڢ)�7 5�ƅϰ@D(���'�Z����_*s����V�'��'Ib�O�"(Ӽ%���P �r���'t����ID�T$ڀ���ŕ&��sTk�g�į:����D��˂�|����U(b$=j�)��,��jL6GM�����>rc�<b/�ຠKDl\"��
΁��I	���D�O�=��'�Ҍ��a�'Ҏ��v��@/���'�J���o�"0F�Y�ʍt*t���w���SџL�'͖����-XT	D(M�J�WAG/�T�q�'���'B�O,B�'��I�4#-b� $��R]Z�cN�@�j%�怍�?��k��	����0�K�y�'<b-(Q�+*��S�
�<�݊uJ	z`~���$�,Dt���(�X�H"?9�C~�7E�@����ö8o*�
��٪A���8ړ�O8� 0!�t�3���.�J��7"O�I���	�y;�\��̼ۓW�X�4�?�.O8y��ÀH�T�'9�ɟ�RF8z`��qyJ��֍Fe��8�2�'�R�U�h�481�U���k�uu"ѯ;
"��� 虆D��0����-�G|B�I'rؽ���ׄ��ܳ����a{����&	wL�K�n�+W��z��">Y�쟠�IA̧Od(ls3�+� ��	G�r���<i�[���ca�Z:T[�X�Й5ղ��	&��$�*��&˙�#�0Ⱥ��͵8��)� |��ӟ���Z�4�7]D��'J}zp�^Jqxe�_o��:��'�J	�rF��G2e�$Ȁ;'G�}BsK�@:��D�E��L�ED6X��!g�L��y��	e7���F'�@�P84��E�8"}�t��I~�樑�=�<��G'��<���ş ��b~J~��O� �R��.J�&,�s�ߕH�|��!"O��h�Дnt(������6¼<j'�I?�ȟ`l�AD�x���X�"WFq����O���OnY@��^5���Oz���Of���OtP8��Qc�ܴ"D�?I����  K�5`��0ȍ�B@RE����Hz�~�O�m0�Kݾz"R9�d�ީx�&9*��НW��$��r6%�����V�S���'���h"�7[�aB�KXv���O<P�4�'"���<A /�8�� H�����dXbc�_�<�B֟zyB�y&퇧?<��%�Ɵ R��4���İ<�P�7� �� $޾�՘�S.U��q��?�?����?������?��O��Pؠɝ�:����
�ld8Z��WNx�i��9�x���@F�e� #?9�D��{�q��I#&>�<�7
%xܰ [�C	9K��k!�B�InP�$�	J��D[�S��4! ��$N�\���a�G����-���O�)$I^�(e�`�r��l���%"O��q�F]<7n���2�}�[� C޴�?A/O���#Zr}��'��i�W0 �FӼf&��A!���/e��'u�,ޟn�j��A$!QYN��Rz��ꖷ�BaAh
��4���-r`�J�E�mb2�^O�\c���x^\M1YwԞ��6�I,:.�+ɚ�c�`y��Ă} p@Ó�|���?���i�*6-�Oh��c��,��B��Lm����V� ���O��O��S�Ox�Rӯ����U��w�f<
Đ|r�i>Ac�4%��v��&cA1+��PT��	��I쟸��쟜��ş��I��D�	�|"���+WLܙ�ŋtf���}�'m��}rBkȌ� �Ӡ�
)��)q� �`��'�x&�����'K���҈AZ�Δ2t$PQ
AK�wrY�۴�?)��
�y��N��?������yR1$뢔�mM$LPRU�qO��Q,�x�Ѱi��ʪ9r:O
H!5П�^wYL���5M�)O<v	�!"�;x����d�8^�����O���o�����?��������y��l��P�#W.u��u�V�=m �8��?i�
��?���'��\A��M��ɶ�I�o�hKA��>M{*LZ��-'7����7��D�O��J�\���'wb�OtFa�P�Q6ˁ�`�X���"Rz����U�dLr�'"uȰ�'�^�d��`M��i��q�E�@���m׷b�.����Q�:��6mx�Īf��O6�6Ҋ�������?��'d 
aB��ڥsn�#$��%���kgȑ�y�׻�?��e��n�OR�I8]�>��S�1Ӈ�,�X|�u��3jӰ�!�h,A�����<���Ο\�I,��?��K6p���B���a">O-�0G�i�d$�8OB|��)c�FnZ�?=���?��Ĺ��pl�L(Z� �O��v+�1�$�Mc�鄮�&��ON6��?�n��B����iA'-e�XVH�.(-d<��J�;	P��ȓ):\���T 4	�}��@HK��n�Ο��'2"�'"rY�8��56 8�va�wK�YAt�h'.��������8�Iß��O���'	�'�D���S����v�f����n�V�D�<���?)��?����?����D�#�@3eH\�i����t�iD�'2�'A�'.�-�� ��GC�('
��:�$qmӟ�'��?�H�d� ɮ`Yl�3A2{q�X��{ӎ���)���<��';��rP"B�8X�0�qЁ?��O�����d"}�ON�~�DM	���lZ�#�8�yb�o��1,R��B�� ��y�֧~&�S��ۨ�ؐ!���y����,i���b����@R�y�+��UF�`ЂڛW9���;�y�#E< 3Ve����9�&y�w�֮��'�q�v�˒Tc� 3�ώ�+.���hU�s�v��%H$$�"�;��Ԫ|a�娵*��kK>���-�&���e��s�az��߽�>�D@��H�wH(��'���G*��|�p��t���Alt�q�\�r��X*��ť�~L�#-G�y:6P�l�7�����nű1�Jdz�����0�-��7�����+J�MB� ��k
��2ts2��,$S�9����Q����~�^�b#�34z��Q�_+N�41xd��	&b�Z���Z2$�{�b�ش	]�Q��[�?Ҷ�F��,Ħ� �'=2,[#�����6/1\� ���	�R���i�Iw�2��C�'O~�X3�^9@މ'LD	����b�b��b� �V������*���?�2s��8�D���Rs�9��+�$���do��E����ܘf�R�8ti�F"U� ��	w���i�a���c�I	BjxxRANB�c,�x��m�Z]nZf��;a�P)3���W�@r��2T��\� �io��'n��ʏw�*����'<��'��;+T.LHeG�t����? 򑲣#Όw���H� �
-�@&�2+U1�ֱ�'��Y��~h���NC8�&�9�6�֤�=0L�S�>�θ������������w#��@�
���{IY�N26��I�B���x� Փu��l#d����yP���y�S�P|`J�*�?�0�{$����~��'^ "=ͧ�ēԌdJUׇ	���A@�+���g�'�8���',�'��Iw��Iȟ�	��*��r�T�\Qa��4l�h��Э����m�q-M��=1�� l����'e����G��
�ܡ�P��pT��Sׅ�0��=!w�ƚ��1KD��M̜�BSnA2Yn��	#K�8!���b��8�OLN�<I1�	t_�ч�^��?����?QO>�,O�O"he;��MY"��S���\�('��<9��#՛��'��	�2��%���7�Z"~EԱxFm/\�d �Q&Cݮ��	ϟ�H���T�I�|j��۔�����)ѹp�f�� oPB`�/ғ!�vDK���N��ч�8H�H���%�2Y����ň�r��k7G�D�֑��C�x��i�!6O�,B6�'�47�[?AdL��@6�8Ō/+"U;��fܓ�?!��TPzt���_��2fG�2��uDy��i>��F���0Ht��`�3g����-�A���<��bX?�	����OHҐ��iB���[�,�^�5��2Z���I ��Op��i����fh�$L����\�;,��!c��@��s�é҄#�Ɋ�:AƠz��xr�Z9��R�ǆL@6�ؠ�e�q���#\D�	��]��؜�c�ߛub4$���c��O��D-ڧ�Mñ��"S�c����2��+�,!���dG�(+�C
`�l؁��-p��E{�O5��<a�@��T�PQ�-�<�@Q��]0�6��Ot���O\q����J����Ol���OGE�j8�@��Ʋ�p�@`aID����C<=�b�nZ6a�p�b�HJ�c9�I,|8I�bZu
2LrI�P�l]� �TA@��&8-��t0�-5 ����U>	[����y�F�*G���REC�A��H�V�������<	�F����l�L<ɑc�9e/�;aК!j��{�'�ay",�'lk��S��.rtF�:�a\��~��'�R7m^禥'���?��'=xA��'��w��'%�\A���E�X�@�Ot���O���޺����?!�O��횕�Uj��$�O�n��F.A2n���ؕ���|5±pv�Ȃ[�џ�R�h �]1g���Q��-S�5��T, '�%�����D��W;r�<��	����;F
��`��+��?���'����l`'�@?�Ȩ!�8�@�7"O�L��M�vV1IQ ��x�@������	Ry�EQ�9�7��O�6���++��2��42��}�r�T�c�h�I蟼��N������|
#������q.��!�ȑ��	�y�q�E��4���-FKTDT锦�n+�<�DD��t0���}8t����+2]6�[AO�
\�����-�&OSbS�cS$!�H�X��!��"�H��	���ɱ6��pɕ̏�r��`[⁚?.��B��
%�p�������-{��Y�~A
�<���4�j��ę#nI�SB̳q������*A��O�CQ.�����'O�S>$;�oZ"��I��\�TN����,S�N��$����?�Ձ�X��ś�/L7>vlT�T�Rl"�n�({�8�4K~s�+0��Q[�Y�?B�$�L��+�._��Ѓ�V.]�F���V�K�����(،��V+^�k)�,�v�[w�'�T�Q��?����e�4ū�Ń�JB�&!Z���<�E�}H<q���&@�F?d���Gx8�����]!w�:8����W��5��P**8�m2�4�?!���?A��[�p�@A��?i��?�]�]?XjW�G,[�̕��NU����Ć�<DI|`�f�i�>a c,��p��ӭи'����b�U�	ev����h�6�1�I��հa�0sY��8V�C���OWfQ�#�O�AL���@/����B׀c6mGjy"O��?ͧ���x҉��K߆xه���4��	�1��';"�'��f�Z>�+dB�R]�t�ʽ$\ ��?��iW~6��OT�nS�d�O��S�>��t �ghȻ�Z%F��$�eM�{L����?y��?Y���b�D�O����)�'�ɛC�H4P!���Px��k��؈u�@$8ʟ'��<I�'A�q�d)!$�I�u�(�a�W�4ȸ����	ڨ�rU��(ئi)�	E�nM��3`u@(+bkڎ��'͂gj N��aM��J��Ȃ&dT��?���'3:��Ǡ������M$?�H��'�LQ�#�_}ذA)�>���H�{�`Ӷ�OJ�gI��E���i�1NJ>���y�E_ToT����?a��i-(��?)�O�p-��b�	A<�z5�ɬ5���j�P-O�%��ǎ�{OV� r�%,Od*u�O&�:[r�i��]24Bxc,y@��]92�(!�4&Q&ǰ<��,���p�N��0��1!�|�5NتL0Z�I$�*D��G R�{@hP�X>gV��b�"ʓ�hO��þH�D��#�p��0��� %T8��'o$��J�m7
�o�˟8��E��G���?�W��0��0'
�#༜2�Ey��'a ���h�4z�-�O�@AQ���{Ҫ����'�ôa��Q���]8�*�p0�x���
l��f���ƴ����=J:�U�$���� #��(#Ӧ�.V�(c䈃]��,RJ<a��ڟ {�4j��>y��u1)�E׷O*�1&��PN��DyR�|bQ�Ʈm~4m������8X�E7ў�S��M�ִi��'�)д�H-' ���U�ؕ�D���
�¦!�	��	,~2��cQ�Hҟ��	韀����H:�� 9i���`��Y	 87�� =�D�ŭ��T� |pt�͙s�L�O"�dX~B�!ib�0!GٜK�x!�&Cr��R1�! fͱG�Z/>8ث�}�OӒ6MW��� ����T�k$�����DX�XM���˓�MkAY������O�2&�8a�%�!Y����&ωR�A�����hO?�$N��L��&5:��z���$��d�O��mډ�M�L>�'�R�O�X�L�]�%R���-��IN��k�(���P��ڟ��	��u��'��'h�5�B�+	��y�%��l��� �@��d���F�GX���'��`���#-�7j�R=��/s��h%H�i���.c�v�Tm�
	?����$W(޸'F^!��E��{��e:q��K�A� ��?9��in�On�d�O��O�7�۬4���N%	$�Bv�ۮ6P���Iݟx�	c؞�Pp
_o�&��0��;�iC�
U��?�Q�i�@v� �n�O��E�o�f7-�Of6�Y1
*��'��!alni�f�S?V��-��Οl�5@������|B�-ho4�eH٧m���*�'�"�Re�Dm�]�`���	_�:��۴v�vUFy2
۹�"A:��ɪ�ҕ!��U#����4y'O�F�B-@������fE���'ܪ���?I�O��B���H��nG�k8�x����ON��$\+ ޤ���Yz��K1�ߣ����X* �����G�Xn͡�ڃ;��#��ORʓ@�UJd��?!��a��-�
n��F.�
0̛9��!&��	�h��O�%�P�STRLp�k[?*P��A�M��T?�k�L�"B��ŋ�y���3�?�D@ ��1□��SB�,P��!Xz���LV`)��I����ν.Z�}PH\0>a^�'����OR�d8�'�M[#�S	a�d���܄z�P0BEI�5�!�o<��*N�i�\��d�
y�E{�O���<�Sjw�R��<"2 ��ب�
�0��iQ�'���E=������'B�'��;1����I��7זH@�+̳\M,���G�K�:0yr�ټ�Z&B�1�1�d�'H�|Ò�	>�(��ș�3�|e��&D.<]B`�E)1�^!`,Z-��O-�j�r����=*~�9���ݺzЦ���'u�I:t���4�P�$/��U2�+`k�F���G�`�C�ɀ\tb�P� ��#�]ȗ�
�<N��	۟x��4���D�>A�l���i�l\�Zf(T��
�0T�0]RL���'�"�'����t���|ZFcR�O	�
M�:��}yaiه#��ٙ3B��c�x� �� �~�Y��{�����lM���:Cݨ�!�U����V��p ��7��UN��)��sB��R�G�TSF�IߟP��ǟx�?Q����0Uv8�O�,V6��{4�p>aJ<�e��5u�4Ã��T�%�#'�RܓU1�6�'M�	"j�\܂ٴ�?a�4f��T`7�G�fHz�8Q+��D(r�`&�'�B/��"�'��i��P���P 흀nM�}a'��UHp�4�ܺe��Q !��{GD�*��Q�Niˇ@�Y$F����_�q���E���6Z�Y`�g)_���#!o��a@c��b�O�؅�',Z�'�A"w���h�M�h����'=�Y�T�,@`�I�C+�6)88\z�'RU�6�Y�_�5*Qǯ�y�D��o��'l�$��l�T����	��<7M�+l+��Qn���d�G����D�������!Gx�1�3��WE�l�r�ɣ��i�~:t-T����*�f�5x,(���c�	"ZJ�@9S��W�pY{�"�gqܺ�D@�2�B]��OJ����H��@c���G�&qSL<!�� ןl��g�OB�f�"�,qW�]�U����@˫n��C≊�%n�'k)�(������	��'`R�<�¦n�	�Y�:I�Q���
FN.��?A��yր�b$�4�?����?���Qb+|��a�s�9����G�8Ê`�O^� ����$��d��T>�9�{"Jބ���9�n�@@�U�,����X��� �F�4g�[��d�>aGb��+��@�D�њx��S-Ivz6͘Ʀ��	�(����)�<a�4"|T���*
�+Cc��F"�� ��'1��'A)�Ѐ�@�T(yp��#{�P��'Z�v�DlT�	%���M}I�#����j�*y�*Q�&M�!n֞z�~�d�O�d�O޼�O���'��Tԃ�xq��$;ƎLWb��h��i3��m8�S�H�,GL�dF~�h��~����͓^o��f�ڳ
���D+
�?�d�\�]�
�҃MqӀ�����:�O�� @��=
t�S�M7N��sb� }�/w�.�oǟ��'���'q�P��)$z�=j�4�
Vo4�O�O��E@2G[6<���+k1:e!PϞV�I��M�@�i:�[�⭖�5E[*��5ce���A9\��O�&��O�OZ�>m��W�bUq7�6<�zf�]�F�LB䉟N��0H�U.�@E��eRC�cB^kT"R�	�ֹ1B�#b�C�I�m34���X�g4b(X����0C��;r�P9��o��:����b��� ��B�ɢX��hӄO�P`(�J�	~�B�	m0�՛���Wy���K�:.rB�I��Z4)��&��#Uh�	wDB�)� L}J1�בl�Ӷ��7ݨ9؇"O���L�dRa�BU#�x��"O0�90#ɘ�����M��� "Oj��%$�-���.�%�0�#�*O�}8G���;�� y��E�.=�	�'l�as�AӯyD�Y3*�<:��	+	�'p���N�,
X���E!�30�� ��'�T�2�/��v1K�ܘT�(��	�'��2z��c�(� XT����4�yb���Jh���� �Oj��a����y�*Q8+���z
^�P��0���M��yb�B/;A�Iz�jL��Y2�!�!�y2��:tq|hp�@�<1���y� :���,I9;C����CZ4�yB�\��ꭰ�%�.��}� �Z��y��Ɂo�:�m0V�Z����U��y�^�Ti�7lJ�NB�; ���y2��%r�A�/�rL|�Q'ND�yҍE�s/N�iw��$5���kcC��yR�\!HX�xj���)Aw��z2S-�yB�J�w�&�R b'6��P�*ӏ�yB�*{��y#�V&,J�A�W��y2INz�,x%K�/u�(�Z����y�մ	<u��	N?k4�Z�gE��yR�ۇKO�\BQ���E�`�e�B��y����>�9��h۔n�����V�y�f�|m��YB�ϡ{vt��
��y���e������Ҽu���"cDG��y��[)A�:���
�\#�!���y�hʺQ!�i�vo�"?Pt�����y�f��$��J��&< p�@��
�y"j�7#�ޡڂȘ/���a���y�I�R�b�KǔY�zl�х^��yR΁ KD�U86�ͬY&6ŋq�ʂ�yre��zӚ8ۦܳ\��ir���y�@�1:���!с>7��a�����yB��q� qa��.;����yª�%k�2��'�x���6�yb�L*y]2��[ -TLc��yN��Ԡ�X�"�6�\�*�D��y���j��h�ˇ�� �cB�(�y��-Cdjl�1$�&{��goޜ�y��ܗPWFM��蝤w��i���ybi;Z5D9ZeƆ�lx�c�N�,�y�
6�ځ(E�	�iUļ�-ͨ�y�'ȄPd� �JdjL���f�?�yb�,:�Ab��Jo6eP����y�d�5J�~YI��
)A��Ѩ�g�-�y�E8������N�L�	���yB#ƣΞ�Qũ ���Y2�y� �)�l���K�~�A�tN���yb��	�(k%eػA�蔒!�_��y"%��\��є�/= q�\4�y��ڰ2Vl�Sc=�:�
AO֗�yҡ�5r�ȳQ
���s��K��yb��t�Ã�%�� �G3�y�&�;XY�EQ��:3��)�y�/B'��KTB�.�qi�N��y��O6g'6�ʰ���J��Eĺ�ye�Vjx�x���=Mg��&N��yB��aŨP@G:\}s�a��y���9���C$I/o}�h�G���y��E�3�~Y*��f$�L���y��� VR%Pf,^:O�AH�f���y
� lU �!( |��E
/�$��"O������?3�\��!�}��k�"Ol��'[7(�,�
�F��`�t"O0�ǀc�U�sEQs���2r"Ov8S.ƅ0R��(�
�Y�b�:"O�����4MI\�y��An���"O����J�i�L]%�E�Ve^�"O� ˡaɚ�h����{T�(`"O ��P�k���(X`A���"O���ƌ�P��q�P�Z�X-jg"O��A��	h���B�h���ܰ�"O*�b�^5F=$ �Ǒ�v-nD�"O�,��왟\BfH�0� f���#"O��6ǝ�_H�#�#�3&�2$pW"O�rq`��	�g�?{Qn��r"O�Cf"��N=E��O��v(!"O���֦�#K�5���:u���r"O�ә�h�bq/V�N��9��c�F�<���6O�^��B&bB�+��g�<��ԬJ2^1�R�Z
3���T�Nz�<�5Œ�:���:�ͅ��)r�<��lT�+�v9����X�1�F�d�<���62��]Z�e��K�A��a�<9���f�V����ެj��	E�Ss�<��`��{��s�	N%|�FQZ�OK�<apQ�/,2�r@
ؘPCP=zV�G�<)e@�3*�$l�dN	*x�r]�խ�F�<��ʇ�v��ɸ4$�)3�h�*�OJ�<�wE��Vd������,/�HMY�-[D�<�Se�;l��)7	+�(��Y�<ipn-=b�T�E�D%�L����o�<qЬ��xsEFR���@�h�<�ul�:}34`���@t�-ȑłe�<�Ua��l�<�#e�L���ۤHM�<��ê �Vq�n�i���#�d�<ɀ�Et���� &ԎMv4}0�fW�<!ScڴU[4,�E�]�>}+���U�<��Hƪ5���ѓ&�J~��S+�W�<�N� t$Ȱ'�C\�v0k� M�<q���̼��$Ã7ܦ�z`�E�<��u$l,酫� pV���FD�<IK�>]��¡?`�,ᰂ�G}�<aF��+je
dP��F�Gߐ��v��r�<�u�M!qeaA ��p)���w�<Q��P;?�Xk��=s����t�<���2>�$�Э_�o�
�G�<�0�ˇEI�`x���91���M[]�<�b�ݧv��BF�l˪@����W�<	�Ȃz^ L��O��Cp['�UT�<�T�-W�9˳�E&i�x�bB�T�<�'hW�Pn)� /�� ��L�<91$��S�h�O�2kf9�D�D�<qf.[	M]�}J�T�\�����{�<QW��8P��G�F0Q!�r���l�<�`���I�|!��$`;�ϒp�<�#�%<$�$�D?c؊��#�n�<1��5C��hQ��$D��`�k�<i&h[�G�E�`@G�i`�����<I�\GƘ������|%���AE�<��DV�J����/�6��A]J�<Q5cP*J���i
(t[$���+L}�<�lL�VoX�Bg(��!;ZXSfHo�<Iu胀t���RG�&G�xaR7n�l�<����mvv��b'� 
���E�Kf�<� B�[0�7f"��EK�y����"OД����<���J���l-�'"O(@R�bG �X#P	P%8�Xi��"O4�`��\�><h�Q����(5*�"O�A��/G"tl���F��� +"OR�fG67,�!g׬o��#u"O�LX҃Q�ɶ)p%���Qo>�HQ"O^M;�������U� j�"O<�3ħ�TS�$
s��9�.i�7"O	���K�@d��AFW�Bw^���"O�Cf
�'�z�"e˫G_�PIA"O҅d㕖(5&t��	��U(�"O"�X^h�%��U@�DgɦY�!���)h�z3!o�K'����$�0!�d�$q%Kہ�\Ě0!����$��'vNA����0p�ˎ�4vy��'Ċ����:�)5��=�(��'L<"5�ZQ����dCX�r�
�'��͠A��S�ty4c�q󨡲	�'���t�L�n)��` 
%uoRC	�'kp��R	�"Z�$
�"R<?ǘ��	�'
�KUdL�+�a���P)C�(*�'�b�-uC��0�L�\=�8Ek�f�<i@�Y��<��-^�;��h�N�J�<���rJ�Ƅ+X�t(\H|�ȓ,�r�D��/�f�a�Hm���ȓ�8� @Hə,>����0F$��ȓEbqh2�	x=p���^*T�清���!���$j�}(R�J-kT}��ϸqQPN׮h����%0j�i��s_�� $�ҿA yWo[)
�ȓ�Jq����p� ���`�/a����ȓH�Py�rE]�}�-��L�<��-��E!� ǆO6�N|�f
U����ȓ!�,���`S�l!nq�be����ȓd�@8�'�T�,��S1$�uk�l�ȓaL��A��z�x��Ο�x2쀅�.rʭ 5KX)��i��k�̈́��V�uR&�  ԅ]H��%cn�<�FKj�HɈ�#[�?y$M+�D�j�<Q��.Lc���`�o�8k�jTh�<i �˿
��`�a�JBDŒ�L
L�<�!��8�ޥ�Tb��>�4���Jp�<��E�&.��y4�L?��MA���v�<�"��L=�{7F�,˴ḥ$�]�<���9l仅� a|N]��ao�<!f� A��˵K�8?N�3��a�<�UE��$i*�@��fX�6��t�<)!�O�<��L����*�t���Ey�<���#nh��J��� QSy�<y7oY�L��x`�j�F�X��Y�<���ϏXH�!�B 'aF&�Kn�<I��(�V9Scg�5|"���t�<q�������"-	0v�YY��k�<aſ`^z���LL�~��5)VTj�<�e&3X�ƹ���ɽAs�=#&�]~�<9�АԜ	���"CᲔh���q�<��+V�Nk>��C*�wBt�l�<�Ы|߶�����`�:Gd�3"O�ta$ �@�	�F�DP�=y�"Ox�3F�Q�T늱��B�B�U ��',z�����GUHl�C��hN�г�
�\�h�6h�0����G_<Qb$AD�l�n��f��vyt�ȓR��ʤ�M+O�6� PB��n���S�? � !���:]�Mᇁ��訂�"O��⥟q�^��!��F0ӳ�#D�ǭ�&:��I��|����a"D��yh�$=�L�s�(mxr3`�/D�Hc��]�j�X�`b�	;0!J�c��-D����.��.K����Eڼ���)7,/D��8�,É7�P����Ysz�]��/D��SS�+e~^��7�ז��,D�,P@g��0��`H�3ȴ�S�l%D�RVGJ�-�V��f�G,����#D��Q�H�I��1�$Mga�#�,,��B�ɍpת��t��1�pL�G̰k�"C�� 9V~�:��	Z�h�1�`	K^�B䉾�����JV�A�r�I�nB�B�	�@�B�p��L� `%&�:1��C�I�+�� �*��$pFW6>��C�ɵD��;�閯=��B0�ʴH��C䉂'�+&��?NTH�2��. �XB�	E9���u�ն9�.������m8NB�)m�*���J�`��1�2OQ'F�`B�I �@h("y ��H���C�	��N�8`[;�����_�1�B䉃?�&l���^�7L攋%�A ��B�ɞ.��)��i�4!e����i���C��3/ܺh1'흦6�����W@�B�	�*���Q%j�vU���&+�sU`C�I�C&P �'hJ�>iH��@ [r�*C��i�LD�2�ǈT@�8��-��Y'BB�'rN8`@ehSE��4�f&�	B�B�	+}��%���� ����V��Lj�C�66d�EU�XKծp�	��ۮC�	�4���	�7H����S[fB�Ir�νB�Ï��h�B�˄�C���Py�r�7E|��
�C�.H�C�	����{e#ݡ}]��+��

 w�C�I�>ez$%�������ҝVM�B�I�P�H�Kₘ�,��I�P�R&FK�B�ID��,ѱ%]9?ծ���M_"T�B�	�SK��3$�6q<J4��-���FC��5z����BԲJ*<��(#t�2C�I�t�r&��f�H(��Og].C�I�e|�x��f՞(�p)��LB�	%v����
��%���"���
;<B�	�v��� ��J�h�
��	>���$A�	ޢ!�c��6w�C�+q!�DF�ujĠ� ök
�M����*?K!�N�8��U����)bo�h��JZ�6B!�d�7�L��E�b]��AD�O�g!��@���b�{ʑ�dC2!��\�'<$5�o��<��I6Ɏ�*�!�H�;d&���._���hE5/�!�DG�M \h�)�6?��إH	O�!�d�j�* k��_\o\%���£y�!򄛝(����7ȡ(Ir�i�/	ݱOZ�@�OJ'N6" ۀ�� �"$�|:b��H[�d� ���$}@�bb�L�<K�?R���R�Hܘ.�*EAg��q��"��?e�D�耫ZĦ�ӈ�Y��G
3}��R�!��>ΔJ#�!D�@�#��.������ 2��t��V��5?!��:b`fT����X��#���X�� �4w~��$�X`p�$��?B�����̃[��`�0�0qf�+���H�N<���O�(
U�E�!#XP� �ŵn����>is�ӯz�a�,\6�aC�)ӡ��
�-��{���W/!!��<�H�;���b���Y���9��B���3a��+��Ë5�&c5�g}bOT�K�~,s7mEt6Q��뒢�y
� Xy��w�����\�!dmX��i�����*Ѱ5�؝j1�D�-k�����A?m����@�:��c ��a{�S76�`CTdY�����ڐ5x"'���j�|sР(8.C�	�1^�9��O�s~^�dD�/fVb�(�䃉5�Fx����N�x��dJ_^������/	.��PIظ�y�ŗf6���,/QrP�3eO�$�|h�e[l�r�'(�M�F�>�GJ�2n�ِ�̑	K�h�c @O�<����-Y>�r`��d��LK'�R�As�!÷N,���Z�I��UK�S���0�`�0S�R��˕�zi��I�v�rx���X?m��u��`7V�0�E�O�F�}�&¯CL�qb�'񒭐�рY����V�6y4��}B�EmwB�J�FdC晳d2�Ӿk6Y�
85��9�ƀ�� C䉀$5d�	w�C-'{�U��̓`5n	IPG��P7��s�W%xN6��}������!֠�1����:̨D%O�!� �Q�(��o�;t�!F�M��6�3��Lz�
����H��*O8 ����8
�p�`�N��f<�3�'�Xɹ�Ƭ�pfOG�I�>�Q �B6�p�Bu�7�(T��+���w*#+�ҵ`u�	"��(��-����`q��ω,JՆݩ��O�Ji�"�K�<M���e�dB!��'/�9yv T��T<K�n������j��'�B�dDգt���qc�	��(��	�,\�hr/�&4��JXU��B�I�G�\AV 4�f�
�gF0٪�:u��5$�R@eg�а=���}g��(b���#�J	�FbLQ������1!%x!5��/p��e�0JJ~d�TC��w���Š8D����J�Ga�����ߧ
x �'�$��χJ�!�#�ԊY+�y�=§-Z�e��n�,��3�L��l������M�"=�>82#E�Rx��V�=�˖�,����'P�����
C?-���*��с^w�$( �/D�(��b��"�����L1�i��j���F@皉��'�<� C-ٱH��E���)��Q�g�I�Gm��!f�C e�?�T�X�`�'L�$�B�[g�<�@�ێE�a���Z�>���U�Zx��9�Q	ÉV�]�H�B�	�?Jͫg���8ax� ��'2!�$ׅY�T����/.�X������L�r\�Q�]y����f��<��>�� �>.EhD @CE�
X�A�<�DC�{�>�c��SmRtK��٦iJrg�6��pHǩ]�.	����I���l`7���t(
�Ý3pI�����]
��r�L�h�N	�7/K�4٤�ζ�Bwn�
s�C�	*"���i�o�s�2�q���gQb����I4(��f�͞%�Τ�}��R,bb�k�]�\��ɛ��Bs�<�e�g!�PPς� ��;dD�2q��px*�)Eu,���i�7�s���Qn����뢁S"�#D�|����k	|�8�B�dJ��ч�v%�/PG�P���\��� �g�'�e*�I��,#���p,Êw�2��Uod�n��E,tz� Ý'��P�Ba/F�x�(��R�g�2�{�D8T��C��2o�]@��
#���Fz�/\�Nģ�A��wR.!A�~��i�( *@$���o႐a@Ch�<q���^��D� ��xE*������Æ�h^�Ck��W/H����i�H�ĥ{@�i �-�aA�YH�'��`��"�$��Q�5%�!��"�L ��	���������B=�U�E���&��V�A.96����Qy���"�N��x�`�ş{� 8fCσb�%��c�'˰?A�.�q����KAG��aa�x�'��&�ă6�z��'��4��4o�z��q �,��`�₸�y�L�[��}[B+]������Ѩ�yr�ϗe4�Y�g�o�)�'O�V�ؔK�����p�)�j��ȓAv�tɱ�T�d
�2�Ӊf�x�O%�am��SM��Ó<&- M�B".t(�� I�n����R�&,���V�DZa�L�Z0�����.[�!�H/$��}C-��~~�i{\?�ax��K8*��O�]�lгn=�-X�by�Q�0"O�#� N��� �Ѧ\e�xږ"Oؐ�DH�&^��d�*!F�Tp�"OD� ����1� )P�X�"O� ��؂�[=<8����T�r�ܸ�"O8-��f@��I���77�Ne�E"O�0
v�- ����!}�Z8
"OJ+d�'�v#"�8�H$Z�"O��굀3f�
���F¸;����"O�p�P"�1��%�#EL�����"OPU�ȼ
q���S$߯A��]�"O|��q�&Q��d�j�^�"O�IBA+ؼcત����eI�6"O�Qs�S�k�B�����)jG���F"O���C�1	�vABF�$P�@�"O2$�GÙ�M��Q�އU�)	�"O�9K	U=,�p	�ĩd��٢�"O4�8�$�T���Ȟ��(��"O*L��bܪ>-҈Ze퀵��9�"O��(�� z�)a�Cų-&�	s�"O�%����h}8���X�Rm�B"O���г6!ƕ�E��6G0}s&"OPPS�h�}z4w*׆[�l$�""O���D�@�{�X8�F�O��:P"Oʬ�DR1�z�a'�&LD�K�"O"��s���mn���lZ�=�ޘ�"OzђWj���ӣ΋̛�&7D�h��-���n�S Ȁ�m��ܹq�!D��a�,��e<�q�e�tي�2D���Bm�	%����IIHf�!�c0D�S��ոikX��!���		L�Zc�>D�d���K�6q���]� �m�C�8D�\3��ՙQ�x����>7wD2o&D�d��+(>L�����,���D$D�h���0�RP��V�OЉ��A D�\+���'���"m|��1��,D�$���$9������y~!�b,*D�+Q��hQ��'��:��� �=D�`x�ɟ,��`d+��t��	�U�=D���$e��wzv����wĒ)HU�(D��S�A��uT��b�D3w[|�Z�J(D�X�S��dT]K%��}��h� D��IVbR38eZA��$Ĺ5�����%$D��;��S�,n�0����C��@CTM<D�4b�ǔ�+��H��NÌt��0��m:D�x�QՄ7���p4�C�.9��ɒ�9D��h��Tn�B��"jT��cK*D���g"�H-��#��d=X��`�3D��0�P:�lJ�O��9���1D�� ďƝ�D�V��/d!Yw-D��C�W���[�U��ūA�6D��2�ZX����A�;��Y�7g D���e��$%����げ&�MY �/D��QG�D8�: ���^�)��.D��1ܺ]��a�Iݞ'�2T�e�/D�����<?��l���[�F�֐0�-D�X(2ʓ�	�څ�R/и��-D�hbcA.V=���k֖;��|�g�>D�x���`�$�B$��h?D��"cL�	���"ꓦ`���ԭ!D��IB��rz����#o�6trh D�\b��F�]lг �Y�&L�@�J4D�d��F�?�9Ǆ�=M�y0/4D�������SM[.d
�l���0D��X���)Fb�R�/�-yb�|Jv�=D�8�s�;�8%zA)�(a`��c�&D��`�(BrR���^�w�6�9�l'D�HȷOI�vz��  ��k��a&%D�� �Y���B`h�b׆5�$H���'� ��e()��!Qd�[8 �i�rhˑ]1��1�O%�Y��R��@0잃I�ԹQ̍	=D�!�ȓ*BH�'�~ ��IR�hdu��mv���g���R�h����ȓ=��:W�Q0�����,�5���"����m��1;B���X!�p�ȓ.�\�����c�a�(�/oɺՆȓ|��H�E�K|z$�S�I�ZQh���l"~��S�']�
2��u�.1��� ��2�
Cc$�b%&��J�"u�ȓoƨ���(�]HB�J�
^��V5��4�@ŀ��$Z���RC����=�ȓX�X%��A@ gE\lZ�[�
X�ՅȓV:Q�֥U(1���3s�A'r	
0�ȓ��1�l�aDm�b# "�d��\�}PG�;yE�С!���]����ȓ9��"��ۨ"��q�˽�KZ�<��Gb~jYXbi�,	���n�<91�Ԏ5?�L;sa��-2�У���S�<9��>6��5�m	<�H�v�R�<i��@쾨��������K�<�T�P7)��c�b٣L!��p� �O�<!�����a���i�!%��I�<Y�揎!du��S��=d��H�<iSF��2������,~
RcJ^L�<iС٢M�<0" �\�r3p�A1NXG�<Q��L�Ux�Ĩp
o�����A�<��!�/�]�B��<�$����|�<y�"6�� �@4},���iDN�<�m<:3�U��%�#|0�1��Ar�<�d��6Y��u���!N(0��e�b�<�"��2�P�3�ዑ2o�\p�lL]�<a
�D���ٗ�� |��v��o�<�6�NLA�(j���7��Pn�<!�5F��Y������)q���@�<!����j�h#dM��U�|��t��T�<)��
��;�@DG:���i�Q�<i�� �Kb��X�+sh�H�<�5n�5m�v�5��g8<P)�o�@�<�S�-{(����,6�и1��y�<y�iL>m��l0��'z�m�W��Z�<��+�G<��1,�#y8	��'MS�<a���x���bfk�$�yp�nCY�<Q�e�?E苓(]��ΑӢbY�<�@��!8�N�Q�h��L��pS��T�<��i��~efp�'�����R)P�<iT�U�y�,���C�w� �Z�M�<�E���-{fd�
�V��dFPN�<ɅMT�X�4t�L�l �1ɰ��q�<�֬S�*�YQ��C�iߢd��	b�<�懀(>��t��MS}�b��G�a�<yQB� T��)�.�J�rl��ƅd�<�1����Z1�dΔEf 
4�U�<I� [Vk"�[��C� ��iA/�{�<i�MW`���1�Ş g(��o�< 
��Wy�h�7"r��@�j�d�<1�%\5,�����K�R��ӫU�<qA�	w[p��U��!6:Q[Ӧ�N�<Y'd�s7��+��!�Te��s�<�b��a�$��-���!�d�<�BT{�%ã+�Z_��W,U{�<	UÌ�b��T��:O���D�Qt�<�J�2�e��Es��21�y�<� �3	Q"u�bȓG^�(�Ò"O�eçH�	t0R��/}<��a"O��c`@�7��Q �-)1����"Oҝ��OԂF/�� `�a�d0K�"O�@֯�qΎ�x6��n��3"OJ ��_�l��ٴ�ސ'�8-Aq"O����o�!� ��a�%Z�`8#"ON���O��l�>�)o��p2B"O
�Ӧ"�_�8LÓK(-$���"OQ�HO'`�X�C��F�A�R"O:X��Ͼ �0� ��{$��b"OFI�1d[%E��P�0��/m �(�0"O��`�L8�n���QN�,���"OZh�-I%����l�v���`�"O���˃�>�t@��U�M�����"Oɰ@�[��f\r3�֘i�8���"O\�SP؅A����z��(z�"O�����?_z��F�U���J�"O�0�уHL�])P��6#��-�"O(%R�Ayb~X�COʁ}m�	�v"O�!qe$�3e9���-+69��"OV��P+�>y1DP��o$� �"O�7aOuͻ��;+F�55@+D�tɃQ<Dm 3��c���)D�������i����4� @A�K(D��`�Dí<g8-�ħ�HL��� �1D�� $iݱ�l�q��#ڊ��.D��� !ՊP�vǔ�)L��+D������Zׄ���&G/:�0�<D��q��Z+4$XA�F�E�`�;D���#
�r���t'��er%+��;D��p���9R�f��(/8�B�fA��yr#B�Y��x�� �����N0�y���KvR� �&ӽ���q�FJ��y2,�h�����NU�F�5�K��y��Q2C�@� �2TG���,S�yR�Bx�搹1,PS��]��A��y��b��}�UFQ.ز+� �y�Bǀ,������Q��a�λ�y��	�*��,�a�QMRY;���y���W�"}�E̗�K'�p��y��E�zVh[��P�7�dABn��y�*�yF���JY��䠊"�y�)�O������0P�1��G��y���44�:�i�ODhrfM�=�yb�� a�!��HR���'˃�y"��3�"e�>(��1i$��y2"�+7=���Q��Q�Rг����y��[DHI$��#CD3E�9�y�
�0x0��߀t�0�@���y��ڕ~	�yme��f�xb���y�Sl+z�	��
�*�6�Ҡ�C�y��A4YDq�a����뇈?�y��79��݂`�P�����G��
��'��{AF��8l�� !���� R�ym�D�I:s�Ȟb�Z�b�����y��P�>��	�a�
(ڸ|R�E�0�y2�Ҷ�xm;��K� w�ܻ��A-�y2C4V�j�)	�" ��*4�yҊ.2�h0�hU/ FhdA��y��V

"�܃�ƍ�zd����%�y�
�N�+�"|����M36C䉀%=X��6!e������78u�B�I�w,d�IF�S�Vv�!��D�B�)� R�iЯT�kTL
�FVۺ`�"OPh!�F�F*���ʨA��{�"O��W�2)��X�$A��zY�#"Op;Ƌ��j3�Hqd��]X|p�"O6lbt��*`�*|�3C���.��9��uص��#ެ�&`���@2s�ņȓa�����A\)v�xhP+_Ĩ��vǾ�K�!M1w%��z��Q�/RD�ȓa"l[��bOx����@)^ �ȓ`X � M��xS��v�S�]�Z��ȓE��x"Lu�Г���<���ȓc�uk�B�C�l;��ɗ"4 8��1���x g�O��Ф������ȓX�d�\�cinEh�������	�"hذ�޺?%6i8�Ğ�sO�̅ȓ.�:���,Zc�u/FؐQ�ȓGc|93d�Q�~�r�ʅ�̣�R��ȓa�\��I�]r�pڡJ�8=��H�ȓ:�r
�e��]k������u_Nx�ȓv�*��E~ZU ��3$����ȓ%�LI�N���R5M��Ȱ�ȓ<t�KE�ͺeD�R�'�<+��ȓrd�AɈ�T]�-7��l�2A��¼��� �r3��; LA
-ΐ��ȓ;eD��C�'�>Xk�քn y�ȓGc&M��O\#+�����dyL���{䠡5C��Z��E�I�L�����>�p� ف I��8�.Ǹ�:p��*�\�k�$��hÀyx�"U4 �4���8�R]���ӣ+�$��҈F/j'4��ȓ]
�H�L�=���	-nL1��p��!ʒ�ǔ^���c��@V��w��٣Ȟ�1=v���%9-"�B��< n�⇊S |`8�����&B䉊
~8�f*��>�P�+���C��C��	E�9DA�o�hp-�"T�C�	=H8���ףs�e[�ᓙJ��B�	����"2�W�g��00융>�C�IL���ȡ��3���b7%�2�C�I|vp��F�*xbs6�DC�I�Ҏ|�TD4u�D+���'S�C�	QZ8$3�D�S��r�L��Q��B�	qR�tkqQ�JI��B@j�] \B�IlJ$�9�M@#��0U�^�XB�I8z�"X�T� %>�������:��B��,�b$� Þ�;JL`Qf��9-�C�	���R�N#��)aA�ȋp�C�	�)�=*sBS!K��h��⅄w�,B�Ix�pE��J͟tjd�2���H�B�I�N�@5���ك-_>L^S|�C�	
�02f� T�$4����>�B�Al��{�K!<���Y
[&-B�I�)󂅐䢑2q�]8v�T�D�"C�Ɏ��qiAa�\0X��S,+G�B�I6@*u�1�2p@b��G%�B�It���!��#U���(��E�o�B䉘?�XS�c̕gǨm!@�vI�B�Ɂ����T�2�Eqe���|�B�ɕE����w�ʰ5�L��mZ�\GjB�6OoP8�ZT�xDa��ה%��B�5	z8�z@���-�.��5��p�B�I"~bj��u�)Nl��T'��*��C�Iy�6��ҧ}|� iP�;.�C�I3d ��!K��zĊ���~��B�)� p�������C�)@/(���"O:�#��6
	�d�D�~ªI�"O~)�a�\Yr��Z��#jZ�p�"OR����L�OS��{�>j��aa�"O��a� ��� �nR���q"OМR�(�K�u���.7�L�@s"O\)���Z��e #�7 ��X�"O�Dy�E&q�aIq��Y�v(�V"O��!�k$��!8a$�:}�}��"OM��oE�Y�I�A�,�`�LR�<9��7x�e���� 7\�����(D�l���Δ7�h�U�X��X��&D����eʂe�6��V	��5	Nl�Ѣ&D���/D���p��Z�~��Ǆ:D�L��B�/�|mȥe��;�����:D�Dy5K˩\\,N�EDl܉w:D���1�/���c��Fh6����<D�4X� �r|����"M�T�"$:D���򬏥oV���W%Go�9��9D����L/rfԴ�eڝ���6D�T��B��
���3kķ(����$�(D�\�B69��@�kC�]b���9D��AsDˢf-���ԸB+xU�ǭ7D����Ȟ#BA��{"� �g�4D����NC�)g�)��Ä=����2D���e� �iX����-�5+��,D�`a��%I���z@�� q�*D�X:�O��Ig ��2K=4�0�" L=D�$5'�_����"r#�xX�Gz�<a�$ҹu+B���*_Q�`h�CZt�<�J ̘����(��$Q�Iq�<�b#��HѾx�MA�nu�TԈ�w�<0��,;�X1JH)Z���n�<�eAK�1�h&��dN�0r��]^�<�GJ-u���R@�"�j��)�\�<��		U�*%���Fnʩ�P��V�<�TǞ1:N-��M�Lw���S�<�t�� J������\��qP�c�f�<y�i@�j|�ˇʕ
cngTn���'x`�#���g��	q��Q^��'��Y�%k~(%RP�S���H��'#ʴɥ<A��l��  #�y��'����,�=^nP�i��֋�f�q�'�鰧�/��)B�:r����'�R������Ab��5^��q��'adR��#��
B��(I�e��'��1�b�!���bւ;�z�x�'_Ju��oo�\"'� �K�e��'��i"R�������A�,��'R��h1` �=�a዁5�x �'>��f��7���b�P�ĬR�'#8�[#�
<0�pȆ�3۰1�
�'�m*t�Y���b׃�*���1
�'B��҃ 䠩�Lˬx�(Y��'�����Ȃ������ڋv*���'�p�!�^>{�(E[��=���'�6pZ5m�#�$��.ݻ.�b��
�'Ƃ則)�>�*)�V��8�L��	�'�؅��\G��F-��.64	�' ��6��-�8���.x�6iS�'l�sp�OA��X5�G�r����'qF��gA�;ZT��a�h�(�'�hp#&ߢ������6�LtK�'9���1�{��p/�T�PKe"O� ��S��/�8r���!l���J�"O(I�%�<W)ʴ��b�$@ %"O���`��R?�-��*�N��a�6"O��@��͔Ij4���
�)s*j���"O�%Ȣkܫ  �>eF"O~�!B�Z�8����  �m""O�4R ė1@�x��+��>��}8G"Oܨ� K*M�ʕ�@jG�P`�#7"O�Pe쉿���
���wp�A��"O�XjuF^��B��ݾh�Թ�d"O�5��:	5~�����4���K�"On$ᓇ�E`���\.G���`"OD1)�-/�<�Q�S�!��yg"OZ�;�(��l�b�)�bؓ0z��"O�e`4�@����bֹo����"O��H��0!���↍_lց�0"OqPn�8HI:���KX_�!P��'�����(XX-�� DC�d=�Ħ@*L�!�D���c�$� D�d�C5]q���E��*@�@���j%9�!jB�yb#L�x�P;�CX9m�!QҪL���d�Q��(��Wk6@�Ѓ�._� /���"O����	@�!jӆ��W!a�&�x2��W�� �t�0i��|���K0 ��"D��J⠜q�ui��^ _�:ծ,D���b'͠smT��G㜭O�(!��,����xh�)ϘT�D��um��cz��4"O�D� �G��ك�%Z�{u�tJ�"OV!P�_� �=��N��^���"OxѪ�����h[�V����"O�$��䑣F�:��ܲ/�� �"O�#C#�nɈB�ݲ(��0�"O�� C�.f�v�s�eۙ)+���"O�Ă����ဲ'�8V!�}�"O����$Щ�t�����"O��#�G�}�� �k>s��0i�"OR}����:���d�[�ch��[�"O�ys+��vyk�>.^�ks"O����ʑ:@�Zu�G��<V0�1�"OH=�ᢒ�h3���H,;x��W"O�!�Wǀ`�����5�*��y�EU�u�2Az��.u��Ju₡�y UQ�:�Q/O�t���p���y�%H�aF�%
R+7.~���`J�y�ɉA�AW X�/��3+׿�y�t%@��g��'��1�C��y"l��^�á��rd�A�ʵ�y�g%r@�h��Ў+�(e��-���y�X�?>-�)My���b@��y�l��X��h�W�Ǝn�~���3�y�% &B���#�Ȏh��]�ƫ�4�y��6�4��J�j� �!��?1�3O����F1^zlѲ�?u���q"Oh2f眯WdL賔 H>3Z�W�ɽL"?�rc��,kT��j�H�|8"(rvj)D��$�8ALd��r�פ�2�l�J�d���ا��h�i��ðr],��ck_�D����"O~�PAݼWİG�H5bP��b�����ɳF����Μv�	c%ϛ�b� ���u��!7&��f�#�`Y-I��a�QH;�yB�P	��(�gAy��e�a�Š��O�"~"�j�t�UkO5?b=;M�X�<y�.3��f!�:.�m��JV�<4��m{H%gh�?g�t��*�R�<� �p��GZ��|�!#��7 *��F"O�}{��N;qRlp@$g�h|��ya"O*�8#��x;�e�!g��G"O�����
%���aF�ֺxOڡ��"Ob���,M1�؄zW�˲T�|�"OV+$�>,��պ6NG<A�Ly�"O�%�������2��+�"O�9�� p~�����U�L�s"O�ő�5X�a���y�U"O6��vcO�u�0 QFAǒ_�Ј�v"O���.��JS���Aٜy��]�"O~�B��ͺpx�:��Y�{ru�u"OR�*��X9R��0!CE�{�Ƶ93"O����CR0`A���4��u"O��xD�9�ؠE��+�&�9�"OLeK�GX�;Ԛ��'�"H����"Od���#ŧp��ak�C]	�4�"O���M�=#���d�L!"O�1!6g��O�l�diU�#ZT"O�  ��3V���Ĉ�%J"%"Of���nݺ	l�t�f�_v���"O�!i���.%��PE#�yp5Y1"O¡�R�Y8�NXeM	gj���!"O�Hi�@A�`$�$F�[f�t"OFH��*>B�����|�M��"O&��(�e)�A�3��jޅ�5"O��b)\k��L�;(��"O���&'O��,a��f���*F"Oxᨕf��ZX"4o�)gbp�z�"O8��R�X�f�~!zO͛+��E��"O��%S(-g|dh��� =� U�Q"O|- ���
�Ll��ִ�@$��"Oh��Ĩ�!�l�Q�D�]}�98c"OzY��W 7R��Ud��m����"OR��r˒4R�DD�B�&�p"O��S���0!�g��(�p���"Oz=�6oƎ �@��~?N-q�"OJ�S�� �Z�C+K>i2��"O�U�r|d���j��x �!�"OZH#��.Q>r珈n#d�"�"O���ud�H|@��iP9o6���'t��CQ�x��=zT/E�	�ʝ��'�Ψi䃞9#�th�I	�~>pE��'��T�&�^'Qer�CTDޅF=���'U&8AU�
2���L��=��E��'C��P�$�X1���;�L��'�^���+�#'������5]`1)�'��V^�H�� E=4�f5p��/D��kC)]2ͼa���n����/D�̓rj[8s���3pN,����	)D����-�u7����D�pώa ��"D��9V�=�����Ǻ��p'�+D�@RF���4�B$��Y3T�ڷ6D���'K�f&D���ⅺE�&�;��4D�����g���� HX/Q�\`� 4D��`$ݛ_H��4�B�^&��c�=D�4����=3]>�����T�(�H=D��2�nΓ�`�h"��?��{F�;D�pB2�B�:���؇c =]��PE
<D��T�2GD��
L�I��E���5D��sV��=QZ|AO
1�>e!'c5D��R���I<r35��0D��hr �?�:�	���`��@�e�0D���j�P�HK���1iG�x1��8D�� (����B�k5$�Q�/F�t�@�@"O���U��36Ūl��Y4:��lz�"O�����ِmڰ�S��-<��jW"Ot�1Gl؀,���0a�\X���"O�%���/R70xqҍT=�`��""OH���'g>�d�.���"O�m2�"L�%>�Ш�M�(��8Z�"O��3'D��&ƿT��Z'"OFx��I)wf���љ#�ƝI��'����'^#�q��'F#,5ȱ?&�p��_#Orh�$�O����O4L��O����O
��$oN�[_谋A�̡T|�$▪	�NH�P��[�ʬKU�{x�d�"���lފ<b��{�(Y��!��h�	ΗT^��� C�b!��ѬZ�'k�h���X?�0@5k�,��=��-�rgv��M{�'�2�'��O�S�6�09*qG	�M���G�=�➘�L>?��I։v� ����L���mN�p�j�	�M��i5�	d@VXPܴ�?q����J�g�.x��L a�X�Yb�VJ����K�ğ4�Iǟ��f-D:�t�����p�IL��K\)F���k���9��<��D6�HO4Y����8|�\렡Ɣ{0ޡrc�ֲj�J��'�[�" ]�6��:"�mR���@�`��{��R��?�i�6���l7�ɮ3����:o[�HBBȟ�%r�2e���?����OS��\/�1A1'Q
S�\�	�NB��$���as�4�M��ߗ;i��*�g	��U�jŻn��7͆ �d�n����'a���O��'� ��		�X¬Qa.�)p��B7-�%�tP�T�F�,|���F0t����Go���?����f	>� %�7q�ՀN��\���ylĳb���.�q�v-N�Q���9�Ư���5�ņ"W��<b1�Z��ѹ�
�MC��}�7MNΦ��޴�?���i��z4*ϓ�\E��Td���*�'BR�'�B]�8�If�'W�.��i�4%�I�1^U��Dy�
�OJ71���42��ם���u�F`[�]{29�c���C4�����?2�M�B Fl���?���?	��4��p�����k� M�����&? �8b5�Nܟ覈�5KQ���דd�Dx�F�<ṷ�sʆ�ker���@J:-R3F��^!!N���߂��x1�d�uy��I9�q���(�e�u�W�
_���ΐW�4��䦙�TQ?��?i���M�M�7b��Qn�PjnaґN�9-�!�Ĝ�p��p1G�-kMR#�9z�i��4,0�&�|��O]�TS�h����tӜ�s�e���1�^͢	�b���T��֟4���/q���	����	�<�J8�!��(q;Tx��.oY�D2����J ����������'֞l�'��U��!lZ�u*X!p��D-y4�:��ʇ@��58�[[8������O�}�G$�h0a�Vd�	Z�R��D��%���Iԟ�?�O xi�K�.{r�����9y� \1�{Ґ|B��%'N���L�"��H�n\�A
�ɹ�M�B�i��e1`��ٴ�?������\,a� S��$���O����n�џ��	ڟ,z���h�ܜ(B�O��D�~z�8T\��#c 6��Ճ�Ɔy�'t�r2�3>.�C۞c�2ACRD��'C�A[%�)C��jW�2
"u�Vܨo���=�&n���ڴ5c�O�֭˩K<���% (
k6��s��g�,��(��O?�D�5M��ؓ��p���)F�#X�|�GgӜ�nZ����e�j�tk�o�0�X��0�!}2�'a��|��
J' x  �(   �  �  �  �&  v-  �3  <:  �@  AB   Ĵ���	����Zv)�� ����'��Ot\8���6^���qc͕<Cz6�ON[ƽJ7陓!|��2adޙ"$ݪc���)!��.C�Çn#D����Z*+��|�"C�>k�~�k�ˁ=M��BΎ#!`�Vk���4�sT":Ȅ�S��4�.H+PɆ3Q��I
�fz!��!G�K���Rẽ�^�A��|sDx�X.\�~pk���
62����BV���΄�B(�щ2��B2L����7-��2b�D��ĩ����H]���PEJ�%���'Y��'1���Ꟑ �Xw � ��ᄋ'�KH0��y ��+)\]��$ɓvb�|��G�ź���`e�`j�f��F�<����pI��+Q֨��F�}��A����0��"á|��:sX�����>�3KƉ|�`��.7���Awy�J�?��i��#=��'"��C"�u��呀�H*#�-َ}��'����!�YR�5�(�<9P*t�޴HL�	t��O�)�(�F%A��TAʰ�G'�����#�������?���?Լ����O��Sw��5CVĜ�5�vd��E-s�&��&�L
u��8Z"�I=n��@;�O����O�B��Q	A!&�7f�=:��� �CP��Ҽ�%� bdhl���VDW��mZ�C���AR��Q�A�����t�0@�a�R�m"4i#�$�-p8Ɖ��*��E:2��[�h�4k4��y���}�'�X��nG�`[ �`W
�^��H(�O��l�K��<�ٴ�?1�����%��l�t�C��\X�7B["�M��OY��?i��?��/F�e�^���Ή��IfB��٤/r\1glS�(W �K�!�l�'�
�N��+wH��� �	�(���N���#b��3�ў$;@&�O��o�ŘOǬ�R�萷!znt�h�8k�v��'�.�?����?������z�^MpAl�4!�����1�D6��<I>�|��R�|zu"�/"�00N��_I�`�H΅��dWZ`�nZ�������4��&�1��ğx#�+��d���(�N�4����b�г�M���Z�"�Q�W�X�2�{WnZ��i:�S�{r:5J���dͻIH�v[�E��3s����L�_�`XA�#�4L�#~j4�ޮ;�,y�`Eʝj4���A���?��ʒ�|�޴B2�)�����(�C���]�\��k»��C䉈]��C�O��,���n�7	�c����=�HO�7�����4���At!ܪXZ0�n�����S�Ɣ���Jş �	ퟜ�I>�u��'���c�HP]����^�*�@��)@��xkw��6����'"!>��!�O��V�S��ēpЭ9`�RI7�}���� X��z��:�쩉g��;�X�ӆ�i�d ^�[�26��>��I�g�JmW�)�p��a啉&�t�^N�\�����	X���tD��5��Ih��Q�B��K�fX�ːxbf�+�M�K¹F ��0H�,��6O]����'�	�bA dTIM�T�n���E&N�`�c $��!�΀�����	���+[w,r�'�R�ˊ/�ʄSä-�R�&�J$�ČŮF����	�+a,��ď�qc�x�����C{�Hf��+P*�G��>	�<��FK�d=�B��=C�0L��CƾyR�O:@�#�'�T(���Hy�a���r��@��h�L5Dz��d��ԫ���E�0��& ��8(HP�",O�<�"ʕ�hg�jE�H%aq`ܳ� �z}�Br�,�n�hy�MH	�&7��O��?���Y5z���S�jv`��f�d�rq��O���OB���7!G�l�pݺ	���Q� H�|���)�d���G��$8���Ct�'�,�ꇤ.�����Df��)��;�����Ɉ��[@cb���	��	�E/��d�O��>�K
��x٤1y�Mь�ի`�>a���p>�+x,d]�F��] "����qX����O�$�����_�h��G{��E� ^��
2oE�M����?�*�^���O��tZ��|&ZQ����� loZ~�Z�a��09�ڍA�_S0P�+Ȭ%����|�5��<4�nqC�eJ�}h��dA��<y1j.t7���E�!yz�	�&�&�n�
d�G*F	�j/�Ј��n�&��ya�\�!O<q��#�Oxi`b�'��O?�%TM�fd�gD��A)���(\g�<�	B8(nth��@���*�M��?��i>E�D*�tK֫�=/h�Q0����M���?��LV�u8,��?����?	���\��������-�5���~g�ŬCg�b�OGX0�2�OR�fe�Y�OU�ƮY��ē}ĔX�I
Y�U�0#J�K&����C��lkRX���4}|<�%g�B���i�r���c??!��[�N��	O_B��A�O@y�G��?9��?Ɏr۟Z0�!ʘ8#Ø� �`P�52���"OH�բ�k���b3�H�y���i_�#=�'�?�)O�
��W	8N֥0����<���Q`�q/̤�04O2���O��D�ú;��?���(Fiq��`a�'36hxQf��Ip�Fy ��SU U�74n��ϓ^Bnr�ٙ's������l��]��O�W#V�y$�x
�в�n߈|�V��d�UTb��]�n2�/� � �P�[4C�6��~�'�O�	^9<�Q+ͫI��IP��W��Ov���Ox˓�(Ox@��P�[D������$J6�i���`�0�nZ��ٴF>��i"�':Zc!έ!D���h���A�S59�E�شk�����?���@R�,���}o�H�$B<=��C��ɹ�e!X�; I��.NA��P�bd�S�^�<	�mX�I`���LDx�:�R�b��d�^e�� &%�g�rx8U!��D����ߙzhb�,�wf�OڬE���]�R��W(�+U2yB�Ń��y�d�yr)�(��6p$��+B%��>I6������sHҐ�+[�p�QE�>y�
�z����'l^>U�l��|��/ ��)T��: @"�Nx����4m�l�����X���*O�_*�"c>	R�)�MPrQ�P�O��\��-Jϟ0�ǣ�<+`��wf�n�Њ�iAU�&����|��ܛcȎ�_����c)��ӄ0)�QBpK�dsV��P�N��E��r��!aT��.x�x�
�cF�c8.�>��t����S?$��������1QF���'�x�4�?����*�����<A���?���N�N�Ok,Q���'*����$�fX5c�3D��	�2�,Q���ų�H�)�8��'(� VI��nA
��5S�l[�$�[��XL:����s 0��)K����Y�9dE��jy9���zB� hgF�U� ���O��mڇ�HO
�	�Q�P��bۋ&��Đ��_g:fc����:TH���ܖ,��<��ˑg����ܴa��.oӊ�O�I럨�6M��V�x�E(�.F�VL���!ҕ@�d���?a��?)7������O��$C|9r@Oң}�`7�K�T	H9��)���C@3,�AV����O��d	�.�6"�HBt�ЌȍN���d�ƧO�&�����7�T@mھ#��Y�/X�?"���$��)HD}����Z6�h���98SL�l��HO�=��`�����:��a���.�����	~�'%<�A�/ۀbN����]�?���ӯO�AoZ�Ms)O�q6
����������2ux�'Úy.e)��'�h�oZ�A��T���d�I	Qm�q�*G����OH�Ӈ`��QWL�qq�E�S�	���=���)A&��S�l>$����,Zk@�*ĠU=x�X!��w�ҽ���@Y��d�;�-����Zɦ�M|z�
tΈC���3�4��W/��aC�f�'��'��'���'��s�Eؒ��TAjD�䉎ҁ8�I&�O�o���M#sNR"ob�as�#�(a��K��@�S���i�@���ئ!���@�I�?��PA^�|��&7hQ[��ɭRVfDhᩙ�x ���4b����LǄ?K|e��|Ԋ +u��1��"�Ӓ`���R�Dd,a�5CT�@Y�	)g�!G$��Og
�1�^�#l�;eE�)�Ė�t� 	Z�uӠLH�j\�H���)i�҅X��?���������'���H.H�$�3"H<� �a�H�L�!�� c�AI�!�c��:`L=Ց�R��i�r�f�&i��HCI�`.ư#�@�m��,�ɷF�
��]럔��֟<���u�'���:��ۀ?�ht
W�Ct��m�& �cn`�Y@h��IZ��@v�֮Dm�ʧ�O������l�.�Ѓ@�/Lޢ�Z�T��H��5�N�
�컶�P${d�����1���x�]�V�ޜ�PaMG$���F#>�ؕ'� ��?����'���ɼf��R�J���!���IM!�e�i��-A~>IU�V�&��l�<�HO��O�˓q���pD��K�� ���r�1t,ćh����?I��?i��,���O��%!mĉ�F�<[��``V��$���d�[,Z+@����Q� ��-�{�'�ey�Nߺ$	Z�����z$�)j h^;��d���ѥL��H+��?6�џӓ��O�p�W�A;a%�����4&�ɲ�¦A�I^���h��vEM�ggzA���U#���akŋ��<��d��,U B�Ը*�����;54�ɯ�M�����$@
Cqph�OAԟ�6��2���A�<R�e#��i���˗�'B�'��X�/ҡl�3��@h���jU�n>YePZ�z	����D!G�"ړ"��ea׀Ңm"l�F!��64 �ӛOsB�W�Չ E~xań_X�	��� �P���'�q���a�� lb���i̕^�q+'P�P��L8����,9�l�j�<)�r���&>��4��|�c��hPG��?���($EQ��\|�C�>���&'��&�'�[>��H�����	��z4�%��r,A0c��Dc�MY۴�lT�S�)? �!i���b%�[?E�|�B�TQ6<bS�����S?�Jd��w>�c��� N�	H �@"Y�!eͣ;N����jT(3
�z�o���C�rW� ���?Aŗ|��I�W�Μ�c��Z���"qc٬��B�I����#V�������nJ;
"=!�#o����" @�z�$�gb�nwFq{�4�?���|7܁�4
���?!���?I�f���OklA�y�H��
XY.���+��2�ʴ���iNj��Vc_3N�2�S`]>�DxbA�ElP�e��^�|0�hIgx "�GH�B������D�>��-��Ukp*�'3p���'�n���b��Ԫ�o_�`�H��(O��JC�'�2�'��O����[z�ab��)�rt�����)FC�06���6��AU��G�7-y�����'��I�;r�`�p	ހL��p�Dҟ{�4��A9��=��x�Iڟ� �����O�@���1b�ڬ�A
9��3���I�fR��/��p���ix�$[5�״��cOR�>㞵�����j_.�dD&��=�0� #�ZuG"��?�� �࠵�N�SP���e�P1����i�7��Od��?����?���IZ)n"A���<���Q��X���<���dқ2J�ljFB��22`�9�'R�p��ɵmd�1ش��H���i��'"ڟ��2�ԣ 
X��1���czq�װi�n%��'4��'Ꞥ@���.sl�l#`�T'1p�%h��?�cS���8��LS�T4��tbRm!� �
�j���52�:=�V M�0�v�ʓ��b�b�*�� �"���yx�!�B�޴d�a�l,����d�l��o�ߟ��'Z�*d�@�]�-G�3�OӫJ��`oZʟD��ٟ������&Dф+a&`s�������(o�ր&�E{�OK�6��%���[҈U�t�I�;�(Y��*����Ҷ;f݈F��w���J��=I������F2h
Ly�ƬS�\�w)4D�H����=2N�X�$a�0l��hY',2D�8�S��O.M:��B�\�v��A.4D����f[�%�̐��e�'[� ��H7D�h+q �0f����΋0?���0�/D�Db�Ʊ�ج���ʎz���c��;D�$[�k��Ev� �#��(�
L��C;D��F��4�<�A�� 5T q�*%D�x��#�#1����孎Y���*��.D�����)�2eрƐqs��Ƞ!8D��HU���|b����pH�0��0D�*����f(������;!DDɓ=D�L�ND2U��Yf�V�Z���;D�|hFk�FS
5���ӕmb>�Ҵ�4D�tdL f}jm�&1/M�	��%D�l�����
]���S��)=g�)�db!D�����,�V$9s�'��0rUg/D����-Kh �0%�K�d�~��0�.D�����W�A2*�$Pt���b.D���t�K�k�ڼ��n�8y���)�,D��ѕ�؀I��b���yD�AA�B)D�੄R�:��]�G�	F^h)�!"3D��r��D�XNX4
���#^d�*#D����B�#�h�Z`F��VL<26�"D�d0��%t��3F�K�u�Ze�p,"D�,�u�S�	��U�S%I?���h,D����?8�J���n~��	��)D��B��O*�
]
$��f,�e(� 7D��C1!T�fX����g��q+�A4D�QҎ�=	ih��(q���b��2D�(����+;h��"��?T��˂J0D��� �R��lk���Bxy� 1D��*����2_.��6&�	~�����>D��IG+rt@�n�x�s��(D�83 ��!O�E���;N��b�3D�h:��4� H�DO3xf���2�6D���0➌�4�c�d��J�6���3D��6�%y���4�2Le��z��4D��d�K�&��*�l�S��LCB�-D���([�ehx�	���/,���7D��x� W)z�Ȱ�w+E40t�U��4D��@���B�"|�qC�*S����1D��"�!��_1������/~��)X��#D�ĐT�B�=biy��E�R����d�-D��!5��an@�(�������B�I�
�Zܫ�h����'���UIB�+dZ�����m�J�s�����C䉡'��u�k�$,\��+�]�b?HB䉶y����π	�J�b�$+<B�IG������#�\�񁬅�}B䉽+�}B��%`��pC��~�B�	2L�X�W
���*����ðB�	�Dp\S�/K�rL�y�уU�EP�B��d(��G�m��Р��>GT
C�I&z�x��i�cc>$�%gP�x�C�)� v ��L�7G��M;6�[�:�b�"O��h��6s�@b,�r,�y�	�!̖�k1�v���A��-�P��qO\hXI4|��!�X�Y
Бy�'a�hY��N���ЋH���  �jZl��Ć*\������5|O��N���a#�B�L�P���	���Z����*�0AM�����&F�H�	
t��v�>�!r��Z�<�G��;����6۱K d���Xyb��L��,��\�;#j{��&�'Rt�d�mաQy��K�mD�/���ȓB��<
!c��Q��$��S��+f+��0r�i��4j���rN���g�7���rS"�
E���8푔u����I�J��t&�%+��z�NE�C���'Ѕh'�]��н��d8ߓv2bY�2L_|C>�kqML-}r^%DbI� ]}p�2��%�t�x����`�#4I���P`��A�i��4� "O0ԠAn9��-�W�0i���1ST�L3��W�K�$�ӥ�D,u�ڋ��a2R�,��"�"�8�{�"O�P��7T���tH�(_�ɠ�%q�q�BAcӎ����"940��qO\��ֆ(�n���Vh2̨V�'u���nʳzf�i7��1v}ޔ�q_�g&<�e�يV�b��%|O�$؆�ϱM�PyeB=
gbA���	����kB�a����%B���!�B��#榜!Z(�D��g�<�����#��ɋ��N�k���' Ny"+a.=�!O��l�2r� ڧ]����B�jK���ċۏNL\����ag��y��Q�$QP9P�o١;6�Șݴ"a��A� :��g�G��Ey���)[���
�Ê*Wd��Ig�BE0���G������I���p���
c�x&L���D��FM���@x����6��A�D��y�����ӤcȆ12���ơ#�@S�fS~`� �ճ>I����"O`큦Ŏ�Cp�5���mF�X�Q��`�D'HҴ�a�Jx; i���I$!��!q���a""d��"�!�D��Q�B����K�Y�ra��HX?Yt�g,�]>6�M,Z�*;��d
nt�0�uU@�'���{�ar��:b��5�V�N&,��-Z5�3s_����DS�(��e��CҲu��0��	5a7�Yz����=�‛���|�#?�e�u<�C�<����F����&���q�d�`�C�I�[�Y�ԙ����^D�e�OV�q�S��G$Q:`���S/*Bl)�uiBN�p��� �\ԡ�$�C9F]��/�<�����}�b�;�k�O����ͯ?ϐY�S�?#<���UiJ�(�%Uj��7�UF��y�)�+(.�a咝|�}�c��^�~웒�R9P�.�˃-�Oj���օXD����!3��IV�'���P!	����'��5$��)Ԛt`��=}�x(�'�0 {���P���y�"Ծ'�~%�I����U�=���H��$��o��01���'�lQ��e�;;��<�ȓy<��@`޸Oa�S%�!f︈��ɓ�M���
m0y�M,�3�>8����2Ƣ	��KR!02R��$�xL�&�߬p�*Q�NX���ݺ�_
!����50k�|B���I���ƧB�Z�H��E<��O&@�n
�JuriS&�Vq��x nyr��ٿ�f�:�c]�f/�C�	��x�ҷ7�,�� ��m�p�ah� MX��d�̟�������Q־`0�؜x� X�"OB��ϰ=�a����CM�L�@*�)��ٷ�',,3�ϔL$�ϸ'g$�)'ݟ&��L��KE1)�,5b�'��Ia��Zjip!��'r�<1� ��t��ȪQ��&W":7M^y����$߿A��K��X�:�� ��	3,O"a��nՑ�CT�X��0GC,���po��E�8qV&Be�<)��O\�!PB�*'"�L���(#*Ŭrla���a�O��#H�S�$@�@��O�:���'�I$�T�4��M���tnj��#�ܰJ�I��Ȅ�?I㮆������D:q ��
2U�n�%@��\C�I�(n���1%��$�M�c�@���Y`��QW�Q�
"�%��	6p70��2zt���#�.Z������r�t���+��asKQ.b� ҂�pO�l)�\q�TC�ɩV}��z�$Z���F�O�R�<c���B�_�9<�h��ۈGnQ>��`�L6�%9".F�O;�X�#�2D�� ��!r���␣�`E 7,�{Ê�8b ��&Yyr�K���d��
�Y�-��e'p�{E�� !�$�#�B���Aؐ�| ��C�!�9P�"D..���Ça؞�rʀY�Ha�M�	Z=|-I!.lO�0E���e)"����Ґ��D˜�9�*����'F<�ȓ/0d����,.1^aA�\�S~�yExr��o�`�F�4m�7�HE@�T�$Bܓ'#���yR!��$�~�i��J�nXy�c�]5[R8K�'�)�����˖?�T��X)�l��)D�89�L�a�@42���C�4�w�(D��y���&*)#c��
�J��P�4D�\�R��k\	�បAc�a�R %D�X��G�=��#�]A�<!�?D�t'g�s�����#A�~KX��>D��H�%�=Mn�x���r2H�2j!D��ْ)V2hY�֣�$E��ڕ�#D� yS��^�Љ����<C�P9��;D�DeK��~<y��B�tj�s�@,D�� ���H��!""bA���L�06D��V�޹[N8�qp|R!a!�(D�d�@��d�؜���"�t,@wh;D��;��.@�h�3eR'/�@��R�5D���Ѫ��_ܞ��gI�'1�d�2D�J��a�h�I��B+�D�B�>D�x[d�[#�Ԃ�c4ق�1�0D�� "-�'0Ȣ���ץG�Z�Csm<D�(4��&��I:����hr&8b��?D������y)f��P��ْ�ч�ya

'C<����[�0�J�k)O?�y��C�7?�����/H>I��J��y��-1N���+y���Tn���y��O�~�,Qb� O#x�|@$�K�y�˂�_���B�l�F��=�yRJ� cr��CHV>f�4!"�҉�y��N0Tʶ}�1	��M��#����y��J��b�:t"E�{͢�X@�Q��y�	"/H�=�1�b��Q9Qτ��y/��H\��'l�)@�ܐ�[��yb��!��`T���,�L���y���.C����m�@�v�q!Ү�yOّڍв�b����b-09�!��,�P�������R��}[!�DY�,�J�[�6I�fM�a/!�$J�&�2p#��Ҽ"~�:���$D!���M �[�`ɞfi��Jb`O�;�!�DRa:��X��/ �
�a�h�-d!��>z֙Z5�՚V�J�m��!�dM9-b�C0&N�I:^�Ҳ
�;g!�$�e+�=�N	�90�}BdLP>x!�$B�0Qj5]e�p�4ˆ2)����wLTP��%pF-���X�X=��QR&��l�#K2�lk@E�3b?��,)�����.yx�20�E7>&29��,��q�Ͳ@	H�qb�1}u�<��X���իA�;�Jc�JO�<�W��0mq�9�� �8 ߪ�p/�F�<�7Ȁ��S.3�D�XP�OF�<�R��(��t*���2R\���]A�<I7��=4�R�37.��&v�Q&%VG�<�a��� �
)*@�
,D�z@�Xo�<9&L��zAf{� ��dU�7�Sk�<I�C]�0=����:���X`��e�<)�K�;H�X ��VǶ��D�<eG�	��b
��<�D�`�b�<� ���P����(b��!c~p=��"OZ��\�-B���źZ@�1\�<���pj
��C�'2x�R�F[�<����.��1-�%g�N�J4-�n�<I��-(�ei�+�	x(����m�<��n��*���jԁJ��4l�<���/Z�J���l�XX��i�f�<q��*�#��)$�
!��~�<��C�r��BQ��f#�
eXz�<a7$��pIJ�7R �A��K�u�<�1cC�8R�v`�0t.x0�p�v�<��J@�xlPK�$
�2�FX�+�s�<�'.r]�9�4��x#����G�K}�ș�9Xl��	���� ��HO��@�� nMpS��7l1�<(T"O8����Ln 5k���j P"ODn"�=�t�PH�
Up�*�1!򄕿?��2�$��=��G�!�$��'a��&�ٔ4|����5�!�$�@��LQwD^63�f�e�U�-�!��ľB4|!�	�#z�����6.�!��	4��f%ίnT4�����!�dߌ^���G�%I�-�B!B2 !�D^-������.+ ĳp�I�0�!�
�U���Y��� �mN� �!�$X9�� ")n��K�!~!�$JR�RH'�,v�0q�Ū�6<�!��Դ0ђ��'��p<̳1/�to!�$� >�q&�l�l( �� #�!�$Ԝ�JE�s��]�p���� �!���D�ӱ��Xffl��MŜN!�Bs�9�&Ė<�b�05i!��@~\�Cb	��z����Ǫ)7I!�d�@�2�в��+$j4�1�J!q�!�dҔ�� ��!��a����jȊ �!�$�v0�ѭ�������c�[�!� N�lj��y���h݊ !�d�:6��q�іqɮ-�@H]��!�䌝t�&�#t&��}�X%�%�1�!��\y� T0��*���{Q!�D�([cn�����4������?a�!򄆜2��t(fW�w�*t��"-�!�D�-��a{��2�0��#Zt}!�K�?�N�����k���3�[	w!��ܡ���+��4*Ӵ��%b��!�D��o�xE�$��:	\Ƙa���L!���|$��)AO׊�@�	%�K!�ă ��'(I�54h0&��^!�dj���$�],!�>�BAèN!����ze��&+f�v�3�ť>�!��E�L|"�"�0\u��@Nϡ.!��$_ ���n}�����E锝��:�IڇE�F��U���^�R-���`�j��(u�1���E�	�X(�ȓzB|AP��UV�5�á�"�&	���򼃐�C�x7�SrKG/gPd�ȓ]5�][�#7|�E��o�fp�ȓf��2�"��u�RٙS�Q�Q��a��B��i�C�Z�t��I�i7:��̆ȓ{�Z���mr�h�D�m4���ȓLݔhQ��� 5���@&M�D�l4��x�4�s��R�?���p�¢��}�ȓC�M+3��	��ՐF�_�R�<̆ȓ qȅJ�m^hy��(!�z�a��Dh���%��j�0- �eǱwه�S�? ���K�a��{6�[�P�@� v"O �Hu/]�:�8��k�Z���9�"O>�#L[6r�8PR�폿zh<�"O��#�*�K���ʦ�U�6e.E["Od`:w�	�������\4�q"O8aI���y9�IM�W/��	�"O�0uc�4�$yR��� ��""O�XSf���&D�
!FQ.R�PQ�"O��ٳ䔔Fΰ�&�� ��4��"O$�C%U=>$и�DJ�HjJ��s"O�q[�n��@�X1$K�AZ��`a"O&x�0&��.�J�i�dVe#ک0'"OI@'ME&}%z8����Wpp���*O\�p�{�`�����U��'�l��'c�Va�դ��M8�c�'�T��&�+d�FҧM�

%���'�@��"qB�+�I\�z�����'��,��!O�&T	P�޼qZp���'�Xt;��C�G21ڷ�U%hA���'|Kb.C�'�}�&MM<`\ ��'���cD�"-7ZT!F�,k���
�'4d��Fוh|����&UҨ9	�'@�e@ ��44���⥂D�uX���'%���N�2��Ԫ���bP��'�� mن,��TIq%&Ո i��O���Ӿ��Db��/d�
�d���!�d�7p�ܴk�m�\��d�ukH|Fў���E���
�bR?&EJ�Q��=B|2B�Ʌ5��J�'�OH)	�&]�r�ɵ��?i�*�!Z2�8ċM�F����JI��|iT�xb�˸���)s���viz�:�k���yY�?B�ZhL�l�ԁ�bб�yrA_	 7���S'��`}:UP�i]�y�$^q�6��tN��W9�ܻ@��=ў"~�>�$"��4�ȕ�A�R(C����%Yݪt�>}G�XR2��n�!��W26"���L2����fh���ȓ�BikT�
�d5��� �1�ȓ J�e�b�� �~XX����9� ̆ȓ4ad���F5m�$T���.U!�ȓ6�Z���]�"�e@tnL�x�~%�ȓ.�>�eB��[�VI��c�K�8��0�J�22j�'&u.u�*�.�>8��H��� ��mŮ��1`T�Z��ȓ��@+ ?e�x$���,�h��c  ��D���)#ˏ�.� ��ȓTE����8�Z��d��I5�L�ȓs��=��M6g0���+@�G��ȓQ2V��b�$����%ޫb.:�ȓ"������+K�ɓk�$����X8L���",)�I��/��P��$��;��Z�B�26�}�RB��t���i(����
^�b%o�38,��ȓ+d�PP�;0�D}Z�N�&��Ԅ���TfL3w��0v�J��Ɓ�� � ��D��s�&]�d��Bc&��ȓ�0�X0�=���[�n�=r�|���-�⌊$HD!��9��-ېs��\��'���2��#8d�"^q#���`�*�+��ݲ��b����>�t��?12�)��N�j�1)�)c
���g� �y2�VL�͓!�Y��;AJ�#P�Q�����Y�zF��ı�U�sk `0f�>D� 6�E�:�q���)d��ɕ��Q�^��r ~� �CŦ"�-�Gꄎ��(p �'c�O"�u�F*I�"T�̄ ��	�B"O��B���l�x0G*��Bx��Yc��}�(���b�z��#�I�qʕ[f�P8JfC�� u�3%H)��Cp�q�ډ3���s�I�*]/4��%Z��9$˾�
��:D��KE�&=�F��AEO*p�d���8D�@�U(������\�.� �5D�Py�-?�V �4��x,Z���K1D�(��fLV���k�(�T���+D�I҄ .w�DU`� HT�P�H(D� ���J6Y�,ui��R�c� ��E�%D���A`_�n ��a!Q�#��Ń��"D�T��- ^n��g�Z>E,���O"D�ؙ�ND�_�����E�`9A��>D����
9|y�"ړQj�,!=D��k�lL�P�0e�gmҿu���s�/D��g(�c���n�!]%Ĥ	 L-D���b��*T��j5䙣k��!s�%D��C`�Y#nǒ����ձ *�DA6�%D����K<�t���b��(���@s�#D��qV'�|䈈S�l�%й�Rc7T�T��]�F�:���C�%%ڮy97"O<�8���"�*�ɖ�ڞze�#�"O�H�lэ&��pPd��4e��J�"O�X+U"�:�Ԍ#ŁP.Gj\:""Ox!j�
М���p7a}�f��"O�(8C	
$"���@�o޳l�pQJ"O*%�t-�|�l�RshJ3J��b�"O���6�\ �,<R��T(Ѯ�+0"O�$QU.@�^-��b�
m$\��"O �
�+�NN��k�
=8��*3"O
a��Ǽ ���5���O�Ҡ u"O8�۶$�;S.�}Аg����Q�"OР��IC�骩a�=:��:""O&�:�����Ysa^�h�
|h""OF ��N�War���ǽ �&��r"O*5(�/ͮG¦nF)tJHS�"O �a�F$ W,����l.ˁ"Op ؆O�>�6����@"e��8s"O�%1�e7nH5�,Y����"O5��O_p%b�X#�=wpmp�"O,x����<�lX� jfhhG"O>I����k�&ò�@cUN��$"O�!��������.�.֙��"O\�BMP2J�B�*@`�;g4j�HP"O�u2�	�3X�&�䭑�|&v��"O ES����N�	`���7��o�!��t$tYH ������A�!�$��kO���VGx�Re�P]�
�!��تF̌��E2^��H��Y.So!��ޯ=���� (��U��1��'5�!��ȓ]�Xl��I����	f�Ek!�ė(Ty0�a���4�@��
�P!�S�k��*w�G�R̞=�[�y[!�M�B\SDɮ��ٰ�$/U�!��l�}�P�X$x����%醦qK!��׏;g�d�Ǝ&��`b�H��WX!���\f�Y���(Gl� �GhR�87!��ߦ4�ޱ	0��<����G���!��I�&N|����� �yZ4ņ�2!�� �:�V�r�ڣ ;�LC "Ж@!��� 9\�c���!x\�6J�F!�U*<=z�L�5͚�hF�X�!�� �Ź�(��MK��j���p�$Q�"O��;�xO2X��mZ�_l��Ie"O����/�A40���+�	h�9� "O*Y���7��8�_-K�`�G"O\TH�.��<x���TD)M�0�"O���đD�� ��c���"O\ԛenQ�~�3�l�;�y�"O~�a$��,y*ɍ�(��"O;6����ϵ ���u�@�~�!�$�Yx�\6
�-Ƞk0+[!�D�:ǜ1��%E��@ࣃmK9m5!�2-v��I�N� c�F!O�!���O�Y@�]�x5P�/�5Pr!����\�u�D�I������e!�D[�?���;�\7Y,0�p�N�%G!���M��eْ���>�BX��V�W.!���P ^�+5� ᅫӹ*!�$Q�~) h  �8G��`!3K��I�Ir�9D��I�p��1 ���
Ǹ0��c5D��z5��Y�\���#K4C����i3D���� 2j/��2���gP��3�3D�� �q�a��#�(:�` �+9�}J�"O�;�iü"��ʒ��>6��"Ot�q��2��,27�׳ |��K�"O��*�K�E�h�p�#ƭ\�hzb"O2��M~��b�L�I�6���"O� 1����k" �K������"O.@bD�Ť)Ѻ�{" R�6E�r"OP�T��8�%Y�6]k�5�"O^����P�+ɺ����jA���"O˕�էS�L��旲}8b��d"O�
�EM2!���f��4@�q"O ����ů-��q6G�9>��X��"O ���"�m<���l��R���"O4���	�N�p�J�lIO�pŨP"OH��r�Y�#$.9�u^t�D"OTX�D��F�}�׃��Y*��'"OA8�
 W��4��b	.p�Ή�"Op��d�Y�w���XuC��N@a�"O`�xd�)$ ƁeҔ.��qW<Oq���,sR Zl�&xH��!5��Dr���&扃mO�,����I��0qf&J�:o�B�I��K_���a@F����	��HO��fA|�;1l�#0�0T�*�1l�C�I"��Y�Z�R�p�2�Gº��$8��'�g?م� o����E͓��
=�	AL�<a��"7=��"��Ȥ]ֹ�w�AD�<�c�=o���њq#@�Q��F��&�ܸ�C^�0���'��&zv�8Zs�3D���2ɑ$1|�ɵ@JB!�����2D���6'âX�P�
$�U	D���i1�0D����$ܹ�؂S/�5lp�#�2D��������J*��(Dx�h6D�2��R�P��-�M~+4\���4D� ���F�aT��f�	:�.t�P� D���S�<��p�L�p!c��;D�����Rt��"���v�ؽa$&9D�P���F*�zM�q�ŤF�x�PK4D��I�*�U�-�a,B�T��� ֢1D�,�dK���H���F眵��1D���b(�*.���(�hX!�X�b*D�ܸ6��e�)(1��X���*G�(D�$��:U�����ڱ^b8š@j&D�ċc�G����+����-&!�fA#D�d�s��|�*�j��W�m�$0�l&D���ؙ#�P]�Q��	"8�7D��=|V.��D�6�� �5+)D��В눘!���B3��64#�L�� ,D���%E���b|B�H[)L�84�&D��
��G�^y�#�ׂV���y# $D�,�w���T=��Ηin-8��-D��Y�#�ܑa�!�T�@G'D���
��j�ڴ��'_�P�c�$D�|*�)IB9��� ~���[U�!D�LJ���+��y���_^�<0�k�O,���	�/���ݢSv�A0&A&F�4��dC%"��'�\���,ϛX��v,ɳ��d)�'�|��PaЪ
�R�5Ƅa��z�{r$�0�O�O��<yRE�m�����0i|�[	�'j�E���܎r����R�rmp���5�	ԟ"|�'Vyr��ӹ}H7៛F�@y��"O^X�v�Ǳe��4r7DN� ��R�i�.Y��(�bd�=m�� ]�mzp���IO�M0X�{"���^�B�0 �� ��C�ɱ&��Z&��r�$�)��Q�\C�)� ��1aխ3C8��D �C[ް�"O9A�l�]������@bP
�"OLx+�	�;�L���Af&�زC"OXL���.`#�O�#���ӳi�h��	[Vq�dP!Q���c�œR�P��D����+�V��a߬L�*M��ՃUȇ�J�69k�/�28�n@ʳƒ�t�d�>)g�3�S��7��(��'�Eu�<�3MC�4�rC�ɛ4�l)��T"%�ĐJS�r�C�� q�Lh��AB��lY��%VB�I�=�V�I"EF�M4�hYG�P	V �C�I>V�.u�F�9Uݐ�+��W�\C�P�����J.a���V�|DC�I���]�E�6@��HH�o~C��3)���a�?f�������/�xC�	9V|D����W:��6�ƻ=�~C���J���1J���r�	�\�C�I�%�TsG�_-O~�"�
��B�	������(m�p��Ԃ�#Z3lC�	�G��E:�N��+h ��$Fͺ}>C�	3Sx��A녠k
��k�Ƌ�kC��w�̝� ^�7wPp	��4Fn�B�I�M[��4:���d�$.�R���"O`����@:]�	C>b�l��"O.�S֋�5W�tbʑ�M��J�"OrM@�R���T8��<����""OH�
"�0A�m�vʌ*�>�rB"O�z�D�D��pbT*T� ��ų"Oj���1c�hЃ� ]p����"O ]h�K'��(B���aZ��"ON�ѶcN)pT�	����&v8L""O>T�'��'I[J��5P."��d"O@��*�Vuj�.ɕ1n2"O�}#F��;Sa�5*�L	�`gx9@�"O���$��?���u��aw��w"Ofp����q���)?fxy�"Oȹ��%Y�Q�$he+ΜZE����"O�!A��H�J�P5)���9[)�s"O>���ic���C%��x�"O��k�*�Q-�`E��b�y��"O�1Mկ:�ꬁ`優,�ڑۥ"Oh�X�m�%����4��?�@��p"O���T�ŷRq��3�CH�ҹC'*OX 6i�n�)�A�֠�h0a�'�E�v���	�d�H���`�b�J�'��à��	
��ˀǀ
�����'Iq�ՂTr�]��яM����'�,��*'����5�ՁH�n1��'�4t�e���M.r!�u�:R`��'Բe�V
^(L*�h��դ:�2=p�'lF`�i��n�\�ʄ
�akЅʓ�(v�X�Mq�Pk��kzD�ȓ?�}Z@@�,�D�U����8\�ȓ=PrdBv�P�C�M�(%RU�ȓB�- �Ƀ�f����fG"��ȇȓ`��p:�儰0��Y��D�D	0,��G� x����%J>NT{Ĩΐ�$��ȓ>jxxsw�D(Y�,Q�b��f��ȓ7&�y�m&7@��.P_l�ȓ*d�(u� 6�~m�p���e��ȇ�|�l)v`ռB�4M�C	,a�Y�ȓn��#f)��:;�����K�&��ȓXQ��b�A]=K�Q(5��*�Q��{�H� ��n�p��.��Vm��S�? �����7t�dX�d�!Ȣ<9b"ON���	��B�� GN�~h�W"O>�X��E(^PL�QU����k�"O@��hS*Z�fP���D�$����"O�L�g�^���D �u�Ĭ�"OL,���֪	�b�N�u��I"O���p�%u����nR:�J�h0"Of��1b�.�%�_;kz��U"O�-Ka��}Pr�q��/x���"O:� 3�<L��T���=5ڂ�B�"OZ C�
�  ��P��]F�/���P`�.D�(�� � 8&"�Y:����*,D���"��l��XG,B:o|���q�+D���A�Z�?8��B��ްZP���+D�����
1t:�˂�W_�Rt�U/(D�t�1�S!^�IK���'E|��(�@:D�L���)�"���C��I�`=D���vf�<'6���Ɖ��
V�I��K6D�`�c�/w2�YGE���(q!�?D� �����mP0=G�YF?D�2v�ٗ%�n�X��ڒ9��B"�;D���v�S8%& �j�U�7����C�&D��x���p���*�.W�2�Ԕ�fF2D��&�O��leb��G2L�xYg�0D��p��N*/G\�k��P�,.�,�
.D����*�
X`�	!`�"m "���>D�ۑ �*��d3�	�U�N�"<D���v$
2ֈ�@�N��$�DT���&D�(���O!���� J�V���#�$D����.�2��t�mG'g����$0D����/
+I^ ��l�&�E�8D�����ʥ@0��AUdN�BŬ��fO#D�ؚ�K�.;�s(K�yd���!D�`���Di+6�Ȗe�Ɍ �";D��`�gAP�*4{�-Sd�F�8D��CDL9;Itu��H�'l9���n*D�`p'!��q*��B�FI��`���'D�l1�b�,>q�u
f+ۖ$�h�R�J$D��pC��� J�Q��	Ʈ*�D����#D�$*B��=t(&�h�zHQuD<D�(@�N�Q%JY�he�Q����y"w`"9��)���֕Z�c��y��&LP��	����HHc��2�y���;&�h�"2���C��(�%��yB�(!�\��V�^D�D��h���y	?6�q5k�#fְa���y"&ׄH���l�)Z�x�	7���y�|��j��I\V�չ5���y�_�Mv����H�=��#�GY��y�!ّ2)v���.N.a�6P���:�y�Q!<rHRw�S
K��`��P
�y�N��p,����0�hU@s#�:�y� ƹ/d �@q��%)Y��AB���y��L=�x�FlM#(]VAa�k���y�?������(5������y
� ȉ�vl��i\ �:�%x̠r�"O�%�n��t1���3%Q�\�t�b�"O������0�d����I�X�T� "O!{3��.$Ex�',���+�"OրⶢZE��� S�0�X�F"O�d�.��0�EB&�lT(�"O��×,K(�����Y�A��Pz�"O��(�X�j-�ِ�

x��v"O�݂f�WF���8���r":��r"Oz��󏌾F���+	I=�x�6"O�5�fJ�M�8p�Ab��)�\P"O������|�����C�0���B"O�=�����å���H�ʐ20"O&a`1*�k�dPBe��&-x�Bb"Oā�%�ԲP�)�S�<��"O��j 0\&N�1(LA�营"Oμ�����K�dI�6g�9�F��v"O ��!B�,��,�F���r�"O���㦒�PPP���ޒ;�0ͱD"O|9�d�pM��� �Nu: "OY&�X�^�(8�d�Ѐ?�b`�!"OL�IΊ���p�(Y��ڝ�0"O*�ذ+�+�@�G�i��(�"O����*Z��愍&�M"O��1h�B��,��KK4c����"O�%�ơE*a$!�jH�]�mU"O4P#
��rU	mo:8�1"O���X#!-���a蚟UZ��1�"O� �-Ny*0�-<?ε�4"O��h�n�����
B���"Oډ���?��Y`�ƀ_W�J�"OB,#��G�"����B�y(�"O���G�1D�p�ǱqM�Ɋ�"O���IN�#6XA l.C
���"O�0�@)�t�5� {��;�"O���𪞷%z�I� 7Q}�L�b"OTe8��'e������mM���"O�s��Ŷm���jQ/ӳl��x�d"O�1�)A-�µ��K\�B4�ܱ�"OBr�M�^Q�DXa�-l�r��"Oq��	�D�"3���#V(��g"O.����	";�h�5ĭL�	U"O�@M!U�!���5�@"O �`��Z���%\�{N��3"O�m��-Ӹ��$`�(N�h�p"OL�J�iT*%-�D ֥�'mSۄ"O����D߄8�����RD"iS�"O]*F�^�Gј��ĭ��4h�(e"OP XgGE�L��$Xg�3Yr��#"O��*�eҸ-��%pK�5��=�"O���0&�#<
�%�!��>��"O�i�b��;�.���'p�R�+�"O(Rj>#z���d�Ɏ��)@�"O�̡��ؗkA�Zv�T t�
Y��"O(�Ӥ��	'�vY�,@5M*hY)T"O����,�3I�
MJ�%ѻz#��ӳ"O6���^� KBI�Ğ���"O�p�r�_��$��C��f���'�$[=@��ػ��r(�xBV7n���
O
m���ō\Y�Р�=>���"O��ңOƘ[��� ÒO쀊�"O5;���B�顢I �50ѣ"Oޡ�w B�$%�'�
 t��s"O~0�U�R�S���@��3k��-
�"O� B8C�+�T�D��'%jH��A�"O
�R#ʌ"rĆaQs)L'!_JT��"Ob�y��
ma���ǁ&R4�"O
�H���<�6��2�H�jJ�ӱ"O��U=S��h��$�Ƽ��"O��Y��}�PH�� A���iF"O0�{Ч�`%ԡ��d�a$����"O�2m�!W�̹Z�¶W%���"O �G��=Kt4k$a�)|j)	�"O�$�b��!�`-�c`Q)BZ]�#"OP��芖sqd)�d���k�A�"OZ$�@j��mn���GܣSvx��T��%����g}2ƕNq�`R�Ŗ0o�E���0=��{�&oLxT� X�"���2�.��\C�	�G��u��ǳ@�Ҙ�թ�6C�	?[�%�d�,��ڵ`��1��B�ɦpWȅ���#=�J��U�^	zޚC�!	�P��ɋ+�l��s�\~��C��?L�����E�6�
��:I�2C���K�&�
6�f����,mG�C�IKt|�ÈG�-xbe�V����=�ÓcCP#�i��}�T�Jflǹ"X�х�X�0�#�̞�����)]�%�t�ȓ+��!�`Z���!�t˚�k`�r���s����	<&'��{�R���a�5D� �l��~Ԧ�[�KQWaN���� �$?�SܧBV��b ʷ{��1C�'h �(�ȓ_i���U`?�x��&J%r�vC�I�~Ͷ G&M�|:� ��c�h\C�ɦ	~����T���c�A�dFC䉻n0�c��9L����
0b��� �	.y���/����ł�I XB�I�\����$�� t��	e�ۗ/blC䉹LRX}�ţK�|���Y��PC�	�	f���#�SKnDp?\ B��	>�~����նUgH��%/T��B�	+S��$s��q�NT����)"��C�	/|q�SGJ��D`��`�}ƒO��IRܓ��';��!��|�y��A�ZQ��'3��!���g
�A�EN�ڦh9+OtO^�S�>Aƨ��0/8u[T�K�;���[-��<)@-To�� D"Etґk���b�<��(٣M� �%��*m�x��Ox�<� �C/5i��GX�st�#�j�<	�ƚ3'"rȒu��5|����S~�<A煙$�	qeݦia�Θ�yR�B�2�r��AD�i�n�"P�J��y�@D ���#�&M�Z�esg�X��y)3ci&ћ�D��Ph�L*g���y�j���z�x�؍tި��BL�y�CV�}�t�*�ܫo�6�`�NA��y@T|� m�6#�Ȯ64�5�&i'D���a��riQ&�Ϯ=�E��G#D���Ǩ{������Z\�e4�yBC(�JI��ʘ?)*�H�睿�yR�j�r�o�=$����ٵ=�!�Ě9xz�ͩ�V>�t�a@��!�ď�R��ͪ$a
�D]�0��\R!�
������V5*�Z1��n�K�!�øb�4!�p��h�s� ��g~!�� q3d�pJ�@�ȵZ���5w!��$��|P�°z%VyQ.T�!�5�y����Y��խI'�!�D�
|᢭�̆$x�r�s�ڔ+�!�� �5��o�$hi"ˢK%.!Be"O*QZ���v3�!��j�#(�u23"O�}�%jQ-<ʹu��J���r	ps"O���VN�d��H)t�܄ ?��{�"O�x�4N�&���(d��3"�B""O��K�Lϖlq��x�n\�O�P"O� s��%kd�*ՋȠWi ���"O0(���U���"�D�nJJAZ�"O ����O)�9!&���++N��3"O�%�`��)�v�4��i��Z�"Oj+f��b{�HkC(]��1KE"Ox�;�j���C��O��0,�d"O����B8@�:l��+O�u��X��"OV�1#�ĚkSp�{։5kXj��"O���j�,L��T"�M���"OPh�'�Z�Z��!�ec�{����`"O~}�#!�U���EEN}�b�q�"O`8�o�|��*J�S\�}s"Od��@z�պ�I��>Xpe"O ���ܩ|"����֏U:"p`"O�D��h�>[[�� �^4��ˣ"OH4X6EY���\/�-0)�(u"O���!_	�	X1��
s [E"O�� Ɓ�9�δ�cL\�m�l��"OH�� ��%P|�3�H�<4l�˗"OZ��2-Y%/�,�G�&-��"Oiـ��{�Qi��ܴE$*�D"O�QuI��H�Q����9��؂"O2�Rv(�$d5`͸����N$�G"O���\3U�	��|�l�w"O
}n
�y��!/��k����'2D�p���#� �q#D�8�n4c�0D��@g
"׼� F�f�r�a� 3D����Z�y�`��#Ęm`�!�'1D�D���#r��$s�	�� �ug/D���V��|�y�rl�*��a��i.D�T�7�l|�l"aj��`����`-D�0�cdܖn�:�G���*��Ս,D���P��
S5]���	�gP��C�,D�����5��% ¡H�D��,D�x��
��-Z%#�&�o�$�bQ�+D�؁c�,��SGN/,�9��)D�\���_��N�"v%�z����e&D��2j�&X�d�WO��h0	�%D���Ȟ$�N8��%R�a�v)
�  D� ��>N����0������`�,!D��r,�6%�eQƄ\�gǶu��1D��
�L"7���±��s`h �3D���4OP;Q�ub�ɚ��"2D�ds'�G
b�XM�+>���u�0D��Y�@x�<pS�"-�\��d�1D�<1�fX7�0�BԿ`��� 5�"D����*ث"zـU+6O�4�q�-D��3r�v<�ȶ���*���ZT�?D��z�O@�_uh�eeH8c���ӗ�>D������b��2��F�(�b� "D��@��	y�d3�F�=~(�sW�=D�d���#~6t���H/�U�u�.D��!%)[�{UX��Cf�ԕ)%�*D����ȅRQN�d�Rm؎S�B�#l~��E��h��H�-tB䉬S�Ĵ�
�>}���4GN� RBB�	�|$Ȉ�7i���tp��O��G�&B䉛N��8��D#e�n��J�[,�C�)� ����R/��@���y3"O< ,NsL�#��W�6��yp�"OAB�Y�b1m�e %��)�"O ��ē�~�R�� �ŏFPB�C1"O�T����-#Ą���	�l�PlS"O������3k���0�%ըQΚ\�""O(|��
Ѽ��j''S�d�+�"O�d@���88V�#ͬȺp"O�݁cj^3/�D-;!g���𱉠"O`a�$� �p�xR�N-��|��"O80zS��;����5��	N�,i�"O���5��O��i��_� `7"OX{�o�Y�ɗM��I��5D�̣�E��J��C��_s�x}c��3D����r+�H�A��Oc,��3�,D�������W��u��DW�9B��3%,D�P!'M˙{�� �.�R�`8�H*D����D���� �w����% ��#D�x8`�/I�u�r�K��A B>D�(n��oc�MP�%I*,���0D�<�1�&9ox��E��Te
+D�H �������ŎEC����c&D��sC�CD`��$�;A� !�t�>D�`PխY�_�BTE�v��@��>D�`��G�D�4���i��`b��7D�D��D�Em��5�\5 y�`.*D���4&ޠ=t`t8��Z�D��5��D.Hl�1�����y��	ng���� ~���z���2bC� Rߞ�R��E+`�U`�m�;NRC�	�?�d%����3o��Ȁ���f�nB�I�__�i�f#���m�ׅD:6�C�	7V�XŻ�E P��X���=�RC�ɭ߶�q�؏J'����`(8'�C�ɂx��ѕ�H�G�J�韭qJC�I,6~8�ȑ@] |�F�P@�\�n�<C�ɂ5����G��0m�L�Ý#`�~B�ɟB����I	#"���E(�-��C�&܀I�)ϐQ�����
�QepC�	x�bȊ��E�8`ژ�
ūn�VC��!�Ȥ��)J��i�n�C�	 �`�F,��Hh ��c�W
m����$Y�"�D�
5Kv~k��Ӌ�I�%�״��X�t�7�O���m�����nTWH��G��/�2%yP*�0���QU��x�$o�9	Y*�e�D���R�M��yc�3x3z�po��g4�Ai1�y"�G>	� XX���s7#�s�OLxԈg�T�01���@�S��B=��'��LA���|�2��(<!���'A�$;uۯ/��E; �;4t��'k��+�����$�M�@�K
�'�&��G6�8!Q'�2��mS��?�S�4��%V�-���͈E����D�&�ye��3��(� ��8��'�<}PB#=E��'^�,�%��}��pi6@��BD�I��'3T=��#��<<B6�]�) x��'>���!O����ʇJ��ݢ�R�{5�{�_m�R�2�t
��!dUpF�8y�"���	
H�w�ăqx%��L��o���!��)*��T�N d�s�������C����y�č/qxi[�hȞm�q�2%А6Kڢ<a+�"<����?:М:���%ɐ9��N�<��C�=��Ւ����T��1�	���{@�Ol�=�}��iK~�z�z ��8|tM�y��(Ҡ�xR`^5Nnl*��;T������'azB̞	w]Z��񃆡*��@E��'�XDyʟ�� �|3�"��pĒD�Q<�!��"O.�K��_�&`*��)�N�(�s��'b�X�B�ļ��1��E�*�n�c >D����D�w��x��Mn���;��-�Sܧ��l�`$�_�`�@��.cp���ȓQߐ���oՖoTd !��CX��?1�Z����`)͙@@l )���N�D|R�(�E�dB\�ȼ�U�<�8c�M	}����MB��+j�>����G�=8�d=� �Ⱦ��$#��ɹ~@ѓSi�����?i�<�_�*����b����axB)T�&� �`�O"�kb��M��Lhu$��Ɓ�ׇ)T7��/�OpU�a�ܩ}{��JϓNH��`�ʓ�Y��l����#w)t��'Ob��ÉC*�ء�I�,%T�ʔ��=���"t!`�����h<�4�
6%�����Nu�h8�4G�$YJц�p8�@��f�w� c cƛG����?�028v�y�O ,5k�]�#��
p�k0cFE��B�f^��Q	FA4�ype؈j��S0�8�O�E1�� 0<9P|�PS^S��S��	#<�1�CE�
�.��E=RD���.280X`��'_V��3uD��?��݌!�]Cӥ�� tP毀J�,s��D�4r�پ�?��,͊m���C"�ϹX&�2�Q�|O �`NM=%"�"��,� E��������{r�oݑ�f�{�{]����ԥ5RBuK�,��`�'�� ��
)� �ɗ{3�P�) ��NK�/��H�W�j��S�Dht]R��3v^M���ʹVNH�F��$;TX���6Y���9�܈poU��ʅ&|���r*̭XW&Q�^�t���7Z���	��\��M�4��
02L�f�ה0���qϊ��$E�%*�I����Ɏ1��šcHZ�:]vd*�AT��|1P)K�9�����'0��a*4E��Cq���D�(0�q� ���Jݞ-����ԟ� a{b���0<�4mؾw���H�'vH�z��2=��H+�g\<�[�˺Mv���v��k�쑰t���[�3<��	�e���Ov�b&`ԓ��`;3E�5(Ht���>�V&
�jR�ʓ��|�4';�IG�g&L@���&S1�	1�L�j8����BR�p\RՃ^�GX�܊��*<O�5�) Ĉ5��J;�3�'ȼг Ǯ��m�q +|ؖܘ�LC?*�Ɣ��J�)�ۅx�6B�-�����.z"��t� �hd�� ^�PE�QJ�ּ�!�>�����
 �vq��ĮOn�����ݗ8�!�$�X ����۴*��4s�܅m�ڈ����:��U����3b�}�����C��<}���[2�@`�����zȪ�'����Ay��^�XD�$>��W�]�3�2�	�aW,]L�R��Pᆘi��nU�B��(e�ه�I#^ 	ˇ�(,��@!Z^PhE����C��=U�����)\�p�lߞ8����ӥ	?z'��
�e��I~>�2��ά_�D1aª_*kU��Y��'J�h��O�b�`	�1(T>[�qv�H�7�(���H�o��(˘1�ǜa���2"#(|*��`@�l��'v*DVD��pF]v���X���H=L9���?���Źa���ì�W����� W�X�� �D)6�.@Bj ;+JB�	;
h^�"��cݙ*�N
���'!�\Pr+�,�Yٵ&4T�ţ(O`���R��D���;��*�ˇ�@Srם&6R���O'�Īᄜ�I�x�yt���6T���΋-I���H�E���b�CG��� m�f���J�O�n�T�'Ҽ�0F�N�v�JH��臾@M�ű���
g�� תD�J�r�+T�_�-`���q���ow��3j��:Ǿ����8/g��BWު-�|��7�A�;������rY��"O�x�L��H,���%�+.��h��>��=��`ݺ����m�=�I�5�z��2�C�!Aџ�����&|��$�e�'K�����ܴ�k��(+�����Փ{y�4a���:7�p�b	�|�V)����ڼ��;���z�O¿%p��$����	����<�e��#�,�{$�O\������_r8�Zw���1�ҭ�,p�Ŋ�`ΠYd`	"S:9���Ǧ5(�#��4���dE�}^�"4ό4$�{���"�T�I�p|l�	A��m��A�b�=�Z
��O ڭ�I�yǉ�;@I�Ѵ�S�"�z����Px҆��'�AP�B�	k� �&HI�	e�Di���p`D�7D�e�dU�~Q>�<�wj��,M���3�B]b )�,��B�	+&�fY�VGϸ�����P��L�q	�A�'+\O���Zd8$���dҊ)~�I�#"O�i�0%P0�ؤ��B�1fjf<sc"Of����9&L�(��ƣ<nJ��"O�L��$���wO��	-��#"O�a	�IVrL��2����M5|�`!"O����\�4�0� 5t��"O�����I-��J��_e�@��"O*�g��6��{��Ҽ!0@!�6"O�\��P�7z�
�&\.O]�(r"O�ai�FHQ��Q�G�!D@��"O��p�C �]��Y7�0D\��xD"O� ��Ѳ�R>!��u P �1��"O�7K0��L��ҞF�L�j��$D��A��
x�tx���.2X���%D� UC7�~�z ��'*츲2
,D���wdH�V�f�Z���d������+D�d�'�4�~���$2'�ݐ��)D�<iP5wm��"Cx��yV*3D���"�2E�Z�"�L]=7%ȅ�6�:D���E��0���	��\+2<�S�:D�0@��/�r��WhP��(���9D��9�lL09����N�w p����+D� ne�P��SV�W�v�y+ 'D�@�D�
A �<or��0' "D��r
���ؒ��[�pXƉ#D�������d�J�A�`A�/D�L�s㗹c��G���r��4-D��Kb-�
�q)g��s�PAr�-D���WA=��P��,%��D��6D�j#�)�Cen�"n`S��4D��jw��G[n@[��Ϋz��MZ!L'D�����ֻ�ju2U���q��)D��!SN[���t�ϛ�*���1��$D�� G��3�R���YP)����9D��x�ܽ�N��F�Nu���)D�����x�2W\?O��t���A��yrA˪iZLȓ��?7�+�L��y�[�Yf��9��Q�")R5Z�&P�y������Qw�N�����C'�y�J� �|9u��5�t)H��y�,�)-�w��%��(筍;�y���48�6���.^�sv zF�@��y�$��(j� #�?y; )�����ȓw���0�'+E<�fS%�t,��F��q��H&ga|yKg��=�4��_�"A�AeJ�6�2��$��.�6��	��Pr�.�WWbu��D��n ������7e�-f(l�#t�K'Jbe�ȓsFx�fK��O��c��)� �ȓ*q��3�D6`ՆY;a�/e����Ifd�9Af�HN֝�&���ц�L���1a��k9D5!����`���/l�h�&��r���p�ψD��l�ȓ1�D|{A�#�bL��.NO�ŅȓD�P��*]����C+��Jʰ���m�d��B(e��͹3k�C^L�ȓ_)��X�'�-6����ǃSiDI�ȓ<��;���{S���ЃA����Z�>�۲�[�:����	E����7��;� ΪC���z5B��w����ȓb	���?�|���S��=��H:�؁���iol���g5�E�ȓ���V�,a�mb"mP�AS�p��m7t�@�K޲L�$4��(P�^��B���p�@�$1�թ�`�t�����UB2� �k��j������6V*}�ȓ0�l8D��#��a�I��8[����VPT+T�V�I�|y��ʫ&�P9�ȓG� B%���y��84�W
:��ȓx�H8R��	�@5`ѡw"�tɄȓ�����n�(�,��EF�M�橄�c'���&6Mi\�!2o@g����ȓQ
�CNXWE�i4�0�F<��ZA��# @�*>ؽ�(@03����2{t"W*,t �T �O	��X]��S�? dI!�(;+�RM����!�zT"O:u+�/�>�x��2E�>/���"O�]�B�7d
�KWD� y���W"O ��fPD�R��F�Ú!^��1�"OjP��$�x�CP�3$)�V"Or"�	�4��8� ��.xa��"OD���/iԌ�G��.CL""O0 ���;a���J����q+���F"O�ēթ��,b��7l٤���[g"OTl萎Q���l��@�6�tȋG"O���P!�({Z� ��ݩ5^. ;"O@���ԛ<���r�d�d��F"Ov���I=P�����Ŋv��`I�"O�T�FG�LUA%nњq `��E"O\ؙ�k�L��ţ���&�9"�"O|q��H�5G������°�޴C�"O:�+B�փIEP�k�/��
"O5q�$¥b�XB*y���"OPt�`A�#V�B�Z0	�%��)e"O
��cI�n�`�'G��W�	�"O�q�`�|Ƞ��H��n�fّ�"OP�qw˓z�$ �'ǋT�$��q"Or1�b9K_~���N�Ɛ��"O2�	��C*Z�����ѠJ�2�Qg"OZ��ăBv�]�r���(�2�A�"O�8j�iR:"xV�����!r��c�'��;�i W����lȃM��tQ
�'ڌ=ءA5J�tX�4�:p�ܵ�	�'�\�seD%EB�@�s�^(rR�9�'/�T���߀�4��a!mҐ��'��qѡ���K*YP��xl��'�%��7:���.[W��
�'$<	˦�Y�{_��Շ�?+�L
�'a���� �m�)��x�	�'�v�����+tax�
�ˌ� ��'�ZL w�Š"��<j�ŉ|�z��'w�L㰏,Kj�H ��V�i�X�b�'X0��W3?��#6b�0s��01�'� �Z!�ƾ[�`���ɜw���k
�'�0a2uaY>,)��іk�!~Љ 	�']j�(Q�D6X��&%�X�T0��'$���� F*rԀ�U�N�d4��'cƩ��L�T'>l��%� ad��'�U��\�D�gn�5PnH��'_5�٘�KT"��
hK�'�,`���1O6Y���_-|w�t�'�l@���1�v ��DX�y�'�v��P�!~d�t I ���a�'���9` ?�	�#�J�����'v�T��)R�c,҅��f�-xS�]��'�R�׉�3y]��U�Z�v�Z���'�J�%�Ȧ`�@�:%!�w6�ؚ	�'�J,�i!	��w���j}ND�	�'S 	icF�X:h��sH��Y@f���'ed<#6�٩nڕ���?9�>IS�'R�����V3����f�� �)��'.X��_jV�`�q�^�&mp
�'3X4�
�u��9!�(�T>i��'0�i V�qk%#mRU�JA��'8�9'��`�r��%���|�����'��Qp��,� �e,�q#ȅ��'��: *7+
d� @*O�q8|$a�',��(@Ň�R����pd��m�<AV,�/���6�B3U�$��#�k�<� p�*��#@ӌ�(vJZ�j
±�&"O�� C��z���#h[2���v"O\)�f"6J_�dj�T�j0�%"Op!"% !`�Z��Qi���ʕ�"O��f+�� L0�2z*��f"O�h#f�:<�
���MP
xt"O�M��/�pX���J�?y��RE"O�Eڥ���~�z��jM�Yn�<��"O��e%�����8C�=�q"O�VlK�v���2u�S�TP��"O�Є�$C��|���^[��i��I1��y�t��vy��B�L1t��4۶9f�|C�	�=V�j��\	[��su��(m�Ҹ�eJQ�W�ȅ�e��?V���&i�k?i.��c�@��)��V�4B��K0͊�2O��RQ+D�~�	ITjqb��>F�l�zG�Ndn���Y���I�fu�=�4&V!�y2,?�ĭx���?$<�X�M������/A��T�A��?��c��r,��P�o��x�M�
�2�Г�ܒ ��Y��#�7l�l`@��y[��D	(��i5��<\�hz���*ڜ����T�|�A���A�1����.���Qe�v�ya����u�w�d�K���D�^Lx�]�PS��x��6�j�+�d�_�Z�[P���|�4��[D��e��<�� �(MI�ءݴ ������ )��~� £w�j���M-	Z�0�a^;��O�U���ݱ0�*|Q��x�V� h\�Z\�1����]D�	�萹���Ӥ�@�����$�]�5���G|R/��)/|H� ��0j.f,��ʃ���$­ɰ��D�*�?Y��J	�>�
a�z�%Ɂ��R�!��hI@0��%0c��i�c҆;����t�ӹY#�}�
#�`�K52v|�0L�)?���DF!'�|c3`Ǆ��ңoʝ �l"��j�Ԉpa�Wx�Ξ�/����_�J$(�[�'��M���ކ,��((�`ڈ'���Sa�R�paʨ@U�M�q��P����U��N͛�[o�h"���I̙�B�?1���VD�l�c���pp��%�C��2��۝I�2��d�J�� [<��b%�]��٠P�)��c�O�h��!ڱ@��%j�n������8[�k�#�O��K��O�f��T��=�"�<����;cRc>��«�3j_�a
���<Z��r��Ňz�>�6%�'2?�}�������Q�B]:���oM��<�C�G�U��Tpu��<���)j���(�07����q�<�N΃U�"Х@	� ���hg�	��Z���OW�?e�"#P�$�lICנƷm*J��*-D�Li��0-b�"�K�q輳�M�R�蹦O�I�E�Y�g�ɶO�U��C��p��ҩϋe�h�'0�� �_y"�ʭ���|jbMA�PB���nу]GZ`2��[�V'CPI)��'k�,��-�:�kr��-Y�E���O���5�|ᒬ�5y�H�6Ƒ�t�	Q���?�;��4��ȏ�ǆ�X®�+Lꉆ��(��(��G@�/��:��7{�b���j@�^y�i�b,q��vo�.sJ���it���.V������« ��D��GʨD���P�XM���$>�џ �r�VA8P]C�'��:���p 
�kRN�7�&�����X5R\�� �'�Fq;�R�|��л�cD�t&�k���2�L�fv��I9�O��8?�3?�m�祍�w<��:���I�#]�+����=5Z3�NX�
w�U�9y6�:Ġ�Jqq�8�r����'��0&�&B��-R���
��Aj�OF}��!B���ؠnɯ�� h�fU�@��9j���M�E2����6Ϧ�E���B1���'���A!w����LA-}]����3)�(!2wI�W����E(Z�:$�r�i�$Us��[���ekڇeW�$�,yw<p���+6bf5�Ɔ��џ�Ѡ��w�Ȑ���'tʇ_�<�$�� ���Qg�Q�n��	��IP�b ��#��y�E��28Y���>'< !B�5��D����T ��?i1J� I�A�o� ABS7x�H��P�[5|��̓TdԎ,����`D}7��dL=Ul�X�0$�^O:����@�	1��	� ���R�!�u�X�af^�5L p�O���Ʌ�y픹4	��Ӗ��9���b��+�Pxb�ܚ��TTcA�id���6oc��Ȑ
K%@10��ơYr�`�&�O(�'Ø'�Z�jī�')^d�d]!e)��k�'�f]���#*Y�CF�+Em��#�OV,�2���p=����F����߂f|,��kQw�<�e�)Mvx ��>9&b���r�<�G�H!4VP՘�Y6BHH IRh�<ArDGz�ҵX���<�@Q ��Xf�<��Z
nB�0y� �R���f�Y�<9en�(����"Bب��5�Zo�<ѧ�ʳo�̘b�]Ȓ��ơ�k�<� �qxkF�E&v,�EJ
$G����"OV Qu
�|��!�&��o�����"O���e��ʘՍÖy<�(RЯd�<�K�	P+\t�@GV��	w��_�<��ؖf�T�!����^(Js#�[�<����b��	uO�i�nTW�<�C͇�:�V�y���i� �5�Qk�<��#�n+���Q�<T5Ҍ��gc�<	�F�'�25��:"�n���FA�<�l��L�@0x�|��IG�<1�[d3��9�	��QТ���J�<���X����G�F�� VI@�<��]�dPȠSAM��0�`��T�<�B�6�J��WE�	�6���K�<�o�0t���I�,w-F�@�TF�<Y#ϝ�����ǩ`���
Oj�<��MF:i���nY4H��b�<q�S?�q���ˎ��8UgVX�<�6�׺ $��'Â&� ���QO�<�D��Y�Љ��L��G�q��
|�<y�]���5��EN�� Qt�G�<�"N��*��$�G��x��m�r��d�<t!̆i_�My�Hӥ.V��:shKg�<��=B	h��w��&b�zG��c�<�Q%
��DԒ(��5��L�5H_�<ن%�<��� ��X0P�J$�aN�P�<�d�%{b�u�摳0Rh�	`kIM�<9Q _���[���-$�<00�I�<)3�5U$`0�f�����s]I�<5MT�hK�i�� U�5LD-YR�F�<��n.���O٦3%.a�RNI~�<1N9~&= �' P|�s�~�<i2!@'\zdt��J:Z^��'�]\�<�E&J���Z�i03*r��c�<�F�~
�S,�,+~���[�<1%���u_�,�v�Ă4d�P$�P�<���L��6�0TM�$�P�!�L�<�H���E��훼}���bKHB�<A�F�<�x�ɷoǼaZY[��N{�<��ȟ����E�O�l0���M�n�<�H�����3gH�Q�~��6k�<!�(ŗ8rl��^"Ur���A�L�<�4lʺY*L�3fa��1kF��na�<����/\NȀR���,W�lY��Qc�<��O\�p�u�E)(#@P)�*QX�<y�@�1����W+]��	�mUA�<Q���}Қ9@ĩ4t�ma �`�<	C�F�}����'�,`+2��Q�`�<�Cއ?􊙩�GR�9C���u��a�<�!�M�-蜥�v�d���X�W_�<�u�w�Vr��V3�,�kSS�<)N۸X�h,sU�ڈL7F��+J{�<Q4�әc ����j�PI2,Vn�<i�(]>o����1�!mo���d�f�<�rJ�O��q�h �CV�^�<�'��>aJ̤�t�G0����� T��YENZ�$�p��@7XV���*D�T�o��WI�j>M��&D�� Qd2uW0X
���582漣�6D�0i��Bm��=��|���v�0D� �!Ba?����JN�Rۀ� ��/D�ls�G��>�6-�S'@��~�BӁ+D��ՏS\�Y�E�_��$�21j(D�
�G�e��A���+%腊WG$D�� �肱님]�hs����fX�C"O�Xi�`֣VY6�Jq��c�l v"O�.�'"�T{"Jb* 	b"O��I��-�X�� ':�`�"O�0�^W�Uj���"O0���ݪC�D�⍐�l��<��"O���B='�Ƭ��K� r�أ"OP�#�(^�ֹQj۷:�3�"Ov���lC�,�ac ��[� �1�"O�㔊"ZX%���/��`s�"Ot��V�OU���YE��F���"O��rC�x�z�*O1v�ŨE"O�iog ���6hE,NN�њU"OP@�3LO����#<"8p�"O&��R��=z���`SPL>��3"Ot411��l�e�b�F&H ajT"OR�X7р.d�"A>8���"O��3�S#^<����N%�4P!�"O�T��-ń!� �KԠ�	O��x�5"O�����u���A?]�ѓ�"Ob�!4�G�yz�`���C�v���"O�)���ғ(�H1�r�|�t{�"OR�&.�����1� �=B0Q�"O~X1C��]��dO6" �	��"O���e�e:�c]�N���"O��a�f7�L�"F�-���"O���v���NMH'�[*a�r%K�"O|�D*cO�ⓠ��Q�B��"O�P��D�L}y������"�"O0����_�`l
����=m�e��"O�P*�ˏgY�d��[4��V"O" �&�<F|����h����'"O�q(����v���*\�<�.��"On��$�1px	���L�S�,Q��"O"(���ʒ�TΆN�$�Ct�C�yd@�XM[�h�L<m��1���%?yK�N�'��
�N[=~����F�7��y	@+蟔X�E,f��K�jE�ǫy8wiɅ^� T�H<�`�2�
oͪ�'	;$h�'�pj�YjG
��n�R̘�c�>Y���Ra�pS�B&��m��i� 
r����$W{���d�I��I��ha���߶� �K���+�$t�G�W�>��,�YI4��S(�@ъ���,����)VPĈ�*T-*�8�<E���e��u��L\�h�����+pjuR󤛫�0|�� E:,rɳh	m���J�-���'���B�\R>�0p�ԓ]�:�jP+��;-L�	�'}�vX��y���!/��ae蚟{y�cE��'󤘑V������z}�З�h��9�$�ДE�x8ѭ��N���(�j�LcIQ$a��p>�&���>��%L�6r���E�d�<���X)�% �!K��"��0!T�<�����1A�εJ�(B��N�<	G�ŵO�����mښUj��)�E�L�<���o&Ti�e�R1F1i�$Gx�l�'������#c�$S����� D�x"/[�
	��L^aܪh��=D�@2c쀳K %�$	�N�,X�( D��X��G�s���Z�kD	 pm�SH3D�p���U�V�턲e��)��/D�t��	�%���8Z���˱�2D�|!�н@S 9B#ˀ5` �v�6D�`c���$8
Ȁ��θ5<l"��5D��x�$"9���q�K'1Z5P�8D��Ҏ��[,�j2@0A  	
�+D������V�Q(�]�R((D�(y$!L�E"�IӢז;#J�a�%D�,�W	GD�$��Gg�=uh�d�P!?D�� 2	�Bc�4G�M`��obXT�r"O�aP��x%�}Y�JI�p�EH"O`EY0�9kn2e�TJķf�H�;"O�`����"GЙ�UJ�4t����"O�X�����Q�$��
��{झ�"OTl3j�(�p@��7�HU	q"O�Q)2��w����.¦Qj0$У"O<@��M��6%vX�u��6_v*=KS"O:)C�D�/�v�Q�Ƕ?t�6 8D��0�m����T�Xj(�;!�7D���Hɤ]��-����dYB1D�L9��@8&|d귏*y����-D�XrD�\�
��D �.7�l�"*D��R�ȍ8n��C!��?t�t�6L2D��i�@oI1r��0z�J�
&D�$�R�ͧ5r0�꧁�8x����!D�К4�,є�;S,�"p�|���,D��!��-�40B�E�m ��6�>D���a��#E6�q�o��\t�AbD�1D�QN���YA�[��%���.D��I6�i�H՘ŲP��"[�?��B�ɿ
RN(�S-0C4����eK�B��#75�<j�˒-��h��C�2̒B�U<aZ�T���4�DR>=.�C䉭�Hy����d���P&�_�,B�I�&��y�gI�uTUi���C䉏�i"�JD�X��ѧ���?�>B�	�4]��񶫚)|��l����t�"B�?���a��;��&O�C�I�*v��kR�ANX�TL��y۠C䉀(��r�OC,�@��B�/�JB��%B�P)�i�3$��3�JB�CB�<@�,�h&�O���Z'��Z�6B�4lO�)�5D��.uR��/�)Q�B�I�mU�\"�a�0+d�)�MV��C��v�^�p���/�,\����j��C�ɟ~�D��"ib�t���éUPvC䉢UQ�(vBƊ^!ƥ	ԫ�eQC�<fIZDA��٘p����L,T��B�I?4p֕�����EN=!�ϒ�F%�B�ɊK'R���#~��㳃�o��B��Y��/m�C�d/c�Vi�`"OP��U��u�I��B�+��`p "Oܵ[���/���)7�P�W̲�h "O|�(&��3`��tJUAa��:�"O��v_-`�z��a�O�P|̰)"O���AX��\PԂ��sؑXw"O�q	���h��99���N�Z�H�"OTxB�E�F8��C#h���be"OP���G*i檅cP@Q�&�6���"O�`��=L�n��p����(s�"O0]�^�����\.Fb\�5��;�y���$lsz�౭�5B�ȓE0�y�拃G�T����99�<��*�,�y¡�>N2�̘�[�aXHM��J��y����k�9��j�1]����C�*�yb�G:j�.e���T��Yc����y�CH�+��2$ؼJNxEp���y���|EP��F,P�z��,:�y"a��a�7N"F���3�y""
3\�$�WM4@f\�C��2�y�B��9�&�*qY9"�|����y��;G��|+FN��,������yB��Վ�9D��h�@@ a��y
� L���h�� ���f��'9�Ty��"O��HAIJ8`��y�ѫ˺]ȼ(�"O~��'ϗ�
S$\Ap
ԪP��Q"O�%���6�� �(�=:���&"O�9���Lm&��k�f�?1J�Y'"O&U����3`�I�%\�z��QJ�'������M�^��E�"�U�K`�A��'0v����`pQeƥ2J,�c�'�Ւ�U.{����cد.��` �'�D9c�ā�?�,a�"�'Z>�0
�'�D=�i �v�~Db����Jq;
�'	H1$D�!�.q�Ӣ�X�~��'�z�q�S9`�vYh��V�x)[�'�j}�(g�L�*�΂� za�'PU6��.ҨR�V90���'u����S������=%�l��
�'�n5��eW�J
�MbUN��/t
8Q�'$@U;E�+]���'�;[^<�'�����']07��r�Ċe�����'AK'�V7��gC9���i�'�.`4Fɗ3���kÇ�tuʙs�'�h�!����f�:sǎ�o88ݒ
�'�p� �5f���X�L\�n9�	�'V�q���;ة����Xt.r
�'�D,�@iD�d-����!�-N��X��'��%aV$�87��x���D�T�6�`�'��D#P�ߪa ����D�c�4h!�'����bO�i�b�a���`�y��'-d��"�+����ą�_��'>��PA,K-:�:h�sׅTĄ���'v�[v*.N}��x���>W~EP�'�%YB�C�q��4����K�^E��'u�}����Ƚ�E+ف/��b�'�>���6/gz)Tk�:)x��*�')��[SJT��\���I+و]
�'������4�d����F+|��	�'/$��ǃH�� a`�ìyBl�(	�'	�u���\w���j�\���y�'
8�aϘx�p0�ե<K���Q�'yF����
���2�.Q�Fm�
�'���h��[�`��$��?s4�*�'���[1O�G2pdQ�d�fp*�'��U��oX]>�)�k�)U��Z�'����w�)P���{��ѕ'�ܐ;
�'&�D�s�0��7M�F��	�' ���CӲbnh*E�V�v����
�'��e�N�fp	d�P�mx��i
�'�^���M�`tF�{�ET�b��u��'j<m����Z	F�s��.�B�8�'?p��2O� ,��<��$��rS�-#�'άĻ�mͶ>ͪ�"(��^�X�	�'[�����	ڽ�AiR9\���	�'�fu{���0l[c�7T6��i�'�6]Z㇆�(�]�2�N/h���'����)X#+].`��� N���'���
�	b:A����Om�y��'ϴ���f�!Y^]C�G%:߀�a�'�N���,J#|3T4�"I�:����'��@F]�j! a�e
��e!
���'�|0�E"����6���W�!��'��Գ�f�dr�y���`�4��'�B���g��Z&�M�u�B�T��|`�'��ѵ+�8P���aE�051��
�'����U�\#4��/_�3���	��� �	#�J5,5�@hM��0i�"OZ1��lF9_�M�ǌ���3�"O�Yy�# !UP��W�Up��4"O�a��_�6(��'
``�̣w"O���GW�J�|]�#�D�#\x˵"O��3!BٕP�Ȓ�nٙIZ�x�S"O�y��+�"x�$��̔(D�h��"O��c$G�}҈��ʈ@5R4�"O�MY�k�*�����jש(����"O� `m�K��=c�(�v	}H�"O�PP56�Tui�I�����r�"O"��ȖHi�Z�HOp��x"O�|ٗ��^�"�Q�B0	��[�"O�A�	D*�M�Pm�/�(�0"O�	*�)S�� ĘRΏ�2Ӿ� �"Obp��IW�W��#�@�i��Pq"O��Z=)�V!���J!k�\�"O^@�W���)��`����>N�� "Of��9� ��#�H�"O��u���
�q�H��J���"O*j��֒v$�T��G�. جiG"O`���$��e��»U�>��"O��QCg�M;>T3��t��!×"O�x��i\#}ބH��ƶAM�DC"Oj�r��@Z�2P�*��a
���"Ofl�רT#}�
e��h�?a���"O�MG
�c22l���'/���"OPᄆ4}CƁJ5N�J��"O��CD
�f�|�� H�|���"O������:0�rpDV�zJ�W"O4���L�4���G5z�L�p"O�V�ޖb�́���F'.!̍��"Olm{��(gh�{ U'm��Q�"O����,`­��,f��у!"OV!�&��Q#�hh�$�I}����"O�ա�a��-QBL:DDN4:n2P��"O��:��<7T�8d��g����$"O�p#5��G�@����*�>IXe"Oz 	�
�6��֊��|�k1"O��!RN	(^u��I�)iS4`�R"O�S$��_��8`h7N�zl�C"O8qB�W�S���G43��aH�"O�	��e�!�b0S�	ks$9�"O  2��ؿBzF�����"<��"O��P�˄8R`�$�Fe=�S"O贃W�"H������-��d!�"O���!/�bl!cFR�w��m��"O�Lc��'_�JӤ]��@#"O�	�ՅٮK@�p��iS(T�s�"OB9Zw��1-���4(��d���e"Oj��`	/�"�S �B	����"OtQRgH@Rz9#�.ۑyhP���"O�L�6ݾs�*���푠?�z��"O��+��2D�P��LE�p�$�K@"O���Q�2A��FnK�X��Hs"O����cɉS��p>�b�:'"OP��S��V�mJ�FxA��"Op0	��B%R1�ܳanM�s����"O�q�V m��q�/\3�ơ8�"O��8�mђ6�B�`�Ϟ$i��,�$"OzI9s	8,Fة���d\e+"O\H���a&n!!w��yLlY"O^�U���0lKI�S4�Qb4"O��Y�,υ'=t�kV(זq�E*DY��$8�4�?�4gӛ�O��@���'V�'f�� �bq$U��V\�E�
){F8 %0,g�=R��ɅP�ٴ�F�~��B*}¦Q�t�ND��d�#L@A�C�"L�	�t�H<S9p�d�)& ��Y�أK�Eچ�8� �y��ђA��?��i��7-�O��K��Y���1��4�~��A�i>� 8@����?i(O:���/��m�F�f
-n#
 ��y�iK�6�%���R��k��I����C����(S�NT�M#%�OF��Q��ͦ1�����q�HC��T�7J:4D�y�4f :
�6D���"P�qj@��=zp��N�#ᒙ�?lґ+pd4��&�\����7��K����qű:LJ�����nc�H����j���'H�`�0;@�+?8Fz<h�4��ɑ�M�d*.}��'#"�x�.�!?�����X3�����	��C�ɊuBȪ7��0R�|�� L��w�i��'��7��`˓� t�ON𰧣��
Or	@k܋D4,����D���ğ,��f���I�x%̐�1I�d��hM:&A��	%�p<2,ȼo�N��FN���<�d�E�]ېt�'iR�iRJ����J��$5XGd�aƬ�7~r܆�I�b����9��G�(��34��2�I��*�����zyB�'��O�O���[畑I�@��6��<G�N��=ړ�ȟ�QJ1/�Kȩ ��OWJ@!dI�M��i�I�s���ٴ�?�����O�Vh����w�e)�$G*�A�s��Or���OP��A�W��$9���w��lZJ�d����RG�<e���a$�&1�Pq���͔	=T�ag(�K�Lq�wm
�H�	���?2F!�Jp�4��'�H��1<����*��٦I2��)ɛH�,���aV,W�n,P7�5 ���?Y���'�B�i�6a��H�M���4���, V���'Cў�S��M��i/�_6��Yx���
;�(�S��삽���U�}~7��O����OL��]
;{�D�O��v��i�o�K.�`�$i �*ծ��lڬ@�'��`����ݴT��SL�4I:}�ϊs�Rl�Ѕ ;��0��Y`�,�;4 �"�M�P�>��zӸE��Nܤ$�4���@��z�J�'� B�������ȗ%���2�I�;�lU��h�b�|����ǆ�2@|5{d. �l0]�T�j��OԜm<�M�L>y�'��޴�ޘ���E�&�n�3č�;���<��I��i��y�i���蠤�=�$���4t������%�I����qܢ�B��5M���S��-B�OU�&'[k�.Q��)I �6�v�<]u��y�)�$�҄)��"W��NSWr��DS���kM�N�4�8�͛�%f4�9aH�֟���4��&�'a�I��$���`���4O���v��]9�X��嵟��������vX���w
ѻR���R�H�y��S��u�*7-6���=t"���&����?7�E	Xh �  ��     {  �  Q  W*  �2  �:  A  mG  �M  T  EZ  �`  �f  m  Qs  �y  �  �  _�  ��  �  '�  t�  ܫ  �  �  D�  ��  ��  ��  	�  �  R�  ��  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p �'��Ih�)§R��L)�'L+��4!`	��}�\��5�d��,�3a�٘1��;�IJ>�(O1�1O���쉌2P
)�`#��4|�u1��'��� p >��F��I��M�$�B>q�a؟��Fˡ��H5L��JEx8T� �ψ��lQ�Q�|�f�j�����"O)QD�Æ[����g��(���^��E{��	]5K�0�����u���ڒ̰�!��f Ɉ1���dV ���(!���H�,�R���s��x�$*|!�D�(D���! �-��-@�D 1�!���3�⤈4�Ԕ-~6 J�I�+!��3�|��EoY�#�p����\V�'$�|�,��p'��e�P�s	n	���p?�4�?!5^�|R�'b��k�H�S�n�<���I�F<Ё�7S�z���g�<9��M�94&��aaO,M+&%r�IRJx�t�!�D�2�h��$��=b���p͔VTHlT�I]����1Ɯ?Ϝx�얺PO���C3\Of���|
� @,��ڢd�e���4#�Hhg"O�0��)_��&�O=Fr0p;3�xT�HO1��p`DA	�E�M����Y��U�O��AK����)T-~t `�Rg�8H�� 	1�'780���d��AI2��B�@�q��7�2���
�M�P���w�>-���0��P�S�iB4H��mf�P��	s�B�F�2Ň78���'��[�n��ȓc�a�ъ	�!v��eB�%�=!�������hr��<?�� ��c�>�yr�U�)$mq�V�GL>0Ç�W��ybEݨb�`�ڡ�S�F��X*2 R��y���n6�h���7����эб�(O���IVk�-��-9U:|`Xҁ�*e"?y%�*�@hKe�]�xd��C��%��C��Z�tE��E�3��db�� sy�C�I�j�\�!�*�7+�ș�s*�4A��C�I�}<�=	7�F�0O΁��,	��꓋p?���-U��3��,۾�q��[�<1����>b��׭بb�`����M�<y����M) Y-?u1�L�t�<�`f��'��D���֨/�H�A�p�<���6��Qa٣�*�0G�B�<!��	dh��N��r� 4g��<q���'"��Ёt�!y��� m�z�<	ΐ/\�eΏ�/����B�r�<)�@����Y%(��n�T��V.�n�<q�#�%���c � ����"��^�<!Q`��l��St�ˊ��Iՠ�Y�<�g �4+I��R��ao.3��S�<�s�_c���ु�:��rG�\N�<A�b�x�l@��6�4Kt`�Q�<��%��0:�2�#Y�i��ٺK�O�<i`�݂t��.�I�H�P�H�<����Q.( R�\0$6HRV�D�<a7P��Ę�B�@7 l@��d�<��$��UJʍ�����q}: XS�\�<)�
@�m&���,��m�@3dLZ�<�QL�N��3Fn��R���!��S�<Iul̐X;���6��4" �X���w�<����`[�����0aM<�*�.r�<1��^�3ʎ�%�/A�d-��y�<�1���Mߞq#R�ha����L]�<!!Ƅ� ��Pa
'{�� )�@�<9P�N5��`���9k4Z|�FK{�<92�	:av��W ٙM�>�{F`�v�<�A��:7���5��,�0�Bg�s�<a��&���b `��r�9t��s�<!r(��e���NBp���A��V�<�����<Szu�ć��c��(�M[N�<���'��g�O%2����b�M�<1NS[�:=�b+�^�lE H�<��ȋZ�J7��o�dPB��B�<QQ� �\a��rg�u�u@R�T�<`mY J�`]�����ް�p�+�L�<yPL����Q�:O�����Hm�<��ٍU*���������mJ$�y�H�Q@��,�4�Ƭ86E@��y�%E�s�l���c�c�������yB��;V�����J^�F	��f��y���E��]@d���j���p7 ��y��͝b��9���	-dQ��{�eQ��y2ۇ�h�����x>90Ve���yBm�}�ڈ�+ԓ4� H6'Ÿ�y
� �!	W���!�Z���hN H�"O�����n^�dN
`$!�"Op�a'�p��hSD.		��aE"O�%Sucb��1, ?z� �"O�H��J�hn �PbX�9	P�c�"O^�e�F0
=��*�,Lt��U"O�Yo;I&�a�+��.�(�v"O�tð!�(R�x���*�@�,��"O�P�f+`�8�襫p��2�"Oڰ���Q��b�I�ta��"O�#!�²:Ƹ��b�?B�e "O|��A��A���rA΁
LT�'"Ot@@�˼
"��Q�ǤHj��I�"O���w��1W�t���/�@Ix�"O�ei@�۶]"�X�-��EǺ)"Od�:3ifm BU	���"O�8��L�3+���
E�S�rV�t+v"O�AzaE@��С��w@� �"O� �M��E��L��;��B�"OD�ޤ����-�)e>�(҄"O���v#�D�}1��	��;�"O�HtK̬d�"=��w`]�"O�}84n@P3��
��%p ���"O�i{F���a:|SFB�4~od,V"O�xhe"�
p�0]���C�AqvAcD"O<�qC�IK��:�϶de��"Oz��B�݆a� �3�L���"O��pd$��`J�	P"M������"O�Z� �u��9�͓o�d� "OxQ���Mm�)��a��v}i!"O�IC5�O�?���ǃH(��A�"O�J�`å]4�X�KR��K"Oj� I�6:+PUXc�A'���q�"O��0�&|by��(ƌ�� ��"Ox��h��6�>�q�Ŧ\�" �"O��b9�(�Ai��Z���U"O�1S�*��h�,gtN�IG"O�u�  \�6�,s�&	 g\`ع�"O�19�׎q=��0"�S��"O�Q�N�VdhAF�]>9H"O�J5�G��6�j���re��"O��@be�%���	�"
��"O�0&e�N�dCN�Eqy 7"O$�#��t�����_�g�p�"OX����'=FA��,9_d���"O�$B@�˰�3� �z�\X �"Oh!@OP�Ѕc4�SH�-��"O��9v(߲M��h�4�
'E&�k�"O>:Rd@�i�=:p�@�L�[$"O:�K扉���� �["ޭ�u"ONX�H�f�����Η�G��-�b"O�q��/�XH�qkA���He�m�b"O�����2���r#�ٿ7RI�"OD� S
]M��	�c��1)�Ԛ�"O�X+!k�sZxt#`%�7l|I�"O��+�mb���v
�N4��"O��21�� �Zݙ��Ăh�Bɱ "O(�Yt� �S�H�Y� �h�"O�A`�=�����G��p�(�8�"O��"�˷j�!2�d�/�Z��c"O����X<jk�`T�B�S�L�)�"O��BWG#�˥���$�f���"O ��S"W˖@���#"� �"O����VX>j�ΙO����"O� J��)X!���7�'_ľP�$"OV��oթ �ra
�EL�0�^8�S"O�hJ��Ѕ�t��a;4��ܺ'"O�	���D34��C����kw|q�"O�1����=3����/B�C_xq��'J��'���'q"�'+�'��'���`�	�,p¢��ʹ��']�'w��'*R�'�r�'���'_Zu�LM�D���@���
�� Z#�'���'�b�'`��'��'���'��Q#G�X�u,��B�Lh�6���':b�'���'X2�'"�'���'N	�ᥟ�q���8���&_Z~�cE�'Y��'���'a��'���'^��'����k�>���ǰ-�1c4�'hB�'�b�'t��'�r�'y��'ft,36���p� p!)T�< ��'\b�'���'}��'�B�'��'R��hQh'�t墦 [�G���0��'���'��'���'���'�B�'�f��c'��q~dzi�
vg�}"�'�2�'j"�'��'�r�'m��'���H�:a.J ���t�XHc�'~2�'[��'��'8b�'���'p:����=.i^	T�J�#*Ή��'�B�'��'�B�'_2�' b�'�Z<��;��
��S�F�����'���'��'}b�'���'��'��x�W�@WP�R6�@�^�f����'���'h"�'��'���`Ӯ���O�@���3g��cFюz�`C%+Sdy��':�)�3?�v�i��9f�P�2-ei)�^-��(����d���i�?��<Y��io �S�CNW�&M�F�J@�1�*b�P�d<��7-<? �^(T�2�;c�1��G(!`1K�Z	Z��_���'[�U��D��IZ�B�Z�jM�<���@���7�T��1O:�?u8�����'�GɂTZ'�עi��%��"T�\|��y����s}��4�N�1���8O����a���۶"η Bn|i�9O�����hS�d� �&��|��/_��� �G8�P������d-��Ǧ�8�i'�:'�(XB��A�*��%@���c�V��?Q�]�XIݴ<T��1O��hg�mѱ<{L�#���s��@�'S���B�zZ��T��4|�B���;E��N���b�4<����/�}y�V���)��<)���+>uB��ۻ#p-��O��<ف�iXrqi�O0�l�N��|bg0NO����Eȹ'<�A���<��iz�6M�Op���~� �8��r�Ν/5vT ��i8peHǫ�r�tpD26�Q�tQ���ގ�q��'�@�[�✘P9ՠ���#��e!
�'�p�J��<�, ��M��a�@LV�rCPA���]�d1����L�J���.�`���H	����OQ�n(�ݫ�אJ���H��9$hB�ӢՒ݈�&�4f�|8{c��+@}j��܆2^���WJ��-2t��æԬ�u�wǖ�[��Œ�,ޠh��U�&�
B�%Y���D���޴�?Q��?���^����&f*����W]mQ�����7��O:���x�R�d7�4�^�O�ZI;�R������ʔ��=Cڴ��B$�i�"�'�R�Op"O����)c}:`��F=$����6��<n�(|c���IE�)§�?�5 ��#���r���X�wB�"?��6�']��'�\�d�1�D�O��Ĳ���e�Ңg�"~�6�(�2:�������I�{����'�b�'���O�)�e�MSj9rq�>�4@p�i�rcC�O剀����O�s����X?^��`f�*<��͊Ѣ?����;�ң�����ϟ,����{����AӄInD2�53\H�+F���O����O�3���O������HS$y
�� ��d�v�r`��%p����h�Iʟl�	����mRnZg*�	P��90I8?&��HU馕��㟤��`�㟠��]�HU�B!k�`Y3��3�<Q�������_���I��D����u�����̟��ɛA�&�x���'���X�GK�`|B�4�?9J>����?��Q�b4 �&�p�B��C}nA�5���2\<��oӦ��O˓v�-aњ���'Y�D͕�5���!r#�=9x48"��n��O��d�O���d�~�c�ٲn �T�"�ނ}�5sgDM��=��ݟ��._���������?���П�3c�ҡq�Ɓ?RT�#7�`6�6-�O����\������)�g?���QF��a���rS	U�1��+�X(��'k��?�������'�~숢D��,��e� �syə��bӊ�:�FN�$@1O>��]�F�%��'1��1�C�6LFNM)ٴ�?���?1fh����D�|:���~"Mee�1��שz Fh��ś;*���yR�Ϳ$���8��O��� r�%�%�U-{"&�B�����o����4nƺ�ē�?������sR'� X�g$W.{�,�s�㦑�ɲUTZЖ'���'��Y��I���#2�2��⇦�C�d�Ҳo�|y�[�L�)���Hj龩�ǐ*<�~ ��Y��4AD���	������'*����i>Ip#J��6G:��K�(!;��s��>!��?�����O��J�m@�(J���3�䁾/�:	U����$s�x�׵=20d���>u,�zQf���O̐K�#�_�� �D�E,e1�(��'@�ɘB,]��%��	_���Y�'�X$�4�̬j�\КLO�'�F��G�C��J�K�S�c�B�%��+�섓��C���S�찹�l������B��%nx��VM ����닍&�"- ��g�\�xPi	h�? l���Lz< T�b�^�i2nA�Ue��Z���Ď��>U3E$:d/��Z�f NU]�s��O����O��q�� ��PK0*Y�d���ؗO�w8qxsM���X�+5Tџʧ���?�ǥT.c����ƍ�������9y�1S��]�s���~����'`8hU�ܵ����d���/����@ƃV�b�h��m�dD��Q�*�BE��xR�"�I���Γ�?Q	�Z��ɥ"X3��]	���,:�����HO|�	�O���!���r5r��0�
=����,�O��$K'NTju8a��O����O��$CȺ���?с"�v�9ӗ�R�+;zX3�#T�<Q��+Kehaz᥇���<q�˔�G��gLT)"����%�E��I��)a���!�R#h*X8�'v�Q�����%SЮ����/�>�Q%(B�p"����		�M�gy��'�ɍ�йz���9���d��ǼC�	ߟ{c�KP��4���S�&������M��i�ɧ�	�<a��͘Dn�f���M���ggW2O�v0X�Ϻ(/��'��'����2�'`2�'�ش�A�еOҠ(0f�i�$��d�\�LVbq�e,ʕj�V��w7M�y�Q�@�k��L�+�/\D��"E��W�]:�L�= #}���b*>�3�f�?w���?����Οl�޴\�\�󣏗�v�yaT�G�T��
�i{B^��	h�S���X�6���b1*G.�F�3c'J��y��+_~`y#�6.d��ek���y�jr���$�<AUE�f����'"Z>���E�;�ؑ`�A�ZX��4��r.��Iʟ��	�j���$�څ	�01�'��>Kk�a�Yl@�2�߭��<�-��|^5��U�V2�L#1/Q1*���Ӝ
E�q�����1
`�XP(�<��B��� ߴ+���'z�S��������f�Vܑr�������U�S��y��5���Ql�^^�A+% �0=I��P�&�nӺ��]���eA�8�Bp�"�B"r��O�t`$mZʟ|�Iw�	\.R�'����}N��4���B��9�b��=(D��B�2~��x�(�
�y�S>I'?牵Rkz��T!x�غ!�S,�X��˷@ڑ��J�(��{�
�.f��ʐ������,?�ĥ�`L��&�ʁ �R��I;�Mk�Q��i�?&>��S�1��h� R�{�4�;T�;d�$�OD�=���F�N+$���D#>$t�@��O$m��MK��d+���'���O�=``L^	0ujA�r��JhL���'���K���t�''b�'���c�m��ʟ$�E-P�r�f��TT��Z!K����Ǎ�=N|��ɵ9�@�`eS�>Ӓ� �-&ڠ�I��%�� UM؞(��\-3�V�Wʙ�mδ�'��"�o���I���<�����L�U(���#(kd��#�ċ3*!�$m#\R�N���N ��3O�FX��4��$�<�e�1���LN�:6b���GǇ'�@t�Gz�2�'9r�'�`�'�'�5�|�b�gɝJ��X�"��!8�
�����8�s���qg�`�+��5���#�(Od�c��݆G�M��Z~%�$X7�P3O���^	����T��Oč��
�OpE)�(6��Ot2v�N0$o�VQ�P��+�����"OB9����{7Js'��=p�`M��''ў$Q�.�W���K4��G��cs%u��ڴ��`f�<jU?]�	p�����:��_�sT�,��M�1Nmd����'B�'ɲ�r'������0AV�:�Z>=R� .I1",�1@�&s肕��1ʓq�3
�5z����搮X�n�O�z��� �˪T���Á+�n�Ȏ�ƌl�Rhxӂ\�~�7$�N�����E�ʄٷh�<Y����>9�bJtn�z��E�8�:d�T��x�8�H<a4��\�@k ��,5�a*��@�<9��~���'��Z>�2�՟(�	��0����,s��&��5��a���X�q�1�ِ\���: ��v�.q�O;1����6?��lac(܊~�h�J �B��b@�Ǟ���Eg�V���#���'e"9�Fh[��p0�ƁF<�1Sf�h
2�a���lZޟ�E��
�RU����0�����HR�5b>̓�?��{��r�D����!q�$	9��Ne�'x�"=��'�?1�̈*l���b�F��T=+�'
�?�� j�h{f����?���?���	��SƟУ��5��*��ٖ_�$��� ��D�*�r	24�F�^Ԡ:Dҟ�أ4X���'���ㄞr�L���Q3t1��c��Ƕ9X4�9�( /(2ezf��"��Dg�!~h������+"�I�zc ��䉃��d��&(tmݛ�'o$}�P�'Y2��,O��ģ<�F�P
�������r`�T��u<��_��9�#�0[�b9`aE��A��x
����?��IpybKn��7��0v�e��N@� j�#E)�"=���D�O��d�O�� 1��ON�$d>Z�ϒ�%�*��G�l�(ç�إZS��*Iݡbr�\-3`�YZǓ}*�:�����=�����@� �N
L����Ō�i���*�/8O>=K��'�7-�90lšc��4Kx�3�& �O�b�l�m��T8�>�I(@����Gn<zz���K��B��ɪͫW�ö5 �p�(ԅ-���	��D(�B�π >�L�c�� Y ��|���"OHLR`�� � ��08x�"ORԁ1��1Q�����KN)J�P�"Ob��U*�qڐF��@�"O
i$ �,]Tf�#m�1�V\9�"Oʬ�2�YQ���L!k7�y4"O��Ss���#bh��խA�1T{�"O�ؠ0M���z��E홣EF��C"O���mH��X�'^:m����"O�i�3�vazU-�  %B�"O���-P�k��=��f�3�l "O�z��ғZ�}�6�	�&MT"O4���R51w�i���Ǐ?� ���"O��"�B�\M;Ģ�	M��YE"OPX2�n�U�qk�h�F7F<�"OR$#W,[�Hy��٥g���Rq"O����ģz68M���ެ?�^!:�"O�8㇉��P��c�C�V�i�p"Oؐ���V���$A�!�/z�ҥ�"OH�q�M�]��I+cay^��"O~L����7�N-�#� >PT�H)�"OHb�V�.<E�%��w7(I�E"O|�g,x��}KA�P�\���"OpIc�ߟZ�-��M�4p����"O.��(hZ.qĪ·N�J��"OXcP돓}�hUY��ͪ<�`�"O��L�;>$�t�T��bv�y4"Ohhh�oS=!"=����&L����"O��c#��>8��;7o�n�n�pF"OZ�C7��5G:ɈЎT�4}�e��"O����!��p�V
�٢"O��J�*�X�ʸag.�(�����'f�`䩌~���H�ⓏNa����fC�дx� ܅g\>��ē5?*���쌑�����?{�U�>����ՋB���3��DSܧ�։��)v
�btM��I@B	�ȓBaʥ�@"\�����e�+�L�:` �S$�U�P��D�P���$:���6��-a�.���J	k,!��3����p��	Afh2@.V�&J�<���&)�,�(����']LK��ה�$+��=��1
�!��"��B���:�Ү8˸�k$�*Xy8�`AX�t� ��'X�iBע �L!���ָ(�����}2&i-n`��M�B4
a2��)�Nd4���ux�
d����!�$��)Ȥ���5h�ɡ6�Y�i�R集D
�[���<�?�2�>a5@M.A6���%�\���g�<������嫃����[g���5��	��9|tr	21kL��I A��ǀ�w~�y��J���?�sƋ>C��H���U�>�(��P0<|
#�Š�H��
�_Z,Aï $�!J�Ϝ�y@���Z�3!�>y�L�#j��j�B�)qЈ��o�i?�}:�
?Zٸ���a];8�޽�M�<-\���' ,te��M�r�>�/H���/9@���L����td��=}�cD�iZ8�r�*i�Pa����?�eeרTSv�w16	f��1$[� �:��i�0��a�hVXò4ġ���p<�RA�6��lq�똓O���+�C�ey��ɏ#�>h�֧D.)�UR���(O������\��t��
L�^��S�i����rXc��ȋv��Dq���j�f�2ЯʘF�6�RƌݝR30Y��c
C}��G}BbCL�I z�9h�R�v�H#VH�6]��3i����{�	h�%�Ӈ8>,s�e!Ou�$��$�����O��	&P���#0ˑ'Zvd��j�/�u-��O<а�(��H|��@��+(ٛ�i&��G��J�,��#�џ���+c�!�ɖh^��Д}�U0aI�=q�m����zeûb���4WQ�#��>�$l�(�����`<�L<���MQ�'�D��A%�?�HG�K.|`�xK^�B��#������ǱpD�F}����.A��GA��ᙗO�}L@���R0D:|��D���?a�@�)��T�f���l�4<03BK��,�Ā5|O��c�D�7 ���-�8a�5 Tf�B6��D~��D��	Ѩ	�S���;P
�� T`�W�Az<�7�P�,�����ɟ"����g聜i�eSS����7MJ�F�J�f�� ���S��3�I��\�	�?h�$�L1�$[7�M�P�(��	n?	EO� ~9����&��u�`� w}�`�)��5�a��$������^0�HOJ	Kvj��!tHE!��zl0�㧜�D'��F�DqB������X�JI����=;Z�<��iֳ����Q�ܐ(2*ܱ�m�3Nf<�뉜*7libF���<�� �RtE��lZ($�-bV�3|O��`D��W����o�"]=���a�Sf�D~�a�4^+���C��͢#ʄ�Y�\��X'� �"wLd��#.G���xF~���d����	>1�
d"�̃��M&��2M�R�ȊM�\<��JD}���
f$h[���(v"�h	�f��c`M����aq�O�i�䎘+^&B`L:\!��^��0
8 rАB��6w�dpC�%�n>�� o%Z�i0*؏3�¹��om,��A�F!C���	��T�.����D�A�<(��V�\�$A3Vf;T�4�0	ߣ�l�E}"CT�	!O����t\6P�$�ǫb��@�P	=�{"N~�%Iň݆5��Iw
]�-l Y�)�	$c����6d�R0`#@�&���ra�M�(��<�®��O4Ⱥ��+S�:Ds�56-	$�i��Iޔ:�H�`	�`����*FP�'�VN=	�P1�K��r���9��m��.�Aq�7�'XV�0ե&��b4$S.)F�e����4B����a���Ty���K.�F0O,1���
c�v\�f��+��OS�=A��D;!㛷��峤Y��"/�)Y_�̢�$���󅮟�>Q#�H�!��
�(��5&eC(0D�4�"��9$2�����R�$ ʓh_�m���G*��~"	A�{�O�p�(Q�>����dB�y���gV�M���O]؟���Jg�<Q@�b�4"��h��[-H :�K��%T�6M!�!��F,�Ԁ ��[8���"b�X��A�2x���ZWE,�<�xaab�{J����cM5qif �C*ٌ2
�gΔ3�Z9�&��#$�B�JE������#�H�WƘ,/LB�I|b� a�
8iVL1��DnB�I�e���x� Å"�p��M_�HC�IPq����m�������B�I�w�r�P�FP8W#N͚�iY)Y�C�I�<�؄(��, �=����6s��C�I�/F� ���-q3�QC�I܉K��C�	�'��p�ӊ۠�89aM0,�C�IG�.Y�􉞳:NX �ƂS�x�C�������|�2x�է#_<C��F B�ڑĕ[� �Ҳ�Q*2#pB�}���7�]2H���
B��jWR}������q5�K�?� B�ɦ�՚g��;,��1�&�H$2	�B䉍AJ�F��E<=�d'ҩ'��B�IL!�|@�	� �2��n�"k�B�I�'z�+�b�p��5Z��C��'!ú�zWNӃz��\C&F�h;�C䉥Ҧ�(P�� (�d��ٳ]�C䉳E��A��M2���#�K�[��C䉇he2�(�*��P��t��m����C��+�ƌY����{�iB`��x��B��o�>���C��aف�>�B�Is�	�d���:�J���5��B䉬{F,���C�h�P��2�7nq`B�Ƀf� :e.:x8j�`�w��C�	�w�P��t�6a�<ݓ�韼<�C�I�~�~i���ùF)�Q��nݮm3�C��Jμ������y+���)h��C��9/�|(1�O�<���p��".SNB䉊M@a�Tϙ4RHZ�p鑵/�B���P� ���[�{�o��h@B�I/�XpqGW>TЖ�yc͗fJ�B�8T~�I�`&li�跎2�2B�I)\�l��V�V�h�� ��1T�B䉵#� �Q`ޕ#�` ��
���C�!��P�Ԉ*gҌ��K #�C�I$<�|���	��w)L�*I��'\�е�� �cS�84~�C��� 
̻D�?�Q$��2@͊A9B"O�mB�O�`20JA�O��dB�"O`�������+�)�6&e�"O������3B&
��C�f�"O��5�D�sHd;��۾^)��"O�J-�3�r\��//Cp�"O1�c�-��L�����	��"O��P`Щ�,�����v��0 "OP� #��!2"PaYt,�6t��9��"O�lA���GB.��J����"O�,i���%ar�!�$/�r9�r"O���Ɨ?��(peT *�:�٥"O�0`�B�
��H8`��<�R0xG"OV}�F$̆*0.�0�O��&��|R�"O�y3��%���E�;���"O����ڶ}c�l�@BX�u�
�h�"Ov9���J�m�l0B���S�E C"O ���"ޣl��!��D�5&�֐� "O�C�K�2k������Z,PXP"Ot�a�|��y�'�>�TP"O�����ێ�,�XRfG�D��6"O��r��|��Ãg �#�
ȓ�"O*2��Q:�:�z�`Ϗ
��"ORp;�	¼Ö݁��B� ʠ�3"O�� 4N��f�E�AiN��t4��"O$l�SM���EaQU�)���"OZg�̿B�(x�Q�۱z.����"O��ɲ�Q�0L�C`�c����"OR�����
�F�F/tPhS"O$P�h�>*0�d%C�D���!"O��c�LݛC����T$O 49:pP"O$��h"<<%)D��X-Je"O����L˅,'��	�B_�Y�n�x�"OF�2���e��!����nA�"O.����"R ����5sN<��"O�X��+�p�<T@`��J[��z�"O�Գ@h�@܈ �G�^����"O��1ᜧU/���$l%,Q�`w�<q��y�D�J��@q���]�<�ש��+pD����Y&6&��� T�<����>e��1����/�(��-�W�<q��ʈu���#@;��*�IGV�<�7�F,0A������:`��)r�nJz�<�scA�
P�̪�O�6�^���v�<QP �q�X��f�� Sup�-Ws�<9�NEK"T#'�_V`) u��p�<��È3+g^xH�Δ;��A�Ak�R�<��埫�^@��.�F�� �w+XY�<QtjK6\&�5iG7]���d}�<!ӌ�[����,<i��iCa�z�<�V�>'���-�8&�h��tm�j�<�E$��)��y�M�5X�q�EFN�<!D����;tj��h�c�ZG�<��-V��Q��AbF�HS�+N~�<I��[>u���*C�_��dj�e�<��ĉ9!m<��Q��,q�N�3�+y�<��(;�|<��B-^� ۃ�v�<��d�2MA�� ���")�d�
2�	t�<yf�.
�YB����\$��C�u�<�$�ѭ@���� hǢ-xP�Kq�<Y�ЫM"h�J�9n+��SORR�<�Qϸj�R��p)�2�<��d�_P�<���) uq_5�����	QM�<��jԚsL8��ڹA-P����d�<� >�@���q@r5#�������"Otţ�0l�ʢ�:_���S"OV�@��f��c		S�8�"O�J�#�!�����Jkrl�`"O�z��]?��(���$4�t�q"ONx�� (yy�mS�Dʬ#!"OL���%W,:w���v猾p�5��"O���A&T�#���J$��|�VȪQ"O���gm����Dbt�^Ֆ�a"Of8;�@S�x�&�ǁ�
�Z8�d"O|	��L�n�$�f�s�~/�y���6(�:���Y�_JҴD���y�̎�,(�T�!��o-ܭ�3k���yr�!:�R
O�<)�E2�l�:�y�@�D�E��L^�Ky�iI��
�y���*}|�Xá�"BRm�b���yBl�(r�uy���1+ q:�M�-�ybLU�o�T�;��"9i>��e��y��i��Aqt���1�����8�yRF:=�X���G��3$�Y�n	��yrJ֋&�:�Ӷb2��@D�(�y�/½1�Hs $�/[<A�g)���y�XR��]��n�]�=�Ȱ�y��Cp�@1dl��T���h�!�'�y2m�(D\�p O�F��1�%�$�y�f@��,c@�G�B/ʴ���Զ�y�ߠF�"AP�ֹ:�pA:5��'�y*���$jf��66�H���yG.�k뀕.Z%�d��y2�%U�X��6� t���Y��yB��:� ����ǣDb|�a�D4�y��GI��$x4LW?3�x��� ?�y���%V�pc�I�&4P8b F��y.�lVa@�Ê:m���4�y���w����aQ�Y̢�[�d��y���@3np[&e� GB������y��V?��U��K6cB���.W�y2�JhR���Ei� 	�~ȹUj*�p<��$�
n��YeANm]�����Wb!��ӏ%U:|��(\> m
�@��ً[N�R���<E�TE��Ռ�w(Ρy��}���&2!�ċ,d�������aB>Y��/�O4P�͇FzL]"��H9F�Y��"O�H��W�1�R�h�O.��[�"Oѓ�	��C�rEJ�Iİ1��9��"O�`
�84q����G8֮��"O
��&��(IQ�,�7�D�<�D<
�"O�=2�<Ly����	�\-����"OR��嫉d�4X��-�x�Z�"O�$d=���bpF[Aς�r�"O��h��X&>���f'��p�",	�"O:�c�'W�z��E:��R&���ZT"On(9R�Q�Zp�D"RnԙU�H�R�"OD`���A	u��is7�/U���"O���4��m�5��F xX� �"O��5"*z��`��O�@�4�����IH<���eL��c1OL�l@�|�Z^�<��a�?tN�#i˲l�x����\�<I�*�?�TX�#C42��P���T�<�U��:)�S2z�*��f�<Y4F]�a1D1\1��q��a�<��یp݂�S�m��C
���V�<I�e�|8.�sk��)BD���+Uy��'�f)��Ò�DuB��5���
��� ������:S
�"JT��D]��"OHta�΂p-$��<<'�����Ic���IS#"��B�OӒ?�X�&�%�!��߸!ݰJsa��E3��²��A��$�S�Oa�zi��wQ�lT{�lt�'ˈ�� �սkC,��I>=�	
O>�A�'^,A*L.�T��;$�p3�'0�ʕ���I/c���A�;�y�,��N�Րq���py
0.]��y���?7�R!3�W~�-�r��2�y��~2aC�KK$�-�S��y��D1Lu��K�.Y�s)ռ�yr�̋(�4�15G�
C�S��_�yү94��%��NN�k����fݍ�yr�Z%*_ 5ڑH�2\|���%�1�y���/O"zx�Q팧Lg>�s�����yb`�b�Fِ,�(P.��#g����yT�J��H���_X�i��C��yb�ѵ�^�(`���X����K9�yL��2t�p��"ߘ��Cԧ�9�y�f�2\�j	�կ��Ԥ#TG[��yb�ۍU>�%��N�t�l�F(���yr
��p7���aLf�4���@��yb�m�ި���N�Uz��@�I��y����u��įB"��`d-�y�ؗi�����N�2	�40�W.
��y��T�J�L֤׳
��c�/�y����٨҂��4�̝�7o��yBj� :���`\�0������!�y� �C�⥃��K)WR��#�6�y�k�Q�؀ʤK�=A�O�yB�̸v�U�����b��\�y2 Q
]����%WE���e����yr"�h��-��H��ǀȁ�yB��3l���-�J#����ˎ�y���p�ȗ�(��:
���yhU"��M��
D�p�,(�����yb搖>�HI�Q*@	R���k�)�'�y��Q�)��H�#ں���g,���y�����=S"�M�bTH�R���'fD� P�	�W��-��@?8� ��'���f�9^x ����3H���	�'��`��V	j��1�cB>���P�'���UTk�<*@�;L{8�'\p������9�ř&$B�^��'c� x���Vp���#(���;�'�K�� uEL`��Q�p�V@�'����Я�5YXt��rIW86L�5��'���S���qɎ��E�$Fҽ��'���!R`4��t��dT&*O��
�'�"I��G��tY�d�9vÄ��	�'�^��b@�9g;�f/�'b+,���'fN�� i�(����K�?T��'~� S�H
)�H�`�Sl���'c����Z���H�uj���'�����޷6o�Uʋ�DrܨK�'.$L��.³?�V��di��D��U��'x�Ȁ� ��[ �9CW�U�jC�Dy�'�o���m���H�HV��"O��e��5
`���H�C#��"OL�S� �D�=���G>�"O�a"4���X���"��)d"O`#a	�g�^q 5��m����"O�=r��j�F%���E✩�"O� �)�6��o��6J�?�L��@"O�uj%hG6;r�XãN�}��,�"O������0�е3���CJ�c"O���œ<=�9g��(){���"O��a�-_�pcB]�=�"O~���&�'WSDa�Nڞ9��HA�"Oh�A%��7�ɨPm%g�L�[2"OTt��%��b�H��lT�rlf��7"O�U3���+N}�����QW4 ђ"O��C�BF��(([�@Y�o@
�"OIa���BtL�vb���m� "O����G��_"��%�Y.��rC"O.�PT���qˀ጗sxY`�"O���M�81^���,inސC�"O���w�CY��8�0oXZ%��"O���SM�e�:� ���A%~̱�"O�T{�N�
PP���0-�T(�"O��Q��þz*���#�)3�l���"O�|�@"�AS��iԤ�)�T�I�"O|pG�G���)r힠:�j��"On}��DهA�����P2d��F"O�
�b��"����f�M
�8""O8��J�pb`3q ��*2��"O>$�L�7	U��鷠�W��ۄ"OHD���	�q��"3�K�qi����"O���A ��b�+W�QM�u�f"O^�i@�(r1��Aա��6=����"O@U�A��K{���  ̙a+��Hv"O�h�JO>$|m"5o�+y&4��c"O�͒U.���,�[��Sp����"Oj�@�'�^��+Ǝ�v,��"OV�IT�J��j bs�̖�4D��"O>�acI�=����7)[�c� �w"OF��Gʿi��Y��IP}E�`"O��h��1mβ�X��0 ��U��"O��*��ˣoN�����E9D��M�"O �1X�$��hP�d�a��N7�!��ǐ7��E��)X3{z�E.B37�!����>4��	x[���8h�!�d��$���kdoŤ@̝���!��D�"��eB�o���#�e���!�䄵]wI��R�h�v�c�$�<P�!�$�[��Ź�Z[�ڑ�Y�9+!�d��4�r�s�N�j�@���W� !�ĎC�!�G)���ι'  c!�䌅����q<#�\����X!�dUd�i{0��
Hj�����I!�$B76���k���p-�mq��QG!�����1PLS)cE�c��Ş�!�Ĕ	\�0��Ĩ��J�8K��Ůi�!�d~��h)R��7P��sW���!�x:��צ��&x:�t�I�!�[�$͸|*E"F4]t,�5MS�!��npD��ӈ�uh����>0�!����&斕Sؕ�� �
�!��
L��ç>hL	�%��p�!�Ą x�x����OJJ�<r�!��T�}�&�<Gb�| ��a!�dͪ4jи��KE�ޤ����p�!��v$�<�f��(�b���Y�Z�!��-��� ��6�:��RI۵Yy!��B�� ���	<�U�J	!�D/m���P����LPGK 
!�$ى9�ZP �.��1�����!�� <�ӄW&dw&�
�a�$�=Hc"O��x�ߣ5PU��`S�pn*�
�"O�;�2p�t� '��M��=��"Ov8�AI_� �@�9��H
��%��"O��iE�3|hn�a`Q5c��$�3"On	�E&�6dx@�/Ky�R��"OJ4�f�\�wඥ���
�??!"O���A--"����*q^Nx A"O�q��.�-t	�akc�CT�Ty`"O�|���K�,h�5��K�3[Ar��"O�h[vQ!S,M(t�Hp6:%"O�qp�O�?W5є��]8��"O�x�PiH/��)MN�p�"O��J��@��I��gٻ&ڎ�#�"O���Ux�0��LHA'"Opq:#�[?C�|��&D�"$�n9�"Oz	�O� L7Dq�T�a޴�U"OX\Xe��l�'T���#B�0	�!��#^(��N��Q��Ԫ�Am�!��23�q32@޽h���@v�$�!�dP�6�0��0_�!@i�!�$	4x	�6oHD�ey��
�LW!�dZ!5�����\�r���&Ո$v!�D�.�@�C��F��'��s!�$T%%����t�B�/��!Q��:9�!�D�?I@FP 7�Y�G�,D{FK��!򄕳f�Љ(B+H3W�ʐs�>���h��e� TJ��� ՗n`܄��t��5Xrf��Uy&��v�ý ��ͅȓ>jD�b��K%I��𡑥�:;L��x
�ȷE�$LS\����U�>WI�ȓDք\Z���x�~]�`(�4bņ�~�D5��� �e���Q�&x�ȓK�6��'����t��fWn�z%�ȓkޔa�iʆck���O͘ȅ�������T�L�B��&O�W(ZɅȓ8��+�_�Y���pS�O�v; �ȓ*4l��kI�:w6ѵ健@](�ȓ٢�Ȅ�(�@�,F?ƕ��"d
�I
A"l�V�G$*O(�ȓYG�8�lJ3�t}��`ȋegdm�ȓP�N� -��$� �;`M�`+�ȓc�T�0'<v5𽐂�W�\��ԅȓr����$*DHP��VK>��ȓRJ(ф��B3�@�@#�?a�~h�ȓ;�� ��oW{�������5.�q�ȓL5�M���E(�9����6̆�$oȤ�c�K�i��\���&�y�ȓe�ݡWh�s�}����Z��x��C.;V,���B [����zSBj�(�`�б�T�YB� ͇�	ԈӖ'+<�d�jČt1��ȓhҵm�sH�K��|�.y�ȓ�&ܰ��H�3bt[��X	�l)�ȓ`��r�〢 �^��VgI.O�nL�ȓ`i���VFK�L{8	�K�'tav����8��v-�k�=!��'��p�ʓ^$�h:⦜>*鶯	ZC�I7
��%��(�W�p<C�	�K��y�C�ڼQ( ��gA:]��C�I�
�R(�c��"(�Bp��2��C䉾[<��NI�K�Tl`�H~v6C䉙X5����䀤PF`S�-c�ZC䉽"��0rIH�8�(95͗�{�dC�)� r4�b�F]\-{q`������"O��:�Q�K�0�Ap�;�~��"O���P��d�᱂�1W��;@"O.�pę8Q�����^�)L��7"O �pQ�U?(.� ��F��#c"O*��Ԁ�8At�9@g�&S@2A#A"OΥ�ū�
�
��X�)7���"O�ܛBJ�C@=x��ɉo���"O����P�v��R��U�gR$yb"O8l��L����'hGd�"OZ����*A��(h�@+5Da1�"Oj����U�1��<*�ߠT�.Q��"O�<��MR��a���U?WJ���"Ob� ���JL��s����pK���""O��k���@{�m�3LJY0�i"O�Ms��;(mqb�-Y��:�"OhU!�+�?"�x�r7G���Qr�"O��Q'�C\\`��ER
	}B!��"O���� =��Q��	ry�pS"O*P��V�eI�p�ůθԳS"O8[v��=bn��k��8bߞ��T"O
���kL!hHS$"�� !���"OJq"a%d���VΑ8I
��r�"OVevτ�dz|�$N[6eeHT"O�H�7L�0B�����E�Q��e1*Ov!�-�jW�Iȅ�(u��	�'D2�jD�Gd^`�Ŕ0X�~|��'�,@Ѩ�%l�rlU�N��) �'�d�rqa����+A�.$��'���H/l-����j\&g�z��'��u�!�ʃ)}(��"#�g�d(�'&��D'��~s�b�]%T��	�'0��3�A�F�0�q�E�Y`,�B
�'S mx��Sxj����ܷMZ�D�'nlP!�D��aB���S���A
�'��]{�N�wRE�D$�.MXHe�'*^�� A$)`m��O�>����
�'x�5���)����gH6(��h
�' j��cM� �Ɓ�wDX!0d$b�'�f��`BK�wp�'�N�,�P�i�'7D�Aኚ 4H@�W	[�ONL�'iytdK�!����R!#� �q�'גpA��Y97��R#'�Y�%��'D��tO���� � 	4��D��'a	A%� }�� l��{~�1�'E�-Y�x�9a�l6�
e V�<�PƁ"���aX�H��	Tm}�<)��Wo�x���|Z*E��F@{�<�Cc>�S�B�#n�rb��]�<���f�-QQ�K�k� Q!c�<�4�R�e(h��bW1PO>dR��XY�<��0{|�E�B[5+.�y��oW�<�Ua�
OrHbF ��M��pb�}�<��R@>ju(u��,r�°��a�<Q��	�������sʒ����_�<��k��K��%���C�9�f�5�ZC�<��X�=U�9T�W%V�E9VB�I�<�#��!Քe�ŭ��<��s&�Z�<�aȡ+�$1h̚?�(�*C��W�<��J2
}>� ʞziB���*D��!A��90ܘ��v�-��*�&D� XR�C0@�w��!�@��?D�0�`��Sݾ1��V�u��yj6�=D��S��L=hҌm@�M�5t&��c�;D�� `d	AA�1)�f�[sb�W��٪�"OTY�����U�"��(v��L+�"O�5� | ���IC<}�$�"O0x����+~��IhS��3��T��"O�M��%��;����E�
� ,2B"O�04&Y7*��|z�	�y'�q�"O�Ёu�5�D�1)O0m�XQ`"O*`Y%V8Y�p����< ft��#"O�p�U��'��Tc�	ϝ",:��"O(-���<mj1gnF���0"O�5���ڟ� ��.G`��$"O�Q����@�Z��"ݟUC@dZT"O��[D���H\c��ǧz#D<�P"O�(U��|�� �K5*LQ�g"OR��D
h"^-�5BA31��Y�"O&HjA���p��F��-<�Ta�"OTQB�[?�ո�O�F�k3"O�Yq��f4�h�!N�"4��0;"ON	����f�,�B�C�F�Ie"Op�ʕ(D-���4�E�!o�8�b"O���ₙ6�4a`暟d��y!E"O2��VH���0$dV2�(p�"O��p��&]`h���G<�h�"O�iR2`A�^ƨ,���>�}�V"OЍ�f]+7�0E	��R�(D��"O���DBF�\u]K^����G"O
�*�OО#`�	Z�@�MАp�"O��"�$�NjKd��P�6с�"O�)�㍌86�f1g�G�ls��y�"O�]97"�{ò�P���MFڔP�"O�5��cӦ�l hu�D#MF����"OD�b�
�"��0��$3��+�"O��8�Ϛ?��1���O}V��B"O:i2c�4�����W�geE�""O�� W��3C��z��?Y`�"OE�� G=heb����zX��!�"O>T��/��1Z�LKJP�W] 4�'"O�a�H�l�qI�	طf���"O���ܺG\:4s�	�6|�"Or`��)͛JT�J�K���"Oz IF��'�tT(��@Tt�M�G"Ob8bԭ?� ��)�L�N�j�"O~�rW���b�*Yr�HA!M��#g"O|� �d<pXل�7c*��ZG"OB�⡉߂d�ʈ�@jX�G��"O�Xs�n�@b�Ij�O%\�a
7"O�d���+�5���$�L�E"O>$*�聁 �PP��mE v��8�"O%�aˬY�V�ȇ'��b�҃"O�Й��G�'��i1G�9GJB`S"O�����Y�	r���k�G�L�"O�J3�M��`p��)�� [�"O��e�8�R1��'
�'z|+�"O*�q���!U�FǃtAZ�A�"O�����6j�!ӀT"X
��;u"O�30�د=������#�(MYE"O��Ġ��*���0��{���7"O��E�G>4"tS#ŕe.��"O�4`��[@���
�mںN��G"O��Hp�:SU,@�f�Z^�c2"O�p:˄:E~��H���0+�>$#�"O���C�R0�ܚb�H���)[�"O�$d �N���􃏈p����"O���d͂�Ҝ�7��oy����"O� 
Ի��ݖ�\����StRԢq"Or�����z��i9L9,]ܠi"O���E�&��y�%+�H ��K�"Ola�g�̃0 �l��O9y��"O�eSTA��Q)(���mF�[e"O�Ex��te� q�+�O�*�"O��	$�ׂXkQx�+N��297"OBh�r� v�N)(3�:� �ڧ"O��k�
�`P��"o�A��"Ob`3��1ˆ8Ѓ =/4�H"O*�+6/�"�F����ǌ)tu)�"O�����:o|�1íH��a��"O����.Q=T5���%X��"O���c�Ȗ"�Y{Ƙ�tƽ��"O�I0�N�B��H�ð4l�)s6"O01a � $���a6aL h �"O���l_L,��#�/E+F�-�3"O�%��k�1�0Q��4}Q0�i6"O��m� �HDP�A�"�:)�"O�I����l�xI��L].hނ��"O��2'(��
b$�Q -Žp�f]�U"O�%h�@LB�����̥_�(�3�"O��Ar���-
B@V�Z��P"O"�A�������$Έ5�5"O����C4z;6��fK�Al$y#�"O�(��O.-.��A�S�S�yD"OPy�ʙ~����n��o�`1�"O�����+��'�Y�>ԀlӦ"O)"�����[�l���t58�"O��%OB�Z��K�F�Rmks"O�Ea�gً2�AqPeˠ#�¨�"Oڬ�d#&our8`gmM�!��IY"O�ŃE�� i�R�9��ؾ<�z�w"OԽ2WK��J���Q"O��Qg��gJ�yԉ�+��$�"Ob�{#@#*"�,B�J�x
�'"O`�u#�]�vI��
hQ�p"OTiA ��"G��y�-Ϊv7��P"O��3�GO�x@�P*)���T"O)�RKNt1��C �\�k};R"O�!Q�-K�`� j�^�� w"O�]k��;��=[�.�)D���"Ǫ�`�# g�DAp��d9�"O �:�(��?#0x���-Q���"OL�8�L\%R�4��*҅$��@"O�9�4�쬂5�Z:I�V,Q�"O�Y �.]]h��ř�Y�"���"O<��c&A�xs�I��
�"OL�"��r�h����,gx�yU"OlCvG�	�eQ d��
m�4
�'��� A��T?��V΅�:�J ��'��ِ�읻��}bU�S! U�
�'m�ԉ��s���l�=NH�	�'1�H��l��m��͠�셍Q���' Z]�G�ޠb�,a�s͋J�ƨ��'`�0ֆ}�p�a�ܵ@=:q��'����C	�s
-�"�D01�r��
�'?0�/�6��̨�f:ZB�$*
�'/|"PH��l� �A��	h���;
�'�hR�G��*� |�
�4|@��	�'ǖ	��٬M��X�D�D%~�A	�'�Z��!U�{ڐ�C�ƒ$k�h!	�'p`R']2|80�S%�62�8�'�z�{�hŧ}�:H��k�"<��
��� ��e�Gvx�3�fO�d5�aI�"O`��@�7UfV��e�0h#�pj�"O�9��)��"h���MT�~���"O��i��4ļ{F@�4j8ə'"O9��?!_�X4C5O�	Z"O�q�m��;���̖B7~!�%"O$���o��t��3,]J4R1��"O|u�"�_T^��@��5%X�`F"O��1�`�/h�J�c�� $�b"OR�B�+�C�I1�-� X 5"O~���E�5M<0=bW�Ъ)���"Oh0�_`ظ���Nה> 99�"O�ͩ�����E�g��\��"O,I�Q$I0$��(�G��x�b��E"O�*���
͎"P��(����"O�( �I)#�����D��2�"O��`� >����`�X��`�"O���bk��L�y�f�Ѭ]�-s�"OL�Y�烔/8�La$�V�d�8UJ�"O�� �ɰT�
�B"�)	�BU��"OB��wÛ>k��a�B�!� - @"Ol���*�`=�p"�-�Ll1�"O�d�%�(I}��pQ� �_��p�`"Oą@PnŊFо�A#S����+1"OZ�Y�,����V�P$�-�W�Y�<�dE5������"���Gi�q�<��-�*��t!��@�k1�Mt�<q�z�������.H@�O�s�<��]�,O��@	��9 & �r�<���8U���$G/�^L�'�Y�<�<\s�H��S)ld"���l�<��[�TV���g����wO�d�<����v�H�2	�`�"ī�a^g�<I����z����ݕ1h9X	�K�<I�I*04 ��ԣF�F	~ܓ��C�<���=n�e�p�VZz�C��Yt�<	�	���2�" �.�pj@���WZ�j���!�R	�G�Z�Q��̈́����[��&:��9$�������B5|�:w���Q:�Q`mv��Ѕ�#��P��o��nli���	�Nt��z��\se��W~L���%Vz2Նȓ7`�@#4��Y�������#k:$��#}Μ����� �̣�����	��:�����	�n�6��!��kg�i���^8�a�gĲ}�3�a�0��,;hщ�dR~<ʢ �N�ȓ*8��2`����
Z�4&r���ar�s�^/�h���M0�\�ȓLN�Y���'y� 5K6$J�V9����u9��"D�{dP�`K�-�4��d�8��cnϔ\~Z�f�'��0��6�|X�P���a�c�N�{���:@x@a�2���c���Lu���ȓb�&Tf��/zLԑ�6nN;A���"�d��m�62�������)��ȓI!~|H&E�:�ȡ�(��2� �ȓ2�f4r'aL�=�ͩ�"6UԀ�ȓgFh�� @��L��&�3�݆�$����醤M�6)cj�=G�!��"���ˀG�Pp	4���0H؇ȓ{UT]���ƠݒaIEF1*��5��.<d3�bWw�(���\�E�X��*g�)QQ'	�(�c�N��p���S�? mi2I�(�fͱ���jwf�C�"O��p�"x��CDE4��"O"���L����z��9w���%"O��#(T�=or�A��1;
0�"O�$6n̙Q���"!L)8�eqf"O���ĪG R�6�`��ظ1��10"O��	��21]|)��:[��|!S"O� ��"�������v��y�"O�0�#a�:r�r �I�K`N ��"O��q㯍�q׺ ��f�7]��!��"O��âIV�ık��\�nHp@"Ò��A�.�օMt��a��"O�%	��T��3�S(F@�D9V"O�Kc/۞~T>Y�#˖ �R�s�"OJA�q��#M��T!`�%��y�v"O|頲�'>�C2K�qz`��"O�y��ӥ�؝/�$[s����!�G7j#j1&��m�
R�@0!򤜐[21�t�E>�n��C$ىH!��'B����g9���&��t4!�����!��7O����3!��
�"�s%�P��6	9�@�}!�d�p!�W�YY�v1�P@���!��>�4�6HS&�tm�n��!�$:
E�0́I����kL�l�!�ɘ7�`4x���)���Yǀ�3�!��P���y� �_7ɴAaE�ԵO�!�D��sl���c]�~�x�p	�t�!�d.!�:ahL�ڹ�hF� �!�L:v��Q�U��'�شy�%͇#�!�䍟'�r���]�z �GF��!��ГsBn���
�5>u$A�Fg��kl!�D�,6��	(�U�Aq���e�)A�!��}�a�+�~��u��
	L!��	ehȨ���^\�`e�V�o�!�D�f* � @�V�<o`\���_?z�!�䔷97\��(o���L l�!��#E��)C"���r�@�A�!��=J�@9p��014Qp啖�!�ϸ;��$��Jɪ�n`3D䟅,6!�䟙w�=ZWǪ��|�R�ڲS!��:G,@��E /v� t���F>!�$B*aO�q�R*ޑ��}Bā�#u�!��E�[�̀D"ͻL���cd��(<�!�R�sn��s+��3t�HH���8:�!��]�/�Rm�c$�Vs�t�qA�5S>!�$�Vቓ�;}�5�@����!�D��Y��y��,�}�P}�DOC�^�!����^�bm$I.��D�6!�Ā�`@�Y�F�`Μ`+�)G!�yE���%ڬxZ(#�gE�4!�;X��Y���X�=P�d�� !�D��de��P�z�A���ה%H!�$����rDCS89��ˎ01!�+{�(���>I����F! !�D�=�	0���1~%�/[/^�!�E8��� ��q���Į�{�!��ښ�xQT�(����O̼am!�d��s���w�޻�`�d�lN!�� �o��`�ʔU��SРjG!�P7<�ЇE
�D�B������l�!�$ơT���s�Ŕ5-�$��d�Ϩ !��0~��,p̄��`Q�*F>I�!�$!KɜUj� ծv9��8��öAK!�� ���p� hFBPhB�ʚH�l��@"Oԑ+���)A��9AQ��:lv���"O�- P�Ɉ}/��⑨K�1�ٺ3"O��PE�J�P%�|�A��a�$*�"O���K.˨�*�d	<z���S"O�̣��Q	 M�����U�2Ht�"O��Q�� ~!¦k�,>�Q�"O���uiWU,bꒅ\*��b2"O.�I��γr�8��@$Rf8�D	�"O�y�v!��,@��S�ºa,����"O��C��R�{]ص1�ѝj}l#D"O4���� ����$�T�*o���"O�ɚ���'@ܠ�a��`n�EX�"O@�Jc�%A�c�`H�il��C"O ����P�(�M	"�Th%�U"O�x�T��3v:��M?PH|A�5"O� ��ӽ\�X�p�ĆT>���%"O$���

T�n���V)^0�\ȷ"O� #.��l|Ā��+Q%C#�8J�"O�=15/	���p�/��R��$)W"O����>v(�Ia��D8w��@�"Ov}�Fǻ2�d�0��2!���"O@�T�3XX<@������
@"O�l����&xX����¤]��IɃ"O�I�lUK5��)J ����"Oj�q3IÄ��LcI��B>�\��"O� ���~�D�F�N�!Zz�{�"O�]�0��/[�����EO�p��"Oxp͇
A>�*͕6q>:���"ODxA��?9q��+��O/+��`�"ODB��Q%nC�=v�X�%��V"O~m��MM�[.͚W��h�*�q"O��,�6>�a�R:OfN�!�"O:�#� Н}��)��K��(�yb�X��X)T�s���!N �ybFO#A=`����#�s�!��y�邃H&�#�Y� m�Ca��y�O�=6(��͛,0�T���y�͊��S�C��𨄏�y��N6R�.H�a�k��;A�K��yrd]���{����E4fK��yrϐ$;�z	�g
��v��ܘ�g��y�*_�B�h8�O �z�3�yb�;JF�Y���jT�`�����yҡ9c1�T�E�i+n�SPb��y�׮��]�-YQWr5�l���y�jP�omp�{�gH�Ep|$���)�yb��j��l@���0n��;���:�y2C��4�
]�uF� C&e�C��#�y��`�}�7�5AB�k�%��yRo�"AI�t
��X;g$A ��[��y��ȦY��!󦈣O�������y����8��a����W�>�y�OĹ,B�r �La�#J��yR�S ?�X5a��]ӥ�^��y�I��{��\,@��9eʧ�y�-� �Y�D�K�ز����y�e�:�����n�<�%���P#�yb�HU)`ↀ,�<C��y���YkJl�F��#�h�����y�FL�t�P�Z3$-h`��)Bծ�y2�S;=^:�ٓk�
]��$��Ǌ,�y2-�T���b@-T-�&��'�yb
O�(���Ԍ7PZ��9u_��y
� �a�&��K݁�I����+�"O��R�0p�^�`��i�|��"O\����%hW���4bZ+	�JؘB"OfH�Cʢ!�@5ɧ�
�R�Ƹ"OԸ�b�O9��tRċH�<�нX0"O��kQhՈ�j@4��U"O�$��6EJ��[�����L3#"OF��nɍU+�)�W��#c� Z�!�d�+l�Pe��Fp����Ks!��y��=sQk��)�P�+��BA!�DV9GN���F3�~<I���n2!���m�L��ʰ$��'�EJ+!��P=v[�!��c\�#���a	��!�Dޙ+�h�
S�ܮx<d���M0�!�DؾV܄��ҊS�4ڠ'S9s�!�\9(��$Ï3z�U@e�4<�!�ߌU�^e��Ah1���0l�!��13�t|���R�:H�P�D�Wr�!򤎷K��t�7%l��@˔�&�!�D©T��tu�~vP��ލt!��
!G�VD�ef�t��`���M_!�$��=��jR�֖c�F��o	��!�$�f���"CQ�I���ZU�"�!��02�2�����5e�x��+�~�!�H5G��%0ӣ!ĔL�1�O�" !�W�A4�i�
�n\."�B�;`���OÆ�b;0+���C�ɦF�\<{�;av� 0�-�86ctC�ɓR��{��˩#T�,.�hE� �4D�q�L�|�x1�We�7���:�3D��@��wY,pjUg�_�d�N7D�h��jS:pv���[3fz��e'D��B��W��h `T�7C�z=���9D��1$��O����%����5�4D�@k4�?*�4�jJ�1�2����3D�P������*]{Q�Ý[(p�(��>D��h6��<*7��� �@v[b�f !D�8�P�A�~(2� )��1�����;D�`AA�2_��y��=]aFh��8D�h��ӧo�6uI�	NOt��!D��X��v�
Ȋ�O@@ ��=D�D:��_3H�0���
�Ot@���b(D��y�O�����
� �i� �b�e0D�\3�U)DY���ӭ�342��P�8D�DC��ۚt�,��B���I\"�� D���/�	Px�a"[%n��UqG�,D�8;�MLfO�8��M�9�1�7D� 21�Qnx:5�I"GO��*Do7D�hr������@{*�jje1�4D���/G������8$�� �5D�����'T�2�(5Ɖ,��9�V�6D���u"B�+$Эqp%��7�fy��a?D�H)�F|b��v%��~&�#2I1D��Ãh�f
$�)w�@.E4�E���2D�@*�@��
Mئ-޴`�n\�5�1D��e�߄BpY[� _�x�U��*D���T�}�|�����Վ5D�`��V.W� D8�[� �\a�F)D���#��w �XT�پS���u�&D�d@�����x��0a5ua�F�%D�Xpt%D6.UŚud]��ȥ�$D�$��gA$��)�N��ib�h��)6D�x��-O�G����u��6.�zt�2�(D��X���� m	�l�.!)X���&D�� �����l�,�yG�%�&X7"OnĒWM��8#
 ����E�d��"O48���
�o| �k��	�\���"Ob�igLTc4Ji���DҒ��"O
�ype�q����bKnb�8�R"O*!a�,�z��{5��Rl�@G"O:���%��j�̳�[�n8�ag"O&��C�8"Z��� c	 ��0"O΁QJ�>"z`ae�4J&��&"O���rF�3�h�"fC�&�q�"O2���d�(��̀�o�'��-�"On��t�֑.`yGZ�f�X-	G"OP�@Մ��{zJ�	�ʨXnИ�Q"On�bB��J����lD l;n�˅"O��s,܍�IC�*��#Oh�â"O�0���+���p�(Ι58�I�"O�H���`0� Qa߱3�%��'�"��Cդ]q<�G%F�?�� ��'�h�i"'�{�L���ܒ;�JeY�'�j���b�v���� a��aZ�'��H��j�\�R��Sb��DlFM��'@��`6�Gݘ ��h@6��-��'��p��DL�̺�y3D@&!�$=�
�'����Jk�4��lރ@��	�')��lǾyH�*�B�y��{	�'��{�nÓB
 8��
o�D#	�'
���
߂G��c"(e��I1�'0b<ɰL߷"$���"�9b�b���'�X"��Ħ/�dh���Y\�P�'��]���G@��R�*F_w���'��q���Ժ�@T��A$����'U8mPҨ�Bb�q�3�߅�X<��'�`QC��Ȇ9x�����u
��P�'\�=�@A�Ј�SBHZ�e� 4X
�'M�M@$,V�ȭ3�B�\��}
�'��@���5A7֩9����eܰ�)�'b�@S�X����c�݊d����
�'=���7�Q�c�4��GW��~�
�'$ݹǦ���@;d�0`y�
�'��DRGÈ<US���&i΄P3�
�'���k�b����0V�[|�9�'����q�ECV�r���&L��ei�'@�ࡥlT�3|�N��xʦ4�'d"�a$�t!��e�O�v�գ�'9�k��"Dm8�OG=p�f=��'6�!�g���'��� h����
�'�z���;��ZW��#f)t��	�'��A@�Ǒ̮e���(gQ���	�'���cv�06Z��	�B[^��1�	�'�2 $�V1�P9�gLFcB�		�'��0	����nD���f�ELR80	�'�y�k�2F,�:~��dYW�G�<�e.,+.����IŤ�����J�<A�&���*y� E�13���x���z�<��00� ѓ�FM�`!<]�E`�v�<��DٰfD�Q�A�K&d����/�o�<���Na�!#`چ����t�<��l�%D}R����̩jS���5��L�<���+�Ei�)�*@��,i�I�<���U�>(�e�-���8�*�A�<�U-��6y��r�mɥ`��]@��X�<	1&ɢ@h���荤iH��+r�MX�<��R�؆,3Hrt� c�/�Q�<)��P�-N�b�
����$�F#�K�<� l(����>#��p��ҴG�P���"O��9�|��]�Q5*�H�"OŘ���q,=ڠl9~�x#5"O�1�B-�0����S�*ty%"OҐ#v�v�Э����[�\x9"O����S���D��2E��L�f"O����yui2D�%��Sd"O��I�J�9e0��h��
�c����"O��*���>ڌ�#�hŮ.����"OV8I�+�l�����O�*7�K�"Olb "�*LE��p$�k�t�8�"O����|���>E�ބu"OT�l��#z\� ��M9sH����"O�=0�a�:F�\p�03)2�K1"O4���Z�~"�B�H�HE"O���>UP��%_�W
�`��"Om�s [�r�j=�cCG ���6"O�Hѓ���Y�  ����0� �as"O�`�fnЬx�V�2`Z�w�~,�@"O�
Ы�1JrX�o�l��L{A"O���p戜~��T�V�Lpj@��"O��ʔ�Q�2��I�-U���{�"Oʽ3�攦#ȼCF��
�8��"O� �G�2!&�I�Ÿ_l)�P"O�)V�uxp �U�P9��"Ob���W���H8�"	Nt1+d"O|{*G��-(�ױ'7B��T"O&��f��E�m�e�L�O�Xm�&"O,0�a���o}V��nS�w��y�E"O~����\�Jǔ}
��V�H��ձ�"O��:s�9+Ԉ�@'X#U�����"O�Eic�͗��A�A蛜;�upc"O�3GK�7]��&fY�*���"O�4���-��X �B����"O��z��< a�@�H��8 "O�d���wO$�`W�k��%��"O�Qp�̔z�-9�.��S�T�"O�UړJ��m��A���Hc��"O.�9����
�ke,H nn�-�C"O�u��ыz��P�9�l�&"OE+�j��E�V�b�(o*@�D"O�<���I2KFD���L��rv��!$"O�9:��x��d���=b$y��"O���R0���bwh� ,�
�b6"O8�c�[�~�ܡ��ŏ:,�l���"O
 W�J�!.DKs�R�6���z%"On��J�H�QP0�]�>`��F"O�Pb4kZ�&�k�@��R�"O�!�\<%I�P7m�:�T�Z�"O^�p @�UV�[7�[�~Hȥ��"O��卺Xf���@�^F�3C"O�@a�$�����@a�3g)H���"O��0���%g�,�)�=��s�"O,��NS3[�P��ِ��S�"Oࠃ��@VZ�p��]6`V ��p"O�E2�Iɚ%�tS$B�GR���u"O�t �"�-%-���
�;�6`�3"O&ɲ�G�@G��A���Q|�ejd"O�Uc��d�Dd8�NV?`x���c"O�u�%B9��
Cg	S��HB"O��Z�W	ELt
T��"�P�xQ"OB`��ʑ�3�ݱ��=�V%�u"O�]�3�W4ZL�µ��@��w"OR�C�AV�vWv-�aϮ�X��"O� ���b'�G�B��a&��
�V"O����d�[!r�i�x��K�"O��"S8�E$��3��m�F"O���a�R%P2�����ͩ;�V8��"O�m�	4\g�iЧ���c�T�8�"O�m�C�((P�X�'��H^���1"O��P�e�3W�i�C�4�X��"O���$D-j{jl{�c��,ˈ��F"O�Xa��^�>=*�	�;;�����"O��SQ挖o �e©DL�z �V"O�y�r���Jh(��^��A�"O���$�=H${�ȝ"����"O�U����Bȯ�F��GNAB!�-�xE�GoZ�x��4f$)0!�� ����D£E�Ĉ��*!!�dI���z��[!8�8�6L"1!�ā�8��괣�Y(Z)%n��b!��/`(ĳ$ U�Tv����O>Kv!�$���ZqPG��N�n���H��/�!�d�<u�x�B��)�2�z��(V!�J�5sxT�e\�4�
+C*��j�!�Dۼ-Μc���;���"p��,!�$ݪ��r5�Ӛh�0I؃�  �!�^12�qk��&{Ym�񇓎Q�!��A#K�\ؤ'ól:R�
GHSm!�$�� ��gME>.0���2�!�ƺn�X����� &�a����#!�$U;q�~����ep���FIZ�  !�@I�bA@��Y�f�P���M/)!�$�/�9@�)9TF���a^6!�WX��qP�M�+@j]c��˺h|!�־W�)��)�+%���,�)4Y!�D��&���h .T�>�H����'[!�$�.~��g ��l�D�s%���!���m����&^~*l��A�
!�]=R�Uϟ7s�%#
��7�!�d�&xXh����m��@�	�>J!�I�C Ñz�8�W�I#M�!�d��Kx�� ��
K�\{d� �!�S�U�̍���OCq`���r!�@�[+
�i6�ͭ�d���lV!�ž��E���۩+��Q3���$!�$A;?k���8[�l	�䮉>s�!�J�Ej� 3�mE�$�܄C�n6;�!�$��'p`�Ӧ��!�^Ȱ׍��!�dב%4�$jRK/�p���-�!�D-G�Nap0M��D1
3H�!�,fU�C� �J�xG%�'�!�dT�ϔT��ӑ�~��&eЃF/!��R̄�P�V�!�^�� ��3g�!�ק%�=9"S���=�@G�!�D��Nn�Y`�5?@��r���XG!����](7E� DE<=#� �/O$!�D@:Ä����݇IѤX2q�	9.!��'�YBԎƁ�^D�g�I��!�D�X[D�1�
�.b��̃�c��:�!�_�`ɌMc�ަW��hÊ44�!�/X��'-f�y�I��!�ϫ/���0hۣU�p��s)�,�!���3��ct�F�\L�i�p��- {!��D���d�@�j.�y#��<!�dD4'�x��dT>~�x�� �!�U�	à�z1�?ܠ��-!�dϣz��@��An��2���7�!�� ��k��E�#^��S��=taj�"O�d�ːg(�㯊Zk\=�"O�HP��3�Дo\i�![v"O&=R�c�L'^�i�hȱK8�ib"Ox(�׆�\Rr�A��Q�63��"O�=�g$A�6������.Pj)	�"OAZ�(16t^y��Ȍ�0T� �"O��[��ܳ��s�'��Mf��g"O؍b茿'�d)'&\�]�@��"Or�9���'�6erc��r+@�h�"O2��G��Z�0J�DF7��1"O��P�hD�!X~$�i�mu~XX�"O"0 t-ܝJ?"(��&v:J�1"O��;d��	)�����-"%*�R!"O�({f��$���!�
�h��"Ohu�c�ׁA<L�FBwL]!V"Oj	H�Ǝ�= zh���̊B�̀V"OJ�2$+4U�|(���
9�xD"O�I��Vur��	 NE��d"OzMX3eߚ8DR� m�6$��7"O���LS$�j���M4� �"OzQ#ЊZ���
�((�V��"O ��Y��ܸb�.�(��s"O�왧�����@$#PF��� "O�%#�F8ࡔ��]����"O�Q ����yG(�B��x���Q"O���$ޤO����!�"��"OV���h|u�]&��y�pa)�"ODlk!��<�a�2Ζ���`�7"OH��AGH�*sT��U�B�|���"Oh	��L[kVH�H7P,%tQ(d*O|�;[X�i�4&Nj{�X��'hѓ ��)(\D�F� ]*t�'�f�R
�yU�/P��dʯd�!��
1������b���s&�E>n�!��HVQ	�$ҕF^L�`�l�;�!��"�B ��H��bc�Y�K��!���X{eABOѹ!D߈(�!�D͡n�z$�7M�<Hyi�D��yI!�$֞;u�$�D'�M5�!�%n=!�$RZ�[��Ԏ42�!��Y�5!�����N�E}LI��S�g!�� It�B0b��#{LP�R��!�dB��A#1iC�.�x�+W�!��[�t���aG�3+�����*J�.���!k���0�^-2O:x;Ճ���ybD��
�J���D�-�Zq*�C@:�y��G=|�� ���!;�����I�yR�S#*��-C�hftD
��T�y�l��vdZс�J|�1
k���y"��':�AX�=?e(��R��1�yB���+9�����%�͹r��;�y"��A�|	C��Q%���Dˣ�y�M�"LN g.ͼT�6|yZ1EvB��0u��]JQt)�A�dʬ%2C�I�I�`hdn �ph�����_�FB�I�Y�6��`�@�rP�BQ�)1:B�ɇi�Ek����%A�E>=<"B䉓Y �9��,�$�9���D��B�ɽ,��Qch[Ej�͒��E�L�B䉒)^X0p7�	�-3��!��^�k>tB䉗~�b�����21Q��/H�B�ɵ;z@�)LF�p �{�C�ɺs��L{`��H�d�a�l�&&�B�)� ��*U�ݙs	~x���P�\�,Y0"Ox�r� _5�*e��H�~�m��"O��b7X�,L���#U�t�3S"O��7*7f��<i�c�i��a�"O����m�r(��DBF\�z� @"ObDɖ)�({���D�U�b�2�R"O8�PU qhX�Nͪ�~|Q�"ON����:w��0�g��Nt�XQ"O.,�aNB�!��M�B�LYa9��"O�4�uf�(����*�P��*�"OH��Lӽ>��]�F ��T8E�1"O��CC,S7.�:ԑׯ�I�x�"O�Y�@I3z]�q�@��x�"Ox4�-�<6����E��Y�ԽR"O �d���EC��C��U\HDٰS"OUX�)Q��@�Y^d�
�ju"Ot��vf��K� ="� ��U`�"O>A�LX���+Ӈ�1>��0�g"O�0&�N�'_R��t@�+��`�"OYCC?l� J���6q���"O�Pjd� I`��+�KZ!e:���"O��D��h2�1p��	Q��dA�"O̍�`gڛk��Y�p�)i��� "O��Q�/ΣOh�B���Dzt�C"O^��VA9�0��j�-j���0t"OX�d� ZE�y�	گ�
ȳ�"O�H�j�&^�*��G�q���Z "Od�b�@:gɼQ;�GE�n�0���"O�-hC�
!�d��P���T�q"O����V"h�����'y�����"Ox�;��_��z�jL�I��,��"OX��grU AaW�B6a�����"O�m��J.(�E���T�$��$B�"OP��
P�bJ�kW����`m�"O�� V���J�ص����u�8ˠ"O>� �hո� 帀"�a4]q"O<5��f9(���"���<~H Q��"O��H��A.7��HA'W)V7�b"OD����85)���< �Dh�"O,�� e�-|fI�G_�\�<���"O�,��M܈$�(���K�J��9u"OƤP�E�9����!�6d����"O�9rMD�r�
�Y�/��Lp�dc�"O��J�TT�\Q%%�y3���e"O����ԳE�=StD���=`5"O��H2��z�|�3��,��\�"O�����Ĕl� 1r��ߘ!n���"Ol�B��_~H��R!_����"Of�3���'.q�p.�\�Z"O-sF��?�J���M�,`S"O���c$F�=�����ZTz""OP�{�o�,M���I��A�����"O�Pc+�$�`��$&��7�� �"O��0��vv�QB���Q3�h@�"O�58���[���D� �z"O��0��ݬ(�p�S$��U�3�"OL�%-Q�w���>�\ �"Ol��n�@����˛Y^�5�"O�y��K�g�X���+@�B]rm�E"O^�SQhI�u�U#��E>nh1q��i+��j�S��M+!��CP�e	�)�'0<����}�<����m̖m{'/�i�c��R�<�c)rp�لE�@Z\��!ĆM�<�"�S�:��,��@�؎���e�<� Z	Aj�9|�`	2B�6+�,��"O0<GZ�\=3q��6���C�"O���!:n���e]�
���iG"Ob���K��8�h��f.��U��	(V"O�E��L��XNh��MY�<��� "OX �P�J�dnl����@[��E�"O �q�M1����SD�Ɛ��"O�A:�a6uֆ��4?a���f"OD�T$��bb���H��H����"O�)Z�C
�NUp1���h|�"OT�Yc*Ҁ/�\ɥ$�a��P1�"Opak�c6=`@R��կ�,y�"O({�"��V2� $bD�[,(���'���_���*qdX�Q��%`��u�D�h!�DC�|�= #��k}�i���fa�����=y��Dدc�Xp��_v��l����b�!��d�8�" �F7=���D�<D�!�d]6A���E߮Y4�(	�)��-�!��Y�
�����'|��
���{�!��	#R�����k�8@b�`�!�$���Y�P
	>i�(ZfG	&v�!򤌹-���b��NH�*�lǶ|�ay2�ɍTp`)�O
5WoFT�$)�TC�	��бÕ��.,\�؆���&GC�	�j��P�Ő�&�z@�ǡoF����?/��=A��o���8%�I|n$�ȓ>�P�ZtLE*��s/H��e��	a?a7%G�T5p�KtG�-�Ly��Z�<iS�̅Y��I!׫��:�����Z�<y��ҙh*|��w���K�Ȁz1E�K�<���Z�Id��d	ek<%r�M�q�<@J$t��(�Q�M�z��	@�H�<��%�x�P"i�9(��#l.��^��HG�\�L���$��T�jMH3�)D� �ܛ	* 1Q��-vM�(D�D*D��<n�l�&�&BaD8D��� �Z68�Őg-M��Ē��6D�4qq�B�/ 6U��ޭq�@SR�3D�����ر��s�9S�TP t�/��ظ'��5U_�(
`N�"4I^X @��*X,B�	]V�C��P=�Zhqg,M� ��;?�M��aS��&p�`��u��T�X��tM>D�����p� ��� {��@���7D��Qs�� [ �p���|԰�A�7D�ܪ�2~L0(����R�^����3D�,+�+���l�
�%��Z���D2D����k�=|.����"UT3 5z�.D�@	�n@!)��t�dI.U��ua"D�T���Q�y2ZR��2]I�A�g?D�p��lՋ"l��/G�M����'�=D��٣Z�k�q���)��3�:D�	%Ox�"�Be�5E�n��D$.D�J�X�x7F�!h]7w�F���+D���5�-I�.ZTe���6�(D�� Q��'���@e-��ș��m%D���׉ �b*L§��1��%3r�!D�q�Be�&�B��GCܜ��!2D�P�A�R:B�(U�Fh�����4D��� J�0���+7 ��n��`�D+1D��іHKl���"��J����"D���d��+z��v��_�4҅,#D�8�th�5~�mXRk�}Cj�y�!D��2�[�8�>@�%�Z�a4����*D�${�[�,P���3LX6M+N���#D�� D�P�������K�,X��"O��@UМo���+�8��U�"O|����§e`���+��`B0"O:,��gE<��|+QI��1��|�"O�y�$,�:;t�����ǔ#��-�"Of�J�c�}!�*2��d��$�5"O�ɥ���!�\@C�� ���0�"O �Z�5\D�t�RD��>-6�۷"Op�ss�Y�9����ֈO0,+,dз"O��y&���&x2��M� )^|ӥ"OF �6LG' ���Þ�>��"O,ȻGl��:����<�p"O��`m��E	4@�'^+#���"�"O250Κ�Un�kf�Z�0�$"Ol�C(Q"/{}��$�:F �P"OĬ�K����
U#�8S��Ӥ"O�kߜJZ��E�@�B���I�"O�K!!��"���ԟ%bx�'"On���&��4f���C�ǽ: `�(�"O��gΏ�/�T!�Q@W�;���X�"O��Tΐ$J!`�' �?J؈1p"O:�A���9�=R�큱B�ش"O�iC�F	%3�����QV6�H�"O�U��lS40���;`�P�;��]bb"Oj�� �B).^d YwE�0>��[C"O<��"{��r��? ֒��"O��C��������\Ӫ�"�"O68P�G) ,"8�p��,��9Q"OT��gŲP��u�#cU`�Y�"O�daS��I;L-��� ?:���"O�a����������\{�m��"O��q�B���e0�/?�"MrQ"OJu�F�4	pR �� ���x�"O0H[��Y�I"�� �j��
a*O�9{RdɴQ��ɔ�'���I%"O�DHg��r@����������"O E�r�OP� ��R.�=7"���"O0��F��&&o�z�GRF�:#%"Od�jk�1��&_Y�2i��"OY�� [c��bJ	s"OB(+��"?�P@�e�m"O��:�G��*D���:���I�"O>�+��#��|s���C�l�c "O>��c�>�*f�ƺt�ࠒ"O�����G#$%p�U�?&l[�"O0z�`�:J���"b�F�x�Z=2�"O��:�f�&y4-��jA�n�T�4"O���q��;
�#g�˂��2"O��9�$��LC�)z1��	Ni8��"O���a(^>M>�
/�gE����"Op�{�J�sk��B�ׯ �\�2�"O����	��pU	3M_9�~X�r"O��2L�0*
 Ń�&�Fe,D�"OLp����#oI�I�� 6?Ԁْ"O6 �Մ���6	�6ǈ&?�]S"O����R:�F��bK�I�Ѡt"O*��&GX�fi�׆�km�	(�"OL��ů$r��2�ć\t#A"Oj�X��W��:�Ҁ�E����z�"O$D.y�`E���O�m�Az����yH��r��q��:S��3n��ybF� xs���@L�Wḽ�Rb��yR����PAE��<Y��L�yBjΩ���8��Q1J���8�M_ �y
� ��TI�_j� 2�O/��E�"O�m�H�E�vԢ����{���"O���A�S�6p���pk>0���"O���KP�s�<����d"O\�ՙr�0`"��/4v�0��'��58 ��TӦɈ�� 	q��a�'��4�R�U^l&ti�i�9zԀ��'�<m���T,OP��@Ӂ�C�����'Z�Q3,�o���r%mI3I�,#�'B>03TK���lP��,�Ut��'cJ�$��'�l�y�^�8p��'�tuJ�,��>�@��d�����x��'ر�.���"���,TK�'
5!�$��A���B��0)�2m��'_�H�f�6�R�LT�ԉ�'�EPW��4H��ʕDw�*�'H<�+%�ğ��ƌ��E����y��Y�S�ޅ�a�_�w31PG��<�y����%|��䉛jא#�����y�hR_�l��2rY����{lzB�	�AG��Z�4Y4%�@�Q#�TB�I8��ȳ��$	 �8��+lrB��9�<ex&��~ڬ�#��b`�C�	#)�5�WmɁpݰ�[td '
B�ɶ茽ز"�$ ?�=(悮��B�I z���8V)_����q�2rB�ɐ0�PrE�ն	�X�9W��<�<B�� tb x���<H b8bGc@^�:">ap�̓HwF��酏@�v0p1��<A� ^mk ��G��=F_hD[�*�m�<��\�RId\�6	:�~��#�u�<�f-ٌRP`1��;\TySh�l�<�saD�OӮ�7���~ɸ�s��\p�<9�Bǌl�`�@h
�^ 3"˒m�<	���M �����#l�mf�a�<1f�$�7�A!L�e��P�M|!��D�-(���e<��)�UƓ~!�dT���p��#J�yp�EڭrJ!��1�Ve��Λm�R���D�!��V�]kv�!�CF�z���`C%W(t,!��W�ƽY�'�	8:|A/ĸ>!�D�v�4,����0i�J�xW��N!�D�hظ���J�rq|%�J�-S�!�D�7����/L'8^�(Q�c\>D՛���~T��$��%��)�禁2�ȏ�9`j� $ƞ;�tȈ�,9D��@�SYb��e���'~d ��T���0�e�_�nD`r��c	J�G�'I1p:��8q�K mJL�� Ђ��=I��D�]
=�ħI0rHaaSaF����7�	']��$[��7d��D�5(vBՏh���')G�!���0���1àSG�D����d_!�WD�����Q+O��q��߳77!�DNNҸ"db�b��A ��=aw!��ӞKB:�!$fӁДL�FG�#�>C�Ɋ���J �S���K�4P ���n��p�nh��)C�	�$Xj��Ў	Y,��ȓBct!�I�;��d��g�:g�U%�`���N<��p�U��$F���r�s4!�䅫�@�"��مr�l����F;n0�O���'<ў֝Y)��#�A��L5�����[{�B�	
|^���Kŝb|��C�k�(���O�=E��镤c�X�׉�>beK� ��<�&�3�ə5\���5oAƢ����2O�2O���$ڍW=0����[bٚ�M��`�'+��Fyʟ���;�Tp�ׇH�YF��7��C�	�Tp���w	Q�#o���S���su.b�pf�O�=�{�? ��zS�߬U�r���Ԇ,6]�'Oژ�5��1r�YhR��/7���Ӳ�L��~b�)�'kd8M� �*`|@Hbd�۹Ukܥ�ȓ��\��nƁeZ�YEY�O�p�&����8G�0��A� �=L`����AHP��D���S �E>"������vg )�/D�8h�OR>#/��!�.ś] ��A-�����=pt�<h���C�0|�0�"O�9��V�/�L��!�@�8�J����'�j��2��h�']Q�����)g$=@�)�~
v՚��k�<�RR5��	�.ox�8�П8�ҐXQ��7Β���;(��]S��0�#(��?�O��Q�J� ��rD��15��pB�KT��`"B�̯Eq$	Ss܀$���A�O����04���w�X��K /�Ԉ3����C������-@SG�	���Cnt,�E�C�{��}���J<8:F0�ơ�\r0�ߴv�|��
%�<"<�[p(�D�]7��d��(-��#=�ԬN�K2 P���O�V-�O��D��#	�+P�h`��R�"C��3����@ԉ K��
��q�%�f������7�d�t�BH��p0�6�MS�ށ
�Vu�SI�Obe���[ Re�!�Xw�\�M��\[�I��@UB�ּ87� y1zF�ʾq/��1�]�� 4�٩*������'���
R��.B�M���8|����	ح%��I�"DY7:R�ӷ�M.K���	ߖ.A�yo�r������R0ZED��6��3���ť��g�>y���Ęn����I3b��e�"�6Z
�Ћ�Q<���r�T5� `��]�i�#II".f���!H�G+Y�-w"!Q�e�#�u�eH��� � fj��!
��~��e�|�'f�y�#��7�����t�h�b��;��*�$�;�l��D-F��ԯ^+bL���3��amJ좐�آL��7�	q��AL��^� {�)�� P�&tǄ�)C�dX�aT�|���X�a�(m��4�`�{��ܸN��	҆*2¤h�4q�K
�3JW��Eߐk2��K�g�h$�třp\�A0F#g�LQ���2ˈO`���6z���Yuh��!4< ���~eD}��-�W�
"C#�d��g���}���Y� !>$b,gA�FC/OG�e�Wc�-����P��yH&���Zz7az�W<%na
r� +
>q��)\;& D�c�K6�~�KH�Ƒhq��#]���T��D���܋�7]>��ӍR�iA��+M>!hy ��"D�|郋ݽ\��1gL:%P�hӊ�?��śQ�{ҨS2EQ7�:x�O?�	D��kRy�;F���y ��SuAK�T������k�g�!<h��l�|�~�`�G
S� +�F�\θ���jaL`�`E�M� =j�=ѡ�ɮz��A#�8����N��'�����6v��1�3l	?�ԳANH-aጐ���� s�p2+���@s��	+N� �	ϓ��Hc��	�or	�Rd�9O�Fl�s	�.u.���#��Y�עRH�t�3��3�XAB(�+"��DIW�d&�+u���d�E���{E��,�hO��i��"�<�ɸ`�� �Ōº�4E�#B4L�#X_8��$nĮNP�,�ղT30͉�EC�K�D��\w�� L�JtM��*R9���1���@٫)2�4�7� G��&�ßZg4KeFݟ��(ևd6���OR`�A ϐ����@�MA��A�Ph�°��"jY*���#Jӛ&�k�Ҕ�AB�"�B	���hO��@�
�Q�dq$��6@�"��\��Z5 IC��L#T�b90�)_���@��@+D�� ;)ɑ�%V�ڠ ��?Q������&�p���ʁq^ayRG�@�њ#�j�2��*�?}h����JG)X�����nR+��ы7����(5��2��y
���:}���c�'��]	�;o>���-�)y�ޱ�l�2,�DzGD6�J\�fk���!��Zd�O��,Ox�7BJ��_$*�z8Q�% �S��L�tI�2���<Qb���^6����(�r0Y�'p��t*��&M(��%&�%>��X��4x�@mS$�����D��h���g	5�ug��.40�фfZ�:�y*��Z�q��!Pc|h��� �r���DN�6>%��F�Wp�9��:�-��}*É�yHX����l~����ܥ7�X��G��K$v��&G�(��u�;S��1�4�Ji�S��@�6��CG��d�r��ܕ<��l�e���9wpM�	�Hv�����U9�v�s�������v�,a����G�>2����ܝn�D�ZٴR���fٻ4���8}�;>�@�+!*�;�h��R�,�E{���R�@��R�O"]�r ٤4~b�ݢ:zl���hк{8<�+D�ʜ0��,��g��X�
����S:¸'������@�	!��i�?|�G��q�DX� ���[)O�9� ������b�rП�`@�.e,�R��Ǣ/�� ��"O����E95�:D�NH-3�d��q�D�Y9� ���D�`di��K���i$�K�FD!��)Jxl���9(���S���kk!�d��@���0��h�6*[�X!��cUz�����& "@"p*�.D!�L�?
Q���\�a�jr!ϙ�6!�֥n��*�jG0�V�vd�W!��D�0�@��(�#���{��ʿ"�!�$Q6JEЬ����<Y�0�N�}s!�	 L�4툡L?CD���h3~!�$��h��I1���z��2�g#$Q!�� RMq�O��)*b+Q% �T��"O�Â�&��-;�.8Z�M��"O,,3�B�'n~�T��ܢNM�90"O�ij�c�ީ��J�=! �!��"O��S���0�P�c4oV�U�P��"OT�"D�@�v)x|Aw�C$_Gb�#Q"O��i�(�*^K�@��×.y�d���"O\�`i�xªp1,U)�̰�"O�4�L��6���`*��*�F`��"O�݂R���nPi;�`�4m�l}r"OV� R� Hr�DA�eӑ;���R"Oz��	]�T�brfIg�@�#�"O����`�;XƘ��!����H�e"On� *��kn�a0p#F8{�F%S�"O��� �
b�tT�%lK�\��U3b"O.@��-	*O�%��垀pu����"O։ �L�eUh9F��,v�Qʧ"OD�Q�`K_�D@d�B�	�Y�!"O�����@UFL�<��X`�"O�(Q�ҍW���J)m.N@��"Ojѐ�Me�d���G�0�3"O̽�D�X!�E�\�
�x�:�"O��z7�-.՞PӖV�<�rq;D"O��䍇.O��C��TH��3B"O$J��ԩ7�I9&�7�&ui0"O��e,���D��k�8R��Hʰ"O��*�I��p���S7�J��LE2�"O���P�
�4%�qɊ$�ȧ"O>���ğ��L�D�� J3ܔ""O�A���81l� ـx�D$��"O`���n�$n K��w���{�"O��W���zy�@dMB������"O�薯�ZLTa. &���hg"O�Kuj@�q��z%K�O#Zi�"O��J$��m�N���陦.�hI�"O�0�A <s�R��[�Ba��e"O�9㧥V>]���:��� Mo옺D"O����J@�5!!��5o�D!��"O���%�d�xȁ5b� ����"O^R�
L �┲���!�>\�1"OT�@Vʃx1�$�˕D�D!2�"Ox�b�KTz�K'ʓg�PI+"OZma��27z�i�����a�"OM	E�ͧ�摱�σ�Ab�T�T"O��I�)�,�`f���"O�TEƎ>!���tşD��8ɱ"OV�h�6�>�����H����W"OA` �,+��=ۤo/t�>��t"O�$C%#ǩMCB���Eܕ$�R ��"O��s��E7c�*Y)�$��DL�f"O���FA��@Ѹ5�|���E"O�e8�-�f�Vm�6��g�<B"OB�;��.�TYF#�1<
���T"O��9q���J�ଡ�#�-$蒐��"OJ�@.]nJ�B`H�%�J�2"OVy�A�ԛMD̜y��A�x��X�e"OT����ɥ��`�@�K5s~ AF"O�Q���ٵ<����%� w�\�hQ"O��R���S,�H��*V��ΐ��"O.�+҃�pada;��ę<�0�J�"O��iU�We���a�2Ba�I2"OV�zݞ�+�M�aI�>h i� "O�����
���qf�ɜmR�8t"O�M���m�
AZS S�(`�I� "O� >m(% ��.U�x���8"����"O��[��A<Z���w��JG� �G"O��q�⎖[�*�h7&nj<�9�"O�a��g�4��TNU�n��$8F"O�9)%�8mZ7��9Z��� #D�8����Q�zΙ�a���&m/D�<PFɎ���iQ��N���8D��!���"�N�T�Ѽ~�1�:D��8���B�,�NL�"��`�:D����m�#`�Q2P��3�r��r.%D���C�%5i��s�'li��I"D�л�ᖨ�BQ���)I���2�6D�W���~|��π� ���P�&D�X�b
��@��A�:�(��:D���cGܺA}T� �_1)o�@qA�>D��{V`�E�&qzA܃7��T�C?D�DZp���\��}���\j"�=�"8D�T8�RBf�J���D>�Y!�6D�� Kƿ����#�>2p嚠�9D�<IV�ZG6�(㩃��:T�P�5D�D�1��g�e!e  !(��x�.3D�h�� ����8( We4r��1D��.I�:u��^�]�(�"e.D�����[+��š m	U~�AB$�/D����ɔ���bG��&Y�4���,D����
�WS��ۦ�@;F��X�!(D��� � Z�\�D�:J�:X� &D���d�,�l4��^>L���'D��H���z$.ݨi��}9� D��{b$��2���{��y"GH D�����Q&�D܁1�T>h�Q�c�!D�p�SIM]�jd#�y�M���<D�(�ᜪ~��1�H�.~���WF:D�lc�նO<0m��7a��Y��$D����`ٽ'�Xh���"4�#ae.D�4iwf��}�L�HU��%g�!���!D���2�96�kFL	&>��a��?D� 2$L�5�����B(�I;@J!D��Rth�7".��A�?��I�"D�� 6&�0,H)����O�j,�B$D�8[�<<+ک)ƭF1�t�k�$D��2�.�(ay~�Ҧ�ŅN����""D���%K�E,���F��6��1` D�<2�f��00+Y	B�t)�?D��"��
���{AoZ;��|sc�#D�\�aֶ<NtӇ����|�v�*D�J��L] xPa��پ"L�L�U�5D�4�ҏӚL@\���V���'�<D�L[��ͼ]f\q�a��c�^t:À:D��k'�F�f�f� c!M�8�8�S�c6D�T���D���i�-��S|�s�H6D���t�Bװ��:x�&X��4D���2�K=A��8	T�&�8����3D�ȓ�ߏ ��+3M��_"\H5$D��`����H��螇R�|d`&D�,�w	�	�(�r�H@�M{�tK� "D�T`4K����T�\W׬���b D�xB�%[�,qq %�(h>�!��!D��u�<��yQ��\�I�A�"D�(C""p���چ���J��!D�(C���X���u>pVx�V�>D�8�1����3��E ��y�H3D����ڬm�DI�A@�_��%��I1D�@�����]��l2T⓶U�E)��-D�� �ڰG	%rz�s�'Í&�H��""O� ��'�/?�AȲ$���5#�"O^ja��?.wHr"/�X5:�"O.Y�F��g��;�o���h���"OF��pBKp���'�N!�Z�Q"OZ,�n��@q��c	�R�
ģ�"O�A+e.�&0d\��"ۧd��MQ�"O�B%!԰r�>\Z�>	{R�h�"OlA�L��c>^X�`.�)o,��Q"O�5ґ"�N� �MŚ]���"OD�Q��5Ċx�Ц�C
XJ�"O�0�	H���lc���$m��94"O<��J�jt.E �Ŗ\���B�'<���f�DX����f�1��f�-6��%�!`���0��>~k���`�Id֟����ݸF9F�ӃUc\P����m�| J���;L��B�4'�6H�"�P��Z�Y�#�:h�I{�Å+�e��?j�����%�4��Ц�?y��?�.�8N3B\˱Nl):��_:�a}b��w1�y(�)F�A���y��!\i>4�!
�w�qI���5_2��&����.C1���f�f�'Ԁ�0�Z���2�^<
�

��P)i�R0Qw���?��k���F,�
vxA����b���֖A�@'וK��}qƁ�`��i�� _�j�16B<�ҬA'*qӔ�(@�^�:�H����4�JB�X����1u��YV&̻S�̼QVCI�,�B� `��ԅ�6+ZP�ē6��Z����Mg|7�?$"d�H�fق\��I)�	� l��S��W�"g�%����E���nڟ}M@�9�HKQ	�W��D�CE�t7l����'�d��M�f. <�G@??H�+�H�a��|�d�NTr���c�:GZ�0m��o�$�i��;{p�h���%�@��'u\����+�֨�d֨l�������9�F 	���?Yr�T� �Ph��j��n���
�$ȯ"������
1��*ɮsL���G��Kr,�P�AM�@aqD0[�b�J�d����مl6͂b� ٸ�I��?�P��++ � F��D�dfE��M���a�I��J�	�|x�0���Q<�D�f���x"����ĺ�M�2j�����{�p��-؎<�F��9Q�8I��������-���?�Ͽ#!LƱ���0�}IK�
�!����E��L �q�h�v�1M�jD8��)
0l��	kZrh��"7��Ѡ԰�a$�	��&F�8�𢀧K��[��($��Kuma�M�??'�)�4.\{߀}�OJ�c�)ݺ=����@��k���@R�!�3e]�0HL��IR9���.�\��J�o�*���S�GR�-��O�M��	� 9�-SfO�PK��"G�I�K��XX2�^3g�1�:�8�J!�4x �-�m�R��g�'���#���9pgf9�ᓔ ��zS�R:Z�\Y��'���@a�VW��٦O>M	!B��6��O�\%���v[��鲆W4P'��(���T(U�� $�����FJ���B���m7�=� χ6{�D��dn��C�h�����x`�w�I���jT-�n�8����P[�	�`P�4�`�w����q�˾!�"�b��Jf������iA�pl<
޴\����ŬqsLt��(�0#��K��R7M^�
�'�` ��Qb`���wi��I$�F#dLp%�M�]x���G�p�i�ؼYA P�
���9��YR�Թ':�!�s�b�^xCC�'�Ρ�FI�?L��{���y�N�Y&N#�u����b*1��E`��0n��.����'���8s̑E7 |�'%�	K������B`HF�dA\�ӎ�d�7���g� �?!tC̰&!�AQ�|tqb�ԑ,k^�{Um�+Z~ ���V&cF5�rf�=T�­��G 38�x�ƀ3-f�@����j�2�ۧ�P�M�1FE�� ��O�2"�lT�Yw�H#V��=x���rC _"�0�+�+N�h��󦘶O�4|�5Oڍf�ۥo�e�! �;��A���)c��u�֎[56���O�Α*F���f������yW����ڵ(���
¬��� Й��>qsO�!0|�,P��26�����&�.\ nπ-}��qA�*O��RJB��M�e��?ibE�)�V*P�0q�ȉT�ݳ0e;2�xF{�ɕ�1F�:b�O�B�M�V��%)��;O؈��^%<��(�Âݥ)��d�X	u6���d�{�M�EΛxq�� *�d_�^Sറ(O��� F���dA�y���П�B��w&倱T�BYXO�C�	!2%ҵs�`^�4����� �^x㟀p2��/Ce�?�X�L�H�J ��Y� @��@3D���EH�-���"�ҳ�28�c�.D��J�S-T����������G&D�0B�k�Z��Bfͅ��}9e�&D�d��C�k�"��'j�����x4�;D�4�0N�Ny�{eσ�!W��y�H;D�� &u	!�^�d��σ8D(Bݙ�"O��ÖȒ�j����J5.����"OL�"!o�8^D��7�_�f�.x0�"O����šW��ݑ���=�$��"O|؋�ǟ�_gH�@(�,�r}��"Ol�J�ES�nv�Q��r��v"O�X*ʖ]xԲ +7��Ш�"O�H�JI����B;lQ֍0�"O�- �)�9Ii�$2���9)J�1��"O�d1doKQ�&�hE�!C���y�"O��׮ܔl���Bb�t��"O���� �z"���$�Ču��"O�p�N� \�bx�DY�W�:	Q�"O�-�����b�; ڀj�E���!� V �<�t�G��h�W�h!�d�V�8U3��P� ���(�/A�c�!���3m�����[a85	��p!�$��C`bU��@�`�p��O�mj!򤃚BGh�[�,�}F �Q�e�+1��䚷O��L+�I�����T��y�"�O`�-�m�<�����hɜ�yr�G ^��в���f���gC<�yr� j��V��Q#xM�3���y�꓄k׈��.E	 9c�K-�y�b?���)�E	86�S
ы�y�GX�r�DH��,U�s�03�蚮�y�R�M��	W�K�N(�B� ��y�eE�=j�m!P Ռ7��&	��y�)?
�!��l��`��FV"�y򫅡<�&�W��(�P-� ����y"B��d���>d*E�7�N��y�Kשi/�=[�f�:"��k7e���y�R35c`�g(C8���"���y�$[�����G'܍/nP��%n.�y����M��S�5Sv�8����:�y�!P�^������̿N��	�K��y�BՌY�"���#q��!�#�@5�yB�R>)�`TzBq��c��)�yRIF�) 4�E됺s�|d+VOY#�y��W3mh~�4E�}m�`�l���yB�O�=G���n�r��̈� ˈ�y¤ 2BlJ$�gD[7r1�%�N��yb��	^��� �.��e�x�`�*��y"�<ckN��VNC *�>x���M��y�Y�;4�c`�
��I{q�y��׃+4��'X/jON`c��Ü�y2�	d�ܨ�^�t��@��M���yBa-��dV�i��5�s/�y"��%L�̀�.��a9�p�gC��y"h��_�(�f�VR��=b��ybHAȜk%Q-H���j_?�ybJP�J��h�`�8=?\�A`����yRd[}<�(�� 4����g�]��y"�F;<�"�m<PP[k��y�K�}�"1��Q�C��ɇř�y���66�,�B]�j)���y�.��D`��0�U�a�9���#�y���%=��M��B�a}�}Ae	A=�y��N16��a񎈂)F�A(��y��¥p�q�iF�!�D"��҆�y���(n	XA&T	�H0�q+\:�yB��U0�x�AӶ	4���v���yB�zQph8R��/��6n�f�!��%���iE+L�H��P��jx!�� �)��'���x"�ū;���V"O�RԤ�B�I#��4RV (2A"O���$�N7P��cI�9!e,�kc"O�T(A�P�It�	bto~:�I�C"O������f����6�;@$�0��"O�$�se�hҢ)@p
B�&�6`"O�И�톉f�Z@0���28D��"O�i�����	=��@�Őv� LҲ"O8u d��"���P1���"O��CR�	�/��˷(ܱY���@!"O�đ��ǁ ��=�V�m��X2�"O�pj!��#дhC�e݃=N�2"O��S�L��39�q�
���$]`�"O���g	/�n�53�Z�2�"O�����(����2%�+T��Q"O���(�;�nM��	m`P��"O\4×�C�N�J�n��?E�=�e"Of�o�(X}�i"5��*i�+'"O�81�D_$���UkLt�C`"OZ����� L��ag%�o+�,9�"Ob��ëʱ!gr��V��fP@��"Oȼ@Ɇ�Z���if��2H��I�"O��1hU�xEP�ۅ�Rw�
���"O�i��'[ _�n�3L]�/P�P"O���Bʨ+
�9����%/��"OΌ���Wu�{dn�4E��"O���m#L��"R��2xզ���"O`�D�̂U�)JcňI�@�jD"OjU�7�Y�x&���ՅG&-����"O�t��&ײf����b�3����"O6�ZdW��b�hV ߯C�tq��"Odm�`D�~��s�aT"x�>D���Vϝ�C#�t�D띍r�B`#�0D���&�I�fě�N�m�r5�Ԯ,D��p$V�	:��0)ʥy�&Y��H*D�����k��p��da0�Q�(�?���m\��< �b�%,� �3�i�ԑ�4'�f/��@�Z<���+�O\<�1��5yR�'�"|�E��-Š���&D�.��ie���<�A,J<o@0a�x�����.I�,�Fͨ&G�]Ae�D�>_z��Z�� �F�>1���W>M��ߎSɸ�Q'=�Z���F�� ��7Y~!(��+4�����S�t�ŗ�J%c�C�:ԥkeѣ��';֡cu.�#�0|:�jݠKHk���lj5Z&�E~����b�y��i�-6�t�b���SnM�f��5 �'+��1E��S0kܐ!���� G�d����3���-Y�
�c������V 𻁂D�t!�2�_�:�Lb��$ ;a���Q������T#��9S-���'"��1C��*J!�1O1���Mk)�m��Зf�=U(�y&a��<�F��}hd�[��g�)�' ܖ4Ad��L��h+q.�0 �ƽ��W�t�0L�-��ᐰg�)<��(�ȓB���+ӈCH�:E;ʇ�/ܞ��;����q�^�@��IAg�\�p9��ȓ{����
7��e[��ۣN~,��f�tU2��ҁ��h��� /X�Gz"�'{�aE\=���Y�J��J�'c�5��
GR��^�JȚ���'$>�jb��4p8���M�>��j�'Z$X��.z�­ڢ�̾B�2ՙ�'YT �f��0�<�)�n��=%l��'N��ҩ��%���C���:�l3
�'�D������q>v�[��/[�z�
�'K��S���>|,��LW�`J�'��x�)*^��XA2�ȏZ��D��' :U�GΕ8��݁aǆ�T�zY:�')���lU	!9��```�?
�h*��� fX�p 8DU@�rgO�^�jU��"O���/L�U���u�S,j��<p""ONM�&��@�|2�N�	�"i�"OTRG�Cp��7N��;���"O��V_��42P��w��D	�"O�[sb�O@(�c��Z�9�&���"O6� AM�-> ̂��I�LPPcr"O��
��U/��ɹ�Lڠ,�,	QG"O4X���3z�mh5�C:G��[�"O��t�F���kX�^�YІ"O � ��	q�!��^��`(5"O6|2hN�$3 ����E�Qӎ��"O�H��ߜZ��+� �9���Z�"OL��B�4Q��g�{4r�!F��!�y2O�0LOh� �KH�s��1[jӰ�yr�H8�x�c��>B�������yr
өrL��'M�D
��#BR?�y��&�n��F��E\p,s%���y�j�r�&g�x��re�	�y⊁�<\����p?^a�	�yB��&7i*�q��M@�Z��1���y��E�z
!���4d.�I���y2��������D H�7�;�y��Z��0�c⃏�:�jM�q���y�O�V��EmF�(yB��VB �yr�ɠ$���s0k_�3趨�� ��yFV�Z�����$ �p����yR�˦�fy�vK����
���y�F@�0� ���J-~-b9��o�?�ybL�?Sb�@��	�L1��@=�y��ɱ�P��o���EN��y�
DC��HG �8$n�J�f^/�y���8+�^����`��P�!�W�y�F&uK6�� T����X��yr͓"c�|)��kޒ7�9��%�yRO�O_�Iz�.�7;�i�b֫�yϒV+����Ƶ!d�� �X�yB��
v�F����Y�qy�dS$ڼ�y2��=d� İtAĔ6 H����y�f� v�2XcH�s>���#�y2�՜c��Q1�V	�8)a��_�y§C&"�Z9���/F��r$6�yRk����LpZ`C��y§�����u�
7{�,ȇ�ҏ�y�!5�Рto���L�����y�/N[x�I�� Y�%�P��yr�8�.\q�͋}(X��F�yB�X�{�\�2��wU�q�n���y��Z�K�}�&]�y|Xy�eߜ�y�̒=Z�84��l��l��o���y2JRӨɢ�$K*��p��V	�yJֵ0��9���@ռ\���P��y�Y��)�i�2|c�Fׯ�y�Kȿr���)��$'�\+��̧�y2l����ɂ��-"��e+�M���y'+i�ޅ` �� m�,c6���y�unlnm[�|������y�E!M�(u��`Ή�N�*�O&�y2�1�L�a�H�X�.`�T���y"����i{�l�2G%t2�Q�y��0庣�S?K6 �I�����y�CԷr��ԯ
25��!�ߕ�yL�\����x���2'J��y�j[	C������R��#�h�6�y
� ��[�bةm&U%��25���"O�x��M�3t��AC�k-B� 0"O�UY�D����$#�1<�,�K�"O.�h.	!�
	���J��F@�"O��ѱg��U��B�Z;�+"OvLr�!��X����7�KZ��y��F9p4d=�BW�4�����A��y2��s�^`���7-f�L*��ލ�y�IN![F8Y�E$c |��ǂ��yR/�=`i�qVOέg3r��-��yr�M?F�vei)��ut�0Tf���ybIZ7X��5��
�)2�r�*�K�'�y"���=�6mX��#s�
 ��y�b�)Z\թ�n Z&�JҋJ��y����=�u�����,a	e
K��yr��(O�@`K�L&��)b$�-�y2��@�J�@��]*$���Si�%�y�O����K�jG�U����OR��yb�����  ��^0Eɑ�yB�S�aB�b�U  Uܰ脌��y�g�'q.�)��p��d"׀���yB�ց�
\ d��?m��6A��yCA�E5��ik��^�6�Lڨ�y�(Bf��rV�[��X�%�K9�y��Y/=P��)�P�|�1U�M��y�'9��T[d/�Z:ڬ����8�yb�M�j��ŉ@	I9P�� r���y"e����ȇfՑF�F��A%V$�y2�[�x�i�qO�&V:�l���E�ybI��z�lk�l�<N�Nh���؟�y���l�8c�nC�0�����y�+�>gK�,�!�<$]b3�dZ+�y�N�!:�"%���$n�(!� ��y"*��G�T�겠N묄���Ν�yB��$;��!êI9Xz�ի�̈�yB ՀJ�lٱ��%]�M�O9�y"�؛Y�ܸc�#�֌#&�y�M2;�0�h��������K�y��;C86�����`�,Qė�y��BcЌA�m�{�D�����y��2k��8�B�7`�\Q��C��y�e��3.�l��ON��9Ʌ���y�DY1_����to���x���ݳ�yBH[�Y?�<	��� h	��1��\;�y���#l�h��K��n�h���Ψ�y��Pv^ܫW�g�4�X�Y�I��D- �q�B�q��*ۤ��I�ȓ]���	�/M����UAݧL[�=��/&@K���&�F�*��ċT�꼅�G�0�ò�c��	�iX�.��ن�R�Б"�I�<2\J0 �h���)�ȓV\�`�P�C�|�9���G��a�ȓQJF��eĉ�,��T�a��q,�1��N�$3�a^#�!Q��̮x����#��*�
�=}�$(g��)H�  ��U-��%��f�@0�d��h @��,���S��#HH,�ťI�<�ȓ50�(��MV��+!)�$Wʀ�ȓ�>�3�⊥1�t����M�e�����.�.��V<��u��A��&���"���IS�E�w̄YR�㌤G56Ї��R)�Vm_ ��!ӄA��^(��L}����Ua��
��U�����u�h�	B��=l1:Q��e������S�? �<�a�[�� I�#nF2U�w"O���tN���@	�c�W�p(@��g"OTqSV�C�Pl��p�L*�\�"O6�k5(�Yz����N�ʡ"O\р��/��,��M�=%�� "O��P��2����G9h�N��"O�#7I?g�<�BkL�|賲"O�-K�&.v�ҳɜ>a�	��"O��T���W�\�K�)�:]��HP!"O,��ƾ��}���5|�Tiw"O���R%@��9a(1��%��"O,���Ba��@�5iE�\��d��"O�E��S�Gd�$FƤw\��:�"O�p!�	�0Y����yW@��"O���l֏<Ș� ����RL*,��"O �[�M�.z�c���x: ��"O��5쉕l�ޖ*R������@/�yR�We��9�� O�X0���-�y�$w�f��˼S� y��]��y�"_�J!�-R�"�Q��U��yR'�,l$���&X�Z���d����y�W�SL��s&�J�	����C�M��yȘ1F8x2��˝q��$�o�y"�D�a��b-b�-�����yR���.�#�L>*I��H�s}!�D�(��IR,
�+=���@Z��!����0�w��"(��
�ND�f!򄎺+I`��o�"�����3^!�$�-6Ehc�>`��S��v@!�$��n�Z�����U�E]�n8!�d�.Ibv�X!��	tNZ�p�h�b�!��P=DX�Pb ͯx�X��MD�C!�!!�������kdV�dU!�DQ�^�#�ܯ�歸7���B!�8}`8:�B���L<0M�3X!�D\�9���#ޤw�tP�PN!�$G�����"C�'�tl!m8!�DXJ�0�:ѧ�h�\3����>*!�D�1V��0�:�x�鶊T�D%!��W�P�*����6\�&�A*\�!�� -P�!�v�O��FAs$⅌"v!�D��8<N4�@ĝU�<�y�`0fm!�ӊ	�$l&�� gD�8���%g!�,N[FE���\��!k�QO!�U9?'uc�ᆮg��:�% �x�!�d�0N���Э��A.LZ����!�D�%1��$9e'�vF�;G�C�O�!�d.^q�}���AT���G�C�!��N�!�l��΂/l�y7B��!�dW�HĂu��]M�mh�Oٞ@�!���A�ZT�`�������q���g�!�۱R�x�gEJ�p޲d*g%�,�!�$Jl�ش���"Dh��	b�d�!�d�>�	�)�(��9;~!�d��L��ha�<;K�8��c�l!򄅭P���p� y[�h`@���!� �:E9�0[��""�>'�!��U�x�l�1 럄A+hŦ^�%�!�Y������$H�b���N�v�!�
^~%����H�jY2%��"bu!��A	 ������`�f!�s�9E�!�S�)����-x�>d���{�!�$�%r
ܓp=5�L�r��^��!򄊤t��af�5-��Mj�B�-
�!�� !4�,&������$��Z"OvU�� 
  ��   <  �   $  �.  �9  �D  �P  Y  |d  �j  q  /{  ��  ��  A�  ��  Ś  
�  U�  ��  ܳ  �  b�  ��  ��  *�  l�  ��  ��  3�  w�  ��  (�  � � : � � �' 1 [7 �= �C &J �Q �W ^ �f h  `� u�	����Zv�B�'ln\�0"Hz+��D��g�2TX��ƕ#Ĵ!�$Ò�?Y6�S��?� ��g+T�k��G	7��zE*Pc��)��oN��7G��T�������Α\,��սtB���.L>ePc��<E�T�;�O��!������+]T�R?l$\��#��ʢ̬;�6]���:2�@�UJ6o���^�9�@R���
��/`���d�'l�H|�2f�/���nڄx�~�������I����I3;Ua{��٧(�R�0�N28_ Y���bj��J�M���?��'oQ"�*���򩟤j��-��ᚇG�Ѱ��b<���O����On���O\�G88s��]��`���T���be��'��h���ߪK����Mέ�y���<i&���=�㟌5��"k���#O�%�R1���qsHD�'{�$"�	�%�RyDG�H��̓qBu�0I�C��LR��_'R������M����?y���?	�'�?�/�󤋗q�(���-.G*"���I�h�H�D�Ꟑo��?1�4�?�лi,~M�}�z+v�BT���+0�[��,#1�� vte)�Kz}�fx�J�����O&�# ���(+!��� wve!�۟4|FB�<�m Wɀ$��Y*�D��V�$` ����tL*r���ll��M��'E�IB86�6|��{p΄?6J@��6N�8@z6��T��XF(U�v�C�M�����~بݴ2��gӈ���J5{��	U��,�LP��MA�36�Qc�K�=xL�n�;�M�s�i�U�% �<�H�	f�Z nzHx��N�x��ǈ�"�I���P�[L�p���30x��)���n�M��DDD:!���H����G'O<b�P$�' �+�<�F��$4��p�i��8�r�!!-�T���O%�"�'��OH=����Lb�,�eL#��5���#2�a���Of���O.��Ꟑ,Cg��Y�P5Ц�O�p��]���|PR���@�0�K3�O��dS �����Ob���
7��Z�)\�z��YJ�����]��H �}N���䁧20��A4�7O�Q����./�E�"�"5�`���%}�>A�1FU�h���0̜?c�ax�I���d�Gy��
�\�PN	<t��8���,�?9��?yN>����?�/OV���o��+��H��`ـĎ�cb��$�O�L{[^B���|R�O�@7=���	��"Q��@�WH��{F��E���ĳ<i#�Ѧ
���'���ݺ
�ݛ�S7r�Լ���҇�|�d�O=j���+8?l1�3kۡ
��An�c�'QC��c,��t��珈�AY y+�O�U1�ɛ�!�|��5fL�IJ� �FU�X��E�&�^* ��"�O� FA��'�K��5����<�'���E�M�-@��ǈH���F+���?i����&�V=2f+:	iF@E�
���G{<O�7M�Ʀe����M;�'��YP��7C��1�l�9.�ȹ���?�(O������OL���O�D�<Yq�قg����Q�g}��{uOԢu�v�Q%�ϓ.қ��E�D��5k�\>ͨ��L�gό��$���P�pv��q���pW+xc�XA�R'�����+:�d�*�q ,�a �B��C�}[@7-�DyD��?��'���|�!�-�� ʆ�D<���l���'�����h��OR��`A �B��Ճug���4�U�'��}�noZt�i>��Vy�J�Y�� IW�D�Kjn�@�+��0�5�w�>Y��?	)O�˧��Tԡm��T)B�ׯn���!����ܹ�.G�2W�iål�#&E�y�
�&e����Y��3'�6����\�'ع:�����@��ryx0ק�r���qn^0}�D��O*�m-�HO\�l0��:RR����<R%��E����	��G{������H�5��)*��	F���'�6�ݦ%�'T���`��D�O�!�2gL:$����6
��P2I�O��Ē�4����Of�D�+'E��K3�"0��Q�����)Ò�]� �$�!����a��F(O$��WOD����br�@R�I&=I���⪞�y�m2�M�d:L�����(-"N{Ӝ}mΟ�B�Id���Ц��7PY���Ty��'���'a�T��s��@(���.<�$�I&ā$��'�����M�	RF��}����..Q��Տ����&�'�6M�!%#j�oZʟ��'X���O!��ʵs)T����Dݠ��E�����'�<�K�"p�ȕ�b�i�N4mZ|��$ؽ	�]6e�1��ױ<�9��O`����Q4S�Q2����!���)6�Q�'�0u��	�A�>�9`�+e�pq䏜�5���5W��������1K|
��TlX/x�j����oI�����B���?O>����?1.O��S��>^h@�w�ڲ�����D�_�'�B��O�7m�O^�m����1%ӭz��L�U�HO�"��R*��M���?��i;�X��E��?����?��yWΎ�L'�h��ˋ>$�0��w�ٺj�&��f��ޛ��]o��y:D[>�ȍ�䇖%�,Y{4Δ?T9 H��M�C�-Q�jĥE�/z����ǒ9��'&�X� �4�0���t�$���&�� �#��j��A¬Od�A��'�1�b�'��ȕ�:��0$�ՓY4�`�@!$���'(��'Rr��>)�(tlM�6'���q�6�Rڟ��ɦ�M#��i��q�R�$��Z�I�|bWKŪ#ߢ8bv��;�D92$W�"$�*��� �?A���?���,��Sɟ��	4-��@��
�	A��A�O��&�ܨ��a�t�D�S2��qP	ϓRآ|F.����$+��E:0������R����胩+���)��=��OH]�����:@2�X�%U0I��)�N��P��c�`�o�����'6��'��?�CP��=Jz��EkB:V��Y"��-|O*b�p�3��%D���ԍ͜e�x=�`J)���j���oKy���(H~�����	�Z��lA&�����Y3e���ܟ�#��Zڟ �Iȟ����&��5���O@�=� p�Bƨ��2�b� 
$\��g�'�v,���*9r���H"{J�!c�H�^���{EjåIΡP#脪\��p6.�m�Ґ�=1'������4u��ɂH��<@�+�o� 9��*�3>(�'^�%��ɴ+v"T��V_�T�K�xm�����E�P�,�2a3,���Dkԯ�!�Mk,O���G����ΟĔO��B��'�|���܃Cq:��`�F(t�0a��'��Ʉ49�4C���rN�{a,�ݦ˧����;3���!ǡ D�ș&-{���qN�8[!.*]>�
$\,��t+ǁM���kW��?MI4�ɽB��BwB��JL��D3?���Hğ���O��D��^0��ʤ+J�s�tR!�&ax!�$O�[î�9�OO��P���3Roў��	�HO����Ð@�{��,p��b���q�	ӟ\�	�>ެ���ß�	���߼KG+GtH�壤�4KF�Pk�A��G���!DBߪx��u�I�E�t�|2��E/qp�Ɇ��( ~�=
Щ]a��I!�Q�D!&Ł�@�. ��M��B�[��77���DrމZ���6
��q̊O�~�y����/O�tb��'}�4�?�O��s�'��X�j���q@	Jeb,D��� 7�f1bv��3E�`��<a2�i>u�IIy��
zJ�����s���2rW liwNW��'�r�'H�'�?��+Btxz��D,h�Tr6�U�[Ŝ$�V�^�(_�T���>^Z5��E�YK&#?���ץ&U��g��J�jШ�CV�1�H���		T� E�T��Zo�y���i%B� ��t}�'�� Ѣ�¦I�^�F�@h2ʓ�&�^�dGĦ���4�?�,O�D�O��d6j��'�\A8�bəUV�yS�e�b����<itNG�y���G�7�:�Z�Hf���M뷾i��I�J򜤁�4�?Q�
����Ƞ/F�i���ԎJS�@���?Yeo�5�?�������=a��ݓ��P�v?<�aNC� S��Y���(ܻaf�6HȜ)c�/��Ey��-��\�`�r�D��1EK����t�Êb���a$A��eBBi�w��Ey�kN�?�ӱi�t�'��Xz�I_�M� ��Bg!�%�L��	1E��M�Ɇ:L�  !ŕJ?p⟠F{�O�v���$C&a@`[�E�E� "75Q�0�@���M����?�)��(Q7��O�`�vA�;^��6��9I�xlS�L�ǟ���3"=�w�C-&����Q�E֌�⁐�}Ƥh�OC��!��%(�-BFA�],���O���j>Vv�7�ł���ף�(u��ԑI?U���r�ejt僁0�6pc�>?���ϟ��4TW�>�ϧ`�r%��iR�F�ؤ8 ��e�rńȓM�@\�A2���xޔx��">y�4|��\��a�c������P�IP&�Pgݦ�M{���$ȯL�
���OZ���O�ʓ1�|���^!1p���(��(l�T؀hM�SE6�ZQA�5�ΐR����i�d@��5�d�)B��(���=Q�B݃�$_f�k�H��������ɓ��8i�(�O�**щg��ߍ�B`�d�:r�
c!�/4��7�T{y��P�?)�����|⩛�3�Fq��Ƿ8�.`xTa� WbRX�`��̟E�T���QŤ��g�
��K���#n3��'v�6m�ئ1�ɬ�MS.��)�|
���4^Щ[�E+CF��s�Q��r�i�r�'��S�b>��f�ء�.9i�W��LU���ڧ(���+-[�E[�Qx���!]�B����D &�n�<�m�GrLU���M��-t�ߩ\��H4�����!_�2��(�v頀�`HǇ0�n�'���`hx4��`�ǻE��a�DZ47J���Ȧ�i���,.��th��梸A�f۰}�"<��	[̓Dm��GG+n�\�SD�8��H&��ܴ�?.OP��Nথ�	� ��&�z��%L��&y�8����ß,�	�b����	�ͧ+֢�*&�ߵYT��p���Pqf�+��ڳb��y�C��.]"�FӘu����H�uv�QM��V8�˔�v��x;u�B�|�E���,2���R�4U�D����<��V�D��ɧ��O�|x��DO�s`�lې�5�,���<�� U�Ȼ|ͫE	�R�]�?1��4���	�Y��%��˟��6�F#K��O��
�)��������Oi�91"�'ƨ���B�9A�Lat��7>$I���'IB����2��?�b����'��)X?(H��DJY�D�^c�`�	3y�I&c��i��L'/:��D"��Mˍ�5=ن�
 �ٕ@��f�T������+���'�>���T��4a�-Y)f���D0#�m�ȓU��L�q���/�bѣ��A�z�
uE{��'l�#=�����Hz�\z#F�^�����D�:y���'/��' 4��W������'��'i�.�� ��N�R�s�[����M��Bk�| Wk��?wl1�#��M
����'cV��e�[���z�n�=I�n�*Q`n>VQ�b�O�W�D�tIE8%��V1�d�_�GJ�Nڀa���ӱa�j���J��:0.��O��JG�'�1�1OF,�YB�Ջ!җ\@p���L�yBJ�2����χ�U��2�Y��d�A�����|�I>sjŁqOU�8}n4�G��&��0������B�'4r�'�ם��$�	�|��f\"}��M��#+��Ӄ�͉/�����_��Q�J�
�6�ٴ���GyR,���� ��0FiG!,J��[ICm�r�;-�D�\Dks��E���p��j�H��bn_�RJ4&���bN߆$�h¦NS�IؠVL�J�v���O��d ��T�O9�(�1Ņ^�^�zWEK�{EX�	ߓ�'6�PDA(k�b0agF��y*M>���i
�[��Z������I��2���:mjl�5aЩ�F�D�P��! �������I���O�����I�7I�"'�),\�Â �Eq�uR�ц M�38ʓ/B=��Ux�#�`�'x`��,��1F�?tݞ5�$`����aR1�U�*�OR�{��'��7�UyB��",kԡŵ��	6q
t`��?a����'�>J��ydK�D
ZZ�T	�E/�O
]n�>y�R<�f��C�"�A�&@�{#��4���\�n ��nZ۟L��K�t	WE}��q��#u�����1�@��Aq.T�	���ǃdg��(%
�q��i�N�*�VHxf��W�4h��RO�՘�Á?2�dt������ME�q���G/Y@�qtO�/ 嶀��X�Y P��O���b�����h!`�=$-B�O���R�'^~6Bh�O[��)���+��Z�C��b�d]6&!�$8A�29�'P�y��Ձ� !џ\0��Ɏ^{�	�"GƦX����@��L�6M�O6�d�O h�/ԍ����O���O*�ݦpT�h��ϫ|���6ő=��&�O�`h^(���P3hF&Qٓ�&�*_'���p�O q�����vQ��N�l�&���ON�(Λ��^�h֪"�ɕd�|RքU6>W��̻btPXy#Ġ^�l�s&�0�(9�4-�I�1�:�D⟊�g��9:��%?$��Si�>Z����ȓG�2����-'�a��"���	ɟ$���4����<�)�3p�� f`�;$����
f����dR�?I���?�����O���7Ŷ��Ć-$N���b��.�"]�"K���c��&^�xq�~�'R�p� iʁ2���c�Ȇ)S�B��\�&�:lX#��V\����;=z(7��4v��>�'͏AΉ�qA�l��X�6�� j璕�	��M�e�i�P���ٴ��'|��8L�=F�4�R��D�1���� "Or�:�,K'8�,ad�vv����|r���v�z7�<�b̀R=�N�OZ�d&^l��@�HRcho�N~���OB�X�F�O����On�ȣ�ȏRN����/N�ds�'�	Y*93��� ��9��۾&��TE��U�U#�H�֋��^�~xC�}X��ː�_:aJ~�f�S'm����5j�i���	Mܓ7�4��	��Mӡ^�`�s�B3a��e�O���yb 3��4�٘'��Y��Z�lt����L��hw��q��8ޛ6d�-2��X0��V��@cFL�9s��6m�<����.j�V�'��^>��h]ៈ��#S#~���BP�6
���o\埴�I43E�񀃥�7)�J��%��:�wj
�q!�dY�?I��đ�c��aS�)�8]��)��5?ATl6F�J�b��L6_��p��
��^��STm2?ג��': fL�����Po<� C��7��}�'��x��<m�v�.�'��$�\$]�dy���=}AXu���;�yB��La<���n�
���2�����O�xF���Z$ 1��o�2.�����ԏ����O��D�_y~�ڕ+�O����O$�d|>M�E�E�ԙq�ȸ�tIp6I��j��9�̑	+n�Hs`j�`������s쒖W����$FTKż��'Αt����%�]�<G`5c��Y_ 4�G��k���v@���&��EEM�A����H�����In�6�]�1��3Sl$���Y�gy��'�P(�kS�md�tI��L�jW�t��|2�'M��Ob�!�Ƀ���ˑ�!i*�#2V����4S���|2�O7��S��RPB�jR�eA��G�0���q#H�Cf���#[ן���������?E�IϟX�	�`k+1hu�"��A�kEZ�l�4l�[q�Y�9�!��!G��`�;�	7r!�ÊU�NC���bTN*%�J�0�ZsdD%	^��Y���uϸ)��hذ^$�O 8F%�m>�I�`�qYN����� ��E��Y'����Ɵ��?I�.�"�R��F�XI�@�.N%�yBBŉM��#�e[�3�Z�DE�+��aכ&�h�F˓� �Ct�iS��'�|i�B5҆u���/`�bT���'8��,z�B�'��I�."W�u��o�'C���OM\^��i����D������]��Q�iW Vͨ9�򄀊I�t��ś�~�R��4�ۚ���K @��U�t�^�M��Ui��v�T�{W̟	��'����V���<�GH�x֜���$W$tZ�Lk��Us�`���%
)lF��H�Sj��*s���D�П�ۢ�כJ�(K��QT|Έ�w��O��x_^��3�i�R�'U��6�4����1�m3P���J�5u�UI�l����fV�Q�J���b%{��9xi|�S�!K�$n�%j%�C�E�l��p�3F	��d����w���4}2��O0Xv��jWYx ��OK\���)��a��mۅɀ7<xL���OL����'��O>U�f�3K
�d���X�4���0S� D��9�߿K�������y�@v�=�� �>Y��H�/��L�Uȃ�.��	�SH�զ���ԟ��	-r����P����ߟ����情�t�:5ab��u|dt�So��Yм��	ߏ��(@��G3�
��|j5�K�8���	EY�ёN�!�དྷ���9,2�Q���'�p-��^���8J!�ޘ��'t]�-8g����� �$@��� 䛣m�/4�$��w�.���.4�2��ݣc2te�3�ǈs�������7�!�Ԁ!o"\)��Q�;iJx��4m��I�HO�	-�$זM��`S��V=N���2S"߳DA.u�pm�%b$H���Op���O����O��{>5�3ʃV3Z<kÃ�`�^P:�	�Q�$�6AH�&t�`�+ȼ���aV�OE�'EZ�Y��0K�L�)�I:2�	�����gvep�8W�\�#.��|�� �|RN��lg�m۶��8�I�m��FOФR���?	��D(ݚA�)��v�<��B��RCn���p���p�߰$4^�� �5.�DQ$�"ߴ�?a(Ob9�S�i���'
9�l�+w�I���� {�Έ��'���}��'�i0M��I��(R�\Gfݫd�6IKE�H�Y�Đу���|���T*B�=�c��
�\�4�O4*w���ԭ����ٵ&#��i‌�|���mZn����-����V��0�	w~��SxH��
VY~�*�Լ���0>��BC�;<�ՉЇ��M56�)a�w���H��W�t��u���l[�%q#_.U�6a��|y�a�l�V7��O.���|��ȕ%�?yU�܃C_��K���a��8�?9�9z�(F\�k�����ЃcJu��Q?��O!"	i�J�L9���`�C�P����O��2�ǐ�+�&%�ȸ-�!po	�$i�uR-���T"����EQ��G��*tad�U���䗏B�~�N-D��5���ҧ0��SW�W" ��A���&�S���/1LB��U��T���,*џ8�ٴk+���	�0��mK'��H���ƅ,�7��O@���O���g�ى(m��d�O����OF��xb~��"M��l�E�� @�)�fB�4��Xi��,B@��7�#� `�OL]ڕ�SJ��[ �A�R��puح���W��!9�^0�!�p���'>)��ƽ!�0�r�<3��.�L�z3��&~�%��Z3e�Oq�1O6�)2�Ib�$����y ��a"O�)2�֜f��S҅�'�*GX��#��4���O��6��6$���	L�6�FP�Ek��V�֝�B�O��D�Of�����d�O�a�ܬ
��J�YL09b�B}.�"a�ިg�p<��eH���xЗD�4%�6G{B	ԫ(i����G\�@�N$��"�GD�t�&�nX�/X����$s0l��d )�"G�|@9���g�)�b�	�e�e�p�����?��$,0"�P"���d<
�ڂ0y���x~1��R���L� H�(�<'��)�4�?�.Oz ��MQ���'�0
�"R�j2Nmj��A��Y�&�'<bA�:`�b�'��)��PJGjM�%������ZE��yfC%r��L����k��I�'āgb��S��$D%�
�e#M�x�H#��T����<8ߨ1�k̈́"G�M��ewӺ4���h��<�������'�j]�����9e�E�#�H#K>	�ц	;�QS�u����I	�͇�	��?�WD�l˒$�&l��@�Q㟐�'�P��"u����Of�'j�����v����1慴f��]a�Aֻ2�����?��n׈bq�=B%��D�  Ȭ��%�AQ�刐�V�l&�QxDLT~2�0B���ۓ��	L�fQI�Ouj�A�z�:E���}<��O:y��?!���f�܈��E�g��`2�L����� *D�@��݋,(r��QMK�3���P�-5����>iZEȉ4B�:��F4Q(|)P��O��D�O>�D]� �rl)�e�O����O���gީن�ĨR��qhg�� e<����}Վ4#6(Ӟv��	a`Ѡ��IÛw8��'?x�ك����j]!!B���
��CFx8h�� j��!�>K�Or��d�K�Z�}�#�!"0����(|B��|���OB�"��̪�P#^��H!����V����	�'�v���߄RK��p'#$.�<�'�"=ͧ�?I,OZ��䦁�X����P��&[J	S��\�0-`�rG��OZ��O����ں����?A�OrAh�(:��Ū��T�����@,®[餰ېm?Z�u��ɘ38�����`�'Ǥ��C�ٮ@T֙0��ӈ�p<@Љԩ`���sgdٚC1�����6�V���E�d�M���䇜�R�6�`�Ƥe� ���'�����Y]�(����xc���1J�!���-�tp�V/�<qR$8�(�pl�'��71�d� ��Y'?1j"�Ǹm�d�!��2I�|Q���OX��?a��?�1�V'���H��H�>�\���'_�u(�b4/�y�'U�5��*Ó=�H�(T�G���9pk��ހ��ԍ DQ���l.��C}F�yq��I<"��$�O�t=|l;�N�=^h	ψ�$� �$����PB_3apL���*y��㟸D{�O6b�$�`���:fj�	[$��1FA��~��Z��8&)AyʟJʧ�?��d��'r�iY�I���)�#�?�?y��]��ё��L5[����ö ��)J�솵�!	L�E pPu�
�}��	7������P���(�G�vO�@����'U6�B�"Y"phtu��,�8#D�'�������?���}�� ��sć��\��9��&Ñ���R�"O�� �}l��dŏ[	4��ş4���DN<	��h��f	#x�nt�j�!%ʓ��_�X46�$�O����O�˓$g�EKd���X��r�ϣM��X�@X&vGĸ���'�"쓧(�=ܘϘ'$�`*�W֖��֢B4p��j&d�2�*tk�%\&X�	)јO}��J�	�>�6��PCa���]��EQ�!�ퟸ�'�v�����?����S�4lU�4�X=\b���fo�"M7�B�IJ��!��f��y�v,Ԉ~��D�O�Ezʟr˓#:E9(�0F^2�����X���(�/���?���?�����+~�e!@K�5V�� `Q�4L2H�a��5�:�b,E \Ն牙��Rd/��S��%�Ad4`r@a~Ӭ9"qhH�S�v�6�}g�h:F�	�s�\��pɚYP`�	�
�:��O$��?ړ�O*�l�M�&!�6��<iB(E�s�';1O����-����C�%k�X�3�|⬦>�(O� ��[M�S�PP��������^��s�&F|�d�<����?1��a�:-+V)+h�|`�\D.�eQ�qnH=��V�pA	���0�0<�l�*g�3�	!�TQٱh�!l@�&DC�T+�!�.	�|�x¦H�\,���z���O���=?�uƕ>H�pݩ��'�&� G�B��N��b��D?�i���E DAN����<��K������O>5�i��d��0��0F�2}Z��'��I
cu:ᗧ�I�|b�HƔ���
Lu.� �+�h����?AT�t�|9"��2>}0�����<�*$SV��� �G;f{ Hu�����B9A�(�)Nпj�x�k��Z�+wJ|q�Ò
�I�5F�l��ݱRe�u~R���?)��h���	6F�,9�W��N�� ��x�^B�I�$�xǃvϰ)2�ߴ^�.�=���6ȑ�H���9'�`�f��9���$.y\��K������I��	~yb�P�p(�p�L9�Xj���ƥHՄ����K�l�R�aA��$z���R� ,d�9(K	�D���$P��?P�R�h�J��'�ѣҨI�C�j���Ĉ gB�i@���I���'WўP��H��2�r�c���i�"՚SJ T�<��: y\\�����ε:�%ڟ��	��HO�SmyB/ʳ
40,�R#Þ�����k]�<+��\-T5��1���f<��Q늱�F-9v�ޥ`�ñ�2��l�<�t��I?x��|��M)&���w�R�'��jݷ��tpfE7\�@��w��y����Q�4�Q
��y��5+���(}�R�=�w�ڴz(�adw�
�*�(Q��u3����#�*� d��Cuo�+1�T��@�\�Ef<l$���@��OX�d)�@:� ��(��`�(P�$ xʓ�0?���r�,x�e�O,-f�]bFBx���-O�U���B�g�u���� re^��s��N��M �N��?A(��` Q�����$		i��%(���1�$u�_�C���YUY,���ߞ
:M�Gf��Y�N�Y�"躛�����)Ժ�:�,L9:�Z=c�ۧ�yBH3g��ШQ�DRZ��R��f�J�*� ����U>CCC�z�X$V$��`2��Z��c�سW)�O���'?%?]�'*���5���O� ��Lk	�'?l`8�i���4D��Б���dp�Of�1X�
)<����cR?&d�E�<
���'��Q�i����'�2�'���'�6Њ�e�j�l���JrxH L6L6豱#@��'�,���Aۉ ���z&(�'�� �!� }��݀�lQ�8Kd�	�^S�-�.A"K���OO��(�fL�0=T���w���k�+	� ��-�w�=
���E���'�ў Γ�����ψ�5R�	�2�T�B5��}c�� s��	Eǌ51dNF�]��H�I��HO���O�ʓ<p��q��TL���uAͬ0�r B�cF`��e02˄�?��?aq�����O���.A��G#ǂe�0�#`6\�L��I�?6h4�Y�M"D!B������(�L]`��16r�(J��`Q����@|��<qS�_�~T="t�7����
 d��A���''�@X�6&�	S�̈́(K*lP���R�F�j-JB�i��#=���dɉ6�.%q���n1!D�ԕ;!�d�7g�챙6�C.8|��E
�	3�M�����DA&ظ��Op�2�řwĉ�U_~�$�)�$�a��'��3��'YR�'�y8$̍"C �J<`�ٱ���U��}�T,�(�����L:^��q�@$)�<�=qCN p
��#_���%u1��T��-d�@ea���+��xwM!z��|�u.ٍ��y����I��p�|2aÏ6�PI`i�T �9GII^yr�'V�s���v5d +T�GF���8��I�D7��1�EfQ)�2`�����2�x����?a����M�$���OJ)�W�̅/�1���#,�=�$��O����(�p��s*�+z�2��'�Ø�ԭ����O������Sk)z�˒���Û'��xF��*�l��h#��l��Jd�;�ߗ%�哫?�zx�W�S,?n��J:bv�I�~�~���OP�S�SF~
� �x��B�6�ze�eb�.H� "O  ��˰f��j��E5aP퉆�ȟ<���0?ָ�p#��5F�����d�O���OXy2�+�:C���Ox���O��I�O0��+���!#p�C�9�\��r�I8ؾj!��:6���+08V�'Lk��H>�#jʑ}TB<�U�I�iP��,���t��D��)Mt�؆��Q����(��i���D/��p1�&� �ǷfhLAc�f
36�I�����ƌ�OL�d?��y�V:h���[`&�9
���+���y��B&L��Pf�1]��l�Gj�,�?9��i>���hy��L�Q�L���ɔ	
�ZTy�^��"E#I���'4��'���� �	�|��d��~��+��e:�����(����b�ͱ�.|;eR4���`}%��D�):����K&B�|���Y��+8y\;�D��3R|c'(b�jm�`��5J(�O<T c�'o�ćw�V����u�T���
]d�F�?ғۈO~@q�j1Y���!�lZ�B^V�9�"O6iI6A�	})�8օɡX�
���T�X+�4�?�-O����<������&�9B6���@U.�
AJ���?ye�N��?����?)���A�(,���Y�ԉk'��ٖ�"�t�납���ŋ�e�? ��YEy�o����\��.�-�4U���	$9����;���ჲPvb�Ǧ(�	� �B���'�,���͛�Ia�:�>��Wl�	*G��,N�c������O��$�)�'�?	�ɚ����G��.���h�I���?��'�ў�'sb�։u� ���NB�(>��[�,�
pbȪpj�<���?����?1���?���?��OI��BADM.[�}33-Z��:�����R�OH��9r��n����+���@�������ēv��ġ~bqN�>���璓 |����Y ;���'��XrV0O�=��'��O
�;O~ȩP��Al���U&@`�"4l�Z�6-�O�����O���>�&�s��D�\cΜ���.^aƝC�A߷)>]ӧ�՟t�	:DVm��u��'���O�2=OZ�+��o�<	}0T$P<��s��?������?��'7r)��M��C�b�	�d[8�

�3"���fq���*Sr��D�Ox�(��p�T�'���O�������� >&��H�Q'C9b`�$����'R2D���'����D<&P��ic`IqW_���[�Tx0�1���u��7�c���@�Ox��Ҳ6��I�����?��'q�{�,�`�n�BH�=�(XHE+���y2����?��G���O���!C��8��ভ@6��7<�ɣw�?@�V���E�Q�J@���<Dk������71��'�?�|<N`�/M0�E��a�8W�"T�c�i���1D6O<T
�J|�t�l�?�����?i���������E��D8vj��àX�c��2�M�ț�ě&ã>y��O��fa��4��?r�Kn��Y���ΐ@չ��� �yR#�5m�ب��	�����ə��M����O\�d�O�ʓ���d���k��A�"$-���R�i5R�'�b�'\*�'�?Y��?��8�%��jB��")�G��
~ 8ء�i�RP�<��˟|��ʟ��	̟��ɾ������A�8�ס��9�%�4�䓛?A���䓎��$J�,]0!J\�3��Eh��o�7�O�O���O���vjMvD��B�*�@���i��	Fy�|RT� �`�`��N�m�:�˷�'�T8�'��	x�Ify2�>1,��X�L��m�5x ��gY_�<��	ֹRP��E���>�����	J[�<A5l�&o.r��.6J���JAX�<��%�: �\��K�6���S�<��, �m���!���<%4�B g_N�<)e�_�:����5��I,zJ��B�'�2�'���'����/�^%����@|�ӌ2u{�6��O����O��d�O�D�O����O���ӫT]��h`A�T��4��zd�l��0�I�L���x��Ɵd��ǟ|��6�D��0\�)K�S���%6 ����4�?I��?����?Y��?)��?��F�E��*&���e��qe��`Ʊi��'�r�'���'6��'�"�'o^t"V�� � SA�ŗL����U�`�\���O����O��d�O���O~�d�OhP��K߃� �ǡE�Ծ��Ve����Iş�������	���ş��I�,{p�E�˘(���
����G��+�MS���?���?����?���?I���?�q@��:���ㅸ"�ju3b���9����'|"�'C��'�2�'���'�Bh߮B\����n ffP����\JV�iW��'a��'���'���'$r�'M���L��c��@��3}�VXH�7m�O$�D�O��d�O����O��D�O��$��H9���7
��skR\R	�':Xto֟���˟���Ɵ��ڟ���ٟ|���#*��#E�R,�C��C�X��޴�?��?i��?����?���?y��"��� ߃#'���&Y�%w�� �i���۟ؕ' ?��w	M�M_�4Y�L̸�]c�����a�S�+�	�'$���?OD��"^�;�`�v��:d4� ed���oZ�<!�O ��� '�P��Q�5#r���M�^���&r��@@�&o�!�-�!qў���<��-#I�-@����i1��՟Ԗ'2�'��6m�?V1Oh� >M
&Hݾ"�$A˟�ځ;E��s}"d}Ӛ8lZ�<i.�&E�7!R07�����&9���cR�Ĉ��ֶpX����N,?ͧQ�8�e���y"��Yw*��r��9��ъC���D�<����h��D�	y8i�%M��of1{E�\2��p�ĩ␓�Ѓ�4�����E�o7�l�#ͅ
1v�)S�F���'��6M�˦���5E�60�C9?I�OM1	���X§t��Y�芾CJ���Aɢyvd�لc)��?�*O�b>AUe�l�x�R��J�^t��'�<9C�i ���yR���+Pf��jFh�0r����!��i3�4�'��7��EΓ�H�fi($J�_��E��i��v�)R'�Hq��D�SN�; 6�0Qm��2��)qF��n�SCč*��n�u���Fةo!@Ty'A݊3V!�$�o�fu���o/�k�]/n�1O�{�.m��&��I�n�`�Cܾ=:��2��N�`�ڡ��hL�T4��<)W2���ƱU�����'G-g�3��]d���V@�s�㲠�"/�qp��˫a�(�wH�!@�1�HW�FQ𽠱H�	�NQj�e� �yj�Ց,���snY�*$`���O�3C-X���/�O�7m�(f3�� ֫B��j��d�<@?��'�.��'�"�'(��O���'��fOQ�Ig����2�NpXCk���'&"Q�h�Iny��'��$з?�Ԥ*6LF-@�x'镟AB�O���'��OD�D)}Zw��;CZD�KP�A�v5p<���|l�q0��'sR�'t@$z��'Q"Q>�i>mm�	0.�`a"�S99�jL����[��8+OL�d�<�����O`�p�@�?2���谢؛ ��;�Kpqp‭��4Xny��^3�AD T;�D�0�
��f������i2�9��)P�@�D�6hxdyW�N�}t��:B��%�I.�L˧$�3 @�A� D�B!αv^��b����`;>l��`�छ�)c���vb��CN`x��K�cB`҇n��tn�Zc�;�ۖ�#w��h#�g�*V"� �É	�V7�� -#l��n�џ4�	���El����|���?1�e�]Q&��d��P_Ќ��»��'�����yB�'�"�'�$���Ȇ�S��:`C� ��9E�'�r�D�0O���O��D2?I�J�7\ �"�K��'�6�+uK�Xy��>��'���'�^�,y�e��M���P�#W�W&��A�(P4 ��i�L<Q��?Q����?1��G�DflzwGV�L��p��E�X�~h��?����?A���?)��?�a��:-��ԭBG��#`� � �'������O<�d=���O>�Ė�a�,���hs�5�!!	},�LhP�Y�8� �d�O,�$�O��$�O����<#6A$>e�gC�6����`!� ��\(�bӟ��I��%���	�Q�bb>���V?Z���Wk��nx��10&W�t�	П��'v���E�6���O����F
�a�ׇU9$`���Q!Xئ�O��$�O䨨 �?! ��;F8��Zև"Ț��J�Oh�8�3T�i��П����ݯg9�}z��3#�p��V�9@��	���cfa����O.T��)����t��CmF]�5�'�N�0ФӒ���O�����j�'��ɡI�t��ē�Hs¤x�mK�*���(����	ʟ4��K���?��x/t��&B��t��	�Í�i*�Xòi���'�r���^O���O�d��O�>��G��9��C�,�>㟰�%�6���8�I�x%D�#3���o�~�
Q`��ڟT�I+N����O<�'�?�����B cpѸ�A�Q�t��!Ӷ;VR�D�O��6��Oh��|�����O�X1�o�,Yp%��2)
=���.L\ʓ�?i����'���'�ĭ��`H#�� ��(��ov��Q��ْt�O��<i�!$����M�s�ܷ �8LZ��_!�|P�!�'���'�O����O�̒�eh�$3�B�wD|��$&�� >H�Ek�<���?A���Dpm��%>٘��� W��$P��$1q���ì�ҟ��D�'J2�'�X1��'��S`]��2L3L���0>3����O��$�<�@��,�O��2� �d�
:3��c�B�[�d(���'w�	П(�I�c��a��r��ּc�L!�#�
1�|x�'�f��'u��Q�~Ӵ�'�?I��6��/�lx��� 6��$H����I���<)�����?	K~J~�Q�ۻe.1�u Y>5�����7�?���ݰ3�f�'�"�'���� �4����a���CĈ�"0;���Oz���O���OL�$��'���B{��%�
�NDC�l 8�,��.�x���:�"m����{��}���@TU��؟P��9s�B@S��� 5���H I��7�<u�	�� $��������IƟԖ'(�eSt��L��%xQ�[�[��%������y��'4b�'B�|r�'Ҭ�cw��ðeN<,�����7C���'ABR� ��*�ߟ<�	��\�O��凞�8����ͪl������|B�'�"�'q�'�"�']Bh�5���^P)pS��;Y;J�9Q�'@��'�'c��'6��'��$X�jy���G�5?d�{ц�4l��'R�'�b�'�'��iX�=�(�b�B�0j�n���	f����'-���O���Oh�O���^�"����:#��m�-��"�bU�gMfh<A0# 4{�����}/��[���d[!0���,�.P�����!���P"S�Z��u��{M"��1�Z;�v��d.� L�����+��e�튰���ۗJ��H$�������р��s�<�+#͓9�v�0�X�R!�H��T�l9��D<��ѐ�ͮD���� \,�unƘh�^И�'�)|#(p#�͟���؟���?o�\8�	ݟ̧]O�p�&�h�Qa��6��U)6��;�DX{�.Y �:պϓ���z"(���Y��g��5���~ipf�,*����X�ԈE|ү@#�?9�46:�z$LG6bX��&L�72�>�`S�'��U��I@�S����M�ȉ(-L��(��] 9!�$��`�j����k=�E��0.�d�A}�\����Щ�M+��?9��D,2���xFrd���!�����Nğs�:y�	ş��I:��h8ǯ�Kf�Թ��6B�O+��*���p�
�@'˖,_��5���䃮$
6)p�I�T%�p�F,��F�~TS�Y<������#wo:ȑ�Ř�wH)[�)Pø'��-���?Qt����iI�i�c���2���w&Q(M��5���O��D�I���	`y�;<D4S�3o�p�c2������	3�M���i3���) ujV�ֆo
�h�Cm˾�~B
&5�46�O��Ĵ|Z�&ց�?A��Mp.Ζ	�����&��������l���� |%l!��ƃYRp�T>)�|nZ�1�Ԫ�LU�rXYڠ(�#r�b7��lі��#o~�U:�hU,^CX��c�TX4�[y��ƪ9�ɉ��r�{f���5��T���iu(9��������E�zZQ��ܭT�@e���X��y�_�W(��p��O7�Y;1*��(O�5Gz�O��Ʀ�x|ցb%��6� ��pI̗Ol��$�O<t{G��8����O���O8��;�?�]�b�N�K�b�4xD1h�L?v�h�3$x]��M>01�=���<Pp@䛎�����HS-j�]"�'��ܑV��|��Q�	�L�'��|+�a�J;á�x)p�a�h�O25��C�O�m�6���<�����=�$�餄�Uj`;�KĘ!�!�W*T�NQ�O[�]�T,0w��8;�pY������~"]���S,���5�G>~��j����Â�Q?a�"�x��~zc�3�H:�dˍC��	*���<1�C�����3j���[��H�a�r\���H�\�8C�	�Z=�aD@O*pc_CC䉫6]h�h��xYT!�:��B�	�_��p#���SE3%u�C�	,:IB !�a�3fj8�e���im�C�	�(�����50����oѭJ��C�ɥE��P#O�"K�0�.@��B�I9wx��Si��-p$Q��2
��B�ɩ.��tN݆JZ���g�~��B�	�Rd��kH�_"�y��A'Q�dB�	=C:i0u�έQ��K�AޘyaC� s��h���;���;�X]��B�ɸHj�I��\!c.���Ґ{6�B�ɬG}���l�;fС�BT�_;�B�I�>=v��d�K	7P�ـ� ɡ]ClB��2 ���pc� rn��a�D�*B�	7|�<��%�q5*=;6�=�FB�I;R�n�
��I�mf$�3��IKNB�ɨ2ܴ�ǈ��]�
�荋+u�C�ɁV!0���jF1�i#3�4@"C䉢-,f���FD _
T�C���lC�I�:����a&D>$�u�#G�, �DC�W� �C����#���#v�C�	�7���3�	�w4�����Ti��B�ɁD: ���郂m@�����T�+�zB�I�/%z���Ɩ���+];�C䉃k�^����1@���BujC�	���P#�큜#�=��'��^��B�ɻ;o� �s�MI��m�r/�0YxB�	!zH<ц��g�>-I�/@=ĒB�	*B���rI�(@���u��>��C��P��p�n�q�)�b �]����@�@�x"��?7�h�Q
�G3T�)*@C���c�)��z�J��y{�XXwG�!3�t��I2�n�8A��̕7)��ܡ�����+S̠*���f@0	�p�Ce"FI��8�]S��0~�P�E���(c�c�D$
��WC��tX0����r��~�EE9S�ru�f���Q �^b4��'7~�����%b�ؕ���*;�J��P�����T�H�(H�4���-��u7�I�t ��r�A��ҹC��[�0����u���fֳH��`� Pӕi'E��aQ�̍�N%(-x�ǅ1_�0yB��' ���m�x�0��N �y"��J(ғ�D�<8�vO�(���T>a�D`�!�2�0�⟘Z�:�ص�*D� �da�� DUAe�<B��i!�O��`��URm��Dh-l	ь�d���N�<�ܩ����4猱�-�ǡ��?l:h-�nK#�����ͧ"^���c�]縤`�K��xu�\" U�m>`9Ѝ�Dת���ED���P�cR�-?Jay���Hb�x���5_r��2��7Vu�2+P�cJv��s�JWTXP�0�ն*�M+��'���r�90D�+vLX��K<�w��15���'\>^�:H�'�*y�@Ý����=(@�U��%f�pb����yB�X0R(f\	�.ߥ1��`B�E��33�%k%"5��qJ�N�v\@H)s�p�S&u[L��w�~�q�Q�9er�j�Jc�%#
�')D\S6��f�hɹ�ȢQ�l%�5d3��06�>=�z�׀{Y�Msf�^�b�Q�Dt��IYJ�㔉�H�X2�i?�K-ZH�bj]�O"�e�g���I�89��Տ�M(FMOc���ǭ\�N���`_�a��x!��
-�r��ǋt	 �p��#(��{��Ȟ_��$�x<<�2I�Dނ̱���r<�pǂ�,��K�M�^�~�P�@�7I^���K�xx�i��$���x�'���yW��W[�{��ܟC$0�ԪȞrT�	e�]����@ 0���I�uD�Y]d�)`nO�#i�;o�֙�
�(�P$�����W�'�F�3S��m��Q%65D�����.B��3c�� WRhK��O���zT���7�.-*�ŷ6L�0�0jK-Eq��k�Z�@�%�ӭQ�Г
W6��uۓ� �=:P�El,R���ʗ7��Y�SA7Z�"u)�a�hx�@�Uc{�	�B��t!�.���R�	�G]�$Xy����Q �Oɠ%J$���n��_�4)P��b�,"�R.��ՠ]5yvH"�y��\�q�ER<}��`��h2�Ec%Ӡ�*��莆�p?���Dw�&=�V�@
�R	;@�9	^�0��S�o���m3����'��p����h��=� L|�U�eIّ$1�`�F��iupaQw;|O<Ȁ��q^�y��	�"3W���P�)<D�9��U+��ZS�˘
t��S$��RtD���͝ 7P���ЇP+9N�-i5�)���	;���У 9��Ӏ����'�j�+��tL����D��qx��G�T?��Y���x���.�8zo����䒎O$���i�:�­�G��hD:͸$�ڟ{����U���Wk0�j�˞�^4���	Y0�I*�R�aШ�p
��P��գ��Sc �R�͋��P�Qh�
\8�4.;�
@H#J4,3�[;S�i���@-�a~r�P�Gt�U�$�#b
䳡�H!xr �Cg�NDh���A��� ���>Ay�y��$�i���I���s�*�0^��9+A��m��4�ୟ���=���
2��+W��3X��� �IP�Ej��tcނ_|��(�.\�-���9K;����Y`�����0Cf���^�\z���'�.�`�I��6�hD$C"L��d����.NyxTA��Z8vI
�(H�F�����!U�Av����'�h�7���S$a�5o,4�QRB�G=|H �[%S^�|��R�I0"8����Սt��!֨Z�
;�#8EfN�@�g	f���P1 =�;�&Ռw��9�h� ^�){2��y���C�dxk��A=3@䴑�aض[�R���70m������'7V���ǗP}"|��ȟ8��qҠC��nl�g�64d���S�';J7-^,����0z�<8�DM�� �*\�vI�&�����4J�,��e�h��&@�)�\8�υo�xyZ��j�Z � &�T�����'4��f )�P ��E�n�|qJ�'Z�4؄a��Ox���H'�j��D��t^�,��R�L~��Ү�&�z�EʃL�&���,S�B㾔I�Ɛ9O�1m���ar蜖1/�� R'	4`$�ID~�V1�"�k5)�<WH�p�2�p�b뗯B=T�8�[Մʧ)����)��)��-1ǫ�}Ԥ,���`�V��N�W9��0�
�+�*���j�%�4�?O�"�`th�:cr��$Q��u2W��Ax2�!��0�Y2u�ߧs���y7
 �̥{�A	`��)���0?��$�P^�5E{P�`�l��Q�: rg�E.PR�E�%̤j��e
���>����O���FþLT���O�_`b<!��I�B�a����2Hw�(t�6j}�]ˑlV�?���!.�}�3�d��y���[���Fa�r�{�A�
�p>�����h,��R�4.�� b���xLpB@V�]�t�ȓ=x$Puh�}���SlĩFcVFy�U#9p(\��IKv��PQ�W�8�T��B�A�[!��5�$�a�u�^e�Qǃ�r���f`�O?7�ς�����4,�ޤ�P�Xlax�-ϟ�铅~�L�)�Q�FG�w^Xm�s�H��[��>��n�lذ]�SE�k> $�g'�SyR������'BQ?݉�.L�kO:]Qv�Zm/���o%D�8b1�H�H\P]�(��&�ŃCb�>�'*R]h���\~��ɭ]��A"�'��!M�'d��D,X먘�2�\�d�dux2 J,0�zA"�_(��D �O�HI�� ����N�5��F�I"VHh`f�I�k����'�����#����!�� �E��`
�1��D���0'����T�\Cc��'�qOQ>]!,N.�.8R%�-QM>A	5�+D��6��0#�y+�h�hGa"��=�I�iCi��I�o�|ӧf�!B�~=Z��a?�C�I,�p8[�͍^�R��&�?�~C�	�^���QV��j�61b�a� 2C�ɍ<�ȸceJ	�-�
5P�m˸�4C��}֩j�d� u�5�D,B�A,C�I ����(6d�A#����M�B�	qwH(�bnX$Y<��9���b�B�	Q2=(V(K�i�R�B��4�FC�	.YWz�(��]�dR�a@�A��B�I�g=T0I$��BT�i��FĚfC�	1H5�`I��ZV�����: �B�	t��(a��07��	0��dB�	�܄<[R�4�H�"!��I�B�ɉ_@���&�ҲK�:j��	LB�I�E��Q���Y��L�gT�JbB�	qr8�sD�M��eԕKB�I�\�� R�Ꮄ]+b`�vN��`��C�	�"P�����U�e�B����\ R`B�ɐ=8y�CĹI�Rp�*�;4nB䉳W�P�ȅ�/<s��G)j�RB䉰M���82(�<k`�x���ȹ.�C�J�҄B��X9+�AR�6[��C䉠�غ��Ҫi�y����wgnC�	;\�y*���&|��e�$�3
NC�Ɉ?���hǏޘ9ӪI�2E��.C䉗6��ł!�8v��|`��`�B剓[�v	yc�58P�9��M �a!�D� H��(0O`I�=�+�p�!򤙴i.6uTe�.�49�	�x����L���X�cٱ<�=�3�'�y�k�;�R���Cٻyi��CP��y2�ѳ$����n��A�&��4�yR�U�-�� ��&�::��qF���y2DQ{pX)E �:(q�KV2�y��cJq�@# -ʱ��A��y�ɑ-;��9�L]���*�+�yr)N"
�y�A?��#��Y�y⩜-B��ɣb>:�I�R@܎�y���"o7�C�@�Hy�҆^;�yrG��S�aM�O<|�A"��y��4{t�y�w��r���!&U*�yb��{���@��H::LY�@A�=�y2��Elvlf�~;�Ts%V&�y�AͲ?��:��عdO��B�U��yʙ�}��l����^Ip�Ѫ(�y2L��sB���C��,!�X�A��y��r3���0��BP�ЄG'�y",T�@Й���Ÿ1ݜ�Ύ<�y",�.� ����� �E��yr!у&��m�@�T�$�L��UΝ��y��B�M�zr�	�<ن�Q�y�/�_~��)�M�R�r^��y�=[���#��3c��q�����y�-V�{0���d]4Yi|$�����y"bT(����_&z4��d��y��F3G������M�$������y�;V�ڼӴ��%)������߈�y�m������*]�R��4x���	�yB%֋ %<]q	�#�2�� �	��yB(7I�9�2(�'����g��y�݊W�\�����Y��$3'���y
� ~�j�(��[��9���`ݐ��"O|=i:6��H���@�z3"Of��"�۵E|�r�O�Z["ObT� +le:"�ؽu��˃"O�-9c*H�_��rTcO�U�<���"O6�bw��
#�Ԗ�� �3;�y��Kt��T���+���5�y�A�:x2����Ȁm�r,���yĝE��c�F�0��A9�yʧ�p�!�$���jp�e���y�Īh���[I۽����C��y�`�(7��<j���q��ʕ2�y�,�.+�.ܓ6��m�ЀSK�!�yr�Q LMd!����a�80�c/�2�y��x�]�c�	�Z�Ҡ��č��yrO�4��rs���W�p9l�1�y�b�8ސy�͉,N�f������yrd�:�d�k +CN%����yrgE�Xr�b���h~�٪� [��y��(~>� EJ_h��c���yb$U.oG�i�%V�]�Z��N)�y­L 8V����Ό�SS����@��yb�:�e�W.�-A%�0���yl|�ر���0:�fő�ŋ�y�ϝ&m���ڙeD�}3�	��yRQ`O�J�ᕋ,ud�����yRh��R��5�5��"?�h�q�˽�yD^�E�V�;�̎�l%��zT���yRgZ�&�����x Ћ9�p?���bv�Y�X(�.�1���1w� CC7D�L�V+BRu8�4$�x�R	j"�"D�� �	�%)�ݹ�@;A�6y�tF"D�|�Po];�0i�2,�1,H�@�F"D�h2�#��8M:�ʑ8���'-D�$��.�-+�4�2��qh.}��+D�Lar�]� ��l��`�>i�����E&D��
�h;g�|x�u?0�C%�>D�pi$/ǟ!S
e!�B�S���A�N<D�H��*P���$�������;D��qi��@*��0zx��@'D�$#v��b3@�r�eҔZ��ԙ�)D�l�Qd��t�����N�~�� )D��ٴ�J�)�N$���dn��q��&D��K���Sj&��f�'�`iJV�$D�lq��J�E����n�2��Vk$D�4jv�0�(PI��ѣ>�nY9Ph%D���#eG�1è����M�| 
��8D�H
Q�&�`��V��^v�7D����E� TU�D��%��b4�`��,7D�L���
[�$��cL�u�iA$A3D����+�g^��Q�5I�G6D�Pat�٬n���ZTaJ��]�0	&D����B:=QD�b��j�V��#-#D����L�2R��-H�G�(A��'D��A��	�1!h����8L�&�H��7D�H�"�P�x� R��B������6D�`J�F_ �"�$Y�kk����d1D��
�E�5
:D�䃉�'1��p�-D���`ē&����H�e�Nx¤7D�,���E��d=b��5�f<�ŀ4D�|�b�?P�ĐSr&��H<8PHB�5D�pb��$*-�tC����?��0 3D�x+�<�恹�k�~�Qȴ�0D�ȵ��V���µj �0�Sc0D�� z�R��M�K�
�`u�/R(I X�\S�[�S�OH�Z��.���ȉ� �4���'�lA�H�2{�Nj���t\��M��� j)az"X��D1���<J�.�k@!3�p?��@�8{��HZ�D��Xd6L���'#F���"D��[c#�* ��$Ǌ�~*����>�U�"�Vf4§Y�J�Ġ��e��|ɶ��(j
hU�ȓl<z@��ǰUʾ����܆U"� ����[��X��C�Oɛ��'Y�N~"�i��gH�nĿy����� [T��B��B<���ϜX$�����T9���F?�훇�'��cD�!�Ai��Ŏ�$����� �OnMk1G@&U����쓳1j@�5�'T$x��˒/NŪIϴ;��B�[%������d�D���d����S��)Ͼ���ɮCƢ�{�@�,\�b=���D�'8��x�'�`�
��u�H��)�=�S"j2���G�U|�T��C�	�Dbb�!RE$��u�KX2^�PI .Fb��%C�'(�)�CHa��ݯ{�.m:�$��+	"LbjG�"�C��=��xT�T<���Y�JN<�	���>�� �H\x04YꙈ�/#�b��r�էK�`=�pgb5�����.���ӽm���*��]�x)�Ո��8V�q����<��}�-X�>���Gi�:�a|ҧ۔$ ��i�<Z3<�
P���ɀ94fy �#�c�t�4.�4DwqO��+�~]0u�u&I:!;����T�y���M�M{�n��j� �KЍ�!\��9���Ą/����{ʟ �Iԅ��y����Y��]h0C��8Kd���E_.�Px�A�F,>���d�'6��,b��ǆ..&9�O�LZ��M]\MpՇzx�M���N�P�,��LC�{L�Q����XC�x���M!�0�B	*�b��4sC�AB��5|�<E`#�Q��17� \���Cd��Z�Ɠ�}��A�0b�:����(}bi�4o�t��QO�S��y���R��?a�3�ܦ4��0���a�|��Cd'D��@!��9�tH"ckF�0����`E�1J��6�.	�l�
�>�I?�[0�O'k2���$kP���n�lO�� ��˅����u!�9��ש'D�)&T�oݒ���#\~�xF�� �@T�*O�3�ɑxz��<�J��wJ��D�0. ��'�+��G$[�xJ��
��X��3����kt^a5��x����C�T"�F��J,�7�<�,
*�� +��:�9x��i�'L��|ۣg^�	l�q�	�'?��@f�C'�z����&B,��K>����,���KJ-$&8u�M>�'�h� V��L��`Ag��_k����Nh��DQ]��i1�n\�'V�3A�_������6ciƔ&�"~���ԋ5���1�׍�{�ԏ��O��B�����C�_s0�x�N*Tx��c��f:�x��e�v無@�'6��b���7z�az�!ՏQ�*� '&��N1,�� ��򄌸|�:Ĳ�'80��5�I��~��L0���Qz�h���)R�TJ��i}�5�ȓe�xm�&���j�L�GQ�tR��YڴM\du�R%�i?I#�'x���!������;
��I�f�y����v�Q�HsK$�O�P
�GJ)4� l�W��|�h �#e�����~��r�p�V@��T@�����'�(��1�F�'��DB��X3cp�4���ל[q���#͌��֨W

vxYCRg���<��+�%IS����n�d�&��eÓ�0<rX�0m,LOL��D�� �������m��Ha�V��xVN�T��I&��:S�='%����~��S1p�k��$�$\��K�y�(..9�<jR�Hބ��-�'2��+؃� ���~��O����0T����<�A��(G�?�	ˡ�U,!A @���'��@��`^%��]+���x�`��
@!���IA?���C
@8���IY0W
E(a$�S�W䀂!I�8K�,) "^P+��,	j�X��ly���j 8M����F��#+���d�

��@�(�7m�<AW�-YE�!\O� 	A�"��cF\<R� 1z��>2Μ�8$��O:`��=R�������Zw�Y8�!�� �2��"G<5h�'#p���iB�JKvL�@#��u�y�4
רZ&���lפO�qO�S8Uk`�d1�R�ےb7t�\�  ճ*i�D#
O�lKEi�0�����a��+ǘ!�*���%׎0!FE6LY(L"j6w8M�>�Fc�&�\�Y�-֯u�vp�&e]Q8�8q�o�?�����5Ũ�C�E�'��BҢZ�7-n���(�\��t
d��ty��VL؞�����L��E"ql��n�CB9}B��f��ܺ'�������Α���uGL�A�6�#`�B'�Yy�X
�y�E�60�)�6G��>������2@ٴl���.�j��T>)ۥ���% �� ����U�]��@�.§k�b�3�
OT�pg'�b(�P��?8���R�]�o�҈#�±IU���g�\���?9�>�V!@따a��Ƭ#�;��WzX�(c�,Am}��G*�p����i.�%�-є"��@�D�`~*K�i��{R%�J22t� _<����G��O�̢ +S��� iR�CI��Q�j�n�pU�e"O����lό'}L�@�J��*.�A�A^�<�g�B�S�Oq�E�ܻ`�$�ȅ�Ɔ(���'�Α�)��*(	p�N����'�r}���`����7���#��
�'<P[����4�eZԒ
�'I��d�]rX\ �$�q�q
�'vX���\	g~�sB��J�D�Y�'D��Q�@83Xp���w��
�'�(b�c�!$�.��ݯho`�A
�'l<���<	�RQ��c�!\�|PY	�'�n���T�Yp,��Z.XDB	�'�֡R&+�<���ѣ�X�S�4�@	�'�`��Чմ��=��LW�x��`��'���+�΋Q趌)po*q޴D��'V�p�"NE�h��x
P�9s��'@�i��j#9C�Љ��o�@I�'X	(�äF�a#�/_���
�'X0ܩS�_�tc�4�B$�7xT}�	�'l���lsߠ��ʚv��5	�'��d�4�V+E��,�R�D�_s�Y2�'?`P�N�C���Xb�g��I�'τ�C5'�Hb�����K��Z�<���f����L� tJ��fmL~�<1EN�oZ�T�B�8t�4!g�b�<	�V�_�@
���,<��f�Za�<�N��&�ę���:,:4CC�s�<��g�O��5�A�$���#a��l�<QEnH�=Q��b5��X�$5T,T�<9"+�!vb��J�UB�P��ŔP�<�A��;�L�E�łs��:2�OJ�<I�ʆ@n����P �̹�t#=T�(H��k�y�P&�w�@I���6D�,c�+��Wv�s�E�-E�9D�����)a��p���v��\#q�+D�@@�'7�lC����*<E�ר*D��A�ԧ ��Y�`�0��,DD5D�h����BYT��3k�h&�����2D�|����~HA���A�4Ḓ2��0D�|����?��A��lL��l���D.D��� �#`����'̗;�R�x#e*D���W��=#��R�H��U�$f,D�����v^ʬ���c���í,D���B&_�8�<����R��:��,D�88Ҡݍ+p|�p �l7�5�'�?D�A�\�b�<�!h��m�Q��(D�\C/֔f}6� �.\��z�R�M&D�����irL��$�ڴ0T�+##'D���V�S
K�6l�E��Z%�Cm$D�h����$fd�"��_���+%D���@EJ�4(���2�G���9b*%D���ȗ�V��ѻ���(�"D��`��;%�}�*�l<���1n?D���Q�_!t�,a���\���, �h D��&��#`�����&/(����>D�hya�ѡ>��ct�ػ,�X-�`�=D��svKr�� �����R0}��;D��+BH^�qZ0��u��u��`Tg4D����ӬF��P��D� 0���A��2D�� pݘN֠|�D�C��X%09R1�u"O�4ۖ%�5%<�#���/?l���"O&�
B�
N-
�3 �L*w5.�:F"Oj3� x����� BP�q�"ONM{��żW���F ]4b�Dö"O�SBH��� `�.���SW"O���2�Tn9S��S:
ո�"O�\�2��Z�\M8#��I�l�c�"O0�Ӗ�͆p�u�V���|.���"OF�:�ҟ`]���J�U�$/�!�$4�vUZ�l��9��c��-x.!�d�JDO�{&���O�(<w!�E�X���Y��y�.�:p!�Ĉ�eZh���L�T �!��o!��>8�b�!�4vz�@Į]2 h!���@BjajT�H�W��m�cڐ;P!�$̋\lH�b�)�8��у� 5!�$M3d�(��RHU�D���F��>y�!�$ңY�Q��%��T�\SG�!��Tҙ�����{� �ЃD�!���/T`�5�MѷO�bX;���>�!�D�CJS���8�~]���&�!��7��80�_�:	�W�8�!�d|-Ҩ�D�80Ҳ̊T�ܩ�!����Z�4����l��<��i�Tw!�$�P�f�JSi�>�4IKV�Q!�T�y�n=Z�I#Q��E@�J�!��ڭ!6���]l�0������!�DUɬ��؄Bsz��dN�H�!򄐭f��lB�B
�D�1�+��=!򤏴� � ���#�L�$�6/9!�d�Ux�I�4�Ӂm�#���!�фi��0/Ͱsc0�)��S�"!���@U:8�p`L���t
n�!��RTI-��ǀ3Y4�Yb��E�!�� 7Tb~<��j�*~��E,�1u\!��"�4�x�ȘN ���VMB,)!���}��섑K���g���!��TNj
�F���q��	�@!�T��	�%�W��z4 �CFo!�����	���%Z�d�3��!�$��}Ԍ�۶�[Ԯ�r�J(e�!��|�@99Q��q��s�)�1�!�d]�6&ĩ�`ܬf�b��QfD{9!��
\��A��G=�
tAGFG�(�!�dٔT��|��o�<!�x�YRDѯlM!�N�r[�X��� n��@�Z)G!�_��a��<�>E���!�d�X0a�'Ƌ`�˅�[�n�!򤁄4w����J��XqR���Py"�ߺIAȠ0hNN�`x{p����y"kּ3��|�c�X�G�BP	����y�XTXZ���Cl:,P Ś�y�A�z�J�S��gΨUr��S�y�#ѴC����πs��4{A`�y�O�1[��T{3.�l�2HJ�ڑ�y2��)���ĤXk�} � �y�g�)cJ\d[D��4��B�D��yB�*	Av�㮂���`&%:�yR��2�
��j��Xٺ�,���y�N�e H�Ń�rî8����y���G�$�6o;k5\ a���y"��+:��#�:Q����bH�y�C̊C��0�u��>Q q��A2�y
� 8��v�Ʈq7��qW��4f,Ъ�"OA;�jA$fHza��EV�xO�@�q"O�`�b�eN�6E��k3�A��"O��E`5~���F��k���q"O�jw@]50�`�כ��@bf"O�UB�׽p�H9P�C�04h��"O~��"N%|�l slN( J�+"O�
���^������Ii�YE"O X��O]H�@U!�J�v�H�"O`�p� �5?h�� 5Bɩ�\�R�"O0���ǁ[ۚ�c� �*�����"Oh"$�X�ﲸQ���|���%"O�a��$�q�'LX�I��Uȶ"OV��Ń�8l�J$��
_�r$�'�D"|O�� ��0u*��M��K{Ġ+�O��Ĉ�~>��i��Dٕ&X!}y!���U<�0��[: ��%�2.�!�D#���R%��G������6!�$���t�2��S�@Ԟ�h�"ʺ]�!��/lI�Uѐ^�ڬs�⇮n�!�d�2�˅�+l��c���z!����r�{��ύ=5�(�GJ-2!�V3&�
����T�� yW")F!���N(��
Δ"���#��H!�d��aҪI
C�+E�H���K�7r!��Z���*��	C�Ѱ@`��v"O��aEʐ(��	{��ɹ~Xfa�"O�	�	y����ĨMv�=K�"O��`1n�����-3�P G"O�����X4d��I���I�]r�"OxٳWe��"c�� ���E��9�%"OryI!
�g6^���IA8"���#T"O���Ǩ-B�V�KfL`�.4�V"O*tq�*Ҫc�"�r���@��H�"O��a�I�9d��As�cI��^̸�"O������!)�89'���6�\
"ON�JI�W�J ���v�$ɢ�"O���T �L)�4��l]>�0��v"Od�+RK��_����V
���Qc4"O.P8d��kN��g�_�4,�ЛP"O&�b����0�w���x 9
s"O�͓��K�Y��xKQ�Â0^�Yg"O�ĳ�D�kS�u�BG]zy�G"O^�:A�0S]&�QǻP4*��"O��t�͉}	�t���Q/����"O.���ì���A�>@A
�"O����,i|��a�+R
�A�"O���,�'P��)��٭H��a:�"O�1Kң��>m��J�OV0�HTI�"O��q�g��&�Z���U<6W��Z�"Opt��$]�5kb�J'.�=1|��"O.����E/X)�u��kv�L;�"O�AtO�.6Cr5s��:\�1"O�u�1�\~~���E�|8H�"O8!�$�ݬ.�De���a��Q`"O`+��O~n�����m�\� "O���p`������1� E�$"OjrR�y��@��C�0T�2�B&"O�t�g�J��P]Q���#�Ʊ�$"O|D�Q��ye�Ěg,�V5�Cq"OȀ�`��&7��8Ǩ7a.� 8�"OƐ��&��E�n�a�Xt!��"O*SU��$,� x��Ŭ�X�S"Ob)A'��g���
��d"O� �Zd���jTb4:�f��O`��S"O���C��^QT}{p��(��@q"O�����,'�Lu	!�P]�\��"O0AI�Y�VW0��K:��UX�"O����,|�j��TL	�!Vܫ�"Op���*�j9����!G�ш�"O
أ����U�V��A	C�X��e�"Ot3$�ЎD�ژ�w��/9���h�"O�\�aƜ<s'V�"*��t�\��"O�@���� Z*D���*s1V �"O�Pr0��!�ތ"o\4q9�xД"Or��%�?\̲ɹ��j'���"O �1�F�&Be�̛R��(#���&"O�xb�A��<n�� +<�	�"OfqS�>-��ePQH�m�щ�"OZ�Ӏ�.FXP6B�#3뎹�P"Ob����� ��q�d/��S�"O�}��± W<͚�O�R<�%P�"O�4�$f�m{h}��)�.<3�Ub"O�- v�$D�:���D�Aā�"O�A���-��%ֺ�ɂ�"O�Y�.�"?�9�D��uc���"O:�KB,Ͻ0ﾔ���<�<!�"OQS�.�(S�(��B�.蘠�"O��"$�}}0̸���l�8�"Oh�*B� �H���� 9fj��"O�qX�I	�~1*0��1`T� �6"O���d0d����K� H9r�bv"OhkCc� ;TT�fK�?���"O��C��c �C��և-��#�"O �[��
-�C�MN�Yl��p"O����2�l��Q���R^)��"OJ��5��,��T{�鈇A����"O��P'g����GjM!.��;g"O�A7�K�N�u�C ��<�42�"Ov����׫#��j�HM�7*b�"O�����L����-B-�"Op�aX�:��5j�[k�(�"OV��3�_�r�I��G�.^\���"O"�K ��(/����@M� 5�"�)�"O~�p &!0즡� Bc���"O��ÖL^�{�PA��!̝8nt��"O��R�! /o�6�!e P'-aZ�r�"OLX�����4-��*��H�F5z"O ���Q�!j����	�9l.L�"O�|��d�6�t�������*�"O,�Z7��c�����5�|lP�"O�qb2�ɱNM�W� {w]+�"OȡQ���1���a��FiZ�q�"O��(�nG:y�2<�W���fDيb"O��'�֗MJ��w�Q
]�s"O�4��-GĢ9sD&�#&�d�З"O,]@�*�3�l�#�D�~����"O2岐M�w���U��Љ�"O��XR�G�_}H완�	Xm4��"O`�y����nyȤ# BBh�9'"O��V�(N8�p�Ǳ*G���T"O����d�p8��
�ڨb*����"O6���D9-hAqm��p/�qs�"ONm�!�V����?�\�"O>�؂��4\K֨knkf���y��1�Bq�%/f���e �yb�ݑ��uhc�,��$�rc]<�y�! �A����+��TqťN9�y
� ��ۥ���hD���<uBv{&"O�}bt V�z� �{q�� '��"O�S��KJ(��nذ��,��"O�]	P'�q!2 ˲��9�|�R�"Opd��F��G��p��K&!".(A�"O����5 �hAb��S���6"OD�0gH17C��&�ުq���'"O�\�ݖ4F@�L?���"O \�+�?G�0Ԙb�ӆw�}R"OF<kQk\+^p�`3�&λ1r,JQ"OvԈCB[��`���~jjP��"O��'mJ<{��@@/�.Vh(��"O�Wb�U�4O@�Fqyz#"O��2���(EL Q@�]�D�����"O�m�D�Є(/�q�īŴ4��|QP"O8��	KV<� 	��z��%��"O���c��j��(I��[+_p���"O��Sv��:���&� ,`>aRd"O��IA@Ө>�bA��IUЍQ!"OB��?/:����i)*�zly�"O��7%�<}(&i�mն{���"OT��&AW��)a�+J<4,0�w"O��˕-�D�`�1�D��w ���y⬉J���@�AO�И� �$�y�oЊ$1�`F��6<�8�[�yb ��j���/	D��K��ϣ�yB�
��<VL�.@����#J��y��-�]Be��jh(C"�,�y����sd=B6KS�_kT��iY�y2fɺL�6��AM2_���҂��y�|���s$��U�8��ȋ��y2�Z 4�,ЈC� F�p���$H��y���
#�x��M�DX����)P�y���{��lZ�-lK�	"�(�'�F�����mƐVkħR�0��'���h�͐�	/�m�UoW;>t1r�'YL�+�E�jl����޳;�F�a�'���q�C&D���t˝�-����'zz`�5iU�ӎ9�v�گ5��	�'^^��*A�:��l��I�?]�Z�I	�'Ԯ�P� ��e�|��R���%3	�'y����݂�yr&^"��I�'7`y��&^�r�ZD��J�3�T,��'��}�".�1G����+��h1"�'�n���H�ZG��!{:�0q�'�]9�n�����L�[[H�ȓ�ZX��C�
R
8�  �G�83ڌ�ȓE�>\���)p�X�ˋ}����ȓ�\��*]�@Z<��oL�0cN��ȓA@����2\8�;w��'doN!�ȓ4^�����4]���
�?��܄�)�"}�0�Q�6@t�'�� ��5��Lʒ�G�
�mJ�8�1.��0G���ȓ �ؙ����6� )c��λ,#6��ȓ!�p�{N�i
�Y�:*����^�X"�ŘR�be�?B����2.�a��ӊ,����:O��$�ȓe �!0w
_P4��`�1�̆ȓ`�������8�2t/ح~��4\��H�%E��"\�SJ��F[���9 �r��ߒ}d\*��<�P��%��C#�ԍP��Q���9'����ȓw^ )�a��n��\����0T��ȓi�M�1j�;�z�x��	+!ꌇ�S�? ~�Q$�89� I����7��0QE"O�Q�$JN�a���!� K���A"Op��b�ꐕP o�$t�(��2"Ov�0��>BҰ��b�Z=k�Ѣ"O�t
@�GA�eI��R0�Bh�Q"O1[��)�|�S�d��b2�ɸe"O�ɒ3<���5$�HD8�2"O�0��A����g�SBB9�"O\}�A,�P	�%+!)4*�&"OPl	v�7���s�ԻFD���"O�X��F�e6`]�(��s2H�(d"O@�0���2:�PM�3環;�퉥"O(�j �� ��ǝ6��+@"O�l����@�Ua��l���"O�p�WL[���U���,�^A��"O��AD��(/+:�H��Z}�|E�F"O�af B�Arܝ�pbg���d"O�`�3d�z֩�w�1o3rQ� "O6$�����%WI�BBG�X��"OԘ	�(�bax����B�%%��a4"O�kУZ��AE��\x��b'"OV�c��0>+@�pt:M]<��"Oơ�c��H���g�%eM�|��"O�p���L�q!%DKO&��kP"O��sǡ
VeJ��/�|�&"O��6�0Mg�Ya�	�d�B�P"O^0���ip6ٸ%@�U<�� �"O|}c@Ā<'MT�!PO�O$�3!"Or�x��L(8z��E��173͓"OP���@=��tP!m�(3�!C"O��BQGB*3%M4�9�"O��!���n�Tp��(z!�,y"O���a,�|�$���`��ye��a�"O ���-Ѹ#n��/��+�đ��"O�؀g΂�#��#�̆z5�,��"O�ex4
�;{�dݢ��>w�L��"O�`H�P�J����?WnP! �	Rx�p2��������`�R����7�&D�����D3[F��c�f�f��1b�?D�X��Xwc�]�Bf+[$�c�J2D�Hצ��vv��⏃�O�b<x 0D����
JuZ��;f.�'�T�1D���6�ɘ9�,���AZ� ����$D��s�D�mؘ���*L����"D��9%F�EpJT��'^�R����sM=D�<bW�1j��Р��|����CC;D�4�! ���Ͱ�m��o����4D�����2zP�`��,uC��[#�0D��0� � �i���TޮA).D�p�I���1�W�¹+l� !�7T�T��dтn�`I�(?���"Oڼp"`TR"RT��N#Y�q�7"O��5LB�����­�� (�@��"Ovt�B+\ft�ȃRv+R�n D��h0$	%e{���4@��w�����"D��Q'�X�Mj�ˮb�J@�M!D���S�L9 D$�	����P|:����=D�|���O�S#�%��犚iV0��G :D��;5�B��i�d��,�6/6D��BRK�	Sz�k�kH6&���2�`2D���
�>�9v��q��VN3D��iP`��������o��d�4-D��;���7<�0����o���B*D� �u/
�{PX�(��ڧgs��g�'D�� �J�B�~�j����o)��"O& S0��9i��}�&I�)c��h�"OX��"�Ԇ�9X �� Xr�z"O��sCkS�{9d�8ǧ^�
VB|B��'��O�m#jC�Z>�T@4d�.8�LZ�"ODPbK�(N-N�����e�\�	f"Oj�Ü�c
,�Ϭs���c"O�|@���=u��Y2�S��f4j��'Aў�ȑA�.%���r��[���c(D�i�&ɮ�i���M.�"y�5�'D�H��.L;a�� $�Z�Z���@)�Ob扫i��2iN�|�Ad�<��B�I�iP���=Aᐍ��fʩa��C�7W����7J�����.Y_�C䉎K��)C �I!�Q�.y��C�ɮE���x�(g$B��!F"vf�B�	M�f,"��e�w��r.*C䉤�����_����S�g+�VB�I2V}�`���IJ�e��ݚAK8B�	�!HD���0wh�cq��{?�C�I��F�C���<�c�Z�EnzC�I�D@��pG�.3p�2��k�vC�V���C4�_)h�XQ�iY )�xB�'��u��/t�X���@�6��C��0n@	!ةdn���+4&�C�	79�����	˄^�vU
2�׶}4^C䉤_	x%��EC	8@�qgΐ)@vB䉄Va��	-/ ��� |�C�I'o��I�R� *�*T�C�I�i�!5�@���Z��S�JC�ɸ$`j�;���]a��W��3
~B䉗a<H	�H@�5�.ǙYzTB�	�z��!����?���zT"�f��C�	�N��e�0jb4�W.ԮR��C�I�6��s-�L��qB�!+ytC�I=;G&���%P<S�&e0��9�dC��#)>r�1fF�4V��{�Gϣ]<C�	r���5!�dxW�	�-� B�I�G�D-�BA<,��wL�$m�C�	  ׀���kG:|��f��2m�C�	�n]�����
*G(ٛF��m�C�	�F��IUD�cR�d���	���C�		L���x���B���l�B�C�	�L�D=!4�6S�����Þ�1	�C䉾;���R�͌L�)3�+C�BB�	�{f��)��Oj���@�B�2B�m��e���0�pɒ���&B�$�F�%]�I�nKY�B�	�-���3�@ю$s谒t�G$V�B��3���c���Jr	����PU�C�	f�"xf�5:�! �̓n|�C�		lЕ�'��a�ŉ�5|*�C��yYP�����+=��(���1:�����u�@�C�e�s��]�t�&�!��e������^�xAz�A��!�䎘p�J)b	L�G�X	��a�!�$�?B|0�葟u��U7p}�"O�!L�?"����D�k���"OP�ِ� �5�zL�劝3`_���"O(t(�"�N20���ݸz�\i��"O���KT��:��t���%���aA"Oh0K���+IN��褧�+�H�"O�z�Hƫ/����L[�5tԺ�"Obt�3	J�
��T.xhj�"O� ��;bh���h���m/p�(2"Op{�Ř"�5r#oA�&6���"O����ۦ�e+�nG�_�Z1� "O��x� ķ7�*psD.?i��ؚq"O���mܰ"<�}yÌ�Q?�m��"O��ʡl�PYN��ՀHX-��"O"8��ð$ײ�B���$BX�"O�x��ĕP��ˁ�/� h� "OL52� �t�P镘`��L��"Or8�FݍD㤁�G�, �
�#"O��ۦ��MfR�3ʗp�҈{!"Od�ВL��rh8I�e­tb�S�"O|:S8<k�9y�"77�1CD"O����jip�y1��B8 �ס�y���L\��!3-�!V�VcW�Q��yBŒ�+#3kٻ8�0��!�yr�?j��y�F��+qh�)�-^��y"瘠,y��1p'��̢)V��7�y����[=rٳg�G�@D��U����y��Z���DKĽ5�!dA��y�:,�"���J�
t�BC��%�yR�^:������ r9h�M��yrÕ�B�|�*Tn8e b��K�0�y�G�n+����]�_3��%nǌ�y��F�22D�I.X�d��B��y"�7g��j$��QŶ���N�yB(�o%^�3a�2���4��y�d��`�q��	2	��#G'׏�yR��?����C�RC������yRVcyd h��7U��J�(�y��;��#֮A�G�%:���)�y��ƽ	+��j�AE�472!�cW��y"N�8Qf�@�^�x80L�O�8�y"GL�pu�}�%��l��5�u���y��c
�h�j�f���K���/�y�Br��ɺ��,c��{�˒��y��|��P� V�#"�xTg�6�y2�^�0�	�0��H�8d9�3�y�쐜���3mJ�i��Y(�d\��yr����T��$�+]���c���yb���)�"�U"�p��C��y�,C#?L"��g�Y�%rUC�F���y�?X�!�Է�*�ʕۆ�y"hR�x6��@��(���׷�y�b
-U��5��jM2�F�
���4�y�(�+r�(+��w�PTy���y��>:��{�'�;z]�1��&�2�y"��1Z&H���;	{fE������yR�ՌU�D����-��%�Ч¥�y2.�K�RaN>�E���yr��*=���iP�ȡ|������E6�y"C�# :|L8��3��%����yB�$o�؉���.K7(
�&K6�y�ŘZfrТ��n�h	;�<�y���I6V�3�bE�B�)��P��y�j�rCv|ˁ�� �Usu���y"�@��4���� �xs���&�y"A�$$pD)���2LH=@q��	�y�*�7��( ��ʙ�(P��&I��yb�ޥ>��Q4.P�2r<�XB��y�	Ǯu��!3w��<\>�Za(	��y2��
G�4����)l�����&
�y2H��k�<X3%�//ʕ�Q)X��y�)UQ��`����䈊��y
� ��:�@�,v�`�w�1y��Y%"O���m�7V��[Ս�n���"O����}R<k�_�D	����"Op
��-�6�X`�X%�`Q�a"O�Y�����w��}`T�@&�ޡ2"O- bN�B���I�ʑ��1�"O�hCH��S�9�B�)>��)IG"O���G�è_�����TN��XF"Ob�i���t�*��v�����i�"O��a-����HG�)q4(�ӂ"Ö
4��O��-��#ƭ��9��"Oxqzdc�:o�h؅�
�u�6���"O�𹄥>%\�A�"�#
?YS�"O$�xe,9-� U�c�}(�j�"O.�a�
��9z�Y�p&i�"OP@��B�4|A^��1��J���`"O��I��͊`v��`s`��=�4�""O^��񊝦����!��ڡ"O�@�����g�tđ�Y����u"OB��DH&c�֨�(F)TG.��a"O��Z�)�wl�)&��V,�MK�"O�E�e$�-xp��w�V)?��"O�E8�
S;*t��L�3[|� `"O�̃$#ʷ��	�$""OHx�u"O�E��.�Y'F�E[�9DD��"O"�w��|8,y16�B�W���`"O��Br�F����t�&5j4"O�\��'f���"�c������"O2H�#敱,L&�����f���
�"O|;��	���8#��*+��`a"O(�J�ސ`ZXw-��0�N]�A"OP	�7%^`�a��[G�� ; "Or4R�*�'_��L+Q$T�8�0EKP"OrLB���7��А�L�#:��0��"O�!��_�x$6p# �)
v��@"O�l:��H"�����J e^�p�"Oȴ�f�k���1����/戤�u"O�u��k�y�>���?Kj�Y��"O�XwbY$s!�E	R�J�NT����"OjR O�EHEY�vE��"O�� �b�PlXmۖQ0��p�"O�xa���%�Qc/͉d� j`"OT�I�/��o]��TC^@�lmC�"O^��ciϖ�B@�#�S&"O8�1c�˿/����`��"�"@!�"O��kp�КƎ��/1��P�"OHD���
J�����U#`� ��"O�I@6Q�.�x�	0,ԊUy�"O�h&�سBZ2d�FÞ���{�"O"�:��ׅu��X5�] �,B�	A�j)X�LTe��RՁ��%�B�	"M���*G/@ vG���.(F�C�I�y���q ��s�l�Ó��ei�C䉐8d���b\.�aj!5٦C�	;.("e;g�� ׈D2sm�N�rC�I���!�Ѣ�/|�d<�Q�0O$�C�	Gn( �BVL.xZ ��E�C�ɉw���5��6l����A���B�:_ɂM�6Ώa�YP7��'c�B��C�n9��ɝD2�K�ᎇm�B�ɰ撐*�k�4D�h�&�N�vB䉬R��ls�/�+^��/K���C�v>0�Z�IN|2ވ��r�NB�I�J]���'^����Ă$&
fC�)� �8���<=��+��*3��|�!"O*��G�1+H3&�
0~���"O�� �$��Yh�w�.E�$e"OR]h�LڭJ��I��kTx�C"O e��;?v�4�F��� #~�r"OLX�$�U�~FH���JB7/�Hr"O.�i�	�>n=��ڱL�>ab2Ձ�"O��i�-5e�<i��� ��MY�"O�ٸ��F��t�6�
�:��H"O@- g�S�!7���T�E�0+��S�"O&�A0�-%�neZE.�!v��a"O��*&�]��D "�m�\��"O�!Sq�@�# \,�_oh���"O�yV�K1vp���m�?����"O^�{�ƕ l��v�J:a�Y8"OV���]xd��G�%�f�W"OVp�h8h �7ωT�(!��"O���"� :shևj$z]y�"O��Z��W�Tڊ��'-{�y��"OАZQ�U��"�2��4v�ȸ�"OH�T���mF��������1"O��U$_%"�i;������ A"O�tX��6)g�:EMľn�F-��"O�5p�h�|�*ȰR�֥n�@�@"O:�{�EQ�K��I	v��,t���"Oh��c@��:%�5OΜr\$��"O�]{gd,g����/��L
"O�s��؁:$l�-,`���"O���SnB�� ��<P��Q"O ���揅\�XQtB
Tbe�"O��X���X]����
�qCQ�"Oz���ϫ(�x���� rѴ̫�"O&h���5�"��g�%�a�'"ORL2&�Y���j��G�1L5�@"O�Dc@ �o�h�Ӆ���p|��"ORA4�L�?��B��)���"OT��1N�eɰ4bĴB��02"O����a�^����D.sW �Q"Oر@��ʀ2z������`b"O��Hȁ#���:��K:J91�"O
ty��J��10rmI�9վ��1"O]9g��$V�U���	,�&��v"O�L���g@n%���=gc��9P"O��b�e�m���R�G��ӑ"OF쫡��w%�X��IC�ȩ�"O���EE�;>���nN�NlR��E"O�q�e"n�R���էv���d"O�l0$Ȇ�6�h��G,Ф5�d��"O����IA&p�!SW�0o�:M�5"O���d��?S�4�7��{��Q!��4"!�͠�Iэ�qiuj�D�!�Ğ.6�(�(RAµ}�vRF]@c"O�A��냤m
�qS��%="VH{"Of|��!�?6�]S�g���j "O`�x`� 
��[Rf�*s���b"OXx"���C̼1��AG�f��u"O���H�/e3n��S�+a0� "Ol��h�(}L�� �o�0|�"O�ШE�	��� ���2\��i�"O&JCV(
Db��'PA�5"O�U9�E��/������7V1��"O6L�"�_�0�2d=t�`�"O� "�I	���2@	�w�����"O�y���]6ȥ���<p[��@"O� �Lk�� f�ʠCD�1T�u:�"O�%0ck�݀(��n�:��PC"O~�{4,�8O4E(p,� C�"OM��/B ����A�V)W���3!"O�Ź�!���,�k��'�ث5"O�)2��roF�D�V�� )"O�0Y���\�I�ÆϺ+��
#"O��J`k���!�#P2B�̉�B"O^��J�}a B�Z���٢"O����$�"\?���ä(����"O�\��cϻ$���;�
&n��9��"O|�y6��E�HhшҐ	s e
�"O���N�r�@���.����"O\�A�גV�t=P��|��TR"Of%�5!א:,�Qbf���TS�"O���Ǆ1E"�8Ⰹ��P��"O2����Z�0�y����M�&yD"Omw��ED0�� d
#.��"O�R��|2�!壆���(�"O@@�c�r��A���O���z "O��z��ͫ`zoܠ-\���"Oj�	EZ�_4��W�ڗ����b"O�y���+&��k��1����'"O`����V�33�q�k��g+l�!"O�Q�sJLDE̸ ��B&<��"O�)p�BV�y����gЉ%Y�8*�"On�i�AM�X�M@FgS�(pn�t"O�\:r��]G`�����9��U�0"O��	��l��9��a��)3�"O�i2C�s���с�	��A�"O4��o&h��qXs![[m�g"O�	�Tn�9��A(��Z�q��٢@"O�!���
g!��[�� �.�"O��s̜:�t�Y�X�v[�"O���M%fP�A�2�� E"O4���`ϙI���IG�£s��I�""OƼ�'��,��r���j~�5`f"O�8*Q���0�$ݪc�=�6���"OPЋ�BBTa�񊐃uܰ���"O�����9#52pj�
ڐ�q�"OD�1�+��K	��Td����"O&���H�]���`��3���q4"O�d@���p#�U�擉J��p7"O
��b��u?2�!��@�n,� �"O m�F@#L�
��Ş:H��2"O*u��!B /�"4a��ϗ5G���"O(N 0�����J/~���E"O�M��Hz�a�W��i8P�$"O�$�F	�mW�@��뇲r ��y�"O*�x�F��G� ��OK�D����g"O(�3���|E�M�7��4G,�cf"O~�yg�D�w��(6��$O/�q�"OJ��% �USv5Y�%ՃKXa"O�A�Wg�:6�d�qD?.�"O���LE:\X.H�Š˹\x�s�"O$��G04��a�+ �<i�"On�!��ֆ$fhx0`�\�\��"O�(�f� 5��!E�˱F�h8B"O
�r���+GP���ܸb���Q"Obͫ���?bDpdr�տi3�0�"OVhc0g��#����M'�1��"O�,��oH$㒙3!�_�!&��U"O�]2rjۅ9V �g��k��$&"OX�!��&�x�B'<����P"O� �uIǮզgE<�S耼=gX=S�"O��3�̀^�DZ�KL>M��"O
P�r�]�Q+4�����{E�`��"On��2�İ$�h�f-�Ĳ "O��˗����ȓ�S"8jV"O��p6�ȍK.j�"�'	�X���"O�u���)���3��;5)8���"O<�`��j�̸!A�����"OZ\Ӕ`�Pv��jW�ʭ3i�HZ@"O:�$Aͪl �q��Ŏ�2\���"O�����
�n�d��0���g"O����n���%ذ���4ћP"O>E�1�C��e��	E6�fm
�"O��Tc�*2�~"r�]��0"O�ЙA>@Gp꒩$M�T01�"OZq1�+�P��Q#�Y[����d"Or��&�������C4t��|�1"Oq	D�CU�
����22��	Y�"O��KD�K�����͓�V��"Ofax�FQ�L6�ɋ��O��,�"Oa �Q�9�!��٥/��msC"OB��"��� ������h���"O��{��2I���h!M�� Q&�c"OZ�dk�7e�t�����5)
��"O�)�e���?4.�ţ�;i���a"O�k�.Dt���@'��K�"Onic�K-�&=��(����"Od0��薟7j���$"�����"O@ݡA��.|�n�I@	\s�,Jf"Op��)�=��:� �hL��"OQ����m��Rv���X�h�V"Of6��ySj��C�K�ieB�S	/D�����p"�!ɜ�D�S�.D��x�o?�M��ϳ��� �W�<iF�~u"��)�� C��_�<�!w��@�3 �W�i�Y�<I��Z4��u��D�" ����l�R�<A7)�0�X�#L�c5���r�TM�<�E*���%,�E?��c��c�<aǋʝX�LY���k[jiY��a�<Y0�aE� � �-Gh^���`2T�K@nP;E�%�fn(�����"-D��zP!�	O�=��&��1�8B��6D��P�J@�g��tI�J�4�r����&D�8r���WR�`�P+�0X���� #D�p���]@�DD��l}��� D��)dn�2/l0� P�"�h๢a?D��d�|?p$�aE\F��3>D��ˇ@��;�tQ�+@��!j'D����O9>�d�; �H���C0n8D��0��W5,��B�S���<�� D��yR	��G}�l���\M0�b��>T��׉��JJm�ƦU's�x��"O�{P�U%3i�-;��P��<�"O�d���G��ك �^
F�t��g"O�5�qD�!H�%Q���<~����"OF��P�I_���sriW91�|�"O��	UdYX�N�H3n�1~n��0"O�P�� G
�qz��d��iS�"O$q�c�2r���q�U�i��H�0"O��&����n�C!�O~:���"O6�Q�L"J��9+���EЀ�r"O��Hd���4�J �	Ͳ}+$��"O�t:qBR��P���6��M(�"O� ,�j�0gV�A�A BDX�r�"OFy�f��{j���	˄Y0���"O��"Q���v$ �)�2$F��"O��%�M��0]@�Ȗ Y�(���"Ot%�☐P��v�1<�@q!�"O��`�N޻	��c�$ۜuYA�"O����K
	Fh��#B*gQx(�f"O�c$O�&����ab�.RL���"O�yJ��*D��I�oR@��b�"O�<	 ������d2�İ2"O�Űa�>7p��إ�V�.!&��T"Oȍ���I�t�rl�����t"O"q�V�شr�4pf�:?1���!"Onд��!�����2���"O��/�#���r>���� "O��XfB��H�^��l_�%V����"Oxe�����KP����IR�L��=��"O�u�Ĭ9ιCbiU��(Y��"O��"fO�rKn) R.�R0��"O`��Ӟ)vihu�#�8�xv"Oִ���@45��e۵��>w�\˗"O���T�M(hZh�A�=�4�"O��5A����cc��*���r"O���/U�RD�%�H�pC"O��8"� q���y0Fث.�kb"O���A�H�d)�p�'y����"O�%���@,xB��`*ܷa�L�z�"O��`hǛ+~�QI+F�1�q"O�d��C�b4��逧\=F��,�yҪ	K�@�h�"ߤ=�6�J���y�S�[�XÅ��5�&42E$��y���v�I��K�#&�	+����yҡ�]�(�B��h��KQ���y�	л\q��)6 ]mb +4���yR&P+m�Iz��gY��S�N�yb���(0��'�̯Y���R�OЎ�y��bn��Ɇ!�F��%�2`��y"�W0e�}���� T�.�ق���yrjr&�� ݏEHR�"�%�/�yr�)F�nM��G<�.٣���y2ɔn�ޘ�$�7�X@�M^��y"J��p�J� ��*\��MƂ�y��wъ���SI���R�A��y�%��E�$���]?P���q�&��yRBټ8V���Ê�C�^<���Q �ybC��8}PiR���,Lˀ/�;�yR�F�d>I+��ɇLH�j��	��yr�֕b��Pf헔�4,[�!��yBFҥf��q�W��Z�ƽP%�=�y�OR���ybf *}98K�G �y�DVi��Hb0d�,��w��0�y"���7�*ɂ�������&�yb���t��Tiì�v����Ă�y�����i�.�J�beV9�y��\�h��d��(*Ph��y�'��vo�m����T*$)�(G/�y�#-z����vg�й�lƩ�y�E��V�z�r�+�e?T@�w	��y��;�J$Hd�\�S /��yRK&n^J욱�Y7h�hP�ץĭ�y�GT�TD���D���	W��y���8f���T��7q;�U��y�,�gyp)���3�P�����y���j��}3��j��Ѻ�)��y
� �t!��ԗ'�>�ǂ�'�v���"O
�+�F	�2І��^9?��pp"OhA��_-�[���)�Xp15"O��;BAU�QB#?&ܡjA"O���G.K�[s�Bë��j��R"O�h�f� �<p��d�E�&"O��vf���7�G?epl�{C"O��@��Dx
ls���%3F\��"ODPZ��U'(����b4As�Y�"O`Q��\<��@"5�ҥs�hz�"O��y!].jH�Sd��;8�B6"O| v�Ć%о����T�m�Tӱ"Oi�ፙ���b��RyX}1�"O@u��$O/$�|B�C�-SHda�"O�=@saֈ1F=�&�ͣ`<�es"O�ы�D�J|�P*$��E,z�s"O��b#j����iN�#��X�"O��YB�A!7�`� $�Nt)k�"O�� Т�(3Ӏ�AŞ`�6|8"O�IRa%5trx�`��+[����"OR�KW�*fV|��bøA�Jq�3"O��"��|�T-�3�yu.]��"O6u����m<��2� �z�����"O���aDS'>Y�/Y;q�
As"O&T���;�e�޴֬�x�"O~�s�Xaܐ��7/�,(�j�""O`!��nF"9�J9�D �_|�$�""O���NK���W�,'n��!"O@@sS�CZ��a�\fBt`"Oru���fRL��K�F]�$�"O�yʲ�ލ��5��S/X��p�5"Of���@ʖJ$��8T�E�.�|p�"O��P0 -B�r�Hu�ť'L�� w"O칉D掵Q�:yz@j׶+��S"O���f@=_ԴĀ�/�m"�"O�Xh�#^�Y�|Ӄ�S6a�Ni�s"O(��1�Ç1���tFβ'����"O,9�РZи���\�*�`�"O�Yq'�S�f^y��%S�
����"Oh�x�d�4y�6��/����R"Oha귢G�C�t�� +��<X��"O�ܪ�G6}6@���*��p�"O&���`�  ��m(���8ai�<Z�"O���iB�>��Qe,țS|p��"OัC���7��p�",�&ZM�`"O:|yU�D��1
ڡ<�:�{"O2�r+��xp��coS�Tޮ�p�"O<U ��{��U.�+Y���9�"Or)�BIF�NT�5�AL�դ̒�"O���A͠>�x������$A�"O�E*����]v�@�\�&�B"O�a�E� ��b@�ox ��c"O�H���k�)@b�Mk��S�"O̍���Z#4p`�!*"��jD"OB̳ �ƦD��)ɦB2��ݹ�"O�=c�'TY��0���I�ę2"O�8�u(�!6A�D�ĕ|lb�y7"O�$��!I�{�I����	��"O��W�Ţ`��Ё��ܱ�'"O�a	��Om̌@s�O�!�
�3""Oĕ��nP�p����P�H�do&eQ�"O>a�1����\�82��#a"O�h�GN�Q�<0e�;l'lDA5"O��ɡ��
��42�����2�"O� ��0�k:=��!�/Ѽ,[6��"O,TP�!��l�6<"�@�<KS91"Od\jw�A�'0�DoI��ұ{�"O�qB�=��,�Ӎu�ȑ�"O��!��C�W�����S��)�"O�E�ϋ�o���#�GX/E�l��"Ot�Qŉ�3C�A�Aɚ,\�`,#�"O�\�h3�đeʐ�!����*O�XA�αB=�\j3�
�j���	�'�HxWNB�y���D��i�<�'�Gl�7yz�C81�~ (�'ņ4��J�<EB8���Y�V�x�k�'��sq�N�p,�Ipm�OX���'@:��ר���,cf��3}����'�X;3B�2f�l�կ�}Wn���'m*}�&��1��ˁp�Ma�'-!��F<lw�$S�j
�Q.��'�DP�b_���E�Pl��'�D����㊱#�<�|$��'l��!"]���(A��ԑ^1����'��$�t�ʡu�>��䛏U���0�'J�iQ����7�r���QSwܸ��'�>�:����աq�uQ��R�'�25��dA?���@ıg思��'(�qS�n	> ��"�2����'�x��$�Yu8e�_�bm>�b�'��u��΁�F��4�<(���'}��j��ٶ^�(���> ��i��'�$q��oJιe��n/�P��'�����&�U�DAº1��S�'���h˃9-j]:� �4���;�'��ĺ��$j�L`�S�K�.zM�
�'��X�'텶W��22/<"�ё
�'>�ek��ٟd~�P�	J�!Wl 
�'���j�*Z�N!r�ۆ�[��r� 	�' �Q'l��9�iv�Q5H	�'x�\ڔ͈^��86��d���	�'���Q�E��Q`td+��B�g�����'{�	Hș�3�jTSS��_��ر�'��"�'H�E�t@�2��6X�@�s
�'�6��3DөKN�����0Y�l��
�'�D� �Wa���Rdj	<g�p�H�'o@���ɉ�a��4FM+	>���'�6�J"h��̈�g�|zԜ��'b�IU힝8����e�sǼM��'�J薁L��Ndy��e�*�b�'��K�a�<v�^i�ʉc� ���'nRH����%�,q� +M�E6f���'��8�Di���@Հ���&�����'����QO%Ӛ��AA�sH�D��'
���I_��*=�Pi��S���'-�hXL*l9�)�EkD1��'�t!�AGC4�ZY��8BQ:��'��(��L	p��Y���Dd�s�'�H�WcCJ}F(��ժ	��$��'6xq4灦
�r�:U�N� �戇�iB�|5�qT���� z Y�ȓ{�� b��Q�|���ֹ���ȓ��9A�E�x	g{��m��U0&	�a%^�wz*uI��W�gSr��ȓ���&H
�2!Lh���Ohw���ȓ^y,p1"K�3٘�Z��7C�ti��Nl�]�'TE�6Ez0�C�$��d��Y�!��eޟ7����@K�YfV���S�? Z���%V"o~ph`F�� + ��"O�1���4t�<�Y�|��9�"OH\g��w��C�똻,�P�j�"Ob1�T��j%<�kf*�(�Q�"O�mz��ͅsG�h��אI�H�3"O�!���&E��0��§*�b�"O��x�7?;�̉�H��JL*;�"O�)4�U�k\�t�ġ09dZ�"O|�	�e^�2'-SEA��S���0"OlT���<k�1�O�3��qBR"Ox���\�4���@�E)t��t"OJaa��ҹoБ��ϐ_;̌�"O����G��W�V�Ka�1�R���*O^X�	��*2��s�/R4��'C�m�l���-r��C	4�@�'�:ٛ�A�.�܈p��5�$M��'��Ȑ��	?|��7獞a�ʤ�
�'�@`PQ%� c4��c֡�?ZƊ�I�'(Z��A̗P�<�{"��Wg0(
�'�(!->��0���e2���'68���Y�� ��̲^c�H��'Z��t(�/$,���h� �=3�'ݼdڕOIZH�pF�հB�y�'��ᙰ	8cJ�[6ЈJ-����'fΌ�� �|�&q u �A���'������F�;	��`��-3D�l0���m7^c�.L@f��s!%D�����S�[T��B.���m�c�7D�$2 �H�@Q��Wi�=� ����/D��0���3j�!+����O��%��J8D���@E�(&��8���Qn)D�\�&�Z6f�4T��k�4�ڣn4D��Xci�O��Ȉg#8���+�	>D��	�Y-y��h&hOWZ����7D�t�q&�&hи���,L�\��'D�h����M �<��N������&D������S�>�ӕnN��-�b?D� ڃ�RL@H�F��&���)��=D�����^[�:��e�s1��zCK:D�X{3��,@�,	WiݍI0�M� �<D�$����-4��eM��EB�uH$'D�$6�Q�l�r���L5��q!d%D�L t�ǃ��T�@@�,Kt�wA%D��Č�?.�\�Z�F��O�t0��#D�<Ktb��4����ET'̴`v�"D�ؗ�NN����Ͷ٨ ��3D�#��+~� �(��O�vXW�1D�W���G�ɩ�n
�/J�i� *D��0e뗦�lI�`܇En��t�#D�����)<�2��]���� D��uAE)u��� m�6<p�>D� �MP<T`Hai4��Y���M:D���6B� O���I����:�l=D�@�k��D\`y)�nU�c+���w*<D��ze�״�s�ƈ2����3F=D��`P ލh�6=�@Ò��:(�e)/D��@�/�S�5Pd`â!i`��"D��Bp��a0(���]�gL;D�D
�,A�[Nv��lھ<���aB+-D�h���a><�Ss!Z%
���:��7D����x�\��`�vr�lHE*O�5��MKX��h8�m�8{\f��"O�ă7�ڀ!	N��PL#f�]
D"O��E�ˉ`7��Y7���b�26"O� ����k��W������{�D�rG"O �{3L�~�0D��$_�H{ԑ�"O�(23K�%I2���pIN*9z&E1�"O�m�&l�x:r��E�� yv ��"O a�$j򄄪��s��ht"O4ᣁ��U� 4�G����&"O8H�"\y	�`�G �!ް��"O�D�-��a�R�މ?�`UH "O��Hő�p��ǚ>af$��"O�e�5�սU��@��H�5�m} �"O p��o�Zy�3�+:�T0R"O��R��[�(	����*�Y�C"O4�q4��3<|y��W)���A"O`)�)U�-"�Y��/[��,`�"O2��WE��L|]�䮆�
T��d"O�q21^�VT
�l
0��*A"OT�dCH�A%R���N!u�Bܣ�"O��Q�"9Mx�z��_g� |��"O�,p��N
o$\:�g�ͼ���"O5���
Dis����-(�!@"O"����ۦ"zJ$���l|���"O@)S��u��m
$�-c�T��b"O�&N�E}nL�d�g�\]��"O^щ��I��p�X%^b���"OށрB͐B�^��3��4�h�G"O�t�&'�FB�X�$��@S.:"O�����/(����k�<N ��s"O*s"�-ՠ���k��yI�\��"O�1���N�=Ȑ"6��4Er}I�"O8��U�2׌�R��ϙE�\8Q"O��0P� �5|0��f�I����"OМ�B�t�(L"U�؟)�5Y�"O�P�Di�:V�*��bk�p8��"OLBt	�(M���І���Qv"O�š�����&E��
<Jw"O���D-��������9`�"O�����Ƭ6d��bB�E�V�t�T"O6�2BV4����Q��kPj�"Ohl�CL�T�y�R�_�a��2�"O<����)n��2oʷ���@�"O��[Tj^KTv��/�-�j���"OJ�B�\�Y*0�z���
&�÷"O|����9Z��{�Mfj a[�"O$� A�R.*�
<�3L��`7$k�"O
x����p$�U�Q�����"O��� 1� Q��K$gk��ɳ"O8c�τ�k�N`(�$Ϣ0Ȗ�0"O�R�oJ]xX1�RLJVV"O�@�c&ܭS�a��}?��Q"O�Q�����R�x���D<t]�u��"Od �M.1>�i���H,���"O�0"��Y�'��a�>]L���"OB5��N�8#"�$Xt"ݘ�k�"O��[��ŔpJ*P@�@ǽT�� �"O��9��������H΁N�ڱy""OY �K�)�Cǜ�E�,��Q"OdE3 �iˬ-�D�B��iw"OT��4��7*�L�1Dωi�l�z"O�9�J�'�$�t�M6�&��"O����B�nP0�#ùV�� �"OH9��)�b�f��AǓB���""O��{���}���V�A[2��"Ohx��X?������F=�9��"O���щ?[� %җcM+$P��'"O� p��쑊yы�BHd)�AB@"O���cA�3+�<D�ɱ�!��"O� �N��Vج�v`R/��"O���D�ջEd�m�ҠR!.=�1"O��д� �-yj$[�X$�B�"O�-����d�j��yTH��"O~�Ƨ��p=�l�'�DD�҄"OV���뎒���!f��~��"O��`	5����RDɐm�L��"Oh�3Q��_��L0�DLa���a�"OH�3�I\0Y-L0�Ճ�/O����"OB5�c�^<ZLרma"OL���˱ky��p�Lت?eܥ�"OL�*�ퟶ���q���.[Q����"OT%��k�;f%T��#�> ���e"O�UZ�?B`X��_�4����t"O|ijagJ	����^�yV\�"O=XA�I�a�n�y���T�!�"O�Xs��J$=���Xq+P=A��"O��&��,m�<D�kШ��4�w"OT�e�5�&��q��Q��M�q"O����t���cF�pk&��"OJ�"#�p���1�� ^�A��"O��C��nR��c���5_��u{�"O���OSF*�tJ���.*f(��"O)`d���e�P|!冲>�K�"OR�!�ǅ�:a#$��L�b�U"O�&��,�-Sf�3v��d"O�x��">���p��[o�T4"O@5P��G��ؒED�<k8��"O~��q���;T��O��S`b!�"O�����,I��$�3���q�r��6"O
D;������h�MD����"R"O>�H��/K�HDb
L�bz&"O6�;ե^e���&	c|@q`�"O�}�գ�`���D傕cE���p"O�X��)"O4i)�	�"B0�+�"O��Yta@�BhXbu(ۨ|)
�J�"Ox-�1�ѹG�H��'[�\�����"OR(£��k��E�!�	�3���A"O(��D�;r��}�`�D�x��W"OBTBǓ1�Ve	��58{p!"O�� 2��d�{��7l����"O�5��n &2Y���B�:9��"OBh��	�:f "���M.��c�"O�	ˤ
�!_���(�/��+�4I�"O�`�.����𨎢RnHxg"O��0N	5o����s��r"Ox����*Vn��BU�;����"O@�je"6.��QAs���&\�Q"Op`b��(V�0��V�nަ{ "O*e4$A%X��I�j�Kh^,P�"O��G�M֤��\-�̥*�"O(i�����-���&�ԥ&�,J"O����@G�N���0�AN�
�Ą	�"O���Μ���!��U�b��"On�:̈́���h�)��[��0"O�m���#H06lZ#N�p޼�@�"O����ML&HY����[ܞ@�g"OP�h�D�W��fh�n־��"O��@u"�)�6��m�5�		q"O� ����:p\�y��(�PF"O&8Ј�,ԛ2K�'6�����"Ou)`�C�M΄�2g���nIB"O� J8{@��y�8,��БBw�L�5"O�Y�Q�!>����� vl���"O��������0"�G�rMf�1"O��PaƎ[)�C3��g��$j�"O.t(D̄?\�^d�/�:��ء�"O�����
t�p����:��H��"O<��օݸ:�nPx�nץ;�HR"O�3$ʒ�j�2 ��NZ�#�-H�"OJ��i��@�.�#�-�0s�t��"O*���O 4�R��ɾP��D��"Oak�D*B#tݢ�`�$[���س"OT)��Ŏ4�܌�p@ܗ:m.�"O�,@��,]{p�(�\|�N �"O~e�f�X
o@՘w��;Жs�"Oʨٓ�M���!��.�$;�B]b"O�[7�^�qx��Y�6�\��"O�$�1��6�����4]��"OL�a7cI� ���$Q�p��G"O ���ȻXZ�8 ��Z��#�"O��:Bm���~�+��3s�q+e"O��cA<q��d�f�ϟ]�l�J�"O>t!#�L*�d�s�,D�X�jly"O�m(�J�t��u웱L�D-�"Op�A��P�r���+L'jE�ua�"O��e�Rb��ak
�ׄ�T�<�䞘(�\�!�䌩@�<� HV�<1qE��o��`�+"�ɳ�mEO�<Y"k��2E�%:�%�#1J�{��q�<����{}b�QJ_4�"�pvC�t�<)%'���ȼ��!ד#�u(��^n�<��҂PJΩ[����x�HYHQ+R�<i�l�{hX��j�6=�"!�F��M�<y0F��C���å��_ !�h�d�<�tB��Y|@,��ŭ![X���b�_�<���[�_	���M\/T����P	]d�<4�Q	���Q�� �Nc����^�<����7���z�@Դe�P�p���D�<�RaI���1�K8,�F@�<9�ɢ]�~lQ1$�*��ʇ��x�<��͔�Lu�@�
*5)�P���}�<9&��);�H���`���v�<�@N43G@r���>��U�]f�<	��T
.�!�wN�E@�	3��]�<a7n�+WSBy ���EX��4D�V�<�Q��7B����`L��r@�c)H{�<!��N�U�jѨw�K r�����v�<9��6X�T��o�>)!��Fs�<Y4⏚���RȐ�	 �y%�s�<��$G�'�(����L;���s1/�l�<��9/��y���3y��0��	S�<���فU���x��.?�rDSa�_K�<1@�Ȯ/|�!Ei�-}}|�b�_�<9����� 񕬀�!�����P�<�`!��d��	H���*5^�Fo�r�<�P�^����c ��v#8l��Om�<�D ��8_����_�KZ|	ӦVo�<qNL'sR(���BY�#@8�� l�<1%Gåyش����Qu\}R�'R_�<��*���hС��5�� �W�<&�@�p4�¶GV��G��V�<!��2�����+�.�R�<�1N S"�`J��!o{��Bb�M�<��ω%T��Ͱ&FL�&��OZL�<�▆j�PI��н7:S��[H�<� ܁[�iJ�8�依"�ҵ��"O�9s6
�i����- 	����"O�H'kLX
<tB�EX8!]p��#"O@���Z�lY�)9��C�FG�@��"O��V����t�AUE3����W"O��D(3z,Ȁ�gj�q�J��q"O�T˧'���2-���v�~e�3"O�%��@=�xP�|���&"O��b ��1VPH�k\�0�TpK "O84����>x&(���(i�ȻQ"O�AR@*ʂgN��@�ͼA�Da@�"Oz���ܧA�54nJ0�tiY�"O�+�N��\����X~�#"OҡhR�DT}c�Vc���G"OnL(s�O�)L�`(��4���"O4�w���8n��9��'^��$ �"O��tkE;i.�#�˅ N�4�T"O8�%� {ŐH3b�I��=aR"OT=g����aH��"��5۶"O>�ҥ�W${b(9E"��G׸��"O��#��,!�5�v�HΈH3�"O�����#N��!��C'����%"O�ݨ�hJ���=0�H�py�"O�q���Mc�I��w5x�*�"O���KX<|�x�ADΛi(�\SB"O�x�v*�D��j#픋3Όs�"O4��nɬ_�d�3Ekʥ��5�'"O`�� �L
|��=��HbJ���"O� �C�j��X�#Bg�"-X1"O��N]�P�Y(G�N��]�"O2�B�EN���֯�^L�S"O ��*N24�r�p�$\�?�X��T"O��agȅ]�")Kg�D"�(� p"O���sɂO���X�lC����"O�d�X�\��A���;O�P�"O��#�E��d� @
$iS�}
}��"OzM���34��I�Ș?,���s4"O��!�MU�x�g^�^sh�Z`"Ox��/U�k�|q���Z��ї"O*,D�Pkwt�����:Z#��iS"O&�JfkL7x���zF�p1"Op�I2l�	Z
��X�\�B��Pp6"O���"�
�������/��S2"Or�ҵ B v����Lɛ:FXɰ"O����DƢ@���:D� I�nhc�"O4��B(�HX�
�j�!-�d(1"O�}�UA-hGh���'|���)�"O�����bR��6I+�lTiB"Od��Sf!��=@2J�N��a�"O��%�'s�M��

H�m�1"O�\�!+̀&�ZL���� ���ʕ"O�x���]3F$j��dN3	����"O�3��F�Pl�f�Р
g���"O��k*<�AB�	�i*��*�"O$�����M�UJ�D��)&Ɛ;�"O|�@�Yt�B�D�BuBIz�"OV�a�d��HA#���(Ӌ�'�ybDB�#�Zs�Ƴ��
�oԗ�y�
79T�V/��V��l ���yB
·L��$�'n��M]<I����y¦)7�Z��A�\6���[B���yr�J�q�p,jA&\�'��M+�ŉ�y��H�+)X��A��,�N$a0���y2��=,t �V�z���,�y
� �[h�}�`�T���,�<���"O<�q�瑳H$rgo��� �"O4=�@3$� �F���~l�{ "O����i�f���P�
� ��RS"Or�qTm��R'����
.l|��2�"O��QU��.6N��㠃[�*g�ł�"O�X�D� ��&��&}J��B�"Ov	��e���\b��Aҙx "O�l#2�M/�ځ�� �w�,�Pc"Ob��?!�nȊ^Ȝ��/G�!"!��J�fRb	�:Ln�=�!E�6~!�$�&e���矕
>ڕIЊc�!��H�5U�M��HHj	&u�'��s�!�G:.�����
�)��Q�g_?Q�!�DH� X����f��Մ���!��H�I%t�e�\	��#��X1 {!�YlT���u�/Y�:]��w!��m�t�U$��f�SϜj!�D�,-� ljcN��H�н{�a��NV!�\?��b�B	�t	f`��4!��&BB�I�h�ި���WC4!��5�T��"����5d��M#!�C-8��!-K�Vrbx㡄&
�!�I�}:	pu��d_z�� �.!�d�	0zܤc2WA{D+��.J!���	�2��%�_r�	�$CBB�!�@��@�� �_Ho8<���\|!�C4c�Py �n�;8f�9��f!�D~��ZQ�F�ob9A����{�!��"n���z#�B�*'���u��S�!��q	��y��3T��3O�!xqO���$�a�P�6N*~��+��)RN!��G�T(Z�������Μ�,L!��!τ@+��wpV�k�¥i!�D՚��S��Is]J��l�2$�!�DҨ/+�t���V�D�n$��X�FY!�I�v�q�%�:9�������0:!�$�?<�i�Y8D�`fڒX�!�D�5�p�R%��u9��%��p�!�$M�[�JX�%��@K\%,�!�d@�W^��J<3��D�&*΄��HE{�>����+dq>��f)��3��jeƬ��o������ݸN~�}���7�A��5v��Y�㕑4�,�1���d*h���]��(fg�&��q��������7I��`;` ���95;����t̓�.,�W�ſ5�P�3%�7Y��ȓT�� ����8BZ1�Qn��!�6�Ex�)rgA�]�d��P& G �����\�<�� aDm�&�N1d��@��\�<A�M�Zv6�C��D�������]�<Y�M�*�����:����a�ܟ��>�Ǔg���"%P� ��ȩt�"���	I���)�;Q�2Y
U�5�Ta��'����D��%��r��&D��|HA'��3�'�r�i��'R6M)���̎3Q���'a�G��(i�����yl3JA�Mj�� .:��pQG��y��P?_2As�bL ju,H�!-��y�&��e�L��/�㺝���ܚ�y2�ʊ�i"����e;0�����ybcƴ1�5� �UiQկM9�y��J'S򌘐gi�>T�$��t��.�y�(�#�ݹc�ܴN]
i��#��y�lRn�6I:��T5J�(�{aH��y
� ѡ��W�B,�b�æn.�CW"O�uk�(�
㤹ʱl��J���@1"O���R�Aw(K�!]�P�p����'�Q��@��X�L,�Y�v��<+\�t�Ā>?��s�8�'D7)�����-܁D}	�ēO�����Ԅ"����L�Pi�t�<A6 ��JO����7�I�4��o�<�B\�~�jz�.#S�x:��Dn<��z\�11쌖RD�c�QMv�&�F{����� �pp�Ԋ��q��@iV�M��p=q�}��[3vw@���㉍n�"�(����yrJĒ�)ML(���e�J�8��	�ȓh���&(�>��̈�.�V� ���t�xw%��Ns����c�zu޵��I}�'!�����?r��"1���Y݌t@�'Uz]�O�_LiB\�ś�'ў�}B��4	XԤТK�7�>��d�Hc�<1P�2�Ҥ� � @@�A�B�E~R�'�P�as&�+@]�ӨU'^E��~"m�d�0B�%65����f���y#��iYt���'c의�C[7�y
�1H�L���K��IвP)N��ybj�'G��d��%�5s�)��M���d׬�hO>I�C$ܗQ�H\1ALY��Y��C#D���
VN����G�w�bI�"D�|�V����@@�12X��1h>��;�S�'Wf���:�l9��a@�R���sg�p����E��9�K#�BP��I}�'�X�� �����zkB�C���'�$�kC���n�f�
���pr��r��9��V{�S�Oo��JD�3 %�򦇉Z�0�ф"O
,胀�w��d�%F��-�F���"O�u���"�2�<)���	5�h���k`d��7����Bώ7o����"O|8�j�6-=��KB��0��Uۖ"O��`�FT
kX��k�,�2I| =R2"O�|�����*�d���87B~��0"O������-E�pd��/&Pp�Y7"OT�@ b *1~���m6;4��"O�DH,u���%�ѵP0���"OZ б#Ԍ#FR0�E�,�(��"O QZ CL99k��r �M?����"O�m:�(B�.<��[F�<K$�	R�"O`H`�e�$�J<bV�ٔJ@���w"O�L���:ذ���ܱ9&v,yv"O���G��43�82!.� ~v�Z�"O���3��~���Ӎ�y�I&"O�x[�پ.4p��+ԍW���r "O�	��`��j�d���
�M� !�"O��KG5t�)�VI�D˂�£"O�蓀�8HG���%�ή	���@"O��N�v �a&٘U�*d�%"OR0����	�^#��\k�"O(��%ңC�n���.-��x)�"Or%N��Tt<;��(e�ܝ+�"O���v�4v.�͋ӣ̇lh��U"Ot��"�j�z��ԀU^�j� �"O�$���~�n Ȗ �r����f"OH� 6�7�"x:�a��M��L`"OJ|)ĭ�̢9(�f��"�>a��"OI8�X�|�.�x����<�،��"O�I�Ӳ`�p�g&�
x �"O<Q�K?BExD;�A���x�"OfM�� ���u���!6J��)"O� ¸�HѤ��]���Πq\JL�F"O�]�s��l�,pʂ%�+6E@[�"O�i�s�	.In�/̤<����"Ozm
�h*(8�f�#m&fِ�"O�u�&F�}'�0�G�K�`!	p"Op��'8MV��u��>w����"O�IJ�	�+B�҅͏[�.�Ks"Ob|�TGj�` �!�zH¢"O`�sǁ��iJb@*gB(��y�7"ONdx���h6$h���>�5@�"O*@�P* ����4Ě7s�>�Q�"O~�k� ְa��X*�G�uy��8�"O������3r���c@G�i�\AQ "O"T�TE�B��D+!�p��"Ot���n�*t�]�bՁ ��L("O�a����b��mrjK��(�""O�Lр�S6�����H� �~���"O(`�r�E�g�4�T����΁x"O��k�L r  �y�&\��tu��"O�a�R�-z���$OX��a&"O �Z �\.G�n,@�M�`��S "O6	J�ɕl[�tbr�X����#"O� �v�Ku��A2��Ծ��1"O�#����*k��ԅ�F�ʕ��"O���$-�K��6$G-oE֨�!"O,��Ю�ll���b�u䲡d"Oh���BM E6���$��< '\�0"O�+� 	}M6L�R.I>$����"O*m2�"Y%�`����7��԰�"O��h㈂�jxUd��4��T�"O���m��`u���fڄ7�X��"O֜�E͏, ����f~8���"O�,r�hȆ:��|T�Ζ`?bi��"O
�q��maΩ��×9\$Ѕ"O0q�Ŭ��x6 SS�(J��E��"O����GȷV��ϺQ��u��2D��LB7xW�0��mǍq��iSa�-D��@�&1]>�e�e���	����U+D���Pxp��RmŤNXv��)D�T��P%�d١�Y�4 �	��,D�@k���2��m�S$�'��$T�,D��X�oŁl��2lM>S�|�e�6D��p�bY�R D��l��T��`1D���*����K�	��kZ ��+0D��z6읇E?X�[ m\�$��M*D��j����`m��֬+*�1#�*D�8�Iz"Y���<d6uSҨ5D�$�ЉK�8���ʦ�ӧd������-D�0ĤE�u�8���B?
���#.D�|�B�T�ɕK�>\fv( ��*J!���# 6F(����(-
��Go�0 ;!򄇾:4F��p��-<:Q��\�!!��
_�6��Wh��/P<h����+j!�Բ
������:( 
S畵�!�D�:j1`�dՐ&� ��O˘G�!�D*��٢ǈ�M�$e Bm�!�.޼<��n&z1�a;Ƥ�s�!�އg�6M"�I8�=Qbd�*)`!��C���)�I�H���@,V!�d\�3�ޠ)�N�7q͚���@V�LT!�d��&LT�� Zb�y@�7!��b;tչ�cP�Gl`�	1V/!��%=�x\��G�-<D�@E �\.!��|�=�# B����/d�!�� h�Y�j��,�3�΁�W"��*�"O��5��5c�Q �G�H�yP"O����ʇF� l��ͺ'Sh��"O�(aĢ�~�����ћL��c�"O�L�c˒�7��I�rA7�6�Z2"OR%�$#G"C��5�`b�<�*hA0"O�IK���T�&�딧�!<�R�C�"O�M��w8��3)�sc�(�"O�Ɉ�.�eĐ0#JE$(�܉2�"O��P5D@M�,�R�Δ�S�ș�c"OT�Ȉ�)��@�a$�_^|J�"O�d;��1 �3�׬\�(R�"Oʀ��LU�XT���&UN�p"OfH��xK����/Q);lJ��"O��8��5nu���#�P�`� iJ�"O2!��
6^��w/\:q��"Op�R� R�]�	h�!>��"O4��*.3٬��%oX�_�� "O�̳D�0f��ah���+T0�*Ob�;"
�1~`Q�,��kL�Ɂ�'�nl��)��t��3�'��1��p��'��P���
~d��*�!s�u��'�Pk@��X>�k�d������'�N�7�Ê J���H���'��`k���=wLLXC�B�F�'��$P�3K`��!`I
h�.�3�'&�{�GX62vZ�� $q5��@�'�na�'%Y���]�c��h�Hd9�'�. Ĩρ,�9CK�:m!�T��'���d#��\��Ï�	d�tl��'������z�6�[�Y�^=��'�l��h��^�f|3���P�n8�'mU&��1v���{)3H&0���'c6|@Rn�#6��&E�~9Q�'RX�)�@8�F���+؆A����'���͖b�Ta%���t�a�'g8E(��!�j�,D�<o�Y#�'��R��0[!��!&�*1B��'�D㴯�9/����lך,�ȴ��'>�5p��i���pu�o@�#�'�e�� ٤�֕�C���Z� k�'�(X؀��3�bëW�R� �c�'j��z��2}�ps��H
��x�'���x(���N5�����$�9�yF���aBO��B���»�yb�ŸG��5C\v�P�Hug9�y�OE?p�Su!Ngx�ɐT��	�y"A��&�d�2�&D!,�lZ���y"�XԼ�{�`�QS���� -R�D*�_)��1�\�~��@��`E0�ȓu���`�K�0A_�h�"�%8Ȩ��m�$#�Dݻ-b��Q�Ye6p�ȓnH�R�#ʜx��A��.3#.��/<%k���7٘q�[7�@�ȓLy��#������g�8܇ȓ�"��`_|���ӆ��<�d��*��jS.�3XmpDZ��� !�^���pj�p6�C�Wj�����5��ȓ+ł��fcF6Yg
��,ղB�A�ȓI)��۔aH�4������_'�P���D+��@�>�&�PGY�P���'xў"|rgKW =<]��M{�T9sB�[�<	��(>Zq�a�_ !ҭj�c�<1�B������
L�\�|2֩{�<� �����>2�
<{���&ef~H"OҸ ����cS��1fb� Y"�c�"O� ���N�(��� (ܞIVƹC#"O��g��*Np���E�v&(0����'��;ғRߞa�C�<|� e����A��F�4�#�H���  ΍���)D��R��	!E ��o�(a>@ 4:D�\IF�� �"Y�2`��4�<x�b9D�P��.Okހ�7
�f�ν���2D��YQd��1o�lxbJHg��!�U�$D�0��)�p�<x�ć\����$�'�\��1�B�<Q0��es2͂k��rl!t�]O�<��ꃒ��!��)�0��I)cO��܄��:��7d���
v�G�:���	w}b.�ß�@ǧ�[$�Z�+�95.��	 �>�
��o$����f� $t��W�ȔDa
8��IO�d1�D� �e�R�24��Ch^!�=,�T�9C)�j�h��'
��!��</�
�����:��`�#���"�!�D3]�xX���� =kXSp�O :�!��Q������LW"1�0,���!�$"���2�Dh�XaZ��L7P�!��E<4���Hցv�}ʗ���l�!�dH�t9&�s�Ϗg��{0g�+x!�D��:�"���Nيnx��H⤟f�!���iw���!`jp��D��B�!��=�J<��"Ȯ�#�^�!��I�"��fݨ%��a0f�S�@!�d &Z�Չ���*��4�#-ё�!���u5���F���E9����� \�!��Q��"�7	��n8D1)��^�!���h|9�$п!2�@*vH��!�Ć k�Vx��� ����LT�h�!���2�l��&�}��z��B�>}!����l)b���\ %*ʆj�!��
5gԖ�(|� ���8���p�'If5�!�Y��P W�W�$9��'�搋�NR���6d�!.z,�
�'�,qۧ��-��"F��-N�&�

�'��!�#Uf:��d,2���'�i��G[�KW<(bw��"Y��Y�'6j9 �I�!R���	��A�L�'3 �z@F}(�i���A��̓�'��A��@��k�(�A6o9�&��'F��U^��X͊R��E?�	J�'��T#�+�Up��k��W�O&89 �'�T�x�H�qE*�@�I޻Nc�q
�'�BE��LR��^I�!C�z8k	�'�}:�	��tx�-Ŀ%�90�'d�R�������{��<
%
�"�'p8x{0��P;V�`��A�s��ax�'���	�Q�L�@�7!ڠ�y�'��rF�΃Hc<�H��ɳh)�	k�'��R�	ǼU�
d�J�(21I�'N�m��`y�m+��Q�u<����'�����"��w`@�A��p�иs�'�Z%���l���˽d�8�
�'��)�I3iw��µ�˶4!�̢
�'��hc�gH�͐�s�'�_���	�'�\��f�2g�2��/ΐ]����'����Nɧsy�͉�A)M��I��'����-W�� P)��Q�p Z
�'�֬�5e[&#'���4#�6{e4�A
�'�Q��)2U`<�����l��d�	��� ޵r)׾(�2a�䊐,W���Q"O�x�=3��9�5
ŀ&��8��"O�a�7���,�6��Ȋs��R�"O�L�V�BcB��ٌEUtM�b"Od`С�	�^�<�X�@	�UJ�	"O����Q@��Ur4@A" B҈1W"OH����M�L
\�PE�\Z&��a"O�)�(��U��H�ı�f��d"O$��Ɍ�9�@ycc�;F�С"O(��PG91I��[�C�t��B"O�=H��3t�0���h��K�"O�ݹC�F*q]�T��Kɵj��""O��c�ݩ/l�0KbK_�oW֝rp"O,���0)f�	�o��BFܰ�Q"O"�˖�ե@��<�eN٥'8 �a�"OB)K��D����DX�j+&E��"O�,b3�˺:/�U�sb��D�}��"O����*	�\q�A�thxD�"O������47�� y�S�J� ��p"O�A���G�?uV�GlS@	@�"O:�� H�S5��#��ߦGc"1A�"O�Sd�K��*�'P9a\`P5"O <K����t �1����[���5"O�X�ԃ��SX���D��[��H�"OJ���px�Z��K��6���"O�e�7�\�b}^�S`�5h��)��"OX=�w`P�"�R�sRI���q�U"OD,��L�T⡒��IY�v���"O��C�C%$�xE�"��p97"O����nwis��M��$@v"O��@ģ,�(@�
N+{��e��"O���p	 #�4�''� ��f"O0
�Eْ|�:؋�G��@t(a"O2�eޫ{���D9zy��"O")��(�d���X�N�s�ɹV"O�2��KT����A�(�Ą��"O0R���"���L��C� �S"O$����KU���c����d"O��D:N�B%P����.���
�"O"�X%�D:#�j� �MI.3��؀�"OF8�K�5a����7͘���"O���e 3q0�S���Qcfy��"O��h�S�k	�q#��zy�ف�"O�h�K�'[f����N+R]��t"OƐYb⁯c��i:fK�s'zRg"O��S��a^��"a�5%x�;�"O��uI�y�d�&*�m �Ѫq"OґzC�3-N"I:��Yvb� "O�0�'Oؚck�q�R��&n4�s"O�4AG���$�`����w @��"O>�{4�CKEVX;QB\4X���6"O��Qr$� u�����(nnV`�7"Ov�k�@֢N�)�O�<P6\��"O���#1�HQ�@�/M��ء"O�X8GD�f�jx iϪ{��Eq�"OX��@/E�,�I�'Иu��eyf"OFp�CER�tV���Iu�H�"O���.��*�Jl 5 �ec� "O�YHR��.�B���l+�6��2"O�ي�I� �\P�"�P8*S"Ot�s�-Ϣ#�0]Z�K
L�>�8v"O�d�V�d\�\)�P�z9r�K�"O�qȷ���I69K��z6���"Od����P���zD �9��"O� �Q�fƠ3Ԫ�0�P�` s��'�BѶ雛�ԃ�*K�8%���&� �N��ȓ
?�$I��E�LdRC(ա�.��ȓ�I`�CT��4�V��ZE.��ȓA�65��&2����_�)�P��ȓ�89H疃V9P��ˉ5�`%��fj�X���,-����3�k�����0��@h�&E� �2a��-��:;F9`2��"n�=  �-�ȓT��cĊތ5��p��ҽ'���� [&��$"!���sFbV�|B@q�ȓ!���았c;���3h��!2�Ȅȓ��Yj� Y�{[�d�$c���.���Ԧ�A� @v
�+5�n��؇�!hh�tm�6��%�bۻr$���ȓ�8 D���v������?/�6U�ȓc5R��'A1Wd��L�[-�i�ȓɼ�JRH	�LbD�;-N��ȓA������>[f�Q�n��&=X8��.:*�jď��X�	�A�0Bm������r�&
=\��E�N(w꜅�ar���o��T�,F��}�"OJ��gE�y�DSr�
�5��H'"O���#[��1����}�:�: "O:88Ŧ�,�}9ׇ�Sܖkb"Op=p���5$�"�Ö#��}S�"Or�P"Y%pi4-���S�%!"O�|�q��1������ɦ7�BMh�"O�9IU!L�
�$��1�F�<�jq�"O��$+��8�
�"Fה���"O��P/(��;�兦r�0p��"OZ%�@�	�_!�i��N�m� "Ovis�E"NN� �ښ+�nLp��'Vvو�"Y.ly�g��9��� 5��-z
�I�חxW���_ <�^�@`BOҘsc�\�5�����&U?{ � ��\-*���%?�S�陖/�n0b%�5K3h�
��4D�$R��8E^ܡ	��O"9�:I���"��s�e]2�(����~	~�}��zfDа�Db��p��N�������V1h��D:pkb��fv��R6���4Fa�]�6��DQǌ)g
�]M�'�X��σ�Y�ϔ�4�![דBT����g�E*a*Ó�|���ñ���`#���v��%!aI��-B>��DU,ibj�y��ϋ,)`�i0#�*=�1Ob�y ���?�Z�چ���҂֙1�˧'�:d����U@�������s�ZA���Y>`�����349�k��<Ҏ�cf�U6��PC"r�q�l��Iq�i0r-�o�2QU/ܱk�䑉2�,4�`��m��8Ն)��m�.�B�[F�@�<�p�#�xq����~*���o>љ���F�c���o[,A�~��U T�z�ay"�_6Y���A�y�^� �l�+-���+�2i�-%�R�H�HQ��bߑ?��A0��'�*D)a��~� Ӗ�ʄG��L<�M�44�1I�-)�$�u��e�~D���"���œ+6�=�7\-~������>�y��Ш]-x!��LB�w�,YfC-/��u��0Z�2�('�g�4����h�d�8�w\�҇@\2^&4����vF��
�'�� �a�d�H����*I�U��

bT��E
t`I�R��7)��� �F`�Q�p�ܘC�l�s�+�=\���h3�?��"Vޒ\�♨�	�B���N�$����g,@�U�Tɋ���Ub�	�iO:�
XHEi�<X����$?�6݃d�I�Z�&`��_���DS=I��x����5��1�O��*�뤪�%^�(P�+����K!hS.#�(A�
ZKZv��U���:�2�:
�'��0x���4W��`צ��2|Ω�wmM���}(�5ubv�H�:y��<X�	��U��d;�&��0xı��w->�@ ��H^ ���,%%D|�A�@����
M)xJF��I����bU	9����*�e�NP�DL<D"@��3뉌N��lb&LM���kt��
>����O$���R�8��#.J�?��h����&i	,�3��>� �C�J;��X��:¨� �C[+Z<p�Gا�s/�&p��HF�U(�h� O�1L�������7��O4X����?�]�ΒF��A�`j�^��yq��7e�"!H�� t�a%�4�u[�'��Y��J�7R�{���XwԼ��I�#/BA��*^9uo�x��S�? ����W�DoDӠ�9�u��\�`a0�����Sp�'h���ɡ1��Q0�� �4U3�wh���j�vD��i���@��ߓ���zpU;^cླྀ�Ǉ�V�N��d)�JB��/@�-uf�he�L��T��d�)��2�F�U�@Ԛ�i��@V��"/A�yO�vUhx�h�<>�ѲBFL��'WΘ��ߦ��X@� }pX���.W�m�Q�%:��(�jVdf*�Cd�V�e;da����p�v��&�=B=~����<��ɗI�,�a*��̭�Hd;����~���� [�e'��
pk�0�ɉI�(�}����FDk	�{����"@P�A���C.
|��I��)

�9D�(�OiAV�Vm��2 �G�?(� ti�gbd�����/kn��acӈF�A�f��h��*���2>�@�wd�#�툿u�$�3����l�R��'J,x㶡ܢ��KB�XT�������L`����`�>��E�j��pIE%�Nl1�mÚ\S���^2X��W"�۞': �xG���� E��E�였��(��Vd$�Ap v�a*TL���a����.�q �b��\�a`ݱc�����9���-[��=�$�+1�	�D�Tb�l��1���4,R,md9Rd�$2��5As��M�.ъ���F�@J�욐3���d�-dr����[3�4B"L��|���ro�T�h��E��%����ڬe/�� ��A`��H�N�G���JƢ� A�}{��ʏ �0�jtK�a&��p�$�Fl�6��[�d�]�]~8\���:wI�B�B��n���䐊�^H#��,;���õ'P��	V�F�h_�D���ˡ-4LS�e�d����L�ظ²�C�&R��f��:i\�L��'�����G;:ͨ��T�05f	���DV�X���dDD=0݈��/04b�5!N���;��Al�B �F(,|��P����=pXА0vm֏S^�h{�hQZ�'犜�7E�-�F�KƂ^���bp�H)xP�|��˔=f)�I�ao�O1��M��X� ��W*X�U�E Z^�y9A��=Fp���<�O��� �֞+�Xa��+^�7,"�d滟X��j�\���A!���0��u� 돔N��i�E?O�X:�w��}#��P/3�lM�$ $޶\[�oY�!;���9�<���� ������E�"�"a*C�L�@]9���9
+��R�>���:�4���e�s@� ���1�������q��(ުAz$Q�q�r}�1F�۸� ���	?Pp���M�z���󄛥
m�AQI�&=�r�{+P C��|R�.F
=�F�i�xps4�DuB���l�Q�R\��'l��;��α	(��a�i͇V5�l���DJJe��#�퓝I����M�
��"�.�(3C�	�8�����^�kb��s�ԛ)��6m�4T�2�"~nZ� 4�1�e	�#,�D Xĭ�2`(���I-I��'��סedV9�ሗ�?{���b��uz�ɣ^�a}b ڂbWN�3Acт,�9�3Cʱ��DF�l��O�~��뚥՞ aBfGQ�r��`�S�<	����'���*u)��P���R�$�I}2<OJ�:�&V��D8�O��$叕k+2M���݃`���ɁL�
�j���'��&ȉ6�T����<u��S8��mL�]��\0�G	P��3�=�0�by��,�S�\��� ��Q��C�F�+U�C�	2G܎-�B"͖�⌣��7W�T˓5^<�c�6�)�'�ڜ:�#�Y�d�I�䌙���
�$�0�-v��8�V��V�6��<�f.ř��<��iС� ����M�PbX]Y���Z�<Yn���r݃��A�2C
��Cl\J�<�3c߀k�@ ��"PT��r�M�<�1��g�:�#2F"6~�H0�N�<��� .İfKXTN��"aC�<1�͒!|b��dO�8�2Y���<a#��-���UN��&��=p4�^~�<��&u8hjsO_<C�a���A�<	U�4m����+�`=����U�<��� Z�ű4��~v� k��W�<as� �q�D�e�Z��b�b�$�D�<q'�Î/�D2��4/�|��#}�<AA9��]�u� �8�1�j~�<���Z04&p�'�E��`]8 @Cz�<A���)Y(�E��'��V�S�<y"��%aCrxj�+L��y:�u�<��a����@RK����g�p�<�ͽ&#d,�B��KD��e@�<A*�)�:�ӱ��&I2�S�*�e�<��S����`ɰ����z�<I,�=M[���U=`��8��C�<� �@��/��KP���  ߐi92)�"O����+9lP�P#l�#"OR�x��"M*����>L��Q"O*s3��S��i�ނ .���"O��:g`χ<��,s���6"u$��&"O
0R�O��[c���R@O�@ "O��$�B,1�X��fR4X��,p�"O1�%E�Y��DPAd�Nqh�є"O6�d��g�.���O	C��"Oxhz��ʝi&��!LFʥ! "OD��'�2�����* $�\[�"O�I�f�.��� �l�(�s�"O`pj�T+	K}`��:`'9�y��A-2d��s�$J�iI��p��y�$�X
�J�������$�>�y��0Yt(���c�:u˖E��C���yReF�u�0 x�cX�T�h�X�!�.�y2+�K�����;q�Dx�'���y�A� ���A�h�f�۷�U��y򇜔��xJ��/.I��5�yb�3�.e�2�F �d�Ӄ
��yhV:h���N���R�/ӵ�y�%��a����Hʺ��mJmH��y��ʐj�,����+� �u��y�A���dۧ�yʧ'ű�ybĹ�r99'��>C���pW�Ϩ�y�B�S�t���0��+�[(�y��t��x8�K�4�V �����y��؝6V��'�ڬ"�� D�A��y⧃�Q��6�Ԍ'�<h����yR��>��xZ�dR��|A�ªC�y��MSxj�(���v�<!��\�y�& ��ar�j�c�Q��^=�yr�ߠ�0�I���^R�p �-���yR�J=Z�*����$#����ț�ya�e��Z&Wa���"�yR�H�Y�%�F�U�B�s��H�y�,f�C���)C
=PCM˲�y�����̑��O)�T蛣�ݔ�y§�T�HpXe/�(Z�� ;��D��y�ۨP�(8��)�[�X9S����yB(Z�<D-�Vi�`��ᐣ
���yjG�b�e���1@������y+�:0�(D�_�_�d�1�*_:�yB(�����sD؋��	h�c϶�y��%T��=��iΈ�D%q�횩�y��yr!y����=*�D���yҊ�2�gCǺ$4f%��(4�y��Ԉv�H�4G����"4\2�y��R�m����]�b̹�LƷ�y2�×b�&�)�"���֘뙉�y�/Ш�3���#�`y7� �yB��,)0�CK� }6�z�ʜ��y��E'���G���`�����y�)^lc��ު�\�S	��yBlϥu}@1�	�y>,z@� �y���#B��xe��f��9��jW
�y��Z�P�vI����=��ʇ��yҦ�N2 d�6�
9Z�츈��T�yb	��]�6�2�;��\���A�'����F1̞0д�ػʜ2	�'�N���ͅ,�t�s�'r���	�'J�ݣEB(L�@D�2�Gn�4 	�'ƤC�
�Rm����A�u������ ¤ �.�A�")��L�-�ε"OR!P�ኖi����d�h,�"O(0�oO�BTlt�T'3��4 �"O�%�gm�0A�J'^�t.ECe"Oظgd�oD���7�D8h[�"OȴT��1' ����M�Tk|K�"Ob�(M�Pp�QK��T�J�+@"On���$@���k�f΃(��u�"O4b�!�&���8��\� sJE��"O�hR��Յ!��b��4��1"O��V�^:1@���seV�
ԭ��yb�G�R�U��.sN��я^ �y�I��Cn�J��0�;�"ќ�y�ǝGx����D̉���IQj[<�y�\�%H�l�����!g����y��8J���ړ䈻4��&�:�yb��YZ�����	�9S��!�y���z���G�4W�3U$���yRoU�����埊<�f�yb$�y����@�\��􅈞�� �i��y��Ѝi�|��J�-Hh}�h؃�yR폕���:���0^��G���y�iلE� 10'lйK�t��Vѩ�yҌ[��R��,S@�4�K����y�\
V1z��t�AC�u�&F���y�Z�%��$���]�4	��A��y��
&G5�%kA��*t�Z��&m��y"`�]Tz8'ݾS��CӪݾ�y�)��'�y��*�B$���ɋ �y�J��>x������K�(3&�[�yb	M/2����Oт���y"lO��P:q�@�Dl@q��c�"�yb�X,g��E�^�G=��@b�K"�y�+;)�v�`򍅝i�ԥ���ɸ�y΋1J�`U�ֽk:��Ҡ2�yr��g(�( ���P�$$��D
��yb�L� n��C!�\`:G(�y��C�l>��Q�D�
A��bu(ٱ�y"���%�r¤uZ����y�.�^	���dV�F�:$Ö:�y2�1Z����D!C8���C��0�y�Ȑ-����o.l��}Ys`N��yRiB���X�b͞.Y�ꡢ2䗯�y���0�p��r&�^�n�j����y���hTА��H%T(�Ivi���y�A���UQ���gR�E.�y�	įf\�U���^���s��'�yB��%xlQz E�V���Pp�Y��yҀ��y�4�p�޽L���]��y� K7ʭbw�ߴ@F��W�yb�E"3,x�y,ߝ:3��k	%�y�F!5���!��@/?"0Y	�KŨ�y��V3�D���$2��{� ѿ�yH+B��%���E,rk$��a��yBN�܌�FN���+�@��y�+䐜��=�	��Ʉ�y�"ɜm|���"h�)R��Т�yRj��-�6��`��f��� ����y�7/�Z���m�+�2�2�����yBő%�
�����"����"H��y2Ֆ'�|��o>&)B���e��yr!P)Qf��+��T�E�x� � �ybY'��Z��ƺ`� �g\�ybF�|q��X����h:䤲�f���y
� �A[�l�X����o�	<H�T�""O�	�J��8^�8�/��OO���"O@ts�nn�,�"�	 YL��"Odݒ�`�fMNu��A�O)��h�"O��m�Pk0!+� $T�,ȱ"O��KV�<����F�w��P%"O�m�do��Z��+��J\IG"O>��p��.7�H}� k�9�(E"O�j�$æG�,��s�U�,=����"O�Q���y���s�d��	>��it"O�i�ez�p�b�7vʝ��"O���q��-8��i8l�A"OV�R&�6{���ԋ�%JX����"O��7��A���yd	֢L�L� "OB�����8?�tQ�f��B���J�"O ���CI�Mk�g\5Z��9Q"O�k�!cR�a���L�b�H`"OP�:ǈ]#&�� b��@:ksb���"ObbD%�D7X�Ѕ%k���"O�A g�=���x%�U>���y�"O��r$۝t�8Y���Cd�d�iA"ON[��R���mP)ǭ�b��"O6\i�H��wD�8[V�I&F�	[�"O�e�BC�SV��A�:���S"O��P����)r���eO1	��0I�"Oּb�ና^/�)��@�j��y�a"O�!y���1+����S _��96"O���@c/x@��ܑ8x��Q"O���
Әp}P�@���Gi��[�"O`�'�I����0c�8`;jAi"O�1[����Ń',�ac�"O�8�%�D�:w��5�B*9b���"O*)2$�ډ	��X#�E'1�$ѡ"O��c����F�fԨ:]�V"O�tY��G�g�:<�fD��I�
��P"O8���ɑA�P�pł'c�v�h�"O���C��:�@��bX���\��"O D Ԉ�X�+ň��pqjQBO�<�c�����7�
�R@��K�H�<��GU
&f,��-�8<D=#�V@�<q�9y)��i\�H����kK|�<�-�5b:��;UMӥy�ƀ�w΍A�<Q$�G̙L���k#	a�< �р|�օ�E(�z�S���]�<�LV�3pZ� �o�%?a�q�FF�<q�ה)��M	���m�SvH|�<qVNK�:�I <�")�E G�<)Tn�������j-+���}�<Q��̢iWީ��lKj���.@�<�U	���i�U�8�$��3�T{�<�T���n7>���W\��~�<�tL�9-HU����3G
��g�l�<��Y�3��(�:[.�� �q�<�(�5��Y��Y4BM�	H�Kh�<�ĵN�������+R����`�j�<�7�U�(}��cޚT4Ku��y�<��.�h\x=㇨� s ��b��<���G�> ��c9t��1A+��<���ڪJ��pJ� �j�IJ��y�<�7��<OXl9R����jЙa.�b�<��2���ɚ,Kl,ӧX�<�qHB�؀�	`Bi@ԠW�<q�GV�_x�9�nC4OdU��
T�<q&J�P�D�eI�!i(r	aTT�<� ��{'��rDs�FY�$�^�z"O�)�sj: i���zv
	Y�"OJ}j$�ϩ"%&���E��j1"O�4�p��_��}�N�9���"O���0jJf"f�YD��\��8�"O�uKe�ַMN�1�#�"���"O�M��dN>CTh�!bH�s�N-h*O����Ɨ?h�9d��iB����'�.2������pNF�X�樒	�'  e��a�V��}Sp�V�*}n\��'n����Pd�*G)��4�Z��'y4���])=�0kGA�7�eS�'�D��nF 	���IN�*���'v�!3���H��xva��]� ���'��U#J�2F�L#�D�%9�Pz�'s�J�ܠ?Ed�㎒D�-��'�b��a# ��$XP��?�`@�'���� ,�>��tAD�3�dy�'b0�Y�]�>\N�8�LݪY����'-��1�O����is�d�� �
�'��x��hIt1�曥_���
�'3Е����:��0,,|�⤫�'Ȥ|��'З4�$�j�H\}���X	�'��Ac�
�
v��� s��<'6�9�	�'E<lS�D�/-��8�nN��.��	�'��U�4BL4%N��wB	: ���'Ҙ����E^ّq�Ō9���	�'Fl�cc�O� v��˒� �<�R�'�`�IGQ+Xo�4��l��~Ik�'��0s��(Yik�h�r�9�'��Im� 2=�e�A�ėe\��'�Z�����+:�h�d��]�:�K�'�zp���f٦|��&YT$Y�'P�#"�,!`$�`ғ]R�y�'��$J'���WN�%KM� WĘ��	�'!x�o@n��x�@�r����'е+�ON2'�F��a�`��	�'ӈ݃ ��0����"���Y��Y	�'(,E���C	<����A@����'�\���=
�ƽrhC�0�'��`�e�$`A�� �< Q��'b�b0�	�G�p5b��L4>��S�'�e8uc-�`ԙ!(D�$��5�	�'�1�E�WlH[v���k�����'�Ќ	�`�.lNV���a��-��'P��z���15,h���a�#X��M��'�����⋘.�ֵ���_^n@���'x���6 �?4��I�`�<T>!��'�z}B� �Ê�C5	�3
���y
�'�]ɷ��oT��4-��v.(��	�'����f-NyI�O��d��`Z	�'��#a^�,�*�"���S��e��'�|��p� �8(��X@�'N+�a2�'$��CH�ٌ9�L=E���3�'L���e�Y�$T+'C�k����'c8�9Q���n��pG"K�_�6E[�'@p�+#@�\��9���]�N��<��'��e�#�[�����׋Dn$q��'��kW���K�p=�t.�=1p�'c���c�	!纠�Ą�<5�@��'�R��"^s�P}ȢaT�6��e��'8��1��A��	��e].q�s	�'��43��Ĩ&svxidE�	�>�"�'�9ђ �#DZ���'׹yh@����� �L��R(n�\��MV�P�4S"O|�jw@����`�a��fa��"O��R�g�)�^ ���Ze�T��"O�m�&B]09IbYF�֍�"O�%�B�RC<8��d�[Q�ը"Ov9J% .�*���U�7��I("OF@#"�����v�� �F��
<i!��	 /�V�@1I&srp���#y�!��ٍt�	7�ػ?l�ʓ� wu�~� ��`8P�	g��5\Y���	�L��u�X�'�.�����!3�,��w`��K�P�0\��?V�y�'Ղ���Og,]�F憙Fc��@6�QT�Њ" ��iel�D�d�\�UEI-(�܇�7ng��ڳݙF�^L�1f�&*�7�̑Yzt�3�H�I<��
�d�~>EC���W�D}ꡥơ�e�B��Tj:�y5m�'[h��'�����M�V�z���;�����M��$����4LU-WK����l�&�B�O�z����@1]��q+e!f� I�%��K���^7bQ�j*Ф���M��]��[X'̢��(}bpm{ύ�^Ѻ�e���
IN��7&�67����!q����IW7f�ˇ�!;z7N���vqk�'>|����O���e`^�A;��B��f�.�[���Q�Q�#ɭD ��i&�>�0|B���#���PЂW�,����D)N�2R-ތ,za��0^+��|�J~*��Ό�D�+٤}�^�z#A�"��Ȑ�a��!��o��Wn&�{ç,u����ԥD�8X�$��#|8��B'Oɦ����W��FTzԢO'�0|bW6ab,��b��zV4qнi��3(`�X,6m�
&��S�L�<B�Ȉ8S��y�Ƃ��!��9D��2&�
>e 0��,]	��*D�\��\m&` s��h�\��d,D�t�%�{ڮ$	A�?"�p,)�C)D�8��K_;(�9SI	�$�"|�A�'D���B�G_/.4��J�'��q�4J'D��H��-��d��ӟT�u`0H+D�t��b%�DZ �N����kQ�3D���mQ8����nM�W��ѹ��0D���/��D�e��� Z�=׮/D�x���7.����q-��\�5���,D�����J.� Te�z��	)%D�l�E������Ed��<(�@8D���H�H:֔*vG�
��� �!$D��{p	݀	�H}�!/ze�Ţ��"D�Tsщ�9y�� ���M%�Y!�d/Q�vU(�%��Lo��5ML�G3!��4m��AS�,
TҼ��k�\$!�$ܿY&�q��A!uB��s�IL(!���z,�ˁ'��g��'e!�$�?�j����R�ĕ{���
 I!�8Ej$�t��+zr��@�0!��R�-�<%A�o-rn��2�i�l�!�d�YB�j&	��Wr�Q��&f�!��wz� X�-�5r��4Fj�!�D��Х���*]�̫�΂�!�d"0�����Ŋ{��DQ�H�CU!�$Z�Ej��eJ�|�8�zHL�U<!�>(��(�e�r	� �Vi��ȑ�'���bԯS�% I[�L+]t��'�d5S7яv�$ᧆ�*Xi� H�'�Q ��'��]�6e�{>�;�'o�@òf�O��PE�w5^��
�'��T�S|�ty�ȏ�`D,M�
�'�>��U�	)7a�ě� ��&�� �	�'5�۷��.r��d��N\
��	�'i�QQ�F5�B�h"��M���'V���Ƙf����ve_(����'.M� ��N����i��x���'�b�����#�X��U��W䢱��'���r�J�)~��t�̨fh���� e���:+�����h���"O*�7!ϣU)D�0E��&tIt(D�� S�>���Q懍hq<!�G�;D�l8�
I�ItT��"��IRȸZ��8D��*A�?��*�u%�\���0D�L0A�Ţ}ܢ�A�F�(Ҵ0B�/D�����Ȭb�v0C�L~7�@1H,D�,hwk�#�l#�L- �^=y�4D��p�)�oS|4衮�I6��F&D�� �)�`����W�߽U�"��2�0D��Y����=栐hGL^9%`��@2D����c���q��#s�T�H�I#D�T1 ��,'����;+�$��'=D����GOB��2/���ۃ�/D�d&OѪb�V!@���>c��ifg/D����đ$�1�b���T ���*D��	����Er��q!!)� t�`�+D�\krb�>|b�Ѣ���q�U�-6D�lQ�׹��qbDL�y��2D�P�'ǐ
W�PS�G\����/D��ӑޡL�L���8HЙ1�-D��q!..��0X6gLр�j��8D��8��̞@�P�c�f�6Bfp�#2�7D�0��"M�+��)�5̛�	�`�ƍ9D�P� o_Z�&4+�G��u�J����"D���
�7<I>�h�3�>��@,D�L,S�qGz�3�ƀ�~
�P��4?I��ᓳ)����ek��q \*<fB�>$�2��%H� D	��[ NB�J��L�׫������jՁ�`C�	�g�Mx2�������c�(��B䉭1�]CA�#�΅�B�;X��B�I�
�j�&�-��8��#��B��&<:�!�L�3#���Q�֤OSrB��;bO�4!gb�2��8� G�9N^B��;�d3�iPWT�P�'�1�rB�	�`��JԱM|xx�c��
s�fB��8!þ�䋛wH�y��C�GQ�C�ɐ?�4]�V�^�~��8���%"B䉵<�*�)��m�����@C>C�ɼ�T!H�©E�u�g�5�2C�ɣ}�Ѫ��G�fN�!� fKm�B�I7!��(Q��D~9�ԣJC��B�	�N�&c��1YN=a�GK��B�I"0<�@��L/U�8�g��|� C䉍o����C�.5VN��TǉR C�	%z�F�Id��+�rL�(D�}�&C�I�h4`����U����V@��yC�I:�dG�]��6YAaˎ0D�B�q[�6:۸��w�	iw C䉰sJ�d��ؑz�:$i6�!�&C�I�@�NxaÇ^f�ȩR7dC�X�C�I!l?N	;E@�9�����¤>�B�u�:�8q�ίd6�0AF���iZzB䉢/�b �dI�b'f|�$I v�C��<]s���K��I�HT.C��B�	u]!b�V-��I��m�;.��B�sm�(�$�K���!� �ړ3y\B�ɻ4���!�I� ����Q"� 8C�	�,\���קm½cu�_�;1�B�I��`� F��5@ �@Q�#^��"B䉊MW��׎t5s��h�C䉯 �R�c�(U>��"u��*URC䉔$m�u���	�@k�-�������B�)� ��jV�Ӊ%�~�l;_b��:�"O,\�!��y�N���C1(U��x�"O��3�"PU�� ���	3���"OT���DA������ط"Oz��)�1�}��k?ql�%s"O�q��D*-��e�B�1NM��"Oz�yC�#����f�U:(3pr4"O\��2`�OP�`ab��f=���p"Ov�����X���T ��{)�� "OX\0����J�� <�c�Z�!�DE�kN�h7 �ό��Pip!��[�u��B�9x��A���"N!�ǧ[^L�uNU4�>�$�7]R!���w@Ҕ�K*�D�s�!��U!�DY+��M�Uh7}>�ۄ�U�^D!�DO�98��`@$��4I:l���P�i7!��J,6,q��۴0,0kc�p�!�$I`0�YX��Q ����M		$f!����E��e���R���!�䖐�2y�cÓ. �J'F��T�!�$	n(ɿ�b�Y�3^p!�@�E�0��ƁRyj}�Ԃ� {S!��Ny���&Gv ��h��EI!��n�ڲE�:c���Bg��Py��5?*y�爛�0�b�)����y�-ķE>D��&/�/����-��y��-\A˶@�1w)�d�Ԁ���y�(��8�3$�j�m�6�ߪ�y �<Z���r�*� \x&c6$n#!��ɧ6��Hv�	M��=�Wm�Y�!��서���^�N�j��c�
�!�d���R\80��w�¥����^�!�ȭH!�B��Q�!x��xW��2f�!�WL��9֨��)D`�p�ŏ�Jy!�dF�~"h	��%�*e0p���� 
p!�Ħt�l���@�.�w�M�D�!��
�C8�a/7]�l���I��=�!�2n��x�wfC5}
Q��:�!�䞀�X��6KD�7�v�Rr.!��:]b�[Ee_��I+ �a�!�D�<	�b��䂆]�����.J��!��9`��PDe�,'Ʈ<d(hO!��-
%Ra���G޴z���=/!�D�	V*k���I`B`*�CV+!�Ę8a�,�AMPqGP}�bXe!�D�x�T������Q;��QfD�0E!�'*��;,���34� %!�E��������� 
δ$"!�DF<yL�R�
�Z�V���o��V"!�D��@� u���+u�v�2čܝ<!�$Y2r�(��m�1F:^�T#�:#o!�(_{��1DL�%B���ۤM!��7�t��F��-��y �لC!�d��e|B��B�]�n$*�a%�D�>!�x�Da��p��3�>]!���|$ޖ�F@���G�
/`�`��
�'�X�#��Z,C��cRj#]����'!, )&�	� 9"2��$�
�'���YѪ�3O+$�Ӂi�}8v�`�'�Z�p4��3�&��RW������'S@P�!�d��T`W�U� .p���'��ܳ��c&-��-�8&���' ���@v�d��R�T�J "A�'������Д_혙����5�T��
��� ��V�մ.��j%��p^�)B�"O��f`P�a � �mʝ~Vh}�1"O�}a���*�(� d��|T`\�"O@�2C�.;(� /M;x��Q�"O��!Sfߴ}������;�*���"OF��uA��{a�	��C�4�&���"O� �@O�	���0nöH����"O���$�0�$Ხ��U��Qa"Oݓ��
�d\��^r�1���y�	Uc�	��֞B� �H����yC��ӄe�0l�3K����h
��y�)�hp���G'�t�j����J4�y��Õ5��ɂ�H	[��p��EQ��y��0���%�ߡP�E�6$�9�yR��UV!�dn^�JrD�Pv��
�y�Rl1�"!N��F�ҒiK��y���90�����FԈ�tIX	�yR�ѽ(|���̙!������y�-�2r����qkU2s1~�"�
9�y��ʯEN�� si�c�~�)b$���y0l��$!D�Y:���!'��y�FD�;'� ��Mbg�3Q��y��0Y�yTl�Vkr��J�$�y2�Ȗp�e�6/�S��E�@%W��y�l�>3�ܘ���F#E ��x�Ƈ�yb�	V�:�;"��X�a���yDV~<H�h͈Bi�I� �н�y��;Y��Ԯ 6�����y�Z2l�4�$mP��hY���y���D�B��L���r�� ��yR�)
x;�h/B���Wd��ybኺvJ�H�d(��UIޑ����
�y"B�&`��D�\@Ƶ � �yR��P_�5�a̲R��}[��/�y��w�PQ�qbڞP�,T��y2��E��<� oLL�F��2,0�y�ڵZ!<TI���H��R���yҌ�3LPв7/P9Ɇ�����*�x��'���B�h��0�iK�a�,�����-�b��N�O����O����ƺs���?���k�\pID��~��I��Ų{�y�&�r\��N�R����W�'G��`sd�	K,PH��#��7���BԎ3d-�Ňȼ ]�p��/@�]E}�QK��Eȍ�-�Fj�e�,$����j��v%=��O��!��=[��y�·�yW��;������I_���)$��%G�=K n-a��L�2�Z�]�.]&�b�4n��&]��+���1�M����M���p�r��1�Z(*D����(x�b�''�<�a�'�'��(����;?F����M���Gn,����j�o�`aR f�mX�z�gؒW��Q��Ɓ�j@ HY����iDH��cmM�h�p8�So�4F\��ӵBi�J}�3j<�;>�����ѦM�'i�epu���	U��@�A8æ�B�'��'^�O񟆤��
��A�T�K�@��,:`�Ou2�)�'�-	�ȇ0PL�d��,���5�A��2���^�� B���Mk���?�,���cmӤ�Ӓ�S�e�0i�Ō6E"<���AZ�� �I)�"g��;w|�����+�M�*�D�'5���(H_�l�8���$c $����.��	/��9� �#q�ҹ��k]%������А�5U�
��C�HK<��kĜx�ǀ��?��i������6�U4#a
���xQ�V���O����D9��Xv��)�r��daJ&y�N��'�X�0�O�	Z��q)�4�ēeְ�C�ǹ/�$|pf�QkL ��zӒ�D�OH���"s�49T��O����O�����!�o֗^t{������B�f�0#C�+@��� ԀK<�ST>�ˏ{�K�W�X!��Gs4H(��%]D�l2�o
�!�	2vN8����L<��W�_heAǓ�zNQ[�C];L�x7�EgyB��:�?�}�I蟌lZ x�
�9GK� h(���Q�� �N>i�D�����-v�¥f�<]�r\���?YA�i��6�7�����I�>	T �B}�mpE�Ʃ]��I�`Aٞ@R�
5zӮ����O�|��Q0	W�ͨ���D��\#��_
>q��&S�*	ΤHN,b�,����_- Q����8	�ԳM�{�f�uAkRi�s�O�IQ  �Tʚ
d�� )"<qq� ��8��L�+�,�xegԘ����%����4�v�'I����>!��E�0�h_f�ƽ�#ʏ+r���'��'��x9��Nq�4P�����~�8y+*�dP�]��mZuyb���r�П�m�v6����ս8��eh�6�$\p��?��K�?����?�wGؠ~�~T�N�+�M�,J�\h���l�dA�dPDR��剓�y#�m�;2jB�  ��W0Dp��PdCZ����+v�DܨW�'v������������T�*���� �4��1􋹟h��ԟ4�?�*f�%��B��m�8����n?!I>I��4�����	
8Q��y�%e�9C&�#��l�K��ǟ\��Z�IK}��L L  ��     �  �    {'  �1  8  J>  �D  �J  Q  ]W  �]  �c  'j  jp  �v  �|  4�  v�  ��  ��  ?�  ��  ��  @�  ,�  n�  ��  ��  6�  ��  ��  *�  m�  N�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6dz���s�<CMJ�(�� 2��3f`2� 0�1D��k�,�!V`��1��:_�
��AE/D����C�qÐ<[��)eî�X�-1D���a��#W`�Z����� .D�dI�j¤E�ɩ�C߃;�(Q�3�+D���k�
��1�`f�<�%5D���u���W�^��2I�:X� �H(1D�ܨ�Ƃ�/�Xm@T�ݎP��V�/D�����[�k���G蛥I7�PJ�-D��p�c90;t�R�X
N�$���9����̝k��ݭB�: QqB�<�W�84���A�uFݩ��ޘ?4�H�pA8D�pR�0YmN�Ƅ� 7T�����3D��n���ySd���~��P�'D�����&�
yA�f׬<����+'�O��ɼ���QQ/H�-8P	����1sHB�	/��E���MB����$Kn�?���IH7
�t킥`����[e�!z!�d5�v`	sK
�	�h�17nB�~�!��W_,��y1��93ʠx�t��Q�!�¿Y{9BcL�JÈ�b"�\7���p�X�>9��c8�Pk.�-�8ip6I�=���`�h`��ۤ+�	#@!�.����x" 8�O�p"���)@�i�J�"7v!����nZA��2�M�_w����D��QV��ݲ[[�aa�'(,�
c�� ��9cTŁV�*�#��� ������p����!'�"�h�"O�#P��C���k!抡$�-�"O�%iƯ��N��Y@�"J�m���"O01"S(EJ�h !�`�q���I#"OVQ��H�y�� �� B�">��g"O�I�1�����8����9�ޤZc"O(�1�S6�N`�E�ے�A"O�|bF�L�n��-��:s�|l��"OR��� ]��h$jD�Y����"O�ѫ7ȁ�:�J(�ǩ���1��'T�'w蠨�J�#]�;�Z3vؽq�R�'Ǿ�8g�
�V���a��K����'�L �0͆=v��ӷl��?��{�'�aR�<�� k�"�!��d��$�6�yr�ϲ/�����,��b l��y���"<"�{�nޝ�FɱG���?9�{r�|�E쁤h6����/.WhqCC'Ev����'_ޱ�ǡˑP���ɱ�`�Ω��'z �c�W'l����@��R(��
�'��D�U��4]�a��
�m^�r
�'\�EY���`	���d&Ty	���k������S�<��L��V��|��i�PY�1�I5<}�`��H1!���<����Ɋ�3�n��3��� �����9X!�d�-Y���шd@��#�% gP�O���D��
Q��-�t�Zi�S/G-?5!�R-VFi�W��%鏌^���B�?$�L�X>�ƵYɆ�,�i%�:D�p��I�$Z�A@W*�:Vm��F8D���vl��q0���e��gm7�Ƀ2ў�O�B5s1���Nԙ���X2��M��'7l�{C����yP0��$1�u�'϶$ځ��Fgt$���sUDɀ��:�S�t.O�^�C��@R �v-���y�#ڈ��:vd+�X�@'���=Q�yb�Q�
�<���Քb6��[둉�y�"C�"zޕ0�<^�Z��w+K��~��O��s��.�)�;�$=����=�(8��$��B�.���j"ѐP�<�'J�B䉴w֖YӊШO~����ą�8Ͼ����O�>��=���2X�>YgĔ�G���]�!4�ly��hWg�� i�����e/IQ��pU���T�H�ȓ8��H���G�VT�G�I��Ȅ�
%�	��h����%��Цln���8:x�Qc�T�DP�XXt��=85&��r���P��9n����&�V'���ȓH�xiqBEԓl��J�AX�7���I]ޠ�Ջ��'��-A�e�4'>���R�rP�	!AMJ �ɛa"zЇȓI�X�,��cF��$���]`���ȓc�x�KSmҖH՞�P�
A�\� �ȓR�(��6{���hA�_�w����ȓMsؑr*�L�`�L�2?�t��_}tͩ�����j+^5y���U�<IaF3U���V"q�L)橙\�<y���a�*D���q�hݐ�@�L�<9����P�]�X���x�I�K�<1S�P ki�̫0g��:<��)Z�<����1���gŞ�T6�D��w�<���!-d@��%�%����3aw�<���̱:�x2�
�x�
"��G�<qK.c)��2��K�%�=�.�C�<�+��.�nP��j �VT�gIMW�<� ��Ig��&!V���
>y��c�"O��n#�R�8����&JD�3"O�P�iAe�!��lN�$3N�;�"OX�0U��J'��"&��$&��$"O���%#�:(Y!��%Z��3"O���E 6�8
�<(m�"O�hRB���io�	�.��с,D�d	"���]��8��G�Fr�'�6D�X*�J̤*�$#�
E}���)/D�L�f�נ[�Rh�LD$7/�d�p�-D�|���LD����ŗS�rLr� (D��p�jX�v�@�� � ^ ���	&D���矔gm��cG(�% �:v�7D����a�gT2��ؙ2�����#D���tO�$z�ٳ/̅j��=�k"D��K7#���쩴��r�I��?D��	�ai��|��T�u[w=D�X��-t�·�R� �n�sg&D���n�|��E��1nR�C�/D�|��뛫�����jC�4f���2D�3r��a� ���i͓~��lR� &D� 9��(��2ӡ�,9��Xvm"D�L�P��6Ȇ$��-E4.����5D�,��Û�yc�([�n�G�:��3D�l�fа%f�d� \��tR�,0D���v��0���q@�6k��3��,D���ĭ�&9�Y�����rNL��o*D�������0TC��?(�!��(D��{ I�YzD�R
��԰�#g�:D��)'�˙PتQ1�o�L�~͉�g3D���R,�}0����X휡���2D�PCs�9� �ŀ[�3��k�2D���a�7-�p���.\(|1�2l.D�Lh�Á� �,��(�(�X��H-D�L"���6���e��}�*Ӎ>D�|��)ċ~#�T�w��	��Ɏ$�!���vjH�4`�#_Ͱ�ȁW��!�D��}1a�WDY%��!�G^<�!��ò2W>q�)�r����$S�!�䄿d=|��%)GQǈУ#FP�nj!��
i� �����>���qFU9!��?̘ f��u��R�1&!�$D�Lk��{��P�)K�8��dP�Q�!��P���tz����<!Q$*j!�R�+�]2agJ���C׽d�
�'��ũ7��$b���)\�i��L�
�'���'JG%^���:�fa���q
�'�̡��-��#
��⒍_8R�s�'z*�7�I8dJPB��n^@S�'Ѽ=���ӹ~�8��1�F*x�":�'x0�"D�!�hT��M4q�����'�Ј���~v0| �+�h��0�	�'��!C�E�(1�}��c�,���'z��S�Sd�2�NP/�`�9	�'鼝c�MZ�,�^�IQ�\"$�����'�6�S�V8|�}����+u`|��'y6`��&W(Qq��ð��D�'��m��G^Kr���ꅍ�@!�'�FQ��d!zt�(�'JGSF�	�'Rp����M�^��󈉦�����'��щT�J�����
xL���
�'�M�����ԝ*c
�)[����'����6���y�Ѐ��Q���z�'ET	[
�'v��I3����ţ��� �ܸ�꘱Pv4�U'�<z��"OΡ*1��$
�D��e��I���"O.�2O
�2"E���
�j'"O���RgS����#��փi��D�1"O�%�C)ƪk$� !�_�-����d�'��'f��'���'4r�'�R�'�,E��K�4tX�� 	m� 䣷�'��'=R�'��'��'���'��`���M۴�T�?�p�23�'R�'gR�'�B�'L��'�"�'5�VF�w��	�&�!��U���'
��'u��'���'��'�b�'�܋��Iʹ0!%=�y�P�'���'hr�'r�'uR�'���'�T��5�&�PRF�S�&�J��'���'~��'���'2�'��'�� �W���]l��g$Ȱw�lt���'���'}�'O��'5�'�"�'�49چeUM��X�3i��(�Z����'Gb�'�2�'"�'�R�'�R�'ID�5b�03����(G�{0����'�2�'qR�'���'8��':r�'Ң�"!ʩ{^zD�p`:l8dYq�'2�'��'@��'H�'2��' ��8c��8t�Z���O;����"�')��'�B�'���'���'���''֔��D�n<�Te�S�&�Qu�'�r�'N��'���'�2�'���'�����oD\����d�r�h���'�"�'6��'�B�'�"OrӸ���O��QoW%H`t�S0n��x�����Nyr�'3�)�3?�@�iʰhQL�a��=�w�� "�v�k�9���Ѧ)�?��<ё�i���7狍+�Q2�IˤR���a`���DԘN��m�4��0�b	K�c��}�"�~:Q -}���H�\�eL*`s �E��?y(O��}�a��\y�#ғ}~�̃�Ɂ曆��=��'=�R�lz�� ƈN�O0��9�a�+>��}@_��M��ir�į>�|�!���Oi���T.�ŋWL�k՘3Ħ��CE�ϓm�t��7c� �a��0��|J�\���[�GYg6<5B�(B}�u���$1�$�צ���1�	�a��	���Ϣ4+��X��
���?�wS��ٴ%h��2Oj�7��ъć6vЭ�@�Y�)�)�'G� !Ǎܢ��u��D�]�=��1��'t��%�*ru���dS9>Ր��PW�Е'���9O��2C%
Iq�(�N�3-�=K@0O��m�������&�4���1#@��@Z� �.ÿc����?O$oZ��Mc��y3w�R~b��R�y$��l����	�6$�Aj�7ky�Y��D$���~RI�*�.,�}&���䆉�Aj�����}T�XT�5D�4�C������#���7? ��f��=���`�3!�9ڳ�Q�ejAz��L�ڸ�Ra��#p����!��0��aȈC�Lh8��T��4����ecn\�GK��dU�0�@�0G���vgÞo���P�Q��d$�2�
�y[���B�IPA%*w�@�Rs�A0&W�@H��
/�L�Wdt�4���O���z��'Rtx�"�%EĠ��k�U�����O,��]�k��⟤�3�DF�gE2��s
L�Z� ��^oӛ�@�t�H7�O���O��	�i�i>i*�W���ոdm�r=�<��M���T2��'���y�'�� ă:F� ���Y6~kNJ7�M+���?��E�Nt)��x�O�R�'d< ���SL��	X�W<�@�s�H�$�O���Qg�p�OO"�'��'. ��$,�̌��S�S�%9��e�t���l��u&�������'�֘�.3n�Mb7k�!�BTFc�~�d�d���O���OR���|b��P�i���G�sF��1�ON����H%��'�2�'b�|"�'��0�B	6ɪ ���O<]z]��FX1��'��'�\��n
���4&��BYD e��,2��@y� ����?�K>I���?�&lB}�aJ�>���J�:wJE�Ѩ���$�O����O.ʓtVTО���Ҡ8*��@��Θaj��`A�bL�6m�O�d-�D�O\@"�i��Q�fH9r�T���h��,z��k�4�?Y����dРh��%>����?�	�:Y�tpɓB� 6�`�agۑ�ē�?���Ɛ
���?�����SER�a��k6�Sg��{�6��O��䞖 ���lZ��	�O�i�O~�&տ7�̐,�So&}�Bʻ��D�O��(��#���?O(U2t��+D��aarKώD0R�V�i��5�yӬ��O�����V='��S����!��K-[�b ��ƍ�Z8�qߴK�f!����?��?��'��i�|C"u��p��!C5fy���L�E֛&�'�R�'d<��X���	�a�Ve���֔'��T'I�9�VO4���`�㟀��v?��
B�`@��� �,�����	/a�$�'}`���'����*Z�m�C|������M;�jp�hI>)���?a���dߞL��D�T�Ҏ#L���d �6}|\���D�I����T�'�r�'�2%%`Œi��KE��k��̢2	 L,R����� �	Hy��K�-{&�,bzLtYD�B�*d���V��a���?)���?1,O����O��r6(�O��X�FQ1|���#��I/�M�V��Y}b�'2�'��	b>l��M|BT�����2"�ߣ(���`/W�L���'E�'(�	@���	K��GCY���Bù������1>�6�'bP��pď�ħ�?��A#n{P�Z��0�����Ӧ�'��' �(S��'�O$�\� NQ!�.؞[l�#�퓢<ю�+�x���'xZ��$Y	M踩���R�H\�ֈȓs�!�_�*=��A�>,��=�ʒ��E�2�H+y�Xbi�$u�Y�N\/:�d2v��*8����ȗ͜�����H�l4������S�웏G�+�HH��aH�9;׆�x1�ͺd��T@�����I2���6��%d<K"��W�@��G͝4�. j���$��d�N�t����OR���O| ���?���8,��Q�2�B0�⁅ l��Z��'��; �	�x(��wF{"��6"���A�>B{�A$gB�o��0jb�]:v
U"E��`�D��O�%k�,f�@��V*��Q/6����R��-�n���'h���|ΓM�.��ǉԖά�ƅ�X�Ąȓ �� ����ɀ�H-U��T��)*-O��8U��M��
 o�n|�u�Щ��/[�Ha��ڟl�I�� ��)埜��ޟ@:�]�{��˴��<�b�@�`W/g� �"��!@�xM-��dz�I����5?�@��6�,*�0�2�˙�k�
�{��C�
 (A��n�c�zY��>W��$0C��Ӹ'o����?�w�/	���v���D��x���"
��'�R�'�O����O�(� )�V`xbQ��+q)p���O ���P�HK�
�ļaܜ⃈��ya�ć禅��4��dbdD|n��H�	M�$���bM`d��8ֶIp��.����'�b�'Af���i��� ����(�x�T>9�@�M�h��dLB�Ec�]k��#�%�8`FϬ~��hѧj�vc����O:R� �H�W ��b�_h�b�Y�ԔB�l�0X��OĢ}z��N�Z�.�:��""(�� ��I�<��'`�������X���VM�]�8aH<w���! �9���ޑ,��g��<�`B�����'��]>AڔI��������d bL�"�d�t@�2�@t��ITN�(�h�pk��0Q몟�'���?��ǅ�U���{%�f� �	���/5� `���m�X	`�OE?E���MLhe� ��U^ޙ�ED�
q&B��V�?ҵiQ�6m�O"#~��?r`�禔 �й�Хr��Iß����7F�g��q��<����d�#<7�I X���7� Ma���J���"���K��C�	�V���AJA�+�� Z�E[:vY�C�	`���c���0�x�#Rϻ@ȸC䉯d�n��h���>�P��3
��C� `�x�M�?=f9PtJE�AԖC��\!.5�ё1@���`��.�B䉵�6@��%��2��A�t~B�I�pc�{�`�; �ȷc��#�C䉬(��M��솚Uɦ@� ���C�	�O��I�m�`�t}+ԣF�TkjC�	*w���3%HHW�ͫ턿)��C�݆��rE�>1�A��䁎x�0C�ɸ[մ�b$��+U�Ҁ`^#@�lC�I�j�x �$C��VX��E�(C��?4t���P�c�h�` ���$B䉜l���3���$��\Y��2R�C�#��l� 1e�rP����9��C��>$-��8��ֆ,/P�M�$��C�&�`���
�	w$��dN� ��B�ɢ9VZQ�(��t�NѪC��%C�3=x���P,�|�^��q�R�B�	�YL�hBF��	��ChT�\��C�ɦE������%. U�p(�Y��C䉤�:����PY������U EC�I�:�bt���X.�-�*��(<B�ɪ/�%�n�]�h��S"�;!��C�?D>�<��	�12|�!�i��C�I�w>��b�k@����B��ƾ�i�lW��� !H��Gf�B䉉FM��'k�>mf��A�X�T��C��<��yX�k��<G�-Z�NV$C�I)h�Ht��I�7|�$\kT�Y�J��B䉁Vq�{d� �X� �j�.k�bB�	=���$L��ec��j�(L�d��x
�����
*�l�G�$v�Xh��,ǎ��fV�
28A`��!V^~eF}r���>y�%���b4H�2j�A2��-D�� 0q#㉒��lC�K���K�4O(h��������� ۗ�G(���p�Y*K�8YB"O��t遼=���j3#׏u��*���d�nV�_k�z�kN=/Z�L�EdY�!�\$1f��0?��%��x�5��#��qȆN3��u���}�<9��H$AA�t0A�e��-���z�$�8OJn\Y��4�4�"$��N��S�D+�1YY��ɂ��ɚ��UJ�=�y[6
*��[�m�2���˭ca�d�����x����J>���d%J��G�ΐK<���u�����y�	�3.*!�ް��A�KX�ЈygG�?b8�T��@'��}]�y��2j���
&�1����l��H�R%:w@mx
(��I%$�4EȐ"��C��l�UL��4�u�#Ǟ�{~�az���?qWn�7Q�z��8����'o�|���o�6�zWC\j��tq&�������dT�N�΅�I�R<lI�{�O��-�GJ����t���	�n��	�'�ܽ��!��T�Pk6.Ց7�!�E��(��9HSE�S�4&űwW әwf��zQO S�<t�� Y,�<Q#�'��x%Y31Q�]q�B�'��*@������>���R�ZLń i".��(O5�����0H��h���'t�Dʴ���"$D�w��� M�	��[:�w�ۇh�8����R����K	�1'�|��ɶ@۞#B���p�V�h��գt���ya��]^<H�&ޖ  D�4�V8��L�/E�S��[�6���+P"O�X83�=3���Q-�#}��{G/��ss��0eÊ��)�c���yC7�4b�ָs��9��D�E{&O�5 ff��sW�����B�M�7�����ɵ~[�-�c�3���r�Q�t0ը
��:F�V�O�,��k*O0QBq��72|@aaЧ?���i�%׷69��X0�T.jM҄N��PGr|i���EH���+� �St�u�$�4L>%���'j.mKDa�(<�6͒( ���^��	]���?�Rw(�;a�V!�i�<���AI�����D6:�
�C�<�2�;~�e�됈`:�����1��O�S0���c��)|a �ՑB�b��$F_<�MKn��W��Ij�Xu.}��DƔdaVI{�AO�4`Fщ�O�Sz�*�V4B�!� +�'%�h�G~���v���b�BBC2�i�#��4�h��S�~}��\+_�&��A�'p<�)㥅�BSF�(��Wj�B�O��6�W9����	ѭk5P���!_3:�h�R�g��k`Jڽ ��i�ȓ��A���F,"�,�j�4�M<Y@@I>~U>i�cQ%>�P�@L>�O�0�pP@M	�����!�����`
�脈n�����q���*��Z�LqqJD=��U̓.�(���d��S�e��E�Dd���Ͷ@d����,�#*S�D�� ��F�i���2 #&|Z�S�A�(��m��@�ޟ0`Ư�e!���Ɏi���"`y���X�G�p1��k�xɉ�e�:@��̮)�� �u��a���b��@Y��޷AWT�q�N��w�~B䉖ɨ4����6�05���V�D*ik��Z]���i�'5�������f_��(t�Xż#��4N�I�Ē	-� �	FB؟�JD$�Wxx؁�
�JU��t*Ӧc���'�����xj�G>^�va�B�B5;rqOV�Y�(�I��@
Ĥ�L�؛�ɂ�DI`�B f]�`����, ��7m^5�f@{�b��q��+ү�"dQ�4S�h�7�� ���p=��mB�:��K�YF��#$�H}�L2M�1�$�9�@��2)R��~��O��IxT� N�bU�1�K;f��͆ȓ
��\���CK]����*�L���ߵx�>���O���C?����]GMM��yg N�oTĹw�T/���bdՑ��?Id^�/�h����<��t V[��n�(��'�P�I'"����T����ӵ��ã��G�%e$ �S��,V<��"���U�ax"	 �2�f��	�~����ѫݲrS��Q��NE�b�Yo��0*�t�1M���$RP%ƽp�{��]�Աz6���WEX�C˱��dVo��5��&��#�����I�OqO�D
>.	����ʝG�B-z���y�c$$��<�S,�;L:qUe�;�A@���3{E9��{*��u��0��.J$M�LH�U��5���0�A� �!�$Z~�4�Bh�/���y�J��/�$�9��>����>�>H�wj�F�c�M�z���2�2Q�ղ,;
h����6ąቩJ/�d�UHӎ`ar�)�*8�Bh��#	�8�~0��ۧd�4��d�	����_��|��I�[��8(PZ9W��y�c�ɟ/Ғ�2.���6��ߤ$�u#>G��A�=�F���)b�T�"��-��mF�_�B�%��ūp�B1N��M�5)��7â�I�J�.ဃ�4By7,�:e`�ĕ��d�?� �E(�����BlQ91� sg
O�� `����"]����� � �	"Þ0ب�'�5��Y��~~��O8p�%l߬P��E0�E��&>��4�'��@�Éa�N�Z2JR��\��P�U�k�'��4cs+  ��أ,SJ���#��d^v7#}�f� g��8��N�Qk�i�|�<IE͟�f��]"0!ڙC��h ��<Q��	+R��)Ӆ����5�G}�<�ã΍e�h�Z�o��JI��\|�<�R��C��H��)z�9`�%�s�<9 ��H�ɒ���<�EG�V�<�_��Rf�"�$8'K�y�|U�ȓV̪�G���rYfH	�땙ge�$�ȓ$f��gMH�t���p�D�[|��ȓP��82u@�$l��9S�l��@����(�=j#()>\2�aU�y���ȓN^Ш��̈́6w�h��Æ1n1 ���^o y3�*�&Jv����ȘCa2Ԅ�_  ��@�Ԅ9&��;H��ȓ\��Q�ĭbi�C��L���ȓ8��b��M�`nQ�
�4��0�ȓx�$j���8�Ԡ�J�B�����pH��H�Z�l�8�	�$.Ф �ȓW����I�,��Q@w'V]e:Ї�:�����"ʮ
�.0��$�'^�@�ȓE_ƙIM�G&T(���;�y��}9�E(�k1��H��9N�(ą��1��Ί�VBԳ��ǳHЪ���W�	�@`ݖ: ��3�	E�,��d��/H"Y�t�ONB��Q�P�9r��ȓ�
	9C��D��̦S޵�ȓ+j$*ܭ(t��%l�G-�h�ȓ'Xְ��L�ob�P�&��]=!��*�Ҹ�KHi�x���GT�`̢���f�JH1��c�~��ŉ���ՇȓRJ�qIQ�^&Z�U@��ӓZ}��U1l��BG������ꊈ;H��|�`���޹DƢ��o�N�>u�ȓ &�UfL���7��D�r��S;�K!,�90@�]�fa�9�V��B��`3vf'ɸ9�g�р}Z��ȓb�.�P%���&�+��T�0#�(��7v�����px��%�	=(A��
����S�%B�:f�\�pN�i����m���S){f�@��B�`,�y���Z%sWE�aH��b��R��ȓO(�)�
k5�p��f�re|T��{�ViRDaPn�+�m׻��ņȓ�>�х��� ������C�"O�1,��x2�8H�q��"O
�r�f�3n�杳r��Q�T �"OR��CN����z	�?=h&�"O:��1�_�g�L�qI�`<`H�"O�y�OηK~ �㴅ڌ!F��B"OH�敎�yI�$D��\��"O��{�g҇Prt$�%z4xG"OP����4",����O%Kc �a7"Oz]y�G�ij<�`oL�s\t���"Oz�z3�,nD��#ͩAzU"O�� ^�n�(��"�bs�!��"O8`WA�gQ�!:ƦV�"ud] �"O�Y[��'��+F��?9���"Oj8#� ��:�:�p��މ:�P<��"O�P
��Ȳq
<X���(�bQ"O� �5:ch>�2�ba �Z��"O���B�J��n��Ʀ��A��4sq"O@3
weu�'��b��e�U�G�<�@�aL�ݒv�u���ˇ$C}�<y���2J�6�@u�J�W����_u�<���G7���ѵ-ʦg:��s�V�<)!��6T������:O�����SN�<�2�W�E츑���"VD�1��a�<Y��\	/k\��o�Ԭ��^�<�   @�-��aK9� a�j V�<�ƬC;P�� Q��_���Hc�P�<Y`�-�RM�w˽Y%�d@��c�<���Y5����W#������!��IԘ�I���%p��Ɵ;!��<��*#ď��tlx"B�%�!�D��=�f��q)�E�fq q��W�!�d2-��)X�,�֜�W���!�$�+mmx32�#��ڷ���4�!�ӈF���sDI�0�Rh��Q�!�d�^��M+���[Ą@��D�!�T(�M�U�)��q�7�c�!�$t��F6U� yw��)/r!򤚥@��c⇨ ZP<QG
�Cl!�9�l\Cƅ<.����LӽK1!�DR���2��=\�hp�S�ä�!�D�Xu�X�흢�D� ��p�!�$�FxJiʡT-	�,�h$��*@�!�$]��ЋM��݈� �=�!�A�:�ju��o��Xx��L,c�!���50o�I��"��Z"���N��!�DH�]�T�kE
� #DB�:�J��.�!�U=:>V(��l��h�,��LC��!�a�w�I�l(*�ib��/�!�B�-U�8J��	o��j��e�!��d/�`s�#�`Y@��'�!�\�$U
�@��^��d�R�O;V�!��ֻA|hʠ"À&��:E#!p�!��$���3�b^63�tt��a�0oC!�䞉t��	�Z�x&�Q@��N&!�$C�$���R�߫\TЈZ�`N�!�$N�v���b���o^� AB@�+C�!��SeʖLy���+mB�۔��2Z�!�������,�1=���N��W�!��<&|VMc�
/v0�\� &Q��!�$ѠLF��X�⚅L����b��V�!���!b�u���N��dd��zf!�U����q�-��!P4��bN!��3Y�l�b�?��8��Ó�!�!��^Q�5Hꀋ$�D@!%=�!�B�p���AVn�]����s�K�c�!�$HZ#��"�(j2�Jq늌I!�D\Rq�@Bbc�ys���(B�!�$��s�(��ƅ�pI�@JE�[�!�$��l5l��E� �h5 -ۤ�k�!�ė(#�����I+_(�TB�!�Ą)��=�P�C�Q����-h�!��Ao��I�Mɨc5"��ч.~!�ج_��AGc �D5#��C�y!�d�`X���,^���ʃ�L%u!��2l�.Ɉa��[��8�bEY)-y!�dG�H�&H�&.{�:H:�C�a�!�D�k 0�Gd�O嶜����>�!�bv����J�O����	q�!��/���J�{��	�[�L%!�� �Q�M�Q���	-�Dd"O��� 	�B�<l�r��0wvv�q"O�5�jΝZ��5����u\J"O�4����p��UC$�R�<s�,Y"O�� ���NKB�3��!Z\�\`�"O,��'��-g��ݙ��,MJ��r"O�q�D�Z�j}��Gʽ,8B�c�"OԸI E:�&Y+�H�B� =�S"Od�@s�� ��h�"O�ܙ7a�(��ݐ���z��xRc"OҩB��R�=ML+�e�3.���"OjȚ�ALD�4�X���|ڥ"Odh��.�
d��Q���w��	�"O�}	t$�DZ��`��ɚ,"O�����)m��x�S9d�h��d"O�93)O�f�X z���0&���"Od��"ܢ*����g#��#�(@�"O�8+�ę����rU-Ѕ=�4<�"O��Ҕd�=�^i�fɄ�&Y	�"O�(W���v�$`���&&�L�t"O)�ЄP�1��D+�B�����"O�Y刖�-�e 1�	I��!"O~�iP�E�b�
���Ab� R"O�̈w���QL��ۧ�?�� �""O<顥�
*`{�QR2�
9@����4"OJ����/fO�(+�g�9H�ћ�"O\�jȑ9�@�EI�Z�2<"�"OF���!P���btD X�V��"O�c@5�HX�rBu"HIb�"O��ȁ٤)�te
4
h��|�S"Ot��$AQ j���oW���{��|�)�;s��;tm+��C��1C�B�Ie]�@x��J�z���	�	S��B��+7�n@�N!o��M�b)m�TB��6<w�A"�ER�C������T�C�+x���S�5�G�<˨B�I���� �ƬB�.�+A��00T^C䉺-�dcP��
�P�F0��"O�Ј���hd�`�q)Ԁ:�|��"O��R� ;�����BS����"O��񒪊"Nw��yU�]�]O #u"OdT 'c�~Yi"���P��,�3"O��U-�} |˴Ò)#���T"OL0ӯ٤H���ѽ-�r�`"O�����):;�Ԓ�H�#�,#"O�!0RN/'(��- q�	�U"O ����T�O5(���^3M2�<s"O:L�,X�]ax���Ö�1��"O!��bY����+ ��"O���BɈ�4�A�+U("I� ��"O�T��%B<Bv"YZ@
WL��+�"O����)��ν�PIt`*�"Ob��3�\�f��D鞰M����"O�ਂ��hҶ�2��`�@j�"O@$DP�P����'��y���V"O�����7�z��&�a ����"O�`�U�V�C���腹q�ظ��"O�b2
۵)���(4'M�J���"OP�����w�|V�L04��[�"O��j�dC�'˴I񪎀&1 ��"OD,�5H�8��1C�@ۙPD��H"O$бŢ�5��! ��>7Xq�SO��z`�G>m���I���dp\��k8D��Y��5��1Y�AK>h�0C�F8D�� ����gB�h7fXAc^�in��"O���m�	l�8�YV��/9h�]A�'P�$Èn�*�*��\�hTp�(�&�$HC!򤒱5�h*@��J7�%iue�!��F�Q,l�G�?Z2�PQ��Ǡ !��6��8�a	 e2.�i�j�a �'��|�%B�O���xƍґu"��$V<�y$�&�� z�'عh�M[7�\"�yR���w�F�Po,NvD-��"�y���:�j��×6��r�U3�yb�Մ|��Q)`�3��ٰ�̎��y�.�J((��
�ĝ���5�y� �1s^\�6��|Ztc�H�G�<��P�E1J�S%��6ukrt�2@G�<	A�� *yY6'��Y�rFB�n�<�gE{�$�c4M
X"rFPh�<	rc�4Z�,��!��[��!�@�b�<�%�>6��ʡ&K�-v�� V�<��Hދ?"�:C'����!�ϞR�<ac��n��03�����<!ՉE�<Y���(:-�| c�]�,a��f�<�T��1n��ت��>�b af�f�<ᄍ�Bj|!b��I;eG< q`�U`�<a7瑎Z�<��u��6x�m��o�p�<��O �~D˖�]p����UXi�<!th�1�@��R��9�Z�����a�<Y�kރz�$��j�BL��ЧM\�<a��R�ƭ+���i�Ru�BP�<��+� �$:�݅Hfx�a�E�<9��L=XzZܻ��� K�D�!��B�<	�E�&[�4D����������E|�<YD&.de�a3H�w3���%��b�<��i�N�`&'
��@��[�<y��Z��ri]�)9�
�|�<��+
�Jt�� �5^]u�ƞy�<�"�Gc8I��G��LW����Xx�<��*�,���
���%\�jk��q�<�D��*HT-��%qn´�f�\t�<�!�6�|l3V�(V��Y�<I7�ʝ���afJ���"�ч͉^�<10��6��I�7�:��q0/KV�<!�'ӟJ\!7��e"���V�ZQ�<��@��nP�c��v+�lCUa�L�<at�
-� ��"GE�����ŐK�<����D��Y��K@;p80E�ZK�<����^���#��4�T�km\G�<�#ۮ|�NLӖ�Ց>(�� �w�<Q�鉎5�ĵ����'N�@� N�[�<�1*�&Z߆H�U�nW���[�<A��t�"L�4!f���s�Z�<i��b���Ѡ�'���.SZ�<��_�$&&�QaoݒI�,��C� o�<	a�fgbe��HP�<AX������<�DH��R�Y�3���C)���wg�y�<��)�R���t�X�dA\n�<!�Ҧwo0�˖扸C|�Lz���`�<ɰ�ٞ*��!Æ��c(��Y3N�\�<�� J�|�\�ؗ@�/o�h5����c�<Q"É?N<� �ɔ�b���8'�y�<A���0d��8v�O._	��`��t�<	G-Y�g�x{6��l��ؐ��s�<�e&P�o�v�Q
�fԂԒV�If�<�Ы )'�N�Yg��/�4��DZ�<YeD�/ �"�i�"3y�\��TP�<� l��@��=t�n�Ps��";>�(�"O�H!���B�����%C�}��"O�hv��=�B�a��ѵ\V| Z�"O����GۋH/�P�H�*,V�4{d"O�I�#Q� �p���R�Щc"O��C����/��Z;R@y"O<�"BA�6^z��z�,�Th�0"Ox$�7��<R�&(�Γ��չ�"O��y��8w�2Q���7mr(�K�"O��T��5�:�����G�0X4"Oʬb����EfH���oոyކu�"O<c0M� .��)H�J�Du`=J�"On��ӻC��ٻw�_j�P�"O.QP�M�kb����euM(�2�"O��a�����4Pb7�!03�P"Oȅ{��������3oڤ��"O:�����>/�4-)��ߞX1 "O���p�l����_�.q��"O��4��ȸ�����\9�"O�uJ$�X1a�q	BFۇ�x�X�"O|�����@�pFeC�t�d쓣"O q�7�Р?}*�a�%8����"OP�$�ҤM��	&��8���'�AH�B#>N��c'��!H;Q�	�'��i"D᛽S�$sjLC/�a��'��=���3f2�ؠ'�!;��i�'�0)p'�E=a�R����0b|)�'P����ƒ+�,��W�	d	.�z
�'+����I�I��o�S�֩A
�'%t�  F.m�$��Q9Ow� a	�'OfA��!�P:�A(���'V�8�GÈJ�Ĉ��Ɏ$)o�d��'���CBV�Q�$��!�Բ�A��'H<��WP�Ed�	C*�'�>�����!`=N�y3�U����$D�܈�Z9}Z����%rg�e�Ei"D��piD�'Q��)K<X�Q�5�=D���0�Rg�&����/`��b	)D�4�T6,|(*I� w�6�C�-D���NZ	J>i�G��hP &M.D��ɐ!�"=�H�� &�\1 m��9D����I�,+�(XQ`F"v�	�7�8D���p�E"^��1����:3����7D� �A��u. <�ĥ �JPB�Z7:D�,)d�M�D���8��F1 �'9D��8�@1�VR'2��3e�(�y�>S")1d�ɿ�
m�¬P��y�X#u�Tm{f��6z�%�oN��y�X,�r0���$q8$�A��4�y�A�5�-�`��E,b+j�aȞ��ybCB�3��m"��
M2�(�/�y�`�5Za�I3oԢE����Hא�y��T{3���2(����y�ݷF���K�M �F̉��yg�*2*y�ƈ�E�4�e�W�y���/#���%9s���1+F�y�nǶ(�4x)�H�@;�������y"䟾��8{�d\'ZD�����yR�xV��FIN(C�+�DĎ�y�-�d!#J	�I���J����yB�% N%����h�`ˏ<�y�n��4���
"ƼS�X��y��t�h��Ź��=1GdJ.�y2'R���Eh�Dg{E��;g�"�y
� d�b"�D'Bf�S�n�{W��;�"O*52s�ы!x$�X��ќj��$"�"OV��a�њ+_�,�3��4�� �"O���O���H-��y�$��b"O���D�i�դ��p�b�"Ole�P�E�UI�� M��z���"O<�#��Mނ��a�,��r�"O2��P�D��`X4�Ѩ{��6"O.ɳ`��ǂe�n�'`�C�"O�sG���x��!t�YPu"O�P:0O���FHa���*�>e�"O�i�VG�>ao�]sD�$@ޘP��"O���`��v�Nu�����;�"OPA���X3%T�9�&��D�h��"O��v��U4�2�M�
��H��"O����ȩ<�p����z�B "O��R"�A
E6j�K�ME�H�I��"O��9Pi,}����ҝrW.}��"O���Z.Zzd�m�ˏzE�
'"Oj���	5���y�	<84RYk�"Ont� 돘'3���aތ,�m:&"O�r�!}0���C,5�	8�"O�i�@_7&���P��"O���l��%Hz<���֛U��h"O���a��{S��T��4qF���B"ONũ$����Aw�:oːR�"O�]󧠚�V"(�:t�� i���3"O���"
C�
��y�E��(�aʑ"OT]y0�*B"��f�ڞN��f"O<<صQp� �Ԥ�!O5����"O.8�&q=�i�Ga�5�9y"Oİ(����*�^Qk&o�0""O��Id!�(q�T�Ҏ��f�f,Q4"O�yc��Q����S�s�0-�R"O8��C�{Ev9k��ӳP0�A�"O$8:`�?6kPЈ�ȢG��b"O�i苤R��4���P�]
μ
"O�@��.z���H�/�=!X��'V��zЎO%�����) ��@Y�'���ɝh���*r�.TB�'ӤMp�D� #�8b"��k��:
�'Ѩ=�a��V����,K0ȤT 	�'��Uӵ��T& �A�� $���2�'��t��k��㔝��'"->�@�'����!5�r�:0��
��U��'�xĹr%X<�h���D�l< ��'d�dxg���IȘK@�g+0���'[�	w���^L���^�X���'��%�-ڔ�#.[Զ���'���*T�� !�i��K�Nk.��'�|s�h�8�h9P*V�9�J�'wx{ k��!�έ�����6�d��'#T`�A�>�ܽs&.r�d��
�'$�6e�0c�N|9�E�X�.�z"O8,��(�!|�|-KR���r�����"O���P��T��x�TΩT���x"O�$
��3���K�ng�T*t"O&�;c�@!�8� �R4Q�~� �"O�`�����v8�����U�.p�4"O���R=��X�)F�~#:h�"O��a�ՍU��g��CA����"OԲ� �4EB�����A,�P"O4t����`�T�EM	��E"O�Y��&��,�����X*s�~=x�"O� �I�pM3t��<P�j�/i�H@"Oj}�1�Ȇ� =�1��V��Q"O��x���2��%'ʞ1y�r��"ORyj �"f�(ZI"U��2"Op��CCضtY\as���'6����"O`�aa���_�P$��9R���;�"OZ�srK]'g�h0P�$
t���"O�l��T� 5H嫒,&a�"OJ��jk3@KdD����a"O`�F�U.3њ�ا�љ4��DҠ"O�Jf�B$���8&�@M�r"O��9$�|�,����72�4��"O�P4a�=lLD��mB�"Ot���	�8N�h!.̃l�r��1"O6(h�i���Ƀ��5���x�"O:|�s���Z=������Yxi �"O��%�zU��0F;_X�Ahq"OBI�'��(1)#�"	r���"O�3�=%��l�3��xo���"O�K6et�0���@�+zT:P"Oڹ 0����ɛa΍�af�5!"OV�Ҕcъ0H�M��CO>Np@""O~��u���8��"R�%�If"O��"T�C�2����!4<��3�"ObA�W���/�,�a��G�pyj�"Ob��$��!r@v��� X���b�"O�� 'E<3���A�!)s����"O��࣎B���	_t X�"OTYB@�z�Z!q��J���k�"O��cU���T�XF�U��غ"On�0@��8H� !vgM3=HԻq"O8H`�, c��W��
v���"O􅫒�Z#Q�F��Ȟ� 'd��'��){���.`�zS@?A��9�''~l���>6>uA�OS�P=�i��'�h����:G�\�*E;PD0�"�'d����=F��k���$HF$��'�F�St��e��`h#�î8E���'�1�� ��̤$�"�Q�,���'�)���U��qHr��+����'!��zu�-[&]�agƙR����'�<i� �3��� ��S R�|m��'�H��!/� e���a��J9�E��'1 Dd
�b��D�u�*��
�'�E���<- �""J_="V
	�'�N�Z���,|���ǁ3L/���'�Z��d\�,��JtH*v��b�'�����6`��Kà�m'�!�'��y��
�z���r�K��s��=�'SJ���"�?i�ȏ:khJ|*�'JR���'Z'�(8�,C:dPX��'����+C"B��x����p&��'�<y� ���kϰQEk�dX
a��'�.���L0+Hq2tcO+d׬���'�u��0n�p��JڬV�<�
�''fI�t�Á%Y�M����9L�z�c�'�6e8�M��d1�!@E葟n\f��'D �@j�7�Z+� �`��M�
�'D��2�!�þ�[5��Z��@��'=����H:Q��y2�)�7M��1b�'�x(V��I1�	�T���b,�
�'۬ś���^�r}�4!�+;��'�p���+��1AE��(>ԕ��'�� ���UV,)�j���L���� (�H2NŁ4����-2:�C�"O,*�/Ϝ  ԰�'�W�郠"O
�b� �CaD��L�9"O�䃷���<>D�����E�$Y�U"O��E��B�x�Ɓ7I�}Ҵ"OB n�8� a��`�Vq�P��"O��9#јBo��0$�֘Ap�h(3"O�D�����:�jeM�Zj&��"O�XPB�3�J��ƙ�`�-��"O( �a��老�3��	K��"O$��!��b��ـ�H	ق`qT"O
x�W/A /3>��aEև'1�	�f"O�����0hj���cU�%��ɧ"O�Y ��)09�����G��r�"O`�z�*L���H�sGӲ8�HI{$"O�kg�Db(��[@زe~���u"O�h�@l�t��@ի��U���`"O����M�>��](4�w���"O�Ɉ��·B>I�󯃽s�~���"O*L��Ϝ�'7�t�U,�^8��"O6���]=z�XD�J�4���x`"OD��us��M01�D9ag��i"O4��f :�,��B@�50�"O�`@��y��0;,�
[8��"O\H�P.�P�i�
ԄeG��q�"O�������_��hɑ�k�!�DB�:�j%��&�_�����MT�0�!�$MȾ9آG�-��1�U]�!���|�r�Q��;b>\0�g�$�!�X�,�<$xQA�-FXi����,I�!�ɬD�80��V�V,D�����#�!�$�j�����}8,I�Ī�1Jy!���>hm���'wM\b�cG�d!���~9�|*n� )U��%\`!���^�zy�ChV�vm����є$�!�d�xxghR�[c~9�h^�`�!�$��_
����lV�;Q�/	�!�DF�<���"S��	
%�Y�O�j!���#�͙�엤-v�K��<2�!���V.䐆�&L�@��1�!�ĝ�
��e�g�J�xقB$�?�!�d�u|F,��+��3���1D��;F!�D^%eM��D	��C�$U��7m)!�� �&F��s�@�d@����y)!��Cb���_T���a	&9!�׏3&��ۅ�ٯC�"t�w-�G�!�XQ�~���k# �"��6��Q�!�>{�p�ԃK�P�����O8n!�DĩE��U�C+�S��]��(O#
Y!�D��cψ(���݆O��à��j�!򄊱 q�� �'��&��H�b���L�!�d+2�}�� F� �*}���W�!�d��WВ<x�J��ƕ��oQ�?�!��b�
�Z)�/����siѵ�!�D�K� �J�m�҅�(�>d�!��]�&��xsCUc��IAG #r�!�D©l��mʚ^������a!�_$��r3�	�z�T�����`)!�dD�S#8�P@@9+����"86&!���,O�P����:P���CC@!��>e�^����P�͸��T�9
!��D'/��+ �_��@tcg�* !�D�#m|4���0�@�h�#X!�$�E��)�m�("�0u��GD�r�!�� r���b�;�$��c�Up<�쑒"O`�2f +5JH3nO0`�!"Ohd귅Φ2$D��4Ř]�6���"O�x3f�4��u�4&a��4"OF�i�+0�T	*��
&~�!x�"O��K�ˁ�N*��P ��s:Ш6"O�a�T��G@ȰK
�p_�1c7"Ot�H�J�?��y�1͐�nQ$`��"O��'X>lK. ��B��\"J��C"O���:�T�0ba5@ q @"O�t����A�r
.M7"O��%c߿+ل�R�#����""O��I��@�y�H�P��I�`cv�b�"O�\�3f��CL���bεMZ�H�"OhZC`��B5rX�qbS���"O��rg��*t��uc�ӱ)J���"O��Â՘x���2iѺ5����d"O��#�̅�nCt0�!�M�z��"O�T�����2�n	�G�:ҸL��"O�S�� ��U:�fȤ{����3"OP�;�̑�U1Nuh�i��{�"O<�32B�}ۺD��L#Ol��4"O��y�jЧ.��QU-�Q�r��"Od]����@��sU�F3g�|��""OR�ʕ��t� � &ń5j����"Odљ�a�_$dk'��0g���d"Odq�!�(��jTaS���"Oq�sB�k�l Gj߇dc@Y��"OL�Td��vn����U`t¡"Of�B�dKFO�$�LL�UB>5Y�"O�u���X���+���,:�"ON me`'ʢ��\zR�r�<��\8B6������HR"@SB�<iE�L#��0�%]�B����o�h�<�D�Y[��窃g��!a�C\�<!��*Wx�01 ӻ2OB�!��Q�<�G��s�ʸ3�C vcl���\O�<Q�']*��Z�g\��luH��f�<I��ٛp�j��ChG2{�x�� ��|�<�F8OWD�1�Ϩ�x���l�<�A�Z��N�E ɧA8���b�<�b	D�[H���
�*,l�#�$�g�<���G�E1�'B�,C��+��Ca�<!��kU�ԚO�&X��-��_�!��c�A�E���4����̔":c!��8'd}H�G9�*0���.g!�A.J��`��0���CC�[�f!�DN.-����J޸�A/�/Q!�DǗH�
qB����޴����q�!�dA�h��D��R�0��7���!�
�W�@���-�'��!5����!�Q"Jbڽqba��Y�v݉!Mȳ�!�d�8n�Ny���M��Li�`k_�!�d	�fx}�&���T}�@B�@�8�!�Dʨ�$	hUOB�^> �$�&
�!��я�x0���&$[l(;%eQ�b�!��>v[x�!�JWL~t� �Щ;�!�P�z�(%¦���?6�ɕ�R��!�䒕9s(Ī���n?���Ƅ�!�$�4N?b���g!�U� �&!�Ĕ Y�D��5B���<�!�d������S�Ƅ$��kW�Ɩ-�!�Ū0E��t��]#R�x&�a�!�d�#[v��Baᖢ3������c!�� ���*h�!�%i�~���"OR���<K�:i@'��z�A�"O�0j#.�wP�Q��/1��%S�"O�$����6V�Գ��X�&��"Ot���E�bƞ)���O0��
+�!�d,�����%�� �T�#�!�D�-�e��!�Uo`�Q%�2�!�*Ii8��W�͵
n���1�"O�}�Ш\ &STp9eǝ!|��3"O�̃Q�� e��T��fˑKr��"ORY���-}~��B�R�|W,(�4"O8��r{�*yP��<AMXm�""O���.��[����b'���0�"O�``��*"
y� B��v�!"O�����I-P�}고��EP���u"OU·8o#*�
E�F?�h�"O�9�p�-:�� �5H���"Ol	Фa��G2d@�q
�5?2>���"O��9g��<'¨��'���J�5H2"O�E8l��=Z�1�D��47�,�5"O��ҥ؄I=��UHϲQ	��cu"O*��GNT�M< ��FA�F	>a0!"O4}�Ti��b��|J���W�P�`"O`�Ñ�����sJ�6T����"O^MJ �MY�D���z���S"O���Q�@�O��<�'%ıL42���"O qT*�or�@`��W-(+�e�%"O�$�A@�)E>ɚ��H�L�Y�"O�0"!&�2{���j٢԰�`"O��J��~�3	^.T�.�Q�"O~5�uM�E�V��ǡί����E"O
��q���6��s3$�H� v"OD�rr'���������SJ��+�"O�;"��5�$��6c�;��Q�"O�1��a�j��$�ϧ"6�P�G"O`ܻ�.6��(�"Gִm3J��"OΑH3ǚ7nZf�Kr@�/��I@"Or��I�Y��ł�D-��b"O��#A�N�2EFxxp%
X��E��"O�����ݷ\�(���Ť6��5"O�$!�N�>F5s���F뀜[�"OƕUE�M<6	JR�U�u�H��"O�`w����1���yf�cA"O�8��ʚ �VqQ!�v@�P�2"O��Qp�T
���!.�y>�u�g"O�c��G����Oޯ6���"O�]����*E߂	�B���xC"O.�rFE�5�nhbA�S�Șg"O�l �J^4S�t C��J�0��"OH �t��X�� �"mҸ^�"��"O|�Y�/ɁP�$Ȃ�����}�R"O��q��=���C��*q��i0"Oq@Q%�\��N&=�&�`"O~-klP�	�nI��	�<����"Ol��`��L�hvhG�\fJ	R�"O�M���#R4�(�lЋ�~]H�"O��I�.��'��p��Ŝ/�bq�P"O��� ��U�B�	3�O�[K*�0""OFDU%E}�4,)t�<WA2�U"O&���S�(話4�W0K�j�"O���Ƨ97V��7��'/� bg"O���fE� �,D"ӨP{f�1j "O��s ^'(?���'(��Msp�``"O���v���EO��+��S�KT�9��"O� ��ʂ��4RV�@Swi�F0)SD"O���� �Fb�ݻ��%3�C�"O�W��-�ZKj�b��"O�YJ#G��!� ��D�8Q�V"O�f��I���0§ܝk#�"O4�z$�F���p�T�_$Iv%�C"O4�9��¥|lvI�6fM�O ��"OrI6�V��B��G �5c7"O���D�̘�<����lP"O�0ha14��+4�ٓ���2"O���b,Mh~�T�ɏ]��� "O��q �c�� ���0�.�p�"O���6�
3z �X�x&� S"ODQ�7ϔt��y�S�Ҝ� Q��"O��*^6�� �%Z4G�H%��"O�U��P�pu��)Q�Y')0��j�"O�!���%Pu�@�Q�}w@ɔ"O��x�͓�wG�4�$O%����"O�аևU�Xi���#�6�f$h�"O�HBt�#{@t��ӂV/K!��p"O�TД�/]3؄����.� ��"O�0��!YT������S�D�;�"Od����.b�H%���]��"O�Ir+�'A����fb�1��b"Ox����"_\!�0�����R"O��P ��.	q���D ���\�A"O� �5*٬�"�HvC��F=#�"O��"� [�
��H��~�&���"Oz���M� ��dB7S�H��"O�qi��M�R1��� 8pmYQ"O,@:�M�O���� �|�
q�"O@\�a,��5� �J&.'�T�a�"OV��&KYRiNYCQ�N
\�X�"O8�1 ZX�&���"�T*�"O>��)��Z>��'Q�nɬ��7"O�5���M�;W��`�V�K�r%��"O�H�0�T�(�԰���I����{6"O��{��O4�F�`�"��l�pQz�"O�9�O>t�\k�G�&/��} E"O�I+�� ���S�C�d�����"O� Bgm�p޲�9�Ύ�$�H,�D"O��C��T���ǴmN�<�"OJٹ�Ȇ�}G"T����)��#�"O�%�4�AXI�IR&�kyV�;�"O���ueZ�G�ȥ�1�,wYz��%"On��aDC�x���{�iW='M���G"O���LDS0��̀N�"a)W"Ol�;Ql�:;�����dܫZϐTrg"O=�q��Wc���PC��|�Ҵ�f"O���A�¬sO���E���R� "O��a*�hFbi c��+���['"O0!8gFS�V��� �xx@!"O�|����sc��{�&�49�"O"y���j���Lˢ�n�B3"O�ѐ#��=w��q�'�̙��uCP"OvĂ��q5��D >�%�q"Ov�w�D� z�y3EjM�O��Hb"O0Mɐ�A�Zq�Q��E�pچ�1"O�Y�i�y��eAUjr��4"OL��%X�;�+I�^��@U��t�<��C�TI"0��.R
B��,+��s�<9fˉ5�L��4�{� ۱MPp�<�UMN6l�Ĉ��A��w�R]i�b�j�< ��*2LE�IּH����[j�<� ��C&Ʈk۔�e��-r�b��"O��Q�O\�>0��*d,ؑ!�L�r"O�T�BO_�'=�Ż���gaީ�p"Oܩ�6�Ag��	S|�A"�"O��ĹK��4���6^�A+�"O���uaP�$tlx0̏�&t)�"OR}PP΅`���Q��{��"O�л��K�l��0�,�. ���"O.=�2�R�U�� �s�F)��cHP�<Q�@,\$my��A��D�E$Dh�<	qc#T2L GH�6���1��g�<��I�A����Y�Gh��R �KZ�<�b��t�t�V��b4i�-\�<UG�v�ҕ��M� X���"\T�<���
,,��!��353��X�Qh�<�`k�H��I�0C�G^r] ��x�<���\� �x�2���S*iP���u�<��C�G��4J��-��d�n�<W�X�9�z9�҃S��*��&E�k�<��Œs����h�����
�e�<�V��] dKêT�<�� �d�<QWH]%�d Q-؝5B��r��F�<���1P�,a���Tb�b��<yd�mf�-6�ܺy}���VbVA�<1�M�"�R�1p)S?���c�a�<�ף��gX�ص%� 8��TI�(	^�<Qs�(*Ѩ��u�B�
������]�<Ѵk���8,"��j\��D�PU�<���F>kH�U��N�?ǀk��i�<yt��x�}��O�0r$�)�{�<ɣOV&#\�y8��ȅ� I!-�x�<a��U=x�D���3��`��r�<Yt�üCVhC���k\��toKo�<��!
@��*b�F�;���Hp��P�<����X��T���ē#��P��ZJ�<���!Ɓ:Ń��p�
<Pu��F�<a�![�N�0��V��7
�[�$�J�<�юT70��X)MP5L>����VF�<� G�3.	9�ʐ]qt����l�<�!��pl��1$� ��B�Ėq�<QQ��=,��I�sG�\��ia��NG�<e��N�vh��m�"�k�<�'��,N1D�A�j����c�<a�gT�i���b@�M��bW#�G�<a�,
�%��\��o@�QE�z��A�<)bF�M�m;V'�Cr�8�+V�<Iu恛=Dу�ƻ���t;�B�I4_���
fV�>S�)�w�TC�I8.�a�^,amE뒊��DC�	Ld�8���m􌛇!�	<ӦB�		Y�LDb��3�t䳶�R��^B�	�AGL�J�O@��d��w�C�ɣ4ߎԀ���F���Cӏ��PC�I�}�n\�rIF�s��3�hM�(�"C�I*R:��C� ����Ua�R�jh��t0����R5l�A����J���ȓf�d��A�IE�Htd\� ��j��EH�H/NZ� G�V:�q�ȓp�X́Ŧ�#о�b�\6(9��ȓ&{L ��@"[�LY� �B�lx��V�0�ӊ2=y�� я�:&�u��w�v��Р�%O5�e m�#cm����7hn� ƀۼ/4: �C���F�ȓL�
}�T�6}��q��G�x�,��S�? ���T)>P��Dq/Al��"Oh�:4㝫+���d4Ш�"O8�cF��1lp1�Vl-q h�"O�	����"=�@EK������"OL��#��*2��]���y��P�"O��HV����9[�J�NtC�"O�����3r�v	"S�޳~u�ES�"O��fN-#	JD�M�@�5"OJ��"艙YC�Х�8�2��V"OjуD��LM�!a���1	���B"OƜ�`��'7�0��V!��3�����"O���E=D݂��A��V��M+ "OZ�!5��2�
�Ҧ0��I �"Oꡪ�ǸR�d�p ��#F�R�	�"O��P��9 ZZ 	Ѝ�#F�p��0"O�Q�"�
/�0�1M���h��"OD��. �;�`\��eV)�(�c"O�9�6� o��mr�ƼO�(̓%"O֥Z���4L1(�"�b�9YD� �"O��@��`[l�`��M�9(�e"O�A���
�0��f�Z?H+ �d"O� HK�	k]Xl#��zo�ݛ�"O���&��c(�hٴ�Q�jc\�A"OZ`� �n:^�� j��Kb��a"O�D����]ul�`IF�`��8�"O���F͋eH`c��8�@� D"O
}31���^����)U���Kg"O��@7e�'��A���E�)OHye"O���!��D'B�z��R�x�L��T"O���fT�`���c�*�/F����"O�`�pcՀb���ǅ5M�z�x�<��A��/� ��A,K��5�U"Us�<�U�.=�JX�r���H
`��i�k�<��씋[a�b5�� iQ����i�<1e�O�n�n�FgĖxn�����e�<�l��<�$T ��*,���cKd�<ᖋ_�P̀d�J�o��+���H�<��΍-,�A�O� �6�r��~�<I�U�s{$tG_�L�z�ⴀt�<����|�b�sD�L>l0��B/Ge�<a�]�t���I�,�c��Pl�<���^�<���L;L�)�#.[_�<�����$�X��<"���!v�N]�<�W'<H,��1�+9$��!�\�<�v�d6TJg��?�}!T�V�<�c��	�,S4�_�;���
��U�<I�Ś�~ �L��`P9w�.�JA��P�<q%��*�����87�5�5�XH�<)� ��l��i����k=��xQ�Gn�<��I'��[U-�?[�������h�<��$=b����iY�R�>Y���p�<� jT$��5�7OG.\�G��a�<A����V�$P�Q��Nx����	`�<s��*f��e	ͳq�|�����p�<q�EҜ <��2_�sц\b�eRs�<�B��=	1��;�W:���b�V�<�`�Nc�.��f �LR�h�" Q�<�F�ɩ,�<i�i@��5���J�<&���M���edŮ@�<P��N�<��l�$}$�ۡ�Օ��T��t�<A�"��N���J�h�D�X���Z�<	�Lu�&�j��ڿI ����Q�<Ѳ��W���x�眲v]�(G�I�<�%mD�*�;�W�`��i�G� B�<� �<Z��@v��9 �֭Ktы�"OX��s�MRw��P�������"O�M�	Ɵ*��Hsf��/��t�"O옃�&�x4�P����S���"�"O�9���Y3�h�m�pz���"O��0�u�$U�w��[xB$�C"O&� t�T�"�����%T�� "O�T�ҁq��]B��UF����"O�$��5DY��1�R0q�씲�"O<e�6h� x�4�����90g:�K�"O����j߁u���c��w���"O�����e� 4r���Ha��k�"O�bSB`a���P�:����B��!�D��h6Q��Nʦ����J�~m!�ݓD��͹����T��PhrR!�d��T�AB�֟sp6��BH@�~�!�DD=P��)�
�NQ��!��!��B�3�Ν��TJ HC���a!��� v��aasH=���qn�&\!��R�hplWcP�=I��[0���`Q!��
�~� ��J�7�r�l�<L8!�ֹ��	�	.H(2��N-�!�81����'0�l��T�z!򄂾���g�4RD���E�=J!��Y,-\��a�@RP�ͪ�Ş@!�$A9���d�Wt��@3]64(!�$S���P�# �X͚1��kw!�$_�6����&��BES��@�=;!�ď'\��!3$ �s�P�`돨4!��I!��!��$4<�C��A�!��~���ߦU��S�ŘWb!�$ۈ64�x@�Ag&���4��:�!�D &Yx�9@G��Y�h�+�F��Y�!�M=I���Ib$�+�v;�N�K�!�dF>��)��Lv��T�W�!��
�q���7o$3{�=GD��Fu!���i���@7�5�����9!�d�6�>�S�N*/����!�D
�E�
�h�5[��x#���!�D���Q��憖=��aR���	�!��K�I�4�]x�<�	�-S��!���8HQi)g29(q-�z�!���qa~�Q%�_�YNX���G)Y!�d�i�� #$�V-��di�d� �Py��_�<�*2�^#4���Qb)��y��N
3��� ��*4��%��JD?�y����29Z'[&)D��cV��-�y�>��U"�a��P:1K�'��y�k��Z`�h��C�2^��8� D���1�=ˠm�Rᗍ���Ӈ(D��HgCt�R��3=|�sb�1D�d`�ˢ>�F��&$=�h �fD,D��*�8T�s7d�e�fܒ#8D�x����+��E�s�r�D ��7D�ZB�7P0���r�
���9D�
5��_��,c��8g�X�E=D��(�
]=wE�Ia �K�_<����";D��ѱ!˷~�`�wi
�DQ(Q�ӊ6D�q3$+�ݢ`�]o��<�@'D����֮\v
����4w"����$D�@��̞#f��B��\c��"D�H�j��P�  ]�x�u+D�d�anяr�K��*
Te�(D��2 ��.�ZU�fG �qft�QV/'D�� D��D�X�&������ݛr��Q"ON�a���1��չfmH���S�"OD�`��r*�z7M��*q|i"O�Yb�FI0Q�x!�CL��|oT�� "O� Uj�3s�l��d*.3}���"OA��c�!q�!Z�H��q�ٳE"O��Ef�g�,�f�?"\*,��"O
��S�N �и����N�8"OJ�J���%	����um��̢�"O��#��yN	����!UZ��"O^ɛ�O0 ����+�9'"O֘!3��H$!��̯�h���"O:4AТR� f��HрBE��x "O�X�-մa�R��)�	EDɘ�"O�q��&Y!`�t\���ߎ_
$���"Op�#V�&n8�;��ر���	7"Ob�bVU�{X����'�=/؞dP�"Of�HQ+��S�DQ%�]Ԍ�#�"O0Ҏ�^
$��I��g� a�4"O���5Q0�vp2&
�"�4��"O��Q��xP�³I��a�^�"OZ�aq"�0�bi�NP(OȆ�"O��[7�W#g)�|À�R6M�p!�!"ORxÅ�V����0Q�޼d�X`G"O(U�6����듏;�>���"OzE�-���U�� Y�P�`�P"O>�s���<M�$93U`G~�֑
v"O8�E�|X�h!b,ʂ#�D�X�"O��s��Y�y�)ؔPe`�9g"O欙�%M�X�~ј6)�j�(
"O}zfb�3�,D;��;�d�CG"O�M��/��\���?|�1�"O�\� C�vKp�:G ��:pF��g"O�����Q4m��P�N��nY^,��"O���f�asڐ:`B�:����"O��á>�E֊$���'�l�@�n�-�,���J�Y㊑��'�2=1��Ň)H��GƖ3W��	��'��p����*vr���Uf΀���'�U���E�/(5`�[#�h��'\i�U�\)3p��N�	!�$Ii�'�����y��e3�/U�0�\��'�����=&�y�U8!��`��'fޠۓmJ�A�]1�� Kz x�'xݪ$��1�n����W27�����'`��+ٱq�<b�)_�E�^tc�'6��`��z�~m���:EY�8
�'v̔Z��E7n�� B���9LnMx	�'��9�!õ��  pe EAp	�'��(�6�ϒ�T�WkG=*<	"�'�U�E%�,�)[�;P��S�'��Z���2"��� X���=
�'y}D�7]m�a'I*,i�
�'�2a��I�}E�ٱ	H/V6ؼC	�'��t�WV�*$6�*V�4%��'Ŏ��C=$w�X�GＨ�',�D��Q�e�N{�fN3m��J
�'�B�:d�هD��J��p�p��'v��rM�^�X�2 T��
�'-�̀0K��"�tA��^�`�n��	�'���T/�p8��L���vy�'cY geցG�	g�M�I���'2b����x�cŅ�>��E)
�'�%f��)�@�c�D�/1Z��
��� ,��6F��L�:��g�#J�Tf"O���Ԉ��y��P��E �܈�Z�"O�=�F��Q8&������I�$"O�|a$�[��1eD�HѰp��"O,��V*@���3^�;*��d"O�(�'�T0^�3g���2`|%"O���nJ�M �8�M�q�"��"O�@'��`v�� �?~�d�p"Od�a�@S._��i)�CZ�Or�H�"O&���ˍ6� eX�!�W�i�"O���a���x�u��чk�RY1�"O�)qB@t������٨;���"O�ـ���^P0��1f��G�N��"O M#���>���6�Z��"O���h�0HW��s�X�Etܙ"Or��kc׾��C�����"Ov8{�`RJ���XD+�C;����"O�AM<�|ȹ�KڡQ9��p@"O��!3K������N�|�rG"O���b
>1��̱�/�	^���W"O�IpEM\��YGɏ����"OH���l_j0[ҍΧӼ0z�"O�980��g�F�2�gM�{b��ZP"O��`��hH��)caR�,\�p�s"O���,��Pئ��pm�x�p�{�"O��A���-F\J���e�$��"O����Z�)8�����/"��+d"O��ɠOҟ!��bM�&���"O���!�/k�L�p�˕5+�ݲw"O�|���ݯn�)�G�0a�0� "O�Y�G$_���8�v�M6�Du!!"O�9J�Q�F�� �0yJ�x"O�L� %K8ҩ��-=@>�Yzb"OT�p�k��a����Z4�E&"O�p����4O�!{�-p�e"O�S��8��}����B*�J�"O��Ð�N�#b6\�#�%F�4a�"OL�1��=�����T8C�*��"OLma���LLc�K�����{`"Otm��T���Ѹ���H��!�&"O�ʒAܲ� �قA$�.D:�"O\h��0�X �4�ѓ%rv|�c"O�iǘ�!L�1S�Ņ11ŮT��"O|i`���:~=���B� ��Q"O:���4Y��;�BY�b���`�"O�H��Q�0Ƣ�ڱ �#�6�r�"O��9sꈋ\L�@� �O�7"��ڀ"O0aS�	��@�;�H�0J�2���"OC���1>���g���b��"Oe0�����:�G��O�8%�"O�P�D�;3��Ii3�l�n�;�"O����mǹg�l�p�ϓ�Ɲ�"O\�Q�L�X�*��X;;���9e"O��ʶ*^-��l����hH��"ONm�2U�N���ԟM&<��"O=`��N�X%T�i����"Ȏõ���+�q���ĢmS�"Oh�
�c�#��E��W�B�4d�t"O��[q@'��i�TChJE�"O �e(N�x�{G���r`!�&Ze��U �"1���*�@x!���2Ӡ��ڔ�
�s�kR1sj�B䉀q9�ucك~��<��!�dB�I�mG��x�ɀ�u]|c���)�DB�)� �]
F���v���"bd��Җ)[�"OВWğ4�N��	�
��T�"O�t&bO�br�p裉�U����@"O5��̄�-���gB��1*"O�и�B�,Ct"���$O�șE"O<�⍗:_���Ë�2��0b@"O���� ���񲐌�~�~���"O�S�GR�M:�����~ò��"Oĸ�(S�`��#.$�� �g"O��R���4nHT��A�,mޖ$��"O�$J�
1~'� ���A����"OB��B�V2]b���f�Mz�.���"O�%g �Jmc��� �6%��"O<�{�@�{�EI����2��t��"O��l�O�	;�`<�P 3"O%�pK�И��ͯ	}���"OJ���V"Vll3'Go���"O
SG��:�L�w�50V���"O��#5B7<|,�@B��-��"O8�x򉌐/�^�¤�R�<�~Ap�"OH���F=��B%ǉ�|��:�"O((��ˆ36l1�W&���6��"O��"h���g�Q�y�\-��"OPySs�]�3���39��iI�"Ǒ1��j���cr��g����"O��b�!3��څ�
�]�88��"O�(u*G/w������t��c"Opq�q�P��ɗ<=(ŀt�V71i!��n�>��dZ�9��7�޹3]!��08\���]*B�� N�M!�d_���LJ*8� �\E!�D�o�Փ�U��T@�͝�?[!��C�c�rqIT �3>�ȅAL
�T�!�d��$.|��e�!0�,����r�!���Q�ԓ1HP���숢	!�$F��L4H󉏞x/Z� ��
 !�䇡A5�X�+��{��$r�J��R�!�$ �w-�� �d��w�U+PD��U�!�[�@	 �8}?�X��#)a!��h}~���c"���u�<;!�$ZN��l�c � g��I��`O!��{����QN�;Z�v����[2#!��f�5��m'���B�[!��&�P��_8(�t	䀒!6�!�d=q9��"�k�5t`��X�a��/[!�
5x#��GmJ�KF&�y6 �0C�!�$�%�j�����x2��ɇ�Hi�!��&>���*�/c��ui���8�!�3 e�S�G.$�B�� "�. !��j���H1�֌"�d剱�>q�!�[�����ƎH��`(�蛂zv!�0Wd "�èb�h�
$}!�$�6�C ��S��H�a�A�!�䙭o�t�+� K�P��٠7�#z!�$�*G�D0tG��z�����!�7���s�ݦU�ꍠ ��t���߃�Б�o�k� ����,�yA	��d�J�K<񶵸qB�y2mW7�~ `q�]9m��
��M�yBgV�Dp6IdI;�A�1��y��V6|��U��/����I�	�yR� �z��;C&H7RXz�	
�yR�]�u:�KǬu�逃�ڔ�yK�&��9�R.�� ��P�C�Q��y
� ����Z�*��"E0y��f"O���`��~$e����2��A�"Ov���	L�0k�X���L�Vע�!�"O����+$�p+d
\�7�
9�$"O�1�G��(��[a�K:p�s�"O�l��dΞ��)CBM�i(<�{�"O�k��M/<�P`�;F�z)y�"O��k�	�[x�1KE��54�H��"O2�z�)Y#}�$(�m�J/}�E"OҀˢEE[�\B��^2D|��"OJm�VO2 7�Z�)� H.��j"O`)�0�C�F�c�Բ~{�)�u"OdH3֠��M�����E��:x�"O��3�[�owL((ԄE�u�����"O�l�E��!���C�P�:Q"Ot,�p��L3�	�nH�$�h8��"O΍۴-��i�@2un�=���'"O�5!��Gq������O(�2"O@��A�ӯtr�-�U�̜8�4�"O��u۠I��yB�!C)"���q"O��UGA,�0�j�a�:!쨄�C"O�� !�
@)D�
=�2�"OZY����	Al�������v=�E"O� "s[�lDBD� ���e�h��"O�xAt�M	<Dp	R5Z��H�"O���D�$o��A8C.�+��ɹ "OJTA�Fң~�R�L:U�:�	�"OTTj��ʐw�R�2BR�4���"O�Mѓ���n]�NJ�A����"O������t��9��@�_qdH��"O�u��m]���4l��!�V�;p"O�E�SF�)e<����[W�>DxU"OJ1p#D
�y1�� �8��$J"Op�������؀�ρ5E�t�Ie�|��'~S*��q@�h
T�W,`���'ۊ|��,:b:I���j}��'�@K�	����䆻��ur	�'Mt(�iU+W[ E�L��m$9��'�Zx��������HzU�5����'�>��
�� � _rN��6@�N�B�	2-�4��K�1%W^��2`#x.B�I� �
yUA6k^
�	�jТPf�B��U,�6+��k&�0��
Ӯ	��B�"�N���Đ;�I����+��C�ɩp~(Aq��'5��S���Rf�C�I9,5�PSKN�8b�p&��e�VC䉋8*�u�r�^���-!t��;�$C�;N����Z��j q����J�C�g�h��F
�q�F�ۣ��Xh�C�	%	����g(�-�L�k�+���B�I�0�ʬ��'7.Fu�$Ɲ!���?و�	@�*����.'�̵�B�4?C!�d2`�f`���ɽT�Ԅi�L!�$ܷbDf��(C�O��A���4!�d[�z�4���%�.�ʴ�ól!�$N�(Z�5��Ŋ*zт=kl]�w�!���4������/)�Ji�l�5�!�$eR����8E��-��KP+h��IZ���O�bA�9B�ʁ���D�`����N.�y�ņ�� :s#�=O ș�����y��S�u~9@6 �83�(�S*݊�y�G�!0j鹰J=\�Z�#2�֎�ybmϼJ��K�\�M�ñ����yrF�tt��ѳ6��3P���y
� bС��Q�֘%�(����vU�$ZS�)�S��f��e"r9�$�܈n��Tm@��y�lE�g�tdL�nO��8��K:�HO(��U�gf�&}����U�o�!�3����O��@`{5F˓k�XШO���M��E~��b�
	:�+��)�R���ń�y��)\�Rtw&ۈ-�RpbA���~�'������D�,h"�C�5;�'�4�
���'C�tR�3N���#�'v��%��&9j02��Y�7v�]X�'��3�悿�4����@y��z�'���k��=,$�A��P�A�,	�'��sA��:<xC�˻8���y�Q:m��q�R�M�S���9sj���y�[<����@n]-QM,��b�W�y���2q���i�C
�Iچ���f�;�y�@���:�BDY�.��� 7�y�G�y�T4�ġ'{��hb���yJ	���}0w�Ct!ɦ'���y2�� p=��6�B}�X��%���yB�EI� (��.�g���/׌�y"�
�����4��`C6%8����y2IQ�O�����Ī@������M#�y�f�,�1�F-��d�CeA�y۷b3rÃӶym�ԙ�����y�g�J�I�ƥ�(l{�AkU����y�雦'U�{�J�N���H��Ά�y�(A���H�IC�H{*�0�j��y@�?3V� ��
OH�DƑ6�yҁ��ko��-�1�x�ԬS�yB��Cz��R�*�	�.�H����yB���*���82�bEdP����C�I�W6ry8�OK�k,�l��jʴ|�C�	;,��ё�i�$)�K�l�N�C䉅�hk��ի@S�	b��ܡ򤖻 ��|s�+̩EZ� $֔+K!��H�Dh|����
z�����*f8!�$Ƹ�(�@��_$�jp�I?88!���*���(y��#G��s��ɷ"O|�hG�im@<�䦒��x��"OF��e�_*�,]��g�K	�\��"O�c�T#j�B��F4}�"O2�q��_qj+g���Y,��"O���l\�c�½�8a)���q"O�m;��YZ��b�A5*��k"OT)��B$��Y�nP�l�(�"OL�`�4����^u�B���3�yb��D�Ңň�oN�F��y���La�A
�l2YqT��y��j�l�vk�D�"3�`]��yBBÃ?�jAA������E�y�m>DY��+k�@��X4�yr�q��=!S˦�tH
�G�y��$�,E{bv��pt&��y��.m�D�у�u3$�ғ$�y��*2�H�x��_8o�2�P�j	6�y��.H�T5)eT+aD~�Bfӆ�y�g��	�*h� Ѱp����B�y���n�Ш���C�-�� �yi�	~���1�<����<�ybÝ�'��0�GŻ,���[��1�ybnU m��H��q&�4��?�y���*7��J@H�>a����� �y��9ԑ�0 ��D�p�#���y
� �G��;�d撲\xؘ W"O�H���[}�0�%L�
\b,�@"O��"D�*���b�.y�Z�k3"O��4e͉f0l�7�S4clГ"O^��bnB�T6Q+�cA)d4�q�"O���5k |�V}�"ȝB�4]��"OdHsSJΠz�NL����:��7"O�<9%W2Zb��שӝz�H�1@"ON-r3G( ��=�S��,����!"Oࡁ�R ��D@�����r"O]���0E�a����E>���"OTD�

<+�(9Z�&	;AZP`"OxM��D&B�"�_%nW�BT"O��8sB	������q><|`2"O$ S� �����e��wl<"O�	@�b����҂8ht"O�Q`�iԆ<+��8`˞�J�"O%8�+[)8�^|R�l��/�L4H�"O��Z�N�;*���	g�N� "Or�pW	�2l�!L�f1hM�1"O��j���J����R�7���"O$�+F'F����B&V5�,u�b"Oΐ�e*)x�(D�CL�
Jx�"Ofȷ��$#_�i���0~G���"O��r$��p=��B�ݦO�f��D"O�9���}�&%q�W"9��:s"O��
äU
<C&����-^��8f"O굈�.C�9T9���Y���@"OZ)��a�%�`}�7ݒ`o�<��"O p�`�[�b����q ��Slu��"O�P�V%�#'F-3���`��"O`��gI`�SōI-6�
��P"OX�:6�B`��=;��Q<
���1�"O�`�n�1�s��?"��5*�"O@l��.�e�>P!.��
��a��"O2bs��.��ѡ� <��	�F"O�%�ƎJ�}�b�q��T�,~�ZT"O ����۝%jP��1��dr��kw"O�Z����BA�1_H0C�Ð7M�!�D�s���1Ԥ��m<�˅���O�!�D�r�����M8� B���)�!���t�8A��(͓Jń���Y6?�!��� �d����ZI�Q�
^!��\�T�sL��:`����k[!��$>A�p�J3\��4����!��W73Zr���B�(ň��Ãi�!�DP&8�	D0%�L�Y��N=h!�ޙ:X*��w�M�	�^M!Ũ��NS!�c���sf��04	����(9(!�df�&�0��/rD!�]�J�!��U���]ۥ��%(JE�ek�v!�����B�ϊF��v��gS!򤊅wE��Gӹ?�*T�ZQ!�d^!v��A�1���lxdX�2N!�d�fU8 �kI5!�b(aco�3!�Ć�­�цK�-���0Ïo}��c4w�~����8vJb��ߨD�v�����.ZB䉻<�j0C�E��<:v� ��3un>B�I�9��Q#B
�$]����H6tx�B�9�fi%(A*���q��Z�fC�B�ɞ	�~pS�(
�R�ҥ+�G:Z�B䉌`Bƨ�Q��$9�7�Y�P�B�	H@�)�"k킁�p�
�?�.C䉢M(N=�r�ApVHsL2�8C�)� 8<���Ǧ�!ܜoT&@&"OP�ڦ��'��a��`]�'� l�g"O�`r�N;|nlQ�������"O��8d,�����P�kD�p�"OL�3,��8�H1F��e�v�"O"�A㇭>v ����"{�9�"O��C4p����D��z��֋Y�<I�O�vt�$kϽ�L��Ӣ�[�<' *v���z�
K�k�<pU�Lo�<yrB��1čx6o\�?s����h�<� �!h��h"u���T�ػ=�!�/ngP�t��$��ebQ�C�!�$N��~����ΈX��<Y��ߊ����4����c�Dbq݆M8U�ȓ�V����Tyu��#RAQ
 ��ȓj�0� Čݕ1���0O\)�䤅�!�����I� &�T�W]\!��I����b㉢_}|x�3㎋�\Ԅȓ^~�8C���1r�Ai���z�4Y����5���� �cߴ\�Έ��:Hd܀��.5�$��d�.K�)��I����&o�3
�b@��M��@�Ĝ	���L,�T�5+/�vi�ȓU�T�"%�gw^,�@��@odT��)�\0��"[�Jr˓}��Hvˌ�m��T�[��"1��	5n[����J�#~��AKV@�-�c��y
�SAl�%@����Fܚ�B�H���0{�mU�j�rm�>Qu�Z<]�aK��!�`���)�)�	{aJ,P�nBF�B�!�m�]�!�,��Q�A�#V*4P��	be>���_���-� %��d��0v��I}2�*y`fEk$�H�}��8"��y��a����L	$��q��'*��k_<��|� "H�ex��c��m�'�|YR�_=x �baMY(f�8��	ϓz$�B!�)e�4��q$f�T�Vy#�m���R!\��鑡�@$�d]��S�A��(
�4�a�S��=u&�$�$� ��y�"T8��ʹK�Y��^#tlx��^>�*��ݗ`�(�JPi���8���G"D�`�e��v�(퐧ğ�z�`j��_��)���}B�
�' !�(d�}�C �Q�n��m4<a�@����[T\<��dV6  �[�8Y���w		�$�
�� �ha�-F(A����Vl��0@�gڑ�8���_�W�^���d�+k������:O\5b���v��mZBo�n��7F�2nV��w�o�Pr �qk�0�^_<�U)�lD��kVB+/�d�2�mG�s\�O��%*[��X6�I�u�\�1u�Q�X���0�@�~�D/�Fٮܡ��� m�`Hi�<�3 ]�"C��R � &l���[�G��;
�}p�Ĉ*�H�&���~�������]�{Ȥ�;sg8ivJ��`��1s��
����v�Ε!��l+�,B7�AUf,Yy�-_��L`ن��q	�1�f��a��a*�	�o,��@@�Sk1O�����ڳ&^0p�@_n�
�9�퉯&'�y��̉�:��~�I+�}VTT�਄:mzF�ц�A%�zh
g	�	�D����l;X
1��fX���d�L�EUb��R�كU~��B쓨K�hA�V/�)h��*�(�ڄ@�CYt��� �Vzv��l�)I�\�)�! ����=]	p13w p�PC��m���U ������W�$�V.��YzP!-{�~Q�,��o���5������W�*李=]L�!��(��G)"{*���ج<�B	�#��- B��b�m�p!�B�
~:�sVOĊ,5D��Vh��7!�@a��9c�H����h�@Is��	u.�YjnlJV/V�u�>8q �k�A�?�� M�j�����_.C�4eHb �;Τ����H"��;����#�ҍ�!�x�����b\>|"9��ݺZZA�g�O,~(�#?9Æ�c�=�T�v�NY�bN8R5f  �AX�Io�hX�(T�b$��k��Gf���Lu�DA��?H,��	|taӆU2\3���RW5r�����@��1K���r�
Y���QqX�14�1@��9��z�(0�ŝD��4n��r�a�� vT��1`�>�:6͍�!ݾ���]�O��yRu�'"����Y<J��Lb�,[>S���	�� �̬�E�t� �[U*YfIH!b��
9^ni�� <W���1&E$��VY@�)��h 4`5�A�WbF鉵�M2d��h�>a���(1ҶU� @��bJ�!��V/5΀�j#-�
p�A�NX�(��v&�X��P�7Sv�y��$+�ƹ{�����Ac����O���M��LXp`7�S!}����3԰U��a�px.5�A�)iY��0��Z6OThHw'�~
��eX�6״�rNʵ'�0�`螵0Խ�DZ.�Ps
��p�HJ��K�� �pf�^\�(נɥ%Y��H�o�ݛ��u�p"�����B��ۼ[T��1$�� ��C0g�q�-�ĩ�W�rh'�'�>e)���X7 {I�)+6���]��iJ5K�$H�ٗdޱe�����\�S���x��DO�9f,ޓ^��qze��&��Ɛm��	4Zᜬ�7͵V����>IS͕+v7|(���?!�x�C�F<6�R�zWc��o�<IIťޓ��H���ի;�T��,ӔU^�)�a�ʖ~GJ��SNԼb�4EQ��D@�f*4|�W���^��hS�-�:��AƢ�~o찡���4`���@�d.<l�g��_��x{�̓�>��!&⟠y�h�� 4�&�ib�P�F���� �O؟�9Վ.m"�d�Y�Oą��艟R�^U��R�BM�m-ȕ��(�P�Jy�f�AJ�m�q�������� ���!̾�h�0����E��8�P%�_�x�F6@H�A��)g�敳G/qwhx;� ���B&k����enNl��"��W#R�bɗ'ޘ�%d��Q�࡫�eĦ]�0���d��C�2��눃a���[w�+�ɀ�<���	��u����	]�"����_����	��y0�� ��B�|\X`$S�t�L?�Hej��H�Y?* (�)R8Y3���󫴟��p��5j��`C��A��^{|���L&<N��rg�(lj��O�g��l�pd)F�iT5ht_� �f�Q%r�Y��P�y*�E��A��l�	*���TA���H���S�my�$ݲ3��~�� R �k� �,#6%���а ��r˹D
$d��"�H		秈��$ЌQ��pHWݘ�d��B��!s9!��:����U�"k�uz�l��#���Z�L=���0|O>q�ы�K�r���Gb�b�)�'�$0C�C���y����Ұ�E$6;�yk@%E��y2@I�
HpE2���z�PE4IY��(O��`c )�'^x�l"Sa�U�yP�� ]���I�_|�d�bd�3]rt��EK<�z���BΦ)b6O�b��g�+N��G_;��eڂ�s .@D~R�ž9����'!�SA \�ҵN؞p�U��mQ� �B�I��V�P�K	�neX5@�}@ �^M��� K#?����͐8KzTxd�G�L�h!aZ�,�!�˗4��`t��a�JI��Y�s��g�k�[��IN�'9@��M�>:�	r���"<�$��%f�zC��H����2�J8Qi���"U.C㉀BC�p���p.N���M�K|�#?	��E
w�"�?�ie`�?X��`q0oߝD�̠)��=D���b��%�����Ú?)ܠ�qa`�<I�gG���(�(��.۹hpSAݏ�&L[�"O��FRRA3�D�4��M�F"O� ���*6���Z�č!"O֐���raI3�I�J�<��g"Ote�iC,!�I#ҠY%�j9+�"OX]Ps��G�Й�'L�j�>="O���P�		QO���s�T���UCG"O�`��D����Ȇg��P��h  "O��i͈!Z]z����ΐ;�Pb"O�̈�*�*@�*��u�*<&<�#$"O8���K?]�X�2�Ȋ^#���"O ����NrP�y8���`�%	�"O�}�ď?�8���JЦ��a>D��skC"8��br��;h�n��1i=D�����%�P�8%N�e�&cp�)D� 9�'��H�-S���p��1�'D�X¤�B�`z!�r�Ǎ/wʌ�g+'D���0��n.X�*���4ʮ�Y��%D�[P����yc�ҭD	���g�!D�H�ġ_��2�ΓQ���RCn+D���GC�t�H)N1�L#�$&D�d�2	Y' Q������A|s��+D�p9QdD�b=��DT�|A�wk'D��v���?m�l�u/� � ���J#D�tP����{AmV'($:���#2D��s0	�kX��b�H(�]�0D��J�a)Έ�pc
bp2!2B3D�$a� W�^�*A
��-_/�g1D�(��IO~,Q�E��XȾY┤+D��ǈ&?��;��ȵr[�����/D��`*I����tc��Fz��b�l9D�� `���N��z1:���$p�"O�!�!e��
�z=�� �=�TP""OD�%�,@Wz��P���$��"O2����:)t婤�̨9�d�hR"OH� g�	3(*��L�4�
xCg"Or�!�-�8��re���&��es"O����P����ᵫ�kǮY
"O�yCR�ɪ	
�k�kW�O̺๡"O�C�Q��"��� X�!H<��"O �1��W2$��X2O��E��"O��� aW��`��E�7/@@��"Oa"���� �҅r3�^5���a"O,U#��ů1�^��"�À�^}��"O�I"���7t�h˖��""���s"O��J���9n扈p-�t}�R"O�����*L.�K�+K�EnP�Á"O��"QX�^S���Sg�yZ���"O,�K�t����-ȾPZ�l
"O���kݻRC�A�%FLGFգ7"O�PA���K�D�d)X�#L,��"O��H0j�Pu�ؗD�J`�"O����ϥ�Ja��E1j@H���"O�����`-
���M��G"O�S��گ|���P�[�Pae"Ot�Z��X�F&�sE�X�a���*b"O�	qBC�+լ��ԡ�9�B���"O�]XၞL;�d� _��4 �&"On�0#�0"��5�ŎN`AK'"O<��#LWe�x�rD�i���v"OI񱈄�Q�th�WC����'h���
1%�V%ST���<��
�'����������#0��	�'�"��1���/�ޔ�眪��Z�'��PP&.M^u$h��*�2O� ��'�Hb3Β34�)��Iy����'�r�!A�vF|b�f��u�����'O:P���8�NX+��ԧn�Lu��'�f��b���İ��V/]�x���'&v���ŮS�!@���^��-A�'R�){��� ��6��'H"���'u"��1�G5����ᢈ�A��=��'�N%��A�p���;ю1:|٫�'�>d�O�a�����EQ4��=p�'Զ�J��X�_'�<C�>:b(�'x��Q ��fy�!�rf�$3���'����3��a �-=pR���'����@�����JD�~��!�'�X���Y=�:S��@"f'r��'�6�Q�K�|!��a�N�k8�K
�'�\$���׬6�.����Гl	B�+�'���KE�ܥ�B
iD�oVd���'h��s�׊�j@2Lć6���'�޽Ӣ+D��qn?�����'L�D
�m�b�I��͑	yr���'t %��M?oi� Z�_2(���'�i�*�S�|eQn_*��$J
�'���I�˄ ���ړN��{�L�0	�'k��(UJ݂QV\�#�Y�{n&���'!\\���02V�\nM���S�"ON`Ȥ�&9�x[��A�p�pJ�"O�@�nծ8��{e)��Zm�!""O���ԥ���Bzf�ֿ&i`uip"O���6#J?S���K3\x,
'"O��`�C�3(�H����
[犵��"O� ��F�YC���r
��x,��"OF,��%�4HdB<�+�}�]9A"OfnΗpi���R�P�$Q��ц�<D���!�3dl�&NCB�x��(D���t�ŗXj����M'Tb��Ѭ=D�����ޘ4S>͐�.�wZHJe�&D��@���+F^E�a��&#:�2�>D��*�ƃ�\�A��@)SO4$�F@:D�<8���=!x٠�ȉl���*�'D�	�A���͓��ݚm�� A�%D�,+�l��"}q2�Y� @�T��'?D��a���)�ހ`�n�032D�
��;D� �@"�0�d���@��XF����3D� )3e\��(H���#��Т�$.D�h���Y�H���J�)�`���*D���$��((j��VJ�/8���C=D��╮d%�!T�j�<��g�1D�QF�ǚ:dT}�e+�#*�h���.D�,)����!���u�_8N�h�3D�8��F�|�U���Ð�!3�=D���1i�p�|M��CÚ�PEjP=D��{ �	���Eo� i~*���	)D�1ǎU�D�SGOy:2��� &D�,[�m��D�FU� ,^?o��Q�#&D�Pc�L��G��q�Ƅ�)[����$D��C�BƧQ?쭐�JhJ:��-#D�|`3��#R�*l�b!Á� i�&'D������VŲŅ�8L(����+D��Vo�#A�갚�LHnw�Q`��,D�d��M�$�tE`3eɳQϤx#�L-D������M:�*�#��D�VI-D�p� ,�\�� N�
	q��{��7D��$��N�x�¦��2+�
�rdf.D�����f���	�g��_x�䳢�-D��X�I*x&iY��>Lz��0�)D�����6#7���=�^�P�SE�<a�
�����i�
h���� �H�<p�ϸS^��C`.�F��G�x�<開�/f܀��s��q���,Np�<����.�J�Aā=<8�ud�p�<�E�Ӏt� A�W"G�к�!Cl�<y���_.��tIB�d�B�"�j�<��#]�*�I�/>k��1�aFf�<	1�^2" ���
L�'��P���[�<��� ���P�!�8]<Z$���OW�<	���?��d".�
�6��TKZI�<�R+ʜ_Jl�QB�ƔL�ވ���c�<�!A��nJ$bC���CÀ��RC�K�<	�(��E�����n�Z�MLE�<���O��83 Q�L���S�@C�<	ҫB�\	L;UǕ�@��@tʉ}�<���~U�����*$�QS�~�<����~��J"�"|$��|�<��gE�Fl���;By"=
���c�<Y�j�:���E��1 O~ я_�<�K�So)腈Q�c>,��1
�T�<��O�-��� �BR�M�ځ��P�<)pA��nz4�р ˅,q�:Úw�<q@	��xu)B�k�	\b<�z���U�<��з^w��'�W�v�"1�PSN�<�e�ɸ&x�2��w,.�&
H�<y�A]�P�r	�*r M2P
F�<��O�5V��k�c��/:Q�wiC�<��!�7��0p�$�7RF2���Sz�<� 4y���3@���3b��wE(��"O6��Z�l����M�*N�a�w"O�Њm�'8حȣ��!&͘c"O�$(��M�.�p�vMH:+$� ��"OX8�A��/uB��k�X4!�]Xa"O"�"�2;���c�ZT����"O���t�C"��drw.�4�����"Oܐ1���\
u*���o�f%�"Or�����g��0!a���&�\�1"O�2'�Í����Uk?[�|U8�"O��[�ř�S��}���������"O<YP&Ύ`��8� \�,�$(y3"Oڼ0L�a����ro����s�"O�l�$�V'J� �җqa��
�"O��2�/�&tN(K�P+"O0����8m�����U�t���*"OtRT�ۛ`㊱� E��!Ȧ"Ox̹"C�or�qg�&	��EB"Om#�g�%���a�%��W��<�"OP̀Q��%Zj��6�ňV�"�ن"OF�0&/Dr��]�dߙW1J�XG"O��j�H�4����#J)lQ�P"O~ك4��1d(8Q"oZ*U���b�"O`�Ʉe�en����o �)C��
G"O��щ��Noݣ��J��Z#"O�����6z,�",K*1@ �c"O���n?5le��g��t��"O�%/Ș6���%
Mb�\�{V"O�<B$�/b��|c��FꬡhS"OM���׽7�r]C�iK�_� U�3"O��8��Sz� �S�-V?:&���"O8)�g)�Ɛ+�C�U��"O��q�^�&�#'�P'dDhB"O��� Mk�ָ�gO�t��l�t"O�y��2)�z��PJ�^�R�"O�$`a�Bĩ!2+�7-2L��"OީhC�Ϥ&[H	��\�uȁ��"O1��K�Vl�"��� ����"OP�sU��,܄<�d�	�pʘA�"O���$l��[��''�e�f�P�<��� ?y�,����� H��ΉO�<�P�C}h��Y1͕ FV�c�*^n�<�g�S�jt�z�C*"�
�:�M�h�<a�W����aj�#TV`r��~�<��o��Lfpa��11.E�E)t�<����?* 1��n\P�y�4��s�<1&���.m�y4�1"bPc��E�<��.�:t�Qr�+��1��az�<!�<ab�W�V}z��O�B�<AFkֆd�z�ymÚ6-�x���@�<9U�E�)t����/D¼i �Nj�<q�W7�Dq���|;X�遆�g�<��k+b��S� ���q�o�E�<��aۅ�L���5*~}���J�<q�bIQ�p5�D��Hɺ�0r	D\�<�1��@o6L�c$��5����u�<�G��6.6Zq��ڭ(Ƣ9s��v�<Q��)=�����F<i�&�S�Y�<Q��=@9��&	av��@�P�<&��&O?Z�qI��_����Lv�<A0D=Q�Р��a��Q��U�<y��8;���a�֢7[��� ��i�<�&&�2��z�M�.��e�h�`�<��a�0n�YcL��v�
19�%�c�<� ~<3sF=�9�A�-��u�"O� @ǃ\�)9��j��K�,�.u��"O�H��ݙ7�
�A��6d����"O��apOK��FTs4�9�ji�6"Oi�0�F!B�<�#�"�2oI&D�1"O!�R�}�V��0\t��RDD�w@!�Dȩ[���"�.�&9Ir��V$�/US!򤉓&Ͱ����|�9�bD�2?x!�D\q@��G�U�F�e�� �AL!�d�>o�:5�#&��aX����P�1!�D!V�各����q�2�A�C�!򤂞D������-^��Ș1!�v�!�D�/G�n!���μ�4�i%�,V�!�3)�������d��E���r�!���jt� �??b��H��C�!�䖫J��4�GцO�B��$�Ɔ)!��)B��UH�H�9�<E��#q!�$D0W]�쓥�ϒK�JC �%S�!�\�	/�t�	O2:�X�r�ԩ$!������c�
zblR���I!�䜝3_��ѕa� {���6L�,	!��R��&4S��˗\Q�I��Z�~�!����8�<��� ܒ+QF��K�Sq!�d��ЌU���I�ԑ�ʇ%bs!�*ńe;�h�&������X!�_�v5>��.09�F(N!�DQ;!�S@ƈ���l��љy!��zG�x�L
���e��C��[!��Ƚ��:��p���M#WN!�c�>���Y�8�t([G��U8!�d\��5��A��:�2�G-S^,!�1�d enE�/�p���l!�䎻"��i�4�_6jƸ�s�φF!�d��$-�	�U��jt�UP�фs�!�q,L]Ґ!�� f28��Lv!��k�L�)F�X_� B��m !�d�\��(���`�D��H�:,�!��~���u�D.c�l22'�ji!�$گ$���$�	�`l�0�SUa!��"S�0<��Y
|�VVT� ��ćȓ'���qW	�:if 1��A�&"@ɇ�b]J0)DԲrw��Hd(րSk���ȓ1)��Ԇ�jE��p/� j���G�]21	�9)|�Kv!J�MW�U�ȓ�ܲFMB�jmk�K[
@�Z��I�(@: �P�`���*e'�
�4�ȓ���[�J��`?�Z�
OS��x�ʓ:4�� $��_���Abވe��B�	�m�ޭ�Ó�9����˳��B�&N��U�V�_�}?�=��m���DC�	���HM�qU�9�v�h(C�I?eQJ!A_�9��C&g�<[�B�^E"-hVÓhn͢Qi' 1�B�ɣ尘��[�u{�lb@���B�	90:�M�R����
SLB�I�?Y�T���M��z�ۦ�ϝF�B�	�oV��М`
*]�gAu0�C�p=��Ղ�(��7��B�C�I:��Y�b�<A�°�шNüC�I�#���U)MX����&H�lC�(�BxrS�V�^r-Sa��=KC�I'S%L� ��L����"��3H; B�	�x�����X������[��6B��"X}j��C�!�$�Tg�WpH�b$!� ��D��V�)� ��u��:
������V���&�|���9W�Oq��؃��Ϯ{���� � :=�負�νxJ����: 	��C��e@�l��|ȕ��&�j��T��0X��Ɖ�\���bb�'4���	��uC0ɋ�w#��H�H�;9H��������q�T�F���D1�Jxi�!&���R�h�X�b���g���ɱ)�"��v��V�a��(?7ƸX���%s��c0CŪM��6�X�K��T��CN�xd�P�����E�ԍ
�t[Z5.x���O���=�V%:�M/y��lڸpZ�s���?�ħqG�(f��1:����eE7z  g��`�^�c/I�]^Tp�'Bb>�Ji�`����`ƌc~|h��Q(���	։�Nd�0�� i��)�j]�t�į�P0]
ŀ]p`ţ���L�H�5!�� �R��OXX {�˄	c�nD���G���3��E�8q̟h~�I�Z9|ga�T-N�v$]��G�.F����$��0b�a��!y~��r@�}b�J
�'�J�;��I�!⎸ ��� @�xL�p��?3���l��бmڴRQ>��T�QU�]?o�ua@�vSf��jE��x2�87茬����� y�D0�y�I
\��,	��&B�г����y���%a�(ЊF�J1}/�x����y2ꀇ1/�pHP��8v�04���y2�N*W�T1��6|�
�1"#��y���HaR��]8)�"��[?�y��Y�"_���P��%V4�: G���y��:b�$p�D�B�+���gI���y����q!(1�D�TC��
���y" u�h�va�B�8��k��y̜5!�Q���P�=pN89�D��y�"[���ud��:��Ph�6�y��� �݃b��/Z�V�+�y�H���b���k��s�ta3�c֎�y�,�9�@Z�ĊekP$��Ȏ3�y��)k�&蘳��
g_�xB�ύ�y2e�8A�� i,\�l��d�y2�6~�� �I��A�!&�y2Ēk�hx� k����"��y�c�+�u���F�$�SE�.�y�e/��\�v��<b򘐊����yʖk�$�cD��Y�T�ˢ ���y��_c�a`�!�m*�/��y"�A�6y��;���|%>\��I��y�dȂ(��pj�1�i9�@��y�KT	]P��*�EC"�N�b�LA�y��F�!��	
mzA�Dl�
�y�l�&�s�FV5��c��y�e��V�("��ؔO�luW�O)�y2�
2o�Y`�GA^h�3��ʏ�y��q}�����=
�D1{�X,�y§׉M��z�㌰}���3Q�Ę�y�%a>0r�薬n��Ab��W�y�&��1)
5���\=����֞�y��*mĸ�r7�� c��)a'�M�yRF��*��h���9/˂PS�J��yb��M�~�t��,��(��Z��y�OD;_�\PR'���!N>�%F�(�yB,;E�]��d/��!$���y�$L��P��ܟ9�Љ����6�y��X0(����� +D�zu�ǀ�y�?��I�7A�;5���Ͼ�yR�8X0IT+D ����5D��y�D-NlD�����w�(h�rk���yC�*D�lx'�v	ni0BLW.�y��֐}�P��`�n�<<�r�Ǘ�yraї1��� 
͕g�nu����y`T�z���6c�_DΘ��	�yb"�{ <[%&G!l��,������y�#�ht�5�R� �5����A�y
� ��B���	1�p�Rj��3`"O2��խS�G����)�@�A`"O�hF��8tY�c^�|<��q"O�1�g�·w��!�o���p}�"O��s�j� ���g��C�ЁYP"O�D�1��CF��`TI����3"O��p��`T)�!J
��E�0"O���n�	�t�1 �*,�ʕ�"O�T!U$��n+nt��a2�0y@�"Ov����2
����� �y����"Oԭc���-���C��R���Ib1"O*��̊,�A���[�<@�"O&�B�����TPc����j���"O�t���%�*�����y��{"O^ ���� ���Sˌ�J2����"O���2ږ$�u����8b0���G"O�hΒ�wN�Y�iSa3t!���G�O���됅@!X�uk�R1;����'��4�U�!}D����*1�\A��'9r��g	�4��dSsj�&����'��XRI�=i�q�Ǥ��!2T�	�'��Qp�띦$�4*���_Bf�ȓb׬T�c�Ӗ ��QJE�V�	��m�ȓs��DR6��"���#�^-	2]�ȓe��� �A�2��	A6�ލ5����ȓZA�l!���[��HT܃CBE�ȓ{����vF��{!���&ūa�8��E��sg*ȭ+���8�O#u�Z����Q��b��c��x ��ML�E�ȓm���
D"��ô�C�l��O�P��ȓ_M���E��. 8=����mb�i�ȓ)ذ̖ٔ+�T�Bl(fv-��"�|��P�hĸڴ�(Wڄ��y�4b"*͉RS���g��a?���ȓ ��!e�@�{+2�0�q�d"�'4�(�Lƴpc�pbB�;:Z<��'=v���%��b:��˽+��0��'�`܀g-�)*eIǡ�s��=��'���b�� 1�8d3�B �p����'�Ċ��G)r�JXa�e�a�< �'��X�4,ާ6���I���;P�'����:E�h"1Ό�}^�͊�'SP5p�H�W�<�!�i$JƦ���'�f݃T��9%��l# �::iBh�'�l��u�Ou!�����2
����'��Ń�
��b���<��+D� ��=�`TR�֤3
����(D���j�'z����юob����B2D�T9wb^�;��YS����<9rW)&D����b�>=-�Xx`�U*3g޹���$D� ��#ԉi��5���k�r����"D�����0��QsRʌӲ��E�!D�hJ1���@"�S5�����9D�t�Ɔ��P����Ȯs/^�bE�5D�$�HF�9a�#��IR�Z�%N!D�����1��r興U�2��`!D��
!��zj�	cG��a��=;%�1D�8�4�P�^g\���6-Б���1D��&)�>hH�B��C�z갽�P-.D����9Y}���PQ:�cM+D�`����;�L��eM�:��ٸ�'D�h��LY,+!��F"�<S/dH�$0D���
��-�`��aE�	�N|��"0D�Q@�O�XU�D9���<d�6��"i9D�� �y��͈(}4�I���m,��S�"O�`����`�G���d�` �"Ol�Ư�s�dC�߆:���`"Op�:��
#�~A�J�p�51�"OP���7H ��>m�� "O�L�'(�-�\����?@��}x"O���*�r٫�l� 	�Ij�"O�a1��e4���Ź_}Jd"O�wKhҝ1E
ȝT(�1�"O�i"�Y�1�m"��H�*&�d #"O��y�hմB�x�s5�ܦ\ ��S"O�P@��JH����N	8�( P"O����ГSvP�@�S.G&y�&"O�0y�J�r~�As&Ͼ�j�"O>�f��^�2<ZQ�:���f"OXQY1
�DV�}��F���{&"O<�8!�^t����*��:q���"O���U$�~X�s�˟Z_0șq"O�D�b̆4it�`Y놕+r��u"OM���1ۦ8@iQ\ppb�"O.���R����HXx!�y⁃�+�5)M�@徼!g�@4�y���8ye>��Iҿ2�2Q)�e֏�y�h*� �FU�n��b����yB�B�'�x6&V�q0<5 ��P�LS!�d\��<+r&ߛr�B��<!�Ā=,�]�R ��\�ZM����l�!�$�&�(�*RCz�fSvmWW�!��fq�k��w�.hWm��a�!򄍝i*�� '$��A��ǂ�!򄟎#���zU�5V�����,�
�!��P9BlX�"`�E56Y4�����IZ!�F'T+��B�g߶E�v,c'd�>pW!�Dԩ_�<Y�#_,m�����]	U!���(Q�P���Η�^��ѩ�Y�e !�D��o�8-��lK��"������:!��-#-�T�c-�r����D`��!���X(�dp�e܉e��Y�/� �!�䘈~u��9���tE H��囔G\!��0�>�iŌ0,T4�#
/_!����L��jG2:�����X!�$׽K��P�:\��8��� @!�$��Eɦ��v희O�P�%�;	2!�DO�sah�T�3�8M	VK�6	!��4h���2f�
Rm:e�"��',
!��k|R����I>_��I�nN!�!5�w��0V2�aa�-M�@_!�܆{�B)�#��N���L� o@!�͑9�t��a�,D#th F�F��!�$�(j %!q%�(}�L��$Z'p$!�D��Ej�0���	<Rʰ��b_�n�!�dɶ��Ae�"p U�WB	gF!�D:}w�0:eHH)v{4CN�TB!�ڟ)����c^4���[�s1!�dD��N��i_�<���(�!�D"VU��j��қa�Ջ�\�z/!�d�y��˂���4Q�l	���
!���F���JT�	B7@��.��`!��	AP��K�ؠ�DLǊeW!�$֦%�20
4�/@Of)�w`��)�!�$��j�)��DvD�ɌTt!�D�z��	f�y�0XS$�[�z_!���4>b`�a�ߦD��P�H9kS!򄋔G�d-��Ĩ�~=#�g� @!�� $K���)��UC��Zzn�+D"O���1��=p�z���e�,q�x�E"O ����5.Bdz%�rkP�"O5cf�T���KA��=� 0�"O�/�3q��IQ�ϐs>�l3�"O���-�K
�C��ќC�0!"O���wjB�{�4b�,5��i��"O*�Q�*f������C%�u"OZ481	��[|��c��$�,!Q"O(@��#AOP0�˪j:!�C Z�x���@����G]�/Y!���k.���+H��h�	��N'!�$�.���r�X�Q�RE)t��3/8!�Dع.�:��N�d����U--!�^`�����y�������Pu�C�I�nC��I�*\��Գ���p5B䉵aܹp�H��T
��q � s��C�I+f�r<�� 'a{zD���?$afC�9_�:�7�E&}�^�b�Ǜ0	.C䉣KT"��)���kԉ�7.x�B�81utl�Ec� ��yw�H��B䉬	��Ȑ�뜑*�Q�w5��B�7&��U�և��V���X O޵]}�B�I�;Wh�"ꑡ1kl���6�6C�I'�88sCܟ_�98�ξe�C��ʠ�F��1>RY���
'b,DB�	2�`Ԉ�h�sC��1A�	';B�I��-)V"�]M
'K3C�+o�����)�Q������0B�I-),~ @   �T   �  �  �"  �-  F8  zC  �L  �R  /Y  �_   g  'o  ~u  �{  �  J�  ��  �  �  ʠ   `� u�	����Zv)C�'ll\�0�Kz+�D�����b�f޵�y2�S��y"��g+R���/�V����C�	^��dl�CMNA�4�۴hy��sE��{���\���:J�	��o�59��>a��D�" J cVʴi�%U2]+b��&O�B���7�>�x��I��i��'�?�&IV�*!��B3� ��V�ΙB�
d��M�
,�%N%aңF�~_�6m�?���D�O����O����� �\�"���,ݎ ��L+��d�O��nZ{!f��'4�j�9hz��'�⁐�O�"T{+�GavJf�W:"���'�b�'.r�'����1�u���\�ld/��~Vx�BS�=.i� ��Fl�GE�<��S�<Hq�\�Op�q�%ˋ��e����
���#4)�:<�~꓌y2�����q
G�����I�=��j�� +<b��삑���$��)�	������<��ޟT�O$���9�i�P���0|_BTxr�'��7-Ʀ)�شog�&�'��7-�7!�Zml�	��\�ǺQ� 3��H�K�����H�)�@�R3��AP��Yd���WCEJF�E�X�Ժ�a�;���H��E^!�đd��� `���K$=D���H��M�s�i��6����'L�Ԙ�5��B���0<���f/Ԋl0}m�?]�q֢0^��S��/����66��aC�iaV6צ��ՈS.:��]X�jĶK�B@2@��?YW"���#ew\��4,�fv��r��2'.\�ā��r)�b�օs#��5G���Ғ�U�U��i�i��3R�T;��즕Y�4}x��k\�/����M,29c&C*L�2в�T�4Y���*�FI#�cӚ�RA&�<�@T;��¨.i�e`te�O��|)�O�G��!��U(W���D�^�r�DX�����ӟ����?i��[?S������h���@-<,���N7L�H�韜��+2�D������c_�8�#aF-$s��xޱ�6�<����\?,��q�3O�`h&�@�j�Hg.K�O���2��
�ew�i�ѭ/�r�b�ޤv4H�RU���XT�c�{
[,�?a��i�V˓$M.=8VH-%(x��#�|��p�I�� ��x�	ݟ��I������|zPM�:b�MW��3#2 4q CZ����IC��u/Ck����Ή�"y�y��{�>�d����J�M����$������OVT#f�j=���rl�
e+�\��K�O��J��k�T#�h;���;wϛF�	�}Ih�`vKZ�P�����C	�J����0�xF�
�)�ȅr�hG!���2��Ʉ�W�HX��D+>�X)ԣ���	W*d�����=���Iu>���B�=I
���.���V(�Հ�O���F�����,�z�`���;ư�GA��P�ўD��M3t�i2b�k�,�ɨ�x䀂	��`����% �$�O��}uv����?���?Y/Oz��!LO,PL�x�*|>V��1j
&�>tUbG�a�	
�3X��OU���C��8e���s�@/"�Fdx6�  �e*�n� �� b�HP�c>�kI<��iW�*0(:D��D�)I�I�7�M�^��8���Ol��7&����n�1�I�V���%���TƒΟt�	`y2�'(��f ,�Б�
(*��R�o׾dDdy��ʟ|yڴ5\�V�|�O���V�����O�#%x����!LW<#s,�۲eD�0����O4���O�<���?���?� ˆ�I �� `�f�hu��{2���ǂ>Q��I��Q�a��y2�Ң*M~ãfҹ"I��@�	�S�|)[�Ŋ(J�)�Q"�T�����N٪B)ў��"j�Z�x	r �,.�P�"ӗA$"���Ц����$<��7�	BSH��%3X|9`e�1��M��h����%?e�<!ƍ	EA����̍�X�B�ݟ�S�4�?�A�i6�7M�|���[�6�'Hb��3��]�T2��}�Pb�R�'�|P���'(��'�J��K
�9�R����ה/4�N5S��4����I���KFA�Cax҂�6)���$�(<zH��\Ǵ�ht���$��Ŗ"6�N�B"f �q�Q�d����O�,n��M��N�쀖 ��L�@��UBǢ��]�/Oz���O4��5� *eB�"Ig�X���/�6i����Oң}j׺i���`�N�:�r���v��u�p�^���Ŧ�r��8�M��������i�OLl�S �*��t��*G.)K�#E��Op��L�:۸,���P�`8�6�͕�M3���C�19��J �{a2�TG��8S��D��C0$��+��)Uf2���-Knh-k��ܿ ���S&h\(��c�m� s� �d�$9)�O�C��'��7��I�Sw�']��u
�O�	]^��D�@!:�P�$�4��m������dy�ߠn8� i\$o����I�#=���B�i�"z�.���-h�"�BBa�9E&6M2b�	N�nZƟp�	�`j�nK�,�u�Iɟ��	��ϻ'tx!�M5j�YB�흍C���FÄB P�ڴKn\�rj����O��^�^�Yv�
�K�<@��Bu�eIV쑄V�D��g�9VP��$gԜ=�-�Ɛ�C�A	B8�n�.���V�Y'H��T��#�`�7��/����5�B��'���'��� �$�g�̵�u�G��hK�'@��'��'���U��x0D��}��5)e[�)r�\�	ƟX	ߴB�F�'7 7��O���n�'�|i�`N�HQ��=�D\X�Ɓ�pZ`����?����?	��l���O��S�6\4��jާ���Ǽ<��X/��ɀ�S��ވ��"J%��<��G�<=lh�GO	y��9f�I\^Ax�N�.&������P���З�� Q,��eF���#R,�k�$
)5��A5���.������� �	ǟ|�?I���M,9f9��$�pP�MZ��{�$L�lW����>M6� C����'�R7��O ˓N
ġ���i?r�'hl���H�'c_�iq����a;>�9�'�2��A��' �<U�Ji�
�-GP�X8�6�� :b�زj�L�JG�.r��1�=��C�r�3��9w�,ə#� W�B��u�^n�่V"��9t�Dp2�<g�.�x�l�XW�➠Z6��O4�%���9'�ZP ��Ռ6pZ��;D���UM�M�������&O R!�,�O6=�I�E2!�`��EoB�blS(��Of�Ӳ�Ѧ!�	���O'b�x��'�<�p�I�#�d�!UW�u��A���'�b�� dpmXn<-m�Uq�m�>ـ���IJ;G��{�N.Di��"q�<;���k���&��O���t��0D�ȕ���ue�A�iI=D,t6��e2y�����o��	&d���_�)§IN`{���1�@�El�<r���>Ζ�A��]�4ѫSCZQ���G"�6ڧ .����8�fm�03��ش�����P�����`�'$��а��|���p灍��}A5m��?���$�d�>��R����'^A�O��s6Ӛ/��uc����(*��P�7]��-�q�Ҫt��<#�1�:�O��#�����qR���#KjXq�b}�r��'X1���˟�'i�5[(ŘWu��S���9R�Aٶ�'��W�p�Ie�g���l�����.$Vx���~b�'d6��ۦ�&���?ɔ'������^�Ij0�F�'b�����M�öI���'nB�'or����؟����"K�b�,$��"Q^}諲�L�]������yD�%�ϓ-4jI�D��$8ʀ��b��!=�c�T�a��L�s��#5Py0сߡͬE��-�,�hI�I>��-��"6m�Ve�3l0���9/���ɬ�M+��	O�W��	��E�A�>D×�Ta�h���']���A�d ��$��W��X�K>a$�i~�7M�<�Ei�2@S���'K"��%<���+�jS�P`�P�-^�= ��'��=c��'�6�"|��)�(F�!�Ҕ	d�oZ'ф�Y䃙4/o�H�#e8���D:&�|�x����@�ґb�c�ͦ}Y�A�؀�fJϺ�),џ\����On�$6?AT�R\ʲ@�{�(�bg��T�I͟���I�O���B'����0�㗌T�n��F{�O������	�6l���8^�xT+񊆩oZ��K�K��M�H~j,�"��6@�ΰ�`ԧ)��Dc�f��tk����Od5���B4aLȄI�b�-v��$�eF[<�
�&�?�#�A'c���3$�RRn>����6}�V90���䅑�4��gΑ�N�v7m��k��Z����C$z&�dSe%�zwJ�{*x~�J��?I��i��"}ʟOK����c��U�2�[^�����<	��?�̟\Y��P[3@��f#�'^��*q��󟌓ܴy4�&�'�6y>����v8�y��EM��l	���I՟��	��rT��t����ӟ��I�k�H�(�h4���čn$�i��/�Zx�?
�4�[�E�y�p��Y>1��NI�'�U� �4f(s�dR����j�ឈ:xz)a@Ᏺ4�X�%��(n�ʧ���,�&�yW��0j��Eբ&`�3v��".��/�<q0������^�L>	C͝�;8ʀH����pL�薅'�hO����՟&�傑hA1v��b@h�R�'v<6�Uئ�$����?�'�|01 �� �-�֠�=1uZģ��%�db �'5r�',b�b�1�	ΟX�I�kJē���,o�6P��A�0)q CnL<�Y�E�'`����L�"gV���5�E;WN	d$�#}��}��Z�h��P�P�K�P5*�C��;w>Di�=a珝8*Pa��+H�,GF(V�X*Y��8�	8��9����"<�%�ҹ]b�����DC�Bu���V�<��3es"�;#H[3�f�
�A�W򉌟M[�i��	�V����ٴ�?���/>��5".1�� +�3b�a��?��=�?q���D�5�?ɈyҌ���ڬ��_[|�4x@���0<a&��f�']���R�X�B�N��5go�ju��i���I��6~zl�'IՓim��(]4NLVɇȓ:�lD�'$K%�@LTYǔ��	�?�c� �B�!)8l�-"_ޜ$��H����M3��?)+���!f�O�}��$>G����7$0N6�����O"��O1���g�T�X�����&�%~�|��j��aAΟ�DQ`�O�7���@� k���R���Z�f�<6��A �@�*,H8�広f�.X`�8�O4^ɘ����Da>d  �P���J�O����'��>q�	�Dc�Ub��B�&R5��o�>g��T�ȓ2�<��K:y�4����s>�F{�'0|#=y�BG�+nec3K��9���Z�_�K/���'O"�'�<��A,[��'��'�󮘧�ʍ�_* ��ܩ�8�F�Z,ѳNq:!cJK�]v�0�`]>��S2�'d���)&X��Ba՟�`�4A��`�:���e��(JEp"��6H%��^>�4c-|��;Y:���MM#]QHh@F���~�t��4c��I�3}������g�
 f}"�bJ	5��ѱ�@�bL,�F{��'�|�h��&]}^��i��m�,1[���?)��i7-:�4��I�<���- �J�FM��/[��T�M�J]��HI2�?A��?Q�����O����O6b�o�.@�>y9&C�+���y�J�1���r��s��)�.�zD��иˀ N�GJ����H�#o��A3�%�`��p���A �(��p��P�?�P�D(@���'.IB4GP62e�B���(a�aRRbՄ�?ad�iB"=A���G183
���Y
^�y�𩌥3orO@���ɔZ���壟�6lI�`�|}�~�nzy�'� S����?�6@̿M �` cB�1I�LG��?Y��a��Q��?�M^�̸5�P�uJ���JG�fL���53�<t*2k֣e=�@z!lD s�0"?����m�P��p�XG�$T�Z�����م;�i6jP�!~,�8�i l��A�Ѝ��'n�r��x��6�x�d����nEX��ǿJ�D��s⌒'@�˓�?���?y�'f�.����&����Je�5�<�ܴ�O�S��M�H�woƩkukJ�(Jp�'*���X�x��T	��$�O�˧s�M��|�l�%�O�\���X�4�����?q�%HKK&	�bDD/�l��U�i�M���n��i2���=�x|�U�c"�IKWeiQ�M#g��p��m[/t"����`O��d���ˆ9P�zH�OJk~2K��?a�i��6�Ol"|J��K�.v\�am�9�&�`����@�'z"�'��ϸ'�ժvjJ������ˊjh��ʋ���O�amZ��MkL>Y�bY�2	6PK���@�&̚����'m�!��?	�eL�q�e�?����?���/-뮌�>���%'�_��	&R���/�*d8������J�݃"�%����y`�B&��9g>T)��T���(Q�E�2Q�4�``_�q�����OubO��p��0'��R%�+Vcx���'S��+V�����Or�=Y�mô Ԍl�w��%������y��Վ or�`��V8�$�1-Ě��d�L�����'���~	�G(	+��hd�
W����	5꘹��ǟ8�IΟp�_w"2�'/�(k�ҌdR-2�I����Y��h��!	�sv��q��I�����C
G* ��2)�K�aY�<���צ�MP������1 tX��$FMR����=8��X�(Rg��yrW���I<)���?H>��?�t1ZU�Q�.h`pps�$0K��J���?��ٸ�?����?��(��.i��,�d�k�|��S"$H���� �<��?���iEY����έ����O�M` O�Oq-q�']"Zgz�1�*�OT�$�v����O��Ӌx`�{b��;J!�xP���1�t}��L[���ٲ$��4�>d3��)O�d�U�C�5>h$駦��e��KT&�-#Xbd�G�{�ՂP`]LaxbC��,��d~����61A�Ţ�# jK����0>�(A�V7��c�
8^��d�1��e���y�H��#���0<E*��YF2I��hy�gK]9�7m�O���|*��M!�?�� ���@H#�	g�����ߚ�?���aLM9B9hɾ�0W���D�yC�]�"��͟��9���o� �C+_0v�nA��x8����W��E	ㄜ�'P�@�'�
s�Ar%�~:C艷G�=���ͧ`�(�9��I^~R���?qQ�i!�"}R�OI*}�Q��w
q�$ �02(���'�D�"�7��1�&J*~�<�����OxxGz2l�o�����!�'�n`IT �n��6-�O��tSt���'�?i��?�/OR�9���W�@�8e$Y(z@�1q�_�c����K�f3~����"c>e�� I$���5��z��	�r���e�'�0`����� Y1�A*E@j�
`�	��0ʧ4�����ݼ�� S�.�J�
�zd��p�����M�U��;��O��I9&�dۦ.�8����-ಎҪI!��ECډ��!Շ�RP*5-��/�'�"=ͧ�?	,O���i��Xe;���[�ꨠ��Δ!��E.<Z���O����O���;�?1����D���.}�bo�Ix���4�T5&���pP��6�1G�ӷkƈ�*qH�?7.��Gy�Ф(�ҩK6�3�(��g��<���K)S�R��	��\�)��,A�^�)3U���	��'�)E�B�#)��8�?Ѫ��	��?y��'4���r��I�g*�2v��qߓ��'�`qAFI�8�P����mvMQN>9�i��'ڴ����sӠ�d�On`�C�ֱ:��hb��''�iF
�ON��F��(��O`� ŤaҨB
� �����z%�e����1��2E;��V�!O����L�>�2��r�i��@�	>d��@ aA�+.����ٴ(������r�6�D�/5)b�+bjK�1������R�!�ڸt=���М��a�Ֆu �O��=ͧ+R�����D\�8f���&�]�� 	��1��i@��'r��x�Ɏ	�tH�t�\<D�j�`*J�A�\]�����{�/���l*��߈0��Tr���s�j����}�$�]�i�����_�L�y@.ڔ08�	.9���cbѭ92�pb�'x�@����Xn�������:T(ŇX,|�EAņk��łb���FK�O��'�"|�nֺE�b���)C�T��pB�O�<��ıb�nd���R "�KcK�'8t�}ҷ��Vn85��$HF졑P��MS��?����0aq⨜��?A��?I��y'���%�#�;@����_�+��qY�hQKT`��@U�?�"É���9��^**�2q-��OBp�F�ֺ|\ e��6�X���"�W`���5�P�X�ʧۛv�P��y� ��02l x$�S8$�=�b�-��S9$����DΦ)���5?'�`e�߾31!�D�b��p!�1T�g�ֈ&�2�'�#=�'��Y�8-t��su\A���<%��%r�u0��?!��?�d����D�O擥P��}��ǬF׺�I��t
u�A@�g�Tk5Hƀ3�JM��']\�'BѡQO��R+�#�J�6��5 C*�A��%E�R��H=�nQ� �R�Tϔ.eM�c����Y�|�D�ҫ)g�X@T�D&��D�w�����($D�C��p��a�ŧ D�P���6[�j�kPm�쬀��=�����%��1D]!����OV��֯W� q�A��lO�<�uD�OZ��ڶ
����O��S�*�z��ӣ�|	��v�#\�z���״3L�;E	�T�� vn5O!�!nP2Z/D$�t�
�c�� �ؕnWHĢ�	�,s�8Ũp�J�m�ax2B��T�ID~�����f��-��t��%O����0>1�Lߴ1aR��q=zZ8R���Z��P���u7 �q��q���CBWy%���	Dy� ��Jjb�'{"W>굄���@���#.ش�6�^�L���e!ߟ<�I�F�q����o6�d���T�.0P��ޟ��'Y��Qb�O�~Qj��a��R,��'�|��!�
,Q�x�2mR,}����2�G	>�ʟ����8�j�B�g��=̴:���Ⱥ���OZ�$'�'�y�F�14:8q�5(Z� �PQ�A�[��y���A�2��I�F�d@�����G�O�T�c��ڸ&���R�7(��Ժif��'�� <�iw�'_��'18�v�RNڹ2�ΰ�EZ.�@1���E�I%kfF���-�3�ɿ*m�	���=.��K1��X �܂��(L�^A��$N3��%�����'_F~��-�м{�+�	l �8���&}���c�K,��~���IN�g̓_�@	�p�*C몰�Q���v���3*�1JR�ll�2�,
�\���'>L"=�'��fl�R�
�5 &5:%*�9���spoHV�r����?���?�'�?�����t�E�+v�;%iƱ~��b�*\+)$<�4��0d�&<��m�3Q��)����}DўP�q+�PeD��Ы�7*R��D��.MC0az&��
.�eñ�Os:<���޿gE�x�Q�o�	>fE�8�7������cb�;Y�%2���OL��.ړ�O����K ~�J8�t�?�e2p"O����q
����dөC�h�"�|�l���D�<�l��Yd�Sꟴ�פS&~͐X���=����ş$���O�V�������'V�xl��mѶ4>�����S�IM���Я��0U��`�.M?a�sc;�ʉ���>���Tf5~���`e�����Y�t����@H+ai�,���MK h��e�OA2��'�����tרG�N��#f��U�r����&��2�O�I�-�
_���#���Y�q�'�l�dÁ"��y�f2#J��S䤌�O�Z�D ����Ms��?�*�d5���OL)q�ǚc`��q�Z)A�x����Ol���,c~)c�J��$��e�	T�ʧ����+�����8Ŷɹ���m��	�}X��p��%	���#JK�Q>��Ӄ6_���ڃ�H5U�T�!7	5?A��Ox��'ڧ�y�mޗ���8gҥL��T	���y.P�_���5���x��s�b����O��G�T`�2�:�Y�o�o(���넽�?����?���.�TKD�˱�?Y��?����y�M�)R{����6|���!�=s���+V��nA(0dX�0��J��ĢU�
u~\�?���eK  ��ǀ��~`���H=<��	@Q8oc���QH~jݴqL @z�w��Dkt�L�z{�ZcȂ�E�0�����$P���'�ў4R"NV�S��9�"L�Ҙj�'E�<�`��?��M@�Rے��agBCy��&��|J���$��/�{Ꞣ5���;G �!d�8e�Oh���$�O����O� ���?�����T�
֘�)��U9�� 9�
�. ��P��J�eW�����ֈ*eM�W�'���p଀,l��l��ď���Q`)\�~��h�%_&>���Hހ7囖��I���${#IV9Fh���2O��5�ޚ<[��Ĕ~��\�Ů�'H0�{uEI)���Y m2D�8��O�FLq�Ѕ��9f�XaKL>�b�i��'b��c2�.�	�''�@p�>M��h�lʦwbS�\�	����	RD�xSaI�

��q�P��?!��R�9��c��?j�|�b�� _��hS+ш(�"ɚg�Z(n$�B�O4���/�&W��y��E5�H	�K��HO�d��'�r���9N�7}4�,�9���'���O���͹ic��G�=!T(�$��-��O��=�''�2,M'��T��IW�P����K��?�)O��A�<�O�S蟜 f�c��Y��JQH���U���ɚ=�@phfb�7O�A�@��?E��2#<��,/���ԋ�>��$c7�	��n�Y� �b��x���	�S⓮_-��i��P�y�pQ�O�����a�	ڟ�E��4O� �1�vԔO�i�Bꓩ6��xY�"O�A���ԙ:=�sv��[�>��E�	ǟ���aP"��A���eH��ѯD�	�����D�	p���$�Oj���O�˓H�������x��MC	Y( ^�RS�L9
2T���'�NU��$H���Ϙ'͜�DFB8Y���"*���4�����r� ⶉ����4�I"��O�,� "��>I�K�'
�n�*�]��4�W�����'� �i��?���S�R�8"�fݓ���R��Ir����#f �o@'I���� G��F�����?iC�)(OL-A���:FA��,��O���/^���d�Op���O(�S�'�	�U�TF
����"z)~Q���^:�U�曛zA����'jN�Q����C �G}� �d�
.5��Yl�H���.�w�̜� S�?D&"=��d�4=+w���:qnhT��C��q�I���F{�I�&�(�A��,堅�� �$H��;�IYaX���"B��S����=<�OZ,�'��	�hPF�XH~ڲG�9�a��C�$n�q�%�ş��'"�'wk1�"M�	�?^�����Oz�zd��g����JB!z�Q���'-�풃��ctJ	�׎ZL����ؾ%wN S����!Z��Q#��qiX!�!)ғJ�)�Iܟ`�'�6���F=�r�D�)�B�N>i
�f ��P�$`�X��DL���?!��4����	.�\`W���?C��Q��ۮUp:�D�<�'��?�O� B?U����s�Ƥ:�<4;RL�0b b�'���@*Ψ3��cTN�a�:��=nip9(�(�RE��K�J���2�b�B�R�4�]���4%�����O�Od`���.��(rK�Ȋ�5��8��O^���'Y���<�c�4"\��##o�SU��2B�i�<�
��_ �h��+CT�Z��n�'�Ҍ<�s�<�D����x���>�
 ,O"�Q�0���?���?�-O(Y�3+�CM��e���8��,p��ґ��#u�Q�t�Pc>c�dB �'PĲh�QON�F�
��Ů�?H��c��F�.�[D�'�c>uw�� ����/�mX�	W�ݸ�đ$|]ғ�ԣqg�O���!ړА���"?��	"�U�(a�Lq
�'�:��K��}�����`U=5|@�
��?!��)�+O&`Z��\7�p�@�;�-1��I""&؅��jӖ�Sg�;Bw�y��J�vBX�ɿs<(`�D�Y�ߵ����8aц=�Ŏ۽9m���'ϟ8���������П�0ff�)\�ܵ�ƌ�'	Դ�����yg,�"6�ʶ_[D�8e���*J������V�p�<�7��,h5I	f�=&P��!�#dⲼ�d�w��\ۃ�ND<Ȓ�ӣ'��<a@�
柔��Ģ=��1EI�$Ā9(��M�6�pI�'"a~"���+^��k�N� #�q�I�:��>�`V�iD��b5f��w�ɏ+R���@ȭ<�&���?y��?�.�Ĩ��E�O���Q�$t|�+�t��fF�s0r�DeMI 1*�깸�FQ�+⒜᢯E*r(ډ�4"�ńj�c�dZ�2���0�yR�E<2U���"���Qjҩ2C$�9�X��3��o�'{ƐʧeVsFX�H�n��U�N �Yfu��Ɵt��'���F������+����`�0mS!򤑯�:�B��JC�rY�u�R8r�ў����)���X}���!X�8�wN� n���O��d��M�Y�3&�Or���O��D������P}��c�R4au��*�ނ�Z�aF�'1Ƒ&[,B�4���)
�*@+l���'��U���&�
0׆J
E�Q{���L�<�Cs���}k��)W/'��I�9��HH��0��ā1�j����(�>y���$?�7��۟���E�'��
'��|aG�9[*=�gĠx!��t9�	�@_C�xD�Y�9 b�$��|J����D�;5�v�� �z,1�����%���-V�T���'�"�'p�g�%����̧����މqd���q-�(���9�ޑX<0+D���(��n��&�����f�:��ēӦ��<�R��eɾU  *���%)+�I��+��9=DTb��䑩d5�F��1�$AQ#ƪ!�
�B�٤b�	M�'��Ac��޸8�Dze�P�mX�'
�)¢��\��$��.ȇZ]��0/O�Hlϟ��'�z��"Q?=���<�lB�y��ї���u���t*7�Aߟ�IϟPsR�=E�XL�����(w���FT/8�&�s�@&M� �1d�����H�.�SQԢ<����z�L��2�ڿ-���aרV�d6Դ��&W�JH�ǮO�Us�uh3���x �ո����{�Y��퟼�|�V>>M��&�W1P�8= ��Tqy��'��� ��>�J�2��I��	�N>q��4��U�'Lv�U ͂l	�(�T��-�q�.O�����O����O�˧iS��X��?ᶣ�=:V�Ă"�<����(�?!c�E�|On0� 掏b�"b�ۦ8H�^̧��M��F�GS:�у��Y�8�� �ף�hF����()�8���������$"��'qnڱ�Q�Q�bs�~k��>Olzd�'�ҟ�����S�? 4d�&4|q�Y;�&,_̽�1"O�K$n�*,�'&(Uj�e��O��Ez�O������
@bXZ�R6bc����'��'N2�yvC�:��'r��'s���'1dP��')OI��0WȘ�QrY�"��N5h�I�R���-������'GZ5�7��&3��3p�t�2 ��"X+Z&��{�̀�7�\e3e��L4�S��MCe���b9k1��˄�?I�洠�A��	�N$�!���qAg�O���6��y��YD�P�H�h
�4�[����x��k�F����(Ov\�`��1x�;��|�����$��u�7�Fe9�g�|� ��-i*d���O6���O$���?��������}���B���>7�� ��_0A�p\�D�68�A��+J,Ѣ�Ȋ=+'5EyrG\�}�Q9��P�I�)h�����7�>}L
�:5�\F*��q��[�K�D�$�%K"H��W� #LP��+'��uX�iC D�moZ�HO�">A��\	��wN�+E|nX �@�t�<��$�2��\�r%\�!x0UWy�bt���D�<i�����'0�1�^1r�(�7��X����4iPx;��'o��#�'d��'L�;0�[�H��@	# g�6�i>9y�#������E�%p���bP�#�*�t����z�x\�nZ���	�Z�0��+s��;��޾C��qQk�O��n���'��(Q@$�7C�R�����>;��I��?	M>����?�,O��d�Op c%�!`r1T�� O���7H�O���/�<Z֒OX�)G�瓟���ջ¾�K��  k`�_�DxFa�<!���?���?Y��?����?)�Or|p
�A?I��A(2ČcJH4@����E�O��<�DmN���&��[lL���"�M)�ē=��Ķ~R�ɘ�-
(1Q��7t��䡥J`����')j��>OF���'9��O�;O�2H���.�ˣ�ɣ6oX���L,6-�O�4i��Oh片J$V�s��DK�\cԼ)QN�0]V��#�Gd��uk�����I;Fܔ͓�u��'���Oj�=O���4�!'[
�3R�ΰp��`���[9I,��'��g�'�����&����u��A�<9+II� �B�.˚L(�FF��?��n��D�	�"i|��������Ov���OrH���Y�.D`w/^�}���ȅ��U�:�F�'E�� �'����B�{��i/���U�ݫ�rL��/�0bT�U��,�26�|�,3 ��O$�^�Rc���	����?���v9 ��EL�yN0��"
���0�#��)�y2���?��,��.�O��ɋ.��u�S�Y�2,[!On�����;QZ�`��5>ϰ-���<����۟��	!Mc��'�?���Q����⑲v�v,CP�\:
�<��iZ
�>Od�a�g�fm��?��	��?�q��=�:P� o�L���<M�r݀��R<�M;�MV=p�vo�Ob6��?�oZ����h�	�6�l,���ӹ!��e�<R(I�ȓӦ	T�/
2���cF�?8l o�񟀔'���'�bQ�D��5�HT!@d�U�2 �5 ܸ+W��M���?a��?��P?e�I���IܟT+[C�����FZ)1�6%�7�M������O��D�O��D�O����Olb�.��v*<<��V�*��r�h�Ŧ�%�������%�p�O��k*��-�
�*��T=�x�i�R�|��$7}B�O����A�2�����ܸ�M�)OJʓ����$���qd��s�LDp塇� v����>Q-O&�O˓��ɷ$�.�z�Ѿ��b��	]"�C�	7f� aGO�ZS�U�2C��dC�IvQ�x1�G�$��٠�]�'@�C䉀3k4�3� ��:�qP�>skdC�I�j0�a9Q�Q�>��qw��
�bC䉍6�*���%�;j�]�͂.&�⟄�Vc��5����@!nd�SI�c-���q��2i��5�ׁq�lQ�bQ!�TactGB6c��%�^|�Y���2W+�p�H%*ف"�B�_w�c�����לv�R�bM�<$�` Df�� �P����+�VЫ&��¬�&S󖁹�L_���f��+L<�u��m�,5[�l�^:�hcw��8o�d]���ѷMؤ�z��C�Ec�����q���Lx*l`aH�5,R [ ��:J��RV@	:����`%-;�f  �n�R�6mn����"�.��y֧��C�&���������QJ�w�HU���ڗ��2���~�򯉽}h�R���=��4s�A�ɂ^	"��΁� ���Ǹg~���}B�.	�?V�����0(�&�	$��%�O���$ڧ�M1F��p&U"��O&kFnXR�9d!���=�@���
�6��0s�����yE{�O^P�<�R��|t�R��U�O6�;a��+�*7��O4���O�hjb%@�?����O���O�I@�X�@1�C)�!��H��F�vH
��p|�ʞ2~�¸h�i �3���
i�|�an�F�z@�G�d)�-8 A-���p��\�&��Hg��x���"[vN��5O��h��(B�!�� nڳ��)��O?�D����\LvA��
R
O*����0!�1�|�u�S<v!Ĩa�>(���OLDz�>��O|���	�!JT�*��̠i�����G�{UFpY�������$�	��uG�'�"=�Hـ�i�	j�x���g��$�l*�A�~,��Nc�ԉA�B�(��?a�� @Y�dY�>�2P��K$'��HsKT.}B0����t ��P������b���O8��M�MNl��&c��]�v�PQ�R�'���D2�Ӣ,��TR#�)���)�2Q��C�ɼQ�6L��t��tR�X�$V�����4�?�(O0X4��n��iEP���A��i����޴&�Ny�S��OT��F�,���D�O�S<Xp�D��R�6����P�
�#�V�QcH�"w���)LHsM@�'�����J�~�hI��=Mo0�9"n�
��i����4),��2���џ(���O4�Ľ>	�>g���*ǫi�~ ���~ܓ�?�˓Q8�$b#�-x<�R�EXl�>�Gy��i>˕J�1�~��"�D�+�aن�MD���\y�k��P6���?Q)�(�[�yӮ��__�����E*��R��˟��	�q��s�m061�[�h��4�^wݖ`��Z?��� Re�Xp��A�|}L	��(�$�]�"(��Y��)AO�1��=�I�kDÐ�i$>��S�E�%)�/ Z�`�(Րx"L_��?q��h��6��8Nج�B�Z�B\b�GM9I��p��Wx$q�O
u�<Ш3ݚ^*<r�i>U8����] ��(w�M�$X9套& �,}�ݴ�?����?ٵ�ܩ��HC���?9���?��0/�����\�"�K&��4����.ՔON0 HgjL T�Xd�ӊQ���O�^y���@����YxY,qv�I+m�0GK��z����B\�xtx�
������M�&`ޡ(V�6\8.�34+�T��S����?��O$�������'��O��t�\�/��a[A�/#	�D��"O�H�#�ʒ?`���d��B�\���>���i>��	w}2��4¼
���_���Rf�A�`�̀8$4g
�D�O����Oʹ���?�����4��A����� 7t�����.�(c'2w֮]0 d����I�![�*��ܘPn���ĻP�~����һTN�@ ���� �f��A�'�T��M�� �����X;���q.��?i��?Ɉ��	�9p�
��DꝐ`"F4E��6!�d�:a"r5���ʅlo� �ɟ�G�qO�mm���ė'AxR�L�~��4C���wA��O���X$̄&WɎ��1�'bh�C�B�'s�)@�v���0
�.}�`8�0b�-4lw�����Q"I�G��|@��.��bt���AM�����)ȉ!`�/1&I� !�r����! � �?��Ş�4d���L>����쟈�I|}R��&j�lt� �3+��x{��C���'~��'�t�s
��I�b�H愤)/x��!��|*$�O&4��꣪��=���J2c*	��h����!o�,l8�OGbU>9!�FЦQp��L%�PD P"X �KfD��?Q�
vDxQ��2�3	:�ᦥL��uG�#G��9Y�����8������5�<O\� i� :����� �|�4&r�-2H�����
��#�8y�	I�Q�Y:�&��E��%�	�� F�T�i���QGO/RZ�e��L�.�K��;$����(�V�M��F�;Z�f�O8O��Gy
��hK`��IӰ�!⤀8G��IK���������O&c�8��W :%�w���1'tz#�O"�	B?1�{���:? �%�� R�Ehމ���	D�!� �!T��b��WD8MP��4Ew!�E�{oL)"e���I0d�8 `!�ˠ?��=�T�έySdx{f	�`!�D�L~l��@�FD�M����
@!��݀j���KV�T<9� �V)0 !��:ѫ���Nؐ'��9F�!�k��m*��Ԩb�\��Sj;G!�$�	%a�tP#�O�q��oC�!�T6)c�%�b$U�Tа]�uoG,�!�dUˬ|�F�d��y����(�!�$�7�НI�M������j�$r�!��ъy;7)A��P� *-+W!��ˮM��=є8�:�x��%�!��0wd<ˆ�_��I�e��!�$��8z�ـ'��@����z!��,\����^4D�V��5�H<�!�DCA�$`�J�Dj���,I�7�!�$ɦSJ��g��n+�I�iՐv=!���:�@x�e��k0F,�g_�	!�āL��h�f
�,@Xl���|�!�Dχ#�1�&�V�5�2DcǏ��N�!�D�'R�2` $�?�� �Z"$�!�8k,P�M�5R�_*y�!�� l,��
�K�И����
a\F��a"O��b�풼�X(q���(vD��&"OP��DB��L��"k٘l��"OluA��İxW�E AեL*�S`"O�UafdЯFV�������<5|�"O�T�d��+��a��Jxp�{T"O���#�Ꙃd���[D��"OBm�cS�z,#��^���"O� A�i�c>�A�W�^¦�
w"OFQ��&?M޼0�Ŗ�k����"Of���N8-�����B��*t"O��:t�OAs��iD���f|qq"O�<*e�דx��LE*gw���G"O��C�b\.P�h$�3c`i"O�4�P��i*h����ZD`�T"O��#&�^:`(�W-��Q�"O�)b��P�T�aϕ pqΩ�"O ,sJS��a7-W3;3v�� "O��c$�*E���3
�y�x"O�K��]9�t��s+
�X �|��"O�ܚ��lݺ��K�LҒ4��"O��K �ݚmZ����N��(%"OZ1��C��g��͠�.�t�dx�D"OJ膇�K�T�J�k&\��"O�9[R�ߘ| �YI'����q�"O��ˁ%�$a��C�/Q�_�M#&"O��g���^����6/�Fb��!�"O����W"&��e�4�X=,X؁"O�!@�l[�D��t*�o[�t�\Yq"O^�R§�4>���EN�-ͨ��G"OX4��Aۓ=QSgj�K+t�C"O��m��a�=�T�� ��܂"O��zVѝM<��� "�"��"O��s��!p
D��d-�.�>�"O���2�sҍ��lU�H��\	�"Ol���DA+e�'LK��	��"O�|�%�/�2�a�
͝sq.9�2"O�x�J�8�����[d&�{�"O|H�c�,�c�G�, <�$"Ol�+ ���C����Nݹ7wf�Ye"O��ʣ*ʉ5 ��C6K�X�H�"OzI�%׽028�h�a����j�"O�p�Q�\�+Ql�#I�cTzMH�"O^�(E� 
;$��������"O�4��(,W��
����S���2"O8����L�J�b�Fh����"O�1�`��O����PJ�S�\�h�"O8"���!����\�Q��"O}�W�H+I���q�����%�P"O ��h�&Z�v����	�,f���"OV����,K�d�9&�V��U"OzH�F,�=��Xb
��*6j�ɀ"O|J�A��+pT�٥Jζ| Ċc"O8ј�gA�0�YpQ)	,{zd!�"O����Ř�|Lc�Jй sh}�"O-Y]��ت���x���WIP��y��S\U8l���Uk1v��7F
��yB˗:����#ۜ/9���q��y���5�4m[DC��>�R����y�A�6�u���s.}Ba$^�y�+��Nq���b��(~��2�B��y�Å$%<l�d፤v�H`�U��yb閂f���s3��8:���G���y�Ң9�ҵ(f��?EY� WEɒ�y
� ��PƧ�,U�釧�h�5�"O5Ӓ$����B�ȍ5�<p3�"O��E��F��ْ!�>5� ���"O y���\)���*���r�q�"Od�X��2��]���@�HQV�� "Oα�1"��1_���Ɠ�=9d8��"O��������裢H�mD�!xF"O�{�`��?%bE��S�`C<]��"OLX�L�z�pb�g�@��"O@@�bcِ]"2��@�3cb��d"O��a�̪^�d�ti��|0���"O�(��-�#^~Y��q�$�
3"OZ�3�F�A���pW�;A�R��f"O&Y�̂�� �[c�WK�v���"O��ە��.��٠aH�`��T"O:l#0aAw�Rm0�)Q	}�%�"O��ō�51�~�9�LY�"F"Oy��ĉI&"q����!Od�	�""O!rC2a��P�u��5+N�"A"O���Fb$.a�,��������!"O��K�C�.2�j�@�:�=��"O��anO8D���c�K�	v�}�"O"yA��F�_��(���8M@r�X"Of�G$æ6���ڒ+��TU���"O<E��Ыo�0�;���'Y�h(�"O�
C�J/mJ�b��J_M X��"OL��4a�	L�~E@h>H��"Or���?_l\��7�S4%��j"O���%(-~�Z(��U�j"b0��"O���7Ə,�H}b�ĕ�?���""OL�q���a���3�L�E5�UC!"O�9�2L�4lq�x@`�	�� �#"O��3��W$N2���#�y@�ˀ"O�p+�N&$0PTB���]�����"O��9�g˯E(4��F�^�x�(X�S"O(���L�y��M�G�ֶj*��"O�Xkn+y7��8����bH��T"OnTr�g�CNE��O�te``�"OZ]q2D$[k$��R�TMz� a"O�]:F�1�=R��J��3�"O���A�x~汚@��f��5"O����W6q��r�-QtzəB"O���#�Q�_�|%!�*T�7���e"Od@r�D�C���6`�%����"O�ܙ�D�;�����+V��1AG"OH	�F�X�C��C�K�\��"O҅�A�/v̈́��U+�-=- "O����?c���jG-z;H�"O�����;86Y�!�ʁ=�8l@4"OZ]H$�B8:�A��5&ޘ@�"OPt���g��J���RȦ��e"O&PB�i�cR���D� �:��:�"O ��j�:�2i[�
Q:|gh���"Orh��#<�y���>Bԡ9"O��rl$f����'(P*
3R���"O�X W�Z������'����"O����
1mi���Rj�T��"O,Y��ǵpp�P[e̊��h]e�<�B�R.gY�%���Wx����Zx�<yP/�J��-!�@�+'G��3S�t�<�d�Ђ*z�dQF�ݫF�L]2�g�<�#!8����+�R%bF�Sg�<i6*߉Ӧ��P P|��	C�c�<��m�"�`�p`D�<|���p��`�<� $@q��ULRV���啦A%�"O~=`��M�N��)� �]-��s�"O�HA�Z�!V�g�<K����"O�p�#!Y%T�y E�V���b"O�`[�懅:����℉
?TZ���"Ox�D"η`kF�)��R�p��b"O��!�h����d�)�'@� ͩ�"O�yѓ,�F��cw��H����"Or���-�P���Ӹ9���y��^�.c����"�O@���bL��y�� -�F�j��E7��3� ��y��Ʊ$��p��Ư^�&�kFM��y��$�԰����\�Nd;Vlņ�yR� �F��PfՎ)8�XS$bA��y�S'J���Q��+%켬4 K��yB +G��@q)��Jv�+3�H3�y2'�9S��mB��OfHLar*���y�FϞ8�`i�!*���#�意�y��
%�08	�kV���`x!fO�y��V����	���`Lɱ���y&Ҥ?B"H*�DY;{��uIDnA/�y�E��N�����@y;�MѶ�ɉ�y2��;,�l���MoǶ��`ā�yBG��Z���ŇˣjF e��)ݸ�y��0��"j�v7-ZF	���y�G3� 	��jɞ��&H�y"�I
-c3i��,Ord�f#�?�y�nP~�-H$��'p�����-�ybk͍�*-�dOr)Z�L֫�y�����M�	�L�p��y��� ��6]4F<��A � �y"��8x�d�i�"�#�]�P���yb)Ա���x�G�rs��p�O;�y�G�%��X�C$�bbr0�!�@��y�h�k������*J�J��"H��yR�U-s�.��aH&7�\���N��ybJC-�	�s�cǀ�i4柭�y�B=`��I�Z���#�C�yR%\=6�8P9E��?#�8K�c��y2�����k��σ=R�ȕ���y���<1b`�ggB7��R�	���y�ᛤs�Ĭ���,��*��ҧ�y�*8\��5�!�Α �j�9�Q��y��ݡ�d��$	�h�����B��y�/M..%�rS&�}c��i�R�b�Zw��`p��'F-�y�M�%&$�PP�<�T9@t�	��y�DܳBy��q��1��##���yB�Y�sa�}��!L�#��Q��y�욘X,VL�p�F (mؐA�����yRI�&��Quiۦ%-L`�!�ɮ�yR̈́2df:�@
 RO&`! ���y��'C��E [�G&��1aC��yr^=��XqL�������k���y�,�%������g��XT ׁ�y"�4B�}	R�@�&���L�y2&:U��+�#��.3�!bW��y�K�ܮ)���!;r��#̕�y����K���A�#�\/zU�B���y2�ޭaغ)�2��P���y�C���y�c�-e%�)s@��DR�x���y� ����PK
Os�u��(�4�y�G�`%�`Bw�C?F�� DB�yjY G����5n g��]jRl�:�y�#�1�6-��e�;�F`b˷�y
� ���@
�;}����F55"Ovp��䜳G|���A�y]$�{p"O��@���6��� �Rzr�:1"O�j� ^i���8ƀDax��"O��P�kV:m����7(m�iw"O���s�3���p�'K��X*�"O���t$��AS�%@� ��&EX G*O8���)��pV� �3j�	ZP�5i�'��Er�hDm" IR3(�GԾ��'[|�R自F���Ӂ�@=����'A`��K��$��B�&� �	�'��j�f�Gܔ൨_�hD)
�'l����!R�p[��Y i���@�'��I[%+E6	F��Xb�A%�T$�
�'b�L�Whʘ*��3�E	�:P��	�'L�Q�*gg�x�V� %r�`�'��D۩:<��0'�^��9�'�mЧ���H0Q�	�`N5J�'����G�Uq�� $�(N��i�
�'5H���/�:���G�C6���'�*@`� �\���튲&L	`�'����j�f2Tq���׳f�,`��'�ly��ۊ]�`-#fM;s����'���Ł��&()Ba@�!!|<{�'�ă:vn�Q
.��I�
�'o�=�� �,0����)�a:
�'v���qLJ����Sg�]M:i�'�Nغ���:��A٣mU	<H �
�'�r�c��5LJehtD�
���
�'` M�g��)x^�<Q�^��
�'Z�A���Lj�%��l¸>GT �
�'rR���B$]�Hp�Z�69����'�$�8��&H-bP� �3��c�'��Afo�!bv(���0�dY�'B1:�Lԩ<a��X&�ӳ+s�l��'h�aȘ���d�
-^��I�'����ܭ�&�X4��!�����'���C��&+.P!��-�}l�C�4R��\�f�`B`�S�#��؃��'/T}y��@�!˾�2���j��
�w�R�#VDE3ި���ׂF$J��Y�[2��1�&Y��-ycO.��f�%�A�惇#a|�q��M?5=��F܋y�8��_�'?�`��bI9%�����fW8���q9�H��N�kan%�v�J��6VLx�RE�R�{�$]��i[�"}�'��(��k��?�Qj_���=R�'�x(r�/�/fٸ\ᡄZ�w�0y��4ete��(�|P��6ax���H���[BK�2ᆌQ������=�S"Ԁ�t5����<��K�B�q���5Ɵ1�
=��M�$l!��	�3��	��-P�m0���&c�OL #ƨ��8N�:q ���@�|� �:J�M)V��9XlY2��yr�Тz�l���<k��X�� 5y7�-�u��n����b��M�$�>i��Κ��� ���l�"�(p��e�<�T˞z_ �ȳ��s��$�ת���@�4=9�Y�`���$��ua�:��u�b�-%bj�SWe�+q�����IT�*x'��$U4�	�2�Y6#��mbf��,s��y��٣�e2�'�	�d"���J�vB��Le�}�LsY�r$ě� n��+�3�S���9���9ǈ�c�m·p�FB䉱� )�1�7-|x��&#� Pp�z"��=S�q����;Kr�6�G���$މ:I-L� :��;t�̻*c!��:���qǂA.,rd�r�3r �V�\���0ɇ�J�,�\pD
,O�-i�j�]��}r���H@B݊�'n�1B@�{Q��Z�j�)��0pU,��
Wn���m��:�D`�pi'�HjF'"�bQ[�FTa���Ѡ�"���S84i�$�YU���Gi��OJL�EՔ�¸
�G�0'B}��'f��K��mP}a&��0����f�1t)��F�= �41��>�S�? ��G�}�L�+4nN�Ou(u�*OdKe�)/��*B�B)�XM�ݴ#)L}#�ρŨ\)�%�)�ax��=����FҥDмsB.�>�p=�pa1to��	�GɟRt�9�N�+�邷���m8�Q�#�hB��1R�> �E�U�\q`��V[�㞰�d#��1Y��X�	Pm�O�jq���a~����,M/��k�'E�L�Ԍ\H�P1��؆pV��V,޴Mȴ�`�u?�OU���D�#?�X���D?i��������d�$$���� â�K!�
>a�<1�DJ)�>�4$
�Tb���D�Aa,�tX$)C��÷cB�az$��a����5)����gS6zMbL���4WM\� �Y�y���2)��q�B� �f�x��Y)�(O������i(�s��)�_Ң5*�MȿfM��p�D�qH!��ȨB�������TK��q�Q�Z���(`G�o/>C���"~�f���� N12�@p�V#��[$�-��&/�H`HS&�$���ن�8 �ɡD4$c�G��
�lZ�Cdb ��샾b�
$��N�V�����I�D_�H�Ǣ�>R��`� �%�"dY7�͘���I�C �C≶}��a��kLH���
�*/�b����ӫ~Z�x8f@�1C��0�}�!�� ��Jק�;WS��y�(Q[�<�v&�7by)�C6����F�F�-�BXs)��"�8�b��'$j�E�,O�4��.Bj�2%�$��!i�ĥB�"O�pՅ@&Nk�X�B��k�x���i.���a;k��=Aq��ap�xR�w50��=T�Y�����0>�F�
�}�$+Î��I�Ni��EZ$f������� К��ix������Of�	ud�-$��x5*�2�Q�(�����ql�m���zI?�pՀ�:b� �"�B)$_r�xAM%D�0Ѩ�� E��w	�44��q�f�����"2y.���N��@���D��4V�.$��(
�%*�8�a�N%kht��njDb�D5%���E�:X �<���O�PQ�	ɘ������C���DҠD�4�Ö�U�t���N�a}��t��H�`��2��XV�#&� kՂ־vAؘ*D�%��~b��^t�#ێ'R����_�HOB᳅�[!��違e�3iez�O�ܐ�b��f�ެ+3GD��ȌI
�'M��H���}�`�Jr�&zP�!���d�~�� �d�\a�M��"~JK��yxJ(���3o<[`H�y�-ѓֺu%�ǯJ� �kd+�_剈_?*(���$� �g�'�H��@Њy�� �߰=p���M�����MJ7|OL�@e�ڵm@�]�/�Ҵ����.��?�%H�.]\P���><�zI��C�H�'�(���!����|��)CG��BqKú<�l���%�A�<y�g�` �-�P�Z�/���A�<i�$S+9�㞢|rQ�)��CT��p\b���T�<!�F�7,�`-�r��;g�1C�@\y�' 0A�."��/�|H�cB7q�|�r�$Tw�<���ˢ#:z�zv�>Hθ<H�
�u�<I�n�G�Cd�>���Y��Ys�<�!e_�{t��0)5`ؚpI�p�<�A��\��׌ݶR��<��l�M�<�SJ�X= ���I�7s�T��o�<�VA� 1jL9�F[4?&�)B �`�<	!�Xm���?�V@&�R�<�B�V����[�n�.a°q�]Q�<!�n]�uD@İ��MҥI�]g�<Q��� 7	;�f��s���KXb�<�T�\��hZ�S�G�͑â�z�<���R׶)p���h&Yi��o�<�c+�,Y�B=��(at��Q�<����q4����GξBP)�7�F�<��c��4��"%�"Lyp4�A�V�<I�e�%���S���L���1"ÏR�<YDm�/vLP�qd;Mg��)�lS�<Y���4"tY�!Ը^��Ȅn�l�<Q�`��~s0y	�F�3[Ā��b\_�<� *�)8k�T,rQ�^�$(8��"O9�'D��JC��Se��2d�z��"O~Q�#Z�>^H���!�M�!"Oz\���!.�8-�ψ
���"On��U\�*R��:����;��MS3"O���v/PU-�<�#��lkZ!��"O���􌂧E��3&�ǉ\�&��"O*��%�hK�9���ǔ;1ʕ�g"O2�0W�E�7�FP�"�^;^*���"O\q�� �&A1:Ms' ��b�Y�"OH��� P� �Rf�W.k�f"O���FEF�+�^����=�t"O�<y��N�4� 	�� ˍ/����"O\��U��#+�~@tgP�&!sp"O @�c�L���F�K�d�y�g"O�Y���k�ԕ��d}U�h��"O� ]+8/D�3BbD)G" ���"O��k��1
JY��!�8:I��"O�5��y<�5 ��ʵ|�B��C"O�	CPM]�T�8JP�+$>z-��"O~q����S��]�Ri��U���Hv"O�P�F�:h'������|M�&"O�횐�W�*H�7.R�0�6��"Opm�k�4Rۖ�#h�*3��l�$"OJ�7l�#к�z�O��ʦ��A"O>qc� 8N�L���`L�;�Tya�"OR)Pu� (LΆ��Q�B�56Z��@"OR٠���',nu��捪>'2���"O�b1!V%���V�T*=8��"O��u��?0B
��q��Q����#"O�\K'�'L�6@�7�N�D�.��"O� �q)L�n���#L�o�\�a"Oԕ�)
�w�,��$F���"Ot�n��WT�xPE��;v�l�S"O0\�鋔�� �jF�`���"O�	�F�S����C��Bے�2"O���k�&~��ѴNS��q�"OL�a!	J�VD���͈�ej4��B"O�8`bD�;>�R�s,����u"O`!��`5$FP5��_1 k��@$"O�Qz3�橳��yaP���"O4�sD��:PꜢ�a׍ Y�Y�"Ody!R	,���c� ϷGV� ۲"O����*��`8N��%#%�ha�"O6	��$R.V3���`
�t��0X�"ON5!���=����ƌ�(�7"O�I;�)�V��8f\5�@x�"OU�4�ɇvhn�:�C=q�ؔ�3"O|���Y�>�C�N+P>����)Aj�����V�8?��y�e��m�@�y���w���s�D4�y�ЍN܆H���Ƒ=�]�����y�%
�$zT8`�1;U"�C$H4�y�BP-w
���Q'46!�X�y�.ZLwP|Q�[�1����b�֞�y�)�H.�M����1=;�����yR��;$ϐlT�_53��฀C��y��L k�&��Z�T�� p �˩�yR��J�@qA5G��=*�`�7F��y2)�������;�����o �y�i�<}�`��(Ѣَ����ғ�yr
ϗI��@I��J�{��](M��y��m_�-�5@�n����a̷�yҡҘS�P ��;j�-��B
<�y2원k��Q���.�I�ꓦ�y
� B�z4�S2�l�I��[uR�ys"O��c�c��(&�S��6oP�±"O2%����j���U$�6J1�(��"ODՓ���t��QRD��Cs�}��"Oy���Φ?�hP�B�.yuN�X�"O����*٦f���A$
�L�:��r"O����A!G�\��3v���"OHL0�nת;�R�K	9��	4"O����ܧ��\���QG����"OI�g�P�-puc)̈Y���"O�sCG������+X�.mpe"O�0��G��"86hS����fȱ6"O<M���é
О<b���W�Z�C�"O¼�5�6@qB�;!`�O���"O
5���/��KDA
`����"O�DZG��<<o�!y�M�b�1["Ol��JW�z6=$,��b4�w"O��s�N�1���H���MK8�2"O��1D��nH������AQLe��"O�d[w��x�Ns��y5�%��"O���V����E!Y�+.� a�"OJ���	��H-��Oђ3M֔K"OXE+r�B$(:Bx�@��")�����"OxA��	�9XВ�$Ӗ4���U"O>���D˥��Y*��'�7"O\|9�ƩE�|��Vh��*Rm�5"O�(P�Eޡ*wT�#� 9�Hв�"O~8�B��:,��3�%B񦀪�"OxM����]�*�J��E�>؞m�"O��� � aYf�Zu ��E�vP�c"OH\ �⃳#0dt:-)��Q�d"O�%Heȷl�`��������"Oh����	�,�N��V�L)�]�4"O� �hL�j�E��G��l�(���"O �Kf�rT䀜�<�9�"Ot%0��޷P�5�Ce]�js�q�"Ohm��h�9E�LKĚ&��y "O� 1�d�e��-�J��(����"O쐑S���(�����!rz����"OlQ���8���R�@u�="O� � D[5!�10E���Qy�"O�9��B�p�E�a��|���s"O� �'�Y��$��--p��"O��x��%t��ph�#� ��"O��RDD۾p�rU��ƾ����`"O������F���ɦg]T'�`a�"Oʐz�Ǖ%k����f�#q
�iɀ"O��!�&�l���B#X�a�NX��"O�0��G�C�}� `�}0y��"O����D-m�hRaN��1fvA�t"Ob<�&�wm��#A���E;6�k�"O��uF�S+jXB��A��{�"O���ć�h��c��6\G���"OfU2p"��
�T�� æ1��ѐ"Oʑ@#���r��a��̀
*��H#"O���&(���3������K�<�)�?2��q$�*�R��d��p�<�\(z`�C�<_\41;�GGB�<9�y�R���FʎE�#�AB�<�Ѡ�v>ژh!��0!�eh�{�<Y`�P�,nu��V�aN^��L�<a�aY#3=�2p�1o���ːM�<!���B�V�b���/S�ɑ�e�I�<�原5bΔ���3~�X9��^�<� ��3d�-v|�)Q-ȯOf��"O���6m�T �ˋ�^���c"O�Ś.��G�V��¨�{jr1sb"O��FٍsT��W�I/0�R�"OX8ʂmI��C�KM�V�x3�6D����×�}��yr��Nu�ܠ���&D�\#'�,��qQ��R�RU�|��o#D��B
�t�&)v̂�S��x��"D���\�I�>x�6��%?��A[�:D�Tsb���qUpP���cp��xuk:D���뚐g��I D��I��-yŧ9D���.�9Q�m:Vc�M~��0��*D�T�P
��s?Υ���P�bL	¯4D��
�����l)����^4r �-D��K��By�a' 
>:2THh��%D��#�JΠoz�ؒ67�4��Ҩ$D�x���f�DX��ćr�$����#D�@�Q+�J($,0��D*�]9�7D��Y��Ԉ�2�1`BĮ_���f6D��2N��T�T�A]���j3D�$rn�v�tۗ� 56�9�k$D��3�ޟG�L ���6�R1�E#D�� *�(Z�5� �'s
� 1�!D���tκw3�DJb
�AG�a�?D�p��a�P�4�K�L�j,�	���9D�Шɝ���q��gL�y��Y��J6D�X��BT�9���S(��hZ���2D�r3�Ӟ{ą9��u��*D����nXk�-��KL'o��ŀ*D�d G�_�x��	��IZ��PsF�'D�����$sB�'�#������ D��aAzl��MȔoV=�c">D�l�唚ግ�A@ٔv��QYv�:D�\j6�0_��+W�c4���ti7�I^��<�ʮJ��9w�R4;�숱�)D���� 7dT�B�Y��5D�,A�@@�9�tD�54nㄠ��4D��顄���U��F�|�(���3D��(!�SC�`a��D�pt�3D�`C�C���GEI�6,U�?D��N&f�����Ŗ$�(sE=D��;d�>(Zq��k�V�Ȁ2&�5D��*���]����BTy���D3D� x��<O/�〧_NtfQ(3D��BwJH�H��3(07"�mf�<9t%H
h/���1 ��r���J|�<y!�]�>�����֜����ϟA�<ɅȆ#~�XF(��AU���@X�<q oZ�s�b\ɱlW�I�����\[�<!���7�zi���Sq�@�`��\W�<q �h2����ɡ��� ���V�<9VO��j�Hc�A7T˲�0�W[�<a��D�Ԝ�����m�R�*Uɓ_�<�!� J�\�����26���B7I_�<��4T�D��@M��X�DΊV�<c��.,����Vg�,>�!�PJQ�<	�	����`�hF��v�;�-e�<A���>u�@���դyM\dA3Ef�<����5vs�1i!ܣr���g�c�<a���a��`H��ң"_l�:�"	c�<���)�|-�t�ˈT�:��k�E�<qu�
�,,BP�ߘ�� ��L�<!VHR�}�*}�Fb�U���Iq�<�bÓH�8@9��J���]���Zo�<� ���U�[�м1 䁳so�0�a"O �%�Ⱦ]i�� 1�l�l8B"O��K�'܆(ǐ�����"lR8�"O��wj�/D�4�R�'ܷc�|x2"O�Y��a��WȘ0��S��)�"OP`�,'w�
<���R�l��("O�Y)�*Ԩ|�:%�� ��R[����"O�<���0}��7�O(>��9;�"O�)R�[2^xa㮈�k�����"O@�'��.B�)��ـgo<�AF"O��#f-W�u��x�"֟gj�Uy�"O�q�׋�	J��c�ēBKF8�"OJ30�0y𾩠�ϚB4���2"Oqr�-U�v(�)1�N
�)#��Ӏ"OT��7�b<:���u��2"O\�"C��b$H�B$���"O��;�
��x��!��?E|@�"O��Y�Iחo�&�#/��9q<<
�"O����7 ���C�$
�Wz��"O]S6��+3���(7��J��B"O��MR:����'FAB�(D"O���V�<�R�Ä��`��4)�';����O	�(�Bb}����+D������x�� 7o�3g�����-D��!�I��>10��L5S�p��C7D��Jc�9l� �'��6I�ܫ�5D�,�R�[�v�Y��S�-ah`�Bo2D�0���6'$���K�2[�h u�0D��PQC5V6��9eb�6a�`x)�-$D�؂���#*۔��eS��X�xP�!D�أ���<s���UI��F@�r�!D��!(��@(�(��F]�С?D����,J5&����	w�]��)D�` ���F�ꗅ�!��"(D���h��-E D�3*�uDU���;D�  �Ԓ�,��4C��V4�|s��8D�p��C�0Vt�Q��R����h8D��� �"N�%�`Ć������@8D��Ѡ�5t�Q��">��4J�3D��P �Z��Ѵ����*�z�?D��xe��u��3d��aH&�a"D�� N�o� [S�K ��V)=D�pR�G�f��¨�8,��1�� D�����r9 �n��0Y���6�<D�D+#/�����S$J�i�~�1WO D��{A���lE�I�Ē( `���*D��`�H�?�$�����D�8���'D�p�捀%����P恪lB`��O%D�d󀍙� ��pq� 	 >�Њ�g>D�rqO�# ��;�Bߞ%�v� r�=D�Ȉ7���va�(yRKЀjJ���.D���5F��-L�Y�K��-.D����gP6,�|k ��e���x��,D�d
C,I�!�l��p��yRBlY��)D�p`hM�9�P��kT�l�Csg<D��C�@�[U`X��?��Eړ�%D�l�`��w~l{v�͛tX��a D�h���ӑi��]�S�K�f�$R�m<D�\sA�F"m�h����_I�)�"�;D�������f( H�N�:UV��h7D�(���
2f��G��>�z���l8D�H{���_o���$I8"��Ŋ��!D��xah�K~xIpP���I �>D�P��hR?tFČQ��#/߶��q�=D�� ��K�
�cvT8qaEy!���0"O~%ҳ \$R���T*��,�\X�D"O�h�1��,kn2"��3�Ҩ�V"OHP��@1a��Qτ,Cƞ���"O�� w�ӈtf�\Y��W4j���S�"O���@DW:1���'-_|�t�R"O̠�Dh�KnL�ᖫDsP�b�"O:�I�h�Vna5)�8w:݀7"ON`x�b�-:�M� ���-h���q"O0�[�KծG `�"�)8"�"O�aʘ�MѪp�J�qL c�"O�� �d� ��ܰ�(�'liiW"O�Uw�Ù5��	S� q}�#"Ol�9��֮{S�@����50�P�G"Oh��n� e�X)Rb�*t��+�"OFUq���g���F�/��p�"Ov�x�F�(|�ո͜�z-^\��"O��3�,@/R���z$vd��'�:��tIȣ1�>�;��X!R�X�'@�P�
���2��t��U�ؼS�')�IK�Òōua��Md�T��'�d}�A$z �}�+S��'��th߸.������>Us�'U��Oy@�jQ��'*x��'� �ǫ�'����)l���	�'#2�"����ʴD c0p��	�'�r��6������L,8M��'�U`����Xq7L�2�-��'�$�F@�q�Z걎��v9@��'5z] �gI%f�R���a��8��e��'Ԙ����/4�� ����B&�ݰ�'�Tx�i�=TJ��24�����'~��S�� o��
��()��P�'O����m�9)O�X`���!�~tR�'�BvbD^h�K��}p� �'�ր�o�6x�La4�O1��(
�'_��۠ �.������9(�0"
�'v��agC 0�P-���#�����''b� �a�-[��a�i��J�13�'�V1W�F4O;DL��X�	���'Ip��j Oh�3�c �tձ�'���q܍�V�8���P��4	�'�X`9c��%a`Z)£Ƣ�@�h	�'�(�8��z�@�"aΔe74�	�'\$t�%犳8%&�P0��5&Tx=B�'|�|��+����Qp*Fx���'#H�C�
N�Y�&5V	θJ�5��'q�!�fX�:�� е�\�J���'1MQ㔠f��i󓨈:G���'6����)�H��#^)�'��xPDG�2u0ACv������'���w�/�LyT�H�ȑ��'�T��@H�k�T���h֪>n�p"�'� ���mE&*ۂ��	:-�=��'T�Q��7o�h��Ѵ+P���'p0m�#��>���AΞ�*?4���'Y|l3�,B	vb�ҕ�<Jd��'�
��ej�=�� A�E Y�T��'I��0Ɛz�$M�����Q#�d��'-��(C�ޖhCp�[SO<eN@�	�'�|���Ҩ,hvmX3�T3ޖ��'l�y���]~x�B��(n����'7�[�!ɀl<�AǄ���1��'A�R`��<ZΠ�瀏�[S(5����  )�ND$��l�t�ӪմӢW��;���Ӎh	��Xq���TĹ���j��B�6&�T��a��/�|,���V�8�O����K�M�`�9��Z�D�mS� S�����O��;�:cKjݪC�D�1���Ѥ"OZ	�UGZ +�uH��;���Z%�	�:��>�`��9�(��(��q�W�-D��g�/a��F� �Ҭ.��B�	�l���U�ץP�
<A�io�B�0f8��%)��W\Z�G�<�O����M�y]����X&M�h\A�C�54�!�_Na�l@�-�ɶMZ�b�(�!��Md�k��I��B���;!�:|�8+u��<H����o׫_!�$H���=�#�?]g* {�m�0�!���!#���`��ܓ{W��R��F(B!��4����[8VE�wFZ�&!�dXj_Q׮�}B��R��8P!�D[0�>�$ν�E����
�!��HDjX���хb�j5A�A߲�Py� T�TI��ॎ :nK�H�PeP/�ybO	�n^��g'J�Htdڰnݪ�y����a��'v>܋0�,�(�R�'���QP�ؼ7�Y�O["ec�-�
�'�`h!�����HGT���(��'ir�H�c�$�@]�V+��lez
�'����C�A�b��Ơ�9L�:��
�'`� 7��0���i�'v�j�
�'v���C�Kv��� A��C|�8�	�'�Y��9���W��<�q�'zr�*�)�5����'�D4����'�*��bp��A����C9`P��'�Z1�j��~�~�va�J/:��'��L�Q�[	d`���k� �x���'Y��9%�W�fp���ܒa��'�vP�'�+eT��x˛����J�'���y�/
C	�0m�����'H�<��E���8��	�h(T��'}�0��Y"�5[�▻I����'Oƈ��$om��p�aJ>2�0�'f�ʤ���-k�E�0��w��̹���=�����w��:���c$E��o�b�ȓv(usE&
��|ܻ�FĪV�t}�ȓS�0񲤄eX�R�'ZS����5���1ħ�85C©�2/�O:��ȓ$5�-�р�:9�z��sE�X��]�ȓ_�\���R�?�!��I\�sH�Є�)Q, �U�[�R�|\����-dbĄ�%�a7��9�iB,5.�`�ȓH�T ��cU��-��G��qtt��q��K�%�*P4ڶ��g��q�ȓU�<Q 
0�:��H�|T�ȓ/��BpD�?z-B�N��\q��sJ���p]o~��u-��(��y�ȓU�
Ģ"�$W�DH##�x[(Іȓ%L�$��4��1s��Ջ`��̆ȓ4�|5�֦K��Q ��L�Ald��	�����w;^< �/�8�<��2,$��l��8ޢ��f�<�H��mלq��A�0��ŜVVl��ȓFr|l�chG�}�5b��\T���8Y�9y��|�2��xY���ȓ�2�`��q3J�,Қv�l�ȓ R@���M۷X�~�bŪ��LXd��S�? ��
U:ir!ec�<bZ�"Ox���I�'�����+�ԫ"O�A��8&��I%T�{L�s"O���rh�L���S=Q�t"O��Oǖ�T՚�oO3t��![D"O���w)®v��e���Λ2�\�"O�L7��a5+��\�+���yR��#��Y@L���`����y�j�QPܲqgU-g�0![�؏�yr�͍��]��/(%Xm[�B=�y��8}��M��E�, �!��aD7�yb%M
yZծ�>:�ES,:�yB�ǝ0tb��N����� �R1�y�N�<��$J�E���S-[�yb썷{��i!G㔋
�,h�B���y�/�y�mX��9�z����y��K�>��ԆO��n�Ū��y�G|��ch'�D�X�y�G"$���fhĒX\���Ӥ���y2kO�S�舱�ڿR�.�k�L��y�K��H_*E��IN<N�<��sI��y�B��c�H8PA��E�&1�áF0�yR_�H.ZɁ��>�$J4@��yr��>&�`0P2"�!7��)�-�y��߫cw�D��@�5��X�v�\��y�#G6�\4&�vQ��r�.)�y���4�ꉳu[���U
���yҮ�͘�B�����B}{e�Ө�yJ[&8�a��"F"	f[ �X��y"���0�s0%�5�����y��<�H��bK�w%N%�F��ybL�?uK���1�Z�@@�d��y�>�>�h�[�x	�UQ���yF8'�$X:��xs�Q�ø�yB@R�,��LV��r�⍁����yRX�\�x�c���6j�u�s���yr`R�LNt+��S�lװ5��m�=�yR��,V��J�h����q���y2	�_rD�[��^����R���y�a�7(�D�ab��XuF���I�y�G^�i�dHR`���'��|K��ڎ�y� �N8Xe���R`�4 _%�y�k�.eRd��&-�:�U���y�@�^8�H�S`5nN�9/�=�y�(�c��h	��.DA"Aܪ�y�L��Z���0`�<X����(��yRh�u5R`HPe�3>�S��[��y�`��OG>�+50���8�ƌ��y�@��Y��(a���@:�ydR�ȶEQ�ǎ7xPU�����y��A.Z�
�A�hE�f�b�K2c���y��Sb|=����7r��л�׬�y2��&l�F��
\<>۶AB��_7�y�+8��ࢵb � P�K G��yō��v���zqT��'n_;�y�⇃f��yk���q���C��H(�yb&J�GI���e��&Y�Y�Ɓ`&]f�&HnZ���l����)�<T��d�Ob���h�4b@��=#��v��I�Eh�;<ԖY��d��k�4l[�dX>�Q�'l]�# *)������g�����4mִBԣ�9*�<����^#�(L��`�+���5�dΎ��;7�ě��Lx���;$؛����?�V�i!N��?9F�ܴ��	e�U-`E@��̖m/�����?!�52��N�q�B���gy� �����d�$�'���b��o�d��?!�;1�h���_�d��]a!��W�"lC�'	Rj�K�q5�'0��'�� iݽ�IϦ��ce�ySʇ~/t�'�T�?Y�$W�̺�a5d3Ȱ<� b-*����G���U`
9��Ѡ�[�B�JQ
�a(fޕi��?��3:�1S�	��9��	[~4A���=U��p�fʲ�R���-���9Ӗ��>��us뮻>Ʉ��2֕.3A젃���a�V��N��h��ݸ@��)]of�Y�*b��-S����M+b�ia�n{ӆ���L�ɤ|���S�(���A�	pb7 vB�yjЧ
��<i��vV����̟k�D��OWAL>�{�&ޘX|f}���n�taa��">�)V�[|�'Wf"�T�p���ql�$��4Ȓ �G"	S��2$ D2)��I���	�Ox�0��'z>���.��8u�ء+�*;)��Y���3N�L7-�Od��?I�R�'қ�#Q�:Z��C���P,i�Z�Z=
�$$�O�TabO�|$4�&鞊5Il(J�O���!�����'��	��o}������,�O4����M�nG�Us�N$4��YB�ƯGF���O"��ҍQ�,{u \}�'����pi2&	�
~t�	��
WE�$#=a���e�tR�i"*��@R���i���K� �V�d��3�(Ѻ����E0e�P�㲙MK��ixL7��O��N�~9��غȒ�
&k�4�8i��'��'��)�矄k%��H�L8ptb�*K=(���G(�O$	o��M�ܴ[��x�c��"?�rç��'�JA� '`Չ�it��'��Ӣ�����ҟpn)xi��JF��%|�t��ů�9B�
�"�P���J�h�4�MK�An��˧��INE?����f����wN x�>������=I��d�n�G�ч@s
5�c�s���s��P5e���e
1u���V�iMT���>����<��]��M{�o� �$����	�f=X3��|?�����'���p�B�L��h�%E��tX��<�I�� �ڴ&Y���|�OT��!��11BB�v<����QӸ��Iß(�"�g��|�	П���֟��ZwҴi��,�($Y��f���s�*�Oh��r�ܼ �� � tas� !G�@Y+�����ȼ��L6lpRT	�,y�����(�k�Tݺs�f��CSy��]�gre!L?S�~A�/���D�)`�r$xӢQ$��	ßh�'�v��V�hi���K��o�J�0�'�a���[{��0*��?́P��	!T���l� �M�L>Q����N>!޴Qnl� @�? &�m(�"O�9!�͑�&�j�K��#��<�&"O���A��#;9X� V�	~�D���"O\tÑ��;S�BëK�b�@y��"O\U�@۝w�����K&U�<��"O�HS��*bh%�@�ٯ_}���@"O|��_2"b!�1��a�U#6"Oj���Bե>Z��W�dO
��5"Otȳ�C����p�(��t��}�"OȀ��+�yLh�@Ü	A�ebF"O�(��]�m��pҊũQ#D<"Oı���	�2� *��|^� "O�X����A|p��#���Q
�@�"OX�q�x����� 4ੲ�"O@�k�13��9��H�o����"O��Hus�M�uǃ�m��ms"O� �p�u���	�:��G��,����"O`tR��_�4Ԁ�ґDQ a�@x��"O��a�D-k8Y2�hP�7����a"O�X�O����(3�N�\��eK�"O<����Hz_�h�6FG�ƁC�"O$�ʱ�De9Ԭ��Í�fZv�*�"O�<"��Hl0�����A�Q�l"�"Ol Hr�.R3r���֌sB�Z1"O��B�-�`e���֮�
�A4"O�& ة�Ơ*�P2���z�"Oz9w�&nWPY�$^3J�����"O�Tyv ��.[
i��҄�Dو!"O�8�B43����(Q%L��d�6"O�آB�ǯyh��AG�ԕ9^�e��"O��[���3)4���%�6e摉�"O��#�mHq���nP�\H���"O&�+F��P���H.��}ۊ �"O�U��ߚ~�4�5- �.���"OvP�ҫޮd�)��~�,	��"O8 	G�5(o�"%��<���"O�P2uO-.,�}@���6�Ȝ��"O��jT�ʠ;A��R噷e}z �"O���c�K�o|���B�|F�!"O.e�R.�=`#ڽ 򋕗��c�"O�1P��[Bqza�G�P��`��"O���b�>	�ü8�@(�A"Oq��N��#v-յ@�0�hW"O�5�A�#7l8I3�L_I^\dc�"O,�B�-EUm�q��@�qb�"OQׯ |8�e�	���"O.M`ïK�'x����Aڜ� "O�)��	Ib�.�x ݱ,��a"O^���0\�ycrO�2��2�"O:�Z	�� ��ŷ ��<�5oi�<�3�Аv�d�weU%�]��+�o�<ѥ���Y8pU�W�Ҋc�T\�V��g�<�r, `�6a�CAf�e9��Sf�<��K?=ꞹ	�����Y9l�b�<���ܘ�nx��茆E�����[�<i���N�`p0�ܨ}�i7��c�<I�dY 17���Φk��PzU��E�<9 ��h���A�&_b���C�<q���*Ѵ9:��P�'Qj�9d�AA�<�լ�,>���� 	>d��uH�<�^�~Y�:w�ٹhD�t�P�k�<��H*J�P��j�1ed�ܻU��m�<�aC8[��9j��۫'��P�L_�<�&N/"�r����&Z���;��UQ�<Q��K3�������J��CqJ�X�<����?�)bA*V\�P�K���~�<�뎏D$v5��&L*cV��%�a�<�G�r��H�m�[�d���,!s!�D�'QsRq1F��=z
��F�6Y;!�dvU�#Eg�a����%mL`�-�ȓ=0�A�톪7Rrap[�[C�@��F�"W���a�cW�D!T(`Q�4D��@����!�fA8�j��?���(�d D�48�IO�MJ��Q-��0 "]�s%=D�xq�
Y�����'(���b,O�<�6E��.TMW�Œ)��y� �U�<��ʃ!3z�r��G����&݀�ȓέT�UeA�(KF��t�lY�\��6�l�bEF�Xh&�`�P��2�ȓw64 : �&Bv��XC-���Y��S�? ��Qc��J���(�JM"��( "O��rǅR �X�P6 :$"Fp�A"O��B�ن�t��$���؅�a"O(�k�]#Y�4�)��C5;�Pc�"Ot��Wd�N��|�R��r�ј�"Om�Ef�0	�MgdR�f�H�"O��(�`)OĠ8X���=���"O�A� zJ\�Rc���>%�O�<A���C����@*	� MH(��Tb�<�D:u|���G�c���P% N\�<i���4B�h��-�K�2�"D�b�<��ʹ-�`M�G�y�P�Rv��X�<)f U�����fP&�P��%�PT�<�˕}������F#�rR�P�<QD���{��)y�D˗Xf�qJG�WN�<Y1�Mƺ�c���M8 �h"�S�<��K	17l0���a�n��^h�<���?ǚ�H!c��X�lD��Sc�<1g!΁(�N��po��*��僐�b�<!X���pF� ;�L!�#�7,����_��S��_+w���H��5��5��~8��3W$�8XP �ƥ��ȓff`B��F��<H��+
A�$��XO�YW��A"h���c�/
��ȓN���N��\���P�+�`����3c�J������=w�!�ȓN\���c#Voέ��M�!����
줅ӐkL� ���kJ�|���ȓ��:jx�a��oy��էl�<��.�,x{0U)�Ƒ,\7m
fM�Q�<	��@�hf��k!��-~����R�<ɃL�o-d��[>7h���V�Su�<�&��=f�|}x�{\�`x���j�<1qG)�"� ���\p� ��|�<yEM?G����Ugj��c��w�<Yr�
�Pz^�Ap������q�<)�K
�Q�\`��jI0��ċ&�X�<	U"�'xA�Aѩ������R�<i�N�"U�u��n^�m�<�8C)�Q�<�*)8��i�W�T�jC��M�~B䉆��b2�Ґli���:rHB䉷4[��0��S&	]�l���B.i��B�I�I�X��A@�C������=M�C�I4O�A"cK�0�v5��اC,C�I�^m���ÁäKj�¦���\[<B��-l&�* 
�2e�H���L�.B�	5��A�D�l�ЁcMh�jB�ɶ'IV1H�jG�*8�=���LXdB䉬U�j�Q�2�~���j�s"xC䉂l?��Fo�H�(�pf�,~rLC䉷'��Ds`����
ہ:y�C�I�'��u�0�Ҭe���C����C�Im�`!����^R�,��Eըi�B�	�	��k#,z��j����Z�B䉣&N�x�U��ɔ�1��C䉴:=���r�O^P�*��8G��C�	$4$��"R7L-�Q�.��C剢Đ��� ���k��
,�!��׬on�����\-�5F�T!�@�u	ᩌ�)r)���A5!��i��ؓp�H2x��i� A,!�;c��' �	:��t�O�v�!�Um �ႫmʲQÁe�*j�!�D]�<��!3��
�Zx6�Ԯ\�!�� �d��/�?)�\���M�9�rT� "O�h�t/��.U�C&��^���"O�YKg�م^���B$'�<�4�s"O��w�	-�2������R6Ѡ"O�`�A��1f��q��[#�d��U"O�H�A� @3���R�[������"O�`0O?�F��P&�
s�N��"O:�r�FMW:� C��/J*�K�"Oڨ�pJ[q���BT� �p��"O�(��J�_W2Т����lwd���"OLa��\1#ĉ�7�Z�+n����"OVy�oL;��ehX8~�V��"On�Ȣ��_��H���VL|�!"O�h���;z�E@��S۔Yp�"OV]*��'�X<1�O�_�j�@1"O�Ա��¡�Jy`'iX�{,�""O�PHWHX K��Q���)�<��"O����(��T�D�@�I*F~�I�7"OqRnU��kB�/v��["O�����A�nDQ�e�Ti6"O�DP3�f3� ��!�Ak�]:��"D��6B�3�N����Hd�A�a�4D�8B2K�LE6n�-�xyw�.D�,�eJ�#=VD8��F:����+.D��� .�W/���A�L���G�+D��R�E۴v��*r�����K��3D�ЁaFӔf��U
�fZ�Xk�=�#�-D�31	��0�d�з�Y�=e�,D��"���
�����/��p=7�(D�� ����q�+.�%!D�aS���T�f��$/���c��>D���h���ظ��X=�Tڒ�;D�Ը��	�
�������Qz�a�+,D��rb��r�� Z���*�^��&a+D����ԪG�!�!-O��
��'D�����&��=(Wk�"Ͷ��r�$D��q��B��$A��%��t��EH�!D���
�8J�c-����"D����H�Z�Թ*�i[�1`]�'&D���w��&�\TV�˽6H�an8D�X�*�;6Z��q�I�vz��ZA&!D�z`��7Og��1�-_l����#>D����F�?LR3���L�h!ڣL<D�|Brㄦ1���Ѕ ��&B9�C-&D���`��%�>`1���9� 9��(?D�$ٴ@�o&�U/� <��e�1D���`��0���"���p0�`.D�r��>F+�4��'�	p`Q�(8D�\+ҡL�v���
>sI���Ƅ;D���mۏif����G|�*��K-D�D҃����\�Z`Nؠ�a�� ,D��*#���\��]�e�V�5�R*D�8@���,����eh-��Qwh(D�����
S��0��иxT�;T�'D����F�q��3�d�?;z��'&D���'.�v|��"cd�~��|1h#D�\b��!��q3ŏE)R�<��P�?D�Dk%�ڃ ���ߤ,!*K�H?D� h�D�/jҤSu
P� D�� �"D��C�GA"$�d���bH3g��+��<D���P�"�yb*��`@�4�;D�tKekN�[� �(2��a�V�i$B:D�xP�j��&�:���e� ��ah7D���C*��3�`��s�Ɩ-X��'�5D�� �Y"�I��w�x��┮s�)�"O�����@�(Ŕ-ⵇ#o�zِ�"O����ܘ^NQHw�^�B�|��"O, �r�2<�6�G� �J	�"Opa E�F88�.P��L��'� �A"O�}ۀ�A�\�cԫљ4��}ZT"Or��Co�>GQd��2�4�FI˥"OJ��LD��=i%��T��m�s"O>Iqa�]�Iz$��j��-P�"Odq+n��Z�A�䀇E�D- g"Ox��b�r��#ƂK�ؘ�"OtPA ��y8��w+Ӌ/x6�;�"O�E�Ɛ��r�%zs��#"O���"��ʡ2d,��cd�y��"O�`��<��ڶ�X�tyXC"O⠋�MO~��b�ꇹWC�YT"O��[r)�k;�X�䆓�0����"O���� �H��4O��Uf�Y�g"O�XD�Vs��i��.SPD��"Odl���0{T}��H	^=�uCc"OH�P��%/����d���Ih1"O�8�֧/Dz[ P�L�
�1W"O|9դ�%��y��������rB"OJD�����W\x�S;Tn,3�"O$�@!협`{R]q�ƍ�gf�"�"OXȆ�52\����ȸX+8p	f"OP��7-�2@-�P(��C#~��"O��#A
W�{�d-���"v��R"O��i�e_TVZUPsdݳ�v�"O^���+� >0"C�o�l6"ORPZ�[x����F�Q8_�t2W"O&9� ��d"B-��j��3�n���"O�qr�NϘu�*U7'�1��8Bu"O�ˣ��:Q�8��PިA
�+$"O"T1��^<%�m`�ƈi�ا"O�y�ۭ=�E1f	$,c< b"ODP��{FDI�.(v|��"O�p
D!Q�	��5�+^�5�>��"O�Q��Cs�F�Ie)Ŋ!{�5�"OL�A�B4Ud�h�V�Tsd���"O��K�A�/Z�9 ��,��5��"O$p�
�1`.@	�jG!vЩpq"O|@B@�s(~�g��xbH5ؕ"O��3�[4O殬�4��s�:�q�"O���)���3$��'�t`��"OV��P
]���2�"�:��2"O>�@��*_kT)�VB«~V)0�"O�xCtLF�4�:1�[�C��уb"O����eئg�HE2T�|��81"OpDs�M�,-Κ�z�-Q?H��U�t"O���M�/p���0�a��d;�"O��v`V3@ `J�L�C�D(�d"OBL;�K[�>2xR�j��Z�� "ORYgQPD�x�T�1��"O*�;��\
'�&l)wH؞)i�@P�"O����� afi�%�%@F��6"OP�@�O�� ���P�@���S"O@Șf	 ?���&��Q�%��"O��1SÑ�R�� B�W��ě�"OJăԄ�=�T��3+ʶH�"O,��a��q�d�S1��.Z�4���"O�(�6ϯVz���eG��Pz8ӥ"O� ÂLm2P��B�_3�P!v"O�yIK[1h�jmx�V�s���6"O� jLסыO��Q��+��m��"OJ�Ac���~�y�	�v�SD"O��!N4-E�y���%I�M�r"O�d�s�*6rzI�� �,>&XZ&"O`<��T	?b���.��b��ȱ�"O�I��^�I	��@�?	zp�6"Oh����
W�1�#eS)As����"O�e+Q*�|(�(��Ka�08�"O�PS�(������V���p"O��'��.-��(���!��"O��qd�b?�0�㖲r����0"O4��c�Ҭ d��v!��6�Z	�"OJ�js��/+$��6:φ���"O�<�F���@Z��H/�h���"O�}�'��w�|ArU�Y n�\�!�"Ohi����!Y~j��ǤV�V����"O��`��JW
|� �Q�~H�Q�0"Oލ���ס]��q3�`��Nx�2�"O�H�riJ�9,0R��B�q.����"Ot�ɦ��Q=�rV��^�0U��"O���7-�^����!�AQhTD"O ��v)՜c�v��'9Y�E��"O����<\����� d=&�[s"Ox�P�I�/Π�p�
�+6�U8�"O��0-�v���#8$�\�"O�X��l��|��e�փ�� ��L��"O֬�S*�=5f�Y��⋧Y�v�!"O��C��o�2�a�����1�"O`�'�H
���i���6u��̋�"O~�gȟ�T x�
�.�$x@ "O����E�D���%N�,���"OT	��kW�i��y�S��"���"O����*;	���I��92�vi	"OQ��O�X3��9T��X��d�c"O�<u��-��h�E��3�¨�r"OXU�'	�V�A8E�6�ոS"Oj$�&�'i��IB���(=B��@`"OB�"Z"���R��'�yb�"OL�����c�t�3�"�m��y�"O&�"6���tVH�b��t"O�P�q�6�����7x�z��"O���`Ȉ�+�H�3��a)�"Oܽ��/��MKC&Ɇ\�� 0"O0uj�5����v��A2�$ZV"O(�x��M)>���k�$r(�"O6����v���z���Yf�`"O��sw�ӷ	�~LJW�	�kHly�5"OبKA� UU:q��(�)�x�1"O���U����v����B��=#�'Ht�0$���l�CF"�j��A��'���"A�N7"��ѥ
ܳL�E(	�''@��q���ʛ�l�`s q�G$D����EX�GJ�"��4�,D����q	>L['F�A�\�>D��`A�7n�=�R���H)z���>D��Y&H�f���@֬v�LU��/D�|����8z @��]O���!,D��"�(�)(�`����ͽ#���q�,D�t�Q"ǕE(��t$NȬ �C�6D��+W���(����[U��*wf/D��7�3>�B\x��=�dT�B�+D��ţƇ���醫̵w����a!.D� 阞h���'C��P`��-D� �"#-0���C�	�"������(D�� �T�5��.[|�$�E?2��"O�0x��@�b:Ĺ	3ͺ.ϸ��S"OJ����(�7���yt��&�.D�@�N+5i(�
��X(%�L9���+D��zQ�^�ϖ�C��S�|��)D��b��k���#�щU�<I�'(D��8�#@�\����`�`�"D�,:��āc)*�)�m	�~�&@j�,D��`�[/l!@*�̂�X��R�� D��s��6 �D���n�;�
� `E#D�\��ƞ^t��TCH�k(� s�$D��KE�M�`p-�c�Z�:e�U5�!D� �Gc�t՚X��m�8
�����<D��
�a�3Ae�ib�D��s�}I�j9D���##6tJd��)�[ў�r�*D��+PO�S�а��}�@A��5D�D��̯�б�E�8�8�e�4D����֟i�F�	ƃz+H1�� 5D���p�ŧ=|�r�$=��#R�.D�DBD�?��$�d��� �S�*D�p+�nS]t�b�͎H�9�D�<D�l��.٫8�LE.�s���kvF?D��`#�*4����AՒ��a>D� �#��@'H�w��85�I�eI<D����,�t!��	�җ1A:Icr�,D�p�5���.3���]�.MЕ'D��ch�|@�L2eϑ!�ڝ��(D� ��I>>��P�0O,p݊4��,!D���む6;@�)��)�
�zjË)D�T#�c׹3^0hVO
54D�s%D����L:bR��
���q1!�XCWrC�b܄,;�h	E���9!�Q(!�Ȝ� �R/��Q��I�
!���w�-� 	q���[�	�
!���t���n׏*�X)A��'q�!�׮?�,K�m�KlPf�R!�DE7c��0�$��$Z���"��@!�dE|69���?L���f׊Z�!��j�
���n��c�������!��Ʌc����%�?&Ξ�a��>p�!�]&*`���Mד#����(5�!��iI�̋�aZX��Y�Wß
�!��<1ޱ�
�#%��̂#�P3`&!��;"m��s���)�\�S��ѐA�!� >i�T)X"��t��ȡ��7!�D[�+�z%����hb���9l�!�Dʤ��Pt)�,gD�e�C��
'�!�D 
~֥��o�7A&RelW:k�!��֗I����A��^	��*���>!�D_*	D�at��9)������!��T�gv"��n/u���BCs�!�ݎ��X��H%/r@U�4"ԬH�!�D;x�]�$Đ�[��y���N�!�زU�Z�H��WRNr�I	͜#�!������K�ϒ�g *��N!�$D�vS.�@���g�q�/�!���.X`����ؘ8B�M�c�q�!�$O�O�D�'��h9>�F�"Xl!��Y,6ќ�A�%�8,6�Y
��^�"Q!�d̃t���`E�S�#w�)���S�K!�O�%z�����sb����	x!�G�C�M���ΝK�*��*��!򄐴t|
4�B�C#P�P�p�[!2�!�N�*��y�F��Z��}yrH�L<!�� ����1tv����f6�х"O����
u�Y�ƅ$l���cF"Od�S+��@(�5��d�����s"O�pA0��'&a0D-c�2d�!"O.��@^�(�T�Shѵ8:`��v"O����<T��	æ��NW���D"O`B�Y,tؠD�ᢟ�U��a�"O��a'ƚ$T6�I��-j?�x�"O�ɣ����R�ⵁ>/pH �"O
�)�*3��Q��˔r�k�"O挻�3v�ȍC���Y�0r"OPd���F�'�s�*X�(���#"Oj�H��6����Q(�n��"O���tk�.cÀ0������K#"OX����Q�4y6��*^���p�"O
��BIh.�Q�dK�7��\rR"O����Mǀ)Q�_
B�\���"Ox��	.UH�U�L�$���2�"O,̠�$ԫ2�.0�A��9*�""O��{��E���H��Ɇ�r��ر�"Oh	�1�A�51�ș5�J���"O�����H>:�#�'�5w�͡ "Od�k��΍<����S%ō+>��б"O��X�!�&��1X��Dd(��b"O�U��a�`OH!�G�?Jћ&"O�Ÿw@��B0qaDa�.�^(�"Oh5"$DJ.V��	fφ?��H"O��⧭Y�;C��ʣM�-�4�"O!P���r7�br�+����r"ON�bV�DG5L��ě&e����*O2<���5� �`!��64d�X��'�褀�½e�*Ix�+K43;K�'B~�c�!۳m��]R���%�
�'gv���K�Ʈa���K��x�'�,��1(�����c,�}*���6T$봄��TK�AyS��67��ȓ?U�����V�>l����tx"�ȓ��$���7��!8G�F%*�4�ȓ?k�Zg��G����
�#�6q�ȓhԂ� ���K�d��Ƨќi�a��.�@�@� ��f����Z^yP���K�X�3��V��h�BD� ��|�ȓz6�`�3*G�ibf0��	��FT��'!J��#A�3bh1W+W%m���	�'.d����*6��Tbso���� ��'(J4��$N�Wgd��q��2�
�'�0�b�a�w8.�c�Ջxz
�
�'���A�G)xv��E*e�8��'��t�_�]1�H@�X�����'���82�4�Bi��T�x$3�'J��x��V�pN�  2.��kܖy�'b�-A��k#���A']fb����'S�u1A��)o�� �b�)'v�r�'  ���%6�����'���'R����6��Xq,�U����'��­59�tC��4Q� �H�'��p%#�"&@Q@�F�|.p���'s���ҡ�>#�h��G� ژXs�'l0����Ę8*�PS���0}�!��'��	�Q"īYNPKG��!�D*�'���)�Ų�RQ��Q�m7��
�'�t���\$h��1Z���S��Y�
�'�4y�Տ�9��A��^�N|	��'�μ��m�0=k��h�%�(?�y���� ,�Jj�&T�ȫ�'M�ZBF};�*O�y��nO)y^��3j�=@@l��'Z�a�%۔>��y���#p�%i�'���� �%	����!JϨb:�e��'+�H��.���2c�gû��Y��'�2@�Vb�<�����-�l�
�'j(�QE�&r�*p�J2V��ɨ
�'�~��cȚFM�	ŌR0 �&�:�')�t:g����rȺ��n�L�	�'R�{T!��/.�����_�f��P	�'���kE#[9���ǁ6b��8b�'
J$�����^h�� �R��}#
�'����T�L84��bq�Hr^��	�'r��Am��x�Q�SxP ��'Ј`��GI�|�9�S!ޞm�hs�'�5�S�ʝQT0�R�Y�7�@-3�'�ڵ�`oޚ,�܉ @_00�	i�'�4�2�M\�hr�YKD�Q# �
�'��G",�.ɩ��M�(�
�'` �1MѹQ�j��ē����
�'� ����;ϤٚRI�9w:��z
�',@]1 Z�!���� $ ��j�'�Jl���/Dv�!��ڄp�l͘	�'�X��"K+�.�׀�
}�|%��'P
<��iïG��z�N5q�JQ��'�u�����,/,���_@����'�2��L��>"Tj�eؽ��'I��6d���,�0�Ϣ�!�'���ȰK�,9,�-��I�d횹��'=@d�W��
%���Ԣ��D&�'�`�+aAC
=�0���J�|�Xy�'���1��@Z�HEBL�y'F�K�'b�*�*-(�F%)�_�y�q�
�'�8�ECסS�Z4 �w�((a�'R�¦@�)�ة�2�Fk����'�$q��[-..C�m�#0�ҁ��'�T��W! �,����_�";���'�n�;`DXY?V��g����(�'�
�X1� �q�y����I�'��rT삄3�n�ǫ@}adHB�'{z�*Co��(����zm��`�'�$=�G�E�'�J"��|�5�
�'����[�|�Ac�z�|�K
�'�<��KI J�1����)	霍B
�'=�5���ox�qJ���E�	�'j �*��ۿn��y�TH�+J��	�'ʊ�RR�	�<b6u!M�Jp	�'ؐ �&#_�J>Z�0e�$`�%��'1��f��y�|��Ԡ�+	T��:�'Ά���Ԏ9��d��!%��S�'%&4�dG:H��\j��2����'�Ą����1O�1�3�F6�9�'A��rE��4H����#\��Lx�'���A��d�����.�5�hQ�
�'����i'B��d��pM����'i a���N�V;��)5♔d�{�'{*=��M�n�X�k�aƟ\9�0��' zj��_�CV��	%����uY�'h�����=z�P�f�&U�J�@�'�а��	�h=Д!yT�u�	�'i�)EK�#Ic�L:�L֡Aݜ�	�'� qs�ӱ*��)#�A����	�'�T٩2퟿Y%�ZV� 2a�թ
�'�� �i��^��C,3���	��� �!8�C2cn���n�.7���"O��Cg�V��Ƞ�7��#�"O�%xs�>`�K�i�/��H�"O��W��hL�)�Ɔ��U23"O�+!�Y�kpq���!���S"O���c-����-�q`��D�B9��"O)�M?o�P�y3BϺc�x1��'�|���.2�Q׮�+m����'Uf� $�E#"f!�WNN�M�]{�'Ehq+ËK�FD�
�Ǔ�Ki��A�'�!��p��S3�tN\][�'G��`�K>n�p(2�f� 5"\��'t��YW7Є:���X��'�t�C�^��܌�>H�"*O����W�p�|cņ� $u@���'v"X�.�l�b�t�����m)�'	V(��S�,:���4$D�Y��Q�'g|	0L�L0AzdJИ~�&p�'����BC)9��ɡ�bĠp7D<��'��� �	�)}�	����=3�����'9�Uz�"׮[<����˃�*w�}�	�'m��2&
0$X�C�%��d��'����7㜑i����JH�"��<��'vԥ�e+I /Zv �4��&�Ay�'�Z�(�E��ذ����P��'�f��S�!�t0�d7�f�P�'l���CO%(���`C�F�9	�'߆t*�נX�~����&�Hq��'j�e�!&M�u$��y!AJ4qlް��'�(��&�3�<YA�'ؕ7�F�z�'���A��]ɅkX�D�\�8
�'/�t����@w
����7n��$�	�'a�ɦ��
:��D��By$ "�'B� ��$��+���X��Ր
�'�x��JJ��dW���
�'����ȒJ��%
��9_��L�	�'�Ҝj0��.{���!G>R�THA	�'�E�Q��z ,ї�]P2��K�'�&��cR�_���v(E�[R.���'�$������T�x��FV�<d �'F^��e�x�@AkG8WK1
�'��y��B,x�d���?W�.4Q�'�A��C'M�
�qCѐBM�)3�'EHٙ�X�U�>�Aq�=��]��'n�aP4��!(B��#��2.��@�
�'�� �@!��0N��ɣÇ'�0�
�'ߤ�z��2�r���!W�%��)	�'4\�0Ea�)W�%bn�-h�1�'�rx)��BIڐ@AAز%�rQ�
�'q6���R�v�Ȥ!�`_�3D��
�'ل��IؠvĨL� ��+HPS�' X��Q�eH�7M�0G����"O���T�/t�X��C��g�$��"O`�$A-� m����� ai"O�`���ǜ@�l�� &�'!�Ѥ"O�� �
�1r�*I��$[�!��rg"O(թj��Qh��փ�Wh*��C"Otı5���E��`������r�"O���7*8�N�Jg��	sǸ]a�"O ��CFy�L�5�;��hs"O�TC �׿Q��-9�&��L�H\��"O���ALLL��!wEZ*ǤP�%"O8ݪ�C�1:\S�DQ�
I�hJ�"O�4�g�
$,�> a�\�uE�l�q"O� ����Y�k�pe �D�'m=���"O��L[�8l�R���Ǩ�˧"OT�P�b�@`U3���f�� � "On�Q��O�]���x�`�>d���"O(�a�C3�8 �S��3 l�Z3V��E{��I��V�ڄIƂ�5��8�F$C!��W6E�)��e�9��}����t*!�D�=`h͸D�M|-�Ũ]�4!�A�Bt�� �N�~1�b&��!5�!�8/��4`��0vҢ��2n!�ԋ5Vh������"�]B��Dg!�ę
�t��0m_�xkP|�M��c!�$V�L�^,�ro�M4	
ի�I[!�d�r^���o[,1%x�ʆ>W��`؟��0a��?�h���'�<{Z	�Ce��G{��I���^X$A��؀���X"*�܄�-�\��х~R���*ùE�Ƥ�ȓ_�ّP�E=N�
`@3��*_�*M�ȓwW�H�w�]��R���ݨt	����HO$	L��'�fو���r�z�sw�1r�1�'��� �͎W�X�Y'�K�gΤA{
�'8q{�a����t�eGҺ[K�U
�'� �� � [�Ĝ�E���T��a@�-��OX��˦o_�xӒ���k>��H"E!}b�Rb�(Z�ǆ:[���ʧD��'H�#U!�O���McP�[�D��RE0q���"���<������*�ɀ�̉Qg6�#a���Z�p9Ju�I�<����O���!p/P�gǜA@�w�"@2/O�m��O,O�g~B�!|@�"2��e������������\�W�{��Ӱh�r8 GR�o�+Х%~�JC�IP��Qk+�G�H��99� O��	O��0*4K�
l��O[�?K�) 'A0����6/�h�K�͏�o$H�i�旛�l� �W�'�Ĉ��U\^z���`��P�&oX�<Dy�B%�`�S�GRd�.����ְ�?i�
Vo��LP$֚$dpTp2���u| ��>)��&�S�$�x�G��>!@1a�^VpY�@���~�,ғ�HO��x��ӗ1
�8�[e݊AB"O@�a�J�zA[	��M9,#cO~�����g�@""D�*�R���8��'*�|BN�i�R�� ��.���N�yB��;+Z�I�D�->�ne��%U�yB	�����k�KK/G|:a�mT-��O��~��឵�R��u$E6��b�M�<�t�ٵz����M �,�2uh�r�<�Cgϡ :����%sʵ�0h�p�&�d��hQ�Wd��щ�2rݾE���8LO"�d?�$J1`�)1Տ�$0�Pb�ƽ/����D{��H}��kA��lz7�@�'YZ�"O$���-�Q�T�cj��1��[��	w�OS`<��hՇA��Tcvp*�'a�1��a�����J�5���'`�Ç�n����N��c,��P�'N��G��@"64��.ϋ&�.eHZ�0=Q��䌖_�����L�2L�PS�ÎK[!�d��Z��5X�MM.I�<���lZ1O`0Fz��d.[�wbH�TCJ1
9�h��oϚ��>��O�p�u�]p^�BA ،0�q� \O@v!��.�L{5�\��X��"O�Т�@�\�bS� �Z(�u��"OL�x䅂�{P�`���ӳ|�,$�D<|O�h�f��p%8Wo�*$�`��"O�1BI�0\�Y!��"�(�
�"O��'��=����(|�r�:�"O� �����O�?�0����2��HF�IVx���w��G ��1gCCe�f���f�ԣ=E�ܴH�.Ձ!ҍhf$�u�,['
l�ȓw���`���`�Z�s�
��cM>��\�����U�B��ˡ�T$s�>�����0A���(ɫ��,5B���hO?Q�p���E���x�O�J���t�"��V���O6��k.8�\�Sc�ì�@�'?�u��/I�̲��ۗK��H��'���se�ߺ^"�9i%B0H��<��'���`4�!���+L�vX �Dѯ��>�OdX�Ղ�uX��V(�1'vW�y�b�=�x}�� 00��H@�9՘'�ў�'�|rR/8u��� %�)nƸ1�!�2lO➸ѥC��L�!��K/u}~��/2D��Z� �N�`qJ� �)�\I�D�0��p<����<!�>���A,y# �"�EY`�<�P*\�\`�	���A&;|���c�_��Y�ў�'��@�Ŝ%�����8��
�'����ޏ2ܦ	)��Ɣ�*#�2OR������� �EÔr����\����
�'/�`��%�8KL�s��B/Rb"���l͠!1�D��Y�I,&��Pn���'��>��[�����k�x��г���U$C�ɫE���)�>r����i��5�B�I�[xɁ�ʁ�Itxl�6���Y2�B䉲 h�]��L�<42m�'V�9��B�	�;t����kˎ /��aEɕ�[�Pc��G{J|bA�BJ���I�ݘ{��k�e�<!��9FՐ9#%�[�3�����_�(OzuE��O�Q䧇J��� ���+ P�)"O��r�*V,3�v�8�H�R�Z���i�(#<�-O��?A2w�[hN<�a��"��Q;@)|O��%��ƥ��n8:��ƈM$U�y��%D��z�59�ąb�.O��`b+%�O����O�8s�g���e��&�Seq�F"O�9r�n�"/�D k+� ~I��)�"O��%i�"(�Q��R�o/�l��"Ǒ����?�"3�ْ d8���O��b>�C�d/ICąh���ݼ�a�M)D� � kB�J(Ƞ�w/S�r��DB��4�3�S�'=�&б�N�N�z����Rf�2U���P�'�� �dH6p�x�
��(`\}��'��$�6O�f��̱g�}!�'}@����_-n�h�#�n�& f2��'�
5�C@9N/Z����	0�6x �'`� �[�d(���+E�-��'^�Ɋ��H�9����ڮ$�(��
�'!�I���
�|�4�C���������*��XND�A'��1����'/C!�͇ȓ8/^U��Ъd������*����	4�pp�O�=Q��)b@�L����q��
!G!�}%�§nм�'��}�-��,���{��x����y�DF�zZ��ÏB�J��:����y"�4�^�!�e��C�[���'�S�OB�z��X�5��*��8m�����'�:5
d.!"]~��gkӑ<�ȁ(	�'��0�@E�d���cD�ϱ*J\��~��V�vYpG��B����b�]�y�iB8Hx��-]�'�T<�Q��y��'kR�Y"���)1��	��!�yrh�z��8�A(B�_�
�q璊�y�Ά8~uL0�gCT*]` �[�F��y
� P���p�<S�)	�#�x+'��C���Iǘ.�� ��úsw( rկR�g~!�䐃�\�ڠ��?9s���d	�$*j!�dӣ\�ʤ���PC��aw�3e!�M�g\�و Mq�|!C��%2!�$�����qp�ƛ_uF��7�V5B�!�$%��9�`�� [�\����'�!���(�����$�*<'*E�����nF!�DT�i��P� 9r{�a�A!�D�;Y�P�+�e�~U)�o��k"!�:QW�}�s&�Ua:\��m�	!�$�8�p���L2WD��Ì�#q�!� ��,��aA�$5���
��!�K�Mw^@	œ�k������_�=!�dN���D�FC�.$��@h�Ï6�!���xϪ����	�z�@Hă�[�!�����&���`aBN�NQ!�$��`����'�6�*�'ڀ.F!�D6o��ܱ��بb�(M�ɚ,?!�DI�/ꨠjsDL1�8�#��Ճc�!�^9p��ԭ�7����G��%�!�D��:J��A'c�:Xâ �E��fR!�d�D�l�����a��M�&��eF!�K>��IS�.@�t�ma�$�t�!���M��c/�\Zx�ǃ��g�!��L�8�
t�;OY�H)�ޕ2�!�X4q�8I�G�0���+���!�N���qC��&`�JlypD��v!���f�b�%�.O�Zً��Ďnr!�d�4�\#5i�
�%��8�RA!�'�P,�Y�腩�9u��RN�X�<��,z��"p�M�I�9�ʓM�<I�!ľ4}vM�� �N�x�m�<)f� C�&H� mŹꈑ�w��a�<���X|t╩ߴVJ�x�Bh�R�<	&�U?:�R��C�!|Ш��SD�<�sCM.�q�'d� lZ���C̓c�P"0fU 88�(���۴~]�}�<��lQ�g}�Ha�ͽa���S�W�<�Lݛi����!I�Td!���<ybjScz:%�����Y���ʰ�@]�<	E��
lm
����13�)�we�l�<ц�Y�b]�c#��G�1"��s�<���A�$�p� �D��xL���t�<�vg�#�Ќ��g[�L���PFv�<� b$P�ء��L~�ș#ex�<䯘�>�ޙ@TkߙSJ����{�<�D�4�-Y�N�8}��� NIL�<9�"�<S��x�!�Px�¬�`�w�<�À 4r�`5S�,8�㨒U�<9h�I6��9���wNa�E�R�<qա�8 ���F��=h 	���@v�<��E���r�)�➶�B�(�s�<��a˼n(�$H"�ӷU��ɢ�
n�<a��l��<1�"��#��y��d�<p(�\P��\�l���e�b�<��`�2|tRi��d��ui���FB�<�1��g`TXdL"k��@�E�U�<���,n��У��}P�����Ry�<�3��>.�#R�S�)�Lh������_�"$qO?�R&�9_�J�0�&�� �`���s�<�c�;/{��J�#H�\8�H�r?�3'�Bd�P��"LO�=f�@�E��iZ���'1�DS�B�,�#�I�zS)��n]�o��q��5���B�F��	��44�
�h7�[-aV�O�q�el�{���qSB���π ���Ly��) �ļ��u��"O:�q@���p���7d�R�"�S1 ]��J�Y:t��h��ת#(V�Y�%л~fi�F�ܓQ�!�D��a��ȳ���pPRuc�#Z�D��b~�Q�N�j�rT[��'L�<`�%K�$"Z�JWo��X�H��čw_��C�{J?�R��R�x�g��uwb-���hy^��V�[��j!�'GV2x���`[�kL����	�`b:0�ݚ�?���.�F�&Q!ԍ�'��mE��آ�Yd�~r�ۦ8�̹��-��]b&eOx؞���U1Iɮ�)��W�M>�٨� �c��D�*v8`�x���,,Q6 ЊKQ�J�#�v>�ٰ��b�)�*w;`�l���Z7�L�G��c��*�ʅ����Օs���RT T;;`D4�� ��3^Y9wn\�|��fةM7��	�=�p5R�`�8i���Zt���!v
����O��Yw�P�;�dj��;l������>?R�D�U*N��A��/K���s#�C�T��D`^=�𒤘(�u�Fp�\m
p/��b@9�� �#���'p������Pp<!�gѽD�H-prG^�隬�Q�ǒ#|�cD.��%s���{"c�iը ��Wqn�����'04\m�v�n�nIq�H�+9�@r�c���Q	r��D_�U8��S�1��hP�c�GN��qP-*sLO�@bv��0s� ��<FZ1w�4�y�E��6��h�F�
;��7�I9����"�ڠk��}������N<(0�)� ��?��D��Yt�E�1х1~@��A��Opl;�g�����
��-�	;���ZoL�9 y�TGF0 p�{p�H)3�Ԉ�#ᓗ
�f�,�`бM��t�����ޔ�r��a�M�־AJw�A�	��M� ����x���Z�p��� �_��x6�JF�	�AC��$pT���"¬ְ0)��23N{�gԺ?%>��AM
�G���Õ�"|L���"B,Լ4�b$_4.0�إA�.w�dS(*@�Y��B�]���g��%F&�⒄^7+>��5L����<����3c�	
���u��/�lI�S�=1ι��O��V�����V�>��ٸCȺ��"�s�*D�E�O<�!��G��2��i��Κ���{����}|tpr�O�5>���Q�:�d�<��Q�*�����'t�Z�s�鐢@������Q�RQ'���
)z��N�8YeȔw�^�c�)"G���K�$T�L9��0������%Q,�� �*� Hݔ�O�� �ʑ�L׀ ���ދ��qBu�
�F�)��-	0�z����H��};w`<|�0	`�� )���H�q ���'�T�'�INuzԭ�����+T鑃~?�p�G�L���e�Wa^΀�#-%$�~���_�li(f�M<��q2R�8N���ݱ_�Yq�&�7p��@��Ry��q3F��1|�r�h -��<�`�w-��biV�-ޔ��S��~��Ys6F��x�d�$� 0�& Y����O� �Z�ڰ��d��%N�(~�:$HPNԫjN4PP�A]�����B �@���O�`!��6aP�YA�|D!*6!�$�L[���4��g�1�	���c"�P�e��h�B�$��Xk�*]O*��q���6)<q��44���e$Í�~tyc�iO$q��&6��H�Q�ݏ)mK� vV1R�C�V���mA=97����2�}x��2J��H�DQA�O[�~ud��'��vlY��P�R�D��T��)p\<2p&Ɨt=�eoĺOR<��� i|6�ǢY��� 7	K�U��(��M,�tLhr�V�}QB�ꜫKEذ)U쑄'b`��GaФ�ډҤ$�W�YpR�=�uWi�p�<=9��3B���� -FP��&��uQ��Q���9�6=��6	V�����@�1�	�'��qS������Y*n�0&�O,q+�jƊ&Q����׋a��h�b��@�~�B%[�\ |�`��N-EK*Ɗ'T�����H�6E���T�v�
D&"�� J�5hT���! �n�0Qt�|2,��o�8ATbҫ��|��鈒#$F�[�<ۥj
!
:��iH�"%F�p��M3\�ЌH2@�Y��Q��u݁1���4 ��4"��&Dv����$#VpA%LA��"<bT�p�d��I`�莎a��Đ�d�+��`��D���8�K2��`��/�f�r�j��_?:�tAS�̅���q�O+[��{���֦�����?���r� �>|'d��R�t`������	H��/Ժ�,�iW�	Z)ޘc�@D/$�P���ph����b8J����� 7�ʑiQ)ڽ\Fy�q��^���k\���ŋ1%���e��I�4�ޡ��۾THm�)O��b�Eř'�����
=M*q�c�%\T�A���PB�賄R�b?�H�����#�o��r�l��̆�L2��B��b��L8�Å%N;dk��YQs��2��͆4Fl�2Eޚ=�'\�(�)X�e[���5��_2��ԣA-��q!��qFC���5S�M��bq�"8h*ĳ,^�4�����mv/��������9#��\/x�
a�
-p
�܃#kJ�S�\��'Wl�{��_\Y���eBޯ�\� W�ָN������*X%��BqÝ� �X�;�
@/sk�|�%e;ΉYD81��n����� gӐ�[1n����a�s�h�&� r�)=@���ab�?t�n�&ߣwذԒs$Ɋ'��K�N�n0�=J��,8H���A��ԡ��h[����RJ�	�L5qV�Km�4��4k�Y���'��|�vSH�d�l�"r�*b�Q�-�j�RE�H 6�Ot�p ��j9��@e�]�d�(m�D�	`�lڗ�j���L��)�������zh��jF��|�r��f ~��SŘ��Jc�˹��I{6`�
=R�e��)1[�I /�hYV�C%�@��E sОQK�J���!hMU�ֵ��m��}���к��8	U*]�;�9q�q�|b磑�&�D�ϓ! l!*�L�g�n��a@��V�%a\x~��5d����;v閴q��W�?pc��:�>�c��'� �H1�H'<p�(B�ѻ3z�c�i.��'�"F�,RG�t�̐M�0��#�uǃ��rp����)[��谆��`h�@f�Ͽ=&���5�I�i�>����b��o��T��$Ccc�<@v��9(��g�&?8x�ր�"=�P��qT<i
ٴ.�Z��^�C�`��M#zx��|��&OeD1g�ܛJ<��-�d��u��s�¹�d��{����Bnר^hFY�]�O.=��l,�n���s]��J�D+@,)`O�1
;L�pBeZ+N��Ez�N�#�����L,�����8Yt͎�"ԙW���'�I IH�B��l1��ß|�(1P�@_&��!�M�*�����O�i��$MR�G�ǘ-�B��ѫ��U�(!��>���WU��qJ�T(Y���O9~7���NK���\9�u�N�c%
��O|\��M��~�N�6BP�<��@��%;�U���՞e.���nϕ~��![V��xU ކWW�p��,B�T�r�eOU�epe%�'�yRm�#_^��@5�UP�X�#�àP�h �Uŏ	(��0�g�A�N]�\Q��@�bWt����#z� �T�ɖ3�Tz��G�)����f�
� S�T�{��D���҄)`H����с1�D�w�~16q��F��SMԏx��n^O��i��9H�9�cY�/q��{C$��}�����Y��O�t���#R��w��� �%��#��bH �`�);:6�a�K�n3��zF���M+�G'8�n�S���[�.� �ЋQtp`����>&�~���/hv�;c�<�Z��`�5�	�=��zu!�\��N#&z����Z�V���,N"�$��"�֟|
i�U�\&��(����;/�h�� �P�[p�y�#�0����	x q�%g��\`s�
>K�@�茓k�
�����PRFBH7Do�|�$�M�I�,�)R%ߥd!�d#&i���wiф4A�����",�h0 �8��9(fBb*��B���c�a�(����dL0�L(�j��r����s�D�$c�Od��1(Z#b�tXK����N4�T7j��fM5u��L�t�PD�l�e�PRH�ࣃ���`���P؞pH�`\��f!���[�Ёu�@ry��IG�L���E�Ϝ[��IT�V�p�a~�
�C�x'�C�-?4� �I½U��CP�H�,���fӇ��F|R�
�w ~0�@E�"}h�x��i��֥�){�j�&N	d���5A�LI��wI�>Q�-�-��U*�T<O�z@3����t���Ҁ���xQf��<v�`S�,C�$Ƒ{�d{���3�4p�(�"�";tI��lZ��E�i�E��@Ĺs�xq�m������>E�k(�,2<h!S6�ک<4\��5�Q��Bˌ�Z�ayr憙�+F�l��$�1!B)�3Ƹhǎ�1e�-7n\����bl���̙�V��z��F��"���߆Li��VP,�t��E��|�6��d��Q��騆��>Nc��86㞲L�X!P �L�B��Ć�c5�	�4�� �X�$�U=Ii��Þ2L�R9�NHJ�V���FC�1�T[��دI�� �2}w�lrFWg�9�����B���#kj}�a��`u���~��㵯��0%�6:�I��`I;X��P����nm�?ArA\�HZD�  ���W
��X��Ky?����s���/F%\�7�9J]T�@���Q ��`�d8'Ա�&U�G�b��ea-:V� �@��:kD�)�/W�Y ٪ߓ|>
�
㬁�gPT�G�77�������=���
(R����Vd�p pE�=ƶ�"�.�nl���w��xر⃎S�n}����eW�}I�/˄����4ڶ R��<�f�1$�B�{�lm0CJ#'������C�(���W�7߰,R��<�l6j5�h���5!�04�$X��N�S�LE���O�4R#���(��tӲ��v�UX8��t�w�~�IB�A-e�*|�E�M��T /�'��rJ�\2��	s�t�iN�,f��I!$�J�p#"�7J��x%&?��'����*��8�9���	jH��ؙ��,��A�CK���aNM#:�^�IU�\��f��H��� �shEUw����FL���1�-�*Q�[� �I��h��e�����BeH0R-���>Vp��@޼.W�K�`UK��x��%����B�������&ܬ8�C���a1��/؈xo�Ɇ�	�a �L����G0HR��m���-��ybD��$%�����]ڦP����@(db�(n��9ȵm����(	$LL3C"���J[�Q��ہ�'�
���/)i�V=8F��9HS�г4�49g/�#Q#��K���g��ϓs�Lb�b���\h��ix�Q.ޫE�@H���
��J���,ªE�90��S�K&���Ջvn<���H�V]��՘D@P�A��zz�Q��J��9�����)x�ɰ�֞y�P�2*��]|���Q�~�ɧ�D�*�����'�z!�%z䩋�������;�t�����C���1�K�[�δ��+G+�B�iK?�����L:�j�����&�Z�ŝ�lN�FE5A��T��A_�����:����T�-�Nti�����A�M�HmӲ˄צ�:49~'F���تk^t�ТLB�B.��7�D;�����*ňvX5"5�ar�I��0<a�`ʩb�� ��J�N�s��/<Z!�Đ��c �X�0�N�Ӣ���+T$Ѩ���uSi��/?����4#��ٵ5�\����@,�X��gZ	���f4�L�'�"�*TȆo�r,ɖh���߄�`ڴ|Lx��� )V�aɵ��2�v���n��j�L-�2�^].����n�DI����B�'�n�ې�H8	�� c��Oi|���s�?	������'.�6���:}l��!u��Yf�Ğ:���S�ׯ�; "�P�H!�ǘ�a�6)��EN3(��!�*|O�<S��@61���J�.��)k1���xB`č*u/��2`�ޱ�
��wD�44�ؘB�"�-��9s�zD D[Ӭ��D>l�R,cdN)��]�{m�x2$J,[���y%��1ta�9��imj�Hu�H�64�͕�O:vD{AƋW"�����R/�F��4�6ln�`�	�
< =ɒ�TI7lh+�'�Y����x�|��F��9?�,Y��I�����/j���˃)��M۱�˺��k��(��\���C�l�h�P�KϟQL��3r�X�v��Qb���A���)��8#ƌIJ�k^�de�$��R����0�L,}���	a��m���g����'
;_�6(X�Q��г���w������	c��q0�(&N�nk�@��R1�L�3�Яc�@m����0��<��X ]�>���wz<K��X���^-Z2��a�3u"V���)_8Zl����e�ޒ�c�;�|��/2���&�yb��pY ���9yDMPc����'k�c ��2,��@�'9v��� �� _N�2�`��'ˠ���$	�:���(�ƍ�6�5j�L��I�̯�|!F�ISk��u��	4C֤P�93�l�;7L�	�i� �	��I.O�@%��n�5>4�ֈ��p�Ⱥ�O��8S#�&�o�N��/������϶C��0��$�O 
�@��]�LM�ϒR'�� Ӌ��E ����딧7��b�	0��f�~�b�)�ᦉ�D�?i�HЌ}
�!��"t@���#�а=Q���1znhZ��Т#��+|m:"��]Q��s��c�
����%%�*H�5��;� )��ΟXZ���_R�ɚW��%`�A���渓h�&X�Db����0`D�R'�@�z�Dh�c�"�zC1�,rDU#���S
�P"�'�1يӱ��`��T� Le8�Db�7/�b���:f�ĵi�M�ey8@�2�<H��{�\��u:>hK>YD���nٰsi\dßw0�C�F	u�*Y��lih<3�'��Q��k�J "7�ģfi�l��+�7(��8��E�v�R<FF�]��UÒh�n�P4J���!el�|�]cִ�Kƈ̮nb�\ �ɗ_�ވ�04lO<����Q7��:7��h�àF\-(H*8�f�^�ڽf��h����C2k�4م�\�k���F]/����  ���GQJ1��m�9(��i��ΊijJX�$�S�@8= � �[
輈�fE&J<,�)�E�^��a-�}�vu�IΪ&2Dȉ�aI��H�ߓ�btP&ˁ?VA��R�2���(`�ԃ�`��bI8��C	�hdHkA>	@u�`o�V�:����E�)����Q{��B0�
�ht�]�ȓ&Q���Y�~�Z!"H{sl�y� Rm�4���. �$��gǝ.U��)]�j���yqn��1IVb2�(]�n�L�a�g6?��" �'~�q�P-Zr�����t�A��X���C&d�es�J�f��Չ�	y7�Iv��?�I&�;��<`��K�I�>p
r+�VC�� "�ꈾ2Μ�ǎS�|�Ob��1#��?���R�(�,I�����9����s	٭q��݊�'��t٥�
�� {�K51Z�)�rH��__����̰F�i>m��N�4�
Q��MM�m���	%]*H@�r.� ��p�D�6'��B�I?��b�&"�|��%k	��I�4� �cU,ܵ���}2z����z��K)J�Ng�\ы���=@L�H�dmx��@�$�-ݛfA�1&U�@�+Q7T�0ƤKz � �5�~���{5*A�}&�й`E_$N`OS��r,��.$�\�-�8cp�ub֦�O͚x#D([k�*�VG&dnh��� `����Õ$����խ*����%�����U-��� �v:���`	0S�B��`���X�!�$�i?�X+��~t�D�_*k�qO8I2�o�5�0|�0�W��e�e��Y���2D�m�<�Ə%�T=�N^�Q�+��Nk�<ab-M�7��EZ&ۻ~d�����k�<I��"\m u9�-�4(�2) �d�<�&c��3$�0��$W�AVȴy�H	e�<ْ�J�X/t�B�,�|��D��f�<�ٲ`\���Ur��hS �K�<y�¡=��i�@]
�P����j�<a�CM�G��H�q+�=Lt� $Do�<A�Ӯ7�J�j�*�>8j�t0'�_�<����x5#� ,&�H�K�HDP�<YvhU��!+T�-0���QC�K�<��C�:jbi��/�Kl�t:7��X�<� ��aL\@�� �5��Ck�L�<��U+RN�X��P,<a(���*s�<�v��d���[�Tʀ�1F�m�<�ƌb��8�d�#����n�<��)�;:�X�kM 4 �Iҏd�<y`f�#}@TB$@��"�����e�<�(K*^��-RؗE���Sa�K�<a�׉�p( 5`�6�Q[���K�<AQH�+&��8�fZRp����R@�<�pm���q�H�� E�R��X�<Y�i�Ap�@��C�=%FX�p@s�<�eb\
;7:丁��9,;�9zD�d�<�V ��!�V-��oݓ,��X�#@�f�<���L���7�&6���]�<��:Q;�P)�ʛE�D�"���\�<QpM�>��b��|����Yq�<��n�#b��ebhE�}�^u�c`�t�<a�&�1����	;��a[� ]�<��R�oB�D��MX�ե<�`݅�
g@���dƋhr���*nR`��P+�˕�=J ]�'̕G��ȓ=��<���yN	���(p���4�T)��DZ4VXPH����DI�y��(���t*��c�Ǖh`����qi���9�,���S'����O5�d�q/�@���Y�ń�p~�%��%$j���%�7����	�++�ȇȓ2`r��#�1Z�9C�۸7U����l��iK�U}h�1N:(��ąȓ�ڜ��ɢm՚�H��מ`�pQ��5m���Wǅ�>>��)���q���I�~wX�����9<�4��t`�&"��Y�=hjԥ��S�? ��@�H�Z���%�ɏs�^�X��O����f��Oz��V��D��2N��d� �^�~X��IP�����cR*e�1���0 �~ b�U=x����Msh<�VB i�Tdj�#@�]j��Lk��U4��JeM������ '�Ӹ>��0�u �=[r�E��%p3�C�II�Tz7�P�b�
L���E��Y�T���s���* ��~��$ ��N,@�ŭ|}�ْ�9D��I�m]�B@���D�h�@= bCwӴ�K*3�ગM^�Bn��Q�̵���3�`x�u*� U�1ȡ�ܛi�qO��j`��j]"S���]�x�p��9ᰬ��-�%!���׿��?�&Y�?�hESL̽@������ٟ��햤1���4O�YJ����X,;�~U2[w���K?�8����2�X��e�,���e(lOb����VU��Q������ރzJKс�v�l��p��(���W��1�%@���� ��z�ġ�w�j7�aج����E: !��D_.{Wl3�{�oW�)��M܍F��,�!Iѧ'�tի�@{>� G��,��l�pCW%EF�VM��qt��r���9h��$Eo��\+7�'��D���� OV�&�5sp�iS)ǝ}��0��f��SGN)�JB�5�b����ʢ
j�`)Ed�S�(�Jci�ݺ���&]@y5$ը��p�;:�,C�%�$1%*|�b�Z	.B\�#oS35X@U3"�+���bAD%>�<!{ӥT�0! �(c�� �������l$��@2�pi �b>gf�< �C$�~��`Ժs�~0���Oi�zsˎQF����4Z�h�!�'Ю5�� ��0J�L�e��H�h���gv�rsk!0y�t°e�+A�`9� M?_YV8Z�7O؁z$*��}���%D����� V��y�s�.)!��#	ȕ1�����Wg�!�ɗ���'e�#�V%��pɑ��j 1�F�6�r�)H͠�X�!V�N�
h2�E<�Jl�L��`l��T��UU䄱�����`vaW�J�t
�E��9�PX�L[
b�iH��.HG�*�c֘<!4m�`/�B�`����!@8v����R��q`$��J@�4J$�כ9$8m��o�B��3dN�4�JyXdW�7�` �	L�2E��1�KU�A�f�!C�q��<r�d��7�XQ ��|�%�P��y��	9	~�c���[R.x!!E��#~���s V�1��1���C_��IZw �,���rb�I�1���j�:*��  Ǌ'J�(Ic�L�<�˂-�!t�p&�����%~�@�$�ӓ7� "�o��|���x�A͢TЈIu��U���7i�g�:���&�:d��:`�(9cь@�4�A#�ժC��c�`��	�jO�D6�A���I)��D4�U�0��+"�~HQ�
�#��8!���㒀jүF?(�R�+�8E�&հ�/B
;d�0�0��r��k;�&��3���	64�*W��:A�4��so��=i��#ҫG�L��s	׮P(G��>s3
�JT�U�?�h������v*�kף/C�@��c��dp �]���`�kP:V���g�rx��r�f�q��=��`A�v:dHw��g��y����\Љ�'��q~��"A�<�D�y�-�En
�~I�8�TKZV ���`]2[�8�g�ɑL��Ex� -}��UN�0~M�0ل��Dz@M�k�V����Вzn	���N���E�Vn�o�	��G�KqO�L�s+��#x���/��7~<��G�[1�}���� ��j���|`��P�.��|�P")�MK�/�m��@�C/Kd925&N�S��]���Y�2f��)'CQ1��\�2P�h�R���G
�no�@у.�8e5�&H���\kU�ت�☫��/ 9�T�ʹW���9i?D�Z�@P I��6�@�R9��Y�F�Y/"@��j���`P;>R|ճ�
/K_��
m�:���S%��h�d��Y�5�ȸ�@H���^5W>h}��,�mh�E`���v�"����G�6�����d�8��'0��q�-��Z��,���N�Y�p�"rcI�f��'��)7bP�`���\�2!�׀A�}�Ι���rA����	��7L]
DZ��S�6Z�2)���'�н���<,�R��'�&�M�7�L
i	t����z�RaRB�P4��z�ViBR��4zqȰ�`��v%(`�u��&`�j�"7���B�X	₆]�Yj��,sX��c����w!0T����ݪ]>�a`���>V� ���Q���aui�;�l �C5}ҪR�ct��`�Ǫ�%x�J75�<�&[,�v��q`´s�ZH��BĐb�T(���,Dp4|C�LD�i.@1��œ)LZ�R�cӚ��ƍ�	#���h%��Z��D�VΘ�S�ƬQV�x����ů9�%�d'd ��	�2%6HЂ�A��W�֌��q��Ȏ���'����ӤJ d�<c���C�|k����:O� 0afN3E��8TA�6%����Dn� K�Y�L*����~v�ӓ,�+g�8m�W�O����'=;Ɗ�R�J��zA��j�A-|r���,Y��T����^&~9��/��-��h����5�(�0��GJ:b��"�I�m��2��7�p8�,O��z(L�K2̔��d�Y�k	�� �d9�Y�3F�"q�*�[A rE0�A�]�=cZRW�ӽ�(WD�6�i�#��v�>�1���V��� �
�!w��{�ޗlN��a�O� ��ܩ��L;"�Ϊp�J�c%J:�ġ2��
�!��zw�[����@�
S�Pȹ3�8R̘)����-,�8ݴ9t�9�����jS+�*��N��F+��.�|9r�,\�Q��I�)W���R���3��Q:���a���U(O,�b,�%S���ݨl�H���w��$+B�͏If�p�� N�D�@�2)�2"���H��lya�H4,��42�̍Mn�l��@�<����<|`�`�7#�D�fA�4q���? ypBĦ��C�&Nr�8�@��#	gR��PM�>hq���nL�3��8���3��J��֬F�8�f����O�?��%�T�H��Π:�bG$�a�!�1-�!
̬�J\0��𲕠(�	��(5��%c�Mͭ^`��� ΢7�;g	���ū��<t��\B���uK	
�Y��P���'� H3d��"򺐣U��=�(h�Ӂ6N�B��9Z�=-	}9��W*[I�8^����#.EP��r�ˢK����;O8��.,P�8�\wo��"7瞗"xLpI�B[*�X��cJM�t7vXJRgE!���ɕ:��p �#�妥�R�OP����̅t6ll
��Ce��a�M�7n�n��fJ��y�6�)tfڝ�M��M^x�\�Ѱ�P'��Ӣ�n��'��X���W�yNHJtX+~q�e
p�޹?�d�:�'ĤG6����X'����c�*vPp�#Y)}t�e0�8:�~�:��G2��yP��ްr�>�h�8�n8�W	�G�'�8��oY;F�B���B�y5��K���9����H�bAx�[�	1@�z��C+Ίy��H{��8-�<c��W�>�����H5eKj��	��Ń 36�"l	�h��#��#­]&?��K@I'd[�Hv1X������!dӆP#7������r���\�y�`H��F�u��"%}&-��KQ��
�1�R$��$�Y�M�����@���M� �l�po��YƧ\
�<�(3�
�	��5q���e~��3�L���k��aF�]� �P������|��u|��x�c�;V>B��M��?I��Ɉ33^�5�����3�/Q���ECUe�`oмm8,�e )N]0��a�'
�݃f�B!,^���EÉPi�@/��my0 ���A+J�P(�#�-$(��
nS��RL��c:T�F~R�%Y�V|�b�c&	�4e�lJш��՟��02nS�J\zЋ&�IMP��A���"�8	��G<hC��d����SNVl�Ӏ���M:���Y�<h���d�]V����۲!ףn%�l(-I26}ִ�a��;-t=�F ��pP�ܠ�d��"�Ą�%D�i
�#�e�+Hp�B��	LUF ��>sX���D�-!�̌謟���@� ��ѢU2!��mB�K$�~"�ޏ��)�oһ^�&Y�B�O?���x���M7K�%i[
��7*�4`��=�ƥ�5,Ԉ�7Y�6���/��!!F�"ϴٖ�(O�*�e���#��E)u���������:a^V�"��+���J��MK��V��kS%�9X%jVnƁ(m�a�`2����%�#d�`�
ۓ{���;l�viY�X	�-���E<q+w��&7����iІx��¦l��(��4c#hh�� �<'&ѧSV�QA�"���'�܌I��G|R*��0�6�����2}�J���i���jL�j(��3"��O�QKd*�7G�m����8!tl6�4X[D
(}2��-��N~BC�ד$uI��mV��R� ����<Yb'P��~�P�D�S۴&J�nڴ]�
�{1�@.������e��E2���o�:x3DM����o�>p#Tm+,O�����%��M����|��<P�,�	Zs�R��\��m�w��c�
���O����,¼NE#�w�VlZ-=B���
!�@�����GY��$"�\∲��P	:H��S�)N���e`N�=���3�D/?�J��d(ڳZ�����I�'��H��烧�� !�(�K���э��+��\���� LQbR�*���F��/���I����c��5`�t���i�=n�����lON��%o��:��P��LB�r�{FK���)�G҇c�Hp�#ݲ[���89��`� �C�b�S��?=��F)P�|�b�֚ �T�1D�q��������=N���X�O�ú6�X�}�t�G�����i��ؗ���Kx���Y��M߼˅I�0�D��G�]<',8	(qo�[؟(c��IN�iY�H�˷ub��gIE*�Qk��
u��xCw�|�B��2�ѷ��X7�˷��'��읒 �~�{ҡ�3�����DΰvI�H�1�ɇ�66���Rv��%or`���l�;gH4`u �[�����G�:�jX�C��W�<w�٨B���l�0dF8ɖ�^�#�D��1��=jE���GAۼb@�	���	$�"����+x��$��Li�C5&8���¤O*|g~�x �����?���ѱC�Q�3��s�U�"��8���N� vЖ��Θ.SZ����"O��4���p�]�ʟ֡	��Z������B#r�l����*8������$ ǎV`8���$�6��nS�y=�|����.,�9�nS�m�8���Η^<��
`��&�4���|;�d���O�8����=`2��"Ɦ����W �`��ɦ>PH��!Q�Rp�I��4�9��+R�mn��0
U�*���A�'"*�0-��&��
�LQ�"�˞G{�%nZ�$��8P��+/Vtm�(����ā�[�
$�F+C�B��s�-?A�͡U��2aǕ�w��0�dK��&��Z�P*t^�q�Oɂ*����d�ڍPX�����2�R+؈OD��`1%�50��@�m�(������d�Q4�GJ�1O����A�mO��Ae@�?y�f��ěZ:���$X�U:�7�0J�����<jC��I% 	�>��W#7��S�AܣI����.�6���Ĉ�9��B�R��`���اV���PX�/B,�iP�i�0�TJC�|�){ ŉ$?⩑6�3L�<��a2U����T�rГs��
�ҨYE�8O����+�d(7F� ��dǃep��p�Q5B�q'��H�|$PV�0��! ��v",4�lgw��(�+�?R�9�"L�r�D�u�B\�V�D�F-@�e�ް�I	[�T���k>g&Ȼ���H�$�}�B6-W8WjP���  |+��(��=9�^�3���	wڧBݍdr�ˣ�D�f x�`�I	4@4����+#F.��Պ9G���d��L���	�!��W e�@p�BH�QK�tPիUw�b%&	<W¬�f)L�[�f�Ck�G�����(n��<�ߓ9_ؘr�
=�˃(!k��d�]o��7��d�X�j2���-A�9��&�"xZ�)��U�'g��$��\j�$���@�T�.���N�i������ؐF����;3:�]�R�O�aE��3
uӰ�R�O�t�^(�um�x�F+ˮ(�����I���LE*��5n����ˉ�
��%+�%qg�LÖKJ�<����=I:��U�#5?윻S�ǟ�ҳ��^��<r�88�Ll�ҭ�(<K8��!;������O#�DSъ�fZT����:KLLI�nJV$36��X[��됤�v�d Ų�O��1˩���9�]1l���9""� 4���1�\<��+�" � �a�+���iP��0o���b�M�0��*�_Q���`a�XQ��D�G�.#����剱=�bѡ�/B�5&G ]�d�RȰ}oแdϏ�HS|*�5,{���_�J����E�  [�@��G��~i赑\w{&��7j��QƋOL�Đ%���b�d��l���Q��3�$���#2@ܝ��������Bd�K�d��PYAL�>�n��$ƿ&N�,B��J��u��f�~���N����w [9�DuKFǈE%. ٴ��>��[�i�4c�l�(��C�|�g@�9��tOǟ4��g�%
�aqǤ�C�*�a��~7�~��2XC@����[��]e/Oň	���K�P��^4R� <�\w�f9�g�;R|7�)y`��,y��8{ �Zh������8Q=؉��	�y7zQS���T�>MA&鞔z�C㉄pv�H�a$��y��Q��Lݺ2�P,@Ǉ��D�D�w��y���$�u~�\��OXm��f9B)N}�-B+t �[��D݈��;e�X����D��Ƶ(�8R���٦�׻:�j��6꞊BA�u��:l.p��#
h����$GV&�xA���5X��Q[q�Ծ"xh �bΔs�uõ�5�^ɯp5,�zqK�tȤ��%lZi������ ����3q���d	��-�"O�ds�/׋l�e�'���W��YH�K�R�l�p�F]�x��Lx�j\�b��t{���f�Q���
�S��Uh���X�+'�Ŕ9���T�ɽk���f�p؞<�烍8f��0s��	*
Jͩ%�O�S�n�0r
5 - ��U�U�\��i��׎ ��@+��\L��EhO�W��O�k�e��9��̭8�vL"F�d�>���
D�Hp(����1����AIX(G�Pd�'�Z�����K�;�&%���-4w�m����޵��1b� ���Z1t�=��˝?��:C�M�<�9׮[�N2���C�˭3g���a�0p�	�ăJ�;�����Y����₰�6����ܬ_pE�ȓ.I�j�m_��t�e���'B0t��Q(%��MX��YL#Ҥ��*N�Z_���\�� ��%@2p��E�\)�4hDb��eX�_��ɪ��']�Uȕ,���L5�tE�<]�<U��G\:3R��)@�
�V�8����\}ĭ;3% ��x0,�?Q��<��-tк� L 
c����*Ǥ	.���A��X�i2�X ǉO��U�v�*�J�D O9�B�yR/�%�X���L��+��'�H���*͏A�8��$7�y86�Ĺ	����G�J3	J�i>�Z�C�,�4�PŅo���ɘPD*���I��R��D�t��C�g��!B ��zD�X��+���P�I���#�g�X��|(���r���ޑ>�.��ϟbA�2��dQt8Q�@D1'��m�r�'��e�RV�8�OV�J(%2b���h|�)���0�n���Ⱏ@�́�v�q��'g��Q*O�ܬР�H�,c�a��'�b��ℓ<-��id� (Ѥ��p�:*K2�ˁ�ߟG�|��/�~XHY�$<����tf,��Ŧz�"0��>���&(��#@	�И��@�'�!�N�NWٖ�rƔsAqO��!#�9�0|�K��OI*m1����DS���`g�<��aώ�T#��ڸHi�=QQ��g�<�%C�
D�����G �l�1$�0D�t�U
(TH����Ƅ׬,R��(D�����	S�D�1c��Q.M��yB(�c���`	L�~�n�&�!�Z�v����>D�8�h�@�cH!�D���ڂ�>>aD���@�\!��� ,A�n_�$���m[#�!�䀻j�~=ɂK�.�����L�D�!�d���PL��.�o�.9"�ʟ+[�!���9D�u:�GR�$-p���0O!�˗CW(�:B��*�����I�k!��2q{v�ɑ�Z�d�3H�+&!�D5T�j��%k�R��ذEN!�""�n�x��S�,��&�q!�$�9l�����{7&���K�,0!�R#8æ}J�aŵ@,\��4���!�P:Z>Yf-V9?;X�b��I�!�D��mĢ um�I�L��#�9�!�!-ĘXĥh.x�C�$\!�D��:@pp�Z�.V�-�y��yB����E�Ԫ�/&	�͝��'�P9���EHI򷥌��T�j۴�tI�(ɠI����ȟ�L)t�J 	�����
(A� C�ύBF� ��kN~�,?��-H���V���,>z+�tb�躟���LT��M�����a���~�P[��%V�Tt��M.��$��<�`/;��S-w����רK��#'ڟrO� �����Z�jsb#tmѫQ4`Q
��T�$��I!k�Q�"}j�B�`��:WN�7>�$�t"�ҦE ���a�e�<��P����3V�X7���x�����N3q��L>�� lQ�F�������'F��=��C���'��9���#���0Q�(��Ͽy�tp[Q�x"�K^?QAN�`�O�왨�e\$�Z����:;n���O �(��T���y����'B�t
e�P���@gO2^l"�n�N���j���S�O�vI���� �p�0`N�J� ��Nה+��c���ç*,��E!S7����,Z� I����� H����	H
,M �l��P;�B�S��O�թf�Ţz�1O��i��W6r�*�E)���[US�����y�S�O�8T�5E`0Qd�Yaٴg�H���T>��'WZ��Zw.-����^���i��&�|��"/�j�L5J���O�>@ЀŖ+Zt�U���(e�� �C�Yn��	��B�*@�?����� >T���+g��J�G�$ 8��_�<+�Nh?!	H<E��C��P���!�&a���J��U�M�#�]�2@�4�'�T���t�O)�P��G���d_;h)Vy��"_���p�@[�^K����B��H�>���d����C2T�&Q1�%��K~��Cv����< K�HR�#_����G=�$1���SԒ�At'�%��rl2?9��Kv�I�$8��-����)X�h�R >�V"O0��i-Ett�	E��yW4L�"OPph���(4�r���"d��I�"O�M��K	a�V�ᵀ��#Z��`"Ol(�$HT�JVAA�*�Px5"Ox��i�_
mZ���� "O�Tuo�ID(�s��IR��P��"O^�1K��p��	�W/K�MrB᪡"OX�sL'A}�m�'��n�u"O�)° E(T���ۅԺ�� ""O2$�F�Yf�d��Fэ��5:�"Oh;7`�rj�mҒ�M2;�R	¶"O��㱊ďe<�Az�G.E�a"p"O���$�s0����.v�F<K�"Ox�:��K��z��WEɻC����"O�f�xh��BG ��cR"O@0ǮN�MXp��`�p7��{�"O���T�A�4i�wi��l,���4"O*��2Kצm$�D

<�qh"O���/�&f6j�B�� ����"OL�s� ��j�*4����=i�6�E"O�����s��)3�S��};�"O�d���R-d��a��=`�P�+�"O�ջS���JsE��9h��a"OBT@07l		/�[�ջ�"O�9�5o�N�P0Zp�ľ7�dy�"O��)C�شM8���.�a"OQ��#��R`���e�"n�(�"OpI���6��)��B��4a�"O\-:5�&^"�؀P+�0r�d���"O��-VM����ۏI���"O�(�2
�I���c��4 i�"O����В%�3��z�D��"O��8�.Z�#���Cp�ґHDz�Hq"O�iX��
�A���p���/�1x�"O��!�% ����m�k �-Ѕ"O"%�����a���|~�V"O� �6H�d�&x��4M�H@�e"OQ��NM@0���G�B"O\$cR�ݪF�B0pT��+_B��v"O~�À�&h����ټ'H��b"O<d1���Yh�� D	*4�3"O��P�h�di���"�h��d��"O��ڂ�&4��@ŦŪ�ZXa�"O�l:A!D�%�@�3�Ӽ��dyf"O`����,�F�1w��;��8�"O|�qf�N�&�����h�T��"Op�b���H������C�qO�0s"O�&��eVX�䁃�C9���R"O@t�r!B+oG��w��>1�f��"O�ta�_'2֔r�O 2ۣ"Oh(�BBmc�s�
���ț"OX0(�#�9��b�TM���e"O�Bh��1v���gԛ`��"O��7��w}��!��;��E�w"Oҡɡ��.������Žp��4+�"O��p��eA���$�.+�2�"O.�y����`�pB�����%"OV��S�*`�pLQB3VlR���"O� D�R BD����� 1&fi��"O�0DD�yg"d�PJ߄TQPh�g"Op���E�A�:b*�)7%�@��"Ol�"V���q���v��6Bj��ڦ"O��Cu���lI�5I`a�{rxi"O���3,A�1H�S�)N?|�$�E"O��xF�C3�M���)3��$Sr"O�	2S(M	]2��HR��L�9�"OP�b��-� 1�˥q����"Oн��K�`��i��+jMΕ�w"O �g(��H��g��{K�@�C"O��s��&����"�ً36|��C"O&`�� �0r�}��;"F��"O����:KM�i�P�N�v���"O���b�(W�,�4G!�D��j�M�<�"�NXF�����A_@����H�<Y�%�#e���oJ�cRx��ÊB�<1cf&C ��$#RG`�-5��}�<1��
k�h�O~x��pċz�<�1� 	 �t�ȝW�� p1�Xu�<I���R��1� b�O���Ю�z�<�C(Q^�냦<R�n�EAO�<AW�M>�8�D�S�R-�p � �e�<	Qf��,가�VO��0��3G@�I�<�A �(�L�spLF@��0*�l�<��!�)N,��&L�y�F��d�<�W�	�X6`rECL�Z���a�<!�旔(�B9��n�����
�^�<a� �O��τ�?o^�:��a�<��$>�N�1##Y�9�zm�� KD�<9m[+i��	VhԎai$ya�o�E�<�򅒵dX�ua�/��A���C�<A�ԚfC~=��H�9	��ృf�<�tKB�a@��w$�[2�X���]�<�CX�\��� �� � \���p�<Q �G�	���"6��4����p�<��	C�0x��co�!-v��sei�<�M-k5-��]�\Z��b�<Y�ȁ	ON�A�!ˢ�����-�a�<i��5�ͻ4O�6n1��I���F�<���S㚁z��ܲL;.�G��I�<�sK �P��9І0k �l�7�G�<�X�[X�$`���2`
� !D�G�<���E�3=�p��BɬZM4$ċJ�<��!ڐt'���c�E&:q�}b!�^B�<	�d[� �0�A@R%Aj�!T��A�<)"�X��$�� F��ݩ�*�c�<�	<,�fa�}24�]�f�!�Ѝ	x~���.LX-%�A4B�!�d��-mt�to@�jt(��T�5/{!�Ċ$p���E
*yU�9f!�4v!�d­LyX5ITH�SN$��ʞUs!�$];�F��g�N�<3�娢 �0Fc!�U� nx�r.Y:��Ľe�B�gN�A��_�I��`a)����B�	��vH��ԆD�HyZ���
A�B䉯j"�I��͕�`
��q,��u�B�
6������0�T�ΦTf�B�I�}����؇[�����gқ	,�B�	?76h�1!4\�� PB�)yvjB�0�0����E1_��5;�!N-0ofB�ɵf�ȇ�H���C�H�"�bB�	��ΈI�IT�_`M���D�!C�I � 1��B��2�P�L�	L�C�)� �bݚ\�T�x�	�.8�i"O(���)k"tj�脠}����C"O(]A#�ƀs�n<���5�L�"Oz�5��Z�8h��ӵB��i�"O���I�$���!���<7����"O����E��P[��6U��=��"O�x0�ј	��	1,�^�@�"O.L�!��G��򠀂�w"��"O���U�@)Gn �8P@ַiL� "O`���aƱ>y�,����Ek�#�"O`� 䏃�>>�bQ'�-WcRܡ�"O>		�kA'x��3WO�zE.���"O2��)�+;-B� �+_����w"Oja(SK��{R��JrJ�,R����"Od��"�Z�+2]�V�N7���8e"O�M�ЩۀM&���.�#)M,	��"OL1�,�	2������L7جJ�"ObH��%Lx��w�̶|�&ū�"O~����O�J�
`��̅0-�	
�"O�=��畐+e~d�g��$Q b���"O� �f��-w����O0P�r�"O��ء��ߐ��SG]�k
�,t"O���ca��E�Hk�c�d�t��q"O��э��y�D"�A����"O���� ZwX[����]��"O���b��Q���1��n���"O��{�#�8r4{cm�<B�b�ӆ"O���χ[���g)�_��"O6��7^+(�WI��P��z"O�`��L�@�!�h{�NL9� D���Ei�GI���a�3v(��2�*D���Y��� 	�N���Ce)D�h�"i��`(�����W�=�����j(D�l[�o�Y%dᚣ �t�x`eG&D��ӑ�V�P�,l��������!D�x:%"Q��:$ZE!�,20�DC�i"D��yFF_#��	�AҦJVUa�-&D�,���[o��m2%'Q��$��6�%D�h0���.peZ}c"��$
�5X�"$D���a@�� S��̗&�����4D�D'�*9,��dZŞ�Qw$2D��ˣ�
�>�	�pkp�Q6�1D��A��B���,[6Rvt�r�I1D�����֎X7Ɯ�7#��`�hH�.D�<AˆWb<5����w�,���	*D� ASo1Ϭp�ŧ�$����(D�����{�~,��J��yT*<D�4��W){1�I��&<{B��$G&D��b��ѝ*�E�D@_�bZ��3�!D�<���Voz}���($fU´e?D��kqhL�"����SJ��n���q �9D����6A�,�(��T����j9D���kE����m�f)����7D����f��\F��r/ȵi�v4Z�b D��h�@1'�%��dƶ�X �# D��"�@V�K69�Ǌ�P�Ҳ�0D�(q�c�
7����M�CHtPg<D���dfRv�ލ��]8��uC�8D�\��k�C���UE['+=��ӧ(7D�4Y�U�j� �x�E��4�����5D�H+�'��gv���)�B��U��A3D���*��,���%MK:K�Q���y2H�)
�	0�� "ƶ�%f���yBa$���b���p4�ޝ�y
� $�PM�f��{v�H&��]�"O��k�GΈ��*�� v��Q��"ONM	���4���)`.W"���;#"O8y����r8�\{7��i~ɦ"O����������[�.�0nYf"O,�k3�R?�jx ��̼]S,dR�"O�=�&�ՋF�p0�R✼@j��+s"O�	P�w-�<��T�J^v�� "OFYK$cV��N ��r��5"O�`��d^{�\p��&��d;D$i�"O(�q	   �   +   Ĵ���	��Z$�wHU���C���NNT�D��e�2Tx��ƕ	#��4"�V����c��mZ18�4��YX�ik���pc��(*�vpP�.J#�Ms&���n�.ԕH3>i'�ѝg�h��	ڟ��6-.)� I�
ц-.b�b6�=$�t�B�]���T)ҝa�y�M��9F�ԥV��I�K�4��h�󫐪AF6]�4��7A�	;:��i���� �L�nЉ�f��rZ���'��E.Zj���B��	$#0pka���]���s�<}�g	�Y��$?}R�׹T,uR6�X�<z2�^�����S��e��E>�xل�[��ē{+�1���*H�\c��jt³l@]�2ߟ�~���ha�=�F�2}r�T�d��H���0}�˔?hL� ����7�1�W�ŀ#p�(Fd)��|T���]?�?O�����׿%D�՚C+p4�Q��`�`��;}bT0F����(!}B�ػ�t�-O̴��߁	(!0�H�Q����p�'�|��#�(8%��A2E�+��O"�@�� ,�,�ǌ��5�!�t+�>b"��@~b
8O�@��ں��9OB���@��?e�.����l�&U�|��F2�? t��L>Y�L�1&d���Or��'�̭t�D�I�J�>����&� �~��G�.��^�	bGN�N���!��ݖ{���J��B*|�^�Ĉ��m��a�O\�Q"�qB���O, u�M<�󄄇2VlA����U�����*DQ�	�\��{�M<���(7 �P�t�|b�8����GH=IT<��U���t��Á"Y�I"$�C#>�����8+�*�)v����F���)����x%�qz��bb�3���:#c�����]T.����ŞK��0��w\�y���̛n���Ė�M��i�'� 59�C���DL�Ȫ�BMS�i���gÔ�<U��!�����D0͇\l#K>��L� 4LVy�<1�f�<TL���E�.@�)Ht�C�S�	��'�*x�@ ������`�
c鐸Iǉ�K�<Q*��y��@8��S
j���̌~�<�)�=d]3�aV0HM�=2Uw�<�VfS�0d<p���/o7:�@a��Z�<�J��]3���&��Z��P�c.�\�<ѵ!ؚ{��D:q�\�t��sw�@a�<���F�9{ �яRp�+�&�A�<�� Kx��$�f�c�Nf�<��� m�%1"�W%F���CĬ_�<��a��       c  �  �+  �7  �C  P  �[  �e  Do  *{  ��  �  W�  ��  כ  �  \�  ��  �  2�  z�  �  s�  ��  5�  x�  ��  �  N�  -�  _ � � 4 w �% -, q2 �7  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF����n��R�p%����I�= j���ML"H^��P�E6d&�B�ɍzD���r.&r<5�f�_��)D�DƘ=#���)��Ľ&�z�Q��Q�Q�"~Γi�p)y�-^��0���,�dn�v(<!��i���!�$����Wf�ߟ���>j��C3�ǟQ�ҡ��� =*!2��ȓ��R`�!]�r-�p�-���'�ў"}S⊣<4,��`��F|�Sb��T�I�|$Ex��D�ˎE�ƕ�AR&@���7�3�y��לs��ۄ䎍;����U��OT��D�"���2Wd�	iyd��ʡ�D,'�p|)�l��Y��M�w�]x�ZM�ƓQ&,��� J�\�� ��+l1H�F}R�6�6�Hs��bd��2�/n�F�F{��'o
m�UJ�6iƅ�ʍ�TI�02
�'�6��F�O�5��˨M�d���'cP��!O�����)X�@Jb �,O��
�8�R�ӥ��O�0��6��2ȇ�M�u
�	��^P�@�r�Тq4 ��2�X�1Oغ@3~�8��@oJG{�<�� ɔ���fR��m��)�t�l݆�A����PGE�Y�n��u脍8J���S�? �����W�p5|����[�Yʺ��"O�@��@5Q�����
���qw"O�����[�\�80#VTƦ��`>O�Շ�	�l�����ʆvzP%�"�����	N?Q
�$\6�*��ͫ3�X��r��%U����	A���L�㈐�h�fUؕ��0r��ȓPb3CLE���[ā������X?��4��S�O�P[�C�x�0e�9f�$�"OܐԈ	 TZz4�ÄN&������A�'��7�;U��l2GKįS��P��K�)!��vc��x��0�6��VM��s!���y8b����2�����&\�a~B[���w��)I�� $�9eH
,�r/0D�`K� 4M"�∉%i�Y�I,D��P���1������z-��:%G:��m?�ÓD�Nl�l�:$#��pq��d1,��uɛO�U��˓�B� wkT �?ae�'���	�G�q�� BgL^-r�<�I㓲���(�V�G�K�9S�E�1)���ȓƴ�0Ei�X�!+QꔦҒ�D{��'�*���7=�� +��p_�=j�'���`��~��K�ђy�Pd�%�S��?��'���SM8Z#P!���
[�<���I�,�p�{@�n��q(|�<�B�m�4y	D�y�Cg��y�<�Pj�6I0L���Q��C��s�<٢���.Y���f�ܗ6��`#�lŪ-��t�=I�S���̢	�
��f�ݠA��B4�ùV;a}��>Y��9'G�0m՗�*��a�Hy2�'.�A��B,U���Ar�T٠���yB�O���ȡ���7L(@�e��fSXC��Ć��E����t��2kJ�(�S�O�\	A�Ǔ$��Y"�E���Ka"O�h;Ц�� B��5�\�an~eA`�x��'������� �pr�_,ٔL���M�d3O���SC�s
9���ҿFL���`"O�AC���}�y+�dT-C�[%�xbX�%���e�i�% ���`���P;�rB� O2O�*v�%Ed�R�a�(fUX�"O��Ȳ.Z9U�P��B�e$\q�S"O�1�gb��T~�9%0!���C^�(�'�ɧ��x2 �?<������t��y�����>Q�O,��C��uUTXs㦓>T�Q�T���'i�y�]=Z��%Q����D�Z���Q�yrhY
&�Z�頃^ �[h�*J����?q^P	�F�;�����<m!�\&8���Q�,[�9ⲁQ�l�_�!�Dگ5�|���9Q�f�&�0]!�d��� C-����P��|tȵ�0Ot�=�OG�D�>iV��.�
�#�O�QF|MٷK㟠D{��I�,\h~�㷯נC
>�S�
�+�B䉓$�ި*f✴g�8HU�½Q�B�In�Xq��♥=`�����(C��hO,e�>	S��pH� C�݊ ���2�[W�<�⎇�ns:s�Ê ?2�R��T�<���I�)T�}��כ@��m�d��SH<a�jO�8��Ś2*�3dQjh4�	%&Q���	ǓTXQ(��a
�W��'aN�I��	M�'[���	�
"^��H#(ڠ�ߴ�Px�g���CϹlj���`c���ē�hO�������ޠ`��5��
E�.���"O�0�\z4���%�1��pq�i���Z�v������m:"�9q��i�!��ay�"˪��0���y����S�? � 1ք�-sh�x��b\�"���`����'ўʧ�6i��֓~���as)�>q��-��V��y��U�c�Hii�a;Z��ȓa�¨Щ[Lr^E���Y�'�H�ȓa���4��G�&�z�$S2/�nh����$-�S�!��Q��D��F�c&E�VB��6�$�g�@Œ��#�j�<!˓D����n�:x--B�C](-}����IR�'�H�#�'h�,�sXH4h��M�N�nD�d�eHV�2
�J���-�_�<�#��QZT#Q�-?�R�[Ve B�<q�f.�!�.��Z�~lKsl[S�<����<	k¤�B)D�bZ���WOS�<I�$.n+\���mJ�Z���r�̇�d.ў"~���\�d8�'�@9(4p����fi6B�ɇM��i���"T(�*��E�2B� ����Q!gPЅx��[2F�(B�z��"o̘5�M��A�Y$B�F R͋�oʜe�حa���J��B�ɿ}��5{�'K
s���"$$��C��*T�ʙoD�|s��E F�-��C�&cҊ�L��"�-{���3�B�I)_i eᤥƞO �廂艼0)
B䉂��w��[���ض4��C�	#/���y�W7fW��S�Ǆ<F,B�I��Y�'ǜT��e�b�B�I P`�Q��P�B�
8���2XRC䉳ALF�Cd�̟
,�3j	�4�C�#P|��XC�s�F�"��ڟOg�C䉅JQd5;�fլ)ht�C ܡ^�
C�I�'28$&�2 "�hҢ��e�BB�I�L����L 9Ӳ@�%��Iu$B�I�0�
8��,�ry2�� 4&C�I�tq��ѣ�0o������8U�"C�Ɇ@͹�BUq�M�r�Ϩ'��B�Ij�}�B@�#A~���f�c�B�!-��q�cH��u��?Q��B�I9x%�����`E0�B��"Ra�(�` 'ʬ�9���7��B��OL�H�&G!�rY�Ƅ̀>��B�ɼ �����DM�l��@W`�qY@B�I\Iu*@��i�B��O�"pWfC�	�)��T;���t��m�R���o�B䉇(��HV&�"z���iדp�$B�/\B `��Ֆl 0l�f
W%#9B䉁N��3��]��ָ1�=[��C䉯5$�m�2��c:�0���Sh�B�I�p]xt�0\� ���� �N?j~~B�I��@a���)Cˁ/	�PB�I��|�Q�M�q~�p`��B�8B��0 p%I�	�U0U�"��'+BBB�ɑ]1�H�4��9,�ͣ��"0sB�I^�N�"k�?d,ʔ�R�J3QAVB�9���A�һ	^|�)��!��b�X�i��./���ƾ!�d˘f�bQx*�/P�Jw��?R!�ǰk��#�Q0y)�!b�ڕ"]!��U9r,�i1"G�	�]H��@.6T!��!v~�z �iҸ���=!!�$ӗN�"9��CF�!Zѭ؛@w!�3k��!��D��g�t��J��!�DX(0+(	qݦ.��u�!���!��I� �Y *�%$���	S��D_!�����&��3J�&T�'��=#!�� ���E�3@	���Q�R��,��"O��.��Q���i���'T��0e"OlȠeG/T�
�[Q�M�[h��"OF4��_�U�l�9C��f�	"O����"�i�C'D�2y���'�2\��	ҟP�I۟��I˟��I���!�AJ�:
�0bl \<ҵ�	��I���	ӟ����@����	�2��X��Ǻ,�<���Ė7�2d����X�I�l��ǟ\�I��@�	��L�	�p�@d:����c2p2'g�eܠ���|��ៜ��˟�	�(��ʟ��I:!��{"ƒ��P���]�~�A�	��4��⟰�	ܟ�������h��73YH-*�c�'F%����}�J��៰���\��؟��	ӟ���㟬���vaPU�a��u�����Y�}����IƟ���؟(�	ş��џ��ɧo�Z��0�ބG��(��-һ#����ȟD���H�Iş��	��L��<�Ʉ Xt��g�G�f)*��F�T�����ן���؟��	ßt��ҟ����t���87p���f�9�Y�#��I��������Ɵ��I��8�I͟ �	ϟp��40Z4�  ���A^�$����d���	���I���	ӟ\��ҟ��	џl�I5j�C�	}�d,3â�9k-b���ڟ���ß�������Iʟ�	����	�E�� ��&����Ǘ-�L1�	؟�������⟔�I�\��4�?i�Q(D��ɢDi�!�ŀ��,_|�r�Q���ICy���O��lڳe>����%V/0�
Gg
9a��[F9?1�i��|��y�Cy�H�ë�?7�D$pw	Q:!�Q'��Ԧ���	���RC�c���.�$i	@7%B�R�Q����Ot���k�� ��<�����'ڧ�ܲv��EU��H��Ijj�P��d�����?��.�M�;Uԙs�M�w>��SdԤ$W��R3�i��7M�է�O�*}(��
��y�(�?4�A��.A�9)�e��y�<l�&8�rD݇B]ў��@K`��#� #ǀ͌+�( �7ht��'2�'{�69;n1O&���ƕ�q ��Z7Z	�K�B"��6����ݦAݴ�y�V��c�N�S=rD�����5�N�B�(�Q��Mn�a�|B���Nhra0��;^����*d�:��B(ކvA<��+O���?E��'f�˓�ލPЄ�cE�Q�uw4���'Y�7�B�����MÊ�O�:<��ț��Q�T�%"΄3�'�6m�����I�m��8��9?� �ƒ<o�yٵ��<h�V�x�OC�������J?���4�����'+(�ܣA�Ĵx� �c�Q�|<��'�j7M�={#1O��i,��D��@l�c9D�¨�	�A�Tϸ>�7�iL�7�r�'>�������ˆ��h��N#Ǥ�"��ޙI�4��@+�>	&%��>dZ%����x����21�˺]���
�+J:.c�-��J�'��	n�I*�M�珀�<ytJ�v^�)�vX������<��i��O�9O��m��M���z���A�=� l���՞��x�Agڳ��QP���\/�n����?���ź�`�~�Y"��H�T�XP	�ɔ�D�5�U�v�p�IUy�X�"~��ض
*h�F@G%'���&��N�>�FNܩ�����=$����! ��͐3i�� h@o��<��OLo=�M��[��	Z�<��>n`�\���<�t�_Q���	Qe:v�X�A��3����4�F˓�?�6��$���������<�I>�s�i�&]��y�S>�X�'�����S4hM�p8�n8?ISY�p3ڴp*�&7O.�
��@�w�N�9�dƛP�P���#��Vv�x��g�����D��9��`jSj�L�^��˄	��Ҡ��d�����蟜���P��?��O��ɏ�M�c-��^��͘�J�~��X�JN&2�6ϓ�?��i�ɧ�O�>!�i�q��lA�c���R�����t�0!l�91	�`�`d`�L�	:�4�H��Šx��'DRh+CfC.p�5��JԪh_����'e�i9nߟL��џ���� �OPĠc���%K���	O,�zk�0Q��4O��d�O�����S���R��yE%Tk���*Aq 
c�4O�Ơ�O@��|�������Qs�@�Γk�f�̂�CO��jEIj��tϓȬ��� T�U�d hM>�+OX�D�O�=BR�*��s&�__�f��$��O���O����<Q�iU�q�'�"�'�$�1T�N"B�4���ʸZ��`�U�|2�'!��r?�&�dӔ]�	Z}�K%7�dL����_�p���
C�y��'���Ú	?w:�HY���3JL��'U��D�t��/�t�����o:Fa)c�W˟��	П��	ٟE�D�'�T �`,�=�p#f�$K;Ĉ��'��7��'��D�O��l�a�i>�]���`�VBZ�G�\}�� ޳ho��	6�M#f�i�x7mJ*nJ(e7O��D�%�|T*�c؃yI|�#&��9d� �RT�J-r֚9�B�(���<1��?����?��?y"D.R�}����h���J��$Ц���x� �	�D�'��	�Ob���j½��=#g�EO��Ӣ$u}��p���m��?�N|��'��A�˼g��I�ş�#t���	=�����P���20{YS�#.j-t�O˓S
@��f�/��$I�OM�w��Y��?Y��?�%�E�S��Y��)�4��Pͻ/H���mڼ^;D�Hq�L"͓�cޛ��'(�i>�ٮO�xnZ��M3"�Of(��A�ߐJO�h�GX{�	�gm��~g����?��G�&�m�!�Ր��Dퟎ��q�? L����'S.Y���-<4P�P3O:�D�O����O���O��?��K�!��0���/=X�:b�h���ȟ�#ش G�'��6�?��I�R=(}b�gK�v��� a�9/�x�Ig}Rn�($l�?�k΍9G���ʟ��P����hr�*�cǨ�*xMӲO�%��E{B�'������2�M�;T�p���O<7X,�Ça�@%��h�4*_R��<����*��h�h}``�"Ä�c��F~�-�>a�ie~6�x��%>���Vo����!�z���%G�\Ya��P�|,4�3rM0?���l�L�Đ �����l@�+��T�����	1)O����<�|�'`n7��Y>��cL+:m�͑�.�,۲��4�޴�����'V�7�F�dS&=JfGχ0�8a�R�,��qm�����  '�����z�&��k�)`�<?�%%�M�@5`�Q=*��e�e̓�?�-O6�}RB�Z8D�(xz�ĝ�P�P(9�%��Λ�+�Θ'K����t�z��N��x��@h�/'��1cE�dδ�m��M�'B�i>Y�S����������7c|���g.�:-",�Â�I/�p�}F�H���]9/Y�E{�O�fJ8E�0���ܘ���!�U��y�X�X$�(ݴg�2$�<AWEIg����P+\�Z�`��I���?yN>�6Q�<��4h��:O"�6
ȥ�Ul	\x����~�*���?���ɜ8�(a���P~��O&y��X!m2	�3OY��7�8x��.�?�b�'�2�'���S�<��k�.�ʍ@�ix����៰:۴Ip��(O�tnZj�Ӽ{ �I+$:)�"��lv�WET��ЦE3�4qw���Z<1��0�'�r�
_��H��N� 8�����G�d�PD>��)1�|rT�H�I̟��ٟt��ܟ��H��`e6au�>��1Q ��oy"�r�H����O|�D�O����?��}��-�|�Y��,�����'9�6��oڼ�?�����*������@�` @�ET�`��H��y�n�O]��#ؤ8���N>�-O8 1coڠYY&����	{���B��Op�D�O����O�ɾ<a!�i���'���7J�Yl����*ķg���'{j7�-��*���MѦ}�4Qq�Ƃ׿\;��hE�Y�Q�fMPQ�$g6�����$1\�]k���D�|��\���m�>4�gdѾd#�d��		�M��'���'5"�'�R�'��ـ�섩@x�-���kt�����O@�$�O�8l�<T�u�'7-�O�˓ �D�#A�I�h����Ħ(B�h��'e�ɽ�Mf�i����B3����'��睺Zq�IYpfԡRQڼP���AvN9(��9aJ�(��|�X��������I��Uȟ��a�p(H�*3$\ � D۟P��`ybEgӊ����O ���O&ʧ_/E�Ʀʪ
�@t�BBT>w�ZD�'�`���giӠ��IL�+�(�+�Ӳ5�����nܺo߬EY��[([]�V�_�������䆵l�re�b�|�%��a�IQ)7�<SG�Q�)���'���'���dW��2޴j�Pmq���3.�I�ƪ 5N����)����Ȧy�?��Z����4w��CV,�� "��Q0�B�sA�iʈ7-Ӝ=���c䟟�#���r��	��"Syb$K� ���kPD4=h2,�EAU��y�]����՟|�I�p��ʟ4�O�x(ӣ��b�p-�VlۃT%��X��`�*5�l�O����O0����ܦ�]�
�P����,�ҽZe$ӊ^)h���4y��$�OT�S�'?�L��+��<9C�=]UT0�&˪ �YʁBV�<1T%��~�M;���%����d�O��Ċ�{DX\Sf�Ĺ,�(��灓+�,�d�O��d�O��9����2�y��' �s_��e QH2p�P���$A�O<@�'6�H������Ŋ {  ��#0uq0<��͋O����OS��S��]qF��<��'r���%�?y���
;�:3�O�E�� 2��@:�?i��?����?�����Oh��U.T�L���2PR�=B���O��m�#Cn�ɖ'd�6<�i��"�	8=8l-��]�"��=2�z���شEԛv�h�0%w�[Ip��6"p�i0�U"7�`Ѵ��a��y�'ܖ��9�6B�L�IVy"�'�r�'r�'s���7 d���	�d�`�pш�剓�M��2�?1��?aH~��t�ꆏ͕d���r��H!J�M��P�$h�4'�d�O"}j��Ի"������&�0��Q�1��e)u͙���d@-FC4q+bT�5�D�O0˓n���K�؀,���c���L�X�����?���?���|J)Oވl�i�L}��#2�qc�ޝz��cL�+R%*牧�M���ĭ>!��in�7�Q٦%30 U6)chx��\'6Y�(+V-!^�f=�2f!?�W���m"E�F���dklQ ]��Ӡn� t�x���>�d�O�����S�vG����@C�&�>U\T�Yt�2�.�M���Ie~��p�v��<�P��7~���!�#�*B��7�y�Y�(�4�F�'�T@0��G6�yB�'0*0���Y�??\����
�P�DB�HՓ���:�.O\ў�}y�'2��'�ؒa���G��.y�p�'�'@d6M�2}�1O �i柰kqo��z�\*��	�`�ԕ��s�O��l��M3�'�O���l
)QD"��U�j�(T���~ͦ� �Q�X�TQS�O��IU���*��7�ğO�4����^D\-Y�瓽5��˓�?y-O1���/�M+��G,�N��G�l��F�N!J����'�&7�O*�O�9O��o�9�:��܊9�j��&A<�
���4�?)b����̓�?�t�Ϻ){�5�c�GB~
� @�z��X�!�[��؃�������O���h��� �ޖk~���4Q*1�5����Ҋ/�	�?�'?����dC�*yZ��'��\�xB�@ 7�V	o���	G}�Oa���'|�yB�A��y���Ju@��
�Rb�d�''��y�T�Cb��Ff	�{s�'`�i>��	�`T��ɂ��T��8³MO�P�D�	ٟ��I��'%�6M*Ci&��O2�$��psF��g,3h�d"��5#��⟔۪O�lmZ�Ms��'Z��\Y���ݑ\�Ryh��H�n�ӟ��e�^@� �Gy��O��H�``R5Dw2�X�Q�n���D6�d�)c].Bj��'���'��џ�ʐ(ջf���T/ΣW�� ��`�Z�4]�X�i,O�Xn���&��f2IXa�O|��u�0.E6�牴�M[Źi�"6�[�>�F�0c:O2�d\�\�#U��a�d��b$��u��+ύu2�Q�P!;�d�<���?i��?i���?��� �'R�Ua�LҪU�.qP����A��`�ڟ���џ<��j��'"�adX=z�P�@Q.4g�4Q%ϯ>!��i��7��֟�%>��S�?=�l jWؤ� �Ғ�pBvm�>A����&o�py��. й���ڕ)��'�	�I�� :GĂ �d\�r#!�n������I���4&��6Z��k۴C6��;�Dx�������sEC3-��"��'���|�O�6���j�j�o�<iV��g�]jHPm[�]m0��E���H}��Iݟ��բ� 2���b�ZyB�O�L֘���0�AK"X��7��?X�I͟��Iߟ`��ԟH�	ŗ�M됍�3�BqI�!^.}�t�**_�؛6�'%��r��Z�7O���Iæ�&���qF�>& ���1NI��hK��?٫O~�lZ��M��?��s/��<��B:N���j��e�)Ky6٢Q(3Ax|�q�ő_�Lu'���'���'�r�'V��Ɗ����#��T,7�2��p�'�2[�`ٴʹp���?������F�6%Iu&�8g����!�!h���'R���ִ�$Ye�',�O���*�%Q�|P�.N�>��M0��M<���`��2b����Z�`���sXx��A�p�ɹc:(�p6a� �<1�� �(���Iٟ������)�jyb��Za��a�v勓�ŏwA��s��=r\ʓ{����'U�''~�Jb���	�ew~���䄲j@2M�Qb�#�T6���=8jM���$񥢔-&XZ�d��Sy�AG=�p8���^�Z�J�����yX���	ן`�����	���O�s�
��S�MzR/�pi.��eh� ��!�O��$�O:�i�|Γ\��w �јC��a`49��u��� lt��nڃ�?�O�)��j�ɓ�g��q��7O0��6�>u^q��҆-���2�8O6����� u�N�<����d�O�$��*O6�ѥ_��e[��եV]����OtM
ǆ����'Dp6MF���	�O��d�@G~0It%ϳ?�T��a���YJ��ON�DZs}�`�rn��?y�O�-IG-�4(آi����4q��U�56O��䕶+xyp�M�u\˓�j(JVvq���l4�dQ"�S�xL��(�ʥȄ����?����?1���h���D�/oBh�#��L��IQ#M�e[�����ص�"?�iu�|�w�N�;�G�:h��^����'�<6Mզ���4sM�)�D
�<���-�r@�w$Q�d�p�" ��[� �`ť����`���!����d�O.���O`���O���&�걘��_t�n�b.|�<˓^w��FƔ����'�R?�d��'�Rk^ Wk����"l���3�jˤ/���(�f�&ja����?��S��ԁYפ�?
W����]�}Y����m�w�'E�e a!��<�5�|rQ�|��z)�6@��fۚX �Q/l��OT���O��4�ʓ,��	��yR�Ѯ�\L�� ߛg�|C����y�'t�⟸r�O��oZ�Mcøi�:�B�Q4�I��J'ʈo2F��#�Q��y��'ߌX�[7(�"7Y���Ө�5�C.&�Yi�W�D��	ؑ�y��'���'�"�'�r�i՜_JP�������΍3V�R��?qѷi^��s̟��lZK�I"=Z�M�T	�u0�$ұ.M&�-����$�צ��ߴ��W�
[�`X��?��G$.l1����mbj|�� �(<W�\!e��	װ��M>1-Ob���Ob�$�OL��@j��� ���<=��[���OX���<�0�i�Z ��'Y�'S�;*lf������LϨ p�#	�m2��A�	��Ms�i���d"�)�����E�չ[���[@��4��:��8�<��o8>���2#D��R�V�XI>��D΄�p�cC�$��]����?����?���?�|�*O��m�xW�T��IR���#�A"���@�Uy�bi����#�O�Pn�;>�j��Gn�%f?��!���) �شb��f/ӆY�m�'.LfmN��eG��n�剣WO�u5�-��ʁ����|���'��'���'@B�' �ӛJ�����%�h��B Q�����4
s�]�'d��	W˦�]�A.�6f�-W��	�eF�M�4��4a�����Ox��|B�'���]��"@͓T��94h��u��y�qh�=��͓_����𭒹��H>�(O���O��`Эէ\�b��D�ڂ`R�j`��O�dχ3��у�I�<AV�i�)��O���'��������iK�,��ڐ�|��'L����Viv�
a��Z}�f�&��l3����/�외�に�y��'ب ��[�� Q����<q��ta�
�ڟH�dΰrq�yGD�eKZ�Q��ߟ �I۟ �I�dD��w
r�	p,M=q*X�-�
����'�'��6-H,��m6�f�4�	�çĶp�L�b�a�i$�@�?O��n���M��i~���*М�yb�'-�l�h�:D�Y�� P�+0�DK�,���D�{�.` �`8��<���?���?����?aa�I"6��QSp%�>Y�>p��hФ��dIۦ�1d�ퟌ�	ٟ8$?�I I3�;^~�ĩ�0Cpx$z�'JG}r�b�
�n��?�H|��'���\ R`�Ex�$�R-�mZC��>x��1V�����
�o
I� ؘr.\�O˓,/����OMT��9ዔd������?���?9��|�*O�n�3A!�m���5Y�$�F �q�E؁�t�$צ��?	0]�D��4}��Km�,e��o�-S��K���WaTH�0m2�l�2�>O��d��n���;Q�
���˓�����hq#rBE�g��`K��]�]O�Y�d1OV��<q/O?9h�恤<
f��V��0hs* 扺�M�Ѧ�@~2�i�����<Y�?�̄bL"�&@���J"�y2Y���4]����'?b�y�j���y��'�b�� �LF]j�̙�> ��
���1v�@ ��V�ў�S@yr�'$��ħ�W����GZs��4H�'}�'��6�=]�1O˧Io8A�(
;S�,h���Ý����'v��}��6�m���	_�S�?�.4J�F�Q�M;\�R��J�V��S5F�*5(J��&2?q�'i`Dt��iG���)r:�$V�Da�pRG�U�4�*O�d�<�|�'�6ޢH�R(���5-h��DH�rG�-Zמ��)ٴ�?N>��<��i����6%��؋Ђ�:4��Qgy�"��8��4O���M\)��f� 9t�ɧzѬX��̪ �,	aI?4�,b� �	yr��(T���d����4!��:�*�P�4a�b��<�����w���1nv� �GxB�l臄����mڞ�Mk�'�i>���ɟ\��g@�KR�	�  >t�@LfJu �dŢ.���=	T���Ħ�CV(&�������'���@�O�q��vhE,?�6H���'�RV.��9	t\��ݴbO�U���?���9?dL�Rf�T���cUG��y�����$�O`-�'X6���������J��I���;b�X�z4 ��'��r���rGh�6^���Ce}�����s%^����³cbT0���2f�XD������D�OT���O���+��c_g�ءc텤#����ӹ�?�׵iE�ٱ�S��Jش�?!J>ͻ!^��0N��eZrB���BJx�j����g��nZ�T���Hs�,��=T&�Kq�T,*J1�̆mE��Y��/D�1��g�y�Ioyb�'&��'���'�2&�(-�>���
<6�nXS��5TP�I �M�v��<����?!N~�t:�hk`P2Ò���HմztTu�Q[��P�4ś���On�~�i��6�Q�(P�/�b(�G�6KƜ�1�=A��x�,�<�rN��w��b��K3����D��l�da�w�	&M�����IȀ*Wb���O ���O�4�4���Fj �)�G�3s��рq���qĩ��yR�n���˯O�Hn��M���ii��{F�t�6+H)\��5D��*�~�H�'�e�q��!��@W%{,�	�?�1\c���)�HK�"�.\�1�ͭVZvx��'�2�'�R�'��'��ڹb���,z.Ah�BS7�>�qD;O��d�O��lڵ;l�IܟH�ٴ��WD��$�R6n$�x!�1[��0�u�'@�ɛ�M[��i���B�>]��H��'�2�H}Wx�K��8X�nD�qGS�]��D8f�ߢx	�����|rZ���I̟P�I����rړy��P��/,l-�Kڟ$�	^y��|��I)"=O��D�OʧAZܛt��16���iֿڦ��'��4��6k�Q�	C�S�?I�g��9I�xӃm,B���q�֒�U$ϭ?�� �'�4�ދ ��`��|��ݳ3���&�D��nq� �P+qR�'z��'4���X� ��4c�H�슋����1G^�hJX��t~�����:��\}b�h�(�d*�7�xx�4�q!@�x�����޴6�J|;�E��<��.݌Db�E޶x^d��*OtQ�E	��r�T�eC�7�,�2O���?y��?���?����򩒏)��=9�!��@#��� �4#q�l�'u>�	ӟ4��d�Sџ̳���Sf�("�E	���>SS�E?�F�k��hmZ���4�*�	��1B�	c/�Pi�ꭉ&� ,hMz��1K��$ٚH���QCEV�`�O���?	�)8�]���
�p%P���fO#_J ���?Y��?A(O��lڞ��`�	ß@���b�d9��OT�_)ܸ��ʇmS%�?yFU�8�شۛV��O���=.R��݅s�I: �ڙ=u�$�O�]x�%�,���d�<��'E�te�Cf��?Q���*V��a�K9V�����?Q��?Q����ß��ՄR���c�B�"&��i
���韈jٴ{Mx��'{f6�4�i�y���(�2�E��|��Cv�X�شy��f f�p;Ҩ��_(�$�ODİ4.	>-�0}zw��_����ah_�R�b9A��\�ȓOd˓�?����?���?i�v�H��`�//R
�B%o�<���x-O>�m�y�"��$��V�s�#U!ߌ[��a�M��fzr�ׄ��S�i
�1�� �ЦMBI|����ꣂA6]G&�g/��p���;V�B&�P��$:ڠ����	]̓O��I�P,b�nV�n������ �ZE����?���?qsC�I��f^�T
�4�~Lλd� �$����Jƅ�\�%���֐|�O���D)�v�bӠlڑIA�]y���)Xj����&�*لɖ&k��	ޟ�30��i+EI���wy��OG"�X	%x)-�cT,��
�O���T�I��\��՟@�	O��pOxdk�+��K��Iȑ��4�>���?���9Ûr6OJ������%�8*�h]!.#X����1at�P�n�%�?�O-n��M;�'R���qSe	�<��YE��� B��ʀ�4���!sgν!G�L���I� p��0�$�<9���?A���?ِO˖����%Ƅ�V��E��?�����d�٦-ʇ,k�P��ϟ��O�*�v@]�U֎!���K+n^ ���O �'�6-��yH���'�
Q� c���s����hi� �5�huA�h���l��+Ol�)ײ�2�3��!��ڕb7� �F�67C��#!-��.�8���Ot˓�?�|�,O*�m�$d�)�A��p���jtB���йHB6?q#�i��O|5�'n 6��M�(��&���EZ�C;�YmZ�M[���j��͓�?���vz��X,��D�]�\�h�D�Sߦ�C�۷���<���?���?q��?�,�p�2�����+7�U1!�T�x!*�} ��c������$?����Mϻz,�`Z6;p-k�O�pd��U�i"�6�Mǟ�ק���O&���ٷ_�Ȩ�'�B�V��R�V��S:mٟ'����!��]�ƕ2�|�Q���	�����
% m�S�Ɂ�J��C�W�������	iyb�e��9�4OB�$�O,`JfT�`�25����K�0dI�"���O4��'�H7-ᦱ����$�7����͊�Ks�h��a�g����O@ع��]pn4�T*�<��'1�!���Y)�?�&�� vO�����E:�lT��R��?1���?����?���I�OP�ZBe��l��{�ɟ8U��p��O��n�y�(�'�r6M>�i�a�'Ͼm�r1�V�8c(Zp�ҏu��,7���nZ��M��g������?�v�3>�P�z�q�`M�(|Ֆ�0qkٍf#t��*�D�<����?����?I��?��+��=B䍠�hD(Qz�䈒%ٲ��즩�3og�8��ݟx%?�	7C0��3��V�>���Ci,�0H�OZYm��Mc�'�O��$�O"d��R"�@�*Ri�3M�p�"͑�N�X�S������f�ʭR1eDP�Hy��^/�D��@� C�0�1��Yu��'?��'x�O���+�MC�K�<Ahҥu|�a�(�<��4x#��<�1�i|�O���'9�7�Aަ��4?��=��G#B��� ���?l��I*ƇE�<x��Γ�?5��3G�&݃�G#����T��"O8Dc�6� ����E B�|̓�?����?���?�����O���b*�*zIC ��r��M��'�b�'��6M�� ��$�O�LoZ|�	�l�R��c��HE�Q*��F�O��e����������޴�*�hƕE��8ϓ�?�m�=�D�g�H�<����
kܐ�I�oM:~wv�IO>Y,O��d�O�$�O����ܿV�6M��LM��U)�K�O��D�<9��i*
$Z��'���'����O�vR�c�ln��p%d߀.�Tk�O|U�'��\k$� >D��*���Q	�4�9:�I �Dǲ�w�C!i�(5����Q���d�>twF��7����耩�ēJ�JX�bcӌn���pꈑ.8i���'nb�'�r���O��	��MKW�(�@I[Ѥ+VS�}�A�$%t��'p�7�>�	���$ۦ���81
��;�+"W,ܔ��ό�M�i�>�ʆ���y��'��(���ܵp�P�q�U���G�غ�"�"Y>���R�`�P�'M��'-��'��'���["��[7����d"���:(�4j�4(�BΓ�?�����<����y�bG�cz0�9�Q)8j���O��Bo�6MGԦ%r����4�v�i��iЕ�O>y���8rkX��A��8��`�gh��,<Y�u�0fQ�$&O���?��M�x@���E#��� �l `����?����?),O�8n�&���	��8��?��D�Q.ǈm�fH[�� Y���?��S�D�۴1����O~�-��$
!k>j
`�b��:6����?�� N��T4�4 ������R�S  �۴1��PـbR�q�n�r��+	�lr��?q���?���h���d�[`P�����YSػF��_p>�$Ŧj"*?r�iib�|�w�ָ�U)�z��Ū1$
C1��I�'�p7��ՑڴM�<00�ƅ�<��3RPlf�@�qm��*��՘zoB�"7E�J����!������O����O~�$�O������vJV�x��C ,�!L@ʓy��f,�&���Of#|��%K=X���;�_� ���80g���d��uBڴ��T�O9��M�03���(B�p�Ġ�V��2N�T3�=��I�u�+�/(����|�[�tIgJ mfxٱb�;-�j����Пp�I͟���ɟ�gy2l��Mr3O�|ôWxxf�"�L�223�	���O�l�O�i>Ѫ�O�n��M�½i��Yj�i�r��E�I�>( UX�#GS�,ٞ'�Rl����r��	�?��_c�����!tq�	K�ᛸB����'�"�'W2�'���':��<j�N�-%9"`�@�I��mM$Kdb�'�`r��A&ɬ<	v�i�'-�� ��2��s���9*�2ђ�b�O �:�֠���	]�L@X5O��$�4F@��!k�w��ERW-H��UJS{�Z�S��7��<����?����?	�#@D���
A�&|���)�?�����ͦQ�������`�OqL+ GD�X���KI�:��	��O��'xR7-�ۦ����'�F��>m�V�r��A x<����O7V��q��[�T�*O ��X/I�b�z�+%�d�S���5�H�]��8��EF�k�L���O����O���I�<Q�i�P�G�P�,�  ��#9�X�"E���̦��?a�[���4
�޼ c�
8� KШ������if6-�s��9*����1��1<%`=XT�AZy���(k��`��b'�P���yr[�����`���$����O�X�7/S.L�δ+i��|4�Eб�bӆeZ������s�'rV��wH|X�D2fv<P#aG�"[�a��n�o��?ɩO1����C�W� 3�� "d$�Z�&�: $$�Iq�0O�ը����6X|h�@"0���<���?��#@�or\͚�$�=V� 6����?���?A���DҦ1p2�~�L�Iɟ�
����bd� .�;�����j��_[�ɛ�Mː�i��$�>1$���@��J��=q�Ms���<1�ri���P��=*U(�/O���]��L!0�:i�w��D���w'�!T}��p�"O �Z� $F]�1�QG\��'��1d��"�2� �'[;�,�ML	FHz��ӥ��U���� �?�d��'�%q����)GȌ��OIRʉ1Q���"=xh�w���d��9W�.1ӲI��~���KƅU��m��m>7����J��nHP@���3CȸQ��7P�.>����&I�L�X��$X$����X�-��$mംL<A���?�M>���R���j\qH����&��i�RgY
W2�'�R�'>B�'��'P�P���C߾qh��9~2&,	F%S�-�Ob���Oz�O`���O�EYbN�� ��ˤ�ի4}<�j�-�n��D�O~�d�OV�$�O����O&�[r-\�|��A�▨xj=�t�ԦI���?����䓹?��	�`�x~��a�!���j0���b,�y�F�i��'/��'���'��1�U2��D�.����P�B�"r���w\ul�ݟT&����ݟ��Q����\1u�S*����$#9��1Ra�ߝ.+�%Q#���S:���Hո#{�)�������&#�j˒�FZ���נɉ3!�D�  �h ��{C�Ċ���s�`��
����K(Py�8�����:�t�e����S�R�<2��H�↋Y���ڦ.y;\��S�[.w� ���/��W�:�p�D��`UD�@�e�J�%(Mc�0ыP8[�p$��,�: Ú �&������?k�a��,=P=�@��Um��%bJώ����?���?���x�{���UQ�d@�Z:A�RBJ�\�A�cQ9H��G�zb>�O�[t��	��i��߼f���S�UpV�������r5,R��q��'ؚUїė�L�Qr����R��F)y�
�'��\���|�����'j�e��d��=6�E��,J��0b�'���/KȠ�S䇖#n�0��On�Fz�llӈ��<Ɇcí.�@���v�0T!@�}id�:�e;�?����?Y��!���O��dv>�8fM�%"�\�shM�x��1Ai�w���2�d�(	�L ´�'�@I��$�D��2�K' М�dB^	qw"  +'��(��$�3�?9t�ϼ2p��!>��'\���C_
xt�axХ!zKF�����?�Զik�O^�$�Ob��Ѧ B���=���+��0c��#D���e�,^"��y�[Kۘ��4�>�	��M���DG}డm�ٟp�i��F��]ǔY�́�06(P���OP�ć|����O|��k��(�'kD�
S�'�R�9"�:PV֩����\�	Ǔ=���8��Z:����O�Q��ȕid�Qw*�7�h��'V8����NS��`ӂ�dZ�?2���'@Ȩ]81��N&D���?q����m'�5R*��e f���

�XE{�Ob�6�;c��`v�NT����	��K�����<��N�=0����'�V>)���؟,Z7,��F9�!�^��	-i���O�8'��B��x����:Rܡ�R����4T>Q�fe�1�����O�r�JTyЪ*}R�S=ļ����[�J�"�`���M��(�:|��0���z�)Z}Kp��Wf�6�(P��>)3�՟(Y�4|���'2񟮤*��5	&d���6Z�<����O���(��|LŶ&�>완
8|���;�O�hO�IV��E3ݴ��2�^��e]T��]��\,� ��i�b�'|��Q1ҼT�%�'!2�'���wf�3ѫP/K�>m�H/L�h���@�'%�
E�%M�h��z�˘�g1�LM�Of �E���	r�(k��� xL�P"bK�j���c�*g�����&�5��v�~�����$j���*x欢aDXcI��z7
�.*�ڴ|7剻PX����'�B�'X� �&@ �h�e�G�YpF��O�x�N	�W���)fj""��h┟�Z���4�ķ<1P�5͆M���$]O 1�c�ߎr���#�*���?y���?����.�OD�dk>y�I!C�n�@#o �N��qI!G�@Ā�W�H�� ��mS$��0��$U�]���hv���l:+�:o�:��t�L�7N2A袭X������ w����D�l�xx��67��l�P��l��4kdᘷ\���$�ƦIx۴�?.O�D'��6m���ծ�]�8-hsh\%tC�		w����p��>6X'K�)
�b���I�ğ��'�$��e�b�e����@rD�?ј]ڥ,ҏ�%.,5(����OV<�ŉ�Ov�dw>����3HԠ$���7歫��/=q� ���51�l�IZ�güD����>"L�9xg���~���*�T
$��d�r0�y��V�<���JE ޡ8@��DD�ظ'��\�T��'
|��j�<<��z�jF�G�^�`�'�0� �H #��) o�+=H&$��'w�7M�
p#�LQ5�F�)�2�ؒ�Πz�6�ObŹb��u�	@�Oab9v�'&�HP�	�!_�� �u^)yP���'�"��i <5 �%��8DhHPg��9i���'��)�0#��kg��?>�tHD@�[j�G�H�����
�`P � }��y��	Ǻ�aJ���t� �h�P2��րM4bm�4�Ǥ�� ���d�O���|��䤱���y*f���\�l���{���O���� �����n*�yʂ�A�g�I��'y�#=y7�ߍ}�(��(;.�Z�!I�x����'��'IBM���\!��'<���yg��QǬ1�lβYyl�r 'L�mԜ�i��,���(0,�w����q�dΚ	ynQ��N�j6HɄ��� �A���T��E�MBV�9B适0
�'�^���|������;/�d%��F�Z�>�q%�*�M�U�iK��֭��,O���_�`ޙ˴��&1>�E����YJ��=����4Z�xZ1P�8&84pč����M�Ʊi��'��I1��OG��6?璈��FJ
�xx�W�h��h�'����˟����Zw+2�'��E�3&��B�U7z>|��6U9�$dκ0�uX���p=�A�I�AJy���<�c��)�d�Մ��#��p)=\OB1!Vn	6��D3��L>�.K�	�/^��Dm�&�m���L�'P�dj�ܙ�%�A2�&\���á�!�px���Qߦ=�.=�t��F�1O���'�	9JlىYw���'�e��L1ĊA���)+�D�E�'��!��n�b�'��)ݩ)u�x��|��ޮ	�>T+����m��-2�ʚ>�p<ab�Q�~
t�&�``�!�63T:��e�X]�  Bc�>O�T��'��'R�vFT�yb�L.�������I����?E��D߾a��y��X(�,qA�5�xB�`���K�F
�,�*�*C�M�E�&=O,�9�������?������_���dM�f~��g�е^���{�JE9]�����O,m���4,Ȳ�7-B�P^Lu��_.���R>M��"�w}j�!�c �8c�4}��J�s.J��Ŏ�2r��dk�A?�pȓ�G�;Y��\ϧcIb%3�+�*L�Ƥ2&� f�}�O�IW�'26�Ӧ���e�'�`8�E����d$CS� 5�>h�<����<y���*~�~T� ��	m��YRB�c�����>���U�C�p�8��b挻[�j�
�Oz�d�O���7'�+�����O��d�O��; YdTCv*iK }���]���	�y�	��<�w��=�
�xBߘ����eEJ|�o��T��ɘ^)���A^l�l��F�S#���M>�C�Fߟ�>�O�=rC�D�@.nx�DL��~&��p "O,h�dIF�B}T��Ԩ��+�n����T����S�&B���{.�P�#��(�)�a�?K��H�IƟ|��柈��(��>�9�R-+�H�c�7<~]�0-W�	�A��&� -�qC�嗬:��c��dЍdx��bg��4Z���8\���d�E)8N� �%j\,R#��eis'b�4&�`asÔ��1�C+`6
����*y�����O����O^ʓ�?���lߔ+y��3��l�ʣ��>�0>O>a�i	> �����W��@V�]�ya�6�';�Ʌ-����4�?���jy�)##سi-�g�Q(q�����?Y�B���?y����*L(�9��a\(MrY�!�
/r�+$�Ɉh�U �͍��^Ի��+�p/� Ack�U�E $��=�=���ޜA	��9�A!$��Q��;1�.����SnB��[�b�O��<�1�S���j'�(e\���LG�<Y���?a����U�9����V;I%����1}�!�d�̦��E�=Ld���t�H������'��@8G�w�����O��''ٖB�)K~l��O��IQ.I���	����?ap�ր.�v���S;K�왣��2!L��@�t��SSX��D��1+֡�����E�8�v /7 �����P�D��' &TS|��1�X���$�J
�!a�0hV<�s�>�S��q�49n�6�' �&(�Y�Q�@Cj}���ɢK�1OZ��,<O�1����Tt��/B��G�'ih#=)���:&�d� #�"����nĺf��k���?��B|�j$�9�?���?���h�NڼE��h��*�3吅C��D�xUZ�M�(��ڒ(7�+k:擬��Q��[G��2�T,r��N�vB%(��٣N�������*7���B�a���O���E較�J�W/�8:V�G�,%F��3�Q#"���K�<�ޟ���?U�?��Lh�@�w��҃�Vb�<��߶d���rd H�L����t~"
7ғ.~��'U�%*�:���ڠ6��P��%7?�C�I/&9|l�wK�O�d�`vdN3��C�l$<a���x�(����Le˔C䉃#�����Fp���Pb��G�B�INಭ�n��"��&i�7}DC�	!_\}�&S%)��+a@F�z3�C�I5s���-�u:���FXJ��C�I?SG�I����5�ڳ� .(�C�� 9`xy��
�O�Qj����_�>C�	/XjHđ������{��>C�bx����낑kY�uYb�U��B�)� �J�'��
�G�8�D���"O��H��|Szq������@�g"O���P���H}X�����zj�i��"OP��KA�Y/��%kV1G��<�"OJ���͐�!�1�
:�ɛp"O�� ���~Ўe;�I޷9}Rٓ�"O �i�.3�(���	G>o��� P"O���gl�@X��ߝ����""O�1��׫>4�<�1(�.�"O\���һ.lt��mҢ`� \P�"Ox�(B��a��;熨_���*1"O����S(U�Ld)�`Y�q�Hy�"Oz�*�̂1�T0��6A�b�r�"ON��E)0V����B)�5l&��4"OܴJa���s�f10B�D?m`6�p�"O��b��	�n y�ŝ
S����"O�0�Lܮ��v+��pC0��"O�1�-E/~Y���L�=2� '"O�4{�g��p% �iAj\P"O>$��a�5t{TVc�E8\P0�"O�<��Z#V���T�֪
�R� "OH�������B�4}|-i�"OJ��J�BS�9[��R���"O���g�؞�Z,��T�;*5Z�"O����l�%Q������
)l����D#Q]P�����"��͙5X�T&-�ShO	Gr �6#��?���@�i�x���t,P�ԉ���18�pA�$G�u�H�ц%T�(�\��K7t�r�[#��:-�Q���']���S��A��Fhr`d�9dB��4g��%W�Z��!@R�P!l�M���[�Uj�ȃY��:Zc���#ß3\ޱS���?���s�N'lO~����E9����O��N�fu�	�	��A��G�W��e�O(ā��6/H�֡̌N� �2�D@�<�%���>�\���!��}��#@"�8�1t�E�N�����DP���O:��cDE� ���(���~�bG4OT�
�N�"�< Å�6�:��g�	�&9^m�Peā/����"���&	j��ŖȰ?ц -r�r٘�Ñke<L�� -��� S'���p<�4�+��1Y��J���gC*����I�f���A�8k��	����+8�-C��
ᑞ�
#j��I�xU��
� P��>AL_M����Rڂx��A�L�Y�'A�t�� ʹl�,����pI$�C��D6���t��n�i� @�*�ioZ0<N\y���Mr�I-	l#?��CL�g��������j�����[?A1OΗV�8�ZPc�'&����%��S�'n��3B <[r��'�ޠdi䎎�}���?���T,.y���a�ݓ�G�B�jd�% ��(�1RL}��	 R�L��p<1@��"j�H��#N�p�&m�i�-+�CW�C��	�o�v���_:�)��0;��9���
}�I�☘�.�Z�	�'J$��P u�~�%kuD\�n,ڀ�>�p��c�c�¨`������Ny"����$�O.4"p$�=q�|ZČ<?�"=�u�'� ��t�ɺj�uRa"�6�,Q޴�9[SHݕ�LŢ��S�eJT �=)g��0�yre�0@��)����J�i&�_7W&�D�2�ɚE�T�&�t�um� ;ў Q��T�D]�U8�$�+bZT[ 0E	LI�{� �� .��r�'	��ra�2��i:����h �I��c�`��,AǓF'��Z"=��Iz�Ξ�����K	 (�%�'��	���Oӧ�O�fH#���(�eO6ymʄ	�S�7Ҡ�Dz��1�v��/��v��ѡ�;��$��y���u&�_�X���/D��� 	��r����E�������^BŪ!�O|����8h�J��b���J�̊P�i�= �I	q�L�S�K��
�:���]tB�P1�T:��TE���+�O`�nZ3zr�P�il�h$�F{2��#�U���,<��x"��9Cp8�� ��~��g�S�~���e(ڗ'ª�{D]�q���>�p<R��Zhr���) ���A�ضCft����pTqOr�	u�d�|�Zb�@$Q!F�+u`P�����?[�B��8�EE����D��yy�Cۿmm��'�h�yV�P�u� �"��G�&�������I���	rO��Ft���K�s�v�Ϛ�XA2��p�J�lV�[��
Hæ�QFγɚ̨t����On1IT�D	��Xs��5"�h���E���u׈iR'
ہFJn0IP�4�Q&���̈́ *7�0I�\�
�L�i	[џܲ�'��	0�2hyЅ�=rd�0���S�3���%��G�H܅�I�Υ�F|�%q�(�t��M�S��
*1��)��6�	u?������OE�6�݂Ԁ �!�F��\{��9��X��P ���ɌVG�@�f��}{��d$Q#/� ���ɑ/31�yk�@������\y�1��?��'k�DQ,z�^�XD'��(,r�D4�,*HW���q�&��46��V���5�R�ݘ�&��O�AL.&�\��� ���I'H@П�`�E10���
F��4�E<ړeH͚���*%8X��ߌs��%�T�Č��O���4�	z�" ��4b� ,��i׍{�� �'%i�pA��	����!��n��+D�Լ/ǔT�AO��&V8�b�&�Is����5Zy
9q h��p1W�_��������HO����Ҹ��ǚX���aU�P��;[�b +�E�:��� l!�I=�M��%kN��1'�"�X�o�,��|�4M:"�������ګF���m��	�@�v
���]y���<}y�"?�3&�9d��sf�K��8�����:�6�\�?NL|�dA3�Mcb�~ݹ����Xm�D���!/"�	�G��M�nY�ѮX�q<Q���*�@���p5�
��xr�3'��䨸y��i<� z�RN���{����˂�U%H�urq�U�,�.��G���<��"AG����&�^My-I��(�$���"`0u���I�d���Y�T�`�D�͋io�x�҂�>
�H�k ꝅQ�t4��!+�l����T�F �XDW(��y�Ʌ@B`�Z� �'2��T�-U�Y���LP�*O.�ƲG��dЖ-be��'��z�"6Z�����m[	w���x�'���@ql�.[J���o�/~<q����m�F�kWkO�><$�ǦΌm�DL�����%IGv�f�jW웖7#ўyQ�R}*<��[>��+�K�W�*����sx��� ˦��J�;Zx�����-��m���Hx����jޑ����i�tȪ�3dٲй�D,D���  :��K�hQЦ +'�g��B&KW<�,�ߓA�l��GҕC<�"�MF����I�N�$\;p�Cb^dC4�Y�/lb��y�n�;qN��ЅԶX��eIV!�z�||�P�L�+�l��J�$��1����J%΅����yM�!#(��/�tx6��"0�����	��'2=@JX	)��h�D�S:�<4M�1,��Oޱ��Ģ��ۃSd��I9G"��wi��� )�+A�Hi^�}z0b�'��X�AB�8�j�ҁE���0	`���H�F��wGD/aL�b�NN���dU�<�Dܹ'��p&N0V��#g����4��l��C0>�YI5�r�iH�L�&�?�qĖ�t�1!�e��t	�m��K^�lXJ3� 3�6h�	'�f�8wʙ�;84��+ �66mʬXgN8t/��|��i�&��O�m��݄y�����W�\ˑ��0�pxQl�+q���b��ו\I8p��WE&���	5 V���
L�dh�@뛙RY.Pd>��y?���u�`�'GzL˧K�l���_���@�}Kr1����:8�d#ǓBY�,���w��pE�Y�^(�@��l�,���>��FA
ve�e��5���ʧ"��1��/���	w���p��>�"=�Է	� s��NQtd:Wg�<y����(�B�Tzxa�Mئ���'�~AC���`Xԁ{���Z(��4��`���?yߊ z�U���;=<�({&l@Ӧ�YH_�J5z���6%O�j�gyb��~y�$�UA
, AW���A�ߓHX��Y��A �sу;t1���%��퉦(���.S��j�*=�F���!ݟ�0�(ڬ&(B���c���3��}�E�ќ>�]�$�xR�X95)���A�J
k�u��BR�ge����	�k�(�oz�Ir�e�	Td�����-�0+BGڦ��DM�A�ae�ɌH����H�Э�e��W�t�a�)ۑ����S�\h�ٰI~�Zwr�Q�J-U���y�c�!@AN�b[H�>Q�B1��{�k� �N�`��W��0���,����e��+�>�)�v��00��8߲��䚞O��}��dl��z�$�*>u��8�	ǾN�� 2��>�uf�=�C`�S9�%D{�.�'�*P`Q$��O�b�BY�(O�$÷&�Z^*˓;,��'*�j5���^����P�yo�m�����S��%�'	�K��~��"��7�89�+*i;�y�-�\Ax�ӱ���	4#>�1 ��	�hT�<j�8��N���D{"
X?´Q�3}�O�)���
�(�z�a�HR�!Q3C��"H{�1F|mO�z�H�3,Z�0�p��!O�UI�	�H�8&oˢEV�7홑j�� �"ЈO��ٶ`��;��7-L�3n�D�oA�9���w��<��}����Ρ>W���w \�s�ڢ=1g�|0"�)�#-y$��\{}��i�I eژ�S���@[>IA�	�t>p�+YP*���G�;���J���0�4��/\��Š��OĪ�x���h����'lR SbH�B�
��쉂B��?B&2A(6�Ӻ�%A{���+ �LI���_?;��\�"5�a(�Y� (?�'�?*r�N�Q��ٝv�	:�����d���~���"��֐���d�=$��O0���ስZ-�\�B�
�):���i�:�R�����0��9O�Q�FbZ��y���D��"�',��)�����:�"��tOԻK�Bx�V�Z��$�

wD�3ړ~A�ɐ�G�^�D��V�D�&Mta�,۱L�~e�a�O�4k������Q�����q#CT&F/v(9B'�� ���>w�Dd`�j�r8�Pr��+�Q�T�D�HTb`ϧ=p��a��S%;�N4K�O>샏����y�`?�8-"q)B�6r�JuD��6B6����I.���V�<9&�\;���"� �"@�� ~�29t�E����;$�	��M;@�
�|�d"v�ʫ�F8�;)�Bd]�Q�pX���Zց�q'V6-��)�,�����G���S���	���'#
���n�N�⥘ҦW)hn*�8�i֛F�Ø8����Q��
�) �ʚ�hORx���@������+|[j\�!U�W�� D�J/A�X��=��`�'N��"w��A�~鲇J/��,�H2g�A�<xEh�0�P����WUP�pF�J_�@�5�|B�Z,_
@���u7U�/5cÁ�C��{C�`�f����	$<
���D�́c���L�\@�'W��5b�JM+G�r"�ۗx*2%qA�LC�U�����Z8��ŀ3A]���s��:��ǙA	�aB�b��V��}Ke�gӜ�:7 �hT��"F�/)���q��ݗ	�ѹƬ�#]��S#��x��6�:W��q���j%�gϴo��>ړ(;�p#��;��3�Hh�;�lG�]���D�P�]���h ��;��O�S�'o��]b�!����!Z��x����V�P`�4���w�x�C��|!�LS���MЈd����T��H����2�~�7E�V�6�'9Er���Γsd��ħ���$�ȓ�F��j�Y�|�5��1�$l�ȓl�A�c Z�~o4�+�h��J)B"OԱ#d/�6 �69����nMz9"Of�3F���^LU:���:�ɠ�"O� i��ӨD4�򅪙��r��e"Ofى��ϖO<j��	���(�"O:,bխU#mT��s��_cR4�$"Oű�g��?�f|�I�"^�H2"O��᠊>.�0	��IL�OZ� ��"OЭ	�� k^�1��V(]J�0�"O~-��@�*WD�p��M+;�L�"O��w�L2>�I���#��q��"O� ��$ѓ%(^�:0�ٚJ�2=�"O�=@�GLh�9׆C�P/�P "OjX����(� �Jg��C��X�G"Ol�Jg�!¾��t�)EL(�$"OtxYh���d��5G���"Ox�p��V5��P8�'X&�"O�a�p��%(�i�1�H�%	�Y�"OH�e攄b\Z͈�� ���"Ot���z�rԸ���2��H#"O�[�"ȢYi^T	��Uq] Ec�"O�� W���[�D�"f�Qk�"O+�(�?O����5��;TV���"O
�96O,%
��߆�|�b`"OVĊ���q&�@��B�;�b��@"O�X0'�$mpP���C���0"O�p���;h�؈i��R�tq�IxU"O u�s�X�h ��g�	EcV<��"Ot��ǯ�+D��9�u��1K��1�"Ox45����{VH�7a�,t��"O�ᰕF����ǥւo�4P"O��C���3]��$A�&�*!�����"O`A؄��7�N	p�&��Grd�
�"O�$�tiA�i�������y\�j�"O�(�PKN$7���X�%^{V2���"O8��F�@� �RԚR$�7Pȕa4"O�L�0�0Y�u#��&NRuC�"Ov�Q�-ZH6��� ��+?��n<D�X�N�f���àm�&�q��.D�����_g��퐶��<ޕ�r$,D���4��+q�H�@�L��@�.(D�d���G3Jh���G0�5��!D���0c��P��MS�e	\��d >D�t��l$�m�PI�>8J��I�:D��0�YN��4�/��r$�!i$D�˦�J�N?~��U�R�:MD W�!D�X:T�ġi"�,����	R�Ԉ&�?D�L���ԁ�E�fִ�1�U�QZ!򄗋eo�B��B�8�ɂCݜ*�!�� �-����2u��EӕG��V�`(�r"O=�v�/�>��)>�:��"O�C�O�A�5�ת�x	��"O���C@[?Y�������&��d�"OvHs���\�:U3���%Q:|�E"O^5�O�'(�H(��$�=4�f!�P"O4�r�a,x�zH1 d+�\s!"OI1l�b�	��C�a�B�A"O2�K���<<�Y7ȕ0�|��G"O���LӱS�R)�6*�o�0���"O��ۦaǳhZ�3h�_뺡#�"OJ�P�N�|vΗA�e2���y�_�\�D`��K�)�:Ȼ�(B)�y�kҲ3�%IϞ
�`yQ�+�y"�ϣ[�f�k�"F�jW��y��e�DH:RG�U���/F��y��	|G�Y[�(UB����?�y�kY�)�4�B�/�=�29y2g��y�a�7�d8bH'RB�+�@�9�yҮ�\������[A���y2�<{g�4�AnR�~9��SA�Z��yB%v��|
���"�b9�@�ޠ�y�I� ��|AV��+mo�d⢢^6�y���2y� +���sjl]8�)��y���81*y��E��j�.Tq�Ώ�y�&��DA��"�!_�f\~�!���y��ޜV�*�(0��tv̬��Iʾ�yREϛz�"}*�O�n�p�+t��(�y�G�#HF(Ȇ-�a������y��
*=jE%ՋYn��v`�$�y�j 2��7kU>T�m�GK��ygU�bV�� uƑ$Z�Dx!����y"f�Z(����W�V��'�_�yO2^�����/��R�<9 5ʆ�y�W: ���GNڸH:%�S�K?�y¯[�(� ݮ8.ڹBѦW��B�I�|z�r�e�[��	K l^0r4�B�	+8I�p���A�P��h]4uQ�B䉀�3ێ��jڤwD4��`^M�<��	���uK��i$���HB�<yЭ+S����	�v$�"M�|�<S,ˆL��LAb��%�tT&�_P�<	ɓ1\>�C����)ڣ�D�<كǗ(<����O�� ��o�B�<�	Y"3��˱�F�i�^qx�/�S��p=�J�]~0�J��=ᖤ�gFPH<I��:�&|0jңIdi��≠!!��~��p���kA�E�� ?p���G��4$@�2+U�o9 �Ձ?�y�aKcb�k�J��d��p��J��y�gO�琌i��6_Y�`����!�y�f��a����O�m�J��b�yBH	0-��e�0�)g�B%�"����y��Ԯp��A렅�+���1b��y�&h�������o�
I�"�	��yr�1{%2���E�n3⌊% ��y���6�S�j��kƘi{�3�y��)�'.�Dcu��8��y��*V�L��ȓ)@eJ��R0,����®8�t�ȓMXp�BB' �U����2ECv, �������5J��p&����ń�p�'��m��&O�t9�U� ��}�ȓRBF��2�=W��h�0Q4��ȓi�}R���K��XI�b�/4q`\��S�? Z�p�j[�[����)q�೒"O 1
Q�K�|8 ��m�HԀ!��"Or�{D��8|�V�׫}�ܰ�"Ov|���ČI���tMÍhM���"O� �%ͺcUL(E�О6,(3$�'d�	�ozt��0o�Z�s��("+�C�I0mjب#�$�� +0!�'.�C�ɒeh���c��!�4������TC�	#��a���Ċr�Np Abɹ,��C�Ɍm�4����[({��� &�<��C�	�M������!�l� �ѻ3��C�Ƀ�J���L ^�^��E�óc�vC�	0m�<�j���Wf�[D��m�B��3Ik���m @M�]�dj��00ZB�	`vY#Rm��C˒W��ܲ��'6,(�e�
9
u�
�"P��I�'-�]�rFT?u�Ց���t#�Q�'�(8�r��r�J-��mZ  ��D[�'�h�R���C(v���߀f$��P�'ňRG�N�������]F��'��9$���>�L��W�x5��'L��Y�F		ygJr�]�|��p�O���$�Y���ŭ�5;��Ƌ=a~�T�ܹ�/O���d��5#���J D���tM*Yp���B��Z� ��J�O6�=E��.�n>B�3��.Hq���蛦�!��K�v{��x��p�����	d!�D	0�&�����'g� såW)p!�$[��bI��_��\��!��|U!��ѴI�f��nS�'6h�C2?��� D{����]�L�T?$���4D�p��Ç�;��ӓ(�nO\���f1�hO�S�ౚ�k¬*�lM"g"Č�C�	 Y��k`��"�fy1l%`{&�T���(M |8�iԤs@5Y��/r��B䉆<<5b�Z)j�q�N�L%�B�	�K��_a@���(=]zW�'��	�E�5��B��=̖��'f�(��B䉳
B�Pq��+�tT��B&cS�B�	)tjZɩc�ѣ8��dp���B��� �qC��CZTҷ��>08�B�	�4!��(�A�2�:���j�!4FtB�I{^5A��[�V��#��O<�C�I�{~���sX.Oإ1S,B䉁�� �t�ƓSe�U�Ҁ�0u8C�	+[Vb�;Q�X�o$V��3��66�XB䉫7:��A���bR�3A.��L4B�I�{��8�Ѻh�={�拚20B�I's�D�fÚ4N_�${���F��C䉩pf��q��|8bL��F�VÒB�	,I���&c$(p�G�
.�8��D#ʓM�z�B�'jM�)�gĖDW�nr(<�a'�!�Rq !�;{��<���w�<A�Oqo���v$�:L\�e��IIw�<1@ ��$�4MPQ!5���#��~!�䏎����^	����Z�B9!��x)n�+�ӧ'hbiqp�/~,!�d�=�0��|����Ť�)�!�d��k����P�D�#ˈ)��"�1�!�$�c�|�b��?�Z�2��?t�!�$@��:��@��;�4r��
l!��"%b���f۟���C���K
!�E9�� A ;�|��ƈ!򄂬��`��Èm��H�"�"葞܅�)� �	����"���˄h��d �h%"O0
t虞A�Rm�T�ŐRH�	"O �Ф)Ґ\%Ҍ
��y,��	�"O�	��	�b=�����i$��6"OY��-��te�����ݚ�"O����E.=J��Eˇ\*��"O� z�N���N4��-�����"O�]9�@�~�tQB�i�{��E��"O:�1�Ú���j�JHfTę!"O���HϮ`Q���� bx�3v"O1�CMW�1d�S�h�L�tUD"O��9BI�6�<ĭ�X���sd"O$�*᫉�]��XiU� n`��p"OꬠӨJhpEe�H�4���"O �S�O�	}qH�*Vd�@���A�"O䰑��Zor50Cɏ��fAV"O�1��l -xxX@ f�EWE�6"O>�%��osA3�W�<��C!"O��"�	Qf� �6��
63�� #"O ̱1G�!
R�G^�=Ş��S"Ox1�!X c���_�f��4���yr��o*ʙ &hZ�/���A�[��yҨ�x-�D�$t[�-�2@$�y2�Ҥa��r��
p~�0���8�y"ܝ,/�Ȫ"�C�vj��8ǭW=�yB�_~)���NԍxD��� W��y��Z?)�/�"�$��k��y�'������H���)���y2���P����)�B+@�+E�Q1�yr�-�xYQ�*�8@��IB�'��y"͛�%�H�ħQ 8.��8ZZJC䉓7h\�I*�B� �zC�H�KC�	2^@L����4qy���F��1;$B�	,}9`.�;DB�85���>�VB����i0�$^)���V��A�B�ɭYv�d+p-U(��u��U��B�ɋt#T협-")��,�aj�2H!򄀆Z9>A�ϓ�<x�g&�.hD!��	���Y�gF�~N�1�d�5a�!�U��tm�&ib5q���Gv!�$��Su��hT"��5wTh13��b@!��(]�P�T�N�^�t���fR,0!�D�l��jfhҰ��hTO�eH!�$�T�b��`&CF�"�J���+P!��:*f.��ς'c��a9�ٓ*H!� �� 
��T��(�`�B�=S!���WD���h��|��\ƃY?9�!�$�q��e1��&(@^p�X�"O`�F$U�B���������p�"O,�5G'y���f/L�1��|95"O�i�0��4��>�|kҬ�BA!򄇛a�UK3料(�H�%L�
|!�dP�X�D����ˊ�D�SP-X)~!���xV=���C4QZD�c+�8u�!�d��Mcޔ��kS�N��Q��#�!�I�i�����<]&����(|!�d~�C�U�K��p��M*V���H�"O^\���Ne��I a���l�B"O�����v.���� Q'�x(�f*Op����#,l������>k�7"Ox�X6I�&��P#Dϋ'�"�A%"O9��D�pA�Z��!`�jt�F"O�"���.�|,��X�F�<��$"Of��0�Q�� �I{�虂!!D�� h���Z[�x�E���4�`"O���c�R�'*X3E���Or��"O�x�tl�f��e�Teу>Q�(��"O4��De����r�cĦ8�tE��"OPQE,
.C�lA���A�b,�0"O��+4A�&lq�����5%�T1w"O��@�H"6�$��ì�-�r�"O���m��MPZ0��H�
�B P�"OjQHd��"�.�y�$ݳ]��%�A"O\q+���b$���#JE ��Q�"O4h��ʓ"�^q���B�"<b�"O|E3EbK�1B<�#(�>Vא�`�"O�U���ލC���G΂s��v"O��2�x��lp5�_�x���"O(�����L��'�����8�"O��)a�o>����[v,�ZW"O����+���}���0lL���"O*�s+P>���+&uP9��"O���/��2�<��I.T�Bm	�"O��Z6O]�da���e(��8��5x�"O����K�7(rT�@p@�*.�F�j3"OVC�A��2'T��6`�Odz��"O�(�0��8?^hmRVз8I8hSq"O�iB�б�����L�AЌ\Iu"Ò �b��6v����>fD �F"OR��q��e��ŒvΑ�Jq�"OZ�&m�W���p.�g�r�Q"O��b���/S���ae�[����'"OX�K1�"�l҆J�q��q�"O,e�'#�;3�h�rèJ�0vJ|1�"O�)!��Q��0�c��o.��"O|�J��ї�,X��QQ��!@Q"Oh� ��XF8d`�O���q��"OL)����y�F���@��ֵ�4"O��1�H	\zy����C��A�"O(�	�J��z .�Q"/N,cؔ�I�"OB�(�[))�]R��H��D�*O���@-�$X;h��'�e��@P�'lf-����8��#�h��YG����'���e)0jΪ�0�΄�QW����'blգ5�[�몉	���:�=z�'�`��`�î ��x��i�9V����'� �c4jO�J�[1�Y���x��'}��D  ����eT�Q~�p�'L
�Q�M7q���(�)L���-�'�01�%¼Q�V�z�!��CQ�UY�'��`��:�ɩ��ǅ8���J�'����i҃\��x��1hq3�'��DZ� �+t��Y�-�/YF��'5����
�� :S��6C݊8��'jv�nB.=��� �̒.oy�X��'�I����?�&Ts�o��2�p��'��� 6je[�Qr��>1W�1��'����n�\t2�֪Z;$FJH��'9�\@�j@�/7�����A�����'�:-��*�"g:��ԃXb(T��'�5��� �v*�<y�"�!v�C�<I���$/b�s�jź/i�l��E�<4	ӝ�0��`!_(��RAm	j�<����g��ȑ-˵\���be�]�<�# Ӫo��p�ɀ�:�B �r�W�<�&��5eX��o�/m�Ĉ{�{�<!7/�o��:w���:�P��{�<����H��bˍS>��7�{�<� �+"���1��H'c�=c�����"O��
2.ԑ�&x��B�qT@ZC"OZY�@��kH��P�8[X���"OBK6��2����b��"@���D"O�Fꨄ�g�G>+(ܥj5iP�p�!���1u6~$҅�߹Zؐcӧʁq�!�D�v���e"�t ,0d�L�h1!���A9,`��!ώ��LCT��Q!�$�58��C���?��RR�F�u!򤉢ff�QR񯎆L� �X��8j!�$	 7������?���;�D��=y!��u��\q e	�8� 8�p�P�E�!�B�Dq�ikΔ.�n�	�����!�D�q.�Ts-1�i��@T <�!��I����
�g��B"��*�!��|ab�B�E�B�b� �!�D�wj��0��G (��\�aӑn�!�.�,���-��v�`����^��!�K�c1|��Ҥ��P�֡J٤-�B�	0^I�Ȃ�H��Px�ٔ��YB�B�I"�ܫ��� {&q�怟�2�rB�aZ������\6�(Dƀ�ǜC�	r;@L �)ŗJ��`�V�:*vC�	->��JK����PlC�I�v��%���T߄,S�"��|6�C�ɈkuH����3vL�s��:��C��~�����_�&�z%[R!@MK�C䉅>����#J����B����B� J�,�R�"W1*�X�@+�#><fC�	��ѐG���|�bǥ��q�rC�9%4P��@�W�`7l+Bh���*B�	�VE@�2��:H�d����B�	'\�P�cUH
)k|�3��X��B�/#X�D��"M�$	��G'+ؤB�Ɇ
fp�����3T��|aq�Z�CDHC�	vB���&	�	hӓ֑lƂC䉞^�rPj+Ӟ~𠌡�U�.F>B�	�`#��
i����NLˈ���'�2hQ��i����G��5_��	�'��T�f�\�R=��n�/F���P	�'��2��i2��F'ԍ�ָ��'�6\Z���4��1���hj	�'�h �G8���Bм~�8	�'yDɩq$�%ox�Y3$V����'YP$s� �9W�|�:�ݺ~�z-y�'w��t$�M�ꘒ1+�c� S�'�`�g*٬B���� N3r��h��'6v �IU�bm�D��k���
�'�T�:w���4\j��\�h8JA��' (����%(tAxF�$vL09�'c����9-R�:1 E ���'$����L�lqqՋ��xzK�'�� g�#r����
w��P�'�T���% ���J����6�3�'�vHʤ�7p⤌�#`�� �L}��'�N��5J��A�rQ!���k
�'������7L����(O#Y�2�)
�'����мl�t��q���}�\��']�����V8"
L%i2Ϛ�w�4D����x��ҳ�G�!��x1gF��y��&D�I�׎ؘ����fւ�y�	 ������6.�zQ�m��ybd��1�|��'Ž7vԓV�G��ybE��n�<E��m×Vz%і���y
� <Ac3�V2D��Y��E9Ѭ���"O�X�3�T&oô�34��a�4QK�"O�-K!ȓ�=d����F]�E�Bg"O�T���*H/�L�#���j�"OUS&�n�+��d�>�S"O\ys%�ЈY��ىb���F��<�G"O�
�J�a�P�%rl����"O��3pC��q\IK�@H<B��y"O�0�Ҧƭ�N��jH�H���:�"O�����@h�=���Us���"O 1eRI�٫%Aی[�ᩒ"O|)p�E&!z� ;t@QS"�E"O\���ʎ�:�
����&S,*R"OplY�n�8k��	�UfL�cK���f"OЕh��RDUh�RŊ�#����"O�M��mѸv`�m�䎗M�<H�S"Oh�w�ڳ4H���A�0X��L�"OF��̿Wrv�A���R�;"Or#Q*)Z�P@f\s�V��"O� ��R! �e����zq"O�����2@���#Θ�S�8���"O��9S��@bT���K�Q�Z��"O$�Hv`�)S��T#���	�L,p"Oڴ��B��/7Z�,�2m����"O�T{0�9�h@���ƖW^��g"O��V�2jV,ѓQk�A&� r"O��PcD
G��� 툾P�,j"O�i�#a�w<�,���J?4M��c"O΀��d3g����!@���L��"O��+�F��T���r�ܞS�Ԑ1�"O��� i�,�P�� @<;���qt"O~<�@�V<ft��*!��Ȱ"O��lNE���Ѵ� �c���"O�u���} 8��&=����"OD5��:=���FƓx��L"Oܝ�q�[�"�X����>U><�S"O�A8�璐v��������t��a"O�B��Ŭ0�A�'K�<�@�"O:��1������0;�n�"Oh,�)���-�<�t\�3"O����,�x��ѡC^�h��A
�"O�D����,4���ҡߨcz�(AB"O���V��.�n�K��z]x�"O�1���6�(� �J�2���"OzL���qk����%{�b  �"O~ 9��Y�r�Ȓ�&�<��`"OPM ��F�P��eE���<��"O��[!EճPSn҄D�%h�\��6"OrqH�e�2"Vأg�	�z�.�HP"O�$��45�X���V�gS.��t"O��x�iG�T0��?0���b"O����/i"� �`��0�İ�"OYX��Y
�|��H�s���F"O�2%�.g��10Wa�F�>�V"OiB�.�PqvE�/xK�rd��"OT��rlֱ���S�R;���S"O�$���Ҩn��iQ˕:]�H�3w"O6%(]>6o���/�؆"O��
%c� xhņ"!���"O:�W��(�#`$M�Q��P�"OV}J�	S+.�Ƅ�~���k�"O��RC}��� ��v0K�"O�i5鑚j�p����C+!�!�"O��B���y�(�"�Bm! F�g_!�� "�9w� �31|9��fX#QZ��%"Odݳq��xx�=��c�;���"O��s6�I�u��u1"�&=��B�"O��K��-)|���ʹs
�ˆ"O(�c��./�LRG�'e�i�D"O����4^z$(��ņx�`��"O�u:���_��!���F1m�L�"O2�I���p�x�1S�� m���"O ���:;$!葎�`�����"Ovt�AH�u�֭а�G:P�����"O�����0{�(h��_3F�j)Yv"O���E�	;r}��\w��3"O@��Fb��E���c)�_��""O���$��,_2� �"�Y5n�`"O�Ԑ�ϙ�k�ɱ�N�B2\1""O�xc�!��<�D)�d���s�"OBA[qǂt��@{�!��(�ā'"O$���C�F�����?�j���"OL-�b@of � �.)�[�"O�eI���B���k�fT2��A�b!�$?*�Pհ���QшQ�'�/v!�Z���V� X��2E���e�!�D�!Bc�= ��0*d��/ߖ�!�T���)#oÇ
|�r �T�!�DP}1j�:�&���6�S�$7H�!��ӏ�N�K�l@>I�p�@�/o!���
��$��"sHt|�4oN�a!�dFj^�"��J�C*ԥ��Z4�!�D�dĈa���:K ̄*FF�o�!�$X�T���p�d=Lx���UG!M}!�D�>�P! ��Sk���W,�!�:C�@�Pf�%DQ�¢z�!�<�� tL3������+Z�!�dF2D��h�$��/:�!�d�b�p���N�RgKٯ�!�ę�}�a��1H�M���Z�n�!���0
���)H	&�d��	ڌ|�!��Hsw����	]?���hZJ�!��5�RD1�ŀ�K�.���FX��!򤔓X�)J���wӠ�� �X�!��>N�7�D2�l,C#�d!��e����C�Vr�(ҝX!�$�)�^��g� j�P��QV!�D� ��4ؔKY#6����T�m?!�dسS���Z'|��6N��&�!�DĜB"b����>?�0�7�!��]�N��+Cƌ��x��uH�+Mk!��ݸ}V&P��aĮ �Y���;!�d�5|y��J��N�<��Xr�&.�!�d J��ڤ��.e�������!�$$Y��K��܇^~�TӅKU�{�!�Y�O��u!�Qqv9ZMT&o!򤙺IL`�[�O\I�xH�Ϥi�!�Ę?a&0,X�`�'qC��2U�
�y!�$S>&ɜUk�-��r,��@U�C�z�!򤊟/�I���42�P+v��	�!�Dύ7�.5pO@3*h���bV(CR!�@@1�U�9^��Wb_)�!򤏁�bLS�a��mX����O�0�!򤓂+/$���ĉeMVD��	~!�d��X$�	L2La�4��#ay!�$ڛ!%���cŨH ��Q��[""^!�$Q$[�2���2��c��eO!�d%KʕK���-��kBu�!�� �%�"��^�&ˢk��n�4��"O�X!���F�䈲i��i��t��"Od@+I�87b0�f���,~��u"O���S	�Iov�'��Pi�"O�#u��PFĹ����7Wܲ|Ӆ"Oʙ���1kUd8�$�/� ��b"O��q.RP��B#�P�s� �zu"Ot�@PKK6d�b�
��%gz&EC"O��ֻN �Z"�_eL�c"O�-,��Zdz��ߛw�Q��"OPa���@�K?��g�E�.��`�"O<�x@��$��Yi҈ K�\�ɢ"O����_�pۜ�X�)�2��U�"O��vƳy�(L`�ꏵr��23"O���J]��I+��҄8�x�:C"O��Y���y�L�
a��a�T�XC"Ob8p��1bm.�`���S�h�"O��Jf��>�uYR���T&l�a"O t�椚b�*�*� �2o�eʧ"O�QS��8C����*�00�"O�u1��٬�����D9'�tH�"Oր�`"UR�܃6c]�c�<4��"O��� �*�L`��"-� ܡ�"O�P�&D�͔pS��0��5je"O�L;��DM�P�
̇{���"OH��� �+#�09�T �~�2�Qv"Ov�)PG�kr`����
B/�lZG"O`� �J�n] c�	L�h[U"Ot�ˀ�R=d�xсb��=/�Yۧ"Of�"⓶k�*#Z����"Oz4���Hl ��4,�+g׼�;�"O�l�	Ғ&�hp�c*ĥ�5!S"OPIK���~."�s�	��Y��ڥ"Oe���;+���q�	�)��x�p"O"}@���R�n-��扅n�t��"O�M�F�x��Š��I�*�����"ODEk�AF�N�k�	�}0��Ѐ"O �p�i�<"m�,�H�z�T���"O����ٺrz&�Bu�U�3h�Z�"O��ـ�F�GN$��E��8UJ��"O
���/ԎO]B� ��0E��y�"O��2tE	x��VJӗ����"O�X`I�[皼yr��m�
��"O>1ʆH.�Ь؄�7�ܙ�@"O�P˒�K8"QPHS���'z	"q@"O��
Dڀf������ݤt48x�"OH��S9�x�c���k�0إ"O�Ի,�~�2� G�P5-R���"O\Y��X�zm�$Q�䕦W�yr�"OB����m���s#�a��\��"O6�;vL��,-Qe�
��%��"O<%��,Z:�|l�Aa[��&���"O|�(f��Lz�`�c`F�,���v"O�yD�
�r~���W�ޕfW��"Oļ�Df� z˲�2�(E�B�"v"O.yca�������],Ij���"O��sEY�#�b��(E�O 0x�"O̼iTH�O� �au�d��QP"Oxl�%��^�>y�
��D���D"O�H��(��6�S���>M�d�:"O�}��śQ�8��	��8Xj�"O�C#'�xv���W�qȂȹ�"On��%�,U�f�r�ͅb���"O0$[aOD�]��b�ЉQ8`�ɡ"O� ��1b��N��(����9-U�0"O����:kJ>���
�u,,�P"O��yV���a{.I�� ^�ԙq"O�UۅR�D!�F�R����a"O�k���;(Iy�'Ҟ���"O�|	��Ԋi�p��L�=� �`p"O�ī��W;:Jt�s��"p
�B"OV��֪���Y�qa�2VV�9CR"O�����]���:qa��pD4��"O�]�#�,i����ȿ.�@�*O�a!��Î[�֩oF	Z��
�']�4�5��8���q��7�ֹ�
�'�r�!C)E��A�w�*l�
�'��bɑݠ�b7B�$~�xx�'�)07bӒE��"��P�l
�-3�'�9EM.ol=��J+f!�E��'h�AT�+Ҟ�cgO1^L8Y��'3z B�
�v��٣��=U��y��'�30�&G���hɻI�`|p�'Ab��&HP���vJ�x���'�t�%'�F�n��5��"KL`�'�H�1�ԁ\`d!V�^�}��@�'/&x�#�	�lVZU��J%r��'��c%�+�buI���<㔁i
�'G��c���R�VDY�� ����'�XIb���7uFQqBkD�=���s�'#2S��G�.<����dȂ(�����'#�=�v���*b!�GkP�v�i+�'I�:E-°h��١"S��
 	���|2�ӴZyx��<�*�êB���C��9;�Ƞ)�i�3Zz�U�� 1ΖC䉳t����.�#! < W#�~pC�IZ��`��"�NE�	��8��C�	�w��� �@�`
�p B�|��C�0,���T� � �9�̖9�0C�I�gF�Tr����1��B��߆��=�.O�#|���2�� Y#E��C(�� aCH�<I#�Y+� )*�ݛw�xTZ���<Y%&ƋF�Hy�fiJ�/,I"D�w�<	%CFT=&-�TL�Y�j�yCM�l�<�'�d=�e��V�"�0��&��e�<��[�C��$ڦ�B�E%��x/�a�<�v�O!@Lr�p�2l�8vJGh�'�?�;G�#a�z�Qlr	C�H�"S�!�D��fD�����/�|A���ױ9�!���>M���R�Ȣ5rbФ\|o!�	�F�@0�A��P�$��Q�Ԩ9y!�[�,���k��	H�Fᳵ�"R�!��;E�.\���݃n�� B����O�!�DT��x]ie�H,d����2f�c�!�ԡ��y�wlˮ��xA�
&�!�Ĉ�y���עK�P���<g�!�$� at�%�c�I�}ȵ�^6M<!�䊬&*Xm���;D���RPA��NX!��V�"�Pd�L�Bറc��C �!򄌹�H�k�숋/p{�I�*�!�Dƀd[�=��Qf�G���Py�k��5S�I����jq[��.�y�	� ���F���D��F�U;�y���6+�fa2'h��u0�D�"� �yRH½����׉�o�`����ݝ�yZIeܹ�e�*\pT0���e�(C�	�3|x�_9&p��F^�`I�DK�'U�I��.�4��ͻ�,�,��(���� X�MJ =�z�ѦS���"O X��4vzH������Pc7"OX����u�^Ti2�ȁyt�D� "O��S`̷\�rMX�����{�"Odib��1 W�DR@ �%Jܴ�k"O|�;�B�Hl����$:���xq"O�P��JΉT�8)�ӈ[
�8`�"OkC�ʺ,r�ж)=�ze�"OM��@�: x@��`IV�b�T���"O���� �>s\�����V�S�"OL!c�`�+B6L5�2��%Bx,d�"Oy2 -՛\�������K Hsv"OX!�����B��Z�I��}3Z}PT"O���@��M��Q�&T�n+(�A"O�D�$�#�>�R/ߏ. Ĥ��"OB�9#�Bsu��%̏�,��0�"O�`����Oڀ�3ƪ+!�@t�""O�@�7� @x:�����m��"Ot��C���P�� b�Z:�9j�"O�;g�ܕ_%�|��܄3�����"O��@��.&ܲ8p��֘ dj�3�"O@tk �יT�}�6�K�2N����"ODEP��5,�.U�O@�gB ��"O���s���X1f����J�=$�B�':XC��n�`A�.�4��P�'}D�����-j��l@��<'���s	�'�4�(��k��L:�E�!�|4�	�'"����Ӧ�Ze)[�����	�'+t}���^�4�=���(Z;�<��'y�������?\>�S�C�d�Lys	�'H��$�*�"�k#�O�&��_\�<�-�(Q�r����	�2���C�X�<	Q��|Q^`2����C�P�:�.ZO�<��䈮{,��a���"󮄒ІN�<I"ձ=F����5� ��1�K�<A��[���]al��wn�M����A�<!n� *v����!>�I!�HI�<!��<=� ���O�������M�<�6"�u]�l�`�� �xӰ!�F�<)��D�q�6Y��D�.�@�0o�@�<I�G��Xھ=�di&-Df�zp��V�<I1	�	`�^�����0p��ċMSh<!Р�{-���$��;JQ�j�%�hO���i).	���d*)E�BQxb�Ӌl!�d:9�"gχ��E�q��je!��
`g��x�ɝ�TȞ<��� �>x!���`(̉�3,H����'�F!���0��h�O�?�~�h�Ǐ�!�<PS�Qa�ą8C^�`���+!�dB�tF>�R��0.�<��K!�D ���!婀�~?����%_!�!�ҟB~r�
�`O�L�CDA�i�!��Ђ&�h�fNK�m��c�' �!��S��Vh߼mz*Ё D)�!�+�\��#��*x�x��iT!Y�!�$L �Ƚ��a�T� ��g&M#S�!�qN�3Ac�2� ȩT��U�!�O'�0I#V*ʹg�ܽrA��!�֋B_ =��m�3VK(�EA�:�!�V�B�B$��aοG��0����bM!�)k��	���>.��cp��!���,�� �.| �/�
k4!�dR�+�8A�ȎLx�!�S.ػ��T��"�i�j̝Y)�M�3��29:B�)� �qC1�%&e���pj�>��m��"O���G�-V�$�#&k��e���U"O<�9�(��9���#�L��%�8t�`"O��*2��!M�qᇥ-�QD*OhIΪ	�@Jȕ�q���'�f��R��3x��0`чܐxal9�ϓ�O����Stf-
uo@�mz�d�\�H�	t�S�$��x����>4�mB�[T�؀��5D�$83
��0Py�S#��xC�Y���>D�$����w`@w�߾o���Tb'D�P��%�M�-���R6k$��r��&D�@�Gٮ@LiIf^+ =L���8D�p�G� b"�j�\�e��|+�	,D��8��߇5�&��7\�",����O���d4?�IQ�J�b� ��3Rp^��%bIR�<!Ə[��P�g�2n�9b���P�<��P�Y?愚p�&X�L(R`�[I�<�0)�H�cG�� r~űJG�<�M�\I�I�� �P!�\�<q�d�<�Pp��@�c� ��`BWC��l͓?���5�Z7v\�K��F�CAX�'���i>5�'�Ju���úQ�6����͎)�<9�'F��
C��|�Z	�b��,{,�`�'�&D9��Z�5A�i�,+��x��'XZe�#�B=p�  V,
�(�k�'�xL�i]������@�����'����[''eDP1���,\T��Y�'�N,S�ȴf6�S4��V��Z���0���R��Eh�rTh�����"Oܑ#�lق;��5��-Z�r�q\�@�'���c�O��D`��ގtӊ��eM9��x�'UM�3�,t��r�I���0Y�'~���U�-�LX���{�1�'��V��:
�Y8RFB�	�0Q`�'&�X��#_ 
Q1R�7 ���'�՘&���Ĺ�u��
�'U*׈݆T�q��@�m�ڥ
�'���u��)ZM`���k?F� 
�'�lh��خlt�p�%vH
�'�Tt#�]�)z��B��8@Q�@q�'Ǻ)�4�Zwf4���a�M��h(�'z�( �ة�	qA�B���'b��妒�)Q�ۑ�� H��P�'7�w�ԼT9�@;��<v$r�+O�˓��S�O�t÷`�|o ��$I<Z�D8��'�
�1��?�h �@��a�RJ�'t��i$/��j�M�4�E�QON�s
�'�h��o�9k���P�Q
N�~����yB��B1�
0a�����ĥШ�y�+��U�K��>�mh�J�k#B�ɏw���bG��%���A�	��D��C�+@K�%۔�BPJ�1p�㍃u��B䉨k��{�'C9a�����F |�B�ɱv/�;��n�*-��N۠] �C�� r�\�'����XQ��ؒe�rC��Mtt}����4J61r�՟��g�	{���4Ȃ�"� x	��A��u��yB� !��d
��}b������D�<)*O�"~3"ʿdY`Y�M׻(� �#a�P�<Qr.VQ����%�7E$H�ENM�<q4m׵=��%2rŞ2h�.�S��m�<9֢�=e�$h�@M��ͫ�,�M�<�2�X�01��	�NЯ(��{ak�Ky2�')ўd�<	f+΢!��X#a�]��#5�]�<� n���P�y�v�bk΂~��=���V�h���Ց�ĭ��
SN�n����,D�h0�N:c����V�OnWdi
�F8D���7��w�P���IB�@�A5D��Zcjӯ{5>�C����5,j�@%E3D���R朶� =j@�R�q�8hQE�)�D�<��]`h�+\<=|fq��!j�T��ȓJ@�YQTAŠ�h��4�K�iPD��H����8]9�8�K&|�eð��&"?\ņȓX>`�2e]��K�B&G�`��@T�X�_�U��+�C֪�Їȓ&k�!�!ÅZ��x�'%+s<���I�'���RT%_	B��)hġ�O]�� J>���D5?����1eX ��3��/$l<R��@�<�'�JY'i[�-_������Łe���?qÓf��A���ݴ[A�8u%QY��ȓ.M�H�L�_IM�i׿p�ʄ�ȓvZ�,���SҘ�Y��ڄQ�1�ȓ#����.�(ޑQ�?)~��`�R��Ʀm�-1��X�s���ȓ�
U*w'��q���Z0�ن�P^ޔ�Vd�Q�=�g
J�:��Ն�HBnm�E�S4;Ĉ��R�����ȓ\��Hu�T����K�jԳ&K�x�ȓ�.]@b.�X��t[�C�1zf��ȓ3z�0�Ҧ
���eD�+~x�A��K���Y C�o�]�PC�"8Nx(��{kX�� o�&?��8y���'6���ȓ�,d
��Z��J����j9��B�F`�/ ���&�͎��ȓ#�y0�'5��L�G�
? X���Y��T��$�'�T�Y@CM�<Xt��_C���"V�)p`����/*0�y�ȓ+�4��˖�Z>��`�(��J�І�G�':�M�� �p�E"�+�4��g"O`0v�
�>�yg��Q��E�"On@���'m&�ɳ��׽7J����"Oz`�@
I!^���J1c��@�"O:��� �8q��H�f$�3G�d�s@"O��Ճ6`�^x9W#߹.Ԡ�O`H�
R.�.Lq���2]�b#�6��0|�� ��^w��W ��w&���m�<a�&_6�H�n<>ٔ���P��W��C���;h.t	d��
jjl��>D��&l^�b!�)���Ũ%S�@�D1D��Z/�V`����G���4�u�+D�C���g�(�	G���o��T�$D�Li$FU���0Á�=(R�[U7D��p���8%�I�2Οz�]���/D�h�����r�^x� ��*rQ �za�<	�r��l�'�A�	��q���yٶ���&�&dyW�!J0HY0cW�$8�܄�o1�}�v�ʖM��%�@�ٍ$�5�ȓ{�A���@�Uj�SaD5b0p��ȓ0ߔ)��-@�I���]���c�X�9�hU��`���]�HC��2r�\��"U;5�AwG�0�%�ȓ/��C��;}��EɖB'�L���
������F�UQ��R�B�����-Q8��L���JG/ޠ-sTa��u���$n����e�v�^�9��Ȇ�	��tS�i�PNքq�	V(I��s6�����B���� �Ҡa7����$Μ�Hf�D ����A�C��L��S�? A��db��RCo�H�S6"O���jp�j�� H�d�x�"O\�#R#�)��13E>LʘuP"O����C8S�,��!L��jM3
�'@�Xg,�0K�j�n��X9(X��'�\���e^�H�����W�H�*��ݖP:2 x�ӆ hb���b�!��ʾf�z�U�r�Z�V#&�!�$��}���ÓJ���.�4!���*3���2"�W}���Ђ�H���
X%1��@�d�3����y@
	������9sXʥ��2�PyҪ�:Ah� ����qDꡊu�[c��,��ryrd�� d}�v�B>o�ByZ�)]$�!��(x$YYD� n� ��.�l�!�A*Ln�y`�	U'PQ ��U�2�!�PJ�����,Pr�k1iھ_�!�D_"|�j��d�D�E�̜���Ƃ �!�S��z`�`*"լL⣧�~)!�d�
�����c��8�p��H�����5�g?QU�E T\K���/�����h�'%ɧ��(˂D�T�hKeKǥ36�a �#D��I�[�	�R�:�D~B�¢+D��a���I���h�/�{�XhS3�$D���tA��I[��i�%/��A�PJ/D��r���b}�2��p������:D��E�������88tU8H;D�@�C�&\��4 e��lDN1�խ+D����V�~	i ��c�.}��*&D��1c��K�҉��IS =�6���$D��W%X�3P�8��аZ�])��/D�0�fD(@d�
F.�d��S�&-D�[�a/p��� @(��fx�g�9��� ��\�I{y2bՕB4R�ဈ�VU�e��EU�.!�$ݳ=��T+5�Nv62���d(!�̰�4���ˋ1GGd88�J$�!�$�ef�)3C��\� ��D2|U!���?t�����~�2����-PI!�DAX�=��U�I�ԡ	��ƴ|,!�Pd<���E
�)�ҽ:��5���)�,O��	1��Qs���E�з��)q�B�� r��5�Ci�k�Hd�D���=t��O:��7LOΐ#�)_06�����>d���"OH��cdŲS\�8QM�O5�x%"O�d� ��,����v��0u.l���"O
]P&%�&��d'�nq�"OE�%^�8h4T��h�3\����d�'=�}~�G��N�l�`n�E���:D.��yҬ˼02X��P4af�m�Ȇ����O��D0LO��8�n<G��q��4=ւdA�"O���g�7:�2@��Ǎ9����"O
��,+�������<�����"O���&��*'n*�JfF�pk�M8�"O8�	�?��!�e-([(�h`"O��í�G� �&�ky����"O<TPE�ًe��D�"7wx"��4"OdAb��V�{P�r��[.
�2��"O���"s76��`&�!/��8�"O�4�Df��g|���ϕ35�jX�g"OF�@�+�:k����1��a8� h"O:lZD���e��p�b����M;�"O�3�Gϛ �Acο+�B��"O����� ���6�U,9���"O�-Ct"U6H�`� Pvm "O� ��� �E!]��mj����xhej�"Oj��@-������*�Q��1�q"O]�@cTΨ��t
wO !�%"OP 23&ɳ=%��Z�j�5����&"O A
�܁p10�gC�9/���U"O$9У�� ���b�2tlT""O����ꚋ{���!wU�Y���t"ON�kw�Řvi\�A�e�Rn��U"ONY�m�o�iEdЊ@@����"Ov�dA�,{�#˰4�D���"Oa�b�&,�<xۆKZ�j}Y"O��)�zh���'�-���"O
�`OM�>Q�m#0��`c� rg"O� �hN�&��y@�@����"O\���ծNP��Q�����HD"O�,k�h��X(�����5RPX��"O�lC�L��V�f���D��{P�QA"OhxctL�I����$�:?�	B�"O��ɅMG
pv� �&♋Y9��W"O��Rr�O�$��.D� �""O��S�"< h�C��?+<��"O��{�#�2��*��9m65�4"ODȰ	X$h� ���'ە��9�"O��)1�N�[s�m��G8V�:I�"O�TI��M�~G�a����8O�"e5"OThȖ��h�X]�S���K��]��"O$��� Z�	v� s@�L'h�8�jG"O�1����!6����	��B��"O�M�c
m�Ėu�$�X�"O^��BH� u,��k�G�ă�"O����a +Q��",M��Ae"O�%�1�ơyE�L8K�TR�"ODm���3J���U-��zIz��"O��c�L��N���L��81��÷"O�	0'H���~�"5l@�v)FQ{�"O���S��$t��F��6x�(�"O�\ԣ�_�(�Sʈ�y:�{�"O�p�I�3"�\�fc� s�XE��"O�2֪�=��p"�,�F�0��"O����W�~� x3�Ԁ
0$��"O�K���#^+���qD׾@�J,)"O8���)�-r��2�A\${���$-D����jE���`��	<�$qs�k*D��K��Θ8�(�!p� >��Ԉ��'D�4����
<��S�A�Tq�Q���%D���c��u-�9!%�٦;���@��"D��`�/E�mg�2��'#Vʲa!D��rw�E:6���ǮхX���to"D����?Q�N=���ϷY�0eۓ�5D��A2��?4��Z.Ы�G���!�$U*k��:���Rl\⒇��S�!�D�_�X��ڔpj�3�E��6�!�d�!xT�!�)ۼp�JE�w�J�a!�ա98�,y����`�Q��&�!�D�4p��Q�^u�i#Hޱx�!���R�0���:R4%bR�Q3�!򄂶@pĚ@a>HD�P禉��!��&=bX��` �5"�EzD��9H�!�Ĉ$@�\=��+�*T�QGMҞx�!���o����Ǩ�D��]j���
�!�DC�1i�� �ŀ���Q!�� 1�`�ƌ#����C�T�6Y!���0,"J	*ȑf���@}I!�Å|5:��D��O�]���^�!�� �!�F=�d����1�hl��"O����ȖqB�%�DgN�G�^��"O���L$#,���%� ���"O�	�j�Z'�pI��9wݮ�H�"O��K�)Vč�L�<��X[�"Ox���#əX�(h ��C�0Ә՛s"Ox<����i�lQ�S�A璍�"O6�Ie�2L�`)�@oȁ�`�1"OtԉW�G��i��Fv�q94"O�@�	$����Ċ1C�1"O@�p�䐖�f\�e�Ҷq/&Т�"O`�A��e:��d�$��Aa"O�)H�IF$$D�V�Ӌ��L*�"O^�Z��.9�����������V"O��*�U�U�&ӅO8�MX�"O�`��&_�pPM"��Y�����"OH��Ŏ9U�,p�-I��6���"OX��@ I��y*#A'�X�4"O i(0�۸D.�񰐪O�� @"OX�2��*넝J�N+`;�!��"O��Peܭu��J���8V`�"Ox@H&:�PYC��ԍI5`\��"O�,b�m��
<����%� ^0��V"O�Z`�Ä � ��G$��B�&�"OI+�-T�̱�s,�~�R�z�"O�,B����[��,V'OdBu"O������	Z(L��`�%[�p��"Oڄr�$5{���y��M��a��"O���c�-N�s���q8V��B"Ov4� �7Rv���
;�L��"O��qѣ�$z�9�®�)��D"O�1z��4~��31.^���"O�A0�k	R@�8ʲ��*�>�b�"O )p�ʎ�؅��I(a��h� "O:2ѥ�@�P�`���vC� V"O��sEN"?��q2�(QX@��"�"Of�Ja��%%�t��ٙ=@�y"O0��E���V	i��Y�zd�P�"O����b��U�`�R�M�q��[3"O>����5+*�#�N#x����"OJ��G G�]� �ʵ�E�H���"O��c��@�0C��0���"O~����=X ��@�ͭx�>�"O�,�N�)>{���B�hä�{�"O�y��aY�Ba���Z�	��C"O�5"g-b�*X�"�UQNy"O ��EUs�����,�
� �"OH\�	�>��p-Z)	}��I"O�)��ɇ#��H���Wt��#"O�LHf��A�&��3JBd9�ْF"O���"��2hr��Uh�"Mt�Z`"OJ�����	^��@�^) �l�"O&�ॅ�YPȘe&�4z)�Q�g"Ob����I�i-�������!�C�{�=Z�mT���C8 p!�D��67,��pE���b�����Py���?i����g� X4b���\��y���0V�RMK0�S�MZ�@ o��y�a���41�c�}�.$(P��yR�$��H�I;v<,<ɠ��y2�Z�'��q��-O̔i�P�ϋ�yҮ��H�c�k��x���Ҡ�y�n^�	x�E��c�,f,(�:�!U�y҃H( ⁻�,V6��xڲ�ҙ�y
� �=�kOG����F�}ENe�#"O�5�炟ui�lk��˱2*�`%"O���R��*�9�F��D0�=��"O�ꃪM%G��H�����9A"O�5 `�?R��]�@���
����"Ozk'`U�<N JQ	��"��"ON�B���ʷ!]��ܺ�"Or��ȝ4A���@a��L�x՛@"O����?g��)`D�ߋ̲��"O� �����T�R�`0 @�o����c"O����_�nٔI�ӬTj�P� �"O�р� 6�(���U��\�"Oj����
�kNu���:�����"Ol��%O�IJѱ��#��"Oڡ!E���-B�3�+!����r"O���`M�sb���g���1q��"OtPX&�F5Q�Ƚy�*�.i�,b�"O�U�LC�s�NԨ#j���N%��"O,Ad��b�$5��(~��y�"O���r-ΣI��Lcŧ�9H���f"O���#��&S�-8��R�x����g"Of���P�4V�0N����*O�K2Ȍ1�hH�Z7c�~8��'*�r���'���ؕ�P3�ҡ��'�8H���zRp%��t��'`*-��N
�	�x�����s&����'�5��ju~\�EΔ6���8�'��T��Ȍ0�ЊE�����'���adMQ�Oi��Dc��U�
�'?j0�4�v�8I)w��\����'�(�`vB֖��k�@�B���'>�(�7,�3�X�ՠ����D��'� �)�Ʉ�z�c��/R���0�'����Fg6�U�P�^W+P�h�'��j���	&0H�p�#҂_6Q�'�n1)�	��7>R�����]�2�a�'�f(X�+ƍEE��C�D2w����	�@ԝlM�5j� �+v�漅�(=Jp��k�5_�1�g�U�`��ȓQp~�X�g�T�E>N��ń�-�f�������ABD�|�ȓ�x]"��,��tY� �4��I��.�(T��8g���� �+BL��f����J�r�RE��G�S��ȓ�¬��A?LP4@Ao� "�Ƭ���<�{$�'�J9�M�3s�|��+��u3��!0���-658��ȓ(Z��Qe+�+ߴ���̥s�e�ȓB���p(S	l�����O��ȅȓ{�|�'GNI.^%j3��q�"D�ȓ���r�lPtA)��u����6��� 㐄u��(@� :��ȓp��!G�6T���բV�Ҙ�ȓ8�k��)b��
U%C0���ȓO�h��O�muf$[�T�K�Ɇ���(��
#p�2�z ��u��}�ȓ*s�5�4-�%w
u����x�y��9t<�RjӇ�����B�8kX�P�ȓ:V�m��OܛR��5��$N�
YV��ȓ4ml-� �60�*���F��0�D���Pޤ�1,F�n񌅠&ȍ+6=����>b�{��(ڠ�9��L�h��h��<� )����8݅�.�{Q"��PHRiR�e��8I��S�? ��d�J,�E�D�ӡ'�$YXT"O�C���r�,���&�d��}`"O8+�.�Et�9��l��m�"O����1vJ�2��Z�7�R��`"O��2��&��ri r>��"OL�R�*d�MRubZ��&"OF�h���7 ͐ԋ�E�
9kR"O��P���7Lö<C�!�S�hXR�"O�U��*��:��5�g�̷�`l!F"ObZ1DY�|�Q"E��r�B��`"OtJY��
C�Hg�e@�"O\�c�� �&�����ETF��"O�T�t��(	,ش��L�D*�9�"O�
G�O��0�ү�K&n�U"O|A�"?Q��RQ�V5��1"O
��P�N����YyT��w"O|A�
%���9�O)0�����B�O�~D�E���N�{��

7f(�	瓪ēb!�L��6gs�<@�
����ȓ3_̅�waR���)�JD:~f���.���ҟou�d9sOV�	�i�ȓ'��d� ��mT��Їb�><Մȓ�̱�a��L��iN���ȓi;�d;��)^u��ê(�����1x��`�<U+�hw(��y�d`��E[|}�p��F�,��)ŤJu���ȓ?�q�f�2=��ccK�$�D�ȓF���B��I�ڭ+�[=�N�ȓb�h$�����@0.i���5a^���b!�j��*U
�µJ�4
�:�ȓy)f}q�Zs�VIq���x|8�ȓ%O��z�ˋh'P�X@hIn�J��HY��ȢA�s��Bt%�/8��ȓ׼�@0�j���W�t��0��&b�`��6�tA�G�-i'&!�ȓ%��Q���:<>�x0eۓ.�t��ȓP���O�b�I!�]����ȓV��k�O�f���b�_�l�&��ȓX J���]�v����,U&ê���h#٩@�Ri�xB��1�p�ȓ�t����_^Z���,�M�б�ȓd�Rx "��,S��b�m�B
p��e�>�iQe	QD�Y�3��θ��GN�C��gS��j���&
8��ȓd\���aG_�e��Iw�X�(|z���b�b�pAݺ<$�	
J
]�j�ȓD1dp'�D�I�0��.� ��نȓ5v�9`���_�n\��cӅ3�^��XeV@�̉�~.�2�^N3����PL:�S�
=7�� 
öesF]�ȓ���3�مC��u��E�q�\݄�OC��B��فSڍP��lx`���4�Ơ#���	 H����ǝ
P؇ȓ�$y�f(ȫT�a���3i<ԇ��TEZd�Js_hh�����+�j`�ȓ1[�`9�#�rZ$s%'N�غ�ȓ'�
�*���(��*���!DȆȓZ]�H�u�O�| a�E���N�z�:!�(�T�1)Auv.0n�P(<1���>�"�(���$e��A���\�<9%�.l=�Ղ��J�;��(! �U�<@Ɛ�0��푁���3�P���Pi�<����#�q��԰P��8wK�^�<�soY�x{n�
�
4��� )B�<� ܬ)�AM�98m��+Iv�"O��*'�Q�ͨ�c���eӖYi�"OP�R�lG8����br�.��A"O� Kg��;�Б�!#�28*����"OHU��父W��ڃ��3mv�C�"O"�j�*���
�2�m%K�l�"O��Ye�(̈́�PG��&�e�`"OHq;���<�ܕ�熋KhB��"O^� �J��x�A�Ne[�a �"O����n_�G���P�O\�#A�E��"Ov)�(�b"���.3�5��"O�<9`�P3s:v{GN(|��� "O(�H�!��K� ��W�N�~���`D"O�tIbD��hx\�Y!�Fi#��cQ"O�h���)D��A��[#q��"O\��*K/�j��daCr����i���[�R�d�ҥ�=���f$�=�!��E:<�q��8�NA���Q�F{!�Ҙo[�*��O�����o��5�!�$ nl����Gr�Xz��q�!�& �x�Z�%��uю��v�KQ�!���(a��uCQ��Ȩ}bЌ�bt!��sVIaT�˜9�(t�f��Oc!�%���%<s�X����bH!����6���L^�����a�!�*ax��B�T&1[�y�©��*�!�d �96R,2C�4_FJ�Hׇ9�!��W�1Ƙacr�Ǆ9�M	�Fg!���Q�,��t��8MJ��F��60!�Ė�T���q���i�D���!�dR��
�"Eo���ص�
2�!�<i=z�Z�)$@x����[�T�!�$���A��i�uU��XW��:�!�$Z�O5�|җ��pp�UP�j\b�!��6��[��R�`✺S�8z�!��@|�Xe)��S�}�bƟc�!�C�% �i� �F�o�2�@C2�!�DQ7	BX����=��Y"0�?q!���e<ib�B��Ei�?!�ͺ��c#����s���dr!�d͇t`�]�����tP���J\!�B!D��Q�c��=>��Y!���q%:��!��'�8�`s�͋^!�D�Z� ���t�"�m�T,!�d���ptf����E�Ѧ�#>!�D�%IU�p����b�����㓿4�!�Dڬl�<���K���PrC:�!�$R�<ޞ%�4��9�RHrMF�n�!�$�D������Vh�] ӡ�5r!�d�&fcl�QL��Cbx���t�!�D5sj:%Ȳc�4���� �2o�!�$�9�Qit�E�4xF�Î�	o�!�D
�Otv�9`��aN�Dx���!��׿mx�� ��{����ˈ�P�!��4^�Bq�)*����F�Zx!��������˜3�T�!@��5@!򤄆B��D�#i�z�b��$�Ug6!���Mƚ���	P��-����n!��R/sF.�2��N�h�b԰�M�>4!�D�<%�(����C�8�q�a!�D��
1����@u��V!�䐍||H�hHKivh�(#�Ζz!�W)/�n�j�G�p�{e�B�d�!�D�8Z}�&&�%\PН�T�!�� 2x��A�65Ġ�wA��<��"O��R���N�|Mk��1n�Jh[�"O,L5S��h��ӃO�L�H�S"O��c�oČ�^�9va�.~��1"Oh\�@dL =�|%+�K�	���"OH�1,�&[�&���H��b�i!"O�-����0�9?oz��-	$[�!�d�3�)��Щ&aU8�kK$p!�DX=pRf���P�4�PMD�FE�!�dH9là�z�N-k�fts��ĉ2�!�KX��'ںw��<٧�.o�!��5�$�Kr��r�(�$!/>a!�ɩC�V���j��B)̱$H!�E.H�.��$�ץs���"g��:!�ċ�(�u��.��x�l("�ոJ�!�$��8v��x��>�b�q�J�*�!��
�y^�|!m��a,�*˔.�!�C�hAjA�ZyF��)���=Fq!��͔L*8AV
C���$�����6�!��4B
X���/ts 혲i.!���� #3g�f��LL�{:!�֩D(0�`��A�^����%QY4!�҈A�LR��Oܚ���=t?!�Dܛ:5<��tk�"|������	B!�͘%|d�0'щ"A�U��MQ!��#.Ɋ��"�H u��4�()���hT�eoм|��}:B����i��S��9C7kЍC�RL�C	r0���&��|���$`�����ڕ�ȓ������(#�cU��U��D�ȓ8t�yh�B�fH�p��s*�ȓ0	�hq"�F���ض�DCL`���(�G��6Eh�KLrl]�ȓ�px�.H�x�+r��c����G����}h􈓶�B�/��ȓ!��K����=sB@G\?.ZxQ��a8������vɹ������,�ȓ��ЛCg=��BN�:4L��F������Ut����Y�HW� ��T%,��τ�V�Z����2&f`���K쪼2ū=K).Pѡe�!� =ΓS��أ���X�(
�U��A6`���N��AP&{@��퉉=�> �4Ϩ2�0�*@�q,��$\�XH3B�8� B�	8��hF�`
��(b�ʇ.\$�!A���/��������~�`�ۧ,�a[�j�;%SȘ@Q\B�<a��H�9d٫�#ݶHtz������W�������|~'�����	1�2|���p��	T#9��C�	�0��ŉ��6��j�+
�~�@`Z��[C�1�Oa�6
�2`��e�,er (1��'e(��?����w����ɒ'"�^q��@�<ASd��S���0Ƨ��۲KIJ�D��N��?u83�,#b�5�T��f��Upm1D�lZl�50<NHI%�>^й�@,��.�����A~�@eF��@�R��ҤDe�!�$W@}nx!���+�b�֧O�$%2X�tm&4�Ă��)���&k��w��*O�@y�G'�ɯa)MqգH�ϴ�K��2�B�	��DP�F�{ʂ}���J�o����ӎ��I�s%RYQvl��O�8x�덢���r��H��\jsǇ.$�Phi��.����!��.����?2
,�fM;�HL`�&�3�'w�zb���H�{�%Bc4���)\L�p�'9��H�b�B������oN��wd��ax2�]�M �O�Q�Ծ~��y!I�E�G"O� \uRTfO�^�z%���,3�
��Ց��Rf��w�S�Og��� ƣ��� Ō��|���J�'1�ɡ�AN�M�ܸ���"'�$}:�y����%��yR%��jFxK��͢7��A�H�6�xrE�>h��Pdď�V����n�04(lUO�HJ�%�dǀ8�b
�gR�԰��'�V5V���8���PP�A8ȹ���/�!�DT�{'��B�CP�fr��� �&�F˓A�q���������85n�Vi���=8:az"���$��)2�Ӊ��{NXz.1O��cW�8<OPYkR�@C2Y�H�d�Y�e�$(�S����C?�<*#��'�<틐#��6��(3�O\�ЉS�(M�/K�r�j|r1�	M~Bj����'�v@���r2wg�	
�'��Q3O�)]�"�*QA�;�d��V��@2u�"�S��92NؔKX��n� Ԃ������ȓ6�$;�g3,���0.V�>�'�DKX�(��gM3@�2���5����e�.4���я�eh�QQ�i�� �:6kM���B�	����𪊎P�>�J¯^�S����dǨ_x5%���GR�c��	"Rb^������+D�p�;mT$2��W��� 5�ɫ\��U��J|�W(�.:��u`����4ӎap�P`�b�P:�J|Eh �$Ta�),JZ�5�҉P��QJ>��I�O��D	a'���f�ϧ�X�&)���8V��B�(��I[�XPc^|Qz���N�-��	4�M��:9��)�����pbe�L2�ի��M'�ԅ���9p�\A2R��:f��ɚ�& ��هDitY��O^�[c��)0܆89���$��T�f"Or���ƈ4s���	Rᙓ0�رr���f�L��'D*�0W,ˆ1�A����1&�ą�	�E.����7t�Q"�fL1�DX��o�b�aSg_e�$�#&�2��$���܂0��C**=)v��!M5Q�8	�H�	�D"��R�c�N�O|h�˂�]�e�H�c_&\���ܴuZ��9j��м��)ps�?��}̓?;�s0��5Ә�ۓ�\8h�~B�.R�wje�qaO�F�@{�͝u�<y�.�Q�@�T��O��Lcrf��%��$�O�.KZ��T銵$b<̖O��4�4.��ʦPI�i._�$ɲ7� �OA�U�� $���S/	8:��C�%�a*^�	b�83󎉨�c�8fY�H�;H�}r�	#��L��N\�NNtGyҠķ:L�iZ�a����T����LH|����xG� �����ɉB3\Y�U"O20���3?oN��4h�r>����� b:�,ۓ&�N��},cv��p���0u���}λ5d(9��5[�L�YViÄ4٘i�ȓ�;�FޚKb+w����dq��1@k���Ć0q�X(@O�|2�&ޛNn�0��#�6`l�ś ' :��I��9|O ����@�w��܂7Yz���%G�9C�C0`�z]�%��{@�a"�ߙ2f>��d�������^�:���/Z/��O�M���/���u��]Z9[`�0���L�H��P-Wԥ�K׆#�|C�ɤ!�Q���ZP����kN�8~lEP„o������*)����s�%'�I��(��vޭ�G�,��X�OY��l���8D�X�4-�c8�A�)L����V7I���C���o&��t�irr�iξg2�*�&"�	�k2H�R�L@+��8�k�0�2���N3r��19�	�9n>P���e��V��A㌹F9� ��S�	S�i"���82K��9LOI���%)�(�'��3�8����EE�0
N��gG�����.�)@$�/���K���X	ޙ�1�$e�Dd�ʉ��y��՞#䬄{4mY��t����
�V�	2.J:Cـղ@�֪�hHq��#E\c�ȼ���C�Ocv\�ֈЂb��y�X�<�7(��
���dm:�aҎ�x�f4�@��M�P����!�$�����mUx�L���ԠJ�G@h=y��nh���I&����I��h%�Y����']����¬�/P]x������OM�`��hJ���b�\�&�L�poQ?d`X��)3�	�j�0q:��I�1Z��a�!{��,��K�B\��cw%ĊY�� Z@NC�S7�q��c�<I��J%A��㥈U3/v�ի��Y�U��@"$�Y�Z�L��'���q�h
$C��'?��;"~J-�r	���,מ�T��m;�"O� ����m�+"N��%�37����Jޚ�L�"��BW�#Cʞ2���-Ŀ)'D�0d��)F��� DgL�\I��L���{�$OE��\�A-O蘉ыY�11��0��G�;��נ���%XcCZ�A;|��s�'i�a�.��@��,=��P��$� N��aC�/T��Y����Z|�h�D��5��}k�"�c�𤹖��Bڲ��"On�Y�J�hw�� G��#y��-+�F�t�l����s��$�g��!�d�y�
V���yר�#�Vi��'I(8�h��D�Z>�y2��y��P{�	��D��L���Se�űJH�w�j9b�kIRj�|�OF���D�d�1�|�yS�<Ȣ]��(Ǉ+�a}"��S��)g���{�z8 P��( ��U��̀Iy*�jǂ ���JU���2�K�2!�ѵ��9ǒ�K��,�3��JC!L	~D~yH���0%�<0�Om�	��� k��U���@�V�L��'j��HՄ��
�[g�)Ilx=@�'L,�ِ��gu�����Eh��D��H7v-�lY ��XX��[�y�[�x�Hة�bV�{� iŨ�u#�=�W��OdQ�H�W��tHO?� �E�Mt�� s.�ZZp�s��<�O��e�Dن5�����I�5��(3�x[�-ؓol���� �`y��L��W�I*���!�ةCz�к�"D�e�D�����9�!��7�h̡���D��1��A�2}!�߂�|��c̟>Q6�������'4P�����S�N�(�$��m�ܨ�	�':RQ�f�6a&�z��7([�Q��'��� ��g\@-sV"Չ^e���
�'�� ��3BT�q�ȁ�}��@�
�'�����w�.pf@�%ftQR
�'O�9H��zD���M��� �
�']v@�������9���$�nT+	�'�X<HJR�=|(IsO\>a��P	ӓ��'�����C�/&u�BG�=}��dX�'T�xQ������h��D2,��'R��@����}Q�ٍH�<i��'��$���\��<*���>6ؘ��'U�� C�Q��8���P�0��k�'b�	��^N�H�Р�Xc����'U0Tj�m1��� ƃV� ]!�'��p�����':ف�c�@4��'�́'O�Nظ:dڋ�>�X�'F�ҥ�G /*y�/�$�R�'8�p�&C�n ��QF�1����'~쩋2 "3���F�2=�	�'� � 5拈E`Љ���1�����'E�0/�$d]Yz1#ؿ(P!H�'�V���!2�|Iǡ��&<z�'�H�"���jM&��掖<F,i �'�^���سN���y^Y>�H��!D�(��(X���[Fi
-!���YM0D�`��ΤS���Z!q`�qg..?!
�M��p���D	Y���	`�oa�)��qa�����R�D��[x9�C�)D��ri��¨IR�U�\c��g+D���D�ʕP4i�5i�}Ұ#�;D��Y�f�i���(v��+����*O\<���1X�lK�B�k�<�[�'-����P)���p�(I�HBґC�'���X��j-�M
!®D�I��'[N�P���_=�MZD힎� �h�'b �ϟ�� �����'*F���Q�n�� 0 յx���H�'�B��S*�PS�}�'OĪ�Y��':�����.%~*h�V&DTT�p��'[ Y�F]ipp!A6cH�V���X�'����5�_8:a�e�D,[��	k�<��"ž) ��k �>�8=c��\�<� Q*�۬y���F �><B�� �"O�i��̓!+\���M~�@<Z`"O$Ii�H��Z�c�fZ�|���b�"Ov����)V${��'2�2��"O��P�*��fl����T�޽�u"OH)0�&���b �Y>\h��"O�0ЕC%OZX)Z��̚J#*`�"O���ώD��,S�J� ��"O�t�T�OG�8;c.^v, �U"OZEH�!賒�Z]��h�"O0:@�SC
��f�=5�x��"OH����k���!\�,j�"ODM9�ğ|��e�O�9�~4[	�'�Ġ#��Qt@b���@`�'d���,	)(b^��c��/Gݒ�c�'���� �=��x�.0��m��'�� ���:7���qd�/�J��'�(��?�#6���#ѶQ�
�'�R� �.�B�0�@1��ny�)K�' ��jD�ԅ����0B��S]��'j�yx����2WPd J�'-2(��' |<�u#��.<���N?D�b��'�@	��K�_-����l��E!����'N,�
��j.�P��>3TJ�'DQz0��}40��S�x`���'�
��CC�(���b
3B�tq��'�n!� �/z1��a�\�>��T�
�'W����@V�[vz=�aF�-���8�'9<E�Y>yFqP$��H�.C
�'����'p9���R���G����	�'��m9�`ph��	¢��mQZ�X�'��(�'�i�`=1��W5q�R�Y�'�.4�/Ʋ9�����6h@�R�'��ػs�ӂe��]��I��e�����'�(0P� �_B�Œpȉ�^HT1�'m��
���
��@�ŉS�I��(�
�' h��<�B��d�*61��	�'��Y����72X���Hɦ!j"���'�0�c
ѯct@��pu��yb]�@<`1�ąJV&��#(�y�h���`\����һbL+�'p���L�/K|rԫTT=��Yz�'K�d�4�I,4m�cۗ,���
�'��m��ܿ.P��2C�/8����'�T���@�Q�Dt2�]&����'6��� �܁exZZ��9.(� �'��e"Q&K�
D�!n�J�P`�'��p�O�;��x!f�%:��=��'w�'�Ia���bC�%N?�"�'~��n*`!�����Ȫ]�
�'��@㦙,-�b�h�N�YN}
�'2��v���N��W回P�"u��'�R�q���w��VI�
0��c�'�ƌh��$1�=
��Ʉ0��)�
�'����&.U�Hx���ϱTE�
�'��YS�L!az���,ɤ`�	�'t�= �m"!P` ��%~T�	�'&�!W�	V��Y(�,�a�ʠ�	�'�N�;��-c6� i�Z����'lZPc��]}�P\E�ѷ ����'˪a���_$���+	�mX��'�ޅ��Q�D/~�37䕌$��\[�'"�,�U$�B���I�`#�Ry�'��������<+vm���[�/���� 
@�A��J�-I��US� ;a"Oj�#�K�j�e�J���"O���ˁ-N�Ճ �S!$���c"Oh�+4�)C fTZVe�< ]��c�"O�!r�QF~5����!V ��"Ox��b�I.X�2f�.0j�"Op�"�b>_j���Z�Y�"O<��$У Rf�QU���33�P3 "O�,��L؀yd�h�F� .��Hw"O��a�lK�k������y(�+�"O��AR�P�A��HGG��rJ�"Oj�g�T�nd�j6c»-"�h��"O��p` #~U��HT�i���	�"O�!"���*E��7f �c"OI��j�5��$�f% 'v����"O���%"�F��e�`$L�E��`@ "O.�R�+�F.R���A�I��M�d"O4��f�a�d�T ���vicP"Of9����cn�{��׵�9�"OB�T���T��a��P�5"OV� �.F�R/8�s�D�%��"O� h�lT�b�)�
�VI��+�"O�:b �UF���0D^�8yQ�"O�}�t+Y�b���BSCW<>(��q"O\h�۠E*vīV�9wB�
�"OBL� �Ğ8�Y#Q&�$o<!�"O��A���&�m�#DC�$��R�"O.ȒA#�Ă��2�Y���s"O�]Q2Ğ>&T�`A��3jW6�� "O��B#ؙaip� &��OZ(�I�"O�<r�i׳)�BѠ�&
w��C�"O����$y�,��Q�S�cVX�"O��
��	&L �ֆ����}@B"O�Ћ�)N�4��ED]�DɖT��"O�Uȗ.�"_������<���A�"Ov��3�U�4y5�n�,�)�"OR0�����Z���G	8qz�I1Q"O251�JA>krx�z�/j&d��"O�s� v�T�	��/5�"6"O�M���4��ag��T,B<�u"O�m�t�īEA<<2!�5t04i��"O���C��ބ #�V� �%kf"OZp�B�F`"\�P������C"OL���0�m��CHXh$"O��?�U�扽B[��"O�u�፞�u����F\�mN�ղ�"O��hqꞷ:�H]"�Ć3�{V"O.����ӟU*�|qV��!8��R%"O����}N���Wg�7<a��"O��@�	_{�����'ͳ6+T�"O̱��Z�B�T��	X�Xt�""O�q���<Zg��2PG�.e?���"O�����C/d�x*��2�N��2"Ov��*@�]kz��'A�9�)�"O
8�e�?
$��8"��i[V�[�"O^ĉ$f\*[��QC@�_L� ٰ"O�MGFE�0�����Jصl�m�g"O� q�'��%�$%��$��ex&\s�<���;VW�`x�
U �̙�@Ci�<1&JE\����E�99츴��`�<EG�hm�`�sn�-Z�Ќ���^b�<��U0d�� +)T�-{#'�_�<���w�0\ǈ��V�����Rp�<g�<Α�2��! �$n�<� qQ��,U��
#.�(*��ѐ"O��10�
�7Ў�x�,Ĵ���Jc"O u�����w�eaGʈ�'���"Of�Q EP$��A���m*Δh�"OY��N��1\���Q.��n|�ۖ"O��ӬW7���M/itY�1"O�!1��=)G�����^�$"OnՉ�BR�E�F����<K��T�0"O(�q��}V.�AÜ}�h��"O�� �α&ரiS�%��"O�i�+�U��Rf�̏z�d��"OP*��ÿl��\�w�ύl����'"O:!�d.� �xRAA0[�4p�"OL�AZ6�5�� P�f���"O�d�톥
hTP!N:[�B"O�9��D�� iem� \���"O|�3�,� ���P4�Ы1s:x��"O\Q@4F�M�:�ڐ�ƞUmG"O�l{��/]��4(�X�}�ʩ��"O�����?8К-S ό;'|���"OR��e��0Z�hs�M0I�$ s"O�b7K�?@)�
�m���Sq"O�lG�=��}���5�4у�"O*h�2n��#�|��
L�nۨ�1�"OT��'+	#"`
5i	6���W"O�l��΍��QqW�6XҘ���"O� 0`z�{�#Z_Ԗ���"OH)y!ކ�·����`��"O�{�"�a�*=���m���"O:�B�Q�&�d�bŅ�"`�:p��"O�m1��ѰS�����Y,h�Tx�3"O*�I&!��t�^B�ӥa���y�
�>�L�+����\��E�e��yb�58��q3��.x�L:f�Y�y�J�!���BĎخ�&�2U����y2b�6"�:	�5dЇ>n���,�y��W�f��I�!��,`4`���y�l�4�%�#Y�LԐ�`Ɉ�y�	,\�^IA��W� �h�Q%�yB�/vH�P�F��<�0��K��y���mN�q�.[�/[L0���ۡ�yR�\dRE	���.}̐y�*���y���R���G�ӈ:>���y/HfO�arC��=H
=�Bd�3�y��ӵ���y�I�GQ�-���I/�yS�d�|�S�@�nI�%HJ��yR#��l*F&�,���"��A9�yR�A�T~( a+L�!@ A
5N-�y,&H�eI�ɐ<W�!�WG ��y�֫u8P!����T��)�[��yb�W/ea����۴6	~��c���y��h�!X�{�����+Ӂ7�j�(�'����%��emԉ�BKԵ(�f9�
�'L�tc�bL���I�Qʓ�#���	�'������`����a�8	v��'ѱR#A u4�0d���e�0��'RvE!�
4|Q�l)�%�Y��'�hR���3�h�2� ]sflz�'�Z���U(#@��2C��-b�����'���0B��Gll}ȁ��-'�l��'���5D�� 9�,#!)/��Z�'��@K���
$��l; �R"k$��'ɖua���)G4����ı
�'<�$���bR08r��91��y
��� r�yU$O���ے�r�Y�"Of��Q�G8�̨T�C�L�hȷ"O��+��1	曁��:g"�@�U�4D�h၄!q�@����
�	�p�9D1D�������ʬ����R@�1F#/D��jp,V�O(Qar�̽\�"�R .D�$Zq���jZ�����K�8*:D��h+D�x`[7!:]9u&�DJ�ՠF�+D��PbH�P�!���G�+�r��2&;D��[pϙT��4A��D>��o6D��pլ�,y��Ã$=���P D��z�"ѸP�آ��ߢ2PHq >D��Ο�−�O�5&�L3�j>D�q��5R�*���H�Sr̀�6D�P�A�K�o�,�ۇ�8{�ް��j4D�d���?o��yӥ)A��k�n0D�\����,8�.� ��ӊ,�x�ca�*D����':�u����9-��]���(D�a��C�|AN�IC�OaGڠ��:D�p�n��W�zefҢ����<D��a'dH�Z���� �FM�T�;D���h��`
~����S<�F�`��7D��0�"J*-��ti��D�@�6��2D�$2rK�(��4��^�u�C�0D�,���3r�@�p"C�&����.D�T�'̴d���:C����2qڳ�7LOb�)�@�{�:���'<`Ҝ҇��*W(�P#���'��zQ��}��F�J�k�Q����R.�"}�'����g̚�T�԰�g��.�`d �O �q�l�S�O��P�MC��薜!�����'n@����L���؀��Y�lH%oB�<l�y�4+����v�Q�K�4r��S���e��d�N�^����)6BN��q&�&<��Y)P�qO�(�*�)��O��� �B�Z�K4�Ԗe��;��1!���.�Zw`�J�'m�d�*�B+�~�`@U��O�>Ƀ���B�ƅ8#X�J��Dzc���Xa8}!���	�1�fY:2j�K��Pa��Q�/�5�?��Ez݉�O,��|��P	���: R�:�H�H`O����i�����T%d ��l4�g}2"��"�����7�
d���-��Isn��?�J�-~1��c4*U�.(�˒i?�a^#���h��$;@�H�q8�r�G2H|�e{��
2��0�?E����.o��{ģ��4\f�Y�m��:�yr=O�a�.��`�Od�Y����LQTذ�B�	]��pС�Tu?�ҦM�<15�Î�~��SL$1q�̚��"��eB<@dd���dR�<aA���~2�SYy�d׃sd��� A�6��x�l\]�r9lZ�^B$�'��7��?=Yu�W�G�t�V�Jw^�� ��U�zQp�O��	�A�a���3��<P�.������/�)~ɼb����ɩ����'7�@ڷ$�))�����4��O��+&�ivn���e�O���>^r̤���B�a�v	)H�G���.�G�*��5�,�>�G,�tC�����(������\P�<���H�F�J-S��#{'��s�
L�<��)ۇ-�t�x���p�eKSJ�<)C�E)o�(W��1G�%�d��I�<���ΌK^^��+���hI�<Q2응#��P�f��Q�2)��Lz�<A�b��$��Cw��vZ\�
T"�A�<���'���1�#�;��2��}�<��a�3w/n����G�:�Bm
2"|�<!a V�	�,����I�F@f�-�y�<q�A#n_�鑥�C�.�YKs��t�<���:�Fd��`ٴ
4��E%p�<)�� fߖ����	�*5)�E�<i%�~LIW��(2�rF^\�<�#�]�8!�ُ%�"�'"�W�<9�2}�Ȱc��K��|��k
P�<� �L�wƒ;G���Ѣ��6�J��f"O���� ;���Y�≁;g.��u"O�E�Z	��y���/�ZMq��]D�<)�j��5.�	�5��)��%9F�@�<9�H�^M���͊�Ke̘�3n�|�<Ys�?����䍏�*�V��*\A�<�'&�ⱊ�;_�䙘���}�<i'G�Rqn�äG��e� ���R�<��hT�6��y!Z�EO�����i�<����햌Q���}�V,���~�<9�'^/JIF �CD��"��Q�O_�<�tɗ�K��i
$O�M]��� b�U�<aC�-C�\в1/��,��g��G�<�ҤҪm����Q�܄��@�+�B�<Ʉ��6�p�i���(oŖP�R���<�.�9�>�Մ^�~�6�QS
G�<	#kX�}	�E��k�Dd��C�<iD��T�2ԁ��Xݠԋ�kLJ�< .H0�>Q%-��y+j��W�QC�<AE�̕5�����!����{%!Df�<�f�NI��U!�:��%�f��b�<12�&T�6)��ჹB(�3��EF�<�s'A�y�ЫT��8I��U��C�<Y��A�U0��K	,<�lăr��@�<a�%2��+bh';��$a �s�<�3Y�c!x�sN�&Y��y��Ps�<���
��%lU;��5)F�r�<a�ĝ*Ō�$+E��@X:WA�D�<�֡X�F�TP$Kv4X� D������*ո0i��g� %2�`9D��@�K>�b�zƇ�F�Ĭ���8D�H�SlF���ljƈDϬܩ�E$D�����ȃd�Xi���´/c��pui!D��ې.��I�̙��B���-� �#D�P*�j:^q`��7LƫKWNiid�"D����jŖ9'��`��=?���@ j D�<���Vkx0{2F\�u�8)�g D����I(٢��NW	��Ts��?D�DA�M=���ĭ��U[��(6�<D����bhS\98�`ӱ*�j�y�(D���Q���f�t��LҜ
���0�E4D��c3�Hz���Q��_�6|�T=D� �&BW���)2��p"4�à=D���F�Ը8����3!�$}&��G�(D�l	��UQ�6�p`œk��9"@(D���g(��i�����&����%D��C�*J	Eq���P'ѨČ��(D���v$P9�`A�O�I�"��j<D�|S���Zǩ�{"�գç9D�L�v��lg���m�7��9�a6D���V���h������HR�t��e6T��j��	� F�'��X9t{�"O  ���t�8���mV�i.2�RQ"O�a�S.�S��\����!�|`�"Oz�d$Sh�ԠE�&��h�6"O���$�r��6#ޗ}�\S�=D�"�ElJ��\�݌�Cv":D���e�D�H9��p2�KR�ܑE�9D��� � ���pi�;���P��%D���k�6�
}� ���@1�D"D��s���:*\�� (��U�т?D����X?`w\�j���7K�`!�`� D���������=14�S�#�>Ţuk>D�\���,C�8�C�O�J�{4F:D�� nѹ%	5^�Y+��G,1�⁂�"O>葰B(m�PH�Pgl��ؑ"Or[�呒$Ez��֏sH�1�"O�i�ɄM�!@�mF�W��`�"O�� �'�j&�CmJخ��P"O\h��'ʱ'�jel{�� K"O,LA��ۡ6���"cȚN��� �jd�J�(q�i�%蟙,)4m����=�4h@m�1B�OK���@���,�����Y�L��B�jV��ȓ\�*�AϞ�J�"�ȓ�'����A'*���g�	$�"R2(	lÞ�ȓ%f�#�f�C��p �"�+
���ȓ2Zi	��]�n�d�� &1|�P�ȓr�T�A��=/x�S�m��Z�ȓh=�-���:&���������e�ȓz�����C8.O(p+WgHP�fԄȓO�ȑ�ӎؠl��jQ+�Toޑ�ȓe� )"��I{��R%�4�tT�ȓ{���FC�������s>����]���
��1�ǒ{P��8:س�ٻPyf�Y!��}0̄ȓa�|�� ��`��'L��$|�ȓg��5XՃP�V����3(�@|���Iʠ����$V��@�dD�v�M�=y�������z�&d墒� شTS��Ρ�y�(M�?���Ñ��b�~�Ç����y�� k�<-���V ��c�H��yܖar� ��Q�HȀkvɄ��y����0]� ��9�`<����y��̻L����9�1�p��~�<��B
z���A�@�<rd9�`&AW�<ɷ�R-3�B,��ȑ�LyB�cB�Q�<ip�έZ|bd� 1�,0#(�Y�<ϓ�:�XÅF�c2_�<)[�w��u�r�ј*�Qct�@�<iQ���l��
��܌�U��W�<� �ߺv�X[�CJ	 zZ���n�<���8W������_F�#g)5D���h�0l��c�����p�1D���ƈ��U��z/R�rAL�Ь0D�<���8s\�z2�;-�$�*OD`�&��e�>q��I��A�����"O�}@�׶�F�ĭ�)e�Qk$"O�T;w�S�>����Ԅq\(js"O�P;�Vi�JDɠl�&d lD06"O`5��J2���+�
-�1�5"O���s*�"M�F�D�)[�zL�b"O�)�pj�pؐ��&._&+� ���"On�Z!������4�Ww�:=#�"O�H@�Ȇ�3)H�DӰ~�~\�6"O�=
&I��?k6� ���"Fn6u��"OR8��BW�}�z��@mٹk��y�"O�m�C݅'�pi���K,IaJ��G"O���BĮu�@�A�P�f�]�3"Ob2�S7,@��Y��� ��a��"O ��!��"�FeQ	�<O�T�f"O�ig��]@4�y�Hǟ`���&"Oj���N]n��j�h�� ��Q"O�iT���(��!A8��*�"O���囐7�z@�a~����b"O Q����^٩��5�8�	�"Or:@Eb��$��C¶[x�$�G"O�˅��	���3� � pRЂr"O� >My2E]d"L�����C���"O�̛�F8_��ia�%a%��"O~I�5/E�z���OU�wp���"O��l�!>�App�H�va��/"D�tcF�֞(�M!�a�D0ir�
?D��)&� ^КL�m�����3a<D�H�$iB� ��8`F��J���2��=D�|:�d�Z0�с�B�0C�X!$�<D�`	�c�?����򄋖_�h�%`<D��B���+�f�J�J�0ɤȊ��:D�����}ք��kH�e��=Yq)%D�T�+'B��p"�@�+h� �h�!/D��AՋ%i�Ԅr�T�V�<etI+D�����\p�fh��HE[ת*D�<���Q:�d�Q�	�����)D�\��J=p���%'�e��#D������U�*�i �%~�0����>D�L�u�ŊT���!c��
pa>D�x9VDF�j}I�!�A�O��U9�l/D�h��&G�d��%a��E,D�D�mއ{�X�cfk�y��!�)D���r����ҔK��v��.1F!���g��mk���� �\����G�o!�]=�T �bLQ���R�ՑL!� ��1��	-~��u4G� h!�D�*�iJ�l4x�hH��EԪ!��cҼ�2%�
v�����2�!�䒬d��a���xlj�Rb*Za�!�$�	h�}���X�8}���q�!���sz�����e���W/ 5�!�Ec��=��:h��m�*�!���V�Y"�&ݽD$���2�!򤅭)��HZJ���N&P��hc�'"� E,@y0`��4�̞^��'��X(�
�VQ[��L`���2�'�܁��� aԒuZT�DX5X���'0�˂�Q4���to�x#`%h�'�B�3j�.^�v)B�
�i��%R�'�x	U݊���1�62�@�'�`D��M�%�a�������'�
���L�\)��"UAR
Tp�'�n�Х+@���垺@ɰ�h�'-P��c�����7�X���' �����3:@�s��n#�'�.�y���2�\5�Q�F��h�'Y�d+��FvD0aI^�p�l$��'�8=(�.��q�2���ES���'i��xT'�'S,�;���F88a��'jRy�r#���v�0��q�5I�'�h�`���8=>�g�H��
�'?����!�>8p��`��rH	�'��!+����z]��xd��#l�|I�'�Ha��I�1�t����ee�8��'��a� 
�.��)d;^��'�,8@  ���     �  _  �  6+  �6  CB  K  6V  �b  �h  *o  �u  �{  �  H�  ��  ϔ  �  O�  ��  ֭  �  [�  ��  ��  g�  :�  ��  {�  W�  {  �
 Q & �- 4 H: �=  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p �j�������-T�p �(VF�e�1`$D����@>8p(I��_�:��*��"LO�⟨�v$ˣT�9�����Q:�j D�<KU��&Y��zU�͕T� �a¥>}��iS��?�����+G�>L��]?�	4!=D�`�(��N�A '�SEp8��=���<aGe��W�� ��!�,U�^T���A�<Y�)�'e"b=�f�]��4��������Cj�Ff��8����T�Mc���'jf"<��  �``��햴@|��T+�"Ga~�U�<�� �%#N�k��E�N� �Fa'D���í��^���%�9T�*�%&D��h��4(=� ��)Wn�`2 &D���Wj�,:��C��-��LI��%D��mڧ=�x@�i�f���6D����!OJ����,loܰ���9D�$�v��4g��)q�ϒn����6D�������sv}:,����yT(�#p#Ҷ!�,0'$ݠ �P�V)Ԑr�-v����{
� �@PB��iP�J$�ćv���Y�OL�=E�d��-A�r��7�ügr�����y�ӽ,"�QP*�'lo8TJ��y���%�HPW�[�Z��@-�ȸ'�	)-)Q���E"c!:\k�(׼j@l��N���Hx��͓�A��%�bP�ǃ�0�B��? �����/���	������}�g!�Sⓞ��h��M�$�]ZCE�%�OL����[`��^1X����s̑-M��O�=���!�"�Mrp�o��W���Z "O���fcǊrz*#�8$�ڈc��IN��&��@���1o�R=H�0-7D��p�8H�������:7�N��3$�O�⟜��>��a�3��%�4A7MS�0�>�d�"�,���,I9���#X�s]&�P�u��LX�Ց}���O�w����'�ў�>=��1��(`��¬P��0�gD M��B�	�;�N����Y�W�
;g�.3��B䉼(��(2�EQ0W�Г4JՈEcV���A�DK�z8�`�.Br�pg��i�!�@�{2�Y3�f V2&��u�!򤆇`�"5��k� �j'қH�1OZ����kY��pI5�tEa7��)�џ�G���602ȨbtDL4G�&}���y���02�����͒EG��L܇ȓ*B�#�3z��t!�&j�a��*�(ɲ%M�RF�	��F3~|$<�'eў�|�g��+�Ikál:�c�3XnC�e>Q#R�@5̰z��:�'d���DQ��8���#əb�!b�ɿ�!��y(L���N�%3��x�EJ? �!��9.�āEc�2BB��5fµp\Q���'W�~�Y4n�=3*��#ǩH�Xb�Xɡ"O�Hz1➿=Vx�����L<�>���9�S�'�p������	,j�Z#&�,�
��ȓT�0 ×A�LH�C��9�n4�>�
ד�F��4-�9;��-���ً$*4�ē��u�&�αi��R�gA��<��^~H<Y��x@�0@n�$&}>09�F��<I�n�T���gI��"pzR��~�<	gG�1F��2�@�� � �`��<��.Q+A�Z|�����B��?�$H���j�4O�d�N������ZE�ȓ%��mٷ�Z#�x��0�T$���3`�����)�z�Jd+N�YH�ȓgr��!��=S�"N�w����e&���.�3I�lՓ�.��G4�=��\ʥ���(/��M) ��#�����n�T5U��^T*�%�u3`���	F�I�xp*e��G�����i���vC䉵�x谩A�S�h	p���|���	��h��+�%��]j@�Ժkf�W	*D�0�A�
�[8���f�_�\H(�i��(O��l%>��6�Y\](�q��J1r.����1lOV�4x�	/��(��J	 G>�xa���<����+��e�W���zl�T[�k˲+ІB䉴jXi[��-;�r(	$�&9I�C�	.1����J{�N�1��R�{�d���ϓk^�):�MH-[��Q�m� {9�D��VKD�e�Zܼe�q��3_XȘ�ȓFj�����<n!�Ui�/ݲv �Ȅ�%�yzE. %����Z�f%���,���OH����7O���B�L����E���'W���?Ad���\����G#S/Kp���-�f�<� (Ѡ� F�.I�p��/Qmp�x��d(�Ş;�ҍ���� .ʦTtK��V;z��ȓ0pt���@�j����/�(5�$%Dy��'*�|�A����i$ �UT���'�"��ħ��
~,%���^�T�=��4�Pxr�6K,,�&*G�9���kSP��y2�2�.4�`��B.��s��"�y"�ͳ��E'9�L��O�7�'����A-?��kW�Y2`�*� "O�8 %�X���h�/�,I��`*�Ӻ#����^�h`�A=I�h��)����p"O�7�:�x�e
?{��27dӪ������?U�g��Y�91�39D�y)�$J�qH.e���hO1�Z����)
��S.���9�$���3lOj0�g)_;�@-�6�E��6=�"�'?�承0��Q�U5F ���fD��fB��Z��y'�ػG�}�d�@z`B�ɤ/f��:AH(m+�H�3�H*:@HB�ɖ~�~A�څh��;�F��$b�PD{J|��I�6�tbc�6U~`8����E{��ID1X�
I �=c��yo�Fy���y�|�4�)�x���('x9C$;D��X�a�8!�H �2l�GHmB�{��B�I�Zv�c�Q�0(NXB��r����	�'��)Z���4	�m�c�LCm0˓H��$:�@	p�4ez�IU�~bu:�`2D���2n����3J��I�h�Ñg;T�8�a��j^�U3���>K@p��"O����I�z%�F^�GOs%"O��p��/q���6��x/R���"O�� �DP7�����j��+B�\Y�"Or����^/�l��Ʋ���"O<�R5�X�>�N�#$@ǅn8��Q"OBX0Q�֩P�
�P��
9a�(x�"O��G3=�J%��4/+� �"Oj�� �-C"tt�\� �b�"O��b�F_�>� �*�<e(���"O��X�d��P�p�i�*�5�6X��"OL0������A�G�x��L8u"O�$�_X��#�i@�(�DE;D"O\I�pkԟ79f�ʜ�h� HA"O
bg�	Y�
�f�A2e�Upq"OZ��$��W<a�7I�&s^bm�`"Op9��	K8�F��X�{P����"O|X��&�sG0�+�� )9 6"O6����/��a���5?��X�"O���.�6L�<��d��p�F ��"Oܸ�F�J2�&qG�Թ.��`5"O�M�F�	{
j��`%�2=��d�"O����=�&���#�Aٲe�"O��h&������M�.$�u�"O�8h��I-y@l53�
�}~�d�1"OJ���m�T ��	mg����"O�X�Pca3<D�d���J�!�̶q{���%"��I��Y��J�!�d�uw�̣�C�$��#��!�\/k��,P��˘.=���`ʵI�!�DZ�vB"�c�B3�<#��[�r�!�D��#.������
ɒ��2��|�!���0�ā��b�D��5�5�L24i!�RU:(����ܥT�0��3.�6�!���7r3?4Љ�j�S�^�	�"O4:�K�mʠ񘃫ؠ��Hȳ"Oȵ��O�-W^݁�I]�
� �AF"O� �3�5bR�T�&#�s��Yb�"O��;tȖ�%��4"AA�ht�1�"O�9�SH��5��0��W�	g��y"O��QU�!L��a.�>zRP�; "O� ͨ32f�
E�sP�(�"�'
�'�"�'���'b�'b�'^2P���A,a���L0-;
 ��'�'���'���'��'k2�'4P����D! ��C#iC�'m
=�T�'�b�'�"�'���'���'R��'�2�[�n��<p�@'dU�Iv����'�B�'eR�'%2�'y�'��'lؔ�mn���%֤pX�� �'���'J2�'*��'��'��'��U�e� riZ�TF  8���'���' ��'�b�'B�'y2�'�fU��!�� �%��	�g��%�u�'/B�',��'���'���'���'v��Q,��.�
9��PyS���'�2�'���'���'��'j��'��������|�%��Q�t�[�' 2�'	��'�R�'(B�'���'.�TH���@��tbS "/�}�G�'0"�'��'cR�'�2�'%��'>��!��T����6&t�v�'/��'��'���'���'��'!�@It%	W�f)
�m�4$t`��'H�'�2�'���'���'b�'F.I ��B"B`���c��$Rd�}�7�'���'��'�2�'���l�H�D�O�@0�J=O�����bF[���p7�@Dy��'0�)�3?Q �iM�<�g� %Q����%O3&X��p�G����Φe�?��<鵵iJ�-��j��>�P�o�(s�DtA��y�r��L"8�hhՕ�L�!��)^\��&�~�g�lg&eA� �~��%[�n�P��?Q-O��}��@��H^��r�K(f�Nۄ� L�����'[�n!nz�=I���u+��!�Q<f\�0	�#�Mӡ�iR�>�|�A Ÿ &-����xk	�]M�Q�`ǜT�ʽ̓2��Mv�	P��A��4��$K�^���(F�~�0�l���ĵ<�M>��ipF���ybV�&�5��;�jix�)���Ob%�'e$7mT��ϓ��DF�,�B��"Nӳ#\J������4U�	�g�8�u�	�8�c>ٱլ��i���I�w ����`�;P��)&!�T�p0�'���̟"~Γ'�vr�T-
�$P*��3L����,ěF����d��e�?�'[������E�K��i��"B0j�
��i+�vq�V�ĉ6Fr������j��U�.���D�Z{�䈧�B'C�嚝�x�����A{�Ha'+J��I���kv�yuE�
B�@n�?/�Q����@ [��Ò�@��r�Ũ�Kk\h��4?�dbVdH:� �����4�ص��̭piВOj� ��*;-fp���-3s<����׉�����C��uB���F@�P����*	,r~`}r��F�}�X�V!�4t�zJ#X��H�l¿Paz)��AS�a�|a"E��3����$�	,\e��H)L��蓀oűLYJ�3#�ҙSxn����[�Ɛa�"��u�F@	�
�0`��i	�'��O���$̴��"��tg��b���+��|l�֟ ����#<�~RR�P�����.��9�N���!CqN�M+��?I�����x�O�ZAh�IԡFC�,��X%o��(j��a�I�<���?��g̓�?q%�^�<�怢F�C�}"�y�7ڥ[����'���'�����3�4� ���O���ǖ\?`XZo ��0TҦUX}�'n؈��'(�'�rK��]yA��:BC��sC��1K�6M�O��9 jUy�i>��I�T�'�9�-�U�-��h�q@�d���zӴ���"~�1O����OD�$�<���p���(X-��A	<��&C����?9���?)*ON���O*�k �E(м�*%B�$a#p!C(گ~1OH�d�O��<Q�����iFtFԽ�F��O��@yu��u	�	��|�I럨�'���'C�E	���*�K��[Ʀ��SʀJe��5Y�t��ԟ��	oy"m�$�L�����@)7&Ή��#٨L�8���d����I�� �'���'�:t2��PC���\)�*�ءiP�^�7m�O�D�<I���^��O����5�lKg^�-���ŋADΩ�3�D;�M�*O\�d�O��b���?7m�. �Z���߲wn�IXf%֐o��T��Z�ƛ�M{Y?�	�?��O��lLK^��uf׆)=\�ك�i�r�'���3!U��S���3񤓾cDqP�&�*xE$����*v�fŜ(�6M�O���O��	[�i>�ciJ�4��1�6��CT41ulæ�Mc�F٫���O4�d�1O`�dC�=��ȓ$C�{���Y�OP7��n�`�	ҟ�"',B����|:���?)E �V�$�Đ0d� c�X�A�I����	�bV�c�|��ȟ��I+~SxH���L��|���S4R�옳�4�?)�i^�{r���D�'�]�L��N�F-2��� "`�pI4̑��M��#p���<���?�����$�t����§��v+��HRJ�p&��+�Y�I��X����'�r�'���c$���5
)r��-p<Ȁ��I���'b�'�W�d	�L���DNh�pAA�:j��8�+�k�R��'92�'��R����̟(�%��~�E �$-��y$�F�^�Q��!Nd}��'"]�`���8^(ؔOx���<�b=S��X�}�"u;6��I�7M�O㟌�I3r0�]p#'񄌌
��\K4Eߺo��!��<����'��Iɟ�CC�E�d�'#��O��D�Y�#�0d�������(�I�h��`Ԋ6pc��g�? ���/P	\Ш��p�C*ar@bS����2v����͟����|��iyZwa�@:�&O
O�k�΄*rr�a�OP��@�ةjd��	�isd�;�$�<n�9p��ϣE�-�b�b�'���'��DY�����3��g
l��C��.��	` r�m���!�F,�)§�?��,�19dDh�kɧ{�ԑUm���'�"�'&`P�P������G?��<bS,ea�ȅ6H�U��_#.�1O�\q�L�\������I?y�V�9��Z �E�$��0FB٦���)ۨ��'kR�'v��Ĉ9h<`�`V�M����F�2��I(t츔a��+?����?*O����5A��	e�ǫ,��``w+��蜓bκ<����?����'OZdr -�g��:yۗ�ږ'����������Of���<1��B��q�O/e����sO�tX�FQ)o��t��4�?��?����'�ȵ� .��MkA�v�(��#� y��A��GFY}��'�]���	
T�>��O;2�L!O�lhT@
/Qo�����YP�6��O*⟼�'��@J<�t�B�n�K���+(.�"��ئA��Syb�'���	PQ>e��矄��<�<Y��J�%��m�O	�PM�p��}RV���se5�Ӻ�V!Si���3���U(02��v}��'v��qp�':�'���O6�iݹ�5jՃ0��})@HJ9�4P��>/O�1�W�)�)��{�X��I;B\�b�` x���/�/XKb�'���'���U��S��h[PǊ�g�*��#h���)9 �߁����>�b>��	�g2�"� �C��d(E	ڟj�����4�?	,OF,c�<�'�?��~r�]���Eh��x�%�D�J*X�#<����D�'�Od����60v����0K�Tj��i�Bo���	џ �I���=���B+	�1+2�t�p � �	r�ɻJ�?�����O�Qfb̘W�~z�+����1%�R ���?����?�b�O�8 A���hI�.�d%p'�i�V�C�O����O�˓�?���ˋ��TE�7��<��鏈;���R�M���?���'B�	9�
7m%aq�������)�$�����ퟔ�Iiy2�'lt��R>�ɲ8˄}sv��������c`�5+�4�?a���'~L��ɛ�ē{Qp$� �*u�K�9�V5K��t� ���<����L��)�����O��	E�K�.`�� 6_(P���ע{A2�>��}w�iBw�A|�S��M� 0�,�I�rݐ��������D�Or=h���O��d�O�����Ӻ+�f*�J�p�����Þs ��'$�lޱ�Ic�y��D��@^��ǉO�L�`���M���Q��?���?����*O��O��F�(19�/P�0F�"����2�N?^�b�"|��?�$�bW�"��$.�@��i���'�b����i>�����n<��T�T��~h�F���ta�DɔI�f�&>M��ğ��/�f��j�k�<%�(l���n�Ο����cy��'2b�'�qOv���mv
����6~��ᨂY�P$�N#�J�?������O�Pq� C�0��C�A�t��J4�^�?,ʓ�?����?ɈB�'�Z�)uc_$D��q�f�-*D!�F�j����O���O��?Ip��(���"@2D�:�T*O��ɒS?�M��?I���'��a�*�X�ߴJ�&����r\��:~���'R��' �ğ �7��K���'�`: h�Dr���.ۯHR2���}���D,����pqN@�O�	Wl�)rN��"�ꍼ@�`�Ʒi��Z� �	�Kج��O���'���X�6�5ڧa =�H�)7���o�c����32��$� � �~"����hHhx5|��j}R�'�6��P�'^��'6R�O�i�ᳪ�2i�����L�u�v�1b��>i�-�͋B�Qn�S�o�j��I�>t&|Y��&ZRdnZ�#�p��IП$�'y�V��ʟ`(B���1�����ƕ�y[�LJ�L��MC¨Z� E�<E���'T�(A#_:f�0�[�kY�K��W�x���D�<!��6��4�~���Oh�	����)$�҆y��@Z7�C�f�~l �yP/��r�d�O���c4�<�YȰvH̃Y���Ct�b�$��bdY���I͟`��a�9��ԡ���3j����v�T��'���i�����O����<Y��S���$H��0�19u�V���&3��D�O����O����ɏ�`2C��.�X3kV�y�����*��?������OL�0��?Mm���P(Ru֑�̤��,i�����O,�D1���k�ٰ�
l�pE���f��4c�Ɏ�4NL��!T����ğ��'"��ɡu�S͟�PP�ωZ��h�L�w^~}P7�ϋ�M3���'G�(�
S�"�J<�ѪڞET���$�D�>d��]Ǧ��	�����ǟ�I[�oӞ�d�O*�D����/�(*�|����	>�
���ʦ��IPyB�'�j��OGRW��s�4šĉW�9�vdۆ̃qP����i�"�'FX�J�NnӖ���O��D�"�I�O�pR0`T�zΔ�	sc˒v����U}��'��5�Z�M�����4���O��I�!H�&c��zvF�/��A�4R���KR�i��'��O��D�'��'ij �Є[�1�4s�j�qZ9+�C~�h�{V��OP�O��/���O�p� ���!�5 D!�Rfb�ҧ�i�2�'tF�Mr6��O*���O�D�O�[1N�>�2�g�+l;�["+uR���'��1}Ab�)
���?���N㶘+�dP�:�D!���ƣ���[7�iM�\6�O:���O����K�$�Oh��b�<`rt�#��_��b5S� c��o������������ny�΃S�̥�r�M=M��\3�d��DD��>Q/O��d�<Y��?Y��W��<��Q8k^�ŉ�dD�H4�����<���?A���?y�����
"�.��'
� �k]^��E�o
�nBy��'u�I���ӟа��m�0(��¤L�&6�0}3�x�@������O����O6˓B$C�_?A���L���AĔ�N�8��WIú(��HY�4�?�)O��d�O��DS(�~�^>7�5B�� �U;0[�c������'E�Z�$8�� 9��)�O����8Ԁ����֘���p^�$[�N\}��'�"�'ߖ��Ο�I]�҄n&��ש��PGT0���ϦU�'���	��aӜ��O^�Oq��T�A�X�o�d���58�8l���ɪN-"<�~���D�^FA����>������妱�#Ɵ�M3��?���:�xb�'!
�!�-��a�I�v`��C�o�*��7OΓO>E�ɎW3����a�J}:�,��ȉ�M3���?��v������x��'���OdA�q��:���%A'iܩ��i<�'t�	3T�+�I�O����Op\1Ǆ���Q�P��t��E#�Ѧ��	��&xK<����?�H>��4P�4eѪ1H0�q��'��X�'�xu(�'��I˟p��S��mNH	R��R�D���1�&�oFI�����?	����?�^ڼ�	��Yt�Ĥ[%��;�,���?�-O&���O8���<�Ў��'��6QT�)"+H=]=�l���G7f"��ȟl��C�ȟh�	�!s5��)*�v�a��1�NTy!�m�V!��O��$�O"�$�<90�E�^,�OhXȀ$�֨'�HQ�\y����z�&��-���O$���%U�/}�.	�h%��א��PB6����MS���?*O���7(��$�����Ek�/�D� Ay�"Q2�=�dp�	��x���HՒ��e�~�UNET.�}qD*á�qZ�$Ӧ��'����d�s�0�O���O�8�[e:�##'�X��a��}}<�l���ɷ1����F�)���$�\!�V�"S��<I��\6��1J��1oZ��4��������ē�?������W�ⅲ�K*i���jw�id��A�����������練PCܻH躨�S��c.�6��Oh���O"8��R�I�����q?)��>N6��D_;	�����F㦥$��+��r���?	��?y�/�Ok.�:U&L(	�n=�A�,Km���'c�):��:���O�D?��ƒđU�T8��}���}8���P�x�S������'���'��_�8�����k�p@ H�
�>��#LS�rFB|BI<)��hO��$�G����-��X�}���0 %Ka��Oʓ�?y����O�0��C�O�q/YBeQe�.v��m���	���(��j���,��2J�b�aӂ���L٫%���1���-h����Z��	ҟ0�I~yr�ϧ ���:8c7�ԅJ�*����Bn�	J7�R��Ia�����"�c���D��e�<�[Gň9-$"�;��c�����O�ʓT66��֐�$�'U�D� 3p��/D'NzV�)Vf^5z�hO����O:���~"D&��ZA�%Ε2b�A��Ħ�'`��`)o�4H�O�2�On��O=�H ��Rw�y��]���o�p��NQ�#<�~��\<8b�U=\�$����2�$E͟<�	ß��I�?���� �O���C2��[�heY�+���h6�n��K�M�St1O>��I`��iq�/�N��ff�q=�Q۴�?9��?9�K؋^i�I\�t�'���œu�R�(t�|�!�#,�=k^�b� �%VT�I����	ܟ�K��Y$�ٗ��i���ꑞ�M��!=0�#���?��]?��	M�I)�}
�ܣv�h��k�
E�1q�O��cY/#��	�|�	by��'+�pY`�C�M\�ir,�3�
��Ư����'���'�B�|��'��A�9E�E����"4�JS�¨l"�	�k�+����O���O|�^�� $1�!���҇W�t�BD�� =�̨BU���I���%���	��0��ü>���{���.(#kb��@Q}��'	"�'s剢5��M|:�ȕ�?t=sr"ـ��uAͅ�7���'^�'n�'}�C�}��]&o-���jS<k���_��M����?A(O����,Nw���H�S"o���P�EI?#��9�%
f���M<y���?q�hO[���)�?�<�K���	�X)s��ʓF� �c��i�2맧?��'
��	�2�Tb�I�2o�0��W'�~4$7-�O0��	o��b?����R:��l�$$�%6��A��q������NҦ��͟����?5RJ<���3��`�s�Z�k�� ٖ�
�U���0�i�x�ˊ��Ɵ�9���M ^챳'�,,�i��)].�M��?1�S|�<[���?�+���d���2w '�T剤�y/ؽX�L���'��#��d�'�B�'�H�)��]1BI���9=0��(b�u�8���Td�'�X맒?�����l���7_,|t��@�HW i��U�6�bK>���?9��?y��fG� �L�ˑ7W�ĸ�� 3|���1�oS�?y������O��O����OŪQ�K�.���H�FM����sK��@�E���X���-O�i��΢/=(D0���Gɱ"��)2�j\�J��Aa�$I5�yRA[�>�j9+N�.�x/����'�N4����;	����k_ah��1nF�s�s`�͘9
4 ����s�f,�n�rP����r���g�ć
��pID�P�b䠐b��G����i�N80��a��P��c�P� �Ā�O��P��7�0�7S�<+���!�~z0x�"KܐPoʭI��M��������bԺ �<�8p�i%��ʟ,�ɗ�&I�䮚>i��!a�0*A�p`ٟ6�'[-��z�n���t�E埓+{�M�O�I[aķ6���MK�N�ɐC�\��qi����Zw	��ct�וE�$Q1vbЭ�O�h��O|�oZ��M����O�RTلm�&!oV�� �ÿwL^P	�y��'{�y"g��a�*<�U͌<i���$��tў��HOhMq��O�<I�r�$ �� )N�4$�����O|��A2N��ͻ@��O��Λ��'���ݽ|��%q!�P�bLpo0�e�dI�'~��2��H��<ta��}�'/���J�&~�hU��b�p�"d�3�R�t�Y�e��!�.ʲqF�隠�W-C	�$	����n���a�wH��h�9��0��#�8h�n<��'���p�2�4��=�V�S,3M
��ȭ0�~}b�O�<i�N�l�X�"r�-a�Pp�(�<���]H�����h�'�j��늠�������p6T��!ְ:��t�P�'P��'2��zݑ�	П��'p�@jp���M�#A�r��AI��d%�Ҧ@�"Xb�󭙗�M�'&w�'2��w���X��"ц5�)�Qh�qa2���,XN��) -��+�f	�=av6�<�'l�2�d�8Y=�=�Â�j~]��?���hO�q���!X�}�Tg	��x��$� D��J�F�tu��0�	�5�h1 �F4��-�Mk���ā0aV`U�'�"Kރ�\)�a煽H0nt1��UG���'�2l���'8�حPbO:|ȨHq&YW�.���oω�"�����1CU꡺!iF�R�* E~2�X��h��c�pWb�'D5�F���?)N�WCŊB:���� � ][���V�I����I�Mk��i��.��|��4*3�� �F�!T�	��<�?E���#l9$�⅕+�=���x�`v�F�I�בJ1�(
����H��G�O�˓%�0��2�����'�Y���	#
�$��@%$�eԽ53���Iʟ��c5m
 ej0�k��Y5L �u��[g��4;lRth�E��ؒJ�#���'V���恙pj̭���A'E�(	��mx���YD�;a�m�F�Sm�{vi�F��Q�O�0��'=\7M�a�O��D�JvN�� "�2�
���4�����l-Q����`.*P(C,"fN��=ͧ$�����G��d�(�EB��XRx�󅯗�MC��?��:�^�
�*��?Q���?)�Ӽ����B{B�y���g���q��̍K��Y�e�<;�i1��J�Rl���tLG.���͓L��J�A�(i� �E>
�$��gS4=p5+U�@�+\�q�@�L|��?�g�Ҽ�#��A��0�&�W�I[.�N ��FӦ��R�Z����Y�����1���3<�%b��~ڼ���8��s'H7c�k0�F3bqHt�'9�#=�� �;�?Q*O	2S!� (��ĩ��μ(n�pꜿk|.D����O����O��d����?�O�pM�B��
�%����08<�)BJ=f䩨�מ>h ����N��xUR�Q�'M��Ĕa~�� ��/���k�9_HNl��ʊA"Ms	C�z�RI�q8D()"�|bbI�o��� C�>ap���@�3��%C��t3�&cnӴ㟨������7G=������UcB��ռ�0>YK>�ChڡL���v��pK��*�k� �IFy"��Ij7M�O���ހZ(̊�Aɬ�z� A�ڴ����Ou1�-�O��D}>���G]3��Q�$[,4�<��B�2O:L�GF˫EA�4����E�F
Q�X#��Ʋ �b�G[�<dp���__�1��OE�i�8�U�	m!���R�o�TH:5�]q�n����h�@S����EƪN�F\p![�!��'�}��I��t�?E���� .`�eMN�.g����:�hO�DЦU�3NB&{UN�q�mә �����J�t�'����r�$��O��'����^�9����S�N��"B,&R=��?����6N��c!B� 00@7M�O�SS���V�~�2Q��HƵN�����^ ��I^��6 E� ��a��?:�M)�]�N%���]�;����%�� `ģ�"�X��O�x4�'�����䦄Iа`�a� 
�P[!�Sܘ'�b�'T�pӢ�+�pL�'�U�	�ΠJE�i>I�����.'��L�{���������mݟ������O0T���ן��I����"C,a��Ǐ��h��%�TR��1FX�I5�@�S��,Zc�GD�'2=�*�j�t2�$���1�˧a�q�w�<p���$� 'w��Q�ӑ~�u�W,�;�򉉀O3(-�w@���N�`S��c�^�S�f̻�OiӨ�'�d����|��'��''�IR�L��H�f��7I����'�(����x�.0���!
L�	�'qB=ғMF���''剔7� �30�ח"���k���oah�zV&JR�`Q�	ퟔ�	��;XwX��'E���� D�&��d����h�:d��{ShM4[�D�A��х�V<J���*��O$]��L�̱����
%J��d�+c��Q�/���x����2	(�$����\� 1��{r�%��ͺP(��Cj�HT߹U$������?iL>���?	����+��&jM�\>���[!�y�%z�JS��	d� ߂��'�7�O�˓��	�\?y��7,5�-��i���9C��q���ƟX�QL�ڟ��	�|
%�A/��@㎁A���Q�Шk���Z�L!#ŎT��gB�)��	QԩHuF�.C2��4��7`�V��3E�������f-`�KX���O2�xd�'�W��B%��@`T �K6݊�h(�	ԟ��-O� �CՈ]&$�����:u�RB�I��M�)�v��E���C���SpJ��?a,Ol��2����蟠�O��� �'����!�'��h�i��Bt�'�'r���� Jq�HX� �B�û#���'��	�3W�J����T�9�ܱ@Bɣ{��?r��ؠ�@�t���H��)��!��~���7��
�u��ԋ0)���4\��A����Ʌ{j��æ�+��i��(`�2@��A�P�e[149NQY�#4���b�@�XI�0mI�_�2�[1�^����/ғZ��a�N��>d���I����%�i���'���]�0�j%��'C��'�Rk`݅+SAɬ`;u�"e�:i؀ڄ)�#	ku��<t���w���'?c�xhw������c_Y�vI��Ý:s���m�v�!�f._1��L>4a[089!�
"l����$���?�u�i��0]���,O�$B7g�z���(ٲMI�Zt$"���� �D@�#�����`3*z����q�	��M��iNɧ���O��ɽ^�J� +E1S�&L�1f��X���H�IʟD����([w�b�'1�ɟ9>�j)9PIӒf�<�V,��1��1�NV�杸1��證���#���Q����ƺ�C�� �6L*L�?�(
�M��ep<h8�����
���'G� �fd+����O`l+A�X�`h��F�w�$d C=!j�a��$���I؟��?I6 L�\]�I��aZ��8�n�e�,'���"A��;��D�1��%w�l�r��0扝�MK����i]�@l���I.��=�T'�8rrNX� �ƎIg�E������B�Ɵ��I�|ꦁϭ^����Nrg~}z�i�9�FYز���
�a�N�����*�F��Ae:ʓ8;|�2���j��4p2�#%�'�2U2��@?H�bTR���`��$��}f����o�O��o��M�f�ʇ��=S�o�'����(Of��<�)§f�,�Jr�Gk�༂p��'%^��y�vN��P�84�F�K����EK�4�ҝ|�K����I����V� �7C�a�MI�.̜B䉝U��8���}'���� �Y�lB�Ɉ����	�>~dBQ��x�<B�	�?��4��MQ&H��&?B�I�P�8)�ҍ�=x���p�N>jPB�Ɇ2:�C��=X ��k��_�JB䉁l���d#�?3	��Xь<>�\C�	 ��VOLh�F�ʧg-r|�C�59��X2쌇�+&&��"~�B�p]hx!#$ܛ��xa��7@S�B��3���u���uN�a�g�!_���vAD|j5#_55崠����1T0!�d_$�ĭ��a^!>;�ub�
�0!���*�QY$�Q�j�bD�d�F��!򤇲�d!��a�x�{-	T�!�č�F0�ʀ�|���)�!�Z�HzBŚ����ɾ/��І�,������B(�^���Nph��ȓg�~�{�,Ym�i�v�,�,��C�<j��M4�ib�/  "�V$�ȓ-��� � Rw��!��]��zO� ���+*L��GLF�j�!��&#�=yg��4�#�.F�1:0�ȓ,t���fƬY.�R� �N?����/{�
�!(UB�����*�x��IB$ A�A*A����mB-����d��� sC8���E\��&H�ȓ V�4*DcسW�uQa���u�Vчȓ{I�s���>`�ku*�Ffp��9�謪�E� �@ɷ�W?aE��S�? 4�i�CB�x�E	M,L�
q"O��H�IҕҠ䀃oָ2'"O`���NW���eC�n|Xa"O
����;��(@ee�yx�"O���D>���j�� �ݨ9�"OxÆ�R�i�|�(BK4Ͷ��7�'�.��rǇ�b���B��O�`�=٦ߟ���B�<�{3�č=� X'f!D���'D�b:�[O�lY���5I��� [��G���u��
Y�m�c�ʼ���<u#����H�,)ir��FX�XP�슧M�Ԝ���W���H�Ȇ;$M{����~b�Px�6��$a�O�H�Z�#V.�Fx��U9}
�D�e��j:يa�F��HOzmP⢍Aز�0rg�?1W;O�葦g�.�<�����6N��f�!)�v����#)m����0v\�$���|�j�Xd�	�`�&
֮+�0SF-QL5�	��M���Op�R�`��\cO����+L�lM���
��9�'��A����3OH�O��GV�`8c�'K:6�C?9�E�O�@��S�i�G��֤a:�w�T��n�}>d�/U�0��-�F�,��]}�L7H��gi�X��Ο5f͒�J�����x�f�5zk�x!R$��p��M3@���|t�-o�<��D� D�����,ғ�>�e���T� �M�O��oڅ�M���T|�t\���ʏP1��°E��^�@׵L_���D͉su�@9��R�k��;֦(|ܛv��v?�����M�4u��&�#P���i>��s�Ya�dҤ;�(eC!�Fd��-9%�Or!Ae�p��1h6��p��k�d��n����3�8<���ڦQVm�y�f�~j�l��.���a��%wC8�錊u ���p"Tx"yڲ�^%��3ǣ�9Uk 	q��T&t(�m�>�(�t�+���t�P�ϕ3S���ic�tr�$�g�~�1a�E�8��Tj�g�'XuJ��U�.��J�&�<�P ��E�d�^D�A߁t�\�	0��$S��6�O#P7��
� �aa	�n��\a�D���^�
�<R�Y���5ְ=�C�S/#P��p���mc:]�SDK'}K���'$������O�,��'1L�K~����yhZ�ɖ+��0�hC0cU9B=�	Ó܅�A��Y+��[��-p��e��ڔc��@����%��8QX�kp�Lϓ[���/K��Zwӎ@�Ǣ#��݉V�T 1��	�-e]��G���e�DX8㧝7��	)K�t�_I���!�ZVw(b������Z1�����]ZҠ�f��A)����O�ӡ-�(.�PXJ�+����3$�`��	E��⃊�ઔK�Ơ4� Y���N̓0�y�T�'��9͓`Up,�o�a��x�4!ǧ5�����d�y6hS2#�'	�r���O�MZJ�6�I@Hq���}|�-d�����h �?Y �4�Ӻ3U"�vx�S5���l�@��#hV8�<
Ó)�e��_=3��$�24�"e�=.��7��i
�ёB([�T�������p3�2Xa��H
=i�t;D�O��`q�!^=?Rv��B�
�wͤ�J�O��pw��5o�Hc��	<h�,����>l���C뒣�+�&zf�y��O�
� Ȝ�6�1�ègࠋq��O������[�T`��� Z(���1�ZI��Al�����Q���	����'����l�Y£�@&NJ񳣬/Y�l�2`�|�e��Ӽ���J*/M��(�	<�y{��_~bP6p����:���(�.f��]Xr�т��|8�l�{�0R�Ҳc�ځ��+ Cδ�>'��M[�`n�
C,F�*��8�S6?�F�(��g2�LY�h~��d��Vġ�vĠ/��I
!��(1�O�L�J^�M�b͓�˚t\��?1͔�1(�)ԧ�QW^��1�PL���ҽ��q�5\O��*Y�4piz�lظe\��ӆ�!�ԋD��7H��Y��'��Mɱ� #� }����8���b5"O�0Б��.?p5���^(V,�Ad<,O�	ht�ӝ,X0ԋ�F�Y+��PP!c��F<W 	!
`����I�B�P��J�|&0[�&�~� e����E�'��<�|�HG��ILV��a��E�B��a��Y�.6��qB�u��9�,9ʓ3O��c��I�n���s�5k���'-P�k$OL�:�P��$�[	_8hH�
E�rĥ��ō¾���ɥv��&��i��0$ �nc�]xe�[�-���J��=}"��-��a�2�Ov�qbg��5+�YRu��-I�R"OZ<	�K�$V�}(��B"|��u�2O��O���"T�gax�2kE>�qw)^?�'L�\҆Q�y2�Q��H�]�y��ɕ8�B�@��$�.Q�bߠ=�r�R�-��f�����Σ>����m�4��O�u���H�g�?i�'j��Z�^��thU��(�p���M�&)tQ�l�F�J�u�u�|�'�ؽ��H[^ VxA,B,oJa��ͫ<�D�hU�WD"Ŕ���d!f����$ L,J�\�wlm��ƤA�1��A�)�4����0i�����	��7�,��DOX����_�վ �ߓv��v�҆w���x��W$x���'��ԛ$>��=i:����"��Dd��?�JۭT_,(�r@(B( �P�2�OP8�b �Vh��C��^��Ě#m��S�r���<��[�yR��;qI�G?����K���h�� ֤�tMTUn�5j��zp�i�kM�WDS�J�V�h��68��S��߁Ғ�=	��x�T�j�� vmyjё$�[�7aH$�b��!g����'��3�h�V�4���n!�� ՉO��$Bbĺ��W�d>%X��M���?�@u��q�p��4f�>XsOA/7���/�|OHIE{"�I�OV��Q�w^�l�u�8HN��+(
x.Uc�-߆`���lٚ ��S�'n��]�����!K�
�G�8�0�7�b!�d�I,�A��I��As�iD��&X���M�!/\he��� �w���iX4�ƍFJ:
1y�D^�f�X���������o�����C�NJ�	&az��-r��=)aS�z�1�D�t��y�S@�̳��!Z-@z7��  �0�@��p��
ԁ7ӊ N?㟘� ��p~���"_.|�Ĩs���L�q	�k��mR���c,W�z���3�E&����A��9B'oJ^�>�lڂ\��c2@�hў��1)f)0�,ϛ`0�����,�\\���S�(����� &�ek�ꊖv�D�`�UX�`Y�S��Oz�(�'ס{ӌ9���͟=����ɲ^����U�_�#7&p�����,��s�H����&x$P)��k
z~�!@����y�Lm�C
�2h=�ɮ���{��p3'`�
3���C��gբE�����2�B�Q�j�rR%J4l�q1#�Ox��T_��ͻd�^��f�.}�l�!��W����	-&H�Ћ{���i$�T�Њ ?7��;�NP:'DXPHC�]%H� �q�'����'���޾5�ZI�+J����4c�}�a(��Qc�����X���,�|��퉦1����˓	��QAD-��a�P�[�$�c�`��E#@�8Z�	�!ƒ3RI�	(pÌ$�O� pId�X>@�ā�咇W�bH��\��O\�V�Ã8H��@���K'���b�\�D���	8h����*n���9�
_eR�'��;�O1%����,�^��J?9��gw85A��1e<
6��*�{p�K!`��=P��R�$n!�E��#�(4C��%�<2�0[l*��8,X)qR�\�1��lW�*���Rq��@�e����!K�J�Fy¥��-"�)G��$E:�%�;�*)�U"K�V\Xm&��Y��x�í�����(���' J���t�T�1H�!Pɽ<�y �슻�N$����)b� ����7$B�����/�$-�Eg	���V�;�Hy�я�����rK�p���dUBC�O���y���?|"<�a-��.`��e#L�رS#;�"٪���T�#q��:"���c�`��B���&��a��>iC�5����Eʄ�Qꐪ6�@i�ӳNH>�Ch�1(���@ ܠV1�<��� v���*$@@k�Ó�>�'�k�i�])��׿M��s(S�^D�] /O6��W�M�z�r	�������/9�0+Յ�	^�|��iȽ�����K�rx}�����^���eQ�(���]*y�f$K���*[y��-Cխ��/�R�>����(a2D���d�.��7��zp��Z�*A hB�OX!Ҋ��I�V����ٵFZ�6���Q@�$�O�����̲7�Ǩ=�$�i���("uL��L�ٲ���1=����Mȍb���)�����`�YL]����Ry�����/�8+|z�A�m����l	�w�p��nٗC� Ś@c��	A�Qx)�x�}x�Q�-|����O���77��cd끹�v�
5��"w�pqGI6����"yKD�����AY.����*JÛ&g��?@TӶ(ʇ�M�ݴ!��Y"f4�D�?ט�2�NՉ�`�8qfyIҪM�}U����[�6�����H�
'��vʗ��lbFHG�����''|�H���O��m`B@W�QV��\!����T��l��7fNQ��j^�#��P��$�����]Fc\�c��Z�6��fV�C���'5�lZ���HJ���`\�K�̸��Ra�5`$4� ݒG` ���h�VY�J����,{ �p?�O�B�'���5���v��W�RX � �T���Ğ .g�x�&U�E�< $@�[�ax2��!&z�����..���c����yb�G/)u�͢B˺��c��|�g���'xL08Sg��9�pm�DnPr�jy��3<Opl�@fA56zX�1D��q���:v��
&�l��ɀ_G��:�kǱ]�ў@���[~l6H��o�2� h�0"X �qRk>/~�,��͟�W�Dr_[;�'?}1c�<=0�B�N��j��|�a�F��(Oh��f�}��@�F��*J�}�eW��%�6P l�"`�%9f>��Gۮ¨@1��k�6X�g�O�4@���8��iͧz�u `ڲ��c�D?x <)�wH'B��,��ڸfH��ȃ���O����,�Z��ЯX=�`��;O(���(
����JV��iݕ)O����s�=!�o��*�Ԑ�%�P?5~�:0��3R�y"�@u�
�x�����s��3�X\�K&-��!��D�O��8�'�eЖR��;ֽiuX]�ӺÃț3}!bhI+�f��b�""FXM#,�/�O�������&��Q�'��O����k�1���T.׎T!��@�[
k1�e��er��J+��O�R��'̴�k�F�dvt�����A����D���t�BbOW�:8��S��M�;]��
 �J�R���8c
7Z��b�M\�@ �(�'&q��cQJ�)S̀�:MA7�/J7����b�����44�P��pKș!��)�Y��K'!��hAEɗ�1<|DJ�4�O�x��+B Ҥ���<(�B�w�÷ap�X:�A�n��ȁ�O���p T�]�Oq��͛�+
"h�f��9� �e�	!`7,ș3!G4L�E����!bH���c��	;(eZ��!��:f'�\B��L#?:���*Eجarj�$�5�Aay����� ZС��^:�YHc߉"}�Pa�"O���ؚx��bTL>�d�R�"O0x�q-�$Yu��W��;n�B0��"Ox��O	�,Y�P�g#��"�X�"OL��U(.�hA��$
/<��8 "O�ݓ���?ehDB$ğ5I$y��"O���;���c�a
u�&ј'"O8p��K���۶ ʘWC
�:�"OR`b��Vla7"��r1TL0�"O��V �,���1A��+M.LT��"Of\r��2G��F���Y��@�F"O��Ca`�vi��)ǿt��$:"O�X�֠_�%��3����F���"OЙ#"G�r;~�SEB�u�z�H�"O\��?f���g�*h
�	�"O�
0���j�IjUg�)��{#"OF���֜�>鉕EèG�\M��"O��������Te�QX�Hs"O������d{0 9F.,ߞx"O�`��Ȃ24ʰv!��<I��"O���Umڙw�������,=*�"O�	ˡ��z��`2�烅X�z��"O8<�D Ej`&\:��1�"O�"�D&J�0�
�֡7����@"O451� #�J�j���7Lz\w"O4*`LE�H5��Ddͧ5�v᪥"O�t�D�� ^����eY�K���	"O )�4��	~Q���7 ��L��"O,]�6��}���C�ʶ=���"OT0
rL�������\'y��"Oh�u!L�(Q����l�(bmP ��"OH*ք�:)��	T�Ŷc�"h�"O4u�Թ:�P�� �^̩�"O:���n�-i��2CI.@iJ5Ӂ"O�I�Ù��(���1M�@Iyr"O|��+��@���' Z$�Ƚ�a"O 6��u���)�%���`"OT%���_=|�����F��9�&�2�"OP� �P<mS°k�&�p���"O0e��/�p9�X��f�m3���"O$}J�?Af�� �eI;��`"O�PI#e�a���م۪X�,��"O�0���г8 |ju'`�V(��"Ol%�B�Si���V��/o�HS4"O6���A�#�l�A��a{����"O�Q(,�#jO�u�Ei�8VV�ʰ"O�yq/�=\îD����F0$"Oz�:�C�$&<hu	���1}��6"OD� �S:O�H(���3e�e[3"OHD�I I@a��׆yW�[2"O���PMQ6�(Q)V��B"Or��&RW���)�]�,�!"O"�bS�U?�te򇃭gr�x�"O�d2��مBsв�$B�1eؓf"O�d��Z�9:�ͪ�d�*c��8r"Odq��*�jD��㷣:3����B"Od�ɅeA��P1�C��Z��4"O��1�@�qђ����&Х�"O��d䜘^��I�.�6t���"O8M�A��u�����c�ay�"O>U � �%%��9g��Af=y�"O�A �mK,	pEY`B�K&$i��"OZ�H�:%��(IK�.+y��"O�� 2 �㒣!$'��@�"O�  �k
J�!z�=s��s�M[�"O@�Ӯ��vI��@#o�\�"Oʍ�s��'	L��E�ۑ.��"OxA�!�O�_M��ґ�1��y�"O�(��Q�u���iR�΄.���"O�T���O%̺M��k ,�����"O:��BH�>L�N��+Y.,�Dr�"O,ئ��X֌<B�	��8���"O�PDE�#B^���H��S"O$�A��O0P���p�K�p�J�b�"O����_�%��yu�$�ST"O�S�nˊQHRy@���*�v�W"O�j�D9b��2�Zi��@D"OzE
�*�_�:�I��On���	�"O0��t�� ;,A{�l��\�(S"O��1��P�V�*�aN��<�r�"O�i�c��V�УR�5�6!v"O�a����'�`����� ��A�"O���vG�SQ���G(�����"O���CѮR~�<�g��	^�t�b"O�D�@LK8J���)�<�8���$!\O12vd�*C�� i@. H�$��6Oj�'h�/L�������u��Píl�<I�K�3��(hu�z|>�;��N��d�'_ �1��ƙog��@D�mTR!��'�<��+H!��Ļ���Pdv�q�'�{��X	�t�1͞�B�08���d2�'d,< ��Iɭt�v����N}�?��q؊���Y.Ų4�$����ȓw9�-pB��,Y󚄙���P����<8���=M�0�rcZ/z4i��~s���w$Ltլ��5��p<�ȓr����C&Y�
�X�ݓdM�ȓ) ��9�mڈG�R�����4#k^E��?�ډ ��/1� �"��S�_ː9���A�p�g"�(�&��-T��܇ȓ.�4�e)N=�¤��U)n�P��ȓ�xu���4�
��f`Ξ uL�ȓ.��	����AS�U�G#��M��ܘQ������`�Zꄆ�/]pd���y��ق�傤N_0��ȓAEB���b���E·%u4H��E�(�Ѣ�K�
��R�KX��Gy2�'�|�zW@����cqH�ʺ<��'4��;Q$�* 8$ܸD-�0���'t^L�u�� \b|`2��׼.���'ה�c���)����e�R6~(r�'�f�y��_�@��L�D	<�`�'OΡ���W4�(��et�8�'���w�D?w��D��k�m�~�O
�=E���׃����Bǽ5N�ꥆ�y�
�1��`w"�-JGf\�fH����0>�P*�*IZ9�֎@;^�t��G�p�<"�G0}�X��W),�-���j�<��-u�^ix�`�19����Vg�<���"J�$�eo�vU܉��Mf�<A"+��>
~@���5\��H!�-�{�<q��D's;�}
g	3]UB�`�]P�<��--r�F ��-�."GJ	a�P?���E�бr�#�8�^�n(�ф�SdCe͚��P��\��Cǐq��8[S4TRC��?C��(���?���B �	�aݡd�,P�l�~�<��g�*d���WT�t!�`Ts�<� i��e�.E�x����Eylm�e"O�%���D��õ��<YtK�"O�Ur� �9Z6�A@iѭ;b^��4"O��k�<��K��o`��"O�thD��p���7�6"L���"O�X��'B�{
Ey +�8��"B"O ���$~30����˹eD�r"O�(pcǄ�n}��G�#�����"O~�����,La؅Fǁx���3�"O~AчǎJ0�Q�'f$2뤉`p"OnY���G_�p��C�:�8a!@�|��)��E+~���E�:'D����
٘\/�C�	6E�$rD	O|��K���;xxC�	+{�De��Ť2���j�GGw�VC�	��CI\�/�j�(��W�V��C��/w2��hp!tl�ӣ-ZW��C�8�ř�E*4:�0�圫{u�B�	<tX۵"�~�֥R@,�;l��B�ɤj�̐Kţ� �n	�V��x;�B�Ib1�9pe�ځo-x���C�~xB�Iy"b�y�m\�[��Yr� �C䉖U��[�#�޹B�(�<�>C��&9F �j�P�!aʅ��/� W�<C�,)�l���!���I��r�,���4�I�h-
��KO�xY���ǃ�b�C䉯ې��g��,�l�H$��J	�C�	�"E�'�M�2��F�Z�JB�I�y�\US	+�ZHS����W��C�	�D0��F&N�X�U�<0B��'� 4+G)Z�@,�Sd�>C��'\sȜآm�zF��D�R7A~�C��"s�:�3%�̌h6���t	ՉnM�B�	�8N��g��P'l9�&�!$�B�I&	�N�(��ɛ^��1v�R�&�nC�	�o2EX�B?Pw���L�LC�	�]��h� �ޭm~�qk�[�>C�ɏ%&������ckpda��Fo�<#<!
�8�t�ݶ5pRwZ�  ���>R��A)_����� (^����G� ���љ��sч�"]б�ȓNݐ*�+��]Wf!Ko�=È��ȓi�17�.�� ��G�e\IE{��O��9�+�(e��%�M+v�l��	�'�4��g��?2������y�̍��'��PTl#{W�1���Gj]����'T&h�#,�?%�6e�b�g>�i�'�acH�7vb,*և�pT��� �5�yr�Q0���i�o�4`uh��yRg�9�RC��-+2�;b��yJ¼Jn�����I�
v���t�˲�y�ꄏDf��u*�{D>	y�K��y-:/|�i0��B{�A��!�y�� h����ϋ�8U�h����'ў��H�3��%� � u�۔?O�A�P"O�r���a�4u2�
�%F��&"O0ہ
�HAJ��ŃE��r"O,��!�۬C�2�C�I�h���[!"OX���aTal�k��D+%��lR�"O:�#K]3B���Y�n�5"OZ͈Cʇ�j
2,�K�$-�,s�"O��RB�-P�
�Qv @�r����"O�C�%H|����!B^3��T�"O��[,�5U�$8�Uj؇X�ƍ� "O��s2HX1I��I͒2�qR�"O� �Y��gژkPsK+O�j��W"O�A���W����\�Fh!�"O4붨�/
+0�#ᣔ�nR�A"O��w��'Dj� s�Bʤ�J�Z"O޸�OW�F���@�QpveA4"O传ȓ�,`�RMϤSw8`ic"O���e�5KX�Iq0��4��0'"O���b�g���h�@�w����"O�}�qd�&<����XA�|5��"Of�ct�Z��`c�Іg�,H��"OF���ś
^_��ҡ+��db"OV4iG�J)X5����A�.vp	u"O~�� �@z� �	�u ��"OD�!�B�6<!�T1��>ax�IP"O��a�îa�V,C@M�Y�"O�e�oWk���퐧)pq!"O�[���.~vj��d�?�F��c"O�����6e�F";1��\c�"O�4���]*5��=+���jV�2�"OP��ע� ��� ��!	9�!X3"OQK��lb4526�E�M1����"Op�� ��"F�!`j�����:$"O0�7��e�X�	�Z�l�Z"O�	$�������'�> �l(�"ON9��G]�u⊌�"�C�S⒩w"O$��$�\�`0`�E�!�V�W"O��1�DƏM��H�hؗ�r�I�"O�y[V��8.Y���T��"v̂i1"O�1i�C�:T���a��/_,n,{�"OB$a�o�o���"$H!$���"O�5A(�UR�����i,���"Ot����R���9�#x��5�W"OP�ґ�ڍ+{��	���-l��I�"O�	VH��v���eP$I��-�"O���b��2AeX㢅S�]���@"OJ sN�3>�|k�ፆ&�" ��"O64�A�&v\�ĉ�E���I��"Oni���ĩO���$-��{����"O�-��I�-���q��1A�"���"O�����3U���s���C�HQ�"O2�h*�\0�q :�hh�"O&���I_�< �ѥ�<�<��"O�+�+����Jed��h�B���"O�e�D��3H�8C��M��<m!�"Od1�0��+D�<��K9$�
V"O�����9 ^0�1bM��
e��"O����g�3T��h�AZ+~�M0�"O5K���#O�x9��цQt�c�"OB(��I�{�p}���ڵ5d����"O��1g�&������)� T@�"O� 2�V�Z?�!�)��>}��"OHxC&��,$�J�i��~��3q"O��b2(�7A��e�w��8a��"O��cĩ�y�XxU�Jdg,���"O��J6u�b�[!�
a�9�"O0Li����8b�Id6ԉ�"ON@�&CW�k�V�" ��Y*���"Opq�I�
n4�x�Rhر#n8|��"O6�p��%a�J0q�iˊZ�j�Q6"O�5��*\b`���Ӝk����"O��E�Km T��FC�$���`�"O��BӨK �;��U]�|�Q0"O-�퉣tf�A��eY�2����"O���@-��`D������9[���Q"O� ڕ�)�)X�0�؅b���2"O0m�!AJ7-9@\*�B�x�
,a3"O�q�*̿>�XY��A��B[���"O��3r�;zx��ւ͢~�>!0"O�aI��U�0�ۄB@ Ÿ5j�"O��Ja�H>[ސ�{R�g�<� �*O���p�E�7ސ2 $ߐ[T���'�^e�M�9."��rZ?����vG4D��q� �&6��
U>���>D��@�h[+FX$[�b����cE
0D�xH��ɛY�\�`��-j�U�E.D��CB(^�1	6��0a\Wؽ��1D�|р�s�8EcҧV&�]�`0D�``�)�0�9DK�[,��j��,D��3v��0��(Ӥi��3j��(��%D�01���#fM��쇝
ƥ#4�?D��I���;zu�L2S�[F \rca?D���C��m|��s���
 ��q9D�,Se��&+��Z���l���7D�@P�ްa�2h�TH>gBAs+D��)�$h@�spoF�@`d�+��'D��(D�i_��������ň�yҨ��1�ҍ�1	�03�~ ���)�y�M�bLm e.Ҵu�ժB��y2hG�.��F ,R�2���y���/0��,Ö@y0P��yrf�1p��H��MM�q�D0`���y�"R�Sh`�e߉se@��&��6�y�f�#;H�y���M�7���CS%�:�yL҂Sz]��P(jsgd
��y2���c�����B�/'�a�CLV�<A4#Ɉ*G��!��$�D�C�Jp�<� ȏ |�@B�*J�`�z��2E�i�<�ǫS�	���?������f�<�B@��.�����$��`��\L�<��	V�)�����$l>�B�D\r�<�cA�+��	+` ڦ3���R�<1&�^���� rmY� ��-i��e�<�E�Ƶ(z<�9F��}Cnl"��g�<�f.T03����Š��պgM�d�<�F)V3*�x*�P�9����Rv�<�����a�@���,�;�����s�<C�ޙ6"!�b� hFu�En�<���Q�m��2  �:��(r�EMR�<A$�] /s&��P�P�/#b���O�<�L�u�4�g�.b��(����L�<I�?n�ލ����z��m�p��D�<�D�E�d��xkÀ�<ĺi�nK�<��n/(~��wOʺ6l�e/�G�<1gfȇ:�l�!�D<<x��[օBA�<���	"��qC����K,p��_@�<� ���kW��R�&��T���1��z�<�e��P�J������e��A�Hy�<��ʚ7|�����o��xj4LCO�<���1b�� *@�V�5���o�A�<q��2$I"�AooI��i��y"Qrlܓ�@N�Ȗ("c�e�<'��hu4�(SC�G�ؽQ�	Vd�<a�nV�Ȝ,����O�0��M<D� ����2eT���P��i��7D�xC�*j���Ig/���H��9D����悻{��(s f��[��K��=D�|���P�a��H��E��|L��=D�`��)qL�tg��R�&&/D�� Ry��̌/]�=;FHH�J�D�;f"O<�2�Ȗ�H�T���-�_���"Od��`��+}٢P���W�cEMB�"O�q���"$�t��U@\&0�9j"O���D�4h�,��Ɋ3-,]۰"O(���}�ܠ��֮����"ORU���g�t�������X���"O��+Q%�%X,uhܘ�"OHQ�DJ�K���$'\�kY�ٹ�"OH`A�@�!h�A�� "O�=��@
7H��<��'�J�~���"O�UA�'�-���vH��N�!"OT���,��~]�����B�Y�fͳ$"O�<�oA*����X)/��|Y"O>�R���/*���f�A���j@"Of8��C	E�F�����!�"�"�"O:I��Nz+4��ŋ!#��Ma�"O���Ї��q���,���Ȓ"OLC1HC=+
걩�
U�2��$��"O�I{���?nj��/T����2#"O��ypO��G�Nm��o�,�^tP""Oڰ�ٱ���
�ٱ'"Ox,��g=:iIp�] ���"O����%�Qi}�0�p� ��y""��c����U�?����!�/�yBD��O`�hb$�+���	C+߯�y҉߳�r��� `E�QiR�W��y�-M#E�)C�e��Y��(r�$��yb�ܫ%>���R�MF��an	�y�%�'�N� q76�Rq�Y��y�k u�HL�&-�>2S�@
�O��yR�	� �0�ȷ�X�x�ڱ�@@[��y����>Z��F�nB����
��y� �\Fɒ�M�c]����8�y�KߟJ�6y�`ѭ'�j��Y�y�	�+*w��㑉�1%NX����yJ@�.���i[7$��%�gaC6�y"BՈ����A�O/�5b�mM�y2[����Es8�+w�O#�y2#Ʌ2fh!i	g���#�ʓ��y�A"I����,R/C6I���8�y��ҟt���pC [�����y��3V6��O��dX(�ݯ�y�MR�V���6)C���u�f�yMR.�e;�b���!��&�yb�5='j��Ǌ�5U�]�Ѝ^��y�N�w�H;��0t��	�y�.ևwh�S�阩s���{&��yR�ʐkؒ}C�-�Y��r&ٻ�y"+'P))��"]~�ݹ�Eð�yH$'�"���NS%B`wW��y2#6�rU	u��|� �p���8�y�fʻ�",AdΈ�t�X�b�,�&�yr��t.�XK"���mb���+�y2(�(f,Ԅ0C�E`��j���yb霯5�RiK�e�?orth��Γ�yҋ_;jJ
�	g�˨9� �:�ѥ�y®RKb՚Vi��1�񬇌�y�&yht���ԩa�h=��kJ�y�'H.h�g�F�n��y+@��0�y2$�V>6<a�
�_���CFL��yB��Qv�9���0[?���R�͏�y�*�( ���%^Nɠ����y2 ,<��i���N�Tx��%4�y
� D���� d�c�bU��4�"O>i˦�1a�.Mj���
7�b�K"O�8��n�
�A���
Z��"OVX�놑rx�:�nĈw�~Y�V"O$(��(�4���'�
��"OH��#�7��c�cP*%��-JC"Oq#��5���B��ȭA����"O,��w�J7��0u�U
mZ�#�"O4�*�+E�h�!:zY&YX#"OZ��/ 3��pZ�f�!r�,0��"ObI�s�$#~q�Յ�4�{�"O���A��5>~�iA$զQ"O���b���F�0t��n��Mru"O8]zE,Z�u@%�7��\�"��"OP2���cV�Äj����� "OFXc��KM�b��*L1>�j	*E"O��Ѥ%�%<2���XY֤�0"Oh)��J��"lAէ�@Z$PP"O�5��fF�,�>�`U�ix֜	�"O��h�ٍV�f$B��Iza:���"O2ī�l&���E�8wlPA�"O�)��DHʾ��A�9@vnlʷ"O����mƨf6���!MT�f�Q��"O&�,�H���Rkц^hh�&"Ot���JO	k�h��]�?Lt-RU"O੐%�� L���u
�1B� T"O��� mߟ_kl�07�M�0\��:"Oѐ5k@�ձ "J�A��"Op�K�1\�L��v���&`�a"OLa	�4``�D�nvi�4"O�����a�Y ��5_����"O��	�bpf�rNZ�|}pT��"Oji��׋��X ��	h��"O�0���g��'�Q��1�"O��R�gM��i@�K�|τ0"�"O`�mW"z,|Eʐf��3�>a+�"Oީ��\�.\�r�ā)��#B"O�X�ɔ�d��c�D�,Y'�x�"O�����K���Y���,Z8 %"O΄��e� �V���4�J�yB)ZQ��٩�g@x�1iţ�yr@�#A��@`0�$�:Ɉ� "�yb+L�S�u�r&
�I~�@���y�@ţ �nhӲ)U����F��"�y�%O�#I�
5D����Jݿ�y"�#7�U�P�ݻ2�@�P����y��5�[!�L����b���y�K��W���3�-�D���;�y�fV�w�.Ԃ�+ǢXXiD��0�y���~8q�v��Qdm��yb�Uea�����~X=Po[��ygՈ#���'�G
f��Da�i���y��� ��X
[;����V��yR�"�Vᤤ�l��Ҷ����y�cņL���hp�Isr0������y���ـ�PBAxt�"���y���M���{ I�o���`g���y�;$�@q�#��+aT�E�g�۱�y2OٞE#���%ƛ>TyUqT�(�y"�����	&�^�D�Z��)���yRH�/_�}Z%�@0hu(�Sj��y�dV6F��D˱/�5-�^��A$�yr,��F}��bO��59�dU�y"JX3�f��EXZ�le��k���y
� rm�6�����ʢC�!�"O���
���,˥!�>�xY��"Oݑ���U��s2��l�x�T"O>3�Q&N�����̀�K�"O�p(�٥P�Z���f��) �`"O���5�I%U.�'.~��l�v"O�����D�/]6�2���.�T��'$����<F��׎�V��%�'�N#G��'u����G��0��'d�-��lU�8�����Q:��p�'�`,c3�7X�����/y�-��'�`����/bVx�a�!�.��':�1xӀ)܈cr�͈O�Dx�'�"-��-ݒ��A�P�
�K�h�Y�<�1a�9n��$I�B�?
��:�'X�<�'��:�z5�Rh���2��[P�<qEM�>u�-�`.2x�V�!��c�<9`G�a�T���b��`�r�8ElZ`�<2�>�#�ˏ$!�l��	Vs�<y7"?��BB�Z�7ʴ��Řl�<w	�NQ�KFق9���e�<1!��1�%���R>;�J��$Yj�<QԨX�n�t�cvm��"%�"�i�b�<�� 0f�j�۳��/^�Τ�f��d�<��b�;k�,t�ӅA�m�L���eB]�<)��)9� � Rk�0��yh� �c�<٣��t6h�JW��1�L�w��\�<y�B\��PF��m9���s�<y��A�5:t3dg�)��M��c�n�<����rH��Ԉ;(*�CI^i�<��FG�O�||X��B9�BUi��Vd�<)G�۫��A+��7l�Z@��`�<�p�V%0׋_�6NX\ҧW\�<�g)�.��������`
u�OC�<��|�B� �h�0���#C�J�<�ӌ����B��%�I�B'Zp�<)��e����#P�o0�0��v�<yP�nXI`5��:��I�qC�s�<�7�I�8�Xz��C���
R�t�<	 ���&�PPm!�$drcF�<a��\�L���'G,�����E�<��eۣD	�-�G^<΀�9G�X�<��煩03R����/������P�<�$A*@wD����%��Q���N�<y�B�}�p�bF�wL�%��CR�<I���(S 5���1�Tp��G�O�<asK�'��Rτd{~ႅ��u�<ɂ���y@��(���>��u���u�<�@"S#8=\4�'oL�(�����y�<Q�	,�D�!�D>Sei�ʀ}�<!�M��4��(�i
j��}�d��|�<	��C%He�`�Qf��5C�@���{�<ᆏ��lb�3�KX"�љ��b�<��A�8�tő��-P�L��e�<���]�lEa$jЧWX�BX�<q%��DߌM*� �:���(KW�<�wΆ�s��x�f�ҢA�(���}�<ɲ�ƽm��	ɰ���D
4e��@W�<!A���\Q�,�VG�%���UC�C�<IcL� }��eo�R�0�3�U�<Q�
�[n���@�IWL ��k�<!̌*��q��>�Fػ��Vq�<I6�+̆�2d>҈M�w�Px�<!#��>��(Aw������Ww�<� � �ud�RV`��W=G���`"Oh��&�]$L����=;w�X"O����*y1�)E�`g�ܳ"OvL���5�lҧ�;c�b1��"ON�)��M&m��:,ͪB���yb"O�L�GKS�..�T����v@��`*O�D�Bc<��I`��Gަ��
�'��1#''�VMPX6*@�;�6��	�'���cfHJF�b�(V���:�e��'>���.b���:�&�B?�9�'��8xT��6c��D�⮔<����'v^@�V��_$m�AD	�.��(�'YF8A6��}�<iO�+��hS�'Vn�h��Ⱦ{t&9�C
�#��k�'aK$��kR|�3�սY6,yj
�'��ذ')p�1�C��$�E!
�'�$	kRF׺j^�P#K�-�@���'�ݓ��D�6=j.��+��Z�'��!8!E<L��LC��U�����'׆@S�A�Pώ$9�(��,�pm�'�^U�/�?�Vh�G`
�t x��'ɶ�s��&X�P�Y2ͅ��jex�'e�Y�4���f)� �`�M�	�n��'>L�x%	4wxH��٤O⎌�'����e�t|h7��L�����'9�e1^ p�ǝ�m:6�b��J��y"ϝ�+i����cI�m>Dшc�S�y�͐,'��l���c�l�³���y2���d�o'X�Y�#��y"L��,����"��k�����#��yR��Cp�D�A���Mz���( +�yB�D,���e+��r�حQѢM��y�Q1j��]�2��qp����K��ym�~^X���M��c�b��g�&�y�,\����A�^IZ�y��
r�<�!�\ ��$��	(��9�CP�<9�/M�*N�Ha���Fĸ�FH�<1 BC]�@��&" ��dx��N�<�S����r�A�8sN���a�s�<aam�e�0��n��^$�gh�l�<١��"s��A����
h�P�M~�<����2���¬U��<�6`�y�<ѰR)@$R�{c�ڹVn����Za�<�&ӻ7'�H2��X����D�a�<a�Cҭ1O~  ��X9SR:��E&a�<�w�W�w"<�[Qʏ�)���a��U�<9ç�#�nm���@�w*n���Q�<ɧG_+R�� �a\)I�� ;�I�g�<��W]�
���ɢtN|��Vd�<���#�zU�DZ,4B��@l�<q `�5r-��w)��[�rԡt��i�<	%�B!t�)a�D[ߌWvC䉴Ksѡ�@Q�}i&�3�A	�o��B�%�=�ekG&}����c5H!򤛦Ae<���fTƩ`QCޠ7!�$L�I�8҃��PN��r���sQ!�ϕD����FϾ=X�P��Oo�!��y���#��;e�!��F3ri!�D9
e\��p��p���#'L5�!��íB�*=0פ�[�1�E��!��a���-k����iç3!�-?�dt1N�*]�t��HS�S|!򤄮m	�d¡	�&�!"I�] !�+ � ���p�B��w&Z�!�� ��d��9���A-�6��;�"O|���"��b�LȀ��	B�$���"O�d�v�&*��dP�L/zb���"O���m0~{d�S�� Q�պ�"OT�(�ʃ�iX������)�@"O�ec�鐼4F]���^�.m��"O��@,Y�>�#E3b.��v"O`�E��2��TA3ᒽ~h���"O��Y���5#�Y�36���3�!�Dدw�-;-#1�4�E��4�!���m��tRֹ{��᳋�	~!�DM-Yq�Т�$hk0��7�LW!�dK���H3����\�X(�#X	M!�D�9`E�cǎ�*Q��;��^�J!򄀣 �:t�j��N�M�f@��_!�Z 8�p�)4 ��*Î]�c�W�!�D�.>�Vi�FΠj�L��4/��!����x���D��:���7O�Y>!��3z]U�k�:H)/�3'!�T)7bL-8���?m|���(�O!�ěd`�C!c��uR7�ƁP�!�� ^��:U��+]��)B��F�k!�䖛���L�nyQW,��_!򄚋4�� �$��0xj�r��j�!�S �r����=livh����9�!�dѣ9����7/��XJ���E��!��Uo.,+V*�� �~�3��I�*�!�D'X;�ds�z5VԂ�hL�A�!�dS�6�<�/�.o~��0�h��H�!�D�%@h<q6m�>)~Ь!��*~!���(j����ӎ�7]e�4:4!� �!��^9A#��[r�hWH���
M�!�$܄+x��M��!l�h94@
?J}!�Tya'���Ƽ��Ɏ$ b���'Y��#3��Bv������5����'�Ā�cd��C⍺M�lE��'���`��JnuK� -����'&~�yR��*��H`�Ңf~���'�@!
4$�S�A� S!T�a��'Aa�Т/k9`�e쟊���'��K�<4�h�Ha�,�����'���� �~H`݉�gB���'q�Ja䃢*�����*O�p�'���8w��	f�X*�B�!�a��'�*M8�H�4$4;F"	�zȘ�'S�(���G��HA*�t�p	�'��H���V�*RT��c΄eu�	��'�~��Q.#ɶ5��jU�U!a�	�'�"l�!I��R6Ü5d��H��'�dqV�S�5N��Kc��_� �x�'�Ja2� Y*ޕ��mҿW!ơc�'SP�B��$Mj�끌Qڦ���'�,���)��bS�)�Ĥ���9	�'HAQV.ԹR�`�K����~6�a�'7�Yp#E7o�` ��ļ*C�ظ�'�)��!�uR�D�	Ǎ+����'�8w5Y��H�kʜ�R�h	�=fC�-@�l�ŵ�IҚ�Cmġ�bC�	�1���nN�<O�Y؅_�{,C�	�d�A�n�xp;�&���g"O�Y� �I�V�`5	��@�a�B"O�Q�����!���D�6˪�p0"O�C��< ����c�-=���p"O���NG�Nɺ�#!H%k�E��"O� rm2' �7��5R5B��	O�yA�"O�P��$��":D��`��rA@�A"O��ȴʐH�Z�£�ͽ�~!r�"Oz�3��'C����LV?�dY��"OD�9�a2T��"�)�'|qz�"O����F:]�����O�q7V��S"OB�{V��#I^≑��ֺ�;�"Of�������r��$W�U�@a��"O��[�g:��Ă��5p��@"O�uzq���}|�*��_�-n^9QF"O��tC�;r~�@�wj̉�"O ��R��4g������Gy��h�"O�zu�Y  ��D�<i�љ�"O�9�O��{ʲ50��8Q\��"O@X�7J�.Y��M��!]FTL��"OR4c��q�����ƀM6Ċ�"O��ZA'�7�<7��b<�}�"O��p�
S��͓ǉR�0�A`"O�5ۤ�	�1�:�k	O�2�Գ�"O��:C�#O3���p�Ɓ��j�"ON-X'eO�V.[��^��	+�"O|(�$�آ5L�yH #Q�!��40v"O�p�C�NW�E�N� �	M�y�k�/Zc�8$JH$N�*�BRM���yRo�yqАY�XM�f�ZF���y��ηer�PAȯ��!��"��yr��3 8���E*w�6��͖,�ybFѕz�@�z�\ j�(�C�:�yR�K$;C���$��dP����`]�y��4`V���ŗ'ce��)D���y����-�x _�
�:�x�����y2c)we�t�Q�C#{�XQ;��N8�yrJ�\��3��(}�u�Q�'�y�a/f4LCLx�S4��y�q�܂��
hJ�`�o.�yB�D6
�����l�c��p2UL��yR �ITa�х��I��������y�e��{|y��-;H֡U� �yҫ��)�d��b�Fg�$ɚ�����y�ٝ�� �h�`��d�Q���y��_�P�
���!ɥ^���`�f��yB�L�T!�<����TZx@Ak!�y�*�4���2Ud� �L�:�%Z.�y��܏b�5+�---Ht�0G��ybh b㶘ʧ7#��@����y�L��B� -I �P��j�
�y"��&7d�M�c&E 98�ha���y�HH
q����m60��hI��y�܍pD��fʉ�}��aZ  ��y���/��B�k֟C�@@0�'���yBoY�ಘ���J�m:�������y�ꎍ��U���$_N��3,�:�y����&/�Z�J+�j��4G[
�yү�u��82��T�_��Ҵ䁘�y���{HHAT�WT��ZD���yr�wJa�ʕݦ�)4j̉�y�*��4�w��!�VUJ�H��y��������&&~��!SC�y���$-Kul��3W��h�hߣ�yBf������s^��s����y���f�D�Qu"ȣ\�2Hj��\��yR&I=l���9��9J�5�3E���yb���v=���7�����yr��1������m�&iI�Jӏ�y
� H�yD�Z)�@�
�A R"E"OfA�1�۸b6��*C���j�.�H�"O�!gE,|)��܀���*�"O�E�֍K��A�EE�{�& 1�"Ol�ƅТk""��#V�:ȣ"O��"�׉X��u!��U�%k�Qʠ"O����GW�QO��t
�?M�|�"O�L��,5�u�@�,�T�K"O~�B���(�*�1d�J5U�v��"O��R5�H/qz���" O����#"O6�Z���o���CeP�Jlٱ"O�٨'�M"=��)Y�	K0
���"O,@�sN�5m���V�=��<�b"OP�T�6i�j9�예}�N%ʃ"O��ks,&E%0�!+݂p��ź�"O�բWh<�� +�x���c"O���a"@�s�l]��G�H(��"OZ:6�Z8[b�pRH�����E"Odm��F�%w0S�G]�PxN�T"OĹh��:2��4��X�S�4���"O~��d�ܢV��Qrr��,����F"O��IB��G���T*n�����"O��+�	]6OR�ݘ�<4'���3"Oh=;�G�0r�4�s��?%�$:"O���VN3G-(��<�lA1T"O�4ط��"��C�N�Lt��"Oa���ʋ%�e��fʠ@�.P��"O�ya  �B12����X�r�p"Ob�ɗ��M8V0�s��U�H ht"OP�1���XmZ�YRZ��"O<��௉+7J��&��� JUp�"O(�鄥��v���z�3@4��"O�%�1O2���#��(1���"O2�R�`z��wd�H��;V"O��C�=�b���؆,ͬ�I'"O���c�F�F%�daE1жa��"O Q����N��,K[	��0��"O�M5���q(��áhP";���""O���ݣ;,�����34F�0��"O�@#NOI�tT�6E<�{"O�x�6������ / �2s"O�id��1���R�C%
"��t"O��1q��n����c[�%6���"O��hsB�_(H��Ad�	���"O*![�E2r�(h3!�3�f��"Oz�IQd_�[��T�!�%NC� �7"O��aG���Y�bU�o��#�0ܳR"O�гDV�q� ��@��J���"O�H!C�	5���ZЎ��!	l���"O��KdӇ�|��n̈́i��=c�"O��j���0��uA���,�D1%"O���G@�0+�3)��C�"O~�Q�#A�&��hV:#�L��3�>D���6
]�c����/T��j�0D��H��,3<�1hS(��	N��.D��p$͂�AZ���s��l��J2D�;��͂N�D;0M@�l~�r�.D��xV��8�ҭ_;0}"@jC�+D���g�H9~�L�a!�	�2  X3k-D���6OK�$C҄�K����B!D��
�BՒCӎ��������>D��B�)A��`Q��K]�H��Z�� D���t��L)������Mn5�#D�� �#'��X0S`[�15,E�m4D�� ���eL�e֬��L�s���"O��[�gQ�h�ƨ��FG |��"O:� �d]�}}x��q�ڂy_
���"Oa8u�ƹS���5��/nE�E��"O{��^��0�҇J�c3�e"�"O(IzG��(�����+�� ����"ON ���(0����a�(�H9g"ODi�ՠ�|Ј!xu
��o��9;U"O��agVN i��ʇiJ ��"O����K�v��a{7�?(���`"Ot�� �.���ٴ� #q"O@��Si*�Fa�!�U;��E"O�q�B���*|-���ɏU��i�D"O�A�b+�="�q$Q�{7���"Ol�J#F��
'�� T��(��b�"O��Y5�ҟ?�$�#��k�81B�"O^��s,��E윊E@I�w(�"O�$���')��TAi٨�(�"Oȁ��&�+%�����$��9f`7D�C ���jx����d:1^8 a�:D��j��ɟb���(ԁ�^x8�b5�3D���s#G�xx�8V�ǒY �a��,D���EI�S���Z�녺9V�	�0�)D���g�7y(����
 Ut��$(D�` ��`\
�p	�{#fź�j2D����ƄN�*�#c��1M*H!z�G1D��[���:-z�#3RT����-D��wS=7�څX� N�BM���,D���@@M"MU�i�7���Nz"���*D��񋝻�tŒe�ɐ,Ӱ�9w�&D����L	(~�1Å!�[��̘��1D�b����f�xzW醽4�*��Pc3D��#�ٸpi&���Ŕ:�i��,5D�liԋ�%<�݁�AM/�ɚ�`3D����f�"����fO��8�jɒ�	,D�LS1�T�#���"��lС,+D�ĉAv�&EP��ޫt��b�(D���_�4rdȺwk]ek�Ғ�"D��p � k��� �ᚿ��A�!D���!��'{6l؁�J�7\d]��e+D���%A�\�b|[piH��~�e�4D��ضo66����í�R��u���2D���m�=D��n�H�,����3D�i���ATnE){Z�z2A,D��a�̝�
��3��� )\")R�7D�0��jݹ5��C��x�M#�4D��p��H�L��	/�.k�6l�b3D����Ʋg�����S�nHh��,D� �5Cي6l�@�F�_V�A�,D�(�AL�&fv�فo��S�q%�$D�x���1K%H|���B=8�����0D����O�:qA�#ƼR&�0�G#D�`�� K�J:��� _ QD�:��=D�8�v�E'x���8���&N �"SB D�PA��4,�\I���*㴐��=D�8x��8J��4�Ɛ�N��%��:D�Ĺ���5��A����2��$n6D������Cú�g,��}A��c&� D�H�d�� e~<�
E&�GR�kv�=D� �+��

0��'�e��@���7D�t����T����!b(J�#p"7D� �dZe|ƽ2���<g��q�5D��8��D0A��MM�SݼU8@�?D�8�3�ֿ\~� {�^�`�I�Gk>D�� ��7S.]�QMہ4��8�"O^��� 3~AD�$� -�����"O����B�2,T`��)��L�"Oy9�h�!��I��a ��h�"O�J��� s�{�bC?&#�4RB"O����D,afb�pV��?x�(L��"O � ��]�r,jՠ�?-�9�C"O����(t�.y(�)��#�9�"O�p�bK?'A�0
P���e' �["O���D��!�D\�!�RZ��i�"O�M0`
@�
���TDď\���a"O<����/_|����9I� ip�"OnH�.h�܃"aG�~�v���"O�9R	�#���ɵ�L T��4�6"O��8%�Şu�ZP�aoW.�>m�D*O��:��ĉ`��s7%�^����
�'�����u{��8GQ��f�:�'H��{`	ƟZ��킃J�g9"I�
�'�H ��<F<���F�/1R�z�'�����ֶ[�f�2�N)�F�c
�'&h�+Q�0���D�P�҉ �'e(�a�V�Frޅ�3bX��a��'�z@�we��1LlLZ���"\ͪ�p�'�~����r��z�@X8M��=:�'C�ip�)� ��Jȓ0����'/���O�>@'��Wl�T��	�'���%��.܄2�OL"�ʥC	�'q�p�!,�k,ЦD�8�b���z�6���͗0-�D�po�69F�9�ȓ<��d��,�9���H� B���0����DY�g�@Y�i�%$ ��ȓyPy�ǡ��j�u86"�/)l�Q��<C�U�%��)O֐h��A�G�(D�ȓ)�p�1��]�@�5�55�8��?�d驡�0Rdb�E�m�a�ȓ'�4���mO7�`�c�mB��X���g���@3�6��v��/����ȓ���!�B4q��m9QN�/H�2ŇȓA/x,�r+پD����g��lȆ�%pj����WD�Ȧ�0a:�ȓI��9夏��½c�K'V᐀�ȓP����D�=*�.ثŖ&\��Q��>��݉�?E_�Ћ�'TU�L��#��xB��A-&�J������D���pl��� ÖZݼ��ȓ{��,Idl��$F�S�hQ�A[B�	��W�  mn��X�
�r�B�	�l��pZ��]��r�)S�lFTC�I�/��4ru�A-y=�QvgQ*�B䉌|�T���$O��Єk!/.XB䉒]�Hkv懶{ܔ��T�:+�B�	�I�R�C��D�*|cq�	N�B�	H��d8`n�7:����F�V��C�I�V� %�`oĴ��ئm�^B�	�n�fu�c�M/5Ex��V�ZB䉑5�NɁ�$Ҽw�Ҕ"dN���B䉉Q)�!I���$ˊ)q�'˴�<B��)B}���a�L�2�A���]QB䉍^� i �޳���
�-H��C�	*n8�ypf!�4oGv��Wf��"B䉩dh��S�I��<ƚ�����Q��C�	92e��h�,ɐ��̛��G�i��C�8.J��.�xa���`�Ħy�C�ɯ�p�C���=U�D+ǋ�#+��C�)� �p��6���C�+h�B"O>���㟚c��2�BJ�IP�"O�j���%5ӈ�z��]"���P2"Oz���5]
�pB��ڪ��9[G"O�e��.�J)�q��jE+Vm�f"OH$�E#Уt�N�;�CFz-fT`�"Ot���E�w����G�I2(��"O2����ҥ}6�����'0^��0"O̜sǈ��v�tQ�Z�g�d�P"O�x	�K����1�!PA���"O�1��j߱p&���/XR�s�"O@!�A�ǎ(0���S`X�ۢ"O�yj�ѝP��ٺ�+��L���w"O�%�")Sz�-���A�tE"��!"O�`�1�*��q��%,S�x��"O�Ͳ$)�,/�Z h⏛�5N�	��"O��Q%�_�F���!�N�`��"O��K�Œ����OU6�xѩ"O��i��T�h���;���"O�JĬ�%V{�,��n\�!�~Xs"Odu	�-�)1�,�@��D%$a"O$QI���F*�K(|�"�"O�]���!���K�"ۆ;}���"O$DbҦF7i=��#�3s��(s"O:�Ѫ�6Vx��Yp��U�|�"Ol5�J�`%�[� ։���c"O.z�S��3�Q� �n�A""Oz�G�ށ}Wִy�M��o����"O��H&�V�U(iC"GݬbuREB�"O��"i�"I�e��+� <�%r5"O�l#KYM�U+��;)5S�"O��@��,+��J�O V��v"O���KR���ib��~����"Oʠ`��e�b �iS�!�9�"O���Hnh4�1)K�J�J�"Ot�x��B�>�4X� �GS�,��*O�0�A�3_� ��ݎg�-�'v�4(��&fnhy[JK�����'AxBF��*C@�  +RQ1Z���'�P���&�YiB<B�޾��!�'��i�'�J73�"�I���r�8�'?D�Fܤ#�:��&���e@�'�<z�aQ#�8��(�6'��	�'
N �l�2H�i*@�V�8���'`P��B��'�\�7[[i���'�p�����5�P�2"�	W�%0
�'r��y�K	�@+�D�
S~�q�	�'P(Jg��?2m�s�	�tuH���'��ma�`׽@r����̃0C�J�P�'��踅W�y�Y+�-ӳ60��X�'��%[�̓4A��x���936H�'��1y'È�px�QE�3�f��'�p1���&J2nĈ�G�>��P�'��S6�N )���S���>9�ndh�'��0+�/T�|����t��0���
�'��a�IE�#?:� 9t9B�'�&��;9xr���)���$�'�X��A��fd%��b\;v�Tq �'��lq��A�FT�P��U8X����'� �� �T�J�P)�sIb���z�<����"L0��J|z"K�u�<�Vm,`�;��Gjk�:t%�p�<)e�&��}�CL��BK�p�<�P�A�j��t@ÉȜP?�(��ER�<� &�c3関a`���e� }[�"O�)��!O�.�
��R#���:E"OMS��I�;�H�PV*A,�����"O�����F�E�V�pɎ#`h!"O0�W���F��<*�g� ���"OZ1�4���\��s�,p2�h9�"O4��Z�v�� a��*-x%��"O,�����	���v㗹wDB��p"O���I0"{�:T���L��8�5"O��ڶ	�={4&iش��<)v�P�"O`|� 䑻!T!�k�=ij���"O�y��*�4�R��֩
<rW��"O�]��j�� �6��C�4lU���"O���qÎ�U�T4�si �~ݙ�"O�쫡h�9?��3��ۦ��؉�"O��p�H�}��􈀍� 'Z����"Ol���U	�f��v����	�"O8t�ƣ�P$��cj�C�m��"O�jl��aꜝ�JT,I~<
&"O�Aq �
(=��ad�]�2��Y�"O�9��.� l�ޔ�T�ߘD��8ڑ"OԘ��
W�X���V���Z��Ԙ�"OQ��,	+����o % �"O���eQ�`�.�9��P�	���"O��0(Q�a��i�bA�cײ�1�"O��"	_1~�p�u��)�Ρ@�"O�� ���Rzҭ�#!Op�4�h�"O��u�ְ��Y"���lL��"O���v`�G�f�aV�At�dd�"O�=�F�^�X���^�a��u�#"O� �С�>��t����|&8x9#"O�%G��{��1�vc��Q�j��"O�,@����72�h;Clq�Dʵ"O��p��т�asV��6t�5�%"O" �V� ��29�҈�!�~z�"O-��O�E�}���ߓȳ�!�"O��
��H6I��#ʑs���;S"O�|��(�Ɋ���8?��̐ "OL�F��"�FLʤ0�`�R�"O���%I�O�6�@f".`z��"O�	�҆Zah)k��M�*6��4"O�����v�4չÃɣ&6����"O;��Y��|�!���YF���b"O���C��!Z%j1�q�5F3�9@"Ohsƚ5h[����S�wL�Kr"O��v�um
 f��@!@A�f"O*�C -.
ƽ��M�7}�m�F"O�uxamԒ[.u�e*U1�,��"O�x8ף�����p�:�"�k�"O8@B)�98�!�ѕM�6չ�"O������Xi�dG E��m�t"OB�����P^��3�S7�ތ۷"O��"wA��a腟]���pP"OH�p�,;dZ�' 	qe�X��� D�T��A�+t��R�Ƹ_E����->D����ƛ P������#�	�2h:D��Bd��>~t��Ƭ�7�b���6D�H{L��^�,���%�; `���5D�`��d^)x^�c���C�-0D�8#�*�p�t����1��lA��!D�8�tN��h�z�
�!ӁS=���g� D�@U���0�Z��F�]4yo\\Ʈ!D�ҁ�^�r����f%��q56��N4D�p��H�.<I*7A֙n��B��7D�� �M�φ56Rl1uj��&~(�T"OV��@mM�zܭ� \�2�T4�Q"O��q���#O�082�o��1\L0"O4�����H�!ŮҾ!��7"Ob�p� ����zD��)`h0�"O�8���)|t��(�@C��	��"Oz�X���" �4:��P�hg"O��y���&W"�;PE
�k���"OPXy&�N=����aJ�[�,�t"OZ�Jt�߿a"l�Xs�M�q:`{T"OԂ��^Yp4����64\:]��"O�H{��[�Tu���b�:.���"O��S�їm��-Ʌŗ*j-ʙ�"O���*N�W���B	�M(J<�f"Ot�Y��6!�T�� 8�T42�"O��2�E�>FB`{a�Φn�L��1"O|�)��X%�m�Oλ'� Th�"OJT��D�%`��Uz�.[;/T����"OH58a�߹��1�B�Y�|���`�"O�0�֊ �~~TMS�L%p0Zi��"O�-���Ƥ�'�� >�=��"O>`
���S� ���D_c!"Oj�U��=�q� %��W��Pc"O�pPW���;Q���rdF�V���"O����R<7��u�:,�{"O�H�!��x��s���:#�"O�I
���3vM�����5 Z�"O ��֡ϏUf�b5��d$�q �"O]�6恻&1�,Xc��H����7"O��s�J̸b
�d2�
*w:9�d5O �=E�dm��oe�Mz�eV�	��u�
�y��H1sx��da¶"yr�1�g��ēJ
R���#~���ʁ�P*[�M��=��6O��D��XQP��@5 ;��jA��t��I!#�b�
 ���x�t3��D�g�D������"Ga�`���sp, �F^iBU�1D�p��^�jݤ���j��n�N}���5D� ��x3P�Ą�8q��=5c�g�<A��c��'�^�}U��1b�`�	p���O�ޙ��C_�cb��
I�<]Vt:
�'g�M�Ë��;�D5З��2d���O$����>Itd"b�L�%�&��0E7f��DΨL�r`B�3#Ē��(��WO
B�)*���DLՖOMN��BO�����?�U�t�s	����SP:�� � 8)C��%���wˀ#`��$�E{����?�ZXc��ɇ/m�� �yr�
�d� 1	�ʋ�&�y`#_��Mb�	K�'��Ab&#��*TH}jd��E��8�	�'zP0�0*ҐŝBZ~�i�'��	��#�'"�x��C�@Wh��
�'ĥ"u��#P+�@8lC�>8��	��h��ɍ��c��C#y-|!:`oO�+{JB䉯dy�dA�E�,᷊QC�Fb��D{��惲7�����?r������0�yb#<(�@��&�Y1eH�!��>�y�-Og�HX�W�	Ǥ��@�	�y�-N�n���*vID#�xY�P��y����Or�=�;kX��D�G�5�������� ������7`T%�8(��qF�ȅȓ2D�)V��#��QA��8�Ex�)�2K׮iʰ֌�jW�P�	\�<ٵ�v���a΄�1��}����@؟���o^���]�'�j�(�(��t0�ه�S�? L}����0�`�%ԁk� ����l�Iw�S�O�$�����p?HpA�,G\��+�'�B�@���6iBJ"%@!v#XMx�'�x�V���O�LmbK�j�L�0ۓsB�O깡�]#I�D���L&*��Y�i����	k��hWE_:f�$ͺ4KJ��!�$W�d��ж(m�bhj���!���&���B$��١��@j�'���gh���f(P1,�:n�P���'�|�HK'8���k1�	�bfzŀ�O��=E�(
4-�y�&悔󀡘5�d�'���(ʧ*hCB.W�_s���s��F���s�"O��Z"FU�CN�4���\(���ȥ�'��'J:!�R�!,0�H�̧u�8ċ�'O�Q��B[<wn΅J���$n�Bl���hO��+�B^D����F�_�0�"OzJ�Q�h�|�&�ǻgyX�*�"OhqbQ�7d^�\˃�ΰ~QI;�	7N[Q?��ت*a.(�sn��g8�Yْ�<����ӻn�N�.���b���E~��ۗ�"D�4��%�L���dM�/�]�!D�T�7ӑ
>�!lȋpH��G�+D�d�w���L��I���G�9��h�dE=D��ӥ�A  $�J��8�BP;�L:D�8U�V�/9^\��*_��(DR��<�Ih���'3�=�a��� A�A��8,ED�o��<Y��T?#<�N-��Xr��%�a���t�<1ߞ?��@����X ���l؟to��ix�D��NQ��ؒyYH"F7���D}��%?`3G�6�s��;S�><��3D�L�%�=^\��7	�5eT�C�0D�����m�A AP�f["���e!D��BZ��L�4�R�}��D�3!=D��7��M߂�7���Wd��P6�9D��*q��.7$h�U�A�~O%��A6D�(�$ A #����	�*`$]��+�|��V���O
��s��']�ыN�U�d��"O�u����+ms��M�~����"Ovi�&ER$jG��R�
�f���"O�I;Fқb��xiB�L,� uB��i�ў"~n�{/ʥ)��ߪA���ғ^�"K�C�	�
	2M�*<荈�mA3O�C�I�b�>틐j�3A �"���cz8#>��RT>iQrd�Yr#���A�+$\O�b�(��쓀 �Z���Ӱ8�RI.D�б&*Sx�2�1����J����J��~��9O�)u�%mU��*R��@��,�q�O��Ic��HO����n����g��2�n���I��<Yу�m̬ �_V�n�"NH�<YУ�@����PX�Mfv�B֦F����PK�q�RH�cb�D�I�Xn�y��IS�_yh1��.~0E:�BܿTd�>����䃖)!�ѰQGC�Fm��ꤏ/��'����Ow�S+]���@��	�j-���A��W~BC�	��f��EP
S!���n�7QyC�	2 �>��ٳS� �
@j���3�D�]�`a�����h�rL^�zq�O���&.d!�eg��N�(�8§�4h!���US�V�J�T�<�	�D��Oa!��)KM �	���l�"q�#5]!�ĝ�K}�8P�cU�+�&Hx�k��ND!�dƔM���WƔ>7'^$��ʚ�#�jC��hO���&� =�baʛ"�N(t�T'v�zB�"̚��cZ g�r���N��C�)� H��.�!_����d�!�NIz�"O��A��L-+�.���A-*	 ���"O��X�I �&�pt/X���M�&#$�S�O���6v�N����65y�*��=�C�I�m9ll�գŇ*���!��ܥSm&B�I�a:�Y�!�Z>C;�U�p�:�B�I	~D�]�Fn9j��Aa'#�7[}���hO�>�ш��6�@CiW�lfH�#�K)D��H!���l��D`s��BQp`T_�����d�vcT��G�@��+ԊL�a{b�5�	�*����!�E�d�Ԉ����O9��=aÓ�HX�UFRR(�9R�^���>��)�	����I�LTH�٦i��K�!�$.B���CR��a�R�(�l_�'UG{8O8�}� ʶ�P���o��X 4�t�p�<ABFuM�8@A܈f����W͒s�<)B�پY�勃dD)
�Q��XsH<��5q�Z0��KP�tD	ǃ�8Y�!��+��X�'�����v-�"�!��L����	��S~��!_1v��d�{r��\)����D�	��B��$[.��0B;m*�I�g�(���$.��t����	�nb,rWۋ�"E�ȓV���HWL�M�l�%� i��ȓ}l�4H�N�0D�ChBz hM���t�c��Mڞ��*��'�P���	Ȇ=�K�'$��uB��"��1�ȓ`Ȃ�`p���>X�"��[�^*�i��=���scN�a�nyB�#! G��ȓq�j]���
E�:f�~�q���zA;�BV�q�m��D��1���0i��ܬi� %� 05����ȓ&�@)7nч#�Z�i�l���U�ȓ	�t��1�]�7� ��ɘ#X�ņ�K%�M�<5��eq1��,�)��>����P��.w�G\'s5 ��~$�0�Q"�+^��@J�����ȓ,��-��Q4z���&7���ȓZ����H��j�d��kE��Ơ��0���i�n^/T��'�3e�B؄ȓ�H���A���[V��0%�����l��%Jw�A5i$-vJFV#xɄ�
Dٓt�#�@ۓ��6�	�ȓK,k�)N 2;�,#���lX�����B���#Ftܒ�i
�Pٴ8��t=x��-�<�bv��\&���f��=��%c'y�VGA��|��.}�IZvEPLc�5
�m�ʴ��%���"� -��G�f�����s�ହ��͞NF��9�!�.���#����:.r|���*Qu8��ȓ ��lcG�p��#6�?lZ���ȓ����@Yk��)5B2+��ЄȓM�s�B�2z��K�Y�.���ȓ*а%�@K�%_�e��\�2c���ȓn^��겉�O����C�� l�y�ȓ�BĹ��Q/B@Xr�딕_$�ȓ20̕������p�d�*�((�ȓ�q+�+�E|�Kg���4�H��/�D�ŊC��@H�dɮE�6чȓ>���߅8���4�Q'!����a5��C H�l�K�m��>�<1`��� !h�c��o> 8�-Wy̓C��8Hj�C�J��cd��9��OQ��p�i�+D@z���JA�\|�P��S�? �Y�C�tG�ҀBIT�(B�"Ot�#�H��J;�A�7'e
���"O��j���Z�݁f	R�1$�\:"Ol]Z��Q���T��(E��"O� �ħ�o�ƙ�f�#r�Ψq�"On��&�����H� �D�֤J�"O�V���;
T��7�!z��pa"O���'��"A�����<=��=Z�"O� ;G((7����/q�8��
�'tn�jT�Ĺ��	�F��`Q
�'����3 Bq:���U�3l�i�'B1���jF�hd�zVd
�'���Qf�ٖ�����wd���'
�%e	��	��@�chJ�~��@��'�B�;2�%<������I�tOHA:�'0��Ё@�3	�XYk#��'�I��'����ɴt���a˵gJ��'­��`�O�Ȫ�-\�	*�'�f,Vք?���w	M?$�2�
�'2d�B�@S`٠�歞�Y� c�/u0	�{���''�疤 ����rC�
����'"Q�Њu�̥1���;%j|���I�@7��r����$F81�" �	'~��u�l�a{�O�r��+�혌qb4��.����U �d��U��f���T�
�9la|�ǫ�`���䖡x�(���ؐڸ'P���%��,g?R�P6�ǟ��3%	�^Ā�Z�����m�7Qp���)#3�v�["O�!)$.K����R��*+yԤZ`kؓF�����4��veO�WnkȜ�Y�O���;J��Q���ԘV̰����B�e�ȓ�*���!a	�{�Ɵ�D&Uұi�R,b �8th�Q$�%�"�f�#d���<� B_?q�P�'FُOd]QJ�d����,G#���RHS��4j��ڡkUAR�F�y���'#Vx!ѡ�R8 e.$LO���d���i�O�-k"R���I�i%B�Zv���>�cV,O�t�����bT�d���1�Dc���I�Ƕ]zƘ�r�/�HB�I=p�d(��c�!̅��n�<���[?u�~�W#���5o�0���jZ�u�v���a�d�)�y7��t�S�cЇ]&n5PW��y��m��`9��
 m����gCr؊j
P���Ipf@�<S�E@�dF/n��LQEO�e�'4d��s�S/'�&�a�Ú�=�Ա1ӓY��(���Q��<�A�\�I�������p=�e��6Q5z��.ύU��pC݄f�lu��H���P�	;7��qѢ�R�d3�j� V�
T0b�z����]$�#�ޖ/�,�Sf#��3z���E�4������x�\�z3�@�t������������6����Q����,Ȱ#�iA�A�X�p ��5�(	Ġ;��Cy�tڀ`����/	ƨǹ6�IB ǿSvl��P�v58����(�(q)0gV�</F�Jyl��P�˼Ldt�iƠT�%�p\�g�	�����Gg�V�ލl�����A�{���`�L�(3C���fmT�t+~�3�(ga�h�LJ���=--b�|1��
�{�@�y��Fl��x�u@P!bg ��A��?W��^%r�F�x��+�Gh��Hʅ�1��vNHɑ��޲!Cr}+��!J�㟔(�/�?6�ce�aJ�̪��R
E��;cN�*u�9��C_��PKmqf�A���;k.̉p��.���͈�<���̗L�d]��C�9���3X:q����
/�#��Á8v�IseR']�f ��b��6!.8(�����(�pF����,�&�Ex��`f�� ��<�B��Pˎ��3@#$gt�1�፣j���t���?`�f�0���ȞK�'��EM���'F�R1�É��y��7���x�,]'5ޜ��Ѐ���Nh�)ەA�Z���� ���J���A�};:�c�6��oȉ�����/ǧy�a�q��ql��`Ъ��?�lHZ0��d�㞈����#BB�@�e�3|�|0�	T	x�r��p[�5��K��!�N���@E� ŝ0y�p �I��y��Y4Gėp(*�Y�I�72,����F{PPaWS� �zl;��'����1Ҍ���J	)�Fu9���#���P��_@���R�G0�h	�4ؘ=�5D
*�PMy4������7�ه�؀��ڌ;GZ�����Z�8�����r�iB��'Y+��ˢL�;��چ��b��b&)γ8k���CI�o�:-8�)ˠf��8�۴6!�-ݧ�>m9�쒝cx�D1��n��:�%����E*FH�W���'6,5��$7��-�0_K�x�Qӟ��a�hl��Ѫ�ěB� �[��K|����G�	�yr*R;vk����x�|��fĚF�.�{��$X�YBXC!m��1o�|{�/��K�A�1e7�B�)��7�25�D��^LDsq�2h�h{�O��N�EC
�����f^-Dn�X��Δ�*�0�����j��b��uX��X�GzR$(B[>Rђ��G.�mB��$'�v(��3�ȟx����fd *OpD@_F��Ƅ�<�y"�է9#�
��O�|�R(G��lm
����0<��@S�F3,�ôҲKr�|)����@��/
V4�%f/4	�T��H/���X��^i0�b�i���5����D��'��� �4����y�%���G��ȣT��Rf�8c�h�����z�&�{>�{�藛}�<h1��F�U�ȑ\�i�x�!p@ԪQC��!e���1O��%��HO�����\��Mx �1������z�h����H�;=����+�Y��QP0�1����s>�.�@��I$S;��4�'2@(0��O,�h�/�}�(����ǑO��cY�|�ɢW/?�r0��>?�AI�g�x�0ْc�FM������|��nZ<
$aÁ�	;��x�D�L���$�vJ���-G+,�q"��^
���!а%�T,P*��pi �O_� 	{"KD �yH@Vǂ�s��dŅJ2���#�E�E�t)��H �]�e���j`ːd� ���I�;|*�h��ٮ�)H��	�v$�DH/GRu`��A)c��iI��]0H�Z��0���b����U��qO�ӑD?g\v8�����=�7�H1L�;f%��$A;��{��(�1��cTx$�a�S���9�g:���t�]x��豌ά#�x DX�,Гg�dw`A�'��ԛAއT�����l��#a6��4�̽*�qX���/�N�""�H�ē��V��ܱ2��&i"��4������qAve@���$/,ɻ��A(y�x�A��c����T�ϰ�Z�Y'+�:/E>�c!o�'�lA2����9J���һ�|m��)�%P��R`��:.A47��L����2R��bĐf��agm��	��9R �e
�'��1J`�^aP$	fH�p�&���O��P��x���d���VME�o�d�EG�* :��36��n�@`Q��5Zq��'B�-ʆ�e�x�u�~�m���$� =�����q��ȅ2��P�� _�\���S%^�-�Hx��O� ����N�:\�]��Έ��ˣ��A�Jk*�R2C�'<��8�I3B��dh��3��">��g�:�����2�l�3E۽��I�SJБz���)W3R�ͳ���<��G�N��~�Y�Ś=��u��j�'|�0+^�]}Z��#�	�8�VAC�Os�'̎���U~�0ҏ0Pڄ̉S�/.x))0g�
b~��&�UZ|�ɒ�V�vޠ0���hQB��g��*`y����c|��F�_w����67�X�(eͷ	~�5�5㐸i��	�5�*�V�֎G�Q�wM�!;Zs�_���D��`01�оR���k3m������M����?1��6m�8x����"�#y��ѫ��ڙ*���i��\���jJ��2t�U!*_�\ɶ)�6�z���(@N9�rE����o��iC��Z��!*\�d�F��=A4���1�K�^����WD�:f"��;4<Y����]}OD�K":���ڑ́�#�P� �@5	��a"�9;n�Cb��|���%t��c�� �T9���6�$���;?a�­���Z6%��,�(����' ����`�<��P0K�/�@�y#W���DBxx�A�N4�(e�ⓟh���E���(%$%.�*MZ�^Ԡ0�ϟ�M����=�@�/S$pd�P�n�i���d�Je��g9艰Dh�>�d�1k�����'F$$�p�G�J���p��f��KR�! O��'���1��_cr�d��0������y�ņ��GH�I��"��s� 	���!}�J�JSiܺ�mh���#���g�D.6�օ��n�E��ϒ�_d0�c�#"�$��Hٻ%Y�97����4&֘y���"�@u(��0a�*Edh����$��E��!���]�J�	�@�`�E;�a��*�p��ըE�$�̫qF�WNВ��\�P�a����o�aku�/�b��6'�:B��V
:"�С{3��jv���?R��t:��s��qMb�W&�%���AwɌbf]�T�-�w`>Q���I���k�N���̌uD�{��ht}��Ԟ�W E�R��o[� pA[udP	p�(l�q%��D��-�a�4TD�8Ǐ�$_� �$|UCe�?���wC\�a��F'%���w��$)&�Y��ę�npB��w�Ep�ҝ6j^�I��% ���@稐��$��yepvM;+���x�%Y5tϺp����`ߦ��Bk�6\�M{�L�x ihFm�:(��� S�X�r��L�@�%X�4ZQʽ0��d0�c�G�L��N����K3� ?�F�/,���*���U��b	V:��C��E���]���Q�2MY�$-M�'�L�PЉ�_�-���L��$CrO����M��i�6Ey�\cŘ�y*_�-G4b�h@"CՌл�b��U" �M2R�Jb���_���#�y[�O�Ll��҇�l��)�`y� �ۑDZ�N�Pԙf[��@�w��?@���Mo��9�P?�X�u���G�HR��1�­	���hW��9ti�$]�9���� N�V�B�Z1;���|���j]���1P�L����[� �� �U!�+v5z����-��^���W��J��G��0��(��Q�:1�^
�,IqOƜe0�����d(�>�|$͈8�Hh�Cه%!���#�3Uښ,ppC��-}H���~a=�fd�.���s�C\)f�H���F��jL���@��=:���7�u+�-��_�����Ε1j�� ţ3̰dB�e��/�Qʷ�P?�=��J�!P�=��
�y�"%pu#�0��P2���(�}��҃U=�UZ󅃚s�sdռo��p��%���!��U��'
�y}:��!L�
ڤi2���\s�h�'GR�.\����0$i� w��9���j0�ĉ;%@(3R�	p�J��(�/_F��3��3%j�4)(�����B@����(c囔_��@p$E�I��5[�e��hKA�D�!���dP�� 3E�^���I�F�9I�e�1P�Eᅉ�fs�}1�c�% �x��GZ[�f`HV <|lZ�.�.x���)bz�QQB#�'����&�sD�p&9)��P$�0�0@j�9F(��{wG�u"��B� �sTBʸuq8Iˑ��0�*@�@+�4نE :�B9��a��x���l\���I� �P�+����ƟN�]�0C]2�D��n�4+����D2���2/؎|%`\Y��Y�> Np8#k[�+�����F`т���@�7���r��x/vh6X99��*���AKgE�{�2Lq}2NZ�q/���c��#eI��;� 麑[7��>y
�>T��rt$�	D�����mj�=��[-FG��0�O�3n��\��F^�e����	�C��5�6�L�oi�5�!۬E���3 �.�� QK�%PIH�U���x6��jI�pZ��ԉW���#p�R�-��1+A&ULD� 5�ʽ�&a��؉{�4���	#ݤpt�ZU����Gp���ɁF�"e���~� � W���a"_��Uc�F�B�y��'Â,�e�]�V<Ua�-�r�6�XB�H�\��	0��PB�T�)'� ͜���6�� �c^n�d1�߳@)7m��Dx�󳭘 .���s.ON�!�N�d�<�v�X����6��O��2��/XnӶL:E������ޫCfպ�&A�j���Ct�LI���r�DW�Xk,�VZ:F��Јd̚a6N��d��O[
1��[�ɵ:��42V��(�p#��G�<q�C)
#bY\$�K42�x�jp(�(c���� �'��q;�M,���
�R\H"��7R�R�j`��a��o��S"nlذ*�rF˕�T�ˀ�f��$�d�P�T2YTR�p�"olܤb-Wp@㵵i�	�MZ�? ��@AL����b��v�����	���� ��<���J'eG���dY����M�qaDa�0�l�ia2'˂M�t�Y����� ��
&|���-vnTU����o�uYB�OЌq�'X�&�n٨sj��@���`�ط{s��{��6�ɰ~J���սz���[�A�j��$"S�%<`�����\8*I��.H�3��l��F �LLӕ�Ҥy�8j�$?a萧��4^<,A��N�0�Ҩ�t)ŕ@��p�e��;z8a3'�(?�vkԄs"�D��.M�:��h�o�J]`�Og���]�aGb�+��M���=[��Ҫ!�ڑ�=f@�R���E�&�*���`Bl�{6D ��c��R��5vة]�P�vȂ�u�f�b�K;4�R���JT�m�"�j'�ƭ��#�$��[(8LI��]�U�\�:����&�`��TaGXp4�0�����]h�솯M|P�U��-��Y�$�j� `��B!~l�!���"^�q3Α�2[�<�w�^�g����ߘ4�u;s��}j�9)�@]� X�y[w��di�(^�ys���N�`�:=J�mD89���玻t�}8&,S#��'�i�ҡq�P�۳�E��1N&or��s�&Z�%{���&�#*e^d���?a���G��j���F�%h~��3 �+ w� �@��"+gT|�f��1G Ȥ��R�:nvٲ�%�#���Mq������(:V@�E�1�Vy�$g�/Z��^[�Xbp�F�����	H�$���^-)^<	X��Y79>��!������r�a2�]�s��O�<��H~�Q�4�ŁA#x�Ak�Yj��ѩM�*�H< T"��������� �J~��f� ���ӢI`.`#�I�-XV I
S��ɰ�f65�~�A1d�c��`Ŋ^�Mg"@ks��_�3����1~�DXt�@�q��,k�a�:{$����B8s�
�0"���G�x�Zha�� ��u׌��@o����.�Uйbf��#	\P9!I�9��9�a)b��0��}Rʘ�7�*di��ĥB ���G�$U�0�2�@�� t�5��Y�|�o�Aу�`�^K(T�e��$V�$�Bd н8X���B�[�x��ì9 ��ـ�  k��T;�L �5ғO�\+�,�*6�٢��5,�fH4��'s�����FM�^�i��Z�
$�(c7h	ld�YQ��7����p�I�q������N�1si=.��;P���C�^?v@r����#vD�E���;"��3��֘l@. J�ADo���mXq��& ��av�՚����B�ǰR� p�e�g�@��
,+?f {u�_�IH��T�(O�d{w��F���p�ȃoonM#�F�6�?i�.�lB/mn���v������K�!ő���]�3}��{��.0̳w�Y�EJͲ3�N�(T ����=yT�aG��9m�H,;V�`A��t��ՠW�P%m��*DG���-7��|^q��fL�F|�h��P�q����E$n���'���rÇ#_���D�&8�PB�鉒6�Ri�!cP�gLV�kr��S��׿c�t�Y�J��d)�x;�֝4�v����V���CF��57$t�a��?�z�l��s��9�돛�y��$[��iƅ�%	�ʩ�a#��M�T :ǮD����;q:f�0���G��xd"����H��c���=�7 �-\bliP/K%+<|H��2�͢�eF���PF}�ʗ��82����t�q�E�(�zM�ɣ2�Fh��4_�J�JЪ�5� �τ�q�M���Ī�zE��+
�-�P[�Żs���*F ������1 d>ث��TKsx]2��
�4A�3>���g�4"㬽�aJ�v��9�@��NztA;Zw*>��I�'p�u��/x�(H+c %ړ��a�`	�2AU����G>�	L"	z��Cco	>�����4� ~(s��,Uk��$�:��'���6`>Y���E��2�� s0DPs&�+=Z��S�O�0���� ���z��Gk����@q�	��~kY��N) ���'��"<)�/Ox�R��|�<脜?#<�3��I�&�Ҭċ@����o�U����G��6xb�b�F�.`�<*Q��qE'g(!�(��ugB�}�t�'��:#Sџ���V	��
q�1Iծzt�D� _>n�Q"O�����!R�q��Οa&4!z�"O�,֗�P�)VlV+�Pۥ"O̰���$�H<2 �ǜP����e"OT`�� r�Y���H8� �"O�hbC���6�R#ru�"O�qB�EU>|}�=�4M�y���1�"Ol�� ͆"d�n���j�F�8��c"O�cퟁ.tn�
���Q�"O�hqb���evfdp�HN�.h�t�4"O�t��
O�>}`tLsJ�Z�"O �Tm��\��	C�C5�Hp(�"O �S3 ա.I���˨:n(�T"Oex`��.$��EqCʚ2Lo�-x "Ot�� �&DÐ\���u86��"O��0Q�H�~�a��K:`Iۗ"OD1�Q�O�^V��G$W�l�����"O�0`IL���	K �M�����"Oz �ӣ0�=s� ��S{�}rT"O�IKO�\)Go>Uaج*�"O`����4�"��o�oBճV"O ��f�Y�-�I:g�40��"Ox��P�<jݹ���L8� 2d"O�Lڄc�#".��p��!�2�b"O� �U`��Q4����Ce�y��"O�E���z6U��nK��%P"O�=�����/JP!d�ף~p�aIg"O�ԣ��Z�c�f��,΃g���B"O�I"�舃X��ܒh��{vd��T"Ol�
��p���\:Wh��H�"O�A���ҾvJ���c���M��qPB"OJs��=\%(��E��-F� ���"O�ى�j��'ڕ	�|z�DiE"OTy�5��v���qm�.�Ĺ�4"O6�ӓ#�0)�8�p�m�>D�1"O&8��	)U���¶L��F$�:�"OL(Q"��Y��������?�lCc"O@�3�'ٺ.\*0�*0H�"O�-���w�,x��O-�h�d"O�5�={����D�\����V"O�C����4`��]�YKZ��y�	\
=c�i ��õ(.d=��@ة�y2J�5���Ʌr3��C���y2�A�eB�(�`M�i�|���մ�y�&K�C����gbܑ��l(r�ȫ�y��ؕiofT�e`���}�����y�HȦ> �㯜> ������y�dR�p�}
򇜪Xdxy�'�{H$1� g�'������FO1r����b��Bț�p#>}��'b� H��w�I�&��;'%&���$�
5hg`]4hP8��d�>��q1�1 /��3��REa{��=z#\Ly*08}�}����2c�Hl�g����A�����d"S�K�a|RL݁a� ��! (��`�EN0۸'q4��r�X,a��5�EΟ<�%gS-q��:���l�8fK;5��K�jݕaR�E�"O�q��׶d0 ��P/�,3�H���6j�`Mv��>	��v�ܩ`@�˖mѮlȉO�&�λLz�C�DD�btC���0fFͅȓT���"X�dy�2�M�7L>�c�ɐ)M.�):��� �t��#�0T� ��٣as��<�C��mA���YX�ZU�	������b�|��UdSI	T���I���b�@�/�j�ҕ��6l"Հ�"�d�2M._8��֑^V�x�Y��"p��b^�%91O&|��b�
 4r)��E_E"�}y���'�c��\T*Mc)��<�$�#���-yՂ24�2�`��~ީ1W�F�8x�)��%�"ܴc!���p h�����|Wz9j1@��{ح�O�u��w���6�ce�8!)�B��}�<�������t���J�!6�ϭ ��Q(��O��]�
c���
�`؛��������T�~i!�ΟSiZ)xaF�4�VX��)5��x�o!����ț%�@hZ�A��M2�DB��?���QB��$`�ĳ�I�W���Sq�[$�Zp�'F���n����C�D�|3V�`�y�1~4F�0�D�y�<)X�n�GP-���cN��w���
`sTN<} ,�e��\�������F�����g_ހrI�*�D��-(2��<H��*#�t0�R���M٨�bcI�aTʤ2b��)�T�ܴRa6�I��w���GR�"�t���H'J��e2�'3���b�ۙo0f��G0I�B}*�Cʫ/������<{���tt�jtT�0�n���֖a�b��$jRR�ШA�5��(pp�Ч8���+��'��D��r`	�Cu��!�\�P�~|��O# ��͓D$��r��%��R��q���q$��/��'+`Ł���\��hr$�=DJ"����]P̒#+�9��DY�~��p�ea��>�v9�$�Q_p�@&��^ZT08��Bp`@U%�e���Q� Q����?�f�� $%��(�'��캅��aT�X2�ըEߤ��/�\i.$!6H%"LN�dm�%NrT9#�^&����Kt �y2H�,] ����v%�H��]�2��I`��eB�;4d_�Y�9{��N�		�8DA�Ml��gm���0���AhI<�(杕O�ۅ*� ^:x�@�b�:�Ov�0�n��)q"T��I��a�ZMH|�VE��Dg��x�^5s�,��IX+-��Q	f\�V�]K'�@0O����r��em�� � �7w��=�G(�3I|:L��d@Z��Ոf��z�~�d�B�|G
Ա����j�<��Hy4l�G��\����F�2{�x,se#/)�D�b�Ǥ�tIx�ɃU1��
A�'(jP�07,Ofȑ�+@z���]H_ZM��J�z�dী�<O�������79�p��k |	���TN\�JYXa�c�K�y�
`��F�D�`�
eD�!C�[/�0<�&�� �J�Eȉd�b%i��#S�����B5��E1�D\lhpu�ߍ3y(8Pcn�PLI��i���a�hΩ�R� �-����@�w"�A(���?7j�o�wh${�Ol�2T�8<��dRV��=)(�㰧�?�a��R1U'�UY�8	���;:btȱ�#�o�(8	s=Oҹ�Sf��?�&3��IG�:9frb�(�F+��"�̼�p)�5鄑��Nʑi�f yM)�\���-�8�&�G!�ƨ� Ɂ�邽�b���p� ��"p��5)$\qE D�N���B4�H* R�iもUD ��i��RVp(<�.L!fЪ4!�+W=piH"�" ��(�-I��j�cW�v'B �L�}�+V<t7mM��<eA��	`�X��ָs�ax�IK�7�Z,��>B�ȉk�&�R��jJ<Q���Þ�È�8�	ΩG����aEAh7�U�pLΦ�9�(4?�w!�`;���t%��bK9W�Z�q�(�$l�s����Ch�oD� �"T�%�Xhͧ<���� !\͊�	JY�r�$*���0�6<����@�4�I�<����P��o��y�� 1$*���k��6��X�&���8F[��R�	�("3
�j�M�#@�'z,������3���:t�M+�N�����/�$EC!�$�8r�ӓf˼t��sG 澁��#K�:e��{�j��~���[^=�,�#�
�q��[@�@�⸉��c��M���	93��EqW,��b�
E�ׁ#Oʑ�&Ί9fs<K�Ț�(�C�D¤Ԛ	��,J�jd0�"hM�z�&T���M˲<0p�G�+��x�'��՞ٌ�$L3d� (�A�G�Z^t���mЎw1����JA�ڢ�l�Ql3&�Ha�ˮ��-�QNGc��u�B�X�|@�6l�%�j] C�Y5*b� �,��i�4c�(�l5i�qO|I�P.��6P�		�����)W%�,�)@)R�!���P@ꈪ{�ri��nS��82	Z�����9�͑��5����&(A��<!��W��AnG�@
�lx��'3��c`T�W��Uj��V�ʔQ"I�= D�k*X%f��y���c-���s�T:U��u"l�S�ޤI�Iۦ���lO6�^�A7�͕��1C��+>��x�G]�6TjX��D�#+���3��JhEiT� ,"4�	�㏟>�&8 ėE�D�R���C<�ԡ�O�Nb7M�_��Ν;�> h��݅�.��pKD�_Ș@�'(M ��'ɚH�g���uH�-�T�ѵ�	�}��H�N���}��� ��aRWj�#0@><��n�5/"J����%t��5�'�U�BBԚ��}zg*�~��A����n��5RL 
�F��p#� ^�j�pM1󥅢i���1(	�@����V�1XT4r0����hd�Ƙ�BI�3S���6\�3�Y(u"z���!96��)Ca;bo�4���:���V��oOtC/P��|����k.�Q���P1<�Z5k�;��!��b�kFj%r�cC/V��T��X?g(��n	w:�3F�O4��[�A ړ�,�3#���9ug�*�QP@�\�~SP��scN�.N iP��)Wԭ����83����DK6�j�G;y_F��Î�/HYЄ�Rs�Gg�/�p`�	ϞUk�D�����$J;֭d3�	��ˀp(�2�dH�T'�b��AS�MHې�O�G
j�+�-/8��TA4
��6�H�Cjh��eE$2�0���/�I4{�T{���[�8$���.�`1'6q4��UlC�]���M�?��A��e
��g i���c��(f9v+�_P��h'��O����PAd�<���I�s�Ve���I'}F@U�Є��_I��`䇔/��)�Q�{G~��5D��Jjh�2 �cK
�හ�^K����D�/��Q��Љ}Lj�����sb��ҥ˦&�-�b�ֻ-6p1��dH�3�T��U���h���ܔ=���g,ҘF4�|����Q�:�x�f�8x�4���O����8ՉB�cf���ǌs�~����ߓ�u�a�5���;^cC ��pjP�BLα�P�� ����O�J���d��(�%��TuH�a��	����5�ؐV3����-��u������J�Y�	y��:Y�&�S7�l������P<���U��=��d%䨙��>!���Q'�Y�7�y�1nZ8S˲�r		qH�Aӝ?}�W$?�(��ڢI5΍ө�
/z�hQ�"��)��S�H��2�r'K�P&���.��'��#=A4l̘N~@�SpbI�uGBIHr�سæ�@qLE:,�@�$�� p�!+`l��J�S`"�sLXqH�G0ʲ��,ĸ$����.Us�4���Tu�����,ثi둞HK�
I�Z�H����8U���fLյt]&�h@O¾2p�x�L��5E% �>�{c�6d�,��j� WU4�8�o�<1x�p�O��! ��wX���O%sR6��\�L�����?!�� ,�^H���;~T��� �rS��)s��n���I;P@��S@>H�b��O��DS��۴<�R�d/�!��NO6�mk��R�VI.P��O�M�W�ƌ"�t���D�@��j��X�{t�X�N?=D��hQ*el�E�g�#�p��Ã)E��V�|j�Wo�<v�@���Q%-DX�$�֯x�f�3�MU<�I��@�J�I7TN��bt)�~�5/ޭ4j�8�a��i�t��rd<o$�}c�H��4%���.B���6B�52g�8��)��l�|���D>k-�e�� 
\���'��VJZ��G�? @���EIy�KVO��08p��2&��I ��j�d����#!��JT�Ү�>>Z	�C�wɪ��,�H�س#U ;�>1!� ���ZH������靁F�d��.��%@�؊�NG�K!ک���,)�rA��i0�� i�8R�R����-I�28ͧ!�H�{�o��߁�A���l�#����0� $�dFR�*�10�V���q9�i �Nn0��B���z�{!��WyB�x���G��3C����)W�16�ȍ{�k�T�Rt�I?mָ1B�ϕK����g��@S��������*��1Nn�z ��+��0�
<�lY�D���	Qmd�� �!8b8o�TR ��>A��M	3J�z�y��� R��JL�oҘ �$��b#29PUo��(uц��M�h�F��W��aѲm�8֌����!AN�3�і����J0P$Q��^\��p��[h��e��Ä�#�������l
>)�j˽6�����B�-�|T�W���LN:+fU�b��]$0IJʾ7�򰛀�,�xX8a��H�J`Y"$�:��%g_? "ŉ$�F#��	�]w��#� �H�xaR�Y�%�8�)�?&��I'�):�-ڽW�
�WjV7w�8��"ˏfӼ�S%K� �|E+�*�X+��(��Z�S�8��*5s������@��Ou�!��dxV�h"(5�(Ԉ�瘰*��i-dJ�(bH�4�0䨴'�0+��u)fg$���8i©n7��T�� }�A���� �v��6Û�K�z8'�&H�V��O�QҶÐ
=�,m�'�DP�@a�A���	|%���_'�H�p�����8���@�yH��T�F$sP*��dˀ&�D�8��ӳ��8�p��;Q��`#�.D�����8Ai��'Xp1�h��U��-
`�)|N��!�V!i���1�`���Î7�䁁@�V�(@�/�4�x˟�*r+` � 'k\��a��0�����bw�90��6&~�`��:M��x��������M�Z����݂d�E��*Y�&p��ؐ/T�L���P�D!�C��~��I:���i�~%B3�U�n�t0��9��ب��V�2n^i��!ˇ�?���i�x5jc'l�ʓ>3��ҴD�>O>E�"��=.�� a���LK٨��&/b��*���	�OL�Уd��.b��ڴ$�d�) 	H���u����Xg��`'����4N5���a̐~�
<��ĸ<т�F,4I�%S `�g��aՏO�? V�26�ИJ����î�"<����a2���O�==�\)�
/F�Z�㑚N������"9������-d9�i���\�H��(2�-̍L�}����I4�[�����==F��a�@,����!ɳ��	�3@xH���;�,�+� `��<�'�0H�C�˓= �6Vo�@F[H�h
��
�(u+�\�g��;v8v�Y!,��W�z�
0`@�qؑgc�����O��S�ieRk�cԬ}&�xQ�� r���CY �&��W��Tx�9	*Ob� 
I��<�g"�L�j����13/R�7i
�(ɄG�H��5S�T�z�
-� �BK�l���I27"H��P	�&�Ԩ "8�h�h�[�eI�'�r  @B�h��yI�-5,<�Pw�J�'C�� �@ADh�˱��|rl�q�蝷S��X��޲�����GD��}�!��o�	��
H2|wf�Y�H�6Q��@�&�0EH8�@I�$�|�Y�C#�D���O���H�K��j�b<	���_2�r qq�?qqBk;Ho�HJ�+Χn}��B���&�֩�DF��C��D�&�/(�}ar]�Kg�P��P�V�I.+�ט-tO��Ño��~]�9��h5B�,p
�9�Чe޲;��IĬ$��'fq=˖(X�O� ����J��{&	I�aᗨď��TC���<$d�$��X�|�D�ȡ
O�I��S�{�Ǜ'�|�[��EO���7lM�Ho�$����:c�Fx�D�A�}�� �ĆH�N�r�[�/��I���Lmݹ)�����qD�U�\�D"m�a.T��2�ҝCNN̓
% ��c�țU�
���	IFbT-e �yd�U�'��e�Ҧ!>�y��"O�L�q��4*a�yXb���2K�Z��+e�u@RC ����&K�� 9w�1��4g		�����;����/B=s$��"ǡ���Q�!��r#���LI&�V��-j����F�4�s���a��X8UJ!q&
�8�k9FaJ�.�U��1�15�����/ǔt��Ḯ+���gͽ-}�X���%?��`��A�Ut�O��T���{�Sj�#LD�+��ڽkofꄚ2��	���Ep���6W34�V�Qӊ"HP�K�{RN�$F���⤀C$��:&"�it�8(I�4��-Vm� ��G� ��2$AE+��2e�� �x¤P*F���d��9>J
@0@�H��Ae�
K�2��#D���O� 	 ��[s*aHP���C'2��J)	G�Lk��_U�ĉ�ǣ	%y���� d����9 �O�*{0�l��ʛ+I�d#�^�P�֩җ�I�y����݋f�L��D�]� �\	��Ik�	�!�Zĉ��"7Ε0�oE�I��	 r�5�4$�����J��0bMj@%�SI|@��H�S�N-�7�%UHHe� ���RUH�z;xy�e��y
V�I�8�
a� �e��S�k�A�d��N�/��� ;v�BP
��d.������ē#l�c�.�t���&� b��R�*l� )V|�nP ҡ�&|�3U������D4{Gx���K�$Vp�����'N�U���V(l�2a*�G����0�7��7}Gd���kr�ř��F <½*��ݍR�f\ڕ�0A�̅��*{��e,�e�'��
�N u�^�nO=q
v!�v&��d�4r��A3,���;@��ik$1V��"����t x9�&��0f�<z�O��P�shS�OA��Ԍ��zF�I�p)ғjK��y)�$'wJ$*6�=���*?�z�����7M-*asS��2kz��SM�K�q��S�3���A�j�fh�'���yel��8�N�����cF�Y�{pR�uKɊ<1��P?xļ����(4�`=A�'&�S�$/��0bǣ]��E�f���w��a�󆊌~{����\%j」PW)\'>j�����Y�̣>94�K�qR�h�

���ց�A ���M�� �,h�(B�v^�p������v��	B �L�S!�2PaRx� g�. �R}�a��<a|���Q�(��0.��*P�R�!SH9�a�GV�&M颡�*e*Xu �"�x�i�.R.^��;���!3�Jk|ry��ꍏA �$"�퉢g�����X��bÓ��A�&U�vų'DI
)� ��=���,=�JBaD�z�ax��\-PP�T2��E7dZ��K��?	%�M�A}2�i�V 4Y��)�'j����?`b��(wʦa���y�
�t<RC�ɬ��Ue�&v����Ǝ�5
�ɖ'�܁Z�N[�,�$xϟQ�t����4Yc$	��<\.�A�'�pX���,�f�����?9j���	Z;u�t�.�z<)��6�싴YMK�ps4�p�'�ؔ{��~�'U�T�5�ԒP��!����	��ȓmH�a5�C�>�@����(<��ͅȓ/�y��i�*$rB�9�׼}ybԅȓfV��G� �q�D�C��ńȓ%2�@�#���)�:9�JE��btC�JP4��T�^0��e��8�9@F͗��L���W�*@|�ȓYT L�ӭI�8��*v���P��=�ȓ}�0ԣq� �����9�ȓ{R���� aʈ!WZ̠�ȓeL��z�
B`�6���S�ḣȓEn��T�xL��aa�^�d\��ȓ�����n�K�|�!�L#�*|��<�52�ň�4���4n�#C����ȓ�Ѳ!�tI��� �3�'�~4�kCK�K���<z���'7��gH�S��Ը!cr���2�'���X��Ӈ!�8ī@�j� �S�'Wt�FC7�Az��l�JT
�'��3g���O���e !�fYb
���  �KF��<�P�I��T���"O�I��6hYt�@"��dk��BA"O����JM�G��X� ��\W�m��"O�)��۳bzDP�M�1a�N��D"O� ���8�|1kp�O3
�H�ju"O�ܐ��l5��򬌿v�(�g�DM<y�ڗ��>NfԹ�C�*/�1O��I0Y��b��R�I�n�CQ��LPT��H�dc��
B̈�4.8ҧD��5�#Ȓ2�U2�h��`��uAT��;�(!���#���W>q��؀a����$�K���a nK7)�	֊�<MC�px��ښ�����~"Ü�"�����ڑh���O��R1�= J� 3v�߼���[�w��!��f�%��#��;�ēt4H�f$�)�S-KG|q�w鞤HB�}"��RF��K�&A��;�)ҧa�"}��#0���N�@ߖ�o$]4i���<tjx�NA?"�ibİ@Crh�S��w�!8a�������n�Ќa�*�:-,m��Bp��FL�T ԭD�4 '( �0�t�(X��x���Ͱ^���MC?)��5tl��rȟ��U�ɒ&D�F�[R�K]�ȵ�fL7<�.mn��zJ�t���]9V}ֈ����'|�PB�5���I#r6���0��nk҉5�_��?)wC+}�O��<a���B\�T�DB�]�h!4.J�;�.@ɕi���	Rv�#|��4Q�.׻R��G�K2��ô��N�p�#�y�/|�v��;�*"|��
�w�YP����ebV�3r��n��7ebT�;�}�g�^t%�D	1]N�j�E�|j˓<%Q��G��Ġ�6]q������`��M�5�S�Oo��0��A�Lڤd0h^�R��1���I3�0|� �܅�}��Z9�*�X���`y�ID�j�~ĢC%�)�C���ҁ)��Z�=5���R��6m��Y;0!9F��3��)�}� 4f��2&�\��C�_r��w`G�)kJ��	çj8����.I��GY����	���I���',�>e�D�zج����5!�Zsr�@����7��S�'H�w��zdi�V�ͯc��Q��'!�p�jDD����Ջ��[?��Z�'@qУ��|��ٵ�����'&
᫶,
4�C��q�]Y�'-6a�F�-c�y��*�R����'3z�R�
W,l����C!K�'�r���n���(��0�]�
JZ�`�' ��4E���ؖ��*F�3�'��Y�T��j>Y��ůwҨ��
�'"�ڕ��T\�i7\�4L
�'�ڜ" �S�� @&j�'',ZH��'Î���P ����*���@	�'��\)�n��Ign,�.��%N���'ň=��ŚM!��k��o&Z���'�Fрꔠ��׀��d񎝫�'��K��I�n�A���	H�2@�'�r]rD�E�*ĺ&��G��I��'��Иw�V�7�L��𧝿1�.��'"�P#d�2]��1x���/&5��J�'� 5k�!��+�68
�N۱M��r	�'���J�4R���K�#M�) ��'��Uss���lU딁��Җ-��'�*]d���4�Ԥ�3��vq��'h�}q��ıe��ĳS(�6�\�	�'��dp����_�,��7��	;�8�'�������F�=��OU�n�0��'N\�!��Íuh��6-�?m����'�N�Q-��8�)�u��-n�Q3�'UX\#���@�&�
��fE�u��'?I�En[9<� �4��)^��H3�'K��c�k��� �(3l�0���'� �`u,¢@�R�ȳ_]����
�'��a��7��8���J7�8�	�'���SP�t��;F,�H'�=�	�'ݬ ð)۪D}�a�PN�:��<���� ^���X�L����e��-e�p("O�	���b�u����|���"O��k�°]z��+��	�njti�"O��r�\�nh�C í4�y��"Or�S7a�4M�D �R@�x+�"OX���ۥ=�f����=g�<�y�"O��iF*G8\�;'�Z����$"OX���ْ���+CF�cƦlA"O�����l\�!5Ɠ(?��}�Q"O 1z�aJ<qH�}�	��D(#"O*)y�GS��E��GӅ\�$�h�"O���P�v�d��lG-w�tA u"O����K��^�J��fk�-�8�W"OX)���Kp�|����ǣ@���K$"OB��e�J� � �)�-�@�Y�"O,�`�BM���A21�_"Bvb��"O����=$$�-8Gj\�(Ѱ�`1"O�}�uؼKr��g��%y%̽�"ObU����2�\Q�����Lx�T�B"OV��'��x���+a�<~Zf1�"O�X�n̡���Ac��Qa� "O<`F��BrZ�h�C@:l_6�"O��(' �M�-�P(=9�X��"O:�
��
a�� z�gN�p�"O4����G�����cQ�-�l8H�"OR	��o֑m�0���A�@����U"OZz�eT� \�KFF0.Lc�"OP��@�`��A��6&�X�c"O�za(�:1��`��8i�g"O$��F́�u"���-��!�7"O�<Q�Yϲ��փ����y�<9�w؀Pj��D�e���Y���K�<)1��\�BA˓�]ߜq� DM�<���,@�0X@E�'X49)@(LJ�<yǚ�zF�٪�!�O��XX��L�<Q7�	��с�=L<�����_�<y6Ď��|�����$��(��X�<A�DK3<��	r�A_tA!�m�U�<Qq4��P��	ۑ)c�و1��T�<��Þ�y���� `J@>.=�k�N�<�fB�2��\r���FFU��%�A�<�1e@�@�f-��OP�7L4]Ϛ~�<�Dۗ"����UB݂|n�i�p�TS�<���_���0�o���D�g�Ez�<�RkŻ�܈����]tL�k�ß_�<�Ղ�	�.UQ�lC�0�����BY�<�wCՙV�H}�-E�;b qCV,_�<aU�:��P��
<k�����c�<�R"��0�Ȉ��J���Pe3$K�]�<�mB�(o���G��m�����R�<q`��*_��|B�L�fJZ��"GKM�<9�DRE~}�6��;����C~�<�GT"'��"'��{-�UQ�<�3	Y�QO�'��4!�����K�<i���5ZA�$�-(g�(�7�һs!�DX.Oj��@kB�@T�HA�#q!�Y�A@���an���*����̡E�!�dƆc�p+��8h��0p��)&�!�D�	2 �tÇ��f�0��G3G�!�DՀ]�Z��&�<"kjP�w��*=8!��!F&DHÁ��kCL �D"�.WK!�d�y^9p��:]��y� ���w4!���>*�tB悭n]��Q�`���!�$���Y�B�hkF@�!V0~!�� ��`6�ȍ�.E:��]�2k�! �"O�Y#Í�#1(DpB�Q�p�T�JU"O����.m#�ɀH�N��4�W"O�E W *uX�B��A�`?l�B�"OZl���Y�*�t�䥂>G3(�t"O"�fc�-� �)��W90���)"O����o��O���� ���ARf9�"O�h�4N��Y��9(7����"O^�R�C2^C�!S7ǔS��ȑa"O�����D�c)dd��낷f�B��"Ott�5��9}��I�s�Q�p���1"Oz�J��
'����ӝ���c$"O���r*�3Ip𘹀�=jK
u8"O6�#S���®	#2��� N�<.�!���l]p8�� 2R��1T�]8f�!�d�-��4s%�n�Di��!na!�ŕ*�P}��a��a���I?ME!�DB�C��R(A�!��&F+!�$���xA)��ȴA
�C��ԛQ!�B=d���b�sY�)���F�6!�D�I�.���톻QB�%�@!�!��;C�l��ż1�D�u�%�!�Ē&L���� 	��iw��Q`OF�C!��,0�����`s � �a!�|�p�j�� 6��PKs!���_�@���L�?H@��gaM#!��]5��0� �g2��8#�Ҵ(�!���.7X�h" ��4)�e���`�!��B�DQ�뎽r$�2���n�!�C>R��%�J�E �<��D��=�!�D.4��e+T�5�q�Q��&�!�$F��H�j�N�;
��P�
�!��N�9:y�7�@�X�H���,\!��>,3ܴ�54����,!!�>%#T�!cc�,�6<K��!��41�"�����82���2�>?2!�D�O�l<��ǀ9�Fa�P�B�l�!��;�� �����/�0@��IÖk!��ʥ��@-he��!�!�$׈1��	��[/Q.V����1�!��[����oBA�򏂡�!�Ċ�?�p��BՅt���g��d�!�%}n�mR��0N��<�Pa�!��b#�����A�@���!�d������)O�YSc�95S!�$PT��
��!D��5$K��!�$ԧJ���8��\@ !���=u�!�P<9h	��K�=^�ք��
E'9!�DM&3�頀�NQ��"�f�W1!�dP9jx��`�
Ym$=q�e��z!�dD�o ����SF���DS�*�!�$��k`eC�גk�RÄ�U:M�!���m�D���1k�T�*��,�!�$
������Y�7f6Ȱ1�U+�!�D��|꜀��<lT�!� ��!��z�Xi�vl�2[QJBR�M�A�!�͜H��9ₗ�y�xV�>x!�ĕ( U*�qEͅlU~!��	�`%!�M�{���Ǝ�-u���fI&Y6!�DG�~�H��5�E;T�i�G/�046!�D՗!*&P҄��9 �����혻I(!��R�I�ej�Ŏ�p�68�w��K	!��ǱDVt��R�� (�!9�!�W�v����P�	�>i(4e/!�� ���ԏ��L&���S�)J&"O���B�S��}�e��,����"O���-��%c`4� b������"O0%��G�*�t9��`�8*D\��"O�EHFO�<�J)# Altړ"O�M1x�F�z@a'fs�-��*O�A3��I+����'��8?�>�q�'��TRE"�V*��c*i�1!�'�(���B9�1���[�	�'HH����j���땫c���z�'�����&j�
���T�	�'[^�b�#vZ]
����Kז��'r�ɹU+�>eW@�t�&=3���	�'���w�N&�YK�OF=g�T��'�ʄc1��Q������1	�R}
�'3�bA�D� ���
�,�1[����':$:����k�Aݲ�i�' ,��J:*�:��L�'��q��b���Tm\�����'|L���ʼ=Z�A�Q�0�R�'�։�U���:4��½��'@���(�;o%re"�h�y ��'}�(�!
7?4)BSƗ}I�x`�'4�x+��Tca[R� �ua���'�,���"�^�xa�Ӡuh���	�'��Mp��O(8���� ϋ�qTF�r�'i��^4@���0h5w�x�0�'q^(#ևő,� ��T��s;�`�	�'�~��E���QCǣO���E�	�'�p!r2���|�PQHv%����9�'[��+��G����⅍R� �ZD��'[��{�JH�z���E��%��]��'�b����$a�r�*FO�<����'T��#�-P8^~M��S�Vd:
�'r~ ��)n�T����D�@uJ�'O
�R  ��   '   Ĵ���	��ZI�2;���C���NNT�D��e�2Tx��ƕ	#��4"�V���D?W�m�'CT`�,�	
zd��)́G�B�J�d���jz���Mc �
^	��	c=9P���*pi���0��k�e�6xa\��b�?$ ��*�?~m0dc�U�����Whʸ�H��IƋ�3k4��i��G	D���1 k����V�i��I�W�lI�c�MV��[Hd�A��ޑ�'y&K��k��m"qN�,A�U�%��b>ެ��'{D�	�hh��qo�n�ӭ�D�'�+cR��uML�B=�iP���'�Ep������Q����w?��bW�[_H,"��ʦ&X����җa?���@��4�H>y��S�h&��с�7��ػC�!2�|��
�+NY�(�1�|�DK'��0sqL�x~�J8~DXP�Ʃh^}�e-ĨG�]PW��/�ēF>�=�q.Q}�Q������Z|}��t=2��:آupш���?1���	"	��%��ゅ̀%�.�%���abE����e�H�k�
�3`���$�tL�hߌ���9y_��ٰ�1�X��L��!!�5�2������0�B������/��<�W͒ O)�ء��O�		�l(&uC�ҟ{�&g��J4���IQ�sp؉�v�@�\r��;��=	��Ɍ�yGln
����$N��"���	���N�(\Q��<W(�SP)�J�I.8*KP	���8�'��|�f�D?�@�����Q����z�N�a}2K8���0L>���Q�8���$�����Rk>��EaG7pQN�����=V��5�|2'"�(M>!'�L9�l� oP�'X��0c*�,B:&i��.�u¨8�e��1_N,����bm�� �?���Ib?q�!}�@���[�w�xc1 �A�:�s�Z�x��j	�|V4�O�����B�pN�'pj�e�F.n��a8�h5:��hi�қU�|�"N>�G-��M�F��<iؽEo�����@�Ȳ�a�A�5-�Q#�'Et�Y@ ����?f��w���WĠh�"O�91ի�+(�\�XQ@N"8��X�"OPm�Ŭǎmܒ�X���*S��]��"O4���C�:-aAKW ��*�"O� kK�4
�u��IʏU�*]3�"OV`�3a۲a?��a)0ɲ��S"OJ���6t��)��Ӵ I�I`�"O��(c��te�u���;`�����"O>�CE��H|Z��wb΂Zr<	�"OF�� ��r4R�   5  �  �  ,   O+  &7  nB  eM  �U  a  %m  is  �y  (�  j�  ��  �  3�  u�  ��  ��  >�  ��  ľ  �  K�  ��  $�  �  �  ��  �  ,
 � % �. 	6 K< �B SE  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��[J"<E�Ԥc��[w��;�ц��
t�!�đ;\��|�1a�- 0�a�(����	Y�}�mú��q�NT�l��@Ⱦ��=	p�@6I(��;�'�:�0ɏ�z�*�S6A'F� 4��'�
�Baj��״�y��@��`�"6OZ�D���P�^����\�P2TTk3d��y�)C&H��IJ��A�@Ь�5 ۩x�6l����s���!S�M�X���{��=) -=D�`�V��)G*����D-q���F9D��P�B΀pF��sp��=kc"yqr�6�O��';a�͇|��p��F%P�8=��'u)���<HI^9P���F[ �I���4�'Y���S�\*SC��ۥ�K6R����=Aۓ���dņ��^��W�T���p�ȓk1��� G�8�x5RV띙F��@��w�d��3�9I�	�w��K�����4��"<����'��dZ�_� �9sJK�)m����Z2"!�dI4����i��;f����=:�ɇ��&�JZyb�>�}�qk)u��3�`Ӏv'�<H�JBX�<�O� �AO��W�]��,�U2��|�>O�6--Oرj��M�$A��R�"������'KQ���~��������4|䵹����
Ӑ�S��'D�̃�g,�t8��вA U)'D�؈��l��Lp�K>}�l�נ1D� !b��!<���0�Ɓ�Xl�&�.D�����#<AX���n�59�V�k�N.D�����Ӛ8-p��<�P@���/D�����<Z�q���>N�JX�%�'D�x�G���zوpA�."JL���!D�����í#����RMy��>D���}_��rra�:`�<���7D���T��	cô1�fAԅ0�u����O���S�O혍�U�*@a6�kXA�⇌��y���j���VE��v�9���/�y�ѩ�~	P�ɛf�࡛��Ϥ�y��V13_�\��l߬)E���Q��yě�4:~�spfPV7,�*��eA6�=�;�hO�TYt(�8�N�s�K�12+J�qg,D��HŒw� ��Æ��$: ��(D���!Ty�ᦈڑS4�ce1D��	��-p�(i�v�:&V!�*D�P{E�=-�2�b׉
x��@	��(D��0�JФa�� ;�!R�0��MK�	$D�ԡ �NT��^��}��!$D�  �#�d�N��7��7s�es/ D�s���s�D�	2�L6VuDܙƌ(D��{����/��@w�O�p�rt� 9D�(30��q�@HSq�Ϣ&��)��)"D� 9��_�U�v��D�N��$(���>D�����&�0�{���`bHx��>D�x������#ËE>J�6�%I2D���ī:	�.X0�B�_d!�0�/D��3�a[
S�"p8Wo_�4��C)3D��c� KV���]t��`j��,D�H��l��f�rLB��m����)D�X�S��0X���'��|�lR��)D�H�S-L.��%��K�8�u�=?9�g�(XF�Ј��Ă6�ԇ���6�I1������^eR�h��2�
C�6���у���@C0K1�ʯ��=yç&� �A��׶Ehb1���7A�8���&T�E�� 
�~���I2�Fc�B�O?��m�|��A��BY�M�r��7m�qO�O��I
B;1O��`!$��z����C� #"
O�6m$SZb���N0/�
��2 Z�}䑞`��	=B4���g�+uy�u�ЀPKˬ��d.�	�����
�R����M�
���a%�@cQ�pE� �JQ.�����j��)�C?}객�-�/]�ʜnZI}��';�I�0�3b��y� �V��=ь��<1��4�'!c��(�/��Sn*��A�Yzt��A����A�8W��؂��ӌn q��IMyb Z����jH<Z�"�S�<����Cfɀ�	��Z5����e�'���d4�@`D��%>4M:Eg^(C�i�7)q�F����?*�|��K3D�@:��	6W��ۣɮc�2Li�K/D�����,�@�AN�*~g��6
 D�������u3���/V6uY��8D�x�q'�������M�i�^���9D��@2¢GZ8]9p
��L$�3�e,D��ӆ���-Z0�v�C�"��X���=D��;fa�*�"E�K�\4p���"ړ�0<� ��sMH>vv���#F�^�@ 4�"�S�'��d��F�f pqʛ�q�ȓ L|��nJ�^�hsI�8g��GxB�O���d�i�I��툤l/L`�تpj�B�L(D�8��E�[4��#q�Z�� �f3�Ir���Af��G՘S�MRd�$����s��yj�J*(�b5+�dN�݆ȓO�!��*DT��E�r�̼CԆēa���' ����HšQ��ʍyA"O�cs�5���-H	B��'�1OT�I�^�����AK�9lr�͍b��B�	�6|V��7�0!�bL��K�{���c�a~".�	&>���F�=5<������'�ў�Oڬ��`	�z[�@;@���7��E�'-,@Y�_�.c.5ӗ�A�2Ϭq���D+��I���-v��p�h�\_�,2�"O(�R��կ*	(���Icf�A��'r�O��1S4f�z����ȱ&j�$��"O��Cc��d+��!��SRZ��e_���<���ԟ�P�WN�!.�0IRm��*hr�D"O�Jb+R����{f�T(,L Tj�'Pў"~��K�AE*��.��U\�
�D[��'���쨟����͗%#^I`4���:D��[�����]ޥG�4k��T�S�T
�<a��DU�y"!��b�M����6�r�����=�x�'�$ �����dl�2Z�6�\��GH�X�'�џ�s��N�8J�� ��2\��� D�<8@+��c��U�U��%�hx� f���E{���0:h�e��0��-Xb(�C��|��)}Rg@|�h��GS�H�04��?��'аcF��)#��;��(��ea�r�'�Id�'ݠ8��FB \�����F��ȓ+F�L	 d�<u��&�1�x��>A۴1�\�>�@?�bn�!;���3G�e���AH���y�G���4��4gnʌpQG7�y"Ȉ�7�$��-&2xb�A�j��y�K��~���3�ɏ**wT�[�閁�y"�U]d|��6'��"�f�R�aڡ�y� ��\ *� w�վ!b&���,�y�߽}���,S�!H8b��P��ybD�*o���s�h���X�ca�Q�y���EY�q��N�S~e�Cϔ��yBNN�W
�P+T\d��7+��y��bײ �.�\p
��' �ydݟ~t��:�đa۶�jW�=�y�gY�Y�N�Zt��&G�`@G�	 �y��E�B$ܭ�����i�ƀ	0�y2.Q�]7��b���~+($K�$�y�,��#z�e"�A�zh�rĎ��y�Y�=�Z���bܲ$������y�H�@���b,H�+�c��ybkLȮ��a���� sq���y+A	�e�!Ȃ������y�m�>1Af�e��<Gj�<3�@L�y�+B�@6��i�C�v�Ҡ��y����A����g�*@���	��y�C@>p>��@�*
�tD���)�y�\���8S�Ϙs|�Th��yb���/��(*���@�ҕ�eᙨ�yH��6t֤�1����S�Ӌ�y�	�dorI�$�)0��!M��y�H�:Vox僆���"f ��y���r[��x�x� �k��޻�yR�ОLаX{W͏�sj���m���y
� �% QmH�=��;/2��	c "O���t�N�+;��B���T��r"OtE��<��)R� 3vh�Y�"OB���ء*H�fh�>)B|��"O&P�$�< shQ�9-`hX��'�'���'=��'\��'���'�,h�&�R%'/�\�@���s���c�'���'��'���'���'!��'�#��5�(��Fl45����'~r�'�������'���'���'[`�T�E�Y/�Zu�ɭ&dM�T�'#��'�2�'�2�'��'�2�'���2�G��Y�&=�W�
~����'z��'Jb�'���' ��'��'�h����Fv��1/̎,&�����'��'���'�B�'��'=��'��ˠdY��ۈgC�����?����?	��?����?����?Y��?1֤P�<�qc�.B��c��?����?���?����?���?y���?�ъZ�w8����B�\Ix*��)�?I���?!��?���?��?���?9�hT0u3<E`���yD��fP�?9���?!���?����?���?y��?QU��.U���{�$P��05v�
��?���?���?���?����?Y���?ٴ��&>��y'++���]�?��?i��?���?���?���?ic���O����+'�$H���Τ�?��?����?����?���x����'4""�UI���!�yn�� c��L����?�)O1��I��M3���57KH�t!f/�2]A0ٱ�d�t~" t�v��s�X@ڴ\N��@Dƥao�q�Ǝ-�x��s�i�����q�OP��i�69��9I?�* 	�iq$��#W�8�xG�(�Iݟ�'_�>y�$��XO��"�'W
BL�[�̚��Ms�y̓��O>�7=�B �H"/DQ�wI�-����Kܴ�y2_�b>��$� �	�R�I�F6e醈Ӆ)I<���Ta@6�ɜn(&��2��h1N1D{�OR�@�<�@db��l��D��y�[��'�pJ�4È�<	� ^�b���ˣ�ػ?�8*;��'C�����kk���I]}b�ʮW��i�#�fG@��FC]"��B�Gøp��OG;lv1�HX�"�ǺDv.��D�]J��9��M|��̯gL����O?�I�hv�ɢȼooX4�6��bݐ�ɤ�M�J~r�p�$���9G�桫UO��D#g�w|�	
�M"�i��� ��[�O\���免>F�!�5��*)�"ؚ���OP��A���S9��=�'��D(��8W�E�wg��Q_��F��*2/�ɪ�M�qC\��:H~�� ���j1)G�O&Sj�XW��9Y�I��Mc$�i��d+�	���d��}���	�e���Q"*X�&v9�S ����Q��\B1������Ք>����0Ca��%]*�ࠢ?|�ubL�x�'u�	s�I��M{��<���+�^���ħEh�!QdƓ�<�Ըi��O�9O��m���M#��E�a[����~Ѓ'�S�ol��Wf�"`>���nS*5x�fܸ1M��j��?q�S16K�m8ZcgR��cR�e��8W)�:z-��'=�[������0�y��X�"1"C�4�DD(��$OʦM���!?���ix"Q��Ӳ�D<iE6ܸg�#8��)�4���<��O��m���M�|X��a�^�<Q�hZV���iR�mcLh�g�
�R�nqvo�2��V��hO�<)�$�V�Q�.�=�Pe¥�[����̓����^ ���y�P>��A�.�Z���ϥ:�p�׋7?�gR���4W���:OH���	�i� H�c���E��6�2���S�z
@��2������t�"gO�hʰQ��7%�8��G΂�Y��	�* `��6�6b�T8;�N��z!AA��f_�1��̇�u�\i�2/*H�Y���(^���qC�	S�(AsE_�5�90��S"�̼ t�E%v�Y���Y�~�ǅ j)�0�#�[��0H����Wr�x�0&_\�n��d@��[�N!ɑk�W��al�X��h�����#T p�޸!�F��o����l�)/N,�Ŋ�.>*pz���.u�$c�B��9B�#�}`�B��ݧO&�!F��N�*	�`��R9rZ�tX��A3gԠI�5JԪX�d��&�K�+0p3q�x��'B�'�����\���O�E�֣ܚQ�h ��ۉd7�M�U�E�	ß���̟��'⮌з�v�kP3<���cE�8��:�&�XD������I����'��'�)�����{���8vb��bU�2e��K�Y���ҟ<�	ry���R�d���x�F����1�ؿ&���U �ͦ��	ß�'@��'�nU	����[>8�x i���v����	��M���?1(O�m`�,�\�ɟ��s�%(�$�$I(L;h
Mq|LS�hӜ��?���5�@F�4��M�3�@�=�fU���M�hPJ���I̦�'����`����O�r�O����c�%����BK�:�� l�����	�/��͖������'T^�LB8'��+C"����,��4wL��дi�2�'O��O��O�i��&#��8$C���*�#��lo�+O�:d�'�2�'B��y��'D��d��>��m���ч��]"��y���$�O���ϛA�0'��Sϟ��	�+���� �$�8��#�%>�Խs�O����OX���O����O���Gk�%A�(Q��*#��1�������>j���(K<ͧ�?����D��DO䥛QO[�U��QǏ3v'�o����A
+�	�|����'6�H��hH4UJ���(�PF�����sd�O����O����<!��?YA� p����k�"�QsDKP7<���t̓�?)��?�.OʤR�g��|�p(��e�>偒	�)x]�@�n}��'1�'I�I���I<�'h�@JW�U�u܆( ꎉ{}
$�'���'c�	֟Ĩ$��P���'] �jf��np�g.�&,9� qӎ��/���l�7YG��OZ�� ��%$���7&��`���w�iV�U� ��U:�l�O���'���@R)nhh��	2���@V [���c��I3h��XCVN*�~�-��d�@ ���@�E�@}2�'�x�P��'���'7��O)�iݕ�G�5S�}�p)O��d�>��n �U[��G�S�'O�(!⁈ݻ~�L�s���5�f�o��*+2���Ο�I�h��jy�O��Q3gh�X���-�=jEΒ�7�T6��%�v����̠�î5��a[vHÎC�}�0�K	�M+���?���Q~t1�)O�I�O�����8C�U!n��bO&8���wJ<Θ'y�Q���5���Of�İ�4�'/�"��G٠(�2r�>� ˼����O����O�b�$�$͉�1��M�
TB��Y� �#���i���?A����d�O���tJ�6L��1�3��
Y��0�f"�A���?y��?و�'�d$��
ܮ�⒣��d�xD�.��tTR���O���O���?F�������W�s�`Ј�AQ5@�T�Z��MC��?����'�rۀK"0�4�ح�r�.�P��W��<��'8��'��I��� �WJ�t�'�ָ	B�D�6�p*��&p�[�*pӪ��?�	����j]Qg>O�A�ԋO�t� �P�w�0�i�2\���It˂U�O��'��D�W��=9FN��|�(�U���b�|�	7`Qx��'�~��j��Tbz��,(�������a}��'B����'\��'8��O��i�	H�c	�l8paa�9	�j!��)�>Q����y��P�S�'	cTEY��FPn���LJ�
q̤nZ����?���?)����4����Pm�$x���0t	0e���%]��nځ( !�q�>�)�'�?���V.@���cN�'J���6�'�B�'�T4�Q���,�	C?!�$v�`0����1�j5$�O�m��K|���?q�'ʦ������e�'
��ss����4�?��5��d�ON���O0��!ю2l�8�0M�;���զ0��E�������IGy��'q8����>/DR�ÐGQ Cޔ����%��	ܟX�	����?��'f��C�\88���%ߚnJ(:�4\�ޅ�'D��'��I�ܫ5F�b��J0.(��Q�X-8����y��埘�	C����$қg��׹.����)F?�
�7bN����On�D�<1��u6n��/�8�\�/O����əXE���c;���nϟ|�?�)O\�ZE�x�$Ýhl����Ϣ&�z��%��M����D�O��3���|���?���3ђ�ұ��;s�@=f�d�� ID�$�<)FMD��uGl�7 I['I�!�
��DO���d�O:�`D��i���'��O��iݩ�4�	�@���a-�&RT�Q a�>	*OZUT�)�	#q�#��RC��O��YA�iQ��R��'Vb�'#��O>�i>��	3I=������)���[pO�Ri@��O>�:�)���x�G%�:BZd�E&0ҕy����M����$өA���|���?y�'�.M���Z�P����J� �i�� -�ɡCw��XI|z���?��'�N��q`ȮU��Y�fbN���i�4�?92�P���d�O����O���82��l�|�x�F�1M� ��sJ�>��L�Jp��'M��'����$em=X��$���.u�!BC({ET��'���'����O�� �M9VN5������%�f�L6� i����P�	̟��'�→�kg���9Q��'g �lR��7PY���'��':�O���O�2����i�Ԭ�[ q�7��8a�H�""A��d�OZ�D�<Q� ��Q/�����r�$�s���;6'&Y��`Q�~��yn�ܟ��?��Y��a��E}�	�M�" Y,6���Ä	��v�>��<I��T�:�`*�b���O���]��%���0J���0����b2�A�>a��[e�a'�k�S��G0��II�h�LL"k����D�O���wC�O.�$�O����F��?y�"��^��U�!숐w��C�T���I,g�d@��`#�)�Ӆ_�@ء3��{�ij�B �p6m�5e���O����O~���<ͧ�?��=YjҴ�Ԧ^�[��s����`��xm$)P�y��	�OҩI� P�F�ȦI��=��1Hd�Y���ʟ��	>�t�����'���O�J��ߙI��T�3�@#Ԃ�^̓1��P�#����'K�OX�[��.6%�*�GM@Z���i���3H�쟨�I���=a�)�-)bam
1ϼ��b~}��D�P,�u��Ol���O���?) �;���Ӭw�0��"��6Ͳ-()O���O��&�Iß�7L��y� �{eB�/:�����b�4�`P�/?i��?y+O|��
.�*��5W�&��FoR�A�<�C�;���'��'*�OB�E��K�i��y��N-��Uj��sw4PJ�O����Oʓ�?	�j�8���O6]!1��tI�f�$%4}�Wd¦���U��?If,m�i'�� �!+�Դj��z��)�2L	��i��X�H�	,9�O�r�'��T/\�b�p�%�7N��2�0 �c���	�uD���4f(�~�d-��a���H�(�a�����'l��r+y�:��O���OO��$��0E�
	f�eꚳY�no��ɿ|�T5�I럸�����S��h�i��A���"�(��R�Ip.��jr��p� �Цa�	ޟ��I�?�S��8��� c@,	�K|��T�46^dd!��M�2���?���?�b��|�K~*�'o�P%z$)��#ONr�dޯJ䜕0�i���'����9z��7��Or���OP�d�O���;w��� ��|2��Q�Y�Li���'�b���k�֥�S�4�O���'v�x�烸��Y�L�R]	 F�k���d� 7:ldlןD��ߟ������ɥ�pHRĆ�5�	�3�P��|z�A�>�� �A��?q��?����?�g�:����.lb�up��Zc`��f�i#��''r�'�l�����O��y�0t�)ǂJ+���t�	�X�Vx�'���'���'�rY>���	��M���9X=t���L&FLF���"E1p�f�'s��'ar�'��	����ep>����81:�-@'�"s�!����M���?Q��?����?���1囖�'�N).�lA#�G�
\m���7d�-&��7�O����Ox˓�?-K����o�$�LfJ≇Q�F=�����b����'d2�'�.;p6�OV���O8�	�m��)wA�'5�i��ǆ^tf)n���4�'7��C�j�Iqy��MQ�e8����Óh�D�$g�ɦy�	֟�x�σ5�M#���?���r���?#��%�dA�d�<$#f�ɶDW��I@�p.����	Hy�O��e�����t�b�Z�$��M�r�oZ Wv���4�?I���?��'�z���?��^�FL�G)8(�(�	bo¥988��r�i0t��'FW��ST�؟���5z��;��+a�( t��1�M���?9�j�\��q�i���'�R�'.Zw������J���k��_[��4�?�*O�#�;O�������ݟ��t���w�����BAv�9&�B1�MS�N��u�is2�'#��'��'�~�m��`T)�c[�.� #�]7�M���3U���?�������?	��?�����M[��ư>���hP��<��չ׹ij��'��'�:�'��$�O�y�%�P4TTpِԤ�Yʀm@Q� z�$�O~�$�O����|��>0v�i��� ��L�G,�M�b
K~�l�H�f{����O����O����<1�$[�u�'yg�y!Ӎ�x8R���b��^� �����������I ,ݑ۴�?���6��}���H��(� ��E�0������i��'��Y���	 �����@��t*:Ei� ������H�k�*	o�� �����	i�vԑڴ�?���?a��FQt�""�ϛ#H��O�B&FX1��iEB]���n����L�ɞl�R�s�`;􇎷$�e��js"d����i��	9.� 	�4	;��˟`�.���X`�,�@�� ��4j����כ�'5����z�"�|��/�!F�49U�N}%���B��M+n˞s����'���'y���4��O0���W�&&N՚���F��@�&�ŦI(�Km�H'�"|���0uA!f��@l�� � ���`��?Q��?��AN��'�'
��G�V�p$��t��| ̊�;��O�lB���O����OX���C��=y#�W�!���d�D�%�I�vr�N<a��?�J>��R��i��K�v�|����/����'W�쨌y�'s�'e�I*|�.���^� �h��oO6Ř�d�P��ē�?������?��d��e�3��p|) jN�MC��C�&�?1/O<�$�O���<9nӻNg� .I*�!͍���@�P�/E�Iɟ ��@�	ɟ$�ɽ �Ɍ$�A��&��ງD)��-j�O<�D�O��D�<9F��(�OxPqb�6 d�9^%�8 ��q����#��O����9$)��>}2(�{䴻NQ-i���ѤD��M����?�-O|8`T}�ޟ��{�ةZ�L��Ch�*v�	1�$A�K<����?��
[������Z&k�j�ْ �X=��@���v]� s�ȃ��M#!P?u�	�?9C�OvJse�8<�( Oӿ���ih��'5FHr��'Tɧ�O>�Q���?6I���+�
7J���4Z1��c�ia��'�Z��[�I���Q�)�09{zI8w+��	`!�M����?�J>E�$�'��йg����8Ib�	]v��	�p�`���O��DY&��&����$�`������!d\����mK �mZ^��>�)B��?��>�Ѝ�j�����%ߝ1��B�i���	z��O����O��Ok,�9:�������#@�t���W�t�I ���Ify2�'YR�'��	�%����E_�M���贉���D̢�ē�?�����?���3����GK -]�1�'(�'Z�M��P�<�*Of��O���<A�囀<r�ɔ8FH6��|i>L[s� �S����`��^���d���ImX���RqR@0�T�"l�@ �X�2�6��'���'��Q�d� ł���'Z�o���4�!(R��^��1�i�ғ|��'������y��>�d������Ȧ`��@�C`�m�	ן�'����)�)�O����J���� V?C;b�zcGɍ�ӛx�'K��K�NMB�|������e����6 �c$K�M�-O��j���ɦ�A��`����ܑ�'�-����<���S�@5���O��������O��~� �q	�+X�p��8�G��	N�:��i�T�QAcӒ��O
�����e$��%]1��s�j@5CF\���]� L�ٴ?��PH���D�L�O�́����Cf'��;�(Q�&yB6��O����OZ���e�O���|b���~��	�_��-�O\0�����`�dc�,����>��'�?y��?	�K��;�B�9Rv�����-0�V�'�,�
�. �4����O��'d|��`��c�X� ��:y����O��!��d�O����O����O��q֠Q��ia� �p��1cD��t>˓�?����?yL>���?A�A6]a&��'!��4�X�ӔBȯi�>+�A~��'���'�剋g\혟OQ����n�a�4`g⃊Ԁ=��O
��Ot�O�$�O��2Z�(�Q
�.j��R��a�b�2׍�>Q��?����ě%I:t'>�Fڻ<��6jփg���Lʳ�Ms����?y�A ���>9R�ԍE���3���(b8�@�@¦=�	����'�"��Є&���OH���M�����ș�.�>	�W���IL&X'�x�	џ�� �:�S�̇�=�5�'&�$��͐�+
��M���?���W=�?����d����K��v<�[�S9�kt�
����������+r�b�b?�I�$�0�$�UƏK�T�  .�O� �s r�8�d�O��D���I�'�哜x4�r.V4�&I
!�؈�ٴriHhj���O`�'k�ŊʖHz��9[�n*�*��|��7m�O�˓E�B��,O���?q�'j�k��e�.UzEU	�>l�PN)�Ib#d�iO|���?��^�� 	�J�.b�d�@�]�rI����Z���ß��I\y��'�'@^M9���@��a���Pp��>I�̛�r�^h�'r�'�^�Т7fɔ+�"���b�SR<���BTWz���J<����?�����'$B�՛.�����%Ʈm� I���'���'Y��'L"����i� H_bM��E�%!�D�Ӡ�֝|�F�'32�'
�'2"�'�F� a 	�M3��Z��)@�
4M�rd�s��]}2�'2�'$��i&*�N|vD\��t�P���Ė�`���6s���' �'l��'
 �}�B��r!H�K�B�4nY�(��B���M���?�.O�A�F�y�S8���r��dà�áI�^�'U\�3J<!���?1�HI�����
r@��Y*F��r5��lbش����`�.@n(����O����d~��K5�\�E���)����S�ܭ�M���?Y+Zy���O�P��>��zr+�K���޴j�����i���':�OE�Op���j���1��0��	��Á�q�^�nڸ/�#<E���'�|���9'��X`��%5mʸ��p����O
�$W�ed�&��	����p�2Ta�m��.�x�D��S�-�I�HS�b� �IğD�	�*�J��
	���!�(\�M۴�?�gn�J��'��'�ɧ5fo��9���6���pw
�p�	��Ė.�1Od���O���<1�愥J�8�@1-�&F+`�
��LKj3�x2�'�җ|"�'���-2QC�J�8]�P����""�l���yB�'���'���'�����' 2��#T���$*�C�<~��f�~�tʓ�?qK>q��?��â||m?X��O>�0��&�$���?y��?)�Ohhisg�~��*o�!�5:ΰ3��J�*|��7�i���'��O���/5�ɼ=e:&'ٵpA�q� ��G_�6��O~��O��D�j2~ʧ�?!��j1�F�~`��e��):)�@���Չ'R��'s���%��"ɘ���W�Tҹ�q�U�i
�zB�ۛ�R��H)պ�Mk�]?��I�? �O�<��ϒG���`��B�N�zg�i^r�'�B�+DX��S͟��3�ĉ$0��-�V &$�&�ڲ��$���9M`6M�O��D�O�	QA�i>-��8(�x��Whl����c�:�M3񁜶���O���1O&y�V������/��h/��
�OT=]a2��������兆��a{��ߖ7�a;E��;WX�I�E��p?� L}^�dږ)rq
�'�}ܕِl[�gM�����ZHz��DZ����5$�JE%�U�5iP�KHQ�� �Jf�:b��>d�
$c6F2
�&��a惧9��=�W-G;w@~���6z
I�4p�Z�2�ק$�D�^�;�6l��'Y�uT�k�L�Ɵ|����D�If��Y��ğ�Χ\}��a&o��2���J��<�ꒅ�5+S2i��Y���=!�c_�FjV� �"G�t���9�Δ86GtK���p��9��U���I�lz�#C�/���U��`B�Q`t��ß$�	r�S��l�8�T���D�WD��KFf��y�n�<k��x�m�-z�Wl�8�y���>*Oh��t�A}"�'���4F��WY�,F���ߘ�v\(@��������̩�5Z� "T��'�+�Q д�a�e������y1����Bt�<Q��I'x�l*�S�NPȡ��G��/,��@�G�P���rB�ʲ�:`h²]b<L����^a<���ڟ�$���u�\%x���:I��P�a��<i��zR�K��X>e&1kU�I�P�m�'tў��ēj,�5$�K��2��[�1H��ϓ���Կi�"�'���
DUt5�	ܟ��I�H�j�Y��Z�@�8]KS'�P�Ų�(˄5�<%ig�x*�Xb>�� H�{Wd� �D 3�W�Z������)@)�ya�J ��%����?�L�D"Y ����1�~��'��0�2Wk����؂j|`�⟀�N>E����y�����}���9&�]4u�����K3���`�Ӂ`�J�9�΃�1y�Dx��0��|���5���
�/a�!!�h��K�����?����N������?���?A�� �4�H�beF˞�|�C�"ہt��ԱQ�OT�'mS�$��l�$� ,Olɹ���a�q�1+�l�@���O2A0	U�kY��b��&,O��ڗʂ�]�N�Ŏ�_W ���O����'���|b�'�bU���Շ��4�X�c�e݁���3�F7D�8a	�p� 8�,�u�h�itiA?�HO��Ny�!ߠL6A�}:���D�4�)p�"�"�
���O����O�ѐ/�O���t>ei�E;�����fG(��Y0 l.��K�oL�d8�����<�gMXr����s�*J4�-� �L
龔��
S$~4��7�ayR&�?�3�in<$B�ު�b�2G�]�Z� 6�bӌ�X���9O��h��''-���CP[
Иh��'3ў ����	4B����X��1�v�d3�O^˓��f�iR�'�哷 �0-��#�9 zD̉�/8#�	,�*����L�	LD���O\*[aJA���?�O��1S�	�d���A?>�Z᪍�$ܵm��}����b�܈�+-�I�v�h4QW瘩i�yE�̩q�Q��7��O�0mZ��M����		��,RcoAO�-s-Χt��)�)��<�q� R�f���D#���2�B`~��i>��J<��V7n��
Pgh�Ȃ��_�<���%	$��`��?�.�vّC�O
��O�|`��K�XPf[c�K2}���brZԊt`ʭ%�d��7(���2�Y�O21��MBW�H9�q*��l�6D��@U�	قTF��1Ɩ��D�MlF�����ƺ�f.�!%�p�C+�
�G�>���f턑�L�.�ĵzT�'�6-���Ij��?qb�H�f�ǂ<AN�а�	�(���˟���I�V�0D�K�R@i�čT�X�c�p���HO����OL�ڂ�	�5��P&k\�,��M�O���P�'��e�cO�Ov���O*�Dպ���?1v�ϣ
��(�aW�"!�\RB�:K��s�E�D6uKD�<%�� ���HO���5��d<iHR�8��8D,֦fG
��@��4��!�푐t���+�Km"�C@,&�$���l�5O$���p`����M�!�x��'cbV�Ke�BH4%�Bl�%U�Q��A1� �	�G������T8E��I�l�����$����<��H:����͛�Z(��ZC�ib��Cr�'���'j�\S�O��?���bq��-r{,( ���&a��N��(x4��	�q�r���n�3�,�?A��K,0a]�ŏ= Xh�P!�J�1LQ [V�"E��6��s����0E��h������B�;nBQ�Wi��~@#c�Φ}�Ily��',�O�� rc��ং��*��ԒU,��S�V��&�BՒXtJ��`O>th��ZB�̓X��'V�ɪymB���4�?a���]��F8��U?{��c�%3�`���OF���O�)���� ���9%�'#�$��|���N���d���Of�$�`D��' ~H���Ux�ݪw&˅x�O`�t����9А�铨�/���c����?f+�'��Ohb�QANT�*G%:4P���܇*�"��s�bf�"$�t��q)?S�eд&�Od%�lY#�	Cפx���?X��� b�LC��M���?!+�2��$e�O��d�OL�Ȗ�?7{�U�gk�-hW�͈�Ɩ[�.\j�WJ¼6�.�?�O�1��_.$��9��ܩi9���),1�~Y�äC�#�;�% &L�`;`k1����A�o� (����V���8#O�u�֐����M�aP���0��K��	2r���Pw�S)"����!z����Qx���N�;KxQ���}t��AV+��� �������C�Lȝ�ah0n���F�NDJ���O"�y#�(G���D�O�$�O��;�?���t�r-�' ̩L�N�����,B-��8��'P$�JM�]�y�4�����R(?�A�Hv��@��U(h9���Wr��4x�D�!
�d9�ԟ*�@̘R��(��>�#�+U�B�K�) �IT<I&cP?6�_���Rڴ&1�'��'�ɖ���K�E��Y���(��H�(B�IןJ���+Q�
�ٖ�^S�>d�w��HO0���O�ʓt�P�A��iN��) ��j�E��%��	��йt�'�R�'H�C[
MKR�'���ɉ0$!�wBÀ>�њ�EB�kE��z��|��M��)�P��p�'�(ZgK��TM�@η"f����$���Qdѷ1�8�k�FZz�^#?)1L�џ��ܴd5&�%'��o�f5�Q� ����t�i�b]�L��h�S�$$N�+����u<:�c�oJ��y��9�J�q�Z_��T��N5�yBEk���D�<����9[�S��X�O8䵫fW�W$�X�J	�bd�D��,l���'�bK�>t�}�G�[#qH\ܨ$I\�;ڪ�'d­����_��9X"G�<g���Dybl��Sk-��	�)o����a�%Q��4'�S�? �p2 �	 �D�����*tb�U%� 2t!�O�Dm����Om�Q�ӎ<s��(��Oմy�F ��'���'C���䆞t�l�ٳ�ўt����Oȣ=�'br�'\�I0&���[`�@Xft0��'&���!v��D�O��'KDd#��?��H��ɹ&Ì����)��Ȥ�ܼt�Q^���B �$�[�ɍ#���"��OX1���\�t�#@ls^}x���3[�����C�ty$a؜�Q?�$�l�~���F'�!  f�4�r<�F�O�=lڮ���4�O%�	�S�>�j���j ���t-��'#|B��{մ��4�U4-�-���Ȫ)h"<����*���]�#����9(�ଫ�@�n:���Ob\�3�>���O�$�O�����?�|[I�D@��h��X*2���{���/1u��y��q̽k�+pڐ�	�l�8bR*�WdL�B�Q/x��Lh��6�V��%�'! P���I�?}0޴az$��A'5��d\�:�bq�*}:���V���֋�҈m�4�mZw�}��=;���(3LE5`d���u(�_i�B�	��h�%̀�iq����"^j)K�8	�Ez�	u�6���<)�HD�K��VnI�!3�7�JG��!�E	}@���O����O�"դ�O��`>hr-�6hmx�@u#Y�etDUɰ��m� ���i�
JX���~��`Qï�* R!�U/�(d���{�MϸH!�;C�'y�E��J���@]2Y	C��1�<��nƞ{��O��$�OR��'FR^)�V啲3�`�6D��
�t���K��hl�e��Pw~1�/��'��	*e?X�9ش�?y����'� E�7e�:a�z2@����@��8���O��D3����(�@6<1���oD A�O�L�0�HP�o�8�2��&�.Up��$�%�� �&n\]����C����ŭ;)H��[���Y��s�Q���Ɖ��!�&�"��F���`�nD%>�ɽ\�Pp"�҃U��s�C�l�^��	Q�S��y��� � +Rc܉f��3�����&��|���x��Z�1פ���ϓ"d�\H��
+����O���=<O�Ę�� ;���U�Er���"O
��օ�!c�dY�Ƿb��Za"O:X����.a���w�L�h��q�"O�|!� [�؄ �(�4q:��bQ"Ozd�XYLlc5*<P3��p"O�Ш�nL�u&�b. d���x@"O�����&
E� Γ,����W"O�h� 7egX���~�ʅ�"O����IZ��,�sa$Θ,� }cW"O������z�C��hX��"O�D�g�'�l|�f�Z4a�jy��"O�@��[�` "2,���)��"O�	S�ڧP �c��ݩq�����"O
��0g.<��v�ב\T�*�"O�xX���ǒ1*��0�&��@���y+�?T�l�t%�)g�%��gա�y���U\E�sk�"�ȡy�����ybOšc�8�k�*"P���P
�yҎ�9SJ}sb� ����Cw(��y�nC+TP�%��	 ��˷�y��U�+:����תt�p�A�6�y�5����kvy��k��yҮ�f��8���8gl �y%I,�y��3/�z��L�jF��۔�X��y"hQ��]���!.�"q�tm���yBC�QM(��#ފJ�²�I/�y�⃷yf���҉:B�X�F�#�y�G �>�D�D�<��<+�mȪ�y"e�4,T �@�4t�鑥���y��#C��3�&�%T�$���yT)q���#)ǉ�lk�(�3�y���S|��(�����D�y��]'Z�Fl�T�� m*LP�����y�DM���u.ʮ8�̀���(�yb�U�IBőR���q�4�����>���=:�Z�ka%V��U$��}��"� J6p�fPpth���"˓hY����=y�xQY��ۯR�䖻ב���r���!<������,L)\�v��o� �I��{Ć�ӓ��RN�=Ӡ+O�T_�(�CdH}Yl +駈��$&��dF]c��|*Z>'��F��U̩�f�ǼObBD��DV��>����8`Ƒ4U��9���<w���#&�HQ�EQ�S_�q3�'1f�c��22`��F�_,s�ȋk�_�!#���-���0I����	��b>!!b��XE�Q���H�i��1c`2b�{��;s�fa��~� Up�&Z�f�Z�a����e�=�#A'좤j��O��*W�OSFI"�S�D�yK�����u�����i#4-Ss!B�9
��e�A,e:��O�P�1� �}8l���P�T�X )�l7\��ԏӶzJ��s�h���#���83��8]2�����v�:�x�k�\��X#C�87T�А�3��K��� ,��9R�e@��	��<��ǎ1fH��D@��]�C�b�9�͋�qwLP23-U�Wʔ8P"V�S[��Y��w[Bd;qX?����l�O��Ό�:T�u�6�+y��T�3FZ����%]'x��[!˚��l%���])c�J��%�
�::�(y��G�,oؔ�	��Շ��1sܘ�G�ɨj�]�&W?R�"=1Ch��}���aElE,qi>I��	��4�V�T(&�I*l�^p�%G��)�n���C��&����G?E��'L�9Q�F��tU�u��h��L��4{�J��H��*>��ǽ	�>��ϟ1ON���+<�qA����
G@�8`���8S�N�R���0��xre�5o�����K�Â��D���\�V]��&�;8��Y5$(�)�Č��X�F7�˱"��9#�	��W9�Q!k7�)�A��r�w	�	b�F�#�z�) � �*��]�W�|���~bM�T<��O �\�Sɋ !Bt�q���n��Y�ع�t����ɏ|���:CJ�,wQ�-p�̢*�B��s���ca�4k�
t���'~[b��4O�`�AE?�c��ecలb��	�:����_���g�iˋ�p��m
F��%��i�6 1��
��φ d΁[6����O��H��8�Vh��7O��� ?hߊ5K�&�3(�xx�L8�p<	� �&��kdm��1��P��H�@; q�e*��V�Xg�$��^�➴���/~�!�ʂ�lP�%�b�X?��ϔ�k�� {ci�<{��r�h
�N�LO�	
e�0��1)\1���CS>���΍�5`:�d	��tvQ��'%��<a�4Gi �`m_
�Ҹs�. "1*�!̀8Vdb��B���!��O�pc4g� �Ū�PCbX��UF;}2+-D�<�`a@!<�u�aA���|��t�eI�>t3���El�I�$��%47����!��q��\Z���a:�aq�I1�"h��݅���򄜬6K�6g#�=��*X�� �}��v�H����va5�Ȫ0G�a'?�ia��f�0i�U��.^ZɱA4D��c��S�"8I��_�y����f�>ĂE&������)�8>�#}�'�8�uΐ)�؉���2l��8�'M|���j:n%�Rb��B�s�|���*�n$�Vj�(�3���<pQ�mB�'X�BOd��$�]������t���)�LF���H4�0�Q��1a��VCX$�%b�d�hʓA�?S���h1�U��>� ��@|4HZ�oW��a�'�ؤO`�1	��'�8xN��i՚P�怀1���w�a}k^!o0T��3ZJ$�Y�@����Bq#޽0[0�?� n8B)2�Pխ8w�m��2	29���!��@�&��B�,*��dA�HA����ƠdIQ��I�1򖱱f��c����-�> �X˓F̎P�2�S�D{�=a�h��%��Fy�cül���YQE��4r0=��E��M�6��r�߻U�4xI'ãJ�T���I�@��!q��^(oH��X���,AD�E2'o����'�2���#ؽ{�* $�G2Z��kS S�I}���%����6(	9�đ�ێa�d�V�����'\LXCǢR���Pt�#1ٸ�``W7�^�;�� I-�O��PK�d���]X����$�Z�@|�>	:�gC�:n����� @T�dU��� �L�m�b�Qc4�ӵ72r�bu�H�Q4�s%f��F�zC�ɥS&!���͍c�Hd�(׊6��\9Ci�O+^�;��T_r�j7.ƅ�~��4&vޥ��_DŚ4�1C]�BBl�JC�7+�f�	�ɼ|�,3�nJ�f�y��iΎ ^���"3i�Ej�`�}��+�7fs�d!��|���Bg���B�i;���dW��=�4a�6��(]Q��馅�j����,l��D�߾.�x�)�1Z(���+D��?��E�\����!���f��_��������'x4���'�3������G4~C˿^4��p1M؇j�  (�iă_B�ؓ�&[
B�}���rF=�!��鲥"Pi�g�g~�	?^�P�cD� �T=p����!>�pg\�@�@�#W뚩�SސQ�g�~R58�b��H��r1��ˆ�����&?x�����%�;=liz5!���p<��'�Q*<Uh�¹\h�	�ƅ Y�2|��Z���*��V��\	��L�Ĩ���O�O95��)�[�ic%Z�q�1x��ASx�h`#B��d{��ƴ$	�G/ĸ"g ���Ɣ3"F��\=oD�  cu��q�*W�$�`���O�t��0�?��&�C�H���T%&�d`�'$��y�x�J�/��S��>Q禟?M��M"R)�
N�P�b�R21��ؑ�G�f��Ц5i�("|槀 ���e�\�X��hV&O9δ��0/�v���-}�.�g}bj��n1�:CN�z����
_.7&���kX�7��%�Gڼ+����V��as�M��fBXi0&+@�?�7�N8���@��'�	`'ŉ�D�����1B8Z���5ˬ�2ө�w:
T���|����R��]Ū��]Njt`7a�N��aSFA�I�$��'ذ��'�TiR��H�
�6�%�ti� B�A�ju�q,Y7~T#�lC�u�(��B_i�J~��S�֑$��1�U�H�M��D�䓟 �k̏�����kW����@�K�����Ɉ,�?I����H�z�cܯK����cG�?�'�^ ��Y/!U`h��	#xy6��X��V�m` �r4��Gԧ��r�-8g"�9u��*��0�j<���.C�oX�v�N..���A�N�{��Q�tU"X :����ϣ�y"�����PAwӨ���Iַ-��o:���ˀ�Z;�0=ѳ*��dB��`�	2O�QP8��� vX��	�7� ��6H�/p{{`� S,9s�j[
g��9�k�'X<����i��P�%�&�� �O\�c�H7~��p�� �-ڡ�ɂ]�]�g�X> �r��8`j�ʓڞ�(�N��q�Tѩ��p)*��	�Bj��G�Z�����R�_Z��>��Ń�P7(,@D�Ŵ.�Z ����<�q��"�\M閥�~@ى��"@P,	Y�`ӄ!J��:u���3��@  �a�m�4LY�'���r����Z�mIbX�,G��#UH����\����B$�1Ad!�e{�q���L�3�3�rA2��V�Ek��S$_���iK��%?Q��hMk�uy���B_�@�A&D��Ie\O����$Y�|��i0Δ� ��D�p���=@�7�\=	.Ҹ�O��!K�,Ι:��	�A�X� AK=V�~
���7���˧[�H-PA*�:��P��U,�(�B�.1��LB%kK.!TN�����0����"9�0]�P��P�K*t̳2ܑ8�z�D|�[>j� ��A��=���y�G-R��㦨��K��0��+$� �u�� a*h�p�'b|���}�@�E�A�ֹ���y�Ų^|8�Qtf�k�]A���M�p���d�.$x����;�l���E��,�t��䆍Y��1�m�I�\Z��O~X��� ��-��b�a��rd�T��l��a�L-��T>Qr�&J�L�'TlArPf۴�T�*���<q/P�M>)���1�P�A�G�L�R>�	7A봀ƭc8��Gh�$H:V�@�U��ǓBn�a�OY#�$�!+��5t�R���f�+.[[���[GO�
U��Lce.��R����`�<u��6R�)i�&Z_����O�T(^0ysD19���I���]����=��ʚ+�@�� �d1���4�*Y1Sm+�����pӌ��/n�mB�mC�E��9��6�4u�b�����ӹKq)C�惯6�a��K.��Xp��̅x��C��G�Cx���S���yң��;E�d��Y�Ǌ4��9(U�����D	���MC-z�'1P���kT8���	y��5�'�Сt�6�qӧ� v�&g��F|8�&ˆu���@�<Wz��|n�y��]4kD�rB��n�#G&��G�d�Is��1�E�6�Hy�I�LB�ءfl�M &��@�*7��Ƞl�?.�V�	&DZ�T���i¦�I6=� @�.?��Xw6q4�r�<�BP�s��qBh�1��zR�׼n���Xc NP�֘{��F�߆Q����5�M[�?O�ԛ�J<���B	�|jV�J�M#�ʧ.���ځ��%]���Ơ_W�l�Dzb�U�Q|�B�˂7��qaT'�	�H�I�XdiC�e��{���j1A���%M�`�V���
�6h0������I�pb�ڤɸ<!�冥�xT)��	B�
̩�H���ݲ��j�>9F�K�y�(����/��'��扅~�f��v�V�w�&�J��?9�py�#gG�//|�8fS��j��7�g�'B�m ����q;��'@C�K66�K"L�$C�Y/O.�ژ'�@��F �)�P烯	�([w�P�Έ)tI�����CFy�&TNaa{b@�T��l�=-Ӯ�k0L�?���Б�Ԓ���ў'˄��\��l�i۾�+�O���Е�ĲNE��ؔk'4jE�	�.�<���C%^��yۓ��a�@��:�Ni0�b@�gή�qb�, �ّ%/W��9f��#Z�B��iz�ġa�ƠtO�\���R)��<�/[|y��M9m����s��a��Y(�DY���'��1SR��we����J�!Vք��O��k#E��?��Eɂ�X"0Ph�G ;�Y�G)�9<�ʡ
���!µK/�@9�2�"w�u�-�9͌� �kЁk!p�M�~blu�|�p�Ce* ��ힾ"NF ����0h��a�ŕ�pA(�m�V<D-�Z7����4]R���燲s :����M��3O��c�G���C�!�9m������t��v���-Ov�4@�aUbvN)2�_8��=iE��	��	'���͑�{�4bdK�8�9r�	�ZY���B�"bI��I��~�O0	6��	��	�,Jfh���1Z-D�X�Է�B㟔�R�OJٔ��
�U��O�����&��ѹvn�7v�ĝ#wa !O:�j��
�+gvyaD�2���?��nʱP�0�ʙ�"� u`rB�U�'0�L;��2&6@8�V��N�N點'��A�8VvZ�arh!>ȶ���A��r��Ms�T����,V>�*k��~��V0�e���E��!��뛆���I�-g*�qp&��,H6�ɊF�Vt!�$ �FC���gޚpI`-��#°U!�$, ��A�mD;l9j���LC;P!�� v	P6&-G�b`�B��̑jW"O�aa��֗	X�T���N�5�b���"Oe�r�$9���R��N��q) "O����_$]���AmԹL�vi(�"O4���n� Tǈ���aٿZg�A�t"O�l����#aF�J� 3c�t�c"O(��A�J t�he�V�DR���"O�8 ��N��4�5�ʙBڡ�4"O�h�U��&R����C΋�6�j�"O�C�G����iũ�9�ҘP6"OR�A"k\�`~�=�"hH/CV�Ӳ"O�X�`@F�C΄����2M��"O��b�	A���𡒎V�`�"O�E�e��m�t�
6,XK"O������P���BbD�zI��x�"Oҁ�����bL�c ���E"O8�Sh֞
��� ���&c�lH1"O`TJޡ#.`RDOϿ���h"O( ����l X� �+1Ìp�Q"O��fʢ,_�i�eO�_"�e��"OR�����^��uM\_�n�k�"O��х	7��9�X"ͱB"O.�H��!(���,�?��M��"O� �oI0�n����->�j'"O�ł�B�%0b�S��e!��"O:L��d��	��0t��� �+"O��1G�߲N.���n�&+� U#'"O��"-L�A)������v"Ob�A�6=��L�$Xkp���"OȜy���9X&�IBKڹb�LX�"OD���]�?�\uXJ�z0�P"O���S�Q'V�x,��iK�eF�%�"O@��&!<|c���H�l�3�"OB4ڴM�9ᢽ� Ż=y"��"O�� ��V��$"0E�F�`�I`"O��`��T{��#&$÷�h���"O���dP�1��<`$�O��>�y�"O|�Q`�ǀZ�TU�׮4���"Of�@ě���] +Z-����Q"O�d�tU�]l0�H��55 -�"O��I%��;7C��0��嘅�"O��ʠ��;K��P�@�-f�X��"O�pD
�>`��X�`ъY���U"O�� �-�L �m6lfb���"O> ���"-����˔�W�Iô"O���C"ԣ+Վ�q*��s�QJw"O���CdT�1f�G�L��ŋ"O8�R�d�'T�FY���%*�,���"O�`��i�*u`�{����~��b�"O8ĊၘJZX���]"ٲ�"O~���V�F�I����xA"O<����H��I�%QY���"O<��D�R�N�4iI Ǣ}D"O5��eM#����U�Չ_�ڷ"O����jQA�t��Z���
V"OL�CEo��l}.�[U-߄T~�yb�� G�� o�8b�00S뀔�yB��,��$!���&O'�1aI���yBF�.Ju�!Х&��6"�ӳ�C�yE��8t�Q T��Ks��'�yB��1;��p �i{G�Ѳ�y�H������!)Q�{��pF��yr�TI�
� ��({��Q�AŦ�yB��!��\�r�G�����"ŉ�y
� � s��ެ!��u˗L�,��ȥ"OzY��_�T�P%Z1f;�r�B"O�\P��D�[F��� L� 7�~��"On��I	[Д�����z�($SU"O���"�7^��T�3�05xq"O�����@��B�1�lt@D"O��Q��4ix��RÁ,y���� "O������[��8"�X�>^8�"OR�a�蓀f3�=� �0dN,��"O��X�B-�N��N{/6-a'"O���(�TL�[��?SF1�s"O���mYct~L�e�H�9#,X(B"O�AXG-͙�F�/�emB�[5"O���m���z���փIo:i��"O��EaR6<��i�'	]4�b"OH�*϶��л0h5:7�H�O��D��%�(G)��q�Є�$�!�Z '�^�C���p�:f1I�!��Om�\�O�6I�PhK�C�V~!��K�"*�H�n���Pp�A�dt!�i�b! v/�,���C H�Bn!�$I�>�n0��-LS�r�P�i�+6b!��hp�Z��Q�f������![!��ȥ&{e��*â^y�๶��c�!���y:�1"ݪtc�hr����/�!���Lݾܻ5��cb`����L�!�Ē&-�#G��yW�9X���p!��M�Dü};1��e< E������!�D�?��A
TeS�9ͦ�*�����y��)�/+�Ja	�E1l$�aTeW��C䉱gs(ѱb��:>��Lp���O��p��	*7֍F&y��\P��PP�C�	8�0�h�GN9��K�U��a�Ɠu�����Z�Y�.1a��b8V���H�x�sMĶ=b�l�����t��~��SW�\�pL�A	
t�p��鮭�W�P�s�����K )��ȓ��tb�AZ5"x��c!���ȓI/����۩���0%O�`�����vH
���^��Ha�E�b��(�ȓ���P��O�N @�)H�fج���k�u8�H�l�^����;�B��9��P�/�(g  ���Q ����K�0�l��xq~q��hS=k�P��@@Dy jW��r�xu�\�v�����hO�>!�᫁ �h��5�Œ��)�3i3D�D���Ls�T!�*��o4����/D��C�%�>Y�U��8R8��xB�2D��ن�ϖ^�&-;r$P!c�Z�/D��ؕ�D�B� ���B��W)�Ԫ��+D�0�"��P�JȪ�J��Ε���(D��(� ڨC�z&��I��j�l$D����	�j����G�0'��i�,D�<�6�nNJ�K�o!"�̈p��7D��{�I; �6� � 
O�B�5D��� ��)U�Mj�Hq��c�?D������ft�|S��$4���8D�T`c�D�|�xu/U�2[����#D���U�P#wE(�b��OY��*�!D�${c�K�slre��MI/��H�eO3D�l��d)P�ց��/I��`hʶn=D�$�M��x�b} Q��+i���G0D�� HL��B��D��m"�	/D����)������B��b���k/D�� h����:*�
5q�E32(L*�"O����돣r���j͠Yv��E�'��O�� �W�?I4��I�C?p��"O^����4bv�
�3?"ث&T��F{��i�i�X�r��=)w�0��ϰ<�!�$�QL���@l�F����^k���Hy��'
KQ^�bD�S�I�P1��I�<�i�Hz�Ak��Mp^0����C��'�d�u���X� �#F?��4�=D�l��tHq�2oߚ(x �?D�T{�`��3���
U��~+(�&k?D�����!z_r���'Q�!��`i=�O��J��S�(@jJ�Q��Ͷ7��i�� ��`�` �`D��Y�S�uv�YG���C�!�r�ɚ5W���v�͖+�C�8.0ڵږ�Պ#4��"uč D��H��	/j1�9��H� ��(Z����"��B�I�U�J��s�|=d|�1�W̌B�/�hHr큛j�HL��'w�XB�	($V��5���N�c�)�-�XB�I(9�$�o��Q��*f�1*^C�IY�Ld�p�� &)3�e�.�Ʉ� �\����/���:���_��ȓVT�i���m�֙
� �l����5��%��6!H9��G�`��ȓ�&ءrc^ ��ɳmW�;�R`�ȓ(�0����85��㶩.p@�8�ȓo=J������Y�q�ŀ[0�܄ȓkξ�P�J��?�:@qϟ<-!���j4ր�Ԅ�	Z�JQ�V�8a�u�ȓo��B�)�%b�|��@ߴs�TĄ�.���y@�	�8!9�H���~Є�
���сbQ�`�����h��M��voX�sQ�����y�c��|��Ԅ�ZD}
�b��#D��L�R&Ʉ�!D����J��,��h�����UȄ�
R@�aa"�������@�4	���ZZ�I�e��y�*d�燅d7B���n���cۆ�b��� 'mN����UӬ�C��7�
P���!7��A��IT�'\�z��R(f�l���ÓBK�@�'#��@f�4�"`c"�&6K�5��'���#�ֻYɢe�֧Q�*~�)
�'I� �Y�8⌥�6�R�$��qi�'߼ ��n�DT���g�ߊ��'����G�/@�1�fB:S�(aB�'~�I��T�Te��;��2E����'������ٖI��Tr�Vn^]��'�H9�a� qS6Tˁ�E�`�H��'𑀧��4`��x����	`��0
�'�4ͳ&�1Ǟ�X�e��bZ�+
��(O�|Ak�`˄��#)ʿDH��9B"OT��"RI�p-����"z3&�r"O 4�A(X=YH� ��f|����"O�j�c�"�p9��$b�����$\O^ð둮n�h��&�tU��'"OzT"R�L�9hDQ2�K�N-{�"OvMCX�ALv���f.#J}R�"ObQ��x2�qw ȱF�ct"O�\���ǢУp )EX�(��D=�S�'cQ�u9�f����k�`ӡ'�䑇�]�<2F&?~@��kP�p$���+��<����io4`��fZ�w|U��s�Xi�`��$�V�J$#Q�d��Q��S�? ��� X	b��]Acj��a����"Of�A�b_�E�@�c�^$}� e��"O���3���*ݸ%�j�b�( `�"O+d�W�9"���aiN)����"OI���i�\$��K({y �
t"O�r���u62ܳ6A����9�'~|D�P���ب��'"EO��J�'�
hꄆӾ>Yԥ*�臋eО��
�'+@��
N6��)��m�cZ �	�'Y�5Ar�P.6(n�K!�͢�^�+	�'X����ԕx��$Ƥ��'�<�� ,K�e�n��-/Q���
�'���BwR9o��ؑ�Svx��
�'�����͜�+���Z���&\2�-��'blF5��pSPH�Q�Rĳ�'K�$P��*冲8T��'V��킋D��0	�?3 �I��'�̪A�
�[��=���8B� �+	�'���  �΋G b	�����9�Hhy�'Z�F���~���.�0y�'	v�`���%:6څ���;�����'N@h4(�:�D��ʪ,��'��;!D4Q�5��5(�$)�'�` ;�ŝ�L�̫eB��9T���'>A#䔕�
��u_6|2�'V��!�ʿ���S�'^�Z��
�'5���SF>R�|A/e���3��A�<Y�ś/4�2�XA!�9n�$
{�<R���r��$��=D��+�͛`�<w�U!,�nѣ�L�b�&��C
e�<ɦb��b�,[�K�I�\���]�<QD̊l6@��B�b���be��U�<��N�-�*�EB�!�Ľb�V�<���mxp��Ղ�Q,���S��z�<9�MX�~:��3�$�Fh�u�<�BF�/82���̏�* �2f�Mp�<��%�!��Q�l��e�����'�@�<q5G�Hb&�[�^�- ���gMv�<���2o����U�%h!*1k�	t�<Aş�h�N���E�)h�B�NVt�<�0E��h�����O�V�5l�s�<qf.8Y}��	ä�.}��9��m�<9��]�THz�bT�~(��g�<)Uϙ,?V�
�,�>:�N�`#e�`�<�"k��>�&]�k��?| =��h�A�<1��׷l9b	ȑ��*gհ����v�<���#�5Ya��#_�DhwKFt�<I�����|�f͓8Cl�:vAFJ�<I�3qa�l����1�J��� I�<yt��!Y���d�Q�~lj(���D�<��ΦSbv���a��"p�іg�|�<����8@�T<�șKe4
.X`�<q���':���n� P��16@�Z�<���Y%gK��`!
��r F��w��a�<QwH]^�|�AVgH���p��v�<�&�0����g�4M�����r�<	�])SLPY���H�4{V��q�<�'F}:��0����h�����p�<�ǯ��^C��c ������p�<Q�&�5ʒ��&CU��s���g�<!v�G#C2Y����+;�$��G�i�<��QQ�`��J��0a�� ��e�<1®]/�l�u�Y8:J%����yb��"�Tp1�h�1Q馠AѪ�y
� j���f·Y̖\�0f^0'��1$"O6-R'��<y���6
�;l���"O$�Ueğ�bM�׫5Y��)�"O"| �C��ku��*�
\< EAT"Oj��׆�&ZKr��w,��o"f[$"O�}�#��	;s
Lu�	#E"O�9��jG,6U��+G��9N���6"O�)���9r������*0�s"O"���!P'D���oɡ'�P�"�"O�!P��*b�$�0ϒ{�&�P�"O\���KVX�p��/dNp`�'U�l�C�2\��eK��-�l0	�'˒1��`(T�8eA��zP��r�'��ܘ��R%�x�90���r�D(��'f�("/�k#����W��P��'� ��sfӿ+[��FJ� ���'G>ũ���o�
c��z�8R�'�A�'�#()�Ҥ�j�� 	�'�F��T��eju{�)L�Z#@��'.,���O"f�d��C�c��'u�QsaȃV�,�c(�(�B�
�'}�l��� YA$���a�	24ā�'�u�G�X�2�H�ƥW����j�'�
m��N-T=�5��o6#���
�'L�|i��H�[�!p�����LX�'w����X�s���A7�ة��$�
�'d�CT�G8�}��'�b��< 
�'�BѹD��!*(@@�b��i!	�'p>��N������W�E�h�	�'=tzUkϜ�4��ak�6\�U�
�'�u��m!&�9�p�	*;�!��'O�]��$� � ����V��#
�'�� *�f�6S6!����:�����')d�it�,� 컠�Ѯ/�8�'�M0����	I^e��� qs\���'1����<ck���F��%�LPc�'` Q�i�%�����4��dZ�'B����BF�r�H��Ri��p�+�'>�tkT*]��� �ØO�z=�
�'�h ��Ë.p��օҖi�0�	�'�=%�l]PKaԂd,���'��4�
V�%���e�OK��
�'[N����;��i15�F�z�)
�'��	��o��o�^��ǁu)��+	�'{��B�ENG:�*7"W�m�|t��'!0�p5$EE��|�EL�:r�p�'.�����4�92e6ly@�`�'���k G�*�
� 2x���5D���u�[�h��1�D&O� 8��4D�8jd�I�$�J]��\)[�e���6D� ��T��آ�^�;(F�5 6D��� �	*6�a{v
Z%�J���a'D��Kp�.;I�L��V�?�U��#D��9թ�(������.>����6D�`C���+$֜R��
�Bkb�3 �5D����^,u�	y�A#h����V()D����ƭ���r.�7#�0�*D���D�Շ;��A�F�x�{2�$D����o�%)��`������K�
!�d9
��i�_�Ŵ`H��6&l!��1D	UF�*6�d�T��yH!�Dja���	�v���0p�`�d�ȓr��\�3	+b#��q�  M�~h��sѺ-��i\�:2�ju�h�i��S�? ���4I�8z�n�ۡ���p��LCG"O���%垿U�x��bAd�l�["O
�B늣Sx���bݳMʄQP"O����CO/Hΐ()���>C����"O:%b��;N��@ɖ�Y�(aB�"ODeyg���x����V�A�` A�"O&�@�P�h�,�#�]%	?�]9�"O�͡e.J�o/��g"h>�)��"O��s�D�e�d����h@"O�#��-��t ����U�0�"OLH��V7^,%;��5P�`Dف"O�#^Xx2D����p�cO�"�!��2+(����3~zD�
���7�!��' {#�K˚���a�,o�!�%������P	1����1>�!�$�;[�r ��HٮY"4J�ϔ�}!�D͂A*���u��H:)��Y�m�!�d�+X`0��f�)����`�b !�d�NT@�H�K��i��!ݫT�!��'	eĜ�%
ݘ"�X�B�σ�!�D�&)�d���-<e\�Q�f	 �!�ʞZ����`��]tT`Had�&?Y!򄁿(Y0���G�im��3G��>$j!򤙵iHؤkC�D�M_T�q�I�F!�d\�/�Ms5�ǹ=[��X��ħ �!�dL<
5�a�����]G0R��-2!�\�:� ���O� @Dp��g�N><!��t�Ĩ�jW'7X�0�(��:�!���ct���v#�u���d��Z�!�ę�	w���C�?Sctݣ7h�7�!�#{�.0 #�\)D���߭,h!�$Ť.�l��T��$T�!��䖮R<!�D��V��<�1��~���IP�W/!�$ѐ_��z�@ r�8��璝 !�dV�_��TB6-E�72HÄf�2�!�$M�L�"X��GO�p���+aE�{�!�$�U��5P (@�r��xt�	Cb!�>"�8��9$�M䃍M�!�$[#C�Dm��E�3S`�'�$�!��^�\kTӁc�!�(�
4.�,B!���9l�($�� ����
/g!��H[%�;�f_1��H��>6!�do���jUDJ�$�~��.�ca!�$P���P1�ʃw�(bC'F5A!����L�{� at��J�K�#P1!�dմM��id�RXj�1p#j�UD!򄔗BV�8A`H*Gw��c"H*�!�D:nIz�
ׅY.Z�Ȅ�c[�0C!��	Q��;��*5�L ���(@!�D&R�DlG#�;>�d�[@*T�3!!��_�Y9�-y$��or��&J�.6!�(0���w$��k�p�1V�� �!�jaF�+�g�#�
��%ݔ!�!��Z�#�C�.���T�Ok!� +����4T�V�h%�̓E3!�DU�� )HU@�	��� �?*!��U:nj�C��/S�P"�O�%p�!�N�n�a�4& 8x�AW�F#T�!�DK�qj���Q�tn���NJ��!�ă�G'��*�E�eT�p���{!�ă��Bԡ`��j7�4H6%�,|l!�d�6?J�\`j� �*
 ES�!��@5a���0��]q(lf��� !�dW�vz�Y@��<:i�����1!�!�� Jqs�/ʼ	M�h�cc��aDr�� "Oڍ���Mx��uA�+A>�a'"O��ҡ�B�#Yر�2N�A�|��v"O���6i��	c͆�:q�"Op嚗�(�J�
��9-��r"O�,��L�z8��q'���&���z�"O�x�V���1�q��:�z9Q�"O���gW�"Zj�`My�2���"O*��r��X˄\�����c��U+'"Ov8�sCӂ��-�1��,EԢ�T"OX�c�"Z�5����
�ty��"OZ��"S�8�Ԍ[4/�F�05��"O����� ��fnR4��z�"OTd;�L��b���+G&j�`,�"O�*��N�
gb��QҰr$���4"O�����?3v�F��:f!n�z�"O���V&"�2���_�9����"Ov�Zbn���xW�X9t �"O��R4GQ;v��bҦޥD*u�"O�L!tAКc)�X!�.r^U��"O8l�G
]<�8ғKA8@��(b�"O�%[0Hܘt\� p�J��K~4���"O��9fH�[�bp�n�2bi�Mq�"O<! ��G��سdǎAKp�
G"O�U�t@�A�$�!�bo�����"O�1I5��Yc��Qd����v"O���٫)bi�"����]�"O��"p�B<lb��PC	>8@BC"Or�jel�9!h�l�jT�i�Ɖ�"Onj�<Z*���5�� Ar��i�"O�	S�
�2`�5��ȇ�� 9�"O� �&HJ+�\%Q�	� KQ��`"O,
��݌y�LL��Hݦ��q�"O~հ��0/��%�.��q�1"O`��Ɉ��&���F,���"O�`�p�<J���e@�v�~ɑ�"O^]�`L�'��M����S�:1�"O�h@�b٠)��ݳ��T�.{`��A"OP����g��q��ߟ!P|p��"O��1�o�	k����T<8I��"O���ǉ�?ؐ�12h9 �"O�q{t�:n�jl��nD�9)��a"O����I�:6���Q�H�{����"O��A�C4�[�� x����"O�i�N��B� �����rM��[E"OH��~]Dl��Уfִs�"Ot��"6Y�UB��Љ���3""O����	�(A���"�1=@qqd"O(�`Ɏ>W��a�F�Ha�p��"O@�(� �0e�*� �:���0A"O �E֝"�6X��n(u��l�"OҸ���7"�`�6��p4���"O��@�ɴ"������EZL�g"O��R��!mO鹳���pB I`"Oj�@v!v��}x�)�1��hW"OaR`�F�B<��Ɉ,�
`�"O�U�q�K��Xx�eHց]
E
�"O"�)F���<���us�\��"O�I��n��4���ȡ��3=�>L4"Or��r#J�t�9j�R�v��yv"O�U�aN��	����7)E�|�v�I�"O|y	��O
&0#�%�)�a"ORlx d)?
���Dԟ$xڠ"O�yI4�ۆU�zy�qTyh�k"O� bh�3��+@��7��+NRF� �"OT��e�iAB�ad��/�)�"Ox)�ǋ^5_ i &	ˈi �%��"O��õ�2Ii6��"B?J�d��$"Orn�,��񬁎m���[&��/R!򄖬o�D�Ke��9�ZxN�Am!򄎀%��
Q@E�'ٞ����;^3!�d��e���a!������9!�D_�/�&�y���-�X]K��G!�D�_�Ti�c�Z�^x�|��\���$B�������:�x1��ܟ�yB'�T�i��M�}��$���U��yb��s<��x�(
�q�"Bv@��yB�ĳ�R�	7���8Aؑ�K��y"ڀ|X����ꃫ3��tRF���PyB�T�3Մ�1v��f���c�I�<Q�
��H��i�׋�;͜��I�D�<Y�P(Fv��fE��&��rTMWB�<IEӆfuVd���l�:t!��Y�<QA�֣YM� xE�3���#�YZ�<�΅��D�3'#P�i[J	�&+~�<���� 6"h9B��F�!P-�O�<Q1+��lab�Q8�N���/J�<Y��;|�|z�E�yp�5 S/�F�<1 �RZ�$�2պ,���c��E�<���B`^5Zp�Z�l��	Ӈ�@�<q֍��a���j����f(j7�E@�<�S8x��w��Lm����<a��C<nO�ٻB�?MD
�Ѵx�<�s";z���䏈�1�Q�AdUt�<���(o/
0��'N�N����i�<�ڇ���
`*Z�F��0te�i�<��
��,��i�t-( ��a�<�%�=@!|�H�LY�O����Á�T�<1�N�$8@4{��_8o"��6u�<񔅎x�`��͖�*s�T���n�<�� �}D��;#�<]`��B�<Q���Gt:����v�1���<*�>� �A��E"X%�G�y�<���Z�p]b}K��־`O�|q�	�]�<�S,�8�R���8%̩b�@��<!ڽ�iZB�,#o�MJ���s�<TGP���&ڦ=D�e8@�Ko�<�3�8q�\�C�I$w`t�b�MT�<qR�ʾy��9r&�df* �$ M�<��4
��J�i-��p`��}�<3%�q ��!H͑'����B.T�<����U� �Z����9��B�N�<��l�T�̩E�B&�p�!�f^d�<����3z�h�"ܷ���� g�<9 ��:`Z�ea�C�� ��BgEj�<q��%��Q�K^!}�p��V�^c�<	�.ȸ `�,S��V�0h��gKv�<���$�JE�C��.�Լ��r�<9Rn^�k\�1c�f�Y5�����l�<�B�T2=w��A�lT�JZ��WEGi�<��m�@�1Ƅ�_e5��F�I�<��/d�b�筎	Og�a@��k�<�d��<�,�(��ɇH���r��f�<��o�',a�'q����ōd�<�3�՗��i�ifFi:��M`�<��d~:�x�aZ���5 �s�<y�Z:
-zA@q�϶�����q�<�Q�B*P�J`�'풰k�@��Tb�o�<� ��GE;Jɤ���a���1#V"O�e85l�9R-zb`E	4�x�P"O�8b�e�1�V������4�Zg"O�xЦE6 _� ��6�t=�"OAʶN� O�u#媜�6/�
�"O�y�
\�Wc�A����<�b�"O��ۧɋc L0Ȕ�KP���2�"O���pLR�sv��uaC�@��HK�"OD��H�#K��-JR�E�;���"O�q���	]t乑�M�tפ��P"O0XM���R�3*�9
���""OX��J04ź��0�͎�F���"O��z�J5Z𞸹�f���BI��"O�i��Ap�d�Hw�]
�"O>�C�y�Dՙ���#FY��t"ON(�%��&o�B�-L�i��"O���D��&x&��SI˿
�� 5"O5�����XH&�_�A�z�س"OPz��F/{̩��Y��ڍP�"ONA ��>,�!���	$\��`"O�L�v�u_0����67R|�D"O�pI�`S	�X:r. lGrQ��"OXp� I����!�OE=����"O��ЧI��o�d)���Ү�Ї"O��a�i�?ZL������f�:b"O4@�j��	-b`څ�׍�*��"ON� ��s�6@둈�>E>�Ӳ"ONā�)�-0�.ͫ�(?���"Ol�hf�Ryjj��t,��$
����"Oh�B'�bV4�b�
��,��b�"O.|���-N=�����#"O�HDG,�:��J��0�l�"O 5�w�ѼVV�9��B#*`HR�"OF蓰�Ƨ5������Wq��q�"O��qg�,gdމ��억G���3"OH���"�%�VǶP�|�""ON��$I�v�z�S!D�gg�١v"O�UjSl��bP�uC�	0d8�	`"O�Cf�_�(����b��s�"O�T ����:��
� �2�!�Ė�\�&�#q��)���� 6!��?g����%�T>{�P�	C��gK!�$��n�"E��D�<=�����05��$@�M�t�yƀ���q� ���y�A��©uj2H�^�X�����y`��%T0X�G��6
,rccH��y�I���d��eƑzh]���E��y2�ө'����uᇶw4�h*�*	�y�!�Lli�waZ1s�X"�D>�yeR�zxQC��fp��yp���y�N�03��c��:\m�MX`���y�ꓬW�r��6��+?��aw
���y��5\�	���O�6n$8	��4�y2���`="�!c�D�u��I�
�'�,D)R�L��%@�*�+!�Z�p�'\�d+eƉ�Z��yQ��J	��	�'�2pID�/}ir�*B�]?KRt��'2���P�`y�mh!�;]}�(
�'�� A��2�0(Aeݦ p���
�'�8Ѓ�ŗZҒ`(�hM�{h&�r
�'s�E��J;�� +�e�*u��
�'�d%��C� ���"V@ʿv}[	�'>�z�ӼC�Ee��2��dY
�'�F�"���(s�t	8M�>��L�	��� l;d�,|7�2�i֓QF���"OlX�7,,C@��wc"_��D"O�j��J�s�l�A�ÕEi�Y;�"O4H)�d��nw��(R�$XhX��"O�cV@�(s.��Е�ͳ3C�H�"O�sj�I\�W=W/��*�"O̤�so�v����M�:U0��v"O>���53VD0J lY�h��Q�T"OB��v�7>�0���H%j�ص�"Oԙgd�Pi�h�F���r�"O:B����	XHƭ�ĥz�"O��@�$�j|!�'Cn0S�"OJ�j���㞈�W��$z�"O>�##�SY�vtJ�,��n�h��"O��SZ�0���+��L���"O(9 �I�*_�z��&����2�1�"O,�PRm�32���h��o�r]��"O"9��b�>�҈�FgK�0a�IT"O��K�HQ�:���{��L M�P�"O��
#�:
�&E*R$��1E����"ODuP���<j2�u���'��IT"O ���ƵX��i�!]�	��hb""O�%�)h�AR�C�g�,�"O8��և��L`1Q��hM<��"O��W���D<x�l���2�yS"O�Ys���*�ժӘ$;���"OD����[(�8|���}���0"O|��r"��
�V��G@�'�Bb�"O,�C��1L������![Ҝ�%"O�9�E�p[@�W�EI|Uk0�_�!�dT��J�jv���`F�9��Z?�!���c4`�[;f)$��`�-+!�$��CUQ"�I(2�f}Z���!�#x$���qH�#%o]�Ru!�F�&�v�� ��~&�0��U�@!�޲CrD�7��=����X4!�L�dg�QS�͚Q�L����!�d� B�*DBU��b�N��G`�RS!�Y�k���`fEV�z�! �G5.(!���PvA��$Z�DL�͙3L�!�dR�;�����E�r�l��Q��r�!�d���C�A��am�D��o��~�!򄗡m��s5�Q�>C���k�{7!��ܥ%�f\����2�!�b��4!�D�U�5Jd&�x�.Hr��ř3,!�$\M��x���:�0�v�!�D>h_b�BA�7� ȣe���5Z!�7V��8h��Ԫx��P!�ӚA�!��?;O���景h;䡺qF���!򤆗Tt�	D(�S6� 3�!�!�TJ`aBO�}�p��pL63�!�D�2?(�+��߇젥
!Ȁ�Y{!��N�v�����oK�RHs憒 �!�Ên�ސ��l���,1`W5�!�d��r�b獍^^$i���Q~!��0O'�P��hޠ/�H�H��t^!���y&p3P�Hu��`���5hT!�$�(��DY�ʒ[�&��5NG?~B!��J7�,�&a�3\�����Їx'!�Ջ"djx2� *f�z�(�	���C�I�xC4U�"#Ò�-��F�)e�nB�I� 0S���>r|����]��C��b��H9��
,@`T#��vC�	�v(R�.�R��A�H��]� C�)� 2�q�	�R�*��& �+]�n��0"O��Ӑ��"_T�@22��.�F%��"Ovi0!(�]C�X�pL߆"N��ڥ"O��xuN�K�T��dL�':5�,Ӵ"O��a#�C�Y���A@�D�v(l�"O���+��e��	]�S}FA��"OR1�#��F���	�\u��V"O���ch7�@�Ζ�(���"O�1r���(��L��-H�pj�"O�<�iۊ��0@Jw����"O�a�Äd�x��r�(���H�"OZ]�i�:T��C#=�QY#"O�xqgH��1�&q�7j�I�n���"OX(HƋJ��nd�ۻ	�mR�"O��3�k�:g�F��F��n	J�"O��*���ڲ���G�t�Ȕ3�"Orl+Wȇ�:v��P�IϬ��"O��iQO�u�I�����"Ox	� �-M�>D�$6}��X�"Or�RQ@2����R�B��=X�"O��Sg��B�i��C3o��E�"OZ*v&N�[�FU��F��d��]"O�q�*Ǯ}:<L�t�L��ر�"Of�i���!#4 t�V	,֮4a�"O*�JSL�$e�ppB�՗t�:��"O�H��KH�(q��0��V=5���#"O�PfS`��`��#}>�R�"O�Ѐ��0�
�2����[j@��"Of��b&Ͻ5>������We6(�V"O������!��� Bܛc|�a�"O�!�	>��aQf���0[��u"O�U�����a����0g?H�u"OLep6oK�b4X�v�ܯi�:�A�"ON�z%A�+�4pT@��,��-r"O���j�"v��`��M�'��S"O��枾�2h8�.�:��-e"O `B��Op�P����I�y@"ONu��A�$k�A�Ơ��W���y�"O\�(�ƒ�M�=�������H�"O�� T�G�c�l��ǉ��+���"O$��Gh��1tJ%BK>�1[�"O��t��%0�x��ʊ
5bU��"O(���cƘT��P)HkC����#D�\
��P
sꩺ֊�Vն�`�7D�Ԓ����s��2
n�S1D��Xw&�H�A��G�i�y⑍4D����[��68zш� �px�3D����數4f����-���,D�XK#C,bn�<f�NS�cĮ'D�$XG�ڳw�="Ģ�6,5���0D�P��bK���R�a�<v߈2p	.D�4�C��!)ԼH	A�]�I� �*�*D�ܪ�f�$]v��y�)GS3�,Q6�(D�� ��w��i�q˹.�,ۓ %D�Pi ��i�nՃ�K�cI!D�t����*~>� "��h�@��A�=D��sBݵ#I8�" ƌY`� 'J:D�`��+�K�D}#�BD�O�d��o;D�jC�V.t
�Ph�K (tE6!1��5D���Q���A���#g��8-*yJ�!D��!�B�u� )� ��M��*�!>D���u��
8#T�UO�g��ɠ�=D�t��$�$q,�x��$(r�<D�\A�+����%Z�À�!��h9��>D�� Pd�	�=��˧H�z\XX�f"O��PW I�HTrҋݑq�Z���"O@���_
]E*xBd�8�4�#"Od��Ι�G�y��$W:X�\m�"O�9p�[7
�eZ�A�0���9�"Ol��ѫ �#8�ӡ�U6!�]��"Oz4+��K�88�8�PS�"OP�ZV J��NH �ˀ3�\	��"O61���芣��	n`H���}�<YE�=Zb0��FH�>�E���_o�<a���:ǲ�� .G��h���t�<��, 2e艑!�)Y�Ȫ��Ut�<�A�L)@���v���x�	���G�<!6@�y�� ���Ɓ�`�Dl�<�C	5&a��-�l��$�R�<d�#�������a��UiS�WM�<!���za�&����F�\w���=��"j c�$0ʃ�;�����:���kg�Ιj�BdlJ�qKl���?0|��Ǝ�%L|���/0�ک��"W\@H�E�~���������ȓ$i�2aC�*'"4ёՄ�3GH���j��x�D�9�J`A��X\�h��'*���g^o���&A�pb`�ȓXTl��-H)<�x�c��1iT����Q�z��7��lʢ����/;l�q��!�P9���%#9|L�*ѣ �h�ȓ<<�ur!�:R�<�Q̖���ń��x	I�ԷZ�]�R�ּ����m�\s'��8?���fK�1~�@Y��a6�-@�)F�`��J�l1aW�̇���t�7��a
����0���ȓ&�:��㙪a �j� ˬ3�����q�!�h�<:��M/�t��ȓ*��x#!߈y�V���aQ�|)��a ���1a��6���
c��ȓzk��"4E�%,T����"O�Ek`D��5f�m
E�F�F���#�"O�X�Ç
E1�ܻ}`lz2"O�Ͳ���B��iŎ�W�*5��"O�0B5�I'U#��!�ޖ[�$��v"O0����u�p�a܇tRh���"O&�����Z���h0@�-[;�xI`"O29���\n��}[��݈�|=;�"O���EKMh���U
Sg��g"O�����1����Í+`�1�1"O�����'k�[Þ�}j��"O��6��+(�ȼ� $Y�||x��"O���Q& �4M�sb҈t�)�"O�����ޑ��e"�aU�t)�"OT��M�8DN"��dG7)貵�5"O�!��Ɛ+
rD�b��dվ=��"O69�ŪB?P��ph��0�&؃"O� S�o�� Q P�7�"`"�"Or�-۞2W��CՃ-7D��"O���r�B�i=l� � (J$��"O��xR�(��,
Ai"9�G"O���'�D���g"�k0u��"O�ԈvH�W, �#�a��T�A�b"O����aS��	j�-02w����"O����B���1���Y.h35"O<�#ŀ�8�&����@�:�3"O� ��h\5 ��}!��]s�\���"On����L8|UP�	�*�()�B"O�  (�+�@�N�����kB60�"O���#�[]�	Sq������"Oθ�m�@жT���L�wꌅ0�"O���Ə�jOd!��͸H����"Of��6����2)A�\��KW"O�u9W�K�j���R�2=���"O~�q&���5!{%��9���×"O�E+��X�X�@4���
5����R"O,��͍�bܣ��W e���cV"O6��c()9H]2>�"�ZU"OZ�a��ܘ#�LH�T�)�D�B"O�r�/D�(����J��]a"O�P��%B<��(<�(���y�:qR
��TZ�
	�V���y���MC�� Ϋ;�� փJ��y�Ǘ�]�0��,24��Go<�yrm��l�d|�Q��1$�];��G��y�ԏFL�x�7�ǊwS썠�BJ��yBM	r�|hsR�iq���̎�y�'�!��4�e"�m����B�V��yb�R�|�[��7�<���'�yBV�~ev�s���x�n��MO�y�Q�6��A��BQ6q��&[�y��ʤkhQ��)?4؂�\��y��Sb����$#H7Rz8��J��y�靴2]���I��*2GZ��yR/@�|z�O�{t��PD��ybM��,0�`�+؃#���k�gĔ�yrJ՜%$pp��m݇��I�U�B��y�G<��t1CA����S���y�Ƈ9:=lu�2� 74���BoA��y��*�A��M�.�}9�K��yJ04]��e�*�U����y��Y�
_b����&}�A�٦�y��^5|JBl�VH�p�����S��y+���}�TI)l����Ř�yr+ћIp��
�	9j:����N��y��G�ı��%�Z��Ы���yboI�_Вu��G_W&VH q�T8�yk��Nn58��	3N��8pk��y�(�2[��X�̆M܎�R�R:�yb�IF�!a���V��G�'�y��}�6XSb@B�x?������yR�̱H٬�4Y�;�򁈖��ybJ!��ps�R�,�L�b�N���y���4KH��bM �%�^!�"K��y�ϋhvr�(d�PE�l9%�G*�yra�-�;����DGQ[���y�*Bp|��ٍQ�~�X���y�S�F�0���?[��=aӣ��y��!T҆a���Xm��x�n�y*�"a���V��&U��8Y���y2-��!�����R���Js�̉�y"�C8w"���$P���Ȣ� �y�(Q��@�`���[ypdS"$���y��'G>zM�Rٱ K���y�X�	�H<�f��z&�[��P��y�"��8��g���b����y���)��P��ײo����AL!�yr
$C�D��¸j��M�)L��yrɗ+i�taP�R)a?�X���ݩ�y"FD#D��>��y£J���y��F!�ڙ���_�F�H�R���y"g̥�(�� �ZMOV�8��L��y
� �aG���'�u�"H	e3^��"O@59w	J}n���f�E����"O��c�G�>�΀xDŚ�7I1�"O�����)t
4�[5��9��"O�Ro��\�&��r]�x`"O�`lľ ����"k��4RY�"O�P�H�$6�$lsrD $ $���"O��[$엣B��hk��E"4�x2�"OФ�����F~�J��R�r���B"O��E"���t<iT��%v�V��S"O$уKQl��xJPc�#o���!"O$��d�4T��!¢ 0�� ��"O��$Ƽ4Ƒ����wY�%��"O��Ã��Bٰ1�V�Ή4�n�qt"O�t��+�,]�� Y�@F�$����"OZ�:�K�0P<���O��s�����"O����M�0S�.|`�Hڍ<0yQ�"Od��u �F�f�z��^2<�p'"O��P�ȝm�t�Ä�/$�I�S"O�1t(��w� D	vU�����r"O���S*ښ#q�0�� ^�����"O��;օ�f��q#2y��h��"O�����[�#�n��NS5��Q��"O>�C@��p���&ȐI�M�!���c���)���;Uӂ��2�
)Gz!��8���W���W�.4c����O�!�$óCI�����B��
�P5"T�U�!�[(*-��H��+<�:���A -!�d�3�&i��dB�z�j<#�MV8q�!�(r[ �*e�Fdp+���b!�2W�<�:t�Ƽz-L<h��5�!�dM�t�2"�7-�	@��2Ct!�$K�-\M��%�x#��XR�U�=�!�DŜ1�P�$)@�]#�/�=f�!�dF� ���Fɭ/#L ��.�y�!�D�Lp�0y��׫Hx��Q�ظC�!�$@�"��dK�(Jl26�R�P�!�$A3�@����&0��s�f��!�D�n�:�v�V;t.@�G��1 �!���%:� �8�\a|��X�Q>!��ȋV�D�02j�]Y��Q��Z�!�䛪n�H���ܘ	*ڀ�PF\�_�!�d��a�� ���܎lsd��,Bs!�$ �.��lД�͏r�d, �"?G`!���>��a�3�	�
��ua/LU!�D@<C�t�2�В����T�gK!�d�?����b�Θm��H�j��H!�$��e�dȉT��zy&�$�J/MD!���1Pr��4	��2��"N!���.R�	�RGW�k�<���5!���{� 4�V�9�:�["EՓj!�d�Y [�M�X ��	�<R�!��իK����6c�DXz��!�ē�Q���蓊�"t�6�#�U�$�!���LP���6!ʞDK`�Ȫ j!򤝲e�X�B����t�a�&fi!��8�hD@��NZ@0kS��[�!���s���P�ʨm(�Y� ��0�!�d�9X²�H��P���ܪ��#/�!��g�`<�P����<`��g�W�!�ē)0��h��цM����fD�qt!�dK�o����JօH�F�w��n9!�T�ot	R����,{���)�#O7!򄚱m�Ɓj5�W.HQH��UȐ�0!�� �����K�+Y�H���?_l8�"ON���EJ�#�fS�Ph�2�"O����bW0�%)��?-�У�"O.���E�P$0p�a���$"O�cȢa(^� ���7h#���r"Oj�3�\�\�9:d,B� ��#"Oj`�#j���0��ӋZ*����"OjMA���qe�����TK�}��"O����J3$��i�`�)&��J�"Oh%0��A�|�����5["O����ό4�`a��D�^��iPr"O
�q���5Al9ӵ'ƿ*O�0��"OX�����|�$����]#	���"O��T9~
��DO�g�QK�"O^M�i^4����Ba�R�@"OL�v����\��Q�4yp�"O�ȩse�R ����	q0��"O�$r��epJm��ʔ,���D"ON����۬zYJy{�)Ц(�V��0"O�p1F(�!G��4.P���5��"O.���J��=�j�4.��� �"O�����ڬt���ӱC.#��c"OU�!��@��AH�6Z���"O@�ͪ dE�2�W8�(�"O!B0�	�u1���g��=�*D�c"O��4kK8jN���M��i�K��y�l�&b*��Q쀟X��1*0��y��W�&<r$�d��;>��<�L��yRς(yt*���0���旖�yb��8V���0ɇ�%�`�;&���y��\�P�88Jքb�
�/��y�(�5?�A�`c@�
i�Y�V��-�yR-�,�dQ��^n���SB�y��8�4["E�N��`�Ì>�y�C�j�p��`��JK`-X���yR ��cm�h�5#E>�]*��yb�X9d}�0� T\��`
���y$�/
��(�5͝~��ʆ���yRDɲl�\�ɰ��*�P��y���kV}b�'H*�а!J�.�y���<I������k���y2�B�7G��kH�~�l�
r���yₔ\��9[��ĐBШqf����yr��tV��dC�)�n�#���y�G)6�s�K�'�ܽ�t��9�yR3)��|��G&j� ��Δ�y�h�8� hj`�R"F�����Ͳ�y"��;�pL�B�ԫuʲ��3jK��y�\à���I:rĊA�a��y�� N�Ma���h���z&��(�y�-޻/TRbMΪf��E�[��yB��cD  8!�ɝ[4�p��[;�y�B�mE8����Y� �
�,�yR���]��,y���W|�욶���yr�Z4���/I��6�Z#�yM�/C�����LEƱ����2�y�,L/AR�s3ƪCdvpyU.I��y¬��=~���^��eC {	���
�'|�As4��/;��E��#Gx� �
�'�n����[�,��Ɔ�e�-r
�'S�ӀL��=�
��5���t�	�'!������q�3�X�
��P;�']���u̍/[0$gJ
�P8|���'#�1��&��S�D�S�O;C������� P���K̋n,T)�D58�tlY�"O��i�Q��,���DY6}:���"O`˂ˁ$�
��7f ��s"O4���EZ�;�^�Id!ӌ)iȕ��"On਷@ʞr7���U`ۂ=Z| 8�"O2��oԍ�
Y�DɃY5�x��"OnP�ϛ�R`z�lM�O4��xq"O0kmP,#�@±�8T1��:S"O�e?���"5z��p"O���T$��fz��i��ҵ��"�"O�x�'jʌ=�m"D��A�l�(�"O�D ��$�@QSE ���rL��"O�Qم�уs�D�sn6i�(Q"OT:Ʈ�*�JM��Kh��\��"O� �@?�����ʷKC���"O�����Be�8��I
[�Lb�"O�6DS	Xy4�)B��zά�(�"O�q�r�^�W�Э����4��]S�"O����`�4<�B
��<I�\��"O�P�r�j4���I�p܄�"O|3���,���듨����9�"O�h� Jՙ<@�@;&TZ( ��"O\�0��JOF�xC���#`�TRr"O�#w�@���nLv��"OdTPp��l�Qv�Ǜ1K�	�""OV����RU��I��EJzhxU"O�1�3$�|���jE냡A�Ҕ#6"Of�'']%HKb0�R@P�R�}�"O�����W$��hBAF&J`8��<�4���B܍kb�
y�D�k#G�{�<A��;�l��&E��o�N=�u�Q�<���H���+p�(k��l��IWJ�<��/,�0�PTe
�p\e��n�<1�U#�z M�oZ�-�6%]^�<�E��(c����K�9Hy���W�<9��#�E��bݻ��u���]Q�<�co��~��@"�8�0��A��N�<�T.���)#��4��(�a�T�<��'[�o߂�i��96��ـ���w�<A���[l��!2'W���]`u%�v�<� �@2)Z1�@�I�~M@�Ǎn�<���3�2�I��Ϸ|k>�#3 �f�<qӁ�o!�	P��6"� H`J�w�<�%��?�
t�ܳ%�i���s�<���"<#r@����r&�d���e�<�1@A�X�J�Ō>�6�CKb�<!�e�?B��4�w�	<Ih@L���UZ�<�G+��F��\� �JY�@)�Ԁ�X�<ib�JM�8�	�)�G�93i�{�<Q���~�&�JoW��yd'x�<�7JH�c�й�%AU�����v�<q���V��3��PaVnS�A����ȓq�ҁ��h�ۄ!1�Σ^!�هȓB��0;�n�26qF��Vb!ҶU��.I��`E�Ξs�H2f�� w�T���#]Z���"ͫo	�RҊˠb4��ȓ,:��g,m�~���n]�HπЄȓP�؄sSg�]�����By��)p�ɗ�R�W�pA5�؎Q��ɇ�z.�9��	U��IYԀ�?"p���n,��)���Lk��W8`�h4��A&Ĝ�!N��40�c�����Z:dŪt��63Đ`��H����fP����rx:������fц�S�? ���᠙_�괮�zfҵ��"O�Y�b)���6��9MP��"OF�*	۬=�)��>>�}�"O�B���e �����E3e/��@2"Ol��4JL�;���ɓ1'"�k�"OT%a�N	���kvK �Mt��q"O�� ��&h��q�Kqib���"OR�ȱ�g����tI��4��ye"O��zw/H�GJ���Ǖ�#1� ��"O�=�6Ir&T1[���d"ޥk3"O<�2��*2��	a�R|���P"O���KD�)�k��':$�WK;�y��;B��۱����H����F*�yr���:$��|d�Dz��U�y�CR�t�A!�#Y�>�"I�!*J��y"�'b���ߚ'��8�@*���yrl�
 � �s�	��$�����yb��e��T�sɪ�.�z�/I��y���l`H��%��$��qW���y�*�>�ś��u��HK���:�y��P2S'���J�q&F<z1-�.�yF'n�4$�4��o0����M��y��=z����L�w҈�ZǗ��y��'VYe��h3��*��7��Ea�'HZ���闀WJ-�	�qu����'1������qk2H�E�۽Q���-O��=E��@�?��)�J�Ц���D��yr�'V�=�����tyi	wK�`S�'~N@P�.�:{��P�ݾ��a�'6@�"A rl`���y.��(�'�>(P ��7G��9��鏜r1b�B��� �H�N�X�Ƌ�i�h�:�^(U�X�n��h�W�)ڧO�&Y�7/Գ_V�kp)V*P��]��eP�*eO�]����H�$,�ADy��'��ؑ
�`i���6���fC�{�l�Ħ���	�h�8!�C�4"X>|�׋��f:�C�I/,J@���0(�$����?Q�~���/ʓ H�Ң�6J�aH�pG�$��IjyR�16�vУ`

�d�ȓ;#^0Cp��3��X�����"|���'��ᓌz���C�ȷi���B�d?^�7M=�h��ݞ<Fl����/��Ӏ�;D��`ቂ�E{nx��&96���(9D��[��ښD2��p�D4z�^$:`�5D��*�U24�X�ӖE�5ÐU��2D�`*W�E�o\�J���4q�`�&�hO?���:*��0��//@]�G	Ă(0a{�$3&`@Đ�d�e��o.!�D�&H�bP���I�k�6�'_�D�a}r�>�QN_LF(s6�D"x�R`���,��x	���A�҄��veG��&�~��)�'FP(�p���4 ���Qj�3D��H��IFyr^���A�C�T �4pPJ$fhy��ʹ>q�Ob�"}�ecL7FP��d�P����wc_�<Iv(R3VH�]{��L�8����]�<֣�0)^pѥV�� %	W�<����a�`� ��?6eh��5^P�<�7�K�$�j��?9��pF
K�<i#��3�z)�6�S=lP�첅%P�<�vB
<" 9��G�WtL�5+J�<!�c� ]@�xS��#=��%���C~"�'N��h�zXѭ��|� AZ񩟝T��h���A�<��h 7>�ua�P`f�e�D��E�<q�C�6�ȍ�F�A�T�]а,MD�<� ���a��(���p��78F��D����ҋ��S�z�Fu)U0	�Xx�@�Pg�C�I�e�2MP�nRa`��/��X�<�a}�₿z�����AM����m@ў�|��O���6+�xh	�t�[�K�(�"O��A�f��t�Gd8E��I�$�<���E�#��Ұ)S�9<��!c!��; ����(."��#��3�B�	�v���gB�#L>����ZC�	�gx���]�\2����[�*C�	%p)��H���vY���]O��#�'l�|��S�O7�M���1f�r�pg'ʐ��*�'I�|��a�&��H�6"ԙ����
�'���afQ�X��L��n�
�tP
�' � ���,P6I0��/=��{�}��|b�ӻ=H���&�R 0`<ţ��Y�3#�B�	)\�į�q)֩�T�զJ�B䉦(����qo�F�d%(�l�C��C��>�T��1d�
�����[xϬC�	�Y4ke�(sH��ʐ�E ]�c�t�>��5�IW��K`�	� �����ƊC�	 gT|��s߸�:7f�  O㞈Z����D� ����
[�%� P4C�Oʢ=�O"�1��IS<��ɐ���;�!$�9��'+��Y��8D�M���3P�֔R��H��o4D��@�k64$�Q�i��A�%>�d*�O�Qۃj� 9�X1��.�l�Y1�'I���'!>�p��ְ=���FJ�,s��	�����Y���Ѱ��b&F�US�m��?Ɋ}R���O,1�t�[�'I��;&�N�#2B9��J!D�X1�d��(F�(�!�ߩx�DXb1�~�ЌY�{��>�g}"hP��d��H��|X84
(\��?y�}R#<�g}bM#!�t�Y��6b��uYo����?�4��<��͵u�L��a�*3k��c���p���=9P/ӵ)φ�(@b@?�p`ɋi�<�Ceϫp�!F��3�@)�īc}��Ol��蟘��l��<M���-c��Za�ך�\}`Q�p?H>�c��O`�{��.��9ťՉE��}Z�"OT�v&�#&
�񄁒<^�L��"O�1#�nr(��z�CA3qy ���"O��p�M��;2��qbخqp- "O(�@��,=r�� ���T��I2"O��K�M�'	`�I �Ҥ}�4A$�':1O����ͭQ�TtPQs�L�%��Y�<��g�1C!.� )�V�@U^�B�	�?�fdj`N�d��|�����[����d��� ��Q��00���/&�� #��"D�tX�(�^v��T����,�A;D�(��o_1��9��K�tո���7D�|���q���	�m�5$´���4D���D(�VD���ՉW�=C��&�-D����Y9L��@{ԂA��ZĠd�-D��Y�+sF�Ր��k\Rx�í'��P�$?�'r�ͻ��!u��i���9��̓��?�v$-T5�����)d?ָ�C�S�<Q1�ɦI�b Iu��:uPĐ;�#�g؟���|��is����Q\�n�1CܘD{��	�A�
Y��X-+������r��}&PU}��E
X谁��2_�Ʊ��g�y� �L���!�a	��6�K�MO��ē�hO��je�HQ�m]Ҙ��ƍ�A� )�"O���ekȁ Rȥ��$�E+�D�t"O5jc�I4�b���l">!�D��.��$(5�o4��dG(�X��S�? t� ��Y�	�j��~��="w"O�4b��H�E�����Y�Ba3�"O<�j#"�47�a�� 9#���p�"O>����>v��E�3�I:(_T��搟����">�(�s������J<�B�	���#%
ҼC��Y���C䉢^9��rU�K L��f��V�=J>��y���><_�0�RiG�O����$���y�ESO����?^�z5�4
Ӌ�y"�J1zw�D(�.	[���P��
�y��.H��Y�aպM0A��'�y�lC�k�.)	�!�->�du�"�ބ�y��G�[�:Qi�C� 1�݀�jT��yRZ�8�E2%b=���k��.�y�D�1|�:�ԨF�A�C�(Q-�?�''�	'OO��M�c��gT��k�'����E��X�4Q0�N7�BIQ�'t�Ic�B`Tv��+��4]J�'���V�3q���P�η8a��'�NY� �*GX�!s%�|:,e��'��9�&Ƒ> �PD�j�
t�:�X�'Wjl��#�
-�B�l'�!�
�'�v$�4@�?� �1��o��S�'��A�1U�����E����N	�y�
ԧI¬��Z�E䴡Cv)��y�gR�
�^������@~�iUΞ�y2(�*1� �q�T�2���[�@��y�+�%�l}0!� +l�-"�E�%�yb�ғ2��UJ<1�@�����y�*K_46�cF�?&�|Ā3/��yR�܏P��)��"��9	���y2�,E��9:E�X�^X5Yg��yR�NW�u���̊	EB������y"�Ak/�O�)`Ƥ�Go@��y��@�*]��	��R�E�����y" +h^�L�+E7�T[�%�:�y2��B}��(!B�i��Ռ�ybϚ�'}:��'��Mom��b%�y��]���aO�J��t	�&	6�yB#I�lm2����3�������y�=\�jM���̯}�v�s�럲�y��@�Q�Ȑ#�!��`	!.��y�ɜDm�� bT$} bP�#���yR˒ �p!jT�yT&����J��yM��f��4ɒ>o+��Sh��yR�p�x�/7k�j0+��R:�yrA<C�b�I_�m�W��yҨM�,ʰ����/SB��x��F��y��ѻ*��@E�=6CP�wK	��y�.A8��Uk��)�~�(��ʏ�y���>��Q�A4Q>�L���ۻ�y"���w�L���,�8Qr��ƣ��yR ��N�ق��íC!jJ&.V�yB���3�d��#�� �q��o��yrB�*d(����)�VЩ)��ݱ�yr^�9�̼���\%��!c����O4qS+[�fÎ��a��r�D��7"OʍX��ɕ��}97F���xq�"O���i i�n@�@f�4�(��"O��@$n%(���5��"O0 ��F 0��h�sΜ�E����"O ��o³!m�u+��!#����"O��f� :p"��	�f�\���ɔ"O�pd��'M���ڣb��R��"O��X��җ��C]/b�D�A�"O� ������3L#8iq�k������"O��!C��9+lx˅	݂n��qP"O4��	Ԛ! �y����9�0h��"O.,�I�g�Lht��^��d@Q"Od�2��lR�p���L�L��U"Ot1X��D� `�@ìa�5c�"O��B��PP�a��ڀ�Έۄ"O<���O��Bր�5��/[�]K�"O�CUl�@������f%�J3"Ox��E�<�ŰC䆚7\�ڡ"Ot���J�}��f1L��b�&!�d�BP@Iz�Z�7���Qa��(J+!�џ+P�ɜO�E�'�����BU�a~��D5h��|3�I�'����g�+��<9$Ή &����G.�>QǍ�J�P�R4ܞ�y�w�<Yg�#gs�|�a*�4'�Vmb�r�	�hM��򔆖$f�(|E��M�^���qgj�2D�ԝY����ێ�0?9��[�IP����%�+�ܸ+�"�20_�q�4��O?�Ħ]?��'�Hk��қw#V��zE��'C��(A
A(U6(zI�v����c�I;72�����M�sq��Ȳ�?���3��N�,�ܨG�.~F���[�pc�������ĸZO�"��5���
�0<�F��{j>8��� �'P��J��Cx CSL���Z���	�2�E��B06��<�O��q��2�3���D��.G��Q���9"A��S�O��� �vO���7��F� "|��螟mR�w�("c��X�FM���Q&T2}��oӾ���	�"��O�h�H�#Ϙ����V�E��I"�Pc�$���On�p�!�!�i��!ʖ����C��1���g��H�����\�(!8�w� �ѤL�Z���ד�f<9##D���틏_� y���<<.�P���)ҦаeІ: ��SBH
���JY� aȣB�|���(���[ ����p�!�hO^,�ӍE�$����&�'{�,�C3���?��u�\7]������T�z�L G�/Z|�U녯�8[�@�׮�'xZ�&?��n�&{^��5���R#�E\"�Y��@��6-�[�lx�h˥4���C��ٚl
u���T!M�l��؈���5(%D��l׸p�:��n��o5Rl�ҢԹr�z�K��*����v�ɥ$$��ȓ��V���&!fvtҢ]>Op�!�!�o�@lQ�&f>���GW���6KE e�.v2lV�)Α٤�I�A!&<3��j�	���\Y�"A��� > �F�l9�Q �c}�)��(k���c�a>H�Q'0uѶ�q&�n=�UHFct�1#�-�~����9a��(���[ƾ0�3��}�'�*ȃ&:g����ZX��$����|ڀ���sk*�(u�щ2[8dp���p[G&ÊT-
�PS�Qo6 �~2q��p2�w�:]�s$��q�h�D��ruơ���:@�X����Ln� �\=�>YD��gP�w�,KQ�ŗ�v��j�=�x�A��2hHT)�)���3q.�"m����U�'���O|�D��.X5�Zd����k��4�O�-;��]E�u��5=
��]w�AQ�O�y��f�	K�ȈȢ I;$ \
�k	|K�t褍M	.	�"?)1AґY�\�;���Qު���մ� 4;Sa�6���[�Z�o�XEC��6>1c�?V߰��JԷ�6sӡ7��ӎO�@P��j�^�`��FP�#<�2���|�Pp�����x��ٍ)�9Χ&��$����5V
E�El�F�1B	�3^k�u;Aч\��h�kE�'���!	���1Q`���y���3H��裠o��)Q��� z�)��_80�Qq����3J�c>�'�1����&	^q��Ï<W7`�3@�PX8U0��&Y:��#Ń�?����%�hÖ$E�d�t`J`�T(�`�ơ�Cw^�J�-��V�ٲ��i�.P���I���9Pr�����7h���A
_��E�u�?fhe�B猹_V�؅*ۤ��O����J�6�fu`����������$�؈�JP	���a�܋?ܼ�;"O�*	���`́�؝�sm:��GC$�IGJvܹ�p.-��#<i��O��` 3
����C��]<2R���{���*c��cix۴��<�D��תګ6���{���L��p,z��n����J?���99 6���B.t���;�S�x��sbR�Z'���	?`)*�'��:%>��M|z�Ϗ�p��@���1���uJX!����l� P��ꀎ^���9�m�џx�&�_�U&�uQ��T'gm�PE#�5m��	�b_�D�FQ:v˃P>���ߘT �}A��Ԥ`o�P%c5m��5Z���K�`��WEҀt����"tij���N�q[*$N�P �=`ŀ$K������T��b� [�\|@�;/ɸTx5��S �!`� &E����,���H*d-1d��2q6�kҦ@>H�Q����k)tQ�k�1w<�1F=N��X��aU8��`n�?}H�иC�A>
�X}����ԓ�ď�;F�`*V�S���I$P�.���+�dlШ�>�dEiB=O�r��~���V�:��t!�+���� %�t9hу�l��-����bSvDY�c?m�-�`���T���㉫(�Ftsr�4�!�3��d����#FhAC���9�
P�A/�)�Dpc2!�0�����`��¯�	PZ��r��͘$f��q�ɚ�Z�B���'pi�&��+U.PEbێE�H3	O�@�x,�ubɼ@H���m �4��RԮ��Y&��[4$�D�ps�)���%	�AJ��T�گO��!��ҵ2�,����O\�KСO7Z�R����&noh92�ĺ �t��I�\B�[`��0`�C����S[�%��@:4 ���y��Z#^D�s0@±b�Ę'�� ���6鑑(} 4k�]�	�ԩ�u"�)i�1���@L���N\�_-����i�,z.([D$�
�ڵ�%�کj�(�8Š����e@�2��tH��'^I�˟�W�,8C +	GX�ģg��:vt�@3E��.v�Є�A�yn��Ǉ�4S�r���!H����FȻur�`c�.?)dݐd =xe��ۂ`��~�� ���
7a AA��{��tA�ғ�̈�" %�"�+rn�:~h�7���]}�H�M��$�h�!�F{��ŀe��!�6��6h@����Xt�Bn���SB�$V�@�f���#<)� P�5Ԑq���$L��;ЂʹF�+SmY1���b)ڤoB ��*_�0���i��]%��i��$�]�����7���Y�i�iI=����O~"mJ�N�TyY��'���*Т������qH��:�M�C���mK�J�@U1פO�"���j�NN
/ڨ���Ӓ9Ƃ��rkQ�l����۟D69�3��*����Z�=��Q�ɦ$=v��,h�ᨕoWd pRc֞��L�"��_�,���"0f�!��
�-i�帵�SUf tz��W	m�p����,3f��5"�>���m���O�l����������6m�t��#�Ħ�Tx���c�A����-;	@|r�˕�B���)��&{x��3����r���f�u�g��>�`@0l�+b��� ' |k,0����~o&(��.�Ō�
�N�
u��gfC�>�H�lФ'�����ڥ;U�X��FY�m�AR���,)M�Y�c%	�[c��6��.�٪Rd�>\�@�ef؀�~b#�?b�~Q��E���5#��p�`8���-nw�4 ��^�15f�J�+�x�����
 K��~��㑽fK�P���$F���ע�2~�BdM�L��p2��z'� ��"A�`G|�IN����1��	�$��`W�P2�� P(��tZ�8�'j�z�#O�����1��"�m����C@!s�̌j R�SN��C�N��~j�hG�)c$�=��Ԓo� �Ö�^�7��"�k���"Æ+FO�~n���ep�����eφ�Gٽ2Vv���L,.B�&lX�5r��K�eV>*���"bM��)�2OM4S��s��t��i�R!���׽oH�@�]� ]���!�e�^�&�48�kN4N>�[�M��0���ٰ$����H��È�2�d�zsHΝ
E�|��N�O:�s��*2����`���\��@�(%ή�j��?��|���L'M��:"��) |:U��On��|�T@��&Ȧ�r GR�=��x��m��K�ŨS� ����ՙ��L�i��n�&]B�M�zN���hM6�z�x�'߾A�L��R���@�e��1�#��%QP�J##�U�Z�����0�y2e��4=\|)U�Ԭ� 9���ű#\ ��Jqh�� ���!P=���s!����x���pl��p�#V0����A�
�贈"�(�&��rϓ?<+��H�!H?��A��{���1,��
sZxi�Oq��ۄoO�g=Td�s"�
f��yQ'�5�z-*�ʘ���T�'
Ш��h�`DD��	�@xJ�i (Z���zF D$+��erGW<	��[0"�6��S��"\�v���g�`Q��U"� ��vͳ ,A8)�A[��ğN�Y�'������n��S*�))|�뙻%u�x���?A����XV�����];X�y�#��d�/`� a����+Q匚;�L$����UW:�1��R�����E�2obI���͌�5V!�<K�xu1��6=n(��@��& �Ի�bϚ\�`�G0,�	�^R�3B-C�Ȯ<@P Hɼ�QK��"�:��#���}^�x�G��
#�	�^D�Q�S'Q�񮴱�N8t)�E��00~�4S�ǻ8N�|	ǌ����� ���¥��s�h��p��;�� б�ϐ-[�9{7�;����#�� 8����Θ�i2��q�h�>重9q̚y�1nC��Ѳk�{�¤�l��㫢Px|��JFK��n�vW��)�� �-��*6��j��[$]�	��
ΉT�p���C٭SE�m��n�#,���խ�9)>��$A%�zh����T�Ф��F�
|!�/@r�+q��L�84H���'�jp��$�8�N�\&��M�k�L��/܀6����#^�B��f��T��90a_�o�.�U���o�Z��CyB�~���`��@�ܰk���}����eC�	�	�͹A��-�7���~�ȉ�Yf���,@?}WxȒQ:��\҄B'C��S��ρy^���@�M7%J&l� ɽ�?�/O�$��i !����@�k�6x"��c˰a���9w,���B�Xf�O^`�HA8b2�E��"E0f_� ��oG��[�C[h H4&EIX��t���0g��!'S*:����+��j���Ϡ~z!Bɚ�\ΈqHpO��$�Wg��!N�X�2쀓O�Z�c�!X�*ְ�V�M�(���D�a��P��lK�X�rL��L�T�K�A�3	/ؐ��d.eȣh�V;��@OB�RCv� �&Q:�ܬ:�ۊS�8�)�Ć�d`�(L�?�����?Af&�=Ud��1e��@�v`cd�Nw�Z�Ň_j%[43L����gI�SPh�ё�2�MSpV���rc͏E���z���b���P���h�%At/�,Br��YV?	�1f�M�Uι<��]���ں(ֈ+B�_\L�{�OZ�����S�����a�f�3!��M�Hڼ�M������-F�k��p�2xQ�=!f�(�$���O m�4����MO��������MX&A����4鈲Q22�)���DԞQb4O�I�� [�cB�JT�i�0��{��PiҨO�W�\�O����đ�r�X��Չ˰NvQ�㯚�(I�ϟj�)�]�|����N<P7>#!e��L�E�>���k]J�=�Ȑ3��'���w���Z񥍉��t�4GR1E.�zQ+�.XԀ@@JK{45# $B.��O�T��<�0K�<S��vlМ ��Pb ]�P�+�� �h��!b��!���+ĽQ��Gx"�]��Hz��nu:��r	�(B%0��ŉ�%%d��&�R�(�Ĩb\w-puΓYc�ű$J��0��Ȁ���H�t��ul�q�Ԫ�(Xz���A�U�D�9q��9ړf�0�R�
����+��R+ ��ČJ>Yr�M)���.#�:]�� ͭ@ά�5�i$���ED֧
]��u(��y��ȣ2"���$�7�0��܉Y߸��0�V���'�:ܐ���>yE�L�t��v,r]۲K�Y���_wlhp�A�g�PY8e�O$#���O���0jJK�H�+ե����|͐�l�y�^�"H��}�Uď��jh
�k׿]�f)�4+�4^M򰈑�F%g�d�'?���wFP��GK�l�dt�u�_F�#0�E}��;z0�/ �3��ܵ@�Rq`Łخ7�=pf�ľ��}K��TW���
P�b�T�ӱ���b����g�ĒO����\�8��0��g� n��r�߶H�ɓS)����O�z��H�*��Y�D]>H�����Oݯ�$�QE �Y�\��Jl����q�#P ��0���(��r|b��O�sT�A(����]����>1���?,�P�!逝8��y��A�(n������ٺ@��b�{�/+����x�(߼W*H3# S{�Oy���!� �2���Ư�6�(��Y� pӨ��v|ܲ0+BEu�ŸQn�A�S�y� V�hˇ顥�ɀ�TX8&�U ��x�'j�r1A�a�g�I Lh�=JE/
�*��eCP���$S��4&_ S��Lْɘ����oݥ���ռ,U�l�O iRsO
�F �x�(��	��e1���U�Rt`�S��1����׼. ̰p�K�F��H%)M,$�D�ԙ#��D���
P���r��бM3F�)�>���� `�v�R�W�
���ɭL�^;���*?�9R& I�.��ɘ�X�\�b�F��Qv�R�� �2��M�����x��J�"�`QƋ�.DѰ�X����#�+CZ�@���"c6�5G��CT��tՋ�%K�-^��+�įG<@� ��<KW�t�bś�prN�j�#�	�p݃���w�^i�Ɲ$z��!�/�e��QS��@;�.R�����/��V龸%?㞀��@qC~����')n�@Ԋ��,<�0G�|2d���Y�F�~�Ӹ �j�+��>�1΋I�d	�l�7}�Ы�  R�\$B�.6�0Q��!ɽ��OJ�b��Q:^IҜJn�as��VH�c"�� ���f�¡	v'P�jb�,A�.�~2n18��d{�Đ��zew7�\��dŕ�<Hq��ڍ�lD���	�/JPP��fX�͘q�G�*TL���d�4��I�D�ڠeF��սC�p8�;��h�JAA��5��c����v���� :�	`UD��3fj<a Z��+�Ց9�̐��d�*�`l8�`8@ Z�>����,���PEݬHh�*�3H�,8�Ri�O���$�Ǣ�Z��qO��r`S'���@6�K4Gr8��Q��,o$�"�`ŰH{��>�8�-ւ0�@XB��}�Pd�a>73�̩�L�� ~X-�׏�6�0>�R��	YL� b& pH����증"qk�aI�pK�@+p�T܀u�ڨ���!�d� �2G[>u���?LL���������7lOF���"5}FĊ���%YnļZ�C�����B�I�h��L+:�,X�k�~$�$��'Zo�"~zu�ƲGf0|���V;����0��'~.�����p)ރ[_q�� a�-�<VҹC��!Q��	@�Od���c����d"�1�3ʓ?��Z�%"V���t�ʗ&:v���V�2����I���DH��-Jb�Z�c�U?6��/��M�>�A��+V��H�԰���'� �9�"ͮe�i*bd�\���4?�X��5�<HO�,h��q"xi��j�ۦU�'�IL�ԟ8��W`�&7L�qa��Y�N�p��'8}�u�	S(ݚ�ʠD�|`P�'��dt�x:p%P��(!�G&�)��R	��@˹BC��'��5�p����#��*f���q��P�~�R:`fX@��I:ȦHѢ"�}~�
Ou��{2T-y�� ����bپU����p�DٲW�O�r�;�]�"~Γ\]p��˛#`�\��Dǀ#`z<�ȓ,��)"D�V3h��k���)ޒ���R��MSWh�e���;	c�5��A�8�4邡ײgB�}��W�f@2�o��PД��DΕgծ�H�CJ��B�	�W�>���A(��T�A�+CZNB�I�
�ĻD�$��DK,�,��B�	;EV@�B�E�~ݻQ�`|�B�	f�*lSE�~t5��̽!
�B�	-X�Lݲ��R
d�$�r�ǔs�B�	�?�t,�m��/$	����(:X�C�ɱ5]n�q􉒐O���`�1/��C�5j�؁��U�����~��B�I1�xc¯�<��=��/�zB䉊=RQ��C�a@< 	-	�\B�6X��q�,٭q��T$ƀj�:B�ɷ6����p(�h���ș_�B�&κ8� �9!Q�I��C�;^�B�I�s����ưc���ׅ�qP�B��JV��7��#_�vaxG�=Q��B�	�9~��HV"ƺS�VѨ J�dO�C��%e��Ҳ�Z�?�]�Lӧd�C�	.:�M)0�@�VX����9w<PC�ɵL좥����{�i�ޙeRC�I�*�X9�e�E�&�����?&�DC�ɿ.�<��ˆ	c>���w�@_B�>w����`��*5�iy�(=/�C�	�!��uJ���_cбI ���شC�%�swIO��i)�A����C�	���9;��3\Ф�`�a�_�C�I=P�������M��)q�քzk�C�I�m�fq����<�X�BQ��1ۼB��+G�͸w-^�P����T$�}�B�\�G̔�*p�Hj��Ƅ+m�C�I�F�tuz6�в' ��4��[�dC�)� � ��4JGؽ� �7<V-�W"Ol�J�.A;��0"O�'S����"O�9�d�
�Scz�2EEP�#..(��"OD%dKPv�ʙ��ڧ��"OV��MΒ%����#	�`��"O �)�d��r"B	9Eaߟ�Ld��"O�����Q�=v<����.E�b3G"O@$�Ab��.�����Q��i��"O
ء���K�d�W	
�>���Y�"O�u�*T�|B"M�Ю1/����3"O⽰�Ã'<8%K=B�����"O�Y`P�����u%� M��`��"O����蝈9pn��S�A�е��"O����I�4-�pJ��͆"�n���"O|Q�0Æ�",���v�I�M���E"Ol}Q��ABpTsR�D9U�&|��"O~T*`P	h� 5��ʃ�u�j�3q�%���v�'���;�a�ڮ���mC	c<^���ت̊��	b>\�J�h5����
f�2p�G�q�Ĉ��5QB�ʂj߂&b����b[�T���&����G�7�J��f
H�O9��e*�� ���(����ر[������T��G�Z��dE�G�]�Q���K�U��+�N$B�|��(��=���+�`�>�ł�U�} %�Q0�Y�gnY(<q�D�|��dKB��o����� $d���ǋM� L�v�y�j~��5O�Z�y� ���4�S�L�8e�:Ór��%�(`��	�(P�?�C+��
�&'N2(j .L�:�~	!�Q?y�!Q�sg��>�O8I9����V��Zw�Jt{J@!���*�.N����l%*�4tF���AT���!�w%�!voP�%���+eGA>�j��AQئ	����t�џT�Ԥ߻!����A$8h�Fm�LF�#��
�Lj�cƒo��瓻 ���B��@�4v0Ѷ�KO�]��� R8�B����cHKĀa{N2��'�90b!�PS\сk	<W2~M"��<V*�%�����#�cפp�<�k���Sx�Q��P?zM��������K2�I�M�ws��c��='�ў̳f��Nh�}S����0H䰡oI<����Y8W��j�͙Y�e�p�V�_D��3.�.t�ք����	�x)�M~��)��~!�;c5Z�-�?|��Q�!�A_�8�lBG�Y��o�<)4V�!��%�f�(4�����YK�,]8D" ��RY�(�Q����0�ȱ#$ ã?Y.�Ō!��q+S�<�|c�HhU��,db�fkŴ
r0Ԓ�&�U@�4��fWo�Bl��'��|ze
+f`�KE4p6��<��@-nPN0Y�Qq�~t"Q�Ѳ9���F�DS��;���\���a����0h��j�#=8\��B;i�A
�I�H!Q�B7[�j�ql���4l�j�!4(Då�~�DJ���ئō?q)�HU.�e�'��M���K
����M�r.�hen��|���ڿ8���򄎶I-6�Cg�#Op����A**E�@�4B�rp����~��Ň}��h+�w(���<D��
��O�@���HD���[��#�/���` F,�E��� �7��A�R)�% �v��B�[���kV�*�TuB��9i&2���H�;`y�a��)�g�'n�0P0�D�JL���PLI276�	aӆ��D1HKд���031�y[w�!��ug	17;�1)SFL�$U�WoC�Y��JWf1E�>$x��&{�&(��+�2��1bda ��$�+j�1=�n�1Q�;Q�đ��׬f�\�#��3��3�e�\�l�R��3:�r�Q����Y�Љ�X?1y4�^'*��iD�X�$�H A �H> R�>H3B胣(ܱ:J���a��|�Ǎ�O�($q��7o�B}1��I�|{̴��Ðr�&E��o�2�� ��?y�m^�*m !�w�p�P^|,���i�<[vp��AJ�M�e��`S�{��ܛ�%ǧ�|�p$>擧�P���,R��Q�NԞp�a��)�	s$��R5)�6�H���^��p7bدT�ў��"͉��a���4FFͳ���*,ז���bU�)�$վ.���&i@�pgYm�q�F�h��`#�単j��I C�]�,�đA$n�VPΔ�V�Y1eџ�
Ƒ:xNqa�F[�ưi����+F��c��λm��������6����?U����OϚǴY�a�z���5�a�J2���� $ʙ0Y�pDxf�� ":ƃ�`4��hQI�Ɇ�=�D�k�v�Ba)]-Q��O�C
=�&h��Z{�&���$����)=H�)��O��S"�\sD��`�x�>�зC�D%>���GE<>"I�w��y1����S�^qF�rd��D2��X3!	���֊ъ!r�S`HP6���_�k��8GYp�'sB����zA��a�8ΰ��U�.�^���D�tH������DyC��a��9Ψ���#(�Q�p/�E�t �U��%|$��쑅��=���"3В� �H?_\�8cK�M�|��c�VĐ�P�T6�,4��j��<��%!�lH?X�A��&�R�Xç�v�T��jyj���X��$���(O�)��iq~��aP���"�(������^%7�a��,,���D��(lz�u"S�ѕ(�f�
Ѯ�,@G>����>��l�DR
f�e�P1	~ �u�+!/$�xfˑ���9@@FZ-ЕJ"��c� y�o�q�s��z�*O@Q�����������jT޶�Q��+	(�ǓQ���#����	{��rעT(�X��λ$Sv5�G�.p%\=��a��P���+�%�1
s��
��+�H娎x�? B�r��J9\��y#�ʂ�O;N���Ĩ�p=��KS�W���C����ž���O.�$jU��:��;��ʺg��r�a��S�h�3�<ľ���Ǝ-����8��+�
��"�C��ֽ�t��NÃ7ր�GxҦZv�i`W�/}.N�(W휄d�51a\s�����ת�<�&�;r�p�8����.Ub�␉�џ�ϓr�����%�+
�6 ��5��Ѡh�D���/h��D��3w1�FN�Ww`���	7F��!3�c�#o�\�Y��.k�P3t,2t4�&NόQE&�*a�αOԍ�ҺHE	�"�@����uq�",OLT"���AH�� ԅ4�������G�"!��x�VJ�Oz����c2jω�n�0���_�#"�mȵh�b�`5*�Y�^ɻ3�P��{B�ս8{l0XEI7m6ޜXl 7d`p�o�J���+Ճ	t�tK���C�p�D��W9θ�쀵aP(tO�O���k��Lq��m	GgǶTC�U�2+��<�2hi��d�/�R����Oi��Hゅ�Lq&M�r�T�(���vkK@"��r"�_�P56u��	 (m��xA��߯#(�3u��~����k
E)��"���8R6�I�{�d��"�A�+a�!�"Ķ!�����Ǝ.�T���V%Lt#b-\��tԀ�. 4-j�qe��5'��%��ʆ/S
�`��u��1 0,�VI����H3���A�k_� �H�A�d�n�'��zW�C�j؎��"ʸe��!�j�ro.��VY;[!��3֋F��$*�F��iڊ��bJ�g��!��� t ���jϱ-��a�5#Tɾ�Qc�J�a������*e����1�4Pe�!r�T�"�'pz`X�1��Sr"W*!�Ne*��2TuG៬J��U�vwvpّ�9rB��Ѕ����i�ף�,yE{��2`	2Mߴ|�P)�%�MS��Yq+�lٚi��"GA��Q���3C��V-�5)(xtQe4;��IiЊM���D��i �C1�~b/A�=�bp(!�L$�	P��@��?�L�>��$܁&"D���;�vTx�O�H#�- ��s�$���1�L�X5H2B�F���[i�~$k���V�� k��׬e�V�r�'=~���PZ~-��ِ
�m�Q���-���s%%V��?1A�X�5n%�bM�TRlR��y�6��Y����Q	�(���E�˲;���H�oF>������'��`�o<��$r�I���L!����9l�ڡ�f��a�4ˑU0K�܅���jhH
FɁ��@!ۤj:i�Խ�f c�|8���b��T ��%r>�q1"�#ғ)4�Q��3\i>���n��0�b��3��P�c�GP��j��6��AP�&ɶ<ur�h5`N�B8V�ks꜇`�D�#�G�R	��BTĻ2��u8�'� ����Y�������L���q)���U�p(�/ʰ�tQ	�0�p)ن
�����`MN���1����Г�ԾQ�yK�	�Z$ ���I��8�Xͳae�5`�V���"��O���Dz��ǜd��Tj� �H���D(V�Rq��ᆈO��bU�M�T�"��t���$���&�L��tM�)U�LM�a�4:yi�ʂ�7%~%��@J���$�M[R����*
VԀ��l
�(���jeD��KV�U�T�Y��"�H%�˹xb��*d�f?����)QR��S#��"�*MR�O>N��N'�����R���ajs
? �-X�,	�5^���'�(�(�2'_�l��B�p�ΰ�r�C
d�"%k$�mj��ǻb<���F�p�CcԚf?d�k����v!��(g�l�j����v�d��d�R�c����t��U�G��0�,��"� 0 _�mǉY�x�(�!���(�0#��r��q�'*@��&���O4���,��H���F�Fb ��D[�\�1�la��;T� (�X��5H���O��Yc&�M�4B�I�X̓�n� Gl �I%H$���(D��b%4V���WR �$����B&P�;E�$�2'J(/��[f�.`�b0�$(q�� yP�TT��s쓁_���HT@��8$�1煋��A"��T�h0�*Ot(C'H�,X����z�I����5y����b�I��0P�Ɓs�� ��C:�B�a�U�bX�0�a�"N��TLPC����p0+p���g,�*��4��� �T�M�Y��&MCv,9ЬZ�drZq� ě�k�ǁɨ�`���%J�q���F|
0�,gzH���a�����@maN4�s+�7t�Q��9Ks���fŐ=��d�GǛd���ӄ瀚ndT�=>�#T�O���)U�6*�-��g�c��Dk� �W�Q���Nt�HO5�c�V�O7��-G&�������C��ǳQ��+��	z�PeD�Ġ8_���^ػF*��,���yލ�7I^�g�h#G�O�0��3�:{��y�!�N6s%�'��m���ϴv)�Y#��%7d��g	ߊ��Ѡ���"|��D�d��/D���'1�S'G
�f|dB���]�`�I�Q�py�lGW�B�@��o]^�*5$ͧft�i%kK���	� m4)����)\R�0Ĥ �+#\�rR�R�9�Ƭ��EQGGx��g�C����c�S�5gJŢ$(aw�A�i�-=�$�#��U�N���z���B����:7cLͺt�*d|�$)����5�@%uj�7f���A��V�~�1#�� U�|L��=?�|�
ƞ7�D!���?����P�n�A�K�"b�$��W:�p!d <K��� �F�1�L�(CFd�ӄ�K&h��H>٤�K�$C�}�n��p�Hec�-�#��j�6s�rB�մrӔ�i���,F�v�܎B�̩��N0?F\�]	�C!ŠAD封�ȱ]�,4�1G�J8�U����<�dU�� ���Y�kŰ�@M[w��
�	�+�F7�ݒ�#��v�@7-\" p���ƽ_:j��FN�*�]AҢ�-�~���G�m중��$���q��JR&IJ>@�v�'}"�$M��l�r����X�a :JV]�	�G�D�[�ԅ.C��yz1�-[R��p���B[�r�ڤLp��5%���'Af̚�w� 1p��*�4U����A2���ጓ �u��S�
G��`䓩��O�l*7O���q�Q�<��l�V#�(X��E�K����k �,r1��e�Ə!������G�s;F��+L�[2��SQ�HFt��#��x�U����z������ �'dݰ�;_k45�j��/�`����JȢ����ͳ}��4��Mר/	�}��l�H�'!��[�l�!;��
ߐzpx�(���&J�HZ2JF>z��!����0��e���a�D��g/Y=%��؀AƗ�H��Ĥ�}��Iĳ^��sh�~WF��g*����O���4����VP��ď";��uY1�(N�<����pC#�y�j��O]8�f�Q䚟��Q-߻s56�x�H�o�Q?1�6a��txq�O�3Z��ZekR"m�Q#!R����.V�.-�F�ݶ�O� �]�)�Qê�=o��)���о)�&1��`�����C������L>�7E�1c��1�F�8�.ESDC�}[�=K6O��:h*�����C�&̭;tņ�Cfl���tǬ�B�I�/bZxS%��VDB����U��2��!�T��P0��s��:U� :U��-��m|�RƋ�=���&���R �6G.c�6��{2#1Z���O��{�ß>���c�J߻g��ձ���Y�~r�E1FN�z�bd*B�ĩ~况��G[e���s�.Pl�EZ%�+o�!
lW�!V��[$nX/z�?!@�A?0|Ȁ�k�d�����GWV�[�;N�,A�k�-�` ž2~�O�x�5Q~���4B>D$m���C���L;������e$lB��L>��X9F-
��ό6���[GMBD�֬� ��݀�ڏxm��!T�d�;���g1豥O�L#6N��\Xe�W�U+V�*xs�l�&`6���a�7|1\�j����mH�M�\�UY'k +���g�:,��yU@Y�>(���ͼr��}��"X�V4�x���ògD�4�fH봟��s��1:�ܓ�烒d}�M�"	;�	�[,ukL�h`���'������w���4��X�`�D�b틤:o�ɂ8%�c	�*���Y�@�j�O|�tH�"2�,���k�c�$���W9B�N0�C9{����B�-z�D����y��"\����S��-q�[�[��,� H�x�������E��h�Q�3�I%v
eU�B4y9c� /��\�Q'P1S�^�S0�t�BΩ?�"�ʀ����&�n�i��ރ9� ]�M��zY�Aʐ#M��	�#oS�D>ڈو��G)B�<�w`O�b��&HT!"��b�F'Wl�@��`�N���tjryz�'��*ѓig�+��7w�)
�b����\�*��a�wJ��}gQ����K�h��=��|���&��"��F�N�E�2�r-�	��p"J�Y?��	X�oS�|P5�RU��X���鑹M#���� ��H�����ɟ-,3�ޫQ[n�2�.R��h��" ��7��}��~mZ�i�Wf�@0!c�Z�3����E$�n0��%��DI!W5l���ޒz*D�K�N�2ŃW3x�	����?�$�S�	H���X&v�ʨ�j��0��)�F�C�M27���O�>!�^f�Q�`G�;E,��򲍂&7�h�oZ��h(([U�q�Ƙm?� ��8C)���mæ��)<}����R.y�Ҍ3�⚌�a{�rnNl�`R}��� ���y?r���iЁA ���%hM�����L�:a'ϮCotM��i�/��	��f{d��&�?qK�O���O]l����D]�PÞ�>�Q��5y���c�/�	3ʸr�@E1��P�/O$�0�j�����x��}h��K�ph���L�D��笞���XX&��^���d�z��y¯C��`�N�8�Esd���k���IA��g�T���eк���bҵVO�	ї�>g��7-�7V�Rl�v�H�%�|���2}��ԑcI���O*����:�2���M	�hxa��'�"��0��r�:�*�N״jc�Yy���m�
��'�<�rE�ēze*A�g`	�O$ҵ�Fj-7�f,�?����G��H��o��%�Jb?U �D�W�P�vk�;���t  D�dC@�.{EL�i4擭mڲ��6�h��d��D`:ݖ����*�>l�� �#>��xk�m�'1|!��ݪi��m�	�T��M�%F��d[&o@�Dx�jG4�0=�.	+jF�"�ˈAQ��a�T\x��A��^�vCƱp�h$�Î��^���ҿ�y�J�{�p�0�,p�J����yBB�=sݡ��k�Z��\�yro3S�`
��(`�$=�P)��y�ʚ�l�nQ�U��:X&��W�:�y�䑜]f��k��E�xa�W��y���ъ��S�3<W��cf*P��y��o�{� �,�B=�5IΛ�y���&�Jm�CΜ .A�5�T��#�y�%5y�����`��+qD�RD*�yr�SIŴ\���m["kU0Q�	�'렍�F�S��Rl{�&w�9��'_�T)�`Y %��x��G��4[�'a&�qƯk6���@`ZŃ�'�|=CQ�`'d�['@Y�>�X�':e�í�sG� 5g&J؅8�'L�!��M�D[��DB_�SX���'7�I�B��/R)��J�J�+j����'x0��O,"���`Dh <���'1t�rB�eRZ���������'st��Ǩǟ���㗧\���x	�'8�
3!�:���P�
 ;/�(��'0"%
5 �V�L�{0)�#k��I�'��y2�M-D�1�F�� �n���'�1)��M$R�,��ՈD���(��'�
au�ʽj�#Y��<4ʞ'�^�I�N(a0��P�.� k�]h����(c�찡"�>��cg��1��ɍHQ�"}� 0M��!� +�p�;�(��P5��9�i0�Gy��)��y�� ��\�S�楋ŇM+� �<�"�O�X�]���%9tȽ4]�T��O��Cb�VP�S�Oh��9��%M5��tm�$3 �<bش=ƶ�����a�S�OH>�j�I�"�|�Q���.jbԀ��(v��b�Ј��-�����'_کI��οq԰���fA'"XJ|����Z~ōNE�"n�^
D��c��+Î�#���H�T�C�\�f�\�`D�@�H�Rw� �e����ED����8��i�,�����O�?M`	ڡH,�a{!��Aa�4 ��b��"��LL>��bO�xd�b��(T�@���۟�h�|�&��J�T$���:v&(YѬ֊�@�&�,Q���0|B��[�b��]�$�NV|1�C�|�	6'�"��x�韮�j�O"�	�[�#GV�9Ɂ(�L8:�^�1�����اH��([�&�M���
��Ht�d���'iD�d��S*e�!x�1��|Rt�ѿ|�h �B�_��'5��V\��i�G���ϓ6"m�PCXR��;��E�"I;q��4�-OIo�I>��	b��1�nX�!�c���(��0�M�s�-�)�S9>h��Ċ�.�����	�T�Fʓ+;�v��_�S�O���Q��.�<�р�7���Z����6#�G�Ӻ#���/%�j��*����u���֍A(��Z�V���'�a����8�N<�`(��m4U�oӷ{ZI�#Ȅ��R<M�p����$O��
�l	ho���º�TT�	��č���ڕ�Z`>Aa�`K�|�i��ʶ3:,9��L���r�7O�h3�������)�mؚi�iO�9F�M�R	�7d!�C�.�P��	��L�ŷ ��"O�	�VG�&q�r��)Oojܰ"O�9 �'��3e�ۖ[J*�z#"O��F�����j��Q2Z8�Q�"O�@f�N�R�"(��l���iJ"OJtAs�A�%���Cҋ�9qA&"O�@؇�!;\%�qL>����"O���M^�>��U,,h����"OFP�$�Y�d+&|v���my*Ab�"OU	f��1*�.���8j��"OJ}rr��R����<Eb�sT"OJ��������xQ(:+G8 �"OV���V�g 4��f�$�X�"O�`
���"�\Ih�N@%\��ؙS"O�$�Ɉ��
��W�{�M�"O
*`$B�/ V�E�*�`�"O�A`BD�p�m��lV&}��d	"O���f���?F�`j�Kv܍�`"O�{���L�z���(�p�d�H�"O.��AJ�s+rtjAh��&�&�3V"O����"�@�f�9���0"OT�P1�==�4���I��#�"O(@!]�;F.q�v@W0���"O�Q��`�^`�Tғn�E�E
7"O�$��T���h�uM�6T3ٲ"O,Ԓ�S�F$Y�0퍦e���(�"O�,z�%�=�B=r�F׽K�t1:W"O.����iXĀ�U�O�d���"O.i1d�V��q��n[�"m�0i$"O�y(��	(����D�5[l�`�"O��dANb,q���Z�/����B"O�a
�MǡI�b�S0��5���"O�@	!I�.a�ؑ���
���"O�`�b=�x��W(�tn��4"Of��a�ьt�Ј��Y�^0qc"O�%A�
Ą �0���W�d�ft:�"O-s�`'#h	���"����#"O2)0��1�ll���F�?�j$@�"O�ڧdD���HPc�Kq^0{�"O�3�"
KܽHT!�6��]�"O� Dъ���v �jR*�"+t�$*u"Ovl:g�W+.G�C"i��~x2=�"O��Z L�c4��ʂ4C�ՠ�"Oĕ��iȅ+����Q�.Q�@��"Oڥ�5+T.oL^q�>2<9q�"OZ�2��=46��2�h�%J�S"OV�YU���7<�Y���"jV�3G"Od�*��ŰH@yѲ���W���rv"O��C!䝐Sk�I15��5�J�
�"Ot��U�ڔ}e:�p4���y��lAs"O�$��ᓈw lS���$��Pa�*O��0�� �41�Dǖqm��
�'_�Dr��y[��r "x`H�j
�'E���Lq�pQy�%ێX4�=
�'<�p��T�3`�qQ��&X��Dh	�'�x\�C��w��]��QZ�l	�'�r�)Rꐖ:���A@C�$��'����5��,0��z�"z	q�'����D�EU4�c	�ƅ"�'} ��0�Ԭ)���R $X}�����'�L�����B�D9
�	]0
�l9�'�P�Jn���1�7LL-Nt���
�'%
U#�'�)O�JE�G�
�G�H�
�'G�q�QG
��>lC�m�(�:;
�'�@���T�<��8��G�*S�p��
�'^�𲌀
�L��o���
�'�n�bwhG�c�v)	�nX|D���'F�!�m���� U�p��d*�'@�T�%.����o�XaR5:	�'�y���X��s®W�k�1r�')�虱柉8�8qb)u�L4��'� �(���+�x�X�,R�e�eJ�'@����;	,d9 �h��]�~DC	�'%4
1�j��q��Mp����'(6��	������a�A,���']�a{RKU�)�A:@�\<�
�'�H�Y��V9|���av�9�$0[�'�T�+�i�+����E�F31�9�	�'?v$(��2f1T)0D}|}(�'�Ɓ��jY�����C�K��r�'w\��.�#�F�%J-9�R���'�hx3"A�*~��D��	��e��'u���P�?v<��$m�%/#�� �'��噐,�b4$��
֯'zl1:�'V�PqǑ}(-1QC�3C�H�'�9k���UVNH�ǖ�~`��'y�ر�)��G� �S�'Pp--2�'��}�1�W�\AfM���P��'Z����[�N��u fhπȈ��'�Z)81�E�K�y���,�~��'�ޙI��n`��$��&_0��
�'��]����r7���C�YvТtb	�'TyR��(g4�asK��[��h	�'* ��g�<��@�"�N����'��2E�<4�n�#2�̚]vPpZ�'�zrm�6O�� ��L360:�'$fAJB�N	ƍ�eM�L(����'L@÷ǟdv|��)�)I�~�Z�'�n��&���P��A�0"�&L~4)Q�'�ظsTg�
%~čQ��Az���X�'�R�CD��_a�A�qi\'o0}9�'�N�&�F@(��b� bP��'=X q.3*1�P�`�F*{��h�ȓD����"<>��@�W�{�L̆�S�? ��aD�.�x�"F�!E�$�d"O�`��A��+#��Stl�JЬy��"Ofm!Q�B��j)�QM � �I�e"O��9�C��y8T��T����lP95"O(	0f��(gRٰu�G�X�*q�"O��[�όa����V:u�^���"O�MP��� ��l#�@	4�7"O4˰� ^C($��� ���*�"O��a�A��Gj�8a�SIt�W"O�4�������M�Dyh89�ς��yr��+�T�Y$7�� MI��yr�I/�f�� L[8+��9Ǣ ��y⎙�n�0�@�-z8N�9fJ��yB��?(�6���w@$P�G���y�L�� qB��ɪ�MD
Ĕ�yb�^�l����9 N�{ܚ��yR���x;��+�J��VBQ���y����3�>���h԰�ii��1�y�J�F�B��m�0P�ԟ�y2�A�(�~��rb��c�\�6��?�y��F�v�B��`��
x���X*�y��*x}y�J�6�U��%��y���R�Ȁ��D�WA]C��	=�yr	S�Q�0���8`ap�"�y2��8U�@1Q��
X�r�c����y�S
+r�P#�9P�zu�!GN;�y��@�x��pc�	����0Q!��y�Ooɐ��� �3R��!��L7D�\2`�5Y����ԽjL��'!D��3+2Sl�s R�m��!�R�#D�`�@ >ty$p��G-^JD%��6D�4a$*/I-�5����D�Y�4D�\4�R23#�M��b�>l(q�A6D��i��2j���j���2

�$ uF5D�رta0am&��R�3�R����.D��s�Z�A�>e*5�&o]z�)��-D� ���.+A�Q*c��M�d�c!,D�p�QDT�D���� �Qv2%�5D�Tz�i�%8��rv.� ��z5o3D�$�r��9wt�t+&��D�"���/D��UL��G$�9hpE�r�\���!D��sgd��z�~8ӥ�Z�'�+D�,q&ЕyS�9� -E	#b
�;��'D�t�тXa�q! %E)�,���%D���Aԛ3U�8`Vφ/qL( b5%"D�p��Bֆ�b�B0&���0|��o>D�8#��W�V���CV�ߊ:�(CW�&D���
[�}��'�h$��E"D��iEB@�j�B��� @6<���d(.D��#rk^�#������� �1�L8D��:��H{��i�k�� ,����*8D�DRRg�l���e�ȔH��dHB�5D�,C��פgKNH#���}���0��>D��{J���Qel�4x�\��2D��r&�9hv�
��_��R�g2D�L��]��m��d�	����sI>D����D���Υ!J�m�{ф:D�P���\�/nx��P8 P�:D���B�# z� g/N
W.Q��l#D�ze%	.0*uk� ���A�%D��Q�/P�͊ԫ�KGK;0}q�,(D�聅� �3�\����_
z��� ` D�lS�n\�:H��o �M�e*OD�i�U�q��t.��[��u�q"O� $����Ql�a�o�-���@5"O�=C�G]�[�؁�ˀ&�Fp�"O�ܒ�щ3�~�R�J�%~��Q�"O��ڲe�z ��`���'m�l�Hu"O����E!GL<��h�&}�� &"O� ��ӣ&x�!q��(�
�2�"On�k�CK(�9٢'�[�hr�"O
Yb�鑯�ඦ�({т�x�"O�59�Hp�M{a,��7��0*O��q�I	=KΔ$����$x��p�'�B$����4��p�R��4x��'\�*R�K�|�H膪0J�6H�'�`�!�A�_B~}p�A�4-�>���'�����~�<�W��,	����'om�A��m(�[qM�>r��)�'�V���!�|�X@mcl@5�
�'Z^��BM�l	S���`eְ�
�'j:p� ����X��؊[�J��	�'�Byq0b��q� �ri�^T�DS�'�2y	��Z�(�6��#���T�|u��'�EjǦRw3���o05y�'-�th��	��`�H�&��8x�'(vL"�"հR�����ƀVe�̘�'�EHPo��%lN!ᇇ�U$�l��'�b���(H�n�8#r��'@�h �'׼���k�5�8<82��*����'䖸������&�c�gG�{Ҋ�
�'��]��N��h���HmZ�9�'�2��  ���   �  �  P  �  �*  �5  �>  �J  �T  .[  �a  �g  n  \t  �z  �  $�  g�  ��  �  2�  r�  ��  ��  9�  ¿  k�  ��  )�  ��  ��  ?�  ��  =�  	�  M � _	  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r{�EQ�( �gVlɦ�M,H"�OQ��Ʀa��#%$�$y\&�+��'�ўl�Q�v�*ax1�:0n腓A�1D��{tCO.]�)X��$\�L��k0D��s� ]!B$�%#��سt
2D��� ʓ+(�)�`!Tft��%/D���n��~���(�ڍbd�0D��aBK�>/(��sD<U"bX�!#/D�8�P㓎U�؜ʠa�IVD�w�?Op�=Y5
B����G�i�t���A�{�<����O���)�L��Ii��c��<�g�'L�O?9AD]�K�DE3R���`��c��=D�ң-
v��Ѩ�&�����<I�  L�3AJ"OF�u`GF�u�����#�|%�j�U}���%Me�Q�ȓ'�i��Ӝv�^�CE�Ŋ^2���ȓ�މ+��*�A�SǇR��-�ȓgV.�a�\�Y��S쓃7㎄����aJt�d��t�Q�+	]����2z�l��Q6��
�)b�Ć�`ob5cJ����p�B"S�2�0��ȓ8��|ӑ��lr��� ئ|���&~L�
EMٿFp��j%�� ��ȓQ�v���GAu{�f�V�u�ȓ!7�s(�"X�@���ɑ@$D�ȓ%h%
g�e,8�chH
ن�S�? �H$�X�/�XI�Ɓ�e�qC�"O���LؾVs��)w�<D�r(�W"O��-�N��a��$B�t�rP8�"O@��C��#�t8�"݊]�\l�W"O6��ʊ����<O,Nt��$ON�!����?��"ׯ 	{ʩe��-B���hO���� �'� M��r�,�z"O�dc�!2h��π,dD!�"O� �W"�V��{Q#8S0,@g"Ol([!��!��I(E�p$؂t"O$D� e	*��;4���5P�| �����E���}7l�0)�����	["�yf�31 �kF%h\i��F��yr�\�T�$�B��V%����M��yR�;Z����f
:'�	H�����'��zb %b�r�Z`�Y�&�LmSj�	�y���-���J��$��se:�y����2��1E��r�t1`�#�􉵙��hO�Z7L�m����!C��9fO�J`�~"]���Q�s#��c�Y{����'8T"=E��4M+ �w�K�n'���� Sg��I�� ��1ғ�� 6��L	1�G���̆ȓB� I�Bh��ǐ�Ih8��'ў�|�ש��/���"��'`��H4�I~�<� ��7��a�f$�%
5�u�b�<��H����I� �6�bDyf^x�tQ�ҁ�'f�p�ɉ	Jd�d���N����/�S�O�0�iP�JE�(��ˊ�_=�4���D7�G��D�d�����G�ӵ<�5�<�	�o�r�!��?r ��p��:x����ȓv��qp撊U��YЀ´+-����a���2�@0#~4��B1k6�}�ȓB�	6�!�8�rjQ-#�d�ȓEbp�J��
1���٣�Yq �ȓ�R9��%˟P�$�y�>r�d!���T:�H5�p\�㌆�\r�I�ȓA�L{��N4#Ĉ0���75/�E��t�ƭ�4���;�@)xa���uAt���(3dtrB��2RȤ�G���i�,��2��,�UÀ���Z'|{�	��tޢ����
xzeQ�aW��H��?9ӓG=fA�c��4^��B���p =����?���I�p����g,�;Z(���h�<�b��5B�֩���16�R��'ў�?-lZ�$�Ȕ�lğP�y�JA5,fB䉘>h���I�1d�X�%@70P�=Y�'RZ0���b@R�N�zv����>ه�� k�$��r�-�#�A6]�q��p}*��t�S��{b���MZ��`���'���B�$�y�!�x
l���8Jp�j֥�
��d�ӟ$��MȾ�óh��Rc�҂'k�2T�2��y���ghN�z��e�ƹl=&��q��l@CEe�<I6��@uމ�4%I�T���`Ci�hX�4Ey�'���<u�Eɘ�n��ĺ����y�)f�@}���L��N"�t�/O�ʓ��S�O��i1� T�n��ĨL�vp����y�F��m�p�a��!:*��$���'�����gܓ@�|�$Nι/+T$�`92��D���r>%
�m�%}�UA#KH*t=�ԡ D��c�倏lͦ�P���(�$��":��҈�����Kܫm\�-[�œ�L����S"O"�+��X�d����j;[�̌�"O��(d���� *��hP��'��	�9�+�͙�~qu���.��#=��S�? ��@\?F���g�< t���t"W���)����F�M����w^�}V�_��
�0?�0	��g��)h`Rk|Z�CoSݟpG{��Ƀ�3�Z����'B��q:��C�I�Zi�Fb��
����g��<q�B䉬V�@����Ƈ�v�Ѕ��}?���hO�>=��
1: �*�)BA��!r��O����S��{��D7(�Ni%�8/���dς��$(�d�A�Oh�4����k� x�!��0Nɨ�3�'Z�	ӅdQZ�){��/��-:d��$]jb�)�'���3��v	��sA�J�l���cyrS�8�C�X�(�|�8���n瞴FO+D����iu��Q��@��$���)ꓬȟ.�e�$O6 �y�E�+:��B"Ot-�uĈ�����`x�E�-~_�n������ē��>q`@A�A������6~0����XR�<Հ\�	�:�A�A�A�0�t�
L?�!$�S�O.��& i�48�!���@m��'�N�;SC�+q�@	(eb�� ���!�'�T�Z�*'�����]	J��pJ>����I�H�1wi�P��|� ��_�!�D���i���l�hi�Vjζf�Q�`��
,�<PR3���D�5��Q�!�B��2�>��Eϓ(_�ya,�#IPC䉀C���r�e������� 9C�	>3���۵��M܄�rc��B�	1x�,���K/RÜ����@�B�	�q����&o<z̘6HO/��B�ɀ'��k���](�2���8dC�I�#�B��b\�Rͨ�����+L��B�I�6A>u�w�M�ca�0�]��C�ɑ�xh��P���a�kߎC�I8/x� ��[�*Ö�2D gB�I8" *s� n%��{#�b�*C䉎
��YH�

�Ka2�o�w��B�	/Z`�1��%2��Y�[�x�B��
����eJ��@�X�h+�C�%x$�8ԏ�f���c�W<g B�I�]��	_26ܒ3�2l∊�"O1+���($��
�	��&��"O�%��lڦN'=�&C,ƘmR�"O�m*%L0 M��E�N��M��"O�]��`#��a�#�>8��$�"O�D�@&o'�@����^���"O&�����}�$�B�D1A���(5"O��a����I;A��(�xX�w"OZRg�H�G0���@�:�L9:�"O�8�a	 ���� �9M}��&"O �c@+�<^����1.
��"O����8�Ā�� �sq�Q�R"O=�d���e ¢$(�a�0"O���3C§G0�x�'�\ WQ1�"O�a�!�<*�xB@�U+Z�L)�"O���A�C' d(�g�x�-�V"O�����qN�)�f �L���!�$^�q��}���hR� � �p�!��=��⢄ՄSC��A�p�!��A'>�X�y�k�-%�Ce �v�!�J��U�LR��Y����!�:c`њg��3�ht�c�h�!�$2��LSBk�6D�>�9�k�!�Ų%F��8V(��=���Z �L5Wv!�+E6��f�1�$-HӨ�!�ƫy�h�x�K����\I�ȸ~�!�� ~d)�!�>^������q��"O��4�Z'i���X�)K�$��Ӱ"O<��B(׵���)D/TE�����"O��Q�р5�� ۢm�:���"Oh]p�#ձ~��as�Ф+ư#��'<��'���'���'���'���'s��qԁH�r�V��TOS!fI|P��'|"�'���'�r�'�r�'B�'=�5�g�[C&�p���2sW9��'���'���'�r�'kR�'��'�t�`aJ��t���7Z�t����'}2�'���'���'���'���'q�#aM�+��Q@��@�r��8�f�'T�'nr�'���'���'���'<0�%��11. M�P�q�wn�:�?A���?A��?����?���?���?qeǻ�6ęw�M}p�0�w��6�?Q��?����?Q���?Y���?i��?��Ɵ
P�5F"(!��[�A�7�?	��?���?y��?i��?I��?I�J�I�V�0!�W�+��(3�[�?a���?a��?Y���?����?y��?3kP3}��T[lE�V�R\E���?)��?����?Q��?����?A���?Y�/ޒ?��kuE�HӀ�-I�l��	П@���p�	����柜��ğ����j����VҌ�hw��L����I��$��ʟ4�I�����������ɻ����$(�@@I`F��p�4��֟t��ʟ���x��ǟ�C�4�?a��L�-�!�@�;>�Sg�:�vd�P�p��Qy���Of�o��<��Q�E��3s��h�%Y�s��Y��<?���i�O�9O,�m�)Ny�,�#i�p�b��#�[:P�|���4�?�T�C�M��Oh��P:SI��I?�3ԃL�M����j�#��U/$�ԟ��'��>)�#���vt����!��rF��M����@̓��O�R7=�D(�.�M�&���Ç�)ސ��aĦ�	�4�yP�b>Y�!�Φ��G�k_�P3�yԥN:RH0̓;��(ɖc��D[H�+��4�����9U�U���<L������<�J>q��i��mP�y"&V 1�z�;��N7����;uc�OV��'{x7-Kݦm����Q��hX�UH�`��nàA>�	%`a�aV�BҪc>�0sa�к���'Y��lNf�.��"�` �p�Q�x�'	��9Oz�С!`�ǡS���5�H�y"Ct�Xt�G���!ڴ����ď�E��=�G䈟O,j���[��y�#|�mZΟP෨C馁�'j%�g�ڹ��eYt퇭w�:U'K](����2��+C@��kn0�b@@���C�˵8(L���b 5
x����&������64&Ф6Ȕ�s޴�aO�
��H���0?�#Jy�
!s���WZ!$H�08�� ��I�Oͦ����RL��\#ë�i�L�[��L�CrT�a�J�>$��� c�U���T��,x&�"w!�����W+{����.|j�`��X�.\(e֏�&Pv1b�#���Uc�&]���p	&�XKT"�<>e2DO >�Z�[�T��U���(�I�?}�ş�Ʉ֢i�lP����.&(�h�������O$���*�O"�D�<�'��S�|/tPsv��H�~`IW�Չ(�z7M^�9�"n����	���S�?��t��Y���eCǲ&��A@�:80��4�P���?�(O�I9�i�O��p�
�+�]a�
q<$��dAউ�	������8��ܴ�?Q��?����?�;_���&��a���s���74N=lߟ�'F`����i�O�d�?���l'@!�����k��\��M��RS� V�i���'�B�'Ԫ�'�~���B9BS��`k�(Nؚ�M��섗E�pqΓ�?I��"���?A��?A����]!Bl��X�,Ir�
+F1�M���iEB�'d��'�6����O&Ѳ�"�81��J��G�-V`!(P��O��d�OZ���O��'3��(�v�i����,�!���b�ͼS��YUo�t���O����O����<1�~&�Y�'a�^��Q�A,=S�U�CeM/%X\!�DU���؟�	����'Bh�U�ڴ�?������+V�45�������x@@�i7��'B]���I�s�t�' ��J�!̘�viژ>M�H�JɨTߛ��'���'cr�D>'� 6�O���O��iʀ�Z��Ɏ�5Fhh��D%N��To�$�'{�D�����|��M�a#N>pz�paI��^��(���	֟Њ3!!�M����?�������?q�O��ujTIW,Y"�2� qQ�6��	��hs��Gɟ���zy�O%�'F�I8�!Vr{@��M�n#��nZ�+� �q�4�?I���?���Y�'M�M¼��xaD+�}N�Y靛[.7��Z��"|��ZUH��p+N�}wT5�,\\�"rB�i��'B�m-F��O����OL�ɠ=����ȷw���Ef��-B�b��� +���@��՟��e-�T2�IX�D�BE��s���m�ڟ�b0*�3���?1��������[�s3bmy�"�r�I�,�]}O���'�"�'a�]�쀀ղ^�<u�^�X_����h1+�N�M<���?I>�)O� 6&^-C���&S�w�������En1O��D�O��$�<�D�8<�)�9Hn̓P�?Y$
�� Z=�Işp�IP�	Ey��˃���L
���ϮJt�|��-�	����Пd�'&�h���.�i�U��� ��lXԠ�b5m��hl�՟�$�ԕ'�
�}jĲA�H�� &��E��9�M���?Y+OV�"�b�O���<�Ӻ��qRe�����G�hoHPrN<�-O�pp��~� ,��֋�*yG2)��>��m#%�i�剜R-8,��4pR����X����$O#b>X�	�W���p䊯:��	mZqy���O���h����:B�|���"@��4 �i���"�'q���$�O���n)�>��c�	9,Nq�u���U­�
g�l�"�0"<E���'aX��7�B3v5�4-��T�Q#kӞ�D�O��$�fE�i%�H�IΟ`�8�D���ob��Gԑ:X�>��KT��?���?En/Gz�(qE�5r-X��������'A$���%�d�O���!�������Ʀ��A��}\9;2[�D)'�(�	���	՟�'>J�(���jVIB��"�sF�!%@�O@���O��OB�ǸX��+�A��%�To̡i\t�ӄS]��?1��?,O�ma$��|��QO#���b#Y5K ԳR��M�Iҟ�$�p�'�H5�On��"���;k��B��6��IY�R����ן���zy2D��9�����k��N	v���0�Z-I�t��������j�I~yc���'���Iu'L+Y�Jx�%�-!j���4�?�����I>P�&>��	�?I�HB��+��'X���٠G�<�ē��}[������5+�}����aR���o�|y���'D,6�x�4�'��Ĩ"?)�hM�u�,i��H#cKN�En�����'g��rc�4��'�,�Z�e�yy`0�C�BB��� ܴJ��Q��i,B�'<�O7�c��Z����Y�,DQgE�@~�� ԍޫ�M��/�����y�'fI���'F�09clگf;lx�a�cӴ���O����~=<t$���ß��ɖR�bx)`ő��DH�.jh8É}�&�&��'r�'�� ?�r��fMSe�  �1L��6��O�L�T��@��?y����*4g�,|�0 ��JH|02[�tQB�#���|��̟<�'�t|��T��9�L^20p~LY�bR�{3XO����O&���<�+Od�9�-�9ތ��!�̴/B�eC���*E�1O���O��<YIY�V�󩆡c=ԡ���qFl�'M��������v�my��Y9��	�u~@����YXjTh�eܤ-��	ßD��ٟh�''0]��e+�	�1m2����´y�2���Y��nZX&�@�'$�ۏ}2@V+\8r�Z�	�=�i�'`C��M{���?�/O�ի�n�S���S#\�@P�%�\�BH\�a�Ơq��
H<�+O�!���~��aHF�Jh�2�EmrH�4f�Ӧ	�'L��.z�9�O!r�O#��{czx�O�x�xV��!��moy2���O���]��iD:=�]pW��8av	���iΪ2'�cӨ�$�O(�D�|�'�����6�0-hT�^�z�#I��`Ӵ-kӔ��C�)§�?��	R=#^���eGW�N�����$V���F�'���'�
L�3��OP�$����Ů�w��a��+��d..��OP����O:�d�O�uY�i	�a�� U=m 6�/Q�=�I�@Bށ�O<Q���?J>��Vͱ�Ȉ�q�H�Kҋ��T��'� �S�y��'���'u�	/*�hkf�=5M�e��J�R�ص釨����?i��䓂�䟖b�~���K�%?�[b���,�����O���O6ʓx�Z���>� �s��S1���;a�L�YzV<:�xr�'��'c�IH�Z�tT:8Z�D�Qݜ���NV�a:n-�'��'�b[��x@�)��'�\��W.+R蹒�
 3I�pU㒽i�b�|�U�@�'�;�	�7�.qj�8AW��٣��C׌7m�O�Ī<7�;��O�b�O�.!x��_TP+ǡ^%�+gA6�<��M����)fj��u�TRP��-V�U���\�xZ�hC�M3'Y?����?5��O��Zr��<bc ��sϙ<n��b�iJ�	2k�#<�~� �֍8Ȧ����<1`�ybCڦ	�2���M���?��������>�|�wL�.�|-0�!E?��$�ٴTf�Gx��I�O���a� �4�$�B��U:QxHl��4�Iğ�`�N��ē�?����~r��C���Ҥ�R��TX�#��'4��y��'*��'��V) �Y?>�9��Ҁ_nLD�e�,�d�>m��U&�P��ʟ'�֘Gt���Q�˜S0-��d_�PaN�N�%�<���?����`��4%�
&�0�u`ٺv#z����N�OT��Ot�$�<Y���?��$�-x"R�PIN�l��J�Ǖq��0����?���?	��?	(�z��e���X)/�H�/M#Q�fm*$e�%.����?y��?	,O����O�H�uW?A
�#�k�i㗇(x0VX���>���?A����M�?�"=$>��艹;��8#F�'����M;��?�/O~���Oz5���?�#X��ҡU�;\
�{���	F��mߟ`�	ay"�ø+�T�`��ꟸ�r�L�#�����W Z#d��Ca�ߦ-�'�2�'��1�̟�i>7M�`[�Ő��:K�4Y ���/ɛ\��&#���M��\?M���?���O�e�¸y۶�W���"5���q�i��	�U�"<���T�\$JL�m��.U 0�"Ę�'4�M���ܸ)����'0�'����>�I0J��X�"��%�����%�q>`��4VPX�GxR���Op� &�ҥ��>|�Ȣ�cS\����i���'�B�[X[O����O��I)Ux��@�)br��T���UK�7m*��ݞuĔL'>��	�<�	���gL��sO����?�޴�?�"��'���'-ɧ5��u16���Q�0�P�@������dg��D�<	���?�����K �J����?Ò�b��?B]��s7�o�����IS����if��gO�ٴ�J�D7�FDv�H�IXyB�'z"�'`�I;�t�Z�O@��+G�d��'��g�R���O��D�O�O��d�O��8ѩ�O~ݙ�/C�	��� �N�lf�A�����OR�D�O �g���ӳ����F��d9�wK�DE��	�2:1�7m�O�O`�D�O"qA�B�O2�'8��)U�����d���JCe�� �4�?������K^<�&>����?�)�+�$-솹3�+2�  3��_)�ē�?	�Q�z0�������_�c%ʡ�`']�<6���8�MC(O���E���u���\�d��<P�'�l�Ӓ�O�1+u�q� 6��)�ڴ�?��k�h�i����S�'�(�Pa\�fCv̘��Jʬn��p�R���4�?a���?���m9�'d2�ǰG��q�$<FT(�.Ic7m˳
;���'��Sǟx
-`V4����;S�y�FÔ�M���?Q�==�UX%�x��'��O��)��}�@M�΀�V���"5�ib�'~Rx�Tj<��O��$�O�@P�AĤJ
�dQ��ǺI�� {�ɑܦ��	�?i�C�}��'�ɧ5Fd*<D��)f� ��%d����=�N��<�6�̶*��(Җ�y~Zw�����M�K���U�B
�±��'��3pL٤EG^�B��R�ܪ��$b�,5r�=���
d��1|m�A8���N��hz�k̯-���
E���M-�JU艭��z�
�^&Hx��b�v�cm���haK�珟qUf�c�բ7�͸w�ξ;z�h`�-[h8W�y�M�)M�*<k���/�ZTԆ�	
��xX�GD,XvM��-e�D`#�aM1Z�u3R�ԥ. ��O��d�Ojiò�e���"ae )l����|22$�Ex��
0�
�q|ܩy�Io�'X S1�r�##+G�F�=x�#70�,I�%Y[Ȥ5��7�fA�� ¬<v��=a a�ٟ�X�4is�f�'���w{
<�@	Da�x�I�/\�W�J	�IO�S��yR�P$6��x8 ��h\����aӻ�0>U�x2L�I�\�H��_�0���¶��y�,֊e��7��O��D�|b�D��?y���?���h	�8�.�
�����)ܞ2�ļѕ"�!��-���Ѓ?�]�(��b>�D.�f9@o��Q(@���cd�k���6���ZF�L�Y~8���.+Ԃ�p�ŧhf��߅�U ]���� ��Wq~��&LX�e�ɷ�M��Z�������<i#���8B? g�M �LY�<���=(�q��)Y7qsm�M�p�'�N"=��T�PAF�B�z���ٞ{.jL���Tʟ��	�P;�]2�Ɵ���ǟ`���ug�'d2Ԍ�d�a��Mcv�R���~" �.�(�qMSH���#��J2}��(%l^-t�d0����i��
0S��I	P�'D|)���"`R^ �5�-w�(�v�'�)F�'����,O�D�<ѥ��4��Urh�* �T��Qi�<)�я��U�-�)_�&�Kv�\-���ܖOQ�ɏ����4_3x`%B,���:Qk
5Xr,P���?����?��/O�?Y����t/D�z��9����7��EP�.�1j��C&7~�~uQ�4<����ľ\�*-�*#J���"�:@�nD��n	�b���a���+Ep%4�_�'H��[/�f䝃D�� "��4�N��T 
)��O����O���i���4�A�iᖅ�L̮؄�Ig�'d�Ґ��7�p-�3+\=RNz�ژ'�7-�O�˓N>,p�i�2�'u�ӄQ�Z�c��-124�S���5Ys�X&Pk��'m�
��R�K�ဝg$Z���	%t>�gZ�L�ip#gΖNKQ�d���T�@�ddT3|liР��w?���A�8x8ȡGO�.Y[С��R>`���d� 0��K}���o���H�O�,��b�.f4�qʉ�B��>$��$�ON��OZ�Ӽ�����4s
��R���3Z}��R�`ش{ƛ��'S�l� �Hs�����Ǿ,P�e�'�&���Q?	�����V"����Of����Y΁�SJ��x{����K2)��{c��,�����>�O31�Rjٕ"�l�T@
����	�0�Pр�.fb�l�J�"~�I%ӈQrՀT&NL���i^U� �����Iş(��d��?qWɞa_~!�q��	 �� O��<����>�e�,��)���>��UP�"]a�'��#=�(��y�g��_�Xu)��:�����H�O��� � t���0��O<�d�O*��L������?�@U�?C��;D��m�E:�I`?��R=�l8�ۓu:�x�Uk��,���"�%Ci$1�s3z�x5����=q�ɔ:B�P�	�+r�Te�����?�*E��?���?�gy�'M剳h��jw�0n$%��)��B��4#�Na�QD��z���
E,|�ȍ��?M�'<4�K��hӖ5��D��=\��1"Wr��B#L�O*�D�OR���Ϝ��O$��D�h1��*� �%{��j	�AP� L!O�4sbmP� <,���. �rk��-e.E3C�	
K�t� DEt�۰E^/3�t��	�Er�� �qA� 4Rw%	t�wV�1��
��M�����$�O��'|���B�.W��,�ֆ�;�H=��K�'P�1�0NƄ%�t��5휹-^�Y�'�7��O�ʓ[�@80��i�"�'9��~X*Iy%��l�
�8 $�n��0�t�ן4�Iҟ����)xR�}I&J�[���|��Ή���5�փ�W�@�Y dLR�',�`�*+�2��'E�m����� ���&٤�:�����!6�����ʙJ�'���8���?q����'],C5/O=WeA�`&^�T02��g�'��O>�'�|����M{�5����?:t��Ov�G~"	n�f-m�(R�C��^x��H&d�_��l`S�� �M;�E���Iџ8���?ٹ���ҟD��؟���e�#s@���C�#+��0�O;S�b��+��ˑ.��2��|ѩ��b>�N�m�}�F�,9��{���I��u�Չ׬&JT�"$֢ <��3�,�J�ϿT�d>,�Gň/�V	0��6vF5C�j����<%?%�SBy҈�9K��h���L����H��y�%ڢ?��ʆ(� �<1P$���OzhDz"��>i��Q<�fʇ�<
�&��埄��xb)�P1�mz5J0%�|�
�EQ��yB�]>(wH�����$���K&��y2)Pc���� ���"�״�yB�0:H�,�A��s*D�aM)�y2��'A2̩�U�m�mQ4	��y�
U�v`�j�!é_��1I��ݹ�yb�� ~r�y��,�V����˨�y�(W���왰�TDU�kL��y�lŞ!��%�^AX�*�3�BB䉱9/H}Y5�� �@�Yg���Z�B��5 ��`��Y$h���F�C�.��]*���k9Ҹ4��(<]JC��%�9{��,�ʘ�';6C�ɎS���e��E��J�jΑ-:>B�	16R���D%C���CS�L&�,B�	�H.ڰs�bۿ;�,�!���y�B�	<4�8��q^ĘS!�Z�J��C䉇Bz@����;L�����E�bC�ɞ8���ש]o�|�O@�^,8B�I%͐�#�IOF�0`"��4O�C�I��a�2�.��X����t��C�I5?�� n�d���t�^�f�C�I�cD�z�,'��p+ZLC��4#d���f�/1�60��͘r$"C䉴|����D��"d�ZU��+�LC�I���X��Yf��(�aȓD`C�ɶ�V�a�.ֵ9}�����7~C�-<p�b-��_@�%������B�ɑt��R���S�)@`�+m<�C�I�+�t�VD�lix]�BΕ���B�ɰq)*�dπH�B1:#Ԛ=��B䉋Rl�}"�I�f�	p`@�*���uΘlQd,С��S�O��q�FT8]��P�(֍=�2�h�[�<dh��
>���Rĝ�	�rF΅b,��T�+}�휼KE.Y ��,��)V.��s�T��7��@�0�r�|2��= ��1�v�A�"eRx8�D%���^���
S Ȟv����(u�"I�ǋ�p�����hw��@��CD�g�	�:���[G��!���C	�1h�A�����5Dj�G@�]�����,�3?��^���7��&r��SQ�In����1C�>Ӑi&��U5����i�]�Y?l�D����*>w�90A�ε~p�d��N\$,���wo�c���d����[� ֽ7��\(��nT#���Z�u�8ڕNX���9��c#w*����\�6��ф���dt�"}"�	f�l0�6�X�z����f��>���`p��$2��ƫՑ)	6E$��v�G�c�m���ÐV�.x!�L����lC�^^��BJ���(Ҝ&�Fm��J
�9~�b�l��B�y��a+�� j
"�k�b$�dR�����dØG�xhȦ�T c&���b	(:�6�{ ���t 0bJ�o���>�O�l"Ң�}��d�'��}aȽV��b��-ӣY�:��\��'D�5xd*K%,��I@1N_�q����ӭW�g�2Tà��4c�)��<ѳ$�6}Hc���H�q�oPX�l��΀�e��b�(�`��@�� ^��h��:
��r��b���=O�٪q�X�W��a���̥ko�1���.���KP([�l��U9��֔t�8�F��ēiitp*�
T�
d	�%�j�՘�B�B�Aw�H� ��DRu��.|>"M�vl�.�����d�6�n���.��c>v��aږ#[�'����M� �Qv ��d#*8X���,.�e	䨛0%���J4���5#Z1�`�u�ԧħm"�0&Eҟ7�8A���+<n@Tڲ)�.#�$�{7�Z������b���M�����2;��T�W�Ʃ�Qe˱U?r�a?c��ы1�~��'���ϻ�p�����x)��3b@�8�|}	{��u7IA	WpRA�c� �,�L���",28�2�կ.�@��q�B���%�L���9;~a��Y��2�BP�6C2q ',�3 ]����B�pM��ϙ�d��&p��c�&?N�$��b��]�]�ٴ"�L��À� �27k�'f�<�v��m�L`�\�n��$N�g�X˓]��Ą�xY��`�E�)?⁕'�L�l�1�~Y�t�Q�3߶<1'لI��['��M�w�ӆbvڲ&�
X����Xw�r��6U?�iR��'D���b(ұ�P�q��@�f��|@`�Po"�<~�Gy���a1nR��v�z&,�Q$K�6�ީ�$��@�����A��9!I?���u�>�R ���Tp�p�s�Q3\w��4&�(YH�<�S-0p�q�A���0>����B�>�8T�5�.���Ԧ�m�<�q�o
-|X�m�<��<ؾl����3P]G ()Qr}s��7pvȠ��b�>���#>F���GŜW�.�!����8l�H���nյ��Z �O�7�@e���+2��y�\p��?y�L�E �U{D�A�l� ��zy�I@ ��ar"K��<��7�f�<fg����O��p�EX;@f��b��I`�]�Wȟ�\0|i�KD�<L�d�D�5:���Kѷf;D���Z&q��]Ey��ߑ[���)W ji`�C��\�U��O�s��&��䦟֝K�<9��_H�S �K![g���S)��s
�����O�H�Q$�[����W!�꼓P$ۤqq���&QB�uZah�	��	�x��oZGܓ�?���*��I*�eB	Pْ�	5��>�b�Nǭj���F��͉al�]7� �S
D�d�B�`\��'I��)�.�QY����dW�F�؍�e��W�Vl����&^�7qĉ��G�f;�%?O�M��Y@f�$)�|b��0��lӠF�%��'p���p�>!K͟k��w��YK��%>���b3�7 ��O+	p���ς7�&p��i�U`�%dx�����S�*+:�G��� ��y��<A��~,�έ����z�x�j�&b� -���,O��������� ��G�s��t�Mj$��ׂ\�>�r�a�/p\�Ik?����=|8�|���2`��fa&lיּ�1��}��C$��=���A�4t�,����7��xC�'���	�3�\��Ө�� Dz��
�<Ff ������
(r����\l�7�W b��c�(# 6�f�RlW�{�� I��b�E���ˌ*��r�1d�ZX2T�Of#<�#'D�yР���4�n���C {��CG�'��>���i�*�b�-E6��� ����@�"�O��=�OR�-λ��+�@=0��ZTJ�/L7�����n-�WK��>����G	X�a����̝U��y���O���CH�Z�����ܽUx� {��'��D��#�F,"�`̯AMn՚�����"�� VL��P4�ǀf7��I�\�($)J�6�@l�rZ q��I	Ѣ�cj�SP�Q���8.|�=�'�y�����2jp�hA�Ȧ��%˿ �r1 GN�V���G��GxRF_�^�9qGZ�"�H0An<3��$i�m�37�}R��(<|y���~lhcnK�oUj��˧�XF{���5��w�����03��-`D!�^�0�R�0=>`�����@PZ��q	� ��M�K�x��C�ĥ���u�0@�]��x��G��O�%Xp>~�,`�#���w�f�����6M-�	����@N�3���5���5_�Ġ`��Ǳ�:���+@\?� ����r�]���2�ŊO�'�B����_�ze���!AT�q�E��4<s���T��O$��7fʂhX^���z删�M>��-@<.���Z􋍽f}!Z!d�M���@�~����o�<*4��%
�u�����������<)U��G*�'����<q��c��c�w��!+`R8H@��� �#�O�-��	'�?��nZ��ͭj�������!���>1%KF# ���C[\���%�?l���K�K�'�\Y�%���<��9Z��陧u�.�LBb�[�N��-L$Q�n��Vn�$F�i�6�t�8j�.��ўd��avb�����<��b�2C��^,�?�����gyP�D�Ob����.�dH�/*�(�W@	����cH;u�F6MU<%j *�<]��˄A�	7,D��&yL�������$*�S���޼3����<S�l���~�xW�XX������pf��R�׶@�P�S�Yg�0�b�)��'F��ǖ #P�Q�2��2�j�	.1 o��u��̢��C֣�HO�u�җ;n�I�k�*&Q���%�O�=I!kR�jf�p5��yɪSC�O����n�(����o��z�T<K%cJZ�'�hiYeᅋqj6c�LٷJ"���4m+,�r5F݆ �(�RaR$Y������O��",�T�p`�E��#��0��f�9nB��E�=�Ot9�&%΂uwD��v�(�,��M��,��-���hO��"JY�ΆE�l���S�,p��gg�	Z�a}��ހS4D�۴��&6a�dH[�t�T�3"''&B⟀��f�`�`@K�4T�1& g�B��)� �MS��VD40�#ڹ9������6>l�(�b�Z�ȓ��<���i��3�?P	�9�.�45,  ��O��H$�A�4� ��e	�t6☂�	U���"'�����p�OZ<P5�7-�dĕ�+8.�H���N*��,b��`�f���uX�)e�nb��+@+�ڹX�l�D����;�؄��Ǜ�h0�K�'�.��M�~y��0��'.��=(��Xj�H��Q�V��j̆剑vTt�u���b��Ԛ���Gn�<�eO֐n���٤��8�b�F��tzt�OX�)��o��O�X�� ��;9hp{E��z� E &��)�(0�s�2�D.�NPb��./h��PD�d���!��Ӭl�M0tc��A�xP���Bz?�'
�7������aF�AM&��@�P�ɜQ
��*��MvWN驓�N�IM���͎r�5�<�'l��vB_}?�4�w�Dqr`g)rf�dQ��(I>�5S�4��� A�ܜL�*1!�7�eMD�X�����$c� ~h�x*ci�ӌ�O���!�~�cU���<�s���B��\3n�Pԁt�ާw�J���� 
����&\����B���n.�H�4aY.sk�ȋ� �&����)�r�IC�~�� |͌,��ʏO��� m�@��dg�-`FN�){H�`� {l 1vʝK�N`�I`�>҂m��^�^V������7vZ�&�����'�Z��'%Ȗ^M����m=�x8z/O܉�FZ����0E�N*���3�ˍ�/�����ZퟤD{ʟD6�'Fz��A��7� ��,4��ppd��8_�L��t+X�@��>��?�n��	�]����Q��k�HI�:�Q�D�'����С��ZH�!J��\��yGa�;N�
�Fy��ȼ 	B��T���{Cid�����W@��]��ʴB����dW���2��|*����p����T�������U���Sc W�2�^�X���$�:C�����K����Fz�"ԄG��<)���#| ��'o��(O�à*Ĥ)�=+���c� ��#W��  [��QX&".n��t#݀J��4��
���>q /5�v�9ǌΫyށ���/rR�RGe��3L�����,� �p���Ͽó���F��h� ��H�]r"�LF�<���2V~�Q��Y�B1HAƠ9���(���O�~�U��<?B0JE
����6�� � E��k �4��y��t��(O(��
�/(Vf����X�r ���#�� 8�l��F)����ğ�ࡰJ
�P�F99R��`k��5�Y�d)�QbL7f6q�-�e�'n�$�b�Z�J�P�Ը.L4m�OP#Ç�'&V� �1ƃ�!)}q$�r�x`fM0X�<�=���dY��I�!E[67-ZT�g�	���� ��YҴdqתU�<F�����d�O�#h[01�+�;+��U9B�|��)��$��d*Dg���6��S��&DL����	�Mz:��D�^�f0�Yj����v��s-=��L�sR=���������u{1/�):���"F��#Ĉ�@d׋l��q'X���,�u/H�]℘8F�X�@�v��<9�ұ���A�W"(���$��9��'z�� ��b�(Y��!Z�~$��yI�KxP5x��2Z�@����/Ԑ��E�W� ��T̓�OTA��#��KB�j§E�xi���E��B� �Ȁf�ZU���*Ok,S�(zZ8 �Z�==�x�w�}T�'�z�Gy���?�1c�nX_����lP�8N�x��!�|L�bF���9CǇ�(&��@��G��D�6MBnՒG7���O�l��"̊en��,8h��ip���lA�D&�+&ȝF�X��D/��ē{B�JŁN(�,*�ؤ>E��?͠t��,4����ҤQ#�,R`�,
���@w�o�4�qA�E�`c?OZ��pg�Y#������]F�]���;M����1J�.\�8!�a��{����i��;�#74�8AM��B�`����s�1�tKC�ST�	+�VX� �v��/N�
1��gв8��8ᥙ�,���@� ��,�����)��[�y��u�x\ a&�t�J1ւ@���>	f��L� ����S1;v( ��ʸk�:$[O�[8�'W�tJ�.�78����Ab�<B�HƔj�Ȣ�*ʆM�ў��Dm��z� D��,@�1��!͎�jȝ�p�ف8M%O>�t�ɡ����;V~jH�q��9�1�a�@�C��Zb�P�EJ��{QB�/D�m�B䉼"8�A�	�Zo��@k֟2�B�I*)�Dp��A�@�2��"�N��B�I?}�@,�� ş��;7P�zB�ɻ:���IP�,�:��a�/FKdB䉯� �+1*%_�<Q��O��om C�	)���~��2��Bd|�B�	�9��@F��4)���l\�c"�B�I�6lLڕ�]u2���ĕ�FVlB�����{�̈́ ȹH`-��H� C�I�_O�&n՛6ҢѺ3���oߴC�ɷ=��J�o;�~�8 ��	��C�)� �9农2+���J4$@6w� �9�"O���A7n���"SR�`��$"O2�)gL�>�L�@�SO��)�`"O��p��B(�����k�`�"O�9+5���k��,
/��B"O~}���F��HaV�0#��8"OQ�P◡\`@
������2G"O^8Q�lR�"�(�3��}�n��r"O$u� J�[H9��=�
�3�"O܉�"M�3/x*!���]/F�88�G"O��`��bŲ��X�1C�pz"O���u��.-}�!�ҳ3j�Z�"Ob�xR�8��x�����l�P���"O�1�<�Z�P��5�"O��H��Q{�{TN�>S��T��"OҀ��� =3fY��	�@Y�Ih�"O�8��h�6C�9�KI�eU-k"O2<2�аK	��b�i�.P�y��"O:�����5�v��'�;?Z	�"O�,X5 I�x��]ǧߐ_l��B"O��cSe�"e�JXt�ˇf/�9Y�"OP�4DV�Q�*<x��(�j��u"O� ��	�h�0�9��<t#Z0A"O��u�E�( �Ӭ놴c"O|9	R�<�­����e��d3�"Oh�hΐM���r�g��%ɓ"O�*2�F��&�9'�ĿW���"O�[S���<8��q@��C��)��"O`�`��>t
�#�3P�r�H�"O<Pza�^�<e��G�5(02"O()�&��;E�|���g
`i��"O���P��(\����6�.r�f��"O�TU :��WE�RJ�x��"O(�FΛ`0���%֖I0�y�"O(���	���T8Q���!
��a�"O|l���Ә�Z�	��2���"O6�JA�E�"�8A97�����"O ȑ%��1#~��s�T9(�dI{"O�1�0��#K�<` 畗~���j�"O��ǐ0o�J	�$B�/���"Ozq`d�[	l�(��d�
~~֔;�"Ofa���E��p)M)~�d�"Oh��(�g$h�0�̙^���#�"O��1��Xʎ4p��%]iPA�"O�EY6�$#�H�ą�`Q2��"O8}96b��M���5��E:B䒷"O�Z��I�dr8��E��^)^([�"Ox ��gX4O��e{7����XW"O����〲0v���j¿9�y3�"O�|�ի]	o4>=@��� gh@�R�"O�x�vf�t�����L�:[X]1�"OF�v�X-\fyX��O@��
t"O��j��2~ת��%	��}�:$:�"O�HڴE�5u��]2BM}�<@�"OXg�(aI)ҍ �S���RP"O[c �: TUⱭ�g���)�*O�t�Bƛ�MT��&e�<�X̓�'����D [��K�c�"�
�'1j� �)��`����k�z�<1�.[�_,�	��
��IW�_u�<v��$�\��41��ٚ�� \�<a���<�`HK�N�82�
�K�O�<�Df����c��ԋy��iJOs�<9%F%T_�`s�܆gOl����x�<� ��U!PGxm�  .A�<�DO�A"��6�ШQ�iQ�Fy�hX�B7D�L9��PEr������v<;3�!D�jt� K�LK1��&2%��{r�?D�|�b�@!P2�T�3�2v#:5[�� D� p���Wީ[�ԩt��P��*O�b���Dz��S"�ߟ{ղ{��������+k� ER�@��3��\��M�8�y��KT�I�"�^FR�	t���y"��H�޵�g_�z8ң���y�Mܘ/⬁�b 	�U�� �C�W>�yҌ�*4�h���D/?ɀ��BbS:�y���?oтP�Uf��EɼLe�W�y2��]p��B@�T�'{dUc�-�y�@�3&2 9[�� F0��L��yB��z��1�B� ,&�&x1���	�y���,��ytŵR��+Ġ��y�Q ��AI��]�����&�6�y"c�?R� Yv��%&��8I��D:�y���G���FQ�":Kaj���y"���e��I"5�I����z��=�ybN�-�.��1���\F����_�yBo  f$haV�͎P8�q���)�y�k�0��l3�ƇZ��\ �W��y�K3`h�yF-�E���2�m��y��ڳ%L`D��bZ86b4���R��y�!��̳ī�E�`h�%	 1�y���8��TLp\�`+A7�ybN	/m�z��B շ$�!�G̔�y��P����/�%T�������yB�]$F�@��\�N��ӱ�#�yRLY&n�P�3U�ŅM�� RD�X3�y�k�8F�}�4B��A����3��*�y]�'��z =h� �#C��y��	�	-8���
�<��ԪWEZ��yR��%��E� �Δ94�S�-�8�y���["�1􏐯!������yB��5/�DaڈE��hq�Ρ�y2�+9f�
!`��څ�Ӱ�yr��<J�� ǯ
�d0��ӊ��y"D�0�D��c���P�Ӂ�ӧ�yB��
Z? �kg!�4ô��E-�y�M2�|�b݂�ac���Py�l�{9���
�:?�����/p�<iCL�����A�L�`5�Q��.�i�<�q�F 7բ2˒�^�`��c�<��-[H�Lt��D����7/b�<AgJ�mh4�P7�ƛ}���['��\�<ɕ�>f5���U�ܖ
���R��L�<QLդp��s�IFpɺ��f(�L�<Aj7M�6�ۢK��U����%D�E�<	FB�D� 8�3�*�0pK�jE�<�A͕6ܶx��/�zQ\m��j�<�#"Y�^�H����@��Jj�<	����b>�$��	�4ժ���j�<!3��
95��S7l�t�1c� e�<	��@�m�D\`�!x3�� Lb�<Y���9>t���
�P°�����Z�<�DU�>Fĳ$D��O��WLXA�<)4��! Tΰ�T
S�b+ m�dD�C�<)�`�8#Ȕ	�"�?�4u�G�S�<Ɋ��+���SΉ�s��}��&P~
���0�	�K�\d��gF�0F����!~lB�ɻ|} % ΍	��9�rB�����	_��h�� hݰd�{�:|3!�ǂ?&=�d"ORqA6Gz��P�H Q�0!��"OF��	�b �*�e�A��	�&"O���P_8'��ʶ&F7
p��"O8�c�.�����1=�&	p"O��rF�[�)��A�GC�Zق@��"O
���%�+�d�F^ '��4�OH :'.��q?�њ�$�Gp1a4�,D��8sJ\1Wb4R��nC"8P��+D�(���M�URWɒ�<�!)r�%D�(���"�{*��myYd�#D��'��+a�&,�Q�>!��I
�
!D�J�͗��I
1�Z�T����v?D���㖑6L���Ǚ{�����=D�L`���\h.A�(?d谑�=D��Ɂ��GH*� Ӎٛ� ,c�=D�p`��$P��,���u'��	G<D��xU��?r�	��I-�����9D�Y6� �8s�5�Ī�1F�ms��,D���B�rԘ�oP��:Vbm�`����nv��@G�D.Y�.�����
6rC�I�f�8c�F�M7fBWb�MT#<yϓT�0q[cn�5�\�:��ȟ07����N�n�'AT�fOr�b��%����ȓEW�dA".�4 �l��:|��܄�uj�(Kb�KM�4��QkP�-�68�=������ک.8��S
�(C�zF.��y�LM�^�n��ȺM2L��mC��yr�*$f�M�$�?<����8�y2̐�9[�5���չ8�H��GL��yG��W`~��I�< ��H�yĞ�k��$KƑ1��x2�M�y�+̊1J
=����.q��3���:�y2·�m�����"�|��U9�ybD�6v��	y X�p��ic��ҹ�p=��}��;'���Y�j������y"�9=��#ƪ�s������A*�yb�O�0p��k;>U�"����y�(�iW����e¿CⲘI�ہ�yF@�h�*���=l��ƈ�.�yrb�~Lș� d�;f��x&���y�H�*Hu��拽]������[�y��_�.n`I-V�HTeˁ2�yD�-0֘-�ǈԶZn�I24�ۧ�yrG �q{X��N9YƊ]�(���yBA0
����\!`� �"c���y��F]y�K��-�rHXR���yr�I�P�FN�	#�`I��	��y�!)=��Ģ7ڷ�lțFe�ybjT-?n� b�iVp�.E�vW+�y2IȒ=�8Xp�_;u�vQ�*E#�y⥗1o�(�����6c��y�K��x+����%[ n�Z5��ybL���^�p�FO:2��Au���y"��F�麱bɌM�ȸ��ȓ�yb��*k����[�rݜ9�JV�y+�1����Pf��2��x)����yRH�8&Ωڣ%�/\�	Q��@��yB�F�Ey2I8"��/QDl9�F��(�y�`X8٪1X1)=x)<�� I��y�n�/H�Hk�GNpT��\��y�n'���9@D�bl-�����y�����@)x�aX�/�X���'ϰ�ybΑ�y2���N�!��r�kى�y
� T���L��)h�S�&��w���"OjԻ3�^-J���de��^��8��"O�ё%�Edj ��eF�u��"O$Xtm�|?�D���x[��R��y�n�&�����?7Ԛ��d�؎�y2oY$t��+�G�C6Ddȫ�yR�gn�p�p�����8֢�y� z���IB���~���F�D��yRo�#Qb��d�| jFM�?�yBI�4R��q��$c'��h�'A6�y��<�<ٙ	�c��;���y��ˍa����!��\"!�6d���yR�Aa:���J�B-�g�=�y�aW<Vq2ÆF߽v���b���y����*A�)�\�A�.�y�	�+�l��g�"����y�+C?R����ș��h�����y�@�0wl�&��J\ aÂ�y�a��&��H!��
�6 i��y�ߠe�I�'Y����'�ߑ�yr郒<�8�'茎��IX`@��yR��fx�BQ��%t�<`+�H��y2��O��9�#�Ǡj��y�R�Z-�yF����1�S��fC~�����yb Ð��@���f#��O��yN'_8	#U
ba���7�Մ�yr�ˁ}��d
q��`��=:2AG��y���� 9�U��\�&c"�yR.F3K���{#� �{,D��%b �y2L������/�z�������y"aF;�vA�� �rbPy��@ټ�y�+N����Va�m8,���y�I|+�q���:��Q�##�y��K����H^7|�L��7����y2̀)?��5��l���a���yr!X�u��t��fK�c�8b� �y���6ff� ��0(~��J���*�y�㜥 �HQi5A�$�zh�Q��y2�P,k����菷nI:���Q�y���R#Z��Ad�
b�<X�g^6�yr8T��H��@�|�;sF�9�y�nˢM��-�#-R�$:�T��͘��y� �.r�l�xb;�D�A��[7�yX�0���c��D���S����y����`�*)� k�&=s�D"���y҉?4v�9B�c
��\BDFԡ�y��Ι+���21)��|D$���B�	����@3��&ƚ�U	[?t9$C��Mt4����ѡ:��Hc4�\C䉺x�vy����v��p)��L�6�C�ɬv ��R�D�o�PHY�J�*��C��8Z�4���WH�������lj�C�I>Lv���d$F����J�j�JC�IBt^����l��\��	$��C���,Ѷ�`|��@�ג�xB�	�vRH���؟�&��r׎E>B�	�v|���I��&1k
�� �,B�ɳKX�%�NS�^���-T1B�ɺtY��J2�U�/y^�)�!@[b�C�	+HR��ɗ� �,��kQ:U��C�	�W�)��v�t�ڲfQ ij�C�I�,�Ɲ��n	��B�*� �NC䉱_E�1# ׂ1�<pb �K�:#VC�	+�@�����s.�T��I�U
XC�)� �t#Wm̿i��D0T+]>!h"O@1�D&�f��� ʁ�gLxX8�"O�ũ�Թ�.\҇���hF,0 &"ObaaAC(�Zy�4�N�6A�&"O����ڙ�����"0 �Ig"O��iIZ3^�z䉤F�}�D Q�"OǪ��i^*pa�,�1x���"O�rvFRZ#�\�Jܸ_���z�"O��@��N�e��$ �j��UzVl�"Ob�#��>B�0�IǇ�Zifh�A"Ox��) N��KslP�(S:Pˣ"Of9����%N ��ئL�!np}q�"O0�z�a��[�<���jY$�JM��"Od��B��4�|8xs
��H�"O�%�Md�vPs`� l�V"O����R
\���N ��%��"O&ĸ�.,>�j)�d�L��a��"O04X�G�~�R�ڂ�����t"OP�Q��yf��kφ�\�%"OV-�$,ޘ"a�%�kL�rf��6"O0�Ѵ�O�\���@�_��|+'"OZ���֭"D!�.Q8�2<�"OD� �$��-�>0QE#[�.<�MF"O.��ĉ'��U���"Ԍ�J�"O��S�d�gR$1؄���fa[%"O(��Β�a�.�C�R6s�1��"O��4����P٩�ȓN6��$"O����A�s`��¤ǅ)Ov�[�"O��+P�ד2�v���$ޯa3�j�"O��G��%3�Q`�ůg>�t��"O�{�oJ�2�����O.��`"Oh�ڧb�%u�ؔP3��!>>E��"OlP"�R�j�:պ!�@ %E���"O��@��RBL҃�_4>飤"O\�h�ŌM���cv%z\ S"O.��m�$1GTi�#�f)��"O<�	%(�)�}�w�z�
�3�"O�4�aT
��Rc%��%|�ĉ6"O�ss/��P) ���c�J����"O��б�Y�}B�]d"�Ak*,:�"O���w��>HZ�0�'�o��%�R"O�������� �5��-`JvL�E"O��9�S&`���j!/R@���"O�t3ƟlVI����g*�2T"O��j��Q22�J}K�ߨ���"O���D��0��yT"�Q���B�"O~u���Щt�N����[�BY��"O�<i��܌5U�A��pYq"O�h(�	!6��hqO'gPr�"O�p����
���z ��M�K1"O�a�!oV=;>M3��
B2i��"O
�{UJ�NQ��A�䒺e��6�*D�Dٷh՘�H�CWLˋ\�`1��'D��Imm~Y� ���!��U#�  D�S�dJ-5|#d�u��Q)��<D�d��ά뢁ˆ�GI��뷥&D��9���� -�|��,F�5�,X�7D�Lq��1J�y��Ġ����2D��r��:u$0�u�L�'�&)b�3D��p��%"����CN�2�
�J��.D���
��zi�rI�$Z�Eۇ�9D�0r��"+Z�A��Wn��'�:D�4{%�ڃD��y�T�8��d�#�7D���D�Ny&�Rd��-x�b<�ee6D�� �����eq��J,�~%�2"O��Ȥ嚈d`9�O��+�"OҌR��"dH~�	��/.6�"O��B�O�*0��H�E*���p�"O�(���8>g������$q�R��"O2'��f�ڼ�qDR��İ"O���EMO�B�z�"cF�)[z�A�"O>�8'�B�^�����Q�ld�v"OƵ�p�8�� x��	�A��:�"ORq%a�Pؖ�$	�2 #\В�"O�!3��îI�n��a�l!R�9X�!����v:(�a��(Em��i�*Ͼz<!���}�<���y3� �F��!�$��!>�p����h�:��Q/(!��XF����!�0\��
�H�r!�$H ���j������n$!�<FB�ƧGҜu���F%�!�� �S)�d)��Ò�6�X�&I1!�D�
%Py�*ӏc粌:cʞ�M-!��W8r�����	���|�`�д'!�d������OR�q���CVG�'!�$�F�|Ap���N���3��K�!�Ą,K��7�1J�=�B�J�!��˲hL���7��%FL�0ˇ	�2k�!�$K�rp��%֜7� 9��O��!��+!>m���jI�D�9`�!��=Ḅ"����E�qq�D�!��J�a
�1���J�7����8|!�D�����R�/K�t�ƹc�ĂRk!���"P��0�W*F�5�4���W�N�!򤆉���{v�7<)d�����,�!�D"��h�V� �8!vf�Z�!�Dlw���G7����B�B,9�!�$����$%�"a:�Hj��1�!�D�	e�I�$bF� &��2Q�@�R^!�ė>N�JI ��X��Q�n!�dC
N_�q�H�Ym��k�/Ÿ<!�Dߓ#����
Y�7m��p7oP5�!�$�0&J��g�"uT�`X�._%#a!�d����Sׂӷ>?ޔQp R�L,!�$C?���ЕG_�;P9:�O�:!��\�!�~$��>Y:<̩'��<!�� �!HIѳʎ�`�<Ԛ�EQ7y!�d��tA�!�":�b�5G�!�dݾ�8���Xۢ@�@��M>!���n��1I]�F�^A`!Dެ!���e�Ҹ�DK�%Q�����XN�!�R��y��:+�P����Uy!�T�He���$�^:i�1R����!�D^9.�����ϥ}y�� �J/X�!�d#�p��̌@�9Hr)�{�!�Ě�e{
IƆ!s9���#�;+!�$�*��H$DS�(AHti�G��7�!�D.[���{ ��E3Dܸ�Ӻ1�!�$��<�����<DS�x��I*$�!�D��EcB�[wZo@P\ !��8o!��H�օ�5��1:��FUYi!�$ ��� `�?e ����Q�]�!�DBy���)P��n���"��;!�ĕ�|3N�چ��
l��D����!��uc����.�u�_�#�C�I�79�(Ae��:"K�����2�C�I�Z�n]`����5@�!YR�Z<\�TB��f!� �wE��]Hzy0n� l<B�)� �%��h� {f1��HA�E�Z)��"O�`rʛ�!4fh�RfA�F�1�"O6� C�
�^R� 2��$�J�"O",��T}�����(�o�!��"OR�� ����j$.F"}�(i!R"O�u��S�I��=`b�W�a��U"O��!����) �Nƛb��W"OP�7hR�^�d.C�k]�q�2"O.,�e��T�f1[��є Bމ��"Ot�B�*	
 �#�m΀��"O蒱�]6 �0��t�U�$�"On���h�e�}JrJ[2[���B"Oи�k�M-p5`7JI#.0��"O���b	H�_{�,�%���ސ Ç"O4Mfhƭ;�ƥ�"(�Q�ZdS�"OT5�
֥}��	ac��t>,; "O�1��E*P�|���F!]�Y8�"O�C���*@溸�2Hl�N���"O&	ZYh��w�?bqB�{���2E!��#|��`�A�{h��2�ͼI(!��0�@\�'�hUv���W@%!�䅁M����=*Gi���
-L!�"�n�� �Z�+"@h�A�<y�!��L�-4��2k�a�P��7c�T�!�$�NL>�8S��D�t����oP!�]&a0]�u/�>h����5�^O!���A+�hX�fY0T���$U�1!�]�em���r��o�ؕBE�ׄI!���{g���P��?K��u���s!�$��%Ǟ8���Ǽf�83CHZ!�[<' �q!թA�ie,^"s�!�D�C��P	T�KE�:(Z� B1�!�DV��`Ep HՆL��L20�D�%6!��T~����U�PgƠ��͚>�!��5g�Z�i"��grz4�e�Q�R�!�ņv���,W�~ѮI�Æk�!� $_��)�	����Р��ݣR�!��@���D�R���2�T�j�R�!�d�V�X��e��8���j�)�1&�!��[�txh�z%c�<2�p�r+�>pu!�%ݎŨ��7l�l���A�b^!��!V�"���(#$��-
�Cs!��8A8�� ��,&�2%�GP�lb!�DK�K2x��%�$ے�C�&N+"�!�dM5���`ҟc�zU�%N��!�X(D�|A�G�va`�$�T�!�
��8 :"N�s���i��&F�!�Ңx��6 �z�ԹSF�޷7�!�BEx��rOHۼtӊE��!��q/�8�4�]6zjI����F�!��eN��[K�E�^,I�n� �!�d��HC$�#!JN��P�:��-�!��
�`�򀙌u������`!� x� � g�
S���.��!���8��G�
 ez���ˌ,	%!�V���!���	d�8�����Py��1\-r���g��&�l9a��U��y� �/�Mh��p�cCgX,�y����]yU���,�
����y���b�ܰe�ڲ
�&�	S�W��yrm��D�����'[�.�}���F0�y�HW�]�\��A��3R���Aa�yr)1�T!��S��F%j�*���yr�E5w'x���k\,�܅� $���y
� 	�Ā�S�Z|�c�Q�8;�"O�I��i��p��O[����"O�ٛ��ҏy��ՁG-\�vrl�"Ox����	E���vLݐ>h\���"O�JR�@'\V�Xde#AY&��"O�U�6���<a �� %�*C!���G"Od\0��\�BH��w!U�r/(ȺG"O"�B���; ?B+����K���P"O���c!/;���`��ظ=|��E"O��D��Q"PJ��� ��"�'�
�rhͶ��i�إ&�L���'٦�ҲgZ 8jX(c��� b��B�'��4�v��$u� ��S䂰	@�'�j����;z�p���㈌F�F�c�'��s@8�e��o��&`��'��(��K�%��1%�R=�� +�'h|}�E]�,a��T�����
�'WP)r"���:�Bl�0�"4:�'`� ��o�c*�U�M�]	�'���qK(Ib��H��
|89��'I@��"_����c�vE2tz�'��,�F�Ig��p�N�{UH��'kҥS�ՎA�\t��H���(m��k�&��m�}��DI�4�"=�ȓ+�:�k��K
�dL7��&]p��zw�c����W2�3!�^1i ��ȓu��Y���C�;?��&���T� Y�ȓ\�� �aߐ7A ��4ក�,`�ȓ��a!^;D	��R�Q�@�l��$�����PQ�g'��K)ʰ�ȓ=�¹�¯]�ZLȡ���,khpA�ȓ,�:���&ӑI��`Ƀ.�?5�̬��*��%�*F��9��L?cmH�ȓn�Zp�[�@� �ߦ#qĹ��x��,��	��(X���N-v.���h� ��k�z���(w��Y8Pm�ȓT�F�
�ʎ	��,pd��<�z(�ȓ~��$J�8h��k����
 ��-Qn��E��3� �Vg�.[@��ȓs;d㓌�hAhe�v־ArP��B�lx����D�R��Rtx�ȓCp�Q1�-��T�p�37 �����������+�'9\^�c��a�N��ȓ
zh���B�2G �Ɍ�0Rj����ƹc�̇8vtl����~�\ȄȓLA$��DfOKx�0��0�� �ȓ}��Hi�/�-*O�yS�'@�T��4�ȓ`Dt�0��#&催eNL@�Ґ��z��yj�a�v��e8��X��Zu��T����⽁�ٌ��ȓm��pJ�L��{@���F#�>[�����?b`�	�K^fP���R���ԅȓz\A�Hؔ	�e@�!۵9��a��>]^QQSL�$A��k��
PÊl��S�tA��i^�"g&x��-�:�^�ȓf�43]�H��d(�<;.$��ȓg�ũ���1yθ�x���"I��Z3MĜ;>����w��@��i$t��.)�\���"�#S�����e���	1��QcW�F�����ȓ?�"P�`�F�2Ԃ���:j����'ʒH�RA��o&Z(E¶D4b4��u�ʈ�%M��3�(��gD1����B殰qo�A���b@��u��S�? �����T�`���'�4)�"O�)�V��L�Ȃ�����+4"O�� ���2@�ՠ�����i( "O��˷K'a0T��<r�ԻD"O��ҥ�dM�¥ 
.lf��"O@a��7��UB��E�>	԰��"Oh`
d�,#�l��$D�!�F�"O����ּh�V���"�
B���
�"O0U���=0b�{BKI>Y^���"OJ���aU�ZHY5,�#j ��"O�C����b��A��+sb8l��"O��A�*`!������b�N]BD"O�q0׈@�^�z	��Zw����"O��r4� 0� (Ȇ��<b^�j&"O�1����bд�q��Y� ��G"O:�2`�rX�!Z�ćD���t"O<X�P�L�.�Ȩ+F�C,Mr��"O�����*�<Ċ̋�q-�=��"O�	��G�,`w��­_�Ry�J�"Or!���&h=L�cQޗQp�	�f"Olհ�M�紙Au�� D2dhc"O*p�@��[�����\#z j`"O@�󯀦�T���T�H#2�`�"O �zW�0W�nT�� _`z�`�"O<ܨp�
���/��T,���"Op���j��a���|)�"O��
�R:wGN|�N֘W�hA*�"O�!F�@�^��t!���q JQf�<��/�1y�9�hQ�<��R�%`�<!  	8i�Q�!V"�����E�<�Q#����Ƞ,`,�6��@�<!��n���hT(��=�����_|�<�����$��5�x�Ĺ�ՊSv�<ID��6F�S�eN����FL�<�Ƌ�Gd��W��;F.��DC�F�<�6D�
8n��I�\���^b`C�	�!�:}�weY�A!��ٵ�?;G~B�i�C�BVER`+�C�9��|�c"$D�L9t)�:�(ě���l�@ȕ�#D�()&̓�?����"]lg`�:�o>D���`oQ�mi@);�Z�'&��X�e;D��6N�K;��*���
X5��H�9D��!6����9���(]�!Q��"D�P�ԥQf��t��0�i�Fh5D�d!�+�(�t.U�ky�d�a�3D�8kB,�B`��(W��8O�����O3D�X��� b���hҒeW��B��2D��S(E�m#Xx�� �3l"|�F-5D�� ���K�l$�6�Z�>0X��.D����)�9���8���2~\P��g7D�*� r���d��i+�1�!1D�(iƭ� z�����c�0�� �o"D�D��� t�H����}l��`G ?D��yU _6G斱�qg�W�`@�b�<D���O�y�y�0f��R�z7�;D�X:���2]6a(W�P��W$D�l�(ĵt�t��m�.���"D���(����C_4F`7 D�$ 5f�2����CHЋ�T��B�)D�DX!�T�Y�!&��P��X�`'D��t�t#���Ռ
����A�#D�H�4H�8%��	��5����.'D�,b�����4���iB
8!�� ��%D�hCücT6]X�K
�L�Zׂ#D�� �P�b��>^��V�x&�-�R"OJa��G
p����E����"O�$p��ɭr�"1����eR�M
"O�B����$�`6F��RAR�%"O�P�$G�;�x�����;�=��"O4�h��J�)-hp�f @)�r<��"OJ�x2�ϔ9Ѿl�!A	�!�t"O�K���.~�Da�n[���1"O��*���0|�6���#�"O`���8��}qcKc͘Q�%"O��HV�ҧ�0��B��:<�""O���e��C�&����d�
tɱ"O.�����?*ġ�� �\��P�"O<�(2��h]�A�g��6�����"O��ॊ��M���%�2�n�*�"Of�b����J�e�����	�0}J�"O�f��Ha���d�Wp��P�"O8��@+P�,�
����C�a�<��B"O ���]���f�l��"O��*�`� r:N�����5G�}��"Of]a�.��a|��I���E-r�"O̱����3D�AB7DF��`�"Of�����##����D��)�m��"O�@�@cL�"���S�B��Zk��y!"O����h�$H�qb!�N�&Fʅ�"O��Õ/D�¤9�Ѡ!4�@Z"O��+�J ���h3bhȒe2�� "Ox �1תgF��0��>V��9iW"O��c�·�x���ߘDF�3�"O����c��aChiB'�ֱq'�X�"O�D*�fƒ7�d
e��H~��!"Oz낀�/H��)��0��"O~P@!�:��hU���F�ЩPv"O���$��5� �`c�
�����"OP1��@Y����3���2mx e"OP�x�T(TQVMP�iμˡ"O�	i�B��
�#Q���@���"O�0`�o��W�P�!�l�#*�^�Ӡ"Ov|i$Ƅ }����W��+Ny��r�"O�8�2i��Y��HQ��$a���"O�i��@=.��`j �ѾbO�@bC"OV��F�S�8�-���M�(Mv��""Ox$H���w|LR�/,а�`"OBDSm�*HT<UH��ߌZ2$ �"O^���-G�W�@ ��\�f�ɵ"O����΂P�a#���/u�FY�R"O@|����!�m`g�o�!�5"O3�c(j��D-H�DTyd"O�=XW����t�"Ǚ?�b܁U"O$�;	�O�޽����i��a�3"O����EAR�`�b�:�zh�"O��3�&b�!
�$˗]l��H�"O,pi�m@�8Œ��cT(xO�陳"OƼj��`8T [�!0L�5Q"O�P�'��\)H`bB�FFd,1"O�9ZP"��7�p��4d�q;~��"Oz�(���+t��֣�%u����"O�1�p���n(��@'F��AȒ"O��[��Ȣ ��m����4��ږ"O�yi���&~u��jC���W���)1"O�CV���@����BD&5�l"O�$#��՜hO8�(�A��cj��r�"O��c��Ϻm'X�yr�O�QY�H��"O����ƾ>�8���ރCBlq"O� R�@(��Y����q��-ph���"O*�J�#V�S��L�VnM>�f9�`"O����{�
u[�Y�2�$уP"O�(�`��t�����o�Lǔ�H"O���w�4qp:�"eήhĄ��"O��	#���P%@�ہ�W>i&�艃"O��zs�_(spT�i5 �t�"O�pIr��T�� ቐD�|�f"O���_�H4�U	�`U�^�~��"OmcA(G-��r�Z7U��]�"O:��I$z�1p�Z�B�T�W"Oez&@ƶM62���,x��)�"O�!�˩q����sg�'��{�"O�-����'��s憑�k��4�"O�52Ѯ�&xp4�6�мK�‒e"O����LX�Y��)P�dC���p!"OV����Wu��BT�&h
��7"OT�2�KΛu���!w�IAj�c"O�`��+�/R���#,&� �f"Ǫ�AO8(�]���5`����"O�%;���a�0ݐ��
]�	9�"O:a�7�*~�ґS�i>�(
�"OB�{�/�/� ���%J>��r"O,�S�ņ,���+ǉ�y:~̀"O�%�2KK�3A��x')�N��3"O m[DEѓ5´��聚�
` �"O0\�&��1gֽ32�ѳ(r���"O��*�f� ��u����*\$ҳ"O�I�wO�	P�R�Fڴ*���"O��Sd�L�A�fmʱd[��� S"O��9�̛6O�&x���#�4�S"O����3l�D��R"U�B���"Or5�[�w-R2BA^/ƾ�h"O@�*#jN:6�Qo�);��"O��.�_,��I��.���"O�,kS��]T�H�������"O|Th4fȞ���S���GȔ���"O���B�Y@O�Y����kR|d�3"O���H��R �� A@\�u"O�t $D��Uz��!W���A"OE�!�V�H����7E�v�r"O��h�*U.��!�(��"O��!�鄗2dܘ�B�D!�j�#"O0@�x�6\�V=!�m�"O�)JVDA`GB���ң.o،S7"OhuP�E/F�1r�j��)Vґ�"O�ͺB
�)�����G� �.@p4"O�,�eC?%�x�\�kӮ��"Oթ�%��N)p�s#��J�0}#Q"O��#��� x�|�{`ҟjEh4#'"O���c�X֎@�%�T��zi�#"O�H2�+�9)I�%��aĖ9S"OF=(�肃3.q��Y�'[f�(a"O��v��QT(L�!��@�Byr�"OF1� �O�� w�ʀ.���"OX����D���A0��[
F�y�"OV}2�h٣I���st>r�AU"O�P�BC�7&5�&#/�p��"OhU@ *P�43@-p�'W�+��Q�"Ob�B�O�A9���&���G"Oα1�JÅ>>��k1�^�}���"O���Hģ88���s�h�}{�"O-ѣM�)7k�ep��^�1��A��"Ot[��. �$�e�4T 8�5"O� ���K�"dJ��b�"�60�"O�]�Վ�6�M��	��oHi�"O����E=8�\�p��U9�$"q"O0��R�}�p!V읿�P5��"O��q��J�c��t��1"OV� 
�C���3��=C���T"O��p�Bw �� �u�H��a"O��{���\^h�'��?�6Ak$"O��c��]<2ݼ�� c�> z�%"OTMs5kțr��D2$!�8C`�l""O�@ҘZwP{a	�\���V"O:\��� *+_B�Y��)��"OV��/E�\xRi��,�3}P���"Oޠ�4@� m	j������h�"OĀ�
���ua���\#�7"O�3d�#��2�2Z�a�"O*�hb� �"���!G�7V���"O^p��ެn�|��FO�wdT��"O�ڀa3mb=KsH4RZ]3e"O���DCʷvW��H��,M8�R2"O�e���ҰF��S�~�Y��"O���6��V���@�*�ܠS�"O��� ЂJ�x*u \\�\��"O�y�af)hD�7Itx�q��)�y�c��H4���V�m]�E��y��+��}bs�N�'oT�á��y�`��p�����@�%X�y���,�y�C!E?�Y�jFڐڵӇ�yi�?ʴи��0E�|Es��&�y�O_��l��đ=�Jp2��?�yR�)�R��Ɲ�0��k�S��y�B�m�:�K�GR�z �+Á�y���De8e��N%?��B"����y�J݁����ٯ9�lS�d�3�yRګ8���c`Hׯ0���E��+�y��w��	�+�:%Pt���"��y2�@ D΀�@�Y�0t���߲�yBD�H)�$3uB�I���h7���yRbv*��Pt1|���A �y�`�)7v��m�^�]�W.�"�y��ߗ.Dމ����Xd&�9rj��y�e�A�zAZ�)+H�𳡠��y��Z��������;��yRk@6�y�б	EZ��� M
�����y�Ą9.|%�@W����`0�y2�_���y�e�Ǆh�0����y��M�4���C`o��4��m�0�y�E�9U�f���	ջ��X� ���yd\j��M��hH'����gA�2�y"��	V.��K��U@�'���y��ǎ"F��Qg��0C�Ms��E��y2�
YBQ���1��L��}��'$f����7x�}�"a�����'�&��7@	$i4邱舟_c~�z�'^��ɕ*�.a � ��ٿUl���'��}#�(�XތiR��T(Fb�Q�'���9R���0["��!�$4�$��' \� �:C0\��.��'�l�'�L��b�	BU���׃�)j�D�'9X)yr#`�8=b�j�n�1
�'D� C�5K���r1�z<� 
�'aD���	2ȔQhP��|z�8��'	�tʆ+#*����L������'7`����t��H0$m�#=�,��� ڬ��"˕^��aF�!J@��'"O�����*c�%Qc���Y�~���"O����GW$@,u�W�5{��$ p"Of �&�A(~"�UH���$V���3c"O���O��i�l�@�l�`"O�I��JQ�a���uF-pҒ��7"O<� ��r�	bSHA�.�f���"O��B��Ԣ�@��,N�����"O�yh ��m2�1���*����"O�	{�_Zڞ\�U��).�$H�p"O@�9�m�;�L�B��!k�q�"O�u�P
;H�����JU1SmL,�"O pH��Q�!9n�˕�);NX�Cs"OptRr�@:. ��r,�3y]h�"O�)�Cʰ: �!��N;+D�-0@"O
p�6#�;]���@R+R5x@��Qe"O4�`�\�20mRS[�s;jy�"Od}���O�&H����ηc5�ԉ�"O�e�P">0���4�Y/+\�g"Ob )wԝ0[45��(�
���r"O�-���9:�����&ʠ�r��"O�)�����
�5X��}𖋋��PyB͍4G�l�pH`�(C�Ɋj�<IP��t��p��I�\媓J�O�<Ab�?g�2��G�����2�IL�<ᣦ�)�"� �CSvT��*�$�F�<�d?x�4 U��n5��
E�<i׈R��pȓA4*,ธ�(�}�<��_�&6����})��I2��|�<A��D9FL�0�fۂI�h�T��t�<)S(wIk�d�&��P�U4�C䉐kr(��䫝=� i@d�s(�C�ɹ{᚝�$�N����#X�
B�ɱ9��f�dIB�� �0��'"O �a(C j�Te��e̯arё�"O�(� F�N�`�vŏ2S�.40�"Oz-��B�0��\X1O��y�lA��"O��si�E�*i�.��~}v�("O��R��5�J�9��E�N^b�b"Ol�#4gS�3�\B+S�h����"O��1�g�*��!�aD_�)O� ��"Om`
T�Y�bpS �� 8��� �"O
�Q���>=�>�:TO�P
��T"O���$�؜�^�n8���"O��! Aɜ������B�,�*�"Oj��	�B%Ӵ_5�]YA��%!�DT�+��m��G��!x��[�+D�'�!��S9V`2��`J��%k���Q<�!�$A�)�h�*� ̳,jD�!�Ҝ�!�$�.dD,� #�e�ƈ ����K�!�dژF��Ċ���Ƽˣ�S>�!�䌺l�b�j�A��,XB5��Yp!�dɓiģ���ؐWb�,V!�͹1��!tN��G��P�K15i!�r�plP��G�u*��H��O�Z�!��L�1HA�B�D*�q�S�!�ݎ=�f���A��C  ��W�!򤟚5��ԫ�@�q��}H���,�!��l�E�Ɓ�"g�~���ȑ}!�� ��=5�Șr�� ���5_!򤑎*/ -9F"G>Uy��4F�'@!�$	}ޤY2'ͅ"�h�a��\2!�䇥��i��Gj�4��v%P�L�!�մIY�4� z�����G�;�!�� �K�@�8���Z�ĎWB<q��"O6�ѰJ[�� �S!nDb����"O*Eѣ�L�g�M�"&���F"O�LkubB,\
x�a�@��b��9�A"O��1��E]҈26.-,xhx;"O^��
�Z@�n3
�H�U"O�m) �>
骘!�HP�q��s"O��۲��#�t�DE̥1�FX3�"O����O�0���8�E�;�^��e"Ox���S$:IA�k�*C{jP!R"O\�S���K<�,b��D�<g�0"OH)q ��jL����G>"%"OH� ���a�yV�ڦe6F]�"OȘ���"/o�(Zg
�$B�Y�"O
�aUA'��I!ě<g)���"OJ�`��Z���YKCa�U�63D�@�p�T+
&�b�៏��ݠ4�1D��C�m�Vi���*�,�@Zse3D��5�̊�ti�w�;lx���;D�,�u���9%�[f�ҦN�
��l9D��Pf$�2@��+b��]���5F7D�L�wLǉi���"��B�oX�	���1D�$��C.]��l��  ��V!��<D�h��mF�	�l�7�t���E9D��8cA 7��}�b��\.��K!D�H �`�Lx��v�߸9Mj5:��"D��d�Xeu�4H��_/F}2"O+D��� ���VцU�#�_l�2��u�'D���3+�\����N� 1@0���K2D�X���(nFA�s�@
zL¸�C�0D���u�Q=����CO�%�lف�2D�"@��}���)&��rR�<�E�2D�\��+E�rB� ��D�Vs��r��$D�<P���4+��R&��-]@�"i?D���� ]��1��+ʻS��r�*D��2׆��f�p)ʣ6mau�<D�(��h+`aH�S�=2 �£�'D��*�ޤ,�X���&{�$�g�&D��
�2M�1�'g��b�D��a$D���s��l(θ�R�ˢk|4 ��K"D���f�%���U-H�WU��y3�%D�p $@"v�&E���[ 7*ԅ� #D��jbS6���9O����1`sH;D�H҆m�^A�	���>#&�MAG�8D�8�3�ׁm�i�Bş C\���n6D��k¿4Ő0�V��!Vd��d�(D����L�o�V�31��
Qq
I�1�&D��jD��X�����.
�	�)#D��1-O	h-`�ZVC�'��A�,D��	Įީ>W  �uE1�(탑�6D��3����u���D�Ƹ�ӣ&D�����{|6����=u�p�g$D�\Be�AR6y{A��]cx�a� D��!Ì��=Fй���)6�Ʉ�>D� I���c�J��̑9$��t`;D�X:tD�1J���A�"dDCGB5D�t�d䊲�@9*e��
`�b�4D�C����b�B�8���	.Б�h-D����#�x	�����iI,D�tQ�d�<t)���!��4~0)�r�4D��3&�]�]-b��%㇭�0�1D��i4�ݬ8�
��B�A"i��!D�d�W�V�J�	c�A�eTBP�7�>D�)���9���#���+�@�9�7D�� �&�'d�Miդ:3�P#%"ORa�^�a�x�8�ɉz'�ɰ�"O@R���"^u�\�$�&k#���"Ouy�M��w� Ʀ�!!�u@R"O,�[A�P�R���+�*
E���"O��Ig�ŭ��iy&�G4K`ĠG"O����7����E@FLY2"O�����ڑ}�8�������\�"O�(3��7&���ǌ�r" ��"O��:��RGu���Q�Z�C���7"O�T%ș�?^�u�U�q�>�s�"Oi�5��,[�ѣ0)̬=���"O:�ɃgN9��I�b�8F�t���"O� �S�f��H���ۍJ�¨��"O��sKL�xH�س�h�5���KV"O4��w��D�JqUn55XLYP�"OҘ�'i^�4���e.C�@!v"OP-�v�v��GȚ�'����g"O��ӆ��'9�)T'ZZ}xx��"O��·�G4C:l�
��Õ\^��v"O:��T���T,��bݖvP���"O�<	g&����RA�"MJ$E��"O�yà�����*W���-�,=�w"OXXفE�}���6s�<��"O(����8ܤ	be	2_l�0��"O@��c.�+$<�ZT�[/H�"O��c���!B�6-���u���*�"O2I�G���I���ߎb��*�"O�h9����x�p�+�/�$��"O0� �̍�v��zAO-&�E2�"O���	(5I␘e�O�^�����'"
]{u@5	hU6 H�E В�'	�˦�M�o"�#�J"?}���'HRT��*U(�n�y��ّ
=��J�'7d�"&@')�z� a�����r�'p����)ϐ�{7#̗y�H+�'De��`��Th�XS�<h8�':�+!�M�Q��������ɳ�'0"񁐝t�&�$�@�	�	�
�'��EBWnłD(̠�eK�Ql�,�	�'(XU��J �c�C'愯IB��':uggֈxF�Y�WdV@���
�'S�	�H$P�Uڗ��#�6���'��,����F/$�Aǁ	�1����'z�a�b�=rL��X�뗟f�B���'����1�H�W����RGQ�`/�i��'5�\Q�,��	C���C�f��"O�H���T�ٲ%"�*�a��9�y�94�LH�*T��$i�%��y�f_'P�N��W��O�T�#��y�O	�tж@QW������DE,�
�'lx�a@*F��c�B#<�<�	�'C2SP��<~�a���3'��	�'|�䡆G�K|~�B(� 	�'���	@�;�pA�
�՚	�'BD,+Dc�0i�����ܺ��A��'ݜĀ$��~����IN�

P�'[�R��_�P�J�!@.��^�C
�'�(�f�xEQ{7��;�
xE"O`�1��K�H��Ԙ��X�� ]3&"O��2�Eҝ����%��)zf�3�"O���_1.��@��JU�-y�"O���lGI,z��D`Swݒ���"O�5�u�V<8�tj��@&�\*�"O� r�Q�&�ps`i(vi�)Rh�z7"Ov��$��%(Hp��uI
��(�"O@�9�퉬���hWi��I�*y�V"Ot`S� �� o:J��1���)D��p�� f��=��*�_���`B�&D�Pi�ۇP��`'O��d%�0��#D�\�7+ۢB�&ă��B k���"D�P:U��*s��  B�N��yZR�<D��
�
�����k/�\���;C:D���P���-Z%�8(vp��4D�x��U���Y�L�L3�J�L0D�PB���f(�P��ܵ1�hl��k,D���bL�s��*��Z	J����+D��S��#��d��z������/D� �'�Ɨ�x�C���e
�|/D��J'�b�dH��� a"�@ش&.D�L:���$)��R��F�h�Xb��7D�4b#�+5/�����3脄aB7D��:�"ɦfn*��r�µ0��8��(D�ȁ�� �e�Aˑ̖���e1D�$� 	�.V���GGӇ�ʑX��/D��8�H�ܸ����Q;��S�"D�Đ���N��3�ϳy��;�i,D�<y#,M��Af�6�>��2�%D��	D`	x�i0#�G:�j�S�>D�쑱˚* D@fO��_�Ո�;D�h�g�	}�8�Q�ܻc����0g7D��S��q��+ǆH.q����4D���c�Ά�TE���)8�`�n D��KgQ�|�&��&d�M�Nȡ$�>D�H�@K�Wr���IH�i��<D�X��#L�L���0_jB�y4�?D�l9 ��/},5p�O~v�@i3�=D���	��PPy�g�;��=D� b��1���a��՜PbfT"'D�d�N̜d!6$X�O�)adH�5�#D�p����n���L�w��� �"D����0Gu�P���YH����'=D��I�M�"��� U ��������9D��H+E5n�a����Ը���;D��k��%
�����Ѿl����d=D�LcUU�bcS�M0@�F<D��rp��x?nЋ� 
�E'���O&D���3���~�$9xc)�(u��� a.D��A1l�_���0`%%A�ۣc,D�,�#	ҽ6\��CZ� ���K��+D�<�+���(�����V�^��Da)D�8�`����rVL�g��$��-<D���$�L�|ޡkl
6|��Pi��:D�����Z�ؤ�cNȡ,���E<D��+���G�ř�O�w���h��?D���*ˠF��-CQIM:&n���J<D�;�
\9���a�˝e�4�#B+5D��!�+:3p���Ht��h��k/D�b"��H,Z���Ƽ@=�I��)D�TKD�ġT��LrC�O�����'D�L��b�Z�|u2�JZ��5�)D�,{lX;~ �4>�P�� =D�$i��N��Z���ilC,�Y�K?D���$U�C��m!��@4q��y�VK2D��9�-�32H�*4�T(?�ڡq��1D���q螲MhY�r�M(%��S�2D�h�,Ϊ'��T��ˋ2Ѭ�ɑ�1D�8�B��*@׎D��c$U>�L�4D�� �h(69H�}!��˼	'�y0R"O�!����	: 3G��J ^"�"O��;�z�x�3%Y�%*>�+�"Oȁ�͂jDprn�p4]kG"O����L��"�_(W��(!"OPu�e`���B�fF_�H7��$"O�Y��K��Yb�J�	0j�0"O�)�Ƀh�ν:��I�*&HK�"O�IR�"��eт��a��_�$��a�x��'�J8�4���a��d�+Ur�U��'��5���T�G�P��;�'j��̓L�H(R��7K|5ʏ}��)�iَ��@���ޭ},$Qp�\�*�I{��H�,鐲kYm\��R"y/�YS"O�6+�@�}���V�4���"O���1OLyYp�h4�.~��rb"O� [1�)�j�q`	)���"O����ق(#^	�gB�BLv�Q"O�} ��/WzrMjD��8�$S�'h���O:Q�jL@��0b�8;����"O��XG�U�$6ՑRaI$'�(�("O�$#��]�F ���[�"OB���R�b-i��?���'��'�2��,�|3��=D3��"���y�J�3�P"�3G��� o�yA�_l[�O�'>��t:�	���<���$�ly`�#я�M{Ha��,8!��-{�L��
KHԒv�X!�䜓8�m��發:D�m��-�e�qOp��DxZj1#�V�x��+�>n�!�DN;~<�-y4�?��@���M�&D!��
ݼ��aE��&��嫗�I!��0	�z��)zɐT�4�<��G{ʟ|հUkL$8{�Xʅ�����)[�"O�Mh��Ú���,�x�氚�i��O��)��QzUO�<�
X�'!u�,��b`5�ث�BG3J0L�'H��)�����.B4p�!�D� A�尶��ʩ��F;a�a|�|BΛrd�1��,�=2��
�e�#�y�Gפl�E2�䂩*J��e`ɉ�y��@<�q9�KIh�����y�H�rd�f��r6L��>1�O�s�í@��|��m�H�@�"O۠dG�h�L;���Z�@��"On8Ѱ�X.[��ɑg��8o%&�[�"O������H�ly�f�?$0|�P"O���)H�:����AcF�v.帑"OV��B�)	�¹��t$8|Z�"OB���M�D7���@�&	)�"O:`#b��9e^�1GM�6�P�b"O�!�w����!.��Q-M)��
O��0�k�5��E�
�[3�Y��'���I?:�"U��/\5PD��	5)��FzP�=E��'a�;V�	4�&���-�<b`��
�'�J��K15פ��4�G%/#�|�
�'s�!���5Y���L�pb٫�'^��"d�+N���X2
\5�:��'�Āe�U�m}NѠ��+��J��4�'I�n�r���:w��c܇C���ȓ�z]�S.I�J���P���ys ��z;�Ւ�j4o���p���x���	Ӧ��U���Zj����b_��Y���N�A8�J � a�W�X�%D���fm3D��gǕ�)6Jm�ċ�*���s�M>D�� ��b��pa2e� %�+Qx���"O섊%.��%3t�{�C�7Ԙx�G"O|ՠ6 �8f�V�16�CP˖���i�ў"~n+g�l+�@���fH�`Ō;+����$*񤕪f�@�
f��q�lb��O�}`Z�j���v��?9����E��Ip1� �� �/`�<i��!���r�㏔wo�LS��\?I��'�X�[c��:��2,��]q�|��'dy�U�
J�:!�3��Wbnȫ
�'�2�ceF�ɂ!��=��R�'H|��E�B#~�1�h�0�DB��D*�����\/2��$�)~Hy�ȓ2��)�4 ܛK��R#��
&">D�<۲K�T0���D� G�8���	�<!��ڠ�R��1� �p� }�b��'<�'�ў���&��kt�V�E u����C[�B�ɉ/��H��NĞ	�x����>VB�	p"�0	�x���$,Q.ZC�	�*n�I��Z�Q
X�4��Ą�ɧ[����ʚ'yx"��3G֐����G{J?QkdN�O�=��ϏKI>k�-D�܀A�2^˨���͈;":ɚ�1�$7�O6���W:?���CK��2��p��"O\���A�*r,s��� F�6X�'O!��[�Y�6` q�ɱ#�������J���G��j�"��X�H�z��Q)�c�0�yB�æ@�� ���pr�tQ6��&�y�)J;x�(tܚk�$`��y����މ9@Ɉf�Z���8�O�}{� ���k�̲+��R�"O�ܹ`d��uJ``�P֤)I"ONMb"�Ɨ�24G�E����1��\>��@v��`A��P�����?D���h�R/.���D؎H��\�`�*ʓ�hO��h (�k?c7pU8w
�F�|B�IA����R�*>cn�sS�C=]��O���]�s���6o<�J5�&�4(�!��
����@��� u��Xxׯ�,"!�$�pbf���)@�(��ձrA�ў��#2(���Y?*���Z�L_�B䉦�[t!F����Xv��
�>|Oc�t��.C�T�6�B�U<r��}���=�O �I�����I�>2���h-E]�u��'D  X���*�A@ש�/*��[����4לY{�G�5���6��F"Q�XG{*�Ȉ��[k���3nO 6�T
�Z��O���'k-J�&Y7pv�J�P�=,����~`���ns�,*�J�:^u�a�ȓ^��4pw�L�go�X�ttE�=I	ۓHڈ9@��|n��#E�7���"���kF�I�S��m��A`Ȥ�ȓJ�#�m�#�
	�C"�z��=��N��\����x��ݙd�)
]��5n�y
���u��y��[�P�(��E��05��"(���W�F� 	�ȓ`D�z֭�PH�a�R�H����74tX��Q�<hn��
�#�������)�S�S+E$��:�;N6��s!��D��C�I����[�%�+{��*qE�P��C�	�@��])�(�)R�yGibĦC䉬L"�X�p��?���rV�
3f7M�<����)�|٪x F4�6M�.��qH!��6L%b����>�B}P�L1�!��+'xD�hE1��ɣ�k�,V�!�� ~�����	H=2nD&>Z*�P�"O����A	.i򡀶�OmC�A���'ў�[ץÙof�P+.ەt�z��"D�dr���<	��:
��{�uzqdk���>I���O�,��ɃKg�񩆜0�0��V"O4u��Ɓ )�4r�����y��"O��ӶMK�Ml�yh���w��2"O���d\7un�E3���2=ɤIj�"O�I3�AL�T��F�!r��y"O�Z6��)f���P��Z9����"O�,K�
F�Q]p�C!��D��ٙ�"O4�1/ƭd�T8cf�WXp�'"O���h��U�A�Z��T�"O��2b�C�]e��#�c��u�E�&"Od�F�PE���S �-pҕ#t"O����*@n(@E��1u�����"Ol�tc�)Ϝ� &S�_Sje"r"O�L�$�*k��.M�E�ȅY�"OL��d�zG�"�NԿ���E"O0\�'
\�;�l8""��3���Qq"O����ڔ��' Y <LM "OR��3KS� &v�x0Ac��[�"Oh	Ye���>t��* ,:��S"O����<�l�
����?�����"O��ƭW�,�Μ���X�I�"l
�"Oh�@2f	.[q��kբ_�5�:��"O�\�cC=�~1���M�����"Ox�P�,7��H��5L��%�"O���u.�K�  0tb���6V�yB����|񓯟�T�\-c��
��y"�Э:�&�k寀�@�Rt𳠒 �y2� 
 -��Ҷ���Dm��ҧ� �y"D�T���
Q�'/��}�����y��\���	���K�Vy� �P��y�L4J��1��>M�pz��,�yb 9�
��f��=IUвH��y������2!�mk3g���y�d�{������8�۵���yB��.ƔI�f�=���S���ybA�/gT<bq�T�rM�����y&
�/am��� ^�$���y" ؟��uH���.����a��yr���s���b�؏%3��C����yBM�z��D��_� �h��6�G�y���%��e:��Ok�(��.�2C>u!r��%�0?���m����1� �{i�I��#�[�<��#"hw�M�,L!U@�Xf�T�<��+E�E�%��4(���p4,�Y�<��NX�T�	{���'#Đ�A��b�<	��ܒUS򵹵�"Whx�2Ю�u�<b�)P����.ݱN46�ҀOv�<�󋇇r<���c���'[$��@�[U�<y�E���� �@�wnJ�� �WR�<Y��U�p���Q�����.M'J�k�<A��WHFM�g�`�����.Uf�<Q�j�.D��{ 		;a_�����h�<a�mɥg
t�����9=Pp�d��m�<�EBܬUf�t;�Z,S��g�<i�� X ����
�z<�X��c�<ɧ���V��!9��9���F	1T�p@�*W��u�0f߅OK~��":D�(@ԥ�=J.ݙ�M��&T�D 9D�d���	�֘�a[*�X\��&6D�h��o�.K��5����]��uɢi)D�� m`¦��`Z K�	2���"OL��t��8i�F}��	őL��C"O�{QAӞS/�qTgU$mB�0�"O�0��ɂv}���'4|�3"O$�07&�3T�S������F"O*i
� �=,�ĵP�	OH��	pp"O|�����eҠZ��ϰU�e�V"OP��ᇙ`H.�"�	~�Ri�"O��"��12"�hū�Dِ�"O�ȵ�S*[��iP�D��\��!9�"O$�
%h��2��8�{�h��"O��eg�,@v�B6�# � ��"O6�a��W3~���&��F�$�"OZH���\'���J�n�=e�:�s"ODs��O� C��`�l�8V�.p��"O~%)w� ��l�[3H�jY�"O2��G]S$YapG�FZ$�'"O��#Q+��KϜ�;'@L����p�"OR᳇@}�z(�s��
��"B"OXq��j�9�E�b	b�B%��"O�×Fg �͠&.Z�:���B
�'�N�`����Qk',E�m���0,O2�Bf��0��=�t`�)`Q��7(��s��^8���6�"{.H� L�q��-�S,��3a�歚�R~!�Da�����aS0[	h$���Le�������h��IG��f�'��KӃ�5�d,��@K�F��ȓY��`�(K�=#�]����{�~���!Y	E��(�c"�H���,�g?�Ec��d���qf&/����
U�<�F��3���H#�����۟0�`�[;����Ab
p�ay�@ő8n�au*02���4M���=	ft��a���� t�d��EW�0<8�ywF�(��}Q��6�Px­W���(�DD-4જD�Ʉ��'&�S���5[)|l Bb���q�d�J�'ξ(;CdܧY�[g"OL��Gl�!pF.�^���Vbğ!jF�����vK8��c�-�?	��>� ��`�vH�����]� ���m�<�ת�,�@��qO�<[m����_¦���%�z2�����"����㉌+ S�AG+Ӓ���/����$��^p�9�2Ő�)F��
��AWj����E�'P� @�[��C� jqN�yM�#��l�	ߓ3��b�Dڧ$%9��a�:7����}"��'�N�Õ�W��X�<���초j��)'�5s���<R�sa
*rQ~}�R�Oj�E��O&l�7k�భ)$���"��y&"O$AfDE����0��ZJY ��'DRT����'X��EX�tĭ�?KXܒ���6m� gm)|O�d��f�!rјl+��T�Og��a`
@����J@M-q+Jl��'�2�����VT |�hf�|�����P�q�E�� r���?e�d�Z@���dE��qQD�$� D����V/`�G�CY�v�P��/?�l��Q��6}v<ҧ��҅��<�b�a��6e9fl�y��v���N~$�9�D� ��\;t>�y�ۓ�a"��;�h@��3G1ȵ�ȓ&�,9��˚?�\��٩z��Q��>�J!��6��F�́VQ^`��?�d(5�(�Z�3������B ��K }H�	4�:pd�P��jv\�
"Gݬ �0p�;U�RA�ȓ9�A�h��Z��t�פ3P!"M�����P��b(XC�=�x�ȓg^N52@KģH�B�b��	k����ȓ<�ش�r�֟^t��r��P�Bĵ�ȓI��� ����N
Veڹr���	�ԕR��>jKn�Ѡ�ɰ}����~"8La���$��X9UD�-U�(�ȓ��ǉ-�Fi�
���S�? ��8�]��f��dF3R��x�"O�z��U�hE�:"��u�T��"O�uyQj�%c��n%���;E"O�<8�L��B�r���G���"P"O҈���� �8���2�4��"O�8�C#�7l��ۧ�¡�D�xV"O��QU�>:��x�o�>�z�85"O܅K�����@^�Pd�|�D"O�Y!���1~Z�Iq���P��u��"O�ث3摽f��0iU	Ԛ|�.���"O�ha�o.�xq�脝p2�H"O���䎑���D�?)��H"O��cD�R������X�
��a�"O4�W�U�pt�AuBO�u�PqF"OXLa�`R�I��(2daF.2��@"O`Dѐ��U�p�*4��@l^�z�"O|��6��05"8�1��ʜH��	�"O�tK�<xnn`id䟙 r��u"O�T#�`U�,�es�-L=l ��7"O��)���2,w�I �mTyd�}�1"O���D��\��a��UR��{�"O�x��`_,Z38��Q�R���p"OB�3P��,;<P�v�A�[��r%"OvŉA/%� ��<G���"O~��  F��m%X���[�"OT$�C!Y \'��+���f��q�'~�hכ|r�û7X�u)vh�)UVP��W�y�㚉7����AH.{�ػ�'͒��z�ă�g-�)��'�N{`�χIt��biй&�$C�I(5��U8� :2x��2����$�J�{B�	L���+<>|*rK�/
�tqw�N�y�|a�ƓMk��ȧC�;5b� ��_=O׊�z�&	y�8��D[6tv�R�⑜O���g_1��y�J��%���u�P cȰmk��A1� �TM"D��9���#���n�-@T$��%�,�$ެCS*���{��4ښIԬ@�6�ڙN0LE�	�0�yBh֨~@L@���;��z���%9��O�5��3?���KA�$���c~�y0���\�<��'�l���"rMHZ�ȱ�c Y�<i�$F����ԡ�x�j�{7��Z��d�?i�O�#dh�Bֈܷb�v�;A�LV�<	�R>;DbhPև��@��Q#�SM̓�hO1��ՊwΦk��Ať]�M�	�"O�#@ə�[>�"��y�Ly�"O��
g��'c�\JT#� ,ؤA�"O��
���1��-'k���w"O����6)�Ȉan�7nj]��"O�@g�C]��l��E�hL�d"O���n���4�J�'�&Eh�"O�t�A&M��үV #�:ՋW"Oƅ����8R��c�I�)���p�"O04��O̠M�\D�2`P�<aQV"Od�gB!r�.|�#-V�"h�4"O�8R�6X��0d��f"��"OX���;lۦ(A�ڍ@@��c"O`�[��Dq0<�)��܄u<X�C"O��7Ǎt��17�J�@�d"O�p�V �:*vV���A۵g����"O�9B���?e-<�����BW�As�"O���Ca
�.~���S�R�;p"O����R�KalI!rl ������"OD��/݆q<�`����\���3"O2i#S�,+|5���-��\bU"O�����!?�F1v��5J�~�R�"O� .�u��|6���7*W��j��$"Orp�e!��U#����C���q�"O�� e��1\F|��h�Y�6!B'"OZ\�C����H�\R,���"Ot���)M��2�bnN��"O�@��$=Ƽ��=V>�`B�"O��Yda�9����jM�aؒ4"Oڤk��4���дp
M1�"Opl�L��uWhB�6g[��"O�x���H���͂��V�cޡ��"OZ�Q��L�6ZN�#R&#]<�q3"O��c�M�&.�QI�ř `Mlq�"O�
�mU;M����۽<0�j�"O𽲷Ǌ	���`,{#r�G"O��ٴ�)����9+ر�G"O��h��/_`�Ku����,0�"O�(��.8	-`e�[�-��Х"O�H�"N7d��x���,�5�b"O�i9�&�78����6 �|��7"O��j ��4�εɆ�^$"ЦB�"O����oH�W��ѓ���!a1�1�"Of�9� �	ci8e�၀4Hf��"O�=y6�6�|2ҀM5$~d[C"Od\A��"x��&o\*�"O0I#c�ҬQz�	�w���2"Ol�`�!�D�j�c�A�] g"OҔ)#iGlJ%��k=�[2"O��k1/H+4-"9�`b,tZB�"OJ��������1"�(x�A�"O^�
v�(f*�Z �ɤj��X	%"O���.�j�,�����$8�d*p"O���kH�{OLm���D�?�`KT"O��:�h�<,��:�iD�/��l`�"OU�ю߈p8�x��iQ�k��bB"O��D�=�V眱o���5"O���E͛<�4�ㆉ��`w"O(�
(f��A�qd��.^���w"O�pJ�N��^��YQL��'E,U�"OP��`�H�Z4cGj :c"B���"O���炈"R{N	pςx��h1�"Ot}#�כ8vq8��S�@�"O�	�ͽ|��T�ҮGMK$H�"O��9gmѼ\MP4��j��[L h�"Oti�í]F�����@�76Ha(�"O@|{7�Z�kc:!si�s�vE#�"O
t��`�+x6�@jb��!{�,9I"O�y�2�C�"7:��@�H�m���A"O �p7���7�x`CᝃrD�dٲ"O]zP���R����G=t���"OHÐa����L��"Iؒ"Oh�k�.L}ܠ�\	 �qB"O!��a�/�dth��X-b%����"Or�!���6�1�=t&8�rq"O��!-���|���*'��"O��i�A4\.����t�����o�<����J	B�	'I̕QGVp���g�<�!_&Y/�IPE 	�}�@�E�z�<q��c��HP3�*?�-�El�u�<Q��.$Ȃ �8�j@�f�[w�<�f�)!�" @Q
�{B�;Ês�<�t�/_oZ�#�Aا
'�#��q�<ѭ�8h�C���"u2x��)�f�<I���)���G#-
Cg�<��]��@"�����P�b)Gv�<� N�fa��A��\�C8J� �11"O��Y�͉��a��
w��xz�"O����0,z��^b�"= �"O�m{vg�� X�9aW����P�"O��S���.mx��e�!,��"Or� A.*��9Fc�)I�5i"O�Y� �0��ʇ�B�x���"�"O�1��F�'�"]��q�6k#D�P�g��)�f��D;_��@SD�>D� qG/f�l���f���L{w�>D��I����!��l���W�MJ���
;D���0C�3>,a�dkȧ2�<�R��"D��X�2� �ې�J7_\$H��-!D�����ʖTX�@R�ɉ9R��K��:D�<�gJ�=
 �3� ��^=�5���.D�X��䞧�.��7�ǡ�,��rn#D��5�T�,h2AEW�,nM��!D��
�k��3�������,��Df>D�L�5I�,�v���#ɾA��T��+D����i�`&�:@L��s��${�"D����b�2��"9䚕��#D�`+��&2��-�� 8�dmwB>D�|�@ȗ%y�����&��yy�,=D����ڄt����R _�4�&с��=D�<*���-C��!�q�:)5�x�TN>D�t� �KM�8�w�P�0��H>D���G�~�4dc6cX�,�NTA�"D�L#�(�R,�}���zF�'!�D�	!t%�@gHw0P��Za�!��j���ST�6s`@SSd�$Y�!�|eR|�3��; nx�dn3y�!�dE��*� ��[*K�\#+�i!�D�9�
0���Ēw!�%J��ȱs�!��I��R1rщP�)u�퓤�%O�!�d�j�yІ� �G"����I]�!��K��b���
�)��Q��L�#z!�$s��� ݄iw�勤.�dh!�DM�Ih"�yL�ӭ�HP!��X9gDBt`��8 S0�t�Ը"Z!��]�d`�C�XHNqC����!򄌋WǊ�'Ϟw �B5/�g!��<� ���nD.}$<)"���U%!��֣fQ|�g-GH�2e� ȯ@!�$T H�V%�c��7�%��f!�R:^���Qr�U�:��hd���8�!��]]��;VC�.��1vM�w�!򤁖u�Y(eK�7� �Cw��<y�!�M'd��P[��0I�v-�s@ X�!�ˋV�͂&'�H���b`�S�"!��]�O�09�D�)~�x�n !�$�f�lH��'L��z��׸?!���"�\�+0IFBq�#�X�\!��8>x,�BE��#aƤ��S�[�!��S�<����g,Q�W
J�h�l�!�D�l�N�(�K�G_dâF�@|!�D�}ר0 u��77ED�ɂd�9Q!�d�8��w�Ѥ"L�����:�!�ċ�J]�qm��;9ꐲ��ϣ!;!�$�)l��\�bd�#<Ǆё �֬/!�d��d4 �$X�Q@$B^�;(!��GO��|�ÀS������ٕ5!�d^75�������?2��� N	f�!���(��'k�-��̺�]�$~!���.8��@� 8p�1&��'�!�� �`ل�T>n�V!��Z�a׸��"O�!xD"�"��Y�$��c�p"Ob}��hW��6=Q�Dg��!�$"O`Y2���7@���� �l��(k"O,eS�ݶ��Л��q�@���"O��!3�6��1�ì�E��X�"O<A�P��IzYxF��ds� k�"OB�Jׅ�~D~��5j_��^qhV"OP}
����9����Q*]�N���YD"On(�3x-�HrP 
���4*P"O<%Q���->� 8K�&�EG�ȉ�"O��2��ĚLD�	j��W2## (
�"O|����^���� (�4��"O0yxO[�G��C�/�/��؀�"O�RA��1|2 !.?!�����"O��Q��>1'F���M�^��@{�"O�8� Jɹ%����a�*~�:<��"O��I����LQ0��G�j�x�e"O��������q��I�5_o��3"OZ]Q˖O��T+��L��1)�"Ol��c��'=Ժ%�30���"O4�)a�Z�<�T�I�HIk1"O�@�2Ȅ2K,Б�N�T�\�Q"O+�a��U%l���j����:�"OȤX�n�:���O�	1�]c�"O*q� ݕQ�9[�M�v9�6"OZY�d,˟lS��1��y^p�"O6�+!�m�Nep `V�D+x)�"O��`����Xȫā̮DtΨâ"O� �S�[�SnFD 7_/R@�%`�"O4pr$�'_#�H�dG�lL��c"O6ęa`_�Bd�'� ��yP"O&��.��6��ذKN�H��"O,M��̂$�9*#Svfhj"Oz<���Z���I��Ec����"O�x�3�aDۡ&�*o��"O�8r�� S8Y(�[.���G"O�0#�"�30���0g�/�5P�"O(�3�J`�r��3VxT�Ps"O�5	pΚ�N}d8jw�@�}m���"O<�q�G���TAPkׁUN�M9v"ORT�G� N�F�[&*�7~<�xÒ"O������M� ���:]@�"O�Qq%�Oq��xpG��u"O�
�#�:x�ԉBC�/vꐵ��"O�q S�?:��`�B�/�"�ʣ"O��+!��eɒ0�'�J�y�$��"ONL9#D���ջ�(_�d_xŢ�"OZ8�E�ڃ"W��c�٤��@"O�\HQ.�3�T��s���O�B�`3"ON���<Ef �t
N4<�P`�"O�h����$iYH��@g"O��6�.3��$O_�Xl��"O���$�PS�&�Jn���*"O�#4��	v���R�ǘ2��Au"O��ʣ%G%����'ض$�0���"O����l5F��"�	�R��6"O�B�JNr"�s B(8�D;e"O��Zw�H-A58�q�
g�Z���"Ox��5fI���D�Զ�@YR"O
����#�8s�*A�ZΆ͸�"O�܃��`�\݂ F�)���"O� %ΧE�pa�2��x���"Od��&E�Au|�p7&�)�N��"O� �<)�d�9J-�CB�1o*4! "O�B�-��Uq�)�#F6I{�0�"O�d�FgVMf|��o9�Q�"OHM�3A�\S�X�C ���`!"O0�b�" �:ug�Lz��]1"OԬ�C��'�(�* #��W� ��"OzA�Ajop�6��z���1"O�`RPY�g L@X����X�"O���eO�?z�*��n\xƕ�"Ofq �JԔ*߸�J��ٯ`Q�QP�"O80���Tj�*��F\��|+p"Oz�" G�]䆡s�,�[�DS�"O(�D�ڭ;�>TҀJ�,��ܢW"OT u@�]L��֣I#c��=Q@"O�x�5+� ���q��K?��
�"O@l����� �x�x`��"���"O�A8""��~ ,{WǇF,�q"O�P�d��6.",ᳯG�X�I�"O������0�f��������Q3�"O�)qsŜ�4��T�@=U��X�"OJ�7�Y)a�̒l�'
��p"O�A���C5j	
$�'70c"OjUhpÛ�$#�Ԃ�N� ����"O��S��܌Nb�l�O�t�-i�"O<�sL�W�$X�*V���"Op��cu��WJW0��<�'��IQNB�n	�L�c�%z��pz�'��1�L�o����BM���Q�'�<���!J!��R�m��,�HD��'=jݛ��Ns�@'�j��p��'��H���E�1{=�U.׋�d��ȓ���q�CӲ!��M��8�8��R�XР��*���pҪ%�����=�N d[�C�������L�r���0���1�R�M��d�chQ+o�B��D>�����ߡvi �Ug��g�C�	�t�6|ч9�d�ԣ:��C�I.6��$�w�@������[?]p�C�(_�d�3����nx���#�̡N�C��5$v\�)&拒`�4�KJ�<�C�ɖ.�\`T"��)A�X��G��&C�	�n�=҃�6��$�#�#fg�B�ɶB��8��H+[���EA�cbB�I:�����/E�V�A3LFB�ɔ!d6�ɷ��G�XB����ZB�ɹ~�n<�q�$[؎� ��X���C�ɲIf���	|yܘ4M�T|�C�	�
(H��!�C℀rb�Џ	D�C�I8����-��0�4�1a�^B�	�D+Z�8Dᛠ���q��%1lB�	�\S����oO_Ŷ$�W��1b�|B�=$���&K�Bh@��ƇPT�B�	�{VX0�K�
S�b�3�!���leĀ.��"?1c�Q}��'{�j	:=Ƹ!q���ek��:�OJ��!V���e�O����tC�)�D	��N*�F�1*���!0a��"Y�:(��k
/|~��Q B���'>F� ����d]?I 6��1�P�b荓6ǉ'b"=�~zV��]#���&�>w�̀����Uyb�)�'8t�i+CLA�y�N�Cǯ�/����v����Ȉ���е$;vŊPiБg��s퉹������
�hh�83
�V��j���<��'MX������ȗ�M��E�V�z;���VG-}��[�����|��T+����4eէa�)���_�{��M�g��P�Ry�`�<E���� 
��������V��h��� �I��'F��� �:�V�3) �H�a��y� 1񑉈 s?j�'��
��f>��Aɸ+�L����@0W@Y�U�1��D�^%uA��0|�g��1xܮ����9=$��Ɇ�d?�fe̶'���)�O����%c�Iaʏ�T�fH���<Z�P�!�ݔ6���B�}��	~�P���B�L+|�a��L\@4��)�'�u�i]>1�`+��� �v���(�hO�����m����&Æy��x[�%�K��O��=��)�W̚�AH��t�E3yVx�A��|b�)�6%,��1�6�~�1Rm
�S���OU���][�C�:����I�dk���N_t&�;D���k��O�?�d�W�c���EaZ�I�И��O���'����}�d-�Y?��օ^�����r�XH���>h�bY�'.ȡj�O��}�	�������ܖ�0Q1U��n�����d@�t��E{�H��6pŢF"?��=a�l���y�.5�l�t��5;<�՘�� 5�y�
f��:Vc�6��96
��y���^l��fΐ>��V�V��y��I����ψ:4��u�E�M�y�� z�Xt�S��=*����0�W?�ybK(�t��e�"�(����ը�yRɗH�l�xb��GY�D磞�y�dN�\��d�dLJD��hj�Ȇ�yRm ;��E)�/:~��!���y�W�<n�y����9o�Ar�/�y�`'"��TX��J�\
D�!mL'�ybʏu�J񋇍Z1Ac3�J5�y2��~�h$���Q�N��e#��]��y����sH�{���1tG�-�"a\;�yR��14�N�dgہt!��� ��y�L��&�@�A�dT�9��"P�C䉸>��Qhn��:���b�|�C䉒�B�У^,6uI�d5)-tC�Im�}c��,Z��{�1��B�ɛ$WV����=P��Dǁ1i�B�I<'�Ԙ�c+!6\$^�kl�C�,!�@p���$L)C�㞢>�dC�ɝZ�H���	��y3�IG	x�B�	�]�8L��ߏ}��uRF� F�B�I�#Sq��w9j�uiO�[{VB�ɫXY�09v%��[�<U+t�RiJB��=*8�x3#���4M���N#"OB�Ɏ�9���6K�r��$�,ml�C�- y�ؐe#��0ZD4�u���U*�C�	�qF8tzAeE,dA2h�c��7\�C�I�`�ؑ��p��e�#˅�6)B�	 w�"����r��֌Wס�dY�|À�	�ES�d��=9�-̉M !�d�z��4��7��}�Q,''�!�dԃc��@ ��	�hߞ�#7���!�Ĝ9�^�����$n�ޑ�df�H�!��ӌG��X�i��/�@�s�X�!򤛕$�fH�D�*H	�C0!�d	 ������,v��у�o!��4)<ʱy�a�i���F@�9!�A����3@G�G�&!Z�N�{�!�dA=_��Ȓ�T�}P��	�q�!���y���jb
�Jx�I�R���!�dQ#�h����-ozU�@%T��!�X.�^�����y?.��NMR�!�dJ��Ը7�I�n<+��r"H��'U�e�e� 8S\��F�ViP�'+�*rL�%��E�b˚�F��
�'9�����(13��q�Y�5��1��' � ҭ֓7  *�`�4���S��� ����?�"aˁ>Tġ!q"OP��􂍀=%P��3K8�"Ob\R�`׻V��j�O(<*d�W"O���@� + ��p)�'&��"Oڸ!���74 bu����3B�,)�"OpY��+,'V���P w��:�"O�<��	�p��e�㣐�L�浹�"O:E�`*\{^����S�Y(XH�"O�X��/�5\s��� ��<����"O.1�W�7DB�&�k�X��"Ofس�.�c["��׊ш�x`S$"O�-��76\z��ʢ)���	"O�ɺ��8�Bz֡ʘn��k�"O�� &HJ�E 
�R"B� ��Ы�"O��8��X"X��A�#~$|�Q"OJI)�JZ	 ݴ�c�϶%� ��"O�4�@�%X�8�Gg�,D�a�&"O��Y�FW8;☘� ���d%<�Y�"O`�B�(R���}
��M-s7���"O�4i��	�--2��.L�)O�Ě4"O�Y�ժJx��=C@�ɟlZ�ȫ�"O��yB���S�hU��k�/T<H�A�"O>�)r��R�̴�"�.�Zu�"OD�8�.�$���j��
(}��}�c"O`�p�N%�� $$[�u~�m��"Oj�����d�<+��	{K�5�`"O�X�����Rw,U!��"O� v��`��p�R,�9S"O�9�������zwJ�w���"O���e�˴g�ҝ��N�v�`\�"O�!��
z5�a�3�' ќ�b�"O t����9�2H��$ۄS�|a9$"O�aS�<S��we��`�"O4I!Ad�7MW^Q(s�?��՘�"O$%	�,؅>R����mG0c��a(f"OЁ���1�*��'�%vg����"O�Cv��38#�h��*�,f��T"O^�
��� �0@I܉1d���"O�)�G�oq���g�q.ht#"O�X��/��2bȥ�%M�ch|xR"OF,���@�UGz�eZ+@#�)��"OR��r�L�'��s!D�.�a�"Op	�cZ�o2�
%s�l�""O`]yd�^��%*@KҾ���j.�yR�Q���yCɐHH��̰�y�a	9| ��y�@γ2  �q�ϝ9�y��
�*/x]ؑFK-�����A;�y�@�
C���)u惬x�r\��2�yҫ��1�hrc��v�,�X>�y"KӠ��A�VA˥~�"�u�[+�y�jі%� �AT-,��8#��y�Iѵn=�d0�jƿ%C<���D��y���!=�b`�FM�P�,�1i��y���#~%~�{��,aU$��L���y�!Z)uN
�i��ȶ"UL��Ad�!�y�És-��[����Q�:��!׾�y2��e2X�C��ηC(�#q�Ϋ�y��ϒF��26�џGR�i���O3�yBE�(?D��r�F�D�"�M�-�y�FG'RC(��7�vg.|�����y��Ѿ9���2(�(hxp|��g>�y2Z�bp@XcP�(c�8k����y�͔��8��$�K�^ڪi桀��y���g~�z���F4����O��y
� ��S͓�Y�j9BV��5��t�g"Ol��4�T�7L �I��՜z�����"O�xĂ�v;Ľ�2����a$"OP	۶��9yX��B��ɶ"O&�;���>R,��`C�
n�y�"O�I1�҈�.aHR�S\h���"O��O	 *ԑ0gT,J��ò"OLh;�Q�Q�C��2'�Z$��"OH�.ݓXy¥h�"ϰ
����"O�X�s�.0��[D��3?Pu""O|���.��͓�Y��rP"OVH1�Iγ(��'gŸy1���"O�X�Q��jc>�t�ѥ90Z�yQ"O�x���2ZT��qE�/Y<BŚ"O�,2��5� .�5J;��b�"O�M2�,�jZ�@��؈g"O�9h�)I@`$�#�z!!#"O>�
�L�5@�Z����f�F��"O��Xmė\�*%�g�"��}RC"O��K� ��H ԯF5F�T�a"O2�P�� 1.9��T�a�@&�y�������o�!C��U�D��y�"W�y����oP<m-�xŦ׷�y�
Q8'�8�v wND�"6�H��y�m��I��Cd��s��pi���)�y�+� �Z8�F��*9�^���]��yh�5Q��"���.�4i�E���y�
Å1�jm�� �!rjm+ADR<�y�L�.ѨU�c�	1)�dS`�I��yҡҟ1����F��-W�Y���A�y��խ`�P��W�Q�%984#�I���y�"��s�i��l�Ӟ�Qa�ɱ�y��˦#\�Y8�+΃�Z=�WL��y�
�&���z&�E���$!T��+�ybW�{q��
r$�r��s���y�O�x����˫b^\ �m� �y�ϒ$���Yt�Z��@�ۥ�yr@F4�^DS7l�6��,3�,�y �̐H�����邉�	�y�U�&Q¸����#pq���a��y�V#tQ,(�� �n|L3�̋��y��A��$I0G��@��+\ �y�Ցyײ�ڐ�X
��*���y2㔃����0쒒z�4���X��y2���i�j}	Ѝ�#\irوA����y�ϔl�<y�/RS�v���y�������J�K�	D��F ���yf���I��J_�>�xC�=�y�iV]�]��B>Hd=�ȉ�y��x\�R�=����+�*�y�dO�}���`OU�5��$�P����y�FU.����al޼�tS  �yr��#�l\��Ɵ�>&Ձ�$��yB�a�<�`��w� ���yB"ƱT��U���L!���:eM��y��B	f n<���T{����,�>�ybb?@ �`?��\�ЫH(�y"Jڛp_�U��aY� �^�����y�F]�L�Bً�Îp�� Q��ؕ�y�f�1	�t@��0iyָ�%�ϒ�y�/��������?`Nf�Gg
��y��U���y�)��U0�q�g��y���sb����&�-K�`�u��yb�Ί6�`D�Qg�7 ��,���y
� B�8S+�6�� #p��)4ch�&"OzEb�YpU�t9"h�q��|[�"O¤�fT�6��Y��ئp"O6��I뒍��$&m�J"Obx�"ؖ]��BT�V)0�2"O�8R�&�|`h�"F�M0��x�"Op�z�ǣ
���W����3"O���~���;�MB�C��	�"O�13P��a�8X����@��"Ot%I��3� ٳoM�j��QT"O>t(�.C2]R�i*"oJ�r�V�*0"O򥡄���b� R�`傅q�"O"me��!��P�p�<<��[�"OL��Bޥ_c��갩�
��U�Q"Oĉ�b�ԶUJ4�0��.��a"Oh�����N�L(���_�v��Y#�"Or�4��4.��5��� ({�8}�"O�	���gުXP�(P�6�R� 2"Oʡn	   �      Ĵ���	��Z�w��W���C���NNT�D��e�2Tx��ƕ	#��4"�V���d�9�AmZ�Z||�jUj��CiڐU�X�_���u���s��0��� �M3+@�>�����W�r��AY�x�q�'�ƙ�y���a0��d&�D��I�e~���g�Py�)��O���k�b>}B�K����ż��lRE���8�\	���*[���'=�e��*\*?� q*Oz=w�X�WF&z�	�-��E2@ �$�锇�*dB���׶�><%��"7Ŏ?fo|$>�@�
�y_hy;�g
�i�5���dZ*$@&�|���7s�*L�L>)R��Gf( �@:��9cL�%�}�`�%jPp���'*�U��B��'�����1�~��b�$���*�`D\(]u�!
Wh�9!ǰ��A�O��Γ>����p��<�'.S�l"Ѝ�)N�4��,��y���>$b�̓b���W�{Dʹ���ĢE�U�����'�>��C<k`ɻ!�K*z��q�u,d��F�����󟰺P�Ou�l�O�h	��H���#$��s�
D8iH>9��(6q%��)5W�f7���c��Ǖ7�<k�Ō
yi�I��P��%(���?�|TP֐>�P�� A���&���N��ls"DL#Re�$J�zy2��O��Q����5��'2����M���#��^�n�dP�w�]�X�$��H���0X<�	��y�힖�����p�3qΞ�.謳VE�$�z��'<AP�a����Q��Z�`�u�	�B��Of���"؄{�Pl�$(	!���Jq�|҅�G�����y"h�%D��m3�lԔ,E6Y9)զ!Dj��!��6a�R}�b �@Mz�OH��W�'l$'� �KP���f.U��(�#������Z8$�6�|d�q�h�L<!��PiJ<a�w�ͽ\�BA,�rۚ� %$DM�ɭX�&� 7��r�O����SA<T|`|�w�A7�^���'���@ ��  @�? ��#H�D�^��'�L
@ ���  �;��
"�R�ȓ/���Qj�.5����n�F,}�ȓD����0�\A�`�q�t���������SS�=K$�P>_�1�ȓt�Zr�K@�@�r�� �܇ȓt�L���gV�Ypd���ڔdt���~�̭B P�f���+U��؇ȓz^�)hx�9!�Rm6���2B�P���.�l�E�ʑ�Ь��vG��� �/��     �  J  �  �+  �7  �C  �O  �[  d  �n  �y  �  l�  Č  �  J�  ��  ��  I�  ��  Ը  ,�  ��  4�  ��  ��  �  O�  ��  ��  D�   e � � 0 �" ) `/ s2  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����ȟ$� ��@��X@Ƥ�S�Ys5"D��8a��+B-����
 Bc���*��Q���'=f���4�HTk.h+��4a���ȓ_�R�� ŊU�`us�1\(�Al�
�HO?7M\�������<�����\�/n!�Z�v��r�DL�4�:�7���'k�Ik~�)�4��"o�!���P�e��y�/�'��T��[�dV��
ƪ4�yb�	�t~��`�,H1`(�c�7��=�y"��b�hݻS��%�p�A!����M�']�i�T7jj� cV�a����'�\�k��]�q����U A�����	�'4JR�I�7<!�7���&<��'�2�+d��(my0�F�Ph�Z�'l�M@��A	y&�÷ƜI��9Q
�'��@c���W�� C�:l�	�'V�)��M�7̠�SQd4���@�'���$kJ*d^P�@���,d����'� �R��B&7���p��8,�x@�'�Ԡ��G����y��ӱ+��Ћ�'�<\���Կ1�=�`�)�~-���� \��f��bm��r��eL�t���On���!d�>�'f��[_0��߷E���?O0�7��Oڨܺ��-v���:�"O�DrP��,S԰i�&IǳI] ���a�O�4�	T��h���Ӥ6,��<��'N�#��ijd2#낪t�
x �O��=E�D��`�؂�jӇ)����V*:�y��$/cVE�t�$
=�&@��y���ĸEh�"Q�Z�{'��Px�i)�	�A�D��♙F��$&w�P�'���쏊��m*D�4 W�X0��HO�P0!Z�A>0}js��V�H�[��IA�O)Bҥ5��( �,8�,X�J<)�'rz�b?ic��Ĺ(����g�.��Cӌ4<O^"<�hޡ���r0�S�MR�ăId�<��M,6l@@f(p~�����O�ȗ'���������$���� HјM;�P 3bCUW��ȓ~x|A�6�3$��qu�N�b�%����I�)`ڬ
5>Z��aHt�C�_���d.?��vӎ]�a �E#�m��H�2=`�"O�<����2J��j�o�� ���b�O��Dx��L�`�1����:v����'%0鑠˽{.fM��!@E~���'ў��D�*9�T��6j�x1d��B�u�O�<i��I�w���U?ETvE9��DH�<y����EZ���֦A���rgF�<��,�48,��"��"̎�Z�=Yɦ�[���9O>Ip��D5x�Q���T9���+d"O��B���Ē���FVWDhcs"O2��㜔+e�-����OO�5����)�S��F�v(\ �1��1	��0���I�-�!�$ݪT��D+c��-�L�ҧE�.0!�,t+�KG �(;�l�Ѓ�H�!�$��2	"̊��ø��K���3n�!������h�%�-��\#��95!��2��P���
�n̐�q�!N6)�!�D�8W�\�4��-
�)��O�v�!�+���Z$#��K-��8���|!���\F�rViȯF����`O�������)��`���^>���G��(q�كB�:�O*ʓl��5)ը�|�h�FaM�{�۟'.���'�(���8b�Q���t��8#�X#Af|C��E 6�JAF|��ӓp��-� �$G<H��+�,`_��O�I�ۓL�0��a�˲�a�B�-�?��y��u>�����1
�
�tq�t�T�Ϥ2C�y��'J!��< �A���Z�H��kb��<_ў���)_\����"xR��A5űOP��o�t]�B�=���2w�3r�, 0���Ej��'if�@s�Dt�'<�T{cϊ~B~�k4�ŁXq���K�#��y5M�jD�x�׭@G���<i˓+C��0J�3���1f'����'đ��Ex≅3 Y��E��K�� ��Ԓ�y�ꁬb@*�,GNh�e��/�y��ڽE�j�V�rK�0zJ��y��+2ݞUs1*�5kn�LbwL͔�y" �s����5�בj��Y���"�y�@P#@9��ʔ�)enx�B�aP�y2f,'��$S��Vh(����y���~�����	P�T��y�ǔ��0?�.O��*I�~*jـiI�]#�c�'A��$c�(� F���{i�*HB�I$E]vM������Dbe�>�dB�	/(U2�rF�_:3İ|[+�91�C�	�7�th�N�#.�8��V�D��B�)� .e����+l. ��
��|h��"O���n�_rX�ړ�F�:{�q�V"O�H���]����B(
���cD"O��p���]�!�[�:_9:s"O�5#0����)���_-Hp،P4"O�%h�W�_5j��'�Z�f>�x��"O%�� �&]+D��Y�.��"�"O.Q�)
�8^�B��q��#"OD��.ٚ4�(!(b���3�R�JP�'���&P�8��` 4"�=��iY��6��D*�d��*�#"�Z�J哃�ӻ!��0Մu�q��ϸy�d�F�'�!�Y�X\	�ĵR��Ȉ7m!�$H.
��1P�T }��f�	�2�!�$���݊c�6uռM��)��,�'���':�̚6�_>���6n�A��	S�'ݛ��N+#WM��>ahz	3�'ɖ�yrnU�'���RB��e�8D��y�Ņ�"~�<���N�d�,���ý�y"L��'c8!�a�,h'� ����y���	`ƕH3�7K"")1#C��y��c�:y�RŅ#E�6����X�y"��XP��`#e�!O-x i"j����?��'$<� ��N�a.��Cd�U��䌳�'on�pqk�	^&I�ӧ���J<��'1��)��Z�=`(;È�Io4�1�'2*���7�LD���#YxFD��'<��3N[�Y���!(���8�'�����*Β=V�ِ���x���	�'cĬ�pˈ�L�]c"��3��a	�'�ƙ1�ڤwq�������K���'�j)Ӷɩu�l���^��4I��'-��{�b�6HR�q$�
��q�'ψ4#��_�f���s(y}LT:
�'2h��  <d9|@&��>��]9
�'Ҿ���n^;:z��fV=�bH2
�'u��I���Pj8�9դ��2��-�	�'Qh82V17���!��6(��Y��'�*Ʉ�Z�C{z`�+կ�H�C�'Ќ��� ��
�
&�:>�
�'0��Ċ,1P����P�A3���	�'ú4�T�3Z:�A2�?+*
�'�$�ۧKC�LNr�@�U�
�LT�	�'���+$@ť4\h\Kd�	:~@|��	�'�dy�QC�`rP�t�sa��0�']���CP
YA�������a�.��
�'�b�BD#J9�zc��;bM���'�`�w�;^�v�kჹZ$���'�N9c'�ҼYK� '�ϐQf����'	�r��P�P`J�"̂TX�
�'P<�`"�v�>�
5%Y!H6<<�'{�<�r���Y_�t�#�-�f�
�'�A ��z�E��������s	�'H"�;��5Z��Hٵ$�D ��'�^}���$`��ૄ�I^�D3�'�ĥ�G
��MÆ�*e���,��'��]"�LG d�lc���M�δ`�'�\���(ȦV$Ht
Z7>|6 ��'mF�xS+�A;^�s�C�#	��I�'
��`A	=�`��]_�!�'������h�&�0���&��B
�'՚iq�j�����D��qκ��'Y젲��Ç&L�
1�P7nE����'nڐ
"�K��%���k�^l���� H��P��)���:5���I!8"O$ �g[�bw:�x2���)����"O�hQ�Şv>P�̜&�L�["O8@�ݯ*�8 A��XT����"Or @\�X��XeO�_�TI���'cU�������֟�����/R5@Fd�se��sV�ژS)����ğ��Iݟ(��ϟ��I֟�������ɥ7M����FW0C�<� �D�W���I����ǟ@���P����H�����ɧ)QX�JuA���"E�ӡV�3k�)������ �Iӟ��	ܟ�I����<f1�Zg�	�:�����Y{wp���럸��������I�8�Iٟ��	�n�n�`�G6:V@���38E�	�� ���4�I럌�������ɟ����!���`0��Շ$�z��I����Iß\��柬��ɟ���ڟ(��1���j�.Y�Yz���dNfA���P�Iן�����`��� �	�`��.�Kr�P=P�V��E��$�5�I������D��˟,�	�@���`�I>X�d�O_�l1X%Z��	36���ß��	Ο���ğ(�I����Iȟ �� ��ar  ��z���C����I����	ݟ������I퟈���X�I����h!��?�51��ȟ/�����`��ɟ��	ɟH�	ğ��I���I�S�8�x��Q8	h��#K�o�X���џp���������ןX�ٴ�?���B�6Źԭ�0%��պ1�߯;[���]�(��ly���O$�nZ��TӖ%](_��hKfk����%�!h*?��i�O�9O�l�0C{�$G8��w��=��+�����Mc��I��'o~bdع	���R�h���� �xܐ�'�̪�2�nϚ 1O��D�<��)<F��s�\#f� ���7�*0o�{��c�`��u��yg��%o�BT�5K�T�N�"&��gv�7-Ȧ�Γ����M:��aU8O���B��J�� 8���	\� �z�2ON��*��f1�HW- ��|z��+����dˊ�ށ��bZ�I<�=���$*���ܦu��F$�	0�8�D�	@���g \�H2 �?y�]�8�۴s���:O��7x�咳�����#�:A�\��'T��1��Yz&�����꒭e|*����'20) �AE���1 I�b(�a�6S�p�')��9O�|��� xy �CM	���33OJ�nZ.~�8֛F�4�V�Xpm�
E+Rq��[=��eYP1OƬlZ��M[���6)�BcAg~�"n��h�j��k`ͻ2���PЉrt��>�a��i>I�'6�O78��$d��P �k%�!4$��O8�n�<kb�D��p�S�[�Z���i]�g$���A�$z�l��OJ8o���M3�'��O<���'�� ���AԲ<s�l��E0~��}�UI�O,��c��t�|�p�@��ē��ӴM�j���3�u���ճZr2��<�/O0�O|�oZ�g6��	$ �`&�n5Ҥ�v�ǑLi�扷�M�����|�ߛvs�
��ޡF��E9W*��a2�c�B�kt�P֬ؔs��$սe-�aE�ѣC��]��O��b5�
��8a�2t��+���s��t���	�T�'&�)�'L ��a7��! �hAɕ��2���<�W�iT�!��O|nZ}�/9�(d�jטk��H��zr����D�ئ};ش�?i6(G�0Հ	�x��$��Vt��37��WfV�aOʡ.#�4��� pE(AsM<y�O�i�<��(�}"�B�Y "Kə;��Γ��=��]�Θ'v�>W�̵[�E*r<�aRÎ;lx�W��	��M��i���5�����pv��BhB�Bjݠ0l�|���7���Ӄ��	��I�?�pB��^Bܩ'��'^�*)p2��sLʘ�������IJyR���O��	9�Mk%�x�D�yC�>z�	K�ˑ rӪ��'��7��OʓO�i�'�47�S��P�G�J�����B�alZ��MKC�v�:�ϓ�?�Bf�{'��/��ĉ�|Yp@���	J���#
��^�$�<Y���?i��?���?�(���y��_	����W���\�dMQQ�֦yi�~�����,%?�	-�MϻN�p��,� �ে��	���ּip7mBğ�է���O�4.>�A�'�ԁ���X�`�᷉J-j��' haE�B��T�2�|2�|b�'�.���m��F�����K�!�THF�'�r�'�@��S��۴s�h��'�?a�tlʡ�� W�t����^��:H>��`"�I>�Ms��iV��d�>q�ǌ�r/zHY�G�I�J|9A��<i�<�yb��D��6y",O��鞼ZaB�����O���	W$( dÓ�ЂMWαR1��O��$�O����OB�}���9�4�22kyd��F.]�����ߛ�	χ����)�?�;2�X����L��|�@g�ω/���/����~��UlڍR^v����,?iV���W�X�Í_�7��(u'2]T��8�%I	t��H>).O.��OB���O���O|�BL��X���V �l|�Ԣ�<�ѹi�0HAP�(�	^�'!��y(uNޅo2J0��O�	�dU RY�|�ڴkK���O(�l�	��K��ۏ#�f��pD3�P9W"ݚw
P��+�<�D�	��q���/�䓉�d��V�h�1��)U�ȩ!F�d����Ox���O&�4�.˓E��6��'�yHRT*ޥb�ɭhX�8��ǂ�y�t��$+���{}��bӰ�m��M�Z�6J܀A���(r ���T�Cs�I!�č�<i�u(��x JW�5L|��,O��ɟ�� ��bX�Q�����L�Z��-{�6O��$�O��d�O��D�O�c>��d��	08�(K2��
p��I�wJ<4��O������HP�f���	�M�M>�eCPd(صk��-��%`�џQ5��L�>�@�i%r6��F����X���O�� 	9O�tY`�EW�2����G�M�V�p����N[��=���$�O֨�'b�����h
f���6O��OB�n�uz@b���O��L�ް$/ش����6V� �OR��'6��ڦ�ϓ�ħ��TO��F_@<cb*܆:�~t
��/P�$���j�� �`E�'���,TeGH��B�|��H�#D���$].&K��Ud��I��ҟ(�����d�ަ�i��Iи�Ck��qVH�$��'��6��Ol�O�9O�al�%E�x 2$�5w�P�@(�]�
�iش�?1�gQ�0���?	Ad��W�A[c�ZX~b&)'r�C$J� Q����gǜ��'��W�`D��`�qY\̙"�
�NQ�@�S/(G~6-�xQ1O�	+�i��.i���Q��&ɐF��R~X��4Q>�v5O���|z�'�?��Δo���6�#�(�,}4mM���i�g�B��r�"�r�1��4�F��$W.e	�>0��	�cY�SW�Ĳ<�O>�V�i���ӏyrY13�n���EťF�$±��{&��|҃�>Ab�i�V6�|�x�'`.�`M��h;�0�$S�bj�b�'�2�ХDo�x�%��4��$�,0���A���dpI��K҈�42�\����Ȉ[lx���O����O �7�S�?�l����#�Kʧ8%���1R� �6���X��Tkڴs<�I��?!d�i�ɧ��w0E�Gx��à�J�"m��'>V6-Ȧyq�4aE�3�(B�<�49)\xI� Z,g6�W�(��Eh� W1��l�J��M��'��	���֟�������I2p���!���W�V�@�͚K�u�'�&7MÅ|n�Xn������?���\�I�P2¬�s��-w|H���B�yC�a�O�n��M[�iF\���������F|�&�Z�*U:$�sfȿ,$V�@en�>�����z����>s�'��I#�h@��/I�P�0*6��_�D��ٟ��	�<�i>��'��7��/0Lf�DR��~�J��y�f��U�F�9��I�MK�rc�>!u�im.6Ʀ	��
$V�-��.����ai�p�J9W������Ā��^XR�EPXy��O���'_F�"��1I����G�?��	�<�	����	П,�	]�'u���qǽgI�e{PD_�a�L�A���?9�"y��R4��I2�MJ>Iu���.� a��!56#d�˧)��UF�\��:ڴ���OPl9��mC���ґ�I�K5@ ��S�;����X�E�Qc)���<Q���?���?��� G�}�."��0����?a�����aP��럤�	ӟ��O�l0��H�0�$MSP�_-4S���Oxm�'�6��Ԧ�	��ħ���OO%A��iHQ������)�d)��B�7�L��/O<����DL\`�O�E�1�S0b�B|0'���%�(�a�O���Oz���O1�NʓY-��B!`�̐�@�t픩c5d&W�#�Y���4��'��e��o�7e���a'K;DT{�G�K�7m]�i�t"EՊ��ϟJ&k�"�h �By�BO�]�tE��&��1����&!���y"_��Iϟ��I�������O|+dI	�pc@h�R��/kO����E`�l-�V.�O����O*���$I���1B�,�H���hZ�FY�I� �4r͛�#�O��S�'�$�zI��<q��:G�ܠ����3D�ɚw�U�<Ir�V���#��,����$�O��D�%L4���ۆB��J1S9=9�D�O��O��;q��J�=^:��'��[4K�� ��<Lt t�F%��OL��'9
6�U���	�������sO�I��<	�� 5oāXn�ɠy�@��qJ�H�'?u�RC���H���#�m�'�
�>�$9�#��3�R���џ��	՟���b�O��A.b�Yw/��fͰh�c&^68R"{���;���(�4���y��2L+�L��D�_J>�SԋV��y�&gӴ�m��M�%MǄ|ǐI�'o8Ⱥքެn�a��e��5>岱GS�Mr�h����&�'s��ɟ���ٟd�Iɟ4���3:x9���i2U�K�O��ؔ'B�7��	����O��$!�9O��Q���TP��wf̋X�굪`�M}�v�F�m;�?���i�7N�t4�b ֿ��mYq�%)��)��U�L��]hб4�]�T�0�M>�,O$���6��\�$߇g<]��%�O��$�O��d�O�<�4�i;,D��'N�h�#I���AX�Z�*�N��B�'�6-3�4�l$�'�27M�ۦ]Q�4_���86	�9Z���/ʆS�����È)���Γ�?$ '�"0	V	�9�����|��1-(
���"An�L����.X���?,O��S�Od�`c�� z�u�a��: ؘ �y�`g��1Y����4�?A/O��s��L�}�V\s�CK�T}�2"j���'�p6͏禭��b�`Ũ�nn�����q�.�j6J�7�h4��fQ�P��}����c���H�S����R�t�I62k�ٲc�¹Dֹas-����m�	��MKG�p̓���'�0l;�')(Dɢ�G�*0p�$�'V��Pq�ƬӤ�R��?��o�&�:��3�.�S	\�qx@@�Ӌ�qQ>�Bq�Q� |�J>y!"��U��G�P6:�����O@�S�g~2�e�ZؙP�1Ǯ�+��~^�RF��H7�I��M������|Γnw���(Eٞ�a��[$Af�P�)�Z�27m�O&��f�K� �d�O�=�6���MR�Ԁ���� �ayg�NLܵȢ��3 ����Oʓ�h�"��!�7g�<!{�U�F�0��G��5��$6�	D�'O雞wӂ�"Ʌ"Em�U*�!��	�\ �1hӤ�l�<Y�O�i�����mK�� �7OT�R�K/G�����\T(0=O�$񇄔{��B'`%�Ĵ<ͧ�?ylٝ��[B�T�W��;U��/�?���?�����OȦ!w-�ly��'��@֦�|'V$�#��&{l��	�'l�'j\�V��v�iӀ���k}Rn�߄�R��nB�wMި�y��'� !�b�R�L����X����#~C�%�7*����0!@�Vԑ�^�_9����	�ş��	ןx�I�D��w����ʩ_P�5P��٧�#��'��6-L>?�˓s9���'`ɧy'�.W�0h��o*�&��w�
%�yҀo�(|l�>�M�����'p�ϓ�?�'��v?("1��+z�L	@rKڣe�.M#�*�>2���L>1(O<�d�O���O~���Or���[7R�����k^=P=��x�.�<!%�i[�M�Q�'z�'��$_>��zg��Ĝ�IC��X�
ښ挴�O�o��MK��'��O��O���Y�l��{������BYw� ����*�N��E\�,q�C6Z�!��k�	Yy�H���at��=���者\���'7r�'�7=��˓uӛ��7�y�˚"n�Q^$څ��@'�"X��n֛F�|�Os��HD��`t�@Uo��X�>t���g���H�0WdɺD���n������vf6<P˓��7��b�c��<��eY��Ȟ"�R*s6Oz���O
���O��d�O&�?F��<`�� Td���!li����ϟ��ٴ[4�$��?aӸi4�'�pP�+�|�uo��.����"��O<�[��VbӬ���u|R��&?O���N_��g	$& �}K�,�9X��!��KN�X�  6�D�<���?a���?����l`�p��-\��f� ɍ��?������}�v����P�I̟���?��*@`�9�"��P ��<?A4Q� �ݴAڛ�*�O$����[vob<"��=�d,vA�Ij�u!��u����e�<1��<�p�gO����hN�B*�@:��1ţ�/�px����?	��?��Ş��̦ѱ��_%��-��П�5�)��]��a·U���޴�?!M>�sY���ݴ͉��,n<t�Wc��*n�T�'�iZ6��-s׾��:O���A�'��`T��o�~ʓ>�B9��_�5�Z���m�7|b�͓���O���O����Ot���|r��!<p���O�A�F\��#qF��-DL�r�'�����'�d7=�H��㞪]E\�C%��j3�}����p�4V��W���?q��0���ie����`^n��H�([�f����k���fA*DB��ef�	jy��'�b�V?������-��t�pʞ��2�'LR�'���+�M��*��<	��?�v��*fLe��.J�t�Ҙ��	��?�*O���e}R�eӾ�n��?��O�i㗃;�`,�4��f�<�D6OL�Dɢo���#�Wd.�����k�:\0�x�G���U��*�j��[�;�z8���?Y��?���h��Ć ��`���t��qH���t�d�Φ�B�8?��i5�O�{�����
/�(UCs��|���ަ�۴^֛�cK;L��؃�'��
u M�'N�)mCh�!a��9G�l�`$ФU�,@��|2W���I����	۟�	ɟ�ۀ�;LJ�"%��(EF�rA,Oly�s�f-�:Oj���O^�I�|��~ � ��+`*q `X!
��Q�P��I�4'I�� r�V,$>]��?mCl�8�L��䁇�w�b�����'
�@��C��ry���o�(�b-6��'n剋^$ %����j9��ad�[E�������ӟ��i>��'`7m�"_@�W-#И�Q�]�M�:]�,�'�D�ۦ��?!cR�t�޴d*�F�埸�R��i��Q�MU���T�W�zQ˜'�2EJ��8A�u(�io���?��^c�ڌ��8K����-��X�(x��'Q��'�b�'��' �0�[�F�;v9�H�!����J��'iR�j�h	�<9��iC�P��C�KK���-R-��
�9� T��?1�OTEm���MC��:H��
���<q��gh�pa��Q>bx���r�y+�Ik�`*����������O(���O����F�p铁�ύ5�)Z�n$��'�S��XشS�����?I��r�'S�R4�k�_B<�����0I��'��x-�f�~Ӣ���B���?!�7�/j��8s��Uh̓����xۄA*���8u%��'&���Y'��b��|b�ȷ
'�-���.gVUq��� ���'�"�'%���P���۴r+�9H����-
�q+��X)Q�2���b����d]����IM�I;����Ӧ�3�'+��%�ŰU�x��F�\�M�4�iH�+�.5�y��'�́֫*�Z��!P��+h��<��=�AAB�p��p��-w���'���'���'B��'��yV��١�S6G�	:c��� f�p޴;�pΓ�?�����'�?I��y��
X:P�3SE�e������A|7��6�I�hէ���O�TF B�j�'$Τ�w/X���BF�^�T� [�'˂�h'�V4X���8В|2R�������:��	�8k���m��^���'Ib�'剔�MKg�N�<q���?	��}�~!c�@B�&d�o�䓞?��_���4E�F��O��{�^ s�L������d?a#>(͓�?C��]���Rw�	����럒��]� ��d@�%�ȉ��ۑf]�3$(`\���O���O���)�'�?����Pe��?lТ�XW&A��?��i`��ѧ]�t3�4���y��@��$d�V��ek2Tq,�yB�n�&�o�
�M��̀p��͓�?���ß~��A��N�? �a5+�^a0A��,�<3*��p@&�d�<���?I��?!��?&ˊ�l^��SR�/!�V�B@�����@[�͔H�I��4��P��'���2�!�:�@Ģ>@��tL�>���i�7�ޟL$>����?���
W�B���Ӣv�"U�@Ĳ.��yP�f�fy�F�?3n�I��ղ5��'1�	)	�d$�hǚ�
�B%�5D5�I��������i>��'ʨ6m�?�L�D"3�6��1��:+˚���͏	au�Ϧ1�?�TW�4@�4_B��'q��t���ڹjRnJ�xvzy��EV��jT! 9O2���}���N@�P���rԶƮ�s(BI��/�bӫη�y��'��	oy��	�9���"�#������ϩ#41ON�mZ�S�l�j�f�|�`�9j�A5iKf�z`�0"	;��>���i��6-�O��3 .T�&��d�OF,0�`�(�F��,h��wo�:I�f��G�j6�=ͧ��D�O��c�Θ[��X���r�����=O��OInړ|O�c�8���?��盾x����So�V�X���9?�US�X��4W��>On�,����4�\����X���քZ)A-�8I�Ͽ%g�� 瞟���zA><��]T�	��h�sUe�/mc����#�~�(��'�bS�b>�;�6#\G�����-Yþ��@�&,��2�O�YnZu��|Γa���mIi���v�Z$H(}jPeW:�6��O��J3���OG�D�O�����0�Hr֐��Psd�XE�e萯H�v�M�ro9�	H�'_�>u��L�1�!�2䆙 05Q��Q4�M�'��}��2N~Z2��y� :w_V8�� ��J��C�fZ�r��6�ʦq���4�:�	�O`\Y��K�Z�󤂶L�7X���녨�hi�4A�3O`(��Ծ[�f��f,�D�<�'�?i4(ش6U88g��t�P)''���?����?������Gڦ��5�����I�d��(ٱwG����MM�!��D��kן'�\�O,n��M[$�'��I�~I$|;u
�?�$�rħ=�����(�q�F�6wp�����Dyb�O���.6x�܌Y�2�З��3*̸ӱ̌�!��'C��'���ǟ��;93�%��Ȋ0kH�T�\Ο�rڴ`�FP͓�?�C�i�ɧ��w�ک�a�<`Ű!�3z$�`�'X�7�C�M�ܴҒH;�N��<��s�EQ$�-b�t��b3���M�3��������䓲�D�O$���O����O��D����0��Np"�kc�E��tX��H�4*�<b���?����.��) ��-6CϧL��J�%I!����'��7����-!��ħ����T�r��6/'p�颷�	?�Q���D'Q�(Y!)OD���d@�Z�Hŋa�)�D�<�"���~���!U$Eq�n�6�?I��?���?�'���Ϧ�q�{����͔���� 5�I>f�p0�~��#�4��'�Z�\��v�u�VtmZ@@�d�0q^l�`jƅA�бS3� -L���	�����V `w�X�d�ny��Osט�0�p �O����#�?l�I����	̟x�IƟ���R�'M8��C'��R���`#,���?i�d6�FA��'��ɨ�MsN>���P�0�hP�a�6<D��!���\��ڴcu���Oˢ����5�y��'Z9�ro�5Ij��l�_�XpY���b���dF�]��'��ꟼ�	�,�I�/�A���^M��c_�� �	Ο�'56푗[��$�O>��|‣�n$L�[�Jр}3&��<���\�����M��i�6�b���?9��c[�L7F���Y�Jn��ZQ�W�f�C/O��I۵^P��2����2��E#%�ͪCd�	 �O0(l����OJ���Op��<I�i��sR�n�"�i�n�R�>	�#��y�'�
7�;�4���'�.7�0a��H�.V!xh ��[(iuN(n�?�M��B� H]��~���
}Ʋ��@��iy�*ޮ�\��aʖ	�l�"%aE.�y�\� �	֟����\���P�Ot��H��"7���P *E:@�|
�#|��:�6OJ�D�O䒟X��ڦ�]�G��dT��E��b	*%���۴\՛ gӠQէ��O%����7���[�'u�=�QFɊ �hq�I\*z�� �'Y�����r���2�|�P��I̟�5����)�阔<�.4�g�L����˟X��@yB�`�c7��O
���O�p#����iB��%.Z�
���ON�OV�ק�7͆�������$�P3}���^��bc ��i�d�Op!�CL�0~ ��4b�<!��xq��D"��?!�@N>.���p&Š3��U�6���?����?y��?a��9�]*�MK�%-:!��)�nI��"�O(���0��Oyo�E�Ӽ�cb� v�T1huE0w��`@�i��<a��i�7M����+���I��,;T��m���1J �%$Pǃ�#[����;T$��'��'���'^��'oB]K�Y�蘹��̀:��'R��BڴXl��͓�?A�����<1�� ˬ�Vbߋ�D�[�"Pe��2�^���<�Ma����O���)�?K��Hۀ�s�D��g�~,��S-�(��	�18��$���7Ңd&���'��aatD	�T�Lc-�-�Z���'E��'������P�\�ݴ� �ΓSsb�a����>�-�Ύ�z�<��C����V}�-u�j�n�/�MdB[�_"��A���eZ���ٌg����%�<��dA��cV�Y��R*O��)�C![�r�@��%�"DǺ�c��<!��?!���?!���?i��4 O�#5$��ǆ��2�ح�G�	�=�'dRz�<��g�<Qӽi��'0p�@� ��(so��jժ!�� �O
�?�V!v���6`)�,����@%)� 6|ô"]�k�ܸ�H,��x*�	\-S�m�C-�$�<I��?����?�c��/��	PU<ym����"�?����Zߦ�3�'m�,����H�O 0�( Cǃ_L�9�C�N¦��O���'�47H������ħ��	ÆX悥k�Ϗ! �Q�W����QmM'DtX��)O(�i�� ���SG(�$�������wI�h��d�I�@��ş �)�SVy��c�&�I�.���P���E�>!�b� g�����MˌĿ>ٰ�ig �q�
0 (
\c�ЕF�*Ɋ�!y�RXm��m2��3t�x����+��`+ҋ�-Aq�'�b H�%�p�$m�v�ʐF���ؚ'\�៘�I�X�	��0�����2PgI��̵X�6ГC�Q:*��6��?b�d�O���?�9O�oz���Y�n�9�Ƃ�{F���� =7��mڽ�M{P�'0�i>!���?��fH+ z���0L�'�$Z�|x�́U6z扞R����L���%���'��'k2��M�f�2��$��|���'�b�'c2P��r�4�����?�������PkZ�
����7�2� �� �>��i��7�ܟ��'v��do��,�<ً`���@�Z=:�'�bȓ'l�[�*��e��?��rf��W�8��9����UC���f�׵&l*��������۟L��O�OpBl[R\�ǆ�v��I��-�R�b���Ԃ�<�i�O��Z��V9�v�Q
3L�I'@��:%�d�ڦ�iڴu�����^< �'L��N�.��m���� �-N���:��
1z���Kp�Jy�'�"�'l��'��&�=!�B��R�Jʎ�:��<z"�ɡ�MSg٘�?!���?IN~ΓT�|D�t��8a<*�1 �{��t{�\���4c�F��O��p�����Y�@��|t6i�SK�=_c�4�V��<c �X��#�<�Ө��F���)�����D@��}z.$�ᰅ(6<����O���O��4��v����ra�e�x5��Z�x�����e�yb�~�h���Ofn��M� �i)���r��,����d�1U�X���~�y��'r�7N�P�Hc�>,����?�Zc���
�$Ŵp�m���7u��ӝ'N�'��'���'h��`�U!0N�$J��kA!��Y����O��dB����,�uyx�$�O+�j�3q�!��C·=����j���(�'��6mB����S��R��n��Is��E�*. `YQ� @#kАEQ�cTu9r�BP
VO��Zy��'���'B2��+SXđUN_�	D�H g�B	Dn��'��*�M3+��?A��?ϟB�@�D?��\��HٽR] �O\��'ؚ7MW��3����Oq��2uM��%E��X��Bp� ��$Y�|�H�1�#���i>pv��'#B�%��G�&���yFF6T�><[uED����Iٟ�����b>�'�:6핋,�J��l^� �x)1�`�!��Pq�<�5�ir�|BK�>���i�B���DO�qRN�`֤Q��] Q�x��m�&;�Dx�m���I�=!x�b��֒E�DȖ',�u[��S�35���P`���4+�'��	�����ΟD��ȟl��z��!��2E��ZS*��~�.����{PJ6�i��O�$#�9O�nz�%����L�~\�吅1�P��@��M;�i�����>�|Z��Y�)������Z2^|���L� ��ϓn�0���h��I>!*Or�D�O.a`�K#�.  v��! 2���Dk�O��d�O��<��iS̚��'�2�'�2!B�l�7;)����B�;t���\}��a��%l���?��O�̠0�V#.&����(?����C3O���/)�F���l~2ʓ�ڶ H*K5�����T���������oL����?y��?����h��.��xB)�c��<}� �ҵװ;B�d���U��h�`y�`w���杳+@,*��	wN���e��ShR�ɑ�Mæ�i
87��S@U�5O���'L�01�Y�rX�Y�'����Y��n�d�&�8���<1���?���?a��?Qf�E���H1��3qe$]��X����ߦ�!�r�P���$?�I�%���[7L������rG1����O�mZ�M��' �>P�Ci��us�πIPtaq"�(U>��Riy��Q�U87(H��'S剽?`2 �Ł3�,ԛ6Kǚ҈ ��蟼�����i>͗'��7�،P@�����#A~E8� �3r� �+0�$֦��?�Q�Aڴ'ț�oaӀ 9 ��^�X�煃�/"��G��u.��:O��R9Kt����.�R��
��1�v� ,䴃gdىE���`>Ob��O���O��d�O|�?a�� A2Kof�0��\�9��/z� �I�<)�4S��L�'��6�(�dP�	���0�e�V��x�w��u�49��O}�j�"4m��?��%N�4�.�Iϟ�j2�S"�rYs$�J-?�V	T�o��3P/4DҬ0'��'���'"�'Qd$bY	<ȄV q=���7����?Y����D�ϦU�A�q�����ȗO�<M��H�jJ�5�d̚@� ���'�R"�>ᖵi��7M�џ��|��P�<2���� ސH! = ��u�Q�ԕ(�T@�B	�<a�'*v\ba% ����B��2wc��33�T$~��P��d0�?���?����?�|�-Oj�l�=D��8�-�r�\m�TL�,Ȭ\A�#1?�F�i��O�u�'�7͑�ssT{'V�Toh�Bp �:=nZ��M##n�p�4��?yt�� ��]�5ˁ���'2
(��
�E�����N�<���?!��?����?�-��U�1`���hx�E��MP�bS���XB�c�p�I��X'?��4�M�;r�(Cr��O� ����δ3l25 ��i�7�P�,է�O�u���M��y
� �̢2E��s3����  U��J�5O,�:��W�<p���l>���<���?�^�q"�T�O�h{4����C�?Y���?�����Ǧ��d�����	П��71R����/[0���I�e8�	�Mb�i���$�>�ɤ#���p����  �t��\~"#� ;!iT�	��O��i�7LI�xb�
��y���z4�ic��[���'���'������Hpu`��3Y��٦e[/��%0`�ǟ��ڴ��e�'�7M�O�O�N{���["q����q""/�x)r�:O8oZ��M����.��F����?��"&��H�,Ă<���@S�>xxG�6R�c� �Ľ<	���?)���?��?�v遒3���H0.ҍ29�%9���������ei�p��ڟ�Y��'����V�n� ܐA����� dϷ>���iD�7�WП�&>����?)[��ǁ[�ua�cz	��C�]Da!u#K��J�#h�-���ٓ/7���J>�*O��Ƞj��u�,Ѐ�cD0G	˃$�O$���O&�D�O�<�ҿiB�QS�'_�(�po�7'<���Ɓ(D� X��'��7&�ɾ���K��J�4#X�&"Ê- �h(���g��1*��U~��PY�����y2�'5\5%-K��()U]�$�ӈ�5�,�	f�4p��OS�S��0�I��y��'���'�"�'�r�I�l���扴tp��%�a���O����צ%��&8?I��it�'�&]�@ˉl�H�"s��r�@��O��k}�� n���	�@�����2O���ݤ+F�i�r�<>��T��d�� �P!
�# ��c�$��<	���?��?ARj�$|�|R͜8L�"�"��ؖ�?A�����ܦ�*er���	埀�O]�Di#ȞE� yb�n��G�"(��On%�'ذ6��æm
���ħ�B�Ɗ_4A����mB��3���*`���C�/$^��-O����p��`iD�?�I�2IAi�FՂDf�4���D4C�I�h�>��`�f��X��Կ�.�?!��C5n+�1#� �0U�J;dX�솔������:r�A�Vrij�O�Td"�1`���)c6���撡L��4*���9� �{��L�b�ɫ��@�h���B�Q�-25�Tl�pS<��K4 pUH�V�D�N���D��r��< ��ڗ,p���G*��B6�p�T�;2�T͢����V`��Bǎ9�X���Ԓ���?y���䓜?q���ά˅��{�ސY2�	25 H\��(��?���?9���?Q��?I��C`2a��i�С�� X/:��\�ecڑG��f��>����?�M>���?��Bȵ�?��������g�ݢ.��eZv�J3y���'���'���'b�B��c>�
!�L�<!a�X�)�Ny�Bji��� ���O��0s7<�D�O�dęh�Z@�ƋѠ[�
��*x5,m�ß �I���l��J|z�����������Q����N�*:�'�2�'	����'2�'r�'+��I{��,2\�h�fF
 `q�'�",H�P�#ǅU�'_j��$��o�
�i������
�'��LB�X�4�\k6H������!J�'sά��#�e��H�PUv��eG�2q�=�'�]�U�<���RMbLy�t
!)ݦщaG� v@Ժ��K�vH�3��.b�Y�G��$��7��H�E�*^t�1�L�j7:1/D1j��x*U+fj6㍝3���u�iĀ� �I�F���'���'�T���\�ɔ1�B�#�*e�ftHD���<�D� ��ǈP(UOKv��q@o�?�=��`��"3H�;4C�uj��
�\Ez��`�}: V:1nlC��?�=)ө�e�du�f�'-�nP)O2�?i�jV'�?�i`47ݟ�Iğ4�'���q�qz�h���	U����'�8�g�ٙ/�~Pir�=Nr�X�g,ғL����Cy�U�:�-6޴�3�H���t�[���&r�������I���)���(�	���C�g&I����.�x���f��u|f����Z��d�Q�Z&��<��`рo�z���W�a���(��#/[�E"���q�&�*ϓ.Y��	Ο�)��+:���U�br�p �ē�?�������)
]_������,!��hJ�f'ax��I/N��"��Je��F��o���I��Mñi��	$Ge����4�?�����	@������G� `e�Kb0hpw�O����O�,�� �g�2T'�ʧb](,yU���1�����A�iyH�Gy��J!R9h(���I�HHCO�X��I�����s6�<)w_�SڴN����'z�WRy�	�9x�lA����dy�x�	k�S��y�c�TE13#ōT����uHM-�0>B�x�kS�1TT���Q�Ie������y2"ׄG�r�'�"X>���ڟ��	��L�W,��Mr��+"��_�9�ŀ� Y��ɹw!N�����N�M,�ؓ���ܩx3,3�O�p����+̙Kdņ* �)3�!Liޤ����w�Ͽ��!�I���S�N�0�6����Jl��R����p�v��1��Tڳ��_�l����W_<��d�~����P�'P�OrT;;[q���/��	��CAH��c�����M�Q�iP�'8���O��h����MüX	���x�0�	�'���>Wd���'r��'�2�jݵ��ߟ��ɹ-���hWc�#Y�I`&|����iœfb��4+\Yx��6j I�F�{�GD�Ul�CKٳa˼�������,�p�4WT��>��$?Fx�h4`�h�0낢R��?�C���?�i�~7ݟ�	ɟė'6ɡ�+X�	W*I;[�����P���I�T�)Fx
� ��:!fS��D��O		h�]��F����4��,����gybIP#kz�� '�D�E�F�+���E�Uo|�4��ڟ ��ʟT�%AJ����	�|��%��MPf�C��� e'\ C���=��	�0�֧{ ؈@�$+\O��نV������X��]a�#J3qx��'��$3��-2�_o���	�M��
�0WpmH�]�KY<��J�Z���'#�I̟�?�Ow�L�j �����$M:�A��'֥��l*	�NK6G$XR�'�~���DУO����;�?�����5U�8*�N� �-WǟN�"+��O����O�A��ީr��QȀ�5�r����|��#�2t�q�D'77~�(�_�'R�t��%�4��ċ�BH�V�a�O�Z(���DKx)�Շ�, p���DB�;�"�fӔ�d�O@ʧWv�M:hYp�6d�<|-i )�O���O����O�6�U�$U���ȷ7��hV��<j��q���ē���`d�Z��d����7��X�`"�)�U�iX��'`�S`(d�	��4�	�԰�vg�s�f��gH�<=h�pS� �h����G褍��H���)5�������w����CZ:�R�K��P�ICh�Ԃբyhz	�P,O�]��	E��;{LN��t�IB9��(��+��i��d��?���|���'b���F�/1����M���'�ֹ�Bě�PNu���@e ��yr�'��#=�'�?��V%^��,����%4Y�5��� ,�?���҄ �?���?��;X��O�NS�Z�L��e�<B�� 1���yԚ���D"U���[�N &
̹Dߟ�5���Ø'��StIW�h��	��'��	sJ��w����PGn�z`i�)���.,^�8;B�r��I
�x�k��
;G�����?������W��@��2�MC��?����?Q��?ͻ �� ���T�n�s&�(Aƈ����?�iN
 c��2� N�x���	�&o���2ݴ�?�-O�\*B�U�ը�@ȴ@Y�ő#��'*�^�f�͟L��˟8�I�QH���I�<ͧ	���ebH�I+Q1o�jy��lߎ1�Z1A#�#������;V��=Q@o8ʓ&�^�@å��jA���ޞ%3���=Y0aȕ���_�@!1q�H�C���9#�d�A������YH���#H��`ʆ%�9|�.=�("D�	�o�#'U�̊%+n��q�>O�=��ۺvJ��*wEY�,q��PN��<�P�i�ў"|�Ǣ��6�VlQ�@c�F�����i�<	#��*I6��rK��2�.�aWhEl�<A�括\`,����Ҧ� O�<�w%Z�Z��Cg��s���g��q�<��� /~�A���b`m�k�<��N�(�@aJ��
m� �S�h�<Id枋o2�DɄ�K}�`1S3�h�<�p斢s���K�/��7���� ��e�<� ג]��Y	�dB�PV��°��]�<��-����G�D�z��:A�T�<��E�wF�:�Q*j<�'Zi�<I�I@!� 1�Gޥq��t#��Oc�<�sm^�C;��Hѩ��+E��C�@�\�<Q��ՐOU�EpPƀ�7.,z�.�@�<نj� W|x�i�eN�2)�y�(�s�<����+z,�K`D#:����&QW�<9�J_GE<%Z��3'�8`i�O�<���:#`a���S�豑�[O�<9*�*��� ��j��Au�L�<)f����0�A;�z-qTg]�<��b8�4#���7|����j�\�<��q�\}��'L/[�6E�q�<!G�G��(��P ]��K1�i�<Y�@�g��A �G�]����%
f�<�Q�ҊL�) ��81� �jea�<�ը�� Y0Z7�X�lL�
��Z�<	���!�d\�#�O�^EbVD�W�<�`Ζ�U�����g�6)�d�6Z[�<� �,{��ҰL�$98�`��Ua�<��
Y�8%a�ۣ�֔p0�Y�<����=$���ʢ���;��VL�<)b��M�f� �4.�@��jb�<	 �
,B@�@R�WC���ŉBR�<���s���8D��8xoJ��f�x�<� �!H`�� �hLI��@2j/�!�"O�� ��E���u��E�_/$��"OHY�&����<���ń=^00i�"Ox�S�*	�mx���e"'࠳5"O2i��9J�<L� d�� &��v�'S$	[ -��	��\Ƞ!�V:ĸ��C���M�%�ћW��<�!�����b�K�� �<EI�f�D̓�zm���+5:�`#�a�;t���=�4n�=z`R���cK�,�\��q�	�-��@�\	�R�$�9a61�� o�d��'�= �z���I�yRȊ�hI�L#���r!�D�d�_�$\���QP�y��ހm��ag�W���xC�^-k��$A�T���#I΋'Jpx�̓1>����U�S�8����?
	R���J�`{0�rw�K�R��hu��<�p=�֭��ZD�)"�8k邴���g�6�g	ì��xK�i$�ɧ�$�0�' �9��i��f�Ov]�S�`�6��HS�+��2��ǆ��qA^�o����� �*�J�(��@C���@̞�;�L�KҚx"��#�����	�#�\���wa�lx���4 �5Jۅ**L@s�ئg��M�$��u���O`�i7-U�wE�Ѭ�^�H�Oz@�
��jk3-����q��M#��4�����&\f�:���`���
�+�u����%��@��)*�$�>�D�s5��/�4�7"�)<8 m:cXT�d�Op�p��h.F���ճtF$;��|���!9\m�'�� ��ķ�HO�|�����\.6�
Ń�'� e�Z�~R ŷH�F�YEk�;I�ES�
�?�R}�0eĻ4f���(Hu/�yB޲a�����9TH��֎��?�F!�p��D�T�)mHP�B�R�'p�v�O_�b̹CEU;^Э8�"M<U��yBMET��'�Z��D@�Ri� I�g�eP��1�,��Γ��X�?�u��?��|Zc t��$��%PO�P( �F�$���jO>)�V�dc����Of��C�%,0�Q��$�Z,	�%-ZX��]u��'�B6M�{�JYb�4 ���j�,<��Fv��H9��]-���ѭP_?n�b�x�K���䛴M�ԀD!�?�O2. �.:��-�'*��;�xb%�B Po�Q�Ǵi{D��t�'Okl�C�h@�b�:h��P��
6�f�`Z���~��>Y��?�:��C�#��[dΕ�=�dR'	�J8�2�g��j���A�l�q�.M�
�|8���{�1�D�0�~��Ol�'��S�Q��yaf�!�֤�U	ُ"��	��EQ���`
&��'"��hAX��*6@�>�XU�{�Q6+g��)����]κXۢ�ٯ�~��'����M~D� ��s��K�����5Y�%�#f�D��R��44'��P�H�Pr�E�j��"?9�4O�!�a�5]��
"cΠ��5��2Y�qS׍�� �����HC8��X�Xy��	�.��T H�G�;b��>��'�����L	Ԡ;&�K�#��5�u��?eu����0o�q��(�~��)�M�\�`� �U��I����w6\���~�/>F����|���O��r'�}X�����Zs�U�F�b�	Аxr��%	����9Tc���'��9w�I���9�-X�dr`��'���'Ab$Y��H`杹�J.M�؝�J>���Ì?�,id��<����n>��� Ѳx�ɇ�	V}�&W�4���ɐ�y��-����r��E��)��cɒZ�xZc��E(#�̽^���X���L���hK>���~��)�~�#��@�L�0`F��`x�F3�p<15ʐ9q�p�@���.XM|���b�1z( �͐�f�܁2PHH�M��0}�HI�E�!��\4���ʢD*��i��с����ҡ{�$7���D�x�,Y<\�����z��1�4jG��'�rk0'߷�mJ��ҊIz.���!�{�|�Ɇ�M[5Aߥ0�<�bRh�2��ZwH,�O@Q�'�#Q�DP�Z_�	�
�;�1#P$5^���=ɑ(��~"�^ȼ{���(C%��KH@����D�I��v�'V����Y�,�Q���70C����3�Ć54K���>��,�*8�Rv�J�c@~��(�^8���$B�=kE� �E���8��V7!��d�S+݀��e�U�p=��BU �vq�Z]P͓�+D V�\P���_�&��1��B/��	�&�afk��9rx�
���+J=�O��	a+��u뾼sT��q3|��䖘Y>��'_()�Y�퍃z�':������wY���u�C��n�X�kY.+�s�-�>�:��Ğ'Xʐ<�A��-I'�t��ߛ]�x���#Z��ݐpJ_�I����D��NAp��s�|4zVk�J�^C�6,����蚉:���  .��/M:B�I�I�\ :⇽ͨ�#�J�;3���O�PYC�7�:}'>c����ɣܜ�Ӥ$	���Ԡwh7�O�����,�I23!O�Qp)�b�	�$�vh�f����?�&���t�SP�U�H�=K�l�P�'e��z�K��
/
D$?��v�B8D��(-�1�~�`H)D�� ��j�L(kR�p�JR���-�7Y�X�VO��db��>E�4nѽ$pࢢ��H�Ј@�m˖�y�ٮ�&58����+Ί���NVfL�ל{����bL���'�$Q[��8D���fo�,o�tD�I>�bg�/qtE�E�5�z�A`	]o�Cƨ9�b@�5#���t"	�s9�h2e��so��X�/��:����Ʃ;�jP�u����<�g-2R+\��  	4*lp3	ϭ>Vb!!���!,�� �D�'=,�C`"RY��A��BK��8��
���c��|�45;煐@A�x�C�9�X�Z��S��x�]� q���?F������O�j����O&ݫ���{�Tن��d�4xҁ`"OF�kWm&@z�0��A�Iw��*�hʓi�ę���h�QS5�a~2eUnP\��n�b��Mx09�����
�**��"P���gAD(S4F�/=�d��R��� -;L<�c��	<� Xr �(%
Ʃ��l�>W6 ���I���|xB�������qa�J;z��$��	W敜~�6!���Y�Wu�}zL>I�+�Ƀ���#o�'��d�^7�90XyH>a�Y�x1,O��c�B!
2}2��
%!J~�Bʫ*���&�c�(Q��,��xR�
#�P�yREǴbۨ����Į"<q䚟T�3��&
�>}���a?!���E�ӯ~�R,q�H�p<9�"_�F��|H�đ�����d�GV"��oҜ+x�p�@1I���I�{�e:N�("AcӜ�y�V��(���������H��,�2��M�TOX�an�n����<i��y�_��Du�haT'�8< A��+�X�S ����	=%xX��&�2��d������7����:�`e�<�h��S.W�M����!� �q%�i���(��n�4�'4F��bR�-M	=�±Ȗ��c"��󢯍>%R����,��a:"ʈ�p<IQ&x�h�Vϛa�4�S�D3�"}���O��	2-L ���)�<��>�������`�m�.,kPm.L}����'ȶP���Q�!80�H����e�?p����0&��0�ူ�_*&�#=1��S�y��K�Jlp�� �b�����}��MP�E�ZOb�����V�>���Љ��̜+�9(��!h�pi�w������1�Má��>&��y�8�qT�s�A�H>AwDӕt��I	��r�yc��T4�4\K���|���/?Q#-КK�X���������B��a�D�4lϦm�Vr���69"7d����۰%�J8�@� � Rjf��dF!.��%Z���E 	�'�	��`ŻZm	u3�tQ6�0��wt@ D
��n�.]Iwf�xr�'�4��u��4�$ܛ�O�X�R+<}Gp��G��P �`p�̙m52�	�i��I<���N}H&WM�N�hDp�1&E�8Y�*���(1�'2�T�CAF�b����9O�KU��^����7_?$9Y�l�d��.>���E��RT�U<��g?ٱI%C� ��ƨ,R���#Ġ]��U$����V���``�p\ԂAJ���I�J�"}�I�6\�^�rA���w���ɷhti�a�EWdHhyǓ_��x��F	��m���'C^������gxn����f?��Ŝ\�	���FQ�����p���4$L����	6�;Ǔ[P�1��ԦG��`��@|���@2�8��<Z�!j��<�mZ/d� �T̨{�����W�?�4�X	���%; }҅Λ_b<�іx��w���z0�a��ܰ`�@��y���5����L
�B=i�-��y�<�ɧ&�p�OL-�լ6��#$���
"�
%6�҄�M�6k�=@�Ɵ�`��R�iC	M��Uh�n�|�'�,O����xM���5 r`
}@��L�crd���I�L����q�J0Z4F���<d���A�Z�mڨ6���._��'��q�C�̇/`$����z����է�p<�g N$���9��R�5��ܫ,~!I�CǴ֚��6�"'q�����Ĺ>A��n�I��[�&i�0���ћt̲uJ�E�P�Ƀwi�d� ��a�إ�E*�=F2X���$�&MB��0t�Ȟ@��H�q�ƞ����}O4�3� ���gpfM� �#Y���1��i@�{o�M`�0�a��?��^�'.4���'��P�P�o��D]�^w ��O�y� ��dj����j����"AD�E�0`�萯3��X�R�'�DX�S!
�8���%lE���N>��$��s�_��Lx{���#�P��i�^8��1��A66hiAŦ�Y��]�So[�QYq�G�Dj�0j0�u��ɀu������'1z��ՀR04�'�����$�`jG 8�����*V<A`�4K���O�h��Qn��`;pݫ (�vQ�%�[eV(�ǝ��S�O6@Ic&�C**�Z��Z(��%�w�@Ha"�S
joZ��^ �����OX�%��O�`0v�/d@�$�F��1ߺ0�O�ereOވKF�1J�ҷE�Ze���A&�䌺`,�d} |Y��E)�epa��q�̜	cA�<�L����$B�I�Z�&a!5NU��bP��僾7�B��)Tނ�$ԩ/Td�D���gMvB��6�Nl�BM!);�L�B��'�HB�I;g�p�E��+�v*��VQ,B�	����PƎ�PH��Ԗ,� B�	x�$R�f�!O��L����C�)� 6�23j��z���Ad�3�D�`�"O��2��+q�Ⓞ]!VƬlɀ"O���gd
�ě�C"k"���"O�݃�,�y����0-�0�V"O`ѳ#�]H���.$DE�	�ON!�䍽hp��I���.�\A �C<K!�d�lê\�d܂l�.��V�Ƙ<!��5�6�8����f�F���
��8�!�d�/&Tp���A��W5��S�i Y�!���/%"��&�RU(aJ�H�!�$�
i�B|�2��-�(liG'UF�!�T�ʑ���jŌA(V'�)F�!򤐙^(@���T�nh`3�!�D�5*�EH�.�)����G�2*�!�D��o ޡ�Ьιj���X�-��!��Y|ݬ�	1޼ԞݓsL]�]�!�dK�h�.t�  ���}�R�$7�!��G?!���S�X&���� Y(4�!�䘜I�b-ѡ#��!o�LiÉϴ4�!� SA��p�k�!h��A�M.,�!�D��Ax����%L�	PL�>ug!���F�h���Z4�p����;[d!�Dߡ"(��2դ�P��H���!�$�U��=�D#ԧ�~EkW�_�!���Q���oW.�JQ�>>�!��FZ��z��L�Ӌ���!��t�M��F�iʤ@����"Z�!��6)����N�4���`���!�d�u���Q3,�L�xi��F�h�!�$ߣrr�a�K�1>���J��@�$�!�$��~����I'��0A�-��Py��ժy
Ԑ�d�ʁY�i㌂?�y"g��4ꦥ��Խ;*��aR!�y�TcB��"I� K����R'�9�y�g�J���HՊ>gP,sb!�y��W�C�.�As N�^��x`��B&�yR�V��@��eȀX����P�y��;M� HB�)
I��Ia`�ݯ�y�+�!�8���$Y<i �ǃ�%�y���3AND�b�Z�/� �yr�"�*t3���XZ��fӊ�y�;u�&Q8"��L��޻/�\��ȓR*a0��ݝL��]�@�$�ZQ��@V9���J9�~iK�Ί�(.���ȓH�L�1o��{��9c��P�M��T��T�h�� -����cA��?�>=��D`����U�ۚ�����O��ȓ�U��gV�;�v�IU*EP�0B�I�/�������0G����v
Ι#XC�I�WL:U�$6��(���Mh�zB�I�;ЊeE�b��j���0ˠC�I����AR(��������()��C�Imz�TÀ�ɡ+X��5j��k�PC䉉_�ꌚ7h6r���1^�`B�	5a�z��ƠX�uq�ieƟ�*B�I�<&�}y`�O �x�Cu큸V\�C�I�����1$��zrԻD&�E��B�	%uR�A˦�C2V�^��t�Y-Vl�B�I�.F�X�,8v��<"D��%��B�	�d{dX{t`@�Pz� �Ʒ#�B�I�&U1"͡sgv h��"HH�B䉛h�t-Z�+5L�zCP��0N�C�I8	3���s�֙\�hI� 
�t��C䉿`�� �7"��"GVE��
�<>2�B�)� �@��ȱ,�&�!��T����"Ob��dNM
UH�A��"����3�"OjA�Q�3�*�����7�ę"O�u�BF�U(N�C�~����"Oʧ��'�@a�$̀"q@%��"O�%�U@�kޖ�����>Z6(�Bf"O��"��z
h �q�Gcz�h�4"O>��b��\Fn9.qy��a���y�(dW�A� əO��l�"��y�I	6����i�!F�{���y�l�15|Xr�W�p�.=�$����Oh��3m37��M��iִ�*���A�a�<�1�ʃ@hx���(�8,��i��[�<��O:�@��ԋ�27�T���Ip�<1f��*-*\�������Țsm�a�<�f�8�BU0�G�QjV$�\�<q�K��J�*,(U�ـh��� �V�<y��ʥA��(2���o}>5�MI{�<Y��فI���n�8i�4ٻ@H@�<15G�)_�v1c�ߜ?�6�cr�c�<�Z��~��&��$ͣ�`�E�<yE̒�P��9IfP/F��ja�H~�<�sӑ%ߔ���i�3u�̌I���x�<A��/!�<)�FD-��%��Ŏv�<�%L�%���5�'qfn���[�<��R��BE!��I|�t(f�DT�<aF��uO<��J"�r,"�O�<1 �._��s�BV!���c�D�<�&�J�-<|�
#�șH~�y[H~�<Y��D���"gN_���Lc$�}�<Y�%�!R���1��^ �ic�AC�<�ė?�R	�aG����� ��S�<Qb͊28SB�����	!K�m����O�<�B5*��Q��N �P��K�<�d��1<(�&@��
�<��A�L�<��B
2��၃�鰢�K��hO�Ob���"�(��,�V�N*i,U	�'c�hfR�hdR�g�%x����'��������ő�GƼ�'TV�c �'uVv�X4�ͩ���'���r���*���dΎ
[��C�'��䦜�.�P�X"�2}��0��'c4��ĩJݚ�"���>uM���'\�zCl���V��v�T�:�{�'g��D�S$�xB&�F���
�'�ٰ䀅q�4��	D�Oh	1
�'��A���Ӂ*Р+��ο���	�'���Y �4P�C2�T��L40	�'���V�498P����P���	�'BN2q��(��U��WA8&�I�'24I2U�6� ��?�*�Ǔ�HO:~��T��#&k��*�^�M!��x�zY�� ,b� !��ѽM�!�%vX� �T(�fy�P�͙�(!�d��+�К�m�Ԇq�RƐ;b!���A�L������|�Z��a!�d5P�d!��NQ��XUb"�F?M!�d�<O,�a�⎐;����!�	�<����
!���fɵD�!򄅺YE��(�ސ�m�&ؤQ�!�d]#p�\m��aH�u��'�L�!�D�!M�2�,��,�����`F&i�!�ʱ
���"�>v�
��c��~�!�@U*�`���#|�ykA鏇l�1O��� �i[a��X�� �#�G�H��CP"ORL J�� $2��A�b�HB"O�}�_�U���	S��q��"O�=��n�����%��>�Z"O�=�C��,.L� �o�.%�;"O��bh�2�pV�	x�"5�Q"OB<�"�Ɛo�&i����t@L{S�/LOp��CF�)p�d�smC�m�5�&OP&cG�$��`����$���K��D�<���7��۰D��t����H�<!j:uND�'��'G&�-��D�<��_�J�Q�&ݸz(䳳�H�'�ў�'iR��xfL_/V4�Qd+�H��QI����aO+6�8�I����(���D3N5�veQ&CPY��S� -Z\��ur���#Ã �JEDҒ|�Qn�s��_��>�?�+�ӤKs�����N�j+6P�"O�]� �Z"<u�@���r"�ݩ�"O4�r�L�R�R�a�R	l���"O�!�τ4i �4��V�f���:7"O�D�C��'�j|J�A^��5S�"Of�1EO�i���"�j�=��} v"O���턶'c�M�S�	Iv�"�"O�M���#՞��db8�QD"O  h���\j����n�+K�	(3"O��y�d6`��Q�e.�??1���"Ox�;�U.�B�M51-��A�"O�A!�"P;�2���K |�Г"Op���A̅U#ޕi	�~��;r"Or�hQ䑑p@��Ӈ"�L��Q�%"O��aߡ�έ��@O*�B|S&"OH���X0����9W.,�B"O>aj��#6Jd ��#S(�U��"O�(�$hB�>e��P���a��es�"Oh�s�g5Ǡ�[4KB)d�AT"OlA�'���s��Bc��2���W"O��)f�]�(�P	G"p(���"O\��(�P<z��ХB�160͘2"O��XꙖO�ܒWj�s3���"O��5΄8�0�����1� ��"O1��DF(]8r��� .�p|�D"Oy8%';��)��P�t��(Q�'䑞��\P#0�b*Y�)���:!D����'�l2M��ݽUR��S3O?D�DA�E �#�La�� �G��
�`:D��۴hH�N�<���Գ#M���o-D�lb���f7��ՅX$P|pL�֧,D� �3&G�N�aR��g}�<;��+D��Z��܊\�i�" �E�� ���6D�DӶ�ј>7D����������5D�hq��V
c���0�-۪�"�?D��q���
P�"mic��]P�t��;D� PE$��_�[��.*ER�RU�,D�d��&^eH7i�:���"�J�<Q�.��,I��QGf�b�0r�˝D�<�� A�g��X���?{	�����D�<�p����v�J��}�6�2C��E�<��n[�Ir�3�F�>T���z�M�~�<�3B؀l�N��U�[��P�JdE�e�<��/@�@���w�λM
�1�V �c�<��	�*9�٪�E5����E�d�<).ޣp����_Ya�I)�L�_�<!!��Td���H�S�~�X�@
Y�<9��?���o�T�`I���T�<� ���W)�:s��*�>6zx��"O.Iڀ�˫B	�lJ��C.H�d��"O�=IV���n,��ãP�f��C"OҘc��[d���C&�	N��X#3"O2�A%(M��Z���#Y�����"OR�02��1 D����۬I���"O��ؒND���|��6 ��9�"O��#�/_J��Ղƙ{�D��"OJ�C�"D�6���CS�b���C�"Oz��d�l�>XS��O7]��;U"Of�S��9(��4��c�7u���#�"O`���!UYH������6�	�"O�E@���d�Ԉ�7�U ����"O��H���#VO�@�''оG���W"O�EDJ��A �e%PWo�� �"O������=�pa����,�V�� "O�@2�%@�r}�'��^�xA"On��5�I�c���؃�&K���q"O� �@�I�����KH%d��}z0"O�0R����p�C���( "O�D���҅&U2�r@� �Uq�"Oz��.]�б��V.u馈i�"O��{�L&:`(EA��=���"O����lϮX����H�6�
�!�"Ot���9 ��0�5�39XҐ�5"O*�i��;�2���L�-Kv�9�"O(���P�G���!��:Lf%W"OxeWJ�o�� 6 ƥL:�``t"O���/����r��+��T"O����֜6�!$nh�a"O}�v��6a�q�%d0����"O���r�I�9��Ĝ�	����"O�q��<]>��f-[]
�]�#"Oȱ��ƛ �0������8�"O0���C�S�"a�Toцقd+'"O|h!��A\h�����?� 4zb"O.]F��.:�x���M� RY��"O��B�̯C��1X�"Mlŋq"Orh�q��3T6�m2�G_/�9�"O�T�t�J+ZG6͊#F�q�����"O�4��� g� H�H�4�2"O4�E��"x�a�t��|���`�"OTH�ӥ�iҜ�HХE�{�F�a"O�c2N�2��%�
 �DD��"O.0	E�He:j}��Q�=�%"O����A-@*��6Io�,�d"O,e)wO8WP~QBG���f�"O����gw��e�0i���
�"O| ���:U�b�� j�Bȗ"O�A&L�Y�Y0��� .aÔ"OD1Rsf��!a�Zp/:;��m2S"Oکb .�q�
�aQn�,F�NUI"O�T�4E�Ru�h�0��@j���P"Oe��+���P=�s��w\D�r�"O�\�5�4G#�����Y\�|��"OD)�W�ɔ)P$�ϬH4*��"Oa�:����ʔ3n 6�6"O8��œ ��yGI� /<���"OJ�#MƉ.\jS�F:KL=��"O�LI�*Z�<��DH�
h�K'"O^����9ONh�Z��_xG|q�$"O�=�霏]��R�D��jl��"O�A��"��w=p;�N��~��c"O2�v���بr$��{�,-{a"O� ¥�$��.KF�	�Nu\D� �"O��1F�ss��k �|�̱�C"O
���g��b-���2'��]�~�Jg"O���u�]ز�@2&J6h���"O�a�ӁRY����*���"O����iϩyɴ��!�>�<m�6"O��$�[x�����S�֬$�3"O�� p۞��xc�'p��AxE"O�Hic��wӤT&LG
L�����"OP�Q��Y��Ԙ"�ي2�~`��"O����/7S�"d*�0v�`�"O�i�!
�%���GH6
R"Ov���� �R����	p"Ot`b��m���J1`%y�8H�'mAˢč�u�N�F��'n�Y��'��4kB�p>zX1U�"Nw���'�����횥z..<��쒴4tq�'q�#���3 �� ��(2�3
�'F�d*֩�-�
(@�W4%@�UB	�'`x00T�E�Y�GbK�f�r��'ȸ9���	+"������ZE���'%4�,�t����I�)7y��'.�"LR J^�����2�ݘ�y���g�s!�K
n
��_�yҢ��<	���.C��� ��3�y��#5Zn��o�u�i���4�y���9H�^)+��6��@�G �y"�R�3x<�aǴZ����A޲�yR�H]b�0��k�OL��e��1�y�5V��ɂÚ��t���Z��y�N�4PD���@(�`�  ،�y��]�P+����8l��ʔ��
�y��)>D9"kŭ-nH0�`%��y2nA>vj�Թb/�+�MhcP��y&��dm�%ZEŘ'ldU��i���y2��J<���O�2��8��}�
�'�r�BԐ{���B��#� 9
�'k�F@��
��]p� x+fe�	�'�f 1�T�tξ�&����,Q�'�L�
� P�T�����}4D��'D� J�eǏz ��U˙�^(͢�'�\�cå@E���%��3v��9�'V�H���ŎV��D�%��r��x�'F�%���\��8+e��-i841k�'L<�Ц�FI���c�b�����'��!�c����I�n��[�l)��'�B���b�Gq�qr%���p�P�'>�8"���F�F` LE
��S
�'�j�XҭE����	o�*s�Mz�'��	���4r�G۰_�@]�
�'��L�Ү�8.D�H��I#T~z �
�'^�`�� 7?x��5�R @HM(
�'P\�'��<kߺ<p	.G�Ru1�'i���beQ�Xf�@�w�O78���`�'�Hb����`�i��MM6Z��q
�'��
",�-|�@�"�녱V�x��	�'�V�˱�B�}��7U� �	�'�����5(&.mC��7����'�DLz�|ITq�΀��Tb�'�*��!�I*`Q�lk�n���X|(�'.T�r�#ٚ]v��Ʉ���i���
�'J����nƖ~P�x��%��P^�,�
�'���`#h� ^��K���<|��p
�'����aʕv�v�cAmT�HT��a��� �ř�:1M`:"��n|U�U"O
#s X�!?XP����vn���W"O�42Wl͐|��T2��شW�
�j�"OV��0��v� ���6Sw\�˰"O�L�hX�I���Ҳ^n�,x�"ORpʳJ�-��jTC��Zb�`B�"O������D�Idٕ  �1y�"O���֨�\F=j�@��'�l�	"O�H�uA���Cg��5�d�q"O����U6N������A��M��"O��A b1W���%�"|�`�q�"O����U�M9�
^�,��E"O)���/s��yc�i\�"�b���"O
��&j��,�1#��!v��#r"O��P�+W-	VYZS��^�H'"O�UQB�S�@����SH�tx3�"OP��Q�>m�\`�K6�<���"O��As⑮*����D1���(�"OX�"3��(�<��cf�a�D+R"O�@J�+"�,�J�%LF�j�#p"OVM���I�����S���8U"O�� �C��Zx,q�S`O�=�,�"O��0��X�h)p��Qe���"OY�F*����Dst�%\l���"O��0�I�yE#�G�幵"Oz�4X3TAd)h�F�d(��"O�H� 
T2'ڎ�KE���r$]a""OZ8#s�5O�L4�5�_�S�$��"O������&U�mq�Ax�؅�$"Ojl�$.�(g��u�DO�2���"O���Gvm
��#M�;�|	+p"OP�`�²u�@�R�Ŧ��9i�"OB�H���`K6�Y��$��"O�p��ʣ3:��r�@����eB�"O<QP.A+2���q e��V�����"O�}�%lݹo�j�z0���F��`�"O��#whU�s���TE��J��"O�h
�gY=D4�hB�ƥ>�pUyf"OPՑq�Z��0��E�n��i""O朸�`Ƴc����!��d��"OU��*qZ��jp�L�c:��[�"O-J��;A��]�e�K�y1��q"O�P�u�*�^���I1]���&"Oxi�$M�n`�,�pH�T,��`�"O��塝�yx��BN��\�"O� 2��-vO��x@��?���R�"O��Z����6�<	�a� e~b�5"OX����'��P�$O�/R��b�"O�%���M4i^�0Ó+L�H�`���"O��#���DF�CKO�g�,|�"Oh�Kс�����CG2��0"O��3��kLB��C�Ak�zl��"O��@`�,p�!��89�1�"ORer�"5>�J�*�82З �ybG�9^���U'M���)�L%�y2I�F�`|�GR�@kb���`ڥ�y��ʘuf��q��Dyh=A@fA��yR�!w���2䖙>��E@)_��Py�FM��RĎ�5W������d�<y��Ý'��%�e��)d��X��Sw�<ᣢ��;_�S�J�	4a��h�GPp�<�#-Asr 0��_�2U�2F�m�<�㈃7xNA#�ARS���S��e�<�"F3H2�H��*�>!��yTVc�<� �x4��N�ư�SOެ78}�Q"O���`��]���@n?N˜4 �"O��:��D��r�(�B �*�A"O� ���hR�9���%O��р"O��&���DZ�A���9@�ș�"O�9 ���I�=��G�\Rl ��"O �����-q4�R�.C~�"�"O�eZ�LXdG~�!�ƻ< �f"O��Hcʇ#�@`���$q�F�X���O�d�<)����IY�P�qc$��&p]���e�Z3Vm!�LNQ�xz��͊(<vL�;U�!���!�@L�3DBN�����3�!�dµ^��y�!�j��i��+5@�!�DV"d��͟�t��x"�J�_]!�D\M����T-`{d�%阯RN!��۪��O͂|���3⧈�%�|�D{�T��E�t�&,��q�-�>]K¢A��y�HM���,�SeDot�"���y�(_�(�x�Hc'Ʃ{���VnK$�y���9\A���N}��%:����y�L�Q��ʂ.�m�α�5e̒�y�,_3U ��dGֳj���ÅN���y�dˋb����cMM�s�5jƪ�yς9t�d!�'� W����ŉ��y��O���!�aKV�H؀��B��yrE�<�@�(�S��ÅB��yB��qTp ��UW���Ve �y���Q�q8�F�8K�f���
[��yR�M�\6�0s�/>�2	1�Ѯ�ybW�9��(��H6���d�6��=)�yrmS�u�j���䎐0ư�HSO�&�y"�P�"����˓�s4��G�&�y2� )	�Hy�PBH�p�
�����y��\�c��82-��G�rؓ�BQ�y�`Z�HR&�(�ݰ6��y��C@"��D2Db�:�o���y��5>�	��|� PCp��y�#��Pw4���J̅E����d�K����?1ӓ:=�A���2�Ti��7&�1��L��e+�+��<�k�Y��ɇȓy����;T��œ�˚����x��@uƷ(2�L�l
�`���-\AP��d{<#ӋW/oB���V�����ټ�6�Z�ń.����e.� ��`U;���{giF(m�!�'��'��@@���OkJLZ5 ��F�$���'�n�p��d=�s�K�m�N��
�'N�l�e(IF�b%0s�qƮL��'?6�nҖ#D�L҂�_9o����'9"�a�Gѻ2��۲mƱa}�m��'����A#Ҧ"�z2 �9	��S�'�����m˟q���	}%P�������?��L����4<�a�`E�0~�|�Cc&D�0����Q�T˘�YB�@1f-%D�`fn5"�lT����)[��4{b�$D��ǧ,�hiР,�c�)a�%D��׭]���)#BűU2V�Ѵ�%D�ȱ�k Gi��e��y|�Kԏ"D� �pc܎>���Y�+�=uz��0��0<A�e��E~��#�v%����m�~�<1"��M���[�l�	v������v�<Q�	����ƨ���P
��f�<1�A��f9R��ń^�NO
�I��]�<��*7���r+��.���3j�P�<� ����#Qx*aэ<W�p�"Oxa8$º���'��1g�5�!"O�|�%�^n�|q�DN�Nw�A�3"O�<�gM5I)�T� %Ms4�:w"OD�:R�]�n�@��2�W�^3�"O� 0�.�$NU��CJ��e��"O�ГT�2e��R�=K׾��'"O�:w��!Ixl�qgR.$?ܰHd��-LO(�1D�?~�(��ő�,6���"O�i�/³i�����Ma0 is2"O|��&莒y��Y��5&�8�"ONy!7�U:bc���ë+Bš"O2l{#�D�Q�8�F�b��ZW"O
��/�	��H�gH�̮9Xf"O�h�T�ٗYK8���iƸ�!�"O����A|�Jᆁ�D� s�"O�K@�&d�0q�E�*T�z��"O�m{��_�I�}J��YI}�hR"O�lA�Mɼ@��<R@�Л-�ŘR"O^m�Q�Un�\p�)�>d��]c"O������1�N%��n�ԙ;"O����ʖ������#��=X�"O&��b��5����7'�*T҈)+"O�=����BW�=x�L��0��m��*O�!�a�e�lA�I�T`��
�'�1�$�@gΙڥFC�@f|���'�$�:��<v�F1��H��>��tb�'V�!�.�ms���V΃/�N��
�'mx�7��V�Tl��
(xs��V.�rh���L=sRt�3aӣ;��O2����H�*������铆`�!��2��	�b���2��[Ǎ�L�!�O6�x��3�٠@�f%E&�_�!�FE��`2i20&\�HcB�0om!��7w
��5�(2�~p�K�Z!�d�'�$)�.�
E�>�:���:!H!�$OҍN9Jp��e/�(oD!��"?�Lq��&�1\�ĭ"�n,�!���`��#��Du&y1#(�E�!򄅝Wu:������9cnݡ�̆�!�d0o�4����hID�� �Bm�!�J+t�r�@qO�QFL�r �\�V�!�Dn@ܜ�BE�RA.mZ�Ϙ��!�$�a��pY .>f:Fȫ!HD>/n!�d�B2$���\�M�E��xU!��Ts�Ր�LK Vڝ`��x�!���r��A04�T7��\�!kؙV�!򤊂IB�5��͌lQZ�I����!򄁀 ���a�LC�����H;o�!�L�nUrpG��oA�uc�mJ]�����;fћW"Q���Tq�jX�-*B䉒~Z*e8��*c=f�rs�ׂD��B�I(;�)j�	�*Z@Ȧ��
��C�I�2�4�ᗁ��=CbX�3�ֵY��C�5:̸����V�
�@�u�
]PB��:=� ��Ն�)Y���/B�HUBC䉴Y�d�QE��v{T:ah���C�	�%�>� b��Am c�aJ�s?"C�I,�Ơ���ܼ��ERP�U�!hC�	2,�!(~�y�T���a:�B�	�x�.rp�����I mC�B�	|$źG���O�bA�B��7��B�	% v�lH��٫%�X�pn�!Ba�B�I Vu����FUH�`_�d$B�)� �1�gOK,�@m�fB��k���"O�aSF���NvZ$�a�
1<�qT"O:���HVU� "���H�z@{�"O ���j�G�$:Q$�Z���"OmA�e��҈)�ޗ]�z8�r"Ol��cF�6_� ��݇I�vСV"O����L !�:8�@�5r��в�'��	,z"�t!�GJ�9!Fb^	A[B�	7^G��*�R�w��1���*u��C�ItY��QE`�I7��뱏1'�C�	�}OЬ"PA�q��u�ٛ%%ZC�I�t��(A�Rc�%���7 @C��N������N؈0Ԏ�X� C�I� Ϭ�1�&��L͸� �b�C��%��5[���,f8m!�����B�	���١��3jy�L3�lP�I�`B�	a���bť��#h����OQ.6�&B�s�:�i��J'=S�\)t�;�B��ض00�=��)1Y(+	4D�<��䇤�`����v����3D���oZ�~3�	�Ҝ3�:-c	0D��Kr��N���2r�$º��r�.D��&�� ���2�*��]
���L8D�P:%�	�,��R�c�C<���*5D�<�lNkX9X���2Jh�t�4D�+Â&~3���"�$5y�ha��4D��!��ȸ�A#ʫ^o4�:��&D����֑Z�b�3�Bµ&�4��%"9D�TЃI�>�ܘI�M�<#4x���,D��p�L�j�^E����;4.��7�=D��P��Z��+�Ĭ�!� D��[&K�:���2cH |����=D�Ԩ�B�~�YS!3�Z��q=D�l����@�i�Vl��@m�h��J-D��X�L19�0�ʴBȁ(�-9�0D�`�Q֠A��c�h~�D�s�9D�@��$�0r��c�ĆG�|TZ�K4D����ON1&f�ZC�
G%^ԡ D�@5�D�;���sLC�h� ���>D��2P(,Bd���@�s��X``# D�d���P!��cfM�<�$�0D��������8��ǚ'>P)��H;T�t b$E8x�*A*g�ǡi�4��"O��d^�u$$���KJ&I�bi�"O��R�C�H�0U!X�N�P�X4"O����CD�$P@�Qij5��"Oh-��%�y%P)�a�B,���"O����[^Rxqڕ��g�,�
"O�0sEA�&i�F�:~\((��"O��{*��R���!��	��#�䓋0>� ��	 ʼY�Ь�,�~��sh�{�<����%Jdl�ulKIA�M�7�H|�<��䐓w���5�ƹL��@g]�<)�o��dB*����n2ɡ��\�<��(T(9âHF0Jhٙ�b�\�<�����h�(�PH�d�����n�<9�
��n�`j#d��ސ��ʌc�<ٖ�߸x":���eY�Wr<���Ft�<���-�V�(S$A�K�|}�$J�m�<�CHכ>��	c� �`���e��g�<)��ȹ���S�#ܖ$  RaZx�<A���3SD��+�9������v�<�I��O��� DƬ�IS��r�<A0�E5J�1����JUp�<� Hd`�O
�:C���ի̚*E�1PE"O��y��e'8���
}1���"OI�U���.��ւ0�|�ib"O�iK� ��(�ASR�"6'.D�hsC�,h)l1f��uS4�) *8D���P�!Tw1
�O��`D�� $7D��Y�K�z��8��� N�E�J0D����1�����S�s����f1D�� s��)W�v��c.SeW�9B#�0D�|#0"�>�����O:�
�#�`.D�p�M��,�@����+D����$+���J�+K6X���(D��bT@˙7���(mߚ\���RG'D��1��S�R��d#�bS�?��	�j!D���׍ TJ���+�dM�!�U�<D��që����lH�E����B9D����)}Wvg(�:!0M�8D�`���`����#�\d!�ҋ+D�T�'nɎj����MS,�R�C(D�tr2�Vq!����G�!E�����*D��w �e�6Y��K��&�io#D��8����)�!�@�( �Ĉ6D�H�eY�.�� 
q�Fv��"H)D��c b޼N5��JR$��L"<U���%D�ЙQ�9A��p�@�q&I�&g#D� (�K
X�a�FcA;YH� ��@#D����Q�����B�.��`���!D�8�  -YJ��H���A���!�L D�Ha� �d)�8�d@(0~�QD#D��)0�./����v��]bȒe�?D����ɘ�'��J�͙�x�V�ӌ1D�Xx��P�&B%��-8k<L��-D���Y�>�"�:A�L�Zl2@a+D�d��*�^��!⇓�R��bB*D��z �����C c�7C��#�'D���4�XI���t�
fz�07'D��h�l�hr4��+�2 �ȸ�F#D�0��jH�w��d�+w�ԛƊ!D��
��$��M2v(�3b��̺g�:D�|ȣ�#;�08��φr�V��&6D�P��8�p+�b�ga"�x33D�����m��JZT�ڀ�CO2D���'��C�����9g�X��N,D��#�#&|��j���E��4��'D�s�f�!>hQ�E� xp�՜5�!� M���{�)__�[�㖠_~!���`�X��`˔UJ���>c!�O�b�^}��mX����*G�lE!�d܈Gj�{휌[U�e�۩_@!�Q�M���@%v���h�뒟8@!�d<`>��a���}��dP!�DH��I�O�Ew��CDM֡5k!�)x�4x��A�*>o�9��ՌV=!�$ =���W/�*AWjY
�_�E5!����*q�6�7&r���GE�8!򤎠)g��F�
OV�#��8�!�$$@�m�skۓ
���!&@;q!�dݨ��5�#Q�XZ�DU�!�F=8� � �M��{t�ԣ I�!���;A���Ea�:�tLk�hÂj�!�d��r<8k�!F�,^q�b��!��o˒��թD +���AAːo!�]b�p�a!/͗y�"��ϛ4#y!��iM2;�J�����kR���dr!�� �j7䊈���r�
Z�q>�A"O���s�1GC���S�e9��kW"O��&�Zevh�C�.l�"O�][�&Z=&ͦT��!Zf4��"O�Ӱk�bk�d���\��Mq�"O����W���̙�h��R&"Oy�Q��b+�
�I��*���t"O�I`��h��y&)Td�
$��"O4�@��N��]�D�F��؈��*Oj0ۥ��]h��m�u��1�
�'T��㛔>z�qp�BH=<� ��'��R�H�i�"9Pቆ�2��
�'��\�i�!B��j�ć)���b�'ONY��DJ����S�L<p�j�(
�'p��q@.I dc>̃p˙0jY<9�'�8���W�:h�0�W�7i����'J^�S��277���G&Pg��	P	�'���"���*l���6b�0Td��i	�'z�L��R�sqq�'�G�Om|-2
�'#��z����+�%MRY+
�'�Qd�-!ځ�$�\��(
�'�������H��Tï&,@�s	�'���1�ל!_���Vf���'H�)��l��ƕ�ӧ�;�@c	�'O!R��N�k�t����_�/*~�*	�'���� �?_>�a�C��y�F�.c��1B)�/b �TR����y�k��3�X�j@���[18�l� �y�#��9 "-���V|]�Á�-�y"�A9r�X��&8Jв����ړ�yN�!��5�^��1��G��yr�W���)���H�>��c��yr�D�%�X4"�#���oO��hO���L0v"Hx��C\щa�ۼ�O���ϊr�օp��õ���g��_�!�4K'��i�Q��$��!v�!�D�-H����B�mڀ� �|�!� )}�ٳ�	���4�*�n�)5{!��_�,|D��QO�
�� ��ա@p!�dtOdكe��|pP�7�Ԕ)�!�[�k'6�0&OB2f�����
{�'�a|��F�I�<�bրV�[H���d扃�yBH�	_F���σ!(�t$A_0�y��1;����u�9gd1nK��yb/Ao7�<�Q`���t�ED!�yr��6��g!�����P���y�.hO����g�z���W��y��G�\9��0<�����ٹ�yb�ɏK/�KĈ��xU��;e"�y���,e倌	��]�]�2i5����y��'H��I*��T\D,�8ae� �y���㢌�֣«g�-�@N��y�I<0��r�%�cM� R����yB�ߝ] �E�`����Íʱ�y�&�GL*5F�.%����m���yr�ur8`[�ԁ&qi2�d��y��A%khȬ�6O*#(�pN��y���D�6����ջ#��bG���y�D�Q�l�E�]8"悽�'F��y2'ن'�4�&�#����&
��y��D@��W̆�Fo�7K�$V���~�'�0a�:Re�X�䇚�:�9��'��U���O���!���p��!����&���'Jf��!��!s�FuKr�܍9F���� ��5��N��T�d_�{��A�"O�a�����z�BvD,���K�"Ob��qCV9~ ���68sr-*P"O��sp�<L��ԉ���Ljt-��"O�%+�f�a
mۆ�K�%~6<�"Oh@��nC�EmX}��b�4s�T�b"OB8ĥJ!tob�r%��wr%��"O� �p���~&�@�RA��*X�Qt"O&����^�L�`q0� ^�n�!�"O^�� �]�&݊qb�M�u.XZ�"O�������sƪ�N^4ܸv�'����WAA�}� �5�Z%rл)�<Q�04J�i2ϑW��ͩ��e:�,��J��!��O�qi��H	Slb���ְ)�.��sw��`�)o&l��o�(��!��0
80�A�U,�@��#	r�4���$��HA���A��A(��P&�%L��,a�O)b���D{"�O��\K���y/��� �Z3���'�
�2$�PN�F�!QcM>GiP���'��y;�`�Cr,<�m��k�������Ħ<�	Ó:`��1r��<��X��b��MT����R�T��T&�
`9�t���#,����nD�ȁ��ܔ��B��L��P�ȓ^-��2U�_=����P��T��|MĤ� .��Rm �gF�p��`��j�&�I$2��U��6��2��IkGn�6؄�˲�^@r!�ȓINȡ�D.ʃ]���� ꛗ,Z^ɄȓT�*@�2?�2�z��������-�D��]���"��'c����Hi�\��ܼD�f�� !�!8�D�ȓ=B��QMZ<�8s��6t����ȓv���ugY�y�d-X�65�X��I�<	Ձ�e]�p���$�so�H�'��y��T��?�T���(��+�Ν�F6D���%O��� }���=eў!)�6D��T��'M�2q�3%Z�6M2e #�6D���Ʈ��U���qb����9��K5D�#�P��������KDc'������P<���C�W�^�p�"O8A��j���$�wVb	>=�"O�9����i��i*�M<@�"O�9�1I�g#��"(B=i ʑX�"OB͠�DȌ:��v&_a�&切"Ox��Gˆ ��2`�E{�<t���	E>%#B�U�\x�1�	���8C (�	Yy"�'a�OZ!14��0�<�I���.�ڤ*An%D���E�l��l���rA萘!�O�ʓ��D6O�q�`N�/�ưI�O�H�Z9��"O�<y0`�+RH�X�%`^�,x�r"O	� ��iN̺�Η,p���QA"O`�z�m�h��麃�����Q��'��l��L�1�떄��W�ܙ �j�<�����>�ӓF���+��J�V9�ch�Y$�B�	�?'�u���B�L��5��(�hB�I�.�`���"4f6�ŉW$Bv4B�	�9&��P�� CQ�(1&�V�W1�B�ɷ��c��K.Wh�xʡ�Q=�B䉟|	F]���� �l��̎�w��B�I�X<j�iH�%(�X8�EK2��ԅ�I�t�Ľ3���M@c
��r�����<���ǖ;���cČI�?:��A�؟8�'#��͟XD|�� �)���0RUDW�y
� r��W@$\|`dC�!��r�"O�:b�5̬p��(HV�L�#"O�i�3m̿Z**�E%T�ud~]�G�'�ў�'��'�h�1�����C�
�g�������Ob� �<9��+y�d��̀#8�B2��m�<9ӆ\�6��,+!� %����D{���K�f5d�q�˙n�h*0���P �B�	�K���@`P�9����b��B䉽�R�u�ς;h�+�X�7�B�:����*=t<d����֣~7�B��v�h��F��tl��|̀B�ɚuҘ���`�^D��C�}�>C��R6��K��E@�4��f �<�B��Q�R���hW�:��l�1�W��B�ɭAĶd!fF¾r]|���%{�B�	���� C�
5�m�t�LX�C�&��q��N�%��(�削}�C��+?���l�%�y�R��-�~a��R���a����X{����gX��S�����O���x��ʂ)��P��J+��E`ӫRq�u��;m�|��ȓu�\@k������RaN�arn�ȓqz�&�	�x�J�1) ����L�|1�m�N
��I1����lz�qk����*} �VOY��>@��:2|`�Ca�7�xT�' �tD{r�'�Dd��H�Q����F�6���'C����,��f#`�a�oJ�TG� x�'gH��6a�Sg ѯ<#V�0��1D���$錍K@-�edͅQ��S�.D�Xz"�R/o�dQ�"L�DR X�a�+��0|�A��`�p���;;�_Q�����O �e'�W2
$h"��z��8Z#"O `�B���v���a����"Ob�@ ��:�|ћ�iϊM�&�qU"O5��K� � \JRh�>q����"OX�s*R �eIaD��9�`�{"Opa���Y�<�(
Ad!t�آ"O�Dr7%�91^���
΋&j9�"O�Q��ݱ7�I@�Y�R�����"O
|�U�K�$*��6�YQ΍S�"O^�`���_� ���f_#7?�9��"Ol10��]^�2-�F@27:B� �"O�|*�.��'dܜ����"7H�P'"Op��W�\��L�A-C%F�)C�"O
�X`�".�JE*mL�0��d��"O�l�i��&�������&i��"O�Hhb�̕Y!Q�e�H��*"O&9��T9i�Й	��Я'���fV�܄�	�|�`�惘�ǐ����G��B�I�E� @���$�f*�{<�C䉛l�n\�l�3���I3";$�lB�IB3�M
C�<8��/��f�`�=	ç#G�t ��C�3����DmE��jy�ȓ0e���!kܘ10Q;��>qs���ȓ�`p�#""��)�n� \����ȓN���£���X�\�q�Ô \�I�ȓ1옽{R嚩KUPDQ���x�F܄�P��4q�� �~��s�ʳ$��4�ȓPƐ\#SkN��c��PAF{2�'E?���*r�0�G�$�f���V�?��'T�������"�	�xD
�'��<J%�0b�T�J���v9LEb	�'������	3(�=ib��?k�L{��� ��x��	n�S'�V26v.l3�"Ol�!��_F	ٹDK�.E�<ٴ"O�3��P*<b��P�h�H.�4 r"O~I�"^.Nq�ؠ�"�)����'�1O�ěa�^:2%�5�B̾xt=�1"O i��a�:1�<�B�C2�:��"O�\���6BD������;���ȓ"O�����)��u�ɒ�x_��Ё"Ol)�R�G��!�cM��N�	�"O�xj��g_0Ԩ
_=��J��'�ў"~�ᨘ,Zff8sa�6XQ�xف�0�y�G���x��oW�V؀	���y�#�A�H��5�)^��=�C*�y2��$��2s�>G��%��N)�y�ۜl/
��͑="�d����y2�ML�~-$nď?`@��»�y��V�����E�XԊ�_�yr�&L�p���#B{e��Iɮ�y���R�T���a�$-&�x񕫋�yR�K�%g��P�F�&#|�tcR$#�y�&*�%��H�	�0������y�k�l�"�QW������g�ʬ�y�m[�n|��fϜ%��`Pp�#�y��uD�=�%�,p]��җT�y������i��G�e�Rd(��;�y��.�,ݠ��ȬU�h�(�c��y�ꊸ<�P�s�S�Iގ!�%D��yr�½�T̑dm��R�>,"FEF��yb�Ɩ?Xl(vϟ>R����D��+�yr�>jh�c aL4H�*������y����zt��OW<p �@C���y҃˔a���  ��U��=��)���y�kN"{L�����0FOp�q�T��y��t�������W�V0�"���7&t�0�B-(�YSV��<e�>م�\�^�[�
@	������u��
���?L�vYxbJ׮)�p(�ȓz| �����P_��Ύ,Vq�H�ȓ=�d�rt�D�-�@Ѩ��z��L��-�z-J�;	�@��T�=�@��p����O�y0�;A��o0�ȓ%���{!��h0��Nٍo|ńȓw�<�4k�n�
`S���
��!�ȓO92uz2��.�� ۥ�S1D����ȓ:A��A']�B���'-�/7CXE�ȓO�`]+`E�)P�epVe(j@��ȓ@�]��%Nq�En�?�݅ȓ'�D�r\�-��ع�~��ȓ7� ��c�-3�@u��J�8��نȓ+��aS1oR#��K�O 5/�}�ȓx-kG��g������2}�ָ��BW�� �>S{�	��_��m�ȓK�6�IF��ik� ��J��ȓ{������c$���:&���ȓw�58�Ε����S�&�`��=�ȓY#��qp��3^q�i#tN	�k����&?B��Aĉ2fS�#!�9x����ȓ5r����m˾�z0 ��̩yc�}�ȓo:�FJ�(v�Ts�S�[��l�ȓK?v8r�oO �X��hۨf�@�ȓ ��-[�^ Wz� �$l�����U����
��6&�	��O�.��܆������&ޛDu���q�E��݄�\D��%���T�x�dal��S�?  0��2"��!��5��P�q"O�8���4F� I��OG�E�V%bE"O��p��� 'c@�D�I,)��}�"O��� H%U,9��H�^)2{�"O��B�m�](����R`�
`"OB0�5�:��Z��ܗq_��s�"O���]$�� �+HL���"O�9k�$����Y'%,5Ä"O��1֯s�`=8@���s�i�'"O �JR��=V��hf�K�l�H��"O���cۜN�j��M�u��y0s"O�d�3.׉=�\ 9#*��w Lq�"O��iD,%���Ã*��c�R�"OQ��D-��"s�\t��͑P"O�HӦF��I����n$����"Oj���E$p�@+p���N�R�"O*��f��+��D ��_���ҥ"O�0�F9}}�
�L�o��MZ�"OD�8�˕2��B���ƙ�F"O���4l;��5)E�^�cxZ�'�b܋��:�z�""���#��a3
�'�ƭ���Æ`��� pw���'�rt��H��8���ѵ!Ðh�>��'i��x�-� c<0͠��,M�P%�	�'9����)5oB81��??X�i�'nH����&�N��aմ<����'�B�G�7>d.��+�$E�&���'ߚ!X#N7q�%d��8ߖ]��'CH ��&;���s�[+�EX�'�v ����N��R��8N*�}	�'�D�Ѯѱb��ՠ�AN;z����'�2�TC��`k�%Xe�@d��'�",z5�<,xb�I�$Hg0�p
�';@D�&�Z5 ��� f@O�k6>�A�'���Ӡ	Z�TXj�@��jzЀ�'o��P��8�	S�<���'�n����;n};5	��x<�|��'/`�0R&@�v'p@�s�p�B4K�'Αx��3�@�$&z ��r�Jr�<Pf+`b�Ii�@G�ܠ��Iq�<	vl	`tF��������`�Qn�<�N�?@*� H��ɍx�L�k��Qr�<�Y&>7D-�1���v���0�Tl�<�a�

|?�Y륨XG@l����c�<��O_*�,�B����XA���r��u�<奙������"�b51ȣ�u�<�fA�~D��C�l��ց�r�<y���Y�zh��eǳx���sR$y�<aÊ��or�\��$O;[D�@"6B�y�<Q��R�n0�m���6::)��t�<!D�ؑQ����T1t���)F��r�<�W-�=R��*E�� ���n�<y֫�,��q��0;��sM�k�<qŊ�J�D���nW�z����Eg�<�cB�/1��O��g���Y�<�f�I"f$�PqqO؏lB4����I�<	A�[ �y��&����1�D�B�<ᔧX5ri8M���W�39��o�s�<����]��ғ�hP��K1� G�<9pL�(0ވ܉b ɑz6][����<��
��e��1��foJ�J7Gy�<��<}�<$��JJ>J���Ģw�<W��X�q5 ��@-�}�<!��N�����;\���SI�Q�<� ���CA�W�d����t�@�8e"O�@[u	  ��[2G�q���	�"O�'X+�|� �H��at"O��A�߬3P2�d��e�"O�����K�,����ҵQ��-j�"O(}k0���C�B��l�� ݾ��"O���$���
HzE��`��l"OΔ:�ȟg���`����A�"O���]3y��3�,�+:7���"O�X��F�V������]}V]�"O
��f��^X ���	�`q>Eq"O��6O�G��I���98Z`�R"OX@t':l0�8ZQH�15G^,�"O�=i�K��NLP�GLP7�a"O��ِ�_�mz#���DB �"O��&��)�{��� Ήz�"O���Q�!��Q���O-���"O\L��텝b��TZw`��Dl �'"O*��-P��Dc*� ���""O�)be��h��xu�Q�N=��"O����*r��ka�^�.���� "Oz�x�C�(itB�*���	���AQ"O�\���	�@�ԁ���>o1�8b�"O�l�%�@+kT@�eª]�B�B�"O2]k ��V<Y���<���F"O6���?OuB���A��a�h�9�"O����d0�p��ah�;u"O@��dT�-�&Q�A��Efa;�"O�m(A�^�e�����L�*Er2"Oj@˓Gփ7�t���	6,�"O�AiBL z�(]��#����"O�ػ3m�<_h��/0kL�w��w�<��k[�/2�i�@��&Ơ�9��O�<��ܥv���3EN�js>����I�<Qg�!Wl8�*$i�|�����V]�<"�%�l!"�&�p�}2 ��<qr @'|��C*��J5��8aG�f�<�bn�sM� �� IӦ����G�<�V�\,m�
���Z�T	2���W^�<)�N3��P�G�<g�Fy�V�<$HP�3�Ā@.�f��d��I�<���"?��U{ ��~ĠHc��Y�<g�G�2�DbѽyM��L_�<A���=*�1c2���P��u��l�Z�<Y��R@
!���@[����m�<�E�Be_j���&�z�\�22�
m�<i���hS������n��@rP�s�<���ߙB�@=r�Ζ�\�4၁@m�<ٕ�,F�b%BJ&*�]3�N�<9�a*1$^�Q��D�j�z��r�<�3�Y�i>�1Y뛱3-l��sAKc�<��&W |�xȢ�I���Qz�Z�<�4��w��x��P�oD����\W�<)Q��	wV�m�6a�.��(2D��I�<1�%�f4.!���I�2[�:���I�<Q#�� �hW#��>z����@�<�J��GkMF�+L�d���iB�<Q���>Vv��ܩ� ����D�<�R���~:�)�5�'4������X�<u�Ύ$��`�!bZ�.}bppP��j�<��(�+K��ss�ٰr����EBf�<A`�((��(��$j9��#6�@b�<��Տ@?���-� �R�	[�<���S˞Q��'�:z,�ZE*TB�<� �#�L�	J-:��en�\�@q�"O��1�5k��,᠋��rw8ZV"O���
V�^�^��Ǭ������"O����[B�)��l԰X��|2�"O$���ː^���� _.0ԛ�"OΥX2�L$DE�m`�����M��"O�8C�ܹT���
oHƭ��"O��PFfˋJ�V��2��*@�� "Od"W'^(��,J!��F?��"O�I�*�-N�9�H�sf�u"O�=J3bҙ{葨�`�$e�y�"Of����8  iCĥ�g|2�i�"O����c�K�J�×�ǥ�$H�"O�L�D�5{����f��]w΅b"O�K��J�U&����'>'��(�"O
)�'M�5=�N�iRm�.yg"O�}A� >���F�ÖD��I
�"Ol49��O%Q�q*�#�/t��[w"O2�PB̔���<�p��iD���"On���#r�B g߅���C"Oڱ�4��hd�5�B3M``�"Ob|�e��&[Ǥ�Z4��)�֤!�"O�Y
q��*��LA��]!?괚�"O@���I��uB�'���d��"O*�ч	0���eL�;L�d��"O�DQ7@� sB�3 L�Rkz0�"O~����8�:@��%��&@p�C"O�UC�hǳC�(����
"E*\d�`"Oƹ��J)!�L���-�1LCNl�"Oh8
0H-D��lp+���"O��ȴ&�L[Ђ�*��\%2��!"O*�#��P�)��J��r*���"O �	tJ $39li�Fصc[�i!t"O��'�G�~�P4/B�aG���"O.�h����(�L�SGZ�Z8xy��"O���J�6b&�B2�2?�g"Or�)��N-���$D
~��"OBɚ�LإRl� q&Z����Bg"Or���n��J��gHȐy�*,��"O*1sƊڿ�$}��^ڄ�9�"Oޱa@�T�vP|�겈7Ѧ,�"O���CNY�3� 8ZpΥPŔ�kr"O 8��ǆf��Pu�,'�T�{�"OyZc�%(;��r�̨���"O�yZ0��%N�_�jy�S��y"�ް�~����߯Rߴ�[��E�y���[L�|�D��x7��˔���yR��g�q����j�M��y򋐪/^�Q�F��k�bP׋Ȼ�y�[
/0޵�C�R)c�e�&k�B�ɠL�D���f��T�&EI�W,o �B�I��p��G�giV�)���=K�fB�	(�iU�����'�ѵ�NB�#I�Pa��KB��yB�o�����'���I� �F!�ًc�ۘ8`H���'q���z\��ޱ-v�83����y"DE�"a�%�$�J%*@��� ���y��O��0x��ɰ*�D�B�H��y�g¤?��^�ظ�:R��1�y�l�^(n�q��<8� Xbaֹ�y�e���X�Q$Yu���Qf@�y�-юTlX��"�'{ˀ]A����yҥϥC�>��@U�yՌt�P,
�y2A�s����4�����H��ϲ�y
� Ș��ɘ!3����rc���"O�8��HA:bµ ��b�P@"O\@C&��#�P�[�!�2iW�ȡ"O���ԉ��mP,9`K�	Vl�{s"O�JЏw�4}�+�%:��C"Op��ՈR����$��yYv��1H!�D� �z�+��N�b��!���L!�DS
C0�9hӇ|R�����$4 !�=z���Qi_�Đ� z�!��^�J�%E15\8Yۀ.U�J�!�[#"�����d��
�,O2�!�d<Y�z(*�ɍ#hХ�	(D�!��/e`xa�4c_�&�.tY���T!��0T֐T��D�Z��4 &!�ĎB�|��F�[�H[Q!��L���Gݑ"&�q0���,�!�D�=����t�\�r�]a�mǷ^0!�$��z<����=t��L�<�!�D�Kf(���وs	.���J:!�$�>[ݾ�DC��
KH<��D�(6!��ƔkN���u���I|塤�S�Yv!�d�s)�l�W
� LƩ���җiR!�$^?	xH��.ĬG�(�p�_�}P!��4r_PH�70\P@5A)WO!����M9� �Evй"r��2H!��P�
vx��Z�b��"!!�ЁTN�C�W��t @B��]5!���7\��`��k�ʑ�6���K!�	�B!
r��hp!�^>|A!�d]�j�9�I_%(Q( 3�@��|8!�T�m�f��8�T�A��y*!�$E�-��Q�"�/ˮ=���g>!�d��C�N�2G��Nn�r���#j�!�$S���(J�� �G*�-xUA6 )!�$G*˒�	爗�/.]�c &!��XR6�S�ˇuP��4!/!��*��ԣ�m�T2�*P�N!�dH;��P������Y? �>��`|��!�)ڿ'�, �䧎#�~-'����I�h�*�Knõ\U
�(�mN�!�C䉝1/<�1S�:I�����B�	#D-�5��aڴ��Bᅊ�H 
B�I>#Uh�����R1�:�� 28B�ɗ,D��P��ʔ���iL ^��C�I�rA*��,��r�m�_�B䉰23�ٚE�� NҚ� ��G4B,C䉱(	�m1��#�VE�bD>vC�:��$1ԪP�<g��S�-P�4v.B�I7h������9=i�Y�%ˎ�k��B�IF���d�!C��P�2� 2gk�B�I�x��i�{��t"r�{��B�	*#~����:3'�����B�ɼ|�\D�O<;o
p��%��*t|B���j��o�V��� ��KC�I�N�Z�(�B8��FF�H��B�_�I:S�G�P�]�(Ldl�B�	AJ��#̃�KX��a�գ�tB�I�Q�@Mh��BY(�)��ʍ.o(B�I�k� KR ː��Qr��:aY�C�0n,JXJ�G�:�T�Æۄ`�zO���$��\�"����F>@�g�X�!�$H>z�hc�-�H����!�Dǿ0����R�` y���ӝ8�!�䈯SWL�c��U�+�V�C� �!�� �!�I���x�*��=Z+R��"O|�B�ɩzҞ�Hp-
gH����"O�%�qh��=�To�E(e�C"O��ȁ`B�&�8K�dO ���K�"O}!�+G� &2]sₔ#g��"O0 ڄHW�z��z��®?h�u"O<��U�@',�91��r*�0�"O���*,L�`�p��1Zn�Ĳ "O���Hݥ#�\��@�+XOb�S�"O�<�qI�gM�%h���'�<y#�"O`�0�H��p�ro��N9���"O,u���������*�8��"OjȆ�1l��#F���p$�s"O�����_"KD^P�B�F/n&914"O�ag�I��8Y��I�8 sq"O�HU�K3xr��UN_�=���"O0TѶ�]�~�`��G�H�Wr�U��"O��s2e�{/�1�[X��1b"O ,X����r1�Q��.T߀5z"O�H:�� ��pxCԹ2��p�e"OZ�����mvɺ@��!/^qS�"O�tӥ%»�f�YCn��HIس"Ov���O��"��Բ#�K��ѐ'"O�h��ΐ"DF���B�'�jh�"O~!�D��74Q����4!���"OԌ3f�Q�x�v�3%�۶"w�q�%"O�%��4@<�� UOZ�L��E�0"OU{D`��	x$��NK?��� �"Ob�0 �Z�P�@��G,ж�9g"O���h�*7X0=�� 5�ؘ�"OP]�5L[&nB��LO��J� "On�;d�e6�ӡ�ܫi���"O�M#C鉓+R���� Q-J|�(�p2O*���h�'����5뜜4n��� �̍����@ 4�f��Y>�8��'�>��2
؁2fZ�%�m�r�ȓ0r��OM�5 ��rP��U��F��=
�dL���o팔`�(��ȓG�l}3&�';� �4o*��y��@�Ȝ�M����YPsa	�)��ȇ�Xz�n �`��p�E��5F��
���A���Mr��X�$E�lP��ȓH�}�B�%���ڱdڞ1�!��EG�?Ųͺu�UWg����&D����)�0A$�(�L��� D��&��*L6�@��խBs�Y��?D�r6n�9~��0�aNԅ%�D���:D�������~�{rE^1O�]�%:D����D�G5��ۢ	_�Ab1�3n6D� ��MސJ��=2�Oۧ
�8���"6D�8;�M�<����6��_��5�%.D������y�L��*�/�q���/D�4P��͓>�^m�T��l��%3D�h�˗�Pl��ئY�����K2D��B�T~���Td�=q�\m3��-D���4HD<f4����WP�H�n0D��±�V�7oAi�*�i�@�ɰ�3D�<�4H�;O5��ؽ<��[b3� �5H#!0� �g��f$^P�i����ӂD�o�^z�A
�c�v ��SE�(B��j�I���$:�Xхȓ{H�q����('��T�F��,�ʹ�ȓ�iZ3�˕��+P�Q�o"hq��	0xA+��ǎ\|"'b/Q�q��w���HG�	��B(J�LC�R�܇�S�? xqㆂ�2�j5�)K�QSt"O:Q3�jS$~n�p6�A����S6"O:8��!�	U,,�цыb�T�p"OF�Ӌ4e9*��a�	9ti��9�"O!�&�=pL8��c��)xF��u"O��
��9��ȩ$g�:ܔI��"O�,�K^�1�D;��ɚ*���A"O�h���B�_#�!;�쐏[�� �S"O�H���<1&���̰Hüd�g"Oδj�a�Q��q2�j֔{��x�"Otb��U�M<�x�#�D?��lsE"O"Q9&Ț�otd8ŕK��U{D"O~�K7��;j@5�QEW	-�N�A�"Or|��@��=���B$J{�,2�"O�}!��O�D\���
1IH9� "O�T`�C\�TZ�:pʌ:q%�akb"O�<�B�+F@��3�Ƙ5uH�"O�!�e�D3(�����"O��cS��;��ZND���"O��r��_�h���%>N-��"O�(
&A�w�\�gF�>7�T�U"O�QK�"�l��a�W-J��"O�P��ݫTh�$ȅ�O�	y �"ORЂ��0
&54�8`��t"Oȅ�0D�h2@�	<��"O���D�[�I9���獔<o*�L{�"O T��K��/+
�i��>,��y�"OeƎ	�Rmz�O;Z���
�"Ov�S�e6f,�)�/@>�X�"O�<;c���m<�ِ�����1��"ON�"#��zK<H�nӟ'�N���"O�騃�U�v�D4�m���:�"Oh-Ah�0u%ZdS&��#�����"O����k�-"3� G�n)��"O�pC�I]yv�	����2i�4��"ODl 3D̷8ġV-�te�"O��2)�)2���e�@/1f|��g"O��0C���{،�"�B�F[� YT"O6�� �Y�P��̒��A�N[���"O�L��L]�#Z����
nIP"O�݉cK�o�zq!4gU�����#"O0�A$�Y,Z;P=�w�[�X���D"O��ʃ�^%5��}��Ըo�n0*�5O�=E�4���a��ze�0k���BQhǆ�y��?�N9ᵮ�?�Jə`�.��D=�O����k\�^�<G�û^-�]@��'��I9�Q�u�|�[	4�FIVB�	�j�D�h��5gM�]0a� xm�#>	��)��W�|TCp�L%�Vl�s��X�!�$�?.��ˆ�r���ơ=@��2�S�O�Rٓ���c�+�R
7Xܡ�@E(D��q��pS\�ƆT*��2n'D����Xg���(`m��B�`���(D�yg��3�$X�ᇑ.����&/&D�����B�PE�P�
H]�)���$D����,�4|����F5eB�@�f�#D��`b�\tb8i�d����ș�	#D��Y�/I��2���!!�d D�����`%ԅu�P ���r҈ D����'�L��!yrO̭C�z��!D�����Z%<C���K�j�Ђ�!D��ؒ�܌}޼p��I�x�hd�*D�����b�*X�VOK��W�)D�@	���:_�&A��He���	'D�� �=��J��^fp"��J�JXʴ�"O�hBǜ"�b�xlT�U@�Ċ�"Orȇ��XS
���0$�Q{�"OD͒��G/@JE����T��Qc"OP�Ӆ�ӊ8���Ѣ	��[\���"OVQ�V쇋\:X��	ȁ{C =(�"O^/l��&�99��P�bē-�!���2
���'O�cS!h���
�!�ьv�j� �?��8��o!��c��8 v W�����")�!�d46�z��5�7\F�!g(N�f�!�$G� ���Y���A��b��*�v\��򤉚�8,�~&�Lz䬇�t�LJ"�{��z�f)�Hr��\o��h��(�2H��fH���		'�X��b� `��CS�z�0��$����m���'��	��� J�9p4��ᛎ����Ya(�"�ˁ��'m��(B䉣0�tst���A����p٣vL.�[N�2�WY��K2AQ�X�1���i5#=�y�r��6	����M@<,!�[�+mVh
�Eͽ��$���CT�����ŧr^����/M�C�Z�$�~���?��^���wE�u��1�j��l��$Z?`5v ؂��	8œ��0��Ł��&]d���#�=J��)�͜9O�����	2��P�(�q�>��f�ߜ6�ў��S�L"5�!r�\6L*��WgM�=#����RKǖ�J1�̷:[��"D�O0!����H̙!��ӯ���87o��Ҁ\`{6��7�ˉw��Aa�K
ƉƇ�o�'�D�q�&*��q7�p�����'���R��q&�86�֊3����ϛ2/�zy9w��`7`����
.��)K� P�!�%}�OL>%r��揕�P�z�ЈW���O�D�1�>��.X����'$�->�L�BS�3ZdSU֜cL��s��.1O8ܙAc�W�f�1Ǔ`�,�{��[%��X��.�L0Xq�'� e��e�d?i�I��I�P}�Ɖ¬(�6��@RR��Q�WU#Z%qE�
�Ur� C@��)[�v�Y�'Y襪�!;��Dk���x� �޴U8tK����m`�e�?�M��Ço�p��M�<w]������AT)*��8�e	��s"�[؟�Y�gB*Q�~�� L�
բ5(�m�l�ah�OF�˰D�`MZ3�0 �F� ��	Åh����A }�מzpʡA�Ǝ�3\�4K�����O����N̛�~�L��E����%��d^&��G�!
�ܱ6R�8d@�*6�ã{�dhK2@�h�*�c�'B��9!l�7����L��4$j���O���ׇ��~���yu@[U��?;f�2�̋*<�WG���"��C?w�z�a�S���q 
O����	�+�R�آO׶2B�0{ҷi�r1���R�ɚ���aB����M֓_Qĵ�_�of���c2i�(���I�Ϻ?J����}�<	� �!m���*�i��GE�\���1PkQ�3�* �r�^6s@h�ŭ�~���� ���K���M\'wj(�(�0S{��K<�O��[W��:�����ϡK�J�4$ò����g��L��,�D(�#KI  ��{e���f�'o��H����\��b���D�����6�r<�H+�p��,
a��\@�.G2���*��5	*69i%�Q���H8�(��L��ɍ)�4-���8Ę�[���g�6m&d���)7��z�P0R,U[ujF��p&��SS�1. �P�g�!���D���H��ȓa't���b� /���Hc)N��8�S�bF�"
в�6�����;��$  �~��d�O�.P�,Z�I�Ŗ|J��
�oXS��}�/�Q���!�m
��s�^�)!�h��	1�<�& *=�	�r���oҞ�'�ўH��JޚX�����K'��۰�*�+������V:k�n��w
�g�:4�b��+x����	�g�p9�E�hhJ8��>��,uX	�@!���o�C�@BQ4O0X��e�?Q�ZI
�m�%C��Ie�ÅZ�?i)�T$6�J �'I��)঑��2D�z#��2�M�#X�5!����L�4�F�qaC ;�9zS���OBr�<��f�h~&�zamů<Ju�R�[؟�cs)
^yB���K�	Q��q�59�^t�ѧD�9�΍0��M�j]��	��ȉp��U�J�sd�e �?)���c\]!O��<c���f�%)�(��E������9u���5D�����ǹY���æ^4u���%?��ͽi9�(���ۋ9Z�0���ơk���5�KObE�c�ݙ2�!��.�v����O��i%JX�#�5��LG��ըa���~&��T @	Qz(�+ڊl"I���;D� �b���9�H�r��ԭU��Jt��>YTjד�p>���ԧM�&�$
V�c�$�)Vf�o�<� ����hQ6p㕧�!nd�=��"OJ��J%M�rmc�	����P"O��`�F�\ڭ0��=�t�Z "O�pk���uw�YSăQ)E�su"O&KwI �iQ��H@@ݹk�Ρ��"O2=�w��i�*��\8F���!�"O.��R�#>BЂ��s�mq�"O��I���C
�Ѹ�R�ެ4"O��e,ơs `�CcR�>�:�!�"O��@A��*`��BN��q/4��"O�@�!C��J`��Is���m`eY�"O�0<c&� w�7�B���"O6���W�*]~�qWC�1a��v"OP�s�J Cr@���L�L�5"O� �4�x�&�C����}�@"O��D&��l���S��KT���"O�iE�.��EA0�� $��Q%"O\���,,!޼����l4�p��"O6Q���*Sd�8�MP#V*�("O����-U�T�Z��"���(h�s"O��E	�+b����N)�^E	�"Oy��nзXP�I��l�	Bf"O�E�BB3g�D�34��W���{r"O���b���+�r @����]���)"O�P1Ӏu&0�{t�,�:U��"O%�5L�4m��8b"��Tl� �"O8���M8,,j�BR�->���;�"Ox�"��&9��I��HG/�P�
�"O��"�+��`\�u�����n�x�	�"O���D�.#S�5��P7rY���"Ol����o��e��&{��W��7�yBMJ��L��2.� ql5����>�y��	��`C��Vp/��3w`���y���$3�6�+��)*N����N��Ra|2�ɈkV�4���V�֩��M���(Om�!�)��-����(�R]��	��lQa��	&s!��A�<s�<(A`'{��Pi�q!���:z�v��f
ՋS���cA�Z�D�!�$�l�\$Sp AT_d*��!�d	�:T��O�C�ĩ�'���!�d�9H�~t�����;�\@���?}!��(pZ8UY��S�f�G��hr!�Pi�����2���K�Q�(�!��X*Bq�D�((�ջ�`W#R�!�!je*�c�I�wg\����!�D�o5v����w��`R�τ�!�W�K�fP0!�	^�s�AO�o!��\�T��h��s��h*6oA�!� &u,�
@.���V N2s�!�DG~a���S�i^�xR&�a�!�d�.n��$�5*�g��#�L4)�!�d+]O����j�;�*���d�<�1��4g�ƹ�K�6�jH�Mg�<�f�S�N��$�3�PXot���bAi�<wD՜�H�T�]vؙ����Q�<ɱ�=I��A�MVA��	\Q�<�ɔQ��
�$cJ��c��M�<���H�K{F��	U,[�r��'�Tv�<q�ឝ?���s��e%��աOr�<9��[-N°@���՞j�>���"U�<y���b�p<S�-�2,�xC��WL�<1���4�T��+�a�؀ 	�`�<��@¾~�( �C�ؚ9p�Q�f�<-��t���0190I���Iގp��S�? ҈*�	B�C}���FDɪR�$�d"O��b�S( ���V��M�t"O�x1G��!]���0�JV�a��"O0A+Ú A��fˎ�R~|<�"OLٳ!Z�Ea�ыΣ0C@���"O��(7eK���A�TB�3|(���"O�=��'ob1��j�B�"O���ω*V�:��&��D[�M�"O���r*��w]N�a��L�b28��5"O��T�D�z��|+�B h��"O�Q�q�C��(�Sឬ6��X"O`���B�<#��A/C1p�ݳS"O�����Q(V� �$��@nV,zf"O�s0�A�0�V��4h��,�l��C"O�}`��B�]��03��B�z�UH�"O��򨞰�\5 ���4����E"O��Qr^t� 2�"�8�h�0"O���F�N'
�r4�I?Q�&XH�"O֝[�X���7L	�zr�%qD"O|I#Ҋԯ`d��n�&Td���"O��x�E�++��#��)J�0+�"O��Ve#.+d�K�K'.h��"OyJ2�6f�N��������<��"Op��q����U!A$�]����"OH���fڲR,�Z��@���Q�"O�̙��C~���ȓ�Ft�`lb�"O�L�%+Q��DA5!�	]��x�r"O���Qm�g2���¨rl܉Ӳ"O�m�Щ�L�f�Rs �p��ԃ�"O�a���m�L�1�`,:v �"O�	�G���7���/�se61Ã"O^l�Wk�V��q�hOzr��"Oޕ+�+A8r�� h�m�#Mx��h�"O�}x�k2b'8��T�͉fR���"O���@DR�9���S��XU�ˆ"Oj5s$M�%�(�i�(MX����"O��W �;��S��g��#"Ol8��X#y�K�dOr�A�"Or$�G$F�q]\��T�ܡ0R����"O>5��z�w�M$ESx�Sq"O
��j�+Z�(�č5~_���"Obh��D�B�څ)I�8u9�X��"Olt 3��B:�K�"ي;?Z�ن"Ol�{��O�5RvP36��-B�&�(�"O�X	�E�V�.7��ӞC"Of�p�L���D���%�L၀"O��
���?A6e�c�N�� ��"O�����.-D0�17G[�@�0Pt"O̜�R��9��$8���QRt��"O�ݢvD�83��e��Ԁ1G���"O씑w+!��E0��}J�1�$"O$��FlQ�w�N4���>N�Dx"O�Ai�Hْ{�|��WD�D�(�"Od4c@�8W<L�d�,^�2Ā"O�$!�j�88^4Bҡ�	r6�e"O�=� H�ҌHDn[�a@��"O�Di���v3<������)	u"OZx����48Fhк�l�M����"OH`��G/@|�̋�DF�	L���"O��#�iԷu�4Q�iRL)+A"O��E��F���%�A6��	�"OJ�3q'U�������!C.2�pp"O�����ݫ	Cv�b6���* du��"O�q�!G��1��a��M΃Z��!"O� V� �-6v�L����~�-�"O����
ͱ��Y����00�"O�9��M�[� =3�����Lp�"O�0ERb�<j���%Y���B�"O�����Ό��-V�J�F�)�"O���SMΙGD�� ��>�-�T"O�$����(Y�q`���D��yR�ȸw&�a���vjd-3����y҅GH���	6K���A�F��y�*P�tjJI�O�	AF�cì�y��5��9H��B�'� �d&�y�'^ p�4p.R(n2	�Ї��y,��Uj����bH0L�B�h�_&�y��C���
AK}�MՊ���y��M�>h���4F��{���bUi��y�J�/#���B�$}���T�U��y"ċ�'p0!�"�ô�uH��y"m�d��T�gQ}�֥2����y�G% ʚ���A�X��JVI��y�A�m��h��f�]�l��ҊԳ�y"�N���0[���6e��qw��y��ww.�����P�F��F/W��y�#ڊf9��Z���a��y��ƞf8��쇾$$���alK��y��>!��o�/&������.�yM	0A�>�
.�C=�)��GÍ�yBm��>"�YB��FEY� ���y"�z�d (7�.W`ʩ����yB,��]��mYG�NDh!刎��yr�O7)*ƍH�^�9�v�{EIȆ�y� �3;M~Y��
��P� ���yR���cy��d�."��ª��y���>X�:�ӣ�F�;h�����y2ڞ9�=�q�� ���I4��!�yR�	�Py�	��pnҨ��΁
�yb��5h�����;w�d=%c���yB�Ֆ?_���5�G2�)�h���yR��&�Ra;t�0e2m��H^��y"��1?(�P��1�$�6*���y���45�MiR 8,n�z�@�y�N+��!zwmZ�U�X`˨�y��ќ<81XG�@���\P�l���y�C�u�1yMS*F�<�X��<�y"k�i�)1��G��8r���ybʄ�0X�l�Vi�6�`Ex��A�y⪑��*�;!&Ǡ-	�4�1F���y"CΗ�<�B���^��[!�ѫ�y2�7��J��UV���(�a���yrǍ��V��G��C�T��iO�y�卼o�n��E	��G�b�F��yJ�9lм��$6�� ��DA�ylآm4�a��"A*��B��y��O�)�GY�.�E�P��y"��TI��b��X!/k���$+��yRh4�윐�&�?� �#�yl����Zb�̘%�PDIq��.�y�h��1�P�90�ǔ�n�0mJ��y�N��O�9!a.�� <b0�0Ϟ��yB�X�pQ.YJ�+�
yc� ��-��y�k����{�.
�>Q2�����y^��q���V�M����ڎ�y �C������u�J�*����y��'��8�DA��F��)ɉ�yb�I�r]�HN9q@R8`���y
� `e��+k �;�k��  x W"OV-�T,�����J�"7�Eq$"OT�[������	@1	N�o
�xC"OPQ+D��"���s�Z#�$ �"OP�J��֠�UƊ�nĦ`�"Oj����X�,M)BnU� <�@"O4���;%�09A���:�0Ĉ�"O�TR�C\�x8�̰1�s0rMs�"O�p��N�*����L�<T��&"OT��BT8i��5����4���"O�`5M�p�(|�uÛ�x���4"OHH���
-����@�*U���c"O6HZgΜ�x����(���vtz"O��N
�_����,C�kpzHG"O"UC�`�KaF��@	]mY�e"O�U8aj�?��av�ܿnX��ʰ"O��V)��Uð�Q��s؄}"�"O�l ���8P?���#�<��u"O4y#h��(���3%�m�EY�"O0 ���,��k!dJ�F�<�"Oh٣vgޗ 4z�:�#�2NY�2�"O�}HpL��a1VU���b18�k�"O�"b�= ���{��	=pd	�"O$	��Z��0ZE��?�@\@�"O2�k�k�6k�I�FS�TC"O��AD++��!hv'����"O`��g&S;Vҝ*���.FzFx�#"O��ʓ�!y�̭i���f�H�s"O,Q�0C��;a4m�Oؔ9�)"�"O��4僴F#v!I��R�Hw�4�V"OtUj�t����1M�!jj���"O����DP���T�� X[��YG"O<�Z���9���:T�ӭZC&xP�"O���Ĝ�'��jw�
�(F��X6"O1�OY�D�H����[�9{�"O0m�Ǹ
v��P�68��"O>� ��/1xP����G"OJ�kpȍ�9���g�c�0�A@"O�p��ȻdG4y��C[;(�z�{d"Oƕ����!3��@�#� �,@��"O���`GZZ$�q�W��"��b"Oj��6.��f�XD2Sa�}�p�i�"O�\z�KB�K)r��)�$>`��"OU`�,Z Pz�L"7��Qq�"O��a��Q�E��m�������"O�y�7L
��~��S�֓3!HyA5"O��+Gh�5���*B&�H",�i�"OJUG�����咋7 ����"O|`Q'ʆ�������*9���"Op�b���
JT^��p��Ќ -T!��nŎ����L����MH�;1!�d[6t,����+"O�͑�l�!��<��%��O+�vi� `�T!��u�>!� �=`��B� 4Q!���;vX�%�B�s�B5�.C(�Py�\Op��)�R��q��%�y�MA�i�O��O�]���A��y���:��U��Η:a�L��Ñ��y�ɂ���qgj��<��2�A�+�y��9g��K�R�Z^��%L�yr��j�0��tO�*.k�[f���y� !;�����r<��+�/�yR㐰c��G� M�l���^��y2�H���8hЊ���	S���y
� ��P������pF#ۯ(���y6"O��&�bd����#��c��	�\�z�8P�M/9*@4 A�x��I�]l*)WÆ0@0�3�&�.jC�I�2�dCq딳W�%���1CR�!C�l�<s(M2;d5�t�S��Q!bV
P&�\j�Ԁ��O�B�R�0�.�ZÇF$�0|�f	њ��y$�\@O�,�pC;l��!�,G�q	�Č2�y��)�|Z"�AQ�Q	��l����L<��÷R���hQ��Ɵ���3�*���O@�A�q�@rb�!�Ch�J���'v
�(� �ۦe�I}���Pb��A�O�)�TZ`�͍2�R�e�����[��㥃�Y�Z�����~��^���O�>�R�U}�u{��Ҕs�	x"�\�E>*}X���i�C>&e:�T
 �&XR���!����?�!D?��pQ "��&�0H٤+�!���z����U]d���[?�TD�J�Ę��m�(|���Y{�$��Q� ��3�3v����D	՘��>�㈹G�b���-RVp��A<��sD�A�O?)9F�+V�1�u- <.L�({3�ceB|����������L�~^<��C�s�Z��?Is.2�x��g��8sx |��dӻL�,�a��&g	���.�[���&ǜ GX�5����d#r4�`s�7-�>&���PL~"~���۩A^J!j�E���p�a��;}~�7��D̶�D[�9��]j���Ա_XI{チ�fC�	�7-�3��4�?a&d�Пx����1�ȟ�=sc�@�Zk��u/�M]�%�ī��Р��[��M�������~ڜO��iG.�]�t�߄@�Zu��J�?>�vP(��5�y�u��o�N�OI�Q�ɘ��L|h�4=�,y{�$
Q?a�'������9�������L,�`rM!�h}I>ib%�!�jy �)Y
��O�U��.�&5��C8h=6D)�"O0Q����7Y��D��y R�8d"OT����)y��fiu{�uHf"OX�Bs�A�:��6��A X*u)5D�h@�JO^��kϱ %�Hp3D�XAD�"l<J�K��չe@1D��Q��\Ǥ����ť>Ҁ)�q�3D���w
�ghk�(о2�ИR�1D�8�0,.4�� ��}\Թj3".D� �s@I���$(��x0���C7D�P rNU�vXѩǥJ*gx��cD7D�4&�$�(�#�G�O*�r��/D����ƀp]
��'�>q6�|Q�O-D�(��V�y̬-£�I��P�J-D�����b+<�2�E �CF�T�`�7D����X�F�P�ْ�E���W�3D����.�g�ax5)�>n�\qr-/D��˥i����u-��NX�	+D�XJ�D�Q3�����
!�X�),D�$AQi�����kցQ{�=y�
+D�|�"'�.�DI[���B6���7N*D�,�umP5��5a'�ΖFN���	&D� �v�ūFi6D���K�a�԰���"D��`	�B�X�j�F����U�*D��QǗ�v�0���G ��Us�L)D�� �N������-A�U�b�%D����Yun6r�D�DJ���3%%D�h�A��*�=�υ�n`P��3C$D�3��ے�aa��_��a	#D�dC�!�;���K��HF����	?D��16G�+hj6�`�΄=m�U��';D����	H�w���УՙqUZY�vl9D�����A�NH�3����7D�HiV��`�(�xs�U"<�LYs�k6D���P
�&�l�(��H�4
! �5D�����!��e�FG�:;g�Y� 5D�����>]��"�`�$�@�1D� ���bt�i�,�2xf蕊��<D�(�7���Zx�:�F)	��e�e�:D�� �x�#�÷8�I�Cl����E"O����Ɏ�o��
"���I�J�i�"O��um.)u0�ʢK�8����'�HՀ�KĚ(��5�O�y�jU��'�8$����%P(u{a���m}@���'W�E��Q"S%��	�k�?c��2�'$�����6(��$B��W�<�8�'Nb1�cF�7Y�.�X�N�"��ɚ
�'6,���/�r��Ý1|"f5 
�'�萹��ێwV�i�bmQxµk	�'���	gn����S���O�Ҁr�'�X�Z��-����EX �a2�'�P�.�,�H�2�O����U��'"� ��y�<��b�M*6�ͻ�'@x��֋F�9���:BfV?N`� �'.���"�^@�:�i89�lQ��'�$:�ܦk���d81U¬8�'�hHbD�:qU ��U��'=\ �'��i���
��>�`Y9L�"}�
�'AD��rƓ7	�u��hL#J�8�`�'�س�ꘟVA�؆��<Ts��k�'2���ޯi���i��˾\�����'��9qVl"�n������Qi� �'��aB��.ʺ���=?� ��'U���VGE�{�Z	���?
��
�'zlq�@ńjO�+C&9^ �q�'�ibd(�ru�U.H�~�R��'��D9�����5�p9J�I�'�n̑��؀^-���ˀk�̫�'"d�K	�N��.�/zB�Y�'�qkT
=j�B�.W4^�S	�'��0!��g�j݋b�
$M6@�	�',�Z4�&6�Q�LIz�(	�'=�uQ`k�q��0W�nm�`��H�<"����eo�It�4y���n�<i�OM� ��V�^[L��s��m�<i���~y���$k�W�HP�<A��[%x�!��J�	{*�[���H�<���<v�P� o�Y�!UC�<!�e'mx8P�+P�O����I�<�"0
�p�	K�UN0Z'�o�<Q���	�$A���<H�Rp����f�<�7�ͶO[H�B�m��
a�T)RC�z�<у�@)$lb%��`ԕ3H`h&��y�<�q-^-Gp�#�*�Gt�� A#�s�<��L0N�ģ�DҏH �X `Zq�<Q�'ͮ9Ք�;T��Gn ����W�<Y&L�������:�Jp����P�<� J5j�t�uCS>E�IXbO�w�<���^)1O�$b�0iBt�_M�<�� #/�5���U�*�^e��"�H�<��d�6�6Ѻ$��u��A�1z�*B�i� ��*{,SD�"E��ђ�'e�1��
&4ȲQ��,<H�My�'����S�S���;��Q}��J�'A���b�;
�&�w���DՈU��'�X��ǀP-#�\���/o�1��'D�f̅�u&\�0W��Sf����'=���$[�n�>��c!,}j4�
�'_Tła ��FC�q�ǅ� �qJ
�'m�@J��ٙ:����E��!�';��
�MC�j�R1.�<�^���'DN�(��K%Z����? 8 ��'S��a��%Z�Fm ���}yx�1��� ��@w�\�AQ.Y�R㟔Y��B�"OB؂��ߛa���$�\�Z��m��"O�c c0@���/��m����"O>ځ�Q(���tm�7
,L��"O�13qI� ӸJ�M�&bm���'�'j ��vGI�O�L�p!�7//1)�'������KN�(�rN��&V����'��Y�#�M#-`r�;��szl��'3 �tB�C_A��?Mɲ��'r`���C=T��!�ľ=���'r4=�A*�=O44Q1�"Ō'�Б�'�HhR(�,67@��nW�R���	�'���)�GO*R{���F��@U�\@	�'�8��Ѥ�3t8�,y�ҧi�����'����C=8ީ��ś�,�|,��'�p�rB@ǘP���*I�#߮y�'5T��N��̩���(,j��'��#U��>0` Ń�(���'\�5)W�\-O;����Z?Q0d�'�V�S�V�Fpˆb�v�L��'�����Ӛ��1�V��	r��e��'���WǗ�c_��E�(�ڳ"OZ���+d���u�K�%�T٘�"O&-{���5�	QG��jw���6"O�rqf\2~����r@�'@t|(;�"Ob�j���]"�,ƅw�ڵp"OP���:�&PJE���}�!�"O�t�d���x��c� /<悬��"Ot]0g�
k����U���2H��"O(	��Fw�����Ǟ5!�"Of̹��ŬeBY �G�bf���"O:�Bd�ļ"�
��2�߃W�*�Sq"Ov��U�3*6��P=op��"O,i���ndd@���Z7���G"O�j�8(�TC�@X6���"O��kD�L��(k& O�q$��SA"O�Ńv��C�xe[�o��4���a"O��0�֕~²ȡ�n��l����"O�([ aI�rG�q���ĹE9�H`6"O��7�����#���L,�)qV"O*MX �9gB�\�s��5���"OZ8Jvh9s"�Z�GS!K��:u"O��@Te��jm�-R�vD�"O������`YIP�V����"O*!kR�6Ƙ�����>~�r��"O�i�D.E�_���Š+c�Ja�C"O�(h�ƌ#z�%R�u���"O��*�'@�F)�GeM;Bn���"O�M`���/����%��#d(ӵ"O����*�9i���e�T���Y�"O�*��ИX�l��AD�J����'"O���iѱV�V��!;@���"O���Q�׹�8�z��M�b$��"�"Op�i%hX f�2�ڶ�Hȫ""O&��!k��C�޹�bφ]*��E"OD����P5/��ΥN����*O s�+Ϫ�\@9K��l8"�'��T�W&�S"0hB����Tp��'�~���u.V�Z��)��z�'����vL��*��&��A�' ��Y�����D�Dh�!.� r�'�&!r��t*6 �s��Ey�����aQ�%}�9��o,��5�W�<���75�N�p$fЇ/���V�J�<� ���V��~�b b�O̊-2)�"O��Ü�{M���H�1"l�"O�Ib�'�Q�M��߽0���G"OT0:$҄.�yIՊ��-���(q"O��!�W6c�!�T	O;AZ.,X�"Ox�i�o�
B� ���
ESN"3"OL��E(��yS�������ZD�Ho�<�C�-t���X�!�2b"T�g�<9�*�4rY�����R�p��jd�<W޽d���w\�)i"�Hf��^�<�ì��ڡb�jH�h2$l���r�<P�"��1�<v6�)�L��)!�$��B*~1�U���Xh���N�%!�D��ld��Kw��<����+�M�!�G�T'���s@��|AT�y�'T�M�!��S4k�Ia��N�9R3�H�1�!�dɞE]�%��!�0j8�UD��!�d����q���?P$�X��)l!���D��-P*h$BT����!�D̥B�����v��b�̄!��G���m-0t�d!ET!�Ě
�N�F#ĺ�4@��
� ~%!�d�	[�j�I`�G�����ʒC!�dT�{����󄓸��h���w!�D� 'P�C�ɛy����H�k�!�D��g(�xh�f��*���j)U9O�!��!��Lx0�S
Ih(�sA�9$!�Ĝ,q��p����	�n�A��̥8!!�Di�hPd!�;r���x`�U�:!�*e=~k���&\�7d\�mo!�$"2� c�$�>a؅ÒĢ]�!��	>� �  �   >   Ĵ���	��Z��w�D�8,���C���NNT�D��e�2Tx��ƕ	#��4"�V���d�9�o�0N�(���P�zԾ�a��e�ր[Q$K�\ ��W��M;C����!�M�����C��8�	�c.���	}$f�І'�fQ�1�4�����1�Q�|����l�zJ�0�g��1Z�6�Z��" vp	vFEGи����(t�	�K�:�R���� �py27�мj:,�'�L婀/��`�"UIT��7'r��̤��,��'$�牰c����W�t��O�r'�C�m_� �rN��Q��$�#�1{(�	�ƕ>ѱG
#s��8��>9��?|��h�'A@IQ޽o�B���Z"l�.���'�J�C-�P��'9t�åb{����S�<�&&M#33��1%N�&d�4�G���&�[���^��" Q��7Gw�S�e����H�  ��,I���{�.�j��ޚ%���0\��@tg_�T;f,���<���]�Ω�q�|�83E.T�a}��z�JW�j@�J��O�U�'��<^��'��F�E8��[G����2��LH�^�\�`!� @��	-Q`��@�,bf2OjK��$�B�;��c�N<��M��uy�\b�ḥ|�pd��"p�Z��fl01�Dn�<���'ppgR���I
~�8D�DÇ�Q�N,��Z�%I
r�X���%�<�&�'}j-���@���	Y�����ڐ	�����B�Br��C �"��O��P`S"��$H�<ɧ!�?+�X�I�|�T�1w��)����Ǭ�&�t�4��5sU,y�ɨ9I�0��-%��[�RFh9G�߯n��R��	�` �b����fb�
�c�V�I
p����c��#.8�(ȉ�:0�Ԙ��� z�H4"�M�&����mM@� �"w�G2'(�l낹��|;�m�E���#�`(��x�e�.^��s!CT&:q$Q�'�*|�t�ݘ'�܉�Ul�L�Iiq��X���
�w��@h�C�҇M$��O���ѓd91Oh�����#[Qn� �ŨX���� ?fRC�ɚ�� �  ��r�WK"A�|Ir� t�B��'�� ["k��'NB���skZE`�`P{?y�wFB�k&	��P�1�
�~���Z
Ó`A�<3��s}�A��"�I�#-�i2�H�y%X��ă�� ��A�$�f➐ ��OH�oZ)��װ8�14�Q�*���VOڬ"�b�'?b�|2�'�'�B<���h�L<��yT   �  �  #  �-  Z8  �C  �L  �R  >Y  �_  -g  1o  �u  �{  �  Z�  ��  ��  �  ܠ   `� u�	����Zv)C�'ll\�0BKz+��D�����b�f޵�y2�S��y"��g+:d)�i��B8r�Nϼ+d�]26�R"�Tm�ƎZd�
���FL�Y��̭Z^R��.	Ќ��ؙ5��˗H�s4ڑ�&)��_������:b���9�/�O�A�(ͅD/��#"�%��'a�ֆO.tz0�+ѐgZ\��u��&�I2��� �$
0"�(ѪG�%[��m�;^0J��	�P��ן\��m��ḧl��W�h!zS���TP&���>5X�Y�4X��E���?9�'J����'�?���~�hwʕ�Cج]�&�,(Op����?���?����?a�4'R��;v�� �e���?qB�	�:2�x(D�ă���"ߧt���I��򄗈z��u���!�v�N�Гm�899JͳG�Y<[��qU]�����'8J�w��h��*;OX�Y 0LBH�r`܀Uu PQ��',�7�O����O���"�d�|*�w�r!�GJB����r#�%(��Ɂ�>�6oq�8|m��M+��9웶��1{��6)?~ t��,�^;�I�G�_�����ۀG`慖'țhpӴ�D�^:�M�W'E1_��yt	� Ga�wݙ(�M�H-���#�
[Z��;��	:Ӥ	�H6��8sE�� �4UE�6�O>T�Ә%L��&P�"y8�r�X��V�!��Je�7-�-Z�C c�*z�&QI����Mk��ʹc�zVa�Tm�9�M���
m�e�& �6)q<H�QL��(?.`ņ� &XS�i��7-EϦ�jӀZ*�	�sB!b3���b �jJT����s�Jeq�!�^*910�D�(G�T��M��i66-�R���ꌛy���Qɟ%ʨ@�/�&G��4�[c �ى�l�ʦ����FoB ����;���Rq�^ڟ��?�$���4m�"��/2�� ��[�II�lʇˍ5�?���?����zPgS2�yK�?A�o�Ѻ��2GX��$�aa�U��?9�^�X�����?!��^,떉�*���Iἓ ��	M�^����wRŉlb�$�ddZ K٨����C4W�P�Q#�@�h?�����o�������v���m�S�8�he��G~�Ld� �'�D1*#e�-�`�`秘0C�� "���?�����?	���?i����T�KW�<���xj�J��C��?��i��!&'A�S\��!QEF�FNdP1�oӔ��Wڦ]��Hԛ�Ms����d�����O���d�I�|hZ򭇮(���Ӏ��OZ��2����Q/�.7-�!��J�ڦ��b!��#�0|�c��H�x3�ۭ���c]�@�Հ�?l��&b_V+��~��ǹ&6Qh�R5R�r��C,�~��K��?I��iC�"}2�OW�e���Z�fc�xav8/=��)���'�?�x���-�((HÏ��>'�Ř6�HT�'W�i���m�����4�y�_*x��pHY�x�i[ņZ��?����DR���D�O�$�Ojʓ_s@0�sꋃ$�.���m�J:	˾�1ѺiCxp�GB�^a���'d4��c�өM��C4�S���A^.������p0�ӫ��Oa�O�iibc�b,0�Q�Ԥ<��T�&�{ӌ��'� �i��zɟ�'6d�'CR��h8��*`c���S�' �[����I�g�DƉSt����s.�t�0�ӣ|	��'�7̦͝�%����?ї'�<9�늉4Y�(XdA�v�~�-�*��$!�'"�'���k�U��˟�	48��ֆ|��KF�qO���eg#`�h��gi�-CԼSB'<O�1X�o��{��!���7q+&@*��h|��\oK�岴���R��S��(ړ �,M�����3�'�K;B$>�q3�J��h۴=.����?	 �H�es:mYD&4$�3@9�?QO>9����'��'l� �%$�.���� �s4T�k��b�F�'06��צ͖OT�$k� b���$�O����ˉ2Nu�£���v��@1���O��d����$�O��	#x��)H�L��0%���K��­$n�l��@���ld":O�� 0�W�5@z�QF`O; ��ņ���\��i��
�te�?7�:)����%ҁ`ӎ�l�H#��\�ݒ�I.3"&���hy2�'�R�'�a����)T4R!���P�*G%��(��'1r�Ӥ�McD%P�m��Ȣ`�|�Y�҃�5
�6�'� 6��*b���l̟��',�D�O8�bը3��qSD��(��	#�r(b�'��!8A*�iX�(AĴi�ne��K�f��L�}�T��0�%	�
��O0!#p��z|hYIG�7C�Hq���׳+iX�'��w�V���0"~B�	Do�2��q�O�z����<d���U¦mHH|"���K�<6�q@�Z;zo�e��·���?AO>Y���?i.O�0��KLyT�WIO�Z�����K�'YrE�O$6��O��l�ן��B��*�R�;��҄)�Pc���M��?a�Ux�у'+ɂ�?����?���yW慮9&\y�Lȅ��d���φW�h��E�g��!Y����\>9k����3c��P��$K B����noF�KUh*�ȳ��D4
��F�+Z��]	i��w�	���O�,\T�iu����A��֦y�U����OPc>��O���D�^*��b� }�(Q���	� B���O��d�O��d5�3}r͗�g��JX�U�����?I�Tћ��c�x��E�����?U��_���9R�ƕ�#�ڦqp��x
_�z�@�k$��<_"�'��'����ԟ|�	�|���_�^�"����0v[ޕ�`���E�L4w�(���T�����
�A���;�G�Z����7�ٌ~��$ʲ�r~ݙgnܘ}�vi��MJ�0�Y$Aݝi�=�L>aA��f���ƍ
�.���0�+�-+,4�IƟ��IN����3$%�6S��5[#��8JF�'71O�qq�G'B�L�#�H���mq|�'w�����<�!+��1��F�'bB���xb
����ɤp�t�	K;?�"�'t�S��'�B8���G�$r�rd�#?�~���� �(�)S[�Dّ1G�:�z�� n"�oB�!��ʔDQ��r͍8)x��C�D�$��R�픖T�iD^-^����)��U����� �O��'�����7 �&A���8��hy��-D��R��!��8�Ef��Ѐ��+�OF%�	2 K� R1��d�#@˧:���O@������M�	ԟ<�O��m�'�'C��X-b0�ѻ!i��O�+�')Ц-��(��5d1*�� бTOj�'��I�(	z �0�?R渝� �8.��ɦI�qCv̿G.�}`�"Yp��W�ҫSbh���ҟf�B��F�x~��`�J[4=�IPu��<��@�Oj-'�"|��l�2�����,G�	�ddT�i�<A7'��,�C�ID��0q�l�'K��}���g�H��,V��$�Z��M�J>9�F�%S���P��Uy�%D��t��=Z��0KC63�t���ʀ|P�7mP�P��be&�|��$�US`٪WA�Ckܔ��˒2HN0�����Np�9W���v�(r��%�dΤAԚ���'Ĥd�ecB�@�<�6��[y"H��?A�'���|B�@�*(�"���S�Q�E�B�''��֟���O�� X�5��#@$f��$١G@�E���'�46�Ϧ�%��S�?��'��u�@]U��6T��� ��,n<����'���'�� g����l�I,۬�y�L�;:�|Q@AM'�b�S5�D�7�d<r�%��5}�I	ϓӸ�{2��Y=������40�$,�rF�t�X���P�H�*�/̯��{�A�cTz�N>Q�A�eܖ<8�Du�&`B�A�S7����9�MS��l�}��[�E��SMhX�$��Ia�y�˘'=j\	׋|iL��C�RUh9�M>t�i{`6�<YD��F曦�'�b��J�2�U{:�a�A7O���'����p�'�29��%�!�׃�LQ�i�,u��lZ8��ۡ��
�*��#�N:���tҌ��g�:�"�s�n�զy���	${՚�0�ŀ�a��AK�'��Uc��?��O~�+�ޔ�l��MM�r�ꁐ|��'�az�ńbG^	�>o��Y��%��'�ў�Ӄ�?��� L9�烏�,�rE����<�'Z��!�@g�f��N�'�?� �+pԢPړ�(9����Ƌ��?	�50��L�]�P1�b�#d�`�p�(��%�O����ɿs3N|4��Y[��Y�����#O�K�j[!��	m��yT�
�M���(5P�m�4yQ�j\�xV��)R�^?uVܡ���S$�O|lZ�H�P擞�ļa`�E"7�N��Ѭʈ�J�=�)O��O��'��m��E�B�U�b �WtƁE{��'PN7�BĦE��(�M{�O�8�X��J�QGfPA��[�u�x�yQ�iG��'�"HR+R$�1�'7��'�b3�X�X���A��t��*�W�������T��Bɲ4L�5�(���	���>��w�V!��AC�j֡5P0�р�A��G'ѹ_�@[��I7�<�UX>�#�4$pQ̻j��E�D�q���#�7,Ԓ-��NK���.O�m�F�'����?�O"���֠=¦��Q��'':�� 7�<��0<q�I\�S��zH^�0��4���X���I�M��i�ɧ���OV�E�j�abj.��y�IҳHh���Q	O�5�l���֟$�I쟔iZw�b�'�j?J�鴩��fMf\j�$� ,і��b�ĀN�B���5�2�E�[$�f	�A��Y�0��c��
f�A��[�)�.�P���W(aa&�_��qO�<��3�H��6��9�!�IW�W���<mz"<���Or�d�E�6jD-
��XX��H�"O�A-�4c��% �'��4:��F�|"Hs��neyrCD�&�67��O���ܱ@�2@k�Ș%f�ȫ�i�}���$�O􈃲��O��Dr>]v��O�b����"G�m#Ԭ7O���Ai/O��{#�ɴR:�`sJV�����E"����䛲P���"�DĒ�� �i�
Af LH��0C!�$�k'�t��LW����� @����O@��D�RS܍����y�L�¤�|�٣BcN7m�O��į|���Y%�?BJӕBYv�R�Lێ%�����]��?)��r%!Q��9ϞU�3�ޝZ6�,�C��~@#��.�q��4���R1+֒>%�� �O&V�[�5����H�+�F�"Նu�y��D+"�X
��M�$�'�O��,�0�O���'���Q��?ٍ���O�8S%K��uJ�"B��@A�'D��Zv������j"���5J$��?Y�	ZD��c�t�@��"�+)����4�?i��?�1h҃ �VL���?)��?)�w����'뎔Z7Z����'�`���i�9A�6��'�ɺ;�0@��K�����<�!I<I�B)!M�sF��u�X9�e�-I����'W \�6LXu1���@�ε��)�y�b�rޥq���'D��e+��	�+w��C�h�ڦ��.O��\��SW�L>!rhL�J��5��bC�TY�E�P���hO���$��LR�(2w.�|�t�qaʬ'�B�'86��m$���?!�'�`)I	W.r搝��k��"��fK�4�>YKw�'���'��(wݭ�I��l��5��kQ���>B�)&� �4��wMŊ�Z����M�U�����N$��O�Hb� �X�2�ȁ~�l��UΖ�J�1A@�'Ǯh�lʄb��1ؓ�Z�#���1��Ǹ'v���%j\�v��6��_e����\9�?16�i-:#=����3�\z���Tْ砈�`�rOH�b/�;D|�"a�wf�S՝|��n���m�Py��#����?��L�8 jn��1'��>�B�"��F��?��v�n̊���?A�� (�u�d��5(��M۴�F�0�v9J�I�X�v�`s�*���k�BO���"?�W�˂b�a��.��ᖷxR@Cn�/w@�) �ӧpv�5d�i��b@v�'z�xu���lӖ�d�C����VKipTY
��c�(��?����?�	�'b4c�H�Vv����b����<��4�O���M[�ՍL� =�a�6z��3�)a��_��T������OʧNG�U��G�	�"$��5x8���p���?Q�g� �μ����C����R�i+�O�4�[�V-����6.�!���3��I*]Y���1 ��1<�
ԪM��]��ԧ��!j�mY��@�HĠ�XB��p~�䃁�?ᣴi��7�O�"|j��'��ǡƎt����o����'r�'��ϸ'l��s�K��7����+p��������OTm�%�M3O>��(�	�=�a���Pi�D3̾����?9��iP�/Ƃ�?1���?!�;��N�%�ج��ڞQ��-S!f܆m�s1.A��dU6���y�,�Ӧ�ēq~Rl�f؉v�.%�k��>�(�e�/j	�j��~e���T�''׉'<��*C��\�L 1AgQ9Y�������d�r5��'wў�IA�X4K$�8 �9�d�qJ�F�<�3��6���ό1���&��Xy!,��|�����$Ǔf
��c gů�\��*E�a%d��1}B�d�O�D�O�����?���?�����1Cρ%�i�$��4&����#��q��ݜ|��y�J�W"�GC�/��4b�H�+�titǟ�jg��ؑ�9qg�y2��7@`�%ՂH�b,ƝK#�J)RNa�+O�U'�����'�L�I�y��<�rl�T�h�K@6!�z��Iߟ�S��V՟�����R�����u7�|�d&O�8P:EMI!�1KWǁ�m[�I��,��4�?�*O���G	\�4�'�h�2���#+��aw���nc�$�W�'�b�Ǎw�2�'E�B8��dy�l��M6������C���`��d��A+�*Ӊvi.�p��'��Jw�W�a�����H���qц�8X�0�5k�2 �B�03	۠�0<�O��>?i��$x���`'��␮�[��f�tx�U�r����/ی��&�O���	�X~��V�c�}�N�<����<yDI�&Y�f�'"Y>9�W����0�$]89Z��S��V�����B���I��H���U2���Rt"ٴ0r��.�/b��O�XJpA�l���ţ�;^�4m�Ox �m�>gӺ��D��[[���'��(ƪ�L?a�!�J*u�����I�[ZR�I�1?!R۟�S�4jZ�>}�'I��V��,z�}�á��1BЅȓ�flؤ���SO(��ՎQ�w�EE{r�'��"=ـ&A	{��d)L���=�!�!(�v�'w�I6d�pH�������؟ �'���Y���(Jm��A����{�Ց*�1�X�'j���p�N�>1�t �3̓��~�GH�o��9h�O�*0�o� ��S�ˑ�?D�u@׏B4���q���V��&=88xj��e����!�Bh���^s@(�ˏ����/Oj���'&�$�?�O���@�Co{:�gO�#���"�%D�$�BV�¡�1��"UY�i@��O����e���T�'��	<>/�x@�Â�8�t��D.ťKy������~W6��I����I̟ H\w�r�'��	8	lf1�%C4Ԍɸa��30*�f@[�5�ăJ����P�e�arf���^�Qh��Z��`�8�����ó�ˡ&6�u���Ր3��p©�%<�h�a#V�-���Of�#׈L;8����Gl����'��m�2�1�Ohu�T	�J��g�Ơ:8ݰ��'N1O
u,D�`w䀢�"�9/�-��|�z��O�ٺc�����	Ɵ���NF%x� !³�˞Z!�,0����Oh0(3�O�Du>�B�
5������\Y���	�+�~�K�G�� g[�5L��d��^<2���D"D��V���� H��1rfY���˪o��z�//O���S�'�p�O&���"�H�$`��C�"��xT"O������6�i��E8~��!��7��|jB�'�P�� Y�"۠ań�1U�`��L>�6��![����'JbP>YX�E���6M��,��cǍ*;;|���ڟl�I�8�����x e�[�&D�!{����T��O�Y��D�j?���ʈ���",��d�$7͌P���_�q6͊�jVH��E�_ �U�O��c�J����G��7\��O�9 5�'�H�O>�"`F!֚yA�-HS6�! D�2D�h�d�ȉIdʽߪ����'���}R�$3�ʅ!�۹jG�u��(��M���?9�f����o��?Y���?���yW@]L�=�Q�U4n��9��i�c��i�܋8����e���X��q�}·�|R�$_����5 �-6�|T�
}�T��&��lb:���C�.{Sڔy�����C֦	ځ�h�� z�Q�db`2G�-�`�A��5�D-�B���o	��NL _����LR��!��:jc���Vlı���.�[��':�#=ͧ��hM�A3��VՒ�9TG%}B0]�F�
d�ԭi���?)��?�#��L���O��Ӑ ��ўh.R��@o]�]-dL��JN�.�u����<�v�I�e�_�'�d�!4�],��2�L:tͤᨂ�5b؉�a*Z���!�%
�P3@P�*�Bc�0i�5ǔ� �)�2t� @�&gE�F,��GI��H�@# �M|FQC�F��_��3�a6D����m A� �3�,AM#a�B'�Ğ�9&�l���޽��i�O����$��z(�̡$MY
p��P��O��D�}߶���O��M\�l����`@�p�S-"O.�D �`��xS�h��HT�R8�	��5O�y:A�^V��ʑfC#M��Y��E�C5�IP)��5=�M�EA_�zax�ͨ����`~�B��~p�x�6�	 ���8U�M��䓏0>y1!��w3h"�<�ܠ
 ��{��D��;�R q�#�e<&���]�`����	DyL�a���'{rQ>5q����@�cз(�t���N��av@����ݟ����w�����`�?j?hH!E]4��|�؟"�'x(�a�l��)v�A�A� p�z��'�<�p���v�t�c0�Bk��{��̎�6��ϟ�8��aW"cx��9q��Y�Ahŗ�dSs��OJ��)ڧ�y2#K�wM�=)�+�*q(:�R	R�y"�F�dP�c�b�Fy��j�;��O��G���}��qXqF\+X�j(��Ѵ5��'2�'E�"�,S�;���'�R�'s��\�N�����M5r�IC�>T
�$�,aP �m��b>c�T��ę�yf��´�K�C����D�Z%F)� �6xn���T�IX�����~҄���f�;E���;�-	(�@y�G3`2��L>)R�����|�<A0	 �4|��f�����`/�{�<ٓ���<̐��'�A[wf�uy��8��|�M>A�JǱ� �goB�D�4b�/O�ĻWJF��?���?q������?i�OJ��$P1@�Q���<n�r��IB�zvЏK����63�\U���'�L1@@ދo����U�M#,8��7C�����J�i�3ѧ̟��zC�S��r8'��bC�� ��<Q��:	��}B��ߩG.���Ox�=����ƉC ��/�� Av�N�ֽ1	�'��@�B���k{,D�RσG�(q�H>I��i��P�bGE�*����O:RJ��pۤ��������O���O,u�>�D�OX�Ӓ(�*x#t*��Jf(��BH8�f���Wp܀�'�\Q�+��^�F���Wj�`�抛7�\�X��\�^��	�rh��t$�u�.�x OP̦�1aHI���'!
)���?q�O(�0�
, ]��xl��b#��Z��|b�'����Ώ;-}U�6�38�xh�y7b$O�i�u�GG�f�h��A�^��?Q.O.�k��Gᦙ����O�Xe�e�'�N̉�f ._i��{d)�`Ո���'	���}�,��KDXՖ|�FD��oy�u��CQL%��G9���RgZ����
2��0dc¼{̚ĉ[y�P�|��Y�c>�h�F��d������g~����IB�O��dªx��e��e_Ό2�_�!�dǋ��8��d^T����eŦџܱ��	ؘUńph���U<�Փ\�Е���?Q���?IBH�����?����?јw�`�BU.'|�xa�	�vx���d� !�ė#��9N���Ov@𙂨�?i�I�G���IE�|��`��a̤%�n���+
��0Ѧ(A�|Z��J~Jݴx���w@e�)Fi�j��q&ݢ
�<������E2R�'TўHIR�N" ��jgL�C���`��I�<)7�7I���&�S.k�8�vdUByr�%��|�����r�8��%��芠��F�Q�a��.pOZ���O.��O:ԯ;�?)�����e�<|�����&PE�-q��
Z[DKT�WJ�~X�"� � |�FCM�~�]Ey���x���U�V�CY޸c�	k4�59#�^�i'(2wÁ;�pM�u�ih�6m*�	O۬�2db�' �lԦ��w^���G�O������B����""�*@/��I�헩2��C��)U�,xx�	B�eg��	��O��o�S�?M8��O~��I�R�n8���I��k�⟠�'?2�'�����!j��EK>\�6H�B�Obxʡ�@�U��ʥ�̪#���F�'Vl}�%�[�" =��`
/5V<-ycԟ}ɾ ��H�y�C�� t�1�d*&ғP2�y�	ϟ0�'�<+�bQ�!�����CR�3��=�N>��t�����M� 8��	NFh���?	��4��|�	�e��}Z,�x��u�AnȑEUJ��<i7�ۦ��?��O���G9foh Vd@:�J\�O<^���'U���HI�n�<D���K�Ra����&X�L�A�J�^u��Qoچ}���Z���Ĥ�>�vU�"�2��0D��O�O����`�]�@ ��)J���x"�O� ��'b���<� t"�&�4"Q: �Nm��X"O��b0��0$<���FOn Jr��ϟ0Y��d��bo
X:A��*�ұ:D� ct���D͈e,���On�$�O�ʓf���ʎ*�IbV��y�X`�g�3XHvH١�'�� �b����Ϙ'
�eޱA+�@P�-ȯ�V�cņJ�b8�j�d��'���ɰ�O�\,�⫸>��k�%2��a�ɬ6iD�ٳ�����'jԈ0���?�����s>l��ǟ m:}���Y�3��C�Ii ��-5_�f�G�ɶ��O<�Dzʟ�˓n���X&�ň�aQl
�2���a���?	���?)�����~d�i���w�zt F�3Հ���ꌅA�5p��6	8̅�vl4!�ch.2�rVLC����&����M3���\\r��n�@�B�(��E�' *��e�y����M&fPx��4�?A��hO#<i`M�7S�ls��D'Mˀ�<�O*c����M �}��K"P;��E9�  �ďD}�Q�qգ���',v��M`�f$�R㋳����Jy��'�"�';@��@�է	�`T��J�*M�~�$�5r�:GA �`�I�Vcax�N�,�jeCC�Y-Rk�Ć(�|��PD�u�B.U^�K��jG#=Rh�ğ8�	f~2)��j��k��_6S1Ҁ+F͆���0>q�OZ�aL�&�Z��b� bdZz��hO��B��Ԃե��c��uqq���yp��ɡ��Ojʓ?5��1+O�i�D�',h�K�gչTh)�`�[eDh7�'r�\�6������L�R�4��O>��p��0-@.M��R��N;?kC�;ʄ�90 �/aq|((�E�<8�8�����9Fu�(��`�<.h� �EY
��$y|"�'��>Mϓn��8bN�`źu�B �<9��Ɇ�$�4��@
{�:���g�;
�G{��'2#=if)	9܍�r�O*��6��'���<I@%_&�?���?1���D�$�Ɂ��'���[�j�un����~�����-"�@ �D3�3�I�5t�L�VfX7�`����D�X�<\Z�p��ڲ�B�<�*7���0�O�Q�g჌QrQ٦`��a�x���'$�	�*�����O*�=�0��sJ��3X��Phxc!U��y�J�4 �8�r�bأBܑ��` �?A��8ӑ���$��,=1����\�3j'L �����nq46͏�	{���$�1(Z��	ǟ��'�B� ��]��������#Q�
�
G 2u0�	�!GD�I蟠�ɴW�p�`�BP;b��a��uڕҴ�=N�hxׯ�h���I1E��DTa�b!ʓ!N��4�ߴ[�@@�c-D����D��N�$� �K,p�j��I݂GQ"|���?ʓy��Q�����|RDQ��R��!!ʙP��3��ny��'�aj�aA�]�@�ҷ��1n`\Es���I*U��T���u������ʓ%��)���?�����}t�$�O�<�6G_vC^MaB�U���@�O��t��l�ژ���o8$b����c>���5�%�D�Z�^���Nt��Ad�)ytr}��g��I��)ŕ4Tl����	�D/���B�$55���H��;���˫*Dr�'��)��1?i4)-I�D] �Q2����[`�<ƃ�!t88�Ӄ�-6>��YT*�[�'�~":d�peP�� Ntp"��R��?a��?1���/<J����?���?��'�?��#�_N������d��<���7RYZ쁖b�%.��iH0G8Y
Ο���
���I�U��#��'�$p�Q�΁uZ��;o�1'$�sB遆�4�Y&a4B�ޞ9V��'FyR����0��AA,@�$��On ��'�����<��+E�'	��YEo��0{Z��`�D�<�5�>��!�	g�ԃ������4�����< G|��H ���f�&ęQ��?j�՘�.��?)��?q�����O���n>�@��2�0�#bDXx�a�C6$�ˀ*��`�6�CE�̾wtQ	��d�n����E�͌{�Li���}�0M� ��c�L��N��;�ĺt�}�'��K��<lEh@�D�-�V�b�j�1!2yZ���hO6#>��I�0�HUhҁ�;a��"�WY�<�PB]�t~dꆣ50�ˢo^WybFd�"��4?��Ċ��I�O*�I�`g`��� ��mz�e:Ԣ��F��N3@�d�O��dFW:h@��}<L�[נG>��,0u��i�D���� 8�.��$_wњ��5�ɘi��z�"L(����&�G�Ht�6͚-Th���4mJ�5En��0N�73�};f`�v�B�&�`#f �On�$$��1&���r\�S�P�cBY�`]���0?��E�����.S W�<�z��W�Ib���T�<�"�Ҕ>Z̪p%� ����kSy�)M�z���'i�Q>A���۟��}����'/��35`���p��	�Ip�ԋ,�*`#�-82��Oe,4h�ן�c>���K��V񬨱dIW�	�B�#s��V�G|��-��3b�-�#m�u���<M���Y]>�q�Ŕ�Z	[��խ1N&ȫw�r�����Or��0?%?E䧀 `�;��-�:��F)�,�B��"OjIp�&S̢0�c�2>�n�{���O�(Ez�OvTȉD�%�Ę�^��P'�'���'N� j��Y�s���'���'��4�'��vnͅ�4ѻ#$H�!�DYxPJ��{��iҌ�+\<����$������'8��9R��^c�`��h�)g, �Ee������E	�=�ZT� GȫZK�ӌ�MW� 6��;*��!aS�;������D�tqJ�'pduk���?���b���a�� ��÷EF��>�qO;4��p���/fRء���T407��֟ ���4�R�d�<1��ƴW�^P�������RG�~7$���.H�?���?i��Q��n�On�b>��7A�� t��D�X$=w �8��C�5�6=��&\�`��pEؐ�� )�흙Q���\=k�����E�B�rW	"!��(,s�ɒ�K:ښ���JƖK�'d���� �f�� �ʳbp�D��^�w�d�hD�iW #=!�����)���j��J�p0S]�%V!���B����$㒠�|�V"S,*��I3�M������O��m��t���|J"�X}2^XQs��*;0y�@E˟�"�E�֟d�	ɟ��p�U4"3���1 �;�-A޴��t�A�i�ʄC�;���0GΰƈO�a���:p���y��q(�''�r��G�H�Ľ3��sG �E|�$_�?�q�i��f�Ҥ\�5��}�)z�����O��$?�D�O����<1��?�6�V$����#X�8A����?!t!P�}�|II>���}ț�O�^�=�L�6\2`rN]��/G0;@� +O����O~���OP�$�O|�$�O��S��
�kT�� �B�k���V�¢?�ӽA|��"��*e��f�=i��ع�2��ɣ�?������)�[�Ph�@	��T�#-٦y��
�9�8v�9��Ɵ �SП��0�>�:�Q�!m}1W��/�ĳR���MC�<��+���y��K"�����KT�?ט�@S��sdDZ8~ZYy����$� ��'a����s�Y�	ɟX���lΓ&q�W��-��g,�2���ȟ��ɸ D��	��?�7�wnzݝ3�?O�����İlP����� �����ODӦ�'��aH�<��꧊?����u&.���g	Dsܩ��T!	T��gȒ�?9�G!��0��Lyb眺��ܴT�<��Ŝx��u�n��AY�����0ԛV?O����'��Z��|�$|��	��$��?^����)�+bϨ��+�m��3V���<IF�
՟T�	7�u�'��dE����Ms�eN2QɈ�����*�Ȫ1 O�� c��y�`���?���Q͒$�Op��'��9���zr��1�䞓3��M��A{ӄ� ��n��Bf���}yܴ����'���K���t��]PQz�H�$IT�D�G,&�� ˩A�7�	ҟTlZ�"۴s���T?%��	,gTmڦNP>V���YQn� ���	�'m�	��K�Wq��@��w��!��4�?a-O���O��D�<.�k���I�Z��c�B�z��Y��A�b��f�'O�'��-�~���?��?��Ug����ci��n�qW�����'I�����I�������Iߟ��dǡ;,���c�>
W�_��MM>)��?!M>yM������7��0�F��WܰMAek�`�$#�(�Is��O�q�Q=����ʗ����S�(�'#�'��D?�7Bµ��t�HͤO�T�񕡂c}S�<'�`�'��}z؁�%CT���A���&|��pur��� #����SK׾?���ȓ�~�����C4$0#撠�*���Z���+٣�mR�n��W3�̇ȓ���藅LZM�z�K�m�(��#��P���a$��W�Uc��?Q�*#a��Bb'�&"��@"aIT4"����#	':�x��8#{l=Q�" ;!�`���8�@]���݅.���ӓ�0\��H�H뎅Qs��(z6X�>�'�^Tb��iR�$�>���D�ą�ա&�
���T�h����'M�S����-��G`�h��al�4Z��0a������Y�\�4�q�8hUJi����#i[������С��(SN)�G'ŽM���1b��ih�dۆ1Z\��LD�6y*�	æ��(2�Q �!	�F�^�l�e���VbD�͞4���F�2N�2���?	�ſİTjC��T��_y���O�S'E�<�i$4#��R�Ĺ5��O���#Ւc�)IV�"�^����)�S	^
^���g�!D�����o��6�O��35�'�B�S��q �Sʹ�4�3x�M��A���xrNݡ\�N�)s��I8��w�Z�<�أ=�',�Q�4�� Ϙ`��ϝz���$L�]��'�r�'-�	jc�7=��'�����f��� &��h�&͈��Ձ!ȡa�`�>@�D�/?��xR�<)�x���NH�0�JX�"�%h�~���͉"X��,sp*
�M�����L<��ܷZ�X��o�� �x�EH7=��7��ky���?�'�r�}Ra	�=���'Iڹ��I�p�@�yR.�45 �C�~��}� �P��~b�'c�#=��Z���'�.�q�?C��@裦�.n{�!q��\)u��JM�O�d�O��$���s��?��O�Պ�l�u�fHK� h���`�i�1O�i(�i�!��� t.��F�џ�c� $�ѕ�W#D�`�C��4@�7�[�):Ĉ��`^t}Yc�MNs�!�V��8w��O���eA� r�a����&%�5�3�[��'""��&��6�:=�U)�L��H��OI/�C�� .0p�_��LR#mG�F�Tj�4�?i(O����K���id1c4�G�\[Ɛ�!S�(���O^�䇆�����O<�#m)��	�̃8 D����(��rc��5t�<� /X������{�'� 1�4WkN`+Ae+d�8�S�#��$�A�D��mUL�Kf���5WџH��'�O&�$�>�eM�$ �Y��j�|"���q��Xܓ�?�^,�5@�L�zư���a�tEy2�i>M#�`M-%G<�Ǐ�rȐ��"+���	wy2M��t�����?�(��� bw�(�4�4*�)�P���RR۟�	�3�<hN4<�	��요3F�5�Zw����[?=cҊ@�G3���f�KR�pµ�?��3�|H�u�ٷM#�����-,�t���ĺöȕoD��GChi�����^b��賑x�ϫ�?����h�(6��?��D`��v�T�a��j���ȥ��=���P�ZTTꝡ6�i>�;��D*
U���L�����EDޭaF��4�?���?��Ǉ*� ����?A��?���5mT���*C��F]
v�ʀRq�(+�@�9��T�2+�8P�h��E�!��Oě��
�?���7/p���,٨{��%�r��z"�S��W�LEDN�
|�!ѵf0��q��:�w���CG��-oPj$:�o�������On�t�9�i>���L�
��%:2Jэ8��!��-a���ȓymV ���	3z�`���"DS��1�O^<Gz�O("\���2,��"���J�!���јwB\1����?����?��M���O<��w>�B��G�f9!���� �$�[�C�v�R1��
r��z�K��l4��E�	В�:t� �˭m�@2f�y��� S+N�9���U� ,K��9�d��,9��	G�V�z"4����[H�2c��O����O��H�~ӊ��7󮡃�(X7O�>�����_�<��
��� `�N^�����Up�1���'��	�T��!���*7��&r�y��f*8F(q�"$ȃ (,��ß�s�"�����|R� �&1Er��!�Bfh�{@Yu}z]K�@�/0vQ��0a�|�0��D� ��ٴ�ĂT�j��'݃7�^A�GS,p��@�
͂���n�O,����|O"���'�RP�� Gӵ<mr��%EE�ZXLt���#�	�`��33*��a*>�(8q �ظG�>�<i��4�2UC�Ҥ)؄ը$�CS����@�,��<�#�׺9�����O+��㥹ix���V' �.���BG�T84Y���O��DMZ�*�BΊ%,F�U%ƚg(�;���騟����P�"�թe��z�d�ڥ�xbJF�
��I��M�U�B�jc
 
����v�h=��Y�� H,�6F�����[�m<t%�ܫ�!�OJ�D%ڧ�M�T�t!r$��|�^ЪuFc��Q��'�ey�(�u^0)Qo]6F�lQI�/�Q��;��=��t�� �p=E�E��~�z?�U��?�����'�x�I�L |B�UI���B�F����y2�O���?!�XF��4a��29r�ȋv�<����*�P�j%��8V���z��Es�<i�/�
{������4gf,R��n�<�fȑ��^�����0Y�q� ��U�<Y���xW`9X!O�,�|�ZR+�T�<�P
N�^ռ8��,U:��ŦW�<	� \6�z|�eE��L���GkL{�<at���V�<`!���c�P�q$�@�<!�M����D8⇟���G�@�<)���0F� ��x	k'"�4@�B�	�t�´"@h��}H��9T�/
b`B�I�c�"��BFT�(��T0��B��6l6�-c�f�)i��u�g�\!�V݊�n�5CPzȂ�'��%�Y��J�̽֣S5y�CL��=��'E*�1p@�f���kt-���b�'ަ+���>rXޘ�DC^<t��,`�'F���m��3>D%�#*1\ k�'���Ť��-�X��aDi����'j�r�j��s,*H�A�ֆg)��#�'ӞId_�����TX�:X*�'O�Dp���6�$tQ6l��XH�'j��kP�_�f`#&j��@��2�'Ւ��ȐPo���%�t��Ȑ��� �-�t`kl�!�ĩS�<���5"O�b��>z<���>>�:$�"OJ8IJ�,T��X�e��5h�ʅ��"O��yr�Ǩ{�|�2Ɂ)q��K"O�Q"��Ⱥb��,C��;Q��q�"O^9!��I��:"g�1V�R}[F"O}p�dXq�㒆*�
`p�"O���@ɼ5��Pr��R+z-�Q"O��dl҉#��y[�`˿o�@�!0"Oj�ʑbՓD
���钔>�$	"Om�dJ,tՋf��鳀"O������> ���Ԧ�/��"OH�"�8,jT'۱e�(d
�"Oj�`,
�J���&|�.�a "Od���K�l��,A�G]F"Oई�EQ;R�T9�FѠ5Jt��"OH �&ną~H`�Bc�l���"O"{��]q��
ug��� ��"O� ���ЭLp��He�Y�^h;�"Oi�%�ݟ�͈2��~�.|��"O<,�ե���I
'�ݏV�P��""O�9���܏��mC���(��I�1"O��( lB�_a�u+���/�	�"OTPsmN�M#�u��@�Q8>�p"O�`+�MM�dY�H$B7z\*g"O��f�!x�m+!	X�K=��b�"ON�@�.[j@T �ǘ�!��$"O��S�*��=�c�Ң&g|�0&"OL�)�CL 
��a�!߬
�C�"O�E�+ٸy�<�� ��i��#�"O"���"��uY�բsfًq��k�"Ob\yu�9S�J���Q2t���"O�}��bޕv/,��T՘�Ի@"O8��N		7DZ��CF����j�"O$4���*g�b��&�M�5��T �"O��pW�ݥ"z���9�Ȁ��"O��Bƭ�:�����A�]S�"O�4�7b�e#�t1n��Q���є"O �7�N	].�qP�CL�]����B"O�̈� @D�n9{Q�ц[�jD�"O�x�@�s䜱��A�@v�1�f"O�"�I�d�%�P�7�Ѣ"O��qT��2܆��P��04����"OL3穕�x�`egI1M�T��"Ol}X#_�5�*�9���-P7`���"OB�㔈�8�|ɵ���T���#�"O�\��.�a
J!"��l��-R"O�#+�;�LE"ƭI ��@�t"O�e��#��#Y�LS�>�3a"O��
a펕~�H\j���0r"O"�����t�6��iݚE�����"O�mPEjZ�k���I�Hs�pB"O60���n��������yT"O�=RD/M�=7	�)�7�D+p"OZ���(Md�rܚpiU���7"O�i�j*�I�/5+j�)�"O`%��A�>O���5/��_�EX�"OzQ؁���6d5�"O:({nQ� "OpE#�l܂)�4u�aU�`��:�"O�b�K'g'v�4c�>0��"O�drɉ��T�'JzI���v"Oj�Cb���\����F<�̲#"O�lH!��N<4�"4��D��� "O�)�l�2c�X�c
ָh�|��"O� *�3t��d~�Ӕ(
 � ��"O8����%36Bt��"`G|l��"O.�#�T�9g�k�ƒ�v��I�"O�=["��1z�@�"�^�n�8�"OL�'C(RH\���"�9`B�!�d��53�D�tm Cy`�S5#Szp!�K�!�n�����s��×bE�Kz!��G�zY��&G3kX)�`��AL!�U;x)>��
XM܈�b��B!��W��h���]�unHs&��m+!�$�5|���	�D�<D��EW0!��ؘ4�����ۜiŀ���bD/o0!�Ŭd�DpS��(L�Vq	>(!�DP�`�nxb��Ж`��A:%��!�F�!i�8cu�R^~�iA�nF-!򄆕g$@`QJT�Wbb �B#X:'!�d�%d�@���!�*B+���ÂG�-!�D�)@B�b�	΍'�U`W�P�!�,��{��åX�I�j�7)�!��©V�@)AD�U�z�(�r�J�J!�� t���	�$P����C�ʆ-Va!�d��u�v߃ڊa4隴BE!�DzԈ��iյ}<�{���|W!�$�:+Rv�e�޻$<�*�F�4F�!��ƶ�e����T�sr��3]�!�d�9H	���ɑް�dA�!��:1�Ri�J�;(�lj �#4{!�Sl�|��A*E�w@��ۂ,%�!���0�@2~6&uy1-��~�!��l��5�"���3���7KP�2�!�dJ�-sd��sB!q&V�jS�L?}!� c�t�U�
�JǪ!!�F+>�r�"���rpjƦ*!��N�Zf��F���LhX�M�*/!��D��a
&�Yt�q ��C�!���?�0!p���;�4X#Ϛ�v�!�D�����Nƹo�N��N�:q!���UŜa3�,��q'��*!ß$F�!��Q�:�<�@��]���6眻q!�$L�E���g�V㼙����EL!���C�<�k����v����E�Ue!���q��i��_b'V�d��!�D(`�Ҵ����/& �Pf�մE�!�$ƭE��4�Ru��"BƮD!�^?J0�C󌐱QL`�� C�l!!�W1X�
a�gG�4�p C$<�!���5(x6��3�Q3�-#P�4Cw!�d],�dq�#�����MU:'�!�d�.&*r �ا0E��A��
6gr!�.+���S�֕Y(t�ze酀|m!�$+m��Ac4�_tlBĸU(Cb!�D[�s�ȽK.>H\�!�!�O!���>�䌘a�n�" �E���_K!�$\.f�h3��z^��2��2!�F�fԁ(�
L.��"�����!���	BI��@àD,O��s�d��!�D�e�LP�Ƈ\�)茠�6Å��!�D)%״�`p�/$9P0��D�<!�Y�h�!c��3�<̰ `I��!�Y�άcD�EfZ����8�!�Č�A�H���cQ�)F._*x�C�'�p�aQF�i��D���bA�AS�'�Q���:=$R��c��=R�����'����nX�9i�)�ٶM�@}�
��� ��	��G� �@j�#ʚj��[�"O�,�E�O N���3QЮI�"O&6�+,����N�2���"O2Y�
0���ېc�ިɆ"O����O�{�V�&,�,X��<z�"O\9R`��J��Q,x�\I� "Or��Eߙ0S�i��+��|����""Oj$(D9T���YP(_y杢"O�Ux7�)X���(��
���{�"O���lR݊���ň5���G�RP�<��e�;L5j̠4
�Y�5!���u�<Q$M��p�~h��Yz�����W�<a��Ұ����s��WO��#%.�V�<��-Y�Pl��{3B�B"(]jVg�l�<�R�^�������ۨ�Ra[p�<����4ҵ�XuP��A��m�<aSeG�S��e�����5%4�9p��}�<��&O ����R5��99���w�<��#�HB�I������%�_�<!�e�*2h)`�Q$���sCA[�<)PC�}�9R�(W*,;���2�Cn�<�"l]6�X!��,��(��@Xt�<�����m�!�A=0�8�!�ĄI�<)6�Y��t���o@c<2���hE�< �E�"���̓	<�����B�<1�B6'�"y腌>3��(���y�<1#��%i�ҙ�%�6.�8�vb�s�<�vO�C��
∘&�ƙ�F�Ny�<1���E��J!��4���:UEN~�<��U<K�$����6����x�<Q����RВP�V�rtL݊e�s�<�"L�7،�τ.f���aZr�<����v��Ƨ]s�<�����l�<�egB�*F�x��ԕ5c�t�1'�j�<�u���a���V�xp��aB�<)�@�JjAH&(đ(`q�CJLs�<q����8�v.��l�����Dv�<�V�߮Jc֭z��ˇD;lTXbN]p�<��k������@���Ǭ�h�<qmI��JTz�$Ăk�f2#H~�<I!Th n	դV8]3����]v�<�`fךZ��b�R�<��ȹf�s�<�b .���G^�x�Ƽ�6�n�<�Bg�j� �{q�K&�^ŋ�n]u�<��@4e��e*��2�l�+gH�9Y�DRTd�x��(��Ϊ��<qЂ�f���1���!��y�r�H\�<�I�:TQj���m��5��T�<A�*D̖ht�S��+��ñ�n�<�SN 0f��ʣ��%~���Շl�<�M�>���`�!V>>�&c�d�o�<�O}�]:�l��d��\a�<�iN72��MS��ĥ�#
{�<��N�+&~^�� ƀT�D���l�<����PP.!��_r-B�e�e�<i6ß%)�� ǋ��5YRa3�.Ye�<a��41NX��o\jצ����W�<�Q���2�,iqE\/H��@�2��Q�<�C	�
�ZIx�Gҕ]P ��g�<qvb_ i@TAp`�+l�lZ#�DZ�<���ny��r�%L({�ţ�p�<A��!��(-%W�����	�P�<�4l �O�2���¤��Zr@j�<��0g#ȣ�ԾxR��#0`�c�<qQ�'��dsG�D��T����~�<� `���� E1���
5 T}0�"O�ΛyZly�;�p�"O&m��t�fٚ	���0S"O��Ag&QdҜcE�7��Q��"O*��!���< �R��p�$"O����)�D���%��!��eȠ"O^2� �e�"Ls1�R>d�"��$"O:@��� Imbi����{"� R"O����Ņ�"��B ��"ORT d�K��x����2\���"O��Q����<[�C�<��<jU"O��
�+�0!�H�C-C��Ya�"O^X²��X�1rg�"̅��"O�����Y%�Jy��hp�Q�W�	I���Q�-B��`&�D���a�,�ybEګ��xc`�	��-�y�/�3j��uq�$ϥ>�^� �iH�yҫ�%�R��;�x�����ybnM�.���樓>
!� Ɏ�y��L��p` '�
r�`����y�:j{��e>�tuy�j�+�yRaTdg��s�%�� c��1�[��yb�^rX��6��.�
��P� �y򤟗U�dh�.��)TF���J��y`rB�ey큩m䱐Yb��ȓD�f1��g�3?��q0�G/�p ��P�j����)��ԈV�|ht�ȓB=*�i��T��ɳ���m�|9��
��)�D�I�)���+���Z���$a�X�S��#^��9��B�n���k�����-�ykQY��j��]�ȓZ��7��;3C��:��B�W�}�ȓvE �*eɌ��|Z� ��,P���!�j<�T*���%2S��? �����e�� �CA�eF6E�G��?y4�݅�=Q@�'@ƃzt2��2���[��ąȓ|�(��WN ��I����1"��ȓ9լ�ʖ�1g:.�Stj�]W*)m��y��:�H�[��̀��B5�0<q&F�42��<���,{PV�P��]؞@�g0�x���H��Ii4��ɇ�r"5���4.\D2�I�xb�TH��`�����<E9�-�1��'�p�tȁ�r=��ہeN�C$�b>9��B.6���A��N�ܔS !6D�I C��
��mrV�Eb[��y ��$rD8���6Ge�4!�q��`F��Ou���(I��0�G��/b9j�"OPL�u�Q3ft�3�����3B�i�n1+bdΜn2�� �g�'X���G"��L�Z�$'C\"v�a{�K�d��J�
	΂hR�bцp�����ko���o�6%n�C���$h:q�;n�؃di���b�X�J��8���̉w�ȸX��D�4Hu��磈=�Hځ- ��yrF[�������ƚ9��x�Bc+'4�+"oD}�aN���Mcg�>��*Z��1�� w�v�r�
�X�<�nQ�h�v�X�jޫaTh=[�ަ-k��>4���z7��Gt�	Ó��`!� ߧv��`3��;8�@��ILFx<�`�y6��
D:}���iٟ`������"�����'5ڬC��ڭ{(P�;V���}��7L�0�i�
�*J�~�8B�(����;�/��,�ԋ�xB��)�t���h�6G�`�4#L=EaȌ��L��
��\aq jsB6-I���$�Q:���Y�I�`z��͆k!���)�,����V�L�5��4��9.�����^�l��5�
ÓY8\��0�� �z�2B��b�	��I?|��PQ��2���'K<��rj�I�@��W匎L?2dA�'��|
���I��wE��n�����}"���=�d�a�-�;s'�9�G6��Hmf���U�?U�帵�ز:�`B�I�)B�Y#�^L]4�B�ƙQH ��(��f��O�M W�i�"}֧� Ԁ`�m¯lp*=�A匨h�"O6��- �T�I���u�Z�9u�iո�p�Z"~�V8��T����&�f(�P�Q�� A%I۔=j�zR�W �BH�2m��J�H���
t*ܓ��׼����ÁY�����p~)�fb��gC@5�񪖳h�p��=yQ�I�ޅ��C�H����Bf2%��dj��%{g��K6"O�e���*����GM<2J���J�9�@��c�
�~b�����I�Mk,�J�h��D�Ʀęh�B㉅�<+cNM1	�|�c�+�b�b(I5�ٓrf����<�����9� ��I��`��cB7 �(��]�6˰��5� ��ɋ ��'��!3ϞK��-9S��	o!��E� �R�'׳D��H���=Q����U�L��P��S�=���q���J��\hUy�!�$��$�i�u��9���pZ��H&��q�ט�"~���=: �	�TQ ���"��4�ȓ[��xi&�H� �`hj'&^��9���&�u��6��ϓa7
�Y
�p����y��	�Y������oCnZ'rE���-�Ws������^� B�	��FR�ԄMx�I1I<q>jc�LPG��Pri%(X1�6p�}ZG�4�J�R4��*�*C䉜&��cӈ�t���C�jӟa��k�v(C�@��?B�?�gy�i� j��iÍ֥"t�r41�y�+�![�^�4�Q�/ ER'苃�M;`�+C�&0H��j|s��d�0e�Q#i��Yu��5��N���Q��%�L�Xt,@�(YP�&h	'�l� ��֯�M��'���VDEj�:����I�RB� ��d!@o��RLU.*:�±�Ys���>��X�!^Ω[��_E!�$��VA���T�S�R�DzD����"X�*q(Q��� �����4���pg��"���	��(���:�N1D���G��z�Ab�"�1t$�|��芰
��fF��ACJ�7(��g�'d@�
*�0���ɜ�Q(��	�u#4QjË��,�9&�	\}�a0fʠ j�qdł�#R0��	�Q"�Ã��>oؔP0��O9���Gz���L���wa�,�(�Z�~j�y�*�Oo'�a�����!���b�8��F��0"�L d�Z\���C?(�	%��$ &�4�S�O�HY ��au
!�ѯʙs��3T"O�Z�%�	p\8��9h�A��Ű<q��Jd�4�)�w���$�~��耕L[�8��5��؍�a~R�V"�`���>_b��T�G�_TZ�ybC5W�Z���'�DU�f��Lrbxye�D	Z�\칌�DD�/���� /����OFP��R�(P@>��3\�Jp�8[�'Q4����^�L52�h�=7 x�/Ox|1��X����(�rȋqC�L���� �,n6�0"O��اiёNa�������r���G���$̕{i�|8���U�ee�2� �ȓ��䨧E"!�"�>iZj0��]�ȁ�c�7 ������:L?���j��X��߈1�*���[3
��G'ܑ��dٻ[*��U N�ZԄ�L��0��.����3v�0�ȓ&r�l!E�1L�ɸ��X�V���ȓn��L*Ҍ�� 8�����`���o�&�cW�ԴBnq�u��,ʡ�ȓsO���6&)$�pA�Q�)ծ܅�5@��bS7+�zD�A�T�)�j	��tKذK��:p2	�,��FJ�ҥ�עd�
F_�/ ��ȓy��l�h� �ZP"��R�21��*�6���m��X�&�X,^�6��ȓl6�01�'E�%F���"V/}3�)��W��#�$(T9��+@ �j���&80��TB��Y�MN���P�ȓ$֭q� A�S�>���fK4A�x�ȓa~<p�e	j/F���蛻&;���S�? T�� ��:C�J�� � �u�rE��"OP�Ks,Y�Q&b���
2q 1�"Or��gN��&�� �8b]r4��"O�$k�+�0f��y �+%�(bB"Ol��Q$CF
�l�t�H)�"O�=	�l"W����E/Kf���"Ola�pkңt�aQD^�-�d+"O�%s�H%y>�dw-�1�-��"Od�J�%�=w0���$��d� t"Oq*�O��5���(;Є�6"Ob"�k�+t��0�A�H�����"O��H7ʘ�Q���b%�$?�h-a�"Od�!�� �W�z�	�Կ3| yj"O��Ҥ�ܔut01�jҌ7h��@�"O|]�)D�q�Ji�6J�:�lKe"O�%�d�[��HB.B�Z�b�R�"O
�"�V�F�pհ�-�"p�}	t"O1���՘]ӧ�Z�I��iZ�"O����ł=Ocu�T E��=�"O���V�GxJ�H�f�PZ�L�6"O����-C=�akk�`�>%�G"O��2e
�@2�@[�L�=j��q�"O��Z��ڿR��0��t��0y�"O�M��o���@���"E"O�<C���c� �H^�j��b"O@%á*żh���0u��"W�^mQ�"O�%����L�d
�[�|�3"O�9ӂI��@����WP)�Q"O�ѹ�'Nr�T<P�b��q�,��"O
+7��<GG��ѥA���$B�"O���D͆w(Ȳ�'�P"O<\��
�!<�q�F��K�X-�V"O:�P�T'T�@e���$?S"Oڨ�P� /x���Aѱ	��"Op�����8��9Z2A�"	J��4"OLp����4u��	���mj�\��"O��&ǘ�p%�0�v@ѿX\�$AE"O����E	'��`��Z7 ���"Od8AM�A
f��2�6r�x���"O��!ě%��&�Ⱥ!J�"O����B�W���hT�aj(As"O�X�		�B�0P���O��x�"O�a�GW�}]�z �	)�LiCc"O��� mG3a: d��N;���)�"O�,���V���ɳ�N�e�ƍ�"OXy+sM�Fq��Ӣ��[�<8�"O6$"�L'G�	jD�U��H�w"O�t`C����psNC�uv�8��"O
�ˢϮ=Gh��͛ic�D�ب*p��q��9�<��4b'<O����M#F���m1b��P"O�m��W�:���,�|
��s�"O`������ޚ�Z� Y�^'l%i�"O�@�V)�;J�1"��,E;F"O��-�\x�؃w��E2&��"OZ���DB�QK:tR�`�34���E"O�\@ 	�9	j(8���Ȼ%"��1"O@����i���5��!0�&"O����*s� yaN5*.`��"O`�x�=d�@y���'Ly`L�Q"O`�X!�,'�n(St"�4i,��"Oz��w��G0�3#Of����"Oxd[�o�>n�|%��nۀh�l q"O�	�u@�E�UB$����"OέKjF��F��)�1��ag"O� N�Ar���0�R�a���"O��9d�WO6!J���"�F��"Ol1���X���z%n_�"�����"Od�����I����F�f����"O��+&�!=��8��T��q��"Oֽ⡆��4SH��֮F�|�b�"O�9�`Gڪ6�=Q猌9Xְ�yG"O��c�4ܦ�2I͈m��t�"OV��4gH�;�� �G�Q���"O,l�Q����1����.�H���"O����n[�TQ��w��#iØ���"O\���ER��%��'�.�;E"O:uز��	�*����"aЄ"O~̡�W8,�>�	1ℕ⬁�@"O�\T�D�1KZ��&�U��@@�2"O$��W/��PO�)�ԁT�`Ӹh"W"O8Ċ�M͛q��5��A��8�k!"O��X�.�8�E�Bo�+fW����"Oli���O��؍{�͈;QHN��"O��[�*�0<�0�����	>�M�"O���r���F
�u'O&x5��Ң"O����		;�r��wF0]��AR"Ol��2��Y~���$ݶ ��A�E"O�DI�I�Y<~���I���Ap"O�u���[u®@Pa�E����A"O� �F��A,,}��O�
I.`�r"O�H)E�ð�����(P�h*��h`"OXxSJ�Dt0 ��GT�$l��Q"ON���<=2� :�g��M��b�"O:<�A�=�Hu�$�*a��ٙ�"O$y�'�¢&��`�=x�d��&"OxT�s��
�4\����.(��U"O��"핅xp�� ��C'~�K"O�I&��--h�B��2"�L�"OQɶ��$UCh�CEC&d��"OD8���Ζp�f��'��`��y��"O@-A`*	�Mj��2��K�0� �f"O.$�Ν;M���!k+]a�a"O
m�F̃dHh�)bv��U"O yT�[	bt~���I�o'PQ"O\�"c�����`�(m����y��	*|�5`�˝F�8-Rb�U��yRڀ0P��c#�O3O�|d㱧T��y2��;����ר7�X�D��y�욙}������4�Y6�L��y� ��mh��(���u���[����y�[3d�B�#�)�#f�v\��fN��yAPC�ؼypk�6e�8-"�&D��yrB�;^X貯ݜ-�����)P��y���>��"��ù<�f�a��L?�yB�A(�$5r�o/`Xa�q)���y���%������	 �3�A���y�Mmc�����&gj �*Q ��y�H�,>�)1u�K�cZLq+U6�y�'+��9��b8ؕ��f���yb�Ɯ~��=�3�K��ي���yr��!O�T9�Ĉ� {�%ʒ�֔�y�OX�fQ��(�נaQ�`�Ѣ���y�˓�l�dX)�NO�*AB��@�Ζ�yI |�|R�d܇#%�l��g��y���4�!�Ҍ^�r����Y�y��s�J��'�,(rI��K9�y®�t��%��#�2���.�y�� ��s�ꀬZ�^� ���y
� 4Ir��G�{S,� ^}U���G"O���f�[fɪ�/I�%P(�k�"O2����[�G�a�oVu��""Od8@,̐y�2�2���4�rXc��Ox�=E��,̥Kʚ�0р_;��I��M,�y���$��%w ��,�Lh[1]���I\X�0���� *U"$��D e 8@��*D�<�H<w�H�!&$"�(��W�$D��#7m	�{{l�!�$LR��#�"D��f�a�<PX�-r��u{�%D�X�f�@�$�܌A��Σp~�0�L#D�d� đ�6�ˁ`�����{�O+D�����/,
�� ��KTJ0)��*D���Q%�-S�%�6�\�P
$q�**D�T�3#W`��(�'��!l��ݛ��#D�$з匲�X��׉���bb� D�<����,�P=!"CW>)�J��S D�Ԁ1 ��.h�T��D�ń��.<D���Wo�=����3��vf����/D�\���-�$i�w������y �7D��"qȖ) ��Y�c[� ���+D�|�֫��By� аd��'� 4�+D��S	�+C`X�G�q�΍h�'D��i� cw�Lq��/L�l`�G$%D�03� ��$�ZF߳}�PD�Cb/D��W+ߺ_l4��oɗ"	0�q-D���a���0��ۯ9���ZrD5D�xs��֙nlFH3c<:p�%���4D�\�⊀�ly�`S��.	R�q��0D�P@��	�f�ҽ� *Ԛ>���g�9D�� '-]�#�b堡�D�#۶�jv�2D�D���E���#稁�օ��y��[�K���b�V@���y�,
��Hd�8vN����ȅ�y���>� P2�V!W�B�z6,�6�yR��5�d�B��D&`U��G>�y��1TvpICJ�K�D��厈.�y�K�Zk�hG��Jt�43����y2ƒ�X�z(�P+
�v|*\ѳmʷ�y�k<�$31.�W�
���yrAV&F%��cT�V�T�E>�y�
1~���E��N�
��G�y�ʇO��|��B�6ԤS�S�y���f�`%���Ό+J��#L7�yB��#A�}�B��T��`��3�y�%=v�T=��B� w���n��yb,�&�2������nR�Თ�҈�y"n٥5dJ�P�;k�(H!�!���y"��~}���7#A-g�T������y""_d�&�������U��̔;�y�n�Hv���%������3�N��y��֦*�|��M	�RP^�#�[1�y���Q�t�IO�z��+�yR�@!?��� ��N��%��y/X<��H�šԸBm�����&�y���BU�1Ư�&7�r�J����y�ƌ%�l�S�̞�]�X��.�	�yҭI�b�Q�޹Z\���1���y��@#r��Ibŏ�H�"X�͉�y�aƚY��l��DM�@EREN�y2�	�b2lTH�g�*(a��@�AR��y"��>b�(���C�o��]���Դ�y�	C�ƌ[p̑��H0�b�2�y"M[=1�� ��t��P�k^��y
� V<��J� RC�H9�ᘶK3�("OؠC�Uz��1��|I�"O�qJŀ����̂L����"O�u���R�%(��.@9< �1�"O	 Ï٘b��ԥ$dD��"O ������-�z`��-πnP"5*b"O4�@�M�^�� z����ET��"Oddp���b�d�Ǭ�F���"O�����,'-�C�E��>�c "OZ$jC� '��3�C�	#�	�U"O.���+��N��x��S1|�h�p�"O��P��� �Tdat�́u2�8��"O,��F�ٸR�0�+Q� \�A�"OV�	�T�6|��!��T���{�"Oڅ) X�8{���K�1.�#�"O�<�`��^���㞦~�l��G"O`]C�
ì4��K�LY�B�t"O�e�$K|�٩GUL��H�"O~9Qm�0/�-�r�ћ�I"O��P��[9��<�S��B�b "OP�9TLީ#qĩ3�Bə���"O�ŊÍƭn�dP�a�G�{��)"O8�{�+Ʃ$~�1�OMB~&]IE"O�<�aC��>��g�?vl=(""O4���Ʈ��9BS�Vv d"O$-i��=[H ����;>J�b7"O��0��Шv*����W�H��]�4"O2hX�e�,l��}3!͂�1X�u"O
���	�Ɗ�P�+ԣ()�A��"OG4`����7J��e��*O|d���M�e�\X1�`�	�l���'^�Ad$�R�ؕS#�	���(#�'}܁{���^�
����G+'4��'I���{6�$�b��:'5.�'jM�g$ �c��Bb�K+�ZL�'�-�p�R	
�X�3�J�-Z���'����L3��0�Ѯ��"�
�'f�c���扚䁐R��u�
�'�(�L).�"��&-� 7�(��'��	2 a�0[�v��k��x:aH�'*Tp���9c���ň�~B�'��,���V2K����"ߢ-2�'�0���,r��
�Œ|ʤ��'N�0פ6c������<eI�1	�'H�a ��?yz<S���,6i��'��:����N�Re��V𬠠�'~��c��+Qox�ǑP?�͈�'5@� ��,!����^�4�Z�'��	��!)��⨀�Z��J�'��$�Eg]3&�d
��6\�i�'X��
�e g�ѷ�ܑYS0p�'�P�[RǗ� ׬	��a#D!K�'df�� �)��[�DCy�i��'o�9*� Ԇ��p)�?r���1
�'��-�	�.��0)1��c�BY��'Sx�(Ca�7`���C#DѼa�
P��'�d	bg�0Ū�S�Q�4��'�����ĝzt��XB ���x��'%\��0)K���1Ƌ� �v��'����E0x(�!�
�k�2M��'�p�(0���9���ဂ#i�x�	�'n@!Æ�[�?�f� ����`�'զ�� ��"���Q?�0��'�}2M�Z�٤.�F�A���� �����a"�j4nV����!"O�Dxsˁ�CM���p���w�v�c�"O&�3BoԲ�*���9\��b""Ov�p��1��9��O�:��h��"O�����2�X��D�)� �g"O@1i]� I��L�@rn �6�B(�y�C,Swf�Xuk����������yo��p)����?}���ł��y�
��^�fqZE�
&��j�C��yB�R��biPB䑅%��� DЈ�y�ׅ:��@h�����컑-@;�y�lB2__^x11n۟���уG��y�N��L��#�@Ո��&�2�yZ�K1�]=~\�����'��DK�b̋GZ�X�Ag;Zu� �'~�� 1f���@1�E�	~2��
�'R�l��ii����,��ܣ�#MT�<9琽j.T�M�'we.�[&gL�<��1H�b�����h���Y��%T�`˃k�#R�`Q��j������F(D�`�P'ЪM�f���R�e����3D���O��k�R�3�E�Jn�#�j3D��a�j�@��� �h�]X�/D�h��h\+T%aGi��?���q"�+D��8�D�TH�T��3��e1�h/D�h�@�<~/��:c��!�"��ç-D�t3c@�4�+�J�#} 
���f)D�1C��&�PhZwF�-l��Hi"�$D�ba�&Go ԉ�g]�`�"�"D�t"ҥ�)Q�^Q�w�L:F� �K D��CѫH�>���K|� �uo;D�����&s�f!듈'G�l�ل&4D���C��-e�n�a�ǪDD��/D�L[��P*k�Y;֥�U�~� �:D��*�-�B(�ZcY��x� 8D�@[e�0�*�8 f�Wo�X��5D��J�c��`�N=��5a�L���� D�@p���:�pI�Ǖo�8�.2D�j�h�)xX�RQ�	D
ѣ&@:D��;�*̂#	PE�֏O>%�#k9D�0��d sF�!�@���&�$�yPe"D��sE�ʉ?=�=��H
-�����?D�������GN�xKZ �P�UM=D�˳�ȪNʤБ�F�j��LQ�#;D�$�r��2#���W�SmrP��;D�4��"X�WL�$0��.�d́�>D����`F,(������0�P�.D���f��%g�d���+�D|�Ǉ'D�81vK_��6�kE��#D���2D�!Ƅ��1�hPـ�ߨ-3�1��;D��@���G~m9�c��>���z%�9D��2GJ5,���HUH *DP��a�6D�����#*<��U�_`G\)Hp�4D����\�n�
���8%E��7�3D�K��0h���I���9|
ڸ�R/2D���be����+�&����W$0D�p9!��@��Mq�a�fq���F1D��U鍾.c�k���Q4�D���-D�$��JX�#%~0���O�!�<c+D�̱&P� ��y{�o(%M����$)D��cDުi��Ypf����$(D�4Q�dJ�I��0��J\V�X�!D�T��	~��f
�=LM Ei?D��᎛w��l��n�4)��(D�� T��U&G�t��� F����
I�!T�H#����44y��JKB���{�n*R�C䉠%JH|	��W�r�@��׍�`TOD��d�-TT����Up#	a �B&�Ol\�v�\�g�l,j6![�+�"O�m;$��$c���Sr��;a�t
��I6/�>%�G�Ǩkb�P�!����AH�'$D����hP;B���oZ�P[�F"D�d[a�	�`�z1��lL�f���8&  D�T�"�H�X$�K��� ��E��c)�D6�O�������1�^yj�*�(>���+�"O�<a�
,10ū�
����"O� ����sT�����u��H�"OF�*�m ����gi�2JT�Q�"O>M#�,�d B#(��Q�"O�3%�['���C ʜ���pE"O��!�K��b |U��Y�+��Pp�"O8@"���1̀�,Z:󾽁�"OBX16�M6�p	��*әO�L���"OD�A�#�W�!a�h��|��p��"O.Qp�HC2g���C�P�q�Mk�"O�Ց��	=Z^�YQ4A͛�)"O�鉵˂���E��
��j�"@"ON�"���e�"��V*`��\!"OK�#��< ��^<@d�0 ��S6�yr����K�I�"�zd�Vi���y�@�)+�`�r�M6\A
��ŭ�y"��|A0�w�?�
<����y"HQ(R9���Ǧt����	Y��y��^�.ƢyxQDۙv5�	Z�)E��y���+��1Xq�*J=y��3�y���[�u)D�I��+W��y�i�"Mµ��m�FNF��,��ybg
�p}�R�A*$Uӑ��yR"xc���U�zrD12�yB���tx�+�|�D�����yR@������"�O`�云���y2��;6�D�ڒ�X��J�	Q��y"R�U�t��$G�3f���1j���yba��W�L��5 I�t�V���k��y��܍[>�p��<%� �F"R��O��~��h֡n�I+s)_�&v�q#	H�<ɔ�V��9��� b`�B��N�<��OЙfn�&iW�w�=	E�I�<��%Э_eV	����<5(�h(`�B�<A�lC>!��1�8B�(hxw.�}�<q�mԙ�䘱�H�P8���n�<I�Ԃ\&rp8fI�
!Z��l�"O������{G��!�������kR"OPi�TL3(�>��.O� 	�"O�z�!�<<6 hÍ��\��Q6"O�(ԯW�jLe��+T��t��"Op��c�F�Y+��!T�m�W"O^�CBKَG�6��"�pi��!D����GaВ����,LF���c"D����`Рz�ʜ�H߱(���:D�����U��N4��j[�,���fF=D��(pO�M�<9�r�X�
n��I�c?D��d⁳?gF�W3?��8M=D����G���"�l��S�� 
 �9D�����;K7���R(�{��bbC5D�P��L7tkƘ?�,��1f4D��#�b-c-��ʅ��(0�Ћ��3D�dbA�E��#����,D�� ��i�5F�Jܓ��5:�e�B"O8Ũ�)h.�e �Å�3/��)q"Op�� T�p˘=H%DX0A+�ȩ6"O�܉��#U�ģ�H:y,�C�"O� %%�4Y^��Fڮ:[�s�"O��
��-{��X��	-mK��y"O-�$>�l�H�*B�
d��"O¬a�Y�n7h�1)��cZtѫ�"O<��їy � 7�˱"���"O�QHCJC&d��( 7'�F�8�"O��Ʉ�X�$80e��7�Z�҂"O�� �	´Z����e�#���$"OLY����u�L �
����x7"O�ݩW&I5<WJyyG��
���9c"O2=bT��<�n��3��Uxf��2"O��vÖ�b:*4z����om,Yj�"O�Y8���[*�,���E�gE�Qh"O�����B"az���)����""Oex�AAv�R��%IҐЊ�"OrEђ'�s��2��S%:CU"OV�8 �_�I&"��@	o���c$"On�RR%%F�)n��Z��ͫ"OUW��8�4�0vmV�A<�,0F"Ori%^�eZu�WM�~L^U#P"O� 7HҲz���+�&��ͪ�ç"O:�R�*��^�<Pp.O#�HP�"O<��LՐz�X�P�["qTH(�"O�y�삒��u��GZ>Ԛ��"O�(wB6#�h��Tp�1 Q"OL��$�-*��I�UB�()���"OR��A�ԙ
��:�xs0E��y¤�-1t��f�ЪzcvQ�W*ڶ�y��4B���)h�wJp�S����yB��v��x)T��r_�Ļ��K�y��">8�)+�K�2�p�q��ߨ�y�c�)p~�i�D�A�d5�C㋀�y���B�B �T�wp�9�J��y2�__0D��	)l��h�n���y�ݿSu�u�w@{ŸӕG"k�C��%�f�¯N#(`���'|�B�ht҈���$"R�I�(�B�	�B�Q��(o�D� �F,O��C䉗l:X�Y�E���zM�C�ɓM_ڬ ��	v��0h�bC�I'��B��-�Z��)αJ=jC�I<+�����@�:Y<Y��)��Y&FC䉱{(����Q4Ny 85P�v8C䉵P��@̸��"�aN�n�C䉠H;V�{bE��PQ�˘p��B�9qx�e�C��/F%��֊�.p�B�	';�lr��S�s��y��C�`nPB�ɯ2���'�����2'�Y�%N"B�a�\d(�&ìW���ٶ*W�c��C�ɱP����`�tic"Q95��B�	20�$1��*���	1���,��B�	;;��%�P`���qb����`B�*7Q��&^3;A���G��Og���;65C��i�r�i�X�'I�8����?q�4;�nUP��N��eѐk��бS�\�7�`�ĈoP���na�h�'��)[?A�ƞ�Vd@�(
I�K�b�٦��B��$5�R�kB!S���H�jA%%��p��1-`�1���c6��hӈ�.f�l��8��P����*O�4�sӂ��m��9��2ÐL;���O>�$7�O\�᫞�+d�<�c!ϧ[�����nA��?�нi�7�.�$����݊�Xe17�W�^i椱�ލ
v�`���?Ǆ�&2���?1��?A���:��j�ܔ��G�`��0`1�4Q���0T��XjPr�JX�� R@1�U&%|��e#UX���0ǈsI��À#G�f8jy��=8S�S�+W�4�r�8I��I�	��	c�7nx�Qr��	P���ռ���lN��>q�7�ά>�a�(<��1��	CMB�C�k�W?����wP)����7MpR�ꚫe��@���ig6��O��n����?��O����1��o7���0fqh�0%Ӳy'��F�'i"E�(NU�@HTƖ0!��P�D�Y��Z *doH����!z��#�u�3��D�hO�D��^8��p�۴�R����eLN@��O��b�zq+SI`�*��T�4���;/��Yc�bK�qD�
E�G.9�*�gj[ܦ}��By"�'��O2��z�<�{�K�:��|x�I@ AX�����H��ɒg�~QxQ샇<���r.I�2���<oY<��޴�򄆗%�Y���?�������/��`�V��`q���N�W���V��$�I���@�æZ�:���O��$�~�3$�{�ntг�P�+f�H��MIi�'�%8a���|O��ye�ŋ[t\�#��2�!W�B� Qq���B<=bD"�H��=1���ǟ 9�4���'��S�'\vy٧I��@Z١k�7T�� ��?������OlEz���#a�A
�i�4w"^E F�'�"6���n�:��ʄ@�<i�FA{� ^<[��I)~�q�ܴ�?����L݆���O(6m��18�ikF��8C�����"�6� q��,R��R��֦�0�i.�x�Ԇ���%(� h+��Qb�V�2cf	��vӂ���'�\�`�$i�����iæ��f�̭B;j�r�W�X3��P�47����I��M33X���*��!�A+p�r<9Ɉ>(�B���E����`���HO��jE��H4��;�(�n�*����D�OJ�mZ*�M�J>��'�u�n�>v��}UΛ8��c�`�"v�n�d�O�Q3sϐ��d�O�d�O�0���?qشqT����A:��xCT�G, ���'�T�0���b����0<KD�'�D�92j�˶��T��<� �aszd�#Z�F�<T�m�~�� ����Ƭ<Ѵ�p�P�ϝ3�L��%�;q�L<�'~꜉��R��f�=���O����>��Y�f�J�!\<W�p���z?��X�D�xr/�/Pj�2tЅ�u�k�n�n�F�I�?���T���у&    �   >   Ĵ���	��Z��w)D�;G���C���NNT�D��e�2Tx��ƕ	#��4"�V���d�9�o�����4l��AՄ�BF�pMpH��j��YqD"�M���i�J�d�<�6�.�D���HBTt;��(.�&Ts�	\��v�0;Nv��X�(R�(�4;V�5�I�HZe��  삱s�c�g5�2`�B� `6/a�	�,�)� Q����QbR|k'f�E����'s>�!�,h�q*�kb@�"��$%�	�'���ɳϤ���X��P�O h��6)'*?,��*��hcN�Kp�D.yZ�>4��L��8@�>�VΜj����'�T���
j�*}��حIz�P:�'��! �U�h�'���5�J�����<!r ��D�H�#���C�GK;_CJ @��|�I�K�Z@���Oⓗf�Phv���)>M3��H�le���YyƸ 8�R��IuL�)I=��<�t�"���y�ol���h[�u�d��9L�Х����O2E��B�`��'m�ڇD����"��8��8l1`d�k�'!ŀQ��͖-��x��$�Dha7O���JD�zPKa��Ȱ�̋�~m҃J��T�bM�`*t����`�p�G�<���'�Psv,\���1��A�N�T�1�#:a�X(E�M�'���X�"��)M���K>�`F6��ĺ&�I���a�1T� ��ek�m%�DI/7��ika�O�Q̓����n���g
�Q���쌧?�8��>����!Ww�%�L)���!_o<�O�tS�h��Ac��@�
y�t� ������L>�df �&�&��.�!��%02�	ln�qu�F�:�����8!�z݂F��\=dt3GHM�\8�{R�W-`w��/�	w �?ѐ"E�7t&�	�Wl��G@ly2�v(*q�y"j^/a*<$��SFg�����2�+<°��@S45����Q(+��D�?��Y��D����G�Aa�AA��{� �c�N4F~!���@` �  �'�"�'�"!vݡ��4'��PˀឰW�&ոDٯ~�̱�!;j��$*�I�A۴����Ӵ�Æ�x�Ε�M����.ۯE/^ԘG�7�)�'
޴A���B��s0��)��=Z��ЦU"�k��<)�C�)�ܡ�'�t,x�	�My�� �?����?i�џ�C ��/u�T�	�C�+�ry��O �����<�$   �
  �    �   	'  f-  �3  �3   Ĵ���	����Zv��	�(��'@�Ot$(Ғ��6^���qc͕<Cz���'�-�^�����>�\�02ﮨPl �E�r}(�ռWn%�"O�(��jˈe9��r�<h�0�� -��� �☯)�R`C�4~�Pr�HO t�):3�(@��C6�	.1����orR��2̀�)��h�*��� �����T�H���
6�V!� ��VSʁQ0��xh�hУ	��� �'#�~��V��`�ܡâQ�<s"��I��jv�}��ᇞ�?y���?)��Va��O��ဥ�;C?L��"@�`�Y	8c���ޒ#^؅�s���Q_���@Q>�Dx���"�����a��N��"����n�H�S/E�V}���O6q�`P-��#<��Z�}��t�	߹~���*��dy�����?���?��bޟ�)�OT�LP֭�,�C��L�O��+p�)S�|Q���D�~���,[��AɊ�4�~�Ŀ<y��ܱP�X��'��QFlʡ`�H�n�Y�c���?����?	��w��.�O6�do>y�ր�a�E+Ti���eaѿ�B���N��v �i�uʘ�mz����Cq�2#/�4R�(�!�;g��D�Q�+G��H �+/�,�'*�X��d�$J�Ŕ�<���C�Z j�����iٶ6�,�I��H���Kܹz��jP%,Y�������<э򄒍��;��c����v��
��	��d�<y�CX%_�������C���ǠI
dk��u�� r�m����۟���$�n�r/ċ'�~ �w�vT���O����^%�%Y��DAx"銎�D����悅�l&��3Ч��r�z�q��v�R-�'A��ʱad�?-r5���^�_N>1�I���}��\ 4Ě}�c�*e¥��m�C}��'�|�L�&,�4A���5b�`ܓ��
:��>AМ�,�&�^%VFbMp.��$ ���O�>1�f�2��V�'��T>�:V�ʟ��� {���JV�1����$�֪�P���48�S�@X�+��#�"?�����R?��|�	T3f�����>��� ���?�$Ƈ�^ 1р��3Ρ��+�h��Ey�D�#)�(p#犎�%1 #�g�O
5���'f�����H�į���cK	.��ѵf�	zz�Q���0D�D��D�0��%�fά4��pД�!�	��X���4���(aU6(JfTr#�
�S�XI�$�S��%�	Ɵآҫ�V�^M���L���К^w�2+�0ЀQ� K>R��5���է�*H
�)4�:m��ꘃxg��JcO�|�ߴo��|&�l�c���'b���
�4�\��$G/&P�1�X��Es�k�
Uz�'����iȾ�9�4Ot-���>V�؄nظ)��I��S�DA�B�O6�d�OH�x��d�I0�������ǥKߦ݄�v�4H����n�S�Y�D��t	U�i�"=�'�?�)O y�ã�.h�pa��mƹ;-9��.ZgLF`����O���O���ɺ���?y�O~Z������k����P�R�Gϲ���㔋cEFD�3�M):�U�j��]P�6���(O��hV�̀B�d�d��X n���Ĭ>���b�\>K&x0�K7jߔ6m܇'0�E�?�������!k��LR���Y�G~n)9���M�����'n�>7͜�P��h32h�:9s��b�(Yn!�d�0bX��@���lP⨑ց�gx����M������;>tĨ�O�ޟ�Ԣ�/Qj"���[5S	�t`�i �C��'yb�'j�8v��"����c�@�z��$H1Ga>�:��_>lF1��JR��a۱�*ړ�jT�T�ˀb�l��P;A�����Op�zA Լs�Y��A��tU*]9��̜A���'�q��5�ǎ�J��*�uC��K�l�>	��p>Y� �M*�cт��O9J�%h�dX�h��O�T�'�P�F�X<k��~P��bV�l#ҍ��M����?9.���� �O��䒐oL�QDנ@+���l�	�Hhm�)dT{�n��E�8�������\���c>��F�S�3n��J�$J5i�����П�#�!��m|̒'��z Z��_�?I�"�)S�BȔO�te��[*"�u�RA�:X�E���'f��*���?��O�O���Oj`�	F�7n8Qt/	C�ވ�"O��Sk^4/1����o�����D�O�Ez�Ob�R'/¶3d\�S-87y~����|�*���O��'�GY�D�O��d�O���;�?yԤ)V�I:�Δ��mP#EY�x����C�9c֊)��]�4ԕ��\>�nZJ�vOj�Y�Pc�A �OS�x�R(�pn�6�t�E��m�2�+��>��̦��d�u��T�,1a��v�6�0_�6�̕'eޱ���?�����'��	�+B����@xB�ŧG�~!���83 N�uY$;e���f�v�"��|:���	TR���q�AN}�Q����!���h4��^�<��)P�}���7�Ě�H�D�Y�<1ÊF�1+�h���L���*�Uo�<��̗jV���0Ӊ/h�)���B�<	��*;��"�̪S�ڜq�Cz�<����pQ�)( �$F�@aI�l�<�F
D�&uԐq��7g��5Ys�f�<�`�+Cy��P��Z��4��`�<� 8)� �+*��1q�#X�`�� p"O�xx�	�!J8(%a|��$"�"O���U͗�3A�IB��2 �@U`�"O�m�@��*GҀX���y{�"OB9c�>+�d<b�*�-i��1�"O�D�3�G�S�<�G�G<`�I��"Oq#!
=&H0���iQ�c�����"O�9h�L"��pi�O^>���(�"O����J��ѵ�U�(8��AT�<�E�R�AqR�0�Z�p�h�f+�W�<��һ��I�(U� ���;��U�<����-�H��ڝ'�t0��	P�<a�`�$7=T�:�|�5k�o�<���G���`�I%#1C2��E�<qу�ȴ�굫 g�`�0�`�F�<y�Ǔ�Ja�<ڥ���t�	�o/D���9B`�!d��f�Bq��i-D��!��Ջgچ�����<�NdzcL(D�,8��F@DeT�A?�@q�)D�D���Ŝm�Z�zs�N9gy
�QGC(D��(@
S"1���S̀N�`��6D����jc@���,�OT��*�/5D������%>3 YڢK��bXA!�$Y�1�-��o׮\`�J��0!�$V�v�h���b���AB!��P+6��-�#�)#bU�/��oX!�d�?U�Py���L"m��A Y6vk!�P;>�,h��͍�%�S�E��1L!�ϣ8�$�#�Q�k	��[�!��C+$Q��N5lK�,����7�!��َ�S�!]D(|�@퀢T�!�Ć�v�"��`[
%DXE�4M
,e�!�d�0�5:�dY�F�lQ�V3"Y!�䟧>��˴C�'�de���$ga!�䏐,�B�b�.Ǚ,�y�-.\�!��W�������7!Z������ !�ӄ9�tX��
æ�Jd���fm!��t�`��H��Y"I�>0Q!�D�kZ�lH(؅zʒ�:��ңO�!��6b�98co�c�H��m��$�!��\.R�<A�����c�q�!��є'�8�KҨ��
=�}(B��>!�ƀ(�}�e�%1.|U��W*!��R�Kp�Ɓ�2~�5``G4)!�$W�z̀�Wm;DȈ�Jsf ]�!�  C����!+��y,R��#���!�DX)qX���`N,X�QC���!��P̰�+�7xm�����E�ȓs<:�#GnIq>�uq2e@
06�G��UD������!i���R���u�u�ҋ+�T�R��6$TLX�"O�������P���C[�<9l(HP�5��=b��0���i�7�Ѣ�F&/s��h��܂]!�ɀ	�������:��C��X�&��z�Z7�I�X(>�� <��Ub/Zɂ�,��T��7Iٍe��"	]BoQRG
~�j�@(P��.i��	5U��P�e�4����D�;& |�����L�q@팍)�џ�I�"�h33�	�v&���Ir���h�=:��u	&�\���&�HpU�R�q�X�@��3��T�'�F)b�K
�RL`�Q��� Rܣ}J%�Q�1�6�1�	>B%�AϙO�<)!/U�9g�E�T��*;�H��'L�2����q"S��M[g�\��I~�=�F��&9>�mP��ǿg<҅j��FC��4�D�ƶ0.q2Y	,�D��n%d���	A���pJ�9��=YQ+�f"١�2��1��Z�'O蘈`��S(HT����$O+���_3_l��p��M�#K���`cз)�!�� ���7oێG���#�����2%Y� У�
2�Z�Ϝ4
�`�ڌ�	�4/���
�,~���%J�x�!��8$��z�'��,<ș F�Q7� �B��Ҿg?�6�)3��4뤥3��D͜5f�p��pTd���)5�RGŌ�}���cEӠm��AɘA���R�+��d�	;��=�c�
3.ɐ�l�8J[��8Ul�Q�'\�̹&G�9��m8��\�!l���]w��j�����I�l�!�DX�b��Jt�S���,��"�e��!o�� r������T�5�h�>�0`��4\;�b>���6"Ox��j� e?�Slն1T$�����Q�'p��۔+��D����qO,u#7�	H�����6?�(��!�'�u!3�X134�p�G!+��ء�/ơӈQ4K������$|OjMyҭ��p.��"���b� ��I�.r¸�C��.pຸ������*��d��XQU��':,P��v�<Iq�K�Ra���x�̸h3�Jq}��/w��qa�U�9�
����u�O}�;@m��hؠ]���Yx�D	�'�X�a�a��a��܃�LǳdbPp1���yyr�]O��C��$��DŚ(�K�斅@��۱�ʭk�~r�$U�ڱ V�p5&>V��1DT�]���cQGS��@@��F)��x1�[�4�Mq�M>�H���*����W�&}I�֗����p��q`*�X��-�!���-7�$��H
 �vY3䬂�3�����RR�Ê'�\��g�Si�B�pA/��	2F�ZԊ��o2C��%
g�QaJ�������m��\�tNo��n[r��~&�B3J�\��93���*&�@��5��!�O�t�Lؑ�D�L��M�B�(r���K�ǔ=	�N��dѿ�
̙Gd��o,�;ՌZ�{�axRh�b$}�d�̉&T��M�Q&_:�� �0C�d�ȓ^�=b�MJ�{Ǟ�AFo��I��'m�y�	�%�F%���7���R��t�]=g��DyT��0d
Fi:w"Op1��FL�>�8����;,���R�9��u��'Z��F)��lU�ϸ'dXd�'\�ht�K�<L"�-h
��E�ȱ�"�IA� ���Ě��N�4G ��, `�Ib�y� YpPM��u^бp�ɒ�.��,Gb�QA
�yC�ʙ���Q�4�:Q2���B5�gjEw"O��y��/ؤ�#�f]�x-Z1�>Cfݚz�>�X�j�z���2�'&i�@���	���C=T���6��0�5�ʁuz��� �U,P�b��#c�Z��	�b��*���ē&���B�'���R' *"0���Q�<�F+<K�f�a�+��pPf�C�!4����gV�Y�J���*�fE�e�9L��+#�*+%�@��o�)+�
k��A��eF=pα�'*��FW$Eq���+yl��6��(�ԣ�&_�^|B�M�S,�&�|@�E��,�`gE����lD���]�"G��E�^I�D���yb�$1&�z ���qK���'�ݕZ�@`Ik�G����:��\���L���C�}�� ��ڣ=��d��%D�|x�m_� 96��o
+���baçw^���k�z�a��'�2�`�*�lbfavY"(�>U�
ד��A� ����ܴP&*���d����V֑ �ņ�"� ��M�ZP��R'٪]L�5�=��d�fo���H����e!��t�#I��0�`�hT"O�FNO�>������4X�t��P��/d�%8��+}��$�g}R�$s�̹!P"��nn���H��yR��_�r@��v�F=IG@��y2I Gd���ɵK^,�� F�'�a�HX�c���C !���l�R�Km�g���hėOS���ȓ��(qq#͂L
7o�A �؇�W��|�ub\o��%zu�$ކ�ȓR�P�!��V0h�#Q�Kt ���.��UX A� ��d ca�=N��݄ȓd��y�lՏ(G���
�v����ȓ ���KwƋʸ)�PC�o�t�ȓ|���f��������X�d�ȓu"0�I#D�*/�رѧ��D�=��S�? Z�� e�yF��Sf逅"O ��/�t�@����}Y�<��"O���������pe�V�lFQ�"O�%(� 6�6�0��V,LQ"Od�"I[���ږ���d�`��!"OXtj`��	S�<��M��"E"O�����mo�U2�	ں����"O����l�`�����5#I2�#"ORY�rbӑ?K$�1+Zp@Zd�!"O�}��B[ Wd��9�X�S�*Ä"O��q6�Q>W%ؼ�7�\7A1���"O�]����oVU:���1T!�x�b"O�@:��*.�ᲁّQ��Lx�"O��{���!%q�e�.?�a2�"O��y�-����K���0>��I�"O �S���<�L\m�y#n��"O~QO[�UQ�,y�㎌��`BG"O��3ЉD���K�ɟ�_���Q"O���'aD%_���N�`��;�"OtZq�P� H	2�J�>9�5(�"O@���ú�U1���1 ��b�"O��Qˋ�l��2"��<�f��4"O<�h�,N+W����(W�`��xb"O~��s)�4\�4K@ƍ9)�B���"O4��� B��rb &9r�A�"O�<b�a_��M�p �WB+0�y�h9d�rXE U�q_�1ztH˫�y�
��;V�:�OCi)|�ӧC��y���<�C���O�1�GHˎ�y ԒA�*�˱K�#�`��ڱ�yb̕�D �)��J�*�^��eQ��yb�O;v��m�#��(F����+�y��)>$��`�B0]R,H��m#�PyR Y�f}pESAs
8`kgk�P�<a�AR4W"��0�N�I-"���u�<9��F��� b í�:��A#�e�<i&`�8^�!�hM�`�����-�h�<���Ӷ8�9�pi�����d���y�.؜/��nN!ɺL�wh��ybӎ�"Q)�f�=�<P����y
�;�=�S/ %�,��X��y� �	O�FL鰫�9��KW�)�ybb��z\{pB��>�1g�y�g��{-i�銱	L��I՘�y�ؚU3`Y����-����V�֮�y��ߘg��LzՈQ�,��)p�! ��yR)�FǞT�#&\R���$Z��yB@{�mY�Ƒ"M���B�.�y#��J�A��0�h�""0�yB�ުSC�!Y$b�:a�5�V��y�lX�"�T��IR T2�y�a�9�y"e�d�
0c���2-��Y�f����y"aU'W��Mj��T����\>�y��S-��z�(�7S&$dZR��yR��"*��	;P�J�KYdm�U,��y���z�q��K�B���!ND�yR�̢}�U
�dڽs$�� ����y�.��L�|��Q���<����ؓ�y�La��̘%-:�5Y�b��y��=E�j���o�*�蕘ٌ��?����!Z��9'��q�h��y���"O�2�I� H��:/ֽ:����u"O((jV�ȧ�p���گyY�'�$I3�mʓ#�@�ɓ
������ 0� T��?5��x'e���E3C"Op��+�2<z���gdF�'\�}�"O�|y��O�,�
	���W�iI�h��"O25��` 11�2��4���)&�x6"O6�++ݶމ�%oŏ�,%��"O��r�BM?4�V�"`�%$���"Oʐ8�ǎ�YkC��2�$�D"O��[���3pJ�]�@�x�"O4б�,ƦT%0�R����:E!�"O��h��3!��.
n�>�"�"O��xB�׶ؐ�ԄƷ�J��"O�iR�m�=#�D�@逊�z�K�"O�L��ٹ1�Уb�F��H|�"O������N])S��4����"OT�W$U��4�ǯ5	�� 23"O
�Y���fh�@��AA!�@�5"O��!���%�R�3�яH*�ى�"O���$
�)�fу����&�8�"Ot�"��,PL� �D�&J���"O��c���3��9B����$"�"O�u1�=K=~Ase+ۢw���A�"Ox���I=~��]2�
���VՙV"OD���[5;)�e�0)�@Є��"O���D�	O��q���90�2�"O�A7(I>V�ݳ��K�*2���"O�i)󀏡y$��;��3DEn)�"O�UrG��J��W�U�`D�5��"O�mS�0>G]����^C|L`"Of�h���9$��)�M�?"����"O��RDdG�5v���!̩��ElE�<�/����-8��/x9ntv�~�<�C��\Y�&�ǡXY��j�m�x�<�S�OR�	����6^BE:'�r�<��"]�9�Z�(a��92mBr�Mc�<��!5Bd�7�ҳ,kr\:R��d�<�E`C�S�<��$��bS�ia���E�<1��)��쨅���T}�&�|�<#�^��m���]�`I�l@t�<A�A�����������d	lAd�<��H�q.�!�F�7��I���`�<���z圜:t���M��(��Nf�<٢�Z&x�!��;o��a5'�v�<��_�l��Qq��:�:Q�dx�<a��DB�|=C�C�=����֬i�<AD�2
�B��󏍍�t�a�kg�<q b�0v�J�PW��!3���H�<ٗ�ݺn���!��>Jܔ)���O�<� hF.H�ɨ ��:n���S"Dc�<�OQd((I��7nR��v��\�<!'�K�Zb�t@��U�,�U��IZq�<�p�QI��%[dI*72�r���m�<��.L�1��V��B�j)f&S�<�2B�hT8����CX�	QH�K�<��싲(�Z���22�%`��q�<�7'7��0�3g�*N��+� �k�<�u曔g�V� W#ZH�DP�<�!N�1]� !R�RQ��I�ciY`�<�&o�y��kc��	�f0��(�^�<as��}�QKU��R�� �F�<	�#�$�*�&������@k�<1�K@�V.��h��t7���P�<� K_+w
<8c������O�K�<y�J?*梤�&
�}�X�і��M�<��N��a��@٠"ʖh�F�)1H�<� 2*�+G�P���3d"�0j�Q"O@y��f[,[f|m`��X
s��[U"O�0
PBtư�� ��7p�Xj�"O��x#�/�~)*���5e&0�E"O~�@�J�nQ�yJ� �.4�{�"O�b����V\�I�/�4~���Q"O��)P��<I��	6NV.Рak "O8�(�Ő
?9М��쇐���J3"O�}	��E�1�|*�K<ΜD(�4O�d��I�A� E�w)W�B7��ȳ(�>^d���4��$3��D���1~�x�o�8i�0B�	8K!(aaR(�;�����P��"<I�)ʴ�E�9v�b���6~,��quC^q�<�q��!H5*�Y�H�2M��p�qF<tQ��F��'�H|Z��՛**&ً���)��q1�'�xy�t+��G[:��G��6���'@�1 �b�2tx-��aȇ\bdj
㓡��pqH�h
p��q�j�R�P݄�^$L"�Hϱ
�.�Q-߬y�ȓ�L���o�&�S&숍�ȓ{.�IW�H_����F�"?l\�ȓm��$ɦ.W��✂�G`��ɇȓ(��S�Г T������� x�ȓ9Z�%Ό���5Y��"Q�ȓ���l��
���p��;|��ȓq��X��/�}�(pp���5���ȓd���
c��J� ��~q:��ȓ3��8c,C�h�C��=����J��q�D�iw�L�
'�����>A`�"�xվ]#��(��L��<8JXb�H]-�$�@�	�e,x��ȓ;��e#B���!�bhZ����T���ȓz�x\�E���"���� ��<Rj���i�pÕ߸f��#�[�_& ��K_|�S�녙�b��fЈ�
�ȓR`lC��L�4��p�qi�N���ȓN1^"��<0E��9��	�%I�܆ȓ���فi�-LV�I�W1i�ȓ.���K���3y��gǱ<.��ȓV�vy �
HIv �凑0=�đ�ȓ�D��r��\���CA�<�,Ԇ��\i�J�;��c`�B�!A�I�ȓK"X ecM�8�Q{�(��(���<��	VmE�Q0���	[����/���p-�!uG�#��f\�L�ȓ~wF�r��ȧ]U��c򊆙Z�ր�ȓ3��m;���H�:M[�,��1��Ȇ�	��,�elK���ͺB(��ȓ/A�����:?��+ףg�F{��'[���lMӈ�	Q��GC`�'yР��O\�b+�$P��K1Eg���'�yѲkX1z� !���09��D;�'�m����J�\�r�,֭4�:�j�'���OT6�*G�9���i�'��m:��D�P���D ؎7*�$��'b�$2�G	�
@�a8$�>`�0�'.(�#�_��Z��'^���3
�'�Q�T!/Xq*��.ЃV�ָ�	�'� 0[�/=G�Rlც��I 	�'-��1�<3ޭ���ɬ?���1�'�Jx��(�H�L�I�M�����'�
�U�ȁKMj��r-Σ|Ҿt��'0ِ´xzi��I)n_~(��'� �Q��:\��eɄ�TM ,y��� p��k� Φ0�$�$��P"OP��$,yRjXx6�!�`y�4"O���b-(�*`
ee�5d����"O����C+��4)t�Q�v��`��"O~�궤֦-6.�;3��m��q�'"O���� ��IH������"Oڕ�V Ю`� ��΅�r�,(�"O�ԱɄD�$�$�Z��@93"O2��*��P�t���_̈́I��"O�r�k'\�� O��5�|q��"O�$ᐄ:D�=�/a�BV"OԼacn�yt@��L����@v"O�x"d��A�zL��OI���"O�90E�]1yP�1��KP�{㈉�F"O�DZt�_w��j�H�^�||�6"O��P�K I5X%@t��[�.غ "Ov�eېpU�}��&4���"O>��%�^\�(Ip*�L�`���"O�8�q��w����j�/��@�"O�p��d �ة��hƑ<���F"O�0 񫝋A��QcUQ"�Pj�"Oȁ�EF�B]�9�֠�`���"O&(�cf�!�P���JA8��"O����*k#����3��y�"O��;�.!%���Q��Ò.�j�@�"OL�I��%iy��s�嘈[���"O�q��w�6JS�M�D���RQ"O�(z"�5t7���6	F�?���:%"OΑ�
��A��xuI"�l���"O��HK\?&�������e�a"O�q�=����%EZ:#q�QJb"O&�آ&N	Y%r��e�V(@Wv�B�"ODC �E+2�ؚA��5a�x�"O~���cF-[�1���3@�!2"O�٢�g���x����G�$�r�'�ڡ҅�ٶH:� ��^����G%D��ː�"	�B�k偕��i 4##D�4�!Nݷ�T�!_�uB֑(�b"D���E�Ԥ&�@���k�94E�5��>D��aRd� ����B�,�xŒ�>D���6�<e�\�B��T����fL;D��"4B�,|,xb a�ziSfg7D�D�𡗼g��up0�5��
u/6D��� �Q?U����"��1ۅ)4D�4P�)��IL �0({n�{wg1D�$�j�1�r�2���:zP�`B�1D���������5"�O�0�{��:D��ɰI�Z���U.Ȇ#�P�#*O�	;&Q;�1��ܮdN�R�"OH�q�S�w�T�d�/
R�Q�f"O��"$ 9�v,���$���`"O(�)�h68F%hD����x""O��j���_� ��N����c�"OL�%F
-mS���M6�R$��"Oty�^VҜ �vL�,jJ,k"O,��t�ۤQ�:�q��^ DpLJ�"O*DS��W�-ňt*��ґ1O.��"O�y!%�?/ch(�� �-V0.���"O�e�Ћ��9n ȧ���,��!�"O�Tڧl�yV�s�؊�^�
�"O��
7˂y�ux��'f�^��5"O�x�o#<u����(��L_`ܓ"OVe�t ��P]p � �j��)��"O�x�`���I�Ьx�FJ���ir"O��-� :     ;   Ĵ���	��Z�wE�?]���C���NNT�D��e�2Tx��ƕ	#��4"�V���d���o	��9Q�?=�xP�FL�P�]��_;(�`��H�M��3!�.	L��	w$�	zZ���B�&��4eۀ�f,�g� "��k�i�f�h`]�X���$��N����ӄ^��D2���v��0`�%+ Q�N�l
�	�""�t%"���>�\Q�UhX��'��Ak�dڔ2 ���֊=���톎+~�I��'=p扤P���	�]�$2�OVҍ����������<���s���s�>�@!C9 �ԝ�ג>a�'έH��"�'���*�e�,�@��DW�s@j)@�'
�p&Y+k���'�Bu�ѩF��t��G�<���Q�5�>Ԡ�/֓�B0Z�hz&�1���M��?+�(�9�'�A⓫_�0�����!{g�'̈:d�nI��ڬ]���U�(Aŀ��E�mjDH�<q6����2v*v��d�Z�OH��¦�"$Af����O.3E"�8 <�'���x$$<��I��D) (�~�MC��fH�Z�D	��	�y�Rm�)ot�L�9O�l ��"o�\��l�2�(��zJ�!ň���l���g���z��d8M�A�<���'��)P��G���	P�e�����<*�h5�H@J00��۠[�:�\t�冚G�N%*H>��'_�VKi��a�;d��ܹ��\u{Tu�0%:��A�Bzy۠�O�4��ıI�踟0A���(v��u�<�(�	X)�ɊS��G�2��N8{Uǐ|B��	<����ڟ]�aCc.x��{��j�ɪx����A�9�d��;|���a(�(��a"�Oٹz�P+���9i����$����658�6�RV:\ Ա��ih��OY�ߴ\:T�{w#�]ȵR��v{~�'B����j�?1c�'"���l�3(�����O�/�<�Z ��:a���gg��!�ʒO�`��1O�9����gP�����];"���Bi��)�C�PjN �  ��?����"O�D:A��<W0=�"��JP��`"O,�����#���q2l��3�����"O­�t��C�Y��/]yBT�"O*��Q�.N�*���@�$̶4Z�"On͐�EՓ/��r#�Z�^���"O�y��F�8�Y����.	�ژ#"OF�ss�H�d5[U��O}��"O�\8��V�Y�w�i]��6"Of��f��O�*h`�
pGZ����	��HO�Ӎy4I��ܲ[��I�\�N&xB�Ik�)0CI��p���1^�=I� W���d[�|�݈����O���n�X�C�k�0Ԝ)�ԎA,qE�\�v�a��ʉv3���ģ����H�RN1��=9l �=.��#iR�D��ӷÖ;t�!��G�F��H�#�&����σ0Zh!���(�:�JQ*֣'�tv`ڷK!�D§?I�m�T��*ab�q��F̞�=E��'����͝�f��mڠ+��M�'h��aC���k���w%����'&�9(QF�G����� ̤n�&Q��'��1���cJ�5� -�)f�r��'���QS撋{R�c�,���%�	�'�LԺ��ͺ�T9�-Y��5S�'L�P�J?T���cI�O����'�d��&���Z����eD�Y�]�'@��֨�RPzH��P#J�M1�'s5��B+u���1G/J�xeR�����ea�b3A�0�S�8D��.<P������Z�h�2đ�J�\-�ȓ5T̑��M��Q�����S�.���%V�a#�G�U�A���U�`�b���,������l
t�N�</4=��p:@�І�V��PF�5x,�H�ȓZ��H2��Su|��ӧ}㜬��J��kP�ن|�����Y�?� ��ȓn�<���ܧ?�Eq�.�d�<�ȓ/Q:���� 2���X �Ыp�T���S��A�C:*�a�'�O=a�b��ȓֆt��gK��� ��l�F\��?��)���H ���aO$�����\���@R�5��s�?($h�ȓL�J% ��[�k��1�7k�ن�S�? ��QD�_&6�t��5oĬZ:v���DKQ����3�l$���I;ĭm���R9l�C�	0�V\Zb �Qx<x�C�	;�Q��D�`���䏱"H��2�1/~LC&�sm!�2�R j'��S�� ����*^z���).�O�@��ʝ�A8��!�BZ�M`��'������՟]�vL"'A��~�$�#GE��t)!��D�@S�Jsퟨ.\ 	I+R�W�O��b��)�)�����rV#�I�t�ӱ ?o!�A����h�V��ږo\m���=E��'�8�A�*�p����f%�,�D��'7�p;r��(����6cI!#�0���'�R@zaR%�`��@�Os�<9R��5@�x
���.�>��0Ύo�<)5�JHDb�aG�<b�"�j�[o�p���<%>]�6K¡wƨH�n���+%+��yboB�y��!��Zs͢�il�Q��@��Y�4���p�0-�A��~��ˢ�2D���$���1or�b�T�5\X��#k�b�����~��6fY^�V�
�T�'\��#~H9�A�P#���u�ȾWtV��ȓ�x�C�璦
D�1ڤ�77x�y�ȓ�\��"�hD�!$�0
d��e���� ��	��H�K���t���\t���H��=w��a��6=���E�T�96��X*��D��=ƴ��ȓ�J��ϐ�S��R�� 2Ld��1"�3a��9p�(|��ʧj ��ȓ*��|
4MԬD���a���h��ȓ W��`ƍ�w�`E���h���ȓ!�|����G=~�8�gݢ.b����ar���#�n�����W�+r0�ȓq�<��!T�HA��n��P�ȓ0�6�� I��-إ�Δ`pA�ȓY�1@���Bw�!��o^�Ѕ�b����LV�\��a�K�tZ���Qg^��Qh�U�><Cg(M6a�ԅ�	��"g�%�p�R�l�6L� ؄�V�pK��@���5{Ǿ<�ȓ~mX`�4G�Rb��Aֳi�H���37�]�'no$�ʵ,�*�����&������R(iV����@k>l�� �Zݓ��^1?�6Ī�G�l����N��XT�D�*����H�8�ȓG���b &@���0���(�A�ȓJ,Y����D\16�Tk�<��ȓN��J�e*I��1����@����Ic��͔Up�@�T]��P�ȓE��d�b�\#��a�g�t4�ȓj�������Y�Й( �p����>�d�[�Ĺ}��@t�цd;���ȓS7��)
�dat�9Q�
����t��h��F�m�f	'�F)���ȓ6H&��weU�}Ø�Q��6Yzֈ�ȓ1����	C�(�D�Yj:����]�!bF�'v��0ȕg�J �ȓ ��F)@
H�H!�@�6 ����ȓE��J��8|��Xq�^�I欜�ȓ'��"�)!b�X��Ҹb(��D q4��! �b��N�Z��݅�d��]3�oA{c)`�'>c݈���Au��4	��jҎEz M}LΩ�ȓ �Ls�M+�����9q�0I��O�pyz�mΝVKhp���@����S�? �*���-Ք�ϊ:8����"OHڰH�6C����n�T ���"O68��=c�K��U�z!���Z�<����2� �{�`�00����Z�<գ
��L�F�.!e��!KQ�<!UE�].v<�E O� u!��ZL�<�d�=XJ��T�Ēy�^y�*�J�<��VP.�*�&��q
�<�R�D�<Y $K��[p���0�1$�I�<� T���� �`[�6Z4٢oM�<���5[�+Չ�<5A4-Q�M�L�<9Fa�7m尀���ѯ1%��2b`�G�<!Ă#Ɉ��0Ȁ��ڑ�Hi�ȓ�B�B���]��
�IҐ�~%��/T�K�	�:aӎ����M�m^ i��{�x���GS.A�nx�u��o�(	�ȓC��� ���x�R�Ifp����&�ť�u�`�p�ă��X��9}��ʅ �L�T��� �?
����ȓ9�Zϊ�vdV\��� �f�<��]�=Lh9�f C7|#G��f�<A�K��
|y*��Cdx�s���`�<���,   �      Ĵ���	��Z|�wI�:.���C���NNT�D��e�2Tx��ƕ	#��4"�V���d�;!��m#7���7���r�p���֖$Ԓ� ��!Z%�Y�I��M�b$0$���*�۔cD`�V��ȟ�i���?l ����*N�a�`��;pzU��yCf��G����I��r�J\����c_��TEL�b��Ga@�*�剁�%;����04 �g-]�=N���'8����J ���w.*>$��[�Qi4�x�+mb֘��
o�\����d�f�@�oN?]�T�U�s��/"Ā�g *���r�;E�O��c��<�hPs��5�D]�E�O��/^���H
-}#ś@�҅sK>Y����R�!�u����38�(�q3�IB�'=Ne�Z7&��O�M��!F�=H2p!�� T#�)|��L
u�x�V��ZIYL>ɒ*��Z)�p2����S��
hr���������;O�����¡��.�q��f�	#U��\#�D\&"~�y��J�n�P�I�ñlS�'��\x���6��'D�˃K��E���
+"��4���ga(?�m
�6/��%���竄=66�'EJ��^|F|�w�ǣx���Qd���A)-O�d�I٢�ڗ�7�L~�� ��A�=3��cʝ�	��1���6��|�D5���Rp?�"4O��`��ە�~�һ!~��Do^�L���������\�$��|��C��D�N>I%(�T$����^T�P�
�O�:o���Ń+��B�}ߊ�E�D�3٪����N.6�P0����8Ζ��Q�kG���H�!h�t��sM99��� ��O�R��8;���2��?�v��51v���c$�(K�q rM�my�Aޕ	�\LQN>�։»5�l,%����K&p�|0ʗ�U�E(t1sgU-Xh�x�w�$��A9"8C��d�>i|DA��@M�+�GP'��Å�1D�0TF   �'�F�@ ��-ޭ7J���_7:q�C�I!U� �  �;  �  � �5 �A�5{H�,�'���谭+.�t��4��*I�`�
�'�8e@�柱����4MA8n� �'D�1ӵ�2f.~|����a<l�I�'��Ax��ƔjJd
uɁ4Xi��)�'�,�1e�@�<xT#Q �SfD�@�'��D�qlZ\�ȍ��jX#NJ5�'�m���H�k�R%�Ə�"I��+�'W�	ȐJ��>1����"I�3�����'�8E��d��.�Z-A��V�&����'�@�0�K6DtC�"J*I��'�+l"��z��R���Q�W9�yCI�4�S&�ݾ!�mM��ybh�$_�ҡۂ͘<G�d(��G��y�e�*��aP��7;8��р:�ybA���#��%w��D�A��
�y���~a��� C�u6г!��?�y���P0D��$�~�� �1�y
� 0HSb!V��X\�iJ��e��'6�O�u� ,Z#�Y�n��5�"O�e(㡐:Xjj	Y�M+������=�S�)�*
	�XE�$p��Yt�̫{�!��Z�Aa>9A�Y�.l
1�q��(f}Dz��9O,Z3���Be+��� ,���S"O��0�T8h.����r�$ȩe�'�@���	�al�z�����#T[�I2�C�ɉ(�8��c�'74�(���3��C�	>@'����T4�$�k`�]�/�"<���?�8CE�D���\M�z]�Ш9D� �� ��00ɢ$�
pe2���7D� �@��d`�&˚	6/�:�c5D��
��u*^@�䮍�@l�}�vB4D�`C�d�i���V%�1X�z�ip�0D��{�i;~@��@M*U��2�.-D����Y�aP2��f#��Cf�(D���V��L��
�GK����T�:D�c�-Ji*��1A�`�/8D�\�bΞfc$�p@�-a{�� 8D�|�w�҂r��Au)D�QhF�!)6D��T
��2<0��q�O�����'D�|�tʡwa����n�Dp�#&D���+�6-K4�EO왑�G!D��	Tꄕ6O��!�V�cq�y( ?D����Dg�: �:4�Y9� D�P@�A=j@�@*��0Q�`�E>D��x���w� ��� p6���E=D�{ @)?�2Ĺ�
ĸw�v�j�d D��q!�%*<0P��'4&t1�4�?D�xz��x�2iO#^�l9P3�'D�Q���'�(`	tm3��k��9D�l���ĖN�J�`�Z�z���QJ5D���V�q��A�̐*��Y�#2D�T:������q�J�ܹ���-D�,��8P��g�Τl�����J.D���*��5� ���8^d�HI!O6D�����N51�zm�c�K$4X<b��8�I�9��"<%>�Aذ^��Q��BN�P�����8D��RHđ=� p��	�.T���Z�@}�'�D�,OBx�u�C�[��r @W�X�8v"O�ܪ�Y/@�œ�l��v��5������I�
µ�%�OV�rmb�eB���S.s@�'���r�GK�5 �L��B�3�y"/�"2U^�J�EO�� ]����O��=�O��x��>S�L(��4��U��'t�+���S������8 ��J�'D|��$ $$�}��dM%fPX 	�'���� W/��8k��:p(`��'�����+Ni�%۲58�h	ۓU�H�OfP�7	P?;#�D�2���Ei*���"O���ӥ��"��A�E�� M�-ڧ�DH�(O�O <`s��P+�)Q-D� �`��	�'��eX"MQ'��U��� n&Ɲz��	��H��	�i���d��3`�j(���7�B�ID���I��d�B�b �Q�DC�!{����똰N�F|�g��!*�hB�8W��0Au�>�
��H�e�JB�ɴbŀ�'�%=$I��·!�:B�ɦ|.�٩��%�ڄ�c��Jn(B�6��ɸWE�O��!t��>!�4B�	C�J0�̩]� 83�(h*B�I��(x�n�W�88�&��b��C�	]\�h�U�I���N,K��B�)� tɃgÙ��[nZ�hk�p�R"O UȺ7�~ �d-�'?D0�0�"O����#��(�n�J/�$��"O�`� �O�\2i��@�X !p "O֬�C"�vK&��eM��Of�I�7"O���j��8ZpK�%��F����"O�i��m�:{�8�u.\���y�"OJ�G 8�PT�C^���y+�"O�U�V"	;m|�ЦKG��D�y�"O�J�Ҷo�H�vL�r���Y5"Oԅ2�Iok����[�lE@4IW"O>tK5�R�8٤R>p?�Y3�"O|qq���"�^�c3��I5M�c"O�1��Q9�,2p��Q/l��F"O��q�L$8�tc�*E9a�0�Q"O2��$�@� n� U���<icQ"O�)���F[����Mƚ=0"O�%iԋ@ ������C@�4�K"O�|�V�ϛ>�&+����N�2�j�"O�a4��n)��Ț#☘�`"O�=zt��z�v �AF�3.��1�"O2�i�&��
e���]2`&��r""O�a�1�թ=��$��ht08�"O<̈����n2+CE�c4b0���J�<����&}&X�N��mJ���)E�<9�ȕpe��q̐Bi�d��MY{�<���S-��e��ɚ.e��b���z�<1��+{L�Q���̊g���P�_y�<A��Ѩ1������Hq��.�w�<�'�3��}����
}�d$@q�<	�J�y5�!�Sŗ;�VPP�hDp�<郏�=:���P"ߴ`�F98�EP�<�b� 7\�P3�l�#"���L�J�<���ͣ4�R!� �ș�p<y��J�<q���f?�q�,:�D�0w��p�<�lT��	pm��-��	��ID�<'KφEh����-�JH�v�u�<iW��	{�(�C�����	Q�IV�<��(
�Os���͊��AK��\T�<���Pڎ C`
���D����S�<qL�">F؈��Μ3����b�e�<٢�;ڐA���F�"1APad�<	�_�.������OS<0q�C�_�<�fƓ;��9Hd�
M: ͐��FX�<q�́�jq1�i�y*�`���z�<SE#ojx��D��}�z�KPjw�<��D��FDL�:�G�����!�G�<�pj��;�p�I0 qI`厚�b&HC��::b��/����$�@C�Inܸ�{�h�p�b��b@�\�JC�	3p�5�d�R.j62d%yIC��6fx�up��<~�>9`���J�C�ɩKp-ˆ		#�<��Ï�?E�B䉚M��Vn^uc�m1��Q,p2~B��"n�5�S��Q��-�c�Âw@B�I����+ֺ3U��p�'�VB�I�@��v"�޲qpe�	A�C�	a=j P  �   "   Ĵ���	��Z��w	ċ;Z���C���NNT�D��e�2Tx��ƕ	#��4"�V���Dǝ���&q�Vl*f�=`�n��OP��HKw,A�a����+R��%��"P�uנ�3Ep���Ïp�r���O<k����\`�)D�0 ��b�'P�ad�+,Oiy�ǛĀ5�O����8z��k`�̴K_����@��R�����]�Z��G
�l���2n^��RչL��R�T�+���1$�pqj]"��#�$Q�~����!C�AyB�J?I��={r�&}���6V�*9��nK���
���(w��0���g�I�]�@��5�$�w]�����O���1��:?���F�!Z@1��OС`�H��O��i1��-m���O�����7�r�S�Τ���Oʌx�o����3N�EK�Q�	���*k��7T<M� ���l�%�a���OJa+T�/J�'�`�r��F/�~r�S^���1�	*O}�쳀`H-W����� B��c��|��dh`��N>Qԍ�,NB��;��!n{�-�3��-U̪=�Y�������l�p?q�<Oĝ˵�۸�?��ЏcVh���޾:Ґ�GA���ܢ�����s� E?��8O�$c%���D��{��	�]Ob� �'Q*(w�T	�R�G�)F�-Zz�'��e�G�����O���0a�G�,Œ��� {������	�Ld&�s �T�
�~�I��y"nA�\�0��o��q�֪�"y�x�"�,�M�'�v��2�E3��t��\�2�Fu�7{���[D��l!x�Qo�	؀X�I<�'��0Z�Z����,Dh�ڹh��k��x}�`V��5��������F>�䡗�0l0�ԁ���?j�(���7N��Y�&�o����F
t(���݆A�Zx�gʛ	�剱v)���a '�dA TqH�+�x��Fԧ �|}��\�9B(�mM)s3d�H>�@O��\#T}�<����T&F�0��7b����胎'����
�'�b��@ ����� d  � @�?�?@�?jg+Q�b��YQFS!RTM��6����2��y�uOv�\]�ȓ-��mK1�ٗu�&�p���G�X��	Y�� �X�0���9/�#�Ԇȓ*T��e�z���)�I+p�)��k,��x%��'Ղ��"��fA�Ԇ�;iI0Q�7�V�B+I,-�<!��fHܴ��F�,mZВ��1&���ɂ����9�V"b�G M����̓�(�!��E1@u�|p�d�
$>H,��Ȏg��)f��A�jQ�����������b�J�F{��9O� �Y��D�O�D`�'b�n���:D�>Y���)ʏ,�Z��3D�%$|]K�)��!�$L�{bZ|2T&��2l���㏜K�D/�O���d�,D���vؿ^֕q�"O�k��=��ez��	>��"OT؁��V�$�X�0�(PG��ţP"O(\�b�5t�A�Hϫ'}�4@�"OL`iҨB�S��pq"�F90��Ż�"O��*D��!Jv���V�N�B0��"O�HMS�F6 EBV犈��,�"OR��P�F�J��e ���z�*u� "O&u��mֺwz$}����qJ�J�"O�0a�,^L]-�iA�Pr�B"Oz$�����d�� �5�W&�
�"O2H5AK-E 8D�#ī&Zj�'�@�'�Xi����k����ʖYjX��'-��A�ˤ�������>�<��O�ٮO赧O>�yGn��62�%�"(Y'j��3:D���"-h� �C�;f����N2�J0w-���>�A�Юm�B�^�4M���35s���'�*�"�-�-r���"h�J"�B5�$�|x�<�ҤK�,<���%O5�PX2��7D���±!2��STnр~N<JWLTh<1�I$�0$���Q(*�Ĕ�B��BX��EyL�F̻�ؑJ�Y[�@!�y�,��J8�� ��F�(`g&��yG�K3� �� �>�¬@���y��ƒd���ۥf�<K�<3$���y2/R�#��r��?B瀙�ڨ�y�&�=U�AZ�B[�B��������y�'��j��P�R&o�:@�ҍ���y�Ȉ�-�D������S��0¢S��y"lفb>��cW �3�)R�!�yҡ�cZ�t�0a\$��9
�y��X�L�hL�W6Wl����A��y"*�B�S@����8�����y�4����w&��	����dJ�6�y����JV���\n�ZX:ԋ�&�y2Ҝ>_
ђ�A�k�(��s�#�y򤉺r"��@�f���CDE!�y�gJ�nnx���΄Y�>�*�&U��y�
��p@(�C��F�� ���y�͑)�\�@�o�AXCM��y��ԬӨ�BaF�}�vx��K��yK�g�*��
�{ee9E�X%�y�(	�0�Dy���k<2�Q�e �y�a��;�  R�f�"� 4���y�+�:��� Ne~�ȸ�/ɰ�yR�F�~�jˢm��]	�`�����yҍ�4~�5ȃ$JTm�iAAd���yR��7ЅH#CH���Ѡ��y�b�='J�Bue�@(y¡��y�E�skX�s#*�;��jrI���yb�
��DK��J	5y����B�yB&ղ|{�)K#��`ǒ�y"�V�k�r�BU/Ŷ��lҦ��4�y�gH��́ԏ���y��*�y
i+�A�Y�X���% �y$]�$Ej)*S�@:L>V8b�̞�y��ږ.bh�%͉�>����ئ�y�ǶR����� .0�tА!��y�i):��;�����{�a�G�!��aC��Hg��CI"�Hb�(�!�D�=�\`sc���I�Ĩ��-�!�� 4��A�Y:Tk�b��b���5"O 1%W�!)�2�!ը	B���"ObIp#��4.�p����>uT��ȵ"O�T ��_�c���r�n�
Ns"OD,
�H

½�1��t< ]�"O�:燊�2�3҄��IJ�	T�'*�8Ҕ��8Vک����{�Z�1��	uB��'�� ��	y��u�� �
i�a��'+�@�lF�
i�v�O�oZ��y	�'��M��oӚn�V�Ň�n���yB��7Ĥh����H����؀�yr
�u�8�#�ڛL���>�y��ˣx*p�j�ば<�*U�$:�yb���m���Ц��0N��q�@���y�ב)��D�i��))F�����y�@2:m�|�'�ك;��r#m�,�y�M�y�2U 6�MO4:��'I]�y��3�x�W��D0.q�V�׉�yRa��s� i&�����U�7�y�/^�9�	�&��;QZ5�X��ybn�6O�!��������ĉH�yr�?`��;��4jQ�EKNS��y�͐���ж�^�pnᘧ@��yR�Y��#�g	��ʗf�
�y�a��1�,���D�U�42����yR��4�Ve�W�I= � l��yB�N��B�ZF+D�rL�ɑ ����y��"A#�hЗ��}��a1A���y�חq����.��Jq;�Z��y�%�����[�"f���
��y¡ֹkڞAbW��?��*��A��yr�@�6un]
�m�[l�Y�G-�y"��4	�{���j�J��p?#��:��d��2�h����J�;��,��$Zh<ـ�E>�����B�a���ȅB]Q�'V��g#Q":b?q(ʇ)	pͻ�腁:5<����'D�<�F��|�&�`a�g� }�U8O�뷬�	 �Qh��"~z�O�
y�����wF�t�D+Y��yb��Y<��)l���������$ą:;F};D�W%NM��ɼ>, ��[��jdƀ�
v�'�t���́ݘ����� ^(���@Åb�:K�'�V�,,�@�)$Ȍ}V-�1��?��g��$��@r�eX6o�@*�畻J{�'n��4Lϫu���!d�M&����'��j�wd���԰M�e��LO&��th
��'l��b�İ�d}��F�O8%b��&n3J[a�G5p��ad�#	��F�b,����'���D6"�c!Ѳ{h����d�86#���a!ܢ����OaV) ��H�`prd��y}����M�j�L�v\[�ࣣoı��O�����7!69i �W��t8W�O���)I�Q���'f�8KB���Ʀ���0 �%H*{n"����I=iP�7gP�-n3/�3;��m�� �${q���ӨYF�`�6*���3�F*9�6���儯Zl=a�X�9,v��++VX�ҕ�V6/������(�y7���d��x�!(����C�R��p?��$	�>A�Yr�'�a�zł�.�)_�t]8�CŧRvV�@���ؤ�%�A;RlG��b�vݲ��(\�xE�'�XxgK�(B�A�e��848��$��t��a�҄Y_�V�[0�@��D@�c�%L��E� �B����;�D��YU�
!x@��;t �J��� ul@��БG��I৚�P���t��r�Ȏ�9ޖ��+���r��&�σ<ܒ��u�Q�3� 9㖤O+�dh��D$g#ԩdQ�lJ�����3[3���'L�
,^,T�wF	V���^)~�B��2E���t�PA���\<�7�(Y�@�tO�-���.�t��S��7>y��b�κ&�h����;�$�CN*~�Ae��o��i򡍋�'8���� G��M;��U�H7�]y��GR?�0]F,��f�ݥ��ɝ#�� �b�H�oȊ�3�Qf��>)�h�*����vLٿ�Ɉ��$��@�ӧ�"Ch���U�<4�pq�Gŗ<tD4RA��SBi��cL�ty\tER+�&9R$���#.4X!��o���~!_7�f=�1�y���e�R�.�Q��)V�Ѡg,ȦY�����W#,p��ۅ���S\@cUH��4��	��`�{Ǧ��g;Ѝt0i������<qgءj�c*D_<��`h����͹S�`�s������@� ���7R6��q�AJ��c�O� )�dH�$o��Z�"��	H!P J��I↹i	R\"r?�,:0)ѽO�.�	E@��!1h�K �b�0Sț0����Վα^4��@!�3V��1��	�Y�� #�R�/
$H��I�t�	�c��	g��ۖl��ʝ�n��9!8�����?k���.	q�����>s���.F�br:�م��T��	-u5��c�;��
��>�X�2��	�:����/aӺ�ۑ'X��@u#W>[h�y#�::o�yc!�T�2t��'Qn�Ss�� [�i%ʝ;;�t���Eǹ2H�1�UnP%W�Ɓ�C��*Z���_�}"5�;=�j���w�,4-�(�ĉ�$���3� aI
�$�0Bd�� �:�G��=�����V�%�rq�'6�5�SI2pv�Q�j׷� !۷C�:��9�q�&�~mS��O=,�@p��6@�9�`O����Oz� d���6�,96`þ#�<Ձ�/Ƌhq���@� +0��!9��'Q
���in0(�fW�"L���TJ������aƃSm�O��P&[�i8��NF<7=0�:��'d��6��R�j�KSCB(&���p�ƚ3o
.�A��ƽ44&�B��b��"�Č<	���u�)>(��"j��6G��`Y\�>��퉘k`݀S�x؀,�d��� �>�衙!��\X6�Ɉe��hS�K�o��Ԩ4Cc��P+L5�� I�f�
�.`���=P�.%9��'�Fɓ�$\�-F���{>��9�D#���'ɍ�a�X��GCI�`N�] �J��~���pF�řz:��aV�؇$�ȈW	��c�V����� .A�u&�4=�}�@�l�'�ث%���2R��kL9.lvt�Z�����
R��xi@�ڨX~��BI��/�dQ�AkJ�Z���'�������W���hI �*]s�➤����c�-Җ?'KP9D�T�p�uG�����K�ɂ�{N��c9.�pWDيo���yQ�	�C�H���T�
~�8D(�
un>P�0iS�}�ZY(@ ։E�F�h�f��p=���F:��|��L�-a��Eԙ({`��쏦�Zl�bQ�HS^���=��p��E�+ e�4ET�)~l��`O_���Y�C��X' i�TY�����AC�R�ѰϞ<Y����;�)�����?�ym��t[�����4FR�d����{��Q�� �o��Ȱ��jW�@�W��h��Y�A��\�1��\<I�O���w�5�hY�&�߅��Z�+	:|)��q�mV6�d�S�V-���`���"cnTk ̀69�~��Bh����q���7�H����*��b�`y��2-�r��F>/���2a�$ƌ�r�_� WvЛ�"+>|Ab�.�:Eg�>�s䅃�+@���E&��p�b���T4b@�C&T�ZN�1�L5.�*�r%�ƴ��<ɴ@���`�.�U伨I�(�>H��QMͥ/�&i%Nڦ��g�@�\4���D�'��iq��?}�<�U(��ir���jN�yԘXӗ�	?v�a{"�Z�h�f�n���$tw �rHѣ�X��p �i� �.�~��-Kab�&�@�>���'ɟ1-�=���Ii�|x�/]�E�� 2��%hB�xa"�	�% \�`�^90���y�@�O׊��`"�Gꉳ�A�n<�A"@��:u���!���y,�l2J��wnX<>� ��яB��f��`�,r��'e*��J�+"ϐ�a�']9)*H�qqƂJ��zBl� q̡�2���l8��djN)$����.%V�	�FÍO)���#O�:Z�4��d��6V��rE��:(4��S� KG�PHC�'��M��j���}q*U0,� ����_���Q�E�^�ڴ?��!�K�=a0b�i��I�J���a��L�|�Df/s���A�Y����FV�q�ܜ0%��3O�D1
�m�70�$�FA�Mk�)(Gú�&��q ����0]Bu(��&��(����H$lR<����%n�����$���=�#��'jr`�3��Ÿs�&x90�H�:�NP�6!��rĔa��5gj�� �#v�9ߴ3h,�fl��\
�h���<��Q3�� l��X��M��~�O�6k<^��B$�"V�ъbb	�y�=+CP
u��./)�hW��l3@�������k��0v��Dj5��Iۈ()N0B��Q
e�]$A�{�����"7M�H��d���%���ax�:�%�=��� ��J.X@\a�O�_�6-_��Tm���y��D �P쫖CX(�Iqb%��iL`ƭ�j|��3'�Q�$Q^����'g��+F苐*dfpcV�x�����S .:e�"� 5�h%��+�>y��[0� �v��<]�|q2I��yy����?��L�7�'FNi9U+�'��>�+L5y�^�9���W��\���+;�ش�D�]��mQ�f�	z� K�Lx�,l��kU���y'�,�PsvSyl��G�Hr)�m���e$27�T1t�ī�� ����t��[�ɵe�,��'8��(�"J؎9M�I{v�Xd�@ҳk� *�����e��z۸8�� �Y�
�CY&0X����Ji<��E *66�Qb3� 	yܪ"=)��.0�(e%�++�셀k��Ϝ�ra��RP^����_��S`��?�R�iRJ�S�� �y�P<��-�LTW�4��gEQf�y��K3�@����q�H�E$�B�iE��q�R	�+�_M��yD��R;�]
N�W��d��T���1.8p)���e�B- Th�%˅7B����bln�Ǔ�]�&�� ����Xj���I�G3�!�DΕ�D)x�µ����PTc�>A���-}�^Q�Ĭ�!֊mJ7j��~��h�Ŧ��Re�c��-BJɌLHYy��/\O��zB#�W]Ȁ��F��|ǼcP��UQ�@2b�չxB�+S,
0��`	�ɦ&�J��gA87ϲK �-ғ*;�!sd�	&,i0��"�#.��=�w��p��-ء7G }yÁ�z�
����O2�#"I�SJ���a��`���2:+��	�d]X����ʎ9'���!ȌC��X#0��.I(j<H
�C��� �)"#��b�Y�#:︩����g@v$��M-!��� �"O�-Ӏ��� Ѳan؏%�1�p۳|�ah�O�Z������ �!Y0���D]�'
牔x DTCv�R��5��/�N������h16�J=!�AC�a��D�� #*}A��פ..�ES�!\E��0c��� yt]ʢ�4��O<A˵�>c�$̢�NTf1���I�8IەÐ>b�&�	�Vb9��'+����iŝ_:z�h��F�!�N���y�T���V-H�Q�P��$���9��8�!�� ���������G�(��Ub#"O�`iCLDK�P��eL��z�hE"O�DX#���M����@���p�L!x"Od�����45�!Xb�1P��dQp"O�R�BT#/��<2TgQ�z"O֜�J�n���I�F� ��"O8�s���|����fF���j���"O8e�'���4U��R�	#��5"O8RGL�1��W�ߏB`��d"OVPCAJ�k�`�7�W�n��1"Oؙz� #O��#���!��H&"O�z4��a���(�	з���Ӏ"O�*�L:�:�ԋ�h�v9su"O�0�� s�و�T9��]n.D�Pb�F�?���� 3�f�s�b:D�p���;�ޤrc#��[F1���<�( ��r�QP�	��i�j�*���(aS�t��I�=�JUx��"~�r��EI�md&Uz��]�ZŦ)��G<p�S�`��36�A4�Ϣ&��F|�(ǯwA  �&@f�'{nv}����!��z�e���ȓ>�<h�7�G�rځZ�����%Γ|dl(��GܪPH�ҧ��Q�N
��^�yW,�<F8X�8�"O|#�&��g�Vu��ʒ$ꤒ񖟼Ҡ � V�qe�'�,�@$*\#Wʐ��t��?��
�O�H��!A�r]sdNV�T����}��Ht�7���J�b�`�Sq��)>��t��"&�Y_�u�'�؎}-h�>Ap��Z��bTF��Ӱ��"D� �ЪJ��B�#��\ <ǔ��
z����Ĺp���S�>E�iY,)�������0S6:�H��O9�yFL�C�Й��*�,�V��ɤT@�͚~X����K�3���OʋV�$	p�/D�\�1m�(Դ��u�O�%;8)��-D�  T�Ed�s�c�q��@�k*D���&#ŏ#�氡�J��H�����+D�쫤���|�0Z�l�:|o�M�U�/D�,J�g�z֊��k�?+�P��T�#D��uG�Y�Jh�H��w^����5D��+U��#%����"GW�y��0D�Ț�`�63����-^z�˷�1D���p�]�e��aƅ_�g��s "D������+m(�������l��ˀ�#D�x�D�D����a�^ #���ѩ"D�����A�l:��G�(`n�ъ�*O�� .T�6¤�*�P0'�t+�"O<qY�*V E�u�҄=Q��%�"Ohi(u�L6P�Vْ�׉K����@"O�0��F�.��غ6�X	gغ��"O`q"�:J��2���>�X%��"O�`�����0��ㄜ�W���""O)��C�mxMc����("O1�DhY~��B׫ڵ����"O\A�'ZFL�j�@Z��-��"O����D�a��A3��C�$h���"O�<�e�ؕ/%3D��G�ִr"O�xK`�=*v��V�'�4�a"O�
Ꮛt�rxB#	����1"O���$|���V��d$k�"O�y�BD��Z�B�<�ji#�"O�5Xt�X0��TzAB�b9LXA"O���#�!3�%�Q`�A9LYx�"O��!s�A�_x*� "):�g"Oy�	J�nR�"3���- �cd"O�Y*�Ô-6M8
�2"�9�"O
��l�=6pH"@^�vQt0HU"O� 8�cL�"��hJ�H'+�t!c "O:�f�Jk�]��Ʉ�V�rh�"O8�r�
ԷS���H��"��c"O��I�0j��}�Wf_i��Uy�"O�@QA,�9��V��@��"O8U�l�^f���IS0��0"O�aBBLߏLva���A���D"O�4v��|���!"�_E%S"O�Iv�P`<��b4l��"O4U��ׄ=	b���Ʃ!0�R"O
���aϒ�p�ـC��3�q$"O~��m��%�Hl�6�Q�^��Ѫ�"OV5+s�wz�a�3I� Ҥ��"O>H(Ҁ�A�z�pi�'jl���"O(`�dF��ȸR�L�+$�T3W"Ove#��,ٲ#�G$Yd"O(�kE-�l���9�M��"ZܩZQ"O�P���dɓkK
CE©I�"O/P���Ǒ�)N6��0#��p3!�d�M�H���kD<r-b$�%�� #!�ĉ�)z�b$�N3	�z�#�)i�!�Ā�	������ίJ�,�7D&�!���dڸ�ђ`�-c�N` Rf3;�!�[�rI6������|u�$G�T�!�N�-{`�i�o�#��1p��@�	�!�$ǿ'���pS���z6���@ 	!�!��%ʌՃ����OpT�J��-3�!�D�f� �Q�H�&Rg�L�ѢY�$�!���P$T�1U.R�jPJ�! ���w!�dނ]�ЁQ.2]'���X<^!��}.�)u��4s&�e�m�!���*IB1�p�t밽2b+ڌd�!�d��P^����8�
�����[#!��Y:���2�G5Y�����h��++!�D}�Lɣ�D7^8��,>!�Dڔ��a�,�,S)�-�P�,;!�$/_&�љ�f�9/� ����P�~�"T��x���?:��3����yy���Q��x��͎_p9rC���<s&��5��O>���b� Dh��~Zu�Y�l!�����(���Q�<1BI4*��A"�O�?M��y��	���H����%Q�x��Ԯ>?E��C�"f��8�gւo�b��3�$�!���"I�@�kƎʄ6�d ��֎-{�ɳwP*�aV���C�~`��{1L�G-�,�29+6�ʞ'�䅥O8abv,�=N1O�)ҕ?I��C��+G���nƱL��u��59}����^p���>k�0e���3y{���3#	�}LO�$17��>�2����$I�DP�On4��?��(�Ed �����S�G��<���'��8�%��)�|���� m�X0 ���.�`y�"L+j��5����Q��7m�,-U��(���O�hJG�Ӎd� �.�:�xP���ɺ{�b8[v��<v?��̟�!���\'l�8
�V,^�~�Z7I{�ޑ��̕B����+�-^�.aG����[����/	�]��$�1)V�~�e�{N(�
&PJ�2�q�[-[\te���S.f}���`��j�B���T�s�V����W-QR,x��	��w��eʣ ��IѶ�s�	m-,�8�(Z�>H�D�� ?,(��B�r��Y�S�U2M׼���ҋh&:��;0��'d܊(���A�A�F���	�/���.O,t
Y w��dD���6OC��`��v�x%�D΋o�<�ѡ�/	Eh��gB���V��<	�oR&��l�%df�+�Mu�'�.�X"�ڒ)�|q:1��?1ݺM3ď�31|�R�f��.��JϽ(�"c�.Wh����	#;����2����O�P�� .o|"�H5L3�4���Oti�c��(7o�E�6��6Z:xI� ֵ:�Z�*Cfنop���X���'Y��=�����w׌1��@̈́)����@�}��Q��
$����!l�́k�7D$�\(�hɻ��6-�z�����M9ǣߣ ��:��-r�W�"@�P,;m��~���i���n�G��(��Z>ee�����3;�� A�hJ�E���M9Y;.�Aǜ�$� q1CH7z�Ќ��S������:���R�'|Y�ppc7�[z��SJ��&
�E�'�H� 8h��G���fM�p+W"_����Ƞ.:�2��V5�`	��m�}�(� �n��� RQ����<X������#\�����O��B���;��!�r��:�6M �߯@�nT�J�*�@�۴(21�iC�Y:��(R�lf09�� �2#�2��$Zd̂�.ϱ@���#g��,sU����_��(SM];sm
�r7E@�]�֫a���3�N� _��]�>�x)*��޼y��A�느~�p����:�D��@ٝU-�������9$C�ț  ؟S%��4�dr7�I�}��� C�@��j�!tG��"�H�����1��j������DG}r��:	I�)O"!p%��+��%�V�!��ȐA�4�H��؞;�`�*��֜)d�SAW���aC��b��K��dʹ_�huJ3(ӢhQ����Cm��@�YÒG^<a� �,Q�$�aD	6+t��CQ�jӼ��uj؊V�T|K�gIh�dg(Y�?P��@o%�O$�a�؅;'���ƃ��	#�hg�Üa��a����o1����"�s22��?/����#>
*�( �3�����i�)+���h�dI�]���'+���D�:��h��*S-2�Y���d&<�c?O6�B��[79��m V�B�?��\�4ʒ�=�e�C����􄁆�ʽJ�8f��59�e#��N�w.�耙�D]
/$		0��_̚]
`��>���C�G�<��yȥl$
\��ڽw{�Ň�ɿ)lvЁ��ߔ#R��H[;[���DG98�E!b%̀B������=/ch��s��&Z� �h��]����R�G9)�^ Y2 ��]ݎ�Yc�ٟL5(��
O&y!p�ІL�rU)�χk����5gӕ�Y�4��@�L�VJٻY}0MY�LI�xU�$φi����E7�,ys$��F�b����$L��4�'� a�"RHؐ��@ؘ�L��phMo�09Kc�M���qυ��ڤ��(������X�B�᠈��h�*+O��ar�.�Zi��	
�|����	�=�eK�Л;ZN�(��-�ըmP�0A�9�
��A����ӆ5��	s���!��)�-� Y c*Z�4������
N�f����V�W�!a<Q��e_�Ii�?h�t�"��RP�q�%^����Ƭ-&o m`1�A��YSWl��2�$�h3$�5+P��N[5�K�3�&���] 6Lt�*��N�zHˑ�W6?ԝ8��X����$뇷�bY{0��'8PL�%
�O�ft�qN�� ;ލ r��/��X`/�?��5pG�\��{R�؂t��٩uLJ�)dTCUd[�Y�j��@�sf���i��D󷋘,!�T ��O/���v
	6x���zb�@�W6��B�n����X�E�O��<�:(S���Նf#�]zs��T�zd*U~DQ6�٤4�F�[�d�:K�n���酽8�"�8p`D=CC������,O�@��S� H�DH�N�p�����RE@F������6��i���J�c[��Q��i�"���`� �\Yx6L=��&�ݥV�
�ۃ���f�Q�ˀ�;s��"��/5�,��qA�Q�l�ڠ(6����*(���b���]��[',�:�.���* +�����L�v��6�ӄR_F)��ۂ��)��Xp6Yu%���|15�7�`e1 [k��8	�,�x��m�"(蝁R$�Y����3�:c�Ț��M3"C�/�z�FQ$bII���ȶ��4K�#PaizVDз<��XK�bU!T�АA���?@�!2�*S��O\i*���(F���IS�\::s�L{�'#*�j$�_?E��H�X.~kl��TE7t�s�/n�f�EOL�9��܁� �{����`��3[���K>��G�X�z�*��RQ�)�d��{brl����+gZ�Q�Y�H��㇆5\�l�B�E�O���J�1}n`@�v�I�e}��-Z1P�0�����(h��0"&�M�=Ҹ9K�S��<1g]4 ��$)��C���E���Vz�y�ѩN�h�Q�	ڦ=s��9g60�I��Mk�O�촋@���XP��l�{�A�>�������GE�9,��a��rwi׍���mZ�61(�)��®C�*��4)o����7ol����&[:��"��b�ś'"�&���ӭ�<_(D�&�	�u�쑰��Ȅ8a�HS�/�ަ�;�_.&xl1�OY(�D0�?r+���B�G֦!�c��l
����D�}SR̠��^1=_�}�ƀ�x�H|�Ip���
u_��5��3 ��]�o���ig�2_��{���N�(��+˛rP�)'�0A��C�VL��v	��*j�ybNX~�*d���Em�.��2f�%"�M�7.�&��O��#p͆c��D{D�S�(/X�Vͽj�XP�h�7CO*��i���� mӖ9�J��p��� 7��i������vĞ=C�쳇�G�/�e�A��)�0=�����$|Yd�,?^�e��F�=�a;��ʗF��ң��7:h��!P�<����,��i����K��5�Ѕ
��ʨy�e�j��%h��P~hu��6[�$�&) e���CuG��U�،1c� 	���2�!fud�"�H�0����qQ�7�Y[� B��%�6,z�΋�G����U�I'�HJ��ib�J�fÝx xh��$}YP<��O��#�Àt�(���ѝ6D9y���;)w�=+' �	���+�XRƈ�=$�u�DfX ��H�҉U�d���;Ҁ��Kk�1�M�/�VjV�	7/F���7e�+FϾ!�fH�&1��h����zU�R�l[#m�6PjӋɴ(I�������McTQ�Ikr9͓\Y8�K�q~�:V�΅7��l����fѾ��1�'����4�0�hp�3$8���]�a��JZx`C�ؑG�å`P2����'ǂ�H��ݮ �ЬŅ;wi$䂥Z�h)�"r��
����$�6i禭PD�H%c!,�
��D0�;Di�1-�:����^�<�dR�F��۪O��"7��!������H��Lidͭw
�0��i�p!�C�43K.��qg�C��(�;r��%��G(i2pő#?��1�r�ʣ^�$����T:�(1�c*�-}��,��|�Z��s铡<��-Њ�K%<��`;A�E!��dZ�F�1pqO0�zCo͚<U8Ł4'�^(��W��(1�ʨ�f��Q6瓓l�(붦���)v��at2)���'�v���*|Ce���,nX�� ��N �`  �WP�ѢFE�xO�,���.ç_��"*�Z����d�!�DΘ?G��16�����%X�䆧���3�͝��D��L"����8Êb��R�M���B|���V�J�Qf zC��*1�qaq�;�O�\���Q�|e�s� ��Ra��k�U�aDJ�"�z(��,����FY$B��
�.��CY��R���|�L���"j��D7pdQ�tg��}�D�#b����7�~��I7HH�8a!
2�F�p7l��-Ϙ|��D/�O�aS W���Yc��ru�l1�"O���Y7d� �p�	�.T�-�1"O8���c �Q������+M8��"O �Ä�(dLNe3ХȨE����"O���$_)V *R��\�Hq�"Oh����%_���tCP�K�J�u"O�� J�HS�-�p�{$Ԁ�"OQ��C���hA��Cȕx�"O�a�m�zVaI%��%#6���"OH­%O�<�CT�E�Tt��"O��8��F'T�i�J58��(P"O��s�@��y0l5 t� f��hj "O���1M0Y�l���Ιx�� a�"OP��u(ϰE`]H����3*S�"O�4ZՈ'1n�h�d�_���g"O�D���ڢS���q��xK[3"O�䓓����9}� x���x@��s��	��	�#���!P72F^�@�<Y���D�-s�DpA?x���N܀5�\�,��B�Y"�m�AҫC�����Y=<F">�q�>(6�hB%5�S�0�8iAD�.���r&Z�rf:B�/y���5F�Z�r`X"@[�F���	Xib ��J�&�S�O�b���#Y�:��@ �)g�Xh+�'��҂���H,�C"R�t���O� a�A���xǓ [��R��>����7-�&x�����	=DSN)�r�#]@�c�`\���𩌴$���
OT�Ґ"Ӎ@�&M3iR8Ff<T�I
RDL���_&jEq�~q�j��e9�!+r'I�V����"O��kփ&R|h�Q&�s6�)@E:Ob)PR%�b��!O�"~�`��97�,i1�ee:$��l�h�<)bn��%R)C&��M�P��w��O�Č:5�ƭ'�",O�+�`e���!f�*��b"O��X%��F���K����j�d���"O��aD�8$���8�R� h$"O���V��n�J��%�-H}�"Ot��Oջ#@�G+XaY�$@ "Oh-���L�4��Պ�iƆu5pT5"O��cs
��U*�����-@<��"O8��$�
m�}@c���FHtq"O�!�p.�2}V܄2��ؒ@X��"O�� C��bQJ��)
/���&"O�q�W���#A�Ȉ���$F�0q�"O��sQhf��j��#4ԼX��O'!�$#"�b�Q �܌yI��d�!��*�|���x�����%يc�!�D�!Ǥ�"`Ŏ^��R㖾.�!�+B����(�3w1je��1�!�V�6�fL��N�<�*�ZD��14�!����(�������-'��=�E�	_�!�$ſ1T��u�R	y��i�E�-�!��ѮV�J$+�ʜI�$�1g̍	�!�D�(#6	3�܃y�6�X#k��;U!�~���H�,X�hb
}��kU�\H!��U>�:Qn��n��03�# bQ!���+lBa-T�%*�,�W'r%�"O�r�I�[�qq˚�`�l�5"OV�񠆁�5��$�#�\�*e�"OF�Z%���t20pX4���^%q�"O|�BR���Y_>`7�0AZΙI�"O.0��ǹb���[@
9l:�(A��r<Ȫ&�I�`g�\j؊w�꼄�S�? �Mj�η18$ŐѨĘA52H�c"Ox8
T*�n�V�s��l���"O`�0e�	�/�x���F�^���"O���2
�Đ:�Ã�w�"�[P"O
�q�?(.m��a�*_̬�z""O~9`vJ�	�$ANɯK�%@�"Oʁ�h֞ip��Yld��lx"O��`W��[\VآD
> ,�`1"O���FGТ%���N�#�"OL�`��jA�h򮝯/��=A#"O��4��+9�����*R�*ِ$!�"O�SB�U���ȓi���!"O�����.ܬl
�.�^����t"O^IP���+��HH0�	����'�l0p�C1X�*�a��}"L����7U/�d�
��V����˦
aF�XEm��]��P#.�2Rz�\���mӪ�Z�K|�ƌá��6VjyqÒ?7-'?ͧV��`4$G�U�`�#��?��`U�� FB1O���.5�E��)�J��jB7r�b���y�J�r�`�~�	 %S܍��"J�V���Do��� Ot���f�	T��U��@M�SJ��a��ۨ	^$A#p`k�@3����fk��&�"~�#&L#y~� �,���-Z��X=c�0���N0�����	�eȟ'�����m�Dp��@B�}PqOdh(	çۈ��C��^��$	�D�<�=��$ "t��	,�v�W���o^TyQ�N�(��޾����=�)�?�>��UB/����4�ڲ�N�	-x혥?�)�'�@��W�U*U� A���3+�4�`-zD^��'��]�A?���XƎ^A~t0%ㆺ<�����Oe�����p�V�ZV��̺�K?�����/2���ꎆD����Q4���D��A'4�b��+"V9�lE���8��տq�B�e*�5�u�?����'✁Γ��bg8l`q��U�:� ���'w�o�,/Դ�'h�S��a�	v�	8]%l�ȜsFX�8Gd��E�i�b�xJ?�O���N_P�)�K��s�������� 1�`�h���LS���<6�eȒFI�ɍ9yn(À-⧘?A���|l�q)��@|pXp�M^R~���5����|���E��]����T�3Wx��W�8x+�ɏL�4ka��>Q	çk�>!�Gf�~ղ|� �ߚ<`�V�S�{eD�G�O��m���"�������`�2Ⴑ h�L�1k;
ec��@�*,��'�؉�W�@�Bh���#X��9��'A2�cT��A�mX�W1��:�'n��R��=m��K�.E�N�
�'�pPx7n�<g��B��[�I1��
�'�`��ı5�H� �J�!I$|�	�'�  z'�H?��J���Ѻ	�'粬�BT%:3�$�Ӣ���h
�'�4y��矒"�>�@����p�#	�'<�\	󠎺k���[�s�p�	�'�RF+��j
Q��p�r�'�x8��,ۤ~9�5�Df��l��Y��'ʂ�D�L�h�/U�g��t��'4ⱓ6鈟T�J�1���!Z�t�	�'֪ܩ���p������_1IK����'���g�* ұK��-:�t�H�'0��5�%?�`���[�B5���
�'�آ�+Y�y�������v=
�'J�
���4��e����
4��	�'���G��"��Q��1����	�'1�p�1�;8���i�̇�+�R�K	�'�,`�Ң)��{�F,7MR�`�'SXl
FkW�Q��Y1���/� q1�'������9\{ӏ�!"
��'^P�Ҡ�^-YE ���bؐ oC�']T��9u�A ��p�'�.I��ĭS����(�9EĄ�'k%9ъ�p9D��i�$�pq
��� �����&-]�Xɡ&ψ5��E`W"O��+ìW"�Аj�K�~���@"O���J�_<���)QK���c�"O��tB��O ���皚Y���A"O�S��5������(�z�"Op9qꅱ,���y�+��R%cv"O�Aa6D9����F+��D�D�U"O�+`@�B'��1V��z��M�"O����i�s�|���0��9��"OF4	��M &�P�+i؏%�VC�"O�xh��S!�XC��X��8�"OP[�&_1��@��/K�Z���"ODE�m�2c��GӲVp>
�"O�t� !��,f��)MUbN�+�"Ov�R��0��Xy�&˺ �R�b4"OĴ���	�x�$U��C��ԩbf"O�]1�f��퐈RԂ08�N��e"O�*�i��c��e�wBL��0�8$"O8��� �Y��TZ��x��H�"OH��V$,q<-z3�*W��]��"O>�xA��,X��@���]���xE"O����T2/,�9���2$�ly��"Oԉ�Pc'#��U��+&dԪ�"O�%jv.^��d�I"�*�3�"O ��cᘫ0{��2����\��"Op�	V��$����'옵a�rx��"O���æ����"�)g�ntB�"O�|���3A4�I���/����"O��Q0��$�h����Bw4��"O(�	NӁNh|��Ǒ%`�(�0"O  R&K �1� �J�t#@I��"O(��7<�4B�5��9Q"O�͸%�Db��Y��F�8�]��"O81ӤD�w'�5"�ʤT>��"O�-)6mK> Hir�[9B6�*w"O4dp�NC$�FXK\�8e���"O=;e�[�R�������G�|��"O�L;&�R�]ZQ�t&��=A��t"O��*WO/WH��6f�K@j (�"Oxm"N��gn���%��� 2"O ���:
�@�dW nb�:A"O�����xT䩫�$�ek&	q"O�r�D�dpq�s��1@hl0c"Oj3���k ���؄ ~<%��"Oz�x7��d�+p�-uiD��"O6�r�aϔ_m��xr*�Q|�Ų"O�a�Z/C�0t���ƬP]\���"O0�����+8X�9�@"���&"Ot���ꖂ��1��K?u|�'"O���K� 2D q�㋓50R�D��"O�!x ͈Lla�`+�1��`""O���"�	P����jM�T���"OT���3M"����o�#
f�c "O\���K����H��H2g�� d"O�i2E%�%@<Al<y��"OX�;��$��,�̘�H��岥"O���E�S��)b땡Dܦ�'"O��0�D33�,Xq�	I1q̈́+�"OHhK�<��Z���$Fv4��"O���@:��4���Q�b�P�""ODD(�	F�M�<�)��ځo3N�@"O ̣�ꎃ,9��!��
�#-�!��"O�|����PD&�i�ލ��*�"Oxx�R��4�B��B���F� �"O� ��f_�M��5�ӱ5*q�U"O&��f��,1���g���"Or� �g�$&�;���J��p� "O�C$IƪPm2E�6�џ=�(%�"OlmK�b�F}��P��_S���"O�mjg��m;� I�/ir,rt"OV�b��8E�J�J��g&�d"O^,A5�[��B����� Q���%"O�<�b�83/T�#S�3N>a �"O~�!P 4	�l��v�X�}/z��"OD����q�D�F�J�x�T�"Oe�E.�hp��<�*���"O�<*ǥ\1V����Ɉ0!��%J�"O�,c��\�RH�§K���p�"OV$��	�8유�h�+�Щ�"O��[-C2��욠��!g��-r�"O^���)�I�ܡ�7����NLJ"O�8�q�P1Pd� �<<��(1@"On��t��}C�`��Z�n�|�Hq"O$��� -NNT���5}��"O�8���_�,u���y�Qt"O�E��N�#�1s���)m�Ts�"O�l�6�/#�J3�3nY(�"Of!�p%� ��]���X�Ax�x�$"O@��Y\��+)��Vvd���"O��v)�{g�嚦Ȑ;[\���"O�8���Ҧ&�l��t�̊;W2$��"O�KƁCxH(��ޒ/\�-2b"O�tAZ�X��ݘ���"����"Ol����$���j�ž|����#"O0�S���1Q��I�F�j�\��E"OT:Da��p���],�c "O�Aq�P�,�b̢b&]3/�Y#�"Oɒ�/q5<m8�N�`Ԧ4��"O2��H!Efɋ$�̣Q(�lc�"Ob����Sz�dr���6&�(� �"O$Mp2J[�D��yi歒�k�ȫ�"OV�ٲ���Y[�}�"m	�XN����"O���u w=Y�큡I�j�"O�qお[:������P�d`���a"O�UQi��l1����BSB.�` "O&��%�T�%7�I�%����"Ov�ynĪ��Ij�CZ81�Z�"O��#p��;�"�����<
�8Xå"O�K�GǾ	�6e�fC�&����R"O����c��WPPDB9T�h�BA"O�1
A�2<��D#s�Z�^�j�l.D��1b�7j�H��@ύ�Wd�볎9D�<��/Y�4��aV/F+09�#D���#�L-�	���7��� � D��Q�	F+F�Tl�A���n,���է=D�x�Pf\-RC�mp��Y�$��$��+<D����E��������7�l��A6D�`R*M�6��|��n�V�J�+��.D���Fg�
�~\�$j��@b�@�,D�`y��T,�Ii�.X<��ru((D���!̔?.��[�V'}�Ԅs$�'D�0@���Hp��zKP#y_�|�*9D�Ĩ�jاNZ��׎ey�E�'6D���V
Ֆx5R}�M�,�����&D���q�LM6���ƩI7J~�{��&D��
�-$�V� �:xS�xp)$D�@{��N�/���F��m��� D��Y�lӭZ�v�����v�d"�F9D�� �kى`x�@�ᨊ$*���ZR"O���M)B����ʑ�z��P"O$4
��[CD6��C�W�q��\��"O�i���	%�Ȉ��QU���"O��
A�ު@�ƅwlY�"O$0S��w�4@óO����c"O�Q�s�l� �SbH���}��"Of��g$^�y�,9d�u+�(H��"O�� g��r����@|d��"Oȅ�fJ�~���
� H���"O�Y�(�2Q�����`��k�~��'"O�mrj�%^P�Z������U�V"O�I(�[��+!	)s\��#k�|�<���p��8��!9H����Er�<1#�I�WF�����#G䘜+�/Gu�<�v��-�"Q;��"�������r�<�4 �R�	�
��匠P �Wk�<�Q�	42�(���DE_�Dx���N�<�S���.��1���ٮeĠNO�<ATʽk��y�&�FR�<�ˈC�<��I%F��ո4r�)#bKEE�<�to§�$2$̅6y�N�
�@�u�<a�D� r� �@�i8If�yՍn�<q1E�1/p&���%�?[��T0�k�<���\�T��=ñF���-��`�R�<AN�j$Z���45۞4(���L�<A��B(YC�l3%�єn���!
�_�<	�h�]��Dɓ�Ҫt���D�<���Z�K��G�X���j��A�<iGH%%��y�ſn��밂�~�<���[)'4ɠÆ��L�:�*2�_y�<��E�7 ђ@����8E!*���O@�<	u�� 4D5��=1�$�� �Vy�<�I�3pC�����CD`���@�u�<�C�=4X�"���r��!��C�n�<���[.srHC�)ձ&�f�13o�n�<�W�G b��-�R�-�����AU�<���7�����V>zZls�"�P�<�$-G�j�(@�`Ď2s������r�<��CQ�E҄�@M-sS�кr��k�<�m�>��t�Se��<���V�A�<�
��i�`� ���"d�O|�<1��O�'@lCw�	�pUp$��@�<�� 8  ��   �  �    �  +  4  .>  �E  �K  2R  ~X  �^  e  Gk  �q  �w  ~  P�  ��  ֐  �  Z�  ��  �  8�  ��   �  ��  :�  }�  ��  �  B�  z�  ��  "�  �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�	�<I������t��v��AHZ�<��#I�JF����3Q��j�<I���!O�"M.R�=ے�f�<aE�İA.��W-��`?fEWm�|�'1���1A�\s��ʾi���
F/G!�D̂6)�qz@AV�TP,D�ߞrJ�'�a|�f _�Mj3�݌w)��a����y���c�pd��@Ojt�`��J��y���C���s%��P���(�jQ�y�Rfܖ�����ATH��B��y�1v}�W���=D�yҏ��M����s�F����:�|����9NT%�"O��c��G~�	���6~'���@Y�(��|�\�d
�mچ�R�`��<�&��ȓ�B��wd�V��M�"��-��UDx��'�(�з��,K'p���m��sM��2�'����F�sW�-X� �-��[�'���!p6RǺx���N���yǓa;Q� �A��0��s���;�F �uh5D�|I�JF�KH����h(�dѰF(D����Z0Y3ܽ��̜�C�<ɴ�+D��j����p��ɲ�����jӐB�	^lйU�Q,�1���NƬ��hO>� �$�O�5���F��R{Ƭ�p"O�Hzf�O�j<R)�mʊ8T��ֹiʊ�Dy���i�6i��)� �-0�/�ݺ�'�:��̉�\V�)�D� C��"OԨ`�ւ�4�w�11j�i#�'n�O~� Ë�i��TɁ�ôQB��9 ��?��<� )��r��8���C��q��.NX̓�~R����m��Q#�e�C?�w�	V!��B�5s��ad��P�*�z��>(��X~��xJ?�3�,�-�/��j�; ,F���n��a	�
�,���ʸ��)�ȓra�0.�`@�F�X�Y���?�4��/"$iAa�=Ҿ�:"Ye�IE��7�	]�"u�`��x��L2�.D����Q�x��h'�2 �Q!EA�>���F�Fi��
7*���c)D�
��PE}B-������HB�x����M�QQ`݂E���!��E��³��Ck|��4�ވ~�ꓬM�O:�Os�g?��T5r�*���*ז!X��JtFW�<��$O#Z�!��F�80jq�֧Z:l�"���������ν���K7D&�4�b���B�S�E0t!��ѩ����'���	=C��~��'tef	�b"oa.A�(����4�INLQ����8Oh��������f܉ea}�S��lZ$	Rf �GC_~D�酢B� B�I&A�e�ע"��i��O&����$�s�'�bq)��.k����C�b�M>�޴meaz"�ȺZC��������|�i���:��O."~:@Y3>�|i%�V.H�h3n�f�<��a�	r�>�Z�B&x�FŻ���A�'�F���	e�`���Q�d�ۤ�!���hՌyшπ6�>8bd��]n�c��F{J~�F��1��`"�E!5�,I��SY�<Q��/��9�苙_�<�@"�X�k��y��^}��p��A�2lDM���կ�y��t*� �@0s]X�cWB��yb�=CߚҥEՅrJ��� ��'��{�쟏Z�$�u&Pc´���A!�y��p�����+)�`���g���HO`��!b(�;���;.m���J�!�D�>^�Pت��#.`%ReU/!��$�Eq��{�z[%��*^�!�DNK�H`hZ v�Ĺ�Ĥ�!�D����Qg�ҤB]����i|!�$�9�deQ¨T .[�p���P�-!򄜀,������:Rz�p�>[�!�ӴV���QB�E��J"	�;�!�$țX�} ��W3��b�9p�!�Ɓ7F4�U#�� �"���/܉L�!�C)�T���$�~��(����:(!�d��9%�i��	M6�h�ꛣ�!�*9�HG:"B��ʜ?n&!�$ǭW5��!��$��(T�ԝ]!�?�[�b`թK��@Q��V�!�d5��X�����1&���7`!��To
ɂ4�B��@ūVJ��*�!�$��1P�
C�kO�50���2>!�\(L� �G�@K ��k��=�!��ҧ.Z�}��$G��ŕ�!��+sZ�JG�
T���W�S�!�$Ł!�d�X�lp�eІd��8i!�d� P�ã�T�Zd�d���1!�$�
Q,�m�dͽ��i��(�"@�!�$��>��R@ .��AGN))�!�� d�a�[�
��z���2cl�8� "O~t w��'j��EA�)�*W����"OfY��
|�z$R��B�8t�e"Ova;F��&)�Q�DW/y,�<�!"O�0��T~��L�'C�*8!��	"O�d˕ȏ�.�f���H�Q��P�'"O0�c��q٨ �Z�m���#"Or����k���k��1F5	�"O8����Ƥ$1"� "F�raZ�I3"O����\�_u��@ݠX0�1A`"O�9�"Z8�c��I�N+�9��"O�8B���"Sքs ���$u��p�"O|�����I���ŋdx�0d"O�}�p�՗'[�S�͎�mT�)"OF�1q�V;��,�I�
aR��Ȃ"O���+��]����Ȁ�p��%��"O�U�P�(iP�~
�C0"OB�VFP==����P�	m|F��"On����'Pu�P�W���#�$t� "O���P��%u[�����[�n�2%Kd"O�ͣ�H��5��(3����V���"O*��1�U(LNj�"���,�"OB�m����>7�Bh�"O�Q�Fה��ɀW�����=�"O�M�VE) ��S`슆=��I��"O���R)g0�ZӬ��5��0 !"O̜�J�=7��ԡ`��J�-h`"O���/�<��E �)��dP~X)�"O�q���Z>j����HWF�<c$"O�Y���	b��m��!�r�UY"O Uʤ�J@!@T�� �ITJ��"O���@dњf���@Y�K5lea"O������=��� ���/GԐ���"Ox�I�:<Z�UQ�G̀�"O���¢�
��_5�=R%"Ov����2��1(��
��<�D"OƠ���|P�e!w��!�����"OP�Lוj���&k��*Z��"O|0�DҮI!�CBI���+""OXz��ʇy'�l�Q&Mm2{b"O�a��]���a%��+aT��F"O:�(�JO�#�!Xfn�qZ�|�E"O>t�5��{�|b��q�p�
 "O������ #��"}�Z@�"O@qRr���5��(�	'ljb�"Ol�aX�N�"��ao	?��՚�"O�Չ�,5  ��/òM�T���"O�I1�A�|�&͂�H
�9rF"O���D眀U����'�$ x �"O0����N�RAbT������!"O�m�0�@)T���Qx�P7"O�<6;n���˚���23"O��	���^����&X�Py�"O�!Q3旑q�l�8e	��%�P�X�"O����( ����MɄX;� ;�"O�mk�i�(yV�ac��݈}.<�Z�"O���A+�#B�Q�׺=R���"O���Cc�
�ph�2ꂽ؜�2"O��K �_�g��A���P�6��'"O�eڃ.�=fC<%��-M>� i��"O
��-�	T����&w8@S�"O��Z&�8z������s^��T"Of����|,��(i� %��Ă"O�A+��W�{P��	�+cC��Pf"O� ����:�j�3�Ǟf,��"O�թs䀗r/��SF�-]��ju"O�A���j=�¡4����"O��`��ٿ`��hJf�Қ02к�"O�1�B���F������J\h���'B�'/��'/��'�B�'o��'{čJ�AK���y����.�ܵ(��'"��'��'W2�'���'���':���!�oS*= R�]�bdA���O����O����O��d�O����O���O¸� .E�*�)�߶s�����O���O���Op���OF��O����O*�B�H�bkB�N�T�,�Je�O.���O����OR�d�Ol���O����O��g
��S7ڝ���M�$�H�O��d�O����Oz���O �$�O0��O�,��"R�kf�PHЄܰB��ђ��O\��O����O �d�O��D�O����O@�'�H�"վU��� ����O��D�O����OT���O����O4���O�0��*�)Jn��S��CG��T����O���O����O��d�O�d�O����O�@�T�X�a]\ݻuK�`>qǈ�O��d�O��D�O����Op���O*���O��&���?oVmYvIVwP�x�C�Or���O���O����O:���OD��On�#G���
<Y�V�2+��0�"�O �d�O\�D�O.���O�d�O��D�O<Uxe��)S�X���W~�:,�	�O����O���On���Oz�$ Ǧu�Iܟ8@��$t����(�1@_����.�����O�S�g~R�m��i�5B�JOV�U,M�Ca��J����lq�I�M���y�`{�\�EMC� ʔa,�&;FZYӄN��=�ICV��oz~R"S�b��(����I�IsE�P�LA">�������E�<�����d-�'���sOB9G�DF!�*9�,!�"�iE��9�y2�Ƀ����(�`y���@��իj�TЌ��4LΛ�6O��Sܧy�RMn��<� "�#j��u/Z�H�:��Wl��<��*ĸm��ź4���hO�I�O��`�i_[^:���2	a?O�˓��TC��!�*٘'#�|ccĆ:Zu,�t�J�p9@�!��J@}b�f�j-l��<�O*������b��I�B�1gJi�����ۓ�D�l'<D�4�&�S�i-�\��"��b}�L���(<9�lb߯C��gy򧈟�dL�G� ���+��S�p+Ge�
'��d���&*?y��i��O�IǊ+nQQ�E 3Nj/ʸ7���Nզ��4�?bd���M��O�/ź2�x�0`��sx5!���,J Q�j5�4���@ޏ
x��abݎ{Ҁy����|r�
�2�돚@��Q�鐴I����ȓ=�\���LLO2�#��v��}�S��9F��I�EQ�7f䑊G�"3�b)��H�^i|����b�ȝRҨ��E}�T��42^�Q�� Y?
;�9��CT�@�B � !��Cp☶q4 d�"��3\5��{��D�(����@H��fb���͂�}^�,!�̔ 0���0�G�T���n�ݟ�����P��	���#6�9���D[�XĀ3��^����'4����7q��|��� l���0��.FC2iZ"�অ�w�ƣ�Ms��?q����#�x��', \�e��`�t(�?"V��zu�j��P�Bm�OP�O>�ɓbT��L),}���H� ��u��4�?!��?95n��27�'�b�'u��� ^n���R��S;60��M�UO���|�BY����F��O���VNI��;4C�X%(ϓG~v�lZ�0������D�OL���OȒOk,ŕ_x����ݓ=?�1�2꜡t�V�'˖l���'X��'�R�'L�U���C�

��Wk����(��@�/1���4�?����?a���$�Oh���O8�Au,]�
d	Y�
�VT�ѷ�^,���d�O��d�O����|���$�L��`�i�2�Y%M�:ee��'��Z1dU��x�D�d�O:�$�<���?���f����n����� ��E�4�:���� ��9���iUR�'��'b�'���3�	�oa�l�%
�3�Z��QE�$a4|n�ȟ%�l��ȟ܉����O>I[4�\��L`�lL���e 2�i���'� PK�L|R���4��H��uUcU�.%nh��jD%|��'\��'�Mh3�'�ɧ�I�9N��$��	E��i`I��s���Y�ڀ���M�fZ?���?9��O���S�ʬX��$�����isR�'��ٓ�'�ɧ�O	�8���[O����Uh�)���9�4O�F�ֹi���'q��O:���'Y�Ӗ;;<1���T�N���!^�w�x�"�4XBt����?q�]d������Oz�Zr�%c�yr�G�+'�8(a�Kܦ-��П���,� ���4�?�-������H��%�>��Ypv�J� �iX�L~Ӵ�d�O���Tx{���O�2�'��ߟD�Bk��hT�mɖ���l$05H��iSRD��>!4��?���?�I>�1el�k&KW4 e@rHҬS��Dn�ɟ�����p�	ҟ���ʟ��I�(��$��K�L�X�����ǴPF �@��ē�?!��?�(O����O$=Ps��6}P�|����Ú𪂂 � ����<a��?�.O���[
��	<�]+��ػ���xQ�X�yw�7��O��d8�����I�{ü�!���9����d�����-;��m'�0��fy��'���6[>M�ɘ8��]w��$J��ȵĕ�bր�`�4��'=r�'��h�yr\=��s�&Y%`&���o׷H��7M�O�ʓ�?�j�����O����k��4;`1��@��V_DL�ы`4�'�B�'g4p2u�|b�~� ��B2>7��Z'%%��0�R����;T��	�H�	ޟ��]yZwC^`���/��*r��LQJ��4�?a��K�,��<���&��0��R.,(���$꒛���i���'�R�'�$P��'&�~y��h�t������ܬc^�rW�i�PH���|ү0�'�?��҄$;�l�0a��"<0Pg�$H���'b�'���j)�4���D�O��(am߇
 ޙS%J\�
���eB�ϦA������I����˧�?��'R�x�p�z�Z�鐉U4��ڴ�?!Gj���dV�T���s���c���B��@���1��8mԟt��?�ԟp�	�x�'�<����</����ȮEG�cT�M�	:O����O.�ĥ<���?�,E��4ju��X��ES�BL�T�#���Օ�� ˛����!�O�'
\dkqj[�.Y6��5��ܱ�ȓ,�μ�@�9 P����gE�=q�(D��.x���/Ѝ���)�jd�@i��bz�@�@�;i*�)�lP��l
!&�px@XS'Q�(�.��
̽*z!�� �¢_���%��θ$
BQ{��J�p� 2�@�9�"�BB��	q`tR����D0ӭ���>Dy@H�8�҆E��#�Al_���I�A_1�6AZ�O�� ��kÉO���	۟$�n �(�xT���ԶA>	�էVb�dR>}�ᛡ	������`b��p�<}�Қa\$X0���"��|C��O�O^�����Z40�ƕ�T�,�I��``n�Otm��M����O8��T
�|}�q�c��9`�P�؈y��'��y�ɤW>؂��K���%� 	�ў��:�HO�%�� ��(���c�l���f2Nt���O�$ۊ\f��'��O����O���\���*?1X��s#��4��4�fH��L����[����L�`�����D	�Z�� �6���5����H3'Ԧ1;"@R`CE'h��X#�I�4xGvm�C�K$6e,LrX>����@����L!�UꗧX�f����� ��aߤ�lZ��4�	2V��i>-������Iҟ���Ъ��%N�#NY{�C�#?����ƓJJ���K�'���:���HX��?��	�M3����$S�-�n��#'S�_��Mz��A�ܨ������ �D�O����Ob��;�?y���TFF���%�TO��B�9 	�r A�ڱ�$�B�df @���
�*�p�Fy.�D��i��صfL��gNǿ[:Z�����	��ib%�`ӌm�$-i��YӤcs�j�t�a�e��b�\(p�_�h����ß�0�4G���'��ϟ��?i3eX�i����^�H�����\�<q���},@Q e̼b��,��C�X̓o�v�'���11mp�p�4�?����ܯ{X��~����?���̶�?����4�6s��a�?�� ��F[���;���Oy������"~iI����	3^�Ey��vy|���%-C��8�E�Z�.�p�"�ff<�Ѣ^3��ဦ�i���2RB"��RFJ���OZ�/���AF��eu�{�]�n�RHΓ�?A������6�i�O<	� t�U���k��xB�p� m1�/A�*�����&�:89�%�O|�]�����i�B�'��S .j�t�	*^#�2ӄZV�ܻ6�ϭtf���	��wc��O�&lcD�1iB��|�-���Y�O߮#���aA�Z�e���>����rPn��*��
��uz���?p�4��ϕ�`TȔ�Q�<<��>V��\h޴S⛶�'��v�!!�^���P����7��O`��ё)��[��2e�$��f�1@5axҫ'ғi�Y���A1T�� ! �Mp.��w�i?��'32iˉg���@�' B�'���w����gȥT�0<�6e�����h1l
�X��NϦ�:��+E�c>�O|!B���!�H`h��U�2!�y��?@>^�/ɝ�M�A`�)?���>�O��1V�T) �!���$;x���ߦ�!-O�(������?��?���#m�x�i���=�s�_��͇Ɠ}V��`N׌�b�����j��P�'��"=�O��I
ݶ��F��\>�|HsD�4@P��%�pE��ԟ8�	џ��^w��'nbH-_9@D�`��j$Iqb:�@ Jц�c��H��	/I�@�s)2��5�I�klE�fVJ�D�P��ʓ�b,��B\�ad�a�W+̖r�p<�r�
��Y"�J�5��' \)8�$�# �ْ�G3k♻@�L/�?��iJpOT���O���S�R�,���Ę:(S��Y��4�O֓O���%�]#P�����?":��s�F�<���K�&�'���%:͆M������>X�r:�b�(7���35�۟Z��$�O^� ��O���w>	Cr�H�7���&���.=|QVI�@OAX"+ĪA:B��ǄV��{�d_�Q��X2K�"v\%�䎊�a��F�F�I�P��d��] ����Jy��	8I!zI{�RID/�?i�i�.�'st���[Nd}�DG#��t�<���<���	n���F�B@��5s�^<C�i)N,��Q�9q�<sEgܙfR�Ú'��I�)C�A�4�?�����IܯOUH�dQ1K��rb���8��aAL:==�$�O���C)� w"�C�4V�ĥ��D@�!u��#��X�t�β��x���w�(���� ��a���ũY?^DT85%%;���;u`JM��X?yɒޠx��t��+��!(�y��&}"OW�?���?���O�Ҁ@�u�u��>Z00�y��'F�y
� ܵ%��'H@�RcȖ>B�(� C�'��"=�C�>+�,���i�$��1��i�e����?)��r�B��wL�=�?A��?��0d�N�>0�=;b.�%�äTMx�!��)!�� n�%>��虤O�T�3�I2R�.����j��i�V�Ҡ
_���f�$b	(<�ezt�U��(�'��Հq3O���� !q�%��+I�4<�!�Ox�'C us�S��0�I��и5��R���ҕvP�	�ONx����i��g�j� ���B0xy�QC��3?�B�iQ�7:�4���I�<�pvrar�%��tKU�$Fbq0&]��?!���?a�Us���O��$v>�6' +gc�p�����xK��Tgx�0
U���j0Ip�*��S��x�̙R�-pqj^�� (A@��0*�y"�W�4mqS��(x���I�_m�J��m����"��[��Ԃ`&��?�!�i�b7�6�����O�~0M<A]�7	a��hi	�'��*,�g$��VeڍX����y�
�>,Of����U˦!�I��tZG�T�Tv�qy�kY�B�|ҵ`A���	0ьu��䟴Χ}�b��%+v��F�L�uڎ)㔹wD4ܪG'Zw�!Oz��C�ޢh��8�2B�1��y1���5��9%C�U����@�p<��t��Gy��@��A!��U���A��y��'�2���!;��ؙ��(�Dqs֡Z9�VC�	��M�S���X�
�MSQQ��d��<1,Oj�"Bh�Ҧ��I�D�O	����'������>[9����2i2��
��',�� TꝢ5�6 �j���"Y"[@"�S��)^3�6k��s-S8"2�XCr.��gv�'�����,}�hP�e"]H���'Q!�R�[?0g&lsc�ȍ?�ry1�e$}҆^��?���3�O4�O�X�nάD[�\k^ft� ��yr�'z�'��I֟��O�N�D�]�(�l1�[�0�Ó��F)j�b��[�E�	9K} $)�	��&��'���"���4�?!��?ŭ � 4(���?	���?�;U�.T ӄ^�VaL�o@�&)�0!0���GIb��x�� ���V��'{�؋����8qbď<3i�L3�@�� 9`��
7$����!F$(r؃���|J��A��j��e��(Pm�
�����_
3�\4�	��MC�a���#��	֒?���p�A�tSTlR�+�
��q[�ʛ��hO$�zp�m܀	�d,�C��-����<��H���x���$\U��?��O�N��,�8u�kA%�30�8�֡C�Q�L�J��'J��'�b����џ��	�*Ě�ن�ϷS�I�F�A�@c��ÀmV_:��:)]�kxXd#'@�';�����C/[L����"� �a�R��>:�zH��f�dXR���!��v�蛈�Z46!�/�9cL�XXC1(��p��џ�B�4T���'8�	���?���^6REFE3��]=Cy�5�Ш]���=�G�^'{�|���d��0BK�����0Jt�iz�'6�����\6�A6#P�T�1x�B��'�C�	2	�\Q�+�q����#J+k�xC�I
s$v)�%ȷmE`yH�6C�ɂ�,���(� ;�>e�!�E�	&C�	828��%����L��YSm�B�I+P�@��K�0���Ue٩<P�B�I�3����&A�K�B\sUJ\�B�I��P��Éu���AmH�I�B�I�[g�c�M�Z���yC���K�FC�I.V���9TG�.���ۣ��0O0C�ɣP���,X#,T��7���jB�	1�V��E R� �^.7^B�	 n
�9��T�L.X X2�^9v�B�	�`J�yP�j��y��Cץii�C�ɈBՀ�j��G&4��$"ƪ�'[��C䉻8�PDyc)�=	�>`v`�z�C�	�&�D�P�� D� ���a�X��C�3�N�Q�+\�gQ��?12B�I�m�V�	�c�(p���@c2�B�ɬ���EJV���ؐ	�V��B�I�Bt@�v[�1¼�;`��(d|B��g�Y�#+�J2L��-��R�TB�I�3T��%4Ra�����E��B�4^6�$��?hY��MK���'��U,��-$��4΅v��h�
�'xV$ wcJ'5Z�)2!&]/�r5�	�'D ��o0�h��M��c,��')���O�,����5/��H���� T���	�%�@͡�=X�|�"Or��7I��bQ�L��"�@ �"O� a��0�1��T�̔f"O6�rE-άv⶝Sf��3]z�*��'g����\�^-
5��i��`���9<'d�Ŏ #3:1J�'K
��c* �,�!,NedDӍy"$^3W�dEѱ� �{&2 F�d��vl�k��(nD ���/�y��}X*��������."M�Pڃ��:x����NPtG��O|+MD0�CX._^�"O��[2g-?��h�*U&|��E�e�K�e���e�(Rd�דOff�a��ˉt<���'\�>>�ȇ�ID���&V?_��|07�O�s�CT�)5>���(�J7pC�	C��
 ��-).]y0�ʘ����ڣY���,�x8`G �(����[9� H %�	'4��8�"O�%����#�d*a� �7�릀M�n�@�9��]��~�(N���I2	�V�jaG��\�ezd��AC�ɻG���Xq���  �[Vg�$ȽyP��U�J)
4	P�%��z�M[48\K�{N�I�`�93�<��g�%x�Č�.�v}��3�═�
��'�Ԩ˅���	HB�	>�"�`kAnF^%P�Ň� c�$R�է_J ��W")60Q>9�GE)Dch��T�;��]��)D����V:a�H�S���Y��p'i�(m`��D��č��(�剟;/D��!n�C�5�=�PB�IT�
�j��H+0�$ɐ��q�N�I���� �'�(���)�T�#3g�{R	�y�$�ڗ���� �	�61��rD��+u5>AP�3}�\�jj|���CG����s�pM���E?d1���D-B���;ҭ5��H'#�����`n�=I�%@#G�41���n݁~&�9	�D�$pP��?(m��c��s�'���
t��<�;Y<�}b�*Ӂ)�Ľ[��w�*���c��`�v*�a����O^�H�x%����GN���Dˉ|��`��t�
6��17�ʪ*Ut��L���O*٢R�̐�M��cM�%z|7�J<$�`(
�FS�(x�+��А�S�y2���'꠳f��)M�џ0�+��n)�@Cr��&7	ļ(���>I�
�s$4�K$�U�t�ӑ�TWy�gy��Ł=���R+��q������C�Z���.�O�3��Z�#8mq�F�f�`R�mP3*��:�c�vy�Aɶ����4h�)��N�
f �E��/)�h,�CH��a"��
&����
ҺEO�
c�՞<>���LD�1* �Y�,��p�X�	%���'FX���� yy�`�3�K̂�Gc��7I���O��#2HH� ��=�@��	R�DP��ia 0��뜠\H��Vʍ�<h�,(>�a���[(<�d�����/ց2� ���䃿S�ҁ�'1�[�g���h��9�zP�+O�������"XP�瓾 M��)�k�
�(Q��	,	&q*�.�x�'�[+s�F��$i�2�Lx-O���gܓ��d mӔ�ۄP��Es�lƖnRj��DZ-@Z�%�@�_��"����?�`���O$P�u���I d��O,���� �'�"�����4�l�2�4b�ʊ�$�~��-�qo�(<X^ъ#����Q-�b��Qi�l�4Sp"�*}�x���?�=OPܪU?5!��Fd�H�'o�E�2CťVH�3�G�U"5K<yc���E*D-h4h�f����0��O)�Ui�0nD$X\�Z���g��U�4��&�~�'��,|�<P���F�'��i[�T!jD���;��|e���1��B�V48Q���D�Zn�$����j�M� �ӹs����P�ll,��	�	�A��@����Ճ	Q$��'@��ɟ�>��X��$�gW�"���6��=fM6SC�R�*��'J´A�%_�<y Ċ,,&��1(O��àĔ1A�X�F�7G�A{��@P}W�p��8`	�&F`Qf :,��X�лcV�<cd(柼+&��y���ġԩk6�����"Й���'�J���n�?��P�O�mʢ�T�Q���4@��%I,���ֶ��%�=,�DiY�Ț9Q�lȦ�$��/X@<Bdn��x�(����L�a~���e:B񳰩��t�|���nN:`<�i�Ck[�xH��_L�'n�u��ӻ&��𲲭��#��@� ����z
G3����D�&Q�9��ݻpx�J �ϱ5�.�#G��r0 XS�ܫg<�h���	/~����b����dE��2/�'��A�nR	��t'd��O1<a�O֑�6J���x�$�^7c��L�&i�c�M��!�,�h���j0��W#ȧ{_5�5bT��Zl�K�=��}��A#�F&��?M�S��6� : �χ,���!�Ƥ���n� �~��z��M�W�p�'�"pҨ��e���ጜ@O�\�B'2�ɳ~���|��BN� �T���� `��x2��
y���10'W�j�����)d@T��ƞ�y9�UY�ܾ6N\��L�;/�4l+�^���i��4�K]�Hy�m��-����#�ON�:��> �ajR���,�W����Wcj�*q��=�@A�Ь�p��idT�C��Ĭ?�����F\]�������tb�� �g�r*�">��Ŏ
4d�=p��R��򐁇A}b呋$؜��#���L�Y�fO:��~n��/B2Xp i�I>:L
��'��h�&,�e���R��8�^RhӁx�Ĺ�dZ�jU�����������Y��Q"ƭ<ifKŶ�Ny�DZ�JH!�@c�Q؟�1�Ć�-W�8�6�D_T�� �\�4�rŚSy`���k��:}Zwr���qY� ��z�4� W�ԩS�Ѻ5&;���!�����	��MC��Q�D�$Da�!�%`)f��qfT�$HH�̺���`(џ8�%dˇ,���Z�iQ'o�Z��>9��*�9{O�|�.O�'a�.2faZ.T�N��6+1��q�� #����DţX	0�E	&(<0z��
4B�����T~b��<a��)?�3���V�>t�IěP)t���&	w�<QC�ޓ-&�`�%�=�����r�I.r�Ј���)�K��)9e�� l�A˺l�!�< ������<,y��h\�@�J�`@0&X�����.�xڰf��)Ɋ��F���|@�ēa����<Kтᠣ/��qBF�+��8�N��dH>.Lt��X���elG	W�y��-E�1O��9A�5>�y��֯����"OXm��2z��-�tLZ7�R}
"O�-*V"ޞF����+�|��L(�"O2an��+�H����u�XAa"O��)`!�N��x��,9'���"O����f��jCtŻ�l�p�@�"O�5SɔaQ�S��W"�C�"OB����Y�!�z�zp�NN���"OX�D���FMH�Cf�%N~��w"OfT��ۚ�H�HcdE
B���"O�r�`\�BZ��5#Ƞ(�1��"O4��)�93�}
UD�b�D�Z�"O�|����f0ճ@�[�=׈AB"Oָ3�!Q�.�z��A	�8z���"O�xkD������#�>\�"Ot)v�6X���*'�G3�H|cd"O�e�	O����Yf����"O�ԩ�k�R�^U
'�т��8�0"OB!@T��~2 ��ŝ!���"O�L�ҩ��xl�P�E �"O�\��j�w'�4{�Ҿn��5��"O�<�t�+rl��(S	�<?���"O�M�c�ު6�`hp��ΰJ�2܂t"O��#�Z7�<�ؕ"�cz`�#�"O,kD Ʃj�҄�b�:s�LX&"O�!Ґ��K_60aU#.a�� '"O~��m�h�T 0O�`Wؔ�G"OĕhT̙�cC�ɩ�E!4LJ"Of`YqIM$d�D�����G��yq"O�L��A��`��	֥y��l��"O��Ñ3�$W8K�B��a׎�yBo�R�D��)7���E�B�y�㔆m x��9W|�I��E�yR�O���-���P�TC��y�Fc�T|��m��!
(R��O�y����+T j�B�
�Y�fʃ��ybb՛b�&d�R�I��̨��ו�y�m�)���xd�4
����1�y����.��y�nױ{����i2�yҀG�$���ŗ�x�|�����-�y2b+#]�lR��;q݌���g��y��@	[:��j#��*c�@9�Ga���yR�,$���z� �����ǁ>�y
� �	���	r=v@��K5�a �"O�l���>�h\R� �:GPM1"O�@���;��]�n�G�)c�"O��x��9k܄���V�{3e��"O
@���e�@�NZ���"O��1�1	�vl�+��c��)�"O�,��ʾ-/��I �?>��c"O�-1G)��fV�٠��I��1ڦ"O$53�HO����I�f��jwN�f"O�pZ��>�9�1f:��"O��҄Ұ�*�Z��<NԤ0�"O2�篑�W 6�A��ͮb\�� "O֥	�h��]�L%
K=vN��2�"OP�b���?F֤���'��o�y�`"OhD�īW��y�uFEh&*�
"O��9�B׫e�쩘�%�_�r��"O*��C�2y�ڤJ�!d�v陁"O(�A�D�v9n�E�	^�n��"ON�'�1
�
��h��O�p$�"O�-1���H� �΋r2�]��"O\B�� X��� d��C*�� "O.y���5y������6�2�U"O�P{����(0pQ:G.HZ��"O�����r~B=��M�6HԤP"OJ5�	ڕNN�}#�Bӷ^Ԝ�Y�"OTUjƣ�&��8(Ǣɭl�H�	v"Or����lN⌺��+���"�"O�PC��#m ����W9*�����"Oh �3�M(~Є����� ��"O��趩	$���,?�ɫa"O�$c��!nT��1�KG.p��ɃQ"Ott�G�9q������5g��2#"OƤ6'	�_q<�����f_�tH�"OH���<r��Q(���, V��5"O&u��d��Z��e��(.Dr4��"OJ��0�]
{�h�Yh�� >�Щ�"OR�yF����x���GH$&�(���"OT�娎�Iz��i�+�"O�=2��I٨�(ү@��H�"O� ��fԓ��t�5{����"O�|��o$b�d��$�St�Y�C"O��O�J��t�O�./Xl�"O��b���zФ��G3Kj�HPC"O(	`�1xB�}Ȣ���m|���2"O���2��.�
Ҷ/Q���K%"O�ECSG��s1��*T:A{�ȣq"OX� a��89`���#�cĴ���"O���'�Ðe�8E�B�êH΄Ř"O6����A�\M.Y�!ȞO��Y9�"O@1�'�+'��5{��Y�P3�)w"O�A�WN��[�6��T�L�F�P���"O��7�,<�l`N;(���g"O�8q��R&h�|1���[�Zmr�"O����d	��d�fKP�hse�"OTi	�p�d�ĝ�%Z�YX�"O1��m�!�6fI�vA��"O���u��;��e�T�0%Av��V"O��dØ$9��y�3M��܄��"O~�Z�	F��t8�A�^
>�\8k�"O�0	K�FȺXC"���{4���U"O60�b	�6I�0��"��	/V]��"O>XPw����6Z�p��P�,�6ŅȓC��`��X����p�釪V�<�ȓf+�:1��	;�2���(å5v���S�? �ݺ��6p���A>3<���"O2%�f ә
�X�K�/�+���*C"Oh��� �I*�I�k��d�N�[s"O��@�ʆ�5�V�k +��Lm{A"O�i�f��
�����  � ��v"O�L(�R �����5y쐙�"O��+s@����f
�S� ��"O�*�,��f�j%+�S�T����"O�ap���<_�(�I%	� Y(��U"Oy#ّW��a�rM.�9�g"O��@�I'�Դ�Pb@�:x��"O>��R,�2&L�� F<�H�"ONe'�ٓ?F�9��..8�E"O��H�Plu���o)|���"Ot��@)��>��� 1�PK"O�5xo:�8i8�	��r�Ty""O��y���	~�m�NH�h�6�S"O�QZ0fE.>�ش����,�&�J�"O���_h�1[��5���!��	T8��($K�28�]�C��2jFd�w�4D�8�C֙w� e�P��6Z`HQN2D���M�Hx(X��* 1�B�i�%D���B��4?O�I)s��l���BG>D�@2c�2��MsP�_�7&���c?O$"=i��׮�^���۹
�F��7��z�<�� �~-z<�7@80(� 0��M�<��վ��1�A�3l�	)Hc�<�錵$
\Y�: �2�(�h�F�<y��RkL�[#�f*�`D^h�<�a�}��u�i�0e��[��C�I�.4�a�R�Ƚa7�q�`/�"3h$B�I�lB-���d9�p@�4AZB�I�c���HM�.9!ǆ-p�����$ғ<�	ړ���}k`=�U�ۀ��؆ȓf��;$�:k� 2����ed��Z�),��"�D��w��?%�n���_�
 ��(}0�����_�3mֵ�ȓ}\���">�n�H�	��L�,T�ȓf�����]VI�� [<eD=��K�t��Vm�r�i9�i/�LΓ�hO?�3݁G�4�97��>3�^Q���1D�$ʶm��pB�H9U!J���2D����e�>��H�E�H�
.�9��.D�Tz�!LoA	��|��#�9D�4ÄE@�~ٔ�S5��<n�ش	5�5D�8ᥠL"d��$+�@�=L7���!*O �f�B�E�lr��tW�"O��8�mO`����5?�	�"Op;!K�%ٸ@h�Ā;��$�mH<1A�;?ӼU@�%�
7�m�&��u�<	���b�V�ە�Ê,nl@F-[�<aq��4vм���B�13T�bB�T�<�k��i�=q���<�䘊P�N�<W¡,󨅱5��#�$�jcMI�<�t,�qߐ�g�kN�"e�-��xbКl�T�#���ት-���y�l@ل,��fX� �d�:fhL��y�?f����]!u.��"6�G/�(O���dނ|�B�Ȓ���aӂL���Z�V�!��΀/`*m��(��i+�����9p�!�N;%��	���۟0�@�0sT���d� ��<�J<a��~sz��rϋ�Pp"$��C�L'��"m_�'�m�C��b��I�h?D�2�Lfˀȁ���#:�<��A#D�� 4\���4z{��
SJU�V��`�D"O&��[+g� 	V�^�9�Ι0B�	u����눼X��Q��9:�Mâ�8D���%�9��Ě�#Y�ؠ�G�6D�D� g�1�`�P`Xy� �!D�h sNǴ�L� ��ô}a� D�I��F�V躔n���Y��g,D��B�O\6F�D
��֔��!��+D�(�O� MAnp����E��i�!I4D� K��ƒX��h8��n��y����t���d�<A}켛�
�1=!їm(AJ�y2ቒ@Cʙx��7f�<s�K�0�tB�I�U���+cmU9%���3�H�0��B�I�� t׫!�esC�0&�B�I?R����T�L�6�������B�	.]��]c(�M�~`�N^��LC�I�{��i���*=rLP���J�HC���Ȣ%k��'1�U��P�
C�I,?� ���ƚ�$���&�-�B�I�u7(D9qD*������/*�B�	Zb�W�Ԃid�Z�Z�C
�B�I��
x;�	Wn,, E������'�2|�� B�[5<�a`�==��i�'�jl!�KB�s t�!�);7j��'���C�S��p1��*0}J K
�'K��ТG�+
f�ڔ	�(�b)�	�'Gr�)�X�=aNG�4�r�	�'���cQg<�!�e�� �P �'ʐT0w�\�uJ0�;�B��0��
�'k*9"W'��u�-ӄ�^0G���'LB�j����,�)O�b��'�|-	�jD	Axl�����a��'2�;��Z�(aCX!U��"�'W���M�k�5��K��!x�'�5���֗(I�ҋ��!
�'�$US�kL/��1��Ǒ&�����'.z�:g�
[��� l˞�5H�'�6jg̈́-p��x�c��69��'��X((ݏ��A��H��*d��'�$,c I��V�H�Ω��Q�'��
ǣ޹L��A��T#w��R�'�XX��j�?���4 A�qJ��;�'�4*φ�$B�ϓ�Y?&���'N�@f���s��䀄��)�N���'0Jİq�S� �n ���ߓl `%��'�Xr-�4r�6�j�.��_<n���'l~0%�2(��u��k?Y��q�'�d��� ��fC�m���"<�޵8�'���)ub�4z���̩2�|�x�'�f�éK�M���a
ي! 
=D�|0�͍(���k�"�;)��D�/D����H�%y8蓐����J3Z/�B�	�i�i�٤-3�I%���f`�B�ɯ[C=b��m��S�g׸?ǐB�>}�1��&�$7�٢F��C�NC䉺D� ���!A��Xyp�	�+�C䉢y���_�uX��bӖks>C�IP`���ÈQ%H��G�y�C�I�֐��o�,B�b��a��#u��C�=OR�a�eE��=�\�`�+��C䉤0�"�R򇂟1<U)ҩ�o�B�l�stJG<jl*��Č4"gJB�	ܴ�B���f��LadC��/*�C��W��X*��X!K4�y���i��C�)� �$��D�*Pe1�N	��(�P�"O0��E�12a���*}ז|H5"O��c�+T�>���b'R��4�"On��F�H)�QРe�#�:�"Oԡ���E�:X$\R��'{�@�+"O�% ���C��i0�O��p�"O�)�0hғJ�J�"&�`�z�q�"OP��k��9�\�	V��$K���y�"O0�8"O�.8Q�bNńG "���"O��	ҤH#F�����=-�@:'"O���h	Mp� ��\�Z�� "Ob�"c�G"�nxX���@Ā�k�"O�XrBO�w���ss����U*"O�9@��,Tp6u���,��+�"Orh@��iz\�1�@��v,Z��"O���b�H����@o�=�ܹ�T"O8���O����O��q��0"O��#臁��l�%-;;��٨0"O�!Ц�F;1��y�ƅ,T��"O���p��=_a\�+�A�7�H��"Oz4����*��26O��y����"O���RTr�9�L���Z��"O�#b��BL�h�*�E�n��e"O�	���r��Ukw��g~����"O$ ����P�Ѓ�!ɬIj2qXW"OV���DǪv\�Y�拺��1�b"O2�1�J[�h˰a�����*a�0"O�$ef�`; �R��4\��P "O��{��|,�(�O? @Z6"O�a(�J�3m�hV�ɤR+�%��"O��p���;2HR����Ⱥa.j� �"O��孂�P�zd���\���"Ov���L�%�\�ҥi�Q&qx"O�X�-��f�z,�Pgܻ���J�"O�<:��|��x��&qJ>rD"O��q3��X*B��T$�P���"O�:��:5��D�����ʐ;R"O�ݲ2�W+IP����0ly"�!"O�=�(^	e��i4^�)?���"Of��k�kU�(�f��."�P�"O��Ƙ�e.^e[4T	2ȓ"O�	1��a��X���~�&�p"O&1[�V����3Ǎ%�j��0"OJi�NLƅ�r㞸?�j�r�"O5qb�m ��Z��є/$01�"Oqb�9b�4\bV"��t�)6"O$%�"(�O��tڀ*@�L����V"O<y�eN�,l4�c�Ͷ��� "O��K.��@�0
�A�i �"Obx"䙷r\�\�U��g'z%"O��31F�Hu���Gϰ>X�y���1Ch�I� K	/��H�q�E>�y�`߆_В��Ґ5nz��ӄ��y�	�'� !u/��*�Tx₌P'�y®P�>����n�n� �"*S��y���\�&��/-*�s��¸�y�B��,;�5��)	2l��Z�U��y��&cW�
���&�V�R" V��yB�Y��`!��
P����"�yr�ܥ'D���֎o����Ñ��yg L�z�[��,��l�#��9�yD�.�r|��?k.�����y"	�P�D���j^$_+���ћ�y����o�x9$�M�Y�Z5j2��y
� �D��NC�{��P�Ui[�3ȋp"OJP��&��f�L4H�N�P@Ց�"OJH���W)Q�a�EnE�yC�H#"O��j���=c�H �t�ٚa�j�p"OZ�����6�r�PC�.jr��2"Ofi���2�*@�9XU�ׁQ!��5����$ʨk��R&�	�-�!�W�%h���C�:9��RdW?h=!���h�2��p���KԢڽ6�!��4L����&�9%`)��"�6}!��O?u">pXƆ h*���N>_H!���n舱��hU/0�4���)��g�!�_e��ML���[�ɋ�Yl!��ť-��ʆI�I��� �IϐX�!��+92�#�G72p�E�i��@�!򤐂?Lsso;f����!��ǣ88�D�Y'v�pB@��!�d;_�0h�'��*�ɒѣ�&V!��	�_v�����m�`P�\7!�D
M�e���*(hj:�ˑV&!�d�}8n���X�����D!�ɸf&�av
�:�0��S6!�*|p����ܒK |Р]�L!�T�#�r��$��>��	�U*!�d�33�$IW	ɬe��HCH�> !�$~���HW�
����v&�*U�!�%^�|�%*H  �%6f��+�!���+h���&+D�j���!Q��
K{!���w�E��:czP1��eN�q	!�$@ 9۠�9�$U�Zw2�X!�$�9f�(ѩ��Ŝʎh0�;+R!���:S'zJb]�v��농��:<!���t�L��)�0Pǒ0�4M�8(!�[�L/��SS��__r\���!�$D���MR �0#VD�
b�M�1�!�dJ)GÆ�1��:���e,
=c�!��8Y�8`�I�$����Ҙ�!�d��ak@mv)��e�����ӆ-�!��ņ��:&L"z�TX�Q�!���>i��1���(F�]�c��'!����i�r�"��LDl����:�!�DS5T�X�V�MPʬc� A1�!�T��`E�ukܽh9%�a���mC!򄐤7Ķ�b�δW��E�ˈ�a!�T/=U���v�H�	�6��#Μ~!�ߛ^���1�/zu�B!�?�!�dF2D���ۦ��&-;�ٳ1���;!��J��&	Ta4x���E�]H!�DV?�r�!!!S�j=t<� C�,>!� �I�mAv�Ӂ��B��4!���!��SZ��[����n,�"O
�C�.͢|�`1��*$��1�"O��Q�*-)rq��x�,�3"O�Es���p`v.ؕ�x%R�"O���a�!k"IQS�Q2Q�
�(�"O4�9��ÉJ��i+��:~�t�T"O�ٻQ��U�^E�r#"���03"O����e�-]�"9+���<�|g"OtI�+�άh@��9��,��"OF�b狏�8[
�ReV�v��m�"O��;�#�ƈ�r�V�����D"O���5$p��b�)c��$�"O��CsGQ�`� ;�*��M�<�h�"O���A��<�<��T/��+p����"O� �D�RK�.G���#�،R^(�y2"Ot�q���3#����Ζ'�&=
�"O�Ś�����Rq�НR"O�}#���/u6eyH�_�e!"OZ��3�Q���f��]�у�"O6���12��|b��(U�k�"O��Β[�UHţZ�)@b�Hg"O6Qa��
1��8�#L��f'ʼP"O^��! <.��@�AI6T�YR"Ob�6M>��X��Fz��x��"O�)�2l_
 �� �	X�ȝ�"O�D��"�j�BՇ�j�"O�\��)Pp� ����H�@x�"O�E3��F/C P�"�Q
��Ոa"O���%G�O=䠒c�|�P "O�՛v銿^ఙ�"�'�%��y�by��ePC����MsU�R�yb�σXT�xP�1����%���y��é[��Ƀ�:Gk��yr��Y���#N��
Q����yBE6-�LƝ{��A�g��"�y�
�f���P��q�� �'ǝ��yb�@,V�N�)�*X	f�Z�I���y�&V|�A8��O6(>Xp�&nI7�yBLS�:�['B��#�6��cA� �y2��N��֋��3���r%5�y��������G�����C��y�R'?�xq� ��.���ҁ��y�ª�|�s�GM�C�n��쟾�yeH ؐ�K1���q�B��y"%�&U���jT눭,3��8��;�y�*��n���Ȏ�DAP�H(�y��H4K�H,2�'
>��pF���y�F^��c ���;� ����M�yb/��T�`����7���[�O��yd�9�b��A�&1?*xy�$J��yr�[�b�*ULH(��}�欟��y�WD�\b�D^'j�<��3�
��yb�
6���E�^b%v�
$��+�y��ykb�h%']&M�����%���y2BĦժ1��Ao�(�	WM���y���7QEPqk���(g�&hYv䝜�y���,�<1;l�-3��� �c���y�j 5{�2<���˟)4p�F-ʁ�yBȟ�CJ���#�M�#�@�����y���օ�G�<�:���'��yR&�#�	���N!�� �,)�y�	Pb��벪=I��5P����y�Ț)׎(r�%J�z��q��y�Iۚ;O^�{�ΈS�.d�!N��y�	E.k�@1�d�R.OWε�����y��YQ>0)bb�:2��ːH>�yBj�67.q@O��PH�-E�y2�ѐ%NȠs�/Q)2t%�ʄ<�y���<-�� qL۟Pt��̗&�y�.�U�@�1��y�����ɵOX!�$�>)6��a�R����Z���U�<	���.+*>��$ L!���FR�<��,JE�P�߲|kx����R�<EHԉA����B�9��@dM�<i�j@�rz�4�D藢Nr����K�<) ��4򣣚!/_~��Q��~�<Y�+U.xG�#�ɛ�{��(PQ�<9b��fn.����Ҽ���K�<� \(C�B'f% �	��ݑ,��T"O �Qiן6�0]��nC'b�nܢ�"O������}٪\r�]�� ��b"OH�c��AJY��
E3�����"O��X��x6E�P�V�Z{�H !"O�˖̬+�zx`�ٱ}���+v"Ol��M�?,�yz�*�I�Luk�"O�e��H�)���a�
ӓZ��%�"O��H�ᑦQz�)�c�#"�0R"ORe#���3E�%� %�"{D��"O�I�R9o�$,�BD���D�W"O�[��lGN	��E���@K�"O<Ը�݈Bh�{wd�� va�Q"O tf�YG�-���^��*�"O���d�?J�Ա�+�� �"OܑY���+�.�p���l�CD"O�9�PɊI����E.�%�F�y��P-.C)\�2�f健GV�y2��6%�(��2&����Ë�y¯Λg�29�IC�"�F���hŴ�ybbD4I
<�Uo����g�Z��yI§x�%�2Dp�X0�@��y*Օ=ɬ�do�	Q����J��y2(�	.��t��N�#T�\4�"�y"ɏ-L݀!�r�~)�6.��nx�ȓeϜ1P��A�~+�d�G���h��ȓr*�2��X���!�e�
l�ȓv��9�P��9Fi���Twz4��ȓ\��ThQ'��Eg p�d
=o����q[�(Y��^`�ܠ㓙>���ȓf.��gK�	0� �oFh,L��v�<ш�\!X�H�H&�#�}��}��'bM5 9�PH�Lcg�a��4I��1(��(��ɢ��@�Ե��_҂��S�Y6�J�ܼ^,� ��p����Z#q���8�@�:)ΞM��s�ِ�V2g+D� �*ʷ@!х��fa����0R1�b�2\�����5�l`�lj���ꀌT/d�f|�ȓ�l��f'�
`)� [C������Ӫ�"��<KJ�P��C�x4(u"O�Y`��Ӏg��D�aޜ�چ"Oք1ԉS�Y)����H�-\�T��"O��K�|QHР6�L�Q���k�"Oҕ�v%�u�|$RG��� z�"O���2�P9�0aq礁�b��37"O�E��	ҤV�
�z`�G�T�t`�7"ONd��bݝi`��Bb��>����"Om`��4krP"���/\����E"O.�4���D(� p���
�"OT�a�FF�&�X�!G�ɠ��M�f"O�\#�L�+'�b�H���w��3�"O�2�b@<�f�6��M�#�"OT�hՅ��f��١����Xµ��"OLK�A�Q+��ٵ��[t�6"O�婶D�:x,r�����0`u�g"Od��:.�)`�@�>���"O4�$�K�T \�9�v�P�K!�dΔ~`�i��T�J��\ۤm�3j !�$��>�B�����l��Y!��	j����%�ʧ��)�ǮF�s�!�d�6W]� ���3��,��� v!�$�!}��a� �:M�J��  r!��Ж��e3#��zd��R�@>X!�� �� ��,&Թq(�  '�a
u"O�����њ+�Z�� T:
����"O���U�v�F���n��`i��{�"O��'d�C�"�'ȇ4`��e*�"O����YH�U���<�,��"Ol����R�`��A���G�~T!�"O�,�`B���R�ӠhQ0^�Zu"OX���GK�Q�sh 1;vra�A"OZ�X&$�:z��ؘRj��Je.���"O��!oŀ`st��*^zT��"OZ��A���\E��Y�v����"O����	2Lx��~q6��"O�}c�._�)���!W�KU<�Z�"O ��!�F/$6,��`�i2ّ�"O�IRA��A �L0lX�/�X�B"Oz$Aɝr�ltP�C�QT�"O�MPp�73w�L*AK�9]S�8"OfXȲ �m�1��O8 ��"O 4�H�k��h�3)R�s| �*R"OV �7�_�R��BV�2Ls�@��"O��r��P��H�g�"9bT8�"OP�Rq���Y ��kRDђRF*�ˆ"O(�RO��
ٜ8�U#��xG^��W"O:q ��L57UbR��IA���"OZ�(�	6���
o���E"O8�"RM5H�~=�ߚ�x�"O&-��@ݮ��tc�Pk,���"O ���hʾҔ��O�+�@ ;G"Od�F�(8��%s��_�;�F��"Ohe�ƀ�8Vo8p��{M\�R"O�ء2fV�kp��/Ͻ	=���"O��SͮcN�۳n���X��"O��yw��j�%q!��+��0"O�
EcI�P8�ц+\7��Yڱ"O�03 A��Y�>�����m�a"O^q�*U�.8��φ@��9D"O�����ʀ4�İJ�+~�8%��"O<@9d�Ԍ	L�I����b��R"O���@�R���	�6��;��z�"O���C�6Q��ᨳc�����"O�#c��"=����t����U#"O��8W���a�Ha�m�"O��FI��u�qg�:M���!�"OV�5�u��8� ����Z��"O��R ʒ+�9�L˂vV�J�"OdۆG�'�����l�Kߺ�0"O��L�4�xPp`lŏoȦ�[!"On��3^HT��˼P��!��"OV���Lb��0��;J*�e"O\��`H$�n�Ua�]�eX�"O�4����* H��:� ɏAٖi��"O��J�zJ-b5iǏ}���5"O&<�t�Ձ�<�4b� �T���"O>��J2=V,�A��C�,APU"O��k
n��A����8b�"O$����ޯ�}����R�p�	�'{�}��fû��qX��ʂ6�`���'����E��<�)�`�*��	�'�)؆2��Zs�K�3$��'W�� '@Fe1���	�*/_&�8
�'��H`�)G�r<�%�Ǡ^GԽ	�'��S$E�, �z]�+G
\���	�'�^���ʆ��#�%�z�	�'攩���ӚX��ȕJ�̍�	��� �ٙ��'���ӥ)�$K�\���"O�Up�ы�ܱ��5Ր@K�"Oja���)�$I�Iׁ9Q�d"O�%x�O7:������Zy���x�"O��I�nn����$���B"O$m`Dљ��]b�l��H5-��"O��;��)E?�t`�Lӿ~`h(�"O !H���i\Έ��L�'��qW"O$�9���24�������j�����"Oh��O�(9\nLA����e��#�"O�M���X�n'����ۘR`�|��"ObP�&/yᬽa�0AF��t"O���!���p�Pz$ $?���"OP��Y8��db
�/B�
!b)"!�D��H�2�S��\�)`�ҡW�!��4?*y���;r�eّ�ιU�!�ES�(A�Q`�Ec�ps�Bl!�����;@c܉e{��*G��5i!�D�b��	I'��>a*�c�ٻ&L!�d��=\����Ė�S� -Z'mV+!�d�O�~�#fLg��v�?#�!�d׈?T�)���6_��P;��+b!�D��^��%ڟ2���b���'F�!�_8wIJ8��H�L�؁�f��p�!��h��i1Q7}�F���B�!���PUwM��5�%RU&��H�!�1�v�Br��7m \]ѯXOP!��_� �xAŏʹ{�́�3ɔ�!�DC�+��E��Y�E��}��Z�!��@��pf�(�tT���s~!�$� l �ĢC�V$�� �C�,Z!�����yW�F:#�@aa�O`�!��@���K�z��H� ��S�!�Da�b�{�Ӂn]5�w"�t�!�DJ3��=�d)O��-�%�4�!�d[�7��pSo��.��H�`��>�!�>EH@��3b�|��DjGB� 9�!�F�xVz�����Ff����=\!��Q2l��h�2��BD\���aIy!��T�fq�i��	:♲� ɯ^?!�DC�VY��2G+�0%��3��� !!�ć6FO�]#ꓟ<b�a�*�U!��#?.uSp_�c
�)q+V�@0!򄈣Q�<5��R		6��d�Dx!�DH���#$"
���"��c!�$^�a���� ]	u ��Y��α�!��9�0���X/~�3U�@.3�!򤀍#���fI8<uj���N<P�!�ĉ�*��M0�l�lb�@��
j!�D�9E�X���>����1B�' Z!��
�����FZ�i���q�Y>�!�$g
x�Zi��M�2"֭M�!��	20��5E��_z�%ѳ"ފ�!��ޅ_g0i*_��są��[3m��"OY��X%v`pY���� �y��Ɠ'���u���/���ֆ��y�e>[%� �C��|���?�yRo��d@�""�?���g/��y�����=QS/ߋI�<� �Q��y�e����5HŬR�?DE��ܳ�y"K�7��Prq%�=:S��C�$��y�搎G;�5�Cϕ�<�X�����yr��)ՖH�q�K.v���^��y�IԱx�|0�[)!��=�'��8�y
� ���ǡC�)�Ƃ��Zw"O�	�T��)���0Ga)*�!e"ON$ycm� !WHKf��4@iru"O�@*# A<DcxYI�/ݝp=���5"O̵1�d�%�R�CmU-| (`�"O�d��?ն�2���.����g"O���maW �B���� -�X!�ˬ,h^ݱ'}��պw�	=�!�@�4I��I$�"m����KO��!�d0l��x�%�$v���	��/4!�.�j��l6E���i��.}!�$ͮq ���K0 2�L+��ޙrD!�-T��1ɒB�?�D{¤�'3!��F<
KX�p��'Ԣ��pdJ�5"!���8e�:*�E�;x��pZ���0!��+˦Y�!��3n�r�Z��C0�!�$�bEj0�g��6K�Ԁ��׏F�!�$�yb����>4�����*Q�!�� .���+K+��{��&�!���	$<��F+^�|�]*F	�MD!��+f>�S"薐-بe:��Q$J!�DN8bzL��5
�87�������!�ds�$�!L�dߐ��C�	�C�!��	��ra%I=g�8y�a�×E�!���+@g�]�#��aHv�s����)!�$۹��ܱ���6Z�v��7d� M�!�$R�Z���F��>�i{��Y�&�!�DK�Y皍Y2�D�0?\���k=&@!�d[/�@�C�N�#[L���K��1!�Dӕyr��&bV	uQ��{�!�$+�h���Hv���Ɏ�H�!�$��*�Vl���#rC��J�GS/[z!�ك5hH���e6AW�	0�݉&z!�Q�<8r Zt��+PQ�0�d��~!�d�R��H�1F�+OS΀Sf-X1S�!��,B�B@�i��\!��qMUjS!�d@!B���R+I��T@�i�/p?!��KE�@c2)N8 *B�K��*<!�$\�6�Aq S�eЀ
�0&(!�Đ�&B�)J�M�vTX���&x!�$Rc$R�)U�f�(|��.[V]!�dV�=��,8U�OH&��gn�4,!�5 �.q�B��%��)���[��!�P��Er����(�KN#�!�$L7��� !B��Rv�C�'sy!�d�2(3����Ȭx\�)��c!��U�{�؁(ti��t�v�KCh�!T4!���~
 0g�-�� %�O�^�!���*8�	�M��c�бU!�dЩvPV8�׌I0k��P��N�R�!�$�s8��q"���m"���anK/We!�$7J�p��Ů��t>�*�"է6e!��ۡ=��� ��K�k�TXb�"^�HT!�$A�6,�!{e˪D��7g�7k�JB䉹($��#��6�)0�dە{ �B�-_��(��cP6��Ms  L2P��B�ɪI���#���8sҤp�P)���B�$b�6ujQ��H	rlq�dg�nB�	��,�c$#]�F�i��	,�`B�	�1b�5Ċ�lQ`��� C�*�C�ɘT���!gE&:\�8� �B��'dI��3���A7>lZ��\/,�B�X����$�� ���0)��Є�VJd���o�%����B��,q�X��S�? ��d��,*Ū��d)�w�*a�f"O�3��H�)��<sPB"���ش"O�2aM�
��X`V�c�E�0"O<�0do�%H ��8u�@&hb�IC�"O���)ܿ���Q���"\�� "ObиA)�zh-�D� OT�2�"O�� R�������kG�X>$@�b"Oyh�.m�t��$�yN��I�"O@�7i�(�vsc�۟
-j$If"On]��_���u2����p$d5�4"O| �F	 ����r��.>�|P"O.��V��=��1C5��� �4�7"O���bh�r�zUɰfH��0L	�"O�Х�fh�T�&�)=��M��"Or�H�I�T�l9F��h����"OZ%��%�+w�A�ß�G�����"OH�1��~� 㝼Jpa`2"Or=��b=��hs�T.�N�Z�"O m�pl��uf����U岱3g"Odq�4���7�x�A+`��D�V"Ohٱ ��N�0�@1?���j�"O���g^��r�oC��Nj1"O֡Cá��7V�b�oи|h�"OH1��]�O²�a���j����"O6��%��0qif�Y��C�	IX-z�"O�� L[&{��Y�͎'O8h�"O�$k�Ξ-	X�CH*NLzt"O�6H��`.X;6�#T�sV"O:}JԊ8N�^<Z�bV ,�`@"O�8!���Ĩ�HƀRX�l�"Or}��F�/��ѫ�Ϛ�~:L�Kp"O�['�U�m���Z�͜>&�4��"ON�"���6몹��,0��A�"O<@3�3PP�y��åz^���r"O��k�٪	�f%�`��Pޅp"O��i�M��\��s�P)P� "OF�"B��3쭀3h�A�\@B"Oؽ���C(2�2愗*�|�&"O��U��"\�%[�È6F���HV"O��� �5ZP�9w En�ƥ�"Op�k���u�ҀHU���HH�"O��Z�_�7L�cr��\v�@K�"O���B.��*mD��-��>a�c"O�SF�'��<�ǫE3cl����"O�-X,C�h`!+Q���*�"O�Гl��8��c���L�f�Q"O:���\���x)%��)m�%��"O�A�3��Q�VI�s�^�r�D��"O��r`�T�L��}pb�ݳq�&�a6"O�=x�
}�$ ���6��l0D���VA�R1���WIB>1p�ɀm<D�h ES�~�z�@K�D� -9P�6D��h1lH9z���`^�p�"Q��?D�d�a�bv�M��M���ed=D���D�^'(�\�(ՉX���Pc7D�l�ҫ��*�Ҩy7�H�J�Pq�/D�t�A�8L!�9��0�����j+D����ҩIV�tO�")b�0��.D��+4��x�����Հq��3�n,D�`�h��C�h�0��0U��)D�hS��-2�b1y�����ã&D���I"�i����;:-��*D�T�1�1DH\E�IS(�rU�"D���&��(gnh؄��T�����>D�� e�3���_���7�6vvL�"O�!�a`Ys3d���1,�$ē�"O`QȄ�Xq9�C�K(x�v)""Oj���ΚL҆�t��8����T"O��3B%��?�:��GBVp����"O�]h�޲}$a����$Rl,A�"OԼ�c-
;��H�b�֨0\|I��"O�)�t��n��#�Ҁ����"O�������V�P���ˏ zT�3"O�D��I	�z��A�=�����"O<��GI�fF<\��V4S*��"O>�bCc��h�l˥��6Tr|�w"O�t˅"��٪�D�b5��!"O�PSf�N���)�E�	R��QIg"O�`#@Y��>�)�eZ,yȀ�C�"OV�MI]��a���{"ȡ�""O$��dą�j���Ȅ����(�"OzA W���w�XZ��>�xXy�"OR�d�(���ѕM�[�� �"O�U�rC]8~z���|��l"�"O���Rư9R���K�@[<	�4"O�zG&��B�ƥà�
a%�y�"O���N��d��4H�>��E�"O -!G��|�x4����鲤�"O%� ��n� 4Sw���D�"H*�"O�Ir��wb�[���VƎt�F"O��� ��|������W���A�"O����W!5YL�Z�@�.�LBA"O�$��*9�pp�"[��b���"On�:C�8W�Z g�N��	ۅ"O��Sc��"pQ�slʼ¼�["OP��4��&|���#���I����A"O����@n�,4�4״%�"O&-�W��<.���ޒa���7"O�I�PH� ���bl�g-P9c"OJ<�cg�t�ˑ�YzDpb"O�ea�D���
O�Z���"O��
U���7LH	ve$E�����"O|�*���n�~ ��Eݒ���S�"O`x�ӭm&��S��m�2!��"O�TQ�ύ�R�n��"2��	�q"OV$�� �@Z0|(����xL��"O�)`�!�
?�Z�K�H]g�}:D"O�x��"�v)I�%sU�	�w"O
�C��˅|���u����Cu�<�$l�0AZ���T����GOl�<�@��	z��q�4ń�X��@ �i�<��懓��I� �'�4�S��Z}�<�2�ˏ"L����NA��X[T)�z�<! g�t�sM_�8��(�Eu�<��КSɔ��G���/(~��nr�<AׂR�E� 8���H��W�i�<�7���
�b5����a��<��*e�<&�ѝ#���#���e,Y!�	g�<��ň&_��#�G *��`�Gk�<A�,y���a�>5����)R_�<����q4�85���#S�� ΝS�<�qB�d�Љ!e䀷qeB@H��P�<����1�*1�L��u�wc]I�<IV�Y�� ���$	��~W�!�䄀E�ey���9IZp����j(!�DW=�m�5��G	d02� 	!�ĕ�����v��T95��!�!�9�P��fF�^��P�UlF	�!�� 0�P5`��(l��-�L��4"O<��Bl�4��5xu�H�tT��z�"O�\:�N^%,$��D��:�p�c�"O\�چ�)5����<�^ �w"O.tS0e���D����@j���s�"ON�r�A�i�	Q���-L䠨�"O
ـ$b�Z���H*N�"0"OjH��G� 6�;5�W���t"OȘ��h�MX<�c��=���"O�pz�	\&b@i�`΋&j($)F"O½X�H�(p��pQ� �_�z1"OR��Q̝,W]��gϮr�r$�"O*�R�'��V����1����"OBq��&LMX^��p@�3�F��E"O\���� HvXaO��*1��"O�)��yt2|`bN�6`���P"O��bCH(s��	�6�	"O����78>��2�JY&_���	V"Ob+�'��D�Jg�߂#m�X�"O�<�1U�&����	^6Sf
�k�"O�:��Wk�@ZI�6��|�q"O�X���	Q�RH�P'��j�NݹC"O
fI͹yH�P{�'e�L-��"Ox��v�͌Y���Ď?�̵x�"O�h(�&�V��0�@�� $*�"O�|��,kQj%��z�j��"O�pyc�:6e��#ݽ,��%��"O�%�"$�-!I�=z�Hٜd�iq "O�@YG���P1p�9���6�b%��"O��)Ö�gH�!R#eP�X�P���"O�UP*�F��-9��N`4u�c"O�����8<�����^F|�Je"Op|K�/�� �����֨� "O��Rk�!`{�Tʆ���:ʄ�b"OVt���ވ|& y`��9ݪ$#�"O�sUoS�fLt!Y�\*��lȴ"O�x��
�4:s"|ڥ�O�gʐ}J�"O�\��S�T�X C4�� ���`�"OzI`�k�(j���w*�;v��s�"O�0����.bPW�Q� �I�"O�*p�L/QG W)>>�Ā��"OFT�Aj�F~iQ)�X���"O,M�$�b��`���S6ƶ� "OP���&�1_bF��2��2�z�zW"O�TTn� I�Pv����d"O^P+E��>�֥u�Ư8j�Q"O�	Ǎ���1b��ܽ)�f("O��H�o;P�B�R�h�:�"O <��LO�S�]#6���oF��u"O�S�M��v��I^/*��B"O0݋�L��*�N44��k��-�"O�������> �M�s%A~�8x2"O�pQE �:I=L���#�2g�5B'"Oh�x�CH�K�����ZeVY+""O\�:C]cA@ "�/�r$��`"OD@!@ ��C4ԙ��?f��p"O�E#&ЏRD)��MV�t�L��3"O��k@�(Ψ`d
�:C�a�"O2���a�6��9��h���m`�"O\!�V ��I{F�j�d�1&��Q"O��O"ZT-`7c�-36��e"O�Y95���&UH�( �P�1"O6���*��hH���u�^�wNPXG"O��P(!P��,�¢^�x��;"O� X�C�.�88��	�4��� "OR�1��w�ȘQR&H�R,�"O��Ce��ee 	B����Ye��Z�"O�ت��M�)6}�V��F	��y���Be
�3#��p����yr.E�?vNDI6FP!#<�"t�D��y��3Z�`X!��Li4���s�ݨ�yR�Y ts��c�|$���O��y���7T��Pӡ���2I�X�4L^#�yR$�&��p�Qn�*A��J��y��A�V�B�F�9'D*�r�@�y�2>��6�C�pBd�`�G�yR*ڕ<�0��W�Z�Töl�$�@+�y"��r&Хc��ߏI�:�k�y��?i|��i���󖌄k�o��y���8$�|����P�����UIT�yr�E�1[6!{%ϋ~V�թ��'�yrC�#	Xy�7hN~L����y�hӃ']t�c�,?|�t�b�#���yB/��n�0�sR�Cs�ȹ�y"i�%���kE�k$�pu���y�L�L��u"�:\�д�����y���4v��i��d,��)��yR�R3�����W�y����`��y/W�0�y�B:f%ْc	��y�+O+J���r�F�3J.4�7� ��y���_�V����$k�)jWnǪ�y2�ٝO�e���Ԑ5���u�A�y"'���TŘf��."ЄRE%��yR�W��;k�p2�-�(R�y2c�	BX��J�D�r-x���Ҧ�y��#��)9�� iN΄i������E6b,�p�D,S&8å�N-*^���ȓ_�v0I&�ģ\	�;�aJ(0.0�ȓ^X�-Ӷ�y\�j2 Ϩ)�|�ȓ:�"�&�rCz`���6L���R
�'�(l��f 	R�xKU-
+4�\܄�?�{P
K�e�����?@.��ȓY��E��75u�d��C�pT8���(�t�ʕO��HXU��$�*a�ȓ{� �0���ݤi����b�ZЇ�qۊ3$
H8+t��£l��,��.�p��- 2~*9�0ɌL\l�ȓ2p��a�q1hDZ$J�<؆ȓO:`p�w0W�2)�&�.jm،��]
b�{K���Aԡ�(p88Ň�lX�K'�W:��Q�;l X]��O,�Y0㈙k����MF�s��i�ȓ��%A�N
R���e
�N�Q��w���򴥃��I����<;�x��q�,�Q�C.6-ڥ�"E�9:��ȓ'%b�br+L,�v����U?
-�ȓ5��24b�#��e#TF^
&���k���@�;q["��7��E�Ňȓ D�l93��E�1�ө�?/��gyހ@��"����K�?$��Ȅȓ0��}H������'�L�vR�a�ȓo��ȑ*�?���U�O�9rԆ�>�����$`x�e��Ε'#ɰ���V"���M�)�JM����+2d��ȓ9�dti���w��Aq��QԠ�ȓdJA;R��I�����֙3&�ȓU�@�3C�7U� eK���X��ȓ.����!CA�y�J��f�J�9Pbu��S�?  ���Y/D�DIk&�ʥ ���"O�a!#'Z.J-��'�5t�RE"O����hֶX0f�:Rr��Q"O�@��HG�wO��y�
.vL4ȃ�"O����z������Y8M� ��"O 4!�+I�Z������V�s�"O���3MZ�3�2��q�h���"OFdi��[��83 �,D�n5�P"OX} �+ƶB	|h8�B0�N�0�"O���` �����`����tx��"O��*�� �
�U����1(�Pi6"O�Y�Nϯ8X c�|�<�"O@5 �-A�u�4�^-�tp� "O��B�1)�8��$̏B����W"O�9�5mִrk�4Xb�D�SNa�G"O\t��(	�{�"�	b_��`#"O��hB!J9�j����=r��7"Ov�X��% ���4g^�{4Ȣ"Oԕ�G"ZjX����f�E`�"Ol;� �[��[ԃC	�4U�'"Oj��p�ȼy�� �o�0�&��"O�%����4�̒�>�|�"O8P7�TK�5�c�G`��0S"O��A�)U�z|��Qڸ�"OZ�� ۫G�D]` �
~��@�V"OpiCBL�d^ ��<e����"O��3�n5@o��"`��HXN-�"OF�����;�Z�����(L�`s"O�}b�h������W&�8w"O���� C]��g��5�pEK�"Odth����E�T�L�q�P���"O(�+[�8	�C$�% �"�s�"O��:slH�[6 �&��;�f��3"O !�R�ޮ[�$l ���R�L���"O��j���$@��.��,�1��"O&䐠��1j���T06h�c�"OzȪSE@�u�b�brA��^̸T��"O:�Bw�'Vl�AÀ�&-dZDY�"O轣'�ȗFDsd	֭s���
�"OT�s�	N �&3W�I�.L$�2�"O�U��`
�vi�@�ń>b�@�ږ"On	�w��9)9�ѐ&B N�9�u"OD�c5�]�V�T��|���"O�����"d�lܣG!U8$YΤ�f"OH�x��%(,��z�)Ȼ%m�`:�"O����ױXJ��"�)7�I�"Obp�EjݺU0�)&"� X�u��"O.m��!�;�&X�� L>Ť	�"Op�� ��e���Y�����4�q"O�PZ��!"�iDڄWpf��s"O���FN��5d��mD�2�"O��"3�V,#ӎD�����ZX�=q�"O�R��*e�������*�k�"O"�d�C"E�z%�&h�+G����"Od)���T�@(�Ɋ�A�:U15"O"|� �f���bI͢'ڔH�"OBH�c�_�A�)�9�@iӠ"O�y2-�a��@���E<=��2A"O���AڭU_ȉf�b@�"�~�<��h�7i�|���A��;K�|۳ �z�<)w�_�H�\�p-�l�<���Ey�<!�i�WE ��q-�w�<�Z��n�<Y��	?8`��f�@>lz�*'G�g�<���ą^	Xl
�LP�~�г��d�<� H)a �XB�*( �GҦ]� $br"O��PN�76�-jG�/�"���"O��9����<;4�æl͇T���p"Ot�A-�:c�ڭ�+��V��q�b"O���0�F�̱g��X��v"OA*�j=jZ���F,f�Z�@V"O@���e�"(�����/�
C�T�!�"O�a�v�Z�Z1nX�����x�@�`�"O�,;V�B$T�s�L"LB((#�"On��W-ҷG�j���@�L*�Db�"O�����S/S�r�@Q2$8�jG"O�Y򦁑�|b�����9,�� A"Ot=�W�X�}�8
�IϟA��"Or+��T�CJͰE���t.��3"O�0ƛ��<L�2h�jhv%�P"O��`Z
3��P7�ʻFعw"O ,�#.��Q��q൅	�3�|�"O���2��� ��s��ý���`"OZ$���:����F�۪H�����"Or�K���r�"�z�'r-�c"O��k�/��vv]�0&���x "O�I��F];a�ZM;c/�\��y�'"O��xEș�{&X�m�:rE�p�"O�,*.R�$�^H҅,�!o>�"O�<15��:@nhi ɓ*�.��"O����;\Iqa�\������"O6���Cn��iA+�,>��i��"OvL�	�#F�zX���!n��M @"O�y@$Y�`5���B���"O荱Sn -)�7� � �T"O0���.	,2y�#��<W�t}{�"ONx2(S�x��7,� ~��!�"O~���%}0J=)���
�
Hѥ"OZ��"Nʌ8�J�x��
��q:�"O���3�$5|j���|�"D��"OJ���(��$u�8�%�u�zp�"OȨs�"�_��I��!_���"O �@�CΚc@Z�A#Y�pG�Ժ%"Oj����F�#�PQ�d�,6�C�"O�x�b/ߵo���դ��wltz�"OJYB�(�WY� �M�1��٨"O�M���Z�a���I��"�"O8����2R�xASDP�jԀ��"Oa�@�Q%df��QABF1d�ñ"OfpQ!�	�y8^%�C�͒P
$]I"O�	։ßo�H�P�/��8��A3�"OY�"X�%+�b��6c�"P�"O���A͞.�.iqKOCu�H�"OČ��=��7�0�p"O�őӫ &���c�O\�.!y�"O�2qg�P���c���SjB9C�"O�p�qHF9��P�	j��R"O��)��'-��`
צޯ=L��y�"O�QB�ր_[��W�t-���"OL�Aǥ��Rڲ=R�nR� \�t"OT����Z�GL�����,m���"O�M ���)��D�&��c�/^e�<ag�v�B��'ڣL�-�"�Aa�<�+^3�>,S��@/~����RY�<	F�_��1���Ȧ��A�D~�<!&�ܤy2���╔2�����Q�<q0A�8_��K�֎T
�C��b�<�È�4Bw���Gv����`�<��@^�1|��L87,�����U�<� ��r3���t�&�	/�E�e"O�ۤ`�)rм�W�в~�(��"O�`�w��0)s%M1�l�Y�"Ol��G�$��<�ǢĊA"O�ģ4h�5�@0���1<��r"O4M*�b��Ix��q@EG6U����"O�s ʳ#����"�ն&��X�"O�M�OM�N*F��
D��j7"O�%�p�&6�,���j��Xa"Ov�qc�U5j��q3�X.��}hV"OT!"�L�[>̳�D-�t	�"O֜��.�3̬��`$��͚��"O� O�&�����jʈ�@T"O0�d��95�T�f�o�a×"O<5�U��L�^A����L���"O )`������+J:��5�"O��it��H������)�Z�Z"O�@xe��"T��BoK�J���B"O>Tҏ%sJXH�태Y�h��"O��IA�[>kr0X4-�8�PQ�a"O�1Y�(\	/�I�6��f%nH@"Od����׹dFt4�#ȕ&"E1"O��7=d!�aI
 �ŉ�"O��P}����d�ʹPLqk�"OP�	J��m�@�6(Xr�p�"O&��$�\�}����� *0��"O��fA��/�W��,8�"���"O�����Jf$��$"Nx�9B�"O�4�c�K�6T� �!�Sj�m�w"O�MP�`R!.��K��Q0�a�A"O �q�b.��-Ӯ;�H��"O�Q�g�DWZ8Z�Qo�XPa"O�w%גLC4y𰆕�n	}��"O�qp�j]5�d� �J	��Y)�"Ob�1�D)lc��B�og ��0"O������r��T��ɘnh`a��"OH���$��I$t"��N��u�q"ORt���%;�ZTօ r�@��"Ob��l��h,@���fP�\fl��"O�8 �����P�@v�� z� S�"O��J�(�9���Aj�#�8!p"O��*S끫<����`C�y�r�Q6�'v�'Û�nL'OA����%����e�:�y"$P0w�8񂠌�!�SЮ�=�y��֓S�>�y�(��1���ȑ�yBEE!UE��P���-��i4���yr�= ����Ϭ(���)�F��yk�XNmS1N�����x� G�y�*� �x!*�*�0�X���y�$�c�D��5��`���û�yBHǣck���PgܻA�|�&��yb��rbr���</�4�j���y�JW�U�A9��$[�*�A�掻�y�i�'+l�yK�b@�Z��r���y�R4t�0��B'^c���:Ab��~b�)ڧ#E@�2tDA9hp(��(��|�ȓ8��L�#�ψN5d���h���@(Ex��'=�9&��&T�
-�1hN�A��m�	˓�(O�<���OA����aHD9y��A"O�����y�q0Dh
�
�$- 3"O���h\�Miv�9�G�
�����?ɛ'��`�dI+"���Zĥ�8�D��'���\�$�m⃇S:6�>�0�'Y%�p��t���X��P>N����� �ͻv@&`�������	v�T�$"OfI�3�ٵV f�kR	Pk��b�"O�*�E\�U&8�Q��]V�x�'�O@d�4�� ɂ� oY�#O��"O�@aӁ xo��p�.�]L0Q�A"O�x��A�md���m�5DV��3'�'��g�B���8�c�Oݍt&(Յ�@��9���c��*�(U�]J�h��a�����_�BȤ�j$b��$V~����0�#B�,P���b�jR=���I}?�H>	/B/`�8Q0m&fՠ P�ECV�<��F\�X��3)Z����se�N�<���5&��M��B̉�&H�Mt�<!�%XI�*��f�p����o�p�<���պO+�$!��u[���b@q�'�axB��>]0h�8Qe�$%�`R���yR�&O}&��V��Q�����)�y�̪,  � p'ך���0L��y�C7t�`d�5��,~� j����y�&hH�����^9@�[1��'~ў�On�0s���KGD�� ���䀛�ĥ�b?On<�cf§�hRV&���T�x2�)�S����I�"��T�ҹQV�-'��B�IB?�ta�e�R��uq�.c�6M�D�'?Q�d���4U^�9�nQ�%RGc/�O�I8`4H�ɦ�˾"�>T��c\T��<��G�T�,�0:>�I��8Gi����^%dp E����F	ȠA��f�h�Dy��'� i��,Bme9(w
��_u��0	�'��� �c������O�V�F��	�'����5�;W{����S�"�!	�'aiGw����B�	���'�Mj�,��Mh欳r�Q��P��'��R�y�i�aa��0��'����f�0��5ҡF����Q��'�H��GI�'e���nE}¶h��'x`L����5x��; ��bT61��Ox��Cm�6��u��τ�H�<)KA"OX��ċQ2L�@�1�h���Ek�"O~�)C��9M
�"���b"O����&d��t�.K��`Q"Ov�;�%atƴH�&Ň �M��"O,��Ǌ�.���6&\.$�Z"O
@Zb�����q��α(�ejS"OZaRO��-Q��s_ uas"O��q�.B�嫖.A�x��P `"Oҵ8m��T���wM6�Z�)G"O:�R%!��]���׬��#�����"O��)�я+�>qp�E��0#"OTR�F=�nt�1�@�Z�&,B�"O���MP���#�$T�k����"O��{DL�/�6
0J�:�\M�W"O�kq�].:�D�j�7�ԍ�"O�)��X&ꦽ��	ĭ��E"�"O @���N�c�����!�@mr��%"O�I��47�^���/�)2�"O�����8 �Y�!Z�%x��P�"O��YA		
Bdv%� ��R{�Y�"O�s���e�b5ST,�[m��y�"O,A�lɯn!��E���1WL�"O�ę��E��-NfE~���"O`�YW�ߢ?"h�By/�Q*"Oh5*���k�$x�!�",�X;s"O�e���)f��x�`��_à Y�"O� u�e�IlU���Ѓ�
Ԁ�"O�� ��C�~��A�鏯x�Ұy"O��à�19p�s)�N�6A "Oޔ
AE]�:H�,!��˻G����"O��1�k
~4��Td@�S��D�T"OFY��b%8�ӆጊNcT�y�"O���� �Qf�� �$o��[�"O�TQrǒg�1@ I��zT�Q��"OZ�'�?+A�u���'���G"O�]Z�H�W v�S�O���aT"O^��eKB;)�R[$L'�)"O���RK��GN����&�+K1ܼӑ"O���ώ�&�2iP��7u��s�"ODT�`��X�pd8_i@�B�"OX��B �+#bt���)ǳ8��S�"O<���}H鐶��q �I �"Ot@
�A�
|Ԏ��� �_��`5"O�h�/A�u�"qðn��t��,�"OM��K\�#�:�+�:w���R"O���#V3p%��Ị%´���"O� ���( ��X2K�?6���c"O�U�s�(�p����k�t��"O1�p�Q�U+�@�%J_��[�"O�%u��
-~d��:X�X�"OpI���	o ����0���"O��H�B4؄���[�)r*�j�"O��� ${X0�&���
h�`�""O�� ��W�E���٢(6AM���W"Ov�%I%Y�Z���LԎ\F`��"O�-��Fv��UaE�P<���5"Oؕ�t�WQ�Ղ
�-p����"O.M�AG��~�IH��Vp���"O
i�#$�|�T=b烴&�p"O>u��TX�p�e��s�!!�"OP�����v`������+�~���"O�+#�	�#v��BB$(Iۦ�Q�"O~��j��;��p
���4D�va1T"O��r5�\�}�sgl2?��H�R"OZ�҇���EM�ӌZM�T4r�"O���HG_��3�j�/[�(#�"OD��b&W=-��@��3fAz)�$"O
j���V�բA&'�<I�"O.i�oݞNAx8��a] ��u�"OV���S�pB�}
wa�7Sʐe:'"O�h9�(��2�pa*f��!\>5��"O,�u��+K���C��.Z�C�"O�M��+�);�t�C��_� i1�"O��ie ���]@�Rd.I�"O�t0�"�J����a�-*f&)�E"O�qiDk�3�e��`��pv��	�"Op�#�!e�B�귎�/"rT�P%"ON�h��:?����c��Ov��1"OP�3���y���D"ԅ~649��"O����8o@x2@ #\xi�f"O�L�v½1���0&�Ǚumʭ b"O�)�eĮ0�̩G��B�@0!�"O`m�g�/Ao��v�ۨf��ۓ"OF�Ъ�A��m @8���8�"O�( �j߸~��ERT/ǻh���*d"O����*̕c� �� (~�^p9S"O�5��l���|k�'[��"O\��r��(Q�BQ����f�9�"O��@��� $� Z6��[\n�I�"O4�·KTs%� GnEh��'�p��k�4%*�)S)�=ڀ �-����(��%��`A#�I
5"O�lXf�[���$�CA��)v�$"O�rQ"ٝ?w2����
-�v왡"O|��ťN>�q
D�@O���"O�<�%�T#&��˲7�}��"OTm`���k�h�4(
"�q�"O��:C��/�Ȃb����S�"Ot�e(C�8�$��+G�OZ���"Oj-6,ֹk?60��-^>]� T8"OBT٤o6UH��Tf�@��1��"O%�	��S0�s$P�8��"O�<�a@;A6�0�$[gX)�e"O����JĆC���DCԵ-��Mؒ"O�UZ�hH�B��ђ�̾f|�)�'���#���+�b�!�1)�r �'gڅ�ekT�3X�
� �{�T3�'�h�j�m�'y=�a��ǃz�Tܑ�'�^��ԏ\
2��8�a�9�:��	�'�����V�u�xiЮʴ~v�,)�'�,�0c�--紌�`#��AFl��'��$�U O<{���� �J�i��'�NI�Fը��UA�kO7~a0���'|���R�4 wDzХ��w���
�'e ��n�978��J!,k�I	�'D��P�~3���b.>8(�'�JA��R�
�u��f�=�z	�'t2E�2���L�4�c�D3�r��'Iaۂ�P�>�D1�/�-�����'޼�A��I�X���LMJ��'(BĀ��2BdI��B�<��	�'�h����NqҦɌ�?�&�Q�'�m�cd�"ǐXZ�c�\d>���'�|���` >&�ݘ �^<Iu@h��'��-Jl۔v����P#ɢB	~�	�'4 <�qi^�ʤp���&B����'�.T0� �� ��I�hQ83xZ��'�Ρ�C*O+�t�&�4����'�fٚv`�.��T�T^�.<^�z�'@�Y��@ϯ|#���K#
ma�'5�\��`�7C���%�AA�]�
�'�Zi	�$��Eǰѩ���(+���
�'`�;�����5E�̅2�N�:
�'߰E:��8M��,��D�4x�e��'E����d�e	ˎ.�9�'�.�B%d��.�m�v,���<��'B�(0W�0 L���P%�X�ȓ/�Q"�.רyz �d�=r�ȓ�V�Zo�*I�n5E	�1&\LH��P
��%W���]+7�/u��ȇȓ��L�`hsՋ,Fa8��N�@� 7�̏6hh��g�P܄ȓ	%�`*S+�2�� #�ϕ)A� Շȓ&��Q��(����W�A���ȓN��S���h���9�/�#b!�D�()�����R���'�@^!�$�>+%H�B�.�n��HP�� uj!�$�[��*����ya!���h��$�"B�:��J0UR8��!&'?�-*T����?	��ԯTcB)�G	��P�� Gn8���Lߥ9f��S����GA��'ˤ�Kt���N��SD->D��8�ä;X����+��P�4��[C82�D�l��	+U@Hc�7���yǅ.5���B�s*V��C�.f]��Z�-�Is��y�f� ������
.��������<��3�4U}:[����d�W}��A��I�H���7�K������u�A��R�,��� ŢR�d�1O��0��R�f�2�p��_�(��
� v�QG�¶�faAь:t��:Ѣ��v#"t� �֖�O��ʢ�ٽ%w�L�E�ŏ1�D�i"E͝\(1����L���Xy���RP4`c�f�DI3��B\�x� 6&lq�O��@�R"̷>ߺ�jDŒ #��cM<��dH�'EN��*�*]L�����7ZL1���jGJ®.����T.P�x�I��u�.�ʒ
Q�*�^��e
4n���rg�?�r���l�>�ݝg�$"BjE�r�@���̶�I&��� �^�1�i�1+܁Б�;���B6�[f��b����-�q��|�b��+q��!a"J�E�&���ǃ.z��Z'���%� %��JA۔?�H���L_6���q��,�xU�sJ��
�O�p���´��K���9�e��WFL:rtBE�ˇ$]Q�BE�S,LVF���	����j�J_ ���%Umo� ١�xR�*��,y�C֗�N�`#)��]�8���Ɏ�q�Ӣ�&�v��$-S/��7a�2*u;�
�?K�"���I	t�!h"ѷ#�x�����N�OtM��❓E0��6\�8�)��tI�  �2:�֜+�^��X�$QL��OD�
��(�`vr=Y��H�\���!L��G��&�(訔�D����9��	�F��N�l�h<�F�y����
T� Y���1]h��O�ngԍM|B���Ƞa�]#j�܈���A=MGN��囮v ��v�9#����ŉlW��2���f�ʸ�@"@�HM�~�ЅY�!��xPU�vǗ�L&d`aQ�����i�Qޢ�ҋQJ0p��B!g��m8���_�8���%��u��B]�o�L6�#�K���Da�F�6h�����#�0���'��#s)G�e*j����S-�Ā��͟,�e����Ԓt�شO*-�#eW�	�>�x⧊o��a�tB�>Yb���)�#t����ꙶK-9�E�������
1CJ!iۄqD�Z��	bB��K�4<��bY�SpL@Pa�D$/�0���B 9 ��'}���DƭcF6\��O�!+�1�W�^OHh��'^��⚡���O(��GL̒� ��IHl`��pà��̚[���D@� ��Mh�̋3g�Ԑ����	��I��b�x������Ȣ�܂?Ͳ��`��o�4���ؐ,D��S,J�����"T�-�2� :Ʀ�'�8K"�H�R��H�A�p�ڵ��G*5��i)ѥ�#hxw-�)8�b�:�ݔZ��0�� �s�ֵ��ǫ6��UA��Ό!N�����4>�veZ�1:��
��ȟ�&XÓf��,@�/��c`\-�#@�)F��Q���d�Je𗊃�^��}�FnZ�4�h�lT�0���K�$k�uӎ�1b�@a��
�\��m�v.T�ƌ�c�0�q�BF&&��8�]B��k����H(-�d���ŉ5����@F؈����ҬW_��M[
.�������iu(�"ר���(�:c�Tm�6�#�$�v�d%C�hJ5vFiށh�
��}�ܐ#`�.!�|��I��,ݹ7�L�>�j�*�2. ��`ȟ�u�TfZ!� $4Ky�vj��0	 �@؋,��d	#d��i��}� �����B�1@M�>�%L�CT�p�bd�WĠ͑��ȃ,���VD�4*I���۟,��o�,nM�T��DL�S¨Ց��H�/���҆$�5(K�ÅjJ5^(^�� ���J�J�bA�\��PGx�kU�h�^�j�A@	@�z%L�|�J���
F�Ե���_�y��w��	lð�Q�h�zo� �<u�j��V�D�ҽ�����&~J�����9GZ��Jԏ��ğ?!��yB"W�Q�b��Oҽ x��[r� (nc5Z?�)���
H�"#��)3�II����g ���� �+3��#�XS蓟qO����ϱ}�^$��/O�t���E��|�0���İ��`:��̝]L��O���n9������\�:�B=F*��'�>G��Y�qτ�g�$�K�B ��0<Yd��y ,��$ΐ�8��W/�k{���Ԏ+L�%��I[u� ��&Ǟ?L�"�ڄ���<��)i��B�lt����O�%ц�F'h�īFc־ax\��B������Ò�[�\��!A�
�mA�A
1�'��8G'����YwnG$��dB@��:gGY���q'�%��lJ���Or�t[7X$"�����"]�+j��-O���G��
w���y�� �ؑ8fi�+{u(�P7�*:���9��I�͕�vup���MےQ��=�c��X?���$oޞ�>�O�"šM	u:�]�r�
�`�.�D�^#Vʈh��[�-�0v-?I#�O�FM���y��T1���H�#hpq�H�}%H�!��E�T��I��5O�/o�PZ#�H$0d��$��r�F�$6e�\*�72EּSr�<b�����A� �q& �=Fz�a@3��05��� y����M�um �X�$P�Ii^A�2a�:��I��޹X[��҃�.����ɩ!|Ȫ�G�1z�eQ�d��'2�'����ɛWJn,u��X���#�a/��ZT3�&�Jv��R�H-�\B��%.T}��Υ��%��mF�X
PZ�"�]\�TQ�Ҧ�X�b�A�g�D��Ow���-v����6L@!h�!��!��={eo�B�D� �[��.�QJ^�V��98Ti4|O$���-��Y����(ӑTC�D#��'�0A%Dt}��T�p1�I[CStlB2�گ�yB�-�>� 
F�;�8�y��И�'����� Ջ���3�V�E�'FNѸ��
)�2i�RDd�t8�"ONQ�ąH�W��Ɉ�EP�X�li�4"O�YP0&�
Cަ�ҵ�ʆ>�d �s"O4xr�$I�Z��̣��z�"O�8G�A�yN^�Y1�!�l�r�"O�1���N">�4�U�ǒ] Ԍ�A"O^+�� "�*��&U�#��0"O�=��$���`��+CH��}�G"O���
P�>�!2$�X6n��u"OYpʒ�iZ���	�2|*�#""O��Y����A���y��}��"O� �쐁�����`�͑Z��3"O�q�C�&�hY3� L�z��"O"��NK Yֱ"@Nƾ\�"O.]K�	ǅ�2u�%�;��(��"Oj�Ӂ"δN^)�S�X�rH{�"O�u�b�(#VF��@�/ ��pQ"O�� B�prJ�Ҳb�����{T"O�{����J��<�T`�:\7��8%"ONDI@� @��4�B�� �s"OJ�`-�tGpA����4Дhs�"O��W�S�O8�*�^�$�E"O0M����A�
\�V[`�H�"Ot��
��>�N��7�9G�\	z7"O6�t�Q#+ӸA��1��ɳ"O�	R
oq�I��,�L%��ò"O�4�T͟ /��xc�L�9\
�8�"O,AfH Zt�����&��tq"Or�Ԯ��I��f�G)P�����"O��@G3pP����2A��f"O�d2�� P��%jb���U���g"OҼz"��R��˃!ǅ�����"Oj0`�����;�O	�����3"Oe�#DZ�¸h� "����"O*( ЧI�wDiN�R����'8"�2E���!3bG�{�ب�	�'b�=�2��O
|Y�VL+sbd-��'n�ոa��1�����c݈^�`��';�#Q�A�y|��*[�K�Ԉ
�'��%x�G��j��c��5\�"%a
�'�p!�/�'x�Q�.�.�B��	�'ޚ0�c!���R���$�F�x�'@HCVh�@]�7*�$y����'i~���ܗg����*N�Jv�Q:�'P)Q�ä%�*P�(0B@}��'0���8DJ�F��3D���3�'��ib�@�7F8��*����! ���
�'��=K��Y�>i�ɡ��CL��ݨ�'�V�
$�J*۰��� ۧO�Xb�'`֥�r�D�\
T�rT�L�p��[�'��Q����5���Y㭛�)/���	�'ylE����-t�8���;5��h	�'���튍RO(�� �FfA��'�\lYA�S/8���q��B�<���'%{� _�g�P*wjҡ1�$�j�''t�k38T�ᖭ��e[�u��'���Ɓ�� ز�5f4C,��'fiX7c*!ZݪT��>��Lh�'�@� �H���1�ԁ�|<��
�' ���HɍE]��d�
�5��K
�'�^�+5A�5w\����)��ق�'�����?w��p)��%Q��	�'��b��7}Y�e#��\X�M#	�'��s�ӱ]��r%&A,!E���'��`�s����R�\9�l� �'�j���F�2�	��LO,B�N�#�'��!�2-��c�d��
KD�p�J�'����2��mZ�p��	("�(d��'z�8�Woݯ�(	����1̶-��'Jf�h�R�B�q���0D�~�'�ԁS&IK�0�vq�5c�8��Y��'l�4���Þ,�i�E�C�6���'�F��r��8�H�f�P*�'����,Ž"�@�x�m�&����']�0C���.�����Ɵ1������ (����A��bGIĞ:�����"O]��h\bZr)��Pu�,bS"O~�h'� ��v���ՖD�1Ia"Of�S��ˁG��iȓd�|��E��"O����C�Nn.L��!�!�"OX9*W�U(z�ڍ87"_�3�ar"O�ӧ��,>>p����z��	��"O�����>����	ք1���k�"O�1��6N�v�$��h��0�A"O,��5'Q��f�QV�m|~�˵"O4Qx#fďTܨp�dĥV�4�s"O�03�ǒ�B��L���x�Ŋ�"O�5dK��&6���ԧ�|S�Pj�"OF�����V�b��e�ByY�8Id"OF<!�N�#��1R���
e����"O��ð,@�C0&�T"*>X�"�"O��#��B)�-���I�J&�{"O�Y�ե^'iW�M���߁*�a@�"O�d����C��/�C�M�"O�y���E��,z'z$�@��"O��s�'ڃp�ӡ��i\@qw"O��*7aݛ|Jٛ�Ǣ��)t"OF�yp%C~�p �%v6l"�"O�G	�FH�'�>4�VPy�"O��)��[�T�y�b�:���"OB}��cD?w%|�7�
�JH7"O�bɟ�S��Q�T�#���k�"O��R�P2Hrh��2� *{L���"Oj����8`�y��/O6p)�"O&�Q%l˃�
 �ׯ� 7Yza��"O�Y$m\+'�mӐ�nG���'"Or�*���k�$l�&�/l�ƤZ"O���(T�+ؒ4�b�ƓI����"O�(���K�+![1��ibp"OH�Y�'ҐE��h�GX ,}\���"OPl@��X�=�RKE��`��T"O )����>�P���)`�.���"O����E�q�l���1@����"O2�n�s,��3u͖#1��1ْ"O.d!'fܯ�.�[1�'"�y:�"O|-�A���T`VA;�T|	%"O�PÇ��`A�$���@�S��X�"O" 
D�ć7��d��Kҫx�>�H2"O��)�.Hlh��D�Kf8%��"O���o�2���Aa�HQpl�[!"O�9��A����p0ъ}�źf"O�����Gf�A���L��阀"OjuB�
�Fb@�)�9!��<cg"ON��$̧	�R
e���L����C"O�]���L� m!T��8��L�"O"l�P%�
�	K��@��""O�h��A�5pvA�U�-G;����"O�(�d��6!��S�˛�M�q"O���[���5�T�ʍ  �4q�"O��"�D�ڜa���+�eB�"O�AZ��X���c� =Ҽa��"O������8cAļh� ��/���"O��r�qӶ�:1 ��^�_�yb��Ul�cW��h�J�O��yR�K�a �t�_;]�Z��S(���y�c@>8�a��!U�5��O��y���4"`�#�.'�(�ٳ��!�y��Ϩ3g��6���.�a����y�n�
����<���r�ƨ�y
� �(����1��e����?���Y"O�l�_�`� M2-��u�D"O��@�B�O^�	Q.�8:a� �"O�`bʽp��PQ֎�IZ>�ku"Oz�81nM-ZhV�t�wO$A��"OR���\�w7�P�_�%��p"OD��#]7~�¡�(L�,�0u"O�MY��D� �]��e�)g8f�#"OZ9h"@�
ohɫG㓑Z'
��"ON���nN	�x,p!�-n���T"O$x��+O79�@( ���m��s�"O�qp��(^4�.�04` }aA"OH�2��%;�~���OG3���"Ozy����H̢2lJfe>���"O"J2)��z�JP��S_ha��"O�����*4���(QϏvA���"O�AI���Q��ktB�`q��"OX�p��&|�4�QQ�ȵsvf8�"O��H�1<���MܴhR`�U"O���$�����R!�?-]��rW"Opl@���P\���>}ݦ�XB"O����d�_.�X)�f	�(���"O����d0�C�/�>ī�"OZ�Bk<�(�C�X K��-�F"O�B�	�0�z����@�gc.4 g"O�C��C��Q{6�AHX�0Y�"O�q�u�� �����w^(���"O8ZF�b�|�0 V�;���t"O����k84��)s�`��+?Ԙ8�"O\���`��N���:�Ж) �C"O6��4b�u(d%�G��w|bD��"O*	�`o^yU,؇�T�o��,Y"O��9��a�v�3��R}�m�s"O�B�k3k���;��g[�L!�"O�MC�ja�I	%�|���N�D�!�$G�l��*�`�:@��IT��}�!�D�&	�m	� �r��I#.I#!�D3oTl�� X<DzzSuN�I;!�D�#4D��2 ���hWr��\_�B�ȓq��ċ��o��:�b�,,0
���7
�i�PL �/�1(�g��7��ȓS�\z�8 ��i��V��ȓ[�Ȩ��MO���l�&�
$��(P"�y#!�!i{"�%nM;E�@�ȓD�d-ɂ'7�	�P�h��`�ȓ0�n��ҋځ0ظ@�BE�@��>�H��F��]���:avd���8y�PA�F�`#�9���52�Q�ȓ`��\¢'�z��cfNJ1|����ȓ
��Q����S�j�5Iɩw�Ș�ȓ&�$9S���5xR {��2G�P(����{6�D˾ Ap+��F�����&���q���w��t��#_2Q& ���vE@E� �ERexc�խ$�襇ȓ?g�q�F��wd�(��C$���ȓZJI	7���>E:���oP�0��g�y� ��(���Ye��$�ZC�|��L���Z�&u)%*�?�B�i)r0���+�Й��.�FT"O�0s�A�2���FI=4�8�`"Ot�����U���hG%��4~F���"O�9 ��W�%mдYEED�4m*�9�"O,}8��U�hh�ψ�]Y�x��"O�Hqa`JNFxT����?J-�͡�"O� <���aٲN�,D�7d t�`"O:��`N�GYp]�F+�ȀF"O\p)ի��1���۰W�%8r"O\�@P�S{��s���Αq"O ݉0����s��R�|���"O������QN��:�'�?s�-y�"O�t)r��5t��M["C�3hRhP�P"Ov0�%X ���F
L�Ȉ�"O� ;��֌y��eS��LY��� "O.�1&a�!g� �	>80�d�4"O~uB�N;�T�i�ΌO
.�c1"O�� NQ]W6�B��&7�!��"O�V^\QT������u� EH�<aa� �hkx��P��3��K�<Q�F�d���1AO
d�`�	�H�<QB)4^�4�{��L�Ö��W/�@�<9�� 1`�hS�ņv9�a�T%Y�<�U-�(`Ԯm��g�Z���yF�[�<��H���))&BF7��9#0SX�<y� �I��Mk����8����3<!�E>��9%��[J�{�oB6}-!�d�/�>ԛ' �+|>J8p��ȸ>	!���5"���2�k�z��Mx!��[!�D�����<����C�!��+C和	���.Δ��j�7�!�	��H�����N�"e��,K�!�d�6`5h��DM9�4a��Ӻ!�D՞'UXE0�+Y3
`�G!�;g!�d��|��K��}�㠚�^&!�d�~<P<r5oٸ(	��*s�\%p�!��S�W-�p*�+4P���N�M�!���=혭9��\ N�`d ��!�$
�L{ҕ�E\�c���@\�k�!���"+r�}cP�7ڴI�d��L�!�ā>=������E��L�#��%�!��GC�rac��	�������6�!���8b�@X�V��܊���� �̅ȓ%��!@#O&+�z��bY�$�Ν�ȓF@�*Gd��u���p֬�RѠ	�ȓ'Y�y�ʮ{W0���m�&H\H��r`��i��]�A!�P����������Ǯ�&LXP��b!�.a�j��ȓY����6!��t�10�Ϊq�P���\d��"��ue��)�J�n�ȓ`�%��EJ=��4!b�	�mM��ȓ�r��ޭ��dmH~�H�h�'x���cϬI��UuARr����
�'B�y��/A� �)`
�ut�eY�'�<�R.E���$(�e©P-� i�'���S�Ȋ�*,�(��N'!4��	�'��dy㄀|x�% �#�&ϞHp	�'g��!��
bl>	z�jI0C̝*	�''����!VH��Í�9�����'������<R�D�Ä)T"*�5��'��ɦ�D!�0�����/Vx��'�&��qhګa�I[�oY�?~2�h�'��SP ��,A�٥#G�O��9�'�ْ���2΄�A��\.B�� J�'	0�k�EȤ`] ]��D@B;H��'L�`�D̔3���t��?
� �'f���-Y�U*�A�$�Hܫ�'�~xP�%�FI8
&��~ �8
�'b4׉��\�p��,Wꨡ�	�'pą�1l �K�4́u��8�l�	���  ��GAC��ȥ��@>E;F"O$}{󬔧>%��2��X6zu��"O���(
5�	����#V�0+�"O|I2lȇLa�Ѩ#�Q B��"O�(�#��~x����&x��*!"OL%q5�Ϩm%N�;T.�Ǫ蚒"O�X�G�$X:J�Ŏ�-,��{�"O��硖����Q-�5ʢ��%�'_����&� b_J�be��;_�`�'�_�U9��;��ÈY}��O>1��Y|��ç0'�,�5 حz����ɴ��%�'�p���'�ɧ(�����c�'f2<�pɈ5BÒ0"��'>�мQ>X&��~BE�v9��e81f�*/��4P��`��Z@��g�S�80d�"�?�9� ծ_$b,�̢+�>���~CѕFeY�ܴZc>���xB�j�c^R ���ܦb���D�R&B��	9�EXK�/��K�.a*4�O.1���/<򖕡ɄC$���bQ��?�3O�z��H0TBؑ�h���(a�(����Y5/�~�S��l����e͛v�ǡ?D]�f��~���b?�Xن#C.C�5���X&ŦOpc����R�G��12r������V��L�����(O�>�I&�A��r�0CQ���z�&Sd�<E��'ow^=Y2Mf���	�@� ��IZy�F0��	ɬi�X� 5�=�y����NJ��E(I�&���tZ��h��>�Z7#
W��\i�nV)�X���H-�?y���B��O���I$N����o�B�F�����N��'�>�b��)^�D�3�&�<��P��!���i$0��I���u:����#P@�i��%1��C�{�f5��ş2�>�vC�6��C�ɿw��h�N7d� ���c���C�	�$#��1a��8�¶�ƖH9�C�	�\F�ݰ��`����H��.x����>�����k���h$(ʠp���l�<1g�J�����nA�7��e�C�<���"b�IcQ�f`��*�e�<QC�4)B�	���.��P��-Eb�<�����q�Ã
�"%�j��R�<I�Ȑ0�l	Ө�3���B��I�<iT挾]�ZM:����4��ł'�Yp�<�p�P*��x'#�"nP���o�<�}g�P��4��pg!U�<�@�U'������h`X$x�o\Q�<a�]?w�XeV��*��5�b�<Q���;~2�0TIU{K���O\C�<�R)U3�5��K�"�j�t��e�<�#ʳvs�|0El��t)�e�<�A+��\����?nze
� Nd�<�b�M�-o��h�ɓ�Z��đRO�b�<q �&I�)Z���4t�
X1��V�<�.XPQ�DЇc	5�\�i���\�<�!��)%��H�PiG*:��q��r�<)�_($���q.�''�f��m�<���˓+=��,�%J���8֣M�<�׭�:^Nv�Y
p�V��I�<��oD�&y QG/܇Hn��2O&l���E{dt� �<m�0��"O�i��b��<��x��޹1�D�:b"O�����	M`9�(J�u��� "O�����ř�ش�Z 	w�DI�"O��S���6"X�	��,[Ipu�"Oޠ+B c'��S�¦kc +�"O���e�Pt����ņ6`b�m�c"O�9HFI�}%(��2":rJ��3�"OV�Cd��i�$�a��^Cj�"�"OL�'"��sJ��q�֒$/� "O�����4s�-I��ޟED-��"Of�2(D�CE�I�mH�|��j�"O� Ԭ�6i��t/4P�d�Ƴ:y�\p�"O6,
����n*~���CK0+�"8�G"O�s��wq8Mؗ�r����e"O(�
�FS"�� xB�K,C�|�8�"OX�XE�1""8��օ:ը5a"OB(@��W%># l)�C�(Y�8��"O =�UJ�EB�a�b��<�"O͚E�U;!���
����M��"O��Z�@6X�`�ckL?v�8��"O�L�M(Y����tJ�/�j��W"OD��nY��}�RĚ�V��*F"O L�t*�J78|{��ͨzD��"O��G&�� ��65��@"O�9R��l04����$"O����.��_��U���n�d`U"Oh�#�ך;��"*ͥG؂�P"O����?G��<�f��%��iI�"OVq�@ %�n������1̨7"Oj��
��j�8�w�� �� "O�e�I��ܪq�S���)�"O���ɇ��b���r�(�%"OP�e�N!{ �9�	��ڍ8C"O>ŘV��	"*���h�@�p)�u"O��6��N|P�CF
3t��"O����ŅL��u��Q�$W�)�"O�����
,>�P�����#EzH�u"O,i�w����tU�F�G�iNh��"O�D�d`"a��lx�؛'Q�Yz�"O<�b	@�E�fUx H4C���f"O��Y�k��`�Q��F�r#:��"Oƨ �F�q�P�t�Pu�Hz5"O���@�,� ��Nh�4(�"O�5�al����pG$�
P����"O� �7j� ,ZCf֕`����"O,�)��j� �s�D��&˚ܢ"O���ge��*&C�=q��"OB8�2��64�P0"Y{,���"O�Q�b�`4L�X6A�&%�y�0"O�p� #Q{��$��<@"�e�"OLL��E�
��	 `�vH�@e"O���\�V�&,�Ro� n���"O���q敷o�(��O �>`���"O�C1��n����2�~\�w"O��#L&<b\�0/Y4E���"O�T¡�0;G���w�P!y�� Q"O&�Ul��y�NmcbfU.'�xՁ�"O�ؑB���-0��  -wh}�p"OZQDE	q@tk���R}{�"O8��ƛ=ɀ���g�.��q4"O��r��K�?���8�G�(J�r��6"Oz�J3	X=�Z
_s��W"O�|z�]o�L�H��-hJ(���i|ў"~nڍ�A��F�E��z�%��+�C䉜&�ҭi1�/=mNq��w���p?���Hvѓ��]�M�Z`
���pX�H�'�6KW]�r!遠H�(|���L��y�b�Gsؕ���<�@\˥e�&�HO���H��$y�-N�up}�$F:Q�B!�E"O����M-��b4`Z���ӳil�	P�S��M3B�Q#"�=X�+�<F1��ٷ+L�<Id
�tP���uh�;tѬA���^}��'�$Y�K:uD �*�eB ��h����	H7�I��)�*�b1S3��T�B�	$r�t�+�F}�D-���<V�C�)� T���Z�%b��W�[�,�t��"O���7�M�� �↷d��Bv"O�h�)�/3?�+t�@xܐ�"T"O�a3����;��ռ�&�je�_�<�w 	1݄�ʣ�ޱRm.	(2(Y^�<!�Z�C�)h�@X��(H&ĝ\�<y�ʂ	k:yJ1k�4EA��3��b�<ƣ��}|��w�-Qy����w�<�7
��6h΅Y� �&0:1��v�<�t�� M<����Ξ?e�ؑdGY�<�	�g�&X�F	?]0���L�<9�- *Ui��r擽kW29���K�<Qֆ�hG�%�*ػ-���׈�G�<�!G��I�4YXBg�6@�Mh���G�<9C���I���[05VH܋ahG�<��KH_\�`ň6 ~*E;���F�<�F��?��Pac�3-u`h�a�Lj�<� ����E�V�]������y2�| �pP�@d֐��`��yS|<$�� ><���J�NC��yBP�yݶh����)-�4▍�%�y���"B
�����ھ*W�]�e�]�yrI�zv��	q�O"�
<E���y���5G��|�$C�a���S�X��yb�ц�H1�Ð�Q`^$�G��yr�3�P���Ř\T�����yMN�qu�x��,i'TQ���ϑ�y�ʛyG�}����g�Vm#BC�y�aǶ=�N�8��?)�8�Q����y��]�:F��	�_��F��yrES(/�]:�a�����Qo��y�h�v����H�~݀�`��X��y2Ė&(=��I�L�,�|�2�(���y"�H�@���@"�A��c�y"�O�W�T����Ofe���߂�y��9��Z�㓖[�XDؠ%���y�_(4���a4�N
1@�z0O�y"�Ⱥf<����<664S0���y�C��V���C�i׃
��H0�y��P!#69!�*��|�n��w$¨�yRbc,�)H��N)I��P���
�y�,�&H`�z4�B;DO$\����yrn߅5�xd�Ţ�!>`�3���yB ��5ܐ��C�W#Nh��T�<�y�E�:~�h�p!�����M��y"晞/��ۡ .Y�rX�3���y"�V*L<��*_O2ڵ��GS��y"�ɯ
	�h% � }<�D[�@�y����8P�q���EEŁCm�=�y�ᆂ:y1ԣJD=jU���y��]�4~(�ѲLB"Coԅ��Ϝ�yn���`D���;F#lx6��!�y�
߷m�<;5*�L�2���y�*G�:��0�A 53��1����y��a#601ᩔgc�Bt�խ�y-�2�xi*���
_�
�q�#�y����8���g��@)��f�y�
[)m�t�i�,�P&xa�Z�yrHL�`���Qd�2~�&���(�yBH�4r�X�nR�{d	�'�Y��y�����bw���fxG��y"��6~XH�(��� R���y¢r8Vhbr�J=?��8.R��y�]	\v�A@P��l�Q���y
� BQ�jY5I��*�'*N0�"Oh���,�Fv4A�� �%�Da��"O��1�hR�%Xr�FNC�q�@���"Or�:w@
	@�8L�g쒍n
��"O �r%��6?���SA��:/�֬��"O�Pa�I�/��8P+N�>�S"O4�C�L܌d|����HL L�s"Ot��T�ތBްp�ā2<C�HU"O��9B��4MX.��Bj�Mb`;"O^ i�v�p��V�AFl���"O�}�!Ď�{����D�±5���"Oj}��"X}�l�s��u܉�7"Ot����^����%'�:G
���"O��斟;C����@O�k���!�"O� ��ѻDZ@�E F�T�z��"O����U/D�F�CeH��J"O
Li����$\����"O�j�Q<*��Y��@Em���"O�d��A�5~� �S('�p��"OT�×�D�Ev����J�"��"O������H݄�@2�N�P�ӱ"O��&���1KX����𴢕��yR��.U��"�6���A�Ə�y��T��BX���8^����$�y"�9% �|A[b1�r/��t�pB�	����-�	4
X@풢{�8B䉀6P:PH'𵫶&�v�
B�I;i
��h��!FH�uj
�!� B��:%�
yA ��t��	X'��a; B�InXv\�D��(��]:vG�5��C�9��e����!U�^�`EcT#N�(C�Ɍ|EHA�7�$];���(auBC��z�U��kKqH<�R�_�2C��,��2��ןK)E0�`�c��B�I(oM�� t�� Z,E�P팵J��B�	�%��x(֡��e�Ec���7g�B�I�/Z^����[�9�!��.y�B�I�7:��  ��     �  P     �+  �4  �>  �J  �Q  HX  �^  �d  #k  fq  �w  �}  -�  p�  ��  ��  7�  z�  ��   �  \�  �  K�  P�  ��  ��  �  ��  �   J �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4����T:
b�$���/_>-p嬖�`��� � Rl�B䉸i�x�K^�o[x��W!�(.�B�I=c�6��B :�R����ɫ��B�	 6Bea�K�?-b-�qL�3��B�	�%�޼h%�,`$n)25�����O���?I�ӗF��s�h�?� �!w�F+ߨ�>q��	M9^���3��[���aM�MC���1�Q�"}�D3�J�U-�)Q�^�0�iOq~��)§gr I�#����cw�Ԇ|�ن���`2N�$�P��R���o��\�=1��?�� F7Y|��x�,�6<Д��L�^�<�v�{sXt ����ʍp�U�<A�7b�j:��,S���T+[�<��
o�l�b�
�hL�j,.{ў"~�ɦ>guQ�C &m�~����/i92C��$:ht<�a&K��)Wd�>�&C��M߲q�(P>kn����#�k�����<c&ԹA��jVŋ��*�R!��V�<���;N��0����: ��Lz��Dk�<f[�O�(��rC�6s�D:��Jk�<1�'Ѳ�����+��L �M�<���%��\`HI���(q΂H�<�Ќ(ҹ@UM�kS�2Ũ}�<���W�	Ƃ�f�]���{?�'�t9��U~�/R�`�ϓF�Ls!��F�����O�7-6�T6l�
�a�C%�V�!�d؞MY����
�n���d�� �!��U/b��I�t&�w�vi�-��]�!�
/����(2ت�y�%Q2/�a{��� �a����_ډ��A+*��P4"O�pf������2�P�\�X�'�'��?n�Q����)ϙ%��\jqM7D���&�x)�dMv]�d�g�u}�xB*�g}�疗O���Y�ȍW�����	*�p?Y�O �:!����&�pV,��qTx���v�����41��gL#}Px@q�4r���Ľ>��4�~r�2;F�9XG�3!gV�bA���y2��6h�E���L�
��-��?q�'�P�`r��-;�H�K۬�m �'j�=���ŻR1����
sA�Y���%�U*	�¹W����o8n �ȓ��@��l	�y|>uiv��6��=��3D����(R*'�H�5h��*��=�ȓ)�������^��w��`܂���2��{2K͏!5:�ISD"k����ȓ#�A���[�����%�O"rr���ȓ ���K ��*���{���H�!�'��ѫX�B9�Ylh�{�K ����	�$0�S�F�R!�0,͟Nф��A-��|��Z������Y�f��_�X�P�
�.А��U��򉕓9�P���+\ 85ԃ`���$mq���S��a�zt���!��&�ú�hO?�dJ>��1%CŪ4k�)��f�)G!�D�>Z�~�1�O_j |X��0!�$��|����"�|F*H���8!����0?�����{9T$�'�$P�	n��(���(ЄW�+�8�H�B�Cv\xj�"O>06�%3�!��B��l��zW"O��	��V�]���o��pfPC��'aqOL�*��G�^�֠�TA��DTrВ�"OFP���(C=��Zo���r	�����[���S�:�����ɜ����4ě�D�rB��U�,�UA� ��Ȓ(_2*pj��6�S�O�F!YD+{g@u�ƕi����"O��r����F��� N�U�N�ѐ����	�P#��X��G!�M���P�q����n��;1��uCgJK�_'����'�[�|C�I��t]�)O�NƤ�*�"���_��h��tz�h�6D_��2K�[JJ<���J�O�dQ�O� _Fh�BpEF: �~u��'�f-a�E�=f�\��f�v����yr�OV��a�D�F��r��.�u��"O�hRw�,&�[�����ES�"O*%i�lǹwZ�HC���\��@�"OXm��F�=Wv0��ȉ*zjd�')ў"~Z�[o���9�"���!䓒�yB��r��0h�]��Ű�O����.�O��S�ӥe>�%�T�^StLs��'��$Ǟ(������mDH��F_�m6�v��4�4E�t�z��"bF�7ϪH���0��hO��=7&�����2 �.�@MS�QY�B�I� �h�E�2$X(�d�$dMr\���)��<�s��3,��irL��[;4=��J�<Qr���Xq6�P�������i�J�<�q��9q��܊w���� ��O��'� #�,Q
2SH�{�`��;h�}1B&D�ԡ�숇xDQj7��'
xi2p�%D����i�MH�r�,A<P�x`Ye.D��y``���Tlc5�^y� �Xw�8D���2LιR���1H	8�04"!D�D��,ߧf�>�àȉ	�@2�#D����0l��m#"��-��� D�h���4Zj�i��\:�&�=D�� ���DB�:��B��O�5�b���"O��$�M�[B$Yq-�c+�3"O����rT��p��!���"OP���$EASzi��DA,�43E"O��;��X%YC*T����q���V"ON	�BDZ�B�N�؆!��(U�"O`�A�M�#.Ƞ�s��4ZԌ���"O �X5%�P]��t�M�.��"OZ�9��˹"wT��N�K�Re��"Op阃	����f��-%����Н>I���)]�<[�d�cʁ�u� d N��?�!�dV�ftxh;��#�l��'��#a���R��%��g�Ն�ps&*д���*٘GavԄ�	^?9��Z1]�.��eh*�(9%�BM�<�A
�}�6l�0�դ[1��9�ǆF���M���O�raӌ�:o�"��-�+�*�Y�'�hm�ckO�YX��s		!�����$8O��KEDeKp��!��_-D�ʕ"O��I�`����P���$9O ��D�;�@�xC)Ìw6@�C��/)��}Ҧ�<'��"ݔ����� ��G��p�<���@�K�����'/x�ޤ�f��kܓ��$:��I����q��g���ՄO.*\4��S�:Q���G����A� �PH�ȓ@��b�ɳ\�`غ�bsI��ȓ^8b�G���8SH5	6A�,F���yѴE��㞶C���)K���$�ȓd���h���-���Au-�ix��'��~��M�1�mےnЁ@0����M��y��7Z�R�q��-:�b0��M���y���K�4�D �|��[�n*�y��;X֠P��aĈ�����^�y���,x����/��y �E9�y�"
�fC|�)QȜ�'-x����yB��0�~�FS�>ͪ����yr�Q'*��H0B�Q��N�i�F���y2����+�_�j@ŊƬQ��y��ܗt�T��
/
�Ɲ)��P��y͘_�z�K�H\ 
��T�b�ĝ�y��VH��R��.Z ���U �yr�X7*���.{���3/��yBiJ;V͌�ڡ% p�����7�y�*��N���v��4�Xy"AK׾�y��C&:��B"��9	��_��y�aH�YA*�uJ�p��T����yB�>�5ye�������Kޛ�y��W�L-�ԋ 65f${"	��y��!?xؽ	AA`�����yBD1*x�D� C�'$ �U
t5�y�倵t�-�M�E|R�c���y���1�`��		h��$3�yr���)��D�PM��U���yB ʠN���" �<�F�
t	���y��׽|(T�bʔ,i������y�!C�':4��Z�L�F�٢�yR��2��+w�H)Y�
�6&�yRB[�$
H-��$�g��!h���yb)UU�$�Uo�:aH�!FT��yҀ�<�D{2ʂ-X���H�mN��y�oY��8k��K)ʹ���9�y"�P4K��40u�'o\`$�"���yr�Թ}�|q2�ʠc��b U��y23>]����U�`u��G�y2��� �"`��B
�b��d��,%�y
� �@
Ҏ&�X�抒'2)�%�a"O���&ӹN������� ����"O(���7W\�p���M��aa"OPe�T��r��x"�e�Y}�""O6(�d"ޛ��"W'0hhv�{��' �'sr�'�2�'�B�'Wb�'J�	r�D�Rk!X "��(��,���'"��'&b�'���'xR�'�R�'�Z�ӦL���Na��j��'&"�'���'���'�'��'�)��_���H3�
20-�ܱ��'��'M2�'�R�'�"�'r�'�ٵ�HeYqU��#l����'IR�'<�'��'"�'X��'?B�R�K�x�Z�x��ƾE�ip��'��'�b�'��'�b�'8�'�=����ܐq��/��h�'�B�'`2�'��'���'���'���8VEܡ[�l�(Їu�Ԑ���'J��'���'���'��'��'D ��.M�ih^t!e�U�:Ј{��'R�']��'-r�'��'0�'���d�O�I&-h�#�/,$�%�')B�'&��'���'_��'��''"�k��;��Yc�	 I�t�A�'���'m��'�2�'��'���'��]���V�lە�̱8��c��'�"�'��'�r�'i��'��'�!I�*��)�F�[F�E�. ���'���'o��'�B�'��w�^���O& AW)P;�2Ń"ӻP:�[�+TPy�'��)�3?���i�4�q��D�:H0�X���x{�8	%N��$�Ц��?��<��i��$���u'���6�X�j�|��d&hӖ�d�b�"7-0?	׃�/����1��Ls5�Wg�.]�x	���ܩ��'��X��E�$���9t�x�aϗW�h�դ	2�z6�H�31O��?]������խ-��=�#�='R�J@#�>=ћ��sӨ�	A}��Tj\
i���:O�ˁM�~\T��W�3�MB0?O )�R��7u�r���/1��|B��>2<i�6��1E��`��^<D�\����"�ę��ZU�;扭2�,���8}�B Ѓ)Ǿm���?	�Y���4��V1O:�Θa�*зOmv���0e�,�'��l����(yH�]����A*EN���ʟ���׵Y�����\�� ��$�Zy2X��)��<���23[ �I+��)RdT�6L�<���i�b���O�(l�\��|6/ظ/A�*�5 �}��G��<��i��7��O�E@ �h�n�* �@qɑb� ��bQ�#O2'�
E�2��yK�	��I��7J,���]�$׀=pw���2��)bFĤ�娳�T�E3�NK2u�-�^�&���-�,B�� ��z���i7�	4X�J +���������p� ��ƣ(p��1�
�t��xa��J��j#�����0(��s��}
��y�i����&��4/Һj��	S�S�L���1�G�
��+!R%)u���v�,մJr��"�&cr~�9����$��	 Z��Š�3s��|m�ş8�	�$��%����]�yhZ�hYbT�w��S���'�b+B:�b�|�J���O���?��\W�"��Ϯt��t�G��M���ֵ�?���?����z,O��'�rl�#%;�rŪt��-℘���i���;��������C�8����݆`m�`'��s�Z�n�䟴�	����f���L�Iz��'���J��@9���W(�(dZ6c�,\T�<�QJ�S��O��'��B���`%�&JĜBF�	���"�:7-�Oܔ����<��Y?=�	Q��4X�*�+��
k�d4�q��;0@��O,�"uB0tz������̟��I��d	�m�Z1eg�V��9&F�v���'��' "�|�'�<XB��� ���/�pe��,�����+��D�O4���O&��O�X��A�Ox�Q���,�"/��k�  jjaUk�O��O$�O�$�O�9
���fJ�� ��+�&L���6I�|�!�P?����O��D�O��d�O����+�|���0WVI�%��)Zp��b,$�M��i�"�|��'�R"O�{N��xM<��,�.p��Ō=�aВcR要��럴�'�RT	7�I�O0���j<��߂r�VH��b�>pl����iw�I����ɭC~c>��	�?7�;��`Z�Fݿy>%U��b��fW��b䇐�McwY?��	�?I*�O�D��9PPAs�1v�$����?	��i��؛)O���?Of��e��h�*�`�nM4��ԓD�i��y��sӌ�$�O,�����u&���=+��%@��)&��UA0�b޴
7J�9-O����O����O~��`�Ɲ8�
9a��,I�6Ȇ��	��p��4-3y�M<ͧ�?��� w�	
Ĉy�K�=	���;����d�O���u1Ox���O>����Fu^]���G&;b�$`�l�D�Fn���p�M(���|����?�,O\]�H�9��3��N�:�!���ަM�	�a,c���I�� �	ǟ����n�
e��V$K���: �U)��E�B�n�D�I�<�I���ɥ<q�#Z��B�)�:���
_:�9�%b��<�*O���O����O�D�
��l�ƥ�CLQ3$���!� �2�4�?9��?����?)O��Dǭ3��DJY�qbDИ*�8��W�
�y�.�n����֟8�����ɅZ���n�՟t��3N�h`xV Gs7��Pa��}-��	ݴ�?����?	+O��䔵6z���O��	7<��̈��4��%��i�e�:7M�O@���O>���u� mZ�����埤�Ӯ%� 0ä�J]�:�PG|h+��ަ5��}y��'�R�i�O��U��s�� �ae�-H�x���;�"��d�i��'ٴ�	U�y�z���O4��⟚���O�X��	Ð�@���6c����Qu}��'e� ��'�R_��Ss�)�pF���&W*V���3�
Oț֧�-;��6M�O����Or�i�f��O>��ETLR�/�hN�T�Gĩ:N�n��}Zr!��Yy�mH:�������O&��G������E\�;
�!�T)uӶ�D�O���Yt�ڨn�֟���ן��Iߟ�]��,���H��J^�E��ͳ�i��Y�$��s��'�?���?g��_��Tg� <H�|����&d�v�'%�뇆v���d�O|���O���OD�d�~��	��հwt�8)A��
Nb�	(���?!���?	��?���,��@$lߴI~��S�~�����
8��&�'4B�'Y&�~Z.O��D�N�8E�	�X��0��fG(zL�%�2�D�O��$�O����O>ɡ���u���,�Łڱ�
�4��0�M���?1��?������O4�u?���(�IW�ء��ŌG��%�*P���I��t���� �I� �5��1�M���?��e�eS��:�l�����l "����'w��'D�ꟴ�Re>�O�]9&�./��!����:WĮ]���i-r�'��G1��������O��B�E�<��K
7u��C A�6��4�'Sr�'Rb?�yb�|�ןΤ"F߫{4�ɢ$��\P\��i�"�'�2e{�gj� ���OT��� �)�Ov9�.I$>%l ��Ԅ*�^�brb@}r�'�\�b��'@�T��K�i�!$�۴��UY��)����k�����{Y�6-�O\���O��)�^}RZ� ��ܥY�uq!o&5RjH�����M��ɒ�<�����2�Sџ��!T�l�p���|`����M+���?������W���'A�OK˭1�$S�a�Tc�nޫ47�O�˓U��9�S�T�'��'�
@��fB�����%u��\˴H}�����"uPmZ����۟��	��I�� �r�X$�$y0-G�>6Xy�4k�>1���<���?q��?����i�S``�s�ޗt�~�(4)�f@�l:�&�Ʀ��Iҟ���Ɵ�ۨ�l˓�?�@���\*������� ~J�����O6���OB�b�>8R�7�b����~w�u��o��j��*5W���	ޟ'���Iޟ��%�~�DABc�o���遨�u��� ��2����O��D�O��jT����t�[o}�Q[1�L_K�M�lU�W�6��OĒO����O�svH�O��' ��HV�\����£Ċ�O�d��4�?�����pV�)'>!�	�?�H*E��!�Ñ0$�����4���?��@}������S����|����tm��\|���M�)O.A�G �覉�����d�p��'���,݄4urm�4�,7���Pܴ�?��X�͓��S�'Q h*�mZ
���ʝ�BtLAoZ�v��Q�4�?y��?��'E)�'��P�>��'&[	���`�5X�6mD��"|��T�e�2�R(Y!�E d(�y1�i}2�'��!H�i�`O����O��	>h����I�FK�P٠���/J6m�<Q��/��S���'<b�'���/S��pjV��4DR*��!
~���'���'*���O��,����h�B]�$l����jH�j\�� P� 2D�ߟP�'[��'%�O��3R��v�1١�N��TH�4ň�%]�O6�D�O��O4�d�O a���j�Z�څ\U%F	&�x��<q���?����ٚ o��̧t���%���B�Cb�L	J@�'�'u�'�'�n�C�'���`#[��@�("\!�l�$h�>���?�����7cH��'>��F�	S��J!��8��+�A��l�џ�&���џhJD����H�O�ܐ䍓9OD�$u���$��i���'��	 �t��N|����-I�#���D��h"\�FI�`&�'�r�'䫤x�\&��e=X�:cW"�ÀB�E��4lZKy2�j�d6�NC���'���!&?�$i�8z�֝��԰0(������)����|�DDşx&�b?�����kԒ8uNV�E)(�sc�oӆЧ�Ҧ��	ʟ����?�KJ<��C}�灏2�Z�X`�@�����i��!ʞ'	ɧ�f�D���]�pES�-.d���O�%Y%mZ�l�	ퟸj ��ē�?y���~2�\�*Rܐ���r���؄�A��McK>�����3?�Or��'1��q�n�"��E�F�3�$")�F�'ZҰ1 g8�d�Ov�D,��� ��D)ٖc+H�A$j�;>�dj!�i��`��RW�HrG�ĝ����v�xB	]`�L���O�q't�X����!򤑢Y�Fx�a�� ��U�� �^ Q�������1@�O_68� a%��'S�Ȑ��a�3�~5���ܟ/S��Â�!+�!kR����K9&���zqd�%+�Ε��х;V$�SDu�qgٛD"d-�We��u�S
C�0bD!O�����KP�XU�Ƅ�,9Q��+G�וe��֩^�7-��HFH.)��3UO�,x��eS��ŞU��D�Od�DX��P(���79� RƉ5x�˧7�б#"�	jĝ[a#ߙgV�Eyr����P�@$��;9*%@�DL'�h%���W�8�����g��(Ox�9C�'����ݔ�@�G�>L���ʭy�D!�O�`�̀�pd�!�nM�_��"��LE{�O��O9�bMx~Tz �@�n���63O�I҃#���ן��O����'I��'�� {P�f�L��b� ��k *0g�(�c ��6��SE�'���Y�s�� ���$C�Z�N��c�Z�^`�A2G��9rț��X��L�!�D��	Ђ�;jټc>��Z�A>D�s��<�ݙED��-��OP�o�7�M��舟�H=��%��iIpp�Ǘ��y��'pR�)�S�R�zv�n�:�y��C<u�#<qпi�<6-6�䝺��d'�I��m�&����t�
^���'2$����� Iw��'�"�'��םٟ����B�p��P	��A���&ԩB ���%�(a�'��N�	#�d�?�=��~_t��E�x��2.�zwLt��'�=�(Q'딯!�:����:\qb$��i՚�3A �	Vn�p-\�� ��r��q`h�� D{2P����ܝN���e� �@U��@��&D��ң��h,b�Ë�,�L����HO���O&�� �K��ih�x��I	P����Ɍ� ��i�p�'���'��� ��'��Iņ9{�`i"�˒!�he�$j�&l(���E�y�����'b�'KA�l���k�DH�j�p5��4�%�ï\��0>G,��������k�%@�#��P{��Q"=��'�t���L�?�O���q��Տi���(ߺ<{�	Y�'M�0��6�4�(�0B(��'�����DR�9h�oş���^�ħ@/z�:��܇4s�L��� �.`�x���'2�'Y���� �?U��4p��\�r�T>y;g��p�� y��?{�Vڡ�(O���&�|������!������)�m��䀾u��4��`��(O4 �'�R����'����@�\2s�uS��4X)��'�O?�	��v,����]n��"C�8`<��d�^≀��a�t		xx^,QOE�$�I�sԬ��4�?����)C�"���O����LF-Z�Ț0Hq�6��uo�R�٪=�l��!]_��l��|����yX�BEM�i0d��#�H��E��S�$��F��e`8�
�"r��E���4NN��)[Xr���X�1�~�HӤԛ�?���i����?uE��h3Qb�N�t��9c_�b�@ϓ�?���� ����@�l�!�
"g����<���k��P��ʟ��4��d(�"���nH�{�
�˟��I��4�� �����	���I<�u��'e	�!V��g�وy,�X����~��$��>�'`�h�|��da�:<#X�K#�]s?Q%�~x���D���e�z��ibp'���0���O݇�	)���N�#h�0��,}�jC�ɖ 1F��T�h+��`���6�������4ڴ*��ے����ހr�Ux��i����?y��?a�ѕ�?�����KX	�?��Z��5(�g��lb��U�X9y��D��U�,��l��ԡ��6,B)����5�P���.B�z�dH��A9O�8R(y�2T�ɒe`�L:D��{3�2A��e���n���U��hC䉩��!��6:9��H�gw�牤��'������{Ӣ���O2�'C��(�g��*�)d 9WV5ҡN�?����?�!]8/������:���Y&�k8�5r2�O&�^� �I����㜬GPr�Eyr�����aq�Dy������0w3��)1)�,�2�a�*��maQMY� 78��9o�'0��yn�>�`�i���e��
����%:D���cV�o�J�� ��'5��%�G�:?���4��T&��A�ɳ/Q���3o�/2ؙ�u9�IQ���`��	`IX������X:D�t��$T!mb����S��7D��S��Щ@� 2t�\�|�B}{U�7D��+���,I�J�(�H� /@
QB��8D�h�d-��Z:Y��e�N̼ ǋ8D�$�� �*��5���X�Z�"�c5D�P��@�i?<IIU��IvPpS'�4D�H�GȌ7S���reЍ �r�0D���b'@{EV��`��ZW�h*O��h�j��q-ʧ fv��"Om�'�ɰ#�~�
���#����"O� g�בV?H��Ƃ�Ъ��a"O�	��  W��`�Z�)���"O�Eȥ`C�����p��.L@��0"O|칓�2/NTEl^�YIB�ۅ"O|$ hN�}5B�S���)��zg"O,��&_�o��H����{k��P�"Or��B�� X�0�*V��y "O���U�IcV���C�N 0�""O� bI��=z���!yK�Y#�"O"��&;n����@��f�["O{�J�Ȩ &� = �zS"O9b �U$���D�k�hr�"O��Y�"ǂ/SB]�ƃ���
%"O��ZFNƷ=�p1��̅�6��m��"O���F�g�:ej���MiJ�2g"O*ɐ��R�uPY��IP	;|��b�"OP���F��FiTȈf(��H���"O���)�༁bq��q�|D;�"O�2'\
c��I�E�e����"O��Z�䌳U|�d���n�;�"O x�v�T9NmL11���:i�H�Zv����)�O�[#U?y�r̔'>�����)Кx3d
�m(�KK��p?��(�lZɉ䊘3
� �!�
�PĦ������ ] hΧA�^wD�Pr�t�	�*�
]��+';�^�p�lMjj.B�'9H�dP�����y�^5<��y���Xf�SR���E9�x�	N|*��Ɏ?��(W���o��|.,�s��+�O���߷]�~Q����:E�}��b�:���ȍ��uP�X��R�Rc��#2�ssM'�0.��b\j�P��D1�ߴx=1Ob���妡��J%C�0�5AL}2��6}ph�G��.z�(���0��l��6�O���!�ޕ,�z��Oٷ(���R�#��<���{�|�&�%��3?�O�� ���C0�@�Ȱ!݀ p�y$�"LO@eڔfP�B8�=�'kR=��
��o�l�r����C�.Ń. c��A��l|�aKǵK�4q2�X���V�[�2DlK@
^�|vX�x`�1�I�<�X�zd������=0�iI\���@�y6��%�P���і�Z6x���*ߦ=8��6�zڕ��OX õ�	�+���s�M�a���ӝ'۞�J�X}ҿi�X!����	<���	��	v�.���˲`<�������p?�-�����!M8V�4��RoW�œ;O"�D�&��T>�iuv� ���#��WTdh�C�H��U���'�25�W��M��Lʈ~��|#홚�$-�pbۆ_��AAQ\�� aɦ����pR���O[6����y,��U�~yQ�
_9`A��=��'�C���MӶ��o�X�I'�|��i�>��D�n}xB�盃mo`���~���O�d��8��� �L��#�1H� ��� LZ�xhĉY�t�� >
�ŬE� F��e�P�|��|*���G" �0acaU�6�$T��<1@  ��'�$-�E�d.��S�j�c,��޴E٢�Óĕ1��S��OX]�%�ĺC1�-+7����O�q�N!0pG�E����#b��'��4T�`7����r�k��	�`��"c�1��dO�f�Ni2S���h����	5Y���͓\�|xѷ� x �Ŗ7�`]���նwD`\�"���s��@��N?��KɺB2謚��ʈ
g��`V��џ�) �ފ)����tΟ/&�n��C9����w��/
7�)Bm����e��;g���aTVy'����B̓Ps���3��-	�)�O�C�H 1�؊}�a�M�S�F,���r%�M�v*�0�'��L���Ѻ;��/X�:� g�Q�`z�(Ӗ��<��أ�eGk��$�G/�wv(i����)rq�	��o����b.��XcD����d�(P�v��d__:X��L6m1���!�5hD&@�����7$�D��<����d~D�pD�
"Fe�D]̓*�ŉr��4Iέ����c٦qx��O�h��!K���:x�;�e
g�B%�
=:�ʅ�r�.H�qI��� R�ѡw�Lkw�퀅l-LO:
�8k�U�ҏ�����S1 ������xJW�ߴ�$e�� ^��a}���
�&���J�/4����gA��&TF�w�T$G%���DF3j��G"��R}|�+p-�@k6\[�6*��=2U�[�E`1O�<�p��X��ʺ`�P�Xw&
q���O�,��, �m�`ĨD`D9b�q���
�}�l�$�mA+VB��'�j���J��)�(����,��A�'+I�ֆ�p)��(�?$xj������:�m��'�$O!�@ n�����F�=�BH�JLj��	h�m��I�z6	[��A�1�����щ`2D$��o��5j��dL�h�d1�f��?���c�� � ���)v��DS}R"s��O�@�t�B�s�@�L9f F�Q�`w�H�ӓ\��ӠD�{r$D��nXh�aPnޚ$GV��c+C*1s�ႍ>�yr�'62�7O���
T��O�T	0BA1�m����hZ�P�}�����Q1,�(EE`�m�-]'�^��]?|،}!����N��� �@W[�@����(�DG�����O"�c%+H�&�9؋N<�2!�2�eh&(O�S0�����,��S�4�鿓�˘�Ǝ��-�YyJ����)u:���e��1�0?�w��1��e�<z�	��Ԧ�M<��.����n�8��g~
� 0�!�ꌫO��8��Ӓc�N-0v�'D��aّ4'��i�Bi���R�)x�H���U�X���]�,��'�G�~��ǮDj��SA���y�%I�j����Kq&�t�0)[���'�:I��%J/~.H�SU�2�1����$�AU����B�/Vr�аhG"�R�:�b-,Mv% E!�0��Oj�rV�U�H$�J�kCN�BL�g�V	'�^t�@�Z�496U��$�4=j�<�Oޢ� �a١n!"UfD�.��m(�%( ����	|��$��C�3K<,�A�#�6�}���ĕ>at�F tx�NΙo���Fܪ���h���"waz"f�#�P5�AI�{���ywH�%�L�ic�
IF@(g[���D_���&��s���ɺ����d� ���%T��?���R*W��u�t��X8p�8@N�A̓�p�:DFá{Y.�p�L'���mz��;��y���N:5\Xh���+.���'�Ҩ��JL�Xp+�'��N<�I����6`V\I@3D?u��8�aPS^mbͅ�<�S��c��k�>A7L_~Z�5�4"�푥Ci�bV�(4�%��2@��ҥ�1����͸�2/�Xc�P)�O��+h���Ԅ���W�ZIy�'F�����<�Z���$� ]k��C*F�P��^����IU�R0@���U?�2͉
2�h���#i�C!�ѩa���VT�b�����O}H�tO*YN��Lu�x���N��W��)��_�[��T��O�)�U ���<y� ߹b���g?�ƆP%5̆�a'��_��` ��!��d<6��!��F�/F��F�@uL��re��9;�b���A��l#�	�n���R=RS�i���3���R��O�':�����#����Wx�nu�w��*l�Z1��"ݲ�蠦MM�x9)%`̢.=��'�z7�����Iq���Q�K�X�����Ő�yEh��T�ʬ,�Nȸ	ӓb4j}�cmF6�d�r�dϷ+�2�ȓf��"f�S�O����ю*��#�$Ө|�8�D���pXg��k��P�4�Ѳ�!��G�L�	=�'WL	�$9 �XDK
k�B�x�4��5oZA��$3.q3vC�D�r�25��X�u���[>!x�ㄉYhΡy�"ړ.��<��*J�0v�y3��7(8��鄀�#;*�5gϊC,q����nH�f�I�'ެ8 ��,��Հ��=B�y�Ś#0�)��	�T�X�`(��:N(ce�T�����8Ƣh��b���Qd$��p��iC#ċ[[�Ds��rm�H���DN^�����(�; ^V�iWOҿJ���{ѡ>����C�(]�����x�'���Zb���\BF��s�T�<�Ƽ��4+�0E!�4%�����!��D��1�'H�	�Bj�?n�\%�⁙�3���l�2�����]^����(��{�f� $fph�W��N��y�a�b2s���)X4:`⧠tݍEzB��.�R`sv`*w���@�N�)d�A�f&'�ƀ0���D�`T�@�ty�܎��Z���'κUM�h#G�F�F������ : ��Y��'IP���7[M �2�
ěI1�4K�ؘ]��|�� 
=C���"�v��?�>�iM̋#>Lir0ʊ�}/2���X17�axbB��1��Ȼ,��*R��q���z�FI��~0
Ҩ�_ϴ�Zw�W�I?�e:5�� Xß<цcͭ;�^�o�� �Nᎈ9w:ڱ��)�}N��'n��`u�K 
;�eQ�ɉa��3�FWv7<��W� �,H�&sl��� *Hz�� J�>�g�ߤ$�xQo��O 4"�$X��HO2��j�
���F�6��i�,�x �`�T�H@�T9o�*M=e�'��O��c!��n��(el�YpU�J�~���#��
a|Zc�,�0�p��u�?=�2d��!Ē,��^�Ba�O~u
]�nl��GT����!��+�,:e�'����%N׮4Zp�ĭ����$!�%r1D �u�q8��U�5��?Icp�72O$e�@&�( 9N��O^��ش�`ṧ%[�d�<{���%G�>�&��{�Ƀ~|��|w�e��r�<��|����!>�MhPq�$�����7��I��a�%FP�D{bPs��[�ў`ae�$o��BU�WU��6v�@�b	ۑ�TTzI<�ϸ'^zd�s�
�':
�#tA18dp<��Wz���{�:���%���<�ƞ�;�8��O�{��]����G#GV<�96c�3�<�ir݈�f��+�s��yrͨDBf�lZg�,z⫂�	<�Irg�MmiNu��I�B���L�����F�^w��Hpc�]=-��ӧ�yrnB��P�x%�ԊO���_�ēU��5�ߟL���
R/d�'���S��9�LC!4��?pg��陾#L4��IS
,(|�s���Q��eg�Y��I��&�
�r�M��� ��4K���L���k�<��'{ҥ����	wq�}1�i�tr�+M�[���r��[���/�.����dJ���My�D¡:~��Iz��O��牷4=n-S���'�4�5�
1j�ڐC��\E�<��d5"Tt�#�G�t
��ɠE�~��,�u���۵��41�&$��c7k@�<� ȯ|�d"�63��"n��<1�h���x��! C!a�L�ӣ"_�	�B�� �OU<~F����'��	���s`�>j�%,4"�n��B,3*8�	1B"A!f�F��D�0稒W�j�>��Ax>Q2�E�X���)���-������TM�P�lA�
Ϡ�OB�[�ʸ�n|�B�ʴ_"$4"�E��%̠�y��벀#a�����0u+|t�`��`}�<��d��n����m7P8yE+E��4dЁ�J�S��X)˓�Rhʤ��*'R��VO#� �]¦�	�V�C7A��*^�X��	ꦥ��E�7Q���ȃf����'�,5CS!Z��T�Q�A<�K>�P�A�����Bt�Ᵽ1�NܓSr8�E�A<5�����H:4������)�>���A�����8@��Ӵ,f��+�g�-@���E��#�:L�fnO�2��78��?])q���<i�,���@�v*Ig������fK"a+u�'�L����"%�@A��X2�xi�}R��|�Z�0Q3}R�xB�P���2�
LsN�E҇�0=�W�y���&��#���⦈3N������MC~���떽o�9�p���<���{<�'�4���aد���ߋh�N��)&��E�9'�'��$8%�B72���ye�	PU"�È}B넷u�x@p/�>"��2��ˇe4NyYK���4n��x��5-LD#砝�v����遻F� �S��T2��6��:{<<�<����d��Mü�Q�O3Skr�Kc��b�`q��sh<iR��(��,�$i��J�ʙ���
eΡ��1OvnZ�M; <O�݂�Vh>�^@PQ�N�
B���e��~؇��T�pcH
yĈ�edr�4�ȓF�d�'c�,[�������I���ȓq��e��`L;f:Τ�ѽaW���l�J"LE�A�Z�o_�Vz���Wlr�80\-B��H:q1� ��E�^I�;�y�)�/T�X��8�1���SB�,|�1I?>E, �ȓ x�J�;V[��󕁝��|��ȓqmn�c�+��fr��J�$�)9��ȓs����F�>�@uB��E�=����0y �'�!"�,m2��ȯCQ�P��rD�02�̍�z6�Qڇ��N����f�6�+V�ـ��`���iB���4B|���l�(�Wa5��هȓs3�脁�$n��h�e�/2 :Їȓ?}d(�ѫ�	���N!�؇����5�Q�=J��bsaMKR����+����l��Gh�Z@��g�u��Gޮ���@ ;�$j�N�&E�ȓn��h�w-^�),$B��,x��C� A�gN�r���h�I<3�j��ȓ=��0�ΘBvN!c�:6�`@�ȓ~�ѐ7e�������F?`s4���R��Ac�%>��kRj�4{��ȓU�(M��)G:D���ꊳRψ��ȓ/�`�I��P��:9J�f�.I	����.h��X��E'c�RI�W �c\fɅȓ5HF��G��mK���7.�D,R��V��̑g��x��� Q�Sx�v�ȓ�f]��)2��H"�Ε0�ȓKF�Qa�+ȹRL��)�(D�$@sB����Ǉ{[��:W�&D��yN�P�9*VkK�5|���O%D��"��U���K�d�@Pf�1��"D��p���_+��҆,6=��#!�<D�\[��F�|�����n�aP�a�(D��Ò���a��l��`�>
$D]*�I(D��qmT��q��7'\��rG;D��;e��,UJ�p�%,e�]@�>D��R�"�(g��Ǚ�*Y`9jc�'D����
A�hI|��!Eac���:D� ɅKޡ�n	�ū��^���BB�7D�x(Wn��2��rG��PA�LJ4D�t��aS�j�&�s�L���t)e�0D��ᗯ����z�r�X��<D���Ҋ	�8qd̊��ҟ(P,j�J:D���7�́o�X(j�jģAS2�C�
:D��bV��bk iq��x�B0�2	$D�xK�
#g>����M�.���$D�Xyv�G�/\(aŌ1��!�a�.D�� � 2�!�)\>��jdD�5����"O��dCX�A��9H��S�1�M��"O�D��
1*<����6t-ʴa!"O��@�/�#�f�ʡ���t?V�`"OL�J�.'�l��Ǝ�U'�:'"O���g��G�����\�n����"O`h�V��9��e�&N[�
{�� "O�!1 �+&Z��G	���BL�G�<�Kݱ@��H[���BM cL�I�<�fN�9���ePC�v\��F�<�DK�.���@F��|�� *��H�<!��V�:�,�AW�/�@��V!�B�<�T�טX��Y��#}x���x�<�GY5�����:�RY;&�}�<!���)}�r�r�,ǖ���s��<!����ңl��:X�3$�<���(H{~��!�ĥ_k�}�'��}�<��6r씙P��ݟ?�q�-B�<aр�zS
���hkRia2��A�<a/��_[�������t0)��u�<AՎ���Pٲ��<��5�s�<a����&��^MB�h�Y�<єFʊDݾEе�/��M�CCW|�'��x�B��K�$yy�aծ#�Ҕ���yR����>����5Wđr� �y��ْ?L��Ac�1����To���yr����Je�=�h�H !�y�����Q��o )|
<u�d�Ե�O��=�O�4� �_3N�cf� -R�K�'u���,P&�`u!v"�4�]��'t�]��ɥZ��y�"�"vd���'3�ɳ)C�T���K�FK&oy���'�U�c��m����	�+i���R�':��!�<(�� 
Z=S��IH�'�+e�N#WUn�h�h�3UE��z
�'-t�%�4��K��_RDj(�
�'=L���sd�iB2�EҺ1�
�'�̱�C��=q[�ŋa� 
Ul���'j�!�#嚬@����wk�4�Q	�'֨��DB�g����S�S�2��v"On����R�D����ѳj=:�B"O�!*�EG8o�}����p-��"On-ROQ(U���K���p�r\8�"O�T���1)�2$��۲ k���L*�S��y2��+Pb��@�NE������.�y�j�J.%�DHɼA������Ա�y�j��T����#�|�r@lY��y"(N�_VԐ��M:c{"0�P�yRH�h��e����'���3p�8�y⌋�+���U+��%�0�h�W��y��I2X��X���-���&���yB ړ]C潊Rbʠ��W�N�y�%�*t�^��dj����d�C��y�x4�q$���lX���_�yB���x�F���S�j��b�ؒ�y"�@�y4,�r�� _ p���y��:�\	�e�3�xy	��A#�y��,v��̲���z����F �y��ޮ[��}���Z
p |L1�hҨ�y⌓�KPx$�DkL�k��c�㎤�y"��АP�
5:x�����y�"S�HҰq���M�����yR%��{#n���y$q�j�yU�m8�AҨZ�_"l��A� �y
� >���B#D���)�$(&BŨ�"O\m넃�*N��p���?M�,ūF��k��U'�7IJ���!�PG�֕�d!D�Ls���H.&a
��N�<s�1��,D�8XpC�F}̄��GK�@��]�u)D���ǀT1tu,�I�(Nf��)�'$D�|5��)��u��B+H��c�=D�X�FBJ�QSFYh�I�r����`6D�h���"Y����R"����4D���q�W~��!+�	��(�e1D��:��� 7Z@U2��Ѧ$.<c�,D�4�0�A�&��ѠeQ�QWl�X�c,D��x�e��x��:�O��j�k�m*D�����wF�(@�ʋ�Q<(���%D�`���	~$��"i+�>�$G%D��ri��bڦpb&)�?��]�%D���̀7�T�1��?G����FCFh<A&'�7h+h �#>`���B�I�<Y l�1/Z�6�	�G<���kZA�<!f�"x�����HE�bNS�-�u�<�Sφ�g=��iV�XSV����y�<�#���T;���%.ҏA��L����~�<!��,7����TK;e�-b5��x�<�GGN�US��ǋW�H�z�9�n�<i"䌀�(aueR�X� 3&��s�<�7)�#N�\�瀽zn��@dCW�<����(,@x�f]�R�qZ��O�<iCGEp�d�XP��	��t�<�3�0���s"�Z�*^�)�#Jm�<����7�R-a�d�E�`Ly���q�<I��DZ���*Katݠd�Bn�<уND�M	tT����}��,���i�<��#���EO��J�P��p�<	��#QX�Ź$Ϟh�|i ���p�<��!�,"J�UE�G��1�"�Zl�<a�qR9 ��6��b��\�<�w��74��]���D��ӠU�<��aTD��уT�мSR�Y�<)a�;$Z�B5KЛ:J�h�R�M�<��I��+���	ì�{����A7D�|*��,��ڀ�O6\���3�6D���rcҙ@��]�qDM	�zą0�L��
�JVU�>s���GʀFƐC�	�)�R�KQ�Z3+�p��<3\C��1q���ǩ�.�0�U�Z""~@C�� M.����C,x�̉�� +C.C�I�	�\�ڶ��i��ˀAB6[<B�	�����=K��pr�#E[�B�	]b�P�jȉP�5���[5�C�>�M��ڌ#��\:Q�Y�w�C�>	;RXc��<k�k��Y-c*�B�	<P�@ FM�l��I�E�bߘB䉢+.u����ԙ(%눹_�TC�	�
�h�s�)��N��~J�C��;5��p@��U�3�A�'�B� �B�I$�݋�*�K%�1҃��;:��C��0O٪Hysg����6��a�R�ȓ.���L�<��1��%�ֈ�ȓ�*pq�F$c&��(��y��,�ȓv��!!�qi� �9ǴL�ȓqà��G?s.�J��-�R��ufq㈚ ,E\Œc��8t��(��c�TP�ଔj��U�2*�56�ư�ȓ(P�(�� _��}��	�+8)��S�? ���o&ĞX���/�p�'!����JK�G6ܚL_"J�XD��o>D����d̈��Y��'T#:dYI!�$!�S��(�3�	��X���$_�,��D��R.�)�E��r�A��T.	>���"�zq�Q@>_���ß)�͆��|?���Ў^��� �UL����/Yj�<���R#j6~�f�CB�R����e�<���E�`;l��K�|h@Z2@I�<YH�$`��	_[@=�.�_�<���8�h��ɀ)<x$��[�<A�Bo�~p+��[�h�&9���Vk�<y��D0�b-��H�-9���P�C�<����bZ��e.�:�h���-�~�<y�#�S�٠��ިDP����<i2�L0�Qy��w��p�B�|�<y���Q*�%��J�X�)� Ya�<ɶ�<O��C�&E�p�F���K�`�<yQ$]j�0��1%� C�MVZ�<I�'�K~-;"���TZ8��ga�<��3L<��KV)G:�l�	�]V�<�q���|}ɵI�.���Ү�Q�<��D��
t�#�#�>�aB�K�<�����  �� B�s{�8���E�<���\��
+15�	�C�^D�<����;m���b�f��Y��!����<��)������"e�tq�B�v�<�ũN>�|��DIp���*Zo�<�@&�Td3�U*�ͲՈ�d�<a'� �,��U�X��iB��l�<���F�d12Ŗ�;��q�_c�<qW�*)cf(ٲ+
�
���0r��B�ɷ��c�k1&����� #�B�I�^�p*��Ƥ#�A"�l��C�I�o~��@!��T<x"��==iTC䉬:����KQkt���JK"l�B��%3�ъ�Ʉ�b�b :i�:��B�	'F�\Ԓ��+�:�(a䆸؎B�	�@����X o�Z4�ޮ87�C�	�V���u	�?jLP�`��2zTB�v	��B�a߉ �MR�-�B�	�W��A�^2�x�B��8)�C�	�4s�Ԛd�U�$��!ˁt�B�	 PԺ��Z	�4��,�UD�B�	 Ji�����-O��P�S�7�fB�ɬά�hRcXA8����E�i�BB��!|�x���2"	���A�T�K�8B�	�@�"aa���9a5F2䩟8��B�	#[��!8� ��'�5�5n_�fo�C�ɿF7T��F �Н���УP=�C��j]���J�9-~� $%�>B�	�T۪�k�*�e\I��mAB�Ɉi��I�[
��H�cњ#;�C�	�y��k �>=S�n��q�C�'�Nhx� B�2��{Pl+_l�C�	�W����c�D�z��r&�I�w�C�I5`�{��Ǖk�Zē&慵QtjC�Ic	P�DFw,��1�֜MoB�ɐ7��dYfB_w.f�*G�0�B�	� �r���l~rp�rJ�@Q�B�I�w9��r#��H� 2d7}hB�ɚS�a�p� 0Q��e�'�:M�C�3����)�SP��ٰaS�^�B�I|s4�Q��Һ7��t{��5`Q�C�)� p� �.B&�n�9���(K"OhIp���h&Q�&�E�A����W"O��a�O�^�yґ� J�j���"O�}Y�#I3$�t�a(U�5)�ɺE"O����J�<� =
�F��7���W"O��
æM+5���l$=��l#D"O��!jL@i�(�U�&w8���"O$t�E�2}y�i�PJϷv_ !3�"O����f
�E�YJ�(^6V��Ո5"O��b7��
)�z	��H�,�*�"O������Ǆ�s�Ör|XxR"O�AHC�V��}�&bK(Dq~��"O�Q@�O�2�|���@3Uub�"O�h;6c�@-RC!O\K:k�"O�PZ���h|��Ј5d�)g"OF�Yf�\'2#>9cC�O�U,e8�"O�1K�c��z�^�(�g�LX��Xq"O�	��
2�����JG�pQ"O� y�k�J0H@�E�69v�6"OT)��t��9S���'%(2ٲ$"OȤ14�(�<��m\#o:��(�"O�¥�lFbT����b����"O��a\fd"ݙu�T��] $"O������>.Y�&�T)f�q�"O���t�j$BE�o#b�"O�� �{r�C �E�S��#2"O��	#"�^����ψ�?��6"OD�����|����D��<��"0"O�����r�॑��?-�\��"O%��E�P<�`���=)��щ�"O�4��J��y�띠?����"O&���^�R\��
��"� L��"O�h��"�	N���g�
=ֈV"O(At�� |(�P��Թz_�a��"O|�8
Q�&��� ��Z8Q�h��"O4x�q�#I��ثUDG9g��-�"O���E��'"�p3ҳ��;G�G��yH̠9'l�Q��V�0�&$/�y⩚2[��'Ƙa�z}z�iS�yr`F#k�8&� n��|X����yr�x������'1N�c���y�do���+,7�� Sc��y�l�<y4��ʳ�����"-��y�]�>^p�pȁ�|�:Y���y�"�/�t��w$�o��	pT�ˡ�y�l�nT %����*3����O��ybD�>*Ř�fS�x0L����y(U�Hı�k� �I*����y­B5�yIG�Q"�Ҥ���yBf����j2;5���,�,�y��߈Y�����^�0B6�ڦS��y�[7��m9`'_8X�ͱ��	��y�	�/>�8!��M!!�¥ ��X��y�҆�P�2���H�@c��yb��G�)9'�Ǒ&����jL��yr���G��-2"�C$x���W�6�y���4�
�s3$\��x���KV�yb��=j��v��(2,8�&X�y���3NMf���ү5��jԈG��y�!R�T��csd�$����#Cˀ�yb$�.�4R�L�qiꂏ ��yb��|�f�S`�r�@�r"K4�y�J�$š�cη���q�?�y"�H0"V8�X@C)�T�*�N
0�y
� �lòm�Y
�AZCfR�V#"���"O��Ɲ>Q2�Eb��˖M��h�"O���ׄ�8�P-��ϟr#���"O��$�.QXµ�Ui�>_�N��#"O:�9fa�]Ҏh�f�L�����"OȤ%ct�����M�i�h�y�"Oڄ�b���"]�aA݊`��P�"Ot9I�۠^n�)�� �B���b�"O����F�x�g�3�&ġ�"O(�V�!|�-P��<��&"O�[�'�=��lеL*�Ԑ�"O�a�V�_��B ��E��NDq�"O��0�I�.SdT�p��^:�\�"O
4SD��#�¤h@�*>}L�"ODӁ��-l�x�����ԉ�"O\͑bo�/C>L�1��_^��u"OاM��P *�B915re�R"O:)��i�Pi BGɐ�y�d"Oƙ�p�K�
��p	fc\ 6QPq"O�@��D��Qo<�g��4u��a�e"O~`S������Q0�!� 7��)�5"O�EZ�n�_�l�� �B�=�֔�"O����	2�\qs� �:��ҡ"O2�� �J�|)f�֝�����"Or�ᣣE��Ph�mN^xH{�"O��D��
S�eJWC@q��e"Odո �8#��jFb��F\H
'"OZ����G^(���!�:P�K�"O�*jѴ#F�����3���SP"O쉸�ݭ�jD��G۳hl���"O�#ƬR2���k�'֦M�$R�"OԂ�X�;�1g�S7���`�"OH��@�K{�x���@�n��e�"OM�`��O�&��w�X�eI�1"O�11 �ƅV�����W#P[��h""O ��ڜu���8qA�N9��V"O"��l@6���tME�D�4@)"OȀ�4ǀ�ax��+e턥d�BԊ0"O�7D�"~L�AB�3nt�q�c"O,9�B�1|x����7e�j��"O����ͬ_e�W
ĥ]w�(�"OF��� �H:Hd��K�S�� ��"Oj�2�E�0D����*��#�`y"O^�*�B�`m�4�֮�"�Py��"O|��qf	3CÞ�BY��֥�@"OfUʳ,�Dv��!�ޥ#�h��"O(�h�h�5C��GQ�!�	��"O��!#�]��������*^��L�G"O�9 �~��AHӴf=���""O��G�EGu����m͢#�r�ٴ"O�ѡrE6X��i� ��oN��"O��`���fB@#/i��"O��8��)nH-A�ی,b��p�"O���"^�:����"d�$^���$"OXm�  V<N-��ґ�K6h��<{#"O i�pJ�+BP ��u�ڨhR"O�)�N�����d�¼��"O�PY�G��Cc�9���ʲ4�Б�W"O8���&ό��x�b�3*�0i""ObPJ�&�,e���R��
`�S�"O��+�$ B�1`�o�sW�D)"O��S���&�\d�ca��WMlH�'���ѥm��E('�ݞSK2�c	�'�r ��39pЉۦ��0`�<H
��� ����W1k7F}A���}��i�"OL��ˈQ!�9��!
� U"W"O��it���j �R������"Oht9�E�/}� `KCI�*�*�"O�e�6�C@�<���x���$"Ob��m,8#�I'�<3�uR�"O�+���{�,�A���#S�DA��"O�M�Z$_�d�%��uΪ��5"Oʐ�e*�f����g� k&�!Yb"O^��1�E�����%(Y�R	�`"O,ȹ"I�:x����\3��i�"O<0A��I �V�E�^�����"OʽY�A�$U���W������"O���GͧdA)W�ܷŚhh�"O��'��0�I�`ΣODu�@"O�-RRGC!s�\�6FX�aJB�Ѥ"O�� E��q�U�N�`I��R1"O�@!����a|.=q�6`%h`"O,b��)���/Q�P`1�"ON��AGΩ,���I��_K�"�iE"OJ�Zk�2U2T��KX{�k�"O�Y�DI���3�b�9Ff���"O����^H��u�@9p�����"OR���Ձ��Up㟊e�=Z'"Ol܊���c�܉�B�F�^[�"O��K�1=�H�QE �+E�P�"O�!Q lθ�ZiHo�8�쀀�"O%a��ِ=��Y{2Ā�o����2"OB��f�}� �Tb�/�����"O,X��c�.V���0 �;��c�"O�� � 4p� ��E>"�b�V"O��3���!(�'?��h��"O(P걉@�y���Hc�-QIs"O��ᵯ��,"�D���T22�
T��"O6qQ4��i�:�Yq�\�J���J�"OT�����-d�mA ��.Lx���f"O΀#�/ۣ}�:�Z ��bG<�"OB����
z�hp{��x?�@�G"O�PE�G7;3>�[��P�2"O�t��j�	[�L�q�CV�d�L���"O��(�ڥ')��ZS��)>��À"O@���͝�7} ����ܼ ���3"O�� Ɋ
�ƀ;�)�4���C"O@�2G䜹=����p�U���h4"O:cb���ƶ)1�-���Z��!�$�
-P���v��%	-��w΍9�!��t��CV�<e��`�����!�$�3�<O͌�"Ċ|,��C�|�<Q�ˀ8h��� �ԗ��K%KUt�<�d!�-R�(�����v���"��Kr�<A���kƌͫ��S�H����l�<	���	Qjx�U-��F�ʹ��Lg�<��  �_t�
�횂jގ�����]�<1C�	�:�&5X�憀%����F�r�<��B���^=�W,��|xX"�n�<��'
�V�م���UF$@��S�<9�I�{Y���w��1;��Ge�<�$��,��X�ϰ}�h��!�`�ȓi��9
��A���DK\�����sih<�So�:$h��B��~�Fl�ȓ6Ahs�f�f��i���,U����z!�	��CּQ+�\"�倐k͠�ȓ*����PH��H0"��GS�p���/�Z!Ҍ�*Sk}1��ݐr���S�? �%�a�U7�܉ED��v,$��w"OJ�	P��4(���� d��M�"O����@�3p���$�7k`�P�"O2�B���8y��YZ�a"6	�l2u"OR�)�Dlf��e@�;Xʒ�yG"O@Ȱ%KYl�>dۀ�L�E�V��E"O�q����1'$!C���%v��0�"O��q�����幔�LkV�m�3"O
��PA�1��ptF
Jd-�&"Ob�#����J9@��>\���"O��� $P%kV�i��Dx�:�"O��f�� ��m�� 9
��v"OX ��R ^�h0����7;����"O��W�F�
F�A��/1A���"O�x�t	U$5"b�����/=7��"O��Q%X3
�$��U(ʹ#-��*�"Ob�y�J��cM�Q!��1R���"Ot)�#o=��3,��j���9T"O ɩ�
!_𸑳�
�Qt�I"O>8�v�̽i����*.�ʱ�"OA�m�0n��t�iH^�0#�"O�p�0i��|�zeQ�E���ī"O5{��_M�"����K�(o� �"Oҕ����l~D	�D�)Y`ūr"O�EQ/�:^��V��jn�ճu"O:���n�X�A���.�DhJ�"O� @N
F�l]SG��=I�lA�u"O*��P�֫p����i�����c�"O
�p�V?Y�,��膫v~���"O��
��\9l�H0C�hG�]Т�"O*!�gh޲T2�9d�5f$t��"OXH����'Vñ�H���]�t"O�@J��;%������X T"O|u9�C�e� h�$L.@����"O�A��ބ&�5�pB��M��"O$5����=.�"�Z��eh�"O@����Q!#L	�ׯ_�(�r\B�"O�,�@��ƹ�qɢve$9��"O6�င���}��\�4��-��"O6�x��Y�uN� ���Lr�"O�h����>%QB��w��H�"O��R�&�}]�b����|��\+�"O6(Âdآ��r�-I��hxJ�"O� ��DC�m�z@P��L�$�Z!�"O. є�ڥ+��؃R�ȥ��(Y�"O�h�%�U�_�FU���M~D!��"OԅR�,I!8*xj�%uR @��"Of�ʗ�mX�z�ыGFj�ؔ"O�qD=7��I"w�X�tӘ(ys"O#��,8�P���B����"OJI�gn_H����U(h��"�"Oڙ��L(lÌ �P�D�[�̨�"Ob�I�
)
�<����^=�B�"Oʴ��O"j�����1~�A�"O�-BF@L�^���&��*�h��""O, H��V�+@j�P3�0p���1"O(pQc�O��m�n �c#�� r"O�Qp!�>-�$z��C�>�e��"O@�cJ��vǀɩ�,N�:�2=K4"OT8���-��:d��:X<q`#�?D�$�),�*6�խ}R� 3D�@�snݳ$�rt��%q�8��/D��A�,
SU$0��;y!E;8D���W�V:B����tN.1=cS�:D�� ��)�ND#
OvY"�^�YA"O0;�`�l�V���W/^�`8p�"O����.�o TXRIx�H�Zd"O����Y}]�uP��C7V��dˢ"O0��H��~zx2�f@�X��S�"OŒ�- 40����Y���-0�"O�8`D��	�T �X�d�乹�"OJ8v@�	�p�H�#��Xh�"O��)��^
H�:ѣՊ&����"OЭ9�(F8b�)�BA^z��"O���G�A��T��C�4�b�H�"O���`-i�.�s��?iԐ@�"O��5������Z+�PB�"O����!��E�d�߇r��8�"O�Lxqb ���w�&����"O����E|g^��-"~W���4"O,���C6�,AiW�	Oq�"O�yS��N�(8\����M:��V"O\A�l� �Ra�K�.iP[1"O�	˴I�h ��ƣwށ�"O�ʀ)��s�bm���S� u:8��"O�����5 (%{4,�_��)�"OR�h��!!N��Y��J8��"O8���^�$��`V
/���"Ox$V	R�gF<-���'�"�U"ONZ���OT����EK�:��S�"OX8�2�S
|� �C$�r𬬰y�d�:�0M�e�.��IS�_#�yb!��y��$�&�*���,�y"nU"\�" ���[dބ�R�\��y�O�.?".�#��>y�}����y�I3�h�#�S�B��(��d��'��e"�I�Ne��k��Y!'}��'�@��V�=,�Y��5lXؠ�'��X��l��g�8��������D �',Z}(�.�+K�b�B"	B99	�'n�� �#Lj�ASC���1	�'��J�V�i��٥b�
)��e#�'�T�ʠ���|��R�K!+��0y�'�@��������sj �S)R��'qZ�0cbF$o�t��2V�>��p�'q �D&\":�h�C�4%\���'ؠ�pB�Y3+�|�j��ƻ,��Ij	�'y��h]� Y�i�o�!Ti����'h��qd� 
acV�[c#/"�"�'���b �x���(2�ڄ߮��'�$�C "��v��!���V:���'K�qR�%�4i���hqA��#xe��'J.x���aa&$@AK�2����'�i�5��w�y��V B��|2�'�T�*�� ��~���U-K���'hF\{��>4RB��舅;�D�c�'&H� BꟹV9�x��1`�
�'?tM��O 
��r�Ԡ%���
�'S4\UCA�_?�ȨA`P�rt�)�'[:�c4E�7���n��i�	��'�6*�
��pȦ�?_Mܬa�'}��`�ʸ{�LI Ul�/^ն�@
�'���H�M�7MK�2�`�f5���	�';*x�shD)�D��㈶]�����' �AP��U$W��=�%��[�2d��'��!Rd��UD���������Q�'1�{f���Su�1VC�G�^ S�'W"�B�("�@XY�!��P���8��� R�k��q�v]�A����g"O����8<b\��&�xxHs"O,�@��E�X\�1AUwo�Z�"O�|@� MH;F���NRY^��YE"OH0ME�p. ��"̊[o�,��"O��32�<n
�@ŋ*f=����"O-�v	X�b�:�R,�55��C""O���֣r�����̐�|xAi�"O����j������儵0�;�"O@i2B�:N��X�P#V�K�� "O��1E�N��hH%��|��D��"O|��(��%| T��x��|K�"O$1`fψxeRx	� W1	o�ܫ�"O:<x�B�.mܘ��:"����"O�TI�,)RQ���́;�r�"O�-
�a��B�0@�d"Q�P��9�U"O��a���A�NL���Œp>؜�&"O4�ZF��:BJ�Ir�Y�^(�4:"Ov�rS(=*���
��F�L��2"O�q�DɊ(0)�D+ݙ�B���"OR�(`�]��p��/o0�zC"O��h�F�0���:�g�[h&���"O���5�����pQ��0\Wz$c&"OZ)�'��-3f�0�wd�u��ʷ"O�8 vmM}���8���G�2�i$"O�]���ݷ]%�d
SA	%/��X��"O�\��	+��)�#���x��A�"OXxVe18&9x�.�r � S"O���&
�5f�T ���
�ژ'"O���4T�mhE�T����ع*a"O�%iU��R�p<���X��v�ڄ"OJl!r)`��x�$�ә(��1(�"O||B`��?�`�r�c��~��LI6"OH����0j={����B�"O2���zbmơ�&V]^�!"O�1�s%qE��!
l���@��Zo�<���ܕZ�\�+�C�	A� �X�ȔB�<�.ģv�r8ڗM�x��)�ӬJ�<���W�v�\$zai��z
z�r�l�C�<�CO@%v��p	f�:���K�J�<��H$(1�	�Q7L�#EjWF�<ae�H{P}�Ta�
��T�E �E�<�'`ڭ^�$�`@��%�A��C�<�0EѬO�f�(�(��w�����B�~�<!ԯϭ<��✏:6B�ס�t�<�s����xc�7v��yR���n�<��K��kF��G@ҋ+^����Gm�<a6��-O��0�+U�\J{B�Du�<yIG%2�.-�Ζ�'�ʬ
3��t�<I׭W�k(E��j�,$��� ��WJ�<-����2����Lߜg;0@�ȓ0u������]� +e0͇�/��k�@�V{���Ņ���ȓ:!� f��<XmP�1���j�X4xD@��L4+�dC�5|"-�ȓ^�,8�j������B��|PɅ�j8�q(�oT"�r��&-R�$�ȓ6�*tB$]/�v�)�(�oF%�ȓ�Z���-�L ��A�;����e�BP�í
=�Ȕ�pn[�C�޸�ȓ\t1��� RA�̱�a�4e䐄ȓ`��}	��V5�����=YE��mϒ)H6�:}Ҥ1'�r2D-�ȓPr�Y@��$.�Q��L��P$-��S�? ���".H�jx���9�6�@a"O�l8ЄC>���!�$o��(V"O^����~��m��T~(�Z�"O�;�� \2|�%	�m����"O`$�dU��M��b�*k�n�A�"O���d[:"��H"k̀ �  �"O���gU�0�T�X K@0k��;�"O:,�ǃ�(nA@ba�T�Q�(��u"O,�K<nrؠ�`�3C���X�"O�Э�B����[4hR:HcQ��R�<y5�Z,n,� �ܪq���B"M�<��c�-y�=8�̭$��x���SH�<a��˙K~�:�ŉ�4vH�q�
G�<�`!�� Y����"���	�oM}�<��2
�t��Ï�t�r(�0��p�<	�P�0!�̻�y��Hs0��s�<��R-^���жB�m1�+�KDq�<��N� 
��e� 4�,1'A�o�<!��K�2<!;���瀝#�@�k�<11��ဩI%���k7\����q�<IT"EP�Ç�ƹr�M�X�<���z��<�5H�}�Dp��JP�<aFl�+�l	�,R�`2��Rq�<�燔O����0��%%9��K�Lq�<Ia��/I&̻w��QM�T��a�<aT�0B.p�#lW`�Psu�NG�<�r�
-���f�b|i�d&�k�<IW�
�%c�J7�SVʡ���BN�<QA7M8Xʁ��ux��"�JF�<!�㟫7d�C���iB1��.�<�3d�>e�K5���G�I�P��}�<y%H˼���O�#=��D�v�<����1*D���*=�����u�<Qr�͹2RHݙp�9�]F\U҄"OdH�+��6LrEI�NA)b(PR"OX��C�aْtCK�9�4ě�"O�h��A�N@��I"�N̴dx�"O��a@���(X &�J�Xô��4"O(b�fصszE2g�;�ƽq�"On)p�ƀ��Yh������)�"O"@rdG�$;�؋U�Ȓi,�Iar"O689�nƱ\@��CՕr옕F"OxM[���r,��ٵdM�[�X<;"O&t�D�L�|x��mT�9�LR0"O~պǭǃR�tqF,œ4*�E��"O��j��N'x0$��ׯ%2`���"O �ѧ��$Mxd���,�*3���X�"O��SW-A�m��ڠ�*t�XhS"O<�0 �;���� �E2U�髴"O�:V��%	>����'�N=�12�"OJXg�Ӛ:E��5�� }$l�KD"OV�C�h� RLEÄJ͵;1����"O�91��2 ���!I�� ���"OЬ�1웴:�x�7��W>���"Oy2� �t�.
Q���-� "O|�b^�L�"!Ì+9�]1��ٴ�y�
AP��S �"l��y�A��yb H�C.��� k�M7~)�S�=�y��HQ��uDD5C3�������y�
Q+g��u�����G���q�y����-;v��ɏ�A��0VNO�y�.jp���Ū�6;|��Ĩͩ�y��۬
7&��r)�*+�����'���y����^p������ %�:�#ԠC�y
� t`�r�MB4��ѓCo�Ex�"O.���(@�PY���Ξ0R�hc�"O��ýB�F�.͆p�z|��"O�s��^h4l3An� <�e"OR�q�MUq�X�c%M��c����"OT����M=N�����§+](��"O���f�;9���Qeıl%�t"O|��Mv��3s�F-V��L�E"O��iELS=D��2!�Ƭ4S��1�"O��NÀC��H�� /A���u"O�tZU�:1<���OһC"�@��"O�sᏈ�QɊ�5җ����"O���N�I}��ڢ.S� X�Aa"O챓 )X=a4���k�(���s�"O���qOV�qظ1p3j%GB����"O~� 3� �lr�ܫש.l0j�W"O��@�嗋v������jм �"O�]��Lܟ��� �
�3����"O�8��I�Ar��ʁ%�^�Ε�"On�
��3�:��恜�9�8�@"OJ��I|9Y���@�e�"O4�s���p�`P�]�H| �"O:��� ��n��,̪3c����"O�	#�J\ uGJ�saڡ �ܽ�u"O0,�6�$*�&UՀ@�i����"O��s%�[�EB�P�f_�85Pa�R"OF�ムʈ^'����h֋1΅��"O`��O�:؝ꠧ�b�m� "O��`�ʁ3��)jf%�%*��;�"OB��Q@�Bv�q���Ak�,i�"OR�j�Gá\.$}����#_W����"OHVf�B�[�-�<���d�8!���vB:s��ЗOGp9���m�!�DM�VI^@���)S$��a�ߛ$6!�䇵�h��B��(����B�q%!��V\:�;��"ӆ$���T�!�Đ�4<�a�#�">� �7��1>�!�$�#��8�X�l�ƌ�3퇺*2!�.Dz�r�K£C���30�߂`�!��w1�0@cN�:�ڍ�E�'y!򄓵&����I��>.&����W+u�!�D\� 'r�rM��zܹqH�y!��C�b����6w`J|@ЧF�/�!�M���Ub#�FNP���S`!�W	p�D��N"E\�[��K)u!�&oLڀ�q%п.�L��JF5QI!�$
T邵K�ǒ^#^�c�+E!!��"1ɞ��$��A�B�č�� !�dòm���F-���!� n���!�ʨ9t�#c��%�	���J*�!�D�"�a��n��L���p�!�d�D����fA�za|��V�@�!�$�>@Eh�Q �ʱQQJH���$T�!�4VJ0����2���F��OR!�DF�(���B�3:�h4�󊖶im!��%it&D�%�ΠM 蜸S�ݜ5�!�$޸7:��9֏J�Fp�F'�|�!�G&�1@��]@�2��t�!򄀠)�n��2���R�L ��eо
!�$�1HV�R���Ej�2D%�
�!�D��`��9�%C.*�*�����!�P�y��Q�R@\=F�@���;3�!��`����%�BP�k��P��Py�Q�i�V�k�dԷ),I{�F�&�y
� �����ƌNmA��`����"O��+�	�>��*�,r�"O�`x�	9�dp�Ǯ$~~�Ɇ"O�(s�O
��婒dͪUb�U�1"O�-��LL'Zl�-9� �"ugH4�!"O�Yp#	�O�jT��o�<_-�7"Ol������D���XB.ԕ0�"OB��a��(s�P��3U�v��"O�!x�f<f��$Ѕh%;W"OvE�ݕ��w@J�*�~���"O^"�e�
$�5 �n#F݂�r�"O��(�-��m4�!�r��h�n�QG"O�EB�ɱpX��tj.]f�
�"O �v���i�l��(�,Xl�H&"OH J&`B�v.f�R`�%P8�p
�"Ox�3 �ܯ ��05�_�J&�)�"O4�ӕ!WKǮ�s��f��S"OL���
DN����D[�z1i"O��B�+�7�JIHS�]&"� \�#"O���ԩ%s�&��@�K0ip"O�t�R�Ֆ8o��yR��S޵�"Oޝ�rOR!`�Lp���jJ��1�"Oބ���1a�����b��F��Z�"O���<�P�νa���1NOZ�<�ǅ]9���Fٶ<�,pI�.Mk�<���%9bt��c���(i�$Fh�<A�f˖Ͼ���D!��<��.�<����Av����-֛tc(	�u�<��(�;C@� ��1Vp�V�o�<�"n�3'lɣ�C:bG�mس��t�<ѡ��#����F׬Fb9@!ǁZ�<�.�<]��P�m�#l^�ڕ�X�<dŚ!���ڑ�� [n:An�x�<�h�W��E1턪
<���N�<	�)�l�S�Y?H ��,F�<A��E�:�Zm���,��D�
�}�<�dF*�l����S?�L�bU��w�<Q���>�8T�����2aR��Mo�<��)�,m���yW�$�[�琴z�dC�ɷ Rh��cV 3�tC�C�+v!RC�	:X�>��5 ±hx&�(%@4u(C��,K��r/��,`�ܩ�%��hBB�� �\�g�H6��`��=�HB�7+3���w�k ��PD��#�B�Vz2H饨��\�I�% WC�5���S��]�Rj����)�5Z�C�	z��@#�C	POf��-k�xB�ɇLH���L�s�\�끬Nr�@B�IO�:�dg��wb����	�<!2dC�	�#�:�Gm�'��%R�H#U�B�	���XC�71N�E�b�B�	�q1����`R�Q�R�³d ;h��B�I�e&n8P��!O9`TCĩ�pB�I*�ڄ��O�Q�>Y��çP>C�ɦ	0ZT��N�7Bb.� ��+�DB�Lԡ��+	[F�����2�B�ɷ@�1��lC�ݨ��ɀ+<�B�� fجb)�J��idDb@jB�	�)���`b�=p
4¢J�F�BB�	�^�V�a�	�y*Eg�T�dB�I�nL�&,G<��P��Ә��C�Ɋ0r�`8�/���H����?p�LC�;rY��`'B�Z��V�Bg�s�'�p3Ԋ[[��@2�Ȇ=���H��� ���D�عQ��tC>u�L�+�"O:�Hg	��{�n0ɢK�*��i �"Oz����]"=窡b��}QrIq"O�E��i_0"Y�Q���5y3���"Of�)0B�1�� r'"Q�@�l�CB"O��:�`J��d��0؂s��Q��"O�}���	t���S�2�l]�!"O�I�h[,X]�27(��U�����"O�Da!(�Sw�hr��^%����"O�cDdTM��=I�\�g?�8�!"O����Z�6Ȕ��	"x/����"O8��B5~ЙTBC�%py"P"O>ɀDD�8��i"���� .[�"OfI JJ�O��t� �=LL)�V"O8�Hq�L�{-z�3�oL� ��,*�"O ��Pa�;&��)у�[��1�2"O�H��Yf@���3C��ё�"O(}�B£�RI�� ��Se��R�"O��σ�u!��F��� "O�I!gC\�2��9�m7����R"O�jw�X�XP<��< �&M��"O��դŴp����lۿ�8\�"O�Ku�D<t� ܉���4�>!e"O�#�ڑ"��[�dX�$� ��s"O�ܡ�NV�#5�BI�|�8��"O2 ��3M�@F֝[ ��pb"O��Jw�L� �ą0�BˋA�0���*OT�S4M��s���`�Z���i;�'= �	�I�*�ZொA/TI��'mJ�"/��6����g�Ӽ(��E �'��ab`b��h���V��-($�q�'{�hat�� �2�
&$$b ] 	�'��2��S5rXp�1���e:�S�'Ɋ}z��\�>���97�'eOԤ+
�'�8�'$X���PcTYY�b	�'��=��ǘ�{��ٲ)��Q�4��'(&�0�ᒕSfЉ	�7O/���'n�WmU�.K����*Dn��'���H@Z���c�fI�d�|i��'����r�r�L�P q��`!�'a�鰶�
P�� �E1b�@��'E�)��MD&�TA�1*~�m��'K�����"<�ƈ�c]5%���'4�AU���4�D�bh�	�'���Ae�!G%�|+�I������'5��դ�qr��C��>����'�p*� A�l
��
�^����'fT��4�A�#�0]�!,:�h��'��x��c���L`
'��l�<UX
�'�%C��
.I��H��OGk�$h�'�b�,�$8� pU��
�'�
����I�:�8U�7
	�갓	�'��P`$A�;:�����jF |�:���'j��.i���ϋ<nw�Y�'�
hc��D'𰱄ǌ�޺���'�t[��ЌR��5�q/�$��)�'���2鑴i�����<4A	�'P|����Fx���{�G�$
l�*	�'�4����(Ƃ��G(�_�k�'�v�X�c��f�m��-'����'�ʭ�)*RV�=[�`Cw�zIs�'����RY0�a�iSsE�x�'�$lA�ET-Ѐ䃥J�bB��h�'�@9��S$��B?bI�i
��� ���J\*J��S˓�7�(M*�"O|��!�HBzH:$)U�(�N��a"O�tpэ�'ZS edH@�/�Ls�"O��������"�@�b�T�1W"O�D*7�X 9Ȧ�����fzp`k�"Oh!�F#�>��e
�*o��V"O~�k��:K���9`f�!~6�"O��k�~��m���ca���V"Op<#�V�P�,�b��9k^��p"Ohx�'#)"��!�͛MG��K�"OB�ťZ�cm���bi��bP�}CF"O�(��l�pφ�
c&�2KE�Es"O��)h��9��ؐΉ?�i�0"O�Q�5Ɂ ����C��*2��"d"On�XQ��� Q��
�2���*�"O�hK�d�r��-� f�	�2yr�"O:�9�L�) ��H	�����2��"O�8�cL�=+���
5� j1"O(AP ��Z�� :�,�:v�(��"OtE(�	p�~͒v�׈5b����"O�ȑ�n�1��U@iO�j�H��"Om�g	W@t�h�!I�BP�xI"O4P��Ҍ1�\r񍇓wH��Q�"O����M>)&�q�,ō1FV��&"ON���lɴC$�����9�"�*Q"O�X�C�/h)�P���PR�j��w"O�(�F��:;H%��
��jPպ�"On}�*�X������MULQz7"O8��e�#=t��sM͌:�ܫ�"O�u��^��`۳Kɇ)4 ��"OF!� �qP�� ⪊n2�!p"O��B��V��=��%4���"O��9�m��vN�,�1ĠI�e8B"O4q���S�l���A��5^��F"O0,{1#ʷ]7��	U��;9J Dj�"On��c��{<`�;��ɱ+3Pl,�yrm]�Ԑ'�U�<���`��y�K����1�	�5�JJ�ԝ�y"�؝@?�z�㖊-1�QHÁ�2�y�	Z~�RQ6�P �R�T/�y�!�e�.��M�T��I�e/�0�y�( O��aÝ�?��,R�NC7�y�A��j���
G���5��h4iZ�y"�\!\_ �%�5��-����y��e�ָhw�/*	T���9�yRE�#���G�w"<u��@'�y�K&D��S+=lp)96J��yb��;t��A�_f�v�e���yB�^�i�&}D��d1~=�r
̬�y�����x{��]�Z�贲��X<�yb��-+�,-�W�N[(�ca�\)�y�$�,dR �M'2���ȡ����yBU�j{�9j》�!�H)�i�5�y��0]�@U�
1��x*Q�y2c�Q�X�*>�^ 8��H��y2oL�{����g�\�2W��J�C��y�މQ��A����!��mzs�Z>�y�q�ܱ��H�XnȲ�f�,�yB�P�EB@��^Lny�r�І�y�-��qM�Ě!��(�Xg��7�y�iB����쌓u��r�d���y�GN�K�i�P���t���s��y�H�ƈ� ��B�
�4mI�y�J������R>?��"t⋯�y
� h�4d��
�X�gnŚ1�<���"Oȡ�4,��5S@9�͹bʔ 0"O�k!��2̶`���[t<B�"O�m��hƑ	� y���"U�"O*�Sr�+s�i�@ֲ����"O�Y�nߓ&� AZ��Q,��L�B"O������_�\5�w퀵QQ�,�"O�#��^�o����S(l�ѡ�"O�=ᢁ�]��e��+#~p�F"O�T�����n����>^���7"OX�r*�G�5p�P�,C��pF"O"�A#�W*̲��
&�*�J0"OzHZ�P7!� �(A����A"O�����:.�� v��+�Q�"O,��L �/��I�F��6��"O~ ����'Nc��Ig���`��""O�	���&nl �)<�)"O�A�Pˇ�B�t�e��(�0K#"O���OF a�I�P��+%
j� 7"O��P �S+p5C�=�4�SP"OR����>.���D';��$�"O\�S0b�?c\$IZWf��r�b�8�"O���",N�4t�q���(g��XZ#"O|��0˒#F
l��R�&�i+"O� i�!�_��;��8iu ��'"O �	O	$k�5a���~k�*�"OR��k�4q��	8&��5YrP�%"O��#�(R'�԰��+A��(�g"O.-�ԩ�4�9x��,B"OB[�k��RE"R�Y-����"O@(ѴaV:Cߌ�a���2F�\P0�"O�}ȇ$ÒhC<$��ZW`���"OZ���
M�t�p���fO�Sm�H�7"O�YX�C (����DE*I���"O2��'��!cθ�r�C���v�+6"O�-+@�Ɩg9p���=h6l��"O��� c�a�|ȃ�@�|v�-�"O�XO(	��C$MrM+C"O�kt��!mn���/ērAa��"O6��b����Ui���� ?B!a"Oh(�@mV�Öjr��U2�)�"O&��Fǅ#A�4�7���sP�A�"O�a�U�D,I�)h�$�Nz��1"Od�O�/i�De�c$�JiD�j""O2h���M�.TU$�0>�`�""O�- bɟ�Xi�D��c�@<����"O� ����G�y��E�l�����"O��0�;T6��Aeމ/X�!�"O�8�o�]�d5�@N�Z�@�"O���ŗ�:㒝��GI Z��L�T"O�d��k�hC�P�f��h����r"O�ek���&�!�S$�x�~�X"O@���<b�8� ���>��+'"O�(�"�>[#��)r�Q	pkx��"O��c���UЫ��s������N�<i��o���Qc�U�2��IR�RF�<�$,��#�2	bbC���M�Y�<����r���⋗R��Z�R�<�P��-����{"4��"O&!ВD�&��A��cK�4u6�k�"O�T�b�lZ~��ra&�`��"OPL��	��CI�����ot��"O<�ȅ?bFN�jk�=:�4p�"O$�xA�B�r"-y�*��O�"O� �	y቎�;X��0�	�[>j���"Ob��A�)3�)��LGn�2�"O�{�ÚaLr��s�hl���"O��A�'��3����P��J^��"OFT"�eឤQ@F�EA`��"O�T�'��
��1 fK�+?t���"OJ��Ш­1&��ҕ�V4d.�m�p"O�$�#�O8�T��#kI�x+
�Y5"O�-�ԉ6V�F�Ŭ�+h*�d�A"O�9zu���	U�d j�>���(�"O��9Gł8�����i�	��\��"O@)��?f�Ȅ)�&S���3"Oμ��^)R�B���%���:�"OTx��$�4L��@�=Di��u"O\�(��m�bc�Z�K+�t9T"Of��k(30��$o�X���"O��	�A�g$�M��O�5!��Y�"OV�����"�F�PvG�*~�d��"OnPsg�y�M�P����: "O��fcӱ�]�c#,O����"O�m�wd�?J��0m�&usE"O&)I%�6rך "���H2�I$"O���Ãb��16�Uw%vh1�"OL �#�yB�ݙ�&\�.2��0�"O���n�%���S�D�i&���"ORu�7��%16d��R�=%bm��"O���b�����d�)m�}�w"O^���-Ofl��Pu����"O~�ꁫk;����!��^c�@"&"O(�a7K�+Y�0�`�@YvC�X��"O,��p�I3p�F}	 �W=|���"Oi�nCF����įϗx X̛C"O�m�!�
���se�E�K��"O���&��7g���A�@����Ey"O��J j��&6	c��K 1l���V"O�z�N�~�<��'���|OHɫp"O��y���9J�eSe�W�8B�岑"OP�òo�z�\ �	/���H�"O��2ʄ���c�cDs���
B"O����
4�z���'�q 5"O�]Y��e���Bd�M�d"O��A7�=z��i2`�Uv�s@"O��#s�јq�r݁R��R�(Pr"O�ze-
H��q�ᝯ"٘��G"O��w�o��0s`�,/#���r�TH<Q1C^�q0dy�mI#9Ŧ��4eNo8��Y���޽%a<т"��0B�2 �	�Y�!�d�YeX`٧�FT^���OR���'&ў�>����7�t��h�J-�݈C�7D�8H�B&%9�dJ�ȇ�\��
(D��j1��� q��)J=Q��/'D��he"�	��ph��Ɓ�X�@q�%D�@�tb�x,4<I��'YMRY�W�"D�d�� ט�)XlQ�4uX���>T��+���)���3��s�`u��"O��SV@����t0u.��`�t�Q"O$i�5��M˰� �����0 FR~H<���˅�ȰWNһW�~+7��lܓ�hO�OI��i&��7�f�K�
T䒡�	�'U������Ap�����"E�P�H���(,Op��ňR��Y���ɒD"O� ��*��1� �@C�S�2��8�DM�Px�mĹah��;%dJvE���'��y�"H�q� ��B���`% �G.�	�y
� � XG�Tagz@I��	j����"O��� h�7MT�م!�H�����"O�M��֡_�"�J�`�5O� �"U�0���v��i���lTT�����E�B�Ɍ/`��;֤S^Vi �� �fC䉲i�rTPnĎa�y:7)Y�y0C䉚$��(˰��B��:�o�jf�B�ɒJ�V���'�3c\�����0H��B�I�u�L����b&�D��ꇚk��B䉽=�Ĵ(�	��Z�iFM� 4�HFz���8p�ل~�����G��Re�!�7D��Yq��	kj���\�j�a*�cy����<�HOP��#u�۞s+��sS�#{Xͪ�l1lO��T���W�^�s�
�;c�C�b.D� ّCY&Gm�<���#:�T���7��#r��>��K/l(�w���Tk��C�n(D�t��M�` Z\�>03n��p�+D����N��_6�L��ǌg>Hv@)D��a�/«Y� ���ƍN�(`/&D�|Єj
�]�y�%� -y��48G�'�O^P͓���4Ð�+tl�' ��,��e��T�c�\�"���� 1j�P��� ����ݧ/��C�9Q�4����O�$B䉦����QΔ�,�hy��J,o��C�	��p�!�Cؼ �s�,:M��C�I�j��@h�Ý���$�I��/��B��G-��1�e]�JD@���
�"B�I<S���1҇G93��<�j&"�*B�5-���C1�S*q/��C!`S9~��B�	 c�
9gͥf�Pm۶G�C�I:}��3���\���[���?p�B�	�CH0� ���P��5c�Ü=M�C�IB��	��,^�&E9w��X��C�I�H�m��D�&Z�Wi� ;~C�Ir��C�N��n�r�;em@�p�'�a}ɒ!R�Ĥ�1�R�]?�넫��yRi�=B��a�B+O���� �y���tN�%H1T����Q*F���� �S�O� ��7T���c���C��Y{�'��6��s�l�B.�1k�p��'�R�K��nIdC��S��(�}2�)��J?����M��t>H$;*<x�!�D��3��6O��Ƅ�w.���!��aU.����'�z�!CI��!��1��XS���1�}A��<O�!�G1`�� wo aba��7x�!�$�4Ԓb��ˬlO�8㜉o(!��N��U�jƣr���E�.!��o�\��ơ����%��T!���J�Ai��[�./$}���4�!�dG0do�tЕ��) R�Co5�!�D�}6������8�U���O�(!��=P�����@��L
b/!��W)7�"�;KY�:��ǄÅ	-�OX��D��J��|*eL/;��9c @�ўS��S���=��
W�昊� ��4C䉺k�d܃�e�5�	��F"P�7͘{�Bl�{���i�ldb�C�$jH5�!��`�H�C�'��Ac6cG2h��˲��]�Z���Ol�2�OP�2W ��xص�Y#��$p"OZ͠q���#�HH�i��i���@"O��s��Cz�QiL=c�E"O6Q+ Α�'���/O�\Q�"Ox��`�2Z��@�j��27� �"O� ����=ShtQ�)I9D+�u�"On�)l�	Q*��wp""O��X�&���eېƃ7U $}	V�'21O:���G~� r�5$��A�"On����M~/�����N��~X��"OTM��kۣh[�xa�dl�4�E"OF\{�ũ�0�Y����D);�"O�)�Ө
�W�Nm��!�xoʸp "On9����\DB0�j�kk6����'N�'�-�k�&q�X2$K��>3ݓ�'�"XAC�̠s8�z�MB�*��ua�'��B瓵>��i�%�r����&�y��˂>�|P۴H	pk�r�P4�yn�=$Gȩ{F��Z͞"���(O<�=�O��������Ɣ�C�2b����'��2�	�5:��b�$VI��'��d����F��e�N].R=@�'�,�1��^���q�X�)X�<X�'������%y�,t�M&#n�-"�'��)���r?8�eh�o;��
�'Z}x�넫*4�	��oN+e�N��	�'p!�ЅVv�i��!V��	�'6P�  b�7%u*�s2�>������"O�M� #2c�Ⱥ�JH �!�"O���w$T4j�<����L`HJ6��)�S�;��A���&�i�����C�I�s �)�v�U)sg�H$2�C�awvXЋЕO���6A�"#4�>���i�2�  ��GQ�ZuDXcdI�o�!���|�z�����\M��9Si!�D�:U8�pE�ZCظ�# Q!�d�)d�pA�3=�,����R�HJ!��@*-��e��$X�7�p�`�ھ2ў����	_��9"��Y��C.;�.B�I�#����(�6�!�.b%�B�I�X�jة֦M���%Kd�e��B�	�b�Ĥ3�,A˒�e��1��B�I \��(Ca���N�:���ҭg�B�I�>$�ك�ۨpYB(�UL_DXB�	.'���C���n}|�dB��	]
���3�H5*�ͪ��M6B�*2)�|��%xD�cTJF�s~VC�	�$��y�Qm\�"�S�^��HC�	�u��
�ʆX������1�bB�I�U���+�&��\Y���t��j>B�{��]�4��Xy�gC/4`y��@s"�i�*ʢ�HG�l�8���-tL���R!:$��O�QUM����A�q޺�8"�#A��ȓ*��@�u�L�7�y�L;>	����l���Ӈfޥ]�~x(��8D]���+0�����(���R��;I�万ȓ[Q`�@�ZUk���#l�4u�Pm��6��PX�* k"�8��P/�R����ax"-݋W����u(_>-q����R~�� ӫ�
v�E�R-T7j~(��ȓs�NC���e'd�7-�|I���ȓ
�� ��`��0�$b�#�섅ȓ_4��x�F� �3���1!���'¡��-� 8���BDDK�\��%G���b�~r}�s���>\!�dŀ3j2�	�D�p�z@H��`P!�䝋"�� h�'��p{���T���!��ɟ�Ę� �F>Uh��P�N��93!�� .Pb�G�^��e��.u:|I�"O*��#đ���=���3oLx�"OVx��Y�nT���&Iє0XN��V"O���S�@�s*^�ڇ�Q
-�^�8�"O��(��3Xd�V�Àv���s"OYE#�+ָ؅�=:�, �"OV��B�1��5��b	���;�"OF�	c3k�M��'9���{c"OrT �c�"i�"7�Χg��49OX�V.H�u��@���M�lhX3�����iDnS��������~�,C�I�pr�
��'~`C�jU8�"B��.6�@r ��� p$q�h��r=B��$WL��w�e{	r��gG�:x��C���3s�͙$��uk]�sr�C�	2'F�ȠPG�-\;I�\B䉱|�BC�H�E��)A�)X9�|B�ɯmd(�%)��Yȓ�*&BB䉜M��}[�`�s��ac�>�B�ɺnP�(A��ٝm����^W�C��=K�t��f)rV�:�J�m��C�+I+m�pdD���5��T4Q��B�	�/�ا�4nd��p��v��B��,FFj �rA�il(����=�*C�	{/V�Jf�Y�j�~����B�	�g�<��%�3,NkS)�il�B��	I� ɰC�uS^(���J�l�B�-7&,�C�� T�@0	���*;? C�ɐHXX	�D��8`�� �Z^0C�		2�2&k�	Ӹq�0�S>C�	�]��@U"���b)�R��19��B�I,�ƭ�b��Jv	Ks�?��B�ə#�����K�J�a5�IrC�	�x'l�ؕl�F�����K�y�2C�=��8����j�  �_@FC䉈8^B�Ar��rrTY�G�*"OB��0f��=�$Ѳ~�2����]P��	s�kX#C%㧞��G��'_Τ@"#�o�"U���d%60��'��`kpbW,
^�Ӄ%S�f�3�4mH��A�
|~�h��'L��e,3���؁h9<t��E&n����)v�W'D���%���|�+b��"S?R|Rt
^[Юt� ��?"�z��Y������b
6쌠E-���'4꜐5��QP��	]ct�X�rN��V���T�8qZ `�ј��F� Ჵ��G�A�<a"ʜ.<�(�2ǄW?Wju����1"��͊㫓�wDv�C�`�&k.SB
/?� �"��8A�xޥ��� �r�2+��I�.l�94��Q�����[��ݓ?��a2j�)G����ٸ3V������%�ȀJ�`������:	�'Cz���Y�:s�	� ��$0�t�)�"&n���x�4��積�[~�<���u3(������<�p� Q?r�����I�]���
sf��'�~P�U�]>I%[p#ΚwJ�x�q*���$��;l��RE�+�~�:'�B� ���\�,Q|�������Lɑ���&)�	H �>e�,eP�/*���7��A��A�Eǚ����$8{JL\(D��"Sn���*K�TD
�����@��q�%Gں�TD��I�`�]�, ���_�;	�ҵ�ˌ�p=�g����|˓\��m'�V��(C�iOd�����x���͔�1�p��f$W&F=��a]"]�R�B�Hƛn@z��OJqÂ�+6a� %�ωT�
��c�d�+I�N�-O��)RJ�$9
'��$aFK'+��e���SDt�@�V��r�h#���>Z^�) Ni"�!3����n�	�`� _ Fm2����!�<��H�P.DB�#�oO0���(�VT��	p%�%=�]���Ѐ#Z��bp$�Xx\*0#XA- �m����X��j�gh��K+�T������Х��&טV��-D#\a05�]�W���s3K�)^��C,k,�8E��1�
�M��e��ķ�$`��	Hω'�jys�nǝ{�]j��hvv���
��"�d���G[�5غ���G֊�nuS��Gs�y"S�Jn{l���W���r��.ta�)�3Y�����	�y�0[F�Q~�>V�
��3u�N�(X��k��2**�U� J��TX�(�rE>!�t�2"�4�Q������A�&\ǉU�JQ���9�	�JW�)Cc�$+��i��n�(M*$�ڤ�\01�e�RF�mTr��T�4�H����+nv�e'�O��	�Ɯ��yj�s�- A�i�֔S"�0l%Pa���;+6\���L�0+4)���Tz#�s�� �!	6��3D���R�Z�WDb�"O]Ci�2u:.a� H۲GO�Q �n�7��+G#S%
��d����K�6����rZ�ɞk��	�� x���!��Hl���i��M�5�"t�!��#�&t>�a4GէZ��X���}2l��B�CzZe�����ƬiH��,^�	�J��?�����C Ta�d��7_6UbN@�lCX���aaЙ�MR�zQ�٪���7i[HH��	�?��������@����5;���#���I^�lybEYGX�D��iK�!]K���OF��Q��԰B�D��v<i��
	�'EX\2ѧJOv$i�M��Wg���$��p���!�P�v}re&_���O�,��o���c�� 3v�����Xjɑ�G'��) &��x��r�#ѰyB����);1Ɣ�w���6!×$N>����cÌ���O�q��C]�J-�	9����u�>qc��'d,��V�U�S��	�T��a����!�S,j��O	Q�1���2�$���&�O40�[Eе�C��;f'M8N։'	 �,�s��uX�g�-�X`�������'"��0�[�&XhH��Q�6�*B�I�*�H�aKE�P6�="�V�SQL̘�!%�XL8�^�0bE$��,��#����OE�)���,g+!�$]>F?8G�/
��`ʍ�U��{�c�qpV��!P���$C��'.ܴ�%o@�#�*�9m��ד��$*Λg�6�`���I�`J�X�>���PҨ5|0��
O`\��)-�0c#ىE���V"O��9����&��!�k:��Y�"O���W�~H�QI��-:���8'"O���R�X3eE��� n��5�4�a�"O$� ��Z	k*�h��8r��F"O����c�4	�`P�L��r�N�8u"O*a���[�1���_�Y��y�q"O&	�j�Fs���!ǃ|���yg"O��[t��g�`��g�1,�,�"O�\�a'ЊQe���D�+i�!K�"O:��V�GF�
�]' ^��r"OB�f��'CRj� �s�0�"O���� �,U� ��ʜGޠ%{�"O��`P-?w�n8t��<I̖�b�"O����̗ a��էP�/�r���ƌ�.�t0FX�Q|a|b@��x��E�&+�2������0=17%��s��Mz����?Y���8	�8 PN��Z�`չ0*�y�<9V�1�UôJ�l-``���Kx�	�m)jx��c˹`�Da��S�;�l ��< 8��1b�"2C䉸"��yʴ�ΒE-�
�5 4Ɣ"�\&O��<A��'�6@30�,�3�$68�>Y���Ň{Z�U; ��*h�~�J ��c��s�x4�ȉ.tJp8���4���h��F/���r�dʹ�P�Z�w�j���iB�
,=�$o�!\���B�hOv|� F�J�<���hV)=3����C�&�nդ�\�����l�>T�9Je�ˀRI2|�5�|�0�	ۓĆ����>����A��(�9PLH�~����Kʘ]L��PnPȐ�ɇ/?����!eE)�p,�y�(Ĭ�D�E�1*�%n���m�tY�AM��-F�2�H������6�V&۔`�"D-r�b����n�zE�!MȄ(L��������λq�dlk׉�-
�  ax���I��m��9~5��x7�??� �Z�J 1^����Ou������R*p�0����)(���L_�8�>�2GjAs�I�a���x�!;<Q� Q��
� :�o��Pq.ͣ	Oh R� !4��9R�lՐXSd<���PJ����+PqѠuӅ%!N1	��A��h���SS��@�Յ:�lh���"?PA)uE��'�Bu�S�Ǆ�B��ԗU^��(R��<�v\��o��9HeyE%�*��J�y��mX&�8�����'�z�G�Z�{��)�7j�=.���*I#}�!���߃~�����}�8��Z0z����
�*���RYc��=ȧ��0���*�����hɇ�,lO<ѻRA��)�ƭP/!j8�\��`ڟ�H9�W ԸJ�8Y��3O��yы�~	^��dmR�o5�`�"��V���5}�I+��[ h��w~��f�^4��'A�ɘgM�>"�v�Kd@�K���i�dڎ}�^�j�aJ6��4T�S���1�+2+�rv�R�M�^�a�e��֥:��'AB��c�!h;�,�Q�B�h
�m�V�T�D6�,�F��?<8��Z�mJ\�St㏢n6����o�]��D�8CY�q�FC#cU�I�0�ץ{B2"�e�g(<��A�#|�Q���',�4�sІ_(�'��%y?�Ix��Ȳ<�u�E���x�m�gcZ !���+���Ԉ�,%�|c�
0�b@� a{F�=5D�$�� 4_A�'N�{�f�
��
�T�y�G�>r�љ��V=q���� ��puN�[W��~�p�K�j\���� bό	.R�qa�@��1�>90�.`B�sbI?6/�T�"$�b�jf@İ?#� ��X��И>� M;�C�tHbr��2�����7T0N�	� �%�p<Q�(͵�t�P7&�25|p�0ɝ��u�ŭY=��6���:PJ7�"7�DȪ��c���0��p��M�#����7+B��Ā��UF�8� 
�'y�q����o�\:���)�Z���G�f2���@	$@�ђ�ļNv��Ҩn�tz4�В*�P���gu���A_�l:�
&�i��P�X���'9B�����.)A|�F�c�~@�u��K����dV�nh��AF,�^�@��u�ǚ y��I�0��[� ݲq񂃁�2I*Xᣌ%+~��@6�K70�q��e���M� EO���U��+Q�D� �&Lr��w'ڼR��h��E�5^YzP${s�ɇ�I�E�(i���~������Z8h�6�P��R�����\�n��D�G�8A�aKߋy��ݒvn��o� �`��g��TX@	����ŭ�(�`�'�T�Is#3`�������b�4���44�)3�쎭\&�%YF�B)<�N��Ù�b������c�6�Sb� ���$�+���rT)�2s�FȄ��03�!T"ڑ<Y�����ʤ��D!{4�1�#E�=�\�J'�>����?]�tb�U��M��e�Y�8��TS'G�%"�����$dy:��v�ȸB�(Ӱ'X9uT�ؖ�����c�oʰ	r���#��l��y�ΘT���Qj]7��(G�	���O¨r�mL	Q�L�����YK>�K�*y��h�p��*N9�����_4>��-��p.N8� �5>dq�PeR�#'P��'�踥�J���p���"�y��-3�:��I����əE�!�ƾm
X�P�H�sC8Za(��t�`��� �	G��Tm�C(sծ6�3�I*	4���K|�����yz�C���h��!D������#2�$���F�@�Y[����L�^�����04�C@�_q��S"H�	�!�d�]&qb�N�3P�����J !�䕜
�i(�ꏽc��̙��^!��:Yl��$>I�r:D�L0�!�dQ�`L���%P�ѱ���N�!����@�P��Y;j�6p����!��	%�q��c�"m��L���!�o
m�M_�@��Y�&AM3V!�$�,]�Th ��D�� P���
�!��K��ph
�j@ <�!�G�N�ʐ�%�G�;��hy���!�$^�_��B

 ��͡Ǭ��q!�D�J��#���U쬜�T��&�!��rơ�4���ؚ��G�7=�!���!.~xQ��"�~���g-J�!��/\tP*����h �X�Ϝm!��\ ��=�,J�:a�t*Q�}S!�$V�S�����1a��.��Bn!�������(K*��°���YS!��:� �j�s��(�Z�k0!�݂�j-�4�ρ%a��sJ�-7=!���2�p$��j��A�)֏\�!�آz`�����Q2PD�
9E�!�$�7��������L��;�hɌQS!���X*�G�I�k%ⴊ5G�[N!�ĉ�2�:��P���)%!e��K$!��k'�����85���B�'�3�!�$Z)��M�s_���B,�)�!��;���Y���A6�I��,śP!�DH��^��5a*X\�uIs���wV!�͞4���0��1LƝ;�%�+G!��C�m��r)6~� � 
s!�䒲;��F�J���b��[��!�Č�!	"L�3��G#�upb�^�!�-2�� 'ֽX�G'�!�$C'Iެj��Q�#�W�"��q�E"O�e��hq쀙���?&p���0"O���אW�
��E�Bb\�C "O���"���d�I�	Ѕ"O~ y���,KJ��!��$vG"T;�"O�����(  H��c
]Ԝ���"Oz�'��x� ��`?4Q��c�"O� �� �S�_PPaP�.Kh��8 "O8��G6&(�ʴa���lUZ�"O,4�G��A�hbD�̗6��E!G"O�L3`ć�_��$�q�
�R�p"O��z"g�@u�pz���94�*��"Oʴ�Fj�.�Lt�T,זV�(|z�"OBYvlZ<=~�5*K$�tL!�"O�(��K�7*n����N�����"O(�����5TE{g��e���"O<۵�-��9�f� �<��"O�	kB��e����v���S�(�Bf"O	��oD`]��[q��Gp����"O=Q1�	-j��Ʈ))l4��G"O`}��"Z�n��sb�����b"O�aB�/	1@�&��b6Kf�0["O^Eɠ$��2	��+F+:~���"Oh�Y�o]�F���䋖�vi��+�"Or�K�^�V*���;U�
�YV"O�q)��ǨS�%�����Q��Y�"O(�0���R�� ��dB�L�	�"O@,�-P�<�̍[d �(�r�2"O��i'E�:>F0�V��K�Za
0"O6̚%�X�?�h9������`"Ov���L�x��e�	+c�@��"OL�a�Jk��4y����_wNU�"O���`��?�
y!%m�s̝�Q"O�󵠘�z����87��|�5"Oj2I����$
�P0G�N���"OVQ!�Z 3�\�Y�)v��kvQV�<��T=i�9���[�)��t��ÆH�<��HI6+q,����$��mX5I�<��
���d���Miޔ�]E�<���@>��1��?\}���DUh�<q��C-I���a�/��S�ը@Of�<�#���"�t=`�+�1~���0s,Y^�<񄌚�V��D�ʲb�
��Cb�<I�HOU��F�΄��3lZ�<�`��(���@� ���0 �
l�<Y�.PQ2zQ�4ϒ�T����Dm�<���Skr>T�Q ��{�䭰Q�*X�:=���%���h��P'J��1�����ԡ������!��̢ �~�B���]�-�@�;a�6��R�#��2DZ��lF���$�q�d����Au�z%��[v(ً%��I`��Qk3 0ݨ���x{���/��29S @S�+	\����(\O�
d�ƖC�D�js�
�7�`uӳ��ʙ5�ni��� C1dp	��T�4���Yc�V6?��D��!��A���e����2IV5f!򄃤E���y4f&�v9j'G�$�(lt�	CjdA!��uwx�K"K�F���Y&�~�����y7�/�2T���ޓH��A)�����x�µc�t���A4❪1b��"T;F��;f�Bap�#߫$x@I`˂4`�`�[���D?��&�4�� �Pp"A�E������5<O�@@Ra��C����`T�t#�����N"Đ1��I�0�4��h�x�L���bM���PK��L�n��x�(ˢS�vh� KΏ��:�+����r��@�d��BeF$�����.F{�jFh� P��E����/u�|�F�;A��p#ui�$�xb�-@ᆙ�#ᝏD^Q k֡g�z�Y:;�̀�D�p5Z�Q�F퐽�S!�F��D�Z���;�� �Tk�=�<�b���f�C�&p���$�Q{Dp��E�@ q;���L�ݰ��D
Pv�iT�Q4$v�̲�K�}ZL�p��G��(,�z�X�1UH�=����Z����ϱWO�[E�X6\�Ƶ�2J�$[|�{��;jz�E��ת[��+re<0�@��VG�=���/�����$�	�2,y� C���,�����'��<;�Ύ�4Q�P��!.��@17������5�^18��=��h����Z��_4R^��2g/�OƖ4f����L�^Q� ��gѩcd�� ��y�����3	q�rƶl�I�E=^m���EX?�Fϻ{2�۲IE.ɒaJGɃh�ظ��<�u�6jSx���*+�#���c��5i�$E�G-�� � h��"<	�e�V��|���b�K��%���	*�戛0�֟>Jf�{ҭ�=����	,tK���'R�	\��� 
��7���v@����j�?4�*Y�`	z,�$�$޿h���;#S������B�dEb�iD;\q��|��O�<����φܘ�
p� ���K06��apaL�=eV|cc��Y��Ep�T�u8��ÆE64��~�W.^�t�A��j�4d�!�E��M�U�˚,:�����k3���,[)���"�B�[Җy�.�kD�^���`#�ؤT�XH��"�!��7�ȱ�B�m�H���A_������H��6@�V�,��!^>���)�2�fH��˦�0�f/;sDp`�n�w�fq�fe:�O�=�/R8*̦��AJ�9!�.��ꔤ���R̛8�*�k��;N�P}�Aߺ/�Q�` P)��z$�X`��=]"�/&� �� 㡀&<��H���?hr �٪���yv1;�5;�����(��Ѕ��\V��Q�
<M��yv�؁n;��{�$3c�I2�h2a
�05�\;1��3ˊ�O&d�4 ��z��5��y^U[�'>�k�kH6:�X+5l�2i�)�2�;��P�q��6T��K��ܠ��O�9p.���c�o��<]~u+#��>��}RC+���gd���o҂P�֘��i���%&���=���C`Ze��.ѥ8������d�s~��1�'C�4v`��k��<�S��ua���/����y���	Dq���;`eW]�i�0�6 X�~B�H8J�hc�G�?߰��d��ē}�y)M	'�f�s�ɐn���*���V�S&f�� 瀎>]��H��`�B�ɻl7�p���, /ԡ �㗖T:���,�$�2����B<|mi��/�S��򤀣]}J�CT�_��#�j�t�!�dɌb֝�&B�"{Ͷ�[#H����0�ݘh&�8����7�lCP�'H��0�_�Di�ō^!GG�ui	��dy�w�Qp_^x0�3g��U���sS\
�a'dq��s�L5��jVA�0}�Ƞ��4v,�  m<D��:�؏	Ĝ8����a&Z0I�D:D��rs+�$�,���,t@� 9D�� a�� B����oX�9,�!��:D�h�t\4];����5���:��;D�P 0��
tl���D��/{��ҏ8D���������){4� c3!-D�Txd΋J����u`t�q�(D��2��_��u-ѤW���9e($D�toѓo�v}�i�8b�*]C��#D��B��/� �P�G~�:-rs!D�<����(i���Y<IT��9D�l!ƪG�u��²�֎��� ֨4D���9�T�Ѱ��0غ��G�0D� B�#H$3���f���C���Bm�8�L"�O�9n����ޱ9�����F.5��\8ӬD%^dazBCW�ct&�I"ү3�bI�\*L�	l�e2���� �y���8�^d0�ɨck^Ii�O���bhV]YeϜl�ժc�%ҧCFH���\*:�p�Be��"4^��ȓ2G��R	Zj.Ț�$ɫV|� -������O��J�!GJ�g�	�_`�q��ï&d=��)͠)�B�I�1��좄��Zq��(��z[~�i�n�/O�~�� )$�N����W�'�����W:^x�,x���;nB�)Q�4P`\"��8OڝPs�N�Weތٲ�ӳJ�(j�l9n��`b��WZlm� B�$�ހ���� $�֑[��Vv؞ܨ1I��5���E�Ƒ  �����<ir,��O�``�K�D:r`Z^�
)�K� Lhw�O�6"	�sJ �Anu����� ,���Q]�<Q�JS�j��#�SyV}��i��*���,�Q�0}�a4N�~�iઓ�i����xX]�t	Wټc��$W�� ��6L����)�\���A�fF&��L��K'"�Zp��� p�w,�b�hb"M�%+���.C�z��xh��%�LT�J>1��Й�<�8��G�~�P���dRo�'ez�ː�ѕ��]*%�CL�ڙ`��|@����9���P/ǣ?����Ɩ8��$�󭞎g�p��D�*J�h��>;��!G���3"��B0gգD�{���	T.� kro*sR5�`dн5C
��`nH�oK�L �(}```���xbJT��dU[��I�h��[�&�0p�Z����6����^�of�	)�jM{��I�i����y���V� �G#� je��� �;��?a]e�H�!�j�]��ⲁ�'aV�4C��y�J�-�Ur��@�F<Z�I!��Z��0�Ba\�fY�?������ޮ`���2�L?~�AD��W�x��QB5��Y�a�"-�����/BG~�۶m�R�+#%�9,4��#�f�A��-�90Q0��)�z�	ea��!B�c�IZ#����ɷM,�Y�!�x�5ѵ�X}v�l���f�  1���0#H�P����+E�U{lB��C�)� &I��C�� �{D�E%yߚ)9�ES�K40��am�8@JBx�WM� ]8u���9��kT�E$z؊q"5�P12���/H���("hɽwy,��OT=�+P�mZ����!%xh�e��<��&�(�b���Q��Ðn]����/�" LI��qw�]>��<�Ua�b����`:O��lׄ*p��;B@�lbơ��
-�L<���#ˆ}s��۟uД�r/�&��|Cb��Dy����I�it�p�g@�	NE���CL&c>O�@	f�N�4`�EmΚ+�4C1I	�f=f���L\����BQ*#��Zх�_h̙)W��)PC�ɇcE��z�ψ�"�.�qF���Xu Ĉ�d���ARC=h��"q+dH��"v/� ��i˨�\��PZ�Y�� �
��H����:]��B䉤WF �:%�� 
X��`t��
S�t��.T��0�p%	Ay6���E�|jr@�#!�O�H[5��#i�hL��C@p�pa��'r�hYe�7S��:pF*ڊTڦ"װJar�[��O#�z0�RM�&k!`-�t��9�p<�O��f�AP(�*��逅&�k�'�:Ы�&�;\{(2�K'q5~��F�=zdlUH��E���S��8vG��X%��EH<�#�Q�c���`!H^1�������pap�M����Ë�ir���d�谈��%[�BH h�iV$ �w��8y!�Vr��BU�?�||�s"݌o�~IxG���Q_h�;�
ǵ=,��&�?��'bUN�I2$�����l�V�1%�9|����D�rϞ؃���=$� �P�Q5�x�@�E{���A0�q3@MW ��y�
�~O:�IbL,�-	ЩƆ��O��[�i��(g$|0��M28�{��?Rڬm�qL�3o�9U#�V�%��x
��B5b7�l��j	��'f���uBO�&R@�B ��r�X����	Ü0�Dhu��/_Kv����4a|!�M���r�ܙr@4�J���F`����м.�ʕm�V���ـ�,�3�I<`RT��'HO${KV��Ѭ�&
`B�I�)���O�m�t�Y�'�*S:�%���:�`t�vן$y����W�`��%���κG��CsA s!��΁��Ls4$�`��hS�Ѕ_x!�$�]U�1J�O��$	a��G��!�d 8E��@PF�\�)�B��!��	�/��D�\�I7.e�ǌ�p�!�P`�橂1jK�v"Lm��L�w�!�䛬c}2�ٲK&3>�S�J}P�"O ��0�S/X�B�����#�F<�@"O�T���["J���AbNʉ>��1��"O�s��FӜ�1 ��o�
��"O����F�JLDQÅ݈�Z�@e"O��(����
�&��/���Z�"OD]s���tP��DV�r��2F"O �U�W�C�E���B�Bj�"OF����X�K0����ǆ#��qg"O�����
4X�'G>s���kE"OL�:�j�:FT�2aA�=Z~����"O���Ł� f��PP�A�Mo�js"O�����5g��(�π>P��""O�ɻ2nS7#�Y��.ϲ]QN��"O=��/R#C�T��g4H�ɣ "Ox};P �=^�]�B��3���t"O�D��^0n�&T�`L�?��pH�"O"�{Ѣ��ax�LH����"Ob��H�Q�0�%�<N5<D;�"O^��T�;oXU!2��<!���iB"O%C����8b�U.��"Oja��O_�"��Fn�&~L`a� "O��a`��)�QM�3_�����"Op�`���L4>�	F�Wd���ї"O���)�0%��7H�(Q�ּ�"OV��@S>sO�X�v� 0��"O� ��JV*Wp(�N�a�"O4��"	�5
3���v-�iU�"O-H���-,9��xb�ұyQ���"OH�yt�V�{	���fӝ_Z~�"O
pe��U�񻐯��@���F"O�IT�d��0����s��1�V"O� &t �o� f�����I�
 ��e B"O��v���9>��A獆x��)�"O�Y���JW�l�(�!ۻ��Z#"O�ᛖ��	�
����|���"O:���kS�V�$ a,��I[�"O�PP�x����׏�Mh�L	D"Oj�#�ۦ� 2mҾ!14�PE"OLi��(-�4��b���9X#�"OF]AF�]h��#��B?�!�Q)��:A�i� �
3�N�[p!�d=i>���PJ�����ݻa�!򄛛e�(�/�Ut�aaO�q�!�d��O���U�c�Hĉ�� �!�����C�:z	���&tK!�D?�|���\GH���&F1)$!�M���H�-��-�PP��I6�!�d�l�Ą񬉏-��1ku�4󤍻��ĠB��0QX�t��T�k�ؼs�4U��6�i�B( űi��K���K:6�qRgC?0�ީp�O8J���C��'u4���ݺ��S�H|���F$��`r2�E/�,Y�C�~?I�%s��Y�"�%86�Ӻˌ�)Ұ R������ K�Z$Kq�_�dʟ���pid(��pu��riI�L��l��T5���sq�;n��n�Mܐ�N����H&!�^zD=i�v�`c!F ��6D��B.���#��SaY$ApE�X28|�:co��Vz������e构S����*t4�	о/Q,�rbA��@��y�r�֓3	�� �OQ>�`�h!*��9�p�	
�4�r�w���J����@�>�|�-O����9[�G��[,�K��>i��� �'8ԧ0|�Ri0�����ǂQ�M����,��+�A�h~�A����>�O��Zr�.��@�K������ߞOb�'�Q1Wo?�0|�bÏL�8� :x�N���C�Y?	��!����e�\�s����U
�P|�c�Ǭ/�:l����^���?�~��⊃��S�O~h���ɛ!18q� )H��"姖�:��s��S�A���q��#H�e�N��R�B��[�R�@��	 	�d�S�%W�#�~h���5�b�l��_5� �D��%r�Z<"�b�R�.T�cE���� ��Y����v�)��[�,�� +�p�ޱ��S�����Y��oZ���S�OG̹ɶ�"\Q�����˱I��d�f��l:� �e;��S����\G��bE��9�����F�`�L��e�?�$�*�a��˓�M������^,`d(�i�<L�>�'�Z��@��2y��n0���I�b�P�C��5@q��3}��ĩ��<Y� ��^��-�ʳL��?�:��ٳ"��P0T�\Ul(3�"uӒ0sFdV�*d�"��ʍe��	�M~r�����C��(��Ѳ��U�C��Y�`�N�<A��^>�(��농Ug~��ao�d�<iG
�[=j�8���eS`���d�<�v�L�f�Z�h���5�F�F��j�<	�
�5NP�f%C$_��LH7�
f�<�"ˈ&:�\����[�{2��D��x�<�����Zp���2 ���95`w�<�"�ـ#��@���e�69�ȓeX;`!
z��=�g�[@�ȓ ..�!�HܠpEM���ؐL	��I�eȶ.O�1�ICM�F��T�ȓ=vJq��#ǬgN���-����ȓV�̝Y�ϲPQ����X����ȓ$V0��'�\(7.�[���$'4��ȓ`��\����<�2g���
��ȓ,:L�Z�唈?�U�W��6��ȓ�R�i�.�;��$ʥ�L,n�}�ȓ8��`s��5Q����C�+%��ȇȓ+�v iV΃(upJ\(��.+���	�@��sM#*�����,�:������SG��`@ xZ�Д!�D�n���	I!�V�K��Q�kX!��
�vy���V��?NL�kQ	��9!�*>��y7�Û#J�E;�Q��!�� �x�v�:U�xD8!�Q�;;��{�"Oށ��ʤ-(%�� ��$F�d"OjL����H�@z�`B�s�.�6"O�4S���-Pْ"OTN�(J�"O�:~@��\X��UK�ꊐ+x!�$�9���W�^	\���#X�3f!�$>^q���uφ�K�1c��W�$w!�D�9Y1�} tJ
�x�T�^�-�!�d "yb<��&���b&͟G�!�D*g��8D��;���j��̌`�!�Dѕc�@ CP�&��D�@�!��_��,�#HF-tZr�Z@�	n4C�ɳT �P���(墀QC�]�C�	�
E^B6N�;$$� !t�	!v�C�I;x��00*W((�j�ꖯܪzB䉮!Ad��uʍ�B�@`z4�4c�C�		V7�eW��z%[Fjט^�xC�I5B����j1q^6����*LLC�	�X�
 ��4F�2�3�^S�C�,^#�4i�l6'����)�1u>C�IRm^�����'	ʍUbS)B�	�D�M1D��a�n�+�BC䉉8l^�*Q��u$����̄�P,C�	e��Ee%ԔhA����e�C�I���p)�?P�&	b�B�?]�B�ɠTҴR�^k��)A�/Ө =�C�	Ehhx��M�M����R��!o��B䉿h|`G#Na�2ѥ%��Y��B�	�Mʎ@���P?kR^���.�/ͮB�I�^|XٶnD���c�m��NC�	/�Q�[?GR��	O�k�2C�I�:�A����z}Ͱ`����C�	�W.�5��A� ��8�S�F�nC䉅ka�q+�+�\�$��4�lC䉺9Y0\�E�#�
��@��#H�B�ɨ[R�҆�56���F��ps�B䉷�2���M^�qd:T�g�C�z��C�*N�|3��L�:\ASC�%�C��_�~%����mB�C��X�fؤC䉤S����
x0���/Y�C���$���!$ɐQ`���gw�C� Y��kPJ͔pY���(��C�7.��ẅ́� ���I/nOfB�ɕB�陑o�gr=���I�"B䉎YuԜ��k�ǆs�Ș�L�RC�ɨ�~�#�!�W�P"*ռ$6C�ɰ6���Q��r6B!�2
U
	�B�I�emp-��E�!��<�,�g�C�ɾ��)UK�6��H����|�B��!!� ��$��(�TÂ�͂I��B�ɱ?�$��+K�PXX 剌�Bd�B��f�Z�B�E�,N~1S��IL<RC䉍.�i�W��4l���u JMfC�ɹC�� �ѧӱh�hT�1�H�P�NC�	�3́Q�ԙUd.�`�%�)A,C�ɽ,�е�	�9X��s΄�V!BB�I;�ӑ/�W�VT#0�WP�6B�	?[zI����|:���.+0B�/񌴹P�¥d��}�Mk��C��1 (���؋<���fʅ��C�	�|��Рc Y�	�U"'oU�i�C䉽U�h�f�էڝ����(XC�	/��!�t�քVNq��9ySvC�I�S��<���>u�����
@8 bC�)� j|"c��7�!�r+	���F"O�	�D$U O&4� lт����u"O���$�3:قB�Ȗ`A��h"O8S�H�{s2�Z`�H,Pت�"O1�G�S(c���k�V 	��"O��!�
Ў[�,�C���
r	���"OJ�[7��3p��8S�C+>���"O^\�U��$SUI ��ɺ�L��&"O�ycFIL�.��RAFN-z�"O�D���G�.4hR寋�gu�A�"O�t!��Z(�~��.Z.Q^����"O��p�� �$E ��:h$=7"O�I*�ρF�$ɓ�V�&Ͱ4"O��1@ыg�Jm�#�mm�E"O�o�T6@�Ƣ�=n�����"O����^�^�H�#�b���iG"O𥺂� xı���I�5 !��"O"�UM�_ �4:��I&�2�"O��F�_�+)��P��0Dy��"Op��e�O��X��d���vmj5�P"ON�KF�,�j��ȇ�5�^]Z�"O��������d!D	 b����3"O��a�E�B�T�"oLVO
]X"OM��bL1|C�La7'D�T�"OH8s�m��9�� e0m�\�(�"OTA�F�g� a.S	?��	0�"O�P�".EEB!��*8�έ�w"O�!I����Z��'Z�d4S�"O&�+�d�}0�)�Fڕ=��}�G"O�qz"i�/F�*�0��[�h �"O�=�S�D(=z�AԏF�nH��"O6lK�����E�&H� �L�"O���c�D�)b=Zp-F\�Rl�e"O�a��͵}�f}!���)kpX
E"O�4(��Y9C{���2
�_ԲB"O6����Ԙ!B����h	*�8�*O$s@�Q�R�=�W1�(i��'f$�:��W�p|�Sڠ8r1��'9�E���=Le���%3ȠM��'�>A��!�0f�|�i۰+�x�[�'H�	 ��[�&�p�r�dã,S(�b
�'�����E߉qe��;� +w^���	�'y<YD�>KP *A�u��R	�'��8�P�%"�q�W
�.7��aa�'�6�p��R%d�y�g��/HZ<��'־$i��|���v��"�e��'*"EZ`iߋ�� !Qo��$�E8�'�>3����@@���	ք �,�8
�'#��JR��j��?x�́0�i'D���M�+ei���.��A 0D���M͡'�{0��JhU�/D�����K/k�6Ԡ��/+Cru�b�-D�X
�A^�c���rp$O-AO��a�&8D�����D8^�lt`p� f�9��7D�X�˙� 41�`^�z�X�� �3D����0M[,4Y�cں-"����`0D��r󉌰c7���gV2	+��#D�X[gn1	��f@w���JTK7D�X*u'Z��8UD��R8��8G 6D���-M'"&�Ւ$�̟$<�h��
4D�xR1�T����c��H|��R��1D�$�0j�O���� �(��li�:D��F�h��m��"�Y�,���7D�<8��ʣ"^.k̜!~�p��I4D�� J[q��F��R@nԘo7ą��"On`#N�1+�
�D�?�`9#�"O�jRlڀF_���C/�):q"O���9C6Y��=jҽ��*O���WO�@�|�p"S������'g�4Z��<���(�ʍ�&����'U89�4X=_�	j��Z��DK�'Z`�5�� p� ��E��ʤ*	�'.1��Ə(#X���P H��>H��'G� ��G�d��T��ڨt�zB�'��M2�n��X��HNͷs�8\��'�Z�3�$Q�d���8ǁ�'zN��	�'48����$)����ցr�rp�	�'�ny��LZ�2r��e&J�^Ϥ��'� �ku$G,��@QuD�OX���'�t��䔄q`�J/ MC8��'�
P����	
�nM��/JF�$�:�''*���;xL	+6k��r�<�
�'hظ�e�YB�]��L�a�}�
�'�Prb�����#�"I@	r
�'����Y�0 �b�ٰ0��P
�'�HQ۔�� 6͈�h�/ˢ4I0:	�'�9�Fҡ`�V���(A��	�'�>���#Խ1/�&n�1%����'�@rC	��'��9���-�@�
�'�\��C� E�xT�uE�.��@
�'�}#LA"F�l�YU���^A;	�'Z(�P$ϙ(����t�
9 Aƽ�	�'�(�c���?�C$͘�`�(�y
�'(])��S�f��]�f�(�F���'t�\�V�
�I�(x��	T2%��0��'R&��e	�o�4$�<g� ��	�'.N��S.�z}�CM$a�t,`
�'����6+�ĨЂ�ʩC�q��'����o�'L��4F�H	�'q��0T%�2���1��^<!&̵��'�V�+�ɜ�[�2��']3~R�	�'IT�����t��j�{4|��'�2D*�ǚ&@��-q�!"P�9�'��͉�d�)|f��a��0�����'y`�pf�ɂ�f�`���E�Pk�'J�(�^�xD2Ɓ΂E��|J�'�^��"靨[����Fɕ@�Q��'�x8����H�t�DU8ظ���'8La��gW4g��Q$A�,∥[�'"��������q�CF u��3
�'�y�  ���     �  <     �*  �5  �>  WJ  �U  E\  �b  �h  %o  hu  �{  �  2�  v�  ��  ��  <�  ~�  ��  �  H�  ��  ��  ��  :�  ��  �  O�  ��  ��  �  a �	 e  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\����IW��~ܖ<��O%[4A7a�a4^��ȓE���g�.k��]&��\\�y�ȓb��A`���@3�}�#�S8I	�D�ȓz�Y+0NU�D�����t؄�n��DY�/�iu�xv�@�7�����c���gB�-~*9��k@�N�V��ȓ	�\�+ҽX��e2ӆ�p� ��u��Aw��e̕q��6McС�ȓ�ؔ�B!��GLaّ���*�ȓj��ɉ���S����%fS�M�Q���v��F�~~�;��q����9\O`c��]�7H�aK���}�� ��'o�'������b ��
hN�[��ޡ"<P��W:��`F�K�F�N��v��!I��D�ɦ� ���JU�q,4R�A
( PQP3��$�yB*P�-blY�ƠI �bL�1��ܦO���hO�7�:e��AP�e{��ZgI��(� ��d�>�e�0���H��Yb���� �����f�N���I�1xb�aR��0��E}_����O���,a��ܸb;��#���x;~D���?����4�0���`\@�s�"�h?����Ӓ^��1���ւ{Oj�J���K�zB�ɹ��db2iޑX2誤�X3}:(b����/� 锭��.ڱY�@�o(DB�	Ls�� �����˝N����rǄ���å"O*9�F�,���+�H^�t�
���"O0)1`�� 	�B�3� �8o�@l�"O�-J�F�8v~�騤�^�m��L�""OP��FL�&`���3��0s��b$"OLݺ��>辐y���?�Qה|��'����RmM���0�Ӧ�nt2��
��K3�"��!�pđ�m-fmf����D+�y��E��@Sc�b!@������?���' .m��c]�<����;MX�
�'�N1:��T�y�P��_�,���
�'Z�<�Є:ƶ�h�=[j�5��'�*�a��� n��J6�ع]n2!�L<�<|O>uӑ@�b�\�! H
/��E	p"O�l�䊅�>*t§I�z��P"OHА�_%L6n}[�M��^���1��'����'U��"&�+'�$�! ߏN��D9�'e�g'4�p�@)�i~萊�D�N�O�2eP�̑5)��pk݈D���h
�'�E�'ߝ.,�	���@g|ͺ�'A�e+#��8Fp����]����2�'���F�06��p��4	�ĉ�'S�����M2��Q ��KV`��Q�'1rD~�0�j��ߵ2�|��Ԍ�y���xr�}�ΐ�u�ă��3I1OR��k�@����R;Z���f��-h������Y[az����r���8�dęb;�$J��ѻI��hO�䓐	P�(�L[c�Ɔlxh��w"O�x�gL���zg�� hZ.��
�'a֘��Y�tÊT���wE\���'�X�pp*�=M�n��&mӂmP�'�����e)Z�r��d e�<���%5���'`�PiRG�^�<9�c�m��� m� Į���W�<�W�D�4�L�9��W�S.X+%f W�j���O�\�b �-f���ӀaK�8
�'k"�f�uϬ��ï�!WY@����D'<O4SߣW_�	� 
�4��1�CO���u�߈x\�X��̟�^ ͱR.7D�0&�X�[�$1�w��n��ȡe�)D���d%ɫ
pYx`)Y�y��$h�C:D�� '�Ơ��H�e�x��D7ړMy�?�w��:l��QR���*�J�Z�&4�Ig��\���^	\Ehɢ����!��i�!�dQ�s�iP3��� 1���X�\�!�ɗjݢ��P�^�|��5G�'���?!� �j!�$ ���xȱ���:�:���t@��%�I�CT�>����uX0�d��'?1"�`���
d⤆ȓx�B1�2���:�T�5�ݐ��Y���� �r#�>7^�)Q���:g>��D0���0H��ņT����`O��)��>,�p�2&��� ��%i��e�'�ў"}E�1�\�䮔4c�Z�P�%Ut�<�&�~�����n�����h��p=���O�p�(�'AX'w�<x"�g�<���R6��+$#��@
�RՠBH�<YA"U-�@)heH�AX��d�j�<��H�eW��X��Cՠ���l�<ٕ ~V��tI9c"��a��Uj�Ix���O�.�	��؉0�$��B�� �9k�'� H兄:Ք�{��1c��x
�}R̘x�h�G>�"z#'�%^Ru��/LO��`��_�lL��䕡O�����ȶ��'��{p+�3}
� 6�`�*�9�`x��hG��P���1�HO��
P�.��C��nn�yg�
!w9���'�ar�,Y���=/ҡ9�'��M����s�J4�\�.�Z��ʆR�pc�"Od2A�Z+?���@m��b"Op#E>P\��PJ�BꝊ�"OT,�r�NO���puꏭ-b��"Oh�X�͘Rq��`
�($���א|B�|���5���[�ĝ�(����1��lo�C�<�2���
�->q�2��	�OԴC䉕<��ɀU$Ȋvw�0h���6��$���~R�&����A_�$����о��'P�V�'m"WF�H�t��m�h��*54�yt�S�Fi{u��8,�W��Gd!�d�=ti����Ψ�"�����HD�'Qў�>����m����5� `��+D����jO�O��$��J�Jr��*AA(D��e·�\���K۬�.��g |O2b���3L�-�ΐ�vf�#�ȹqk(D��kW�S���xy��Z�S�i��&D����*9F�RG�l*�[n?D�T�P�ىb
�$,;X{��'>��mZ�T6(,�fZQ�! `��xB��?[n��+���w���r%e��٪���0ғS���	��]i�5�f-��8�F���
PԤ8� Ԍz�3neH]�ȓ'\䝨A��>9f(��Į�2Z�~��>1������q7��	�1�*6N��y���&<x�8f�
(�6�QЬ�!�y�����BT'�-&�u��P!�y2�?N�v����e� e
�yB�*L�8X�uq�Uڒ�\��yb� �,� 1�Xc$�,�!(���y���F�`��F��I�� �yBG� )��]90��>#� Ӑ*���y"U�Z��ab(��:Y�T
�-�y�#�:4ݨb�i -�P ���W��y�.��<�`�ɤ�ݯVB$��0'R0�yJ�-j�h��!�EH�����Y3�y����:�zh9���6@<��'mJ�y�n�	-��qH���=�DZ�C��y�Ζ�{����,� �B���K��y��X���!!3#L�҆l��cS��y���.Jr�IׯU�$;f�Z�eW�y�č�;�h\��o�;}��6��%�y���V�.-P�Дޑ��I��y���$
��`��IDnYk�R��yRc����@�p`8Jn��9���%�y�)�B�,�S�\Ċ�C-�y��G��(�E��"O�r��rO���y�e�_��qb� �Q&	b,J��y��]��t�2�de�1�Ô�yB@�2Q��U*�/�
1�|L�q�Q��yr-/4�s1��/�j� ����y���"�dx�"�I8wY�@�0��1�y���gp��q/?<Ť���I���yr �R�F`)�!Z**7$<ۂ���y��ոv
�0�]/¡��H0�y�E/fν��'�3&`Պ���y�d��1)攡6�G�A�����y�g�Y򦀲��[�p �[ �F��y򎑪;�T�Eą�mAحK�"E��y���.8|���_�{�%��_��y�ņ�'����!ޖ
�
�+'�2�y
� ��"�D�^�EC�Ga}f�a�"O���uY?�t�u�E�El4�b"O���"�!:�~���M�]����"O����<>l�R��ؑa�2�"O���m	TxR���M�L@���'�2�'��'j�'yr�'�r�'� ����p����5iE):@����'�"�'���'�"�'���'V��'�z�Y��&/� ����val�'�'���'�"�'���'[��' ��'�,)�U��y�p�9��J�:���0�'���'���'z��'���'�'�,m��$T4'� (cp�ԛYĂ��'ZB�'��'R�'���'��'*|����7}B��P���hX�5�'N�'z�'o�'.r�'��'q�m:B�$'G���'  
d�y�'���'��'_��'��'J��'�M0Pg�+MZ^ܢ�L�`(�iq��'��'���'2�'b�'
r�'2�8��H�W��)p�ȅB������'q��'�r�'~B�'A��'�2�'��kf�t)@u�Ш�3d:<���'~B�'��'��'?��'n�'p����!�w��a%�ԱS��Z�M3��?���?Q���?i��?����?A!�k�Y���]��[qc�(���$�OV���O���O���O��$�O���75&`���Aϧ ��	')�*���O���O�D�O����Odo�P�I�YUp5��*m�<Z��ӱ��I�-O��D�<�|�'��6�O�$r�4.�>��y�h� :<���c��0*�4�����'�@7��m~�`�����^`�%�1 ��l�ʟP;�$Q����' L����OI)�4����"�@��1�<��W���;�Q���Oʓ�h�\@r��~DSBC�$43�-�!���uc0�#��K��\��w��1U�G&���A���m��z`�}ӊ�l��<y�O1�����Fw�r扥X��g�ǝ6���(N<Z��
|�f<8C)�Q�$�G{�O��
�9�2���� �x�SqD"�yX��%��2�4]�-�<9�D�jR����N�>���(�h���'���
S�Ag���	w}��/⼱pT*�	G:��4)��ɣ4�:����%jc>m�˞׺���'�� � Ι~������̫wzܙjU[��'{��9O~=Y��pM�|hr�Y�9�	2 <O��lZ�3
�|���4�H���
�r�Hss$�6���	�4O �l��M���_����4����f��YrCԝ�NxA�;L�rE�@�	#$�d�<ͧ�?���?���?Y��\�'.$�aŊ�kc��r�A������}3�ӟ���џ�&?��ɶ9N���A,K�=?:E��E�X�,p�OJnZ��M�'�'!�O���Oly':v��@��'ء?����N4ў'"����		��mK$Q��
`���$���Ӟ͎4�U iv�0[&F͐Iy$8�	�i)���'��o~�|y�fC�Y�Ȑ��E �����e.�p��LK�AfT����/|>���D��*i⭣Q�����' ��eW
V�Tj���`E�����*MN�A ��AḸ�D%1'*i9���/p�=qU�GH�`� ��yw�IC��m�h��#+lډ�4��1:T�0֩ +7�s��;��BG�'TR �3�4���1 \	��@�Wp�b�(U�#8M!�ȍ�d'���JYkZ�R�D�S�䰢�Th��6�<�����$�O��d�Ot��s:OҴ��б ��( A��C�H��ئ���d����	�ؔ'G���}�B���OkL��D� �!7�)YG�	���Q+B���'��I�\�I�����|��'HI�ϰXk�q���!JT���	.k-��'zR�'/j�Ȗ�o���$�O��d�����M�~�����:q��&�æ��cy��'��&X�����4`��y�l�Iج���AߝY~Бo��Ɍ6
*d��4�?!��?y�����^ �+��Ǫ[�|ԙtN۰e����^�����e�)�I�������~�r�	�P��1��c�ڦYi&�ݿ�M/�M���?��������?���mX�0p%m�q���ۧ�% HN�9��i�F�C3�4�1O����4F������E;�;vj�/��lZ����I՟�a��'�M���?���?q�Ӻ�e�_�.��$+��!Yj̐�5�Kͦ���]yr,���yʟ��d�O���p����R%t&a����u��6�O�@w�Po��$�I���<��ɾ>/E�v4�p��ЂK����n����'���'���'��S^V�����J�h.�BB�E32�p���M#���?q��?]?�'����)i\)Q�^m;���6)]�Rl��'���'U,�Ӓ�']R�'8�Х*��7�+�88��b^�t�AR;e3F�m����Iş���T�'R	̕��d�
iZxx&�+��xsSH�
�6m�O��d�O��d�<�gA3U�����i!"�(1�F Au�@�n���>�M����d�O��d�Of��55O��d�����k�~��gj� 1Ь���r��$�ON˓\�1qP?��	̟��7K 5!�aY=�P� �+|��qc�O����OZ�$�'*��d�|Γ����[i���	��(T��`��Z��M�*O��p���!�	ԟ����?�a�O��Z�s�Xdbv��3���K�	�?1���?I�I	�<�J>)��D��%{�!� Aԣ>G�@�JØ�M�Q�a��ش�?���?��'p�'bGI�����MZ$D,l267D3:��"|��KQ�!C6*ʏ��,�Ϙ;NH���i��'F�+�4q�fO��d�O��I�rkT�r������E���'�Vij�y"�'���'jT� ���s
�*732`A� ե$EJ5���ix"���+�b���	p�i��P�"�^<	���HQ��+䎼>��~̓�?����?�*O��WGK�s�2T�I.Z���⇅��Dz$�$���	��&��'K�%��	�{� ��
S(~P�q.X���'2�'�"Q���6����$�O�#� m:�hݒ$a$�x���$�O��$!��<+�}�#;�����І	Jv��`�(��d�OJ���OD˓<4�%�����>G��zs�� -иc�'2P�,6��O��O�˓�X�>�aK�8)tJ�Uv}R��Δ�q�	ȟ��'��$�%<�I�O �Iݸy���!@���t��M3p/JQfvM&��'9��b��T?���gQ�RW����-ڪ3�,�㒋{��ʓY>���P�i���'�?���k�����24�X�4�t)����xdF7Ͳ<I�i�d���O�<����Q�W�]Q�(V>rtHq@۴"�� Bƺie��'��O ^O:�$2�2VᏉ&ԉ��f�#xҼl�&Tl"<E���'�]y'`Ǽ�H��E!�&i��X��`�t�d�O �$��p߄$�T�I��{�����A�t�R�6"����L�>i�Rt̓�?A��?A�4.��G*6lUR����Gg�L7��O�Xzu��J�����Io�i�y�q��9��%m�4B�ȵ&:v�s��<����?�����d�j:�q�)�/yv܂f�̊<(dU��g��?!I>9+O�D*���Y�0�X�hX�i��Y��%�y�1O����O��$�<ѕ/��, ��%�aC��y@�x��.��۟���k�[y��Ӏ��D��|���4���!��I����꟬�'�����"�-tn��`'%R�XE1C��V�hyo���d'�Ԗ'`�	ȏ}b�j
-аDڏz�^�q���M���?�)O8����K�Sޟ@����P��Q�yޞ�P2��[��BH<�)O�����~���*V�Љ�~��YR�Ŧ��'7�-�6�r�X�O/��O�,�h6�qB���jmDː�[��dnZ~y���O��H�K�,a@)!�o�O̕�R�i���Ol���O��d��f��>�ϝ6�Y �K,|�zQc%�U?)d����O>��	��͓R�%k����v�&W���*۴�?����?���7f�'�B�'O��N5T�)�a

qj0��9/�O(�����O��O�8#��EcFa c.�X����W�ᦱ�ɛ{�e)K<y���?�K>�1uK����˘�p�ɐb�@)���'CtHK�y�'2�'"�	.)D�k�S�<m���2��Pѩ"����'�2�|rT�@9� � ��أ�nʟpC���A�� )iXc�����L��}y�iSk��7[�J�)G�Cw�L�2�G�y0:O��+���<�cbPn}"��W$�w���8y�#�
<����OH���O�˓_U��p'���n+a �}�bN���XV� R�H6�O�O4�'�
P�>Q�M�s�����!+.�9��C��IߟX�'|̻�7�i�O �	I/�l0�-C7W���WH�Yn�[y]�ԙv ��ܴ	��`zw�]<$#�h	�LL4�mWyb�`B66^���'��>�B M:c�L3.�-��)S��ڦ��'F<db��4��'rd��`b�lLL���B�B��Uj۴"������i<�'��[>c��pKS�<�!�A�9��놩�/�M3dh�������y�'�F�xC��"n`It�1���q1�uӮ���OH�ď!V�&������,�7���#NP�?<���%K��3?��>a&RG��?����?�'�z�`�ӗ �x�F��Z����ش�?e*�kӉ'g2�'�ɧ5� @�@f6��ǧ[R� BE�X����u�1O��D�O����<	d��Bͪс���g�#�i�Y�:�a�xb�'2|rZ� 	ebD1�Kӕ)�<	���x�,�c6��Oh�$�O��/m�g>�P��K���:*�dBp��4^���I���$�Ԕ'�����2;D�Lc��ߓa5�,�a�����	ӟX�Iݟ�'x��&�I�,��튤m�|\vsH&0m�%oܟ$���'5�5x�}��;:�D����m���� ��M{��?+O� 3���]��p��3:�x0���l����v㔽��pJ<9/O0hR��~�� ��A�W �4\,D�[a �٦Ŗ'U���~���O���O���L�]s'+[X�ᒡ�;*���nryR�%�O��ȑ"���໰��&܂L�һi=!�a�uӪ���O��$�|�'Y$�)���B7=(�Y`%A=p7-C+)�����@��՟p�	"5�(	c�b�m9���
#k��I9ݴ�?����?T4M��O �D�����֫K�V���9E���E1��NF,b����ߟ���Z��A��Q�4�#�SI��5�۴�?��_�'�O<�$ ���bQʷ��U��a�!"�[]��	$P�� !/�������؟ܖ'uPE2b»/��ܰ��C�Z��;`C��$&O���O|�Oʓ ��C0(� ����E\`@┳�L�f��?1��?*O��0����|� �̻v��*H�,j&�R�/&���V[�X�Iӟ�%�\�'���"�O�����;�����*L��ђU\�P�������ly�oP-V�����m�1�:��v#���轢��u�IMy����':�< ÅИq�fx���I6��)�4�?y����$��&Ν%>��I�?� s��y�B�
d&Э���:t�����3q���'o���/��?u�� )�'M�V�l�ay�Nˌ�u۴-�������'���_8J����+[�GX�ء)�P���P�\�&�%�S�Ps���ݨ~^	Q�J�L�4�oZ�jT�Eݴ�?Y���?I��L��'���V�^&ݸ��ſ�n0�b`�>6�h7M[�;Y�"|����e� �	
\pK���R%L�6�iZ��'j��H�`O��$�Ox�I�}��urY��Z3.Ϩ �c�1$�.��l�����j��@.;n�$��/�����M��E���x��'
2�|Zc�*�s�&�B�&܃�&�3hhc�OlRv�d�O
���O|�VCX Q���m,��PWM�=]ZH�0��	�'x��'�]���	ߟ��Dؠj6�R�S�uU`Y��cƆc�c�T��֟���jy" 
�\�'T��8�ǅ�#����w!V��?i���?)O����OX��@^?�kd 94� �"�aS:"0`�!�>���?Q���Sk��a&>��@�l��1�p(��K^$����Ms���䓺�Ăh��O��a������DÐ��~�)f�i���'��I�!1��H|����Ⅱ�	�ٲ�eëx/�$�f�E�K��'��ɲ��"<��O���qD�+V�D{PR�q��!۴��۹Y���o���i�Oh�i�x~"h�*����*�� H�'mY#�MS��?IF�P�<IL>y���c��ikBǮh��܃W�R+�MKv�=��'���'���!��O�����ĒP%@�Ĝ�d�8e����Ʀ���c��'�"|���K�8[a�1b�
(��FՖCW�40�ibR�'2��WZO`�D�O��(j�"\�A:#��HP��W���4���d�SB��T�'��'�"�B��3
n��Qݩ
��� �jӬ�D�7:�'�D��؟4&��X?�P@P��Αu*Z �6�ҭ?�.�E������OZ��O�˓{�Y�K��Q�Hs��h���s�^&��'��'�'��'�H�K�Gj1Ru@�01^�+�ϕ?��Q���	�D�IFy��!%Z�?
����A�a4m3��T�@��?!���䓙?)�� P����	z,�#b �^�dEk�"�}�L;vR���I�����qyK1oEZ������J��,R���..8F�ݦ��	^��ß��	f�ID��Y���Y�O��I|�$�	�-`���'&"Y���5�I0�ħ�?����i�'��4�R}�q�Z� J�C�x��':B����|��Jj�G�rq���“�<衼il剤k��u��4;��S����S�����gz�ڠ��%^�H�J�ڎ>Z���'-ܳB���|��I��5���B�7_�E���̙8(���	��F6�O����O�iH�	ܟ��t�3Q\1�*͇h������(�M��%��<�H>E�D�'��G
X�&�9Ć��xE��"a�~���O��$\�=v�)$���	��$��|&�p�q�6r�Ҙ3�k\:`���oV�m�a�O|z��?��-�к$IĶaI�ݨW3��X2ĸi�r�&�O,���O:�Ok��-^��*'% �BX�Eh�A���-pb��	ly��'���'���#XbIq�h�1�G�>� ���$1>v�$�T�I���&�P�	���S`�J1
�$�ό�w�t "2I�O5���By��'2��'
�	U�8�O�y7R�g@@���@���XQ�O��$�O,�O���OH���4Oʼ�g��@7�֋t����f�Z}��'�r�'~�6��uaI|�Fg	!NV���O��i^p!�!>%����'M�'K��'�:���'��YNP��1�4h�V�;7�ru�	m矖񦩔'(X%�5�i�O8�	W�R��PSC��.c��D˳��K��|&���Iʟ��4d�ҟ�%��)�`T;���p����v�G3��;I���jŐYl~)L|�>��')7�T!	��Fz��#�Vw�<)�m�Ԫ��4�ڂAs�Cb!�5'Ԝ�h@��(EC�}���>*:ӂOL���]���߈U[�=�"�;;��dЀE��ժ5ݯ&4f��0�L$3,�J�U�l���ʂ��.���@�2�6�k�إ26<±�K*/�)��gE�.=^�[$D56�ĴZ���az���DJ'r�u3��(�?)��?��9����O�����@��Y^�`���hǼE����Q� `�6oA�0=���ĐM���9��L�D�r�iQj?a_X1a�BζAײ��$P4 ��@�2^��2/�l��D�Լ���O��ԟ�Ɵ0�'�b��7E�/�B`"r���H��k	�'IrA+�E��p����^�;w���`�(ғ��ɩ<ц�ɜ+���M-?���C�/Vă�E>z���'��'=�]���'7��`"�e�H�nq񡭖�{��U+���{��Q�R� �p>��'SSl͂�l��,��x�͊6uo&iJ&*U-6R����T��k��9!�g�Ȏ�C�!������+�S�I����IV�S�� � ����Im�fF��^sp9�"O^��G�e�lycF�hV��V?OΌ�'x�I%pC&$�4�?����	��\�~A�і0Y�� �%��l��m�O ���O0S3JA{���)͝� 

U�ㅯ|¡Oݩ"`���'�'Fx����h�'����I�@���!J/�)�.��Ȑ%�O����b#'�Q��`���$䦩�	�x�OU��I�/߽y	�y�CA	��m(E�'�"�'32����퉑kUl<J�K>AԹ�smSZ6��$B`�	6S�!(!-��B�����h�O�0�4,
���4�?����IK>p�|���Op�d��~���*0�޲\����R�֑J�ƙ�DM�%)R
��WL&?�O�1���R@h�b�՝6
�Y�3l�67� 0Qv�҄��З�"~��5V��# ^N�}�.�8$9]s�NI⟄�ܴG��6�'�?�$�?rn@�w�KY�V<2�&�,p~�d�O�����Ty�$�PEW86@���C%���X���%�~��mN�zu��t���G�D|�'}"1�ѡ	��'��'�v�]ǟ �I����U� Q�h��>U���I9`�h����F6�Ǔm�rT	E��e $A%��t�p{ŏK�j��ؠ@[b/��BT,q�`�i��_V Q�UĆ�vX��2)o�lX�� 4$��	Ɵ&���Iş��'F����	�(�{T�C�"A��'�ʉrwG�y)��r�W4	@ɲfD#���I�<����1P�fb�44��Eoڑigh\{�(��Z�d�O����O�(X�+�O\�b>��/�� �����;�Hy�Ī�+4� QB�H-R�ҽ�@�Чw���G2�G$тeK6�N)p���A  �}�d�i�c�J��0����C���JV�_H��
w��oܓ%�~)�	
�MSq͉�~�1���Mq�ʗ*KՉ'."�'��O���D�q���Ӡ �܈��:��C�	{���/>p��XR��.B���	��M�����ז( �p�'�_>q���J;�`XȰP\@�"�� A���i�7m�OP]��M����<�OX=Ђ/��t�(!�S na���\>j*�#�7\^��h�g��`%��Pc�'k5���?9���?�)�J�Qe���;J�����nʴ���O��"~ΓM^�8��Mt�����Ct^X��I��'����GI	]�t��ӥ��j��Γc ����is��'�ӗ TL���럸�ɀN���U�mJD;����7�BM�ֆ��q���@��u��PA�S����'!u�r���n�)��R�I0P�B�RP4K���5K�F��ߟ"~�Ɉ$!��vDX#�  rWL�<$f�@B���D�	П���J��?d�ޤU�d�ۂCY#K�nP��σ�<�����>�6hQ�V�&Ld)�:9�{��^X��?�A���?u����>�ۑ�,5��u�ǥ�;C2���fs�PP �F��;���3#�؉�ȓ/�D�x�h��c1���#�)��Er� F�4YxD�RS��r	<Ą�}��a�`�\L�(�jQ������� �"�J�!�]��Ta���ȓs���E@�%S�R�i�@T��4��ȓ��`�GU ��C��(}:Ćȓ;)b�I�E<I*�Q	���v����S��������/��I�!K�5�"Q�ȓA�0�)�Հ[!5q�+A��8�ȓ
��1¢m˜QJ����_�n�j�ȓ7�l��@� q���Ů��>,�$��.�xFQ"A3�i1�
N�|�~��ȓ{��M��ȋ)>�X�K"�L�\��ȓP>��G�)Ct���GB͈ae�=�ȓ:�hy��ϲ'D1{�����U��q7L/~��	Ŵcȇ�>��9a��yd�"5O �W���ȓp&�@ C�t�D5��	�ox����B�Y.@�ze؄lK�>N����h �A�m�(���¢��Dm�ȓF�8U@&P�'oD	��Ɉ�t���f�`����Wn�p逤͂qhr��ȓ|B:���H�<����R.¾�����r�`��/��` 4e<E��ȓ{��9���+�+�*��V'��ȓz��hqCđ4r�t���_�	��S�? P :e1~������p4��"Oe�D.����QB�\��ˣ"O��B�#<u��j1mBb���ۓ"OРi�(��VL	r��}�48�V"O��R���)oT��f$�=,�D��R[��S�
��0v��%��|�w#Ƈ��G�
�F��QrG_X�h+��~~n����x�(�r�Z���g�B�n4�',�rNa���s�H�r$�ڡ�>��Z��O
>��
J6p�^�8��
�񟸑Q���!��9f�̔(�$�э9u����۸#��MD�$��b?O��i�� *V��G ��9��x�i	�vyl ��j�9� 6mC1�>�?�Ӻ�%@ҿ?kB��R��^�!'�?�$���.�~(���?�p<�1*�DY�v��>=�|if'�X�@��+����׋޷&��q�M���N���w`E��Ģn�,���F$n�-�$�'���4_�Z��i� � Qf�)�b4P��%��BрFA��({�ĕ�A��9p-@<6Zm��Ý��O�hB��$�5`��w�<���j�#�8}Ӏ��a��,�ט�2�s݁��O8~KL��u�
����Th�V���P.��������&��Y0����aZv����z�MG�E#� Z��%���8�����Z6��e`�ӧ�I�;7^�W�I{i<Q��i�$,�w�:�5��΃1u�����F�pb����Ş��"�l�^�z#^
Yk�`�R�9?E��'��\#Al��T(�B��o��\s��n�R"�\7E^�ܻ�b��+��i�]ԤT�� m���8��0�y�MB @�d�R���'��h�Q��1}���eG:x��.��~�Ip�c��R��4&�D����'%k �S�T�d1T�_i���qP�ɠ&0��J�HL�G��c���<�.x �U��'=��"4��=����=��`�I>9p@�6~r ��ա&�n�6C�l��)G ph\h��^O��x�L���ԧħ	p����- �{1�>�I���99���V	@�W�.�A��Dr��SG�:!��A��Z���X7�G.Uh@ᑆ�=t�8�Mӆ�%?��<t��#c���m�ؖ)q
���9DzZwF� ��/�c��,Q"�.�ޔ1'ӹ! ���EL�yHA�u-�2�����v]!&�2�`]	���g����=��ɺՂ�=
�<U���>��FƍV��P�
Hz	�V珢?c�֎�jc�t���H=A���3HN1z7|\Ԉ� ���um;�W��7@^:�|]Ѐ�(@0�'����-v	�@#�%��~|P���
1{�� �6�M3��j3�y`�+�-:,5�~�F�3l�J���. ��d�
��=�R&����� C__*������Ͽ��N��0��fU(x̊eJ�>ilD��1.֥���%?���x���Y�"�@�; �)�0K��]�n�C���� �H�@��(�4C���y�ŝ��b���`W9BH��1f
�X�6�\p;��)E)cpFb���		#�FM�U�;Q��ub��R-�e�&�2v �i�BP�h3#%�a����D7Bw:�[S��O�6��h�D�FV+VTB�Cw�THdeJ�y.�,Gk1O��t9ZWY<O���P%��in�(O��P�٪K�I���9je�	�!�].5n�����������;�^�S���+���?嬻e2��7��
m�x��X,�Q.ӛ;�\��r!P�����)Т�(O���_�t��ơ{f��k�
Sre��9N\*ѱeR���Ӻ�L~�'c���f�?*����]�0��X2. �Q��i�j�����M�p���Z�w?�)�@#іWH`���=�DA����>�@��MS�{B�' ��#��_�H"ՄLE�1r�R��P����Ay����
�yxG)^6�H4#��P�1���:K�N�%$K)�V
�*R�!��@�O�P��Xhsb�a�JxZ��`�E�'��B��c�ܴ����(L�,M����T1�!:�󤻟�க&��s��#4���$&�"gbͲ�e��y�6���d�� gjݒ���(OklR����YrK��l[�h��A�a��Ŀ�l��e�#F]剟��9O�S�4 XѲF�/:�M#���_,�U���:qо�2�L:�~��[c� ��_+=�fEs�����yř!��ı�(�S��h׫I��(����k���d4ň�.[�p�XH���XM�',XJ��i1�WUIbER�%PX?A��O$@�5@_!>/�xSa�L$���ķ��{�'�0����2Px�S�i����s��,��h�!C!"&��P���K��|�T@��	":T��킣�`hϓ�~ҙx2E�F�:|J�Ϛv{�b� DӴQh`�ӇDy�}B�L dJ�kC)>�z��E���E�H���G{����wS�8����KK�8Bd�-lW�9
�X�-qb4'1.�3�/6+u`@�)��j��AH������1�'k�`A�!��*��@J���O*eAD�xXB���:�Z��r鉵�!�*$�,6��WOZ���^�ADm��()�#�7B>����O�E�t@>A���5m��T��!�2퉳0��-�`��0$Ȍ]j�cп&��6-��e�|��Q?i�B���Mϧ!țv�ծ��+Dx-8�� 9ńQ;P��b�t�@��ǢS=����.@�lG-�)g@MZ�KN� �*�Lh:bҢ��@ 6���y*�9�F͘�l)�q�,�l�r�'�l8چ�B؟�)CBH;�
�q�ܡT�&�u�^�r���Qԥ >Gl�H1e���?�q�n��k�)�%_�XX����(h�q"��,ғt��4��"�g�? ��a��Q�}��!Ie��0B�z����O���aY
'��Ӌާ,O�1S��ɗ�5�i.����V0=��6L�|0l��{���q�� P6��Q�[&0���:E���5����;)Ϫ`�մiǠ	�j�^x����ꌏ�fY1hX%>�jYJ�>1�J�C*�R�ژ"Z�sq�W�<�s�ʧ9/�����H�b�*�����Id�`�;0�'���3�� �%4IKq%�3z^���}�Ϝ�o�AD�ti�fP�	'�بR(؂�HO=�0��,�y���?�lU+4O�[�D�$H)���@�8]����F��扴B|�����<ap[�O$�=y���0�ؤ
�#��C�l����צu���ar �7��p��,���
�+�v�	 �r�1RJ^�C?vT��C]_��oZ�s�Jȩt�'�Т�O�v��I� B�S��c2�jz���N���IJ�y�nءT8�%�i�E|ay�
�*�>���F�9��Л�ɉ�� �
hZɕ��O �̓w� (�'����Ұ��\�t�'�|pI�h
)�h�E'&AÜᓌ����[��H��C�z0��Oұ��ԃT��5����>�i��迟�x�Q�V����G��XP�V�1ړA���ȣ��1��R�(S�(�]m�7Z���;�
@� *dhM��kX��q�'��H��nʞ��S��_�n�����dߞY��'+t,[D��s�l9q7L�>���Jג$x��[����C��y�,5Q��,�@�ϝe9 lB\��>ـ�t����"�^�y�$��C��V\�b���$��O,�I�9$��S�WV]�f�ѱdz��D�'W@�zЩ��6���ci�Rt�����郋F B<��H\;�b���t�֝!8l,A���vh�U��(D>�	do(�)�HӎZ^F ��� �@���=`@�4K�\#@b�r>��QVc��)�b!΢+�H�yGƗ{Jjm� Ȱ�\Gx��Ʉ0��i�̕z=&2�M�'M-�M*kJ�voa}Rb�|�mk.�+pJ��3��5L!��V?���T?Y��'Q�}B��!u<rm �Թg�r�+�jx���K�3O*�S Z��މ�qf�>Lf�����7D]ʰQ5�hy��O��)b��[��UT���9oD�:G���L@H5�nփn�x�Rа�ēG]�|�f��!	�А�&@��~��\�@���RM�X|$� *�	'%��?}"�)g���	ۿi��UI��7�D]�76~M�g�vr��:�h
�<Դxg��$�6b���8P��gm$��o`�c�ɫ(@��ō� 5��lڻ!�1{H4a7����I�/�kLj�eJ��FY�C@�[%%��'���KEy�!)��O�H�嫒�N��d�a��'w��GÞ�>���]S�����T�nN(�v�zD�S<�Pz@e"� ��!���䱟 �=�'b
 ��)�G�>��gH�$=��Dc�2F�戓�A�>�t�EZ�0 3O�N���1�f���T�>�f�P�M���t�B;nߢ$�!`Fܓ�?�R�j�e���p�-Yoy�,�6Vz�ٹt�I8Fo�=)e-ք O�ma�O����)�S���i��� ń�hلx��F�7Gʹ�*«Z,̈���E��	�tyq�DK�b<Q���w�a�Ņ�/l[е�&�L>:󔀡��D�<����+z�HQ��,nB��lλA6��#��'��?�JU��.¤�dޛ��n�$)��ȓ	ƻW��1ia��P��M�'oў��V�\�b�$iS������
��l#ts�@B%R�@R�l�S�ԙy � 
QMH��WD5�����fK)3��(�C�=e��Dy�	�,G���n[	s4�)�G�����E�h�z�mV���)c�2�0Y��V�W[f4��	�<tx�B/*N����X��Go�lt�0��_n�\y�Ԉn����Whxx �.xJz�A�ЍvV�C�I�6��X�$!v1���Ř��N�_���Fy��Ͳ`�z،x�G�~�Q�eɕ^��)�� ����6$=��r�'�>(�'eXj5,�8�"W5�x ��D|¹����XydJ�R��L
㪞�r�ΰʑL��O�\[�熩e���աXn>�,� 9�	צ-� (ɕu�n�X�.��d��k9?��熞"e����ň'��P���{�n�+V�ɨ|P�z�d$���٧˧$�f}:'�B���1d&A�=j�}H&dƇ3�[ ���)I t1A�G�&Oh���#-Yd�F���O���o�yN��q���!��A0�'��8���Q?/H�и#w~�c�䅙6�|<*3CT6,l 21  ��cܓr�Dd���S��a��-4�ݛ&ڹ�~�2 ��f�6�O~��6Ј&"6�@w(͝)r��ɥ�$�1T��le��>l��0�	�T+@b���4���@A���&&X�AU�6��=Dv��B�M�Q<&�i �I�Qz<�A`�_D]�8�k�Ƹ'����ˊ?T���3��n����O�9���Gm�C�����O8��X��⃥�z�4��P����O`h2���I�
�T�x��/��Y�E�������+_ƾ��c��6�%����`�<�
cnj��f�]�H��J�H!��T�D��������bG�IX3 �`�(�PX0�%*�
b��'0`5IPDTD0il�Q���*�C'K�E	%���p��M��e�"�4q���N��(
s�ˤ�&�~&�� �(�gS ֮(`�%&�3O�p�6�d�"v݂�a6��ps���iݭ��l�Ut��@���QI�!��*yOf�SAOZ)t��9�LBX��Zā_ m:̥�a��O�NY��Ǻ��Т�L
]�X���儕��)�)Ư�yw��pؒdKR쏒>wP��E+
(ް>��F4<���� }:PMZͺ)R�DO�x(O�tQ� ��q0���#�Is���,8�nU�G��?/ў b�@U#$R$G�D�\={�������Hk^@k�S�%$�Ա�y�C������%��T��(��bH	�2��[�"O�51t�@�]�QJ�ѯE%4-�S"O��m�*Ӆu�"�rfn�
�!�dO�t:\LR��z�
P��D��!�$ۚ}���`H��Vr�m�5��!���C<&9���՞�Д"�ӷ�!�DIR�@��#�Nv�R$�	;�!��
-1�L�3@�2o^��3�ǚ/7!�d��5�%���[%� �Y��W�!�� t:�):��N���2�+�!�D��d���G�$-��a����s�!�D�r����$o��
x�4Ӕ�_"�!�d1H�<p���]�<8{��D3�!��Z�NI�<��tj�ͪo��!�I�Op��З�ϥ1��)0r���!�DB?bm�H�g��	P��Uu!���Y�Yb ��M���3"Ôl!�ě `Z����bRs���+0�ېQ!�'xT�����?
{<l�⠙:[�!��tW4L�v�Z �s�4d!��.A�A�O&l�
��3�"�!�S�t�0�rR�BB��UAb.,Z�!�	/]�Z\��e'9���"���!�D_�FjI�ES�G}6!ӕ́i�!�d%|Nr�c�!@����%�
c�!�+fr}��)��Y]j���OJap!�d��q�H�BoE!E�M��/��{!�$�-#d�)�+ɑuP|!��ވ[!򤗥
1ufě�Q�� ӑ9�!��Ͳ�$���U�+���JW%�1(�!�d��
خD�V��I=K�D��7�!򤒱[:d�`�,6KӞ�bTD�=a!��h�;�Ā4~��@��b�&|O!�[
�(3Gc�;�`� eBB�D�!��Z��P'�L�c�@!p�O�Gt!�;pκ���: /Z�CB`C�6e!���6
��A{���O-�Q#�J� 0!���Z��#Ҋ`�(a�(�L!�D�
���z'̈́�t�p��d!�=V�@�+ã�
<i�%@9
!���Y-�!:T"
+S(��b��?�!��}���5߄F�2-�eO7�!��T0B	hmi��d�ڟ]�!�Ď.<��	#�lӒ
� ��qg�49�!��E2`�ѺB�3�ƨc���9�!��Z��iJG��7/�4����Ԗk�!�ğ/B��)1�X��@����!�G(6�j=)�D���m�Hp�!�$܈S�VHaD���:p !�Os�!򄎏j
�<PS�J�w����]s�!��][�X	� �I�C��ly��V��!򤋅AM00B�c�4<���Ƥ¹�!��&#v�Ъ�P����8v'%�!���lN\�Z䥂�9��5�wbW*!�!�� �Ođ�jI]�ؘiAP%'�!�䖙w�@M[`�İ/�rc�%D+X�!��Z����
F�W|DXiE�Ts�!�� Le0�F�!�a�%��Y�""O
�Qb��W�t�J��\�D�"O6�a�S�	LX��(��@�R�r"O����e5:Ĳ�M׈D��B4"O�<'OӒ"ut$��K&�����"Oԡx��"N���Z�<�R�K!"O2�� �iZ}y0�2!ix1��"O2�#N�Q���էT1z�ճ�"O�%�c�#��$��F،���"O� �Bo�$����eBQ��9� "OZY�FD����p�Cٲ`��展"OX�Yc��K����0��%�.iX�"OD��&HC������Qt�H@3"O��Y@ހ}H�j5��9`��"O��yt H��BW�DUj���"ObP(6��$�A�%'Ѐ>e��4"O�ă0��(ظq)D�@"#F"��G"O�|�s�bm��4e_`�Aq�"O�����@oT(J1EC�c	) !��]�U�|�1��#> �#B�Z�!�$��c��L����@b��j��?�!�D �0)�DaJ}�5��!�DC/{��m��&L6AFL�]<@�!�$/HƠ��
�%K��R��Q��!�d<iFDj�&�#@�&��s�J�N�!�ē�:R�� :c�`�����G!�dN�WO��Ab�6T���rBO�%7!�dO�4�8PH/�6���M�U!�D؉}���:���m`PU��9T�!�O�E}��32i�u�0DMn�!�$ߋ���c(G�t�`��%��!��� r�Ag�,O�$d�a<?��O��=��.0#�*�R��4� ]&��H�"OTH���>����>N~R��$"O�P2G(��J~p�k0�_@e�a�"O�-��a��5�L;�@7=���"O(��&%�� C�
�HU�b �C��:�S�Ӫ�H�9��{�
�1f!>v4�B�ɢ\�>D
F�	sa��E�=s�B�Ɉm�1�c�vZ�);�lD��C�I�NȈ���N�H܀9XC�÷n+DB�I�S&�丢�
�U�V�ũ'i����>�I�Z�,�"�H��v@V2�<B� �PT��K(��q91�442HC��3��XY�D��Jц1�!E��0.�B�B��вb��+c��06/0��B�	�[3 Cm�Sg `�CLsG�B�	�q�6����cǬ2n\5o5�B�	�8���s%�2A��e���q��C�I9V&Y˒�O�.T�0��ڶu�C�I:m���G�b�0���D��C��<q@��X$����#��7H�C�ɧ�1�c��~�es���-˶B�	(O��,�D�_��E{!�B�"вB�ɝk��21ɜW��˒�n2�B䉿ɼ�Q K\>{������MutB�	���k�#wni1�@�2B�(h[P$A'&' ���f_�,CTC�ɏW�Ψ��_f����@Ȃ:fLC�ɘ@Y��u��	�������8p(C䉇d�Zc�K�5����#�ߕ~0C䉻H""<�3f�3~X�u��d%?�FC䉜Զ�	LQ	
tI���V'Y-ZB��ßQ�,A6HSf@
|��`%D�� �RV�8U��q/T��L8"O�=�V�5[����,�&f����7"Ot����:��ɠ	]�h���Q�"O�+d��2�"l*2jM!)�}$"O҄��"f&H0�R��$�,���"O�`���@�g�u��*�m���c1"O���+�5���j�^Z�i�"O8E��T�b>�� '�F"XZ:4"O^A�S �"m[ĬX��N1UMp��""O�R�co��X�ܮZ�½�"Op��d�� v�=��S�S�T�E"OXP���F�G�1#ҡ!��"O��8�ǈ6L�������J,�QQ"O�S�b�FE�����o�1Q"O�y+WMߚ}�4�"��9P�n�S�"O\��Rh�&V.��.Ԣ(��9��"O���"����p���E���x�"O�ͱ.�-\�M+��H1j����S"O|�����4��Y����nM"�"O.�6��R���їb��s�M��"O����# �P��Da�7��y�"O�\�凄�I.Q��D�h�hT#C"O�T��Đ_[�����W�)���"O`�s�7I�������R�*�Ѷ"O�!���6 ��{bK4-�����"O�J�/t0��AJ�$����"O6lSH��f�~�pG��M�V�b��'vqO&]�f��	x��Hyd&2�-I�"O��W��8j�5s��(���'"O��Dڛ*) ���������"O&���ƃ$���3�I
� eI�"O$����кpx)��j*3�2���"O*�Jf+�v�	Q���>�v,��"Ov2e͌�pl���%����#�"O4�C�-��z�%��	�[)�"O�\[���.^��;D��:a0f"O�]��ȖF�fњ�cܵXqt|��"O�}(��B�f!Sf"�R؉2��O�=E�T��G��!4�����K2(ľ�y�_'U��ə5jД	C(�(�G��yBGo�Τ����-c1���y�/N�7u�i������G�1�yR��/&*���0n�j(dC��y��Ox�XsU�Öm�v|��IA��ybk9s��)T�=�`=je��*�y�lZ�E50�1�5T��S��G��y"+Ȕ$�*�Q��3뀔�3��yBY��������0�½�c&��0>aM>�1�U(@Ǭ�ڦ�ܒLDxҡ�{�<��,	��1k@d׎oΐH�0.�_�<���Сs� 	��s/�3o!�DJ�14�������&.�&�ԆēOp<j7'��X���G>i�DU�ȓ$�Ȩw���$��l�d�;X�Rцȓ,0�R�M++���"�`�"ц�8���:Š��)
6�fn���݄�O"��u!Z�g_�y)��Bv��9��&/$0�M��5:֤2߰!gX��'�:�#b��(k��$��@�|�P�'���Y���V�Ĕ �l¤E&��'R�h��Q����z�ݑ�'�@(��A������+G��ʈ�'o��M�7`��h,��}z���' >���i�Q6��n�,U�� ��� j5)u�E�brEs�.&MZk"O
PpF�ͅ	>��&�,>����q"O�5�N߈\�TIg��~����"O&����׈];4�"Ir�97"O��Ѕ�Q2R ��zD�q/�<H#"OPT)�J�h�r�W._/h 8d"O���C-׵.;j���B�c,��*�"O�1�d�0�n(�F�M51*K��yb�/�>�"�O�|����#�yB˄ a�rX9#���p�a� ��y���<S�,,2{�b�hA�y��x��K�"�s��(��N��y���0¸k�-�u����6-��yRn�K���Ч�̑>e��SF� �y"��L(���JĐ<~X0#�M��yb/�(��10˟34�"�8Dk�/�y�hf����W�Ղ,y�2�X�y�#%�8����ۂ���y���m��tʁh��^��h*�f���y�*��s�J��b� &^`+�'���+�l�2�T<J!1�P��'���rī�;Z�4�$�&w����'�$��@�-P~h!�
j��'R �B&���I!!J9}����'_��J�T�n	a�b��|�2���'��8 ���;�X�c����m�Z�'x`�ȥQ������ >4��'�R��cI�9��Z�C^# ���'�.�2L�y�(Hȃ�$',�/D�0�Č7����oL�z�z<i�F-D�h	�*_�{�n�z5eI�{<Ta�,D��;�M�kО�c�'|�2(z�'*D��� gէM�R�M��d�ѷ�&D�����Χ�dDS �a�,��#D��(6GZ8w������D����"D�D&�/������X�j/*#W�<D�X��ꔲA6!K�N	^�t�v':D�0���Ϛ�*��u��;ZL�+cB9D��R'�Lj�(��#*Y�a�MK`�,D�<��.�,�82ּ�J���,.D��C��	N�\�K�K�jl.��p#(D���s��UE��@�bӂ�\9y��$D��b�lT�J���c�đ�c���Y�e!D�\s(�*h��Q��k\� z���� D�����`��G��+�0�+�?D��X�L�"���$F'��TN?D�|���w��y�v��x)�@#1D��h���' � �����yMX��(!D�X@(�N��8i�%9Xs/2D���f�ӋB+���A�jc9����b�<��h�QQ*dÖ&8L��d��g�<	f���r";V1�v(�f�<!���~���厞;�e�e��`�<���7;�H,1�A��+���7�[Z�<9��I�/�1��Aa���U�<��V��q�V�pYH��a!O�<�mC!�T��-ߠ:� ؄�J�<��!	�<M�-+�+ϖS��[R��G�<)gO?	�$�f��O�t��F�<�¦R<>A�-�ef�����wˍ@�<�t� hQxe�y4�����}�<i�g�D-	��S�%�P��&D_{�<�$��	�`���&^m��:F��P�<1���/�ꌒ3�U�`��<K��L�<� dm+���)�Z�#�F��f!�"O1�D";AC� �vDH�h�b5"O��y���T�b�B�_Y|�1"OD�C�����%!��>nx��g"OT���S8�t��#�gjhq�w"O8M��L�gW�l�BB^�RS"O�*s��y��� ����$"O��"���h\�<#GoH�i��"O�ݳ@��	@�t�IE��E��� �"O��#��|�VT�`��C���kW"O���T J�i�Ţ�3'��b�"O�m�GO�n�2 ��.M�@���"Otl*̛dF6Q�E͚>��y�7"Od�y1�\�H�0I�g�@�)ں���"O��[����9�� X)�><Cd��S�<a҇�_��a6�M�(%��S�<�bg��"�-�Íjb<�d�Bj�<q��+���JR��'��z��k�<1 똤i/:�i��U�|L����Dc�<9Q`�W}���J��5G�`�<���T(�V�:c,� �DC�<��ңg:0ʐn�;_
}j A�{�<F�Y��F�����7_@�$�6Xa�<a#�@p�!r��,�TYZC"@`�<�T��#x�Tq��L��Y��^g�<Q'�[�S���Af%��g~v�	&�Z�<�v�Fz&vu����|,�$(DU�<�@h�X�<)��fԲ^�@	Hq��J�<��Nۍ6��k��G����dcn�<��5�>�z��G&u��І�l�<pQ�`o�yc-¥a{8p���f�<ɗʍ#O�dɋ6�D�;�F���{�<a�j�S
X��"U'x��LS�<�3-�D�xp����#�1s!iLD�<iW���1Z��z�ӎd~�zv�WC�<��N7nJNQ��[�r|
��|�<Ѵ��>f����$D_�!�F�v�<�Sj��(���,H���Whև>�!�$^2��5iB�'��Z�H,Q5!��7i�2���+:>hm�S�{.!���0I��eX�aW���ޚ_!�1��R�ӳS�ePa@�+�!�d��7�0gi�"C@(��SQ�!�$��0ֈХ��訢1��]�!�Δ0Ѵ���������ߛB�!�č��n�!��O�R:�IІ>y!��A���0��ɔVK��BġβU~!�_�]OmzS�^�)M�}�G�̩'!�˒$�����h
X�-�)!�$Ã���*0�9M� �FjR=U!�$Tm��*ċV7 1Z����rH!�$�=�9̗6,�U*�!Q!�Dż$����4 ��x�yvjW�a�!�DP8)� r&� ,� ���!��9��E�b�]�_���b��~K!��? B<1F!R:7�����J��E�!�$�Y�H���"u�|hZTHT�N�!�R>F��2n�&i����G	�~z!�$@�x� f\�u�D��K� �!�D�!K��,�%K�!c~	{'dՈO�!���56�Q�ad��3���rPS��!��%Sr�sd�[;g��p��Mw�!�d\�qL��R���d�f�Z%/A5)t!��
�F�1��"�I���NW!�� ���CVf`�p)� ኑ��"O���7��8��m�(E&+���ya"O�\i'F�iG<�9���pJQ�@"O�i⥄� ;ɺe w(Exd�-�"O�y�Td��T_���1G�8>z�¡"O"Trf(T�R�4��veT�^X2���"Ore���5M�zy�P�U�co�yY�"Op z��=f&�#��hWX���"O�p+DU�:bC#S0Qg"O�x��^>v���C�9C:���"O���E%SNv䱓���B��9F�!�$ǬN&�X���|�F����4v!�BY2u�@�u���p� F!��4} �)���㊙j���1e>!�$��!����C�(�Y��49!��&{`Id!Αd#*�h`m�&I'!�Jn�ʤ�����B�]b6�>!�D)v9b��q���`��͛F�*�!��,V`�P3�3i���kH"s�!�4M�vl�4! ���ȵ��F�!�ɥ\����R쁏t��7�H�G�!��(��a�m�8;DN.q�!�ěO0�b"@O(m�0�'#	�8!�P���d��jlk�('�өs!�]�ذq��P]LT�92�ōO]!���*RYȸ�`7A��Pɀ��E!�:T��UGȰy����P/�%(!�$��gZ�W[�������+3!�dJ}�$�B���:�>��5IO�n!!��J����'d�2~�`]c�&U�J!�d=C܅
���>,��@� �H	!�̈Y*�P�2�6�d��/��{�!�ޤ�b=��h_@����%���!�D�A����n�!Q�t��$���y�!��]F��X�3�Xky(Q%Q�!��0YZ�9I�oQ@0���<N!�O3�z��,?|%����Z7!��;_
R�)F�%�Aqc�9-!�DU����c$F6g�
��#E!�SZ��Y����x�֩�0�Y?}	!��m�(%�� ����� �3�!��Xf<)�@�ڗ5��]�5Oو5�!�D;���A.no|�xҨJ&�Py"���]8Y�/T?4Y0�3+��yb�X�#��]���O�3{�Y��Ŗ*�y�ܐo�Xԭʃ2���"R���yr�K3
\!IY��e���l����'����FB<�t���e57���'��xS Y�u��IAa��x�I	�'���r�m��V���"����u�TJ�'��cG&��QT6���`�p���'J��ś�}��HT'N�TxZ%��'�f}���j�E � h�"OnV��<P����DQ�+2k�O�!�/+̰�dDT����1˜&{!�$�&e���@�E4fݎ "U�P�4�!��&��2bR`�^�����?�!���Ra �M�.u�Ȥꒊ�3r�!�DB1jQ������oR�Cp��1R�!�O� � Q����!�8@�A+E�!�d�ٜ2Gaz��� CY�${!�Թ;�p�`" �$��H���ۖW!����O"���dDD�R,��[�9�!��*3��z���3���a#㔔?�!�� �|�L�F�2�c�h�K+�9:t"O8ub��Tg)�1�J4z�"O����b u�,Z��;-, 䪃"O����M��!^HH�f�S�^z��u"O: 2F똋Z�l�h�i!_�B�"�"O���6NQ�,P:�a�'$Z��0`"ONq�e.ң�Bͣ�a��*(��"O�
ecC	V��.Iݖ�"o��yB㜘n1Ȉ"�)�^�8}��Л�y��0G�Y�6J޷]Z�,��yɏ/@*,���K�Uf@U�Ư���y�G�e*<�H��Q�J:���2,]8�y����l����G�����F��y2�*|p*�n�*:�� s'�4�y\�N��9�䈗�:��%�&�yROг{��5Y���? &�;�BT%�yb��W�tL��k��Ze�􋅏�y���-ݬl�`�M��&l04W"�y��+��bE��?�ZX��	���yBa�+ HxT�P�ݰf��0�F��y2O_�<G�Ś�iK�c]��C!�y"�ŧ�F�١!�6[~JK�$���y�k�#}&t�� ��<�Е(ǡ^��y�	�;[8jq+��Kʒ$�#��/�y�)�Ox��)2h�	=ӆE+#�ȵ�y�$�S��@R���?5��[�HT'�y�Ob���h�N7z]��s���yb@A3\������a��"�$�yB�&w�Ȫw��^�����䀃�PyR �S�J�@A�2C1�JA/�P�<��d^7 ��l�4��B	z \B�	3C�8�aIZ'8����㐿!ZbC�	"���KW�"iI\�`U�L)w��B�$]@�J�+|@8��$ʞ���B�I�h��J�k{dh�!J�O\C�ɷY妑ɱ��~wvܱ�I��v�"B�I���EH@o�,�@�%mmI0B�	X;��0��&2���aA�-O%B�I'j���Qi�))�ذ0�K�<8FB�I�Kh���l'���4�Ή}DB䉅;<�x���͌m����f	��}S�C�I�;\H����M��A'����C�ɫ%~��1 ��C怞>�C�	"?�mx����ؼ��I*�HC䉿9��lZp�L�r�SÇ�{�~B�I�F�ٓ�jMc�hj@�J�3ADB�	�9�.�z֪@�)Ppȡ�#� *B�I8.�z���n�jZ q���#�RC�ɋ]��,sʆ.[L,�G��lLLC�O�`�_'���AE
�SS|��$?�[�̵�R�T2(v	��[�)�0���x/
��R<��t �!�����1i����H�>,wp�� |�",�ȓ�v)��+=�	x�AzF�ȓG���J���e�tX��1u��q�ȓ]��i�2F�[����)׼<�ȓ ��A�!ϱXr5�L;����O=�	��W��u�s�Y3v-����y�A�bOD�{����{���_^�<� ��wΔ@�,��z�*��La�<��f_�T�A��X��iW.�F�<ѳ�B>(<���O	F����WC�<1�MM����/��]^��'�<��C=#(�d:��
 D4��0K�b�<� tb1�T�/ݔ���i�\ؔ�R�"O�SP���q�tQcƘ���"O��H]|�4Ԛ5P�x��l�$"O�� ��'a�N �NKq��hb"O
�BAjB�Zf���WZ�n��q5"O�,��/׆m�<x�a9qh �:"O�5����K��`�1��8tR�@�C"O^����z ���0i�0p��R"O����ɔ@?*2�^oFD��"O�����!Dب��	i �"O,�&f�a14�K1�-$��r"O8m�&��o�s��f/9BV"O �0�n>,��꘬%�v�E"Oȹ����J3�Šfޮ�t8ۦ"O��sӃ�l�}r�Ä8Ѻ�yP"OX4�T�D�(���I�y���q�"OfPŀ�7�$Ģc�H�PD̻�"O",�!���!ٖO��4�@!#"O
qɆk��]����DJ(c��"O�<�T��+���cğ�L╀t"O��@��j�8uh5CL4`@�\p�"O*ؙsL���S��0*?��"O�y#�͛S�P��bD�,J��
e"O�Y��g,?������W% ��[�"O�|s/˵T���W`�h���9�"O�������;���2\�*@�!"O�Ź�C�z[p9�(J�4��"O�x
�F8!��y����C���ф"O~0��Z�4,��� ����ұ"O.��ǅ�c�p4���|T"O��0�����G#ЉP� ��"O�}��mZ6*X��4B����p�"O�A�S�̿/z��C �H��TL��"O�A�2�N�14ɛ�.ߤ���"O��g��]KH-��M�9���A�"O�4���+�`������V>$<�F"OfQ0��ߩ<f��laְ�C�"O^M� �W�qc� ƞ}���"O\�)ER
Y���Y@@D��`r�"Ofx1֫�%w��3�eR�*�r���"O��Ņ;!�6�b��?E�$�`"O:<h�/C�v�(�Qr��lְ��"Ov�K��V�1�b�j�!�"Ozp�c�^]�\��BE�k���@"O�yȳˈ` n�����R]r5"O�b&4hq��"m�(PV"ONTs`$T3 Db�AءSB$�`"O��k A��o����oM�a8�\�"O�pI���t�f���/��aK,8
"O��A�ʀ/i�(�6�HC_@��g"O�R�Ą�	b�����V"�k�"O$!(b�F)�b q����X�"OP|�a藲�`I�LEm��!�"O~��V�>z�P �`�G�˔}ۖ"Ozm��	^�](���G.? Ƅ�'"O.����/�6 ��ӕp����"OR܈�!ږ;=�P�8C`�B"O����b�?H����N��1I�"Oԉ�h�I��� �B�̥H�"O
i����o��Ѭ�3	��Ҷ"O0��6O�Ȗ�*�Ɵ9���"OB��@�G��ܽy#̅�~��"O.��ȼM���ī�/>�����"O��ia'#nՠ�!́Q���P"O� ���M�e X��@�S��m�1"O���gK�Fz����v��hg"Oqb!/�\�9��
�O�L`�"O@�c����P C�4A�����"O��cF2B��˰�x�G�#^!��&p� @Ѣd�\����!��J�F `;w�ϙ���I֯!��G<LM�UCޔ~�4��iڡ!�q���L�}� ��c�J�r"!�Y.���RF�EM�Dc$�B�!���&��ڱc
֒D@r��(�!�DD;�lAH��ĉd�����F�2t!�U��H]�gK܏\� �K�OO)U�!�<��J��]�EoXQ���ѳh�!��8����%i�l�
T�%�!�ٽ&�&l�2��P��['x!�؛Gg8���c�#��\:t(�.o!�65*D(��o��v�#T�Hj!�������,=F��`�ai�$c7!�dб'���WAV�^��c��\�f!��PT��[�t$��c��[�!�D��Pl����I��/f�\J���k�!�$]zH�cIO�_�XH#v�Q�!�䍿V�t@��
|�m"@�y}!�@�o�4SD�^�C�U���zg!�R�]�&����83�dD�&`��hf!�$V5biG
Îrg��c�Y7"N!��Mr�<���6 �c�� ,6!���50����Q�L� �ы"!�$�;v�D=�	�hC�hP�OR-y!��Zu����ױr)����F�d!���Qۄ��Ǐ�HL���� !�ٻ�|`��!7��3U�T*�!�[
(Fʄ���4 ��Ȑ7� l!���#.�EP���l=�D�՗]�!��.��� X���ԒE�!�Dĩq= E	�#LL�3�f�9[{!�E���'�ڒ`��ѹ6�R�>�!�$¹0��*� � ��n[#Vp!�]0R&��##��u��䑥.�	!�RSM*D0��PL0@(�-�	
V!�D�NM� H�KQ�d!��"��0&!���$
Q���C>q
X�#!,J�`!�$�*;�؛t.��\t�)!�Ɋ_!�dEc2�1 �����A�@ s!�
�hU�ـ�ȣ4ӊ%R�?�!�d�+)���#�%,��Am��=!�-J#�8���N�t�:u��Lɽ�!���)	j%RS�ܗ-���p��T!!���/]x��qT���Ԟ�6�!�DҲ�@�#�n�99�t�y@߽]!�D8!�-�vO��s�V�g/�+{�!����"1\Ԩ4�Ó&�<ha��

z!�S�:�L0���Pajбʣ��!�D�,`�4H�����6�c����f�!�L�ӴC��LȆ��b�]]!�9SM�Kv��0�ruC�d[�>!�Ğ+wt٘�F�!{6A
�K�w#!�D[2W�4�Q��l�"���K��n!��H�rl����r,�@�1�3�!��	l�FO�%>(���w�H�f�!�DPs��K���9(��J`k��A�!�D;;i<y�O�S�v�PA!�0�!�d,=xv����We���0�f�v�!��  �p���P�P��u�\�
[��9d"ON�9�J^�Z���
-)J�y#!"OBms����ذ��^3b��G"O|4{�A� ?_�rҬ�3zA�P"OR=2ׄG�3G��xBL������"O��"�)SC���ê�f��@3b"OV\SW�$�I6Cӵ;@Zy�R"OpE���4Dj�UdN��Ty5"O"����5�4u����@WDAb"Of0����qd�`�+���h���"O|��BdE0GXzD2d���E"O"Q���$)�l�9��ڃ.�ΐ`5"O�Gh	!;颁�!�����"O��!BG;E�x�J4
��Oq�X��"Of��+�">W�x�pb@�
E�"Ol-(B��z�I��P�K�R1�u"O�y�H�/,)�l�gK�9à �D"ODQ T䌒�,���CM[̒j"O������
��Y��1�"�""O0���U4��Tq��W7Ff�裠"OT�"臌 ڭ�1�S:f 0�"OB�:C����`3u�_:Vx���"O8�p�$]
"���&��	pTb�"O��iE��~k"��a�&C0]s�"O:p���;<Ft7��g4Qq"O6}��G��o(]k'��%��hc"O:�3���\!���h��m���"O:P���9���h!��Y�6�2�"O��3C޴E�ԥ�%�����"O���'�}���h$�8T2�}p�'�vl:ም�㲑���̄E�Y��'��<Ȣ�6*G&e ��;K�2��
�'�R]WN���n �.Z�?Px`�	�'i�%ӄ愵̒T�`!ٺm���		�'
�GL3v��M�%H_e�����'m�Y8ШH�B�&Ye�P�[	2�a�'ۖ�@���x�.����	Y�P�'�L(Q�߽	��T�4�[,PQ��(	�'Î�Ǆ�f|"�!���X��M1�'}R y�G�,7�8'��;>�l�'��)�*ψ,z*��k�%'y8��'(�1��ѷ+<�1E��,0ެY
�'"e[�
��V}�E��##|j���'{���J2V#`]a 
1�6L �'��(ڧu��� $��$�b�P
�'�L)1�g��qI-�`X��R�
�'���)�(�1b�{��.�,y	�'�ĕ���$�Zh�Y����yb��O��x����(��`���y�&�&B�,���޷�$�0F�y�˘��p!�T��*g�{SA���y���k�����
^<!����� �y�L�ܺ� P]�}V�����
��y�-C����Ҥ�^B q�ի��y��/$��A�f,W7�*�"����ybD�բ8�ڀ5�(��Ð��yr�0Kʹ���H�8D:�����yB�,�����R/��0!�j��y2�C�BۂxQP'żzrf�g��y��I�h5D�ϖm��m�gBϳ�yҭR3'k�;�3_�I�C���yD�Ӳ�H����T�v�b�����yҤ�#�PcuKG �z�F�y"ꖦ#Ƙ ��=�������2�y
� �m�gZ��UQgK5�pU�w"ORm"�Hʾy��(� �G�HjX�93"O(��.O?\��ɛ�mD5Zq�� �"OB��b��d�ܔp�+�;\�P�U"O�1��ƒX^l�j��7�*�+�"OR�A%��"�>9��o��.�S"O¸����M��9eH�B�|��`"O��YX��0��r;�L9�oB=&!�H�>�X�(O^-�1�gO�
�!�R/7��œ��X�; l掆7S�!򄟚/��E1ӎV�*�Zmr�c�!��H�j��\��� �&Ű3�W�D�!�*���D M�&8XT� �c�!�͛7J5����*3�di0���3l!�䈴_G��!�/֒	�jq��C�!�DT?�~}9�h�),������V�!��[��.e��A�ن]�0�E$*�!�ę%���T�+k�8�E����!�I�@2 ��#$M�Y1���f�!�$��!�t��4�R���i�"�!��)cTYhqB�{�*B�h��"e!��](G��)���� N��)�n[wd!�$��
�������}>��1l<UT!�ˍ�FY����Fq�Dj�K�eK!��6�.az��St�$��r!�DVȪ��۪7���Ȱ3�!�$W�W�YؗfL'$t��/w[�'Ŕ}�'��`/:�1�H7o��)�'�z���Ud��y7D8XjH��'���wN32�婱���P�EK�'�����f$����N/Ch����'xt���F�V3`��0j�a��'���b¨�~�q����d3 Z�'\��X���`��8ա�+�2��
�'ɚ�"6�J�O���2$-ӫ$($��'���h$�A �(�EE������'>8���*<���@M��G}S�'�6�"uI��5e��*�a�'	R����'���""$T0Dz�tʇ�Z�����7R�|��UH��[��2c���ȓT�� a��ͻSo�l��ǰ:'�L��u�x���Ē�_N���VbI�u<D��%%�>2Y���̃|9:u	�'D������O���JgOWD%6�:��&D�H���5e�v�SD�B������I%D��J�Ոoc�������d~�h:�!.D��xŇƘ=[�T���C�E�Ѳ��*D�xc��n��<�d�$C��VG'D�taT�Ь��W9j���ǣ7D��yBjEaǾ����G�r��Ps�0D���3H��W���dE0m��M!D�,VΊ��%e�D(0�aO�(:!�$����ɠ%(G�$%��bW�Z�!�D�_����dRrix�ߠ>�!�Ƞ0��d�UJZ�L+HY��^�{�!���+K���ر�RA�|Z0C�t!�DJ'N`ꑬ̫�(�бǊ�
�!��4�H,���vوĀa���}!�$�W�L��&dD���1�^!�ʝ	�DmXч�`��0b��7�!�$�+W��9�(ߌ?��C$�[��!��	$���Cw�_�5w��i�g�P�!�_�C4V��@�:%~vyj����i}!��<�nIA���v	�%�#�ƌB�!�� ��Sծ�hE�����^�yz,\"3"O���3��'bz��@d�b����w"Of �$�W ~�������9q�~T9d"O��c���<7 �kv�Tr�E#3"O�ݻb�Ȟ�&�R��K
 ��y(�"O� z�
I	Cl�DQց}��t"O��Z �C�&M0B�A0[�
D)�"O   �l��\-�ap���JP��"O8]�%�)Y��,a��^1�"O���",JC<�3�EQ�!�>�a"O�U	�n�:f6]�D_�C�R�"O��p�ې{�h����*_34���"O���+�N��{��6LxY:�"O��;to��CA6�XU�Q�Q�lՂ"O ��C�*��d�T΂*+�|�c"Ox0��Β"�vD�C<V���C"Ol��q��G9p�ZҢ:9͜p0"O�L2��Ԥ$����6c����9�"Of}��ۢk����5��y1cc"O����*���jQ��B��!C�"O�tс����� p�]:̐�E"O��2�؂f21�D��1��Q�`"O>�R$�E����pd�նv�<0�"Oh)Ac��00��5šFr0�"O�I!#��2���P �20���"O���
4s�j́�`��q��$)c"O(K>z�!�.J�Jl a�W"OQw�)l`�Gn�4ftX��v"OP�S�Q�dX��mO�"g4�B"O�S��8L&T��Sm���R"Ofh�HZ=/��``$��_alD��"Ov�1�A��*�+v�ß�fhKV"O�8��AR�8�<#�0p`PJ�"Oڌ0S'�.X!l�������"O����%Ʃv�b�Qa�K�c �MB�"OL��bҔi��t��ظz�k"O�`���ql�i�@�r��Y��"O ًuJَai�N܅Z1̹J�"Or��a'��&�0�Jm�=<Z�y�"O�<�B�$L����"듅%8E��"O�(�3�p��`:8�Tچ���!��Ӈd���Q� �w	p�!ë�u�!��i&�8Ҕi��-MpE�� B�)�!��|�p�Js	�?? 8��@Oˇk9!��� Vg*��J�]���W(�G!������Ḷ��s�l�'v�!���b���Kb�<�b��rk
�3�!�Ѭ)�*􉧧R�K�^�ɔj�+!��Z-MbL�P�Q��䠲�Q�j�!�D�,���C�,�B�	���W�y�!��T�u�|��"�Ӿ3����a��1�!�d[�/*&hb��=t����B���w�!��9K�dQ䫗�C�(4�t��Fx!�d]�E�b���Ł
�v�k����d!���]
H��ը�#!������ϲB!��e�P$9���<Kzqb��5!�d�29�l0��I�6Y\�G�ӧ�!�*mӲ�(%$Y��k!�ғ?�!��\�i(�\��AKTKVT��,$D|!���z2�t�b�L-�-���]�vq!��Ebc�9�sK:~��x`p
�>K[!�´~�R����#��}�P�j	�'0z|�G�
���9VeC)>?��H
�'��i:�@GH�Ai�W�jY޸��S�? 0 ��j�|\B4N�%�F	C�"Ov���+Z�#����b�_� `R�"O�		�"�門bfl�.����"Od��4�ΩjǼ�����;�JD0Q"O�s�Y�RQ^%�&!Ō8���3"O&(ˁ�ݴF��0���!C�B��"O�yy�c�.$�!�L��p�xC"O�!H��GP��c��w�A�"OhQ8�Ϟ�#-�tKQ#4wlx��"O(�;�IB52Y�a�QqU��k "OU 6L���d��!�V9><�"O�и���6�����\7�Ce"Oέل	���}�����8W"O�H;�b�0�5 ���>t��"O�A�&$Xd\��DƲqIX�AE"Of]sabHeаpe"B����"O8Q��&V~��}�ѡ�;|c��b"O��1��^�$w����
^*x!�"OJ9xA���).6۱���,���"O��1�#(+�6�fc�^}��1E"O�ӳ�M�z�r��?1��"Op��� 
�E�]�~��"OFy���ݾ|LDaEd���D��"O����a�,����N�Sx���T"O��s�}��p��ؑF6l�
�'">����YP����,�=v��
�'`�e�w�];?�&��S.�Z.�$�	�'��9h	F�J$�Ӧ�7��8	�';�}{� P�@���y�`@�����'pFd��b\{�Q!��p�V���'�y@�Q�Z�V����mj��'+�$�p���*��ѯ|;&���'m��J��D�yX25�5n��q��'��m�#�[�&�a�U�Ҥ	�dh@
�'�C��
���Tm�>���'�Ι����;T3~�Ҥ$��f����';����N~<��dmǥ(
Bu��'î�B��[u$�0*#W��T�K	�'&ݪpK\l�`�<n�XJ
�'���R��A�m�����.{΀
�'�u��2�R��D�ҽ!7V��	�'�����iJfʰ����.��'���!�ϸgj�-c��`�,R�'@���Ô2��t"05�"��
�'Y� `�k���`�(I�M�
�'�H(c�S�h�J��%g�$O�n Y	�'?x��G��aR|�*�4J���J	�'~ܩ��E^�V�\h�F�1Hv��	�'G،�ːq�!چ��2>��'�b��w���mk+Q/i4X
�'b�d10>L�5�R�MP0���
�'\�P�tLӎu"��
�u��-j
�'�}�AIӲ|�B�:tEh���'aR��3˂+<x�+��^ s� �2�'�(T�3:�L)���� ��Q��'��s��X�^�\@1P��?�Rܨ�'�f��h�ApbZ�ʝ�� #�'w��9� �9PXj+�\�`���'��@���y��Y��ȟ�TX�,��'�\�h�h����Ж�I9C�6�P�'�8E���2C*��%��;κ�b�'#z�����|�����1�҉�'	*��D@وA-���A
W�d���'���1TE�8fe0A��'��J�L����� N��ǟ�AA�\����!Ks�H"O��#�eҡ\��i��QId̍kV"O�T��25ej���ɏ/[^�k�"Ot�!&"�{�Y�g�+zU�<�"OL�h]h	8qj�4<�~80��F�,�!��ӹ5܈P#` �0p��]�R�I�{�!�D�)/h� �@�p�z��̏j�!�Ĥ�Ĭy6�� �Ԉ�sh_�[p!���_ad��#�%D�
�gJLcW!�8>+��R�.\���c���!��U�g "bD�G �:���
}�!��+20�P	�s6�A"�/W3#!�$��c��Xce�O�ha���!�Ğ/(1RU���^M�ԙ�߹!������.Q�5ڜ"����!�Y#|Of1�ԊJ�90Q��
�v/!��"r��wcR&1o^0a�� �( !��0	t�I���Λ?W��[��z!�"X�Uz��3{��5�!t6!�$_y��R��b��c�O�)5!�d�/�hy��J1HΑ������PyB%��=�4��M�z��u�Æ��y�_�&.d:��j3����C5�y�,�E�8����H(���B��yRṃ+g�l��ܽY�fU��g��y�G=M� p�S���Z�N� �O,�yR�@sW����$ЈZ���+�cެ�y�(�/�43#"U8\�ԩ�s-� �y�I��;�<�pBʑQ$��	��˝�yBi�YpVL4�0�($� n���ybOϑl�V���3�yB��M�yrK�l���^�����T$T4�y��1|�H\ �%�L)�k^��yB/�j�hY�m�5	��g$�y��2I��a���O�`�*�A��y"���w��Y�R���0J���y�ŝ�xU�h��"�:<d�EX�K:�y�ς�MÜ%Q� ݒ]�ޑj�$�5�y��W.�tI*���?k���k��N��yR��J��0c�Y�xz��*F�y�+Y,���Δ42��dŇ�y�l��f�����z3�m�"�yrkL�y�p	�f���D�PT��=�y",�?��ȲEK��o����c�_=�y�lX�|K���tNE�j��%*�I��y�B��Ag�'C[k���Rl�!�yB+�2���jCg�M�^���/B�y��ӫ���� �КG��Jb)�y�H�.�Tx�
ͩEF0�x�%�y������'�8#L3��A��y�ǋ�(i�|yT�C�fvt`�C��y2�D����dL�:U^V�Xq�y��%�t=��lFW�����j͵�y�O��:��i$;D�4!0ƎW5�yB*�:ǈEK���r�X�W7�y��,4v]pP��5}�L�k�8�y�ZKʢ@ڗ(� q�A��ߝ�yҋ�$I�y�a��fz�=�&I��yb	�G���F鏨3hl@G�4�y�)7�B��ӧ	�6��wc(�y"A13$�zd��46J��߻�y"JD�[�LCB�Kf2�����y"Ɓ�g��TR��Q\vz���y��&Id�gR�Stl(� ����y
� ���B��4� ")��cJE�`"O�m��"\�KS�P��o�м2g"OHt���Ád��8bЈ�k�i��"O�����?P*%BDn��Z�Rp{Q"O�|;�_I
��M�1���1"O��Ā>D���#�9o�P�s"Ojl��NM7����ʛ[3fi"O�%%A��{��m���F�p�6"ONP�m�O�,� ��q""O>ñb��((%���R""
�P �"O� �%P�y'L�S�H�;����"O 5#D�&dռ��
�<�T��"Oz��"��l�v��s�P�R"On�7@ϫ)�D�B]$��T�"O���P힭_U������<����d"ON(z�,�1�	��E؄S��q"O��&(�>�ĉ�B&ʢ97�A�"O�Y���mV��RT��;4�h0s"O�A p�G	��A;%L��P҂	��"OJ�ԎU�"BĉJ�/�:t��"Oj����˂$��S��%����"OZ���#�R�s��� '�Fy�"O�+�ڽ+��Pt���̘�"O>�JA�	n�"�9D��`�xA�0"O��l�	KX��2��`Ȳw"O8���@�/@
8��[�p���"O�0�΄/oH%@��K�+O8aq"O��'U$r���"m�� ,
(ٔ"O� Ia��6�`�B'����R"Oz�yT�)(\y����vY��"O���Q�.10|+cő*�j��'"O��$f"X���Gx�}ɵ"O���sE���n�.\S��Qsq"ON�i�Oð0_�9��Q�E�H���"O�p��7 HxQ�D� ɠ��"O8��CB�?^�$ؓ��%%��ً�"O�x�OO�3R���䒟2��Y�r"O�l3ţ{O�� tb�8C��@�d"O\��d�7�6 !p�σ%�0+�"O�<	W��J�V<z��M?4�`�"O.��A�el�HDj�0JL�2$"OxY��ޤJˮYQhO�J(���"O~�a7�7{��a9���^m��"O8H8��	��t
`$��c�>{�"Ot� ��^�G�~�B��K\ʎ��%"OЀ�@	�%C�Є�_�GԜ�"O�9�	:|^%##�O�$|��"O�%
�Sn�!�a�� "i,�d"O����E�9:)Dt!�E*_2`�"O�� D���'_��"�=p-T�s#"O����'�>h[0�w�����"Oƕ�#�������H�A�.���"On��$	܈$�t��m�7t��b"O\S�!�.6���Y�@�9k6"O���waQ0u~����(����"ONbb�\Ŏ�{�m��)��%�"O���D퐥4��uy �SF�� q4"Op���B�g|��nȋ4�jg"O�,��I�>�x�.���0h�"O���p�\u�.�{���iv"O*�Ӧ��q��My���/	�Z�00"O�T�E���(Ӷ���`�$��"O�e�2�ԙI?|���L;NxrS"Oܨ��F?'Ӱ�c� u�=)%"O�  A��fAm��a���\.0^�d�"O`�0ǋ,x|���p�٣fP҈�'"On��TD$C�:�@� ֌�RQi&"O����?ut��ńþia�"O�8�IҲ=b��:��>����A"OT�����r��8Y eM�]�>H92"O����#+���s�X�")�1�"O�D*�ڪz�<�R��V)+��dI7"OhD�VcK5L޲�r#B_0���H�"OP4�$��'p�D�����i�(�r�"Ozy�'J$z�^\�7����"OD�I7��=:ϚI�oI-@zL�R"ODAy�o��LT��u��	>R�"O�P4�H�	�JĻkM6}�"O��%�Z:��4�X?x:"O̬j"�X�u�.M�@G	�u'�&"O�j@'���q	�߱@Pa��"O^uqfil��g���YH�"Of�[Sd�$��U��ڪZv��a�"O.����Jv98,�V].}7���C"O���&�49�&e�WhS&
>���"O�p��fܢg��5Y�,�g�3�"O����FC���;D��;+r�@�"OB
�!��7�ɡ
�GHr���"O�C-��T����C V�Z�S�"O��A۬r`�(S�D�%�]�1"OvЫ#d ��1���0�@H�e"O�ԱF��Ar����ݮ{� T8�"O4�@��9E&a{���?���4"O
$����=afT%�JT�V"OL�zQ���I��aע�m�2y�F"O�Y`0-�wݸ����[��)�"Oz�1��4��`z���3�J�"Oj��!H@"�Xa�N6O��}��"O�!�n%4B����.�r�0YP�"O���-��GM%+�: �c"O�M�"!w�X0lN"Y��M�G"O>�hvc=Y<�a��(Ok����"O��j�/�y��q�d園 Q�e�%"O~�	�G5%a��U��+�޹+"O�]CbG�L�M�RDƲA�����"O~Pi�	�A�^�
�b^�[}J�X�"O�C���R�d cc\�jX�-Y�"Ot �F�.�YA��<W��`"O����E�)��I�A�8|���"O~���攄uD��$��'U*Z8+�"O^}٦#ʌI	d�j�+�\���"Om�m�%^.����)"�"O��P+�6=�RiSw聭"ڐ`+�"O�\IC/�Ip�gȕ�Ÿȃ�"O<�8Di�\��'��g�h�r"On1hT�9�t��6�:���"O���`3P�R���ԓv��@("O&�d�����W]D�4�9%"O:P�PHP���)�"L��P@"O��z��)xԪ�B���x�"O�M
�. h�@(Z���4f8�Z�*OPD�7�[�0�"5�B#%�p�h�'�:��"�37H���.�"�9�'W�ia0E�2i��9�cF�!�
�'�q P�{g���B�P68@ܐ	�'�!Ӏ�0ڬEG�\I��3	�'�HK���,�l{*��bB�I��'Y�����Ω|.p��°V|Tuy��� �˥�#|�hF�_��l�3�"O�<s��GK$�
`�P�2pP�"OBy!V�\̎l:�m�		$��I"O�LӰ��'vv��RV��3��m�$"O��v�H`iJm !�������"ON�H��ɀ�VŻ��?:���"O6� �˛=_�����J�?��w"Ox��WcT�VUX�f���%F���"OBM�D�[J`-���y&��N!���4)A0��I��5k\�B��\
!�	g.�|;eEH�V%Q�ƻx�!���u���UN������ �����.
�V�P���RfVD�7��9�y��čI��Y�.܍Jt0Q�E�;�y"�@��ĩ��=id��֦_	�y2ʈy?��d
*%D����y2p!^�h��:2����E�E�yR������4y`Ƭ)GƊ�yb��mں\µ$ם`u���DFJ�y2�ͼ���K�4a����1ǧ�y�Oպ|9�oJ�p[�]qA���y�k�4	6���@F�l�����y"�ّ}bVQC�h1g����$ �y���(0������A�X���#����yh�b}r8҂i� ��#���yB)�_��5p��y��81��ޔ�yb���DƴK�n�<\E];�H3�yW;�L3���d|�qsʒ�y���p~�;3X�a�@쪒G_��0=����W�ej��≗�)�� �J�4�yRʉ!z�Bt3�ա&��4�(��y� ]C�Z��K^r!0�k/��Oڢ~B2I����paΆ)���i�hR�'��x���
F\���R�$y����ybf��?���3n�	X�Rh���ј�M�#�'q�����Y������B�����'e�$(�������1=
GT��� 	 !�$�6���c,��n���"�F)0�!��e��Uk
R6^����4�eoa|�[� �	-H��K��`~���H�aL���p?QV�at�z��l�xa����[�<Y��L�ytX+ �ӧ"�h�@doW�<	Qvެ�˴k8[���D(
QH<I����v`D�cie�Ε1�O�@!�d����7��?���h!c��L,!�:	�E`��AX�ZB�oA�C��F��OFީ�1��]X�=0b���y�lT[�Դ����H�����y��Ł*	�؂�I�2b���qJ��yBO#f����=A�P��M��hO�����4�l-�W��j�����oH!�
,�������*�����A!���xԐ����fZ  g�
��!��f2�맋"D���Ӊ�;�!�C~����A�4&�<��)K����)��}��j�p��� ��AW�����&4�����?���� 5RqC�K��KM��Um��O�p���8����Q~\���-ڽr�Ji� �5o>�%����	��B|B�͍^ݐp� a}�B�ILJQ�4$S�0��	��#C����>)���]"��&""j��҇��H�<�m�T�Q`��D;��	�oXB�<��JQ"8LHhV5Z�t���-�Z~�xr�� @�j�Ȃ��y:%�7�*��c"O.L��	��v2�i�S�G6��u�s��j���I	9=N��f���N����I�&x�!�R<n�&�{�  < �"�Z�'�!�D_
^��ѦDՇ��A��M�:Q�!��P�RY�x�j���ؼ�%MN�#�!�D*m���`�Z���H ��9����'�r��n�����J�.$P�e�>�y����S F]:3��U8%h���y2��6R�+�`�@�2<�s���y��tqb5� ����q)�$���y�����"=�"�_�60����X�y�	܉yU����m,40`8vl�7�y�㚐R<m ��Iw��[���yb@��,V|�ǂf�����߹�0?)-OB4�q`nS��xR���ƴP*"Oa�Bɗ<�JD�f��;���*��'#�V7O�=x�GU�u��)���	i��˥"O���GM/ި��r���q�B䁃"O��8�C�2g�H �AO�{$*��"O* ����$m� ���!�A�D|q�� ���(�r�^0���Ȳz�����:� �ȓ*X�)+��-v֮�*v�@�l\�O^7�?���'f&������!���@+���	듷�f�L���*%U��Av��@�����퉳���2�i�X���(%l>�P���.�M#D�W�3u4�@pס1>��a�B�I�<��ǌ  �H(�%^�`<�Y���I�<Y�-�9qި���[#�|L��'�@�<��m֕v����T�.���a�f {�<��I�U��'<k�.�*�"Hp�'�VDD�ԩ �{�i#��1<
x��E��ē�p>�&#���2���2R�H��h�P�'M�~:$J�(^.l16�r �	"+�M�<�`$5'D���֎n2
�;g��E~��'�;3i�f�.�)ZR�˳nBm�<�ӄ���xt��4D;�9�"h�<Q�#�'a����'9^dR�0Nb8�$Gz�DA�uͦ�"	Z"x�ejpO���?I�^C��B�X逬!"R=��ȓ9Sҍ+e⟩{�H�7(	>���LEƕQǦC-d<@�cB�W�r��'���*�S�=��y[U霶-rj�mO�I]nC�	$"�0�`,�;.j�s���/b�B䉎t<�����xl�`S!̉�/�B��+^q���Mސt昜b���!��� ��I
^.ƐpW�^ ւ�:�E�
����$ �	�?��!x��ܗ�(h���e��B�?ؘ��a�#j�:�Z��Rm���I�h�?1����&f�R�(_)`��x(�K+#-!�KjN*�kv���Xl�1Fz�!�Ӟ@� �2b��1A��hc�J��4�!�dCA}�(q3#��%�.�J�O3�I\������ ���ȱ)Y�I���𩠟TE{��)��f�F$��L"�R7.եl�!��'ޕ�"�ޔ[��f_��d:�S�O���a�\&8��I�$a .�#�4�Px�!�1X\�
惘�:�h�Eϻ�?�������i��D��4�`l��A�Id��$�@E{���OƮ��)7�Łt�P䠀��~��'y�O#=��;kV%�1��7!v(y��Aܓ��=钧��*d��Xr��|`8A���|�<!a P�8���!��� �!gFD��yR����X ]AB�����V�>�f�'D�� ����G*d�	YA�1-�Ai5P��G{�����'@0 �O��5���P�,�3!��N.w$Q8��@�m�ұqc�؁{��G{���'m��i�.KY��(@�o �G��t�O�<E{����i�ȁ��*^�8d���'xa{�͂�"g-�"+6E�oЋ�y��MR%�*�CJ�t�b�Ǉ%�.C�Ig��<`�Ogy@-"'G��!�^b��F{��$�^�I�4�֯�6���;u@9�yb�P�
�*�S!.*:a3�����yr	�X�����1$t���i؏�yHR�<˒���E�T�+'ꗌ�y�M��q�7g�724���ΐ�~��'�r�CV�.~�2d벆(�,ё�'��aǲ%{����
�<��Q�O ���m�~�ʢ"�X)c��(IP!���d�j��z��M%���
�'�DLh�m�KG��â��JS����''�!�EG�
�z��ȋ@�Č	�'�(�1Pl ���u�)8�j���'��d�e�.n���H���T��'�`����a�΅����h�H�p�{��)�i�B�Tɑ�V�f���"��J�!�D/q�*P�ӆq�5a�,<��O^�D=OR]�WN�c�����ſBeR"Oر�s'U�qr$S�뎃N�亐"Ov%[`��-	s�;��/�" �F"O~�P�D:\����J39��+T"O����58HT$��/�6��}rP"On��&�)>8Zt:v�F�#��(�'&�T(!�������e��'����'Ϥ�t3RL�a��]� %�E�'o
�H�#��<Ex6&�rZ���'��݊R��2 �}a6��J@ ��'&heK��ӚO���X�"�Tq�PR�'��ec��6dϬ�[��J�P˸9��'<Re��D
�XA��@*���1�'=�}���)�������Ш�'�tP�gmZ�"p��h53�^���'^4ˀ_=r!N9y�BF'-n���'�a�,���!vn�8�k�'}��SA�J2,T+�$�&% �'�R�� i�O���QN"qژ��'��}�p�ǫ<d�)�n))t�J�'��2�NJ ;�����1=��'oX\ i����y����D``�'��s6m��
��q�$�p����'�ic�*I�#������R�Wf0�0�'�<�2b��n�)p��ڙG���Y�'A"=�HM��f0�5�Z�W!�t��'�|���`�s�T,V����'�]���6{���* R]��'s�P��XB�Fl�)��h��'� Ȃ0���G�fL��YgL��'�0�$�C	!1p�vN�:/�
��'+��3bϚ\�=Qs��8&c$�
�'i*Y8�A��}��r�F])2�H+�'b��T	ԠJ�x�)����Dm����'�$��5-R�_aL���
<o�@]��'v*�9A�[� ���E�(\���'+6��c��� JTC[�~��U��'����J3�b$H�	z�F@��'&젣��A�U�Q�J�p��qz�';T���J�$��ɻOY�6����� �e�d�k�^�j!�6���ꜥH����V�'&��(�M�rL�V����'*���:`��e��i�,;�	�ʓXԜ�Ku�S�5"���
�"s�Z���9�d	GnB"��I�I���\�ȓV�t�j�
2:(��B�RӘM�ȓ��B�-�#)UnгI�3G:v��)�!D-1<�b�M��M�B��ȓv)t����P��h\��i�%	�े��>��&��|�ҰY�j�-7����ȓNʜ�V�G�j���+�"Vy{zE�ȓl\�x��)L"2 ���6l�>��܄ȓ1b���CB�/�4�ZiV�5��i�ȓ�u�%�.?��Æµ���ȓ&� �2g��K���'�%K]�ȓd�aa�iX�E��M��̈�R��ȓYxDѡ�F�.F�V�C���m�ȓ{�
�@a���
�ư���~������Z��A';�~�r�Wj
��=���-ƞ�i9�
݋���ȓ\��,� d��Ur������D��`��]K�@Vm܀"�*���h�A�����it�5���־3]B��$��*3��I�ȓ^̤�q&�V?�@D�R-"��M�ȓ-h:0�u���t��c�B館��=t�;D��,'�AK���z��H����s靍7ΰ���tz����z�� �NX����_�(������fG�Z�����@ۊ2U�(��$�\�f(�2A��j�
�t�����]]��,,
�2ǏK5
�A nMQ�<�T�I)mtjthQ��
X	p�Zu�<���J�f(p[��O�W�Fŀ���r�<iaI֗TO@�2�)�'Q�ڜ���q�<A'*F>R1����͢`�� ��nN[�<�%�
�G��
�陜{�(cg)�V�<�R�J�!�����X D VA�OP�<a��ǋ^�=�fl��I}���@"_I�<���	X�d���w\~$��D�<��B*��s�7���e�~�<q�Q�c.���̇-/T)�1�YL�<y'�[�M#0�#��ܸ p'aAHy�*�F�tt��	=9��|�BOT����h�I�x���A& x�IpN&=˰��Z�\�Y�r��Q �k�'���i�%y�h����Y����ڣ*<�	���H��?U	���p���ǻ)߶b%D��A��؝T���h��^�Y��F��e��q�/�$�^��'�>�	*�<U Y�C��Q1�Y0s��C��6v�M	%'Ƃ PLH�pHT1?E����RtlH�Ņ&�L��X�L9)��mH��kD�N+6�Q��ɴ~���)UC2o�~�Z烞div@�eZ0t!��#�L�}t:��+MBT��L�;}��!���jU���>9��|}�i���0A��0���O$1�Ru0��A�f���H�B�0�y�Dų�(�B\(��U��T�0�s��ű�2�*4$��_p�	�	��H��ɾLv� ���3M�&�b�̟�	bB�I%?��5�O�&A�*��*�m�[�#X��]z	s1�6�p<��"_�T��J`�":"y贎�c؞X[t�G&
��ԧD<u�>8���Vq���C���t��M��s(<���8A���F珛0�V��D�j��L4�!
_�M�u��K���O���C��,>g@��"�B }-����'��� ҉W�,���uC;ڶ���I&�l}��/P8_30t����H���/����b�o�8�:� Q!1�C�	}d��b���!�i���";��$+d>�X�o��O�R�9
��
\�%�Y:d�h�ԄF28h��ɶON`0Ca`C7�P� ����KH�<BN��w�Q�-�B�QA�~H<	�
5sh!Go 0>����΋P�'P�u1B�U�o� �R����{c6���oAS��ak��;5!�E�b��-��d���,S�cK�n�X�9&��:LбjP�>E��aP�tɓ@$�����)Q�g�ȓG`��0ѝA���A�ԣM���'v�R4�FY؞L)�h�ox,; �	S4���"+D��8&BU�M�l �"B��{��ɂ�2D�Tps�[�MD	 �C��.��:�.D���A���4��.�	��,��6D�`�3��Jv�,Hִ��� 4D�� �'@(`�
q� kaL�2�%.D�0	čϗ)����p�٦X�F�Z3h2D��9W�ۥ1�PE㝟#�f���D-D�<c'�zb��qr�ڳhl�#�k?D� Z���(P��7'�\��I&D�Թ �ڲd2v�[A�"�$�Z��&D���4�؅	 0505& _�V1k֏�<��@��0>�hγO^R��%�7�֥����JX��ceǙ4��nF�P��q�B�{
\U*qM��y�E\�%����#˺Ũч ����̠���V�c��S�i~�̧'���3ǐ�g�C��l�X`�K��y���HUOZ�d� 6��h�Q3�����)�>9�eĺ].PX��1BG�D4�}؟��G�k�9ȷ.��J%�p�l̸'��L��?�$�ȵi���IS��3�x`�`���AB\��&`]�dJ�tF~�Gs��t��51�I���][��4������%Ld�l#���47Mh�H�HT�,����J y8'�O,g�z��'��\H�ȚeKb*��C9X|�1}>d�S�ɗ��#��-o A�ȓu!�����&J��ł��ĨX
:�%����A�Y�O8�P�@)+m���$M6����'�XlZ�%��(�t��@�&��#Q�$MQ�bjd����a/@����� ,�"�b -�ax�6�Q��4cdI7d��	qef�L`5�ȳ��?I��E�vc�����k�i�!�[��;�l�ȥ�<9�H
��-)��ُx��pa�HW�<q��,r���@�\?HAD��L�=J�<�|�B�W�16B������`�Mh<���Y=d��OV���s����m���F�c�le8!a=6�N��$��W�F�����k��k����2�azr�M�R�Y㠖�_����5�8\�5�ܹ={�s6�K���A�5(�<˦Ȋ�JT<$��@�;�O��2p(D�Ҩ�;ʧO#�AHpʲ|�~��jǤT$���ȓ[`��k�f�Vv֨H�)ףhF�p��GDH��CF7D�8����W���d��N2\��aL��*l�%�u��wSh��f��Z�)�E�h���%ߥ2��L��)@q
fMًC#J�a���1_.h�ȓ�t� ��L�` �O1c�D����<����/�]��`А2P�@��`>��@�	������Y{����4����$̇c	�<1���i􄱆ȓ`��R��)Q�v�Ȑ���)��$�ȓ
l�����fT�`'*A�N1�ȓkX����X�^!��%���P��]�гu�X:-U�Q���A���ȓ[��4:�8P��elQْe�ȓtZ�S�Jm����- �쌅ȓ8��d�֢��%qCG+t7z�����lh�T�d��I˜4��1��T�\J�P������z��O8�(����wX,`;���c�X"OnD ���� � �B�Q��g�I�6�:����"b؂!���@^�]J��]	Vn�C��6*B]����m]qw�"IS�}X��qO?�)� ��B��\sT0"îώU�2��A"O(���0g�&��w��$��%8O�#F-C)�p>a �V�ɂ�� �޳�f���a�E��F녿��$�8u�4��$#���;P!�4>!�d�#nJ訩#���G��;��ۭS�Q��"Rc�O�DP4��>s�F`�ԃ@�H��T��'h��
��'�`�K$�̙1�0P�'�t����?�\����f����'.��R�ʞ8'��&� R���'~�Y��!�p�k�2U��`��'~҈��� �&E9 �S��\-Q�'�\�٦m�/���T�O	{Z����'n��{��̠ ���"���j�p�J�'e���#.��Lw�L3���=X�[�'���Ӣ���`s���1d�)�
�'I>�0�E�M��ИA
W�d~@��D�b�����->��H��U(V�0m�ȓv�����M S:x��r�P(2V�ȓ1��0�KG���F%TJU�ȓ`�fa�(Wj.��ڧ
;6jq�ȓv<;W�L��hۃ(BK<���2&�8�$�L�l(��e)��՘��ȓnKjH "�6p?(@���5ְ�ȓI-@;��w����ę����ȓ|lA�Ǳn�s1G�\B���/���qd2s�,�gW*#��1�ȓ3�&����6j��0kĂ:Y�l��ȓ ����/?����e�r4����~��dx���,����J#C���ȓ>�R����l�lqҤ�R�y�$��f����bP����Qv��H]vɄ�A���3�E-�ȄQ��+���ȓc�|%C�LA�����%HF�㾤�ȓ$s��P��RJ�� y�@�-e��i�ȓ7g���)^ �n� �%ۨu$��<�BԃA��S�FE��LI%z�-�ȓ<:pq�"iP	�@Q�Ѧ]��,�ȓQ(ѡk��~�1BW�^�,h��T�$��%�l����@G�`����sT�i��|�@��+p*��ȓ�H�#���0JYx6�C
O:j���#F��b�Ř�^��HB�߿J�P��_��
����q�N��I�<򔭇�p�j����n@�W�8wM��u���K���-A���*�Lηf�d ��E��=S��%Z��wM�uX���jUč�" [`MJA]�\4���P�R���i�4t�t҃gҪp;bU�ȓAK��{�ذ_Y0!R�+��)h��ȓb���@�OA|� �a��߿Y ����D�<��vFޅa�����E��<:��ȓ:�V�*`���q�(Y�BV;ht�����+�X���yP�ɝ�R�!�ȓ���X�o��}5�+�샅0��<�ȓ�l�������1�7N�n�D�ȓcC��k(�^N@�R%�ݺ_W���d�r�s���8���SC�>O
z��?�͘��;H޸��#G�w�i�ȓY�d��q���;�<B��ƙG��ȅ�<���{��f��1f�M��6��+�!��X���)��J�7d<��ȓT�H�"l˂a�X���Aѭ���ȓy�,��jS7/rL(v ZY`a�ȓ�A6�Z�-8xQ��J����S�? �J7��,]���6�єz.0<�P"Ol�Jc#R�s�����.9�4i�"O�����ܶJ�v�p��-?��@�"O�T͆I�v(�EO�/�HA2"Or�k�o0�%R�)�R��@"O���7n�=qЉ��+�'��d��"O(���2�扪ǩ�,��A�S"O`$��KF5BD�khд"���"O��3
��B�0lɠH=b�hd
&"O.�C�O�Xa�ɺ�.�!2��"O����d�	�����/�f)(��e"O��m��q��٘,�H�B�I0"O|�ȱ`��V�Ԍ��дn�����"OL���L�$,Q�L x ��"O:�X gWY����KG!l�:�;`"O������uFXm���p�,��"O�)�T�jp�c@�ȭ�z���'�<ɱ�E��4.
����U�9� �	�'qLA��)Q3T����?y���'i�xBBB��(����8ؚ� �'6v賣F�7�v�����4���j�'c�Ԛ���&[�V���Ȇ�-L���'cd��/�l�6�T��#�N@�	�'��hC�>Q\��C̓�|��	�'��1��"��q�2��;-`n�s�'��C�
4Bc0pj3ʉ�z"T�
�'�4���.O��qS�׈a�,��'c,��� V|��7�K���:�'� ��H0�^�Q�_1d��'��U�io�,�vK��f�6�[�'a�A��R�-{lܢ0e����h9�'o�Y�Ӏ�5eֹ�Kц"S><h
�'s��ca��Q$Y�"�S�U�<�h	�'f,Z#� f��9�*s&MX�'��-!W��f�䡢��A%wipɋ�'�P�2�N�;�����(�L���'�zL�@G�$-P0R�o��rZ���'�u�R�K�l6�����!k��Mj
�'!���n��"ᮁA`E��cو�*�'z��p�Iмu�� ���(�P�8�'E|��#/���������
*	�'?\3��MO6	� 	*儹��'"�PD�T!08�����\��;
�'|��Ar���#���MK�I�dt�
�'�.�3��E�T�<�5 ,G���		�'�.ġ��J�7��mse��2
\Q�'I:��d���$e s
ք7#\Dh	�'���P�u%�<��H�*ƶ]��'`\�5��T���j����4M:��'��UcwC<��q���#9���'O� �t@WJ�� ��HJ�L[�'m�5(�d�%Y�P��;G�v͑
�'�b���-��F����c��?b�
�'�dDaQ&	�I������7��*�'s<� %b��N �K6��_P�Q�'���"u$ 
^	��`H������'�2u�����]A�9p�8
����'�r=����.n�dy3fL	i�4�0
�'A����M� n�JU��c���8
�'�ɋU���0e���D(����	�'$� V`Ҥ$o4P�f\y��C	�'����r��#*�Y#en�	{�����'�b���JK��LM[@f )�L!	�'^X5bP�:*�5�dHשZۊl���� ���V������
���ڄ"O��c5-�L2�(�*E�"Ory3AC����M�!cp��j�"Od90�AW�R�|� ��Y+lri0�"O~�ʔ艆_I��Kf%��B���"O�p�w��d���&$�|?Ƅ��"OV��b$�}�,Q�#Ư)(�ɢ"Oʸ�w�&B5:���@	�i��"O��b� Oq���o�X���"O�؃�M�,O>t�@3�|��"O��[Coְ1qr�)���Q����"O:�"FG�xa��A�:����S"O�0J�͚�"�ƭ�g�ǲZ�t��"O�)�ٻ d�hqBK�+��4"O��r��)4��P T��}XH�j�"O\Qz���!K�x��&��2r]+�"O����OިVjV�z�'jYФP�"O4��a��4`���d�E�< �"O�-{EI젹�F�#	�-��"O腑6hB�Wj-���џ�XD�"O ���U�)�v,�D��n��a"O�aAU�]�pu�8�`���$�Q�"O�-2�&ٓq��
����2"O��/�O �!�Ԣ� �"O)+��� yڪ��!��.`���:�"O�`AE�8yCd�z��?P�"Od]��P_��`�Ǐ?<�0"OF�c�O��@S Y�_r�u"O8lv�\&�����JV��Q3�"O�e
u&��+��M"�Њ�"�P"O�ҕ��:7���d�˭syV!S"O @ċÒR��ʇ�]�#T����"O��3�A�0_���E�G<"]�H"O�Dzs�׫Y��q��7J�p��"O�=8�F��VےP�J�HN�u�1"OH��T!\��P��ʙ!-�x�T"OB�� !)&�*�
p焼q��i�"Oh�x��Pv���bB�D(J}�cq"Oȡ�A�%��!�2E�7mB��"O�	Ԋ�Y�z��c�Pr��u�
�'����1F"AZ�7�X�Dll�(
�'�@�U0X��k����9?�U�'^�d�"dR�Z�N�ٶ)��n���'ւ-�`e�Z
� v	G�U!8���'��j�|*z� U��+��'h��U��Z>ĉ�*�M�҈ �'��p�7�
�5:��q��:�%�
�'�rU
�j�K�� �2C8��	�'�* �I�
0�c0b�)���'��k���O�\�C��]1!�"�S	�'EjU�* �J}H6lZ�K��)�'4�q��H��%8B��eQ�(�|��
�'�8�P��/B6��F
��z��2�'��-�$P)��pc�,���	�'�n��`�1<*&�� �R#1b���'��pK�)���p�LJ�5Z��'��J���.��9�� <WH�'w�e��(BZ�@�0'&d�
�'��)���,!89��6Z-��'���ìUp�\}IQ)�S�x�S�'�Ƞ�q
/'I�@�V�eB�'����w�6E�֡�7IY��b�'��Prn�C�"xz���'6|���'�Fq�sL�;�JȫӍC�F��I�	���  �;#�T\����?W�ؑy�"O�5#7ȜI�MyqIG?1;>� 5"O�B���57(�!����N�V̊T"O4Ѩ�ʡ+�>��p�X�+pD�c"Oֱ˧�	#I0M��BLi��"Od�{p�YO�0�[�!S�l���� "Ozt��� $[Y3 ƗP�&�Р"OB�cK�5��y�u�ƥB�r�#�"O@ ����m%2�ϒ?�u�A"O0A��hI�[a:%P��"h�t H"O0��S�ץ�@��g�e��ykQ"O��0���/=��Kd`H���c"O�\CU��$6NpRv��('��"Oj�R�̊7^Ta�
�.N�����"O��CңA�d���(1��hr"O��h6��8Ͼ���<W�N�
"O�3*���R#��iw�y��"O͹6#9t4��b��0�`"O�Ł���n� y�T��� �@�"O�6��V��]#w���X�"O�a_�8��e1b�23�N�g"OΕk���aq^Q��bD�Z���	�"O�ds�L�c�|X "cE<$����6"O֬Ks��i3v`�4?�4�A"O�q�!��y��̉&���N�d��"Or�`��>�t����[���0�"O���eҲ*(��蕔/]qB"O��IR�Hb���G�͗t�e��"OB�'�#h	�ؖ*I��)Y�"O�-�t��
@6���1q
�m�t"OR"�!^�-B�����݁��0kt"O:T���[`�D�d��05��0"O^|��gU~1qM,I.��"O�T���^�� �ݜ9��� $"O9�Q$�fi��#5�RTf��"O�4�`J��`��Y �/U�}��t�"O�a ��~�b�  1T"Ob�)co�+):�Xkv�ߋ-�����"O����ʚ�`���*[1Ġh��"ORA)c�D!�(��,̀h�"O@��K��9������gL��Jd"O,��5A&/DT���1^T��"OF� ���y���B�匀;*~I��"Of�K�oȤ)Q��Dݱ5��$��"OڐhB�2V� �@"TlZ�5� "O�� ��з0�X��D��5uH�!��"O��X�dûi5� a��ז$��ii"O����ש�����Z="�h2�"OH��RA+ �8A���U��pj�"O�pAa�%PB0�n�s�Z�q"O����0,J�k��������"O8L�ƮD��a�&'A�b��"O:!a��6�l+��0R�NsQ"O^<���5t�4q���=)p�Y��"O�Xi`΄�ux91q��2g
��"O�:��"+����J�D.(�v"O�ɒ�^*d�*x�p��"6X�"ONS���t�����Ž((u@&"OJ�r��֨@h}���&;sLͫ3"O���\3Q�0`:��^+L��t��"O���
��l�{��,VJ(yc"O��)�)��T�l�6@4G\ "O*��nT�vx�1���+M�I`b"O�@�WΌF�Va�%��*0P�T��"O� �����2n��BF�	b:\m��"OdJ��V�xX���R	�35��0q"O��Q5L��@���{'�Ȉ�|��"Oa��P�(.R4�����;�"O�aJV5L�Ҩr��'Q:6�`�"O~Lá�I�P�:����*@ԉ�D"O4y�5�Ǐ���f曈y���+$"O`���
K+d*��A�'9l8���"O`�s
��;F��a � R=R7㇍?�����	�)���?�E'J�4�.A�A擿V|+U&p}b)�������z��G�`�ꁮ-TMxa�%���8V
U�?��*� l0s��j��	�e���5�$�2Sw������h��M�I"�m�2�D�x���'�D�I���O企���$6�5��:d�pM8(Oڢ=E�� W�
S>�1��QLD@��?����S�;YN-I��N
$�����)<~&�=)���h���󪉊2Y�}�3��$�⟴ړ���?��?�(�P��)a���4@��aԌ,�O�\��I��ª�O�αȤC�R8��P,)!R)s`�i���Jph�G����OQ>0�X�r�Q��F�^��@L�^�R|�Ihc��O��֧���a����?H�:h�v��[�!]�{Y���'Y�) O�G>�R�ž���U�^�u��i�b�ܯ��$�z�ԡ�	��0|B��Y�^��)�@��GF�i�P��J?�dl�K�8:"o�����]�ޥ 6�`�ݺf�WF ���b"r�0�}��)sc��B�gC�k�p ���[���8'�)�'�u�\�B��pY�ė��ְzvB��hO����L�m����5m�~7��h����
"�OZ�=�����GI#y+r䪕�S,g�Bs�|��)��=p�G�4Y�=�ՋQj��ʓ����Z�\�b��eX�R�x�ӤB0�A�U
V� X�O�?UB��^�<"�XqanT��̸�#���'�| �}�q.�L?Yco%,�̰�d�U�cr��(�52�T�'���ٯO�}�I~;�l��ˏv
x�Ҿ;{F}�C��@�ў8y�f־N_0�i_2��S�[�DX!�������F�!B�@�3�I*�C�(��e)פ
���*�Ƕv��C�	<R��Y26G�W:��i>u��C�	;�B�
�'��Վ�
MY�C�ɑ�^ ��˽km�5ǃ�j��C�I��݁��S$*�0�C�ٮ%&�C�	0C� 5�堌G[n� '�A��C䉈~��m) �P�H�:�Iր�V�C�ɫF�ީ���B3J)\����oDrC�I�YAʈ0rc\L�.-Zu�Z��pC䉋1�r�AI�n�J��e�EJ`B䉆
���1vOM"g�.�;������C��G(F���'� �&�y�-H�C�/Φ2��Z4&PIR�n��C��� �铔W��0p}��C�	�V�20��1oưy"��2��C�	�7A�ȋ%HH @z�L녭M h��C�	�#J X�%̐ .���fg��gxC䉄Y7䭋U*��uz�P���7C� Z�}B �H�:�:c�.s�B�I?V]��8�"T�)%Ě�r"C䉸8/�;��f\��ġ�9�"C䉾J��LZ�I��.|�A�L-��B��:\����B�M���Hq�"G��B�I�RĬ���mW�/lA�	'(B�(>_�Ds%��o5TA�����xs�C�1��a�qMC;}� ��-�e#lC�	�a��x&�ƿ�НCJR;C�	�	t����ƀ>r�EPA!C��B�ɮq(us��(��Q�%�k��B�)� @��qiC6=!B���Q�	��Y��"O�Y#�@��<tk"F�4���"O���dG~] R�+�:�X�9�"O�M�"���?bp|��V4;��i�"O\�j!#�)��&�  tI"�"O �W H1A�J��$V�Hdބs"O��S���!46&!G*�>-,x�%"OBl1�����B���cPu""O�}s%F�k�4hё�̀O�\�2"O��f�G)xΦ�#f�X�I�Ƽ�"Oj����̹udh�@�� �Lp�T"O��d�I�:a<���؉B��)p"O�4����*0�feP��L�o^y��"O�<#��ڈ7����D��:k�0��"Ov�z �%dP�8�'T6���"O.���˟�wX�Eð���x=΄��"O�Q�!,���պ�\�u`���"ON4��mw��(��
�n���0"O�C.�R P�h׈�N�}��"O�Ț�@N�?Y��W&��̚s"O.L@�[�� + %�#4ˀ��@"O�pd�ؼ�bť�5[�e:d"O����͔/O�^���c	
�α�g"O���֡� "�t�S5"�'� "O�Y�1��!W��B $��"]d��"O0ia�NA�-��yX�HK���@�!��E�*��P��Q>��?@�!�$L64�6�"��f��A�G�t�!�O�#�N�" BC�+�Иy��!�$�<P���b	~�,���)!�^8~��&K"d����aP�"$!���1R��A���(�V�ӄ�çG!򤐐&�u��O��:��t���24!�D_��9��+��`���  +!�d�1B�X�@DW�R�F8��d� �!��
�r)���ɳW��Psd��!�2"}dy0����(����S-R#�!�dG$m5��;�*��,m���Y�!�ċd�Tp#Db�7lZڵa���X!���g0�X%�]5:�i��/��X�!��O�,�(��� L�y�A��$�!��G�-��m�N}T�І��$2!!����0��B�Ox�\y5 %bb!�Ju:�4%�#c�p�a�Q�L!�D	f�<%0�V;!O�����)g!�df��Ha�ID�����B*Gf!�ӵ1Z��z��2|�UG��"`8!�$²x�p1�n�k�ԀU�@$jJ!��G��A���9
0�to�t<!�$M3aMpDp�P4qHQ��P &-!�$P!`$
4�����j�6�#�� �!�$�<_
d1x��H :�ʰ��}�!�dĕ,X��9C�C D8-Y��͐8!�$�dF6��Vj�}X�Z���� !��[=�V�4�ј$Tl�sƯ���!�D"I7��3�%s�(��.�	�!�,��!AI�7�+J��9�(�ȓ+U�A�&�J*D���,�74VjՆ�[�J=�4���g@�&)	�Z����ȓW��R� K9��A�PᅸP��ȓ$p�L{BL^R���ɀ�ߴvR�$��
b�
W��1e��qq�Q�/80��"z$�3`��@��Eq�"�V�ȓ~4"�:��S+	dP�A������S�? �m��J�r�>��"�b/�Ѩ7"O0[��^�M�L�Y� �'L�HA�"O�4�B*�<��U&_�4�T��g"O�(���ݘ�R �Qe/z��Yiq"OI��ÿt� r���*�h "Oj��[�F`d�U	Уw����"OP��Ҏі>d�x���Į<����P"O����. �90��@���-}T� "OF�cES���cF��ؾ�9�"O�<���^�"���@�ܠ��up"O4%��Q<J�DZ��� }����"O0A�'^,�����-S?p�6�"OB9�U�7�u�m�)F�=P�"O�Z��Ko`�܈ƌ�|v["O��BI޿#�PpÆk�v�T`�"O��fE
�>��|`Giق]��A��"O����)F<����n�4��2 "O�M҄�$l&�@+.F�o�"O��s��^��Y`�oO�J�0��"O4ĈäMs�]���ȝ}`��"OR4HAi��(��,� H��"O�q�-7ȐL!@�8S�:$ZC"O�Q�B�M�1Xp�UI�/�X�*�"O�=8%�> `a��]m��SC"O��`t	�?��;Qm" ���	�"O��B,,_J�T헸+��(�!"O~�Kcԫg���3�Mȩ�����"O|��	 �-�����A��j���"O�!��i/�����D+[�0�"OB�I��2PAx�)s������!"O0�X��o�tQ3!�$��=	�"O8�!�ӢZ�ެ@�.�i��)�"O�S�o�[(�L22c�d3$)�"O�,��H͋3@ ��@��kOR�S�"O)p �Ѳ%�JUy���T`��J@"O�y1�H��d^��q���+[|�3�"OP!(�G��H�ed@*SW�4�"Oj\AČ�k�(|���,}a4Pp"Op}Jsi��f�^	9��^���D�v"O��8�-Ƒ-<`tyt�N>\��"O��QVjӯ)�b��ġAdЙ��"O��32�ø��(F������H�"O��D���J�Pru.ݯL�D�X�"O�2@-�[�l�(Qn�-�b�C@"O��� �V[rA;Ӫ�?RkJdX�"O�U��B�`�pM���ٰ V�`�"O,p0���zE���͗ P����"O��;rl[yUZq`&Τ<j���"OB@��"V�|}�qHFG��jH��"OZ��Ѭ�r�N�â�&2��1"O�p ���C��9[��V�Z�%�A"O��YD�ǽ���bP��af*2�"O�YRK�2h鸉B'��":��A��"O�⥂�KŎy�e�T�D=�&"OV5�S�!4�X���-c��L�""O���j����I��Dݤ1��h�5"O@���� �ʔ:�$� ĺ� S"O��v˒,@�����U�E��Q6"Ob<���@�%:�5��K�e��+@"OF�����	R.&�X�h��kƴ���"O<���̎T�^�%�1�y���3D��2���> D5:J�05�b,���1D��У�6 ��&NQ�e&n(�#-D���5�M?t<��F`�%v� =�B�,D�� :��fJ��ʀ�@�(��!q�"O�\�'o-�:lS��N���+6"O0�⋗]��Ys��M�vQK"O�y��xh�[6uM�a����z�<QS�˟0n�S@'�,��r0�S[�<�e(� e�F��&T�apq�U�<���ψ�V�S7!&C�]�T �i�<���T�H�"�_������f�JC�ɶ0TI��HʛQ��`
E�È2�C�	BC��	�C� V�`�e�#	��C�	����Ō�3����!T
u�C䉯#�b�
�5?������={prC��+�q�B5e�^�ӕʃ��tB��:K3�8�V�њD1jU3%+��FB�ɔQ�p��I�)+�^��P��R�`C�I�x+"�
ո?��qꅭ�i��C�I�h�[�'2v�x���E^�C䉊�4eX/�J�(c/��m)�C�	�8&P�{'R*D,��cEL.��C�IG�LE�	�dْ��=��C�	
n�4�����o��K�)/�B�ɂ�N%`rj[>^�`�f���2�|C�ɭ��)@�Ŵt6d�KүB=�FC��0'���I� |�Y`!Hܤ:.fB�I^3��p�cT�lXDS�)E�:B�ɫS�n�q�+�j0
X(R&C�kx�B��#ҭ�0,�cX�!�� �D��B��b3���Г f����*S��B�ɣ@V����I� $;�)�Rg�B剉[���6��M��2V��� �!�K���e3`� �� E�!�ē-u.HA)ɠRn��;��ʥ<�!�dM����I���#7|E����M�!��B픸,E;�����A.�!��7mF~@��g�,,�8��Z�!�d	3?��J���K\(	e<A1�'}D��r년/�2��'�4U��qh�'� ��"�Qs.l����X��0�'�z��  ���       �  m   �+  �6  �A  �J  �V  �a  �g  n  it  �z  �  3�  u�  ��  ��  =�  ��  Ĭ  �  I�  ��  ��  |�  �  ��  �  ��  �  ��  ��  Z - s � �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��	h�I{n��Cv�ݨat�����R�p�<9a#ړ�y��P�k}dț�`������
��$"�S�O)~lYw��Z�>d���٦D;�|S�'*>*C�1��Y�w�J25��PK�'��b��8��2�Y=&�HQ�'<�u
cC�b�`�:!-ǅn�>yi	�'x��h��3
�T�(�U�e�jp��'<��%p�D`�ц�,�R S�'���"-�%@�
-� ��$^( ��'7������>T1㯕�"
�'��!hd��
N�*�朴f)굘	�'�~|����">	5o ����'��Y���8Q3�a;���4�8�Ó5��	G�	;F&�S�;�й��J)o���d:ғBL<�A�A�T�f�#Ё�##�����~��I<H�t��
��V�(��C:]��M��IG�w$�眧,��7ٿIJ~<��7��8�N]�76m;���:� 5G{��'����ċM� �±�ϧX�{�'i l�R䓩,�J�4H�+[���
�'G���%*|�F�2�N���U"<|Oc�D���ȐN�T��v�X�Vq�
?D�`���ώ"��x��ͩj�pӢE=D��襫>���M7L|I��&}2�'����cLM|uH���H՚$�$Z������t�6]+��P��@�B�)~!�D�J�4����1�hPD#ݣ[�qO���ȟ�u��
�CKJ��`��>1��I7�'� {'�5���t(A\X{e!6D�L('��.>���'�]"4��1�(D�� X����ǺE	Q-B
_�F�"�"OLU �"��/�4i�-���~����'��LXj�(Al�x�� �&�j��!<D��1�#P�i��ܚ��3�r��i4}�)�S�6<���>��H	�`E�7�C�ɻ]}N�����1�����-s� �' ��	Iܓ��'m�  ��b9���CB�%4��U��'�<]�cOU�	J=�Ҍ��R�Ty��"O�\�0�C7���ɠ�NG>�
7��|��w쓋u��I�,�a�P�(U��-���P�j�!�
 �����ŶI4tB��U��'j4�R/OF�<�Ӻ�DR7&n	}�H~.���������V0
�lh6���x����'Uў"}�1�RB�ȌѦNF8J@�5
B�U���OVm��8�|��R��6pʩ��'i�,I娌�m/�Q���f�$�Ǔ#>�"<�&	�Q����	�<����#�n�<�r�4#�|ɵ���A<�0�B�b�<���Ǩ^DT1�Z&WX�]R%G�`�<���	�Zz.$Pc��&`DJ+HZ�'�xr��@�n�hg�I'��=����y�lH�V@~�cS�Z�.�e[�B�k��B�	�6���s�BҒX5��¡Ο$���Dg�ȩb�\�ɔ�:�Zg�C�/��(�`Ͽb#^C�	(
�2];����t9,�Q,R#<���?1�2%�+O�F�X�Ȼ���!K3O�#=��ңO, �8��(g����HO��}�xHJ�i6ꆼou�yB���\�R%����ui���_L�����h��g<	� W�&1:��f��.�C��l���O�%�:��':*�qvɁwPry��1D� �q-���bU� �j`Y�we9��MC
ç&�M�ፂ5f�ԭ#`F��Q|4��ȓGQ+6��i���a��D�H|��^�l yScо0�EJ��� aJ���ȓN�yY &<�Rr,��Ϯ��ȓ;�x�Y�Ea����A��=��IH~��6.DUKV��*L��B�G��y"��
�h� /B�6>�	J�L
�(O`�=�OK~-R�Z$ǦaYFJ]'!�R1*	�'H$�0
��y��କ�N��u���(�S��?yǦ��K@�O؋��
� �D�<)��ۭ%���ҏ#�l�%�؟�Yr�'�0ٷ��x�8�1&�S�{"��Y���TI��<��f��f�f��r�ԟ��q�l�e�<�@�̸G�dzEʚ"�,����Z�'ڨF{�O]B�ұGȄS�.����3	d�9K
�'�N�c�C;�8\��V�k��r�'ў"~'�8\t-P�╎ �!;tGbh<����m�Tm��ŀq��l%	#��$�>�ۓj�@�s���֥P5K�&Ntz��<I���IŽ(�~h;lV*=n�Ѩ�c!�D�6`v�9�e��$*)
��w�ϼjZ���D{��\�gOܿD�V�I�OS+v�x`��'�'�*iy� -$c����H�.0<�H� D{��4�f61�3/�%!�E�yM�W�hr�0y ���M��yrf�g$*��n�\{�EDo���'�	o��~B��%B`@�����"WUdd�b�y���#X,���M. �8��K��~B�i��IH�)�,O����El�j`"Ƒp�8�pq"O�ͱ@��_�Rݺ�i��6�Zp��>�����S�O��Y��bB-G��EsB̋�u!�I9橘Bk�#M���
gÜ�!�� �BE
�T�&�*�IT�3�ȑ��|��)�F�Vx�`��5�(QH����6��@p�'ZfL�v
Ϫ.��Q1#F�#�`q�	ד��'�(0��!	nR�������6�B���)��G�$���� �۟��1[ ���'Nўb>�X��΍g�}[�!��^ ��Q�#>��v���")}�5�W��]"��j�DJF�B䉺y��� E-�*7!�=s#ʓ|����0�S��8O�Di-O��	7�
Y���ၒ�/9��"O�Y��.��/�l�+�ғOɨic��s�����pCvI���X������'<�{��|d3�،�����^��$��BAָ��}�����	
 �))� M�kZ��jÄ�-�^B�ɔ@�b���!1�t�A�&�VB�	+u�d��J�!%�^!�� �FB�	⦩���3V{�-�6�N5-sI&� D����kКDHX�(O�V%& )�>�c���'C�ċ0G�0vܶ���m\CaPT���s�=C�E �o
�m�L���fK��@$Ey"�'�p�BbCU	����j:0�HQ�}��)�IA�f��q���Đ�^���E�yo!�7Q1�s�u=H�9���bd��$�=_��z��]�K�J�+BÚ-l�B�	�=��	���B�z�^� �`�@^���J>��������/,l�G��U�VxE�B��y��8km�	U�S
Q��������y��Vq\���J9K��m�%I��p=��}��	f�*� T�Ռ;���@L�y������5/�=�(j+ƅ�y"̋�y�X��Cʒ�4�,�U���yr̉!<��i�  �-&���J�#�"�y��J�ub��\�F< �Q��F��p=9�}�H^�dK>���M�>��)B���'�(�GyR������X������iZ"`��(+D�����8+90����*-��mÔ�*D��J�
�;(`!B��ݺ<�,H��*D�ag O8��k�"�&8�U1��)D�ɔ�X� �td��j�0W"@�[��&D���C^�[K,(���5�y�G/D��ȇ�K>-0\@xpCّ��غ�/D�LxsjFId����K����z�H.D��jJ= �����E&#�!�-D� yEfׅtJ����!���I�,D�����G��Zԛ A6Җ��P�)D�ɗ��,0�*��]�1P��b�&D��y̆&�(8*�!�(ژ䰃�0D�D�㩉�j2bQ�"N�S�v�kp -D��ꇨԖ\��YX��W�(D6\B�,D�pȓ�[+~F��a W6NSր@�I8D�D�B/6|ˇe�1�0É6D��p��_D�\�I���8)��7D�Hl
b\�8�K�����y�
5D���w$�	���zSi
�?�d��&1D�����H��Bւ�%0�VH���:D��
DI�r�� ��C�����/6D��bb�y��	�d�� ~}����3D��� �ڕ+s�D�������XH �1D�0#�,O?)k�5S�W)Z�h��2D�h0�"զ/��SPi�+gr�U[�#D�X��L�*$�r@��!ZHE��$D��[q��+G&e�w�P�[/@!�N7D���0��9�$HXWIB�g�,�j�4D� �eM��mWXe��,@$w'B��&�6D���T�U=yH�=˦#2cwBxI�0D�� ��p5�do�Pyt�Z�A"T�A"O���� /Mz|�f�\�)] �"O����A�����wɟ7?
�Y'"OV����;�@�PiH&6ҜXI#"Oܽ�D!)Jv�C��	Q�uX��'�r�'���'%B�'0��'���'��d8�G=M>��3�#� C2lj��'���'R�'��'*R�'!2�'�ȱ��BO!|��Ez� �lsw�'&B�'%��'���'���' �'2�R`�KuPx+��GZ @��p�'���'
��'a��'^��'(��'��е��r¡�w��W��s��'���'-b�'"�'J��'1�'�P@�
� S+�}	w��rE+H��?i��?����?���?I���?!���?u�޽W��u���ǘu�ժ�G\��?a���?����?I��?A��?���?D�*\��uڔ��,E_��Y��9�?A���?���?���?���?���?��!��f}�A�Ό^�,$�������'���'b�'�"�'%2�'���V�o�@=@A��f��1R2�'�2�'R�'�"�'��'XҨ�^֖%P���T
Rp*��0��'��'J��'�2�'<R�'r�ǥ5^���jT�c��;"�ߛ�'���'WR�'D��'���'�D 3@�t�3x���֨ C��'UZ~�F�'D��'�2�w���D�O�\���+_�xbj�q&rHF�Uy��'�)�3?���i�����[9*�pz6��ԲTA�jI����U�?��<I��iWV  �F�����x�L֫-�"��rIe����\�b�z���Dp�Ǯ73n!��~RqD[�	�h����EF��2c��Q̓�?9+O$�}Rf̌:w!�؈�M��z���G�F��-D	��'��0�oz�i�����n�b��^�J�(ЊE���MS��i���>�|zd����͓/���#k�c_��B7�ֹ7)�|�$�]�U�6w5ȝs��4�����>r[X�Щ@_��,c��K��<�J>Q#��1���<�q��>w��h��	&n$npr�O�2��'52��&�P��<O6�lƖA�g�viԨCU��.j ��'��(+W�D�~S0DA����ŭBU< @��'b�}�s�S�:c�!'!��(3��a0V���'2��9Ot��C惪N�l�`/ŗN�9�9O�n�!2�� ؛��4��3S`ٔmv�X�h����#v8OHmZ��M���rVr-B�a~�C�R=�9���؍"b���j؎Z��2�Ji+��W���b))F��X�t�)��6�F�Nf�A0>a�ѡZ�o0�'Y>qG����l�d��cBnh5�4Ó�+"��a���&#��<���/R\�� s��}�z��� �ݣ��]/��1�G�֌}�^�� �1 ��
s�D}�^V��01Z��ةč�2N���+&8�L3��<G��h���%�`��D�/uP����C�xA԰Y�
=
`|,�F�6S�XT(V��c��#��(:�`aЈ�����df�"i�nes �Y�?`ݣ��z�����O`�D� U�'H�M��ɏ�%���#t�@'L��`X�4��D��Dp��f���,e�\�!¢v
|�b��0pś6�F�P�86-�O��D�O����G�I��)�k�t�vyD�G�8��qs�\�M[5cث�����y��'�E{wIۀQ��a��� �����r����<��%
���<���~��	@J���gw�L"�f<A��b�� b܃�ħ�?����?)�Bφ3��ġ�S8��r7f�*��F�'`<1�&m;���O��D>��Ʈ�@p�qBp����I�tലaZ���u�9�Iʟ��	ڟ��'L�چ�	��aS�*
%@��$S󨅜vp�b�<�	T�	eyr�G�2���c����x	�H�"��,��yR�'��'	��'6�0s��'���+$ʇx(8�LE<p��ӳ	`�L�D�O@�,�d�OB�$X�?r��#��i�:�QЬ��wR�q#�ȩ�(1 �O��D�O~���<��*�.Nm�Ol�6���16D��g$���J��E�]�����`��{y�T-��'GHÇ��H�� ���8#O�}+۴�?I���?�6P(I.��������;l����[��e���	�\�'���'�0A��h�������@6�d�Cf��Rq ��.�A��V��1����M��P?-���?is�O��3�憃}�"�i�k]��S�iG剞��"<�~��CR�Cw�K.a؞<�Ba�Ϧ�"qG�ş��Ry��O�Sy�$¶3�����
J�	���[�c��6H?e���������R�²�:cMM=@�y�KB�M����?��y�ȐH��i���'�2�'�ZwD��1�$��ud��	#�S�=ꪩ8�4�?9*O8YQf<O��֟��Iٟ�1���B�&�*G`K>SR���a���M��eפ�	P�i���'K��'J�'�~�#��D�ru�8����<���ň��d�O��$�O�D�O��'r�6���CJ�9+∉��C����ɵb?�&�'���'R�~�*O ��- �έ�E�<T�d�9C�U�%�J�=O��d�O.���O��$�|Mńp��fn�*��{���d�p��BM�Y�$7��Oj���Ov��O4ʓ�?����|�1(9�������YF �i>~)n��,���L������\�I�t�|�۴�?��N��yPA����UT��&���׷iKr�'�"[�(�I����쟈�R��`Hf���JT$�!��2I��eoZ֟���ʟ|���q�Y��4�?���?��'72�"��� ������m؞���i��_�h�I�Sr��S�������t�? �mH�(�F��K�K������iH��'���-u�|�d�O�d��@���Ol9�K�C?jG*��]9�0�"a}B�'�RL�#�'6T��T�)^*D@֙(BA�����'�ʈ-"�֋��.6��O��d�O��)�*�$�O������b�`⎡���3L�����iϮ2�'��Y��p�ȟ�q�B\9b��T14-��EӢq�5��M���?��XL,M���i���'��'�Zwf��#g�U�p�x�#K�?Re(ߴ�?���0��tY��<�O��\�M��z� �p҆�(m�J-�U���@$��"���?qUiN#v��'q��'�bŮ~r�'m�e�3h�?������[�Dr�43��p�����<i+O@�i�O���O ��Ң�lh��νB��	q�G>B C�Y����ş���۟xˬ����?�0'Еf�u�!B�(��ѵ,߃x 8@�<��?Q���?9�[?X��0�i�:X��Ν){�0��V*D1�@���w�2��O����O��ļ<)��.0:�������4��!x�H��1���^Q}�$9S"�'�r�'!"�|����O�p@��E :B���,��k@��3��	�9��Ɵ���fy��'j��j�O���'��0�a[�0���w�=)��y`���@7B�'���'�����{�b���O��D��lG��`P
��ć����
���U��~y��'u��(�O�ɧ��4(�ƈ*U
U�V���V�?=p�]l�؟��ɱ,���ߴ�?Q���?Y�'���N����$�E)`}�D�i9O�>�S�_��ɲo��}��hy�C�-����~R��/?`x���ҟ5z��Ce���uQ�ʊ��M#���?Y���R���?��?���%hXp�[+Tv�s��[���ϕ1��|�O��O�R�p������~���y���$��7��O"���OHa8�����������I��i�%�Ԅ�	�$B��L�sV�y׫nӈ�8��`x����<�O����'��3b�U*�f� ,ܚ<�Ӯ��B�7M�O8��ↄӦ�������Iߟ�p��(�I�vA�8�ɋ4I��h����ժ�u�(�'���'���'�b�'U��G�0(��P��&	��+Aaa��7��O��D�O���q��S�����B�X�c�e�>�ޑ�83ն9�gk���Iٟ�	۟��I_yB���6��S5B��(Ɍ4#�,��v!ؑR����?��������7L��I�Z.��iS��ZJj4��oTp���?���?�+OB�2H�M�S�m�@�5�"�p4*��I�r�C�4�?�K>1/O�C�ă-�nHr�ɰO���Z�hK!���'|�Y�����,�ħ�?i�'=�vͻ֮�|찈33�E.C~ (�@�xrV���9�S�t  �T���r�M3 ?\l�c ��M�(O`a��Sݦ��X�$ퟨ��'*@h���
��ĭp�R�����ʦm�'Z�]Џ��)��u��p�B�Üo� � ��E�B��v�/u�.6m�O���O��)E�	����T�0~�%�u��ŏ�M3f��E������S�s��Q�@�f2�CE)˖	��<l������Ɵ� l�-���?���~R����6a�VȎ�Z�B ��FF��'��ɉy�'���'�
T�%H�w[�%��j֔r���k��w����.L��&����%��؈D���l��f�<�@ф^��X�g%��<���?����d��0+|���T�Qb,2��ڶc"nՓ�aG�������x�ty�(�&B�Vlp��\NJ�Ш��X�=S��j�y��'H��'��I
ON��*�Oւ����
{tG�W�ZYđ�OP���Ob�ORʓ_^��'��@�b��?@�N��L�R��Љ�O����Oj���<ـMB�6҉O��Q*�d5$LA�+R�e$���4cm�B��"�D�<�!��V�ef��;tÉ~4a���̔62��m��x��fy"�('������ޕcFH��fy�:��B�uD�d�5��Q�IEy�	�O��%W
���@��X:��IR/J�C]�7ͪ<�ǩ�.R����~Z�������0�h ��0R�}Sj����o��ʓ_��dGx�����+8 8�b�@ֳkaN�@�Mk�b�*&o���'7��'	�D�-�$�O��儊�L�H@�ǩPHxLȂ��֦���&4�S�O�B@ΗtX����	D�C�4��L+I�z6��O2���Ot��CJ�O��?��'��Eq�oV����s���$PEЌ}��'���'	ō�y�:dC��Q`�ڔkFNQ� ,7��O�ykgυ[쓿?qH>�1X���)��|��I��&,���'�\t��y"�'�R�'T�	�]^�E��[:F��⊒
b�rx�(Y��ē�?!���?A/OPʓp�`� ����d���X���!�?����?����?)����<<V�lz����N��zCH��>��ā$��O����<�(O�T��Z?��Nٞb
��{��;��p����>����?a��������5&>�S�"X�v�HreL�H��Ho���M���䓛��ҨRB�O��ȑ��=�.�s���B�v@*R�iR�'剋+0D�O|2��2^w�}3�!�<.�J���H̵�H�V�*�<�!�f���)��'G4�r&��G��apw޳%C��T��3U���MS0T?�	�?M;�OVI��!: �-��[h�`!��iC�"�."<�~�gEQ�?{�<��H)Ȑ��!�ڦ�˶��<�M����?������x��'�� ���3 ���
*F��]hT�h��A��)§�?�C� fɈD�B��P)���Rn���i�B�'��G	$�zO���O����>�H�V�CzR�� �0��b���V�!��Ο������#���-�uEmSz�.���h��Y�6m�O@,K&le�ퟀ��N�i���-P��pq�e�t�=a�b�>���{̓�?��?�(OJEG�^,0�P"Fi[�C�&)UKѲ�~�&�X��|$�\�'�y�%J��bp�#� o��uY����'���'�\�@��������B����G/�/:��<ʢ,�����O|��5�$�<i`jCO}�+	bqp�`�,	I���da�����OL���O"�4G�9�����x��� U(G	-^��$	؆7M�OJ�O�˓!=��>��ޔ
���z5�	����y@E�)�	��8�'�⡹�*���Ov��ڔA2VU+vm��=������k���%���'��j��T?�@��4vb�C�'�ke�(k�jӊ�0`���i۠ꧻ?��'S��1-�RX�1�R-U���؁$ܡ	`�7M�<�HL���υֆ2	^�+�O�("ntxh���$�M�CB[ƛ��'"�'��D�8���2Ly�G�p͔���ϙ�.�! �4j�\�Fx��)�Oz�j2��L�(�#��#��e����Ǧa�Iԟ���	,��t�}b�'��d�
=a@5:�KP�5]��As�9	�On��q�D�OV��O��a��1|�DZ�q��CáW����	�#AD`��}��'8ɧ5f�ǳr�V��W"H.2�-ґ���^Q41O��D�OX�D�<YD�F	R�8��F�7XF]R�BI+ox�M��x��'^b�|�X��	e�د)�-&�8F*4
��H�6��c�����t��by�.9e�擥hN1r�R~��lʲ�U�c����?a������$�-#����W�l�ѓ�C.j���H�X�Xꓭ?����?q.Ozp�\4l�
�ZQ��i	���aF���T¦!�Ih�iyr�E&��'�MQ��[�b{n����8I`��4�?����_�g�v�$>����?�Q��S�v�c�_��A�a�=����DǇ2���'c�R<`�ƂF��ly��B�C(XlJy2A�o��6͉E�D�'��$!,?$ ��*�*Hq�����rAa�ئ%�'�^qc�������<���H�(I�/��J��F�]��$7��O����O �)Ad�	� p5���6�,ŀ���6y�X�1椘��M���x�����$DI\Q���S�7L��R�;4�T�m��|�I�,z����ē�?Y��~"i� 	��*�I�rv�4Jц���'xP�I�y��'-��'�$��Ee?}�y�f�g�1sf�dӮ��0HL&�T�	�&�֘n�t��*�Mu�5Y����.�`����<���?�����־|���R��K"�|�9�MUTxR*�n�	���Id�I|yb�P&"�� �$� sh�þĄ��'G̓�?9��?)OP=q�S�|����c��`���Sz���b�f}��'��|�T�[4&�>i��� j�����>A�0����m}��'X��'��	tZ��O|
œ�lQ��3w

��r�Z bS�T���'��S���I�h@�m-�',���Ò�	l�DX�L��	Pt�۴�?Q���Ŷj���&>��I�?�5G[3
8�X�I�vat��7��Mc.O$���O���s�?�nzŅ���ɾA�T�$$yG��h�4��D�
J���oZ�����O��)�|~¢2���P�IZ+2��8Ѓ��MK��?�4������L<� n���H]�P�_� �Y���Ǧ�Un�M����?��"w�xB�'�$t*r#P�R��k�W7ƴ1ǯaӂ��a8�i>c���I�@{쐖��&��Q���3F�L�ߴ�?���?Y��E�5�O�����u!�s"���#b�R��TJ5�;�I8Dc���	۟����(&<,x#�C6P̸�R��
4r����4�?�5�: W�'
��'Pɧ5���=>�>�q�&llQ�� ����\�qC�<����?yJ~����
k\��/��A���R�nup�x��'��|��'��l�`,-�CAA@�p�F�X洡C��'<�����	ٟ��'h;� {>�ہEܪu%<x�@�[xx��>��?�H>���?Qrb�?�"�3z�b�j���$���@�L�*�	����Ȕ'��P� 
?�IޡlV���ԯ��G������/M��l��t'�����$�Rj?�	$3�0S«��@ܘ豐�+@�$6�O����<�i��mV�O=B�O#�P�  �����12�	�yZ��C�:�D�O��d�9|����(� bV�}�(��E�'�:�oZEyR!T�b6-Z}�$�'q��B&?��F�(R�R�(TJ	VղT@b�Ӧ��	ʟlбOs�t&�D�}*�lл*.PQc��\��/V̦cc���M#���?����E�x�'�޹93h�G�����Xo�ƙ�5��
�*�?O
���>��I�-qp�$��a��l#�ݼY����4�?9���?�C�i��'�b�'����^��ԛ��*A���%�<xۛ��|Ҫ��yʟ��Or��W(;4@�PC�EǺi:2���CZ��l�ȟ8i�%^��ē�?y�����{�c]�� �I!�����J}�AҋO{RX���I͟�	ayr�,� ��Q@	�B��������'@���C"By��'Hb�'��'Ir�'wr h�JT�v?.(�i��xNdq� L��S����ɟ��	OyB�J�
�
�7JDu��ɞ*8x� B����7��?�����?���,�q���&�����(��R��Y��Y�T��p[5_��������jy��ۊ9x�n%���1X~�˔�,a����
�����D�Iԟ��I�BaD�Ix�dL}V4���-��p"��:���'%�U�زck�;�ħ�?��'}�py���
4�(��kÔU$�a�x��'�"� <."�|���K#c�$>nx|��.��f}��@Vπ�A��c�'����U@ǑX��ϸ'��Q���`h@Q��ӻi9 }�'��p��ˉHc����
'�(��O+@��lP�^�t� dc�o58A顇M�����ZnH���nP���^��=�D�۵QF�xq��2K-H���ՆF�-�䇌S��� �r�8����޿x*T����V��0�zk��s��0ٴHzG�G=��IHT�Y?%,4�BM�Oh�d�O��D�к���?!d�γ�d��bG5_n�\�bb�u�b�K�Xы�`�'G>�g�'��%�%iV2T�7�e%0)��FQ�\x�4:֤�>T��y�$�����#��v�m���`~B��[F�;��С=�����=�~B�ܙ�?���hO�˓T󆨡v@ 'H7m��/5J��� r�Q��׵8��9@'I7wo��;��i>��IZy�E�{@7M��k�J=� ��
$��ע�����O�d�O�12h�O��dl>����:��w��# f�q� ��K�8���a��(�3b�`\�D���Q�~�@��@�<�؍СI�9 ��Ez��M�9��l�Ю�۰(z��nN�80*Jܓ$m���ʟ���A��8����5���@#'�w�'�џ��d�O-��&,էN�Ѫ��7D�@�4�',�&�TF�,D	2�v����4�?*O��OUL���'�Shr���ʛ����xH ��R5�ԇ��X�I՟@	�9x(8����<3��@�S��g�n}���0Y&rMR=ɀ%ݓ�(Or�h���~pU�b%U�F#�=��
~
��Č�ؔK!�V�p�d��tT�(ON9Q��'��IT�I�A�+�?݀�b���s��D0�OV���A�B�<���L�uT�B��'&OVq�R�#�,т",ޥ	f�Y�6Oj��Q������Ob��x��'���'*IpЊ
1Ě� d���.�lPf��?�h�Q�
����|*����T]��E�9,�<!����f�ԍ�Ph�9ZXR<��MK���O.��j�<B�Pـ dTtv�Y���?�J�D�OR��?�D���]mr��숓�9��"M,����?�	��L�(��H��!23J�/ĺDDxj'�S�4d�:�.#�� }��@��G��'0��S������'��'aם�����w��¶)��]�:<����:(򲉮�J��QrC�Y�/ ��������dk�|�'��@q�o\z|�8%�;$�iuɁ��e��
 &0�ȀF���/ʓJx@Z
.K��8��Y�r<�բ��w3ҠP���?9����,O��$�<	�b��ݫ�!����������hO?�� 8���c�V�5Pv!�ڕ��I۴xh�&�|�O6��W�x��)ا�M�d�(O�ҝP���#V4�"RFN��?����?��:����?I�Og�%�s'�X-F�[���Vr ��Xml�ʰd��N�D�MyɆ቏*�윸e�>�X!TĕUb��a��%��e�X
w �YF�#O" �'JV6�	�v6B���$�)��b�T�>ԢIl�K��c�>�	@��[��ݘ��0aCR�A�C�D���C��En�`��K�:)���I ��D�<�@d������'�B_>�#���8��P"
�,��4ᎿB��H��ʟ���`f(TJG�ô+_�8����M[+�8�ڰk?hn䝳B#�]��q1�	�%���m��R2-�a$EⓉ[|��AAV)f`� $qa��<7�Kݟt�ɿ��'�?�" ��~�&����@�H}�����?i���9O�!Q�	o�FU���2��]�#�<|Oxo��M��c��`'�3:X��c7�JX���z��|C��i���'���j
��������I#Z<ԅuL��?�t�p'����t����i�dL���Φ������i(��O̱aG#���T�eB@�nD �@ÜOQ@5j�LC.nR�6���?E���U�u9��[29Z�c(X�4�l�`�]�?�i���?}E���h{�9r�Q���Y��C�1�2U��?��j��%�%�Y_J��s#K �0�<���q�������,�7�,"�.�@�ΐJ��L�����	�( �������	��0�I�uG�'��̘�7| U� [մ`:c���R����-2Hp������"u��O��f ʄ�,)�ddX=%�RT�1 S$ZtJȩ1.PyD �+���#mr�S�q��LR1N��I]�,�B�ލF��S��у����A�b�d�O�On���OʓK�-kQǑ�\p!H��!Xq䥅�`Qౣ0�E�|�[��)J����i>U�	Hy¬Ա$ڠ6�;peb5f�U!�T(�-�8V�$�O���Oj(�R��O���r>]!�*���P*T� ����	�̾�Q��ћk�6�9"�*�D̄�I[��T ٚ��6��5F6�A �9:�tZ�a�RcRQ� bR�'������[��MV=6� ��#�� oұ��o 8n7M�OB��?ɉʟ@L��A�0L�����B�*��Ȳ��'ў @Wk�!�~p@�dBZxr���ch���ݴ�?a-O
�zt+F�}��ڟ��O��|�rSg�p��B�`N����E�.���'��%�+/N���םP�p��JAV7&��х���hY֙a*L�Z�B\�U�$�9��$�Xun�X1��qE�Q��P�a���g��)jT[dmE9�&���,�NDؠ)
�~���%��IS��O�m�(y�z<��R�� �;<�@p#�ݶB���*CV�c��'��'��'�[��"�*�9��ۨ\�����9P���hO�)�[ݴ�?�a��d���ht�H).���B���P�VB�>��\��?I����3(*�?1���?9f�n}��c�dS ?*4��C��k��T�@�+M �% 0%O�MZ���hTjIj�������V�Y�g'\p)��8�x!l�QQ�y����2"��1FG#��-'��<���ǅ���ws�H�t*ڱ�$�
���~07��4O!�'s�(pm�ꟜE���}�ԥ�#r��J7�A,�za��?�*�H�(�,S>	:hg�a:�	�<)��ő�$�S՟��%�8D�U��_!@ �!��t���U����E�d������I��u��'����~�̻��`d*
���f�H�x�+%�p�}�K���$2�9x9I�h�|j<%ke(�6
)�8�ᦛ0�����&a�����%�C�F�%��	�2?��o�f,�A�'�ܠ�А��}?)PAL\�޴����G��m\�OL�}���H%g6(5��ۙ�y�eD�i��<2��L�Z�R8��#�e��#=���i�2R���Ǖ�M�Q%��]( �����j�R��V��?Y��?Y�[������?�O��l����+3�\J���%$M�u�&̛�K����òC\���A��^�џ�SUǅ�9���(󋓗j�F���Ϋ~����cEC1Q���8����0o�HsJ�!m7�%8%��D�Φ� q-T�+vT�i�HS�X����4h�M��R�$��<�-ݩ5�8�9EL y�AW��T�<��"E�Y��;E��8"i1 ��<a�i����"ҧ-'z�Xc �#�\�ȷ$&	�}���&�ڱ��&��8Y� ��>I��g�(�uΘ:C�@��C׎j�d<�ȓOgX��˙n̰��T�43���ȓI��򆨍)L�H��ff[�(MhńȓD>���e��0b�V�iO��za.Y�ȓ�4��d_�Y�`��) �&0��o@8��Դc���t��{b���ȓm�4�.��[�f��V�I��̄ȓj��Lp"UE��)1�%�(�*H�ȓ����ᚶvcmڴÐ�p�H��1k
��T,"D'�h��W�Z��ȓojh\z$*%+� �,0;�|���}0M��6)>�w�A*j^i�ȓ&��Tr6OI�u��Y�d��4��ȓ�`�qr ��Wr���Vbx�ȓp{2��ʋ�.��p3�l�-��	��"{�Y�뛮l&|8�+Yvr�5�ȓn{��2Ɉ&n�fM�a���L5��x�KY7c��#� Ӈ<jI�A7D��Q@�P�P��s�*�r�6D�x2Ń6�����ۯs��{!�2D� R5��8�������tq�dj*/D�, ��/�\��jI�t���$�,D�XpQƒ3Y�I{d���)1R�N7D��Z�������J4aھ�$I6D���C�5�Y"f�S)r2�%1�8D�4��K);�����8V����0D���6��D2&�q�� Q��D�/D��2���#B�Q6�,?2�Ts�0D�M'yf&|AͻI��4��/D�2� �^/�A8aA</b�9���<��%]p�q����z��$���ky�Q��	�m�dĈ�%A�X����ƇP�!��p�'��	�^î�	��X��%�c�XY��w�~�*��� *�ʦ���K�?x���� ���h�*�a�;8�E�v�ENN�@��Q��f���+I�.w0�Y���*4��<����[���t�`�0�x8�"�>9A������π ��1@'�.}�d�b�
3.��I�>C��<��,n��e�f�*\�.��1�"�ba_J֑��C�"1��hw�d�8M|h��S�{pM���S�5�����/S -� ���0����<h��H�E���y��ں���]�y	�4*wCQ6j2�����E�Gx�@R� sIkP斂,Td	�����^�k267%0*H`�P�"�-�~��qE��� �:ʓ�O��F��v�dؑ�Ѳ6c��rQ(X �-jcB�=Y ,i7N�W�"=)�wpd�`��K�P�P��,ǣ'J萻K>������u����dn�'՜���kηJZ�[C�'[<@��l?�|R�wP��Ġ��S�X͑�H�A
�Ȋ"�|rB�y���%�PU٠I�%@�a�Ҙ�dJ*\��e�G�D��	�i)p�x��R�8eуlȚtfl"<Y��L����#IkX�.;6�<Ex2��g8`�����~Ґ�b���	��DU 1��9+���v�ɲi�7T����R�<Gy�ቪXG�C[�rN���F6a`��qA/q��4(��̯N�`r�J���ݣi��w_6-�sr���=�@O2�!���I_�n���h��8b���N�/~����&��?���`��x���F�o��Μ� ���'�0��tQ�l� jSqO��s�A ��?Q�f�(#P&u3�e_�D���;Im�ɪO9��.B�t �Hhw`^6h��ö��O������V��P(	���2��>�I�F�nV�eL����D��0�2+Ol|��eU�5�9�#�]�>��`��֧�V�[�ÀC�S�O}⼂c�;��I���Ct$p�'�x��ݲWB��9�Y3@O� W�����;�,pc ��JWF����ߤ
�pl�e}rm<I���	d�Dџ�i�-��b�o�$d�rAP�/>NŠԬ�2x�&��䒀2�|��E�I���%" 7r��r&�:��D�F�R���`�	,j�Rܣ X/�(���[�Q>Q)$+����D���&L.��
�<��g)r��1��C�
Ȉ¦Sg~J?�x�� ��\�Z�{�F�\
P�z��?4\�E8��OA�Y��;��d�>1�&�i1�ƫHp&��Qc�
S��wf��V�n��Ol�"���Wm�!�ĪxV�����@dT�����C�h̦��a��	-��BB�*z�>��d�Z���]c,
!!��_����R�t&���OV��1)����ɏ_��k���[�,lЍ�aaY�S�(�І�`<����-��?��eiI�)�Ԏ� ��N�$K��t�0�X��4(FDT���;@ƀ����!�r�S�'���C��1J0�BD�E]d@F�����4b*�,�&Rzd��z��8e����)�8S�FT�"��K�D�I��b�CJ�<�㭖��t�	`ݙ�3�
5aG�y���U�a��&�&٩���a�0�zbB�>uz�Xc�a��J�� ����JF	O��l�!��$l�i�#N�lI��(�e�B�R�BҦq�8� ǆ��`[����! �hǘSEǺ:�J�xrI@���O��{���E�2��cR����H��Rt�7��H@��RL&����=O�[bO*x��`61�0{�L@P�QçO���I��'^@�A��4j$��B�$L�4,����Lםj�1�t䑧S�X	�@�˺bv���JR�aG���<��BB�!Ǌ�;Q��N���)b��A̓�}Yظc�U��dĦ�J�J��ǟ�:3�W:��M��M�D1|[
Ȉ�0�I�2�T�ፎ�O�R|c��XT��*��Y�\^�Y� "�'q�>�=�%�O�Z�(����!kH�#W�A�Fj4�)S�$�z�Z��
j�N�z���0��C�?3�ؒ�ŐS�0�w8�ɫQ��H�(U�س�Ʉpe������و+X�l�5��$f�V�6,Ζ2azBC��qo[*YOV}�����R@��w��ۑ+�1;	|7�pB!t
�Gs�0�RDВ7�ٕ#�{�|lrT�#ZH�"'DE�6�t�eƋ/�':�0��� ��Ƃe��Wh���L%/M�U��3&��84t؍��Oz���#�}�V��Eb��8�������Z��%aN�*�b"aĩr��իt�����U�Ԩ�	b�V�h3 I���ԟ$�:Q�'U�X�Q�.'O̩�,��4h�`��K�"���1tȅ�. ��K�n��=�Pf	�Z����JX���a�6L��I<\�*@�R��ğ�Z����P0*��C�DyRf�0�X����vx AG垅}`���	 (b�ݱ���`�v�x� �#aZ���
0�F����[;��dT�(�ր�4&��O^�I�1�"�XΪ?���(�8c��a��;Lߜ��&o�~��u��}�O4ݤP�ӏU�Wn0|qVN��-n�4��|��͓��ޅ���z($PZ5��~�&� \g��@'�ʚ���Aڦ"��OR���5`ٴ�
g�Z�	�5#w)��Z|��IcU�L:������t��ѣ��S@�� ��&W�z�r�EA���� V6�hߓO x������k�G-ޥ�@ ��Y��-c�'R j�&%����3-P(Z䨭2��=�LB��'�����a?�7%L/=|P]9��G-�&T���	 ����e������d?��O%��Ir���t^�"lÒ1�*��2nM�Y�ɂ4�^� ��$@3Az
P���T|����؀�?��%�M�剟!_X�S��}��ȽN�\����J�Фpb�V���^�K��*�)곎��;�NT��޻3�0���h�CBLL���44��S#m��)�� X��67�t	��ˎ٦�7��~}rA�?�םTB�O��ws,�!�G55�Php�ܛF��Q��'���yנB?	%� M��a�7T�1s�&�R�VU��L��>�6�xGm
w�"�	��0|3%��
v�j h�X+(���r�J?�)����)���g0�Oh�f(]�D���%�J4'� ��4cQ�	���b>�T��l���g�U� �1ِ����b��a�N�j�� |��d�4S��	�rFs>�S@Z}YP���lCi!����Sq?Ɇb�'�B��D�=@%2�yjC�e0��Թ,<���'��,��a�x?�s��= ��|��nB�_�.���(�{	�L�r�'��xf'��Iۮ��V�M
7���
�n�)��U�f,L�k��@1.�Uy͖Q�
���O���r�@ۧK&�qBmĆu{��`��
�S�b������f. �d��Q��샣��<��3�T0��
0U�x͔�u�|9�,O�Uc�m��4�Yw1U2��j�`����$ ����
@͂jr�"ɫ� ���)ʎ@��-�"_��3����<�gƏIVи%��� |���#9��Y�pim��|�@!�6>&��7��H�X õ��G(<��p��LmH�.4�q򏗊9�az2,B7Zv���C�<<� �Q@+���[���=��D�k���<Y���Gt�E�c�m4� �u-A�}N�M��o�M���!ǉ����'
��#Á��oWE��Ȕ}F�ۈy��v�ʠ�S�� K5�O��@�1�_=V���b�~%J��>�d'����Ć�	z�R��o����થb��(���$5LOR�R���2?�<䎋�qB��-�
EIA*�k܃n���~�mb��	�@}�Pc�(1���Ɠ��9 �O�-��yQ-F�y��,ӓV~꽪�����àݡQ���8fË�v��9�@ʤ{�,I�牑6�8�D
ڄ;,H���?�̕b�E�'�8�� /�=���'%��Ԏ�I_B���1Sf��(O�	��D�K�y��˫~R�h��ɜBm0`C�\��"fK�}��/���y ��5,%�L��K�v?������G�xX�V��.M2z	�g)%v�nd�5)@�� �� ;2P`�↑ �~P��	N����/ԕ��	�5A�<%���0~�:�'�xH���I��(A�f�T�@�:�b�+8�)Se�"��?C�n �~@�8�j�7k��N�4QS���aCO�"N����>�qOXI��3��?�� d��i�9KP�
Z&��%�8=Nű�OP��6������u"�=GZ�$�W�4�&��㌆�+VEB��v��Y�`)��'� ��Z6�Ze�V�؄ .O����P��r�6FB2j�x%k�ϑ|4�3$�`�$$�i�8II���O?��eH� p�R��*o�����cݾT	c�� uZ���X�����ͻIv| qu�M�`�nTqꏇj�&��	0��u
�V57 �y��d~�O@�5�pg����3\b��T-�reU��'8�U3'�J�Kd�n
�L<��/A+���F'P?9=��c�'}��t�)����۟�E�BPrp�����4N���C6�
���$V&BS84i'ɴk\��N�<\��|}��4}��ڒ,
�+f�xCA578�K�_�\�'�q
��ےDcue�,Q�(���OH<��D�)g4�R/z�@�x��ԃ�$�pB�@P�S�O,<�j���[��y[u�O�F��P���V�.(��������i�A/%�Q���wk�4v璨]n���b�/=��!�H��He��J�S�'L��骣m9/�|0%&�7*��������HO�N�62� M�dB\2/��!�w��S�ƿ<\
 �d��0�UЏ{��8'�O����p�(��G[�R��e�C��X�F���P}�%C=Z�$��0� vN�E맥J	�O�.ΡQGv�����Lg��	 �nU|�'Dܬ�s`ı}~��>%ω<���0}'@\��L�
 �y���ߗ-���s
ԥiN����D(�c��������c6h�$��2�@�i�h
�!Y&�L ���HO睨,���"Pk�;~���	��5��O��=�}�$@9�X@1�(��5�t%
A��9�đ��9���s�#A(R$��+V&U���=b��Zr��":ȼ�$����H3�NZ@�7n֬MhJK�]ceȑDӓ�
,#s�Hty�)W2�v)���	bQZ���o�8�O��# %��
���B/o`��&�"��RCHZ6`���%
Y�^>��'�!�4�HBTm���	V��3���.(� L%��O�e��B�5}j��wjɂVh|pG�_�!(UZׯ�<'�-j��'1���<����q�o�CP��2���ėx"��i���O����E��3���ʷ��F,8ZW�ߚ8�Q��I��s-��ȳ���8	X�w���qg)����0��<p���{BE>x|�O�iո4�J�B�̏�>8�ēS-� 8�(]���^}�,��*Q��B�-lV�!k�OH?����E¬tv9�@���X����E�&_��Oh��Xw�f����Y&��'ƌo.h�9@��܍	�T�!`V�1LV��G��m��ܚd��S�F.�@�G�����g\5���h`�.��ɕ\�?���S@Oj�'��N�q�
�XD �,
�*D��ˌ���&V�Ƞ��R$�~�S>�'8=�s�^ı�Mٜc�x���C�~".g^ų�Od1�6�Aܒ�II�@|#��#�y
� (	�V�O�'��dYvGͼl�"O&�[〟����	-[n80�"O��C�?'ư�SԿ2�1���a�<��EA='`1�JܓY�����\\�<9���*�z���S|������r�<if�ލ%��C���V�^0���p�<! K�GGnU�R�����aLl�<���T�y����L�X�R�E�e�<Q�������@�
�����]�<���vZU��
����c��[�<���E.�X�!ܜ~ �ۄM�Z�<i�MU�2�)@�ٓo(��cp �\�<����'Z*�$*�@�|�Hӷ$�b�<���/\
B��j�l	L�k�^�<IC�%_cD��$Bͧ	��k�]Z�<!�#��x��ɹ��!G�v���kWS�<�`iJ�Q�F-1F�ǚܸ�9ҭ�H�<I���ؐ����,i ]ǋ|�<A#Ş3QD�!�h{�4��gdQ�<aQ�!$���D�r(@�jv�QK�<���%dUy�L��7$&��T��E�<q�ĺ :M�!�Ӿ�yf��C�<�%쓀$b��1��4}\�X*��C�<)�M�w/2��󊘊 ���i���A�<���$Q��_zV�y���s�<A�ZdH���a�O<�1�2�n�<�W(I�6�(��i]/2������P�<�#AJ��t��M	,�"�:7��e�<)�D�2�<�'ϙ%Y<�:#�2T��@�$ާ	��	�`�~���N8D�T�ׄK'w�Vj� �2��E��5D�D)�EЎC[�՘��("L>U���-D� �uȗ�T\��Ucx �(�3Z!�&�m�3mK3tPDQ�.G�S!��!VJ�d�sK�CJH]�k�U-!�$M�l�
� �hfQ�2�Ð&!�D��;��&P&�Є���1�d"Od��@a�UQ��w�>�s "O���Ư�.V�8c�f�D�"O�pW�-.�D���2o�H��!"Oj�+Ӣ\v���9%$�:ni"���"O�Fc�E�Q�qᄘJ��٪z!�A�e��i��_X��œR��}�!�$��f$���J�c��� �kU"n!�dD�⸘��@oL-
b���=!�DJ'�D�9B����RY�@',!�D�x]��Q%-�/@>q�FhQ�=_!�$�%t�����Ą��/D!�Dڶ4Bjx�È����hfl�3!��&b��� tc������ �R%a*!�]�@���i �J�D�����eN�Iz!��M�R�����ǜ\�F�h�%ı,�򄁏Mu����#X�g�S��Õ�yB!��@k��T�f�$0�����y�G�r�^q�ĮUӊ\���(�y� ~��'lъC��H{2MB��yr��7u����ۤmp�����y�؎9����K�e�#g��y��H#��G6f��Q[�JϢ�y�i�*l*���d�r$��\�y2&M�o���`���0���+�N�y��W�w4�%��(�� 
q�'�y���/'���)l����g�Q.�yR�Ϙk�r]p���g�
׏C�y
� ���F+��/����Cp�t0�W"ON k�K
0+@,�*��L8v'�2�"O�\i�ɗpF`�R�bb�Cr"On��G�K��0�Ԇ1�P�p�"OZp��)-��p`���\��"O�И���Q�Ľz���y��D��"Oh��g���s��Yu	�y���&"O����X"lm���1ń����3"O��:b�^-;�i��G����
O�7�"K9QR�VPP��T�!�$K<kX4�E덠���(�:J!�� h��{c��6�"t�W��	b!!���|��
�d�I;�N.S !�$ͣ���1��V �岅�CN!�DM�/�LQ�Wo�IJv����_�!򄍶4�X��&@��}FJtJ����!��ځl����c�F3R�ϋf��O`-q&���a�1B�n24��V"O`���ҮMc���c돃I�"Onah���2A�JX����:���"O���椖p�t�U"�M�13�"Oz=�� �rFa��?
�C3"OT�� �7I��Q���R��D��"O�䪠�@8X�PإO�r��١W�"4���1���$��p��W��1H�#D���0�V��)Y�ʂ��qba7|O.b��0!gE))���H�'�b�	�e�3D��;�C��ju2w�m���0D�蠡�)/̠e�a)�{.ɐ��2D�ps���>���
ť�8�@���+�O`���3 �u맪g�B��4,��yY�B�I�7�D���(�.P$�[�P�Z"C�ɠ�
es�J��1����+�C�I�W�&��P`9,]��kªƐ~�C䉗�x|�sN��iZ��Yq��� �C�	^m|��h��,�`MC���C�c��Չ�(��,b>A˖- �z�B䉃S�@� oY�XnԡR�'^�S�XC��
�y�%ˎ�s�ʍP��ے_b������O�50w@Y�O \���ý
���a"Op�צ�#L:���D�C�v�@W"OF�3�b�i渘�R���+� �R "OB#��O�K�0@n��>t예�"O�eIӋ��D۴hs�M�N[!D"O�u1�I�@�ХK�f�a���"O���2S�	��5fYD2g"OVPа/�?$��!qt�F�)a��Jp"Or$��-φ7�XMq�[$[:P*!"ODԢ���j��Ѓ��U���T"Oޠ�a/�	$Q:�Y�	@C�ͩu"OҩSaE&=4���ݛNV��"Oh��#J��΄��RǞ�N׮�h�"O��	E��}Ve�Ʌ���0"O�ЪV��1n��-�w�G�88�r�"Or�(��G��8�f�+��}�s"O�[�Õej���@đg�l5�"Oz���_�g��oG$P�LyR�"O� y�O�=�=��H�2��(�"O�x��ۥ6�2L�`�L?V}�"O�]�v���jQP|�4�R�]G@(�"Oe�_�tQ�IdFȎ6#� 0"Ov�xs�ԶL0�X���<2�P(�"O.�N� y��I��	�I��(1"OD�[#G�8)F��e�ī�D�xR"O� ���s�"#�ؼ�F
�-5����
O7-[�$�B��l�%\l�tCT�_"�!�$�Y�XR��G*qR^YA"+:?�!��ұF���稔*yD���*�2�!�C,�&A�䮝4he@'�B����hO�t]��-?y��ੵB�?�x�V"O�90�-������P'��$�"O��[T���6s���eɃ�p�$�"O���S��8%Q��
W�T�Q"O�}�l�4�J��' �d�t���"OF}A�̂�:���alГu!ȍ(B"O$�c �clm6�UO�љc"O8e`�`O#j�uS1�ݛL�s3�'��֦T}.�ɐ�C���p�HS�w�!�䓃T�,�z��N�|.(� �*w�!�DN�1�|�cO�x+��+�a]�E��D/�O��U$l0{��I����"O���D#SO�4ʐB��"��j�"O���̗��!/yi������5��'a{҈ u�\i	��(
�\���K��y�H��,��(�z:��q�[%�y2k�W�ԭ�`c�y-��� ����x��&M!X=f�U]�j�r� Z�>!�$�3.y����΍#pN�+���Z!��/xL����f�Vę1��5�!�$�2���d��tL�J�H{�!�R�y�RHZ�a���\�JG��!�K�W�`8e�/\��H��G�#_0!�DN>���C�ԭ���@�@',���%vV@�T�4l�lL�sB��yrK����,��f��c�n%s	ϓ�O�9��ɟ+\l}���E�5d�"O��qAK�52��˃MG	�48yw"O=;F/ܤJM��A-�1Ep�(c"O���qg=O��-v�X4���yD"Oj]!�`R�:� �j,�i�"O���C;���ٔ��1f��`�V"O
�2R�fΠ|�(�5xz�	�"O �1��O*5-t�C�'�1_�tp"O�2-
�y�X	rglU�(+�l{�"O�0@#��7��Ċ��W[0~0S�"O����A�"$s(�U.B�1F"O��)�M����]XV��!.8BO^	��+y֬��oM�s�<Hj�$D���&�JhD�-����nI�W-D����e�RdP!�;�>���.D�����%-����ԁ8�@��W?D���4)�,ƺ��cG��&D;�B=D� ٰc�"#(A�mB�y��5D�p������,��r�]�Pݚ�Ieg>D��p.�$�2銤@Z�PI�O=D�,��P�1*B�(��9�d\ʑ�>D�鱇�#�F��gVe�m2&;D��3���1� =S&��?F�����o&D�dH��oaB�D�(�b�2%�B�	+4U#�q3-�ԋFOZB�I"WO�9B�ԏO|j�31��N"!��}��Fd_�N�1r&!�D�O1��ТE;m�v	�eh�Q�!�$C�!�t�4�J8@D�L?.!�D�p�d93���,A� �K!�$_����N�'~j���@�\�!��Y;ZԆd�:n�`6��!���K� �b��ASv!���)sP!�� `u�g�_�E�)�����7o[3"Ol�*���{*Z skDd��q�"OXY����@�by+c��9(P��&"OB���юՒ�2��6q�l9�"O��QbO�W���j��j"Or*�M����8H��N�G>d�u"OԬ�o�F�F	����2�
*�"O8���E�
[�HѪަJwLL�"O�l��G	�\�V ƥ4\�A��"O"�J��֑j��	����m�pM�"O�r֨H�I6�P�˓�`�:���"O��B�M:��$����d9�"O��
��=5Z�	�%�� ]>��1"O�tQ0��!f�2�Y�Gͼt3�a"Oq;gɈ+�T�2 3Gp�b�"Op�{tE��Y��@�o������'"ORՃ��q�DP"m�2D��2�"O�,†ȎHq>!Y�KQ/M���"O��J"�A2����˧l�B"O6ȡ��#�b�ߌV�L��"O:Y ���~Uz0A�+-�y��	�=TH�`z�mZ4!�y��Q>c���bC ��U]`|�3�R�y�%&!D��rm��%��8�����y&ޮ+%�BE_��|@��ɿ�y��� /HY���!��̺��y�c�,5�0��ft��[�*��y��A�i�x���8s%��Q�,�y¤N"oN��s���^�ҠX&���y�^\%hq�v"�-Z�&�I+7�yr��]��}����_�v�A��I��yB-�]=(�B׬ߙU���p# ���y�G��6�ഫFI�>�"AJ�	�y��ͩy��x��.36@@�`å�y"��>ݲlc7��1	�\H��/�y��Y�hb��+�ˎL�F�%��y���=1H�ȧf��KE
L
�$A=�y�GV�_�ٱ��#5
�p ��V��y2MM�HX��J߾3�8��V�y�E�&�e����1���BN��y���8Hi����C�U�lƗ�y�cW"r�T����#��qY`D��y�?��QB�[�#����e�-�yB��w��lqdCM�~����tgΑ�y�F�=�ƱHrgZ&y��S�V �yBG^]�p�rE�0u��Ѻq#���y"DݗBaʠ$a\l"�2��yo�:x�z� ���0���F�ܾ�y隅/v	3�l]�#�4�	��ҝ�y�
�-o�MЦ���]{�k_��y�H
�*��Ը�*�"-������y2NŌr�Q�1-,�⤙sf�y�δ]7�YkHZ�K�������y��ː#���	��H'��p�D��y�/�:l�D�ʑ����;O�-�y¥L�U�@m��
���`*��y���{�|�`ԵX�I�cA��y�CM	f��U�}��͹N���y����G4�B�l�)��g�y�"��.tJ5OC�J�-�Є�yr�+(@M�>4�Hb ��	�y�6<���S �(@?����y�B�9:HD�q%*%6;R! �Ě��y���֌=c7�T�.�0*T@P!�y
�  M��$Y%>�>��v��Nv�`QW"Od��2ǃYRN� u=sB��"Oj����+i���S�T��6"O�P��ςQ�Be�� �o<EC�"O&9�m��r���BoS�(k*�B�"O�e��OT �,䱱��3UX�,��"OH��d횬RW�0R��7:.�*"O,��	�
�p]+ELC8l�iW"O8l+��F�Nک�R��O���P"O��C��[�i�Z􁓐|�P��$"O����(�ȉ�@R�/� ��"O
�S���.+:�!��Z,�(�HP"O���%�A<��<k��̽��J"OZ��� �,�Vz��;*�!���+��#��@�t�c2'��q!�Q5��{ '���Q*�V)2�!�d�,ksJY�CgUt.ܩ���' �!�� P���d@�&�*(�w�Z09!��.1��}�+S{Ԕ((E..!�dݎ!îQVi �"i �R��Ƒ!��ǃ?*0}�pc�� 1K!�\�-/!�dat�I���Z�[��̲�/Jq�!��R�{��(WÓ�Y;�8��/�m�!�M�r'���@�e�#nH:!�d�r5�d�A�sI��� 
�r!�)(����7Dc���րJz!�䖓G�6 k��@7|]�Ⴭ�,Q�!���n��!���}�ʡ@�y�!���o����_�Z��I�qKܕ9p!�Ă�Y����aM0x����bL�KZ!�D�e�0����#ʶT ��Ie!�$�	�x�1��2�f�Rb�?eK!�ۚz���1�*6�F��.-1�!�D�8[���K,̹�r���-��!�DI�>��M���6.d(����1[�!��K�X��1'ԒiM�t��dػXl!�$]�FS>������J7F��#̙!I!��ԍi���h�-չS��a���ߟrH!��`�t�A�N��+�,��`�R4f�!�D����ܢ!ʘ��&F(FV!�䛲	� ��)�� ������3!��M~���M�9_ (�����}:!�ć�q�$-H$�9�F�Q�,D(j�!�E$V�!���'1�d�Hd���!�$1cb�u�*y�l�P(�-k!�DY��,,�w&P*Dࢩ���	lH!�B�Vd$ܺ�i�z���h�k��^F!�d|�*�����
�ڰJ�!!�$X�`-2��ʡa��PY�Ȍ� !��9ҢiSG\p�:���Y!�Đ�U���p5������x�oSe�!�&e���+OˮW�\Lk�M ��!���U��9���a�`��u��!���|#�P27�K��p���P�s�!�dJ�\dJ�C1�%��1g��
hm!�S�D�T�:���Nw�E�֣�0@�!򄞓8�n,j�iZ�Vg���FDӓ=�!�d�S�J�(!ѩ$��ȁGh�d,!�2E���sC U�̽�d�	)!���?!y6ذ��ʋ ��#�$��a&!�D����ҕ�2�Ner�c4v!��-K��$ƀ1k��aR�|!��B�.���@� B��G ��	�!�ƛo����Pc�(Ĩ�nɹ !�� 6Ty�[Y�mi@a�)
���2"OJ	3�J�{%b�k�ѥ}���	R"O<T���!n�V�ӧ�D�U�R�"q"O�SkԚyO �9�@[�}v���$"O(H�# ��I��𓡋;fk<݉�"Oi�2
U%DBh�%�vh��4"O�Y��*�#�1��<s�Ѐa"O����@�O��݈u�T*FL�"O��rq-ϳ0��T���I�	��y���%)4��"�<����a�A��yH֫(S���2&����@i@n��yR)S�T�"�H2�ҋq��lCÂ�6�yr�I�"�tl��@�v	����y��čX?x`�R�[-:Ϧ���l΂�yRB�>ɤM���̼/���P��D�y�bq���@v�ݛ.?���5�^2�yr%�0S �1��6Z�*����;�y"aS/c���Xᡆ3$X�w ы�y2��l�r�ˆ��dQ���ybH��Y�\��u�D9�Ԭ�6��y"�73}�����H�s#tWg
��yҁ+SJ2<�э�BqK�Ί�y
	_=z����@$2M�y�M%#H`1:�!�,z4�����y��_�x�qH�)�)N|9`�-V1�yB̛.���Ӗ��l�u�ư�y��47�йFG���%�]��y���%�@�ؔ'�t�l�2$�ʱ�yңKEVJ`�@�@pn�͚��ӡ�y2��1QD�e���\�0��m	�y�b�����s�Y�x���O�4�yr���%��b�Ċk�.ݐD�3�y�V�E:H��S6�l��V@��y��RV;�MS����u���,�yR��!g/����!q�~}��"M/�y��DlZdP-؞4��;@���y2'�'.sDI8��,st��w�]
�y�j��t����i���Ht�e���y��Hav�ACƵ=}�*�g�y��@R�H���ň� 3v]b�X�yr���<XÎ��yQ����y"���$X�6����̋w���yb'�u�<�+�.�/|�\����yrj�=��t&M&;�	x��G��yI�{���"�ٗ0&!���;�y�jT�z��x B���yBK�X\ڡ ��N���ς��yR�	:V�n��u�{���;�+��y�o��<`爻uOn�@���-�yre�O
ҰJwk��g��h�BGė�y�I�� Ny�D!A�0&<:���yR�Z3$�qNŗ,����Ҳ�yBC� sҺl�2kT ���2i��y��@�Q��	z����\"aĶ�y2%GB�(hRɎ$�"��A�њ�y"͗إb[�J�q4˯,A\e�ȓQ����F@�#*ܕv�,/�"مȓ$wa�ɍ*_$������,MO䉅�I�
$�3,K�x��4�lS  ���K�(]��&�,l����f�쁆�u��Y��dԞ^� ��2G6.�T��*,As�#W�T�BU�	�	%��ȓ!�`��nS��1Z񄓼M�N��9�X�0&�+��,*��?c�d��S�? �	�΃K��[҇;�L���"O��jW��!,�ԡGG�Q�8i�"O�@����h���H�)���T"O�������J5 E��_'����"O��t�E0	ӆc�+�(�"OƱ`��L�~������r�*Ƞb"O�P��� �r|�&���>��"O�9j�-Tg�����N4p��#4"O�@a���%z���ʐ=,�RU��"O�\P�$�蠴ڲO%�fL!�"O��Q (�4J~��ɗ7L^�+�"O�lXu+�.Hq�Ȓ��6j= ]s"O2X{�cƹf!�+�*�E"O"��րā� ���jޣ~�!�"O
0� �ݮp0�J�*F�68@B"O����m�Y ��V�?)� P"O��0�'D�9?`��3�
 1��Q@"O�ᷨ�
<��i��g�2D),@�S"OjE0�7*R<�W�F'\[s"Oư�A�0P�p&ĈqPU��"O��Ѳǐ�i �s@h�&gF|p6"O�H*�A�_�f0J�Gەm`n�:B"O���N�q_���֥ϥ�N�"O�P;Q�� $�r��*Ox�|� "Oܘ� l�py@0�D$Kl�͡"Ola��	G|<x��bHL6.^���s"O� ����,�����H)(D ���"O�$r�	ΉJ��șfߜk=xq	�"OfE9�T9F ���F52. �#�"Ov������5�4�c�J�k%F|��"O�9�K���y�@��M D�s�"O� @���.���eG�b�{�'����q,ӷzԘ�`.�5��@��'v�S!��d'x�0(ѐ��	�'k� W����M�Эӡv���;	�'�6T���3I( �ֆTe��',\턒w�NL�&�ɰGf���'rЪƢ	;e@�0p�
^9� @�
�'�cC�],0��R��_34����'�����DoS,�x� �� �h��'v�(s@��vR��0۾���' ��!&�V�>B��R��?>dB�'��\HU�`�W�҄��U�<醅ج_�p]��FŠ ��x���k�<��A+J��CΙ7z�� u��B�<iE�( �ԉB��Q}1��Ȱ��X�<���$�ڤ�gD�S`�x�U�<�t/_&?[�g�^m��9�j�L�<�աR�J�ddFx�ڕ��oL�<y���HT�AC�X8.`��`GND�<�D�����5��j��e0FF{�<�F� �_T�)Q� � �t��b�`�<�r* 75�� F�0M6���b�<9W!�n>�݊c�*"Jh:�N\a�<q�B�"'D$}z1���{��łf�<���%S��`���ݷ�����Ix�<�f��d	�$�����
����J�u�<9cY;
e^$���>Zu$1j�
�t�<� N�   m����7�y�ƕg�<��cS�0UR����6׌\"�n�d�<y��B }�n�����	:�@j�Pa�<�ƪ�	S�P�$�D4�
�������錨]�̘��C�@4�ȓ���1s�Bw8MYc@sHU��S�? ��Y���m��	�2$����;�"Oƴ�v��P�Hՠ5B3(�a;�"O�����
klX��Aޠ6� ��"On�̀zKU@��F��AqQ"O���U2N�\��!��,�<�Q1"O�x�b��A%�c��Q�by�)R$"Ob��&��9����ƉZ��\��"O�@���CjȐ����9�BM3�"O�(�p���=�t�8��`�h���"O*�R��.�� �����"O�<B��.w�l���B"b��Q�t"OjL�
kf6�:$��?)�����"OR0�@R�L0��B$$<ofP1�"Ox�J1l[ _���Rc	j��|[�"O�45ꞔ �x	�T�1�2��"O�Ui��1͛��3d�T���"O�<Ba�\\@UPPoy|(TzS"O������F��-V�Me��d"O�ypl��	��(:�E�.r��2�"O|iQB�6v�l��c��PTrc"O�}��"#���q��(���r"O�Q �����:�i��ګ�`4�t"O~�ӱ��v�f��"b]J �U�"O��+��:;�j��$/B8�D`�"O6}�������ǫI��ni�"Orx��[�?4�%�@�nȖi"Oĭ�e�= ����/? �)ST"O"l��.��
M��(7N#�Pir&"O�,�ЮޭD�b}���6%@=ȴ"O�y�EB�%*x�ɣ��%��Q!r"O}#(݊*M��ᐍ7�`�r"O�h�N�#m]|��@V
���W"O`�j7ǄUH8cQo�	({�Q�"O��b�0�)�A�	|ػG"O�����&]����̿_�R�r�"O|�:7�� $�N	[p���l\� D"O ���Q;>44x���;7 ��3"O�ɹA�ջ��AH&$�&k�U"O4�#4,Y)H�L�V�H3K⤰�"O��K -D'E ��Q��3Bx�B�"O���.�"~R�at� ����"O���Q K��%��G��a`d"O���q!C����3�.1IKp��"O�}��@/K��q9���31l���"Ox�R��~ٔ�h*ܔC�P�c"O~Ub���6̺�+.�\#�"OV�$�_l%n��W�>[���c�"O"�@U��~\�9r�F�}0�"O���Q��5O%�٠�BQ�=ܙ�7"O��z��T7�\0u�X����"Ov��'�K4W�.0�&���X�"O. [҆Ь`4��B�.A�&"Oиr��!�N�z��׫a5�5"O�<Xǧ��Y٠UxP��l` ��"O�bH��p�<R����"O5��fȒA)r]�WBw8衫"Odd��$@�XV���U�nK�%��"OLS�j�h�� #�̚.��e��"O���$��$���_�R���"O䜙3��+4���7k�h��ة�"OB��`�Y&~�4|�d	\�rE�"O��ĤÜ$*�Y:)Z9x:M�q"O�eH�-�
d�>J5�S&UjR�"O�Q���R�'/t���R;A.���U"O� ��A�A��pWeW�D�zS6"O�I`���;����G�� l�pQ8d"O�X�b�)
�@����U���a�"OB�A����N��"M��%� "W"O:��uKމa��C7������"OrqNǋ�0����v��8��"O����V%@u(�K-Ϫ_����"O���2���&�cǫX�`/�,H"O�-3���Ed^Y�1凗zz�j�!�d�%L�8��W�qVz�j� F=b�!��8�*-�q��;P�e���J�!�$δ@��YU�Χt�\y�1��p!�d��᫱�˩B��9���ě3�!�$�
Vj��C��TLd�Ag��3!��9�DhD�=��S`o�"8)!�ظG�<B��	!���e�Đ!��3]�8C׃\�.a���s�!�D���ёw��5GYB�� ��:}!��Ϯ6it��B���Vưv�� Q!��K�&�F=0�j�pR�<y`��.�!�d]<����-^P�����*h�!��0M����J�]K�=���5�!�P�M� ���b�4d�A(gH�@!��?+)��g��3r"��1h�Lj!�䖾y�l���A�$�Z��G�´O�!�D@�k'h�H�I�?��`�r�χ�!��@�4����D��S�Ĉ��C^�C�!� L*���J�� �x�aW(]f2!�
u CRŋ��8��'�<!��.�<Ӳh@�v�0��Q q !��!S�؃#�<%����(��v�!�DE ��X�ę�L��(�aHߞT\!�*sڔ��_�{�z�ך^?!��F�A���ҙDb�	(��7.!��E��f�r��xR8���?n�!�$̥����ʙ�-hܬ%�.B�I�V,�%À��va��h�I��6B�	'ngt�h���!��%2M
�^B�I�I.� ����04��%����dB�B䉪S�}Hc9:�������D�B䉕M���```�Rr�(s�<C䉵')�ؓ�Ï��B�(��P�KC�	�c<���Ņ/�VqQ`Y�a�(B�I_��;V�.X<mpq�B�<�dC�I�=p�arU#<��\�rBߵ�0C䉜 ,0�Ы��7�� � �ނN�C�I�O�>	�aJ̆j)b(i��
JgC䉽m�q��̓j�N��ID7[FC�Ɂ7��x3V�U�-�>$8�gA<J�:C�	,K����J��Y�$,z��^Un4C�I6#�����(?�����׶T��B�I��Г"سPĚ�q1`�&R�B�	�#(�8vK�,$3��1�Ӌ2��B䉣n�5p4�_����b��ޣ8mFC�ɲO�N��uj�
;v����'T�C�	8hd"gM�iQ�ɛco�B�	�e$���O�g���9G:~�~C�	�#�e�b:i�@���^���'P��AvJL�>2Nq;�`�, B��'@�mIwe���G�ax�'��ږE�4[,|���bY�j�p�'}j�(7�O>.O�<�ƇP�_�8L#	�'ƨ\�F�Ѯq�h��H�Q�b�'��id� �eq�a��lӰ3��h��� qxM��uݚR��n� iQ"O���Eŷ���g �!�<a"O�q[�eeji��R4�v"O�8�p+ڠGH����/5�"��"O���_5��`��  $�8MC�"O� �K޲@-hUZ���c���`r"OD)� �('P��b�� J�5�
�'�z�@���2l���U�=�|���'�2���_p�@*bn�?1�"Q�':ؔ��,]�#��-�6)��S�<�	�'=��a3L~�y�&b�Fpr	�'I���A�/1�E��?��<;	�'Q��Q�`E	H�����'�D4AA�'�$��Wj��`$`i��Y�I��'�6��!
���( �Ky튙��'҆y�Re�m��q��$�v���' 6��/�.��|pe��>(�'��)!"� �^��J�	<ΰ �'�H q��ՌK68�Ѱc� �����'@��*� ji�!��Ŏ�(0��'�&���f��5���r�͸�rT��'v��sS����u r�ݢ ����'/�mc�@�g�8\Y�Gw$�A��'0jU�eLG'6g5���n_��H�'`>�`���eR�����2��]�'�����nO>���:�F	�.�`�
�'Ӗe���0<)H1;�KؾO^Z�9	�'1$�pK�cth���>��a��'=�Af�
@�0���Մ4� �
�'�¸0�/J8��䇂5��P�'[�RB�ͯm@���&�Z��
�'��\`�I��.����(�	� m��'�T�6a�����7F�i�����'�H�Y��xH�)�A�R���`�'10ճq��E�P��.F��{�'H�(��РH�f0@XF�"�'��;�g �^ھ��2��.�M�'��0�E��VH��!�H-�� �'|��	��I�`�҃ŀ"8��
�'�^x*�` /D�+�h��l��'z-�c*��Q� 8`4��	�'�т��%ʤ���a��(���	�'�N��E�� K`���F�s���'T�E�����;��Գcf�{7<B�'����G^B���{��&�H���'����"-�l
�DT�M3,�
�'��ը�>Y!��Ũ>�*,�'e�)���N�9K ��'��26�  �'�M��@\Gٚ��\�=�t�J�'>��#���<��K�얅-پ���'}�9c�e�a�Į5������a�<�p����2-��ʏ.6'�]��f�<�M�J2l� g*/JM��P�Y^�<!3J�LqnU�t� (��U
�D]]�<!D�'p�&�s��!P��rF�O�<I�J�R0��J�w<��b��J�<��e�N"��@/z&�L�$hD�<��(+\������w	��&�)`d�C�	1u��͂�k
	l��|��Ɏ���C��<�`h##��� �2���ʇC��C�	�;�{f�ɩ6�M��"J8<��B�ɬa�&��ȉ5u1��28k�B�I� �F�8W��dX��!v��r\B�ɻge��R�#��T|i��ٌ�2B�)� RP
��3���G���S̲�"W"Oj$�����<����L�y%J�"OޙK'
] Ǟiy�K7*x�"OT��q�Q�
�	#K�
&�����"ODQAT]�S.��[qX��v���"O~8h�nEM|U�G_�
��D"O������ry�3P��,�b9�"O8G@ƺHL��) ��E�p-��"O�Y0CH�8����#BT��,-�Q"O\��bEؼ"��}��>�=[g"O����d�<�bq�2`[�><��"O����J k�(�V�� ۶s(!�ВV=Ak­��f�@e��	!��8`�0,�Qa�05pb�Q��P"v�!��T�J��]�iI9[~h��	��,�!��Q�N-��"#�qs��b�ڭ^�!���y� �*�B� eN�
� �>�!�D[26���Um�E��MY� �)x�!���2���$P�"�U˗�E�!�P�y|��RE��4�ލ ��K�!�Dʓ"��VE]�d�HKa��!��#�"��	<	8b��P�
��!�D՚i�zp�'��e<�s`�~�!�$�1�n�p�`��c��C��3c!��w,b�Ʉ�Lw�D���*Y!�Ē1ҕb%�>�
��EO�.m!��$.1�Gj�$3�-�Ƥ��!���+b�n�8�GǙt����r��%�!�D�(�$�3F�l�@ �P��<&!�d\t�\��)��m�eiހM5!�DՂf���2�O.rɖ��ǒ-k�!��_�<\r�A��
<�HcS�P7U+!򄑞;L^�` ��5a������[0!��'(֌e� ܍6�PP���I�!�^X[ !Z �(7P�L�uH�>9�!򄘚0n��{W�LN2*A���C�s�!�
|7JU*Q�/f+𭘓ȓ~�!�DZ����J�o(ll�D�I�,�!�č�@w���!���2�I8�BV"E2!�$Z�&S����D[�A�j]�wd��!�݁f_̤�tM�.T4a�5��@�!����<�
�-��3CD�v��(�!��F#=��p�$@k$64��
1�!��˃W(�$��c1��ѣ�'h�!�dբ	i�{E��7��@㧉&�!�DٝT�(�Q�)؁�ζN�!��S.qjN�8���BT���M�!�$�R� }�7�B6pR|4r&%��h!�D���H���\1$4���G�O>f�!�Շ5$*ࠂ.C�t:<ɢ,.�!�����[�@�iM�I�J,�!��u���"M��lJ�p3��<:!�䓬D��-��F �>I��f���m!��>�m�$Ӵ��%H�,�	a!�D~m1��4��#B�9N�!�W*l��\f��,��xR��^|�!�Ĝ>U�E��-
'�~������#�!��6	�h�(���5WM�<sR�'�!�d�I���а;��RS�D�x�!�$J�4�Hj��ݯ!��d����.8!�
>�^�34@�%ޜ4Pf��7`�!�$°x �-[����Q�
`!e�G�E�!��Y�<SС���t�XD��\�q�!�d����a��7�X`����Wz!�� �EA��@0iϰ�C�N���(u"O���F&S�&�{U��O8����"O��C��{�d���,ѻ"O��Ce?(Ĩ��D�٦Jv���d"O`�k�L�!w �	���hsƕ)1"O����,6����B�vb�"O�[�lf^Z:��؛\�u�4"O��"�Z>}ZxG�;z�<��1"O�+�=q��။��&��4"O��$��']
ƅ�F �h�i��"O8�ض��n&�Ԑ�L��Qv`�"OBhr%`�;8���6%Ԯol�'"Od�S�&*�2�8�,3@Uk�"O����"=jv!K�H\�wb��"O�E����PIм����K���"O��: ,@��, '�S
���"ON4�S&�&5�<JWK��d�*!"O�U8e$VB��$���I��^�i�"O�U:@�b �A(^�9 uH	�'3��"f	�c֢hXD�_�~LV���'T�`a�ꞻ65�A���O�F���' J�� W�#�p�R�H&::F���'� �:�ԉG7"i��2
	r�'j5)׌J�L����A$'@��'(t�9��ߛ<��(�`�[�.��5��'����@�]��Zp�]���
�'��x��ə;j:=���ɮQ�f��
�'#�Q�������&A  �%k
�'�(2�� q��Jv/�t�\�	�'��x����Pzx�El��s�����'�������<Tf�HY�Ό e=F���'��|����1x�"�(fCH,/স��'N� {TE�&q��=,H��X�'�𽘖$e�R�Ʉ���H0�'���C���A��3����P�Z�'o�D
&mӪQ���ƙ0S��)�'[�h�b)�r����N��b�'nVء��({��)��G����'�ڴ2���C�����Ϟ�����'��@9uA�&1��bA��;!^��8�'���U����pU�ےht��'�����_}�޸#����d{$m�
�'��q�MB0y�L|q��	�q��d�	�'Zh=�'i�1 ��d�-�=u���3	�'f\0B�B� K�e	j�V�"	�'?r��D�ħq2B4h�޾iA�k�'�Ȩ��P%A.����¡a�~:�'i�qc�Ċ&���p�koT�ȱ�'Q0Y�I�n���ّ�pa<���',:|�A�
bTp��vh�r�'����6$�-0�T)�C�S='�+
�'�l�Q�l��;+��H��L
��s	�'�Т��\%}# �����{왣�' �i���D�ڍ�p��G�<([�'�@x�A�;zr9�� ��?N���
�'0�d�7뒓7ʱU��6�,8�
�'$������g�8܈�K�"3���	�'�Z��c���I��(�bI�4a��d��']p��v˴]�&�+�3T�`1��'���I��
dW\�b`��D[�2�'���* C�B쮥R��\�@ j���'�b��&7oA*����H�����'n(���_�8pJ��Vb3C:����'�t4�p/R8H�FZ�C�R����� �HZ!�X	(�v!(4�޽$xb��0*On6�c��y%L�6�H��'�bQB���qM��Tb�$E�<Xb�'m>�IMD.8��	�elӲK�����'�D�k�,!s�� ���N)F$,[	�'�D��' �G�
p9��1=`�}y�'�՚2K =0�ZËX�'/��y�'��iJuŢx���r���N���'��<B��% ��	���#yH8�'�T��O�ug��h�`GEqvT��'*N�Q��9lu .(7�(��'e��1n� L�zǎ׏,�>0i�'f�ĳ���)RT����%h�$�
�' Z��т��Y�Θ:u ��l��\��'נ	�Qcخz&@bӏ��t�����'{�Q�ma^�ICLΝmKB���'�T|���p���n��,�	�'�L 3�D��7�dQ��J��Zoz���'ڰ�`T�^:.}��e�W�H���'��Ū0
YK`��j��~��m+	�']B r�i����x���v����'(p�j�����H#���Ap8���'i��9ӬV�\*V�"0�S=C����']ȹ�4�)C�&5���%5E�M��'/�]J%`�@*�C!4�=S
�'�j�R6i�.	�fl��D�}h�
�',P�C�nQ�Ck�I��K�"( ��'���hw�� [n�q�Z!QJ���'4FuI'���[n����oįN,p��	�'�0	k�M(�>�A1�\T��D�
�'�Px�Oc�n4��R^(b�
�'��]X3����ʰ��R#���	�'���B�'u���3���=HN�`��'��9j  p��`'�C�=b�4��'�p04J�V_ТL�J��`��'��1���P!���A��G,GI��S�'�ڭ[#*?Z�*T.\�p���'l���\�@�@�\ v7Li
�'�L�_#P����
�-]8n�j�'����JN�?�֥y3*�6+x��'Zyj��NR��}⳧I����
�'�r\�E���B�k����~���9
�'�d]�s�F�k��2�m��x<��
�'L�(�s��6rxrgo�^-�=P
�'�d�*�(�*��}���ݟV�N1�
�'|��V�Z%6�.��eO���ZЉ
�'�@(A�^9	U��8�.	�'Q4���"˰j�,�u�5
�<���'�Ap�kH���em�/�4�
�'(���0��<E,��(FH��-���p�\���Qe��6�����p��
�
I$	F(���ܐ)2艄ȓ7x*�S��Ģ>���IP�ҵ�݇ȓ1�, K��Jz�9���&h<��ȓ$D����X�p�j�+��!��Q��]8��iM�p�(���L����ه+6�"}���&4�̆ȓ���XS�V!鐽�S�8��ȓ�t�C!�	J����L�~b<�ȓx�6�a��Y��a �ě���Ʌ�/,XB0�F�m�-fA2����
#�Щ��<�0�Eٰ.ᠤ�ȓ_�&=���3�Lr_�݇�i˨�b�⏺2oB#I��Q��S�? 0 KO��vF��ӊN?x��(��"OJ��̔�<�:IӠ��]T�)�!"O�d�	�G����gi 0�0)��"O^y�,��\�<!���:�xq �"ONp��L�v,�H��1/�D��"OA[S�΀[�AW퓜[��U"O���BY�g�^�i�K����S"O���T͕ �L�R�J��g��7"ON��`�-2����'�I�Z��f"O�-���"�$�����3��qE"O<dK	#��!�ѼDD�}��"OZ�����$�W�M�t�t�3"O$0���5.�@��+��9�����"O�*eΙ�]�j@��(Z��yd"O �SCGj������.~d��C"O@XR�B H�<�S'�HN��"O��{b`�*J"���b�ǪNE��*�"O�9i�敢u$��	�在pD���s"O�r��=~W�H����=}9���"O�8`/�H��U��E!F�Ѳ"O���@��/C� D �:�1�"Oq�p�U�G�m�d��[c&�	p"OЩPcR�U�)#�f�4'�a��"OL�b�莟%�R,�t��Z�p(� "O�0X�A�"�:Q-�M�����"O:�A��E0+��8A��^y��"O����)O7B�hQ�,c�9c1"O@��#�ѲS�PT���dNT �"O��"��C@{p�8�rh`�"O�I#�OW��0���GNa���*O6)��,'9cpe��ɽ-ր�
�'Ȝ���ʒ%�M���B��քa	�'�H�!�M�"5�쌒����'�����ӟI�B���/�h��'B��D�ȫ5�=�を2�i�'s�e���žzB���K
˺�8�'((Y��g*��؅o�'��$z�'8p|Zfl�"���BfP6v�q�'���)�����kY�E'����'+�<�T�0F��⤉�6 ��'����Vk�	�(d���#����'�V�b(	'7�t��*BpL�Tx�'��P����A^�9d�Q�z���'8:�(���2R4^�	Ee�?�&���'`�1�F=PfQ��O� Kz��'�di���Ȁ 6tQ�t;`�}��'^ѓ�mӜG�P�`�KRx�%��'t�0+�L�)�b��͑�N�����'\���-���
��G�R\�	�'����Æ�B/Dْ'j�Q}RXR	�'�5��R�<b�X�w X0[*����'!�9�E#L*V���C
N�U捳�'��(bS�ٿ
�u���I&���'���m�����M�#���'[B�	HT�v��p��ϩV!���'K�A��BӘ8(Z�A
^'G%BP�'�BU+�D��>����B'B@|��'(�x&''�`+!!ޠQ4HYY�'���`ӧ"���F��B�̥�'r��ƉcD��D�2f:���'�Ҍb2�U22�t�00��=`�선�'P�HQ/�= �"��G��Vv�8
�'�P���@!ԕ�%-�P@ra�
�'��c�a�֥�e"Y<L���
��� �9)��Z�\�Rh��ϤD�n���"O�hK4oL.y=Ĕ0�H�51?�0J�"ON����4Q�M��-8�6�y�"OBE����f�$�eLku4}�V"O�� ����6(W&r��0�"O�@�5���0R�k+�jK*�z�"O���A��(�		Y��"O�� F�S��q��ԓh�JI�"O��$D�L��H��s�H��"O��Ja�U *$Kt�R�S��q��"OY8�L O�xU��O�,��"Op��s����m��z�"O\ݠb�EL��ы��4�B�"O4��*�r�J�
fk�"�>�Rw"O,�`e��;V�)0H��R��س�"Oj�lx�`���{\�=@B���e�!�D_�G���x��2\�,����Ǭ !򤚽`li�čdgh�q�� b!�D�>]Ҡ	����z[��j�FJ!�Z5r�ڔ��@I��ʇj�:cB!�d�P�^��T� e:z����!��_W��Ӫy<>UA�P!��Z>jΐ�D��i�
������r�!�N�H�r�)��y�9�� v�!�$&�N�h�$]<d9�S�AJ4�!���[l8AjT�V 	2��r ]�(�!�Qy)����c�
A�H� �!�D�:�ϐ�&���w�&t�!��
!J�-9�f��Cp8L��c�=@!�dK�V�$`��ψOc��v�X��!��Ǩ[���5��bZh8��ރB�!�VR�	���B57l����YX!��)ʸ���"6���#��IM!���]�ue��"���D�kd!���"�`�8�@(v������*R!�M����e�L�s�V�_�%�!�$@�nz� e;�49�6D�}�!�$�>Mz��pU�I�J�8�Va�6k�!�$V�<���C�Ƭ:E��f̠sh!�/L�TC�N�z� DKR�Ġc]!򄗮�tp��e^|�(�#�>!��,U|ԭ[��/��vL0!��2?n�SI�?�����ͭ"X!�DF,42U���F&d���)� ��'!!�Y� �Hs ��%�P��0`�.!��?EnxJ��6�� CL��!�Y�KK	Ӕh��^�a� J�&!�D�f�ŰG#O�P�䙧/�[!�יI��Sb�6�p}��ɛ;N!!�Z J-p�n�!F�&�2�bG;@!�$ �xU~<hՋC,�" 9b��% �!�$V�HU��� ��`�>��Q �(B�!�D��*���fǉZ�(�Ni�!�D��^�@{r$۵D���t�8R�!��7k�()$ 8�P�9��:�!�D7��X����z��AB8Y�!��Л!�P� �욗nr,��P��t�!��58�aqG-A�so�{#�\n�!��B�K(��2g\%F2������!�D\�ZM���n*	ȳ���!��	�M@�j̷dR ]�g_l�!�䔌�8`Z�L O����%Ӳ�!�2p�#��% �����ĝxѡ�H�o���s�ۅ?j*d�����y
� �	��ޅm �
�ƕ�,#"OD�#J<S���f�S�'Yv�Z�"O���ɖ' d�ܹ.΂Upn�;�"Oޝ������SfH�{:�D��"O܍�C�?����08���"O2�K�L�Yq�D�1�}*=)$"O@��Hh��%��2��e��"Od����N�rQ D��6�����"O2ɹd�I/�N%Qd��l�8��'"O`�£�P��܉��
�>^UY"Od-8R�N8}���cBC�JVX�"O4�B���Ҕ-YWAP<]���@�"O��3�CV�kV�4��rΊ�t"O~�!ҳKit��ȓZ�X�a�"Ov�1���]�Dqs�	��P�1"O@�Ze�G1zz�I���r`�$"O�AS�-�:tG��ç#,TF��"On8�UdN%�J�f��',LT�A"O(8��Ȱb7x F(_�~K��q"OJ蒣=V=0�I��')M��'�\�&��Đ�d��#�JA�'�xZt��m�ܵq$*W3p��9�'���1��$U�64	�h�y�����'F��`�%w���W�O�qKlŹ�'�4���Ί)�H�2��&m�xP��'�H��*6-�|��!�E�hh�YB�'�T��SL��'�,�X�#�]���A�'��I�KL��sEk�Yt�42�'�Nerr�K"/ Ɲ�4��Q͈�{�'��L"�C_�G2b\J���O-J���'\���hU 
�R����AO���8�'�����	5�vAZ�I ��	�'��i����2`�R�8%G���'��D�r�c�ͨѯ�#P�}��'*=�d��9y�F��M널�	�'������V�9ג�[�D�/�Iy
�'�<0� �c�ε�we٣$�s
�'LE���9!�xh��!�r+���'Ϛ}�Ц�&&�M�t��("��=B�'Hz��Qo?�H]87  b �
�'k�9�!eF9:��bI���M2
�'�h�� Y>0̑����r\�X�	�'���E�@��U�#�ߝ&^)r	�'�V���Јo�ã��3	���b�'�n��7�#r@�O�|X.��'6��i���iT�|�Շ��q(N��
�'���Ʌk�~H�� B��e�(Px
�'�<8hb�ŰO��=���0p
�p
�'fLCƭ�ld>!�'Ï&$t6-8�'��Yi��Z4R:,����
���	�'�l�S�O��b���Ń`��,I�'q@�3&��L�X������R�>)��'��-I��6�L��95��r�'�R}K��O�2�;�G�1`�[�'����A�[랭Q�_�0h�P��'2���	=8��� `�.��
�'�
83	��q��9`BD2�d��'�t�A�	�=�B	a	�~���'� ��{n�Ж�Q������'gz�8�C�o�ҵ)	?Ǫ`��'�y�Wˀ�r�a!p�*b�(��'���d��]w�����S�*_�9��'��[�a̾t]�����1c���'�� I��=6��ԓfCw����� x���s]���+W8*���"Ol��!�SnNEЁ�ٖ+ё"OnM�&oF��E0��'2�=��"O�Y�Gh1E`t���(I�zY�u"O"]�7�����j÷g����"O2���9_>�[*j�r��"O��&l	%�0р��p��"Oz=b ��u��!��e�~\�#"O΁�c�1;vM��G�]o�p��"O�-��W(CR�9�H�<�ac"O<D��Is�y�c��:x�+3"O1`�a��~l8�UE��<w �Y"OB��Є$-�J ��b��6���9""O�x6�]�b_�ȳw�غ��`"O$�qcOK��j|!C�Q)�� �s"O�[eظGG�\فBұ	�\|h"O�]�ǌ͜FK@YBPb��1"O�����L�{���jc!�#n*�!�"O���b� *)H@� xk�M�"Oތ(�B	�py|A��PG`M�t�'��D�<�F	��U|��N$%Ɣ �P̓��=�c,[8&�uR�ҙM5�@a�L�<�B�%w��q�$U�h�������E�<�ֆ�(uBخ<���E���'��h(O�O!��1нb�G2V�lȪ�>��p�ēM۾��Eʑ�fьӔ��|:t풕��`�O�p�,y�D�d�*O��[��u�<�Q��:�2�F/ ���!���t�<1���(�%���K�1" ��6���Vī��ַ>����듇8�c�"O�T�Ќݯ9ȊM�W$>p7 ��5O K(Oj�O~�<!A,��__:��R�ǓS�D� ���S����<��+�*f5+��C�|p{��H�<�6�ؕkd(}��E޲+�����[Y~�\�0�O>E�$+=bK`A!�%�0p�VL����y���{h ��i	�i}��2�;�hO��$I2N�����hZ2�����'v��	yx�� $#	X� �`��
�B���(z��q���|�'_ўt��ZBh���WG,Is�%D�������p�L:��㶹�t�!D�h�'�D��Q鳍��,�����n4D��r	�7?��$IꞦ4�.4�B��>1�'��{RF˵�x��#5\Z5�@ψ�y�@A�	�Ҡ��GM�Nh5�R@N��y��R�����ȂHgԴ#�^��0?y)O���;v��A#��B�T��Y�"O�y�&-�/vp�ɂA�r<��3"O8��V��WB�n�x��|���ɓ�ca�}R�U�m"�$Z⫅�Pf�'��|���=��a�刖���x˗��yRl� )�10�N¥s��Pu���y�$�4]�� ��`I6}����f���y�AԳ: �(�_�x|�0��'&�y��_zs��3��A�o�pA*����M�	�'�~iSQ�;T�T�A#�!T�Ii�R�.�S�	R	�B���F�rV2�3ŻyZ!�䃻[>�{��֔>D8�%ЄpX�xFy2�ċ�J�G(�9�E�U��0��#D��V,�]/z�s�F�LP��n�t��ɘ��,���)	 �Y`�B+W׸B�	`���C@Ę4��X�΁#J0�B�	��½�	�rظ��wG �e�^b�`E{J|*S�Z9YX쬘�OS/+4�k"��q�<I�$P�3�i(en��,T�sA��$ў"~�)� h𸄃��R
z���'T�i��4��"O�L �U!҄��4j�E�D"O2=s�f�:��2�c/;�-�y�Ô�C^ބ#\	J,�Q�B�y�dM�P��X{2Β/B�[��+��=��y�E�.3��b�$J�K�����y"�)�T�6�i研�	���˲M*���'�ў�|�)�v��ݺ�)ݣG���Z���s�<���OAZ�`1�ٻ9|�5�*��<�����d���JE�J��as穉�^J�B��N[2D�偞�g70��G�?��B��<(�P �%ԊRj8�%B����8E{J?�	���,�D�q�h����a�/9D�PC0�l�,]��^?[��]��5D��`�ɕj\���]"����.D�$�U(B�)�+Ĝ��I���0D�xPq�J�Pn�hQb˘�K@�)��l/D��s��E=F6�c���6�t�R�I!D�h���R�Q�S�\��f>D�TqG	�����䙡s�r�xa�'D��PQ�	�5������,3%a9D�x���F<JCd�Pō[.����K7D�( !ـW���d�Ya�)�.!D����f˙q����	��vJ�]�Т?D�X"FH9l,嘷)�4|���=D��2T� ��P)�G��@��h@�*OV�s�$գ��A�p��gO:9��"Oz��"*X� :���&��/2,�y�"O�U�хl1�lX焞f���"O�(T]ZD�
 	2=�LL ��'�ўH8��N�n��m�Dï* �M���.D�����~অ�T/p���
,D��+�J٦x�Z�
+��E�R�$e&��\����;�U FKF#��H��m\�	W��Dp�@�&�S$����!��K����6sr�@敫$�DGo��Xj�C䉵F�恘7���<�L$sƦ��1^�C�(�$ls"���|��5����%�'��'��`�`�E (�0�!MB�+�lyr
�'��+�B�a�:���ߪ#3xt �'�|�YM	%]�>H1B�$gr �L.$�l�f��"�J�x%���%x��4D��E��9I�X��AA �BJP�>D�x�l�)xY�9O	 Q�.4���)D�|�%6%u�����']L�A3�(�n�`��8§-@�V�$"2TB�I�o��iCWˍpR��9#�N�`x��ĥ�tH��� ��i���?z�v� ��:��x��ħ7o>��*�/w�~]�.E���xoZl�������g��A���Ԑm����J	l�C��@4A��3a��M1#=���T?m����&~(fAk`)7TL�pZ3�%O�#=�4�D�b��#2�[9cv���D̓�hO1��;���M3��B=F��e{�"OJ�S�n��)��/E43�,(�T�|��'@<�ѧ	�V*䅢R�1M0��ȓ��䚠
M�|�y#a�+&��͇ȓs^��� �Ũա$!�/Iz�G{R�iў֝	H.�
'B?$l`+�.:/�C�ɖ6�蝁�/3m��u�'�,rC䉳N]D14��?Q1��B�_/et�B�%<���)׃��e�*�B3��1k�B�ɬCT�h #�C.@�ц��x�Z�'�ў�?����" "MT僝f�`p��D8D�� >�9��^}�,�D�:}(��T�'���t~R��L���3A�\ċTǊ1��P���!�!���a^D!5���t��]0�nذQ��'��Oؐ
��D4Y���2,��&)�M�
Z�!�$L-F�dp`��؜6ٲ��Kƒ�!�d�=u��9�bgY�H���J�!�$�+�~I��C *��H��;!��=*��q����T�aV
 '15��yR�'�J)BR�O2�K��!@p��
	�'��!y$.�-�@9IqNދ?����CO�G�ў�
��S�l��h l)���A�`IO�b���}��'w����� �lm�D)Qz�~P��'�����* ���eιv�>��I��E{��N��|M�]S(<B'�c`&P#�y�F�$�������g��H�����'��O�˓��$̕}1�lY2D�3(�]!4]�X��$ �zm�����*S�%[��M8.$`��'zў"}dW t��D��ظPD�^x� Ex�0<2|DH���Q,�I1�φ�y�	�6�8�ˇ�Z�zx�-@� +�y⪛�n�*a/F�e�A� �,�y�b�1%TV0xpnBa5f�k0�+�y��Y�}��ģ\� ]q�θ�y"���XY�h�g��N�z�bB�y�놰Xo:�+�c��@V$1)�$<�yҢ\OP!�n�?2�`�b!m��y���45� T�v醫Xp$��B��y��_>@x��6�׾X�d2Gϝ>�y⧏�/����A*U� ��5�ո�y��F W�R�Rр�F��e���˅�yRO��wSd�CBNrd��h��y��RDp�-��*̞:%���J��y�h�:r����pbݑ1��DA2fϰ�ybE8r2@]9�d�	U�ZubЋ�4�y2 Z�BLf�!R�"X�d��G���y��N�xʲ1�"�N(�z��@��y�o��$�l8�4���21���v�ݧ�yrDW=>}6�'E<|�4�֍�-�y���:b!������nU9踑	�'2�qa����9mt��uKSb�\�;�'�p#V��1����jE7q���:�'��y+  �9Bwji��I�_���'�m0�j�0���hS�_&��'�йf[�nH��J3�U<_4�3�'h��Z6�	(7F��
�(�0c0zL)�'h�<�#�^Iw�������Y8P��'Ve���\2# !�Q�M�W4ڝ��'�x���J�7pO.is�"ۛL�|�
�'麽&�E"�P�����I	�Y��'��a�B��G!�i�-@�t���'p���C/ɗ�2t9�oǼh����'16A�f�T#[v�Y�r-B�_��8��'��A��	�9sV�89�'j�D�
�'�P��J�,<����'C`��Y�
�'��V1~C��A���!ޔ��v�4D��Z)0m�nd�2�ڀ�`�S �/�[�<xV�+V�ic c؏p>��Sf�A��8au ��!M�KRh������QdF���c���t�a�ȓ2���G�W��q����$~L��p��-ڡK�^�ap O<B�j��4�Tdyԅ�	b�2���ۼ?F����ԁC�^��]�E�Ugɞa�ȓ>�tX0L�?z�\����;����+:�9��պ]��I�3)Ddل�S�? (��ReN�>�H�a��/4�2(`"O��#�/�/ ���OUBV�{�"OVt"�#G��; C�.ʱ�"O�����a�yc�-j�\��"O�� �ȼb�t�������X@"O�d�
�1kp1�&���1�B�j�"O� r�(��ƚ�!dF3h�:a��"O��3%�&�(����S�
|S�"O�\C�hK�H��D�$x�$�r�"Oฑ��!�@�s��՛����g"O�эQ�,�T �t	�(x	�iH�"ON��E�RK�� �+7
o���!"OLt��.�=6�\�M�!W�d"O~��5I��R�ȹ�a�ŋg4z�{�"O��֢��w*��0D��rN�	�"O��*f�y��e)�cNr�\Ȳ"Or�!@��l�N��AT�f��M��"O�lZ�,=������Z.wn>�cV"O>5��ʶ� 9��2|����"O��ht�J%4e6=3��"�¼�"O.�#B�B�g��{'<q�E��"O� ��ˊ�.�f�y�FF�BqD�!"O�Q�]�n\��J0�Oq�3"Op��@���*��s�I*t(�R"O� ����M�$��gɕ"��ẖ"O��H"e�8P<,坍d��9�"O��'�zh�a���~�0��!"O�䠗$*/P�I���W����"O��� ��WD�b��r+�a˴�'46Y0���d�6�&4;� ��#ǰ7�p��,D����LÊ_�T03��ńuc���&�.�I:0Dn@�'�'=tI�f�4s`2�C،�r�ȓ?SR��Ӌ\�)��ܳ/��l8���e�(��m=�F��OJ����	!}�<�"0�I;Ƭ�R"O�@ $C�;0�jT�p-�Ud|*B�E9r�[�*&�O�܀6�Q;/.r���M9hH���'=vH�睶'��k�b�P��9��(��U"@U�C䉴j�����[2ET������,%,Nc���r�R�&+DAG��np~�D�F�p�N�V�C����z�<��Wj�4B��@;��3t/+��pmH�1���p�/��4�1��P�H�5���0��/%y���V+I!y�"Q�T�P]�l�B�'*�OV�Hn]�S'd����ľ#^$������c¦>�b�o�LpG�*5r|�WB?��T�Z1��o[�L����ۇY�az���'q�b��]��W�*B��i�pDd��($�zFְt�ڇ
B��a�"A�$#}�'�4H1BԆL���iƦҧLTUۋ{r�'�������� sA<x2�K	������+GP0'��&��Ѭ�M�ȥPD�� rC�02�m�z�0b��D��;�,�#!����O�2ţQ�A��-�(H�N"��8y�(`��@�&чd� h��'��|�'cS(<�U��nV�>�6��J>��.��<�<���	{58���ߔH�n���J�~�CA�!�h[%
B��J� �Je�<��I1@��@�B͕Y���燁�c��;t��+�L���/ry����D�>�杲]��P����
SqUY%ᆏ'V�B�I16��%zr苘f�$�[�bΚs�9++Z�$���)�i�>!&��g^�!��5R(KY�'��0�6���!LV�z��<k�=Z˓'A��2��==p��+j^C�đ��Y�p� }���N}"`Qk�;���!�hP�p>a�CF�+��D��B��u��R≅k02�۲�ޏ �j�P��ޞ-��|�Fc��,����L�D��\�K&�����H�Q�ȓ?_D@)�%L;4�T`��]/G�\�se��wUڄ#��D#��)�RDO�=\@���	�2�OļӬ�'n`%ug[�D޼����@H<��i �c����� Ѡ5��(�Hų$d �8f�߻y=:�A��t�B��@�`������� (`��r!��0��`�cHU�n�ayb�B�Agށ�r�Q�~�H�qÄĒh� ,5�Q87}��v�Q9�z���S��k��'�.�9�fʓ
�F�B&n�2�"0�K<��̜#5b�e(&g؆<��t��\�\��1R����DဓT<�`���)Ԇ���y
� ����M�~���vD�8amR�bC�̿��!�	nK��KfF�*6v��H~�+5s��X�H��$����%F�|3%�1�!�dR$]����w�l_�0���:�N��5k�|l6EHl����#��_������.�R�h�NZ<f��p�e�v���	4yȖґF�:]%�`S�j\.D]`-qVo�a���2���>Mo�1[�Wc�:�1���h8��B���:�t��c��/v�ڝ��/�䂵^蠭w��}J}K�G�q8p˥Z:r�:���K�B9j�K�BP�9;�`%%��B�ɽc��@�B�0IJ��t�ԁ!R��fMQ$�%ä �JoX	 �b�OfH8B��߱i�!�O���Z�꒼]u���POqXF�Y�ߠ�h��%;�BA��^�g]y���B��y��h��n�yKvL�ٮ�<Y�k�����q���cW"]lx��	!��s���[�"\�A�&q!��=�>�#���!sF�K6-VC����lC=C�a}�j�c����Q�y���ɇ��(��y�����&Y)$�x�L�S���	�}j��'|c`ܣ1��/`�B8�@�7Q%��~[�M;�W>V0��x�m�1X�0��%��P8v�[u��t��� N���O��y�w�(�ʕKK�c����!o���'��V���j�(�p��ŧ�7���K� o���Tʄ4_nz���l?u��"> ��-gϰ(�a%�x^�r��U؞ 1o�_JT)�r�B�Y�؝Y����rN�\C"男P�"Y�r����?:Bh0vg�:@
��hoR�m��H�m>z|�� l·t�4����D	�*O1FM������h����yrL��6a����ص�Չ]��֘��ӆc�`���+]���9OȽk$�L$�^a3����Z��}"�"O6��o�Wl�)���P�K�Y�ȰrͱeGl���*B8���f�.����a�T8iw�!�"<O��Q��d
�}X�ԝ��d�hH$�	�����$����}�e��n]k��_*1OlU{�]/n��/�\Z�lo�7}��'\x�2�cr� iwN�!_��\�ȓe*��b^
:��ˑ��&?�bM@�!j.꽐s+P:�x�s-D�O�fE̓o�8�!qF#ȴ=��Z o�� �ȓn����B�/��ز��О2��9�&̚p.���bϬ	O�	�(Zú������J�P	��<^��(�4��<y��{��I�xܳ�)��H�X�Tjӳ%o�difg��A�%�f�ՑK�29���r�Ɲz������B�s��D�Vڜ��������%�)��"�塅�=)���:�!�S�!��&�H8 bl�e��y��O�7n���D_	B���̒�/�)�������$(�SL������(D�(Ғ�3k�#G�Q�2z��Uc)D��cd��y��C�N�]u��"��$D��;Po@�8Z����O�
�h�2�e&D�|��� t(2�"R�V5n؆g'D�|�����"��{��Ҕn��Y��'D��0�i�`�����.E,��$J��#D�����4*0Q3�%;:��3D� ��D�=.D��K�k��(����*1D�(��-*D�ؚfgӣ\y���:D�x#�o&T�kÇP�-R�İ��=D���6lB�Ej�e|��G�9D��!uI�
����.���4�C6D�xSF��1L��`�X5Y�`���:D��Z��^�4��y�S+W?Xw��
c9D�|B��E�Y���$��(O�Ɓ�b7D����~�Vű%�?�q�7D�Z�jC��H��g��M1��2��5D��`�,��D�E�9���x�c7D��cW�@��2�%�@?`�Z���8D������F�~ ��j.
��"4D�����v���թJ9Uv���'�3D�X����k�-	�h8�\��l,D�����L��ԃ���Yo49�B�?D�\	 �ԤZml�qR�5}����&D���ׅQb�6-8D�@1����1}R�H�`a{I�7e��hA�G�*���*س�0?E�K��)c���h��9�''��B�Z�o_o�<� ����jI�Fgޡ��Ëh�FRU�	�=UH)��,�'f�
��`�G�FT�]I0A��꠨�� F����F%8�Xy2�+
S<4̓Y�~h��U�S�Oc�yA`��	!R<1ȇ�U^�%�
�'���bD�/2���f�P�@�O�E�u!̎ �az�l�
eTm���0
$=d����0?�&eP(�r��?QB�ʶC��dz��Z4KHD�<��(Z.��YҢ�F.\򱒂�A�'������STL⓯��0I��b��;=�C�	*ol�@uK��H,xt/�&$��C�	,M41�H[8h�*d�2(U2��C�8���#e�S��B�4LdC�I% ��БG�U18��y��N'}5�B�s�,Ѩ�<�a(X�SlTC䉭<!4z��+*������$C��;ȔxVa
Rrԥ�V��~5(C�	
?6}�F��:ؒ�Xp��C�ɶ*  ⦑�P�Q�4�ٿ��C�	G�PH RL!7�A��֫vhC�I�B�9Qa�?�a�.��8��C�	=I��t�,��F4B��0+S���C�)~�Yq�d�:�N�Go%�C��a����ߠU�]p� [�PAtB�IFub��3e�zع��V�d��C�I,M���D�,�����!֩f�C䉖UL��#��@�D.jȆ��|�C�	;9�dȖ�M�nv%�%k���HC�	g���K�!Y>#�JQٷi��w:�C�I�hzFlzen�.�2eH+�)`C�I"��iAՓJ�<]���Y6)�$B�I�,�)�rhلO�NM��k�IyB�I42|]`�*�9uo2��+1?��C�	��D�V�L7i9b�	h�C�	'A,�k����u��Pa#A�M�@C�I##0ن,�5	��|{�&^46C䉖,��)7��0qV��hB¦C��3k��|����k;Dt!�땓m�C�ɴ� x�e!�O�B�;VG�:��C�I2��$�1��?�&��0f7�C䉂-���c��V����ҷX0�C䉭"f�5�l}�<�)��?�C�I�u}֨�+%I��źb��J�rC�	�i[�2t-͹{d�
���6%PC�s��|��U?z@Ɂ��"�RC�ɐrVt)鷍�@��f#��I4C�	0Gn\Sm�����6�B�ɣL��1UM��GL���#[*PX2B�I�t�p�' �h�"���	EB%�C�	h�!����e���8uJ��@B�I�:J$%bS�U9I��TɁ.�tpB�I�AZڈ�4��%I`��P�F7lC䉱q��I��mR�
*����R�3C�	n���c�M�(�j]Bţ-kCC�I�&�i��U�M�\	S������B�	eIDI�P��o8&i�t�YSh�B�	=��mU9%�e��f��P0�B�<vk� X�-16�&�QJ	La�C�	�np�r���=� ��b�2��C��4�Lc�E�k����-��C� O�t#�"��!q��18��C�	�&2xx�e�;ݴmp��'b�:C䉫�$�ס�(��؁�%ʪ]�LC䉿0�ak��*#TE2��Ĺg��B� ��p�ՌċVq.��AO� %9�B�)� ����Vt:R�Q�IQ�6���"O��X�bL<^h4��'G�!	l#"O��������y+՞M���a"OD��cM? 8ԸJ!
R�G�<�і"O�xGğ9��q�AiֆC��e��"OFfI�''ep;C�_�0d�mذ"O8t��O�.%����	`&���"O��t��VO`M�a!��m�D��"OY�v��'��	#��ڐ=��e��"O�YVdL9WT.��b�L�6��DA2"O��U��^5胋�G��P��"Oz�:C@6z�H��kՈO��sq"O@�B7$�;�1p�$�`50�"O����.uX�a*��
���Y�"O���K�%��3	��C�j4�%"O�l����t)�4��)�H(�%"O�uPs��;s'��E��:8F8Jv"O`� �������@�K��)@a"O��J*�KJ�P��OΌ#�&��p"Oջi�#u�����L��(YU"OP�QtB_�?rhl�d��?׶��r"O���+�Q�9�pj�s��إ"Ob}�d�X�p���S����|��"O�L���P�c֦$YfjZ�X���1!"O�$�dOX=#ռ�6��Q���f"O޴��Hh�y*��?Lu�HHG"ON�v�o#�ݒ�O,JR`�� "O�t1u-z��@��^����`"O0�A�ѧz�ҝ�&jT?d��"O��3"Ǜ|��X0o�2l%6D��"O���wNpAԽ�c��L1�"OĨz%%�	�c���
/,<"O
�:��֨ouT�7+έ�ƨ���'����0����F=w���B.�e~�:��5D�cQ��d��Iѥ��~. ���1�ɿ���S�h8��x	�L�󯜕xi�qAc��p����ȓ��J�jH$-�I���8.�|�A�� ��/ �`E��OZh@�EQV��Px>�sd�<I�i�}0�ZTN�%��)Kf)F)�������>��T�}�������ĸ�2% S��P��(��gV`��'2Q#C��
`�L�`̓-� [	�'�P�S��]�]G62�Bـ=�ˍy��Y8�	����+_���كm@%�
�60�ʬ� "O�y�V�8�	�p��ֈ_o�l�O��&�3?�$%DFM�Tm\�	BF��V.�k�<�q$K�cO�I�e�� ^:A�u�%@�(a�\���>�@��5I�nm��̍�2����@o���J�&�NR� �'~n����  ܨ*�� �-�l�R�'~�"h�6�V����K�&M����{�E%YN���I��n|���(I#:5h�F'�!�� � �P�.C�N `c7�l�.!R�5�g?Y7eJ(
>,���"���)IHf�<�6F�2B�|+���6UҕfGT�<�"�E�m*0��(ٯF
u(n�W�<i��Ϩe,n�P�D�%����P�<�GB����$@b�Ώo���(4��S�<ᦈ��]�"�����z�J�H�K�M�<��J�_(�H��*���L\�<av`ٛ��@c���M���X�<����]�x�1�]�Э闇7T�Hd�@�+������$ �X�`n<D� j@�Njɾ��"��P����1D���U������F� �K<����*D�P��+b�¸���Z90����,D�� f� ���zQ�p�k
�L6H�0"O,٩��<e8.Dq��ݪ�c"O�)� �y�����a�
~��1��"O���r-�0��-�&`�/��Q"O��c �N';�����$"O؅�T��\&[� G.~�p�"O�p[�hB�Z&a��EN�oƍ��"O4I��g
l'���2��#). �F"O(�� Z�bL�ٷL�$)FВ"Oh�����	��Xy%��	4��h�p"O$5�"�:�qqj^�:�d�@"O<9�rA�w�NDj�	��U����"O�Y� ��	l(#�ǈ�Q0�� "On�˓�Ӛ,�)�DK�0C*��"ON�YmAT���ZM�>���(q"OjUx���A�q��mՏ��gɌ�y&[80��uj$ I,Yz��H�
�0�yB`�m��83�ŏI%�c!(
�y�l��!�JP@���5B��9������y2��"�$�teN�9�����!�yB$J�R�B�aa"ӯL�,uAP�Y��yG8FZ<���Vi?hP ��p�<�F�["���"G�f��+��Bf�<	U��w�Š���|�|���E�<�GHd�4��aJ�3u�$p�S"j�<Q��Z�m��(�#睮�Ľ�S��m�<�Q�ܼ0tڬ��B�<P���K�d�<��ς8D����:{�H�J���g�<��m\:<T<�'C�8���±ǜe�<Y�o��*����M��'�D�<i���aK�٘�I-0�,�6�E�<���O0��Lz�!�.8�2����_z�<��H���L������X��*v�<y�H1k���B+_* >*Y
w��l�<Q��s��e�B)B�"M��� H�d�<	�ށ<ށ��E�a71 %�^e�<y��.除
�w"�T��cIk�<�w�L-|P�<��^{�Ȉa��`�<��YY�z��AH�~�BHIrb�<��ɚ�S�2qR���?D��i !Bb�<Y�Bܡ9AP�A /p��L)G��a�<	ůâm�~*�H%i\q���]�<i!�R7�* )ukOF�Z�x�BV�<Ad"�2��5�����8�N�V�<�� V;z��e�W�k��9����z�<I��ى=��9��B� g�:�J�m�l�<�Xl=68`�5M侭����c�<��
U��(��1J�N��B$�Y�<�JW#U)L�yd�
��9�w�CS�<�'�$�,��sǇ��� �`&�N�<���� CF+ ���@Ұ��r�<�'��2����Lb�X��D�u�<9�!L�R��`wMA�sw���K�H�<!���K�lE����|�d|�uj K�<�U@�$$�B���J	��m(�a�@�<��㕐q��J��
yrn�����}�<yr`��7���q��i�$	��{�<I��S�@d�h�l@�er(H���r�<!�/S������&���Rp%CG�<�n��H�������ɑ @�<�4�'z�@�͆8f��u���<�q�W�U��QF�V9[��
��b�<� +�(��#�D�B �4i�G�<!q���E��M�Q銱2Ѵ5�IZ�<� Vb $R4x�ʳ�̀}2� "Ol8
E�SO�>��"N�;q愑�"O )a�؛��e�5co���1"O��H�+�q2���*St��`"O� 3!R�C�ԙ�F԰1j�R�"O��ՏVN̪��'d9%"O��6��D�L��C�	K��rC"OL�(�i�Ve�0��ސN<�|&"O��aEL2C�DYG[<u)�U�d"OA�6���r�� ���,$�E8f"O8Q�&�^�`k�a7�؇N�L�(�"O�M�g��=4�׊	�`̒q�"O�]Ɂ딂]���v	O'*�  ��"OV�v�ԨZ_a,�ҵj��y�9�i��C?;i�=�dE˸�y�%[�J=��Hs��7M@x��a��y�"Z�N2�+ �_��܊�,V�y2.V��D)�"��Y� �����y�k�����BL8][.=���Ԣ�y�aM(.a����j�=<�T���̓�yҋ��:�,��>q�֩I��Э�yR��)TY��;2i�+u�Db⠘ �y��D6��Y0�Iɨ�&�󐫍��yB疍��p��n�!�K���y���%R6X	��Z�\�����P��y��F�[�*%�V$�UZ�4rUˁ�y�Fn�qI�E��-�g.ڦ�y�ņ�"N�40���K�.h�7&G��yb���&	ހ��Q�vj�A�C���yR%��6�&�9s���RGf��U���y��� ���ђ0/t#4�=�yr�M:�r�QG���'1F�z$gQ��y�;`�T��`��8	� HW��y2�T�vQ���������珯�y�kUe�����4�Q!vf���yD�w��`��E�5q�Ę�F��y��	w	����!��=����y��� ��dK5o��jAHD��y"�U��6�)4�6-��(���yR�ҵi�X�##	/� 0huJ�/�y���#�[5��R�Lk$��:�y���!Qq����.NQ^���V����yr��#��̺7b��b�MAg�:�yk]�$W�%�PGɛ[z�i4���yB�70�vh��X�S�<�;s�Y��y���P��2v���Y��9+R����y�	1	�tA�E�b�阶,Ċ�yB��87�p�Ӣ��e�~��eCL�yb
\�*V�p�ƛe�|P ����yr퐓/?j×�Ց���A���y�C�44, �{�h������y���H�H0����	>L�ѐ�'��D�r��i/P(�F8��P�'�Ir'*��U��d�6����p�'�����2r���	õ L 8�'�n��Uˍ�uUjaj�c��I��<�
�'�^�d��! @�5
ҐF��D�	�'��)�k�hn�s�9Ҩ��'�R�a4!M�QX��AEߝ:�Z���'�2	�n��i���D��Pq{�'p���!Ƭ42gO��K�6]3	�'��)�6 �[�I��Hi�Ztr	�'}�i A�ӽ<�܍R<q��j�'B�xjd�V'h��6镹e霨���	H��X�#*�.�:�BW��r��� 8�z��<;Ԗ�x��%�@M���d'\O��1��4Ϫ�	�#�g�a�v�|��)��8��I�jF�.Z�㥈�,���hOQ>�Hgj�R�q����%(�d�w!�OĢ=E��o�O�TH@�읠���gdÕ�x��'O`�`!K�'~����!y���ʌ}b�)�Y�	��Q����!�,8W�Z�D �{����hX���Iޔ"�.�S +��I��HO�N
Qܓ2q��B�L�C�8b�͟s(޹#J�D�����鎚Mﬀ�������U����[�����Ҙ[��>yϧ�R�1m��<{�p��8�8'�t��d��u �'';<��#��~p�aB��4cs�,����i��G ���)r�B�_�����m?�"�]�"�H�@b ߶9��A{c-9��7�P	I�'5�$�'X� ZR����c�G�pA���%�/�	p@�Ą�S�l!8LhC��*�RI�d��7W�c�L�tĄ�W�qO��#�.A�Bݨ��^�n�D\��<�ĝ}���O��r�
�ޝRG�S {�R���'�|4a�n�1��p�U/O�� c�'�Q�0E{Zw�xm��a֛Y���%�Ӧ@5	��ybKی%/ #P�W&` �˲.ȓ��'Xў�OКL �����,���(�@�8M>�������'�B��C�O6)���fŋ/��Ie��(�d@q#�L$ڠ�2�B�Iy�rU8O���/?� �M2H54�0�F�U2����H�<Y�o��U4 �Ǥ�Q
��IfL�B�<�ҁ2\u�dNL=��SԪ\z�<����bƊVʓm�� ��Xdm!��A�zƄ"vb����wK^��!�џ|�eȠ�G;O�̘:B�I!�$K��\̓An��n���1���u;!�$�.����n֦�r�§���/!�DıRe���\t�Ap��R�r&!�$H�������}|�X�6-]9`!�DBi��qѐ��*}�"��*�k	!�è������$]V`�ՈUo�!�$��p�2ԭě6�I��C3�!�$� �:uI��)��z���8bR!�$�9㚀��
�x[j!���?U0!�Fs)Xkd�۪O�p�%ĝ�'�!�$R�N�]a(�6h}��-B�N�!�DF�@�>�(@�=��h��@!�d�}�0l꓏]�p>(�bY�,!���[�ʝ���&#�
̰񯇾�!򄌖n\���)_�+x���.
W!�%� ���Ts� y0�O)IM!�dP�p����g�L邭�&�=p8!�d� #�>��af���|� ��7m!�0�:rwe�9s����,j�!���[�@����؍z���*���!��M�/�LT��fA�l�h��-[!�څ^�ְ��l�\� ِ�䏿oE!�$���#T���mrm�ED$؄ȓK1v�#�P?�F�iEI�����Y�0�XR�'2���qI�1!G ��w������ۆNϦ��te�#�
��ȓ/a�R�%4^�IQE�M��a��i�:�슀^3tM��͘�U���ȓ"���92BO�)�;6�/lЮхȓ+W
�Ju�E�;�|��A���PA�ȓg�*	s�o_�*�,�i@� \ Р��<��,b�&�%��M�xB��ȓ-�Nm�p��0>@�hѫ9s��l�������e#�@�hqd�(����S�? BdR�ℱ\( 0��aȌ@���"O�s�n�=#��kcCU�b:��B�"O۱�I�$�P �"V^t��"O�	����Z�T����M=���"O޵2N�yNd ��c6�u C"OӀ-��	O�]Q7�R�!Č��"Ob��`��7`���ᅇ�!5@��r"Ova���
J*S7�'HE��AE"O��u��L_��i!�ЬNSj�:�"O�ḷiѹv!�Q�5�	�KY()4"O�T(��%F���/�=財��"O����cTS�����^HߚY�6"O����Ѣ7F��K���&�<���"Oڭ`E'�D@μ���V��<�f"Ozt�D�A��dR��s�$�!�"O�[q��qa�BDʟ(�I��"O�u�$��9t#n�ZTcπK�ص��"On�R�
�Rl[4�&~����"O��K�Z9�0!#bTz����p"O��@`�Z�Hø}��W���I�"OF�yu
�� Hh"sm�?�J�;d"O\4��JUi���o�5E�u�g"O��	��/Ir�#�͸gM�mX�"O2�c�L�di�EC0� $��(�"OF�Y�)�(e0=��%�4X�y�"O8 ��_ a(��Yх�r�e�"O���$ �0��)h�DɝD}"OJ�3e��k贰gnB-.�ƝҀ"O4x��"�U}P�!pΜ&	�f|ȃ"ORu�iT�?�xh �mׁm��1۷"O��c�5���[�,�y�^�"G"O�踃�תw��Y���*v��@��'�ў��bo��N7&XaG�+Pnt�,D����݌Z��j���E�4a��(D��Sw��ej����Ef� $`��%D�x��eW�mj���FD��K�"D��;�)�+��a�r䀋e���U D�T���A�qU�ٶ�B�4umر�3D�p��.ԚZ�吗�")���&
<D��b��߃���i�92"i;D��Bv'�#J B夕1�͢��3D��i���.	�T1���R�i�J��L�<i��@P]3w+=��,�CGs�<��$͜_~�1 ��~�*}[���o�<aFX)i��`zW ��y�f�e�<���q�����O-bY��xB�OL�<�&�N7C����7�̩ >%j@oM�<Q��r��b�Ez��ElJ�<Q�*S�-P��΁g�<b5�	{�<���>'���9�����!�箞l�<1�j�	"��d���Դ�^��
�h�<i�ꃣ<��(Q��%*l@�I�@|�<�B�ԚnҸ��IZ%���F�w�<�`�B�G@\�j@<6ɢ(�m�s�<)��I�z�HkҨ\/������o�<yb+�΄-��薪M�ڤ3�Jo�<J^9plp)p�]-usV�q�g�<�p�2���a�I+";��P'�a�<i��yG�R$'�UjX�"Ǎ�g�<���Se�`İ��E�.�2���_�<���ң4���	�G6�|J�k�W�<�^���@M�Psn=c#{{� �ȓXy" ��µ!~�[��I�O؀��q*zE�bH�sՂi�DN?T�0L��S�? ����` -�� �"=2""Ob<`e��[���۲-R��U)�*O�i�vBr��ٲ6c��qr���'��"��}��k���0��P{�'K�D9��%��,�BÜ�{��9�'�z4�&_?t��Kꋒ\0�@�'&Z`��g<;r�U�Z�O�l���'�D��c1QǺ!04�O�vm��'<�k2�C%2�����-^j[	�'�-*2C�! ��Yb�G"^�,I
�'Ѣ�y�E�.0����!�+E�P��'�x5S�N�]�V|����7��0�'���c����j�ӣ	��*�'����MG'y�`�X�Ż�ꐢ�'� ᇧ1���x�F]�|6��'��<�	D�eD�MZ��.��'�!��N�	� 8ӣ���R�����'<谳�E��)�q����Y���	�'/vp�%o�I,�I�Q@[�U��K�'� i!�&�/3%`[E�A3���'�����5�5��D��V�C�''l�I�Á$�6��aC	x�̝#�'x���%�//�!��`�'8Yk�'�vi"pnH�R�b=�!͈���M?D��gÐ5��u�� �K���h D���S��Q-9t�Xj)>D�̈�U,;��9�j��6�a*�*'D�챴-��z jF��/'�B0K�@/D����I��ڀ� k0P�Ze��$1D�@��눠?�Bhu�T]��r7�+D� q5/�:3��,r��P�	x2���*D�$��`�z���j�D�k[���#D��DK��ިIv$� g)�%��� D��`pȜ?D�45�& �"=|9��-,D�����ؕLD m
G�eܪ�"3�<D�����\��x�P�CY�5��-D��
7�D${n�eQAo��%t�66D�ppD,ڵ} P����	=SLBF�4D��SҠ[�#���lF�d�P�)1D�����S)q6�:jO���4��"/D��0�R�������J<R�!��:D��� �[�@Hg�9L��lCG�%D�4j�i�4hw�R C9EIȔ �"!D��K������ FFҕBt� D���p���1K��'9W��(��<D�����5Eג9��m?�Pm�rA<D�>��`T(.Ui�lՈ%e�C�I�0̐Xr�Eۋ$�����'T�?FB��
�����Z7@�<��	S"G�"B��Q�YE�/1����wxχ�y2��a7��Iš1cR���ND$�y�-^(V���:������e��y⦌�TIT�bR�\�=J"��թ�3�y�!��@���t��.�ĸ4�ۂ�y� �:HK��h5���8�H�Ë��yR�֏�$�%e��4L���c�4�y��K� ����K׎50����Q��y2�Ƀ&�Ha�цW��4�j2�A$�y���7W�R�`pꃁ{���r��y�`�h��
���;���K���yBO/�x��� bU���!.�%�y���	��	qH>`PQo�'�y��:2|$�sΟ�V
�l0`�Z �y��@����w�F�Nb���g
&�y
� ^U��l��d��a2P�&�vq�B"ODX�@b� ˒�����T���"Ov|)\��T�c���>�(�U"O��6��m���WV @"O:d�U,�s�0=8��TduR�Z"O�i�v
«d~!��Jг��FRG�<(@�5➌j��)~�l�1ȍx�<Y�LA�x�^��ۢ'�%�Uz�<q0�X9,�M�R*^�:e�t0Åt�<a2k��>�F���΋m�T���J�<��/��\4T����%I�,���AE�<!$&�5G�Ahb�4��L�E�f�<�� ڸd$�R�L�9*� ���\�<1���6I��ܢ��I�>��|�P�<C�	(>Fv%rPi٧w�"��ͳ9^�B�ɱ1�93!�6-XiejL!0�C�5�V���
9uV�m�a�.��C���֤Ч`�jѲ�Y�M�'bC�ɏZ$(���S%V\´1e�C�ɥj��z�M6����T�{E�B�I�=�ayh�3Tc�%*�#W�6,�B�	�%2DbģO�,/�1(�"T�wAdC�ɑb��}� ^$P��J�?!�C�I+5<v�@���ո����O�'uB�^�2���dK��0��%#�C�/A-��I`h��J\��C
=U��C�	;��@aբ�� ���Т���{�PB�	,h
��7>hQ\]A�X��C�.~��|���1� �q�\��C䉐',� @  �"O8͠"���"ՑG�ݎvw�X��"OVm���
�R��͈ёShj��"O���
�O�>4�(�z���@�"O,�9���+ ��%�q�"�2�Y�"O�1Pǡ�)����H�<*�"O(0)�D p�b�`f�o�Ɲc�"OX�2��EAru���ֹ1���"O�Hs�ɍe�ܽ���Q0b*��"O� f][1o�D��J�E-X��s�"O<�J�+�K СCdE��U�V"O���9gs�h�KK�b	�"O�dZQ*�1<�	Ye���N�{v"O��$3ru����Sܾ�"O�!�C@�S*h�y����a�|��'"O���v�H�k�&��E,�!/Tk"O0u��M�w�L�q�l�m��1u"O��zcH�C?d�+�X)7��H��"O��H�zQb���+�29����w"O�\3��	:y\h���SqD"O�e�㯑�WѸ�
��B�@!t,�"O�Ƀ��-,r�J�	�((�(�۲"O �Ǒ&PA����=�ڸq�"O���㚹`�0De
:O��@�s"O�Dt�C�
�ĲR�X m�.�`u"O���`�K�"��L�N�J��ܰg"OTh� #ݚ-$&y;w⍺YH�]3B"O�UP�j�kz%� �#O&�ّu"Oz���$]Km��RsZ3C�ⱒ�"O�i���Χc`x��HD&&��0CF"On� ���*�!�"^�#��,2"Op�P��ƾ|22�0cb��e��$H2"O�ɻ�V�{,|1���ʏ�T́"O����d@�XZJ:R ���,�b"O�����i[D�+�&K:J��0Kr"O��1���
���Ś�w��""O@I�iƥ���"��AU�-"O�tBU!� =��=�R�B�%_���U"O���5d�>�:֭ڱ���� D��c &Y�.�����[�,�l!��?D�� �ɻq�l}Cp%��v������6D��u��+$6 bk f���`#D����L�j?
��` 2�@�M D�xФ㖣3>�6N�g����a)<D��z�
F�0 %��8h98q�I=D���6�Ȉn��`��Z��c�'D�@Ҡ�D�;ax	;s�O�B9�-��+D�,�QG��#_�-{�C+ޙ��k&D�p���94I�A8U�ͣ{�ڕ�r&+D����BV���ՋH95�5K�(D����,3SR�ABf�<7�H�3��)D���.F�=�*��Oǩ%(2P��&D����I�*]ֈJeF.�N`�$D�\P��z-�؁�P�} �j�F1D��W��#a����1�/"C�]S�J0D�p��<_�^�r�͏�ǂUUf0D�P�g�)%�=JB�;Z�z��tB(D�P���7b�\ �aG#�|I�rB+D�x:���i��#T⏉|n�M��h%D�ģ1*@�*��H�mЅl���'#D���1�h�|2�O�WھŘ�>D�x�턷-Y��@Љ
4}b�CQ,?D��(��5BB���e*T#*H��Z�j#D��oB�6L11$�aEr�a� D�,��ֲ!�h�Dɟ/r�H9r�L?D���%HiӞ�H���%�|4�#D���!m�"{��|�P�ǭQ�h�ypA$D�i%m�.Q�	�B(I>U���Z��&D�p)��0Ql��AbS8!�4:�N$D�ػ��&�։��bN�:fx� �h#D��`�$�gK2 &P��\����>D�|A�Ò���!��P H�С	�$9D��W%�Kά����v���7D�� ]�#��73PP58��ŷN���P�"O�\0�M+��iÈ��e��$)�"Ovu(C��%2�d�S�K�=B8h0"O8�����3p���#.N,Ё�"O\�zǣػ�v�� �X����"O !���|�XAm�:.�����"O<�9�)Hb���X�I�|c�"O��q�ႊOP��*��$o���*�"O���B�@s�c��={�"O���E
��uە�϶�. u"OҴ�@ݏo"��c�e4=�r"OD|�v/��"���������<i�"O��"2�$��D�8<���)�"O���f��l�!O��ɛ�"O���&�M�}��,(` D�2��9�"O�53 �I� z�ܩ/)G�,"O���Ľp]Q0��p昑�Ǉ�P�<1�)�`�d@�'�X񺶭�V�<)��+q������$�@'T�Գ�+�-�p�5"�;F1�9J�a-D��Qf�����(ˁ$�5�7�-D��i�IW X��Y&K#\�`��)D�8k�I\�9��YM!��g�'D���$Ǘq% �cP �5H���c!D�X�t*�SEy#�R8�����@=D�|�«��?clg�К 9��g)9D��	�)B��BG���6}��#��5D��k���V��t�*Bʩ�
7D�T����&-L80�6��7��]A4D��J@��&9��� r N���l2D���5�	_Q���O;9="����3D��PSj[fȁ��H\b蹫T�<D�`K0�L���Ar�b�Z�tS��=D�lHG	P65(|�`g�v��y'�6D�,y�i��~dِ�4��Yy��9D�Њ� R�r�*��H���7D�@�+ &"�v�8���3F0A�� >D�(���7(i���A�=i5}�?D�t!�F�=v��bSІAo��p�;D����ݦg�5����1䨨ǋ%D���@Ҝ\�uz�I]l�D²� D����fL/QW�����.p��q
%D���#J_����6�G\"��L D�h��E�3O���N�T�.�X7M*D�d�5j�}����6k̩]N���&D��͟�P�����15��p�#&D�P2IRF�8�i�']s�H�C�;D�\��#�$
�� 	��Ks�T���%D�H�O�t�ܝ�c�A�+$�D�4##D��(eE�
.$�X�!�'@h۷+<D��ćJ��������:'0�yU'<D�(3�N�MLkF�D ��P��&<D��)�2QYL����1䌈�v�0D��j�+��9$n�4�
|��a1D����J�����[/X�	�Ǝ-D�Ȃ!�آdG�ؐ��4՘����>D�� f��o�:$�U�	j�n���*O����m�|��o��T@��K�"O>���Z=L�LEq�@��cG�-�"O����l̓zϰ���m�J ~z"OR�R� �|�(4���L�^�EH�"O�|��B�Sa��r�F@k���"O�-�ՊL<vQ����@�.�x���"OB�R�)Ӌfj	
v`
�
<�"O� �� i��d�Qx� �J��U��"O���p-Q�1�"�	g���j|-˦"O����iUcP8�N��]"< �"O4�s�!�3C�v|�GL��^$��Ц"ON����:�,��+�a�C"OpQ�TmZ&:���Z�ȑ�6kf�%"O
AP�!^'����"a��2�e"O��0"OR�Q��0Q��b��� "O�i�G�_,wn���$! �b"t�8�"OJ\{�� @�T���À/H4�R"O�1�c,�� ��q��*�<�"O�Ր�F�q�`IU`ɭN��H�"O���2+V7Qn��b ɋo@)�t"O�l�	A[��d�3�;�mj�"O	��KL5�< �EY�\���3*O�JǧE%(}�m�r��
� ti	�'
`ݡsD��sxt�I��� �Xe��'�ƁЃ�E&&� PH�a��vWT|��'~�j�a��26�@��C;|΄�'��U⁄D�<���{�[�$Ef��'��TO��*}-���H4� �'ά�1�(R6��yy��҇��}��'�^�
5;�DAʗ��
H�=2�'ȪA:�Ŝ�θ`1'��xV���5|R a�I9_YHԑ�g:.��هȓm̄��N ^��A�%�&���S>�(�-W� ���4�I�a����ȓz�塥!��l���Q���G>�t�ȓ	���`�.I�M� )	�|$��<���(D�
G�j��u����ȓ�lil�=㌀��$Ì#Ө�ȓH�\���:p��C1$R�:HL��ȓ�E2d'V�4D�|㖪�u�؅�RP>���lԤ/L��
���%�����Y7���BQ�2�2soE��I��&���)�A���apǉ%��ȓh�8���ج_b����Z�~� �ȓ����/͕޺��N�:����ȓ�`Ѐl,*��
؉>��ȓC��RR	�V|���k����l� (��E�-݀@��C�q�(Y�ȓr�֭�G�-X~0$��gY�j�1�ȓ6�8D	�)�4E)
� ��B�%a蕆ȓ<��1s��wJD��b��}|�-�����
��M|i�Y��<�N���'@�m�ϓ(p��B��p_j4C�'�&�)7��@� �*M+!�ک	�'�@���� �
m��I��v���'��@h��[5Tx��U�8м��'uJ)t$��(~�s�%����'K^*��S,~py�Goǋ��M�'���� IKD���g%E-P�0
�'�BY�&䊚~*�z@�;�0d�'8�9$.
��&e�׬��A6�ea�'�-ӓB�
R���hZ,4R�1�'/�����N 8�#Ʉ�s�T���'`��c�g'Ye���@��3ab
�{�'�|}BP��-a����P�P��1
�'O^�r�G �^�	EG�%�
�'x�0�f%�o��-�-=�F�
�'� @��Q�
��3��U�X)*Q
�'Дz��}�2%���P�+|��8�';N5�%�6Q6����''����'ܰy����X�|��	���z���� 8��� ݉^�ȍ�E��1p ��"O�D`��-1�AH�B|z�B�"O���F�6j���ON�h\Hq�G"O!�N�@�8a*3.�>�����`�!	��������㝿b��҄�zS�#>������,U����,�|@!�����6�S�4����~�X�-
�hr�lP���'sўb>ez��ľ�4����(R.���+7?a����)�.Y� ҭ<�~Ti��1��Q����*�$[+7r�Hc�GP�D'�e��H�˓�?Q.Oa�T��=�r�� �;z�l1�2����y�֚pn�X��BR}�㰌�6��'�ўb>u�b�
"ݰ��!#]�	�.�Ð#,?����9��T�T�X�|���Ô0�v�	E�����L�fg
K���
	+[4T��+4��mם5���GQ�d�k �%D�<I7�V�nr �/ۡk>��{A�$�a���Od�-s�W�L�j���"H��O&�=E�4��g�2�'!�%XUr�TE\��y��)�'Yw괺�h>5H�� �z�ԉ��''�ɶ��$#�ĥb�D9������ŏ?�q�D�
:� �6I�\�D�<�(O?�	>��\:I�6}�v �˸�hO>=��OD��9%K� �YdIg��D{���Ś���$LI�	�
E��(&X�=�� ]�����T~�2C�VZT#<����?�)���vn�ex�kנN��uRD/�O8O��Q� �1<m���� �r����|���� �p������5 ��I�SK̭�'��6W�69&��7:B�Irur��w@�@<<Yi2�]�0B�ɑ/d�=(���>6L���a�K�B��!�"O�~�P�i�fЋ *�C䉔IT�!��2o2��-��E�C�I8t��I&��#_�@���މ`^�C�	6}�*Hd�\��Z4�!,�lC�t�l�C�005�q��)2!ZC��k�nm!�N�� p�"8&C�	�-�����3k�
� �"sV C�	&*ŊL���׋ry,�@4/�;]j*B�	�<�v��	ѹ2\�j�E
aB�I�0�+7h̊A��)r�֌)U�C�ɺ�r@���+v[�]��k� h��B�+^q��+Y���BVb_%jӚB�I [i輢wf��R� 
ߢEfB�ɼ[����+W�A�D�Jv��}<*B�	�hn�5�ݟkXD�xg��5��C�4�t;�!�Z���A�eIT�&B�I,��c�E/Mr���#�!30�B�	)E����.F�v�y�E	�{��C��"[��1�-ܕHJ��K[�t�C��
;e�9+�C�;�H80(W�o��C�I
U��*ȝ?2����&���}ۘC䉦Y����gco�!�"�� }dC�I������?z��P@Z� G&C�I'Xr]�kP5AN�(�9��B�|�V�� e��M�L��#vB䉐���r�Iڗ ��
�pU�C�	(� %sǊ�xK�UiJS~�B�I(J������
���Y��.z�B�	�x���d!�3��� �̩-�zB�>i�jȸ6`M�G퀘��ꄠO�B�	��e�`�Y�x)D��"ZB�	yP��J��]�u��0
�jB�ɛj4�0��޶ᠡ�te�6�RB�)� ~������<��i 7�G�}��Hh�"O���w�U;1�P��u�_�)J�K�"O�y�&��;f_6���D��.T�˲"O޼��J�
��7m[�;�%]��yB��@�,�a�Ȧ����j�=�yr߶1�Ѱfdֶ;����S���y�G(A�E��B1�+T�3D(��N
��&"_���Q�ǈ�7g-���ܝ���d<���e5U�\ ��'��a�SD]���T4ZP<��r�p���]�(k��T.{_2L�ȓ<sȨ���Q(tƪeC�$�4ov�0��R�iz��݄8�2��o�2ćȓB����Al��:������Tی]�ȓ��|㳄R,N�V�27��\ԾՅȓD��U�&FP!a��a��+������<�#�vs� ���-N�^���]�кE��a �R�O�%n?�ІȓNK�$�P�< d��R�J�"W���ȓ��{���P`�E�,i�̄�{�L]���ϕ.p��dUTe2��ȓ;���	@��*>FT(	��s�z��J�.�!Ԍ�r���@�V|��M�ȓX�~�%��"���е�L_S���ȓB�L�3�v��(�Uk�>5<p��K�,UjE�۷W8%q�J�2#ڄ��F�r}r̢4)J!i2O�x=~Q��3H���C�T.B *�adK�A�:���t�d����=h��LICH܄P8,x������;��iY���!T�0D�X#Uj� N˼�S�b�IP�q�+2D���LN&b��i 7$k�n�0U�<D���e�
#+�!�U'��&t��P��$D��Rb�ʯt٢�Pu�b�h�v�.D��R�K9$���qe��.-�ġ��!D�,�o�E%�a�3��� �:D��ӁD�pv:ى�Q5wߐC�%D������<�B)z���k*bd���!D���gЋx�JE��*��=9R�K,D�,���'���Z`�`�`��(D�$��OH%Ra��aC��|��P;`�!D�T�D���E(��Rl_@���4�$D�\��&�2��u�qF-=z��fK5D�di�j�V@�ת �t�l 4H3D�(S4�J-k ��c��qKt9U%?D�Tz��I.(�.Uh@܏\���H�i;D�x#�)Q�(�j�:�@�'�1s;D�@c! ��"� ���;W�E�"�.D����QP�I:f��rf$�ZG,D�h�e�>r�\+��ŭl*�R�%D�����,*	��c�bŵ$��y�+$D��R�8Q#���GP�E�-��` D��h�e��Bz����
c��aє'1D��R��ޫ��)����9!bt![^!��Ȩ \� ���� �ʬ`�'D0t!�[>y:^��Kڝ$�XQ	�(�E^!���ta^�*��'�P=a�'K|N!�ѝ7"4��w"��a�(�# �EL�!�=7 >�[&�R'0���G���!�$���!ڤe8�l��$)9S]!��M�S1���O��B�pqS'�/}�!�Ĕ�CܘH�rB�$h��y����T�!�D_5P5f�E�/cz��0j�!�ɶy��郶�խTR��r!�؜h�!�� <m��+�~=BU�M�`H.(��"O��@���w�^��׏���y�e"O�Q�PO�m�4< A�Ag�\�g"O�i�w/��I�6T�b�ÄIl|0R"O&��'��&:bT���2V7@�D"O�$��֫TG�A� ��8Y0xAr"O��Cѫ�h�&�Ц+��""Z�c"ORXbC�¢B��08�8
��A�"O��v�"eӇ*ŵm�
 �"OH��'[�y��H�u,ڡ ����"O$y��Ĝ�)��jS��;�>0s"O>u�� �N�� �-i�Hb�"O���s��Za�ũ��@["O<���!�
����A�'\,��&"O�]�&̷>����ƈl�z@:"O��9�CS'E��	TC�1�2"O�q0N̍4[ڼ�U��7-;�T:�"Of:�j�8ar�� �D85"O>i����/5��b�4~E섒"Ohi��έ}oܨ�'����L��0"O�= Pd��o��`�R<^<�B"O��A�ظ�V���d�.`�m��"O.)ؠ蛺9�(�"�=�t4p�"OP̒G,B�yS4Ea�LD m���� "Oh��C�~}�͑ƥO�:{ Lc�"O,T9a���Whjd�΢l�i�"O~L�3#.eH�I�J��d�=�"O�x�QK~	]�p���e�MI�"O(�Iv�L'4,�`'� ���x�"O� Æ��<>�I�ǙXȰ��1"O"%���%n�`�CdZ ��@!�"O��� �J5y ��Dg ��� "O$��&\�t���K5%E�6p0Y�p"O�����_�\e2�	:;l�ɡe"O��;�Xx	r�J�M��z�q��X�<Y����
�l���dY�s��j�<	'�ԧ7��lK�ێF�p�� `�<�4�V7Q��i���z��q8��QB�<�����ք�dO�S��]8"ȟD�<)�뎒p�*��t��:��Z4L�L�<鱠� ��z"
B��i@�p�<��M�R^<[0X���vj�o�<�c��0=S��[�o����t"U#n�<q�H��R�B.X�6��cF_�<a`�Ȟ6aKt�Ĵx��y��TX�<�c��Gʠ�qf)�-Z���7gC_�<�`\#Hڔi��9T�%�T�<Q5˟� @�`d-Ⱥg\�X�fN�<q6n��5T�1�dML ��a�c�<	��l�*���`�%T �kpI]�<�P��%V���j@�[=Z���Q�V�<�����H{��w~b��p��x�<���=R������!8�)�q�<�W�����2G�Ba � 6̏p�<9�PO�+'Е<hX<?Z�P�"O����(-Y �A�%ŢZ.Vu+@*O�1fM�p&XHam- ��p�
�'�� �Q��i}p�9�K��u�'�:��`L>Lc����K5�~� �'2��ab��%'��iA %��	O��'�Vi�0��Eڭ['[� p���'H"���j�� iND;GG�"%j���'δ���zQ�$�&$���J�p�'7���(A�p(�ö��������� v0QH�s�$�9�59�r�C�"O���C)�bw��H#b��xNM0"O����)�<vv�(G�X|=�-�"O���V��R}�ܑ@*U.t5�y "ON��P&��U���x�V�63��r"O�p�"�T�7�&��(�'I� ؅"Or�� ��/#�Lu�sG������"O lA"N�? �.ei��-���!A"O~ ��V&CF�Ã�)�X��"O��Rw�$=�� DFE" ɨ���"OD$h��.���B�+��9�R"OV���\�G�lL����4[�XD�V"O�-CE�N��渻2�-���"O4�* �(a�l�)�HI P��Q�"OT`��)~դxʱ⟈|�L@ �"O�
�ѐz̠��P�U�7Z�`b"O܉(�iC3}�:|���
[E���"OhA&�*,U������h�HSW"OR�"W��.�P���<q��1�"O��31�ӮZ�����HQNE8B"O��jRb�%E+r(۠2�)�"O�+deG�Ф#�g�*�59�'c�	�4գ0��@Щd���yf_�V��$8&�C)d~فt�(�yB��+/,��t*hyD
���y�(D7B%�xGhY�!,����y���)0�t9� 4t�ȑ3�� �y"aP�A:�p"G��yāѲ�/�y2���5l�A�&G[Y0Mb�T��y��ԗ<�*���ױx��B�2�yrJ�bVe�߈Z޴D�	�y�덧[��AnX�"|�w�y/�x�	��y� ) M��m���?Y�O��~�m��O�,C׆ �2߸�b�݉^�*Qp�i���"��wn�<�K��:G��S�?
P��l��˓G�
A�`����\Rs�D�Mޙ2��-�(Ѹ@�̢	�lP#��)���r�M�֤���y� 
�q�옲�.s,��R���0^v�'�ȱ��� �x�b�'}Ҷi�:�� L^t�Y�aG�H̨Í��*�S�$$
\���b A5jK<8p��Ķ�~2�p���oZG��?!��Wyr���<s�����<A��ɸGCd`R�h�$��d�O�̩Q#�]��D�e�60c�
�bؑL�z�^�0��*tz<YES#Q�8�'@�@5���+R�s"�
���%R��(b�g��Q���y��ަz��SV�;�f�$݃
��v([|H� .UN�x�ǯN,|n�;�&jӂDz��Dn�~a�u �7j� @`��$�@�u�	HX����Gz���#];Z�ҔxA,J	q��F�'�Z6mX���i>%;����M��?��4-��Ya���09[_�~�@т�'��ɛ��'K��'��U(�,^)I�p1"��'{�;	��h6	���ꢇ��_�VE~��Y����#"�T2d��EuN��&!"@}��n#y��� �p�����M#4�i4��u!O�t��b�s	�ś��O��$*�)�x}���7Pt�F�q�QAC̞%�p?I�i z��G�υ<�д3d��3%]���	"~r剕&R<Xxt�K��(�	s�D��(�2�i�����D��a�$��R\��j�H�O��Y�	"i���`v���䘍���ՓV��T���|�]w�"y�/Ȍ`�	�㢇�R��}��O�P� ��N"]S�+q����	��)�J~���DR�������uW	Y}2�ܔ�?���i��7-�O�"}"͒0'R>��R��>�!�1�	A��O��=�N<Q ��}F��r�߮gDn<;�%y�'m6���A%�0�f#AN�Ƀ���;@��L��Ej��	_yB◙#�7�1�X���6���a ��Jt 
37rhoZ(�xMsr�;S�4X��
��$�O!!C�����$Ⱦ^����E)�\I/����ťN�� )�l��9�bU+�^�?�H�O �%Ε�& �i�FP!�E�a���Ҍ*OF�P7X�Pԇ�O��K|�	Ο,�I��m���j.�X���R&1�@	��a���	@���HO��U��]���1��ÑC�0�&�O��nڍ�MS���?����+��+A
w�¼�S��(]��s*�$�9Si�O����O ��ʺ���?y��2L$��ęuaR��#�u
���8R��D � A`�]#��u���R�'|����	�m���㌋�za����.p�x� ų
W �`��
(vm�DG|�'vV���t�? ؐ��H�2S��,���e�3�MC�i�bT����n��?�iq*ͻc�v�"�w��f�!D�lY/�+r��#wi]�Z����̻�`�I
�M���i��O*�D�>��.�< 2  ��     �  �  �   <+  )6  R@  �J  .U  H]  [i  �t  6{  ��  @�  ��  Ȕ  �  K�  ��  ҭ  �  X�  ��  ��  �  ^�  ��  ;�  ��  W�  ��  �  i � � 3 � :! }' �*  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��I�<��!�]*A2'-l�ĵ���@G�<���%.H]�CV�+J��Hg��A��X�?9Q��;� i�;CO"���	YE�<��)�2tN�P3"��Gp�I���h�<��DD�T�rĮ��w����JN�<ف*'1:j�Q�^;x7��E%D��1MM�)<M9$fǭRu�1�`�!D��SwaT:ir��j'[����2 <D�4Bf@��&��-��I��rޔ 2A"6��y��>�ꅁ�dC�l����F��B�	�7&��)q�ΤW���YC��� ��a��h��H���74���9��<��"O���C�x�P3���b�e�7_���I�}[z��Ì��S�.�@�AiC䉋(K � N�AS@Y�3ϗ??��B�I�:JvԂtc�d�*�� �}DԢ>������zp0�CY:XVƜ� �]
9��6�0�c���S�?񄡢�*�o܊ �N�'Df �$�B���'��dEx���ṃ>����h@��Vɇ�Q3�բ�*�a��fË�x�����*�X9if�_�?�����	VBa��G����ME�c��(q�H��h���Z3��
�͇+M�� ���jч�9���p���;���"צGSx.���f<� �ah�� �D(RR�d�b��`�<� )���׊T�@��t�_�SH��"Oz��1D:z����Z�5+����"OVx{"�x�A%_/!`d8�"O��B�%O~&�q�J�.n���"O��+�H
���%�ѽ8G��`�"O�}�'�M�Ĵz���4G�5"O��i@�]ɐ%���T� ��"O��J��ɓ:]Ss��4��Ԋ�"O�e�f*�E���rWf-q�m��'�qO0 �H��^��(@U�gCx�I�<D��1#*	Rp�y�T ɚ#�h�R&,�Iy���'X�� �gE��l��c�:��m��Eֺ��6��g
���7��{%
Ezr�'�=%��*$�C��1:�ԋ	Ó�O�6��?�0%��jP�T]�E�O�z����$�g?q��V&�&l�voȤXW��{%�l�'L1O�b���A�	.0�(Ȉ��V�<�3E��7�y��'P�Q�"�N�	���@�H3��ܸ��Y��G{Zw|F����}�5�oE�z��9��'Ȑ f��6���˔}QfLш�'�xp�hY<l��Qo	f�6��S�'��O�%�mء,��5i�|��x�'�#=E���CR|$i` V�Af�9��AY`�d,�OP��>�:� T � P�aR��'�1O�d�T�F�ct읓O�h3d"O�4*�ҏ�,���k��E������$�S�IۖHn��$�D?���i�l��+!�ߌ5͞�rPI�oӨ!�KZ�p!�d�{��8�ʞ�@ ���f\!���rZp�f�
<f���I��O�!���A���E,��C���E�H�!�D �#J\�3C+�5,(�YaDL�x��}R��83F$�*�i�@�(WhH{n3��e���S�0��p�i�����䂼j8C�.���8��T�Q�10�C��A셭�8������+B�PZ��hO?٣��=Ql���A�$.m��q�UE�<�v�D�kȾ�AsEϋd��u%H�~��4�<�gҪ%�H�cI��p��٫�)�wx�P�)O�����Xi�l1a MPrl���d>�S�i��l=*�j��[��\ʦ�O��Py�:�fM�� F�t�GIM���<���$��C���p��-���0����x�!��8���R�jĞa\l�vo�:}�Ib����j��n1~(���
%_��!V�-�O��O�	� ̻{+R����	=�l�fo�O?A�����T]��|ZgEŷi-cF눇��$�2�Mc�<i0��qc��P��E��m1A�T^�<Q#+W�k��P����6D}R��$�
s?������� [��Q�i����09��d���d,�$(�9H9�G����t����Ci ���Iߟ��u���:!@q�ȅzf镉$�6��'ra~��dv�����ΌO|ty鱈^���OTO��O����pN��7�u��戏Ģh�
�'>�$-G'U
9�1.U!��و��)�t�ʭx?Lj��]�Vd
��E2�yB��,~0��XQ�?��5���y���2M'���A-C�Ԑ�36�p<�.O�O���B���1�z|b]�w�(��"O,yz�b�(!#��J�&�0������'ω���4TlC[�R`	���8t��"O$��!��A����`(S�/�ppx "O"L��^L���!Dn�Y��"O`��#jM%��p�_3>���I�"O� 2��� ��Y�`�#�:a�p����J�O�y��Jވ�B�C(מRqN]��'<:� ��)V=��#!i	Ϥ�-O��Ez���pp�4� *W��.�!�$�
:@�:wE��x#f��w�_�5����?+OEGb�Z�X��9��$���ҊU��0?y�X��L]�zٚ��AV��0��%D����
D�r$�wn�\��Ţb�"��hO�� N�,@����!|m`��1�U3w�B䉁S�0Bd�_0��6T�G5��F{J?���I'C��K�Mߐ\}J�#P	6D��9D�@62�H�)W�
��W���<�}��9O
��oGq�P�E�o`٩�"O��q$�׵B b��6i�+~d���ī����8�	{�'"�Q�`_�T�l��O�
6,��O`㟼����$��t1����5�LT`ӣ�G�����)D��:ť��b9b<�4�1�^9�$�+މ'U����E�	����
҂��m<�����n��:�D@fdj�*�-�DM�%�:���x�	�h���O���z��Z��F1c!>4�@�r��(Oj�[�G��UZ�jI�0Ȫ|�����x��P�NܰǪ�>:t�fD[���?�Q�>�˟�aX>�յc�D�H�A�y� �ȓG^�b�-����W�+,rP�{A�-��ګ�0=ْCR�_1XQ���K"pX<Ta!��m(<�شan��R�� ���	�X۔��=ѝ'��x���P@� !@_3$8��r�+"��?�'��a�4���pL��8"���||:8c�'��1�H �hO�����m
���'�
�27(�D��aGb��g_ A
�'B��{���(��E�g�Y:\~�9��'�4�¢��S˂@4���M�X	�'��pҗ �{�˂�1&F ��'�^�*�#��C��L �D�#U#|�Y�'�޹z��͇˥?�δ
��x�<��"V4�ܔ��<9}���c��s�<��G5*�0  a�NBG���dMXY�<y�G�{���*Gobi�tb�^�<����(��@K���" M��P�CE�<�sÖgdPI���Y��.���[�<�P��>�Iw��64He8��X�<�ce�V[2��!�WK�ۣ#p�<a7��l�Y����L���"o`�<�F3} �X�r@ݺ4��	)AdRG�<�X�9�r�Z#��33�0��'_�<!����E S��UB�ДF�Y�<a�M$O�lA�e� B�YP͉W�<I���0�ZG�7ݔ�;!�AW�<�sl�>O(Ii�C=e��Y�m�O�<�`2/
N�KMŲ^��x��w�<�pG��E�2l�PoG�t��p� ��H�<7�߬)��I�'��P`��
��FA�<�mܪG�~�h�B��~p``�I|�<��I�5?����ݺs�j$ꅏ
u�<��i/H��,Z2JR�#L�P��G�<)�#�obaq+[�M{�����{�<y���:}����S��+�H�O�<����r�>`b�)GHP����o�<�NSs��Q��焏��(Q@��Q�<1�V)5�}굃�`��	1���d�<!���WP��(�T����%oY�<��̀![�����mv� ��R�<ǌ:crJ��̚� ���\M�<�5�C�wO��%d  9�ɐ�q�<� 
`OP({�NT*���G� (�4"OƜ:�"B�a�@�@�'���U"OU����^�9�B��7�P��F"OR����!zѲX�FV�|���"O칫���Ί9Z���8����G�'�r�'�B�'���'�r�'���'�l"�j�8f*� "�ᜳ`�g�'���'8"�'���'i�'Hb�'��`0��Az3�$Ce�T�ij��'�"�'\��'���'�R�'p"�'��|`gJtEp�J�iŪ,ˢ��f�'U��'��'���'B�'���'1�����TVZ�H,�>'�n=[�'���'���'�2�'O��'�R�'���z0�+%�JcP�7�"E���'��'�b�'���'���'��'Ƭ]��e8�~� c���+C�+��'R�'b��'���'�R�'���'u|�k��#�	
w%2���`�'c2�'z��'���'���'r�' {7E^�E����$���8�Br�'}b�'`R�'���'�b�'��'��:@		/h��@7��7m��A7�'���'���'���'R�'���'�UA���<-�:6� w�P���'��'�"�'���'R�'}�'��	�䂨L`P��C��}��;w�'_��'O��'��'v"�'��'QB5��L��)��$J�<�U�7�'�2�';"�'�'P�jӮ�D�O�p�q�e�pQic�^�r}�UӏZGyR�'��)�3?�ѱi�쭣!��c��u��&+��H���^$���榭�Is�i>�I��McR�g�Ԭ[�H�9!+� Qh�cd���'M�Qĵi(��O�RFn�!�������HЧ��� 1z
���EwLd��N9�Iݟ`�'k�>�ñ˻��=�-U*(�$���ٳ�M����y���O�H6=�"�q���%D��0�7�]4wN%�v*ئy�ܴ�y2]�b>9�d�M���\ܣ�%��'� ���DE7(V���^25��OÆIH�t���4�
���MY�l�����]
�L�ʂ���d�<YK>�C�i�C�yB���P���c��,��[įϗH��O��'��7���̓��D�p�<�0)��v\����S��:M����e��b>Q�3e�ٺ���'� :u�C�#r,L�R�ؚ7���2[�̕'���9O�|�P�U%'�\*�I�YL���2O�nZ�K_��c�v�4�Rm�'A�$c}�ŉ'��I��"�1O$Ln�	�MS�N\@�4����&-rv�U7V�țSjǵ_��ɂ�ʞ���TG!ѐ�r��
Tx�鑉�'Ei@�P�L"q�Tp  �� �����E/��ġ�$s�����D}�)�� Jv�`J�(y���rPm��\�t�bu�ɵ �t��B(������և{y[@��/�2,�!Ϝ�G�XX7����4}�s�ſ ƴI�eӍo7f����Q5��y�p��aWhd��M�d�p���n��3�p�D�e��Y��E�[��M8ĻGO�p� DqmR^���djW����#�Qyx�0Q�I�r܎��c'��7�7��O$���O���矬����$X8�{�Q;~)���@#)x&h�'q�D�sb�'�i>��H�R��h
�)@�ވYuH��$�i��5�R a�Z�d�O<�D�����O����O���mݩy�Q�S��#���Zf� ͦ-9f�㟰�'���1�O��O?��T�2�p�T	�+W���uC�%^��6�O:���OV-�5��ߦ���ڟX�����i�	�bB3��]	C��5,�\�iWm�J�O䀩W9O�Sߟ,�I���P#R�}��%���#[�F)ڂ���M���*��@�S�i�"�'�B�'dj��~�jU1w>��S��MJ�ʧ�Ŵ��D�5=�1O����ON�$�<��ɲp*�1�d�,~x���֥��ːR�D�'N�P�@����<��'p�i�)3M����̚'��z���Iܟ��I��t�	i��k����6MH;�`���M4v�.����$0	o�џ���ݟ|�I��'w������+�S��R�-٬&踬�+�yG7M�O����OJ���c�$�&! �6-�O��dK�B�8�d��&Z��S�F��kf�oZ�����ßt�'��������'���̃=&1�r�F�(�d�c�X�YΛ��'F�'cb�� �(6M�O��d�O��i�2�)�P��x�Y��%T$!J¥m�,�'�2�������'��i>7�W}�3w�!������[����'��/��5q�6M�O����O��)�V���S�.�Y���ŀxZ .W�378�'��Zl���'�i>ᦟ�h�fd �H�NQ8�J��x�F��u�i���Cu�z�$�Ol������O���O�Ir�U?u@RlC'v�=�v������Lʟ����h�go>�$?q�s�a��\��P�$r�tH	&K����	ǟ`��3|I�t�ߴ�?Q���?y���?�;k�يE��5s7�)H@0n��Д'3�@Ҙ��I�O0�D�O����O�5ܱ�sD�8@ �A�D������JT�h ߴ�?����?����K?� hۻ0���
}�����z}�h���y��'�"�'�ґ�t��9g�@���V<<�H��4��*<�9dd�|��O���O���O��	ן��wˋ�U�j�w��3.��Į�p����?Y��?9��?��&��� �i'Vq��/�LV�*�B�d ��af{����O���O����<���VH�'~�^,�3�I?q�d��C�Ós`�Q��ir�cCcSR�'��I�6d�E�O|�3�Hf��Q��a��(�pt+�� � ԛ��'��'@�I/l�Lb��r�-������6f� �B�d�����O��R(��!����'���/�!f:шH�(���A[1a�RO�pd�yDx��� ����~o���R�G8,����i�剆S�� ��4#(����� ��d�-k.I�����p���kŃO
�v]���d/$�S�'v�40!��7N�X�[�.$��o͂��4�?I��?���e߉'�	6E0�)���u���rÖ9D`�7-�6Z�"|"���<c���a��a�R킥>�HM;��i2"�'_�	T#npc�d��K?�p/Z�BL�7E�.UNRm��"�i�n%�)�<��?Y�h%,��)��R�$ݠRkI�>���p��iX$�.�lO��$�Ox�Ok�ѐ$U>�iB͠J��q;u�^�tz���2itc���I����iy�b�ET�E�?z��=�2h�?�(\(t-%��O���>�$�<��EחI1㔀\�N�3,J��,)�<9��?�����@-<��e�'6����uN̡X֝ۢL�|��8�'a��':�'`��2C\����j��0<Ֆ����ʚp(z�'�B�'d�S�L�Eۨ��'r�P�J��$��H�JF����i���|�Q�����7����v� �$�#L�a���mo�6�O���<yAc�5��O��O�v��1�Ζ><�)��W'e� �Ң$�d�<Y��L����[1Rt���U�j���0�Ĭ65�VZ�X��/�!�M�RS?����?9��O�hY��I�Q2�ɛ��i�p�i��I��"<�~J��H;,��@�@)=�L��c�����1����M����?q���7�x��'
 u#�/0�$L�2Jэ@��S��~�%L�"|J��l*0�Ѩ�4��h�g�O2���i~��'����Z�O�D�O����3GBm:�H�z���x� G>~��c�|�t0�I��$���	��Rt��a�I
O��)	Ԇû�M�pK~	יxr�'`�|Zcu>��&��V�p��E�m�xa��OP,"3��Ov�$�O���f�!&�c����%�B�a�E�2ya�'"�'��'�I6 -�����&v���E�S�"D����@6�I��(��̟d�'�f�ѶEg>�SJ W<D���ߞP�`C�A$�d�O��O��@�	�'�F�dX�MiZ	݌��$"�O��D�O���<I��W�O��s��NV���%��:����Fi�8�>���<��j�q�_X�ʂ(��4�vI��o}��l�ß���ny�n�(�z�l�$���
�M�n˘Q$��&b_:���d�r�Uy��1�O�Ӧ	������b�.��7٧o�6-�<!ӌ�*˛�-�~r��ꄜ�4+�Y7���+P P�P��oӒ˓��aFx�����sL�܃��0�D�s���MK׫̔3���'��'���&�I�s:�J��/�T1�2$��FM�Ip�4XלGx����O�G�H�7�����5���BOڦE�I������=�^�RK<!��?��(���AfY�>�\��SBx���"�d��j�<q���?���d2�	3U�X����Ԑu"��i`R��3��c����򟠔�5f%X5M������{	�qv����-�1O����O����<�L�H@�臤�K=P� �
��+�V��2�x"�'���'���pyR���q�=HHR(l`L����Y��L[�y2�'���'��	�~�x�ЛO��u�a$��p� ��Ɯ)8|�(:�OZ��O�OX� �t,�'~@�1+�0f�TP��
|�&��O���O:���<9b	F�~��On��+B�K%���	#��eD�]r�.}�(�1�$�<��DZ�j0���g��Ir�;�d�l����Ity���a^�8����R� 7g��O�`0�ܞ>%�q�v�q�yyBHŵ�O�өm�P��`�<SK��:�Fc��6��<��>5�6-�~r���e��hs������BR�m�@��e�V˓|�vFx����2.�t��`N�$SvЖ0}?8Ml�j��4�?����?��'G�'�B�K�H�T$��~��cv�^��7m�1M��"|*��h �Q�I�Bf}�A����Z��i%��'>���WrOv�$�OF��-+3�p@�b
���`_�:I�c�����/��ɟ@��ڟ��M��m)����/	��09V$Π�M���?����x��'�r�|Zc|2͈Ǭ��ds^Y��I�*$�`Գ�O��" �D�O�D�OV˓'�,�1Pd"UO@Ӡ�=��j�FgF�O���=�d�<	�&_�3	sbE�:W������ۚ�ll�<���?y����>}d��'�J0��!|���FK�8���%����F�IHyr#]���dC�=�ޖ��aԮ�I �H�O�D�O���<�6A N��OzDYi#�ŚSV,�Sh�O��ܢ�o���d.��<If�X�Spf��0��Y����ҕ���mZ�����by�(O�?���(���&��C肭d�`��fD�U�4��Z�DyR�P*�O��"w��J��&"gl����<�7M�<�a��\�VM�~����:���X��n϶	V�V�Y�u��<�D�`���B�VUFx��$�X�^B�rb:Y�x����M[� ��;M�f�'���'����)���O�l�^�4ـQ��a�N(����ɪ�n2�S�O�b,� R�����;���VMO�J��}(v�i�r�'���Y5�O��$�OZ��"k��%r3�R�n�H�:R�WPl*����O��d�O�}GB;^���rC
r��I��N�M��Hwph�I<����?�M>�1/~���
̙k� �IU�`�eF~2�'6��'��	TIf8A�*|��UC��\"R�񆇡�ē�?9�����IR(r\{�&�,�T�;��S> {�c�4�Iџ��IZy")ѷ'���S�����d����4���O�kݢ듡?������(O>��)��81�H �R~�(X��[�H��ʟ���VyҀ�(��Fd�4������uNԯP��
}b�nZ��%����	-�u f",vHe���q%7��O��<ѣIR�vىO�b�O%��p��N��@�o��>�D���3�d?�O̐�k�N2H��sB��n���_�,Q�]��Mcd[?a���?%!�O�u��AUgp�Q�U3���R�i���'��}�W�4��'�*qS��>@jhH�2i� ��޴}���1�i��'u��O� O��ē����ވ$�@!
ܕLu�k�4 ��D���Ϙ'��`���R�PU)T�z�)2���h6��O(���O.�1��M�����	ϟ�JA��Gvj��`޺&Lx�cq�ԭ��'�%�y��'2b�'V��3H��`S�qƮǿr>�r�����U54�(��>y�����K���7R%b�a3���%�`.}}�����'��'f�X��ҥ��+gh�2�H$�081��'=a2]�I<a���?9J>i��?��K�� +ʉ)���Ԫ=��	9w����$�O��D�O��\��|�D7�dDp�*�)h��5��,�f�j�X�[�\���p'�X���� ��ҟ�c� K/�y���O�\JD�3@�)��d�O���OJ�94lĭF�S/%��2h�'.����mt}Hݴ�?yL>���?��Ʌ�<9K��u�7+��a�A�PK����q�J�D�Ojʓ�^��ו���'��t����<ժ�GKn%H)�E�A9"DOH���O6�	C��O��O�;">lBt�"�D]8u�$��V�i�I�c<Pͺ�4L��S�����$��n�F0sE�o�"Y��S����'g�/ҡ�yZ�"}��삅}צݨ@��8þ��Fݦ����M����o̟��ӻ�ē�?�`a�"	��
Ѥ�(�0�(�^�����y�|��i�OJ4����'x��g�%2B�Y�Rgڦ��I��x�	�?s�[K<����?��':mz'f� <�<9$& hd���ݴ��nm�]�S���'���'������@XG��|���hӺ���P�}%�h�I��p'��،$�4+�c�Rj����}���Ghi�����O8�d�Or�M�$�-)X��ǨE�7�0��C�=#�ļ�I<Y���?�M>Q��?Y.D��'#T�;� �a��;T�Q����d�O��D�O�˓4�T}�t5���JSc�-x������M^D�x�x��'��'���'u��S��'kj�2ve��K�ʨx�IT�N��0%�>	��?Y����d� ��&>QY�@��X�0lU�K�z�S  .�MC����?I�le�Q�����<YQD�I�/ĭ}�L=���'O[ 7m�O��$�<���Z�\��O���OAD�a�K h��3pf�&ꢈ;d�1���O���������7�T?}R�*�/��(�S�T���Au/o�T�#��h�i���'�?����Ɍ,��u%��o�`y��eX$�6��O��$�M��D$��i��s֮�T�ry���W�I���҆-͔@��ȁ'gX
m%�l��C��q�������I:%)d�G�$gk��,4P�5)s�2a���e�:*�)��C��C��f ���-ӞM�Q���28��H!��� �jP�pnߙ9B����^PhkQ. ���Т�� P�;u�,Fz���.˚k�H���Y.�2%�s��lQ񥗒)	 @S��8~
}QF��CFYy1RK�a���T��i�֏�����JF|u�A���?����?)��F���Of��(D�ޖ"�n��GA9̞�� �E�C֠�L,9�����'u����jޭu��А�
�?9���Q!ϥ>�@s�I!|O�L꓃��*��W����M��N�=ro.�O��X$�J���ś �˥Mn~��P�'X�'=(��M���E��
23y��yB"}�d�OvU�����Iٟ  A��3����1̉�w��@����֟`�I�/��x�Iǟ��I"��Y�)��M����eQ4��gUD����6X�$�U�D���O��kեV) ����K$.�@hƫٟ`�04��E$?_�`�%R��BY0���8k6zAj�{�F���?��i�v7��O��Ƀ��?c1�܋�ᚌb*����<�۴��O���I�P:����<��aɌ�1�az��'r�I��M3F�K�syL�����=?q����C+��V��(F�)N�p5���@�O �=���'����%&ZR���ض,��Q���'"ƃYUB�T>�aJ�h�t�	~F�Ps�NDI�O�0��)��9y�4���J�k䠋�Hn��':���z�ɧ�O�(@�)�E�~��c� �j@��	�'ה���F�pP�9��ȏ)*4d�	ÓHU��� p�6!Ԝe���P-g@Xӷ��`}��'��(3\Ԙ�r��'�r�'��w�$�K���
�d���F8!Oйi���� 8����O�<�a��V�1��'��q����&m{r�s��6}�t�"a��|�lݛU��O��r���7����P�ڴ���L
)�p}��"�"&�p͛����ą El�O�ў���n8]�x�'ŉJ�ش�%�>D�Ļe陋y#R��� C $zK�=8��Ƀ�HO�	�OR˓4�����A4j񒕰1�T���&B�
�p���?!���?Iŷ���O��?���܂x�z�3u` �GO0�!��4���oϒ,�䜰�G#�%A�Ĝ�Q�>B�	�.�8��C^�m�`=HB�A A9�u��
�OPl��	�d�X����{���'��&C�ɖ7!{q�W�7sNi�"�ޏ{�Xb��K�}��4|�P7��O����e݆�@ë��`�z�qd���` �d�O�iە��O���|>�9 ���MѤ)gO��V X�Y��%7�%��@�7tZy�7O���A`���	0��h�Ț�O�����)��p�1b�LH-I�qd���
�_�<�U����'�݊�zK�'Fx &�T 	X�x!n	ϺaP�'�d�3��������	�2���'*�7�6v��1A�I�)��jAL#���Od!�1D�]����ДO��i�d�'iڄ�����R�Ȇ	߉M�
	{4�'9"��Z��M٤*ݫG4�'ד++
�����IR��t�ӆ���g������s��<�D9�W��-���#���7N��mi���C��ZPI>]��늨ZajQ���� @��@�
,}2ï�?���|���ބ	3V=���þQ)�T@S'Q!�y�EC1SF�"�G��M�X���	�0<��I5:I:ic�أ\"�&��t�"4��4�?i���?a���f@x��?1��?ͻ+($BEW�o���AA�܆6��1�r$�:T����tԁ 	��1�I+��Og(�'���;V�� ]8�u��@�@�QH�R�L��E��)(D)����>=�M?E�AfE-8B�.γ|�v���Ge�U3�*�. �D�O��d�3����Y������&�9GJ��o����E�O��Ɠ�h�{C��*N�[��~|D��'��#=��'�?�+ORu{,N&e���m`D�8�g7��ᰁF�O��d�O��Ӻ��?�O�� 㒭H6F�4��!�ϋ~j�Y�ԣ��x�IE-S*��;��H� .`�H�,�z8���'-��3CN1���X�h̤U��P���9�?9��'��E0�J��:������1>$��'F�G�Ul"�;s�U(|�Xy�N*�ɝ<�����4�?���g3�캗ʇN2��&#��Ko�����?I3���?������ s���兕�wz����5~���X���"t92o&S����0�)�0Rׇę]�H��s&P-]�\Jc�I۴TSڕ�(Z���-�Zl�-E�53F��ɖ"�O��d�<�(�J�@��"<a�C#��<����?����Ӻ3쒅B톷~�e��ֲe$!�Ŧ��@	c���bTI!+���C�H�'�����*h�|���O�˧|VM��*=�H��c�l|��P��^;FۀY���?A�C��&5c6�4�T>5�O������/Bب�����n��sH�X�F&ל6���"� `�O�NC�(S��C/Cy 
M���'&�OJUl��M����O�xQR�ǐ�,)��M� ���b�y��'��y�Dݗj��LI��]�!5Υ+P+��0<�I/YN���5v(�u��<�Θ��4�?q��?�`ML bF�J��?Q���?��;1�� y� ��q`v��
�jX9�Ju��� �	�R�z��I����O��'h�0aDL�	��Y(���:�f��b`�q�4 c��k	H]�0*Hn�hg+�|Z��i3T�̻g��K @A�ezP�N�+D��b�|���+�?�}&��S�HL:!ԹRĆ�%�*��6�"D�X:��^"�p�H]:w�ܴ8p!b�d����HO�	=�D
0AK��!KA�6���Ԇ�`B0,����O ���O�Ю;�?q�����!k���v+�=��0��9y��3	�',"\���5_� ��Q��zW���x�h�� ��X#�!F�X����J#j���*��1saʐ�`U���2M�
MNLI񯇅�y�lY�T��@	 �:����^̘'/b�hyTč�M���?�c"���b1�2-�u1&NW,�?��l�����?!�O�Yc��T�;W6� Y��p���d�}�ҭ��J�QI4O�J���oиB"�>�3O�kyr�0�ѡ �( b�a8���"�OZn���dq�r���O�>|���IL��O���3�)�'K�zI��-�hg��� ںn߬	���4<�&`��z�hiâ��/Z��a��?�yR^���3	��MK���?�-�4e!4�O� L��Z8,)���K�M�֏�Ol��S�j36!��dP�{��Ŕ��I�|2��N1z��q�bf�P�e
R��).�̅�!�Y-��e� F�k���"*0�	��_��t��	�?"�.����[,��|@�M�	���S��a7p�� n�T�J�0�:w�8��.Ud��d^[��|իE�r0�ቷ�HOu �#\�*:Z+B.ђX��J�$Ǧ����|�ɕ����mF����I���iޱ���2e���4�-9�����AƜµ끚��p��H��h���%?�.���8c���iB��MJ� GX1�~@2׌���(�5�JVoZ�q�oḑaZ-X�Oi�=���ԩj��1�$�"�P!k���(�M��]�� ���Oq���'�	T<E�,���T��B+u���v��'��{2F+zL�1�(�u�d!�s�ǃ�����e��4���|��'���J,l@vݚCƛ�Y8���kW>=��4xÃ�i����O�d�ODٮ;�?������H�aX�ݢu��&(l�9�/|f���~�����B�2�,R�2(Naat�ɇq�n�hFA��R���G�0E����DfZ�q+�œ�+αZ'�*k��E�ɎS4x�d$�1�@u0g �.ypd(,%��#�Op����:�fEIm�3^eˢ"O�E@R&A�k¨@���,<VX����DӦ�$�Ȉ�i������O����Ǧ2J\���?.D�a���OP�Dޟ�@�$�O�28:MX��&>�x�ݲg��}CI	�,,��"�ʔ�Yb�]BW�5O���r�D��M��"*�La�LV-+U��(�o�L���B"�V��ax�D1�?	��i�`�:�P�N��NP���b���+��<	����<�PN�A4���� �b�c"Ne<A��i�l-�d�\�0���Q�h	r]B�9�'��	�0���޴�?����)(�0�<�p�b���
#��C����O�l���/���w�Gy*�X�'/5j,ڱ)�)�8!!�].Ӡ9�O��#ED��o( �Z�#+����:V����oI�39䕤O��E�'�p�O�mc�H$�D0a��q�NQ#�"O�,�wl��"-ȥ
R,��$��L+q�.��|�鉉V^�e�&ꅔ0�04 A 90���`ݴ�?���?AVc@?M�H����?i��?�;:\$R�@��J}�D #�ȰXdYi�yRū��<��ß�\����=l�g�\�,Y.��+:�4��փ P��J7 �˨̱K>qw ɟ�>�OpmF#O�N	N�RT,��d�[0"O-"S$�$\Zt90"� w��V������S9^�~�j&�����v!/�^̸��U \( �I�����ȟ�b^w2�'��	B!ab�U�� `G�}��l�<wN|4�aO�YЖ�7N����ڑ ���)�!�D6N R��ЊI��$��˚�i�l�E�']���DѰ=# �� -\(bO:1���@!�Ċ4!��)�d& *VF	x�`��1O���>QA�Ȃ"����'Z_����b�2�ޞD��1�	ϟ|���ß��	�|2��>X�� C�����TN�@��.
�j�)f�̂0��x���&��0�4"�8g�I�Kr�h	4�ȴt�6 v)·CA^��J�\�	��ē�h���ȪH���sDX^>��+M������=��ũp�EʡFx��i>��ݴ2�0�h�F֎ >1���Z�"K>!Ҩیڛ��'HRV>izuM�۟h�����E�PE�'e�8%��*���Ʌv>l��	B�S��OZp� ��a��q��,�^�*��>)D�l���Obvt+�!��E9���n�,oݬ�J�<I!j�O�\%��?-J�&t��$�7l�|H��ҶI$D����^�⃎+M�fI�m!O>�Gz��f�X������X�� s�7��O��d�O�D	�o8��D�O����O�N˜�8��G��:K�9��ʹnt��+O1^;�$X��8��Ge+��DV�����Dn#K6�d`��*A�Bs	�~��0�ggעBv�: �f�ӿvq64�6��Qx��ŷ:{{�o͏}��Z�J�Ŧqiܴ�?a�C�?�}�'��@Z*�B<�S��c<vqg�$[(��',��˟���'ߜ�� 5)�.��\�t�2�r�O�0l�M+N>t��?�'��%�3�̈́*�TK��$�L8puԕ>w4����'�'���mݍ�	ǟ�Χs8"4��F��jP6���
 =�� �e	R:J�ɓ7b��i�d �0NC:o�L��Y�b%��^��� �&P�ܹ�iQ�>�H��QK�O��I�a�ލ��4)K��OН�	I+M
���L�4պX�B&ۃ:���-�O6雰nջT�љC&L69�X��'i�'���� ̦%L}����+[V�C�yrG}Ӵ�O`�a���z���'&��`dG�T�0`cV ��d����'f�'ը`	b�'�	�c1;��ԇ!Ĭ0�f��� ����d"�1��ڹ�%�')N��w%A�s;���� ��?q6�]U�2@��'3��,[R8���T��O��lZ��ě�d�����y��lz@ŉ~01O��d(<O��C���% L�dp����&�0	"��g����`���wŏ�c $y�A�%wy��$=O"ʓ0�z��p�i���'T�#�-��V����(J��Q�͔V*����ҟ�0^WT�I�#�
X�{G2O�T��Jݑ@Ġ���o8��n���I%;���p��r��9r��%�'�RI�� ۃq���gG�8""ɦO��1�'�
6MPu�z�S>��ƦT�u6�ضiY��c�@��Cx�LSa!ā5��pXTI�S�`�ƅDu�����2�gy�11 !�	0��P�v���*�8	y��i��'���[�L	r�'N��'�r�w�xU�q��C� �@�Z!G���M[�=&��#ׯ 7}�9:�� �1� ��O$$
��֪R*��q)W< ��9�p�ϻ`@�1c�dе�U�r)�$�d�Ħv�D��L���ϻJ���b􄘛B�l�i�2X�8���i�ʓG��I�i>���J��`�-P��%:	0�����ԡs&n�R�����ڵ�'[�"=ͧ�?�*O�ȑ�˗ 8S�CGB{�`%� +��J��S�E�O����O�����3���?�O��+ti�;>��4,Nj���V-ʂz�PB �Ϋw��{��غUM���c�]�ʜ��Ϛ�1�� �&b��*\�1��� 9�f9:�
��1���4\٨ro�0]�J��#M��hP�47W��'��Ο�?�S��
��˦
L��XЬ�O�<Q0�;+�z8 O��6��aY��M̓EJ�aQ����~�-�OZ,U#f���ȳ���v!�h�O��I���'�����'��>�D-�@��Cf�1��&y��ʙ� �v(ͼ��4bG/:Ѧ���2��O�`U#ۼ"����pɛ�8�����Wx�Ub�lŬd} t!P�F�Yjd����,5��et�6�')�kU�[=�6�b��*WJ���yr�'�y�bQ	���b �BJ�YY���'�xB�n����,�F>�ȳߨ^6Msw*�O~�k������i�"�'� w�T�� *��K[�	��#��>�~5���乲"�O�X� h:}*�6�'pFdI௚�wȡ��D0��OHP"4� Ţ��'�thR��ש,gNq��чY�P�OȔ���'�7��d�SR�E���xrk��13>�;AR|(b�t�	Kx������t���u.�-:��+&OrYDz���z�p�7��`sJ���* 

7��O �$�O�0@p�<��d�O&���O$���	M�<�g�+C��(*V�U� c�$AרJ(J��{�mG*Uٖe�'�Ss�I
!-\dq%�-ˀ��4��N]� �a�i�b�"CT�)�8a�Nś.#�t���q ᣓ
�yǧ�B~�0�ȑ���ܓ �O�=w(�O�̓`���D��¶7K�I����r�d��Or��gO	|`�`���u��u��?9��i>&����f�?��9�ʊ�m��8gɌ(���[��Qޟ���ڟ�����u'�'��0��h�ЏȎP���DV�.:�9�I��4������j ����A?<Oȑ��.c��(���"t�i��R9HmJ�(���� iA/U�Q�҄9ړe�R(E&<:�z�Z��X8t�����<�� �0��G
20�@C�#Y��:��ȓP0�V�@��AH�u���<ᶷi(�'s��ULo�D�D�O<���!�
xaL���G\���%�Or�Dý%�L���O��O��àu\ ��'	�Iq�h���AW�����5nέ0&����O�ۡ	ߤs��`(�(�`�Ӯ�(��D��ڵP�
����P�����F$p:j���{"�8�?�C�x�Jno<`�WEV�jx�Y)�.J&�y�J�V�`A+ʓ:0hn|H�f(�x�#uӮ��BDw�lU��W���y�*�䊏G���m�ןD��b�DN�~Z�k��\k�'	�d�F@H��I�q���'k�a%��|fZ43d�]�>�T>)�O+�1
W�����FP��XN�p�gޔ ���x�j�9+"Z=E�dG8O��1�
%-�-��ڭ���KZ��$��y�J|RI~�"lK?`�e�W͌D�P*�ʂc̓�?�ϓDБ@ ����zh���F%��ɽ�HO����z�dQ� D�6�@�E�ئ��Iş���[#������� �IП<����%��.��	狊�+9�d;t�l�^%Z3��
KǨ��B�C�p!�|�`�>ـ U�|&�7LʑjЄ�! A�:n}�$�#E�V�oH0f��ر��EU�ӥ�M� �h�-{W �/�.�A��Z^j�]�A<��]n�M�)�3�D�H~ε�d�̪P�.����1H�!��̫=�jq!��הY־I�a�E��O��Fz�O��'��E`sEO�?�mQ&GۀN�����Y=(��\���'jb�'��do��Iٟ�ΧN�|�r�c�ʔ��S��xVص���5q$���L]��@�tm��p��� <"�۟z�aC�	���S�.��3V(�Y�&ɕF��q� ��{0�քv�$��k0ܞ�h9�� ?_L8�!$��s���D_֦�H<����?��"�&y�<�2UN	&OjA9�GJ �y2"��M�A
E)� �����=��'YH7-�O:�g+ȥ�R�ir�'-,K%�0%�;1�'��@s�'A(�&��'�Iޗ���B���Ha �'	��wN	1\p\A�`c��(�v��
Ǔ��	�o˕;z����ߟ�0H^�=�"�3w�B������(O�D�@�'c6m�䦵�I�au�ђ�cϔ(�(�
Sg�, |ؖ'A���,�h�uTJ�@���HFDB�I��M�s�G	f�*�+�Ea��Y�uh��<*ODѢɗ������O6˧)7�؋���^4	��Q��摱C�@
��I����?��kP�A���M|~rQ>U�O/��"���,@ʡ���g
}sI�h��d�h��� H;5\`8�ǖyUJmPJ?9	1�m¬X��ٛo�X�P�"}�䝳�?���io���'�'��Dś�t�- ����uۜ�[��ϸ��'����?�$G�%t����� [�x-�2#͙P�axRp�0l�����4�?��hL~��e �r���CTOF=*���'�'��=�O�*�r�'�"�'L� �?
w��U��'6��.�k|~5�K� a�iR1d�b>�Op�Ca�.������ѵ-I��Ѱ�<p�B3L�2�;�3�$	1ben:D�� <���֠8C�b���O�d�=l���Y��I����@��=t�r���ʕːE�Ɠ`���C���8mT]�7d�%l^���'�$#=+�T�ʆeB��ޑ3c�+�"ݠ(s��:�4g�)1���?����?������$�O&�ӉC������v��te,Pr�@���=��T�L~���,�� ���(bF���C�ɍNt4Q�鎗�ƭw��#�4�e��O p���#x�����Rwh����?T,�C��}ߢP3vk�6�"���Q/.ئc��P�}���, &�7��O��Y 7�c3g+�Ȃ�� �$�On�`� �O<�~>�a�O�O�����)
��r\�ep�ˑ�'4z�����D�2�P6A_�y�	Ɓ��p<�C�ş�N<i��\�n�)���T�Z��uQ$K�<Y�j��q�Lz��(F�l1��\K<�G�i=���FlX�E%��bP�1I
�'g*�a��_;�%Ȁ�	/�"
�'4 ˶fYo#��Y!h�--jV�h�'��pA�6v��bE� ���j�'����㚟����>i����'�	Ѵ�T�Uuv��Z�LA�'�>����)�d�Ɂ�Ň�&�
�'�XY��\9dT����f��1
�'�����=$��"�OC�܌�	�'~�L
�l�0 *d� ���r��'E��
��ԲC�+���H��'Vm�M�l�^���A�'?P)b�'{��xs&	�yp�(�AX&4��1	�'SP8�Q���wҐգF�W{�8�ʓU����a�?
��Q��0�
%�ȓ{�Jy���%z,�1
7I@��j��ȓmM�Taf��%���@K�* ���F�q	E�}��8�)�#"^
���{����

oO���"V�C <�ȓb�(�ED�z�Z��%Ϝ}��Ȅȓ+�b�i�e1f*�@�� �M9`̄ȓ
�-�V��Pt(% r��u'���ȓ�81����!e���f�T(d���&t
`�3A�N��I�	r۔��ȓ¢�6c�A�|p3���
L���ȓ'�� F���w/80{B� '�p����&�2�@�K�j��&ǔ(}&e��,���Q��gbb���C�$z����(��xDm�>$�Ő"r�bم�*�����eP=��%"0�H����<4��dI�Wh�9�A�P�����d��r�E2	!&u�@#C0
T��S�? $�C�%�-A�fE�H��Y�A�T�2�0bF$x��d"t"O�%���`}�����3���gn��}G��r�!��JʓA���É�HT"(���Ex��y8ƩN��P�KE7; q�>Q��~���'�x!A &~Հ����� J`D�łW0R�`a�SȊ�HO��	���w�N�F��F�J9H�b�.��0��0.DL⟢�D5AB���$e�p�L#�A�GS��AH[01T�2��M�%�̉P�֬/V�{b�^�L(Dxc1黟|���s�S�U�GT�����e^�7�ɋ������r -C���i%.��(�^��t\GR2�sU��~���'�����C�4��Rh
?/�U8N�h��4>�^a�t$�>��A{f@.��?c�,xt#�57а����)r�1��IN������_M ̓�I1j�ݘFkY�"`j)���	�1���nM���J����wF�$FѼ=���`���E{��I[�xJ�[2B��$�$	S%�%mTZ�s�I	4�F�җ̏a�峠�Z��牧8����NŕKh�����#2�����!���
�.��*.ȹ��s���̹P,�a�EH͊&m��:�i]��	�J�ԭj�N=�����b�葮D�	J��s�U%-��I�H�6�����
�@���A�V��"<y�٫���K�7�N�[��oң<A��ԟ��e�4t�~(��
e(�u�u�Z�PMAc�G�2���<��*%��t�q1ﺁ��ϸLQ6� ��[�6�\���i�"�Gy��	d�����EF\�gF�t⡂eH-���8(`Pw��
�s%LԿY��OPj��B���k�)��<TM�Q�O���.��?���@>j��*�*@+f<	�$�5��1
�a<Y�J�g΃LQ!5��p�f��A�4,O�e�U�\�4|�LI�*:K~QcƟ>��fE:4�����L<�ɔ��p��s�lMx���;.��W�ő |59�Obx�̊J����k�&qД�R,�L�̭�p��j:F�<��1P��V4�F��o۪N��z��2۾Jql4ғg�pԚߴ��O�z���L"w.\,@�D��#. �2k�I�Dȸ��rJ�r	���6O�\O#E�"UCT��\�:�R�j�	Pr-S7@��h�Q��N��� (��OT��e
�!W�|Ɂ��1o��I��F�D�x���L�\.!��	��~�+����u�*%�I<A��x���СR��a!��\yBG�J�	�yH~���	�<zz�O�	���\<E�\�4EW*t�"��eV��O*u�&�4�m*Z�fE��7)f( ��Z�	��x#�n��v0��4E�<X�5�
;/Ң<��:Gm:-b-�O����圼+��m#1��3i�8�/-�p�<�.*��\��g+�	n�(���Ļ
�`�W���^� �}B���  ��Vh?���\}yB�i�v�x@lU�U䲥	T��64i3�'+�� �-]�2&�P��s�@iG��C&v�z���X�4����C��b���	zx��FC�?��D �O�柸u�-�Iψ��q$f�����j�67�'�BUQ�'��ۈB �p n*��*j��q��i����0�԰sZZ��B
'X؛��'��rN[K�����52p�qq�j�"C�|�Hm_��L�{׳iR�R` ��\���EzZw��0��M/=�k,7"��Bo�,��y	��S���p!V�N�	�Fˠ�>ͧ�qO���@$Z���� �k�A��81�O�D�6F\'Bh�(r�'B�,;E�K#Du#�iPP�e������m~%+ற����*\�SSʜq�r��**7���	@;|�
�DdV"&@�,p@E�h ��C���f$`��2't��X����$��y��<Q&�\
�܈EMZ)��	(9�����X��37g�gJ�㟼���?4��p�P鑳� e��}Κ�BQ��/��		�>*�Fw�h�7mΨp����Jt�L�C�0S�CBK���<�S>4UL�A<�X%��F%.W|S�&@�i�1��U"Lq�U�p�!e*�ԛ4T�`�W�Iº�	J�6dpS,"�r\���Ga�\����U@\�(Lؔ�U��E���C8zEDq���ŷW+�))3p�
-
�[�$����(O�����	�/�B��N2�X��Sz�\̓� ��`k��#Ak<����X���(Fހ&�jS6�J#=�̀��'t`i���~Z�Ɲ>g�Y�&�T00�hyp��`�D� �����b� +�Ѻ��+^�O�}k6��cD�s�� ;4�s"ĠB{n�Y2B/Z��yb��}�	�Ot�w"H�I+&���m
�u���`iP'?�����jH����e�5S��9N�z�KX�(��]	j� F��s���S�,L*��}h�R��Ey"Kڹzl��`��C*u��u�ҋ��]�>��*U!W갻���"N)T��M��.��Qp�����҆�W�0�B1q��.jH�<0g[�DEy�*\���,���
2~���XFB�Q��0���2�d��F�H����h�.�!+W$Q�+�4щ҅C�1��3��>a������{%zY"�(R�M@6Ԁ�H7	 �^�m�ˁ.� }�s�T$D�?���]
ExE��bTq�3Č�A:>`�G�X�w\�a���OD��	��6��;|Y�f��6�#�τ<$�(�#�ˇ-�lp�e+1��?�!�ǔ<dX��&4,�}��b�D�
C���?�l@��'1{H` �Lܺ��d
6�>ʓ5!�E�`̺a�IgNe#T�T�'�м�>!Q�t/|�5㖱g�h�;��H��zD՛%��+���Q%��q1A ��~b �
Q��	`y�O�\	���@�~�H�H��!�V�0�� 6k`��b�|��aU��b�w@-��l�1����eR���`� �piU� 8�G�% �8zVBPmyB�?9˔ ���I�9��"�%=��O&Q���ԭYyb<��nW��&1Qt�i����1#_lx�4C��3CL�������Y)Ȧ>ao����<�Ӭ(�7�V�LPݘ(n�M�+g��{C`W�*���N��8��O��<)O�� \:4{~��A�R*Mx8�d���'� ��ǈߣpi���F�
٨5�-O�6-��!lSB.E�$�^��򊋤}����22�B���ԟ�y���n�x��`�	�X5�V�߯ �~M��&��*ɚD�E�+���4�ǔ��g����<%?�ʀ�K� ��aؑeI�S�����DG���dW�eMN��6�3]!2a��"P�-��OXQ����LJ^(K4$<?�!C�Uy�T�#G�~��)�JD��#��<"\-r0MI�C�2QX�LԪx����'�%��?-p4EY�&�N�8��5p�&��pR]��3%��*Y��h���]�y�l�d�9���sS$ߜ7Lc��3�&�\:����:��鹧�=���*P,9�aj$ ��!�G��
A�I�'Np��� #��S&�R0O+dA�a�rgV�1�䖰���ѣ^�� +sn�<� q�Ef�[�Q���'�J��Tb�?|��X��E��@)L� ���;b
���V�A	RJ��$��%&`ʷC�?S���5�O�o��\`���?�S2�+H=�)X���;�Ū�^��,��^P�[��r��.�����-o�5���Cn!n�0q:%�^�(�D�O>�=E�$Gç$�08�K��0�����e�*�� �>��BVg@�I�0���eRG�w�ɹ9������L�U��D����@ʓ�(O��;eqQ��x��'Pg����=z�1Ê�7_�E�k�+}�a٧��P���x�-O�y1�#<��<YQ �
�|
W��!Q7��m�C��̅"n�$�G�
�YE���a�O��0p�6S�����/+"0ۓ.l�&����	�&F��<�4�S}1���Ʀ��Tpi`�cߣ:��k-��?��®��X��Ĩx6���f�Z4�lm��'���@��c�]�S�O�:r��, � �!7O��t�� ����B��t
�
��@XGf���	1�L���SOV��jq/�_K��I,}jy�?�'k�t�� ՏeQ�h���b�8R��$�l1�$�>� a�\+�d��4����Ë�N���g}D�Oo�4�N L�ػ�.͐���Y0D�g�F�t�F�B�ûa0"<� �K�:��@�<>�����K��Hp�	�8 ��.	��;���?7-[9}'D|�����z��;f"X�.�p7픨oU��SU�ǡ�(O�t�T�F�z�(�9�ٹ6���'e[�H�b0�ס� Q��O:�	ғ3�l�D:��-aL
�1䢅�&!���̇8e�O� �%F�"O4�0+�'�Bu�/Oh7mE"qYD���L��%��a��ؗ{��%%��,ۀ�O��SΓ��|Y�oU1����A��*Fy"��t��k�t�b�O�X�N�`�/��X���;�dL�C�$O���^C�U�'I"_�έ�Q�>�R!^r?�Ua��J�hp�1l/�	�b��8��m΅"��A�$[�?�$a*J>A�,K���O�I���O�K��xT� ,k��0���܀�M+s�S
�a�#��?c&C�A�0�D��	���)"C�l�<l�`bٙkD�G2�\�L��'n&����|o&���N՛7���Jv��w�21�\��%(n�����w�0O�rJN�cJ���Ӻ�I��>����(G����X��K�⑐h'�-I��$!A���-�<}2=�W	˲T��@�O |^���/�c쓄�@���"�F�+TH��V�E>����O�1����<�l,S �7$�Iq��dʹg*ɨ�ݏnܱz�����M�ēkh4s���O�](M�ʽ��VW0)�,˥�(O�牼Wʼ�;k0��b��BcV6,ps'��CT5��X{F�kwf4�9	rc_���0�8�I���	���"^�,p��>p>$�'���$�<����ʚ��6�x�'��᳐�ԟ��[aEN��t=�1�D�g�,0')D?	���3�o�[5�L�u��"3B��DB�y��Q���I	T �¶�DIh�����d.�'�v�݇{H�]*�bX֜ʏ�LƯ�Xq6�J�F\Hڄ�� Id�<��ԟ`�����=."� Q`�%z�(�Ɗ?hm��*(R��#=��y�J�U,�բe��{w��rA��"�;���O^����
���'/�Ԡa�Uo.��3@ě>���&�~d�#>���U3;��y�ƯL8P^�řE�\�<IM�J$<�`�C6zn�!v��}y��|r'I-�(�򀃝.]X��%�ȍ�~򅗵J��[�W�pA��,v:2y���J��-����q�Y�]��{��������,(�5q Ԣ�����ʲ��D���<Piߵ%a�}�-��f�����a�!h�y�wG)>����"eY
^�=r�O��%)h�}����`is�W�y�
�3��2SN���v�|D���Q���7��ΐ�%{�Z�����>�ڹ[�hĉ,��7ML�Pp"9@���O��M~��a�[;c��{�/�C$rb��I�� �\�48���/m|���!�D�>������	@T��/�?_��dLu�N���(`�B�ȓ���&���Dt�a��Ӵ1�4%@e��;3�l�@@�	6P�>L�DC"޽1�J~��#-1����O![����T�ď*n¶��!��i0v%�!n �=7�O� �ݓ BѺ2��h)2E6j��hQ��]�m��םd�O�ځz�Dݣp�Ja2�C�?�䔪E��W��<S�6aS�����R�+Q3�8%*d'��|L]�Tb
m�(8p�S��"��9OV���'�)�|�J?�Y�H�i�$��E��H��2D�d:�$Ng7�I� �,��x�B�$D��"���x�:���3�(c� D� 1���c�DQ	�b�Jnԙ�3D� ���҅{�t����2R"8@*P�;D�0�1nP�X��QJ�C=��`��&D�����QHZq�0��	3Ϛ8�':D�H"�!�$K�>eev���U&+�!򤞒W�@����T$y)d(ܵ<�!�F:!a�i��D�9�`�s��p�!�RCP��A�ԖU��AKSǕ��!�D4V�`�Kbcڥ�ڰ� m�A�!�d��l������4J\R��B�'�>E�#�ɯDxDi��p�
���'�6-ҒB�F�БY0��X����'D0PQ��M�B�����cx�]#�'��@��/ wD�X��+qT�Q
�'V�Q�B��Q��� �,X2�	�'�N��F��r��4!����'�kG�
?i�`�3F� �02�'�u�'�Kj������b��)�'���5��++�e�b"��U���!�'��� ��Ko?nt�ҌƶY5�$��'Ђ����C��YQ&\�T_0���'�C �^�F��*&��^���'�T��q�8���;��;+O�c�'�@|y��n�Ρ(3MʮV�~�k�';�`@���_��y�B'<n4��'X9��ʃ�5���q"_�a��z�'��a�(�=+�䙐��$���'x<��a�e���Ӱ��?7f5��'K��S�bEq��S�*�E��'� ��@�dܭjЁʫ�*[�'�(D;��_��7�K�J}q�'�� �O�D5�	&ԋ2�]z	�'Zp�o��;�p��̿s֔�9
�'j�E���׿R�&��1aU�w`�B	�'��p��Lϸ[�
��7pi,j�'�,�@�Г_��Q@	R�;��s�'պ�)�Ɵ�'��i�1�4���'�4a*f�ؖcN��@��
�0���']V��cM����m��L�
$U��'��nQ'y�H�.J����'W>)�C���2��SF���Ф,i�'���	 H> �:�"Q��.���'e|��m
��A�W".<��'bX,� �ՃkT�,���O����'��@�!bG,Z��ʡF�*A޵B�'����B�1��|��Ǘ=#@<��'�@�k�M�-]�U�v��$ ;�'���k��_5��Х��l�
�'u��KL8n�.x9s.2DS	�'���pbC�3x�p)���+���'�J豗���p�`�*IRϪ�c�'w�i��Ă`h��J!E(�4`
�'��=���\�L ��G��KRԜ��'��["�	�z 8ԉ�!�/�����'K�XC�#�2!N�24JW5&����'�j�	�\.{�%��@�o��|��'i�p�$_(@�Y[w�>z��a��'�D�Pf�u?�w�_	�<�;��� �P`p�K�g -���x���"O
1����$O\�ȨVf p���"O8�cV�aB,�0�h�X�"O,�)pÂ�P�8pr�Տ9�|1�a"O�T@B��с�OAϨ���"Ony�v�O���T+�#�)�"O�9V��(-2��J��J7 ��t��"O�)З�Ga��9���ď��Q�"O��6G�e>�[�/��@�����"Of�����r�ӷ�τZOf�p�"O��# &L�,��l�īA
D4j"O�E�i�'6���_)gR�Xy�"O89��)BW0\҈I$a�(�"O&-`��['�Zi���K���"Ov!׫Lu��� 3댺=3x�C"ON�#�
�e
5˄
CL�TQ��"O�t���\�G���EHK�+�P�2�"ON�Q7�ڬj�ʅ��-�JӨHhA"O�������
�V����Њ���"O,D�do�$U�j=����{Ǡܢ3"O m�#��LF���#1#��PS�t��	d�v��o�`���JBk��a�ZB䉁o؈�%�(?��e��'(aB�I(�m�QH�Zp�p$J����C�SEzd�W�5	�LQ�`[�
-�C�	�m�B��.z��t�%KF�=�C�ɊU(z� @�2��k�*+v�C�I�3$�j�b�$dX�HGE�2x�L����;��|�'����b�<odX0��+Y��ȓIΘ����ޛKF\�UF�O8-���"���	�=��e*��HO����ȓ:�؊�`ػ&F�ʷcߎ&qL-�ȓ�(\�c�M�~����mͥrl���U����r�ؘn��e�f� 8Bٰ�ȓQ�����ſ0.������ȓr���Q��@��a�T���1'P��ȓB�-A��ZgN諐�Ȇ3�^<��M��hށ/�\��nD)��=�ȓjCV��1���D�l)�'���D��U�ȓsT���aN��i�����>i��M�ȓT=�8	�lS�&Q)�W�_o��Y�ȓ�  A���m�@pq%�Y�;��$��C�V�
�	J�X�� ����	��T��x��PB��8`�l���&��Ԇȓ>~��
F1�)KԃN�e���ȓ]z�{�B�!K&���+������d�	v/8�4����cf|݄�xI@0�D�B3��Q��/�T���O��Jx�eٳg\�Rp�`��'9�Op	8�,��9��9*p�L�TV�)"�'�!�d��3�<%qFN� V�M�az���]	\��,�4�@�|H��Y���9!�D��:7���d�RP��H�PQ��G{*��4(v'ڣ"�ޭ ����(�rG"O6I�w PO\���K
hs����"Ob���B6sm�["��{r��P�"Oj|��jұgk�lH�KU6zI�,�b"O�aCf�P'Dr�d�F�� �"O�%������4�7j 1�u�"O4 
qM�>�x�"j�:'� �jP"O,��bJ��غ��SU���"O�XI�K���`c�*�A�6��R"Op�K�m��B�"�`��M-k�b�`�"O��V���&P,(��.UҤ���"O� Z�1F�L�@UJ�]!#*h8)�"OJ=%��k�
%(`Νfe��"O:e ���,|� � �o�l��F"O�ݰ�̄\x*T���y��}1�"O��)���V���"?�H��"O� 䈃n�y��(sS�uYP"O�"2��!��KXwHL=��"O��ZS��l��G(C,=2zQ�"O����G�p8���Ѧ��)��KG"O�Š�!B�[߼�ۢgL�F�6$� "O��a�:x@��j�f͙R���!�"ғǈ�� c2�i�J��@ -����D6�S�O ����˂J]�mA���5�x�'7�u��n��B�J��u��u�ع�'�y�6��)HPE��l�5j�����^X�\R6/	�F�^�����Tp"�1D�l������)�$M�8P�w.�O��=E��K"x�V�a�-_�����r� �ў�F}½ih�ЁaEƌJs�� T��9u��)Ȏ{��'�r�Cg�N�B�RHRC!^�z�����'V4���؊j$a���&v���S�'n��g푣(�u��[� �k�'��$З�JW�r��U鄚}9ƥ��'?�&� �AQ$i����i	wK����=�S�O&�L�	�b�᫡.�g���	��hO�=#�i�2]b���=�.l��"O6 '��R��Dq��F��]C�"O�$H��*j��2g�ՒB+�x�%"O��#��)z�i��K�(T�����F{�O��'2���s/F��6�H4)����ʓ	�\�gˎ".��y!��,}2���iʞ�0B�;�ʄ��ҼQ����R�̵��mK��ĥ�$	 h��O��D����%��q��F����G�}�/\=�%!U�*!.X���MX����ňxQ���!�+y&8�'Xa~rO�W�'�	�"_
t
󢁨�yB��
pM��Oš LA�2���yRk�?]&h���#
�z�������y��J���q�N�7( �}괪̙�?9�'�n9�n�j�@Mx���}�(�	�'"�����~�U:�cpl ��'W���+�-U�<P�aW���X��D"�S���B�D�xM��j��(� �C��>�M�QVN�/T��,rΊ/-� ��u$9ғ�p<������%�1n�s��Rr�<�d��֐!�/�"��-u��v�<٣���R#�չ#@'^
h�hţ�J�<ylL�4|BI25L	�E5�Y8��G��H�'-��;DH*2�b|j3�
����H�E{���(U:B�ݰ���3���RÁ]��yBcF!D�d|[�1�4�*�O�����6�S�O�tQ��J$$> XagHZ�=�0���)���=j�z����ԏv9�)I��	a�&��p>y�bܮTA�1�7���F+{����>������<KF(����;8W���6`V2pt��$ƂZQ8���	'|o|�K�*u0�,���'8�h��Dr0M�	L�Pt���	�'2�T��&�q�t����F��Lb�'�r��!1"1�"�!?C���b�)
3,�"	4:�&(΍*��z����y�MO�kf̉�d�.P4ٸ���*�HO����b+v�Ñ�39�ls�H�f"!�DD� s>�#��3?Dl�W	B/tqO�=%?� P��@�2U\U:��)�Pqg"O��@��';4�$�ܣ.y�x��"O|�X��X�6T"���3_��"O�Ī��]Z�r(1��Ȱ_Z̓"O�Y3��Y<7�8�@�	"UQp���"OJ��$L�u;nq�IaA��yRM��]��x&I�)<ܕ�G#M�y�.T�.�6�*C�-6�h���g��y�(=1��"@޴zjti�c����yb�	yVza�BΑ�z>r� �I<�y"�׶0�Π3*�\��,z����y�/�"t@]c�D�"R��Lf���yB��g�V1�6GM&Jn�U�%�� �y�A���y � �B�\8��\ �y�	�?�̴kӃY�@��(�.S;�yюX&L�a�S��Р�3)C��yb&�}&u)wW���{D/�/�y��er0}�!��n�5T��y�,{�x@Q'J�6���Z��ħ�y2Ι2[�$��"+Z����W�y��ë=���h���'��iK���yN_�k�B�J�aQ�����B��y�ʔWkQB�3��i���<�y�gM+s��X��Q���IR�U"�y$�1i�L��c��NXP	���+�y�ʐ+py2���hI'vU���3���y�+�m$�� *߻g��ÇO)�y��թm�x�*"�,[���s
��y"*�e4�-"dI@[=⬘���4�yb+O�5Dj4����bD�R-�9�y�gG:;{|���T�t�������y�ώ)n�����Q؞ɀ��&�yb.�|%����ҞK��UJ�����y�	sx^ysUf <��x/��y�(D
&�=��Oۏ0;����
���y�"a�P�T�4q#���&�?�y�n_�/xt)Y�L�p(���N��y2Ȅ�����g�1j���M�y��T�N�(H��V�g�v(#���y2`�H�����Kæ]���'��,�y"(
"Ԩ��
m���b**�yrhĺd:���Z��@�'���y��G�l�.ت��̳N�Խ۶��yr�t�H�*����A��'��yF��~czL" ␰	e��c&�ұ�y�nI�1����J
�z��1ǋ��y�72B���I='P�k�����y�I/+R������||�l�`G
�y�gB��LE8J�yV�]R�D��y���+�Z���{n�����H	�y2&_|��B��_uĊQb�dY�y" ��zE4�;f�rf� p`�7�y�1[
��f#(W�4�b�8�y��J2\�1pׯ�<�p���Q�yb�ޘwPM�e�\	�(�#���y�Eخ!԰�Q�79��R�HR�y���,�Z!�a�@����4냛�y��++�b�r��¾����yb(DV~f�����s]�,��ݝ�yr��B��Pn
<s'��HL��y2��x,�a�C����mH+�y�$<\;�8��h��^�D�hA�+�y2�F��xv��W�XԨ�Z��y"�ұ^�LM�g�3V� ��b��y
� �qa�M���0��^�a�t�"O��Q��߫&���`�"�7ad�e��"O���G e��liG� F���T"Od�1pI�m-�0�UJz��AC"OhiPb�ˏS�<Q�&=�bJ�"OD�`�-R)h��LjŘ�x�PE�r"OiF�	YM�t�dA�l�ޤ{�"Ou��A(|��0�N�$Cd�"O�C���
)�mY��V�[b�T37"O�h��6���cu�� K���"O����ۼw�sF�L7x�#"O �� �����Ť�14F<�Xb"Or���]�~,�����H0��"O��"�BL�}95��qEL�;2"OV��%�V�m��2qVMB"OvP �Q��a���$�q"Oȑ�ӧ̗cƅ��Ⱥ ���Y�"O��3q$��{��8���J�U���	"O�m�C(6�L@�fE"�"O�}4h�i���h�X1;����Q"O I���&�fU���N�g�*��"O�I
Gc��8�P,ㄥ�fi���g"Ojy�� �:3��R�N6]�,(��"O��dKPZK��ӌ�?��Q1"Ob��O2p�RUY�LF�;"OFLXЀC&K~>u
�	�3?�
!	"OF����FZ�L9�cF��d�1J�"O�����'d�d��ǆ_fh�%"O�QB���V����[�����"O*!��@:�fZ@AQ)d��PB�"O�k�D��5Sb�EW�4����"O�07�AQ��� j��s`��r"O)Ѯ�5i=�5�r�Ǆ*]>X� "O��!��6Uy �^��T�7"OrqY樑:`��=b��P������"O���k�G6��B҃��d��U"O�=��5�>`�LV�Ń"O
�{��ɱk���ڃ��
��*�"O��˔o�x		"���~��4"O��P�m$�J��8u���"O�A��d��S'Tm�A�V�IO*	��"O����C�Bx���?$f�@�"Or���cˁG�T S�3�>
U"Ob`d@C�|�����/V�7VE�&"O��3E�*�����;"����B"O�1�׶-���TdΕ	 ��ң"O:�pѫ�#���Z��M%P`��!"OB8�#�Z2��@CeV�N�L=ѐ"O4`��������E�Z����"O
@�6,��t�S��� ;��}�"O<�R@ζ�����ϊix^��"O�ԡ���	 �)wnJ���5��"O�i��`�-aB�:NIb� �"O�r�O�b�	Ƃ[������"O܄P��ZR:�&�I�w��T(�"O.�3%c�rN�-rFAG�6�2ЊC"O��C����2*�jŪ	�����"O��S����|�k��:j*4�%"O�-��)�6'59��ѿj���"O�����&l�ksH^@���"O�h��vhP�����/\�,���"O���1m�<��IP��9Z�f(x�"O�C�K�-��� �N!�<<�4"O8(8����`������8�c"O� @Hڕ�5By�l��	�k��"O:���$U*}�Jc�)��Yg�� "O8�k#��6x
5 dHQ8A=���U"O�]��EDvV��C1kR�p�W"O����C$~�] �e�O�d�q5"O<�I����8���9RD�(x"px6"O$�XcbкLa0����M�e��z""O>\�I�~��c5C�X��)�"O��wLR[�~�أ�T�A��0"Of�2)Ɵ���d��Bq�0�3"O��RD�cu�|��P6iY��"O�i;�~�@0e�uSL�2"O�@@`��5]�� ��k�
��"Oʘ[BEN��5:�t�D�rC"O\�� b�,�8-�6'08dT$c�"OT1Tϊ.p��z�/d���B"O$�!q�A�-�@��b��wIHr"O�����.M��'hLx�
6"O��Zc�s�59TFؼt8 ��"O|D���<� �I��-!^:�"O\Q�O�1o���A�2"�!B"O�ٖ�'=�>rÔ�o�R V"O�,�rn��[�Buy��\�vj�"O�PV��7w�*L�㪟�(����"OV��&W�X�:y)vD0y�ވ
"O줁D�j鑖"�#q�r��"Oj�r��Y�EX��($��2p��%"O2�Y�.ѿ`JZ���ݱS��h%"O��,@5tM*��H��e��"O^��3�Ξ|�K���t��"O��"�S!�ZT���@��8��"O�h��[�"/��*�
�9��Â"O��X��"��d�p	�5�|�qR"O|m��#�>\��pPH@ �6��"OD�:�.��p3z����M�04"O�1����MX�(p���-�죓"Ozx��R�-T�*�ƅ!w-r}P5"O��p1 ����i%;$:B}*"O����$����d 7S18P�"O�͠��e��̒a ��X1Z���"O��h�m�442$���O�hC��["Ol���<,�2��% aQ�u"OBbA�
7Q� ���K�kYV�� "O�A���23���K��-IK����"OX��[QN�L����0.,U��"O�4�DX�zmD ���>�a"O��S_��`	c�.W'v�8t��"Oج*v�a�%�d��}�J���"O�١g�U�"{1��l���c�"O$�*ӆǡ_�D:5kˁ%���t"O 0#���*JOH�*�
��
7"Of����'P�> y�+H&D�"O � ���t*��RF��(.�!z1"O����%ִwʦ���˻DƚH�"O`aX¨�?���9���^��T*�"O	Q�EG'u��$�����"Ob�sg�Z'D�[C���]�Z���"O���#l�Zq!!I**��p"O���!�7A��:a�?����7"O@�6흏'���um�~��[�"OB�F/��M�.���n�$���"OX1y��T�؂ ��D& ���T"O\��REW�9$  ʣ�-sZ�8�"OZ-�0)״XC�u�ӣ3dt���"O� &�)����6#���-N�TpE"Oi���9V��A�C�1=J��+G"O�!p�j�*P��������Ҵ8�"O~�B��~8:U���݃D�֭��"O���� �3T��:��8�Å�"OT8R���8� 85"'�d��2"O�I "�Q,�l���B7	�h��w"Ov�
������KsR�s"OP8�bI�>�0VC�Fi:�h6"O"�A�X�o34�S)hTB�"Ox���(M� �dNL�u��4[�"O����(ߺf�<�(Ս¼5!�Ph�"O��ڰ�B�BZju��+��h�ܣ�"ORY��Ϲkvn���ٞv�D��5"OF��Be_�T���F�X � %"O��;B�'1E�E� @��J�cv"O�D�d@��<�T��Ѯ��D�P�"O\y��&��l:�^
=ɂ�!#"O� ��MЃrF&PSP�F.���"O*�T��:G��jj+]����5"O��j#$T�6��!�V�+�"O
y�V�ظ(f�ysfBM���pU"Or��D�@.k�)�cc�
Q�2"O]Z��נK���D"P��n	Ɇ"O���ƪ%a.d)g��2���@�"O:5+j;��x&�y;���B"OB�$T[ԾP�G��:y�hA9Q"O~l+�E_0/Q��bC.�1{,�d"O�,�Fۣ���(���^o��9'"O�M�bh��,��9�pŃ�2z8�U*Or� @��j  ,�񪍵ۚ�S�'��1!��v��E#� Y��p��"O踁��.�r�C�i���R��'D��aG�]� �4�0���ZmX嫷�2D���ԧP�bV����0hd���F1D� ��O8�$c"��4�B���-D�p�VBWQ�l9�̈  ��e�+D���'�Q�@��{�郯=���+D����새7fN�R5H0��L:3e*D�0��#$��X�� �`N4�Zd�(D�xH"�5]�j,�#�	P�6�A��;D� Y���x:��I��xB!%D�$Y$�
��R��U�(��E#&D��!�g_26��3J.Wڜ�"	&D�("5,o)#FiK6��c�eB_ơ�d��9h����.�
M��P��y2�G(`n��L)z�p��7�T"�y���+<z�`���p��i2GJ�<�y��ۖ:SNdB�元��;�W��y�M�/R��1����7�`%iL�y2���Wo�q��	��J��Pb&�y��Jk�V`�uaWx�l��n��y��z	"�(�,,$o��pE�
�y�B��8H���ͮy:�R��3�y�*C")I0��M�1.�B4�$ ���yrB��Z�x����&w�:������y�燀:gx$�ek��|(N����yrHξG�ɚ�MN�qaV="�ɴ�yb�[����ޕ^�V��b�yb��^f�(*5Ä#S��"�,��y�jѬ^�dx�1�%+:��A薫�y�P�uU�ݠ��5.<�VK��yҊ�5�l��׬쨵ؖ�?�y"gQ	��Y���΃z'�hv���y
� ���ӊ�2j��$Kdg-y��h��"O��@4��l��3'`�KWlL��"O��8��,T~5���9-�"O��'u�N����9H2���"O�$�7ł������C�[L"Q��"O�B�G��o��Xz'A�.V�<q�"OpL�M�G�E��a��>^|T	�"O��*DE/'����f�.TP��0"Oz%[P�ӮR�
%��g��̅�"O| ���B��Z�k$�-+���"O~X���թff�3��5��"O䑓 �1(. ��s+G�<��-1�"O:��(�U�u��U+Xz�y�"O�l�TF�qTͱ��T0j�<�'"O�`��,�Iש�jsVxR�"O�PSv+��\��a�T��"\đ�"O*����?)�@	ؠY��9�"O�5�ե��oJ^I9�	֥ul��(�"O���@�`�*�ƿjH��"O$�1 ��g�p���I�<����"O�!����@FHH;�E����"O� 2Ѧ�=:�&8�d��.�PH�"O*XC��F�>�"�p#)I��k"ON���k��q��Bra/3V�yhd"O�:V��*qu<��t	O���A&"Oġ�!k��hmjwG�x�v虐"O�Āe�6o���M_����"�"O`钢�EgJj8H �V��ؙq "O��YV$��>:�qxpLW,5R`��"OpUX�g��X���XP��ũ`"O��X�G�h2�Y�s�ۘ=ݔYI"O@����*U��Mz��$P3"	�Q"OT8!K�g~ٱ��	G�Ј�"O>T��C��0l�h���F�Rl�9e"O�XS�߃= �yu+�1}�A"O4y3�O9ǀ`��Ț(%2�V"O:���C =CA�(@5I)	��Ɂ"O.U�#EuP�j5"�&s�L��R"O���`o�-��b{�̉#�"O����@̀x��i�w��g=��1 "O�Lq��0��ƀ�
sG����"O�CQ�0隈���D1�F"O���䂕�c1�R�
�Q��"O��y�l@aŖ�B��"Heޅ�C"O���T+1�f�RΔd(J�y�"O��y5�*X"�B4:�"Oz�ۣ#D_HT�a�H�! �q"O�`"� ޘgVI`�@��i�0�"O�����_:�ֹ���\���Ͱ�"OKR� ��,��[�Q2B��"O�a� h	�6�L}��D�"6�"O���7�+�����S�����"OX��#ʱ^��eJ�L7p��"Ol�ӵ�/C:��*b�ȣjY�Q"O������y�,���J���"O�)k���=W��X�&�ډ)=���S"O�A�c͝8����cL�N��#"O�A�D���PB��A�LϸCL`�"OU�%DS; �D��?fƾ$Hs"O>ԡh��3���R���X�p��"O����/"!� ���GL���"OY���4]��aw�W=ȑ�"O��uI�,L�b(+���&�0B�"O���X	A��p��N�5n�S�"O� ,y"�I@�v߲H�c�Ծ]�6�Y'"O�%+��[�a��x�'�ܡ�~��"O���c&��C;4��wꕆ�b���"O`���'l�VȺ��ޠ��|;A"Op"�L��G��ܺ`gG��|�"O���.�8^6I���Q1F�X�BA"O"�إ��=0�8�ӦC[4JA"�"O��Z�͑�t�a�A7Z0�k�"O����oU*="`�c�Ś##b8�"O�()d�P�t��\��@�	[����"O�!A�슀�@	��	GB�X��g"Ov�A��B�q�2x�"�V���a�"Op���˓�)P�4�Bhy>��"O���wH��h�p9�#�B�fẍ�3"Ol�#�˙�&X[ƤQ'e�,�w"O|�3D��&��pn��]��$3�"Ol�:F��%7u��1WM��Ui\���"O���d�eg:y�u�d���T"Oj�ʥ	6_�f|J��ߑa�HC�"O$1��h�y>jL�E�VL�E�@"O:Ekq/��Kᖨ��C�}X��G�<��D��a`�� �:�Vi�2(_T�<ac� �&԰��ө�%C$Xh@o�D�<!�a��W�(��&֗���K�l�U�<)�i�$�+�(�H_�H�E�FS�<c";DN ��EX'�� u�'T�ؙf�0F�Q b� 8#�i$D�X��d 
9��A�D=g"��á D���P3�
	#r��{����-?D��`�C<�X�;�gL�� � 8D�l��\�Tv�4�����'dx�p"D�$vj,ΔTy'�D�W[H�:�$D��Ӯ�3�`������n�� D��acKNq{���[�`�H��WG<D������n��F��+>I��>D���U���R�(����3�����>D�8��5u�ѡ���8�d���9D�|`��ɜE����b�b��F2D���28a��9y�:B���hV�.D�@B6	�	vl }Af��6x���*D�<�� L!h$3�JT	?�\��wi*D�d���Q�24���L_2���t�;D��g�N*�V�-���$�8D���6��a��)�!�$7D�ؠ1��H�z�9�(C�.�D5�4D�����V�R+!/�F>}c J/D�0���W'T��a�ą9�%;D�xW{���{��95�M�9D�4 ��Ėw|�L���F {h|Cь#D�<���۞g���*��,R�*8�6�4D������!\b�	CJ�(���=D�@[c� �<���T :j@պp;D���dH��D�C�^PB���:D��C���vc�ma����=D�H�1��y�t��Â��Q�d9�V�6D�L`a�TY[&E�54ah�3D���+˨{�,��� (��@�k,D�����R(���*�?L���q�+D�@1f�-� j��U3#�x��'D����'9�e�V�����ү2D�X���Y�|��f'�Ak��1�/D��Bda(\|�H5�4v7����"D�hY'�->�"%!̖6�.p��>D�@8���rNb�Ƣ-@2��ag;D�� �$2��ມ[�Q�����S"O I�P� !f�(�*`/X�j�ʜq�"O�\Z�=qpXS�'�H����t"OD�Ƥ�`Z�����T>��xP"O$�ĒT�j�k��)�\"O>�Ӕ��>����_�M�X#�"O @ ����X���$����"O��#�ː�?c�yaփ�F�XP�!"O�tÄ�#g�6@��\�:`(&"O�<"�/1	b���1�F:x���"O�a2�+Z��$���b	�a��i��"Oj<�S�^�F`��Ƃ�t�"O�=s�)G-ݜ�g�ܕUK>���"Oj��s$��l��eDYX�"O��Y�������ǿP�i�"Oz���E�m�D��e,��lo�峐"O�)K�?Y6|�TK'{��'"O��Qn@A���ǩ۽Mt�y#�"O<�X�F��<�ZlC2銉sZ����"Or�VO�.@��0f)A�UF�j�"OQI�G _��आ^�#;��B"OH�SQ�G�����ԍw��9�"O��7��� ɑ�C��SfE�T"O�jW`B�l�4�0�#�0t�գ�"O�}�l��r��, �O��u!ƕ8S"O�b���I��UAuV<��"O�9c�+�(%5~pB��y�s"OJ�r�aH*S`�lH#C��W�5�S"O`j��׷�,�1�@��~�s�"O4h���#4&�<�wBL�d�T��r"O�Y��^�kw��"�ì<҈̹�"Oz���?v9�HX���vk��
�"OX��5jnM��X+/L�|y$"Om��Em!2����I;mҬ&"O���G)�:M��dˈE	�`�c"O�ũÜ�G�,�	7��?1��X�"OX��N�@}�Cː"��u�5"O�	0)K��@���F2�|��"O�Ah�%M�uRb�ˑ�A���0�"O,@��n�	JД��t�EL�e�!"Ou�# �{�V��c�6,�h`"O����M�Kv�����U�I���;�"OB���,�f��D�A-��u"O\�[f�: *���ׅŘ0�0Xkv"OBI�� �9(�$Q�t�Q� �Dh�"O�:3�^8cՊ��V���&ͻ�"O��"��#}��Ad%A� �x�C�"O,|�gmۦzC�1�Å,��e�(D�ds�����:`�f��:t
��j!D�<��)��)P�(7�ݥ���qU?D���0k (�,pa�i��{T����=D�THf�!);2P��� @�L���:D���Bm<(�H��Y����y.%D��Q�G/OF��f`�sg��-D���UF�q�����ԟ�|-
g�%D��3�n�!M�<���B�n����'D�����Ø;rї)928���'"D�,P���3�,�"�*ה!P���?D�d)֯�SY��Q���$p[��>D���"�/���`��1,ڐܛ"�'D����$H�X(
���'T+C?����/!D������r�.T�3�� ��(s�  D��a�2��`{3�S�D��-k5�<D��SV"�4U8���bnАfͰ��A�9D�� $�͇R�8L�4�ںHȆ�h6"O���d%z���� Q��9z�"O���cR6��4��$�*9��lbC"O�E�W�L�rT�&��!��-b"O��1��Q:5�x��`T�x�	q"Oa�C Y,�Eϋ�L<�PX"OL(���s��� � jݺb"O´B �,�P6����,Pa"O~8��Q1y�Hs��3�
\�A"O$Pi�➤M��PD�I�2p��"O� )���Gi��ĕ-�����"O�iX��̭:W\A�ǠO*�J�""O��X�	��j�]:g�_�[���!s"O����>� -����?a�:%�G"O	r�L �
��7f�$5�,M�E"O�Ⲃ\�w$�<��K�,��p#"O��C�KW��HRj��Z��Ց0"O�x��^��6	�-jqu�%"O8�C3���0p��g	�f-��"O�!qf�)'�v%��A4�"O��Y��_�_ ���P�^��@ W"O�����C!}�䩊�X��"O�lۂ��^���c�I�1� ժ�"O��CdM;nz4� �ܑQ��hY"O�3V����ICjJ�`��%��"O�q�ڂhx6�"�U}�\�J2"O �`j͹�D1Ch��S�P��"OZ��C	�_�ڥz��2$��q�"OP�G�D<o*��j!ݐ6���"O�釐,I��CA�Oj�q�s"O|���$�$�!��8��1A"O����c3 ��#�)pc�kק/D��X�K&)9) g�y��i��o#D����A�!t�(JU�ƚF���F�"D�|0'�̮i������E������
?D��Ҏ�6?����aD�oV�]�e�/D�d��)�c����*C�Fd|�B�-D�4��_�|�4��u�35W�8�+D�8�c�ӚtIJUAC�>�d��(D���ğ7*��h7�ϸ=��XP�;D� �M
5�x���j�|țs�;D�䘕	Z�(�
6���*�t�p@�5D��C� #!ޜѲ*D�)��z�.D�|4Eԃ�A�a$���F=��`8D�
G.��H�ʶO���̨�.!D�<���	q�D��ϔ7�p���1D��P)�T�&�&iv���W�"D�X��W!$��Y���;,r`��R�-D���U�),[0�	1�Z���0D�@R��W�����N��Y�dq�<D�|�V�!|nbı��[������&D��sm�yNJdKw*٢��9�W8D�k#���H"�(�	�J�F��5D������dqZ�I��x$x�2D�,@ ��5IW��x"�C�+
H����.D��8F*LB� 4���S��j�u*O
�V��e�'*��>�B�"O�9j��d?L	��NH)z� �F"Of�9�~�px�M�5D�tI0"Oz) c0���+ďM�(�*W"O���X�j����g��z���"O,��GI=>�J1A�GױY�,��Q"Oڜ��DD��D0���_��\۰"O|�	���)��0"�J4,�(�p�"O� l��Owj�؁���&�6D�3"O��0�F�=�z��@�FB���"OF��wgzYx��}=R��"O�p�9��T���M&/J8��"OFL� ��-����4��4O2��"Oxd���ÿ%34ڧ���+��@�"O`U���+f����Y3���"O�@�fQ�/!(�6�A�GR��1"O\т_��p�*�+x̱8B�ş�y2�,��˒�S��n<r��8�y"��4�I'�1a=Θ:��X��yb�R���Ɩ(%�d|�,ȓ�yB�ƛax�� �l0R,K�P>�yb�8>��EA5bCDMأNê�y�^�6����J�"ٌ���HH�<A���?�d���-N�4�(SX�<aE��;_T �u�ғ}Ֆia��LU�<�DkJ�f׌eڣ��s_n-I�dQ�<Q�,F�[L>)���X���`2�J�<�Sl��-��Sw��I� � D�<I�@=5I�qJ�A_47J�I���@�<��G؎|���Q�mV�lʪU��d�p�<1���@�����1D�����d�<4C�x�l�g�Ѫ(�4}3�LUd�<��H��lp�q�7D�7b���WW�<��bG�{�F}�*��=���EH�<1���5a�'�JT�i�OC�<�b �6X��� rLI�"��U�g#AB�<��d�58����4���_��Hs	~�<���Gv<M�K�F�z<�!�
O�<i���,JE!�n0P�y�dJ�<q���,"`�`%�x`��H�G�`�<�ՌK���#ѣw䚘бN\^�<y�%���8А"h4}�N\��h�\�<)`%�='�c e��MDIh@�p�<�g"R6(ؐ6�ަ&E|��&�e�<��b�Elp���L��6�V]k��L^�<��I5r
MS�
ɭwV�y�G@�<���@�\bFyWJK*'iܐ��aYr�<����k.��s@B��b=X�s框t�<a�O�@V P���̲6��Q��f�<�R��[M
�a�C�?���gD�_�<EI��k;��J6P��Hb��g�<��JՐw��넍R)G�d8��l�<�e��9��n�&d���9�e�<���5z#���'A� r_piY�FJ]�<)�L�(n��\��oJ"m<t�����N�<ar��0g���S���oZ����FHI�<mo�$�r[:�2�� !�D��v<�Yʡ�ۂW��Y���քQ�!�ē:zL,���J7t�"$Sb	��`v!��>sǲ�Q�̋�|����&(�=\!�$I�z|
�hE��(��K^y6���ȓ1F�%����r��z&�J[���Xu~a�s#YSK(����,K(,�ȓ `
���U������EC�t }��v�������@�2�� �"��`�ȓP3�8�2�0j8$�%C�合���^��'���ɘҪX03\�-��7sd��*D�3v�%j�Y8��ȓT� P9S^)�xD��*�%N|�ȓY*:�	$�N�
`��Du�<��ȓ�,1[�I��l<r��K�#,:��|<�ag�V`&J0�C��(YS(���S�? �A�]�d��m1��H/w�6�p"Op�s��Xai|X�`-�W͆���"O��z惥oYnl���ݻd]�K�"O��z�o��9�~]��+jl(@ �"Ot؃q�G�P��A���
T��A�"OHt,�>0�RX��4JJ�-�B"O���0j� 3!@��1-ޕO��H5"O099��L2,`ۅʞM��Q��'��I�3��64H #�i�5/�d��'��tF�a0U��\�񠑀�'d
h�d��=�}��lA�R�չ�'�D� �G2`𑍇$U��)�'��Mi���6ͤ0�1'[�	�*
�'>�E6���7$�i�/�!�\��'�V�����M��x��Ő7r��b�'����s�M�Z�D�U��)w��9`�'&�e���Tp����ԨANe��'+ƍȅi�Mz�ȳ��<8�����'����Tm
s��!���+��e��'^�(�j�[�^�ɣ.�0����	�'>�-�t��=>������3Zv���'����(֡|;04�
Q*�b�2���j� ��	�K��l�FE�s�<�'DWA�qR�� 4% �A�Ff�<��
?W�dAc�9���e�<AǦ4;J Ȱ�JYlL�����`�<����-��M�b�-��ȳ�(�s�<A�.;��aKf	�5d��S��D�<!cϜ�zy���� �2ծ�'}�<�U�іI�pa�6��M��5���u�<�DI���1E@ \��&��[�<i�Ϣm{�M���ar���#	\�<� ��6HV��'K�TH��[�<AFlK�
G ={C�7�ZQ�7�
Z�<a���/j���K���%TLy��)�W�<�c@1<��1$5D�r)j�C�n�<�W��
���Q$��\B�i�<�'�J�0I��.M��Hr��h�<�#Ǚt��`!��'N��e�נ�K�<��G�z!P�bT��-)��P��"�J�<iFҚ'��{f�ʧC��c'ƈ{�<�oT�E:�q�5�
ENF�s�!�n�<���*0|0���)�*Z�hXs��h�<)�(�C�޵C�L�(X����d�<!�.��q{��n@E$����UZ�<��� ~؜[�L�s������P�<�$&O�ʩI#MS~Zz=�K�<ٰ���4�D�o ��	D�<I�����z��'x �r $���yR�A1ۦ �F��L�n@a�-���y�(Xv��xu�D��Q�I
�y�@�{� Q[d!;��B����y�� 4F\��A�D�J�a�t��
�y��
nn��%��@u��+!&���y����6E�4g�$BЉP�!ϣ�y���0��Ed�n
5��,��y2��+�i;N����1��;�y�����lK7IF���JcI2�y�䈇t��@'`�U2�(���7�y"FO�y�8��B� I2�zbB��y©֖��T P�'��x����1�y2���2��ma�="1����*(�y���5�u����HY�׍̍�y2�3YF�8� �p���y
� 2�����86<�-�����J
l�8f"O����OR2�ܕH�Z(8�ܜyB"O����֦ �����;B�4ɩs"O�(��d�R��BF�Hx�u07"O�$�`�!{�5�2��&��R"ODd2�9K�EŊ�J����"Ob�������Y֎m��"Ox0HA�OK������I�Z�@A"O�X���A�d��n���&D��"O��@w��9L��\QD�c8��'�||`��<� �Tɢ���1�'H�0�B�$�;4ʛ���"�'�*���F�	 8ݰ��vƼ�Q�'_�TG���3~�؃D����
�'�*h0��Y��z���&,>@I�	�'����`_{�x<���D�n�J �	�'���t��!�~hi�3�|��
�'n�,ڑ�v<�e� �&E��'��D1(��>\"�gI�g(����'�xxRc��kVhY���P�_6H<�
�'8�ء�f
�2��(yf)a
�'#ڥK& ń����l��D�q	�'�\�P7
eN�E�D!�z� �'��,KϘ:l�LKc71.@i�'gV͢`�DN�R8 '��,���	�'Ȓ!�EI�P�>�8�L�4�����'��R� �F�)피-xbPp�'%�9�H�;3��
��@�{䌜
�'<F�� X�gR4)*1���u����'��|�n�9K��8 M�{�h�j�'�p��4.��K��L@҂�a�BD�'��pR�ˆomP�qhݠ0<xi�'�(��(�ji�C �%,&���'���[�&�^� =� ���g��d��'�u��)�*r������Ya��8�'t�$S�K� �T��վ>���'�,��� -|��%�� :IO��'"���5�z TY#Q&��j�Ҥh�'�,@(�n$:��b 	^�8bD��'2V��1푴��T" �H�\T�P�'Py�(�*z�"�E#(��5�
�'��)�կ�*8,��Ѹ��=s�'%a��ˋ? �i��lՑm`A�
�'��!C��Ml�aYЫ��^0<�
�'4����-ؕeN��;�S�XF8�Y
�'��-�ѩO2��zgj��kv��
�'��h�
({��mivF�w��
�'VJxiմ�*i!V��}���	�'�*In-P] ��̞f�5��'�,���&nFq�ĕah�6"O$�sgU99VU��l���!"O�� ��  6�D�l� ��z "OLyA���=���0��`��+u"O�yrT�V~������A{Q"O�� ��]��ѩPgS�!�]_�<�@�PЀ��7�G'k�����!�@�/2:d9TaM�?�|���!�D�:J�T�aG*�w0Q�°!�!��G�z��̙ ��)8hp�Rr�־y�!��*w�J����5�`]Q䤜�/�!�dT3G^�M�S�VP�^���1`e!��v�N0r�L�o�zi �DR!�d�`~����Ōp�ʴic��� �!�d�+7D5��K�r�tU)F�7h�!�� ���f"�_���`�JF)-�iYC"O�T�k��=������&�h]��"Ovh�g.�����˚=��v"O�����[�'A�	� � �(��"O���T�&	b�u�Ǉ�;BŤ�S'"O8e���	C<�S-�>����"O�I���E�eYP��l�2`���	�"O�٨To�k�A�AD48��qQ"O�ljRk�^ݢ�Y�v�B!q�"O�e����6l�V�!�P�i(NXT"O�m+Ι�f8N���	�R�X1��"O�=J�iY��T��g��+~�v�ٷ"O��fҹ:yD!ӳ��>	���
"O*�`0A� [�m9nZ��!"O�)j��^�?��ԂU����f���"Oj�V���C���B�ꖻ_><C"O��a�"K"Uh<Ф�2)<("�"OА e�����3���~�er "O��[f��,,��R%��6�d��"O��1V�=T�$�_�uŴ��"O6p��6*���ЫJQN�Ӕ"O��N�-=n���5���c"!�s"O�4z�e�,ef0�@���+��!p"O��Y��P@�u��D֟@��@�t"OBt*֬�(j���rdM�R~�@h1"O�"A�:$I�B)͜���"O��n�u��2%�V1�ּ��"O^x�p+�G�\\��V�%ߐ�4"O1���I�d��,4[�|�N�s3"Ot�bL�-'<�s�֧U�^5��"OZ����ݛ�fF�:��Jv"O�Ls���|O���=m|M��"O�k�B�*�Ārw��aN�x�"O�|��!ߖ1��)��-D�x�vUb "O�q32ޑU���͂"h����""O(�C��gҌ:����?ID�W"O�R��eh8B Ç:X�0� "ONu��Fʖ	&$��o��� �""O�%�@�R�	������֐_��x[$"Of���ίS�$0e��H�\��"O�P'�Z���0'�Iǎ�P"OP�8��B�#�)2e�.���"Or�h �N*"�I8e^�A�H0��"ON�("��$JD*a³��=-�&S"O�if P�F�*�Č���L-�yr��`!X�!���8N<!��oL��yb��8}�j�Y��G�D�LXר�y�[!5v�)��A6���`��yR�G'\��IB���e W��y"��"��=�E�|�Nj�cM �y��Q�U^�� ��?t��ْ�ʃ��y"�J4(�Uq)ُn�Ԑ�TJ��y�&�!Kt�!E�h�"��,5�yrc�Jcb�g�[6�m�Ĉ��y�hތdq8��W�N 4��ȴ�8�y�ݙ')��#A�A)Jv�`���y�$:%�hěT�NF/�i�mH��y��B<)�ʤ��E�8\��C�Ɗ�Py��<hT��;w�Ĳ	G�@��-N`�<ac��mk2ES��̨#l���.\�<��'#�0� rA�#sV>U���\\�<IB�Z�1��e��K�r�GVA�<)0a�+~#�Y�兜[c$\� �{�<i�E�/�>DP��I ]㊼��dJp�<� @}�"kV�4��͘g���p�pq�"O*@3F��yz��Z��;m�eɰ"Oy�����[�zeء!x�Q��"O�`�5#��G�W85��%F�ϱ�y�G�{�@��w"�(kD̪��.�y�Y8��S�n�1Wt� �yR��Df|1E��)D���7�=�y��-@]� I�DN�&'�S�����yR QBnB�T� �u���fG)�y�+��bwp�XqM�]�&8ˠ�!�y���2�n �Eą@���$���y�õ��۷�'��y{ԍ�y�N 1�F]�UC\�W$�c�O�yφ4.����F+.zt�SF�ybǉ�+Uty�0�B� �lRc�Ⱥ�y��G�t�r@�/^
#(B��2�y�CK5\�$�4�~�X1�'B��yr��-������3w�N�C�&���y� I&HN�yQmL�g4�,�6LB��yR�Q�.BPL����� �{����y2˄�I!�y��/D�u> Qf���y���+:x���.��Z��0�)�2�y2�	&*%�����c�Rd���N4�yr�8N7��qTK�b�L�`��ܠ�y��Y�O��#	���U���7�y��]�Tc�Q�r&мD��!���y�d��1Ʉa���a����M�y2��N�\T����-~4 `�&�S7�yr#O�q�b��)ZẍuÖkR��y���;�R��دY�TA��3�y���0c^� ��9P��AZ��Û�y�"صdon`��G���{��$�y�D@k|��B?��0�@�-�y҄�e0`�[E�
t<��g/���y�%͑q�j�!#e[�V�	2G�^�y�m�V�Ztz���H��T��G���y� L	;�T+�
X$EK��q�K�#�yC�)�<�RRI؝o�li#,�y���LE^�D �*bF�!�ՃR��y��0Q��1����Y���R@��yR�ǜJ�y�i)��2���'�y�aW	P��頧��Di;�O��ybL̨7]D��'��c�A��y�!N� ƘѤl�9~ap��!H��y£�rv�mH�L��_��\!!)��yҧ�
9�Pe�S(��h��=�y���8<ݐH�!�ш0������y"��T.-�Q"0.q���v�S��y��5�H��1�T�<��c�O�<1 b�"\*��W��z!��8&HK�<! �V0u�vTj��%��їK^�<�cb�X�DDpR-Z�k�и��Ir�<!s!6,�\$�CGE0����#$�k�<Ih"B�^\J!���f���7�yB 'oo�P�@��U��.�y��BBqܡ���֨.�٩ӡ��yB�$�D܈ħS"��s�P�y"/D�i�\���lR9+��˂i��y�[�h�!2�j#�HY�ś��y���G��jӪ����IB���y"C�7:'�thd�&N4�x��Ֆ�y�`�e���a� ��IBWCZ��y�OKW?>�(тA�:�i�-�y�FI�(GTĸa��{7F�QW돍�y
� �)Ę�^0f�a�h��.tZ��B"O^Ȋ���KB��rc�ȋM�c"Orq L�!�b�EG�fH�"O.�s��):��� �ǭu��Ȁ�"O�ۄ�]N�v��WgҘG����"O�uA�H�7v+f�[`��;Jv����"O��z�I%Q�N�9󌂇7N|Y�"O.��S��-r \)@#kWPA�؂�"O�	qpѡ4��	�R0+
��1"O��#E�U ���F�J�z��"OF� ��?��%��X�4:�X�"O�9	2��7T��A����; ��U"ORy)A� %�4ِm�>�h�"O��"��F�\�z�Í�>r���"O�(�a���\�Mm>�"O��B #��V���$P�H�"���"O�Tbtf/4���QK������"O���ƈ�w�1���I�^�2�zF"OT�����'5p�i[1~���2�"Of��F��U8Wk�;�`���"O��)�ķ}Tӓ��<w�Q{�"O�C����6�&����"dH�Cb"Ozuh�B���i��I��K��)��*O��&  3.�D�cB�!`ڡZ�'�zH#���Uβ�02M���2�ۉ�4�	XV(XwO)�@9c�┉���ȓ\	jL�W&�q��M��_A@U�ȓ.2��* ,�,ie~E �A�n���e/8kJ9_�X���&��Q��d"?����"W*e��$O54a�(W��0fv!�$��V�<�6B�
>ʴ�5�Z56?��d1�S�d�38��(�ǚ�/| ;�
X��yB-�
ȴ��Т�COdY�@'���y"�V<���9s�6 � %���yr�A�m10yJ��ճW�-R����?Q�'�r��㇛�+�P�1e)�Mr��	�'�hd��ն���!S).�b�	��hO2�!QdZ�f��1�5,�.[V�Y[3"O�A*���MI�JZ���`�i�ў"~n�7��Hq��!�F�2U%[���B�Ifƴ�!�RwDݘ�(M�6�j���������
�� �f�,h�D����3	@� �O��"D owƐۓJ��;����g���vN��HD�.�bu�ӮٳD��{����I�+q��J����!A ��!\ +�l�s��)�矘Se���>��$��b_0E ���d5�	y���)�O��"t��-ڄ4�՚w�P�`��O����6W<�: H��[�`:��R(Gga}��>I6�n��Y�F6U!*�[�#�\�<%��r�"y�U2E� �
A�KP��hO�O
e#���	l��գ��Q����'�����Q��y�P��K�q8�'�L��懬-�~D`�NE�B ����/}r^������Ц��5=b�Dܭ9�v�B����#Tu�&Q�Ne�p$>O�"=�w"�:�2P����&k��\Q��N�<9!�Z4DiNA�X+2|<y������;��i�a���>�ص�I�W�����8�A��Q'y����n�#	���ȓ5-�[��V(l�e@Ԍ��1����ȓP6ˠ�@*T:��s	g	�rm#D���2���v#�ps��"b	���+D��bP��~�d��� �l�.�;�,>D�܀�*�78���Ch��$;,����<�<�S�g�? ��٥� ��)x�G��X�TI�"O�H��V4�zq@� ك�(IH�"OT� #��"<BJ	xS/K}�tK"O�|���� su^q�5RaVHSu"Oz��=Q���UB�q��K�"O\��4.M�
����gԗ��D"O���&H�"u"�0���F1:������_X��+#�69�|u��%�<���xu�3D���d���h�`��c2��:@&D�h�Kկ
�� 0��^yt�2��$�$2�	`̧�?�K�Nd:��n@�5-t��g��:i�B�I!d�H]0�c���>��6�\�(+B�	P����p"C�OA����U��C�ɴ[!t�$��3<H΅Y1�� P���?�HO�>apGnɗS�\�� N�76���,0D��r0�M�}i��7�-lu֐ �A.D�p���E��<�� E[c�|˵�(<O�"<A���
��(�vˊ���Ș��t�<Q�&MⰩ�gY.D�Z��gHs�<yG��e|����)m�n�#KKm��<�<�t�6D@��S�@]�N���E�Tl�<���N�oӚ�+q�T";;�x�#
T�<����N�d\��]&dMhY���R�<��K�oYP���I�\��i0D�L�<u�ЧDb`�P�F#K���ȓG`�Y��M�h�ðj�(�^<�ȓ@��xȥ L�f���d�j�ɇȓ4�x%JG͚�eW�Ѩ�hQ:���'���D�����7I����##�	W%��Q��&es!���P��p�Rn��W9����']!�d)e�4("D�=m��e���L���D�$+U?#F�q@�нt5�`�����y�oܛ�> ��a�!�ݙ�����y�kg�<:3�J����T/N+�yRĜ>ĴL!	٠ZX�5�A��PyBb�c_`E��H[�D�����D�<���9<�0$aC�>OT��.������z�"�Yр,a/v��p������:f~	����7�A��%D�Mf����[�"	�`��x�d-�$�A;a�X��ȓ[�phU虓N�j���A�� �Zh�ȓ8>����U7CQ�)ґ	�$Zp(����
'ў�}
AeΒs�$ل��K��c�D�g؟$KW�'�@��D�A�����:'R.�ˏ��6O�)��ςyɾ��N�M=:(�q�	u�Oi�b��#��%8r��j=Z1�'T@���
�"T�@A�3XCP�*���If����H�4��ʑ�� DB�	1\=��bB�J�m"d0�j 0".B�	?N�H	�p�ej&�x��C���C�ɳo�P��bnތ	�"��FA?Q��C�I�gצ\�'$5{D�Ёe�K�m����4�ɦR9Zq�\\��[��;�6�,�S��M���
�]K�Ч�
��P�KR�<���z����D�/N�D�Bqˁ�E����(�ɦ*F�BgD��p*�#T�[ ��C�5N���+�/��d!�&jא}�B�	�x���.�ԐG��C}�B�Ʌ���'�Ԁp� �Wl��.L�C�I9�����DmTC�'��Iq"OH!	�8"r�X��1р�"O0�a�N�)��eV*V&J����O���W�rD��"@ӑm�`�rFe�t�IQ����Հ�8�QjT�Di�x�8S@.���)� ���D��T���hc@�;��f�O�b�PF{�������0z�R� �ѽm,`zg"O��(��(8Z��Ε�h).|Qg"O��r��>B�| ���(B�;T�$G{�剂"/aZg�ߪ��H$�
��B�	�[��R"�u��P��I�m�2��^؟�YuoT u�n�bK� �F ��� ړ����Dh�h#�Zs�"uy���As<)��<1��哝	6Fi(��T��Ih�O�
lB�I6A��Qc��
!���C+mƞB�	"{}vI�cC�@"�(��ܷ3�h��hOQ>��pdԥ{��)D�_�^r0��#D�dz��U=�@yS+���ͫgj�E8��Ez���0�")"�/�$��Q	��
�y2@�:_n����G��c���M��'�̠3ת�n���P�D�QM�H	�����Gv!��J=�I�
րvB!���,i읺�m�8�șa�ɀ�E:!�D�?�*p� m� �h��c��8*!��:q�L	[$���.���&�Z�6!�DV�o5TaR�.C�{��<"�CM!���4�T)3�E��H��)�v�Ҿ����7�S�O����㟩��DDG$*'،#�"O�A�`n���~p�'��*vig"O��&�;MV橸��G�%=l�ۖ"O
���X3���`�OIW�N,c�"O(��^,`~��c�DϮhhz�Z6"O��؜��� g�ʇn_�}B""Ofh�@�»},DB1]WJe��"Oj��g$^H�ڣ�פ9:Ir1"O������Z��Pcq@�%M�΁K�"O| ZQC32���(�R5�1�s"O0p�EEAg��˗�`���x""O��:�DS
n��:@aW�P��sB"O6Se�h���oR�o�v��R"O�Hȓ#��f$��F�I�S��@ڔ"O�PB0#=R�Pq�CޖF;$Uz "Ob����[�V�Li��6A2�qs�"O�K�������v&�(yv"O�� �XGʕ���T����"O���w�ƅ�����5���"O��)W�D��5��'
d�ȓW=L��b�I�L����[B,�,��r8�	��.�B�`�;��ȓO
��t��d�5y��N�U��=��qo.���@�P�8�̅�eu�ąȓ&} ���N� ���ʀ�D�ȓ¶�	�ޗL3xA��KGl��a���ヅ��A�tꙃ@2D�ȓBt���s�Z�\��p;#*�-Ƞ��ȓl�:E�F�[P�mk󯐪jn�ȓ[�h�IB�+?UXY�v�')s�ć�/��U�e�	��-�!2�й�ȓK�tQ;�	&;ʅRE��$8^��ȓ:D�a����J���p�C�PP�h�ȓ��ɓtE���� �$�x��4�5H�`�nE�IZ��O��!��2+tUb�f�Sn��ȓjV���	ə3h�dPf刿ފ���DTT	�����<v��4, �ȓB�*`�a&��
�L�t!�d͔E�<����	cyS�Låi|��`�g�D����5�ўUF��i���,�Q�ȓY�����Un��I�V�&Q�Lȅȓ(R�HJr�[;6���rV�����S�? �t2�I�\Q�G�E�0���"O��Xb�	8\�l�âU�Q�dj�"O�rG)_�Uc�Œ#!�K0�ՑB"O�uZ���?Z��@�k�.$��"O�}8�O�J�ʬ`�
O(j:r�`!"O^A)��]��D�f�҆`-Ԉ�"O*�ѳ+��3/��1�]"1zy�e"O�qhG��&z>�pD���␉#"Oܰ1c��m=�`�E�!<�i�"OB ���¬���E� ,w
�;�"O��:�ßMa�!	1�1R|Te�"OD(#�[�^�(4�d��;2�"%f"O�$T4z���JsB̕�ex�"Oܜ���,NR�p���tȜ�QR"O��C�ʂ_*H�灋8U^	�S"O��(Q��,^<p��1x���"O���u�ۭ�8@�w!�"O��D�4"Oh��̎�k!����Rh㐔[S"Oj-�Ud��xQ�φ�R�b���"O�PZR)�;'JhIs�HAS���z�"ORpqb�]'��Py&홱d>�R�"O��s)G)~05A�mK*te��A�"O*}bA�Ϻn���2`%Ä^Z`Z�"O�6�J�9.P5q�/^�4rh�d"O�tSB�771LM@E�-%>�V"Oh����9g�B�AG�^�tI�m�"O�0avE��]� ���r	I� "O<#C�ܯh����%�%6����"O�Iӡaù#����� #&~t�"O��Hĉ��H��F�H�ur�"O:	9�E'0V�2�cCt���"O������-D���A3(���"O�)��# H���)��q�����"O�P���*B�,�+rmԯ*|l�{�"O�x�+�;	��\��È�[���s"O�!���=f��u�B\n_���"O$@�����AR�@)��R"O��d��7|^�s��*h�H�"O")�u�+J^8Z�N��y���x4"O@�D석#�ZB�="Kdh�"O.ѡcA�p3P0SGd�3o�P�"O�� �"�1H�A�3%���S "O��V���flze���}_X��"O�02�'"t��E!� ʹ�ۢ"ONa�U)	�"g�؞}rҭ��"O(P�#.[��M`���<����"Ox�0�b�~��""V�:˸�q�"Ob�3��Gs��TC�l֑%���3"On����M�Q���G#r���"O��xw�;kЕ�!\�|�E��"O���t�p/��CG�'[:��"OF|���G2�8:�c�4ml̸��"O6e X�x�Q�VA�%[j�I�"O����K+B�\ٓv�H�(8R�I�"O����V�XMvl�"�٥R��*�"O4���o[5f��k��B�:P2�"�"O�\Q��W3+P��؅��0yQ�͈#"O�Š��^)Q��u��&Ј(vD`x�"O�\�7�D?ha#V�Z2A0�p�"O��SfI�#����̖D�Xdp�"O�YY��)Q���Bg\�NR�ar"O����I]3���ש��Go>�"O`}�#�>E"�X&�P0|&Ta)q"O�(9����p>�
�'9s6�	�"O� $�*ELC+\U�G�0�"P�v"O�����G3\�n�0�Ӊ%_�Q�k���|<˵���O���u�]y�e�v#�8d�19"O��c@�ĀlQ5!^�"N"���'uH��P�T����?=����ڎ\a*l%(�)y&�{�6S����7"?<�X��u�\�k�J �@R��k#D�,���Ѽ���޹eu�QPS�>;� �6����̘��Ӯ8�P*7�+|��=c�̀Zt�C�I/"����C�HQ�%� ���غ�B��UX6�$e���ؖ�<��b�ZꦘhUGU9]�h0i%M�O�<�ց(9��`aDN2s�Z9�c,ҽl���Sj�#J�w-��<��Mc	��:�����L$Ӧ`�x��хւo,�Y�i��fj�t��e�2!�BOƈdE2a���wh<	����q� �s�dD�Ci�r�nX� d*65�U����O�P���舩��td����'� &��@����j�#v����$a�g]�QZT_�ϝ�����6J.�	: j֧m6�q�f�w�.C�ɻS&#4'T�r�\5C��ßJ3��`�B2GxXaB'�T�G�>�特da��ڗ�ƂA
r|iÃk���D�?����0P�=#C�M��""ƒ�K K��Af�	�O��P�)֖a|���Z0ްq0e��0۾Qx� ڋA�ly9F !�S�h���1fE1q�]2���h�B䉕,#���� �Q�*Ԝ��@�b�uS�e�AA��T4�<q�B��{�
Ī1�'gs�U��(I\�<qUcZ� ��]��c�!r{�1���X#W4�))�)�I8��'\c�����a�dT	cFѺ6��D
E!2lO� B���J�"T��#Äf�A" '��kj8*���iG��)�A[C$��P�NT{�eϑK���?1R� �3Q4L���(�'��5���B�v�8�"f �r����ȓ�n�[��(�p�9v�\j=����V�D���=E�����[�B�&m��S�%�:D�<�T͌�5N�C�ĭ��,�d�;D��A`�=���z����Y� 6D�tP1��A��=Kƃ�]��r�c;D���-Q�v���sELݟ8� i�a;D�awo%m��iUD�I�QX�b,D�����0���S�+K,tD��s�,D�ܨ�lz����-�<�|����1D�`���ߩ{Vrt��E�,]sD�-D��q�Y�Y���Lϱ*$ �%*D����T�Jq�R�*/,���)D�����$��)�I����c�3D���!��xQi��Z��ʅz��.D���VN��N��� �O׼nv����,D�@��ǆ3(}t��P�\&\���%9D���ǚ4�U��g�-}�X:F/9D���E@7"L4hC!£aˤ���*D��0����P�i��J\Z��)D�S�D�rԘ���z�vip1�-D�$���
).u<����,ِ8T�'D��{�k�9߀ٲM�)�| cf�$D���4�\,{�u�pk׃�@\
"�#D�K�j���m��Ò�jU�>D�`�W	\�Rl�PPl��%K�)�E�+D���"농:)N� WlO�ԹA�N(D�,Y���[f��f���p\0g�(D��p�"بO�~�#�K J�t�G�8D��87O�0"b��X�`4�&��	7D���&��TrD��Uև�����&D�$kE��|����a��	{��ւ&D��D�ǒi�@��щ���}PM$D��qkԝ#��]K��]0�}9�m9D�tE�}�q�G�֠n>pIɐ�9D�\��R��:L�艣��:D�� �N@���@�k�8
��"�"O� Z�Ŕr�왕C<��-y$"O�$�)�X��z �UA���K�"O~-+q���:u37�@*F�ի�"Of�jwmwb��ㄐ���` "O ��ET�z(���A�a(Q�|���ɓ]`Sq��=�$�A� �!�$[����JSԓ<������^	Ӱ�=E��'괰�2�9�4I3�Y 6x�z�'Ls��	B�2|J7eٶ�'��j
�N�����߱h����P���0>iL>����%E�d	��Q64r>x@B�D�<�s�8uz[t��$�0׌TC�<�elY2	T,T8r)�+4�0�/ E�<�`IߖO�b�apH�;[�DR4�GN�<�C��pX��Μ$��͘�,�I�<��I�7?�4�'#����t*�	I�<�cCRi�@�`&�>A�r8Z`�y�<AA'��HZYV`V56�y���w�<q�jӃ|r^Ly�IP��|��Aes�<���J;G�=���:�}���s�<	�H�21S�W.+���2�[j�	�]T"#<�~�S ��x?�(`���7�'B$C�I?�v0i�N��E$�X�&ŎEf�㟠ȑ�'Z���&B%`>q���I&	�5;�'ZZI"��7	����O2p�Y�O�����^��-��H#_R�� �'
�O��a��)tt@�b�5 	�"Obd�%	�%Dڽ�'�P�
c�K�y�?~�^	�@ǔ�^���pG0�y©C(_�^����M=Nu���/�y��ҏs>ȭT*Q=����GD�&�ybbR0jdvL�3�	aW�@����y�Y�+j�4�K�g�<9�G
�y�MY%��٥eYS�ڴP�%'�y��A�J��i�$(ڐN�ha�bF���y�d){ʬ�Г�+w�ֱQ��
�y�B��}��d�;x�6tqD"��y��0M���R�����l��ӯȿ�y2���T�n�8#�	
���Z���y�Iߒ�
���J��x����R�F �y��B<A�<�6eA�{�Hh�����y��-U��"�	�|��)�(��Py(�9y�P(�%ț>P&f�Bl�X�<��
5/sZ@3񄔖5�H��C�<1�F�L&�00������tM�{�<)�Oפ`�rѻ�O�+�H��J�<1�%��t��#h�����{�<y���ઑq���z�� �%�[�<I`A
T�d��C č!‹���M�<1ꆁx��� �����$���!I�<�� �\���j��*O���I�J�<	¥���q%	֜;VPɊs�@�<1�+��`�oF�Xvv�W�k�<�'�^�}4�p��0�I�0�]�<)�k^�����@c�k6T�)&��_�<�CjW����R"
���#�S�<��ꅹxB���Á�&�MP �r�<� �Y�nK@��g�H������Z�<Y���3z�a���ђ�̡KB�W�<�PI �H�ɥ�Vo��5Sp�J�<��O�|�9ʓKF�bv1;�IA�<�d��@��P��8��,�RMX}�<ɲ��w�<�K��̕'��t�*Cu�<� �D�(�hH U�G��RP��"O�1�6��.�j�{s)܆b<F�"�"O�i��\�I�"P8u�Õ4h��"O^��vf�9MU�5Q�Nb�LX"O���c�6*��ˡ!��6p ��"O4͘�l��v�P�Z2V�"O���צ�-]=�bKҳ)�aI6"O�J��d �	�B��8)pp�Q�"OX�5�C!�Q��+��q"O|Hs�K��*0G#^�֜�"Of� �j�QKP�2����"�  C"O�Q��铯|f�F��.Q�\�7"O
�%�x��jC��2gT*���"O$��L�@!�X &�ɊF10�"Ov��K��c�xjfeQ�pL��`"O�mZ�;�Zbcߛ]R��"O����S]�Pq2`ւm��H�"O��+EI�4|zi��E��.X�W"O~��D!_*� ��d�<���	�"O���I�d������]�lB��"O�����8f��r ��$���"O���5*́c`����Z�cs���0"O��"F�u��Г�+#�D� �"O ��e�	0��Q3Nek2��"Ov`Oۿ����EkZ�vT����"O�����0[�`W�Ѐ	[���"O*=�Rg��<��5i�X%�e��"O�0Z�fS�1�d��шP�:�6yF"O�PHw�8�j�e��$�����"O0����;��1�v�I'^�v�$"O�H��N�+01L(5h�pTB���"OXt0�.я2���BGN+&@�$0"O.mb �I�w��x������"Ol����I�RdI�T��D��8s�"O�Ԑb	�]*Ȋs���9��!�"O��S��.:�T��ȵD�$az"OL,+�c�����Á��@����"O\���E�j�� j�4��]�"O�uqN5<+j��T<{rx��"O�e�V�r|Bf�ѬS���%"O�p�a��h���ƨƲ�Ε w"O�IS&cV(M�Zi���G�8h���"Oґ����IBL��ϐ�vn�� a"O��;��ja�/�'\��)�6��)�!�DX�o�����
ɂ`٨�����,z!���p��������`]�.ԶYs!�D@�n�:ؚ��\�[�txH'��[!�İ bh(�A��|<�1P���:H�!�DG�	|�Y#pJ�/*�HU�H��!��%J�>L�V�1�d�O 5�!�8{툑�ե��W�����}�!��;E���3``�,qf�i���k�!�dr��a��f�7a(���KF�!����q���O�k�t� U
��!�D� *�Y2��Cx�	R jM,<�!�WNJ�����֜\6�\����(!�$�|��UXU��,Ҡ���1!�E$�V��1Q��L3!�	F>`$r�fQ�[㞙!�e�3�!��*)�h9�� c�f`ʗ� ��!�D��Z� �h7l�5�,��eϮ�!�҃F�ڄ�%��(��C׈ �S!��ʋ �pI��3|�6Pˆ钅^/!��v����)�z��§��m!�� "9�p&S�FE�����ȯgix�2w"O�ɱ��;Xj���T�]N "�"O@��"��l����	�`"O*�p�拱H�F���L}����"OpL@ ]�[o�%!��چXP��"O�ERf�U+&��uaJ�,��L��"O°Q%�G�jmҨ��I��t���"O��P穖�V�,p�b�N�p�"ODu���^�Ҕ�W<���%"Ot�0A���8�.�;1ٴ}��"O�P���8��킳���'"O��Еh�k|� �.7�F���"O$@ �ED�U���j7�<S"O�� R�;��Z�j��qL��HT"Od��fG�;Ls `�i̇%@�a�"O~��ŉA=���Q�hT�ސ�6"O ��O����X6D�`�"O���E�lߖ�$$ !$%D��"O�uxCk=L{�����'`�I`w"OD��G�.9��-���ԭ(��G"O"�E�<�HY����0��<u"O�T �'5�|`Di��H�"OhTSBL$d�eh]�A�v �"O$� b�oǂ���lO�d��� "O 	�&�4M�@�Y@�D!Wp�L�r"O�$��Fݜt�"!�R	ۭ*��]"O,ջR����Yk�ȭ8��4�@"O�y�@�8}��U�xrb���"Op|d�P�w�hH裬Z�qa5b'"O����ɬ���[�Y�qX�"O$5Y�ϔ�����
F%}�q"O��"/7��Qgʁa�H	:�"O<[F��RH�u��IB���W�yҡԛ�f@��O��:�
$:���yr�H)g�B�2��ߋ>�I�teU�y�G�V
���͉�,Fh��`I�y���84st4��œ)��e�$ᙈ�yB�1E�t! �F�)�0:�h���yB�A9�օH3(-/�9��H��yb�p%>aUH�"&��i�AK���y�@�C|��˵�+^��R!����y��Eh�ȉx�e���Z�L�/�y�Y�m=Nps�
���c%��yg� ��H(B%���f �y�
��� �ɸr0�dr�hC�y��ǻK���3���hx^�W(�=�y*�+h�hRw)��a
@�V ٱ�y2�ցGf6����U�5FnP��� �yR�F�D��\ �cϦ6�N�c�i[��y2̅�vq�!�ц0<��1�J�yB�]=<@E����;�4�؀���yB#��4w"��%��x���	�-�yB�Ò.�<����n؊��0�Ͼ�y�"U��*�j��a�T�者Y��y"�\�l(�Hb%��c
��'����y��Z.0¦�p0�
5\X�HJ�$K��y�o@3T��zwmY	P� I*UM��yR��.1��ǅ�K�uP�n�	�y�� kF������"A�M۰����yR�ٟr�D�W�=9�bp� �'�r�Q��שLU\��ȇ}����
�'�
�hgm!~�>HZ���m����	�'�ށ�D��Y�8����H�\�|�I�'�Ь��!�/	���+$���h��� �a���?*r	!T�өDK��V"O�%�&�P�����M�6#M���4"O�4��a$���8��9t�9�d"O6����,b	+���+O��U�c"Or����QbHZA���58��@B"OD��I�-b��tCHQ$đ{�"O|e����iv������
���r�"O
@�3�B=] pQZ��ތԜ�!1"O.�C�MP!gr��#�D� �t�"Od��ۈ"���y�xƒ��B"Oh0��ي#�`�BU�.�^���"O�tYCm	�$�hi����0H,�"O%p�[�i�j=�T�� a8�bw"O�� ���<�& �U��
��)�'!����2$0�͈�7?��a�'�|	��MҪ'�(iP�e	pwB�k�'�H5#����l�jY�&�LjE��b�'��y�oɛ7��z�NڮY4q��'��+TK�����������'��$���֘/ލbS��/����'Z���E �7Zr�}q#�[�$�r��
�'�PD8������@I
�'-jH���[�4͔�2�T��j�Q�'��9����?[dD�f��s�d�)�'�����ꚦs�n9��u�,�z�'b�(�奊Ȇec2D-3�$���'V�=d,ʫnr-A�P-0`���'��M�Q�����s���yʬX#	�'�M�4��0Z{,���mNi�'_�P�WBՓXe股ӵTO D�
�'Ʈ�;��U#M�v��$��7W����'��ѩe�' ��`&�,@��#�'v)Rf �=!]��pEӤ$�H3�'ΘBT�ɩ$>ɠd�߀$0�Y�	�'�(�X���>��U��`9�&��'XRE���N,(#Jl�u�_4p��,8�'������ �d�Eg�{:V���'¬]��ס�K%�[�i�@<��'�b�O�l�>%k�jV(`u|�	�'Ѫ���X!;��P�OU,s*��x	�'����N3!#�I��Fh ̀�'�Ģ7%��)NѨ`�ɵm�J!��'�\��Z$n�e�֊ݝf����'?�L��'���@VY"!H�'X-2 h��z�J���o����A�'Sp [���9K��x2�X�'��DA��:#T��$.�	�ͳ�'���K��نs�DP�hސ��#�'O*x�u�K1,m��Cژv(Y�'�0��
ZV�F �㌵]t���'9 mH��3I���+r�j\uB�'&Y��K9�`$��IF�\���'��)סV(V�. 8��h2(��'^ԉjf�h�y[�H��X3�'�Ni�e�f�Pp�H�<͓
�'��iw���eT ��gꒄ6f<!
�'0H���<[R�*�"�<&����	�'wx@��B��;���hŬL )Y�t
�'2�9E�ݨ^�N
�˝�+� �Z
�'h� �d�;X>@���ۗ"5��!	�'^�Q"K;6¦��#�A1w9քP�'d�m��d��H6Y�)�,i�L��
�'浩�Đ�4<p�0��e����	�'H�r���4�L"�o�8PA�4���� �ᚦiC�X�X}�O�H��YЅ"O��
�F
��Di�đ.��b�"Ob|0X �SDfY�%��vh�V�<IC�́9�dX'-د�j�1���P�<)Cf³��9S"ب�P��_Y̓�h��ޚ5j:+Q�_�4+���<�E�ܱW��!V�]�!������T}B�'�Ѳ���"�H� Ǽ@� �����hOQ?���B�+8�.��� ��Ѐ�>ړ�0|���B�:.��ª>F1
����z���hO�'���c��D�5�䴻�"�Y&x'��G{��DE]�
���iU��
s�z :�����<1��0|ڰOK!|�9Sm�N�Бq�L�&�ԅ�	�Px�"S-ޚ[ *б�K�O���Dl�$
��xN���Fȁ=_�~� ah>��O����9YM����L� �t�HOcΓO�=�}2`"]�uI�GY�N6�����Oy��)�':@h�+@$,H�`x�pŅVN �ȓ;Z}82��)'�Q�,ՋDàM����<1��H2a��H;SlJ2~�dy��m��hO�'n��M�������⎕���/��<�S�'u!�a��f wA�sO#�`U�'�ў�|��QF�1ۢмc�� �B�Q�<Q��Y�l!��鈮n���tPcy��'��	c>�"�@N/]q<�2��$0�C��<�(O�=���9���Ӣ@�p�5C=�ʴ@Н|"�)�'Q�E���Z/)b4�V^�U����hOQ>����M��� �mCM��P��Oޢ=E���ۦ")�	P2�2���'E �hO���D�6 p⵬A�>-US�i�Q5Q�\D|2�ƶ*l����4Q�����
}��p�'(D�l����#r��pyW��7&!X��&D���j�L��`�MZ��<ȵ%D��Z� I��rO�{��8�O$D���r��QҜ�B�AD�.Xn�s�&D���	�+?mvE�`�D~�*�;C�#D��1ac@�T�e���3��x(#D�+���V�8���,7?���'�6D�ı�D݇& ��r�PL�`� ��>D���R q��M�p�Q$.� ���8D�H8 b2w��,BBS�!��%��8D������!���DcѮ���32&2D��A�%�-qv�۔AO-��Bq�1D�@آ�ݮ�`�(�
�yc7�0D���!��l^�U�i3����,D����� %	PP��F2�5�1&-D���s�S�^�i*����w��z��,D���FV���B� 80�ܠ�-D�P[�`��|]�=��hY�	[p!�*D��i�.l��6����(D����),@k��&F�->nhT��f&D�l�#/�5�+!���1�TtR#D�$!�^훤�ښv��# D�TA ��R��s�m�	�tQ���>D����`V
]$���#��1C�<D���A@}:�{VBY6�`aZb7D� ����^��qH��$8���A4D����D��4����s�<�$$?D�,s ��9�����Ɂk�r�x��1D�h�0�^8D���!%��h�i3�+D�<���L�l(�� EG��+d$D��#E� ,>���#w��a�4/.D��Q��٧
�F�if�!�'m*D�l�w���Yh�UI�Jp�s*$D��J�!�	7�\1b�H��<lY@%D�� �y�g�Y�xx(��ԐR�"O^����ϕ4\v��G�=[�0@"O��r��9�>iYr��8�x��"O�}y�����@ש���� V"OP�nC�L_Tq�	[��hXٳ"O�Q��H�2.��(ۇ0���"Ob��,^�{d�	�3*�E����"O�up@'X�l��Q�
�?ItM`�"O6����"+����ᩎ�W�İ�"Ojh�$*5Ȫx;�'�&�I�f"O ��*N�����e������"O�� /��zԞS����;&|�"Oz�� H�v���g��,x�V�r�"O��ʰ!Q�j�
��S�
ٸ�"O�x�A�H�0e�����>R�)C"O@ER7�Ӵ��Oĕ��"O��A!��.6��t��%}Jl���"O�a��Iׂq��ɀ.ɘ/́3�"O𨻇��&2���M_+%�A��"O>]�0Ć�9�����'T�r�"O�M�  �^a�MC��Y��$�"O���n��v-�RJ�
"�L�"O`a@���=8����6��h�}��"O,A��ŗ �"Y *зa��c"O��h%IY�C�pP�*G/dh��`"O�L����k.|A�ת�Y�U�"O��4+οK�`8g�F,�����"O�x�ע�>	N���=1k����"O�E�D	�Wj�h�̈SWRٙ"O�\˔��n�����+����s6"O���"�6a�r�h�=���ѣ*O�(` �W�2��DٓHJ=H���'u���'bW�~x�C��2	����'K�(����1b�Dj��	;^�%��'�����̄�����(,�Dec�'��l5�A�X�$�Q@�&����'�&��@A"42��(%�U0���z�'�l��tLC2$�$;8�t8	�'�aY��>1" a]h.���'�U17��63`�$��d�<���;�'��Y{�P�$��t�H�}> ��'����Iҏ(�"#CI,,*<@�'A4�Pb ��/���z�h�'��t��!~8��c�C��L9s�'6Z�����SǺ�a��:r�4�R�'
V$�@MH�.H�A� ɚ5k>���
�'�Ή��̯>������VX�0P2
�'���G,S�ݸ��!�Z���'����
ér��Q��eL(!Q�X��'�~١�],z�9��ƆD����'����%��|j*;�+���'m�E�"l�4zŮ�{hZ�]�i�
�'E@��w��Y}l�����}����'�4�1�×}��q���sۘѻ�'DB��"Ƞ$�zD��:{�*J	�'�	������.�F��L��'Z��P��Q��r��۪9Ȕ�z�'g�m8�T5Z���B��j(��'G�e�C��gV|��B�%?T��'�P|R� +7��iqfC�����Py�d,ͨ|�fBP�&�8��D�e�<����Y��8u��s1��g��f�<�ǡ�1�&ĚҩxWZ`�@�We�<����2|ّe
�8HC&)ef�\�<� ��J�gԉQ��j�cOi����"O�u�t��4QD���"��z�B(�A"O̸zvf������RE�K�����"O����˹+x�
2���T�"Ov�m@Se*�j3 	�hת8�P"O�q	�MB�u2R����ܿ6�T��"Oi��)E�
έ�V��7j��e#&*O*:� 
�w����G:�� �'ºЩRJЩB�\i����?/���*�'7�)�̚(�nlQ���.ZZl:�'�TEJ*oUڱ��aƧq#訳�'�Z��h���Ă�6��;�'�,E�g�(�传r��).��a��'� S>�U�EH�,B^��'�ҍ$��!=��
ɽQ�(��'��IIs+_��fYP%O�N���
�'тW��YkT�p1"��iY`��WJ)D����Ėmk��Cb��*
X���:D�(0�܆6-"T�c�ɜMU�H���7D������1)�B�`� �\����4D��`p��8˴y��*Da6�c�3D�Y�l�=����P���a�$#<D��z���f��lJ^)Rx)B`:D��x 	��_�`h���c���ą6D��97���fƸ�q)��cꨕ�&� D��BG׏ĺ���#kn@��>D����Odn*�BV���XЂF)D��+�ʇ�;>� ��
�83�C�B;D�,����$����G�{�.-���7D���f��[�x��En�9��2�5D��x��Ĉ"���!E$�

����L!D��B���R�(���,ŲH{,����,D�p�׍�O�2ii4�B�)�L]��?D��!B猑�\xjW垤C�>��b�>D����݅3�!qV"]��<���<D�y �νp��=8��M���5�:D�la�U�U
lIh j	� �F���8D�*��˰BѮ8wŜFR,a)d7D����k�$ ������.�愈�/D�|�RE�&�2([���
$�CD/D�<��薁!2B�h��ˣS�4�tC,D��"D��<�9t)ɢ2!����?D��D��n��e�e@Ɇ�.m��(D��
��0	�1�W!ǙN��\�T $D���#MC�?-(x�b�R�'q8E�5	$D�X(�f�	�����Q�6&}b�&-D���fd��G�AA%��9�!K�+%D��&��&�����I�dWp�`$D��$[;s,�TH��P�d�� D����S�["�q�&�Q�5c D���T����;�h*B�X퀑,=D��;`ák5Lp� v���R�(D��c2�}���jŹT�@!�H&D��Z6aS�-9l��+H�0D�*��#D���P�� !�E��҅U<F�c� D��1�h	60��I�CI�'�
��f�<D����˓l�Nx17'M0�P�d6D��#�.�4n.R%�@�I��'D��h�胟g�\{�c��7�(���"D����&�� ,T4Kg�x�*���&D��C��
W�>X��眅2b`��1D�ذ��G����y��Z�S!�8s�O/D��)�j�.K;�A�q��V��@S�0D�#�]W�>��A�ۂ�\a�TJ9D�� 89�&�_�#��pJ&,�/sC|t"OB�W��8M�������LX�"O6dk���:.t�hg��F��bW"O��IO���1��]&HۀC�"O��9ŀ��g ���Y�)�n5��"O�وA/39o�@�����y5"O��(�*_#� j�HC��P��"O\8� ��U�$51nL�}�H "Oz!�!O��88T�އ��� "O�x�r$%+o��R��@���D"O�P�_??`�X��'uJ���"OօR���J�[��ɧ_�d�"O�PB����s���P��:Cj���""O�	ɖ	ԥMlX��A0/n���F"O4uZcg�8��0_NX�Q"OA���@�\�b�E��F$��"OlA����Lb %04+�k��0�"Oظ�6΍�*2e񧊜�6,�b�"O�Q@�A�6�AQpK��`�)�"Ofm�@�E[Q"�,�YL�ٲ�"O��3儂�?A��`3i۲\P8�B"O2% 1\�`��ai����z1��"O�h��;���(���P^�S�"Oh��0��-c�Y@�d��mZ���"O*��i�u��A��b�1?����"O~���H�&L"u3w��5%Ȩ�:"Ofa��^�,�����L� X[g"O�Y ���h|�#�L�#�p	�""O�%�t�����e���z\ �"ON�P5�եz�L�'J��մ� �"O�	��.��>���G�3f�HP"OЭ+ӆQ0.�n█�/N��{!"O�s���@X������x!���"Oޱx'�ۗZ�����S�(i"5��"O~L�    ��   �  �    $   _+  7  SB  �L  T  C_  �h  �n  u  c{  ��  �  8�  }�  Ú  �  F�  ��  ȳ  �  J�  ��  ��  ��  ��  5�  ��  �  A � 0& �. �4 ; ]A eA  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1R��G{��雥|���m�P�K�.�.�(�'[��xB@�/C��f�Z+w�舰N��7�' �QV!B~ACį�a2���'��s�	�R��h��*��Wpxp`�'������ ��ɻԮ��38q�'T #08�R̪4I�i��ȑ�'�н��;���u�з]�.ٱ�'��	����a��iY2
�>��	�'��4���O�Du8�O&tnޭ3
�'��R� ����(n���	�'�D�YeC��}�6(�q��>U��"�'��Xi��)����g�'�
���'��`�� ��,<��0!�;�l(��'�:�#�����Pc�ڟkX=��0�a��Bǀ<բ�$ԕ6���ȓ]f��1���)�Pi ���7n�.P�'"�\Gy��	��d�T��g�+r��TÊ�B�!�Z�)�|��îE�\ ���>ǉ'. ���	6h���FW����3������+񄆳+r��p����G�)����i�!�E/u.����4(,��v��� 1�O&82��~��G�?YvsA���f�ScbRI�<�p��%�^x�,E<+�����b�j��p=!�ႾN����	X�� h'Ue�<!'P�S����4��GP03�K��<��N���	�B)@X�]a�M&bV�E����(����m6H���R�%N\Ȗ��yBA�:|�v�¯�1GZ�(�(Ѷ�����(O>)�Ud^',MЬ�a����l��"�"��X����e�N��@�[�×��Z�8�G<D��B�KY�Ti��Tm�&�{ʛjh<���2L7RL)�+��k�aU]���?�Wg��Q@����U�[F�30G�W��H��\�ɠ)$8��CF%=.f�Ю�O	�B�,: �}
��#S`��P�6}�ܓO�Fz���M4�M3�l5O^��gΈ?wd�l4�c���	X&�9ٓH�U�}I���&m��I�L�?��T�	�y"�)O�&��J���䢙���D<�OF]J5�H��(P�(`�t�Փx�V�xDxB�8����5��� U-��j���RH�<��EF�U�D$*�)ڎ}��I��˙ڟ���B~�W;����t���V� #k����&1u�'�����OV�b������v��]9�'p��PF�2(j ���NO�y�
�I�'J�����z���b����u���qߴ�Px)Ma���D��8��ȃ�Ř�yr�ʙD� =!c��c4"��a��y�+��[F��p�U2cn�3t!�/�y�e��<�\�"�&��N▸�DJ��yR+��q�⎐�M#���S�����YQ�O���O�Ϙ�� Ɲ[S%ԟ*�����IPtB����'�r�'>p�x.�#d�љ��Ӥ6����'v�@":��� Q ��2&�H����F �ȟ����ܤn׊I�T��ld�D�"O�`���#�(�{S&�9o��Pj4"O�͡�I��0)n�	t��0j�5)�"OĈ3�
��}F��G�hެ�S"OH�K�[5`���K�c�AvQ{�"Oxe��d��0��ˉjb�!�G"Oеx�}�����1#U���i�ў"~nZ	T.�07@D-:�x����ԴB�I�"���#��۫7nH1�6Kȣ\U�B��-eD��bV�H�oU*YᇫƴK+�B��9�tع�7�V���Å�^ơ�I0~	��a�L�O��hKsa#8�!��Z�BE��PɁSY2}���[�!��7VnT�aI�1z<��cSeԉf2O���۴##���,SE/�32t�J�O)ED���A�>D�X�4.�,���j���H�@�d�,��x�H��0W�+�i�Qn�[���/�Px��i��1vb,o��*'jɓ[&���'��A��\aL ��&��pU��aǓ�HO؍�@Q�>�Zǭ�3r�b(�e"O�U#�$°'�2\�4���f�.}	��>����ɔ��@1�@��
V �ccc�7u�!�ґB����'k2l�'���x�!�D[!�V�8E��N��`����ql!�D��7d|p������'-�%~Y!��5#��DQ��@�aҨ���Yv!��
#
Di(��=��5�АV!���`�b�Â�.z6P1@�.48!��I]��zr��h�����C1!�߅Us���/_�8t���֘ l!�䒂83>U)R#:G�LD����!�W�xB�TY7N��*���bL>M!��ԬO�]y��%Cq&�Ӫ&>K!�ċ�6[��R��_��cd��,!��6����犁	;�ҍI$�*!�DΛF�$�H�/�ftL5Z���
^!���'�x(T���'/�\i!�"X�qr텏}���2BU�Yi!�d6m�a�� "�$�A���
M�!�dٱM��d�GM~�䫀�3B!�;@V��q�!W X���M�>!����.My��F� �T`E��
!��$t�&�%���[5Bޖ-�!�O:'Pu��U>S�(8Ç܌m�!��ܬ!�Z4�_�D�D2a�Ǵw�!��'f(�R��͡>� Iѥ��!���M��l#��5��չ�Z:	�!�䑌(�RB�Dd��S�m�!��qy|\��L��iD����m	�M�!��C�2��U��7����_>�!�D�v� ���I�"� �Fa�c�!�ċ4V ���C��P����O�3>�!�$��q�x��C
��hӤ��A.���!��5]��Џ�*#�l�4NǨ}@!��AA�܂G=W��Q@�K�D&!���u*uC��n���X �<!�� "0�;��~�` ��IӋ[ !��]�|%4��1�$	�g�(H!�,e�t��2�ƒ0��Y`d�I$�!��t���2&�H�j����@Ŗ��!�$�QԤ@�5Ä�E������"�!�� ����@�&��w�M�~S�$`c"O,a8���N��a�3�R~��"O�yR��Q�ny3ED�VQr͒1"OT	�`!i�`�c��scd0 �"O��bf�G.x@P
^��j�'��'Xb�'�'n"�'<R�'���Wm�zΕS#�66�p�(��'���'K��'���'t��'���'ݲb�A�0P�=`hC"[ȼ�Z��'9"�'���'���'��'���'qz�,�5c��*rM� ����'���'���'���'���'���'� m���đI�\9
����tYC��'���'�b�'�r�'���'���'��H@�&-i��I�mP�Z�Ԑ��'��'���'dB�'Nr�'�2�'f��:3KA��t����
�&?����'�2�'��'Q"�'���'~��'�(�j�%I��Fs�(	'��E�t�'Gb�'���'@"�'���'���'I���ȰK��L3��SD(�c�'!��'Db�'�B�'P��'Y��'/�A��,�3��8��IS/��%��'���'���'�"�'���'���'���#K�P�%�,�2�Y��'��'�B�'��'�b�'�B�'
�< �D%dNj�Prm�� ��E�'T2�'�2�'3�'X�'���'Z.� �쎊ttY�0�+؈U���'���'���'��'�o�0���O��1O^�|b�動L�� ��rg�@y��'�)�3?�зiMƩ���6`H���ǒ2D!�5��g�����즁�?��<�%�iv0Y�E�'6),���\D�	b+s�B��H�f{~��R��,`�cLa�0G�~�w͆�A��ř%�P����іN�P��?�.O�}JA�֍`L���3iD=V��=aq�щ{��ɐ�'(�nz�i�6�XX�6�J����i� ��6�M+�i��D�>�|*�d�  ���6�E����,� װ�.��O���z���(����4�Z��%���1�&L����,��(]�<�K>y��i�0s�y�,&�����)� $��d2o��Od��'66-���Γ��݁Z�	9r��FH�s��eA��3V-����Y�V��c>q�3�֧U˸��ɛ)��%hЫ
�|@`,�w@1x���'��I�"~Γe��=�-��^�f�����&eL��ϓ|���hތ��F���?ͧy������;dK��r)�d�$�\O��@i�������3��D��R�@b�[�Ϟ	˒@���Z� �P�9���.|v��%�앧���'1r�'�r�'a:D�G'̗t���gBԾ&?��R�W�(Z�4'�<%͓�?���:)��ĝR�
)���C?�Є����yy*��'�7U��I����'����[u�ȣ�n|clH�M=3g�= �ݒ2����x���3��@���A�w����r?�ed�<A����Yk6����v���?�?���?q���?�'����U�Vk~��c��E+��rŎR='X�;D�|����4��'��xw��Bq��=o*C���b�N�+,'n��ptn�'9
Nh125Of�V�D*�gM�Κʓ�Ru���4:F΋�K�����Tf/��b=O��D�O`���O����O��?=�U��&���cFL�@�ڧ*Eß����YڴQ�j��'�?ҵiw�'T� B��/m�09QL� 8�4 B!��Oh�b�6Dg�4�IX,b��e(�;O��$U�����R��~!�'�shL�ط�X�)�&�a��5���<y���?����?��I��n���2hPd��U֢ʾ�?	���D�ئ��Ta���	��O}��d�.{$8�C1ێis�O ��'��7�G��I����'�b����@p>��el�T^l��*�O�jL����s����-Oh�iE*k��/5���~��TrRG�z�����t]&�$�O����O���)�<���i����<Z'<��(�Ms`y2�Y?Cb�'x�7�.�ɠ��d���]RS�T���i��*�5]8$b�܁�M6�i�
��eM��yr�'�f,�GΚ�؀��Y�H��ϻZA*\ #a�(��I	a�x���'>��'E�' 2�'E�S+x���� ��^���ba\+P׺��ݴ}5&���?	��*���Ċ��]-w��q�dBP�P$���#3�չ�4.��6h�O���|J�����L߬O!L͓W�r0���L�w��-bՄüP���Γn�X1��H٣h10,26lA1n���,(��mjւ�%i�>D�g�$
1�24F��*�,��7iW�3��@Ђ�'Iw,x�aOO3G瞵�`�>YP��A����d��oZ���Q�R�`�ғ+@#.J�	E�[$
-�ĸ��60�2���CD�Q��Q����^c�Ts�*�!(J��5�"6�Hu�H>!�zT
F�ɿ/��xB��C���0�B�n(��[b�Ò��љG�E2��Kťơ�|����w�tdq`I�Bp �w�#�<|����m�q��t{!�RM�������f��%�����^�&�s�ek����O���Ė;��=B��D9#��uϋ��]��z��ןX�	�c�j�̓�M��j�l��E�ydS�OZ<r�H��i_2�'KR�'l*4Qr�'��'��Oe@��Ԫ�W!�Ţqb��*������;���O��d��I���!�T?�)a�6	��ӌF��I9��n�n���O�9�	�O�D�O�D�$��K�K���	B�X�����צ-�Iԟ�[ m�A�c�b?�x�g�,c�ޠ�Q�� �����%t�@2u��O����O������D�O�˧sx��R�9�!
�-ۛC�4SҸi����H������:�DC>*�hH�%	&�f�R��66d�0n�ȟ0�I̟`{���՟��	R���'F��2l��pb���P�L� &ǚ�4{���<A��D5K��O�b�'�r�-� ��s5�Є�4t3��܈P�r-x6�i��$�f��ɲ����OȓO^�*J���.>w�亵��D}�$��(��B�O����Of�d�O���8�i�S��㜽�� �mE�S�b�OX�D�O��O֓O�$�O��C�Ɔ&��l
.ï6�^X�2@ٶ/���E����៤�	Qy�n�	"��6::Pak���<5>͈3�W�=����?����d�|Γt#���Ocn����L-�"�:�E���O>�$�O���<�3�� ��Oc��b4�L�1r���$��*�CEGz�f�$.���<��CMy�'|n �g��|"bG�C8�AoZϟ��IYyR��?����$�k�A�7qډ�捔�~�<JU��̉'�	�g"|:�O4���<�v��vM��@��Aaش��䀊a�(n����O��_`~�ӊ5 ��q.�3^!���K��MS���?A�/���4�������'�� (�JՕm����JKʸ��4w�|�ʄ�i���'���Oq�O�iE�:�j|�Ue�?RI6���= )�0o�|�'����M�{̓�?i�!]�����[����"4H�F�'!R�'Һ��G=�4�&�D�O
�����n�M�r{ʐ%�[}b�'i�րĘ'C��'��B��#>��
��p҈��&cX���6��OT�O�Q�i>��	Ὁ'">���R 1AR	"��>R��D�bw�$�D�>b1Ot���O��$�<����=r^��Q�P�3-LI*��[7��cЕxb�'/��'9������I?,b|�!��@�ZрX�<�Ph��i#�I�����ԟ�'3��!�s>���M��x�|�����9�
�>����?!����D�O��dX#��;(�
5S��^�D�,��,n �ꓣ?���?	)OR)�iY��BU�X �L�"la�4�B"é{�T�@ڴ�?I���$�O���	)1����v��_Dڹ��VY��s�ͦ����Ж'g�1�ƍ)�i�O����DdzR��`��V�T�aӱiN�	ԟ���#lɼ#|r���e���`|�y�����B-�@���u�.�[ �Q�t�i�^�'�?���:t�	�T"�V�Č59��"�hZ��D7��O��DW�Gj�S�����Nq�3�X�2�2ذcϱ	��n��ฑٴ�?���?Y�'C1�����ܣD�T=k�b�N����ʦW��6ҁm����?)����<y��T�`,!@��(4H<�ܟ�~<��iP�''j�
/�zO�	�O��$
}v�ʲ�Ƹ+���ې�U��Y�'4��'�Zx�yr�'�"�'�D�23o��bФ� [�,�P �f����ʋ7G�i'��Sş���py"oM9rYt	Ke��p����U�έg^6�On
����O:�D�<1��R�	��ň�k��}
'i�q���Ҵ���O>��O~���*i�TZ��퀐A�L�2$�m%5� �?���$�O���1b�?у���d�ը֪t��5�Ѓkӎ�d�O��D=�I{y"lԂ�M�CG�J�09r"�)+A��JQ �y}r�'��V���	�a[�%�O��#U/0����F�D�"4�T8���i���$�<���[]�	�R��Ya�)ڋf�hb�`F�XJ6��O
˓�?�F�-���<!��|�����I�:!���ÕM�< �a���$�<!�E��u�.h,�Re�@'hrNP�'�F����O�:c��O��$�OH�d����Ӻ#r�L�~�FJ.,�r�ヤ}�[��0�6�S�-3�֍���՗q�d�����N��7M .��d�O �d�O����<�'�?y�N�4!��@���4��݂a ��I��ɥPf#<�|��0����[���E��E��Mb#�i���'ra�:A}�i>��ݟ�����<�%�αa��m��Ƿ4�XӖ�ɔ�ħ�?q��~"�f���+V� (sND���Ҳ�M3��:���(O����O(�$ �	)�`�(�79*�y�@۪!x4O��5�������'yRH�Å�2E��HC�֡q�|E05�7K��I矄����?��h�~�Z��P-"���2hZ��43���(
��(�'5b�'?�I֟����q"JA����w"̆.=*ժ����	ޟ ��a���?!��0-6xmZ� ٌE�OTf�*��σ]���?�����O�$Cѭ�|���nƀT���1x;(�Yc&��"i��b�i���O.�Q�R&;1�'�� Av��$@(���Y'D���4�?�+O
��N,Ds�ʧ�?�����Ψ9Ԡ;?z�H�M�9fg�O��D��Zw��ʘ��ɗ�+"���Qc*AÒ�*��I���@ ��ҟ���ן��	�?i��u�"�1jh0��&+�Qb�%�����O(ŀ�j�4Q~1O��PP�� �?��|s��PBEp�i	��b�'Z��'��OG�i>�	�H�h��n�bLH��!��Tކ�B�4*A\<��c�v�S�O���11oʄ�7G�D�6t��)]��6m�O��d�OXX��J�<�'�?i��~��A%::�k���=pP���3EӹF%�c���L�ħ�?I��~BC�
4�8��1H��e_�8a�'��MK�;&,-:)O��D�O.��&��"|7�#㯉�E��� ���#�2��%k�p~��'�X��ɂN \�ږ�hD20����6h��R��ny��'@��'��O����8�t�23��g�9��]�1)f^+�X��?)����D�O����#�?� �$�c�A3r
P,!e(�1t"2����iw"�'�����OT8"$�S��&��<?���J����:
��u������O���<��'9|�:/�L�D��'�8`j�cީq�.%�3hݨ7�(nZߟ��?���9|Cc#_�ɸ�F�T]���V@3~��6�O���?�1�����O�$�����A�~��1`"��87Be��
u��?��ㄘr7��<�Oi\��G���
���׌`��'���Z�]���''2�'K��_�֝�Q(6��-��x����g�U,B��?9��	�@<�Q�<�~���v-v0{���6��r`�_�����ߟ���������?������'��D��N�'�<���3z��
�Bc��9
Qǃ/x�1O>	��3E��P��[
A�X0СO $�La+�4�?��?�P�ԭ��4�.���O��	�"�4��0'�.����"C�^Sf}эy��X��֝ǟ����T����݇���S2�� IxP�A�۳UV6��O���4(�<���?q����'�v���<���+��2���ʫO���tD�&8�Iڟ��	My�'�:�0��5~m�TNޙ"P�!yV&Y$��	��P�	���?)�#)�0b�C�Eֈ�B.�>l,8{Pn�y��t�'���'��	ԟ��2��C"�)�4�ڐ���=3(�@"�����Iٟ��	A��?�$mB&#v�m�)�ֹ��h�X��+��,tz��?1������O~ j�|��'�P�"���w�b �7��]k.�h޴�?q�B�'I>��sO�ē*B4�P����g
~���_�e��o��ܖ'��*�)�����	�?)�����>,|�rɍc��tJG���'�rۏ-M�y��H��0�I�e���`"�3}�����^�(�I'y��=��ܟP�	���wyZw����j* �<)5CI�Id٢�OR��XJL�����	����Hac��P�1� Й/B����!["�'���'t��T��ןT�FC\�!ڦ=c�]1V���D��Mu-,�`H�<E���'���)qa�9h�0Cs�"���	��hӨ���O��䅶2�0��|���?A�'':`a�*�;ɶb$/�(H�U�M<�ɞP3֩�I|J���?�'�Ȉ�Rڝ���#ZKl%iܴ�?%�Ӹ���OF�D�O�㞸��˃	��zRn��f):Q+�>A���|���'�b�'P�	�4����!'�Ia�"֜c~��q�Nݚ4	\X�'zB�'
b�d�O|l����!Knݘt�+#� YԄ "��E����	ğt�'>�f%.%�IM_���6#ʮIlHH�f̟U�v�'�"�'S�O�����N����i��Qa��1HI�<#��4
�4�O��$�O�ʓ�?�эK���O�0��@&%}�y0��Ƀr��)��l�ɦ���t���?�EN(Y�4l$�ȲE�]��91r��)lc��Y�od��Ĺ<�0HN�*�����Oh�	�,;�r�HaN���E�*J;`�0��>��6��2v͚{�S�T��Q���sUr��8�fE����O$��G��O����Of��៌�ӺS�DުB-pm�u��	4�����F}��'4D	����'����O�1y#��qN�胰�&pL��4k.����?����?�'��4���d����"�@>+D���V/	��Tm�U��3�j7�)�'�?!/ً$<@Q3�/����
d8��'O��'f��ʑ]��ן�Ir?�% j����W�.r I�q�A %=1O�!��!��S䟌�	j?��/.b���J�\�Xt���Цe�	Z60�'��'-R�\�6��LQ��9y�����!�"K�ɹ�T5�c 8?���?�*OZ�$�z�ह`eߤ.ОȃҠ	Uꞁ w(�<1���?q����'�bDFVK�F��	������%(�$` �
����O<�$�<���b�)�O_~����[a�h@`�6$��)*ش�?����?A��'5X�8WG(�MCIK�b����F p�Q�+�@}��'*"�'h��'%^A�Miӄ��O�1��	=-kFDʆg�kk�}HǋǦ���̟(��Ly�'����O;�ɗ��ё�@�a�Xk�h�+x��P+�OF۟�������I�Fd��4�?���?i��0:��Wk�4'XHI���:)�L��C�i�[�L��2���쟀���ܴd7�h��(f
��X���dS�(oZԟ��ɞ���4�?����?y�'�
��WZ�-3))?�������% 젢GV���I�,���}�i>���y�cM�>M��8���J`��i�6�Z�Fv����O����,�I�O����O�X+Q�$E>�n�=���ܟ�M#!I\�?����4�������'�Z A�>J9���;Y��mZٟx��럤"Gj�M#���?!��?�ӺkM*T��4�,�i#,ׂ7�"��A9�~ʟ���O:�d�>�q�fL*4P��B�c@n����+�' 4�M��?Y���?�V?���-�>�a��8��t�p�S./6�m8J3ܼ�T$z�X�'%�D�'+r�'�2&|/ K4�ɽ��Ç�P�^��8Jw�`�$���Od��O��O�I�4�aEιC��Uh��B�@�A���,���	ğL��ڟ��	�D��ğ0��Ñ��M3w _c֭�$כ3.z�@a�A�<ߛ��'	b�'8��'�����P94�>�c�H�$l]�厸;L�XB����M���?A��?�uS?��Č�M����?����'��sd��,I^�c�h�y/���'q��'���˟�C��q>m�'�6$)T)Pt�!p.�.���*�-=�2�'���'؍Z�Gp����ON�D��
� �a� ��$)�-����\hw�ib[���I��~�����6���s�P`���[=�����	�8Z@�	�iS��'2�4�wgh�"�d�O"�����	�OZ��uK"/ĕf��q��|��
�{}2�'�l�B'V������O�T+^�2�c�$�@h����A~��7-�O��D�O��i�0�d�O��пn|$<k�d6N�L��@��o��5�$��������������'9���3ʠZE���004�}��av�Z���OP�% ��n˟��Iȟ��	���]�wJ^�� ����Q*�޵I��7m�Ob�#����S�d�'lޟ��+A�8:X)��&��E,^���iMHZ�o�6M�O����O���OZ��O�XbH��"S�}W�U�o�|"d]�4`�&l�h�'E��'��]�p(��xe8]�C�)�ʡ#�FR!i��O<i��?i/O����O���C0T���v�R�I�"����G�$CT5O&˓�?i��?�,OB0�J��|: ����4��K��J�a�w}b�'>BS����ݟ���>Pq
�A�P!�wϘ,�Dp ������'�b�'��W�l�-��'V�p,�⋓��Raxg�Ro��P�¶i;��|��':R�N��y��>	r�V;#��!�G�:y�<*r�SӦ��I��,�'ŜU1��=�i�O���T;)��t��F�k��� �G�3l"�&����Ο�:��r��&�@�'%|��Y!�ÇXs��(c��W��%n�Wy��W�26�[b���'6��N#?��[�]�� N�<�*���I�I1�{��$���}��N�/tL�f&�Z�v ��ݦ�A�D2�M{��?	���1�xb�'��Ыuo(#���+�#�-�Ĩ��k�������Op�O>1�I�ee�S4�6P����S�<}&[ڴ�?���?��.��H�'��',���@P"HեZ��
s�C4A�6�|bg�0j��d��Ox��\&���%K�(�
 �vD�c�^�l�T�P�X��ē�?��������<8)"��#K,I��-`�%�o}�ʠcZB^���I�$�Iyy�L�]�2UEdY�3B]ЭP&|�RE3�D�O��(�d�O��$͕n�v��F/���cV�[Ɓz.�Ohʓ�?I��?�)O���a��|*!��I"�L_�4(dTKA�b}r�'�2�|b�'��d�����D���Hg&�0��{�����������(�'-B5���?�(2 H ��P�W1B�+1"GK7�IlZџD&��	џh�Ň�ȟ�O,!��ߋd.�
#oX�dA�	���i���'`剝I�0HI|B����VYvAӗW�i�����2)�>��'S`8����S��*I�T�>����i���W����%�+O�e�U�W��=P����䟪��'�`,p2��n|m�3$�^z�U��I��,��	�(���Oj:�*vHőf�)�O��r�8`�ڴp1&����?9���?i�'�?I����]1 �y�!�8\:�9e��^�l+�쀫�h4�)�'�?��e�
1��q(�v��3���' r�'C~��!�4�F���OX�¶I�y�R1ơ�$+l��i���La��?i��?IZ��9aԡ ��X U�_,��n���0�S��Xy���~j���jN�����B9.K2�Yw��{�=!�V��#	t .��?I��?�/O6y�JDu2XtZ�ϋ�V[2 `�Ҕ`���%�l�I��('�h�	����6l<b�0�0ѭQ6\�@�I��)��c���	�����Jy"�Ƕ<L�擊J�Fxa�(@AH�mҜ+�Nq�'�'@�'�'̶���OF��+�>Y�H<�B���?^L8u_����ҟ���iy�
o������=9g�Qx�Ŕ/$�`��!��}�Iz�	x��>d��b�����T���㆟^�f��C�v�*�D�Ox��LG����'T���Ζy�Tx
�2UL�K�ɑ=e�FO����Oj��~RFGʈi��e�7J�*�9!L
�M�'Z�ءKmӜ@�O���OB��7LjU��\Q�D���5���m�<�	�N¢"<�~�@�8�0��UkO�< ��+���kD���M;���?Q���ZՖx��'�pZ�!��jkѪ.Dpy&p�V��)§�?1��h4��!��!@����*�ћ��'e2�'>��t҉'���'����,T�$	��ޥk�0 �'�&1�OL�#����Ot��O�P���Ȉ)w�^�{;ZѠ�	���	:�� �M<9���?�H>�1�@]Ic'�,a���bP�6ک�'�Ȍy�'���'��	+qk��Y�LƵD�^<X�`ߘp�z��� �ē�?A����?I�:��3!��;T鲤��^&ɰՂ0��x��?���?I-O��aF
�|��i��&褭���8���5���ݟ���e��ݟ��	�ib��"��e�*(�0�ua�� ����'ub�'�R�'���{��� �ˀ^[�Y�r�YB0i�'�,�M�����?�[�XU�>�#�ƽ)�x-�b���7A��*���֦��I⟔��؟�z�f�M��'g��O$�A2�"�/wl�d.9�J�Y�H*���O��hN��FxZw�������	R�Is+��HK�{�4��D�PشInZ�����ʟ�������ƚ�@6# �h�2���تu�x��'ў\�O��I�E��h�G���2Op\:��i�J����'�V� ��RyBV���� n ʇ��}�UY�A>����սi�DKR`՘�(�V)�'wa�$�= �.�	�
�c����&�
>�~r�K�P4���7k��*���p?YS��,�N��hA�}�W�G�W=��	�ꃊ[�>��Լd�T� ]��Vx�dkF�h��֪B�C�e�rw��s�_'q�`��Շ8���{�ҟ0��%rf*�Az0�h�k�moH-i�
)m�j��d�Ѝ,��I����^�l�0�߉*������0��0�̟\�	͟��	�|j�����P�'�H$�#���h��S�=w����؋G�Ԁ�F�1ɸiJϓo�<$ꥧ�*8�(�q_��I��^:Y��PH˫�TPx��� ��<�`H�㟘�I�)G�����گ�܅P����QF{r��'��L�F@C )C�HBAҰ$���"ړ*3D�C����`I��!�*� w��<͓[���'��.$��
�4�?����	F	0غTG�
i8��A2�(�c��O���Od�`���,T�'��'".��" !XgT!8��Q^�Dyr�#Vn�a��8ܒ<j�넫,����A1dyV�<Q�g�埬����Ip��L�-@N�!�Mþr֎4;P.ʰ����s�ذd�aܶ2���8��>�OHh&�P�6 C1KM9���Sx�qҒ~���ږ��D�O�ʧ;J�����?���9Z
A80��
N�
����M����@7��,�'��^�Q�W/��1?
���ΘϿ�P��#Z��̑GŒt1����%�����ƔN2l�H���N>"A��M?h�~t�������wp�A��ӣ&�s5��.��` ���$�2�'1�)�� �����
��'�N%��5�� A�!��F�Ix���`'�;D�TE��
ӶE�1OX��I���t�'�ls���%R�ޭi��ùt~�
 �'o��d��R@�'���'{r�s���	�x�ED��2)�'/ҙK�8�ҭ��?風�H�b!�G�����3�(3�l�,ո���_(�E�ӟx��.Hq!�)G2��I9���e-�M�Hz���mP�I�j��OR�=Q)O�%�`�.j��}+���(f��Y�OH��83TT�t%�8�#�iO�[g�,Fzʟr�\��D�i�ؠG7A*Zq{�2ERYp�'zR�'���ؒ1���'5�	)�P���)��g� bS�Y�c!K�7�vU�e�]�(��$��ب혔 Q�?vB���С�>SC?2)�q�3��U����?2	�'�R	����/�r5�sb�,���
��	z�'>�:��G�[R�	���ڠ&zA	�'<�Bi\!���Ek�m%T��'k8����K�0;�tlş��	B�t���Rwd�QAn�W:α�����N�@��'���'�јB-y��b�ʧ�a����E_ �ړ���uDy"	� r�?�Y��4���2��L��PqUd6�UGf��	���'?����L���0d�0�VdJ��,c����I[�S��yB�'y�L�iG!V_����8�0>՗xb����L��!� RG�L���̈́�y�'�S�6��OX�Ĵ|���[*�?��?IA���%�b��n�H�vr��CHŵH��8&�ʧ���?a�%���S*�Z����LJVv�h��ɧ�����o(�T��E8
$]C��n�|��V�'�\6����	��?�va֎րSReԽR���7�X�<���>q#��6?hE�A;5���2���q�'��"=�+�)���ێF�a���%~� ��+�O:�d^.N�.�r�O<���O��dM���?�a�M�&�	�	�6�jq��+%��д�O�|�|0�z����g�'0�U�G\��$Ȉd�-#�lL['�S8}N�k�X.J]���)����䋏EJ���I�7�L�z�B N��d^ N~�t�(IDz�Y���!K�k��@kû��p��/D����e��,9��TÀ��y��%�HO�Ky�h�d�7��R��цE~�"<9v$�T�����O�$�Oʀ���O��Dm>q UCM�� TORQ��mc���Mx�iR*!	��1���'?\\����H*��ӻ�iB*��oQF��f�W0w�`i��m�z������O�uor���	�iΪ�Z W�P�i6|�+ߴ��'��#}�$X�4�,M�9��M0E�U�G�؆�u<�%J�(%DN(�ҧ�.v���`�	Cyr ��_�6�O0��|2�kS(���QbT>Jg�e���:U�������?��SY�p�n#+��O�$I��h��
=8˴���.٣ ��<i9;,�Щ��J&(�x%8c��+.Tz�K�-���I�>p��C׳YҠ%�I�i�J��[զ]�4�?�.���q���qS�d蒡�(h�Z�ؕ��O��"~�x�N�9�K���"D��d[�p�؅��*�ē0��%p�I'h�t=8!��9O�p�'�b�'�ybg�x:�Ā-~D8vB�y
� �-� e7wm(l�7�٤"�@eÇ"O�xS�ND!���K�
C�	-q�"O͉6#���I���B
�Ÿa"O\����W�0I�1i�?�
���"O���"_�b��P�'�0MJ���"O`q�v��
v\�QUGI�Z&��k�"O� ���Y C�49eQ.;��J�"O�����'ؐ��i��x_�x&"O�p7��<_�n(3I��V*"O^��C�>��[ӎ�6_Lv"O�}Y�NMĜէ��&O���c"O�4�6pS�,�?|�-�"OZ�+�e,0�j�5E�:l��;�"O��S�G�8X�<��	]���� "O*l�I��s�M�fdD!N�]rU"O��ir�ևP)VNT�  �]�$"O��3����4#�X��|x�"O���ÁA��&��D
�L���2"O2�h@#_l�Վ�1A��-�A"O4�2b�]��ȍqd��4h�M��"O�PAB�� �D�sA�y��"OB9(B�y����B^(����"O:|bE�ٰ��`���$a��H�"Ol ���
r�u����&1��1{`"Ob�{7k�&Sb�*���*��q�"Ov�萏
2P	qB��w����U"Oh�r��"i������?Xx̵rR"O�D��JS�8p��-�X�@�i2"O,@����%,���g#�8k�f8)f"Opd�gFO۔U�i�D;�i�e"O�H���N�b� )�Q1vP�a�S"O* #EK����!���d=��"O2=�Q�iT�1t�B�e��"O�5� Ħ��Yɠ�Z,X���"O����Ŷ��i���d��"O�IX��C�y����4b�$�4
�"O��@��4
L
��vaݠ[��"O�Ty�`ҍ�����
��0��d"O��A��\�W�d�J���@x��"O�5�vk3�PP��
����"O�4��.��d8�\����7�5�'s�u�q�י�J��h�0r�K�=(X�T�w��8U"OT�K%眕���@�� �w:�0���s*9ӰBT�Pz�yE���֧Y��-�a�ƎHg�X�W��>�yB�G2U򈬃�)_4.����];�h���8|���:��D��O���g�̵�ib�.O�$�$K�"O�)#Ԅ�))u�(:g�6&<`&n�0FE���ǌ�w� ��퉐5g��Xs)��ˠ�= ����ĕ�SӜE���|ϔ�m$k7
5֤*6��՘��"\�RA�r�@��?�����MM<����ɫ.�x�/Ce̓*�h�Ñ/B�_ȚT�'����&�_��J�>:B��S��%<bx�$O+�y��D;�Z��[�=�d�fГ+#\�a�\4�U�gB N���4��3DG��ݗ>�e��g�����	¯o)(ņȓ+�"���M5���El_�jh��!S�8T���H�Z�&p�Q���/�2ԉG�7,�n���`A;<@�
W�F"���Q/ؤ�r4a��e<$�36�ғq��P�7�&�Y�K#S*<����0h����0�6��AI�E�P"?)�IS�}Ą���/Oʲ,��:���FǏ�	�<t�p�˜+�Y�"O`<�.�$l��ͻp���v]��!e�@�_�ބ�����+��uZ�S=(_ԉ!�lF�m>*`�#'��C��=n�z%˖F�[}*�P���@;r�ႡG�,�`��կ)Ul�K0+6��dʫL{n  �·b���H%� �!�dڋ���`A"܍\x���fR2C8(c�'�*R���ʁM��&��	�r!t ��k�r6���a��s�������5%�,�v�i�Y٦� �h8r��&	���x�L�9��s"OL�I5
ߊ\���S%Ǩv~�0�e����!�Z�e��cBÒ�})F�Y��IH�"�蘁K+
�����̃T-!�Зd�i��Q�
�ԕid�æ=|K�)��V��l��r�\��6�3�I��f ��R
�(��J��������<��=���~U��d�38��h6�a' M B�_&-�68�
�&C,r
"lO(L���YV�ȑ`b	�3�!c�d�H�� a��L=� �a�<I���?-�'��Y~9Q��BY�n��J$D��I�gT����.3��9�7dT��%�7�a����s$�8�3�>%?��g�fޅ¤O8$���X�h���@b6g:D�<�	<Dt��A  �d�.�0F�3?�q� |I\�e�Ї'�<�����n�'8���/D�C���,?�05���8��_M.�Bo� Vx���Qr�d��d�%/#FbAi��
�#3C6�O=���8 ��e�G��:��ڦ��6X���آh��;�0�$I�>�J?0�Ƿh����Q�n�)'A D���\�rc�$��dрh_�C�
��s�s��5��<òiB�����:�'{F�#�@P#؀��T�,���y	�'�58V��'6�6�9��<aGT���#�|`gf�L�rL�!:m�4F}���n2f-zPȴw�n�c�E��0=)l� ?ΐ�U�G�^\t1��l䆘1F&��2�����PS�0�Bfx�X)G�Ъ*�� �O挐�~�4�W1u�$qPm�/!g�բ��y�a����	�~QCuP���)�4�O�U7�0S.B"*�h�X攲c�Zq+se"%���V�e�N(�����>�ӉݩK�l�#�kʌ	��,пȼ�`��B;����h��<�ׁ͉�O`��[�M���O�J�]Z%���C����A��2)�����"��b
m8 ?Z����DE9����N�-��Bԉ�z��D��}G�$��@� ��m�CBU_k�)��|�ȟ�4E�M�l0#�J.m*�p��@@��p<�ńH
q0���F��3�*W\ߪ��RhV�@���u�*rT��ʯk�ڙ��s$*VW�Tj0��S[e���1Ñ�D�ұ!���l^0c��#���(� d�Q�J]�iI !m����C$���c�[�j�17��e��{��)IQ�'&q'�ЈQ���s�i$}r�Ͻ.�t�됏����p3J�?����E��Nyhؙ�B�-�yr�ߝnUt���F#p�ƛ�e�4�T�r��?V	��qA��=�F�r��Y�m���!���8W�*��IR����JO�"�B���D_?�$�	5���h"/�.?���QuFR61��S�'�RɰwDN=�4��;Rj�beM!|:`�DH�2V�p�'�'���Al�Y#�w'\��q,55�����<�b	�w�E[GrQQ��a�� �8�L��)�<5x�~�����J �,����kH�p��|̓+�H�Q��.`Xx� J9}"��9Tа�"H�Jlɛ�ܟv��S�H�^J���$̇�m���k搻q������>9 ���/�m��BʴZ��e�u���C����I̶8����M���d�?�5�4fKD��#$��v�}�'X�
_��c�L�~ʒ�*Si�%1�����*O�y���J�NJ���t�x��斓�O��J�I>ͧJZ�Q5�<0l������YvjN�aaXՠ�F�w�0H�Ǔy���cQ�R;a0ވ����I���5K��<��$���o�:c�Xtb���ʜ�0a��"f��}��3K���a4s�ty�nUe�L��u{�fEnp0���?�'�t���\�?�<0��50f`�@�����wF�#Ј@Ykd�'��ɐ*+�Uᦂ	B�2e��:[J����M5.��1#�!COȡ���pq��Q�	�T��NE�3�i#�'m$�$@U�kT�:˓^Y��X�*�<)൳�B��K�������Ƭ��7K.����r�L3ϓw�.���	�2��M1����%�=T�Pt���
"i�X��T]�堤�X:a֖� ��#T�2��iB�V��}hU�|k1O�|jQ�<<�Z=@� ,^&�i����y��<�N�]�������"YIqO|Q�Cf��d� ����0"��0��|2�O�N��Q�V�L\�¢^8e���#�T)\Ul���ԥm��yR�Q)c�p��7���E;f�ff��0�W�=�(y[�kF>*�����ܽ��[�B�	":�����*]bܼ���@.����+e���S����	�����҈�0=�FKʤn�杒Z/>�aC�ы	��H���.c����$I�c;���ƫ��p�C
(\��%�/�b�@���'��y)c�(t��]���M�a�PX�4o��@��KU��1ı�"~nZ��b�����1��i@�GK)E�VB�I�1P�jġ���F9\�БC�	��6F|��5�<@ᴐ��4P�?�A#K�-z(�`�
��fy����HD�l�Gh�4�'�W-�"բ�����^�k�#�\��}��D�A"HI��Y�'m��ᕃH�oy	avZ���7팜r�J���O\
U��Q��P(�?)��:i~ĤR�P�L9'�O|6���P��`މh�oؒ���V#��
��P�0?9��^%�����qz�}�3�H$XR�Ly%�S�z� �B�'�5��T}��iP։1��h�^H�Щ@'���,O�  Q�
�gg0 ���+!��P!= �x�'�\
�������ɹAL�c��BX� ���n�n,C�M,r���e�}p�����4Xd� $�@�F��+�x�'":i��w�9��yn�XZEs�Z`s3�ت3A:@��n��P53�wS��8�3�i��@E$�h����9]�aY)Ģ�G{�"&�`%�BB#�AC�wT�uSp��3-�t����w!�D�O���;�	i}bɕ�P�"p�&���Ol}k5AQ5J�ܱaq	-I���'T��`E�>�qh�쑝m&)�B�v�.@�a*�V�����cR
dJƽ��/�fpl������&��ybṟ�B�l�;~R`j�[��4a�F��3�;=.��D��y� S0cZ#p�`��9n$�<�%O"!sF��7�ָ�5��'A��hi�nȨZ� ���P�>��D[�5�F�hc �E��ˉ�$/B�CN�+�l�� H"A��h�C-ٳ��q���Ψ(� b��7"�@	�'/�%�^g��à�]�y�`�[�*P<�ўD7�ϫ)�IhQj�x:V���1� �E��g�f�@�/� DE��Of�B�'� �1Of�pF@)�����IΎ�	0m�(22��ύ��d�U��E!�+c��95��|��LQMVv�3Dˑ�qhD3�C?
6��USlY4�re�Vc_:�E|Biцt>�`h��>)�ĩ��!D�)AZ82�㈡R[F={�� ������3s{+�aܣW=��?y���m�W��h�1�j����X��a�a���Oؔ���H(�)�� ;��n� ��cR�ׁ2ۊ0���dK1f�PX�W%�.��dG�8Έ$�� �+nܩ����T�v�����P
β��0̅:*0�9J��wN��S�/�#i��H��nr�!�|@��.��#����D*扟%���YS�Z >>�S�ɺ}T�'��}��F�;���hI�w�]��ׇ8*�![�ǐ�
�T{'AL$D�xp��4/��5�Ʃ�8��E@ �7?iH>�T#F?(ޚ�%��.W�]G�� ��Ts�xэTy �d�q,�+L$p2���7���&Gv��5�  i�L�p�s��,�0��%��yf L[�i)��O�!"!M���&�̻(T̨�B�4����e�BL��B͜oL@��&��$�|��h[��m
���\�Ν�G{����QL�'X����օ,\xz�OYN?��dP�
 �a��`3J��j����8�4n��u�'� H���|Zc2-���S�5Тhye�M�OD���O�D���$_=K#�Q��h��L��0pV�c@�Y�)��X2���j�J c�Ft��FB8��.ʧxn��a�Գ%7�� �%��. ��� 9[F剷~�1̟�,�-����F��1)B��@J�1��$���@B�[�ay2NP���{�b�>e,ٻ��&�y,E�~����� F&eB�n���y2�E��F��'
|>��"�;�y2%]�f� c��&t*��R�ϋ�y2 Bd<pY!�cB�=T�д���y��4!
������Nl�T兔�y2*ۣ�n����Ӯ?v��S���y��^A��ѐ�c�05��yc�і�y�h�V�F�q��O"4ԛ�J-�yB��&��0d�<l�a �V��yB�W�XG�I	�5B0�/P��y�f��#.�}����txY���W��y2�W�)����#d~\��,�k�<���`�F5�R�C�`{^a9�LO�<�D+P�q�� �HT�I��@�Qo�<9tHޛ(L��)7J�� �O�<�JE���bt
��D��B�<�ኝ�A�^5����Rݦ��a�B�<�v��4_s�-�� @BI��,�u�<�uG�5/j��*[*@@ڤ�]o�<�R��%2D��@��֣[�*$��^`�<I��
N~�ȲF��"�<����[Z�<�IW!te���7��Sr�4`�U�<1d�n��(j��.��I@�Q�<�1$М	�6%P��?�㶍t�<��'�#2�9آ�}s����\�<1��J=��(�QeZx��y;gm�W�<QRlC�`�F�5��N��wf\�<a5ÉPTƙq �޷Y��](ע�`�<A`���}+<	ie�v_�(���x�<A����KReیyy��3$�r�<�dKĭ���@�釾-L�	���k�<Y�lC��e�R-=G)J�37�Ck�<ɗh�`�@��-U<}�ŋD@�<� ��ÈV&Z�p�"�_e��$�b"O���%/�U ސAqW4U&x���"OV�:R�T�%�`	 ��,-t5��"O�x��05���{f'��>��� "ORix�/�+P��l��ݯ�T��0"OxUz��Oo|���N\Pǂ�6"O�8А�׸)�DK'��OƴM�q"O`A��
�%"F��������!��"Obr�+��DJ\V�F�L}�7"Oh��ei 2|�BZ��H.'v�)� "OȍH�%ג\��Q1B#g`E�"O05���9.�}�UƑ`����C"O���3�?�8�z 3:4��"O�Q�R�]9��|θ��Q"O0�;�e�`bX�!�Ű4ZD��"O�-�ӥ7�`��+�7��(A�"O8�eMO�3���0�K7�RĢ�"O �D̓m^� ࠏ��P�"O�l@6��j�r��qOV2VѠ��'"O��aG�Ҁ;�ht�"ϑ2n���b�"O�����7'��;b�K�n\�d"OL�2%L��W����,Ǹ\��|1�"O*0����Z$��g��'�&��"O�MKӧ�3u.Vpu��?>��a3"O��p�V���|�$�%I���"O��T,C�� �U%��T�3"O����o"�y��E!� �"O��e� ����@�Al@�'"O���I=[�bIRo�5��%"O�h[q.�7M��� W��=0I�'Q� KM,~%,0���Q��bI��'�ƹ�BbR�Xp�}��M����
�'���Ve�&���a�=(�'=���借7�lb��)y�Ji��'�`P�KL�l���� Q�j2�l@�'k^ �V���>��u�a!��i�9"�'tH$��[?+Ox�:���*3Լp�'��D����[v�{���3`�mb�'�"���ͅ;3H�����#ݐ���'6r(պ9(t,��-��J�Gm�<y�&=N�0eC�$?�Y�q��l�<I���y'�A!�ޖ`���l�KQ�<9⯈�b�%[���|K��� �D�<�q	M�<�P\�Û�'ܖ�*��@�<�a�� s�z�ט�2�1�Z@�<q���<w��Q���N�ּ�w�q�<'/@+�,q����GwD�b l�<�t���$�mXv�Z3$�pC�k�<A�+�u2�!�Fj�&�A��p�<q% ��T<�s�^�(�pҥGh�<aa�J0$�X�p�ǐ�B�a���Y�<����@�<	2�خh�|��q�p�<���jn23 G�0@��&l�<����h,�2���A���C���d�<�uCO<b%��Ia�
��0-Y���a�<A�j��X#�]�B�K@���S�	\�<!#,׸j�&�ӓ
���`��^�<�SA_��H�0Vă�H̒]��f��<����SK�zu�p��s3ҩ�j�
k�C䉋zc�t�2MSv�m�PD��D��C䉽%_.�)��L'���+�W�D�FC�Iq���)��1x�d��V�;�bB�ɱs��`��"��9 \���S���IV����̩z၄/�Z�r ��7`�-�s"O� (���A�v@�/�A"O0ȇ ݱ%֤H�e)R,!@5"O�a�A(	�իHZ
���w"O���J̀q�A��:R�bQK"Oε���K��r����]%�j͐t"O�	��HY�s8|8�+��I�~ܹ�"O����ϰ��sv�t�V�0�"O���pDϙ"�h� 5�I�9Ɯ-��"O��ȳ�Ȓ^v@�E
�Ɔ�S�"O�QȊ���\x$h�l~PY�'	�@�d��:`D!�� U�
�'�M��ɔ�Ԅ|rR郒%�j�;�'��H������,�Ҋ�`���'aXõ�l�
���M�)e�h� �' �E�p2��5:�A?]tRa�'�&H��%�'9$D�W��@kJ-{
�'z%��K�!bة�-N�	� ��'T* ��	�%<�P+�#�nX���{��)��X:"Uw��=4.���n��|+!�d�+	���J
"7PI��N��S!��If}9����%&́���"�!��&'Դ��T�2H�@Ϡ�!��ŵ��9�LʮHj���!�<U�!�$��ƈ@�'9=�zX���ՕZ�!�۩5��AA��5�By�6C�I+!�Վ,H 0*��%�h��P�ޓFy!��Ƀe6 ��Aj�#(����j�0XZ!�
W;F����.U�J�"ǀ�"n2!�$2 *i�O?���ҏ�!�$ܑc;q2AZ�"�艙�N�,%�!�$X�z�w��2t��H�1n֓4�!�� 
=���Җz��Уv BM!�$ۇ{�\�{s���dJ`AV��4!�d�#%6�q@��:P�쀗�8T!�ܫWAt}��ƀ�t��	����!�I=8k����x$��N�!��ŷB�Jș1�׊}�(��e�8yc!�D+$�xl�-Y.���>�B�I/� �2���p�����)ϼC�I��@�3��M��L�4N�}H�C䉵$`;�ܩ'z�@p/��dŮC�	o���5��6 ^0M�$�ٌ\G�B����N h��i%�N��a�g=D�̪2� o�P��F�ʔF�ZY+ &;D�pj��*	`��f�;$P��s"8D�XЗ�X:(L9��Đ�;*��pH(D����I9G�Px�䭏��<}"w,D�xyT�ɔ)R�\c!Fθ�-Q�*D�t�PJ�t����o��=��PHţ*D��X���*
��8kC�|��P�'D��zUM�	���ش�\{���cD�$�O�	�WMD����V�d�x�%�)	�B�ɈE�H�C�)���D�Et�C�	&��H��͑�5�����8�B䉁 r�K�N	�R��f�)
�C��ߟX�ALa���:�Nm!�M�!�|C�	x�A��"�/s�H7M��u�\�=�N<)���Oĭn*�2�"�(y�eK��y"葇lo@��K�?r��0��C��yrlT�a`m�Q)N+G��P���X��y�ya�qJff�w��)c��wl!�dͷ"���K�旨a���k�*)�!��O`L"�� ^/���\�)p�"O|�"��ӫɰ�8�����Ȳ'"O� @P)���F��c��0!�����"OR�谏S/�5g�� ��E�"O(�Iq���,��|�w�����"OX���t�X�����j�T0r�'�1ȧJR-�Ҍ��E�n^��'!��c�
�Rrvjߗb�x0��'Ѳ r�%Lb����
۬1�'��c��/ �RIIgH){�';�3%K�\��u����4zU��9�'���`3�̖v�b�X7�Q�k���2�'�*��Ѓׅ3�p�����P6&��'(��RD�X3i�f��HĠ�¥A�'g�14Ƕo!��rGU4i���
�'�,���HbRh�s�Q0&6$�	�'�B�s���R��s�-���	�'V*)1V��2\���
S�Z�����'@*���y�{�R-*�z��~�<���ъZ�$0��ؔb�b���F�<9�#����w�|ul���Di�<��ݠe+��#�\�B�`ɡ�OF�<���8D%F�	�&�ζr��a�<�p���I��9��Ѽt���)Dw�<����!n$.4�B���{�9P���~��O�ʓ��O&�C`͔��a�l���0 K2"On�;#L�'K��ab�
թ )haJ�"O��Kb��4�1ɳj��=|ta�"O�Ir(Z�O�^�[W�@F� I��"O�K��|��6ҡ.�V4J�"O>LnD�/�t$��PX���"O�i;�$����Y4��{�<HC "OąĆ>_�ܤ���J�]�@��C"O������Mc��,|&QJ�"O��r`<:���#Af����E"O8�12�p�h�3��]��<�B�"O �b4GI :�B��mT o`-a"Of�IF��3Jf���'�L&���"O`4K�(�'�ddy��(8u��p�"O�iP�Z9s��@��Ǆ~����@"OnX���$S�����8����"O�ܹ�E�wъ�Xb���N��P�#"O�)Z�g]�A�D>!�1�"ODEꡩ�d�B�:Bʡ�����"O޵�4fC�{tD`G�X��L��"O���cR:��pᖅVA�P��7"O0�0��%>��LK�� =�6L21"O|Q��䆞&#���H8��hy�"O���Ū��vnY�N(T�`��#"O�Hde�!���w�ŤM� В�"O�Ś�k��wm<��w��|�|�rs"ORT�0�݀i	p�R��h4.���"Ob�2�J@�`X�C-U�+U"O*�� I�_��I�CO�/�ԑ�"Oh��f�9CBa`"A'H�dX�"O���`bA+�29�A�,$�ԣ�"O�0�TO�Ū�U��L�٫�&z�<����Y���c#&�Y�l�k4`F[�<�FJ־u��ĩ)|G�c�G�`�<9��"Q����o�Ba{�gH^�<���	0��%��ٜ��d���^�<c��3�bxSG�L�n��!BX�<!�*m� �]ɼ�����V�<IP�߶e��h��/���#��P�<1f-L�3Z$��J��#��D��C��>��s�*I�U�T�k��ξbG�C�)� H����%��K��s��c�"OZ�e�#}���T�N�eg���"O�9� d�7���J�U��"O��C��eR���ܱdT��"OVɊ6��3V�^�鄨F'+@`��"O�̪F��4����#Ȉ_�"OH�@1�U�3c����ɇaH�"O����dY�i!��زdB�-��"O��z7,��m:��O�v'`��"O&�1Cń�R��V ɿu�.��1"O�@��0��\RRj�g.="O�����q��AQ��Lge��`"Oh!� a���r��tY�}i "OZ���,�sr� gB�*�0�H�"Ob�2p J7�d<!��P�E�N�PE"O�pԟ�b��d�Z�2q"O�AR�/N����*X~�x 1f"O*Y�p�>|gd�i Qm��A�@"O�����S:0���$(�ޙ�B"O�Y��Â'���9g�(����d"Oz��wB��N�����������"O��P��3z��:sJ�0���Ȧ"Or�)�)�.J�g	�ڨ��2"O�<F L:X��k���Bwh1D"O|�� +O�5G��Ҧ¾Yx֩�p"O*�0bU�rB�DE�C����"O�x2����p%�u�(41"O�`�%�><��BF@F�N�c"OPeR�Kذ@c��a�N:M��V"O(��䩕�2����0�EKb"ON�{2M-~��1sS���`��"OT(�j?��p�v�R�?��o>D�0;Զ��Q��BV�gA����
��y��+]����C�o��h�#O8�y���L�� k��iE�%�ƃ�y��Q��J!��>[�ȥ2C�ث�yb�L�<(~q�'M��9*o)�y"�֚4�t��5gJ�@n�X��*�y�I�-S�R���a
�
�����y�̀<2��!���;qR\1H���y�"#�0H�ţn\̍�gm0�y2�������{iX�0���y�#�*cz�	�E�"P�Z���y"�Vi�Hm`��($�� 3�I��y�@F|S��`5h
ܰBÑ��y�(˒D��-0g�K��T��5fW��y��P����
�I�PӤ�ݪ�yr����n0�����̰:˰�yRA&,�&�ے��Y�><s����y2�A'|ص�@#L�$M9��9�y�ԟF��H3�Q7J�>��C";�y2�\'^YD���A�G�������yR*P(-�D]���P�8|Z\�A���y2Hخ�r�0���-:"�Y�FL��y�j�"��h�#�����&�yra��E��H��# �x�@)���y�N�a��(�TCP.w�#��ͫ�y�命&8*@�  6r�ڄ"�5�yB�F�j�U
��l�H/.�y"DNhJ![�i�7���r�G�7�yb�
]��7�fl���e�}�!�DU!'ZI��uV�l0��H,d�!�D�R���@��j�H�sRm̹�!�dX�.����(һ
����&��w�!�� �dU�S�D�d�@�b�ac ��"O><�o�3%Xt�GØ->1z�3""O4Y��Oh�	�������"O�]
���>͐��/���eX�"O �ۃ.đ)� -�ՠ]/`<YH�"O����:b�j4�7`�z�PtC�"O��quB�#>d�¨�5~�6�i�"Oљ�(�}}z-��	ۺC�VșW"O��p�s��z��	:�NdHb"Ot�vL_���  U�٢"O���`�ؕ��Cu'ѯ}P�=
f"O|؊��+QT<6f]�x 	�"OpaU��X�A2FO�o�Z�{"O��Kc�J��堖.ѕ �����"O����(Q�� ��\{~(�"OV-	��"x��}����N��S"Oҁ��	]�5� �V&��F��m+2"O�u�!�C��̣��&�lh��"OԌ�T��39\��C�&n�Dp"O�M�D��BY�cG�U]X0��"O�H�R��kp.�s�iF�WZI�6"Oz9Xtk
�P|��B;P���"O&<���C�Xu˒��7$8�L�@"O��he�ĨX0t�8�$�)E���E"O� p�ǐ{@H`�c^�Qؒ�"O$�*ΰ~�`�av���C��Z�"Oh2 A�Jk�T����s�6�{w"O��䜔\�X1+߼8�Z534"O�u&M�="HY�a @�}��(��"O�@{Cʉ3w}�XC�)RBhTH�"O@i!s���}���3[8��"O�q�� �,� �A��/w"܀�"O(=��$�?�VI��h�В"O&����2���"f��ð���"O��)C�V��jA1�fI�i�2��p"O��;6!�;��(��.����"O<Uђ���f�@j�'BN��
,D���dbR�L"�ъ���,s�z�X6!(D��2��.�2|��D�lTF�V�'D�8���0���PUH��$��$D�h�C�2�4k"�=8;F���=D��r� ��6��m`e�E89a�0��/D�L`�I$CP��3�Ώ���g�/D�Љ��w�,x��F�ca
��J;D��i��ʇd�&�Q��	u�\�"�8D����)ׯ7�جR�P�] �@B�7D�00s.�/�X<3f`Im,zJC�6D�|80�!��D K�8T�
�x��2D��9��"u�d�!5`�Bx���:D��� J��1z�(2e��\�0#&D�Dq�
�A�$�����a �*#D�(8D/žm�&�� ���.lYö!D������0�]�ÆO&6kH��p�;D�ȹ��Ӣlt��p�+Π6�<u�A�;T�lK�a��u���h�$��#輔��"O�]�i�t�� ҃�'�~�"O���#b'�=Z""�"�RIQ0"O =�UE��L�`*p@��(T�1F"Ob!R��$�d���X�p�K "O�dX�ؚ��d{2G3i����u"O	�C �1�Us�ȃ�z����"Ot�yU�R	(��-��ޥc<��"OĠi�k]K$��n� 4-Hiq�"O����x�F,Q$N�3���q"O� �,y��XUT���je��	8�"O�4��!7�.��3�c�T���"O04j6�[�#ȥ�6Gt���"O�d�iR�A���I��ך	�fY�S"OƱ�S�Q��閧D&B�l��"O�����͙x���'�)0��xBa"O0r��RT̈��g�
�<�"�Z�"OZI[��P�'b`d��N�L���!`"O��;S�5|�a�I62!�Hۀ"O<5�d�Kv��4`�oO�W3�LE"O��!�c��@���g��vJ�LC�"ON��6� z/-�D@��8CX�#w"O�e(��[�%���2p�uXƝ�U"O�X�th�0T � �TAÞyu,}�6"O�M�"�.vN�PcO
��½�"Ot�2@��<4إ� ��N!^�1s"O��*a/ܜz�`�-�#vRDS"O ��Tl�1X_H�Y�mX�MrP�;�"Ov�:wL�,��\c��ϲy@�Q�t"Oz@�C`	�N�\yʒ���Z9v�"O>���FD��MISa :_|�,G"O��k���D��U��,yf����"O*ɐ"�V�G`��ugI�E�r�@E"OPd�!`h���VvF���"O���C���~�F=��Dͫ/W���C"O���ʍ\	veH7Mv<�F"OL��&N˴&F���DK�C&�u*Q"Of}B��2b�pCA�<����"O��$��X�ȁ��.a���z�"O��)!����Zhs*U"l(X�!"Oui�l�Y�6�KQ&W�i��"O�0+�
��N�mzuE	�{��\J�"O&��#�*b��@1B̈W��,�%"O~��7Ɩ%���#A�/Z�YP�"O&E���S>��ZG�+jq���|��'az��B�U6P�3�2j�!���R��y���'B���N�LT��G��yB�Z5l\��vI�9sAP�a%���y��
*H��t��=ǂu��M��y2�M-:�Eۤ�����6���yr/KP	�lIeBѩ0�����y�U��Z��Lx��
 � ��'���?���hA�"�L�h0b�:d0�1Qg/D����,��6��쨕i܉b��PBG D��:��D�|�!�K�;Ð@j�a=D���ï6�!���#I� ��)D��X�bF�[������/��	s�e,D�h�0&9;j�ɝ�p��]�F+D����mD�l�t$я~W�8s�"*D�,Aq�% �C�¢;�ܤ���&D��'�\�Iv�pA1�D���H���'D�P3�ռz��g��A����$D��s#%ƛ6"�hT�C�\�J�iT� D�3��[�c����� ���d@=D����ԛ��
���:B���d>D� Sρ"4;�Y��0U0��<D�Lb�H����!�聽v74��:D���D��# ��"AXQT �2D�VD�4] �����/pXR(���.D� �"@�,��[p+�()b)��+D��ʠÖ*^��dEB4Z����a)D�蒓(ڳc���Ef�M�v��/2D�P���MH�^9���A�:i���%D�dA�-Y��܁b@_�]wB
��&D�� l�ZS%Q+�mB����m��"Od"h
�V|�$U�Z���r"O�${$$P� Y��]�a{ "OĀQ%5��:bb�8���%"O�ЀF��66~p�8�&�*��d�P"O�*
��QVn$����+̌�a"O.x6��;4:��s�9#�T�G"OPUP�Ǘ6p��)sa
.���AB"O��8�l�ͦ�;C�	(.��1""O�ɱ�n�5���ɔ@�9l�ࠓ"O�aI�A:@/z@����Z�x�"O�Eg�Z�,L(Av��5bN�"O��u��)�զ�Nq�5a!�|��'Z�	����9_&����0�t���'��	���Y)!�i��ʕ�|Yt���'���*P�(T�z�Z3��*s��p�'X����ɲ��ʒaAo�n�I	�';��`%IԀR�H���A�_�� ��'X�b�h�1p諦��Uf���'x��ࣔ�b��tss�ɱQ�h:
�'��m(��\A3|M� �[&G�Nu�ȓ))P9�%LM�!1�)�!`�"���Q
��h>��P��SB8���rTx�Q�a�����fF-
D�ȓ!D�v# %z ��j1��rd␄ȓo�l���)���� ��|�ȓ5�y ��}��b�wܼi��uQ<�,�*Q�3��V���4��wt#��5gf�p[EDV�,�2<��V�Duh5c>(�9�4Y7e��|��o�x)W��F�z�4ϑ=5�4�ȓ������>2vfX2���q6}��^Դ���X�rZ��!d��^���T���k��K=�A0�F�3�l��"���R���^���!�m]��@��L���*vH�\�ֱ�7·�0c,���VΪ��q��.K�:�A�낅x��m�8�QB͋"�,���I��u�ȓT�����?7��)��S�s�ԄȓN�x�`s�� ��D"@c�aNY�ȓO��%Sgc]@���h�T�eu̝��O�p����P�>qfR�H�ȓtE���v��7~��}�7�W�I�\,��^����ȠE!�		�Ƅ�����ȓHȶ�@�fD�6y�9�a$u8��ȓ=�k��0Z�<�4��2M����`%Q¥�x�T��2L��Y5:��ȓ
Fi� ۟=�(�"�(V����/�fh�aK-sl�@�`� �P��`�x�Ȗ�.wxA��`C�|�q��T Z�c-r���U�~f`e�ȓ6}���@gύV�*�ϗ�D͚�ʓv mh�T#�(�#��W�~��C�I�P�����)؂P�J)JǌU+��C�	(%�L�����2^!v|�N�4�C�I�v�����*j�>�Y�	�y*�C�		t�4�q�`Й,�J�* �h��C�5����	�t�3uL�/rB�I�?&8PqA��c�r�1Ɔ�e~FB�I:N>>XB�ҩ IB$�i�4k�C䉀H�l��R,A1f(��1���Q�C�IO��K���$kP س`C��B�I5l\4(DR_�e�6��j�fB��<S���d��E�L}b� _�f\*B�)� ���Q�<\��u��H�/&~���`"OX=j(�3`�1��]6{H���"O�	+2*�<�e��É*8B!��"OT]hQ�/V,�Ѐe -A=ʝ��"O��#��	9��٠�i�eל�Z#"O�b2枘@͞��4Ɍ�-�T��"O�qShT@,��H��b1��'��Sis$13���Hĥ�(�C�!�Š�d�����J���� �!���n�1 ���vD��*�&�.#�!�D]�3�,����9%�,��@Q��!��9�@8Rs�Œ��8{`��y�!��#X����+G�T�@�(�!�$ @�,���.@$��%<�!�)d��m�$	C��G5,�!��P#��i���6UQ`�r�%!�$P���u�E�?N�Y)$i�-h�!��j8�y�qe��@_Ȑ`�Ĥ*�!��*{z���"� �fũ!�ĕtz!��(� ����ƮI�%����Ho!�ā,2�X���j�(�����;^!�dȪ`Gpl8�/�0+b]!����!�$�Q��%�B`�$����9!��<F�B���茞)H����6!��/SU��CF�*UZ�Z�隮t�!���S?�8��*2�t�W��0�!�R�|�VQ���X�,, ��� �!�dQ�n0��D�N�r �5�=�!�D�&Os|�k��M�@��'��.2!�$�h���`v�Q�$)�Qh	�Q�!�$L�| Z� ��zΩ��"iz!�$T�HW�J�㍞*_�AZ�)�� W!�PC�e��E��XY΍���Z�L[!�S;d��� �M��;�焊?I!����z�(�6�G3�Уt�ΆK*!��<qs��	MP$�6���OT9"!��[3A�  ��"
��!U.I,^!�$��$s��Z�:�8���ĉ!�DW8(�@	y�&�(m����NC�!�L������%��%!.Cs�!�DG�;
Ba�gHO�훂�^!p�!�DPT��
�,/�Q2��6g!�D�-��	"GϬ}Ty1C
��\�!򄑈gnD	�iZ�d������6N�!�$F�M n����%ޠ�9BF�!�d� �,q�JՒ�,����"b!�$׻%N�r��_��a��+� tU!�$��S牵
�
����D�!�D�0O6F8����Xf�4�`�L�Y�!���H3j�T!@�'Wv+��Ψ:(!�D:%�\Ě�eT8xGd���`ȑ '!��+bD��ڕ��8	��kD�@�f*!�ܝ
�L��I�9�����(M�u!��x�v�qԨ�.F�쑀��qI!�$�_\����E:�vBĭ�'!C!��9Ir�2S`��Q���R�lߓ5:!򄍹���ʴ`�R̠%��K�>/!�$ �9�%B�M*�v�Z�$�7o!򄒙"���@���}�R�#��B�[7!����ԁ!(�/F�d��!��$!�/Yav��b�H~�Yqx��I��R�e�^�v�u+ݢ2a��ȓ)9� � ���2d ��l"�ȓ�ZH2��ǫd�ڌc�<$ ���S�? ��S��.�IB���F��"O�Ա��� �L�)Ê�Cav}z�"O��K��.N�B�vi�;`hxbF"O"�  �,�I�jޒ:Q��"O`H&�)C��YPu�KRD"A�u"OD�S�c	^�EA1�P�{1�¢"O��r���D�IX�aM7`̋�"O��K&CeKp�� ���)H5���"O$=�����M��q�2��M����"O�A�gmF��L����}頄�0"O걊W��A�.I0R�Ɲ�^��$"O�� u.��]|��FK�d��"O&�:��>�iJ�fڬ~�l��E"O��э�1^Ji �f���tQ�%"O�iؤ�C
qE�L(0�
���"Ov�+$F�QX�������LAH�"Ob�A�9P$�*�ó"nک��"OBcE���\��u���+[��t"O�����bEp\0��&�4��"OC��#�p�A���� �@˥"OT����T>��e� I$*��YQ�"OB�Csa�jt�o�Xʴ"O:���틣@��M����4�Ȩ7"O�H�Z*��c���)���+č�y��1��Yw $Ģi����yR	ގ?V�Q![�0B��se�4�y2�!��0��Ǘ)������y��W��T�1�T'
F$P�yBJ��UNd%�d�S+	��ua���ybo�8X����e@X4/0h��C���y2�ݯ^���F)�^(!p�@=�yB��g�T��Ā�%@�q���&�y�L�z���L�=5��$X2�!�y��|Ȝ|s ��vC����'��yR@*d�� w���~f���9�yBK��*pxIq���{�`ѪЂ�y"M˴^�qQ�K�x3f�c5�U��y2���`�̀z��<���]�1U���ȓ�U����xА�&,����D�� A��W:t��A#����B�	9![lК׆�J~���AUd�C䉎~��8`j̓om`9�g&эMB�<C��@璃�J��7PòC�6w�ZA�iN�v�J�r�$��,_@B�ɇp$�!��I��w^7mzB�	�t��-�ӃʜX��&�/i�|C�I�v�aKc��2S��0TȖ�7�xC�3�X�D6�(���YK,$C�	y@0���j
�?��������8��B�I�d��� cʄ,*�(���HC�C�xB�	X��Y֯-zF�=�ܥB�vB�I�7ihqh� �R)��kA�Z-o#.C�I�T���	S:��ZSN�C,�B��r쐱�,/bT���'WgC�P5(��.߹MJ�4O�&K��B�	M�D�PU.^!B���t�Ŕ  �B�I�y,�a�HRS�����:5�<B�	�R��s�ʒ&o��q#)@L��C�	�	$Z;u��zo��ӥ���2~C�Zpv�+��� �Vm:��P*XN<C�	�2�h!zG���^�<�CLE��C��B���@�\R�4��k"M��B� � h�E��Cg���'��R�RB�I(O�4��.�4����SI�;b�FB�)� �[�*�<w��EV�ic'"OV�p�e��L.xH�b�G	?ͫ"O2Hrq'ϋK%Ȉb �N�(��RF"O�M�P��x[FCjJ��>T"O,���$q#$ W˂�q�\�G"O(}xB��PK�����!�6�y�f��z����%*ڴ~��@�1Z5�y�A�w��D��)@-P��`"�y�5y2�M[�~�V�i蒸�y�[�B�~�`HLs��9Z�쀡�y"���7��3V��n �	Æ��y⋞.SX\��qG/<��Mr�Ο�y�7d6�=�S�J9ߖ�bV!W��y�i\������h�1x����_��y�*ŗ	)�Q��%�.�X�P��yB/Ԋq�> s��4���Ǘ�y"�ޣf�楰,��:"ƹ�Aky�y�g�"s�	�3*�9V4��%�D�y����|82�Z�/��T
����y����P� b䀽
��E+��y"�������(��謃�N]��yb)śO �W4	'|(h�̔��y��*R�:)���z�	`��9�y�'ƩQUV����ZzK�D
!!�yRI��r*�h���q�jx�����y��"��&�֮i[,8�Ī��yri�v��(����Z��!�y����h����͂ ?T@"����y"�ūh�@���f��Xք��̔�yh@�x(��9'�=~���tA
��y���bI��p;��@��W/�y�S��^�r�F^^&�d����y���+����IT�\a@�q�h�.�yr��{*69���VM`E�e��7�y�g
�nQt�W�7�n|!u�M��yb�R�Ps�tz��J /����씇�y�o��|':�3q';#b��h���)�y��]����Ώ� ���Sw��y�c�8�����3g-ů�y���8
,�4Q�l�
Zpusa�D��y"畯MG@)�Qe�}���pB�ybE	"AR��&�{;r(�����y��V��P�pf�Y���yB`F�B}�l��v�H�$�E��y�-��� �*սn�ڌAB�B�y2��\����I�gp1�C�$�yb.��l;T�'$�:\IfeY�`_.�yk�?G��J�(B�Z.�`��h���y2h�h�,Y��ܥ
�����yR埛"�N�t�ƽ.��u��b��yR#�7C���[P�W�%��;v�(�yF�+5�h�ᨃ��!i�2�y�I�n��t"�w��u��,�y�	��^@	��)G�q��a�S�yb�I�y9�� ! �p�8���EE�y���T ���|x(��sM�5�y�!�j=�[PJX�s���)d�:�y�k�">����f�w�"�( �y2d[P��an٣�2)�FJٵ�y�dY�LPBfG.�� �j��y�/�v�i�CF	�)n�XC���y���g�X-Е�R������.=�y��E9����ں�洰��?�yr�=y��Ur5+�����l��y
�  �W��6 ��	�rN
v��	"�"O(%I3�\�P�T-��L~��r$"ODDWk�bDb��W��2�X�2t"O�-zWԒ]}�i�2�S�c��x�S"O��+��1DУ�.xa��sc"Oց(�dY:\�J��rf@�X�"�@"Od��ǣ�NM!�+@�S��5B�"O�I'�͌ D�q���_w~,�E"Op�:���1�:��#�Q7���"O��9�+�5P���� �M��V=��"OԐ��Β�$���I���:"Op�k6��}�� � �/?���p�"O�q�Ԥi�x���I&H�X=�"O���#�aBHH��0y��;!"O�����D��vU�G]I����1"O�<���*��P�����Rhc�"O|\t+��Z�����iXrS"O�z�o_�-�h�CO�<���J�"OdhGσ�̠1	$�W5��hy
�'`@�E@��!A�d
��GQ�D��'��d��i��	˸܈g��qYR��'��$i&B���f̈ �4y�'�¡�Fc ��C�I�iW�p�'�0�+��D)u�Q�c�g�0�'�z<d.ûrt�����P�p��
�'�����iεP�4�ԀK,K뤼��'�\�b�nē_F��c*=�.���'�x��6��'(/�0a�-�'X���'�T�6 I�N�KZ�T`��'���1��rD����\�	�'d�2���<VS2,C!g��t�jhR�'��p84��JFu��S�|��@�'� ��D�U-���G@!���	�'u�HS��3�S�d���v�h�'��X�͏)>F�����o�u��'U�qJɖ�a1Í��$�K�'@��$�"IX���8��J�'�h����E��kp��y0�	�'��Hж�[��|JAG���]��'2���{��〨�1�v�'>6,���"kE��()R��0�'��}��V�5�h;���p��}[�'�'�V5ofhҦ�˹h�T���'_����̋v��pɎ_\�	�'�1�Ã)�J&��+\<�3�'�!�r/X^�]���
��\��'�H����ii��s��ź3E�x�')fQI� �,(G���scu�V�H�'2�8׃ǋq~	:�j�s�^P��'G��I*�rt#ê�~�I�ʓ<=�P��iʼ)��9)m��CV�ȓ>�
(�eD�X2�"g�zV�\��"4J$�p�T�� �����2���LIP�0EȲ.T$�nL�gh����;�J��
5.�$-�`�&t@�$���z���Aҷ:�����5�$L��_*��鷬I��� bȔ+J����"+:��iW�>�d�s�Z�x�0��E�#VF���� ���nL�`��d^T��.\k}�;͂��4�ȓ*���!oٚ!I~ J����m����ȓht��q�-Q ���o=M
4��� d�Up��W�@�`FH�?<�@��Ga�E�te��,�P$W
f��Ї�S�? �,�Q"��3S���J),&�(�"O�x@��ffRĢ G@(�"O\lz��iFU�U�Űj+B�z�"O*MX�+�+P�v�*_�`��e"O֐���B���
UF^�S� z�"O8�*��(or<1�%�[�	���Ӆ"O�5��G�w���`+�G��*�"O��0�O��J�k� K��	r"O �CM��W�.��1Ǟ���"O�es���$6�{���A7@x��"O��E�FD#��`"���7CJ�1�"O䰋��x_V6̢D.\Sb"OnX@B蓋�X�+ġ	 �D9�"O	���]�T�Dh�j���H!i�"O�����"5��#{1Y��[J�<1�Ъ<�ȸ�g��~\V�X0B��;>Y��*���)I�X}����hU@C�I6pY���o�W�v�W�b?C�	 �0�@o��s�����k��%C�ɆC�����E�b!hT� &N�B�I[R*����S@qj}�кA��B䉺0�������W�X��#�B��B�	%e2��C��
:!@���#>^�B�5��d#V���#�����,��"��B�	�rs^��h	�#�ڐҠ�T�B�I*R,d8y�.ލ#}����@ޖ��B�ɯ:�x��Gˮeڠ���/	|J>B�I".w�4y�L(9��<����>�B�Ɇ7O4���i4A:���ARf�B�	BK�����"F$8�e
��C�I(Q�􀓃
�W�m�eN�nC䉪t@�����D�#bBܫ�˃�=�4C�	
>b��icљviHp� g�:S�B�I$ڽ㡣�G���¡G&�C�	��=��;YM�d�4�?h��C�I�>08����Q��S!(f.B�/�~�c'��{�H�G��=�2B�	(q����í؟|���b���wB�ɢ
P��s� ȗSQ�YY�&(C�	+�A�7�T�F<��C��κ0d�B�,]wz�@a
�;�F%�a�O3L[�C�	�d�r�����X0�Q���q�C�I!e�pR�B.ql\���Cu7�C�	J<�9h �B|F�
���HB��)f$�p�HF!
�{��,+�:B�ɝFF��`\�AVʸi�jG
mrB�II�f}b�	v��KuL�:Z0C��\��Ӣ�=7/� �%�[�t!`C�I���-��F�N�@���(vGB�I7|�X� �)��H"A+S�Qt�C�	(�b%���?A��sżw	�B�	�\ :�����msPY&	�~C�ɱ&�|�З��3�6e�u@�9hC�I�w|�Q�t	ǈT�)[viȫ
�B�	�(tZ���O� �Ubv ¤תC䉦|�>ar��ۊ#c�h��R�p��C�%w�*J@ԏ��O6��F�^�<��Ȁw�0����7/�Y���W�<Q�H�J���IP��.��`/�P�<a�)V
+�b��0��V�@A�ϋe�<�sGFh�\�#���NU�l�'�I�<���K����`�A�Hd���,I�<qj\D�r�ĉ�c���MWM�<It�W�!��8�\;m��G+_^�<� �A��H�Z����B�"O6�@���*��EL�&
���S�"O�@�Sf�,Ha摡q���(�W"O �k3�N�OB���8pc�| �"Oje���B�80R藫>�vp�G*Ole���ݰ$.	��E�Eo�C�'���#*� @\u �eی���
�'+�T����I�f�Bt��m�q
�'~@�Y#�90�b��3��|�ΐ�	�'Yf$��,S����ͦs�V���'��5ڵ9Y��(L*gw���'ᨉj�S?Ģ�����1x�uB�'X��� J	<r���'D� zA�
�'R��+ĺǬ��'�Ȇw�
��
�'�����N��Cj�1O��g��Ԣ�'oV�bu�M�X�,�P���T@!��'e$��S�����H̯K8���'Ǧ@㑃��r6by���	!s�j���'�E��B��|�Y����c
��'&(ق4@Ͷh������BHF=�y�N/dX��Ǆ�3j�p��N�*�y��;{��'ًrȸ���4�y��P7.����/N;5��Lx$O���yrMW�A�.����#���EE(�y�ѰIh2T��cͨ"�*�	6���yR�Y���s�T=��(sUM��yblX0�|���jˏ��E
UD��y2�ֶY��:?�D��H��yBoG<E����`Q��c`��y�j����nO6+*��#M�G�C�c]�M��F�%[+q��7��B�	�Y�((!�E���Xs�מ
|C�I+h�<����sk�p#���W
C�ɠ	tu���A4jH��P�D�3t^�B�(sv�#a�Hу�pC䉷I!v5g�ֈ:<;�o��wDC��+EN�ɵ`��&D4��Dψd8�C�	�]ۆy��2$��������C䉯k�T�5�� ��\���F$բC�ɇ���jP�VJV��Qx�RC��S� �qo�5	~t@���7zJ�C�I�/~b����;�k�';�zC�I,Cd(��$&^4y���Ç�.�VC�Ɉ7��X�b�9+�M``σ+_L<C�I=]����F‧3T0���dy3C�	�\��@ҥƂ�BM.	�����'Xn �GK^4CGȸ0�ʝ�|�x���'���8f/����)`3hU�y�J���'TRA�Y��(i���?o�5!�'�x;��Lr��,hԁ��L	�'����GބO�2�J���B^<�'�sЮ
�;�d3f�y���'��\���{$*=�GJ�"Zպ	�'�2PztB�*eR�j�ܞo���	�'��2��]�a��P��F�_y��[	�' ����&�g��hJ�כVkB���'��3���P٪��5o�.X�� �',zu!p�\�r�PQ6^~k��	�'`��'���Y�v��z|�)��'�DP%��4j���աD�_G�(�'�R�9w�ƥrмU �Mͫ
�����'��r�/�=kS���'�/W�b
�'�����
	X�,���[�nٳ	�'s��T̙$f��suO�"U������ �(IV���񐐬К ���"O�l���ti �R>��{�"O&!�7̔��<�ۧ+̚Cd΄�q"O��h�	��e��Q�6	+�[�"ORU��)��N�H\cňG>kB���"O����ߑi
���&�4>)F5Q�"O{���WbyHŗ"lʑ"O�,��M3Y�+�4l��$W�<	F�ULaH$qI�8-�X���U�<�FX5w�.t�ŏ�G��!��X�<Y����f���I���=g�b��K�<a�k��K�|�J'e������ks�<���H�#���B#���@ Su �k�<I�+ثZP�-j��̪om�Y��KA�<ib��	���F�ךOt9xaO�}�<Q�Ȟ:�\{�Sh=�	}�<�T�Ӫ���w�
z$( rN�v�<Iv�Л!�p����-I��^[�<0�1j�T@�KR�e�n1dAX�<�A�K0m���ϑ&w���!�T�<�w�B	n!l;��45��|��@CW�<�Ej0n�>�r��4K�Vب%��S�<���Z�q����M�~�f��&�h�<�䌆gY:l��V��behGb�<1�*9Y��e�4'�A[�<�`m�S�<a�a@-r	��D $j�4ɉ��M�<a"�d�D�a΂�k�`��)~�<�`�P��1���U \�����E�x�<7)
I���ȴ�˺~~��b�)r�<�jY�B�]
��!�aȗ�C� ��sE!@�X������c\�C�I�Èy�¬�����v��<4�C�	?"���Z��0oD.Y���)��C䉪X�\H�	�
!��J��} rC�I�����s ;9B���aS7G�DC�I(E$��Gk�v�J�(�Q�JC�IW(d4��U(o��B�M�qy�C�ɭ/cL�����6�ҜFn��R�C�ɹ:<�f.d�|����]�$J�C�*�5���]�PA:V��%"O^����Wn&��bQ��}��"Oz5k!��1�����f�P"O2�#���*ښ�Qqe��k�n��"O~��@d��P��$B7���6��@"O���#�Ŧ9�O�@k�Q5/.D�l�7!��<ޮ�{�BB67$ EP0� D��s��
 �0A�c�+9��JE�:D�� ŕ(�q(�{��l��9D��*d��8/��+F'ʠi��f(8D��jĩ9F��#��F�K��;�N5D�|���+�xl��K��/4��y�5D�t��)/�x ���b�y�1D��2g�ШV<J��t��91��Ӕd0D�`�b�ej#�������k(D��ȳ��1��!26�A!����(D���錾6Wy����1�T�1c:D���F�]ܼhT�*s�\�{��=D����˺w�FlH� �Z�Xؙ#�<D����Ǵ$��@�Qn�)��=���:D�P;����A�EV�� �`7D�t֢\#M��c���p},L���5D�\Rq�:QO,�J�"���2A��4D���\�����rnju�'&D����h�:\:h)b���dI��"D�� pH��B_r��@CFԏ33x�S�"O�0KI�(j=�(!��S3 R�k�"O��J��Ĵ:KL����Q�h[q"O�dq��
�Fՠ��IظY"O�h�T�P%Xp�(P6,�[@tA�"ON��!�(s���$|>P��"O�ui��ë�Jdb�)�.,���Q"O.������qi�)b�e?���R"O��u��#`{Y
�$N-|K���"O,�X&� (I�]u��>��L��"O�홄�˼�,��G��G>B���"O|�(��]?N��x�׆©d8zHI`"O�1*�L�+I�:��A�U%�u�u"O��(s���X�N9)�Ơ)�����"O�u�eNӮG�XE`v&�J�T�bU"O�\�b	�(0�կZ�	�5"OJ��DM\1'L�qČ�ج�7"O�Y���Px�y�#O�;[��S�"OXdQ�_�T�J!8�b4H���"O�0����{�||	�l9vCح	�"O&��'�ߏu�J,0#�	�L��"OJp�q�~B쓑�շd���"O��FlL0?�T��1�06� "T"O��z4ȅ�#��̣HԆ�>���yB��e�,c�F��5�X��"	���yB� �Q��9��$y�t�������yW�T<�TS��pв=�7,Ч�y��ƺ+yj�#/��l���רG0�y"��5W����ŇlN"�N(�y�`�68p�񋀨��k#~�����#�ya�,���*��R+آd&# �y­��B ��j������yb+Ǐ&�V�c�-P�o,�d�ː�y"�D�Z��0�DJ�%}����ɠ�yb�QMV�a�9m�)q����yb"_�KX�����`�f� �](�y�MR8�FACGE�$�59"��(�y�ςlRёU��4&����^�y�R/#ʆtr#�N.eT��-ܽ�ybF ��0	�o�F�sp@��y�H��^n,�è�d�X���C��y���7rKڄ��݆ho�����y"ˀ�v5�|`c*9tg|`H�E��yĚB�(+��� �L ���� �yrE�7C���4�ӰMcF������y�J�C/pmZ�'C"]�j ygAF/�yr��<���8`�6d�N Kp����y���</����1͍�q�����΄�yr/
7��C!�A�oD����к�y�EA!T�j���BVa
�42B���yb�V)'�.��i�	�D(�y�)P�L|�9 �ٴxtx��+�y�ᆦ]�:��� XҠ{�.�	�y��&?fq�Ë�&y���y�f��yb�;}�LY�!m��x�4k�hU�yrN(}�P�ɰ��v$<D���:�y������ۗs{��i�Ԟ�yI�*[�	q��hJ}T��y윜
�h��g���cƔ��� ��y�od@��K϶	0\p�%��y�Ǘ1FI�5�r���QK'-��yr�I�0�9�� -�|�(��U3�yr.^������hӟ#uZ�ժǙ�y�
���\�b[��<��Y#�y
� �Q�����8���i��]w"O��t�C60�d���j[;CZr�"O
i�F�9� ��)�&F8�H��"O�� �Q�t�z��Ҧ�,�(]ڐ"O&옒�E
�7H�j�"Ojܲ�X2�ѣ�̖bta��"O��ҋ�6Y�N�R#�,F��"OҨ���&� �r�
1L��CW"O��֩H< ����&1 �c"O�i��A%;�lq�C�ģd��E"O��bD��2'�F��o��0�"O��aV�F��|m�g��O��6�"D�@(��F8Z�|HB���|��b,D��1�(�5H�<\R�V�
FDƈ,D��{6��8Ac��G;T�D�5�-D�0�$h��`W&�VB�=y3�m;r*-D� ���D- "Y�'�Y�gU���l,D��o:b�hA$�`�pi5�-D�HB3��pdݺ�#C���d�5),D�H3� ��
� ��$��+�\䳲�-D�|�0K�o�- ��_�58$��)D�T1ㆅ�b�Ӈ���wv�� ��'D�8�Fb�e*p��#C�� ctf!D��P�A�:����%K�2���[Q�*D�d��]�.((h����\\����'D�D�1�V�&T��p�8sj.�B��?D�D8���bh�r̎�-W,�AGk0D�P�alH2?�X6ΊxU�I���2D�0�p�)v���G*`�ɨrb2D�<��a�%<Ŷ�)�#�,%��A��0D����-�+b��	��$]�=r�	+D����N4P��0�
�#.TU��'(D���4/�%>R܅#�(��z&8��;D�c���cO��R�撪~i��k��4D�X�hI�,f��{W�ω[˺�I4D�� a���P���l�$`bX�`��0D����ƙ0Y�|�d�[�)Tq�'�/D���3�P���8F�ם2�p �d0D��p�͜�d��� U5 ��9%�.D�0$�C�~�D1q�,�4�,D��h��R&OCxa���_ �X�!*D��h"G��'ᔐc`���p�����$D���`�xV�p���1@�
�[��$D���Ag�=�=ˤ��zO���!D� 	3-T���i7§!��#+!D�T���Q����G`ߔZ�,�v�>D�P��l\�X��I#���V2�"=D��Qʄ3,5����f� �-s!�I.FLt��/+D��iVfBEn!���"l�1�`F�"0DXi"��A�!�[X�q���yͨ�8���&J�!�Ė��Xa�.](m�J���̑�k!򄛏f�x�_r�PM@�N�^!�d�:|;�/�?����c��	[!�d�ycF��@��<5���QE�3?!����IL ��E�1|b,�bKj�!�$Wɒ�L�T����A9r$r�'��)C�H�=>��܃`e��0_����'��L��D�e"�A���!s#Z1�޴�~2'��0>!c��2�v9A&�;X=����Vn�<�3�,+�(ě���8l@h+F�<�����4X,�#�C�IfL@Q/%D�dH���_�l�2�U?� ��#D�P`���7{2�uS����3��x'��(OR�}�S�? �-��o��,�(�H�E.�( �'Lў$���6R,8�$l�4ZRX��%gӞ��&%�O�-; +��O�XP3��3�A4����'�đ~��fN�R�&��SZ���.k�<	��N�S��{P��&	�("�M�^?��4�?�y���
4Rf�����(;��dkt!�d�T�(1[�(j�ѱ�P�da���'T�~R��)A�N1+�*P�*��Iz3�X��0?i�4�y�E��{�ƙ��爊L. �����yB&�]�<ѱ�@�7��4�$���'Q�M�'���dL��EyH`��"ҋ~Lء�撰�y�HK�-$��s�Gqu><�%�N/��D;�S�O#�Ԛ�� '�z��C<�2�'��!V�s@"����=����'HV���W**�!%V��@|��'�05Jb��;@:��!��#���y��H��]�f�L7��Pb����y��)�<t�'杔[���!�HO���$��J�rsώ%�@t�Ç0n=!�D�]e�<�5G��o���څX�����#�O�z�n�0�r��3i��Gu�I�e^� G{��̼$R����F�"�(U�vE��L,!��=����v&��pt�W/��:�1O��=�|E܎/��p
PF�`
�ЃQ�t�<a$O94���96��+g�ꑓ1.�D��a�xbq �4+ԑpyp�p7'<{��Ia���O����`h
����,�	p*[��y@a�ra�Q ̐v(4-:�P
��S���O3�̀����Y'��?+Pv�X�'��+��ί��$[���'){���ڴ�hO?7�ۅ"/ƬJ6��P�Q��)�6>@!�ݏ2>Ȥ�G�6�dݠ��?!��X�#Cfఓ-�(��|� �ۂ a{��d[4nr������L`isp&Y�e�!�$S�$1�o�� �L�RGc�L������O�r��T?���_""JZ�iF�X� [a{"S����-�&� 4�B�u�$��#�ڇJ����M��i��m2)Ab��_�=�����R8�%�E)���!��΋kaB0�ȓt ���f@+޴�e"L
!��%�hD{���l+�r��e��(�2(q��T��y��A��F+�8or�b�EZ(�y�i�� _*�1�ߑ+�Dp�a�!�0=	�B���,��t)���:�Dۑ��8�y�X��� ��ӡ?İ�)1�]��y�$�(�8u�D��D~d�0 ��y���o�!`��_'�EI7�H���*�S�O�ҼQ�(�8%y�dKC���qb<a�'�h ���ՂG�X�%�9}B<š/O.��þ	?��W��v]��26���a2�O�� '�Y0`�4�9���,A�0���i3��{؞�[D.1iN	�PiH�O�<:�%0D��p�K��8q���R�5D���q又�(OТ}�����$\��I��"b��Ez�_��Ez�ȅ�S&H�<9�9�r�L�`��<��I��|�`ދ\}LT{�d֬#:��ȓs�ּh��H�&�4�@��,3��,���M��0qS�����.L � ��NR�<���=���HSK�/�P�F��t��h�'���+Ŭ��P�H��$OɻY/�`r�'A�P�D�]a�PAI�1 �ݠ�'�x�2�g5�^��B[������<��T��[�b]#2k�AVL�Y�̉�O9D���̝=-ht����P�
����6D�� f��W���q>d��$Ҭ_�]��xr�)��J���!,�x2v�	Pn�fC䉇=jyI�����-;���0A� C䉤\���B���
n��q�c�ǷJ#��?y�'W��'���yZwD
D�e�5�~ZC�ф�T���O�����A@ݑ`a�
��I��;�!�d�Z���·��N�$5��BB�s�azR�i�^�O�4���"Gzt��"�(d'"�`U"O
-,ILhT��īC6��ȧB���O*(Ezʟ�`�J��e�:���g׏@���0T"O0��b�86���I�/Ҽ��"O�Ubw�����|q�
� P�N�;E�����ia2e�MjDI�`U�<����$)?�$a-}2�S�e��� "�	?��k7 G�e,B䉘8�0%:T�Ⱥ��'Ʌ5B�Ip�����	\��`+DF��C䉩F`��d,Ϸ=P��fL5��C�I,:,"�A�L�L�R��A˅/C	�C�	$AALA:B!!l^�0 �ߏ~��C䉞T�� �Wd�9� �S�m_|֘C�	(�HM��F�5x��!.�)8p�C��,��ce�+]w2���ڪ@��"=��T?H�]G��4�Ï>�8C��)�	h���ӷN�м��LB2!��U� �NB�	�5�xaA�!�;0��L��l�#vKB��1��F�t�	at i�`H#ph�"�U�m���p?)��Qx-�dq�I��f��=�t���ݚ
�'_D! 5-[^\,�G��BƤh8�'pHe�DoBj�082��uT�C�4��R����yb#�O$lE�a��-�1�(ϭ�y�#߼g�Z��u�ij����B��y���7z�`�/qp a��@��<��{B�'��X ���TpS�ǃ'n�lS�'M�8��ݝm��ዥ�T�"���S���+O�	k*��X�x�/� 2�Ի#"O����ˡZ��9���_?a`a�v�iȲ#?��6�ɦLv���6�:s����! %�>���<�	H%n0i֥�%"Xv����]b��B�	0S^n�(Jŝw(�$:��].�b�<E{�Of�D��g@���ܵ99�$�T�]�A9�'4a|�$��BѲS��[�)�F�>/����(�TA�΁&:F����@< B�I�%8 Q2�f����2O
�S����O��([&h�(e�4I���3kuhX��<D���7�^$F\��Z �̶<fF�+'�-D���gB�L���S�k��VR�	��,�ަ�Gz��>�4�]�9��,�3�Ѹ<�P{���_�<ɐ��''bx��Պ_�W�j��Qr�<QS��URZ��+)|+^|+���o�<1���Gn� Xt�ơDab����o�'�Q?��Pe]\�(j��(g�i�Ck(�	�xXQ�����1��>I@����ݑY�>`P1�is��D�:K�p��SD�&����NS�Y�!�9H=ސJ�)=*�1�N5}!�4������#t-��� `!򄐧.�* ��#��M! @�(X�md!�d:f�\���?1����5S!���kM~��RO�&pGP�@��
A!�]u9&���A 7�Y��e2%R!�$W�<�<dXe��q���)+�;!�ԥ��`D.�,p��9Fi¾!�í��]A�.��.��|xe��2!��3*�l�q�/C%d�XjqA)S)!�=�8e���iJ6���	!�� .���� �c3���7Z���`"O��K��V�*|`���]�}�좤"O��A�h��'���dO�O=�"Ot�G�U48�ؑ��I�$>�8�"O�9b��� q�|�Fi�#��=�"O:H&+
�v�����@?*v��"Obu��ǍN�.��E�U,vs���"OdP{�b/���S5k\3"O�D٢,�*GO|Irp�b�26"O�pH��|.��%&)s��qzb"O�5��
N|����'d�y�X�� "O@-�'I�OC����6w�-��"O(�ÖL'H�̺$"��J���S�"O��cu�E�+N�����T4i��7"OlL񆂂?���#_#NС�"O�}��0���5�ӜV�.B�"O����l�L,\���þ̊|�"O� @�dr�����#j�8,�y��}��ծ�&�I��y��E<j`��o�#���rT�6�y� ���
H�y&�fCJ��yR)����Q�"�r�iZA��y�6��k�"^*{V, [ug��ybJݾzu�ZA���B��WJ�,�y¨�%P��ciC+k�xxG'�=�y���W���GnM�Q��5EKL��y���: zś�k�6�X����y�B�?n�� ����B2$8�	��O�|���Xn�T�s��O�7�d<��"O�&��Q̜��Gi�b�5�d"O�!�(��oV�4��O*!�~��"O �S$]�l�ڵ�¨��
�ڼ�`"O6 ZC�
H�b��4��1s&��a"O���Tɏ�Z�����M����B"OZ��3,P�m�P0���s�I{�"O�U�@���I�����U���#"O:UeM�,�-:O�U[D"O>��׼e�8@�1k��.�����"O�����ɅZG�m��7��%��"O�K#"�I�b����9�H���"OD�s���kv��N�<YH��V"OV{4!�$P�h:���9_��ۀ"O�͚�d��q�4m,9�=�"O���"�"l�� i�?v	#�"O$)�2�H�0k
 �E�0y.(��"O�D`�}��,��-�
b�"O�����e���,�@�9�A"O�\{��Ų9���{�j	8=}.�sC"O�p�҄Ը#IX� ��Ð�Z|aO�ds�M��L>\ɥʕ�u���A�6��}�פC�]�X]Rۓ�r��"c���Q�,ŷBS~���Ɍt8Գv)H2�A�B���,Hs.ڇ�P����X���2"Ođ9�n��$
��!T�
8&`)М���s(�rI � ٹ0"�9��[�'a3�U�ucQ�SC&\P���Ćp�ȓ^�L�; $�3�L�3h��$�J�%�: E�%�pH48�~<x�I@�49��'5nm{�
�;�P&π�H�=S��Ė���]�K>AccV7y�)	���2	yR�Jd`����T��p0-��#�FX�tF&,O���ꑦBmԩ�#mS�B�XX��'�a2�&]�?�2Q�'P\-�$��80v�I���	nIf�c%�)�0x�
Di�q�tm�
kR��
O�E3dE�%?��ء�ө=�$$�[��z��H��� $�.|�u�鎨,~��$��Kf��`v,EPp�Tp��)���><�j����"G��h����I4��Q�)ȼ_.������KOnY�Éc����U��=
V��DDS0��Y����y�B,}bK��*��(Q�
%eV�xs�Cؑ�(O�����.��!1�%dT�|�S?�����'�lm�Q�ǧ�N��!�JGV�Hz1NW�XfH�Aj��u�8`�H2�����N�=��D"r��skX$�c<�|�coO�!R2���Һ�#C�>������I�Ks֙	Ad�?6� ��SM��mDDqS��%j�����Px��إI�d���BX@Ǽ�wBσq|�I�$/V;=$�M�K%�xw��&L�p��C��E˪$����y'B�h��� �:4�����K��0>qP<U�y{q�ܶ%^�b���6� !`�'�85e�m�u�~m�rF����\X7�M<j+^�Re�V�-ntR�ʏE�dī%� �*A"ᐐ$��0b����ۊRG�	R� T�B�qC�\ݺ/o����,Y�]�����0r �H�rL�Čً��ިh�.!cw���.�ay�o�� ��Ӓ�TRTY���R�[�p�0�*ܲ+DT�p5���k!:���BG�V:^!�m�
HF`��B4Y@�;�-bu$�q��>�XI��'&�=ʣ�B�?6��4��m2�Dڡ�">�*����H�,�Ж���!�)��+±=?��Sh>�t�a������EY�g���G�0�BQ�5��>_az�MX�i�8��qގ+����`�����D�`W�<H6��4�P��@�jL�y&�g��1� `�O���D:}���g����)^��٦됵�Q�P�P�F�c���QtO��]����˰~Z%X�p��dM��DV8�HEJ��a �0 �ɁI�(�s$C�V��l�'"Q��nѕ��'"O~h"�f�)���U�
3��#�G& n�%�"�J�\��i�*�{��?��aP�x�蔀�F1c�d���E�X�6�10s�<D(����'�Z$�!��!l���hVG*�0ѱPN�6�:� �`b��8��!m���@�'��T �"��m��� �6b����i���&� �|i��I����� U�yjv�O�0�:�豊**T�CAY�d������Ω�ұi�&8���ui�]����8TW:�b��ЂrhA&:֘��6�׈�G}I�-)�`�'�B��Gd0JV`e��Q��0��B�i����n��	�!Ƀn+�Y��/P���m�)�'
}�:q,K�3ӎF�w�.�Gy"�8x���
�|��C��}p,(�G�߬&b�ǄX2J9�u��z��*��P�vA���O�ÅJ��5 Pʄh�8���K��1X���p [�@H���O�<���K�6Q�%'�U*��P0�
�
�nF8B��CE��U��}"@؟+��%��ĩGXt�`S�=6����I�Y�Z�:4%�
2b��c �(����OD�GZn�8&<�y��՜z�T�Ќ�)[	��G��0>�B舩x4F8�b*�I�����!�<i�Ų�O	'68�Q�4)�J^u�3f�l��X:ã��M��Ͳ�A�&=j�ͪ�/ɧ7:�U���%�.�v8<=
%[�� "��GxB��bC$q�L�upt R��ӀF#f�1椓�u��lh,\m�@�s%E::=:��N�V����6�D�UUt��s��	��`x%�I�F��U�ĤӨ\��P`�M�n"hqT�]7J@ �����EU�D�Fb�E��M˴DS)^��@Hd� �F"�E��-��`�D�@6�L
z��*r�ǰlh�! $�O�%9���!BMy��L�Xnʭ�PW!J\@ٴ(�p��̺u�����
&B��"����ʴc!��Rd#RA�4&�t�X�X��3�-u��x��_�o �xa����������L�8嫒6Z���ٖ��L�H$+�K�U�*a��*ٞkQ��L3�F� e�4_����6��H�F���.�<0	�
�W-��7��A@˓l�Z�`�+(�Au�J%
F���6I�4�֥j�I��TԬL� J2c =��!@���#ӳ$ʰ��&S1u���S���=41[�,+�D��a�B��&d| (k�[�8���h$�]$.?EV'�3�M�G߸���%�K��6͔<k	����<p��S�,�)5?�P&l" �-��u��|�L���-˵�����DX�"ֱm����$5[�
��L/f��DPx��P*��` ��2h���#��4_����c��P�4$���H�KŌXZ�'I�Q�I	�JK�Q�ռR������5V4�Eڀ�X�\���#qe�9�*�
Ճ�&_�I����Z\�k��C�T7�Y� �6Z���{I>�d遐3p^�Q#��%�l������<1#g��F9 ���*J
��˴I�6zN�y$��!�x��d��?L�$Y���7xk|�����X���q�R� �a�'��2�5M����<�Dɇv\V��,�0(��t��ɔJ�l�0w�T�J�x�2�4?�JE��醌rVB��l�/��p���ԔM�t���L"{VT�1�/�2�@(C��M���$r�"�	EG`t���P�8������  �E�eŋl���3�]�6 o�^�V��V�:���	���"��a��
o����\63L�Gm�f��	��@j�ik �A�|�qO�9�� ül:��m��(V�03�A��/�/�|!c����|�A��^�J�`��P��D�~I;�mG;�a���F.�x)sL״�r�a�c~���T-
>S7Z-����By~e��	b��+%C� gbeC$�V�Z�4�Ä��<V>N�P��4@|tqoZ{��a��,�f8�\�#� 
��SB`�<ʛּ�A�3� ��kB�\=�(Hx��$:G�����?$ ����w��Y�e.[����вOA0�*']�\��+̞3� %��t��q�N�_���AC.�0Hm`�j%�:�$���VC�uQ熉/ ���σN�DAd�wh��ҁ��	�4�L>١��
�&<hE��>bv�C�2 �RdB�']<m��&;�M�!@@R�d�PK&.y��W�Ρ:`ht�ɆB�L���&gE�A�3�6���!3I@TA:��[?1ܓOPM�[;9�1YC*Q�88��'e�T|H�g�̴�)2�G�8¦ �$�Ąql�y��J&yvp�C�ʢJ�DX0`�����r'�%<˴��d�#áR0u�T���1tI�L�����+�&
�]H��{r�������I8g�`�U�ٻ J6��`�y�<I�U䟇!�p���G�+$E�4J�F�[N�i ���>nq���D�5g l�%D_� �r��[�&%Q4L,��F���a��-e�$)2$�zQ$���M��v���$N���Ńy�����[�f�0R�	{\8�����*kd�H�@`!����P�� b����F�(��6�0�{�$�Z���2(��݂��0���SMA�X�Y�`����Lc,up����5ˈu���/m�-�t�S�ݔ<�z��1.C��tF�/8x�#�Ɖ�88 �£����tL�8Zd���k�����%3��I�Ʋ_F0���i�),S��K�4�f��$C>j������0��nM��j=���[&i���
�X+QY����n߮c.aaw]�`���;|�4����4:���Iꕔ)�2����LU�u�sk]�U2D��*A�R���G�3c��_� �����v��ad�ڰP4T��j�+	U8��g[B�U���C��Q�L�hl�_tPD�G�+�A��W�F�df�Ux]F�H�"�N��Y�D�ok�_rWB�E�%�N�洤��E�I4w��#�wE>W����F�N<}��,�{O6_������ F�N<}��,�{O6^������Z���d�R����9N�X�,��U���l�\����:L�W�$��X���k�[����6G�U�,�P�����-qM&�t>&W��2GEOAڀ��*wH"�v?&W��2GEOAڀ��)sN%�~7._��6BCGHЋ�� |�<�K������㬶2����4�A������孲>����>�I�������8����7�B��iֈ����%'�|�j?�`Li��i։���-.�v�c7�eIn��bۅ����(,�t�b5�mAd��d��]�M-�s����Ѹ��	�S�O!�|����ض���U�H)�v���	�ܵ���U�`����
�|9��G�㳭�h���� �r7��@�翯�l�����q0��J�	迯�j��թQ	��`e��	g@ȝ	�vO��X��gm��oH���rL��X��gm��oH���qI��R
�<��A��&�P�l��WOW�9��A��.�S�j��]
ET�9��C��)�Q�`�� PHU�6��N��5�S�N`Hq���'kE���v��7�S�N`Hq���'kE���v��2�[�BmG|��� nC���}��=�-�:���Z�p��}+B=~&�9���[�s��w&@=s-�:���W�y��q H4x!�0�~�86�6�@�>i���(R~�86�3�H�3b���-Wy�1<�?�J�;n���"Yr�4=���G��0k~�G�����H���L��4gq�M�����O���A��<`t�O�����O���A�]U��2�v�j�����XQ��:����j�����VX��?�|���j��� ��XPd�<1u���pj3���7���a�99���}`;���5���a�99���}`;���4���f�0��f��b��.8��.IB姭�j��m��'2�� IMﯦ�c��`��-8��#CH訡�jư7g��W���l��Mo�#���<�7g��W���l��Mo�#���<�5d��P���d��Kk�!���9�2b���Ҟ^�`���}��u
 ��>���ܗP�n���s��{+��<���ݓU�`���v��x-��6���ך������,�q�3+@�5������
�(�w�4,F�1�����/�r�1(E�=������T1�7+�@��"�~ L�)�Y0�5(�C��,�w&I�+�^9�?"�K��(�v&I�+�^9�)��r|�c�}>�ٰ����("P*��s|�b�<�ٱ��/#Q.��xv�i�t6�޴����'.\.��p�����,8��v�Utc׌�qZ�����$0��~�RrgԎ�qZ�����$0��~�RrgԎ�q[�����"�t�������@����[5�$�t�������H����S=�.�w�������J����\0�%�q�^��*��5����eD�q��^��*��5����eD�q��_��)��	0šz��fG�p��^�.���2է��x�Q(,�P+���5Ц��u�S(.�]$���7ԡ��s�Z"%�V.���(Ww�<�-|�b�3h6��y�d(Ww�<�.x�g�5o1���`+Vw�<�-|�b�2j2��q�n%Zz�w�B�:N	p�9�l���ɄcS�p�H�4Cp�?�l���̃kY�}�E�>Ku�<�o���̃kY�}�Ew�(�6j"�$jm����C��.�2i#�&ii����N��"�:g/�.nl����H�u�*�������C����=Fy}:�=➒����L��
�8C|x?�>�������L��
�8C|x?�=䚔��!��9]�<k���ua�9{�*��8_�5e���}f�:y�*��	0U�?`���xl�3s�.��p̯���)�͞����
tή���)�͞����	w
ȩ��"�Ė�����t�\8G�И»A�$υ�����_9G�՟ʱL�.ā�����U0@�ݗ¶K�(�������\8G�������m��Wdz��	�������d��[hv���
������m��Ta}����/��d|��R��9z"z��/��nyt��X��?}"}��&��f~|��R��8x&��&��o�ö�Bѻ&ڏW�SЈ�d�˱�Fһ"߈_�Xރ�
f�Ⱥ�Hز$ۋ]�X݆�o���T74��t���6eFF��ƽS0<��|���<iML����R0<��|���<iLN��ſX;���\��{}_��>@�{����W��vrR��=B�{����P��~{_�	�6I�q�����4�p�����|�S��h��q�> �u�����|�S��h��s�:�r�����q�X��o��r�> ��|

{:��Y�����f�v�|

x>��Q��ʦ�d�}�ww3	��V��ʠ�b�t�|
�:,����ǜBGL��Z�;.����ϕHL@��S�?(����ǜBGM��\	�=*���H���;�3��oi�{����@���6�>��dc��|�
���J���;�3��oi�{����J��H��5Կ&1�sW�L��"<��O��5Ҹ!9�{_�E��(5��M��3Ժ":�x]�D��)7��Ht�6�0{�{�ȿh}�F�F�6|�1�4s�w�ǲdv�M�M�?t�4�5s�w�ǲet�H�E�5~�=���I�e���cB����&:����B�o��dB����#?����C�m��gC����,1�����NSw�Df��μ��"Ӵ�^ϗ}�Cc��μ��"б�VƝv�Hi��ƴ��'ж�^ϗ}�-T�@�/!G�|��t}S��U�(P�B�/!G�}��w{P��[�&X�J�#,H�q��p{W��R�-T��U� +�"l��U��Wb3!�V�!�/a��]��_j;&�Q� +�"l��U��Wb3#�Q鳈%S2	7��Rf����2��/�	*S3;��Zm����8��.�-[:1��Pf����2��-�-[��Ft��<wM����$����O|��=rD����.��	��Gv��>xL����+��		��FtU�Z��P�򚟧��l���]�^��V�������f	���U�[��V�������c���X�P�)QS��o�Fj�����憎#]_��e�Fg�����根&\_��f�@m�����⥲(T�	��I��=Z����D>�{����L��<Z����D>�~��
��G��7W����O4�~����C�}�-�K��Gi6.L���Iw�x�/�K��@c? F���Np�q�%�C��Db>%A���C���CR]S���(��H���Dt��GWZ[���"��D���H~��FQ_S���(��H���Fw��KX��Vpk���
�宝P �,'<g��Qwl����署W&�($<e��Y}g����箝P �,'>d��Y}zp�F�-�p�]9����w}�L�+�x�U1����zp�E�&�u�_9����zp�F�q_��3�t4�A6Y)2�q\��	?�~=�G3\,6�p\��	?�~<�D7Y*1�xU4ٰx;n�<'�,޲���?[+>Ҽs7e�6*�!Թ���6S-;ѽs7e�5/�(߷���5Q!7ڻv%�#�-�ZĹ�S��l�Ͷ��>!� �/�ZĹ�S��l�Ͷ��<"�%�*�]̰�Y��f�ű��< � �"��n�)��5֨�٤��7V�+��j�(��5ת�ܣ��9Z�*��f�/��7֫�ܣ��=\�"��?���J�9Pv>Oثv�mi?���H�:Sr8HУ~�en9���J�9Pv>Oثv�mk<�����L�?����G�l�1��v��A�>����E�l�1��w��D�9����G�l�1��w��D�OL@�n�O������W��ϚHID�l�O������R��xȝOMB�j�I����Q��xȝOL ` �C���z��!j3F�G:O��9���!%B�C4����@!�\!��L҃u��L`S�ĈP����@`_� -p�Ȋ�4aH� -O~-�\w��Dxc�Q���Q��O/ᦌ��ʄ?8^�)�ҫ�`8���n_���t� o}��^$C1����U2��� ̋9*�M:L�`����qP6���'p�.�!Q)nY�% @,D��j�j�*#p�'E��z�*�#q�?� '�v��ɋQ�H���@��Jɥp�N	i'�'���.�t�2�(1$ItR}h�'N����Ӵ)������[�B��� �']ZT`1���� �79��C�'@�{@����%�^�#�	ū	I�<y,��7l���CN;_g�iR�"�F�<a`bǐ�ٹS�E�I�ZM�'F�C�<��J�*��B	��QF8�ȓN4��a�E'yA*�Ad��t��y�������A�m�#��ه�"Q���r�M��`=y�oڌ>��Q�ȓ3�v�2ՋPcq��a�D,Ɇȓpw�ТGeݽpfu�"Q<8�d��ȓV]���G�2R��m���#�h ��������c0�[@��5 	 �ȓ$�r��_!jԀYa��3kgI�ȓRժ$�f	�_� ���N�W�f�ȓp�xUpB��	-t ���	[B���ȓ4Ֆ}aDJ�,L�|u�G��\hԅȓ	Ra�b�
�- �-r���ȓ�"��� �#$����բR]N<��ȓ\.�@��5d"J��`H�v�чȓ7P����)�%Gƚ�!sˋK�]��0Z~�#�,X d,�]�0��2��t��Hֺ�h'Vq�J�0�ĳ��ȓ.�M���U�J��U���@ T
)��{�� 9�@# Єӡ��Af�ȓ-���I A$�{F��'�&͆ȓ���d�Z|�%��>b�b��ȓ3\����
76���b"T�J�0�ȓN9QV��	,�t �!V�	&.�ȓD��t�퍨"p��m:p��݆�e��|��%�+L�a��/=Aj��ȓa$�����R�,\�ߨMÚ���0�e��!f��u� <,�ȓ�H�.�,+C$���L�w�$Ņȓ@�n�
�J[tN��쟪Lt��_Y��c�K\Ȓ��"-�-�ȓb��1�����@���t@@��ȓar���A�"d�0�׭~�`܇�;�V-���A=��)(B��5y����ȓ$Ҋ��G��,hrĻ�M҄i�R0��D��"�51�>( @ԉ`@B��ȓ��ՉR�& ����k�x/\؇�t�ԑ DT��(B��N�ȆȓTmRuaf�y�����Ó�V���ȓgO#Ԡ|G�ݱ�.�#�TՇƓ`8Y��&ǉ@z@�3ccǥT�d��r��nkp��GD>27t��D���	 M�9(tB"��֭0�x�g����1�T�Z�D̈��Z,V��6�C%Oy|[�L�N^4���"���b��ƊE'�i�򅙭*{�H�'�JL�EK�YP�ȹD�0Pi2�H��)֗����	�<%@p�*U�7!�[�:��GM�?BQ�� �×V����P@�)x�(�4�u4`Q��EAo�0W:�0�f+�� ��#L�[ZT�>y�C��.`�OPS��L�U
I#�/�;hc*�k
�7�<�%���q�Ҙö��3.��|h�w��E��ӛ>�t����Փ`.v��	$*�>��,�y;�ɾIR�m:Cg,�d�*��D8�p���̐#|_�=V�\Sd< �W�=�=�-��+���Nq������n�vԖ'�6�AC��4���끉j�^@�k��0�l����[2���&Q�q��uk�jZ�pbe�'�p>)2��{��q��<� �����?Dfp<�0��4Ƥ4��@ N�$�+�fF1w� �,� ���_?A��fIX�D\#&<.(�jĪ*�X�;'�
�HODD�GN� @U╕n.���|�f#K�3b6��`�K�ЙXpK��M�`@��R,n ��D���^�(	ǓPv���aN��o�z����%t8E�؛�q����(|�TrǓ���F8Eܨ}�e�ނ&����H�emҜ� g��Y8�(���]�x��ՓE�	�Px�#��b�k��K�q�G�ޭ8�0E@1L�t�XA�� ������ө�(��b'+U6N�Y��m,�y�����X9�F$ο<2*�3�B$�0>�a�\$4�!��VS����❶:\�yc@N��D�Da9U�a�\���
�l��X�+���D:ow��� \q�$E� /���e�#˞�5$V�p0�̒D�F�{MD��C�0@
��U��캓�"��B�kѨ�$q��8B	��@�S��&��Ε��R4єÙhX����Q)I���C�Uu @�8�)�>^���T@��;�J�(��E�&��读D�")�+�>R2�=XaH&3�t%[�N/R�\����ڱӰg���B�y ��Z�@�60�p� �(^�i�wb)E���9 �<��e]�{%��b��Q<&�SЉ�.R�Y���<���!�
�bQ �V�-�B�3�*:LO�yQ%�m��1 �؁ICn�S2�e�����&�)��W�'D��A&.Q�Q�t�SrOY�LH~��ɚd�ѤO��9��,��=)S]>����i>ʓ;�����(��!#�?����O<��� �P�#V���Ҭ]VQH9�9�G�9S�&��%����d�T�F��$��d/V�x*!AiI�8<ȍ�RI��}�`]��⑓w��\��#��,�0ӏ��')�QA�'�uCR(s��v59Ђ���~�Q�!h�@�k�@���ʛsמ�a�oV�j�h�\ܮ�1�4�M�!@��C��=��G�w��H� ۦ���\ڦ�y�-բL�}z�Ł�4Y��K�h��@�B���&Z�y�(A�D����- 8\��@5���"�dS>O.��0�5�f�ױ%�p6�B-"=R5���A7����N�D�V������g]�c'�&��O��"e�,�b�e�� �,"�ģGk��+0h���RL˼z���� ¤N��d�`MA�#ƶ��ӂp���F�@�{6��#7�ؐa�J�<���r���&.@ z4�c>� �ʎc$>�`�(_�tI�񡗎q��0���'����A�֧n�g�'D�̛6,U��(��f�ިZ�dEE$�k�\%ّ���lP�����O�bQ3�$�?o�B�����/`�f,����N�l�S������'�0a�U�j��gN
 *.+g�� >�@TbD��=p��X0��p�z��'RJl)��gΊ&8	'�g�aR��@�*(k��3U�F�y�#�O���Tb�9(�� ���plB�o�C���A^%jV(� ,�&g���s��߲(�h�"	�tdZ��=B���!�$kR��#`r��{@��&�n�����+��p�&EB���1G���=H��Pc��jRb�XT�/m��+f�K�7Ɗ�9ūY>\]F)��[�`S��R3��W��͓EeU-n��G{���~z�04��d���@VkƖM�&=�'G@�E�fp��\�e�lt��3||�Ti%e�ʩx&�FO�.	�ǂͮP횕s����f=���F�L�W$��2�.�9�0?�!�Ƌ%Z�q�!D-7�iZ���<�x�Ex�2���F�2J�x���C�O�0�6��^g�=�4n����s��]�@!4�$����p<	1�e-�8x�Ȓb$� ��ũb��hը	d
�Ɔ��ޠZ�!��W��T���G"gbp�QLͫa��(E�t0Zv�ǁ��d�T�tyK�^l#֑���1"��	zW��@wnTd�S�i�=X�@��[�q�TA ��I�4�J�+!e"O�|ٺ�AЉ3z�b^t:�вɑ%V�z����X=��Ë��O�y�o��!l�`1��]�\qJ&D�Ҵzr�Ќ26-ѨI��ᛴ(�UN��ٴLh2E�ܿ~�
�S3�\�R~�����u���)R�	 4��a��	&���-�UK�Ȅ#K20�2�P�ݶm���5�\�N8�$���O�I��(��PD��
�6�$�b'6o���h�ݮ'B�����8/``��`f�.}Q��bbd�����r��

l�\�#E��*U^�P�Ƽ <\	��f��l�X)�.AXx�c��m��f*ԑ[�8��'�$H�,m3נC��| �8���R6q4��AI��=��OQ�N�:Es� �<}�Xp�a� =���4*M#��B�S���5bW�V�EFU�TbY)� iz �٢tn��D
 �!� !V]f����)%��hP�AQ$ �9
��(,�J�
���q �#W^x���!A�$��d0p�ͫhѰ���`��G����O���G���'ݜ�t��2�0��є�ک��J�|����`�#	� q��
Z����ק�>�<���ѕ�΁��|{�����I��x���k�U��2U�	'9v`����B$�=��#MX+
���J(Ř�R�Y6�x��;���Gᘏ	�]:�#�m<�{�H,p��P1�]'A8^]��:���
g�،�y��U�MK��80Cm�	V0"'&� �>]�2���АD�to�A@2�RBQf8h�M\Dw�܇�M�R�
��D+�� z�ˌ�($t�C��Uv���y�,"T%�ud��	�j�`B���J� ARL�hN�!�rOژS[6��
0M?�����+���iu��j|�<��C�(hZ���O��VP.-���˰L4��������)�LC��,H��-@9b(�G-�*�4(:0-B�(���cF�u�by�⌃#��'�fiȒ��!}:�a.��.88��"S�n�}���?�|��2�iYPl�S���*\�TʗB\�4SdH�E&8����E�y"���Ł��w��y�rx�� �#ۻ_�Pwj�w�I;^�	�j�5-�BT�7�J�.<�����=-vU[T �,:�2��0*�y'6峢A4G����kR����ȇ⓿)ji#����:�:��
��z"0�;q[���e���:�(^�^E�-���p 8�L��ujC:+�衉�n��
j�3�l-X�4�o�<	9TI��P�B��,Ʀ�L0��〖V=- T�Тk�v\B����3@Q���C����'�T��i}2\I0mLc�8H�i�Z�Q��� ���i���t������w&t)��e� ;���j�X�IP' [�����7�-�F*F�eY$=*�刪N>�I�-� l�r;F���tS����>�	�(M\m��/�;4e�� ��YY�����Q;k�Н��H0����*^�4��ӆ��2j�� ���Z���j���;j��� f�8Vj��I���D�tH���Ge����plt�7�%���� >\���a��D]YSm�`�P��Rb�4�.	�#O�1ܾ=a���-"tL+�H=��TQs횑`�^��Zw�H��?]�t��Я3�@�oD+jz�a��h���۾���ٷA#,��@T�̀%��[�j�y*�A�M	E�ܔ���0o�%�F�2 V��3J�hY��Xc�Y�tn��s�E�>�Ҽ�ƅX�0m�1 W�
4-L�ҳ�M�MK#��=Ln�"EU�_��| RK	5���d&@�%^@5��kH�&��� ��H?Hf �AR�հ_��d r뛊2��K��L���ڤ�
4T�^-(D�_1�D	0�J�I@�t;�oT�F���(sፔ��'���#!MaƮX��i�F�J|q��C�~-i�l�|�ڝ4�ė,&�W��`Ʋd�I�@�HH	q"�-A�LKe�8���e����0k]ĭ¥��0W���Q�BZj�V���idB[�
�����ܨX��8+��?8��S@d�9G؄]a�*��Z�����N�E��C��X�v����%i�>8��Kp	�Aјe��m4x]j���;����a儩\�u�� �tN���'WJ��e��e���d��j�����EE+Z�Y[, �qE��F��R��ǯ�+ߴ�"�e��nwr�Ag��K1��+�LX�2i��X��ޡ0��PUB[�\.�x���,�~��Y9:&���U��!c�1��+ʺ^𔁛�J;]+T9j@&��j����E/��<*��Ӆ���n���i��K�G�sn\�"�1-��j ���2�{' �)�8���ʪ�����3�	�?�A�G�AgS�-�%%��=�u:T���P�R�!%�^Zf���&@J5X�k�eP�)�Յց<
�]t U S�V�!�Ŝ�75�s���'���V� t�4Ibs�!�Hod,�GN�C`*��*D��E�t��e�^�H�C�0�\�s��"TavU	V�U�U6�	#PK��;�:R&V���ك_���^RD��5�X�R;:\�a���T��ɉ�q��5O4��N���B��_4|��N"�@���)�/r�5I%���0W':RT��0K�#��� @$ӰV,0ZD	س�e˃zwn)����'v̲OR�K����} �)!�ӆO�8͢w!�=6�ԕ��� �8i�$�/|B�C-�+{-
�A1�O�:ժG!�=6ܪa��� z����a�>� _���jrGM�W��|8f�#���%�F�0n�J�c4��>N��Ѕ9��0��*պAl�Ի�@�#]��
�l�@��ɾM�z1"Q�<����*ջ:�Ĵ%���{�Թf�N��ػ�����[�j���oB9�ds�)��yr$[$)ѷ�Ȇ���!��%K�LC���yՔT�P� �m|���A4r8�-Ȇ
� �����M�l{���>-�pL.X�z y&��B��(r�'�t͊���R�� Je�J�` �k�,{>�4U�̠R| ��D� u��(��{?d�
��&���;gL�1NB�����-D��m��Ȏ=p��0����}4p�JL>��6*t��A�>X���� J�L6��oԶ6��r(�(�P�=�f��p�[�Pa7�� 
8 ��,�:�pb&�z����w�
=jʴ����
#n�l�7I��}џ,��� ,�ԀJ�I�d҅�\LْH��f��T���Y����p�Ė)�j�h��j8�%K�>RX��h�(e�bNO�x����V�~d�	�Ǔ=\��S�
.�#:�������!`-i ���M�c��<�h08�f ƺaza��'2���jF�"h1���$
��]�C���ce�!s�.�JY
E�z��d��R�\RuK�"LRtaiE�mh-0����*�d,:�J�Tฦ�VpR��'�bI)5A��ob9���+����/��@a��"̢�*��T=�"<ᒇ�MVz�� �.N�Ye�G)/y�)��J��t3d�P�:,~+Aޤ:�4�4/�5E���c�11�Y�/���O��"Տ�9�{#���$�pUQ�KH�P�������31�4ҫ����*ſ��\`R��ʈܚ�E@.#�F��"\�B�H���1n����U*�99T�'�	0��� -ppcuN�=�Lт�� I��PBF4Q�,�3(��+�)���-jX+��Ȑ8�l�w��ȃG"=׋G���0�D�K�԰�d�%_F��Wb�I9ʜ�$�\�\� �Z�.�*NP�DC��L��q�eIQ�Q�L���E�M>���4]>�EJD?I�h�x{|iHA�
T�
`R�O�K��T=��ȴ�߃A�[��	!D�s�jz��,ܖؘ��[���-���/����I�3���qM�]��芪-ؚb�X�J*,ۜ�h�+R,&d�$zqL@)����F�B����Dk	�#�J4[Ъ��yj0mڻ����1�X�w�ǑG����īR�R���`Í5g�J(�wo�1Ta<i�̨7�'��t�� Sf������)�;ebN #�`�.�)Q��	1R"�rr)��D�4�Ȣ�ܘ/�$[�"##�| H�(S���qr���,T�And�v��.eXig獝3�LM2���jU����$`�)��h�ʋ�R`�dl��v�>���
#]�!E�L$�,0�J�Z$����Pc�l
��ą��?�� �x�iǛ>z@d��$�1��X � L�f��#�?L���(K�t�\���G�Ǧ�;�wvr �.W�L�:��)~�TT�� �6�"�l)5T���.ė�uw��uyR�+y�RX�� ���)�$�T�^HZ���{En@�2�3F�9q���GR�d�4*⛖��&�������
�����6b4�x�өZxi��*��Z\֍���ʄ<��i���<Q�N�.�p���8�e,?��Gm>��EU0Փ�O�7����lϠcl^�X��Y���aH���<JF��
P<
��լΟ5��� ��o�!��A��(���
7���	q��;z��q�`L�BM�qtR|�� ���O�����Z��RrDˈ1O� Z�l�4u���)��(#I��@#M!`��Ps'�[��b2$KH��.����(AMW�����.H�>�R���Q��d!�@���Ȃ�oT�Ug�]5\�.\`�G;#���3U.�ٟ�:j��:��P�#h�2$}�J��߯ T���ǩG�&!���eݭ��[��bԈ�}�B����u�.l���M
T�B �'��w��5-\��t �~nY��_�q�B��	NT�z��֥��R���k9�Q!��M��!ʔ!(�0�ya��CyrhJ�m���У�w.�r'�*V�����Ol���߁R��@Q��Y_Ξ�����{U����ʒ���)	v��ǥރV��hq��y+&�Ƽ��d˟E)�1zQ���E����	J��a����IA��`������ĸO��]x2�Λ��P�$\�J}��X�}���9��ˤ-D֍�t�f���'����`���*K�,�yRσ,��؂DD������f�&7�&đ�΋.LJt*0�ڋLa�][wx���2�J���v��z�ZcD�:t��
<�X!�c@�t�L���D*B�	�`Ï�77�y�h<�u��x�`�G&���PT�v<q��)A?�P89$��\�����Gҕo��C�FJ:�U)�=~&�d ;�X<DĒ1X���Q��	(6t�t�˓�"�`0/�3@nȳ�÷K�1Ol���6IӶ1�k�
� <	Sd��� (� �Q�K���b�#=>4�;���#�@��K(>,�C�U�8�@b���O����'6&�k�?��`�Q������-5GB����'��0���Z���$ո+�p�q�I�9dma�״;��y���5&}�8R(A�3�bu��-߆�Tk�'���Ekm�:����d�uذy0%�w���EdS^-xMi׍[2PHy���\A:�إ�OٴuC�At���%��I?��� �*�㳂�k��-�!7�y��R9<.������џ�{q�H8`�6�9���'bFĀ�BQ����+�Sa��x{��
/��pJYyy��غ������;&�SUWjd2��j�5o��>_���dH�Or�q�T@��ŕ��/cܶ� �(�==e,0�Q�'��{x�@Pl�����Dw�I��%�u�
|P���98  `�7��L�8:
p�7�',���s�!�?W	2���s�4��;@��d��8�L�*�`o���P�h�z�!�dٺ3LBi	UlU�N��T1�S�!�D�
xV΃�5��P*�l��_�!�d�S�`�W"O4{��)�m��L�!�$�'^	L��2�9{�^��-;!�d��L��[���8���n�*~�!�d�"�h��Ac�:0��-̀0N!�,"Ȭm�eL�mU��lԄ+!��<M�j��!�ع;ZZ$ە�AI!�$mi1a�P�$\���#g�!�$��s�p��R���j(}� -V�@{!��H��@�
���t��j�'b!�d�D�dX��i�![��ic����{W!�d�g��Y b�C� ����W@�9.4!�
�>�����`�r����m�5d�!�<m�v��cC$Gҹ��&ޢb�!�d�AXH��H� {H�X��� _!򤑞'c|9t
|A�$�'��fG!��D���jGƛ����� "˃oH!�� b�f1RԢD� ��|'�ƤS=!�d��BH�5�04�"(�q�^1g ����+Zd`��J�@lq�陚�y�ղIo�	�K[�=Aܘ���_5�y�,L�YL�H9�E_!@"���$I�y�A̺ z���24d�@�1�G6�y2L�#e�;����`X��̀ƈO4%��EZB��	��\8n��v"O�@wHɲ�cD%
Ą�"O�A�5�F�.�~40�$%RD]��"O&8$I�-�r���u�6}r�N�@���}J�O$�E��EBV5$�H�]�v�V�U�]�t�F�9�BLn�	`�c(xBG�
��̦O�T��&μTnm%��?A��Z^T��ŏҫY�fe�w�R�����e�(]�*��?O,����#��:� r�`*��:��ȹj���D�$U��Z��I�
8ҁh!�����ä��#@�騐]H?I �]�U��	
�'(|� ��
�N�0��)�z��Ɉ��O�q�y�%!�f��*��ū#�Vz�çA�A��.r�1O�E���|�&
��[�zL���Æ�m:��y��O8�𩛦<I���ĩ�!<6	��Z�)��'yn�d�5���?�'V�T,B�팳R�fA(��_�x��'f��R$���G�ر[rb�L�́���#G�7mW�vJL�"~���֜>�����ԪuՔI2��4�n�����p�G��*�j��X��3urvz�a����d�
����ː+��)ҧv���J5�
=�fa;��X�&�XnZ^�d�K��լl���>0���?�9����F�Q;�<��)ʧ:�ܼa�G��L�|`��Ͳ������d�}��S1��p�-ͭ�@�"5���^��0�'�$�OX-��
�y�#L�77D�#Ũ}� �ɧ;ö�I�a)D�S�),�V2Lk\�"u�д@����΃?�h!oڋ_�L�(P?�#�S��I��}�`�Ǭ1jl�w Ͻ&���Kf؟h��E�A;�M
�nE�\�2i�T@.D��0b�ʗ;3֑SiD���@tm/D�X�$�Cw��+q��c��Dj6,D�x�c���Y�UIUհI�R| p�+D��a3��7��!;��+S����.D�� H]��"ԙ0f�˵i��7D�̲C"O�ت&&
��&��J3^�@i�"O>��6�T�X��x�o�x3"O��c�c̬2w
��-[Vp�=��"O��0#תKNڨ�e�J�6<F0I""O� �P�iy��W!:�x��"O�PI+�a�j�X�F��1�nD1%"O�@8WE5"\\c��<=��y��"O���e�+M���!G�]n�8q"O��:&�4s���B��s6��;w"O�9AG�-i* B#�?��x�5"O�����5d�+�cO� ���Q"O�1��I���xq�B1v��I��"O��qq���'jmZ�Q0F�έ[�"OV�j���!L���f�U���uP"O �Pcl����z�jZL���"O5�3M�	V)��3A鍏n�6��"OB��k<RV�aIJ+1��ј%"Oڔ�Ua��;��� *�����"O�����a
���hݚ>��+�"OD��pȒ�&�n����J�!"OȜ�態4l�I�*�..�VD"O4\ЧM�$����ci��R���!�"Oy�Ŋ�gU�HP$�X<+ZP @f"OiWT�8�5�@��}Hd�[�"O2�x�b��w�lD�n^�.Bv��"ON�&*F �H׮)}�N��2"O�	0���c��ɸn��_w"�	�"OP��	�����B�#��06"O �A��\��,+�S�O��@�"O�@aʃ�:4����+��#ֈ���"O���QmZZM.����M�J��4Qt"OR�q�"ے��a�'��z�ٸ�"O�C�ʇ7,�إadW�!xP� "O��[�$0 ~
�w�L<@�Z�"O����6V��
���C��0�A"O�q
�!��dS@�n�Xyt"O���1m���L�c�{@��"O�y!&H7��鱁�N�&i��R�"Ox��@M8��ǄʐuM�\�"O܄0��W�F�M�&��<.L���"OrrQ@ߪ	��5�`� 1|A�"Ofu� /I2; t��b�h\��y��i&���wN
Jp�x��'�y�K�c8,`�^(5���&W�y���@�=��E\�$D�P0C�À�y�g�(uy�M�B�S�!�!X��y.�7�ܰ��I��>��eN׋�y"�/#ft<�!oΦ�J��Ė�y"��i6
"� �J@XgY��y��b~�)"DZ+mZ�9x����yR%G� �ʴ�����l#�K�O���y2�%O�>ݠ`��c!�R�I��y����mY\���U�cr��$�%�y��J,&�	�,,2Ō)��ѧ�y"m�)W���zc���`	��˕�y�͚
kl�����JX��rc$�y��^6� c`dَ��W�yR(�)��U��]8`�t �C,
�y�$�0����"h��B���L�7�y�	[�X��y�t�P>@�<L��F��y�b�c:ص` Ǎ�3q��:��#�yr��a1:ʂ&'֜sA���y��TLmS�ᔀ�Z|k/�y
� F�˕�׏��-qp��#�<c�"OB��LD���҂8��!92"O���j�Oy�@�,y���"O����ܽӜ�j㡚�f բ�"O���F�w�ɩ@ǜBQ���"O��$`S�(�|�z�"�� � �p"O����)Җ~G✺���M.4��
�'��� �Ձ�� J5�զ�Z�q
�'cHMr�+�/����S������	�'\��äL$)��d����@��'�P�'���m����B�L�7�Fę
�'`������ .��鑊�\}�)j�'N�-hDA^�r�~U��VXz�r�'*�`��R�2,�T�`�SB���'�6L��8>ޚ��I;DSV� �'����w˞6a=X�"�c���^,z�'v �ӆ�׃9���v�� 8��p�'�Ac2�ԮA��z�)��qb�'d`-;���'����% ^�xj�'�X���hB1�R�8 ��Sގ,��'�����M]�o�@1��B�I���
�'5Va�� ]��jĀ�fФ	� �
�'y���T�4b���q�Vxc8��'Jb�8�łk��	��T�r�vq��'I�Ń�Iǰ1BQ���Q�S�tI��'6�Պ�7�`���C<vRe
�'����nS-9��'M_}��A�' �dG�C(4��PJ��%E٨��
�'�񑤙"ߚ��sD�j�X�
�'�R�c�O�`<pt � &��K�'����3M�p�й$�Bur�'.,�!�OZ:���@������'J(����Q�`���¨q�L�	�'���$��?�����Y��^	A	�'�����X�h���ԡ\�Ih�]H�'S�� �e��5���i��>�e��'��ivk<+�<8CR0#"����'��At��1�.4���M�'_j��'���$-	�v���C�	O=F�A�'N����A}_�u�^d�y��'�� ��/Hwp`�.�(/9X���'+���d��U?L�Еiћ&���R�'���gf �*����S3g���
�'��������
�g�K����'����@��cq��KB�Hd�ր�
�'H�c4��)v!x(��@�q2蠱	�'��	kF�&�2�(��(h-���'j�Cb�: p��āY�n��' �ȇ���X����_F����'�4�S�A|����DQ~`$x�'��u�և��ht:c�6[}�=C	�'���������( `B>J�b:	�'��Z�&ؓ�&T2c	4J,ؤ��'yIĪ��q�^��HAJs�Q��'
�I��@�2Vʰ�� �H�(��'wzU�@��54�(e�S?���'���K�I�3g�p z4ᗩ(5�A��'���E�A�fvp�#���60N�p�'��4vɃnY��c��<���'���lL5&�B=�0*I�K}�,��'�����#'"h{�F�\ub�'V���W/��o�ց���%C[`���'��
��(Rb �����A�<��'-�(Z�Oݛg]8 (B"[�@>4����� �9+î�h�%@U��'�q"Oԉ�&��!|n,��b}���"On����� t�bP�S�)<h�i�"Oz�	�F�vգc!T6fk����"OdA犅�5˵���~Q���"O�%����)H�e0������a0"O��`c��x6���Į]�jf���t"O�P2�H�KE5K���yc��  "Ol�r����@XTnP*>�p=�"O`�#�`)>Z��u��=+��!a�"O�x�1�F?"����	NM>�� "O�Py&ap3��Z'	�	f��J&"O���#�����P�@��"O��A�	*9����\(�@�"O"�Q��D1~��DފTG����"O� ��U�#)��`�S,�`0��"O�e(�-ڍB����7���B���"O��Y���[��D2�*֕)���C�"O
P���zx^�3qkD9{��\r�"O�@bV��9���w��Dx es�"O�� i�$PyNXyԉ9o�9(�"OZ��J�c��ո���|]du�#"O�ݛ�E�$9�Q��'��F]��r�"O�QB!�<�a��CPD["O:�;���'�"M����A�<�"O8Ѩ����+Z,9J�E�Fbi�R"O"�+Ĭ�[�����c�$a�6���"O���k�4��M����;�X���"O���V��2Ox�� U@���x�"Od]�G��&'h��i%�P��|0 a"O���baH�0�B�ڦ� �:��:q"O^p2A�8]�:����c�1)"O��D�?}jV,(g�3 ���P "O��B�"�"N�(`�&V�_�&D�#"O�����!�VD؃�I��`"O�����i�ⴋ ��?�|p"O��j��? ܔ��K�h�@Xr"O�`��< pq�!� lZ.mQ"O~h*t̔*/b�Q8g��u"O�%hQ�;�M9�M0yQ0�8"O<%�c�rA����s�n�Za"O5���>GL�9�we���"OY¡�X0pLN���Pe�ԭQ�"O�����t�JPN�u�I2�"O�}��@�/R�����a]��"O��h)E��P����8gSNt��"OT)B�匔d�����ɍ�<xQ��"O�5�m�0��X����,j�t"O�t�%��9ؐ�IH<T6,q5"O���4�=���pg��6b��Q"O�1��� T�:���G�n�d�C�"Ob<���J-fx����^��0A�"O�\(#�)Ln�I)`�Ғt�n�I�"O���`���������A*l��"O��s陜/�f�c�+q�Y+�"OeS`�3f����gK ��� "O�����nK�	G��1L��u��"O$I��J�� DN��o;�p"OJ��%BT� Q��G��wD�XW"O!�s �)GĘ�cG�L;� ;�"O=IT���l�`Ɔْ�m�@"OVP���������SB"O&AI�@�{� P����d�uц"ORؐ#L7�d4#7�2�0��"O�~�s�   �     �  D  �  �+  .6  �?  IJ  ^V  ]  xc  �i  p  cv  �|  �  +�  n�  ��  �  5�  w�  ��  ��  A�  ��  ��  c�  �  ��  u�  ��  { � � � $ �(  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@Eb�?LFq��J��� J �ǍR��B�I	_h�I�4ę3C�����`E+.ސB�I��{�n�u���ΗiU��F{�O���D�̈I�e26��a�ŒBf!��̡*I��b�η#�I�Z�-���'����ۤX�nB�kc�p���!G4fC�I 2��XIS��E��UQI�$V~����'���}r��L�Z�S�K�O���B'K�Z�<������	PiΗy�~,�L�a��v��:�I�C@ d�NƤu�}`E�-D��)��a^���v����fTx`�/�	X��z��

X"�ys㈍�()Nl��#�IO���O@����@}flB��J�5�����'*�1��
�')|�S��Սw��y®O�b���I����y2�Ƌg��!NE�`��S+S�!��!4����ΒҤ��l��n�!�ʻv >��>H�t����{B�O��S�? �UX%��wB�)K�D� �D���"O�xqD�H��鈒�=	z�t� ��N�O��%��آ!��(@w�N�e� ��
�'w�`�3�O�;|lȉQ�X�*���=O2�����A�{� �h��@�P�����	D=!�DC�LP�o�����GX�!�$�-)ˈx���A?J��rF�  1O�1ڴ-����^;O!@���8A_��QÅNTU!��_�(]��b��{�F��䙼d�:!��)��<qr,S'o*	�P�ܧr�8� 6}�<iU�T"e Nx�`b:i�H@d�Sxy��'v eB��`�Z���l��V�	�'��KTC�F�Z���fGVx Z�'	�<�Cn
(p��˥�8w��J�'���@V�3p��U�h�����'�2�Ѵ`W�P�b�T/x ����/�pr&� ��J��j�A)U��%�ȓ%1 H�F^
-�6�g,�9u��ȓ�-r�JU]� ��d�y�X|��8o.���,A>s�
Hs��D��Ⰶ�"DPI�2AӢ����
�%��%G}b�i��>%*F�]�J<X���Ě$@�A�1D�T �g͋8B�#�GN&)���*�O�O���DM-�\P�I!Rtp���"O�|�uɜ "c���!�<_�Ƞ�"O�,�Tm�E���i�� ?�K�'D�$W��!2po���.���Ǟ0��;?	K<���'u0�RWDx�Hv��=-�>�m�E(<��I��(d�k��<k[&a�5%ޯX��b�x���,8o�8��� , <
Mzf��&eb���$񄨟���g�qyp�o��$�<�"��%D�0)����̘����L3��z?��b���Oh�s�aD�Q�HL��^?a y�'V�<@B�%"���(�:����b�6D�D��j�  ��LN�P�D `l)D��H,�>��d(TIL2C��|��(D��ہ�Xd\��'�����+�O|�r��f&��\.�Qs답|݇ȓ/�2�b]�+1���CIQ�p�ȓ@���yvʞ�>��S3B�>'5�ԇ�x�\͙e��$R ۤE	�~vL��<=$�c#Ϛ�J-q���K�^����~E�4D�aj�L�p���]�H�͓��?a� ܎1s�f��4�L��b� a����O��!�ON�xTd<��(�Z% C"Oj�Z���I�:�`t���	041�V�U�Q��F~��>��xئ��$o��31!���=Y�y���7�a� �E/I>�C�/��'a�z�#�6l�H��L��I�1A�ӊ��'ў�O6f�:e@1��L" L�}h�+�4GC������3쐥J�B��?�዆�ĥO��Gx��@Q��~��L�p�ia0��u��j��[6�ybˎ'��QB̆u�*��4�7�$b�m�F����wht1��m
7_�Z�I�ʏ�H�����'�D*��ܶì$0��X:�}r��d;O�}�p�I9d�0�Z nGr
�@��"O����'7J։2��C-K����e"Oay���%�b6jA�(�X��d<�S�әp�>\���"pe!2��:2B��3X]^�#��8')DY��.	2"<��'�2���� c�.�$J�9[
��
�'�\Up�
PX��%�֤�&8��@!��eH<�P��8U̬�B��Y�H�h��OIx�<Gx���e!r��j]�"��$���y
� �Y񥞰
O���ccl�`�"O�Cw��	�Z0��)��uN^�+�O�t��9I}��CEEo�Q:��@x�<�dc�l[�-2�NN�L�%Z��s�h%��A�O�@jfE�>�MҠe�.�2u�`6O�=E�DLH�/	|RfF��+��K���O@"�3M�>C�VaI���}pu���Q�<��B0;˲�+��$M#5�CK}��)�'a��|�F�ܞԸ�#��(R��\������mC0v.�)箉�����'p%p���;N
0�q�Ӵ1q�(���ybo6(R`DP����ھ�yBx��ĻM�Wf@X�����y�$�/^�jbH��U���Z7���y"�D������L/P[� �_��hO���iY�Q`Ș���K�_u��`�2�!��8#���K�O�	?f&I�Q�G�R�!�$Ŀ$�EY�����QS�OÀL�!�$ F.T �S��cϢx2�.��!��H+�2�9���5؆��M�<?�!�P5l���a�
�D��j}!��0A�B}�FJ�-�u���A~!�\-�Is3�?�&0���B�	�>�����'�y��`/��`��B�	�B��50FB�-Fc���(Z�^�C�ɇ=�a���O2~�����X�C@C�I,Q�L�V�i�HKƉ-�B�ɜEj�a1LS�	��kw�`��B�.]��u[$k�7�+��V�O�B�	|�\�x%�M��n�"De
L�XB�I�E#��At�K#..R�HW�ɔ�JB��@�._	2�h��.�vB�:�l!Z��$&$�#�
'Wu�B�I�n~Bز�ߦ:��<�g䄒G�B��1-|��:s��6P<^��ݰi�C�	
yp�8��j�)���K� �y�B�	
Z�8e�sO����qeG9TxB�I�f��Ի�άB�P�k�E��vB�	>:Q� ��!B"���e�6�RB�	�`��L���J��H�����X�B�	�El�KB��~�H���*�<P�8B�ɢ67�Jա��I`�ء���I��B��Pr~Yj��-\�$YZ#��} B�	���`�P���� jrn;��C�I�h�vd�CI�_p�lP���YWB�I��r�H�Bيz��@r̜�[r�C�	�}�	����8`�$�Èٛ�vC�	�=��iP �� W��h�h�S�:C�	�1ۨ���O	�`��c�\�`�TB�I�ܙ�,P2V�,��D�G:~P�C䉰g�Y{��wt"���H3{�"C��S3Nh�D�X� %8A�c��?aBC�I�C�a��k�;�.��TB�I�`���Q���q߸��Q�C�w�ZC�ɈI9R����X��I�QD�c�vB�	�v?*�j�٘2R���6%ک/#�C�	�S*� 3�_Z��(�.��;��B�IJ
�p�&XV�zِ#�RzB�4$˴4�e��g�p՘Ҁ��ÊC�	�O�f̳�� ����d*�>Ki`C�ə1c��`<N��i#�ۗf�B䉮ry�@���O�nA*�# &ZB�?;r��v���@���sc@�&B�I
 �T|���Cb�� �ʗ>��B�)� .�Y���Rw4�04O�)Y6~9j2"Op�BD��,�6l�2.��1.r|K�"O�����
7X[u�plƇO(܁��"O��` C�-m&�U`ÍV�}��Qq"O̭�Ab��-�a���(t�91�'�'��'�R�'���'_��'O��yd)ۃ<;H@��	;���v�'���'�R�'���'m2�'NR�'����j/Bܐ��B�Vu����'���'���'�b�'
��'JR�'�����-6�h�����<�[��'>��'���'�'���'�',
�Pb�?S��'g:U��(f�'!��':"�'u�'w��'l��'l����4p�m��Q�K��pJ��'N"�'���',R�'���'���'>���f�1k��)!�/�`��B�'��'R�'LB�'���'�r�'����������X�[��j��'^�'�r�'���'���'�2�'M�@�E��,������;DPX���'��':�'�B�'�r�'NR�'�� �A��)`�k0�
-$**���'+��'���'���'vR�' r�'%����㞰u|��5�`u�H���'�'��'�"�'JR�'2�'	�1�7J�+)��t9T�_ظQsW�'�"�'���'��'�2�'���'�\��HE�P)�=��L�;�����'�B�'�R�'2�'�"gk���d�OhH��lڲf�ʀ�1��k�d�"��Dy�'{�)�3?Q �i����l��I���ۂ�Q?-�U�ǌ�9����M�?��<aмi�9`D+�=�x�UFȳ,���Mx�B��O�=�y��,�F�N(L��!�~BR��($*4S5%۾DeF�:tG�b��?1,O��}��eG�q��aw}�Gm�^��	"�i☁�y��	���ݐP� ��P�7Qn,���3~���4 ��F5O��S�'T��@�/V�<�u*��.ݒ���%B��aB�F�<�p�.E��8hBd��hO���O\󐈋�g���En(`b=�`?O����"u����'F��%��Luvyq1�-.(�h ��Mo}"+v�j�n��<��OܣФ<`4�!��8J�1h1��hhF�C5m[�X�g%�S+hQ�h�b��<��OQ�K|B]�(�>\��k�� yyb]���)��<��J_�_P){a�E,�杉�̈́�<1��i찚�O��o�i��|��W#�5��+��zwXĘ��\�<q#�i�r7�O�D{���S����;�|����+��T�V�ݬK������X��$�v�U���$[��$?!s�c�Q��q1�-άr���7?!��i����y��O��OBD��鈹|�b���>X3`@�>9��iI,6�i��%>��Sޟ�C"�!2fŮ~I�5Ї����+2$�>q�>���З��	ш�'(��SFܱ 퍳�,��!O~Di����<aI>!V�is����'��e��'�������Z�c®lr�'<r6-�O�O�9OpXo� �M���p栥rC��+2jM� �D�4_��$�T6$Γ)A^t��
�L�E!c�?M�S�/���#_cT�����m���!N8(�`��'(r[�l�����5�'OA,:��j�/��7AV�Y�S��m*�@*?���i��'v�9KN��~���mT����+R0O����&o�d���3j���3O��D�.c("L��CO�Y�%�m"�`$M�|G�`;��|R/O��d�%sq-�P$��Y~jd" .K�<���0�$�����df.�	V��DHz������ �Z��fF����ZE}bjc�m�<�H|��')�.�(���%��BK,f�LT�r�F
c��uo�K~�O���Y�m�*+���(�+֕2R�S"ʞ�k��PÇ퉰u�n(C�Dʹ�8��u/F,N�Z���4�(I��ɋT6Q� ��%bV��{3+S��?	VIül��E�ӯ�2=P��c�G|	RFÚ�>�8Qk�&����D�/ �Iɀc�������L�WTL���Ƒ�6L��y�m��(�C�1C�$r St �غ�[Dc��O=;3Xe!�"��qU���qDB3|��P��E�Z]�B !>��"���`��TiF��=C�\�I�!U'��Q��N/���?����?�/O>���O��p�O95&��tR�@�g'�c\�O ���O��ľ<�Hݙ 5�^cM�A��H��O����p���þ�˯O&��OړO$���0�'��ݐ��P�r1�PΕ����p�O���O��D�<I��*r�O3�L9��ԃbc
]
Ġ�ECN�@�z��$�Oʓ�?i��M���|z`j[ �h�Ѣ�ڡ������U�ӛF�'Q�B��:�ħ�?9���sd�8¬\ٗBH&>x�!��i�'C��'.`���I�EB���o�.��D���ȑ�M�+O�Bu&NΦ)X������2��'�� QH��g �*��/p�3ݴ�?Y�x:ZQ�-O��?O"�$�\!Wh ��M *�̹��i2ͣD`m����O(���ء%��7!;��-J�e��(��CY����4%���+O����OL���O��ƢLWP|U@L��.�<,!�Aۦ�������6���s�O|˓�?)�'���� b�,M8`�$ �$�ڴ�?�-O��a�9O��͟l��m��I��^��/�!?�F��"Ԧ=��*Cԅ!�OB��?�+O@@��h"I��M	����t���O2J�g������O����O&�'�ΐ�&C*?�Ȉ(��.u��+�NNQ��cyB�'=��㟬�I��t�	� �aSkY��̍`u����>Ě�<���?����?�����$1���ϧf���b��'o�>�2*���z�oqy��'��I�D����Tؤcu����!gN�+t�[<91:��r ֍���O����Ol���O:���,Cܦ���ϟ8r��]����a\+4�����/�M���?a����d�O�\��=��'��7�_85Ɏ��R��5�9Jٴ�?i��?��i�qR�i�"�'jr�Orā�s���&�x��V��L���Bc���ġ<���Y9+O.��|n�BK*�H���Y��|@6�\�boP7M�O��$\و�oZɟ��ٟ���?��	�
�IR���l��iaWl�� V�0�O���I�i\L�&�4�L�OetH��Dm<yB���utDJ�4bY�,闽iS�'���O�$�'��'�x���С0.EX��D7wm�
�Co�,H���O���<�'��'�?�EH
�3޵�pmB���!d�/��f�'��'4��q�r�n�D�O
���On���dȰm��]���A`�s�@��rU��'Y��i�O�i�O��$�O�Ev��Y
D�k#j���3a�Ҧ��I [TM{ܴ�?I���?��a���}?���D0
�FurbI�"z�n��qJ�L}��^��yB[�|�	�L�I�L�IRY���T�̅6�ju���hTN��d��M���?��?qY?]�'K��Y:a���X�I�{��,��Hba�E�<����?1��?Y���?!��=��"V�i��xj��1����A�
D=d�k�-bӬ���O����O��$�<!��\��a�'U;v�hf�F�N�>�S�Hl����Q���IğT�I��0�I�g
�۴�?��b�C�eV��F�zj�8h&�i	�'��P� �ɐ8����<��I?��j�e�l  I�[��̅oџt�I��d��.c�\�:�4�?I���?��''�p�+�nQ�U'z�e�P�e�|��i�BU���I)Y���՟�����491b�/��Dyp,����!�"�����՟|za��M+���?������'�?q���Z'�y·��:21Xm�����s/�I���ã΅ݟ��	my�Ov�'@�����/CM�n\ �Ƌ%:5 �l��mAޭSڴ�?����?������?	��q�̸�g�'X)��B|�!zA�i�H"q�')b�'жe��O�O���Z�Q�jD�cW�|��53�r��7��Oj���OʀYR�N�������	����i�iK��\1*	N�+�K�[�"�i�h{��d�O^����(E��?��՟��#sLX\�l٥Fp*�r�@�%^�iI۴�?���(M�v�'�b�'���~��'7�q��՘U�S�� g����OV��R���Iٟ,��������'�I�R��d�wh\0���	ӕ&w�3�4�?Q��?���h��SEyr�'Av	¤�>:��� �6�13��Ǽ�y2\�P+0#������L�I"&��ٴ��H�f�o�����K��pr3�i+r�'�b�'oB]�`�I�!V�S�0˴�6�Ħp�T��Qʂ#L!����4�?����?������d;��$>���(���QhK�_�`	��(�M�����?�O��������	�,���Ŏ�#m�V7-�O���<	�b~�O�R�O<��"b= �v�i��F1+�2hQ��/���O�D>B��8�p���<��M�W,F�I�m�Wy"�M;j�6�Y[���'��ԣ!?�I["����]�'QxG�Ԧm�����'n�p'�b?���F��H��-'Z�e!��|Ӿ!
� ����֟t���?�#M<��U5�ia��ǑFf�RD�!榔Ar�i�L�����Sӟ�7"1�`�lP�k�Y2�Ȕ �M����?Q�A�8���x��'���OШ�`�+1ڮ0J��i��i��i�'\��X�����O��d�?}	�R�M;���,WVj�*��j�t�䋬�f�&����ϟ�$�֘e|��҆�(�����
##��F2̓��D�O��d�OT�<�b��Ϟ�HM�bN+m���&��:UC�'�R�'��'�B�'V�9��kX�y9���f�$:0�qp�"!�y�S������8�	OyBc�?�d�S�nO8�;�(�O������nn(��?)����?!�}�c�%�h �G�_m2�ّB�x�
��?���?)-Ov�j��B_��1<�8�j��\�8s�U8T�Ե�4�?�O>a���?���<9O�L�K�*(��s/�@�$Wɛ6�'b_�0�p�A���'�?A��P��|�'dN�_�j]�A��Tg�iz%�xb�'�r,�`��O�S�o"LQ �m���n��-(q6m�<y��Ĭ��C�~����
����(  $�>\@sH��Z
�Q�@m}� �D�O�!0�8O��O���ASt���4Iv���fߟl2�PѩV�L��)��ٴA�%�A.&��.���hO��3F����d�~���"O�zU�_�U��	��;�Bu�J��]ԥ�`��Z��pز�Q�p�ܹ:��Z�A4�ɔ�	�'�2��H��I9��B�b[7%h�E� M^8*��}�fC(=��B�[���5�CK�*0U^p0 \�:TԥA�ٷ6����dF"
��`F	-x$��q	A4=2l����'�+Sg�O����Op�dF����?)�O�@O�/-H�0�/B�zGȸ�f˓�h���� �#�����'�� �6�ѳO�>����_�t���&I�^#Ľ���O���
[�0<!a�1}�ft{����7ݤ�a$�w��ɵ�?�"��PD�����	�$�"L�D�<!%f͹$Î�	P�X�UE��+cA�*��O�Af��	��,��ԵMe��2�C�1X�q�T%՟�I�Y`��I����5dT�È!�����h��� �� ��7H2���P����I��M0O���{��8pEk��\������m=�hѨӭ:�+�Iܦi�q�e$���>Q����i�4A����'O��������&�r����'b�'I2�'L�O~b�'C�3�5R�L[�ؠZ��ċ�x��~��t���ȇ,
�̉%aO"K�Ե��m���}�'`�[6�i�����O��')�\s�X�����3.���Ư��(gNlJ���?�#f��\�J���@Ƚ��T>A�O���o�bBL��W��>�i�O��c�HȨ/�,���4�'X�Hq@���_..��F�Z�[
 a�O^T 7�'������\4���ɍm�6y[��.c��!�<����<�A/��\P�T������Z��?O��FzB��S~�I�	�/ͦ�r)�.q�`��?i�n��yBԅ�*�?���?a�ֿ�R+�
 [�<�2�5��ѡ ���r�	Q��3�l�@���)eN�Ҋ��L }rE��{e�ׁ���,��KU78���E@L�{x��X(b׊�p��d�%}��Ei�*�[f�+c�:����T�i)���h��O�5�x�0-!�Ю��Ģ,މ0�l���(��:g
{���&�p��8��?I��)�/OzMЫ�]r=�sBC�|�zsA��l����O���O��D�к����?�OO�@��kI!\[��MW.0J�.�:A�r�Z�'Ȓ�0>�ĄY �z�ڶ��9h�)��DѰ~���rLð}ytE���cʐ[���E���(i���>��"h�O�|l,�M�����O0���̉A�IF��3��ȓ��2D�<�4�&5?$0�� ��H�$�1�ɚy����<��H;��ڟP!��
2٨F,͐?����P�Pǟ����U��<����ͧ;Q�8f�H��y��F\�9��M7�[HA.��%�K�a#��󦀎M�Q�574�P�ӯ3,���C�:��ݨ��?\M���	�����G�/t�i�'��0w����a!E�J5@dt�ȏy"�'k�yB[	?�� ;P%�b<�HQ��U+�x��dӬx�চ�6�.��w녒W�T�X ��On˓9�6;A���t�'R哝%U:m�ɳd���!&&�d9�EѪ	�	� ��X�3�q��* ���S��R>���lߚ`��h(S&g�p�03}�a�:{V��Eg\�iW\%*@� ->���a� m� :YHZ`4A e�$�W���'��>WkӠ=��m�'*
Y�E'��V����84����L��AP��!&�iza�Lz���4�,ғ`Vt�C�N�7���[ �;C�9 !�is��'L����2�؁ �'9��'rcnݹy���(fe50�L����^�^������?9�NY�Ȗ��|&������%�4�0�6I�A��n*����L�>��X���`�>�$��3�6�f�ڄG��ˇ(������)�3�đ�Q����5��78�q ��գ�!�D���c$�G�/)�)`0o�q��D�O�yFz�O��'���dQ�(���dέ(�tQ�CU�u��qA��'i��'(�Eq݉��؟�Χv��@D��3��`Z�`��?���*� NW<y���;]�h���qИ3H[9�-���^�L7-݆J�͢㠑W�1�����������\�:ש�4P��m��%4��܅ȓT���2&486ܬ��c�-5*0y�<A2�d�I��o�ڟ|�	 ��Q
�� ����U�X�>��	័�WL����|�4L�ܥ����j��9�4����(��5�p��u��>Oʊ���0!>�Sv(�1�ع*��5%��=jb��=p-�����L��.��n�ᄙ:A�qOt�pR�'Gn7�Ԧ=��4A� ���^�$�3�ǚ��q�'K��S?H ��d@�'���ٹ[ɰC����M�P���"H5h���ׅ\��|I��Sy��AG��7=�,��|��
ݬ�?������y�(�w;Hl�1)���?!����L�$��>)�b�s��ьmx7]>��O�=� �g��ř�6bܬPM����L X���?w�D�I�L�`�y�Ԡ�mQ>	p�Pr��gi���O��Q�'F�6��Z�O��m�LI��`e�G�bM��ksIԗ�y"�oaTo�[��'�Q0%��;F�i>)����PB��	s�?j��	���ŏK��<l��������W��8��l�	� ��͟�]>_��U�1��G_���W���|]�6�P�/��	@�efQ>�h�~�'Q6>E!R�s��
ef23��
1j�<lȁ�0Ǜ�cFڑ:�./#��|Abǒ	q���&A����i�KO�|�wazءF��<��Z�6M��W�g�(��'Ќ�a��|�����'�X����'cJP�g��"6�����''�(`�c�&bӶt�	�&*�T�'24ғiN���'t�,l�\0S��y�ĊJ_�U��
��M*I�	˟T�I�h8Yw2�'5BM�,8 U	;U�Y��4@�ET�1�� �b����M ��AQ��a���� b�0@B� i�P�h�Z	���2��	��!�Vq����FذAE�� :�'�Qł?p�Q�!@3{G���A�]t"��D�ަ$������$���I
bqH�Ԡ�\6��g(x�DL��hK�>�90�,7yN#<�N>�A`S�L���c�L�4\�4�v�,��dQL� m�Mc(O�u#�HLЦ1��ß��v���p&�\qS
��5�"���	Sğ���>U����Iڟ��ɘVGpz���6��5lZ����J)���Т/��k��#�p<yeƧ:+|S�� P���!A�G�@-�i� h��LSFL�,�����f���0�7'�O���b}҃T&d�s��G*�z��ִ�y�'^����-F�*Ūq��a*Ւ�N�<E�f��e�������M��Jʝ;�r�H o�����S���U�\��o��M��?�+�((�a�O��k���gh\�2AU+>����O����a�!c���_�8�S��X>i#��ZhK��M�\��l>}R �GNz�Q�'�'�蟬��e���7�̝9��z!88C՞>1S�P��G�SE��O���0��@����@�#��c���Ivx� �GK�?1��`Q��
�!��e[�$O tFz"H�
3�삑�3'r����)y"�'<b�'��i�`ǟ�>��'x�'��D��wFL}12��0N8���`��#}U�'9q�#L.,OT�[q��#��s��̒a�����7,��)(�ϐ��MK��L�E���>�O��kw�٘k:��en9M������M�4�?�Tn���?�}�'^��]oG�Ș���ad%�ӂ�Y��R���E�
�}��H�VLK&�����Ms2�iX�'L��6�O,�	f�t��'ѻ@�l�:�K�:Ʉ�#s�ݧJ/������������Xw���'��I��@�\,p���l�b�� ۽(��y���AX��7Z�p=A��݇�T��W푃�I:`��H�����v¸q�I��9�j(gԜ�pb�5�	�yF���>x0��O��50*@����O6�o?�ē�?����'��q��ؒ"�(�iˁ�4��'U^���F
�bl��v�<%�1�y"Hq�H�d�<��$e����'�)> h(�`D,RN��҈�;b���'��Y��'�28��ǈ��#>��Ӭ�!T�\7MʹL��C�Ǒs�AA$3Y��x�C�)g�|�Q�	z�����i��D��l"L.������
�8J�l�I%�M3T���"'��${Z��)�Y��\Z�%i�8�	�� �?E�DN�X����Wc:h�!I��x��q�j��ӌ��D�B.�X���6Od˓L�X%"WZ����z��J[282.B4�M��:�t9���&�"�'�"�9�Κ(ՂQ (Y���+UZ>�O�l�EH�T��pk��L����H����gԂ`-�]�E�{�H]��M5��<W�0�@�욿t��a�ą3Rd��'�����#����5ҧ����ڗG�z@��T�d��zԁ����xbf��B/�<��N *��0)U�̹�0<���I>�\}Z�AN�"�h`Y̅�fI.��4�?����?q0'��*'<����?���?�7��2�'�3Q�v��@�I�?϶Y�s&N�G��t�I�4A�h��˗0b>�OL�7"^"#�I"�!��y̌���ٓGG�*R�9vs�-��lĝN}�c>�ӄk��u�Λ[
*`Ǝ� F	�da�mZ���$�%�����?��e��,� a
z��,�e��Z<��'q��rn���p(��Ҥ	/���O�Fz\>��'@���V��x�͚�ͅ��N]��'Vd��@�P�D>���1%A�Z��y��'�B��kW|�々�QWx@h�'���ç�ua��(��	�TG<ܹ�'�-��1%&�Y[�b�"��'�ݻ��(n,�8�!���y�֯+��1�O=4�vЋ�eK�y��߲4�8K�D+(Yܜ�G*��y"MP?b��i���;.�9A���6�y�'*Hr�j��7Ҁ�T���yr�By�y�A
�����yB�Ǆx-:����FrsօA eA��y�A_0)�툒�2n�"Aӧ��y2�9<�^Đ 
�bՀ��߲�y���\c��z��7_o��$�� �y��,YP�ɑm��cR�f�4�yZ>U��V%�h{�M?�y"+5\$�
c|��DF��y��-H�>eJTўn�X�Q��7�y��ʟ5�v�����gH��2�I�y
� �% $�ŘY+0�Y���5�X8	�"Ox�6	Է'�: J�q� ��a"O4� Q�W�9���X��Z3'���`�"O�Ar &��d��#�~V�c"O¼p�G��R򁣕��tSb�Cc"OV��-� t f��T;�鹓"O���CN., \�$i�ښ��"O���m�7w�X�;0��m�8��"Ol	�T$'�f@�3�<^R����"O�0X宗>S���a��!<4�;3"O67�nP[��ťT;V�!��"D�|Yr"��UE�-�"FDg����=D�@jr����`�!U$,i�h�r:�(��o'N1���$䅛h�ͺ֎V��ơ3���7�y��E���k7H�2����,F�M[����5m�#�KV;\�)�禁�g�L�6t��RcZ,;�Ԉ���&�	;���'5	d�2��ڒ[>�(�Յü	�R��		#8�,��K���8͙t&�H�02T�BB�� a�.Z	qл��#U*c���S��M�x���w�i����FF��2���'6��ِ�g���,0k��?i$Dܒ ��b��^�VST P��?	��i��TAݴ���|���+�((�M*ab��1�Б^��|x���4��@���k�'�� U��`���Mp�5�iF� IC�	�3�b9UÊ>O�����?���C�� 3�� v��5s���V�N�r�暉O-g�9G�"�uWL}hň�s�8�8'h8Fz�e��h�:qN��2m�f�@9/؆��e��Sg���D ö*���Ó2�lh��öB�8�+�-+.�+�ǖ�y�0m)P�'�؝��Ӌ"�yR")B����͉��>!$?�6��Q�A#��j��8Q	S�I���'�����z�6��UO�D����i�(��p!��oLax�O�F0��ŗ+A��|a���)b��8�Q$?RL+T �b��\B厝�[śƙ�ܘw	��<���ïTS
ʥ�(?I��D�2�ޜ��	�o����a�Eyr*֏f��x�6.ڧQ��d*U���(O�4�!�JjA
�	�RPSaX"|��P�����Ґ�0<���h��q�E�*�Xqm̠A�܂r$N8G��h`�J�<+�����8�G��B�n�a�Ip^��e�<�O^���35v4I�!i�\� ͫ�l/e�,��?�$��s���'s�5Y*O4H�a�,sL$IP�
Q�9� ���o{�'2"�'��i����=l~�; �ξTun)�e"�ۊĂ�i)be��IQ�B��D���r+��Xh�	�/ ��W�B)2�L�O�
gv#<Q���n�^*��f�d�V'�"���Ӏ��DE	�$��q��� l<<:�Y�$����`�Ój�����+é���$��O�2H�e�/?2���O� �h��p&�T�|�'�a���X�
�s�Z9;8=��6��>�;*h����
+Q0聠 S��Y���k�	4�Xo^?��'� �I�ߍP�]�- ��x���+�H���@x�'m:m�w����F���ԀQ�i�.�aS�����F�n�YQᲟ��M3�v��cW����B�}��,O��V�6�2�$/��a"R��X��1e�x`ҡ�3QO`x� �)ғ;�R�jp��. �& �"� �h��&U�F��� �b�,�0��"?��m��J�)<�b@0��#�)��͆
($���$6�O�%�0F'qώ��a��c��1�d�'Ɔ$�4�+m��츲ϗ!g�m�q×6/�����̌/�l9��܄?lI����ɇE��l�uˇo&���bg͎KȤ���
z�� ��paxB.m��QҷD���nׅHWD�q �	;�-Z�K><Q�E��Mc�cF�A�rX�F�n���r�H�-V�f0��ð0����C�V�hgr����A��	�m���QlZ�K���4$?m��I�f�}��`��%��@ا�½%6�	���U�y�<�C��9B:��K��]^��C��Sx���.�:!�����5���KdJA�~jr�v�P���d\ W��k���Bm2���YS�����a٦_��A�g8e�`IDh�L��$ Xc��&�$6g�ՁP��=���dĈeZ�i"�X-���I˿EN�6]>A*��>��0fL�i
�����-�b=�u&ܥ� ��c�ɕ-�is㉍sa.�
�]?�7�K�D� J���7"I��$���i��i!08r��G&>2�� �A�x���C
�'�~e�L<�K$dft�t��,DG��i�f�$8�A EnV�w���'C$&� x��^rK4(���p��pЌ�D��$-B�T@܁���K��ZD�
R"J	˓ym(�@�,ʂHT�V��Z�A��i̓RҒ`�S��+0Ų���k���oZ(s�Q0��Ud@"��V'�,@֚�e�*]��{b��0,��Ё�E9$���9"�´�N�Ft�pP�ѫH�gZ<m�A�Em�.x	G
7�M�wL��)?X�*$��'kiX������1l���0$�H'S�����I��xl �.#X. Y�'Φ�r���r1&U�A���B��]�J��Y`)�����[�ƙ�ѡ�Od0$�aj]�𘳉y
� �1�4��1F�s"֭wXY�#���n�7hDg�`��y1Op�8���}
�˰l�J<Y�&�]� ��	E)Uc���Ȃ+��	���	az�INn�!�U
�;c!$�� � �M���=�� ��"�F˜0 �Za3�,�`|�6�_�u�i�9vt�ځ`~���a�'�yLa}�J_�[r�u�O^,
F �'/S9@�
	���c+L���ӂ9�"�C��ѓD���q6�uӌA�����]�c���gd����Se�Q�W/����bʿF�n�aT��p�'CT�z���+0����sʼ�s4ň��Q�X�Z�q�;`th@q�#PΦ��T	1�@�3��/lfh%��c�9@��yҪ�;�P䢜�n��T����y��!��h�b��TiQ��}~b]�n'Z1�R�	�O��X�"�&� Q�"FTfz�xxuL�a��M#&�l�Dc��'�J�C ��>0,DxBˈ�a6�1:�4:��@��<�q���� R@\=\2��D��18 �tݱ2ᬁ ��"�ִ�l�1!���>1%�}�9i4`��Mld�@���D�X�Q���4s�	�@NG0�0
���a�(ms�4���'	�����)f�.ݟ�Q�'GWL��@�7f����IJw@��'��ye>O�3��ʆA�&�i��~�\���?7䛶��&?�b0�&�^�O�b=�c�ͷIl�W C�	�S���) mF�"�4�� �Z�b�	�BPf�+�AC/M:�5+@ ���Z�tuiR�Q4/�Qr��8�h{��ч�f��Aaopx�'����|JUe{��4I!�RS�Wֻq	��i�eYvEBH�P�Դ���ʒ^슅�С�mM:�.�01E�V�\��ug�308���[�~�IxV�N�0?)v��C���;B,�_�ȵb��e3`��B���~®	}�ہk�V��6-�	[�뎕�z��̂1��?Ȏ0	s��%
`�(rW~��1&�XR�Q�\��	�Bp���:#҈t#��O�8�����Y�%���(2�r�ifK�1^��V"ʼ ے�Y��H�{E|�sBCq���	�%9�I.V��s7A�/J=)G�P5dP���i�X|BV�Y� � ��น���7D%��!p�
R}2ƚ�PP�`Ů����U&.#��I��6l�bM-�0=7��0��9Ǣ�\TJ�����1sP����wdZ��G��x;��'�ؔ��#�|6������r�4]�S�%i�a}§�/,t���^)qC\���`��fl)w��)�D�5�>���=[�'�|M����-T��,�Dr���o��c#g�5P�(A�4���HO4���A�W`����� m DR�le��R3j0^X$i�F]���ٷ,H1��J��8�7gH�X�F���d�֩�=�D\ ���J1�I����K��禩K ��$7�1�s.�&1�"4� Ꙙ@�hs�j��bl�Ic?2�L=0Uޔ�+��X|f}k$ۥa#��W�]9:�����'��s"(Q�
���B��~t��� g��T�H�E��L��5FNNt�����I�=��L�"dT�0?6���
��S��m�\<I��ط-b6-[�K� �ax��Y�tF�l�a�2��*A����aO��Q�9c�*ɗ,��#>�&j['3�l�q5�'V$���Ӧm�� �*�H��N�4��tJ���&�ē
�L��D׷�%bWM�!B�8��>���)N<��"�J�P���<����3�+d��-�.)�����<�
����ّ��ʋw�|�	f)�Z ��ʄ��=Y���z3�� a{�.�#$����NE0�BVk�<D*��?1s�\3l�xZcu!���7~�4	*4eђ~����^��6�)1,M�(%�"Z����"�?,O�PH�U��N 	AbN�0BvO�P�pmŎ�P��x�bX�'w��	��l��!���i��C��(���Ca��������*}��'�<r�e[��MaU�=�(�p3� �ɩf%V!B��8;�@���iވ,:��	�@����
��sFe���D�R+�=	fG��P��X3�U��,xC�]� ����a�S|P��'
���>�N�*�$�<R0N�3�Иq�����#��S4��I� �@���a'�v����������l\u* R�.
B����G�),OUB�M4l���s���3���������2��e�-A#�h!Q ]U�'���3ԫC< �m�!`:m�
���'N
��ƌ�.���� -�2lW0��N<��	J�%X�ax7�YS[�0��	V�d�BI��b^1h�y�n�K�j}�O��G�־7i�x���Ʒ$fBHD|��W�P^��
F���H�@����%Q[zT	�-� �,��P$lOʀ�i�/��+��Y!!l6�3�(=�Q�֧5�⒉8<�v		�C���n�=�0?Y3�WL�sDKҗ]�FDR�b�:f���Q�<�a�ɨjZmP�č�}�x �䀆�omH��0�W�K�.���`C 1�����Oc~$���
�M�,!A��$/f4򸸒�\%F�\�U�9��'h�8�(��D���V>W�R���}R��!3���3h�*Z0�4�6.���䎙 �TЀ%�ԦI�V��s/�O���'qTi1�`Q���l# ��e����O�6#�$���B@>��D���z�2��3z���rfN����3�O�PP��� 1�sJ��bU(@1�(����q�'�ƀ:���y�Ų� lk�m���)7���ݴv��i>���N7p'����+D��5�CH��F}PfG��*$ȱ���M3��O|	�r�OJ����vRR�kb8O,��$hވ%��K�4�^LI�V�x!���	St�x5-:K��=�&*�k�~My�͘�D�Ps��y�8ϓg_�!U@�/uG��o�"'Vd�����d�R}
� ~��d,RꬤK�%Ŵ�(Yv�G���� ��ZZX�p�ӯ�4���BF�u��AS�l�O�HQEb
˦��O�p����i>5K2Kzf��ac$0s��0�g�h�<�Ǎ�)U(�Ӕ$�
s���YU"�p��RX��u�!Y:UfȤ���T��y���O+
	U��x�QG�R��p?�нi��|����xpċ�)R�{�aԹ�y�G���'Mڀ;�:�8���s���$ruR���F�@��3�͔$�a��E>�Mc��
}���dY0�y�H+&>���SB�>��ч�	�G��P��?u$�Q �H���B�?��>OԐ�B��m�)��b�퐗���NW\�1�[�v���-�$��\)a�	!�(�g=�P�ȓ�΅c�`8�@�7 z<�ȓT�ti��Ǜ�tq����(�\�ȓ-�,Y�'�(Z�|hpu��9!��M��#�rq�*�#�������;���ȓ( d1�ݟ �:��A�	~��x�ȓ�>��L�!���8�ԝVͅ�y*|0j!�����"�՝)�J���A��mHd��w<��Nu�Շ�j�N� 4i� J%�(酩8�ޙ����*��I�]�)9dGJ?���ȓs��xBB�#sz���Â�~����q��커B"v�@� C(l2I��k�:	��d�1 %ceFB0�*e��P BY��ꎝ�6e�V��/G�,H��L��E�f��4�F�z�ɧj^n��ȓW>�I8����vQ��� h��5��Tn�<JF�G�S Pȩ珋55��5�ȓ��q`p�?�2��U$�3qv��ȓG>�\� �LX�4�԰=U�م�#�V���U T  Hf�Ϫb�`�ȓ	]�՘�(���n�#�<4�̘��k�B��̈39y�Y�t��Y'
4�ȓ@�νɖ�#<��Er�M��ȓS����g꞉w�4�� ؠ䪍�ȓ��T�6��u�d����	�X<�ȓ4�$c�A:���)"���p �a��EQl�JףC�a6���,Z�$"�0�ȓp�i�!IZ|F^�R�]\��Wa D�G+?�*\�/�
���ȓ56�%���z��ǂ;�8�ȓ_�T���M�MY(1U�=y���ȓG�ވ33��Ϫ��Q�ܻq>���.��R*	�Cw���M�w:���
?z�8�'��MqTX+qJ͑^�Hl�ȓ#�qp�mZ�6sPs�$L�(Єȓ\ɚ0p�F\
Q�R��卄�Yi�B� a��X���Ga����4�B�I�����ȕL��ՠ���O��B�I+C��B�gB�,zp�����X�B�	�M���#��\�{���iY2�B䉔D���H53I� �c�B䉎|"A�eAFh{��{�H �B䉣|�;��	i���ć<y8�B�	�A�U��B�:��6`ަ7tB�I-X��D������Q4�Ϭ#:B�	!o^���-F�~��9���S�e�*B�	8xy����3��u�@�';B�+�t���ɓ#m�j(!��B��U���c6��I�\	p2hD!:9&C�I�N�x�;1�.�B��e�])!dC�ɤ(@񐣈ʭE;D��pgۃC$6C�I�3_�� d*�B� M��j�=S�*C�ɘ@NԲ�%�&����!��Q}�C�)� N *Si,<%�m�DQ�5�5�a"O�E�'��Mnu��$S�&i�6"O����ڈ"�j���I��V��U��"O:��⥢���J�� ��"O\Yf��7bXP�H�D�����"O�"' �@bM1s
ߚO���"OLm"�&���6
�<�͘1"Ov��QOӡ):P�i�Zk�(z"O���Bo�NY�f�"*%��"O��1�iٴ,��쓤��m��e"OR����z�J��V%��(�"O�Q�!iH�'L,"a%[�n���j�"OhQ4J�/��mxq#L�Ko`U2�"Ov;`F����Ј������"Ok���	?x咃���$�R�xG"O�5Z��C�-�y��JD��	r"OH��3�ـRۺ!c��.��xjB"O�ؒ���N�iB�Ö1v��8�s"O����CJ!s��BD��T�Pٹ4"O4�[f�ۛK"��E�E
'�p��D"O�X�]�A�0�q����hp����"OL��hI#��l���Y{J�g"O�4�����ux#��nQ�m:�"OUp��O64��f+L2pFxYV"O���A���vߐ��iB&!��䉲"Oz�wcBj��Q�����5�6D�,pf�� ��� �,��s���"1�3D��H�C��!;���Q���3F2D���.Isl��h
�%Vm��*D�ؐ���n^F����-+�&Y �(D�+p�C�$!X�)�j .#�i%�(D�\���k�~��q��-uVU�w�'D�<ȣ�ŏ"���p%-�,�F		�)%D�Pu�Q H�����m��S!//D��M�+:�t�W���2��E�.:D� ��bV��q���+�Yy��5D��)��8e
���k�9q��͢Uj4D��XF��mn6Ւ�-�+}B��`R��<Y��?�	h�OJ�+���`@ʝJ\'����'�2d�q�Q�A�E93Ć"Q����{r�'�$���3�TH���Q ��HH
�'��D+%(YG�+��] u�9�'���Q��XE��P�D�]��'������	�A�F�����y��C��Z}Q�-��|�i���y�+Kh2����ă�D���H�9�y���f�py��č��"i4�y��So�%k�o�4�Bu�dmW�yrk��U��p�׶o@"X�vN�.�y�F� T9P�	{_�xb��ׁ�y���r>sO��	&�D�RAP�yH�`���&�&w�(���JM��y��)��&�j�f[&<��a��^�ڱ��bN&9ۦ�X�>�w��}�L���N��T�2���H�c1�@?O~`��ȓ?�P��Uh:
�Z�@�j�9w�d����\2r��r��i��A�d+����{����.Y����Un�y��3"l�Iz�O0D�@(�X9��8k� EzR��32�OfC���B������>5�B�X�B,vB䉋T"��$�D�{���!&ʃ�O͐C��9b� )6��	@d�8Z���8�C�I%u����p�D�X����֢AX@FC�ɀT?0���:�J�����gR�C�)� X����v������B�S�(x	�"O����q����a�*�8$��"OP ���P���@�vB�\��"Or��J�{�$�7CL]HQ�"O����$B>�ƫZ1^Q���"O�]��E&Q�	��߮lFΡ�G"O�p`�:~�0P9s�
j��`�"O<���m�q�(h ��	*��T�@"O�]G@W;+\�q�QlŃ@���"O��Q��G�
�~���{;�<Y"O��pg��1�HH���!!&�聁��`E{��)0 f`�+��^�7�6Й��ԭU!�dA�J�̴
���S�8��e�W�)�!�$�A<DXî�B���q�!�*^�l���~��ƈ�P#!�D�v1XƠ���tE�3r!�͙x4��`�+V�hRC��}�!��,ʮ�J����_�^Y
���&!��j6((.:)v�H{��Gr!�dH;0���K6E��T��#�+�!�@&<
hU�`N�i�`9YE�>�!�3|����ᙳiۖ\�V���6+!��D�Rf�[�d��[5.��a�-;&!�)T��◄�+��=�#��~!�d��}ʒ-��J��Qp.@Rֻw
!�$�#R=2D�#�0z��U(�г!�!��$��ာ�k� 1�-�=$!�DAp����C7i���s��u#!��+C����f���[�D��!��C�B�s��J7\�v@�s�C�q<!�.!d���`�ǀ.�0�	7Nܦr�a|�|bGs(*%���C�TQ������d��&�Y�'X�b�b;0��E�� 5<�Q1�']jԡ�@�}�H��6�&[���OB)�+�
X-�7v��<;�*O�}&���BH 6��t!8A�	�'�n��鋁x�*�Y�N�s2�Z	�'b����� k�0AH�?hbZJ	�'�8��&��NEV٣��_��~}���D9,OUju�נ6�� ҇W� �"Odt��E�$��H� σuY>��"Oܼ+ �_>X3Ji�K �5���/�S�> 00Awi�J�jE�d��_�B������b��&@.�z��ْ&�*C�I+M`��ӈ��U�:$�PLJ�3'NC�I�[�va����[�����'M��-��6O�\c��3���ҠɠE�ⴅ�G��� ݵb�$��E� r\z���4^(����F�m����b~��=��A�,]�Еr��"��~$hنȓ��� �ѝAq��B!�E$_��ȓ7|���)r.��*��7n`F����T�xF���G%�e
E1b���ȓ{Q��҂Ѕ`% ��ȪG1D�E~���97��3w�F)2_U���6�B�ɼ�0�U+5n@�H�h�" gb"<�ϓ�Z���Ȧ]�8zP��+��a8D�t#@d^&�`[��f�<�c�O:D���MS�@fd��������(<D�TI�H!_J�p�'��7!�����;D���a� Q��Y�ւ?�~�I��.D�(�)]4�~��"_�(ej+D���j�N�ҥ��j�.A�ęs��)D�4�@!/*�N���[%I���K3D�� n��a��[��t�E��{^"�4"O��bdP7pN�1��g��ѥ"OnИ����}��p���R`QB�*O�s2������$����R�(�')�`�U�V^|����
�J�Z�'�����?���0� ƼY�ڸx�'�xXµ��I�h�B0�ѣX�m

�'B����T8�L �����{���	�'z�1���#�lhX����	�'�*�P"@�5����e�(�<J�'!X,�1A��͓�ȶ��iI�'4b���:.�� ��T���'#8-9�^8[���H�?��@!
�'����ġ��!�
�� ��
�'z1��H�*�@�%H'<Y��	�'�H��!�W�jhi�� ǒJ�<� 	�'w����i� K-�����D�E��Q�'�l|JV*�"T�H9'� p�'�(��E��;K=8T�6%�s-�XB�'&.e5���K�N�$(�e`�Z�'K,I�S*�.���Gb����
�'�;bMڋI�
`��C�(o�p+
�'�fp��d؅2�D �r#�5gZ��	�'���$�"db��Y�AE�e�� ��'V� �ϕ7�YxA�J22�2E9�'��(�g,�8/68�ȋ�#�|؋�'��Hc����z��,`����<�
�'?�ݪ����k�8�.1�"���ʎ]�<���I隸Q�lL0��|��SS�<�6ß1k r���M8,��Rf�R�<!rm �1P�
*0n|��+Qs�<A0���9�ą{��@�$����r
	l�<aS�h��XJ�B]�)�J�S2�k�<�"��>�L�h�OJ�r�ٚ�a�M�<�2�.���q��C���!�P�<I��ˢB�̘�uL^�X���5mK�<9�� �a�eA:�:��C[�<�3�A<z�
�`C
:(�`!�N�<�1'�,��@7&�*`��LT�<aC��;P���vJժ&B�l�fmV�<I�lߴ}���)d��&un,t ���Q�<y���(B� x �&&���S�K�<y��ЙY�x�I�!U$+\^�X%m\N�<	ΌG~��R/Uu�:*���H�<g#�m#h�X��U�w��Ru��N�<���6���
��Z�:��UQ�<����6i�@��O��X�\}�r�P�<�E�[�{�R|�##�5iH���L�<1�@��<�2H�+���2�K�<i�#h��$����(�@%�D��M�<��NT4�'���hYtpa��L�<����8��	�"a9�Q�IG�<��#�Z,	��e՝[4DM����B�<�ҫ>!gH	ǈ�Q��@c���A�<	�����*#	�SU$M��C�<Qm&6��9{�Ĕ�o���G�Kh�<���U�oi����듉W��D�w�[g�<aĆ?k��Z0OB 7&�ex��g�<9�N�	��LY�BA�%�\�<I&��dgƐ�a̕kw���$m[U�<���U�EH!�d�����P�R�<a!������D��Q��l;!�MG�<1�)٨GB��D��0Lǀl���I�<�6��\@uja�/H�x5[@L�[�<� ��K�Q����J�+U�>h��"O�	#H�Qvr�xT*��\���q�"ON�0�NN�`Y��	K{����"O0�)��*WNT��	B?Bޖ]�"OH�S .<u"�a2tO��q�I{�"OT0��E=l�Qɀ� �S��=��"O�h���['u�,�xi��q���E"Ov�#G*ծ����_*�85�'"On�*p��ju����Lyy�)S�"O��(W?_��ecr�\35��	7"O&Hj�� A��a'dؿIq��q""OfՉ��[%:�"�9��"]Ot��"OdE�w�Iuʾ�)4iI�ބT��"O��ja���@R�$Y��1"OJ��!JA44���9�&�<y��ȫD"O��2v�>�<DʅfM*��0S"O��рH�"U��E��\>c�`�Xc"O��[�k�!���в(M�#��l�$"O����a�&Cg�1�e���|� �xW"OZ�Ո�/Y��̈��4�1T"O��� ݖ<��{D��'� R�"O.q{�,�?B�!pG�&q�:���"O0���'�7'���רK�B�6Af"O�����U"Ǜ$M,��J�"O��P3ę/�vL�S��g"OZ�rGS�@�pѫQ.�D�B"O�բԌ�R0�PMĮL��x�"O�`S�@�6�ztQա�W�ڡ� "OPia��9v�x� /˝!LH%�T"O�HS1`À�>�3m�CZ4)S"O|�@BoX�9s*ty��5G-N��f"O��B#�P�&����Дl)�} �"OR�v�-�
�&����G_�<�ЌG�7�D�@�&�:�:�[Ӏ�p�<1���)h�لGX�R����3�a�<B�Jt�8K���^F�d@VZ�<1'� a����J�3b$e����k�<�8"q���V�m�R�k�<y��N 0ܚ�����qw����.U{�<1�	�2�e���-xAE�P{�<��h�s٪و�'��G�@��Wx�<�f�K�(�`���W�~�����^�<�b)�-l��X�K%T�>���r�<�$HȚjCT�م�O�W�~8�'�p�<9Dm�,5^x$*2�5l���E�l�<�r�O�B˴�Y0��]��Ҧ�UR�<��@�24"� 
�&\����j�I�<1�*�L�n����0�>�81�n�<)B ڒ6Q:��戆$Z㒈�͊v�<1hH�k�c�.P&òQ e Am�<y!�_�|�2 aP�J�Z�6 ���l�<q�,S�:�.�� Ò�K/�ܛ���`�<�P%��"{�#�d!+���q��G�<!�#ֿK���"d!�#^q���Xl�<�f�+]���i�-��W��!f��O�<��Z�5lũ����~k¼�£�M�<D"ǹ�j�Ő�tP�M`
U�<is�,M�ĩ�sd�8]! Il�<�v��~��`�S��6C ���f_g�<y3/rP�^8�*Q3��e�<91��].ڸ+�Q�p.�t�`�`�<1AA&��HI�m����B\�<1b�ޟc�H!�c���%�B�<W�ӓ�z�;#��+A�2�`oHT�<� Z�@���t
�A��M�eL�qRF"O�$q<v>��S V�<�A�w"O�ᢜ� �	�]�4��z�"O���e��6Z8����@�|���"O���e�H�*Ő��D5`=�U"O�d��_B����jI�?�n�i#"O���f�I�=J�x�	ռI��c�"O�
��@�:{VE h�hh)�w"O0�b�AMat8���aڬSI��P"O�X '�ܽN-h�
��m�`D��"ObIfl�3t^�� ��,��)�"O$,�Sa�%Z��h��I�#Ԑ��6"O�M���Z9���X����A�y�e�W3|���\�MV��Q�β�y�!��5���� �u�t�����y��C+m>�Q��6�ͣƫL�yBFF�w�*� �K�#��AU/��ybL@"��t u+�#��� P,��y")IF�t�:`@M&ʴ�*ʽ�y�d��|�CcnƖ,�Tx�c�y���V���G��$:�!�n���y2,̻�Y�fH�3 P��C�ҵ�y�Y�%ӊ��-��	��	�P� 7�y������q�
�(o<: ��/P��y���0�B����G�3�h؇J,�yB�� :�T��C״%&NrwI
�y��sLv��Ι�G�������4�y��1n�8�"�^e�e���y��x���oM5v�fyd��y���|���I��p�6T#�,��yB+Ҿl�r�Νt��m�$*[/�y����� �c͝f��y;$-C��yKF�#񖠱@�Աc���$Ŝ�y"��:7?���U��赈ABA��y2�ǮAVЩ8s%� hh��oӤ�y�曭p�f1:�B]L��x����y� ��T��!��̟R�tZe����y���"ir�q��L�Rĥ��O� �y��U4d�.���(^,N�*�!bd���q�轲t�Qz�}A�H��m��I��I�|�p�H�U���c��1%}�ȓH�1H��S� ��t�Q�[�p�ȓ<����WAلI:Lx��kE����� �4�W���W�
ńQ��fu�ȓ;Ev���*Ћ=
���F�Ec��ȓ9�HpQ�e]�35H��)��Fq�ȓ)�>�
I��A���3e,.^�&��s��M��*��J��a�bfG�y>�$��I�ڰ��愹}�$]#���iuj��ȓ��JQ#9F#(8+��H�C��0$���gĐ�{�d��.I�G�>B��g�l1�עn~xP��Ơ,�\B�I8>6mH����?�$��bj� 3CNB�9}̈́��5�<-���9C�K	O�C�!#��$�� K�i����l+B�Ɉ�*�� ��-�V���hj(B��'-z{�g��9rx�MU$�DB�I	m��Iw��/E�E�"�͛f��C�	&g`,���F[�8�q�����A��C�I�KMl-"uƗ�5J����C];dC�Ir��	X���6H��pke�@'+��C�I7P(�SU�B�f�`���d)pC�&e fT�I|`H<��V�g��B�	��8��d�c�n���A��4�B�)� ��ː`��f�60&�H�@��QU"Ox��wO���~@��燻C�f��d"O�3/��b���І$Щx1�4"Oĉ�&�̈́�^Q�D_4U�L9�"OY���:L��m0CH )M���"O�CB	ܒHW�%��-1/��a�"O��C���>x"�\�#�C%2/z݈�"O�!��BH;|j�H�%T	L�xyP"Oh)KR�M�VGNH�d^��吥"O`� a@�9�"�bS���ԓ�"O�g���-J���֤�:o�4��"O�5p&�Q�[��U#�����F"O4hbA�2e�Pq��#gz25)�"O��H��;ew.�k��[��l�@�"Ob���!@�%���B�O����"O<�8��ߚk*�M����C�m�p"O���` @���!��B<�ə�"O@�{�Gz_X��/
,`,�}�b"O�s� ��<uk�-�9'�(�"O���9��CRL^�t�p�#"O�R��(}  �v��i��Y�"O @j���7>ri!��L ��sd"O�1�!�4Z�tx�	�F�t�1�"O��:vWm����������%"O��lD�G(�l���ԁ��(�"O�a`��B����'$J��;�"OT=S �%0k3��0��"O8�S���g��������Z3�"O.���f"���\�����w"O���B-'��R��/�ِ"O�t��G��W�(PcQ�L�	�hI{f"O��/A}�@=;WE�H��8"&"O������(��TZ�+Ҧ$�ک�"O>�@qfh����
W=N>�z "O�$&��8p7�@Y�k�MAH��C"O��1a�E���Q�	�<)0�@@'"O�xb��St:B7���0��C�"O��'�1m�`hQ�f�B�����"OZHc�NI6>�D�yc��0Θ@�g"Oj�@R)QR�Z a���:���H�"OHA@��w���`�I�+u����W"O<��V�1�rGnK�EB%�!"O$��p%`���d����0"O����j�4>�5����{�Vl��"Oi牂C�T�5ɟ�y�
!`�"O8 c�މh�
�3��BD�6�b"O`d��W'T\�����&~��ͻ�"Or������I:�*�1��\q�"O�"U�SN ��a��Ѻc�L�"O�I3Do�*�y�Ad��Q"O��cr'N�8��� �NuL���y��@�����ro���{�B��yR�L
7!���S�ތ&� �� ����y�S�C���i��	Ń��y��{�j��Ŗ5x�2TJ=�yJј\�.�˞8	S^�A�LS"�y�-Fa�<��1���tj�ի���$�y�N �A��I)r�ÚX���yE�@�y�ƳO�-f���r$kKH�((3�'2�5�1��@�T�s�j�%G����'��(�#KƐd%�шtϜ*@���'Itp�GGY5&��Bc�2����']�er�j_
�\���B
,O͢	�'U��P�EN�<�xh�r�Y�;���b��� �� ��Ɖ:�� t�[��� �@"OD}y�h3x�hh�+���T%��"Ol�qe�^���i6�?I��q�"O.1P��ސah�|�(�@D"O�D���.@�Z	�f��{�p�q�"OBI�F��m�(��̅�6��!�"O��)0e�c���hת��G��� "O�XJ6IۢM�0�r���^�9�"O�3eD�<��:a�"n��|��"O�������,9 g��4(�"O��#���<9#�]�F���2c"O���n�E��	ሏk5^l�"O����	:}��p1�,.�XHR"O$L
��),ƾ��qF��6�1"Ot!�lǝ?����a�S%�h�XV"OfԛC�SṔ���`�}b"Od(9��Ao��A���ځ��"O�L� �'�H�J�:M�\i��"O<�07nÛ ?,��ޜUi\�%"OD�'��4V~ڤ�&S��M�V"O؍���I%o�H`g@L5_�[ң"O����60���6P)T��ae"O:8�@�0���󫊶6[	�"O��13�ԧÈ�a�h�o�r�"D"O:p����K�*$A'�F5���H�"O��D�AB��� �/_�T10"O��;v���=R�X�OR�i�"OQ� �՜1`h���,ůwN+�"OZ5*5j�*[��Ahu�	�L1�C�"OHA�5",:�5:��Z-֐��"O@!�u�1��pQeߍ��s�"O��!�L��+�f���c�+1���"O�Q01�N�<҂X�9K�LMy�"O� �`�W��A�M^�>܆ax3"O��q"��)V�:'^�4y���R"Od�P�k_,rrpY�dM|�M�f"O��	nU�;\�Xh�CI/F@"O  ��ԧ;�\�EƏX��18"O��sسOe䝳�$΋!��� 5"O���pѕ���Q���%J�ẍ"O�M����12"�X9�HZ)����"O��`$P7#�ܸ#�0��Q�"OT���,fIč��G�q�@8J�"O�9%��	�x�S&fԍ_~@p�A"O���d�	�OU&d�c���OӺ�KQ"O�Z%�>v�D1�s��`��s"Oڼ��kS�u I��L�b���9�"O�9"˕XW�R�J�w�r��Q"O�1Ӆ�^�,FBY���k�2�"O��8T� d��h�lY�����"O����P�z%Q���;A~>4��"OΕjUf �5L�E)�&kF`�2$"O����7O��I�mM�s(���"O�x�g +d�*T���J61�AS`"O�a�V$Ϳ]yj�r�B�7
Qc�"O �����q�8Y�&�6<�b�B�"O���C��|���8kN��\c�"O�b���m�|;�Ȥ2:�I�&"O$�k� X�
%��o40<`�"O��f`�oDe��05�"%�"O<��=:޲�%��o�V�XE"O�Q�r��=16
�z6�On&�b�"O�|���m9�[6�޴P�hH�"O��2D�QNT�[��69AW"O� ���@�}<8rbe�t�
u"O��2WM6.z	�B���!�"O:M��Jխ4\К��˛y�L���"O
X�B��?ai��x��R�`�h�"O���ƨW^�,��B�$4s�#�"O*=Rk�$l��S�Е\Q,�is"O��,)�zM���Y*:ق���J��yb!ܞ42���v,�4evf�WB�y�C��`Uz +�Y��TB@�M�y"']�C��!(��%R"K�:}5Nl�ȓf^�l��A�i���j��5C�����O\❑C��'f׾8��J�|����C���c`*�+r����H�u�>؆ȓV�j�ɇi�T�Ɓ��k¡D����8v���`�R��y1ZB���i��h0��� #�r� �+^؜���\��'@�8v��?\7�|�ȓ(�$�E�&z�p㕏��O�(��ȓ)��Qa4@�#�6k5@
;<LԐ��Nz(	qA# �>QH!��޶0-�M��$�YR��;_ʝ�v �p6x(�ȓy���Ӏ�W�.DH�2����ȓiq|���I�=����'�O=�d�ȓ즹总W�"���X5KM�ȓ��r3P�l���EnV��T�ȓ4�V=����5_~����Ռf�*���l#�x�e��+iT�b.Ȱ,���yh8Q�1NI�	-��S�%/��܅ȓ)����c4 2�p�roĻDF����_�P����1~)�5H��,��ȓϮ�2���#n�Bբ_	�L��[|)A�M�)(�)۱� ^Ē �ȓR����i�(w"�����J�!?B��
bֱ9�MUqdL�Ԣ��(�Ԇ�o�|@#$nB8��\�Ѥ�؄Іȓf���Xs�
�fG��{�E��`�I��+B���1��)X`�0S�хdri��~�M8��9)�	Si�8Nt`��ȓhrz�� �^�?���Z�"�6=E��ȓc��ݛ���%	��9��H��=D	�� ���i�C@<Px#*Y�R(��ȓW��aΌ'�B���	$���2�Dq�!��`X��&��X��ć�tA�ݙ�K�
f���Ge	�l�|�ȓ(#���䣇1.�le�P'Ǘ�2@��m���K���4yEcQ����ĆȓjR��5E>��MHE(Pp\��e���C���d�e��m��5�\��ȓ
d�
#opz��r�~�x!�ȓk��EN"P�-�!�b��i��$s�)@�J9qǆ8����<<���'����$ΟDӔ��OR)�~��hz-s�� �ob\8��!<P�ȓ'Wx��3&U�.M���T8\d��ȓEY��Z&��J�Z�CK��0��M�ȓT|�8sK�yܖds�%�(�8�ȓN`�Xb�b��,�D5A�0	�ȓ��̚d㓟R�,��5'��B`�y�ȓ-0n�1b�]:8��I�3FS��$]�ȓ|��!!F���	Sp�� ��4����B4�pؑ�B�L@<0�+On��ȓ2��s�H�@(�yyFL%7�V�ȓ2�Q�!'
��Y7*ܦd�u�����c�;�4=9ƙ]�y��S�? *�� N�]6�t�1��XdD�i#"O�4x�.Ap��!��G,{T�p�0"OB� ,�Z�Z1�]�Nr�E3C"O�g��!�|��$$�E�q�"O@���/��l�|��wA���Q3"O� k1d�gC��������t*�"Oҭ�tg�(1g�!I�LZ:&vڹq�"OTA"���*��ȃՁL>;[Й)�"O����,6r���J�On��@"O�1�þ �z�q��X�q�ba��"OV�I�d$d.V���I�~E42u"Oh�ʸq>��@+ʱ=H!�"O8Hjb��"`��Ū�jIh�V���"O%P%ͤs�|ZS*�4��$9f"OHyäҞ(�&��S�6�V93�"O��3&�d>P[�l�,tV8���"Ov�c��rΚAQ���-1:���T"Ori��e˝j<�L�¬�J
��y�"OJ�rClQ�\s:�'aw����"Ob��V�B;k�L�go_�+�Ll�t"OV@�GIݑJ��q�NJ�ZВ1"O������?4�@FMK�!�ލZ�"O� �Ň�T��rftm~�A�"O��`�j��E��๡�?�0�6"O��`s땁E�^��]�|B�eK�"Oy�/ǓxJج���ʨ �F%	�"O�)$�B7o*tM�Q&�+N�HpA"OD���ˆS���C������"O�4 ���'\>a f��3�$%�"O�@"�HL;a���u⎍;���Q�"O�xC�OGya^��R�M�!�*(��"O��x0O:A�pp'�@�,5�""OjQ�M@i6�R��
r�ԹH`"O�L;�X��=�m�A�8�K!"O�i3�8yP�}� L�(ډ 0"O,U)�%ئ4�f}���d�,�r"O*�@��$bDΘ��� Q�ؘ"O���H�n\zscA\�A�"O����E�7u��J��$��i��"O��I���4�6m�CAݹ#����"O���c	�>4,�Y�A�	)?lz��%"ODY�� ]I�j���A\9�@"O�QBЉ	}K�0�n��!����"O:�(�C�|È�P�L�]���a"Oƀ��k��^����L"�ġ�"O�����P$^PRTpD�G�dQY�"O�`jefH5���/]��vJw"O��$�҈[�J� ��*��Ar�"O�I�)�E'*����(+Ԗ� "OL��D�7[ĝx�߸L���"�"OD�AS*�0g��� (U�d���"O�m�6]���h gFє#DF�{�"O� [���({�:��0lJQ��8�F"O�T���D��H%h��;����"O��ٕ]Z�h@�#�V�DzR�""OȌ2�!(�,")�9`
���"Oڤ#��!7�~���b����"O��2���=��-���2h/y�w"O����� ��8s�E�Jbh� "O~�����:I
a�ҮWU�8{�"O��&���T�r|I�KM)�q7"O0�G`Cb��S�	��>ؤt��"O��:�. �$��㇆N\�-��'�,1��/}�J	�����|	��� �.J����'�n$���"O���b����$����"FTy�"Odh��J%/ţW��7S�D���"O�l����\��W�/�XP9�"O"�`�m�4��h��-P�-j>���"OB}z�&�%�V- F�ʬlN��
�"O����]j^ 0�U�t�h0�"O
��.�D�p�1��C'C�t��q"O�Cǀ��v����G�V�T��h�"Oj4���ۥT��dq.ظ��UaT"O��6$���<�z�,�(��\ "OH�ql�+���`�1L����r"O�@�6�_�b�õ��%{�y�"O��7Â%pm�����Lh���3"O*�XG+�QW�\�� \�Q8�z'"O��e�ԟ`���qOH���qY"O(|IU��
w�ʡ.E�S�Ba��"O�ys6`Y�%�8�'��?K��`�"O����������-�
�x�RA"Ol���@ �m���V  ܼ���"O ��B�Ґ=(Ȭz�`��+Q"O`A�Ѭo���쀭[�0@"OH�1�
�6�X�4;�f9Ҁ"O��:gV�{�V8��D�����"O��2��Dtc�+Ѕ��5 ���"OZ�Qs��Em�������e�E;�"O��)0�L	��(�����j�"O*���oYO?Q3�H^�х"O�C�Ȁ$Z��b���&	�rq�3"O�����?^�n�b�V��1�"Op�j��֗w�2��An��%����U"O��S�p� ��E����yңǍ �0(*r�� ��1�)^��y���2S r��"���y�D��t�Z#�y����W08� ��\�NA�0-�yrb+?��1��T%y\�c�6�yB,�A���jL N�pH���y�k�"R8��Z�>��9i`ń	�yB�ښ?�<ܺCʃ*7���g,�1�y"C�����eŕ�z[���#hƒ�y��4�u��,j��|��M��y��΋li�5[&�۲l!�%��S#�y2.�:��Aڂ�ב`$��F�yM@t�r��c�Q� �z�C��yBj_;r�aK��&R�np��o۵�y�-[�s �P ��F)�@xb���yB�J�}B��U�S��6 B'J��y�/�"��0W�ݜ_�aZg��y�$�&sqBᣳ�̆+(�X���N6�y�+>����w�A�%^��@d �y�*����);�n
*f �\��j(�y���u������G�v�ƈ!�y��H�:9�m�-�4@�P��C^��y��³C�\��n��>r0 g@H�y�ꂳ.�X,"��,��a�^
�yK�q±�7�ϷrZp��&H�+�yR��:`J��k�J4�䚐�y��ǣ54����F��[/�h�G��k�<���A���!�\�^�s��x�<��'��([vʙ+��t�a��w�<�d�T�wtH��p��i2����W�<1gl��Ly�B��4������Z�<i�鄢(=N�($��6o�E���T�<Y���#�rYr5��#��L�#�Wi�<� V-�%��3,��-Y�,���"O�k�X�(1��)�O9[�D��"O �%퐘' 8th�ې1�,*�"O�!б"���rt��"O|�C$I�H��T8g��em��@�"ORt #Ș.@��8����"��)��"O��8�&�)T�eZ2KΝg�j���"O�5�e� rz	Y6�� �&�6"O(�J%NhOn�@TeT0cD��3"OP��C�uը�壊���c"O��A��c�)[D�4B���"O�Sef
�0�B����R��9S"O�i��ǻP3���o�l"��k�"OZ�:��X"Q\&`"�oۆ##� �B"O��ó ��n���嫌��l��"Ob`2
ɘ�Rdz�DF�q$"O��Ps%�!��`Z��X�*�0"O"5���P�=Y�X�F �H" ���"O �f䞾	�&@�� &�
�"O��"��<+�<LrQ�����P"O�XPD�D�4��}r!�!�>H2"O�@�1*U��)#��"s���Y�"O����#q�.Q�7x��ٓ"O�)2ө��e0�4Z�A, �Tht"O� �Q%�9���*���&u��r"OrX��AX�Vݢ�/�U]@��"O�P�UJ�60dT5��fF
=��"O`];�@�!ň��#��o�xEP"OhlKZj��E��	"O�-��A1�B !��!�T(��"O2�a���$M���];b�r�P1"ONU�I�2w� �����T*#"OZ���k%-�� #��C*]a�6"O`��F�9<�|��RJ��?NL��V"O8$�&�U]8DK�	�C6t�Q�"O��ҩ���R��M (� "OԜ��5>.�E;�i /\2v���"OT�b6G@": ��H��j���R
�'����1oJ=��aRu���^�t�	�'�J�`v��o~M�'V�^M�0	�'�f��$D�+�©��.Ι[T���'t
�f�D��PP�t��-Q:��3�'�~X��#]�(�Df���d��'��Ԑb�Ҋ'�����	�>)\ ��'�V�j�m�{�4`F��!:��UC�'�q*�m�`v��av���:�ꬢ�'�xA$� �{��a3��+(�*d"�'9n��t&�����](�b�R	�'=|� ��hX�HZv�N���'+N���W T8�b`�?=�~tK	�'�������8{�.A�&H��8J��'��k��K�*����ܙF�ģ�'X:���@��l鄪ʦc\���'Ѵ}�Pb��L���$�Wv6l+
�'�Z=
@bX�Q�z0 �MO�W+d�	�'���x�	5d�8����.��t�<�S�9�9X��L֘В�UR�<�Afzٻ�K�G ЃSX�<A��O�([:�
@gӼ���� c[�<�U�ل>�,�i ځgx �R��Z�<yQ�W�J�H��"��<ɕ�M�<y %�	-]������#baHa�⌙`�<	 m�+&<n�K��L�A7숪w�T�<�FH�w��=s�h���.�)g�Jw�<� ���w!G��b����(2���"Oj��2˒�Ad8��Q#�38"�}��"OJ���阄T�`Ƞ�c�D��"O@	���G�jaR�S
�/4슑"O�YZ�* �m��h�X�V$�#"O��Kc䆌DG� 
���g���3�"O����G�0w�|�����7Q�d	�"O�)�BdQ"u�au	�S70ա�"O\�!#��m�N��I9y;v8��"O��j �"YY����g����� "O�ؠ�;Y��b��H���Z��-D�0!F��1��@c��9|`�ը�g*D����*d�h�EK�(ڊ-B(D�(��)ȖT����%�"V��6J%D�h1EdM�*�PLS"�/�X��#D�8!�@ҏ�@ Ӏ"�"RD����!D�܃���hR@��#�_8T�Kb-?D����i[�,�
1{��R4���*s<D�����R�'�N��HBQ� �[/!��6B� ��J�,	��X��.g!�d�=!�2ȑ� 0Z̎�9��U�gr!�Ǉv,riT�;B�6����$b!�$�VI4k�/\؈rWNM�R!���U[x�1e��v(6�!�-]�j�!�d
�lt	�#��?
bȊ���F}!�dg�`�T�*��ăߟ{!��6m�h�Ib�'@�"��I	y`!򄃺T^���	�7؂ik��_�fI!�D�r�r%o�RĒ�A�<!�d�W���t�U�N&:�
��\�$!�DC�v�P)1b������w��:t!�DQ6i�%�'oB� �4i�t�S!�!�Dޜm�ɨ!Ʌ�D�P	��,E��!�D�3��I�NJ�&�kE�?�!�d�)s���L�g��1�1�M�!�$�J^
�S`�)w�n�F$��!��4k�U�S��5����3�N1<�!�Ęng ��e��&#r�ad�V {�!�Ɯ��)�����mÖ.�!��ς#d%I7��5�E2���|�!�d^=w�Q ���M�b x�ϓr�!�Z�}�`����ٶ��EH���al!�\/�0�KD���E�1�4a!�dג'��!���K|b�m���\J!��!���Q4��rF%:H�8:!��>j��
mŽ��ȓ̘!j/!�DT5;�q��b�%�ޘ�u+V`$!�dI6��]pgZ1�M�F�C8!�d^��ڂi�Kݠ�AB�:G!�DJ�:r��JI���	0��$7�!�D�KA�$`M�P�B�O��U�!򄓗")褺A��/��S@� U�!�$� X����κ(��1�J�!�D�6fv61*���h���yse�5-�!�����%��.��p��9S�q�!�$�Q�e�>�$��UK<p�!�dݓ~�d0S`
�2�hXSwg�7+�!�ğ!E$}{F��;���arŘ �!�d�E�����ؼ[e�Ċa�D
Z�!�d�(y�<�q��'U4Ii��kZ!��3r-���b�T�q��鏕f!�W� �5J�6dQxa��SU!�d��;��`��cZ�I��X@�
F!��Ӓ"ᛗ�\��� & �v2!�� �)�E��dTb�Z!)���cS"OR� Qc�>u��(� �(\&0W"Ob���)ٶ�$nG�6Z��(�"O��8�E)l̠��J�
Q$�j�"O��c�F�%TY^	 ӈ�?��7"OD�!��N:
B�x FϮ98&|)w"O
u�`�	*M2Da�_+*.���"O����Nce3�Ņ�(��y�"O�Da��_gAnP �G�w�H�Ɂ"O�T7���,�C���cl(0"OF�b�(��s����ǭ�� u�๶"O����׼\k.��@�K�Z�Xu"O�e
���D�U�V+���lP�7"O���t��<�^	�ʃ
;�1i5"OD�
�J-4�~��b�T5�p!"O��8�ɩV�<s��+1��ӑ"OJԳg�X:uK�H�N�p�"O@ء&�ܚh���P0�*U(:��"OН ㍵GY����K�k!N�Y�"OH�H��Ț9;����'��v岅�"O��Q��ٻp'!��'�YӒtZ�"O(	D�I���SB.��rC"O`J���6j�k�d�'d�P�"Ot 	#��+#G�2P-�&�� �b"OҸ�D΀h�6XB�7�4ك�"Oh���Ƙ7�L�p�*[�uJ�H�P"O����ǀX�u;E�I�
@j80 "O-X�Ê�>�M*�/	'�s"OVdۅ��7ض��f��-��R�"OdYa#��Y9^Qٰ���k��(��"O��*�v����pD�,&"O�Y+mq'p�#�V�!;�a�"O��( *_!Y�%�� �1@���"O:���m���y���N�^�t��"O�L�D�_=�9�WM��9�
���"Oj��gXo��2e!R�,�\5Q�"O��2�,xJ�h6� �LD�3"O	+�ȗ{~���1�(��ƫ,D�H��&��O& AR`���
�"�+D�ȣ�N֐<5b��4�
3.���h'D�|�r�(O!�u����m�� R�&D��{����?��y�#�l ����-#D�����]���RQ�"{�-y0�"D������
�@�����-/�R�yW� D���C+�r�ZH��Wa�B��Eo=D��a�)a���/Բ$^(���;D�px`�N�{�P���ԭ\e�ءAo%D�TU�>��5K�
]�h����0D��ZԧӃm}؝�B��	���ō*D����%�(a��@w�Yt=����&*D�HX��J:nv��]�|S~#O-D��3Ϟ�X�!%�ݷ;m��%*D�ܠ,��r�d�@�ϕ^S��'D��w!�1X�C�JSj�J�O%D��*�/^�A��0��1v�ʐK" D���G
�(9N��2Cܝ*6�x�S�<D�@�b��r�ܔq�O��M��<q!�:D���d�1ip�B�kϱR�����:D���Q���*�\��*Mj�ْ�7D���c�߅2�`m�/�	Tv�8�c6D��y"�*xˎ��%�G��lX��m4D�  �m_�6e$��D!v�JL��3D��ԪF�@t�EZW�B� ��,� 3D�����X�1��Q��oA�F��z��1D�� 6� ��Ō ��f	w>H}�4"O�@0�I�?}�T�c&�ԟ*~x�"Oj|�u�ǔ ��]��߽+���"O�չ�\�0.���C��{$"O�u��Ц
s6̘�J,_�$!"OD���GS>�����G�E�`"O��5�A�qo�{�g�� �	��"O�-80ƉUs �2��C3!i�U�@"O�!*�+ȁ	��9K���"I��af"O���%ʚ,x��Q����uS-�"O���L�!ה��%�+_>�I�"Ox��$�F?2(~�9+W�y+�IR�"O����N�h���>U�I`"O����3df�\q"�c�b�"O�X�g�ܴ]o���#�ؚ@K�I��"OjIp���7g�����ȃ�U\j�s�"O����%ɯ|{r�������A"OB�J%.�5n��#)��XM�"Oz�yS���1�t��h�8p�>y�"O:z�ID/"�j��-��X�*��yb�W4eB�I��`ٴ�x@a���yb ۩,0��C��Y {�N�8��F�yB�_�P�޼)��p�&Ă��֝�y2h�-gM�h���«`"O%�yB�."$��k�I:j������y�O�2x�pt�$��a�S�Dӟ�y��0R���Y�&Ί��&#D�`�$eӇB��)���f9�����$D��0b�~0����7d�dd뀤=D��Fm�2Ԍ�ҳ�YK�1�s�)D���U�٦)�j��f�̯s���p�(D� �A�E������#OV��%D��LTr�F�� �hw.��g&$D�8�tLÙ;�JɁ�,��0F6D�Qc: sxI�s�g��L�`�2D�x�� �&��\�b�7fr�ȱ�,D�3�b�
3��8�P��  �d��w�4D�, �цV%����с�Ir`�&D�"����e���t�1a�D%D���d$�?�]�&l�:f��(Z��-D����+�\������(���+D�Ȫ"kC�B�:h�$�ת1�X�&�+D����*M!x���Q�b��C@��<D����F�.ZTh9v,�7,����n'D�`+�½���(�&�/�޽�G$D�4�o����Ꙓ?�]K�#D���ǀ�uN�A�I��Bk�U� �-D��2qk��G�`��ҍ�&�z+��,D����߀<j�}{�l���C�'D���k˻z*�a���|,.}�WL7D�(Ӵ�A(��'웗;�h��@7D�x#׌�3��-A�Z3|�XC��6D���g�0>������I�\��1D�t�E@]Ap����.s�:D��@��-�Z�"똋+Nlt�N:D��K0�]�6V0����Y�@8�G�9D�T�c,V�^��P8wGɢj��a�7D��8s��?08;U��t,�܃p"9D�D�B�M;J�B�e�"�� c7D��ѧB <�6t9iF�I��5 �N7D� B�L��W��q����=x^��k�D+D�@���=$8RA+���'}f�i�*D��
�$��H�Ftက�C&�g�,D��Z3��iV��Sfn\�Ĩ��J+D�� �Jԉ�&`��c�M�?Z�miQ"O�����Tl� y8È�G� M2�"O:��	�I �d�rƞ�s��a�"O0y�r�͌m4��D��>|�dx�$"O&�:1�2S�`�A%J7�q9�"O�%��O�rV��䋃9ږʡ"O�Y�e`�Un ���I�rXH�"O�����)LK�H1ꚝ4����g"O�hP��N�vԛG�
bپ� �"O�`���11�*UHA��^� E�"O�i	M�X�yZ��̘^��(S�"O�*t�_�BZRy[��"m �f"ODT��#�� i�dC���Lk��"O^���h�U��y�DC�!PK�"O���Ɯ�I�⣬ЖEj�"O����,,�����"Ź&���R"O�b���<M�Q٢�H���c"O|� �֨/I��ҏ���z�x@"Oơjw*G1ss���nF�5�ҝ� "O��@7�]�?�~0��h�(P����Q"O�����n<}�c�D�f�x�0B"O��	 �թ<��܂�+@�*���y�"O9�ъ��/�< ��)�$6���
q"OٰC �>��x6��;k𸂒"O�u�aMȀ#c�L�f��2FS��zg"O����O2B��xb�K��#"0n"OJ�Xu ?H����j�&>��au"Ol�����`Z�0[ר��'8F�p"O�<��a)OsF�b�
- �R6"O���u-<Mc��&+��#�"OP)#aO���)�3`�:٫�"O�L�U��a�x���r��K�"OV���t��Y�/QD�¡��"O���k5S��Qω�>���"O\\��'�0�"��R�Ԇ;�e�U"O�e�5J\H� 
�r,��B�"OR�a����Q�R�&K�9�"O����E�0f��N	�>��t@�"OD��e^��(��o������"O��r䌕�"���Q�Y�oJ�U�7"O�x@7�S�;�DM�M�,A�@��"O<�;VK�&��X#��C4a�"O�}R�+M%N��(���%٠"O*Y��ȅ�@��=�� 8%4Tz"OI"��4�&����60!b��v"O��Y1&:B����"�G���y�"O$�;��ȖǦL;A�!�<8"OZ�{0�ٕ^~����<!�Z�"Oh��R ��)<RL�'�L���: "O��J�
��~V��`,$ۚxK�"O)2��	�b�t)2
�.�<�؄"O�l��n�d�sJ^;qL��P"OȴAd�����j�/K��{"Of���W8>�	ۅ`��l�!"Oy!�%z*�!����<�q�"O.����x����͒�Qqr�"OԙAs#A|@���<Tx�u�g"O�I��& v_�ax�EJ�n�!�"O�%rç͜_K�� v�άly���U"O~)g�����StC�.zBޝI1"O��k	�
Ab�)� �2c9b���"O�8��CP���}ڇ�%,
ܫ�"Or�oӾ*DX{� UA�z!"OJa�deˁZt��E��>μ�r"O� �m��$���@���g!6�u"OhQ�KԚ(�lqѣ�&]v!K�"O� 1�%#�b-4����9�`"O(mё�@�/�QB,<$�L�d"O:�(!&��_�$�`��-L:u�"O,l{WM�Ti��� ��p"O�lY�*Q6o�f��"�� �l��G"O @��E�#�B��P�֥8t����"O���MɰT>��h Ck�e�C"O�����É^�p��2�N^W�m�"O�iV�"!�2�)�Sz=�f"O�Mc�eY��0%;�G�1_9�:�"On8�E!�q"�F�X����"O~,E BO��e�L�y�)�"Ovᰩ�1t$��*w��a֔[1"O m(�aI�m��H%��/�<|
6"O*y	��T�t�����l�.}�f"Of��eU~e���%b����V"OLٛ֣W�ڡ�$CS4���H "O8!�C����r�lZ@� �B�"O���� WY�p����2}x�U"O@��L�/3L��3 �3`X��1�"O)[�e��%��,�pO��I�x�"O8	��֥8���q*0Љ�"O^l�`��,s��:u*�6vH9�	�' ����&a\@�j���/�Ĉ!
�'�(假AY���P����7�U��'y�ฆ�Љ��ŨU	S9&�@��'4�t����]����\�h��ܑ�'�J��q�O�?�q�
h�6���'��I�F�ȍCϺ��N�e!L���'a�DJfh֟5}�,��%G�Wxn4��'�08� ,@��Ĕ9���TxQX�'�؁�r�Pk�Tx��m�O.���'B��9�-�|����"U�5�|u��'���L�O�x`�%N�3�:]c�'V�m�0ߚ �#R>5�,8�' tubc\�>E�z�#̻IϦ�C�'w���G �}�]8��ւ=w�$�	�'�dꐈɟL�[��$/,��'=�4x&%��ݳ��ЊT�T��'� ���F�*ṱ���"�
�'5`Ȱ�B�+x�V�;���f#���FO���nc��0k�5b`��ϑ�yB�[�m/��&��<,���+P*�y2�W.x�A�Tڲ Հ���dυ�yb�:n�����*\Jx�nު�yRNɟ����Y!��Y���yrU:5�,{c�E��4eR1	�#�ē�hO��8iƭ�|T�h5�[-XT�"On!�� p�ĥ��G \\h���)�S�'U&&�C��r��Db�(łS�.��ȓz4�zG��+-��i5ʈ6/q&Y�<a�4Q$�y��;V<ý'[�0���ߩ�yҩZ�t-i6�̕�t� �%X���?{���"�Ȋl��h�AX���TF��	��D!IS�
 W �¸�B�I�iZ��{�+�9y�dh�gC�#}�~➌��I�A�0�p��X�.AaL�1$�ZB�I�(���2�JR��-q0^�ѵ"O�$Ѓ�:N�bt�.O�+/��!�"O.�ɐ%��J
u�rN�IE��iU"O���#d}����*�҅��"O�����z��ѐa�Q4F$�"O� ��@ G�h������ �`+�"Oީa��gn� ��T���b"O,�0Rj��ײ�1Ǭ_=�<����D0|O�K"��'p���!l� }Ձ2"O���V��&`�RDP"kI�0v|�S�"O�\x7��!J����aJ�1`,�ˀ"Ox@ʥ�N�$,�3u��:��pC�"O���S����:Ї��#F�X�"O�u�s�у1��%��MH�L��b�"Op��j��Sx�lk�KV7p��X�"O�)(�➨S� ��E�͵�.�Bg�$5�ŞPF����- 2U� �/W�d��C��c|��M7�^PR�h*Ud`B䉴Rk��hFΪ24��"ƈ4RB�I">c
�#CE71M��A��m�B�	�6R�	�b�&r�b�A"��DC�	G?R���Y�~�!��$JUC�	� ��a�N�7`���)Έ^��B�	�|�8��h�P#fL����"O�|�2$ �j)���D�1͞�	7"O�	3�aÈ >�0A�p�T���"O�lGFѳv���s��=#�lQP�x"�'A�q3�j"d��eS���2~���
�'>Τ[7fսd%L��@Ø�{ݨ��	�'�z����r�t�喟�਄ȓ`g�mP�fS�X�F5g��n��Ɇ����2�M��n�j��R���[kX���,̖��A��x�d��5�ȓY�xh�"]����f6l���ȓVNr���16p|�Gg�5(yZ �ȓ� A�%�p�J�$Η1ad(�����Jdgѩ 'v��CP�h��]�L�C%>/܌Miք�!)���'�Ԅ�I0URI�����i cF'er���<�v�k��B�)+ I��aޢ5$���Y��=�c�&�©�6C���%�ԇ�	
}B�% ��!�񹅯� e��C�:*�)e �	L0NU��C�)|`�B䉉D��BGL(C#��1P@��C�B�	�u\�ܘ5�]�L6d�5�\,$�C�I�afx酥��7L`�
��'!ӸC�ɪi3)�Ǝ߈|�\x��G��C�	$�*��f
Y9n�$L�D
��*��C�4m������.�6�CN=I�B�	C�V�a'#ϑ:�4�h4�4`��B�I�zV�H�e` �+q<A`$ጝ|s�B�!w2qR�O!w_]��eL�aLC��>L@D��`���"AÉ'iC�	�?����퍅Z��{��; C�0V 6,_=��dш��6�*���r��(|�js��Mk�6���*D�{�* ,u*,!���<�BL���*D���nͽk��E�G��j�Jl�fA<D��� ꜊B~|��6�Ǿ8^�×+7D���F�K^�X3ωc 김�6�O��O���/�� �ZxXu�ѐP��mA�
O�7�HW ���؏?���0�ļ^�!��?r~8p�d�G�i���*4폛�!��U��!Hg� b�@+���H�!�=���i�,��m+~5ؖdÊU�!�ڝ��a�7��_+t�AЭh��	Fx��@X�;�� PfG±wr�HwC=D�d�taҬK���0�K:d,B$c6D��Sw��t��=��L	�@-F�3�3D�� ����66���ӡ�n�]u"O���D`��������?]��@�"O �3��X�r�@2�L�tCJ����DD{��)�m�`\�d�x�0S d��U�!�I�z}��u"_<!5�I�IШ	!���4^�b�b���0_(RLp�c�!�Ya
���UDxsa��DI!�DL
I�=8�`��Cܾx�cnD�S��y�g!�I�L��t�b�&e8zM���U:�C�>AB0¦O=}�>��lQ�&��'���;���	�w�0J�@�t�D}{��ƹF�!�$��(�J��R	Kx���5��0a,6mi�b#=�.O��P��g��hYE@X	D�[��'���($"|	 �6��Y�/J>�!�DB=T�,�� �
@4��n�@�!��-,6H	�j��*�x�w�^*�!�G�OBb��TjF���0ٔ
F2t��~�[�������R���_�OVR�Z0�6D�Щfn�5]yxpi�]Y`"�b1ғ �
��vj݄K�p��ᐴd�`( F�Z�<�f��	l��و���!a��ڣ�U�<�����𭡴b�Z�٢��R�<Qs P0r��Ƚ)zD�g��L�<i���>��Ȃ��u \�rǄ�D�<1�F�[�t���]�W�f�����g�<G�1U���O�L�L2u�d؞�=�\8XI���瀩�0i3%�b�<a��ֵ7nU��N�8/�5�rLV�<i���5������ U�L����T�<�1]��n��amP$AWf���N�<s�~��P���'F2��nKA�<i&�Bi���D��#i�f80�~�<�a�zd�$�S�A%b0��}�<�a��in|*�L�2<�)���u�<� n�8���*q#	�����6n�q�<�@ʌ�I6��Ѭ3@��ڐ��m�<�b��|P�B�й/M4E��oQO�<��%yk�~��'��(`��Y�!K�<��a@:o�f�0Ga�E?�yY��RO�<���
�$�3�_+@j�CfF�<�ŀIh�0�c��(ѫW�]�<i��_-C�iG��p�v�bU d�<��%�A�!B�h̖]vV�j�H�`�<�d�!).(�
5�º@Z0!��Z�<���3=i�5eof�gB�A�<���,Zp>%��I�@��(�W�Cs�<i�j\*<�tͨw�E�4��@`�t�<�F`�	20���J=��#5̔Z�<9!b�����#�@�dbJGV�<��흋o�z����=,
Xq���R�<1n0R\D����@:a���K�x�<��에KRp��E\������Fn�<!$��2�2����lF%*�O�h�<asř�G�8�qqn�-Q�b�i��f�<�C��b�@�+�D@�6�橩��F}�<���O��Yg���v	�W���<ٖmA'HH�����"���B���c�<���l�ؼ���Y8��ab�L]�<qt��6�)��W;*�ux���y�\�l[��y��ǽhbLm����yBk�
 @�?\V�A1�#�y��Le�t�bF��Xn����V��yb`�QQ>ժ֍��O�f��
4�y��P�j4qb+͖K�N��"����y
� �}A�g��~�$�2g S�c"O�CfBV��lJ�D�[$�D�"Of]�����	�L����!����"O�,9�����0��N^�ɸ�"O��y�m��tB.��J�b6ܫA"O��J�ڳ��x��ޯ6Zj�"O|���Åm�A�FnI�DN��95"OH��q.�E~f)���u"O~A8�G�;i�8��e/��1�|Hx�"Orԩ� >�z�QR/���0M	W"O$���i�'K�@��J�@����"OL�X�jï �p,S�b=;�A"OF�z���2=<}ꁧ�2�j	A�"O�H�g-��+�"��3G)>D>��D"Otq#��׮a��cb�����5�c"O,��mI�~�xQ�g�ϗ~Ţ��"O.��fbӞ��yt)@&����"O"����3Lm��xP۳�.�� "O���e�ŝH䨼��R8�� ��"O��i�IؗX���`���oc���"O^8:���I��J�&ʑJ�D)"O>)W�Q0M�h�
TEM�]�нc�"O б�(�:^Ġ����w��	a"Oh��|��1��Ņkst'"O���(�!�$�
R��Y"O�RF��5j�黣G^1>E���"O�[���7����mz�z$)�"O�����8.� �v��8�D�T"O�����1g�|�Vk̲qF���"O `�o�)t��ڑA�66��X3"O�jS��V��1�j�;$��A"O$(�AH! � ���J�p3p���"O���!���P�8øx��S�"Oh[b�H� ��*L&'�\Su"Obp�p���Z,�5P���?���y�"Or	Y�� ~��x#�LN
T��إ.�Ec��G�/�O�)�*��We��U��D��{��'AČ�����
�>Ig��94�XFoՋ9�
i��l�C�<�d��:L@��EiӋ,f�!z���5LT:x��'�4��"��#d]�D�T�#�S"g[�PϻL�`8uH�K�h���=Оi��Y��Y!C'BKX�ے��%3��@S��10p������TF�k�����L��"<��h$��e�ٻڞx9%,�r�'U��:�e��e�^pK�eT�]Ȫ0�"e��`͌�(� �������?fl�KF�Y	F���0l*|OZ���'���F��#A#̡h�P�4���X4Y["�
�CGx|�}�u�P��^�`��O�@Tˡb�BP�M
��V/z�&b�'�����g�/�U�2bUFO,�9��+x��Y����(/H�9�D�B�����7��Y�b�՘EG>�q�w��Uq�蛥+~$��Ad��3���Z�{�x��gL�l�$3P)��u�F���G�m^h�aN2�(0	���Hw �V�i�k�I���'�H��r�S�{���nV>"�HȒ��dF=��<��͟:D����U�ɳ�h�k���<�V�Y��Vq���e7��[��DRbz�xp��{��x�r��P(
B�ْXj�����O�"ea %/��U&
�lg�]�
�)Tr�b_g�8��f���]�0`c5V���9Q.;D�Ȱ-Xj�|]swԩ1x�����֔Q�i׶p�H���H,��9�Э�׺�5�T���Q��J��yGHq�f,B���q)�����	��xtbO;>1>}��čqH����+͎GW*��3��c�\�P'Ĝ�*��� �í9> Ayf��'�:��A"T�D�O0#�6������M�T]�thǖ7ޞ ��l�8H.:�d��-Nm04��'o7v�2��E\��f���(Q�&�n��$��	�s�[\�i֧�b��+
�9�:���a�`p�XV��d��<ڃ-]N�!VGI`���0=����&��b�.�5�G,�PyB��x�<�*w˄f!�50�C9J������/w�Z�PV��!9̠�$/Y�:7D�b*�	H#̻�~'j	:bJ$\C�Qi�Xl)@fvx�d	 �K�[���k�	�_��qrT@��^@�0���$��]���ܤA @�
ė~��2i��Y�̣<��6-���ݗS�����L�'2>ٹ �Ga�G�U�u1��:�R���q!�82f%�1%�=1`�h2�ݕgDP}�ֲQF��S�? �}��bƑ)>�(d��d����',`�b�M�D-Zh� H�f5�Q�w�.1�Y�"ĵg��2���z/���ቖ#N7���c��;�-��"O����E^�`�O��C4��
������	����B�x�ń#.�|P��p��=R�w�x���P
4~�ɧ�ǩD[z�k	�,���P�#���sRN�~q�=����J���x���<!/�ĩ�g�xF�=�Z��e�^���ӌP=!�azD���M��g�:�NCM]��a���M�'}`�!1 A�0�:���؛6��$��M����dJQ\O�0�2oCYu�m�䪝�J���E�ϱ*�:X�5�Z�K��͈�j�XF�����U~b���ot��A�]Y��Ibn����[��ؒŭZ�v���I#���I�b�8?�vE˶��9s�ܳ��Z>x� ��`GT�~��8rà'3������qH5�wH�"5E8b:��nͲ<ʧDʦ/�FY;��W x����fL� {E�@�R��t�b1�	Yh���d�$+�Ty{7��z���ض�K"&w��8��߈4������v�^RbJ�~R�I@>>蒰�I3*`��$W�!��Hd/��$�ش/9��:q�|@��!�"|h��-L$1i`(�M��8��值f,�	T(�D
��1� r�⅄$��D���wT �ȅɔ�7_���C�
w�0`�R	_�@K��N0Y2�mѰgO p[>��u)U30P� �U�ܗz�$O<[�niTd^�eF�Ъ��&KqOl���#v����"&�Z[2%.W	!ڴ\�Dh)��s3˜6#�PꥯΊ#*��䀇:y�18���'[���x�8ψO�]��푝����E�m̃#-�7j� �Q��ZYpL���A�<��a�V�i(0Q���K�� ���:mҮM*�쀉Sݰ�`q$�X}�ʝ�4���M;�ON��qltx��!��<F� ZO2~8�!���<1f��9��4v0�|4�8����Or��#X;:�:�H��M���Б��LNj��$�+*s6����R�����B�)F|�q�"ZK,��Gc��) �r��&�~B�_?z
X0�hU�8�&}iqe�."�����' �<��	�=~$l���O�+d�B���`�B�|%�Y
����K���[��ͅymB��b����ܴ�I!L�2�Xp�b��� ZZm	�OK�j{��D$+)��a`Ŕ���E|F^�C%n<'$ԫ<"N���J[7Jf�=b�B�vM\����
H��E�䦟"D*pODA�ƹi�y�2��46��Ɗ;U�4�KcAO�/I�PK��0�O>�S���ą�&je�q��M��= �3U�ʆG/�iΓ<��m��t��6��
`����W�δ~�0�$.�&����$!L���M��V�r����<(f���V/�{G&y��˃�밸Y3Ҁ
�Q�Y�n�86-5i� ��s��0J�	�����Od @'�b��D��P�����k����_�TP�Or����?Ѕr�킁Eڞ	@ł�<k��8��4v��3�� e����k�̠ KA7�*�i��n���i��s����!GO�:C�S$��l�(��	��s�ؓC�
�F�z���@0n��Y��N??J�03�	Wj��F��O��&e��V�6(C�ԼX�4��p �lT�A����j~����4;Er��ЎBd�%�f֩>ܘmۃ��;�8�� F�od7��ow��8a݄6�t�;+��	�bۥ{}x�����0�$��	�$hLy�Ե ��!� @��`�Ì3y�J�ke�P1
^ �4mp��8�/�t��)�� ��J���'X�`�&˓=bX���:f����"��q� ]Fz"��2�n\A5�ݲ\i�\�%f�X�0�i3�G�v+*!YQk��A� ��e}�W�%q$4!���"D����F�Ac�XFR��Mv�xr��ȶF��!"nĉ#�n<���%s��L+$޳$�\�@�.�0Jy�@I�A��{��M���d�FM�z� Ԑ�R	Nlaa
,,O:	���$���ڴG���� �O�b�ؔ��d[rɰ� �Μ���li6(M�}M���A���lڜ/��QgO4%�A�w5�lB�kڸ[�����X���{�W�B�t����]����Q�z*Uk;��P3eA��c�D����M�x��3���5Q�!
Vd�r��� N�~������ð�u�"$a�1���<�m31�&�ҳ3����f����,�CCN c�*53��iǦ���S�4>�,z��S16������8��eX	R@"��.d��[dJĊfQ��`�D'4�*�:6��<A�H�x��Z�.��
d$��:�����Q�N����BJ.FL����,���d�[%��B�4O���A���<�bA#f�^���iT"V���K��(R��%�O��"To_�|����E��3v��%Q6��pC2�بr�X�r����c�T(G��8C��:��/W��	1��H�q@*-���+u�F�*5�[�e���ے�_i?B,"�_�u^��O>1&/�vY��@��ܿ)��1��cD"�e̟�*Ud��%.�v��P�e�<nP���b�9=;8!K7�δX������:"줛��0q��d�ծؾkF��SN����J�d��%)doQ(J�z`�+�/=����쟐G���4)'s���3�>c��Q����M�`LZka����0e�>4㶮\�$�%�7E\�HY$:���j��!���\�a�%��Q�Q���N�Kl^سC->t����$�'~�RT����:�p�����h̤~�PT�$F��>��+�kəJ��T�W�'J�����!��2�<�z�`	.�B0�ؽNQ��2�l�s��J�� ������_�gܐ���/d���+Q�I�U�M�`�M9|n�
V>̊�0�^�mȼ���V�a���S�l�	X�i�64��̏iv�Ip�O�ē%��d�``��*��6��>U����O������܁jg#A�M�P�J�7@V(d�d2f�e�o)3�(t�7L�9[���I�\�jS��6BR"ʓqz逡ݍr������%
�
�'�	����H8l&
�Y�"�+ |d(�pA}���f���'�z 'ǐ��`" g�c �S�B��:YZ�Χu�h��߳c Ɖ�#Q%��O�p�A
�bs�t�,����1b$�F�F���H�����K�%�P*E�e|Ȱ$����2�ǈ8�x�:Ag.������jA���G{����I�Ag. ��+K�I���S���Q+����Q�`�g��p�ҕX�IXI�с��U~���p��(_/�םFS|px4cz�0p����e�0�#� ZVh ��l����	(�DD�n���tI��?��:�D��^����AL������&Dv3�c3�>���l�.�{b$1c<�mZ�d�
�B͟�B��B�l�2m�Yx�� }ꕂ;�,hDa�(q��+�h�P	�S�� E��zg耽u}%��
T<����k?����U� �� ��i�B	c�`#�	�J�L�H%�Q#j�H���O������p<g��Co^@3�F20�t2W
\.w�8�hd�0�x ac�����桇#1��I�'>�;�on�I㦛�cZv�xS#E�t�E�G��6l�x������:D�_VqȜ�&m�/#~�1[����9TM#����A����ĆN�sj�I�]C` �&���1{�+#�R7^'�PYB$�lqI�E�_W��8&�0�/+ar� � �Dk`h�� $�҂&���IBȃb���h6��ExQ �45%��'�40�p������Q�F�2y�@c�/B!�2��O�	��Ǟ8q�x�ء�ߒyRHcDo�^�3wm����G�D�@��-�'_�v�f��Q[���Ѭ8�$��O����«��4D>��6�S6�J<0���'��|q#d8� �O5r�^A��?l3���'��v��pc�l�'.;���v��>�wG����:~��H7x�D@��M�/2��r�3,L��'�'<P�@�/�3{�Ё�� t�z��_��Ti�'o�� �#Ul���0�
C�?r
��v&0J�6Ϝ�e�*����A$z���*j�?ef6A�բ��>��_(&�|�+���7_ ���a`��}����gÜ}|�c��Μm�.4�"f��|>����V8b����抃�*i�%�q�zb�VI��,A�Т�+�ޝ)���u�1����A�Fn�I"ܜ��(@�>e!�j�Ш��M�y�l�iS^f���'�Z6w�FH�d���}`����>yۼA3׬�NB� �牬4���fܻvV�2���_���*��Lo؁��A� ����.^/3��8�&ݹuR�J���Y���Rs��"3��<	��T�D�=��J�Qf���DTl��h�c)�0�~qµ�PtϤ)���d��U1��wӲ 
ӮX�!K���Lռ�!7K�-*�Д��Ho���MK]Т$r�o�)t���)�l�6O� F~2E�:~�@�Ku폛a<�� �gQ�n^�S�7�$sŇ�oV���Q<�6���㊱Ps�d�`��<,�%���+8�"<���߷4�jq��^�������dy�F�j4t*B�߹=����GM)\�p���c�&r��oZ���0���?�T�lG�	���4g�	a�,���	ő.��|�g��L���
>v)y��|��4(6�&>�N�(1�"��I�'8O�l�S�
<p%Y�_�y'G��1�ĉ`DP�v� Bf$O��Px�fI�JJ��A9?0�r�k�#e���4�	6�r�)a��:��KN���(S�;"�2&.}�b�6@ԙU&�0@Q����/�0=9#�!+jdX�,W*��-��̑"��Y��NZX`*A9z��0q��[������ �ayR��?`���vN$$t����^,��'�V`i3��!x\�1�N�5gy�i1+D�0�l7m+>��hR�#Z&6��!B[��O��k6M��z��6"�)P �0�߸dל�A�.��n$L�:U�Z9���[޴:���ϻAΞ��'�4��8g��	|Ţ������#G@�G��\��aӒk�d��񋞽qS�xTHL:<5�6���?�+gE��F���,	 N���R=0�%@�6Ќqkr� �$��4h�ne@��+Xq�U"��]��jVF���؀B!�OF$٤ᇸ*�9���X;J`��4�'㨬�dS�c�,�YB��d�//h0��*9tXl;D��� '">ȸ�H�he{,2D���'`;� ��o�-s���H�>D���bӻ�VA���w�P��*D���C�8tI�����qr�7D��)u�ה�Dm� ��SF���m8D��9���41:�s�Gk<<Ƀ�<D�xa��>)8��͉r�<��;D���*�(q�^�IuȊ}~T�8D�L�u�����[�1���r�=D����ك�:�r&���u���⑤.D�@Y�Sc*���*��i���&D�q�'�u�1�q@ٍ`U^���O&D���C'u�>�T��  e���'D��9���$��t�ՒD�Rl��6D�`X�Td�j�%���ED�{�6D�t+TD�G|T�qg��_�0]�gI1D����@ޟ>c����ҁg1D�H��iϚ0�&����h�2��1D���2�$x�ЩcP!p@昙S&/D��0��$;|�X 0�W�,�"��!D�����2L4u ���7k�$4�>D��UA��3��I�i�,���`��=D��a���s���m�M�V���8D��W*~P�B���y� �
V�-D�(��oG&��쁾% ��ge$D�����s� (�Q�H[3 D���Hƚ~}�pd�޽Z�4<;��2D���.Ry�^A2W�� ?4;�A1D�� �����  =@T�K,s&@`5"O�Q�c	ϝc~ ���Q&o��%1�"OpX*@C���5ADW�u�0u2�"OPQ�˫)�0rʎP��T� "O2�"V�ؗ	4�3@O��g��|@�"O�	�G�9�^�3t��Z�|dY�"O,8� #�Ej����ϊ �ı�"O	b���}s��##�.����#"O"�)��V�qT-�a젱#�"OXJ4�Ҵw����A<asF�Q�"O0�p�ݬ�a�󅂪a����u"O�Q@Q�GR"��;t�0��"OzTzS��.��SC�g����"O��@qd���B Aq@"�vA:�"O����ط`�X}�r�&D��Y�F"O�4��l��3tf^�kX ��a"O*ERKF7$��8E�}B�l"O�8��Q<����I/[��"O�;�'M������uL0 !�"O�1�ڶ��M��CM�p N�S7"O`x�SLÍt'� ��Q�Eơ��"O(�An	�q\�`���|
�y"O���a���
�f�@$"O��@R�D�8P�(� 7J=R�"O��&:�h��`T�^�q"OX ��#��U���S��,+�"82�"O��YPm 8�ne0�E�)�l�"OX| u�qCQ��ߧx���R"O,9���ȉ�^���D:6�j�"O��wOӻ��!�����Y��a#"O��FS2{��D��Īu� �"O�����I�h+ ��pO��>���Yv"OZ��3�ۧ;T��.@":�(���"O���+$L���@;��t"O\* ��d8VH��-�[`�e"O�A�b	�8�A���-Q_~IC"Oʕ)���"m����M4C<��"O��
B#ҹ9T�K�ꑲ^'��U"OlY���xm��{��$'�h8�"Ov|avA�"@Q�cΊ&!lm��i��f�1!4�OU�ֈɑt��at$'&N0!0�'p�<� ��$��m#�r�å7��h0 �.�bh���t@�vW�H��Α��Rq Q���ybe}������b>���o�Ǽ�R
�&x �XKV��h>I�4�}H<Q���:mͬ�Y5(�L�����oVR�4��挊V���n�7^���2�^�wޒI��
0~r%J�ɖ�LGv��W%�9E�2D�I�Z68镎ߔg�a�t���E��R%	_�&t:ň#�L��	Mo��>�nԉF�'�Ve��GG,5�H��DN�	37Z�;�Of�����q}B�����^�4\���Vm,Vmz��*���'~dt�IW(l����X�g|T}�ȓ�L�ZFL�I�> 3J���	���,f¼�����6�� � � 	�@�J�O�8(S���-�;Z������D�����n��@���7P|����Y�z�N-��W�)�\(�������Tb��lEKD8|����(�XY�VI�q��T3��P--ՔX� ��+�DE{%\�?�܁c�+J�c
� ��$W�!���D�C�Z%�l�
>�䀘��O=	�V0P�I�i�T���.|O�!0�߽=�F����g�lݣW�'"���,E		�<�F)�|��=1PB�?8�X�� M�.a�~��i��=��H�Ojb�і&� Py�8H�"OZ�q��Y\�\�6%\3kxV�#HD�Ȍ��E
���3jzR�3E�D���֝-�iQl[�V=λe�CƁH.
xIE�^*>$���(0 ��f�3v<!�C�		�D���qh��BA��<L��( nJ}a�Uiwگy"��$ȋ��'��9��  ��=�$)���#�hOLm�g���<���G����r�%zLԨ�tEK�8{�`�m����%o�$��%�/=p�@�Vn�j��xt�ҝZ<���& D)�U��Ɇ�?�4g֎#h�5p�ꃖ+U�P�񀐗N|p��&��6x��%�O���䁷m̹��������!�Ʈe>~}��.��"�ȡJ��$~�"C���uhr�* ��y)���/d<�Į!�ޕj��]!�� �x9/ױ-z�� qD��(��u��'��m;en�4����̤:z�����n� dm�9=I�t�S>i4蕑��@F����d�'�(O�	�sFɆvR�yQ�G:k!�9�b�	1D��	rܗtU@T�A.�y��<����vbf�r`�̝WB�SUH�(ӞA���%��*�ء"4�'���hQ:z>DKG��<������6q_�a@0W��8�ι}(`7偙	�,+�*ߊ�T	9�K����{WBH��0�y��̮lx���f-ȻWkB��dO�I�вV��
lސ�;�f��pR ��7?WF@�vd��0��lI2G����œ,p�\`t+ڹ�Z젂#v��X�Q�ۮ-�j�c���)D���[R��NŻP��P��$�Z��xa@Dv�D�K���4/Kܼ�%���L�ǹ�V7�]��̩�4K�8+�v)Z�]%Q���pnM�����!r�|���u��'MLb�0I��0_h��Q �5-q���tDG�b�:�E)�A�B�ʙIEp�Q�i�+3Y�	�ը��!!Z�����<y����t��U��\�����l�����͖
]�j���%_�X��4�6����b"N�K�.)xa-�0���� �%��<��m��Һ�C�;�	�puJ�H����!^,u���°h$��t�T Z�$��EN�ZՂT��5F�����]�E���M�� 9�E�|�𲴪Q/Q��%�L�a_@��D"	�a�+	&���G ԣO(��` �U��A��i��J����A�#��&D�-z�o+A�N [d!�e��Ź�(�8Q�r�Ѱ�Ơ����	�m��t����T�@SdMϼ/��CN��qڨ�P�"(~�2�����=�ؠ(�MJ*欪׫>)�%���Lvն�8 �N�x�(�I� 	��D�Zn�Q��٦(�v� {���x6L8 �n�r)��
���13�(y�G�i�umS�X��#��u-BѢ�@H�D�*��eL�3g�HgBկ �Hc�2���Ika�8^��8��įM��` �+�7�����@ʍ6�ZЂdk���uoڵv�P����
Y�bU���׿o�U�e��:ur�DyYT&�Ǫ��<�
��z���� ��1�:�B��Ɖj�t�b��ҽ�+c�c���6��+T/"��@��(r�6T�@��Aw�Y^� �`�����oM� ��z���+gz�#c�A a b}��D��)`d+:��ȃ�Yo��!A$B?��,G���DcW�H�l�
�e�\�`ع Ll��q��=�،c5��<�P���-�M.�m	6&�6б7��(nɠ܉t�Y�b`f�l�|k~=jf���,٬`�ӣE
K��F a���"m�?0@�� d�{d`#>�A.��mA�N�t����T���lQ���S� 9���K�F����7k�'�>�0�4:[����Y(��� �T�W���
��ϸ*����'-�2gF�H���f��4bI�$B��vo�U�Aa��[S`v�@���i$Qp�O�%��(���R��ĩ+�i�(i!�����7/�-鳬<lOt�ۆ�]� v���`�~LH�7e�:S�`�M��K�����i�����4|�Us4�Gy%l�I�)V[�p�� ��Dt��'�h@���aD4ugc��k�� 1c*�ԙ�xʞX��n��#Z=kb�ݦ2�Eȸϰ��2�>th)Q"TT��s!�Z9+x�홓���h-R��D�� :��zU�N#@�4�s��V�_�P�*�c�,T��(:�B�"�x������/S��j��¹!�v���'1��/{~l=����.eNk�\Z6Ya' _���SU-Z�f~a��aЧ%o�����SڼI���(Ib�	)��{������C�MMҼ���D�뢌@�E� !&f^�.��ы�YX���'��$0[�	��B�W{&���!ǝk\��ߴ,&�@շ��mZ�oH�ZG�7+)�%8��=l��`fĩwf�Ƀ8���s�$C�*j$��4y_�"=�rd��D��c���<�L�7�[?(K �	ď)���I��B��
2kr+����	��T����.&����b ��S�e�oG�]Q�L�s`R*8M8�oQ�(�f ��Ŋ�<(���aT�Y��!Z^�p�����	.ylZ!i�2 �C/�>Ds �iå˱C�Pm�̃:��b
��N��4��B�ީ[��ٿ3�:�#q*řJ+6�n��
���j�:�M+��$�ڑ���{n��Y�!�F�%'��-�`G&YL�|����ri��׃����h҈t�~I��N܊m����ڀ/�.�lZ/k�έa͒7f<mc '���F\;��I�?��Q�PJ�i�liJr#��p#<q�"�/�el޶�J�ɦ�W�":�"!�
8���v�ԏ��]�AP��T+�)�mHR�ЁIږ���ye�7A�*)E�޷Oɤ�b� B�rIf��	ٚ^l�e�l��0>�RG��>����f4Hƺ��'Fx%�cIx�H���א;5����4���:C�I_rI��'���s �<$��Im~Sf�X��\�a0�k��
�d�R��%�U����@C�%��,֍ԍy\x� ��gӪP�F��(�0�0S	��p�vpǓ�<$��L$GY����`7-�a�ӡA9n,R�{
���F��>�;����#���w��j��\�@�d ,6��� .�<)���%	������Q��2��V~"�t�ƕ�Ԯ).����A�9/b��:wST՚�"
�O�R|���&�<����M5fg���%:֬Dڡo+@�`;�f��џ�aR�P=G��0���+
�,�Ѝ�%����ދtՒ��� ��Z�Y"I��D���-����@�ğ!�E#�T0.��2&�7c��@c�ABm���
}0�kʁXD��J6cK8	p��z�ߥ��$�U.c>��ېG�)��}z0+˃\N��Z#
�}���i&�� �u�׷k&��zAJ�,kwrܸ%����Ozq��*�V����_y����o4l��=��7<�,A�Vi޼�,D�k��Le�s�j��ɣ��s��ipl��?�&Q��޽��f:ɇ�H0/����	��R��	�E@�Yq ��I#ʸ���L�4���;��Y��T���"�(��l��K8e����"T+S�V��RBO�Ʋ�k@߸l%T�JU��--��Q+�c\�E�5.?�0�#�5�Ze�Z�M�so�<t�=p0���gT�]�e��;�*��#�\5 �Zv�z��~|dʐȈ�cA*�H0	�%AyHػ�E��i�O#� �%*A��c@�B�K�'�R�]� 2e#��*0��PZ���(��-��O�
�I����2��P`tK�6q�T,�Bf�-�T�a�)Qݢ`q��H�'f~��0*-�Ьj%��� ����.��-1є9ʰ<SV+�V����k[sE�۴`�r��Cp`Y#��O!/�E16�Wj�ğ<!T�	b�Ά�U�ĥʑo�I��2v1����Δ{�"t��_�-�+���i?�T!�z��|���8<p�a�G�E]a�ߨ~`�K1�V�01n�34`�R����d����aꖛ[.��e���Y���0i
�p��ub���~��1I�X�P�+l��"Ơ�Ov ��W�G\@4�
Z��Bh�A�v}��I2+��ɢ"H�9�)�  *N��������ɩ\i�G�'�� BBPjR�%w��7��v���"��Q�$%�2DX�BRhD+'��b�'��i)%.s�c�̚�.9�����P�Yꢜ�C��?�*��HYNlL��6�L9����	D�T�"\7ni��ٵ��g��T@$��I�J�s����>�b�� #'��	T���	�K���4P�G
}������R��	
t>^�C�K��o�6���k��X~�A(��L|��Ł��Y���%_Q��|��I�TdhA�a��\M ��$��7=Ը�0� ǔp<��e$��N��=���H�t���Q
j`�a�#:v���&��^���'Y'�a}B��3M1�j��Ŕ1�php�W�M�"�� @s}��Ӂ��e�7)���࣢J�i2.1xA�%|���s�@��;#�X��l�)������	@�б��g%�H�:�� b�<��x��\8JsLd�$��/ �����M�H!�N�) ��""*ڪ9�XQ��|�r�ZР^�'����s�@�V�O<!��K�E�Pݓ��	�p��Xp��t?��*^�{E豓ug�0q$��! E�m�����;Xu2w�[Q̡��l�(G"�
���s�<lP��U(M�Ԕ��S����g�CFx�����S�{�����w3��М)� ���l�O-,1Hg�_83�݁rJ~����T��p>�s�.�>"�l�[`���M��g���i,�O�H:3h�0}�d�i���FJ|d�#���rE�6m��!�V� ҩ�.z�X���DSҍU!�����萀G�����Ĺ_q�̓#,S�fm4����=O"�ᲃ�ޝe��	�@��S����J%7&�I�g0Z�:"$ B[�x���BrX=�D) D
p�%��88�1���<���M�y;��u�C��剄6Q��ӧ�� *`����u��4tz�lr� ȱ�;w���N�g-f�`�D�kgf�P 0��p�t�d��OR�}+N�06隉5���ǌ�2݉�Պe��� �Џ�yO�(L� ���7���;.(��@�@b{�胏��^��<���E˷kJ:�d� � ݰ&�r��G��7x��԰��0�=;����{Y�H�׋J�>�v�H3 �2"����a��1O����bm�$"B���	�G�lQ�F�Ǔ&Ȁ�	�(�Xy;�/L�Ru9��B�}�
-Ђ�T5&��ݒ�ϕ@�"H��t������4H�%��GQZ�=�U��++
�s��	?7�h7aӭ]ʢ�i������)%.����t��0h������x��םCv�,3�H w�	) �Ae�t�$γb$�X9 '_7�p�-Wܦ�AF��t#y��{f�W
 �p�#E��x�q�w2D�����l��t� ���H1`Cӱ\ <�O��-�P� 08��B�m��|� �Dʌ9��q*Eٶu����-z�!�
8� ���,�	݈�Jk�yT����R�,ɚ����-�a|"�Ry�.�W��V������p<�D܍R�^U���o��dȭ8(R���/E�F������I	6f!�D٠h����6�!6c�$��A��T�!�d$G�P�F"/�Rm��Ͳr�!�d�[������d}Ph���P�3�!�B�WA$-���>Q�fc��!�dJ
_���I�j[�yw�x�=0z!�?�Ѝ��B���P��jMU!�$; �Fd�"�$��Eђ
��b�!�$��?�$1���3O@�Cb3Q!��i�q��τI�0dʰ+
�u!�ΚC���&ɘJ��K����{!�S:t��ȋZ$��r`���i!�ďdH^ �rj�%.
4���Ǯ<[!�^:�2P*B�_*a�4b
6N!�Mg�:��%��7W��a��C&y!򄀝Zϸ�iaAL�FS��[��-l!�D�	+��)�Q�R,
��`Ʉ	�!�
�S�(�hu�) yC����!����~��Emi
�R�ĦQ�!򤕩*�>eӥ����"@� &A�WF!�$��].P��+�J���e���@�!�Y"���	F@�H�7Źt�!�$̊LӬ�*�2��z�M S�!�G '�40x#�,(��)�`̅gu!�ڜrL�u�+K=N򴨠�j�h!�� ���F)ǔ8��Q���\2���X�"O^В���n��
� ɎM^��c"O����g���y:�O��|K����"O��1��?�~͂Ζ�e<~��W"Oӥ�T�D�:5c"����d"O@$��I:@����b�=9�J$��"O�pB�˪S-�0�E�C��y%"O�0a���@G�|���P��8LZ�"On1"�/�0IFa��G�~>�`"O�}�S���F���/�>����"O�풔��,Z�� H� <�Q�"O���,���40�r��$��A��"O�H��ւC�d�`g^:Ԣ��"O2X��	Q�VT��ƦOSTP�"O�������<��Q�Vi��ͱ�"O��I���g��
Da_�Ɉe&"O��Ѳc��&���{� zWxU�Y�0�u��qO��tܧ0�
 �)�)vH�����L�%�����(:���'>ð�甙�YF�ݹA&9�'��pP�G��Z��O�>��G�]0+�is�G� )�D��h�ʸ�F��-cL���\}���A�C��X3��I�,D��PE+w��2*ʵ#�� ��R��#N?!�~R'E��u�#$M�x��T2�
�uS�M��{}��ҙU�2�'��*A��@�!I��ԇ̯x��q��2}�O_,� � !* ���'�t#��Է;Z���ʑ�?txz�'�Ly��eY-<�]��O?uA3NY�V���㘹oΌ�KwbF�4��p�Q�S��y���<� ���ʩav��R�IK$��s(Pk~��'�J4G��W>e���()���$'lN]sgA���dt�:e;`�ڻ��N?���q�!8hd��M�j�b����M����M��p��_����S1TRz��EϣD�Թ��HI6*�>���Z5�8Blݫ��S�O ���q���򍛤C܁s�x`H;�H�x	�x��O�P#" S]�����H�|Z��B�N�"2�O�����OO�����>U(�r�)��o��M[�	O~�@�_� ����O`ౙc�?�m
� �=^�y*O2� �	�|��|i$���|���@�A�� ct�ю`�a�I�͟pԯM�F�� ��1?E��	0��4��H^)q 
��2%�-a���'a���!FBɒ�0�b8۷��k*p�l~�OK�a��� Y�� �tFM&x��l� +siT�'�\��T!��a���[�x/P��b�)j��Pph�<��dF=��Ar`�!}���@�����Q�J@k�(��雈I�� X"'��HM�e;8y!�\�J栋���i�%�O����a�n%)����(h
�'f%�V���ۨ�"�A�,D��	�'9j�"'
�5�@a`Ĕ4d}��'�.t&���,tٓ�eV��5��'�jr��6 ���K�,��'�,]��P�K't�S��rM�q�'l� 8��W�#9�e�G��m?D�P
�'Ǌ���`��$KWb
�]{���	�'�zSn��3u�Xa�
�fU`	�'��m�t�\��������2#\d��'@Z��#BPM6R�Iv�C9)����'״��uo��Y�� ���T 5`�'�,�"'_F����5GS8��H�'�V���-�9A��	����}��l+�'`T`
tH8xGX�P�={K�%��'t\��H��u* ͪ�K
�z�nl��L�v�`%��;e�&T�6��:o8*4�ȓ/.�i�σ7V� �w�	�[�6�ȓ�^x	5`�jYӴ͏*S^��ȓ(���z�Ң*��GF�W�^��u�A��F4J������lɇȓE��kU���*{A/ǖ_}��ȓ���Q��h��x�'�Ŕ p<��&P8Q�F�m�Υ�d�:2&���p���bBV�w����a�>�����S�? �d��!��c�܀�)_���r"O�U��/K���E��FP�L5��"O �gj1��=�eJ�y0�)��"O�l�n�>���ӥ���V~���C"O�zg���v�x��hh���"OpA+��M�u�����"vK�8�"O���	T�LP��Ta� 3� "�"O^��iV���yw�T�)BY�"O�k�EQN���v ��Y�<��"O���Ɇ�w���z21�h���"O"�be ��ԁ��	74����"O0Ywl��|�ܴ#r.�>1�
D�"O�U�(]%T��zD�Q�E����0"O�=��!6��NV�̴��"O��Q���0-hv�:�\e�r�"O��r.���K�6h԰
@"OpA:���(f���2+�BZ|3�"O��`V�	7�|9�$�7dB<� "O�X��/Q; �i��쏞r'�=�d"O����&�pX�
ګ"'61;�"O��[��ɓr4�`'�+��{�"O�|��G�{��C�(�	b�Q2S"O�������h;�0�uG�$BT�D��"O,mJ��?s��!S�.w;l���"O�}@�☫i� `�&��g.�"O��C�W�I����0EԳH˔T+t"O��0�ˎa��!{�j7/���(T"O�M�!,s{�鶪���|��"O
�2� ��4���	�x�P�$"O��J��>�����)�7��e1�"O�` -�����@�U�C"O Ѡ
ŐN�:4��"*<򼔃a"O�1��L`����0K�F��Ț"O�y;��	/A�y�*3٤��"O:�!`�Ҋ@�p�Xw�L�Uľm(@"O:IZF�ЕGlɡe�ۂE�*��"O�����8\fuX�暪%{�)(T"OQR�O�`ovUH��/��D!V"OD2GɂLT0hz'�]�Qq"O\��A!��"N� ,A�ܺ��
7�y��E	�	�N��(S� t`ΐ�yB윿}~Dk�PX@�L�Ǉ5�y��:�E��,�6b�� 3�P<�y��Y:/��0�M�)[H�"f��.�yҢjaN]S`)_�U�4����y�HR),U�sdB�A�H��Q̄�y�瘶
T���%�,k�0Ȁ�h�"�yҦ�rjuI媈�v��4bF��yrf�'(x��p���gJ*iU�מ�y��8,���X�	�e+�yX7�X��yB,�'#P�@C�a6�q��H��y"*C�1N�`�K���T�O��y��]�9��	�c�R�݈-[$CA��y2��4F��ǒ��u����y��S+�T�aԮ2?n�x�,Y�y�@
#y�����oK��P;�/��y��:d}�x !�yc�pZ���,�!���1��ȃc�Z��-��LG5>]!�آ�h�p�/]0K e�i9�'��!��B�Ϟ=�0f�/K)$Ղ�'�KÜ
�����k��S��$�
�'y:�SW���rۄU�&H#c���ȓn�*���=x�@� �pO\y��qDh�K��էz0�8`��@�h���S�? -[u���.�hG�î�v���"OX ��
������_��p¤"O��c�#{��u٥�^��(��r"O�As��^�� ��L&��D�F"O��ГL�g�Pi�	�$rBܐ "O&�R6+Y|��`p� �7�x|T"O^��@gW06�>a�/�&=!
��"O ���DN�1�t�cs���3P"OPXȵ�B�v<�����o0�{$"O�y�	�^�zD��'V�_%"O�(ȢG��7����f�$!��ըd"O(\�)ߨ[����$�,��"O��MPޝ+"$�\��Y#�"O�q#Rg�*"� �cW>�|�"O0ИT@�Y��!��;����"O�9"I��2L �Ô�rg�Ś�"OM��W��2�"v��z:��	�"O�)����4�*}T傘	>� �"O��2B���HB,`�eՊ\Ti��"O�`	�0UI�aBe&U ��Ӡ"O�pt!�Wo��j���t8�"OX�;��=J�T���Σ.
FE"O�u1��/�,�V!ƛP ���"O��� nY�{�T�QBF�=��	��"O�1�`��4D�< b�gƴ�6���"O�s�bţ�ά��(˰
���w"O���Nƴ}L@3�����
�"O��	f�
��(�g�?s*iI�"OrE�2m�n3V����1U��=�s"O\53S���&�JA)�?m��5"OLpS��� B�"$s/Ʉ: �"O�]#�$�Qź4`@, F���"O0�I'ň0'�r��f�Lp��"O^��]81��U�J#`�i��"O�t�32���# �U�UD��"Op�Y	V:(���о9v��"O�!(fɛ�D�*t@�k	4�ӄ"O��vjS��!�ăU��)�"O��bXr�@��?C�{2"On��T�{���d"�?Ǫ1��"O$@&�� ]2�h�kܟ*t� p"OP}0��O H�����(g�MkW"O��3��Ց Uj$�C9%�ђP"O�	F�A"�*�����~f�D g"O�Ċ#
�bМ9&�{vf 31"O~d��`�<�p�R�B@�St��Q`"O�E��&ȵou�HI�������Rs"O�i�O��0�0C
�l�t�2"O,C��
�Vm��D�� .��"O�Ua�)
2v$(���8<�P�*&"O̸�� E ~��ǒ<"�成7"O��ꢀL�	���V�ߪ*�J�x7"O�\�����g���"�Y��y��"O��LC�7��s���ʸɉ�"OP�7�+X����U��aiS"O@!�	��5R2�+c�ץX���"O<����F�v��F�ߣ,&:I�"Oz�XBG�J#l���ۮvs�t��"O.9dہ�f��@���ZML1�B"O��/Y�d��{��ܮE9����"Od�@�O�X���C	Y�A��"OA�e�q�>��([	K3\xa�"O,�b�#^&2��5|$�Y�"O|Z�"�G0�H��?w��0"O� I���-3���;��8pX��k�"O��ȕ�D�GH��DB���U"O�X��G�	��u`���Y���"O�s��Ӏ�&T�w%LzL�EK"O���d:��@[3�P�C��P�"O�-�3Ȑ V�J�����HAt4��"O��E;|�4x��Y:���"O��X��	�v�T�`�G
9��r�"O��fO����y#`.��X5 �"O�pCф(tdقG-�<=��l�"O ԰w���qM�|Pc�
&{�|��"O����.ɝ)�e^��<@�"O�lPΗ�;c"�P�΋��x�7"O6�(�Ҝ��As"K_.z� <"u"O��X�V�V���PŪںu�lH-�!���v�z��Q� �N�y��I@vR!�$Y�nP�\z��Cy�4.Ե:�!�X$k
�j"��Nm�T��M *k�!�D�0��=HpƉ^db�J�͕�N�!��A=pB��8`N\�qP��[��C�!򤅻C� 1ZIV�"$���=!�DQ:F#�uYDOAbL�1 垀+h!�N�bJ�b��[DsD�M!�d��.ĈQ�c��6]� XB�F�XC!�B,Y�\�� /� G���#�Y�N4!�d^�`]B{U���m�~�1�(VNP!�Ĉ��^-9Ƭ��9���2�(Y�Vb!򤐠�B�"��� _2���Ļ�!�$�,P�a��־X���0DK�s !�D�+E��طlC�
�i�"$ؓx�!�$Ъ��m��ř���a�HƜy�!�%5���/s���2����}�!�D�K�H ��� %x�]�A�!��w�vuD�H����T1�!���@�H� 4A�h�٠��\�!�D̈́d�2X��d�#+����L�e}!�ӵ�4�`i:z���!��хȓG,��+���_?������Y�B�ȓ0JZ���	��6�(��҈
<�v܅ȓ�`CH#���@��"l_`e�ȓW|�p���1,�>�a Μw��ņ�.bTJ���; L� IaHY�^6����4nHBᅅ��%��H˻Ms�8�ȓ/���BQ$Ш��ȡ/7M,p ��&!RPP�j�(=�M��.w�~���iY4   @�?�     �  �  k  +  B7  7C  BO  P[  jg  Us  ,{  !�  b�  ��  ��  A�  ��  Ĭ  �  t�  ��  �  M�  ��  ��  �  Z�  ��  ��  +�  q�  � � � � =" ( ]/ -6 q< �B �D  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����ȟ$� ��@��X@Ƥ�S�Ys5"D��8a��+B-����
 Bc���*��Q���'=f���4�HTk.h+��4a���ȓ_�R�� ŊU�`us�1\(�Al�
�HO?7M\�������<�����\�/n!�Z�v��r�DL�4�:�7���'k�Ik~�)�4��"o�!���P�e��y�/�'��T��[�dV��
ƪ4�yb�	�t~��`�,H1`(�c�7��=�y"��b�hݻS��%�p�A!����M�']�i�T7jj� cV�a����'�\�k��]�q����U A�����	�'4JR�I�7<!�7���&<��'�2�+d��(my0�F�Ph�Z�'l�M@��A	y&�÷ƜI��9Q
�'��@c���W�� C�:l�	�'V�)��M�7̠�SQd4���@�'���$kJ*d^P�@���,d����'� �R��B&7���p��8,�x@�'�Ԡ��G����y��ӱ+��Ћ�'�<\���Կ1�=�`�)�~-���� \��f��bm��r��eL�t���On���!d�>�'f��[_0��߷E���?O0�7��Oڨܺ��-v���:�"O�DrP��,S԰i�&IǳI] ���a�O�4�	T��h���Ӥ6,��<��'N�#��ijd2#낪t�
x �O��=E�D��`�؂�jӇ)����V*:�y��$/cVE�t�$
=�&@��y���ĸEh�"Q�Z�{'��Px�i)�	�A�D��♙F��$&w�P�'���쏊��m*D�4 W�X0��HO�P0!Z�A>0}js��V�H�[��IA�O)Bҥ5��( �,8�,X�J<)�'rz�b?ic��Ĺ(����g�.��Cӌ4<O^"<�hޡ���r0�S�MR�ăId�<��M,6l@@f(p~�����O�ȗ'���������$���� HјM;�P 3bCUW��ȓ~x|A�6�3$��qu�N�b�%����I�)`ڬ
5>Z��aHt�C�_���d.?��vӎ]�a �E#�m��H�2=`�"O�<����2J��j�o�� ���b�O��Dx��L�`�1����:v����'%0鑠˽{.fM��!@E~���'ў��D�*9�T��6j�x1d��B�u�O�<i��I�w���U?ETvE9��DH�<y����EZ���֦A���rgF�<��,�48,��"��"̎�Z�=Yɦ�[���9O>Ip��D5x�Q���T9���+d"O��B���Ē���FVWDhcs"O2��㜔+e�-����OO�5��"O� �L"t���6ڻr'�Y6"O��a
�UϞ����A�^X�s�"O2q0��De:,�Ei�4�j� �"O�lF��E.�ЃG_3X���"O���M"h�z=	�eV�"OF�X�/��{� ex�̏X��4n8D��z�`T�^�m	@�E��]��k"D�P��͑�:��J��V�ȥ/!D� ��^CPȰ'¸0����둞"~���n̨+��J�*�05I���=PB�I�4�8Y�6�<ky�p�(]n0:�	ݦ���/<��z�3z��P)0��6.#h��H��y�#8�:�zw��/�`����'�y��#cV�r-��*:QP���y����r�F�K����.!�u�N)�yb��y��S���#	�ԑP �y2䅬�hA���� �9S�� J	�'Gr�XeւJ�v���a�Q\DܡM<q�W5�2(�"Wx$��KE0d��ц��E�	�P��p�0(F?zE�Wc�9��C�I�#���K�h���W��
�bC��<=.��U�¹'�A�%O	Q�"C�ɫ+��e�� �<,�}��H��B�I*l�ɣ��@�@Hdh����B�N#`�;�KH�V�9�@G4��B�	z�����JB@��!�C7~B�j�(�Ѣk�4�la�ed/BB�S,���c�$Ga
�zŃ��-1�C�I�\�Ё��+̀%]� �!؋PQhC�	�.�^���催S���AV�jJC�	�<G���!��0e���x��F�)�nB䉖V���+i�b�ڄ�� C� B�	�*c4�1�F6,�XMqj�7EW�C��>Q\�`柶Y�1�1J�=;�B�)� �tr�ǎ�/�����<#f]zg"O�m��E/p��Ʉ���,�g"O�q�&��,1�$B��_�B�1V"O��I�ߖ<⨩j@ S�@�&���"O��SV&r!x�)r��I��[v"O2x� �O�/.�81gl
�6p���"O���G@��Uu8I��k�49)���"O~�� ����9#��ўw��Ƞ"O^Dz�`:U�
��p
����i]�yrEV�y�)B�/�Mw�0�H
�y���`������G��a�^��y��� <"��� f��4�:����y�^<M)�q@�@�Z�i�kL�y��]�@�VD+vc\�T�4�15mɚ�y�lR��dt@�,�~iP퀅�P��y2��]b� pV!	����K\i�<�Wn ��`�D=3���v��G�<����*rR�u 5m��|��9f'C�<Q�ϒ�&\$$�Rbde9aIV�<Yf��j]��1��zq2H�bf�Q�<��GJv���	�bB
!:(��h�w�<	�)b��h�j��0c`��u�<Aũ��^��w��fpA�u�<)TŐ�2xr�p�FN=\t��bcWu�<�G[�L\5���@��Vy��C䉩m��{/�5O��2jF��C�	8�4�(R,ғkU��'�;7��B�ɱbP�D�P�exp� 6��B��KHr@ږ�\�y�@���8o|,��)�09�A���0P�!s��${ۄ�ȓ
�(���R�Sj�����0=��ȓ;�4��pƺx ���,����T& 	H�DC4./ΌS3IP�Z-bT�����ω�"s����`�P��1D��`U�ܲ��HY k��FѠ��/D���I�_��V薫G���e-)D��#$ɳ8���1��ߠ���(D��C���#�X�Q��x R�3��'D�0�C蕔Y�H� ��%�|բ�&D�t�E��<�\�1�I�X�H�w�$D���<�z�i��< pS�i"D� YV	�&¾lK�/2��r�>D��eHT�dz�!	 �#=	�i���<D����5�T�2�kT�I��5D��R��fV}P�^�Se6���?D��I�R'@<E�Ʈ]	!N��5%3D�8�0���n�������
�O��!�D����Q�s�K5P�+a�/%�!�dÐP�"��Hp���bj)G!��pwLx�����^؀$�ů���!�D��@$d�A�2���S�ʋm}!򤑱�`�إn��Ѳ�P�"¶4q!�$�����;O��X���ه?!�$H����ĢS�eojd�uʖ�7C!�SXDXk��,�@�S'��s!�G�<�<(��Q	O|���ܮE!��M�G�����Lqn��6�I�[�!�D�NqF #B��-g��JU �%p!��ԨE�J���(�3hz��3�a��!�d��}�Lt�P�kv	X0nݥ !�ǰ[�r��42=��,R<N!�\#=#�`�у�?8D�=j�e��8?!��1��h�%�ӓ�E�p���PN!�Dm��at$�"��-�aL�8UM!�� �p�G���5��a0'��%ۤL)@"O����9o�@H�&Q�Ę	0�"O�x� ]rE&�K�e�4_����u"O�u��W8~�Pt���k���"OX|�,��Q�Z��0�@�~��|�F�'D�\�������������t�I:p����װP��JSm��_�*���ϟ\��͟$�	����I֟�������ɮt> +ba?2��]���v����ܟ�	럤�	ݟ���������	�j��թJ�e1����AP�� �	ߟ��	��`�I����������՟0���2��A�kA����&$_�4���۟ �I���؟���� ����I�D&�u!7�L��1�vbއ:f�p�	ퟔ��ٟh��۟��͟�������	[�,���aH�	8�π=F�5�	ݟ��IΟt������ڟ��	�����Aæ��N
g��� �÷u�΍����,�Iןh�	�����ϟ@�Iǟ��	�b����(?O� d�ϪV�4���Ꟁ�	���I���	͟(�	韰�	�H^��� "w~�9�n�'��i��Ο��I�H�����	��,���T���T��L��nɵWZ��4��t�����D�I��P�IП���ß�����P��Bz��&"� ����B�>����H�	��H�	՟,���X����	`�|�,��⅄=(����&�Ɵ`�	��<��ܟ|�Iן��ɒ�M����?�`İGô�q*Z�Ri�Qu�S-a �韠������FŦ���9gQ��)����5���G�+S��	I��4��d�զe(��A�b��c�յ2�6Ys�_6�M��U��@�C�b~���b��p�mLj�	�	\"����Y��E��b&�1O��D�<����ӪR�\y�- )��Ha���iRunڕ+̶c�x����y7K��P��֫W�E ��J��Z�&s�7Rݦ�����i���dYk�5O@�B���!�b"q�à8Ɉ��9O�@�/�#O2��8��|
��>�j�C�U0b]a���E.�uΓ��"��ɦ��"@#����q�F�{@*�Y�J� R�?�Q��z�4��7O$�Ң1���Q#
���Q����~M�'>��P%(4E�X����o�6y�T���'4&�r��#Z5��0�Ј\]
TS�Д'��9O��Z�T4b�;C͊����Q<O&�oZ���%��&�4�(
#-\�49$�"-�IAX��P<OB`o�4�Mc��*=i+(�p~b�'��q�%���x��7�L>�B'ܚBP�	v�i>ɔ'3�O�V���m��i)4�J2z�9�O�Mo�*J|b����\� ���0d�w��Ԣ�ud(��O��oZ��M��'a�O����'T�5��E�*½K@��#<�0��0-�{���èOᩆiS�U#�=B�O�����$|��]�D��'m�qR��G'�0�$�<�/O2�O��nZ�0���Ix? �3f�L#��JE���h>��	�Mc����|�6��&z���A�]d����L2�X3��c��������yz�W 6���9CN��夐h��'mf��B��Ʈ��#���r!�2"E'J�r���;On��<�-O?�¶̈��"�{5��6n.��[��"�	;�MK�&E~��q�ړO�tJ��ߨ#@b��A�:�X�9f-m���'� 7mۦ5��*l������}��s�̚�N)L���'�v�񤓴y�P�K0��/ljj�Ari�A��g~�O����P�����qB*��R~����q�D'�x(�4R�x��<I)��;�$�H��o��w�jhR%��@ �O�mn��M�'ƉO��4�r�T�ӿRI���R�"�0�:�Ò� h���ό�����"�{���yM�O����H�;�`b�H/"7`�����Ob��<��Ş��D�妭�$ƽ#�8��d���Th�I��9�f�&��'��'�J�Q:��剱f�N�q��,�~<�h�&z 6�p	rԎ�I|<��'��ԉix�
�/�'��I#j]��/J1'��Ѥ'��*��Ey��'���'?��'U�\>-�V)�V�����gǤIN�	ҿ��o�*V��I���Ib�s�����A+��p�b=`�h$'nI����=��
t��8�II}�O���O3x=�uB�5�y�+�7!8zy8�k$N�\�:�O�!�yB��mN��#�	�C��'L�'�ҥܶ^$AbkZf�@(�T PXrb�'���[�1.�	�MK2M ��Z��?iH�"C� 3[�8y�lrp�¡���?I5P���4sD�&�O�?��\K�'e38�b�c�)F@0 ̓�?�6�Z�	2��q��������Y�)G��ď�+������D�K�X����g�'���'�"�'E1�\ {�M�'{B��'lW�՚���s�Ll���#bh��zӬD�U>O����OO�9��|��"��c��N#T��(F�Or�n��M���i�¤��۷�yR�'��s�H*~a�=Jq$�uDH�Y�]�n�5���˅3>�'���ϟH�������۟��I�b8�@Qv�W&8��Aq	�,ժ��'�T6�N
���O���2�9O8D �+Q%���S�+p�(亂�L}2A}Ӑ�oZ�?����=Y�8���Сt�L=�P��74��тS*��3H�˓)�P�[`OC��n 1L>Q(O0h�"�,����!��o�,���n�O����OD���O�<���iD�p�'ĞX� �p��g��,qH�`"�'�L6��O�O��'7.7A��uc�4i�q��F�i���e���M�`��ܛa�`4��?)$
�:{)f���L���$����q�? ���C1�P�&o׵*�:� :O��d�O:��OX�d�O�b>uĀ�(e�m�3C���Ɋp+�����O�D��3E�r���ɥ�MCO>��ìu����R��5B�8)�%C���>!V�i�B7�� �@@o���O� ���
y�4��uF׍�J��U�D)
q�����tg��=���$�Ot��'>+;0��i�;��8��0O��O��mڌ4�b�t�O�8�tU�X���K���H�O ��'�6Yܦ�͓�ħ��A� �T��u�,��k��{�P��!F� �L��'��`Î,���|�d��9��N�+_����CrI���x������O���fD�?�VTR&�5y����hZa� �1Л6�'\ɧ��'��7ܖ9�ҡP�8���C �V��hm����	�⒙t��	ȟXC���%-{�ys�*?a5���d�@��������m��?�+Ov�}��)��$�R��|���G#���&f���'�4��D�b����[�$E���<i
�D���Y�o��n��M[�'�i>��ߟh���~�:�I;oJ�!�ЯR�&Ǥ�t#΢8��]4%;�LźCf�(F{�O�r���pՙ���8�=�eA.�yrZ��'�Dr�4|���<!c�Ϫ$ǐ�Z�-�> ���BQ����?AJ>�t_� 2޴ݛV5O������d�1q�ã`ӠF-��?!'��,�8�;�@�V~��O �Y:���-"��*�Р4��h�����G�(���'���'���S��Pl!g������0|!�	�ß���4 ��'�l6M6�iޱ����3���
�d�.o��.s�Xxٴyț&�{�(� ��T6����nN�}��(��n^��A�%"��ya�BS>_���D!�`�	~y"�'���'��n�:��Ĉ8p���'3�v���=C��k����?����O��?iH,'o;���H�[F�p獁���$L�A��4���SK���{�닫T�lڤC-Y�*
��X�'T�d�B�xU�j���k�IUy���3]�D`fDJ�C�1$�~��'B�'�O���M+����<!��%;�-���ɝyH(@w��<���it�O���'Q`6u��e�.S�	Y1D7��)��6j��cb- �Ct���3�`ѹA��9��@�S��5�#Ąk���s�ޱ\��R�R�y��'���'*��'�B�)��g���ITO���~d�DW#�F���O4�����ɣS�WHyb�g��O�D��P�#�dR#͆-NO,��
ğ �'��7�צ�S�~ID1�F8?qa��c���*����K�މrOޅꗠ[�)�X	bK>�/O����Ob�$�O� ;"�ׄ� )�1�6C�b�O&���<ie�i#��0Y���g��O�7�G7+���j�̞���N}n`��dlZ��?ى�t �2az��j��"� �0�N�1/;�蔅ܰe�F�p�[��S(GQfm+��t��<z��	`�&Ѝd�f�2+ʄ6�Tu�	՟d�	��)�dyRLx��|�AU,y�Lʒ�h���FRD<���Z�۴��'v��Bz�v�۵^~e���P�#��J�p7��æ%��h�?�h� ��c�].���-O�� �4�re�� �L�7OD��?���?i��?����iO7H1`��<���W�"$���m��������I_�s�L@����Ue�q�f�@C�t��:� l��i"r7-@͟l֧�OJ`ݸ�b��y���L���j�J ;f�T����yb	W����.��'U�	�p�ɥ$��5�����EGFh0�	?�h�Iϟ���ʟ��'7M�"'P�$�O��d	�a��!��cG�#!f�8�bI!Ԇ����Of�nھ�M���'>���z��@��!�����2�H�\���0l�#`>�"K~�*� ft�z�i�������� ���V9����?���?	���h���$D�~B�I�DQ :��h�@�ݟ5�Z�D�Ԧi��7?���i�O��[iw�\h�DR��T@�m�{��d�צICߴ���Gr�~H;�OZX@Vh�NҲ�t�D�MVz�BҢ*V� H�հs���Oʓ�?���?���?�� |�����b��q��FI�����*O��oZ�6�.�Iן��	q�s�(a�L��dX��"/X���?���D⦙`�4]���R}��@7��9�n���O�G�:-)Mv�}�'�5��.5zԍsd�|�[���F7e�)���7H�R�K�䟬�����	ɟ�S|y�t�8Q� 3O�P�b��v���!��n������OJ�n�_�i>��O�EnZ��M�@�O��2@/Nx�2 ᰃ��u�dH�&T- ���͓�?yP��*Y^i /D��d�Jm��A��$���7�0!p��#~d��?�)O��S�OV�0K�G+4X��ZѥU�F�y�fsӼk����޴�?�.O�z7��IN���K�@�<\Hc�h���'��7M�Ŧ���� �<��lm�x�	�AO���@�ڿc^��УQ<U��o��^X�� AQ����X��ɖA� ����,a����A�:"�^�ɐ�M[3H�D�����c��`�v M�O�@�f��gTp��'+ �U�v`qӘ�d���?	.m0���`�!3zR,�ԇ���"���C)0P�������Wj�8dFJ�I��`*�TD��M��$ͩ'�є'"]�b>��� f�da`�%�c%ti��aԋ7� �r�O"anZƟ<&��s�<	ش[��} jƈf��d%��K
�	C�i�"���Jl�'w�/�$�a	G�%��� ^��,�$�2��;��Q@��Oʓ�h��"��=&z�S%�?�l��5���1���"�IB�'���w�ЌS	B� ��j�j��;�F���%mӠDl�<ɫO�)�����/$�(�0OM���N�(��u�C�J��E�42O�$��ֵA8�(�(<�D�<�'�?�1H¾Nh�F]� 4`*�9�?���?�����Φ�C��
Wyb�'Ĩ)���f�Xp�K�
0Ȁ �#�'��'|�� ���i�vM��X}�Jw��XR�E�Fk�9�j²�yB�'�PT�6��4bx(���X����"_@x���lN����Ъ��xpvYX���	Ֆl1E�Iӟ���ϟd��ܟlE��w��§L�� dd˲��ªup��'�x7�U]��+)���'.ɧy�Ð��9�e�-�@�0'G	�y"wӒ1mڿ�M�r��w����?���DRnQ�hD�Yȶ����of���f�K��U�N>�(O��d�O���O��D�O��2W%K%^��D�a��?k\HK���<Ys�i�0x��'���m6-�|���a*��kK��bD�kX����J}�Ix�$�lZ��?YI|��'�r�g�:�:tjv"��LRjl�ī��k��]�	W���D�jMX�;������OZʓ2 Lꓥ�Fq04�unÎ 
u;��?q���?��|�*OBEo�8&��I1a�2�KDo+K�y�ˆ�UZ��ɐ�M[���{��		�M�&�i܂7m3<���ɘ�T���B�_�����	�^���Ox�n#4j0�k�ɷ<�'9�k�������1�P�ot�d"1A���D�OF���O\���O���8���lFu;c��pV��B��'"�r���L�	��M;Bd�N~�Jx��O����IJѲ!3R�A��Ͱ�ڟ��'�v6�ަI�ӿ|�5Hf�h���ɰ56�I� �]�8[ѢT/ڀAJ�o�c�x�匃o�ly��'�2�'�R���uy�pbd��H�$��U�p���?1(O��n�0�Y�I������?]�SV�h򵬗0I���W��;h�f�;����MK��i�~�$6�i��D�񤈮d�<٘���q<�I��`M�}B�9�Ik4ʓ�ʒ�N�%7&��K>���ـ7p:��6�W�
)Խx�b��?Q��?���?�|�)OP�oZ�|�d��=Y��[F&��O7L���J�py%}�R��7���r}��o�j��7�\�DF �����lr���q�4"{DY�f(��<��l��dЗ	�(-�(O�$pp�C#(�{�ꌉo�D��=O<��?����?����?	����B�h�u����2 i��V��@|mڕn�J�Iǟ���D�s�������!U p�I���M�|�TY�b�ENy�bc��9�	b}�O���O�.���\��y�KY/jx�S�!I�qÅV��y�����PP��Q\��'������k�X��%L� c@�9;B�_�c�b��I��I���'�7���v��d�OH�đl��ԡ%�x�tk��
㟨S�Ot�l���M���'�	 ���֡�+vx�8��G@ &���ݟ�b��žZ��|[�My��O
�ڑ�I8M	�^^P� �4?\�hf#�����'I��'b�䟬ql�������gTx񠆡�ٟ��42BH��'ߘ7�?�i�Ep�b=����E*ޕtf���|����4P��e�<�A3��d�O䠠�N(�.���Ԭq�	qUd�+,�}�p�\�HE��O�˓�?a���?���?��C���q/�;�!��_�BC��X.O��lZU��I����_�s���EU�Sy<1b��ťZ��D�Ü���Y��]��4l����4�O��$C�d���Q�(!�Nd`�LI��tu�%�m��I=%ɨ��wkC�+r�=&���'7` x���4��ٸ6̓�$�����'�2�'�����t[�0Cٴ}	�I�_�A�f�=A`Y�1��^JTl�|I����Z}rGq��l��M�!�8_>����0x�IѳU�_a�*�N�<��>���h�e�&\8J��+O���O�c��.R�����6vn��`��<)��?9���?9��?Q����+xs��C�RO��9���=��'0i�^����<a�iy�Z���PO�m�⑐7�S�H�8��u���?ѮO��oZ�����2�RS	߼Y���O p�pb��r?�Ҩ�1xȥ ���5@��s�K r�|�O˓�?���?q��y��oܪntx:sJ֯M�Tmp��'{"R����4xn�����?y�����k�\ � �,a�\(q6䐣Z禠�'v:�:��v�v�L-�	g��?]�����M��<?m�@��iZxitq3c���ph�'9�D��ONf���|��P)3b�t0�����b6�ͽ
��'�b�'����X����4YD�	���҉=Q6(0sjT+\p%Cd���D[����X���DȦ1��q��ܸU��h���2�\�M�'�ioJ9J�1�y��'����ь�<Ȯ�qP���5˃�j����ƨY��H�$J`���'P�'��'h"�'��S�|(�i��Kl4j9"Wi�q,��y�4e�ly͓�?������<��y��3X���{D[�t�&d�7�Ϧ�����4������`�!��$�Y�:��t �I2�F�D�&8"�dN@Ė(��� f$X�O�ʓ�?Q�{�W��_)��;dl˄J�x�j�O|���O����<A��i��� �'"r�'s��Q%,�)I�����FV��U�D^B}"x�Tl���?Y�O 4�2�Ρ:(Mi� �:K�6�Q!4Ob��ҔFUd�Ar��=R�ʓ�2Bķ}pTH	�^(�5��d�ZH���ݾ}������?)���?����h�z��ΊD	�ň ��]����/S�S@���������By,a����%	y.A	EH���<�Ԫ�$��	��M��i�$7ME���L�s8OL�$��2ZЍ�n��  ���.Mf���0FU? ��؁k=��<Q��?A���?����?��o-$��[�L��m�|\�G�
-��S��͑�dZ�����ԟ���v��'�����'�wܘ�)C��S��t{e��>်iDP7�\۟�'>	��?���˝d�dA�F�� ����.��x��({��Ly�F	{6}�YdVQ�J>�(O� ԍ� h���b���8eP0,�O�d�O����O��<Yg�iM2�9&�'{�U*��ˁQ�r��\%8����'��6�4�ɐ���%�ܴ<ƛ�	��RC�(3��R"�@�B�Ǖ$���`*�2�yb�'a||�pf�nE��1u[�t�S��5��}+M�EùB@�F�E�y��'Y�IIy��� �;����ހ���g�?+-1Oj`l�0�^�!!�F��;�kK��JP��JN"�>�B�i+�6-�O~h{U�J�b��OF�a�'AQ������ۏN��ɪ$!?Vb�lA5*T?��=ͧ���O�%J���
(�,�	R=�0�D4OX�O\oڷD��b�d���?Mh��%����$�ѸxX����)?y�[���޴i��v9Oz�v�I|tJ���/̸L�\�U)��h�Q��gθ'��C�����ӂtE(�i�_��4��&FSce �aa��z��(�'|�V�b>�>8�v��(w����F�p8���i_� g(�`�O�n�f��|ΓS���©_!-XFFٺ<Ծ`��EФ�.6��O��:$@����O<0ZE���p�eI����В�G-�<��0�������@?�����'��>!p�/̱zDhd��̗�p|��A��M�W�M̓�2N~Z3��y�!DiP����f ��$H���t�@6�������4�$�I�O�T���S=&��D�/�`(���P��P,T��D�"1���z��� �0�O���|�`����I�8V�ֹ
�E���}��?A���?�+O\�n�k�T��ߟ��Ii��J���4�*����):����?�`U�i�4{����O��k�X�5�J�O�|��U��_��I��?y���=��n����d�������
:s����	>�;�	��v�X�ʨ��d�O �$�O0�*ڧ�?!�R$n�6�c'��rؘa����?I7�i�d5�s^�@��H��O���j_�Q����Qk�z��G2��������48����7u�
U{�'�bйĬ�kG�/����ؤo��ؚ"�H=-�X�ם|P�p�����ҟp���Ps3Oǆa��tR���,Q6���g@\dy��w�ԉ*B��O �d�O<���$��Q��D��1+�t��·H8ju�'�D7mT�������'����o�X|�D��E��m�"aFa[l	���8���/O�m����[K씣�g1���<��C�1������L�)���E�?Y���?����?ͧ��D��H����(v��Ҩ���Ԑ8r`��3�4��'F�As���f�JoZ�t�ܼZd��%%��)c%�0"��)f�EF��ϟ`#��'At,�j4�yB�Oa���H��p���J9n�i���D���Iן4�I�����şd��S�'D�d��ԅ�K=� K�c� Z��P���?����N�$�剈�M�O>9 ��;pL�d����P��F���y�T���4~+���'
�8J%�yb�'1@�R��].c��!$��{pn-�1���X��%A[�"�'���ȟ��Iџ��ɣi�|MzEɐ/���g��)�0$�I����'�6-�4>��I꟔�OƠ%"4�_�M��:�!�f=�D��O~��'}`6�P�i�����'�
���nY�YS� C�<Y�E"�������·@�
(O�I�>�%�/�䑢t\IDB�JOb��
� ���Od���O\��	�<�Żiz�=�\>�6�B��=at��5�8���Ϧ���D�	=��D��y��
4�8{ �@eJ�p;�xoZ��MS�
Iw-P���?�p��4Ix8�1��)���L�"�� ��r&~���bZ�0���<����?1��?y��?�,�>��a�;�����Fk&�|�.�ݦ��*g����ܟX&?�ɲ�Mϻ%�NI��\vhv���+^�9"}[��i�d6��ڟ�֧�t�O����ѱ$�pDz�'�,D����}���R��7'����' �#����8r"�|�X��������4�ǥt���S��-=r��_����������� �'�7�R#�����O��$�?BRxu��`��Cv�\�����R��	:�M#��it��$�>1��E!�%�i�-)�U M��<���y����QEQ�z�	b)O��I���M!��OV�� �8H�D{"�}�t-,.m��'
��'�2�s�r2ȄRC��y�,��l`p�%�㟴��4.o���'7�6�$�i�r��	4���5!�?V�>Lv��	�4y��&�u�6�㵩�3E���O��:$dq�!�fh��ڨex�J֟	�X���H}��O�ʓ�?���?��?��}��FBV8��+PU�a�\�-O49lZ'Z����L��h�s�ps���-�|	q���*:Լ��0l
��D�.��Ը��i�����i韦`�6��c:)��ҵS˰5�⁳4���B�<!�l�4-��19W옊�䓭�� �H��ۣs�*u�F-�ha����O*���O"�4��˓t+���	��y��E
r}<�����E)<��4F���yR�wӴ���O�\mڈ�M;��i�E�p��y�z<�S':W4ҝYC��T
��'0b$�	��kJ�y���?�3\cZH${.�Q�V�20��J�tS�'���'���'��'�� �
�m��~����I�;9�V�E�O����O�`oژBê@�'HL6�+�D�$a�BN]+ky�i��j�#�`��`}r��v�m��?�%,�V������8:�'� �8��&�Z��#g�Ͽp�Y�GA>q���7�d�<���?����?�D��/Z@��2UoR�~�"9�r�A�?�����L��1��w���I��\�O�FE��"E�����A�]�@�C�Ot�'��6m���������'�z0i��W�	����x��Ƅ��
�Ƭ�抽 �\0J,OR��������>��1�Z@���ULX�&�z���O��d�O��<���i?hقVNQ mV��6��*x���p����d��9�?��Z���ߴ~��!I�L�')w\!��&8>�J-ĺiw�7_�%���?Oz��M2!�D� +����?P,PeoE-��0Qd/�1W�VpΓ��d�O��D�O���O���|S�Ɩy�r%Q{������@8*��6e���yB�'�2���'
:6=�B帄g�'5�p�C 3A"��-ܦ��ٴ8�bP���?�S�v>֘��ey��,9R��@aE��R���&lx�`#%�(w�>x�*�o�	hy��'�rI�4Z�h�yb�_"���%�Ãc��'���':�-�Mc�O��?����?E�Ӽ\��ߢpO�-X����'���p��ni��9�I[}��0K@R�Ae�V�o}i�Q�� �y��'cjU����9ۄ��gP�|�)6�t#&�^۟��Q�Ҩ�L �+�l�yī[ܟ���՟H�	ȟ�E�t�'	���Q�V>l��u�C,o��H�'�7�]�jʓ^�6�4���R#�$���L��!��<I�i|6�¦���UUJ�П�P���u�-b��5�Puau`P��tf�B�$�&���'���'�' ��'��}K�H�%�2�b�hJ"\��(�\��{�4TR�����?!����<�C �$������3�5أ�Cc&�ɿ�M;5�iy��d$�)�v��ū~������˔\p��է7R�%KS� 
}h�H�N5`0j_� nb��J>q(O h��JE%hю��Q�@>K�Y��O\�d�O����O�i�<��iެAq"�'� �5�i�b� �ˊg���'o~6m7�ɶ��$�Φ��4n	�&@�f,`fɕ)p����Q�p���B&B��y�'��m�4|�j�b�_�����5V�F�'Td!���g*�Y#tB���yb�'b�'k��'j�)�-RÞ8y&���U�\/���%myB�'b7�C�=���M����j Z`d�-�<����[ y ��'C�	5�M�!�i��dn��0���'w�(�G�o}r0��j�by�}����&��Ph��c��#&�|rX�L�I��\����t����1DdY�l�	�b�x�M�����Eyb cӤ��2��O"��On�'c�	�0�ՀqO���
��G���'W��b#�f�p�*��	[���G-�_=��I���#�����)�����X���4�V-����0eP�O���Њ,=��`�D���:���H�OX���Oj���O1� ˓jO���W�06i�Bǃ.K09�e�^�6Vz�+!S���ݴ�?�J>�Y�\��4q�P�`	�~�F1cG��
���a�i"6���C/0ݑ�=OD�����: )V0p.(�+O���B����1r��5h���K�8O��?���?)���?���i�1��l"S'		{����⋑FzJHm�M���ޟ �IE�s��@������-?��=a�$ � [��9v��}�rT��m}���oF-N8���'on�QQ�13n1�D�߳r���'� ��i��r��}*w�|�Y����ݟ|sǅQ/���y�kH,Tej�铈O䟐��ȟ���Ly"Ie�$<���t�	�p���R�JANؒ���E�FL�d�?�Z��޴՛f��OX�N+�s���z���kУvq���'�,�X�$�1U��t�E���kX+i��4���'w�͹4&��>�(�C͖�g`r�9&�'&B�'�R�'2�>����?�T�w@H�\�����U�Jm���ɹ�M�K\��D@צ��?ͻFxP�"���:6)8d�$��E�M���k�
�l���҃j4?�u�V3eŪ�Z����H�cPN  ��j�b���J>�.O��D�O<�D�O����O��X���BX@�T�ϱy��$ �f�<�`�i��y)�']2�'-��y�hԭE��`+�jLQvD8�n҄<�u*�An��A��a�O�ⴢ_��ɂ�=D'0��F�yj:�u�Fy2D��?�b(�+ցwa�'��Ie(��+[7c�L=*�#HK�=�	ȟ �I� �i>��'��7��N�v���<\.]��J�-5j���\|��dEͦ��?�tQ��ݴ-�&�Ӛ�y��!-|2��ųq`e�K��_���0O`�U6%�nD�p�Z����b���}�R�D]p�=/�Xd0�9OL�d�O����O����O��?���³=�J�!��F/3F�1a��l�8��ߟ8��4�l��'��6m1����#�4�b�5S��L�
 Bh��c}b�i��mZ�?U���7Ik��ʟD2��O8l/"U�4� [�<b�.�z@�T$�$K���%�D�'tB�'��'s�@��O�pd�aD�`�\c��'�RZ��XڴC�)��?Q����)�^�����k)�@�ȁ� E�������Ӧ�Iش~�����O.`0I���n7�q� l�3��lرJ
EhD������?�;����}�'���v�K�y�Y��S�v����S��� �Iʟ<�	�b>�'��7��Txhy�
U�3hށcd'B&8rp(�e��\޴��'���<Û�k�Ԍ\���J�@�&�i��6��G�p��6O���W�ݲ-�e��}��{`ٱ��כV'��{'
+��0Γ����O��d�OL���O���|"�߾�ZhX~�,��2��9iW�FÛ<�y��'\2���'�6=��x2�-h-t!�'Bޏj��l0@N�ߦ��ߴQ�S�b>�
�뙉��)� ����/<�@rś�]\\��<O�¡ė�/�!��*��<����?a�%V�f�r�5�d4B\! ,R+�?����?������U���Fi�P�	ԟT�҇ƜWb]R��;~r<p� IG��]l���M�6�i
��ĭ>Y�H��$1|����5Hx�a�(�Q~2.�=E�jyC��P2+��O�т�eP&+��Y�Y��eɁ`O2]h) a�F+*�':b�'���Ο�1���+B=�g�k�@�բH	���	��M3Eo�W~��tӄ��4�4�&�8Vg�U:Zlz�':WyЈ)5OvLl�M÷�i)F�	�Ǳ�y��'�ֹ#�Iēx\�cL̅n
��)3oE5��@�!��'4����I���П<�ɓ'�������Q�ք:���5�~�'M(7-�W��Of���@��<9�۽p����a�?T��=�G�B�9��ɞ�MC��i���?������#]���sζ0
έ�A���CI 0hp���P����2�0��%�F\��ryr�^�9�����;0�@��:6���'�'��O�前�M3��<����iNU8�+%Pv8����<Q�i�O�1�'
26���%{޴6�}a7,Q�BȌR�hNj��ыs�5͓�?Y�N�NA4�PW,[���������:� �+��!o��a���p �]��?q��?����?����O��-x5 �v�Tx��&��߾ٚ�'��'_n6틷Q���M�J>9���&z-.��,I���H�+o��W�d �4+f�Oy����l\2�y��'�|����]"Y:"�i�S!2`y�S�	�UZ�S��f��'�����ß��ɮsI~�p�DE��h  ��NZ���IƟЗ'7�9r=���O�d�|r��T-`Ai�(H�Vy~�M�>�ĳiN@6-�˟@&>���~D��↜W�. Z��!#���G@��S�eP�� ~y��O[ʡ�������'E,�+��
	�� O�$XH���'j��'�R���O����MK�I��Pp|H�fMY(=	$�˸d���'"�6�0�����$�����a2o�t�����ӄd2��M�׽i��9���4�y��'�:3��8A^���ы�H�%+PhS��1�e�y��'d��'���'�r�'����^1�̟&0��OU�fW֘yٴ1�v����?	����<����yg%H*Q	�F�x��'&��6MZ���x�����Ƣ�Z���5O:]��J, ���+�E�.F����4O��BNԢ;"X�J!2��<���?�������J1�:$(b����?y��?���$��Qg"AПt��㟠�F�!��ҷA��+E ��6�X�+��ia�44�����O���-"-N�~��� $#'�P͓�?Y���f�4l��������j�B4�ˆ:Dp��B�=�}(�k[3!��T:r��!&Mh��O���O��$ ڧ�?Y�x��I�/Ю7�u��aW��?	��i�����V����4���y�֨y�`�U�ăG�d1"7摒�y�!m�lmڷ�M3�LB��F�ϓ�?Q5�ȮL�uC'���#���+��^�_��L�����L��`I>�)OZ���OP�d�O���O��WOZα1!g�d���eA�<���i;����'���'���y��/1�n�)��0@����@.
�Z�X��(g�&�	K�S�?���� �*6/�L@V[�%�iF�Q�`V��'�(�&J��z���/����!�ĺPhw�nm;���+�"���O��d�O�4�ʓj훆hN	tG���?&X�,6��Rː�����9�yBnӖ�@��O�l��M�D�i��C��G�`#���g�]��,j��y'xԉ�O0�"4�0��,)�i��SW�ݥ$֌b'b��}����<��?q��?���?��DNОY6x�a����8���y2�'���{���q��8��4��y�u����1'���TiC�Qx%Y�'�I0�M˂�����"ly`��O��c�)n�ȉ�"C5��?�� 1aΖ> tB� K>9)O��$�O����O���E�h�n@����:���1e�Oh�d�<Y7�i��ɛ'q�'�哑ވ�AQ�ƹr�ZP1�e�$+F�)��ɴ�M3 �i{V�$8�i��<�%,\<J(�Qz��Ѯ&&�p"�#|�����!�o��˓��E���s�[pL>y�A�*%�]�ek3�����҇�?���?���?�|z)O�l�s*�ѯM#I������ÚPX���"?)&�i`�O���' �6M|85�R��6%~��ړ��^�tm2�M��D�u�����?��(:o�@�jE���ĚD2 EQ�^Eip쀂EY<s��$�<���?����?���?�,�l��H�
"��`�d?q>Д�r�Ҧ��d���	ٟ�$?�	��M�;A�
��`&�a�\��U.ʎ"�X%�iP^6M����ק�OkF<j#"��yL�r��ɗ��;%d���J�&�y#�R�$!y0�V�+��'��I��\�I%9��Y�گ[���J�=?����˟���쟌�':6��-^���O��d�>%H����8j�89bU��5K*@� ��Oȸo�?�M+��'����8�¥�n�*_�|xƯ��>�� ��i̩tr���cyB�OUV�	�C������=�	ڠ�H7p&!��l�pj�',R�'���Ο,ʷ+�(/����!;�桚�����\��4+�Q!,O~loe�Ӽ�a��(���!��j���<���i�6m�ߦ��G!	�I�����`ݽ���`k£e�d�&�j&qH�T��,�'�x�'���'@��'��'�(��y^]�����=ˈa��U����4<���I���?A�����<���[,_O�Ő��S���$���T����M���i#r��9���.�)�t�� ���f%V� 9���%��N�.l[r(K	:F�˓*�,z+ۿ/#��M>i/Op�0�Z+z����"�T6hTX��O���O��$�O�<1��i���@��'r$b��Z��9BFǤ&���Ý'��76�	�����צ�A�48���Y-7����'���QS��(W��	�B�!�yB�'�����91��&_���Ӝ�5�+�Q��Br�ټ#�+r���y�'�b�'���'"�	�[��Xqu	�x��ͩ��5@|���O���^Ѧ5�6`yB.j�����<�t���&Ya����K�U���d�'L�	��M{�i���o��K���˟'k"ꌹ7�`��b�ޟ~�V�0ܵ
��TpA@��P�i�7�|bP���	П(��ɟ��(
�g>�E�F�{{�%a��	uy�Gw� ��WE�O��D�O��)���å��h ���F&��H��������O�qm���M# �'^�OJ�$o�#r�x��e��4��=�����*����i��VF���Z�����I`%�q�I�xԃ�ܣ@���b�e����P��ퟸ���@�)�`y2�b�&�Pm�� 3��RET��>��f�Ւ�w���DUU}�i�:X�!��a/�Bƃ�qDt�K����4]m�|"`\�<��S���M-�@*O��2�J op�H� C�	D2�A9Oʓ�?���?A���?���i@n�hYǆ���T5Y���yj�m��И�	����A�s�$����ՂJ�Xg�HBaX�2���`��1I�g`ӄT��A}�O����O�:u+��
!�y��	^����B��\#�T�y2j���Y�g�1y�'�	ޟ �	�w��ٻ#*��m�0 i��x*�����D�I؟ĕ'�6-�6X�ʓ�?	E��5�ˢM�a���`�5��'cT�oe���w� ���J}��ůi���snH�� �����y�'󆤑#e�YF��bQ�<���x���)�DKߟ��ŀJ�@��qd�� ^b�����h�Iş�����F���'�hh��'Z|:�P ��L��2�'`@7�ʓW`���4�fI���(e�0�#u�=b���p4OLo6�McS�'p�xI�Sn~�f��p�Q�ڎT�ȁ5��[�<�)
9�ɑ�|�Y����柀��쟔���L1%�DH6)�刻�*����Sy�Oi�l���O����O�����C�x�
�� .�#�@�'����'�$6�⦡(���ħ�����pUj2튑8�b@�mM�)�,���4��Y�(O� *FńY��D�b.���<�`�tʺȲ�O�9t�3bF��?���?����?ͧ��D�Ц}�ğ"6�Mn�P���oa���+�o��$�����?)�]���ٴ|�^����/��@ST�� fP3�cB�_�h	P+4�yR�'S&4Wȟ0���Q�X���S�5F�*8N��"f� B����4����y��'J��';��'���?qlB@:f��1RuP���/ *˓�?� �i� ɟ2�o�G�}���5Μ1T��q3�O�78����������Xش��Q�4q���ϓ�?Q���@!���1a�,���l�������\0�I>�+Of�d�O����OHc"h՟ ��3����L��fc�Oj�Ī<�0�i���0t�'T��''�$�Os��m�M��e۶n�Eb�O�1�'�
7m��-K����'�
rg�7G�iI1�G�2���I�/�w��dg�2�z(O0���4���,��߳��k$�˪F@>�kQ�׃Y����O���OH��<Q��i8�3�`��V%�Qr�"q�I��M����.q�	
�M[�Γ3[!��Qb���,Tr@
3u��&dӨĪ�l�"�d�O��V�*�f8�U!�<AeNE�5?&��s��%w�Z)h ��<I+O����O~�$�O����O4�'0�>�����<&�졵EI>\�n�2�iL���W���	Y�'���wneRW�1F��"��r�A�j}��`n�?��O��������08R�3O�u��bB ���*�� +K:��c2O^p�+�2 ����>�d�<����?iTkő�.q����|f&P	qn΃�?���?q����!h�����I���/tf����w�X!�NG�M���?I2S����4W��F��Od�u��,���.�h��iQ*��A�'9\4*���z|����:Fz
u��'d2�	��'A�t�37cA0a�'���'g��'0�>��I�_H0鴄�6P����$��P%b��ɟ�M#�f�4��$Z���?ͻ>�\�*�D�n_�Բ��R ��U̓B4��agӨ�m�p&���7?A熋}����m�$��D
n�$� �c��b��I>q/OF�D�O>���O&��Oȑ�J�
��"懊>"� �
�<�'�i��<0A�'T"�'���y�& C���$MC��.�P��S���	~�gn�FT��|�O���� �p��%�(�1q�M3Q���g]�� F(^�\�f^o�Hyr�`�a$�3/���P�뇁N��0R��'"r�'�b����V��J�4_c�9)��_���A�gn����J�Wx��
=����G}�e}���lZ/�M��FA��x��^-��`C��e^AI��s~"�.� ��C��4o�O���qD�9�e؇4l2��)+Y��	۟�����<�	͟��T�'>�*PR��	9sl�B ꆟ����?q�����B�|剔�M�I>y����cp@�1T��. \ڤa�΂6:W� ��4V���O�^A������d�
�R�Z���\����+O��K�/���y$o$�d�<��?����?�s�MŦy���<s PS�"<�?�����Ǧ����x�Iܟ$�O6:���+� ��h	�j�=4�2���OL�'|�7�^ަ����π V���X�]	��8e�!RM�����B�Mgx����1A��|"iF� 9�O>�r)��
2&�I%� t����Bb���?���?����?�|�/OЄn��.8n(!!j����a%H����dRyB*pӦ�@�O��l�' �\�P�b�b���EP���SٴJ��"��l��ORih�-�+1IH��b�<Y4��*M�r��D��i��`uB��<����?����?q��?����?I/�4��Gi
Tc���oX�U����¦�Zv�1�M3���?�Oʮp��?a�ӼsԨ�&�F��1N�11a�u�5'"gě�p�F���ئ��i>��se6M�?9ߪŉ�9Ow�_�$�ظ�sm�z��%j�'�UJ0����X(E�1���<q���?)DꌅE~���'�� '�?����?�����D�̦�C�h�\����xW(W�.2-s��$9�H%��n�L��^��I�M[t�i���$�>9呭��D�2�Hн�@�t~Bf��*ԓG���a_�Or�|R$J��a&r��(�ޅ*Н/mX�#�4�'��'��Пĩbԟ)8%��A�y;��rGߟ Yٴ �n�'��6-)�i��c��S6P����
wΊ]S��f�dJߴ��&�}�~ɚ����u����v�0�p��<%�<��� ـ|�!�Zl�d3�BW�	Qy��'�'n��'vR��"C�� xT�Xd�z���n��ɰ�M�+��<Y���?�O~�D�4��_O�]��JQ�l`�RT��x}�{Ӕ�lZ��?!��ɑ����1�6v`k7IW+טd�SG!0 �C��(굁C�`HK>���?!&f�n�I�+_�N�R��ؼ�?���?!��tK��O�$�M����<�G�3>���:v�T6}��tic���?!����|B+Ot�oZ��Mw�iT���B�4��� f�[2$�h�c��00Р˛'�����(�9XR��4��	�?Ui^cQdu�4�Y�K.��q�Hܙ2	�����'B�'�2�'��'m1�l7
?F� �u� �����=+���Oh�dX�����z�0��ϟ,'�Ċ��(Z�x�(� :��4��$*�?�ݴ�?ҳi8�7��Nq�#���󤡟����L6+��ЗO� k	��$��q�N�rq�}��IП�����I̟���� X@���T������܊$ϛ�K��	��@y�tӬ�ic1O�d�Oz���hM�A��2�B%j$�A':]�%Pr3O��O*m=�M+w�i�7�|�'\����e<l��8a���D�z �e`+Y�d[����񟄨�Эݥ3^�s����"Dtp��ȇB&���"D�� �+vN�R1b��g>�џp��P,H�p4\7�⽻�A#h@ڑ
D\�V���(u�������BJ�TPW(�/{���P���1��t �lNK�z,$�cg�p�r/I+ �틕-ژJ}�C�-�2��dB@!ܵN���	��7ZÚ��M@�2zV�bwh� z�j����U"�G	f�r�I�\�S���B�@ݓrd�$�(��⟈&�,��⟈�A�X�c�z�KS�ni��" ���b}����l�I�T����֟!���M�t�ӛ.圬�Ռ4�V	��/Չ5��П ��`�П$����f����r�� qe�("[���ƥ� iLhH:�4�?���?���?��?$�i���ŕ9��a���T,/�4�$?X�6-�OX�O���O:�@���O��$�OR�[Ҧ��-;@���(P��5w�X]���'��'����=1�*����:X�$�J-[�g
@
��e���k�I������)<�d��۟�����\����H�@j�+٠�I�C��r�h��'8ª�"��p��ɒp��� l��%KB8�ÇK3V�C䉭q�li��G͝~��&*�8��z
W�#h�$@̍`�j��!B�a�(�Å	�V>�,��(�2�x��	�t��BD��3&�H C��[�d��q �4rЍ�5G����	�!,J��Ƃ�%2��0�^�x�xy��#�C���h @�?��U��+]4l��WM��M��%��cݖ���?I��?���X�d�O���0��/Mѓ��
#0��glWԟ$�bަP����^6����A:�$� ���.Rd�f�*�(��/_�bM]֪x���?�=9D�?S�x���xe$p2�&I&�?���?Au�i��6ݟ���L�'��ĺ$��P�܈�E�G�=4]I�'!�*���'s�L�*�0o�U���1�p��Eyr�	+?��]�X؈T�c�?|�����c�F4x�Iߟ��Iݟk�����	����G��(S}���*�&�Dx�oY嚌x7��	]�y1c����<a�aJ<}�0"�5B�P�S7�R�n��H�4.<H��"����<�.Aٟl��-ך\YCL�� ��]]P��J<1��?!�ʟTU!�̄ ,&9P�$I�c�~��D�' ў�!�ө�|�I�g���B��w�`Qش/���Q���鞑�M����?�,�"m�CK��@�1��b͸J� �D��9�����O�R s۸ҁ��R�|Z2O
6\�UXg�:�����Ǉ~�'?�TRqIN&`{�>�!B)qF�p�Y2}ߦ�a e(�Q�0�I��MK�i�BW>I�'e���r�<
�0���S�����s�
P�
S����ˡ����s�=�O� $�Xb�/[�K4Ĺi��G
}���{�|# �������П��O�T�A�'xb�'�j$�ћR��[��A-?D	F�Θz&�)�!T����z�x��˧���<	�&Q���jRn��3~؅�c�p(��P�%�����R�mB������X�֮� ��$��F���o���ߦ��4�?a����� �:!�̧[J �s5ƀ�+���6O���'���'�ڤ�V��/ _�E��#�!&P:5�y��'�7�^ߦ	'�D��?]#@#Ӕ���J��̜V��hOڟ��	>}$�$K�h�̟l��̟��I�u��'V�,�@`�0hF�_�c��]
u��<�y�ĘQ�05�X5g`�y��
Q��,��]�8}2Wi��=?�9��J{��d��>c�NK�OH�K���
t�:1�i=N��3�*Y�{b�d������J��e��t�'sRV��Ж�gLrdI��˱��x0��Ky�'�����#|����僽$l�2E$�,���ߴU���|"
�|:+OL�b(R��䅥�.(�2�߀?��	�S��?���?y��O��AC��?��O�<�����?	�CR�x�0X��`��cG�UJ!�Ns8� p���<1E"��a�N�'B��L�@����_n8�L"u��OƙlZ9�� 
�&��/�1��@ATC䉀%\*��e�#m��U��CF��C�ɕj1�L����Z�� Q�h�3*v��	���'G � C`����O��'S��`�ӊ�8-hR<�7B������D��?���?�0lU�2���2�ӡ;*���S���R��2�I��} PI�����(O"Tˢ���b��Y�]��O�Fly4d͔-y����G�y$ ��B��
m�"�m�ߟ�O�N�(Wn����AyF��p�'��O?�� ;�\�$��51�u.ܢj�V��dBW��&%Jaj�̑�*��EAE)P>u�N�JU"��]x�d�@���j��`Ɔwu�db i=D��`�'
-k֘��iB�b�H��8D�hR�0A�H���[8$QЅB�k!D������!N��!HĲ,M��j��*D�`�#b�%�,I��`��Z6zI�,(D����U�`ݔ���L�S�l���%D�Л�"V:�4�a�GE�Q�iC�$D��@#[�/8���B�B�,�TB!D� �*\�!ɲ܂��K��Q�7�=D�|���"vh��$�@Qt�W�<D��6nX4uJX��'��L�V��b=D�(:b�^�lO��녥��#P&�Z4+1D�hPԮE�l�R��6��!#�@��.D����|�P��d-ZS��T��.D��I�V�p"��9֬0w D��9�І)����Q!��e�d��B:D����D<?�t��"�ɱb�x�"�a2D�#�&�[Ў|���H�F�T|@�g5D��a��c�R���C7%D|�q�8D��"��h5i��	ƂzW���#D�̋��N2.�H���	x0�w�+D�H�� ˄ q�ya(XJXY���4D�P�%LߡtL(ܩ!
p
:H�B.D������!0a�6U����/,D���#��T�4�6qE	5D����ǉzp���G�h��(2D����־X+�Q�+�<?SPtQ!�.D����j�3/��3�JU7�x$���+D�h�d�P*ΞMQ7�ތ0|����-D�4sc�L6
�6lr1K۸%��ы4�,D���W!�E�8e��- �1�bO D�T��,"X�W�#�d�X �*D� �Dl�6�}���K�Y:�ӳ�(D�j��ު���\3m���/(D�Ȩ��3d����-Y�E��ؑ-4D�Hq�[9a<��z4��0뤤��-D�Z���>P�(��%~P��*D�<�u�\��<�j!a�7Gf<h��5D������4�:d�iZ�\K mp�-3�I�e6�ؒֶ'�����)�8S��O�q��J�E��9� D�E4�+�H
�{��Y b�3N�TpZ��'"�!�
L6,��� ���87����(�;R.�e�fG,B���q�'�B�Q&h��{ NH�bO����ԝ^="��h־T'0Ũ�,?LOLJ0cO�SbUS��T�/��z��Q-R������I�L(DQ�	ד'��`k�)*l�@D�=� �ܠ!�S�7��G <V��R���FAz(z��-R����x��'b�٩q�2M�ȰV!@�/�b�x�{��71J=��^�3��hx�L����2�@)ꑬ��T���a�1e�$�*w��^I�x�$H	
��Q
ϓI:f4�WH׷.H��7�Y�r{�A��kV�;t|�O�=�$(����H9H3�ʽbR����+�Qt�Ԩ��$4�� ��@�G�����;+�x2�'M.p�� 2��|���ky0�/����䊊��>�	�A����Zf�;|OD��%�����Z
N�<�0�Dކf� ��\�3��'M"�	�R�.-K�A��^Ɣ����	"��\��-Pu�N�U .y�æ�s�D�Fxb���8��Y�✽+ ]�Ə]�of��B��
â�F
1㧉ZIj$+�A�p��`j��>�ԓϓp&Q�e�*2� ��b���S�i���6N'Y��W�"f�� W�q�#=�_w^VTb���@����R,jt�L��O�����L0���R�9Hja[1�0X�ˈ��O�e+�u���w�$��Fo��d�&՚�ȁmZR���y���,-��O�ܴT�0� ϋ�wk4��a��g�x���ڟi�n�y�NC!�?y��
�'�V�y��\�ɒom�Qy��S-Z��i0���3^-��{bk�9�?i���+|j�@�G���ug>��iCD��-o��2���]
I��0CD��m﮴l2u��T�xZc8&�0�lݍWB
��f���R�0u��k�>V�3ݬ���K���%}Zw5��,����Ҥ��5������Ȋv�(��$[�6���2Ꚏc��h�D.�[n"��7-Q4Pm���!����.�>S�d3}����DŦZ��e	Nؼ��i(	�l�V${N�q���P�	6v�}�B��a20�%IR�-Vj㞀xԅ���J���ʃ?oA��SVKq?���?	vΞ�2؊<��ḩ/�LP`�ɏW��9�*�q��h�2�8��.�͓���8'J@��%��S���p��
Q.�1�Ƭx��=���24p���:c`j͈��h���%�'F�����dȸ��J1Դ͓�I �y��>�����$�P7_�"h0eA�' A�Aw.O||��Ʉ%�#��x:H��鉜n����l@�d���%(�N?��'�������s��$��ux&/Y�"qp!.��|�nm����2͉'y���O?"�$�g�_N��$0�{���4VY`F��&jhYp$��P����Ot�ĒC?q�j����ᢃ�:��	�`1A�A�8� �:.>��t1ST���	�P�џ\�'�X���_!7����i��t��1e�=N�p�D�,\�H���5v��Vl�(E��b�]��N����O0�h�O�F�p ɍaG@hѦ�E�)uQP�'���M��Wu��K LQ�����nC�x�%�铞'�������ĥO���#�������H�,��ٴ)۟��bS'��3NN�cF�ǧ��_眝�Ä�6d��ˍ>���=�%�а[Zpj�гl4�{A�β4�-���Ǧ���"�H�[�N	�%��7�ABO��&����n��!9"*J:CY�7��//��0��
�c"����{��3����\?YU���&]��Se��hH2�A��L���j֍Kݦ��Y|(�xZc�<1���	4`%����%0؆i@I>�@��'�~�QGH��#&�.��2T?�s��7x��S�Eq���\����ă�"�~����_�r��JO�?[��b�M�eӡ� �d��]�?A(���ɝYt)"� @��mS���"_�z���U�S�mI�� W݉'���ٖF�.��S�H�u?֡��{�Ƌ3�p�#W&\%r�/�R�3G#?I�O�w���{7n�&n���HǬ�K�IV�yp�l��p�T��穜�6���cqȊ'Lvy	CG����'�<����d]�pn0x�pD�'���a��@���4��J��}���<����FEx�	��e�z�kG�
�\]�ȑ�|B���Oq�01�4���#=JV��#qL���#,Oz�80��/`��
�i&f�
��"438!0���#"�^	���6���3��	���>?Ad��'����ɕ�\B1���UMP�'W�X�,d�$%VX؟�	�n\	wJ��`�X$04�����2b~Hq�H<}�B �����ԀB�aW��*S���D���y ʗf�����R�+af	˗DƘ<�ZF���yBo&i�-��УҒ�6�Ǫ��d�0fD�D��`����)�'A����Ӌ>̝�'��)#��M�ȓpm�t��c��󡈉�5��$8N�H�O	#=���JN|�>�fc��}M���_�K���)��m؟<�3��m�ԴX��X�!!l����B�.�pqK�DU�%h���Is��} j�#(�ܸrlJ��(O��+��Y%ah|f�k��ݺv�O�n�k��h��� Q2�AV�B]!��H`d>a)f�E/T_�"DAǋ[��B��"6��A�IR�t��]�b?�JZL��0���n�H	�f�B�B䉠2���ahQ�w�`��I�[D	�%k�>�8w�Zܠ$2�|�2���[�=9��sw(н:JP��G؈`VV���I�BF��jծ|TxX�7a�� N�p�#�L����zN���5#�S�? �Eb�kV�CT*�Bv��4,�XA��7k�`a�� ǜ4G(UK���4�X�Ӻ�C�Y�s�F XGAS]�@��ˊ]�<)���'SV{0�T
@���hL�r�||0aMP�G�L�����%�S���6��=if�a��m�V֪-{T�HM�<If�(Kg8��v�8�l�(�'U�$֐��)����5�֮�R�'�8�DxR�Wv�@ٱ��	j��r��?�0>QwE��8m�*�#[nS�(�$���B����G|b�����u	�Lp�Z���R����hS��QR��Gx"B15pȻ�
	2�N��*�J"�S�>Sd5��du4r���lT�%�C�	���0�M�
�*x�h�FP�7�6&�Y%JL%O!l � Z����f55��\AKހ|��V��yb
^�2"\B�mR�6C��a�7(&��%+�$_&�i7,��XJp�����t��ȕ?�v̩B�"cV��[��9�O����ϓn_�d#Z��  C��Y�~&��Cc����d�u��>1� P{v�g%��"o�@�r��X�'��(
�N׾]��X$��;gP��'o&0̓���f��B�ܺXj���N������=j�j�ǂ�;D��A��7.�P!R�V� ��*��yAW����S��i�9z�"O�0���
�=�����E��RR���%�s~��{%�}#�C �����Z@�UX0��5<H!���o!�$�,�e@bh�*Rźu�H�]�A��)�O����P ��h1b�W�KL �W"OR�"����XY���0K���*0"O�A�a �9=���E�S�~��1"O�pQ�j>2��ec�e,h "O:4��o5��)�d�'G&ui"O��'�V�P�=1ѡ�6N���"O2���P�_�` ����;t�|���"O�Xq��@:ffAc�C��h���Z�"O,����0l�����N=X�["O�E��r�L���z��e��*}�<�w+N�w8�@�-�u���gg�v�<!V��������I]�8�k_q�<y��"}�4����=�$�Kp#k�<�!��&�����N�=T�T���*�A�<9dbZ"��HIB��J%4t�%/LI�<I���z��Qԉ=3�*�3aI�C�<��(:���	rWA:����@i�<9��Ta������3y�k KR�<I錶I2�i�B`~��Ќ�A�<������Pԥ�$�6L3Q!�f�<1Dϗ r��Ზ`ߊ;�n��� Yy�<)(S�\��U��Io��`�g��q�<1 h��EI���Ɣ�@SM�i�<����}9�т�*��d�R�a�<�7-���bWHY����JV�<�D��vƖta��h��1� ��y�/�0.�R�"���<��T�]��y��J�
��p�*P#*���0�I��y2	6k��jb!HYjH��Z��y��Q�QBT�u�<5�~<�Dǯ�yRiJ�N�ВW�\�:�V�	��I��y�$K�S��3��g"���FȞ��y̦'(S�n��R͉ۋ�y�/
/`l�Mq`�5:��H������y"���U�m�E��6-��ci���y")Ʊ-�Rua.��p����a㇢�y�#SW�`�9�E�m<zi8�o>�y���3���w��l��Y2h͠�y2K�b`��#	J�b76�q����y�G��x��4���XCn�`O�y�C�]Ԫh(q�!޾t{�c��y�$��7E����[�v���ג�ym��bE �6n
�^.�US'��+�y
� � Y*�m��djǨPA�I�q"OYp��gDJ���K,(�"Op�7�[�&|�[A�V�J����""O��x�P�6���0%)ǥ�RdS�"O��2l�9���z@g��6C$P�T"O\��,˞><�$�t��f1�1s!"O8T��,��XQ�%h46aY"O%x���K�P#�f���|a�"O�IɆ�ח]\lI�uO��
�L�3"O�9�%E�?	�8�;u%A�}��d0�"O.Բd*ƞs:�dsg/.k+�5�"O�Ib�]cx���n�,8���"O|�P���b����Ȫ ���p"O���*��^��!!�@9:5"Of��@F�I��ʹ=�q"O،!��+,n�sC��+ ꚝ�w"O��ڡ̘�TD
!����:@:J@+b"O�1���~����c )0��J�"O)A�@"LT�1k��L�0�msg"O���q�I�!��0@,��"O��ӆ�ʐ I��D8��tP�"O��� W�0�}a�	@�^0#�"O(����E&q⸔3+�4Mq�i[�"O� {�*�>����J]2��"O��2a��>�B�c*��X���t"O��D�].�bh+W���ڥ�"O�{��@
\}�t� ��17
X��"O���A)�m���Q'Tz�W�y��N�h1΄S7��*`}���1�΄�y�ʗ+eh�M9e�A�U�� �Q��y�#˵%�L�)6OF�K��;�y$ͻ��ႢG�V�ڜ11�
�yRP3R��s�Oں#���� J��y��c���K�ǅ�e"$�ŧ�y���#;���`U[&N�X��-�y� c4x��
C�E^tK��y�� 0 "(
��6��p���yNF
N�Ե{�P���O��yr�]+G��?�T����y"+L���y����;�b�Y�j���y*܉O�*�$����`�"۷�ybar�쓥)�%
�:%3��ҍ�y�R�xIh���τ���ҵ"�yB�B�(ڪ����#h���iT���y���%�h)E�#.'*`C4!)�yU� �sd�)(�R� ���y��زP!� T*ux=�C'^&�y�$��r-�u�Q���Fтn	��y2�[�.(�%��٧Z�,�'
�yrB�;�0��D�ܱ~��K2C���y���1O�*�KAo~!��ę��y���JJĈ��'S�FD�W��
�yB�_�B+0�R�+H�5I���Ë2�y���WԾ)3�l�/EBp��V택�y�.E._]�}P 7���&�P��y2��h,Z�b�'�a������yr���

x��I�V�XM�DF"�y�ȿy�L�Ď��P!TL3��y�K�;k�Z�z<�
ݳ�N�:�y"eˏZ��!����:��슆O]��y�#� �X���^	^��8��y򈙋b����@U�`���©E�y���	Y�����(Vż���dD��yB �2�f9�Q-BwF8 B��A&�y
� �x��˝�+�`�s���	
Zd�;O&�=E���.�6�K0�À,Ԡ�2���y���/X��b�[I�^m����y2E�tZ�4�,�������y�+a*��A��\��!�!��yң�$8ԨYS�@�@�A"�C�y�+� m ��rvc��
��l�P���yb�X.�1r�ޏ
���bQ���y�+��f�X���9k���"� �y�� v�(����:aB}y�ʈ?�y�Ȍ"i��Ы��
^��[p�_�yBĜ.9
h����� 9"���y҈Ƌ$uҼ��83�0��R5�y�FT!�h��vRܸ�'��y"L�J�:8wM���A!Fߞ�y��D"F��S��K6�����y2�Z�h�F�ϖ2���z���y�,�V�2��ҝ���hȜ�yB_"A�Q�RE��r�L��̂�y�g������G 	�o�2�y�&0�yCŢ&��=Q�d[�Z��P�B��y�)   ����@ė~[�X	��0�y"�H�cx����b��i�0J�9�y�R�v��p�/.��%0��B�y�݋�*3n-*�j�PM�y2��$-��qC�k�ځ�@j4�HO\���G�����ȈЙ %<�!�䊗o���)Y�o�)�oU>�!��50!����+�±��Oo�!�	~�ՀVoڃ_{�x�Q���E�!�K�%4�: ȅ�#x �{g
4rs!�D�"K�VX��Yf�aӦ"�s�!�ē�����!Ҩ(X$h�c�	E�!��"B�%#��>FP���]�~,���W�h�D��Sg��e���yrC7<j�]°e���p���k]4�yr�H&Df�H�NF2�n�C�@�PyR�Bl|���̶~�첥#�f�<)q��;I�X}���sn�"&��{�<ag�H(w��m>Q��áa��y2�M*p�� ���GHtY1�@.���_���O$����Vo��;���R���Z�'�p1�Ēq��A�ѵM�H�ʓ����v��=�<!!�Z���مȓe0��x�
�F�y��o���> ���,�q�S�t�$�](B0�X��7����2�_�dAP��4i������ȓ6��0��k�@��0����~e,�ȓC�<-j�E�%P��m:�&�jΞ���_�(E�ɜ&�L25	�}>dm��8���z$��)�nV^��(ȄX�]Z�|�Wf @)JH�� D���so�+&P\�i�&N��0��k?D���,���P���'{�Bt��)#D�H����"f�x�=	���`,D��P�Bգɶ ���ʦ$c
<�p$0D��2@�`��P��[� pЅ�/D�Ic�
?Y�h@D����Ҧ�3D�P�3W�Rk8#��;K^E�V�2D� ��d���<��㒕W�QQ�04�D0�C�[Ԕ�r�_�z�P�4H�]�<�����/p�Q�`�%.Q��j0ftX�$Dy"��z�$�Sׯ;B�-�C�%�yR	X(b�V ��D	�|e��S��y
� 8y I�hx:���
�p?�s�"Oz����F�(��X/N.Z�yW�iў"~n�/����Kd�|�8�I	R��C��6Jja�b���(�;v/@�}��C䉇t��#N
��v/�z?�B�I���*A�dc0�9�$�E��B�ɶV�|Ժ�Λ0?>���Z�s��B�Ɍ`Z@4c������|�)�.V;�B�E�D��h�\[mWϕwj➈��o�F`�ϗ>O�M��MV$>xC�ɕ�X, �ڧ�4 +�
�b�2C�5)hpp�K�/�(t��oIr�"C�	.]  qe&=O�Z]���T&�C�ɀf& `4Nμ	��D,���C�	$@qԄ�֥[�
&�]���O2��B�?	I�����H�{���jF"M11C��.")̉d�<�@���@�~��B�IHݔ)�!ǒ?(��6�D	Y�B�	�Ov�C��	�!��q�B3�&C�I�5�>|���19��ȶc����B�I�lv�PKĸQh����)�6d�х�R>�1@�_�c�p4;���3,Į)�ȓr��P��
9W@5C���he\���k�f���nݾY7��"]�v�f��ȓ%A�=˱��92xvÔ,���q�ȓ^��蓂��w���"f��_�t��rHL��O3���� 7�؇�L��tr&�����ADT�v��=��
}|��$��V
xEyX����_p�<a$Ã���)�,X<�̲���l�<�F�*5�ah2M�v�Ji���g�<�,�
	?�u��/v|�1��e�<���& H1�s��}|���H�<ɑFM�PfTuqe�o��!�`I�<��c��0�J�) !��27]I�*B{�<���!k�q��؂o�ФqtK�s�<����5fD��F(����kTp�<9����a�Q@�s�$�[Sj�m�<��i�%54�݁�	ԡ��1�F�T�<�i=G `�+�U�����[�<ᰢ�< ��L8�ǈ'���a�C�<�vC_�Md��֥ǱSq\iJ��C|�<�cH�!礩9�C
�"!@����@y�<ٖ�1�hzaD˧#I�XZ�D�t�<Qu!7l�
����<E�U��+�|�<dl�.&u���6��l�N�v�<�l\5B�ܬ2���}Z i�ū�Z�<���J�>�x�Ƈ��!�U�Y�<�p�	o~EgI�(as��U�<Y��٤`DD�����Zt3J�Q�<���ܨ6�n�� *	B�~��3�A�<���/7��i5%��A\�S�v�<Ywn�	?Ƒ�VES��+ +�p�<iaDK�>6hpd�_1h$RQI��AU�<�w�ˎx���B�܇-e��v��v�<��L0"��`H�@-]`�0�� Z�<Q�fV�n*��I�>w�MPbo|�<!4�/g�P��vhҶm؉[��Ux�<�Y�B�"��o�(i�l	=�!�'!���1N
�=��P� �&V�!���0>���0�N���N�1�!�D�V"��8E��p�02$n�@�!��*vD�rR0`s(�=`!�D4Jt�*�M0��p&�:NE!�� @a8$��Z��9�UB��f�"O� �i9Rez����3�D�  "O^Q����re��Ң)�3"O�	(E�	��ޜ���tL8�"OV]����R�qAq���OĠ��"O4�Ȣ�R.�<-�n��bV2p��"Odi�DŌ F3��5�Aj�UE"O�ɛS+�!�B��W��9�BPa"Oy�1��X��=�IY#d�Bd�"O.�	�+� ?Q:����,�t"O�����;@�,�Ɓ�5�F��q"Ob��/�9	�  
/ �x"O��@��ۨzЖu������g�!�Ċ�.v�,*Lϩ"����n_��!�{I�ܛb&W�'����Ҏ�.�!��@��H(�,7[��<�cΝ�7�!�dR0Ez� u��M~�Ф� \�!�d
$f jT�^X����9}!򤀉X��A8f$D@���U!�!��h|�����+Z�E �Ù�0�!򄀴#��]�p�4`h,���B��!�$�g~�|R�!Z4\_4 �EM�k�!�D��K`�!��ɀ�Je�)3R�ݔ#o!��
�hB�MI�I�DL���%>Y!�Dޟf���Q��%� <	�`�(E!�$��pA����/�/l�jd��DӘ4!��V�r� 0��D�<(�h��"_�h.!�Ė�Lt���v�H5k��5b��i��"O�䉂�GBO�`��Ɯ
��2"O��Q�씍Xa�ɋ��ȷD�q� "O����u�z�s �4�Ȁ�"OL�$ㅥ*Ǩ0��a�)Q��B""O�����G�dA/~&��4"O�=��֡D��%���!hh^��"O�yPV5G�B�3@�l2"EAG"O�@JƐ7��a
�� ��!��"O�����Ҳ?�d@Wm��N�Ri�C"O&��tƁ�J�
�׬فU��Q��"Od9U!Y�:=bՒ���7P��ٚ�"O@x!uO��O�X9�`j�D�.)��"O$e���	:����a���n�<�R�"O.�8�J&Q��]3	T� �H���"OJ�`Ԡ��b�N���H���HE�"O���l%J���Ǒ%�����"O䕁W'&.���"��;4�6�"O@uh�F�Y��%:� �2/9V4��"OD)�r/#j���[ň:[X9�2"O�T3�G�>}hv$EM-0�j�"O6X5cR��x�#A'21�e"Oy���F�'V\�	%��|�x�b�"OT]b���k|-�U I[{��&"OĈ�AE�#΀��H�*g?����"OD�3$��^�+Gh��E�*���"ONMbGı9��y��W�^�� �g"O���A(܃Ka� ��3Jf�ő"O�UB$�){2�ջ7��>,����"OФ�`��D�`�8���*r"OJU��I[
�ތ����+Pq��"O0Mp���!��ȱ��9��d�"OZ�8�H�RR����n�< �K�"O�kF䚳���t�Ga��8�"OPmXė�w�>�q[|�6�	U"O���Mݼ��q������*&"O0���0�T�+7b[�q�8��"O� lp����pYJ��q��l�P"O1Ȕ���B?ҡK��Z� �t%8U"Ov�`�%J?a!�� 5��P���ʆ"Ol� $�M�|lt���"q��@"O�a F4`�,x�M�F�d-��"Ol�(��<^7*�p�2��V�Y�<�5�:<�b%�I�T ��K�X�<i�"��~���|���r��U�<��H�Uz�I��)D����T�|�<�D��>
JvH�g�G�7�~-�3�{�<)t�������eҙv[�B��u�<Y櫓e~�ö��(�T-P��r�<�pF�-<�K��3=�H	J'�m�<�BBG/0�>=I���Pچ`�ˌe�<�4��F��(Aa���uo�{�<�d��0�4i �m�˂\Җ*Tw�<�@��,lB`:".��=�zң�N�<)��A�E�2E�C���9ҳ�d�<y�,�)wѺ=
Ѣ�""�}��D�c�<A�ɀf����`��gW(mA�Sc�<!�JL	�|m� +�Z9�}�f�NI�<i�M��[�̱�4a��R�}�QbF�<!B�� g�� �0�\�-7�xYa�@�<	�.�'�a���8Vd�w"��<)�ޓ��H˧F�\,�+� Us�<a���XTn F��uH����G�<)�ꏩf�D��m�w����uA@�<e���2t�)P댜{���U�Ky�<�@)Q?!>� h��АvG�0��b�t�<��cN�/��%s`g�3(��dڷ��t�<�S�Y�{a���N-4&q��g�p�<q��I� �>1�3�\�w���bF�k�<v��/�����"�Ųu��l�<�*� z������|��Y��	p�<91�1���s�,�R���ANQ�<q@�U�`.����<8�X�y��L�<)&��bV !��lմ0౹2aI�<QPDX�K�E��N׳!���Ӡ-D��gվWg6}S ��Ô�Y�`+D�4��!
W�BTN6R=��SA&D�l���8U>{aI%;Ϯj"�1D�����
���+��1D\���R�.D�\���HX�I	�.�,\�!u*O�l�3�>�8��-�+�R��"O���q�%�q[�	��Ce��@�"O|���U>^h��P��_%W}���"O��#�DO.s$�3�ɉ�G6��r"OlI����U�X��`�qj0y "O����C��\:H�	p��(���"O��P��+&�$P��лd���"OjL�S�f}0v��s���h�"O�Tj ]�81������=����s"O<��6F�r��i��
�+u���I�"O& ZH�
	� F����M��"O��`�d�'*������Gj� "Ol�2lܫ\�$#Q\�}	Dp�"O����@�.qL2x8E�/%>�"O����*�3 �$�� ���2UE��yb��:�"��W�b���Y��yB瓊(KF܁f.�o�f�h�!�8�yb-%C����A�A�:́��Z�yR�� 7l�C�`�0�z�H�cè�y�ㅘkF
��r�2��A�%�y��F1. M���@�_9��6 ��y
� ~�����a�8�BlΞ��e��"O0�S(�9U�������+Լ3�"Ohp��ϯHW$��QoK�j"I�"O���Уn\��c6�Y:'[���"On �cA��[{��s�c�3YP��"O�q(9e����e�ѣ"�V1ɱ"O�������� �_xx��"O^� �iƖ�!Sg`^fvj|yA"O,��f��o����c}2ap�"O���*�(S&�!E��	cla��"Od4P����9�"P���V�.=�؀4"OJ�R�J/D8u��+��3�>$��"O���F�ڈ=��0s
�[d (�"O�pߘ[��A7�'/,TL�׎3D����9Tx�D��k,8�g�#D��BB�ؙ?L�1aς�y�0�9�F4D�\�˗�n���`}d� �+5D�d���KzQ��%�)[�,ab0D���򄉫@�f�"�FA�>Eb%.D�(P��7U~D	cK_#-�q���0D� �u� BG�q���פ����.D��S?<}�I �JI�#���� � D�원�ɶ,�*s�	�=g���e�?D���@iY�|�b�Ѓ�0@�t�б/:D�t!�Ɏ%c���xT���0�X�-D��2d�;F�> �`�IB�K"F>D�`R���6M����x@��R�*D���tk�(Gt��,9TD ����'D��! ��!Cp�i�Hx� S&D���L��\�m�v��4�!qO$D��@U���^\��Cզx��S@L$D��z�I�N�1���,���+w� D�phU��r>��/� yՄ��7 D�����Q'2<ᇍ
�..p@�K:D�t�U�5\� �A�!�7%.(鐌8D�血k�?g�ҁ�P�1���7D��8�V#a����f�5(� �60D��C ���:n��*ڼO
<ɡ�-D�<��X�` �S�I׆K|�}H*D��җ�L�z��`��!}���%D������M���⁧.̎�b�L=D�L���0rL�)�6�@����b�:D��F��8dK���V!�X�b}��,D�l(4�f��!e��B@H�Hcm-D�,�,q$�J�	^,X]I�B�)D��㣒M~)��f�)>,D��GF+D�Ѓ��:7�(H�@O�$a�9�V.*D���6������dG�5�a��H&D�D�1$�
a~���VM-��s	$D����k�(_�rB�ܣS �h�4�"D����Ɋ�p_P�Xc�Llh0��,D��7����\�u���/��Q[`�+D�H�-��YM �`�	кG+$9G�*D��B��X�A,P-�ը���D���!4D����$.� ��̝rI,[Č?D�4���I�eP!�	 |� 6�)D�Dp�J	-��=�v�D�/Tp�x�G)D�,�Q@j��\B��C�WŘUK��<D��ɦIF`hV<��瞆J���֨ D��J�Ǆ�	�����L�0�$D�H2R��-;V��/L' �0е�#D�\��i՛q�pP�ռ|��D���-D��!�Ԧm�(�@���@g�E)���O�ĭ<���h�~�I*��� ӵ4�Z%��B^�#B�)� ���P�W,k��[�A?b��"O�)�¸za3���9�����"O����L�� /�#�6�p"O�٘�UR�8$E+�f"ON�A��͠R}H�y�Ν:X$-#�"OB��Є)tW�Ѐ ��OЈq�'4��`�)�&U�����Q$L�60�F���-`�TI
�'T�, Տ:h6b��&�A���	�'��Ѣ(SN�4�u��	*����'l 8�$f��v.�I�J1]x�h
�'��,y1�E�x t�&c�,*~��	�'#
e����&5b�
A��̈��Q+J8X��3N�h!�B��/k��0�ȓ)]� ��bZK�(��%���ȓ~�6Q��kӧ3^�a�ՏM4!�ȓ;+�@�'+��U��Qʠ
ъ	*̡��S}~��u.Y+{ơ��ݝ��ȓj��y��#&���`!���,;X�ȓa�n�SS���8N&�@B��TT��c��"�cK"��]0 /�1{"0��?q���~RC+�,�Ll�r��?oХ��H�<Y�"|4����;A�@�b�#N�<I hT3c�x��V��l/��sTGN�<��'�.;
��q����FOJ�<��c� ��B��� \����HO�<�%E��j����:_��4����E�<AUŐ�Q�4�RE�8Mt� C�`	y��L�I�:�|��C"��l��M���7~�]�ȓH0�p�+k r�����
vM�ȓ s.�q��EH��F �8^b���,���! ��@��L���,g8�	�ȓJ����5%�a���A�Q�"��ȓ{���3��eG�)E�͜W
i��Q���q�d����1�@|��I쟨ΓV�d<I3ߔw�bl��ŤQ�.E�ȓtaA�ӥ�M�&"�<��ņ�)�fѓhU.m����kG�J�@���*@���C����`#vO� %e�ȓ
jTy��w*Z|�#	�����ȓQ�p��e�D'$����g��IE�!�ȓxr8ly��6fuc�T8xOv8�Ɠf]*)�"��@� u���\��d"���?9�p(���F/_M�1.�����$�ʤ�x��b��+�vH�ȓ|d���dc��p���ތ��ȓ{��KՈʹ|b�R�f�`�ȓ3�LȚg�ٷ#�=�υ�~���ȓ���a&
�D�1�*�$o8t��D..e�.Q{:���*Q;��m�Iu<6O�/FҾ�)�oˀ+f~d��C�<Qb�	�5HRػDhٕU*^�sp�~�<ٴ��	$h$E VHP�ꜛ2"d�<Q�a�d�n@���5���S.Df�<y0�� �踋e�Hej� �Bc�<��-����qQ�AG+� d��E�<��g�mʆ�+��)^#(�˲I�x�<�ׄ�cOf|�3 T�WGx\k!��t�<9�'��$������6\�V�S�m�g�<�U`�{!�P�0^,����%ZY�<�'$ �w؎���&Ѩ _���@}�<�.��J�s7��n����.�yh<yd��7��s�KXcK"A��'H��aȟ�5�x���mO���' "$�ԧrzi���W)� ��S�? �y����U���7G�2���%"OH�[�fZ�\@�he@6r��"O@� N�jo�I�%*Y�vb��!q"Oh1���"�h𺃏�S]|� E"O�t���Y((��CA�?���qU"O =��N�@��1�R����
6"OL�c�K�Wh�Dh�S�dݨ��$"O܄@v��/�,�* :>��Y��"O �����g$��#�E?]& �"O��!�@Uvqh�d_/J�d"O*\H�8��؀!Ů�h�"O��s�i[P���π�nx��"O�q���%G�t������*d�8"O���JY�-�Œ�H�:�����"Oz��Ah�(5��j�l�##"O���i� d���a�b����"Oep��+�Ȍ���w��=`p"O~	 ��
E�||� �+����"O�Ĺ�MX/r�$A���>��T�	_�OӜ����0b�Rg�����"Ox���AM�n	�	ǣ!�TY[�"O�#�jJ�ocP�GT3	���8"O��z����M^1�c��'U���c�"O�,�wB��Up���b	�^wlZ1"OP��!�Ȩs>�$�`C%+it%�P"OF�w"B�A��`i21P�!X�"O����Og��'"#x0��!����y2G�*hKV)�K1l��p�j^��y�
��2�ܠ��ӌ{�I�F��y�`A� �X�d�׿:��R#̮�yriQYU�}	'ӊ4�(D	�	ل�y�kW)XdU���3��A���?�y�ϣ�<���`�#)��`Ҕ���y�(�/*����J�D�EkR<M�*B�I%J�9��S����A��qB�	�w��'�;O�|��CF
�sB��*7�.U�F���I�����`Ig��C�ɉ&%��H�& � ��u�$��(z��C�I2D�6�9ga˙hL�lrR��8s�C�*]�ʹۗo��K�9��9Z����7H���Plʲ	�$U� 
�f��ȓ;�%���ڽ{b�M)� �������]�q�Hx����:R�2D����d�9\��V!�+��H��,D�ȃ7F@H��*!�� Cu�*D�0�JH ����@f�wB&H
�'D�P8�N�-b�hLɁH�Z��%�)D���E�ҤT<2�	#���AA'D�l�G:d&�3�%
�;����N%D��Qr��!y� �C��Z�jrB`1�5D���E)��x�2hK �O�bX�� D��썀:t����2s�$�g D��(A��/H:�c#?6����D
=D�xʰ�[�Ax*���nƭ5���RG?D�:���$T�zB����|��8D�B��X�b\8��A��(N��c�;D��FH	A�ص��*�j��� �'D��R��[��}a��
�A��� �#D��գ�,o�R�"�(n+��Z0�"D�h3�	^���U�1m������H!D���!S�����CBJZ Y��!��0|�V��
:��@X�Cɣ`ɺ���m]C�<Ia�؊��0 ��F m�>�`F�G�<��#D�k4(��W�՟BI��0�H]�<� <��.NV;z���FQ���ʤ"O�}��m��e�`�hܱ��tK�"O�DIA䑀dJN����ְV�\�;"O`qB��V�mBjq �àsϼ��'��w��&2��`�OM�H��=�'���(��ڤU)p�`ŀ��o��z�'� s����m�(���D�����'?�,�p��^�({��4z���'k�]`��4G��!�Ҋ�;}*f���'s2�QjI�-��d��A�?��EC�'���I���i�0��b�;[�j�'n��3�<�������8^B�X�';B��$'�\�tH�I\8��=i�'��|K5)�<.b���|~���'�x�nKfB�8� gݜ~F܀�	�'D�4 (F�[4��eR�r̢Y�	�'�>Q�EK%��d���"`�![�'�����À MɪF�!�Y��'����!?I�� $�LP
�'|��Ql@#9;�ꕫ�*��'L�`�.�)k=H���2E�T��'���Q�� z�E���y8�Xi�'�����΍�?;2�A�ʻ%π��'��q
�囫e�X���/%�F���'E�gN�22d��!�C�:�8�'59Ӄ@���P���LG-?n��'��h�f�\�,@hIc��J�I�D[�'r�Q8@���C�lh�a��+}D	�'{������ }b���0��I
�'�|�Jy�T=h6Ӝ)�fD�	�'Mt��Tb��Xv:��4FĨS���''��h�BJ�|� u����٤�2	�'ĂI�*�4	´�]�H(��'��R���8��q��)"N���'d8���	=\`�$!��G7�R�'~�٢�/z:�y 4��-@�Y�'-�4���R��$e�L�`��	��'��̹u�
%u�~{tKΘR�`r�'E�󭀆h9����D0pP
��y�e��v2�Z��29�fT�C��/�y¦*�(�W�ļe7�1� �:�y��;b�<y��$aJ|t��(T*�y�HO��kE��*pJ^��֯�y�"H�j��!�dA�jG���pAF�yB�T
S�&��c@�4��I Ef	)�y�l��^3��`���-T����[��y��ͥ\Z��4��(=�!���ѧ�yb�@~��h�(߁8vE9f���y��(V�N�D���p�vX0C�y���J�jx�3�K�g�X0kͱ�yb�1i��;gGF`�0���d��yrLR�	W)��JCf���g���y2Cˢ�`9��ýVSʱ L�y��tB��۲�^�w��������yR̈�7��	9���o�� Xaϝ�y�IE&-��Ў	n˂�(�+5�ybOŉU�F�+W%��|�� �2���y��DW
ݓ��"h��PJ�W��y�D8R��;���4�ƱkB��/�y"��Y����A'~Tx�f�E�y��G��nyjCE5!Ɍ��G�6�yrdZ��ţ@�%wF\"u!�$�y2Ł%��tyD+H	jTχ��y2�N�z�lg/�d$!Ѳ֮�y
� ��酇�<A'�2Á��4��l(�"O�����G��r�Q����q�h�"O�%!�;��D0�c�!�
�"O,��C�Y�{�)3��U<7�����"Ot��#�N�(�.e��a0 �r�P�"O�yv�ɡN���n�`)7"O��0�5A�*<��T2����A"O�L�!#^�P�B��4V;l�"Ol}�TB�a�n̓b�8[�`*e"Oz�Se��=GA:��5L�<U���"O �!�o���5AG��8+�"O:T���,���v�Q�J�
��S"OF����Ͽe��HCf]�R�H""O��Kw�L�I~}XFN�d�*-K!"Ot��I	`a�4H�2[��
C*O(��0�:��H�OHJP���'`�hg/�8
��Y����/HP�� �'�j�+G����A�P�B�C�'�xy`U��k�����Ől	�	�'�"�33�հ���[G
"����'��<���'?z�� Q����'��1!��YjQE�� !.��'!<Ԑnض$�h��N��M,ʨ�'h8�/� �P�1gm�FM���'������E9'����T9Q6�{�'�,�ɛ�y��r��Җ0��T)�'�lX��/_u�}b���%ߒ 
�'ʨmh�.� 8O��p�B�KC	�'ǖDb��:��� ���3�t��'�T8ڱ� &_��$; ���d$�R
�'lr�iG��:L��S�aS*悵��'2,R!�:)��U���¼t��a�	�'ȼ á �>T	��&�֖���y	�'���ƏO�6���U@/�(��'�HhK���ujh9b�cR�x��
�'⪐S�Iݫ���	Ȟ]:�}r	�'�<qe!�!��5('��l^���'����!lT��g�A�;�D�'X��4(�5%ҽ�A؜rYn��'�^����W2�:�]�7(D�K	�'8��Wh	�tE,d��]?2�^!�'�Ҽ��l�8G��]�F�Z�6\���
�'�j��F̴[��Ě��j�I��'��؋ ���&� &����\�
�'(�M�w��Er�� ��u�T�+
�'���qȊ.j�8Ї)�X$>c	�'��b�g�p�F.�#y�r��'���k�h_(�P�!���$��0`�'�)2�ɥN���V֒K��S�'��49��͝!���Ʀ'�XL[�'�T1�LV�w�TDх�<Z���'S:���o��#��֦nux��'��Y��E+��;���2xv�+�'��3 �՗����T�Y�&<���'�(	R��$4>u��ӦWh��
�'H�q#��D����o�fXy	�'6ZH)�#�#l� �@�K< L
�'�M�d�Z�ۡkXl����'��A���3U�Q�`�)ed�)b�'<P=���,.��c�mR8a�<Q����y�K�>D����fY� �5��%�y�kYf*�x��ʘfA�d)�I��y�^Y��$zb���0�:��R��y���Y��3Ň�%"3��P/�y
� �`���ږl�a����-+���	�"O�PY!o�5f)p�ja��1�ֈf"O��� �:ְ3s��*2�f�9�"Oޝ���?L誔�@A ��D,�0"O��E��VDX� c ܔ+�8��"Ol|�7�	g$R�Y���X�\���"Ot�&�?M���b�I۵�6hp"OԀ�#�# E�����4k��TAb"O0�ya��	-l�w �Xal]��"O�9;JL,}�����A)j8Y #"O��,��\'h��bOB.L��"O�1"M[K~j3���+�Ґ;�"O\�T�٢M�����d��^��u�%"O�F�p��iD�M�M�P��"OvlAP��"��Y u%G���sE"O����g��b���C>�pIW"OT���K�Р�W�ԋ�LX)��'���܃[��%��!;&DC�a_��!�D�'E� U�J�7\Π ��̵�!�D�#>z,��4�ؚ>�u2��z`!�$]&,\z�p#��qDR�m�*8!�ܷh�����C'�4U93�-!��w6����=%m\4 a	��~(��)�
"0X��� y��M�%N��:Y��3�'Ȅ�W��h_��TǮ0�
��?��yrn�	E�)['���F��< �"J��yr�ק0�$H��� 90D���&
��y�)�z��\��л-)�9P�
-�yr��*��A���(zu�]���
)�yљT���$�?�֘�p�<�y�V�Wq��X'a�"����+�y��.�*�l��2�Jտ�y%K%O:]�wO� ]�!u�]!�y2々~�ZQsg�
�8�t��?�y⁂o�@����0,� ���B��y2�L�w����'��&�<Vg�y�*�~Ȯ!{���Y��bGM(��'�ў�|�_�}��!A���%i,ܘC\�<���[8�J1ۄ�Ϻ?9�ŰNVT�<�f)��Z�\M� `�9]�(r��H�<!��-|<Ѳ��2#ϾK1E�<�ҡt���"�,>��Zb�A�<��B��ga�ԁ�F]9�)
��s�<�t#�>�C��4�0x�3kG��h���O�R  �.�c�T�c�{�̂�'�r����N�Jo�ġ���|x���'�&��b�B�V��(�����	t�"�'�@��	.}���{A!C��H�r�'�5�!�O9^)��� -q�'-��`�ˇ_���� z&dY��'e*u K�z�r�2�g�6��Y���'��'�B��K�Z���8W���5�`¦	7j��Od��DC^b�sFŗ�h�\���_�EϚ��&���Ѕt �3���s�A�p�+D�����֗A���h��ŴD_K�AG!���ɬ�q�^�*�&ŉ�L؄T*!�d�,DT��G\�6zF�ȥ�јl�!�D�w�NmY��ͣX^L�Sv)��+�!򤆚D�V��H�R��I�����!�$	�i�<Q��'���Nй�w�џ��?ɝO<,��c��V�͙�JĬS<x����1�O*�قI��`Ԏ�Ї�C����"O�h���U�%��^*v׆P �"O��Z�Zd=����@[�e6��bw"O� d1	P��Sn�+v�A+o`Aض�|��i>��'���j�/��|(�F(��&L�ȓ:���r��=������źm�^�z�'�f�R�/��6)��-J�fw(t�ϓ�?�yR(ܿe9T��%K�?M\bh�E*��y"L�3x�<� ,My8��N�y��A�8�nɨse3��������?��'�^�26%�%{�18��6�u���Oڣ=E���� ?/�!�#��e��T�Ӂ��/�!�$H�t�~���B F�\����&Y�џ��'��I�|�T��R~�|jתL�i���k�-S����?���ވ���҇B(|ܰ����ao��"O�CuD�9CІ�Kg*D�:Zd�� "Oh���F�%�$���9F�{�"O� Ҕ@ �.A�S���, q�"O0��L;��©�}"p�"O(䘰��	u�əG	аY	�5��"O�i����,��&��e�.Q��	ß�G�J��6ELSdd�s-|݃D�-�y�e�1�����]5n4��R�n���y��E�v��a�P���f�� ���ׯ�y�ˆ�6��4
T-g�&�C
��y�͖���sR��c���ߋ�y���i��qz��4�b3��O"���$y>����E0'&b�����:�K��O���0>�SR�0�FAْ�	l���4BA^�<ɥg���3g�İ{<^�4l�s�<�&�9�ܐs�@ί+m>���NI�<��ܤT��`���(k����F�<9Vg\<T��gd���.�Ly��)ʧ"�J�G�d�1B�hF	j0�ȓ
H0dE���Ie����ȓMJ����=�&��W�'`��(�ȓum�)#D(YjT8��@+��#}��w$��c?@Fl�h�ƍ/D�tل�:�MK��R�x�rˈ+s���������������z��}X�bU�8\T�Abƣ<�����(�d��J³e;�6
�p| �!��'���<YM�@B�
"�R��0����ҟԕ'�a|�d��tY���8+����]��y�n1$GQ
����6��E��.B5�yISo�)b!oP'5����  �yrL���(1a�A�/ۊl#E����hO��O<�IdC`Y"H�74lE��VyD����d=��I
`u{geM�N�Dy�c͑�D �B�I������,FJP��O� o��C�I�y��E��Q�f�S�'NT�B�	�wwz��`�H�8ZJ�
f&�	l!��^�q��`Hr�G8�%a'#��ig!�Dm�$��V�ҿ4!�" A%75���h@�i�g�.��y)-��KHB�I>M��8�'O��X�!�!:Ad�?!(O
���ԮIKt-�!ʊh]V0)w�[$�?)��?��b����ah����Y��-��q����F�����[�5�x���2F�:y��F��9�l *r�m��m�	]й�ȓN��%�a'LUy�g%��D5�0�'p�	v����;��<1���9d,�F��$0H;���'b���5t�պ��R�,�6�A�'}����L�
ф�)VM/0��=)O����D�o��y��oόw�q�����n!�Hid,Y��N�!����.^t!�d��r�f�`!��
F,}8��-a����"x`�+��Ǧ�@�hH<��B�)� Ԩ��C�v� 방���q�q"O����bӯC�8�	��RaP"O�Y	�m˚'��AC��
uB3��'	�h�T�J���tk���NE|/?!��2Z�trw�"uqV��b[�/!�D�>�0�p�	I
���1� ׍t�!�D��"���q�J��m�f�b�)u�!��	!W�dD���F1���*�K+kD!򤕋N/���f�+I5�M�䎺(!��(�lp*&/Ǚu6��ףO�&�y��	�t�~��W-� $U2�`���7�rB�I�`��%�5<^H����U?XB�I4X��H�e�Ә`$�1bق��B䉙F�C@�q"�m 5�..TB�I��.���#�?bl=�P�ױLq�B�	e�f1Q�&(!�����$n�$�$'����GH�Fy�͑� �5M�x�1�+�숟�!��]����B �43��̩�"Ox���^#Wt9���Z�di���"OxՃEb[.F�13櫞KO~4�"OJH��� w�I딶M>ąc�'�ў$G{�O�/T��u@ӛn��ћ�B��o��'ў�>=�Ct:�hR��� R��>D��4i�#1�S�JL>:�*#f=D�p;p��
-����/I2B��AS'-D���6��+$hp*��0"�=`�*D��R��I�DP�)*��)D����	ƪ7p��)��M=.標���'D�T2Db��y}�R��#�څ:�&D�X�w�Hg�5��CC$2t�ە�0D���0/Y&lFqPE��%P��Q� �/|Oc� �j� F )v�[��Z��,D��BC�L�)�,(b£!8Dt��H%D�D��i�h�R�R@K���R�e/D�,��']8β�������"�12�/D� �p�[��> rĥU�L�(���,D���ũX<f����G_7�ح��,D�T��m�� �Gh3\� %�=D�8(�M�z�¬°�/)����C;D��@�/�qT>��/`K�8;t�7D�T1����X;�]��'ۤU�x�{�*5D�t��"�3�N�U�ڷǆ`��,�Oȣ=E��Ǟ�.	�u;G?1���ECɺ<���1�g?�ǏCsQ��QWx�p�DIa�<
�a�N9y�FK:@�A�G�gx����d̓d���耯�2rָ��f��)z.��ȓ	;h�vHX>a��Q
�bG4@;L���'A�蠐�ѡ&����a!�0V�tt�ȓ-��(2[�!�¨��"Y/>ɾ|��.�؁f��Q+�y�%�� :!6��I��h�?�O1Oj���V!��Z���hL�hb"O:	tI�
�@h)UC�w7.����՟�'Y1�����¼�~��SÏ+8��`��"O2�B!�*7����W�hknъ�"O��p�&	���(y�m4aLȌ��"Ox�L&2�: Rv�PGKf���'�!��'h�,[�C�Qq<3�ŝ�b�ў4�� r&����W�=��;��M�+��0G{J?�#� ���%��;!�����9����4§N��P�HQ��`0p� L��Ԇȓ/o �².�+z�H@�N�?
2�ȓ=���8�Ń�ܬ�����m�ȓ#�B��G�c6��X��|�Z����z���f��*�8vCĒ�H��S�? *��r�W�D@��Q�%#>YPU"O�q�C�ŭhT��@��D�N���"O��V�R^�0�uAQcj���"O �� �,��C�:\�u�"O�Yq'��������ίvG����"O����"U�	�V8�)��D��l��"Obs�W�)P�����ݙ^����"O��#섬-��0��^2 d�pZ�"O��`F�I1L8 �S4pX`�0�"O��:qCB��VDP®ĭ%;ʙCe"O��ʗ��(l̘��'-Ô=֠:�"O��������v���{0T��u"O�p���N�v	��[ i ��`�"Ot��bOt~�;R��&s}�m{p"O�U93���*Р`��ɐ��'"O��M^� �B���_�b^�I&"O��� �E�$����h���5��"O2������xL�vHH�۠9�Q"O� �J��(Τ9h׍��m�h6�3D�Hi��@)J;~�R���8�h٣�e2D�dRƌ/jK֝��S�a`u�e�#D�<����U
dl#��1ST�2�� D���e���A3a�M�D�0����=D�t Ӣ�T�JxǧK�	��㒊&D�D�an��wDN��A����-i$!�DҊ|{T�eƋ�^"
��T�7�!�dȭ<����W�5���'�Z;[E!�$ݦM���z1��d�� ֌�aA!���4c1���Ä�Kw�8wC�U!��ư�J�2��+:if@�Q�@�f!!���.،�	"�S<p���E�!��|Y����ei�-c� �^�!�$�2G�f��c��%([�lqv��r�!�d�t�8�a�Y�GBx�b �`�!���[5��Fm�H�RC�W!�D��`.�}Ô��7�r4���!�r���J����, �,�G��fp!�$�?/����B�Dv�2AC�E[!�DV*95pQzҭ�D�
�
���tP!��9hp�9D��M[L�`dJ��-7!�լ`������9h��%��L!!򄋺,Z�۞a8Ȁa�f\��!�
!K�\��C�4X��iq���g�!�D��,�������l�uBʃ#�!�d�-@2䁏� l�I��i!�\�
Ȃ��*l����# �(�!��/Yuh��ph%o���ĕJ�!�dM�0��E �!��]�����0�!򤝄FN|�U%N
D骽��C �!��4}���-Ϛ4��a��P:!��ףI((T��P�6�P�Q���d!򄗣<̒���X`�%@�bX"S�!�$���"l��ʗo'��w"�!�D�
	o �����X ��`�қLv!�đ�e�(�3�n2s�t���ɜv!�Ĉ-\m.�*r��i��Ɂ���3!�D�A����Dըc� (��d�!�D���`%��$ɋ6(T$�7�@E!�d�**[�0'��{ X�H��R�!�$�:����ݖ9!�b��V��!��'�J m��}��8 @�E�D$!�Dމ#��$J��W�?�D��3��Y!򄃵DxmZp��N*�\���!.�!򤞍B�0"e�4C��PR�-C�!�� ]��K̝k(��iQ�L�cѪ8��"OP�U�xf�*F�_�Z�D��E"O���U�0������;ߖ9�"OH9Y��8���[�@�(ljd"OҰ+�
-v�����L/� �X`"O�qш��#(�U��eQe��:�"OFt��D=[���Qy\��X�"O�J�M._):(�veZ1�� d"O4�F� ƍ���P�,��"OB�Jvˀ8n$�[q�D�6@Hh��"OB��Vކn�Vq��+��u�@"OحY��Հ2:0����T|\I#6"OBQP�
1k�2���� $R��4"O�B��]�E]���F��dL���"O܈BEM-j��M���3�|@#"ON!3b�
�/�>�u�ɷ=��`5"O�d�gi�(0�P�P�.ˢK��:�"O���.ˈQ�6l��V�D�A�"O�qY�� �b�(�fbO+~}L�"O���3L\�Z���a�R8.N�AX3"O�D����T�: sGnL ����"O�� �RA��E����X ��"O�m�a�
��u�%��6m��(�"O�k@�CZ��x&bB�ƀ+�"O�D[B��/����眪 ��#"O�8KD@?��)��oš��؋�"OB��U��2R���`�g3{0���G"O��'��]�xA
�f��,��{u"ORɀ�՚;�`(xv�Z�^j�+�"O���	�)E׮�k��N�=[2"OD���|N%SF�TH��&"OF����ܽB�e���í��EZ"OXu:D���J�@M���S��zX"O��!��_�ޝ�3&^�|АdI�"OH�6ѥJ�beXV�7S��Ac"O�<�0�^�)�*@�S�� o����"O�e��Çi!�I
4f�&]3���"O@��q) k����cgȕ_�H�0"O�QBA���y�4l�i4l4"O�Y��A�5�.؛�h(���"O@��J;x<bE�t��l
dX�"O��s�-�k�&-9���)z�&y�g"O�Q�F@���D�W#�����&"O�It�š~��ɪ$�W�[q�%�3"O%;h	G�t���G�nm�R�"OXS�P)�p��&�2a����"O���#�lKH�:��!4U��V"O��0Vo^�n�Y1
�CP`H�""O@
� *Ym�mB�T�'#f)C�"O���Z�2�DZ�/�!M.�:"O��Q�C��?̀�r���b]�uAa"OB9��*�u0���E6F5�<��"O�t��	 %a��QF>D�,r�"O�A���x,�	"�_�=d���"O&��s&Q�h � ��훦a�Z�P4"O2h9@㏇k0h�qslW�+QB�Ȧ"OԤە��0$��+�EN�!@$!3$"O:P���{�\��V��k#"Of�ۣA�"	Zހ@�	ʏ_�4���"Od�9�/3W�Vda�g��79k�"O*T��l��W��L� ���>>yQ"O����L:j�ܽk2%PNӴ�["O&M2�J �e ي�� }�`"O��������ӗ��"�4"O� 4��A�]�RdK��_s�0D�B"O��v(<{�l��F!�_� �"OR���J��g]�2� O�J��(�a"O���/\+��C�f�0
�왠"O��8Gb_��QY�%J�C�h��c"Of�C�X4Q(�M�c�T#�t]P�"Or-�0ǒ���hc ��N��ˁ"O@���¹.��1��Һ��xx5"O����!�/�4��C"G7V����"O��HӣU>,�P�rhZ�;tt!�"OP�J��:)S��ͫT80�%"ONT���U���+���Z��ĳ'"On=�jJf5��-Ӓ9��5�0"OȘ�6ME�r��SnQ��8�"O4E
�!�.�� ���I"L58C"O��-��?
2h(T)��H�Ȣ5"O��9�G�!�6�Ic�6k�έ;�"O���/�>�"��Аp东y�"O�	"�h͑iB�l⑃߇0θ���"OxDge�2->X%�C\9#�0,��"ODy�gE���!ʆ _z�P3"O��!e �#Y��2k/'֕I�"O,}ړ�q�ʱ�� V�11T��W"O����a��%�-���
�;�T,�T"Ol�Q��#(�>��($~Z�'"Oʴ���
K���a��޻wNNt#e"O���B���.5��J���"�J��A"Ox��vjH|Ԭ���fO�R�2�"O��+ P@:QРE���ͨ�"O��n�!$�!�
+8`���"OYK )�13B�#�hF�p_T��"OFYI+�_�a�WG��X� �"O��Ňܜg���C%M��p"O�q���EO$�q�"a�p�V"O8 Q�Nʗ�8����_V4�D"O<���@.���s�۽r^�0"d"O�5� ��&�6��D�� NN"O����/ǵ[Vr+ς�dT4�x�"ObE�߸}d�X�S+�<i�G"OD�qd	��<ז�
�靍a+ry)e"On-b�&��c=�,BԨ];^	�"OJ`	��,m�ԉ�	|� ��q"Or�sr[X����I(H�0�80"O���/N�!��@��;���Ҥ"O�,���[��U{&O۴1�� �7"O�����A�v�
�gȻ_�$�&"O��k��!j5���_��)"O����E��Y��]Q�F�C�J]"O��*`�Ը���f�W c�lD�f"O��ש����b!��Q����"Oz�R���y�$�h^b�1"ON�r�ǀ;oHt�dC��X�l��"O���s�Y
/�4{�A
�I�д��"O(���>G�h��c�D�j^��"Oʸ�#c�;"��sq�����I��"O��J����]K�H�4m'[�,�t"O8(���@)��
�����"O  ��->K��Tq~Ȱ�"ON�{�`O�mC�i��E�}�b���"O�}� ؝Xe0)�рF3G���a"O�$f!Ziv��q��E��5(�"O��2V�
6˼(�GD� R���"Oޜ�@`l!'��4.����"O*hAU^�)j���.Vvh$#�"O� �[L՜*�64���gc���"O^0:�LO�H��E��*�\"�[&"O�Qk��ԍPr����+�*,�"O&��aM7�=ڢJ�I��7"O����oW�
8��Ǵn.�|U"OȔɇ��k�����H*�K�"O��c�R2{�H([bĀYr���*O�1h��Q�~���Id�*����'��TZ���O��+U�J��h�z�'�i����x�Az��V&�x8��'���c倕${읪 ��@o�<#�'��]2w'��U��z��I�"�����'�v@�"�P���gb�jLݰ�'v� ��`�$�<�WO�9� ��'�.aҊM �240����:�,Q�'���Cd��u�A��ά5&y��'�
u��i��,��i5Iܲ&S�!3�'���H�JI����e�U~&]��'L��e'$C�J$�5[J�
�'&��!Ώ
M �38P�
�'���;/TB�<u���.,�$p	�'n�P�VC�$4, 1���\�0��!	�'����V�vgZ*2i�t����'� �Ń��!������l��'���9�J��sfع��U'sn���'���
V͏�Jw� ;�埈x��	�'���u��3AЮ}���Q�{d�i�'X)��o	�w+�p��K�*��9�'P`�����A�D1e�ۻ��		�'GL	��� �^�$j� (P¸�'˒}sE#�R\,�s"CJ-.LB�'��!��ոv14�"�+īXn��P�'g���E,܊c��#����'�A�&bPA` ��!���xk�'\��`\8 �$�ʆ傊I2u��'�ܹm,3�h`!��-����"O���!��uY�l�`�VI^ny�t"Op)p�@_ m�`���Ή+K��"O���g��-UT	���[H�DS�"O�"��R�&�,��A�j���J�"Oՙ�O
`rD��"ӓFW88�"O���$ ��_|�Dk�Ꞁ(8HD$"O�M`�$۰T)��c��( >���"O��3�o�&e]ʼI7�Y�\�!���,�S�IAB�Ái9	�*�aT/�14�xr�&0�z�c���+<`�Qs��ݫ�B�	�0��x t�H5���:/H�3��C�I�� �R�������#�P �C�I>�!�m�1&�^X�f����lC��u�,����"�0`!�oڅHXC䉬[l��q�'%$Hz� ��[LVC�\�8���#0.Ȝ�ၜ��B�	6:�����ǁ<U�aKZ8w�B�	
��d8�B�W��ؒuN��NB�I;w[ mYS� $I��
EkL!xW8B�	' �\�r	��'hB�``��{�B�� ���'�n�2���-�u�B�Ix�x@�@.�Y�H�6rB�I�k����aD�q��D�ʒ�x.�C�ɿ{l~a�Q��� �X�E�&����X�C (������J$-���	��!�d�M/�dr���=϶�{��� �!��;�n�����("ıc�e�Xu!���7��l7�җh�(psę�C!�� �� d!�/B,��J:�6�Â"O�)�E�I*�6h���I � P "O�5�Y�%-�B�xL�"O�� ��$� $�B�]'����"O0a���*��]ءK�"ڸf�!��8�J�,x�܁B��Wh!��+��Hr�"�h���J�\!�$S�m�Ȅ	!  b�a"�ފKE!�D�ڒa��;]V����)sA��*�'p�q`f�Ȼ��Mj�3����'�"�H�o�v�ŅФJt��''*]�P�T8U���sG,^7p����'s�,S���!" ��)�k�_$��'7Ʃ��S�1���]Z��)	�'`ؔ0Uy� �V��)Uk�\Y�'B6hԡ�5�0����ЊUg<l��'R<�b�JG�����E����'H44���*f��
E#��F((��'ꪡI���:�@��4�ΙS�Z]Z�'�l���t*y���ȮK�4iX�'�f�7��,���[r�R/,����'8���@P������'WvB `�'f��x�ڴh��9�gӁ_�����'~��ؕ��q0N�҆�PQJ��J�'{�A�HK5�ޅ*��[�N�Z(
�'����S�ݓM���*��D�!��'�|��ĢUh,H��W9�R���'����'iH2��sr��3wڀ���~re@O�eZ!�G�X\Tc��J��y��i<�5�pǥ$5�k�Ę��y�b�F (t�ȋ"���!��y2��6�@Rs��/�1���yb���l49�0��(V)�f���y���t�3�ȿt���O���y���$����r��\�:��M�yG�=Q�fIC��
c~��@���yr�R䱠3HY(\��H�	
?�yb��;��jTJ�N_���Y7�C��jCd��-P�&�mCRnU�F pB�ɖV�b�
�;5�Q:�g�MC䉔dT�8Ԯ�3�}C)S�0g�B�I?/������� D.GC�B�ɸl�q0v�B�N�Yv��D�PC䉮q�^!*�MHE>���4�B'Z�0C�I�<�li�r"�$2����g¹dk^B�	#شP��Ï}^!��J�-_A�C䉜O�lE�dH�Fɳ �݊*�C�ɴK��e�!��<LYᬞZZC䉘5B8X��nN�Z�ĉ�q�\�� �����쩖���k^��%���u����y�dϊxV�$�f������*�e�`�<�`'�,j��&���I�#OB�<i� O�a�|@�ե�l9�eȰ`�{�<��.%S��1���R�`8�V@�<1��G�E�.$�r��y=Hu�l�y�<!��W�b�:d�/��Mh$�m�<	�AW�$��V�U_Y�cDl�^�<��N�����l?i�K�*�[�<�D%\�[�\�ꖤ����0���r�<!�� Xz����oL�H��ր[G�<� %	4Z]�D���Ϧ�����}�<���C{*�b�G#I�T��d�<Ъ����)P��H���Q�b�<��LMW�!I1.[�"?�\��)@a�<� �I�����~�2��&j�m8�"O���NR�u�$@��!��#"O:\ᖉ
�Vʏ�
�bg"O|M[K yc�و�C�Y,�h��"O����n�|�� ���X="���5"O6����P1L�>8rA-ض"O.����R�2��]�c�e |8�"O)�QB�2˘�u�ۂ;�f��"O�Ez�lS"%��q��Үe����"O�����ٖ7�T���6C��X�"O����g��+��`� �8k��9A�"O�ҡ ��7`�q�0	���$ܫ�"O}:���q\��eiϭ��y
s"O���@O�&J�̓��K�j� "O�m���u���H�̖0f�dW"O\��׏Y�$��zaL��.��"O��r�Gݕ;  y�Df@�(7���7"O����2�u�BK	U��p�B"O�Ъ��D��lYBŎ�[�̸Qf"O�=�r-�8YXlؑ�T�<����"O���OB)NX��u1X��e"O:� k��$���T�W�W/,�E"OD����X
D}��^J���x�"O�4��� �$ѥ��3>P�!�"O>��l�l$�	0ѡT ���"OJ�"�=p����� �D
:Q1�"OR��%V�0��m�r �2��m*"Ojh{�չ}����$�ρĨĉA"O�@�Ɔ!j92Q ���s�ذ�E"O���"8,�[�
��,���i�"O��q�lՕ1�tؘ3
]r����"O�t� �OԨ`�	�&�l1�"O�p�EU�Y.�:�n̑�6U�7"O�Lh�����e�-�� � W"OJ�#��Ơ� %�w�H%-nX���"O>�r�d@�Q���0�^�
2��"O����7d���kň;2��T��"O�0C��%�l��$Y<F��x�"Or%��ѓJ�V9CߦI�,��"O�9�ǣ1Lv��e�B��ԋ$"O�,�0aF���%�
�`s"ON�����7rZ1���V�v ��D"O�T["(تF��{�aQ_�ju��*O`y��	 x�எ�b��I�'�l�#�Ȋ�Lt��,L�Z����'�4��睛A��B�K%<x���'+
�x��O�g3b��H�����<���� �I$h� ]̜��(��<���C�X0�5,��,��*�V�'���"V>n����o9~)��'o��2�m�XW�%#p�� \G.PS�'^�/R$C��0; � �S�^���'���b'/\�� ʂ	[�R�{�'��!�%��q(��r�6UK�'�f���N ��B&X�WV�ő�'��8��+7$��2�c�+q�t2�'-j��5�ټ2C���� �;iT�9
�'|�����Y�\���҆O�	�a�	�',@����C�P��)A�lI#�@�
�'洞��+�%ݜ��H������'�B-�@�=�&�;B�[=-����'T�x�7�K�n�&��f�!:��y�'A�A��8
�F�q�����R
�'�l��m�w[��k��K�c� {	�'��1�珴T��)c���vP ���� ��Ӡ#Qɞ��E��<���"O�躖��2s����oG!E�(��"O��th�J�X� M"Z���p�"Oxԓ�BO�8<�Ç�?$��d"Oz�����ä�(0�y4 ��"O��� �	�,�rIԎMD��b�"O�Tط'��~����.XB���"O$��V�=梅��j��xMhhx�"O�tcR�D�lZ���>�ޅKg"O4��NŵV�0�稛����"O�p���z�N�#�gÖ��|
�"OTMa7��<Լѹ�Jy���ӧ"O�u��a��H_L ��+�:^��$��"O�@J
i����áb+!��O!Q٬�Y�N��cp���/!�$9YB�9vL�~S5;�*]!���D#]�ge��@�$s���I�!��ɳFtJ��r
H�8�X��QD=#!�$�-]�&���.�H)\ɸ1�~!�DZ�k�h�ڐ�ݤ���F;7�!��!Ԓq'�G��ấ`��PyrᆤF�F���$_>2�(ɗ��7�y��;-tx�h����7���ؗ%��yR��W�P��NX�S�Y�e���yrG���d�'��pC��S ��yB,J!
�╫�G�pn^���`J	�y�� 
��	��n��r�"��b٘�y��ևr���F�1[j`p��F��y"e�P��@2U�L8-c�2M���y�
t'N�1�خ�lyr �y��˘gA�pId�Q=��Є7�y�a��Tn2�`�� 7fE���W;�y���M�!J��D(�6i�a�
���7�OR��*s$�h���B��2�a~�W��Љ�9(��%�w��%S�`����9D����h��W��)��-�C�P�5�����aW��O�D�N�of\�!"O�<�Մx�KR<iۚ`�Wo ��y��)�0�Y�������`�ڵ �����d���wJ[�w���l�B�0��'4�}B�8~�%"�OE�E���0�F��yrM�(MZV���K���9����y"F
>PY)e"ʤEUD�K�K���y2.�%N����8nc����i��y��;%�bű��\D^�jGψ��y�&1]FJ�s�O�Ec����'Z�y��G�t�2��\&d`�����yRC+u,YJqF[8W8����HU��y�i3qʪu��HJ�W@�9����y��D<�@x�� �?Վ��q�ِ�y�O[*q%���4�%ї&�?�y��ʒ&���0B��L�[�I���y2�Ȯ�����c�X|u{�-�%�y��ݟ���Qq	F��DXf-A��y�B�?~`5�n��x LP�բą,�	;-�� a֋X�g�'C�a	����u���$��-]w�|#�[���v �-"(UQ�! ����W�>��`��4f���&J�(@��~�@ӭ��b��1Dy�j��%L�D��
�x�P���\�$nڤ}��u��D)�R����(�y�܇G<����u�f�����:��u`t���;�Hr��V h8N!��sޕ2�M:-���DM^cF^���H/D��:�C:�h����A���UD��aR>�PF�O�Y(�h�![@����:�HO<����7da;��rH⠒d�'&Rȫ�	�V�`0@V�CW@<�UR�g�<�X��Z�sˆmAed�RA&h�Χ�  0 �`]	~8(uǍ���L���Ɏf%�i�d@���D��1IS9m���XV�7��ԡ����U��l��`�Q�B�]��yb��i$�b��Y��eHC��4��R*!�(���7v	 �C���O��̻B/��b$�Bn� %唐:����ȓ{C(Y�nk!��Ė0���-N�#� a�%�V�\H���I����b�ґw]6�?/�<Dv��E@�:6���0$"�r���2��}�6��#��%�7%��uШ�\&V�A��ТY
� 蒁Y=>`Da�Q��Uz���눝IQ�$g0��2U��h 1O��*o�>k'�����`"��ٮP���&�������`��ᒤq�-�;+��|3"O5����'$-2�,C�CGj�2XI��(�B�!�*�� .�u�%�%�.�	1v���ˮ6�&�R��J#c������Dg�!��7~j��1jN>[�����B�/}�U��V/�����m��j �͊�Q7|f�ұJ/�	�z���	�B�a֪T{R���r���C0iP�!���T�J�E�5�(�gcD�J8���q��\2TH��#�y1J���#(|O8�3��R�F�RH	T��r�`yF��ӕp�|AƤB�f�4����E*qGN�eG<�i�v9����a�)0�P�����)(K!��W�O$�����E+�D��YEr�����8F�B��E%ʎ��p$�M'ʒ��ّ 4�6�taO+t�~�����.�.$rq"O���Ȅ)�@%Q�BF!$� 	℅�.{�L�2lՐP"| *b���KR�ɊW�*�Rc��n�[@d����Ny^�rc,z����D��>+T�	+��HO��b��ƪ$,��+��Z�:;�0r��gt�b�:Q}�ŉ��,�z�' �D&��j
�<1r�:y���yb��8|��9���&j@�`N�'� m�Ç�q�t-��Z�ڸyӢմ<~����D��	kX��{��B8���ye��c'�H�W�<U&��	�R��ih�ͦ~ n�[��Z�Ӥ}&d杔f�>I0NX�t��;u�d|B�ILÌ�ѩ]�qHp�&<^�4������Z$Vl"�K�MKʐ��i�o��M�@�͒)�x	��#VS��a�^@��$r��"�z��`�3C�q��k_,l�ЫC�\�]��1�`���=�˽;ua|")xU���$9u,� ��Ÿ'�|Q��#J/�ܓ"�#F�1�3	��)�'N ����H62��
�G��H��yZ��7GһV��0�싢c��Ԃ�%��}v(�[�P Ͳ<v�-xX��?��w�ޥ �"�"�V)��`��3Y5{�'�hda4��HI&e��-�2�j��G�Ms���fT����C(�bD!?ғR��tAT$\|�j$��S�)��	#`G.�ڠ��Ef��(�OL(+E�U
<�<<Rき�0}�ф�rx��������-H�JE8���&<ʓ1k���.��	�=h�*�8�E�?))�/@$=���E��-H2�&D�d(����f��G�.r�ͨeOd�VP�ԣ|�� �ξ��D��4e�-s"� V� �8���V�Z̆�G;�)�뎣�v��*\�Y7�Dz,O���/�q�b�P�?#<��m���ACS܁�$�X�<�w`����ܓ��9ܦ%[�/�U�<3�Bj� k����8+WeQQ�<IP�(@?Z�<$�~��ы�d�<����;bժ ��߿.P�LC2�]�<����UVx�d���~��]Ç!b�<��)D�-,4�(�AHQ���Z�Ba�<����2��t����,�(_8�B�T26Yc�hƢZ��WڴW=C�	g��\�rMZ�1�a�ب۠��8eLN�S�S���`��2	�T���4vC䉔e��p��I�x��@��ߢ=�6C��8I)��0�޺{^�`�1��&E8C�	�p	��yb��u��qɵ+N�^v�C�8O(,Q@'�2C㜭����Zn�C�51���[����/�( `4�R�>C�4o<ִJ�	�A;ؘ[��?t_C�	T�j��`��'Lv��З�9�C�	�P��vj�)�`��m\�S:C�ɦ~<�������w�v��u��/�B��|�b�ʒ1�
ѹłJ�Q�dB��E"0��(���WN=��B��U������#w�H*֊��B�����"׻�z�(��ѷC�b�� ���7�ا�π �D�Rr��R�l'k���"O�q:�eD��4��M�j}��"O�(��	im�DZs(��*�vH�`"O(U�p&61����� ׶��"Ov����̊>�ТIR�*��"O>Ԙ�#�
o��[���;��y"""O$,&���J-�-��iI.��J "O �A�m_�� "H ��Ld(q"Oh�q���:�QT�ˎ\��k�"O���PD�9����
<����6"O�0�7 \�LO��#�P&�䜸�"O�00�Z��p(�(pf*@h!"OR��
��b�e�w��V�4	�"OЇ!*���qօ;]���2"O|a��h�D��	#䃤p[���"OV%�P�C�H����)�/�A��"O�I�D8]���aƩF�48�rG"O����9p��p�ӥ��q�u"O0����-4�� ��'{$�6"O�{u�U�f"�
�刍^�T�2�"O�]�4�^�s�MG"�9 ��`1"O�\X"/�8�D#�(ߢh�z��T"O,\נ��vA���~��PA"OHE��R�"r�ui&�~D�is"O�����4zr�L¡D��	^�+V"OF���eܭ�v�yE��'�P�D"O��d(�t��bI�~�b��0"O�	��RM=�EJW'^��Y�U"O�R�BV�}�dU{�	��zP"O=#1AP�'��t8�*Q�4��Q"O�$��/]�F�2�� ��6�b��"O�ic�E:�zm1Ei�4uw�p��"Om��
B,`�܁`n�ȃv"Ovh����D�TA��鏩&� ��"Ozy�&�VG�D�V�_�;B��"O��
���-�P���h�Inr�Q"O&=R�]7q�ȰH�E] 9c�"O�Ul�z�L�ň@�~G��H�"OJA��L�(u�ɒw$��m֞�"O�x�+ԎiW0T���
�|���y�BDyOR�[������'-�5�y��_AM�XY�f��o��HG����yb�D��@U���āa
R�c���y�D�+V����e^��yg��y҄TBr���Ĉ^�vq#�\�y��
\&20 @aBV1�)K�y'1\������L�v�l<�bA��yh[ �%D�ø224���9�yR�)gV9�3J?�*���n��y"͇X0Š�P�/g��[�O���y"�210��[� �
��v!J��yR �:)&�4�4�Auh]C�iB��yBҒ�q��F���`��C��yB�U3v��(q��7!���U!���yr�\�D�*����76��ce���y�.��i��k��_8%6��5��4�yCI ~	j� A�4a4��Ԉ@�y�À�cR�Y��]�	V��6&��y�J��3P��G�_��q�آ�yR�� ���Ô,Z@ؿT�Z2�'�x��ť�L0���·�~�С�'H��� d¢WR
��'� h�)a	�'۸��� �ji� n
�@��'P�TY��O����\!S:e 	��� ft9U�G7x�t��S���k����5"O��+�l�aN�s��р*N��E"OQ�a	֞c�D-�d ڜZ�^�a�"OPHa0	 ���FI�E���7"O��H�+�L��l�mۃ#�xu�w"O�X@нn*��@,�/!��}`"O����j�"д]�2KW�_�2���"O��)�&.��(�*]�2	�D"O�ݩ ��4Ò�#�ۀ%`�r!"O�l�f"B9>�B��-i?�ej"O��[�W$E;jɲ�ƻ��D"O.|q���en�������U��"O0d��AX�@d  �m��Oa>)�s"O8� �H��Y�)h3&�8M@"O�qB�P;bjR�[H ,=2��"O��J�É�Lgn��� ae�(�d�~�<�2�P"ƾz���:zr��"��x�<!w	��l��e��'�*��@�z�<�G$Ҹ (�x�GB�M0����w�<q�' ��h� �-^��Z�Z ��q�<1T!�f�Z��ćB~��".w�<)��C��pC	���	æ��d�<�Da�15��u�YIy$��ҩ��h�!�$^2ga���SaٿIXL=�a✨�!���8�ЕcŧE"I��	Q�'F�!�d��I�A"�ύ�$%*Nљi�!�$´=@](�\�5��I*�ㆋC�!��C�21��	�g��sTBN��!�$ǘ=Œ�K��Z�:���7��\s!��L��Ļ�kӑ [�ɇHȫS�!򤖷N�� �j�@O��	U�Ơcy!�DdvQI��+]8�����+1!�č�^0Z��4�~>8,��%�!��N�4y�(��OM�5���/ӵ>�!�$	1
�I9��l�L"���U4!���8K̲7�R2����g�!�ɵp��Z��̖!�x���띱w�!����g�c{�)ɓ+G�!��[�'hRk�E�PY���ͽ �!�G�`L ^	]gB	G�T�;�!�D�gp�i��O�WUڝ��"�13�!�DN�ɠ�c�kP�2� Sub��!�$�]^6����6&!�Ђv�Ϣ#�!�4P�e�� ^P�	ĈC�C�!�DN�b��!ǉ�W*�a�#@M�@�!�d���4��F�#*fn9�1aI��!�$��w��D� �U�
`�I�!�D�+���%iG�"SL�S�jB3_�!򤜚OI&l�׮ڝnJ����� �!�16�� {C�D�7�1Yp�*w"O��䇤~���@���$/�`a��"O�R�� �pb��T vu��2"O�� �ʌ <Œ<A㦍a�h��"O. �q*�^����UF�U��X�""O��C�w9�(�����%{Q"Ope� ���!Ҳ�����o^�X� "OmY�Kٕ2�l$��k��6"OL!:�\���Ac�+5Y�b�`E"O4��)�@c�)R ��,�\��%"O�U+�7~�Ԥ���"�����"O��j�h�w�����HɃz�f!zF"OPAC6�J%��2�����Z�"O��ag�����@b�����"O�Iٶ�%'�z	����M*;"O� �lK��C���x8hX=|�X#"O���S��,��$J�*�S��ȳ�"O�I��˹J��j�)b\���"Od|*��,���*�iѷi3��e"O�� ҮժMF`��!�*�p�"O���$̘��waͪA�uq�"O�CE
Ԛ?��ۇ@O9lh�r�"Ob\��-�h�隅.V="E�;%"O�{m� #�����?!��v"Ob!�3%)93��y�l;oBp���"O��ŮǊL��(��� `�\Kb"O��FN/���������"O8��g
�`��Z�G�L�"O����?@��q�@g� ��ezc"OK� �p)�&Ω5q�R��D��ybS���2'��LHg#@8�y�̋r8)3%K"D�I¶�ܾ�y"�]�	�Jۣ'���"�=i�!�$@6�� أ�޿cz� �!u�!�P�c&�е �9L@��ޯ�!�޺@�X]�H�)He�w���1I!��'C����f�<j6x)��2!�dMw�������Z����m�!�ۺ$ ��7*�f�a�ʳ&c!��@�̰����@�Ȁ���aвh!�dҌZ��i��m�#��xٕ���!�dωvp��!�1v֝b��0�!�֡oK�8@�-N�x}[����!򄖄cy��
���i1�ݩ���[B!��^�>�z��ӯ�9:vh%L:�!�Ni��r��˲��݈C���O�!�O� )x�2�U2jT��i��b�!�DI�o�����S�b(�l�1�}�!�D�B�Tp�.H	�`�0-�!���4.�><
�Ln�u3��0Xq!�D�=�� (��P�.�6X*Ivf!�$� ��0���ͰN����pc�'u�!�d���Hj��@<&e�F!��Ey!��\�mU�Q�eۘ!6ڹБ@E�uX!�^^D��"4d�ĸ3 ��7!�䅝,Ӷ��%��1>��H���"!�ă/	U�,��N�8jdAb˂'!�G�-I.A������0�E��`�!���""�^��HT�Z�2`@��8Q�!���-�qi�C�9�i��Ҋ)!�Db-��a���O���O� U���d��p�䁰ҡ�Mn�"�X��y�n,���ZA쁗=��L����yb� �y�S�լ&-ډt����yÜ$	l��)B.-���i�#�y2k�50���.�6����B8�y���xRp�PtĔO%i�se���y�*EUd&PqƯ������9�y�J�:"V5��>D� �d!۹�yR�6��E��,�A�u��▟�y2��)v)��,]�.�,�Y����y�"A;<�D�˂}���O�;�y�o��j�N�`pJ��UL�ҳ��y�bS�����4HG�|�����yB�g�-�E�taV��q-�yB+��E�d��לw��"�ڍ�y�F���3���l�L%I5(���yb�Ź1Z����	g=p$;���5�y"��S���i�@�aX���y
� -���D��l��h�(� "O�x�������5dه<� ��"O��X��4�Mc`�HG`���"O
dЁ�*��g�@�#
M��"Oܜ��$Ն/XE�/�P)J`�"O��п�Ƶ9b$qT��"O�,�`M� UH}Em9*�h�7"O
DN\���L�p��o�n�f"O@Ԋ�	M=q�a�ce��+���k�"Oܡ�����U����$�6nƺ�AB"O�x�$�	f��:�D��g��"O�̘���fЊ�	A�oXR$"O((��KK!<��Ix2a̵s|��)""O\8:�� OXze�g�P�3��#�"OV��B�4G-*@��q5H H"O���8|1�5�.
Nu�"O�E��LνL����L
�$1�"O�uˆ��)�j����ؽ^�bL3�"Oh�䣈bI��&��2�Lx�!"O�EZ���&o��	3c㌋&|1+u"O�=xrm�&Q� ={�!��\@"Of�1Ud�+*@�*�@ޡ	Ҫ�P�"Od���':,F����MI�.�3r"O��w��*v�%���#El,� "O�my���B�R�f���"O�@A5�ڜVk!h*�-�Л�"O�\��'|%�=�#	Y���Cf"Oh��
 3$"��E�C�g�̭�"O����L�m����!c��
�"O�8���������K�.�)W"O�8�jS�`9�@Ia���.�>9�*O|	�T�PU�.��WH $aQ��#�'�����*ƪ3!��ad+��aN����'����'H�7H����郖g��09�'f	�ܬ~Ɔd($_�^��T�
�'��|s���fӦ�!��#@��
�'��<[��N�O#����F	o�z��	�'���ZҐ��%��B%c7�LE�<A���c�|�š�Cl���G^�<�"��#`-"`
��� �*�"c�S�<	� /�j�P���\B��Öm�I�<��6K����rjĳ2�xi���
^�<� �(��y�dje)��+!� 4#�h�I�OHMG�$�A�Ԓ8 !�:)���$iʘhI��QAS�o!�Dȍw�l�;S��%_����]�!��/0N4A�P�ܲp<��`V�2�!򄞞-C��9B$̙@�OU�0�!�N*e]��C��>)B�/�2B[!�-fpf�# �>s$���M+B!�D^�
����Ӯd��f��5�!�K"�Di`��º.0�d�Ba�$6�!�d�4K|�IK�/�>e�q�`_�!���Jq;R�_��;w��a�!�D�*c�N𪖊�87t��"��!�$�b�JX����`~�A�s��o��DE�&2lqgއ:�=�V��;e�����Q�Q�0 �nN�f��2�5�OH�8 kN� }��Hƿ �\=� ��x�W
�4Jf���#��.y��hI��'����]9 $��y��|c��[R�11�O�+��ۘ�bؚ
ç}�zDb%�4�� �%�R�+��ӟ'�%I3�O ^�(1b�"�x�O�����]��ܳGm]?�M��l̋:������?��/��;�ĸh	çLU��!�ۦ "���G�Nf+�Y�DU� a$�Jw����E�L�ʧ7J\Yq��^�ide�AA��V!�=��a�����'8tB0:�-�W=�qC���@���Ox|�"�)�3� N���U*��AH�m%ڝ��OB�J@�>�)ڧ6����Η(�l�)s��<�x�jc�JP��O�?u��I��;�2�� HϵX�U`�o���'-��;Ψ�l��m���D%�Ǖ�Y�+7��0޴b�h�jq\Mp���?�'��OR|���"y��I���)�`��O͋�>�I� '�|>=�"�w�0s� 4۠�N ��6�w�8c�[�4ڢ-O�?ux�j�	LC��bu�Ŀj�9��G����$��V剓��g~��l�j�V�),<YɐCޕk��q£��*V�j�'����g3��u�)�;J-����T��ڱЯC�0O6��CO _���	��3� 왒MO(7dU��D�?m�Ql̢4�'N]#�\�VV)�l>~r�'I2,����(a$Xpƣ�<L9�:�'��5�6,ԓP�J��������+�'�4A��l�2�8��N�6^�H��'�Bᦔ}��Q�%�C�* ��'��yÅ�Bi�ä�R�$�R�*�'`�ۂ��.	�T���O��V�{�'0j���]�R�Ĕ a԰|����'�$�d ���s �ߨD����'�vp�쎙T�\��Fn�r����'�����"[[|qv+J2e����	�'���ypdR�k?�qq�N�?X$��'jP��"�^�^�>�����SX�]��'�za��bC�p�\�Ѷ�ݰK�z]2�'�%��#��q0$u��JW�{	�'��ȹ��@��	G�(��u	�'��ȣ��)\86�1�lܭa6�;�'"\ ;r�>U�^L*skMIP=��'}�衧M�0JvT��rO*q�,(��'&��s�����S��Y0o��$i	�'u'[W�jQJ7�ij|�k	�'�����V�
��N�9𶉑�'��EQpȌ9ND<( ѩ���4u�	�'�И��`�)O�,u�)߻Z��3�'�x0BPkZ�d�(�@��~>"�8
�' ��d� �U㦭߆j!�t��'qBP��MR�I��8�g �\3���'��\T �Qlx�G�cێa*
�'#�*U�
D�Q�߈����'"aq�%�77jՠs� �>r4u�'��a��Qt��;C�ý<��A	�'�X��e��RL���iwz�'��L�'�
 '.@�a�ȓU�z,�5��c��R@X�̜��h�tyZ��
"Z�颣%��yk���ȓ#�x$R�-,pň��Ԅǋ9H���M�ECdb��	����V�p��م�E�^dc�)R�n����	�+�q�ȓs�<�j�㏍X ��p�)C)n}��r�, Ү;8l��[TF��*�
���p.j'ʝ�`����q)kפ6D��s��e���P6H�IdH!bR8D��JF�O�2���捔wc~a �M6D�d)3�ǜy���E�U�Kj$@DB4D� X�(�, "�h�/Q�R���cA�,D���7F��5ق����D/�q��.-D�$p3 ��'7&��Ve�k�����B7D�8H��Ԫ4qg<\P���5D�HQ�-�J^�0��ka�@P&C8D��*��\n{���f���j�,p�R-6D�t����p�$5⏇m��Kd1D��
>��P�S�B,�ص3fe<D�pz�C��;���S(�%�򐘠E<D��(�G��p����̀&,Ԕҧ &D�� n$���(:��jR/�)[�-۔"O�q3$)��02(Y%O�k߆��"O�e�O��}�,!@�Ҍ���9R"O(�@$�  dtYs�C38���	�'{"@x K�7|q�y"#F�[�� �'uZ�[Q��4�^P �J�VĪ�'0�t)3dĹJ�Νd��Qu����'��4����"AZ�hc�ǕQ�8}I�'n�Qf.O�ܕnዒQd���'<��;S5��T�UkrC�}��'~I�#nH���YVʃ>lt��'�X�ѢfSS�`�#S.M2�49�'?�$�V�'#Ϟ��t���J=*���'@��cӦN �(b�� �1�
���'jXCg��'f㔌[��80�*XR
�'��tBN�X�q�P<t�©�	�'Z�uB�n�H>݊t/�kV���'��hQBKW�F=8Q*�g�2���'���f���BS�&Lv���'-L�CvhU�	��C�P6<T �' py��.H3u�Fa�R	ҏQ�``
�'�l����U���@��I-sEXMR
�'�
�"(�#бsGǐ��8Q
�'&HY���o�
QI���/y��
�'!�ȓ6͌�z�j�P2(M���	�'z�;���fꚠȂf� KEy��'r���D�B�mgHm��iQ24w@`�'�a��ƌ
p|��N���9�'��$դ�7
��!�B��uz\}��'��O��LQ��
s�Ad�DH�'7�(��,ԋA���"*ׁ]A�Z�'NJ����q�L��^/]>���'�8YK�ŀ?��9*w&Z)Gx��j�'�r�p�D:`ְ�"YU`��
�'fx���"ĄU�`C�
�5vP�#�'Q�-c��zY �q��[4����'���p��ї\��EdY�+�"��'��#GfA;]������-�����'�#�K��QH8��膾$ޢ9��'��ts&�� |�r�`Q�	��Q��'?����周vh���� �z2&��'JNh��(	�����e�ȕ
�ڸ�
�'ZxP�M<EbP���[�v�Va��'�VZJ��q��x9Ӂ�8o Q��'��`Y���:��԰�.V.y$I��'�zH�5b�G��C�@�Fzn�h�'�
�ʠ��!�x-����"@��i�
�'�����ȥk��쳡�ּ)�B� ��(O���Im�h�eLs�����g�<Y�L56 � ��4	V)�G�I�<�ƙ���Ua".��p��pr��M�<I�f�YTB\ ��`���9�Tc�<�3�٩">�8ģ�LFp��ok�<9�	:8U���Ae��1�u;@�Tj�<�A����S酒sd����i�<14O�u�����"�U��փ�d�<�V���S|!�I�  ����b�<YG
Q^���:���Z).؅ȓ!�=���Ǌ����_>���ȓ�2l���c�DY�� 082�������K�wlP+�^  m�q������!'�����E,>, ��,n�y� �ct�Yc���$�ȓ6�|š�`B&a6���ǉ|jp���S�? |�@�쒕+\��ч#L��"O��!�O×I�0�+t�9U��x%"O���POܖ9��5�bk�H)�[1"OB�x�G�-#q\Y�t`Bm��X:�"Op��"��@���S�`G�-��H�"O)P#��	���d/W���@�5"O�3u�ߍ[�t�c����0lu�e"O��ڢG�If�"'�+|0�9�W"O�x�U��q�$�I��>�"Y[�"O��R��F1�i�C�$䃐"O,!�(~�UC��T�f�Ւ�"Oh8�pƒ�Yh��Aлpm�H#�"O.hXu錊Ii0��W�]jn��a"OX�8�oͩe,�QB?	M��"OL403#Ș4)��
4⋈9ޜ�+�"O� e���a�(&
�<�é�A�<	��Ȍs���r�G�l|��ZRjR�<��`�R��g�/u����c��y�T�u�`�4��1SQ0�|W�C�/ek�QХΟ+|�t�㨒�F9�C�	Iۤ8
B�?*f@�2&�4SC�C��$bSx] dB� ��E�C���u��N�
�����p��C�	�;Ɖy@dɻt�(�V#�8p��C䉏CJB1�f+�%�eq'�Y<KjC�	�Cdl|�����x�y���3,�HC�I,1�:�  #L.s�x��r�sidB�I�_����T͆�`~С�_9dB�ɤCՠ���倷ղrr�B�Ih�x�@���uߦ�)���5;�LB�I.)6}�aJ����S� B�	�,�3*�0��%I�*P��
B�	(y��3��a����H�M��C�I�4��a0#�̄mI�b��+�C�4R���bZw��q�1��]��B�I�pb�tOX��B䉎v2b|�5)�;H��ːY&S~B�I5-�x�eB����pf�2k5ZB�I�b�H��@K�+X�b�Zt�]�C�	�-M�K���OO� �W�ҏ�&B�ɂ �Hd��˶o��U �9=�C�əJ�>! �F�1Ď@9��	�v��B䉏7Yۉ1O�-0*�L�f�F+�VB�	: UV9�Q�F��r�A��:	B�	�s�>}k����\�fDR�U
�C��7TRy���Eo�,�[Ag�1ѲC�/, �É�-���SF�)/�<B�I�k����a!EО9
1�'�B䉺_"���t@��tl`�9ԯJ%	�8C�	��|� �C��<u��)�6G�6C�ɓE�6]aA��UF���5�pB�	4o� A�fc��k���a���3" �C�ɚn�A	 � ���E6j8C�ɎL�x���@�`d��-??C�	�@��!M�8F3b5��V,)�*B䉘o�ʩBV�� �:�biV�Q�B�ɑ"�v�)޴P��zpLU ��B�I�E����V`�+Rx�=�WAȼ9V�B�I%/�4sw�ОVߒ���v�dB�	/n�tYC)��V���åV��B�	s.���ٝ�]�&�k�B�I/bNbi�&�CK��Lj�K�l
�B�	+u�RW�M�����C!��i�B��3�$�I�l�hi�i ���pr�C�)� Ņ 	5�ԁ���0$���Q"O|��凴֘]� %=�����"OZ�Ke��z�p�q��-�±k&"O`$�wgT04x���`΁.��*�"O���FCĸS�dMh$��e��aS"OT��fL�7P�	�����F �z"O(�Ae�; ����,]�Q�"O� S�ʑ�S�"��!��e��J�"OTjB �4����(�A"O��j�fJ+�	����ታ"O�x�M��M��QiDŹ@�� ��"Op��p#�'\y
B�PzhF���"O�`���C#`b���S%8N�0""Odf�Z6$Ṱ�qNZ�5N�Uz�"O $J���EŐx�fn��L$��s�"O�@s��[�n7�=!0���&Epw"O�$�&w$"���/D(b��	"O�A����}��uK�-̬P
��%"OqJ`́�A\t��@�Vͪ�"O8����sʊ�am�#e �hi5"O(HsMX�7���ƍ.%��A�"On���   �<�>���M��#�0
�' ę4e���s��J�
�'ւ����Ѥ&�r�ql[�wZ,��'��x;�O�OF��AƝ���X��'� �I2g�L�!.]�x����'�hLXp�ŷ@��``�Ĉn1<0�'�J=�ԫ�fi)�� ֧5,�	�'�P�ʃ"̌.RC@��3	  !�'}Z𙰏R>��!u �>}BH�+�'�@pA�*֫B��9eC}�ܵ�	�'��dm��PJ�P�D���T�	�'7��J��ބqϮݨr���v���'8� �'�	�#�Һ�<Y��'Y�Tp�H��B���e��Z�ș�'`��9�b��3��ɄL��VD4�'^�z �"dI6���A�~����'�L���E�0T@J��Q�	�Ű�'r`���"�)Q�dT�iN�}tU��'��#��אU��"q�Ȋ����'�,�&��x6�Q3�E�x�B81
�'�.E)�/m�hm�"�\�<��
�'/��[�c�>Gj��Q��Y�J�8�'� W��8_�X:f�)K�H��
�'��=9���6����AÑ41׮��'R�IgC�*>,F8q��^+�	�'w��"/d�d؇�zx�ȓ_?�d3�$�.<�v̂#�Z<{���ȓe�����X�
��J.g�E��s<x�K��X�)������!2����s[��!O?t���b���b���?c�M�V#�
fn�@�TiS�	�z�ȓU}n�X"	� `�t�ip���I�zd�ȓ��0��/o��@�W�~���ȓqx�hH4��@[�"o��T��:��91B��SLx����`k�e��1� &-
R�	���a����ȓJ-�i��].%b�D��$c�X��>FlKr� ��T�7���R�x�A�ҧP�Ш8b
�	���ȓ$�+�L�F�8(ȕ�]�0��qW���CN�����3f �:�u�<��G:=Ӝ�!�JS�8�����_M�<I�eP[, �0���
�f��FLJ�<y��ӥW�^�!IJ�/�����DCG�<W͛2u��q��-D����iX�<IPF�����`D)�N|��{�<�6�K�x(Deˀzmz�q��}�<!��Ԧ(���C�/>,��-E��hO?�	�o�8�%"ǜ7h0-k4JN:C�)� ��y�@�552���j�s�"O.�v���P�[��1]{J���"O�SUJƃ/Ծ���]�.c(�`c"O	��	X�)��@E��a-��)p"O���(ƣcK���%��K�"O���Ҡ�i�p�z�L�B��"O�
�ǚ�x`<��ڨE�J8YQ"O�r���w�x����:��u�V"O�AEلb�V(B�ٻU��E٤"O�|��m����t�����C"OV�ah�3U��E�qA3.��y��"O Dq7$!������*۰�"O�y�Fk6�ܴ toؔmΠ0��"O�=����Q��P��Ti�0a��"O�L��Ϙ.8���c�:�!p"O*��K�,PG�,Q��D'Q�UbG"O�<S�E#%��ز���-����"O�ճ"�6�Q���@$���"O���Jޣ^�(�(Q�+\t*�"O�t��n�E�(P1h��C\�p"O\��dG-R��EÆ�U3�=ȴ"O�-@��+i� e�<4ed"O� f��0mZ�Ia�$:�JT"O��3��đ|��a��5ކ�!�"O��JB�oda�4��l� � "O�kP��P 4�S�<6����"O� š��^�j��S�D
"��y"Or�Ca'M��� #�ўX�d<�"O���d�_�t0,R�S{�2Րg"O��'.�\V�����޺��'"O�����LK��1����0}@-Æ"O@�x���4j�^+&)Sc��"O���&M۵2J2ѱ�"ֽVF���T"OZ����&R5Yc����09^�c5"Ob)s�I�b���e��aז�A�"O8��C�ܫ)���@�H�'�L�k�"O�̰��3h��Ԝ);`"O�09w���6�6Q�&^9oӦ<�"O�)1��`"[��Á�
T�d"OXM��m\�o��5�P��D���c�"O�5�wJ�~��u��@6&�̙20"O���`A�y�@؃�K5	����"O$�سj���ѵJA=7����"OTi�MP)Vp(#�C#x'p<��"O��H�"[�[�����ė$/*&A�&"Op�r%K	s�%(�c�d�TMK�"O��S���^�B� �+6�A*t"Or\�Vj	+Cع���M�[̈�Z'"ObmIħ�K��};��IN���E"O^�څ�ͭ;����!Hہx�,���"O��rp��=�LC�L	���Y�T"Oΰ��(��P�T��=w��[�"Od��+̋�z�ea�j��A<����هz��:�F�>�h;��ט�!�$�&p�rQ�ʩ���D+�!�dS�y
< �W>P���jϋ!!��%�t80Ȑ�ռ$9��+ !��P�i� [�����F�5!�I�rt�w�S_��ڴ���7�!��7K�|S�Un��	ċ	$�!򄗼A@T9JGrά��
Y�)�!�D�������N"l9B�g�!�$����(p��*�8�g-�3D!��C�Lˣl��lX����4!�� ��k�F3	TJ��Ǐ�}P�]��"O����d�j.b��p��?^�#�"O��bËߣh1�lx�g	�����"Oz)�k�(G�հ���"|mc�'t���H]�x���C ��|���q�'��9"U/T#.|�z��M(K����'r����؛`�����`�B�Of�<�/��FĞ�7A"	e �Pkg�<!�X�%�E���\ڇ�A�'�B�I<NtAi��C�CE�����[4PC�I�x��G	W�Ƥ�@�R��FC�	U�
�I]�P�bN��m��C�I�l�t�jD��"A�6 ��V�fC�I1)�zٺ�Ǐ:yF��w�Z�T�|C��=V��uyW��,�6���� �JC�	�F�< Cȩ-,����9��B�(p���qE�*Op���Y�1��B䉼0������4^s�"��ԨB�I�.�(�D�A}]�}��%W#`�`C�I8e�<B�ʟ�:��-cQ�J�O�8C��2+�ͩ3�A�aj^�	�ĊDq,C�	�C�.�w��AJ��.ԹJZ`B�I�aX�� ��H�AK�I)+�VB䉴iR�    ���O�@�;�?�������#)��@���n��ؠ	C*jF�8�$[�3�nX�E���:�0t�↓Q)lMDy�&۟��,��B�-����x����V.I�.:$�2ʓ��*|�$�i��X��)��"�� �*Q�� �+�<��\ٖ!�O"t����/ ����L������W��,C��1�"��D��:�v�z�G��Si,�O�Im�B�ɚc��Q�J~ґ�� w�d��v(ü/�X��w+���H�'���'�"�&#�t���( r�$m�֮�O�uj�h�,[Kh�G��9?v�p$�'��	�E]�]c�٘ !�9�:�yקP��ř5���j��0��7ؙ��0ғD��L������'�����B_:V�l��b�Z}�(@N>��,�}p�+�u!��8��T�w�|��?i��4����Ɂ/Ԙ��4��9�z��O;���<��aU)��?�O�ҤՀy���i@oÍ>h�q��93Fr�'�`I C
's1��M�T��S=Ey�#F�&C��J'茲cCr�d��H:vHV�p�d��E������O�O��� ��4;	��ǡAwZ1+�O���'�r��<� P�Z�+]�t7�e��� b�>�ka"OL5褬�8R�|h�OF!U��|���	�Ԑ��D��*:�<q��}jqSr.Bʓ��ğ�g(�d�OL�$�O�˓9����c	�,RD�3 ��W����/����Q�'S^�2֨�6�Ϙ'�"�2Pjډ>|l�f�<n<��U*�1�~9���G�SX���	��O;�5��>�d���h�&��hXX����X�'ְ����?9����.�$ ؕ&��2h8��1��!g'(C䉸)��b��M�
�4-
i���$�O~�Fzʟ��f��TYv�ԻLT�=���zA
ۗ1k9����?���?�+O1��� �G�e0��
]�v)��B��~=��8S�^&0��,�&�ZKx��A�S��I�@�1C۰eC'�+-zh6��*4�	:�N�-_(P`6#ASy�����e�'_��;��ǯH�&q�u��������O�=a��d]�/���A��@'A��rTca��{b�D�8�\PP�?S���Ǔ]��'�����d�'2x�%?IX�ᘕ���:W�� S�h��O�˓�?a��?1f�9M�U�VĆ��͑Q�'�<��A eh�B�Lә3�D�
Óa�:��щU�^P�Ǐfb��Є!Fp�I§��j���"�ᆔx���a��Ɋ8���O�J�z*Z
��zDK�E{�'����0 ,��у
�=�t�&(�*'Z���F{�O=z��
+�$�q"�_20z��VOb_��[�S`yʟfʧ�?yw*��R�:�y�g�H1�1��?)��_+���%�&�0Ha�գU���	��):��Y�� 1xExf ��%2�I�6"���.�%�ѧ��89�[��'-���Q�'H.}��<ږJ��&��'���y���?���)d������ ��ȕE��J��"'D�$��Q;O�����N�/�eR��'��?�#��#F�����U{ƔM���,p�]�'A剛9���	�� ��ܟ��'���y!i��1�r�	'@�x&ҹ��CE�3�T9R@��O�+�� iU1�1OR}�4畟����n��o �ȸ'��l�I�3�W8��`���k=1�&�Y�$W} �Q�R���+��s��9���?��O �s�'L퉨�,��%��'�����8�@H��Y�ܡ���Hpu9�/��Pb8�	��l@���?�'�:� !�y�� �պ9l �	���7�6�R!	�pu�~j�'���	�(hJ�*�`�	B=�!�1��$�?�L+�?���?��%*�(1ҕf��x\2��A�����W��4y��@�DD �E�T��OE�'D=_T�hC�n��t݆ʧFt�Y&��=>��m�Iu��D|��4�?����O�,]r�n�tD���<0���)O���Ĉ�B��R�'U�I2D�ؕ'M�?�}bȲ<q�,�}N<�k��5?��y� uy�%ѷT<�'���x��'�"�Y�(�$PGA�l4��yԥH�
�")���ʷeƔd(R��I��θE�t��\q|x��e��8Е���y"��H3����-�gE��!�h�x�)�ӄMr����i�8?+���0�	*vr��[����O@�S�m~��78��DX�	�&�.0%��yB�X�0�c�a$k�Vm�5"����'��`9��|"P�tP�� C�'��!����?�(O����D�O2��O��d�<�'X���E�^I(A��CR�SEJ��&'[�88��\.8QdVfLW���$�	�jO�����4��E# �\]wp�����_Լ�C�'�=��)d��!_j�'P�K��Q�bX Ƒ BB��O*ɰ�'�b�	�<	@��$�Z�W�$��"�\h<� B��bZv�M�fZK	$�?a��i>)��Ky��ƾi#T*$�N�6�� �W+5���y��'R2�'Y�b>�`W	3�J���n�m�DLHA�̓w���A-�{ˊ)��M�&� �	��	�_��`*U��9,J�]��O��b%:q�s	�0\<� �� ֎_�t�!]���p)I+�HOTU�A�'&\��ӡ��&��݉6�*G2I8r�'�ў,F|B�Y7|��(�1'ͦwL\�1f���<���L���P��陓2�l]�3h�i�I�M����$^�8����~�we#Ya6P�F*X�*�y��œ��d�Ob���O���o��:4�)��ز<Ftp2�G�uw�&_q� H�l]L�L�
o����O�@cw̓�V-��n�2Li*��c"6L�r����E+�"��ƈֿ_bm�w�JR�'Q�Xc���?ш���2w�	k��I�b� �c�����1�O⼱#D2l�а�aF.(��`�|��i>]�-OBi���.���[Ƭ[v�Zh��W���6'����	Xy�_>��I؟p#�*��L=��Q��U@���Jџ8K&�"����čIń1��é{Z�>�S�O*KqX<q2IA?p��Vbh���W�sN��	�XpZ��±xq���jT�HǞ�����
DTՈ�$	��y�ى�?������4��� h�0��X������Le3�"O�
��Ǜj�PL�T�� J�|`��d�O`4Fz�O(��1��Q$|��áA�p�D�'3�I�N����	����	ٟЗ���O�7}�����_X��l�&�*�,��%m�X_���6�Ǯv
b��ʟbL�>��F�V�L��ad`! -����uB,d��a*���O m�rmP��&�l��O�yq��ЪD����.Q.S���`���˥g�O��D&��y��ɩIV��r�E�!nuPuJ� ��x���9mQ |Ic�2$ @ ��ދc���?��|�����.c��¿}A�7&L%'�!�ॏߟ�	����Ify����I���ʄ�a�Fłu�O�>���g�U^fa d�Y7H�z���(q�'��|����dv4e`��]�#�`iC�ZS��[Aח,5z +��@�n����6ғ��!�ɳ$`���(��	��Wqߌ��	s�'�Q���Aֻjꈲv�T_�d{��'b��J���sBa1�� V�ܒ'�<�s�i�V���U)E�Mk���?��O�|�)T��s��pl�6nA��\��=`��?A�آ�*�A�N�����>���/{�ɺ���b�2��������%�zX �³J��Ep��B�O����,&lܑ
�S 	rv���+ޗ6�6ّ�) j���h�	�O^L���G�G��`+�çFl8�(���S�<1$�3��h(�G��F� �lQex���/O�a���8�:"2T�X���Iԟ������	y�4�?� �Ʌ&FU�I��	� @2H+��/O6�=yT,�/����`U�|'�	���Z��vx�%���~*�
�L�-�9h0�S�j]~����[��"}*��$�97C�Hs@�}��h�o�m+��U�"?�ї>���N�$�S⓺���jb�ޔ5���caI�}��C�>9��O��}Γy��c���	�퀥��	Z*D��'F��y�ĝ7Q�.* �I;>q��04����� k��I�$x&�'G�4���)�
��C�"S�h�����V]��L�Q��e@�_�LɤOd�o�
D�Q�h����R��%X\�O�5E���oTv�PJޏZ�����(4���9U�ӧ�9Ol8`��|#�ĺ9�}��06���s�YD��`a\��'���D�$��V��a�Q�JLĨ[��?!A	����F""?��y�h7�~B�)��J�3{X KN��?�n3�	Ɵ��I؟��|���R�O��$zP̒;H�rt���_R�<yuK�T�ި�Q��F��6�	Ǧ1��Zy��'V8ꧾ��|nZ���� Gc�'��q��77@��?�/O(�=�O;^��W��,�1���>8����'��v��e0�)�,�\a��$#O�}�@*f�tT���[����$"O�ͣ7ϓB�<�5.��5���id"Ox��a�[�V.���,O+5���T"OnĚ%Ԫ�Ѥ���P�Z]�&"O���EĬ�G��8g
�Țw"O�D�GBAj�Y8�i�*�;�"O��	%)M'
8�!�蛴f�ܒ%"O^�
�l�*�h\�b��*l��"O4���C������"a.�J�������柜��՟����
[�L�b-�6tbU�!�M{��?)���?i���?���?���?qb�ނb�X��F��&�I�	_*��'V�'��'�r�'<B�'�KZD�\�t�י�Jix�P7�J6��O����O:�d�O ���O����O~���� �X�s��fg��F� ]lş��Iǟd�I՟L��ڟ��	ǟP�	�u:��H�?Lk�<RE �/�H� ش�?����?���?��?���?���d� �3He��+��W aU2�▾iV��'2�'���'d��'�b�'"!�3��W>)�!�DJ�`cf�|Ӻ���O���O��d�O��$�O����OnQ	��m�ԅ��+�#����E�ͦ�I����H�IΟ,��˟������ASi܈y��PHĻ�z]�p��<�M3���?���?���?���?����?)t N�Cǖ	��P�q�FiEOX�r���'$B�'�B�'���'���'�b�X�;�b��u@��6��ӃݕnA�6M�O���Op�D�O���O�d�O��Px�"��t��0u�N�<-@�m��l��ß���֟��	ɟ��Ix�	8l��p�J�s�H��mU�jӨ99�4����O�����j5 (Ԝ$8\9�F	I�#Q�q�`���$1�S0�MC�'28��'�K;�8�S��J-0r6�i>6�c��'�O**Q#w�i����)x�����aX�{�B�>*���9/�J%�rF��G.ў���<�r��hH<��Ň�am�$�'S�'��7m��<1O� r�Aݱ'tY;���q�Yð�d�o}�m}���nZ�<�-�L��#�L��RQL�6FJ���\� bb���.��%�(?�'W̨_wF���E�h�C���`rt4"��� @�|˓����O~�}�_����C��zt����	�M�t��c~�p�2��S&���7�_�w0�9����a�L��I��M��i[NA�xϛ曟ā�!�e߼�p��.����S�F�4�ĊP$W�Vt(��I۟d�'�1��X�bX�<hD�:�) e�b��$S��شVj �<I��$��#�Hx�Eں9~V���)��Lӛ�KuӘ��s�OW ,�揶Z�椀���p�P�0e�3"��,r�O����aE�b<��=�J�6|H�E�n]hHÍ.'z�݇ȓ�V�� nB
� �'`))����=�PJ~\���v�0� eK��f)�eeĀu5�t0b��C��|�'NB�_���\�
7�x��ϒw�����"z[(�I�d��w���IM�c��\BwQ�>_>ܑ��U7��# 7��IW��S�R����[�6����s��w�����P?��3 H2���W��F�I����"O3$���&It�M����XRt���*h�3�ԙ/����C��8sK�<r8}t�YB��(�� �Ul�kB�s�,N  ��`U@Wyr�E39��\��ԃpPx-#ELC�vd3�)ˢ75bm���9D�`Z�eC7U��1CR���p2z�c���N$��(��h��$�!Hk�"bL)i�6ть��DZ�M"t��7H���TJ%fܑއN �1�Dř]h�ؖ�K9`��F���s,n�"ٖ�lX�6�i�b�'x8�pԧ�J��h��I�=��<��'�"�|S��J�+"�I�޼1S��%�:���F$i�����O����<!�K�Cl�O3�OO�5ca-$�$���@7�ʨ`�|�P��2��,�S���ךL��r��	ʜ�#GH矨�'�0�
�|�T�'�?��D��	�6�Ễ�	� ]�$�~����'�I	A�P"<�}�G��,\i��H\�AM��� ���ADcP�M���?q��JU�x��'�d,زX��a-��W� ��B�'4t�����8��\.3@l!��U2~��Y� �#�M+��?a����X3r�x��'�b6O�5#�*j	RKW�O#�|����$ÍUF1O��$�O��F�q����dK�k �#WlA ,�����O��R�X}��?!O>��g̐/<,޴Wy�p��HA4����1O����O.��<Y7)�Τ��d\�D1:Qz����R\*לx��'%"�'��	sy�I�'�(=��>T]��J�	9J���yb�'h2�'��I�G|:D3�'��ZE��3@��ts����%R~Д'���'��'���+�0��v1\�bф��cP����t*&��?����?�,O�4�t�jⓊid�D&ƵY�8��ŮR  ���	���'���'J�A�{j�'C?H�9P�yx5p�dC*�?���?�/ORD��O���4��)�`41���:�ݐ@*^%�:u%�ؔ'�����ԟ0B�odU�cJ2�fe���'��ɭQ���ݴ���O&�	�ly�.ްXX�u�͊z��*ţD4�?�-O�<i��)�S�\F���0�շV՞eZP��>,����͡4*po�����۟ �S����?AF�Z=1\�h&�V�y�!X&�?�q�V�����d
4����a�>9u��*r�^�c�����ON��O����*�<��?���y"�A�?t��@Q�oÊ��Z&��'�ڭ�Ր|��'�"�'~�XJEػ�F=� �؎O��V�'U"�Н
��	ğD����D'�@Y����v`Q�*�,.���K���Yyr��g��'(��'��_��x�O� ��Bd�!�F��nԱt�:��'��'F�|�'G��J��b$�dh���4�ǄV1F���y2�')��'G��	kD�̧Q4�#s �+MD��̄�jǞ�������	��'���I�D�gm��<�1(N*�b�!�Ъ(T�����Isyb�'�B�'�剬Z��O�£6v��pK��A�p�Dd��MO>W���'��'���'�ȡQ��D�5O�E��
&6v�B&デt���'4rS����S�4�'7�Oo*-�t��2t"�c֏�,+4�ҝ|��'*BO�:aD�O�	��)��x���LM��I��"uFr^�$�������������I�?��'��g'ӒY N��tgC�@�X��1�'w�'�Q������.y;�I�Ђ�8<w�TA�+4�*��' B�'��tS��	ğ(X"E�%N�*.��@>���	�A o�S�O8���t�H�Rg,=4��,!׎�%X���'���'Y���[����`�	�<I�^*JV ��D�$y0J"*@H��]���!I>���?��T�)�Th�)���##L��Ld���?9g�ӂ���O,���O�O.Q�E��� ��Ƶ}Ni��<��	���?����?1-OF��n͜jTx`dkJ� �FA;B8��%���I���IOy�'��H)bR��FaU�h����.(���'?�	�P��ԟ��'R�y����:�� �$���d�q�bE��Z�0��x��ky��'
�S����e��]��yԌS(_� 3%h�ky��'���'���,E�&%�M|��KI<�Ќp��0B���f�B#�?���?),O���|R��������P48�Ǐ�Wu���-�)���'\BW�,A�Kł��'�?���� �qxS�|@(�#vH
�CִaS�'���x����,�I[�s��S���$aS�T� ��z?zx�S�V��L�'V�m�Q�oӢ˧�?Q��}�	��
M@�i��7���	t�ǸA���OT�d�O$��7�9OxʧB�д�0�i�^��J�4x���
������?q���?�����?a��
��}�L]ڣhܰl	V�`��@y��P�O>�mT8Q��jL/GI�,�rE�<��֟���k<Z4���� ?��`��y�ǢW�\�qg�[<���Fxr����'��'�|�x�KX� ����'͚�pؖ�'������O��O,�D�<� �ٚ)*�Z�V8�vk�6�?�)O����<����?!����D�P��+�.�t��H�΃�~U(�`S|�Iǟ��I�@�'��'��F�2]�� �6Z0�S�	P	kH�\�,�	� ��syR�ӣRu���7F��;�jٝje��JE�R�:���럔��E�kyrG��r̈́�.	P�a�(G�6< ���6��	�X�	Οؖ'Vxt3 �&�=������ �
$�X\��d�O�$�<i��?��
�*�?I/�0i�ƃ&{;�hZ�Ǌ"0�Z��U�OZ�d�O��'�r�ങ���'��N�9Ð�!fͻ�F�yW�y�"\���	ៈkq@O��<%?�;q��$��KЮ(cd$̚m+�l�	ryr!�7��7��|�����]��br�Y�U�*m�p ��]�"EBԧ�O����O�ݸ&��O���f�	�|r�� �*���Ǝ�2v�Q�����?����6�'{��'\�t�=�4�:pv�I�EO�)k3�-DT �;%��OH�
!�OJ�$�O�����˧�򩂤8�
�kbJ�//����K=<J���O0���O"�PD�<�OP�I�;��uq���2`���[[7��B���	�2a,�?i�	�<�Gʑ�~s�i�jKt��-Yf���0�ɉa����'��Y��r���s��)!P�l��,:"$�)Ox��*D:���ߟ��ݟ`�'����1`ӭcB�a�e	�[��E�%�6�0OR�$�O��d�<A��?Q0�D�-���E� �Bx�	�Z*j�����O�$�<y�H&੝O��U����=W��E��
�v����?)����'���'_����%OU=�.�`���$	�24�S���wo���|�	ş��i�nZ
�:���4�?)��oR��(u)�-��qO�n�$����?Q���?)O��D,#c�I$?�f��!����c���7� ��	ٟt����ԸPAÛ�M+���?Y�����!4
�\]֨�
Z�i����?�����O `��;�r�Ģ<�'
�n�z`eY�D���3J�N����?A��sh�1�iob�'���O����'�6�&jL�I��`hW��r�z��`\������*�	p�i>�O���j��ِ�p��+ɵL��L��t`x1i�iR�'TB�O�4�'g��'U֨�w̋ � ���M<��l*�'��2��'��Y��f�Sޟ�$��*$���a�#h�\���O6�M���?!��x�4�	��Zo��4�	���I&oQ"�94�J�F}�Ň��l4��	ݟX�	�%�6��$��l�S�?U�I���1��̥4�lT�V�ЇW��3P� �p�I�hl�ٴ�?���?���{ ���<���Ջo�hB7D�7j��|:`�ȟ@�a��r`6O.������?����?�4��2A�Y��L��dx�E��S�08.�S�i>��'��'j��'��$�O:�
ͺl����� Q�pB�L���'f��'N�',rV>-�����MKC�^�D((9P�H �y#B��?����?����?!����O~	=��#P��_� f�{"��[�ȿ<Y���?����?��'�f%;w�iTr�'�=
ū��,��1�ƍ'3��
�'�R�'h�S�p�	�l(�Ly2"�,YHQy\Ұ��b[#9�i�f*�)�?y��?���+m��nl����Ob�d��u��g�e(�_�/:jD+��O�$�<���?���'�?�/O���|V���&B��|���D�_.�D�O�$�!a�)n�����	�����?M�	�{�dq+�I�+P��&OF�0r��'臋#���'��.ի���?	�&Z�Mr�|A��ߋ_Ԡ�Z��O���gצ���������?-��	ퟨSv�����t�1r�,��L蟔�Ai�ȟ'���H�S柴�ѧ6X�Y�@i�&Qܔ�r����M���?���=e0a@�'�?A���?���?�ԋ�}J�`!�!/?rd,���-�?�O>q��_+��'�?���?��m�
d�8#�HA�Ps jM�?���e30�H#�i��'5��'y��'�y��<肨#���}A���cT���D�&?�d�<)���?1��?��@e�I�Cj�����)�(�����PF����'��'>��~�/O~�d�+Q���W�D� �,�X��b�+!p��O���O����Oz�d�O�uSbY�m�ρ�lРr!�(�2^b���OB�$�Od���OF��?�7@��|�@�M��4�-!r���R��E5�?����?���?����?A�"ٛ��'�i�)�0)�F����!˔�	1J��'{��'����@��m>=��ҟ���W4M��qa�/F��3�ȩ����ן��	�D8��I��M��?Y���
��� 3�ؤ�a�Rb��X,T��ٟ8�'�*f�	iy�Ofb�)��D�Fm�5�o"��A;@�'9�Id����4��i�O2���|y�ji�ܙ�
A�{�ԅ:uO���?���?�w��<AK>�}�׈M=Ϡ��`��9�}�u�ݟ9��˭�M���?���z�xR�'�� �� T��9�~��f�3+�b�Q�'��xk`���H�U�8��j�$�/Ir�L�qM��M����?���C!F��%�x��'��:O��@�e�/
]h}�7$�:4�̭[#�'[�'���� ��d�'��9�𽻲�^^�^�9�ă+^d����'X����:O��d�OF�O�$#�/B\�ʡj��R	i��
�J�<���=�?�*O(���Oj�Ī<)�i_*��	;�"�3wj�<�C�3����x��'e|��'d����A@W��t�;t��'a*@
�'�̟d�I���'�N� ���U;���:�B�0��ˀqR 1�U������p$�������c��֟�+���}�hX��U�i��P���Uy��'u"�'W�++Bu�N|��&�C�	!�.%s���?y���䓶?q����,������y����$kεI�f�����6���'�b\��C5����'�?y�'uT�=�p�ޫI
8��ň�w���{O>���?�[5~�2�ԟ����4w:W*0|��⟀�'�H5@�`n�n�'�?q�'{p��]���N��n��Y�C۝}Jn��O�����9���6��iߤ�\�sI��G�8(��h�2!��84�6m�O��d�O����V�	�x�ED�6F�fx⃪R;Q}��"­�֟t��!�矠'�"|���u��c�$�_+����'+�Hꥻi���'E"��NErO��d�O��/(��Њe '�t�Äg�g���D/���4�Ғ�z���O���;����iP%=E,�9�D�&t���$�O����M_�ן���_�ɗ>��+
  ;I*�bP�kw-�'���H5�']����	�p�'�P,I��Vc4J�
a��Jk��t�#�hO����O��O����O�!��F��ߌ�B�*j����l�CF �D�<1���?i�����dƦ�S�d�2�9�K�L�,�H%��D���?������?��k�ιb�N	�ūU����a�˛>p���,OL�d�O���?5I�C��ħQզ$�t���w�,X���Q�apH��?�O>���?1Η#�?9�Oqa`Aω��wK��e�����'Gr�'�R�'��0RA�'���'���O:T{��F?D�1 �2r��%�P�|"�'�a]��O��S:�N\�福(YK�I���7�R���O��m$�0m�ϟ���ݟP���?��	�E�>�C�ўAJ,Ԑg��3C�L�'z��GB�'��i>�O�Ll�6��?�X�"�ɉ6�N}��7����i�2�'u"�O9�4�'���'�����NkD�*�J�Y��I��',h����'��\��Z��֟��Ä�nG�	!��C$_�$�@qj/�M����?���m*�Q#���?���?���?��D@$nP@�k@oB:�>�r�.Ӕ�?�����2#8~������OJ擗c�(L@f섥C���A+Z3,O`���O�QrG�ȦA�I�T��Ꟁ��t�I�^�ƅ�$*�!�D��G"l(\�U�8��'/��'�R�'[��+E4�`��4wjT�!���mZ�8�d�B�M����?���?I!Q?��'.2J�#5p��_�wXT�����:)�X��'���'g��'.�\>���eO��M��d�:I(�P�F�� ��.Z��?���?����?�����$�O���:��Ј�)�v0��凰oٰQ{aJ�<����?���?A�&:A�)��DU9r�`�!�G/%�.�@Sa޹I����O\�O���O��8aM�K��
�,�.��~��@�P��4�4�	՟$�Idy2A��;���'�?1���Z#�?�]+O�EC�{�FZ�?y��*�;!�O��."`�LI@ R�y7�E�)A$,e����O �DA��V���O����O|�)�O���M� ��I��piH@C�e�f���O���Q�f
��1���ФE?L ����
�ȉ�n�9^7�(O�n	"�'�R�'����'�^>��F
g8|�{���'%��q@��ޟ���1��O 2�h�����oL*�d$"5!��'��'�1��R��?�'I~�Y'쏕L]�% ��C�Q	�hk�#�	�_��$?I�	ڟ��_by��M `x�ig�\�~�ҹ��ПYF`FUyBR>��)Γ"5�T)�����`�a�R�D�{-O����X>d����h�I㟔���$P�,O�KJ�tiD�#f�\��&�>d�����4�?����?���6���ay��'�Jr)��a(�Mݴob��S�=�y�'���'���'���'�z*��wӌy�R& @2�+!�WH�����C�O>���O���OF��<��(,е�'p�ܹ˄��,#
���K�9Qf����?���?I���?���j!؉���i!��'����l !L�/d$�Y#D�#���'1R�'���P�b�|>��	�D��끽n��8s�	j��0P�Z30B��	ڟ��Iß����M��?1���2Wi��S����Ti,^��I��?1������O�L�w2�����O@}�e1�N��c݃I�Dț&���Z�ʜ�%��O��d�Ore2f�1������I�?��S�PP���'TVx��V�X�F���gxy��'�>��%�'���'���K�O"��T���KKq��M�u.�'U����G8d�Ιm�퟈����L���?��������,5�Bv��+��Y�jB;r�~�I�-t����矰�I�J����O��?�ۀiL��j̛Fꉅ)i�Hy`��*�M���?��_>͚���?i���?����?��,����̂l߮�U��?����$ۮ<f8����$�O��$�6"��MH�r9�)W�׳i��d�OXxidcA¦���䟄�IӟlH����)� �,p���h �M�fN�@���+!S�`{��p�T�	̟�I㟌�	���I��J���#  Fy �)e�G�| �6M�M��?I���?a�S?��' �&��w���@
9�i�@^G8�(�'R�'��'��P>!��$p6͓8�|�Q쑉#��9�Х]���O�d�O*���O���?����|�2a.���Z9xt��T��)�?9��?Y��?I��?a�ɗ:z{���'���бD�2f/O�����2�'��'~�蟈Z3Lw>����<�Ge�?Ff)x�唪@&laJ�ͅ។�IП��I���׃х�M[��?���z7����4@�g]&{�(\�%W�?Q������O2Ua�6�>�P���ϧ9$:��
����z6bе+�A��?��%��aÅ�i���'b�O@�4�'�>�%e�MH���,�0�Y�0�I�_����	dy2�^;��Ԓ?�	Y�@�$���'��aq���H�䍴z�n��������?��ԟ ���-.!� �F G��r�nP�9ob$��#9� �?�g�J�nh�G�tX���th
`e���؞rh���$ڭC�\�x�8�l`�g��wP��´�'u��'K��Q"���\;"�3k��u���'2�'|��H�'��'���'���$	�����&�53H�!4���K����?����?a������_7]@��g�X) 7�=�t)U(�o���?���?������?�m�L�n�wg�*/x\��po_-����K�nwa��;�O�{eOO��\ф�� ��Yw�'1#�N��c��U�!O>�~,�`iț]���@�M ި���i����L9$���U�
�2 5��0j��5G&yk	������ҩ� QA�$fH�A��)�V�-z@��!켂GG	P����n�'V��[�C�.r`���&�āx���sCg�� �6E�� !��K�ktn�$�O����j���D�O��ӓ)��l8%�>	��Nne
�c���y�����B�p؞�:B��&��dץ~wt8�4�[�c��@�$�a{bLP�?����MKUDZ
:�YFB���D�8eDD�TD�P�$��U�S��0ۀi����y*�to��r�$-��]�Jh��9	4:cӨL���eC�>�+O>�2 ��v}��'y�}[�Ij�(ڲ�ұ��&��.}��w)���l�	�xi �D+N��[�*�/ � �����҄��G5Wǚe9EL@�����E��\�E�5��!�7/�̉bUÙ�21��^�bRM�?,���1J�*P����N��a��Ov��'�'��+[��<���ۜS��Ы�`�n/H���'�@k�i��:h ��OM-2�X,��z�qO�""����X m׊�(q1�瞗;\�O�D�O��e�R���Ox�dv�^i��	Ѷ�h�Hl�$�|������ҡ��Nޓ�6�A���2y�I;�>�j�K��\�%
�%g���E��}�4��W��=|�(�s�ӰZ]�4G��O��Y>]ˡ�͉ih�m���F�b�'���'h�E��OfB��
�����R5@~�*�d��X��	�'�Vy�̠-G@�c��G��́��dӣ�~��i�j��W��P���ūz����&��On����'�~�$�OH���O�P�;�?	�����C��p�˃D�� ��)>�H��iO�Aq,��B憈=��%�p��h�ۓH���''�54B��rZ��#�ΰ�p$�vW^� �D-j"��c���uױiۚ,*!�"�	J�Nu;�mA({���Ԏ�>	\r6-�nGB�'�ў�&��[sj%/�^h	!o�)��IJC�#D�󶡝�`�ua�fR>A�-j"m �Y-���'!�I
J��b�4�Mdֻ �L�e�@�M������@���'VR	/y`B�'=�	��q����>fż9��$d��P���Ƙ!G��g������
}��}a��	?HL�k$ˇ�]�vL�e���������|��O	4	*7͚):�Zi����xv���H/��R�x��dn�b}3� Ӳ"�$Y���'{�p)��/I*���<�����'_���0G�	J��e�J�(�E}���s�2����M�5:�jI�SS�C��i#�Q�!@$����O~�'N_�СQ�_5�之m�(@�ZP��$P�?9���?�ĬȾe:B�p��Q�3�8%�uk��|��Pjv�݅�u7�V(6�fY����p-�h8!��'��'I����N�`�<�����"� )1���2�+��V56�4mS�$[y��	���=Iv�c�}HO��?���?y����'H:�ɢ�C5=����r���9q>%A�B����	��	(����؄�b,!@�<�� EܓV�a(➢A��!�ǀ�0��Pڠ �47�7��O\���O���s��d�O&��hӨ�sA�ƚC��	�"��tZ6�&�T���b@��_'b�{�ʑ�w�����Ȓ,j1�.Mλ.iP�Q�M8zu� ��gӚH4 �k�  �*� ��F�@�{v)���.���R(#�i�缛��a�8Ea�e̖#8��"팛���'V�	63�"|���8h�%I��RӬ|y�$B3�t���C��h��I�R�@qH�D$7������/ k��z��4���dr�XQ�֥l�`H��H�\((��Bҟ�yQ��s�N���ɟ��IܟL�Sߟ�����#��ֆ{��p9��IdD9; �i�*a�sM�	>�.�`��D3Qs�xr ��3�̑�
�<ݖp�2����M#��Л)N��e!�^8�9ǓW��h��@$[���4�C�]kbl�6M��D�ߦM��4��':�π �X���Сy���X��@�z��i2D"O�0c�c��.�9���g�����I5���4�$Z���7��:M�2���%���t-Q~�������I<~���I��I�=u\AR��Z�R�eM�V���p"�<W����EG�T��}lR}��6���R���{��\��e�	g�~I�A�jN̐�Dk���O�u���'��7�'Z�P�B�r� ����C*_�]��Oʓ�?a��ĸ>i��+ڄ�+֨ɩG��<��E�a�<�%$�Lc�ء"J��!X���TȓX�\���䆓N�r��'���'����ɔ'l��2���$;dF�X0C�
jehp�'�B�'#�$1� 1VR��>j�ma3R>����@����r���XÈѿ'� L�>�Ʃ�>>?^L2R%�<`"=ʄ�!�S'/��t���߶:������Xc_�O�-3�'��m�R�z��"\�<���'�' uv�`�ư?�4�E�"�1��إ'������f?!��4�b��=���
o�(@�g�"/��T�ᐸ|��ӽO���'����ԩݙ2w��'p�i>�E���Rz6��#�T3g{��
��V�;߶T tCO7�~�x�I~�'�ΥXn�J�*��b��:-��y���R�p�g(O�r|��4fӑ>�5$D���$-��% �I�UΈ�XC�'D����$���n�%W-|�irG�
iC����"0��O���DMi��mI�$F�a$>�f�%^�����צ���~�'�?y�4rЈ�#�2�Rl6�Drњ3A�'�����D�-g
R�'yB�'�P֝�����9 F20��5��
m��у$�i
���@�?.ꎙɢ�� z��x�ʄ������a�����(A
{ݤ()Q�E��\��I�}��0�^w+��kѠI:G�nqc��>9�
��^P�W!�)Lp��۱l[�#�r�;1�'9�6�Kצ)��jyR�'t�'���yQe�$]e
�ҥ�	=��ْ����T"��f-�$Y�訳�%�?�Q�d �4�?9(O@U�b@�Um��*J9���@�A}n��f/J�e	q��?��$�x@I���?�O0�5iA�C8 )0�$Yb����W! ��5�u�G�y� �QL��Hzn��L�h�'���v.K�C��YvꁊW��@���M��M
P��ZleyJ�|y����~"㟸K�O�O���lӀuڷlث$xx�ȣ�ӊA
 E�矜�'<���d��)J/��BC-�$)@ĕ�yB!�7 �����T�7`9����-d�����<�F�G�f ���'�RZ>�����,D�H@��8\��# 9@T��	ɟ��	�j~Y��M�|D)��˞
=5aP֟|ם�r^��X��W 7�����-�Lc�L�&�7C��5~�Meb	^\L��o�Vk1�[�7e�P��+[-[M�i���+4~��H>y���П|�	ܟ���\�-	�L�2��&B6�`�7͊!�J�b�����M��cGo�kp�,#k�3�(��{�����1�Ɏ����X�j��{��P?'�pՌ�a���'������EW*T���'.�imm��FK6*�N�rÔ:2Uh�1�!��\
�(����=*�������D�<�ҁ�*�"�SE}�YɆ�T"s
�a��ĽR]0uQU�эZ��"gS�,*(ĻM?�3�w͐�P2=Q;ڼ����mQ�r���O��oZ�M��A��#}�'����G*V;�BmSp$U�[��h���O2���G6/wZ����D 7�=!�	B�qO`mGzR�Opҵi0�4��a�=���h��R�9�$�s�'�a��.=�:��3�%�Ѝy�瀜�y�#�����#��K��c5C�w0�u-��?1G�%^��[ m]�~:\��I�r�<U�
2�:R�Obb��A&P�<�d��^��$Xe�<c���P�<B�
��`�Dʍ?~�VIÓb@i�<i�'ȡd7��З�ҾU��0�Q�<��+D�K�T	`��>	���؆��Q�<��B� c�@`�U�L;x�XEP�<'�ɽHJ����N�,��
�g�<	��,c�"�P�n�
�ba�# ^�<)�B�xƂ5�EM[�h8dE�X�<��`T)�V��GN�'Q<�۶�Ha�<���D�;��
D�"V|c��a�<�pF!Pa ���4.H<�U��c�<	T��a�r%{cE��p`a���w�<9i'g�슷���3!H�<1uf�!�)�'�c��`�7zj\���v1�*2�|	zp��(!�,�ȓ �v��r�?o'�=�B�!z��}����Mu��c�h����b���S�? �}@%�A%8���Cg��u6�!XS"O�J���s㖕
ЎA:�tÅ"O0�a%	J�R]��mX�F"���t"O��G��_��9�"n��91"O���AԌJnhTCᏃ20��1{�"O��S�ND*"��AN���1�"O�lӇŏ,�8����Y�@��<("Ojy�#BPD�yR�_Z�0��"O6��c��a���బ��\��p	�'�P��(Ź:�aq�?w34Q�
�'G
cs�BA
����a� r�'*�W�,)��AR�n&��Hc?D����E��-���(I%���Ã`9D�0ْU�$#f(�䄆'��(�W.6D�@c�H_�br�lᑡ@:���
�/1D�����:�����L�0�` 1@;D�|�E��;!x4a� 
*/���ȳ6D�H� '!6�t��VGHWb�p�	1D�HK&�S�TQ��þlj��#�/D��9����J��R���� �~홁��R
�����ax�dC1�ɳ#��+��Bo�Xi;<O�#���'@j�P�O�8����U�����ՠmKj�z3"O�@gĈW����˄P:b�q0�xcZ�
�z����؜�Q?������	���V9J�4H�B-D��ڦ�G��zm;�kN�M3�a��D
�h�nlYp[����I�����L2ĥ�64�Z�A�/�-�0]��p�H ��3g��#4f��x���K�g��8f�Q<�p>��Ý���V�g^��sŠ�YX�|�c/â,	�*�}?�P��3R�r	�iW�(X,5�[�<Y�MR�}^�Sw�B%IV%Fz�O �p2,K�"�a�2�'L;�4[Q�L�jJ��$��	iH��ȓ0�D)�ѭ�C�h���J{��Z��ٮ�(&�q���x���Q�~�@$�M� �RЇR:��x2"��(�q6k�X��؂�	42�ـ�o�d��)��'��p�S� r����#wVi�ϓr�����"uT�&$M����v�v9Y��5N��ȓZ�2(Q�C��&+z`�.��Qj��<�#n�Ph����)Vk�K�Ӥ �����R'2�Ifx�4�g��5_�5�a�֝:ls,$�O���'���o��8�f�a���~� ���'�N)�*D3g^����$��(Q"����i�O "��oV�9=8iRS+�{�|���'��������K��R��^�@X���'Fy��)�Dtzӓ��e/�-��L#c�!�䟅	m��cCR�<\�HB�j�I�12�|��).���c�cBB@\�a.-�0?)����a�A�! SNM�U-Q�(7��1�'7D�@) �<t��� �+!�"��a4�*��~�0���i6et �#q�����Mi�<)eI� h�X0*���*FB-�����ɥ<���{�H#�";=h�p���/Y2�$*QC���y2�V!0�ԅ 6���T��i���0�f"�n]�b���'_����(O��g��u���� Y�r.>QR����9��M�s]���t	�?1׫�B���r���Љ;�+�r�FE4 X*+�|��0���3�
^���ũ���~�.��W���� �O h[�ןP�{CÖZ�4���OFXT�'eF�*s�)�B$YP�&�[�'+B	H�k�^��afʪ_g��s�&��Ѹ�E(c���妚9,H��<	C�U.1���S�� a�@B��2�x�(�U9��I*�숦	�l�kY!&.��DÕ p>�՘���02�*A�O �˱/�����dW�Pn��:ǏX�/����r���E����g���]��C�5O�a�؟r���ĕ1GjXر�*^�z�lG�mFD)f��p>�qCO�k��d��|o`�����<��.��OO�Q�Fv��Qc�?E"��ʼ2�`Y�P؟�1�"E@[H���ĕ�H[���w"OuX�J��H��31@���'��X�D��'+V�p�!
M}P��y��Ě�M�'؀ ��#��.<�x� ���;B/~����'�fh�`��LsR�:���
������Y��a�3u"����<�F	�?���e$��)uBZ�;��͛��J�?�O�ŋkɕi|�Q�,D�9�@P�U'~>�T?%�)ϸCM��J眨/��,7#n�4�	W����>ir�����)wD�MRDZ�M'�<i�щ�pB���d�$D=ܠaJ~���O���-[G�u(��A�=�����k����M�ZD�]�ԣ�.:�h����%�4�DFȤI9`��3햋HjQBAQ}�I�7X������{�VXbb@O�X� #?�"nL�O!z���bR~D�r�OQ 5�F��<�i '�+c�	s�'0�ip��*��B,۶]3��q�Ⱥo����cھ���-M$G�e[%��Dv?Y��>2��d�aA-����D0?ـ#B�Y!:��D�Xf�`i�JȢ��,k#�UsܰF�G��(�!�M355�$��~�'k�����,3ǜ�9��
|� ����h�
�6tI��j:0(�
�E�\�v
u0��7���74��diŀo����츢�0�i>�S��%o��F��<�=(RA/�rhH3�Č�^8�#'��@"�)��\l 487��j���۔�M�i{���r�d����/�)��Z�@p��Ji�P�2WplΓ$�4����$D+� Ƥ�R�H���@?��+VD��w�z��"m��	�C��$�'��pX�+,FX� #U��q��J���a���z��	�P�P C���-��)+?�GЧ�M���͒7}�@ZC�0�����
j��C �UJg�$�aML/%zmH4��1Ou��H�oU����
"�F�z��JE�Д��u��t��L��t">yp)�<��9�q��h�p���C\��rΗ�=nv �� .���1�mA�<Y�H� &~��'�L�yD�!� �<i	�s��, Q��X�j����h�xy�3��Wh�h,�����D�i�!���J�鎞HҢ��0�<�*�DY����M�*CJ$a��n���%�\���@+��|�
3�~��čz�z��e��D��+񉈞I�⩊p��LW$KQ=�����I.� Y���</�x:w��
ԣ>��i�$kIVܳr@O&p�6�Y�`}>!z� �%�*XaB� ,"��F;D�C7�H� ]�a�nJ�r?,]'�>�m/rUƍ�)R�;ۊ����Ă2� ���O��9C�AX�.Ք|�!����֣�H�@:��3v�©�')ON?I�dҨm��SL~�=�L��(�|�R��_\L���F<�#,A4+���	'
؃G���2��>*�j �"�J�r��5p��~�a��9��f4Ox4��ɆOzx�x �A����V��		�w�����,���C�ɲ�Z !��A�Խ�����Oֹ�.և����OuV}����.G��I5��S�hu�'�ty�cAO�4)�s%ٓ]Lb)�'�	���="Ĭ�._��b	˓7y@�I�+7�dH�A���	�D�b���Kc��!�و7�!E�K�AK,\5�'��1�ƌ�8��S�'�d��J6GC�(��(�t	��_r��cۄ .�H�����7}�bF?3f)����yB�3\�4g�0&����fY��xbn�
7x#5��D!�m��c\�\l���@ 5VE�����:�Z��A�6J�\�(��� |����d��A"�a"F"��ISL򀡰W��8��&�]˪C�	�[����0�B�ū ��-�1!$?�$䌉QN��c#"}����gz�S$�A,s�څSW.6�!�dαG�P����T0/�z$s�����kL��`���,!�c>c�p�GC`V(`�H�\���9�D�&�T�8����2��mT�-����H�s�@I�E��H��
�)�h��Z�s{F��g=\4ҤX���1mN�<3����>����1ƅ����=z�]q�D��PU��+@	��i�">�w�7.d�0�2�*�S �����/@p��2���~�L�_��@S��4��ӧ�.�
���	1��1� T!�jC9O<�����L�I�"~��
W�ZX���@f�t;�B#<���'6�ԩ֢,Ϙ'�� �'�W�) @Ձ]�:�X�Oz�����:��$�MV�իV�W�c��XC�GȂ��H2UJ�;i�v�+,OJI�4
T#r�z�J�K<%��b6@�y��
4�-w9��G~'2���Cu�x�Jޓ�A{r��y�T
4�P��Od��U=$9 �V:۸O�ԝ�ֈS7[�0I!��Q�U���RM<�b��/���b?� v�{�OX3�j}�R�Gov풴)G�d��W�*�p����$J'p18��Cm��`�2gL�?��@�$n�2}Q>���B���P�W����>�ȴ@n���p. �~	:��+�M
�xR�Z$d|����l֤�|$#$�[�?I�˞?�nEH>����p��ߴ<j�E��lB}��p��Pf��#�N�1Y"��ēa񺕹c�-4+�|�Q�;M��`�'�l�i�)u�e��Gʳ~����q�[y�Y>��F�r�`hQ�͡6q����;�O�8��!��3���1�,T�=V���c����JcC�(s�N�Å��O:"�'��>��74B�WN34�F�Je+d��"=�$�����9�S�34t���E>3���E�ʈ"扜;\��CI�^U�zB�K!��i)��?�E C�ޠ�M;���?+*����<}J~b4L�x�&��ڴ(��̣v*�q������P�$}�ȓFJ�U���B�,6Qg�H?ar��'0y�[;A�#���#$�.��=�O��)��-��PK񮚧i�b���N�,�:�;f��c��,��eA�@F~��D��C/4��
�f����C��Y�\,U���P-���z��6Ur�z7�I̸����nHK�>����ɹT!����!��u!��
+E*����'u �3R�\s�ɧ���Ʉ�/| �����a���Hwd?D�H�peDe�]����`'b�Ƀ�)?���I'3�L���h�扡
�G$4��j\%-!��? e\���K�<ˎ��D!�)I�PE.�sKDy�b�!��ۉA����b�>�Z�
��ˮ�!��_�Gj��e�����ȇU�p
!��^�ܢ�zE@F Һ��f��]�!��7��=h���<�Ƽ9�T�d�!��<�p�c.چId�m�e��j�!��K68ʠE��!CRQ�㓎v!�D��F+�p@`$[�EH��c�`�S!�d0)QS-�1>�1B �!���?�j���@?� �N�K!�B+B���;����L�|�!�>^#^ܙ��R{&x���J�$�!��:F^="�JP�s�\is6��* �!�DߗjxS!�K�����JJ�*�!�DƜ'��§��'j����c�.H�!���B��b�b�p9��p!�$�53x  ����� ��߷RE!�ą:Cj��is�2	d��q�'	!�I�vI"wo�rmƕy@k�%!�$I�~8.h3�Kè3Zb�x�mI*�!�D�$/v^�D�6C3���M̓}�!򤀚cq�=�D��P	4dX���:�!���Tu.%�5�\;d����퓢|	!�D�e�Z,���W���@b���!�^G��J$-Y�ҁ�ƛ#S!�䔀g�)�ө�5�l�W�@�N!�䘡��舷�Y�LQ�wa�EO�%"A,,�O&��G! Rr����I(4����"O΍2D�º+� r��+]�B�P�"Ot��W枥y�ĜՋ��k�P=��"O���^&O���گ;X��v"O�qKe��Z�Q��ٯO5�+�"Oz�Q���d��@;	�'�\
�"O�9���ƘO��qY�'�9f
�!�1"O(}�gJ�%<z�(��X�y�Q�e"O>�0�̕�\s���t�Q�[H2ac"O�d��!�`��W��9@���"O�kş~Kq�랥t',A��"O�А�&����p�@�uF�}�"O�лm�>'$8hP�� K?� ��"O��{��� |��h�dd	5�x@�"O���񏏖/���s&d��o)�HS�"O� �a�d��2�\@�VE]=i�����"O���̔q:�qіF�3Qގ���"O���7	� j���{�BІD��yR�"Oj���i��
�2p�Xb�r{�"O\U�W�M"n��Y��I���j"O1xf�@>
�:m
�
R�,�QB"O����M�2�F� Ԇ��5���p@"Od����T�#��S�E&c��x#"O$x#�A����D[��xj�8"Oe��M"�5ɠ�Æ$wh�6"Oj���ө2A�ĢU�%Æ��"O��*�hK�}�Q��i[*\���["O�(�u���z�TB��>5��m�q�ɯÔ�����!}� ��g�:i���� �đ��X,���Ä�U%]����ȓH.%!���XFe���]�2�$�B2b�*ʄmD=�Ё��&S��?E�����LK���6�xˤ旷/x�ȓY�,;g��2H�ʚ�Z��8�����?)����$*�ȫ��C���y���<Q�(H%<����ER�hrX���HX8��Cd/b�T-V#	�Y�򠝤/9H��S�ؾds�0����%m��H���'U��	�a�S�i�96��ء������%GI.'TQ��pFm�v���ڥ�ѯL"��!O�>i`�$;~���ƎJ��
��^6]N�6�m��h��d��La7�� �D/S(f�d� ��p���t2t�j�<�}�]�>+��[8���J�<B_6��39�(��'��<PP�.?(.����S�$�cA�#EE��'>H�(����|&��ꕢ���p�l5Xbnπ:2�t����C�	+6���$i8G.u��(Z�x��F��=Ɓ�t�B�=�ԋ�Ɏ�$l����iz��#��*L1JT�`#�c=<�#���K8�PC�N��$����L/#���WD�{��0+��߷,��@�
���Ӥ�6W�\��O$�}�I72)h�@@>eI����L2|�\�O�U!Eǉ6$���"�VE�	ʋ��F�+k|�8��^�N� Uj"��8q����ws�ԫ�C��p=	���d˨x{���F$�؋��� 8��H��W7�ugd�%Լ<q��EH�e�Q�JN�5PFLD����Z��T�Bx�xe5\O��x��xTe�@	QM�mX%�Sb���X7g�3	�})��Ȧ�>T"����5��9��"��&E�M��Rg~"�?�R�eڻ=QҐ��b�(�>ԲW�;�)>�z��A%��k[�틖�ܗW;D��󩆝\b(�6e@�b�q���c�T(!6��	(dk��3S`�y�"�X���j0�3��yB^�Z���!*����bX�C(�أ섍!��F�΍_���{��9�^�X���A���'�?�E�X�oȅ���V�D s�ՙT�$��L�9�)!5N5�p\�ϻ+hb���E���T�h��um|eoZ�J.�hs ���P��=�S�r]�T@Jh�E�O�}�t`�+n�̜��D�RZjDӇo�3/&Z�Ks'�!�S<R��m4*J*ih,x∉&v��#��#�'i���韢����Тg�i`������v<4�P�C.?0�c%*�O�yb�K,uk05���"r��8��>�����M���'�ϟ1Lz$�	Ԧ�p��'~���7�Y�D< �F��������2l���eV�R�����^�V=��)�Ȇ�[f�)�E�_O��iI���O�O��a�!�����-�&4���^1��A��^���O��b0�c�՚�jүYOt��V�K 4RZ�`�kN�+�@�¨�|��Ik���� �F*[r ��Si��}`t�J8�hO|I����\�fp�PNʃ;����w>����i��@Ӕf�+�������m��Җ|��Ο�	�q���;����+���3%��0!�x���h�r�T�d�B*&�ǹ�*�F��k����T���;�ߡ-���7�̿:�dnZ1�;�-˜#uƘ�S��)>�S_�'���;W�C��0�5H2~�ԨD�L�3�8��C� ��Pm����
���Y	sL�����AF�Ui��F�x��2ߓvzh刜w$P�bIM�Ң$��(aN��"C
Q��V�d�E�O���uM��s
rI�r�_9m�8�y��I�c|\�f茢���SFK
N��ͧ	�B�!� /Z*��5�G�	x���'<hʓI��'���1�W|~�MR��x�i�C���б�N�#�?	����&�� ��
=+l�8��EBS�g~
�$;�0=8��N�Ըe�Їw��f��G�� yƱi�nX3���0����$�7J�8:���G�R=B˜Q�U�X�9#D���)�=�1OD��>� �'�n��柟8����ė�-�z�{p�F�����'�ߩ�|�ێ��H���8��	�h�G��QrE�;y%Hё	�����l� S�9�HГ1︤����5qѦ����Hu��W�I=n)� eEL�)�t� B�-=��q��"v�>�&P�� ʓ ����9dEU�P�(����u���O�R���P%5b ��ѥW�z2���]�TP' ^�z$�3)�GR�g̓4�D�ۃ �6T�|�Eyr	�DZ�P��A�3�M�7@P���C��{��I.}bc�=<���0�Y��ЌKc�BH����"�IӚT;��/�d�R56
� �Ix�B�a!A˧��/~��z�ȉ�W�Tj �<�����Z�g�O�9�0�qe��7�: ��S#G�B��6�x���	&}.,�?ͧd����E�C-�=���]o���K�N����:Z�y ���|^`�%�:T;$M�d/�M�r��6gK�[��R�B�ʟ��1���25@��T[	XΞ���䇄"���A#E|6���^�~I*�Ĝ/Q�Re�cKi�$���	'ɺd3�Y]vU��7V����J4g�5��W�H覠B�nY��ARH�=�}���%?��ɂ��EñŌ%�9E�@X,y��X\��)S怈�sԎ��(���P�Q�x☡ P�Z����~)�G�Y5D@1�h�-m��Dډ�OvKAp��H�veE�
�� �+Ь7qЀEO��~�Af���4�D	�>8�8�*�?�c��)5�ѱg�$U�Ue�y�J��?��O�j=��k�&ɪA6��~�Vg/:��h��hT6E����r	�)u&�����y��).����g=��D/�]@�`Z�	|�,[B���	��s��Ԉ�A�t6Oj����X�H��g
4��0nT���HV��d)fT�D)¦A�๑��ޓh���3�F=D�2LZ,O� �6ƕ9| P��a 8�$�󜟌[E�R�+�~��ã��UUPuh��ǘ��I99�*���bǟkhX�u�/r�x���X�끱b�fQ��C�+�H*�J�999i�d��$˴���b)T��>�O�rp6���>�Z��P�FI�B@؆��)\��(�A��oul�p'�-Șï�Tx�㫑�?�0M�����?)g��c����U;�^\#�Mٗ2�xx�=Ѣ�{>aCg -� �H|zb�S�bp^l)U�6��ق$[�g&�*�͆re^!`Ӌ�/L꠵8�Z���].6 ��R�).�1�.MR�2�[�fA�1�x�i:3j�u#a"ӟ����}��KP-�5
[+"���U�B�X�m +���HB�;i.H�*��a���'n�h��I�P��|��З4���A�O�����P񚁁��=U�aq��O䁈��v�h����.Z���iI���:�č�1�x��%F��|�m��g��i[���$���؇^qO��YO�`Y�r��X8�m�q<��B��e (#1f��3_�,�+d!|�"2#�Yzse�05��� ��ԟ���5?SȌ9��-l]�!��hA��`�Hj�8����Fn�)G1�p��V=���)/��C�W�LU���q*q����b)<P�`����<�C� xP<�Q+C�W+.d�Vm�	d���$��Ry��R&+UV�BeH֨�b��S�dL޸(���Bw$���t��A90aE�$Y]��%!Qw�';$%���?ra���	2�Z�Ol��v�ùY0����*ڄ_ˀ}I��O�̀U���Q��[��B8H��d8���V�,���Rt}��#�܃-���`��g�`s�O�2L�<�� �,f�qO�s�y�b�,i\j���Ć?(���爥oi�����JHm��ꐯ
:��)�j#<1�� F|T5@FEɺh�^%���V.� �=yr#~>1ৢj��b>�!�2�^�A#�F.L��CiZ"`���)�qO1�w��Or``$8rhxI�]yp��"Eߕ=�6��m����H<,�I�sm߅M���S�tmוi�xD؅�{5�)�%	;ļe��/�:)��͈Q����g�2t���Q#�Ĺ i��"���r��	u�j9Ð�9B��5 �
.\4��	�<���R��vh��'���5�"|��)��L�e斅
�
͙��ͶF��%c߄�nX����	y�mi�))�|λQ/��˃��wp0hy�D�<���N��\X��r�vy�ɇ�ֈ�M%��$db=�"�����P�⃊rJb�����Ol�����'�H��_.�7Ծ8L�+�'9h�eЬ1ɧ�i �=�(�0Sd��C	l�ۧh�;p�4	��� ��T̖�=
fM�/_�@��Ӻ�O��	��ʁEl�i��K�&�*eh�)�4�B#���1.��F[~I�N-w�\��wAǄ%�c�퇤`�j$`�r��6��"��8E+`��C���a�B
� ��'� A��
נb�ܠ�fE<�.�!HO�\1( n�-z�V�7�B;bP��� �c�S�T�wv��/ϵ>-��B��0*����y�]�ת_A�ď R
���^���|b�I�61�� �D%6��d��$�&Th�=A�}>���Hn��g?�&��ٔrG�+����X�<�M�"C�4ٳN>�O�4���!��x��E�2���I��K]/]�xyh3�.s��p:�B�M<���A���r������	O토�af��
u�R�&d����r!��3�^ѵ��ds%�C?�6MǾݾթ���,.�}���b~�.G�!����>?�x�"�� �?��d�9�p��`�Y�+а����^;!��߸	��#�h�$Î�{���,��t��O�J6�Șw(������
�������^Đh0ȉ�$�贫���;EU"�mB��	�>� L �qZ��,�6U�5�q_>IS�wYZ�X������q$o׆|���D��1O��T�Q`踥�[=rvlʓV��8�LK�[�.�s���S��Z�:�D[�Y.�q���%P��e����W�O�L�h�i��O��YÐ��";h��cT�-Q�P�X�4+�2�Y`ݴ8�A��U+|%�T�`C$?���!~�!���N�u�*��%��ݦu"�'� @*��4O�?�Ro+��<��m�n��l���%]���"��VZ^����@߶Q~�	S�O]��G�V&|�;\|KG��zP╣�(Q�X��O����#W�"���K?��~Bu�՗sp��S섐M�����?̜x{� |�		4��8��&,8��a� q 6�?��!��[��p��\,%�<#A)�Z�.㞐��?���`b'��[n"a+5�<�p.&=�R�)r͟c��c"΃Og�a��&�bW�X3苑~��<�|����
{�)qCf�7dq�9A$#N;���㨋2w�6|A��b Ȋ׆PH�I</��4��x#�� �ʭ�E�'�"-K�4/���$C�3h�秈��e��J6 ���D_�K7�yP -�� �����~bA��hY8���?�S��-*�i��O�X0�G�ӌ.��Lj���t�҈;-O�Mp6�Y>Z���I��ObN�`Š/� ҵ�"DK�F�s���J��l��'\�(JD`�@c�7HN!�4cݤ���L�|:�"�d��]>�����R�;��1���09b������)-0�H|�Q�/,��P)��;Gf�T� �B-����`�2���q`Y%| �iL|�<��kP�j�%��M� -���2Iճg�� ��csӶH�-�� �8rd��~����ɓ� ��!Y�����T&Ba��=M�X���( 
�\Eb�P��a1�^�T�(�p�A�@��qBG#���k��K�X��q��VzxO���  3e$���i0b�`K�CH8�ē'�v�	j_�,���(|�y�c�  ��S��!0a{B�@'�"9bf'ǘk��`�'�Ïs��r!�&�r��Be�}Z.⟌�,�klɆ[ꌠ����.����r�T9h¡�DMS��eK�!ݑtnn���S/Xjj��DS�ci��"-G�0��Jg"B8U�M��#�:$
��E�:LK�E���d���M�˔D�W�̴C@�!`��X�����E��%��1'/�t���)v X�s�,��(�I�9h�P2��!�~Q�f+ٱSp�O~P�b#ɑ�p$��)e������!5�5za��-2 ��w�Be��P'fJ�WƊ٠%�_؞���J� n����i� $b�"G;+�ಈNp령��2,Ok���Ү���>.��c�  �i�!��Ԇ;�¡h��:�ڔh�O݌��	��hW��5�58��ޅ0��S���5��{W���p�X	�$,ŵ}oa~��ʞw"k�wbP� �&S���+v�˄.2Ɛ�u/�Hɧ���DQKTr��7b�.��ŀ�	09)!�I�=Ŕ�q�?%��JU=zD!�D
�k�E���� f���;�'5N�!�d�>O���k���9�d�;d!!���dV�ѵi����1aR,
�!�d��L��ݹ"ǚ$u�u��d�"�!�d�0���;����&YpXiGD�)9�!�DӋs�A8iהv;,���"Q�Y�!�$/~l�\���9%J�y tL��)�!�d�rUJ�!(�(JI��Ӳ��A�!�.�>ex�@ʙg>B'�O�P�!�$�{���Pq�Ù=
%��1M�!�D6�b�XЉ���,�rt�OIZ!��Z�/�NP��JKAs�H�f��	X!��B��TA���,qp�Eb`!�>)@�b�㕭d�e�'�	d]!�dD�}(�ؒ�����P2�"W-l!�ā$Q�BQ��Y:"a)���Z�!��q��\ȵ,�2�l:aaG%"p!�$ڌnMf�i���bH�� ��!���d�Nݳ����ԠJ�o�>�!���UN�<҅)fͮ$�		�!�ߊV�V)�ܢ1e�$A�!���xjd��Ӕ׼d��VF�!�D�?.$�US��ȕi�Ʃ�%���!��Z
&T2�ŏ�+�B��B%�5MA!���K� �`u�Bz����ϧ]�!�d�q=D%�"�"��ȣT�u�!��*9������&��\�6�ϩ(�!�G4k�5���	�4�ʽj�@v]��ȓ4�IK���"H8l��Q͞�n��T�ȓ&����#��OYT��5A��$��4��@Ȥ Ŭx|m �k�v��	��G٨E��V&(��!���JFje�ȓK�����&J�3~ `��'��:R�ȓU�|(�-II���7N�3tt��ȓv4@:�čBS�}8H[O�V��G�pzP���X7����K> ؤ��r����0]I��Մv�&��ȓ ��́�A�6'��49矩(qx̄�~g��R�V%u�-�"u�т�I�<��FQ	`���Q��8U����N�]�<�c��>X+��%eK�p`W�X�<94��4+�U�ca��G��1��N{�<�ƯV���̐%�\�����t�<� �쀇��#G. 2�h�0�Jl��"OR����}�L�	V��rDs"Oּ3N�:��a��A��r��e�C"O�����Na��qb�� 8*�[a"O��ҌL�`te�0)ǪWF &"O*�Q�|�
� 5.�>wH�d٠"O���#����Чn���q�"O|p 1IK�lG�`�'-.r��4a"O���=rs����e�E}�<ɶ"O��GZ�&#���_0���"Oir�fj�XD�@4DR�"O����陀(�㐤�_)d� '"O�xAq�W���j��]�E� �A"O@Mʐ��1�S��uC�L��"OX�p�����-K�a��m�pPr"OtQ!�	�4Vr`�)2&M��Ncp"On�F%�C��� 䇤OWjYٓ"OU���	;�P��̺CA-	�"O,:f��c�6y(wCN�yʞ�:�"O�X��tk���&)��!�"Ot�Z��?2��Dc�*���r"Ova$b�f���Q��M<Fx��"O�\{��R;a��$7
��Y2|�c�"O|Q�p��{C���@hCM�4�F"OZ�Ή�$ږ5�D��S.,��"O���H���H�U*J*�ّ"O�X��˒)GC
��R�P�/����"O4�ؤ�\�b� Q����i"Z���"O *#Ɂ�hx��6��_<8�@d"O���b��`���
,�l�2�"O�W�!<[b�8�&C�x� �i�~�<��E� �-h�U�"���t�Mx�<��H./���UN�8Po�x��Y�<�s`VZ��;��4k��Ӗ�FX�<�!/N�@F�Sg(�$i�2���Q�<����A/:h��F�� ����_x�<Rd��!r�����R���Y�*�_�<�&$�1&���@_�M��p�M�Z�<I�#��a�j�.R!�U	a�<A���Z!*b/E��j@*��[�<Y6�Zw
�#��͍  �MXVB�m�<R���"-�|#��M�)�X@��B�<y2l�=F�v=��=fv�ۥ�^I�<ђ΃$E��1��!/��(k� �C�<���Xd��y�lԧw����u�<�@NQR����T�I(2��#7O�{�<ӇU#�u�!@�
e:�&�Fw�<��$:9<1�NA��H�� bB[�<�t@ z\��#��:�9�&�TS�<�Rt־���D!�ْ�oQ�<95<W�,h�CG�B!0a�N�<Y��3<D��jܙ1�����N�T�<�pgKi|b8��Й}I�ț!kf�<��GΜ
�\�Z��dͤU��V�<�3�"B�z��%�אsޚ�;�*�{�<6��,�
�S#.ёg�����B�<����	�$�&`��>����
�@�<��F��uh�ҧH�/�<8�vLQW�<�@F��s`��,9Gf�Z�<��O44��軵��!Ap� ]�<)"�R.i�X����a��Dӕ�X�<yf@�6H���k#P^�d��O�S�<�@��o�ƙ��N�$:�r�E�z�<��2�e�t&�k���ԍ�P�<� ���gl�%��뎕vQ�ii"O�|�TA�.*ۚ��t�^L���v"O��u�и����B�4R�E[!"OHls�Y|����ǿT���0E"O��C�3Y/j4��*�"d��a�U"O�����+m ���G���XQ#"Op,�f	�7	�`���A�1�z()0"O�sf�r��2��6����"O�HHT�_6K�����̂�� ��ybk�jM�T�@��!?�L�f����y�k�<K���A��@;�H�%b�y"��7t�`�"ԝ
΀Pbp����yb�/L��0fI�4Ϊ]p����yb�0*d���E���(�B8�v�K�yb
�;j���V��M��xf��yrW$}����QH�V�z@G;�y�HD:(��(�#k-I���R�&�#�yB�_����eӫKy�q)�ʈ�yrO�?~��w)�E��I�C��(�y�j�
⠬y���&)�(;s
���y�-ׯj�
9{�ڤ'?���"���yr�E��h@����8iR.���y��I�6�����'��q�=�yB��3p5��Jfj��z���jE��yҊ��JH�x�"���Щt���y2m�� �Pp��u��}p%��#�y�E��%z�`�Ê��y#��B��*�HO���d��_C�a*��ܹKj��N�/>!�$�{�y�q��x��CΕ!W�f
Op  �nP�k�ƁP�M�1+��5R�"O���1 ͌Tu>M�4F�?H�hiG"Oډ��GN8���0��<Z�"O��֨�&؍�c�y�`!�"OD)8��N4/ �-Q��-S"ON�Z6��"���S����Lc�"O��s�K�L�a�����ZD�A"O�\8��4b�v=b"������A"O*D�W*J�H��My2�V��Lei0"OH��V- �]����vΌǖ}IS"O�tC"&&3L��c���9T]:Q"O����A9\�cdoH5~��""O����GV�D��X�-��}R4�6"O�<�2
P�4�P9�A-PW��"O.�B�hK6��a]iyO>x!�Ҟh���J՜5��wb�#(�!�$ʣo�f�{3���I<�!ā�5!�D�D$�a�2��'9�� � �!���X�m�#ιE|�2��;Cp!�d�/n3�������	0�L��wR!�$��c%
p
H�r�.�	�ִ/'!��G�}!���� )�aү��J!�S ?�H9���x�ll�����(/!�S�-��MY@i���3&k�y%!�(]�̢�G����Q�@H�!�!��T*�����x��5i�E/�!��G56@!zäڦz�>���ƧF_!�U��d#�,O�� &��F!�?��Bݸj�0��#d�)!�DL ��x2Q,�H��i �,η|%!�d�Z�~����&��Y�RE_�5$!���z�'IO #��Yy�S�@r!�DN?�)AA�#_+bi�ec�  �!���T?`� �/N"��B�!�D�bp�\(P��3�|ñ��}!�� �m���Q>K���i�I�.|�6M�"On�)U%M7r ��I���"O e�`��l4pq����;�,�KD"OpE� �}l��S`	'9���A�"O�2��_)]���c���z��"O���bB�	���
T�L�bs�e�0"O��P�Ô%n�LpW�a8�ف"O|0�N�~�ҵ/�f�Z�J"O �a�:G�"�����0	;6"OdUbw� ��=KG�[C�u�w"O�I)�����Vn�C�0�i�"O��2tem��qk��H�L�K�"O*��@�5Af ��gEP�����"O��ԉ��c Y0I؎����"O��iǪ��Y������\���&"O�`�E�m([5eG;W�Br�"O��2�g�2���s���N��Z�"OB0r`��)6r��{�*��$�&m�G"O(�l��
��L3���":�	�'"O�0�j�"h�^�����$t'd�U"O* �@'P"���߄O
��E"O�a�p,;s�%)%ΠR����"O�h��^��z�mD3��u��"O��i�H����c�X�O���"O�,��+��8Z~�zaˆ�@�|0{�"O H� �0��SGJ4%��]�"Ona�Ν�N�t�v�I=�`q�q"O�8���N�J�+O6���rd"OX�ƄϩYي5�El��Z�T�c�"O�Y���ԃr�� kI�e�& ��"O��3�/��K�p)�J=j��h(v"O�<�E2=���a	W�lx�T�%"O���(�2tǐ���FɌ{�\�f"OΙ8�Z$>��Ja�S�t�Q"OlP�q�a;�Q�F�i�邢"O���G�A�T).`g|sXPg"O�\B�+J"F��9��V%5��D��"Oz��d_q�P[DK��(#��)�"O�q�`MLzb�*���� 6x)j"O`��bퟏF~�sT�	p"����"O>�ʥŃ3V]�(�(��A���"O�p	��7Јu9%��S� e�"O�\ر,��h�Jhس,�$"�t�2�"O��éR ҴY��ɴtFaض"O�-Z��]5*�PϾk�
�B�"O��5lVS��!�b�طa��h�@"ORa��W$R�0���mF�n�~��5"OX�a��Ol�J���B�Ш��"O.����#j��X���g�;�"O|��iTB��K�.��b"OơC��)�|PRLӆ���*""Ob)��鎜v %���X= %#F"OTM�p��	<�-��A�{� ��"O���v�ۆ�ٰ�CR�L���"OTp�҅��莡�E�Kq���"O�ii�����dR&�J�0�R#�"O>Ya g�+~���K�]���A3"O����
�'�x�[3��i��]�d"O<�@ �߽�ԳҌ[�$B��b"Ohy�m\
V�>tsE,X�jt��B"O�����Ck��a%��`�M�e"O�e�f�9<���!K�d[��"O�k��T��!���@�O@Zͩ�"O�lڶ�@4z�ɉ���]t=R�"O� d|�7jڤP�*���
�G��"O>}:�e(x��*ϯ4L���"O�И�/?�qhej�81��´"O����A���%��. ~1qw"OZty'��-5Fa�����-D�0"O"�ʓ�یo�"����$8�1#�"OĹ�ƦM;=����L�I�dQ9�"O�5cٴ�c�kʪi(�	"OJ�C�� b4�94
�Ze*�"�"O�����l����W�
6W֜q�"O���o��p��đw:<`�5"O�	���&e����S�l/��c"O0d������3q�5B���"O�ݓ���;~�9C,GŠX%"O��Ңh��\Ś���6WZ��C�"O��	�d���ˣ)+�x	�"O:5�c�&yf�*�C���I"O���5� 3X=*���3�f9��"O"��aC
J�Tt�A{�Pi�"O��0!
��P�ـ��'.a"O����ɊQ{f��G�	�r��"O�y�fC>���26-��g&HQ"O���4�ip��mB�8��� "O��J�"��>�T�K\�q12��G"Oв�	F=:,�gKԷ[3��"O��XV��!9IB�R� ����"Ofd����j�@q2�*�7��
"O��s$Ë>0��� @��UH&]y`"O�x�ؑet2�puOۮc���;�"O2[d�7-�4�н�DbQ��oܓ�hO�O%�8��b@ ��[�r��tk�'\RA,h(�P�,X�7\������5O�=zv�F.NYfd�"ѥg�dbaO����[�5�q ���WZ�Ĺ4�4D�p��GZ(:�.jX�	d	 D�X
��N�<���e�dt�b�I=D�TA�A�'���1���8��0�%D�L��KDG%cǝ?Wd��M�ybcO�eƸ��
Qt*T=� B��y"��P��lt" �n5R%"�A��y�a[�5*ܠgb�j9
����?��'u�,��h�E*�H���A�0�
Aa�'��x��(U���B_V �{�'L��qլ�5�����ī�̀���(Ozd���H9rI̹x7�[����"O`$��ل���� C��ǖ��"OT�5�!&U�逫I5L�"�"O4����,���tD:{���KW"OxMA��N��ؘ�n�%����"O2�Q���'���
a��G��	 �"Ob�k��O�$��I˖��0��v"OT��Ǒ�Jp�8��f���u"Of0h����:� ��7����"O���EQ�F�~�#���$;�"Ov\!�����d��
�Cb��"O0L�4�[�u�6�)2�_7(N�k�"O.�('%��TRrES䦆�h��"O�i���;(�cd�ݾn����2"OP	�$B
7 �ڲ��%r�:�"OZ�2S�K��@� �.�"��d�4"O�-Ʌo[�|h�bNV�y�l��"O�`A@ŗ;:�D 	�OͷM�< �r"O��X�J��f��)�ōK�E1D�s�"O\�!)� N����j�&%ڠs%"O� ��8'h��!ʃ�&�l}�e"Ol��'D�tc��Re�=��"ON<
q˒&AI�M�8�&�t"OН�#��e1ldx�E���%.���yBHZ� o  �P�:�R�q���y���<^���k�ŔT�Aɟ�y���`�W�JuLl%�Fg/�yҎ;Kg&�Q#�i��U�_��y�
4"�u�lDd�D �$�y��u�H��c�F����Ը'n#=%?�tœ�h�������{�L���?D������p,��KP/q���s�O)D����K&8� @@�f��
�U� @)D��ؓ�^��I�-�E���+��'D��UC�!!���F��*>��e��(#D�X!P--t`Ĕ⡎�2Eƴ���3D���6G����w�D�A����,.D�`d�7wQfi�U�@<y�2Џ-T�h�0�9;�����	'T�,�"O��K��W�C���a���%X�*��r"O41�tkL���#��W�2t��FSCH<I�㉎R��"�M��bn�`;U#�Y�<yQ��|(T����b��F�S�<��ګX��x�` �)_��)��K�O�<��gÏy�:�z��R�=��J�<� �H �Zڲb�#a
\�q�[}�<�˅��[-Ffֈ�g"�}�<I�����j-�B	D�Y@�f�`~��)�'$O�q�Fa̕Qeh��©/�؅ȓ0�j�u�T�h�l���Ɖ7�B��WG��a�"ݍj�����04�Ą���q�V��	��i["�_+A�ńȓ��h�t�6'�|���vZxхȓ��zV;��օ՜a	���D�t�t�v()A�U�(N��F��1hb�n� '%�R|��'a~�D�?\Ш�������aG>�y�ڹ��)��+̜�� �D� �yr#�I�lyQ�O� ���ᛚ�y�AA(&@D��g�eDukAH�+�y"dӎ)y8���1J]��X��yBƟ:E�諑��LM�5����yb�� ������7k4�X`��yrG��_�H�B�aNt���mV��y"���#���h!׾h���y��B4��.l�YE��~6iK�"z�P@�ȓf��U�����g��a�v��7GՒ����*h+`�ˬb��b�kH1c1j�ȓ@�����Y�*�|��0`Q�q��ȓ5��e�&<~v2�zse�c?|��ȓk�>u��J���@�z.��
J4�ȓaXKW ��h�jr�F�kʞ��ȓ`�:��X�T��R�/����vR��+Њ/cpD��#�0,� ��t���ۤM�>V���"�b�Ubj��'Vў"}����<Z��2� *%ҵ#7��L�<�YI�"�
2cR���cI_�<�5h������Ά4��Y��p=iҠV'zC**��	H���qg#�L�<��\���Ҥ��R����FXG�<�$#� ^'��9'@D7E�pX����D�<��ōfDh�� ѳ"{��� �D�<ᔧ��%��L����f5��J�%Lh�<����!�����mI����BnRe�<� �ɀF�G8�hTk�L��|@1"Ot��E'Ȍ'Υ:v���p��%p�O��D�h6L�s��9	tL2mF;!��P�$�c'��+p�ꭻ�BɱE�!�d�/�h@a���Sp��� ^#|�!�d�7m|����Q�B�`��1�֚"!��>b��ipQA�<_�Iуj�5�!�$`��׌ғT�N�����J�'�`�gM�D�@���*�5����'��� �c�F�z}(6�B�.�P���'S�A�䩈65_,���:)|�`I�'���b"��&O�fE�A�^-!à�S�':���GdU�!�X�����N?zq�'j 51p�@����j0��<^�y�'ݖ(;sC�m�H��,�PRu{�'�9�t�T�V�zu��Hީ@c����'K J3̈́�?���4��&��  �'8�9Î�sL�V(��1��M�'vўʧI6�$7���v'�DRÄ�
*�a��~�xE����m\�I �L���Fy"�'�"lȥ&ɣH��D0�{�,8X�'��mc��U�d�獓m
���'���6�
��j0�S�o��X��'��@��#x �
2�:T��'��	3ʨE�^�@u�N�h��;�'Ԧl�ŚA?��{5g9���[�|j��Ќz uìևM1�Ѕ�d�yc�gNU�a:F���@�����UVd@jc.1�J��֥�5hrm�ȓuNбj��\�i�gjJ<ea�9����=�Q�u�JE��e�Q&���wު�[Ќ�&BKN<'��Mj��?D����/�!�P��^�h"��8B=D�P1 gN�m�F1�g�@h�%�vm9D�,��ɲtD��%�+���P�"D��f��1:��� �cc�p�""D��� H52��A��
I�r�g"!D�ܱ��߁G4A��'^4�FF?D��!�ρ fD�p���T*����'?D�D��ET"cG���������<D�2&b	��$��J^��9D�8�g$�!���G��D����5D����	00�â'Uy�����'D��35��8}�u�e��(w6���%D�\�*4ufp(�ɗ?8��(��j"D�@Qcf�3Xa*��X�+�����$D�4�jV4�<,h�H�P26d$D���d�(�Ѕ�" �o��]���<D��9�(\+?�p�t C�*Dy��:D�`Ƞ *Z���B&�o��@�:D�ℊ۽%Lh|1C �6+j����g4D�$�$�5!�Fe�J�գ�2D�0qd�/�����	Q�D�1�5D�T�6�T��2�KoY�\�jq3�f'D�D�A"�>�~R�K�1�٨D�9D�\#G�C�LJ��È$�%y��6D���c���=��g%T�K*vQA6D�0�VG�a.5��҈mT\�bc�4D�$q�O��nZ
���f�PJ�a1D�䨂-/t�NE�@ǒ-�FE�4@.D�P��U�{qz�C4N�1r������1D���s�LQ��T)#��(e�x{�*D��觪2l�:w��|m�@ Di>D�\��$�H����G?T3X2��1D�� ��s��Q�r�0C�b�zCʈ�G"OP���l��5sDb�#�@��"O*�qC�;L/hA����4"O d1�(�0w�DJ�Y�=���E"Oz�"w�H45n�BV�'��K�"O�m�fʌ+�tD!�KS�-�45��"O�a�BٶQ��ڣ�J�.�p�2�"O�9�N�
(��c��B���"O*E�2��5�'ߪA��|��"O������Hl�e����S�x`�D"O"̓g@Ͼ)"��jG%)�&�2�"O�t�SEJ��`��	^�cp�L�U"O~�8ր��|�����Y�^�"O���'�_��k�G�.|E�!"O�M�%�.+](T(635�8T�"O�,aê�!�n%�%����=ɢ"O��he�&Yf�R���7s�~�V"O����M�S%8�%`}�ț�"O�3R���f Z��U�\��&l�<�PL�{��1rc�3�R)�f�h�<)3O��(���4b\�I�L}3�Q{�<)!�?OF�I�lծ�.�˂y�<ђ ��E2�x�݂$��ْd��Y�<1 ��,��ip��ȇd>��ˑV�<a憧,��A�!����X��+G|�<�탳 ��{`)�>Sr�ջ5�B�<�ߍ:a�క�57$��HPE�t�<�WCa4����/p�&9bU�<�oV�d6D$�4)�(L�"���̔X�<q卞�h$h�d������!���L�<�J��xH��Ba^�[�.ԉ��t�<�sb�>FWz0���)9[� �$	�s�<�2K	8G^��q�Ý#���ujw�<��Ϗ<D$�L�B*��0D�R �
h�<1�(�n➵��X�:���'��c�<)�b��Y�L�8��M=MF(���g�<��%[gꪐ�����|
��q�S`�<q�+�'xƴ��A+}D���o�X�<	i�$4�����;i����&�I�<G�Ёv���㳏��*�<�! �F�<y�o��T�9p!�����D�GG�<�dşh�<y#�ڦT�PѴ�j�<�3�W�S�9�u
�g�̰ �b�<1Ck�Md��d�ס{g|<�ĀF�<A+݋#����4TMdV'�J�<��K<Q�=zW�2+R|@	u��Q�<�j��xbhh	 �+,�����Hw�<y񢏝6��i��n�2M� ��q
W\�<� c
� KV�E�(�j��%U�<���� �(��C!�R#$�U�<!'g^�t���#�*3����fR�<�q��y�|��D)�� �����@[K�<�p��6�hi��b�Y�Td1l
D�<Q�&ń3��3i^z8Hm�dK|�<y�Q?K��ad���5j�I]�<	$���z�f	s$윅6�4�T$�M�<	�	�x��:�(�>��G�b�<)����$y&4��mBy_�؁QEa�<q��[?h�+D��b��,�2d�a�<������^X��ȚB�yR3�K\�<�����#�@aِ�y@N\�<Q��ąZ	�����]{�@ْdES�<�ЮY�9�Dh�-Vul��DS�<qr)#1��²E��C�P-�D(�O�<� ���N�br���,��yV"Ot����5,}�1+DK
.lc"OX�r�����ƨ����4R
�1�"OLa�ԩ]!W����]=?�� i�"O��FÇ�����)�r٪�{!"O�#��g�S�iW8|5��A"Ovaa�*N�JiR����P)"/��p�"O�8�3/SQ9�BƘ?̴�@Q"O��SbdlU�s bT;Z4�2tAP�<���6V+�M����'�������@�<�tE�[����a�X�0��~�<a��M�,Ų��DBʜP]Р���Rz�<��{v�E(��/O���cs�a�<�dZ:"����4$R�2�@�`�<�d�5�4�� )�,_��ȡ�D[�<��4,�҄�N*_��큕(�]�<��jԚ7
��Z����
;�T��^^�<Au`�>J��ɫ� !e&�谫V^�<%�R8N\�e�qiI�H����0H�X�<Y®ɢ?�A�H�9�L�xaN�W�<a�H�j�)�L8
�^���P�<�@Ί�0
��Gǌ�T���q�e�<�gE�:�b K��>4��l��A�l�<�U
��Qf� �CN�"�̸�˂m�<Yb�A�U(�����H����s�l�<!��C1���a��~Q�h{S��r�<����`���"�q[ڕ*�n�o�<�7f�~��,�Da_g���5��n�<A�d$aS�)�#Ƌ?wj�Ӥ��T�<� &�z�>g��A��Y��I�<9#�:|�P�ʔMl��gD�A�<��EW�68�M;��R�v���P�|�<�)�2:��K�WcP�aa^�<�%k�0���cEm�l[�)�jBp�<!ڊD4M8EM�&	�-1���S�<� i�!g�t��V����4��BX�<	Bh�('��1R�+[�o�QR��W�<���L5N�/^��dh�U�<�N�2��M�䢅� r�8H�ŖV�<a�J�6�0��c�5~�A@�E�T�<QE˄����WNZ^.�I��z�<a O�I2Y��[r�h� Ap�<�&-��=w��ЌErÃZl�<� ��%{*�(���*���{��^�<9�C϶{��9S��M�����FZ�<�A��]@�7ߍ�x�J��U�<��D
J�"�81!�%*p�Y$�=D��o��=C���b�Q\��	�'�duZ�NX"n);�Y�R5v�9
�'묰 �C�N]��P���I��'�^hj�/
-(��i7(Z=u����ȓ�BDh�hB1!BxS�K�7nGh-�ȓG0P�q`%Ա+�,���@��@�N���NO��Z�̃�A�P�
3#�,u���ȓ���Ź_S6Ы�&�$�l�ȓ(0x�e��J�n�#A_ JA��>�ص
柕N�ԁ_�4p���L�<��J�;ÖL�S��{%tiǑG�<��	�!@�3�疳P���0�\~�<I�Z9`�n�)��P:}(�a(B�<��/܎�P!�Ι-fM9V��T�<�P�K@�&i�գʒu"�@q-�Q�<�d	 r��T��l�$tNb(jOL�<q���$LjM�eE�#gH^}�#��r�<�  ��΁	t0h���(`q�"O�=�T,ۏdG,ɓp��mGJ"O�к�4̰h�mS. ]!$"Or�I0�Q�&
T�h�.
G����"O��b�E��64��U�r�����"O�3��Y{F��p���R	�c"O�FJ�$N�l UBN� �T呅"OR�k���+ed5���W ʤ��"O"8����a�����.� ��"O��Ӆ��	�~{�(�6iU>X��"O � re�R8���R�̫d?�3�"Oƭ(pHP�iAJ�	 ��|'�}��"OrQ"�)�R��;7��'*=��"O�,9��	�PZ����u��"OD5�Rn/x�����F�`!�'"O�DC�.U�h.���1 ?n��4"O�%�=f
^�
6�[5/���:�"O���3�B^�F�
�n�N�$"O:p ��<mc�)�Չ[>K���@"O�E��ʙ�ܑ$#%x��r�"O����7"/�H6؛4��-+�"O:�� g<vLLeq�F��tSU"O���b��&�|���|�n0�"O49�v��6O�)ɂ�Q-�l4"OD������\5��-R�k��X4"OF4 HI�V8����7aQ�\!�"OD���@ϗw�pE��
X:%h�*�"O�T�r���6���A*�*FeR|�c"O��B�T=t���{p�>qa�`�"O`a��Bi�q�� Dg5\,k"O2���g3ce���dv�93"O<=2���U\� @E=z���[1"O��K*_�>��X�Uည?�K�"O��� �@�2L�9���J���2"O�
ʁ 0��@�(F�*p�,bQ"OtP�c�1����w͡pH2-��"O�Q�NȽplĄ	t�9{D"E`P"OR��׭¹4�:��c
�"���"O��� ��|# YYԈ� k�ty�@"O�@Z�D2��@�'�����"O~p�R�^��&�0Hi#�"O�t�cO6>�I��F
���g"Odܡ��
�$��\FF��V��Z�"OJa�d�1�&D`&�������"O��4Ɯ�Wt�����IS&"O���́�N���3��9X���0"Op�x7�D#)�2��a�A%[�|@�"O���cM^�n��	+�Ɔ�|�"O�������68sT`ݔx��y�5"O,���HU�\�>�H�ą4 R���"O����$^�2�öC�XH2"O� '�W�P�K��2X�>�p�"O&�3G��Eإs�b:��A�b"O��'�0�8 �A_�u���kC"Ohٳ/����IAq.��Ij�"Ou�f>;l �b#�,&�8��"O���,�#M8��92m��p�����"Oj����l�p��F��Qi^c&"ORi(�^к�B�E�8Lh��"O�ِ��>S:�)􄂼L=�E��"O�,�a -:�{�$ɣX����0"O.�R�oC�n���Q��ٔi�D"O�Xg�0S�X���ES�:�*�@b"O�<	����tt�qS���(����"O� ��s�� � �1��N�j��R"O�U��"Q� �I�a�i��ej�"Oƴ�&�}gNĪ��@� �"O��Y#kB
�FXx3⑬`�Y"w"O6Ԫ�L^�.�8� ���y��"OJ��@FC[p�@�D0({ M{�"O֔s�O�0��]+���,ql��"O��
�G˙F+�5CeO��V�}і"O�(R'���D�0���P��T "O���@��/`^��J�#�bPA"O���Ƈ��:`�I�#�P;"O�M�/J�e�tな�.�~���"ObȲ�AB0�v9�b٬�y00"O�9q�Q-(X�1��1H�0-A"OQ�0�����GK�bW�ˡ"O\A��e�u4>��d���;p&8��"O�u��1x������MF�,0D"O�3��I~����#�e�]r�"O�M�P���k�h��R�#1^z�a�"O�R�&�-5�����SEʠ��"O5�'�ȝG)�Atf��4\}R"O��C��ΐWxNx2&U�&Ɛ��g"O�٪i��o���b��5!�8A�"O�uc�G�V���H�8i a��"O�ii���X��eR�H�J���"O�e�\��Q\>nx�4x�#��~5!�ď�"n�٩����Dđ7��0%!�dSD,�1��!T.�C�g@7	!�d��-��5B�@ԲR�8����f�!�M�iN�)+H���dIR��4!�$ׂ5��ʕ�"%�d�� �RG4!� W�D ��͹x�D5I���!򄇊?�\�p ͗�vV�C¯s�!�U)y�2�ʛ�P�։[�c�3!!�D��@�h�H�$r�!��"@9!�Ɇ�"��a��m�(����"�!��TSPa��T�{�5*�H#�!�d0~�&�r�HL��2�H��f�!�$K0�^(0�-̀D�r;F��l!�d٫�f�ɵ�O�hњ��"
�m�!��ǵW���h�&Ӷ���$4!�d�,��4�@�Мeʨ�˅�A�U1!�$͓g�)@g�ڴW!��1��ܯQ*!��_�`Edps@Gu	D�s4ǌ(\!�S rr��U�U8R|p*2	'�!��86g^Q1 ���-C&5Ze�W�S�!��B�BA�e.M�m96��"�(�!�D5-��a�ӤK�'���#�d�!��C��f@ۅi�@'6q�Rc״�!��ɍ@���I�X*��r`ʽs	!�`��ɱ�^3VZ"5	��A��!��h�a�d��PpX����9�!�d��z�rd�Q��18��9Fz�!��w���A�U(cվ��7�VQ'!�$Z�T����� v]�e�w�ėV"!�d�'tb~�9s�L%XVvy�J#s!�$�q�(J=g�q�6i֊ !�䝏hB�T5���\*ȺӮ�h�!�D� [Y�Xk �ȈcI�1�Et!�׏9~�`� ���0sCȇ|!�Ď�nxf�ZER17c�\`!Cǈrg!�d�"4$�q�G�ts�<�#��7L�!�dL�Br��+� ��>s����|W!�+�&yI&�&>�5z��]!�� X<z���Q����7+D9��"O��Q��|���3b��Z���"O� �W��EP���)JMܘ�g"O2��� �4}��h��=�Ѵ"O�� G��!�2�F7Ӳ8�"O��`�.�;$7h�&��aZ
8�"O���KUJ8�x1�:Ji�lh�"OX�@�3���hei���v�@w"O,H2��3u<��	�>�\4[�"O
�#`���n!3�N��L��)"O���)_�6O�"@m�"�š2"O,8����:`6��"�=V����v"Ob����S���Ă5��"�"O����+O���PG�ّrj����"O�� Ca�fs�A:�`ھq<��ۑ"O|lhto�G�}9`��2�^q��"O���G�G�~¶U�A���b|�h"O��٢�N,X�aA��,���"Ou�����}Z��"H^�"Ox�8�H��-*Ҙ��U�f�֍��"O��r#	�F/pr$g�
&����B"O�q�� $�h��&ҳ��Y3"O�y9�%�.��ĥ[�n��<��"O���G��k��S�e�0�T40�"O�񚂇Y&W}�0@�d&(|�#�"O6ti#A8U��Q׀C:uN�"O ��(DPC��B��ː\�L��`"O.����ľ|�"0�.�`w���"O�)��`��T�.DA��[�P� "O6eK��6 � ��X/s�\S�"O�͓D�  f%:��Ī�*�q�"O,p1C�E�;����
�87�f<K "O���� ��~�U�Go�R�4;�"O:]1� ��8t`c ��.�0D{�"Or��P�4ǌ�(S��wI���
�'��m����k��]q��Q�M�ژ���M�EH�,��-��*v"�"O\��֓p�f�T�ȶG�1�`"ObB�-؊��hc��$e�d���"O�M3���t�	�JJ�a��"O�$��d	1FD��@�!�Z�*�؀"O�,��+��&�fcޟ0����g 2D��PV]�_���X�N ��6e"/D�L����JĒ�ؼ U6���H-D�l�P������#��W��A�R*D���5L�p
T� .�3ATyڒ�:D�a�*��a�6��Wi��pA�<D�(�4E6Q�/N;#* i���9D�P����SJ�۴��]����'I2D�l!���+_�^���G�*M���Q�L0D��j�)�G����v��c�$��"D�4@�щQ��Q"5zl�I�H?D����^b���P:>�R��?D�T�6^�2���׍������Tb)D�d����2HaɊq�P�pڈ�G3D�����U���%�
�T.$\Ҷ�3D�`C��7�����-�$0D)���/D�8%琢'�
U[�J�X�R1�E D������v$e�WF�I�L��=D�0��T��kϠ���q� &D�p�S�u��8QA��X�-���%D�Pp,ј|�Z���A7|�љ��?D���ClK#&&Y�Tn�AQ��6g=D��ɦ�Pc"�	7F�E�v�`DL<D�� �Lae�'8F��׍��<r"O41���%�����^<�,3@"O������u�����!8��`"O`8X�a��r
��u@\ jM��v"O\�-)P6��@�J6g�B\�pb�(�y��I�����	\�Eqa�^��y��%:|Xa�(�ON������y�M�j�xpM�L�$�����y�	�NG,�j��'L�20�A��y�&T*Ƥ+��(BHI�����y҆V�>�q�&9�Z�S�.� �y2�D<l�d���߮5�����#��yr�Y�E�20���-pZ�E-M%�y��uǌa"�o����Ҩ�y�A8I����.��~�a����y�E��n�X�⁓/z%�,�b���y"���W�D�§סp:�)ģX4�y2�֏f=(uYp#g)36Iߏ�yBΆ!W�����Aů�@��e�M1�y"K�g3��Iv��RNh���F��yR
��;��`�s,ԏ5�I��U��yb; 
��o�.	�4�ƢH�y��]>Pp�UK�� �|��R�y/��j�.��1損I��)YW��-�y"B��Rt;�`>C�
	!7B >�y�FČ%�z�QGdDfΖ�G�["�y�G�*f�-2��	,5��""�PyR ۩@<�HY�A?$�P�G��R�<�FgD�dH���lȅ|�����h]G�<qG� /��� �!�,$�d	��F�<� I<�b�*�m��#Hj�z@M�@�<���DG.���*�@��Gb\w�<��J�.)�҄1���5�4��cMt�<q��õa�8��NWx�Y9�`�m�<1�/O"TgTib��w_M!��<�ңA+[�nͨ���::~H�1g�o�<q5Ď��DC���` JT*E��t�<���F�E�q��:��(B�K�r�<�g�]�w��ġ���$��	�	c�<)�H
�>n���r,R7��MI���b�<yCƙ�ҤhD�\��0'v�<�4&ȝb�(-�@�V�OFƜ��h�p�<�H/�~� �]�=�x�x���r�<a5�J�`�y�@Y�;�^}���k�<�d
4b���Csϊ�9�01xc��d�<Q�A�:WW ��Ǆ�S1
�k��D`�<�B
$��砄;
�k�G�<��l
Ԋ|��AM�H��X����}�<I���$TF��`�-W�ؐ��}�<������`h�x� ���bݺ<�!�$i�ٰ�c�E@|]H��P��!�$��Ps�P�R�A�}��a� �N�c�!�$M�`2N��c	����i�v!��AY!�$׻C�, �G��fA�&�6�!��8Vy�(�h�*�|���)0�!�F*C��Ϡ:�=
t#B�{�!�A�V���%�P��ʺp�!�$�>�0HfA
@{���P���P�!��'&�H�b�S�$��z�*@�P�!�́�2%ҡ*0��+0G�#!�V\�\M8�W>'�<�vl��>!�@#G�Z3�ݼJQ���a��F�!���$�>Ix�L�=[T}���k�!��4A��d�V�H�N��b�Þ�%�!�� z���J�v���z6ܨC�"O��sP�/W�9
���|1T4J�'�L��G#�1(�ʝ��J?,���'&T4h�%ZL^@8�J�:#�б�'7�%p�':�� Z��

�P�:�'�:�ۑE� �r��F"Е,��P�' �Y�"�9N�+��ӎ��
�'Ұ@IʌmVp�Ӂ�ߊ+xi��'*�@Ѧ];#�-�p���'n^�:R��)��Da0#��e�5��'$X�GH�4j��L���\��lr	�'������Jt����O6Y"����'��e��\ q�r"�DG�G�����'�0iq���^H���<`$��'6H�RcL�{T�5�V釭	l =;�'�l������/	�f��'�����V�g���vH��Q��'����aGJJ�f"3�@�oZf�"�'{� ���̩a�~�@�lz�<S�'-�@j�=i��)�� ����'
�	��+��/o�i�MDa&���'JB� q�^�N�Ęu)�6�u[�'�Č��L��J+@j�'�&���s
�'%��1U�U�K�V���R���"�'*X�!Q�UEґ�e���:����'�d�� �$W����T/G�'�6���'	z����ܸe��x���M)%β��
�'ư�C�MM�?�j�D��,n�4j�'�􈆏Hl2�H&ݘm��K�';�@ # �)����Ϙ�p��\��'d�0��44���B�V�w>NA	�'r��φ
�4IP��.K6�q�'��AP��-*2��c�b�~|Hx�'�8���j/�lb���~���I�'�fM�^%z
P�8lY�$�x��'�tb�n��X�
�+&��$�Z�'3��X��X���҃��t$t�X�'��@Go]�[(>Y�!�)p��e�
�'�B �bܝ�,P�Ąj����'��Y��|�0pJH�bY2���'l��PV��!a'�Pr��cI�|k�'�@x�a��>mf,�&��U�(�'��UPrᙴ)ؠx�t���O����'����5�W%�������5�����'����A$P�mkN����,��a�	�'�Xx9E,><(�ᵈшV6L���'6\�&�V������ٟG!)��'P������:O�J���9=�l��'J����P\hQ���ܩ葃�'�'���GޤC4.�E���A�'���K�l��?����C��F,!�'������cI|���-L<���'��[�b�Ep�=;�jV 0tE��'	İ+!�G35�pu��
z�ڝ��'*b�)���w� �hd �2 �Z���'����&�X�+8>�iRh��p��H`�'�&��˨<0,��D���ri��' �+%a��MJj�F�ȯȲX��'��(�e�;>s��­~�h��'�Ȱh��T4Z�hh*T*�dl�J�'����.J�4J.�b�`>L�\��'�R�h�ȟ� �`��CI�F��ţ�'Z�8�SN�:uÚa�bϽ.r:b�'�"�y��:/��	K㪞 �U���� 0�oրr�6y��
	g-����"O�A����B6~��cdWW����"OT���CM�Q��]2W�˯�.(qr"OR�k�4��93�*k�u8�"O:���#F����,߽i�N(B3"O��2t������ C���"O��1�UP����7�E1]�$١`"O�X���"�.�ѕN��Y��Q`�"Oxd6L��9�V �����X"O2%�sb��)���?�^�"O�%���U�xZ!B��pf�)�"O���1Q�����!��9Z�"O��
0F^�#�d�H�m_���i�b"OP	P�ֹt�U�ƭäo���"O�1��V�wP$"1��/K�i��"O��cw(����U�RO@�|�@"Od���
�&�=�qD��h1��Su"O�]�E���'N@��T$����"O��isD0��{�S+�	U"OA��	�6o-�ճ��ë=`��'"O�P`�ȹZ1ش��o�S(��@"O`H��&L�!rx���l�E�"OH�avc�3<|=FL� xh��"O�I�V��%�l="��	[�
7"O �PŢ�fZ�� >r^bD	"O��i����\z�`L�9G�ݢ�"O���gN
�(�ԍr��%bW�$
v"OZ��Ɓ���Z�����+T�t2�"O��Zŭ_ a���7&ϿgC4,j�"O�L�s�����ȡj
�)D�@�M���y0�.D�mU ���o'D���Do�)�>��"��8>D��q��(D���pʀ,f�\�"d����+�&D�("e��9��%듶}��U&?D���R�Od�\�C��,C�����2D�`R�g�a�()�C��)�j)� �1D��z�ǉ8(��1��
h�l`�v�0D��� -�TyJ�r�Lm-9rr+-D��0#�F %�>�!0FJ;�ج��!D���/�
B(��Ba�6w	��� D�X8"m��E^"�dH�7��0Y�<D��8�&	{'xT)U��;�d,*�&:D��J3���p>�9�V�G9_P8
��=D�<��F[*;��"$��.�v=X�:D����h;��t�^�jU����u&!�d_�u���8B$��"5�䪑���E�<ią�P���7B�s#hdZ��D�<�N��"����PgАR'lw�<9��T��y{���>#z(2O�o�<� ��v:�]��M06�&uAVH�T�<���_����%�^�60�1�Ri�<ģT<ߒ�xKpȧ��c�<�Kǽ=��(@fռ���`��\�<�����~]�̂���<�̳��^S�<I�e��^x�σ�Jl�)e,�v�<QCG�y�v�QW��S洀�u�<�����Fd2AJ7�O�5X:9�j�{�<Y�F�,F~)�cA>�T����A�<���m�0�Ӣ	�Gx�8��g�<�Q��'ct(�I'��#�.�Q��Pb�<!�Ň�Z����#+��!�pI����[�<y7`��,�Bq��?=�p��gfZ�<����'��Ö�����T�<iĆ�)8� ��*F�~i]c��P�<� ���2e������/�ap��w"O�hb�ޯmv���C舠
�:�Q�"O0[���A�P�6�ҙ=��̈�"O8�q �	F�V%"�� �ZAH�"O\���B�0߂��h��)�0��E"O,��%�U�V$���������"O����_�~Vh0�A��^ֈ��b"O����,�8%�N��b�qQ�"Ouбb�X;�}�` ��;�F�"O��
C��S�BTy��+k�:�[d"O��I�BWz�4�R� O�Z�ȅ"OZ����J�/5��LW/�(�@`"O ���Ĕ�p,���d�%0�re�F"O(�+�Ƀ�:,�0YwDK�P||�"R"OnTc����$5Ԅ�P⛮�Tѡ`"O��`J�f6�SS"ȊXy�h�C"O��PcB¨%�v�  �,3;V�R"Ox�!�� 4Q0)�w�E0��ۆ"Of$�tD� 14�3e/�2�H4�u"O. B�fS���e�V.b�8��$)Cs�<)G��oQ��R��i�0Y�M�p�<��l�]��!�ۅmx�aE�<q���z��Z�e��M0�!�Z�<���F�f[ �����?	�]�@@�<Y�� �&�����
AEe@H�"��g�<���1GUl�@W��Ԭ0�Q�_�<�Fߗ��Af��[[�Qڃ�\v�<� �S$:|�b����_!���6�Tw�<���(�(�R��r�V�:��~�<�w�L�xH@Г�!��QF8�dp�<�+�-�Ny�q��x�Q!Lc�<Y5��2�1��ل+�29�aFg�<QT�R"n� ��Ģ�B���Se�<��_�¨�4f��M�'�	��a�ȓC)p�۳�v��Pk�g��ȓN6rT�Ri�t0(�'�e]Ն�g\�YcꁽN۪a�2���۬T�ȓ}�0��@�L����7/P�OY�t�ȓ�p����7�����΢^��)��V"�����7T�JÉ@�^�D��H]\�i���~Mr ��
ʋzl"͇�������_`�\:Ԃ]E�������A��
$ ����� 4�襇ȓ��ac�-�0`l�tj\�H����yn�E���[�V�2D�1Cl1D��ҕ�!�B�9Ƣ�"���u,0D�|
���0����P4 v�.D�@+�n� $ |bҤ!L�gN
��ȓg�^�愿m����MT;Y�-�ȓ����cR�3�
}Q򩋹j �a�ȓk�����lT�ƹ)���t���ȓk�Hh���.s���a�!�4���&YH&*���@�W�1=�h�ʓ9C�=�5��
�L���¹e*hC�ɔ=h�|[w���-b�H����dC�	��(���NzHhd��k˲>��C�I�8�e��i�*,b�@{�'G�K��C�	�.��A"@ʹ4hu���ITRB��x���64��L#T��[�B�I7,�*��E��i��i�Ҭ6NB�		k4i�D�W$VF����4QB�ɸ< �a�ظ8�.�2n˂+�����O� ��Sā�I�6��J� ��I�ȓ6�\}�3:q�<�'Ǎ9$EJ��S�? ܙ���ϻ;80#�A%��"O8`��L2&�P��¡P�p&���S"O� cv�ZV�rDa@+ !����"O��匎���i� I8Nx�)�"O��bD�^V��9Fo˛.I��2"Of�{�B�IM:���G��.)\��"ORY'��4p�Z�A�L�0��"O ةW��$���Yw陙O
��"O�mg�J�U�,�z�a�VԜҁ"O�`ḿu���� �%^�=
�"OD8�Z�8<��� ���ق"O=�����i�hp" 4q�>�G"O6�ٶ�U��l�i��]ܬ8��"O���K����VO��$mE�6"O"<C, �\P|�!$N��?��l
�"OL�*$���`$�`
�����"Od���K�����ͱbD"O�̩���x��P�e�ܑK#"O��yRf�+�`�R�i�RKx �R"Ov}�'�ՙ)ʖpY�(O�A����"O,�P�m2"zt!�ݴXe"O�h�_5c�œF@�8+��Su"O0I���z	�4�5 ���ȝqR"O�M��
Ƨ7_�p���$Ǝ�)6"O�,;�� ��()���b�(��F"OITk��s8��;A�۱�`��"O*�J��I }ʈ6���4��"O��Z1�>j���e�>��́�"O�mQ�@ˋ.�4����(�
ع�"O� ��i	�.��0ա��0�~e{�"O&�*ccޥSƩ���=p�F��"O�iQ@JO�$4��%��0�fE�A"O$���
l��Ȩ���>-*@C�"O��G�P�2�*�q�(�	0��3"O�ybnɇ+�������F���"OV�«<����V�O�lp�"O2�����
�\�:G	G�ZAX�QE"O<%rD(M�K�hD�����=�r y�"O����c�:Y����>V���[s"O&1���K�U�t�ښotԄ{�"Oab�&F�}�p��b	yL�Z�"O��&���u$ʨ"�F����W"O ``�瑴z6t93..�@�"O�4��N hܤ��+�"Wx��A"O��ɋ%��H�
P3]w����"Oz�H$�@-!��(���9�2 �2"OȬ��G��H�P%Xi	a�`�`�"Od͓�����e�ff��"O��y�`E>9�X���J��t ��'"O��j���lW ў_|�	B"O`�qcJA�bd �%��*GF�""O�����	�p�,�pgbĦ7D}�Q"O�M��:S�<�rF��1#$-�"O�Rb�ف/�Ƞ&��z���"O�����&��9×��QX[�"Olp�A�^�3TM��!�3\m44�g"O�u'@�؄����Vexq�"O�����#]y>�� mR��v"O�L`�)��2.�Q� �&>��`�T"O�p�p �\�ֹ0Rψ8=
x�83"OF�ú}��qJ���X��"a"OI�����h���Q+�Qa�\��"O�4Y�T�)�\`�4L]�$􆸂�"O���¬�E���%nҲsP� x�"O� �|CE/M`66���тG�Z0B "O�8�'�V(�ābBʖ�T'ȑ�W"O��Ʃºm%��Ɇ�*��qv"O��%F��p9�E`�C(<�xI�"O|	�R�
��)��#N��KW"O&U*�P7ά��BD ���PT"Om��۫sNB��r~ds"OT`c���P�|8'	і-�R2"O���C�	2�p6g��B��á"O��C�	�	P5%�	�ΐ��"O�)�` �[�>u{�΍> >�I�"Or(��m��T�(�C�$*�9Y�"O���W�Қ&
�%���߄�ih�"O��p �Σ`Z�Eq+Ė:6��c"Od�Ï�0^�f��ꐍ$g���1*O"*T�72(����e��$̦���'.�S��� *����'y��6�H�o)0��唥���:�'���z�GI�E�U�(BA�U{	�'#n�c���6a&��!Wh��h�t0k�'�Ĺ!�K�;d���V�_ti�q�'��`{vgьJεڅ(�:hdΩ�	�'I��`0<&�FA��3�Zh8	�' ��`D<U5�Z(Xz�]P�'T�A0K�3(�CeO�N�~�
�'�Da �o@�Ұx��O��F���'�<���#��Q��;T�.h^����'#T�q�j	����#��UT��'3
A%�Z�$�@%q���a��\s�'cT�[���`�*��,!�'��k�B�9 �%�tLM����
�'��b���fK�$��oղ|OHA
�'��aB�'3\����g#	�4P�	�'S�A�g��cD= Uȧ	Tu��'b4ɪ�@�dXH\��@ؓ��;�'n�A[���1`�M���l)[7A�T�<��i #
붙[#]��%Q��e�<�U� >�	:�%K"UuN�Ӵ�^v�<�S�{d:�ؑK�7Aԝ��o�<�%T�&~YY�	"�t�'%b�<iPc�yN^�X�j�'me�V�HH�<)��ϤQ�p�5�L�St���V�O�<��E��FM��� ~�;ծ�O�<�e�"m9���Ō�		G���Tl�L�<ٴ�G:,ލ+�۰X>ڑ)h�D�<I�GX�sUO�-b�~���'�X�<	ëڿZՎ��^�҄�Ǌ:8dh��^=����A��:��
�Ą�2��VE�L-8]¡C�M^f\��@-t����j;�J5��QZ����޹3�D�	��E�s�L<@ҠT��&+�� Z8nf�H��,�0���*U"��K�-�2Ԃ�ߍ<��݄ȓ)�Ը����`)�1 �K�.�R<�ȓ9|XKU��3S��ă�ΌJ�|	���%k�-�tӎ+��$�.���c^��%�$� �=x�8�ȓ3Kd!P��ϔ�F����q<$���+E6�gN^ 6����F��5-�Y��(X椱 h��]HMrf �2���'�|Ѳ�bW	E�@rP�ɒ&���ȓ/Ҏ�7n�s�@�t��{`}��+~���4{�-ѴN�C#��ȓ�&Lz�A�'H]��8��
V�0ą�S�? Z�B�T����U _���"O� � %�� �?�L��!"O6�rE�F�����ڐ��q"O�h�U��
ug�KЮ±~�e;T"O^�S�M��Yۆ� d��!�"OL�����I*�I�kX�d2*���"O��#�G�"M�C$�H�@��$"O�,ڂ#I+,qve���)��8JW"O�5����m���(�<��@b"O>����,�T5��KF2�V��4"O�h#�,޺2����ŭP���$$Wt�<��j��O��8Qa֬4j�h�5�d�<i��!8���(�LϟE�V3!��_�<��V"%(�����ц$MV�J���X�<� (�PX���wv���\�<q��ǜ4���2�ށBB��2D��\�<Q���r����5i%?��L�6 SV�<3!�1
D5�¨�y �5R�+�T�<��@ǈ-<VA !�2�V jD&�V�<y��# ��8��`}�}���P�<yg�ˍX��B@ł� �%!��J�<��a' ����+F�zL$a⁜D�<�#�.0@K�І'GF���W}�<�䪊
��+�gl�%cBh�R�<�cڰ
괒efR�T���JrH�i�<�JG�Lu���J/K��*F��c�<1�gʡ-�:%�ԁ��^��bHa�<�r+׶����o��������]�<�M	>��HH��ς&5,l��KX�<qb�E!��@ǉ;o�D��`�X�<)S��b����BQ k�$�0e�n�<�v��
	ΐ�%�٧<�()u#Ei�<Yc��5�~���IA;!4��d�P�<��ϊ�M;L�P��,�r��M�<��F�;Ģ�6��<1��A�<2��))�Es�	N�]�����Rt�<���L�g��̓�.���ᰤ��E�<� ����mh�OV#n�JDң�A�<1t�D�&�.��5�Q�J��U��E�<饎/<`�b�X�&����"��H�<QpN�u�� �}Ql5ZE@M�<���.�%K��We����^�<�� ��%E¥FڌM�`-;���X�<�0L�0�>t)���j�L�*u+�J�<	@MĐg݊�hEm�5=˄!���H�<�p�K'M�$yS�	��@Q��n\o�<��ា�
\�҂�23Ƭs�(Ol�<����	w^Qpe΅�o�$�A�Aj�<���E�:7Z/�]Aa�Qj�6C��,l ց ���q�by�)��]$�B䉩!�ؗ��$FJ����>��B�}���"�<O�8I��K�d��B�*%{�!���XL�a�ߖ6-�B�I:�b�ɢƋ�~�>E1 ŝ4&�C�	�{�-k�䉋e��pxr���x��C��a�p@x ϒR���:.�!N�LC�I+{<�j��91������m6C䉁]g@e1��A�	��c��+<�B�
x�<*���Rx0*�B\؜C��5a��5�d��-
si�6D%0B�	)� Q�fΝ�Y�!��3*"B�	��x�� H�1v��a/�9UC<C�ɴI�ȳ�ʛ9by<(�����B�	�; LEo֟R�@�e�M�C�)� بK&���!�>�%
ɷA�L)��"O�²n�R�P�SP�^�����"O��sS&A-LR�аF��-�"嘆"O8�ɤ�&q��$��Z��� �'�4����8��5��ḪS���!�'6��cÄ�� �ۦNԺ{��e�
�'˾��-���1#*
�{.��+�'�ʹ�aF0f�4�8�aϣ=Z]h
�'��Ui���"�lp!2���7J���'k�Y���)G��R���*�9��']f�1d#�82�ĵkыZN��ܢ�'8A���Ըt!R� ��F�BH��'�	��EN��ZtxQh�&7����'[~yز�W�ty���+*J�{�'V�H�aY#-�lc�e�L�*�H�'1µS&�)���y������B
�'��"�l�T�f�	�犀6~D�	�'�i�F@Iri��U�fż\�'��s�m(V5�H
5��b����'�n��Ԧ9J�����n����'�� ���]*;�T]�ԬK�`W���'Þ�����l��
��C�Z����'�^�j�7db`�]�@���i�'	����H�g�a�N�66��Q��'W��u���� 䕫4��
�'�(� 4��00Zܰf��u�6���'�^��1c��+fڀ�eEN k��!�'��9���ٛ�~	s�*��mD��y
�'����T��N�(��k5e�:(@
�'U�!$�V���s�Ēb�LZ�'/|X�(�3�@��O��(}��'i�x0k^i{���%eT�=��y��'АX`5��J�f�p�DA3; *X�'��ѹp�,|RQs4l�6i¥i�'�zP��c@ �Ӷ4��ȹ�'%�Q��:SP�����E2/SpH��'�f�hƍC5 n��d�
1sф$J�'�Z��ҷT��r��T>�)��'Aȴ��f�,����_��tA�'�@����0� S�N�eS�'���(C.�0_b���a3�@!�'�b�i6��9 �w�I�,�'�^y��`�S�lՈ��Z!y�V%*�'ELdi�䝥�l}еA��K��	�'�������!D��� ���(�
�'�����O�U���q,�R�'�r|�t�ɂ����: �HI�̓��y�A��@��N43����_*�p<I�%_bT�;���^φI�1!R�"Җ	�ȓIt4H���'#�X��b
*%1vT'���"�io�Oq��D{��=,�@�.�1t���;�"O�����~X*`�W?b�8]S��'ɰ<�C�۽pߦ���58q�iYփIR�<!G��)e�\j��/&`!")�<���5�>|���D:j6�����"�a���Ը�e��pT&�2���=����6>����恇G��(����B<�ĆȓlÄ��'bڥ[��!X���I~��'��c	�h�<%���!�d�A"�ff�G{���]?��`�pf|����1 ���]�<�dEӱu����H�-���O_�'�������T#,m���K@� 0�%F�- V�O��=��:�jG.LL-YìZ�_3�C�)\�\�ȓU���hGc�&S��e3��2��l�x������ ~�a�J�	1cp��� ��524�4"O�A!D+˨!8AOӼ���J/D�4A�8 �l	u�+ ��y�!,/D�Y��==��0y���9zδ���I+��OZ�b?y� őf�浀��J��Dpr�*6D�˧���J<cb�o� �� D�4�W��F�4%:D.�����q�>D��b�H	�R�>%�.���Ԝ4@>� l.^q���uFE� ��!�ʡ2���$�
��'ל�W���.@T`��*X�x<!����?�h�H��f��8i-h�c�@�214�P"O 5��[`�Q	2���bVйB��T�'�ɧ�9Ԡ;hxuS�H{%��aP"O�5�� �;9;F�c�#�$���"O6���J�x�*��,֘1Bv}QE"OV��դѪV�<<��_�%2� �?O\�	c��hO��Z���}��t��W�r��'"O`��G�J�)��� �˷���Xd�x��4���'6F#0읰%6��qU-Z����'�V�pQ�^;wB�-q��#dy�<���<>�Dj�e�_pR�1'��x�<��蕦ŀ�z� O� ���!�Y�<yuh�!�X�
�BI�"����$�Q?I���O�V�Hz�	�s8Z��T��- �1��
L�B�I�:�.$ 5�M+%���R���DC(�<D{J?-��C4X ̭am)_�b�3�E"�O���=J�̩k��X��c�ӏ8mb����	�6�$��O��&�3C�"���g���=ѣ��
[�~$ps�ԠSǸ�"R�E�<i� ͦ�L���	 (*��¦�M@�'-ў�'=d�eM	��޼��'ӹG�Z��ȓ^�RY� �[�Ծ<��*�`�Gxb�'�����U�@6ؼ�d��WN|hz�'t�r��÷<VlXE��=h(HN�4̓�ا�O馨��	�?Cg�9�ĎI�"�@ד��'sNU���i���؈��M��yb�'rJP��J�g����@� n0���'�&��+�Phv��/#f��ά��<��&[$��g��+),0�r"� /J`!�DNS��"�]�B�����,�"O�bB^�p��!#��Y�ܜ�4"O�\z.6 �ZQC��)R"O�Y'N�T5�a3��4�`�y�"O�`�Dǰ7��U9�P:[�6���"O΄�T�(a~4�JP�f�dmx$"O�Y1קH8x�<�aפ.��`��	e�OZ���gǚj:r�)��
)mS�5r�'�\`K[���,����$aB�P�'v��bq�h���bMZ�t�	�'��yR�_���SЯ�&]X��'x�m��J��p�[��Z+�-�'�h�"qH�>+�,�W�-")�h��"O��� ��	GvH��$Q�<�"�ipў"~n.�='D��D߄n^d!iC���y�)�'
߬�b��s�^�򀦕/|]��1'(UH�K@A�.��%�սO<�'�Ć��������Ɂ4r�	w�*/q�}���)D�8	�J� 2UPPB�f��8ӫ$\O^c�\j5΄93qꘛ�KˢE��aQ.D�0r�#̾/>0�2S�ǵ	*��9��>��?Y��i(k�24���./�a�4�"-��l-�S�O�:0{�FB���Ŋ'�Z*�`��	��0<1�\6>$t���$f04]�S��|~�!�Op\�
E����AE�UK�u������>٫O� �b��<>�, ����=5���a"O�q����H�5O[4c߂0I�"O�(o�]$�Up᭔�4zh5��"O$���Fս�,�㔊�Nc^�I$"O ��<Vs���oQg���:�Q�<E{�� �T,*D�K�8o�������'Ka|b�ށ8�Dq�1$C�+}z��#%^$��vX����O�G<�e��6�p"0���&�a��:9	+1
ˬ%��d����O"=�.G2rK���VeD�liX�q$��<��Di>ɘ����� e;rܐ�j��>��I`��N8����O&�"|J�����bi ���a��+�WX��hO�OjTP{�*�CO�1����}��$Y�'�Zx��G�1ap�ñ��_��+�'&��3�e\u��1�R�F��!��'�$���Yp����vMªP ,���'�d��K�[t9���N�H@���Q��+&��sj>��0���0i2��#$��q`׶Xkn��&��Q|Za�'���yRGT=U9�@�㥟������
)�'�b�i�D�H��4����7��Y$��AT� ��;��	`��!݈!�l�#�V�dj�R%���?9�'���J�\�/�l��`OP�L�J&�'�Q�$�D����f0��:F�E�>�c�Id�'�(�j5 W$� #YY��N<y�4�O�yR.@�8	:�R&��N���D)�S�ON�)����/{ƼYb��12��r���+5��?��ɑ�@���H��]d�F��6i5�dt�z�C֧%�L ��	7̰9�t-�:�0?�&\� ���-\W�H�rlK�}���1D�<җ��w|�Db�$�)>�ֹ��1}��'���
ު!	�ݢa�*9l��k�eM��ɭ]��B&�8W�)�Vk
5o۶B�I����5L<N��,;5G	%,4d�>��i�[Gmv�&\TD]ˣ`.7�!�O�IܡS�l�7C���B��Ι��{2�'�dI{Z��ٵg���B��Gr!����D�R�B�k��
��%JYqO��D>�)�I:A�D�9p�8�H�a��7�a|"�|�԰~Ϧ�8��VYp첁#�,@�=E���1��I�@��:E������
>�L��ȓ>�ʍ1dO��p�򌇰2����}�8�!�@!7�v���Ō(6����p��<ځ�?E|R�+��U�>1z�ȓ�B	�����Ƒ+Q�C$j��=��g��])����K�h�"�ʙ�0��dV���`� ������k��Ą�~�(�K��&eM����אr~��j>��2�#;l�r"�
g���ȓeKH��$9����D!�B1��ȓ<��t�B�<F�,����O�c�F��0��S��,p}9p �;[�H�ȓ���Xd[2B�0AU��.���
*��Z��*r QݼD�ń�9 �}�"�ׯ�X�Pw-��q%V�����Y'/�'���kT�ӭ�d����U���B�,�ƕ�-Ѓ+Xt���o��@�Q��+�:r0aZ��Jy��
�
�����d:��!g�ߣ9+B4�ȓE�(��g�v�r��D�a�0�ȓ/�Ɛ��헒(0hd���K!f�ԅ�h����ӑr�u{�j�Z�2P��-d���׫Ԭ|Z�bv�]����{)��/I�<��R�5���S�? J�+1X�[.���	ƨ!�B�3""O��!�ƀ����������w"O�m*�+��u۶1��(� W{��5"Ox̹�j�p7F�s*D5���"O,���1I���{�I2^�z@�"Od �k�<��K#��op� R�"OdA��E�5Pβ�xQj�	xd0q"Oډ�b�3	�C�H�8�J`"O"�t����:�5��(:��x�"O�i�e�4j�5��A@�Ix<H��"O�`���;9�r�)1�ւ:���W"OT��bR�qQ��fh�u��]z�"O��k�$-:�
�GQ�㣉1�yBIH�#��0wI��pl�9
ER��y��E5u�Rћ�,p�x�cF��#�y��8V�m���ūUu��CC��y���'@N���܋%_���v�,�y�_�_�x� f��s |��F��!�y���a x���#ܦĉ� ǣ�yRɐ�/� �ؤ �R�T@�]��ybB7m��A4숕aO2��ǟ��yr#0 �JA�r��/�q�Ӡ�	�yR⋋������;@�X��#��y��,4�����$t��yR'�9+�}��W��X�`�� �yBN��
�*�����3�!2q*5�y�2*�0б�HD�Zm*���yr,�y������9k�~�3��0�yaHpL���a�1�ƙ�y�,�:N ��`�H�>�;dA�>�y��@@g���#��F;*Q#%C��y�.�=v�6	)ii�A!B�y�E�CJ�2�JK.K�:$�Aȑ��y���2e��0d(�Nn>HSd��?�yB�^���LXr���t�� ���y��L�1�\�kS��]�J��V&%�y
�ٌ0��g�[����t���y2�ߖ%<�5��cU<@��E��y�eI�f��]"�[�W_V�`��y� n����ïZ�,<
$c� �y�%�M�0Q3�+U8��sɆ
�y2E@;j�RR��{&xDF���yr�Čx�6�_�j����J/�y�������1b��+h��@JG9�yÒ4FvDP��"��P"�,��y�%а=V�|���݅�IIQ-�yr��Gl��(f��2��;�e��y�F��%��%ݤKTd�1g�ybM�yPe �7Vs^��`JhBў"~Γ"~0��_M���d�º|�ޥ�ȓ*7��'��E�*1�/ôU�~e���?Q$N��:�N��g�đC��Q�W�LT�<!�L�-�)�+��Ų�US�<����J�b��/�f26� P�<�oVc�TYA� @����c�e}2�'���I��L@�*DP�	ODx�0P	�'?�icc�w�����7�na	�'��%�v-κ�'˜)�����hOȈG����B,>�b�ǟ�_��e�2��=I�yr�N�0�
hR��02�㑨�3�yB��* ���S��C�����D�y��� *�"�a[
U ĹsB�E���'4�{R��"[N����J��r�R�xb�'T���#��)sXTȔ
�,I7�ߓT�<O� p���HB��\:�Ʌ2�2�3����GL�}B���,��4����,�y��a(<Q�4? �UH�5Ȣ�q�X I�YoZ~�����Fc^�^�H�t%�c/58����yRAl����9U|�����yrޯ$nB�$��3G�h,2pI����$"�O�dՎNr� `����|��"O��XG��t~����L�t��3>O��=E��]]�8d�Bξ�Y�A[��Py���y��A��2�X��	�<���y2�x2퉕_��)ё��*v�4��c��b4x�'��xB��H��+3Wp̜����*?a���T�2�X���\�P�h���]Z$<��Y4
C�?���SDBα�t(�)�B�	�E���"G��2&�]\fB�I���R`��b�,A�1�$7$XB�Ɉ({�]�r�!��b�"%D"<yϓL@u��-��`I�h!V�����ȓ)Ʀ4�BfWSi�ՈYa�t��ȓP��U����,d�NI�B�8,�@���U��@#)˼���s�V�^tA��i�A˕L��`��e�BE� ���ȓL���Ibj\&���KN�cZ�G|��ӽ �������j��R�td�ȓx���w��/$�����OԺ|?:����t�'��;���,ԮY����3�'�HI�`�3>�}b1ʇ����'���ꁂ��>��
��(���'�"Dȥhfi�uZ�(P����B	�'I�����&c�\�"���'��MX��y C(y9� ��Lwn�2�� ��=E��H:R�ʣc�o�, S�/Z�$"NyD}2 p�O�+��.CJp�R拋 $��1�'?�A��g����ᦄj�( ����'^ɧ�O� �`�:��)�̓^�Z�ӓ��'i4�{�.�șK ���X�>����0O�)�#
X<�'oB @�pբ��'=�	̟ *���jT��O�M�����1D�0 Ӥ/��0��A��Z�l�k��/,O��<���;(ڼ� \A�us�oQ�E<�B䉥6��m���8901��͂�O�9����O�L�'�� ��e�?��C���z��1	�'��b�
T�q3�q��铐1>��*�bC.�hO�S�)D���w�Ϳ(U*�s3�f�C䉥3���{�ppsoF�xp]
Q�)��<	u�B/m�Q�6Λ�R�`"O�]�<��'bD���K\�\"�q��/�@yb�(�O����m΂G.9��V.2h�p�'ɄO��.S��N��b��ESƥ��"O&t��P���zfC�:FDe��gBW�' �^w3Q>�����t����D����BYp!�D�;���0U�]6'�Zљdǋ�#k���4�)��<i��}����'��t�8;T"L|�<�aB $�v�X��!�z�b�N�}�<�OE,J ��Q#�n_\B,���hO�O�~-��"Q�U�e��ԹLqP��'��.7pj�i0EҶZ5�!��'t*xɐ�^�88��!�*��D��'��P��j�5S����N'L6�)O<q	�h��a�&F^��"D#&lتHA|�Ey��'�=Sf�	�mql�����K��Ly�'���'[��i� G�yM"��A���D<�����?��
����b�T^��"�.;I`B�4G3Of"=�2�
�$�7
8SZ� k�O�e�'�?�  tX7�\Q�XA��V�n�*���>	����T�H��;b&G�����z!�۲jY����0u���0��$!�$�!Z�� �֓@o����J�.a!�$�4(�,��7-ϋ�B�Z�h�8}]!�;O`��@�m���C�IOm��F�t�ˎ6��0K$B��<2�ݸt�Y���)��$q�ME��ڄ��A�/E�� �l��D{��I>�h�؄FN���y��&P�Q1�m�Z؟��uʃ�J�x�ra�=<���`� #lO���~��/�tźv���H�:�`u��yR�{1�5�2GՅ�IU^��}��)��!�đc@�9YX �� R�!��Y�����H:7���W�\�+m�)�a����J��_[�0�����Q�	ۓ��'�|��&	�a7����߭=�I��}r�)��"\h��{B��	/�T��ϳI!�DܹD���Rs�R�k�F,��P�l�1O,Ra����p<E��:q���CL�f�u����Q؟l:r�~Ӷe�����\qJk��aFh*!�d%n	����E�`�j��5�p��C��i�dt���L�AXes'�h�\\�2o�4��'1O��|���qKHt�Ң�	Gb�hq�Fx�f���O��I�)��;��<cwa\/�8x(N<ٍ�����t�6��!��g�>ѲG	X�!���*tꅆ��U;U�F�K!�D߅j�E �b�)W+|Yy兙`��yrgU#Wv1Oh ZKO�zQDES3��;6'�w"O��Q�� A��qʤ�Ųc&�X�%"O�l!���4:��R�	~ZH�"O�0���BJ���x�'ؘ�@���"O8������X�W��\�P<�'"O�H���ߗ,UR!��/^�]àٰE
O�7�*���aSa;1�\=�� T�]�!�$C4[�K?)g��Ǭ�9Rt݋�'�P�)$kۥ1�T������7�8��'����b 7<L�|!�Ν$�(��	�'��8a���
���X�&_�H�\-�
�'�Dc�Y�����.R�C�R��'�m+�F�e(\�i��E&d�dm�������]���0G�F�8ਤ�q�@Xj!�$�>H��	&�U�2�z�$O�fbqO����Y�a�`��AL��1�>�[s$���Py2��%S�8�G.^w��q��e�&�O���d޼M�LC��3AX�r#b��2!�ދU�.�fD�xd�����Kf��D�;���k3D �tC����&�S�O�z��Z<@V���7�0����'VJ@jg�K�j=��Q`��4 �����'�4���&E�0ZPLN�.|��'�%�WHC�-�Aa7Ȓ����
�'�.-S!O��F����.8���'�l�#秜#X�=�BD�?搙�'`de��!WZ1nPcBg����	�'���ɒnF�wtջ�N��Nކź�'4�d+gn@gņ(��.L�b��'�1�%A�
���Q�,#"��'�$������ R�-]�ep�'�"��t��+N�ҕ��D�7U��x�
�'��!�G.�.�)�+�� �
�'q���@���b Ѵ��(a[���'ˎ%���!-Jf�Y��U�P���'&,�����2��Ш]z�N��	�'�$�VΩ|"��� #ֈ:�"Y�
��� ��r�@�P�pAeO�+[r�Z�"O^�G�P�0��k��u\9B"O��4iܭ�6�	�bn�!w"OK'&��X���/7V�y�H)�y��P ����<;\@����y���&!X ��G
G��A����#�y��\�q��Z���Bs��`��D�y���3L��<
�"�)@��up�����yr��vJ�)7.��'!`qZO�)�yr�I*?jT���[�!�!��y�L�bMJY��"�"�AE��yR���buI )X�E���a��yb���g��L�cjT��p�߉�y���2�*hy6��-��O҉�ybg�$j^������r`[fF9�yB#*4fp�r �{�`�م�э�yb�Y�4��uh}��Q6^o`�#�'���f�ͼ?"�2c�P&ܕ��'J�}���̺o#"�0��Z*N���9�'��T���P�yQ��?��MZ�'U��ٶjɑT"93�M͇;9��j���

�ܐ:�%�d�R"͹�y�L.1��賔ĉ���Ј$.�yœA��Y@�+^>v�����y2&N�kWPI�HPa���F�ɵ�yb�7N�������W|�ȓe���yB�<E�T��&m�EC���ғ�yB�&:聫 DI�@�6,x�C��y� 'U:,�Ӎ�j�v�P%� �y�JCC�
�R�D Y�z=���P#�yb��2i�2�0��!P�j
$*��y��A<EO
��F�=R2ąR�
.�yr� <VlL�2,�@ p��H� �ym�)���n�v�Lhy�ƌ%�y"�6�,UsR �mL-�����y���?��H@���!�8|)��3�y�jS��t�Pd�n��1h֧�y2b�!�.Y��Ζc��̙��_��y�(�9l�U�eNSHN\�Gť�y2��.��a�-C�,{Cn�#�y�BВ�Z�9 F�#Z�|-b����y�FQ[��hS���VZTIY�A	�y�珱h�2�Ⳅǂ@��-DGS��y���8P`�����)A)�����ʋ�yRnׄ}�2��a�߳;���B#M��y�)��r��(Q�I �^t!Ra �y2ɸ>i0���vht��FX�y"�μO�$�u ҷzV�P��@��y�i�/㤨cN��9�̰QJT5�y�`L�{�q:Gę���ڑ��<�y"�x� T@3��<``$�p����yrÃ�L�\��jOY@� ����y¨�
V�(U��k�#]��Pb�I�5�yr��!Z\@`QcʏU>�J���y�O��$�ҽY��A2O�2�nZ��y��Z	+����q�ФE�̜8t�ߙ�yBA�t��`(T��W���CL�$�yN�J���f�F]21y�-K�yE!�@�W���I:�-y���y��ހ�z(��d\Nΰ�ɩ6x�x1�2N�}b�_��,h$��C���g���<aoAA���G�>i��_����N�sD�,
g�|�<�*ĸ8i�o�+Rk���$��"B�'��(iө؏8B�<H��ӡ(0��\!�&@�D���#u"O� ��v�ճQvБCQ�KT��s���o�T--O�=a�GNS�g�	�sY�0��'"[�dZc�6_��B�ɖ2��׃RvPihW��95D�U��w10�0G�F8���S
�)<���RC�"i��4�2,O��!'%G�C�4s(��\ٓ�V���l�j�0`XѲ��<D���'�޵����v��ySFh���>�
����Ћ?=�@�~�I�+ ƞ��i	�4�ty��-L�<i� �,1'�ͺwO�ieM��3�DA8�@�<Y�f�7x����'�ʵ2$��6J���6�>s!�i�'��J�Y&;F�i֧��ʤz��G��Y£�g|�|"n�:"�I���ӎe��R i���<���g��r I�>Q�Ír,)���@�uJ�K��]~�<Q6B\/=
Ax�#F�2E�v�@̓F�6M�VBU�����@X%'�J����٣w�h<rЖ������O�� �U���X���R-$�����K}�c@52<9��ݎ\�$	sHA��y�O�bA�	��e�Qn9[a�׈O�mG�$%�5�p\"���y�Z�!!؍�yr)��P�@t S���XӼ����y�OG����(���M�M�t�z��+
Qr0�Q"O�@򰫆�[�2!a�IlT��d��hR��'�`�CH#
%��@%�%%Oҹc�&���I#F�v������ؓ�4ZC�(um ��3��e� ��aĻ ~#>1��-�'a(yS�#Ԛ:�z���
�Vft܅�.V�P ��$=���B����I��˓�RӃ�+�'
(� P� XA@4����9Jh��
�'��ܩe�ʹZ
��#�J�� K�
��Xd�L��`�p}rFX{���E�!��9',\�of�T�����bՑ�qUL9`��ɓ���S2VLZJ���/#�\�bH-�� s�d�!7�6t�"�'��Y����C/�,YC�T"&z��'��R!��k����6x���Ř&c��D��"����Ȃ1P��a�떡.��s����y-Cy�~\��lכ8=@�ɺ�?�ǈG%z�r����͆��r��Y�	���D}>�[�(�9&���t�ܲ�a���W��T�2�J�B��)yD]&N��bF� Z�j�¡B�yʔ��g���V�&��,���(O L1���/L��]у�B.%�d����+A�͛Ei�<)x�$V�5q�)O�z3ĩ���d�ؠS⭄� e���Ý�ic4dP�k�y����!�겨��1\~t͓	���z�A�--�>�Ii��S��j]	t�Y,=�IQ�mPR�J2�"yʥ�Z� !��ڰ!900R�F�(��)�#�ՖY'�C��e^l����!=�Xe�BZ0���'�����K�|�a�Y>md:�����>�d����2�0?ɦ�*>��I3���5�<Q��� mh�;!���BЖiI���tH��>� Us��(O�ڵ��Z�Ѝr�cA���R��x��G�7�5�DY�B��`�'K]�P�������(!n����
��I�����l�eD�_V�U��ɒ���#�Bƾ��!AF�UF̈ 	Ȝ�R.l�s���d�^ix���R�S��~r4������B�-ȉ"�t���'?�A���9＼S!��j���'�!J�ܺ�N˺�΍�F,O.q�J���O�)�ЍWyh�슂��)+��q��I�o���kS��7DIQud�k"�a ?v��tnX�Dl�Q�O?�#@����h�z����duB�SDF޹
���1�O�,�S��#1��IE��	#�TQ�����#0�D�T
 ���}6�ɣ!�`�'�������@����f�M��]y��:;NR@ ��1]k����o����<�G�J�������	�X�s�CE�q��\hr,G��0)&C������]�jV1�Slƴ�e�M���S�	1�c1�˓y;��{6�,�i>�ctMG��`����[#4�nP��*�y�������4\�U;$�	�JT��'Xli�ް������
C���g��!��i<�)�b��L���9f�����$��L\ΓX�҅S��X>E)����a��@���)�$�>p3V�̒o|(eC5�G�M��I'��L��'Kny+FIK�GB��j�#7|Ґu[s��f��tb$d.D:2Y�_/�����X41Hj7��x;v�qGߛc�)��ID6pa~2B�0�탡aܱ}	�4��,"�d�V�#x�!�W�ɡ>���1�'����ѫ�z�XҪ�z$L�a���?u7t���MMB9K�o�(0�@��Xz��#K�-(	����!�$�{��2
=?�JD���[ )��𻣁@�B�ƈ��C�y��}� Ny�W �'[�s��� ��e"O&`��ÓǢ����ߡ(<1�*C�,�0(P,
�
���1+��T��]X��I5Ҏ-Єq�B�	9�a��Ɏ{�|yy��LZX�8񣜾dNα�� �=2��P�1��9��S��'�Ĝ�TÕai��[PB�D:i#��dL	N1V1(�柾"*th�����$ᐷRڴtQ4��S�P�'���y�+�&H���Vᗸ{�F� ���$0���+U*Xs�(�5F3�'&�A7&ߑ;��x�R�؍��{v<q�I��Y�tp��NU�L���7�����4w��qj� �����<:"挂.Rx,
�B�!�$@��P&��L~��Ϟ(�@%0�nOg6�,�ć*�OpA�0g
�,B��A�L�v���� �'A� �2G61��Y�'%Jb��L儹�&�ɀ)�~���'Av��׆W!P&�!3���)>{*��K>9����>z(��>�)3�I�j�{aNĹ*��;WA/D�P�w�Z�V�2Ԥ	?,xP�-D����"��Q5�BD8����.,O((z�I���q��xV+C/o��Yh&�08 I�ȓn+R�šH�6,��d+�pI�$��k�k�R0$��?�
5��(y8\�1	
r��=��A&D��i��ˎu��X'��*Q���s�����U��#��@�g̓'����к`�����p��G�}<iB�A�X޴y�BlC��=���0k)�E��+�B���9J
�p9�
ĥt6Y�[A�	�9Y �b���G���'|H�ԫι"zV�:a��]��'P��:����0�_`�`s�O�5��
�(l�N�"|2���i���0� &E�:�AM�<��O�*�l����N"S��H:O� ^���'��m����ĘϘ'�x��v��=��C5�0uvZ�@O<ٷ�a��?a��ϵ_@������5g��`��;"^0�ńO�K�N��D�����i�eʍG��,�ⅉ#C�tI���$u[�"?�W��)C1��#(}2�@�t�0�K)��1��H���O�J�� t!Ȋ�T��"���0橃&2V6<�5-������Nn�\�+��)§CfLI�aMb|rq�u�۷t�9͓بXvg�[��ӧ�����ԡR.�]:r��"ڮ�0��J��� uC�u��h(�3�	��| #`\�x=����+�"L�������AdL�Z�uJ�����XX��x���L�9&hY�[�pkT]P���>�J9v�׷����bT:-������L` Y�Γ�;(��lY'�ԭ��a&�Lc׃��E�����0-�x��#�e�'| ��Dm�#"݃�Bz�'^2ʠ���M�V���/�9�T8&��z7��4crqO��:��E�i�u92��
m� �� �C��Dl�V�Е&k����@)&~��k�!J�Y�us��(�8�ϒp�Q>�[�j@�Sb��XVEHd�lLR5&a�LU&��cY��y�
�%Tb�xG@�3��;Ō["a�l�����?1�M�8Qɰ-�I>���d�taLL� 6��bV�A���:?�ɺ�o@'"k�E�ē��)5���o_�9'�?%'�P�'Ph˲�8b��%!��J|���c@�vy�T>qS�S9���a�3�>�p�>�O�m���?k��rC�6���3��o{ʝ�� �,3XH0C�X>�H�'[�>��-m�63%��?_e�D��o��"=i�^��*��?��.�0�q ��<�,E:#&��n���,4�s�2c�z�$ӧ�B� @k��K��h���B�M�ģԊp�!�2}J~b�	�	T�4��4^��x����B�(�#\g� ��;�$���o��v5��(GOJ�$�'���w+�=B>�pR�d	�T�e�=�O(�}5A$��Z5���z;P�j
�r�z�8utsTJRSiP4��H_'I��p�N�9mY C�I:~x����Ɂ�;u�9�#I�ru�"=�����?�����`=��L|�\��h�ʖ�k�o�^nB��x�R�8��bV�1�m�0T(Y��*=��՚��S�O)��W�ûg/�u������ţ�"O�U�s�-W��A(5�*}�8�w���p*�	U�z�����c� �b�8]�����y��C 8�	�����I��}���y��]�
���H7�=�(@A��y��Y���)@o��=� �H�+ӱ�y
� �؃E�8�D��§��H� �"O�A�ѩ�b�"�J�@Y'[Z��s"O�$p0���*Rv�
#� 4;�"O�UV(8Ie���G�ŭ��8�"O��"�L�.(�`³ꕣ@�@�d"OT�o\6-,P��O��2�n�F"O�-yD�r~�@�GXa*T2"OԌ���Ѯ'N� @��y|�3A"O:��CƲ"�H8q��LBΨ�"O�в��ˍ|��Å(
/8>�b�"O&�CW�Y+`��eL�~B�H�"O�`Z�f[���ͰX�v���"O��b�R�I0��$51*�Pg"On��	i��<H����x(,� �"O�HsSL�#�ֵ��.���T"O��:'�C[�ċ7G7RtЀ"Op�[��Lf��@���63��]�f"OH�K���F�`xe�3[���"O���>��Xا‛N"��"O����K��ڄ��P̰8�"OJ5��o�j��D��K��lp(4"O@I�eQ*!OBLzF	ŵ0Dɰ�"O�M#W`E�~������k���q*Ov��`��H��G+C���'J���(bh� �)մ(��M�'�,� g;��a*Ԩر/�T�8�'�f)
��0n\�QĉX/W�%��'�d����AjP�n��t��)��'a�yK$��K%��XToE�n�>���'*p3f�����P�s!�]�����'�$T��.�n��M�HרS��J�'�00�	J�P�X@�uđ�<!�ȓk���+��?z*,1���O��Ňȓn�^�I�W&�ea⎡f���e��|3��I�L�|����*0ԝ��hL�H��#Ҡx��|#ubQ��������;䋁���$K���Gb݇ȓ+�d�3H�4}T�1S��R�_oN��ȓfHvH�ĨxZ�j mS;�)�ȓd��D�(`��b��ѩB�\�ȓ���*ӔIj)*��KA NI�ȓ)И�U�)
�Q 1?XN)��je5��h���R��,����V^	[1&H>p������/Jl�ȓoH½�je�f���I�<a�3D�`�����\   ��Cߒq�:,(6�;D�$s�oʁX*��	GݿY��a�$l*D�H
��'83\�z��Q3s�&D��w��5���Z�3G���{â"D��i1�,��5Рe�Y��5;V�#D�����}� @����}�F-+�, D��I�c�4c��C��W2�Tq9�-D�x��$Z���FF�=.��D���(D�\��@Hu��uIMe1h���3D�쪕#�ܦ(��+Ă{brT ��3D��x!n��4����({�Y2 m2D�\���A�Y|�����5K��c�3D�$�)�=S�X�0�' �d��0D����bLD&sf�@t� ���M*D��*$��A���Qp/ЍJ
�D�*D�<�`Eըa,��5�d�ְ#+D��w�Y)eRP�J�3jJmЁ�&D�����":aH��B�j�|d0�"$D��A��� ���t皣.JZdy��Du݄@0��Jx�� �J�^f��3Lͪ��3�'g��c�+��'R&Cw�ϑ*�4��&ő��Q�"D��!%�<r����s��8l�h8D) ��Fs�n� h�7��~���6J�����لg ���F�P�<��>]?hQ���fH��u$C
N���#�<1�nד	#���'=�)#A��;@3l��	ޝd � ��'�Bx�We�5+_�����O`!
�-AyY�h�2�	<mo�|b
�d,��8f-�_���H�(����<�!,��L9�1�?�~򪕞RF�%2)�g*N�1Å��y��]� I|!���P�@(�@N����\�0 ��MJ7��-^�^13mY;gѠ�σ��B�I%���͍�֬�'��u�����3�	<���ˏ�L<i���"=h���!ܛ#J��i�tH<)�HƇ/�}���T,Z"^m0 �]!v��
�0��2jVm8�L9f���Iޖh;%ٯr= �+<O�`T��.z5�O�-�Pc�%�� j߄c�T1Ҧ"O(qQ@��FQ~�a�J��z;�����d@�{9�舓�2�'�B堰EYX�7�0.9�q��WhAj�A½I��T3�J�/\��ȓF�k�CR&E�=�Wf��]��[ݦ��Մ���Ѣ#f�(L��.�,{���g�̉�6�Ȧ'� ���s^����QO�M���R��1�ȓ&l�Ѫ�{��a�К� ��ȓCk����ފ~���2'��P2,��6�������Yތ$1B*Y�M[Tm�ȓx�X7F�~�		vEG;eDB�ȓ��4��d)}�
���<G�� �ȓ:i���`�B=q0 �3%X:��5�ȓ �<Ċ���_�T�Ӕh�0
��>�B�C � D����P��4r\�e"$�RQ�<A��*�bW`��^�n=�W��vt ��q�|B�H����_�i�'L|�a��ǉ9ő��� ȓ>`�V��U�B�#��mK&Ul�DsSK�\�$���_6�p>�Ee
���QhF�J�$A�D�l?�&�@6r\JH>�S�@5j|�%��&@�D �ЅqG	Šr.<�Ƞ��L�!�D��Ht~9jQ��g)�B���.&5�I'�^X��ZA~�Z4�>�R�����S�9Q&$�1����2Lɑꖣ[�2���q�K�-Xy�"�4D�ڑq� T�����T%x*�XSL�$j��*M�q���^������>i'���Ɏ1y��">)��U�����w�$�;Un���8F���`mM�0ry�#�W)F�=�C�'.y 3cM|�p-�glZ>_�8�'1�(�G��|���O�I���e�g�ް�~�㌵1D8TX�F��h|��%$�y�b>\�BbBpj�[�|�O��@�U� !�h�FdE���	�+Np��ݟ|�)2�	�:0 п\(���'�J#B#ϓ��5�J�"^��� ��N`�Μ�b���OLh(�n�s�gy�ovF�$���~aT��*\���OZ�ˁ-	"�.<���d����d	"��i�l�[�F4�M��#Ә-C��d�(/l����ԙ]*@�P� Țyf�$��T���r!b&��Ӗey�H��\:h�R��nȞG��B�	9�$A��D�=Qz�0�B�MP�O�@A����<9��Z!fkz��'N�O�8Т�Q�<��b�)RL;���q�Pt���
D�<I�A<VVda*���i�@�Q��F�<Qv�ݽB�1�"F��DZ��A&�d�<�UOO�I(V9[`�9^lP�!�J�<�)9��xW���l��=A��r�<QS�5+z`@��!f�ƙP3lw�<�܍k���A� M�cb�HxS�l�<Y��<k��� b�5m��`��B�n�<1!�L-N�i*B�C��<�D%Ar�<)���p� M��`:�n���M�r�<�S��=z6���l���P{�'�E�<ieBH�%��a�j"1�����<� �	�ԧ�>.��M��Ōi���I"O$��7��/#o����A�?F�J�i�"Oj9q���A�^Z�aJR�X�v"Ol��˼2B��+L7S��iP"O���7gU;AP9xH:Z�8`kV"O8��n�pC�����:h���"O���&���6����K^h�J�#r"ONݨw���O6����-%�08�S"O��٣�)ʈ1�GV�1x�s�"O�0���Y9(�G�C���"O@H� c��X�`
G3��%"O4�r� ˡy`jDk4KŰG!��BF"OVl ��_ H��gjX_b��"Oi�0钉���`��P��@"O2�⦣�hj�T���D�k�USt"OHX�5�2bh��*� t�e�b"O��hS�
�H�ɃT+�Ud�؛t"O�!:a�2>ڐ%���jU���"Ox�d�)h��ps�U�NF��A"O�U:S��O�4�s��:z���2"OJ��QB�)X�F}��eֺV���R��'���pA�l�I;Ϭ(��i�3`�X�9�~B�I�SfDer���|^���$fD�=vH�'��La��̉izɧ�O�
�R��<����޾���C	�'�,k5�O�<�`=��̓�	��=�5��q����C����|ҕ��hL>63J� '�x!�D��)�tؠc�x1�,Q�8���N��*�_���Ic�N% ,��U�L�܄ه�ɚqp>1����-Hg�~�D�� ���j�ll��S�bЅ�g��*��ם!��5�냩5)p�'AR�;��VlX�O>}sb�J�l�i7��75Lj9�ď/D� �Ԯ���ٰL�;�j(�EʡH��s��R��
V�g̓"�-9jA�E��l��?L4�$�<ɔmD'�џ8�-�*]��[cf�d��qW�׬s�P��:7da{B#Β\�p����,��52v	��'����	֋h)��2Lt !�>�S���[IZ�j�#k�X��$HN�'q.d� �!JR	�}jA�3r�2�ʀ��"�D�IQ�CD~��W�8H��8��G�ᓜ^y*ՀQ/&�j�{UE�wA2�	�P�2"���UW�S�O?��ɖ
�3g!4�t��".�`j���_����F"H�T���Z�yo`��B� W���;�ͼU���@��'.�2o�F}b퐽4-p���ؑ	XMȣo~qx�c�����.1���Pg�,2���P�*�B,@�f�+��it���Oh\iF�A�6�&O�y�Ε;l�$y���Lx��I�Qg�,z���(q�nU��i���&aC�I�]�&����81}�'��E���k�S�F���̄�u�h`R���R��y��D�X�G�$6^\�)��<�eNz:�ԁt%��^���u�	P�'���Y`P�O"b�N����qe��"�0��'��:��	Rф1���JS8��j�B�o*  �-D
VSB�����O.,��Br�@�O����pcOV	V(HH���Ȥ��!i1868��L!�dT��D);�Ò�B&>��r���!�	
���b���8�_�G���!Y���O�yIAÂ�9Q*؋�m��H�����R�\5Ie�|ai��<����3�\�CZ�M���X�@��г��^�8�=�O��}Γ}1�ѪM�X��e����@���Gz���;���8��l��gݴ���
@1\�,�ˤa OJ|ϓ)�
��)>N�����**:,�g�1G �XbhE2'�v兆@�R�s�ȀD����#� l�t�i��Z�[��"Xs�iK, ��h	�'ϰ�u�@3����eN��T�u��O^�)�f,uк�b��˅fZ�Բ�{����:��D�2�*_�-�)�1�'Y�Q�#�5X��X"�k�9���QOR<'w�1�/eh<�1��|fh6�B#A X�`+�K�'0X�(�i�?0�����3���!"���0��C�<1�	^1���3�^��]@�c�3�-_:��%�"~*֎I#JK�0:n�+M'���`F��y�!Nh��˲cP�L �TJ�ꛓ��DG�G�D���S�? h�*v� ]Hv��d��>WE�źF"O񁅿�\@.���*�dd�؄�)!�pQq�[*|�����;{�@T����بfa�>Qw��K�i7:UF�������Ъ�,!�M�Q%T,y=���X/��1���,H}�B��/l�hL��X�t�a�]�x���s�������=f�B�ǉ>�s!'�y����v�R�̕@*�ԫ/�P��T&��Hp�n�@;`� 4�6����`��͌�6U���MVUBl�ȓ<L������+O��
$,N<�`L�ȓb�����A�C��Z��P:Cp�ȓ>S�9K�� <��$��4t�r���k�d��p��H��̻�J�	P�5�ȓ+����(V�w3p���2t���ʓga<e��\�� �F˒`�xC�zmN�s�
�a�M���R�fB�	�hkL�֫��i�~I*C�	6D�L������ر4��-0�C�	(~�6mB�¯$d��#���0,�B���ݚ����(t�0%|lB�ɥu��06�^�]��A�mɯ`�6C���$z�/۠2(�,Z�ɛ@�C�	�U�
�%jЬn���p*W�1c0B��WD|Ȱ'XI��}���	u�C��a��
�WK�`�� �V� C�I.YH�Q�t��>�D��SW�qC�	�f7���c�..�
����J)0.���^y�
�C?9$�?�h���� �RAP����s1� �vϛ��~�u?q$�}��M�O)� 9���2��B���H:h��':�m�'i a��'I�#~ʔ��8c]0J���<ݶr�!�L��Sq�p�v�i �O���7���6X��J�
^H|(i�G�N>��P3T�<E�D�
��`Yx�� /�u��%�	��t�1�U(�0|�2OT32X֤P&�w�t���F���'�v���f�A>�IAGʯoJbq���E�X����au��	�.�6M�����>]6:!i�/�j�����-r{�SR?��]��%?�S� �z�=Cg����� ��$
�qOD�)��h�D�X�E1����;uL�[g�'�O��Ezʟ� ��W�l�,��e@��L��!e�d�H���O�n���]#O,�Sb���k$%C�O�qr�)�'T� �j'��=>ܤ�8�b��0@5+R(vc�O�?�2F�7����%��&5nV��q�D/��'?���S=j��+���"�X�|M����A_�S1~��,���M��kq��z�X�'��#=�r#�Цj����Gֻ$S�p�2)EN?9��'��|`i��s^4����\SJ����d�!����IFq���c���*�2z:d�Ҳz;�{*�.����G~��(�.ݚh^Q�f"��'6Ҹ�p�<�i>7-FFy2�Ҁ[]����
�]l�Q�j�v��I�^���S�O�؂��4��3g`W�,� �s�8���@� غ�~�$+������?	�X��a�l�
��6��\|��Pᯟ`3E��51����
�'<��-{Qc��5�v,JSJ_>o7&UɃ��25}SC�>��O4��d����W.�e"��r���+-D�xB ��9�6*���~���!�+D����l�7x�8��0ᖗn>`qb��(D�r�'Tm�hC�VX�X�(s+:D�Bw���n� �@�)8Yx��b�9D��D��+�]pVH٨kL<lA&`-D��YF�#=�	�v�Q5���A i?D��(��%~���ՌN6d�v��';D�l
�,�p�z)�un�~�FMڴ%D��KЮ�ZMZ�d�>x�d�J�5D��p����GH�R�g�{�.�ڃ2D�� ��(���@(a{m m3��"Obt#��l#r�Z���*2�	"O���3 Y�q1`��U �%�"Ol$��b�1"�v�ؗ�V�=�H	*�"O �Ǣ$]�t�B�|��"O��y͊@����N��Ӟ� 6"O��i& x$T����ż�`P"ORiraZrU腰E-�Y���"O��H�
��+� A����$��"O\u*Ӡ�8v�Pځl�E|89V"O28��l�4:��X���7&���`"O��Q7A�<���u	ʿ�B)�4"O�M�B�֚m]����C6��ͨ�"OF�#NT�P�:��f��2ɮ�8�"O~|���ׄ��	�7�֟��Pa"O����5��=��E���$(�"O�S�C�I���5�I����&"OF�Y$�H+DP���u�@��<��f"O^��0�S�jp���u-�n��X�"O�h��P��B)0��B�!����Q�Sh�1��A׃�3m!�K�>k$Ḷ�G=h蔡�E��9l!�D��d��HG���0��1�пz!���(~�� ���)c.����J�h�!�]Ԫ�{7��3-��ܹV`�u�!��	�hؓ�)Z�����H�e9!�D� ^�a��8Cm�آ��<�!�I�kl�a[���JFM�2�*�!�$�-���k���`�A��w!��+0D�=+7i�!?�8����!����`@�"�)T_���w�E�*q!�>�W�M;&XP�ʴ�U8!�䇬}5�|Ӈ5-T���a�:x*!�D�-4����D� �G|�0�쎋[&!��D�Xz�̃����+�r�����}�!���n���$f��Zz��%�ܖ�!�\:"���8G��-X��E���9Z�!���,q�}BUH��|����G!�$.�$%�f��;8R��rmJ�*�!�3^)ZX�W�X	O���j>t�!�c��m/G����)Y'!�$M*��!��I4	g0���)[��!�TVh2Aԁ�?o)��z��Ա�!�d�/NDִӵ�y��VBї!�!�dB'R�:���3T���R�Pyr�O<�-�&dF*Fۜ�3m�,�y�!5��]Y��N�24��/�:�yҋ���0	����R���ó�˕�y�B�_��E"'dө}�.���X�y"��3;��TG�y/dy��NŦ�yo
�VY�A��>Ĵx�o�4�y�����U�P "2�<m[5H�y�o��+5"�Iۋ(�t4���1�y¨�eF���v�T����>�y�4JKZqӀ��lYz���aO��y�KӹJ��h�	 	p6�9��)�y�aeU���e�;n��]��$U�y2� p҈d�B�X-3NX� tO���yba#$�ܝ�gh��'t E�SBI��y�&X	�̡RF�:QX@�M/�yIL�"^\E)���,�����yRL"n��Mځu\�L4�yBc K=�Xȷa՚�1�	���y���p�P�ͰT� �sS`��y
� �O��m�@`��۠+W�<X"Oz�����N���	w�	�:H�Y	�"O,�٠�ǧ)��q�2��+�xܚ�"OR4h�lNF��1m���S"O��c�BdI��-}����"O>4��(E?%�� ǈ��ڲ"O,�� ��(��-���|�`A"O�(rI֕5�����{d6�b"Ot�p��-QsnD�5*�q��1i�"O�� ��o�hx��&F� �0�"O^�
d��1���tY�S��"O.���h�)R%�fa �b�"O|%@b�?�IXC�^�LlQ�"O2Љ$.�b4:�H��J�n���"O��FA�2���"�A�����"ODA��k+��1��3�v�Y%"O��g5o� Asc�SA��L�"O��x'�׋t><�	A�1�\�4"ON�r7'"�DY����mu� @�"O��H�<t˦㜚LtF�*�"O�2q���nͰ#\'q�,��"O$`���$8fl�s�Mpl�)"O��!��^L���n�$?c8�p�"O�U9פ�JR�JR���ql>�	�"O����M��,.�)�֚95l���"O �
��K=&^4Z�;")n	�e"O�=�M�2LҮp�'�:#"Y( "Oޭˤ���][d(� ��=Zx�"O�lC���W�f-��T&XpNtJV"O�$ �k�
=*1��-C<U`�}h�"O�-b#^A8Ĥ��Q5c[扢�"O Q�D�m���ʰ���i�4js"OX���:K�88�&� E{�"O��	��q�>Eq�X/g}v0T"O���M@�.��q��]d�ə�"Op��v�14���P%�[H(ɲ�"OΡ�4牅=�PHƕ�k%����"O���
U�@E�T	$��"��9�"O�y")�}�Q&(׊�1�"O`ХP)1Ө�5�
3Ӥ��t"Or��o��j$�0aQC�-�8ٓ"O�\��C�j�䔛�(����"O�ycBɋO��i�e��0\A�"O�Y�f�B4"��m���7��Ջ"OH�x�D��~\Dcӄ��=�j�r�"OBݒ �R"�2�:#c\-B-���!"Op��J�2-!����S�^ (��"O0U*2Ǖ�d0�Jp����(�1"O9�$aI�fΩ	u��k0���y*� �����	�|FM7�y�FA�v1-4��% )}J���'�P��C^i"�L��0F����':Ҝ�R�٤IJFxY�����
�'�zp�S��`�����"Ȑ�P3
�'�ƥbG�=����#�����'�|mc����� ��4'Y�J�֤�'�V��R-U�R��"��C��H�',~�1�QGT�rp�ϲ6��i�'Y��BC�$�����M#)��Y��'�,�#��kP(m��NՃG�y;�'����׀HKm���*��8��h��'���#��?)�`�� ]�-/`�j�'A��$tkČ��)w����'�l��dDM�7�@�`%���Y��� ��X�$Y�[�z��sኀs�Vų"O^<�H�Zu��B��� �"O ����ܒ�(�gW�|��{�"OҼ0�(\�Q!`����˚N��,�"O4=)%���E�N�K�d^�4��"�"O�u;�-֧c�*�j��=t�:�b�"O�bCY�Ur:ثwO��0���I�"O2MӒlV4z�U��g �n�Z��q"O2���g]�?e��̞�n� �@"O�p�4o���$��d��A���"OLhð�̃���H�C��l�c"OH���oˢ �8�LF�'8�s"O�!;e��'T���
��	,���"O��Z�/i���	�f���"O�-hs�@�zHk��#�ە"O�`�`�$g��}i�G��/�v�ʣ"O��A���c���a$E�0�3�"ON�G��f���C@={ɪ1B�"O�z�#G.^�H� `ūM����s"O�@��J��9}^�s@�P�Z�n��
�'2���P�I�=�J��Iį@��I��'���p��c�l�36�Ŀ?3��K�'@ �#p!׍H����`�B03����'�5��lS�[�@)@�T�p���'vn�+QbY�
o��y�,[�S�@9�'4��*ZUi ��sI�""K`���'q����G�" ���pᎭ`6���'�1ؔ+:^�<����д�'�b��AC��$��qq���(���']�l�W,�?���	'���`�'� ��"��-i�v�P5Ƒ;$!,�
�'q��	����,�c�B������'���7i��LX�pƌX)�z���'� `/�>c�ؐ�����.�X �'�b8�7��8��!{�O˷��E�':Hu�敘c�F0��J�=T��)8�'�b��$��~{>uR�C G�X��'o8�	פ�*�V/�
M=����'����0�&'�jm��,@G1�(a�'Ԡ��f�)ЫS�=���'�x�֩�.�P��3�f�k
�'r����Vf���іU�-<v��	�'�h��T˫B�����D-&��	�'{�!�C(|+4�+�i�"�|dI�'\�J��<.nl��/TR��(��'��P�D�ov���∩:����'�QQ�M0 �հ��Dt�X�'+�(Ap���L@�=�CX~S�\��'�@4:��޺O����O��m�d-I�'��P�G�?B�q12'P�p����
�'�ֈ��γBIh��-
�'���Rd���l�Cl�*'+ lK	�'��Є�׸a�&�Iwa��d��')�ň�Mv<�A��@��&�&i��'HHX�t��Cu�t0���`�	�'�}(�m,r�<<�!�G�4T�Z	�'p��t'�%ef�a�d@&~�t(��'K����풕iu�U"�E�~� ��D�O^7m��!{�e�n��q��?����?��ܟn�k�
��{İ�ٕ��h��m
�p�D�ܴ<�Vț#&�N�D�ӏ�(OH��g�(*�v��iŴ]��I1�l&F2��A)	�I��آ&�P����'*��1�O%d
�����H����̦��	�X�Ѐ�I������OB7M�*�j�a$G�d��] ��J/���'�O��8���9}�sk	���3S��<a�4Fk�6�|��O��\�<d��D�:��ɍ9��+%�!�^1 ܴ��<���tm#��7� D�Hb@T�d̨\X�/E
�9��]�g��H�Gf����C晞m��<���+�[A�ΞC��Ĉ��&tFf��g��*<7(M�~����	�$z�ۋ��B�M3a�+os,E�3�N���8p�,��6�3��	˟�	n�IQ�th@�b7Vd;���=_��0�6��yBˁ�n��|���"a�>m� �#��I��M���i��	!����۴�?٭O�+UP6�\�z1��"Ҵ��	���]-��|�b���8K
�3��*e�P���g�kc+��_X���CZ�I����	�-3���`)�;o,,�����YLX�b�O,��Esv�\�_���
�Iv ����,���O �m�����5fL���	8��a�e�	N?�j��?Q������f���Y�8�Z<�B'�*������Mc�؇T�z<FB�'�=*eiQ<c�(}`/O��!�*��)����Os,��'��Vh[���Уs(ę�YjFnJ�t��I��h��]�\�L��Į�Ŧ1�O����#��'�Y��B7I�(�S)z}R��2Hth-9�dQp��P�M�8�Dd�4�i��J�9�Yƅ!.8� �ON`���' 7mU��(������8��17亱*�J��� �O�� �I� %�4�0�Z3�dh3�AE/ҡ�7�.ʓ�?� �i�67M�Ot<lZ~�d#ɞKC��y�ă1��9���]<A6����O��'i���{���O����O��$^>�y�EL?O� 1��A��XX�ʑ*;���)Bɦ=��eزɒ��ן"EyK�_$������7K�ThᶊR� �:P�d�0�Ȋ�GW���J|�4��S≛0�yx E�gWЙ�Ѭ�>yR���iR�J:GBIOJ�<1���MEJ�A�)V�?���  �D?�e	8���оMRz��u���qP�0O�6��!$� (tl��?!�'X�`Y��F�ƤH���7'���+BBD��~6�"<O���D�@-)F�Z'dX���Z 9��'��Mj�C���3,!t����*Jrp��3�	T*rT���/yT��  ��Q���=�БE�>t�y����:����P/.�\�Qo��U}<���[3&��)ˍt�Fɻ��i�v7�OZ��?���i]dD�W
J��Hj2��3T<�0���O��.�Opm
EL�u�� ���@�}� ��"�>� �bɛ��|�$���^����   ��   2    �     �+  �7  wC  �M  X  Ne  �m  t  jz  ��  ��  >�  ��  ę  �  K�  ��  Ѳ  �  W�  ��  ��  =�  &�  ��  G�  ~�  ��  �  � [ �  H# �(  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|���K?I7��.�� K`�j���k��H�<)iE>'l8�7�&��{B!�|�'"9D��g�P�8�3_f�*���yRiWC8����	
��Ms�����O��M��}���X/t��<�lȱC"���m!�]��e�X�A��� aA|��x�El���'�ſ$��x�ĳ_��H�d(4�$����?h74Y�ɚ�^b���+Lw�<	��$��G�E�<6�h��X|�<�Fp�v��U"�YE���u�<�G��[�ޔ���TK�"Q����t�<A��KSG��$dD$�tqKDeMV?#�'�E���C��PP{��D�1��e�}B�X�ɌK�.��� ��<�1�〕Q�B�%`�PXPc(�:�n����?l� b�ҰB.�S�'"~�Z�l�KHd�Wɟ�W����O\�=��ne�IQ�p�H� �b.�%��.�a��C�I-f�f(n=Ƒ{!"̀d�r�<a�1z�p�� 
K��(�i4����B�Z���*&&����K�*n@���=p��{5��?\P���Rm�����ȓE�N9��h4q�P���bI�@�:���?q�����<:&I�g�ߩ1�pA��̌	�!����X�"V	�;�:L
�+T
�!�^��eI�D(`�F�ƣحT�!�$ɅS��u�V�� ���K��Έ)7a~2S��W�ʄ<��H�Rk�%* ��W/�	%b"~zUH(%J m ����M`�M��LS�'��8��ӁL� J[�Fق��E8wX�B�I���Sd���`��`9>�D�<M>E��� V�#�+\�Z�bUMi�főP"O�}�� F�6�P8�V��]�F1�"O�ܸ�BЙv F�� �"�2H�"O�p+tE�5)�~�+�َ��-H�6Ob�8��	����Tk9؞��!BM#g B�[� @k�E�N�ͳ�I4p
�����HOZ"=�'�Y�Hv��X�n_'�n���N�S�<���ŮD�PI�e�%C��� 6OCv�<�T�(c��P�M]��\�`�)�r�<�P�ʭd�.�	����v$�u�E�<ѓES!q��I�˚ĥ è˂�hO��i���>)��џ;V��ˀ��)�>E�WF:�y�I�Μ���I�8AWM����hO��xt��Z0І��Aߊu)����'�'�fQ�f̗�6Y�)Yr��c;ɹK�T��	����S�	:�����MĞ#>ɞ'֑>��N�i�!X�	ݓ5��ɁI2D���0fI9*X@J�)�� ���/�X���-'�x()��&,��퇄?��$�ȓd��@C�b	n}�}��e%O�� &�p��IVz�um��ʐ�h�B���Z�'���#A�ڑ;��JCǖ&J6@@��'��?�)� ���.wD�0q�C��KJd��I@�'��rs�U�5����N&3�Bء*O����8	�*my`�I6g�6 )��VKa~�[�0C'O�)��D��ٻ2��xZF�%��ȟ�4!��&,�T�I�^c���"OL}�o�4 @�b�aǟd\M:�"O"ԊT�=SMb9 ��I� sX	�&"Oy�����F%ԥrw��Ab.���"O�h�5\�B�Q0"I�p��8P�"O�ȨU��"Vu�Aa݆]�vqI#"OTA�O�*%p� I�2UBd"O�q��%t�|��@�ܿv��x�Q��v���		/L4uq�a�s�R��#��	ij!��֦��E�w��E�}�H3�!�$IH�������Z� �E
�!��@�-�����<!�9�a�?E�!�,2�-S�!�߈msa!�:Tar�OQF�V1vOp�	����lu�ġ�"OnE9�k؈n�^�+s$V�pe�l��	^X�0��LT�s$� ��
�Xu�ҍ/��0<Q�b��NP����Ùhq��P�g�[�<Y����?��0��.x� �v��X?�	ד���φ/�L����Y�3�ּ���I:@�!��M�xКp� ǘ%un�YK�(;ax��ɎUư�ځ�ײ`Lvq�CF�=}�C�ɎwI�dZ&��� �X��#-�nc����B�Ş��hb��dK�d�D�G�1�|�Dz�A!O���6��)� �%L@�P�K���V��Tʳa�*W�MyEaA�Ff]�U��O�Ą���Jݛ6CԳE�L �A%ߏ%6���t���0>�J>�"�0ka�9�p!�_�4H�#mRl�<����@@��W�)9t��7�[d�<!� F"n\���T,Vh��h��Va�<iQLK1{F$��E�q� �W�<9�dR��U(_/-��(�j�cў"~�ɰ@��3�.;x��rC�2�*��p?� �C	j�4y��F����)�rF��<���P�lU�$�0k�e�'�'[Kvm�?���ԟ
�n�۸�b0kZ<%W@�y��/CS\#>I����)�\��un�&��4"a���+ޑ�P���H���$�"an
ԡ��C���ů2����O\�"~j��M�q]�A����1>D�cÆ��J���π 2$
�/�)~��t*�mz�b6"O21Y�o�G�xXBL�Ze�eK&"OF�)� �.����Kܝd_2�p�"O,q�a	f��8��v��a�"O\A���
�v����cK>r'��÷�	�ȟ�u�퇅��5A�S)�D�(e�'I�Ƀx�E��n�m�w���A�"C�	��,=J�@�9
�� *#*�,����?Yݴn�:UExJ?"�O�+f���Z6��a^d���'�ID�@�'
���f]<,�T��镈:��	��~"5OĴ�	�gIJ����A]Τ8�#%꓅ȟ4�Bl���j�HZ:8t�:1OC��O�=��UXT��ToF;M"N���kQ>{HL���Mˊ�T?a�<���b˜��@�B�{�o럐D{���͢ �F����"�����EճF������h1�S�ӒO6�Y!F�%p_��飬β+�rʓ%�����ֆ/�����H�u���慇�;3�{�-�D�|i`3P�V�2WF�vD�c!��8}�J�1��Ӌ>�Ū�m`�0�O,�k&��~� ���&-���	�''��&�� �B�j�%��b
3t���d<D�<����24�r��Cφy�W�>�hO�-i/B����R�
�+E INm�C�	��̐��A~���u�ȓug���dR�'�0p�KQY�`���8�^�Q�'�XAR�[�:�{,@�u">H�Ol��4�)§yX�YS�K5'ɸ�Î�*�����t�'��a��	�Z��� �-L���h���%<OL�U$�(Gѱ������&"O��ᶥ׶2���A]B�Ȇ"O��2�-H9Nbȼ�^7�&�!�"O���I��[
���O�)4z���"Od:��T|ⶼЦ��$	�\8[V"O.�K�섭o��`��Oǚ.)ID"ON%�R�N�@TV��O��(.�s"O(I5¸e. |�%�T�5"O8�:��̵'L�4�wl°#ܞ��"O�HS��ϧO &�I0,�e��X�"Odurũ��
"�%l�bʴQ2"Ot���.�79AdmS�h^�\3����"OR���F 	RL��;����S/�M�e"O�PJu�SG\���T�,�+�"O�������@��Aګv�X!"O@�X#炗n�\���V#<T���U"O|e;�ʝ�2��u	���/�\s"O:u:Q�� E,��ǥ�+~�ԅ�U"O�I!��VK�����ֱ)���b"OT�v�	%(��-�ub])�F�)�"O�-���56>b���ʑ�w����q"O���� L�p��Y�F� 3����"O�0�R�O Kߪ�#�KJ
�Dy�"O>��ȏ�t(~ ���I�Lx�(+$"O@)�"V�����)%:g��P"O��03T�z��ՀeIÝadl�"OJ}� �!Y*�-{wf�*Q�5"O
��D�J�.�b|H����XM2���"O։���H���1z4��0
�x}�E"O���
�?Z����ҷ���f"O��� "I.����l�G�L��0"O��*�����#"Ģ'$Z�z�"O�0�Nʴ�l"���2Ը�"O@p����%q�J�
� P.Ȑd"O
��pLÌ}Z.�Bg��QO�c"O*�co��B�T)��L�Z<��`"O� 칺qeH�uS��pӬP0Ui�"O����	Μ>{Z��ӭM�lr�"OJ�p��ۥ_��w	�&yF8�`"O8����?��Ja)P�7� �"O�t��Ô(.�u�.N	1�IAb�'�"�'���'���'Gb�'/2�'��@��H�:��	C�+qjղ��'���'���'���'���'[R�'��� 5�ܮXM�Pi�ۨ8źHcw�'��'�b�'���'W"�'�2�'��9��/C�B��Y��97��k��'���'�2�'�r�'�r�'���'/��� ����g$J������'R�'�2�'���'f��'}��' ��)CH�>r�`1�G�;��Y� �'��'��'XR�'/b�'���'+�L�@#	Yޞ��2@D�u�6]�#�'���'sr�'Z��'�R�'���'#0=97#�k��d�L�	��<���'1��'nB�'���'�"�'_2�'��lv��8�f�x��C�I�*�{��'1r�'R�'T2�'���'���'6� �0'��9�tȲv�� T�xt�'l"�'��'���'��'^��'b���W�q�B��0xu�C��'u��'��'��'���'B�'{ ]	V��&
�0���!mu��V�'��'�'B��'���'��'Ĕ	S7LG���k`a^"Tq"����'���'mB�'.��'?�J~�b��O�$�6���Z0L �Ҭ.�n�+�EBy"�'��)�3?��iA�|������p5�#�$C獼�����i�?��<��i�X�{�L�(���2u�J%���:��uӺ��U�J70?��`��C�Dy� �8���*~����Њ^=_r5���͘'�Y�\F����\����
�[�,�P��Tm|6���+#1O��?�!����3h�'1�i�A��7�t�;�g�1X��&ju�F�	`}��D�@�QT�7O��+W�G�-���ZVK=����#6O(����W�`����n.��|j��8<��[�� �����i�H�'�'c.6�P)vx1O������^�p�S1�9�,�ГC;��4����զ��ߴ�ybQ�H@��27Hz��Tsq����7?�4�ͪ'��Q�GB̧(-��Yw	&�D;!`@�t�_��}1
[�@Vʓ��$�O?牼d��4��LY1u��8*A���Wb��I��M���T]~rk~�x���0S5��z���f�Q�b��I�M#G�i!�^�m����,�fP�hNe1# �F��IR���;!ʘ�SdZ�I˸��7�P8\kZ��$A30Q��xtؽw�$5�t$-Rxz���f_�]��m�ϗm��h*��0x���p�~JF�1ժ��8�r�����-F�g�Y��B�� Y�ru2�c�cs6U��)D1f,�!î�`Y��+A�:AA�FS���J�� q��@�T,>ylU������6)U�J��RE��c��H&�J��y1%�xR^�e�@�^�t��r�_�G
a�d��W�Pԉ��A6���9�'�lz.��	�\,h�#�i�@}����3 ��Dq[4�\�*\+8�aiѴi��'CB�O��)�$��̅����n�e�im�Dy��N��O��aBQ/��4�z-g��D��x{��i��	�xӦ��O����0'�8���zr�BL�f,�)�Y�L���ߴ	{P�Dx��i�O�9�3	�?���ȗ�m�ԠU������Iߟ��I�N���O<����?1�'�Çg�<1\����+\�/v��}���.��'���'B�V[x�䃄�;\�9�(�
I�7��O�0�'b^K�֟h��t�i����C�6�H�H@JN0�@�Z� �>�৕G��?���?y.Ot���g�<Ta����-7�i�G�jq�]%���	ܟ'�ȗ'�`R�F�1h�i�o�  �bV����'R�'SS��z�oX+���`Z1@��^��m����$�ē�?�I>).O%{�X������py&p8�Gx|�u��˽>9��?!���7 �"E$>y���I/&��A*R7*�=���F5�M��?a*O�˓M�(�����J9o��(�ˉ3o�p	k��[�+����'�]��#�@����'�?A�'���@�)a 񳅧Ǿ|T�0��xr[�L#�"�S�Tʚl����ިF3*�{�i�+�MS+Ony��
ۦi����d��8��'w����F)7R�����e���ܴ��
3��b?���f������gLH�zݻajk�ҭ�Â���)�	럜�I�?���}�d�(fx�L�D�_�7ݐq7㙵E��7m�A��"|Z��b�Y�+��#v���S�rd:�Q�i�b�'2�Қ;��Ob�$�O��I�5��p��,�(�A�Ô9 �c�\u�"�I��I͟8�6�$>�ĸ�X����+@�p@l�n��(J׏�ē�?Q������(	&���!��
n����Fg}�P��'yr�'��\���U�]�6f�QG)�k��x%�ŪD=©�'R�'*��|B�'+�UfzZ��癍Ml��f���q��|b�'��'|� _*���\<�-�WN�W��9� �כur(�lZ����Iڟ|&���	ڟ �s�d?��A�`��Q���,����l�I}��'���'��� ��|�O�r�1j�����77���p�O�,6-�O��O���O���5���/9_��V%�Q�`Y��H�\ܛ��'�2Z����&V\�t�'7��OR���q��@x*q�5��+y��q�$�D�O���ZJ���g�? �ԳTʐ P2��r�֊0�\��B�i��I�(�H���ƟL�I韴��TyZc�$؃��\�X�(��Dl�D ��4�?I�,�Ɋ���������'�Xh1���?�M�����?a��?���r-O����O�e(����Y�\�12�ϷrO�����Φ1�"�^k�S�O���^6z��vFA�"������
	�F6��O��d�O�E��A�<1���?���~�<5�x@��[�al��8"[K��e�~9JI>	���?��xj�;Q��+�����W��k��i"��%�	���ß�$���*��<q�	�s��ur�ȁ/��yU��[O>����?�����S�t ciV%�*p˳)˪+!�`�-�<����?Y�����?Q��rpg^�!Xh�z�M�n4�e��������?��?*O�I e�?�*�˒�s
�LAvD�W�X�Ru�|���O��d=���O��D�:���dB���t$[����s�� ����?���?,O6q��c]q�Sei���.��!�� ��=9t�Iߴ�?!����$�Op�'�?�J?)!�e]�	F��g-#h(����m��D�O�˓j\,����d�'��\c����$~�6!��IE�;Ȩ��#l��˓�?����?!����<��E&�b���11}$Q�u��?t8Dm|y�$B56�7M@T���'����??a�&�?	��1����b�%S���I��h��ɟ��L|���i� ��FGԂ*����b�J-�0��46� �Be�iOB�' �O@�O�)V�4;���R��=8[ZDQ�Z:[��dmZ�h�	��D�	YyBW>��ٟ�c��*i�*�۳,
��.����>�M��?��Y�8���x�O�"�'��%��l�%D&����Ո<�8�)��g�����O4˓z?��I���'��d�=b;Ș�� �=���Q�Ρoɛv�'� ���R�K��b��q	'D�PɹǞ�w�hxh��ݐ�ēZ�,�<Q����D�O ��,6���)՗(�4cUCP�� ʓ�?9����'f"�Oj�1�ϟe�8�C�j݄b�
�7�i˘�O����O��D�<��+L=��	ޏ`���ԆB1B�����(���������D�'�"W>�I�^����Ӯb\��2/�.
J�1�Op���O��$�<)!BX�Od��t޶#ϐ<���>�xxys`m�����O��?���N��0����S(5�vݨ�M�Tja���y6��O&���<I�X�0��OOR��5&��P�I�.��R�:�:t���ē��ʈ�t��+�i�?�h�㊒=�4�(B퐈~�(�q�d�~����XƷiOL��?�����( ��L#H�#�F��G��Y��6��O��l��dVZ��'��TZ>7M��e&�qǠ�#mgx��w��9!S�Va�	S6��O����O�iC�i>!3Q.^�9�:P�AdB$u"茋�嚴�M�C�T��?���?�����*��I�9�j�PI��"���Z�ݥz{��q�4�?���?Y �G�����'�2G�W#^Q��*5g1렪E�q��6�O6���O�ыT�T��O����OD��4�Ç��U���Um����Ϧy��H���K<�'�?)���� �d�A�Vp�P�A��;���n��x���Y۟����d�'?������u�@!*�/vk�.Tk�M�R�e�'�R�'}�O����O�[#'W�Gx|ezq��;`�m2d�Q"\$�ȃs�d�O ��?QT�]���P�+g��u!�+W�^-I5�^0�M����?y��'�R���F>*}��4<"��ⅱP`čZ $�)gX�'.��'�rP��V���'	2B��)�����i؋t�`4��iB�'��I����5Ymv���p�Ik�����`�ah��%0��'$�	��j�u���'����5VbZ�x�`t0 [<=�A�n�0���?	�U[�es�`�s�S�djW=Mܺh�bӢ-�!1�)N�M����?�e�0qE���'��'����O(�@S�K��I��*�x\AFą�V����?�hʴ�?yO>ͧ��S2���@0�߼*������<>��7-�
&0�o����ퟴ��?���ß��	�p�X�A�K9�T�ѥȼӞLh�4&.H5��?�/O�)8�I�O����F_"�Uc!�^�Hꄘ�5�E����I������v��\�޴�?y��?����?�;6`ځ�� (lHUFI	���mZG�I7ib�)����?I���DY���0��%@Tz�1F�i��n߃zN6��O`�D�O��K@���OV�z%��t�r5�uO�d�5��T��fu�<����X�	�����l�Ʉ&�KF`@��!HȦE�^9���C�M���?����?ɠ\?�'n�P�eȢ�
�%ژ)�\Q�h�'�R�'k��:��'���'��1$�7-Y�	�T�J�=F����s/ n�ן����@�I����'�GP����
��}�0�iW�
c^�2U���6�������?���?����r,�F�'?B�>�RXb�|
����
�6�O`�d�Ohʓ�?9f(�|����~��ʹW�L��U"�+c� M�M;��?y��?	�Bז����'���'�t��AL��� �hi�$
�7�|7M�O\��?���|zM>��5��g��{�:�pe��=}j8c�q�����O�q"��ͦ�Iܟ����?��S����5�1��
 �z.���pJ@����OzTKc��O��Y����'��S�6`jT�5b��7y�-Z�N 7��?S�Ʀ��	��p�I�?1�SϟH�Iş`���� ߎ@���^5|���,H*�M+AP��?I���4�"�� ��G@�? Z�c�oD1:��L�P��y�<MP�i���'��F;�6�O��O��D�O��K;zz� 1�� �F�l���'��	�������	�f���O��9Q�ѳQ�RH���%4�l��N	٦�I1h�.x�ܴ�?���?!�g��P?���� �a�M��(iVc�R}BC܇�y�T���I��	ҟ(�	�yJ��u��>l�PA� ��œ�� ��M���?���?![?e�'�a��iba�><L�P�b���x�'�	ğ��I�@�Iϟ�����M3���"����Љt�ҩy�mǸΛ�'K��'_b�'N�I���Mu>)����/O ���P�@��;֭ ����O��$�O���O0��(���I���j��e���� �7Gб&"ܨ�M����?�������O`�+�1� �$���ī�42|mXU��� B����v�����O�$�O�������	����?��u��0Q��0l�,�,X��o˯�Mk������O�yyR5�,�ľ<��a�dcW0y<�����]�6�k�n��O�\�b������ϟ��	�?m�Sߟ$����'p�PT�A!Oͮ�9"�ɦ���O�0�'��O$���O��Q"?���OnzArTÇ�!�� %,��Y��4��� �i;��'��O���'�r�'��ȡ����d ��J�%�
~Ӿmy�G�<�.O��S��"��6���EPQ�d)����M���?���F�~� �x��'��O<�w덻\Й �\�7$L,ӷ�i��'h��+�����O���?�9�o;�6���XW��"w�����/[(&���Iӟ$���>熥��E��y+�,c��͒y2d�p���SI>��?A���d
4+��)Qr>6�ذi�b�6M`�Q�FR�I�D��I�	�@�I�.)��� �p���O&��l�E�b���'���' �O,��2�v>i��
�\pc�OU�<t��J�>���?aI>����?����6�?QO[�|/���A	0VKF���q��OZ�$�Ox���<� ��vŉO�^�o9b�SR��v�R=cia�6�D.���O4�d��p�0}�bƯ�PA��b��V2L��^�M;��?�,O����H�����ӫ�č%�ٯzg�=2\~;(�AN<q��?��� 5�?�M>�OD��9�.N M������-i̦��ܴ��䒳M�8DoZ%��	�O����t~2-� ,���K``���ڮ�M����?�BF�'�?�M>����8>�BY�&�_R*��@��MK�˒+ۛv�'���'��d;��O���0)�
����%8h�+�ۦq �*v��&�"|��N�Ё�F�H�'^��x��2c:	�4�i���'I��&m�O��$�O��	;V/�����S�<T���ɼy�6�%�dۣy��?I�	䟠��5xH�F�S!I=���1�[�CB��m���2N��ē�?�������Ê�TW��K �
0��T}f�9Yr\�@�Iԟ���qy�E
o�p�9��7>�x��B�u^�`'���O(�$#���O*���	
N�4s�O�������g$���e0O*��?����?�,O�	�˓�|�i$w�p�-S3lꈄ�U��W}��'�B�|��'��NƮV�r�)0�dp��*w��!�
ҹ;�ꓤ?Q��?�)OD����Sq�S?$!B�������B��M�*H�ٴ�?�O>���?�GH�>�?O����Ӕ �d��+<T�*�g�yӶ��O|˓^���;����'����
ze6�:4��".���J�rO^��O�i1�O̓O��bb)x7ȅ\�y��ΐ��7m�<�q�F��6�~���Rf��p�0�
J@^lj�D�z��8J&�m���$�O"]��*�O,�O��2��B!0*���G�.��f�i�����'-r�'���Os�IW���·'� Ac��\�AS �	FH�7<R2�x���DV����I(#�d�%�� 2��1�׻if��'���S�a|7��O\���O����O��C�s�Zu�Á)N��'�5���'|��'v��)B��?I�s�Tx�aM�'�q0.�t�@q �i?"�D�	�7-�O����O�āx�D�O�a���Ϟ��d�>�4u{2_�܉fey����ӟ(�	ȟ���_��˶Zu��p�ꆕ�\pZDn�	=U���Ոy�R���O����O:1�O��I͟h����'òu����Y���)�K/It��	ןx�IП��I{���'�I�G%r��=ҎޑJ���SR��"'�����[��������՟x��y��'<�|��MKC�S4K ���%N�_b�P@��ۦq��������{���܈G%������T�V*,0W���<�j]�P�>�MK��?y����O�\�A<���$��@� ƬC�� ��Q6M`� ��Ӯ�$�O0�$�O��̦��	ğ��	�?A��ꔟ
���"̔+;���'���M������Ǫ+�;��O�i�|\��#Z}*� c�t�Y��4�?!��u8�� ��?����?��'�?i��[��Ne�8��ir%�}o+Ǧ��Iҟ�s��Ge�b�b?��ծY�xd6�P*��e*gF~�z�vmƦ9��矨�I�?m٨O˧h�B�P��*5 �u���üu�ڠk�i���!F�$�֒O�$	� <#�O/N���:�A�q�� l���I�����(Q_y�W>�I[?�`����䘥I����GtY1O���f��~�S��	ҟ���*�7_���)І��7���� 3��ā^x�����O>�O��B3
���0҂!%rਲ�}rG7��'���'��ǟ��	� �щ�Ȑ�-p��I򇌳^�^�iW�Ӟ��d�O~���O�s���'�6\b�a/\�5H���(	Ҵ ��W0�9�O����OX��?i#��B�!L:NE��P^ :�D�QC�M���?	��������	}��Uy�i��h��Z8Z�lT����#��@�O��D�OL�$�O^����Z9��l�۟��	�vnʍ�u�L�-�[�-77��3�4�?���?)O����V��	�O��ɮ6Z���B˥{j�y�c�/X0f6m�O��D�O~��>dbd1o�ʟh��͟����g^���E�*|����І28���ش�?Q-O4�$qv�ʓ��4���`P�%�P3��h� ����M����?q1!�1�f�'[��'����OG�F�2ⲕ�b�����3�ߌq=�듳?7'��?����?��+�|�K?=RE��`P��S-�~HF`|�D��㌜Ҧu���<���?q���I����7�O�2� �jU)W&nb�B��M+�M36�N��?����?�R���|
M~��'e��0'a˔ J�<*����$�
#�i���'�R�H�T�B6��O~���O�$�O�L��y�S�Q���qs(ܽZi��'.���.E�R�`���)�f���O0E���΃"�yrW�_�������٦���N�t0�4�?���?����o?12	ՉYa�ŋ��R*#C(`�%�Ԧ]����-12��I矠���?��I��p�O$J �iO4-�j pGɑUС��HU+h�6��O��$�O��^��Y����k�	5�nYf���@�iS��s�j��	˟T�I韰��Q�4�w7�L�1Ʉ�I�E�0�ԋ���13�Zil�ퟜ��ϟ�	� �'>�����"`����U�Z[འA�B�v�6M�O���O^���O���K�f�oZٟ��ɚj�<� �O�b��anόs9ft*ش�?9��?a.O��$Ĭ��)�O8�	�T���Kq➄|�����ܧDYH6��O����O���ۻ� 4m�ɟ���П �:'��ٹ���ch���֘k3�,�۴�?�+O������O���|n�5�\(���4F�QC �u��6M�O2�dTev�n쟤��ğ<���?��	�n�Z���F�,x3�\�*�^��O��n� ��OX��|H?�� ��(qn)�qːq�8��vӈ}�e�������	�?�����	ܟ$��J[�@�1O5=���K�_��M� n���?�.O\9��1����鎭=�e
�ݥ8s MW�P]l�l�Ꟑ��ß�1$M���M[��?9���?��Ӻ��Ύ�j�p��!\�uk��������'�Q�t���yʟ��I�OJ��:��j�@�e��{��o�^1m����FM��M���?����?�P_?��3��,(Q��j�.@h��G+�8�'�Z4z�yr N���=wJ��OJ�ݻې$Fh� �/Y�AsL���"O ��jT�nG�� gNμDZΌ���ɷ[�@��䈏t���#D�,u�&�e����ӗ�D�v��Y3�Q5@��p�3k���'@O�;$����7˦��O�B~D��\+|�����i�b���j��w��z��3\z��;� �:��)�'���IWhlc��ϘO���:0��/G�vxS����hTpR�+\	��iU@���A+QD�+��Lb��O��D�Oĩ��I����c�ʧz�`� l���9�\d�GyRe�#I��~`JH>}���a��w�0L�w�P�'�Z ���?1��?�/�v�q&�êS��B�O&�;�#�O�"~ΓTΆ����HR��h���#%tu���ēQv��*�nT�/��)���	>�6�̓h���V�8��z�4ɮ���'�!�,l2$�s^hP�v�=2�k�&�:SL��q��
�YI��y�Ɣ�,s��C7��w!n]ِ��!CV�vhX�c��u���7�Х3��	9K�D�r%/W'3X���:t����+F�M�R��3ޮj[�p0͙41�lh���'��������O�M�5�;� !�����I%"O���P䂒"o��jC*�Z���bቩ�HO�i�ON�W
D(=$�"�L�l�~��A�O��������j�Od��O���OD���'j~U8v�	&ld)V�6aV$�Ap��SW<��gRg��#4�_�����ƍ9���)סP���9K��*�X��m�Ct��"(��T�`�Qҟў��T-�-%:���*N��̱�A˟�Zb��ӟ������<�����ę�Zn��P��l�
��H�4(�!�d�)"�)!�D��0	���K���DzQ?�*On"!.Ѻ[�k#ZG����$y��!��ѝ�?Q��?��dz��Q��?Q�O)zXU��2��g�b�<����5G?���.�B爝P�Ƀ�<%�P�g��Z�'�x��+u�Ƚq��ЬK��p��FϰXר	8�"]�E��i˷L̞-�V��.6��������Or�dW�mX0R�(�A����Ň���=I���֩j
J���nY�w*����Í>�!򄒃���PV�^[��y�E3J������	wyl�~��7��O���|�b*G�Ѻ�� �ǅ zb�)fI�9+��;���?	��*'r����H/?������k�>l�0�@	z�$���+4�B�#�
4L͙�C��(Ozh��o��*^=�6,��$�YgF#���*@�%^d��� ��mj�0�l'��'
h�H�sЛ��j�:���|
���4�)X6W�.(1#
��?)���9O\$3���>�`XT�� j�]����F{�OB�O�}�r,ڍ
��T���VBL�U4Of�	�d�a}��'��� X�p����8�	Q�@a���P�H927�	��b ���
f*�Dp���GR��2�H�f�@��VF�Y���� �a�B����`U���%0�U8�۲��ت����U q�ZsVt���<��������ZQ��ǐo�5яچϬ��a�U�?9��?������i,h�pa�c
�8����y��'��}�D�J٢@��
,Q� �p�π�O�	FzR�OOR�[_th�ȗ�gRH$Ң$έw"�'�V����+A��'e��'VJ�]ӟ���03�q0�<Z�<���͇�17��*3�|.��&���X����%�?5�p��^{1O�DR֠�)M�x�یeO�Ɋ�CN�Uj� ���d`h�X��U5
O�ig���8倖W�I�,ۤ����3�ʹ��_�J�.�	������O�O��d�O�˓@h����Y	��$j�L&��ȓ:?:���E�K��xx���;`a
�P�i>I�Ihyb�ҧ��+1�0��� ��]�Wn�4�2�'��'ɐ�Z��'�:�0�$
��&�r�p��0�(�0��-# �iY'ω	d���x`,<On� ��MW�HH#J��SȚ�kpd���@H�#ʦY�4 BF*7<O�LH��'326i����=D"�;4�ܣ�0�m�P� {�>�I�z�8�+!h�?qd4��d��7d�LC�z�`�m���Y�TB2ez�I���$7��Ħ��I��ė'��C5��OL��g }"�l��Ά�Ro�'f��{��<���ϕy8��j��x�dʧ?�b sǮͺ~���L�%w��Ey2�Q�/̈�jDA&mf���@'�&���5�p��2�RB���&	��~�Ģ<�Oߟؚڴ-
���'��ә+�ƈ�G��&���{&Z�#T����l�'��O�?nO�Lҗb�d1F%8&��@a|�ž>���ؔz�@�#oK��zS�(;�̓>�ʉӦT�(�	̟8���U�d���Ο���}��UٓA�z}CE��0�<I�ʓ�u4�H�"��<, B,�P�T��'�P0�`�}� �塒���Ac���ze��&&8zw��R/������+ŮK䥸ulT�]�T2�AG�.�\���'Q�������<it��T�� ���.F���5��Q�<��H�W���#��N[,tBe	LT��?���i>������,AglX�|h�	���/�|x�Iٟ�4�ÿA���������՟�Yw"�'$~��1��U_�����ƑG?|ҙ'Bd�`Ƣ�������x8�`����9qUm����8A�X�����G��F9v�,�P3%" |�g�'v8�g)S�}#g̘�\u"<{�'��H����?9M>����?	-O��J�$�(h� A�Me|l\x��'�n]9�y�i�\ܘ
N<^0`��U�-za:7�O�O�)�O��͈0�$�iʎ���m�
=`\�×]��y-�?Q���?Y�>�f�{���?�O� �Ш�#w��t�����;���y���
ҸD�"�M�~ɻ3�'�f��Y�9(�d�$\Jt�'�9�$eP��E4L΀��@
{B$10�e����ugB '\�'���:�1]��M^�r�&8����,"��T,����7�O�ʓ�?юʟ�8�D��
Wv	�.{N�!��'�ў�H GԜ�s�������hq�X޴�?�*O����Q���	���OP���#K�\�h��	ԉ4u&y�Č�95��'�R�۟z������G�x�����؉��������8� ���fɰԉF��<A�m+��.s�8`!�̎v�~@E�]3$4�]�:Q�b��%1�i
@H֚:Ԏ��D�M)��'�������?���?�-���I��)yD�Ē j؄3���(vk�O`�"~Γf;d]8�V��3h��xTE�� ��k���:����0H@�Yd�V��l�Γ=��푓�i���'��S��I���ɑM]n��9��%r��N�y8r\AV�5 �h)�?1�D�����z:��&���B�+���Dy"�˄�۾Y����,�V6*�K�Ï�LNP]���F2k��D]w��q��]�W�����2iW9'���&ST!��aEY�.�����O��$�O�#~����^`��O���ځhu@�	ş���	�h��H���y��q���Z�5Tb�x��%�HO�)�O������fM�)�҈�i�����O��	E��E�O����O����պc��?�%�HcB^�3�l_�����D�x�J�x�T't�*��adR�H̠���Q��3��=Y�5�Wl��>t�D�U柮!��t���u�|�x"�̘^	���?G��tZ�L� �I�Z.�upt�_�6�! ���@��ɅG����I��M�����,O����<���̧E�D(�D-� xѸ,��FKD�<9��G/��%��=0��r�������Sȟ�'��A�L�b�b�-"�%��rm8B�?@mr��3�F�V�,��	
B�I6cj-�T�_�G<<ԋ��_=��B�xԦ|IY8uO�H�1�H5>W�B䉷"K�ŊEaBqeܤ�s�ǒm��C�	"~>�IZD��Tgd�F��.gɪC�I5)'�E��j��X�~���&��X�C��N�~����(
̎��6���LC�)� P=�b[&X��'ț^���"OR`�"ŌZ"@c&�*��yz6"O���`H4ydt`J$��K��i1g"O^1y@$^��F��gޔ`!j���"O��3�i�uE�Q:��D�Y��"O8}�uB�.R���F�<.W���g"O�0`�	�p���@��%����"O�P)��f�cb
Nu�4��F"O�(&�݌P�X�K���P�)SA"Ohy �>f�XoJ7�&� "7D��rT�_h�>A�u�Z�x�(�3��6D�������;rAC��j���`�)D��3U�=k=^��J�S���%C&D��:a)?�1��[�dAۑ�%D�83�šD@��.B�B�a��/D���G	��"Q!��ȅLY0��d-D�x��L3F�Bٰ发�<�F�k�)D� ��-K�!T~������p�H��'D����Ć�]o
�؆����0�'D�4ء+S8:�$��L�K�(�4m&D�D�A�	'-���s����MyS)�r?�6�W��0:�h׻
ٔD�E��H�(E��k�^%�L�sj^)s��qbp"Op	0���|��dX��<=fe �� [����'?��Q�kF&R8��L�qO�d��$I<]�$��eE2�v��!�'�Nɒb/�-e}>���_�;"��
Q�_�����!H�����)»!d͓����O+4�,n ���sC�
P��ŮO�'�4�.r����wK�*c�		����h�+ԉx�Ꝫ�+Rm��ZrƟɦ�x��N�=qO?7M�'.����	D8ՙ2CU,W�dρ/@%҄�A�i�T�p�I�n�)�Ӊ;3����FR	F�["l�8��z�b�R؞1�(ΣRp]���Ӭ(��Ū3#Z0�=(�	�<!�~���M��\}vdK�i�t���h�������-�����,����laL-�sb�W���+�k�<:|d����|���{qa^�r?�̡�Ghi\�3�?�P�?Z�h�C��6U��S�2LO4��%FM�j���J a���:Y��nY�r(vQ�2��K�<̳���g�4ijj�Z�'��>7���l$�qÍV�_|t&hH�g\1O|u"`X�'�*i�B�p\h�����R6V�n��I� MT�5Xw�����:	:H�&�Иg-ay��°2�J% �K!o����r.��,)�D"RѾ�"$�.g��z��d�ڻ<0P�$E+
�j��
=���*�oa�P!Rq��.&�M��/��+Y�D�[>���c��8��&d���4��ѭ|V���w/��/ʆy�Ğ�\��!�4 ���O�hHw� 'Q$8�Gx"�>�H�j�5h��%Ӕ�!"Hq�3L�&$��P�� -��!�G��B��Ha�I1��-�ր�3v�D��h��^.~�C�%ϺY�Ҥ�d�38���C��F0���#\���8��BX$�~�A�-ߚ9ҥ��y��,]��˂c8b�n �*�q<��� ��h�v�a���u����d�F�ܘ����ga2�]2*�!j0ƍ�TP�;�&³eE�%��8�ܹ�C�>�'��qb��և J٩'�t�^�R$�
%��Oh|
f�����m�:�q`%�� P/�x�`�"K�#ǢWk	 ��o����h���!êG&+B����rp�8�R@��	�:��r�%��Bz�M����{()$MXx�I+$���OX,���/�T�r����6�ȫOyS�<\,�ڲ�W�%�]���O�J��="��uQ�U���_Pq���-aX=RMJ{(�1� �In�ܬ{���ʟ�82tH��Z���`��D�i��g ��x� 	.vNE������GKO$\�2ؘ7 X�*�j���<4�E�є>������MCT��O"���gG'�IH�"�3)��	1Qm.�|��:5DR�V��HQD��*�F]ɷ#İ%��	�n�>p����!�b B�d߿Pov�'��T����J���(8﬑��ǫG����$�[�p���I�U�<����y_ʅ�B_�lV�dz���C�>�Vb�0x(I�)A�B�>��mVY?�DA�O�x�阼.3�E)�`�?qڐ�D���y� ʕՌ�(wEL"jHd���	�W��]�W�ȫ2��%�����Ӻ�S�T�B�s��j$Л=>��D�&Z�,;�E�� ����#O6��;3#"AB�|�� ����:���27*�`D�5���>�v	ʘ#Ԡ��V   40����%֖B��i�H��I pI� ��F21�Fɸd�
4pAK�!��'I�����j蒶���� W��Y8Q4Y�|�C)J0��ɩbp�����[<
т�j�o��~,�&?�wwTD{a�� ƀ�s��.!�1�I���n��0{sO5�3�T	bd�4c������w�]2�G� �H1�HI>,kj�t��ź��Ok�E9L{����FB\Zݪ3�	��^����-�n"��ōz#��D|Ҩo�� �)KV�ǓTw�HB�KV�|����� ,�I�<v��')��'(:8
�$I1Ee�	3�	ޯ:i�A�ʸG�&�SP�,�rB�y���W��d��6恏Ib�i�F�X�2�=Kpj���D��qJF�'��'4Cg�۸Nt,����R2I�(ϻ0�mP7�^�>m|��u��0*����'w"�k�+��k��P3��&Xw6��}�'h�$���ǂ|PA��ԟ[SV`��'��� �>`%�ݚ�
�.t���J~�'�M��ZmS��-X�h���`")�4X���2M�/Y�Ԋ��D>��<�R�R�N���1���&�l�[��i��Y�ҁ�ҥ���f\l�Y��I���\c\f)�����3�騖�حX{�j�{r�F�}�4�	����?�.W� Kh�� �="^5kuDŰear���FZ�S�$�b�^4iqLՐ%���N�r��P"IR�d���K[�2A�e+��A��e"�ʟ ��R�|����H?7t��a/�/�^�Ip	�>��C�.;9�|{��_�`��h`��|�<�bK�K��򂋊E4��J�O[Y�!����I�n6D �0�
o8��S<Z��ݠW6J!F��No:xaAbQl&�xa��1"d����7V�qO�c?���g �V�p���|(d����O�!"�b�-S�~\�J�~�|����ԟ����)�l��QX�oN_X�L:�	�o���	"��k��I��_$Ky��b�.I�������=N�ً!B�vm�uY��O?������؉%J쟪�⢣\�֔!��5Q��$����n�1O��w��	j��� �\��薤�˼s��wr|y¡lI<]���E�_}��.%����cm��h�9�tH�[��y"�S)AA4=B�D'GQ��A�.q�.�R�Dұ$�ZT2,OĈ�PB@0O�)��A4*�Fѹ��O�}2��y&�<�a�Ű-,��M��|M�c�'X���'�T|1;O�=����N3�6���ST��pG���?1�c�Tt�0��MT�M��k�F	f��5���Ac�D�5C�P�iUd�,�챪�$$�]1 Ż��}�N?)n�J4�w�)_�z��b���85P�O��rA^��â!X�xyu�T?qh�b�4Me��j)���sl�(E�"��>g�,�;��.qG��S&*�!:J�r��W5��R�d�:a��	KxN�λ"vĨG���7YD�N��P!� ϓ:�h�z�M�@lTy

���'@,�y�x���CW�I�uΠt�:2�f%j��Wp���gK�eI:��'���`Vj�h�����\�	����'!���A
����B�8����*��y�h\�/�,�W��/���!JFb?�c� R�누��T;q��H���O �5�Y
pP�Qs!��+� �a��T>A�g�*����@f�J�Ό��\9֜����)m��X�B�ܘ[A̔�O�4�a��wk~%q�NM�oD�X�[(F�Fuӡ�ͦG�|$ȀG�=��`�{*����K[��>�:Q�ČR7|�7A��B�\뇢%!L8!wǏ(PSԸh&�ܳz *pRb��Qy⪈7G�N��(�x%��>2��q�5��*󄂫B��!'�è���>�(��N�.>@���2K��\���!�t�4]�Y(p��ȷ^���0�v�����gWj4�f W�D�.�	�`��K���|P���d�H��	��Ol�f/Ǩf#vXAP�G8�$ۅ�^.6�O�@�Ӧ��$GMR\k��X�Ȥ���?Q�C��f���@_h�ʠ��3h��h�=�O
�р�&Z3�ڌ�`�d�΅+5-8$2�#��(}���B��L�S哚v�t�4�^~2�ѡ>�P嫵-Y'r�ur0h��i#�7E^�S�TcK�d��H?a�s%��?�`Q����dZ��� ��"9���(���C�͸Hp�⟴��{!ǁ�C��=�C��1_V�s0���<9���~4��mEG����|�iM
c�8�y'˙�Sf]`�B_	5��Hӧ�T�]��`9�e�Uy"E�*���L�9ט��SJ݃�����|?m�&p����4)k�ۃ�<3���Q}2!{�ۇ�s2���F
��Nh����O���[(���1䗚(Je�bDY-%�#��[�~����D�nƔ�P��K&踧�闓B8���a܏�l���	2W�9(����F�+��זLޞ!q�� �U����<�N(��PA@h�l���H׈4�f�B�RM�u�=�OP������؛Ih�hT�z��<��..��L�J��2g��W�p�'�*@����\�a�	�w�AX&��P��TJ��'-�Hp9b�t�l��\�d��}І�>�{���c�@[ �%`t���NI%:������ԓ6,�PL�d+#�
�#�X� �.05�(�@o@�r���8��<qgȐ�z�͉Ł�/<�8}���U~�3}r͍Nj� 2+W�����`�
���	P�"�zG)_�o���`��`	
��#B�7�D�������	��8�G�M�1�dǊw8����#<t��z/+��I?Cp���w���'�q �ʂ6ZrEnʛJВ��Į'p+,i��{*��4;�̴���i��5SpN/tV��i�*]�*O�%�gV�]ڔ�O�)�-�T��E�&�xt�Ν�C6�UXt( �n� !F<O�;`�H���҃0�~Z��IFȈ��	\�/���"��"aP��fiX�4o,]&��S�iY�p�,\���9l��,M�%�
sƲ�̙�L�Y
�Ո��/>y�!U
޾]C��I�h��	�y��h�&C�R�')��$�4�ޑ)���W,̀QR�i8tC^¦�96͇�9b��4BZMn�I�{*� |Y��Ѭp��l��놧�\��$�O�J��<ny��ՙK��}[����0t�L���?�����3�D�q�v�����aa�I�J�D�[C����"�Ȭ��k����)I�gX�8��Dהs2�,����I���#�^*�tL;#�ڢ9�M��c�2��4o�?���M���cG�iԢ��	t�a�d��=�SS��	�\�I<϶i���@u���2D��I�t�O��r��O�)��O	!.FQ� �ߘscX 8Հ�ҟ�f�'O��{����6�r��Mˡ'@~c�! ˘W1���$��X��3n�?��@��&�ĊG�8/ ��:;F���gB-HQ���<'o�����'�&Հ-��i0�1v^>��3F��3,�1���#$�e3�?y���_�	& ����N�F�q̐�1�4�� Ri��� :�p�Ysm~F}��/�&jJ��e�T?���nݗ��s�G߼'�сh�~hh�L�p���qR��ᗦ6L�#��l��t�g~rH�=s��J0
�4�`�\&��ۍD#PE-&G�D��D�3��'O�d��'�j|��D��l	��˺d��Y��o J��� ~��I���Uy�����$b\�"�
0�����#�j
&�Хj��'�z9JN�����-���]4-U��XgIY*�I(!bBE��O�(�TJ�h��$>�S�TMPx�B��Ʈ� �������V,P�l��d(@"F,F�h� ��s]�a��l��u�p�O�"%4:�-v�S��d��_��$X��.��ݧx��{g�i���ۤ�����\��!
�7�|!���
x����O�؛+J�r�ތZ3�����)�ztA�'��̪1+ϑ/��V�V5��g?�֤W7�J� f�E�xY����K#�0s����6�Z��o��Pٻ0�g��$�8�<,���ܴv�@�� P�J*������4V��}+�Ub?Q�GO&o��Z�9 �B G�?E��iiyr�<��8�!���������A�cp:vǉ�x�h�:Ó-������%cM|$������ٶ�[4�x0��W?�\�������'���'�$}�!D�Iqdܺ�%LM�tc�'u���^ԡ��Tk���/�=��O�%�OjPXzU��C�����?v@��m�+g�L�:���:�|���'g�P�Uφ� �ԁF��
@�q-n����ADۜ�h�$*��-N@��P�+��u	��'��U�"��F*L�l��{F��a%�O����NH)| V$�D
�p�B��W�xr��r�\%0ea	wj"ɱVL�<~���"��E"�6�r�.�<+E�yB���#�=��؜f Ti�Ȓ��H�9�b��
~��kJ�p,��"t��M�>0��&&H9��C�I&}Q���B)M"}\�;��ܘ}�"e�˓F����sd��q{��.��gs���.�
�e� �δ~����$�8O�1j�	�#\�{E��*/����bJϺF� �2��U�����N�"~nZ
1E&�a3l�!_怜P&
�Oģ?� �ݐ���L�T��5w��$���
_H�12\�ܫW���*}��	E�h����!��A�L� !�C�ɘG�\���߬sh����&A�dC�	�?+���$B� r�x��0��B��<��|9U�+z%��8`�'[xB�I<f��|���B�@y�ѓ/D�C䉢y���X�E��y��ѓ0f���,C��'W;ԅ{�J�9Hv�e�2�ѽ;C䉎'l�۵g�V1��!N�{��B�	�.<tX��űQib����q~C�I'0��<�� �zr�
�whC䉛C����7n�2����	&��C䉤�U�Dg�
R� �P'�L3�xC�	�W��"�a�0<�#��K:�C�I�M��$z� ڭy�5��[ĪC䉨:o0�B�nҒV���8�iI-4>C�I6uh����D��3I��RM��.C䉍9��l`4��,�ف��F1��B�ɀ)��@�ˎO�>y;���
�B�$;^��M�#O��"��9n��C�I�9~x�rMB�if�$��̕!6�C�ɘE	~�i7�Jb/�1�Æ�5�FB�	�$Դ)���1|:.��s*��B�	�vSY9a��g�j	%�]5+�pB�I.�V����ǤI�H����t�VB��2n��0 d��UF�hS��K]8B�ɼ#�~X��M!qO49��"�y�:B䉶lw �A �%,��YE�y�HC�I� x�B�4kM�h��
�	4�B�Ɏ
�H�Y'�M~^�Le�݊RԀB�ɿ]��@@�@ׁTR Uj�c��p�PB�/}T�}�fp�M+�gΔ'nC�ɠ;���r+��%������b�B�ii�a�iZ#GL3el��d"O܍�Eh� xP���Ӎ��+eVm�"O��@�N�Z��5"�΅<�R��"OFP7���Y,�L����7>��p�5"O�,�O�lfX�0,?x��"O� `YP .�	_tr "I%}\
1�d"O����N�c��o+Ó3c�l:W"O"d��N��R͙BE�t���U"O>i�7Ϗ/W��7��=(oF���"O���Ȕ�C��E��ړZR~� %"O�H�f��#ը��F'�!J`�1"O`MY�O�
zb�kG�K�`��"OL�"�:	~ �`����L�JPk�"O��!����=U�8d`ʴ,�9Ӱ"O��pp�P(�:��$@H=��J$"OLus�IҖ@X8���X%r��� "OrqQ5MH%8�N%�ƭ	���L�"O��4M� ?ݤ�A�JX==� QQ"O�L�vAmт(R0�6q�dq�5"O&���2Z�<�"��J��P �"O��R�#�'�6AJ��5/�``b"O�ר��GN~U6�ԣ=��<"e"Ob�H�G�p�8Y"@�N�d�x"O<P�v�QA���2gJ\�՚��"O��rPC�|BP
`(�d���:�"OT`��- 3�R���U<�u�"O,���'J5qEA��(? ��"O��b�d8N6)r!��;\!�"OB{��rQ1���$I3����"OP��4��!D�0U��gE����"O4���'���;�A��p120K4"ORX ௄9���G/ 4p����"O��X �# ?����}���A"Old��Q"�2D�'�\梔��"O6�*�II�A�x8��D�8��8'"Oh�s���7Y��8q�$UPGP!��"O}���F�$#�aW���آ��"ORQ�vCD Pv�E�AC��*�iu"Oj(3�����r%Ѡ�Ǩi|�6�(�S��yReK�QA��!�H�9?a,`��!��y���B ��x`�č�������)�O��䭁9�`X�f��0���B��'�qO ���D�*_�	� ���a�"Op�
%� �ʐ��S�d��y�"OT%�� r������8|C~L��"O����ټv2�H���	�I(�*O4HrLpm:ũ�;%���'������~n� e`�$A�(��'Aā�&��+�|���DN:�x����I�Sؖ�2��(w�����,��R)C�I54"��(�/��8*p�9A�-P!@B�7;0�Zpg	'NP�׆;X.B䉋>�x(���H�,,$tP$�*K�*��G{J~bA�CaZ����H�==� I�	�u�<�"��"j
�`��>`��Hc���n�<�L�=�XT�v��<G�	�s�<�d�CX�t��iJ=7���j�h�<�A0k P=���Լ��l
e��z�<��89�x�H3g�$�!�&�u�<��Eowm�r�R�R��$9Ҩp�<�d��*g{��e��*AJQ� �n�<�tB��>�@��S@�YĤmYg,_q�<��oJ�E�>�	DF�P6���Om�<�D�ӛ/�,�R�%M�*/B��BßT�<�Hϧ�^����ס^W��1ue�T�<�g&S=<n�HxD�Pf@�Y&D�R�<����4>�~��.[�J50��peF�<���G$EL�mO�V��E�4�XW�<����@�)9ҋ�NqBq���n�<� f@)5/F����E���"O����ġ�0؇ˏ	4F�1"O�ݣ6F@/T@7M۲+�hi�"OR(��N�IU��	�,��(D��"O��PƔ���U�&G�=b"O�|	"�O�9�L��\
;�	�5"O�5J���?�@���E(+te{�"O�T��F[cd�XW"C�f&T�K�"Of���%5R����E�����t�"O(qQ�nM����rh���"Ov�+ĴN��h�]5�^�x�"O|@Cȳk���1�ǶF�d�c�"O�����|�I��:.�j�R�"O�Lq�����#V
�`�`%�CO�I�����$�/	�~�	1�W��=2p�ڢ�!�$J
 2�Q�V,� 	����%X�!�,n�8���|Z�L�����!�DI3{���2��y*]"�A@>�!���\E�0"Ť��BEX�x ���7�!�$�&��eQ��S��r'�4@�!�$��1��9b��HU�՘��T20}!�d��I�"�R��	7N�D2�W�	v!�$^�p��኶1J:�M��c��[
!��Qs'|��u�ݑ�,��8
a|r�|�؃|Z��N2&�$���V��y�#�4X�ʇъjTHH7)���y�O)�R,+�B�c�����c�y�������@勖26���ĠR��y2����1�/��59��'��y�7mlx؂�l\�aR�yb��(�y2�X�(Xy#A���#rA��y��'P�HD:D�8{LThɧ+����'�az��9� 	�H�R��4�?�y��Dޒ�`�A�� 9�M��y2���D�Cg\�1ބ�3����yB�.w��9A1U6#x�lH�)N��y���v87/�A3,)"�+L4!�\bp�Q�ޓ|n���:U�!���]��b��_�e��:��߲p�a��O6q@$��G������=���q@"O��	v@��1��Q"Ɖǘ{��x�c"O��1�Ճ!��
F鍆>QJL�w"O0����l=ddqN�w�% "O����Z$%*򌗑X��!�"O>��"FF��<�bR8�����"O���G�M�Ga�����/����"O�	`$��vXr��`@�G���E"OHYC��W2$;�9�� i���IT"O��K�$�SX��g�Z 3��)@"O"�tJ��|*�pk��J�e J=IE"O�$;��J/ʔ����A:M���@"O��i�ςq�r��l%O|�PV"OX���]<Q��X���R�|5�}´"OvxB�/�"$���Uj�"�n$@�"O�YҴa�x�j���fZ�k����"O����5�z������	�@"OBuk��A�����-�sn�H�"O�l!@K�T#>�������ܹ��"OX�2�a¦,�R
�"��}F(b��)lOX�qr퍒��ui��i^<Dy2"O4a7iǽ=k��Kы?l��eQ6"O�L`�ȇ�P6�rщ�.�p��OYH<���0ؾՊ�Gğ{��bgC�B�<��B��Mx�I㥈�"g�5*�E��<� �Pp���}�EG�s|�B"Ot%�g�\�@�$`2AhS/+Z.��b"OXp�&�3 s�u�VDM�J:���1"O�02�ɍ<��ߺ5�q��"OR����@�B�V)XU��AH��Z�"O@�����*ǀ ��9@�|����'��p�q.ۭr<�j�I�>�U�6 1D�ԃb��_�jD��΅�^~x�A��3D��c��Y$4z����PZ��2D�|���X�zՄx��EE�4�N%)D,/D� `���9`ҜSC��MMTx���"D� 2� Y�]fhȀPg�:b$�l�&D�b�Q�;��l�E��!u�ZDЧ (D�Irl�I8�Au"g1
�9$�1D�\�g���b�д��P8�0;�2D�,+�)M�FrD�g�Y�n��i��<D��@Y(X�$sA5]Ò��i.D���0b�Cm|�i�#�bh ��d�+D�� ��܊jܕ[P��������h(D�ܹD��d�6�PT�/�1�]�yb�з�*P`��ֆAL�r�a��yB( �y��x؁��>�TUYq��y��)�C���[���'
Д���Ƀ�a	f��ar\�bÂ�,P?(�E�/x�̓��?�����J��Q��]�JR���E��A�<��e�4���"W��5��)� i�A�<��."]��2dO�����d�<�"̈�#�~�W H^ɢ��v��c�<Y7��b�n=b�_~R��0�b�<��̐'t��է�j����t�<IU�>^б�Λ;b�&�҂*[o�<�U�0�T�"U�ؿ4V���@�n�<�� Y�q�ʄ��JH�8��`���i�<A¬Ш>����D�-��� �e�<9���!�@ +E��lc`l�b�<yRSJм�bbG<ZJt
��i�<��螡#6�H�NһQz�����f�<і$1M>���+�N��5��
M�<��N�)7jJѠ@k�a��FE�<i%�@�P4!tJ�*g&��L@�<��!0� ��*C�T���'��~�<A�
��"�bTi��;f�Y5�V�<1�d�����#)���F`�H�<�#�L�L<�!��?M*���h
H�<�b���n������n�����fE�<�r�'I��0"���2�D4��'wS��ŔQʰ@cLuƶ�K�'H���E77@�J�r�xPC�'K��C*-'��(Īčg�l	�
�'�H=B��^�T�ft{��c�"�j
�'�MhA�mˢ��2���0I�D*
�'�&=A�%�R��0����,k�1

�'7 ��G4%�txy�bJ8'-���'@��A7[k��3+�3owB`��'�#�%�-�1!΂lX�a��'i�Q�E͐�_�z���k,��Q��'7�} ϟ�-J&U�`�D3oz8X�'��$���t�(����
�R���'"0�*��*�>�� ��3`�la�'��pqc�a�Z)�%�]?XJL���'>Q���G�n��H�t�!;�8�K�'�,��	ʼh�6`�DF�.?�����'�4�$'	;��s =�$\��'��)�OY)n��U7�F%���� x<�n	��@L����<�VX@�"O��pm�������)4Cеs�"O�-b�	�1O�TI)���h/(M0"O\����4}%b$@/T#�3�"O����M�4W"%�� e����"O0A��ĕ' ��Q;A'��q���"OIGL!9��uӰƊ�G��p"O����4(��5s�F�-��59�"O�ГЅ��,Ȱx5���^�#�"O��Q􏊓>����cOM�%��T��"Oؑ��N�`�'�߱~�4D@g"O,@�(V^��A�����kS"O��+�L=3�t���	�f�:�"O�Q	�"O$�0l�r%�-Q&�Ї"Ot�LX,eϘ�{Y�1[�䛷"O��#�%�P�q��E-N��"O���«$��3�$�CGZ�"O�0�w�Eh�z�c�c!)`$��"O�0 ���>&pJ'�ɭ?&(c"O���ͩ���3�-��_X���w"Oz���De�0h�^�9U�[�"O��u��.i`M8$�A"|cHL�5"O��q��ĶOH�)���	�@�9"O�TC�M[�]�Ȕ�y�и�G"O$)R� �DD��ԪE��샇"O�j�A��Z��H����h����"OJw�_̼܋S�7�PLY4"O�IjNI>{�ډ	w.Q��jıw"O�m'��.���Ĝ�mԮ!��"OI��/ܠv���Q"	(l�B "4"Ox���
o��*�ڷdϘ@��"Obl(�G�z�i�Pީ�M�e"OxKF<r���R!��C�{Q"ONE�&�Ҙ�� Ο@�Ue"O�=a�+��G@<ʂN�08)8�*"Ox�I�J54V�XvT�S�B	�"Od�HĨ��=fୣ�΁
|0���c"O�-��o�xx&D�Э�90<1��"O���#C�u&�ặ��{Np�U"O����l����y;楏�1!^���"OZ��f���:Ųو!��y}l�t"O64�s��*�D���\$ǜ�[!"O�iz�䘕u���aD������"On�Zdƺ"4����*\��qi�"O�t.W�X<�(#ƽ�� "O@�A%��x����b�4J�6ȋ1"O�5����	��U��.ݞ|Ė�!D"OTL���"(��M�P� 8��hC�"O���d�C =ٜ0��!3W'*���"O� (#��)S��U��E�3}$�h)"O��x��ĞQ�.� �E#i�Lɑ"O�쩥�	�y�\{�(�$�*��"O~��r�Y�+6Pus��)�D��"O��jG��(�8����
6
��8(�"O|����%}L���J�?���"Oz\�� ��H8�%��T�(�Kc"O�lA����u�5����C��#�"O(��c$	*^�NF<h�Ny�"Op�a���Z�0��F g��EZ�"O�L둬ݑb����ٽy�`�q"O����o�:[�����E��_�fp""O�y���{�)Q3�Ϡ ��P�"O�T����% tɓsB� y��"O��iB�H ^��@����S�RX�0"O� pa��̐S�T��рH�~U��#"O��ˣ��u���@��`"���"O��{f�
�bL��/�6{z��"Oz�V'�?7a�Q�F���G۠aD"O>�����4jI�1�T7{���"Or k�,D1G����� �Q��"O���s�Ĉ��u)á��z�
{�"OXq��@ؤ��6�S���)�F"O~�`�̒mf�(AkB k�%p"O� 肫�: �\�`
%� e�"O��!�"�IJ�U����a�1��"Oj��eO��?�`�1 D¬?�r��"O�$�a�@�u�>����ȬjV�[c"O�ܻ��-XG,�H��#I�r "Oȉ[KG�	hЬr�ʓ�2+܉�"Oʜ��,ذezF
�:xT��2"O��a�gĕe����G�R�d�I30"O~���E>J�i�RO��q<��E"O4�!&VLu�4iEnlڜI�"Ot���ƥW��
iJ-c�d�g"O��b����]����	g��Y�"O�,��Ï'r��i���;[����q"O�`+K?dĹ��B�a�U"O:��ަ3��q�D&:�L�AQ"Oy+e�,F�^[���&AO��k�"O`)�V�!s�h$�D��8�̉�"On͒�]S�r�`���4eJ�"O���@��;�$��oL����"O�q�5�ұC����UN�F�=��"O�H�GZ�6�`��P�y��7"OxL�'N�r���Q-�7E\Ƞ�e"O�¶ʁ�=����4+S�:�`�b�"Ox(0�Ǚ�k���a$ń Rw��a"O.���o�E$$�D$ԃWq1y�"Ob]Y��H2 �B	Zv�̺�~���"O�y�voY�w4�1HU%�j�Z� 2"OThHe3p�0�Vd��n3���"OH`( Fqp\p���42&ٲ�"O�IA68>pŻEB��8.`��"O,���,YՈ����	�x��d"O�%QR�͍'pD���59����"Orw��rW�X�rl�հ4�D"O�5��2H��`ꆸ!�~�h"O LJ��}CD�Xs���l��qi�"O�l��cڰq9�zf�Ea��3p"O�lzv+�2 ϔ�Ce��fU4���"O�̈ff�H��مA�VEj(j�"OB�xŅ',�$�$��Z3�Q�"O���1.�(Ir��4�rb"O&h�uD��Ċ�j˖4�9��"O���0I]�J�!JQ"���x�"Ob��NP0KhZ4+k�7�=1�"O�U�hFt詓�GIT���y2d��k�b	spƖ����9�\��y'Do������+�6���ş�y�a�?������$QHؘ#DK��yr%
9v�������bd���yBe̽g�6H��H�ojƙ8n���yRd��x�J�m��5���)äV��y"<�Qz���4�$A�u��6�y���!!�Q:��V:f�Rŭ�y�L�G0LK��ߛ+�E��X��yB�T����1p
E㊁�����y"�vZ���mM-@J����y
� ��2v,�l쮄�`��.�� c"O�x�����s/:P"�=��Qx'"OH��ǭS�L��8�
��A��"O�Ц`ά3tLL���&se�c "O���dT$\^��B�rWTt#�"O��0��+r��C���468`�"O H��F�x]I�
5t�N���"ODY�#o	��N��f�PE�"O�lPe׃i��Q!���4�<U�q"O���$-5 �iw$�� ��r3"O�(�P�ͭn�<�A��:Q긡�"O��:s�ϰ�5Z5��b��`"O��Ҷ���X Sg��{�FQ��"O��e��#���Kq蓶M�HM��"Ol��͆�BcBhŹN|tS6"O�$C��U����W���	0"O�D����r3j$��W'��mc�"O� 9r��?=�����jyw2=�U"O*�S��p�<�)iB�ky����"O��Ԡ	G��0N�8uu��Bu"Or	��.�<8�h�CS*Zf����"Oj�� ��c�-
��7J�s�"O(��F�M^� ������$Ʉ��"O��[��~U�dJ��(e���T"O4y1T
�2�6tC�S#c����R"O�}�rْc�y#�nE+84~}�"Op��A��^(�&��s�n��"O���‐�dҀ�B�%��V��Q�%"OHEa���!8��Q`�J�[��!*�"O01��Y�^x��$�'E�<!I"O�\���y>"�����92c`MI�"O�!����+�8���[0WS�ŋq"O\�*T�_�x�Y�H)�,;s"O��.���c&��+j�q�U"O&]#c�β�؁:��i�E"OQi��ؗ Z��sU��"O��@��<�m՛x�,J"O%iP��pS���+\�(�:}Sw"Od���L�oYv|2�)��@�"02�"O2%b�n�^��b#K�u�r���"O,=�`�J�(jl�`1阱2��%�v"O> {�J�
:�n̛e9�N��s"Ot$k��U�n~�i:a��deғ"O��)��w�	� �2a�"OdI�R'�(Mn�����-(a��T"O� "�@ƾG���GWYP�@�"OJ��qk�#��|�'g�^J&��a"O�-,]@���M�9�z��@k��y�	��>��$�]�� Q��ߪ�y2L�,�Ҡ�QcK�S��� (��y��I`��P#E�C+Q�`������y���
@�ek��Dw�	�w�dE�ȓ�d�z�C��/	��y���q����E�ڤ����E�t;%޴`�DT�ȓ)C Ɂ��8\��&J^�;:���ȓBb�i0� %.%�
K�G��!�ȓ,�
��$��Wb�Ѥ�N PBD ��X&�`3�A`ज�/ٚ.�>1����1/�0��(ye��p���F���E`�� �F� ��!�E�2D���g��KX�ؠ�	?W�����1D��'��I�P�慙K�̵�4�5D��!�
h@,��N֨n��a�.4D�h����>i�hj%��Zl�"U�2D�� %Zg\w�(X1�"
�2�Z�Q"O�4J���fM��`H��@@"Ob�[���65N�g��)3Ą� "O�q�S��q���ЅF=d>:�2s"O:��r&\�lz6���$	�c"Oj��eY�4�d��۾0�X�P�"O�lk�H�g+� SƀآMs|���"Ox�p�% �P��a2gk>���"Ot���H٪)�4c0U6UA��t"O
E�@�/����ui�c���"O>U��ֻq��x���<t|���"O�4*B��64G<b�'��z�b"O�T��T�R��b ��|���!C"O�����V�a�/�%&p�đ�"O��R�
��6 !b.KCs�q��"O�E�A��g}���K@��Z�"OriS�ϝ�;�(T� ʛ�eZ.A��"O�$�@ 
�9J��c�8Z���f"O���G�
�`�⬡��=?K>�`�"OB����!	�ԍRq��� +�컰"O���L�j��q��I�ȝy�"O`mӴ#�~���nҍ5��
�"O���J@)p�"��2Yo�2`["O����	�|���.L�p��	 `"O�Ɋ���?�Z�8P��75�$�"O*a��(YT����a�x1"O�� nٺU� ��C&�+v2���"Ozx��/��<(�)�ę(���"O���!c�*-���[�$��"O1�3lߞ2��@B�v��ɂ"O@�#aW���@�ɔu�k�"O"� ��� �8��``��#jx�"OD�uA��	�����OZ�Z�V��"O�]����+.<�A� ᖣ��B�"O8ФʉP�d�&酎J��IAA"OxI�
	0e�i⑈�!��Zt"O����*Bz��е��	:�R�"OؠXǮ¹9<��*���{�0xk�"O���hʇ+���e���p��U��"OIR��v#�����38�f`��"O���ц���`��A�ٗ/~L�Y�"O
����¿^��i0�O�hu��a�"OP��B�W~h�Q��N�YZH9�"O�h�BG�_Ji�Dנ/0��"O��k�U� Z����<~ F��"O&��#�4���v쐁�v"O�u�A;'L R@ɒ�|p|1(�"O��@/7����ҭ�0��*�"Olݨ��iżHr㗒.�J(�Q"O��u@?U�,��0��?A ��"OL�IP#�HǨ�cR��8
� �"O*�j�nK>4�ݹ����M�xT"O����X�$���"�	�5�~@�"O����\)�����j�i��"O<"g�D�jҞ�.ӄg�H§"O��ڇ��fv� #��$�<�;�"OL�s�JGp���q�b>=��:d"O����X>�Ub�?��l�"OJI�mоyg2m�a�*Q��̓�"O�t����%i��,	��͘{ڴ�`"O�|2� R�MJ%kOѩ
��Y�"O��`bh��\+�!A� 4A�L�("O^I:�-�(|�&� �7�Xɚ�'2q�aE�Xz 8+&`��R��m���� �)��FoJ��i��V���: "O���d�Y�:Hlh�(�'w@-Kp"O�H�@��!:��bU��x� X "O��$��H�8S������"ObXI���%p���&E܀N�Г#"O���3J^w�DTC[�jZ���!"O~��wB� W�=J��N�5�zpk�"Oļ�G	����!�օ1�Z��"O��p��Y�V<����n=�Y��"O��'�Yf��'��R+(=Zv"Ox芗K�(��h��	��M��43�"O��T�@�,��|���_o�:ԪV"O&0wMB�w[ʈ���R�.�d"O��e��y�Jԛ%H�+�B� s"O���'�PX 05-�5�|P1�"O�񵦇5f�j�,�X�bY:&"O6XR���1sj��_�dQ��2�"OP�+"J�V�,�)�e�} �R�"OUS��\�y�>����\�^^���"O��0��fZ�L���ı4�� 5"O0�f��P5
��.2�F@��"Oڔ�"o�
+i�m)��\
V��5J�"O������+4�q�E�L�TR���"O�A��
5M���Eȝ6�0h"Oxܙ��F�j|�s�I�|���W"Or�F�6�4�Q��D��ڔ"O��vDٲ>�����uC��g�!D����."r���E�f\��$ D�઄�)o������]�y�b9D�� 3E��S������֜
V>�*ǌ6D��:_�{%���&�T�h�lD�D�4D��H:�T<������c(D�x!�Ǒi应�B�Bn�̡��*D��� ^0HyFS� ˓F� ��1�<D�K�?'`	F�|3��Rj5D��@�&[$e"]K(�O5�)��
/D��sAj߽r�(�Ȧ�?�p�0SA-D�Jo#2��iХ��hb���v�&D��s�o��HAc��R��8ӫ$D�Ԋ���9r^��B �d �a��#D�؋׊U	s�Pj'nš YƝ��,.D�@��m�4Y��k��D�
E��d�?D��9���w+�����.N0�(���9D����Nt��ݚ�J����Je�9D��a	�%��*�*��d��D��$D�pp����|{̘�@kT5��0�.D��)�nɓri
���#�R[ ��i+D�tp�$�.1M�=(d	A�~9m���)D�4����d�2�3E��*J�]�$D�(3��Ə 94�� �z�1j!D��K�B?e�4b`ۼ9b�z��?D�|ۢ��>a��)�	���$Kb�<D�L�`�"P�� k��>6�$��5�&D��{�@
�� r�!�����W%#D�ċa�(�d9�2Z�hL�ť5D��H�&�:��0�yʅA.D� B��� Jq�!f�<@�̩��M+D� �"P�Z�P��r���1�}�&D����Y�24lXH��іea.%�,%D�4��ڈ��u�T�'����$D�����U#c�65��O�(�h-÷
7D�p6�P��Zb,`��6D� ��\x���s��b�-���5D�dc�ݖoX�l��ۂ f� �`�1D�� �!�VI!f��Y�&�V<o���B"O�C�-p  3��Jfpa��"O1Aw�2&�24�M�IGpp��"O��k��M�t��]��ϗS�@'"O�L0���9��pG�D:S"O���a..�B�SGK�h��(�q"O|)���^* O�1ǣ_�q.t�q�"O��	E�@�01�8����+N<�c6"O���� ��jbJ�#bF�)<pȋ�"O�IhP� ���9� ����=2"O�4�� �j�"�p� ۲h(UQ "O�}���[.Ȝ���)Hkv"O4UI2m��*nx�Y�/�c�f���"O�٧l�'C:���S�6N�4sv"O\���@׳N֎d�L�aÈ��"Of�a�/�1��tE�C�*��I�&"O�p��-_oj&�`)��@+�"O0u�S-�ب��g+yT���"O�T��b��I�THJ��E7}��s"O�Ie�E�!�~$�5�%1��i "Of�b���G���C��/���"O�}�s�"�Te�w���k��,�!"O���f�/-pj��gGA�6��"O��H����u;p��P�O"�jI��"O��5N@(F�D�h�*�0u��1��"O��#u��=;��<h���m����"Ora�mܴ_���T�W8T�j�!�"OP���ƃ�RXX�d��Sx@IBB"O�M���3�6K2呥9���"Oȱ���Q_��ӱc=/��@�"O����#T	,N���Z����G"O hXb�/\��<yS�=Tx�̃�"Oj��q��a��0�t�߄{�Q0�"Oz��Ǌ ea���apfR�Ja"Ot�� F��
N�T�`�?Q��E8"O0(�P��p�iÍO|�.��$"O��`�F.v��`�����"O|G��|҈�v�^�)��A��"OE"̃�&Æ(�.}��)b"OL�+��2�Ҹ�2LS8:UI�"O(����3A��p�,ٰ^V�)�"O�Ȩuȑ�?U��!T�Z,K^�@{�"O0m���i����ȍ!]�$!"O���cA���ä,c��P�"O.�����Ԇ(e�ih&iCG�!��	Y6|�S#��:;�6���C�$�!�dԇ:�v|y� ��6�雵&�(�!�� &}�rDR��&��%�H:Y�!�Ğ4�Zx��j�?d1����CP��!��:]�X�,��L&����N�o�!�D
:��@Q�V�\�8Y��B�B�!��S�uV��ࢂ��.�j5ʵL�p!�ԧ���F+�d�J� ����!�$[l�����[3{��`�s �%(?!�ůp�&��CF�*�<�Ⲏ�/!�d��Q�`-�q�P8��1�c��?'!�$�W�M{���\�P�M8�!��ZAZ��I�F�uL��ū3�!�/8g-K�MG8M���8��1]!�Dq�j<�&-�����v+A)e!�dP9*u��ZƏ?���Ӷ	^>{!�d�H��b�fS(TDL �B�we!��W=4�~@I�H֣Bf������xv!�=~&2I����,)BQ����;a!�� ��
bFہS�Z�@�;OH	�b"ŌQ���As )��o�T9�s�"O� ��X+�Ο!��`�p"O�� &�0{�QK��s{VA)�"O�=�g$-*��Dc�eK�l���#"Oկ}3�q���(kd�:�"OT���
T ���.�
V-p0��"OХڰ�Ydth����<XЁ0"Ox��ӄ�m`(B�ê��ڧ"O�`4 �uXV�r�ޚn!���2"O�%2�ͻ EF=�%�3nju2#"O��'���F{ltra��.\�"O�P�6
�7}]�l�"`�5?�y��"Ol���@�HƜ̃�IŎ&�5{"O�(1RC� ؼ��h��x�r�k�"O�:����fH`�<A��aҲiJ��y�O�x��d
,ȸ8�0�+��ʷ�yB�Q�1�,��ҥΟ.!�LC6�.�y���&WVmS�ߖO�����"�y㞓#!Dh���CH�U Ф ��yRe�?.2���s�$Li�Q�/P�y��#P�,��͙zw��b��	�ybI]�v7(�q ��8n�EB���y�@й6�2M�#ω`2�)5�+�y��N�1�@%+�M��Kv�G吗�y���@n�I���#{��q�oYI�<Aq���N�|�	�O4-���� Öm�<��,R"5Yn`���y�]�潐�ȓ& D8b�Ú$(�cq�J"Tq��b�\���& <,,��j��b���v�x�$`�)���sɗv�<��q���(��A���
t"�_�N���~�݋�����}RY&8x,�ȓ{9�I�5&P�z��U��F�>~��ȓm�B1�sȁ�JdD��q�����r�~��a�Ȩ��#��Yw�<��Ҫ��ЎN�66x�SpB�h���ȓr:��� ��0��[���>���ȓ-��`q�X�l�0@�7a$c�
��q3v����_�9�@�+�ǃ	{����6�Fy��
��{��;@�4�L�ȓ�6��r$�M8>�z�C�+�8y�ȓo��K��Z{Qq����x[l͆ȓH�Hi��3%p,q���~׶D�ȓ.LJ��){XՠV,�*i��~A�3(�h@���&DJ !�L�ȓ �24�q,K Y�B<@��!BD��c=�����1���@2�V%��`�ȓQ����み`�j\��k���9��B�RA��dJ�(}e�beX�o�����)�Q��� ���'�;e�����V*�@{���1t��h!���D�FĄȓ j����	�g���s�jպr�4�ȓ��)B&K4~+dL�DL:yv�ن�}*�Mx$�/}N)%N��]�P�ȓg���!�O8b�jx#�͝�S0@��~�L�x�.ơ[r��[5�Ƅ"��e�ȓ"fl���n��H*D�:qf B�*I��2a�x�%�%D���Q���U�ๅȓj�lԻWKå.�zU �;3t��ȓ_����K��LrJ]@���7,�V��ȓj4ZqI�h:>��"Sh�|-��?�\�7��v�$aJ�h2S�z@���:b���'3����Ԍٰ:k�<��S�? ��cB��9K�ʩ#�Ǟ%F��y��"O0�r�żB�웦�ޖN��X96"OjxrĨٷ$`�uX��/��5	�"O��ۦ�ҧkRP�k0O�59Ta��"O$��rCm8�����xR�A�"O,`QqhC*D���Ή6���ʵ"O!bы�#��܁w���,�\�E"Oڹb4��"yF�"c�T�.θq	5"O�|[s�V��<�ǇQ�Ca"O�X2уџn&E��G�{.DK@"OJ��JG.�V����[ݠ�"ONp� �VY��ѵ!�42>N4J�"O䍂5`��ڀ��!�n7"Y� "O:��#�Nj��R'�D�z/z��1"O�0A�%%I���,�:+�b"OHyZ��\�\h��T�.>!�p"O���6IB�8
n���#��9��Q�"O,qBV�A
:#�W�F)r �F"On�ZN�	|)����+"%9�"O<���E�s��j�3��i�`"OPX��܄W�EK'�:qV�e"O �PT�� =f���ڡ_�����"O,rG)�{zL�qW��(��y�w"O��B�%_�~�u�VcǈG�V�Yq"O�Yy��D�,��5 ���7�����"O2	ړ�&�n$r��Ji�ዷ"O�$�'�N">a(t�Ae�5�"O����C�36vؒ&��Rr��F"O���텵hZ�2���S��d�"O���NZ��H�vk����(Q"O��(�Y&@bZ\�EJþW�y��"O�\1I�wQ~����ǃEV4�3"OTP�E�ܖ��0G�1Bt�:�"Oj��P�=��%puaYc��ò"O&t��
Ynj!��oЂt���K"O�y�HG|� Q�_�i�"O�X�U�ԑ {NP����9� �"O����N9LJ��-B�Ȥ�s"O:-��˝]d��H��,���7"O^q�@�u�rq��$H&t�"O�ܱHإ��%aG�RF�Tل"Ole+dj��G����z-Ba�"OX,H�d�7{axa��e�R�815"OT)��	-c��xGJщ[�9�"O�M�P�';M@h�8 n�[ "OJx��d��(�L�*��6���"O@���/��ku�5�H˂x��pH�"O��*�n��#A�9��gY<zۚ��"O���ϖ��'U& ���(�"O~��a��.m�$��Xvo��S"Ot�
fDI	Q�20�A�Px���"O��w텔]kt�#�?7�5+�"O��5�2V� ���F�l"�Q��"O�\�U���Ĕ�2�O�}�Es"O�$j�bR�0]4|8�C��jg��"O\�� LE<+K�CD�,(�l�"O�����-p�v�����o���S"O�h��l��L
����&�,x�d�R"O��(J��rM�HC�EӁ7���3"O�M���iZKҵm� ��"O���H��Z���ř�jW|$��"O�Cϖ��y`���?Qy�"O��)�!�9q�Qw�Ғyh��{2"O<�P'�V�,����j�5Zo�!�"O� ԙ��+��I�$CN6,P���q"Ob X�`ր2��(�Sa��I,��"O<��(ھY��HD��ElQx"OPi��#�q�� xe��΄H"O^ h�B��m����g
Ƥ�*-�"O6�I�h�/Tn�Ps.�2;�`�K%"O�ܰ�ǔ�JL�!N�7���"O����銜KpɃ
7A��h�"O�)��� y�@��k�v��D@"O�q�Q�ԟ	���P,�mnJ`��"OrdJ҉��r�l�� �>ˆ@�!"OnJ�I�]��C/ʕ� ��"OE��J"M��=��n�1'�"���"O��(�>k�͉�o�'��L9U"O��T�[�?�JaJc@%Dt�#"OBq#�b�.�Bg.���8B"O ��� �$Z��2%��j�y�"O(�#v�r��m�3��8}����P"O���a!�&P���Q
��[M�5"O"x#�GQpH���)�(c[�X�"Oΰ��'��upq��]�-j@�"O`U�@H�}}�,*`	J�%��L[�"O���	Ȁ0)�,�ԇ�&o~�;�"O8��#��*X7�x r�ٚ2]�@1�"O ��(O	<R��D
�sL��Z�"OhmE���D@ʈ ��84�]Ё"OV[`f�Nq��%撡z9P="�"O<�CNQ���ȥ� ��e;�"O$�� ��j��ALj6lRc"O�����\�1#R\Ӥ�٣V,��Z�"O:���Ł+m��K� �<���"O�)G��+4�	{��	iM�� �"Oޕ���ީ]��12�3`���"ON��Voݩ �*M��*Ҧ*-�؊�"OH��`K��4��	QOP�7*�u�"OJH���;/�)	U�	�
l\���"OXɣ3'��:��Y(�5';�	[r"OHr��#]�h�2!���.vĪ4"O��`TgA�RY�r�$m���4"O�6� T�bӍ��"Od� ��5f���H4��6Jh� "O�D`�aO�A� �'-�X�*,��"O�t8�AQ�.�x��f������s"OT���
� ��p2��'�`�4"O��$<ݎ�"��9���"O�p"�BO-Sb�嫳�X�qly��"O��q��\�U�F�i����5��1�7"O��ӇGu�P�ð�s�vQ��"O�"�_�R�H+�(����"O��'�"� �����&"O���2@C\�$%�s�|�e"O��Z"H�Q�f5[��Êv��ّ�"O��i�мsE���R���3�>�f"O��;j�5md�6�R?I���K"OZIx'�D�����L]y{*�@"O�D�� e߂T1%�K�3Qpu!�"O�lS�=������J&y���ӷ"O����X(L�zx�5n��FK�="O^Y�A蘳PF�p�rgW�c-.�KV"O�9	ѪB�Nm���F���j�6�)4"O6��'��
�5ش`^b�]�v"O���6�:��ڒ �$���"O��Z �S-Z�8�A@a�&U~�,�f"O�qRrC\5^��x�����D�D"O� �	R�h�z��9ٱ!z�)'"OX���X��4Ѳ�D)co8��s"Oz�*�M��_]�)��Y4\�q�"O�%uO]�&)�t��9�FTɕL6D�XHDf_$9���#��T��-�$ D�|2B�N�Bqk1oX=_��(��L:D�80G��2O�#��Ղ+b�|��e7D��"��>�4�U,	S���dl:D�x2f)��%�e�C��:}o4���9D�tQ���8
�4L{$d�5H��z1�8D�t�(Ӧsն�)J#6�ШC`8D���EYlr��@]�0�~��d:D��B�+y�H�Ҭ��x�4�%D� ��Ϳ^i^E��ֶS�PD�Vm&D��p��74]H��kTiaƈ"D���&=U�ȑAI��VTެc��-D���ՠZ	+8��E�1u�Լk�&D������(.J�%l�|Er��� D�|�gf
2s��Ϫ�<A��?D�����G�s�ҭ��Уa�l�ʦ�"D��ɉ�H��`��Z�x��`�!D����IJ�s��؁a�̓q�U��(2D����"^1[��\C��G(f���@�,$D�|�QG�30maI�oA�4/",v�-D�Xfd9�($�#�^q�a��7D��Y��?�MZ#ޯ5f�i��""D��
�@Q
a���`������r�F$D�0�E�G�W�x�aG����; �"D���cHI�O�Bd�
�#��hq�h D�Th0��;�ԑ��&}�Y0�
֪�yR,7���+!����6�Z��y2U�V����4�`!���y�e�%��I&��=mw��I���yn��Ex��E��`��y�ԽOH\�C��&&�����y��Ν �`-q�(5�(�0���y��g� ɂ��U��yӁe�-�y2-4����^�c���JA���yG�%�B��g�[8n-��� !P��y��*,�
P�����i) !������yr�H��iY��&�j��T��y"@ܖs�L�Z1�v]x��_�yBc��sV���I��F��SLU%�yR�ǌ"�Z	Bf��$�� qÏ�3�y2��$R�}�3$�3��i� �(�y�#R�`K�ʅJH��)��T�yB/lJ�L%Ջ��)D���yb%ßSb�IA!N�0�~�@�H��y��ϒ8�(���)��d�@@�*��y�.$0��!�DOґ��쒑�y�	��� `㙥%w�H����y��˘�2HBw�� �ʘ�D���yr�&5���p�EǻjD��bQ��y�Bc��k%�5b��9oV:�Py2�
.qO���ćM+",xQ���q�<�e���{-��1J��^��T�i^m�<!��S 6����,��c"n���/Ch�<Q�,+J��H��'m��:�)�g�<Ia�C�F|��ɢ1m������`�<i 
�h��(�m� @J�x2ǃ�_�<I�fk��̡q�V�F�tǀZ�<q�d�C� HW�[v��ĉTS�<֨Ǝwm�����A��m	J�<�@(��Y:]@�(��H}r�K1$�E�<� �9)PO�/A�pcAy�ԍ1D"O&�Y�O��i���ɸ�R"O"Ms�ٜ2Z첔�]#C��\�"O�0���6�� �F�Zu�"O���d�Y����N�1��9��"O�X�2F9Y��@��>*��I��"O
1P��ёF�pX�e͈g`���1"Ox\�BDO�__�th��е	ZhZ�"Or�hq�ͩdA@9�R��2�f"O�ɠ��S�x�01�Ħ'�:���"O�=�`�_�#% �*�j�"O�Z!a�4�(�P����i���#"OX|ؑ偰\�`�A��Y�*"�"O6=2���{��Ѩ 7k�.�B"Oz-r�4[�9��W�Yrb��"O�I!��ف�Zy0'� �+�J�sR"O|�Ѓ��!Ѧ��Z�J5H'"Oڡ�Gd#/Z��J�C�w�HmB�"O�i%ԅc1�����-�V�"O~�"�K,�`�'C�$h���[�"O�`cE�4�Pb��
2_IL�z�"O����=t2�e����<��l�d"O(93��5.Z�)1��
�D娷"O4��q�&KO�=���̶_opy�'"O�XQT��?���re�02Z�X�"O\|:���|b$x�!d�j:�#"O��zD���N��p��62���e"Oȹ��+Ah�ź��T#�X83"O�E� �'�Zt΁!`vA3"Ot ��.B�e����-يb�͊�"OD�x����8���A��8^A��2w"O�ݓ�C��e����d�2#rU�"O\$	��h}Ȉx�A@�)CT�S�"O,��Ȅ�X@�iR᝼55>,a�"O�r@e2D����2�PJ&��
u"O�H�P�  wΒ,(f�ơm8�
�"OT���J3�HDNX���"O�-˰ S�~`\��tO��S�f���"O���]�C��y�`�Y�2t1�"O�\p�?-��tA���8?���!�"O��!壄�b���6L�z,ȶ"O�ew��#K4�E��/C���D�"O��2���a;�ASBoW� ���R"O
� �N��I�7��t�X	Ip"Ob���Ш 4�q�K?O9��"O����:̠��0��L���"OP4K�IP �D�8���"O��[�H�
h��VI��S@���"O,1thY9BxP���o�:�Q�"O�<�n��,1Xe�0Z�D���"O��Qj�A���k�%E�3�:(Bp"O Ӡ&��n��Ka��3����6"OB=A&��/-9֥
u�	'�� I""O��A�a��85���H�|/&<i"ON����f�Q���6���R�"O�<��'Z��e�S�]j7<�.�y�"T;8%��A��91	�Y2��!�yR��&�\��#�,�Α�6�M!�yB��0K����1@���-�Em@�y�a�?i���*��]4|b���L�:�y��A�dIB�6,ϕ{��Ѐ�oB��y�)�b��ҳ	�d�⁲S�yr��V�4P�eL�X$��c���yr�<	К�*�Ƅ�P:�TZU@��y
� ԰R��K<P���I��f]
d"O���f�8<rp�k�����g"O�q�"W)aZ-�t�Dj )8�"O �CأI���-˰yc���"O��j��}�)%K��i�:�Z"OB7_�.X�하I4>e-D�(A �$m=�`"bX�HT(��?D�p� �H�cw��8�葾H)���G+D�$s� .u�%�`Z�?ΰ��'D�(
rF��= VeX	w����4i!D������y�6���&A*q�ë?D�, �݌.g�����ݾO���am"D�XAb�ߟa������n68�>D���Gl���(�*ժl^e�@=D��7��DaAS�Z�f���;D�T@T���(�T c�+��DX�q+��?D�����V�4*Q���CNRQ��m8D��iu��.�~)r�DP�Mㄴa�a8D����!� $���a����N�n�qTm;D� �s��l��k�	j�`0��&D�\�5A�-����T�ԗNd�B:D�LbDOD�s��ACT)F��y��;D��P�@�fh�0����ȂCC'D��aBK�<�vx�Q Z9/b�1�3D�ĉueG�O�48GY�z?B剔,0D��҂,��Z:��@\#f�6�Ɇ-D�l ���MٍQ_�Y�0D��1�����4�ʗm�tPV%;D����!��T�"��s��S�nԛ��8D��Y������)t�� /����8D��mI�pkH	k!o�#Z�*x�נ3D�L�C(�`h�qc.&pʗ&0D�X�� �'t���υ"��{c-D��!�q��ru7i<�ut� D�PA����!��C�����t�!�I����fQ�A�4|0�BH.�!���&/���CA�#H�D���Z��!�P*0�����Γp�fTAwL'_Q!�䞿MT�r�e�<f��XDI�2B�!�<R��l�cD�b��rVHS�l�!��S�7,�s�.4W�
���%��?�!��N Hq����QɎ`�C��Nm!�DBJ�f���ɾwۺU��c� ue!�^���
v�1���%�̜NW!�d�Hg��z�L�e~V��B�27C!�ƘE�~��1/��ooX��!̑I3!��58�l��d�hlܹdN-D!��\�\ٛC�ñE�����-O!�A��Jl��D]!H��xQ!k�2[U!��>R,-�c��k?��I&
�8!�DX�W����	�86�%�t	%!�d��I�왿_+�%����,!�-
v��冈�
�x�f�<&!���g`����A�  �8Q�d&�"f�!�Ă'�8Ej�
�5�BYr`�T>Cw!���6c4L*үx�Nui�N�Q\!�Ą(u�ty; c�&
����-#*!�dY,�*��԰�?(݋`�-	7!�[cl5SKB�A��H�`l�*_�!�d��������6�s�kX�9V!�6	܄,�rB��H!��j��yB!�ʥ �`IPT�΃|�v����/!�dɷO��E+��$@X����9 G!�+"�p����x���{@.P�0>!�� H�ŭP���$q�2���"O��+�΍F#uD眕	�ҩC�"O&4�D'k�����7LŪ�`�"Oʴ"��ˇ=̸`@��8�p��"Ov�:��,�1�gM״$��$�q"OpH��a��Z#��{���1	�'Ǿ�X&�^9>Z>�i�P&�1��'O�}0I:���A�6�L�
�'q��w ��}p��LV�	�'���eͅ!�E�֍�h~5��'�N�����o!b��*� 9:��	�'N�Љ���V����`C>XS
�'����B�x	�$��1Mb�	�'$e;d�|�
��@A�v����'.V�j�a�07����-��?�Όr�'0d�  jQ��h@:VvY"�'��D�C�� A ��'��?%9��+�'�����|���"��Y��u��'��I�u	T�Q�x�v���vU�e��'�$I
FD��2n���f	,��� �'�^�)L�9B��;� 5d��
�'�` ځw�*�
��Ջ0;�h{�'kf��a��2ь@i�@X�U���	�'2s�%�93��P&��3&x���'��h�!fٺb-�mB(� ��T��'��͛���6Wծ�zEԬf�1*	�'ٌtbC+F�8�4�х�[�e�'�b��3(��4T� Z^�L�9�'����l
UO ��#.)ظ�j
�'>�ysB<(M��8E��(�pH�',$ɰ�!�b�"U�7�RtR�'�t�C�-GN�
y�͛�^��'z���*�x�H=�0n������'K�c�A�1h<u(W�O�}g�T{
�'��<��K��Z�T{F�R�{��\Z
�'Ƭ3���n�-	1I��s�L�!
�'��H�#�-ͥ��e�ys�WM�<�����j��
K(/��r`�L�<!�'	�ʎ�h���@�j��'$�c�<9B�Ύ{*؄��2'l�ڵΒa�<�͝0��J#�F�cvYr�,�`�<�E�F�!�\�s��O2!���jKXY�<I��K�\�ʕ�ԫ�o	r��@�<ɒ��!n:F䚇�5�
��F���d^��Z�nX%,h �'�!T��OX���ƈ���Ô�H?h$S
�'38�x����4�2��De�j�$�	�'��8W$�<m���c�`r�u�	�'�H�v�6;�����R�@X�(O����ՊBC�8�
Θ��
S�ѽr��}����ؑ�ֳV���k�OVHC0	H�!#D��P񋖃tu�ȶ��<~�T�B) D�$!��[ǸYh�Bҹ6���?D���S���q82ܫPƑ�h�̰�-=�OV��� qR�Y1j*T�D�8��be�8'˻>� %zl@�ȓD�p���$R��O�Co����|��	�o�j0h�2�eӰ���y��',"=�~0�Ӛ9���+G���;u�L�@��{�'�ў�6/�4�e�ļ�$j�ꍧ��l�ȓKYj�1Dk�=\�l��5(����Ɠ*+�8��lM�D�
ɂ֨�8Z�ě�'M����+�Q7���d#�3E�Z\��O�x�Ń 0��4J@閈#�Hв��"b�?� �$Q��nB���(	 ?̸	�e��R&�7�S�Ov�=�2�,08G�ډ�IB
ӓ��'�J]��f��� ��ʋ��4�I����!k6�5"��W�f(DT��M��B�I�MO�!�Vi�:�걠��%c\t��ĵ>�ℋ��>q��d�'�M3���b�<�bC(G*u��'��D�D�2��^�<Q�A�\@��xQG_"=�� Q��X��w��p��F���H�YU��8 p
���y�B��j,�캅/UxK��z�.�g�'�azB�'�@1Q�׎W���i�նvxfؚ��!�4.P�9����F*T;t*u��h�'w���������T|����'N0���[36r��%��v�����'h�3&�դ_ͨD���F�7j�qy�'#��Df�4��i��R��TՓ�'���4�	�w�qÌ��p1����xr�REnf�R1o
&x� !�K���y�d�'��cS�F�4<�2��yrAP�B�� *ʑ΀���'���y򦑻���ւVB����`�ޅ�yEԋYޚ�`L� 5[
� ��X�yBK n`�Z���'�hR�a���=��?��=A��[h��[��X�W�@�#A�U�<q�	��+Y���JU�Ʋ��ӁAP��hO�O���xC��,`l�x@a̭���	�'*���� ٚnv( ;U�։�T���'侘s�R�]�$
�n�*-�T��'�B��jN�8��4`��E�N�ȝ
�'Y�`�$�ұ/v�T���,F�P$��(O�B�f�GIz)Aϗ�Q�(-�כ�`��	>C9�}�"y�0KC�ͻ	���֢<E�"�&:,y{3��>+�` J7��=��y�#�4qH5R����E�~��B�� �y�|X�b>�9-�y��٫%�Vm! �@�j�^�?����~*�E!W�A{�Eܓ+{`��Q��N?���RL�D]_�%���X=a+`G|�P��D��
����9rk�1Y�x@BM,�y2N�
�`I'T�J؈s�V=KEN��=�����t�9%C:�`CG��%t��f�M �Py���9{��="C�Vk& �	�.�(O��f��2	B0$���@m�r`�B$Tm�<��'k �dqK7� �ԩ�ݦ�R�+/�S�O��G�"�)R��_$iu�X�'	B�x�MR3$�p����Z�s��0�*O��r��V�Qa��!���8�戸Y����ɉ�yrL] K�p���
"�ՠeÒ�y2n�!6rȹ9��K���Z%LC�hO�`F��E+�1!���?n�Rf�Y��y�D�vj�ҥc���t91�~"�iz���>��^�'��<��L�A��1p��&Tm��_�z*�h�
�2��bi�g���'W��'����/ܚpe����%d�L��'�d%�!���j�}	Aɍ$g��R	�'�Tl 6�S W�t�5A�3O	p�R�)��<Y ��[��y���2��҆
�u�<�&#^ G��'��w�����j�w�<1@Z-J&@{�@�5g���R#�j(<9�4"��ء��"&M"��gRH��ȓvx�I��ɼ��)#�A��3�'�a{��'��d�<,�P�d��f�����!e�!�d�(w�E��Ơ+� �跈�4t ў��	Fّ>ő4����|�a@Ԡ/�4(��<�	C���Og��
�)B��2Do-��q�O<���� ��(��ՆL��]{e���Dܮ��ix��RV,Ԯ3�6A��/��u��"D��h��Q�$�;sa5d�,��T "D���U���'��f���8$�6% D��8�)Ei�>�Dʴ��TpdE2D���"N :��ё��aY�lp��<Ɋ��S�1)�)��n�0����g�ц3�����>��W.	6����-��XYfi8�-VP�|�'��ؔ'����B�V a��Ԓ�-�<) �C	�'��d`�¼�lD��-�1k��z��D�<���)V����)�"��^`4�����!`�!��	�-bD�ؓbC#��C�ʬc͜`F{���'e
UI ��t*@ ^Bf���'c��;U�įO�"��W�<~(�AM<�VΌ�$ýl���R�R%�(5FyR�|Z���!H� Cеf%ư��&��e~ў"~���f2��cuJ"pizs�Z�6xC�I�T��u�Rȕ�N��BC�-l`��IE]8�a�/��Y^��/B:��Q䬐��p<Q���w�q4$9�q�P�1CK�a
$��]&�ԃe�W>�j�(���=p��O�Q�شL�0�%��?�s @��{
2-�Cd�%s� }{��Zu����s��bQ�]~״����t��P�Bj,ʓ��<ٰF>l���"�H�	]6m	%N]Q�'�ay2���Y�����.-�� ��y���9�eRnݪ�D9��י�y�"<pٺf�u�aE&A���'�D=I����$�$:Dl�G/Ns��;���5�y2�ٷ6�4��IC��c��?�yR��U��"&�J.6[���n���y �l�,�+$��Y+�� �yb.['R�d���E�%"��q�h��y���<�D� 5$���LB1�0=�bKO�U@qH�"�3(
�i&�Cq�<�4k_�踓��P ��kW�W�<� )��^YA ĜJT�9Pf�T�<�q��eP`���$8� �s��u�<a��Q-s��{ AZ�M`���m�<�"��|�  x��F7<�< P��a�<��o^�O�����i�(�y�rk\�G{2(W�j?�T�$nʨ*2d��y�kL� J�yy4ᄹ`��A�*���$�@ ^��P�2�GB!�dJ!<��8���!f�ѐAI��i6�OV�(d�p��3r@�'z���"O6��0bӓb�d�
���B��"O��qu�M%�}pQ%�Ƹ����*\OP�zD� i�A��M��u8�"O&)���0T*R�Yp��,2Ŧ�c�"Or�h��$:��gE������"O � ��C1m�KRe*.�"���"O�m�w(��*�Q��fM�sy��[�"O`y�d���^%< �Cf�=mf�s�"O�(�V�V3n��в��U*�KV"Ov��Gc�$#6��t!'g��1"O�PQ�,]-��j@n�	V�,��"O�9B!H�)l�$�Ҭ�?��r"O�	G� Mvժ@����%Kq"O�判h��HXɁQ�:|�"�"O��ItF�,H�T�+��6U]֌� "Oj�W������Ri�P?8B�"O.�0���\Y��Jo�l┺A"OVa �O�5'J��@M������"O���n�9$PYæ��O��љ�"O� �ldIG����I@�G�q�~=��"O�I� �U���dh�_Z�� �"O��SAJ]P���V�p!�1�"O���!d�Gedt���.3��Q2�"O�`q!�_-{����qK�PS` �"O�"��X�;��� -�E�qR�"OR����Q�9�UkZk��	��"O�y���Z� h���O4P�x��"O�K�&�qz�B/����(@"O���=oj��a���ȸ<�W"O�t��F�~�ˢC�?@Ūe��"O�<PE.�2�LiYu#Y&~�Y5"Oz���'��*X4�ZD`�2U.�<��"O4���Ŕ�hL���E#qD��B�"O�e�7�߾0���ÕON�(��z�"OB=C�B�.(C��;��}��"O��*U#ՋM���,�7b���P"O�ik!��u����L�/]�H��"OEyF�пϦ�xBL�DڡӲ"O�����sjrX`Ckӭ#�a+��'" ��� 8Ji��틧�� ��<j�' ����(6�Q����}��H3�'zD��Gm
E;��f��j:>03�'.ܨ�l��
��HA�oΆ_'��B�'�DX�P<�<�`�L+K�
\�
�'�FD�g���x�!��MF�D���'�H){V�_	z"������>9����'Ð�Q��&gH8�*C�22�@��'���Ҧ�ߩ3<ԐY��Ս&M�1��'d�Af�n�t]��$E�7�U��'�pT�CV:{�Yr#e�Nd���'	L<�v��E} ��e�ڡ	l:YY�'�"1R��2�(�Ph؝�f��'�@�5I5FMd۵�	z��}��'�m�R� �Lq,D��̍<j�����'���ǭRC��h���ʒW�J���'��pu ÚHOv<����t�*�H�'~��2�\�7����ln�i�'�~�c끥V�Tu�aI� L���'+��u��6�nAi]�`'�J
�'����B�\Ǝ���R�X�C	�'��X�e��
<�p���d���'N��IH�V�~��6�P,SbLb
�'aZ�P4�}K��vd	! <��'�21�@��S�(`{�(]�"z�q��'[�Tq*N�)�
d�ME�k����'����q,��`��h!��cm�-��'��� f�'V�bGI�,����'ܝo���#�-	f!�&%$pL`�'�Lhd-Y}S������Y����'�̙��G:7����#���q3�'D<U��
D
G��l{��R��^9@�'�U�d"�;:w�<���$X�إb�'H�t{��L7fB�#T/�/Q��r�'m��$���&�tI�L�3I5�tx�'����R�k��!�X�Cz��r�'���9�ğ�(��	�l�)s��X
�'_R�Y�!Z�x���$��t'��
�'3��� /CS젤wg�'irڬ�ߓqu�u��M
�yB)>/��'ٳ}�V��s� �ybb\�m@���2���A��.ׯ��'��㥋�s��E�ԩN�5̌�J�\�3RN�z
+�y�KN8&��E-�&5@P8��8��[���,S� ˓dB�|�']�yC�F6k
i �B=�&����� ,�Z��ߖ<_�����6����0�R�w/�E�S��2?r���<�4���)OV����O#���ĕ�v��3ȅ>@�6�S$!�FԹ�%O�X�7ꖖC�!�D�&x�m���>V�Z5�&��4�qOp+u�͙O5��.+ҧ+J�Q� @�K9�1b�dΦ>Ϫ��q��6Gĺ<1x��ڸ,��T����gP��3S��R"�<qW7��$���.�S���n�<��N1�6���gEG'dL� ��\��-�>~tFlQT�'�p����UY�`�k0��P�tW�0�4ڍ14�ݴHh� ��h�51%�5W(��zPFq�$��a��i2~M���>�i��U9�4ڧ6�4��cO�$<Y���2r�0ņȓw���9U*�8@��ϭpJ4k�HʟR�6�'�0G��'�&tȵ�Xzẹ�dʰy� ���'�����M�o`\�@)�*Ȟ���Jw�O�^t�wnS����7%
;<�����'R "R�D�?�d�1'm�=v��X(O��Gz���\6���������H�gܷ	�!��W�kt
�bSn�/|�TEHF��'}x��	�I�K�*G��UE�HȲ��D���M�q�^�[.���`�,|�L�brTu�<"-'�!�S8"N��'��w�'?��G��X�t�pj�خ[��p�E8�yB�ح\vYP'��`��Q�% ����]��(OQ>�[��.�@����
n�$+D��fU	/���Q�,
�K�&ApEBAcR����hӚU�WY����'AH$� �� {�d-� �C�3ɰ?IfI�ɦ�����"� xR$ݝo���X�t��)`BI%A�م�	�;x|Mc1��&Ľ��.�4}:�'H�k!-N}�G4��4�E�v>��˃ɂݺ�S�͹"EzȲgC;r����K�u�<	 '����i'�14l�ex�g�+�~BF�;�MK�&�Gz��Z�'
���O8(��uޝr �+%䠌#R�/s�q�!2�O �Z`+�*i^��ï.Z�r��?U6
��&���m�6���*�~r�U5,v]�g�>;p���fW>7C�Sq@�""E8)F�FJ�Y��$IW�E�<���Oκ�C�*PI�9���ڷ`��ys��ޟ�*儞z�a#V�'8Y�G눴LH�hU��Q*��+O65��"T��U��<��ϖQziJ W&�9���s�*1�Z-.L�s��20�$9�A,D��Ð��#潀vNI�`�D0��I�<�yr^�h��1��]���̍����'.���6�j('�W7,���ȇ���.}�#�'@`x���5|j�G��vT�Ȫ����#�R��P��E�-qg��l?I��;�3�Ʌ4�bas΋9E��X�4˞' �?�1D�;*� ��"mr�4�d�O���oˈ7�����)_�xL�'���P��+k��{�,�b,0R��gf�Ր�!����ȡR|���6��y"�B�T����2e陻MM@��fSL6^����*D��� NS0.�YZ#K��`V&��B��k?a�<O&�b)Dx1�1OJH�eJ�p6���'ɛ���3
O&�"���N]��P`��^�B4���ƥ����O����B�E��=*��R0�p�[�L�N���p�D��@��>��S��-5'�V�Az�t��k/��3@~�|��	1i����gG;(�X	@Dh^Ӱñ�I98}p��2�>E��%X7I4i���b$^�ee��t�QH<�RI��ll�H�>g.
<SU'�Φ-��@@�Of��׬�g��I/|T
��ė>"�L-�d��^��$�$��c�:����<�l��E%L���+%j��K����UDG+�t��Ƶ=�$��/!1dt����.��I��
��4/�\c��� 8��4C'�@S�l���ʄU:��~2$A\��hd*A�АwվuQ�@U�	tߨ](a�'ܦ�F�`k�qrm;������deԁJƆ�%Ԣ�P����R�d9F�
PgF���.aG��bW/�Kq�B�	�R~�)�䗁|�n����ϒh�2��aEGAl1���*l��<���O�(R�!��x2��IB��i�|-r�FֆZe��$)h�p12$_n ]�WI$QZ43�E��e�D��D�f�P
��%����@ՠWv��"�%�,sD�j��/�.vH�"'�*oB%2�G�* X0c>��V%�	nQJ�"��v�Cł,D� �2��,4]�-I��
�>�3À�.���2e�w���У�01	��?q秀 j�J���d["���]	���B�O���F�2W�>��PJ̣T�er�'�i�#EoB�	���h'u{����8�,`���-��
C�J`��yr�*��R�E˚fԆa��n�/%Ɍ���`%r�� Fƌ{�rQq�+	r<7`V'�p	���ϝe����O�a�	R�w~�!��z���|����O	�����Y,�y�o�F�<�A�A���@ˢ�)���)����@0k�6(BN��ro��c*����OD�q����K�@xh'�#3���c�"O ��!���1M��Ё��8�pBC���YC$�81��	�	�p<�"����yP�>\�ꐓ�&�K��88Ԇ_�Sr����9������tz�o7#��B	N?I\����&��y����^�Zh�dL��PrqO6Pf��):�n)�%l7�b?�����������8w��%� (�y".�'�ܱ��f���p�(�?��Y2n]
]l�2!a�O@���Y���,�61u�a�W�_09�h�c7D����F�dLxU:Ѥ�0��q��~��́��	�H#���3F���<��ޘy�b���A8@�Vu�	�G�P����$�#�I�Q����4�C W��h��߬7\�]1��ڄU�rbf D�ЪR�vv@���kي 2��S,(�t�$�$"�*S-*�rc��w��6)Dj�ȕ2��E�U�!Ova@fQ�{:���-	VZ0ei ΃�bI���ؘϰ>��@Jz0���H�>�ZD)�Ax�8���M�.�zdY�d ���*%[����A��q-qZfm(D��ZP&�!�����N	��S!&���
��(q�����ȟ��c*�8j�йr`��.Tf��U"O,����?]�6�E�̑@Ix��%+��|�t��O����7�3}�-^�	9���S�i�(� !>��x���sc�Ђ"���3��12� `[321 %��ɞb���� 9�X�z �Ī/�T�$O9j�џ�K媀���t�rY��٧�ݭ\��WIٺ��c��'�x]��\$d��'S��_$tL8�e�$M�@(�N>�5�&K�X �f�?�'����B"�֐j�#��a�E�'�r�����c����OQ>A�uϖ�<���p� D�rn7Y�b�AI�H����g�g��,|����:O�����F1#�ɦOZ=s��gJ��1OH)ʡA[�%�DCp	��kYJ�s$���M	2 N5��<Sd�"��v#A�3�&�x�Kը�N!#4A�n=�)��D	U�Z�·M�����'|�\��f�r����鎣A�����o�h:ΰ!�nS��'l
����l}&��w��M,�m�<�WL��O)�eʎ��� @�`�pĉ��4���b@�M�_�"HVD���
�.S�l�S�O�Rx�d葂^�&��F��R2�4Q i'H�qO� ���Y�x�;��T��h�y�rB���~�'�BY"�8�����3ʓ^�`!��ЃN"�Mk*�I~��'>�(�h�S��&��2b}B�E���Jn�I7KK @�Vty�V��Ć�I�����E[ui"�x��� X�O�L��`�>"��c$�Ԗ1��}��M���ԟ�����8�e�.9uN����'8�hJ�/�}`a)��BN�,4�T����8�W��088ā䌃�I�,-�'Y�>eA-�yF���TbB�$��k�*Z]�'�z(��ĈH#.��|Rc�_/�X�ᥨM56��#v��PyR�2�̌:�XqX��v�ʭV�*UA𯅺A_��k������%��y!��җ>%>�!���8��L���v8P�+��]�T��d��6A!�E� bDl@��%IP|�j��R68�K��Т%�'ot��U��	l'�擰i���;/!��c�+G+������?Ⱦ�s�쒨3=��yV��#5R���M�*� �*�#˝fg\h3�{���e��y���Q�tag��?.Q��q�H/ �1�鞃"�]"�K�NY�@��t,!�ǂU紴��,ȝl��+�#��F����'dG�x[%؁��)ڧp�<y��O�Ar��J�.�q��-�ȓ@F�3�MH�FAl��!왝dyp�$��z5㘲9����I*=$T��ɯy�r��E�	�����*< ��4-�%��Bj�*SK���q	ːx�
ABD��� \����� �y�h�ېxァ�#J�)C��Z��yCL:]r���D8_ilt�����y����f�칢���\�z)
1����y
� � "�#��^\"ĉ�
]':ĩ�"Ov$�`*#���Ɗ�C�Ԩ��"Ó9ц2�֡j�*��� �A�"OzٛO�S��&�?��x�2"O:�)�XBf�Zt/L�u��u�"O�9�Ц\��X6�	'��|��"O�yd�ځPڬ�x�Am���	�"O��	w��&�`�@�E��W3\AJc"O�)���S���$��,.�Bu"O��kF*h#�����δY	^h� "O��y��C9+�-q"O�����"O\@sQ��zG��pdD%H(ړ*O~��_Z/�pQ��Y�'a��8
�'��q7�͍G�M�����.��'Z�X���9d��a������p��'&5�8}��ɠLޕ��M9�'�����`�(U�p�l�r?�80�'5�0*�-�8KI�y��j�+߆��'&^���g��%��@wQ��u��'��u�+7Ly�D��"�sm��'��hbV��� ¼*1�I�F�*�'UȜC�)��s���c1�#7����'%,���'z�$�#(_8x`}��'���2��t��`XtM��jrŀ�'8E-=/��q�h�|�EY�'�8�
�P	�`h���Nr���'d��Ȇ��7E���_y�8��'V�:Ț03�U�����xOh ��'b��ؔ����Ѩ0��	in�C�'�
�""'�bL��
P,�:?��M��'�ث��9p.��W*H�1�J��'�`5���Vis��J�5����'�Z8Y1���"@�)�_ND�Q�''h�Z� �9�܃���`i���'ʄ�P�
�7*&ڬ��.��o?t�C
�'�l���\52��Q%���O�R]�'�1�DF�����d�+G��B�'E,y1�!N#<�́�FU(8�� !�'��X�'@T�7&L`�6�G�0�fh�	�'�Z��4��\����3��}��'H��jդl��un��Mz�'�*A�T�\a��]:n�
t������"9;Ndh�W�2�� jġ<D�4æV�z���c#�^���`JW,,D��x��������\�P"d ���?D���TK�C�L:�n��Ejf���=D��9��^�6���`oZ�Daz|e�$D�P�0�3@��X�A��H��|�D&D��#1��3e����镐m%4��e�$D��Z��U FV��͂ |a�/,D�,����1P	�U���(7z<��*D����f�9��D�-m��M�'D<D�L��O^�I<�HZ��۞G�Y1�d.D��ұ�у;��+d	Jq���VE,D�`���S�
 d"���$��qJ�7D��K�g���t�0�T=�{�.D�̢�o ���X+ėnMf���!*D��{՝i��l��c�2�v��i*D�p'�M�r���2��=�&C�B�I�	�\;C!�>L�i�S+ ]��B�I	�8�f[{�q�1����fB�ɚ9�Z|j͈�.�"�����rB�d� ɳ2�� %I����N�V����H�`�TOe��IwfZ/�xB���h�"�2 7D�� ��+"-L?H,6ɐ�f�m��:t�D[-(�I�w/4�h���$ ߑ]:���DZ+S�� �"O� ��ɿu�ԭc��f��h�3ِ�k�zyb�]���֗�� w�Ht��"拑�z3!�ė�'���(R4Ob���Aգ:L|[R`3~�6m�D�Q؞����
{�p�s�
	}��0�!\O�ț���?,4ԕ{PFo�NY1�,�x r�]�c�4�;q"O&���
U�r����ķ��������X�T��A�W�"}Ϙ�8]����>Kf�b��L�<���J:()❲�	�A�6AZ�aO3<Ǵ��Rb�i��I?�Q>�c���b����2|���<gbXm��-�f�4�K��x��D,E�X\�����-D٨\iэ/O�a{rl@�r� R&�`��ITB�p=C�~m�(��N1�M#��O_��L3��/#�~dж�[p�<�C��ȤI��L��T�C�i�z��>�0�1c�1�
3ڧq������}����L�U �$��*[��1D�u�z`�U �2�.��E�BFd�'�F��'�B\�g�[�V����*d�z�'��IV�i����u�<~�*�*�'�"�ʎu�Vx��'O0A���C�'�� 'ȪSr��4����9�
�'�z%��!ͯcnB��#P�4u�+
�'Q&���+H9�GIѴ*�A��'���B%�>r��-�g�[�'���'��(�E�܊	x�s��\�#��
�'a��Y�Y>|O��#Ș����'���B"��8�P���\;����'#lqp º:r��0���&X\���'1`�c �kI��
�i�͞=P�'��a� $^1�	��
1~d	�ꝖB��{���'� e̦C��e20"	�Nt���'+2̒�A�'.����g�>H�3�'@h��

�)}�{���U}�c�
�:z,�"�ǿ��_w>�H�����|��K�� a޴~�XB`cB#"���+¥f@��ȓ\X2!�e�N ~��ͳ��ta������Fy�	ɗYR"9�E�>�p���y��7�n� �N#�Ҝs����?Q"'�%4;8��%i�zp�@s�f�,�b����ӝX���W�.}�Ǧ>� )�}�^�]
"O\6
�Jx%�� j�hFR�=u�<�k��h��[V`�C�O0f�<X�����"�DF���=V�����=��eJw4�5:�Q�ܨ���ey�H.C1|`�B�4�~,��fG��"a�����0��
>5�T�!FD�y�TB�I�!����y@��@��_P�D��|'�`%�½$�-N� x�J�Ǽ;b']
��Qȇ�ɾs=��U�K���g\����ĩ9q����M�ܖ	�WH[:@�ք��>07w�<�>�� ��� �R�p�y���:�£?	��
YB^u�1�)�IP<�a�SO��'z��AÐ�5��6=��}�P�7|O����+���#]�B| [�\��B��w���>�O�,��<qe��	T��a��&�̹8!���ȓ<x�`(�o.L�0���
�7�<�K>�����5�4�|�<!�j�\�P�Z�ϼ_O  �Fk(<a�̕/t����J�k��]Ȁg�5y@�a7��#�I��)�BPq�T�(�7D�P���A�e�j��i��}�Y�4D��Pc(S�]�5)��X�v�����6D� �g
kW��k��B�]��U��5D�Xh�E�6s.��8nC�`у�>D��r���*U�Vp�u���!�T�o=D��v%\�9`���f�1 \����8D�Dh􇏂2����oW5Vz4P*��3D����e;}�bt* J��ܳ1l<D� �e�N�2LI���Rԉ7D����ޖF(�Jc�ZT��b��)D�K�탹�X��pꆴ'M��Ⱗ%D��J"��<(h�
��UÔ1@2/!D�� (�����^�ݳuiѢD��y�"O`\!%�
�2D�'��8Xɸ��"O0��n�q~Uc$���;]�f"O^+�K�k~�p�eD�-08�2"Ol��b��~���9dbJ>o��G"O�����tް}p &�bl�D"O�	��H?�2���3:S<G"O(���\�^(@$i���5d.�L�W"O@سIB?J�0�@��K�!�>�-�!��F�>��bn�r��i�^(�0�"Ob����ݔG�00d&[F���"O�]H��Ђ7TH��d�Ql�*'"O�5 �)�ά���k���%"O��p�`ՄS�`(b�P.Q��Y u"OZz�M��B1v�{VLµ_�`�PU"O���B-�9=�a��%D=ɾ��d"O�m�c'^�a6����T8M�4
�"O~�H�]
�H�Y��l�q�E"Oj�10K��#ڪ ���H&�N,�#"O %�$�3	JYڃcȼ�0ѡ"O�i����{OP���i�.x�h%�d�D�<v�D�	�'���U� 2$X��O�8wL
i��_�&���E#Zxx&=9y^����R:��9{V�F��O���ǘ h8��

8�)��O�$pW�އs&�RBn��`22p�����r��:�r-��I$�R��q��]����Q� Yv����^�����N  ��dB\��`�Apvޕi���X�!���|�PY��F�b}f�YR/�\L�'l�	���YKd�D�d��}��!b��:юu����y��j��x��N7{h!	���bahؒ&J/}2J��(���B��C��˃d��A�˿k8��{V�=B��ގ9���i����hu�X�0e[!"7�Š3	,|O�2�,A�6��RB=e��yc�^�ӄ����
�R���s�̀��V'k������S�p���laxr眞Bض����|Baw)��C��G�_��$p"X���^��a���B"���z�����Ď�)@Rx��B
Ay��8��y���K���/4h<ǏO-��1B�@�0����c���	Df�5��O�i�t�$i��0)q�S�8����Ev��ئyy�Je+����:��P�КS����h]"��*0��;=�)ϓ���læN|��&qjdq�B�ɥAO�\������O�i:Ǧ�&.T�O8��G��+w�3a �7
�QiC�I�:��mX�eO;d,��I|Z�C�9'�,����8	�0ԃ�)�b̓	�8����"��@<��/�l������ �(�|����'��M�
��k�p�"n�_?E�ԯBr|�Yx�D��4�V�ib�Ӑ&!.�1��Dȓ�(��ɔ]�����F�)8�:%�a�ڒ.� \��'`F�Yui@݂\YdQ>�<	�i�3g�ƹ�U���+ܴ�"��^y�b��t�=�O�¸�G���8Ȑ�`a���慌<{j��	� *	��P1��r؟��6`=$I֨cQ���c�}࡮<�G>�D��cݹU���Gd�w) �y�O�	�*$i$a�Sˀ!)T`5pB�۝D��~bgq�'n�d{d%�'�hp*t��4�\����FU�+r
�G`@�Q�\E�t�
i�2�� 6mЙ��g��
�Q����+�)j�8@����,d" �6a�&a��Y%�B��I�wq��-c��i˓&�R��Q��9Ba16��	�����j�YЊ
3��ҧħ,�y����<��(ȑ�Y%�ȑ賍Զn �$�)$�d(�T��%J��,m��Y�L"}��]֞a㰫�*��" �0���|����00 ��-��+�0���EK���I��`�t�3KJ�{,����ͺ> 
M� �Q��0���J�J�qO�>=QAf�j0�����v����>�`�Q���Я,�*c>}B1tc�E{�$S�2f��3pN&D�����60�̅��Ѵ/+�H������6��5��iI��>E����	DђA 6��� Yܼ��A���y� ][nI�P�P7m�f0��aC���n�&�H�EC�p<�fԹs8(A1É� �X5!��V��l�FHT�G���e ,��3`��}��iDO� p��q��q�2|��-��_� �"O���$�=-�	���*>��J "O��C��<H��J�T7\90S"O��
_+��6��}&��R"O"��BbH�J���1�&Ԅ|.<�H�"OT@y��l$T��%�:w|x�$"O�4˄�E8=��1�-Ѫd���[�"O�@Q斜:oMˀÈ1St�x+s"O|����0=�͸����Pn�YK�"O�l�a(��4��g�3��(�Q"OLk';J ztF��>P�t"Oji��y���F*ے*k�0� "Ol������W��aE�	�	���+�"O|�(w&S���ij�ۜ��"O��r���z��qi�	w͖�R�"Of��R
8.��`���O���s"Oriq�� :y�`	� +G�\1�q"Ob!�M��~������O�
PEzT"O4�1�A��U@������b"O`]���4m����o�� �"O���u��yl����B�N� "O����RtJ�����Ԁ*->�P�"O�tX�$�\0 ʎ�Fl���"O�iz�Vc�H��Eせg�NM8c"O�iS�\'d�J��&Oo�:`(G"O�bF�R�:���\���@��"O���^�(�`X*�M������"Or�� �W��tl�D�����!�'r��h`#�vN1�D�(?�l�{Tȋ�K��������ItÞcyB��W�C�h�C0��7��p��EP#W���V�R�yK�'����h�c��?o뮹p��)2q���O�v?"��ɋ'o���蟘a��mSK�*Ar�#�uZ��҂�Y��M�r�x�kK�tӌ��[�m@�9�aa� �a͓l#�➴����[��>g>@�s"@ �UP\xHb�Q)zu��	�'tS�%�)�xr=+b�E9tHŐ@��}�$�ѐ�3"GZ��<���)�(��%Gѡ� L���~T7�^�,2d���d�`5�H� �ʭ+4�QPd�\c$|�v[�X͓s�qO�>A��ɐ/��Q��j�*/�X�b/j�|牻�HOQ>)����C b���5(JF)� ��O�Fz����doI��F��k[��1�K���"=!��@:��RS01�BI��Y^QwB�,���GxJ~b�DD-�l]�2.�V����"��D~"E�0��O>1z���0B�v��ҧ�"�F�jg)m�+�L�_�S�O���w(k��4�0�K>y[�$���1��a�$BQ�2�V��p�T�l(����'�O��Fzʟ��qAG�1G���g.@�!�^0Ȅ"O�����--�*�KAM��=�he9��'�:��"�~�S�OX>���V�NG�8���O}�u`�œ0
j�4�Od8#|Ru�ׄq��&ʮ!Q<:fޢU�Ō���i�$"<�; �v�y�^3\�XiƄ�gH:��'����$���\�Za֤Uz��h]F������ w�|�e�T4=���Hq��=/�	�aG��~��Iӧ)��A3,ϡ?'�!3b%�gS6y�"N
�4���c�O
8���4/ّ���X���
�A�u�,p��b�D�@��'���u�CE�����r?����!�9*"J�'�(D�ت�P��	'd�����j�bB�I��č*�#R�d�Ju#P �:x�>B䉹@a Y��!NxP0�ň-��C�	F���o_�V@�A�-}��C�	�(�H �A�׌u>2Pp��Ճ.8B�	�wT��RG�*jB�k��Q�F��B�	��X��q�@+0��Q
��Q"߼B�	��d�� \	�������(1�C�$Ú [C,�2o0���e-C�I�-ִD���Kp�� ��.<`�B�)� ���A3+���"%�#���aT"O�]B���0}��D�� �"Of�2Ј�#*j��P�ϖjH�8��"O:�c�H�����q�	q���Is"O���@'"^�!f�}svx�C"O�1�Ǩ�N������0�|��"O�����$�(�k�i֒(� u:7"O,i���\�,�T� ���p�D�j�"O���bG�����15/.I� "O�0#����#h�A�˃�  ʕ´"O�5`R��d+����8�MQ�'=����h����dH�8b4��'�P����!�����!
�� �'t��� Nόٲ�%��I2B�H�'&�q�� ��D�P��	J,G�"���'��cIO'"�0�cM]-p��d��'\����R�,~|b"ʅr/�=��' �$n�34tU��aR>H��K�'�((�ՠ�'\�R���Îc���
�'Z )e���#w�9G�E�1�:d
�'�H�Y���o¥�ql�,����'�2L`B��*X��N�*�4{�'2(���d(�)�L�#�'P�|i��K� X8�bj2R��	c�'v����[�ZIC�˿N�"X�'��#ğ�>�Ha�F�8 b�9�'zZ �_�:���E��KR���'�Z�@*�H(�h�%��'xY�'u0*!�Ҝ��M��b��uFp�
�' ��k���:�5YaNӀ@b�$z�'T�=���b�� �� ��*XF���'��b���uĖ���L��-<���#3̰I"+��R��Ց`�JdEJ���J
�|p��#qv��1c-Ȕ_`��ȓ? M��/�a#4��@gW[1�Y�ȓc^�ѓ��A�0�q�K؎�dD��R>� E��5+�T�A4�L%nxZ�ȓwO�PC��U�PV��q�MŞc�A������í�huB
�"V�؅����k�@ $E�i�S��.�t��Zt���c� ���:e�0�ȓnq���\>�v��ߖN��|'(mRu�X�a�eE
Q�͢���t���d�ƃa�,d���K�"�v�ȓ �#���ATDjReS$��D��:��v�+��#�LZru�݄ȓ]��X���8#l��*b ߻XW����J���RL�W�J�f(��=��i��&���B �jI��{d엲%�tl��0��`�$ɔ4�΄$�~��ȓo*d`3b��%)��&�'3�l���m�Jt���8Zp
`����t�ȓd�",�Py�B�Dg����"O�=IG$I *����SW��"OvD���;��3�6@M���"OL���Iѱa�n���iYDzH�"O00�gG9n"�I�(�JźV��y�F��X�5�SLʐnX��C�&*�y�N�(k瘼"v��!_�QӔ/A��yrZ�'ѐ��-ۧaV�ʴ�;�y���n��Y˵��MP)a�`��yH�|���3g��>�z�P��y@�B��h����*>�ꨨ�':�y⯜�oL*@ 4��*ƚ��� ׭�y
� @��fV���]��$Y�b:b��s"O2-	��_�}V��R��&.���s"O�]v��7,�����5S,�"O�T����5i�x���fH�B�j��W"O���`�ʁ]������.�ر�A"O���ϛ�o���������A:�"O���Ğ	�H����Y��*� b"O  b�%$����+��'�<�y���!w��9�R(0� ;����y���pC�$��.�f���%�yRe��"����@�<�R���mC��yr��OX�d��X�4�Le�Ug� �yޏ;x2<;Y /#��ŬM�y�����R��&�$)Kn�B5,�y͋�E�tA��!ц<*@�H��y�S)~�t< ���7��@��O��y�' �H�Ya"�N�!{����yR���}��f�U)�107����y«��@v����oΌH: y�*T�y�i��|�U!s�j(0��$Hޠ�y�	1K�]P�Kڶ�S�F�yb/�4	�j�+%�Q;Iz*\Qc��y2��ua !�U�:G ����[#�yC�
�F�;c����H�ɝ��y�!B@Y��SG��<	��Q�ֲ҆�yB!��@�V����:��񈋌�y�@��p�LB@BC��ksƑ9�B�ɚy#U����7��,R��τf�<B�I�Y�2m2��Y,έ��c�-g	TB�Im�"鉄�,u�����X)$p�C䉛d�|�P�"^�B�V�*��x��C��4|<I���,~8�-I�<M��C�	�!s��A ��˸��%GE?q�C�ɬ{�^���@I�3��,Y�<ĴC�I�|h�P�m#}�l0�W�%�6C�q�S��sHa����VnB�I���@�FQ2KHq��%ѩkB�	�R�lv�0..iʦ��=9��C�	a�(5�W�U%&U밡��.�pB�	"B���ƪB+��xӃ̟:�B�ɭe��7��=h2�4��
֊-]�B�Ɋ;=\�p�❅����1*O�O��B�I�`��H�e@�\�Z�r#a:r�B�I�k�LB%K0|�^��M�2�B�I�~.�,�R/%u=:@Q��<}2B�	$7 ��Āw�X��t��g��C�ɟ9Pp����]o.` "@�,��C��,A�Q�d �c�*ƕ�}��C�Ɉ:�e��#Y�IM.%H���:v�vC�	�S���,] :$A]�����"O��{��K8SG������8ƎI;b"O=�p�3���2�������"Oڥ:�(��/l���4O%y�P�"O
�"h���T�E-�'�>�a"O@���@�je�`�k8i�h�[�"O��s�%|� ����Ȧ"O!@��@�4Ϝl��-�.��U;�"OV�lK$B�4(�l�h�0)/�y���[�"�J�\�|	�R��yrə3q�̔k��U"����[��y"e�2b*�\k�/�&;�������y���.�`.7(�� ��ъ�y�n�M$���&�����\ȝk�'`�i	&C@�2�ح�F�9D�2�*��� �T�щɑy�h �G"��Av���"O:[P Ε����!U }^��8�"O��	�k�(+�D� Ȟ0#Fu�"Ox��PkE�$�zI���/�jd�A"O��;�Οv[0S͋+Y��$"O���ƯҾ'�9�ЋK�yy��"O�A�'Ѩ5p!��H�Bv� xP"O���,�'G�}���S�&mB,20"O0)J���'�0�:$��D]��*T"OB�"F><��Y��H�mXqX�"O�;(]&%" �H�?�v �@"O�(B�m
.�=����l�"�p"O@����	^εr���+��[�"O� �������h�p�2B"O�(�fG@4K���
�ᐅ5H�"O���U�^I�pMB���" |ȪD"Ox�+�쏛K���b���o�y�%"O��2&������*��"O0�RNB81�K4-E8lG��R"O�Y{b��L�2�ה (���P"O����S�������: lAY�"Ob�i l8QPk���j���"O �y����>}rsH8Q� ���"O��"��10��	��fF|�)h�"OLP0J�XW�q�d�2n |9�"O�	iS���1F�=�D�.yr�X�"Op
��1�x@��º3r Y��"OJx���\#v��@A�#xH�qX�"OP�h�(�&w"�e�� �	;$(�"O2��w�8$�Љ�#�ܴ'2���"O"��-\���cDHU7���X"OVy��G����y�,��SԞ��W"O�����\%@���p��)ɒ �"O�iƈG;X���L�T�P|"O�EpŅ��I)B�bF� $���b"O���e�=,	�`U�T'Y����d"O��*����h�n��0��	�X$�"O�`������ܐ�pg� �R�"O$���l+n��e�Wg�J���xP"O��x�)t��$G�d�Xr�"Ox��3��'%z1�g�	m�q��"O.}�6�'���&�4)A�bF"OL媀AѨ8��!��ʤ?=�,�V"O)فF�#��PS�((��)�"Oa	F
S=hH`���(a��ٲ�"OpD�F*I+;�~�	�E�I�e�`"Oޝ[����t7�X���+�(aE"O�#2�, �L�6�B�Z��e�2"O9�u(�< 4i�V�֛G����"O&A�Q+њ�*9i��ٽ49Za�c"O�Ū�deR�A��γ$�8��"Ovq�'Oώ_�<8d�W�I)��B"O��ʑD  LNN��R��m��Y*q"O��v��'m@2�T��,.�xU)S"O-
"��3A���A��<Z�t�P"O)à���-�l�b�/@!<�pd 7"O1r�J��i��	�5�<l��"O~4�s   ��   *  )  �  5   Z+  /7  2B  �L  wU  9`  �l  t  ~z  ׀  �  Z�  ��  ߙ  !�  c�  ��  �  (�  l�  ��  ��  2�  ��  ��  E�  ��  m�  � ? )# B0 �7 �= (D NH  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d���uܓ�(��U�R�O��=�]�7�y�ȓ=I����7/�ňǇ�(BD��4l,��jX	~!�����J(�~���mo�kǤ��Y&U��C:�T����`U㡭
)3W2���l��^�>ͅ�,rҌ�(U0BAƱ{4)��a)}�ȓn\��2�D�q�.�C��E�1]^����ēp�8�ѥ��;j�j���9Ec2���Zۀ+гM������!x�y�ȓ<TL<�G*|i��
��4Y��ȓ+�Vu�E�"b�
��KK3n7f��ȓU��#t��$�}"��R�"�!��� �RaD���z�J()�&��O��M�'lQ�X��Ez:��c��Ox�>���Ā�dȄ��ڟ$�Lё��Yj!���O����m�pq��Cuh��P�6qФ�|R�)�T�x����"]d�Ö�P�]}���6��D���)5�L��X�zM�ȓ]BN�p�/�6�L���!/b����2�)�'M���b�#)D:ɡ�xH��n<���@���'�&��!�$ÞK؞A�'�	�X�[d� ��*$(�c��B�I������/�0����2b�8�Ӡ�U�Ş%\�����_Ц���O�uDyb5O��E�d�+��d��L����"F=D��ticc�#?ɣ���;oVd�b(�.�T�js�^x�<� �(��e��;(��Ѵm
(3������O�����Pef����Aۊqr$�7��y`�r���I ΡQ�X]�$#�Tfj�jt�6D���6Ə	'D�(���K<�<(jSC!�	W����4J����H2*d��a�E%���=��S>p�6����T)P�<+�ɓJ.��Il���r��_#km���љtXx��5g���E{*��O�
.�j�c��)�V�Y�"O�$P��z\ܰv&��M�`��"OR�Pr�L4ġ����'p�9��"O8�Bp!-G+��SDc�a�U� ��E�S�O!.p�A�#�Ca�.�|�	�'<Z��#�3����#Ĩa��1���>AA�#ʓ��'�bYq��]�r<XYg��>B�@��d��Ë���ǺQ�
� �S8sW }�s+���yR�(lF�1Q���i3�(�3aE(�ē=���b?�p�aA�R%��v��5M���-;D� a�"G!2��@I� ��C:�I9eazR�$%^l������*�Y�lر�y�	�[4ީ�4���#W`A����~��)�'-�����NR�.~�`��	 Fd��<qJ��E��ǈ>C�FX�A/O.b�$�5I1��'azbo��yj i�!c�
`��h�����/�S�O��[�bǡD�0�ɵ��;� ���'x�֋A�)M2�q�4	������#�(OD�=�OnV;�`M�^�.T�E��e�1+��(O&hR#C�X�M��] �����i�W����_=�=j��+�J�i��Ҥ�ē�hO�OV�.5�}���?r�B��6�y� Z-5��j.�3��g�����'f�y�&�r&;աMN���$�1� B�	�G8��;�R4� h���WH����8�SI��p�(<iwh]�''jc�D��\��t!���q����u�.%����I^}2�'��)�.E�� ��-J����]�J,��'��Y�Ć��$-+��W�~ �a9}R���㉉�d4sӤ��A/X��)��6�PC��>c��e=� II��R6�&��{槅�\6�TL�.rC�\���$}B���Nqp��wg<1�DqF�͌j�n���T?��F0z���n��!Ht�����'Kў���!��$Z�u/��1��C"}�l���"O�C�,:m.t1���E$ir<h0�"O�թ�ʐn��E{rPW��B$"OD��5H��c/��+��Қ00����"O}�5E��\%�APU1,�S'�'0�x��dS5%�09*�B�Qr�9a/�'�!�D�9CmV5RV���`o�Е�E�"y���	T�O3.Xs�⍇]�p��o��u���'�Ѐ�"��7 	�\�eh	>�>��}b�'%R�@���mfڑ����6��yr�'F<��H�u���Z�E�"]ꭘ�O���U�B�J�CS(������JE$Ș�"O�� �(io᱕a�;&i*�"O qb��b}<��C��*%�M	11O9����/��UA��J!V=F�����] B�ɜ
%��y�)Ֆ�&������&�C�*
Q0�§���0��g�s�tc���I�o.��D�N�x�JĔT�6�Ie��0� m��1��E�WJ��;���̨O�L'��XH?��I����d��,�'���J��%D�D��m� 8�1��ܧ�XR�C#ʓ�hO�0nE��qWF�hf�a���]<B�I�*���3UfU�y���J��l��C�)� ��qH�.$=]��m�����V"O�ӂA�6��Z�&�:�r�"OFax�k�5r�Yq%#��N�j��%"O(���A�<�n���0!�����"OZ�h�%ΰ�Ȕ'}��
�"O2��F*kjШ����V�6�B��'I�X��3�E
�89����>��z�*����_> Aa�\#|NHԆ�GZ~�r� ,��}�C.��3a* �ȓv�l S���VhrC�;}�܉�ȓ)�Za�f��>np����l��[�2%�ȓcᳶ���gV^���fłu��?y,�a8�|�G��?�l�Jt�b��튄�>D�ȩ�D"�����Z�	���+�����x2��/+�:�y�E�j���zb�β�y2�\
W�쉘�� ]�,DBf��y�:jh���a\�\Ihq`#ݬ�y�dM�o�<�b猟[�F-�􂖗�y�� �Є���ڭM��������yBNTHJ�"�Kv���"�y�eŹOOʀ��;Es�����?�y��;.F.�#&�E�����ጽ�yrc<%�8�²�s��(I����y�+׋{�Ρ��i��D8d*�
"�~`�>�	�3*�q��I����c��ڸh��	g≪Kh�,�,�^k���r�Q�OKjB䉸M�| )4 խS߰���ʐ�v)\B��*("d�u�>�lAPpAP,~�C�Iw��\r%A�.p��@���K�B�	"ߖ�"b@3����CE�]��C�Ɉ�~Fa*LN�(�(�4
.�C�	"�XP��@#-�x�J�EA)R�zC��8|�ъ���Y%�Ը�!�-5<C䉠���4fR�1~���ƴI
C�I2UFȄ��N[x�h|RR/�3y�C�I�^�
���Axp� ��<�hC䉖>v
�j$�/,�r$�W<`FB�	-A\:���:O� �yQAcD�B�ɸX́�ᆶ"K����CT�=!pB��8y�R�[U�\g�f�Pt�ƨ9.B�Q�����-^�h(q@�L��B�$pvว��(!:���6Y��B�I���h�l�N�d2v�15dB�	��Rq����&��@4zB�	M!\,@v�Čd�����W_#^B�7_��i�.Z�NXTD�g�41cC�	g�Ȁ@���?���unXzpC䉜)Zʴ[����w�$�s��,�B�	Ad85�a���>�0��Q�\��B��)@�ʳ���~��}C�ꛐw��B�I	`���u�s�t�17MN!9mfB�`�^��� h2�MW��-FQ B�ɳ3�YBs��).6����S�>�C�I=/.%J��y��)��E#c?�C�IJ�A�V�ڀ3�	k�؀Vl�C�I9j,����2H 9$b��kg�B�	P=��$O])|y�1��W�-�rB��9C��{��S
P��	�$d��q��C䉽nN�ꆤ�1#Ud��hóUT�C�I�؄!���,77���"`C��rB�	xO���U�%�t���L #t	C䉟S�~�ؗ�S+5F3t��J�>B䉝Jx��I�fL�=}Ɲ�w!��	fC䉿m�llA�gJ����F��JG\C�)� �uQǄK�'T�iB%K�rU����"O��#��@�F�e܄-�Q"O�г7��Č¦@R����"O < �Bߝ���� /�0O��q�"O���QB�?E��aY���33z����'#r�'J��'���'���'r�'k|D @2R��p8�#�
9�T��'��'~�'X��'��'��'|b�[�kTl���ѫU�T���'�b�'L"�'7��'���'�"�'^R��fދR*8�Ag����3��'m��'��'lR�'�2�'��'w��Ӏ@��i�r咖��s�X��v�'���'$��'�B�'�"�'��'e<�i�-�6����POJ>O~܀�'�"�'���'�2�'���'QR�'��8�V����/�=\�%�0�֜�?1���?����?)���?���?	���?iU�ԑGY�s�ݲd���R�C�?���?���?1��?i���?���?��jA�@u�u��-Z<iP&إ�?	���?����?1���?I���?A���?��䂩TQ��R�k�G�b|+tʙ��?1���?���?���?��?!��?Q���iB"�B��zFh)f�ۢ�?����?���?Q���?����?����?1���3%��!�� �n̄!��S��?���?9���?��?)��?q���?��MS��;-��<�r���K޵�?���?��?���?��c��'��ċ}'�ң���ޤ�-7")�WR����Ty���O��m�!���`֚^�5�)_:az!r�8?�лi��O�9O	mZ=l�t1�%$�u��� X�1�l��޴�?��L\�M��O��gώ�?4��J?}��ㆼ���"�(���J!��۟��'��>�BWoW:.%L�2E�d�hW�ۗb��nZ6.�Hc���Z��y�,©8�$�x'�I���/��P �i&6�`� ק�OH���R�i]�D�>c�$�jq��b�m��̆K:��F
�p(Q�ʢ=ͧ�?� �X�T9��ŷe��y���<�-O��O��o�T��c��q���Gb���������P,CY�pA�	$�Mc�i��d�>���К����}�ڌ����Y~r)ȫa/�X�aO���OW�pI��*P���5��	S���oK`2��E����'��	�"~Γ2��jsD)RH�:�N[!?2�T��&A
���D�Ԧ��?�'m?J��P�ä=�az�/W�l�Γk4���q����"FŎ6-:?��/��!dl㖃��c��8;����Z���0K	M���.�.jl>����8w�Ā�Z'R�:��d�wE�j�Ne¥BT-��C)p���m	�����$��\�\�W�X��~ ��iՔtZ*���˲wA�J0h�$�>��f&��t��ֆ_*X:��k�D"�g�J����P�_�H@aE��re.��*�=S. U�4	
bl�ʖe�mS$�W &d��J�.��J�H�E'�1��Y@t�1Mդn����c6*N��Q��A��<�
wJ�Q���#�^I����"V� G(`"��� f�H;g+�@W�e��#�<;H!l�џ ���t������PmN=�קK��q/�,��'���Ǝ,��'�"�':�d�~�
��^0թЎ�\��S2�Ʀ�+��	�Mc��?����U�x�O�l��eO�+*���aQjJ ����|� �+p��<����?��g��?!%!�O������H���Ǜ��'���'��b�8�4�����Op8u��]^�pi�� W��-�s�Am}��'"�ӄ��',��'>򌃢v��D�h\���AS��_'�7��OZ�*�[�i>���Ɵ�'��|���/@wZ���i�dE���)vӘ�dYI�1O����OT���<5G�"['�̹���~V:��F�R�$l�B�x2�'���'��ȟ����-��(�"-|�f}"f�+��
� *�ǟ���ǟԖ'Y �0Ed>��vG�^�ڰ�G�ŀ(�8<�@�>����?�����d�O��d(G3���	/2���Û���o� ���?9���?�(OJ0����B�ӊL�F,�p"	�)Lv����}j=*�4�?�������O�D+�1�h� M\�1��y���88#��k1eϦ����'��<��*�i�OR���nl��T>]��"헹vȊ�"w�i��IП��	3U��#|2��Q��I�����"����X����e�0˓j�,a��i�^��?��'L��	. ��Q5��}�zT�O�${�6��O���X"	����|����&�x�@fϫ9�xpsg ر"7^AzQ p�D��%&�Ϧ��͟���?E�I<ͧ'{ �A���C�H�!��F�6��j5�iMjqX�����(�3���@��ןb��5�f��,�pa���M���?��	}\�{בx�OS��'4����%��'t��gB=XpF�{Uš>����?� �Md��?����?�M|(�s��k��Ό#i��v�'R(�h� �4�&���O�ʓ��r���"%ɾ�c���ľhRR�iO�"=��'d��'��P���]=2w�p�C@�o�֩�Ҫ_�k1�u8K<I��?������OR�Ċ�h4y�UG8t��Ո��ay�����Oj��<��}���q�O�6��!��=��1@Ն�1|k����4�?����?����'�Vx@Ì��M;1+��A�A��N#hn� �W�V]}��'W�U� �	�/ ٕO��@J�3�� AN
�:��qb��!>7�6M�O��L�I�8;��c)6�ү::(A	�-�Y8�̌xl���'T����e˕N��'��O+t��p#���	�H[?X�VM���*�����A
2;��c��g�? �x��ƛ(w�( ��q�-��T�D�I�*
j��Iڟl��՟$��nyZw�za��䍨8�e Т�7S^�OF��:eBd�������N���/E6,@�ZJҶy��6O
!_���'"���?e���$�':ek��O�.�
[�/Z,��ll�r����*1O>����?��U���	U�Ea��0[-x�)ٴ�?y���?��A���4�����O��	�;��v��(bb"�u�M)~�B�yb�M%� ���d�OJ�	-�f�I�ʜV����$�Eh�7��O�ȫ«�<	��?Y����'f~��ƫ!�ŒPA�7P���O���p�I;u���˟���Zy��'����V	W&n��d�P���	�AL�ep���I韀�?!��+`�@[b�'4���*�r������)Z����'�R�'��	�` �'�d�d�?Rl����&^Z�������I˟��IO���?� _<tXؤl�++���BdK���D��-��x��?I����D�O��!�|r�Aф{���R$�D��\+�i����<�F�~��D�$��鈬U�ȭ�@�q�7��On˓�?I�H���)�O�����I�t�H�.y � �3�^�#��Q�����7w�֝~���(��
�B�N@aen�:ndb��?��nN��?���?���b.O��&����@�27�AJ�"���gybc���O�O����4��� ��|�b�4�59��?i��?a�'��4�n���6k��As� ̪ ��Y��Z)Z0X��'�������)�O�A˕�
su�-�`cL9eU�]IU"H����������K�h@���$�'
�O�ࠤW|ixi�pC�v��)���q�'��f���Oh��',`�t�0Z0P]�ՙOM	l<R7m�On����<����?����'}�487�M.dQcǕ2��<�K<�U)QT~"�'g�X�8�I�O� d�C'��bd��LI�>~��f- by�'�R�'��O(�I�d��M�QN�x����B�)T�|7MBv��������Iyr�'����ߟ�vƞUv�A��K�	E�i�R�'�r��<�e��MP���#|�p؇���-��-���>1��?.OZ�����'�?Y�
�mj�����2���ؒ �
b���'��Ov�ěB�4Ya�x��4�9"'�Z/X/�IG��M������O��F��|���?��'^i^���Tq	���
��U���O�E���O�1O�S.$����E��I�.-PӪ�6::~ꓪ?i�Ş�?��?����r,O��s�8����4U.�} �⌧d+����t�@��j��b�b?���C�i+R�E�~*` ��a�r<����O���O�����*��|��n��h�e�:r���2`bC�5�\hհi+r遴!������$�z���
Y�5@����L}mZ�X�	��P�&!�my�O�R�'���
: ���!�p���h���'DV]�<��l�;�O�R�'5�o �˷g�&��9�@��6���'�[4R���������L�e�$="n�5���P�'�,\��0�'�ֵZY�����O���<�����24��T�H���D�--�n�CE�����O��$�O� ���.t�ϙ�k�<��ą�f``b&K��ob�?�����O4�
"�~���A�02����D�5n�H�r�y�h�d�OX��/�I˟#�d &�R7�ȯP�����ЇY5�\EEY�h��I����	zy�'+&�r [>a���e�g�W \�֩Ȁ�R�2u䠺�4�?����'w�zU�ܩ�ēHx��� M�+��6K�>B:P�lZܟ��'s2�I�4^�џ����?=q3�MEE@RQ��z��ۅ`Å��'�Rl�������y���qC��H�)�M(�-�+]��P�H��P���	ş��֟(��]yZwf�}I�lI�0�(�H�GB  �V���O��d�,
���C��iΪWB���@��Bĕ`*5�Ѹi��u�'���'7�O��i>��I�
��x��C��$]$��̪y���4.����dKT[�S�O���5>�SdJƜ �pc�&q�6��O^�� +O���O������$��cm��G�ؼ
�9q(���'���%�i�O��D������#-]�X���X�k����`�d�4�$� 'D<ʓ�?���?q�{"�M$���e� Ɋe{�������T��H������������'�I$M/`H���S"^����"�A@� Z�S�<�Iʟ���K��?	��Ԫ(
��1#ꓑ���#iFk9֝rU`~��'�R^���	�)-�\��?�nl�3��E���T,̘Z�,m�ϟ$�I۟��?a�r�n,K��ۦA���8W���L�'4�h܂��>i��?)/O<��C�Es��'�?��Z!�殝{�ڨS1�]a8�V�'��O���.BX�T�x�BI��aٳ�A�RA��A��M{����O�S �|B��?��,��D��+^�bV�|8h����O���-\a�1O�S0Xc�92�³>�b	)��@�i>���?�'��?A��?	����(O�N^�o�`⳨P7;�D��W�����Iߟ�; �� }�c�b?u���;y���R6�($v��*dF�O��d�OV��ퟆ��|�l|����%
��n�]��<*�i�
�G��=昧����n�? ���% �a���M�1|�aAU�iZ��'4rj�$��i>�����>�,��0)�o��2�D̊Uj|����<(H��%>�I�L������[�ܩ��� >��n���h�$a�y��'��'�qO��u�Q�6b+���"xZUCBz}R�ϸ��:�O.�$�O˓�?�b��<��l�t+ �#�r(����u@F����O��$�O��@�ɽZ�p�"�!�!�,���j�E�"'H�]��?9���D�OXQp�	�?}�sl�<�X� Y��^4�W�cӜ��OF�d1��ȟ$+�ʑ>q`
7�ϝ�r�`��7W�lJ��3	+�I͟��I�L��ǟ�x�ș��MC���?�@L2 �p<��)@�8 ��+4b�[.��'m�'z�	؟p��g}>��Im?���	'T��-� h�����J���ޟ ������M[��?�����)��+��E��̖7F�lc �.��f�'�Iß�pG�n>$��s��2烒�g��M:�C�
h����i���'2��б�a�"���O������	�O2��fl�R͒�N��U��}��dJ}��'�|�c&�'���&m*�x��]�/K����� �����Hꛦ��*��7��O��$�O�����D�O ��̒>N4qӆ�O2�@� �X dc��l�;Cֱ�	ӟ�I$a�b�[���?���ݕi?`(�@�����'��M+���?��\t����i��'6��'�Zw�J��3�F&..�3�o�\l�ٴ��Wkxm�S�4�'���'�����
Mb�t3���4P��]���rӬ��ł}��0l��8��ן<����)���臢��=�̨QD�����@ ̮>A��J�<Q���?����?9������R�*��uԋ꺼cC�Q��:�ĩ]٦�����	ߟ�+���ʓ�?B@�'0B���$)X�q�Q�� Lp0�H�'�R�'�"�'��ӨX|P �ٴ0B�5�U�Rpv�9 �G'6�
�٢�iO��'f��'Z[����4q4�擬j����'���b4>؊�`Vrf���ݴ�?!��?1��?����<(x��4�?���� �S�ȥ!b��� J�t�1�i2�'}�V�|��	���'���l� �f-� h�iY %�9o؛F�'��'
�̒�1�7�O��D�O�)ٴ�R	�3(V�&i�Ă��R�
�	o�8�'��움����'x�i>7͝�n���r�өN���o�G���'^�(��V�7��OH���O�����~�D��R�N�z@^96Q @B��X�;�"��'��B��iy�����2%P5�ք=��h��r�ʅE�i�L�r�b���OP�d��N�	�O4�$�O$����<F��s�$��q���a�����]������	Ry�O��O�2n^4x����I[�L&�=����;A��7m�O ���O��J6)���)��ٟ��Iퟤ�i�=;W��pp���'zw>�#Bc�>�+Ota�������I���:f��`�"uA"�D*w���� ߢ�M���HшҾi���'Q�'A��'�~RdA�Eg\-c�	�n� `1������ί{�d�O��Op���O�ʧ:� �x��E=�~PHL
�s�!�V�ƉK����'���'�rh�~+Of���>%NZ�gk�!CĆ���Y5^�%3������l�	�h�	П����	�McE
�0Lƕ�ૃ�u.P��-*��v�'��'�R�'h�Iӟ�+u,y>�a�*�D\hzCS78�~(��
 �M����?A���?	`T?�
paQ��M[���?��L'd�$�K�,}� yB��7���'Q��'��	��n>���[?Qeb��8�.�1]j���O�٦)�	��@�'#*�1�:�i�O��i�i�^�6�H=*�Ů�J�:vm=�$�OR�d�$l�\�D(�T?���H	PS���QMҼs�DaP �z�:�"a��3�i�맪?��'_��I�gt������s� ݛ���R|7��OZ��Ww�z�b?�d0(���:"ij�:��tӮ,�gR¦��	ڟ����?�QH<��a���Kn���&R.Oɘd�t��˦Á�d�P&�"|���X�t��v��2X��aҊ��n����i�B�'J��ӿwÚO��D�O��I(-���
#�uE�5�	�T��7m9��@�G�Rr�ܟ��I�0�L��d�9��E�zx�(�`T��M�I�����d�O�Ok��oﰔ+ L]�: �-��ݧF:�I�5����IVy��'�Ҕ�4�X5r������9�$o�Tȫ��.��O��)���O��d�;5���;�AQ�\D4�mL��
�A";O˓�?���?I,O~�"q�]�|��m�Y��1r��(3�A�U�ϟ��'���'?��ث��3m(%�!�]$jeA�P(�x꓍?����?�/O��)���m�J:�ir+3&'��:䇀�
0|��4�?�N>����?����и'G"�X���aE.��3M16f���4�?����D�%0���'>���?�X��	VYԃ5+@2<�Z�E����?)�� � Γ��S��M��_O�R�7���h7���M�/O� �������~�D��δ�'
ڰ� *��B�^�{�iʵo(\�q۴�?���_4Ex���
W�g�b��a�؝}Kc�N#�M��4���'���'����&��O�={���dV��
�h޼+� eq�#���k�	d��'�Ԗ����O"�H�GCw�>�@���h��ҳ�Ϧ���矈�	�#bt<�I<)���?��'�N�S�S9k���M]ID,��4��2+�Qt��d�'Dr�'��3䌓�46�A�"T`�8�
vӚ�DJ�M!�$�<��̟�%��XG`�pR�E�'�����'$�C(l�͓��D�Oz���O0ʓ)�� �L�P$S[�5���3}e�������~F�'���֟hjB,1G&��G��7����O�?�`��	uyr�'7R�'�剥Q���Os\��p��=m<`���5"���O��$#��?᱇<�?"!Y0����P嚃[��K#ă�-���'!2�'Q�U�PE�C6�ħ1����,���� ��2���SѶixў��	�&3��	֟���i��`�.P�SFT�ToM�l�֟`��ȟ���%h��	����'��D��?[��z��A�.����4�� pRO��D�OЌ�Ì�&>1O��3Bl$i��h[j9*L�P�2QVl7��<Qk�Fܛ�Ķ~R����(3	��K�A�gL�1A9�*6�*3�p��3񤞫05H�e삾���d��<$��FG�,*�R�'���'@���'�Y>���æL�2p������Ɂ�Mc�+?���<E���'�B�r�:vF�eH�`/,d��p�iӺ���O���v<%�$�I��|�m<~�K�B�"20)L�0n+L��>Y�b^R̓�?Y���?�Q1N}���1Egkf0@���;	h���'���Jc-��O���$���x���"Ce��
�F�d�xK�U��1 �4������I��$�'[V��@��M��ǫ�e��Ly��H,LO\���O��O^���O�!y��?���*�k��?bIұbE�
1O��d�O��d�<y���a.�K$;h���e!/��I���On������[�������a�"���J�h��Q�L�ʨ��'2�'}RU�PZѬЇ��'	(PŃ�"H�+�*=  � O0`���ir�|��'RgǾ��'��R��S�>v��R�(#MJ�J�4�?���d�2H`Ԥ'>����?IR��ǣE���\�*����m3���?��: $�Ex��V����4r���V�B54)�E�i;�	��`��ٴRD�̟��S����J�>�N��s�
&[�9�b�22���'r2iڧ�O����b���fA��+�m @�0�i%F����*�D�O4�$���'�`�	�rT��L��,T�xP�F���D�ߴr��8Ex��)�O��)'����pa7b�;�Tm"������՟`����v�bN<����?��'|� !L��`��$
�؎Z�����}B����'�R�'���\��Drê�	NV�djv�e��7�O|��ȕP������o�i���0!۾6� �RT�å3�<XrdĿ>	!�z̓�?	���?I-O�m)@�ȍo��0�f���AGY�E|�$����ꟸ&���������h� 9�wA��C�GP�0Kpb������IPyC��I1��S�˜QѱJ���C�,�P�'B�'�'R�':�T�O�!��-�w���b��?#�.����l��֟�'+�H�q�6�IO�}4��R��Z�Y�@��)��ml��'�0��矤��:�	�A�ti�u(e?(�!�11�7��O8���O8�$��w�����Ovʓ������/�5R�-����$@S.cމ'�V�P�B.�Ӻc�K� @��6&H�)1()��FK��͖'�6 q&iӂ���O����^)է5�������&΂��%��f���ē�?��9}r�O�)�B�a���Z�D�dD���M�G�,�?1��?Y������?�-�BM�M�8���Q�G�f�|b"��F}�/C3�O1�����8#'�A�v��_U�M�6G̓�^�m���D����xAGCTOyRY>��IK?q���'n�b�Ґ�Y��@�.�3��Z�����	ҟ\���ќr:�K7N ������ݟ�M���uLօ�5�x�O���'��P@zQ� �:q0t��g8�	�'B�A�y��',��'2�'��`�TL��S�bYZp�[-
g@���ų@���'3"�'*r�|2�'+��	8!&��F)��Z�(E��HM;���������OT�$�O�˓I��:�^�ä��0Q����c�	$�@�����O<�+�$�O>��K"_��	*�`�ҩ )\�Ʃc���{t"��?9���?�+O�jx�4X��(p�&��Qz�D�e�ȑGH�X[ܴ�?1M>���?aUe�_�J��ˀiHp#�" C�F�zXoZ؟��ICy��J�������㟼�[GF"y<���V�b�p[���?��RgZyDx���]��'śv^��qCе\ a¢�iR�ɯZ����ڴ8�����l�S��$&�Ღ�W�"���� C����'�R��>�O�� <�T%ɛ��)��͌|�P0���i�U��s����Oz�D��L|&���ɶ*���+����2�"`Ԧu�r���4?�j,Dx����O@�� lLO`�e1�o�&v���H����I������	�m�v�'��S�P��U%� ���]ʺyI"#��L��m���I�ħ�?A��?Q�,�+)�2 p��˴�ps�
�*}�6�'zD6M�>��W?��	����O���R
�j��2dʓ!o�F�pr�xb�|��'�r�'���'d	rB�I���3o2�����M�/�b�'���'-b�|��',���)B@Qa��R55�!�L؍B���ݗ��D�O���OZ���O���f��?9Ӵ�Z�픀JE	��a�5i��x�����O���0���O��c;b�mZ�H�=�WY7(��h�6`͆P?�ꓴ?Y��?�)OY2��Z���'�� �a�,úo�:@س�M���<��iL��'z�O���.�I$J�(4���_8��x�ey�p6-�O4�$�O����7C����Oxʓ��F�
�њ�c	q�r�x�P�mK�'��T��k�g)�Ӻ#q'�b�0tb6"��Y0�B
�+
�yU)N� V0�K�\\�$?�ʑ�xB�R JD���JO�G�Zu��c��y�'X@����Z�9Р/�|uJ5��$]>VBK�'�$0Wo�0��Hӭ&;��̐�τiٞ kҩ��;�,��	.����vC�(%�$Y���� AMM'mx��p��
;V>T�1�]
���we��O��t��'��#n�P��5����5�4�-:�x��BH�t��4˥��x�B�'x2�'VD������ >�ѧM�//	+e�Y�zT����OT�2a-ƙ~]����K������"sg�h��!1:��"��(d&�������cA޷>�6���Пў���XHqy�K�#D�X�qi���X��Ox��>ړ��$�(%�t���ͥS�mɤ�M�b;!���O�2�9+r�D�rm�S�0(�ҋv����'q��8zNH�;�4$n��H��<g���8�
����?9��?�f���?����j�\�lX:�`O��[�@[�hӐ�cq%�j�:����ܫ2n�A:e��',>�Dy�&�^��a����9
�� ���Ft�nA��	V�N �P)A_�l��+[�a��mЃޕ8��'�m���?)���x4a��<%Xׄ�<�hO��?�e��:��z�
�tPx��{�@D{r�S!��[��n؉�� ɟ�y"q�V�Į<9'�K��џ��O���S#�"����n_6}+:���J��3S�'����� ĺ�;�#���H���S6GZ��]�m����o�|5�w���5��pŊ%�ð8����\�池d�^w����F	@�5p�ѸJ�EdZ�@��P����O��d$�/_�1QD��:�u�S�G%���b���K�G��~┥+q��w|��/�O@$��*3��=�.��Eg�4*�����l��S0��M����?�/�|8S���OZ���O��D��o΄l��)޻fiJA� $]�9���E�k�<BE�O��P�矤r��5Q���&�Z��m9�DS�N-��r6��\I���&j��"~�Il�(��V/�1��U� �PX.�v�Bϟ�:�4_��)����z˓V|^<#V�#mٌ�dj@�2zq����}��[.=K��J����FD�Ex"�=ғF#�	�E)� ��[�&�~�c0d!
o�=��ߟ|(nU7@� �	ß���ß�kXw��'�zP�e��qn2t�A:�����'��z�Ǟ�#`��t����-|�^@[��	dI�=�N�dR��f����牆ez�P�U4�̱�q ��"؊�I:<�0���ΦIzJ<a���?.Of��0��37c��"Ovp a�Y�xhA�� '\X~|� ��x�'�S_yRmυ1:6MQ��9s)�";"��P���
�$�Oz�$�OАb/�O��k>�Q<O��]$#�Z�q��a���9w.���\��w�@ي�i�(-��iPB��k\|i��ɉA2���E���G�?vrE+JA�o嘍���>�M������O���'lFa;�b �DF>M:b�I�|ź ��9����!�74q��  u�B	͓Y��Icy�$Ю��7-�O@�d�|
⍊$u�lP���L0�y�	�.�|2��?��?��M�1�M����a�n�8��бW�,I�!�B.Q����;S�?�1�%��#��j^R^�ђB�yQ���G�O��d6���O<@ÕE_�yd}S�������O��"~��B��,_��@YS��[���q%�S�$�O<Q󧄣g��d�"��	0���R���<��.��(��Iן�Ox�S��'��'BD�֩�#5=�1�b;c��(a@�Q�S2%�(N�5ԧ�'��Op� �Ĕ�E���`��o{zyȖ W�=�	YS��h����O?����B,|�0iX�$NѺ��L+���2���O�qoڬ���$�Ou�I�P+����A{W��ق��!�NB䉬Z6@Qf߲)Ö|�$��#d��#<�s�ɣ��D�:U{����Ȋ,&X�IA�p ��d�O�����u����O@�$�O2\�;�?��|�,ʖg�`����U��P0�;����6I��h��0�С��\8b��LHD$��JlP�i�h ��>���	��RUF{��	$�r"B�O۴���B�$�� O!'$��'����$�Ob�o�\	C�FG"t[ؕJс�-��d����?��c�3h�0�33�m%�;���0��Gzʟ�˓v�TA�ĳi�Q!,&:f�lk��?
�޽���'���'A�,R<j"�'x� '3��u�צ=F�}(���_-�Ԑ��O,�"$���vE���ą4!����$^�D�04ůg���5�T�$��(�	��w]���%'�b�5`�/@膓O�9`��' " 6C��8�[>n(l�x��X8�R�=��<����b�D!C'�>]�n���"W�G{
� �K���~PLb�����8y�5O.�mZʟ�'�V�	�m�Z���O��'=T� R�a@*w��#���j&�I��F#�?��?)��X�*x{T�L���T>Uh�%��Aq�t�E� O��2H)��p�A�G�,uZ����0��*T�D5w�29��[g�'p�u��?iJ~���H��
�,X�a�(�r2���������ð0�
�a<�\J� Q�'�O,٘�$�2J@���3��=01O�1��@Ԧ���柜�O�",��'�b�'Xh�YE�ۻrLD����-}�ҹ(��Lfg��T>#<��d��
�6I��F9!�b ��˝;x��2oW�1�(�O?�DT,l�b����-k%�Uz�-,�D���,�O&�D;?��l��?��{��p�� ^�*a�	��<�����>���4C�8�0��U�3�J[�Ms�'TJ"=�O�,�i��߽ch.��q*�[����'VB阚"������'���'��
h����,c�)t�. 
�h��v�8���F��?QUJN:y�F,	��ΪyV��3ړt��}���L�l	���'j�Aj�8$�'�(�å'R�T�4�9ߴ�����Z,Y=���/�^�}�&_�AI��H�b�j��$� ��ɟd�'����$ڐLtX��0f
,�e��'��ӂ�W�o�����.ܤLV��!5� ���)�<��&�C����� U���Q#|W $xWhN,@�R�'~r�'	�k��'e�1���1GC�V���`�A�kt\5iS�K�{��P !]�>y
գE'9<OLa�С.�U��,R�r@�$9^��-z��[�/��0d H()l)F~"ѻ�?)Q�i�"5("�. QbEŮ��h�,pbA0ғ��O  ;1(
�	���CV�N��d�"�'WўRbl¦_�@�ՠ�$"���ag��ڴ�?1.O�H��MЦ��	�t�O���� �}��Yjw%	D+�e�BT88"�'7�㔽hO"�T>Y����-e�� pF�[�i�ά	4H7�c��D�����G&j4p�`Ne�� sb�#�(O�,��:Oh"}��"��s�^�9��'�������f�<Q���2�*EB�)�\%���g�,kJ<��jS�[<:�X��ܤe�T[����<Y���`ț6�'��W>I�����ϟ�����eG:��%�N3Z� ��X&dX��O�l�|��C#�s��.��b>�dݺ%l�yC���O���&�W���!���r��09`��~���4�h�G�T��p�sg��Jk��;�I�$tH݁q�'�6�_y�'���̖6 �:�#�<�����F��y��'�}�$�>�%�J����c̘t�T�<��b�����ҟ��ğC4�屖�͝4��ypS�䟸�	�A�dk`�ğ ��ԟ �I�u��'��H�[;� J�(�#C�������~� �}�\S��'���v �GYڰy�!_Δ��'���[��I8a{��԰H!a���$���z�NοJ�R"P�|�R�'�����O,˓],��G�I0I0U�C�͕>p�Q��T���))�����MQ�G�&�ɇ�)r*@(J��$���F��Yk���y���1%��bCTn����hѸ�y���)SD�x��n�1w��T�q@ӹ�y�JM�W!,�� �h#��r�.t��'Y~Ȃ��0K4	���0y֐U�
�'�r� �ꖇ'2(�2F�(k���S
�'-L���,L='
bH�k�'x���
�'�,$���E(11cO>#}")Q	�'v�m��,J$L�gN2U�|��T�`�X ��
k���c�-Y0Μ�ȓ�t r��z^*��I�4z�U�ȓR'.y��T0F�
u�J�r����ȓgZu���@��ꡨ@E����ȓN�����7�1�Rf�k��]��VI���BH��jL"`$,��g:�m�ȓQ䑂�S�N�|u�!!Z�d��مȓIC�	i4D5/ר����!K��ԅ�q������w[(qAq�ן :�1��H)�\� 5'��2�
֘1	0����D�S�� ���Ra%Bu�8�ȓh2t$"�O��|h�'EY��Ԅ�T-*r��r��pq�Εlu\��;��l:0'*]sP��ǃ�7� ��S�? %��BM�[2�MQWf�I��q�D"O:����E4�r !Q�#�X�"O����o�X���-�*;?6Q�2"O�a�d���Q�D��1;#�t2�"OLy�j�&�eS�̆j�C�"O��Ѳ�Z�"�@��
�sh�	�"O~���Ф"���#&�UZhب�"O�1t��;謀�Ɲ��q�C"O.䨡�Sr�d�H������"O����1Jux`j�m�>Q�Ԁ$"O(���%(n"��.ӫ\�z-�"O����aN�G�y�%��&'�NA�"O��B�ɞ� �~�� ��Ir����'��9� OJ���@��\�:��"Ǧ��&����� VR��ē*�.\҂'��nA|��,M>�n��>I��q�U�tA�x�����G�,��K�?���ck �p<	�&Q�W���y��� ��/8���cK�I�m�A��Ϭ����|V���p��6X���:�g}�'p�`�2���/k������$U�V���/�F��q� F$�'@J,sr�4>H�Aa�@���TlZ�%�.}���u��*tj�q8�Z$�9WZ��'昜3��fhQ����u�E؟�;&�!���;t�N)s4�����o�3���\K@E�FG^�q����w��:��?nI�b�W���Te�Q�#�\���4h�z�ٵ�Z5��zf�}�)�	�#n����V�n�Ы�N��ÓE�����Jc|z��a�p��"�n�X�a�I\���l�/� 9!f��Q�v��@�I!hK��s����.d�,�6��|Y�q
C�l�I�kx8	����>Q8�؁$�r�O��TO϶}t����%}�"شW��2��u��໠�R��p<頇�=Y�!�@�B�dS��I�J�җ�2�?)��P�U'>]Z\w��'� �p��e�%85ID�jbł��,�p?�ݻI�R,1�H�	
��P��7Q!�@$�07b�U
����HE.q{� p����J|��X�e�:�FɏQ�P�GI�W�,i�I�&�n�X��
ʼ��	9.-���ѩ��8�X$υPA���V*Y��RԄ��r�*�g}��U�bI�@ӈu�R��@L��$��Qk �Be��h�B� �b,ڧ& 4i#&�� ^����\f�Jm�-Dd�Y�����)ǤGiX�t�$���l�pk�H9B3V`q��Y��Z��.�V��dS��u� ����'�v�禩K&_�Y�N	B���Rf�����t��� ��=�]�y�B��q��y�.U�5�'�"��g.U�o���I��$�N��yi�3)��9��}ڇ�ߢ*<�76O�����@u����ɝ10N̉�^T�`�'^�6l�uI%��4;-������K�y���@��	֎]�n)b�՝z(8i��[��@�VK��*���[�=?����}�(93.�-��uISk��<�W-��7�¸�I�~��@����$&�	�99Ҩ�'D$b�!_��F�˕�'v!�G��)*�ɳ/@*0����E�D�H伐��û|{� '�h�x��'�*����'D*�Ha"F@��E��˖F�	�@����gJD���.��Sb<�+�@R�Q`���$��yO���b�\��:Kv6�QF�#L�Xa"aJr�Q�Ph� CfFE�C�[����tO	�)L� ����.��d��k�% N7�H ڒ5�TU� �b� iI�LB�-�2���'P'PLoZB�*�x��EHi�u�B
 7W�f�X�I�(����0+7L=�ƺi�T���~R�F*+��!�HV�o-�ia��I#
h��2r}iE#v�P�Xw�V�G�	"d�(I�e⋋N�@�V��T!@҇�����`d�:@qт�# @���yJ|
��L) ��D���Ӻw��9�v�Ҙp�ȕ�`^�,>����U��A��v�"0�ד (=��!E5.��@�O���'!�����]�ip�R�$�:�s�KRz��WC	��xR��l�Hh��"O-5�$���.ِM�t8C I��iO��irT�*�d�o�c 4�Q����f���S�嘔q�΁���;��2�'�/k��s a�� �p��q�� �0<Yw�#IS|$��\�?l(×�ЗM�F�P���?K dce+�}�=� �>���F,{�xyZw#`)��`��e�qO@��ĬC�&�C��_��P��, ���>��p��2�t�����'Ѭ�qvۅ4<��	8�3�>'G�\J��K�P�����#^��=
�j��dD@��冊-=�=�`΃@,f9�DN��(OD���H1C"wr��vOL�!�2���*�O2���کT�d=����+�n��dm^�5�-�t�8�	���2X�mS�?]#�@^�V�VR�I	��IN�~u\c�#�s�I;&$ńD�E� �P�z����a�f���$��9���� �;=s���!c6}��Q67���y���P\ZM׼,p㞘@�M=O��F!\z����	_�� �J�!�¤㤏��, 
���|�ydEA������ � a���F�T�l�ЕY�oS�J�J���)�JT�b�'�P͚���A���i%H�u�`Ј�ŌY�����
�т�	�<p@���*�g�? ���恌�AͰ4Jԏ˞k��'��uZ�(��-u`H���/� ��vk�%C�< ���M`�S]~챀h��'� ��S�Ovn໲țv�8�;��
#1��@�d
)"��#<!AL�lp�sJ�U�b�A�B9�T�)z��3q	�<7����5b��JE��I3���3w@H�ȪXw&�(H���lzqO��D�UU���Ћ�s5�h��X� ���SQ͋L=H�2Sk��[���y��8i?R8�[wܬ\�܃
$��[qcU��0�����<�DJ˘U�Vt��	#T�:A��2IA ]y�7M�� �qA#�N�C�&)
�#�\�4�h��~�I�+��IP����83#m�@�8ݰ=A���4hc����-�*�C���8���+SVH�n�3�2O����˚rU`���F_���d�U�0���zVd�=݊��q�M:���&c3�I�;���p�I�qp�u)&Fׅvi�O~���S�K�6�22�Zհ�O*}e$�Ҵ�e��aˁ!çe	�㞨�$�5(S�X�)Ƶy�,c%ő��RX�6͑�b]9�O���T?c���.�W�� cH^�#uȄ3�-�� n��Su��+p��:ۓ�*��D�,Kw���$��82�h�T���G��H�Ӻ�K~B!'Sd8����$y�%f�¥��=��,��$@�Q��R>&r���@�-*
$ذG��0U�D(���Dh�D)��OI�e�Fi��-,��pj"��{��	���	U�r��DŎ�l$ǡ����L�/L�V��韆9�'��3 ��y#l��Z�|�b�=�(3����)��<�(��|��x c怪4����4#��N�����'r��H'�	��)�S�y��m�f@��Iȧ�}������y�f	�}H�+lO�	H4�����*K��"�HQ|y�o�L�-ׂ�º	X>G���T>�	�s�����N�.��d�"��6����Ā�L�$y�NPgP�(˄++��0�#ɿ �JTٗ`¼j�M��J�,c���	ĠT�=�&�%>���h�_5��i���!J`h�LC1��'�Z,�T��=h~�*7�O�����b�)6g��qS�B 3�Hz �@��j�	v���sW�R T��Iz$�@F��O�D9T�ŎxY�d�p�^�Gg&\PU�^�Z튓MZ����>�~RQ<����̬Q�0�kɻKs��Kُ����o@;���0O0�p<�gؤ+0�X:Q�.3U$���æ�pV:�J0�a��D�S��&��z�1YU(���%G��XwHW/|�0��Q�2<O��Zs@G<0�ͻq=�4"����r�u�Q
���d��
��ވ{�q:$e̚Z�
0駸O!bY��6(v��y����8�ы}"c�	��a�۞[Q>E:Ċ�K,�*5��o):��S I�$��5̃��~�a��B����3x����>QGҀq�������x�H��_5� CD]�<�.˓>�>%ӯ��h���̈́����sh^�l��5��j\�mz�]x�4t�F(�p<���N;Tt,���l����̦�k�����0�]p?�Ý���LU�å�z�����m�� 0���
���"���0=yC�׊I�;,~��0���9T��S�߇%���O+��'-�!Jc�^	W�,�ɸ2}>�*�U?�Q$(�* z��h��1E��+dA;>,ii�@@���i!)�=���'����ߔU���`Q�\:����M_��la	�O�4�CdM>j���'�|���g~��%�b	���˕8�(��c�g�X�Y$��ix�]��+�j�F�rJ>�g?���>���A�ƣW%ج{�	F_^���_;[<|8ъܘc`e��'ǔ���/ɵg�<`��k�,1�LQqDI���P��MS�'ɮ<�Xv��Ag��'B�6��,U�xԡ '���M	�h�T��A.lO|)c���C>�S�Ă%!�dU��L�a��)_��M� �O4}�O�Y(�i� �F�`e��uh�����&Q��x�r��J��[c��\�'c�=� �9O���VӐ;�l��'ˊ��e��7e�(�6@ӱw����� �~�xS��AC�x���K���a��eg(�2���dx��1��o�{�d�@��m��Y�>��ܙ �:@�0lᴎ=Q�' ��O\
)	���ڢ)��
Q�p����� 麌R�!��Ho����G8� 8�`�!z5v�3�
ϊ \�a��f�c���Sk�c*�
��
�Ki���dT2J ]K��,͜*b��0��]J���ȫCRͪ�'�FE`a��%����.�*	[�]�I��Ԥ2�$�ٴ�]�?�(	�)eH�%���ATFDb��XҦ9Q2$�pT������.YGay�lX.Y`�1��!:����CK� ��h�Ɩ6dk�-�"���f���쀤)�I4��"LBJHj�T�D�i�Ά$�,�3?�Si�lj��؁ӍiP��N:��ˢnX�]H0�j���;l$!��a�(�X@ ��'�����(��PA� �6b�ȕ`bD�':�P��dd'@��M ЄE+B��y�%�'�0� ��	A� ��A�y�F�E�H�p�d ~���Oh���CB+�2vb(i��~�X��D�:j�Õƅ�$�������p=q�"Ye� c���f1���� ��m{`L�':n��'0�Q�`�g����g]�8��L@C�-u˦r��/Y�V4��%T�
 ��aسjK|�K#�S��""<	�HM�Z�&B��Ӑ'U��2�NO�D��d�%hC#�~Q �Q�"�Ω�1�"4.�b��R���k4�:}#@@*F�JFInp"�!��OB�)���/=@4�����	��'�2Y|���T��������R�k��^�P�7����w� ���h��(q�p3F�  ���mL6��䈱�
[8��)t�aPN���h����C ¾O`A[���e����h�O"��!�N��
H���A$ʮ"�H�nńyd@�DJ@~Wr�&��d*�z��ϵ?���&��Հ ��P��>0+p��V�M�P%�ܚs�'���A7
�/���Hբǿ$�R��.c�����\������K
�K���"�	�;Ӡ�`�.̡j-��d�I�v�I�A.(7��@��HM�]J(����"4����9����[�nB�����Y1�
�Y�G�>�� �?hh������E��g~�a��\�~ȫ�K6d`ʽҤ�T�V��Yɡ���.�eA���N�*!i��n��a�Z�?��#rd�
�݅�%*�:$�p��	�����u��\�t�[�j�n�Ǔb��+��є���/�C��)b	˜F�
m��M,5�2�5���|*���t�ő�A6f�a�/����K8o�jسu�ǖ 謝��'6N������¦�>p`ʌ�`�V�%��`,mZT��D.�IH�eă[����ڶ%��PI���OF=�����5�aѻs��`���!���7h��C�
���G�u���D�3w�13!
,Đ����`(J�1�']W�P��I<�O�<(���L	̽�ы��K8�=0&��GF�\{T[V�y�)�ħL/f�۠�Xn���p��f1�$��N��䘄�|&���Os���&�:3���DF}���R=����ȓ������7$��a��V�=�u���bP���0;i@����Y�'��<�ȓ-R��C�l��7����d��0E�J���a�B�p�� �)LnH���4�p��j�R�`Y�K�dp0�5VԆȓ1�n� A�F�!��Ȣ/G+�����B����!+��s��3���1fa܀��8-Č1�mͰ)x3C�Q�F���4�1�.:�ܤ�'k�4ux���Q��l��Պ`�. ��(@�JU�l�ȓ)I�\�&� �w�d� j�%'Ѭ$���2������bJ��M��9��<�ȓj�䐄f��w��-�E�A����~삤!�dʒ��GD�+[��=�ȓC|���C��� �� �ʪ@�n!��IBBi@MI�R�%R&$��O!���ȓFH<���!P��ձ%�@�x �ȓ_����X�jy�e!BI��bŅȓW�*&��4`Ġ�BJ��+��Ȇ�wJ�+R��`d�$ D�1�b<�� 584��#�6���@"�֘B&Ԅ�ϸTҢ)�gۄ��m�]G����{~����^�E������	P�����8�T}�R@"e�p!
w���|l���ȓ� ��h��N�
2�˒!���ȓR���f���G���p.Ä�6�ȓA��RP`�#��1Ӆ�,T�6�ȓ+AdY��A�R���W�)cG�M��h�P%#�-*�52%@Z�ga�H�ȓl�6�g�/3�
�S�9񮼅ȓW��	�S�'�ى��,4�х�sc@����U�J��1
�]�l��� ܐsL�b-��]Wٲ̇ȓMβ�"IĤ;!�ɐ����u��OH6�ʤ���N0U(S��{�NE��A\��SJ3YXD��B���H�ȓ֪��E�#ܞ�2NֺZgY��m��A��_�~y:	*�	�7[{v%�ȓs�������4����Μ�9(����(RA��i
��!�䔅�9>��c�M�T��!x"a� y�8�ȓ ��Z�F
�, ���i[��ȓ�hY��e�E�ȍ�䌵\?�M��8�}��G[�5f��7F�,H�ȓ-U����G	 Fࣖ�f��ȓ;9�X5&��(}h�����jr���ȓs
\�rE��'�V��&����݅ȓ2�rY��F�'����bL�X����EXxe��n-t�5�R7�:هȓ{4�����,�f��2Ӓ>�",��S�? �]�CgG���ЌO�UCʄ8�"O����з{XЙYgK϶
)4�7"O%��m���VJ��������g"Of�`�[8	��ܪ���R%��"OB- a� �s,B�g��{��R�"Oz��2���P��P6S��p"O�}��M�T) 	T�wۤEZ "O��a�M j���R7�J v�|:�"O^q�Gkۯvn��{5���-�*��`"O��Q��<����Ͷ�@�f"O�(sM��'�<!T��#6�&��"O��3��!�v̀�eʋ�Y�"O*U&��,���8]\�y��*9D���!J�SH8���mv�p�e*D�t���Ǝ+���r��q�rP�H)D�< ��D�w\0�LՁ8E�q�G<D��"#b�_��L
#L��i�6�j!l8D�L[���o��h˴܀��Ac (+D�,{qL�]�)��M�*
N(��)D�8""ǋ��R=Q���Cڅ��+D�4B��ɗ>��Y��S
��9`'%D�he+�*�:!�ԅ�j��cGI#D��Ǡ�+!`:��N*q-��bd=D�PP��̲!A���+W-.�
]�A7D�X�D*�l���kR����:�9D��ѳ�E��iIa �Gb0���8D� h5�-_��ٴ@@#nz��@4@(D�ّ�D2,Ru�Í*<�)#�n*D��`S_C��Y�3� �R�R��'D��z��V�B5��,�'>a�fc!D���!��|`)��ݴ5�J�g�:�I@؞�S���=��(@����4�Tm8D�(�TD���iT��z��ݩqK7D�p�A.�.O���Q%tu���7D����K���4�ɳt�:�bOu�\E{��)�$H|bw!E�\Bڵ��](Xk!��S�O�tK� J*N3�)⧢۝X!�$	P{rX�σ�D�����ˁMU!�d�X�R��$Kj!�j�#Xf���"O qk�.���~aPéV8w�����IV�O�0p&��<$�4z��%ߞ�x	�'�f)��J�C�(����+S��S	�'���P�GĔJ����g�Z�!�̽{�}��)�IF�@�f�I础�����е>+!�A�*��d �/L�<t(�`�s)!�Q!��!YW�]��y�f-���!���=��ySUf�5c��X`�[{!�$.Edy��ڋZG�)T鍐)!��ӀUg���ed;<3��Y�� �-$!�$6!YމK�$�-J,Xm�ea�6O,��QK�7Mz��K<z5V\��"Oj-[ӭD�s-��K1 -sİ11"O�m��Դl�j��Ǻ |�� "OF���nьl�xb&kS�E�V�R��ItX��Ѳ��R�E�>rJ��
Ў(D�t���1,�rʔ¢.Xj�i(D��R��Y#Kc�W� �����uP���$�<���,������>2�j9 ֤��<)	�]��j��m��M��'��N�䑆�K��J�n�56�h�)�HW�c����?�a�ƾ^�����#ۙS
h�a�!�]�<Y&.��R �	0�K�+ZĀɡ�FE�<y��V�*S����Aۿ>Q��c�[}r�'0]��	1(�u��M'k`x����  I�d��z2�ܚ���~ˌ���"O@���o�%�vE[�hʽ��t�D"Oa�E��HnX����"�L���"O��"��ҽ�ы�}y������s�dI�
�r^:��׃I�O��|CE#9D��q'i[<W5*���dTq��H26D�d�(_��8�P���?�4'D�x%f�;8�����EH�TE�� &D�  �K P�b���.�=N|��&D���5��}:Pa1�舚Sh��2#D�x	©�j���%��*�FQx��%D����O̬l� qed&��A(�/D�(���I�iW�$��M�*Q&�m`�)D�cb�ǖ}�2� ��H�G���	��2D���r`Y,9Gv!���1���>1
��|��."&�R�	3�΄x�#�U�<q� �(x��8��MҲ@�8a�gi�w�<�яF�f���#Dl�1+��,%mp����^�E��s���̻(��ȓ����"j̕"�0�2bi�3>к,�ȓ=��\�E胿0s�P�';h*���ȓ����J� yK��GIן�F���bɈ`�& �OL""tɜ ^�ڝ��nO�H����:*`�pGF�q������E��-q����m�;�Fy��'U~e���4� �%��uaL`	�'� A�פ͗&�L�H�a�2x��h�'7�1p���-(R���� q!�J�'��e���r�J��g��_y�5��4�hO?7��:�"��	G�`bh�8l!�1Au�x���78����&
���'Zr�AŌO�z��ѓs�  =��+�'e��g�X�`�EI�BW�M%`C	�'��q�@�?�MX��>Eڒt"	�'O��0�+3Vmu
Uj�$C�H��'Y���W��/�"xXt@�+fK��
�'<��`��8]hhJ�g�h1N��'960�Ԫ��@$��y���<`ZH�x����$(|O���Rj]��y��^�~0��"O�%�  �����d��s�^�Y�"O���IA�<�~�ׅߋu���"O�AbT��&����K6���p�"OBb��N._?6�i� �u���"c"O��Ъ.}�a0�N:r�P"O�M���D�V�LE�/��4�"O��d�[,l)�=��04�J�f"O��o�(Q��|QU��~p�,(u"O�QbNQ<������mw���"Ot���1h���"n�bg�ə�"O��@�*��B�����Q>M���"O<$�#쎕(S�勵A"5UX��"O�x��Ş�^9@FCz�Xq"O��'HM+'%��;���/P�5��"O0,��V�!$�њoѓp@�A"O<��T��&&��� 'V\E9��"O���N�!��<�ᄝ�B!P�"Ov�P�ӄV�Rܑ#� �Г�"O����@��Y#m�%ېK��1#�"O&ا
�(h~rē�c�J7Dp�"Oq�GK��mC���0L����"O�وE-�.J=Dx�@$�0����"O�Рb`�@o�)3�L���4i9p"OB�c6#�a�D�� 8N6FA��"O��EΡUL�Q�J�o2�\��"O� ��)2'=.�*={0�I�X%T�3"O*�$̾t;B�����a!"O��ZI_I���PH�jh�a"O EX�F ;+�F��7
߳B��b$"O��!���$~H�� 7�ְ� �c�"Of�
u�Ե{�hS�I�.X�%�4"O�q�D&�=R��Tz4�U}MqQr"O�uc��՚oH����=d<H*�"O�J։�("�9#`+��$�5�6"O�0)M�*By�I�*G�W��� "O`�5�%1�~� PIR�-�^���"O�x���C.0��b0����ᣔ"O)B�H�>bJ&��G�G� �dP"�"O�4�r`�㪹�RKJ�ް�d"O>� D@+�Pxڧ�G>L�k�"O�5�b
ș��e��� n��a�"O����.$Jp���Cm��k�"O�q2R��&S��D�"L��`�"OԨ��#R�(�r|8䁃�O6Q��"O.��&ME�/��9����!Ó"O����7A�-�`��%�F�)�"O~��� ���U@ǎ��P��(�"O���`�A%9��a��&a�N��7"OĨ��L@�8����P�˥"OX}����@��4�RH��ؠ�"O��K1�GAR!�s��,�h۔"O6���e� g�^���'�M%��p"O��BLçz���"�A6x.�1Y"O�U��G^!��,���J�z ��"O$�����S�b�o���L1�"O� C�]�����El�"O��,�x�3���gbHcd�!�dѤ-Y\I�0(��6?H��`��e�!�DS�Խv�_^�����M�!�d�z-�'I�@�����!��«v:N� �Y�$]8�g�^�!�D��?U�a�N��y��Պz�!�DU4S����09����g��9!�ŘE_��a��"v~B��ЅGJ�!�0!x~%)1m��Pv�8�Q˵L�!��7��	p!.�)[`0rb�V�P#!�$�#m�,
���<$�����!��]����fQ#����t��K!��"���*'���Bw�Ń�A�y !�$߀F-��Y��޳&Z��+cCQ�`�!�DXd� ��F�NR��HB"ۇ�!��I.X���OK|t�t�9�!�V(m�B��ã_��@��v�.Se!�d�/\ �A�IXO�lyTϏ�VU!�D��Ҍ+2d��I�q(�.�?K!�
Vx�h��i��[Ƭ��ƌN�O!�$;�i�b���K�?W��i�'��E��B� ����G�]Ŵ���'����:!vZ �D@+Y�'9��[1��%�2��2�S���	�'5���q�[�0�Ң���YJ���'�fkw��QM�����L����'�d�⇞�5�F��v�C:=�T(�'6YQb�S)x��@k��"
t8��'Tp�!IݸlpE��HM?fl�	�'��00��)�T�W�rlt܈
�'p �ӣ� s{��#I�Tw���	�'�D!fK��V���f�[���	�'l�[��Mv�L� i�t�	��� f�R�̛"���!��S|�n�"O:yCA��[,0�{��@���ܰ�"Oҡn+��d�#��j����"O�����θO'�H&N�1�-��"O�<YB���V7VH:Q'n|���"O�x�ׄ��!pdd�7-ʥu�v)R"O���f�->�y9�N?A�賖"O�(Z�BT'1�X����R�]{"O�`a�Z�b�`5a��Ңi����"O��`6	L�-$t@1ė&�J�"O�����_�.H3���\�ᱲ"ON8zPF����UMԸ}�4��"OL1Y'��aȄm�Ќ�$\R��"O��1 �=�m�2��.C��%"Ol�q�h���zt�Q�ֆu$4\c�"OƜC�%�&CږA��&S�t~��J "O(a{�ؓ/�x`�Y=
Ӧ���"O�!%i�o�%�$C�}-H�34"OP�ʤ�Ůf~�bB��R7���4"OF5j�K
�Y�9˶�7b���C"O�4��±Iru�p��?���"O����$xN�d���ع�*�!"O�]zEϳvL�%���__���w"Or�8E�7I���Rf�̍#D���G܇S]�uX��J�q#�bTJ#D���㝛	��u9��гR*�[]�C�I*;�2��"�IB<�Qb�ll�C�I>L��XV�E�Mud��g��R=�C�"�Z��d䘛gj�[��rVB䉋OF5�������Q J�`��C�I���P�`�ɇ.�������C�T����L2#S�tI��?n��B�	.E� ��*J%_��� �#|�bC�I�G%2iu!�+K�1:�*�8B�I+Z�R�8�� }�����-���C�ɇFbę�4��`�(�y��Ψ[��C�		T�BWF%G0d<�s�X= ��qk�'�1*SE� 7��5�S,�y�>���'�(�ie��1��fN�m޴�r�'42Y�F�A���j��*q2b�@�'����`@"E�f���	[x��1�'�.�q��
>X���1�;�'F��ز��$b'��sn��'AK�'��M�%�H��i�2M��%B8�+�'u��t�	!L�m�Ř�% � �'y�q4�>E�<H����[��'�2�P�@	��\	�f9	�'\"��!�(�b�y�DB��s�'��aY��$XF���S1 �a�']T�I�?�"�k�AյKbb��
�'0��A �p���BP�@K�B
�':������jl�
���5�ĥ�	�'l��Sw���B�t]��_ ;,,YX	�'N�郶�:2�\E�3cNhO��H
�'�fj�G�6v�Y�R	�d*��	�'qF�Z���&k$0�"�����'�^��$���0H�BEI�|ԩ�'� �H!'W'`1�@��<�q)�'����O�yZ�t�Q�zN�8
�'���{`�G�
��F�Ct��m�
�'`b��Р¥��L��:o �
�'H�P�c�/r�ڄS���10��i�'�ܰ0��& g�ٓ���5��'�~�A�)Q�&G�8eQ8����� ��[v�@�ِ�^>V+ڸ��"O~�Y0�̀A��=X�	�,2]Ң"O�h�qeڪ�'T�zT�P�"O����oW%H�
�����N�r��W"O�qK����6|ʹ"�dΖ5���)�"O��pg��P���1���Y���r�"O�-�5���� �B��&@��r&"O����B@	I�ܢ��C�a �0�w"Or�K�o^�k���B�Aۙ
�]��"OƠ+���g��;��;��	�"O�p�pNҡd��<0`Y�W�>���"Oшa	H�)��B�ý5x��x"O�Ѫ�Lߺ%�2i����	QZ��C#"OR�1��0���j�%3>���"Op ���$D�b���[�_�J�A�"O�8��iPIu�%��	�V1'"O�$e�4GOrdB&)ȁ"�"O��K��WFn�Z���/O? L��"O�]�sZui�|:v��=��-a"O(�˖e�޴�b�T���"O��j�u5�h[p!�?XxJ�;g"O��e��oCn�r�O)]b"�b""O�� ��ѾQ� ��5d�nSzP��"O�/83�H�	���7AH���"Ol�#mJ�)b]p�2O�yq!"O�=" #��V�J[�a�r	�l�<Y�ɺ�&�3�LK���J��g�<I���F&�Hp�m7�L��^�<�Rԃj�v�!�e�;m��Q�k�Y�<q�;_�q "a�4cČ)�LR�<�U-L%0V��s��V�QF��r�P�<ᰋgm*����֔6�2��"��t�<�`�Gk�$�׎��'�R��!hFt�<Y� �"unTr�L߶p(��a�Cs�<��L@�<%��$��<���)�g�<�-,�Xp���F47��� �M�<�u��m̖`G�î~��| #ÜT�<�0�߄#��[�&��:#��!2/T�<�%)�~����;p9t�N�<ѐP)&1
1b�<p���{
M�<�%GV�8���ĩO��VSS�G�<����j8p�#Š�	K� �i�<!'�U��ؔócC�D���B�b�c�<��Eңzp�M���1vEҘ�D�`�<�eP����Q��.#�֜���^�<�s��52$���-!O�*�eZX�<y��I���`��AU�g�XqpF��m�<�o	�4��=���R�bl�J�	�j�<)�nX9K�h0�Le�H���i�b�<�����HT��C 9�C��a�<!â���"fc�2��Y3�Ʌg�<�M��c� 5��M�}��dJ��Ab�<���� %LYA#��0c���\Q�!��̨ޒ%9�
�8\�a��&9�!��)y�9ە�?P�(H�O��!��M®h�t`�P=J��Œ9K�!�d�1;�9���\�f�Cfkԑh�!��ȱ���G�H��t���ѕA�!��������V�%�d���S�!�j%0�8h
��hL��P$;�!���%�fȫңM���s�EM/|j!�DP:�����%s튡�֮EN!�L1��q��>
����D�#8!�$C)���7Μ�+��{Tl+�!�� ��9!�W<%��H{�(��I4��"O� �Ȁ�y��� h�=@?�J�"OD(�֦�3Z�h�h��\%~NNez�"O���ua�J;�hp�c��"2�t��"O��S�����@�I�#d��Ȱe"O�a��Ӧ/v�t���� :�u"O�|�w	��*�R�'
���RF"OԵ٧oΕ?d��
��P�=�`y�"O��8E#Ô$\Y�"�&@��"O�݋!HS�z�fԱ��O_��Q�"O���  �j9�ԋ���,�@"OJ�&�H2!%�e�B���D=�i�b"O� �ȧcr"�(���R�����"Ol�k��M<*\y�e'����x��"O��� h41���P¬�5�>TR2"OT	Cb�Z-ij����Wh�X�c"O�4�a��5��y1JېY��T�$"O*}��4�f�H�H��5r����"OH�����)i�iq��ٜV�Xc2"O���R�]�l!⡷�)aVc�<��d����	�7�O%9llA�Gz�<i#�+���yL 1��@C	�u�<�w�I�U�=������fd:T�An�<!�a��Y���K؈]p�A0��C�<!pJ�l����&A�)tX�E�S�<Ʌ�G%_ǄY;���*6�ބ�dm�E�<�ӏC*e6��i��ŨAJ�+�Mj�<�!K�|f ����֢*#\��'f�<��(.q�[b�2I�p9"��^�<fƇ�h%s��Jh\�B
�\�<qD#Ǹ�B��� '\D*�s���\�<��a�*���Adb� @��{ra�a�<)Vg�E���Q���Ib�4XS�XG�<�Uc�"���G!��I��C�F�<���˲Ё�QF�8�+TcE�<)��U-��� ��_=T+�$~�<���;H�@�c[�2��=ʆo
z�<��[!���P��-R�R}D��D=����
0~ 5�I/b[2���{�<Z"+M�f�"i�"�(,s����H����]�3�Y�'x���ȓ6��A�P��?�4��#(0`l�ȓSN2�Җ$X�=JnT�e@�9M/�D�ȓe2����
� W^��%��=Pi�`��~V��e�
0M���ђ�#n��h�ȓ]�����aҚp'�YS,G:a�f���B�9��b�$�ح��(��F`z����0��
i�l�w랝r#
Ԇ�8�|j@Թ+������/�8 �ȓV�ѣ@���,�AN]�|��]���&ܠ��֑�l�[5U�F �ȓ|/���Ѩ�j`f��І%^p���z��A�R��(��K)چ���W���a )Á{�N�i�D!8c�i�ȓ]�
�*2�P
n� ���_�!7�T��@��%�1əO���$�� �����Z�j[f���Q��
B���dZ��7ǘ0U������~���kg�2w����Y�w
�46$�ȓ2���2�F�>��9��&d}���XH��2@G�lY^9�Ĉ2��d�ȓo�&��0�?%���d�[�MhR��ȓF�y	�l� u ��b-��|aȔ�ȓ;u�����1 �0��M	>jz���S�? n8�H�5Pډ�&�$.�̌"O�e�1�F�	�F��4%A�O��]RV"O��[�-��NZ@�����}��1;�"On�Eă6���ͣ ��5 �"O4}@FN�3�4���';���p�"O�=�!Ȕ'��uzR��: y�"O��O8a/ظ;���T|
9�"O
��� ?����Ȉ&i�Y7"O��鲃ώkC6�#'XJ�t���"O�ە�N��9���]�1�p$:"O�IyR�҇S��Q	�ț�.?� R�"O���q"�-�����B�L
!�Đv�i�S��rC�Lh+D�g
!�$�Y�F���K���
�o� 9�!�$�(�4�{u�4$�[�E�R�!�d��0�B��-޻wJtI#���J�!��N�t4��gG&#?�A�o\9'�!��O,L�,Cw��>r*��'�wz!�J	*�����/߽.��1���Py��WE�rc��/5{�0	@�y�[�T5$����\1��h���y�O9`�"(��	��4���d���y��L��>}`�`�	�N̋��ِ�yE�01�H�!���U���j��yB"M*Q)l�&`)N���t	��y"�#f��ŀ���q�t���y��V6{T�%2lҰ@�U�T!T�y���+�j9�5�:4&�Dѧm�M�<�aE^�b�L w�_X��{�y�<!1fM�E��Z�N$�:Մ�v�<����Q�*U6���_�p���p�<� N:8�B�0��*7Q�A´bm�<�s�N� ܨ��ݐ:*�u��oHk�<9�kA:X��
!"�N��`����i�<a��O?n։8�ÝaIXX�s�g�<����/N��	� �
)|��V�`�<	�iΣ.�\��cFI�	 کӢ�\�<�S�c>|�se͜�X��j���<E��B��!@�N�iKy�<�w"�&�� �g�����r�<�ŧTQ�P|�OۻY�̜(p�m�<�ףE�|]���oZ;;�hy��HP�<���Y`62E甌	�&��d�A�<	�OM�T7>�
��I�\Y"1��g�{�<�Q�I�]>���Q� �~e��e|�<��a��ҩ2��L�^Z"m�@�u�<���Z"���S4�R�\z��b֏�m�<�Fk�}����HϦ�2��L[g�<���ΔW���"���<x��@g b�<�HK�>�@S��(:��=��C�`�<y7Gܢ=�$���K��(�!Pc��Q�<Y�h�h��*�:4�.Ջ�JK�<�AV']}.�Ӕ`ָ*X`�C�J�<ٳ��3��̋ ă3C�����H�<ɢɛ�19���1O�@��G�<�� �i8 �BF�L9�h�P�YE�<!ՏO!;�:m�΀0&�m	y�<��zJ�ɺ�x�s�<���l"����^� �H} �k�C�<"!��b;*d1���W���)F�<�i�{�y�Kȷh�@�����\�<��Ý6h��!�Z���&�
t�<�Gd��n4��Q

+�:r'	p�<Q��`i�5�cJsѺ��c�^`�<� ��!�ȯq����G�RDzr"O�(0��ۼK6���E�>�<�j�"Ox�*�a��+J8mc2��|�)�"O�,;Gk��a��G��I�-+"O�y���2e��� A �:�6��"O0��P�d�AyHb�꣡F�yB(�;�4�P�%�w�6<#�D%�yR�:?����5s�����'ƃ�yBD@"|o�ѲÕ"l\1�����y�ˋ���i�#҇$����� �Py"cA�I�}h3l@	Gj�)���u�<���ЍO�Z����ԊD�&�3 PH�<Y5�HQc�,� �  D,�z"#RB�<1�OL'!�6�B�iST��Fj@�<�� 
->������װ0��t��M�}�<1 �V1x^�ܢ@�G�L�D�J�}�<�`E6���
��\%#�(	hu�O{�<��f^$Qr�cVa  �Å�J|�<0�Z�4Iji"�FɎ2H���,�y�<A���7�`���MQ	�@Yr�u�<���Y/,�̢ 㕇YF���2��H�<!���Z	���"�h�ZU��Y�<i'�#�����P���A@�GW�<�Nʳ4V�u�uB�oa�,iF�k�<���c�ݰ%F)5�eh�ʜa�<q�aS(S�����)H�x��j��#D���So���E觭�OJ���$F>D�`�D)�B�IA��A@�%F9D�xC��V�PW\@HӀ+�l��!7D��k5�	q�izpC/b�:���i3D���A)�y\M�6�;,�idh2D����6?��k0'S�Ƅ"0g=D�	r��r�^L����yf����=D��;�L(���䧖��j�B�e7D��w�FmK� ZR��)3~�v�5D�@�ǝ/Wr�� gWX���"Rj)D�L�k�3h)̉6�	�>�3b�'D����FN�	�Qg�"v�F��"8D������eFl�D�F�r)�C(D�(���M�Wp���V� �?L���);D�\��ռ�.��s��w���u�8D�,��� @<۲C�|��E���4D����NV�aH4@q1J�"���1�2D��c5Ś�c��źA�ܔy�8s�5D�H�*�o�i�B�+!����+1D�������8X���Z	+�ڄ:��3D�Ђ�B�I�@�סT}���%�<D�rqo%脑�tȑ�%��@!�;D�t�5̂48h�`�R�x��X�ӡ6D�H�ɟH��-Q�8 ��Hx7�4D���� S�4�bb���O����"1D��'&�u}�\�d��<S�^]�c$D��M
+��m����N� o,D��3A�!q�� 3BW
6��	7�7D�|{�D
�+W, �Rn�&u6d�i#D�� Wb͒_��� �o�l��L�#� D��P�ᗚ�ڵ�5陘Ab��R�*D��0Щ@�B�B��V@'���s�)D��w�ֿ5�ԡr'$�X��3D��q�?U��y�F�|�D1+g�1D��jwA"lV6��G�1*��#/D��Ðl^8q��R����B$�$3��-D�����W�2-`u�$V>t����N(D�4Є�u3|QB0�U���ə4�(D�� :�e�ĉa�D�B�hk�@ya"O����M�&p�!&h	E��2&"O�����7�xc�ƃ�%�4 �"ODp���ѽ
x�E�#&N9>Xi��"O~��`k�I��jBE��rE��"O*�� `,6S����×��xP�"OV�� �;(���B�v�(`�"OHŀv��Kڅ�#c�X{�� "O I�$.R��2�@��Q~���"O����$R�R6R�	�I�(;h�zV"O~��� r�~]��ɴI"��D"O�BBW�X0x $�ل~y��"O���SO��_08�fE3 ���"OV����P������
#�Qj�"O���Plh�2#�e�	P��!�"Oloܻ`�ȬA��1�x�7"O�(��)���qY��ǘ%�f�a�"Oj ����ހРva�(d��"O���Ɂ*w���{DJZ'M(�:�"O�(��af�aBإcU(� !"O�M�"��7�L�jgf�
IO����"OB���mŪ����Ae({d04�"O&��O������ņ�5^u �"OR�zA�֌z�<� ѱ#UL�q"O6-,X����^�?��h#Ю�ey!�$׶ETx�&�7J����m�!�� ]��J�N�=E&��A�Ӊ7�!��7�<��ǥAiYg-�F�!�DU�W7bM�נ׳44 �v�ȑ}h!�Û|�:᠀Z=<.��"�j�wz!�D�,:^f��0iF($'����F�4b!��y
|�*��[�D"���j`I��'(║��4e(0�{�A�
U�$��'Y�q	ୂ{r�`��7G|�x
�'je�S�6�����c��(
�':�A�&Q#v\}��&]K�
�'3>��Aۉk��Ȕ�P1إ(�'>D}�hB?7u��ǥ�L�lA�'�`!7�0S���ۃ�Ի\��'���@jםm���A6�R@%Pa�'ƎyْÁ5�Z�#foD�eF�	�'s=:��s��q&�� +�$\C	�'Bi���M��8kAOT ����'�p�z���<D�E���ʞ�*�K�'�й� M�'4����,�j�8
�'�@��3C�}��eB�K�2��q��'s���2��{6L<�����7�Xp��/�, C��ZBi��Iy�����  �0���R� �T��ȓ��c�-�x2PxЄ�ȏc�
�ȓn���xh�� ���K"�T1X���ȓ� �J�Y�8��㓑�؝�ȓ1��d��^u�j�@ A�3:j8��?��}!��'ǰ �fI�(Đ݇ȓ<G�A��n��8�����#3l踇�h����d�G�,gJY�FIb���t5"�E�
g�~�8dE��Z��ц�_�FA���M�.�ڐ
ސ.<D��O�[P�(l���C`M�"4X��]u����̈f�����cЏ |ņȓ�f٢`��/h#n$�W���8���oYH9	�)=k��":�a�ȓ0��wo�e0�d* �6�̈́�}�܉��bP*N��B��\%��S�? �(ˇ/P�~�=*�Ko�E9�"O��iW���N��7�(Cuȕ� "O��8�ǐMU*��ܘ��I��"Ox�*��Z�D�mVC��-)"O<i�#�ϲU$Iɑ��*��<3�"OXa�� 
�)1|͚4�HK���Z�"O�q{��3S�R��Ū��?:��b"O�$���
�3fʙ��F�99���2"OH}��¡�h(�©ŚXH�0"O`�'��x�U��-P�V��1"O�<���L�Z�@�8�M��g��y�6"OrAÃś���mQ-W	'���"O�]��S9�`��6FJ�z��5A"O�����]9f��q��G������"O� 7E۵0�ȁ`M-���"O�mYs ҏA�L����?��(h"O�幷i@@h���+x��dI�"O�r)��U�Ñ$�~)*$ȥ"OxH)E�HJ��B�
�Zk�A"O�����0��ya�fF�'Y��A"O�`sR ��:A���./K���0"O���D��5�j��e� �V�D���"OtyX��lJ�D��X=�1�s"O��%Ή6�V�����d4(�"Oz���i���Ĕ��mϨ �H"O�dJ�:s�p��fI� I��"O����K.�� &�j�����"O�sV�ɝ+Wj	�֧�W(�u{�"O�X�3�#g~H�KQ�׈^��i;�"O��Y�	J��У�
ӥ7ޢ�t"Od��7
$�e��K,����"OH�
sj�_��rW��m�����"O�����-���Q�ѐj�"O����  �'G詃�dC�_�@4�F"OL�K'F[cZ�ar3��P\�-�W"O<P"a)պ$B�C��ͰIZ��d"Os����x듮Y�MO:�s�"O�\���2(��xiA(Q�A_T�e"O��v�D�x��P��iJ�(�a"O�����J� rU����g�:�"$"O��	_opT�Y��� ��nc!�D����IiK�Oy���r���}m!��)nRJ@�e[� y��KQe;Gl!�/���p�NvĠMn��
q\!�$�OXȡS�	%=��-��͑3nJ!�$ħ}r���--APi�W� A!��0w,���f�S(B*���:�!�D��==�}b+�c'�T��d�-b�!���U�b����A�(�!�H�%�!�$��2X�ea������F�
�!�D�! ��i�@�A&�3����E�!�$�9>H"�x���!K3xm�����_!�5Q�`�:�ђa+H	�2 P�!򤞌/'r��Ai^(['��A@�ΟhY!�d��+����͌&@}+��0I!�пR��i�pm�/m)����4!�$šZ�����c�� ���S`�(!��>!�2��1�N�hD.!򤗋|�p(�5��;F�׫K�!�$;kz���Y#x�Ԙ�m+�!�d�r�D�5�����4n�!���I�
E�$f�h��y�i ?L�!�$�[VE�@-T��t]P�	/�!�Ș�"�[�f�um�\p�J�!�� ^�*��޶@J!J�BJ�?��`"O8%��GY�ndI���K.�rv"O~|���;��G�T�VB�l�2"O����:u<�|�1m�>A:���"O<��L�?XF>��EO1D-��2#"O��C!�:aY��
*$hK�"O0`���3|��*�)
&V��!3"O.��b��"�|���茚(MF�"O��-i��3%rb��Q�v?r�ȓE�j����0!�x�e-�1O����ȓ��|�TLܝ4�>�0u�D.E21��v7�$�U.�!� ���	0+_�	��F�䔑W`�����37!Ψjv�$�ȓx.�yЄҢ$�L����K9.t��>C���G��e��Jg����m�ȓVH�,:����.,�TCݾM�:��ȓI��E��/�c��#�c��.���ȓ24b)q̈\\,����%$M��U���&!߇jaX�J!O�t�I���蝋�-I�	d�z)@�]W&y�ȓ {Vw)�?ȴ�pf��nCH��X.\Ad��T&�}�	 ݊�� ;���G���z���"ܠY��T���p���
H�P"�Ç�gZ���2���oJ%:��P����6�3�'�����O�`�T8��!|�Z�'���󧊓�~�D����5pW�Պ�'�Ĩ�A��M���1�'ȬyC䌠�'j��ZF��*j��ta��l\���'N]�#㆚z��P����7��ݡ�'bTp�!|����%�>=�H��'[�z�D�U������1;7�@(�'�H�R��"1���%�Є{��8��'���A.ǁJˬE���Q�lu|ݻ�'�.�:���+JLp(;�b@ZKHe�
�'������F�rU��2GD Zݨp��'5� �1��R����c�@rJ�q�'.T�`�b+,���3�Fg��+�'�d�6�13��Hc� �c�Fx��'xx����Г1G��b��_�S8Π��'\|ɡ`���&��W��:E����'�Ԉ�Sh'$������(K~B�#�'��QX¢G�B�`!��eO2]R=��'u���-S�n0�D�%��<��'�,�s���Du�Y��w�b���'�4c����věхC�m�F��
�'��3 B�mK|p��V�zj�'�:��S�.���P慁�?�Рa�'�̋%��>r���pG#�ȩ�	�'�.�EgΌ*�xSwo	#\��[	�'�hE�����O�܌�#dl!���;V8�,��O���~�[Qh��w7!�$I�fMBt�F���;eYG�7")!��<{��%R�.C/^/�=� 	�(�!򤄜>�K��2!���ύ �!�D��` 塕�:B�.�����Z�!�D�0K�Te�a+��O�p��$$�"�!��Ö\II0���0)�a��Y'�!�D�5z��|�2�W�:J�"6B�q!�D�5�`Y`���`��\�0A\-K%!�$U8�x�Av�Ү~2q��!�2!򄇱'�5�FAxZ5	���t!��?e�n����k\u�`�ϖ~!�/LG�͉aG�c]�pS,�F�!�� �D����F|�d�V"��nV���"O�P��u�",��D-m� �U"O��Sq�u�%h�G����4D���v�$9�v��������5G2D��z�c��7%���&�>c]��	�5D���W�0�\y(���� @I4D�t9�jԜe���"��?85���$@2D���a�]1w̚8+FU���h�u1D�P�H]9@���M�H0����F2D�� �%N���ƞ� Ũ0��,D�Lb��L2��
�
�{��Ԋ0�)D�ppHO�I�lpxVE~Q�	��(D��{#�B*���� A��e��%D��8���Z��|��k��T�b��I"D��R��	�2�%�D�V�`�d6D�l����?������M�(aȅ�1D�H	��M+H��_(��bFn4D�`I��2fe�P�P��2{H�"�F?D�25j�3-��ԍ�X>�!rW=D�����/`V��6�3\�BA�p�:D�l���3�9�ᇗ�](Z�ѷ!%D��24"�A<8����H-a�b\�I#D����EΤJf��b�j�N�5�V�,D�Tꥎ�)1L�H��既L(�(t!>D��W��5� �r���+z�T-���=D�4�T�Q#[: 9���'T�*5�v'<D���`l	Y�B��pa�ء���9D���ND�ͱs � &�a�r�7D��΁�>?$�#��V+1@zj��:D��0eLͳG0@�FH�e�p�R�8D��҆HK�,>�ie���=����`�4D� �@Ǖ�>Pt�"1DA��D3��%D���ǁKpZ (���#�x��"D��"R�zxh\أ��(�ܬ���:D��� ��Y2nز���X)���S�"D�w��<��|���[�J��&b;D��ɳ�޹jD�
��?%��P)&D�dr�I^2,B�Is'�
�T䁂D8D���׏�dG8Պ��W�"Z��J&�7D�p $�ɩJ����!G	S'���f4D���5`՘�dUyw(I�Ye|t�%�2D�L��H����0�۪Vиes=D��S�6p@qz�� ��)��e&D�� `\�D'�UړJA4'<h��@E&D��q1�s��	rO�!?|�H[A-&D����" ��rp�"jw��y4�"D�\����$����'GZx��@."D��s��qy~L�����0L��!D�h2"
���,��aoL�@<�8�?D���˧x[h��C ��DN}h�$<D� �d	��ɐH��iʯe~��� :D�,�JU���Ip-ġ<.D�PE�,D�л�g�2$xPa��z8�p=D�8)���`B�(�4��1Q&�,c��'D���g/ơU^�3�h�3`�8�*��9D���rAЭH�:X���D,EF�+B�3D�[�)у�v��%4)��Y��+D� #�����E�I@�.|h��*+D���r)Pf�"�P�8�x̓��-D��P�9A��,�b�+lSP�,D�,"�"ސ��l0f��U5ht��a,D�(������Th�K�o��=��$D�0+�J-y��=1��A�|#��QA=D�0��IV7L��1�f"5�͉��<D�� |�RW�<G03��:�Ċ�"O��X���7�Z�v�G�=��:!"O(Xq��H���3�L'a��#�"O�}Bv������0u�ǚeX,�"O��w�_!Q� �Q��O |��"O�R�S9$0��խ��H�ε�"O�ih l�0;��ܸ�{#pY�&"O�U0P�\�5�����ڪb���"On,�U"�N�,�w� �#�hH�E"O �b�G�	P��kD��)�4���"O�C�%[Fvmcԉ2g�4�8 "O��)��]�2��#�� ��]�d"Ox-���Ƣ/�dфG�<�,��"Olѡ&�JKѐi�%����"��b"O"��D��4lp&��R�
���"O���'�LWqԠ!���l%�p�&"OV!8r�� �"DK'�@2+%�YXD"Od�r�T%��xqg��D)�c"O<� Vi\�8�~�I�E�=���C "O44��&۲i�@�C.�5�Q��"Oh���K��{^�˗�3�Q"O(QjA�)?V�Q�"ٹ2ͪ]�"O(���"\�~40YAa� ���!"O>��@�\�}��H���F�Q���"O���/��U�hYs��T���1'"O��҃�+3��c�L�Gl��Y�"O�h�5�����TQ��^j�}��"O:���̐�t	��ѓA�+h�Z,Aw"O��a��M]��  ��K�|��R�"O�0�V��u��6�U�Y
�"O��2�]-�
Ѥk�?A�b��"O���,�	/4<�C|�N�@"O�����a���#&Is߈5"Oġ���ʾ-��P�-�:6~��+�"O�����n�c猛��ty`"O�mK��[�Ey�$Z"�G���,�C"O`]�c�P*J%��	G��3z����"O��*��J�K�J�Sr	�BfXXpW"O<�RF�^�.i��.U(H�H�"O6,�!�)P(1as�(]���2g"O��Q#*�6MR�� �̊[��z3"Ov8����N�5bb��( ��y�d"Oڼ�T�
Ni����f��Y�"O�h3��X	m��4j��8\Mh��"Ox��B#k� ����`@lK�"Op|y��
KFX��s� �����{{��4N7�ŁP�����"O�a���I؀,�G�Y�0���"Oq�
��B�B Os3����"O����o߃L��� �O�T"�=�'"O΍��-�~�zH2��e��P"O*���[�G�)��U�-�$�"OB�1���#��t!R#QsŐ�W"O$�cCI]��H��⒎n]��D"O��:���>��aA��X?�� �"O����f�7��j��[*p7�8��"O��JJR<�.��􉘃m؄�""O���b`��*l���)�t��0"O<�G�A�rEpE�5�V;=�x�F"OZh����1JH��0b�"<5�$"O�A��=D�~)B�AT���2"Od�+�DR?�]ƪ�1R�Y�r"O� ��đ�M�#�D_�R��"OX���"�Yy���3%� Rl��P"O� =��	9Y�dx�	"(C  ��"O(�CVdF,A~d���V4v���S"O4��1�G�Ɔ|��~�Ե�h�<�3�p�&10t-\5<��ub�\�<�sG�I��Z2�1u�a�g�W�<1����+B͐w2�tK��I�<���M�mV�YB� �D�.�{��P�<���L�F6�y%���0�(i�2A�I�<�C*�2�Q��9����U�L�<au͙�m_��bE�A�k�pI+A�T�<��J�i�����Hd���7@ID�<��!ٰC�B��#�Q��pz�ΐ{�<IӅ�vS"��5+G Z�:�H�y�<���Q�L4V�*���k�p<�q
L�<ᖎ�{w�Q�qb��|��-i Kr�<�"hC�u<^�"c�Rc)��BTG�<9�������J�%M�P`D�z�<1F�[��2�T��0��ZHԔC��M��Y���TC�hYJ����"��C�ɬij6�"CK�qW���`
ÜB�XC䉜Q(t�X� ��)��3JC�	�3�x�k��� b���rABU;�FC��8@�6��@��i�D��N� ],C�I��"@��M��	�QqCR*v �B䉩P$u�+Z5CE���F�?6�C�%?�pы�c!qa�qhC,Ϳk�4C��	l=�%
� ���$-�5�E�(�C䉴��Q��#��p��i�s	�B䉶/�R���)�N�3F+��N�B�	q�9b!�Õ1��Qୁ$K٢B�ɪ�ʸ��e�u��)�g�1x�B�	�z��I�7��a�(�c��]1]B䉕1� e���b�!F�)*�C�	�LG\H��b���0p�W�a��C�k�h��8��8:p��&9�B�	'�x�*���b$�H�3d���B�	�t@�LUjЩ�1����RB�sY���b�H�x����L�/|,�B�ɶ">0!F��-��0w(�"�zB�I�Y�D�)��9z ��hK)zB䉥5�8�$
�P���y6�D\�rB䉊]��P���B�dPbu�L@�o�TB�	�z�JĀ�<�tk���x-�B�ݖ<�T�ʴq+lS��!��B��.?� R�>@����w��B��>��bȞjI`�:�O5oL!��= iбUD�T1V���0
d!�d�4�Ȉ��I��q'-y!��T�2��4���;G�a�7�R�(s!�D�M3"�;�lE�&Ӏ9f�7aA!�D˖3�q�Eɔf����I�'2�;R��%2$J��T��;B�܃�'�"�{v��2o��d�$!��5k(��'�DKGⓌdu
�#tI�<Yk�l"�'tL����l�A{ȋW~ ���':�Y4ڪl����V�ҝU�&��'Y"��@�t���*a�K�R��0	�'jrdS��	^�J�3�f��n $��'�^a��"D�)���JO�lX6X��'Ӕ!R��uo��P��exp0��'���YPfD�;7�P�Ñ5]^ȓ�'*�b�G�6q�(A%$ѼD+�'_�ܨV�9�Θh��-"z��'�<��iиpQt@��Y�f������� ��X	��� ��2�Ԥ0�ఒ�"O�9�3j� y���sDL���X��"OS�,ӄj'�A2��-e����G"O"1�U�ևb�&��"*��6"OD�F�ӏ+�:�
�H%W�DQ��"Oj4"V��L�j�����%�j� W"O�	��2o�x�� ��|�PC�"O\����� ��wjO�`��#"O� ����11��:R�4'��I"O�ك��&3�bRg�Sy���'s�Yk$뙁J�@!:4����'�8��RD_p `Te>,�{�'ɶ���.�1	��ē3P�54"�)�'Cj�z2mG*M[@`V 88$,���'B�i��Z�u� X���C�H]��'�Z�r�QR%�5 6}�0ts�'�1��H<��)�a�+�R=�
�'d�����	v],`��͡'ErA�
�'�n]H1� �-Ԙ�悎'�^��	�'�F��'�'�z�Q����'��1 
5z�����HlFDQ�')ڤ�Ձ�:��s�s� ��'���2��f�*X9�m0o{�5I�'["��M�z%4�!��Z자��'R��Ɩ
x#����Ǉ�Q'��)�'Ap�pE�+��x kR\$��
�'����c�W�ذ����P�(�
�'3  E�?9|���T�D�����'+�-��7�90��B�v��'2�HC3̄2Oz�I%`�;�XA��'�f��cˉ�Fܴ=��d��;c��s�'���i�d �Z�(���9b
qy�'����QYb��
7@�+
�'(xѨ��R����]r A�	�'L(�yG �+z��<�$#I(Nˀ�Q�'�6��mF??�#DƆ���|�'��u��K�i����S�]�p�I��'	�53�B��3�,��x�'��	��ŋ.8�"a����0��Q��'Z�l[bĢ+HF��;+�D%��'`LKr�_�Fq �
���:S��1
�'�~�/������Gx���L͛�y�A�O��8B��<fj�e����y��U�,� dȹ3(NŸ���y*Ogb�;�,G�?���B�6�y"čX(��"�@X�;b�@��y"ƅ�).��k��4cV�@��P��y��}�����/��@f���yb��u����ŕ>z4��uʆ��y���j��Bq�Ϛ	���ˁ�ν�yrL\G�p���
��P�@�y���.o�$+RN��zV8�C�(�y�C�&3�0��E���{w�)�y2LƓ{C��DʍN�~ Z��п�y�6����r�H�����#�y���~Ṁ��5B��]x����y�j�' a�	?��(��d޼�y����c2U#��γF֌���Ԩ�y�*�+~\H�����?6֨*2���y�n�'Z[xH��[�4���qQ)�3�yrM��K~~4*�M�</ܖ���A �ybb�8��b@жO��%C�Դ�yR��	!'~�H��_�G�ͩ�K�1�yR�̯Iy%���D�9��=3�#���y
� r]�q��.P��w�]Č仓"O�,��
�{�&HRF�7p�H��2"Oh�z�)Y�G�R���� 2R�"Obe�Q��8X����	{*���P"O��b�IG2��Ep �ς4:�+"O*�� Z	�~��� �n! �"O��g��~&��eΎ>�.�K�"O(�R@��D��FM���`��"O���!�J4 ���I5eV�y"Ot=y�'�y��P!�ğGl,ӆ"O�<�רN���y�M�c�1sv"O��&��n_D���;kR�"Op��U�E5f���$�:�b"O��ئ��B�0`CR�M|Dc�"Ov@�bG�)U{�h�� :?�hi�"OdՒe���n
�qr��0Ȋ��f"O�9��
&A�j�4��)���#v"O�x��?�lS��a�d��w"O���􅌏e�p�� �@�d�
� "Oh�J�G)jҜQg�S�v|tZ"OTH�R(I<&�����f�p!�.b<-`�*=	x����ُf!�R��X�Ş��d�Jb!߿zT!�ā�9���	�fC0�� 3c�ʙ,�!��)�2��"��Q0����X:`�!��ي4t��5ƒv����C٨J!�䍭td��3�d-�raW�f!�dҵbB$Q4�_,z�"}��B�!�V�~�	�0V$l[t ,D�!�P�r�Rx��;[m�%pω�4�!�$�>}0��u��;UX��#�Y�V�!�D�0o�m8Pȃ
C@Z�rF��1!�dV C �ce�ђT��B-H)!�DA�>�,Q�kV.K��Р�Gn!��n�J���A��gB�x��F-H�!�ĉ*S@�q2	ĭo��� M�;�!���1tj�Cb�E	�RD�4 ��5�!�+H�r`:R�/�Ăf��3�!��;Y�4��r�+.��MB/3�!�D�';��iKr�K6:rq���YH!!�Mp[��JS	@�\8� �f!�!�$� Z���.J�rpI#W!�Z>V&��p�="�P`C/��s!�DQ�&{��˷J��ȑ	x�`��'�ў�}rE�1�܈aBoU�v��dc�Ɛz�<���0@��1�N�=� ����\t�'���G��lؙ|���Ȕ%�H�����y�Ǔ50<>l�A�N7����p�H��d#�D$?%?�O�*�y��
,s��u9 b׈e�,�>��$�S��;�A26FƆdI�Gա�����>٧b��U���%65\��%E�<������O���f!�^�*Q@�W7Kg�ಢ�Hhf!�U&gr�St�̻8gt�׼f�<�It�O�
��j�>j:�a�	�J?N,�
�'Ij� B�&�ֹZ�#�G��e�Or�=E��J��bd��t,�?�z�	S���y��b|!��#e�d�C��*��'��{��ԓy�4<	�]I��AC�
��yR�~�'��������A�(:p�Qd�
�t�ȓv�"8
.�M<<��l�n�a�ȓ�T)�⊩r4�ڒ�V�I'��ȓX�p8�)I�n5���- �o��|��B
��B�O��+��ʵ7��Ř�-(�,!	�^�(�Hv<dZ$��zA�0�g�]�R�v��S�? ��k�vl��1 �q��	���'�󄫟��9�bmq$��m�� t�ݫ~��Q�����x�m�g�I�T���ܑ(�HT"�|�Ey��9O
��LP
*J(�ZF�H�%Č���'�ў죴b��x�V	�w��=�8 �>?�J�H�W�i>� `Eʮ�ִ��ɜtT捸�?���IX~���j��#�(	�!�-̬7fi�t"O�e��
SO���nQ~��L���IӦ�G{�O��h�OV$O�Pq0$f_<<r�)R�'."W�J��(�� 3�D��#����=q����`!
����9��X��dT�K�!��=@>V�H"G���+1d�v�K��dc�N�
n�D����e��a� �3D��J!OÅNy̹1�Ӄjl���J|Ӽ��Px��BP+��q�^� �<}PEp�a?D�hpt�*c:qɠ�@:�X@!���?a�r|�=��Ȫ8$�]�O�,Q��x��I�<I "8r��Q�iʨX!j( ��p����'�a��B�<�8�S��ŝ*�dr�'D����kA�_�Ȥ�d�. ��p�'�����Ɛ	� �6e���@��'�"�3Sl5�(�	��+b�0�}�&�S���'\ü�b��a�0L�@OϓV����ï3�m�'Qe;�H�����U��@���>i"E�H�daD+�X`�T G͌D�riA��y"���(4hh9�nO�4>��q�¹�ē���%�)�Ӑ4	z��T.XG^u�P$�9�\C�T�D� "DO4�6�ױR��IX�����x��0@w.� ć�;�n����iFў"~n�'��$`��.n������V���t��	o8H�#ăF�O�@X�/ԓ��C��x�|�5$.a�կ6  �C�	4E$�)���oB4� ��J�RB�	�R�vM��f��N�0 ��ƺq9�C�Ɏ!s��i �F6i
��]^�C�+#C�U:`i��.�����(l�"?I���Q�
�J���萦t�ٚ"�Q�8��'����	6*�| (�AM�M��� ׫\+S�$#<�L� Ey�%-QI�����-'���_5��x�L�P!\ݢ'��U���Q�òC䲒OB��Dm�Xc��<����O �zE��lG�4�[�������B(v<�.[�y�!܉`�H���MO�?XaZ�L����>�S�O�L�b�(� ���� jƚ��'n�,�CT��Y"�]�t�8��EN�M����M���.��L�iƩ�jD�A�N�I����ȓ*I,�#�`Ѵn����/'E��]��H:�!�hMz���ِ'W;b�M�ʓX��qb���7w���2�n�Y�0B�I�;	��R�/΋y�vm���r�E{��9O����۸�ꥀa��c��p"O&�(�/Y�iU
u�a�N�>)58"Ox}�bl��v�F��7�=\yFТ�"OB)+t�ǞAM�*�Ȃ�`�n�pѕ��F{��I�2n>~P�'NAtrd�g-��l�!��UX�P�W�ؗ}��y(碗��\Yѥ�)��L���1Z�+����G�V�.D�$��(��P)��ۂ/�ݻ�K(D�,��'�P�Tk#gN��iW�)D�<��݄p~���VfZ�_�����ô��ʧ]r&���f�'Cc��r�n�]M���O��<yT�Ǥ�Q�ޖ%P� B���W�<Q�� ��yQE�(3���1�$DY�<��B?w I�ɯ9��laE��;�hO?�)� �ԃ��s�h�ْ�B�H�̐a"O�(�bd��O>��C	�&�Z�;D"O�$q�$�K�T*�B�<�fe)�"O��@4�ٯc�Ω�!G/=٦��j��x���'nz��V�'�ў����F�!S;�5���`u!öD�<�0<���$��v�0� �1!���i��Ev!�䘲0�]	M�R]��7�!�$�&R���P҂�"W�Q2gZQ!�Dye�za_?�����Q�tu ����<����k�<�뱩�q��]�� C�<�����>g ������Z�z�IAɁB�<9$�ܘ&�pɳ��M���ȱ�_h�<� eR�Nd���0��jRĨ(Bg�<i��|V��aX�AȌI���G��hO�O���yU�ǂh�a���V�|s��c�'�ʉˡ`ۻ*�D��?h��O>��'D0y���>���X�b��̒���y��=n�A{��,����r�D��'�ўb>aђE�D6�$b�-��-ה�"U�'O,�=Q�nPA:�B�f\�9��T�U@�<��J�!xi��nF�щՂyy�i���|R� �\(h���H�l�|Hz�ev�<����5i��k����J�\|ԇKp�<i�L�8b�n�C�Yy�5�s�Od���Öˇ �2k2j$��EY�>*E�a��=�[����!�Q���y*�%V
U��p���`�$�D9A&@�*�9��ikxM13��H϶���GF_�䠅�	L�)JݔP`d���"p�[q
�4 �B�"iڦ�y#�_�Jz��z�AV?#�����&�I�w�N2Q���ڔJ���,o��C�	�_�����#�#φ���Iϔm͸C䉯}�p#�DZ��zsa"�YB����1}� �2�d.=.P�2rd�K�:B�	�I���פ����qbÑ R�B��=ܸ�t/,Ri�`��ۓM{�B�7z�4�*:���� ��'܌B�ɇ?��D2G��p݌�Br�\n6C�	.q��0:�$�lt�E*��yR�C䉖�{�(L&0�o�,He�C�I^�����MֈgP����

X��B��)a�b<��C� Cݜ�k%G^*��B䉋p�4�0ખ�b[0�����C�"B�^
�B���p�n�..RMa��!D���'I�w�,���K̟L�ib�#D� #��H7$>���D��N�f4K��?D�lKAʍ�gw�X8���A�@D;e�=D����Q�Ga��9�@G�@�%�:D��' �;_jأ�b3PE���4D��ɧǜ�#(���$��sf����&>D������o]�pq��=�� �&7D��8�j2���;��B�bl
}z3�5D���SO�98*� ��@�*��K�4D���Ը����l�ږ�K�J6D� S6OZ�/�}�(�;w��M�.2D��:����8���I󆐥kv=k�B1D���v`����iϯw�N�+�h-D��Q���$�M����V��e.��݆�G���0�d�|p� fD��n=lE��"�I)�@�5yR �# ���3E���-��L�?D>��4!!D���ȓj$0U Ճ�� I*��dm֚Wú9�ȓ?�MR�Q;bkӍ������z�:��a��$��
E�A�Խ��S�? h�hE܉Lz�X�5&:�ڑ"O���@E�Ut��:#�ؙK�>c�"O��8 ��x�>��GOz���"OB�b	Т�n"�Ė2��z�"O��w��=d�� b��<Җ�ۤ�'D�Q*E��?\�P��8�S�K�rI��'�"��q/V�a����

�v��	�'����f*^,������y�ʽ��'5C���Q�ΈY�b9��u��'�(4�U

�����,,l��
�'��0R�D�>a	m�Ѕ�-n�R�'�a!�Ƒt �u���!����'�>�*��j������H4/t6���'�M�&� >.a"G��"�t��'M�Q���+2	���F�Q�VЅ �'�pM���'{��}�𢙼R�@ؒ�'ԃ�CC�I�(��/
S8.Hb
�'��3�l��ub��[��1�ڔ+	�'�:M���&���㠉�C���h
�'ؠy�PlΫ��c�ɔ.15�u��'�"���:8�@䄇>5�	:�'��H���I����kGת(頰��'��@C��>fp�;P�^�+<Ԛ
�'���ja%��t-z0�P�H#�5��'��� �bVD����F7��H	�'�
ق�J��:L{��C�0M�Q	�'�����H\��SQ�8V���'ܚ$��
�`캈;��,1ͬuY	�'���P�R\o"9S��X>[�6�0�'o��څA���싧��9S6#�'t�hڱG�.`��iAw�B3T4����'��	Y��I�+H��Ō�'NB���
�'��T�F�R�D{��8E��B08��'Q�p�<�0(��ׇR�,���'VD9Ze��pG�����M�r��'�� �(��<�)�d�38�<��'�����\3(�9 ���[І�	�yb��7��9�"�ε�6�X�̃&>���(H��_�g���X/�T���*�� �D�3'j���Ŭ�=��Y"&rLIZ�̅$��=�s	#j��-j
�VN� 4e��NF�;�� �R�a��AQļ�=�S�(`Ta�H��&�$y�BL+&�d(���C�>������$��C!
�Y8���I�|�P��&\V\��$�<�x��4_tm��4,K��+��v�X�O*�uiJ?!	�@�~sS�D?q�$�1�G4<O|cs�?s�.���ԒA4Lx���.��\�DK�$p���xP��4�b�q-��L�ZP
�.�?��PD"׎ω=�	)Lo̱1�D�x�*�JfV�jB�O\]�lJ- Ј8�)�84��$>Y�w��A�S�%�~0 ��
��x�^�:]y򱪆6��=�  �t��i���	�te�,���";������M�{~}s�f�|�V1��M�Y���Gqݑ���^�R��@[�F2���-|�i�&�ܴuqaD��+�ꌔlJ���-�W�lsb�*��ȁ����1���ִxG����E$u�a���~e�H)��ș����9��̖t�G��z�@q#��ԗ)"z,5�3�p<�mܭUS���@տMŖ�a��=NYn$�3K�&�la8�LR6vt�T�<��I��Q�,�C&�[�?2�u�O�ju 7S�yn����
MF�0%J�bE8p�N�=��'�"�ڰ �Aw�8��H�����I?�s�LB���,�L�w��y�n.C#�5	L ���(g��Z�|�Z��t��x@M-�´,��+�W!���ENC
\*pĠ�̊�:�J�;ebK�[�>��e�FϺۂ�ϮP�J���׻)j��q�Ƴ*�rj��].ش	�L'x�J,# ��#P�����[��0"���=6��j.�.3�<��ЧIEJ�3��)R�p�R��C�t�th��>7��Z�'0�8�����E��\�Wkf��bىe��2�ΨO�Qk�&�*��`�I?%�h੄i4V��ЄL�<8�����$����-^m�4ɂ]����(R=G
��L�R���C��-��;f�	��	Z���b4A�!	.���P�h��u�.D^���c�))�j�����P��,� I"'���!nq9�I�$RlH��E�T���Pǈ�%�are�Sa�NNO�'3��	d�¦="@�5;�ȑR�؊� �OC��V��4s���6O�lx��Q�jo��`��KffA8�gA�>��%֦ϸ�Ne!�-�'s���b���F�K�m6:$�c��g
�Q�5KG�f��p��LJ�%�9@�`��]�n�
��Z°Thq��b�q��f�x���kY%@H[�,!� ��0�U#I���r���D�`�cQ�I���pe�T!M���j��F�j�KaJ�S�6s%�G9`���i�M(-|� `2PS|�{�j��e�����	w4 CUe��c���!��L�-'h�@� C��Sц@�v� $�(s�	�I�<i8)G.K'IB�7NAb���s���v��dT*v�
0IF)ʿ`�g"O�Yp�|#��\M�"���8-v1���5W���D��wsܭ��"7ғU�``@t�W� HjG�&��jҍ�B�bWMd��jT3<�8�@hE�q�&T�Զ�eaU2?�2�����6tFd���@XC<�Is�n_$
�\#�D}�#?��Z�r�4eX`����X���I�\ƈ�т��#{}���0i��)�������)�����X�����<�"L"xx������;6 ����Q;8(��y@�O��Gx��?adTC�C^�syD��cD�,����F��S�ܡ*�
�jZ� \+_�@Tr�i�*G�D0���	�y��'c�ЉJ��lP�X���)Z�Zh)}Ӵ�B��r�A��R�d�����*��	�P�F�!�<Y(6�X/��8�"M}���!h�.�E,��DPi���7G4��[�kEz����Ɯ�;r�];�c�?�\���ؿg���G��A?�"=�EY���
*۹`�*]Gϖ9]�Q���� 6���{�)��w�x��c�Y4��4#�۹c�.miׯ�8X�Ec"aD;4����)p�^1Y�J'"V�{��P���O�u[����,��@�L?M���'�d��a$�G-~�ԃ$���wh8�	�B�l|��ͼH��5Z`�'��i��/{���t�8XФ�N���&ezr�ՄL�Q�D��o�9P��Z6.�5�0Q��T�H�Ɛ���G�f��ag�@+<�>A3�)ߖ(�nHp6o�r�����"��Aق�Gd��u8'��+>�4U�)ޔ,���n��$2���/�lY@���j�h��v�#p��r�W"����ϗ+j��0�nZ�,�bEp�(ݏk�n��ꄇ0�Q��,�7
��I�f��JFl�q�]��6|���{)����$!2�D}"�RK �҇J��D�d�$�=˴dyud�x��H@d	#J��A�
SI$���j�f��?��D15-
0��IC�2�Z�"�劳	��9���O��q�"T!�HOq����w$,��*�2f�eȄ�+ǀ]�y�r�Y��Z�JQ���AO�w��W��6l�Q�4E
� �{w�}�dբ���n��§_�ݮ|2'��-K鑞\BWǐ��F�k�/R�hZ �sE�W$vq�1C�x�i��E0� �N0rr�!��Q�*�X6-�aC�	3fN=��5�H��VL\�%�|!��0E�: �V��0�Rp�'��y`�Z�(hn��fB�*,�"&���ְ��F�oI��FU�q]�Y3��/$u�H3kT!�MC7N˹mJ�T�E�id�I�pY�yc"FZ-!}�X��������*s�ĬJ���R�6y�D���57=Z��
=*+�\���U�X�i#�OP�ei�Z�F��6��4����
X U��(�b�DY���U�
��$E.,���o,�mg|��'S�G�������4��&�*t,�0���/)J�p!
zi`�Ra�i�t��%�b�� �^���B�N�(y����"�>J��[5"<���^&�~H��(�	anf����G��Yk� hT�QA��P�aATo44r2���Z�0(�G��]s� h^�AQ��F
$��#dE][�#I1zU?S��1���-x� ����D�P�`b��[�8����L�?��qĂ\�|�y�� \�?�^`�'��/3/Ω�G �N�y�s.�|���"�\�}�Y�d@ݤ:�Rt�w(�>!�����`��8���������q �D���	8��i�� J�� �'��j\5 ��i!@��}o(Ѓ2�
&2�|��@�FXb���=)��|b�N�4m�,*�,��OL���ZB�*]��a�X@Q�(�Sb��h��cg|��/�$�F�1��ێG�<M8f&�b�^t12h��Va�� �M��I���_� x�j��w�L��	��p�i�h(s�� @�^�Qp��]>��nQ0��	�Ś�,�C�8�E@�J�E�X�I�oJ�Y6��#�����Χ*���� ̝�<46g���<� O�2A�ǂ�:�\�b ��'6��H��d��X�VKQ�MH�X�3u�\Y��̗o�E�4� �u�B \���eۯ���++�~4��iǘB��<[�kؒvqqO�%�e�I�=�Fe17��I=�2^���ݨ-�$wj
v*9��䜸_BX`Z�hS3t��� ס�-Dн����'W�2�?i��ѻC���Z�FM�<* ��
,
�c4�H(d����bRL~�hR�P'ʌ95D�6�eQ�r��uK�%K�L݈c P,����ЌP������ j�(��c�1	$1��ҿ�M�ܴ-Jd��/�J��d��W����$��<���d`�)H����&)n9hB�!E:��2��7cF0�
ۓrY��r&� UH�"PE "5V����]����<I?D$b�Ԉ%C&���E�9F��$��#7�H��rP�6���d}��A�iП9x<A�#�r�O|h�!N�*5���P'S!=p�6m��.>���!)6��T�R�,\X��T49D`��>R{%�Ç1!Xq�#�F�d���7z/�R1훌aL �g�>dP�W"�۰�8� ��u�гi�N�1����@�/�?/z��u��,-�B�2��3Uf�Y�$Մ�<g�H��s0O�)�������:aںO�V �H���	p�n�rAS'��`i��c`)Q?������q�νX6j��i�H@�{}�:Q��:&ЦٰR�.��4T����`�/���:'Ӯ̀"N���:��71�> !f$�TI�VK�-gZd+c+�gL��x�KT5o���"栄70�4<a�d���%4�  Q	�?y��sƊXC^|I�J��:�'a�<a��IL?�w�>r�L�k		+F~dI �i�U�ׄ��\q���&��F [�}JE�`
�5��<�V��#M�\j�J�	J@�A�O�l�0���T�`�P�����5i��$D�h��
Ief�<qN\���ȩʰz�+ˌ!��%�f΂�
���Gb�{V͝7*�	�`��!I��jU"ɣ^�U;a�T���+҄�-R-� �E߶�T�ـm�'C��rubI�\�E�U����]�n!@�I���C`� �UT��O��c�`Ԁ#���[Ђ�/ O��`3�i��20Օ@8�% � ^m���+^5;��{�,S�ȥ�L=_��yKac�=B�"���@�Ze���u+�w�jCC7�<� ѦU%uq�i�d�;rh� Pn��?I7'�hFȉ�F��(�@�f�%r�eɆd];DL�R��%@l�X��[#4��i��*Cr`b�!�
4O���$F�Թ�PoV��>xi� �l{(�9c]��|� HC�V�(�V��b0�S�F��J ���:��6-]	���AWMPuH�J� 5'i��[��'��t�Â֨ ��	!S�1"}� �m�F�D/��K��ܢF=�\I�B�5ltR��"�
��K��~���f��i(�+ZJ�P��`"��H�o2�B@��RjY�'������������{����&	\���/�P`����(F��m"���V=����BS� �0��'1R�p�
�Lu���Чs��)�Wc�N�	�L���"�N�
#��� ,
ܣ4+	�堘��BQ<���@a =I�2.
8)��c-,	���H8t碑閎��%#_YQ0P+'n}AڸO� XpLܠ}S2"?_c��M:�M� lh�X�mL2L�Z��ƍ��y"`	�� �d��l��yJW�Ohx� �,�$]�}O�3��A7q¶m��a	��=���I!w���.�5H�.lґ��9�(���,.ݢ�u�}�\�ȳ*^#E�ܲr�[,Vھ���M�I�[��}�s��sN�t��`? � v��D��1KE�J#R�4�'�F�K�O�C�T(����th���8c��d���  �d4�`N�F�� OΙ]�՘�N4�2���1m�,o$�������k�>���"y���v瘣+���vOȍM� �c�H+i}�ҢJ�h����8$r����gY�.�����o��J��;�gɫAPbLj�(՞~����fF��n�#D�F�6F���hn�؆��1CUўP�a�N�/�X�pE�:=(,b��-��*�[�ӓbR� l��"�N�.�^�`�9;&:�Xz\@EAݑM�a�2��$�(Ys���S�	�� >�Q`໴�@�'n����*��%���1Hz��]���ptz��C,ѫ�
,�7�F?�3;O\�x����w�0p��
:>�B�a�TBuv�a��S�.b� c,�X�tM>	Cl�Y�x:5�2�,局�F�2����5��&Rrx�Y�J8r�0i��lH�>���ģ��B����W�W�����d0���T�s�l}�E�?z2�A�ƣ�~�M�Wȸ� R��	�ҿ4��X�,ۜX0U �Q(���f���B	C�a�ܐ��)ޚev�P-�H����%޼=^e��藚ݔI��(I+Zi���c�+�p�y�m9ғo�"�0H5M���2 �e-��G�8��A�t�=#��F��xĸc�HڶK���C�`��c �qgͺ��9@@�E<R٫E�°O5�[U( 3P�;��I�����a٥���j���#䔒R��A�=�d�ޓU�v��u�O�/(v(� ��1M)�)u.�>Z�䜲BN��b�T�r��%+--!`K)��Tɂ�Q�|$BU����ҥâ2����9@Au�^�/S$*A��E�h�#1��r0�K�W��b����7�.�yC�U��P�ȋ"1�1S�C�2.��aU+�7T��J��!2�4�!�'�H@@7�K	J%�!G$�Y�P�#ꅆp�K��¤K�)�/F,�YuB�:h^L\
� �&���
�dS-4�37Ƃ����ab��F�P��e�ۗtj:�����"O.1dJ�X+G�(OЭ� �@%d'��Q�*�g)� �ù	GTZ��!���f��r}��������%w�� �c�
�. )PI��!A���%�&R�g^�H!rD� [�����ҏ����oK�'�8ab��;�(t�6��=9��4S�
ɖO�p��j�h�|ѳ���S��P��M>�"d�^w�� ���U�'].YHseO��u8�h����1"����l@�O�iaD��I.��� d�2o�#B2K�D�����X�7�B�p��R�,��΀�)�lsčC��@e/Si��� "ɵ�R�(aD͏W�<���#�-+��	��T�`p��a&�
C���"�НS�F�H���oȠxdX�)�
�Y%��dz����f�N�͊��6R�h\�@8�q
'}�^�s�T�.��酭�2��`��N�'9�L�eD/hRb��1� )z7醑DP@����M�93���!v�`IdeĬo]xôZ3 �:��CX^�ʖ�רw�@Xa��Yp������n�~�r��DD$ْ@K��o�T���I�t�����H� ��c!�$gC �Yׯ�2N����>	cn�4l� �a`�!}w:p�4��4���Y���.��u���N;VPE6��{��*t���@�ȯ��	�E�;o�>���g�)Β�j�/�"[9~��i/x舰�"�0"�����)O�������
8/��I	�{��Q I�-}����/�	�,���"ȏjn�`!��2��D�bၬ-����� 	���b�('/��	�of� ��
�3��@�Ba@�7�ؙ£R������e	.8���(c`ʟ-; �9��'Rh�P�c��`�8R�ª{<�(�D��Q0`|y��Z�C(}<���dVU;vt	O׍'=<����H�Kl�H��8C'�t)cǕ�L�,E �%�2p(�z�	6Jm�+������QĪUQ1E.WE�|�*�y,0�k���U��
���$Y�$(����Tθuia��SO�T���B"{)����;2���NH�_쁺d-���p<�'׹"�ne��
�ZD��2����. CIׯKr5`��*���I�*R�3�r��4'w��*H؞�&D{2�5/��T	^����9������I�O����,@n����"}�&�ˤ�Й;f��/k\�M�u��0~�-C"mA'��	Q�	�\T>�W�'��I�k��b���"Q ��-�pw/��6��Lޮ �`ۢ�N��򉘲z�L@�-�By�c�*y�Lq�e�;��s�7��x2/O�/Ҥ@�X]�Q0�HT?d�����B��e�:l��eޅR�B�S��'�B��G��exB���B�Z�p=���GB���.���fHK�P�h�x��Z�|�̹rCȟ/�xF�#i�h�sM\�E�v�K�yd�(���U����ւS5�y��BX�*aŞq8�Ḓ+&�y����;	<$�3�;eZ(Ċ��R��y��	Xp��΍Qee� *�y-;sDx\Ц!�	=�0��ͅ�y2�] ~��b���&>�>��A����y���g�B|9�J�?-K0���@	��yr��;�n�*5+�
R~88���y"�& �6|JBá^d����K��y:;�l�_."t�P��( �1�2"O�ɣ�͌�`6Y[c)4O�t�[�"O� thV��bEb��V�]&V�T|�a"O�ݘwgORd6`!�2����"O��R�Ǘ'����#l)&�)s"Oz�T�B���X��͟2`p��g"OȵQ��Ѷ.�<��S��{�E�D"O�A�a@[&m���a��V� �"Oށ9bf^�"�CE
�	�N�i�"O�Հ1kؔ:r�$�E/;y�ܕ�"O��{u��#�6�KD�	j�t���"O��;�%P6A3n\�d�A��e��"O�+��Ŧh�&a�ǀ���L��"O���p���nަ4)�j�5:��h"OP�X"��|�D�qHڱZqf�aE"OBt�/�=&М���(g2-x�"O`�3r!���f^6r�����"OD8�&bI^�� �e^�$:ұ�g"O���F°y͚�r��)ns���"O,���ʺ���0]k�"OrL��,R`���ǔ8*��1"OF	$$Y1{��@BT.�!��A%"O�ؔ�Z�cf <�H.�6h#�"O¼�7�G���,3q����i"�"OlU3��{�͙���`1jЛ�"O�H3U���,Sn�"�עh�~EB"O�{CiJ�<mX�{@����H��"O�A蠨��t*��[�,� �ZP"O�Y���U�*7��p$ȌPu
D�v"O���!��=2�T-���� �"O�hѶ�:��a)J�4�И8�"O��Ç��w�ȰtJ�+� ���"O���0�8I�"��cT�v�����"OҬ1�!-}n��C4'ʊoږ *W"O�Q�`���#��l��]�S�l�!D"O2LR�.V����ʥe/Ŵ�"O��EHiN|�i�D��ɴ4"Ob%�E��'q���BvM˝\[R�"�"O`ݺF�5��r�G%:�d��"O�!�d���&�Y׉�9����"O$TІj��C���[�GєM6�%��"O�`y�@׉X�\آ�+8��ٳ"O.ڶnݢWQ.U3Dʆ p�"O�g��@���iҭq�Z�	�h�G%���L�$:w�;2T�u+f��$�SE0���TL.��JFaD�3������Z!A����bʪea~��ؚm ����էW�`D �(ԉG����VA����� (Ǟ-�4�JEC��E�J4�w,M� a�tAw�E�̭B�Z}�G�!c�pI��
l�s�As\V��'CpJ�M�	:f�<8ǅ)}<�1�$�%f�{�ܟD�Ӄ�~zo�p�8�����QH�@ax�<�� PB	�A�@ ����m]�FA��[���!���`���"%��Pd�?˔ B(P&x	&?�_R%|ΓyR�jta��/�������&���G+W�8,2D���\�(�J|*4�ޕ�p��i�/5���2�&��
ǈF�O����-&�|}y��-s�b$�tI?ړD���� C�_�~=�P���xTs��	8���ź4E �l� 
;��]�[l��Ak�,B�	;� �l����<��2`�G2^���[怂+���s�, "|,��	�
�D����ӂ_$nX8D�]����C�)'*���B<����
7L��҂��"��)]���O����ַF�Z�@��­|� XQ	�Y�q���u��e1B�x����߇(Ǧ����*>:�Y�B�	Y4�M�,=����Cڔ}#4��͟�p�G6-�J|P�;>4�U�$)2r@
I�dĚ�5��O� �2II6qd�5�'G�O�*�Xf�~"�/�y�X��'��3ed�}�(0��Q� �Z=!r�Z3VL�I�G-��E%0 �US�'� �I���Zs���l[��}����R�D��GQIβ.�M�_wkT�K1�WCh4�Ư�:n[�ejP�ԎeHdX���T5wl.�PCI�	g�� V�N_FYc�cApT���=)�� pӔG�L>�t顇?-��`�D�H��ȗ�r�ثr�OA2E�Q�����H�}]b���R��Rv.�B|Q�@��e�[. ���Ɏ#`���pT��%^z��pmR6xı��IA4��0�����,�!G9m�l�1�8�~���<��Y����tq�ر��we�{�`�# �
��۫��5Y�g�L"2 ��Ao���K� o�(;���"��U�_ΐ4�dYq�? ��F��O��8R.����-	�e-��ĉ�"�A�!]�E���y��q�'	�=��O�2 ��AK�Ye���`ڑL�$	c�+!���Ef�s�!�6����
Xc��`7��M�n���d�?y++��\� 1�6`[9��))���^��R6	����(��B�0���'��[�ّ�Ә�*<3�Ό�v��Y��a�N2,���B�5���C�}�8 �Si�'01.AP6Ɲ6oWT��A�*"�.p�C�C����<y��l_ t�G�B+ �(|�.��e�f% ?�(��	���^ق�H &0��!�#�!��2�U�l�j\ =�&�(�� ��J��6��5��	��4]y����44����/Iɪa۵睑jQ|i#-L�]�� ��Z�_}����46��<�5o���M�E��&m+��´S��3���|��xZ�)Ӵ<P�@�۹V�j����L� �<Ysq�??Y���F�m̖��$L۹u ���e�8j5dّfLJ¾�Ga=;S���ƣoɚ�����u:ɛc%I�q����d�?fQ���ؕX�����>kJ<|���B<6¾�J/W�;�T�hF��1k��3#ˈRo���e���f.A�6��@F�p�N�hf�˰i��$J
Qh��A�M�b�=���Pr~A1����Q���I�+Ը*0�\"<�,�Ҥ"��2|��b�ˢ��}�&�.��-e������q��X���,4���Jf�a�l1'�Ho(��rs	�/a�
ĩ��w��h�޴�tݚ��S-��P��/��=����-0.a�BN���bN��dŲ���/��7큑V��3��^< t�"�͂���#�yl8��Cce�03 �$�(���v�� �K��HO($�%	��y��y �����b ��Y�d��J4䒔��.�#$<ʥ)V
��q0�.H��1:��C [�sM��b�3�oOI�d�2i�2#�Z���n&�=,���띦D��L7-�?��x���9;���Үu۶�c�-O54��c��I�*�R�M�=��P��9;�
 �4O�/w޼���W�-�(3%ƚ�IlԹ�I�L�'�2� �V�%� k�f�Lv��'IRB=|m8���$d��`���ʠ��e�� ��{2�ݐ��d��[��) ѯ�?&a��P�Ϭ�����<i׋�i0lP:B��+v�c��E�v���V�$ 'Ԍ��g<S�B�;w�j5d\R�L+(q�C��<w��
��dC��G�
�Ӡ�\�}2��p̌�2��|i��н��G@��	�΢>���[�1��t���|���gK�:?��	x���5)��ٗ`=|�`����ۂ0��l��O
����K׸:��-�D�>C|H3��Ȥl�< ����7Ov����'G$m��!Av�'�%�ҭ�&%jM0DGM"ޝ�e��:�m{��V�Ct�|��b�
X.�����Y4�pyX��
H/ĩ����8
�E# ��F�R c�"yP��Х+]
j��CZ��HO )��
��*�T��n6k��q�͐�mc��G)B�tQ;��-V
p��a�5 �`�R4.״"@��j�O28��& �U����Ofx�� �!��8�l�%sF� �R!�2#��K�$)�#noPHA������Į	�FX<�&�7�*CM�8B��0�h�Z̈	f�VĦ��rH��r�C1��DO:D��`T(^Ā��M�G/d��y�����I���H�ȃ�1~Į�K��&^�e��a��;�~)��O�,�b�H�'p6�[<\M�g�����)Ѭ�� a�E?!A�=s��h�����("?yխ	�n}���ǋ.T���Ǽvф\�&��;s��
*��cc`�c7m�4jp�v'N�Y�@!�i��Y+b-Z&�)
���]��M�!�%��E���"��Or��W��L�T�v)�a�6�Bsk� ��t g�H�9��ƪҪ7��x#��Jq��@����!j�4�J�K6!��x ��8�.Z*I��D�䩛0&v<ja�܊k�$P*�A:I �P�Z'L�t��Q��Btäa��ծ}��m��XҘ�I7'�(j�Ĉ��;0�u�U홟ur�a��&̏��ׇ�h_bACf'\�q��Ys�)u���1/	`mx� �H���2@�U�� � �5�̚�)
� �H�y���3+pM@��'��� m� �*���)&�N�Z%�_ |����&�l��Z"�ԬT�� a'ɛ^eZ���*����O�=8Fgہu�-�5!�/,�@ @VM`}�=��X���B��eװ)&'Zp�=�U//�F4 �� e~��P3) �6����/q�}���
�6�ϓ5_�0뤇{��P��߇@���1Ü���m�WM��?�a ���2�] Ю�{�ZqXpC^D������u�gu������<k܉�g�f�8,�a�ܫD�yr���g�20����(B|��&�T}&��S���>�Li��O�n��Ta�gÎ;x��㌔�;��d����U|뎏���cIN%;��	]U�G uY �Rҥ�w��,�b�C����(�$,0�����ɓ P��G={"l���]�_P�z���M	j�3�¤.����� (T�)E��L�>R�@���<k~�فDΔK,�����"�j��X���)Eb��Ǎγ?���ђ�D#w�9,m�(��7��,�R����C�K�Pg�'�v]	&j��:M�Z�� R�m��4�M���F���$���B� 9/z�Vy�W�ɡWG�-B�J�#L��Ί�V�ʵ����2]�����91���ɗ ���s�G�D��+�"�&A,�(���>�$STMԶ; H��S	��i�1CO�A�PA�ӂA&�u��#|Sv��S,�wyVS�*"��F�`��I;��'�|,Y���/��-y���t��f�Q�%���1s�pdaE���K`�O$e�^9c����P�\��7�2��Xr&�5O��B%��,�4dP�G%F�� ��V�J�ҡA}n@r��Kq���rݴ]8�I��ΏL�]yb��W�ε1�OD�|úX����vA����*O�"�F����6�~�'��	��J�Q�ZU{�nP��̭�c�^0~���,�M�N�܍��ޱ~���U��3�	��\
�y�NQ�C��cflM,�L�@C�;��'l�i��]"K�R5�'�@��L�%�A��]��,���'L�8U�07�͸ ���:nt �ŉW��(�у��� <�s��-XO�5!L0<{P]���+�:t�@lϋZ���gU5��B1>.��O+i����%�_�*���K�9T�y�ˋ'j���� k�62���{�.���d���ؙ
����� ~Qʹ��K�v}l-�`�\��7���|Eqׇ����nKzY֝� �V׺�U���v3h��2��s��@j�ߴ$)�	I�b]R+ܭs�iKTT;����F��NW�I��� ��
c���#�L��޽����Ȉ@�
P)>,�$�h�:k���`�
b���c���Ν�f�w�JA2(ҋd��p�c��p���V�>�dǭ?�8	���+mJYR�,զ逕G�%j���MI�h��������5�S��ꉺVIڊ�nXq��;�5�A�m���ȑ�ѱO� 
�"�̨����*Ej�S�A,.IҠ�A� +X���6� ��B���� $H��)Gv�c)�,.K�Q�@�6/0%H��PO���螔�\�1�� ', �{P����"�����B�-선Ӄ�^62dC�*�-d��pϋ?9<`�O����KLy^��ٴ_28|3�x���	�RE`oN�Y,����5Ip|h'�Ù~~����ݽ)^���8Rs"�ж�K/f)��g�2y���BS�\i�е�~��U�(���EʚF���Y!L�H��D�!L\"_����_�&��'<�(Z#�J=|@f1X�iԓM2��s�C"2����w��f�H=�,]�ek�Gα!-�ӂŏ�؍�'Ō��B��>~R#�-G�����J��%�,u≋7}OV��%���`���S$��P�gdZ��X0 -��z�"銴xE@���H
��H�N� X�hzS�gUI�g6w�Jh���<�!�OyZtk������ľ^�y��b�/=l��:�LX=B��9*��⳦ڨqʐI�cE�P�Y�SB,;h�'ln�`d�� }��YK#,0k��R���-r��3�M�35ʾi���].e8���MS��Sd͋{���i2.�����HY��{����|����<i��}���9�[���X���5%��P�o�qh��ʂ#9?9�̟�o��ȡ5%F��@(�v���Ř�L�YTf�a*��4UJ�1q�[.�Ђ��&s��R�y��D�p������8i�B����zm:Wh׏T~М� B'����w�`� 5gL���-J�b�)�nAZ���Qwİؐ�ޢE&����'�h�����A��T��c�5��A��(Ƌ;���p���=>̱Y�D3XT��aǝ/P���E���Z��4�c��kl��eNY��l�uK�#?��X����.P����jMU≏<�4!�@�2LQ�(�Q>i��]=�`��"voJA�IN�fϊ�;A��2/*��(0�F0h����G	�$R�b�HJ?�G�x��[z$��O�.Es��1�[?J�19G숽kl��H#LC~�'m��Pk��Bz��� �wÂ̛��J7��H�G��I2t��\�V�d9%g+�X8yR#}�R5p� b��L�������-��b��QB�ϊR�(X9�L�4K�t)���'A� �m����h[����~���n�x��Z�'D�C���'w�ԁ5����ƽ������H1&G�]\�P ˜*Y[��˓?�k��;�� ���͙1���P�ܗF�Ș��O�NzЌAΏ#
��mI!Ȍ;���D�̚0�� �D�؀3Mk�dJ�kI��s��5���
Ǔ(Ҧ=��bΗ
F>̀R*J�(F��H�
@ [���t��B�����b�4�uɊ�Mʔ	Y�Jߟ_1l�v*A�X���d�XC����E�F	`�<������AO��3��H�� ?9��ޭL1t��1��D���1Cҳ6b����:�p$ ˝@p��fH��C�0H2Y�GX�a1G+h��Q�.˂ Ɇ�TE�Dz����D��橒-M?9�0��ŗ�#̜x�l_+M���냮R�zWxə��͋�ॊ4�;:�"��G%V.Ĕx�LG��.š������O(`l�I��ӝx�����	�>��A�^�TZxQI���a�n��uI4y�8%Ev���FR�~3t�d�O:�F����
d>%��c�,M�ӯ70z�"tC�Q���UbJ�Xax�V z����Ǐ�[��z� -.X J��^�f�"r�	rf���4�������$Ȣ���gV%0`c�
�]�`�
lˈtvɨBC6p� G��X��KJSb��O<��'C
5�����~�t�R({8�PI3�Jf�$��A�!qA�����Ӝ=0�s�O�KQ`Ǥ*l*���C=����MZt8B�Ϊ�(O��#�+��ɑ�A��Z�����-42����]��1��?�R��.����@��^ə �� ,70��$�"} ��n�s��-�4h�<C������p=�䠏�W4]��GF�#��aC���-.��G%�zpf@S"�5"`����LyW(a�g�4&��ABAƌ+'����eR�2c��X����*�,� &G��Q��I67��@���9Xp@@��+%��FE�jA��ڥ �K@�)����n�XP��d)}B��x����m��R� ��I�'��8�g-Q�_�jm��E=���Q�	�lp��'9p9(�c����+��-l����'� 70����6����a>�<'��`,�h��	3V��A�u52(����S�б`caD<ܢ<�acǒU)f�r�%�@	zY2�3|<A�B�+f^H @4�F�"*��cFP$|�*v%�Dh y"_�3x��ϮT�������7'�r�X��Z"���k
�*��֜#d@�Ϝ��n�s��^`�������&��Yk��W;�`%����#dx�o5�~�S1LV[j��� �A*+j�����4�t�)Ӕn�|��M0\c��ɜ'��P�U`I����RS@
.T�2PUA�'JK�~u|�@eW�N2�����$ Bp��g��W~��4�*z0E0�i�b�ؖ(�X��	2B#ǺI̦hǓa<h�ۧ�	��()�@ݪ"���Ċ�3m}�q�F$}]�|���W8JE��"�FP��l@�煌&X�v��dDJk�'r����@�Cd�쒗��-=�U�L�h��:g\t<�d�N=>�ZH��_���S��g>���X� ��3aL�%�H�	CD����ܘuj��;a~ �
JR�ebD�ǒz���	�a[Z����&Dr8���ɟ�Q�(���+$|Ft�'<J�I7��,DT<�z���-\C�'����B�;3�=� �C�8�I��\�\#��+sH��2>8�3A4 kax℅G�.���Mzf��P���p=I�{6���tx�jS�CFN@�4 C$d<�2�l� אx�\�>���`�o	�4���7���y"��n� �ڧi�9��ɰ���+�y��̈́F5�{@A�-`|�a7�A��y�d/e�H؇ĐHa4-/)���ȓw��g��z��1�p]!o`>��dlP �S�uyj@��L�yƈ��H�*��	�D�|PÓJ�fU��ȓ,�E1'�U���2�$���S�? �\9�D(��!Q���@�mH"O�DZw�X�n�2�i[�j��mВ"O�����
tMXd8�gG49�-�"O��* �=,b�勳��,2+Af�<Q��<l���p��Ǥ>YJ��`�<!T��L���P ��!S�@`ǩWb�<V"��a��I�p*��i&�m����]�<�r�6A*�K\J��-�W�<Q��`�@�kP�K�/���qCǆk�<y�O�y�����ʒ	bz���<C�I�	G�HC�(	�@�r�H�ZK�C��g9`�1�+t��"a˔j�lC�	:X�vݓ�"M-*ZV�*P�K=H���Dߧ���
E��:74ų���-����s�a|R���'	��բj�D�(G�E2�vy�V*^�C`VD�����Orҧ���7�S�Q���ంNp2x�0O>�'��S�O;����B�%����d�8>6t�z��>�O����[=���GZ|H�����,^��	�?sj��S��-6.qO��];���<����3�U�'���3�O����mḧH��*�HN�CMzi*�@š*K���%�i���c�	o�S�O̦�UG��{S|@CG SY*���LʠXtqOjdF���|JR״ �~�r�	�?@�zX�T�W!��'�H�"��Z.i �#}:2��Z�4��厷I�eQ� ���H�aY� �Z>Q�A�*".:�!�̚$3��à>?9S�O5Hd\Ex����Қv�Vy"⥏,B��*�������Y)�"|�0�T%��vh��4b6��� ���pHE�o�S>Q��	fj6h(%��
p�R]Jt�V�@izb�XBd�6��<9�
װjV�hѱբE�I�F@� s�r�O��)�H��S N�,�bG-hDZ�<O2�I�<��O0���R���OAޠ�@��	 ��d�7f���OL\��L`�S�O�$���`�2K�D� �}����4P�Rvi>�i>-G���í9���2�?k_h�;���L�<�r���AfBR��>F]ʼ)� ن*��dQ�����=!�ɀ__a���s���(�2債`P�I"(�0እ��	�u�vԪq��9,|K�*��u��	C����a�j�)�'���$�
�a���ݩbxVAn�R��]�4L�^�)�'sD������Y`"�\� m:WdJ�>��Oi��u��Af�'Cx��0�d�q��d�c-_'O�"��ȓ6N�Yu O r~v���Fr�A��8�@�it`�\��@z�-]�t2�=��1Z8Y��m�"-��R�dؚ6sp��ȓz�J�*�
z\ܱ��3H�ȓ��µ!��\2�YE!V�b
1��B���#G��>��\a� N�!b��/�L]�6a�TB�ԛ�m�m?������y�ÓMt9��޽VW���ȓ$?̥+��P/���Zf�N�!S�|��*��Ӡh�}�|�Pt*�/�|��ȓ/|�$
c͆�`�i���0� ]��;>z a��u����E��E����ȓy'�YYu��#0�𝠔H�ZP,��}����Q�ht ��أFpx,�ȓV�x$��\�ђ��ɇ�#� lЦ�f����n�EߦЅȓ^9�٣���'=�)��Óq�"H�ȓ?*�%�R�ʡ8�l���gH'"N���8sZ#P��%{�31䎭	���ȓ't0%�m�0��P˝B�$�ȓe��A����%IT��.��@�ȓc�4H��/�
���&!T*Y�ȓXO��ї-Õ#��%v�:m�����!���Ȭ=�4,	p�	�1'݅�lDh�Xw���?�$�S�D�xU���c�8�J�BN�[r�����S�? ������/��`�p�M�"��t�4"O�����x�� B%�	s�(��"O\y+1�I5[��XŤ?uHa"�"O^����
%"���U�Im�RW"O0}! �U�Z��&�&O>1��"OH�:Eč�K,��18?X��"O��f��P���G��_;T��P"Ot�a��2]{��KE���2\��"OM��m]�k�e�A֗F� 쁱"O�ܙ$,�0�R�(�G;��� "O���M߶V�U+��Q1q�@%��"O�:`��7&].���FH�k��ѻR"O��`r�Y��8M(�OX�qӲ��"O��c�>��=�F��*�� �"O���^Z���L�Z�Z1�"O���B�(����Ɔ�\���Q#"Oޅ�E�3eȱY7&��;��E��"O��c�@�F]�WDY�0!"O�<�� Вv��y7d�o�=t"O.!��mH�z�� �U��g��Y�"O��� oظ)5�x{7��}�B<��"O�$1���v�``����N��p`"O���!c�=m��h2�<�N �c"Op���ۍBr�����3J����"O�Mk�a��*��ڐ���3�r�hQ"O� �׎(�x(��H�X����"O����-A0V� Q��gϞ{��<�"O�)�Ղ6���G��'Ie�q2�"O$�z��m������"xr4"O���@�[p�6����b��uc"O�1*��J�:�P�+��߫l}�)��"O�u���Q�E'ka�)sg���"O���RΑ�1�q���;�Y�"O�$X���^�x�9F
Ҟ8�r4a�"Oj	�K�!��-J&��z!HX	$"O�͙W�A�h"�4��W"E��"O09����F�6�	1G�1�X1S"Op��Ŧ$n�5k�E�3���)�"O�XÏ�%F&�Г��1Ro��"�"O��Ĉ��m�ְ�CԹN`�e�F"O��jf����pʡ���!A}�"O�p��'J�|A��`M�&�"O~ � ł��H�R[,�qx�"O ��b)Ƕ �Zƣ�W�`"O� �PY#/�B5�T���.���"O�p�c ��/{���D�p��QJ�"OpZ��*t�,�`J>ZW"O��30�S;P1!��q��իF*O��!���x.�=���˄Kz��
�'�8{�bE�2�<Y0C�y���
�'q\| QeF7C	�(��̝�h�H ��'o�1a��e��ђ\+�d"Um�7�y�Mߥr�lЀ��Q����y����'�VD`�1Dg� H�,
�yr�RUPY�� B�	@\��SFB��y
p��,`DMN�{���{��B.�y�Һ2�6�6���kFE�*!�D�*H�ceN�8z �v�!�DWD8�V�	|�<�3TC
�G�!��̭1�h]X��H�!��@��^(h!�E?A���YU/Kt��W�D*!�4i<q�&ͽ!��u��x!�DA7;]��d#W�5��ŋB*��0	!���%+����#^	2�p7��$a�!�� �!��"�P\��.�dغ�Х"O��D�t̠���Y�h��(�e"O�}8"[M��Y;t��0/��'"O*X{����d��C�/v�X�"Ox��HV���c�
=a�)Jq"O�����ы!��%�� _~H�hx�"O����M�� Y�.@$,�A`&"On����|p��U�1��b"O���.��lrRd����!!yF���"O���1�΀>Z���!�����U"OX���[`ޒ�P��!z�D"O���rI�3z���&�Q�ml��"O6X�7�^>\>����;x�"O�]���D�x���Sb#�*� �R�"O:�!uj�9��Xdk܂UZ��(�"O�9+6�O{��#&�W�=>b��"O<��!"�mY�J�"�!"O�mz窖�G�����
��g��d"O@��Tl�"�%�٬O�X�S&���y��4g{r0��nv�� 9k��y⥙!�fL��&˅y#6��Rb �y�G�z�y+�ŏ(�
�S�$��y�A�| >q��l-u�X�:���5�y�ȉ��4D>z�m�����y�*Ȩ,+�����B��"M �i׋�yrȞ�h�^L����1F��y��5�y�Fͅ@��h��&�AF�A��F�yr��G���R�����
��s���y"h�~�t!� ŬN^y��&�y"�̍e�� ��63��jA� �y�L^��D��@U�>a�X�SE��yB�)7��{�g�5G_Z
Ċ��y��	�g��#��	�dl
���2�y�nЦ^��Q���5hۑ�Z��yB�QDr��3(Й}�lpە�W�y")�c�x݊�m+#���a�L[)�y¬\>{�xP�����{�DC��y���->T�LCA�D;��uz�	˖�y��;dO,�y�$U=Ly���yRi�8pҀ)��U;`⡁���y"*�&}�i�w烢|s��PV�<�y��&Nr�x���r������ǣ�y�a�{MXY�a�"o�D����*�y�h�
l��(B�چj���3QD�4�y�d�Fn�be*S5W�u�pmI#�y���B�p���@�J�l�a Ɠ�yOݚ!O$�bQ-����l���yrbƯ&J�1��v��#���?�yr(	yS@t��E��fU~%H&Y��y��=%?옊����\���H��yB��f���S����AU�S�y��0Gkv		�\%xb��0���y��k�V�k⋰zU"ilͬ�y�bֆ+D���1Df¦T�����y���,7�R�p2MO�4�Z�I�dW��y�� d~��S�b�.�>�I��R��y�	�5k{n�b�/O,Z����в�y"aH�#�L�QUj�V�fa2`�
��y�GN097�鱓�P�B΀�7k�$�y2��9q0H��
6<����W
մ�y���~���u��&7D<�q)��y�B�u��dZ`&�(�&L"�d���y�i��{�M��5{~�xp���yRI�+6AH�Yd&��G�JAp����y
� ޼B'$�:AAp�N9R�)�"O  ��J�)?���*��p�"OR��&צy0��Ч��.'ƁjS"O^)��HLaxLR��*/2!�"O|��-�,F`���!��E��z "O��j��qbm)��U��`��"O\y��#�3�`-q6�Gf�H"O�3�Z#X��p��#)\���#"O����U|��C#�H�{�T��"Oڑ�ÈW�1F��0�ۥd��騒"O�ٲ�#��zI���/k�8Փ�"O��:2	��n�"�ȗ#�7tB>�!�C?u�zy1E��4~�F��c�&�!�U�b�V�K!e�	V ^a��Q�U�!�$ޡa'�#�'�2kJl�@����'S�4��·K�Z�P�32��	�'q�0Q��$5���+�8	r����'D��瑅]���I����|L�$a�'>�q�G�C5 ��mX�o�x�'��5I�ӆ��Q9�MU,jK�X��'�
�)�jBv���dg(�j	�'�)��	^�2�ʝ�F�5J�,y��'��Xjg@^	+�����b�0~�X�'���!��t�0�i�"T ���'&��rc�&`T�J��C���p)
�'�ʸ)�'�y}��5c .��Q��'
�� ��]�tG��*�)�����'���0��C��%ȇ=����'pd!!��.F�z �E ���9�'�\P��%��E��ȝ*���	�'7& Ied�+ �VQ��o!p(1	�'�p�9T"�{�	(W#S6���	�'� a�#�Q�5�.m�Sb�7��2	�'�m�7 c���J��r|�'�01"�R�1�FU�4+ =y,��'b�#ׇ�0N�ҕ�c�N7�FAZ�'�>��	Kfj��IM��,�´��'��u1n�`���#��!:0��'|���c��&(Y�bѓD����'��;��H�h0K�jɚ1td��'��s��Xx|)c4ͅ$9�d�'VN0��:G��z�C�׮��'�
  ���   
  �  A  �  U,  �7  �@  bK  W  (^  �d  �j  !q  cw  �}  �  +�  x�  ��  �  D�  ��  ˯  �  Q�  ��  >�  ��   �  ��  M�  ��  ��  ;   Z � V  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��hO�Ә<4�0���H�m��z(P2��/��ȓ��A�EX7w�,Ѡ�C�(�A�ȓO�`|�c٫f�j� en�$ҜЅ�u�j�Q�]�I�#(���!��S�<�����o�ep#��;~�x�x�U�<���O/5�B��	�|M�OM�<�&��6�
�(��F�Dd�s��l�<���+o�"�B�r�����"�p�<���B4+���R��5��ps�jUT���hO�U�!�rNUu���:�c1�����9ۄYiҪ�5D�Z����^A�ȓO&�\�d�� ��$J���+rFj���ༀ�*�)[�Thq��	�L�Х�ȓ8�X X��*VT�f��0d�Hx���q�'`<��㯉�:��Qg�C(o��MH�'��%���8�Q���z��(��'?8;f��cyd1Hv�<#��p��' �\ v�Nk;BP����0�����D�L��2�+�)���V�ܷ}�Q+*D����n�&`�X���*Bi����O�B�ɧ�:��HA�wߚmq��L�f?��Oޢ=�}R5m�=�*��R���s'�y��!�ڥw�$���"�($M���L�|+�'ўb?��e�6^0ѫ�銭�lA��!$D�L�Ǎ:�ܡ �\�z��S�$��4�O$��`�g��WI��~�|T�!�Iq�O��� Z��f҄}�.�8fFM6_ʴ��d�94����(���ࠦ�0w`jQ�t� ����<��{i�Q�p,�/t� �p�k#��B�	�uZ���''Ř7}�������>����h)@1Dz���F�m���PL�� i7
Eay2�ɂ.���t��.W�h�ctÍ+`a��'a}R���T��`!Q=Wt�)�#�L�yLM�U�H�Ў���z�2���yR�:|:�����RBG	3�y�Ʊ6���zԎY�0yp�Q��yҊ�?>��p���Z�o�����#��L���Ex��'����;;?��F[�&�#
�'�v�(tdߝ[3��#��J;X���Q	�'!:�����9[.֐��kͼ�v�S�'�y �K>q"�I:q�T>C��0���~��'�BeB��L"8Up�j�&Z�M���)ӓ��'���� �9�A�Df*�	�'oV��Cʍv�6�� Խ@�.Rڴ��$"�S�'%^f� �dL�it�Q���+G��T≩d��`˂'�-���Ґd���(��N��h��!tj`����-γg�vm�l��<!4o��.���ְQF���H}~��'��T��L�>��h�J,h�2����d���d�(��I7YIB!D�Y&!�H�s��B�ޏ�RU�_
'�	p����d,P�Ψ!QGU4{��=��+D��A��L F'���& 8iո��B����<I$�>I���?%8��� NЅS�M�O�<�$!�5��IU�ʃ#�`lK���f�<QqG�/�Z�b�%�(�ڜ�P�Qe�<W�
�=2L�`GQ&d0XE�T^�<�GB�P�䱂��>�"]AhV��d�)�Ts���/��9���@��܆�^���9Qgه;�Q����m?6,�'U�}���{N��DѡK�Jl�Ug��y��݂Uf�,��������*�yª�7@��9��*\��+��̪�yB�'g�R��d%K�	�D�
�E��y��@�`!H����!�v��Ra݃�y-V=��S��۝=�I��/���x�Ȝ�l��ٓuᜂ@�.�v��"�r�)�B�����_1�鑇�گs��E�'լ��`�]�|b�ZG��z��+�'����8^(�a� #��^-��];!��Y�M����O�
 �Z��nխ!��p^��"��l�Hs`X�b�!�d,N`9�dC��H=�[��!��2b�<k�h\����;-,R��D>�S�O�.t�a��A�"��A��gW����?鐬v�rL!�DN�W�؄��'��:��Ϝl�<QG�� ����!�K*pभ�o�'�X�D�D�ڂa*|��7�Z./o�"�9�y�.��3��A`��
0�N���Ή&��I���(��O����K���5��\��)6��X�<�� 2��cA 7t�lHgk�����sӊ$�'B�$5&�����*)�O �fH7�=��k��	q!�K�< �Z!a �����C�=��]�Df�KX�8�Oָ���W�\�h�`�� �Z=;�"O(��paO�Vi���U��t���I]�O�@T��L�(U��p�F-  �Q�'=�a+�jӃ]�,h���v�� �/Or�=E���Q	ޱ��k_�X�
ݱsɷ�HOx�=�OKh�&h_�(�|]�L˺>�I���� <�o*��H�
�Vh (�D�3�d�<E��'��!�O��zYY��h2�P�@�'�PP��e�g�́!��ʣ�ܱ��'���!�&�ve�J���I jB�y�!ͧUU����
�bȹ
�����D"�Ob�ۑ-�$
0
Ĩ�@�>R�ָ��"O|��%M �t����"�̹_��T:�"OR�
Y��pp��&���m��"OM�Rd��.µPVk�Q}��"O�kQ@�)CEF�Ô�ݰ8s�y5"O4�H���4����8j��\�!�'��^����3�6e��ZBO��xjdh���?�ьus�YYtN�2 �b���a�'�ў�'g�n	���Q��D��m�;`Ni�ȓ|��4qA��0v�2y@i�/xQ(h�ȓ%��H�f��xY��+;<�`��jՖ�ɃĂ�"�t�Sch�+J{du���8�r�7",��Vۥw��ȓ*��u���8���!G��MٰO��������P!�.tRTE�0"O�� ���/���RM�0�8��"O�|ɦ�ڟMY`��劣�������d�>%?]��EH�T�,S�ɘ_X��bA4T�|ag�� f��ieiC01Hh���>Њ>�S��	���QgX :�VmS��j�%��2$�dpb'l)�K6`ޢЅȓv.��`��fDL���jG�?��I�ȓ|[E1F��(���0֪[�5`����_'��)1����ڳ�-`�� �?����~����u/���W,N� S�ݨG.Zx�<1�.ȗt$��F�Ǳ�t�h��Ko�<�Rb٨�^��A�Ыl��0cN�k�<Q�
ߞ4��P�С}�~��S@��<i�d���x�R��"r�>p���}�<�'�؉,�6����c'l��
^�<	p(�L��0딣PF�����Sb�<���G�F��l�A��>0�p]]�<�N��C5�MR�#[�nz���'d\�<��۠w����ˢ]f(�'N�T�<����A�d�1D��[���glP�<�%��58���g�v!<��̟f�<����5J6��jTZ��;b�h�<�ӄ�$�-���A1B(+�h�<�ĦF-h���ҥF.b���B���e�<)@n�����I��E�0iv���hK\�<�DL�:��+@"�*mgz�j��W�<)Q�ǙJ�`�KĤ&��Y��S�<9�Oi>҈�(@b�8p��-�L�<�խ� H6ba(�BDh�K�<����fa�TKcG�4}�����D�<��OF'x.\�Ђ��{�f��&@{�<��	c��(+q�IO68�Sf�y�<Q7�)�z��bd�t$�ڰ�K^�<��̫,�� a'�ԝgw�eZU��V�<��nh�b\J���l�p��FCS�<q3���%�Tb5 ��"f5�էd�<!D��!t}��cR$�8f��jH�<��m��}��̻�)�3eC��B��~�<�u��<|��9#‹(�Xa�-�n�<	���-e����Q̕-=v�1!��g�<�#�U.q��@��^�j0�e�<	�%T�'�l���)+犜���d�<A�I��=�ՁS �0\�BA_�<�k.�`#�S�q{&eЦ"O� NI��=�����Ēg��MI�"O>h�/��ǚ=z!B���9�"O~eC�A�z�rD�a@�$]ex=2�"O�e�:�9{�DĲV�"�"Oj�;��[!+.�QpB3N:,����'Rb�'<��'$��'��'pB�'C���sA�%�4yņ[�*��)$�'{B�'
��'���'�2�'Z��'��p�V�'��x��q�~���'���'9��'���'s��'���'�֑�.�&ˌ��/U�d�4k����6��O����O����Oh���O��D�Oؽ�t��Y�-�M!:oPx�F��O��D�O��$�O���O���O��$�O*�ip�	|���H�RT���b�O���O(���O����O����O��D�O��j�!�#�\T��h�f2!��O�D�O���Oj���O��Od��OX�{2Fܕg�$�R�l�L@��a-�O����O@���O���O���OT�d�O�yK0�<<�zipS�X�Р�a�O���O>��OH���O��D�O��$�O��i���ffQ�3,M�H��к`��O����O����Of���OJ���O����Oʱ"���x����� Q���[�2�'^��'���'�R�'���'��
�$S�����>]�.ͫ��F2a�"�'���'���'���'��'����[u腑Jų]� ٪�,E�N���'���'���'��'7��O��Y*;��\ؔȪ�R܊b��A����'�b[�b>�Y?�6H��{�&َ	��DS��ԼU��m��Op�l�K��|Γ9ӛ&�՜(x�)���U��S��M�^7��O<�s��s�<�#�T�:wǏ�]�$�O��`z��.���*E�G�\����yR�'�	[�Oa�]k���}���	E%�8JZ���grӺ����,�S�Mϻn��9�r�2wL.�U蘬8����g��6m�֧�O�hY�5��~�cN�:F�� ��E�ӪO��扮q�:(Y��<�J�E{�O9��W((I�3'��Q��\��`S��y�P��&�P�޴!y&��<�'��t�(��0�(3�<�k��[���'���&Md���	A}+��0�YrJō��t���������K"v@8�˗�(�1��hhbwݭ��� n.�k�Ə,���J�m�-�]*O���?E��'AH�ׯ��#�PlCed��`z6H�'��6M
G��ɝ�M;��O�Ј���6��R�
ѩD�T`�'�Z7�
����	�:�\�o�{~b	�<�|�U�͌]^�cSNߥ���d�>y�R}�F�|B�'��O���'�R�'<-�R(ФY��I�R܈�1'�4��I8�McA�B�<QF�i&�����O[vC����a��$b�����O,�n�/�M�Ľi_r��������`��P��<�1��3Y؄�:d�()g��$Lh�0�m�+1��tb�Ay�	�H��QW�i�u�Vȸ��*�8Y��̂[y��'3���dQ���ش0� I�L��Q!��%��Ui�@�qBl	�
?���',�'"��6#�6jm�")nZA] 8��FR4@z�c�	P>o$�$)Eߦ��?	��O�v�B�A����$ꟾ�1ki��3��}�5A�Wð�����?����?)��?i����O�`\�a�q�.qy�����)�'f�6M�O��mZp��	T�$�|b�]:�("P���:~��OH�b��7- U}��`�.�mZ�?yP�+N���͓�?9�.�E�|��f�R�YyR�!_#]Hi
���m .�pO>��?y���?i���?�
Z�YK�-��G�'`r�s��Y��?�����BѦ=
�y�,�ٴ�?y(�h���́:D�a�.K�E�LSg���M�W�ic
6͔Z�S�?-H �ڀ20��hćџ`�Xxc���t��`��E����'=�tO�?rq��_�	�/ ��ǯ@q��*���=��	�\�I�L�)�eybIoӸmc��N0&�i�嘾K'pd+S��6N�$�զ%�IN�'��7�E46���X�Z�Y��;fƖm(�M�"˯�M{�'�bʄ�nJ9��O�]q�I7��șb��/ ��UX^�}����S�E�#B��b�Z�/��u��!&�0�����%4�Ƶ�C�Y�a��%~ps �U^~@�8�a*&��C�	>�T���Oj�)�cS6:�p#nJ !ZĔA��H/nU��!� -����c�J~�`��5`T j|0�l�w�����oD+j�Rx�O�V��P��:C�~�BF��"
ŠT
���[��\�emA!~�"��H�J���Ye���6�
 �D�J�bQ ����+x��0śK�6��Or���O~�i�U�i>�+`�����׺yA�2��b���(H�Iv��џ���?�%�8�ɱW��U==�82m&8��ܴ�?���?u)ؤ`�����'���o�D�Cʌ �zXkMS�=����?�����<���?Q�A*����Ǎ_#�ԃ�lǑ.�J�{2�i�2�(}��O�I�O4���<���ۨG�̢āI$D�6������'l��yB�'-��'���+>�q��_$'���kŪS��,��¦�ē�?Q���?�,Ox�d�ONt�G�%�=�Qk��U�&X��c�,$1O���O$�$�<�լ��U���l;ZL��+�e��)aQ@I<=��Iϟ(��˟�'<��'`����d$k��	(� ��EI�:k�ȥ��_�l�I蟄�I|y�O�5Q.���E�/>`�!01n��!�^Y�����x�I`y�	��O{ȨZt��G�x����	�^>M��4�?Y���򤖲Vk� &>��I�?��7#��t;5�μw�ĘJ��$�6�<i���?!t�XĶ�?��� \)��M�'Ts<H���<|H��i��'޴�J��`�v�$�OB�D����I�O�u���F� �h�!"*,͖5:�{}R�'�2��\�ؔ���O�nٶj��0y����d]q�睛集o��!��7M�O��d�O��៖��O���%�j��lJ%�4����a���m�
̻"O�O0���<�'��'�?!������s(�6��u)�Ŗ5v�F�'E��'0��F!`����ON��O���Μ���N�m�!�9:L�]�p�'j.4��O���O����O�=9AjV�nc��",R{�!�G�����I���۴�?q��?���<b�ST?�W�!o� ��N�2p<��n�j}bkK��y�S��	���O:�N�)�����Cb�lK���^0��.Q����'�b�'Q��~Z+O�����U������)��ha��J�u��Lw;O
�H�((��?!���?��F؂\ЛV�̷'H�ቁ��M�X��[(l�7��O��$�O`���O���?!0n��|�Y�#�<���]�Iȡ��.+�V�'���'p��'D���S�7�OJ���?<��E�O�7tϰ�x�Ǧ;L�l��h�I֟�'�(�����\��q�J5���h����{�h���`�Te��ǟ����Ģ��T��M����?����j�FH0t��ز�B�q.�� �H9B_���'��Iǟ4�� q>-'��sӘ��6"luʪVb���D�ƴ@P��'�� ^Q�7��O��D�O��)��<���$ f�� &�<o� lI��;p��e�'X��ٖ���|�O��3 ��2rG�5b��5]��mZq���iش�?i��?��'���?��|�=;%��B6:��x�+��z��6����W�(�f>&?1�S!)j�4	2��'/:�0	����q�4�?����?���E����'`�'c���u7���_:m{�R{`� &��MS����DJ�K��?��	Ɵd�ɣ_�����"���#��ĽP�`�2ߴ�?Ѱ&����Ioy��'�	�֘�*�؈���^�64�M"b<��w�����?)��?9��?)��?I�/^�%z
8�M(x�J����4M�Nؘ��i<b�'���'�����D�O�V��04��ir��)N�p���O)"	�d�O|�$�O����O��'V� ѓw�i��(��"u���zg�ox*��T�q���O���O��D�<1�t������!G�ܣ��
/�X�0vH�����	(�m�I������4��%P�Mk���?9G�@�y .��c�
gI��V�=I՛&�'R��'#���T���b>��'l�u�&˘�|X�
ы��&Q�*���b�'��I tTh)��h���O��I��Z��-��֖	J�呀i�$��'�r�'�(Ќ�O"��!���6Ȁ��<�×�_�LjJ7�O��آ���o�՟ ������?]��?*���dʻc7���l]~�R�ةO����9v����'�4���O���񬖰<�B� ���'���	ڴM�2袡�i��'��O��4�'b�'�Fԋ����%;4�Q�Ҧr��P�eӊ�1�G�O��d�<�'���?�W��$6Ƒu@۟"�6���J l��v�'���'p�z �pӬ���O����O`���J pQ�INl Ǯ�G�nD�i��'�@���)�OR���O^A����s&"E# �b��<!������I9"���b�4�?����?!�TL�SY?Y�e�&���[/p�uz� f}R[�yb�'a"�'7r�'��ӫ"��,��t�1�ڹA�8{D��M����?q���?Q R?�'��O�76je�2o��\};c��L�Ω��'���'��;s�'��'��͋	4�7�F�
���Q`��,�����R�L/�lȟ��ȟ�	��|�'#"�ѕ��ܴ� ���mefFM���.�o���h��៨�I���ɽj�,��4�?i��E}���&�#�R�BT���D�t8��iSr�'��^�H�I�zؼ������ ���d�Ώ ԋ1�׌eDp�nП�������I���5*�4�?Y��?	��:F��bŅ� [j�ɓ�>3A���i��_������������	&_��s� �9�I^�d��[`N�q3�\�з�e�i�bb?4.`6��O���O�����
��'.��Q���&��d��5"���'lb�v��'�2)����d�~��&!T'�7쓤_�H�R'��M���x���'Z��'(��O���'G��Ўs�D!S�*�QhFyc���+TX7�	)wZ��-�4�Z����d��T�biz���#{o��U�ʫB���d�O��D�OB�2�@覩���L�	П\�i��C���_�*�욆P$ވy��e��O��<O�������$:�٠{X���`�_�o��l�>�M[��j�@�K��i��'�B�'���~R鋪4�|y�PA���4�� N���$�BD�D�<���?����?��_�ĥ�����Kn����J�o�޼p���)w��f�'�b�'��/�~�(O��ĸt�*�a��I��u,h��ڳ��%���O����O<��!�	M�Vd��m��Θ�v�ԋn,���3�������4�?1���?���?y/O(�$Q&2����U�����b��L�T��
�Z��o����w�����O��D�OP�K�Ѧ��ҟ��#@_:vl1���9j$aq�&��MC���?1����$�Ot-kD?�L�����B 4�"Q"D XI�M���z�����O
��O���.X���Iß ���?��G���R$KE�ILFTC���9�M�����O �I�7����OV\8�<���D�L���b���LdF�4�ٮ�M����?y�@+
��V�'���'����O��"S�E����̆M�E�Ã�H��꓈?IA�R��?�.O�a"G6�z�O �i#�ٹ7�Ԋ��<G�nD��47�	³i���'��O��T�'�'{���4���D��`J��)��j�k��41&�O^˓g� ��'��'�"S� >�A0�4������4N\%[V�iC��';R�Mc3�Or���OF�I)'��p��F� :�c%�)g�7m4��>��?���ӟ��I(3��)�'`[�:q��8Sj�1�v�#�4�?�`E�nd�'��'�ɧ5��J�}*���̨V�މ�2����dED�$�<a���?����6���Ā!f"���+\-��h�G�Wn����0��k���4�ɕ-V���� 2��(�#� `�Tċ��
��'�'��O��(�Aj>X�A-m�v�SA@�#<~Hir'�>����?qK>���?����?���qˎAڑLYj^�b�H 83@�6�'>R�',��~��i�-i���'�nٚU�v�b%��B��X����Q��7��O��O����O ���:O2�'��j��C�E��ݹS�Ś6�d ݴ�?)����!��8'>��	�?MjvN��FH����/��C]�@���?�ē�?��H�:@̓��S�$�]�A����g�6�"8f ��Mc+O6<��I񦁉������t�'���襫�,j�Jtq�"�W�5Qߴ�?����@����S��n��`���Zf�iS�Y$bd�lZ�=�	޴�?a���?��'_'O��"*��|����5���х����7�\(g�"|
��y\4���7��2��(�B�i�i���'�Bȃ�7U�O����O�����(1[�$�6�Rh�bcϮ Ӯ7-=�dA�XU�]'>���˟��	;J7�ۗ�*_� ��pȤz����4�?��"ɣK�'�R�'�ɧ5��W�c��9�`ӰE�̃�@�;��N:��<���?I����!%�𠪠�]�*i;ÌׂM���4�j���	d��	 
1��@� �/-T�16J�8�,�*��{��'��'e�[�Z2!S��G�s� ���-H,Z^�ꧣL����O���7�$�O��G�iL$�dù\�8q!�i���B2�4XG�Y�'�b�'�2\��[���ħ<N���&"�$�#�@߱6����i�B�|2�'���H
z��>!a����l<[`&��M-W>�7m�O>�$�<��^�:��O���O�$��Q P�6Obh0R�Q5-wrD+r	<��O���V�y�)�T?��S�ط ��yХ�Q�9��Pc�n�wb�
��Ta?Y�I�6f��~��G���\��ɟ5�"H����r���ôc�h�lC�I�M�2����N� �"�s�@y�D�R/`Z�*�e?1Jl����]�vE�@%å,f��QR �o�0�y��U2n�J�&i��2�t�cB�L4M��B5(�X�>����9(�ᓅK(B��dHD,��$�-�3�*q��t+M�j�Ι*��ٰ�le���Q��(k��S�|0`�a��5#\*���������,�Ywnb�'3� ���<����"n@�"�,i1!F�$�A�3�Ņ?�ʤp������dY/�и[B�^�6B��А)40J֩�R�A/.���	�$�Z�j�ҟz�0��@ 1,����O䱂�&	a�>���b�3��R��OF[��'��7B���?1P[?�#��D�v<��ĭĦQB��)Ţ#D����X�r-S���R�#VjT��HO�mZ۟��'X�9���٘"o57T�5�5�؂W�0�ʳ��OP�D�O���������O���g����qmޔ)�F���ѥ'��ʄjD�_��q���XN��s��3������	�X��p�͕X'��y�ˋ0j>�=�$��]����7�p�#�D�~�����4x�	�H>�Gmן���4Wp^9�"�*}<����% �M+�����O���'0Bx���4d@�q�G0! �!���]�'�����)@U:m�e�V�U�f�(�'!�7��Or�oJZD��T?��	a�Tl������M�EȐ��tJ	�2)xɳP�'^��'�4|� d'�T��#A$q�^�T>q1�S�%G��F��A@�.�,K�H����(���a8?FI����
q�E�gT���d��̌�i�漁Q/N9N��ܰ��O��d5�S>q TsbAY�}�Ĩ�ԩM�U���u����5�ꚱZQ��;��Mؕ�+�On!&�@�ń���,�FG�lA<%�C$i�<�L����O�ʧn�(��?!�x/�%g��:��@��v~��g�aƄ(RPU�T>��|�I2V�Xa��^�W͔�1t�Q:i�$��i��+�H� ��%}���'�����`�z��᪏�@�F(�7��LN"�'�R�'�?��V�_�����85�]�ŀ�X�D�O���䜭����I�:�f���딮Zs�`)����|� �D�L�ڔ��7��Q�+
��?��
��sOU�?����?�����.�O���X	M�����/M��m����6�^E��þWILYC��S?��h`ٟў8�0"�&1Z��2*�

���-�92Z�=�@;/�X���	�z���	e݈������	gV�Q �R�#/��ӲD�]�T�I�h�<�dLҦiJ���<9$�M�[���R��4q�<�g�f�<����[^�4!A�J8��RC�$D���'��+���o�SZlk� D'_�����A��w�	�X��������d���|*�F�~H�3'��[���f[�h��bԧ���,��(�$Ux��䛇'���iB�&E��ٲ��.��iX����*��bF��PK
Ǔy=T����H��k�S�:D"k�4]2�,J&����@�?!��9O�#v��&U��e����O_pT0��'�ў� T�â˞:*�@�pd��6J̼�#<OTlZȟ�'�.!����~
����	�|	0�iE�ک/
�5J�.��h�D��O����O����l�={$�}htn�1d�%�FL��D��;W�jQ��K6�`U�Үm���Fybn��`���)�Ώlt�a���Y�<$�����u���:50�����=�d���Ɏ;��d	��k��D-���BD��F� S,b�ն�y��'a�}R��+E���K�%\=\��T�G@�#�0>i�|�+V�&Y�Ĺ�%F�(�d�<�'��"~��'X"X>��0�˟����0�HW�2�D�Ab\#t��+7K73�=���@�&P�Cf���p�O���y���dN�i�I��X�gJ>x����f>@�h��N"�X��i�S��?��3b���vl��P	�����|
�8+��O��o��M#���ħ���Oz9�e�%|L\��t�i��,a�:O��d �O����\4G8<p��`�U�5�&9O���<�`�i��7�<�i_���T�(�����t4՚'[�B�b�'�,L�'@�5�2�'���'&ם�8�I(�$����	#H&��@�Zc��I:��+�ߝ���dȰi�4BP�!��jW�FU��C�+긁�-�/n��y��G���w�[4}��5 gmɕ�~r�=�?�Կi��O^�D�O�˓R���P��`)��`�N\�1��b#�T
T���ؑ���8�y���	e��U�܈u�4�M3���*��蘁&��l,�!ES��?����?��g������?I�O���)u��P�5A4��
Kn��	f�)n�L��fDR�	���THp81q A�'T�P����e>Z��#5+|@%���֐
��}k�A�� ���±�>H��SOw���q2g:��ޮo+"�'uD�zc�ïnM� �1i�l��-�A�'�T���	`�S�O:E�&A�!����OJ?�0<y�����i����i{�B�T*��(z��EǦ)��Iyb!@�#*8��?y*�J� 
�**�-	�왰>�e� '�� ���O^�d��<�"�O�O:�x�˙�ʧ"z)gHK�#9���WH�dEy��Ŏpz�6�9\d�
&���/چ.�M`Ǥ�%�Ȳ'ڌ�(O�ɘ��'b�'��W>x�l��`��acv�Y!Y.1J�ɛğ��?E��'Q�= G�etj�V�_DWt@!�e�'�\��ĥB(�P�b�I�M�� �'�V�� alӺ���Ol�'_l|����?�`�9R*�7��9���B"L�Ԁ���?y�y*��\DJ�@����5#0��Хb�x�	䫃o���槈��d�^�t�"�	�t����<x�q��'���O?���+�f=Ѱk�(F���#�Ύ�!�DO.0`A����v͛�/���(���?aa�d7O ��
�O�-w�M�o�Ɵ ��1LPU�[��T�	�X�I��uW��yw��m]��$dM="�2P '���~�A���>1eˬX���������:�Fk?q��Qvx�HӆIB�+9�Y�5��>β��5���Lف�On�d0���Ot���<Q�̜L�((EiA�9W�܂�jTc�<9���W2ؓ�� �"MR�b��lT����O��I=~h��Pݴb���eFP�2Z��4���0��ua��?����?�C�?�����T#�1~\��'���0�X�`��a��C��
�/�́Z�OX���4G)PmRF�T?ErR �S�'��Q�כV�5C��4�@�-_+�:�7��O�ʓ�?)�ʟ@��Gɖr��5Z�&_<QL�iЃ"O���Q�P0&� X
��Z�t�X��=O���'_�'x|"}*s(�KEd+��C�&I��@r�<Q�`�.�Xw 3O���JGo�<q��t��Y�G;s8a�O�A�<Y0�\<	� �@��qv�	�ю\t�<y���Z��]�3̓~�p<ZE�l�<Yq-@�$l���H��dU�h�bj�j�<��N�\�R�Jٷ	����A�<y1U�]Pa�]�?_r��"�}�<Y�@H�R��l���٬t���u�w�<�@M#zL�b��L�'DGx�<Y�K��Tl�E�A⃁	�����LK�<YAN(�\���ԼJ�^��F�<����2R����h��^J4L���@�<AE�0��Y �+G�z�"$2�-v�<���ʥ&�H���7�2g��l�<�D�L��
9CԠx���S!OS�<�g���|�d ���A�|+#�
R�<� PA3g�Ӿc6�h�Q�W���B"O<�e�4v�X���5�R)bV"O�	���M(PA�����0��ӡ"O��m�?"�]���+]�l$8�"O�]q�<p �YF�ջ"~���"OҩyE+E&{V��a�8@h�p�R"O�A���q� ���eL�{��jF"O�(�FL 30����#�O-fI��"O6$0��l!��\I"��z5"O���ǯ��T�`Yc��V�����"Oh�+�j�x! )�{�.�;�"Oi`uA��Ҍ0U�QS�\Ȱ "Ov�a�GV(F���T&LPҦmۀ"O��cY�yUj�Q'�˸d���Q�"O�9x`/L�h*8�3�מx��d{���Gv�7�Pe�'q��l�CY8-�������]v���Ɇ����<���,����;j?*�����<
b=i�j�I��ҩ8�8ɡ�(�s�)����6��m��Y��h�T'��5����i�,�i~��u�]�}�J��dI��B�hH�wش�C�T�D8(0I���y����ߙ
1�ȝ6�0��n��PҨ�2�1�O|���N�YL��s��H���f���
��N�mTl� ѵ�H�X�S`��j�p��^�M���I�<<���!T+W�%����nԸ>Z�a��|�fĘ~Z�`���95rX�A��y����	W�g�b����ԆL�aY�KL	�p�{�!ʦ��t�YlKr��$	&FxBM���<���_?���-yT4��C�8 ����ˠ<�}�Ł�|�#�_�dZR	��&�/�@��3e�{��J�-���p>��D��Lj� U�]���u�h�Č�E)�♩��6������6mT� �&��W�^	��t�e%�$�3B3LO:�ж�2H̒�����:w��� _�˷/;|kj��F�@�<�j�Γ1���ѝ<{r�ͧ.�n.n����ī?�
�)��@Zf�O
�+��P+?�f��r�[?pN��W���'����I��ڀ�3
�: �\��O(|2���)Ѐ��ڏ]� �I�U��I��-ʇ��[��)frZ�@��XZ�}*�I�����Ӧt�&������4���S�'�4lJ�a�H�yJ����f�(��3�*W�l�`%ؐ z?ы��O\�	̟�Bs��6 K!�ZT�4ț�!�@��(R˓N(h�3�S�[ V�S� #�&=��K�.I&�x�$ƻ8^Ll��$֛�M۲�iO��P�C�)u�<(��7�M7�'9��7�-t�ʘ�T��
e	�xRM<1s�Ǧ%��AE.n�rA���y�J�>��&ϴ)#DR�b�'_�R�ȱ��d��mٶjP!��|��'�\�az�A��u�����]�p/�"_<X���O�]� ��!�O�)���O*�*�hD%�p�'���BU�҇f�ά����j�h���"Oqb��3��8Ƣێ,�����Fj08�ŷi�HT���1��'΄��+z�p$̻G�L�;�f]�X�v�*�cܩ_�D����"N<pa
�,\M�FنAdt�&¦4�2@A�4�D�	��Dr���)�)�4*��S�'�r��E�wF>���&R�/�2Q���_�\:n�z捱Olb���䛙T"��;20��CH�8ڔeZD��on�@���i��%��EI�t������Q��k�.�;��q�1�E�", ݳ5Fb��qc��f�JV��{6�IZ�>O��� k�`�H!�'��<��G�]�h�PY��Qa���3��́ҫ�Nx��#eJ
E�ࣁEo@T���v�֐� ���A���	5��5����؈2T%#H���'����m�
Ɛy�EݐFu�|I�b�G��PP�c����Nؕ`&fO�9a˜�oI\����#>���v��P6�(͓,zb��E
G�Q��%z��
	6P69$��I���5R�mp�M_�{;H�
1�e�ֽ>���Еf1�)�Ơ`���)Z�h�})�c�0*�z`2�^�8��2���"�����6$�
U�r���giέq���c�Hҋe> #�ix,̻�'�4�H��06�
�'{���*�e[ M��N��\Ӵ�>-!�@�����WA��]��-q��.-���S��>0��'V�)��O���W���rUA
�ؼ�:~�`��'���{�7+�t�P�?.*����ێG����,��K��5�#i��< ���\�**����'$	�\Xa�A=	���,db��3�@�w���B�pm�'o�Y���C`�]���R�Q�&J����O���B*� �0�S����^���=OR	���5�8��1�<![���F�	�_��0��-���넷Ph��a��N� ��)J�^1�v�#<�O¦9S`�L*e�HW̔T7*t d�E̥��	5Z5^�tʎ	z`)3�$D�R>�䕰�(O1�B�*A��^�3�ћ�(I�#��}�F��-=LO��u՞=#�qӒ�)~phVf.~Ѣ!sdk�p�p�`�S�D���x�KK�r�p����ԁA�C�y"M�ȡ�b�C�'�y�%��ۘ'��x��497D�0��T�L|Jp�'��)� �p�U_(Gtrl��%� #����?O��p@/�&(ْ	�4�Z;j}�q�Q�I�uҤ"��@���q��
L� �$]
R<p}��?G�.��dQ��=���6��k��:_Z��)��T�`���ȣ����[���9Rm]4z9�}�dC�x!���F��~��[:��'U�D�����	Z��n�$p�=�p��TѾ���K�a~���Kl!�fF�q֠�+�C��`�Cb��&�~�N�X��� 
7�������?Y`��O$�I�nۛF4��� )I����&�>9�i$$���n�8	�����.�1�y�OS�扈x����T�G<$����_LVn6mĵWJ����T�#X��I���-Qq��(�����u��5	�B
!A��L�i��(*��Z�GL�P����޴\��=�)��[�Q��i8��G7�0#��<޺T	�ӼQ�6R�� S�
$�  ޵ep�h'���d�I�d�Ź�O��e#F�A35P�%A0pJ�)
�"���3��o�b��W�^1R��tL��`M+0)�$BR�`���Zq}cJ�	��ɕ"�(S���?I  ��	�Ƀ�X|k���z�<yF��i�.�u�z��^)R\zt��/ ���uߴ�y�� ���pgԴ4��"�iL��M ʆ�<���"$:��!b�'��]��-� _Bv)0F�D�<����ʵ}���!l�"��']�f��x��'���!$	��=��s�OB?T���ɱ�X:a}�;��	��W�2Zx�E�%B'F�`������O�A�.�J�j�4m�.85
��p1ѡ�v�.Xy4J���p�� �X��1r�ڃ�d�R0��Oę�T��a��AA�!v�� K��y�Ei�eY�Oo��Zdh�W}�(�0{rVm����+a@Q�x 8�+7��M1�)&�(?�Sf9b�;WD�1b�)hG��?!�o��$s��j6
����;�bb���I޴M���U{lN��X��O��{�A�!C|�Ě��Ǚu�x��J��t0��X�k�yb�K���E��!s���U"S�N�wu"��E���0>ͻc㤰#`�J�إ� �se�DB���.5�ər}#�͌a,�ɪ�)��h�01��.Y����DF���\2D˕�A�v���o�V@�� Z#g* � M�PY"	2�O���䓐M�4�u�J'�!�]�P�"2�7Ox=h��
k�zTa��J<U
C�����`۵|�<y���G�tCeI��=D���22��h��|�d%: ��At�V�Q�W�3�g����1s'�^��OX����
����X�i# ��冕Z y{���a|�L�DRx�X�#@o�A�Ѣ*>O�9B �Wk8��ݹ��xC��"B�qX4NT�x�*�lD�xA�Oƈ�GG�3�:��։��(�����)�V����"�`8�4�n�t�X|lZWAt��Dث��K��]|lQ�v ��:b�:t�O(��'���;%uE �4~6�P9hX}}��N��\)6$^����j�B��I� ��������!E���x׊��>)�8O�!Q	k4(�aN^�j���v�' ���N��Yf���"��,�#���ːz����'a�
]�㉂>S��� }�p��i�<�ɰ:����9O�!��\$���5oU�RQQB�
Q[�REƧyWA�h'r<j� 7#9�ئH���~���O8O��y�@��Er7@�0C-�[8b�ˁ��p<)w���n��G��gA���]nū"�
z DL���Лxx �a�1O��p' N����J�kH���r�r�I8 ly�CG�n�4̸��.�I�.t4ͻ��`%b�жG�t�ɬ{	�p�o���d!tN(�����!& �I+�V�E�:H�(f
/H�#>����A�`JE��?y�A�Vb�0\ZP�-�4D������*-�)������aH�"�����S�Ȗ�4�~����y�z8[d��Y���o�j��сX.
��|�fB2����TC=X 壊��܇q�&E"� �D�R�g�p���N¼U�X��	���p!mƚ,��"�G��z"h��v|��
�*63LN�z��Dě( �<��_~�tI�9f'�I7#X��N��c�l�� �~2�b���� ��Du0�-��jo�X:��^����#K\�M�b*ϝ\x�c��/Q���N�廷�~�p-��-V��k�$�F>��U�P �|�S�`�ݼP�f蛙:U4�Ǘ�p�T�
�N�>��Q�;	yP�����1�paY^#�f��FR>� %����Pu'��6c�����ƤAg>O�Yh1b+ړmo���`h�D#��^�M*
�@s%�x��P��ȟ,���D�k�����&G��b��U��X�);��YC��Ȇ���|��3�y��5`����7a��y�dH��~b�
���t�.H�]�L��������e�vF�p`Fi���=3�� Ǒ5�裌حB�J�1G� \�X�%�N���=!�b��l߮�Z� V3#6�yq�		B�6����Z��b4���ﮄ#E�ф�z�+1��M�]@CO��!AKh˸Jg��ʢ����T.1O�e)��?Hc��YJ�����Dq�`�;B�p��e`�T��V̣i̼��C;f,�b�Ma�e��@ Hd�	s�Ĩ�b�B�1� طHb�,6���M3Q��8%� �Y 	PK���IMu�S�D�R: qX�M oxR��'��1�� ^�7-�4~B Ы�����i)�扨*���Fc	6�b� �m�j_��h�J�.���c�"+��=� �yRg�a���A#�Oe�F�˃�ǟ ��<t��S�d��|x��.�|~J~Z��@�d��]y鰧o�nH<�J�
n>�IF޼��a�H�l4�r�i ��,O:d�L|���[9\&��'P�Hxc��W���Hkѫ3��a��	6=��J�'M��P@��DL�Ѥ��WFv�B⃦&��6��	4����؎=�H}����q��l��"�ֱ*�@X�6��0q��&���F~��E	GBR�k�O��s��Ħ�Pߘ~�^d��(�� �mA�@�]j���WY�)H��'�aA1�؇Y����"	�+3�XS�O>�F��V���l��'H��*g՟������4p�Jf�o�n��R"O�5����-�V�P��04!�U��Ҳ�t��'��
���4 �>����RF՘��Vn�0�P�}��ر�4D��q��-�Dyq�F�.dD�8�O�������H�@u�#��6e|	зJ������5G:m���K��+�CГD��Չ�H�*?�:p��Z4ӎ<Kd(�@	c��6D@N��S'Df�=��F$�p�(lA �i���>�`��R.=ֽt@�6J�z5 �J!D� �q�V�*��3�
M>��ef D�̂ ��.q����`ۇ��|(��1D�<�C��*g5���%����Z$c"D��A᧐#e� ˴͖[2fQ��<D���s��'f�9�6�5�Z���B5D����)]�Hh�� ���*AVg1D��ʴ�1�:9�%S�(��}8�I,D�D�a_�uf���`�)=�e1�)D�0ʖ�U�A���0���W���!D� ; A7� A;���4QaT�(� D��I�B�)�Fd!�@[�OT��%�0D�x�#�x�vx Y:x�T���.D�H d�Շ��0�	�l� Ku�-D�XN8x�處�V�&E�U���7D�0В��	���XE�S�%2���&)D����|�P
�P�p�=�q�(D�r���v@y�卮<�1��:D��@���D�YS�&�2(r8D�D��I(T2����j�.U��6D���m��mG����"�ch��64D��I�!��T��3,��xR2D��#3IC2e�����Z�b�	��l/D���`Js��܋��]!4j3��"D�8	a+������]!A8��$�#D���ӡD�ڭɷ(� ~�ؼ��,D�̢֪��\�p�bh�,v�� ��*D��97O�'i�Pq����h���Q!(D��`��[� � M��㞩z��r�!D��i�F�-U.K�� ��i��"D����
J�A3q�XJ�p�c�+>D��r���<Gl1�`��#�=��(D�tSP!�5���+�n�<D3U�&D��*3�D�j���h2�΄Ds��AF#D�4�en)sNf�p�i���i��?D��#��N?4|Z䂙�v��î;D��"�ƓB>��&�	c"=q7D;D�<n�llT��N�:9ZT�g�G�<Qb��0�"q����?���]F�<!�"�)$�d�g�ȯL�q��D�<��	[���y���Z�����a~�<1+�&L����U,�",�@f/�T�<A"��?m�(����S�p=(�Q',Gz�<�SFݯ_S��P�ǌ@�<4����m�<�qC Y[�o�z����`AS�<y��ْjR�����B!~�JH��M�<gX�1�M��#V6L�݂�ÈG�<�u�3m��y9�ΐ3q�p���FC�<iU��#�`x˕J([�8���AZ�<� 6�YSeC+]
𨩣e�:�.a�"OD3r�N�{�Fpʰ��a"O����G',8�	����(f����"O�m��		W��Q��GM�!�R�0t"O�L�w�_� �~!
��fs����"O�,��+�5�5(sf��x�"O�P��,Ê1��"ȅ0|�i�"O�%�w�H�IQ(�YF��.`|d�b�"O
���$�Q�x�f���@fF��"Or�ca�\:�����U2>1���#"O6��G��*z�d�5D�+h#Z@��"O<�R�*@�R"œ!c��D�b3"O�4rv�84Ռ�#��=��d"p"O�ː�Є<[09ځ��0�R�c"OR�{�D�Zc�1<&��% �"O��٥k��~v� �DW,TyC�"O�L��I&T�@Qk�_$�	+�"O�a��0E
MT���"OR��b�I�wgڬ9r�ǢaP�"O��B��L�=�6T(3��j,�M:�"Odh;Pϛ�Av�"!!��8��"Oz(rөܾ4c�Jsóm���	�"O�y�N%n�����/Z�j�H���g�O��H;4�՚UM�i!�TC1�x8�'�P!�$,Q�lJ�*��N^��'�� &��'�P�V���>�ґ��'�hC/��m���3�V09�X�����:<O����OL%R3 <�7,��VU�xk"OX}�waŧq &l��I1e܌�"O�9��,M8o����O�8#R�i�"O�rS��O�Ũ�,���d�"O���p �HM1�Ǆc}�i��"O��I0��	�*���j��JM�\;��	G�O�t���
<gBa0U�L-��)�'C���6�I�B�D	9%ە6�Ƙ*
�'5��S1ؚ��a�`a�&�`�
�'>���ꎹUkޤ��l�()�͘�'����s� � �`�.����'.�\������5�Wb���za�'Ɋ��pH�dN$Q��IB��B4��'�.�rG��$+2<D��ޫ{�ҡ�
�'�^�QSf�L��Xկ��u���Q�'G�������p��'h4���
�'2�Q�a/w��!B4N�J�t��'��	vmH�[S4"��?z�M��'j!���<3�U�$,מ �� c�'��`����0T��rK��b���'�d��׮�>�5kd��l���'mH���$y��8$�ďtf1��'d2�Ā֐sq~����	:�
���'��X������ڲ�ƍ�����d.�S�d$޿3洌AV5�����A˅�y�j����p�&.|J���̟��M���s�S��I%���s �Y�"O�1d�͐a#��H��W���2"O��5�UH.h��$0�^��P�'[�i�[�.V���V(ܪS�ꘄ�]���k��^�u��HP%'�j��<����#��B�cQZ�4*Z4�!�>}T��Y��%,�P
0f�!��1�z����T3*�K��ݠI�!�>��d`��A�Q�p#�&	�!���8h�F�cO�/d!����Car�O���R/#xjF�)P�1mk��#"O� ,�6��/�X�3��ϾR�`�e"O$!`D�"R�M��Ǘ_���)t*O�`���1 MQ���P�,�z	�'���2�V/%p ��r�ٗN�� ҈�9�'R��I�Hաy�zဪ?dw�I��0	s���a��X9!1O�0��sz��k��i�V��嫕�wdd ���0���a�� ���/0~F~���&!�a	A"�5<��jd���-�ԝ��a���e�4@\��g�Q�Di��/@ب�F�de杰��ǳ&����/�)`.�1+H��Ao.3笱��(*<�(^" ǜL�j$rЉ��~2���^�U��D�&�0�t|�ȓZ�{���?6����?Q���9�VI����x�E' 	�.������'��=-95E� �i����o<��ˤ�;j-�E�k�&@X��ּ��+y�Ѩ�"M9�V�ȓqޜR����'��`�l�k�r	��W�z�²�.3x�$C��x �ȓLf�I��o�u�4��m� O�P5���
A3��vz$9Z��  <����2)��6� &>����#�5f���u�D�s�f�8�2)"@�8+�}��4�n����C�6*�pHE���oI�	��K~����R4"Y��+X� ED�ȓ3�dp@B#�$g���Uf�9��a�ȓdvT|�C@ã]7�S����;N<�ȓg*�a���7F?�����)��ȓ.�˗/��,Ⱦ�cb��=�XH��7�� aE�6vִ��c�ÚN)����#�8��ܡ]�l�E��R.���UR�	��6�=���
�>"�U�ȓa�d��u�ɳ17�A%L� +�5�O��!�I�:N����W�-G�8�	��^����"T��p�в^* 8t핪	!�Q�~_	��f߻fJ�4j��P�9�!��߀"�����3;n ��A�;'b!���n��p�N4ٌ�����},Q�@��I���]���-t]�ɑu�=7&B�ɰa�<I@'+�Dw:�A��9#�dB��$X����wb���Uꎧ4(B�	�D����M�S�T�yvE��H�B�
D�0��O�IV.� O��uZC�	�"���+V4<��8#��b��Ĵ<���M&� ¦�P�-���9s�Tm�<��Č��N��"���jΡYQ(�g�<	UF�M��f���_�F��|��U�xh�q��$v0"� ଒8�`�ȓ��i��J�J�B5Ӑ���X/���ȓ��� i��>b�A6�V�-r�y�ȓl� u�q�F-R%�^5u�9�ȓl�ZT�`�Sw&��i��OG@؆�z?4�1'h�"^�"A8�-��k��h�ȓ5p�9&f@�fC�Z��y��	��, �-���qn�
R�8	�ȓ f	Y�������c"�0 ��=���h��C��� '� �f-�"'�8�ȓ���D�.]@Xؓ�E�}��|�ȓ`c\%����D�=`�� �$T�؄����WCY�\r4��˜inh��x���a��2	N�sw�]#�B ��A[2L%�N�,�Kl�7<��S�? Z0)f��R�:�B���x�52�"ODԙ'FY�����M���4�"Ov���@�%Lb��U�ُbc�Ac"O�
��L��F	��D�YJ0#"O�|�`�Q:"�x�� ^ |Ux)�U"O�x��HѼE�(����0n��{#"O>u�	A�vi��O#~ ����"O@���I�F(� 9�E%PHf�X"Ol1'��'<o�0��"e���q0"O�6Ɇ {J�@��A�VҙJ "O�%�d�Tm���q"aT� 񰌘e�������=�*���v�� ;d�Υ �`B�ɵd�T�%&THD�t����]��C�	�*���kS�����S���r@B�I�xx�����U)_K�آ���"eB�	�-�B���9 B�j�M]?QB�	;Op�C��<�zl�s�٬N�C�ɵK�n�Ქ	Qtx\{��(;�B�	�Z�n������fD����/YOBB�?1S�D �Ō1_J�"@�t�$B�I	*�!Po��)$�,�����1�*B�4�^��%4��詴 A�X/2C���xR�ެgC�P3fTw̺C�I�i��	�Ђ
,@�Q���̇`k�C�����/C�!��#�
�_�nC�,,�|�bQ#
?$H��#�C
�yCzB�I�^�츀���3����-K��RB�I��dՈw��y��8���/�bC�ɿZl�U�7"�.���߬4m@C�	�b�,hG�\�Q���jR%�0C�	�nV��JR� ��́7A��(W�B�=>��T�Q��rX��:��׃��B䉩(��pc�e@V��*�S�/��B䉠�����Κ#*��X����L:C�	>h�X�`���@�p��Q86t�B�IL���������PC��B�I�w�@��eC����F�5vm�B�I�2|&H��O/:}���c�#vO�B�	#g�\�4�71������c��C�I"Q#�и0�Ѱ6��͈q�A�U�C�	,:�(�j��	�<�^9F�I�\C�	�U^�I�DU�A�@5�b�M�=VC䉞�����M}���b�힅W�NC�	:���CԅZ�liy��cC�I9_�j�*vK�"Dj�1]�l~�C�2���谡��
�d��ƈB,|C�I	�vH��+�y*�!�fX$f�B�	�(���胆|��Yz�c׌F^B�	LN=��+��Kw�>��ȓ=S��c�7[��U�̨��ńȓ4�a���q�j��wK[�nv�ȓ)}:]��K���*�.)	
����f�`lɤD�(�v��Ɖ�`�Hņ�0!�9@$nG-^��DXǄ1=X�ȓ�<��˝;����c��
J���3]4�z�đ�Pq.Ų  ��V�,5��/���"gj͋U�bш�-VPl��@�P�+��2���!�*#�Մȓ`��<sǋ$	�5nڤ����X�Œ�aڈE��s����[u����s�Ze��M([�!Z$#"��ȓv����1
\��-c&��
`�,�ȓhi��)�*���Fl��uz��������90Ծ�xB"Ԃho���S�? ���9J�XC����V�#�"OD9!2�BwV�h16�B6X <ՠ7"O�1qV�Ɲo42A�@�J�e�tѸ"O�U���V*@D�QI�}��	�R"O���̅!D7>��s�ȫ:_����yr�ƕy
0L��!�C{�%���/�y�DЇn8`�04�P�4�M(� R�yB�L],F����0+@��K�9�y�Cޯx�8+��ײ$/��{6�֟�yRG���ހS)��F��y����y� D*%;|/d��ǌ^�n���'��Pq�AB�#�Ł��*����'��U	�"�
}���k����'��I��+��7?f�H�����DE��'y��D�۝`$�qe�0N:�
�'�6ѱ7��j�T����֥v�t��	�'���C%j�=t�<���ޒj_8��	�'JV�C#mΔN�V`�I�V$z�	�'���QT&���6N�K4���'�1��R�9�uˏ�Fr���'u���N4|�mR�O��r��H�'ʚ�KRO$l ��hޣ>�,�
�'F��L]-3,R�s�F�7�0�	�'^��	���.Y��;rC&Cxdt��'����`V-B��=��Iĸ�`p��'�4�Ï��0���tA�R�:��'z�0ʠ)�xc\�
e���[Z�B�'�N츀�2���a��
]����'�v	Yt"�$[7�}+�K2��R�'��$�5ɐ&�eR��MT9
�'���C7n�2B�݂G,SC�L�	�'�*Z�̶Q�Z�5)�f>̭J
�'�T�M�J�(li)N3pu�A
�'j� f��C���*2a�.qJ	�'���Â�H�����,9
�td��'�&Dx���;K�������%1�'Ӏ��W䓄x���*[�L�~�	�'6򰨧�U��� ���CFU���'x u�e���\bN(�fg�@�F�'��Q��A_pqi�B�1�,���'�$
�l��N�ب��Ɨ*��R�'��̉B��!�t��a\�5��ȓd��r�`�<huR 3&�@5J.���'Q��)5�؊ ���
I��)@ܑ��v�p��B�X��P��3id�ȓh��\���?��A�� ����I���
�j5`?c������^l�t�ȓh9a��R|H(�k�lN>H\R�ȓ"C�D���(P��1�m�2T�b��C�2��!O�6S�t[�.�++^؆ȓY���sW&��6�� R�凰M�}�ȓ#���s�/�J��c��V��@��`iJL�1�Rb�ʰ[��G(/ZF�ȓ%J���'��[ivDs�@$6@����xK���~j�̢`�؊1sz���'j��⁃�5h.�j`ǋ�3[���ȓ'{�p)��9'9f�{��P�(͆ȓ5�ll�S�&@E��ya�y�ȓ	��8"���jF�9�e��RF�T��<E�{gAU�.b���D8_,p����8i#@����Ia.U�q3��ȓv��8�4j�1�^]��� �M�Ё��XX�#�=J>���Oc\�a��"�L�N�J%Zp���g��݅�S�? �٢��BYz40������"O��q��r}���E�N�@QsW"O��P�I#_X�9�ȗ�U�"���"O����A׈�xz�����QH�"OdA)��r���Z�gË��*�"O�L���@7gBuig�9s��=�"O�T�-?ň��U�Fݺ8*�"O�}#�LG6ɪ0F�X�%���8@"O�5p�g�"4���Z�AƇ5����"O XXӆ͟^�B�P��K�tP6"O��+[�"��&�M�6�tQ�"O�Pj��b�T1 g��:���"O�
�FS�J�4�8��xCa"O�a���Z!A�9�&G��*�^�cS"O�p!�O�o5](�ȵ w}!򤊜d*9	��7X�,�K��EBW!�Ä+d��@�?��㣣\��!򄕁{�Qk���XT�1�	
 t�!��25�|a!�ӭn���5I�$�!�$�9l�D�"�� |�z��?�!򄜩2�����]8=H ��^3G�!��O-M��z'ܞN�PbaeؐNz!�K�Pr�����>j�53D�T�!��ωe�PxY�CP56X|��6�B
)!��ݿm�TI#��J疵�%.�PG!�� � �!]�Oɰ�1f��zE!�Ge��z���,&���wJ�X�!���`3&�8��B,m H���7c!�$�.1���f��)e����"gf!�$X�=��9(�	?(�٢C�T;�!���y2��d_<#!"���SrJ!�dI�
H��`E !��i���V7!��&;�Z���MV�u�FтCK�%�!򤔹xH��2�2&�E�F#=<�!�C�I�Ap�H�8)wźѯP? !�5�PT���XUs��Rm\+`�!�̋��Ē���;n�	*"N�a�!�$�i����蔛x��R��|!���SK�yq�
*\8��C�Z!��ω}!�sCX���y@u�,�!���/InA���۞�Va�+A�!�8�d�� '[�pB�@љ^�!�$R�@�)E���e���]�!�$�-iD��q#��@���+ՇK�h�!�D�7.mj���/��`�V	9�!��ޘA����'�]����1�s�!򤂶}X�U��-Ol�h?�!�W�H���y:�� ef��&�!�Dƒ�x� &�C�48�e�R&��\V!�$�'N��A�ݰW�LS�ė>:!�2j����!���-S@�U�!��_t�B:�n-%�� #J0�!�$���,��0l} ��:HG!��9D� ��?.���E�,4!���i*T��+�>v)>����ţg�!�D���H��I�1�8!�G�1��<�f.X5u�R	��!��2K��ǣ�<�`|�Hg�!�$/��x[���k�pp���,a!�Ά$�fec&�̄`����	�Y!�$ޙy6�'���������\!�$��~��RA��BH��R�Q��������8*�K�.�
�����	�Z�`�$�'Y��:�$v蜄�S�? �t1��%5�-*��B�G NQR"O����ꜥZ֊���'�"��̡�"O�E�����Rs�W2p�S�"O섈'F��E�c�8'a"O� ��+��+����O(V૥"O\eI�ي9(1$MW<eQ*)S"O(�A�'�T)��댫*�T|��"O�s��'���&-�������"O^��f&��2�JG�_=d"Oѧ�ɻ�0�����K=0U�"O"�v��b�ࡸ��B�R��5��"O�a+F���n���;������"O�YR�ޝ��=Z2�����/!�$�&5D.m���Ǒim������!�$��f�dڑO�4Hq��3S>�!��߻xcD��2-� [��!F�E!�$�#@�p�5g�Ka"QU��(Z!�^e���QB-��RJ"}c�C��T!�
�*�"ɀ�#�.{n�C� �D�!�d֦��}: C��cX�He�9 �!�
�
ʋ �V�	p�µzu!��Y�c�4��X"VD�p�͘�+`!�ď�o�慫�KۙS�(є!D
}S!���/"%PL�e]�s�t��"�0q�!��Y�I ��M)�j!ɲ"ͻ�!�p���K9@�Fe��a%�Љa"O� s��t
a	�,XvT�"OH%��.�#�H�����*��՚�"O���A�3`�lq�f��g� ��E"O����)AI�&��B��I#�"Or̪�@�$�������F�Ό�"Old�Z0'؞qBѤ�~�RE"OL1b�Ƀ%K���@f̏&uF�[�"O.��bN)2K��QGK̀�uu"O����K�"��|CDK�����u"O�� !-ߪ�^eR�	Z�@�� ��"O�V�����Y���+�0�p�"O~U[���v�0lb�öh�� t"OJ��d�r���C\�.�"T��"O�$	������d�� ���"O*������Gg�(Qsb�=��	
G"O�\h���f����@(X�썚r"O�Mx$�F�x�!o�8�\�4"OrTҰ�y�ļ���02��� p"OH��6�|���?Q�b�s�"O$��У�����"
H����"O�L:��9\p��d�P��"O=�"M� o��z�C��N�zg"O�i���:n�B������S%"OJ�b��	��
��N�����"O.ѻ� ϋRP�P�S	�v���Y�"O��p6+�'f0�L3��7Sr�4J"O�M����<DL}�aj��%_���w"O�@�L��6�ʐ�*L�\P^��"Ohm��ʏ�0,xa���4W5V	�C"OF��ԡʌc��cǻ9�����"O����@ƪ�B��l�S"O8ʣ��.K����P�i��p�s"Oؙ��nF�"��Qk4��4��"O�Y���	�L@R�ߡH��<aQ"O ܛgIO��\DPGY�W��%k�"O��x�OS�)��la � %�}2r"O"�e*Aqi@���mL�j�"O��Kgς�$�zDACΌ�*9 	�`"O� l,�&��"�5(��Lܵ�e"Ob%�D�	>j���&�5��zC"Oh�Nq^,H����j4n��"O�P�QҦ+|�T�`D�	I8���"O����I�te<�%E�;-��A"O��U�H�&T��v�����"O�@�K� � ��%��t�x�Q�"O,�)��GR�����]����"O�4*�5x�XK��-��a��"O��Y�����!0��O��8"O�3�d���,e�s	V3bt�ݙs"O���G�H���ס���p"Ol�zr�� gz�r �6Yx[A"O�ū�HN1w�<�B�K�+X�PP"O�JD�3Xꘁj"kǠd�E�3"Oh���LuPy�q�A6t��B7*Opu��F0#�0���
�H
�q
�'����u��V-��[AE�+>Z.�1
�'�搋a�_\T"m�+����	�'��R�a8_Zp��Q�%�U�	�'�	:�J�~�H\JqK_�3F�E��'�0aa���+jyTTH�e>$SN��'c���Ü���<�0hI��D=��'��򰅚���ij޻!J���'�D���$]R�%j�
�B�9��'q�p���_�a}��
�%X2���'<J%2׫�*��[���z���'�PC2+\�@A)ȍr~�qh�'|��&��1@֌��␈cŞd��'8�"�>�6Th�@��a-�-(�'���ہ�̹JT���V	E�9�'��} ���6X���Q��(Ӱģ
�'RD ��ݝa����� �=�&��	�' E��̕�HyqҡX"����	�'}�i;�b�	P�܅��M��~�⬪�'<^]ztC��%�ę7�۾Ls*)��'|�סR`���)�f�Jtt�
�'4!s���:Zˎ|k���	>��� �'��"K�>L��!@��80�:QR�'�d�4�=z�(ER���RHrq�'�Ƞ���]�,�&M*r'�P��A
�'��|�t�S���1���B�Y��'K�q��ϊu(b1[�
��@
�'��ZQẸb�t�' �1���S�'s��#�2��$��A������'��|���2=�0�V͜�b�x���'�\K!��;k��'bL'�:��
�'�L$���Z�7�2���/F�0	�'N���ύa�p���V>nŴX!�'Ą�i�ƴP*�c�[�g�h��'���@sL|Ţ�Q� b�N	��'��:��Ԩ$��1��V("(j�'
�D��[4}TX���G?*�;�'�D�8�#%<[��sΜ�Fg�5��'0��*E�����t���k�<�惇�*X&q�O���M"��a�<��_�1%l�`����\�ar�/D�T�6*�0�l�$ɵ��ԩM-D���J nr�����g"���,D���aA' 8��?!-]�Rn8D���Rz��A��)x�HI�4D��cq�ͨnN:m��R�e9l�`��$D�T��g�5<�}�4�J�4�1��"D��A%L�x(�	��>2�M��>D�� ���	�`��� viS����0"O�`4&��I�P	&���n�"O��J�O×~�����ә4�$�@�"OV�hWi��1��&0	��)3e"OT�b� 7֔��OO�=Ϭ�S"O&P@�b������A�n��%"O~�`猻V��BS�À;�Ȑ�"O��k��V
�|��G
1��C�"O
eh5��e5��S�ЏK���H�"O�@�
&�`\Ѧc�Gk>�{�"O��T/���4�1WB��>���xr"OX}�F!�o�L�ӎI*�8�)&*OD���	C�7$iZ�' �Yǜ�a
�'b�Ps��� X�w�4;����	�'�. �&k�[�&!��Ő8� A	�'
U�ڸ~��A�� �7�m!�'�x�2���-��=�%�GYLY8�'v��
�A" n��ܰQ�T�ʓ&�
�(�(��Ggj%۠�:1�h��ȓjn��I3
�-%��
7�R �y��c&P��J���ht�ƱE)�5��"�И�CL�;y4�a��.M.1�t�ȓ&�\X��Q-.�9�T��&+#��ȓ7�8����!���2H��uh�ȓj�@�7�FA��� �瀏6�<ȅȓ$��B�E�L��dp�B��x��*�
,�&̗9;�8���
�`���}��HyG��$1�Q��>/f<U��y.�,ӕ�:�32&��](�ȓ� S�j��Uҹ3T�K�G�$�ȓ
�*���@�E�����J �u��܇ȓb��l�ӯ�*�n���o��}f��)r��ҨC�͒d���I�Ț0��Qw6puF�*C�$�Ѧ�	;�,��#<���	�d�p�GB�vz΁��5䮨��mW�O��)2!�.���W��}��'I�!�����_�.n\��4t��Ђ��=Ǧ4�/-=2�M��RKnq�*S3"  4cʬ	7ք'����]�������3����.w�DC�ɌJ��r��n���be�%-tB�I'�X�x%��2��f6HVHB�Is8��l��z�Z�"�D�:S��B�ɑJBt�ED-�n��ͅ�"C�	�e\�թa-?|����@B'XP6B䉘@��u���ė5c�ષ/E&j X�O��� LO��D�>x�|[�����l"O��ׄQ�%��3a���P��"O��a�k��b1Y��/�(�W"O��w"�^�r1� ����i�"O��1C��0Ҡж�1<��$"O*�R�a�?^(�u$0e��H�"O$�锨�4&��J�c�gTr=���I|�Lɡ O{�mZ�h�%���q�=D�H!�,O	|�~��v�1�P��/=D�t*���Gs�u��E�/
#���w� D�����bf�ȳ̈.ua D�� QH�D�!���F�F�[b
?D�$�NG
ւ
�c +�p�HcD=D�8����NWP�`ς�x>@ʵ�<D�c��s�DEX%_�k�Lbb�=D��y�n޵{Y� 4e��E��*:D�\���Oa_H��fX�E$|0I!�7D����nՍp$H�+#
�S�&=�%5D�� �\pF@��2�B0;���k!"O��ҡ�Z�
I��A��13�"OB�Ȁ�7o=��C	K�j����`>��G�ƾD�Q�D���n%X�i"D��,ڸi�#��pQ6Ū�#D����bS�8������*q�."D���!8Pa�K]1F&��$K+D��sU�&eHڈ�����'Z�8�)D�`PPm~P��y#��7}�*�i�E(D���'Ɗ�e�,1)�ILI�c��&D�;�K	(o�V`8�J�L�,���%D��{UP��h�(ʝX���ks�#D���Fh�&]< ��.I1J�xA�o D��x0'�<{��e�EH�x��-?D�<��'�+�Q�$��J9�`�=D���� F^�&1s�/ߨ9�|yaT<D�����"2D4�f��GϠ=��$D���s��-b�Q��93~��h D�d�7�^�D��! 'M�=�Fђ*O�CR��h˪���n �Z�-��"O5���É^��+�L��t����"O�HA3���2�4��W�A�}�DAy�"O���/֤pE�A@�KQ�Xh��"O�Mr�i�YD�H�E���~p�iڣ"O��������|{'��hV�uRu"OĳcB]�-vT0ѡ�%9��Ԙv"O@�Zr�F%��` E��&�Y�"O �:�B>y`�q�D^�aX�"O���hV��S��#/���"ON�W�1*X$�@�AҚ')���c"O�2�+��v��`#qa�i\�f"O����̽1nb=�Յ�!�+\3�y2Ǌ�j�@�Q� ��%�>�����y��Gx��e�!��m Ǥ�
�y��ے8G���0e�!M�1š��y��+
��%+'d�H(�Ԉ���y-].BF��GIY�[�mJ�j��yr��_��A�/�E�b��CeL��y�M�#MGy�r#\�
"D���V��y��\;�p!S��Ѵ.RdC�*���yr
U���+3�t�g�Т�y2�^�.w��V%3A@0�Q�0�y"A�"ΉqFG�3xI8�c
;�y��'r�����Ґ��	��B.�y��̕Q���
y�H����yb5zӞ����Ϸ�zd��h�	�y"
\ �e �mO.R#��D��6�y"��9���`Ň
8INd[f�y� � �PX�`��0
����Ƃ�y�o��p���;^	���yB��	)v��B4��3a̤r��X��y��R�6��HK�ㅤ	fi�aȉ�y2a�
*
�de넑����-��y"h��SPp�F#��	� 8Sea��y�!�'B�̥�WM�41ba���Z��y"	HB�:���+�C6�=A@� �y��w��)qG�<��:�i���y2�P�B��\C����J��eX���y��Ȫg=�l��`��`+"
��yn<P��z%-ޕ;�\6c��y"��b�%`A*K.
"���e��-�y�-@���u�4Oʜ��DN��yr�T�3�:�yt��H�bMR4`\��y"�9,�ŪT�޻Fb%#!+ �y
� ��X��)=픉ӇՎm8吤"O��DB��\=B���jh�Ȃ"O����A��M�!"f$S	�(z�"O,=�g��+67��`�����R�p�"OD5���*��X�ǣ��)�PaS�"Ov��3ޔ��J.k&8���"Ordpӊʲu�f��s
��K~d�Cv"Ob��s �I4��A��؈G��+�"O�\bA �$~��C�׹V
��9�"O��@��h��1ysLW>}�Xr"O���&�V�GV>���jA�Tu�B"O� K��/Ax"%k�cE�A�҂"O\<{ЂauL�!��؊^�b�*"O*���ޭn�P�kB��&%�4(i�"O,�(�I�F�� Å�M%D�����"Oj�K�-Ъ:?4�:�N�)c"�٢"O��j���M�����Alur�"O���C�vv�D𱠊(VgX�H�"O��c"�M1(#�����I5�M��"Od�jC#
�`�G�W�f����"O<���J�iά�d��>,��"O�Uȃ�̦A��I�4�������"O��q�۠Yv�aQեg=�Igo�n�<���F67����Kd"�෮�k�<y!��ޕ�����]آ�	i�<!6�Y-O�Ft�5��E����@�<��+S?K���(�>Bb������d�<��ψg���ۡ�P=QD�;��w�<@�� #�\B��606J�{�g�Z�<�E�6#v­@D�5H�^���k�<�6Iʘ>�8�� �r0]ꇅf�<Y@�%aY��<OJ�t�j�<yg� �hz��VC��"�A���i�<Q�L2!(���V'ț -*���b�M�<a�C�}�ȱ@�G�F���*�d�G�<�Ђ+HV���營�a�l�A��N�<QڮM�`�Vc�!d��Y:p`�I�<����5X���Xad�!���i�DP�<�c";+:l��A�M%h��D&RJ�<I�aP)rh-����H� �J�<�!؇t~:��,�7|Z�x`���E�<	�E�j�t�4�(q`�cR/ZC�<��#�=��X���&{�Bu;G
D�<�������!6&@&Q�d�@0��~�<!�,B�t��)тMF
#(P��F�O�<1`�P$O��(7L� h������P�<!�,��9��0a�L�b�LQ�_L�<A�f\�aP�L:A��VQ$ �ğF�<��B\�p.Z�"�� �I�<)F/ٌ�(ɲv��bp��Q SH�<�W��1�r5�e�%����Dc�[�<�pO7%q��a�)�_L\��Y�<���<
��q��F>(FN9ó��S�<��G��i��>1?�`H�O�z�<9�+[5Oȼ��� ׅ,y���V�o�<a1�	-�> ��;��"��t�<��˖w͐��V*S�,��+�g�<�d�25�����ą�s��ʲ&d�<A��63xn�QSAW�M^��Xb�<ѣ�K'��H]6�@�F�\�<a+�~4N)bcŶb��H�(ZV�<���.�����g�2L�@��
�R�<� �!B�4��Ԥ��p�p�X�<�c	�r�0�����Q,�4(�F�W�<� �	�& W>=r��ab�,7hXz�"OP�@!۟[Xy�ԏ\*cM�-�S"O�T��C�#�`�a��`����"Oh��b�^O�@�u$?�� �s"O����ڨ904��	˃Ph�L�@"OP�{�&@.Dx���GH'}Dt�+�"O�-I��S#�f��5r7ҥ��"O����M��i(8�S�&T�"��&"O�X3��6$8}3f̍/(r�"OnTK���4XNp��S�F=��A�"O��	T.߃J]�`�ϐ	"���R�"O�h*�E<z�HR.���f��3"O�T�o�&e�6=�֮D!�����"Ot�9b��>�0�t,�7jۃ"O�HH���*�Q�W�ӽ�0]!4*O�q[�@
/@���a�4Sy�'���B- qbxa�n�&+����'ͨ%a��\AG��0�Th�2�'adL��@u�p�Dć	��0 �' �̓�Ǔ�v��<ӂg��$}��'���:��<=[��aH	�-ӮY�
�'w���Q� 8R��Հa,�7��i	�'3�%+e�۵G$	��X<Vq�'��ԋAgƨ:OFH�P�^2�����'a�	"Q�'w��@Ɓ�3d=��'�"�Ae�$W�.�i���y�@� �'�*���M$��;'�
n�`8x�'�tQ[2
��w�����
�n�jX��'{V�j�f��w��pX�s0lD��'�Z���Y�#Ӱl�p�ЬU\H1��'| �b7hF�4sA٦��V�P(�'P@��͟O��,H�jL
 G`1�'�9�c���:���A1�ZNE��'~�HH�ȢA$Dh��_CR��
�'��!.ޚw��i�/U�
�m�	�'0�<��&֪a)�S
�h�#
�'�r$8dI.)�t�s	$pX	�'�XLA���� U��Ї�A��y��' ��� �N4k�&�cJ٤C^�2�'��Lc&+܏""���N�qH��q�'��,�7�	V��Z�@�Z��Y�'ĠI �H��p��L�
 X(H��'��%�˛o�2t����yl"���'LD����R>J�\�����	��'�X��s�(a'����c��W����'ErY�Ҭn��t���N���K$��Q�<�fC\�}��#�X�
�<�1�x�<����,tΌ����ۡ>]��EƓI�<��d�
:����'i�>j܌�3�]�<���D�xC�PQ ���\P�^a�<�b_妝;"�
4�@���\�<�@oV�j��a�ńW����&�UR�<Aa�0b�v`h�j�5C>@���b�<y�GaK�U�o\/)��5{fj�s�<U�FHX`Ce	MA6\U�<	�"��wzz�bD��8JDr%��[z�<� 㗠s�v9y
�	8�V� 3�s�<�T%~�2L���U�}ȅ��r�<#�1z��9*A��:l��A�dEo�<i�,�	�fi2�C�*x��cA�<p�����
�D��|N،�U��r�<�B��].�����l���R �yh��COx᠗����*z�/�.�yb�W0Z�5�"�W�q�lڂ�
9�y
� ��S�	��H�24��
O��"O*��Dź������d����"O,��G=H�����3����7"O��3g��"O�q�C03m�0�"Or �a�
|ܰ���й{g`�`�"O����؏y���g▙HIp���"O|�Ǖ�DkzD#�a�*@H�	�"O
���ۧVU8��v �I'(E3q"O��%�2
}�G醔h��mp�"O@ ��Lv�k�h��mG���"OTL�ቇ�t�� @���.9��J"Or�JS+ә1pM��E�-X���V"O �"Ï�.�r��v@�;;3�pcG"O�`G��_���{�n�\�R���'�:D+T�-xI!G�Ύ6�6�0�' ��1��K���6-/1�pd��'��A��ndH�ő� R�M��'��a�gE��5̂��qL��vK�@a�'��!e�
p�l���.�<�x���'�� j5�Ԭdp�ɺ��]�4���'{���="6���X1z���	�'��D�'���2Uˍ!u���'`����;�Ҵc ���"�'�$hk���zU30/�i8q��'��!�b�9I��iAg�Ԇq���'�z���AF~(����D�2�X��'�ҽ���Ӛ�i�3@�z����'Mv�!��;.�HL	�g�?m�H�	�'VLP��&-etHH���^z��'u�u���� s�8W�G-���	�'j�a��ܬ��t�s���O�DDy	�'9D�#s"O�֞��ÅًE�T�y�'Tx�Ct�X*�:0���7x���'c�L�¡p�&�pk��)�n��
�'����4n� l��(K��25y  `
�'��EzEi���)���v�h�k	�'3����4xt8i�h@&m ��)�'��@vb��I�V��`���`IN���'���5dD���-3�h�3��[�'}��#�,)f�����y��1��'&�q�7��=k�ѣ(ArC���'V0�I��#z��T:p@
	q����'@6*�MN	TX���/_�n7r4c	�'Z�=k�.:����ADJ�m*�$`�'E�)3%!�'�~�Jr��zC����'vx���Ȕ�J$��`A�
H�q��'.dx�a�d��5ZԊ�6?�'��Q�$��)8L����'��-��'I~h�!�@�d���
��`��'
����L��e��a)9c`��R�'EYe��0��pPa[.-]��'�@���%��gz�Se%U(0�S�'��zV+Z[��Eň6$���'�L�c�	�[�p�Dۆ�Vx��'�PX���]�F��a	W��q�'E��+�eG5/�t�bQ��1p͈
�'�Ҹ�`��s�@�0͇�f�T�{
�'�$��'O�I�t 0dʟ1���a�'KDؠ��[2�7χ�/8,pX�'u(�k&��>vL|IR�! ;#�� �'��H����%�2�j�h�4,,21B�'�����O�ԉ!�� ���H�'[(h�bX�R�Q�A
�9G��pR�'�� �!­2���Z���7�T�3	��� ~����4 ��#��זf5�аT"O��;��֘�2Y��R� �T"O~q:��8Jے���`��y�"O �[ ,��zR�@�� ��@Ik�"OV̈&'��$����]@�Zh	'"O6�!Gjr���`֡������w"O�P���8b<X��S���X84��"O�bRݦ!6�ڧG@�c�hT �"O��Y�I�2K�(��$���F=(#"O�=9�o�g/�|���ՠ+t�x�"Oh�)Q�}׺(k@��#w�}p�"O��s���	!�.U���-Oh�E�"O� H�H�!�m���d��ڠ"O�][І� :����@&^B�"O�I��V�I[R�@�OS�,Mj`��"O��c�de*�C�)߿>+\��P"O�m#��וy1���"��&q? �q�"OdrcM�nO$�����95
���"O�ik��:J����`��XzD�"O�h�7�w���3gӍE�\���"O��M�rC�AbG	�a�Rq�"O�x@ B�:(�V�*7�A-\	`�"O4T��膺b+����	C#�6�pF"O~t���W�k��@&�A�V6���"O��4��0�l���U�D"O��4LK7n����7vӸ�"O�M���:#llP����Y�t�a�"O�=�1�߇|�F�1����"Ohp*b�4��%����k��Aȥ"O�|A'iҋ;��@+��0 eg��*&!��i���e,�L�h�a C�i�!���^0H@�V%�"��2���!�м*��
'��7$�kRNɫ{�!��Sy
]@�# J��C�A
!�˳8�^�����<	�p�Rɕ�s�!�dd�2Ya\ ^�Ҵ;0+�3v�!�@:�<�喺z������)�!�$E84`�3�[�3�= ��Ɋh�!�dL�܄(q�E<.����O�$�!��̇!�0�@16��%aƀ�*>�!�Ď���-P"/
�f�@sB@K�
�!�D�@�(lX�$^�?��-�b�ʎ<�!��
h�`Sœ�z��}br�]�`�!򄃅Y~h���R-K��]����/!�-{��,Caʖ��)R W�!�EE��h%(	>��h�n�2r!�D����JE���,�*� c�¡[w!�s�JmR�`�Y�r�0��L �!��,49j�c��1�B�Bv��-_�!�\e�
d�h���Aj�!�C���!̚*01#�㛳+�!�$:#z10�Ǖ�d��QL"�!�	8��0��!"5(�MM96!��ѰKlM"��W?^�FLCW�Ӡ�!�!aX��q��3q�<}�s#ݓ(�!�$	�t�����G���TIYF!��;GB��ӅWnP���
<64!�DL�hd
���:pU�8�F���{/!��L[�n#P���=I8���(O�u/!�$Ζ1	�����#Z���!
D�"!������`�*GA@ʙ8  !��=\I%
B.Ϸ=0����i�I!�٠cXP�$�W������(@�!��S�s���@P�j\L{�-�+1�!�� �e��gY�n�*�"��
	�ș�C"O
)+��9��=:œ�$�D�K�"O�=�m�J��Z�Lx$"OX1;���X�bq�+G�V��x�"O(US��Ȭv:��gJ��L���ۓ"O<��Ǎ�w��Y�hǣ�h�b�"OH|I Ϟe��,�ҧ�?��=z "O&l T�S"1@~|$�E���!��"O(�P4�
\:$�h@��<x*���"O2�!�@�;|Ż�F:\�U�"On�)�Oɽ=�6���DV�|��"O�$�Fc�QDb���g߼�B�"O(��d/�%8ty�w�q�VQ{�"O�aءh	�:F�(�P�"9����g"O<�!�HRwРy'䇈I�.}��"O�\񣤑x>&Z�3yE`h��"O4��'-^I.bx���q�Lp�C"O �[�� Ǌ] �Q�<�x�#D"O��w��+�LE��'�r�j`�"O���!	�p�����M�FPZ0"O�����[��'oUB�^)�t"O�LZ!��(No���&�޸y=���D"O,�@�g��Vș�N��'����"OF�w)N�W�Vw5bg�̉�"O��i��Z$5��@:���?g`na��"O�I9��)s�Ѐ��3E�=�'"Oh݀��\6D�X�`.�/0��iv"O6q7�A�˄	�U�Y�L��"O؀	��
s,���B#.�H�Д"O8���b�:-Ԫ|�V!�Lᄭ�d"O(}�0j
ضt#�I�,�h];A"OFAR�7!���a��
e�<�"O�ɘ��*^���
��!0�(@"O��yAÕ�?
d�C��<9�Ī�"O(tc��ֈp@�X2��.�,2a"O^��$LϪ^A�����_�n5�A"OАK&�NrF)ѷ�:x����"O�9r��C�@P9P��_��l!�"O�������J� [�-I�5�j���"O�Q2��8\��R}�ZX��"O��)Ц�5)t��I�*�?{" �@"O��0u�O�M9���2LL�����T\�<�V�*)֔Гg����L3��LU�<9 E-r(�b����,�ܘ�F�v�<qG�V�}DJ�Z�zg�p�<a�@^z!x@��d�=j-h�� @q�<1"�ӡWݦ�h�"2�8���
l�<qC,
�h���Ҧת"��쓱h}�<�Ѡ��R�'�����}���^�<a,�)j��|k��&ʮ�+���X�<Q�/T6�l��6�w�9c��]�<Iuk�H��J�C�dTh�2�BC�<�ԣN�vu�I���A�,��+^D�<���މ<嬐i���z�՛�dw�<YF��q�� �p/��󎈪\�FB�	7:2z�R������R��@�VC�ɕ"1:���5�(0Q�T1o!DC�I=z2�6v�H�A0Y�:٫ �/D��;�c�dZU��@�p�aW�-D�$��͝
�R8�,ƣ-�\	�>D���B,�W��c�E,m@�,A	!D�09dBN�
2�Ze �:����A+D�LҖ# *���	�$*�(�RrE*D��R���т����d���(D�� �
��P"u��U�3W�И�"O�Y��Y�r�� ��;7F85iR"O���t�ػ?���K�C��c�"O*�*%H!J@y�r�޳F�,q��"Oj!R/�<0�a�h�16�vD;�"O��q.�cN!Rt&Z�u0|�8�"OX���"��u�� F�(
`ܡ"O*�A ��]�F�z��� s��j�"OY��B�T�F4� %[���u�"O���&;d�N#�
�4P4db�"O�U��i̧
�����"�=1h�"O$Z劔�pR�rt#�.5��� "O��whV%�$��J"O���,G�q>d!�q`�1]��Z1"Ot��T�54����*1cz���"O�(��QD�X�ko:Hh�9)�"O6A�#C�8
�T��2q\�y!�"O.�{aMO?m��a'��Z �c�"O���Ië#\ CU>c��A8�"O��j�O�/[�}�&��m�,��"O��3�H��Ecu�;c�\�U"O��0�d�A��	�Aǁ�e6n8p"O��K^b=�&Q�jh��"O�@c��"5�>t��%M;2�i8g"O4]h�/!,Z�5��^�^��d*�"O�=�r)�WxL�k&&ټ6d"Ovm��m�O$T�ED�SJ�h�"O6��QD��>�����b9n/V��"O��{ӏ�UQ�E����-�U�"O��¥A ( �¨@���djx)"O�k��'?�b5�g��2����"Od�c�D\�?�:T���^�[*��"O��
jJ�����HH�쨓"O(U@�K˿a�~ȹ�`ϑa6����"OpYІAVN.����� lM�""OP!%�7�
��g��T���3"O�`[�,�sT�$�(���.�!�݃J����a	8H+d@&�Z�!���I�m�mC�B��h�fB�7�!��
d
ѣӮ��͆,�Ƥ��6�!����&���i�1Y� �Y����'mp��s�Cā�a�0n?S
�'�x����=7\�@0� f�*���'2]��+� 1%X��·j�,��'�q8�&�S��"d�`�f��'̮1K�$�2/��YЀc�H��|y
�',s5B�p�ҕs�
,JI2
�'
v���ǰZ��A�PK��b)"�'f^��ӖSL$����՝����'��僣o�'[��Ô�I��l���'�fIˠ �u��(y7�X�4T �'�fQ����)O/R]��n�'{f)H�'�	����dq��cо��'�����#� Hv`E�P�d$a�';.�B�H�$V�i@�i��<�f��'�b�S�CA�;[t����A�j椒�'��@�IӉ5����#	�<0y��'~����'cR��֣Z�����'<�hC�ЎL�\,�f���f`Q�'}��p%.�!��,XF�ߜzY6L��'���@<5n6{�˨��I��'��i�b��$,��Ί&�R��	�'��h��U�"$�I��AA%M��y	�'�2xkP��? f�Yã��.������� �}sяa6�!�	l��:W"O�1�Q�P�����fٜ]���1�"OXi0e��0�414%M5��	"O(����M:	�D=���L�8�7"O<PqN�"[5��	v'�(sC�,:0"ODP�GgD������2Qi��"Ol\�v,��D4�P���GnQ�"O���5��:rQ�°L�"���K�"O4�[������Eʣ	]>U���V"O`��Pl�1?p	�HB�Qڎ�3"O¤�ц�2�,B4܄v��9��"O*����'�U0�R��d�3W"O*�����1x�v��a}� �"O�80U.�"s���vG$9n�	��"Optc oE0ݶ%���lg�\z�"O\5��Eή!�0��#F��`�do"O
AH��!&C�)Jc��*I����"O�U:#S��ޝ��DU�?�"O��z�1��9�V��Y�Nj�!�dU�<2��Q�T=G<r���\�|w!��ʈh����P�J�QZ��lR<!�d[?&��H�VMn���ӊ=D!��	�2,AaAg�*�ض/W�Z!�d�$ͬ�˧ 5*���#�<I�!򤜾F�|T	"�K�eV(�ѭ�*/r!�N�i��|��S�,$�˰�-o�!�Ѐߦ8�m.9	��Z�����!�$�!6�uy�A.40���jآR!�D��y��P�aC� �ϘAn!�]?:V�ɫ2`�nUI��O=G6!��H����6mR5>	� ����"3U!�Dӹi>�Ԁ��0�,V�Y�!�*2��a���)��\�2Jތl!��M�%�^�2�%�)K& B��عaZ!�$��D P�z4ͤ�
�W*���!�6f,�M�0�W�w�F䳤iQ��!��ucF8���F�,�ڳ�=~�!�$�DF�M�'�܍/iiHR�\�3�!�d�1� t��ϙ�j�f+3L��9H!�dJ8n��s���M���$۽*!�D�:���@!$�ԩ�C��U!򄚖4����ԇTh���H�7|�!�D^ �ő�8=Q�eё����!��B��zu��C�5M�Yk� ߡ!�$�ё��em8�C�e�5�!��1a�L��Ҏ��Vb��˄1'!�Z�P c��A�nA�5�-�'x!򤃘Q�&��6������k�5�!��P�޽��� Q}0�r*��l�!�$D��ܓ��7[u���N+�!�dևde���oA7t�@q�Vh�-F�a~r�>�qu4�hĉ�fްuz�,�p�<ivfX�H��-3��2��tRÅb�':�?�(�m��t���k Å ��$�,D���"âm2�Ô�!)���r	�>i#�0�S�O2��e�2���y�eX�nS<��	�'>l��΍'6�R�X���k�!��#������M��V�&m��E����Z�́�4	סW���$�>	@��)��xb@{�1ه[�<��aR<�zi��!�p�@%��D|�'�8�G�����i�s��0sr-kA��y��Q�R3�@�U&�16"()s�@X&��ęA��(�`U"�b�{(�������  ��%"Oj���OX@1Fi
'dxIsr�xb^H��� ��HU���r�B=d���jtc�OH�d��{�*8cR+�4_�  {%��td!�$I_��p����G+<j�! T��DG����c� �"2�]�	�����τS�<aWj�J�bՋW��;*�
q[cbk�<�ğ?Þ����^�yrSge�<��&A�Xɺ-#���/q�,�A�lJb�'�?���lW�F�qJq�7�����1D�r2�LH�`��P
�vT}1�#.D�<��l3H�&e�$��ޅ�r�+D�L��L�� �B�R�VFŤ��&D�4�ܧ��Ml'�	c��@H!D�BG�@�V�ȗ�(�j�:b�>D�ل@OB^��Y�)�9$Xp��F<D���!��&<qv�EA:�Z��4�O�'�ܡ��AI*{t�� �x���'�U��a��q� ���ƞ�<j����'h�{�(S�;��Ы�.c�va;L>�D��{e����\�%�����E��$kֽ��f��P��%шC*q)�y��;���Ʉ���-���aT]�9��G{��'����a�bl��ۇ*�,N'�b�'�I
t"W����QG��jƉ0�'C��@ʗ�^4z|9��3D��
�'Ҙ\+��H	�����ș;dQ�
�'JF	�A�'*��9C���0���	�'��٠�OP|�XMC�FW��Dpy޴6-!��8̔��Ń\B �r��{�A+�DG �!P��x3x)蓌E/G�!��F�qQ�8���K	Ғ(���2a}!�dDQp����7-�lA��Mt!���3���� �:��ؓ�a׎,g���>�7�X�(~1!�E^�T �(��FX�<A���3M�ԉ���<K2P
f�R�<�'�7.2�sad�!=6`p�n�v�<!G -uf~AKq
��K�PP��Z�<�GFܖ{ ����F�+��a'�Fm�<����+�&	Q�H9����"�N�<��l��M���i$��k�5h�f	J�<�@d@Q�l���JfѤ�iV`�'��'��O�l
�ğ�s� (�tK�>�T4c�"O����$jN
;q�ԴR,JLr`"OF�qh�
�©j�j+q��%"O��;�Ņ$�� �P���Pw�$NV���_��٢i� 8��,�����&v�ȓ[R!Z�!�E���k�*86)EyR�'%�9*���0h�P\+����b��N�<�0�B[{Jܻ$a�P�>�a�^L�<�t�۴J#��q'��!C�\��Wq}b�'*8�0�^k(�s�&Qֆ� �/���]#�\Fl�C��R!	�ȓT�`�S�ZeD�c�Î7��]Ez��O`�}��C61��`��͈�~7� �VJ�z�<iR�P-V�,�ڶ���{Zq�A��r�<�����l	!����F p���u�<Yq(�_O(hxv�Y"L��e�fGl�<��-7�Bxb�j�3��]���Bd�<�@�H\���1�K�;�����b�<�,2/q)Z ��?>㐩�ah<��gĘ\^ڌ��oJ x�q��y�I�+�
�9��m�2ٓaLR��yR�P�+ƴHv/ĝd<�B�mQ��y���|Ŷ�@E�=d�l�B�i�6�0=�B퉪^ �<
&�\�nynɁeJ���y
� ��+���:�'l];,w���"OL='�4���DK��UZ���"O��Y���!���b�C� OJ����"Ov���ߌtqF����9�PY
�4OTc����i�i 	2j 55�	;���h�v
O���6@	� ��p�p��&��d���O��<i���O�9b��֕*�(����g���d"O�����ɯX�X}{Q�[1�L���6lO�Љ� xO<�#$I�77������'\��I�&��0lX%��P�t!N�<�D���>)v@Kdu�q̒�K� �ɇ�F�IX���O
�ɥa
a�mK֫�?1���(	�'��YQ%`�9*��NB1��aP�'������54_�ѺAJM���p��'HJXha�c��a�@M�C��s�'��=���';zw���)��9��C�ɔ�>!p�G�k��p�hG+0�C�ɀW�91PK�7B������Ŵ�C�ɬd�"���@Lg�!�eb!1�:D�d���ԥ')2��\)6�{#B&D�ldd��@?��'������3#lOZ�'W��Dø�ir
�N�$T#���yB#��"TH0�a�]^Jb9����yB`]���q�r�D�Q�����F0�y�[�,Ǣ�B4�՜�j|B���y�O!mp �bĎC�|a��(b�G�yr,��!N�XC��O*����5�yB*�8D҉v�߰a(	3��=�y2N��Y.ʄJ��J*�B`an���y�cҐj)���B(0��� l��yrBP���6oʀ>����b�U��yR�P'52J�$�@�bbb��\��y�����Z!ˇK"�X8!�'�ybƑ�<��%�� J�B�zT�$��yb��	����%vdPP�'�
�y�M �<�fmB6	U�M	�ջ3GT��y����zFFA���N�D�0�z����ye��z�x ���D�puӢME��y���l
���,��p�nY������y������ӦǕ}öAұ�,�yb$@M����s�5h� �3p.Ϛ�y���D^���3sX5���yb���n�p�d ݎ"�8�1bIX8�y2�"�&�[#,�?"~ڈɱ*��y�hؠ*JzI��O�Cg@\0�@�<Y @=��3�h���Q�p��K�<!����H�D�YK�ꔀK|�<Yq�ݟ-mT�Iѥ��mv"i�6�Yv�<	�n��s_Hr"��0Dl�q��m�<QRb�$�Ġ2��ORtP�i�<�wo�K���2��ѕC�N@:�ǟb�<i�j��i!z��.���LDrbT�<a �K2�t�0�N ]�\��Lf�<�7�q�p��Q�J��Aue�<G�g� ����˖mL~���_`�<ɀ��$w�T\��Γj�$A��'�]�<QgL�W�*�e�6s2i+�d�<��ѪBM8�y�ڌnWZ)��nT�<i3 ݙEbĩق�07��x�@��u�<asn>� �T芖=�&!;'�v�<Q���?nz���*��X���Fs�<��Ǐ"9���p�ĉ{O��Z��p�<�����A�p	��EЁwyNh
1"EU�<q7�׬O8:��c޺Q�x��Nh�<� 6��ԇ��h�&ڛ���"O� W�!��9$菁r�t�B"O���fC&Z�8��H�D���`�"O�I3w��]�\���@W:h�^�I�"O(=�7eڑj[x����`�N(T"O:��ƪF�#Z��z�*P:2�"�3�"O(����
GPЄi�ܪ}�%"O�h5��2.u\�ydFQ(�.�9�"Ox5@Ι����ht�>N����"O�\�&F���Z��4t�ų"ON��2eĚY��
��C�e�(����	�T�� �kC�Yn�I0Gl����ڶ
h^Cڰ�h��Q6/a|B�����F��{mZ�2cE��2B�ɼ_�������0%8�������B䉧hP�b��'#
x���B��	=6x�H#(L�H���́1|�B�}��%[Ć4Wʘ����� �PC�		9���33C��i���Ï2�C�	_��2���V���L�FC��L�@9X��o\4 ���T�C�	����)%�X�P��k��XaWC��	f��h�2�í5�4�
]�pFC䉫M�tA���ߖ<��A�S�� 4B�	�m�.C݈|�����D�C䉔�N� ą�XU��`3",P6B�IQVJ5����D�t�3��/v TC�	 6��|���ۣ8(X���HW-��C�I�b������z�] �-R$2��C��EeH���	B�J��yAb�RѼC�	�.�Ԕ; ���i��Ĺ��R�!��C�	Ԓ �$c�� ���\�4ОXD"O ��G����Z��ȱ(�I��"O�9yR/�g+6x��W�f���:�"OҐ��e҉t2zlI֭��8�V�[V"O�(�&X8h�퍠"�F�R�"O�9pB'A�� t��-�fz��@�"OLb��ij��SrJ�4Ξp$"O})�ȃ��-�CK_5��mH�"O��w-
8��"�
;�f��"On4s�$A{��@8��U$B��封"OҤ�ԃ�##|�cSI��GdpaS"O�M�1oK�yF���L�f��"O�t+ďK <�<�rRǆ�}�Lܣ�"OfTe�shs!�]�byD��"OUK�Ѹ�B�X&�0sf��
w"O0M`��^*9�ġ3��G3�V��"O�e�FGr�Y !-Z�$���"OJ�j"�#j�z��.�5j�ݩ�"O<�p��Z:i�Rt�ÌC�f�F�c�"O*]��Gϖ ����!��6=����3"O���Kˤh p;�D2� �s"O��cO�r��`ۣ�7�y�s"O��+�)^��@E��C�U�tmH"OLdp��ȯ2�y�a�B�re�"Oj�"��A�,�H � [�a��l�"O �a�S�ua0p����Z߆�r�"Om	����^@�nG�|p�u"OR͹W�Y�� ��Rn�>т40$"OF$p%��'�p����eΪ �"Oʱ��K�4f��XK񌍹���P"OB�	����e{�a��H@+�P�r�"OP����&�9a�(�1����"O
��ef׍B�كb �Z�Hzp"O�DE�8զ�h�f��&"O� H}��C�+!V����w��3R"O��RH�
v�k��A�8#��"O� � T�^=*�3��G�v-��a�"O��xá^h�������]#�H��"O�ѕ Ҧzy	` ݐ@���"O(��g�A9u���7E�P��0"Op�QD<(�|P��=jtɢ"O�4`G��9�(L�!�c�H�C�?�y��ܼ�D2����Z�؂�Ȃ�y��J��1#$���+ˎ<y�kD��y��R�d�x��Z%�N۔BG�:XZC�ɡ�
D󥄔T��C96_<C�	%�f}���9E�@�4/v*�B䉬�|r��W���ŧ�QG�B�	}|��r���%���'�<b��B�ɀ>.��Yw�Ї$��y*�� O,C�I>+[��#"L��9C��b�D�R�@B�dP�Q�'ĳ����&���2�>B�	3v�>;p�1@L��D.B�~B䉣:�^�5OΣ+W��i
2�C䉓.�.����W����%=Xp�C�5r���k�F��uB"�B��x��9:���T����WBq��B�	�fn13k�:�n�P��l��C�I[� U+WΗ�K�>�  !L�O��C�I�H:�X��	�-�"Ń���C�	ZU�"�"Ϻ%�� -ZB�		1;�AbR9X:.�Ye��� �B��6{�l�Ӣ�W:�:���OW�B䉦��,q6;����06�PC��t�Ұ6iQ65X腀g��%H3DB��q@��gU>9��R� i���"O�H�u.�e"\�2�R\l��XR"Ol�I፛�
�N0ҡ�ٸbd�2"OP0�,ǉA��i���*
��!�"O�Y�qGW5j��L+�(W�f�K�"O̝��`��|_
D�G�M�"���"O��	�G��PU}NV|iT"O� �S/�<^�N�.�536"�H�"O\�ԌX�5�)걨̿	FN=!G"Oj��'�Jՙ!�1X��"O `1`�|�A�.0X(q&"OJ�R�oKz����rBA�B�	5"O�uB"���	��� �b�K���@�"Oh�5È>P�^@�����Z�"OJ�{�.[� ;(e:�G�d��ѡ�"OR�{�
2��ɶO[��Ƞ��"OL�2w��u��M�A�}���9�"O<X�c���p*�dӥ	Q�b����#"OV� *�&���XH�%8�̠�"O� �Î�V@�%��AR0ϢȋF&N =��yy%d����|�ºi�dx��A�3��Ě�h����S�́b�I�J�?Rz!��	�+��䉣�6K�p�/��
��9ސ}kٴ->�U�a��D7O�|�!�?y*łC�N��8��ɉ�03���sI6|O�d*cCH�?�ha��Æ!�Ƒ
��8��KA!Ӄ%r�}(�(��D۱>%hB�XF�3�ɦe�\��s,�y*����Q �xc�4jTH��]��aJ��N�jw��U�>5o�GiN���� *߼�� #	��4�@�T�-���;�O�0[0#��4�@�Ɇ�D:i&iّ�̲: (�*o�@��޴-8Z�i���"a�VZ�ල`ԅ�+��SӧDi$�ǁ*������k(<�sb͇N(z@���ƥ1u�0v΍;�^}�ǵ]�plC�i�ȉ�#�)
�\찦kXNh��q��]�u6Ա���Ω����$S)d���
�To�����C�J� �(=D�!V��ua����K�l%��Ơ���$ɧ�J�|��x���)`��P�Jz��𡧋M�n&��=�	@HF	��fO�B�p�[`�Il��6y�R�K��iH��8seͣ#�h)�Ǎ�d��=�Ƥ4\�$��X��>!��K���}X���UK��"�ұ_�z�	8|O� ,���k���(M�@h@�`t�D(�^���/
� �� �N�.�����/�6q����~t�t���,ջ%��.M��;S	�&��'��̑/V�&���o��u=�����	?c�N�iBi�X��@	�*��&+T&��<���s0�ĹP�Ƚf�X�)2��"/�~ك�#�̈́�9��:.�E}���
?�qI7t�����)�d���U� w�`�u@Θj��i	� k^�v�HC�o�KD�8!#�8@8��?y�*6�#W�/�w��<iSk�1q�|t���O���!%�ҩ1�1[�mǗ+�⸊7hTf&�
�Ҏ	���?�Ԫ�F�0��`@J�VT�+��'�&��ăC�<��'X�%=�}�Q.�3jD&I�`	�ot��R�[%�*ۆ��F��Gخ%>��C$b�2d ���o�܍���I�Eb����'O�A��!��p�nģ¢��J��Ԉ�N�(�ye�>/'��4k��k�����W�bB�1O����v.�<!�Mǿ,
���т� <���.H&c��Ӎ�dA;Z8TA4����)�B$�}����C�dd��55���C"Y�m�<\��'�,l;�k�?(�1��j���v@�T-B�1���O���P?�	1V��r���:O��!���f>��[G�˽.�ⴻ&ڝU2�5Y���>w���Jλjd�980-�I~Xt���3L�ȴ��i_ �|��T焥lq�,�ԯ,<O%�Ӧ؈o�*�P�d�'Y�h��Ѐ<e���Fi��b@�d�U�6>x �&�i�6�&T���Cȁ�4��m+ �D:j:�9S�
$ ��S��'	��{��4(l	�ǂ0)<�y�&"�!yh}�B�~)�rC�%k*9 �O�{!�Y�0e+(�;� ��+�<4��4���M�+�S�+U&dk�E}B�K���A��\}j��7�� ��	�5.L(I��#/ے���lJX}B��+EE�f$U�`\�Ԁr��)���0�T��v��y�7l�c+8�K����Z�r�	�`��k��^((��Ȳ�k�;u���C���2�⑪���O�Ąg��L��B�:3c�[�I�L0��YX������5h �k��)<O.���΀}���kBFȌk�\8@�#��}�� ��I?#l��ȶl� 18�'��z����&	�n�N��|�bũ�U�$)
Eh֦۸�dq�4g6�O8Ł%'=p:�,�.m#3�Ϋ
��J��|"��Ǌ�55����O�'�b�ᡧ��~�*q+�Ϊ	��(2�מu0Ĩr�N:������G[rP�0��P�'�6�Җ"��@�a�aM�$w@�ē�NQ#y*�Z�Mt��X)���x!ҧ��`� i	�j�E����+ i3k���c��|� W��K�x����
ɤ��I37�D=�h��H"���wor)Sc�}�F��×0Ob���E�S���O�\�p���W�g@xQe��Z����5I'<OvD�fآ/��h2NƗl(��
5Ot}b���s6�tk1�ԩ}0��xÌ�\�da�
5�T��7��1�YцM
,��M�V�$.���O8� �Z�iK�-sԐ*�o� 0X Pp%�5r��B��L*5�4p��I�4ϧZ�,�1u�ށ�t�Q�HA�K��#�����(6D�Ȳ&h�y|��PV��`2�c �O�l�"Y�Ǉ��b}XuY�C�� ���I�'{{����5�	<���YPL�'E�"��Eзl����^
]�Q�O���!x$$�&S!��@�R�:�����ÀAO(]Z���
"&E���'6~�A%��"p�%�7���"PH�"��D�	Qb�P�ĨM�x��O��lF��uG�E�9���zr�uX�9�F��y�e_�&8^���>)^(ɢ�
_�	J�#U�������(3�� ��_!'9>�n��
�4}��"J�gn��@�ס+!�[�-_�;LD6����#٩$�����8S�BtC��^�_6��r�Y?����޷2*Ը��Y{���@�B �}�#��C"�u33�F&XhM��䛦NXL��2��`|��EV�8H�e��H�.I��Ι^l|�R���a�D)��2 ���2%V��t�S.�� Κ�<,>Ԡe��9/�ܜ��Z+p�Ql�k��U��)�27w�@'�P��iI26u�D���)\�l*\�U�
�fpe3��6/5!�dӔ`�^��C���r5�f	��.!��J�`�\��a��= ݨ ��
�.ha!�d�1{���D�B0���CZ�c!�D�`r0t�tLJ������!�D��P����7$�&o�dX��P�<!�dD�Bx�f��_��bg�WU!���H����V 64�p�NY�|�!��N��@(1�Fě^,�%Y���?r�!�D��w&* A��>U�� L�i+!���3(LD��7��&�Z��Z�9!��
5C{�p��UTQ+@�Y�^���'8�=J�iJ�Z�����ɟR�r���'R,@���Lk4�R��߬L�~PJ�'}D$��b\�<c�p�m^�;��"	�'���e�(����_�;��	�'C���d�hR6h�Uc�?���	�'Ӂ����U�$.	������'�<�!p�\�Zg$�`TE܁-^tXK��� �it���G�X	r'I�R'�hJ�"Ojh�$/֫Ul��f��U�G"O~��#T�-0-��Y�Pt-��"O����F�>D�#r'���B�"O�@a�kE91�d�e�8�0<!"O���.��dr0�bec?&��ARD"O�[��[	x���3ɴy	��B"O8=�� �`�B��b�ɏ�J�:�*O��3t&�8���`#U�j��l��'�֤�w,F>y�X�Â�@Y�e��'Jd:aa˃)�ް0a�R�bvH��'��e�s"�2Y��(�����[!
�j�'HP�(/Ƭ�6L>]�0��'= Dr4꛵|1���VK	65+43�'�y(�ѱ�[a.�,�� 
�'˾mJ���aC�HYv�G�. ����'߂5��4�0�h�/U�7X�1�'�v q�Y��d���mW�<�i��'p�4A��4Ҵ�5 Ad3���'�<�s0�]!(� L��� )h�p�'��ӆHcVN)�E�ڰ#�H�@�'މ���XLܔ��H�o�6��'�������H��I��Ɍ3�����'���·>_b2"�B�.����'��	��+[���� #�s@h�[�'���� \]��� �.=���p�'�%��`޽~׶�h3	H.osbu��'[�����1�F\�B�MT�4J�'�M '��f����rE�1l\���'�0��p��
nR����+����'�h�ړ�G',٢`k��KUnY��'�8ܳ�NO�l�j�s�#�8Y�!Z�']B`�W��*5�-�FN�Yװa��'�$�)cNE
t�fY�v���]~fM�
�'�~�� DĄDr�/�/�h	�	�'(�3�:F��q�J�P�R�!	�'��p@adR�W<8�-\fV��'����������O]�
���'�.�1��N�/�l��.sސ�'?��J��4a�`#���z|�	p�'�A2��R�4Pj-!�(5t�&�)
�'O:ā��N�y�+ �STu�	�'��(0� 4inM���\4W����	�'�"�"���+>b�My5���ʓq���
�-ރK<�i�%锊+��-��0�ʬ鵋^rd9�0��=ش�ȓe	�Q��͜��=�Eć�X������9��%]�?I,����(=�i�ȓ"�����"��@�B�	^�.�Ʉȓ{M�xg+�2 �Ơ3CI$�X�� t#�Fվ5
\�,?���qRlgB�93	��pe�O1|����)K�m)���?%�p)����ZT�����e���s��#)w�цȓ4��� �g[@��SM��l���ȓW:V���#!����!˿p}���%�r���c�?8�T��p';; �P��d.���bJ�7,i4x��`R�Іȓb���[?ez�+�_'c��M��G�x<�DO<�t�'�A	J�Vi�ȓH2a��Qt<D����t��=��,��x��A$��$�KKy��P��1䡀'z}<���5�h��|�X�Qf-W{�Р�mK:x�D��S�? 8�ƃA/y����C�0A����$"OV�@�7pErF�ԑR�~��@"OD��H�	�h�ڗ�!u����"O�iك��9@f���풞���{B"O�m�I� F:T:����;_�M"O~�1q�L5<��E��h��"On�Ap �L���q��3��ie"OH�]��z�K�4���E�լ5!�͟z� ��dc�=Smm!�dـ*��S��J�/���-�8�!�D�%�8�SA �����,ʩ@�!�D/9P^x�SO�<d��d�V+���!�d�+/?��٧�H�I���2�[�!��"f�j�ɦ�G�2�T�W���!�D�?^ܥ@ ��&�c#�-K!��G*��I��xO����Fځ7!�ĉ'XJ�H A[;!80�S�&�S�!�NJL~̀�kʼ|	� �C	�'�!�K:>@���ֻc�~��� +&z!���g������ںZ�vu�R- �QS!�Tx�!z�(Ŕr|Z�y����'2!��� -��pڶn��gj���A���[�!���6v�!�g�G�h1Dƀ8<�!�DR�,�:��k@�ڊ��b �'�!�DQ�]v��@H�Q&���Հ�0�!�ğ�JĶL�@&��df�i�� .b(!��<7ID��A�X/H���$�!�V�x�BX` &��lf����JP�!�DB�F���B�:f��: ,H�e�C䉼X��Y�R�����ª܍n��B�I�7RDӪ��(L�QA\��qW�*D���f K+�I���Ȫ%����`,D��T)r
0j�="#h1xE�,D���
E�h��y��-ք)AR�b+1D��p��W<!GF9s�╉'�d}ys.9D�����ũcX^�I�z��L;��4D�@�c�X������1d��$#��2D�\хB^:6� {Gˍ.0�$�2D��*A��K�IӋ=Y<0���ޯo-!���1_��� �b��aچ�^�$!�$��@DQq�	� � 5�h��!��R�.z�)��ٞ�L�җ��F�!��?V���+6���f���#3,תs{!�R(rX�-K�H�
�F�)�L\�v!�T�|�>Y���;��9�W�O7|!�$ÃD2ٲ�5%�D��L%Y!򤋂Y�#&d��| ęЂϷJI!�dۮM� �`���c���� �+'!��SkxU02j�_��,"�)�O�!�-G�H8ꐨ��N�m2F'�2M!�_a�4�s�*��)ª�����7,!�֯9��T
��J�/p�R�h-!��O�=4��A@P�,��a� )
!�A�wCb�B�����5���t!��E %Qh<1���/���5�!\ X2�FB)�%�J<�''������������-`���x������@�
O{�!�$\����t���h���J��󄞽O���4�T�႞,��� �`���?�;d�����zs&A�t�$�7�=|O8i7�;rEԕ$ʊ'/���2哪 ��A��і4w�i�rk�+Q�Dޔ:uy�g�3�6*La�6'[���ez���&.��c�,"�IK�eݦ�[�n�
�'VϼImړM���ʅ&	4Y�q&��Q��!�Dk/_o��`�E!�O�d�1%ėu?�=fA�b�^=�͌�ZPXg��!b|�1�ȕx��`�q���M3��Ì5��BB�Z��i�p.Q*
��a1�� x�����=D�xS��܍H��S�i��l��٦GY�d,���TAN�$����Դ&����,���,���l�\a3��O2o��� ,}���Țm%Q���3��lA4�'��	`lD�4V
��DE�/ц����g�V�9g'�#C��DJ�-�N�6�`6�UpDZ�j'׊����s�㟌�`�ԇj�rI��g�q/>��#<�I��n������$x�竒�=|��c�	V���i�*ѻf��Y�m�/{P�E"�*���s�����G9|Oʝ�w�"K�b��d�@4v�����N��z*����O_`+WJ���ȕ��٠N�|�ʔ��p��옱��� �'��6�5��d2�:e��"O�dS�-�OOF�W�ϊ?���+�e�^��T$U>s����AX*j��pCƍՏJC\�k� :��ʦ+�6g��@
ҫA,�ڐ��AZw�� #�'%�d�ք�?9���Ӊ	���}( �F�(������]c���Ѩ�>����+l*�bsA�(086#�T��nK��0�҈e%�a��!R�\����=� )үrhvY3�'F:�XSAnB,�"�2G��6!zdp��`ߢe>݃��2{���B�H�*�2&#��{](!��#�,S��Do��9䢑��H�)R� �d�0�HD! �y1��% � kp��Ad��aT��M�$d%`�|1''��-�V kH�/,*��C�'i�p��+P�:�ye�L&b�#F�6�\�r�)�T���Pb&�ba��U�"��/� m�-{��~
:gW�[V54�ҷ�&�c
�@�&aK�	��#u<R�
��,-�@��l�	Q6��c �(���,��@�c�= �JT�2�-)$�d�rL��U?�'1�h�n̝]��d�R:����rb�rܙ�H�>��q����'q-���AG�h�\%Q���;+~� �ˉa����!��r�F��2�֪	���0�9<OU�sn_���뜳91�hK桑<��9#��?������5ba���^1����[��`H��q�~Ѣ $�Ш��,�N����O��iu�/!�܄���։[���'ZQ( �r�͌��~��UX��ba)בiiNx��/E�`�k�w�ubƕ�3��]�	�:/0r���t]f�����#+NFԢ���0�!�7�^9��H�VV��U@=,����55,t���T��㲟|��_#i���7�5/h.0���8�hO����5�����mJ�����nJ�x���dCVk	���@�G.@ҴV��"�"��e&�`b6��p���牪��r�ޱqr`	&D�}�^�ɋi�+ c��$A���F*�DJ���; 6�8kR�I=o�F� ���v�I��(h���"B5��C�/=8��B�2�[W��,m����A�/([�#��J�q� ��jJ�0.��"���c�ꃮi����3K�D���о�¡�L eo�����e�(�8�3F*Q1�-D/T���rϑ��^�q��B�P8��E�/+�`D�0A$uiDͅ���v3�e���.�(<��
V��F��·D�l(��ƪky&l��ki��0������7�T�D�Z*�j��$4�����I�zX\�x��%<On��e�W�t0�X�B�D�����Y�4	N�Q�x���H� n� E��E���y��W�\����n_	��<��E���}�#,4���0#�0�%�CoIJb�d9��	4� �1>��$�ĦU!��#1�!ϧJc�l)�Bo�I�d�''���D
ƫ[���s!D��R��������V`�qbfC �R"~)��M�)�B�9�Fܥ`9�������rh$�	�e$�PeQ9W�R��dJ\.0���)K��ը��Za- �h%*DUBe��&"oLvmX�J��P���*�E>h80���'CR)�իT9_��й�kH�z�ˌ�/v���j6K�(q�
i�Ï�	���j�	���
-��EŴn�����<�+O�P,d��j�608��BF-{���a�|��pC�H�`�Pщw��*���Ȅ(��jȉq�RU����y⌙� *u�J�<Pj�(�n��6ɖ�9al@ R����C%V�!︕S���FxR��2Z5(P�aI]0-6Ґb7&��>i'f�u�%��iǡ{�(հ� Z�#�P�+��Éu�z�WHҌi���	�D<�Dp�+�`Dዛ"����$ǠW8�	+��6G���]�@X`p���	U�4	��V�dC�	�$X�H�BiE�%�pS��z�~�O�`s���{�|�G�$��0n\� �/�(���O�-�yBkR&3ݸ$Ip#S�{��hH�yKB�*,�¦`@�q�"��y�X�K����Bc8��&�y�2`�Mⱏ��o$������y�&@���ȃ�a�<����O0�y�j��g��m��'	2:+*��(4�ycJ�=��k�*�9�A%��y��ݓX��s&��&(DH1
���y�n���ѵ��./�� ��ޟ�y"#R)2+�EAE���j�����
��y��f?�ݲ�	ăt�Y�6&��y�f���>�@1�͝:.���a�T��y�  "7�J�as.Ђ"*�I� I�y��Cp�Kqd�&���( ��y
� � �ck��p�m�%T�U�w"OL�R��Nx�&\��72ԣ%"O��J�EA
2�(y�_4zc���"O�M`R��32ktE(%���0��"O �C�l�)������38�J���"O�%Q�n�l��]H i��1ˌ���
|�DJF8&�P*r��(����ȓW!�ٙR�M�Q,�U���K�V���4��@��%QV��3F%9m�T�������m;zx�Ռ˔L�@���ڊAZÊä>]j] �NY6���m �	����,W��ԫ�L�@ �ȓ*sD�'f�d���N"�8����SE�����A�\$&k��ȓ�vJ��[8�MH4#sL�i�ȓI��Pj��������5J(��ȓ!�JqQ&��3$j�`�"�1f�
�ȓ'ՐT�c�ݦrԒ�r����,#�	��w�DzG�VB��b!� 	�QE|�_F��`#�	�WP2�a���~b�P�c<�@�(vĐ���pF7Ml��PSZ�� �O駐~�o�iJ�M��a4�ч	6)
�	�m���	_�i>	oZ��ēT\�r�ɜ�g�~�V�`I��iQ��W���s��|���e��h*3�3)���xp�
2al�Xf*�f�I�2`1����H)����G�\E��A^�a��h�«�"�MKٴW�t}��Cر1�������h����3j�m���s4�Q�g�\��Z��Z��Gt��zq�x��	C2S����A�(p��\ؑ��#=��D@��
7O�E��8"|"���K�%�6nP�l̚����hZ���k�j≧�'��O��b��u���Ք5 �9���6Q:�OhD�c�?��"u��*զ�4�@���?lZ�"B'������D��öEȠ���?��O.,���@�9,0�j�V�f^���OZdn�[�)$��E��aҮB��|)�\�!:E�iA:�?!�)��ʑ`�3}��$,�|beD�<Y�g	�NX� ����VG�����ē�0|Z��Cج�"$^���Ƈ�u�m�I>֧�Z>�����:��H�gN#B�<M��j�[�	�B�>I��J,��$[���t� �ԇK/d���T�l��k�.�j�9H>��P�(���:�fP�2P��ѵ�� =ߌ��3ia#�˜]�䧈�|Щ f��o������P'�`���G
a�l�f*J�yj�IH��x�OU4�j�#�0E��,둯F�zU�܃@e�.6>�'T�؋�������eY24+��R�ؠ��5��R�O���@�F�yР��5���	¢W�T�@p�Ζ̹C8OxqCe*tӢ�0����ɮ��9���.Nx�	��6GL��u#NY�eoZ/3`�����I�Y�l�E�dӟ��iգ�N^r�Lܝ<�\�1Cl�x�*��#��92Q>����� $��\#�J!�Z�E#J�h0k�Aa��1|�ze���DL������M�y"g+U?�%q�f��Q��A3�$��y2���;]���,u��pS��]��y�OO-�T!ڶ��JH00	�'K����� T�����a͸G���'��L���F��bȋu���)�'Y����AF8�0rуE*�E��'h�*NS�#�j��D�n�D��'	n����,4 X�0Ћ��{�|��'O�(�ǁפ	�DLYg(> �b j�'ь	2�GѨ;��9�g��/^���'4r�jJ�d��-��D��W�D�
�'% ]��j"\D����z�Dɺ�'Pn��愨[�8��������(�'�(F�ѓ,2�Q�O�+!^�'_tp�쉜@R �"U��Sk(4��'OR�Dl�3E����t�X�;�zX�'�xY���˵}����p@�6�N���'̐8�O�L�H�0UJ�2=&А�'�J]k�J]
5�j-p�DX<�< �'�xu�f�r�b*�6b)r
��� p���[(���2�\K�̀�c"O��YP*�(��9�E1)Ӿ�
�"Ov�Ҵm�TS�q�ĮT����q"OL`k db�*�WN�+���0�"O��I���	+�!!�ۻm�T�q�"Oё� ֮Jx�����F�4��{�"Ot��P%��k��ʣ7!�ң"O��!�kԄe@�D+Ee��fo���G"O��Q�dZ�|ufAU,(K�"O �-�%M�\�To^�2��Y "Oڑz�N���!���1���0�"OD{0j�>{���P)�T\�ȓWc���Z�X0fIӧG(���~����6,(���ǋ�nD�ȓ$�<tz�+�*�8�2#�
Z��0��#Ü�``e�P-c�	:���ȓ>��AZ@�M�`AԫPNft�ȓr�0AA �R ~	n�!%�Q�\�ȓz�΄��d�hf�p�%{Ȑ��or �b��|(�!e-��a����-�А�qH��%�P;�iR�QF^d�ȓ��UHW0/~�bn�� 
|q�ȓ~�xd�䯋)uI�EFΖ
܇ȓ.��p�� E��9%X�#`Z��ȓ)�3pL�5�ʘ@�j�&��Y��`�h3wk�:D��)8ڙ(!�B�ɾw�@�gҮ��S+�T`�C�I:+l)���@6j������J
,�XC�I�g��iÅ�Gs?~p���^��(C�	����-�,*�{pm�7(VC�ɷI�pj�ٮ'a�@�Z;�|B�	�p�Xlh��ۮ, �+��U�MOBB�It�Հ��ˇRT؀fƁj B�I��`ˣ��&D�L�q%��I��C�I,�*�+FW#pȩ��6��C�	>k�
,@0'�:w�4�#`Oт#��C�I,H����� %��!�@�O�wbC�2G��܊'� �0�҂�P\�,C䉗j)�z�ϒB�V���jM'J�B�	bF��Av���\���� �~C�ɹ�$�D-$5�9؅GEN2B�	ke�$kK]�pјe��`ƛW��C䉳7��XA�DL��+EI&#�ZC�I�0UI��ŒOWx(�%A'W|B�I$m ���GƯ/a��Q��)f-C�ɰ&f���6�A�C���Ώ�r��C�	0f��L�2�t1���Q�t��C�I�����Fkz�XmA�c��B�I�&]pd�p�BT0�K��n��"O��{�˗��\8A��A��b*O��`wL�|�R�ӆ΢k��pR�'*�ZvȞxp*�A��V�dH>��'𨹘D��Wq��Hr�M#r�h
�'b��R�RV1���3n�>���'�؄�%�vp�}a��isjɃ�'lR���cҠ��:6M��c�>�B�'U^�#�#�+	�
в��M$c��}S�'QR����:pF�˅b%Y��B�'۴�'I
�k�`�"eh�WRQ�
�'�6�F�
 ��műpvxx
�'5���eØ�s:���W� 	�Y	�'J@�Iż(� �!�}Y��	�'�*8T��p��K�-!�"�	�'%R�5�˯G�¬��ʌ3n����� a(�n���������-�n�s"O؁r��F?c]ꉀKA);�"O8̺FL�fD�1�Z�#�6��"O�a�WD]� �vJ1,w^S�"O�A�1��+0u$3	��7{�<��"O8P���Me�z6�аrd�� "O(����פ}��dj1��"O����:+V0�`d��4�
"OX�B�o�=�2��MFJ�h��"O�47���qX(� g�EfgXp9�"O���ch�����eQH0�"O.��w/;N6`8�ѾsT@-pr"O@�A���S���N�U;�DC�"O�)�`� iG�ќg# ePa"O�-�F#��tkX�A�Z7%.8T"O
�3C���j[����=�"OP����iTP�@�	��H�rl""O��#�P���0K4g�+f���"O��0�%/): ��%Y*m�H�u"O��ya�E�����P;��t�"O���g>g{ ��䞨-��mB�"O4� *R�
��4��x�XR�"O��F��$G�����}�H�z�"O�ysBQV����2�԰D�8X�*OA�$h�ߔ�y��A�2�~D�'��x'�ʉT#��6�D�*xR,��'��9aD#)�|�g� �Zޭq�'`b�IT��m^u[$EK�eΒt��'�Rd�P�f�ꠉPAP��K
�'�p���L�/�(1@'���@|�	�'��ȢA�5![��Ј^�"��`#�'ԥ��Cȁ
��1��%,!/Q �'O��b�K���G��9pvbu9�'�R�q���\�&��L&氈�'YeAMt���F��s�t�'T"��z��ݓ@]�y��X�'I��1cG��:8��f��k����'����1 �Ul4͡����Z]���
�'��@�P%�-i&1A��� 2>X�'��h`@A
5�6Ԃ�aO.��'���貍7xZ �烐UNɘ
�'�đ��(S '������+	�v���'�1�c�4A��mAsHRwA
iy�'!�
A�σ���2�F�i�R���'9�m�AǊZ|
5�㑔uߤ���'S�D���0<��P�	B�`e�|��'�:l�p�� �XP��U=�4��'`��A�mIP�ݩw��Op��;�'�PKT�ӄy������%/ 
�(�'=(��5�A�<�0Ȅ[ �h��'f̀C�'(�РI��t0�H�'.DX3q/�U�NQ���3-�|j�'�Z��aÀA�b���g�ȊQ:�'�uA�H->��䍤�%��'��:!�N��рgj[�u��P�'� ���ȟ1�\��q�E)n��0�'I:5pAk�f54����Չ4.8���'8>as5i��`z��Q	|pz�)�'9ʩ�D�+gN)�q��w5X��
�'�@ 2���&9�p�a��t!|�	�'l�̫&I�j�Rr)�$c�<�	�'Nb�H?b�.���%�>`&�p�'t0r��{����W*��L	�'ˠh1�N�Q�-��\�� 
��� ���bC����P0̱TC��Q"O�� W����X�3F� &h�ʣ"O�5`� 
/�`�0g!'�n�9�"OL̊5�
�v�L"�� �Ht�"O��RS.��vz&����	�"?��s�"O.0��	9�{���3
�xq�"O>k L�yuX�+�I�?�(��"Ov �Ɔ��f���acN8_��j�"Ot�)�HP��*��ש!M�� "O�}0ӄZ�-�R�;2h�F�Ha!g"O,lX���;%@�q���Y>�q�"O�(K�o��i`
t���W%��!	�'�vX�u��=L"N��BS<e��p�'�@!��#�g*NE�eʼt(��[�'Zl���L�Po �׊O�t����
�'����C�G�u�N���4n��	�
�'����P�2 �nΛ�^�	&�}�<��!��z~`�$�]�ѫpf�w�<�W��Ow}h��?b��E��@Z{�<ɠM�7r�NH���״4������Nx�<��"�<aY n��<��F�w�<)�i��VJf4;���e��
�!�D�"څBg�E*)d�@f�!��Y��<��pMC*Q��Y�ӏ�;[!�dK(v�rp��� �.Ɩ��G�@�N�!�ς�<�9��ձoO�@Pg�d!�\2U�� ��i'
��`.Πn�!�K0&�-��lp�e ��G|;!�	u���#�/0G�`y���#&!�$�kQ�G�Es|,S�G/�!�D6N"�=jT�ũPgʸ��N�$C!�d_-2 (�q�IB��nѩ$�!�UQި�2�9#q ����!�d�$<�`��r�_�;="Ո׎�>y!���
#ht�tH�1g2�8�T�	�8N!�d؋mz�Z���24*�q �C�d1!�ٔ!�A�eÀ-�P5[`�S�!�ƥ	3��G.�,���B�Z.gS!��϶4� Q&��CWFK!�
�0��Ei��Μcy�u�a�Q�`G!�D��*�D�H#���qF�G�	�7-!�d� �~�,村�ǽG~Lz�*O�b�/}�M��T:'Ґ;	�'Zp:��p��K@9��f�U�y�)E�p]aGC+}!���@�yrӼF�U��Ɔ�>l������y�2obp��*�,{��`F����y��Q�D3N�@�M��g��e���Y�y�o
�) P  ��   [  Z  �#  .  �8  �C  CP  �\  i  �u  R�  k�  �  k�  I�  @�  �  _�  ��  ��  (�  {�  ��  	�  K�  ��  ��  P�  ��  � 9 � > � �% , �2 m9 �? �E EL �R <Y sa �g n Pt �z 3� v� �� ��  `� u�	����Zv)A�'ld\�0bJz+��AI�/C�2T0���OĴ�����?Y6�S��?� ��g+`�J���,�V�	u�>RG��@Wm?x��$�۠Su~��@4�N�Qf��IT�j��#
6�xS)3��e��N��>4v���H'9Jz�3�&^72�R�Q9��)��O��`���R����/b����F�A_><��S%ý\���X�JL�y����DA��!0`�2
T,ao$WA�A������I��Γ;�|9�JL��x�O�.N���������M�+O0��&u����O���=CH�c�P�)����w	��jP��d�OH���O����OJ�D�.V�d=�m�AOQ�����K��+pZ���c�"a�%P�/�)�y��<�6�?h���$��Tb�9׎�%
$p��G͗mA��'��!�I�% $|�աA�T(�Q�g�@i�v�ٹ�����{����9�M���?���y�'�?y,���]6,l�"�WOd5+�I�?����L����4����w���$��% v�H9�MS���a�� ��Gm`.y:q�7<�z���DY摞�:�%ö0�>���[t�F�xai�m��` �Jq�@�Z	�(�qL�tyzq�@�����mK�N�H�4v��Ve������|�׋\��M3��ߩH=H�ώbBN��O��M;	��[��ՙWLةLx"�	cHi� �t�<[�7-@ަ%"ܴJA�4��8M�����肪'^H塒�O�B���h�(v��v�k�XllZ�!��mx�j9F.T���)	F:��cgIt���t3 � ԃB,=��X�n@�H.Y�ش���o�2��$b��aP��!,�Ѱ��=`u���c����02Rm�;0c��oZ8wjl2���%Fɰ�r��M{O���~��y�� 1��ɬ(ֽ8��\
=e���oUK�p�����?Q���2�';_\`�4K�e�c��SI+��<h�u¡��'�^�H3�O���� +���D�O2��̀�ܱ󍃞�~�1�@�IS�:|7 �kE��F#����'�E�B�5"�҅s�
��T&0��&�~u󃁛=s��`p hs�����+y\�=���ڟ��ܴ#��I�d��f%T��G2gz���O��d?�$�O����O"��f>�R�lG:�
U�7���H*�!%�O^�n�$-��]Ad+�L�"�+Í�Z�ڴ�?ᆷi=P��aAdӒ�D�<����B��-|Z�)��ڵ�21+W�b���C��?Q�
�(Q�M)��ӧVZ%X��i�ʐs�G8EJ\P�M�T�<��'�1?�R(��1���{ĭS:bޘd4��2�����#q� ��gϋU,<��*V��d^�r�uӜ1F��6�Fp` Eٰ�l�)E��>�"LS�'G�O��r�^�r�F�(�l��J_6���T>�hO����;�4�?��im�� <I
��� ��<v�1���8�B�'��ə|�d�IџX��şؕ'H�)�ք�99$D��Őc;���@�/](��۰�m���Q���:~�ʧ	�O0���޼?�℻q��U�����!q�@���(�M��1�:%%� ���A7����ȟ?v`��������-O��S�'��t�?�O�Rˋ&$f�"0)ӼJB8��v)�O��$�<q������I 5�tY14n�/��j6��-#����O��nZ��M[J>�'�.Oz0�^�]��3�AKUP���f:O��d�O���]�;���?��8b��TlA�t��	
�
>�Q�a!R�"���H6L��� L$6��y�P��5q�.�	�!�-_�@q����I�RT"�DPR6�Z/�ў�zĢdb61jd^5	���{oW(W�h�d�����d$�	`�Z�	��3�)�I_#K��	R�	�$?�<4E��S�ܩ�"�	�}��IP��ן:�4�?Y��i�B6�|vB���f�'bB�M76A��҉;Wx��Q'
2^�'y$�u�'x��'@8���_�b6��ҡ�P�n�\�"	���13�� ���0K�ax�m�Sh��I�
�X�[��F�h��!�g'�)L��ث�N&�`p����k�'wP������jӺ��^96��-��D�@Zn�"dȅ�2�˓�?����?��'<b��Â��O�Zg��hذ-�?���h�mZ�{��Z�]�]�± 匴I�4�?�4�i��i��i����<q�'�
��HY���  �h(�
%�ǟ|4���?��c�3b�<���坔�M�T�f�2�?�i����44���(@"�Q��w~�
Ře���Qe�[HH�RAG��n�^���.�bl���O��x�S"����C`�R��A��O�)���'�7�@�[�'E���(Ll���[ҍ�_�`'���n�	֟���gy�狝u<����Q��e�D0�"=���I�i��Kl��� 7:��É�9��rT T�G�j5mZşl�����q'�Q D��ȟ��Iԟ��;7u��5mܐuX�z�R~��Ҹ|����M;��3�\��.����?�q�H`�Z��#z��[��Г&�*ݰ'��1w8��k�	�_�9P2�����Ƀ��)R�2�.�E��Q�:,�F
J�>���0�q�Ұ�O��C�'�1���'���	,Xn qZ'
E>)���ǥ]��B�'�r�'VR��>ف@'(�h�zGf�X��mi`�J��h�	+�M�u�i^R'b�*��������|��٧b��a3GFǤ!�,�BF��9Ȏ٪dT��?	���?���d����O��$|>m"E�Ԑ> �(�K�&��~�Tx�v|���R�day�G��0� %��&"�Fxa!����Ჩёg40�b����"�Irl��xF�4��'�ąp�˾6���[�@�:lᙂE��?I��?Y��ᓛ���!��T�F�e S�|I���$�I�Q��z�_�{�4\3��!S0�Oʡl���'̢��/e�����O��b��X�-��4h�j����8���O���[�Q�����O���p�i&��Q*y1��J>�P� <�A��+W&��Ja�_d�YHP�=�AÄ	Y�퉹F*t�EN�VJԀ�"۰1�>E�V��u����_)pł��]�^��\�]�?A��|b��)�L�6��%]d00��y�
�5Q�x��ؖ@.��X�h����?D�'F>`��m*5(ЬΩs���H>�thD�|���'�V>mAiǟL��Rfi�d�A�]��D�k�B��D�I"9{E�PM��u����R�FH�;����9jJXa#��7p��q{AM�3y5\��'�����b+w��pYd+-��%i�*W\���5�HW�tiR�}z��0"(�0iX���2i`~�P��?���|��ɜ�eN@�D�WV`�G�^p!��Ȇq��Aۇ`��QN0��� I�џ< ��iWO�8qBW�@R/̝Bm�1fAt7�1����G����'D��'��	�j.P	�ƌ�M�:��7�ӑ<�p�1���_�Z`�ߴ���[��.��Ɇf�:���d�]�N�ཁ�Q�|JbI�P(� ~��׫R QR����#RO̧��h`����?���;�N4j� �޴!�I�u������g�I�G�`-�VL�1<�I[͚2
��I� �'����>ac`�N�2�Pv��'mVMH���埨�ɱ�M{`�iɧ���O��I�v�Bq�iY�R��3$H�;�N}鲣��z����������ӟ�^w���'��偔qe&Ź��
4Y����K�/��M�RdR�KYBԒ�h�$�p��$�|>l����k!�_=S�ޙ����6'č���0h|�2I�!Qh~�zr��2i�V؊��2�d2i�􄳕���ޤq�G�`T]��'1X7mI�'b�OX� 5)D�`y���A�����#|O�b�tjrD��r�����5I��{6�<�D� ߴ��D�#1�o�ȟx�I� ��p�"ܤ8�B�c��.���	�<{Њ��l�I�|*@�1�8R�̟���:#�iȁCV�݁l9#6���p�@�	���X�ݪ"T�z��1��vN_�HLA�E�ӦE��8b#'��џ,)!�O��!?����mb�xG�[#�r�X^
�O���&LOj��3'����%��3)����&��|*��'�,��̟:t7�k��W.:)xi�����$��*�Ԡl�k���'��ĺ��$2%��oK!C�Ẳ�'+Rc/���3�J�>Dt�&FG*]�HfU�'�8`:B�^�U���lN�Ee�Q0�O�EZ�"劤��{!�z�,�榹�Xwա��O�")Q�LV|���TE�A�tE��O�ęA�'j�7�E�O��I/9�A* �,52x��'=�ў��'&R�']��*`��A�A��cN8أ�.Ȯ.��=1�/t�&K|�0�$��ͧT)z���$֢s/�@�pb\�p�VB�4�?)���?A���}���Γ�?���?��w�ʜ��D[�j�A�F� 4j਺�I�s�J����
 A�	�T]�O�����_≐sk� �C<3�L˗iӭ=��8Ɓ�;�����8x��:C%V�I
�$�O�(7Mڃ��-�6�b樚7:���,Ͳ�p7�uyҧ�'�?��'���|�l\�Q'� ��j�(�#FM+R~ў���I�U")�҈@&m0�Ś��6�X�d�O�1nZ��M{N>�'��*O��*[�IZ�����9?@]����W�V��w�O����O����#���?9���BZ?Ѧ�80�φX�z��D�י �Hu���'�O�5���٠&M�����+s�h�@l�:3�8�Òa=�t�d
�8��y:0��mDHH�{��݊0��0�(�,͛4���k�"�'PC��i�EGxbNԖ��QQ��մyh1�dӆ�y2j�Y�lɊQkΣ��c2Gˆ��y5�րm��˓^bG�iB�'�੡%�Ӑk_����ɲj�t8s�'2��1���'g�)�]�r��] e����cö阑����a�ax�K�7�O���ǎ��/��|XgZ�!/��z��'�||9�|��'���a�ȯ�(�ꖰ~�"T�':D��@�N�\|(�2F+#����§��9A�${p�+]�D�{@�ړ��!��=T�i�r�'"��]��l����|X�L	 	̤g��
4���ߟԘ����G*p ���Y�#��x2$Pa[w����?M ㉀�q ���%jT���1��>?�a�jU~5R%I�&2
|Q�����uw��x�~{s�����L��3&<�9ai��F��x���d�s��O|�$$�'�?I�a�D��p�@�Q����y«ʕJ*d)�P�O1f	Q{&)�.�hOX�DMu�'�4xH��ȹIL@C�Δ! d�Cfnc�"�d�OV�D֘V�6�C �O<�D�OD��޽BV��7$�J)�,n՘E�"S2t�0ra[2��<��kU�J �˧���6��°p-���ǭY�O8Tp��a��b������1A���łz~d2���-@_B�'<u��$ި�y�	�	}��b��*�F<rr�K���%�<��ПH��x�L>��Ί�r9x�r�bȭ�bX[�k���hO�����'���`v霈K�ʉ�d��I���'h�7MC���$����?��'n�dcF]���P��*,%q~I�ɓf��2a�'��'��g}��������&fDi�uB��}V��P���`Z2(�ĤP#_It$�dG�"ml�	��N���O؁��� r�x3k�p!�tk�%&G�R�O]=��'��+jYp���_�5�2I0	̳ɸ'��$��P18M^h�DC�����3���?��il4"=���$�g�Kªр)"�P���~�2O\��dT�i�`�Ӄe�F\�#�|�qӌ�lSyR�I� ��?Q��C)p��u�P�\��qb���?���fA$İ���?9��p�L��L�~�!��G��$K�Iɴtx s)k�B�͟"q�Z"?�!%]��TYRb۹V��懔!0�p��Q����)��3UN��зin��k�$�*��'o����{��j|���dJ68z���\�B�`�!����?���?)�'�ā�(�=f�I@2[�m�J��<Iڴ�O���M33 �\U�,X��W�r� t�#��]���M*����O��'5��`�W����4Nm�p��ʨS���?�BA�q��1�.��7ϴ0�D�i�SB��ͣ?8,��gK��k�[��!i��ɕd>L�Č��k�&}X��I>f�l����hI8�l&P��� V���:�~�L�V	����M���i���k9��uA��}ф�pcѐ��O���?����gܓj�X��Z�_|E��<��1D{��'?h7���='���d�0c�Q��nA�'�F�� �j8h�IƟT�ɷ!��	g%���Iݟ<�	��u,�=z�`���O�2k�r$Hc�˄|��\3�H[�!���� ��`����)�Y�	�{b8��a���99����=q����#� %��a�ФSie\ab��6��ēC�P�(B8�( r�냮LҞ��	k~��ׇ�?���hO���w�=�LS`� K�q2��0D������]��q� G��{_�$sϢ<�0�i>��Ky"㙤4r�(׌��#�^��U�J�J��ht��'���'l��������t �GF��/���0hX��B�\<�8{��������*��<�ǁ�O-ε����>n�@Dl�!Hn��%$P�q��� �ː��<�$�b��!��%�j��p·�2Ֆ'��ON���O �O6��H!B���z���T���5=�H�d�O\�A��O����OND�f�E�I>�Դv�f@ W�Ęw�@���˂���O hmƟ��'�
��a�~��UV�hC˾��z���	v�����?ك�"�?���D��#	7���K�;w�	�§�6���ڔ>����P��	u7h�@Ó<�NP��a�q��|ڂm@E��x�"� ��8��N�&XJ���& W�� �'�����A�Y�q�8y+�o]�~b	c�(��=�O�x�T%��D{�ܓ�N��(L�R��'�V��I�/J }âD̍Q�.���cݽ|#�Q�d�b
M��M���?�*��mQE��O�0R�	w��P���63B25f
�O���ߔ\�B ��
p���3��B��!�`��,0�\��AZ�+E ]蕑`I�ޜy�'^d b���wy�!ZSm_0a.�q��fF�{��R�j�3M~}JD啒_a�m����┨�Or�o��H��&$F3 	Z�S��x
cV/RI B�I,d 9��F�C&`Xx�^�E�=a��?q�� �%ߐT@��zᤎ�vq�98��׆�M����d\����O��D�O������H��D�q�@�IL���F�q�fd�#)+�� ��%��N/
b>�����yA���&�%إ��KN�h�B�"'�,�X��P�M��#�&�4%�o�o4�'
5Z��g�M����*�4~M0q��5��}i��U,�MSP������O��)8&�H���٢x���s�0%�Ĺa��m�<�@�J��lm� �gȌ_�����͟0���4�����<9AŖTX��O�GW��ڀ�
���Ђ��?����?���_Y��Oh��k>�+g`�3}�Ɛ��Ʀ7�Ʃ�E�S�d�ܘ�W���pi���l�3h��p%L�3J�Q� �w&ܠtR&��.P�҉�`Q#�di"�"Od�bF,�mĭ	!` �~�SG�u���r�e��7�%�7�_ Xd����O썇���99���� ��*4�@QC	�3h���D"�"a�V�����v�8 	D�D�u��O��nI�W:����4�?��
��
��5�H��V�;�bm����?��L�8�?�����d�Y�J�g_��bɸ��'>Q'`ҵf=�-�V.5&�$9Ó"�v��!�D�[Ht�l�Dwr�����%e$;Hf銖C	t�����-)��#5��ĢE�|�3uN�>�´%MY<�!�_�j���Z��Q�H�ڗ%P=?��O��=ͧ��Լ�ԬR�j֨*�8"����7E�٢�i�b�'���>k�] |���h��ɃS|h�#�[���	џ|��C�J򤀖�E�`��1��:=|�Yr�Q�T"]f�CQlÉR11U�_���	$a��aH˦(V�iiG-��E(X�I����jpꨟ���o�$-��oy)H�!��� zv��OB�&�"|���:Q�L[&��[����R	�U�<��o�i
P��'���c8X���R�'�Z�}J�g���bd�Y3�n515L�lҟp�������.��%�	�������λ*�aB�h؁v����6U�����R;2��=AD�\%3�0`�Lg�'T�'�xN�6�Ν{���n�a	`��J�l�!��"3� ��aX'����$Y>q��47���{�? Jԁ��7z��86O�!S̴8��&���!Ub��[�j"�	�{P`L���<_!�D�KW����?BYj\�,HkR�'~v#=�'��rv����X����C�՞�2����ÛJDVb��?!��?I��N�D�OH��9�X����(O���MG
&Ǆ�y���%MMT��A�3y���1k�F�'��h�^�+�Ԙ�dX��萓A]??�cA�E~=ZU ���	uԥ��%S'"M�b�d��I�^��L(���� Ә�IAN]�~{���@�����l�	�*#/��xȤ�`M.D�|�'A]l� X&ș,;WҬ��>�$FӦ�%���#�����O�a�b��K�2��B��H莔I���O���YY-����O��ӄ|�HY�֠�X�D$(�jT����r���z��Ҥ֎1�H%�7�&O$hZ%�Ћ6ںI�ĥiz��0�!����Q�*Q8��J�)�(.ax�캟���B~��oL�b4DLh�H�����0>� �@J��Iτ��cS	�u���h�w*���Á�2z��T;e�HFq���Iybn�5r�'L�X>��!����qN�I�������:ɁE�`��2g�؉��q��{�h�z�|x�b֟��|Jfɡ�Jidt��*P�u��'�8� �Y(��
�Ʉ6�R���K��	8@��ȟ����W�TN��-��MO�\����%F�O���9ڧ�y��T�ɮe�!��1rh�B2⟴�y2�40rY��d�v<�l��nŉ��O>�G�DH�#x�����W����O����'t��'@0��XLR�'�"�'���ΫK4 ��cP����h@�Ci6'�,+��݀x�b>c�42&�U{i��;p�S8B"\�Srk[�Q��5��`΢7RzU���%����~2�Ή2r&���;;�f}�B��)p��i!$X:��)K>Qa$�֟��|�<�F�żp�i!��$7�d�83(�z�<��� 
{l`�tQ�`#��q��wyr�-��|�N>!6��+M=����^�pl�[��Z��`2#��?���?)�����?Q�O�t�'j�J��p�9W����G�Kf�jp��h	s�X<�h�Kpf���I'-�&��T�V<*�*"�*���n�}�`a��C��b5s�7�
�W	�t�'��W	_�cu4��`&�oI�LzCH��e���OP�=Y���c�ZP�+C?.7��z�y\!�d�'7pD���S�FZy(w��QN�'��6��O�ʓ	^y�%U?��	�4
���`D�	D� �j�ħ[��	��(����<�I�|
�E�z$[��li�-r�@P&T�$L�7��N��P�pl��{�8�K¹O��<y6�Ώy����s�֜Lm����_� ��E#ͫ�-�yVŕ�^���c�4*նx5�D����'���>zv�$ ���FD��ٶ�-r�O���d<	�f���	\�&�3�ݩ<�����Or����<!xI�T�^�b��+��'H剗B,�U��4�?�����	5E(��$0D^�:s뒟u�4E#5�_>v����O� �k�/eC }R �	d8K`�|�ϟ�Q����$c�)Y����G���0���]�]:�+V%\�8����S�1\��AqǷC�jЃtB�`9v�l����OZ�}�'�\��"�.<s�x�0�к2Tn���'�ձ� I�IDn�P�^�$1�q���$�}�OR��I�B�1 �Q�����5���B��?9��?���%7������?����?Q�w����I֌\QT�a��G &�qs��Ř(��͸fCU�B�xԋ�����OϤ�+�?I�/M=y�~�qdHۂ{�$p��
��HP���t�z��6�LI*<��I~:ݴ���Y�w��)��bE(nO����T�4������ !��'PўX�DE:5���
�;p)�TKJI�<�%l�Gw� ��˔5u�� ���*?���i>]�IDyBήdU1���ɐB��	�M�I��Q��ɴ?���'���'Tם��I�|����+۾(� ��&=?���)�.W"Y�-B	; ������"�*L�䑈+���<��mB�K�PX� �
a�p�4�R(nf�a��Þ,*�,@�{��[�4J����D@8~�
�M��;ۢ7F��H�DP��O���I�oS��@�V<��P�炵_�C��a�䥫�)îEON����A���O�<l�C��=Lx� yH~�جTDx8ya
��y��Ě��^��?�-O��D�O���):�$��Ѣ-�.���lAޟ�@��
�{���Ga3#���p")O0a
�I�%�lYh�''� s1D�h��}�3o�
l���ó��? V��5.Ul�'�d����?��O�@�����.�b�:�$��di����|��'��G��>:������4�<*��i>���[�P��޿B�  ��Rd���	Sy�AC�t]�)J(�P���bxr��E�/���B��X�$�O�P�Q������*�Tnu�)§P�8�Z�KP'���#-Z*��'F���폩q<�t�Y�a|��W�Q���X��P�],H)&`1a3��%�W��P8�b�Ol��4�'�y
� �d����~{���Q�j��Xq"O�=���ҍ{}�x#��R5��XЇ�	��A��DW�K�ʅsG��Mf��楓.����DN�W����O��D�O�ʓr?�]��7#� ���Ki�ĺ�eۇ��B�'�~!�g`A$ܘϘ'08E��)G�g�$k%��G��b�$��QH5�]�I�ΘOVb�����>��*�m�<�2�6@5d4�d��8�'�l�h��?�����P����E��b�A��хbw�B��'5!�(s5���)V�B�m��/\��D�O�DGzʟ˓����É�\L  5�X�Wp����?)���?y����N*dFި��)i2��A��r� ��ƨI��\����O3sȕ��I5*Ɏ�Xpo�--&H�Sd��Ck�$�!ieӮ�򷧌�X4Kw(CuY�	�R�	3�%��j܉Y�����{�B�O���9ړ�OV3'��+#�Y
Ҋ]��!���'�1OZ�Z,Y�O�>ɁP�֢R� �Ɯ|�h�>�.OP3�C�R�Ӡ_ `�S�L98^���ak\�|/��$�<���?���X��z�ȃ�Y.�;���l���.Ji�裐�f� 9F`��0<���Q{	\�*���2
t�Y<:�����/S�1ж����I:� �@�A���������O��d*?a��Q5v�D�%@B��,qs
@|�Q�$qG�.; ��iŲ9�l0S��<��O������O���Qm�q\,41�oE:��g�'���	_BH�����|2�j�"퓀M�j�����*3L�3��?i���q&1�Qŀ�Q��I���������"�t�EdڍS;<ԫ"����D��,�����Z,f�
Y�QH�J|r�#E����N�d�pw�]~bg�#�?���h���I2Z"N���� y2����Ù?~�B�I �@��B%�|�".�.���=9��o���0hU>8G�d	r���BR�X����JyT� h'f�Ο��	П��IFy�o%-�b�`��Ɲ<�p�J���8yY:В@ʗ2����.��4�f��dΫw8��ʡ���8��i�C�]�*<:�%P1(�����?���iЊ|���'QB���+
M:�E
�I�2Z
�EX���S>�Uߴ�?����ߋl�bq�:�̸�a����C�:_���f돕)�ģbM�l�����O �Fzʟ�˓*^�]ꡂۍIjn2Űaz(��쉅O7���Q�il� �r�\@ϸe�i�6_
�Ė>U����m��l�&��+<!��&�x���Ot�Z��Ob�$�Ol�ielJ�ԙ ��J�-O8y�XVӜ�񠆋�<S�� U
փ8Q�|� �F�sZ!�Kҽ:{24�D͘�ePl ��	ƚ��%Ĉ�4� ���u%Q��AW��O���.�ӑz�DAsf
�t#��ad��9i8��0?�‛�K���aT0N̈�� "IIx�\/O6����),$qt��"���СS�#��џHQ���ş<�O{`� �O/�M�/!�J�h��ǯ->̅	J*2���,��D�P���k��Ư�5aҍ
�?1� Y�$�	Y��0�c�D)T)ʩB�?O� 1f��((��Ǆ��P��Y���H�i�$�������9΅��W�D�H!b�Ӗ�y�\�?������t��d���̋;���+ЮM���H*�;D�0e�L)t�-zS�	|�`�T-9�3�?����c���kͭ+;�i��$����ԸaeE,��@��֟,�Iɟ���\�䋀S\�P疝L=��X�JI�Z,l�ƅ�tD����Ӕ���O@4�`oJ|��ۆ4��p!��ÿ"FBt����q�|�`�8R��������[��?1�ㅓYQ��"�;`o��1��CH��J5�'d>�)��?���o�X��n�P�l�� � r���m(D�X��%!�V���
:)�(�A��OޥEz�O*�T�X�ǏTS$D	0��]Є��*ȥ)�*��5�CП�����Ɉ�u�'db>�x��X>� x槗�;�
�&��	~����W� �D���	̨_�DE~BI  >j��"BE�R�X���b�&��8���3F\���I�(�#�&����6��z�-�3�\��V��=-B6E��K�'-�@�Bd�21����My��Y�l"D� w��'$!�2� |�9���<is�i5ҙ����]���'��DA�(B�H�5��$'<����m�yb���["��'��M��oP0��D�,YRI�@�O$���"��F�Nd0⚹��h�t%M\�>�����Kѐ�1�$��;�6ع��	j��<�,�"`�w�N�q�� ��A�-��l9#b�OE�O�`9�'����[]� `5�,�� ��U:h��It��0�3*p��P�f�^d¼R�c6�d0��|�U�ȱ�[�W��R�(��u�P/�<I�eP�?���?�,�$��r�Oh�W�v���ɤ@�5��AUB��P���
{~L+PnSDcnii&.F�Y��O�1�L ���V�8@6(�b�@��T�X&7O�y(��9<��ěc��u:���dO�ź{#��=;���.�(��4m7�)�&�	y�ri	7OH�A�'Dғ���R�S�? �R��.���`qI؁@�r�"Op˔�V�~�4��A斚6dm���D�O��Gz�OX\��h��^X1��I�2\%"��'���'��Ap�W�$�r�'���'���'��1�h��`��݅PN�Җ�(p�����	4!��	b N|�����'�\�鈁K�BԂ�=��-� O�/�L��RG �p6d$���;��ӆ�M���o���;w�>Q��W����`G�N���'�VX���?Q��m�,b�A�5#�5��@�c���q+=4��x @
x������ BZ�p��Y��Xێ�4�����<A�MÍ�0��#�� :XQ`ώ�ܸ��λ�?	��?�e���OV�Di>
�a�>;�4��"�Ks�ƄȢ�M,G��h3t뒵;�T�P�-�O6P�/Ĭt�Q��3��_�䊈IS� eK��j�'�s��фN�$���0����s�{"���z�Q�t�gh�OP4J�N�3@�c��*{�0D����㦅i��D.�� �p5f[�J�\�2�,
	����'Y0�A��lԶ�2f�W{aP�'�N6��O��t3�d�i���'��8�0��g��<T��H1���\kR��z��'X�gQa��6&�4w�V�0a�jD��x�<�*0���P~܈�42M�����$�y�<8+�G��s8���O*{� Y�Dʐ���I��X�j}CJ�>�����O�$�O�����'_�?1H�Iܜ-`���#ϻ_5X2�)!D���S)��SprU�S��=8T�3� ��-��|�^��	�Ѱo��|ʓe�8Y*�<����?���?����?!������e0<�JEˆ&lsF��#-�џԈ��鎧k`p�DJ�{� �2.�U��O�e"S�x��^����Ol��h�υ�W��a��#����d�sӶ��1u���ɜ4�����Op���O��I�MH��jO:@!�i�N1�nMCt������ɫ1/�����<��anz�=pʟk샪N�:b`g�6��TJ��F�6�:���?C���y"�����O��I�O8�4b������8}����ل2���
֡�O`��)m������%I�?7����J�'�<2���Y��d�P��h�di���'�R}H��?�Ư�%*	������I�?a���~��d�7�L&b��؈�KA?n�K��|+Ș��ܟ��AK��t���`��$���K	R|q��`0��*|���aK4AP�sݴ�y��N��?��u���z��'T��Of����D00%\N���B�BU�E��V̤�I(zl����O�1���?�'�Y���O��&mC�$� ��]�TU�� %�z�8P�'&�{�R�'�,5�ɟ���O�I '�N��lBpk��U�n�TM���y�#���<iT
Q��M{"�iy���'��D_'k��鋶R ̨4��	
6Ж_�W{T7�N��Qm���ć�?�l�:��,O�$� �bc0�a"˕�sxހ�6����C䉅
>fI 4��J,�d��}�T���<���?������|��dAZ]�q�I�}�H�MÒ!���n����ӟ��I���	�O��D�O����5H�aӀ^���� ����!'�n��0�'���'�"�'b"�'R��Ͻ]l��$��)dqfe	G�7M)���O ��)��/}�*�n���,�b�ó�M������'��O1z@�a]�v�,1nKi�b�m�By�W��&���'��D^7u��T���ƧW�Z��1DL�xO��\y"�|�U�P�'���JÒ>��\�Ԡz�d0�T+#D���֧ϮL��S���&�Q"%D�����^6%<pTpCCU��x�A"D��2�3o-�pUD�  څ�?D�4@��ڀb�R�v�D�����5,?D����6$�(S�2@����f8��?���?����?y-�`gd�@f�>Z$�� SB��l��F�'�2�'e��'4R�''�'"�;h�y;���v�\)�"3�d7��O���O��$�O@���Od���O0��� Yd��!����.�l�',	��L�nZ����I̟0�Iϟ��������՟��I�:�Byx�.��I;�tH���i���4�?����?!��?���?����?���ϰ�B׏ 8��h��F
=��7�i��'���'���'2�' ��'���� "�<e�H�3�d�d�I�j�h��O���O��$�O���O��d�O��`���330�����U38�D�z���Ԧi������Iϟ����������	ܟ�y&, �`B�x�C�D�\�6$��*��M���?���?q��?����?)��?��T_W.`�1�P�d��YX��#T|���'���'e��'#�'jB�' b�
�G���8��ܶ>��y�C�+Y�(7��O~�d�Ob�d�O����O:���O>�䕿v^ �Э��D�hX9��4K��mZş����$�	������T��ȟ���4 �(�1�.R(E��]L�`0۴�?����?9���7��O\���O8���O2�u`�=5TS�D(@��18��Ӧ�ϓ�?���hO�2��[��T�q�(I
3F^�YaT �ڴzd��'��O�����x�ߴ�yW �NJt�0���T|��*B�y��ei���I~}2��DF�Q�VE�'�&�
���=�*��s�ڌo��4��e� 4 �C�<�������$<O:d��Kݒ���}�7
��9�џ0��4sj=�'��� lH���+v�`��4�8m"6�j��'N������OYl���M;�'���0����JH�o�\�)"�p�4���*vbU:� ��ԫE ,�x�@�0O��)LG=�"��*
��攫g��I�t���+T0���РKp$!����O�qn��Q7N����Јش�?�(O�i�����k��m�"@8F��!7w��y3I�OVnZ��M�K�P��%^b~��3<&��YG�F���L��k脰0b��tY���Gn��?����hO�8��F�)S|r�[�M�8c̢��o�<A$�i�5�Ol�����'�?)1h�(� L���B�HF4���k����M�R�i*�9�'y��R�nZۀ��$c��q�X[���'�.	Cr�
��\jǝ|b�'��M��hB��O�f��`
2.[�!�2�'���'���'[剺�MK�M��<��i�=��c'hE�T��D���?���i��'�bf�>Iw�i�z6���(���(�}�a��Ef��3�[/K� ��<OR�$ـ&(�$�O  ��˓������r�ϲ5�P�ꥍ�	k��ׁ�O��D�O����O����O�"|����t%Щ;V��>:d���ßd����d��4e{,A��?���i��'�fX:�.ǕPm�m!�Y�LUP���Ov�X��F%|� �)��4h��1O*���k�0��a�ΧJ���ulV$�0%H�-��-��d*��!�d�O����O6�d�OV�D�/0���;b��Yx0�:�� n*����O�˓2�vʗ��y��'���?�1҈^�NLq�'Њ\V���G�O��$d}��p�t	l�9�?���TDM5=N�*v�޿b$��pk�_ED���),�{-O�i]�Wް�w�8�Dݠp��xum�l�!�hH�Ir��d�Od���O$�d9�i�<�7�i�Z��g⏻	��5�רL�x�	 p�"�y��'R6M �4�"��'��7��&,�	��#V�:>�����Z?�b�lڲ�MS���s�hD�'�}��#_ؑI��?���JS 	V���kI&/s䉡�B�O6���O��$�Ob��O�$�<�'Hu�`aaFJl�@UkDA��4Q.��̓�?���Z)�|�D�ݦ�ϻLbai�/�NOp	{îO�$��4䛦��O�ꓤ"����Vh��<6��,Nz (�O�A�2����$r�[��Lax���j޳![��K>����?	��?�%�ZN�p:���3�����Bɺ�?���?�����ߦ�Ȱiy�����<�'�o�%����)�(QB�E�I��l3�O\nZ��M� �'$�S9x�b�Ȗc��g�6�O^�_g�d�O�(zt��Y���z���<�����m�����ybȘ�o�<�¦٨ ���D@�3�?���?���?���	k�@)W�Q+M���0-A_)���D�OZ�l=8y��I؟��ش�?�/O���~i�犆�*썢�~�����O��l"�M��i� x�?�yb�'Y�a�L�sa8�r�@�5��)���.5Y����F� �'X��'��'���':2�'�Fp�C��=N�۠��1 :��A�^�0��4�@��?A�����?Y���+����J�R�Q� �j��I�M+g�i��<�'^��Jgd-n9��;���O�zm"���SBv0"-OD��gL7�NYè;��OB��[1n@R��H�Pޜ��IV�7�H���O����OR���O>ʓ+����Y��~���h����E&+��(e�T�?���i-�'���>�$�ie�6�O�` �!��q��!h$i�)}�E9���,.�W=O���S�w�X̱&� #�˓����������X�`b��%�R"H��h�O��D�Oz���O����O�#|��6$�u1�X�?,a���wy�'�R6-͏o$�$�O�)l០�'8�B�K�y����e�n��Wf�O�����GbӼ��ؼ��3u0O��"|� ��lB�|�`��&���z`ТE�}�&H%`#�d�O*���O��d�O��dƿ�`iX�p��c�,���g ��"Z�81ٴh��Pϓ�?������JW)v��> AY�	�B� Q[���?�W�ߴ���r��%>	���$hFA�����	����n4
�J�I���"�\I� *vy�O�8�&%��X��'���JD�@�+qp:#�)W�S�'���'$��'^�Ok���M��`$g�<hh�CЋ	ޘ3�G�)xP��?�T�iɧ� �>�@�i�@Izqٖ������o$�LkC+}Ӥ�l0����#�|�l�	1|�Xp3=R�q�'�z��3� I'x���?�6$���'��'���'���'mB�'��ӊ{�|���O�h/���C��ll��wp��I�����\��)ٴ�y�@�z�X(f'�9h2�=ؓB�?B�F�sӸ��	L}��O����O��;�`��yB�@<s����K��0ъe� �A���(Kp��mX"K�'Jr�'J��'�L� B�Ӱ;�QbB)@���'���'j�P�<kݴz����?!�vP%{�((�܌�b&�'S�]�K>Y��N��3�M�iR����|�N!1'��î�*< �F�؟��I>�0�B��-M1�i�'-��E�8��66O�5@�H��m�H�գK�}������'�b�'h��'/�>�͓b�<�:CC\#+��h��X,h��1�ɥ�M�EE��<��%��V�|�O���4v�Qi�g	o�򬒑M$��̦uڴP����ت���K�'��KP%HoZ$�2,J�z�u+������7(�j�v)q�|"�'�b�'���'�"�'�"��q-�Q�CÐ7(��&��")��M@��=7����6.�OR��?���OF�4b�3�����B�$`�!���p}blӘ�nZ��?	N|*���*PaF�"�(U��OYpxA�AN1�̌*R�X;��$
rb2%�`[�I��I'� ��ПXbl��<�0-�6!�p4e�0fG����	����3�M�&�i��I�M�Z����܀ �3�%	/��s���2�  ���'��6m�O�˓�?1�T��"۴@I�f�zӎ�q��K7��� �Za�`�;��ԝo��]p�>O�7��q�
�CA*��	>��'���I���ªD�W^�a��wGHqa�dϝ�?����?���?���?���)��JH`��f?K����n] u ���� �4l�6�ϓ�?�B�i9�'H@yQ�҆]���H� <���@ �O,�d����g�n��X��@	5O��D(K56�h�o^0y"L8c	�,P�<e�`̞�o��ےG/���O��d�O�D�O��$ԈN֤	�_q˰���Ċ�y]@����?�*O��mZ>���֟��Ix����{Cf�`P��0{�&�r�)��?1��I)���MK��i��%�SOM��RÆ�&��j��>~^���"a.{X�LHǬ�<���%�Ȁ�S�	3��$G�ؙ6���l��R�Fxd���?���?�����'��D�ݦ-i��	%��hؑ��b�T���Λf�����Kܴ���|BS\��J�4*��t�E�82�E�,,��`Ң�i��6�A�*��`��8O���4 �p�d �;�d�L�b]ҡ-����.I�)ojIH��?����?����?���?�����	�2]��z$�� ��3Ċ)X��6�9V��D�O���5�i�O�ilZ�<�$I.N)�ݠ��5̀#����MÃ�i5��d�>A�����+�<�c`�<��l�3kf� ���&��Mj0K�4�?Qg�~w���-�$���?����?���_���ǩ�nGZpXw�8}�t���?I��?�*OԱnZ�"74��֟h�I���H�F"3�޽�7��4j�L�%���	��DB��%�4^��Y>��L���J N�|Z���Ģ<��*��(=!�����'h�� �/ܜ�y"��!���8�BҊ!R�L���?����?y��?a���c�t��d�y5t�0c��Vs�\�0D�O�An��j�ܟ��4���|�'i�,��$�`n���&��_R��)v�@aӠ�l���e	*?a7�Ç"90�k�p9�C.��є�ڂY��8L>����?1��?���?A���?1�ʕ'�DxZ�䞌s�ε�S�T���D�ߦ�(e�L��ԟ�&?	�I4-vR$�5
�7m98lsB��X��O>Mnڦ�M;R�'�>U�S��\��KCo�F�A׌��P��e��edy�"\�,3��C�eW�!��'2��'讄��"	<2ҦuR�5:LQ3�'��'b�'�bP�� �4_h�͓:�"����� )5�ϔu�L�����֐|��'�T�rz��*~��Q���$]�,b1�0╩6�4Q����g\"+��:h‍�4�D�F|&�%?I�^cU�� uJ'F�(��Ϗ~�u;g�'�R�'��'��'�>U��oe���b�o���k���?����?�Ǽi�>܃�'i�%l�ܓO�pk����H<(I�����/c�Q�'n�����'�n7P��	�'�V���d����	nm�8w���<ўYa����5��k̀R]j8���k��� ������ԟ����y+:@"���ܴ�v)�Z�n�����'���yB�'��?	�@�
=��I����b��dX	�O���W}� j� -nڗ�?��$Z�.Th�2� �{¦͸1-I�{2 Q��c�4rW��{,O������E1��>��]�8#��4�S�\�� A@�KĄ���On�d�O��d=�	�<�V�i���!@���@D+��Q�tX�a��O�y2�'��7�"�4��4�'�46-��U���
�Ŭ ��� 5�A#j��l�5�M���½m8@mΓ�?�+Ukئ՛£�(�����f�iC�BV�v8�"b�v���$�O"�D�Of�$�O2���O$��0�Di�	X�ȳ�I��ر��<�Ms$A��<���?�N~��tz�<O��s���
����P�÷5j��X7�v��$o;�?��O&�)���	��p|���1=Or����@�i�.���cɐW�j�g'�OtD��UF�Q0�+���O����O���0_�D��bWS�ŋ�%\8O�����O8�$�O��F�ƫE��yb�'o�*�:!�3b耺\�,%c��j�'���>	s�iƜ6m[��Om~�т���3�F$iƠ\�"��%Y*O��C|(
9Jg&�I�IP
!�Gi��H��#'����2�O ,��q�1��O��$�O����O��}J�'|ر0�P�]+�k��&����"K��hE��y��'R`6��O��|j��+�&q�s"�05���"7�Q&���ZC���{Ӿ�o�� Z���5�l����6yG����,G�[6�xcT��7mt(BG͒&��M�W�G]�	џT�	ݟ�Iퟴ��ʟt��5;̸���f���p��E��'rP6m�+��	ΟD%?��ɯ]�A�`�0[��Ar��_����O Ho�M���'��O��$�O�0��NK�^i�F��<Z@�-2@&ܬT��5s5Z��7$�E!�a���r��x�I2�$}*�P��zI��Ι�,cz����8�I���̟�'�H6��<��6�\D(sc^7< ���GO\�:�d�$Uצ��	Sy2�'6"�F�&�u�B�	2abE)�#B`><�T��6�΅��"ޔ"��O��*���{n]�c�<��'
uk�V�"��t(F\��Pi#oB�X�Z���O���Ov���O��D4�S�?�A烕I�B\�UG��I[���O6���O6�l&h���ڴ���b9Q!�
w��KE��Q�bQ�0�'�I��M3��i9����T��y"�O�i�(q朿-sʙ��������Ofn�I>���?��?1��?Y���1y2�1�ICYzP���X��?����ʦ-x�bx������OK�p��	ԋ�bpф�U }�	����?�W]��:�4)���O��h�	�3Bo��@e�7w�����"/Z<#&�è"t�t��I�?���n��5&����'A�r�Եzp�C�fP�SU#���(�	�������'?ݕ'�7-<� ���6�?>��\�UdZ�� ����y��'�6�>�4���'/X7m�:}���W�Fd���s�ˆ	+*=n���MS1�Ω�\Γ�?��&�"gz�<S�o�.��$��#Icc�y�@�F���$�O����OV���OP��O���)�3EIr>V��K�K����ë�?�MkW�D�<���?�N~B��78��<O�m�hL�u�r��u��0��yW�tӒl�?�?9�OJ�)����i��<<hs=OizAD�3F���Ņ_�<UD��O�8#R�ޥ3#\@�P�>���OP���Or�d��d��c	�;PvXJ ���� ���O���O�˓؛֭Z�y��'��:5|ђԯ׼ {V�uG��p�BS���	:���������44�r^>��^$B
��˄z@�J��O����051^��� �)$���Ҡ��ț'x)���):�w$=arV@:��?)��?���h�v�I�y���{҉T(>����S)�d/b�$��� �!~�@��+�M����4�Z�iJ�w�����+��qМu�R��p�����Y޴H�����K�����'Y��t<�(�flدùmI�	����ҫĝd'�`�|��'!�'R�'�r�'��FV�KNv�I��� �
�23��;�Mkԅ�<9��?iN~���hL0 k�lI�n�XB���B��zP�t��4t��Ɖ�O�f�����%b@M�9*L�u�V"	P�r}��͑5娈#@�<)�-�Ot�B�
����?���c�rQr�h�_�:��4��gN�a����?���?)���?�(Ov�mZ%&���I�]���	1`�0�Zu#�$V_��(���M����d�O���'�6-���	�ݴ<-Ne�%b�?& ��Շ���<�r�J��x �ϓ�?i�΋�m���Eb�?��$�����_9>�32�_���@F�,-�H����?����?����?q�����R�_�Cnl8b(CKR�]p&�'"�'�R6M�88���O��m�m�I^�,1��M�tB��1�H�?` �����ަE�ٴ�J���R�d̓�?)Ë��]��qYv�Ch]��-T��ձB(�e!j �O>����?���?���?1D�D�7��<�a�$K�H�2gE$�?q����D�Цa*�ca�����D�Ov41s��$	���9���`\Pk���?i�]��#شvk�V��O�����	=~L�8�FCY���,ޚ��ȢA�ƄLd�0Tb������#�O�`����5#� 4��mP�'L����+�O^���O��$�OL��F˓K���.ŕDc��À]��+!a�lT4y�'�ig� �O�I�]}��i�FqS����b�2H�D�-��Q2��{شgH�ٙ@��<y��iP�� /����,O�9	�$T8m�����P��Q�C�OF���O��$�O��O����O~�'8](�"U$E��r�$Y�i ڴj�j�Γ�?A���"(�h�����̻UFФ:@���%T��i Ш�d@�7-�ئ�b�������)󟞍��"�3��$���+�.�
,��E� �rc����&��Qv���ܒO����O����O��SPL��G�V�q�%E�4�r/�O����O��D�<�c�i�tM�'R�'Z�M:D�V�a�rpP�W�@�e�|b�'�b�
���di����l�D)���B��A5� ��[��?a�A^u��"�o�uI*O|��Ě9c�I��f�лѯFLH\s*�n@�zfb�O��D�O��D�Op�}��'2�Y�S�U�j�ԑ ��W�ܹ��)�V�\#�y��'D6-(�4���)H2A���4��8����i�8@��覕��4_F��)�>��	�'�b��'cSdh��4�n9�� �6Ymd�"䚃8d�R�|�'B�'$�'m��'�BĔ�zx�)���Zl
�Յ-~�I�MF ��<����?Q������O4�2�،cRRy(q���u���r}�Fo��Hn9�?YN|2�����i�Ed��x0���z�޸��ŗ2P����$Q�r �a�1(��j �O����O�J���".�t��# ,[��Ӧ��O���O<�d�O��$�<y�i���'�p���B�D���@�`޽6Þ͐P�'�6�\7͡<���9����M��iVr��Z�W��ݪ2���.��q�F �n���D�ۭ�y��'n�Ԭ׭k��I��U�H�S��5&��T�@iq��}�>�R�Q[!��'�2�'�'��������0(��*���y����O*�d��8�Ns�����M����^'W5��k ��t�A%%��q��N}�*g��o��?���(AT�	�\�dF�!�̸��E��B��V��+GW9KAƃM��D%�0�	ʟ@���8�I�� �ԀQ;��YO�]�EZG��ş��IRyj{�^T��8O����O�:���EHT�kk4D���"��I��HجO8�mډ�M7�'��O���J �%�� [����:��Lǥ�@��鍽^#��ˠ_���S�d����$Cd��.�,�4�3�Z-@%��������џ\��۟|��u�SIyr�m��K�;�v�z�A�.�\i���^�9:�D�O�no�i>Uh�OjDnLT<���1g!h-��,QU� �ߴf��a�p��Ź�O��J��G�Y�d�� ;b�䒨X�%��+�ɔ(�������ӟ��ڟ`�I��\�	ȟH�O�|ZP�)ẁ�"gl�5 爰�2�i3ni�'���'y�O��mu���I_���8wᚳG��)�D��s�>lZ��M���'����?��S�?akQbII���I�=�d8�ŋ15�������*Yb�l�I��� 0��	L '����� ��Ƽ�"d�$2���3��
1$rH�5&�џL�	�\�Ra��Xky"�j�X�\���O�-��CCc�6)i7,D�[y�`� 3��O*e�'��6m�˦� �S���]�e��P�woӼUd������?q��x�����,�V>�<�/O��I��0Z� ��r����ꉀl�2p��Ɉ=GP5��O����O����O6�}:��� ����X�6��胼90�)��'��7-��8��D�OnZg�i>E�S�X�Hb��ʆ'�$1:M��$�4�	�Mӷ�i��7��+2���9O��D���@�@4c�-�T��1C��$:<I06��r��h� N3���O��d�O ���OH�$�OB�D�-��猑[-6�����6	��+v�6)D<�y��'}R���w�<��S��9��p��L�]G��H��>�e�iIX6͋���$>����?���$!�T��-�T��	�^ 9s �ߗ&q'�������>C_���C�|��'YRi
/%��<Q I�81���:�bD=9l�'���'9"�'��	��?�n��
�E�"U�)�[�vu=P0��ǟ�J�4���?	QT�TKܴgn�� �O4�&��30���W���H��`���ZA*<Ú'�r��I��EE-�0����?�\c�Z��f�L����܎k騱���'k2�'���'B��'�>��a�J04�^eZ�V�D4�hA�)�O��d�O&%n��-o>�Iџ��޴��*��` @��y��(�E���	���'�	�MSһic��+�`w(��'n"!�"԰�:�:c��I��O@�o@Q�A�O���2V�|��'�B�'���'?���5�L%1�P���*�cfS���?a.Ol��Ju������K��σs8�\[`�yT@���ȇ�?��ZM�	��Mkֺi�r��)�i柸Qp�K]���tdܔa|it�#�t���A�?��
"��u�>�/O��I-�$�Td�=h�x�`���r���O����Ot��n>�H�;���"|��g����KԮ]��-�Jfdr�{�'�b }�p�O�Yz}Bn��	��mA$CP��̛/fNA�v��⦽P۴K��*����<1�jx�+Y,l��.O$48��ۜe�v�v�X"DEx��f��O����O��d�O��D�O��$�O���`>��:"�x�#w����A�v�i�,p���4���'��®�y��'66}���b�#^f�EI^k4#�ƍʦ�0�4UdrV�����?9��xh*)F�j���QO�e������P>�1g��ƟDjP���~PpH+ �SF�џP�	ƟX��5� �A���P�,A���] ~��	ɟ��4.y��P�T��4S�TI����?��TB�C�*I�@�(V���M>���~W�	��M��i�����|�0� !$9V��鈯!ȎX��m�� �	!\�4��AiC���H�'��Dm��1�vt[�:O���Ź_늼1�K"L"�8��'��'���'��>�ϓ>7}���ҲN��Z��h���	��MS����<���91���'��i>����W 8�R'���HpJ�8�(q�I��M�3�i� 6m�2Q�N�A:Ov���sw0�p�N[*8�
�!�.?�|A�E���[�r(�g�7���O~���ON���OT���O��$$^�&Z�D�\��B nD�~B�˓u8�����y2�'����$�'Y~E� �_�UɓDZ%c�L�qa˷>���i	67�^ɟ�&>)��?��Q.�n���2d�ܡc�B\�Xd���AwyB���_��9 e G����'��' Rj�"�I@UꐙN�h���Ɖd��	��������IJy2�pӂ=)r<OX �2�ӂ!݆�)��	!8�t����O�$H�?�'吼b�O�Q��~�oi�14�V+k� ��f� yXȁ��@_3[�Fɠfg��lZ9V�ů�3*Р �O�A��=�5F�ύWU�P��\����۵(\�F�B�'���'���'�'��S dP�lb�5�5�Q�D� �9o ���O>�l�i�
�I��`ܴ��@��ɓE
ߴ~��Y��E<7D�w�'��Ɋ�M��i�����g���'|B�ЦWB�\�P!��"�r0y�}�X�S���'�2�'���'5��'_�	�S��@^P}"G�&4t���'�bQ�Y۴]����?Q���� K�0�#�雫2_ڸb���\��' &���)m�xe��d�'l$^i�T���3B�$g�� *��<#���$�7��$��%)D%|܄�Oĝ���f%����$�ige�O����O����O���$�>�Fa�����ЩY� 2!,�
eL�K�'�RsӤ�O��@f}� v������x�%�ːOh���' Ҧix�4G? 5���<)��b%��@E,E���-OH���q�R!���x����O���O���O�$�Ot�$�OT�'G���� K@�vR�Hi���9���ݴ~�̓�?����'�?�Ѱi�d�??@�8���蒉J ��|"�7 ���r����D�
�)�T82�̀s��u����BĽ�7jP.7���d�~�B0p�F\:S���O@���O��D�O�Q�_��%���?�~���a�Ol���Oj��<9T�i.�es�'�r�'��,���2+߂x#ՋQ�H�rAフ|��'p�}V��	a�j=n����� G��q��H'��s�h�(A�r�'h�䘐%�1n�>��]�P�ӪE�H��0J�<Q�d��FfNи`��N��PB�����ş��Iɟ\F�$8O��P���,��٪*]	j��!�'�����y��'�R7�<�4����\�*C��zh�,��U����v���P���4c��֠�{׎Tٛ'�R��i���e�!�L8���Y�7BT�H��_�𳖍3�D�O����O����O\�D�O��dF�F�i7�M6J_���S�;���/��g��<����?�K~*�^�B) �߂/�$ř �i:E�_�|�ݴie���O��Z�����q��aȭV���nV�U�W��1W��B�ò<	cD�2c~� W�����?�~�䨃 �6ʂ8��IqԐ����?9���?A���?*O�0�I���3�0���yw�D��hH&���d��5&�H�	���֦�ڴe�b偅\=�hض��:^�����GH����<��5���Zb���_;~h-O��i�?fr	jVL	$ba(��G���4^�H�!��^�~�[աLdx�� �-�2D�"]����iZ-Նp��'�!��
S�9&J�O^��@B 8�!�u�w�ܡZ��7^=\���O���ЧI�[v� C�BG,`"AQ�
���a�"n̎�>17L�n=Tt	1�3=Ξ\��h.n�LpJ���b���K�~�"fI��|d���)�$`���#�.*��{�m3��؇ȓ � �;�"��;�����gE-p���	>)l����O�L���M	.�(H�Ɍ=�p1A��B�G݀D@s��N��Xqҋb�r�۔�J:�x�Htˉ��Q�u�I�s�PhrD�W	AEf���E�7X=���P��-Qh E��@�Qb|�#��'90��ŇPUm6t�e'ɡtgX��ę�a
�a؂��`���A�ǈ%L �<�4K�O���L�#u|U&���I���&�ܱf�\ S2�0�I�u]�%�Wȋ��@�IF�J��	�4�Iǟ��I՟4�	���CJ�܅Q��ã3$�i	� �3(.&$�L<����?�N>���?�S���o�h��f�*1�@�� k�d�J|����?����?Q��?���?����$l��s�|�۶d���L�с�?���O��D%�$�O��D.�����>����KC�^)iDb�zâ���ON���O���O���[|�$%>���N�����.+5�Ԋ�
����Ix����	/Pr��I���	� S8l��R�v��B��/z\nڇmu�d���S�VTZ�鄅@�C�<x&̀���5D�:��h�:(��"T��X�1�I M��j��?1I>����?�����
�"]���YNP
���C�M�h�
,O����OR�$1���O0�$�OdE۠��7{E��I���,|	��do�8o�?y��?��'��'�?��b��#��ԉly��`a����lBe`J�X���	şZ� �t�3��O�ԡ6���K����"�`��C�2���BM�4_+292d��b�� �oμ,�.u��*#�h��	
�?�ΜkBoW�Nx��a��v�ȠYBl�&-Ӥر�c�� OBp[�섨{y��s�ʅN)�1�	�#�f�W&�<�tx�!f����SoQ�3p� WY�5qvi�`��m+CY�c�B���W�E��kU�i��ӧޓ?�b�'���'� ���9�@���`��e�I�,�=6g<��zu�'�Z�J�)��Zf��O�xhd	Q�ЬC���>2��Г�MG}�$(��u7r,Z ��k����'4`���̆j�fX��a��m��E�G�����I*{88���)����$�O:7-Q�,آ���-Q�dA��(F��@!��O>^0a��׿!ì���oԐV=�d�|�'U�����$Ϋ&3���u�	�H�F���J�"O�tT��D�O��$�O���?y��?���Tv��3s˝�c��(�F���q����
%#�4����8\�y�oǾ�t�Pd���gW2}��� w<(�p��v�R�Qu.,��yB�͖�M[��+�<q����������K�YҬ3���OL�D&��z���P��%����R4졉��'��O,�`�K3?�D��ˀ�B%�5ڄ�>�w�i�7�<I���2sV��'��i�jii�G��p\��@І��O"����O��d�Oja��`�^|$��݇A��Yar���]��׀9g��#?A7(G�Y,����t�R�6b\Qb�C#�X�I6�:��O�3�'��6�Hۦ��	��ʬ��KѬ�
�R+p`TT?������h������!rUY� �".���a��'�&�IZ*N����aNd���+��$�)O�%
s��O��D�O�'^�v�����M{��ăGrq��X�EDX�gfX�W�Ba_�$UR��P@�~^�1Fh�*�'��'����&���U���.�8�'0��ɥI� ;�P���b�њ��S(S&u�� +Z���BI��������	��M3p�i�R�̲e�$������Ҥ�ОyO|�'B�i�	�$�Ji1�)�)'�v��g�0uʤ���؊�4A����|������펳��3E����fM�����@����_��)��П�	��|�f=�h��H�4|�0 �bf��[�HF{y� ��:{��dk�r��d�&7�֕2��ǱV�tj5�Z܆��P/�5cA���móX`@떛�􎔞^��C�b�6a��%�a�����30�rӮ���>D?B���;��gy��'�f���R� %���9:�\��C�ˊHF���<1��?�|&��꣨�Q�D r�K�\Xa)��pI�4��v�|�H�\J)O�|K1��[�H7KY&1��@c@NQ	DҴ���H�O����O4����3���?a�Oi������`\rt�
��W0NEc5�D�}������
q�.ԅ�I2�!��F��Q+E��+]�&թ�N�d�� ���%e#�z2Y��M�A�%>�0\:�O�<BB�AV�0N�7�Ʀ��	Ry��'
�O���V�b�֍jQmC�iG�a���L�y#�(��D�C�Y}t*�C����I>{����<	Vٓ|����O|��f�<�񇎇�@?�Y8`)��9~�u����ڟH���Ɵ��Iߟ�iũ=yp�9������o���xŉ�D�|I4�ω{fP�g�	?t�l!S"gћ`���	�(���1��%�r/V�2�y1�GR��E~�A�?��i�B�'��S#���"(Ӌy^�} u[|K0����<�	ğ$�)}�j��i���J�)ʟ$0���K+�p?9%�On=��� =�T� �,�/bh�Y�$�fyR��}��7��O���|�`��<�?)ش=*P�H���t��;�B}�S�'��ȒI/�r���Z�-5��Cϩ~BM|� �B0	@($^8<GA�I&�b�W�<�g*MIs��.	���	GI�O�h��s%^$Q��5��	L�l��$ìO,��&�'�X�O�>m���ܶ+(r j@#�Iݜb�/D��!$��$4St�9��I�!�9ʓ�?Y��韀�s2��14�:�"�n�'
������$���(���QCO����� ����ę2�@C�@�nx� ��X�/��0�҄D�"{@h��� �2J��K��?�O����cCyr�T�ꕩ�H��PP��䑯j���c&K��$-�C�	WMҵ;gJ�|�T�KgO��H�irީ���A��H�c*��Y3<#��
�?��4���z�'����'7��'���'P��R$X\�@���[BX��4�V"�y�M˘.�zEh2��=�F�i�C0٤�D�{�'�N6��Oj˓)b�0��^r����ǅ��90�q�g��<)�'m�O�O��ɭ0�k�C�,IWf,ٔB_z��0>Q��XD����<,��* *^�8B�I�m�����6�l��
 |�B�ɈR�l���q�0\��"��%��C�I�U�Ե�t�)���#��@�k��u�ȓ!�D�A0��v@P��A�]Z�����r]	��3fCܜstkwJ
X��^�"��h��m���`Ɖ������*�NEi�@x�`�D����І�-F�������ȘuHފs%�ф�hvA���#�.��+R
Kn�ȓ�EQ ��\�=���AJfU�ȓ�z�R�̚~�>p(#+U���p��a�bD $��� �̗��(ĆȓO��3�͌����C+S�p�U�ȓ2v�1u䗯C�
	5�OLJb���*��c7o^������ă
����6	�,�s�3Q��`�MĂ/�A��(-�!�rG@�tm,D����";sfȆ�P��qx֏�J��d(�,'Т��ȓ�6�����
�
d��m�:|�ȓ�$<���k���MX;K����@1N40�H֟8�T����a?L���E�IpŬKm�R|Ӵ-�Fw�D�ȓ!�����~K$(+OҔ�ZQ��_��4�偗�<��j��G�h*,�ȓ<(t�P�D�F�hl�áx٪%�ȓkHD�H7�H>� +���,���ȓ)]�eȖ�Z�5�iy� U	I��8�ȓ�Tp�D�m��*VC��WJ �ȓ�R����d��qB�վ?����ȓ^�TQB��V%D�w�� t,���,J����i�d��c�����'*֠��-�K���h殔�I P�a�'cV-!p��ez���0De��'B�x-�';�@�B�B3��*�'�d�b�م�Pj���1F�����'L��`�E?9��:g&<Zj���'[ƅ����MLVU���_�@�zPC�'��s�,�x��mT�a�'h ����W�8�{3���P�����'����	�ke��C@2<��'<̡���2~L`���1-�q�'�,i:�
�=ʐ���A^ �0���'�BCsi��c�<x #ΙC����'��T[�g��j@�|k��'D��*�'�J��6W;����Q)�?M晑�'����D��TN�x�фɛZ�2d��'`�c��Ō{4��$�J�W��u��'^pѡ�
ϣl�i*tJ��V_�Ǔ�HO��Q�ֳX�Hd&�q;<�ڷ"O�4ia ��0`�����=_���>������GE��;���5!�F�ף�U�!�� �����U�T:R%�R'M!51��Cp��0lO.��:y��x0%cF
��|br
O�7�G�X�(Y���ܤ(�����L�!���XkxH%J���H�J�gOX!�x2鉈;�Ṭ�ײ7���*�vZ$B�ɑV �����gOr�zЎ^�7�B��Rɬl�3䍙X�D�g� �.l B�	�l.�+��=F���js�
>ZC�	'{��4"�*�J|��J��m�$C�		>ț���2�8�v��-G
C�	=U�X�ceM���CP/8�C�IP�%�ǀ��%�����ʳ/iB䉜'�]S�О%�@�a�ʩ,�B䉚?_�m��i�	^�`ȸ��*/*B�	����Qe��O�x�s�m�,�&B�	#�.yJ�&��-�H�ӯ-8�OL�'�/��<��D�#7�4x����3 ��-UB��d[� ����m*c͜�:�������!v�<��%LZ�3�!�DԄq�a�F^�5F�`U���H�ў���9FP����Q)�O=~����!x��saeK7Bnh�'Ai�^Q3� ��a_�I
����4 �ܫs��"0��)�qّ?7MO0UN�b��χc=�Ը�	~��"Od0��Ep!@�#�x�$5���ƣ�?�g��V:n�7��N��3�w��	�i��Dbh��e>��e��ɗH{����/ Jh���@�	���(1�_(E�=H���L�h���'��;�mԽH��a�d���u"���dR?��{-U�M��}�4Z�����I/8Iwg��b����^o�T�ȓ��=e�\�(}�\{%���OJ6 ���2S���b��R�8U��� �h���WQ� �!��Ǥ)�z�����0!�d&ElpAK�ѣ8tH �� YF�tr�״v?����H��)�0�r�=Ar �I�Q��q.�� �f��k�e�&�[�&��b
C��M��&?N0U����(�> � j>�O6ؠ�kG����+`�Φ1�,l�'��L��q��c֍;01���Og&]�OO�yz�,�&t'�%��oO�IBV���'� �:DD�T��m�0��@H�@$�P4D�Q��Q�𤎨DB�X$�s���jخlV4�h�.o.VC�.D�cDe�x�,B;`;2�1����3�F�Iv)�|�6�kf��V�j�_yr�|�HQ�ҽ�%��6�z(�D �0>��#�&��9��<�����8e)�d	�&T��Б� k��)OT	Gzʟ�	�'[_�@��5B�> ��e����&+ݴ �Z�R��U�ƿ��Ӛ�n	�ƋJ�F�� gV=���� �)��<��.���$�"F�6�P)�6��1[�Fm1���(j�!*#��op�G���)^"��Ҋ�v ��®Z��x]ϓ+�����$W<	ɤ �������-��hD*�L	�aA�(|�n�R`Q?�}��e�'I|�J��T�d���/v�\��
�_�v�be��V�nXRc��1�~��g����D�$75�hK� �#(�S�t`EG�I��^�}��	R��%�hObH�р:`���_��ħIR��ҵ#)j2z��Z�D��e�l����󄁼�PK�dPc�`�`�F�$�$�\3WE
F2��S�O��(T�J(P%��E��A�'Ѣ��(�«G<d��bE)����	B��>�ժ&\�KL~�*�&���E=EkL�R�I_��$�R�ܳ)X��M�	���FHB�=oRL���J PƼ8��I ��B��qExʟ���u�� <�QJ @ݺS���S��'�Mrp�]z�I9]jƐ3��1b�� pȍ'f����&,�S��yrcO�\�䢅+�\���ј'�Z��"��IL�Z������;FY[�eƧu4�+*�a~�?�&�����w�r��a�P��0>���M~��%�H0:@�Us2��a���yr�^.c�� ��ˌL���9��ƶ�O�����O"}��K(b���'���eB�Z�<�A��=���H%'��� �)���������S��yB�B�_K�tZ�������1B�=�y���dq(态?��q84IL�yRG��~���� y�4��z�ST���#a�Z��'���'����� U8��K�Q6J0�� �y T!d�EI�+Ģe��qzS,U(�O���O�#}B�A�K�\�q�]�9�6��q�<�qn��b��I+�h�6���ȧ��t���S��y2�� Z��x�!�}>�;Q/�=�y"F�>,�bJ�Ns>5	�f�/�y�&�O:9cG(^tb��E��Q�H�Q�'��'����5`>i� �e�*V�,�	�'�b!z�Ѵf���%��.[BM��'����բ�1,��d��K���#�'�<)�`�� 76bm��� 9����'���/��z�.��ac�2�du)�'U��� ��%fA.I���y���!�'MJ�Z��ƹ���� CŶw#�'�|�
��	�p~.Ѓof����'�,!�%�T0Rp�A��]�B ��'��\�G81�qx#,Y�JK����'Aܬ �`��\l*e�]�E*���'�>)��Y/Eb��w#@�8�L�8�'﨨���O1����&�5�N(!�'�~1B�Ϟ(�H�S��!#�r��
�'J�1ꐃ
D$�ʔL�`��'� #����
���C��.��D��'�E3VhA��p����"yc�'-8lQ�O�>fLBV�v���'� %X�/�+q�qrVK��mG���
�'n�d���	�E�a0���o/���'�d)21��hK��Sg�^�����'z���!�hP"��Ȕ|��2�'��$���ȳS�R��%��h��
�'::��+�[��q"g��}�D���'�J��,C/#�Puc��Gr���a�'�Љ��CI�#�Ãl$4���' ���N Aְ����[@@�'N�тo��॒2D��K�T��'	`���X�<�{�n�I��!�'E8%�`W� �HI��.	Y���	�'��8S�.�*4���)Fℭ<�D�	�'�(�!g�2.�lh�u�H$�� 	�'R.Pa"��	���]y	�'�\$x���#�,t4*�h!|x9�'�6�1���)oN����Q�:���'�`�p.� c�$���B��h��'�ʁ����
��1�2M� j�d��'��v�H�G�h���������'��iU��$s����Ȭ�	�'ghH���Ux%<X���V�S	�'s��3�b�6-�!��	�&qf�#�'BJ I�D.` :���G�nH����'�nD��f��_Fܣ�ǅ�p�0�'�h�����^�X�	�Γ7|� m�K<��=�S����Q��ظX="��7��1&����	>6	�C��0%��1����q�YZ%�%��'�]R�e8��Ґ)�u��`8��s�5�%D�|buŅ�B�tXW�^�Q�#�!D�����@�d1f%6/كnl��8D�H���%�:�#k)P�R��"6D�H�5O
�YZ@ԏy�"`0��5D��r�d�ANɶ+֯'�
�Yŋ3D�X3�k��P^�I��K2L����$D��s��ˏ_P8d��c]��V,㰍#D��5�%\��TR��\�T�7�<D��q���D�����G�)$��t�S�?D�� N���V#�f�k ��G�8�"O�}��H�N'������<C9���"OvLie�S�N �᳑�ӒI�~�C�"O"�Z`n�Ia(�T�����G"O.t�`�5��&���!���!"On��`.V@�`Hc�D �B8��"OD�kE��<�ֱ��Eχ~���6"O�l� Ȼ:�fE����(MjE+V"O��4 �4CT���=&(�9$"O� �`cH�d@�BN��Ɓ�f�7D��h�@P�m;(qZti_��-�`�&D�|[��Pt�D��@[�Lt��C)"D��B�fþ#������=��`c�=D�@jfN�%I�޵;�M��d������?D��6(W�^�cO�3:HEK�?D��B2�"�����ƣ(oP-��"/��1ψI"��bt!߸[1���9^!�d���@���oƏ�X�S�B#Pg!�D$�68a�D�7X����ր�<���dAIR0�a�M</�0�����y����c�m�%��M�g��yrj� ���q�AϷ$�x��Iҵ�yr�"�*srn%�ZT���b���8�,�:B�[�v�8��`fl6��ȓu�l���ڥl��f*�.�����$s4*�+ɃB���xG/�8LY�t��Y����!�_ 1��8��҉b����ȓL�d�9��L�5�zA�D��k*d(��D�*�IE���N�(�"疎$� ���A�j<ˁ�_�7H��S���06Ą�fwL�h��0>3���e���b���ȓ6�fqpg��PUd)�"�-D��ȓ]Ǹ�{5E�"]���[���'tby�ȓo4�hA&߯<��`��h� �ة�ȓ+"L�0,]�&<���H4W�
���\��4�J:J��D(G�P� 0.�ȓ9���\'i����r0l1(%�ȓx��[U��E����w�H.��Յ�p��-'nY�A�XP���-z&�ȓXt�옖��Bw�T9��N>0@�ȓ5�*�{�Т=�<Q�J_60�|Յȓ9��hU�	�7$���5a�5T���ȓ�L�H�������nY&"7"�ȓ9�X��T ˎP������܈l���ȓ^u�)I�MB�#_�T����~��ȓv��K@fڢؤl���Q[��ȓ%��fhUW�� ����~��i��Z/(�tK�.k^��	U�E�v��M�ȓB�0 0�V�H� (@�M?e.���sڮ�H�+�'<��,��6�ȓ3�j%��)F�\��#BL�~%p��W�Vj�Ƈ}�B)�e&˶M�ȓ8�\q�j��d�X	�& e ̈́ȓe�p��(,<������R�"u��c����K�R,��rU�)��Y��2�
�A�-PKv�Qš��b�"�"w�,Q��y©��"P"�̻0dE�C!"B�<�2L£m喩����[�,Q�\�H`hj�ʅ^ز,P�I��\𙡌��p�4�	b�R,��� N['nx�I0U���w'];�l����/�"=!s��j��չ����06B��c}B*H�)����e��d<���ư�M�2��sU���u)��'}<��Dp�'a\��QF�62�H�:�F��aT$�S�4��)�B�)�)�6��;�¹D~R�W�!�����#܁ ��S50�xF� �OT�yt쒹W�61� �J��5i�F��G.���	�N�5k�w���J� %X�0�.�T8�X���Z3�_�Ԁ ��c7�!\q�pD˒q�*h�SN�6c��P��?���Vܓcږ�D]��6"B����%KT(dYD�K����NT(vC���`��l�6��`	B�:30=� N��<�rE�i�(aP#h�����7h��.� �dɗV�h*� ���Tm��!�A��Ğ�b��9�UEŖ[��)�bٷ��V�	�z/n��bA�lD�L�("/�HQ���F �?q3�ҘfX�x��K��u�:��w�,�k��m�Ģ=ͧN`  ��9�Ь�R`�q�\@�c[IpXzr�''Э�VF~ �hcvl�P :$�tF�O�lc����O�#���b�
`��"�OF}�� \�U �z���h�z�r4�'ab� �ǣ}�D��+��#>�R�2X�bmr b��OxU�$ʸ�MCE��D�3V��
E3�\�'����ϛ�=�3�F�Y� ���'^��mڃ~�h���R9H���Ǜ�?7����Sn��� &·�ثǩ�">���2�YyX�l�S�C?���P�1�����o�F��f�
tǆ�a�(���7O@���u���?��iL��"P���d�7�xxPoϻ8���{�W5c�D����'��s��H/�|21�H{b����>�`�i��
yf� w�+�M�C���L���30ռ<�Q�2X2�{2���|<W�ۓ_��-Q�-��g���o���?�u�Oռՠ#�\뜽� 7�� ӌdӄ��c��W߂  놖[����E�	+�xYk��ė~�t��i�S.2��#�d1}��O�ӧ5F�B ;�D�T
L87�>h���Ɲ9�*�+>,O.|�"��{���ĖAXl�S�hx���"�Ao��'p��G�]s�D�?7���fɼ0�m �~����4�J,��=ѳ�X�Q 4Dx2�C}P9sa���X�y�o���M�b�
'���(��Lb#K�l�$�p� �����O� m�+F���p4,�&��!�q�I�O� 1&�����P�@P����2#"(�[�K-5�����!kL!2 ���e(0�S�L�<�;c"���ҿ#��y�	Dl��H��ib�7��%,��` ���az&�I�P� ���R�S�y��J�4ht
1D �)k�8�˘�O�햧u�ڟ�}y!T?ט�8Sn5����UD����ƬY&`I�7�F�p<�C�[3f���w&�1�bN�q'8��a�#s��� b&��u�[�;Pf<3E��i�O���	28�2��5��L�`ք4��X7ժ<��q�?Y��BN�~��JьI�|�f�5������	��q�s\�8������ ��'��P��ß��	0 yp�u %��9����C1��R���Z�P����X���,>��8�^�H���+l	�uyBF?�R����D�\��`W�?a��AWM߈4 &
��amE2�T7���/��f��2`mULTp҉�$�qĦ-�oK�ZH���SR!Ah�2\��p����8J�q$����d6����5F�wDR�q� պ?byaס���xΑ#k�]��=��+�l�']���*�(ˣ8���v�Fx��O��BI2<���n��i��?)��i�q��E	>%��Z`�۬kK�� q�ک���!T.2��q�D���J�W�A�Eꈕ3��8E�D8�,t�FE!&7:��bƂ.�dS��"��!����K�,��\E�qO�q{L|���:+��PsP��3�`����ژi����&�G<�tF:�.����
K2xQpV��i_����?���_�@�����.Ŗ��o3�M[�'L �PMX�j[�*���aB�o�'?�5#EF�.�I�F��~*���Ar$� ���Á$)�؊�J���4E���'��P�p��;*T���[�8`@Aj���OG���D�/,u��i��S��)t$�	��HՓ9$k�+.%�BEƐ�K��=��dH�f�2�y��ٰM�d��hZ�:PP�Z0O5��-��*�8�?�T�P6G4zt��"� j�;$dC k��erF�O7jۮ��&��[~<�$F�T�[��r���}�ɛ.P��w�� f�z��DX��:���vKx0 l]�z�F(��'�#��c��G CB�T�`�"
���9���-��3&`E�@�)��/q>u����8PD�4m�/b�d�aD�N78�܁��U$S�� bA<�uEr�Dj�zɊ�l���ޕ��,����	Υi�"ʣn�(��5� B֯���(�!�R�<���@b��x��c�Z*r�P�$D��U"r�>Y��Y�����ɏj�$<1Ҽ|Qr�i��-o�B�$f%֬1��J�t��JV��t�d�`Rj�:s�UJC�'0��h�J�$nb.pC5��(|�A	�.�.qA1��"L�|�4T�i b�
CNJ�z،I4F<�ȓ0��a�A�Fڢ4�˃�8�@<$�4�Ó�x1@=��&l�C'-���4X0�f۠f���Ē�t[4���3J�D��/W	-LTۦ��~E��8��'t�s���v�a�
W��T0�AH�"��26`OA��F�+�
Z.ȫdL��X�D��O2�h1i��8�ě%�8	��TJu�I�KF����Z�H��̐p
�$%�*�`%.t���  ݰ��}fV�R�R�A�(�K�9`�]�cn%O:4���"���2@��@X־iR�C`i9��J�K�AK�tj��d�pG��Ѯ� ii
КGQ�}�f��'��p�@��8���a�K>��,:��Hd���ė�n��Ձ��x���A�Ɲ_-��`�&�\�I�@�6�O����؍~�h���Bp0�PBe�(aZ��׮�U�8zڔ����M�tJ�}#�OEK��Ȋf�����fQ[��ɒ/	���BlU�@]�\ӄO"s
��S�? ��ق��5#��I�
���cۿm�]16gС^ԁ�tD!�A}����l:��q$h�IbHxC��u9��EW�v�0�Q,I�bi��&W��O��F֞IR�Ro�H!z����~��l���O&H�K��Au�'��)`v�<#f)2�T�|�QR��"&���d�q�@RC%X����r�W�_x�����(@Ҭ+��>���i�ݥON����,ݚ�P��޴7Ҽ��V
j�P�#�d�0q�?�N5n�{�K�TT�BC^?q��%FX����j����s>��'����O>�Pf��a_L�4�J�����L`}R�G2x���@�x�ul��e��t$��=�`pP晷�?Y�'M�����Yc��M����(�x�S93�.��w��Ħ;Ɖ^O�|(cN�%Sv���$h1�&�t8#����%�Hq{b�S�'������"<[B`�����<�LYL��M�%��6�	8����@�x2m����m` �w,� �,�:����P�f������)PJbѨ�b
:��O�8�����6��q{��֥L�M��,HGΌ}��EiȘ��e	Yb��|��G6�)���%/�� � �!3�)Dz"E�[l�������[�� ����� tr�՘u��7G?Jj�n�M�xB#�N�w�|q�OF�<�U*@�5�@m��p"Q�C��E	�,+�("�o�q U�S��E	�l��*&�ߣ��O���nI&oW����Vۘ3��'a�e�r��{?���?�f`�|�O� ��K����P���8*�G�5@5|�Ǔ\���S�xz�S
d��!��D�,^hp�+^�5^8�B�a?�N����&�hO��b���C��M^�����B��`l�\� �Y�����"��t<�>A� ��;��T����V�֩H��,����M�UJ�F�d�c��R$|����;U����Bֹ���]�=��J����Y�8h%l�+y�؄��/��$���$9�����蚱��M���*d�y�V=#������@�O.��E����cx�����P�G~��E:�H�0W���ɠ�N���F�	�2�&�)/?y�����]&=�:b��4�0��ҡݙ s�����eǤ�I�n��xbb_ ,���/��t���澕��)lm�L�4X�X2�,}2�Z��z�I�LOr� �MY�~��Y��iٓG8�a���W������R}h�V�Ò��' ������K�����T����1:���'��J>	ф�.�ħf�����?j�5;�B�1#V\xe�ډq[8�oZ�&�Z��0nԊ˸�~���Ms���?ypxAǦ�-z�  �H='�'p��@]�g�ɉ0���قaQ�$�XL�ł[XȝnZ}[0-H���X�g{��=�3�	�<ɖ�6I^z���h��
�.Q�0H�,i�`���'
*ɸ@!� ��.�� �4"�A�: �pǃ�}�9
��OԢ=QG� ��I9Z�Ib��R^Rɉ�Q�*(�i�?�Q�-r�З�\7X%���e�<�'���%ˡ
<D��6FG�i>�ؕ'*��#�8])���OQ>�J&A�����T ~���JU!��$�����!�N�Sَ���)p��v�1Zd�J�!ކVN������I�M-���\�3�ɿ09"	��S��9��I�,�|�	��O�@q�ɾ2a+��O�����4�FH�U)E��ơi/���C�`��R%��	��y��㼃�ǖ�o�╺pi�}�R�0ㄖ%�l��&N�KQ�<�O{�'��y�O��%t^����-��	�b
Ha��b�C��Hq���~�Ob��UF�j�e읲@�pظ�'p|��]�5<a�F�2:�=y��P��Y�� �)�| �7)ϳ�M;'�s�)&a�nm�C�xn=�`l;D�`�҇Xɾ�*��ش#�"���!9D�,��B :b�k��W<(R�Òo"D���v�^�ő�
�'{�2A�f!D��KE�G0CL�Hg���%��*�!�"�,���>x�(IZ$�ހ-�!��R�-�L���4u��x"�#_3!��Â�rv	8	Ѯ�*�fC�E,!�$BGz4��2�*(�c � !���*��+��9_�-�f��!�d��&L0U�#F���Pw��+!�ʴִٙg��![���$>e�!�$ǽir��  �䆶-���+6D�d2�)�1�$zb�D2 b�ia�4D���7��!a"Y��juٞp�2D���MN,>���n��ptp��.D�x�
�[��`b� �,m0\���6D�0��o��P�U"R]�x��6D�dH�i%aT��$��;���)�.3D�l�Ň��3��2��K0u��ؙ�)0D���6(ݹT!&���a��	|�Hl.D�� �i�*I�]�p[�A��u5^�k"O�P�i�.L���$�'7,4T�R"OԐ q��!鮔q��>	�<�"C"OtA@F��S�B��6�[	:}����"O" (P�����o�>xE����"O�����5�ժ�ɸ99ށ��"O�<��@ϲR)l��وa��=�6"O$��wb�5*�d-�C��%i�d��"O�XZAdC.{�|`��3l�(��b"O���o��@t��ϖ]q%"O���FAN-�����C��!"OvA��B%Wf<�Qt�V29�tuB�"O���� �Q��L�eč�r�Q�"O8���G�Z_n�P�"�u�\{�"Om��/ЪApH�" $˼6�ڶ"O,s��
*�}�R%�L��� "On�`2�_�N����1��+�݃"O:PJ�޾650q���N�Ql��"O^e:F`B K�ha
�*���1� "O ,��Q�eJpDa�l�MdD��"O��tf&�����J�;�"O����i��d��lM gZ��d"O\��s�ٶT��܋�`Y�jT��ڰ"O��:sf�5�F�ZS吢fj���"OVs$�j,��#N�? aF�	�"Oy+�n-�� 6��	*�z!)�"O 0���0+l`a���ڒ� t��"O�-��m��yD���+&u�ڹj�"O:��$QL����)X#'�ޜ["O&�b�!ٳ�V$�g�K��m��"Op���6.��p��}�(��"O��cpb	�SDղ>��0�"O�i8�_�M;6$�^ЪF"O�$iP�����P�K\z^�"ObT�R��Y�.q�3�N�]�R��"OP����$I���*�9�b�R�"On��d�A�VV��C)�r�A�7"OX�ȡ��
��iY$�5\��M�"Ot�R$\�_���7N ~p`s�"OL9
�׷hA�5��F,!yb��"O 4�cmN1u�h�e	�mS��Rw"O����&�?h�(��0Lfl�"Ox9�f�L`lȹ�fH>4���a"O��qD!V=DU�T1_�iż���"O��	r��EY��R��I �4��"OX9a�ޡn��a����s�X�4"O���7X���N�v��3"OzuAg�\�%7>��N�0	p�kV"O�0�_��Xᑎ�%�0�p"O\�Pʜ� �	'Mݥ�tI[�"O�m���s�)¶)Y���"O������1h#dD��oV*Tj�ٔ"O@���AI�<�d�($�׻,>�C�"O����.W�}�pK@�b3Ĭ!"O0�C"d� �#�aL%K�P
 "OF4��iX]�q&fE$a\����"O����
!pmS�Ń�=�r�Ȱ"O�('-�~�*��K��TR"OPJm[�*:*U��o�#�r���"On	[�b�#<h��Z"�0BVĘ{A"O\���Mbz4�QR�#BJ�=��"Ol�r��ʋ3���
��A `�X0y�"Oh3�����8��H�"�b�"O���+��@<U@���4(� q��"O� V���`��D�qc���D�0�"O���"J�:&�ηn�T"O���GM^�"]���+�j�i�"O���ΐP���"a�=^܎�(�"O�4�!A�&~4���o��zyΑb�"O��R`�>"�x{����m�`XE"O6dx�I2I������9S7H�"O���	X�.��x��ㅦnI�h�"O��C"o_�:�a���O22���"O|q�+��|�)#)���Q`�"O�8I�g2��0�]�r阃"O�1�S�]!���x���+��0�"Oz��ŁW�x0F��g��}u�Q�"O:�A��Ȼ2T�J �V��86�/D��t F'	����R\I�ia
*D��af��=�Ll�TaW,@MfE  *O�p�lʕ@���s��w�$� P"O�]��̔�*�T zg����"O^�r�A�^�nm�3G.r�A%"O���3C�%J�@`� cl���"O��`��G���5��F�je��"O �c�lE�1$�S�:�QǏ�m�<�'���t~�� V�I�DB�-w�f�<Q�t���JPm2�Dl��Xw�<��l��q���bρ=�z�3-Wu�<�6I^�'����W#k�@�i1kw�<1bEW���4��Ň�W���� �~�<!D?m��J���*z�\"$�{�<��@�m
r���Y�#�F�Zf%�a�<9AĚ;9���@�L>aּ-�5�]�<� FS @t�)P@���s�A[�<��d�F�)��k;WYt�6��V�<�B"�k�:US����"�V �r��R�<)�[�Rp�	�t
6F�i["c^M�<Y$ϑ<1r]��W#�B��v��E�<!��jL,��ݕ'h�pR��w�<	�`Y&�T�!�m\m������r�<�
�!w7�=�,Ȍ9��M3D�l�<���ڠm=�0�C���"�^E�CP�<�� ֓:�&ysL
&�X��&�R�<	e�_�2���^�b	�#s��LX�`Dy��5�D�s!�	�M�Й�oԋ�y%�{����C+�06��Ч���y"&J�xJPPx�m׼8͖�����y�o������$�oXP	�C@��y�eڷzy�����HP�R���y�C�Xq�A�F#4zG�4X5Y!�y҂ђp�6����"e�F��#_��y�ȵYT�qh ��5a`�Ȳ@ъ�yŶEq��^9Ws*�²�ߔ�y��P�"�m��KY�
4�.���y�!ǂa��AEL��6� ��y�-P�P�e��&V�s�̭��g��y�BI% �Z��3��8l3$A*�����yReĺa�&	���T�m��-r4��7�y���,Kqy+cd�m�L To+�yB)}���lTHt!s���y��h�[Ï�7�,2���y2�`l�3U@�a��
�KȤ�yB�BI$`C7-t	ك�!�J�<q2�[�vW��J&��!�����w�<� @�>*pE�4l��a~����`�X�<a��L?��������HQ��	�jU�<�!��f��)+3�"YA�(2.�j�<� �t[��_�,[xB�H��9�l�s"O�YY��ߕta��dg�( �dل"O�ect�ͷ7�xUZ��δ&���
"OL���ώ2B�n�p㓞7���BF"Oy
A�ӻf��IZ���3��"O�5��oA�;>>�h�.��b�C$"ObܣGIÕB1�ps�R�10H�6"O�u�������a�P:� �"O�,�dV�7�a$��')$���"O�����_�-�)�# �9"O�q3s��i�z8Q��U�-����"O�)��HK2g�Z���k��JY��"O�����?H}G@�-�����"O2�T-B;Y�n� �n���b��"O^9�w+��>��7�ޘ'rNҔ"O��B%�-N	��O�hc�i��"O��K�Ѣ;��n�-YX�h��"O�Prf"��_b��x��\%!�3"OL!bl(+�`x+���.�t"O=2 ��8,�"�Iۗ ���"O���A��c�<1� Ə�"�ic"O�Lb�&�7j]����~�.5(&"O�Qϋ6hH�y�$�o���"O:��G' �7�n$G��'k�(1�"O���l�`��(G�ލ1J.%�$"O<�C���$R0��)%�7C��Z�"O�,�cm�6}pِ����~Th���"O��"�b��y������
�YH|I��"O^����<q�F4ۣ�	�v�<��C"O`L1� �48ː��c](s"O`"0��E}p�gQ;OXM0"OZP���]j��`�e�:eZ�"O98��W��d���L)}�=��"O8Y�e��7 �D�1��R%N]��"O�Z����.4��$��	e((Qc"O|����4�y�� �A��*"O��B�~�5As.X�0�I�"O����Ó)~@)��[�i��1�"O���ǃ`H��(0�Q#o��(�"Or��D��5}-6[�kG_�i� "O������bL$\��G����""O���.( �0}!5I��l}tD�s"O�iR���&0��i�[�n�ՠ�"O�@ȇ�&ڴ����]�Rw"O։� ^�9E�� �L	�mTH ��"Ov��qK01�J���솨D\���"O6$�G��l��ʦK��2��"O��P,��J��t�)0�UiW"O��v!�?H�������"OTQ��jA2F�Zԉ!��{p��"OJ����:5�X�q�Br&<�"OV�.�#1>���+�5J>��	�"O��4ĝ8n+��@!��&:ԅ�q"O���2f�\�N����$�"O�%��V;<7ܭ:EA�<�r"OJIq���t!CV�� ��"O�qt΅Z���D�4j��9"O2�I�M� K�,��b���g��S$"O4�gżr�uA0�L�F���+"O0�	��<�^-XfA�)=G��:g"OИB�l(n��@V�^Ԉh��"O t#_,��)(g��.81����"O"������lA�]÷/ء|� ��"O�q�ޛ+�8P2�.R�B��y�"O� Fá�ͣՒ�8��8�\��"O<9jǣ|��Hk���1����S"O���8E�yЪ��H��"On�h����@g�lR���;.pH���"O՘Цݞ4�*��d�-m�a��"OE��W��Ҳ��vJl �u"O�a�Ab�"�a�seN�L.�Pt"O"5�g��$^=���#�5/��̮�y"`�r|-�"�D8�V�A`F �y��� � \y���M�|T�7�	��y��Ȏ��!��mq����M��y"��&Y��`�r�aB,8�ƙ��y�;j� ��:f�"��3)_��y�9Z��e �'�+Un�U��o���y�Y����QRA��ㆉ��y�͎D�=�u�I�H�6LF�yb�׏u����	�<n�ze��y�i�,K����5� <B�����y��3F�eQ@�%�)b&a��y�%K�(��D��Kx�a3䂪�y���_���+b�8?¼���g�;�yҡ�6v�����!"5}��M�ȓ'ZZ�!���+$��U�ò�T��ȓ%M��T�&�9�3�K� ��H�ȓ#��X��N�ow�@��*!�Z��� |a�Uf��z�D���'=�ҭ�ȓv��c���w��p�?C����I08�J:V1bhA��$Va��Gb�5x�k��\�Á/p��A��P�~�
RB�	h�ݙĆ�ZL��8[�jC���_�4�Qe��=7�Ne�ȓ�@�BT
�g)vh!ѡ8����ȓi&]c�F Z�H��X�\�0���;��(���V�(��̉�}��l�ȓ-�>T�i�<�8%�6gK�z��H��R[J�{�2�"���
��q�ȓfx�=��AU��ڵ� ����H�:	��J�S��X�F�)�,��Pr%;ToD�d2��"��/־Y�ȓ9^H@�J��-?E��l�58�чȓLֈ� �0����"��������d���x7f	�a�
�|`��"f�A�1�(B3��ǮD�i{���ȓ[��i�P֖�S锉U����:�
��קW�U$���|���J�'-�e�'�r�,��Qn,����'�r�@�N���pm��O�"�L�'mdԓ�!�9E�hJ�Y�d��8a�'��0b���|3L��� �b�,�	�'���p �:-yh|��L"(l����'� �C��Qe�b�̊�K�αi�'9��I%�ʒS
��1D��~Q�ȓڈ	+
� z �$:���D��M��paᩍ�+Mx|j��h�<A��P Oxj���t�d�� ��a�<I���\���ۧ�TͲ87i[�<Y��HsD�hs�0&�afÝM�<��I8^~�[�c�	���H�<ѡL�e�#�YUK"�sw��B�<Y7���J�Z��3s�<q3��H�<pl�?�fXk`�	�ݒ,�šTp�<Q��۰Z�ȸ��A�<hq Un�<!�+��iL���ʫ�:� �J�j�<�q ����=��,�,ka��˅g�<� �36J
�T�U
��}��yD
O7�'ZB���w��,	o�|
�©E6!��`��L�rhʜQ���B� `=!�d��{@�@��n��"�q�A�C�!��H�E��A��Q�v~��Q£@<P�!��ù13�(�'n�z�h�u�ޒIi!�$D��H���:Ṋ!�_-@!��ŝ6�juX�� u8�@R�YZC�Io�>��t�^�l��-@�>/�
C�əv��)��U�J���K�ry�B�I>y쌉ڦ� �C�H��P��-��B�I�W���T�	�*D�Zp߫(�B�I
M���1��X0KOTi��Cώ�NC�ɊE��m�"���*�s/�]JC�I�s�lXj�"*�$ѻ��ե|��C�I�A0L�ӊ^]�9`�fN>^B�0"�P�ó���|���b�`�0K�!��:ôA����%vj	R��@E�!��}�|%z�ȇ�e(�{�̀��!�O�yAJ�pcT F#R�cwʚ� =!��l�:���Zo>j�k��JD!�dP6L� 
���>j
5`�$L H�!�D�L��r����M����Y�!��D6n�ӡ!L�"͋�D�K�!�dK�\�R*��p��иt�I�z.!�i���'�##ڲ(��� =��}b��x �f� W.(q�bނ y�E��*O���@�ݰ>� ȁ��u��L��"O�yCv+�=j֬)�%K	����"O�ɐc[,JA�M*�j\��|��"Oz���FN�,�$<���W���HA"O�Ez�F�W�@r���%%�B5Æ"O�9�4���_���d�W�s�8U"O� q"oƿ�T�W`N�>lj98�"OʽHs�E�5TQ���yF
ɚ�"Ov}��+V fj�k!dӼ��"O�|3"���{N�q�V�A�j�dKW"O��A��c�����&��T��"O�a�H�7zJ�[קӯj��� �"O���EW�p��v���0̎-�"O"m؅�9��1q&�W�K�PA!$"Ov����V��EKF�ÌY� �˰�i)��䗚wv�$D��n���1w'܅r!��  ��:�g�A��"��&!���F�vE��/ġ-֒�T&�&P�!�X�p�q eҒm�`8�*��"<!�3�R�K�~C|��$�M��!�$
�~�����mO��iB�#]�!��ai����ۂjH��w&��M�!�DƑ}�@�{QoZ�䅠�F ^!�dA#�:��c�e�0�`b��#y�!��F-S��ܣt�me���6J�!��E�
H4��ˎ0g[2�䂀 �!�*��%3w���O�$�Y��H�qOܢ=%?�
G��M�F�*�(('� T��z0l_>x����7
`�Dc6D�4j�!�> H}�"�ޘ ����	(D������k��9��'����k7K$D���UiX�e����`��U点��h,D���ԓD,�u(s,��{p�{�G,D��x��̊@��2�o�`V9�pI$��hO��� �4�X��|�����-~,0B�	XF䅻��>�H�I�`Y�=I�R������&[�  ��H)'���S�? DXaAȄ?d��PP ���� �"O.)��e��[�d騲/ܓ5�� ��'��ػm�� ��bF�b�2]ʃd�*�!�ػ�>eRqjO�L���r#�%�!�D۸ d��#XOuh��C؏�!�d�_o��y�+Y�v]b}�c��/�џdD�dMʜ,�x%xu�	�K�����y ���U�t&�2�0Z����y�JW�i�mz���z*ƥ��L��y��B+5<��v �sa
}�ǃˠ�yBĜm(&y��ǌ�<��(��mH��yR*C=���N�:�^#�EK?�yb��$��K#�]�-�R�B,���y"���O��1(]���ᎋ*�yɁ�V��q�m� a� �Q���y�n͙r7�𑤨Ǵ(� (��yRLM9�b��C�L
�P9d�\�y���&E)������0 �>�8W(�,�y�K�mz��ʃ��"t��K����y�>�6����`����P�O��yB��<n4�fAM�\K2q;S Z&�y��~�pB1e�� �>�yR�YaVz�� �(Qs��\0�yBB����ç_�{a2�+R$��y���;(��h0aK�mW��	���y�n,e����L����N/�y�3���5��#m�}�D���y�Z�q~��sG�V�vŻA��yreʋ=����e�·g/\)�#m�y�տA��Ȑ埏\���kC�3�y2��8 ��5�3`�@�X%�����y���_���1q�ڒ
b�{ө_�yR�ϧ?��䨔��Ml�!�kD��M;�'B���MڀJ��p�e��4j�h�'P&q��'i�u#ķ�l9;�'�ƌ*r�D�z�N��0�uu����'g���-_$�X��5��;+��Y�'��$���
�Q"��J�:~nlB�'V^����#Jac��F~����'������� ���.�}��J�'��+BE�4$�~���م���`�'��-�5D�L(�	�[�WyJ�'׮����Ҥ,���g/���zl�'�U#�O2'>�ੇ�N���@��'�}��� �x��J�U>Xx��'���_	:��RWN� U�0�	�'!���e,Z pH��a�L�k�'j��()AK[�s(��pp�'T<���晁A��=قˀ�\H��'�T���K(p2Ż��FT݊�j�'7���!J�RѱE�X,����'�H��ӌ�q����@#�����'Hf����\�>���{�S-��q0�'hJ�U�'�L�Y'(��(� �k�'I�����n�\��!�ŚH�U�
�'$f@c�M:�|���{��
�'���bDŦ]J�<���Z6�%oM|�<A��H�|R��g-߰cy�Y9ba�z�<�)]I���q�!O'JY���҃�s�<�̿P��P �LE��P��RE�<� �h]�ı%��m���X7d!�D�	O��HA�rO�"V�Œ@U!�)��Q4	?7`t�9uH��NS!��¡v�,y�, K�X`�6�#K!�� Z$��&�H�$% kB�}��y3F"O��B�ݛX6���F#�z;G"O ͓TA[/VL�0�)��N���bd"OR����:41�=�(�tߘ�x�"O�1`��6H���Z�V�C"O8��! �Q��ڵE��JOzuҲ"O����B�1#�u����:-C��sd"OƄ�V�γ�N�@W��h�m�7"O��k ȍ;��)#��ݾ#��"O� BЭ-i JA 2J��v0�h�"O8�
F��4H�e� GU9Y�Ъ�"O&��鍘:��P��E:fO���"OHI0��AnE*"��YY
ui�"O��ږ�
�D�����fG�>hy�"Oґ��b�T�@]���ǉr��9�"O����BS+"a
��H9:�"O�0S�a�?{���Pk84}\�4"O�i���H�oM����I�Ik�	��"O�9�+��i�&�HD'��La�
�"Ob�6]@��٩��&W�z�12"O("�a� ,�&�Q2�Ĵ��"O�P�FW�$�cd,I6PcTe�"O�l����T(D�B�P?-Ex�Y�"O�����<U(BQR��R�ؔiB�"OȐ�2#�=���*5	�17��	�"O:���MC���h��H[�7d�Qa"O
���L~�Ų�(yԜ`k"O�H����O�z���9�"O�S�1b�^�J3*�=�&I� "OhM�W"Zo�aW���B�Q�"O������B��@ᜳ:&��{e"O�mhW T�����`ځq���"�*O���íX(�4��ꅶ&o~���'_.��Gc�)7�E���F�L�	�'~ �(EEP�p�4`� nR��	�'�N�@���'e��ݘSD�� �����'ov�*!�03��3ä�ހĻ
�'��Yt!ǣ����1FI�$�����'�P5�n��n\�a)a(E�t��'?�m�G��@>Jd�e�ߣD�BA	�' ذ�F�޷/<�Z��֬>]����'D�ؒ�G�?d�`���n�1�h���'r�	�v�*N�YHDGϐ'��u��'=�9)��F���s�ˈ'lPp�' �se�P9��e��H d�͘�'���8T�ܴ/3���Q��?�B��	�'aڸ1�蕺VU;,F:IQ�m��''TyyS�+1v����%��N�a���E�X�i��+B��`�GF���y�6�*�i��7&�(M���M��y�&S���Ǝ��Ĥ:��4�y�lb_Z���G$����F4�y�G̈�4	�䎚��f��y2��)]zY��,5-p�XGH �yr!�"O��@�T���ƙ�y��	�N"(�`�� H�P}2�/�yာdCzM3�!��V���s����yB��r����kY`%��kI��yb��1<N^P�1/��d�z��U��&�y�bW�E\�X�cY*/�-ғf��y�E�E]��R6"O�x�N	�Ř �y2lF�h�j+��.j-B�s��y��[$T��ɺ�'��b<LрRĈ�y��AlL��%�&Xͬ��C�y
� ��Q��!k�zYbG	E3=.��f"O-��f����a�ƝʨAs"O�	8��/��X�GU5]rd�v"Oΰ
�I�8�}�PeĹ#����"O�����D(זQ	2���p��� "O"l��FP[�8�bԮH(��	E"O@LK [� �aa�۶9Z�H�"Of�35�8#�X��!Y�-n�)s*Op�bU7��}qa�9pP�P
�'~e���
�v|���ɛl����	�'X�hC���
[,���� �b���'Q�Ӱآk�,�i�1_��U+�'��GL�d:`4�8aI �']�IXT>H�$Q*�
B�Q��\��'�`��ӓ(��Q����N��I��'�l)3KK�;2�&U$LTš�'��d�̿vݼ!;�n�9J���{�'eF���/�/�.��5�]�9{��K�'��E�&�'8�Vt�
�H\fX��'����'�q~������Kt�D��'�$�
������PX��'�NѦ�<*�]��*��J��]C�'�.`׀&l&^�T���F�`��	�'&���e	��e�R�bK]�>����	�'̒a $���6�QcM��ua�'y
5�&@�K�dm���pP�'�T9k��6��[!G�/rI��0�'��y��}����7HJT��d�	�'�rqP����8��#mH�'�,â�L
(,��T#��-k�'`�d��T)_~(���۷²P`�'@H��d.R i� `c�,IF��
�'�^��%��zvT0Qa��9H�
�'����aNɗk�Έ�Y�Di���h�<P��?��$�LİF)�d�<a�}����r]6�����z�<q���_�Ub
͛]00�hu�<)UC�>v����!�:�R���s�<���&�xS�MۻizY&��h�<y��4��"���:�@GFd�<YA"�4A�^hHІ�-;�Ѣ��I�<�DY!X"�8'�^�C���EN L�<���ǨW�^}�%�	x����K�b�<9�̞V��b����i�JEȀC�b�<	"b�0y_�5���6�hǄ@f�<�\,P�r����_�T�s�QJ�<I�-ߧ7ԸH�5��1+��aь~�<�Ѭݫ:_�%�D*�-:�<M��a�<i�� �F"�V�X�����nCa�<!t
c�d�وE쑠 fZ~�恄ȓz���a0.ƪ!d���GK� `�4��C�,�:�O����՛@H>%�x�ȓG�^E�U�K�R��{���!?vy��%������]�%f��W�ރRD��Jk�+S�@"�I���+H�u�ȓ0*5�a�U}��%��R�������"�'��:}���R���}P�,�ȓN)�l�X:Jx�m�A�i�̴�ȓ1
Z����{�xw˛�?�|��U�\����c� \`BfC�_:T��ȓ+S!{ቌ�@�xS��9K"���C�&\���
4@?v0K��*K&�Ʌ�J���A̬$Dޡ�%*3��d��<�x�����/� ��&V����S�? B,��d�@QYb!��X�aK!"O����EA�2䣃��*���"OuR�f҆G�L�����9 �Q��"Ob�ۇρ�%L�Q6��tZ$iH�"O(x� X�?�4�����"6&�@"Oh�A�-�>i��p�f[����i&D���&�Ӵn����^z� ����)D��!�T�.@���#)i�#D�(أ
X�\F�L��cKa���� D����!��B�!H�=(�TJC?D��� �L�S"ԿlSv�p/+D��w�^�� �4��9Y^0z��)D�D��F��=��Tz��d�<̀�5D�8�G��b���n�wF�o�<	�+�<w�L=`A�ϭ}k�t�3k�a�<�1@����C�B$$j􁳡�S�<� ͋!`�0��g���w�T} mEL�<!PLǱ;>R�ơ��PNJ [B	H�<��NbKT��O�|�,�Ѓ�A�<��v��٢f@&���p��Sx�<q�Q�;�Li�p�R�(�Z�<I�ޙu���F�7^���:B�US�<Yף�F��P�����0)��L�<�d�+i���� ´�H%��L�<��և��yx#e�+)�.����]D�<��a��^�4��ЏC�BGl0{�+�}�<y���
 ������G)��"�Ev�<��nO��q�	�~05Z%_q�<�B.7+��cх͋aF����_m�<)c�h�d�D��c�|�Y��n�<IFD� h" �tJJ�2v�q���t�<�Ԧ�� P��0��K#v��B�f�<�/�m���D%@-@$��r@D_�<	D'U	&�􀃠��-���B�<���-r����#�Q��Ʒ I�{�<�7G$s�8m0w*D�ּ�3�Gw�<�u�"?y (*%&I\2x;���k�<Aϝ�� �0IR�W��-#/�C�<!�d�.��3m�U��B�N�c�<)�DW��t��$�qv8� ̔X�<q5!B&!�E�AT�p�"Q��DVl�<�H��*�<�@5�6{E<�U	�e�<Q�)�`lA�Gb�3ch2��k�<���H�p�(�C6�>���O�i�<age^�/�Vy��'\V	�9�(��<c�w�� '�ՠ$��I�Lv�<aU�Y�h�Ǉ&z��3%q�<!5I
�-N��@#�<��2A��k�<��̟7D��89(�9�lA��(�h�<YaE��M<��d�W���l���a�<��ɍ�f�X��%B�mb��w�<�����>b�� eL�p��ؒwJVu�<�PM�$M���I�mMm�f��T�t�<Q��D0I��I��$�:|p�oo�<��W�vp�,�h��oX��d�Un�<I��Sc�d��SFȹW]�%�&�Q�<P̒�KZ͓��_�YУG(D�̣#�n��d0��eg6�#��$D��ic�ӆH%�D�e[2����&D�l��jl��
5��> �a��c!D�(9��J>J�D]���:�IqA�=D��bB×�p��A�悭9�]ZDB8D���nB�QB2�rB)n�.m�q�9�O����O�Z��":Vx��M���Që�<y����=� ��/�do����S�GSt��"O�DxD+��z�ZP���^�A�XLj"O�X����h_��c�2l<b<r�"O�BE͌�A�� �dQH��Ղ�"O t�Gƙ&h�$	;��/>Ĩ��*O$@���:�8�!�O��1�'�� ��w����#�?>"�ç�y��'!Z�c���#��^�ay��	�'w� �*0�i�HSR��]��'t�Ѫ�c�{SZ�IlA[�'�N� �'7YP=�"D��<�B��'�m �'ΐF�vqyA�W?9b����')"\�U�'yfRQ/Ξ,��c�'StTj�E3;N�1ؗτ�:B�ݳ�'��|� (�2dU�L��ʒ9d|@
�'l����#)?������dA1�'!�\`���_�h0�TK�r���X�'p4�D����]��n��Œ�'f|pJ��:�[��F�d��s�'�Xz��,qg�h��@�+[��!��'����f���r=Y�_�
��]��O���DV�J5v����P���Â�d�!򤇓�]ZP� p��$a�8#!��$%�%ic��!sP:��f�E!�Ȕ$�=S5Ϛ�T9�H�G�(~!���vbx���SH&Jiq�Č�!�D]�1j��!"�7' ��س!�� !��R�)�t��Gᕹm����b.���1O�D.�)��/`�`+�<	��,g��C��''�D�R���{8�q��6�C�	��[�C��4�:5���
�xC�ɄZ_l]���\.��@� 9$B�I�8X�9Iv��-y�@��'��8D�H(qOޣH�&�v"�-gݢ��1D��3qF[55�d<�U�_8Uj����%"?������	�
�*$;�aY`OR�?�4��"Oj ���Ác��1@��^�}�z��"O���E��8���
�⨠j"O����ⅻUYx��,W�;�ƴ�W"Ob�3dƐ�4j
����c�d��"Oz�X7.�Js��!�n�3~���x"O�{AO�()��4}1r�ǟD��h�O%���W+C�s�n���Y:&�Y��'�X�ؗ���>+4Ii�`M
<-��C�'�����*zDR\2Vc�g�l�
�'mr���%B[DyK�ʁ%f0J
�'|�"O�?(z�jbE�~㎨
V�'D��I��%1�@SM�~�`�KG� D��{&i�#Q���9��CN`y��?����|K��ǑmEd�z�6�� #�"O�U�&�ѱE@�&NRk���(�"O$0�E��1�
�Bv��I�`,V"ORd��o:+��0K
w�^qB�"O��#r�K��IrF���cd�i�"O�I�a��~���ʒ�%G�&l�P"O�1��Ƌ:v� �EЈ-ش$Qg"O�݀��Ye3�ZĔ� 3��x5"Op�Ҕ�R~�v�a2�
�V��%��"O�;��\N9A�ڪ<���ٱ"OxJ���XC�5 uM��J(.l+c"O�{ 	�_�*�0���-4����A"O$9� �/�zt��� ���	M���)͑S�p���=掭�I�+�!�ά t>�T	N<yھ1����P�!�� ��AMQ�kX�e�U�ڄb�UJ�"O^��
�$$9�(b�h���>�C"O��@�@P9_VH�R4�I뺌��"OΘ�!�T<�J∔7��	"O@�����4#p�͗bf(��"OLx�GJO��+��C��d��T"O*�k��j�z-��b��Smj`��"O�T�W��=r�P�K�!�M�.uh�"O��:f$�0=<�;�3����"O��a֮�'�t��0��F��G"O&�q7!�I,��c�׊me��b�"Oj�`��3ڴ��Ԡ�)8�9f*O��q�@Ls���d��TD��'�:S�H�G���V,ݭ��=��'��$S����3Ga��$�-��' ����!�`���&0�C	�'�� C�`ڊ/3��@ժD�v��c�'@ Ɔ�KҐup쏨B����'zDcr���:`z���gK���A�'�Y��阐H�yb��#��%�yR�'�ў�L���TMP. ���J�ȿn���ȓM��Q۱F�P�l R���5\iR��ȓ/+"�!�ƅ)8�hV�ٱS���ȓB����V���m�xă��/f�(��T�	���"Q�Fd��צ�ܜ��p��� lR�-�y�ҙb&̆�*�)�G,�b��@?y��Y��iUHz���Q���R~�Ņ�i��p�7�a�X�d�T
j M�ȓ�PuЃ��+s#�HЂΒ~����
���c�I�������F����K�IJ0�n�^����k��Q�� ��j���\�C�B^�LK���ȓ1��!	��V�A�� �	qr��ȓ_��<JS�	6w�|��cF[N�e�ȓ`e���}g48��X;�|8�ȓS��aГ�ǆA�@�A�x8��b�*� P��@��I ?V����n����+f�07�.�Dx�� *��2F���I1���45�ȓ|L&՚"�4H��8�bNFG^����s��rp�� 
�Sc�Ć'UF�x �1D������`�����.!,�.�("D�P0Œ�����/D�ΠP�M D�\B�� ����5TĂ�I%- D����F +PC(L	E��<�r����(D�H�e���Ph��Yq#խC�@�G�;D���%���y�dpa�&N�6�hԭ:D�T��ԍx�ԡ �E�j�,l�.8D���FMٷP�v�åa�	���8D�����,P:�0�r*�&N ����7D�谈֨6V���U�ߠ*��+4D� � ��M�N��w �,����e4D��`��~�ͪ��S��ثSN1D�Yw�B�Qo( �g͎|�nqc��3D�h�CW��v���˥FYX�9�G0D����2L�DI�NȽJ�Z�m"D���6�[�pV��A�z��\�`?D�4�gL}p�*�aG6B�"d���8D��
7G�/m`���co3��*D�Lkҧ���l�FL��#���En3D��H�cKbѪ����6Z�Eۄ�;�i����/ͩS�R��􎀟�����;D����ę�#�E+
�'��R�$D�� �A�A8I�ɐ0��c��<�`"OҠ��D�'+x�	B�DY{r���"O���,½Q�MP�+I;$��HA"Ox��4�Ԣ���zR�ڞu�&x��"O�L�&�*�n�� (�����"O���Ť5�z�0eژ׌���"O���^�	��Z�
'Gtr���"Oj`Q��W�2�����ɦ7bHPs@"O��f�T +t�lC��:��"O^����bJ�x:��W����"O.��&lV�`��}���Ӈd{�I��"O�3!���" v��V�[�OaȬ@"O�ah��ڪN�I:�ؚ;4�"O`���oF�:ֲ+V�ܠ4�<�X�"O|��g�2sA�����O���S"OzE�e@/1��|3�L?X�~�"O�dx��L�8)���eȒ�Tq��Z`"O���5�be��r��x4Z��3"OZ-�0�ӸW�1�@*O?6Py�"O�`�G�^�o
J���!z�"̻�"O�S!��H�<�hU��d��І"O����ۘ5^X��1�Ba�r]��"O���Z>w�rHBb
�l��ذC"O��rʛ�~�r�a�h��QĽ�"O�(@�%uN���N[�h�pG"O<��v$�%1���.�#�H��"O� �1��	�*��1�ȶI�<pb"OD���|�N���r}�x@�"O*ԛ�!DJIC�=lt!3"O���v�|���p�EI� ���"O	��B=���c���>1%>y#"Obժ��M+u-$L�E�ǮU�`�"Orܻ���o�|�k@U,A��$+F"O1Bu=&`[s)P���"O�i)���)C�ҥo�>*ftl�G"O�\����'B�P���2`|��"O�� &��:�`��H:( �"O���/Ϙ0`á�,4���"O�,C����� �k%|w��P3"O p�ˀ�X�����,wX�uq6"O�8z* =#�� �l�
T���"OJ#BΒU�z��t�B�
]�@"OZ)��bPv�R=�w*�3l$l�"O>\ٗ��Y�Hœ��Z
{Wy�@"O��k#�����5*S'עN�LAۂ"O~���0x88���HN�@� ���"Ob!�V��.Kq4�b�+?�,�"Ob8�U��$-l�6G��+*Nu�"O搁4D�5��4s���6D̀��"Ot`@W)4#�����چW�h��"O�1ר'V��kck��X��"O0(�W�Ժg�0��I�ڕ��"Otɑ4ó��� r�ھr��� "O��%̀'>I�t�P	��X`��"Oj�R�.�N}k�(�8c� �pd?O���$���*�LT!/O�����NG!�$��?@�`bg'��E�堣��$�!�G��ɤE ;��C�&H�!�����E�ъ^�d����u��z�!�DH�HQ�'I���S�A0�!��4G��)UKT�	izU���@�B�!��/����$S�XV�X���3�!�H� ,2};��FEr�*vAA�Ff!�dQ0'r��E�&�8�#��4�!�� ��1���/!yn��r�~��`�"O�g�L�f�R����_�l,:q"O( !��v~�k�b�;���"O��1�`�V��ʓ_
�H�S�"OBi���� �q��8���F"O��{���H�tS��֨8��L� "O\�1�Д)i��"e�2|���[�"O>��R����1���H�L��$s�"OJaH`�?t�F5�%ۗ0���	"O�	@a�)g��9C�����b"O���ֆ\V<̝��m~��p�"OF4�b�5|��h����Ct`A�U"O� ��Lǃl�V82W��7W�4	�"Oh|xf�Y�u�5 O˷���Т"O� �`���5�����/ǨEk"O��BD�
>Da��2$���4"O���aov]v	A$Y�����"O֡(1���<"T��B*�,q6��c"O�a�o �Z�l����h��I�"O\!����$ZF��vl��"O��t$�C�@)vf�M�A��"O,}r1�
�w|:�E�f6�!�W"O�����b�`�S����s ��B"O�dr���N����p��	`6X0�"OP�kƌ[�:k���/N�Y��Q"O����H�t�f`{��%��8"O&4{SBE�AP�<a��K_猔8"OVaC�Q$_��L��C͞z�*�"O�h��o�?7��l�6�ٹeb� 7"O���$�+���H#H�K�L��"O&����qh�� '��b�(24"Ol1��n��9�����G�DS��"O�ȱ!
	��}05@9K��8"O���3�� ר|�%C�)X4#"O�M���J ����B��PѓV"O�%�AB�]�H��r)Cp"O��*�,��o�u�'�X�]^�"O0i�#�ZR�4�I�� Z��H�"O�u�6��7���d�F�?XB��"OH��"e۽K� �`u��A��h�"O �)F. ����(S�K�Ԫ"O��c��4�b����.85���"OY�.-O���c�-���Ч"O29 eH�1uh���K��Lպm�4"O���w��!B�z�*�(�`Q""O��V	ԽU�F`�V�-R�2� "O��"=����W��59�@)�c"O`�sS��+�������$�4!�"O2%�`N�+3�2!q��ѐJ�,�z�"O� �6A�'��P�wߵb�����"O�`�чW�]~�����5-���E"O��"d���\?F��E
��g�����"O���'�U;y����d
Ҝm'�z"O���G�D�)E����gӦ1*��;�"O�DY��IQ�E �^��`�"O��BT�o��L�`/q�(`"O����,ko��`�!B:W"Ory�v�%'�h,X��"o�vHH�"O6Ej��Su�V�H�Y���4"O 8JwĈ�9n�0@P�֭a����`�<����i���P�l�l��%�d%U�<q��d��C���|#v�<��LG�z\��v��&l�(�n�<�AK�Bb�k
x1�qK�0m��S�? \���`ӿhQ��)��"j�>�	0"O���VA�.���CO Za�A�!"O��[`S-iq���0��Tq@"O$@���mˠ��V��W��t�U"O0uk0"ӽ&�9�'��2\�.�2�:4��d��x�R6%[�9��ᕏ;D��B�`4F�����ޕd+&d&B9D���f*K�=�	{I���keA"D������<|�b�a����Z��;D�Pñ4А8sU&R.UP�u��:D��8���-d��ʯ@��KSo<D�L�E#{	B�+#Ɗ"�T@�E$-D��$`�Y6���`Gu�z��o5D����ί=�]+�m�fb���1D�(X� M��j}����%'(R$���0D�t�� '��K�i��V�(��*D��8"FD�|D���R�Z���i�L'D���S�ĺ&ʀA�b-�]4:|j�2D�8k��Ə(�0P1S�ͭ����.D� h1�aK�!U*o���Wk8D��Sd��i�bI��<U�"��!D� �+P�M/t��t���$���)3D�h0��<z�l�!�˅�&>y��2���I�r3j�S$�3/z:$��P��#<I���?�x���i�$�K&���p� �O-D����.*���V�נac�f'D��ܜGR��(�#��y�'D��Pq�߂r��ܓ��J�j��8Q�#D����a�Xf9x�*��L�ƙb h4D���e�=yb��7a�}�=��3D�ԉ�CF���G�Y�`�B�C&�{���O��}sp�^���!J�qC	�'���Ç���]� la7��B�db�'�9�d;)⸭�"�4k1�x
�'�.�ǧ��k[��`'�^6j�;	�'c��[d���}�0  ���A(��I�'��T�GDJ%I�p�{u�ʥp``
�'� ]	V'ŕ6�����1\�
�s�'��!��> 
�Y.Q�w*� 0D��P��:*�\0�p���y?���3D�� ��E�&�$� @PO�#��.D�Y��s�,e�EJ�2y 仔#/D�8c�P�ppQrfb5g��q�*D����,I�/��Ț���(q|�r��'D���b�&�
�va_��8�Ӓ�$D�`j��(_��q�۴Rp3�"D� ۑMX�e\�����>%P"�@:D��!N�&\+�x[�GY<c(
T�" 9D�x�vg�:^�}�櫙�y��!C�E4D�@��
̋T�p�y�j�(BXx��/D�D8pO��������I�6�P��,On�=���W�hi9� �5�@�X��V �?I���?%��ze��mzt���77�b���:D��� dLo& �5
��@R,A�o-D���BD-;>*�I�"� sv"��P�+D�|)D��q���AA,5�JIz('D���&�E�*D�C	��|�b1m&D��!a�	�#(���D+ݜb5�s�F$D���E�S�0�������d�bi�  D�8zW���q芍)����.5�5@?D�@Z���<�X�z-�j'��eD?LO��8�E��%\terQć7hR�@�>D��X��QL�x�&S�} �;D��r5Ȝ�E��8�0dH6���h8D�� Ȩ�)#�p	3こ#E�y(�"O`Y�I�B���Q�(A�#60[�7OF��9�S�OR���_���Yɓ�²� ��'&t���b�7�h!)#cҖ�%@�'�� �����jh�I9�!�w�<K�'��h"S�� ;LU*�z��]��'_\��S�fE��/�	"ޮ���'˜h�=_�q��͈�+~(��'�"#�a¢Q��"�4g�I��fC��O��=�O8P飢c�Jy T�]<G�=��'א��oNN��
tŌ7��<����'�=��k˲�j��	�=҆!�	�'(���s#ķD�"���˟�0¥�	�'�`�+�/N*ƒ$S&�./��	�'l�����q��5��(8X���'�^��c�G�}�����e\7.X��'g����ZK�h�I 0cd& �'���`�T�7�H�!/G=Si����'�$r��� $��!��`��@��'&�<��(�^����&[*���':n�Y���<���Pw!��Nt���'�-��H�� ���H�?�h��'K��
���btb=��-�.���H�'Y�@�� ��0��,����U� �',伋��)��A�֥O�%3�䐚'�ў"~:"RF؍�f�͉tp� �H�O�<ѥ,C%vsb��O�-A�Ԕ�%��M�<�CD��q;<�!f��1f�Ը�+�K�<ٱ �.FUph�aL�+܅@�G�<Q2.L�1��i�+ɟa��@3��G�<��'³W!y�mU��8�q�����xB��*�:�HU���u��Y�5C�����O�T�?�Gi�z؎-�0A��ZD�"�hP�<����)6�X�q��3Y�& 
��H�<�#N�A1�	�JZ.��0A��k�<	`�-1�%�6�ϫ/*⸠w�Eh<a��g�=�BfLo�jt*�F�\%�`Fxb�)��'Ga2�
Ӯ
�S�8m)��$�?��� ����$<C���"X�<d���$�<Y���γQ+���JD��"
b���s�80��J�;$�I¬���H]���,� aK�r.��	��^#5��C�I7$�m0A�*O6p8(��ݶt��B�I5'Ze�VD!W���
f"H%vX�����H�S�O2��H .R��Q)�����V�8��	�q5�P��[>߰��PH�d�B�IX�;S�U<>��T�7	V�r��C��4]$��3"U-.�V��a�Q�pC��2g3J�P�KG"F�D}bRЃ
D^C�I���i1�G�;rJ���΍(7C��1�x$�C�ů&�0d�p�@�q��"<q���?�ӕQ�:��m2eN� � �ì,D�H@�ݎS�(=���Q�e��%X�K%�?)������TW�{�X��1D��Q��`ʓ�y2�]1^nL��
&_��z��Ǫ�y��9(n��a	�HH|�z��Z�yjV&p(
��.?�(���k��0<Ɉ��"1]&`@	2Ar6C�N�WZ��O����d�<yM~�SD� 9Z4h�j�c �-�k}�<�"ʠ>�6kS������#�{��D{ED)O��9�0d�(�Z�P&�K�y��_Uu1q/«/�PE�F��y"�B)��Y�$���)�l���@_��y"��R8���b�~��b���y
� HX(3�_2V�PBE�TlT���"Oz��c��<n=rr��������"O~=2č��(K�z$�C:��(�"O@���A�������w���ɡ"OUi�KH�
��ɱq�RO?*U�""O�TsU��(�E��@P���&�l�<�	��
����cŌ�!�|۰�C�<1tb�0}[ȴ1I�=T�2!a�Vf�<�A&R&P� T,�%��D3g�M�<�E�ڡqb��Έ�<6��B�F�<q��60�X! 慃X1�,8�d�C�<!A/$%8�(˒�щ%�>�B#){�<�v'��[,@�3	�W6�I���s�<��X�5����$��6� ��W�<i�����L����X����G��Q�<9AӀ{1�Y�$�B=j�(4� b�P�'��?��`΂r� Ls1��|�\�i��'D���^�&<[�n�"�<T���$D��蕍ҶV�@˥٭�@ ��C/D����P!y���&K&�<X��,D�c�5'36q��
&p���P+/����0���@]�
T��B ^��"<����?YYF(Z���:�iڌ4�z���jh����I,t bP�F�KeX�[5,A1�B�IJ�,��(	T�H(@"䝐:��B�	�xd4\�b�ȔRzH��b�[�pxNB�	C�ܳ�f8k�F�x"Y4*�B�I6;\s���ftfh��g��z�.B�ɞK�R�Q����N4�m)�ӵjLC�@l ��,C$MۼAqeV�j9BC�ɂL�<� "	�qBs��&C�	6c0 -x�L\=6���X�H��bB��pB  ��O:C9��;�oF*QWPB�I���H�J�0�t营cD}$B䉗\��E��K��=�(�{��C�I']��t�/�T�ĵp�b$J[�C�I- �:�Q��8)��3��
�C�	1	��I�W*���(�$j�5\i�C�6ylLF)��^]��#.�� �Z�hO>�2EbO���$��K8��@(D�d�ԭ6�
�Bݕf�lJPE D� i���=��4� ]�W�L�Q�j=D���.6.� E[�G,�
�"!�P�I���u)�iQ���%g�g��B�I�ʘyE�ų�F)ӡ����B�I3q������Y`0՘f
�.uu�B䉤#X�a�qht�RUq���L�B䉟GH�<�1�I�4��+��T��C�	�]��u��	+zF��%1rzC�ɬ9�tj��S5Ӷt���E�VC�	�<A�*�x�J���J�e�$���c�ßhD{����
���6��UT���!B;�!�D�-z�����m�)8�NԻ�!�䖮<���b��ID��I�.��`n!�$R4m����O0�b����!�
��l����5���qD��n�!���7����Pr��r1B�e!�X0V1qL�=�|�q҂W�`�!򤘠2'�u3E�� :�$� a
 ]���ox��xS���7A��S�� ��0�( D�|yQ�Ңu>�@Z� ѓt>��R�m8D��&�f- 5����Esde �)D�x�P�ʽ���h�h���8��&D���,jR���ĉ	�K�ȈX1�8OZ�=� f�`p�P5 �(��Q�� ���!"O:)�G!��\�2��b�P�D"O����������+k��$��"O��{#�JL���2��9+�vK"O���t�H��t!��g�4�4"O�`A�ܢP�Z��"g�����"O6�����n�^ԁQ�.��E��"O0��o]@v�1J'�W���p��"O��ҀG�>`�J����؅UE�+�"OFa�,ҩH',R�$��6�T�"O��)��4bNt��dG�.�"O��O	)f�Xu5���{%"���"O��&ƮM�@�Af�C�RT[�"O*�y#� �g���j lμ9��aZ�"O�@A��S�$T�x��� �E��"O^��;RbА���m��0ʵ"Ox �ӒY�E��KA�gn�1g"Or��5I���P8�F`���"OV��m�&����␦vQH%E"O��!"-C�L5�0A�Cu�8T�q"O�Y�G�~a��y�����  ��"O��huJ�*C���:wB����塤"OЭ��mH�9ܠ(:A��)#>���f"O�y� �D-^Q)pIȰ}Ŷ��"Oz��0`�V�4\fΎ�s���ʠ"Oz��7��$"<
�S"����s"O�a1u�er�jD+�'{�Z��"O�ir�̓�5lheٕ����Jq"O\�ҦH֟.�\<���>7e&M��"O��"�G�a�ڝi �A��lr�"Oh���6?{`��5l=� 0��"O�����M)n�i�K�)B-�P�#"On�ٕ!�� �uI�-9h�+e"Ox�ۼb�F�قoі�4��*D��J���>�`��g�ΑR{2	��-D�� �C�o0y��%��c:5pG�-D�\�ׯ��=�R�Q�D�r I�>D���-#�*����»'��؛�E<D��*�P�n�M7k0zĄpR�$D��xp�S�N��! �Ƽ#7rE{�h!D����%�QbX ĠǦU��$?D�Hu���^��cp�Ƨ_D���c�=D�x�� �2�9G�ߺp7�u���:D�00v��B`"G�ܢ����:D��U�F�18����'Z�1��i�D�+D�t�wBΊA�����U��C�3D�4�V
L�3x�i[��A�F��(0!�d�)L����*e�P�TC�!��M>J2���%O�Ճ1d�U�!��C)�Q$#��,Np��!���*;nȹ`h0+`J���X�W�!��W����n z�(�t��	;�!��B��U�Geʵ���@��(u!�Ą<h������M�@�(%���,�!��PM,H��B�z�;҈�;*�!���0��h�Aj��5v�@׉�2R�!�)gJ��a�Ɏ�s�Ȩ�a'��4 !�(�*�ܴ&��z�f� p�!��@�%��KV�T+�1�Ce�s�!�$���T���<�hU��ُr�!���*��|T� ��$��-��5�!��9�^\)S��� �N���왲k�!���3��!Rc�_�<\�6�Xh!�d�8m���Q6� d��d�:'!�� � C���0����@�>ު�"O�%pvaIF]Ȥ����U�b�p3"Ov� D�Ä�"M"����uxA"O$�ǃE"R��qpBJ�W�#�"OfI�u&�7-�� d���b樐�E"O"���E�T�%g<}&��"O�m)g��E��̪�o��R^T��"O.qp�ϏJY�@萀6P�-�"ORHBa�͕f�� #b���v"Of�XQ傧t��pˤ��l��hC�"O	)$.�Q����co�%���b�"OΌ:v/ĻY���@d��%CV����"O�t�
$K�|Ā�j�8B-Ȁ�"OV���`��>#�(c$�2&N�;"OF�i��]�dtBV�BV�*a"O*�Za��J�N�2��B�Z�\�F"O�X��!W(�(�aZ26�B��"Olsv�/;M�MP����:���"O�xX��ɩ^�ƨr��M�m�
�a�"O �*�J]1_����� �D�jd"O�I`��ԙx`EЦ���`�ˆ"O�m"��6SZj��c�A!4 �q�"O��`�oQ�]��΢d9�@�"Oj\Hg	'!���*g��8:v"O��JD�}��E�U隭"Of����IҠ�3��&�V�K�"O�q�!��!Y�iPt&۠ �h��7"O��0�L�B�Jm!u�%��"O�����ƴ;',�`����DiA�"O:TjE�^$ d�f�05��r�"O�9�L*�H9 ���&,���"O ���*���H ���4�2�"O���!iQd\�EAV�]�v5Jb"O8'΄e�@U!L)�le8G"O��`e�_x�D%��e�84a�i�"O��A�cŖvV���$�AY��(�"O��w���޼��Z sSf��"O�1do�>���I��]�4n����"O��у��z�hm�P�؝Gj���"O��)�f�J����Z�-�xI�7"O� h0����ؓ�ޓy]�xP�"O}	G��ܹ�4`�@����"OV��eH��X])Z���.	��"O�l!WjG7B�tM���Ȗo�p��*O�(Q�E�h�N��V��%P�\���'
�:�0D�#��$?����'�F�f.Y�c� �Ӗ<N�X�'�j��fk7��i����?)�zt��'�� [�/, ��^PՂ�K�'.~�1&���v�"�E�<,�	�'�B]k'd����`E%�0����'�D����P�(�$��ā�+B�0��'��y����&h�p ��G�3ɰ���'J,�ÒG÷�&��j�))񒼚�'3nA��+��v���Y2?���'�鰒�ԑ^Z��@�՘0��ݳ�'EMrb _��)��F�%��1K�'��� U
�.nЁe��7S�p���'<�M� E�@��y���|���x�'bŠ0  S6�a�DwR>�0�'�z��ӨBm� DËu�Fh[�'�(E�6N�8qz�:�FP�_�`%�	�'����x�6��cˋ�ay����'SL������tm�2�С��X��� ��v�E�{�ѰE��-w ����"O&�3 L�>�Y7��0j�.:�"O�	��K�o�4��O�*u�9��"O�esc䑈'> ���Uwy���"O�D�b�����XPMt�S�"O`\�f��)a�Y��MM-2��8YU"O:�!% A�洓��	�!#��`7"O�@! �J�>-��*�0SdȌ��"O�uxA�'3(ՃQkP�iP[ "O2���	� C�H�	�N=^	��"Ofy�0D&\�8*�v�v�Yt"O�8�ӁM(0s�<��	�5�~��a"O���)#�R�� ���][G"O��"�R�PB�;� �O�v��"O
͋���&HJL(q�N�c�"O�`p��L�V���-
mR���"O�<r�	�@��;�k�P��u"OBQ6��?ad�5J�_$�3"Oʈ��/�8_�D��/�;�9(�"ON��ڛk�$�R���2C�.Ma5"O����q�<1�ՇF=N �K"O�2�M�H"`�Xi����c"O�����rvxQ�FB0^�n)[�"Oܘ��+�?|D�;ԧA,�`Ợ"O�m�E�VO̜ZF��p� ��t"O4���v�X�p�����CV"O(���JW�'��5S'!W�\�l�#"O�=�lQ�(�L�fT�2LLMrG"O�Qc��˟+����˖�DFF-"O��`��?G��B�ֵ�!&"OX�j���.Q����_�g�"ĉ�"Orb!�T��*S"�0�B<X4"Ò;��ą�p��C�����T�V"Oa#�LƗ�� �'#��! "O�qÊ�6S�֐�f�mN "Ou��ȑ�V�&,P`>fV*:�"O��r��&d���R��ٲ1��Uӳ"O0�SA5i#�I�g���`�S�"O�]����GeȤQ1D_�`=X�q�"O.����p�XǬZ V��@h�"O�(�u��Z�L�z�l�%k�]0e"O�h2���uh>-`��B(4u�܀�"O~0pT��b�tx2�<!Q�8 �"O}��`��LN�ݹ�bU|6\��3Op40Ӈ	MwА�ED�S>^�r	�W�<I�O�[#������*��V�]U�<q�
�X�y`J�U߶�б�BP�<�O�N������#czL�!��]K�<�"���4`}�!�^�B&xi1�AF�<a�H�
i��T+�C�!r$����W�<9"و:{�шQ)��k�\쒖�R�<�ǡ`��)��?�`a{�DN�<��C�n�⩡��ɊlT��7N�b�<��IG�E��y�@�,a��%��dg�<���J7bWB��CKk�Ի�d^a�<���ۭ3=Vu����,����R�b�<A��O��b_�YI�S$F�<���N�*	��KCnZ�}�zK �D�<a��
���y��Kw��Z0#�[�<	 ʀ&��pd��26�d
�d�b�<I�NKR_�IS���(���F�<�&�R,{��У�I�'.�%��� h�<�'(]�۴���.H��e0w�Q`�<��G�
����K�t\��6��^�<� ���B�S�P6�݁�� �<qv"O�a�P>`�������^�F��!"OZ�XÃ�;��aQ6ɀT�"O,���NB+>m�ԢT) �ްb�"OR��w���E�����R�R�4-{�"O�����
��Z,�Uj�0_��E"Oĵ�4�a8\тi_ P�R�"O6���:��Y�GR�!Ӿՠr"O&pZ�(H�|%��f�O+��P"Od\���o�1*g�Q��:"O�����]��n�S�̐M����"O���7E�躍���Vrtᱡ"O��F�ſH��1�+���J�"O2	�eˑ�HaC��]��p�"O.�q`)��RȘecC��:g�*�t"Ob�B�Y�XI��k#0C���zR"O���bF�@�*A2������"OL��צ6Q��҇AD  y�=�"O�,9�%R�rpTL
��'T��"O����I�B;���E�*�-��"O0�0�%֊M�tz�e�9O���"O`�I���dV�)2���kT�X��"O�ط��#=ڲ)����5!LL1��'�2��s?�*�ʋ(rU�H�W�Y�!�!�F�R�H2jiYX�@�S��'ўb?�2ƪ k^"(kbU{�бjg1D�\��� ĸ5���L3��FkM�'X�>�	=ug����o+y����ϖ/�:B䉟/r(PCKW�l��P��?	s2�D;?����I!yntQ�QAdYy��7,!�Ύ!l�p��.39�݂��D�!�3���9��42L�4!S�� �azr��̄.��1PG�?��D�sKK?��B䉎@N�đ�0�̃E)˚O۠B�I9_�Za�x^M�!���-j|B䉀D���cɘ���C�bI� B䉗 J <ZC"��5� �$Ѷ��C��'a� ��[$��X�Ѕe��B䉿um�,[d�7x��cUAʯS�C�	Z۠u�3A�`��f� >�^C�Ɏ�BUKB흴h"�Sh#5�VC�I�k��BU�Z�)� VF�*	�<C�I�Y����	xO��EA˳}C�ɾI��1B�WB������B�	Mbnx��L��!�~Yc�`��3_x6-8����IG�`��H0�׎N���'0�O�ʓr薠+6˟.y#�B��K]����d�>���Z$���m
�$�9G|���0C��0щBN�X�
� ��B�	�W��R�h��8��( ��G�d<h�IZ��h��5� 2Q�~pFN�DV��QD"O�4�j\S1p�	��д$���Y�"O�%���(RР������ %d�'��d�B�н���݇H-��hV��%a!�G�>0��g�K�\��1P-L{��xE��E���H�GH��bX�*��hO���ޣ��[ \�S���c�ޏ����<���S�S��B�^�H�90DA�`vF��(ړ\s���f��>�V�ك��$]�p��a&T3N�23 ��Q�=.�M,OL���y��3����֕���H=��x�(E�*!�"g�0q�`F>(D�P#fG�E�	tx��*���p�
m��[�N��@�9<OL�#�.�	->tqcqnF�f�Iag�$w��C�)� pez���6	+�,�����n�ܵ�p�Sy��S6�,I0 ^#��A�����<y�C�	3�Rp���#e���2�$��D�)M>)(O�b���O����>c�x�R��P��mrp"O���e��h&5G�*��(�T�	~8� ��#P>8\�O�0>��@f� D�` �J%�F$�
$��X�G@��'w�E�,O��3��څ6Ę b��$$F��"e"O�<x�e�����ӡǫ(*�D�"O�1�1ꑉQ5���E�$�<�S�'c���c#���9P��(��ȓ_�Xt��I�zp.!d�H�o��p�ȓcYH\ж�z���n�B"Fh�ȓm�5���^�gV�񧃪+�����$M�j̷-��i��k;B�X���s�f���JG'��iJ�b�x��,r��JuA\�?0�P
���T�ه�E������I�b[�i��'],(�h-��v�J�*�ުZ�`���z�$As��D�l�����7@�A�v��~tY��KR��|R�x�h�3:�8�	�-��#$d���N�Mc۴�?�%��Op���D+?�6*.19Xp��E	�z���dVA�'�ўʧ9���s�Ɲ=�t�2 ߐZ0ڨ�'�"e���81��]F^�(�NI�"��V�qO`��3�$��$��牱s�2����0I&�]����-����Ɠl�������L�}s�F��W� Gx��OF��)Oؒ����Ф"S�ڼ��ڌ;����"O!#��T 1���Ƌ@3FӨ(�uX�(2�Km�1&>�aK,2
�8 ��Hr�����$\O�b�q�X%,2��æ�>D���)"��q���)�Ē Ij��j]��.Ar����Fz���x�:��"�����K�MbՆC�IS���{��5w�̺�N2g�C䉮N�B �����G���ۢ�J�aj�B䉡?!$�C�'AeYl�{��
2��B�Ih�.���.bL��M?:�B�I�4Ze�T�ߵ Hb @�BA�B�!͆XK�/ּ]ZL���f�2.�B�I,>:���<]v��@�&���?�dD3o�t���
2M�,8D�Ɂ<�a|B�|�ხe�N���Oo�y[�,L�y�ŀ!rH�kqoOG��Dk��3�y���)<�r�XƂ(�X5Y����yBꔜ$ˆ4�E�ܭs��y�p-λ�y���RwVm3Vi�i��Qp�F��y���'+ �8C��5-\��Q�K�yR��#}ʡ��gľ���Y��y�K�-�F|�`�ɒ�y�qkɊ�y��5���v� <�z1 �F���y�h�8b��`�Gު|�����9�y�ȯ���� �pI4�{�����y�ϴK=��y�[p�d�;`L&�y�a�mJ8[�'�):��������>aJ�$��S�A+ӂ}��bN+lO^��¡ �\����X�J N!��e5D��3�ӵm\.Ђ�!W[��)%I3D��Plݘ&hΠ	J�;%��xs�0D���oT�	SThЩԳR��i��-D�ԠA��&�ne+�MߡT?���!Ϭ<��4�p>�EkV)����E 9�6݁�ʔV؟�+REP���xP�VA�)�����  ��V(dAs�Y�L�-��N��;!k�!��8����"���=���!/`��4a7$��q`���S�? �Y�p�Z��:���3F7$Yq�"O����$ss^m{���c�"O��
�Pq�Δ�dA��ILA���'��ɑ|a����/>�(��sC�# -�C�I�4i��sFB��;�AՊ�#
C�C�'iۺtQKR�r��3I�	BPB�	53�h	�M�>��G�\�i�2B�E65�Vb �l�%�?K��C䉂'�U�	�3�@��I�~C�	?U�l$Q�$�$)��E%׺x��B䉦^U�4���A/|Ǣ�C�h.C��/Qµ��'�Q0(EP�	��B�IUn$�R���.�(�mӅ!�B�I���'	�n# 2%��-̤B䉩e�2�!4��Uf$:bȈ"�6C䉦I�H����-���a'>VB�F�p��u�͠	O�D0�!E&�NB䉵OPȝ��g�'&����d���l FB��%��RPD�#�*}�N  �^C�	�HƠI��i�b���c$�$�@C�	�B8���Ƥ'����lM�~�LC�	*�P���Bĕ"��
���!_NB�IK��`�.��\a$.1,x2B�I�=x�0cN�9
ļ�fkF>��C�IW��5a���Jw�Y#0m "Or� ���o<h�BX�Gup���"O����3)�)
� RP��T�""O�@e�J�a+lɑe]IƬ���"O );D���3��X5� �#�"OF�WI��DU4�"��Ĉl��i�"O�:��5p�f��>zBQQ"O4�KN@6F��(�`��`�l<)""O� �6�3:�l��N/5vʥ3%"OH�hd��n�.�j��ӂ=��"O����8.Ҷ)��+�F�x퐀"O6p;p��-a�R�0�"���"O.qhW�Ԥ2|����iE�DϬ�H$"O:L�  ܭ;v(��!B��x�g"O�)�T�!k�E����>����"O��@�G�W����P �%2��(f"O\esg �
�������.`����"O�8@�'Q�|	Z�@р��)B@"O�9�뚇�܊v/ق
�@�t"O�P' :{� � ��<lP̢�"O\�bPn��>,v�a笔�h��Z"Ov"G�/ �BiM��Q��"O�`5�֞#�~x;�	d��0"O�\x�C9���(��
v�I��"O4�hA;-�pœEER�y9�"O���J P2�p��I�#�Dq�"OL=:����D�N-bth+ub�8&"O
ٚ��ەTu�(g��b�ހkT"O�e�¡�tܱ@��̷o���"O��j��K1�0�l\4k=t��r"OP����p�Zr�uؐ"O4K$��Z��(��Ш4�v��"O,�"� 3��X�"@̷v�����"O����&˥V�,|�boR�pb�q#"O�y:�a��b���s0	��JU�8�4"Op:�M1���P�H9L��i"O��R
�h�U����S6�`9�"O`��L�6�jPJ����!DPH3�"Oԅ��uSB���e�)wق�3"O�| g)7s��)�"�B�{�h�S�"O� �}�J�6<��|: l8��a��"O2��n�73�1����Sҽrq"OP@��+	_h$Al�b�:8ȱ"OZ�$�A�g $�`�	t;�)�%"O�4���_� ��P�cNE�p���"O�3�M�h�2I��`�6q�"O�p	D���rbz��M#6+ >�!�d�Ж���$?5�p�:tOL�x�!�D�}^=�d���[�6XH�Y�5e!��DQ̨�&V+�e���
}�!򄕦^xD���@B�걑S�n�!���%����%�=��ə�0y�!�>����ϷRxd�1�̪(�!��q�Q2�/��=]`��eT�
w!�3^�5��b��o(�Xh�cR$UO!�DU*0" ��`ψ6bC46lY�-@xB�	�1zxa�Ӏ�
#�~\�௖:B�ɱ.��`�v�P<hi��� �rB�I�n�� 'ޝl��\�c'��f�B��5�t1�s��&�X�:ׇǣUe.C�	,~]��yR�2��E�ᨏ�?��B�ɷb@��)RAM�N��(�.�_I�B�	�f	�� Z�M8��j�ɟ Y�2B�Ʉ;X����A�_�t�+�a�k\�C�	9�& ����+�>-i�A�WE�C�	"-最�@cʈi�d �6�^�g�pC��,�E3h���\\��"3E �B�Ʉ|�B��7ꉓx5>`��*�E�B�	�gy��q�	�p-�ڵ2h�C�ɞ$|����� �|�
�.V�l��C䉿@m�a�'��,g�� �� tNHB�ɷ^R�IQ�EV#Rup𢷩� 1��B�I-V����ӯK"
�>£'��b��B�/(1p�G� 7�
X)����B�I�����H0N���3�Aȗ"��C�0i<���B�J���e�c�\C�ɯ>��}+1.�9��k��D�{%TC��
f��I
�.޺�i#'�H�C�Ixd2%�ٓ0�$��h��C�	{J^M���B�����ǍJL�B�IC��4Bg���IЕ	��$ݦB��	� ��2�E��%
�ȆX�B䉖*$�S�G���A�6� 	s�B�I*	gtrPi�B�`� ����S��B�]-�(�0��7wĚ��sbZ�!�TB�ɝk����L��(����]�B�IopMc�@�<b�*4h	�6�B��)��q�
%Fj$W	M9hB�I�sd������ i#/!_l��>��)ǲ=Ξm[�	^s� 5Y��_�'e�x¥�*�xdS�B�(:��*r�ĉ�y���,S�8�Q��êd�ddA��y�)z[-���@!Y�a�?6�"O<��5��U��`f�¢n�$|B�"O|Q���5b^4� �։ݜe8&"O���^�S�0�����C`� ��"OT����t�H�sL)u�ވ��"OF�c�M� ފ�++|O�D"ODM��Z@ߔm
$�?-�}��"O�+`'ܞ^���p��׫c*�!��"O~�	4�R7��P���?|%�݁�"O��;0	ˊ`�=Kw!H�l�Iy$"O�	;&�U^ HXۇ�W��p�"ORȁ�bD<&�����m�K��§"O� h����������m��:|z8x"OΝ ��-@���y\�x �"Oe0�^��X��_5N��$"O�͋�@�B���")[$��a�"O��򖄐�U>"m��L�
r��d"OޠEH��z/�L�Í��`��"O��a�nЮN� ��-\G*�1�"O&��'���[EP��ӊ ���#�"O�����"+�B�	�L�V�p���"OTtC�m*	�%�3 t�"O�tg(\�A�x�5,F/5vXq�"O��* f���$���k��%���"O��qB6��܀$LVF �Ѓ"O�0 ��G�
P �4
�,<��"O�8f$
Lf��!��H��Q2�"O�H�ԇ�=V� #b��`H8�I�"O�\B�)�4�RDj��X4N	��"O�'+�}\�0`҈B$h��d"O�U��%K�~���Ə�G����"Op50�D��K��ձ�f�z�:�1"O$E2bO��� �KY)R�8��"O�5ae|��r���% ��8��"O�cQcK�Qm��CV�8�����"O�]p6k�0E��@��敡D}��$"Ol	۲m߮�Z��O�(X0r"Our��I�$��[g��zh�l��"O���E ?�,!�ZR��qc"O�`У���)�l�	5���s=���e"O���F&�c�҅{�,ɴd �Y�"O�$�y~�бv��/Sv�P�"ON�b)EQ�r}��d��}���"OF�����	?I�M���ct�
"O��pI L�,���#�.S�@�|r�)��z�H�7�˃E�����-1�B�I�L)�8Ӓ�I�����d�	!�xB��"�X;�IF9�1�0ɆdB��"M�D� "��6W���8��I�B���b�����I�~ى�햇	��C�	�H7���m�6S�vC��T�nl�C�	:4��pzJ<wZ1`%f�zF�C䉮4����+ӽW�����Y$d�C䉏y��Y)%l#[�P���Փ]�VC�	9om�" ��27�Ƥ�ą٩K�$C��*�x��������� z�C�I�OՂXSVc��ߌ���矊x��B�%gXx�LԦRAh���靣��C�	��������0���oDC�Ie����@&E�9�Ai��F�Z�C��'C��Ԋ ͛*�>�`�Z�|4B�/?)6\X����s� x;�D�xk
B�	�~��K���@"�J�^���AM�	I���\�0 E'X�]!��N�hy@�	6���;��:�!��;�K�S�fl�sI��� �N>I����G�G�X���j|��ر �%-�!򄂆�(Lk����8^��`^�!���=������o�}##�Y=:�!�$V�7�&����F�܉�g�ݵ�!򤍬'��=	���e�j�@����Py�	2�X�citj~h��Y
�yS�=�tq�4��*l-�r%M"�y�*�-/@L��p�E�]ż%ٴLF��y�H�h�Ra�t#��R��s��E�y�	B*���Z��X�!@�p{�A�0�y
� �\�C�ΏT���f#ڎt��e�T"O��ڄ���i=���� ����epV"ON��g+�-H�:�qA�� ��#"O�b�E�[N&{�@05��P�"O����R� �iV!	Đ-�W"O��i��Js�R���B�=�>eXr"O2A���'9�eT�Q��x��"Oi#ƍB4|�b1�pϊ{���!� �A���Ön����ӊ�!�D�:Cr���%����&9��(F=R�!�U*,(�)�iA8b��Mr���6�!�͈&���7MS�k�$�2EǴ^z!��Н-)�R�	^��CĂ (x!�����u��L������!,wp!�䂎t��xǥR'��LÃ�D}n!�U*k؄�G"E/h��8h#�N�xa!�d�4/5���!	ι�܀���41�!�䈧j�43��Κm$n\YŃӽ`q!���+��%9b�9^��,���-Z<��$�4��F��!S�5���	��yR��zV^y��#ԬII�a�v'�yB�/A��mf�Q�D�N��v쐕�y�g�;3B�\+�/�=��l6 .�y��9RD��玧-��X�����y��+B�!s�'5䅲w9�yb�F�68�a �0�L};�AQ�y�N�R�J �/�6̓����yB�]z������z&��6KJ�yBH�l����ܖ>��t5K�y򮋝'�6=�nW66aT ��O#�y�H+���Q�]��A��y�� g�H��c�K:	cvi#uJY��yr��1N��{6lǘ|9�з��,�y�L z7­ �Lîa�$�pG� �yr�� '��@��V�Ԍ�V�ϋ�y"(M''a� ���M|�BF�Y��y2l�l<��ir�>���2��ϯ�yOK���	�H=
$@�	��yr̎�|�j�{��� 6���#���y#���	!��+"*�q��"��y"�97zT�*��c:�0�#]�y2��~^�;���i����D��y�hB}�<�w(S3�\Uxpn��y�
=���	��ύo�Y�o���y2J�t��ŒeIF ��(�Ꮷ�y�ɟ)v��&Ǹ!(�p���(�y��<�:��EQ���`E�<�yre͡#՞|�AKԦF�b1�^��yrbF�M�� ʐ�
CWM�A^��y���4��0(d�4��cpI�2�yr� ��	�앸6�0��4�V��yh�,.��q����1*�@�#���Px«�u|X�R�H,	����.��M阵���0�bP�^8>��Y�Ѭg�R���a�n�0��,>��D�d�+~P�ȓjv|U  ��G���P�jڣ5~�Y�ȓamZA���O�aF���$	�]��Q�ȓ'dR�K��a�ׁX�o�np��/:@\�WeP�`n�<H��W�Y,����,�Zp����WRh]���%$d2)���24�r�h��y"�Āj��݄���S���5�hbDa�]�2]��H�*�b�ä{ ��)�CM�(�ȓ}�؅:��^�B�$�#������S�? ~T�R�	d���%�&B$�"On�p'ǒ39�CdR:m�H�$"O������r%|�۔��Kc��w"O��������mͻHphw�QK�<��Hօ[�X ���˲S��2��Y�<���ŧ'�`t�g�V�8��|zwD�Q�<��)e>Ҙk�Ɯ-Mܜʲ" g�<A����boZ�a�'nnX�0G-D�l�cN.J�B��T��5>d\3�I,D��SA��G��LQ��W;a��(D��BN�>R�Y�g�ɥl�
1���'D��S�(ش""���c�=p\�@��'D��1���?[��tr���x|���$D��p��XCL���K�p���b�#D�tS6� �Y4��X�i�UQ�Ki*D�����:i��qa�|�21�4D�8q����]�"a�4��4N
�AM/D�D2�(�*�=h��(uy���8D��� �O�f��Ń�&�<���2D�R���=Z! AP&��/�|�1�-D��Q�cO(M�X����x�|�!6/(D�T��dW5JV-JS�S�<e�h�	)D����+AS���'bΦ
�p6�5D���Pg�XV&�0���7Ёe�3D��`�쁉_b�M�⯔����R5D���3�[����`p%R���q�!D�4
���fQ�1'F�'>��=�T�*D�X�q�_X!ʅ����=+*D��S�h�m�Dj���d����0�/D��qT���#��E�ǌ8B�zr"�>D�tB��~�d9	�LC�4��"(3D�����,v=`D�-ʧ>O~\*0A2D�<82"A�N���
���d!�-7D��!�72�\�x&�����d(D�L�߹$y�p�䛮e��I�� #D����K�~��9Z$m׼/�Ji�K#D�Rq�ų|��bc\yq� 5O�#=iB-�$s��*n4rUgL�<�LR!&"���ɴH���U�QQ�d3�S��E5����09�{�>vK�a��n*��y�@�i%�K��J��=�	��&����-hD^�jFOQ��M{�dY*i�\A��+ΪhQJ%)�y�<9�F��(0���Z4B�Ĩ���c8��Dz��� +�M��,!QʜG�)�y�Y�P�d:�G�#V�Iq�G��y��@��d��)O�!�?�y2�ɨf��q�����v~p�$F��y2�G?�X�5��c�"hۡ+I �y�
�'
�j��
hD�g����y�C[<�~-i���SD����A� �Py2��mDQ$� �%�ynRC�<9wlS1-p T�f�кG��J�X`�<1�����x�@-e��r�&_�<���<4�~��*\�&��{Ħ[U�<!�!�X}~MJ%��5�<@�*�U�ɒ5�>D��'}$��w`��h�A��R���
�G8���P���S�eȔZ��i�p��3�b�Aq�;��@��ͪ!a��c�-	Eh\4҂�&ړ9�a��Hu�t[Wb1��C���E���~!��@��22,!�D��;J� ؊S��� 6o��M#�F ��@�s!�T��@�i$��%7\Fk�aɷ�I;��w�ٻ�y"�7j,��g�����Sh]�U�	���	��2�ڑP�����sLJ,nh����@&d��-p"/�O����`	�?�L$�
� ��!MG,ZV���D?�ȭ��GZ)�|Ȳu�'�Ѩ�x�:ł��'j4>��C1 ���Ŋ}�*ٲ�a�'�����(9��q���4I��TG.���O�36@� ꟬�n�Y���z���P�����aϗ����s�����A�/]�2'�(	��Y��h:D����4���ٷF;��4b�Lجr��I� ��ybP�c���!#Ô��t�'���A҇< ���CY�4<��E���'��,w�bĀ��� WjQv��Ozq�W
'>D-� %�5��>��I� �,�"e�>3@L���e�'d�t��Pe��$K
ya����Q>a[SX�+\@�q�y���Ju�0D���w���5����*��@����'"�zc`�#+^�:��9Q4艮~&ĀF��w�IÅk �]��dz�(�O$�)�'��5�7D֟D��4�ӭ�����^"~Cb�a4��9�0�������$T�\'�H�c��rv���=�Xi ƃ1�O����0�0�QA��z����gL�z��Dh��A��Lt�
�:s������P\�q�!u��ȁ�k�� Fy�!VR�9�q�����B��ŇW)H��ݴ\��\��A=>;TxDy��9O�#�EG
h"cJ�3���;��P�>�PAD���":��	è��B�Q?���릕�U��F�Qf�<I��ډ�p?Y�ӓh(6�)tɎqÌ�fcشW<�DS�@��(�$�h0�]�����1f��	(�Jya����$D*U*H+dي����W˺Q��Z�sC��;����)ŔG��-�5�P�6�z�'�S��?y���(��$I�'�L8rtl5�U�&�0!���0L��1�G%�I��2�{��%6,��@���~�|)��)��<�b�Ի�))�G�x�(����`?) �	=�hܐs ���� P3Vd1O���Zp0I�܀�I1�����%OMH��b*W�v�� n_�
66M�O6T�?+z��6@!!�<?y�)D=S��3��MYSԤkAm�Ah<���?v;Z|z�K�pz2��GCD�r��3��%�$�	E���'8����-�|�8��0��<G�$��	�~�6݃�x�+�옊�䆯g�@tҧ˚2/�k�!�S��yb͞~р�0A��bZ(�V���'\8�v��iB�2d�9��%�,K���U��D�a~"Ƞk�lp��X ��3��6�0>)`%Y~(�m!�-��HC�o��+6�2�'���b��)VT@Z��[�q������Җ9��$?ҧ8ֲ�h��C�ܠ�5Ğ7Sܑ��9�F����M�S��#P)X��<%��J��8$�"~�*Pr�_�w+�����A�K���ȓ3M
�����*Є���ٗx�-�k�t����=YcG��tHs�k�E�jD��a�}� �w���m,A��#�Ԁk?D�
�W�T�B�Ʉ-4���!��!�r���aӨ��#<U�>���V-��P��
#A����I�;n�!�䏔Y���S뀵KP\�AF
��H��@��O�O?牗y�� )@#�%��e�ql�cD�B�@���f��_�ʝR�aE�r��	��?�R[V��c���t�pI0�	S��'���Ƌ�B�<��W�s���B@�$D�h�h@� ��Z�$e����e'D��{�b��L��r%ծk"$,��6D�|c�K/hz�U�wf	#ܠU�4D�`�G�1]�����݋1'�0�4D�@��])D܄Ԣ"��3x�����`5D����G�r��d�Vq2A,.�>�ȓ*�����dL"��F���z3�"OЍ������"�^�8���"Oڑ����`x�"H\�m���9r"O��`A�O�S�&�k��ҋ{|���"O�����]
8����� F�ˠ���"O\����E:�E�� �@�L��"O��1B�Xp��`�81��ي"O�uᰨ���r�Ҷ	�5(�"OB��/WE�F��a�T�\�� �"O� �P��aĬ�Bs��6w�j�"O"L�cJ��t�[Ak��7�����"O�Z�G_(=B/O�<�P��F"O��,
bx&ME�g�5+�"O�ذÃG�3/칲DFVmv��"O���U��?r���§k֩C�<�5"O�`�S�6l� CS�D�X]�Y e"O��p�'�h��1"H��M^l���"O�:	6�,�)��F���$1s"O��;���<.�$�b�G������"O|�kdb��o�T�P�/brp%�"O�<Rs�M1x�U[��V7O �*"O��i�-�j�I���a/�YA�"O�!᳣C�9��+ǭڋL�q�"O�8���@�x�XH
��V�lՓ�"O���j��F@`�'�6nԨ���"O:��.Mq-9�i�2A���2"O�q��
�Y�0�H �ټ]U���"O�A���R��"dɯ+�H	�"OR��$j���9�a_*�T��T"OV�D���YQ�������,q��"O��1���7 H���-�,Pͱ�"O\R�F�*�*���-n�@c�"O��(�d_K��S`�[?J��8�F"OF��0l��72���"��	p�"O��Y��D2|s Lɧ�o]���"O8�;�!0w�>��!�`H "O��b�(��h�%TJ��M�D�x2�h���Oîph���H`b��ah̍x6H���	��Y��F�B�@a`f�ͣ�4b��;v1O6j�!]�p<��F�;wNI�V�Q7I�<�u/X�<�`� 5!�C,3��;���W�<�R	��e&N������ ����GS�<��#O�J���D$ȃ]��q;fI�J�<�NS4o�n��A���uk�H�~�<	4&!dhj��D���o�8�����z�<�uf%�C'��FѾD�b�p�<ٲ���eX��C��q��P�C��o�<q@�R�2�Z	����HN�J4��A�<�W!� u�blH�-� (;���w�<��\༻0�K�(�����m�<A��};������4��11G��f�<�1��
 �r�7��9w3��X�*^T�<q��
|�`5�qhT� s���NFP�<��*�:M+����~lV�9��^L�<-�j��dZ7Z\��+��D�� �ȓL��!��Eƽ
��<Ec��+�d����Q�׍d���B1�TIZ���T�W��
"\�Zg��x�<���
�vp "֯Xa�5��g�8rE�-�ȓ~��� JȎ#�RX�`^��yB�<D��z L�+p8b��V����!s��<D��C���!�n�y����tH���a/D��J�nԹ]���Z�"�'U��F D�TR�L�l����H�3��x�:D���S���O*-3���<!�FU{%�9D�Ц�����勠G
,?XI�L(D��8'��pH];B�^�[LȰ���(D�0s6-Ӹ%���5ŝ;Q�� �'D��炖O���"X�WH�Վ#D�lc��\�C��pꗉ/"����$D��7�ϑ@!:�kƨh���2��%D�|�փ�x�Tp ����)#D�pH�&ț,6Ly������0�%,D�� bmX�-��4�bw�A}���"O���/]Z� ����?f�0Ѹ�"OX	��!ݑ8�,A��4��P(�"O�#7��m},X��=��$�S"OĒ��׼��DI!�`��8'"ONX��@e�0��0a�(�6P��"OF��Քx�����B��Q`b�"�"O��z�/�?��;QAWSb!��"O �C�G�%�!D� Ij��"O��g�Ό<�y��@�LT��r "Oʝ2p�T�O�0�օǋSD��&"O��pP#9xw6��M�F�p�@�"Or��`�E�1t"�{s孊q��L�<�`֫|H�4h%���U���!�^S�<A��"0��������^m4a3e��K�<����+.<�v�O��t�B�!�G�<"J����}�� �$�#�nv�<�-L�r!�4�Q�
,A|��g�z�<��NȔ#m ��Łe�:e�3'Wv�<��$��F�$�A��'�4aq��<au���`��_Fˎ�x2��q�<���N�#�P9�a�I���c��h�<����<�ryS$!�y��H�STq�<Y�mO�J��D��/v�(ɺ!ϟo�<ɇ̟"Z�Ȳ�'I(E�MB��f�<�K�=6%���%�]�
���0��e�<A��y��0�\c��,�s�?D��ʁ�R*����͝a�Je�e:D����A�˒=�ڕ.~^�v�8D�����h�.т��J�,Y3��3D�[�)ѓu��6��2�v����0D���&����슁.A��^ 0A�*D��6�	��4T��%:H�q7 $D�X�6�#B6��gÝ$CEd���%D��,YZ����k�$��vm#D��i�d�I����B(�	�@9��*O�5�M	 `HV����x�"O��0�*�s�l`6GG=i��d"OZ5I�NC"�d����P4�Ґ��"Olh�(�q��P#t�Y�;$` 8"O�U�7'tH�r��P?���"OT=�5�Rx�q�O{�RıQ"O4l ,��~�B�k�;�:�(�"O����MNl"��gK�:V����u"Ou9$�	�}����0JΞhjD"O�D���9{$6��d�O/B�ҽ��"OvE���Y�7�>A)sȕ|	^���"O�� �vVy���:��UH1"OvA���L�aT�1�BƯj�� a*OX�k"��:B��+�NoЊ ��'Qr�;�lNr'�,��Bߴ[��*�'2���@�VD�p
3EE�e�y8�'˖��̊)]rj�(��A�p`i�'�zgC� 8�b�u����'���`��hp`�qe���
��'���)����q��q���DA�'�*ǝ*w�Hx�ȍ-�����'��ik6+X��dh%"Ćr�R=��'��8��
�2�؝ibB����	�'�`q�t�C�2����x�raB�'��I��KB@��pB�*�>c�n�2�'ٌ�8@��X�Ó��.	.� 	�'�� �?rR�P�C��t��'^���iW�H��!]/����� $᫳�ӣ��l����T�(9��"O H �L־o58��Y"y���)�"O�̳1�Q�&܀L`gLN�=�t�Q"O����lݾWP�ո	�����$"O8�4��G����ӋQ�
�ݺ "O��:��
�Y�V�bcJ\� ٨l�A"O��q��q��4ǩSh%l�	G"OE�fl�#}�1���6WI�A�"O��`�I E/E�f��"+�-av"Ofs%)O43L���qc��iDp �"O�y�A��+Yb˰	��p�B|�"Ot�2��@	L�(��?���1�"O:d�	�%.T�BD)�e��u2�"O�):�HҲ)��,�G�?��m��"O��#�L� %LU@��R/h����"O�Q" �>,�(�D ���Aڒ"O~IB�*#<�=@�O�cz�E�w"O攂�j
���h
� ή3���s"O� @%
 Һ���� D�b"O�-�d�7/�1��N>\�v��"O�H����sT���yNhj�"O֜HC-Ȏ��dr�6�P"O\�'���-�<#e��*8�&͉"O��`�86� :�ɇ6dH���"O\4�wn\8J^q�(�n `�e"O��3e�#v�`=	�L�<?@C"O���F�؊j/���j�[����"Of�	5G%�e1K.d��=AV"O�U⋬����� W,z��p�"O$s���L�]3r����ԫw"O�h�)����
�T 3�e�!"O.{FLƐV�E�-�6�p�S"Oμ����Z�&Cۮ7�D�"O�i0�f����3U9>#�D��"O��"��)�]:���3�	P�"O�Y��	L�C�ܜ�%���Th�V"O����Lai�эF�|� mX�"OpaHvEއ:��D��\�:��Y�"O�����c�<:D�D�O�p�"O���v���P'v������Sx�"OL3#��3�D���@{2d��"O����h�1���c�{.��"O���&g��x40}�sBӄg�pd{�"Oĝ2I�'�D�6� �x�"O�,�SF
)q���p0��22���yB�M�*�( ��H�D�nm"�.�%�y⅜�	�"|	B�M�^ء���y�`��
����F.��9�@0$�M��y2H�&.C�u�'(	�1���RӬ���y��2	zBHr�]!$� 0��]2�y�f�?���҃m	G|�b����yR[9��L	�m����b��Q�y��F����u.K�-bt�]��y�%�/>�K�M�!��y����yb	�"1�>4 �H�T�y��ܼ�y����c�y*�?�����"O�4yr��&�ѹң.bh
c"O�t0��ğ=\��I�$v�""O��@����i��t��۸�Z"OL��(�)o����N7'�p��"O�i�&KL�D��JR�,ǂ1��"OT��wLFH��s+ƬW�P�B"OfdV��z�����+�����&"O��)"��2��|P�)�9}�` ��"O� ���L�(^!��U�_��Y�S"O�m�4g_ ;���s�����ԅ�"O��*�Ɇ�D�����3���"O�][*�2n�F�����:|��5�"O� �f�C�}�U�,5V��8�@"O�MX�"ɆTU����������"O\��C�B��ݘ1�Q�_p$D �"O!b�Q0?x�S�"�l�W"O���M�z��(��B��ApX"O�gJ�*}��Lأ�B�'NRAA�"O��o��F�.����ӑ�Ja"O:y��Ƒ|$|dX����s�v8�A"O���Q Y�dqHӇJ����"O��wN�<�	Zb��(��Y+�"OT(���I/�&�3u`X�"���h�"O1�ubσ�l���抌�X�$"O����6C.M�Dj�v_�h�6"O�=��#.��1���B7-��"O��㲅�5��l�S��~.�X�T"O�P��ķ�X9i�$�Q ԙ�"O��B�M��}�H���;�"O.��K48T��k`'�h�x�v"O�Ċ��	 OPH��UG�<讴��"O�TSWJ9,��J"�p����'"ObU��!Y	O�,�������q"Op���Z'�Hq����!�Z��7"OD+�AQ=���!�d?��F"O����Y�f��xf�C��B�	g"O�]`���gB&��w�[�Bhab"O��b�D�$�u��N	J��]��"O~��P�_�[�nXR���<|�4"O ��%������wE�/tX<�X�"O�HzaM�0�Sa�å%BD�X"O��c�L�bh�tZS�V����"O^�i ��91N����Z��Xt�&"O�}#&�N�(��ο�\h�"OL��`@ƩJh��+Z����!"O�������>播���� 5�"Oz!�AٲH��mz�Ċ�/Zez�"ODi�.��Z� zt�Ǩ,�F]�&"O�`���Ej!L�S֞!�"O�Q(�E�|l�k�H���q�"O0�H��89��"oыe�b�j"Ox�s�G�l�!B�윢1"O�ـ�ˢe	1�A $�ҹ�F"O|[!J�-��x�N�:g��@�w"O�tKW:y�4�#Ԍb��qF"O��@�h�a�tJ[�i{j�i�"O�`bsi�iN~���jA1a��R"O�ѣ׋�%V2h�'7�0�P"O��[$�$�l����ǂC�x�1�"O��0��'�L��C\}��d�"O��RCFeK��+�(O�=�pD �"O��
����XJ���\�O��r�"O��(��B!1J�:!��5��9+C"OJ�Is���U�Y�^%
��xT"O�Y�"��.K$�=� ���a�%"O�I1�j���1U���h [�"O����AF"I�����,�<��1"OJ��Q�U �aӃ�5]�up�
O��Ps�-x嘠�d\'��l��M��y��@�.E�(W�Z
��Ŗ�~b	�@�`	P��_.��	��A��y��d��&�JI��O�=�@M`��d�|[�]��`��j�"��ӜxQ b�Y�<����"2�6��@m8$でA�?�"���OE�3� ����,B���ct�82߄xI�<� 0���\�F�>�+�G�a����V��C�F��z������%<��Z�dh���4sp����O�>f�ۮ*2B����ړ_���T�.�5'���b?y!E#�^G�$*7�Dn+���\����"��I�?E��eM);��p~ڥ����M�0E1���ȟ�x�l��c�p`+��.��A�sE� ��'}����[�nj��뤡77C��`5WKL�OZ��E�2�)�i�� �V�'�D�m�:nω'+L �&�;��~����31z�4D'�����Ε;	o�Pc���g?�6�O�v��Mp�Z3N�<Q��S��yb���i����6ma��҅�6X�c��p�S�O��6�M�8���6eG�!�l]�eϐP�+�a�Dĉƌ3F.�e3¼ �N3��'.��������DW�2{�]��ȕ�b����%Ʀ�����i�A��x���#�M bΑ)VK@d�	W�+l�0B��Ħ=:�JIHy�h%��	`��(vD�	(E,�	��*�/߀v[��j/O$��Ê�~����->���bHa��1��ɛ&Ԏ��\��p�'n�T3�t�4��&�1�2�2���	J�p}A`*�1�ZP3��i��9QI~��R�'�N=&>%�O��Ի�D@�������10D�(3��1�&gD4j����L��`�\>a��#J ���RwDS�E����+�	7E�����+�lPp@��Y�0�R�
�n� i�>i�F�H�<ad� 0�� ��
�-�[�o�y�<�R��?3^���/��}St��Z�<A4D�� �@���{�$��V�<i�ş��pE��g�2@(�:�K�S�<a�d�)c�`(��އր4��D
M�<��	ƛczd��t�8�G��L�<Q�o_�/��TQ�ER�0!P��J�<aQl�(Q�������U:`���_�<y �H�$L���FI�3�\�8�ɘY�<	��T{�L���Q�,MR� �NX�<� M�/op� �1	`]@�n�<qe�?��ˢ��|�`C�S�<�dCߐ>\|��Y?p��4yÃ�M�<)��ާO4V��`aG6�l	���O�<���"���T�5H����r�<����^]���cN�39\����M^S�<��
�_8����Z�D����	Q�<�'��$�Xu襍P0=��T�M�<A���O}��I�a�v��d��G�<y�EQ+ �02��8J،���y�<���^Ek��QO]�FU4���N�<��
�!)��1��l^1.����D�K�<Y� �
�	�5I]-qL)9a IF�<���`:,$� Hí5d��ka��C�<y��L&0Bt��BO�&pݪ����Q[�<��O��oc�łe��c`��T�U�<�c~G�١�
��Dl
�2dP�<AR��+��)�G�)���$�QN�<a��L�yM^<R�@AT�x��B�<�ES�{���sP�Ŵ������C�<��D�yZ4 X��D�l=�G�}�<q�HK��P�K�L�Lc����	�`�<��E�?=�>�;�!�.Xs!m c�<!G/O�uzU��I�;I�ذ*�L�`�<恍'4�<boй] %�]�<Qv�L^2��4��@��yia��W�<ëN�w$K�&�J�ht��ϑ}�<��-ˉ sB �7@��AF��SG��{�<�F� ��)jf��"�RKN_�<DM�}Ҡ$#���m�Y��`_�<� ݷN7�L�עDP�NI! ��X�<�ǥ�!Mp���"Xw��R�Q�<yV�*t
V!
2�	�DIYT�L�<As^2c�j��SF@�F~�L+��R�<� �X#`f��$�18�l�)5Y&d�"Oh�`�"�5?j�Ȓ+�L���ic"ON��P�Di�Ω��k�D���"O�\���,A9�����z�Z��#"Oj�+�C�~u��ӌbx�S�"O�Y�d���u��)�v��,Y�T�"O�P:�	ܓA�8���Á3M�y�"O��TN�Fq(�M�q�`,�"OP��І@3�8%2��/��-s"O�-(e
����q���9����"O��*� �L��w�M66�0qW"O<�:�i�6`�N�`a�.!�&0�"O�4B��G �X���U>!�"O��FF8�Di�� �(2@�"Ob�'"5���!�VAz���"O�����+�$#E��=/�lh"OTyJ��`��&�Ǣ �P�I"O��"�cH�.	�t�j��W�d�f"Ohdk0X�4�$��q+\�v��L
�"O<XC� Y�z�V�� �JuJs"OH�T瀱=�␘��C
w�Y�"Oxh�I���=�+�tA��h�"O�TS�f��������=(8�"O&1HR&�)�hLZ&�V�&� �"OVH�v�ND��%O!�N$��"O��C� Z�j���+
�1�"Of��3�M�W�E^o ���"OdD�@��k
v�ۑ$��P�(G"O1��î	ԎR�Άs��D��"OZ��kH�N�`��c��l��M�"O�����Հpz��;��؛u"O.4�u��)c�h-�2!QI� "On	(��ʔL\l��PA�$d(��"OصJ�&��V�ܙ�֠K�U��T�v"Oͻ��/81�P��4���"O@\{�*��m������8_�%*%"O �௏�y-�M Ql	$qZh��R"O����F�>X x�6�ן9P~�@$"O�)��٥>���G��?;6X[�"Oʨ�tl,$��I���E4��
�'y�!е��Ou�a�/^�H�P�'���P���fؒ�QE��90>`�
�'�j�A��r�\i*�&��(3
�'����kفMa�S���
�'��Y�&L
�Rɔ�Z���9�Y#	�'���Qw�JR��83���)�b���'���@uhF�*�@­�("��e�'��Q�E��+_]�u{�EU>*�NA*�'���w��/G�ܕ��I�!%>�
�'F�`��CP X�(%�C��<ܻ	�'o��X4��0A֪|qQ ��:|�	�'���V�c� ��:nBq�
�'|8��P�{^~`B���3e�X��'8ʉS��ǖ%"i	_�hp�'l2��%��R�q�BJ�1e>�0�'Ҭi�@<BZʤi%lW�kQZ��	�'�δi��; �&Q����4@P	�'���z��;u�nH���|��}#	�'��|a��?��!��Ł�m4��'����6B5Q�H����w��'�����J�3%� )%�%7��`��'(t�y�	E�n�1��#^�55J���'~�0�s��*�u��Ċ�,|ؤI�'X��TdA�pT�PQ��!��q���� ��k����Pa�4%���"O�%b�I�K K|P�2s"O��1�s�f�D�&9�D��"Ol%�h9Cn�x�Ĭ�x�"Of��G��/�j-��ǌ-�h� "O�}�$"er�ye�˾Ls�@�%"O���C�@\<H2��z�Ru�"Ol2B-@�`��c'M��ҭ87"O���,_7z8��7't$ ��"OXP��A�z �ܰ�EВ8v��
6"O��H��%Бc�qϪ��R"O����ɺ2h��c�)U*B	P�"Obړ�Σ "N�1�\$L���"O0��b<!���V'7`d��"O��i��Q�����l̋n����"O hR�ޒQ���+��+�D��A"OZ����*�v��S�	_x�Л$"O�	cf�P�9�����pw�͒C"O8ը�$b�^� 4��b��kG"O@�C��=@�3H\s�°��"O����h�7!�9�r���"O�=c�GSQS��1�S#+*P�8t"O��q�,�8ZT16i�3xp���"O��z�8L��-�Fh���`�"O��S.Z�< ��H�!јgx�$�"OL�d"��E4\T����}�l!X�"O<#��l��!h����Y�8��a"O��2&����� �S�#�h"O� DMɯ*Q�ч���A���q�"O2�Y�EQ�L(�x���2���"OB 6/Y3~pr�XP���Ǻ��4"O6�������2��@�V`�ȴ��"O: ��V'W%��vA�h��y"O�T�d��n�8�3C I���"O2	"՟{]�����]sی$S�"O�@�ĩ����IrcXo���&"O84Y��ɛ(�ŀ�B����"Of]��!�4O�*����`P<�x"O���݊B�<+��?&�H"O�p!����K��(B� Q�
-�I��"O��AE��
�J����"�`�p"O���
١;8*��@k��6�<�Ѷ"O�m:��ڥm��̉$�T�qy,a*"O����1'�=��A�x]&X�p"O.���Ȇ6��Tq�`)-zp:D"O���f��.^��Q� �;�SG"Oh��ߐE��B�/�'�"�3�"O��I'i�(�M ���LM�q "O�	���\.-F`�aK�F%�"Od�������p���>Cؤa��"Oy0� ר5���'2��`��"O0��N=D�1�b��(��k�"On���%vVq�fۍ� ��"O�����G"���Z�E�5�.+5"O0ps`��=�^8+��7�ص��"O��bT��$���AO%+kEj�"Op@3��vH>�(��_/?����"O�i��#��E���Q�, �E��#2"Oڽ���akȩ�D�A�T\�"O����ĦB������=d�Z�Ç"O�Z�ȍ�A̮��2��S�ƽ��"O�ڲ��2T�J�7}����"O,�)3�E�j&�����|^l�q"O�|$J�<f\�!ɓhdr~�JP"O� ��ע��"p+�gɛW����"O(�	��&����M� #:M�w"O������+�08���ޓX(ۤ"O y�F��f-�Pƛ�pf"���"Od��K9����q"�$0��"OL�D×����Q�AB�&�6�(�"O���1g�Y#D��&[=P.-��"O��R�S��x�"��r2����"O�X�!��U�cO<� )q�"O��
ԟ:Cn��)�(^� 5��"O�	�Ҡ�r��d�凉�\!��"O,�R�L]�f������9�""O.���&Ӧg��蓦@�_;���C"Oą�"�0���U+K���"ON�2��5v����פ�5g#���d"OƤ"�/>Fv�8R�N�uC"O5i5�C�
u.�"�摙{���Ѡ"O,[�#;\̪���%IAȌ
"O�Aء ¼-oʠJ�Fƙ}�ص��"ON���-X�"�X5��$�� �K�"O���W�	D+���4��8p�\E��"Od���"H�{ddlY���C�,�"On��e@���b	ѵ��4�����"O.��D�@�X'"�#C�p�
���"O`5 �.�qnH�-�p#��*D�4�R$6l ]�4�\�YRd�� Ʋ�M���
�KiJ�bE�'DR�'��hg�a�IҟPm8d�`�s�Q�=\6�+a	�	ZT�{p������C��P8���'���*��R/Zd��O�)=^�q�/�%�*��VG��&�����u_@���	  ��rU�F-�,� ǀ�a=�6MB2_��w�`�&�������%��H���C��ٱ"��<B��f�=O�X񑘟�']����Z?��X���|t�p�e�ɦe'�p��4��,O�q�D�ͦ�m��	[���W�K(P���S�XMB98��?9�C��!���?��Ko�s�/:v!��yڴ!'Le�@�H	s��|
A�ΠH����ɏvH�`��وu"��u�ٿV�}*�ڥ|�%`�#2T}Krc�<EO^]�TF�	6�qO(i*#�'>&7�.$Td9"Ӆ��/�tk$�W
`�YJ���	7.P�?�;���{q���6J��#ڐ-�� Pn�0�O��*��3p�ks��8.��۳f;�M{�i�2jh�z���O�Ŧ���}y��O���hr${"��4(�i��I�[f��?��O��gÌ*6J
U8d|����h5I�-��?E�$χrd�౶�R�њ�,�	^�f�K��-h�`V�=����M> ���58Ӳ���U�Kg�Hx6&,n��c���+�OXYoZ��M�����'mڄ��Y"*�\��j�d�Ӷ�d�O ��O�˓�?�ݟ	���*��@��ȑ��Vo����O埠lZn}�D� ""m*���'�b��9,K�(�ւդ!lH���O"�4��hf�O���OD7̀�G<��� �/�|�1��:���s�����O����O<�<Q`��?�2��4f��}�E���+<B�\��(ܡI�,��X>���ZC�)��AO?e�w\�1RDXH��p�@�&A����e�Om��Ms�9�z#}�'R^�@�'��U��L��d� %��O����O���DW;.lj@��*Sdi�4��@Z�"�qO��lZ��M�O>��'�z�4|�d��U"/�^� ����V�F����'c�lr�"�$��'2�'�N����0�Iߦy�1�@�j�����íw<���3��j�AӨW.N���3Lq�i�Ǔ"���3F�­I���S��*?2EQ� R5�[�A���Q*0_���ON����.z>N}�S��A�^��a�i��<���/d��,!�D�Ov��5�"k*q��OA&D�`\�gøc���=�Ş��A�o^����Kٚ9��<�1&C�dzD��4��J6���O2剬xuh��4�?I�AW8)a��i2��V'b�8KN��?����?A��ˈ�?���?a2*����Y��c�d1�GU<"M��MR��a��?lOr횃.��
,�L�!�*%�d���@�>,�Q;�%�dv��;PoK�;+r���5Z-0�؍{��-�?q�i�&Hg��?�b-:��Qhج��t�N���O&��/�d.���ѐL�'�?.��/	ltp�"Ovq����	��x3qD�pM���m�9�M+�i��'�B�'��'ڛ&%j T  �R#�<D��i5�K�ss�0Y�UH��5
�6D�d�H�̀@`�ѕ/F�Q��!D�H`	S�_C�qrIՁ<ad��o D���v�1\��Ȩv
W�pe`}ɷ�>D���ïȁxi ���(W������0D���"�ܵaJLF���|hc� D�H	$��L!h�$�Y���s�>D�L*���"b�Z���.i<E1=D�+�/��\C��ݎ� C-7D��	��̳?r��%h��6�Tl��b4T��X�/ X��q� �{�Z�"O�TǭC#b������<�%��"O��1A��W�|���B�ര�"O��ņM!p7�R� ��)+��2u"O��
f�3�$��F��+I����"OJ@�c_�ka�PZ��כG/<(z�"O��Y���;�������D�s"O:����H+~`�ck�V����s"O�����DD��L��,�<�(��s"O�s $�*P
(|QVL�$?Všs"O�uZ#�{��IP�VRD( 4�*D�09��ѽD�6	5�S�#�<tIU''D�(��_�X"ܤ���V>1tB��(D�� �5�&��Y�|�')�@�:�*�"O��Pc����V)/*��xB�"O���)��j��W̴<�y��"OR�����-= s7�P!>)���t"Of������	Ȇ0������,�"O��U៖IԝJ%G+6��`�u"O��$G�$v���"hՕ{���3�"Ol�������ae�!d�,;A"O��3BD�=>�5A�Eٗ*wnu�F"O�a��.��mP�b7���tɀ�Ru"O�X��%T�T�1*�c�y�8�*�"OH]{����\�2�I�]���*�"O�h�dhū>��+`��e�2�+e"OB��#W1o@���>��E:"Oz�{P��U�0Ex�'�10FF�"O�e��dQ�%���8�/qZ�m�T�֦����8a�����?���?1��j�d�O06-  G�6�2P�Q&}2X]5���f�74�XQ۴؅f��D����#3IH1qp�4�X4^��c�m52�X �ˈ�B�B��纃 ��?�(O�L��H�a�@ �r�$J�,���i	!�R��+��O��$<�D��DP�*�.F	-���̀#}�x�DW���>�C���t��̚���?�3���<Ph7�>�ċǦU��ny�	�h,6�s�T�0�m�첑쐜 �d!zDM�ß����X�T����ן�cj�?{�>UW˛٦Y���k�*4r���F�H���=lO(��Ѳly �a�]��X��<x�	��ő=v�r��bgE��t��И 5�a��{B(L��?�d�i�N�ɓ�[:?��i�q�
�n�SF��q���O��ʣ*�i���Oc0	JE�M�R��!hY �͈�'�a���. &��O, �Xa����Q �4x��V�'K�6-J0� n�����'�D��B�%�\�=#�E��h�8:&���>��q{��c���Ф��`��}Pt��8{&<��n���Q�S�Al�����%!�
c�d:N̨qDR-�DȆ|��	8B�> �F���u��iR��1���P)x����E�_E`y�I$�M��i<��T��(�� *A��$8J�a���n��	ß���Ly������ᔠ\�@l1P��@�P'ni��x���M��O��� �*!�2�H�j�5HB(L2%JD�r&П��	ӟ�ӊe	=�	ß���Ȧ�FI�iJP�VhY.M_�U!����)�*�>���R����4�(OzYSaƍp��9b+���X3@�3YF�L���g�)��݂%<"p#%��!��ݥ����;^O��[��R�w�&X���o�����':>7�����o�>�h��*�
�L�&)x,�؊��'���'�a{�#�oˊ+�r�[��V���'Tv6mV���&� ���?�lZ+Pq>I��:0�d	3��8��#�`�t��3�?���?��?����O4�$t��r#�;�f�x���9ň݊�G����Q�i��Q:nZ�l��x2.2tzZ��P��?�J�p�� ��-:���155�x� 	W�D�S3�I0o��z�CI 2�`	c��(n7�ֹA%B"}Ө�%�\�	П�$�DҠb�/wD�䙯A���`ū��|G{���Z��R�g��V�Ĺ�7�K)cW��r�N-)P��| Ӗ�	�<ٗi[�'�6�i�-b0@*3?� +L�z!h9�T��O���O
]���Od�D�O�a-��]a��ʟ'+Xi��S�"��R�"ȷ?�fi�pƞ�`�Aބ
�`�΄�)K��\��F��#aZ�qm�l���:M��"
�	`@���O��o�<M{�a�v��/oJ� ���0)HB�C��>A��?1M>a��T�۴��C�+��B�b@��y�gO�p�0��pÀ�@fđ6f��mZ��M�J>y��?�H>��4.5��� @�?�~\m�ϟ�O_��zrJ�,(� �B�$C�@�Y�e�O2�$�O�S��?C.�Lܖ�UB��j�k�l���զM�޴�MCe+ٻ�����WUNZY C&�E?��C!C��f�'�B_>��П������Is)N<�����〖j�����<�<��ՓFS̸�ݴT��7-�|�.�,��LI���E×>bnu	�*��B�Mn�50r�Y�E�6���QV��s�Q?7P K�|e� �1&��R�+b^�V	���?A��i����?�E�ܴCĲY`S6*�ᱡL	bC���	t���HOJqs�����	��F�;j���bB�$�Oj�n��M�J>a���uG�W%I�2��DY�J�P��kX���?�wg�+iaX)����?����?����D�TH����j�4�A��n���˲D�ğ(�c�F�,��$�E�'@!�?'�p�p ���s���!$XvQl5��+�5��=ʷO6��ɗ�mK������"���>��7-��w �`��fB ��	�h	&�Lڦ�AN<����?q�O�m��dJbm�`!�%kO����O�����k�XY�E�M6�B�Y�"�.�A�4k��f�|�O��|�i�8 � ��b����K���1���1��-2�(C�1c�Ԉ�JțH�v����@�8�vp���G�
������V��Ov�<�o�͟�$>���B5�!7cW#_-�q  � �?������O>�=���80�Dr!�z"(O�eN^E��I	�M3��i[���\e�$#�nA�i���x1Nלhc�)(	J>Eᛶ�'�2���� ��'���i��p��ץh�\�b#��AH�!�N��6	��Uiy�V��4|O���o���3}�J�!�����!�ּ�U4�F��.�_�@P3���mB%i(�g}r
��"$����T	2e��,�@�ĕ���,O
h9���O����Nt�c&I�Z��5RT����d(��L��
�K�C���(M�(�p5��b��?�v�iY7/�$���g�䵱uiٚ!v�k��@���bfC˟Xi�`�=�d���4��џ�+_w���'l��.Ӻi��Epf��F�Z�"G�W:D�0���/wK��	�2��X����I��T�D�C��#��_�l��A�)Cq��SF�]�[��M��֤T�>�G8��J���Ķ4z5憓������?�"�i��O����O\O�A!m
�:|]��	غl�#&mH<�� }�q�R��䅱��Y�a?*6�.�R̦���O����Z�1� �  ��˃>�"T;u�U~����O�H'״�rt�sÝ$��Î�鈹p�`�_�w�l�ygNAV��+I�����C`�~���A]�T!t�4�ޣP� |JVhW�������?�}��B쀓QAھ<�j�eE��(O����֦�i޴���uwa�!`��d��!Җ5h&��u�ʡ,���O��ĕ8WZE����OX�$�O|�$ɣ�yW�l�b��(֫�r�і��~�'��]Q�d�>zv�Ѕ�ɏ"�!p�(�O��P�6�ĩ:sx�hQ�w���n4i��
!$S�i҇X� Ve�ڼ���O-B��L���f��kT,]�l˓<v�IY���?I��?)�4l�N��(�'4�¹�Hz1�ɧOb��DG� �(h0�K�B��u��A���C��:�4�����'�ē<�ơ[��Ƞ��LdԴ��O���   �ǔk��USc�?|�nL*F�|�B}�"!
a�6�r�+�bqn��$�a�T�#��O�xnZ#�,��MH"���"���13�he�ßd�'2���Op�d`�<d6'U<$����rD.$��CuH<i�cSJQ�
��6V� �S é� =�Ey�������������O.ʧNȩQ��Y�*I��f�ܜ[�џ�?���?�f�� 4^� S��Iw����Zi�4�C}r1 t�ʦ{5 ��$|i�xh�E�%�5	���#��<X�gFon�c"n��o��<�����'z�Iz�qP�vOc�8��:��>NN:�	"h1*��E�=O�,����L�'���Y�ؙg�]"?���d�G��}3��5\O"�n�
�M��O ��lMx�j"�X&<�,�+��%ضl��4�?��?ͧpn�$P��?���M+��v��$�,$���O�hւ�i�͸w7�cIɦ�ѡӟX˧B�l�����<)��d��b��j�P"�tĻ�CI$���#4D�X��aD��O���CA�$	�da��[-��a��\؟H+ٴ@F�ɻw�#|���-0P�[�BD��0�f	-H��H!���۟��?���O%��	���xִ�c��h�PXO�p�I��M��iF�'����O �f;/�� ���p���̂#A�"��L;q8x���OD��O��$�����?��4
�M��l
D�]R�Bס,�M��i�>�l�)�~��z��X��d�B�g��Ќ�4Oҭ��"���.J���;z���]T��d��͊CQ�'&xպ%�H�>�ư��NȾ2qf�0�4[�D0�ɦ�MS1�x2�'��x�P��n��Q������c�t��C�I]�H�(�FL=,p�I	��ˎ#��uу�i��'}�6m����O���wkTU� @ ����=V侸�	��L���iglJFL�39+&�I�._�h��c%��s�2g�'�Ԡ�WiԽ+�qZs哂f9���b�A�m���p웣2>a��>>���K���5�Z��=YuoFß��i�pДhZ�͕s	����'�o&pII<Q���?�H>qI|C�ȝ7$0CSO?�$��3��U�<Y@)Ҏ����dY>�~|���QI?q�i��79��O�d1��E� �  ��(1ge�"f:<8�"O�@��ۚG��H��݀J%�l0#"O! �霏ؚEȂ��
�� �u"O���q/��'*؈�� "�>X1R"O�E�T)� l��Y�i�7"nI
A"O��r�Q�vyI�G\	"��a��"O>���$��1%O�G����"OVd�"pE�$y�$�0��*�"On:���}��� ��p�"O��#� 1S/B��M����"O���L�>R��Cp+_/El];�"OE� -��/ʰIY1��j>�D��"ON���D�"X�gF# |S�"Oh!	�.�+g���Տ�"?�d�"OtIrB%��T�	�P�]����"O� ��?l���M�:�4�1"O��IC÷&�6L1&P7*�"�x#"O\J�M8#d���n��)H�"OС� �W(;I�q"��m^��2"O(L����N���A�,<��`�"O��
D �5�`�
ƻx�|��"O�U��C$1ƴȐ��ԉL����"O�d8^ɶXceǅv!F�1�"O@MA�N���E�%-�*q�:���"OzEr1�B�����k�6�J@t"O\�a�oN2M�p�I�(�*-V�s`"OLATh��9� �p手USq��"O��r&$Q�Z^���O�*����"OXH�B�G.H8"t�U��	J�"O�e�`��'p�Ҍ^�]�d�:�y���
�^�i��Ό��&�Z0�y���]�` k�-3|L�!Eጰ�y
� ���*T_�. �%ڐ'����"O�$���x)p�&d!$� z�"O���+�w�����Z3C�:'"O�T�f���}�8P��X�F|�"O�)	�4t���$�14m��*�"O��J׀O.�m3�m ZVLiy�"O��dA�2��(`p.ٌLGL��#"O�kg��^܍�0(�7H�J�س"OU�&�=2�f��?(c�R"O�=Z��N7Eq� [��Pc�@Ș�"O��r�*֑REכ��@�"OnY����v���R�Ƀ-%Tx���"O��x��܋ U|:5���`;v���"OZ�#�P���C�B,`��W"O�Ip��зnl�1��8v�Bt"Oq���� @k�c��O-m��� w"O��Ab-=&r�D��dI�E�e �"Oae��T��r��S� ��5"OHláBT:T
4���A�])�d"OL�0��ٜ�1Q�H<P�>�"O~&ɎS���PD�0H��p"O���t�[�$�C�!7qh,h�"O�8 !�ȿd�<,ҡ���/va�"O̔�1���Ԑ�G�'*_ ��5"OHuC��U�xFL=a��(Hp �"O.�	�.�������% .9؊�"O\�2��ۿ\4[ʏ�a��dA"Ox��L|)�	��g�|qz@��"O��2��2:��gQpx�'"O���0
��1��զB��Ur�"OVL��K��5Dڸ�b<#����0"O��!@72�W!_�x��e��"O�[��µ/46ÅT,xC!�<t!D�
��\�;���R�R!�d�?&=�xg�
�j��j��Q�F:!�D3J@�Z`���HC�����(!�ǟbW�E:���:8=�E��3|�!��o��c��]<.5D1��m�Z��$���ѣ���ZFI���y2ݵ7�&�J���A�%hC8�y�#ţ1�P�p�ɗ:���4D[��yM�����5��!/M��$FO�yrF�X� �R$��4��6�yr��x��!bS`��E�pA�#���y�]�YY���Ӎ�)=�:�3���yN�<n<.!&�+�Vm�3���yAч� ,a�*�8��y�b�Y=�y�-d/4c3H]�^�tXYB��
�y���z�������>]�8("Y��y�d@5l��2�6&9#B ȳ�y��̲:�L��ʊLi��C�:�yriʵQ��GNBlƨ�@�H��y��S"Z���ԃ;	J���@Z��yb�_�]1|P"��	�����	 �y�A�:\��_4�J��mT�yҏ�:nJ��b��e���J���y����X�z	94��%l��{e���y���L���X&�(Oda�'f�y�@U-�eɑh��E $��9�y2
�Z���0�-X�E����y2JM�D�9����u�@=ҥMҩ�y���m��X�S��j訽r����y­U�f�� N�f��X�T%��yR��KƐ��=)Ťɲ�W��y
� \2��ջ@��Y�ā�iF�*�"O���eԯSA��r��܅F`�̓"O�|
���;DO�1"����$OF|;�"O4<�eE[�e^���>4n�	3"On��t���j%>�2�	V��%�"O�)�sa�xX�����\���kv"O�dpBG�n���#�!sa�"O8�'��%}V��!���2`��Ѡ�"OpY�$���tM�Q&���B}13"O6(��T�y�l�[wn��zAư��"Oz�bЂ k���`��Z5rA�P�"O��k��׊lpZe懼lY��i�"O��1Ҏ�(C�yQ���'?�[g"O.%�wD�a�p��S�.:.z@�"ON|Ȥkb��{т�#B�a"O�ό
k�J�r���j��U"O�5��t����Ã^8q�"O(�"���)M�,��W?A���"O���wB��?�l�ˑ�:A�%{0"OP|『�oW�@_�R��"O����NS�K �I�C�Hlj��"OڤyR!O�6��'�, k�%�"O���H��j*��U��"O(���"O8�,mr�(.�8T�����%�y��7)�XJ�����Ba�F	G��y�J&(_,A��ŋZ����%����yB��Z�4���N�K�1 �6�y�nӗ!J8��m�3DQL-�W��y�*R�I����$�'�iÛ��y"����Z�(W:�%�1�I��yʡ`�����r�;a��y"�ۉzT����@�C�*�']��yB҆e8 ��旳$�!5�y��2|�(QcM�1�Lq��0�y2�)Sp�kR�</X\Q�'X�y���l�"D	q�7'Ί�:�"���y��Q�5$_�rg�xr��܇�y���nH�FF\(o���C����y��A 򢜚�Od��P�3��y2*ܧ
]��D�W�Z?�5�����yb@�������X�VB5�Y5�yr�<�q���g�p�cM���y��IU~��;`gY�a=t)�c���yrO�,m��ɓrg�"y�1'L���y@��h�_�1� A��N4�y2� �2��x��JI%)�̠u.�7�y�T��)���A�3{�}�$���yB%�z6��K��5���9�J��y�G�$��
_�`u���sNR
�yB�^+;�-Rt�0/�\�Ӓ�k��'Y���T,�_�T4�b�W:+ ��{	�'8��c�R���Q��(�����''�`���-c�j���C> G���'a�jp���f�x�<B6��1�'3H�8 Kƫp�|�G,�9�<S�'��MI�E����\k�H*�J$��'Hj���L��q	0�Q��)��y)�'�YB$قZ�pi'��D��'��I�E-߶?�-;&�& vT#�'Af���$�
{'�]╠Q	 �� �'z~}�6̛�&+Ϗs��	��Έ^�<�F�U�V��-�DG��jj �z�*	s�<�7�'Z�HqpI�"r���C�A�U�<Y�N�U"L�"A�	*��01�EH�<� "-#jKT("��o1
�av"OΝ�=7F~p2�T#��K�"O�����܁d��|��ƈU(C"O�lɱE�/6�.�#ԇ3e"%�"O����,,�*�����;���8�"O^�C��8 A��� �*t"O�8�q�Y�I!���!	Y�p� �r�"O�tȁ*S�q~���h��\.J�F"O$ �  ��`6vY���*�DIP"O����M�L%�J�=X<��"OԐ���J-W/h`q�"ȝ����"O� �ƀ��N�X��� M6'��� �"O>���� ��E�`��	(Rf"O4@�����Zt�
�Zը�Z "O ���D1��j7gCE,45�0"Ovݑ�C�]0��ehԙH�9��"OdtcՄ��J�±1pF;P-$E�"O�Lڠ��0����$l��"O�0�R,D�U`|��7��g��=�"O�E �O�*!����G_;y�9�"O8<x��ޤpaU`̉U�I�V"O��T-� X�ɋp!��n��"O��S4��Tr�ţE�n=�|�"O0�k��6�`��0̾mܞ\R�"O�t�4o]6�\qfŷNش��"O�D�oJ��8�B�Τ��"O��mcѸu���I��~���,_c�<��A�?G�j	��)WWh�:5�Xg�<!�˳B���i@ҕ2 ��c�<!�I�;Tz`���O u{��y3�G_�<��iC�Ͼ=�&E��!YG�^�<!b	27o�U�@������s�@^�<��+�v����`��v�HNe�<���]��\h��L�x�[W��G�<qVj��B���˒*�!b>L�Ŋ�\�<1�
]��,��S�4@6���,�m�<i��I1N�D�"���n\h��S�<	&��Lޞ�c�xx���z�<�h̵'[Q���I��F���Lb�<�	�J���\�BU(�
A�V�<��%OC�����U2��7d�F�<A�+k�H9T�m�UP��D�<qª�;k�8�����Ft6X��D�<i���F��6`�$
`��_A�<�S��_-�=*�o�'�\yp��t�<1f���A�{� �/?�0H�� Kq�<A"�YwL�I��̮g,�P��fIV�<�UB�?q��yɰ��2	��&�Zi�<�#Iw
X��W�=�:��r��f�<.��z�H�[0֦El��vL�a�<Q��ڤ.��P����7&J��W��Y�<!TJL�e� ��c�X�9�L�G�W�<�g��TÄ�
���D�K�<!G��aY<�)�,рeS�Ͱ��M�<Q���<k�L�k�H��l�
��AL�<1�V:�.O�:WT͓3�J�<Q�&�*� "�L��>�d�Q��E�<I�Yuv��k�&<�&S��EG�<���������ƺE�(��"��M�<9 G%~���aƐnΪ��d��M�<q��ɍ=���knAnݰ�H�<R���={|ppń�rZ��x,�B�<1��I�L<p4|
ؕ@��A�<�d�$f��c��_�<)p�f�<� 2�RD �I���C�^�Ԅ��"O�y1%����E юԋa�n��"O��`Q��4�!���	/�	9F"OV��f�� ��i���:Q H�e"O�)!���+|VɛRg
�=	���"OP!3BF�&B�@1f�;���Bb"O (�Ʉx	ö���n�J�x"O�(p�A�H��q�N�ry�q"O\���%��#`)�!�ؐ�"O2���+ �uY�ؘ�0���"OR�UG&w�$��$?�8d��"O�D����q=
�N��pSP�"O�0���~4��Ƀ��6x9�=��"O���%E6R��`����@!����"Ol�sq�]�Q�*��M�*P�""O|%1����<��1���^���rs"O:Xk�d]3`�
���¨%����"Oz�cᓹƅ�.�[FI���!�ڮ�������S<Bp@��0!��"Q2E�AT�u/ne�B�9t!�'/.�p��ںj��Ч焾Br!��Ԁ|Hm��
6:��U����/hH!��@�U듪��}k��3��	�W!��^��m��l^]Ă$:b�1>;!�d��|Q��X�A���@*�6.!�/ ���U�w�u����~!�B�9W��at��4os@��ȇ$�!�$��f a��5qr|!F���(�!��P����u$�Z����W�s�!�0��!�">@M�I�8��� "OP	K�N�Cm�l� �.�("O ����3vf���s��~���cw"O�T�E!:�}0vƀzn��b�"O֬˴`:(�Ƞ��?A<Hء"O��S�Ew$|�x��ǉ�J��"OҬK0	̞i�|E!���Rа ��"O8|�b��<0����ʹim��k�"O�}����r���e��	 �×"O�Y�����mSJ֗KK�|1p"O�)*�h�'��(1
E�rANթ�"Oh��r�>�r-0g�!a�0m"O,��CN�Kk�	�D/�<G{����"O������2�$4 H�N}xp�"O�Yu�C�~F�C�Q�Cfr	��"O\�q�G�!\��g��)`
�Ѡ"Oȱ���؇c��	'��r}j��""O&��lA�^�� 1� 	�w�Jt"O��I��E  �n����6F�
s"OBD�!]tXhѫqOֈO�@�(!"O��r�!��@��#���@�"O��A�o�I<�1�t��l����"O���Ǥ��P�\i0��s��ixc"O��R��eH����AZ�@H�"O֕�P	��V��Cp���=ӂ�I�"O֥��<O�T	�'C�omP�!�"O��vʙ�Vo��zw���kb�#�"O��#��0c�6qH'�̢u]��$"O�q��@�-Z��T(�[�Qj�5"O��Aw�E�s�􄉈
G�(��"O�Y�f��NZ���E^�b���"O� �;!�h��pD�62`�W"O�҄��TIF1�5�ɯ/��Л�"OZ��F�x %��B�;'�00��"O�0�����6n��27_��up "O� .�ʅk��\�.�Rg�G��z�s�"O�`҃�&]#q�{���R"O�	#��C,��j#M�[g|��U"O�=��8�jp�G�)�2|�q"O��cbk�'C�N���\�4�`(qs"OLu	��تe�v,S��H��d��"O� 3���?~B�Z!�#Jx�u�%"O,���h.,��d�ͯ`¬��"O���V��>�	�Nи9F��@"O�X����)�涬Bq"O|pK��Q� &��6� ͜�b`"O5+�ިNsl��gV��<�v"Onȉ�BZ2��d#��J��ԋ�"O��c��&V���J�+s� t[�"O>���+� /�
i`G.gF�e�t"OJQ�$/M7\��Ź�M)��a�"O�|�uNN������@�Z����"O����y�d��.P{Y�t@�"O�Q(�c�R�p����(^���"O�4Ύ�kK�} �lߡD;��{"O�<P���\�M��,��G6*D�B"Oz10/W�s��M��jZ�{�hbu"O(p�t�I�Pِlx���D�b0�c"O�ha��9h,��PW%Ei��aqR"O�� �� E�V�i�Dه�=�"O�A@k�jG��{ 
X1����s"O�L�B�l���PD�*x
�"O<��đ+9?z�k�f�3/#���"O|(I���R�L���J�)>1�b"O���҉�2A��IK��q4"O�	��N��k(�7f3h�p"O$c!j�$t���J	 ���r�"O�����ސ1��A[2"޾<z����"OM�1�;�m�疇UM>�ٖ"O�\8 �ۏ;����S�Ӳ\F�j�"OJC#�%&�>���& y!��b"OP���_2.I �[%A2]��"Op�Y��8�����պ10�(�2"O��z�e��/@b��5$ׁ-�-��"OJ%��bO	{�D�Ʉ�!��"O�YXtl�:Usz��Bh��* V�x�"O��0M�1�^�`E04-�p2�"O��
��@hjd%	E���ap"O�i7��(�d��ǣ�7��;"O����E �I��L��嘽Q��W"O��zBe�������MP�ARLc�"O�4�$�P�V:�T�W��?^+r���"O.yM���BW,�Z
D#"O0`1��G-��(cJ��G �ٓ"Oq"��؄����)Ӷ"Opq�b�%Y�*�ԁ��D�y�"O~0��8 ��D`M\���y"O�T�bS5s8�[�,�z�x3"O�Ay4��7f�����hR�+�"O&�3�W	Z�8=Зe�'^@.D��"O�ٺ�!��*@���	L1^7��Y�"O"\I��&Q��!��b��|�"O�Q(��͕c¸I#�bMSlLl��"OBX��j�?^�D��A�L^R��"O��:���R`*��Á%C�D!	"O:4�lΚD�5p�G
$� c"ODa��S48��X�J���"O�D�!���F�P;�fǈ|TL<��"Of��q�K�%l&��&��-?\ �"O� ��¢M'����'v-��*"O>��f/P\z,�!�F�<VM;�"Op�c�Vs��'(���"Ot���:.DAР��<[&�D�6"O��Jo��f;n	ƀ�!ԣt"O``����&d�n�FM�2Y�-	�"O�&�Zp�:��Yڐ�""OH@cb(C�x���{�T*a�4c�"OVD ��4�&|b�g����*�"O* �Q"A�����DF�����"O0 ڠ�S����Ӆ K�����"O�a��%&GNd(��A��8�#�"OZ��K3B�N�u�M�F�"T1s"O�e)mA���0A��O5=��(q"O����#5-��HP�]ʼ��"O�5"!�3<���PcȾ*dT�"�"OBq2����#!"rŤ��gO:L��"O �;�&*�͕ۗ7HPX�"O�qcT���L�w�-�|�	�"O6����.��qw�ũ+2N`��"O&��&O��Wg��z4�e��L;1"O�3&�K�< rl� [��q�"O<����=F5��Y&j���)('"O\H����16��,��I���b�i�"OL�RE<�Es"Ո�q�"O8�0�̒	�:���fJ�g$���"OD�D�� ���`7�O�贄��"O`���7U޾�q�a��R��"O�P���l]*������"Oڵ����<�\�&kK%Y��,y"OR\��lR-lZ>Q����{�ni�3"O~�ňG�T��<qR	M S�4�r"O�< �	�3a#"����:x� �u"O��gEG�l1$]�qGX�g�D�"OnS�ꊌ�.D�R�G�SN��[Q"O������NE��E�<s5D�`�"O�H�f��O�,�dR>�,�@"O�őЄ�[ohT�f$��u�i�"O%B�'D�T�xU%i*�!�"OXX8�#N�TO��Pg�&/zP�"OB��	�m���c��ޯJ#�yP�"O0D�J��4�ލ�'C�2���"O�Գ�Ù�[�,Pb��4��tB$"O�qRk�-���(��f�6���"O���E�ӷ+�����D8�2"O^q�Uǐ?(��Y��  3��ۓ"O! �e�
P�t�pq˕<�Y�"OHy��W�X�L�"T	U-G�b��"O$�ꕩϧ(�F���=�4<i"O���C���aE����'�'( (aT"ONx�E��k}~� �h\�(�l�"O��%�}�u�2hT�u>��d"OZ)��\�F	T�K�E�.$ˇ"O.�BР�6*�Ό�G�h`�q"O�l)%�K8T����qB ]�E"O�"�Ɯ.)E>� A���̩�"O2��M�<6q��Ž%b(���"O���t�g��8@�m�u{,\��"O@���
ٯ1��X�,��%n|,�"O��g��8��C�;oW]�C"O&�3f��*Vm�У�1DZ�w"O)���2-�֩�T�¬@��%�d"OJ�Jc��"W� �ʖ�j,�u�w"O�]���ĺ]��=�@�BGу"O� $u��B<O��x��V0").��c"O�E[�J9P���N�<"� �"OV�1ӆ��a��JW@��YPm�3"O�ՙg�Mg�@1��#+� �"O`X1��<Tu$�:f!��'�Ly��"O��8V�M2Y��y�T��G�p�z"O.L�v�ԏװИp�
4�p��"O��$ Hɢp��^�*��iyc"O"�8i��B�� �/�=Vk��Q�'��%��#�1ŖZvb��-�q��'|J����zΨ�@���)޾���'���2 �ܬp��9�E�Ͱ)s��J�'�4���׈t�ɉE�ߺ 3D���'/dq25D��^�$G�AWB@��'b���SCY�X��px���/)����',��#���^�R��#!9*T�'��}Z��P�/��� *�67�̨��'������u�Q�c��29�����'���B���<,ƌ���g�2=(�{�'�쐸� E$R�x�kcb�#lĳ	�'��d9���=&��<)�.ػ"�d	�'F4tƧ�iM����"�,���'��9�G�
�"�����ڜ��Ɂ	�'=����*�$T$^�����|`���'>BI�V٭]8T��%��z����'l=0�mۛu]
��a�HkH�K�'+�MA0�8e�0��Ti����'�^:L:�,�H��)`H蔨	�'�T᠍�o�Aa&�]��r	�':�i��!�,n.�D�PG�]�����'-�I2S��5�~���&M�2A�
�'��ifeY�Q�$�qGF1O-�IB
�'r��f��t,ڜ��_*^�4
�'����Ʋ$V�����
Vd��	�'ǲ����/ZJ��SP>(ك	�' �D0�Έ~�TXOS?��!�'Э+U���1RF	emf�P�'I�"m�=1��5�@C�S��@��'�lCƃYX�� ��������'F���W)�-e-���d(�BB�"�'ݪܡw�1������^�E �4��'IR�bph�G� i�/·iZZ<��'3
�1Ɔ8R��2��0L\X�'��i���@N���rP��8'�v��
�'�>��
P�g@�����<,c ���'+�}�w��Y�4pSnY� Sr�
�'"��d��!�y����C��j	�'��[F�K0.�z`9�i��=	���'b���
��L�Z�pF��3g �	�'H��� g�[��9C&@B�7i��'�v�q��Z�a�8�eH��`����'/BQÖ�P ���eF:)� k�'����䃇��1��M:OT,k�'~f0�L�iXz���kL�L����'X�	��^9j"�`��l�w� ��'�d& 
O���i!�+n��<y�'pb�Y��ϱ.@�Y� 
5P�~4��'펀��&<�:�;�LŘG���'�a��kܺ��C�C��1[�H�'yV4�򨌄7<����=F)��'�d1��H�u�lmsd� Bw���',<�Y�甩{$�"�JR,3O�Ez�'*yz�M8s*��z�)\�#QhK�'��T)-�<7XEрE� |��
��� �U�K�k����D+Ա=5��D"O� ��2�<l�p��-(i��"O�0b�F�-r`IR�j \�BA"O����e�H��h��Ȟ�^��� "OՈW�2O�����V�"�!�"O �j$%	!qȜjU���r
e�"O��C���P ��ǉ�@dʝ#U"O�3��ȓ�F���Qb�3�"O��*��?jĵKa�lB���q"Oz��H�f8R��cA]7��Q"O��xB��qB>�:���$'�(P��"OBĂv�+	�ԭs��O6c�t+�"O 5,L�(D��b�m[�]w���"O��!g�^�i�X��4lcZ@��Q"O��2�΀D�Mb+ݱ`+��`"O]p�IY&!�u�T�S�U(T�v"O\�� � O.`���,,���E"O|qرg����	((�@"O��"�aA�e7����W�
�*Ҥ�y�n�I�����C"���%�y��ެr�L��`H�5񄔻W����y"F�wt4q���<'h�uK����y�+��"
d�r3�:b�)"#��y��=o6��g.�Te
rh'�yB�R�V��A�||�Ôm7�y����̴`���L��ah4���y�$��I�d�0��4&�D�s���yr�!=��:@o�Z�b��	�yr�ѝ<�u��� 8���/�y�e�_oa����Z��3$� �y�'E@���T%�	��p3��
�yBlY�	�D)����y�����ǲ�y�ǜ`�(�$��wo��ӑh�9�yrꋖI%&!j��3AN���!Z�yR&�;-p,X�N�=����ۊ�Py�0vmK�LRF��L� ��f�<��	�w$8�z�m��Bxa�Ad�<�6�W��H�ir ��(��p�b�F�<!��E ��i!�ˑ�NL9����L�<� UO��I9��ӂvd��a�[m�<�S��)G�԰ٕ��;�B�3rB@k�<Ip]�
Β4�cKA3+�V�� �m�<�g����0��.yvz�)Q�^N�<3�\���0��VKN�9"�M�<!F��P����Ε4�Z�)SA�G�<Iu��",��K��l�j��cE��<�׀D���91�^�4�s`�C�<�dmĶ!H<��M� wф22|�<Y�BȅE����&'Ð_�M�W�B{�<�GfүȊL�Bӊ#��`0a�z�<����"~�d`{DK�DȄ�e�y�<�g'6��X�B�3J4Ա��w�<��ҭ@g0��T��Y��	�5��j�<�S,Գ,��-H�E��ݩ`�Wb�<�U��*@=G�	B�e�<IeF7�ͩŌ���i�I[^�<q�I:S�,��� �4���`�*K[�<�N�=f�5�5�[�f�48uj�B�<q����`SLi��Z�W��ː��~�<�d+��j)�"�b�ީ[�H�y�<�S��_vrd���g`Y��
\w�<��� ;��1R�bܛ]�ybV�Ks�<�� �[H���C������F�<�KV>MY`���Ɩ|:���Ō��<� l-#6&��6t�EV�P�<�1"O�m�d_�\X�2d	0s��)�"OЌ���ɔ����ǩhA�"O���Vꅇ}I$�Gc ?B��e�"O&���/�,j�B49V�  C���"O���f+x\i��V�G���"O�Ez��G'n�t��@�W�@�A"O���UJ�R�C�N�eW���F"O�Ȋ5
�8Z����V:E�pJ�"O��K�'U�yX���������e"O�I��6V>|�b�oA� ����"OD��̀����g�#&��E�6"Odl��M�.iHLh�&�	>�h�"On�s"-�#��m�$���1�v$;c"OH��wI�-ֲ�X��ڵ�*l�"OD!`s�W�Y��ٗOˍ�e�"O0���NF6Q����%6�	�"OB�[�����r P��9�М�R"O>d�S*_	z�xH���&5��9"O�����`ʂ�SgdN�>(��"O��&%�e�P���"K+9�X�"O�$�Ž_eܽ�r�ć���:�"O|8��l8 ��Z��Xy�"Ozݑ��@^��o)nkB���"O���n	+w���ƳP���Q"Otb��O�-��C�1}:�)P"O|y�E
]1e�䱑�㗠V��	@�"O��1��J8���b�9cq6��"O40QQ#X�88���N��8z��['"O�DKD	 �C2��)�j<w��`Y0"O���"h�^
��
��FZ��`�"Ot)��N:���J�UR�9(t"O�0�F�Ïm#��s^�*0��"O�{p��p�FD�fA,`t�'"O��#խ�i�H(��.χ֖�J"O&��ck��c���ڗ,uh�"O`�҂� -˚��'\�Z[�a��"O(p�#n]7��2�ZP��E"OĐIUMCS�� �w��
L����"OԹr!��9(&�`��NBL �p��"OJ�G��K��a��5P�EX "O8쁖�ϊ1�L�"ϿHPE�3"O�"�E�%d��Za�̅n��Hc0"Oy�1���t�pȂ%��	1�pŬh�<y��L�a ��R ,,g/���$IE�<iՂ��?c�|J�#)F��Z$�@�<9�)ҽ]��`�Ћ�;Ą�����x�<I�F�77L��F�=-Hθ���M^�<	�ψ;������5^� @��/�Z�<t�Z&>��Ԩ�#�1{p�!QŎk�<��A]�\Ř�M0#�n,�Uhmy�)ʧi�$Q�@5���*t� NL�ȓ.8PсqKO=h�`��@	�*��!��m���A�2��VAFgAvȅ�JB���R�]�_��}�(B<�<(�ȓ����c#��v��H7%r���?���)�C�X���M I)A��9�!��(܊(�%�',�!�&e�6�!��O�z�� �W�\.�٩ e�4-�!�͝y��QRĄ>p��<�Wn_,�!���/�
p�֩ڠ)Z���.��f�!�$ܘ����� o�U�b��H�!�$J6J��Ԑ�O�L��);QΈ�>!�$����a�Uђ5{�/F��!�� L��R	B��%�Z*&�>U��"OLx2E��|���1Ê�gd��T"O�@��\"ڢtA�	�M� �"O�Z��ɀ7�r9��JƬ��	�&�'���8wbu��E\+h���(/��!�$�F����GN�U�j8�N�>(�!�$�o���C,#y�yrw��	�!��ͿSp|�rn�8F�,J�F��v!��ћz�0+6h	?�$�'FT�bg!��+Y@��g W)}+���Q劔$e!�$�*
/x8�3�ߘcBl�3b���UUax�퉇7�DD���J�F\@)B�B޽�<c����I4Y)��sC���>~����ދn�C��($�| �Ԥ��6���8f[%X��B�	?	��%�A�o�
�R�&��B�	1H�L}���4c�H�4��"S��B�ɮS��)9�Dֺ(����#O��vB�I�{�X��
��>���3R��R�H�?��**�'��{�H!0O4��1)Ӓj t$�t�!�'�
Ԫ��J#T�qA���L�\Yr�}r�)��P�~�B�,1Yv�z�Ĉ+8�$Q�
�'>ȩk��	R� 8��`�56 ��:�'LHx�OR;��Y�� �@��1h�%� ��(�6D�8Jf���1T.�H!�
�3�� {����hO?�ă<V���q�*�����ш#�!�DG�.����K	�Y:xTML!�$! ��Ż�N_�k������*F!�Ě�j�RI����G��j���G@!��2�HE�GLS�fQgBw�BB�I	*���)İxY<�X"� *1�C�Iͺ��ĥ:�Dq
f��I��C�Q|����L�q����*��C䉏+p�1X��	�v}c�	P^B�ɕ'&���3��=#\�i����bCZB�	�8 `�xV�PI� ��B��C�0b�������p�J]�TDԚ��C�	�t0b�RVN3'�"���FP��C��!l:�	���Ҍe�E�(��G�C�I?*<�Y5,#Sd1��R̦B�	&(KFmK�޾j���֍�K�NB䉯\JN5¶�B���Y%��
:рC�e 0h��QC����VM�0>�HC�ɤ3�|P�Wi�/�X�B方?����5 ��@#���҉�JѸ`�!�D�w[Z�Y���w��<�@$��!���GJ��umOp���&�Z!�!��2��E��*ն]^Z��qOڲw�!��%	� �BڰQ<�W�L5I�!�D�8*�$�`\por�O�H!���r�,����R=m��83�3�!�d
�nAX��@B޼RqM�!��E�'��,"�����:��;~w!�$�Q+\�aE��j��p�Jk!�$V
@��I*p���X�dtӠ���f�!��5"2\��&#�����+� �!�䃹#8,���'�`���Y��D�=�!�Xc�HYC�#G%|�dCto��V�!��+@X�9�-`p �p��}v!�č�+�P܈�K��xq�h�5�Ӱ0\!�� ��e�ՅJ-{����p(!���o�@�ۣ�No��au��!�d�(��⏋scJȨA�E�dW!�2ZN�*�l�0+�;�(�.r!򤛬h�tQrt����H�`�F�j!�� ,R��m[v�eG�rw�1��"O�e ���8Y�<�v���x7N�2"O���$0��#䉩x��hi#"O���fŔ�#�$� ��)�ƀ��"O\�j0�H�vnX�P�A	:n�ژ+�"O`H��D�f6��灈�PS��j�"O"�G�d����R!���Yk"O$�Q��A�#v�X� ]	M5*���"O�����@v��W���-�4y��"Ot�QfdV9~�2�g�R8o�bE� *O�H8@� �R�lU(��J�=��D�	�'��	aIH�D�S $�3�8uS
�'P�`y�i �)x��p�4�f��	�'ŔEk��_:` ^���%�,汢�'��=+l�>44ȝ���K�up�r
�'�h,2�X;G���Q5�D�m�&p*�'��� ���1;��#���u�̌H�'�bu+�g^�P�n�K#�&[���+�'<�U�w�O4m�",W�<M��'��IuH���h8H5�"0��!��'~�@J���,M 1Q�!��x���'.PEj!+K�ra:У#�M���'�����B5`�z}0�$\)q��X�'���"-X�fqz��%Ex�����'�5:a,�h�	���yI΅�'�\���G��B����`�!f��@�
�'Z�h5i�v
�H��+X��Q�'
r��b�P���]�0�"J���	�'��ݢ�A.;��8+`N�;�&i��'Ѱ���Z<��ՌY$]����'ѨȱAдUi��ߑb:��
�'���s���8��.iԑ�	�'z�rG�T,]ҨC��d�c�' ���«ٷ7Mh�""Z�X��'���[%YF|� CL�Qn�8�'Y��N��Eqa(�2+Rqh�'����n -��q�����`q
�'5z1��.��� � &��|�	�'>i�uf ��M٠�
0ā��'�����$)�p��n��1�'��HW*	�O� ��(�Yp�'�`�a���g�,� �-u��\*�'�%���"{���
*t0L��':.�����O���8��2|�V\��'������I�d��C��@lթ�'a��׏I� �����n�U��'�FjU-C-P��;!�V_G�p!�'� ���H2 BJ�
�DY+�'L�퓦�e���1r=��'^:@�ŋ�k�	�U�[�b�H[�'$�4	B Z�|� ��yO�H�	�'��Y`��+g�������X�'���R�+��Q.6,٠K��RlIJ�';& �ϖ*
�`80�H,�	z�'�H #������WF��{Z���'��ٲc�P13��As�Ꜵ|!��S�'�`foĎ���`�iz��i�'p�#'
�{�P��߸^=���'�8��@*U���,d��T�T��J5"�&� �\��!d\#]�`Y�ȓ%N �����` �@̾U-}*��-D�T(fAĦX7�mb���G>8J$.-D�(�p�ܿW[�i�AU#-U�����.D�IC�T,N��-{���99� -)0a,D�� &e�ehT�N�\���m�y{����"O�q�-��8"�5h��[�"O`1j#���6�T$x���@Q�	�"O�����ڼ��A�d8�H�P"O4�9fM�
`x�0��	^�ca"O*����(N����f�T�>�2�[u"O~�8�FN�I=2���Ƀ�B�A��"O���&�!�
�SFi��#�8�)�"O�����E�����D5s��c�:OF��ꜮXVVhK�H\�Q���U�	�8�di�,jq�@eML	�VC�	�^�Y�=oT�F*��;w(C��fI y��
�#6�
W�ܠY��B䉮Vc4]�`^�b�8\�� Z�(=B��(�4�@�T6�^���_�t��C�ɡXK��т(M����eݺeO�C�I&=���z��ݭ9!(��a�T�"��C�I _Oؑ��G��h{�~�BB��Vp
��I Ø\q�/�3~^B�&`�,���S��!IA��m?B�	�R�D�Hbe[�$�vEp��X��C�	<�iqb��2���&D���fB�	�|6� �B�4�%�?O�NDJ�"O�!˵	C�/,aT�7�Ɲ��"Oht����"��M����n���� "O&�8dү)�L�QG*�� �R"On0�p�L��h�M��'��@J�"O���-��z� �`�?��Ѩ�"O�� U'j�@B+�?zq6p�f"O�����HM'p��R�2D�YUeDz�<ɵ"�'g����,s����^�<A�A�WLd1s�,R'\�(š�@�`�<Ye��ʽJt��Y�&���\�<���P��SU�>:��h��NIT�<���%j���5= 6Q�q��P�<)C�
~@��5�:�IS�<y��J�z�h�a!�7�����V�<�p*Qj�8� ���-2��a�0ɘQ�<ї���R$�&d�-U9�0��V�<	�͌�K��EEƅ�F`(���h�<1j@f-�D�nֆm�ʅ�Vk�h�<����|4� �,�8K�Ɛ��N\H�iЗ C
�ֈ�d]�"~�	�=H���e��`:�}��	ցu B�	*�yqdg�.�S�����FtB}h��Ѱ�V� �>O���!�K:��D&ֶm���1�'���ʆ�#U1���uC/Px�̣@���� �CF�_����'�|���HB\&Ri,�0RCԢ&���t"�	C�x�C�#�8�j#iD�1%>���޻Lb}�g �V!JL���"D� ���I�@���yf�S�N�N J�d�\9��8,�d�4��t�ĢN�#|J�੟S	 ^��g͉m(�Ah64�ж)�9u i�U�HMu�ń�m��h���_M���XI� ��I�V�'C���Q"��k�-͝W�A�˓:�@8!�fۛ8��R�H<g`0�%��i35��,��j����Z
e���1�O�į�5\�Z$�3%��Q�h�J7�x"'�4%�r���%����K��u�TSʗ-S��)-x����26��ˋ�$�!�䄥}�V����^�u����0�WaBD��H�?Z����/ɾ�v�!� �~�T�'~���s�a�)ńͺ��k񈁄A��![�@?��r�� 	H |
1ᝇ&���0���1�� ���C'�Q82�A	�(8!shK�N.\J��<�I�.����իɹQk�m!��W<e��D�/'�L��ǅ]�Z��Ih��
?c���$ˊ���ܻ��Â |�|є���J��� -?x��{����-�T�ê�&x��I��ǵ���L�6��r��n}dD3qBouL�t/�?+�����<�"r�ϫ���0���"�&��F"O�H`TJ�+��]C֪G=}f�5�¤�C��������b�l��W�\3,M�FhW=�����{�Ā[�ei���P��`��3 OQ�y�˦m'�O�ۖG�	��8v��+|���@�I���T��%ޏc�>��W�
s�a�*�V��héx���(��&��S�? �=�#�J�pp����g��s�]8r�#Ռ1�cCJ�rt��Бg˝v�iH�m��99F��D�!$��[�LV>��S,�|N
j� ʻ7�l�Ї�C=�ax�Ji U[c��]F͒(i-T��Ԧ47C"��5��*�pI���Mg:eä^AٲR�V�k)Z���K  B`}��k�!Pe�|�"FK�`��2�'�0Y�g��yan�Yr��zP���!�@rlЗ��#j��Y�I�(a�� �xaj�yJ\���w�Ԁ��ĀV/���R��2�MYߓ.�lM�@�ܖq�Ġ)�jU;h޼��o$Pu��'� �M{'pW䝡�� >�t�B�蕫u׬]A�E�N���sWi}2�>h��ɀ�� �K���H�n�5��'K���F��y��Iہ�A �py1��nI𭃧-C�GHdf��1kL �`�֕~&�A�@�c�D�P���NbE��BY�'�F��\I�N�:"����Ұ˔/?ҭȴ�/G)A�Q�̢�Rɚ�A݊M�^�
D���$�0�,81�y84�&����$H���͠��A����	�d���/��ś�A�zɌ�i�!%i�"�"�^=�-ȗY�D�vN��.����@�~π�؅$sqÕk��G
٫e��Q��Zۓ{���C`b�;\��$�6+�"x 0墎8%��T
`�V>|�N��`A�V$�s2jN%n���id��A�}�	A��S�������x�[�홌i��1��ݚ^ 8��>a�&W�M�F<���a9*��#fзult�ؤ�Ű�����Ώg�aYD��#B!4�s��+	���@�/ДCjB�R��������ϓ7L�E�$L-�:$���ϛ-c�(AC��]Mޠ���B0��bO4K�]�e�/�20��+m�sD�!%���
����@V�ɑ]0�"�٠�p?	ծ�	AÐ0P3LG�3�<4֮��R�2���2�h�r�.�fઍCu�B
Eʊ8P��7�(KVn���P�I�(���*W$ϱ~~��ir@��a{07K �Y���e[�9���E� ��]�&��e���#åI1O�X8[���iM�TK�i\�2^�۔n�1!��M�vN7g���;��O�MJ��>��d/�b��T�"�"�O�u1𬋵M@��f�&x��3�ĚξT���5I��l���<��l��kX�f1�6���2�� 8��D�Rk��e4�P�����0��5��	�T�b���*5*� C-�(� -�7�Z!T�D�b��1��9آIS�U�B�!.<>�@c�/u��sU�	(0l
 _�1��r�)�p؟�X�M���R�O>?ʵHe�ݦɠ�,7����Sa\
Wf��h����B�Ϗ��MC�J����&ϭ~�;��G�s��5�P�]X���T�h��{�GV�r�&�c/�X� ���HM8��� �M 9������Ѐ�Is�"��>���£�W�,��ܛ]���EyrhH�?�����mڔV�(�|R�Й�V��㉓A9R�$NV?��*�K��тH&ps���d�Z$6j�g _0�I����;hR"C!7y ��%#�t����/v#��:b˄�C�H�s5w>>���%[7} b 2�'��pr��R�@����n���kJ��rC'%;���K�' LY(�{�':�p�Z�@�P���I��J�*N���b��TH�	E���Ԧ΅mcȓ\h��;��Q��!�K.D�p����hAe�DS��yV��(M8n��ȓ[^P��VjP�}�x�������ȓ���z#��F8s5e߯)�D��a��T��NO���|�(��S����XM����(EA"�!�8ɇ�Uz�H���Ηh|2Z�n�!0ڊ��)�B�wō��,�a"���,
���I-�͓u����6+�� ���X�܄ȓ��������
��Y1
� ��pFz�'QMp�G�4��]AL�J!�|z��h��ҏ�y���G�(D�n�/kX}�$�<�M��чm6��"~n�P�� ���6�@1��O�u�~C��	#6P�;�\�bJ9��L:Y��j�D�H#J9|O$,+`-%P�\+��S�$�M�P�'J���AXğآ"F3s\���g+Q�U����¬3D���0'L7ek���
*��9y֌0ғg�Nl�C�;�'���1�͢HT�z���&S�,�ȓ`jdIF	A�H�V�6��oV���e���?E��_�Bm�<cU�ފAԘB�F�'�!�䔢3����N�lڠ�e$��R�!�Č�@�F���J۸9�����!���R�� �0m�(.������!�%T\f}�$ʀ�A��ZG�ܵY�!򄛾H�xՊ�e8؜��.�%]�!�$Ȳ(�&d��	6jŔ4�M4�!�1"p���m��x$񐍎�p�~r�DBǊ��� 5�*Q0Q��I���2w��[�<9���x�� �!�6�YpU�]R؟�Cb�ɟ�� |��g�65ԑ�1*���� ��74���e��(ꊅ��+W�C�.|z$B"D�����)�&���T�sF(����"D���#�52�h3ϐ�3�ƨ3��>D����C��]��R�N�xB,ڷ�=D����e@X�lk�J��k�x��g7D�8�É�)��)����$XĲD��E2D�|�u��"1D(�'�*o��@S6�1D�Tأ��&H�U�e��$:d<��.T���4@����y���63���"O��{2`@	����՝6?��y�"O><�A��tǰ�@�ՙShU��"O~H!v�<h�F-!�E[ 2�PB7"O�h؅�%7<t}�t!Љ"~Ը�"O*y[g�?�ت���x� �0"OZ�eK��/0xA6�N*@�ً�"O^�4FGtYt�� �R�B�ʰ"O֬���Q"���y!�E
&�v�S"O�`{�F�QH%�h�1т���"O�Ѡ����8G��!�ϸwǀY�"O��&Ā� |��K�G��>)�jr"OH�G���L+�\Y2̗'����"O�M�b��t\�f���!;P�
t"O���UB2~*���p�1%Q�"O��@�ʇ�t e�s� <?��Z�"O.���8Ė�� ��E)ҡ;�"O�U�'oÖ*4�M����5R��|5"O ���CO9\��1��'0��q��"OH̪)�F�ʭJ�9��K"O��R���P�(Hh�,@-D�P��!"O����D�E���#�����r "O$l��ʼ4��B`�$pi˵"O��� E�t��zF�
��1&"Oڥs�gX
S��r�!ڴ��"O�โ���EZ"�ݾd��9��"Op ���M��PD�C��m�l�i�"O*h{����T&
<[s��Y7B��"O�`��&G=O�a�l�1DɃg"O.��OS,c��i��\�!�Ry��"O���Sa�����&������`"O<͛%�̆"U�u�6l���ɳR"O��8��4w���ŉU�U ||S""O���OU��=�4�|܃#"O�K��Ĳ,��1Qg�M�p��"O��c��,nCE��70n�s�"O�pyÛ�F�[2�!O���d"O��*2��8�L驐�����!e"O�t"a�2;���:��̙B�~��"O�i�`A*JX6\AA�-A� �;"OlT���U\}���ǒ���"OL= V�N�)�n 2��3���z6"OX�*s �0>,� ,:@(�}�6"O�I��N�1h (5ѳk�y��pW"O�h�a
 b4�q�SJ=+@]c�"O M��$���CF�Ҝ�!��"OD�h�GW�6��[���{�,8�"Ot��D��v������<�����"O�љa��a�0Xq�����#�<I�o$x�I��j��7w蕉w�l�<y4���ML�H��$��t/�Pɰ��f�<A�j�Rv� V��W�,D��U�<�C&^����(��F�y��j�O�<�@�׊q(���c��{< ��5�@�<�p'��yO����L�d��%P5&C�<� ):��P�omR a���0�2"O>DqGf�+	/T�h��f�ИY�"O�����	��|
�OBK�})"O�8�I�'@V0S�E�' ����"O��A�J"��Q��o�hw"Ov�+��K+�X�T�BjĚ H�"O𴣄+��K���C�?\��A"O���P�F1Ct��dWz��"O��0��ny���E�T9ȡSD"O��ҕ%�"!��x����!'���"Or)뒍�8(�&H��Z a���"O.9Ib�E�W6�Ԡ'挭�鑧"O�� ���`��R���"O���W��F���Sҋ3 ,��P"Ov�4�ɵ"�@�!6�+aӦ"O��b ���83t������s"OVp���ۧ`\Ԁiģ�\��"Of���b��-1�UJԂH6z�`��"O�!crJF�v��Ӵ�ZoL,�&"O�(�Ίp��(�Ѧ��u\"\a�"O�Ac�%T�M�7��[B��b6"ONz�޲�l��֢W2c��1p"Orq	��ͅ!#� %���]�`�"On�����Q�h����B�=!�"Or�*�$C�`Ѻ�_�E���"OX���bF��9R�� V>�!3�"O��D��!w^�����ltV<A2"O�T0��H�U�Dy�A�Zc<��#"O01�R�Bq��	J��S53d%��"OV����G�it1����r<���"OM��k�{R���.^4WGb%{�"O�-��� z��@��1O�<�S�"O�	� @Z �y ��+ִ�KQ"O�H(�!�:� 1�RS���A%"OtsMU�B*ތ8��,��ċ�"Op![Tm�0X;����� -��q�W"O\AI�9���C�)�<�B"O��P�����������>U��"O�ic@ [� ��I=���D"O����*��
�h��aG:Cޥ9S"O�9�g�\(�������Y��"O��R�U:��i{%���/���"O��ˑ/��	6J�s���r��i�f"O�8��d޹e�&��V�|��Љ�"O|�q�f���m�!x��P�*O�y�U�V,��1W�Hs>\ �'y"��Z�*MD�w�#ua��R�'oT(���M�4G�Q�H��)�'Ll��G�Z�y�Fa�}Y����'�Z	X0���+�S(��Z��?D��J��Vg �a���=L���+wA=D�|����=t[�A��+�5B`�r�=D����06D��`,V�K�@�s�>D�Ĉ�C�I5h��IN�s�>D��*�F΂Ri�u��a��#
X��c?D���D�����<C�8 !A�:D��iaG.�j�ri��XFB�C �;D�@B�*�3=ځ;Q.�B���)5D�tA�ڵEk�}qG��.K��5D�X�#j�-dD��c�	�94�Y��7D����aJ,,���$a!�-Y� 3D�X@��I�e��i`��̇	���uL1D�D@��
z |!��� �@e���;D��ba߸ ��p�`M��A�����K%D�� v `�H����'�*u1"0"Od��v��'V��I�L�)-w�Ⱥ�"O@Y�fլG*Ш�lĬvE$�(C"O&I8TBD��,%aj�/��X�"O�ѫ4ǘep�+Ťɶf`L"&"OģuF��%H:�� �@�]N!�䃄L-~�V���i�r����A�x4!�dȳ$ �u+#�|� ����:!�� &>�"eA���4`TB�> �!��wI$�+��H��SǢ]�t�!�D9]hCI@�P%1H��U� m!�B�T��F I�&aԫCMC�1>!��	�()#��7B\v8%�
�x�!�$�6wE�Zb@	�Zdr��*N�h !��R�l(,ҕ$�|f�(P�^o!��%i�DrJBW���f�*F!���mP���;!�*�!�D�F8!�$ڈ�:�ࡧ^�?�t��ƍʫS=!��6���0%�H�<�����!�d�	|�|p9W��w���I�(#!�dƴX,~�W�x'�ΰBw!��2�<)Ѷ�^�|�`�;ׅ[2n!�d�h�n !Ei�T�&�r�D� �!�D�[j�s�Ǘ,;=��C�d���!�$�v�
R$ Ё`n���=t�!򤏨&Q���0K�>a��<(�!�䕃f��K�a�7CQ:�ް`��B�ɼP�0h��I?l�� �%P�Ed�B�I�@�\u�6��6#�\!#�01�B䉹#X�y�ܥ���:�%�i�B�,`ު}� ��|�<=k�b�J�VB�ɔl�L@ї�ͫ	�A�"��?(��B�	$d/4}�����2��Z�ʂG��C䉎A^�Ը��1<�l	�Î�<��B�	�/�p�[�Li �YVn��/{�B�	�k�1�eYV)���?A�B�	��\�Ц��/-@	Q�k��C�	 v=�8����_�U��B���C��"jY\���K2oq���%��qe�C�	'�YE�"s̐(pf�^�B��	Z�bE��i��6l��"ɉ�|�B�|2����v$2u�'}�@C�	8?ip3�9V2̘6(T<�C䉁
�<ey�h�,T���� -�&B�"D
Y)vMG�,+�	x`�ˊ��C�8L���B6�
m�|���F"��C�?F���T�A#21\ /C��C�IC�$l��ؿFj� �M�:�vB䉊y��shܐEyz�A��bFB�	�"k^���%� ;e\}X
O"V%B�I��z�{@�O�&#~�كo[�Z�FC�I�KY�1[�C1PZ,�����8�^C�	s���"���5�k�\>C�	�-b��
�*Su����
�C�I�luJ��eCU!� ��K$r]�B�I�/�$ء!��>n��ũԝW�B䉰b���!�D�I�RT���^�B�	/n"N�9AC<:�*��f� �JB�I���(R��B�(�fE\�E�dB䉕������T3P��BC�6xfdB��9)�� �AJ���	�cĜB䉟Q����>:��q�2XB�ɶ���z�L�rG�ijB�	�ȡk��${�)+�cF	G�C�)� �ѱnI#���#@H]c$X�R"OJ�CD��pR�D[	�E)P"O�9	֏@��F4�'O��V��u�$"O@���. (0���\>s��X�W"O���h�
^h`M�'3@���"OP!#BN�9�@��@�YKvQ�t"OV}3P��1-�T��r艍�|��4"O8�(b&V H�^��S)ֆW��!2""OD�(%W-0�`5�敯����"Odl6oBf���>w��h�"O�Yx���,%�2�����m����4"O�@�RK��>�^Eqg���E��`p"OѪU���<�R�� d��q;�"ODMs'K8Y<1�a+܅ڥ"O$Ey���:���AdŗZw2}�"O�-�۽k��Y���$2*��e"O̰Jbb��3�ᓣ�9'2A�"O,����V�Rh���-~�("O& �v+�$_��e3��5�IPD"O��0��D�Z��d��z�A2�'���bY�t��O�+v(j��'��1x��K��YI��Û�����'����h�EW���%�#<R���'5J��1$�*-K�F� ���@�'��m�����g�P�yyV����yrA�=�}�� ?�B@z��y"(Z�%�4^*�P���T��y�-	X�:eI�эT�HК��yB$XynDk��A,p��Yv,*�y�D9%V�p��ₖv�f]"�O��y�I�ju��#��6~m������yb	Yfha�)Z�y���Q����y���
JҸ�'�{Ȳ� #��y�a��QcC��{���kqd	��y���up�� ��E��!m(�y�'W{`�3��U\����yb��"6s�́�)M.I���[qN�y�" (j�y�NX<3�4�����y�O£Q �$�`ID!� h�W����yrE��0�n�r$�&l������yr�W�U�d��Q�ӻ	䞵6�A,�y��WމIP!|@�����y�-��4PS���Ɯ�X(V��y��͂��ի�P:2�M!E���yB��	BE���P�@��0�e��yB���9g�,�媑-)ࠢU'��y�d�>"s*�
!��?,2�je�H��yb.7n�>�)R�W-��P��D���y�P�,��u�p@��-O|���y�iӡ;y�x��l�P��@�� �9�y��/:�z�JȡKr��׮J�y�F86@�9��4C�b- G�D��y2+
8 4ze�V� ��%ֳ�y�	]<5��xD�!>4|��L�<�yBA_�>�d�:V!υ(�=q�jA�y�aT̅�w�G�T~�����y���ؑ�c�@�@M�YY@���yRe����b���/<k�e��/ٕ�yR�_�q�Du���ѫ7��Ɋ$�y"/3���s�AMVX�@�4fC�yb��3vۂ�Q���H(�]�@��y�Ĉ�&v��
@!��V�!�b���yB��Z���!5��Au�R��y���t,���!��r�xe:bŀ5�y
� z�ѓF�Ŗ%���/O8H{�"O,���"2������JGT��"O���IZ�*I�:�jګ&^���"Ol�X�I��p2�h�I��Y]8
�"OHh�eh $'+ũ��Z#@��"O�ݲ'��k�)3���^$)i""O!&aÅt�~e�P'B�l�E[`"O!$G/o�Xy�bH���� "O̀��%V��H(�4�Ys"OXBT�M����2(�&��g"O�Jr���:������ �&"O.ȸ�ͅ�$�:<R�j45���p�"O��ra.ګ|"�8����9J(dͱ�"O��0fN�r1��zBA@`��9"O���vD�*V��x� ��&by��2"Ox��3�R�.���+��˒~���1"O�X��b��I�J����b78O���K��9� uX@ ڪq��d��M��M�t��\FZ�ʳ��	in ʓ;Qpa����]+t�<S�!��g(.��0OD�ܱJ�)��%��q��B���!0�O?hݺf`�&L��:r�
<�+壖-k�i��I�O�T�C�0�0|��	��2�:��4ď�a,MY�HU�/�� 3�'B����E�Va��jX���_03n�S���x��������	#Æ�(\Ł�..��`� �2n�r�=+}D���K�
�:$�f�ު)6�ܻ�g ĦyE���k>�ZO@9tBP,SfE�2x��i�I� �nHʦ]��,^)p�Eb��)ހTa`���o���Bc�Z�A&F���1�n>*5d堅��P>-��Z*9�̪4�Qs�|�Fτˮ��s��,Jb�8����k�N��	J
B�"y����@O��!��(��'Ўe��������@ �O�5A�ᆁ�ё����^��s0I�l0� [�9�(���]�B%��>���2T̀�QpL���D�T�l��3�Z�C�|q %gӶ� �'z���p�Aed���ֽ=�����ڹ��Xvaf� Բ�����t�O��0��HQ%2;tL �A�A��ъ2���5[ax2��m�f�6Ǎ4�x���y�k��3"p�$'��.�z]ڂ�Y��y� �0�x��a�t.Ѣ$���y2L�=��P&�:<�]9k�6�y�郦YR$���Ҕ��18��F�y���zKеcg�ϴ�06�¿�y��̓R�Z��� �b�{�@�y�-��0p�G.�.�5N��y���,(�Q C�Y�b\i�	��y2�ȸ�n�����%|����!� �y"Eϭ*:����n�f�����y�E�)wC"��aܐaR�P�>�y� �UO$��O��1�24(��B�yB+
�Y;x�B�*$���i6@Ʈ�y2%Єn-�5���Y�k����D��!�y� M�j��q@E��z�Rœ%l��y�f�-?�[��؁wόl�����y��Ǳ%�!�&kA��B�y���< ܎`��@�>��8{t�W:�y�B0�R���V���uQA���y��S�,�a�G�=D�nH	1ȼ�yr��U��iH��@�@�����ǒ��y���mrP�i�BY�3�$16�\ �yb+�*O����,��2� �"*��yR���F>V�a@ǋ�0.�8�"�y��F%X��9[0k'$�%��e@4�yb�Ȑv"������4L���H��yr�Y"I|���EH�j�p�I3�y�n�<�Ȝ�@ Gn�"C���yrVK�d���4v.HX#R�"�y�&0���9�h^��z��\4�y��y���B�+6���:����Y��,��-��Q*�6���G�Ъx����S�? �}k��ƨoa�܊eHE/b��@��"O.�d���[�^{���04�l�K"O�U�ҢK�M��8 M��r��y�"O�0�(R�u�Df��1_���5"Ov"�ʛ�=0�EH��ņ2U|�KC"OF���,_
#�P���lI*@^�9)�"O�hz�� ��0��<E���"O�͸3	�="�-�#F	Un�A�"O�� ��4U	�1��TL� n"O�)�m��K�RE� ̓sL����"Op}�3�$��kF���0�"O���ÚS��l��GT %�C"OX|hԡxs����U<=w���""O�ԃc�ʩ
B�A��r���"OJ�-ެk��z���-A��ZE"O�]��MӉ)�L��1���P�lp� "Ot����^%u��);��Bm��"O�d"򤁻O��	u&�.BQ~$��"O ]�CV7)NN�1[727�e�u"O�]c���l�hwd>:h��q"O�#r�AjB�(�A��e/�X�3"O�ͱg�0z�␕?.P��u"O�ȳ�@H�&����,0~3A"OL��׹!=T���8K�P�"OԽ[d!��P�T�s���f\��@U"ON�1*�C���J��5 �p�Q"O�ȁ��Ƃq���Jf�\��}�""O�m����RO4pR�$�':��t��"OZi��5j����c	(j�2�"O}��,�4]�zQ��E0-b���"O�t)��;!�p�w�HIGY8"O2"�f��@p!HB̨|F�țb"O<�ԍ�9�d���\-)z!��"O.1�&
}�Y(��C�e:����'r��"/�pyvb�:s�Ru�ψ�s!��_�)�V!I`��!y�m�.�s!�$��E{b����� 
J�Y�&-z!�ċkL1`a"
�4�RY�t���2_!��ʓB�$�b���$��4+�/��w[!���_5�	{6�I ��I2$R��!�9]�z�����%r�� `�ҫ8!�G�hb 4�����r*��Rd#ãK3!�D�v\~U�t�50���Θ!�Ւ�����gy��4kT0(H!�䘎Ƙ��A�\�b ��[�YQ!�dH��-#��J�${�׿[M!�U�,s� ��P|#H�WLb-!�$������Т v`[���8~8!�dA$�Y����@/����cC�SG!�d�]@*�BYa�Q`���4:
�''^H��D2M@��Ԫݎ'T�*�'i����FS��Π�iG�v���I�'er٠�HBV�8b@A�2[gni�
�'�h���,�#qΤ��6��a
�'���k��K� M�*V����+�'iZ1���ÁB,�I�I� X����'c��2!���Ql��K\{BF��	�'���SGMM�T:���sA��	�'�4m`5@� /H��؅�^q�њ�'�\���E8]��b�E�$��'�F�,T��ضⓘ�������yrʞ=,A�m��"$�$1:���y�ɛ�v���	���+0����:�y'�`J\1n�|�Ӂ<�y
� �p�kC/^ƈ��A
n�y�f"O�)+�L�NIz!Cm��.� �:�"OP- �&
�L(@����~r�
F"O�T�e�	�A ���bQ"Op4)��2M%L�s�M*�5"O�U��C�F�n]��!��bE#"O��t�)��8��:]��a¤"O���D�C��4�m@="���u"O\�w Z/C�XHq��,Q��X*�"O����㈊
E� k��±[�"O�T�NL"HP��DG4��ؙP"O(�B�Ƣ'o�<�$Άq�>��w"Ox|ې�-.�U�WP�P�"a� "OpQ1ee�(V�z�X'��14o�iK�"Ovy�p&�\����[-8Xz�a&"OX�zw�G�}�H���ѸM� �Qt"OV�{S�8,�X�����k�"Op��+Gu�	���\�6�H�"O��R�K�=-[c �C�T�kc"OTG��z)���@�TM����"Ohq�6��:�>��T�^.>|��"O��X���	d�Iq�Z�KtP�"OL�X4��>��� �������"O�MR7L�q���I�%��"�8c�"OjE���S���4A��K��`�;�"OΨA�M�++c��s����r<["O�-�.� �<�"��61M�a�"O4�I��ū��~����gBU�!���
��4��W4d��e2�A1 �!�l=�hK���4ݸ�s"��\!�D_�X�@݃�\��4� ��}S!�Ɠ_��1B'N�cѨiVEa:!�d%'���@�$E�n�7!�� �125E�8O�03Aбq"!�DJ�T�`�£�58��}b��T!�� f� ���Aо��a�L�U�!�]1:w�Y�ʝ'���Z<#@!������#p�hsīМ~�B%�ȓh#RY����E�@�A)��M���ȓz�|
�B��u���b�ǔ5j4؇ȓ!H&��raL�)��īoT+����ȓv�ԣ����x@�Ed�X���ȓ,�V5§i�*�(�N*|¼��"l|�1�����b%��N����B��4�J�b$CCiE�B*��ʓP� Ca�uX��	[7��B�	�u�Ƹ t�C�C�
�0ͅ�<��B�ɭke&���	!P��2�)z�B�ɟ2���BIa��(&�@�\��B�I�<e��3AK��	�p|�&7�B��9P��5*��V���)��٦{;
C�	2ZVt���/��f�%S#��/E4C�Ɇ��,k�j\�X�A�pXȇ�Eb�@#-M%���Rw&�_^��PB�{F�������
�^=�ȓa����U�*^O�X���8l��؅ȓn�hA��BИ}����G��Q��C��}bӍ'��ː�ό#*F��^lX�Q���7h:�1�d�%�01�ȓt���w�E�ZY��XHF&l��9M����Ԛ.�Bx��  N�j���:o�ݒ �*Cʺ���MR�Z̅ȓcv�3� �V�EZ�dM*�X�ȓ7�,X w��CT�̙e�]�'�q��S�? ~9��#͡K��w	:'I�]�v"O>�bp"͠Ud�b7�^$C	Bذ"O�!�f�גCc��R"��ʝ`�"O�i�K^ 4�M��B�UZ�	ؤ"O6��BDN���'�Xg�T��"Om�ցX9�<��a=,���y"O��@���py��rV0��"O�Q�n�%ig��a��Z�"�I�"O�XҴ�>�p����.�4��7"O�[e�T�u��RL ��w�{�!�D�����Ew VPҁfP�Hq!�D�(u��i�#��@.��C�猟l!�2�,͙�S25Re���w!�$W/800�U��00an�1#��"MK!��E'\1�B��ˍYN�'{^B�	y����fCL@�0��	VE�C�I�l����qˉ�^jy��ŚCڶC�ɼ1��`8!�Aϒ���k��;�VB�I�2B�b��1���E�Q6 �B�	=1X;d�ÄWyȠ�3��B�I 
�p0Ů<4��R�J6b�C�	 K���r�_�er]��oM`c�C�Ɍz���3�oЊ��Z0�]-��C�i��?΀���	�?+�y�q
.D�x҂�K���٣�Ľ&BL1#l(D��.K$_�ra�c�`�9�%D�LqUG�,f�REO�*cX��Pa9D�$K5��:sy�ȱ���8A�H�+6D������CP��y�AU�b��Ѹ$�5D��F� ~��5�rō9^l���U�6D�zcĂ�0�&T� ˄_D����"D��xc���8�ȫ��C�s�ơʆ !D��2�d������l�jhp`�>D�X��K^�y�ݣS�Ƒ;�hh��`0D���CjG�O���a���ۜ��2D�0��� �`b��Ǿ9���s֎1D�x�p��/LKbJ[�`�l9�P�/D���Uq�ѣ���EvrlRE�#D���EBϑ1M"�§�W�tؚ3e�?D�����ܭo��@�SM�4�j�*D�X�6�!n����
�T��a�*D��s���.���Ԉ�m���r�(D��KH�G����&�7d����k'D�l�u
r<�A(�
�rBC%D�g`X7%�@��c�G?tK��
d1D�8¤�@� 6)��K2t���) �/D����   ��   T  >  �  �   w,  7  tB  =M  oW  ea  [m  �u  7|  ��  �  G�  ��  ϛ  �  U�  ��  ڴ  �  _�  ��  ��  (�  ��  W�  !�  ��  ��  ��  $ � � # i! �' �-  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b��|�O���;�'t�4,`v�K)�����Nk� ��+:�Zwd�gIv�:�OD��|\�ȓm�@ � Z�n��=�䢜5P^ȕ�>9������C�z!�1��ϫ>��!ҙ�y���pE����J;@<b�Q�A;�y,֕~�詑s�d�� ��'��y�i�6���.�	�I&�A.�Ң=�;�hO��T�W�{�h��/W\}z�6���'�q�"Y�3G-LJ��1��W�|�6()�"O�)23��5�ڄ�p.�3{��[��'����\���0�E�
���V?f%��}< ɓ�d:�r�$�)�8�r&b�'y*"��R�D/v���@^?z
	#� [XC�2m�D��#ޅLؐ��p鎹kR<$ϓ�~��퓟(�	�S�٧qFRC�� �V�IH������W�qJ���h\$]�p4L��'�a}�,�*�a���V��<�tM�<�p?��Osd ��9Dp4�5.�.{�zB��|�'�~�86l(1�,8��Ύk�(���'81O�u�|rL~Za�%�lm�_���/U?p��C�I�Cw�xY"*�GN�qJ�'���˓�hOQ>A�%'%�x�P�K$!{<�9B;D�Dz0l�^�j�4�ڵV^��DW$���"��?�HI�jݍY�����(%���f�<���L_��:p욫,�$�⋈6~�R��0?y��!`p�TZ�g�B"�h��{�<y ��,E�`b�㉙-}F512��k����'�:�Ѡ�6%j`�i��9U^hS�'OqOX��d��_9Xd"Q)��FǖiEL�;&�!�� \��q�W.fk��Z;2��(w"O�Y�t�X��"�!� ^�����'��V�!IG(��I?!�T���j)D��A�H�X���'fG&�.]�
"D���kI
T�v̒ab�K�6�#�O>扔	Z�L��LG-k��a���1X� ��V��h��`�ɡy�!2�N��pxXD0��'J�O t��AG*d}��9���<?�ɻ�"O$�4.Ư�^��^�,*@���'�qO�!sk�:J��qx�O Ud!��V�܇�	YRXjWA�*�\�m1g>`�<a˓�Bx��nH?ŀ�f�5WX�5���F?��	�<!:�Sbb�)y�� �o�[��B≊+�FQ2�R5h��b���4C�	�6�̡:��C/:n�����,cVC䉂iX ��@&U���v��;,(�0>��4%s�`�rB��� � �@!Q���ȓH�hp�A��uL`ȐFY���4��C�4a�"c�V��ٻDN:/�,�ȓ?|�i�E���д� �A�~;\8�<�����01��� N��u�
�
��˳O�qO�����L�O�ԭ@�{������rD���Ѵi�8��	#��lQ3�>o��A��(=XJ�<���;�$�.kpC�`#Y��H�yb�ʿ.���H�b�Hb���oA���+���>}�V̉�>NlJ�	æ����<D�Lr�H�=(��sI^JOHi�CF:��<y.�y*z9Hv������e�<qn��q��T��\)9<��F�L�b��"~�s��YS�C�� G����\	�2��)�����[6`�!@��,�X隷�.D��S��J4ν��`қT���`@���hO?���=3�`�����d��ȃE'�;�!�$U%!0в$��*� ��"$Cd�!�D�Yڮ$ȷNA��X���E�'9�zb�V=���{-�>W��i�6��zL!��],���3� 8��y�&o-�	�<YW��O4�S�4����S�N���&��@��CQ�<!�F�' fU�ll�(#�+*�@X[t��	t������G}� ��h k`��o�~��� �yR��2���`��C(`H��,���y��&	LY�B>�Y��k[��y��\Ψ��੄�{B��������ybJ�2B�p��I$xJE��O� �y����T����̡"��eK��/�y�!9�~�17 ��iv�A�M3Ǔ��'I�R�(M06�1c����%�y��Y6{C8��1-�0"I� 閧��'�ў����j!f�q��O[-	�c&"O Hj��۳Zdz�YQ�Wj� 9Q�O��:�oL��ˆ�&l�D� ��Mnp�Ey��Dܖ��)�]x���S�TS_��c$�ҋ%H�5�O��Q�&� i��1���9���4�IQ���PCΉ�C��Le:%��+a�!�$F�R�~��(~��5ԉ��#�fp�ɖdQ�"~�d@��0�9k���#
�		��4�y
çu�.���+� 3eJ�RE`��y�A��Du�92x`���͈��=1�y�`���a��Zy�b+��y�	�&z\l�r"_vT`8"b�B��hO,`D�4��:��=:��%�����y2!���sHM�t��D�PA2�M���)�禝I��8
v��	�4g��]F*(D�����M�:D}���/8Д���>��S�? �4p�H�We��ys/_�'S��Q�'�1O@���GE= `�:��'1JȕQU"O�	c�����@P�+E��|�>	��I�7o[�\�/ξ\�\5Ȳ��|'!�Ă�e�} M�8xje��d�7U<!�A5ʞp�R��i��t�3$
�9%!�d��s1�4�*nڎ�q��"��;'OxH1�U�蜸E��7)�qҰ�'���:	�!z��P7'�]�h�r(C��RJzУ6���E��2.� *C�ɢ5P��`E��*�9���&��"?���	�!�ѱ�eI|4@ic��Rl!�d��m�d��D��Fŉ����8Q�Ix���佸�T�!|<X���b���v&"���"|�'w���D@�c��};��� .|J>!�^s��aG�'��MQ׉�L��I�բ��Ď#��Jѩ�G0�{�f��!��\�We<��d菞5Q�lЀ��E�|��x�`۪`r��S�xT�qB�ڥ�yB�0��P"0�׹���g��y�D)*�t1S0�.y����#��1�S�O("x�E�1*�|�aQiַQ��01�'��u"��*�� �P��{�"ݡ�'��y�ꘓa�Hi�G yN����'ab!ıY�n�X�jN�j���W*_�p<��O<�'������-q���t�`Êy�����
���@��h9uBރV�E"��O��=E�"�I�h�'�Ȑ|���5hE�^V&l	J�8���]�˦j�uu�����p���OD%�=I��d����샵���"=���@@�	1!��I,DXG݂~!D�2N�Q�F�To��m�ܩS%�\���&O����x���7�X��uK��6vy��L	�K����>��'�2��i�'*Q.e˃=�P))d���!��*=I�cΒ���ȋ�!��Z*A\�@��Y�d���b�U�)�!�"8�Z���fK�N��|��&Ia�!��G$�|��O3�a�0慐\_!���#�؜	��g|@ydG��!�2$�x��a��K�]`g,�t !�
�)i&�Y�� �lB��".�3)�!�Dd$�����ζb@ܥWo�!a�!�$ɀl����-JR���5��r�!�,zԈ
Gܽ�*0퉏n�!����
�t���E�r���-�&�!�D:�l�f?P�HD��,2�!�$�	c~ ���I/
�D5hb	�n�!�Y��`L��o�9v4��D�D�h�!��@�XTR4KKd<�C�Ou!�dΚ��ġ�S#�ɨ�uu!�D�6,���0�[qCN97n!�ǝOR����Gä+�	���z����i�t�c�.���<1�P�ȓ��S��=_fq{4m;R2�i�����cD�_������.Za��]\p���l��3���s$�,:�V��A��h���[��[��߂0�j���Y��06dG�++��%�X�@ *���.�!f-�q��@�%:ir �ȓ=[�0��M�?_�p!Ʈ�2Fô�ȓ�<�Iw�A�d04��Y,/�X�ȓህ�Z�!�<C���%,걄�K�����K�$�ؑ�$T��l�ȓ��8���m��a	!B�8���S�? \E;Ǆ���k'��Ci�	W"O|e`�FJ�b�s�D��Sx2j�"O�lq��U��Y�c�b9fY��"O�(0r	66�����<&��5"O�(@� GN�� EI�4Z<|��'��'��'#b�'�b�'��'P6���Z�*Af�*��E�!�,��'�b�'���'J��'���'*B�'������G9��ؖ�����Q��'��'��'N�'�'���'JB��"�Y0T=�	��h�&Ղ����'$��'y�'?��'J�'���'8N`��C���)�$���dB��'"�'��'e��')r�'���'"Q�@f�9l�P!�� I�.1�U���'v��'��'�"�'�B�'��';�4��ͳ0�@$�3":P�A�'t"�'s��'���'�B�'���'�� ��O�Z�l3��:�5i"�',B�'wR�'[2�'���'A2�'o�`��dH(��p�"H�2ٴ��E�'�B�'��'"�'���'���'� �2�-�H&�I0@�
�]�2���'�"�'���'�2�'�R�'U��'( �
bv֨XJ�JK�Mb@���'��'�r�'���'���'h2�'|�z$��9���Hր TD�b�'��'�R�'���'�r�'
��'����±Z%�� $	T?f�	W�'_��'�2�'���'��"t�L���O:����D���$��D��9�<	��]zy��'��)�3?���iw u#T�2J�z��'�s�qag�)��������Q�i>�ɡ�Me8t
�y���G�J� ����'���'�^\`BH])�y�'�|cr#����#�O������+MP�i��$�%y��2��O�˓�h�Lmit&�k�4�&V��2�b!,�Ѧ��Ҫ0��i��:��w�
-�Gen����(T�P�x�P��p�(�m��<�O1��1�g���b�$���,?f�� I�OJ�!�18�3�
�\���=�'�?�!��,K�(�(�9 �틀N��<�*O�O�XmZ�FKLc���g�S1&���bA�Y������]�j��I��M�Ӻiv�d�>1KCU��b�i͗	�ͣ
�]~b��2(�Za��T��O�NI˗a��@U�� c%ʊ�+��;���hy�����dU�rd
}�Ơ�o>Ԙ�%��o��d�঵ s�-?96�i��O�i�3v*���!E
#hhp"�d��Ev�
٦�Cٴ�?�1���~�ؽ�'8��^ ���:���Nj�HF��[+ƩI�@�L��H��Ȕ�L�䞟^���_�~P����Ιw|�		DB�t���Ğ7���⁁��ze���7l\5�� ,5$t�X�'�9t������#���VM�l��. x]1!�*s��4�7oS*\�I(�$�M6�R�j� q��R�䞁\Q� x��Q-c����f��#t��hT&
�Q Fe�v��		��q0�#h� 穀	�а:ӧ�1�#fA�|�2x1���%Q����	5|*��`f��ӠP�r#�.�H�$�w�xA�@xB�Y(��ۧ~���B���M����?�����>�b(̤G�$�� <>\� z�˓�qDx�O9�-�.�C�����I�#a��>In)oZ�''����4�?���?I�'{t�'��`]��4��b%�(v�&�aG֎9R7�U���3�I����d�جi��!3B��8]t��L��M���$'d��O���
�4�~R��(ĉ�!�@(1�����ǌO�b�H�#�3��'�?1���?�嚋VM�]��F�U�s����"|���'��5��*��OZ�$:����iZ����%���I�2U�-z�U���`2�����	ǟ��'<�H�(��`��H�E�;2���̳CEDc��IY�	Dy����b}��,7ΌCRi�:�B�y"�'	r�'���'�`���'b��Ѫ�>��A��NFz����&o�R���O�=���O�DW�uz$
¼i��ˑD����1��Wfs}��'D��'�I36+�`�I|"�#-.�N�D�B�'<��W�v0���'��'���  �hb�`%��IpR�����lU63u�y�&��O����O���'
�|B.O��I�Q�p����I�&C=�@�&���	Ɵ�Q�M�1(Jc��fyۀ�ÀWV�K'F��}��n�`y��6��7�h���'��4F;?	E
�DsP�}�~i��nZ|y" ��O��~��c-W/@�e�eB�sNF�#ǹiX�(�5�')"^��S蟠��yyRy�4��B�R m^��*�>/��7�8c֨�W�������+5F��/W�������M���?I�:��BG�i���'�R�'�Zw� 5�87T�A�ə�K�@ѳ޴���ѽ01l�Zc9O�S�?����$��|e�Q#����1r�^��M��d�*	�V�i�2�'3��'�J�'�~R øbY*��O?�4�Y.ڔ���MC1��ԟh��Ο���\���/\�T`"�i��m����Њ&�>E��'e�8�d�O����Oڤ�Od�I�8r��֏�p�� x�ذ�@��H=������՟���۟�O�N�Er�|�C���b��jڞ,���$�ɦe��۟���䟔��yy2�'zAY�O��,�g��<g*��G����09� c�����O����O���O6<�b'S¦U�������蝗kd��#ƾ	��cS�Ԝ�M���?������O�Urr7��D��l��ۻd���A퀨��'���'>��'%р&�{�,���O��$�T}#���P �C>�QY�D
(�xo�ڟX�'&2�ɖ���|��M� �<�6���'<�|�PÍFp�5��i���'S�5J�dn���D�O����f���OH̀��0)��0B�G$b��!�
j}r�'�\IT�'U�\��Sq�	 
i~���*����CI4V��v��wr6��Ot���O����
���OZ�D݁'��i����r�z�1�U���0n�\&��I���D����'�!���n`d���׼q��i0�Gt����O���z�nZޟx�	ڟd���֝0`�ĴP�_����3��Z6��O�˓+s�%�S�T�'{��'��|�X�c���p7*�V�8&$hӂ��`�Hl�՟��	ҟ8����i��L���Ue<m�u�CX�����>��CF�<!���?��?������Џ#H�9��
D�YKE�\�&Z�Y,1\�6��O<���O:��I]�^�p�I7y�������<X& ���	ʂ���a~�,�����cW�Gן���ҟ��)[�``�ش8�93�Ȣr��u"���_�P��i���'���'��V���ɦz����Q��LY��[��b����݋`�9ش�?����?y��?���^]@��ֻi.��'X�ػh�,D�\MHǣ�35���/`���d�Oz�D�<���QΧ��:u�,�`o��-���4 �/(��6M�Ob���O�D߀��Tl�������!Ȟ,�Sk�-G��3,]�%b\[�4�?I*O������O���|n�4����'O$n� �I�F��9$�7�O�����N�ZmZٟ��	ޟD�S�?����g 8 ġR�ay�D��nP���OH�DL"W����O�dC��I!�4�8Ġ�+׊�$?J4�(���M�Td�����'��'<�4�O�2�'��N�q�����:����$Z�V�6��f��$�O���|bO~b�.���%$��̑��Z���dJt�i��'�j۠KqH6�O��d�O��$�O�

w����2�,X�X$?Û��'���=z�x������럸���O*�93�Ľ.������<j�X�ڇ
Z妑�I3Pn����O���?�+O������s�:�����hV6B�H��i��m:����yBZ�d�S����Iiy¡˚H��Eh��K�4c��(>��D��>�(O��<���?a�����pwF��7P�����|���3G���<�(O~��u��OB���O��D(	\nڻ3}���HR(0�V���!$�(�۴�?A���?���?!+O��D�F��7qwZ���+��#�0�v IaMBY}��'��'��'ݐ\��b�t�d�OH�H�$ �r%\`�$䌀�@X��\�����ϟ���wy�'��%`�O��O�Us��լy-���f��H4�2ҽiT2�'��'Q�fjm���d�O0��㟼�Y��7�jd�&m��*W��������ry��'zeɞO�ɧ��4r.L	r'
d����A���]�xYm��@���\�Tѣݴ�?y��?1�'����,��������.ia�F*7�P�Y�S�@�ɕoM���	j�i>����C�DP L9*��+"p�t��f�i�$�y�Dg�8��O��$��j���O<��O !AůJ)yv��BN�,M�����SԦ�b/�Ο�%��N�� (u��:4���{��QT�@!4�6�M���?��6��1�i�r�'��'2Zw�*�!��0���ha�����O�ʓ��Q��D�'pb�'mHT�!���A@Q��!Z'�a��$Q�&:�l��P������I#��i��$���*���C�P]��2��>��)��<�*O��D�O��$�O0���?Fb�@�A��iE�f��P	���$˦��ݟ���ȟdc��˓�?���9-�Q���8S��:�F�89:������ON���O���O��l&�}sZp�/?�,�A��F*x���@�e��d�O2���O��$�<���:��|����E$^�I#�F�w�D$+h�����OJ���O��O"X�:��f�|��Oҹ�猠+�qƚq\$D(2�֦�	�\�I{yr�'D�]r�O���Op4���7E��(���æXHˤ�i���'��&XˆpHL|������Y##g���4^�˅�T�8|�'h��
I��#<�O	�e��6\��L5GÃx�	��4��$B>@�)l4��i�Oj��@B~"��O��84a25v���N��MK*O<�s�)�S�z�XL	 ��J�Z�{�#d��6͐P}n�ퟀ�I������?��؊}Pc���&X����=W��Ȏ��O>q�	l��ݱ`��n��0���_�����ٴ�?q��?�qf͝==�'�'[�*t3Pl:]D�)�/(hM��}��@�ߘ'���'��nƖQ;�I��) iǼA�W�]�)��6-�Oxl���Aw�Ο���K�i��Y�.�,(���02ҙ��e�>a���R��?I��?��O���EY�+$)H�F��;�QjZ�v��c����m��Ey�O����Yr'�">Q�k�LZ�FzP�)�y"�'m�'v�;DIZ�O9��@72��قC��1dP2hɬO����O̓O�˓e��m�'7ą�n�� �T$+N$�O4��Or�Ġ<��D\�5�O��8��=G��P̴��e#�J���'g�'��I7dG�c���#É�B���Y�LK'28{��t�H���O�˓t����֔���'M�$���\�2�O	+ۖ�aS��( O��'� =Fx���3E�8'a�1PR�;b-�D�i��I�l��q�4���ҟ�����D��l;L`�fO�G���d�s��]�$	R!#�S�'5����@�&��)��ʄ+�,0l�<3�1��4�?���?��'B|�'r�G�tҶ�:F.�5
���� {R�7��r��"|��|[� ��`��l�x`G�ڐL��8:��i&��'���$@��O����O��
р�㗣ǅv���8Rń�f�,c���G�0��$����@���xOp���`^m! 0w��#�M���*e��땝xR�'�ҙ|ZcL�����0#lahFӟl\88٨Otq�����O�D�O��AHb�䦁�>�����E�R�CB�#(m�'�B�'p�'��0�p�cR@:i�abC'P���>���?�����Ǳl^h�ΧF�<�kri؃<3M*`c�b\�'���'C�'�Q�P���N��tY�S�P7��U�E��>���?�������s�&>!��K�-d��Ӳ�8� �G]�MC����p<�eT)�$���A$^W2Y�̈ݦ���ş8�'EX����4��O��iP)&$��s�	Y�%6�p�A�I�T��%����"|�0l�dȂ��%V0�6M3?A�J��M�T?��I�?��O��,�&�2�VoK*-�M:�i�ɜ<�*#<�~j�I�t�8�"�J 8��0�	ٟH���W���ٟ4���?�1�}�w��d+U� �P��c���w�6�T&-��"|"�{`�9���N���vE�.Sy��x��i�'�"�[g�b�H��Q?a3j�H~X�)��V�̨��Gv�E�F$�<����?Y�1w Mʄo�0]7�L���Ζc��J±i��h�n�c�8��M�i�����π%� a�`��/L���:���>Yt��Z��?Y��?�,Oi�P'-?��4چ�G=L��c{{���>��������ߎYB��Zbi��d&�D��F"��A�$�O����OD��ư�e0�H��ő*:u��
���#��x��'4�'T���x�5��e9��{|��ti�'�Q�'���'��X��1�A΀�ħiY(��v&�z0���F�m��	ᦸiV��'�Iwy�"P���Y��S�����e�J�ki0pc�-nӮ�$�OR˓;�(�������'C����Tޔ�I�S�̓&�A�(p6�<�*Or0{S�?��|nZ�T?��S(WU>���e	�'V7ͧ<����/k�&��~
������P�Ư�/ ��t*\�n��-�p'p���'>m�����Lk���$��r�KZ�m6��oZ�s8��ٴ�?���?i�� �'\�lH5�fiH'�ĐQ�p=J��6+j�7M���"|��k��#�ܒ�޽� ��8].)���i�"�'R$B��O$���O<�	$�L+�$��^�4yX`MO0)�c�H96M-�I�(�Iٟ���E�HBu��͙�BV��`��ʻ�MS��T�` 3c�x��')b�|Zc���VE[&P������İE�d���O��g���O*��O��bxds1���$J�"�v`�bb`�5s0�'��'��'�	�f�*l�0�L ���	�*�����/�ԟd�I� �'�����b>�(2c�`j3NC[���Č�>1���?�K>9/OB!��]�8��>[4(��̆t�t���>����?����,K;.�%>=8���(W�@7%�Vx�dC��M�����$]�Mo�O���ᖸ5�j!��͋�� Qиi\��'[剧j!�H|������/�R����άyR���ɒ�+|�'��Ɂ?�\#<�O�x2�)��m��k��Dv�f|0۴���L�P(2�o� ����O��)
{~��U�t�dX%n�B��3����Mc)O�d�C�)��R���Q5ί|��  5E�?4J�6��E�<�m���H��ҟ���5��'��Rv��	,�Z�z��r��Z�j�D�Y��)�'�?A`(�,�x��a��ӅImN���'���'��e�#�)��ß��]���!"�')D��R��$t��d�>	�KXz̓�?����?ab������w�*F'DxQ��#+֛&�'�F0#E�$�Iҟ�%�֘
p*��ф��(g�4D� o��`���U���<A���?������%QD���N�@��m��v�6u��A]P�	�l��r�Ily�&�	���`��@�v3&��c�Ƈ8{���yB�'a��'��49��LZ�OU�Y��b�W(� �S]�i^�Q�O���O��O�����''��*3@��yZ���R/K�@�F<H�O����O�ġ<Qs+U:W�O��� ��Z�AB���7��#����	v�:�D,�D�<�U��S}��H��	��阆�S�E���m������py��9d�8�ퟒ�&��=.��D�A�yp�<�qPt�CyR��O���#8��6�dF(@B�FU�P6-�<�e�	Z����~����⣚�@{򌘓�>h�q-�^r4�� ~Ӝ�ަ�Fx��Tl��^�ȴZ�IG�?�������M���?蛶�'�r�'��dk=��O����/B9���',Z�L<|(b&������%(�S�OWB�W�T��Ջ&,3wQ�0P�v\7m�O��D�Oڑ�%�Xk�	ԟ��Iy?9��G�0���x�j�Ao`Tjs�[g�S����<���?I��	�x�Q�ڝE�	j1��N��Y$�i3�BF�@O`���O����<��1Z��q�E�'*���&�;��'�Lx�y�'���'��	�� D�!i�"f�&��3�tac�bɳa��'3��'��\���	럨@W.ֈ=��1� i߬~��i	@̌��c�d�����ICy�Q+7�@�.-d<�`�c{�T��%#l:&��?����?�)O�d�O@!��\?�lO
������0�E`��[	�I�@���ؖ'�x�v`*�IٞD�
��`��ɷ��l��X��Qy��'�RAZ���Y����Ƣ&I�Z�M�.�@�y!�|� ���O��_M�I�M~���B� �$<��Q;Kt��Ϗ�r�'?�I.;�� �?�O��C!Kцj�P`+B%۸{� �4���^׺�o� ��I�O����}~�g��:Д�W0�����&�Mk,Oz08��]ܧi�����l]�p�v���]e�`l�5dي��ݴ�?y��?��'j��'w��DE:!aӦ�kAB-�r�G�T
6-�
�"|"��/�.PIa�Ð�I3��2!.��u�i=b�'e¦��5A�O����O��I�}�=3槃�a����/ɻ<&�b�l���.����0�Iϟ0p6�^3t'9 ��'|ytl���*�M[��Ri3��x��'ob�|Zc�V�c��-Y�}��ɩ4{�-x�4�? �n��?A���?1-O8b�f�w\��Z�eޮ��@1�(��"d�1$���	П'���IП��ǋ�*р5�6�M/`�6���c5DL�Iby"�'e��'���6GR�h*�O�"���KB&9�0`���(���O���O��O���O���;O�p��h٠qC�a�l��*'L`�n}��'���'��I����H|z6H�s� �rc�L9�dz6�J9��v�'�'5b�'�.��'��b��w��h�:�g`�zμm��	Gy���s����$���E��8D�b��nЄ�xU�KO����;%�>�?�O#b�8P&P�T@TJ����(���4���#~ Nl7��I�O���A�D�mbm�n�z}��{'nܳ�M{��?�@��?qN>�~�Ć́:Ȋ�qB	18�\�0��ܦ� dȘ��Mk���?Q����x��'k���ٳw��1�w�S�aQ��ȑ`Ӗ蛅��O�O>���(fTrͩr�	�]B���_�%vl��4�?���?�u�_�q�'�B�'���1��truD4R,\	A/��(��|"	(4P��F���O,�d�>izvH�g�E)vp8�LZ�x-*�nZϟ�J�����?�����۴��:K��8"'�7��)��/�O}b�!4��_������t�	~y�Ą<.B��"J�A���Ub�8N� 0aM4�D�O���8�d�O��Ĉ�Z�@ۡLK�V<����2w�l��8O�ʓ�?���?�*OH9���|b�H�(���V��LŮ}MHh%�(��Ο��'e��'(4�#��B鐱,SsfP	"� ��.ap�S���I��4��{y"A]F,�`,{��O�xd�@� R��p`�ɦ}�	˟�'���'�X-y̟�ɳb\�pY�?� x��̡`k6��Op���<���2Z[�O���OL�t�!I HR�͖�hIT��z� ��?A�������4��6�4h�c&�ѼH^�Ъ�C�0�M[(O�t����#��������'T2�0�#��3E�H c9*�ΐJܴ�?��16��*���� ��aST
y�uQ�'@t\o�Pc��;۴�?���?���d�';"M�I�'�ۻE�<�P�g�sV6�E�t��"|����&J�i�05��P��?6a��i��'�b/�K��)��S��Dѝjp�1���C�"lF��L�)��b��!#Z���'�?����~�I��	d$ �&���pUͶ�M�]�f= (O�-�Oʟ�$��%��˦�Z�<T� ��M��\�'z��NU�����Ov���<i���(@@2G��mt�I��V�|��!�����OH�d�O�s���' Δ�0�].��d��d�x��&�/#�"	�O�	�!B4b1���Qˏ|����2��C<ϧq��C�.�	*��$�*0���ȓ5��y�c��3���T��'"�8��=�Ԫӑd���V�
���h�O�p�M�V �`��A�Q�G�J����O�*�~EҀ(J��0���P
�bM���sïD�-��e;G���FF�ÿc���Q�	:xv� �CFP�"I����$�`tÁȵ4~>ʲ ��T�C苫%)h��p��A�혲.�:�@T3B�'�T�ƈԩ:��yS�i�W�d����'�"(W/��p䊚�:�~��U�X�:������2�]��l�X�h�#/���Ox=�"6)�pIcB��Y{�xく%��!É���TEu|�iI��� }/�ؒ�M��@�\��ۦ�Y��i��2E����m�])��S�I���24��"Kɐ4@ �$�WM�ļj�!OxYFzB ˉ6�����>PP��g�S�A�7-�O�$�O`�+���T2���O`��Oܭ;Eef�*��ܹ6��ʑgP$�Hx"7`�<2"�شvP�,*$�_�1�R��O�%�"��:kr �6!�?,�����+=��%�o����6D�;n�d�B�"0����8N��ͻu�D!ݶ6Wބr,U;lR*�(����䘪v��O�ў��6�P�[�8��bH�g�!s�b%D�Ls8ƣ�Y�\�C�����]l�����'��X�p������Y��C�*A+�y0�% [r����ٟ\��ß �]wu��'��0}��yb��F�1����SN�!V���j�az"��X�? PZ�"P1oeйj'>V�V (F�H&G,%�f����9J��VQ��['+YeqO�i�wsh�! cZ�	�x��w��$�������?���q2�����qӑLLO�<�aFX'e��|����6�� �gMH�i9��^y2��Z�p6��O<��6%�bI`#K�Ȑ��@Dۃ4���$�O� S��O����O`	0M�!�z8�@F� ��Z�O��`�f��'�H2y�P���Y�{q0��䄣dLQR�%	�0X��NN�E�J,3�E�F鮸1diS�=n�l�+/4�A���ΑCO>�T]����M�.��(�M�27���Ck�4:<��(O��$/��؟�����\��6F"ҕA�
�exXX�'N4KB�	��M��p��R&b�+<R�Pi�;U��6V���O��M[��?a,�B=R6n�O�iC�	N��<�[�n`:$�6(�O��ɗj�b)�d�;~�(�p�"�П�'���C"2.��ؓ��!>��ų���6��kvA��0QM0�A�����H�4���U���󆂧����>��͟��	N�O	r���hdҐc�)93�\h��I_��yb�\�BMz��1ψz��E��0<���	��L �UH��"�A�b�<��Bش�?���?�sE3>ݐ�(���?����?�;l&pR`��l�� �ѮU	L�T�z���<<���+fV�qÂ�%�3�D�� �|Exq'�4�z��a�H!)�$���Y]y�J��@�}&�VäB=X�b�.2�$aI��ӌ.tb7��˦����IYRL�)�<��
�$yxf��L0\Y#�Ղ*�.�@	�'��̩- &&��p�,��T��z�O��Fz�[>��'�Լ�5��%�$�3�f.t�t��-Q+�8B�'C�'���s�!��ӟ ͧNÖ%s�L	iDJ$9�́�*�X�5kL)}��d����=Y��M�0���e�
�}���R�O��n���X�ܣ��M"n������O,@rGc,�4@�)M�N��Vf�, ���'T�'�b�'J�OҲg F=@��$��E��5�g�'y�'l�̺rg��BZ�Bҧ��ZFh
�y"Hs�
�Ī<I�$_O����']����`=*�^�_^��v�od��'�2A�'�B0��KD�; u�a��i�>D��;zb���S<S��q8�����+u ���MM}�/��x2�M�v�ʽ7�F9��+�+�p<v��ԟ@
M<�A�ƚEeR���)t��I���e�<qb��0g!\0����/�l�
0�E�'ў�S��?��e@#6ݺ�ۑ��(T�c��s�<k�$�۴�?�����)�F��$C,�&�b�+ԻL��9A0B\(�d�O`�O��>�(�a�^}[>��O,�����UUOtݚ�h��b���KO���FnV��Ȭfs���ME6o��Q!M?I $��_�d�y�?�ti���'}�&���?1�iTf7��O��?��&\��u1UMͨ]}#K$�Iퟠ�	j���D��%X�KY�[-B��ejѣT�zt��	��M�7�i��'�=I� _�XM�xk�jO/l�*�"&CZ�D��'�b�N3[�l�!T�'���'v�bz݉s H�[�9���];��p�b ǥU �Fᐓ:; q���u���|���>����/�
�[5/=��1D�ۗG
��� "g�0J�N�{?�M�Ɓш��S!�M[��f����jW?	RZx�$
�U��9��lĸ�M+�i��$U�{���,OH�D�(t������̺o@�أ�Lͬ	6B��!Hx��o�*�(�a�K���՟|��$�7h�X�İ<y�)� ���zʓ;\���s
�+4t����N��?)��?��.���O�Di>��!� ����J
�@ �@j�@�k�+ @���Nkb^�;C&��8��c�=z���cgAY!@�pl!�'����Q���i�-I�x��]�/E��?鷿i�7m�O���?ى���B�\Q
$�SuQr�3��/�yB�"ξ�a/D(f�^�dj[��'U������D<κD���?)�J�"ͳ$ �XN�k$� 9��ap��?�Ģ;�?����T�{,p03�! �6�I�+߼*��:ƊV�!=Z���O��<r���G�YŶ}Ey"�֌=�	�p	Ԇ<�@c��6@�Z���#LD�@�1���QW��hȂvVLq������'QLQ��#щ'��P�Ӧ�Z��q$ㆷ+�F���'�t����2
̠�s��A�[I�u�
�'g�6-�'%���I�/cM�4iV��|Jp�O�!�TԦ��I�O H:2�'�"����!f.�(B��QoR�b �'_bZ�0���٣ ��uC�O�[�Ċ�'q���R��.��Q.��&jF�q��	L[�����J�O��L�Ò�^yHܒ5�T<�ЃI���%��ON$��?�xU���nX<��B��s��8�!$D�<���J"EϞɦ�(I֤<�E�5O��Ez"	'C�j!J`
E	\�9���*��7��O~���OV=y��s�N�d�O��d�O�n�(NF��#FJ�[�P�H��ٯL$��CwBU�Q��Ų�.��p?@Y�7D.�����M�ԎY�J\��0ǂ�!,f�L�c�T�J�~58���g1�+˄�?1/�VmZ=�� !!��P�s��]:D	�M�J�"E�UҦ���4�?��H9�?�}�'�bF �#R^9��ΜF ��I&֭N��	4i�J1Θ�M'���Db�80�D�Or�Dz��OL�[��Rs,Щs$&A*>-�(#���ri����t�������.�u�'�8��ă��ü"3�Y���U w�%�%;U�*�e�-nz��[t�]��p<�юA�hZ�mcs!�����-��EG���-7=���%�P����
t<h�g�P-'�>d�#FȉB$j(@��'�*7� C�'	�Ov)����b�����O�)i�Qzt"O�psc�[�U\J����6IgDQ�c�d\ɦ���FyR�J1@�H6��O2�$ˆ=R`jW�u�Ir旁2��$�O�9�g�Od�dl>%��䑞T�ء�]}�n'q�`�c	[��3�#�p<I�.�>V`��0�����'/*��D���"�B5v�L�Ǔt�u�	��@�'߈�X5F4>~��
�	L�i?`%�'�r�'��O>mC�A)��jDm_*i
�Q`"�&����4#E�=S���'4��F�K4f�Y���k�|�mПX�	T�D�D�K�U�L�Z8�RDμt�D|�U߬	���'Tb|2�,ɷH�<M�r�Yx��8{Aã~".�LjR�'>��\@t�D��N�"��>��OD5z0�&�|MXY�����O	���ɰ8�N`y����u��EKJ������O@�D�\��k�S���eJ�?J��R!ɐ[U*��?������'o��"8@������)j5h�Ó'��x��OR�a%�X/x�|$�%�P%$�RIZA�ݦ1��ӟ��	�H��c���$����p�i�	)��ŕMN��R	d��"şfXH�7G�1+��Q��&*rf�|�>�'"��#�Νe6�e�����y�#�B� R8�i�jQ2i�?1Q�S�M�-v��z��=$L�mسC�1�EZ�+k�f�<ٰ ���>�$�OB�D�I�~eif*� ���	��A�r��C�Ʌi����#j��^DA TA�f�2�	��D���"���<ɲ�^>">� �"�X�İ��+�9]��B6����?9��?Q�#�.�O��y>M��ת"��҂N� b�pH�ű־C�	�v��q�&��R��Q���L�B�z����3��y�F�d�(�RK�N\���D�S(XW����O����O0˓��󄙾`�2�m�/B�PRg!�>H!��Ē@�ڙ��I�������V]1O�8�'��I�6HV�y޴�?)�A�x�c�,
<XSt,��.�s�,�{��?!"!�1�?Q������D&fH���j]�B��		K>ذ�AJ�5s*=9�lҩU���䐛�>X��ƌ/Ȫ�(�-G
ݫB� �3�c� =;�u���)u����Od˓K"����yx�-c6.@2a�|-��?������&�0�̬�~����0k��{�O�%o�r;"ͳ�i�Q�DP`������Iry�
x<6�Ot�$�|B6�S��?�Ul�!�2k!��U�X��?��.]�����D�a��Z�ʧ���&�t4چ�؉D!�ՠ��e�5d�k��I���l�����-xs(Lk�lؐ}��1`���-c�� ��a���M�U�i2�i C��;'�̮c�B�Y����d�O��D�5�4���͜ Ѷ)��E��d7آ=ͧN2���2��	S �����5ю �|�F���O��X0�X!"L�O����O������I���#Ą��E�4Y 0(�MU���!V� B��q�g�	"N"��BW���	iǅπf����x����S��}&��iB��/1���XǢ��6#����T��M;�i12��C��,O����23�rESf��?4�v����a��C�I-hS��r�A��3���HJR��z�����O��I3,��M�&�Mvl�as�	jN|L*p�Ԕ�T��Ο�����<ڮ�n��h>Yy�l�#��*� ^!U#��T�Ӳ<��1��Kh�36 X�~������o.�X5啊J)��y�©t�J��ЂEPB��bP�u��K�ɚ�\�-�G���'���� =5� a�w��8�%J���?����?�����D�O"��j&��"�2=�UP���` D�hb��Gg�bkG]�2:�t{�o<�	'�M�����@� m�O�B�[�(̮Q���9>3��Ts$��'�����':B4�$�����/t���[�A6h�CN���7I�,:_`����M� �F~b�Ȧu�Q�a큟}ꑐT枘$�t	�t��c���`��ua�H�Oרtd<,�E*QQܓ1�]�	��M#W�<zU�!-��qM�1&�X��&�"��r���s�@�2���F@ԜhfDPXd� �8�ݴ h�i
�"	6��L�$�Q�<�?����9O��k�h�#T	A
��+&\`)�"O��`��+�4��X
?X$1��"OT\3ƯIZ��* $)�� "O� t��3)_�9Vm��l�)>���@"O�l�hDV�5�2�;X*xER�"O�}���t�څB���.O�����"O�$�ÍN�;�*���
�|u��v"O�}X!G�!6�8��;PBt���"O��he%��p:vt����#Q�ѳ"O����ϥ^��M �YWf�"O��ы�{��T�$�[�%F��"O��ɀ�=x\�	b"U���� "O�Ժ�KO-������L0!"OT�6�E<ie��c��V�pې`�"O|�*�Ǩ\���I��R?%����"O��X��ߦ$V � �>I��|�"Ot�+ BH�oZ�{�g�wæ	��"O`�P�"I~p�hb�$$�21��"O��T�Q�\�����!����"Op�E�Ϫ�2I��Y�3A�A#�"OT4YÄ��a��%4A���"O�ܸP��-�ȑZ�OV,-����"O`)�/�.C��=P$���_�Z�h�"O� +4�7I��HIïW�֝A�"O����ϊ�V�`��c�,u����"Oά2a!����X��Үi�	� "O5��і/���Zbc�G>���2"O6P�-ڶq� ��Ed/r)ӕ"OR�Q�H�a�n����ˍ9�E��"O��#�J[��b��Eƕ53���B"O�0�
�y9���� a�P+$"O0�j��@��`s%��Z��s�S��* �7�b��1G���S��	Ɵ�aq�޹|��m�3�� ~�A�׫5?�Boq���p�Gv���9��V�'f��JBmZ0
}�	Z碑-MS��(e�;i�p����?	Ӧ)
E��Pr�
ؿ���`-�-��R�'(��Ey��_T��d%s��q�L�1q�5&�����ʶ�2�8I"k3 �^DX#��1#4qG	P*e��O�P �BI�ML�Qyi��:Fp��d�x�[MXxbPf�6J�N"!��6��'玑�GS������-��9BN�-��!8g�G#M�  ���Y�̅k��W�~5�0i�`!�Q�L�fq*�F~򯉖9_�H�r�Y�m	s(/9������T}�`[�Yx�3�oE�O��u�Ĥ�,��'Q�m�&Ժ��$)2h��E�ر��-�mCV�[ud�����H�@�E�@a��2�&�Bs���.d
P�
� m��#=�;F��� ��cޕ�a!LƂ�Z�i�2ʜk�Ǿ�`s�(ݠh����TCy��Tn�����T�_3��e
 S�g>X�i�}��/�ڹ`�B�?M`���!H ��B=� �DD�+:$�Y{��"�W��$:B9|e1 ޟ���fM߰`	���#�!0z��k���#eMT�Z�ҝ��W�c8vP�'PVD��! ͹�z"=�ק�#8s8� 7`��>��&K�Cn��$�.VKVlS�{�d�cp���ـE��b٪m�*|���dM#z��TŁO#4e��(�/ ���Gy"bU-L�����kk�e��?��-��K���\+6��!�/��z-�D	!�7�2�e����#�'���y�����RC��<�iC�ë�?��놻}��0��Z�d��{����"\��5,�&�eɗp�:��AB���`R�芘F���4�O�e��L%�pQ`��+xj�B�+AI�b��uAf���+t��P 8Re��5|�\�����@@��(����@�ܡ���WQ 1k��ӎZ"pѹ���-�z�!
�6�:�!
}�'"���@��	��1�FJ��"�"f$ک3�6��G%$�x�/�	"Ƣ�8�aS�Hap9rPJR�w|"⟘�E%-l|�ɱfc�!dI0�r�˙	��81��S<~�hh����c�`�O����3��E"��36Q��� )O��m2�K`�Q����:s�6P��wL�xb�B�	��YQǇ7o�=��l�t���75=�X�dգ����y`A	�y��ej1�A9��������'st�A"d	��@���ܟ�N<p܀�.1���	m�@�5��  7��� Hʒ��-������?1HB�T��l���=0�D�H
�P��P���i��"2JQ~��
�Y-5�Db�e�7@������M�Ch����x�\#LJ����Ň}��PQu.�P�H5��4b��1j*΄��&X�MEx��ԲP{ļ3��@�R�p�Xe��>*H,	1O�9'�4ku	G����ɂ0�D�2��H�r��iޙ�-���z-V��:�"!ƉmӠ�qp+@��p<��L�DX��v�AN�5��3�E�ӄth�'� ��C���dǑ_dd|У�>�MC�hj�q�C@%e�r�!І?e��=rA 3�B��#��<�����E������c% F+;�ʠ���ԛ�6��'���CՉŹ[��$<,Ŗ'g^m��!O�@����V���)n�
(���k��q�����D�5D�0�GN	LW�e����~If��  �P���O^dyau��:e6�"�O4|�&�Ky"L����G{��ƙ"gz��)`<d5�2�B
�n�+�.ТuιB�CF�lS*���s��<ͻ�¨�D���@�f���iR�\�IlZ8uht��'r�x$E��X� �ǂo�Ճх�p�pQ3GÕ�O���N}�ͽ>Y��R�>���␎,jfh�̻#]tH�saχ�L��L��`b�Dzkֱn����'A�hT]�]Ϫ�Ҧk�����S4�������v�M������s\�H�5�� �z�[��p{&I�O�)h�ٴy���#D�f�X���'��LY����8B�E-�䈘x�D�c*OJ$��D�8p��)��z�pqq��F��C#D�Oذ�2��IS���E�6/�5��&��֤��^5j���ai��Y!-�*Q�,OP,0�� b��i�i+pa��H5�����8���#��&�O�@V���[Z
]Z�bJ�)�x:��F������鈄�?٬Oe�Te�JO��IRW�닏�<���QR.Z$��UXu"ϸB���S@?Y����L�^�����4?��+ai>h�6k�8�6�����8;'�D�>�/�	/���BH�OZ��X3�׏	q"���߫&.�*qe�^�H��9g�����P�R� ��D�A�Z�1tnX+��O��V�`��W�N�7k�u��e�K�hPp��ym�z��H7������%GXp����_��(O聡`�Q�^tK�ņ8o�N=�V�p�L�t�'�NTDŇ:�ħH�A�	�"pV(��$,����
4!�+o5���@�6�����%h"ZD���-p6nБ� ��PD{����/G(����T�X���*�ƅ���iz�J&�P���!ω61z�CQn�+�X�'��X �S����-��-�Ҩ(OL�,��b�)7zzM����65�� �T��"F}�E�C�k�J��C�d��Ib�M�z�X����!8�d�C���D�����y�hl"c-��ol��1 �<�剕־�+bcԠlrHi��M�Zȣ<i��VS�E�4�U�BV����e�Ojt'����m6�Ӽ�DH�$V�M*@�����U�lȑ�CfMɄB$�>Y�%O5pL���;L2���õu��Hȵ�� �h��,#�~0]%�h�;8P�PC(F0X�3�,�0<HEx"��'i�<����n?1�$�P~e�PV�x)s	W�R�X=� j�����%�' ����'?X<�b�!��(1�K:*��%bD�U<D��S�c��!ĩ���F�o���O��%�ם��Dԛs��"�i?L���E�;��	�d00˓7� �xw��HO괊�?2��m��$ġSr3$�$ԁ\�r1 �^�X��!���ګ)|}�r,�XN1�s�($��|�`�)@"����i�V!!���f�z0��V#F����a2"HQ����&d�zC�n�Aے����R4|I �{�*,7��@��֠o�$#��O �y���lه(ԄDu{tJ�@��s��4}���J�I�I	���#?���q��Ķ=B�B�j��
}�(jf�� Ѽ�q�D-i�ԯ��&���׬s��'���J��A0��
�t��f�HGv�↰<ѱC�{?)��s�FԁV	%�G�B���Ȏ_"dR��ک~�|�s@%DI�ɉ>|�>ͻr�����̗<�4�ĩ�,9S�+#�n@�}��F3�j̐7�ؼ���|�sW͇�]N���џ�'64�2��G�~���ط��M��. �
Fl�D��2<����6��bԘ��M \���(�
v�x9�'�T=�1�IZ��i'�L�N��H��'�0�su
�b8Ź���aLn\��FœX��*���z�.�NJz�d�Q�J`�)t	ف'j 렬�>��'��I�J:uI@�O7kI��˲iW	f�C �R� ,�t����lv��dn�D�*T��^W�'8��Pi`�4�����,(��π��'��	d��2��ޱ4P�t�a�,����Ȉ:N��I�_'.�6Aˎ�D������1︡��F�'�dt�C)I�C�(ae�'��	NA
=��@��"|���-v�8����53ذp�G�
@-*���U�PpR#L_+�`�4H�U �	�.����� �pG?^5��'���y�h�H��G48)@!/ПD���C�F�4�5x���;���
�!D?�� ʒ-լ*����"�� �Be�w"�lYR̨��$�>a�ӚoGJ5�A&�3�V�*s-A�9� ����UY�=�aՈrW��¸+�ZGzBꅮ1�N5��E���IB�ڻ$^�W�D�Y���c复�a䮼�'vU�#�����4�0��G��򔄒���F^.,s&�'�.-q":Oz�wďO��sV��8���F�����X?�[0V�����"0N�i�:+��n-Y�,��JP#E���S/�6�������4�剣6����O�(P��ghĉI���G��8�+�@}"F\�v&R���\i)K�	�Syb@2#Tr��ɬ+x�s���$����&>^<6m<.2�/O6���i�uy���"c7��')n�[&ND�D�B�ȴ��q��'��$J�<�p+խ1KĢ=����%���j��N�jpP­K�K�h�YR����I��O�./����B�'4�V�CР8l���2�R)��	�F���b�'�d@�"c��v���X5F�E��ET}2Fȉ'����`�<i�o�Q��ݠ>�V��w���Ix�)��(�B�f�<A�CI'p㰺inj�а��@bƙ ̎��^h��Oč1�}yR뗦E�x�/�м�6��Oz
�KG�a�V`�f��jy�&�iap�6��JyRÃY���!+�O1K���a}"��8l��%W�0��2�A7/�Z��4�O�;�@�iy�a�-��D{
� ���%)0V\��U+@5�D`�/�!!��Tٟ$R��X$���|��y�j�2R�P�д.T<�$�YA�E�M[B�
�]�"?Q�A�UX�bn��h��G��=��
�j,-��D��ɾR���$�$��4����b߸(!,RD�ܴdpX��$$Y��qX���=c�����2S�'G��&��;�ܤ���ՑE�t�a�Oи�?)4�'��)jql���b芐W��!r���J�7Ȑ�i¼C"�>\��°�`@Z�t�Q�4�'Z2�������5���C9O7�zH�\i��ϧ2n�Q�H[�2p P��%�I�d���4�|���X��=Π�K��*�Sz�*O*)�)�f/T�;�L �P�'-�v�2+vB亏��O[L�@ټ�׉U:@H�u.��G�f|۶џ�F{��)��S�8i�F.�!!z.U�E�Þ)�K�}�o��:D���
�l��Pi����:uC�@�2>:���#��N�
�'KQ�$���ߧ�0�
�×9T��Ѕ��d��ԉT득7��|�Um����H��]�5>�{W��'U6�DyR�����!Yj�|F+ÿS����p5}�F�?'d8����_���# Cݲ��' ��ڰ�
UX���&&"��b
<��hO�靹VVtXz�`0���2H�}|ޘiaM��'�Ʊ��0��?��6X�=��nP4G�ְ�qF�@d�t�%�X���$�& ұ���ױ@<��V&�Tx0��}��5^��J�7Gz� .K��ē���h��>�}K��'D9�Ї�	�I"����%�;8�ZFg�-` [?�8���ڞc�n�9��F���Ϡp4|��[䎬s�S��LR���,h��`�@����'��9�CɈ�x��(Pg�	���!��$�jeI0�HJ�BH�$e�1 ����T�"��]�Pؤ�	:7��c$�OZ"��YL(mP��{���!d1���#f�Hx$�O�2FX��Ɗѷ�
B�	� �� E�T�^�s���8	���S�$^"r��US 1t�PpyE�վcX�'��Y���Cz�څbgG�j��d��O��@i��=UǨ��AJ!�����2�$����U�)��XS��[�~�,!q4DRl�\d�6 ��<�W]&XF�q�%#ʒKZ��Q�^v�DV�e�)!���,t��� �.:�OB�	V��'?ڙ��垞_��)�,�|ܓoo�iZwA�#~��h�C�8H��B�c�� �8�@�4���.5;�����E��y7�[�:�<9��##6VE+��#�t�w�޳c��V��C�ø�M�'RK<�K�O�q�~�"�Ԅa��q�,�q$&�w ��:�^QppE�ȓ+�R
q�A�y��x�����E~�����7o0.�ՠ4�ܕo�h�'W��P �	{v� TG�-e�ΙP�'�V��G�$�"h�  Ć���*�'Ò	��8S*�����!j�'��&���UVj�r`�����lr���6�	*�XZ��7�����AQ i�'*�]�����F2��ȓ���cvf*�0�	DoW$���(	�(�-��J�P����B��ȓ8��Qe���g��A$G/ �ȓjG���QG�����捗!���3�="A�ͫS�:I�򌝷D�T��B�IƠ
�q���G� �Y4r��ȓ6�)D���	��+d ��	6���ȓ@t���Ŏ<d	���Z
�U��;�faK��9`�0�Q`��7U� ��g����s��$��1�� �$}�ȓ�40����˼�se�'I�B��ȓ��E���˜rA\9J��;~�D��D� �!�ڈ�:R���!8�h�ȓ$�pi�OG�+er�Y�K��G%�T�ȓL~�"�퟈
�4����_�,i���I��}�0�_o��y��˼\����4M�5��9��@����+�bM��h'8���$��`5�R'< ����8�c�LH�GM<���j��o��Ȇȓ�d��ƕ30$̀u�$O_�ȓ#�Ф@f��u���@�ͼJ(�ȅȓ ���I�G�B����i�;Z<\t��Q;�M�3�S�w��ӯ� "Wn ��S�? :� W� (���/�	���Y�"O�2�׾g�|�p��L㬕�"O@б+�!��d`V/��U�D(�1"O\P 3
��7S�[�j�YY "O=�G��D��u��Bo꙱�"O�*�G׳E�p�F�6���1"O�#��T5D������Od�ti�"O:,*v�Zc�x�Z�#W�-�V�{U"O�Lzb�6c	ly��AK���H�2"Oj���CJ�JzrB�'�`�"v �G�<dV�2>��FOT#��`R�A@�<��*�!�ڄ�Q�fxJ�*a�U~�<�����3 (EB KN�T�p�<I�hܶ\<0����j洡��R�<�*Ch�L����r��%
E�b�<I�N��4���Z�`�A�`�<����&�T�sqeщw�����B�<�@����iЗ!��`�ʱp3e�~�<�QBq3j���!�B�L\ �(�P�<Y�a�;N#�s+	���q��u�<����6�x�C P�+pio�<�A"�f���R6�N5&�-ʄ�n�<)���^��!�fN5֖A����k�<!��O/<Ѻ��S�z�څ�Cc�^�<q��?eN�r�Ꝼ�a�g�W�<皃[x`śD$��juR8Ч�U�<1� �$:�caޓ)oB���o�l�<�Ѫ�5z�����g,��ps��O�<9�⛛GV�遥@PVk�mWa�<��d�M/J
f�ݺ):d���ȗx�<��O3(�Hj���}�J��f�	t�<�7�ȭE�
���憍dN����$�q�<i���:�6E�W�C�wt����'B�<a��X�rv��P�Iݚ@aVL#`��~�<���'^�8)'�W,W�H��c�I{�<���R�E^(��e��!�����m�<��j�e�Tp��CK���e�c�<�ߢT�8����ۓvl�0��_�<�j���u�f�x�XD�0Jݟ�1�)ڧ.���z���!�0��TM��9E,��oo�I��W�4>(]`(�$�=��V�`R���JԪ�90D^"�|��ȓL����L�a5D+c�[�^�B��ȓAu
%ё���+�(ɚ���3]i��p� ,���AX�A�qv 	��$2��w�H^9D}���BAUͅ�T/VA��<j�~@���lr̩��*� �-�$|P�t�%�f�d1��&T�� ͼoF�ȗ՜B��A�ȓ1f1`�׍E����/�k���0u�=B� 4�t�k�B�^��P��`�Ƙ	Ԫ��G,4,*ƢO�v@�ȓ(/�!�0��Db>�1@�

nH��?�
�	QP�� (�(4ɮ5r+�f��ȓu�(1bw� CM�}��I�Fb:���S����
�*�x-:5���
M��	�������,�8с�U3�ąȓb�L��ë�,��ȶ�җ_rI�ȓ3�,�%N��Cu�}PR�V	Jjm��m�*���$��zY�5�UT����ȓ
~ �Q��>ew����A�$��@�ȓu^�]�ض��E�&��({�<�񠌅Kv�;F�?�����^�<������̅0�kɹ* i�a[�<�  Q�#�Da�F�#D�<cG\Y`"OV�s��-:���KL;.g��"O8����߁Vw�M8Š�l��y`E"O� ȤNޮ�q஍�%��I�7"OL����X	�Ջd<S��x@4"OBAkbEI�s`�QYR�A�Zy��"O8D���)e��6c�v�p"O�����p�
���S�X���t"Ob�`�dE.1^���g]M��R�"O� ��/T�~~>����<E��"OYt���:P��Xg^'5� ��s"OV�{�j=<�� �E�cqȰ��"Oz@���N�ʁZde�Lo�]yc"O|0�+�-��@�dS0�x��B"O�@Ō�2I(|D[5
��0�hh�7"O��hӧ�j��J�\�����"O^2������S��?�^��"O����G�>,���ˈ�T���"O���@�Ӗ#���3țf�fCP"O��� w�Ή�!B�+)���!"O�`��H�t_���	�Z���F"O�a�Ŋ�l5�Nǡu�fa��"O�U��F�GjX`]0��e�2�'G�(�d�����W�\�{�|(H H��^!���$tl`��L>�� �%V�k!��C�M��P0�� �T�e/��+!�D�6��y#����u(�L����Q�!�D�fm�Q�ޝM���q�/�2x�!��ҰS��=�0C��X������-!����i��1�>��W�ø4!�[�.�4ڒܹ�H����a�!��	'6�f�Q��z���fU�!��	}���nX�"�h�PƘ�]!�dڠnXp)���G�l����+2G!�$�/n�6�R�b�|���C��A@!� `h<�0�m�#V��<�"�@[��L����X�M޾q�T|9[�>%!�����y"���Fr��h΋O�N��#�D�NB��3=�d
�̆�*�3e�?%���$	H�2+�Y� ��Tْ�AB�ۂ?�F�m�c}r�$<�I�8��ّ\�%�� �� �������ox�q*�KX���d��y��r�� 9Zp
���,��Y�ȓ!�.��OR�D��#��Ѭ|&�̇ȓ4��Qs��&T�6y��%�)`�,�ȓm�R$���&|���Fj�(H�Ā�ȓ_��+6!����V w䤆ȓ��Ԃ&b�(Aƀ�t�Çv"r���z�n��1o�����J�C(l�ȓ�h���0R�b U>����	K�6W��B, ��>���]�d�.|E}���/��بT��2i�~th@.�19�B�3	+�ش\�<%:�`�A��m�
�'|B���F�-���*��� ;�!
�'! �#�Nؽ��љc�4';��A	�'�n�1��K>N���k�(n���	�'X¡1f�P�M�b���x�����'�&�u�LrI,�p/ys4eX�'�Ԑ������b�qM����':p�Re��k�j$�O�bt:$��'ْu���qئ`A%�9ll�D�޴�hO?7�^1. �RV�Og�f����(O�!��W�f�5+ÁZ�#��h-
�[�!��V+D�e�@�9Y��tAu�M�i!!�� r��*�5ra��MC6R�T��@"O���+Z��V�r��ߡ�� u"O�z�H��Ij(���aX�ݰ8sW"O�23�;3�ޜ+��J��6Y23Oj����6zbܐ����=��(�r+Q1�~�U�L��ޅNDܼ�TIʹ&E@�ۆ�&D�@
��O�S�0��D�A\.�zV"&D����_��=�Pȇ9^q���?D�������İ�#����F(2ړ�0<�P���6�x�Q�&*��-k��Ax�<��a�,0ïM�Bd(�(P�<�*C�5.IXc�T�'kژ��mWM�<��\9����2.E;0���&�<	Q�يt4�P���٬ҀL�ѣ�a8��&���@�W8��z�V��DQS�;D����E/Vm���b`��_k�p�%(8ғ�hO�{
�e�c+h�l��c
)�pC�	:j�|eh􈝋-��c'II�`�B�I�}xrXr��\t�p�!c�y�aE{��9O��+ �	cJ<ɠ�<�@�ː"O��T����!���N	k���"O�)�HJd�|͸1*6!����"Oh=SŃ��T�´kqb�0�\�""O�qH��4�8PB�9\)> ���n����W\C��Q�*���0EAE!���|��pQI�IRq��)v!�ĕ"r]+Oخ=���t���!�$<��M��D�4?�.#��K2H���O��(��9dE 3�҅wHV�ZJʵ�t�	}�O�u�d����%X9F�,`�'-l�ن
��鬥�C��3.9:�����'���i5�Ɔ*p��:`�J)r7���'��Xy�cقxZ@����z����'���H��j�K)B6B5��A�'���� bTz#�i��"K7+&L1	�'l��S�`�� � �.�dj�'YrԈ�--}��c����4�8�'�r-�J�u�� 3b�,$+�'�j���h\�/4L�"2,��T��
�'��	��Fѻ趌��L��L,�
�'R}b�]�6w�p��r�ܭ
�'�2����ab�hG���mNd��
�'��p0g�ߠ.����a�g̜p
�'LT�#h6kw$I�m�2H�2Y��'r����N�)��0��-[�wr�0�'?�h!��%v!xd q�}HL��'v��R��f-R�P��\�k�.��'{b�&kߓW�51E�f&<j�'�Tɻ���#��H�D�Ө)��D	�';�����ª�@<�H� Y�	�'G�	����.i��ЬH�<��0��'þ�2����6;�0Q`�ĕ,2�k��U�K�w�H�j����E�?D�Y5�
&X�i���K��)0D�`36=�Z�af�4>!��3�/D����A
.��6ˁ��v ��L+D���5�6�ҵ�+ob���)D�䪥b�$��h��i4ȸ7M3D�`�Q�'b<�q���"����t"7D� +2`��C�<]"��8M�ĝs7�/D��2� ��1 �v�ȝ|�!)2f;D���SJ(��Ĳ�`m�F!(�7D�,�Eǒ��`8���E;
�9C�5D����BY�7�t�j�)�R@��b	2D�� �t�Q-,7"eq���/���$"O� scT�Y���4$�X��z"O��+q�(.�E٥��(Jl��"O��IB�@�j4��K��V�4�z�"O��{�a3�.�rsDؽXH��"O�qJR��$
2�9 ��#����F"O2����<Q���3B��	rn�Sq"O�qg�^��4+��7a�uV"O>��Հ�3�A��	y�B"O굢v�Q.~�f�C'$��H9�"Ol�9��Q��Y���JE��х"O$ԙ@��$��=�N��y5ZԚ"Or� É�|�~0�W�O0 L��"O�lj�Д'�2��E���?q��8 "OY�ħ��6H}�Q�B!/o���"O�B��[�\�6����fTE�#"OP�)Pl�^Ў�hΒUI�,�"O���va�R�n\��"��	<��c"O�jr�J*J��bF�1���"O�ӧa��.�b��\#�}�D"O�IA���t�V�/N��a"O�(���Op!:�:�ȫ4�=�"O ��Rh>"��0��8�cU"O�XVX�^��A.^�v����"Oj�@ܕ��pzQ&�]� A�"O���1�?m�$��
�#^M{�"OX9�������H�3Xj�"O^���¢��P��DE��YA'"Oҽ���?U̬�e�TLʱ�"O�0��G�T*	@c�)S��u��"O��[�,�,��r�ƦR�h���"O2���!B�� �"e�J���y�n �K)�I	pf�����*�y2-*
���ԊJ��Ty��D��y2��0x���)��d%��EӺ�yR�ۓBf|pZЎ������d����y�b��\n�V�@A�����OR��y"�ԭ
Y�|�u�V�=�V��o�y2$�%��`	��ý0@�=�2�)�y���l� �rI�<�J� W��yb��>���o�>D�d�*����y��
�*���Y4��9�����y,�۲�S��(e��V΂��yB��3,�I�$J�P�QEe��yB�M�g7X��#�/bp��T㟮�y�O�o�ܽ9b�H�lu^8�+���y�ߖ+1�r���]��[��y�"˧#�<q+c�\ |�����yHӑ�Tk���?ɸ�����y��R#x����ƍ�b�n���y"k߱f|��" {>�-�%a-�y�kW�Z�0�,�{�����['�y��Wln�2��>x��<ps	��yBG�)s+��>`��)���όu�$B��!BV M�0��@����[��C�.h:4q���E��[!�H�|v�C䉿A;x�)4mսqbj�kR�?��B�	�l/&)3&�_#�\1���Ƶ<��B��!>����&`Ak�:�(w!�#R��B�iE��(O�R�*���aȌ#|���'��d�o,C���p�!N�&b\��'E��I�J��ZF,����(ҚiS�'-���E_"�̈���3,x�'^a�O� �*�;ъX�>������� �-{v)��~�h�#���$zw>|��"Op��t�U�U�.<A�a��Dh����"Of@i�M�*1�n��ҩ��p���Qd"OZlٖÜ�Ht�](g��r45x6"O`h(�I��:���
p뚉!�<��`"O^�ѡ�Y#��f��.�XrT"Of�0h�=�
]C��ɠ~�DPr"OZ�(�(_�_k�@CA&�R��9�y"阿��L���$s�qi$��8�y���3V��c`�%�"����
�yBFS�{��{�Ԓ}IXQáP��yB�ڀq2�l��$^4w3��!�S��yrĞ�L��!$#PdL����e�$�y�	�:X��y4`Q�̐�y�U�&s���wN�0��[a�;�y�.47P1�žt�4�hU���y¬�4`�bA��#��@c����y��Sx��a��G2Έh����y"0I�Z��C,��`'̘*�y�`ݵq7d8S�k�
:&�qd�V�y2�E��E�
��1���fI��y�(R
O��@���wJ �7���y"�5� =1�P��玽�y�9\Ǻ�f�
�]�����Ȕ�y�/�$s,Z%�0��Kc��"�ybǞ�sbDc�DT2	���i���&�y"�V-V�{���Tl�(�V���y���(��c.4E��bB��y��F2%���kd��∩#1�ל�yr �=�E��E�^"�@0�&�y�l�29��A0@ʜ)@ͳ7�]��y)�5w�~�g�S�Th�tA�n���y��׈��q 
u���S`L��y�e�O�]xw��m�Z��#J��yR�ם;��+BA�k�;G"�'�yb��Ca�p�'��)v���ԁ�y��U�hd���f�P��󇊪�y���"z3�PC� K�LD=9$�͢�y��U�oѠTj"��vTm�F%ǟ�y��$��� �-~u
,	���y2�M
�q���<q�a"1hA��yRƞ1�0l;c��ph���[��yR��	z訠KA,Z���;d���y��_�V ��"�Jh��z� ȥ�y�O
��`P{4FK'<�W�	��y��W=�|��AфvNŹ�D*�y��E(d��̅�t�@e*�fU��yM˽X'V3��کe������޸�y��L�qY�X��^gPx���y�5t�$ @�\�J(�w�۸�y��7wma��c3Sk�0�g��yr������$��N�xP�����y�*K�K���cwl>��KJ��yBG�T;���D�""��1���yR���KEF��u�丗�@�yBlǄN�V�T����ث�$V�ybc�#���f���w`*��'�)�y�E� ^�֭�7��1nq�Z�B@�y�ER<= ���@�g��@œ�y��U�A���t�-t��\�$���y��8 c��Ҩۼ{˞��4'C�y��|¢�q����%2=��¼�yR+��#ZhY5��+-ཻ�)W1�yB*Z�k@�c�M�O���D*�y
� �aأ�7 <]!t�0L���J!"O�� 0o���������x�<hY�"OH�ە�
O��LO�2�q�d"O
��CA��<��e��*Ǘ2H>���"Oh{cn�kO�,(p�֑TA�l��"O��`��F&mZ�K@m�"%.л&"O�а�i� '��)I��U�A���U"O�8!$I)ϔ�Q��ǽ���"O~d	w�'�T����#��x��"Or��Ö́,���3o��g�4M�3"O lr,Q�-�Lz�O²q�^y¤"O$��直0T��9@���2"O���a<?�6�{$�>&��p�"O�F C=k&�;�C�-�r��D"O^�W-��J��=Q�ǐ4�L� �"O��B`�M�
�X䓐�_<j��[�"OB�pc	�_���Z¡R*q~���"O��I[Y�(<���խ��\�Ru�<�A� ���C�&E�,l�ٵ�Ok�<�dl�3��cF�*�|�� J\�<���@�Sz���I)N9H&G�T�<Y f� �V��1��*�mu�<q� ��LZgA�%
� �t�<��M\Z�=٧fݏ��j�J�r�<Q6!G#kr����2ܤ��jEr�<�&IT
u+l�T��/ʺ��t�I�<1c��1?d���k��MP��W{�<��e\�Q�.丠C\9��J��t�<a�A�p�H	��F�Y|� ����u�<�2ʎ�G�t��Fӕn�`�S�]p�<�Hк
>��J4m�b��3���s�<�#U�_`�a��P;g�8I;�A�o�<���@�R�x�P#�ԝ0k�l ��b�<̚�Wt�@bd-{N�8�`_v�<�$Et2����xJ`蘢hZp�<�a406<ܨ��ڗ.��Qk�a�o�<����h°�C3g��6<�tE�m�<�$O��m�����!E�;˴�2��Rk�<�a-��,b���s��O���!�g�<%&Y�w����ǰ_��P��Io�<كE�R�|�Qn]5Y�D�᳋�j�<�4�|�d�+c#�.���J�l�e�<�4��=O(�5�2��-$5:E����V�<�Dg�+E{\P�$%'*���xn�P�<��/S�K���Z#M
:�V}x��S�<��H/��:⍆!���uL�T�<)2b?)*�,�$`���� 1v��R�<Aub��o�E)��H<g��Ѓ��z�<�ӉҪ������5'��(U��{�<q�GB4K}H��gP]d�9�!Go�<�q�*-v37c��b�ĽS@bd�<�M�24��ĉ�i�!Z*����b�<�b��&D�����G�m��9�iF�<!%%3\�w�a#��Z�`�B�<��$�6l��&9�eZ���A�<9˔6p�h�bF��W�Ĉ"��z�<y�G�>a4`�[� �!|M܍�d�E^�<)sZ�`�i��W!S�N��Sf�C�<��(�K�65ٱ�Z3�I)�L	v�<I�
_�(:@Kҗ�����Po�<Q�hT�u,�8#B��d�wHF�<��-�6x͒-�!��6fP��%(H�<��j��vP�ȁ
���P��FG�<Qro�$㚠�jגS<2����@�<� �{��R�x��9 "�ي{s��"O.�P�ަ��qgL�Fsn\@"O�0��r�<<����,&j�0rC"O����Z�SxP���mR�s���"OVC�*�),'d�� LP>��*"OИ
WKj���+" C�o���"OT$;���;F`:�.
�E^��s�"O���#��{h�I`�-A(j�;S"O��0V�R�:��mP	s %��"Ofq���U*.�fM�P,�ff�D)�"O���g(<x��1�E�_Wh��"O^��p���|��j���9��p��"O�D
0�Eb�x|2F!H��,ɒ�"O��(ˏ)�@� ���N���"O����`�
F`��OY:�� ��"O�i���;$>��o���(�t"ON����)S����CUɊݘ�"O��j����a.$E�a�C!5�"O��)�B��%��b��2!��(0"O<���*ɘ� �YVo��Xq�0"O�,i��޵w,���ؓ�عp"O�}xv��5*X���Ί� �>��6"OL3��[�A$fE�"G����AF"O�I�#���*��Ap&lz��Q�"O@���c֐����*K/��ܲe"O�K%(���r�Ęji �s�"Oj03@&[9/��X(��zE�"O��3��88���sĊ�	���"O&���P.Y��)�0JT�q�v�T"Or��T)V�Y�Pl�a�X�[���#�'P���!8����F�75����'p��$n���(�aĢ*��Mr�'=Ha+R� �����]�1��'0>�Zs��yL(��@��a�ΕC�'~0-b4c�
 f�����6H��r�'v�)��P@�����<<_��;�'���:'��N��p��C0:b�r�'�bUA�P����O�-�LP�
�'���M��a��%�P��3� �Q
�'�� ʦ%�0%$Z�Ϟ7A�M8	�'�4]���@d���e�1LƁb�'0m�Hw����R�:Ι�
�'{Fh k	H�	��k���
�'���Dj�4b��(�wǋ�܄)	�'p�٨� �+�v ��*ϔmZ>���'\�x��N�5��d��a��x�'>P�	G�K!0�$ȹ�ȱR%,I3�'�>@at�y�B큠�H�M�2�',�tF�TN���+�	B2|� ��'��Y�r兑�0�-��6���'U�1�&jX�.80��v�Q�
����'��E#n�G؀�E�L�9͢�Y�'�ty����vH����&��0��q	�'p�4�uJ�%E��+�����a��'���@�ʗ�A�X�zT��?dh��'��(�G#L��R�Ha��!]��բ�'��S6�Φ.d� ���,����	�'bnDX	��٨'��&4*�x	�'�J�)�M�2	���\�պ�-S��yb�X+?�����˝�7��µ�$�yrF�K/Љ�`�ԙU����yBG�/i<�i�G��u�������yji�Ō���M�$���y���*+�rx��d��pag�y
� �x���0 H���w��k�"O�MIp�Fj�P���@hh䱩!"OT�k�vWh����0a��V"O48����8G�����'5E��ʱ"O<Yg�^�V�T����Q��l	@"O�Q����i�x���ف8�R� "OlQy�	�� ] �'���R|rD"O���#� �|ꣃ�&҈�v"OdLYS�=?���`aE �Ԙ�"OZ,x!�U��eoE�l f9�"O$��E
�1:��:3�X*p�#�"O�9�C22\�M�2�+(ʹ9!"O��g�M<x�k3kE�A>օɱ"O��)���:[2a��*E.4�8�"O܄��T�I�2�/�,�8p(�m�!�dٺ&_���H �|��y��)H�!��J�T��D�F�	v�H�fV!���g�1öJYl��8Xņ�E!��D�T�,5��"K��i�&�e�!�,u�e�PC��w�@�3G��X�!�$�LӮ��C�� ��)b�O�!��יR�bD����$P��C[v%!�d��� ��Rv6�T���ƺ
�!��_�0�`lC$d�6{�ZRb�>i���0.��+O��1a]��y�E��<�����h�|����y��d!�<�f�G?XO|�k�$Q��y�鍿rʸ�� �:L�Z40C�D�yb�'l���#��x��!�qj���y�fK�5Ƚ裃M�p��X�M��y�.�c�Y0���V�0܁��!�y"�8��p��ǒ#cZf����Ż�y�U/j(���[Q���I�3�y"�Y�j]����Y>��P�*��yR��R؀��B��R;��p��yB×3zR� ��>4�A0 ���y�gԥa+ t��K�:�f�0�e@�yRo2?c�z��У"�|�Gf4�y��� A�p���o�4k�_��y.�JiZU	�@эgb	k�a��y��]>����'[�uv��Q��8�y���M:�����i��y�BE%�yr� G� �f�$����yr�Ѳr�X�xvK\�_(�er�cO	�y2F�wq��S�
�]��JAf���yB/U����kR	F=�I��y���~p��TGZd�)��	���y������kJ7<jQ#vF��y���S����͖(-,%�U�H��y��z���
�EF?�n)SF�֛�y�k����d@��sf Y�� �y�D�8/�(#��-s=L rVEE�y�Δ�gD�#��^�98�����yB���R)H��E݌!�<��0�]��y⬗�>�
\t�U�=�5�g(ą�ybD	X��ą�r��u���y2l��~�4�`��1?�x�N@��y�A�" �d�I����k�R(��y @���XAc.a9X�*�E��yLܦzr�7$ʢ0�^������y�����"����ӱ-n��a�c��y�+�h;b� _N���A%�5�y��8?dְ"�N6M3�E[1���y��\�Xu��GƋD4���@ N�y
� �qR�R�I^3RI[�$!�"On٫��� ����GMl"̃�"OBi��l�)x7z�"@��DnrLr�"O��V�B�`���	7J8I��"O�	�Rc2<��N"x>Rl�e"O�:1!`|+A&��,��`"Or���f}>,�z'%�O����"OH��c������y� �Y�2�!�"O�q�BNS"E�z�s'�5��"O�m{#΍c�hM�F��ͪ�"Oظ!�GI+����acrڤ��"O��h�$V�3p�A)'(�a��\Ȃ"O���$E'Nt��	Rg�}Vp��Q"O��g"%r�V}KU��fO$��"O�Ųrl(l�x�X�'9�a��"O�QaCQ4y��&BɄn���G"Ot���O_�(��!�M�K\�� �"O�Ʌ�!T*.��D�Z4��R3"O��qB��S� Cx���T"O(��,���:�Q�B�6NT�Rr"O��t����b@ ���l����"OV����
-��=atj�m�@�A"Oj<����x���'�yb9�"Ox�2�n�9�|���h:�K@!�y"�*��a���'(�@ȅK��yr�T�0 *��=  |D�dI�
�yR"��
�y�oƘ�1C�F���yB'�6s3�}�3�S�vކ���BǍ�y"�&T��@�B�j�~���Ï�yRGA�z/<� UA�$hB�+Q+P�yBgD�d�p8*��9\���+�G��y�.) ��SBdS!(�J� �e��y�'V�b�)+\y���С�zjC��2oBnq@�E]�W[��xEd�%�tB�.�����|���N )�:B�	�b9H��'��E��	!�o��qP�C�	�u���BL�E���ҩ�xz�C�I1"_F1!s���,ٻu��8v"O�$���%(��}����5so���"OL���BߊF��@͙�^<��"O�3��F���mR��I_�h\�@"O��7)!q|�������guv!�E"OH��'�2\na�d��sp�}`�"O��#5�*f�Z%�6"j�X��"OL�w���A�f��b�*OZ	B"O����#m"�}qd'G�A�"O~hYD@ۃ*2hp�H#*4hh�D"O�\2&�B~�ሆ��	Z�
"O����C�[9����ۙI��0p�"O훐��]�P�*q#L���q�"O�逖B��S�4��B�%�v��"O�[E��O��BG��,�6=�Q"O�<`WA�!�Pg�f��C�)D�� d�?xܜ�"��&u��:�%)D��Pf��M���3s0��!��4D��y#�׋n�j��a��<5^�!(D��ՀB<W0�`�
IL����+D����+*vm����!f��58��$D�L�oJ>2m.��b<Wν�d�$D�PZ��F-s,�4H�H�J�Θ0r #D�p����h��ї�ۜq\z|�5d D�P�1aȠz�� �7CZ)�:���L?D�4@�gУ94����T:Y�PcW�;D�|8���0$ ���t�Q2@�����8D�� ��&�z�v݁4�2C�F,KE"O^��W�W�G��paH�1RDLK�"OH�;6m߲2�8@U���Pn��"O�ɈejX*41�w�Q�k=�h�"O�0�@�J��bWN=-�;c"O =:L��S%��y�n�2RAb`"O.��3��}���3eB#��q!"O��rQސk�|�v��8�L\�"Od]sbE)BY@�KC��t��"O<�	ƍ������
���8+�"O��2a�%|�y����@pr"O"�a�n�	�d�a%V8L��x�"O��%Z�|I��	�p���7"O��KG�Z�"�X�+5�D�@u�U"O���?$9��vM_� �j<�"OXxQ��\������-�ĵYS"O�8AC(ӆ4�(������E{T�"O�(���<Ffȑ1�˟Jp>�*"O�jRA��t(�!�Z�{k8Y�5"O�$�����!�*�;��rJ�a��"O�u
)J(ie"�w��!e�\��"O�@[�矋H�b���ϛ�<��H��"O��P����.À�Ά���U"OX���#�,T2�"��tʁ��"O����(\�ڜ�R���S<$53"O6�V��*`(��%K2���"O>�'��2�6Lapd�9.pYj�"O�I���#9Et��I�J��"O���ט	��y�b��2%�^�c"O�����γ$q������x�>�:p"O���L�>lQ0͒��J0PB"O���'��4�`�2�� ���"O��;s��2$���"�"'� ��"O���#%[jHs�"E�VuV�{5"O��WdP+@�� 9�B��ym�$"O<��`�؞Cި(��
�>Rd$ucg"O��K���57�5cA��LP����"O�M���',���$��>6ȑ�"O,��� ����	A��1Q"OPl�p鄺d_�9뒍�=\�>s�"Ox��C�$A��;I�!"��"O����G4|䍫q�U�W���!�D	j�\�K�87\	pA���!��U.1�(�U�X�9	�ArS��}�!�* \L!��D.��Q[;�!�$��r��s�J�褻�o��b�!�\80�d!�0�ă@�(��!ʔ@�!�J&_��p hY�@����Vm8!�d��r��d��
6��H��P2!�d�&(Z�������b�%E=!��P�nYb��c��ŧ�f1��'Y���&"1F�ѡ �M����'t�%��HL;ڐL(�@��d��'&�-*���|�u�&њ
�x���'��Y��o/15.�Q⛹xy�!��'���Cf � @�x�O��`���C�'Q��3fɚ�?s
dk�l��V��L�	�'�R���	'�B,j��8Y�(p��'�Hp��e_VT��F	JT�Ƀ	�'��0$jŒO�iZu,X*0�lI	�'�<�Tz������� ���	�'@���Q!�!d��PB$�0��'�rE�q�7�B�ӐKS����
�'Z(�3��C/X��9�n�Oh��	��� ����H:c'd�+��ۢ����e"O��*Q��r%F��$GEF?F��1"O�[��m>���GZ!�3�"O@�5C�<3X幠`@�X�A�@"O�Q-�4V�f�"0OG�j��u"O��AD%�0E�$���<`_�,(�"O�0�efU	]鲕S���zUd�3r"O:ݣ$��uC�i���A8W`�i5"OVm�A��y��]�SC�5E:B�x3"OĈq"��43�(��(6R�""O���|6��J��L0t|K�"O����x��YAʊ�rH�A�"O�$ P����IAR'�� H ��q"O�l����7��T�F%m!�B�2R�!�ݾU�݁@��.5�D���S�w!�D�4�P"$���h���_� =!��+h����S,Mg�z��!�Y�&���)��M�.: �q" g�!�ą�%�,��'��J���q��!�	GJ�C��۬qE�,s2`�E�!�$L�
�� ��*G���d���X�!���=b;�0LO)ܹ;!Nɒe!�ę�a��u�b��MZ��*��4<|!���y�ش��\�fE@���@]�d!�ǮjژѲ���&�J�X���!U<!��8�����؅E61(v�R�	'!�$�7ΉhG��Nj0���d�5x&!�L�C]>tQ` Lj��酤��P�!�?Q��=���Jl�p3dD%z!���$�(R�+��%{nS�C��9k!�0 /d�)��פ4���h��ۏ\�!�G&+���'ș�j�q�ē�~�!�ړ*�L� c�c֥8���5�!��U�Q��'4�|��	�I�!��>농�DoȩI�fY��ň��!򤖕nNzu��$��d�.�!�D��U����G�*�ni�FA���!�X�["�	C0+e���Hrͽ�!�d\�F�}qm�TyF<���Y�e�!��*Q�LIyd�%m��a�6	λG�!�3��1�-E�6q������|�!�-Ez�z����	4�d� n�h�!���+|�9è�L�ք��
^�,�!��"��PS_���y'�L	�!�$��mm��3���!
���hߧ#!�$����Y�HBs�H�h�[�!�d�`�$��E��2:ܐ�!��L@!��u�n)�uOB34�ɉ�
6!��,A���/VO�E�e�:4!�d��6$��Arm��F,�\82��!���2i����3%\���G(V�!��3 ���t��X�䨔��!��l�l�q���v�
A�0�T�Q�!��);�d���m <F�ډ٧��2�!�䛥�R�`/(a &�Z�!򤑭x�p|y�L��L��a �E�^�!�d�:n�Hh�G�-��ztDT�L�!�œ^����X#e�*8��R4)|!�䃯R|8T����(�$���H9!�dP'2����#�Tj-dкaH�0�!�dB�&1����O%�9z��Uw�!��3Uv�z � �(	v)Y��S3�!�dQ
&M�$���;3�L�P%D���!�Ν":�A�mةN���[Gcŷs�!�� t����3u�i�'H��j���"O���W)��I��p*wkJ��� e"O�XrU&��xqz�qp!����� "O@ �2��*t	�h��0K��qh�"O6���AԸp�B�@�o�,��xj�"O�x�(\�Hj"F$]��L���"OJD"��A"j���[���&"W�x��"OP�RiS�*��b�N9�d1�"Oε�E��dt6}1�F��81q"OZY�T�A��^Ia��/>����"O��'&�80�X���ň	���+�"O�䩐��S�8Ȧ�U�Z�"�1c"O��k��D�� ����2�>�KE"O���7I�/B��q	W"%FY"O�dK��!,��!m�;���%"O�X��N�E �B����P���H"O��{�Nw������KR	�L��ȓ8n���w�%1l� ���� ��ȓ^|�f�1o��0�E�*2S����`D���E�x�L0���|D���ȓ�ɳ�gC�l���;Q$��{eB��:�����M�{��%�b��3�B�	�%s$���kͦ���w�GR��C�I�n�~݃�#\�Q�rY��k�ylC�I-2��z3��b���%�?r<C䉮c�(EBt�A
uZJ���iC䉄M4��#�X�q%(��&��FC䉨im`c��L�>��ؚ��;&B�ɕjF�ͨs��2ǲ��ML3a�B�IR�b9j�NѲS'���+���B�I�1q�0�v(Ɲs��Ӊ^��nC�I����!u)�_�dx��h
��XC�I�n����Q략gj>ԲT��r
C�	�V��aåß#��9�Ը7UC䉬g�EKp�Y"͎U	�����ȓ{��I���*Vp@�ݧ�
ćȓho }q�R�ܥ�N^%��P�ȓI��A�)�N���zb��$j
���z��5Y	�Bgʧ�H�2�T�<1�����	@P0JՍX�<qщ��z�� �!�0k�^5��
�Y�<y�N�r�^�#�F�3�Z͉dY�<q��f�~����[)u�xhင�@�<�a�h�-���!+�%�	R}�<��g�V���Ƙ�;b6��y�<9e�-c�r�ځ�U� �BI�7��r�<�C0�4IWH��	v�hGn]x�<9�^�H�X�JE�9!�\�"FO�<������P��5~���%@N�<� �[�,�k ����E�p��c�<i���n*f�bu�g&�-��Fb�<Y�
�B����x z��Ex�<����/�a ��	U�T��p�<�'�[�s��(�I�P]���eRo�<aՏ�7*�`�CR9���J�g�<���M!T%+T��4Q'vm���a�<�?sf�蘷-�����	6��a�<	�N�Q�h�RG#�'@n:x�f�
`�<!�
٨/�!:B�cN�"l�\�<i���1`�A T-!&+<@�D��t�<��#ڿ9�t;�2n�A��Fq�<q��P*&�����ݻ�C�l�<���B�Ӓ4ZwJ�t >�[f	Rh�<qfٝd�29��n؛&m��QVK�i�<� �-��/,�*"偮SO ��"O�Ize��W�\0��
Q�3 ��"O���EHЫCY ��ki�D�K2"OXu���D��.���Y�_���``"O�0F�1U �q%)_(Q�¡Z�"OԬ0 MP�P����4<��ɘr"Ol9x��ݣc��XhsGP�����C"O�\��h�Y�l�WF�W�Z8�3"O�!��l�o$��$̩er�ɕ"O����"�\E��+z�ѣ�"OFذn]rzQ��dB��"O<�C���Jib�M���^9��"OEIVH�$f �5�6@�<B0"O���ĢD�]Rxx']�9�6u{4"O.���k��]�~,���W�ls�"O������Wϐt+`dJ�o� ��"O1*�m|��[�b�t��*�"O@�:����8pX�! F�5��"O���R$ .5j!/�1�#f"O�I!m��ʔCB�������"O�\˲�ݞ0�8��ǂ�\���rc"Oț���������w�n) "OD�*񬅘��p�dLV�2"O$����Ww� ��CO%m	��"OԜ��"�fMSVg��q��`��"O���DߍoF^]1��Q7;Ra0�"O2d��呧xk&8�Aȹk<��q"OPܡ��#�PH�T**����"O��d�>�6� '�Z	;�X�T"O���&ā��P� �N�����"O����N_�����×�:�>��t"O���Տ�r���'�q�p�;g"OT�+�ₚU�N��Ñ�d�2�"O��Bw�W�(ɨ{�d_	;(��ӧ"O��%�1m�)���
M	�"O���fK��6	z=jS@�
9J^T��"O��j��=c��<
��	}p��""O֕;��R��m����9Y��Jq"OB�[Gk1,Fp1t놌a����t"O<�WFA�^n��bkB���\�e"Of �H�p���q���)�J��"O@%�U�O.?=��hN'TΘ��"O1�ԡN�2�N<���?�l��"Ol�B�fװlL�����5cp�d"O )�e�Ԟ K�P1�L��\"OXX���ԣ�xis"��>���k�"O�%����4��٨��^�$�e(�"O���� �nJ� �����w���@�"O���7"�oS
Gi�4"O]IG"OzmR'	l��LZ�%��$<:��U"O��!�Z&t��*�f��1�(I""O�0@��89l�B��$xR����"Op�0�H�G,�zE�Ce�p"O��Q�BR�>���1C�v��EX�"O8��D")Y�,��"��Q~�qPp"Ov�z&C>h�̓%+JCl�ae"O����A�% ��qB l��	T@�"O��1T�c��%a�\�p��P�"O�jc���a%��Eǆ��` �"O6����i��� �|lR("Of�ȁ�%z�*|C�ɰ��9D"Oh�0��[��򷡏�;M��1U"OXe0�,�7���Z0��'�=��"O��A�
��N��1,�(Z�TaI�"O� �����'�H�ZS�EH�l2�"O6	 7'�	�`i���X7rs��0"O��8�`��
���"�IR}W�m8S"O^��'	*+�6m�6
Y�S��z�'�v��˻\z���4*�|q�'�Z}��j�1O/��#�&k��I�'�0�؆/�F��pC%C)��xX�'�d����:+�-�hϴ�2��'��E+S*L�j�|��^�)f�j	�':���&D��)f���3��ȓi�qi��Н9���IsN�$�f$�ȓ4d8Q��/K��y��'ҀR"��ȓmnp���z3��RG�_�b��7z�p�.�4d�Xڴ(=���ȓ[j���E4�����!� �^`�ȓ3���u�̚Tx�T��,;m]���ȓ{l��X7�_�|�ĢaA��v$��ȓc�r�:Wa��^�<C!i��JkX�����]2U��'��p��(�=U����/j��8�c��q��S&�q܅ȓH��@qON�� i��B�L'�مȓq�uH��L c�8��H.l���ȓQ\�(aAΎ�T�����_Ӣm��;*\ @'�1>ȵp@�#�6���)�J���ᫀ��63fL��&|E�C�Y �>��-߂2�d��f����@9fG�mC�҂}�RD�ȓ>w
�iҮN�K
n��c��V�Ju��;��\���з~{vyb���e��B�ɷn����6T�t� �� RdB�	=i�z��!�0c06�  �Wnd,B�	�3�h�Ҵ�[&l�<��� T�?��B�I-vj���΀XQZ-��,W�C��49Ղ��wO (8Dq���m�*C�	��ꀃW��"r6e�P�Æe�@C�ɺ>q	P0/�3���$��b� C�>\q��1@�L_��Cc�?�$B�ɯH��AP/dD�剎�E��C�I�9��-+P��9% �'d��C�	Gv��gȒ��� btd�2~D�C��6|�(����%	��D�P-� Y�C䉊
X��@��~>�\���,[">B�I�1�6D���.���kS��Y8B�	"sXZՊP&�9eP|`"�@LD�C�I>��a`�ùc��ѲaW��B�	�BU���DT !�`i�HƂ(7�B�	�\�����^68�r3n�!,-�B�	�tB�D�1��8~azR�ަ�~B�F��(@�`Ml
�كL$?~�C䉕R6���)Ԃy�Ԑ �.g#�C�	�A���H� �t )S%��[�C�ɺ%����K�q=���O��.C�ɤZ�<�ؐ6J��9 ��� [C�	/jjĒ4��@v�6(�5mC�ɮN �`X�㘪M���	s��u}�C�ɤH�HY�i�7m?�T(a�)H(�C��i��H��� d��d�mלkֆC�Ɇ)p�����ǜ6���a��	?a[B�		^��M(S+Đ'����s+�	��C�ɲl9���N�Hm~�+�`ƜE�C�ɺ]BΥJ舏?� Xd�% ��C�ɜy��,�!
��a����e؍M}�C��([M �h�Ą�i��%�Ճ��B�:�e9FG��E��P�A&m�nB�)� ��g ^3���POH��"O��A/�P�h4���qv�1�"O"L�.�)s[>�H���=BV��B"O&q���	'֞��N�����"O�0�Â�F}��r�mȗ)�,��"O���a�?xH���I�}��@��"O�+QKP=&�:�)2�ҩP���D"O�8 a��
\kr�
�v ��Җ"O��� �X�"�
� �v-�"O�m�f&��#<si<S܂\J�"OA�S��4zk(�����(��`#�"O���E�
~ތ%#���#�:�`"O�(��0��C����1�b"O�Tr�X1R��pI��\괌�Q"O8Hҗ��D��ixA�$s�p}B"O�x�K��2"��r��D*)ԮM�4"OX��C+��NlLj��Y4Y�� �"O�!#s��g݀|�у�+A��! "O@T�C�H wi�-�$t@�"O({���&9���3�')`\d�A"Ov�s��]03������ŝV����"OJq"A$ '*��]�'Ȏ�9@t�'"O ��k@'�fh�P�Q�@��Is"O`=�p$�u���yG+I�1:���"O�q+��%�5`H8c�L#�"O(�1�3-G�݊���$����f"O\A�0ƒ�-�D!Pfn٦"���R�"O��S�@�Z� �9o۟Ji<�"O��z���1eb!�M��Xz��@�"O$���#U�k��$�c*K�/\dy�""O�%0$6Q�)�uHG�D�0A�"O^���) �\�q酀l�}ҥ"O�,���>+��y�����d���)D"O� KӦ���!fD��"O]!�d�D���q�K�f�V���"ON�A�c�<l0�jԌ���z@ʶ"ONة���u�`�4�ӑf��ɣ"ON�
� Ԯ����Fߎ^n�X�"O��3Հ�p���uٸat�A"O�Y���u2��"G�\�,r�"O��A6�M"w��̣�G�	Or$�F"Ox<��i�N�~u�3M��d#�"O޵����UF̈a�Ř�hz�՘�"O$�:�QI���
W�Kvd��2�"O,eGDّ'䈑{ n�oʽS�"Oh�u	ɞ('�5�A�i&တ"Ox�dM�=~�i� �v�)A�"O�9z��ڬ<$��i�%�2i���b"O��hs�СL$|(i���`�֤�S"O����)?N���"��A�D��"O ���ګ5�q􂃁�\�q"O
�1f�$s@�$�R>1E��"O����-W���w)/J� �:A"O�����	$�Y+T�ˇt.�:�"O ]hC�����GH"!jp�`t"O�y�U*@�AԠ�!��ڨzKPD�s"O:@b��
6L:�h��O}Dx���"OTUI��P&#�P�t�P�eGz�ɰ"O�����k����A��5x�!"O �{�d"U�ed �>4$<�"O<,+c_v�pH2��j��L�d"O�X���9��
�Dڊ!h�TXr"O$	�s*���n���(]$��К7"O��bP*F1B-
����þm��`"O� ���H�y�Uɧh�>��h�"O��"�l�Xsd��Ǉ�k��Y�c"OX����	�
�����{����t"O���(��L!��'%5:��u�3"O���o��Q�8 � �BX�(<A"O�h������&��ec��ve���"O:`�2��<?���2eD=d���u"Of��v�OA���'䎺n\>���"O��q�	U�|���4�nͺ�"O̤K�3���@���n�b䫡"O.Y�!KҭjT"%�"A�'t�Da{�"O�l�B\&^�^��ro�C�$���"Op��R b�����O(}Xڍ��"O�-*E��xQ�*N>�R"Od��$(Ӎ$S<����U�'>�r2"O����rY`����t#�Ё"O&]��Z�o�\��@�P2s�`r"OtL�u@�A��@�)�'�J�b�"O2)��/�,`����v�>�b�"O�(�㘋�����<H@�1i�"O��CЌ�oz�-�k,����"O���3�s��9�O�Y����7"O�񨆋
$Xq�:4KHD�^EJ�"OT�y��>Sd)�5���L�"O(�h�N��{���CĽy�.��c"O��b�˛ �<��Pf��P�>��B"O �����K����a� r �`"OZ����"-��8Kw��#�V�� "O���]k@�RV!�\T���"O,tc&g�2G����F�O�O?�}ȶ"O2��@��B�NI��8�T���"OL}�"�غ�a �E��2�"O 	��,z\��@�D�*���"Of3Q	U��� �ћV"u@�"OX<9�!Twp!ڣ�Z%n�ڜ"""O�X;'�S�j�y��H#9����"O�r�f� H|#%`:J��r�"Ohm�g �<\C�	sD�-?ބ�F"O.L"���<��)���ގ��*�"O�PY��K��|�+�a�\Ě|��"Ob�EzҠ�����V����"O��*g�o0,�'ꜻ=g*	�$"O�y��e�=#��٫Ĩ�5Ie�(�"O��橝�9&r-x gߐv+�4;�"Ol�9���4E�Z\A�/ޜI�Δن"O^)�����*�����A3c�Lɻ�"O`P���;4P@*��ACyL���"O��L
�L��H�
Dc�Y7"OЄ��U�x(.�x�W)]H�1��"O��r��߬*0����[�$��8�"OTQQ����?�H�ҖM��'��L��"O*�������5+1�
�E�f�c"O,��+Y!9DhܸPD�*��PU����=a���ϫ��Y�� �'aNd���
!bS��
O���N<����S><�U"O�1
��8B7<9 �.V�XG�'��d�;uQ
�������ϊ=k��&�8D{���V:_e��y�i�9���$����0<�J>�*O,�ǧ�C4�)G�-t~��B"O1*P��g����F�+l����'t���}��	k5��D?p���a�2%t�00u��z��?�2����f��-��="��Yd|��<����ïT}
I��C2m�f�KFƟ� ���A�0?	�n΂*�` 9B
A-Ok���`��ݟЄ�Ic�� ��9���;#N,��W�S/�l���"Oz�P"@0���P"y�,A��I|>ȡKgQ����E+NH��m�>�yb��#��Ǯi�tmH�" �>�Zq�/D����ӌ�P1�����K�0اN.D��rH�#�����/x����6�<��.�ڔ�TaډJ@�:VS�a^uI�'A�O��?A%L���D�{��T���i�K�'�����}�FBWT��#%��^�x��m�O�=E��˘*.���k�
�l�:@�?o�OJ�=%>�
��A�%k��yQ�(4,[��&D�@H�䘬A@]'ؒ;%�a{� 1D������~z���B�s������$D�@����,˂��2�B4)�\�!#0D��� �Z.yg�4�2�@S��0�-D��A�5%̈��`~�|L�kk�����%Hzh�h�OD fm����ΘB�ɒnNy#�֤*�<�3��M5OnB�	%yfv0�dLծa�E�w�Y�C�	����X����UA�Ɲ�,p�B���@��KJ22�ڐ��NݖER��O�1ۓB?��[E���6��qs�A�T�$�ȓ8�d�p���� g�B���ȓy��ݪd�5vHXR@ӻRӚ�E~���?���K�_oҥ���j�آ�o$D�ta�ȏMP֝cjn���Ф-D����[:-����K�CH�IIl+�O~�(J��$��-ؒHk�5QT�%�(E{��D�"f�>}�c��G;0=kѫZ!�dS�&��
F�O����i�'{�!�d��N˨�V'�J��RJ��!�d�-%@U���δ
�z �ɜ!�D�<��Y�2�_� ����׍7��{"�J�9�|���"��uW�a���	�a}ҕ>�ĥ��38aӢb���b�W��%���ݓ�%�P�Ɗ?Tt��)D����G�<,򏄟�N��� $D���'�ȸW"��{R��Cb!�ǩ.D�(J���7�]��߄{	%��J)D��pr�ܯ���a A�� )�4�I>:Q���mr㖆r��x!�B�.Y�p��"O~�*��L�>�<�PU/��fT�d�1ʓ��<y�߯=���A��:K��D(�]�<I�@��D!��z�Ց@q���w�W�s�C�	�_ 4�B��6]��%�<�*��D#�IZ��@��[g.��c��,+�C䉸E f��A��z'Rы��H
rc���:��v\�@�($!K�&���,B�	(ST��)�dG2��`�#<���j��h����wjM����t�w�@�"O����cʬ,bSN�q͸�:�"O���(T,~Eh� 6NW	 ਁ� "O�-
�ꞦW=���  �t1��"Oz�T(��aZZ�16nږ�T�Ke"O����Y6Z�����C�f��!"O��;$T"jt��d�X91��`��xR�'/�z�#A�Qn��WA�1~�"E/܌�y"�]4j�q��h����*������'��{��"B����E,t$kv����O�"~Zsȋ��=�e�[�hJ=�C"�M?��Zf���R�(D,q�æh�@�$�D��	7IL���X�GDUQ�̱z�>���(?Y�iҬa ���kĹ!M��(�+O�<����`�
�	4H5_�H���˅c�<� $$���	-���p�� ])BH��"Odk����������� @�!�'T��0��N�b��9�%���V�@Si�$�=E�ܴ��Z'�ԽA��=r�ȥL-nP'�F{��D�=�t9�D˪;�Ha�T�I+�y2�M#@��g�ߴ.춙��Յ��'�����Ʉ5S�ȫ����	_��;B�P#a��B�IE�TM1+ �7��k�>P"<�	ϓ7��m�eg�gA]�v�94b���	���C�\�Â�L�ZtH|��! ���O�%�
[(e����9p��a �'w���1o��D!��	G*����%�O��I]���堄!V�P��E���	|yr�O���$��;E��-�!݀HA���t�&D�0�6�/˔�jl��m�Z�h�Hd�ܔ'!ɧ��Ĥ2O�}���0�@�g�A�~�!��#Df:�+3�M��ؙ v�T�d�d�=E��'e�
B9m�@�Z�M��h��	�'�и C��t1��-�n\b	�';dぃ��~��@�q��)��`*	�'��,A'ӎRm�`�����¼�'5\��l�:E`<[ᇞ�����'�l��CU�7�2@��97V@���'�m� ��^	�)5��|@�R
�'䖼�t�&s ��JcD@�wkTH�
�'�zEk#�R,|Pp���'l��}I��?Q.O꼑�fO�7x��҆ܥW����.LO�Uo*l>���Ń|O��"O�J��,�Z��&�
|j�$i�"O��zr��l��Y`.		���%P��F{J~b�O�(9���0�Ρ�G×r�Ȑ"OX��X*U�z����Ğ���( ��x9p�)��?�\�B�`���P�H#+����扲~~a{����؄�ן\�4�k�$z�bm2�0�?L�������䗦K�- Dl�0a9D��j��*<�B��=|�������=W��@&�l�u$,D�x�������%�G�A��p ��+D�l��&Q�=x��ԅG�>d� �f�*D��3�V3xj��l���S�'<OB"<�C�[�|tUڕ��R.J�`uJ�K8�@$���"@�(&-	���Q!v��q"$,O��'���O���b��R�*�iGfw�,��� ?��ٌwͼ����ҼS�Th�S���x���P��}a�jMGܬ���P.�yb�_+�X��L�BYH�pf]7�y���X�z����F8@(� �P��p=)�}b��r**�|��48	Ӵ��xF�2|�#wȓ|�Α�3��(J!�$�6Jg~��/V;&s�Y�C &5!�P�[��q`����4oz�?y!�d�{`d�F��^�@ �FJ%��y"�	">���Y#�Kb��diP�	.\�C��4
l��a���#Z�Hʄ�ɚV��	�HO�>�i�&���@��gI�|Q��:D�XGj
vTx� ��(2Lx`5�3D��(��`��Ȧ
M�;�
I g6D��p� N�I�RFI6��t�5D���cu��x#�j�aT�����2D������"����������=D���E�ʐ�k��B�$�r@&;D��`�ɮ\ǲ�I,���89��8D�� S�6�A2��	�'�(�G%9D�D���(x�!S$FҜI�h#�L5D�DddF�6ܙ0S@M�c�,I0�=D�� ƕ"�%ޫ^c4ĒA��3s��� "OR���l��M�<j�mҲFtJe��"O:��W�ҩxa)aF��9en��"O�4��H��<�nI�dQ� �"O]:����o^RV�LO�f��"O�m��μ<�U7I�7D��z"O0`K��Q)O���r��[���"Oy��n�h�p驱Aߴy��I��"O"��sF�/Qox��j�ښ\ڢ"O���BJ1���wi>[�A{�"O�37+N<(��i�aF��r�T�2"O��Ã��A������F�FYc�"OT��U�H�N@ZIJ��BT�<��"Ovl�0���;e���#�Jk���"OV��.ȏ ڎ��\l�"O�(�,�$q8u����w? U��"O��ڐeQ�i�4�;ao�~Z���"O��×��8Ax�P�ㆁ\#@��R"O�ԓ�O�?a������
��aw"O��2T�)Z6�`����c���@�"O�<�`i��<o�)
2`°X�|Yb"OҤz�
l�DP��E�U��T��"O�i(�+��D(��ՀI�@�"O��塝%R���f`��C����p"O@|ۢ O/xؽ����&�H�����"!�V���4*���ga�Y�1OX�ДAͣBw@r4�Ž?��z%"O��+�P�_�Y�(ܦmr���"O����.ĭy��<��
�8q"��"O��i� �?F��K7;u(u�"O��a�Iͩ:�e3$�\�M~l�Ѱ"O��r��`r�J6���v"O2����.Z&P!���"r����"O�{�Fǚb�p}X�Ǉ�7ÀP3W"O�m�17C��"���o�:u��"O�;�:{"�,J�k��	[@"O�	0�@�(}L��J2XZ��C"O��� &<�09�ݖQ2�I�"OB�����;�L��ͬ1"��j"O�5��/W�Diu��N��[�"OTlH(1�F=9��u���"O�<���D����1�b�'2D@�"O�h��=Y�e
Sj�X�4|�'"O��Y�J�E�`iA�a���s�"O(L���}�!0u)	0(��}�1*Oh��`������P�J12�',j��D�ýO^��YQO��Ntt�'���01O��zERq6F�Ɛ��4'���t�Ȋ#���(O?7��{xY�GC����(1��N�!�$���`���O-�&���ܦ'��DK]���:���_>�ea"(��l�A���z��QڱC�4���I�9��� ���n�Qs�Ȝ	gLv(Q�iL""�*��k��f�ȑ`��'N��J��4B_��� 3?���}Ҍ��bE�)�ǋїz�:r��9М~ZEi�I�H�����Wi��E+Gl�<�F�� dBf����2�rd�\<R}�P�#��|���فe=�hJ�I5ʧ�V�ɞm�n��5VL�0uf���*C�I# J,��1�8��G-a�!
�����!oS�Ҏ�9Vh#!L<F{��(B�1�DG�p��L���<9��E�h����&PG4�ҡ/D',�C'L`C��!���@��j4B�;v���d��9���'�L!0t�1@�Aa�' 4x�q���Bfh��Ë=~r|M�t�C @D�OT�*��N8����L����K�'`�P�)D\G:���II./ �г�a�PЈ儂�:�����>d�$?���b���y�)S��|P���:�}�h/��x�.�'���A� J��	�
���z(xr���,�d��e�4|�aN%��9�	22�i6O�=<��{��A�5�2��D>z|�Mه�܁'a�I8��D�? ���'��>h��eE@�9�� �/v\��Æ��p>��X�8�(R���&7| �wE�y~B���If�p���v���Cë�Ot��$���`��'���;���L}�]ŋ�np�ȓ�\���7N��4OO�'�x�C0�O'I�E�����J��ha҉����O��ᑲd���y'X�x��x�^iҕL���x2؇��A�u��f8�r7b]�F���Zd��16C#p-
��+U��Y�ƛZ�'�Z��E$�CZH�����
%(lXb	�#)"��Դ\�D �c�^�J�z��UD��ă�c�2{2L�pGAr�Nex��=?r���	�&HcD�$����ւ����I�0KF��uM�y2��Q�['Dz�XU�\�P ɗӟF����(9,�)ɱ���k�7#!�4;|�	���%I-N��S�сm��a�c石)�Rh��*9��֏�4��S)PxL-���)?C֢�B�� �H:��!��#IG�L�Ӷ��'Ȯ�@5�(3>�yQ��D�hP��#BlKR�D�RC�_�@��&�I !�6��2*�	�j�yWI�*���D�Q�\x6��fA�1NQg����t� :����̋
O�5#a曜J���jQ��p>�aꅙ7,Mˤ��6��l�D$�m~�IS�l���piH_0X�`SFB�o� �� Z������D���!�$�Ⱥ J�V���� L:$K�b[�T�q���U.K3p�3�DC� "��E���=�L�T�=!N8�Oq��E	��y���t�(�aA�2]��5E�5�x��i���a��gC4�9v�u��� �
���DuAF�Ӟg��y���a���!W�'iv���@8oW��0I8Ws�9��M�V%��w��CEGQ@nx���JZG3��GH� �쭃T��=1��}(��\z�����љA(dԡT�D� ���$H�@���ɟ1$)��)
S�E9������A� �OId)�[�4u��� c����y���J\@ PO�#�T��U\n�H��������Ų)��(�^�ѝ'�:��d��>C�n� ����n�a�'�f�P`S��(�g�)�46��U `�"�'��[b���.5�%�M+��		�Q���~"(��I�,�|\2����!�]�Sf8g,��F��v�$�׈;fАk��'��!
���/�DA9�aY$��Dx�����5[$*W�I]Ɓ�b���.C	J�����#<�R�Q����y�?SQr�H�/M�+@�Z��M�w
ʮ��Y�@E����s�$MB𢂳bà<A��!Us���"O���"ȋ.J��,[��Z�pj��{Ĥ�/��亄m̳7ޠ��F�FMaxR*�z�Xт�b z��V?��=	Q��A����0M��^D�0�$!EEJAZ�O��Pxb�
,U���J��N�v�dQ��7�O@p�f�^Y�,�Y�&5�S��m�`�������%FE�C�	 .��r�G.�E�]A�)rj�W�AF�|�'
dب�
O.D,��%ʏ�$�� �'���2'��3{�*����T��H����pu�-���R��R�霏)iXQ�Dʠ��U��I�Tܘ`IT�Ćc��8�D�&H*x[��όWc!�Ė�]��aR�蓢
S:h��a@�5P�'�\���ooɧ�O���"c�)CtĉQ���S��}�
�'a(Y�`Ԙ>�Ĺ1fM�%d@�5��O�h��Q�g�I���	9$�ɷ�@`��ǆ�zB�=u4���w��[�i��"J�
�b��X�z Y��I~f|��� �1���uk�3u����f��Ë6}����� *��{�:"$���yR��"t�(�Zr灂�.5{��͟�ē��q2Hؚ��S��H�p�I�X�j���k����pE���VdJx��bˇ�Ь�S'�1���׸��~&���킗gwR ��ɔGg:��?4�T�w�O%i�U�G*U+�&Xч�S��HZ�F:�O<ኧ!D~qk1DГI�<��'�\-�ēeӄ�A/��j�LhE+�`�p������,�)+�p��,ج�e��R�4�SN�!o[�)�C�
(TL���g���Ի�LҶ�Ȥ����ȓ���B�'ڐAh1*�.�!j�
h��LȜҦ�Y�B�`�qji�����R���Q�A�0m4T{d�_���ȓo�|a �J,>��ZU)�<H��S�? �(k��
�NK�qi��_0cp�W"O����D#NM+`��_}� �"O���úL@���3gs4mx��>�!G;g����?����6�AZg>Z,�$�`9D�H��@�2���{�GȒ����5" ]�% u���@�g̓c���9��]�"���a/0ͬه�ɽb���yb-/]v����R�3I콁��=$���ْ%y��𑒬В����n�zj!H��<��COV��F/9R�%��P>���Y�	H��Pc�6- ���)D��s0�Ǜ#Q(Y��.9h6��g�<�4�N�@�����.͟��?���Ʉ�@R��n>&B�h[�B.D�x�#a�8i��ݳt@�����$쎔;\��'86����%g{�ϸ'�^,�e��?B��u� fТ+���	��a�P�U�ôZ����S��0Z������6i"|��**:w�}�HH�K�ޥ��"X!����Q�U���O*�J�^�f� pr�#�y�t�	O�ܱ���(ؐO��yr�F�As����(m�Uh�X��S#
4�9���\d`�G��NB�Q�X�sP�V4^h���E���y�M�#Fߜ	2 H��U+�@�&'ܻݨ(r�]��s��v�jb>c��� �L�l�8���+ѽ`ƈ��n%���@�M>�Ƞ"������1D'��//l\�Q��'�yq`T�2�@��o11f.̸��؍�w�W�}Ɋ�'�UI��b���Z�%G*��J�'�Jɚ��C7\��T��\� �v̓J�0�P�O8pE^�$��?��ǊF{b@��.�4�ԩ �)D��٠�ı-Ԕ����$7�V)�-�]ܓI��6��x�ĉ��8Bb�-U�jd��EԎ�yߺZ�0�f�@����C�R4�yR��=~� �S�32��T )�8�yۚ0������/�6��'�8�y2O�r�h+0 ��T�X	�'$�9�y"b��\�P��T��A; ���3�y���)~\��P!Hӿ=�	��"���yR��
]:�@��|�iC��7�y��O�&$.���&�p��"��@�y���,i�xi4�YE�PR o��yB�M�YZ�բ�Ą/%az�Dʁ��yLkL`x��T0Q��D莮�y��f��1�`��: H˳Ğ��y�ӯ�&K��7#�%���y�n��x���y6�2�CZ�y�	υA\~%��arC��J(���y2#9[Ĝ�S���Q5~��u�U%�y�!?�$��diȮK,0��)˂�y�1$<�����$ ��?�y�`�������΋\C�5����y��<�ɡfY��|ܳ�i���y��ڇ-�B��eŁg}~=��դ�y���`�5�ɔ_�0�[��ʬ�y�]�5\��p�ӏHR� ����y��
��%Ag�U�_�99���yB�O�}��X@�~TL5�y�COWN�	�ׇxk�@�m�y2��(Ⱦx�BˈG�}�"�%�y�j�<�$EC��?��� ]��y�_�f~1��ϸ7LrQ"�yrH��'�T�Q�.�,<��@�.�yreϋK�@�Qk
"p�d!㬀��y�G�X��� ��Jjdyf����y�oŬ{�͡�n��Yp�*%��$�y�A�dAq(X$d�8XT��$�y�o�	n�T�䈜8�0d�S/�=�ybdͼ> ��Xva5{tlH�'��y��D�^"x��셛j��p��A��y
� R���-a�ݫ�L�  <9�"O>e)��}%h�J]�
��k�"O�����.pT�
�*�;�z쪵"O��꒳�ŗ+	�Y����7h���ȓ%��zLs�R*ɖ2�Jd�ȓJ]0Mӡ��w�p��d^�d,F�ȓVILԒ�Ν?%���w�%^P=��;Bj�@�f6BŃ%)��r�|4��N��M���,�X9��!��/���ȓ#q�8a�OG9?�ְ��⍹C \h��i2�)��]���X'�Sw�0x�ȓ����'��}�&a�&�]�Q� y��$�}:�)J5vg��9Fd�/�����5�E1$j�Ly8��LA>$����ȓ8�9��@��FP�(�-�O�F1�ȓ
�� ��^�>��l͜��؆ȓ#"ܣr
A�m�x�	��M`�A��v�����F^�E@�xi(�DJ!�� ��$���F������ǌM�*��lb��!�$�3$��(Hۈ3w<�ȓI�����H�\*ȫF���xY�4��^m�ecM���e�e����G�� C���8~N���6�a�����sJXq�Bv��a"N��W��q�ȓW(, ��I�51Vi����4/��,��=K�
� ���J�
e�c`Yh�<��eҁgr,��	yV\E�Ī�a�<I��#��q!.��p����c��^�<���t�(��G���v����i�Z�<at��L�	��l�g���kb��P�<��5
�up��K�n�,Xc�`�<)E�_�h��T:��B9U��
vK�G�<Y�) �>]��b�/K����e�<Q7L��]+n%5�*�Thr�So�<��X� �H�Z��h�yu��Q�<�Uʘ�u0���ܡ,w�X!dW�<I�'�=Y������{��̘4
L�<�d�8C �!�d�`�m]H�<�uꟈO|� ����4��e�D�<���ěE��ă�D�P�$H��#�D�<1�	�=�,p�BL9>O,�A� n�<�����xLt��r퐾6�0����Bn�<9�g߅!����Oâ0x�����j�<9�ūEf��sfے66�yxU�Cn�<1D�Žg%1�2.�o
 ��ˉV�<Q��C�y1��N�3�بwGCL�<I4��D��}�B�P�2�&I�<�W�T?c�lE�@�7F��x���K�<�3�̃et��kpk_�
;Щ�P�R]�<�hh�9���f���Ӡa<�!�ؽwh����#J�)�  `��N�_!���((��[��o��Hq�V�6[!�D�/D���'�,�\P���[�A!���VfM
U�	cc���� G\!���L�ڌ���{@Xä�ʺG_!��[-([�)Y�>�AR-�(i!��3��!^�,�eH��\�!��T�/��]2%�ΑVT���I�r-!��-)Y��P�-�o���e�7)�!򤈸9\�l�7/��L��D�5��- �!򤔡Y$�7�ѕ
��<�����DM!��P�{�̣��O��){��L)/#!�q�(I���2L��ѐ�+C��!�	�W=RH��N���U��уo�!�� D�Q6�'glrȠ�nA
``2��"O�Q��x�r<�!�	�K�Y�G"O��+҈ڷ'~��1T��:ms��
�"O^|���?#K������o�}��"O|��Q,"����"��(�a�0"Of�a1�I,"���PgS�x;"O�ŉ�a�7u}��S��׻]�T,�6"O�m"`̆nVbXbpM�:�6`��"Or]�&L�5��l�BF�F��CW"O�Y�H� Z���f�F49���c�"Ou�n7}n�уގ9����1"OX��O��_�L�"3b�=q�(���"O^��dQ+.PB��2$K��P�"Ol�͇�_$��d����4	�"O�afJ��<��J�-�Z�k�"O6I��_3OJ��ХK �p����"O��OF�L��a!�����a"O(5���]X����?N�,�+�"O�]�7�Ȇ8.�B�/�;]��I�V"OJ(��oX�Ti@5���K
	�Q�"O���Q�J�n���[9 ��)��"Oj�)Qh7e���[0��\�\I{�"O0D�#o�9>*�:�K]�9z2��"O��3D��Edp��7jA2t�,;D"Om�&�[��PrD#ɫrQ�y�A"Ov�����0C��
N�H3"O:�:�.[��H��=]%�YY�"O�i�	O�4��YƩL0Lܣ�"O`��(ʈ u��zՉ�:`H�g"OЌQ��.b�|��,0x,j�"O~I�Cᇽͨ��莕(8�i�"O���V�H<��bQ��,O��Xz�"O��y�.�����=f��P�"O�`F�Ա���U���U�B"O���iل]G\m��&�uK `cq"O��C��0(���dC�F2*���"O�� �.GG#viQc��kޖi�f"O��u��7)J$�V��K�|�P "O�q;����/Տ7�©B�"OhU��҈ l�1��Y@�^���"O���ل�q���9�L�	w"O����	+K&�}X��Ж�@9�"O$= �
,C#�ɪ�P���	��!RC�`w0�|�'0���×�{�ԑ�f�I�9�Le �'U�e���
=H�PU.�yٴa4�7+��T���!<.-PaM�26LB�˶�˷ :���	4gk���7��W��
�Ƞ�z�ڡHD����LF�i!�䄺Kt2�-W�8lC0�E,0W�' ~�6�	[dɧ�Or��{-U��^��p��"+�dA�	�'i��N�9<|�G&@��bJ1�P�I�|5��L<)"E�$@:�w�Ό\< �rLIH<����v�ܹa�$_-m#��{3�=G���8�+��p?i&HԿ��u��HR�0�s�J\X���d��>m�O\�Ys���}�"�ej��)Bd�W"O�{���~h^����f Z���x㑤
�^��g�|�����WV�]BfI��	��[c�6�y��$3�,��4�T=?�<|Y1�
���L&�tqA	�����K.�E�4斑t�|��QZ��Ɠ)���w�P� �2�qC�"0!ڍ�gL�x0��	0��Ec �6@���`	�e����͐rs8OV�£���Xl��5�˒|E򨰀"O�h� W1zmJ�:8�E	�"Oʜ(��BCK��p.�aw"O�r��ʪ]D0K�jB/$08�w"O� �����D�LqP��i��amd�"O������B؂<iW�Cu@�8�1"O����P΄xb�I�5�qɔ"O �q1b�~��B�&y+���!"O��8�.��q�3*��"O���Sǝ&�N�����%��mh�"O& {��ٮ4��#b?�ja�'�>Ag���:}.��?���%���"��$�K�\a:�9PK2D����n�-;?\\�S������G�RM��'���e�g�:7�IPa�����X�lM,����I;2�U�PMPb۞xҌڳG4�܈������@��x���R)b������C��q7�*�J��u��bW�WQ 5�VT>My�ǏYN:�ZU@gV(�R)D���4��%xm��8�T�Ӫ�<�孀 Ht�0�oͪhw�?mCqJ`��(���&,��Ѵ;D�ԉ�!I�?�xy"Fίf����5dZ�-���'pt)�EmD�'��ϸ'I�(@�O�6��4�X�|�4X��oL�  �,��W��Ҧ�N��%[�f��-ú�%a�)o�}2�T\dd��P	^8#,�1�Ɉ���Ot��U#B&~Q���Tg�f����h|ш� �3�~�����y�,3-��	�C(N	�3C������, d��u`%G����$5�� 4��0%i��y���҂��C
�(��2j�\�҄�1]��RGɫ{Pfc>c��&D��)�\)H+i�t`�5��FDP�%wJ��R(^��x�zuaET�6�
ҧ��/����D[�y<Xdz��@+�D9wcMt�ax�b�^T݀�d�y��ch*�pˍ ,���d� 4�!�J^�������d�n,*Q�M��1���p"����S�'7+�]��)�5Ly 	���>�L��GQ�e��dֆR��u�釜u*z�{�N�
�c?O����)�.}W����A/k�,h!"OnayD���:aaД��+����"O��@�͞<���⍒�<�p�"O$�2�)o*��1�FE�X��"OR��.�<��,�r@�Q����"OHc�� 'A$�	�*�pؼ ��"On�)5�Z_����7N�.%��"OZ �0*äDⓦK�ZJTU"O`5�p^�yƢ�H&&��i
���V"O�mP���,q��S��{��HR�"O�8��.��*��x��M�U�Ա�"O@0� '�d�j���6F�NX�w"OD����_����e]�XԈ"*OP0ʖ-S�l8,�p�׵k�=��'e���D*��[EpE�ѥ�:P�d���'���J1��Xz5c��:���'�T��DP/W���@��~ ���'���ɥ@�6[X ���S�q��:�'�(	�F��9$ �b�A7`��x�'[$�H��_����׮βb"��
�'Q�m�e���|b�&@ٙ+4TT�
�'� �j"��
0`:�ʖ�X-3$Qs�'�V�c��6F�z0�˄)��r�'@f�V��YC�]��&=&�K
�'�=�')XD�fQ���[:�֥		�'�J�Ǡ�5'���de� S>�؉�'�f����wՐ-�%�Ķ�F��'��� �g�9�x��#O
y����''*��&��_�hY�� q�d���'\�9���5Dpy�Gx-�
�'c^�5��X���	�F�<8��'ܴY�F�P4��r��+<�$D��'n�8Á��Ca��`Q�%�⑲
�' RLB��V+<�����L�	�lB
��� �1*�� S�h��%`Q�YX�1��"O&����`c�����m�m��?D�`ZfDO�#�L�f���UL/D��k�@�O��:��o���W�)D��Z6��>�H�	TB]* �`��bH!D����֟m���4W�$���8D� �V�ڭtY^u�Wb�3_,P@*D���-̊�̰�Î�xz�5(b�<D�t[N�:Ү@)q��7����i9D��2EE��/����C��3V~TH��6D��*�i�%f�� �V'��K�<<j��1D�D�}x��qmZ�n���xV�5D�\���D�,�T��WĎ��ԫP"3D��dƏ*-�����,sf��GK0D�쓱"�4Sب���\T����2D��¦_*G��D�Ɲ�3��\o?D�(���ք`�.�[@��-i�6(���<D��) dQ*�~!s�K�{�u�#J=D�� ���cs^�;��D�t����Gk?D��`+�An�����b�t��%9D���VEך?=� 
`���8�p�0%�4D��H�)6a��m�E�Ћ`
��8C�)D�X(�F�3+	 ���b�rS�$D��zdcگ"�ʁ�,�AF�Z��%D��zjW�i��7#�:@������!D���,Z��� �`/�5 ��I!N>D�L2���.�L�У���}�����E!D�T��D݉ͦ�aMM�(Atɂ�d<D� c���ED4b@��? �1�*O��
�k^�R/$���X<u(�+�"O�D�@�"9e̸���5�Q��yR �84��Tb�h»v,
���)ҝ�yҩe؜3�o�n�D�j&C���'�X�ƃ��=�fY!�@L:d�(Q�ƙ|BN"A(d�i&�Zg����V���s��(�^=�PlT5|��P��1��s��'�ў�~ڐ�@�rUi��+WT��D�\�'ra����'����!_�2F�Yc�K���'�ў�O��0���R�sg��U-�8�V��O>����)�e�2IJġ��n�+��3��I��Y~Zw!��Eb��,ۈ-I@u#K�G�b����֏ʰ�Ђd��8R+�o?E��&�Ӳ���?�9R�*ۿFo`�ɬH���l���O�����e��fu�ĹrȂz�4�p��=D�Q���d��!Ȓ~6��r k��V|nؔ�x� �H���O
6(���̔lxxE�J�9�^�8�O��h����^�����`�n��ՆSeZ�ܨ&!lӠ5�*O8(�*O�?M��D�ڨ�� S���(i��Dy�&By�+Z���'2��I�nQzv�8�G�5��''��EyJ|�R�$�������{H2Ī k�J�I�N�Q�b?�3p�9�J=���&
�2�Jc��>QF��M������F*)�V!���A5�)P�N�H9`��rIUR?��O���~������c)ܺo̬H[��6{�<,��K��yk�'�����L"#�ϕ.UF���*��h�^0����p���S�l��aі��$ypׄP�i�O&�=�}��- [`t�A`$v
���	Zy��)ʧ�@�P�	Z�ȑ)�dMU��p��L������F�ۥ8�^y`a�փc2�-��	Z>��v���� �G�%���J'�&�	㦡Gx�'t�j��f��d��H�ߑ��@����!j��C䉐�<��늼9��ę� ��MB�C�I�n���׫�X;~<��יO�C�1�Բ��cX��Q�S�\�dC�	�8U��0P!ōu����͘w,�B�I�6�Nq���P.k��b��FB�I#Z���7i[�v����g�-64B�)� L�,�w��{&	O���"OB�y6#	�Љk��4]�����"O��4��
d"x�I�EX��p�"ON ��@Ҥ�T4i��J`����"O.�� -�$)\�6 ­Kz�A"O*�i��S�B��d��+ɸ�ɒ"O���3*�&��H#�-G	��Zt"O��+j@+J��P7� �!"O�hAS�W޳B��	�{�<����}}<�����8�F�"Q��t�<�%���/GV�C��R3",�$3�KE�<)c��
OL�:�Ɉ�,�:8ɑ.LA�<iA�������vI(�B��q�<�E͈<DN��G�K���xv�f�<�U`�>X�.a���M�H�H�Ma�<I��K�/�`�X�+<>����D�\�<y$� raQ5\#`�u�U&@�<��O�\�6ia��J�d�n�;7��g�<1�0R�~��s�o�$�����`�<)�ȗ��M�cJ�?DiK��R�<Ap��ebt)`@mL�Eմ0s2-�O�<SdG�l�H@�8.ꡉ��F�<I` 5�.�Y҃V�>vb�4�[L�<q��˰�����`��n<�U���C�<IujK��ȴ�Fč�~�,��H�<I�-X/;�40�Ā�1"���FD�<I�^�i�
y�w&��aT��
�$E}�<�u�QS.l�0*˧5@�*��s�<��_�<����&B�|�a�jI[�<1��2f��Y9�H��U�ȉ	�f�K�<q��[�/| �3�� CJ��r�H�<Y��%H������"t� Mʇ��G�<��`��k<�I�6�a���2��Z�<I�7E�Q;��wf(ç�q�<)2�_<k�2%�F�
k<lô*Dl�<1T��65���IE)Q�)���g�<��IIW����(��� Tf�<1��'#���2�惇Q%���h�<)�ÔHG|ܳt��j��$*�f�<���MS!͛�<VQd]'��W<���!+���TCΗu��S҃ޅ�L��=�<]��cň	�^��&@�0ưE��mb(�r��kyVq��F�M��P��+`0K�)F�?j����!��iȢ��ȓW���YQ�Ӣ:��<k�Lt����lN|}Q���=kj�"�'�'Sf͇��`�3�a�/%�d�:@��#�܅�g��s-���¥��/Ey5�0�ȓ(3���@�uL"D�f�>;U���y/P��ukW�h�n��4c�uH�݄ȓW���w�]��:��r�͛�VX��f!�P���V�%�P��� 0���ȓyoP9�Q��\nn܉BF�0)�5��9�iꁫ��^ܤ�4/�2[Τ��ȓH�1��BJ�aY�@[�☇�H�Ԭ�v��!s����F�E�|͇ȓQ"ȓ�K�p.���B��-x�\�ȓ�6n�&��K�U^���Vk�<)�g���t����k���"���l�<!��](>/xT��HP >��dL�j�<i�Ɏ~����;@} ��3�i�<Y) �D��y`��9H��E
�y�<ak��]6�@��V�l�Z�I�D�w�<ٶM�.*~X�8�,ώ8ʲ�Q�Lq�<� ���B�&~z4p�G�
�dUv"OJ�2q�W�!�B���\D�x@"O&�zrM�&�.R��Y�r+h�Q"OR�AP��\�8Qʠl-T��"O�9�6�
`�ْܑ� :8sF��"O�ī�B]�/�<(�8\Z���&"O��BW��l���`�5#@�i��"O��&%M>~��(a�Ê4008I"O� y!��D�b���N�J��pp"O��@��<���s�G���43�"Ol�䎁j�.勅C�v�z���"O&��lE7-��@�L�E�T8!�"O�Xb�mW!^�y����]��(�"Op�BaL��Ia�@�lU#-D�S�"O yQ�FG�j{��ҥaC�2��"O�y: �B�6�ThQ�o-#"�:""OX]'&�t�b-�7nI�1�"$"O�-��zBT�����"��x#�"O�a���)v���%�̿'�h���"O��G9l�CS����@���"O�q�E	-��P9���720 "O ��X�Za@ "B�$&XБf"O*��F���-������'P���"O���X�6�"���0����"OZm�������a/�!Ƃĳ0"O��0��<GwT܂�n��^��0�"O�Q)�"߄�V:޶�;!D	�!�s�\�2��R�����(�14u!���%Q���Zp���vKJ0y���0�Py��W�&^fM��h7O/�i9���y鞓T�"�0a�S�ޅ�7LW.�y2��Ӕ�I@�0;d�:�i��y�&E"nY|	����0ϰ�Y5/�)�yR�A�Aq�P{��]�V䲝�`�yȄ�x ��20,�� ��ht�y�O�7'�Đ02���с�@���y���X�$Sd*�w�D�(�o�y�JP��$��El����-�1�yҪH��Hjfk�U��O�y�DK*# 0㒍X�9��"�;�y�Ċ�}ܰ�8�͓�"aؑ�y��#.����� �t�Y��C�*�yҩ_�s��t���	q�z�{�(��y#�<u]6i�� ��U��L��yb��!�X��v�~��s�4�yB�ʅ `9���|R��Z ��yRC��tVD*�$�)L�p���LŽ�y����%�ǸB4�t��$6�yr'X�Zl��w/r�R-=�HB�'x��S�;z�<��ڛ0DHl��'$M�5�̅Oz��JA�לtP��	�'x)��ǅc�� ���L"��pX	�'
d!��T�,��aE7^(�'�T�7Ś�	�Ij��7M��b�'TjU�1�^?U�Lܙ#�X�Kr"q��'��P��nU� ��̱���?�4��'@,�
��P�i�Pɐ�4@��X��'4v�j�/� h��U���8��X��'c<��׌�0�D$脀�2-l��	�'v(��$lϊD~V�q��R�$� 	�'.�p��V�Z;t R`��2���'%�m�`�ќG�&Qrd�\��u{�'�^�jp%O�H��`Ď�bĸ�	�'GV��`gO�n��q�x�4ͩ��� .�!��=X���I�g�E�B�%"O����N-~��1��ڪ Lv��"O2�wi��D���f�@0��#"O�Y�� 5����w��!$��8a"O��p��� �A�ɓfg���A"O�8D�u�9�J=_�8�"Ozh r&2>X�IF��z��8"O��B��g��'�_��@��"O�q���l��@I�Y��u�A"O�9KqŐ_V��B�¾	��ԩ!"Or�v�C�iC�QU%[�JŴ4P�"O&��0đ�x�F���D_�&�h�B"O���#M�"$���*��1"Oz�*ҩ���8(��`ݢ��Q"O����	H�-�~_�-�"O~�c�IpVZe@��OY8Q�"O�U��1cpY���H44>���s"O��c�R=r�:��׮RA�\� "O���0�T"0�Z"����Jrl�"O���&�r�����M�C�0`K�"OL���mbP���/	��@�A"O6�떷<95:���*�2�*b"OI��/ƾ�"=���P�'�*�`"ON�8r��4U���*�mK�v۪�!"Of���%Up L����d���"O,�8t���>�v��ΘC�BŰ�"O�=YF)���tuHT�]�F����"O���fB�%��p!���	A�����"O��*�M��-~���ߑ���Jg"OP��6kͣo<�����Gs�hXU"O�x���c��틠�Ȗq�P�b"OrM��Ӵ���Fћh,m�d"O�9Q�Ο�t �! f�<6wVhQ1"O��1U�IY����!��E���iw�(D�l���ˉWt�X�F�q	XP��%D�l�f"��O�����"� l5b�.D�ܢ���<.p��1�E�QNT", B�	�r�R	`�L��3��Go���C�I�^v��XOX��j�QqT,C��(3�p`R��p�hQ�Ͽ�C�I�KC2����͛1C�@k�i&X
C�Ʉu�$I+KM�.��;pʂ'��C䉘8��=���ϗ~�Պ!.��i��B�	�}�){�c�ZP�P�#ˏyZ�B�	jA�ԛ�Dܗf���D≿.^�B���Z�@��̄v���0�/�Z]�B�	��B-c���1�	�c��,�DB�I�M���ڈU@p�xTk�"|C�	PEN1sK�-w%��z���?m"C�o�L�M��BV���D��c�C��#d��@oT�dhP�g�'V�C�:Je�0�w�'#fH�I$� PA�C�#%txytj\������?6!�䜒 �˅�E�OP��F��;C!�DY47����� uԉ�ūÔ=3!�Ą R�= p�F2B&>��a��E !�D^"/lɃ��(C�T8�&(+!�Y�b��t��&(Ĉr󄉞|!��ZXv|�Q� �5&ځ�#B��!���,��<q�H�$"$�"7LI�P�!��K$L`��:�(�7�J'
!��^�8L�t tl[�tݢv`�B"O	a�   ��   5  K  �  @   �+  �7  C  �M  �V  Uc  �l  �r  `y  �  �  /�  s�  ��  ��  :�  }�  ��  �  F�  ��  ��  �  ��  ��  �  ��  ��  �  � � + � � @& .'  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h%��G{��Z4H��q�&�/5�Ph �/K��y� �g��ps`��&�ʈ*g�[#��ĺ<1ד.
��[C�56��r�8N5���ȓ<.���O rh�X��[�%D�d8S�3�ڰ�Cnʲ�XY��� D�(c�Ԗe�b�1MS�hʥO>D��#�!�0<�%D�B�`��W��W���s��J���BX�D#�DN_K�BG�:D�c�'<S�|٥��57\:\�&�w�X,���i������'K��Q�fܪ2� I4LQ�Q^����'�L��Qɍ,q���uj�<���'�DZ�OC��^}{ĤS3zxy��'4���|�ĉ0c��9��k�'6�����6[2U��FW�^Q���	ד��'�
)S��(�~��׮�!O�l���'t�d���A�� �fS�W���h�'��Y���e84�����T�4��'�b�',��j!H�iO6J�	�}��'V*��a���Q�ѫ�W�'8l[
�'�x 
dS2Y -�D�M1Ki�а�
3?I�'�a{�MO�W��}Q@ �D&��H�bH!�p?�O��년�m��݀b��W��Q"O�!ɱ.��pAH�Fsp8Xҗ|"�IS�'�rU�N�=(���>�����d�
���庤S�,�1�'��T���'A��I'��W�V���,�+�p���hO?�+ӠN�;\��t� �(~>���ᖐ2�1O��S�g�,��8��zJX"n�6rٺC�ɱo(t��-�fǄ��Z���C�I�ABZp��:U���bhLL��C�	����k��B$,P�1��_�p�C�;(�@��	�X�P��rb[0p�F��0���&�s��)y׭΃̊I��4D�� ^h�F,!C��KB��8อ�t"O�)�DDC't��YV-��iɗOB���g�a��TH��5�f}�*6D�l��N�-m�J�:��d���o7���z�b6��1�3=���Pm^,S�8�<!��T>����B:mp�)�5��=��Źs=�hO�2+v�ccL�l��Q�c���} rC�ɒ��xYb��1�!"V�f-!��"�S��?��&��4��Q)��F�\>�X��o�t���hO�''�
���+�2%!�ix2)��^Ύ=��Sf�ܚ����-�8�5��:,���ȓM���ؓ��WH���U+]t���*=!�Eع}�|�C"�D*��I��ٰ?q�n
����l?͈`2@H�\?!���S�<Ld��W�G@k��zq$��C�	9("�qJ��	�	!xt 1��%=�4ʓ��	VX��0"���%��kq�ߨ8��
'�,�O��Q�h�c�NL�N8!`��'L�j85O�,J3�ĸA�xفA�Q/%bi3U�k?9��)'?��W���d�E������q�2D�P��I	z�X���]� �~LP��+�Iv����k�r�#qI�>C�­	 �ۑ��'�a}ra�~
�yQ�Y�sZ����fʴ�HO�b��n���ĊZ�pݚ@ ?2q�S�Cw�!"O���㙏M�"y��ƙqXL����xb\��&�b?�9��X�e�2�� �M��92�?D���	�Q����F�q�j�K�b}��O2�S�g�I�\��hZP���;�\s�)��C�I�U����G.�+Y,��s��ǋ�Z��hO>�y���c�LX��J�R�6� �8%ax�_�g����e��N�XzE��yB�GT�:�#c��u�|����V���Ọ~n�U�J9�҃ɴFz0eC���w����>iaʚ.�r�!PKR�8�΀��	�N�'��?��cϋ�~|��A�
]鴱z� ��hO��-E���d�J\�5��&X����H�����L�ݠ"�^$
���d�� �AM�M?!�{2�I�r���HB��ʡN���P7JY`}�dP_x� )�' ��aBc��	����9�R	���M�)O��AdfY��id�Aئ�����>!-O "~�㭓�oq2�fL�����S,ԏ������p!��iS0���y��5gn��e��_�R��(�b��d(#
ٳ��?GF��T�x�'iɧ��x�ĐN^H0�w([}���a)�Od�=�O�t�-�y�Ly���"�6��4�Px��W+:�#�늰`�l� ����Pyb�Ƒx��p���*j�B��kG�<�2A�v8���*H��@l�H���<��{���)�*Hb��̧CR��i����i�v��*���K$@O;�����L�h\��'C\,#�B�;!�*SȄ�;y��#�'n�("f��(|�(H0���:�'śf�	(��c��=%�y��/�?�y�*�&jׄ)!AK'"��Y�B�9��O��Čs�IK��h>,��j��M�帗Δ��yb�����Ą_�q��`�F�	�y���A�8 	U)�dF�j��@0�yB1~�@ �]g�:a�`.���y��C�nY|T��-Ɋv¨���+]	Ρ��K�R`�P��F��$L�1�1OH���?y#��NH�UZ��OE�L���6D��K�X&5�:@iwA�N/$�se�<���5E0�)H!ȅ+�	�p�Q4=��B�I�5X���؍8.��
��(�
B�)� 6��l�.n�y��#X�ڥ��"O�}R`�X�=j,=�b�l�>@ "O>��%�/N�z2��_��R"O�E�C��h�t��1�ة��<�tO&-�C昸O�\�cFɘ'`��r�C-D����7�`���D�� �I8D��ۧ�J�C>�rPc���8D�"�
��~�B�yDM�9N�6�	�:D�p1��:��\Q#H^?&oV%�0j7D����*��ST��/
��BTl0D�4�fDđYU�U��e�n1J /D��i%�m�>P,��t��+H�b�O���$W�Cw���㒢0�fm"jC�x�ip��P}�CL
�f\�Ď@F���Y�y�+�8~�=�� >E����׉���'2���}������@`���ѱ��)f�!�dĳt?^yZ%��Do����n�'p��]�0nN~ʟ��~���H�<_�|�q�N�O�
��D�/D����R�8!��>`��dƋ���'e��Y�x�Ј_8�|�UL�KƂ�@�;D��s���4v5�ǉP�jM6�i@e�؅�I*p�Fqb�=s��ɖQ]j6M.�S�$�$�Xh�	[��1{���SH�kJ!��1_�4V�5%�p�\�s��<��E%^ɛ��62�#�+-���AK���K�-enQ�7%ս-�؀�':1O�}���Z�p�M�@(��� �95���ȓo3�+s��h�
y
r�9�����ٰ?�@Gذ�Μ鶉ΞW^���̘B�<�C�W�g>���V���wsŕ`��<��+�Ef� �FSZ�ZmQ�%�u�<�b�K�<�� ����T�@�����[�<�7��.
�8�f"
�kV̤pcW�<�7�.c��AbDKǙ]��͚|�<��	�j�X��$Ua�tc�Cx�<���G?m���Ũ9!.�!�,t�<�GĂ���+uLԀ�Dݢ��Us�<իT���֧�:>̺d��Qn�<�n[eP]���>�<��a\A�<Qs�E��.C�G�-2�f�9���<IE�3W[>=Ze��,2�HX���^e�<�`i	y`ԉ���*{�HГUK�c�<���(N6�"B��W���ӳ��I�<	�j�2ԐQI��0I���S�Z�<�e�R�"��Yc�aF�8dZ8aWiR�<��H��s��0�!L��|�D@N�<��N�� ��!3͡R��X��r�<1 . <���r5�%���3�MT�<���_x�ܐqr*��L���p`�R�<Q"��@݉S��:�,iPЮGQ�<)���RP�M"���s��H�<��$"r�,ه�� (X0HI'�ND�<'�Ƥ�0%�v�ѻ#���A�ΙC�<)��T�ބ`RIڱ2�VE��dH�<�5+/l�H���/yzr!�ӃBI�<iD��vI���4�Y�{��@��ƏP�<!2�[�Zp��ԯϣI��ˆ��K�<�q
I	����E8j���O�!�$�������%(�X4h��T94C!�V��5��K��!�e3��=!�!VkZ�A�B̉5��e�#.Ҋ3!�ùK��p ��J# ���3bZ9V!�D��V_
A!�Y���0#��m!򤋔R[6�"!�D"��1���	!�� ��ԇ�y.�#���v	�e�3"Or�bq�R�z�&�1p�� �b��"OJM�q��:6l�8�UꋳY�� �"OZ����!S����*�"�}�!"O�@
�/P4xbũ�� >�f�@V�'�r�'�R�'���'���'e��'��d�\Jj�Q1�kW�9�>$c�'���'�R�'���'f��'��'��A!�O�-1�0m
@���G�Ĕ�r�'���'�"�'�2�'��'�r�'�d �E��X�9w�� :�,��f�'���'�"�'���'�R�'�2�'�>��@t�����ڧ5�����'h�' ��'���'�"�'���'[��Y��H���k�K�6�8�'���'�B�' ��'�B�'��w�&��RG�<.sL%+�Ή=oJ����'xB�'�R�'<�'"�'R�'P�9�������D�74�C��'(�',��'2�'���'I��'7T���g@%OCn-{��ߴ8;���'b�'%�'���'���'���'�b����[��Q+�L1�8)j��'W��'���'x"�'���'�R�'Y�Y�!-rL*V�v��AK��'.��'��'���'Db�'�B�' ���7�p(S.Ʈg�mX��'���'���'�R�'�2�'��'� �!��Nl��f܈u?6�g�'�2�'���'���'��#|�����O>�0i��$�V�;�nF/�½#oDky��'��)�3?�4�i��T�$�s<����V�e=NQ�h�������?��<��i��(��d��E��L�b��/���b�dlӲ�$��+fv6m"?���!vk�� 3�"����^��͒҈Ի	�p�0�G�Ҙ'"\��F�4�ח:k�!���"G{B���:�7m� f1O��?U!�������`� ;�A�/�.9c��H��@~���l}����I�O��6O*=�#7��lb���7c֔��0Ot0r,A$S��8�1F-��|���.�zA�w�A�XRt���ɍ�{kv�ϓ��D.����r�-�	eo<��fO*3���@u������?	dS���޴4g�F2Oh�ywnQi���3�����0̌�'M�=åi�&xl�p��$.$C~�΅��$Y#��!H��XB�V?_���Ry"P���)��<��Ę�N-�:a�)�N��`�<iձi��1�Oބmk��|�㚄"���p��ӻ24�0����<)�i.�7�Ob�pS�kӾ�-4�Y��7I���U\8b��ï+��u���������䑂Bľ=0ÏL�O���j6�T_�I��M��*թ�?i��?y������\���,�/�հ%M� g��E��FyӠ�O1�Ph��#�5N�,�q�C��g-Z�з�
r��@3�ͻ<itB�*}Xv�*��\�p�8���WqI>��䕨����G�Lڱ�i�c�	3���ITl�`� �g���v��5���1B�xr��.|��ZO��F�tӰo�d�����28[��yc�8Y��	GC˕h�L=8�ʄb~���ӧT�z �,i6M�Z(Eq臏;�x�d�Pk���WM�V�Xc
T�KR U��ȍvM��0�Ҩ%��_ W����Zo܀91�I�"���˂ p�L1D�'�D�r���w���it�C�(1 0�E:����-\�t���$ h�R	x�f�-rg���k	7���l�������%�������9��~?fe�m����0��.�6��`)c}��'�b�'�剙{��O�bHA4c�4	�QD??�R@k#��*q.6-�O
�O���O U�WC7�J��E�r�C��$hb ��
L�6-�O��D�<��Ȧ����O����� ��GU�x)z� �z^�c��^�	����I�"x�?�OZ���d�1Z����n��F5�H �4��dZ�FX�d�Ol�d�O���<��p��+���B%����"��B�m�����	�wx��?�~�&Ƀz�th�.�VH(�3-���
��ɟ�����0���?�'��'/���㜟#-� S�!P�!���3.x�ι+C�%�)§�?�pNR1/Ì���F"fnؑ�.9j���'��'nx�Zw_��Iџ���u?�@fN ��=����`�0�H4�r�R �d�I>���?��9�0���Җ r�{��-2� `�B�i�!D�w��I՟L�	矰'���}�d��4^X<�d�^�Ml�JS쥢H>����?����dϠ<��$X$ եO�h0�.9 H>���*�<q���?������?��n��a�ڴf�r� R���3����
!�䓫?����?a.O��a#�?����4����@�b4��&�iӶ��O �D(�$�O��߼���:!jJ��P��	�:="�̄��8�'r�'�V�Ȫ�D�g���'��-r�*Y&��Xb)�"\-T�v�X��8�$�OZ��F�c�2��+}�f݈UzIc��(z�6�P����M���?-ONi@@�|2���?������*fꔮ2�~192��Պ�R�xb�'?RO�n��O�S%<�v�R$�3z���ہ	غB�7�<����?9���?����-Ok׎4�1�&��6�� �N@����'�2fE"��O�����Vǀ-��с�bƪ�Q�irL�	r�'�'��O4�	�,�ɻ:�0���藁 &����+?N��ٴr:nz���S�O�R �l'��@����i�\A1�(Ee 7m�Oz���O(�)���`}�S�T��c?9�mUR������-�u�^�.ur�J>����?Q�UM� >��A�l�$��		Ilqcs�iBB�Ev�8O��O��d�<ҁ��)7R{�材/�-��)32U�&U����gy�'�2�'���s�q@ee;gA��!�>�$	��*��ē�?��?i/O��D�?��ȇ5JG"�i1E�
^V��ZPv�B�D-��O�d�<A�k�F�󉋳`/�P��aQ�&��pt�E������0�	��'��P>M�	�H����ƿyi�}�vC(+�ỨO����O�$�<%B��;ۉO�r	�^n�b=�F瘅Ŵ���E}ӂ���O�ʓ�?.���=��N�2LeZ��Ԕ`Υ���M#��?�*O��B�N�Y���D�s�aU,M�ӌy��0�Ve�Cmlӈ��?���?I����<�1$�p���%�O[�8]��lPK}b�'��U��'���'���O��i���u	�n���a�_r�Y!~�,�$�<i4�u���'J�:ջf��r쐙��!l`��oZ�<T�8����x�	��t��cyʟ8�+���oBA ' �	��B}�坿�O>ey��"AJ�H�i>#U��r(�M���?��s�h=-O��i�ڕQڎ](�� -��(6S5O(^�Fx�:�S�D��"�j��6�V Sِ�3 �\ }՘�m�hP�ZRyb-�~Z�B��&Q<ܻ�R?�f��_�|~zO�0#����O�ʓ�?i$I1Q�:pYu"�2�0�k��,-O(��O.�$��e?�uKC3r��=� A�-"�:1��O���`���O�˓�?	�G����Qn^`� �V��%�HХ�M��?����'�	>Ў7��=�h������i	ʉz��I՟T��ȟԗ'tQ#�2�B!�@�ā	++��
��>/��m͟8��|y��'5�����O7�U��a��(�T�۩����gӖ�d�<y��{��\�(�����O����*� T��.��AP��T�x2�'��.��"<�;
>�@�k�E���4��n�gy�� _ڠ7��o��'��$c:?邊F�fD�ԉCr��l;ƁT����П���ݟ<�L|���i��`�AI��<�@�D/g˂���4B������?9���?��'��?e�QgB�Ir��[q��Z3PE���5\{�b>I���ID�ʆ�׹�6ěm�-����4�?1���?���Jr�����'�.۪i(*��q�&>`4���M�-�6��Ol�$�<AEP?�֟��柤���q�F���&��E�)H��M���z/
���i��'B�'Ӟ��~�mL3"4���G�/i��1Ч�6�M��k:�ϓ���O����O��D�O"(b�K�}d��B��&�H)����$�-l����I�P������<���|���*�1�<���)V�Q���<���?1���?y����i@�2j�m�T������Y7�bj�c�$�`HX�4�?���?���?�+O���S�i>R���m�/H�� V�ϩH�)x�4�?9��?����?)�1^x6�i�2�'-�r���7����R_���q�����O���<y��4p�`�'�?���<lYǭ��r��"̨T����w�i���'��'��2�{��d�O@�$���q��bV�=��T��ͫ=vb�b�
�����ay�'R�|ɘO��V��s�>m9�HO'����˛K��s�if��'e��
�&s�f���O��$��"�I�O0-B�/�ud=��ǛM�z�@"�V}2�'7��X��'��X��o��޳F�L��Ȍ�56=7lL>�?ASG�2q��f�'��'�����>	/Oj��2M�	"I�� _��j#h�ͦaH�j����py��I�O8���J�Mr�!��;Ixب�ަ-�I���	 |��`۫Or˓�?Y�'0�4�0	)�bd8��(���ڴ�?1-O��8O�ȟ��ϟ0�P�6��=1
6Z�0��nD��M����]q�i���'�"�'0n�'�~�M ��|�&�#��$�������y,1O����O���O���AƄ8�E�#UID@	�� �"��:�LWæy����<��ʟ�j��P��?��U�8��	4E3���4B5����?A��?I���?)���?9���6a��*�2����%,\�3�6�8�CB���7�O����OP��O˓�?��.Z�|N�	Sz�#�������Vy��֟�����ğ��D��;�M����?�0�1C\`����		I��Mq�#��Zu�v�'�2�'Q���XX�b>a�	�L��gI�=X�@>u��pH��M[��?���?9dj�Px��'���';��eO�`h0*"�Z�Z��:�F�M��7M�O:��?C��|����4�����2a�������!GJ���M���?�VZ0f���'���'e�D�O���$�5	�@�g�F�Ũ�X��꓆?Yu��?�-O�ʧ���-.2�h`ɍ�z�8LA� �oq�6mٕ.v�mZ���Iޟ����?1�I������L� ��ǎ�}�lɹ�(i+N���4/�И��?���kP��d�S柔�ŋǢ	���ǋ�~t �Y��-�M����?y�n�Z�c�i�2�'��'\Zw���ʚ�f�*L&b�  ޴��3�t��S���'"�'�d|#����X���i0j�NlU�u(w�$��G��`n�ӟ���Ɵp����ɱ��ZFkܑb9� ��C�����O�>�eN�k~2�'���'f"�'���	J�d�E"A�a�A�t��T�i�����O(���O�=�O�	�y��N7X�Ȧ�W�`� ���0J�Ky��'R�'/��'ݜ��jlӸ�� �M��׻��z�m�2tA$�i,��'���'�2]�<�ɴa:��S4(��{��*��`K5�hY(�O|���Ov�d�O��d��yW`�n�˟�	�'�݋aP�[��+��	5�����4�?I��?�.O.��ӭf�;}"�@e������;�B%����M����?y��?����o����'�2�'�d�\@Xщ/M�d��S�ȔM��6-�O��?鲠A8��$�<����boԓ�.e"���t�LMyWJf����O��f�L���	���	�?y�S�$l��d����D�(UX����2+����$��ED����	ry�O�'R�����#T ��w�C�]���oZ�YtB�#�4�?���?��'�*���?��}^p,qexD ��I�V@82D�$�M�Ы���D�<�g~�O�2IF������Ɋ?��(A�'�/1Q�6�O���O����&Uۦ��IğD�I���i�Mj����-䪉�Vv�p�
h���D�O��D�zl�?]�	��\�	2�I	�A��s~L�5���0��4�?ёBC�����':2�'[��~*�'h*9���Y ���T�6���[�Ob��<O�ʓ�?���?y��?��c��qn���~(�m�b�)��p�p�i|��']2�'���D�O��n�`o��A4�bpP�ы@ ���ݟ��ş��W�DNSY�7M�J.�ؕ�EJ"}j���udf�m�����	�����̟ �'�Bn�=�����M��̚�J�X����dG�gѮ6��O,���O���U�4�_n�7��O���U�E^�C��2@H���k+��]o؟|�Iɟ0�'a��	���TT�`��@��%��rc�� n��iR�A�M+���?���?Qe�M	SH��'	�'.��e	4?��(B��
 j��2g�ү�*6��O�ʓ�?I7	 �|�J>��]PЌ��ʭ��J�` )D�eӘ���O��Z���̦������?��П� 7+���Pj�!T���!�\���D�O�`�O.�O�i8��,M�o����U���K������Mca���v�'���'���Ov�'�零4~|34e
Op5ᵉ7U�7��Ѥ���O4��|�J~z�?D��d�Y׎� �!J\t�Z�i�b�'�B@��Rz7��O����O��d�O�NJ
=��sg(߇)H�HR�U�9����|R,۹�yʟ����O��d?l�X|*���,���óI�q@0�x�T�dő��y$����ҟ�'�֘�*��,��,g:��"�)�h�6�lY�����O��$�O�ʓ��l; 	��yRA�ƍ"�4!�	���'GR�'��'FB�'c�]ڀ(�yD�)�H�&�"�S����y�W���I�p��^y���bR�ӎ|ٹ1bL R:�⅛�$n���?���䓒?��YPx���$�{�f��T3��p���/L��;�U���	ߟ���iy��������qG�I�n�9��P�s׺ #�N��-��i����(�I ���IV�$��,�Z���ˁ�V�<؉!�_5+��&�'��Z��;�+B���'�?���$��ې���� K��e#���x��'�+Ԣ�y��|�����HL4G^pP�Ы�]p�Y�i��I.$=��4/�S���ӽ��D[-7��m:a���$��laŠ����'&r�N�#�r�|��T&h���׀E"P"��S0f���M�5o�5<��F�'���'u��>���O(�%����<Ēǡ�$!n��A즍ↁz��%�"|z��df�AR�\2��@��Z�hq�	
�ip��'.R�P�F�dOR���O���x�.� �#hޜ`�W�r`79�O���,&>a��ٟx�I�K����I�1ͺ���^���X�4�?i�&��(9�'A��'Aɧ5��-%�a��Z+`��H�a�6��d\:���<����?������1���'A�
oH��� �$�5�⃔N��ҟ��	m�ҟ��I�yJ�)���1Iњ���ӄ6�����/|��'R�'\R\��8#٢��T��B��\{�=z;�T���۫���O��8�$�O���R�\�D!^�:�᫁��6Hb��Q*!�'��'�BY���Eؼ�ħM��"eD���I��� ��T���i;r�|R�':�)4"�>��ߩr`$T���M��m��%��!�IП��'�Bш�4�)�O��	ݩ��� #��pj�*�d r &������<���ٟ�'��3��(j��B?E��	�w�@%i��m�Xy��$��6�N]�$�'��4�)?� �,M��w�4g�}�!�Mڦ�Iڟē��o��%��}�EjI4j�(��K.$�Ē���ئ�� K�2�M����?q������?)���?�-�lȠs���l����Ɂ�)V��̃�^���'C�i>=&?��	8��H���M��ĉ��O�!�P-�ڴ�?����?���ש[�F�'��'T2�u�\u��!�#,q� j9^e�m��4�?I(O�92:O������PzRB"�L�{q/ �;��A ��Ʀ���K��{ڴ�?���?���tO�w?�3 N~����a�W�x�H��
�B}r����y��'���'�R�'��a/JP�ŶI�!ᖭ�N�6YB�Dž�M���?����?Y�^?�'��CO�O� dV�6HH@֭6x�.l�'�"�'���'BX>����MsR��(H���R�����*5�B�h�V�'Sr�'��'��ݟ`+�n>y���

H�0��`�0I+寋 �MS��?1��?�_?��vg-�M����?AAR28���%�$w��m�4Jڇ�6�'���'i�؟<�#�>��O�5z6��$tIj �f�
_��u Ľi�2�'���'^��tf�����Oh�D����� F�hĹ,���	�d2���i��\���ɸ���s�i>7��(����f	�v���$F�#!Ǜ�'���K�eG�6�O��d�Oh����2���&BC�A��f�7(N
=R��R��00�'�B�J�4��|�O��+�t���=k�`-��]�,��Umڗ4����4�?)��?�'�Z���?��A�\�w�O�������Ҭ�Rӹi�9[��'�rP���ģrӬ8��'�1~re+F!�!���Ё�T0 NȒ�`�+Z`<�����)��%��	>Wvs�șL�ܴ�TOɂX����Y%.�T�A�i��Dp��	o6�ȳLF>*�^��DF�!V�VIP'��35�4#k��XH�L�{�h�NM(��)�o�4�ĕI@�ܛH7�Ei ���!�C�Y���m!Š�(<J�h�lZ�+��q�1�ّ\��)���FT��B���Lz%�ڴ+�L�����DX��'}��'h^�"��'��1��x 0R'�t����`�$Ժ������D1%���� ��Ox���ŀ�*�>��i\<kZ���2kN|i��<'j}�fXtx�t��O`��",$�TX�	œ0G\Պ`d��R?��=я�$U%+" ��`J�t54Lp�F�ax��	}�h���m�w�I�Ah����"�M+����Y��l��p�IQ�t��$�.A�A�`�(�����Fe!"�'"�'O|��T�X��na����W՛�� ]�N)��"ɡ-,�9�P-S�u��eH!�?)�Q��2��E�=CT��_A�&e@R ���ᎆ-@� �~�����- �B��B c��Nb�����O��'Ae��9]�����.|�5�GQ0�?����?)��?�'�hO`T{�f�<�`2�eգ}Uؑ�e�'T�O���ňpޱY����eA E�;O�����]���	ϟ@�O��Q8R�'��'u�В�&7/�JT�DMM,&7���UF�6S,��lH�o�t+��Fezh���,�1�g�W�d��b6ʝ"R�P�*�K��]v����N�:v��b�/�1Ҫ��6�y��#�N�(���ߑ�f�.'*}����p(�1�)k� i�I˟(�䧝�+.}k�F�(	�#�I�	��܄�������X�
���1)F�mYeDxB�4��|���4�D�
���8M��ȹ�!۴t �����?I`ʉe�hy��?	���?������$�O��D��������W2!�� "g�O�@9gc��L��8fA>,O��P���k�P�����Db�@+��O�*G,ɌF��{@A4,O��တ�N���F��!��!��O�|��'m��|��'cR]�`RUj]+^��4#nM_)L�9��"D�X�+"!y��X�0�H��_��HO��_yB��_��7͏$�j9��]���3um/q�����OZ���O^��5��O����OʵZfkX�N��Ab.2LX�����Y�(]f@J�\r8��C��x����?VhQ����@��oR�p��ƪo��"��[�u�`!�� άU�|3�`ĴF;H��X�|d��?��L��<�	
�u7.Ձ��M��2��@�ǂQŦ}�ICy��'��O�ӝ�A���U�ͥ(ɾ�h�����,E{��	.�L98�M�goDJ�oы_�$�̦M�IWy�f]qd7M�O&�D�|j�M��+r�����vpH��tE��@�x<���?i���֦�:tSR�ѱ�>4�F5�@S9l��5% 
P|�b,^�U�F�[r�Zs��<����e���0
Ra���[c$Q��uG$M#^��A@K�(���T+́q@��%�	�i<��]֦3����*ά���F̤FK���Q#ʹ�yb�'k�}���#4=h܈�U>�L�b��0>q��x�ɝ9w�4 �B��8.-�q���Q�yB$J�-�N6M�OT�Ĵ|�P�Q��?����?��Y�<,x��KV�p�JH���S�P�j@$�3=���q��i������רd�L����w�P�	E?�������<.�|8Џ\`P�la��ǁ7a��d�0����+Q lCH~��|7,��F �����3"n���WÂ��i�4h\��`"|�	$,����f�� ��9x c��	��������
�n�07o@�`��J(:�#<��i>��ɉz-��DH��<�!ʓ#�fe�Id�gmԢKN��Iğl�Iҟ�
YwM��'*�l��J��\��Di�K�]��,��'N ]�� �|x�PC�	]�MP�B� $|�Q!b_�%����v{��!�f�l��	�t�tXE��_h
�C�Jϐ%�ɄTe����M%���,O����<Q�@G� }���U�}�J\��D�<����
]g��U�𰖀BR3��iW��%N��<Q#�Q�	K�E�#����nL
<%�$�7�O/dL���Ov��O��H�F�O �dk>)įЦ���$~6Xa7�I8F�D�FoϳMF���d�!
���` . Gn�4H	Wg�	��I�,и�$�OdlSd�L_zD�෥��\��К�D?���O��D:�)"A�N���Uǀ�p�\P��ng�<�D�`��Ih!''u�^d
����<��V�x�'Z��X�m�X�d�O��'�<�1d��7r��Q�#�c�1k��?��?�6�}�40(g��b6��4�@�k�.�6.0@�K�;6�P��'0�\9;��ݫEU��9[M�B�2R�iTش�!!~Ƙq�2��XLж��I��GO2'#�t�З|�gO2�?i���?y����� �|�dm�8{�����ʍ&_������On�"~�=���%˗$l5z��P,���'Aў���ē5���0Pi߃T�j�DɥEQ���PX؄��i���'J�Ӟ0���I��,�I05%(���п	��!��˛ RFDc�9�}:#�_�h�d��|���&���*��3�;!�3y�`�ѱ��2 �\85�2��S��?��-	&�"���CT�%�Q`�0OZh�*�`h�6��<��V��?�� �,n�豭ޏ�|;%���<����>�4�B�!�6(q�8��t`F�Be�'3�#=�,�dbth�j���"$A'_�Q����Od�䇆qX��n�O��d�O^��{��?�V)�zr0�S��L.E"�];tkG?	��D���
ۓZ,L��
�G��̊b�J����$8���'����=�C�(��s�.��%��� 5 ���\�a�I����?��?�,OF��`dZg����Q`�&$�ά�4"Oẑb��4cYR�#�JeaƵSNS���i�<��f(���M�2t��D�ጵq��ذvj��'�'Ꮉg�'��6� a�蜹B�I�&.�-n^`� �L�} >��C]�k��=� 	0��G���(O`���EYY�j=��]%14u�&��� ���v\��`A?^�\6��\��?�тR���I#;8��� f=(ܹ��ݟ&y�]'����ڟ��?�O�9��FT'D:]�Gb��pIr���'�v���Q�kۜ���I"]�����'��6M�OX˓n�^y�%�i���'���r�����oӑ���E���m�J����^̟(�����$
ٓ�8��-[	��T>Y�4���L� :0Gۏ��ԡ�E2ʓ0�����&~."������_?��2�a.hf੔�Ф�(O
I���'g�6�H���_����m{��d	�_s"ɲpR�(b��s�X�C�;�f}�DCW �Z��'�)�O��'���ả(i��uR&�ԢW2TX���f�l��(W�eJH!��ƟĔO��THe�'Vr�'��X��K��?��� ��� ���r�.�?��Aa� sV��	��F����q��qpdQ�ɂ��X��h����./�X���41k~<9(ϵA5��~�	7HRl��ȍ�jc�ax$�xYRp�4�՟��4b����'�?�dԛ{.\E��eJ�/�jD����VA���O���$S7��00�,�e},U8��H�$?��r��L��~2�F'�`Lr��E�<�R��G+a��'ͺ��{}��'���'�P�]ܟ��I?5|�Rt-L�?�"� �U%�l�I6Z�L(ˋ�����'��dp�EӉD$X�QD�� H_�X�'Ɉ�[L��McD\��q�� ֬�t*p�"וEOn�u���@�S��O6<n��Mc�b#�~��,���J �ߩ*���R'Hc�<	�����艘�-D)9���#
O����ɫO4�Hw�W�Ҧ��0%�����Ւ���A�L���H�	�l�	/o�>�������'+�Vi�EN  ��Y'Ӻ3Q"�"�ꐺx����
��\�=:2�O5��OD�;$EW�7l2Q��[�u��=��%�9�V��V��8'�T	q��Y#3��?I��[�D�4�N�rO̟S��1�g��$d� ��?y��?���?����䧋?���*L�؛'��Q!.t
$	L�<�	=�8!��l^�U�QZ�I�<��R���'����f�<���O>�'88|-k�(P�.�&����K��x��o���?����?1�A�o�l��y*��P�.��+2���W㊒
u����ɡoF�ȳ�6��9Pb�mQH�	�L
�ڣ<�`�]ן@�IB�Sß,��fV/p�ຂ.Cz~�!�A�Zӟ��?E��'K��� wN�j�	_ m�j���2�'�|�b5n<B_쭓��	Yh�M�'� ���~�\�D�O�˧m����?���m'���[�K9��{�
�%_E��XF'�'���	g������&���2��O�IВ�T��vё�_q�J��g�\6�� �� ��1q�i�П"~�	$���X�ℭMH䗼+�P�eI�l}����O��D�O�"~�I�~~�#�oS1|Ϧ�[SLV"sr�	��t����av�yX%��g3��hv$�Pih"<)��	J�$�a���X�hX6-�6|�"�_A��'~8�"/A<-���'���'�4�������9�*�q�;=F@�cGF�`~&�+�/�Q��Ғ�ș��B��?1{��͔VIH�0�/I�h��	ض�
��`V� W�D���(�_:Y��֟�$GyR��&<heJҎkk���Jҁ�~2KS��?��i["7�8�ɐ���j����yd���F� 4;�I�	�'��ՠ���,�%O�њ&6�EzB��>�.Ov�U�\�Q��KJ5D| � ��2'�f�*We�����Iٟ`�I�I8�}�����I2޺h��F�/~ؤ0b���z��-����X�D��6m5�O�IZ,W(F��,ځJ�u��Y��� 6���)� �R����`G��p<�S��ܟ��	�5�Z a�7LӶP(0ۊ|�T�C۴�?�.ON�d:�i>��)� \t���o!6���@ʸ<�ʍg�����$�R� qcNR���p2B�3c��$����ݴ���(-�f�n�����U��;���c2Z;Y�<H+U��K4�Z��'.�'�%��W(,�~u���ʧZU���=}�,�� �ۿX�� FyR�B�l9��Y�%�&��On�� �n˸�.�Hˏ"�T���D�9�'��Om�-1bUZ�1W��>Ͼ A�g�1~����s�h�q������͌�w6��<�O)'�|�VmLw�I)V)	�¹��C ?Y*OL��Ւfݤ���ύ!r@bl"�lR�C�!�$˘�Z��S�3�T�r&��:�!�d�18
�`��)�r��5!@�?^ !�䑺F�9
B�ųQ�n\1���>�PyR�X��=	�m��\EF\q�$_��y�J?dI
T$
�fV���5�ybǞ?�t8q(�+a���҆���y�iӓhx��"A�Q�h���͕�yg޿"=��Z��"J����A
ǔ�y��M��ya����I%��Rq�H=�y��y��)�'߻wB9Ha����y2��*<��'k4�8FZ)�y"i��4s�h�S����)���:�y�.�b�4���`߇{�L vO���yR�.Q^�УL�JI�z�B��y�IC��Ʌj��;���ĝ�yb�_��"O�"*�MҢ����y��ȡ<�4TASA�= �ݣR�M��yb	� f�00c�	OΔ�ȉ/�y���h�>��l�*�,�ԟ�y��	�qx����+�>m G�B�y�
[�0)�H���U�^L��CP5�y2C�� ��y�F�b`�����yr�גH���ڱF�����	5�y�S(d�nM0�+�"�<�2'Fȫ�y�	 ���Ц-et���̃��y��5i�pԺP�°o�jL@�yBhY�P&@�E�TL�tA ��p>1���O�<X�*�!d���¥/\�:���+8� 7��ݸU�	��g�xoH���R�c#Z&���WE�>d�"�$ d �ʡ��>4L���"u���'Ϡ4�)�/;$H)��,�;j[j�Q�Z�}"����%&�L	�R`����n�1�Y`���o�6@��Q,n6��*��?�?�j�#���6���	���o�����}��%�4z���in桹$%��ެ[��XC�������qR��AwA�|�	?_&��H�F��>4��:������ƑM��b"��SK�[U�����4I�$ȣo�Aa�4O
�Y�]�4˂=�"�t}R���3<AV�i�䛧D���A�d��	q������S�'V1{�J�	�(������99�O�`�e�Z�����&UYRY�o�'���S�@��qڬ��qn�*��m.���I�	�1Z���uf�j_�l,���K�kħy�Jۓ�轊U���R�����@����E�2\\�� �M�����L	U�Vu�C�V-�8SUcm��RI�p*��ֺ\���+��̊��h��xb,�=C~�5�Sϓ��`t���F���c��V}�V�I��LBd�i��(�j��0���chO�s��@i�	M�r.���ˏ^�'����茕uКi̻K|��Y��6A����A�;:�:�͓EXla�O����)�~H�����O����� ��%�X��`�D9Ȃa2����`�zhTw�'X��сǄ6���r���7ida:��O>]�pMjߴ.���"�̟���	�1�2�i��b�i�(c��1;R�
V��%Q�
�0Ҥ�c����]�y��KE�P�"H� �Q��
�T1���� u���$�<��J�'ž#=����D4LP�Y�a��d���[���<���LQ�)�Ӆf��@s�ҨlW��(����B4�]j	H-t.�Ȋ��H�2��9)@Kl�͋ӫ��C��P��|)f�)�Mh�(9�	�(E�LAÓ�>�~�"lN�5�=����$r��!�h�
&bdـ��T�l�0Xy6�O�	���{G��U��};&�5l]�%�0��*Eߎ�'��dc�E`
�oڮI�DYS��4h�O�h��K]X��I���U1�L��w���*8�4�!E�$hX$G�D��(O�t8�I0��k
 �!я�/#�hҰ˱D��y��R8R}�`�6�M��4�	_�����(*zP�Ն�Z@#��韚����h�q�� ��hW&\�2\���nD:�@��[ vd�1��7��zp+©�y'n��: P�"´3���v�%�y�"U�"M9������;
�̰�H��/°�p�a��=�t$�RbH�6��	�=V搒�$[�a����,�q��m��Q���h���(��dj���)iP��'����LýR&�z7��YM��O~� n⩳�!�0�+ 'Ҡ.T�M�.�{�P0f ��F�2,���InC�睭r� Y�l �R��ГD���2���(�
�J�)Q�	d��+'"����gy�'�|�#�ᅉn����
�5K\ U�/C&�N�Dzr�U�n�k�*�~7�ыծQ�S��|ҥ
K,}�&��s��Mkp�~�	>9�*t�it��C���y�WQ���
�*Cc���F��y"ۊ(���=%>��N�,�xt��
6�z8��n��$�BP��CZ����
M�4��p+��L�BZ�NB/q��g~2@V�N���M�,���*�J ����hٲ�9�V2&����	�S	���[�Ow
y�B4 �(b�ύz���p� �7�(E����a��ݪ���O.w�<
�ia��	!6�� e�F?
��FiA�r�L�9%̖�_ ��C�r��{2����C7^�@�@�4A{�b#�ѐ�(O��S1@�D����O �|�ʍ�Mnf�B�O�i�D����?��nV
Ę'!�9�'DT��2�[�y��v;@C䌘�6���,�y�N�hjWI�!m��ɰ��x�'^�tx�o;T3bE �)9&E���u�	�|B�B1+F$p��aV
:g�a��/�H���$�07�p�A�`Qh����	w�{���4�V9,�Z� �t��Q��A�>H�p�Ӽ�u�׉[�vi�q�عq֩R�Dƻ�x��Af�&YG��si�
u͑�֝��y�D�?|^��%S�(���S�e��u�$��S�yY"��2O�1S�I����)�qw�m[�m�������(Qp$��
!rݚ��`;�>Z�!"�$�A#@�K��mmz���&].�%憷l�P ��f�Q,v�{�&�{��Y�P�=-�xQGb���!q�Z��M��j�75��n�|�t
�O�pY��20�F�!���X� 0���-�C#n�6d�<��O��s�Ԡc��6��� =��i؄$�j�Pd�]0e;>�(p\�$kP��(���U�#���0d�?x�Ol%�5\%8*�swa\� Yd��%�FS�T���'��t
�Mޏ|����DX�"<2�e�~�w�U#Y	1��X���{,�b��Q���'��um,����	NT�=�O#���0��/	��@��"5h�i[��,��ܻDV4�-S�ꌖu��4яo��zy2K�%h=� r�!�b����� �X�ҋ����	S,n���:��<��	-OY`#��ҡ@Y�0p��3vm���!2��=K�H#7�=b�b0�ɑ,Z��!�uG$\�v����%;fj؈Ijz-�-g\�9�M�#&�����Ǣ5�$]�	�s Z$8`f��-��[qHڵ1V��� H��D��p�)#8�ԥa!l���,�I�O	V x��C.�N���6~��!@%R�%�l]t�`k��G�<�U�I;�V�@�^�R���-XrV%�|
㡆�cT"P�c<��d�4j�H8B-%?�vA��^�#���6�|����@�|��#Ќ*��s2��9g�� F�ćh}�����-'S�r�����̋>l���l.Ĵ�����~/Ƚ���T>�`!��&��h{���<�!�S�Z�xdЊ�2o 2�C�8���w�O& �X(b��10�"<9bַF�dtɇ%	E���Y����v����")G4�yb�˿��(j�'�mrE��-)�~�@Q�!|h��/�L��)I�/{ݠ�h��"TA�,�aڻ�Q��I�;]��j����-�i����WBڿ(,�09�͚�Vth��ޞ<�����ʾ>ѵ�K_�v�('�G$v���~r�+�}
����sR|�0Q���ۣ�:��3#�*S�q�#*�|B�͘P!>%�w#�	��d�Y�[�Pqj@q-O��}��f��X�s��b�lE����0%Ak��wH�ʧ}D�؈6˕#~�J��'���`���vc��h�EJ�F���,6�Hh5��f$Dˊ�$[�Q}d�v [�o�<(b�
94Y;�!�}���ɣb�x���K��s����c�N�B���'����̍fś�A�+�B	�r̃,u�N0��I�?�hO�a��ր��$C�S�`u���O��J��3㐡J6�6"؈� f��T� )87�|b��t��O��Є_83�Y� �2��v�Ҹ7��#.���%S:.�,��u���ٸ���ˀ7=X���a&/��+S%�;*"�B�	4j(�c&Ӽ|0p���CGNA�҉Bf�qO�S�9y`�Ju�.B:��-��<�  h�J�	ˢw4l���ɂ7�l��V!ܣYO��`C��=<�m���ֆ����v$�����Ɇ	�ll�4�_����F|BD�P���"?bm��M��hO��G.D$Ad�����ϯ[�tч�O"T�@+U�:I���Unލa�<��#R�O4R䫗�'�.!�t��&0�
4���҈nl�a�
Wl '�P�_�,���.�=&y. �=�O��$�+۝aih�����8Rz�<��	�,���G�ti�$S�(��G,L4awǯ
�J6m�R�S�ԫ.lX�j�����ڛy�h���ˁU���0f�	#o�V�?�O��e�ʻ9=ܨz� �68�Zp2�(c�DLS�>O2m�g��a���0A�%kܩx��I8Q���!qBE,V�M`��SJ��O�Lb���O��_?R�T��cݟ*Q��'�����W�eDKo�6��N�ԉ@V������y���uR|�K��s� 5ۡi��j�}R#�G @=�Y;�@�]VI���!ғu�.�c��>�>����fD�� C)"8�i��撟u)h�dV�x�0� ��O��hcO@�tP���d�WV�M���E���&��d�h��ve�|<6MP�AJ�I��ď3gj�x�j��y���'��9q�n��',6����Ш��)�IY�� h@GBG�d�9��@GP�$H���<1�琬X(Bh�R/�!I`X6-I�'N�<�M~�4ˇ�CO45(��8qk�􊖣L�	3|I$�􈒫\�|:�LC�B�����8}�B"W�I�u���!�44K̋�M�� 0qO�6�M�6��b��Y7��O����J�TD�g�3-�80Ƭ�"��	PEU48��0�6��##L,����`�'��Xs�*ψ��Rq*��s�LU��K�s����@H/�27�I?1C"ުO����"�����'�ܸ����2�j��D��'H�Lǝ{�������X��Eq�
��j��4oP��~�$�+���*P�_�9z�$��O���1$E<j\��)ͭ:�\�C�D�ذ<� �C���OF�i�O� M���.�:~���C�cT�6y�'Z��A�;���ঁ kҭ�K� ���ָ���1@Nh|Ȃ��<!�n� %�8��%�`H���I?�O\�9���+p:y�%e��5���Ņ�H������xY�qX����B��
���#�N�@��+X ,U8��@��b��������Ob��O�}�;딌` �Kc�ʱ
�LR9aЄ������(�L�*r@�[W���$6�A�C�6I��?a�Q?Y�I(1k�1z��6��4j�<���ȋ�H� �
�6k|�E~����lD�`E�_�X)��?�	#�+P e���K;��k4`�~?� Xl�\ڕgO�A���?)� �T���9��T;�u}¬oP�ɓ��ʑP����� �����	�i���0��Scǈ{ޚ-��6�,���ɦn��!� "�:a����J�D�6m�bAM��P�/O���䇞k|٘w,�McP
�;���K*yZv�1��LaDF�4L�1�We:V�pM@��(�(O�DN	�t̚0�SmtpLDQ�H(�.�3K��lS��������)lO6ٲwj��}�4�T�M�Fr�D	�n�c�4�4+V��j$O_� mF�2�BP��H�fmL���O(�����<�j`��ڍQA�͛0R������*�F�3g�(J*p���(?�}�P��ĉ�ҭ��Rc+��cŽa���>)�h��!��B�N@�	|	���J�6�r��<L��杇 r�c�LK>&8�� <ZB���DX<O���Kq��W�q8��� �(!�E_�'�R�Cb��'1�N��0��	
H�d��'RƵ�E��YEz��.�~-ȏ���B�&Y�� �U0q��cQic�f�E�
H�J'�(73t����ݭ�?Y��č4�ވp7K�*���Xg�Uh�'�l�7o�-#�����n�1íOn�a�G@l�tr7�	�L����3�iM C@�9���s��
J|��XH�E�'�8�;$犚Ŭz�;|Q����kT�*O�D��~�YㅠC(KY��r�'��om�trՅ:�O�Xၨ�Fx�ㆄ	�:e'���b����<Ӡ4���d$�I�D`�	{1��'��t�B�?^�]O�1��+�'�m:� �1$D� R�ʞ=t{�1�px��'Ȉi���;h��a�逸��O̚wJ�;66Ԛ�Ļ;d �	��'�|M���7��A"扠sN���hJ%� ���R6,�ؑ2(�;�E��ɖc~��!,�Te_�~�OX��ۜ��.l����W��T.1`:�.S�4��2��+�yr˞�{�P���eԷ/#4��(֚X���'�F%j�K@�q9�v�4e(���f=�YdQ`�hL��	����`�f� ���t#����X al�+kP��(p�=}ܰ��c�*�yR�Њbi, �(݇gxH	֌�!�y�L*W,��k��s�x�A5�Q��yR��|�B�xs
8d�D3�DB0�y����'�Fi3�,�Y�<��$��y�*� ���w@�I#ށ�"�0�y�O�qĽCnO-OY�T�@ǘ�yB`��0Er�ĄK�
�����yB �pN��˦m�-����c�i�<I�M�-���@O��Y%��˖J�]�<�#�tP��f�98����&)PN�<9�b��ງ�A�}��5z�AN�<9S�݄1Rh�!a�.\����+CM�<I���C��,�֡ԾG�*x�q�b�<�f�ʀ.�H���;$���q��^�<�Q)�b���X�h�/g��{Ԣ�q�<y�-L�n�6�E�X-�M�U��m�<q�H&@N��M̪	�( ��J�@�<	��:Jp��`�A��T�TYhE�X{�<�2��xa�]3�"K�x�>)�'�z�<� B�
�����Ҥ���x�y�"O\�{�nԟ5��M�'�% �
p��"O쀂���b��"��7M�P��g"OhaZ1�LT�i�}�A�"O1�+H5c2��p֧��00C"O���%�4h��L��ހ'�0�0"O�<Z�� �K���n�� ΄�	�"OƩ��B��,�����#�(U"OX�AQc�`��(�gb��<�<�k�"O�|�⁞�3R%A@�ʜg�.Ew"O�\p� �9��ăW��>:c�H�t"Or�C��E�:Ϭ��6�T1q`�SC"O�����_�:HAЁ
�k�L��"O�A�G�[
�3��;I�ܬA�"Of=���,m=����ޘ�E"O�* _,I��`��#�.U�&"O�}��'^1%l����B�
*��9k�"O��bƚ~�Vݓ$L���f��"O�i��B۰Y�8�:&ꉪa֐��"OH��Y��P���ϠQ����"O�(S��\}�Շ��.�J�8�"O�x�T��D����H}�|Lb6"O�p�sB�O�ҩ����5[�u��"Ot]ybL�X�l����%~�TyB�"O��
��Rh�S�W�z�W"O�sƂǅRA�aJ����[1"O�����Ò`&p����0
�Lp�"OX�BP����5�J,	��g"OxToՑw�j�{7
�S׀�"OV�gH�-@����%�Qc"Ot�R��� ���9�$���xD"O�(���@��,p����<�6i�"O�l�$$D.h+�AAT���?�baY"O��Iq�E�thNi:���-i��B"O4����b$���K'����Q"Ol�qD^8/dz�1u�	.L1��"O�t1�3~1�p�ff��a�����"Or��foN�@5�JׄV �
E"O���]�!;2�A�L�}�2��`"O*�r��_{踛��	�ڰ"O�dC!�7~��7�d��FX;�y�O��?�h��+G 9����C=�y�÷TJ�傣�.JJ�k�!�y"Ã�_H@q��%��PG僈���G���O��AZec�!��R���oi����'8e��O�v~^��E��1%��x�'�2�10 	������ݚZ�\}�' �<�EHN��(z6�S���	�'Zl��P�w�4x 6FH?Nǆi`�'�~��2���)�������F1����'{ў�}��j�80�`3�F-}8�RƦ�^�<��/�O�:�zŃ�1&�=Ȁ&T��#�f�xp���p�B� ���+D��[s�
�}1ƅj #$��%WJ'D�����c~u�d�3!z��X�G'D�L)f
��lHAq 6���"��L�<�j�,3��i�jɼ\'��z�+t�	N8��� lB(�h�v� �>�� 8ӫ7D�4���ӎro�Q�7� �p߬!в&2D�`�'*�l�dsCޱ[���B;D�,���E$(��*ݣ��x� 9D�@k�!E�`�!�ț)=��)�F4D�́��@z9c&��g�ŪC�4D����O[~.!xQ�����M�%F=D�� �X!%Qe��9w�V|�"O<���'��-2��#Վ�!)j��'��	G8��1q��s%t���_�a4B�ɨJf�x���J]\�0���YR�C�I$�ݛ�
��]�f�{�eF b�C�I'n���.�FhT��B�9�C�IV��i�f�L���v�	�"V�����<E����Q�� ����0dB<�@U>�y��)z�Ќ�(Z�a( L 7G:�y��H�M/��t�A�&$}[e.����$6�S�O�V���.�5_0�s ��?���	�'�Jx�1i�/�M�&�;; �
�'�t�(t͌�1�P;&"Y":Rv��	�'O�)2Gʎ�C7n���-I9vh}q	�'�* *���>�Fy+�(����j�'x|����V�
q�	Oh%X�'l\�(!��Vs��A �D��`���'B�-C��^7�88���?{�"qa�'�l���( �Lv�C`eL�u��I��'U��{Ç�a�x��U�n"��z��y�d��2�� qƏ�E���ņW�y㔉e��q!�ˡCa��)O���yr�-��q �.��Ȫ�U��yr���^��HKe�#D�LH�ʊ��yR��tF�KE�N�&��5�pB�>�y2�@�(<��2`�1Nʐy���\7�yBl\�'��k1� L���(���y����#���b#��<�H�3���y�DY�?�fM'��1���E���yKĤ{H I�B� 1��](����y+��i�&�Նo�{��y�cB�M��1�Qi���6�c�f��yR��;ή͓��W�y�^��S����y���e 0HA<���G��yB*Ϻ)&�H!R�>}�F�A�\�y�m�p�4<��A��bB�ը�IP��~�)�'�M�$��6[^ �"تJ��(��F�<����|����LQx� ��kR�<AG$��J���[��� ���An�Q�<��� �d9�`�\��B�f�<�Ię�j�R��+.��`#ɞd�<��F�
o� AA�ė=S�����#=T��A�آ��|y'��BDh�PG$7D���p���m��숅��^�4�{��9D�dy��Â/�||���܏s�(,1�D:D���FC�7P!��U��/ @��+�O��I�p���U!I�8XvH��9dl#<����?)W��6H2.ő1�D h�b,3c�5��h��'\Q>h����� p�GM�W|Z�O2D�tZ$��i�m!�O����U�2/D��Q��ˡW| �H�>!�)��
,D�(J���04#�	��E�Zu��#d�*D�\p1�3�T͡#VFN�S��&D��aT��.os���C�.AM��r��#���<D�N�Y����6Ǆ	�(���:T�����rcJ�R2�y�p��C!D��)�j�"x��3�L��/�^�ʵk4D�x���	5��]ۄ�Q� 1�xZb\�І�	<)H�d���R���i�K�8�x�'Bў�?9�»�,��vg�E����7D��5FӞ>�L	q��)�m�a�(D�����7|˲�XE 8=I��q�`'D��a�Q�?�,�7b,����t�(D�@�gW�_5�`��پ�f��2�$D�� ���g��5q@,�B�%~�>���"O�P����J��Z%��<{����'*��{1�Й~^�cR�Ƿv�0\I�'�Z5b���d��p:�O�q�����'�`���<R8��#�&z�"���'���@7�(�0�2#N����c	�'$X�s�*� 1<�Uٞd/"9R���$#A�y�wa62����Y�O�!�$�4G�\GN��O�����*E�!򤙻���ga#4��ƤJ�*�!��ے!fҐ�����s�Zt+�A��T�!�dK��x�lm<���?$d!��@5"t��q�[0|�XpV���w�!�D����#J�6n("�9 E��!�䖕Is�Y�JM�/�����X�N!�$�Tj��'�B tqLӿ*�!��R�X�^|SkU����TbW63VRB�ɽ*��lJ��݀ui�� �9g��C�	�pR�}�V錾9v�"�뀲=�C�əL0�@"5��=K�H�� �zB�IV��k5��.vĺ�����7�dB䉵so\�xWc?��XWK�Y%&B�I8$�+���!F��g���M�B�I��ha����j+dbT�|x�C�	�Z �/P$�@��" S�B� C�I5n1y5�D!
[�9�Ύ6Q�B�ɣi������ �(��
�I#"O����a�ĥ�b0;�v�Ҵ��!�d�(`��I���L�/���4��(0�!�DZ;M&� �-گ�R]�iH�!�$�.rf�p�M�����
2��qK!��Bn�U2$a�2we�k����.Ob��Z��0�c�mړQ�|��Ń�K�!��#�����K<=�ʥ��jׅ�!�� 	�v�g������L��!�Dݣp-V���*ч �:���7�!�$�%��Q�e�9<�Bi��+��[��{b�\3k��p$nӗ,q�ݑ�ˁ��!�dE=&�p4�É�^^� rEL�?�!���XA��gT=Rz��sꝂ �!��� x�R��P��_I��H�)A#~�!��
&)�X[�
�CI�R�D=�!�d�1,X����FL�e:k p�!�(�}J$�R��e�A/!q!��'?�!rňޫ`����� 4T!�֌��%��e�\J��%��cB!�D�Qޤ�zR
ڪ-�9�F�5nL!�D�]u�y�/T* E&JQe�
@5!�dS�L�N@�'��-s� �E�(!� '���U�F�������!���k.��Г�X7;B���2>�!�D�'�^�(o؛���p$I 
�!�Ė�_mFԁǤ��BQ���2!�!�Ts.�9�pd�@	a!�D��y7���s�U�.p%:�(H��!�$J<o�z]뵁ĘaO��:����!��4�H��#�Jj/ ��7L�OB!�D�u��9�!e��U䐻3+

�!�D�(
xpSg��,��u�g��\z!�d��^j4����n��8��� �J!�$�]r�I�- j�޹�Ԥ}-!򄆸$��hH'�2�d�m9!��(1�h�Rɕn��$�^8.!�d^�L���h�t�Q7k��:{!�� �x�  6� 9K�AX&���yb"OH�k��ɰq� �s�e�{���0'"O��a��J~hqY�#�=rnv��"OF�Ô+���l �A�VW�k�"O$��,�)2c��؃�7���F"OڨW$�8rD��.@�s�"O�xHg]i��#m8�p��"O���%�P�8ԌyZpL�k�2�C"O:%0��/j�s��!�.�a`"O��+��ʺ����Ee�{��PZb"Op����JuH��W�R.f�X�!e"Oܥ(چ22L�p�G�D|VUA�"O�(��ʀ�D��L��'�Jwڵ�"O�Y��ء?�2���X8'�z�@"O�\�2l�L~�1����@rPI#"O6 0�#�a4��3�ܳq�D"O����xa�ɚ3� 'W+��yb�Ӹ�~x�����P��O]�yR�B){许0!�ڭ� q ؛�y�n�sm��$�\>��4L���yR��0k�6h�4jM�����s��!�y2a�����W�Thp�c*���y��",$�����}�,�hv�Z��y§_"�ԑ�SO)жpsu�J
�y��%AVEf:����4OJ��y2gr�9pK�1�����V4�yB/�49�DY �#��B�f���
�'}<ɣqn�
4���Y�� 5��
�'��-��G�938�s��F�0� 8�
�'.��R��Ԯ5!�t�&�_�(�.Hr
�'��d�����A�."��J�'�*س�F������蒤'q�@p	�'x4�+姅�lh :P�T��+	�'2�����۔ 6��K��_��\mY�'ɢ��A<X���B0E�K̽��'��H��+LL=I�� �� ���'lD-i֊K&������^lq��'�� 0��܁k���Q�슄�(���'��T3�!Y[��)96� �����',����#ȩq�ZX��� >�i@�'�VP���ݴ"L���"αA]�V4D��Kp�X<%�8̙�㊾B��!d�2D��k�֡u�ތYd$�=�ր94i+D�4�s���y�������a�*D�8�����ܡQ�%Z�|���c�&D��� 6;qt��%ę�4gf\k�# D��*'Ͷm&E���֌z��L���!D���֯�$Q~��Ye�+�f�2��?D��i�S�[���J!�"[H� 7)>D��f�ƳF��,�a$�?]�2pz";D�89���r:q{��Y�S���ze�:D��a��-�&��TR���Q@�$D�x��i��@�I�J�Rݔ$c�?D�\��fF�wE���G
(�PA�(D��C�@�d|ť�9f�,
[^!�\� 	 ����M�`��,tze�"O�8QC�K1.<��a�@��dI2�"Ob�&
H.��)j��,?�$p�"O�ິ��PK��P�)�9����R"O�9	F�1nm�$P��YD�"O���&�3f屗*�j���J�"O�ɘ�A��D�XIX4�	�Y���	3"OVݺ`��	� �֨�A��	��"O��O���9����vT��"O� �ܻ�`F�#)�1!�D�s���a"O�t ���Fr�pč,L/�� �"O����6h�ã�^�+���g"O4i�7�� ;Jp���� t�����"O>�Z�	7@U>������B"O���`HU>k ZCk��t%��"O^HQK�8�f�#��5O*ಥ"O�� RK,@D���B��-�ĸ�"O��"���%����a�%I�q��"O|�1�횭|�>��3�ߛ"��
�"O���O<�t!�s+��3�r%!�"O��� ,~��e��;</�H�"Ox���"�:=��I%�,i��"OԨ:Ġˁ��q���60�hz1"OKG�j%:@�AM�9/�����y2#ɩ9�Az�
��]�Q���Ѹ�y�
�0˦M�g�&(Nڴx ,�yr.F+����E�77.А��A�y"�4G���u�^�)��i�F6�y�'Ѩ+�D	���"�`-
WF��y�#��q:���"�� FP�5�;�yb������F��-�B,2���'�y��;��a)(�t���O6�y¡�<l��ad^�C��#���y�En����j^5��0a�6�yrlȃ U$����
�&TsB���y"��<�z�
���#;jj�[��y2A89�i���ش��I�E郡�y��W��a�V
:u\�iI��y ڋJb��-����Pz� X�yrD	~Ō0���y�D�`��P�y�H�,k�=�a
8��L�F��y�B�t�H���A�C�,å��y"gN�7�\�⡆F7}��-���ߧ�yrDoR\袳�D�oM��eD��y"I=Y-fl�a�3��]�dFTy�<Q��2)q�*j�+�#�Nc!�ĕ�#)4 ���Q��m��dB 1L!�DG
n	��Y�@�P��7�!�D�
7��-7T�I
d�_3!��߹��dZ�h�-~0p1Ei��&8!�d:������܋Ğ�X�蔷H�!�Q<@���+˖#�$a�W�N0n!�$��1������j�Y@�8Y!�$):�2�;vԹP�pBg�8[�!�R�8d"�R!�Ӌ�U��N3�!�,x��M�`��O�`���l�h[!�D����A�W��������!��>b*�P���1]�p0�CL��0�!��,o��q�ƿ��8	C�݅x!��	X��0�ʞh�T�2��(_!�U?_ڠ)���ukV�s��y�!��޾s� 4�S@�E��ܠr���!�_�C�xa�J�]MT��a��=�!�L�mA������F̙Rr�P�m�!�D�n�xQ�e&ƃ�z�z�B��!�d��s\D)3� ��0�t�)Gb�<l�!���=u|as�U���	�B�]�!��3�
��V�3��)�� ���!�DL���亃���0��|�PAΌU�!�$ɐG��!qb��7�`1!4j�<�!���WV��b$�X�dh�D�@�)!�# ��]!���Mm�X3\A!�D�+5����)�^�(P(�n�k�!�� l���J��
��9�ե��o�f(Ku"O���ra��~A�ɷ�⵪�"O���uh��������
8��G"O|�� �ѫ)��Pt�S�p��t"O��aa�3C���Lth4�g"O��!!��0n3L&aO*,�޵��"O���ghU�u�^�`�9xv�]z�"O��K��Q$n���ea�`�"O`���5	�^-��ό����e"O��FJ�9�p�,4�L�#oQ1�!�D�#���։��!�����v!�ʧ.k~��B�؆@�C�E�Pj!��ހ4�
�(��C��F�'b_)&f!�D�0;e�yJ��L�Y�bYz�`�nT!�Ĉ�s~P���0M�@x!�ԩH�!򄘘0.��c��T���X!��Xn-�!zФ1t�u l[=Wx!�ʙ@C���B��<'T�ã+SW^!��o��ͺ3�T��1V�I t�!���aS.�ڥ�?�6I���8u�!��eJr�+�a�9��S
M�!򤍊w���K�FM0=�Rq��εw�!�іP��4b��ܭ#�����!��$�j�IF�N�[�Q�AAZ�G�!��U5K"I�FɾZJ�`&��N�!��	V A�ƣ�s\h�פU��!�ă%Z;������f���EN�U�!�S�l-�℃�c�P�"�ʋ�r�!�$�5��|��O�6K{6HZ��b!�DQ�4X�]ȗ��}L���.E<`�!�d
(+́�ˉO�:�*��.�!�d_�&���)�D[�3�L	U�q�!�	n����3/],3fʀ�sG�r�!��\���6�A�@e�e�&;�!�$�#c��Y��˒����p���!�D����	@M��)�4��>%�!���7���׍��u���9�%[W�!�dÛ\��L BU�`���[R!�� 1�2Ed) nl"�I�5!��Ha�$�Ԅ�Xx��H�N(!�Q�Z���U&�-\�����#@!��z������3�b��&G�|�!�ĕh-J��D�B*i�nܨ��V��!�Ĉ�q~\�p׆�:KuHy[�!�!��1{RB�M]�fe��+���	r�!�CB�F���,`�Չ�!Q"A!�6O�>훢(ؕ2u�UZ�&�=K=!�Ğ?&@:ѓa'R=q���욃<!�ď	m2�〯}�"� wk��}�!򄆷I�:T�.қ~��ѲSk=I�!�}�
RWᖆ0�RD�F[�>x!�D��@�ƴ�r_�4x�
�!�DH�F�J�5�QK�8Zw�	�<!�X���ñk�,	�th��l!�S�}���2��;!~��fE	{!�䕐xXm�sm��=�4�B�IƲ-!�DA(/���H7���Q�):��!�$=�4]��ԟ,�����_�!�H�K�0[%�R9cs5�'ۖ}�!�Ĕ;pHuPCA�n�0P`��H�!���%628�3��p@L�����!�$�r�𠛃�ܰM��)րG/`�!��X%����u$W�V�]���'&�!��"���B�2�� ���!�� �Փ���'g�I�rfF�{9�j&"OU�5`_�b:�s�e"4�
)6"O��D.��.#ؼ;`cȹN��%"O�-!@AF�#�� �cBͽ��ѐ�"O pZ��İ��-�A�.��q�!"O\���Κ5#�2�)���G�,�ӣ"Oޑ	ś�7@��1AבC���y4"On��J*Z��\�p�8�>�	�"OƭQE��V@"$o�4����"O�q
2O�Z�V"S.�d���"O�Pi��3X��M\6Qu�Ċ�"O"ѫ�i�!`!�)�mW�wk�$	�"O����hZ=w)�c��R��A"O�*�7#����*��o��};�"O��a�._wH�Thْ{����D"O�Qk�� 7~��J�甆#��7:D��RDKC��ձ/H)B�]���,D�Lbvjؐ|�X���A�dH� �d,D�Bf��)~@���� B�<�:A+��-D�Ԋ��֡t4\���L�KDD(w�+D����o_�s'�QI�����D�|�<�@�Ū5㘹a�ǒ:~3LU�p�_C�<�1�H�}ҡ�r�]�=R�h���@�<�1˃�x�����l[����ˉr�<��F8�t���#;��� �ar�<�K�>�$E� fȟ4�(���lu�<�rG@���ꄫ� O��9��M�s�<Q��%`{&H��9.�| ���V�<A����`X  	�}l��2Dd�O�<����r���N�ok���%KO�<Eș�B�hYpP͡C��\zыQ�<9���Vd`Q�6F�WTB�@�gTR�<�4/_&	&n��3��i̱Ar��r�<׉�5%���+��DT��N�k�<�*��k5ā���F%^�ܑ!U[d�<q��܁*�n��aE_�{E
]�<4��8D��9;ٚU.\d����[�<�$��>���@��2KWd��b!�m�<�q�@6JȘ���2�>�(�Ηh�<YTK}cD��vgP�0�<H�n�N�<I�酋Nkh9�e�&W���'�I�<�`NF��K��ǓX���9\B�	+}ӌ�	!ػ렕�`(�<�C�ɮ>����qf�*.D��
D�n�C��)Hq�/X+p"NX�If�C�vp�B��[�)��pD��$ ?�B�	F���3"� `����`ج jB䉍����QK�Rf6�
�$`�lB�ɤ0@q�N��sx���	�&B�I"9Hؚ�jF�Cp�e�҉�B�)ڜj1�T
b��q��+H(B�u��,��i]+j���Emٯ".C�I)����%"A��"��-�:B�	��F�h��ϥ(Ό�ӣkә�8B䉡O��P�
7�H�" �2HB�	�!���p��:TQ�#��a(fC䉢R#L�@@��g� �r�,iC�	�B `��(�P�4�#B 5Y�(C�	�;P��c�HXJAǣR 5I�B�	'~�����l�DuB�L5a��B�I$�tr��Mq�>uy�!f��B�>(�R`; ��`�z`SUi9�xB�Ɋ nQ �Z�N �1�s����B�44�J�J"�хE�R� �J�.]�B�)� 4{��+����gH�kb��T"O�4'D�p���̡y$"O:dKP�� %��Hh�ċ>qj`P�""O~|:���,zd�(2D]MQ���b"O֠��U5�,{a�3�*�"O8t03���Zx�Ā����
2(��P"O"%���0�XM���ϒ_ �:�"Oj)R���>��c�d����F"OR��@�4,�XLW��!M֬��"O�B��,4͂}1�'�"���c"O��  Q�4��������"O$ 9d�ػUm�X��FI�'�Th�"OX�-8p���r�:W�De"Otɒ�KG�o$"���B�7���ZE"O�Q���;Ez�CC�3R`�P"O�q��"T?\]M���Jl��ۀ"O@X#Df�5	Hq���V U5v�zq"O�ܰ���NM���.�*ȉz�"O���)�\+d�U,8.���"O���jV�=}6�Qwd��![�]C"O�0"ݲ>�4d8���	>8�R"O�Ipf�̇]�������g%&R�"O��[4'�n��U:��R#\je�U"O�y�t�з:�����E��zaȁ"O�	��eУ%�٫`j۸7��ɩ�"O����@oFYf� \�Y�w"O���/�*EJJ�:�ۈ4��!"O�-��2P��Q[W,�s�����"O�)ӑ�B9Ϙ�s�~�U��6D��j*r�Vq�Ci4<0`�J0D��)�ƫS(����#{�����M2D�� ��T�P+@����Rf�1D���v�X�@Ȇ��S��c/�yR*O�Sj@�[N&�"uD�2��h��"O�t����#W\1��HQiH��"OBu�jҨ-O�ɺB�ڼgm\ y"OP��qh4������6d\�3g"Ov����3M޼QG&��svAJt"O�
��ۉ �蜣09>�l�1"O�X J�s��C!CФ9��i� "O�و�C��D����Ym�D�3"O�x#�N��*���Q83 q�""OZ�9�)M1Q�����E" H���"OF!S�����x4n�*	��;�"O��� V�D����g�e�l�a"Oj�a��T����LӋk�Р#"O�83*z�,���ˮz�\�Q"Od�S���G���Q�f�?^�j�26"O����KP����Dѿ'نy�"O6p`��2~�L�#��}r`APt"Ox�(
�!oL ��vd�5j���"OX,��m�\Z��ԣX��r�"OZY��@A%`(������ij�E "OT[S+P�?�����0��Mc�"O�e2�R1~�M�7�� ݼ3�"O<�:2T9d��H g5x�n�[�"O����N؜5� �%�<7����"O���L�?|�ҧ��|�ژ�7"O~���fj��0�߻�yx"O
(�f�˴R�>H{���>�DЂb"O�3R
�ne2HHC�ΘU��M��"O��#����|��Jˮ`Q��2�"Ot��퇉LZ��"%q A��"O��Ţ߆2XDU��' �X���p�"O� �]ce��q�DL�p��rq"Ov���)-������+��yy&"O��2�U�j���ǅ�b�0��"Od��-�f�ڒW�Ԕx�"O�@$	0d�\h���(��"O 9C��8
�Ճ�	Ӊ]�,t�"ObX�b��Z.�����n}��B�"O��GiL�E�%H@&Ey�$PB"O��"cmA<S��E�pE<����"O<h��/��l��Ʃ&��Q�"ORU�L_,{�|�KbI�s��:�"O�� ��];�p���[�4@&"Of�ѳ��g��˒�F�M�|`��*O�,��������w�H�p�J���'�``5ϓ*9F�ݘV�+i|t�y�'  X��Y>r����"_v00a�'B�����6��%Z��X;TdZ�'Q���کo8�Y
q�42�q�'���D�1$CJ]a@���Jy�'�h�qs$�	h�a�6���g�<�	�'�FM����Yt0h���3\J�u"	�'��ȁd ��d�୨§F1\��i	�'8���K�'aD���r�T4?f8	�'��
%�K11��� }K�1��'��ܘu��[�^�8��Ò,���i�'�
�*�����B��R�x	�'����t�/2`���'I����	�'�Rl&EF�abPu�H�*Dr�
�'b*��υx�8!�E�;�(�'�����0{�� k��,:�2�)�'D����]
$�
Mj!�&/�؀s	�'��.�f(x���#�/-�2���'o���^&Bzm� ��%\6>=�
�'�h�@2
6�2�'P�xqY�'�}z�!$bM���Y���
�'��e[�mͺ~!��ʥ�I4X����
�'H&��	��G�T����c����'��t3��2�kB�Tl�9
�' 
�U&G�����b�Q�Z�C�'d@(3��A�G���C^$:�	X�'���B��%g��J�--�<��'Ԕ͛恃�jo�Ѩ��V)��D��'�~2��Ɋo����c��5!t�x�	�'�p�8,��(j`�>LЄP�'u�1*dB��^����'�8Hm�h8�'bH�!�P@LK�.�6{��k�'�>���L0(�����O�0���c�'	~�(��b���a+�;�����'6��"-� +�u��.�l��'��D��g��̐��H�S-���'ؚ�0"ݪ%�.m�T%��#�	�'�t�뛸b�`l�J*Gnf��'���S5B\L(�CL�>��x�'T�=�N�"vx� �(����H�'A�US���'�8}6!]�iJ��	�'	P���.-@:NݹDҰ����'a��xE�v�$tb�/֍d�8UB�'HF!�r��=3F�+%&٫\S���'N�!��E�?���"��K
@hl��'|ĸ �N6Ds��J�G����'���WI��I.�H@��
�{� ��'��( ��L�KZL�:�g�l~�|��'��X��� 5ی�T��e�}c�'�������Eqe�cF"d����� �  �K�>i��Y�f�Uh��"O���@.�;�`�sv#Ym�h��%"OP�@$͂<�<8��b��
�4y��"O�T!R��>'�X� U��7�T���"O��p��c�0��;��͂f"O�]q%���Yz�"�:4�&�z�"OD�#�
V)�0(� ߠI��\�"O�ȣ"��M�Ո� �"ʊ,ӓ"O�m�iֈo��	�fO7����w"Ob��A�"]��_�k��)ʠ"O���!��#.s�H�mL!9��<��"O�Px� O=�t����O�v���"OJ���(�`@ڍ�AF�4����C"OP4�Ql�H����ge	&.y��"O����g��0-R�c@�q��a�d"O�X)F�5a�2 ����I�`IA�"Od�P�VK*�j��+{$����"O(` ҆=�@p	���%U�!��"O60s ��$4 ��K��j0"O~�y��|�DaC�,uMi�"O(Xj��	Z#8��ω p��"p"O���v A�),���6����"O,�Y��Ҫ����&i4 �S"O���A�]�J����C�Y5��a�"O| ���V3<��I�C$2�-)�"O�գWFJ<H�0Qw��rb|�R"On}+���G����G�Dd�`a�"OD	���A��\C����gQ��"O�%�P.�: e�'+��"�YC�"O8��ƨ�	�&|s�O ꬱ��"O晊��+9=^Ȓ�/�{q�XE"O��z	�{~�R�OҌN2Z8""O��J����_�*������"O�\��R:����H3*�B��U"O�2��7U~ k�����J�"Oi@��
�2�@�;U@�b�:A�w"O���"aD+���2�n!a�|�#"O������)]\��-9{ߨ,�"Opr�L-uL�����3)ъ��B"O&���WVy�x��У5��A�"O-�
�J,�L��w�f���)D��B6Kݤ;Ͷ��󉙭3:&p���)D�\Hu���c2��6�����!�&D�!w�Q)���ݥC�$I�%$D�$�`@��S&(l��[�5�ƌ�J"D��h "_�Ʊ	AO�8>a��p%;D�VIg��Q� �Y��µ�Q0�y���'Ж@C��y�r�!뙴�y�Ő7`��R��Y��ljg���ybm�*� �����ScmLM��y�JC*5��|�����@�X,Ҡj�/�yB�;B��|����+q���"ĉ�y/
�Rt�0��6\z��jʥ�y"���a:��@�}�ไ#�y���LHEB�KL7&jl�BE�#�y��Y4I��� �ħqD�4M��yb��!v�<QJ��	�� ����y��N�|�*f@S:˖?�y�䎐>��:ȋ?�A�ƨJ��y¦Y�r��ɜ���G��yBD ��D���v.���t��9�ynʅ#9Z����ja��[�E��y�ȟ&C��QC�m<L�,�`v%��yr���vb�����=�x����@��y
� �Ixbթa�8(s�N�@��}#G"O�Ċ"Ģw���0"��������"O<�q)\�\���Ə��b T"O����	Xf*���&K���"OL��! �[1!UD]6 �@�"O��a7f5�ؘ`4��T52A�d"Oj$��I�{H����&� *�L�Q"Ox5S�ɂ?en�a`���j��@5"O����L:p�
8�댽~fz)p�"O�9� �|��9F`V�u` 8#"O�� ��=o�DB�.
�!&�%��"O��5�D)%�!Z獇�!*�H�"O���_8{��u�W��_n�h��"O��$�ECj�ݒ�Kچ{iH8Y"O���`�Ƙ���'���Ws�؃"O�A�ʄ�|=�yp@��5K����"O���G�=��n<60�3T"O\9��.	-l� +��]2#���"OxD&��U�yč� 4=*O��Pp��$~ri�7�I>s�XI��'kV���(h�@9Zx,9�'X�Ȕk�~`�e�w*b�@���'�BeEŎ~� 8"7�#m|�$Q�'Ĭ���̄kVц��k�=;�'�^p�oX�NR�=�u��n��̸�'᮹�t�K��y+6�0b���z�'!Ą�t�N�%��b�@[�64�
�'���`�LI���}sr�DK����'�)sFA�Sc�(�L �>�@H�'j�MQaײ,.�HP<;N���'�|ࣰ Q�#�)�A�_�As��'W�1��|�dIؑ,�?�P�ʓ>���C_#�>h!�e���ȓV[�Av��_�jM�����k!Xфȓ5�� `���97tu"cmΤG����-�hC�"ێH��'	*-g�5�ȓ{s:Փ�J"nܴ�t����n��ȓ'�P�At$�9��<�uR�V$��ȓm@"E2��B�c���ԁʧ"�X��ȓ�6�:�� $$tڰk)D�Ņ�Ol�U�Ӑq�ĸ@[�O|0�ȓ2}4��&'":~������{x5��4�h��� zwn�� o�����.��D*]�� $����
@N+D�t�@ Q�)&�qb���֤5�$D������e��#%Ӝ1Ƞ�A�m0D���')��E�.̋M�~�q 	<D�h)���[�LX�M��P�Q�8D��*������ K
�&���4D��çʏG��X�D-v�0���0D�x��� a�hZ�D#T�)ö/D�8���E( �šХ߈$�&����+D���MHc��K�l
%Sb�� +D�������\�*��hZ��@)D�����E�u��*E�B�r�� �`''D�X�+B ((9M2$�	�1�&D���S��4y�T�`��K�8�.Ђ�!#D��Cm��;r����H˴{
���! D�XRA�Ǟ�d�y��?GJ@�$�#D�dY�!D,:��qWi�b�,i��  D��cEn����6�St=)��<D��ɣ�D�f���ӨG�_K�=���<D�pR�C��tj:+X��듍 D�0��[�C$Vx��鐋P�n�Z�L=D�� t�rd .�<I"U=���2"O��b���1�^�+%�Z6���B"O�c�̑�W�BP��F�c�&-��"O
PJB?Sv�%
�%3i��8�`"O&̸��הE�0 ��$t��Q�"OΉ�7�I� ;����?�p�r"Op��@��Ne5Y���v�L)�p"O�!
cl��r��%`'�G64�Vq	�"O���P���J��ڑ/	�)���!B"Ob��`C=[�^e����>�p�J"Oؐr��	�L��{�J�*z��
�"O:�C�x� 1��,�)���U"O�1�'�.[9h��$�@��	�p"ON�3.лx(�j�.�0,�*E@�"O�ԳB�	�5�Q��Lҋ �ʱa�"O�Y�!��u�����KԿ��0�"O��Ғ�F�)�@�dIڳS�,ma�"O�д�.~hI��ҨE���5"O�}�FT2�(	�$�&Q?�Ur "O��D�W&)���ab��*'��2 "Ozu���W��ز`�42~m �"OD�)3b�DTX�J��!�U�""O��%(�$`�ι	W
�k���"O��2a˸Z\�C�h��seL��"Oڄr�,� +��z��Dc40a�"O
�X5�ɻ6+F0��כs|�h8�"O@X���
60@�f��"Rl�Y�"O���_�h!���Ghrh�u"O�������@��
�1N��r"O��CM��{Md��wI�s�f�S�"Or}�@E%>�t�էP�Υ��"O�<PT��W��}�a]�>���"O�<�D��R��p9p�����urS"O\a@��H�;t$Q�G�Z´��"Ob��b)H	o[��sѥ	�^�+0"OP4�Q�֣-@E#p�%h�L �"O<�z�Z
_c|��c���-�5"OB�
ѣ�?Af�3F�B����w"OX|�U�χ!9| ѥj)+��Hh3"Of����אr~��1C�\�8��0$"O��Q����T���E���8ֆ��"O �t�R�/��t���Ky��X{0"O2����&q��2���G�4=Ht"O���B�C�2���׺T�D� �"O4���'��x�#��7j� t��"O��
F�'��x�$�#/����"O�#��N�3��\�p��Jle�"O`�C�lW�9 �P)�!�&#���w"O,�wL�E$^�ɒ���V���d"O��k���:v�N(qA�(�`\�"O0E�V�C���ᰱ��vh�E:Q"O.D���: �abGiY�R ��"OJ�{��	w8mqd��iCj�;�"O=�J�WL���`�	�'�lل"O�m�%�)/f��b
�p  1[�"O�B�Q-k!�	����m<��"O�l� �͜RQp(��؟l_2�@�"O���P�&��u�D�z����4�M|�<�׎K��b�d�G>�R�I�I|�<�YL�R,�cN�+�~��ǁ�o�<��KZb��RJ?RXN��c�m�<Q7�B�sFР�����4�_i�<᳂�"x��(d�O�;�jQ!��[�<Ƀ	�! ��P��I�51�%��R�<� zhhaB�S���bыW8i]�Aj�"O�-0V�*N.����
ɉfQhm{�"O��"fS%ZV�t�ʏ4�~Y��"O֑���LOT�A�BI��I�][�'��P�1bJ��͸��Æ?�H�'(����,zx@�'\�t"��	�'FX|)'�Q<^#���$�, 1z�'�J�SfbY2����C�(,�!S�'�z �!�E��k�E"f0�'�!@�mM<G*Z���.������'�Đ`3D,0�~MX� ة�I��'�b����WZF�Zf'��w�c�'�d�%��%X��\07cշn r�Q�'���L(Ng�HY&�cp�'*�&%�qH�pUMűb��9�'���狔q|h1k�Bn$	��'�8�K�O��l���+��V�m��uS�'�~@YŁ0H��@�k�D�S
�'�h��&m��, �ZS��o�rp�	�'[|�[so��"<*I)�`G�l��'Ql�;�/[�&����3^w�T��'Ϫ�;%R�t	�l��m�F����'F���w+�US�F�'����'k$ ���ˬj^$��𩂶 q�]Z	�']J��DGJ�0d��@�^�EY֝(�'�a3���;7�pu�Q{]R�'\��w�P+���IE��zY��
�'��"öt#��HB�3nl�	�'�X�� �c%p�a��*H�D9��'tL���@+"9V��ŌA�G�$��'g�I��9[��TK%@76��U��'�h�����Q��S%+2���p
�'Rb�FR [C��Ȅ��/,��hj�'(�[WE@�#�2�Z4�ަ �Uq
�'��hPvi�p ����D�}�p�	�'ݸeHWBy�����D�A*�u��'�i�c"&�.�W�D�2@��'�y�w�]"��=�ցȩ?~&4C�'J<AS�ng9�&$��';n��'OpmY�IW�
�d�d�W����	�'��{��ǱW����� �����'�<�21��;���Z���L$��'V��ڀꙞ���ŭ,h�)�'�PA�0�W=f2���u�S�{U�LJ�'�L��rM�_���`��D�l9���'{>y��偱GT�Ѥ�̇8�����' �MZ$,�vD�S4��y0���'nBM�AgA�9�t��guD�H��'Zx\��ɛ8ۦpR��k��	Y
�'����p�ШTt�lq��L'2lb8Y	�'�|�7�̀Ijƭ���B�U�,��'����A�,[�c�,�X�H;�'�zA @�.�\��� 9d���'��� 6��a�����Aگ�H�s�'������(�E�
�:�x�'�R�ȶf�'Khd{2���9|����'ÜX��dȷ=�d�Q�+@h���'Y:d���-Iɂ!jEl�[���'�&8�K��Q@�st!I'���'R�]�aD64 ��� �
�k�X���'�Τ*�J��Pp���
�)p��s�'2��"�P/*;B�񁩒�b�:Ճ
�'/�a���3@��Jd�őT����
�'����AE�4�鑐MjLU�	��� �L� �B�A'9�"��d[���"O�m m�S'����`ӊKL
���"O(Y���4"���O2E9��Q�"O�u�M�&��ȣ��%.�I�"O@5�S �s�0	����"O8<�1�ʮ*2J㵤��>�6���"O��{C� z$zؒ���J`v�j"O��87�T-;[�2�R�jn�"On����I&nl��B43^��q7"O�8�LO�;��?&O2�@�"O�����!R�0���ќ$��y	"Ot���E�oP\$`�F��C٘�I0"O��ҏڧ��IVG%q�H��"Oљ�b�'���J��
g<�[ "O.���a&8􁱨H�$�d9`&"O��XukI9���'��(��"O$Qڶ.](?�ڹ{'�P�2�H"OơA�&O(u�-�D�@�c�]�'"O��zCn]+8����/�"Y�B"O�4���O�.4���?S�\�W"Ov���ϵm�@#eڑx��	�"Ǫ��bV
��iªILŨ�"O�4"�F<��T#I��bCL��"O�H)0���}�ȑiԨ��b�G"O*����".�ɒ��;e��5�"O�Rf��9T�a�Dٗ��Y�"OB|'���iM,��B�#��A�"O�]�Ǡ�}�:�Pc� ���	��"O�,�-�N�� 2�����K�"O��
q�֊I`cN�7UX��g�<��%�J�:�	�"cAje	�c�<��Hl�j�KVo��a�B�)�$7T��$Lݧ(�ȋ�+�
S˾| �1D�8�0b�>W<��`�6pv|�G:D�H��
�,̡�&.l\�k��2D����OV�G������Qb�a+�3D��z�"FM�~Da��A�V(�Yrv,6D��Q!i�4i6�<$��"�>���i2D�0�"C}xܕ�ʛ�~�-{�#=D��R�B	f��i	��+*�hA¡7D��!t�ݦ5R���GK�)t�ZBE0D�l����N<�ЅkՐ�Pt��3D��1k\8t�;��ӖG��u�1D�l#)�:X�l��� �[C4@hR�<D�H�6�^����8�@$�b�c��0D�\w��g(�$pC�"?��rP$-D��˔���[��}��A't��js�6D�����08U�(�mݮ ��`�J)D��x��](I�d��b�[�!А��(D��"EZ�]� :��޿E��T:�+D� A���<BR�rC��&K$DA���(D�ء�n�p@#ɐc�8�2� 'D����eM�n0�ల����Pt+&D�� �N�T�L��FڑY1�1��)D�|U�����ʖ=2ܶU��K&D�(��×nv:]���O'oҰi1�(D�\C��) 뢅��#N>{��]@D9D�k2�H�pC�T�p��W� V�)D�Ҵ+J�R��ɳ�IȈ�B%�֣+D�|�cd\�6�ݘG���|5��C�<D��!1I�oQ&]�NU*��Bi:D���F� �0�HS�[q��e5D�� A*�J`F1��e�o���h�3D����ؘg(5��� �(1���%D�� BX�q��N+�`��C�%�H1�"O�ɨ� �%�̸� (��9ٱ"OR	�WW��k1��C�ݣ�"O��Hr네|Kpr�T���M�q"O0��tOO'>��9{��R�Dae��"O4��0E3�F�@VLȡYJ��"O�51W$�%�~��q�N1D��ۢ"O�
f�@������	���)�T"O���I�v}�
�=x�A�r"On�AQ�܎EqИ��ȝ5Vf���"O�����ޓ/�B�z�fQ�$y�
"Or�1�.Ⱥ*����Q�H0L�-k�"O���w �@��E�1$M�tF�T��"O>płJz{�ؑ%-Л71�0��"O*Ei��S�-ꪹYa%�%<T�U"O����S�E�x�Rb�F�sR(2"O���e�95���X�$�����$D��1�h�!2MF�H��X�Ύ! �A'D����h�/<$IB�X�MI"�ssj%D�@
A^��a���Ӌu�t�%�?D�ت�G	(<���lQoH��J2�)D�(�F		wD��0;Vd�RU�3D���k��{��$�@���P���1D��0'�5�T��Cg�=9�vt@�1D�hy��[/R*�
�k�8q�q�g4D�@2��=eg�C�[]0�1�W�'D����+M�(ڀ$�GY�:_zġ �#D���u�C�C��RQ��a�t�ҋ?D�X#�� ����!X�w#t亦	8D�P�P�ٴBU�H�Q*SD�8\tO5D�;�X�Ql�p1�̟^����1D�d��l�"��C�<���I,D��Z6�I�+��l�W�I�L��b�.D� �fK�0T�l��B�F�f�:t`r�-D��;c��i�rFl$��C�-D��[D
��c��=I�BE�'I$D"Dm+D�@XR��W::�!Oؚ��x(*D�tRR���?Jl�K�)X�q(�%�p�(D�
�d���yYJ��{*8�k'D��IŬX
d܄�+�B�/z�h�9�G D�آ���Y#�Q�5f�*@��5�<D���0�\�WD-J��ޘ5�89���(D�D�rg�8m��:E��-��1D��CkP�2�bE���ܳr;(���o*D�Īr`�� �P,�q��Hp9x��&D� �b,O�|�<�c��@�Y��!'D�d�DՂT�	�A(��tf�Qc�,$D�t�$�����z�ۦscP��H&D�hy��IH�q��Z�e�&qJP�$D��(T{T��Ƣ�
I(]�$"D�����ȦB��]�$��'���� D�ĀT'̞&�^���Nu`�}�� ,D�@���B��D�`�$s�̭��+D�Lӗ��?���;�՝pjh�׭6D�����G�6� ����1b�cԈ5D�r��>��� V��e ��3D�4��� Q0�/@�S����d(?D�tI5�o����Cߩ�n��h=D����ٛO񒄱fꛝ��2�;D�����E��cw�؟h���(5''D����	ε�R�X��>\ \����$D�Da�c��S�ܘXġ�xUzQ�g$D���꘳X�x���"�d��2v�-D�8H�*٤o^,D�`ώec�Q�6D�� �={�	5�.��熎�X�!&"Ov�QӌM:.�:l��D95��RV"O }��ĸN�m�����`"O�E���B>S��]�%� �p��"OJ�i#˄G�٣������@�"Obb#��N`�d���i�bl��"Ot9
�cC�?���P5�%%��"O�p!w�W�_�����]�)Ć�P"O���]�R�z5X72�U�""O��h�N8A�4)؇��
}.Ј1B"O�0��R��E�Rm�	���i"O�5���C$5v��ՂV��J�"O���1��4~�A� �Q]��EC�"O��{�J�z�4�5䝴K����"O~���jWP���#S ~f�K�"O���7�6C�r�;ċ�Yu��"OޤrA��i��
aBR�;Ń�"OR�KF�F	!'��:b��%7�i��"O
] �1`�ZQ2"����"O����MԐr��2���PܸC�"O�p�nY4W({��D�I�n)�"O��PFK�����~x�D"O����I�^;��Sm�#a�\(�"O���,D�d�zqX�� "Or���L��!���DP"�2���"O8�!��y(:MQ6)MR.}C7"O���6�@�)<�׉A;z�	�"O����Λ,G����/-)<A9e"O�)�`F�����'�DIt�m�"O��в�ΧRжlbV�W	a�0��"O"}Q'� ?]�d8�oƟv ��B6"O�c����ZS�nA89�(9	u"O2�p�G�H��F�5>�d�"O��b��
�	��HY�HL�]�v�0@"O�l�0K5H��	��h�,B�T�V"O*��'D
P:���i�?=�$�+�"O�s�R�T�3�聿f��a�"O�RFM����8�&W6#� %�W"O��/��>d
%��q^�'"O�Yӵ�\�k�9s��?�J=�"Or�����UTذ����^��ͪ"O 0)��E�.�4�3���L�"O̕���4a��af�2?��,�D"OB��S�^ =n� �C�"P\��"Oܔ��@$}8���7f1�I��"O�!2�'�3��<#���&L� Y��"O�`����O���X$
�{�ZP "O���EM��I�©�A�TP�"O���W�O�K'�4Y��$>ѐPq@"ON,�Bᇂ$~��A �Dc�"O��H����P�w�ވ�nI�'"OH�0,�tF�j�Æ�2��ы5"O|	���T�ah� �/� P��%b�"O!����
*�q�T�B�[����G"Oh��"�,�,�Ҳ!�H��"Op�����"xj�m�6+�@x�"O<�b�.���C�-��>�n�)"O��S�b�%��|q�LT�K/���"Om��Ξ6=&�"'�2M�t�"OT�kWb��A�R,�Ǜ	dc���"O��C񊍖6�d-@�o 4j~2͘@"Oj� ��͛-�.�Z��̪gv� s"O���4�{�( �0c�AR�Yѷ"O�x���"x�×dնg.�|C"O� ڡrS�G)�~�	u��*i�^!��"O�����k)�s�D��>�XP["Ob�Y���&�:Nt`HI�O��l�]�L��.J^��	�-�I�jB�I�|	�u��Ę_�.�So��#>�ߴR��D��F��	��j���}�ڧ��y�L�;�R��ũ�'K�����ø�ybHS�]�����1D�$"6M� ���"�O0@h�呻�&l;D'�IÆ���'��	�8�0����x��KVa��C�	�Ȏ��a��v=���"��t�C�	�2X�y�+� ExmX�E+�TB��(1�~��J�nK�x0��<!PB�	���U���\?o��\X�!+�XC�	�\�pKT�Z HF���1}
�B�ɬ>p
��hX��8i�c�1_A6�'�ў�?�&�=G'�p��ď�3VmZ.#O��0����	[j��F�1i�$ݣegԣeqO��$K�G<$M�NI�,�2��ƕ�\��M;���IP,1�:����S�D���b�%��o6!�Ư^�^,�.��A�e��D�6V!��َ"+\0�S��0J���R��z`!���>T:<Py�(D�'�6�� ��S�4F�ĥ@� ��UYGO�:k��rfEJ��y�,��ƙ��Լ0n�S6m���p<����[Z�=�r`B@`ZȒ�Jѫ0r!�@9)��T�a(�e_x@(K?s}!��P���x�թL�X�]HVl�'K!��Az�0���-9�|��Qk8��'�O����C�B�Iփ��D!��"Oh(���ܺwu�1J���Y� � "Oj�ۃJܥ��e
EDG�X"tx���gX� I��-eИM��˄�S�PJ�m2�O*�I=k�6�x�D�.��&��7Q��C�'� �0$�-���8 �(�zѓ�yr�x���`��ؗA]�k�P!�3�P�w�6�ȓ+#��@��_X�-�7�*}p����M�0�J��Xs�`~����(м5��� 6��)��f�!n>�'����	�S�(��E�B+4�s�a�4S��C�ɩ)N@)��4
��K��9���mH�����V�K:pSʬ��w>
X��e0�y�.�(9���bD��Ԑ���C��y�����dbťňF�9���yR�V\��Y1)�*!r��J�
�>�M��pGȻwu�I��G�>p8ۃG.D�l�⇰24�8[�n�vV�B�+��hO��*h�y�̏�W�����5y��B�I�x�4wLT="Ѭ��&��^$�B�ɱ�,Jgㄙd�nLKW�6v�`�yy��',� J�'� N�MX�ɎJx���'8�1�ØY56M�F�59������'$
�AWŖ �)���~���}Q����?�O��][ht�p	M�|��ıu*�Q	��,G{J~�r��n�h�P�]/2�,�k`
�x�<1�IC?z~�<b�(�`��q;� N}8���M�pڲAR�-+ ع�.��b��0��(D�´�/�
UBWb��*�Ч%�L����'	�Y�g�7.V9�f��:1�v��ȓT���'ʞ;�$���_�6�mA�����&��G��U)�f������<�yr�T�!���X�=:D�����ybb[�T2���7q�rE�C����f���Ov�z�-�-Y��)���4���S�? 1;�gQ�1H�H�CL�"[�Ͳ���"lO�18��U_���Qi	� ��mHp;Oڣ>�'1O�%�� aJ"��7��U"�9O|���ɢO3R���D�2cp☢I�c��O����|�H?i�C�V�\*�, #&{s����i,ړ�0<��*(6o�[�o��?�$�aWcV�'�ў�)׊Q#EŨ�0]��kv�� Ez��Ynڜ{��9�)�.Y��p�� &^B�	�$�b4pu!�3Y�lK���8���I?����� ��k�IX�H��d��a�|�i�ў��,�*�Ԭ~�\E��LƂ"�zt��O�=�O7�	�B~j��놠?�0H������� Oy��쓼3�n)q�Z�P�����'Q���`(ωT��y�W�T�r$(��x؞�GÁ�J\y(4��:�h��M�>���M�$����Yf�T��lU	!��S�<�V�d��s�ӝ3�,�Hi�j�<�1�D��i�
_�#GΌ�B�[�<��a���C�DE�Rk�ݣp��Z�<yd`�o�ԑ�NlE
����D�Gaў"~�	�`�J��P��W��[Ql\{�nB�$/�鴇9j���R��Y�"=��M�©���9Q�X)z��.C��%�ȓyx�x�c�v �
L5Vl�mZ��x��ʀK6`�(���ؘ��7��=يy���/
���P�	O@\QŪ��y��޵V"`�I��J�څ�ǉ^'�y�J�7wc|Y�# %A�n�"��ɐ�y⡊�<����@�I>��!�aM;�y��Ͱ �Xb�\!<���[0����yB�B�beRy���]��� ��2��O.�~ZТ��BzP����Q(5�,֧l�<���Č@�:Ua�+�#'`*���F\�<�fKй1k����kJn�jTӆ��Y�<ɶLD<�\hP"X�:�"P�m�<)�H[�+ZuJ�
�\bx�Ri�N�<�8c�D�fO2(�┺��J�<a��Nc�u@��_�Sr`U��_{�<�S�Rx�����I+ d$2B�L�<	0$�,�A�͜'	 �A���J�<��!+B��0�`���.Ȱ��C�H�<Iw [�r�,Yf�M�Tj���7��|�<q@��w��T�A��TFXap�|�<�a���2偲!�I��<i���x�<�U��!�L1�l^B$E��H
{�<��ɘ�v���@2��>P�U�D]<���U�H�c0H(U!�r��ή�|=��2^@��[,q/~��2V����	F?ٱ.<O��t���ѝdAD��B��F�<�5&�Tb��K�΅�`F�cl��<����t�O�p��28DiB �:���'i����E�Zr<<���@�8�������M��$/ʓc-^�+�N�6@�9�-��6���ȓ\������E��1��B�|L�'������{�l$��ŕ$vv�ڴ�FX�'�ўb?��D�?(F�1LGYX�ej D�4�"		[H����_)`�6�ȡ�=D�cK�  6�Ҥ���:I6��$<D��1��M0*)BLC�M��Stf��㨶<��/}b��s%��ta��w&�(N�d0�u�%4����Ԛ��预�G�=p���KT�#�*�1���D�!l����z �1C��$T��y��'b!���.iߞ�{��Q�BB���yr��`�<y����=k�#����*kN�Ex��� ���mÔL,����F[�a"O���D}��C�JM:d9>yi "O�P���*�������b�"O4X�Ā
�"�T顨��}��5"OM*�1M�A��%��fѤ( %"O��ڠ"K:?8e��"�5+��Q�"O�#C���</���ТR=�#�"O*��Y)�L895�V�w!
|cu�Yg�<�O�?�q�+���<�s��`�<�WLZ��b1�a�ض4d2���f�^�<�R������rЪ��2rRh���e�<����/N���K��}W�- ը [�<��
��թ�ᛶJ2N�qS��T�<IT�ܱR�E:vK�����P���U�<I�jK�G�8���E�����0nZ�<a��V�W8`���	�I
��W�<�VaK	h�lQ �� �X���� IQ�<iqI���@Db!(�H�9t
�t�<� ϓ�]7N}��;� �Ʌ�Yi�<i�$����%g�?rv�(	�oh�<�b��.WV�0�da�2��-[�,I{�<�q�E.$q����ɲ�8�3C��x�<�ǧCQ�t�Z�U/;�n\�Qw�<��,d(�Y�*R+)�Ȥj���G�<���ҔÈ9Y��a$ճ[JB�	2U�5���Ρ)�u�3��*VC�ɀU�n}����,�s�R�K bC�Ie�A�F,j�\U���+%�zC��:w<�����o" �ud*o@C�!(��B��^=!��C�z?hC��i2r���MkT �o��l�TC�	&/�tp3덢ay���͇j�jC�	�_,^�A&
œz�}[aJ�HC�	t�� �L�1��P�퇲Y��B�Kͼ�V@ܖu���֏�!)x�B�Ʌc��H#C��"K��h��j��	3=�PB�_�f�hU�)d�">1��] c����� ���*c��Q�<ycd�L� �����`��c��I�<�5DD�7T�����A[�P�� FJ�<�7�E�*�ؼ���F�����ǀE�<be�X��`��$ѝy�R�Q�&�C�<�(/zF��aV���N�y�<���U%�X(�Ǆ^�Z�#&��y�<��G�:��I2��(���a�q�<�E���/o���T�5l<Ȃb��p�<����}�ʬ*���g�����_`�< �F��l:B��dNF�x��Y�<�6�S(c.����R 8�|���[�<჉	�#u�q�ᒊhx����z�<�î I���Q)ʒ�\���R�<Q.�(�Ǌmݾ��w��H�<�`Õ�o�+B�C��� jEK�<�4H�'_]*�p�ŋ�?e�\C�J�<Y�d��
�JP��է��qȁ� D��k#i��n��3�(:@0 �!D�L:f�M�S��*tM\�$� ��+D�t����Xi�� '�/o��&(D�܉�.R�qI��+h�3M�)��%D�P����:(D�h�B���W�$D�tѕLT�b��$�"��k��?D�(c�-��Ӝ��N�	�bx@��<D�,�g�K�Np��A�F�8fBNX�A�8D�!��"oO
�b���e�(4��
7D����O^8o;�%2����Ȗm�!�� ��Y�)�y��IB��6Fi����"O���4���H�>!�g�u�~�xF"O!"�H��"^n��� ;�8U"O���e\�=�:����H�J:]�u"O��3D��Q�H�K ��r
��I�"O�a� ��(��$�g�f���"OTq�A@�	�t��1[�̹g"O����Cֲ%n,sQD]�sԨ�SE"O(�	 �g4>|B��b�H'"ORT�w���+�x�P�
mF��w"O�pQ� 	�qj�	��ÓY\�B�"OXd���9�ՂU�IK�M�&"ON5��	>L���蠡N���"O�ȃvi@.���#j���"O�A��O-��ӕ`�?0�!BT"O� FH�NH��O�Z4�"O��X�x���ʀ� ��Xz�JO?�yr	Ű�pbE쏮Q�F`��H�7�ybm�FmQVmAT�)�Ǯ��y�&_	A���R�MX|Uv<��
��yҩ@�ux��90H�\ � ���y��(� ��.���0Ƅ�y"b�9���"G�z��S�I5�y���)&�8��MM�h�E�0���y2l��z8����F�Q@���(�y.דtr�A��+�(�ny�I:�y�Ճa��5�BUY�BD���]��yr�i��Q��*�$�%���y��8�6�k�˪/v�aR�/�y�/߳F�����H.�zP��M���y"�ȃD��lh-S&�JE�')G �yj��N�����(^&޲ 9�K���y����}I�V%	BR8sV*O�y����,���g E�ʒQ���y��Z(�����UF��-�y��2oa��3OW���l��K��y�鍺_��QCV$0���&ϧ�y2�	�Kn����J�0�dO,�ybLӒ5�V	�2:̀{7,�!�HO�8�I��h�}@m>�<0c��Q�6ڜ� "ON��M�%��fəy\X���?�bIb�����)��<Q�'_��2AIת�o�6�`'�V�<���ْb�I(Q��nG�h�LH�9Sr�C7!bb�����yH�
`�3�ӝ�j����"�p=�T��X�4���hF!(�U0�e�S{��׌�81Y�u�"kE�R[`0�G�(pϺ�	X).���'�!��C�#��dza�<d��0�{�&�=�z  ���ur�t�ɕ2��p�g%F6s��K����y�^� ��N�xT`l��ιv������,S{T�qG�%7à�(�D;U���
5GDs��IZsl�R�B�K�[>�	�+3F���/<�@�1�*�&�Z��)a���I o[%�f�y���a�� �C��,@^�Ͳ��Ѳ��̨�i�9`r�:d_.n"
á�H^��9��f��F^���fB����ذ�ٟ���TNZ�~v,��*�o����'r ���k��<�"YN��B�mŘ.�d�%jY�RuҝJ��{����+�T�U���Qp֝*BZ.U��Ow؁R@��TFo�೵ ��м�@�#��ܜ����
QZ0T�<X��Hm���׎byrCDR��P��� �>8n�X6�Ѡ4N<I�pMT#�x�#��HO^�b� ����J��� �֭r��īC�a⑁N�unZ�K]�D�Z���zD����]�P27"��,�((�n\�?��r�n^�T���B�4��}�Ӎ0�O�P�T� �`Ȭx@���,�6�ZD��Ju�I&L� :%���+CI�L����`ɬ` ���,� �r�ɅHp�0�	b�,�����?>&��"C%<O.�ڣ�:5>���D���
A	��5���Q�Ňzh`bDŪ�pH�+	d0JL�G!��rMT�"�6���y�#�jhJw�+�M�s�bQ�@�R��� 6U��LX��!<M�v�>���q�ŉ6+SaH� �m�l��'":�JD%ϊ]T�mB�fԪ
��My2 (DS���e圧vnV���_�"	2�b鉆P7*��2o�t�<�(g�!J`tH��Ø*��8 �*SPu�c2DS2.�S�V�j����\�&40��!�A0,�l����_�4-��X�XK81�B
7jm����m����g�#���)S��pt8���]�p�Bq�^1�*ǡl��������9s��`y
� @L��D�~V��Ŭѡ Pᩒ�'���B�(
��t	t�Ҷ%�2	0�Y$?���$���q���sli�u��!.N�<pH0'M��	>]�1�z8��#L1f!�(#kA2���Q��*��#�K�q���G9q+�Ȓ���t`��S~�ڇ�7B��|��*�y"$R�x,�zw�F=,���5eT�!A*�a�-u�b��BPZUJ19B����O�� ͻ�:���ѡZ�N-��E�>�Єȓ(�~�Zō�O�f	�� Z�c��Bo��V� ��	
�1o���q*շ�(O*LP��3{���BD<D|� E�'#�a8�Kǩ[",@�G�E
vYR����G�r��AJ��?Q� %d9*��DFf���钀ВDr-fb�0+���\I5�F3SR�>MȖ�ܳ�F�i�EÜ���e<D������I��Fd@�����<D���e΍�[�H�FMܱ8���)K:D��y�j��&z��įܘ\�T�� 6D��c��Pv1�FK#O��L��"5D�HY��/QӨ8��%W5�"4��i7D��1s`"g��o�0z�<@[RB8D���4��NX �!R�T�%P�*D��0��_�SsBȑ��7D��0PF�f�I3��d�#6D���F��N�lb�iZ6
��	��;D�PX�M�m��`��D֬G��e8D����E!����r�׉{���� 6D�P�G�)�n�pd��372�y#�7D�<*�P'�j<�Q�7� �`�./D�*�� ������v�\Q�5�*�O^Y���!�M�Dj��w�j��vk�����:R�<��HѦ�1����ˮ4��L�'odHZ��STQ>�s�eF�e޵��͓&�~�h�g&D���W`фe��,���!�2u��≻}U`�KN�9�|ӧ���N�K
�3C��L�t���'�y��D�BX��3e����V��~� ]�-�,DA��	�$,�<��H��8$�c�=.R������x�b�I
+1�0�$�l��0�7�ǧ%��yZ�'c��� 11�84���%V����^Bi�(�g�[0����3׉�2&�r4
�g`2��[D"O�V�S*��P���z�ȸ{#�\�c�.�⡩�7��S��?)��/R:���FO�h�E�®{�<��	L�#6�+�F��W�P��NPv?	�I^+2�x��"�:LO��vb_����H�D��o���
@�'g�-���0���  �L5�kAX�i$5;��J�<�W��ɩ ��5:i����G�'~:�� (��N�Q>�#� � >�p����	�`>D�4ئiY�"��$�*��C��`El�O��9�kɲ𸧈��Y��/�����)0��;�<��ud=D��'��:7���Q��L��!8�d=D��
r�ɏxfYA�8p㈹:Ϩ!u����{��,��L�"U:��8$��ghZ铢�9D��(�D0񦴨G�N*Ib���@`Ӟ�(�����*����8��+Ac�lz�@2ˇ�M��z�c�e���� S�<����$)��:#B�k�Q)6o�)�ȓ:��m����Q6xl��!�$�>0��@���=}�?���*Gy6&m8��M�zfN z"D�L�aL\DI�ɞ1;��Q�Pp`�͏Y@�'��ED�,O��Zu��[��P�$�BX��"O~M�pd��3
��C�.Y挢R�W4@rX@c@\�S8a|R�"S295�7!`�p�D%��p=����:P8y1)d�i&
�;��AŬ��L2��*֧$D�,�I��~e0�
4D7��fh#
��)ca��JP?�[�S�{`d	)�D ��E��%D�4C@��&>I��E10���	@���3�qʳd0}�RB���d�0W�
�#woVG�9q-��n!򤌾�H�`��#5R8���ُU�& �� a�'ܺ@��X���/C�sq�-J���~�� (7^���)� �qbc�J��h�G-$��"O��dM	8���P�нT�t��$"O���bk��#~�� UjH�r쒌�T"Or��*�C���sO�?+�t���'�-c`` �q�<٪�-�,y`���'~�b�. �u�F�R��Q�%ŊEP�'Ϙ-�3���PJLmq'b�&�RѸ�'stp�h�I�ģ!�7p�x�'@�]s�¹����`��(,h���
�'������/O�-����&7�N��
�'E������ڈ��쌧n|E�	�'���y�@�1��U� iK�w���'��A� y������8�@�'Ԍ��V��J�-����5v��Ъ
�'`��q'��'*�2�[?���
�'W�a �%��Q��I�RȀ�!	�L
�'"\�A�ح!���*/$x0
�'�,��pi[=?(1��U�&]�P{�')��aq/S�.��\������'�*P���ZY��pCGK�J���'�R0z�@˂B�����K�g�N���'S�!��M�h�g�	C]���'���H��m�td��(�73�X�
�'���� ��-|N�r`�((���	�'R�m2q�O,�>�Ap��{��պ�'f<@b��/,���$l��p��:
�'��x�Dݡ:}���Säs��D�'�"���(k"lE�ԅL`�v;�'�i�fJ"u��s7���a����'r��sHu\���v��'eN6Qk
�'TxR�̙�}I�ȧ&W$�f�B	�'ל`(RZQ�(� e;1,D"�'6
y�Q�V�Ee&�zo�6@����
�'Ǣ��� #*�Pq��j���䰱�'�FI��	C�XA��ߟQ���'�x����ɒx ��B �cT���'&蝸u�^4-&�m�b���k58�'��QRW%�- �R�aB%i�,qz�'@>M	�)�y1�� U�rK��p�'�֕H�[_��y ��,�| �'�ź�*̏)��ʂ�N	j`[�'�M���P		���(y��P�'��u��e���1�%qj�K�'7r�k4A�6�ؘ���`� ���'�����P!kH\Ix3�!ӵ�`�<��@��t��n؛S1J�*'�a�<�`�B	e�V�B�Zg��"4Ȕw�<��cǽ+)j%u��|T�.�k�<���B�t�g�Rc�0�d��J�<�rJ��.�f�`��O�( v��K�<1V����0Y
�
�@�X�<�s���;��#�Y2GRס
[�<�%*F���a� 8Y0��gFV�<9$��;�x�� 5?^fA��J�<	F�Lb?Ҽr�P0K�4�Ū�J�<Q�/�� /Ա�� *Xz� ��E�<Y�nʾH���kE��&W�j�Q#\A�<����H�ub�OD	4���'�]t�<9�'43~;a�MWژHGRx�<�J�>k�%YRd�Epp�+@��y�<1���%P�lp�T�ފxX�q��!�~�<�#.��DlH��юAz8��ġ�]�<�`�^<i���1Fi_�a�lL���LM�<A1�O��m��F��,en�M�<� ��H��Ul'j��g�D�Nu�"O6�8ѪvUV�!��W�xb�@&"O0��`F�aq�dW�Mlb9��"OLE2�DݕT�z��J?��dY0"OX[��y�H�qg������s"O`p�0�^'R���p�.4Pz�Q5"O���1&��(^laV�K��ȱ"O���p�Z�R&@%�z=I"O1��XE�z���]�5f{ "O��6�
 I4�u�g�>!�@JA"O�U���T��A(P�H2�z0�"O��^81�w�ş"(Z�*�N�c!�ڨVB��{eM�r/ҸS�L�R�!�$��$��ZfN߮E$��["k�G3!��H�{r��r�C  p(����29	!�$]�w���"��1�����	�!�ą
�|!��!P&(�aC�*�!�ư`yH�#F�n}�uB��T�!�� �ܡS�Ԟ,�~e�DO���!�ḎP	B�K�)�]w�!��i[�y�!��h?�y
$D�*n�c��M�!��΄`����J�-[MRQ)`�ʩw&!�D0T�  Bd%��+7�9@�m�d!��4lv���TV�3ED�[�!�$�}>pڕ�;D�����<�!���&���3%�>��3dnr�!�R�%�`UZU��*馀�c�ǒR4!�͊p��Hc��6e�dUXC
�$-!!�d[:4���p ��� �h�R�	ք8�!��P�J^^ac�H֨X��Aô�^�p�!��	\$��K�\�nd����<�!�$�*&�x@��j
��x���!����jn�]�K��ZU��	B8J!�ڢz��KхY��q���B�!�N�]��za��*m�����j�!�ē�5��p)@�<}�G�!�$����){�J2l\tI���3k!��(����U�ݑrQ^�	���tI!��&M��� �S���a��E�lI!򤌆Lr&K���Y5i�E?!�U7N����&A��͒Ƨ�R/!�$�~�vS'�u����K�,!��*R<m�̏��D����B!�d�;2L1�Ъ�+k4 0��ޔ9�!�dס=�l�B�aK�
tFH�!���	[���d;?�8��cF*g�!�$O#r����E.A����CB��w�!�)Y���`��=B�I�����yF!�$�\�&�b!N�=f |�zT�N�$9fE�%h�*� �s�O`-ى�Y�����y����cƄjg�U9 �"D��F�̣7c5N�r�D=��^�hp�(R�Λ9W�5��Cx��u@ǆ&��-I7-X7_ފ����<��d]�a�~㟰�fL[.l��pB�/ԩ ?n��/
5Y���@A�!l�Ү/�X���'fT�;f!T\�`�:���$}�V�BN<��4{��Uu˙�qX���Z�@!�'���T����S�F1�����y�tM��%��~�%ɤg@]�@�C{
A���\�e�����Z=�,,�'�'L%�yb��l��� �S��0k����i�.�bE��s�(�ړ,J�]d^y�����+U�.�j�M����'W�����E*e��1��l[3W~�ib�)ʍjT(�j�)�![��#E�$3�����2ғ@Ndx�Ä?ym�e%"Q&�F��'���#����6���ܠ����r�X���E�T�	�!��$i���@Y.��\�Q)�&J!�}�&������If�N
��W���bG zd$H�N�QK�F�D�R��/��̵p�
,':�toG��(�;o�q�h�]F̜���
l���� @d���ݾ	��h�&̖�U�^]�pFǦI��p	l�n�n�jhH�$�?�t�V֠T��d��N��oڗ:�`8���8Y���Q��"�Z�>����V\��e��*�ʀb�e>� p<�U�P5Y�H���a۩kD� !e`ƁY&I�u�����植Vr4�Bt�'�XY#�Q�^Œb�o�)`1 ui�'����к}fD��(J r����'$���S*X�@_�K%��b����)ބ4ľ��G�+4����*��E@�1
�@R)�2~��b��<��Kc��%��$oZ]H<aJ�����Rg����d�5}�	�zY
5ϛ����D��Q������{[��DȕW��@$��8�'�	O�R����C�ta� 
�y��'���|jPǅ�9�X����V
>�x��Nt���K҅�
/���3=O�a�E�/R�[��{<Y�"OF��牓o�PQd�جu��0�@�DV�HZ�]P
�7����a�"9��c҄�'}���[r"O�e�Q��""���Y'L��c~A[�E7 %*J>Q��>Q���305��u�@-�`�pcQN�<!`� Baj��M�#:p���c�ğ24�֮0�a}��� q��"�!@�e��2E���yRg��E֊%�ME�Z`d���(�(�y",ت����S��F�pԩ�y���<Lt�a��%���r�Z�0�y��*v���WN�t��r�A��y�E��X�9�NT�%� �1����yR����\��i�d���`a��y�Ɖ<��{
�P�����ӕ�y�&J�#�v<:c�J,6U#�
M��y(�&�&9��V�`z`o�y���`��H'N�B�:)�FfQ(�y�I�c�6���Fٺp�'Π�y�ɿ�∺"C�J��d�6/��C�I>XO`��$��}��U�R�
"?R�B��1<��u��|�!�竈�zkhB�I�*�+�B-lr�a(�&HZB�I/	]�����N�yb �OB��$E
MF��شX%�xY'N�p�h�dXr��܅ȓa���I�� WLR9����
n��EzB�ȱA��4Q�S�0���qDE��}0��a���$|r�B�ɓ0e�1�^�Fa�g��-־<s\!��=9�M4}���'�H�@@���S�����%r�-s
�'���˄ּ����R������'��-p������Մ�ə7~Tj�$TJ��E{Ⱦ?^4���	�#��H��ͅ��ر� �K�`�b�	-�0(�'��D�<� f��6�0q���DS�I��W����f�Zs�5R� M���ٛE$@���"O��B�˘8�0��i��U���b�����'��}�O?��T$1��!q�T�"�ވ�b�1z�!�d�x�8 
�ˬiX�ؐ`AY�Bh�DQ!Tre���0=A�)��q[�mM)Y�����i8�`q�f�9m�\i�+	�6�`�B��\:���;��U�`4!�ğ-#�,�1�W��*��`j�m���lۤo֐z��D��W2~5X$ۙk��Ժt�1�ym�G�:�dޱZ������?1P�٠I��"~:�J����M��#�I�Pر��D��yBdZ	Y �A��Ӻ@��ŉUJ߸�y�F�|�T�) ���By��VBA�/n �Чj%�W��~"�ߜ0�L�r癱>�
��O�6�y��A�}��p�5:�p���L.�MC�oB�QU��L�w.T��:|4�ߗN�@���ɣ
؇e8,�� �ii�V��ɓ���iz!���Sxj���Y�/�XݠW`�hnqOj����62b�ҋ�I�$P���p��O�d嚐+0I�0!�K��V "���7)�xQ�D��� i���*ģ`�4Dܢ|�'��A87��:B�X���3k t��'9L�7kR�|�٣u.�c����Ŀx�>y�`�<�0>1/]R�Ba1��T�/�j���EZ�����
�\��!P�6O��2�j��j����W���3͈���"O��������\2�Ǐ�h� Ās��U5nv�iE�爟�L(p@�,b2���æ�$�VA!p"O� P�"�
�:P.�*��0i��\ʢ�ծq�̹S�>���7�gy�(I�$�^�p+A'<@`��!�y"�ʨښ�#���X�'�@��M���!s,�t$FhuC �n���O�N����Ɏ��,��_��[���%H���B�4'���Uk D�l���/Y\x��`·�:��YA�j!D��90�O&�:�+d��7
�H���c8D���E�b�L:�HuУ� v�C�Ɉ0ET�yFM_�k�X1��"ū/�B�	jk$c���R���K4�W��B�	����D�!���e@MmLC�I��x|�"E��/��U���N_�B�I�mАM�šؐF��x�M
�]�B�I�P-6��P���=��$"D�
�b	�C䉬U��p3�ʚiO�x�Q�F"UC�I/T�b�k�_tv��a�	B<�B�{�F|p��iYpPXroɷ<�B�	"
���"m�#s^��1��!a�B�I_�D)��Ѧ<�|��E�!w��B�	���1�G��"^s�ـ`F�-��B�I�y&.l2"���b`�+i�B䉓e�1�_#EP	�R�zK�C��#Y��h5�E*!<���4��4�C�ɱG_�Ixg ɐ:���l�=F�C�ɟq����I*F�l�U��,fm�B��2e�Pq�b�;~1�a;��ͬ���'���� '[ZX�u�)վ��'}��ˢ�R�)|���.�!ui�!�'���Y���r�M�B�/w����'����L�Y��kPc��p�Y�'â�3��^$W�8�{������'�s�.�2FnĘF��`��x�'��y�B$I�n<�CΘ�X/ ��
�'F� 	̉

@�+�*|v���')�T9r@�&)�3�ݱ1w�%��'�l�!h֖l<���a�\�����'�)��X���af�*y�6��
�'3�q+�@�F�	)@,܋fg�z�'��:�P�Xcи�G��$j�v��'�H�:`%��Ai ⠙�*�r���dE.!SE��UĦРcE"/+�Ňȓ7�;��X�X����O�j%���48����~��;6��#��)�ȓe?�E�F�~aTA{f��z����*o�͑��������wO�b1�}�↜ynJ}��O��!΋�kc,����3p�@���C�;��-�&�/;�~5�'�����O($��4�|����GR��и�i�䘖'�8X�����9O�$�oՊ];D� W /�J�?OT�Х�i�b�"~P�����.� Pch4	���=4����j}R�	 ���𩓄V��㲋F�Q�Υi#K�L����>�6S�`�S�O�2��Y{^��&&UW*%��O���"���1��Y}>�9��)�2-i�d5L���K�F�>1�I	�<Q��O�dD�ț'/b0�c�AB�XB$��C��.�M��eL�<� �O���1��O����]e�3c뛳[��Ir�)v>\�=����Ć�y}�H����(:���A1!�dߐ-�d95����u��Nr!�>*�D��I������!� �d�����;�|��f���+�!��8�郣�O�y^���U�)@!�D�=`�|js��W�X�
��>a{��D�I��u�d@S
\��	�C;Z&�L�>�1�]��y��˅n�"Pc����wk0��6��<��wj2�<�Ou�����;�&��h|��	`aHN�}�\�'��oڡ9��A{��O��=��.ΐ�b����πEܼ98�O� ��=/|(���}לXb�o�D��E=}p�����tt\%��l�,\�$��'�O,�@W�5��E�� X�@�@n�`l�c�:?	�)�Ӡ��Tƴ��=Od��� �2:a��KSS� �&&����/_���9�'njdj�K�{��� çf7�1h�C1ܪ�@��_46��V2�Ѝڋ]�QH�A�>f6�5ԧ�O�P�梏�E����gA�fX�X�(����0;�����0|�a���B��T��d����c �g�<����>F��RF����X�PWd�<�i�	]<ȸ��ڟE�dXsc�a�<y7�3���xLKarFez%W�<y�nU��(�E�@�f�*PE�R�<	u,�	C	��W�vnu��C�<ɣ�S4uZju��@�$ӜH�r��I�<��C�C��k7�IGY�(0A��l�<scG1d\���Iռ>��{lj�<��lG�6�
)"��= ��CsK�z�<I����Rҥ���6Ɔ����r�<Y&��TTi�&��E���m�<p�=/�����imU�c��B�<9��Z�R�����
b7f��
Oy�<!6(Կn+b����^F1��}�<!�̕E� XE&τ Hn�3dk[v�<�5��H�F��f�"s �sg�i�<���C7O�p	ǩ���P��)�[�<��K'^��}b�܏�i
�@�<Q�L^/.;���bH_��XB��Nu�<��AX��~��O�%������r�<I��^����o@�(*�q�<	 <x��]Q��X)���Z��Pl�<Iu��>@����B���AĔ'k�^Q��v�,!�!�`�8�!F�z2��ȓf��L1e)Os��d�4���B��Ɇȓ3Z���PoM�U�>�`��E&7��x�ȓ;Ό�/)p˒THGN��{!�d�ȓq�TAJ�"� C��d�
���(�ȓ0V,\ ǋV+l��K�#8�4��-J0���j���ـ'��5 ��ȓ�T�� Gv��֬��m2�1�ȓ
�ґyfF�<@��E�ƃM�ل�>X|[惉w��|�R9"t��ʓ-��$�5�]�*��a U@�=l<B�I0\v��C��Q�(PaaO��k4B�I�Tq��� ž<�α�P��,�C�I�q�\@�F�^1h܄}b�)��C�I�,e����$\+����AX<E��C�ɢN���!�Z�7m����U�JP�B�	�_�8`�����@1!�Q7^o�C䉔Y�就��.wz��	"�˚X�C��6AĒ��S&%���1�ɞ-<�C��<���vg˖�@L���	-g"�C�3z����&�#.02�ٲ��2ӾC�I�*�f�Btf	%^LZq�fJB(n��C��Tl>�Ѕf� 0=����D�W�*B�I1ǚ����Քv�d��ᎃ 1�C�	�.��)�L�'X�.��L �3Z�C䉩Y������zW ���${��C��E_&�	���?Ȣ	��hϦ>�C�I�t�օ�&��&l����3��ϾB�	"p!���%�lK��]�>k�C�	=j#��Y�cߊU� =����ed�C�ɦ|��������@�"h.B�I.3� b@��s��&O�o�B�Ƀߞ�� �"2�bqbmW'fj�B�I�V��a��$F%g䎌"�!Q |�B��(q�,8j�"�9i�R��J�;WTB�� <�d���&� �6�b���EfB�)� �0�+��E��䡅��E2�y��"Oj��g�M,�`٣F�!\L�q"O��p���תrBM�	.�ı�XD�<���N�	���*���~���2*T}�<��G�)/�:H(�j�({���r�d�<	�Ā0$����bӪj����iM_�<1���.a
�zQ���=���/D�8�G���/yt-Іm�Ɛ�#�.D��"Q���YiD��:9HzC�,D�tłʖ%u<��U'�/tVX8��5D��#ցOI�ƘH�ֳ:ɦ�3�2D�TH�lD"�ʬIN(!z����2D��z A?6;�$�e��(&�V/h�JB�	�Ԭ����*�\ɢ@@�hC�ɡ��ҡ�Ɂ`<5`s�T�Y�~B�I7e׀��E߮L"��s�"nwB�ɶX���� �8R��T��+T_Q�C�	{"�kQD���n5���M{z8B�	>W�VM�)	����"!
8RjB�I96=j5BdJ�i��ݒ!O���nB�pV���c�L~�	�䊚�b�C�	�f�@:���M��	j�a��s��B�I�	.-A�E�Iz2	!T�/^��C�IEؔ��]�yc!��+��{i�C��*_���D�EO�d���R�zC�	�f*�	e�š5��l�"���~$lC�	E�����KL�9�`����9,��B�I�8�HDKt��e�z肠�1W��B�I%��5b�! ��7 Y�5��B䉙�z� �D��VpY�k��P��B䉌�	ҖmQn��Q�0h�e�rB�ɹ����(�[��@eH0�B�I�{��$[&'!�=�`B�yH2C�ɺk��E��Z�j8��%�S+�bC�	8$�d��ի�&�-S���wD�C��:(%v}s��S�@���]�ZC�;W�ҙ�Q�7k��ٳD>pD0C�I�(_ZDJ�b.X���R��lDB�I{�4�eKG&6�U��k׫I	�C�	%�@�%e�W�D̫r%֦O�C��SqV�y�ۣ�>�EoUV�C�	jp�l���Y[�&<)ϓ�V��C䉽mr�xP*O.S��\��D�C䉲3�����@W2N�K"/��2FB䉒\+ �+Sg�9-��=*�A��7jC䉇
�z���%q������ JrjB䉉r�`%R
4j	`�/�
@"OX)���=� M+bꁈ}�hB"ORPw����1w靲DUFl�P"O�U�ĥZ�}�0p�5��?{p�"O䰋��w��4�)�7A���{f"O"�c�F�N��5�$;�}K�"Ov� v͆M��Wꔖ|��x��"O�`$ɎbB�P1,��<��EsW"OFTcB�?�Ê�>��|"W"O�LC��?e�$��HW�HR���"O~��G(��gA�\�c��"<9�Y�e"O�	��ź�ڬ(����)+���""O|}�SM̒e��2�D�$�3�"OƍqHΰ��!�d_?n40�G"O����V�-=���a���g"O�� ��G�"�1+݆%��|r�"ODU�@�ܒ�h�"!��B����7"O6��`#�� %`0����b��"O� X8r3 4��[	��F"�Z"O������
릈KG>06�f"Od��r��=_�E����/!�n�"O�E�,\�y�D�𐢛c^��#w"Oެ�U� ���(֦&u�X�$"O�%��a�4�AE�[e�Cg"OԉrS	Uhu��@��\�yU� x�"Oʱ����*�Lx#`���C&@I	�"O���P�6
x�	��W7&�y�"O><x��J�� �kK>)} K�"O�d9�DS�buXQ���2�f���"ON|�d�V�l|A�_06w\��"O*Ey�)kq��k���q�� *�"O� ����\>�	�$E�w�h @"O*�B�(�,|2��P�M�_?�=�q"O�x�˗5GUl��]4)P�4�F"O$���&C^�$�8vGә6N"�AP"O:݉��M9UK��!Ǚ�O1�ب�"Ob)ҵF�&������9D��T"O.e;�� TbɈѨK �)�"O�UC�]�5�ݱeB�#*���q"OX��VV�^�>EhL�>�A�1"O\���U�q��)3*�2-�P�Ac"Ob��G���p�\�1���s"O�I���6K�<�C #Ĺs�~0�"O��2V�ƵI�����W,c	\�"O0�J�e"��:"L���L-�"OB�"V�Ѣ*���T�D8-Tb�y�"O��8���_�!�B�95ڽk0"OD�E�\�7�-�����zYia"O�Pr@�q���戒����"Ol|��#[�xl���8s.y`�"Ot��)�?����G3"Z�a"ODL��*��6E3(Q&�B�s"O��gF�"vT��㦇@0G�5�"OL���B�E^�3�F��6T+�"OI3-��3�lңO׿"[�����pK�s��>?�x�# �(.�dمȓ3�(��]*M�:�:��#`A<���"����B���K��m:4�%n��9���u���)�rX�&Cػ;Ӳ����B &(W��h�ץ��`�>���N��d1��],!��r��j!�C��#]
��噤'�*��g��0�DC�ə �aSE� �0��zFG�7�^C�I>0H4��l�G�ɓ��%hVC�	�f!b�J�q�T�t剃&� C�7N�xAC�ZYك�I�H�B�	���� /]�n�"�rQF�#X*�C䉭0O� k�AT�N�M��(Q
�C��׈=jB!�/�����:��B�I�!U�:�a����C���w2�B�ɺp��A&� V��P( @]0B�I <_�C�
8����B'b�&B�I�p��1���0�fw�x�"O�$�[y�5�O��]2�1�"O�@7`A�e��� \�zM�c�"O
�yWN4�J(25���uD�q�#"O����D�&6�����\�%>���"O-�V����`���j�$8<��"OV)J�I n��*s��+�,)�"O0��� ���p�3/dB���"O"ݱ�)Ǡq�ȑ�a��	iy2��q"O�1�u�Q�p�.��֊֐#�<�k�"O� ���A̫y�$"��D�C��HYq"OH,��8m^2�qb
�W�\L17"O~���LX%,���2iȀc��,
A"O�(;ag�;-36!�脌_~�q�A"ODiN+zS���"W�વ"Oy!S'� 5�T�����,K�-zv"OP�#!\*Ƽ�f�ߧ �,��"O
aP&��%��ʞ�I,���B"O�`@�c݉��(dJћ!�|0�"OV���   �